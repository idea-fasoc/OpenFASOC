* NGSPICE file created from diff_pair_sample_0254.ext - technology: sky130A

.subckt diff_pair_sample_0254 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X1 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0.11055 ps=1 w=0.67 l=3.31
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0 ps=0 w=0.67 l=3.31
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0 ps=0 w=0.67 l=3.31
X4 VTAIL.t14 VP.t1 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X5 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X6 VDD1.t2 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.2613 ps=2.12 w=0.67 l=3.31
X7 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.2613 ps=2.12 w=0.67 l=3.31
X8 VTAIL.t7 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X9 VTAIL.t5 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X10 VDD2.t2 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X11 VTAIL.t6 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0.11055 ps=1 w=0.67 l=3.31
X12 VDD1.t0 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0 ps=0 w=0.67 l=3.31
X14 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.2613 ps=2.12 w=0.67 l=3.31
X15 VTAIL.t11 VP.t4 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0.11055 ps=1 w=0.67 l=3.31
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0 ps=0 w=0.67 l=3.31
X17 VDD1.t5 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.2613 ps=2.12 w=0.67 l=3.31
X18 VDD1.t3 VP.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.11055 pd=1 as=0.11055 ps=1 w=0.67 l=3.31
X19 VTAIL.t8 VP.t7 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2613 pd=2.12 as=0.11055 ps=1 w=0.67 l=3.31
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n48 VP.n12 79.7913
R38 VP.n84 VP.n0 79.7913
R39 VP.n47 VP.n13 79.7913
R40 VP.n23 VP.n22 71.1565
R41 VP.n65 VP.n6 56.5193
R42 VP.n28 VP.n19 56.5193
R43 VP.n56 VP.n10 51.1773
R44 VP.n76 VP.n2 51.1773
R45 VP.n39 VP.n15 51.1773
R46 VP.n48 VP.n47 45.6811
R47 VP.n23 VP.t4 37.0501
R48 VP.n52 VP.n10 29.8095
R49 VP.n80 VP.n2 29.8095
R50 VP.n43 VP.n15 29.8095
R51 VP.n51 VP.n50 24.4675
R52 VP.n52 VP.n51 24.4675
R53 VP.n57 VP.n56 24.4675
R54 VP.n59 VP.n57 24.4675
R55 VP.n63 VP.n8 24.4675
R56 VP.n64 VP.n63 24.4675
R57 VP.n65 VP.n64 24.4675
R58 VP.n69 VP.n6 24.4675
R59 VP.n70 VP.n69 24.4675
R60 VP.n71 VP.n70 24.4675
R61 VP.n75 VP.n74 24.4675
R62 VP.n76 VP.n75 24.4675
R63 VP.n81 VP.n80 24.4675
R64 VP.n82 VP.n81 24.4675
R65 VP.n44 VP.n43 24.4675
R66 VP.n45 VP.n44 24.4675
R67 VP.n32 VP.n19 24.4675
R68 VP.n33 VP.n32 24.4675
R69 VP.n34 VP.n33 24.4675
R70 VP.n38 VP.n37 24.4675
R71 VP.n39 VP.n38 24.4675
R72 VP.n26 VP.n21 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n59 VP.n58 21.0421
R76 VP.n74 VP.n4 21.0421
R77 VP.n37 VP.n17 21.0421
R78 VP.n50 VP.n12 10.2766
R79 VP.n82 VP.n0 10.2766
R80 VP.n45 VP.n13 10.2766
R81 VP.n12 VP.t7 4.87875
R82 VP.n58 VP.t6 4.87875
R83 VP.n4 VP.t1 4.87875
R84 VP.n0 VP.t2 4.87875
R85 VP.n13 VP.t5 4.87875
R86 VP.n17 VP.t0 4.87875
R87 VP.n22 VP.t3 4.87875
R88 VP.n24 VP.n23 4.39145
R89 VP.n58 VP.n8 3.42588
R90 VP.n71 VP.n4 3.42588
R91 VP.n34 VP.n17 3.42588
R92 VP.n22 VP.n21 3.42588
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VDD1 VDD1.n0 236.849
R133 VDD1.n3 VDD1.n2 236.736
R134 VDD1.n3 VDD1.n1 236.736
R135 VDD1.n5 VDD1.n4 235.221
R136 VDD1.n5 VDD1.n3 38.9966
R137 VDD1.n4 VDD1.t7 29.5527
R138 VDD1.n4 VDD1.t5 29.5527
R139 VDD1.n0 VDD1.t1 29.5527
R140 VDD1.n0 VDD1.t0 29.5527
R141 VDD1.n2 VDD1.t4 29.5527
R142 VDD1.n2 VDD1.t2 29.5527
R143 VDD1.n1 VDD1.t6 29.5527
R144 VDD1.n1 VDD1.t3 29.5527
R145 VDD1 VDD1.n5 1.51128
R146 VTAIL.n15 VTAIL.t1 248.095
R147 VTAIL.n2 VTAIL.t6 248.095
R148 VTAIL.n3 VTAIL.t13 248.095
R149 VTAIL.n6 VTAIL.t8 248.095
R150 VTAIL.n14 VTAIL.t10 248.095
R151 VTAIL.n11 VTAIL.t11 248.095
R152 VTAIL.n10 VTAIL.t0 248.095
R153 VTAIL.n7 VTAIL.t3 248.095
R154 VTAIL.n1 VTAIL.n0 218.542
R155 VTAIL.n5 VTAIL.n4 218.542
R156 VTAIL.n13 VTAIL.n12 218.542
R157 VTAIL.n9 VTAIL.n8 218.542
R158 VTAIL.n0 VTAIL.t4 29.5527
R159 VTAIL.n0 VTAIL.t5 29.5527
R160 VTAIL.n4 VTAIL.t9 29.5527
R161 VTAIL.n4 VTAIL.t14 29.5527
R162 VTAIL.n12 VTAIL.t12 29.5527
R163 VTAIL.n12 VTAIL.t15 29.5527
R164 VTAIL.n8 VTAIL.t2 29.5527
R165 VTAIL.n8 VTAIL.t7 29.5527
R166 VTAIL.n15 VTAIL.n14 16.0824
R167 VTAIL.n7 VTAIL.n6 16.0824
R168 VTAIL.n9 VTAIL.n7 3.13843
R169 VTAIL.n10 VTAIL.n9 3.13843
R170 VTAIL.n13 VTAIL.n11 3.13843
R171 VTAIL.n14 VTAIL.n13 3.13843
R172 VTAIL.n6 VTAIL.n5 3.13843
R173 VTAIL.n5 VTAIL.n3 3.13843
R174 VTAIL.n2 VTAIL.n1 3.13843
R175 VTAIL VTAIL.n15 3.08024
R176 VTAIL.n11 VTAIL.n10 0.470328
R177 VTAIL.n3 VTAIL.n2 0.470328
R178 VTAIL VTAIL.n1 0.0586897
R179 B.n634 B.n633 585
R180 B.n180 B.n125 585
R181 B.n179 B.n178 585
R182 B.n177 B.n176 585
R183 B.n175 B.n174 585
R184 B.n173 B.n172 585
R185 B.n171 B.n170 585
R186 B.n169 B.n168 585
R187 B.n167 B.n166 585
R188 B.n165 B.n164 585
R189 B.n163 B.n162 585
R190 B.n161 B.n160 585
R191 B.n159 B.n158 585
R192 B.n157 B.n156 585
R193 B.n155 B.n154 585
R194 B.n153 B.n152 585
R195 B.n151 B.n150 585
R196 B.n149 B.n148 585
R197 B.n147 B.n146 585
R198 B.n145 B.n144 585
R199 B.n143 B.n142 585
R200 B.n141 B.n140 585
R201 B.n139 B.n138 585
R202 B.n137 B.n136 585
R203 B.n135 B.n134 585
R204 B.n133 B.n132 585
R205 B.n632 B.n112 585
R206 B.n637 B.n112 585
R207 B.n631 B.n111 585
R208 B.n638 B.n111 585
R209 B.n630 B.n629 585
R210 B.n629 B.n107 585
R211 B.n628 B.n106 585
R212 B.n644 B.n106 585
R213 B.n627 B.n105 585
R214 B.n645 B.n105 585
R215 B.n626 B.n104 585
R216 B.n646 B.n104 585
R217 B.n625 B.n624 585
R218 B.n624 B.n100 585
R219 B.n623 B.n99 585
R220 B.n652 B.n99 585
R221 B.n622 B.n98 585
R222 B.n653 B.n98 585
R223 B.n621 B.n97 585
R224 B.n654 B.n97 585
R225 B.n620 B.n619 585
R226 B.n619 B.n93 585
R227 B.n618 B.n92 585
R228 B.n660 B.n92 585
R229 B.n617 B.n91 585
R230 B.n661 B.n91 585
R231 B.n616 B.n90 585
R232 B.n662 B.n90 585
R233 B.n615 B.n614 585
R234 B.n614 B.n86 585
R235 B.n613 B.n85 585
R236 B.n668 B.n85 585
R237 B.n612 B.n84 585
R238 B.n669 B.n84 585
R239 B.n611 B.n83 585
R240 B.n670 B.n83 585
R241 B.n610 B.n609 585
R242 B.n609 B.n79 585
R243 B.n608 B.n78 585
R244 B.n676 B.n78 585
R245 B.n607 B.n77 585
R246 B.n677 B.n77 585
R247 B.n606 B.n76 585
R248 B.n678 B.n76 585
R249 B.n605 B.n604 585
R250 B.n604 B.n75 585
R251 B.n603 B.n71 585
R252 B.n684 B.n71 585
R253 B.n602 B.n70 585
R254 B.n685 B.n70 585
R255 B.n601 B.n69 585
R256 B.n686 B.n69 585
R257 B.n600 B.n599 585
R258 B.n599 B.n65 585
R259 B.n598 B.n64 585
R260 B.n692 B.n64 585
R261 B.n597 B.n63 585
R262 B.n693 B.n63 585
R263 B.n596 B.n62 585
R264 B.n694 B.n62 585
R265 B.n595 B.n594 585
R266 B.n594 B.n58 585
R267 B.n593 B.n57 585
R268 B.n700 B.n57 585
R269 B.n592 B.n56 585
R270 B.n701 B.n56 585
R271 B.n591 B.n55 585
R272 B.n702 B.n55 585
R273 B.n590 B.n589 585
R274 B.n589 B.n51 585
R275 B.n588 B.n50 585
R276 B.n708 B.n50 585
R277 B.n587 B.n49 585
R278 B.n709 B.n49 585
R279 B.n586 B.n48 585
R280 B.n710 B.n48 585
R281 B.n585 B.n584 585
R282 B.n584 B.n44 585
R283 B.n583 B.n43 585
R284 B.n716 B.n43 585
R285 B.n582 B.n42 585
R286 B.n717 B.n42 585
R287 B.n581 B.n41 585
R288 B.n718 B.n41 585
R289 B.n580 B.n579 585
R290 B.n579 B.n37 585
R291 B.n578 B.n36 585
R292 B.n724 B.n36 585
R293 B.n577 B.n35 585
R294 B.n725 B.n35 585
R295 B.n576 B.n34 585
R296 B.n726 B.n34 585
R297 B.n575 B.n574 585
R298 B.n574 B.n30 585
R299 B.n573 B.n29 585
R300 B.n732 B.n29 585
R301 B.n572 B.n28 585
R302 B.n733 B.n28 585
R303 B.n571 B.n27 585
R304 B.n734 B.n27 585
R305 B.n570 B.n569 585
R306 B.n569 B.n23 585
R307 B.n568 B.n22 585
R308 B.n740 B.n22 585
R309 B.n567 B.n21 585
R310 B.n741 B.n21 585
R311 B.n566 B.n20 585
R312 B.n742 B.n20 585
R313 B.n565 B.n564 585
R314 B.n564 B.n19 585
R315 B.n563 B.n15 585
R316 B.n748 B.n15 585
R317 B.n562 B.n14 585
R318 B.n749 B.n14 585
R319 B.n561 B.n13 585
R320 B.n750 B.n13 585
R321 B.n560 B.n559 585
R322 B.n559 B.n12 585
R323 B.n558 B.n557 585
R324 B.n558 B.n8 585
R325 B.n556 B.n7 585
R326 B.n757 B.n7 585
R327 B.n555 B.n6 585
R328 B.n758 B.n6 585
R329 B.n554 B.n5 585
R330 B.n759 B.n5 585
R331 B.n553 B.n552 585
R332 B.n552 B.n4 585
R333 B.n551 B.n181 585
R334 B.n551 B.n550 585
R335 B.n541 B.n182 585
R336 B.n183 B.n182 585
R337 B.n543 B.n542 585
R338 B.n544 B.n543 585
R339 B.n540 B.n188 585
R340 B.n188 B.n187 585
R341 B.n539 B.n538 585
R342 B.n538 B.n537 585
R343 B.n190 B.n189 585
R344 B.n530 B.n190 585
R345 B.n529 B.n528 585
R346 B.n531 B.n529 585
R347 B.n527 B.n195 585
R348 B.n195 B.n194 585
R349 B.n526 B.n525 585
R350 B.n525 B.n524 585
R351 B.n197 B.n196 585
R352 B.n198 B.n197 585
R353 B.n517 B.n516 585
R354 B.n518 B.n517 585
R355 B.n515 B.n203 585
R356 B.n203 B.n202 585
R357 B.n514 B.n513 585
R358 B.n513 B.n512 585
R359 B.n205 B.n204 585
R360 B.n206 B.n205 585
R361 B.n505 B.n504 585
R362 B.n506 B.n505 585
R363 B.n503 B.n211 585
R364 B.n211 B.n210 585
R365 B.n502 B.n501 585
R366 B.n501 B.n500 585
R367 B.n213 B.n212 585
R368 B.n214 B.n213 585
R369 B.n493 B.n492 585
R370 B.n494 B.n493 585
R371 B.n491 B.n219 585
R372 B.n219 B.n218 585
R373 B.n490 B.n489 585
R374 B.n489 B.n488 585
R375 B.n221 B.n220 585
R376 B.n222 B.n221 585
R377 B.n481 B.n480 585
R378 B.n482 B.n481 585
R379 B.n479 B.n227 585
R380 B.n227 B.n226 585
R381 B.n478 B.n477 585
R382 B.n477 B.n476 585
R383 B.n229 B.n228 585
R384 B.n230 B.n229 585
R385 B.n469 B.n468 585
R386 B.n470 B.n469 585
R387 B.n467 B.n235 585
R388 B.n235 B.n234 585
R389 B.n466 B.n465 585
R390 B.n465 B.n464 585
R391 B.n237 B.n236 585
R392 B.n238 B.n237 585
R393 B.n457 B.n456 585
R394 B.n458 B.n457 585
R395 B.n455 B.n243 585
R396 B.n243 B.n242 585
R397 B.n454 B.n453 585
R398 B.n453 B.n452 585
R399 B.n245 B.n244 585
R400 B.n246 B.n245 585
R401 B.n445 B.n444 585
R402 B.n446 B.n445 585
R403 B.n443 B.n251 585
R404 B.n251 B.n250 585
R405 B.n442 B.n441 585
R406 B.n441 B.n440 585
R407 B.n253 B.n252 585
R408 B.n433 B.n253 585
R409 B.n432 B.n431 585
R410 B.n434 B.n432 585
R411 B.n430 B.n258 585
R412 B.n258 B.n257 585
R413 B.n429 B.n428 585
R414 B.n428 B.n427 585
R415 B.n260 B.n259 585
R416 B.n261 B.n260 585
R417 B.n420 B.n419 585
R418 B.n421 B.n420 585
R419 B.n418 B.n266 585
R420 B.n266 B.n265 585
R421 B.n417 B.n416 585
R422 B.n416 B.n415 585
R423 B.n268 B.n267 585
R424 B.n269 B.n268 585
R425 B.n408 B.n407 585
R426 B.n409 B.n408 585
R427 B.n406 B.n274 585
R428 B.n274 B.n273 585
R429 B.n405 B.n404 585
R430 B.n404 B.n403 585
R431 B.n276 B.n275 585
R432 B.n277 B.n276 585
R433 B.n396 B.n395 585
R434 B.n397 B.n396 585
R435 B.n394 B.n281 585
R436 B.n285 B.n281 585
R437 B.n393 B.n392 585
R438 B.n392 B.n391 585
R439 B.n283 B.n282 585
R440 B.n284 B.n283 585
R441 B.n384 B.n383 585
R442 B.n385 B.n384 585
R443 B.n382 B.n290 585
R444 B.n290 B.n289 585
R445 B.n381 B.n380 585
R446 B.n380 B.n379 585
R447 B.n292 B.n291 585
R448 B.n293 B.n292 585
R449 B.n372 B.n371 585
R450 B.n373 B.n372 585
R451 B.n370 B.n298 585
R452 B.n298 B.n297 585
R453 B.n365 B.n364 585
R454 B.n363 B.n313 585
R455 B.n362 B.n312 585
R456 B.n367 B.n312 585
R457 B.n361 B.n360 585
R458 B.n359 B.n358 585
R459 B.n357 B.n356 585
R460 B.n355 B.n354 585
R461 B.n353 B.n352 585
R462 B.n350 B.n349 585
R463 B.n348 B.n347 585
R464 B.n346 B.n345 585
R465 B.n344 B.n343 585
R466 B.n342 B.n341 585
R467 B.n340 B.n339 585
R468 B.n338 B.n337 585
R469 B.n336 B.n335 585
R470 B.n334 B.n333 585
R471 B.n332 B.n331 585
R472 B.n329 B.n328 585
R473 B.n327 B.n326 585
R474 B.n325 B.n324 585
R475 B.n323 B.n322 585
R476 B.n321 B.n320 585
R477 B.n319 B.n318 585
R478 B.n300 B.n299 585
R479 B.n369 B.n368 585
R480 B.n368 B.n367 585
R481 B.n296 B.n295 585
R482 B.n297 B.n296 585
R483 B.n375 B.n374 585
R484 B.n374 B.n373 585
R485 B.n376 B.n294 585
R486 B.n294 B.n293 585
R487 B.n378 B.n377 585
R488 B.n379 B.n378 585
R489 B.n288 B.n287 585
R490 B.n289 B.n288 585
R491 B.n387 B.n386 585
R492 B.n386 B.n385 585
R493 B.n388 B.n286 585
R494 B.n286 B.n284 585
R495 B.n390 B.n389 585
R496 B.n391 B.n390 585
R497 B.n280 B.n279 585
R498 B.n285 B.n280 585
R499 B.n399 B.n398 585
R500 B.n398 B.n397 585
R501 B.n400 B.n278 585
R502 B.n278 B.n277 585
R503 B.n402 B.n401 585
R504 B.n403 B.n402 585
R505 B.n272 B.n271 585
R506 B.n273 B.n272 585
R507 B.n411 B.n410 585
R508 B.n410 B.n409 585
R509 B.n412 B.n270 585
R510 B.n270 B.n269 585
R511 B.n414 B.n413 585
R512 B.n415 B.n414 585
R513 B.n264 B.n263 585
R514 B.n265 B.n264 585
R515 B.n423 B.n422 585
R516 B.n422 B.n421 585
R517 B.n424 B.n262 585
R518 B.n262 B.n261 585
R519 B.n426 B.n425 585
R520 B.n427 B.n426 585
R521 B.n256 B.n255 585
R522 B.n257 B.n256 585
R523 B.n436 B.n435 585
R524 B.n435 B.n434 585
R525 B.n437 B.n254 585
R526 B.n433 B.n254 585
R527 B.n439 B.n438 585
R528 B.n440 B.n439 585
R529 B.n249 B.n248 585
R530 B.n250 B.n249 585
R531 B.n448 B.n447 585
R532 B.n447 B.n446 585
R533 B.n449 B.n247 585
R534 B.n247 B.n246 585
R535 B.n451 B.n450 585
R536 B.n452 B.n451 585
R537 B.n241 B.n240 585
R538 B.n242 B.n241 585
R539 B.n460 B.n459 585
R540 B.n459 B.n458 585
R541 B.n461 B.n239 585
R542 B.n239 B.n238 585
R543 B.n463 B.n462 585
R544 B.n464 B.n463 585
R545 B.n233 B.n232 585
R546 B.n234 B.n233 585
R547 B.n472 B.n471 585
R548 B.n471 B.n470 585
R549 B.n473 B.n231 585
R550 B.n231 B.n230 585
R551 B.n475 B.n474 585
R552 B.n476 B.n475 585
R553 B.n225 B.n224 585
R554 B.n226 B.n225 585
R555 B.n484 B.n483 585
R556 B.n483 B.n482 585
R557 B.n485 B.n223 585
R558 B.n223 B.n222 585
R559 B.n487 B.n486 585
R560 B.n488 B.n487 585
R561 B.n217 B.n216 585
R562 B.n218 B.n217 585
R563 B.n496 B.n495 585
R564 B.n495 B.n494 585
R565 B.n497 B.n215 585
R566 B.n215 B.n214 585
R567 B.n499 B.n498 585
R568 B.n500 B.n499 585
R569 B.n209 B.n208 585
R570 B.n210 B.n209 585
R571 B.n508 B.n507 585
R572 B.n507 B.n506 585
R573 B.n509 B.n207 585
R574 B.n207 B.n206 585
R575 B.n511 B.n510 585
R576 B.n512 B.n511 585
R577 B.n201 B.n200 585
R578 B.n202 B.n201 585
R579 B.n520 B.n519 585
R580 B.n519 B.n518 585
R581 B.n521 B.n199 585
R582 B.n199 B.n198 585
R583 B.n523 B.n522 585
R584 B.n524 B.n523 585
R585 B.n193 B.n192 585
R586 B.n194 B.n193 585
R587 B.n533 B.n532 585
R588 B.n532 B.n531 585
R589 B.n534 B.n191 585
R590 B.n530 B.n191 585
R591 B.n536 B.n535 585
R592 B.n537 B.n536 585
R593 B.n186 B.n185 585
R594 B.n187 B.n186 585
R595 B.n546 B.n545 585
R596 B.n545 B.n544 585
R597 B.n547 B.n184 585
R598 B.n184 B.n183 585
R599 B.n549 B.n548 585
R600 B.n550 B.n549 585
R601 B.n3 B.n0 585
R602 B.n4 B.n3 585
R603 B.n756 B.n1 585
R604 B.n757 B.n756 585
R605 B.n755 B.n754 585
R606 B.n755 B.n8 585
R607 B.n753 B.n9 585
R608 B.n12 B.n9 585
R609 B.n752 B.n751 585
R610 B.n751 B.n750 585
R611 B.n11 B.n10 585
R612 B.n749 B.n11 585
R613 B.n747 B.n746 585
R614 B.n748 B.n747 585
R615 B.n745 B.n16 585
R616 B.n19 B.n16 585
R617 B.n744 B.n743 585
R618 B.n743 B.n742 585
R619 B.n18 B.n17 585
R620 B.n741 B.n18 585
R621 B.n739 B.n738 585
R622 B.n740 B.n739 585
R623 B.n737 B.n24 585
R624 B.n24 B.n23 585
R625 B.n736 B.n735 585
R626 B.n735 B.n734 585
R627 B.n26 B.n25 585
R628 B.n733 B.n26 585
R629 B.n731 B.n730 585
R630 B.n732 B.n731 585
R631 B.n729 B.n31 585
R632 B.n31 B.n30 585
R633 B.n728 B.n727 585
R634 B.n727 B.n726 585
R635 B.n33 B.n32 585
R636 B.n725 B.n33 585
R637 B.n723 B.n722 585
R638 B.n724 B.n723 585
R639 B.n721 B.n38 585
R640 B.n38 B.n37 585
R641 B.n720 B.n719 585
R642 B.n719 B.n718 585
R643 B.n40 B.n39 585
R644 B.n717 B.n40 585
R645 B.n715 B.n714 585
R646 B.n716 B.n715 585
R647 B.n713 B.n45 585
R648 B.n45 B.n44 585
R649 B.n712 B.n711 585
R650 B.n711 B.n710 585
R651 B.n47 B.n46 585
R652 B.n709 B.n47 585
R653 B.n707 B.n706 585
R654 B.n708 B.n707 585
R655 B.n705 B.n52 585
R656 B.n52 B.n51 585
R657 B.n704 B.n703 585
R658 B.n703 B.n702 585
R659 B.n54 B.n53 585
R660 B.n701 B.n54 585
R661 B.n699 B.n698 585
R662 B.n700 B.n699 585
R663 B.n697 B.n59 585
R664 B.n59 B.n58 585
R665 B.n696 B.n695 585
R666 B.n695 B.n694 585
R667 B.n61 B.n60 585
R668 B.n693 B.n61 585
R669 B.n691 B.n690 585
R670 B.n692 B.n691 585
R671 B.n689 B.n66 585
R672 B.n66 B.n65 585
R673 B.n688 B.n687 585
R674 B.n687 B.n686 585
R675 B.n68 B.n67 585
R676 B.n685 B.n68 585
R677 B.n683 B.n682 585
R678 B.n684 B.n683 585
R679 B.n681 B.n72 585
R680 B.n75 B.n72 585
R681 B.n680 B.n679 585
R682 B.n679 B.n678 585
R683 B.n74 B.n73 585
R684 B.n677 B.n74 585
R685 B.n675 B.n674 585
R686 B.n676 B.n675 585
R687 B.n673 B.n80 585
R688 B.n80 B.n79 585
R689 B.n672 B.n671 585
R690 B.n671 B.n670 585
R691 B.n82 B.n81 585
R692 B.n669 B.n82 585
R693 B.n667 B.n666 585
R694 B.n668 B.n667 585
R695 B.n665 B.n87 585
R696 B.n87 B.n86 585
R697 B.n664 B.n663 585
R698 B.n663 B.n662 585
R699 B.n89 B.n88 585
R700 B.n661 B.n89 585
R701 B.n659 B.n658 585
R702 B.n660 B.n659 585
R703 B.n657 B.n94 585
R704 B.n94 B.n93 585
R705 B.n656 B.n655 585
R706 B.n655 B.n654 585
R707 B.n96 B.n95 585
R708 B.n653 B.n96 585
R709 B.n651 B.n650 585
R710 B.n652 B.n651 585
R711 B.n649 B.n101 585
R712 B.n101 B.n100 585
R713 B.n648 B.n647 585
R714 B.n647 B.n646 585
R715 B.n103 B.n102 585
R716 B.n645 B.n103 585
R717 B.n643 B.n642 585
R718 B.n644 B.n643 585
R719 B.n641 B.n108 585
R720 B.n108 B.n107 585
R721 B.n640 B.n639 585
R722 B.n639 B.n638 585
R723 B.n110 B.n109 585
R724 B.n637 B.n110 585
R725 B.n760 B.n759 585
R726 B.n758 B.n2 585
R727 B.n132 B.n110 535.745
R728 B.n634 B.n112 535.745
R729 B.n368 B.n298 535.745
R730 B.n365 B.n296 535.745
R731 B.n129 B.t20 307.837
R732 B.n126 B.t10 307.837
R733 B.n316 B.t15 307.837
R734 B.n314 B.t18 307.837
R735 B.n636 B.n635 256.663
R736 B.n636 B.n124 256.663
R737 B.n636 B.n123 256.663
R738 B.n636 B.n122 256.663
R739 B.n636 B.n121 256.663
R740 B.n636 B.n120 256.663
R741 B.n636 B.n119 256.663
R742 B.n636 B.n118 256.663
R743 B.n636 B.n117 256.663
R744 B.n636 B.n116 256.663
R745 B.n636 B.n115 256.663
R746 B.n636 B.n114 256.663
R747 B.n636 B.n113 256.663
R748 B.n367 B.n366 256.663
R749 B.n367 B.n301 256.663
R750 B.n367 B.n302 256.663
R751 B.n367 B.n303 256.663
R752 B.n367 B.n304 256.663
R753 B.n367 B.n305 256.663
R754 B.n367 B.n306 256.663
R755 B.n367 B.n307 256.663
R756 B.n367 B.n308 256.663
R757 B.n367 B.n309 256.663
R758 B.n367 B.n310 256.663
R759 B.n367 B.n311 256.663
R760 B.n762 B.n761 256.663
R761 B.n367 B.n297 246.089
R762 B.n637 B.n636 246.089
R763 B.n130 B.t21 237.244
R764 B.n127 B.t11 237.244
R765 B.n317 B.t14 237.244
R766 B.n315 B.t17 237.244
R767 B.n129 B.t19 209.901
R768 B.n126 B.t8 209.901
R769 B.n316 B.t12 209.901
R770 B.n314 B.t16 209.901
R771 B.n136 B.n135 163.367
R772 B.n140 B.n139 163.367
R773 B.n144 B.n143 163.367
R774 B.n148 B.n147 163.367
R775 B.n152 B.n151 163.367
R776 B.n156 B.n155 163.367
R777 B.n160 B.n159 163.367
R778 B.n164 B.n163 163.367
R779 B.n168 B.n167 163.367
R780 B.n172 B.n171 163.367
R781 B.n176 B.n175 163.367
R782 B.n178 B.n125 163.367
R783 B.n372 B.n298 163.367
R784 B.n372 B.n292 163.367
R785 B.n380 B.n292 163.367
R786 B.n380 B.n290 163.367
R787 B.n384 B.n290 163.367
R788 B.n384 B.n283 163.367
R789 B.n392 B.n283 163.367
R790 B.n392 B.n281 163.367
R791 B.n396 B.n281 163.367
R792 B.n396 B.n276 163.367
R793 B.n404 B.n276 163.367
R794 B.n404 B.n274 163.367
R795 B.n408 B.n274 163.367
R796 B.n408 B.n268 163.367
R797 B.n416 B.n268 163.367
R798 B.n416 B.n266 163.367
R799 B.n420 B.n266 163.367
R800 B.n420 B.n260 163.367
R801 B.n428 B.n260 163.367
R802 B.n428 B.n258 163.367
R803 B.n432 B.n258 163.367
R804 B.n432 B.n253 163.367
R805 B.n441 B.n253 163.367
R806 B.n441 B.n251 163.367
R807 B.n445 B.n251 163.367
R808 B.n445 B.n245 163.367
R809 B.n453 B.n245 163.367
R810 B.n453 B.n243 163.367
R811 B.n457 B.n243 163.367
R812 B.n457 B.n237 163.367
R813 B.n465 B.n237 163.367
R814 B.n465 B.n235 163.367
R815 B.n469 B.n235 163.367
R816 B.n469 B.n229 163.367
R817 B.n477 B.n229 163.367
R818 B.n477 B.n227 163.367
R819 B.n481 B.n227 163.367
R820 B.n481 B.n221 163.367
R821 B.n489 B.n221 163.367
R822 B.n489 B.n219 163.367
R823 B.n493 B.n219 163.367
R824 B.n493 B.n213 163.367
R825 B.n501 B.n213 163.367
R826 B.n501 B.n211 163.367
R827 B.n505 B.n211 163.367
R828 B.n505 B.n205 163.367
R829 B.n513 B.n205 163.367
R830 B.n513 B.n203 163.367
R831 B.n517 B.n203 163.367
R832 B.n517 B.n197 163.367
R833 B.n525 B.n197 163.367
R834 B.n525 B.n195 163.367
R835 B.n529 B.n195 163.367
R836 B.n529 B.n190 163.367
R837 B.n538 B.n190 163.367
R838 B.n538 B.n188 163.367
R839 B.n543 B.n188 163.367
R840 B.n543 B.n182 163.367
R841 B.n551 B.n182 163.367
R842 B.n552 B.n551 163.367
R843 B.n552 B.n5 163.367
R844 B.n6 B.n5 163.367
R845 B.n7 B.n6 163.367
R846 B.n558 B.n7 163.367
R847 B.n559 B.n558 163.367
R848 B.n559 B.n13 163.367
R849 B.n14 B.n13 163.367
R850 B.n15 B.n14 163.367
R851 B.n564 B.n15 163.367
R852 B.n564 B.n20 163.367
R853 B.n21 B.n20 163.367
R854 B.n22 B.n21 163.367
R855 B.n569 B.n22 163.367
R856 B.n569 B.n27 163.367
R857 B.n28 B.n27 163.367
R858 B.n29 B.n28 163.367
R859 B.n574 B.n29 163.367
R860 B.n574 B.n34 163.367
R861 B.n35 B.n34 163.367
R862 B.n36 B.n35 163.367
R863 B.n579 B.n36 163.367
R864 B.n579 B.n41 163.367
R865 B.n42 B.n41 163.367
R866 B.n43 B.n42 163.367
R867 B.n584 B.n43 163.367
R868 B.n584 B.n48 163.367
R869 B.n49 B.n48 163.367
R870 B.n50 B.n49 163.367
R871 B.n589 B.n50 163.367
R872 B.n589 B.n55 163.367
R873 B.n56 B.n55 163.367
R874 B.n57 B.n56 163.367
R875 B.n594 B.n57 163.367
R876 B.n594 B.n62 163.367
R877 B.n63 B.n62 163.367
R878 B.n64 B.n63 163.367
R879 B.n599 B.n64 163.367
R880 B.n599 B.n69 163.367
R881 B.n70 B.n69 163.367
R882 B.n71 B.n70 163.367
R883 B.n604 B.n71 163.367
R884 B.n604 B.n76 163.367
R885 B.n77 B.n76 163.367
R886 B.n78 B.n77 163.367
R887 B.n609 B.n78 163.367
R888 B.n609 B.n83 163.367
R889 B.n84 B.n83 163.367
R890 B.n85 B.n84 163.367
R891 B.n614 B.n85 163.367
R892 B.n614 B.n90 163.367
R893 B.n91 B.n90 163.367
R894 B.n92 B.n91 163.367
R895 B.n619 B.n92 163.367
R896 B.n619 B.n97 163.367
R897 B.n98 B.n97 163.367
R898 B.n99 B.n98 163.367
R899 B.n624 B.n99 163.367
R900 B.n624 B.n104 163.367
R901 B.n105 B.n104 163.367
R902 B.n106 B.n105 163.367
R903 B.n629 B.n106 163.367
R904 B.n629 B.n111 163.367
R905 B.n112 B.n111 163.367
R906 B.n313 B.n312 163.367
R907 B.n360 B.n312 163.367
R908 B.n358 B.n357 163.367
R909 B.n354 B.n353 163.367
R910 B.n349 B.n348 163.367
R911 B.n345 B.n344 163.367
R912 B.n341 B.n340 163.367
R913 B.n337 B.n336 163.367
R914 B.n333 B.n332 163.367
R915 B.n328 B.n327 163.367
R916 B.n324 B.n323 163.367
R917 B.n320 B.n319 163.367
R918 B.n368 B.n300 163.367
R919 B.n374 B.n296 163.367
R920 B.n374 B.n294 163.367
R921 B.n378 B.n294 163.367
R922 B.n378 B.n288 163.367
R923 B.n386 B.n288 163.367
R924 B.n386 B.n286 163.367
R925 B.n390 B.n286 163.367
R926 B.n390 B.n280 163.367
R927 B.n398 B.n280 163.367
R928 B.n398 B.n278 163.367
R929 B.n402 B.n278 163.367
R930 B.n402 B.n272 163.367
R931 B.n410 B.n272 163.367
R932 B.n410 B.n270 163.367
R933 B.n414 B.n270 163.367
R934 B.n414 B.n264 163.367
R935 B.n422 B.n264 163.367
R936 B.n422 B.n262 163.367
R937 B.n426 B.n262 163.367
R938 B.n426 B.n256 163.367
R939 B.n435 B.n256 163.367
R940 B.n435 B.n254 163.367
R941 B.n439 B.n254 163.367
R942 B.n439 B.n249 163.367
R943 B.n447 B.n249 163.367
R944 B.n447 B.n247 163.367
R945 B.n451 B.n247 163.367
R946 B.n451 B.n241 163.367
R947 B.n459 B.n241 163.367
R948 B.n459 B.n239 163.367
R949 B.n463 B.n239 163.367
R950 B.n463 B.n233 163.367
R951 B.n471 B.n233 163.367
R952 B.n471 B.n231 163.367
R953 B.n475 B.n231 163.367
R954 B.n475 B.n225 163.367
R955 B.n483 B.n225 163.367
R956 B.n483 B.n223 163.367
R957 B.n487 B.n223 163.367
R958 B.n487 B.n217 163.367
R959 B.n495 B.n217 163.367
R960 B.n495 B.n215 163.367
R961 B.n499 B.n215 163.367
R962 B.n499 B.n209 163.367
R963 B.n507 B.n209 163.367
R964 B.n507 B.n207 163.367
R965 B.n511 B.n207 163.367
R966 B.n511 B.n201 163.367
R967 B.n519 B.n201 163.367
R968 B.n519 B.n199 163.367
R969 B.n523 B.n199 163.367
R970 B.n523 B.n193 163.367
R971 B.n532 B.n193 163.367
R972 B.n532 B.n191 163.367
R973 B.n536 B.n191 163.367
R974 B.n536 B.n186 163.367
R975 B.n545 B.n186 163.367
R976 B.n545 B.n184 163.367
R977 B.n549 B.n184 163.367
R978 B.n549 B.n3 163.367
R979 B.n760 B.n3 163.367
R980 B.n756 B.n2 163.367
R981 B.n756 B.n755 163.367
R982 B.n755 B.n9 163.367
R983 B.n751 B.n9 163.367
R984 B.n751 B.n11 163.367
R985 B.n747 B.n11 163.367
R986 B.n747 B.n16 163.367
R987 B.n743 B.n16 163.367
R988 B.n743 B.n18 163.367
R989 B.n739 B.n18 163.367
R990 B.n739 B.n24 163.367
R991 B.n735 B.n24 163.367
R992 B.n735 B.n26 163.367
R993 B.n731 B.n26 163.367
R994 B.n731 B.n31 163.367
R995 B.n727 B.n31 163.367
R996 B.n727 B.n33 163.367
R997 B.n723 B.n33 163.367
R998 B.n723 B.n38 163.367
R999 B.n719 B.n38 163.367
R1000 B.n719 B.n40 163.367
R1001 B.n715 B.n40 163.367
R1002 B.n715 B.n45 163.367
R1003 B.n711 B.n45 163.367
R1004 B.n711 B.n47 163.367
R1005 B.n707 B.n47 163.367
R1006 B.n707 B.n52 163.367
R1007 B.n703 B.n52 163.367
R1008 B.n703 B.n54 163.367
R1009 B.n699 B.n54 163.367
R1010 B.n699 B.n59 163.367
R1011 B.n695 B.n59 163.367
R1012 B.n695 B.n61 163.367
R1013 B.n691 B.n61 163.367
R1014 B.n691 B.n66 163.367
R1015 B.n687 B.n66 163.367
R1016 B.n687 B.n68 163.367
R1017 B.n683 B.n68 163.367
R1018 B.n683 B.n72 163.367
R1019 B.n679 B.n72 163.367
R1020 B.n679 B.n74 163.367
R1021 B.n675 B.n74 163.367
R1022 B.n675 B.n80 163.367
R1023 B.n671 B.n80 163.367
R1024 B.n671 B.n82 163.367
R1025 B.n667 B.n82 163.367
R1026 B.n667 B.n87 163.367
R1027 B.n663 B.n87 163.367
R1028 B.n663 B.n89 163.367
R1029 B.n659 B.n89 163.367
R1030 B.n659 B.n94 163.367
R1031 B.n655 B.n94 163.367
R1032 B.n655 B.n96 163.367
R1033 B.n651 B.n96 163.367
R1034 B.n651 B.n101 163.367
R1035 B.n647 B.n101 163.367
R1036 B.n647 B.n103 163.367
R1037 B.n643 B.n103 163.367
R1038 B.n643 B.n108 163.367
R1039 B.n639 B.n108 163.367
R1040 B.n639 B.n110 163.367
R1041 B.n373 B.n297 125.82
R1042 B.n373 B.n293 125.82
R1043 B.n379 B.n293 125.82
R1044 B.n379 B.n289 125.82
R1045 B.n385 B.n289 125.82
R1046 B.n385 B.n284 125.82
R1047 B.n391 B.n284 125.82
R1048 B.n391 B.n285 125.82
R1049 B.n397 B.n277 125.82
R1050 B.n403 B.n277 125.82
R1051 B.n403 B.n273 125.82
R1052 B.n409 B.n273 125.82
R1053 B.n409 B.n269 125.82
R1054 B.n415 B.n269 125.82
R1055 B.n415 B.n265 125.82
R1056 B.n421 B.n265 125.82
R1057 B.n421 B.n261 125.82
R1058 B.n427 B.n261 125.82
R1059 B.n427 B.n257 125.82
R1060 B.n434 B.n257 125.82
R1061 B.n434 B.n433 125.82
R1062 B.n440 B.n250 125.82
R1063 B.n446 B.n250 125.82
R1064 B.n446 B.n246 125.82
R1065 B.n452 B.n246 125.82
R1066 B.n452 B.n242 125.82
R1067 B.n458 B.n242 125.82
R1068 B.n458 B.n238 125.82
R1069 B.n464 B.n238 125.82
R1070 B.n464 B.n234 125.82
R1071 B.n470 B.n234 125.82
R1072 B.n476 B.n230 125.82
R1073 B.n476 B.n226 125.82
R1074 B.n482 B.n226 125.82
R1075 B.n482 B.n222 125.82
R1076 B.n488 B.n222 125.82
R1077 B.n488 B.n218 125.82
R1078 B.n494 B.n218 125.82
R1079 B.n494 B.n214 125.82
R1080 B.n500 B.n214 125.82
R1081 B.n506 B.n210 125.82
R1082 B.n506 B.n206 125.82
R1083 B.n512 B.n206 125.82
R1084 B.n512 B.n202 125.82
R1085 B.n518 B.n202 125.82
R1086 B.n518 B.n198 125.82
R1087 B.n524 B.n198 125.82
R1088 B.n524 B.n194 125.82
R1089 B.n531 B.n194 125.82
R1090 B.n531 B.n530 125.82
R1091 B.n537 B.n187 125.82
R1092 B.n544 B.n187 125.82
R1093 B.n544 B.n183 125.82
R1094 B.n550 B.n183 125.82
R1095 B.n550 B.n4 125.82
R1096 B.n759 B.n4 125.82
R1097 B.n759 B.n758 125.82
R1098 B.n758 B.n757 125.82
R1099 B.n757 B.n8 125.82
R1100 B.n12 B.n8 125.82
R1101 B.n750 B.n12 125.82
R1102 B.n750 B.n749 125.82
R1103 B.n749 B.n748 125.82
R1104 B.n742 B.n19 125.82
R1105 B.n742 B.n741 125.82
R1106 B.n741 B.n740 125.82
R1107 B.n740 B.n23 125.82
R1108 B.n734 B.n23 125.82
R1109 B.n734 B.n733 125.82
R1110 B.n733 B.n732 125.82
R1111 B.n732 B.n30 125.82
R1112 B.n726 B.n30 125.82
R1113 B.n726 B.n725 125.82
R1114 B.n724 B.n37 125.82
R1115 B.n718 B.n37 125.82
R1116 B.n718 B.n717 125.82
R1117 B.n717 B.n716 125.82
R1118 B.n716 B.n44 125.82
R1119 B.n710 B.n44 125.82
R1120 B.n710 B.n709 125.82
R1121 B.n709 B.n708 125.82
R1122 B.n708 B.n51 125.82
R1123 B.n702 B.n701 125.82
R1124 B.n701 B.n700 125.82
R1125 B.n700 B.n58 125.82
R1126 B.n694 B.n58 125.82
R1127 B.n694 B.n693 125.82
R1128 B.n693 B.n692 125.82
R1129 B.n692 B.n65 125.82
R1130 B.n686 B.n65 125.82
R1131 B.n686 B.n685 125.82
R1132 B.n685 B.n684 125.82
R1133 B.n678 B.n75 125.82
R1134 B.n678 B.n677 125.82
R1135 B.n677 B.n676 125.82
R1136 B.n676 B.n79 125.82
R1137 B.n670 B.n79 125.82
R1138 B.n670 B.n669 125.82
R1139 B.n669 B.n668 125.82
R1140 B.n668 B.n86 125.82
R1141 B.n662 B.n86 125.82
R1142 B.n662 B.n661 125.82
R1143 B.n661 B.n660 125.82
R1144 B.n660 B.n93 125.82
R1145 B.n654 B.n93 125.82
R1146 B.n653 B.n652 125.82
R1147 B.n652 B.n100 125.82
R1148 B.n646 B.n100 125.82
R1149 B.n646 B.n645 125.82
R1150 B.n645 B.n644 125.82
R1151 B.n644 B.n107 125.82
R1152 B.n638 B.n107 125.82
R1153 B.n638 B.n637 125.82
R1154 B.t2 B.n230 109.168
R1155 B.t5 B.n51 109.168
R1156 B.n500 B.t7 105.468
R1157 B.t4 B.n724 105.468
R1158 B.n440 B.t3 72.162
R1159 B.n684 B.t1 72.162
R1160 B.n132 B.n113 71.676
R1161 B.n136 B.n114 71.676
R1162 B.n140 B.n115 71.676
R1163 B.n144 B.n116 71.676
R1164 B.n148 B.n117 71.676
R1165 B.n152 B.n118 71.676
R1166 B.n156 B.n119 71.676
R1167 B.n160 B.n120 71.676
R1168 B.n164 B.n121 71.676
R1169 B.n168 B.n122 71.676
R1170 B.n172 B.n123 71.676
R1171 B.n176 B.n124 71.676
R1172 B.n635 B.n125 71.676
R1173 B.n635 B.n634 71.676
R1174 B.n178 B.n124 71.676
R1175 B.n175 B.n123 71.676
R1176 B.n171 B.n122 71.676
R1177 B.n167 B.n121 71.676
R1178 B.n163 B.n120 71.676
R1179 B.n159 B.n119 71.676
R1180 B.n155 B.n118 71.676
R1181 B.n151 B.n117 71.676
R1182 B.n147 B.n116 71.676
R1183 B.n143 B.n115 71.676
R1184 B.n139 B.n114 71.676
R1185 B.n135 B.n113 71.676
R1186 B.n366 B.n365 71.676
R1187 B.n360 B.n301 71.676
R1188 B.n357 B.n302 71.676
R1189 B.n353 B.n303 71.676
R1190 B.n348 B.n304 71.676
R1191 B.n344 B.n305 71.676
R1192 B.n340 B.n306 71.676
R1193 B.n336 B.n307 71.676
R1194 B.n332 B.n308 71.676
R1195 B.n327 B.n309 71.676
R1196 B.n323 B.n310 71.676
R1197 B.n319 B.n311 71.676
R1198 B.n366 B.n313 71.676
R1199 B.n358 B.n301 71.676
R1200 B.n354 B.n302 71.676
R1201 B.n349 B.n303 71.676
R1202 B.n345 B.n304 71.676
R1203 B.n341 B.n305 71.676
R1204 B.n337 B.n306 71.676
R1205 B.n333 B.n307 71.676
R1206 B.n328 B.n308 71.676
R1207 B.n324 B.n309 71.676
R1208 B.n320 B.n310 71.676
R1209 B.n311 B.n300 71.676
R1210 B.n761 B.n760 71.676
R1211 B.n761 B.n2 71.676
R1212 B.n130 B.n129 70.5944
R1213 B.n127 B.n126 70.5944
R1214 B.n317 B.n316 70.5944
R1215 B.n315 B.n314 70.5944
R1216 B.n530 B.t0 68.4614
R1217 B.n19 B.t6 68.4614
R1218 B.n285 B.t13 64.7608
R1219 B.t9 B.n653 64.7608
R1220 B.n397 B.t13 61.0602
R1221 B.n654 B.t9 61.0602
R1222 B.n131 B.n130 59.5399
R1223 B.n128 B.n127 59.5399
R1224 B.n330 B.n317 59.5399
R1225 B.n351 B.n315 59.5399
R1226 B.n537 B.t0 57.3596
R1227 B.n748 B.t6 57.3596
R1228 B.n433 B.t3 53.659
R1229 B.n75 B.t1 53.659
R1230 B.n364 B.n295 34.8103
R1231 B.n370 B.n369 34.8103
R1232 B.n633 B.n632 34.8103
R1233 B.n133 B.n109 34.8103
R1234 B.t7 B.n210 20.3537
R1235 B.n725 B.t4 20.3537
R1236 B B.n762 18.0485
R1237 B.n470 B.t2 16.6531
R1238 B.n702 B.t5 16.6531
R1239 B.n375 B.n295 10.6151
R1240 B.n376 B.n375 10.6151
R1241 B.n377 B.n376 10.6151
R1242 B.n377 B.n287 10.6151
R1243 B.n387 B.n287 10.6151
R1244 B.n388 B.n387 10.6151
R1245 B.n389 B.n388 10.6151
R1246 B.n389 B.n279 10.6151
R1247 B.n399 B.n279 10.6151
R1248 B.n400 B.n399 10.6151
R1249 B.n401 B.n400 10.6151
R1250 B.n401 B.n271 10.6151
R1251 B.n411 B.n271 10.6151
R1252 B.n412 B.n411 10.6151
R1253 B.n413 B.n412 10.6151
R1254 B.n413 B.n263 10.6151
R1255 B.n423 B.n263 10.6151
R1256 B.n424 B.n423 10.6151
R1257 B.n425 B.n424 10.6151
R1258 B.n425 B.n255 10.6151
R1259 B.n436 B.n255 10.6151
R1260 B.n437 B.n436 10.6151
R1261 B.n438 B.n437 10.6151
R1262 B.n438 B.n248 10.6151
R1263 B.n448 B.n248 10.6151
R1264 B.n449 B.n448 10.6151
R1265 B.n450 B.n449 10.6151
R1266 B.n450 B.n240 10.6151
R1267 B.n460 B.n240 10.6151
R1268 B.n461 B.n460 10.6151
R1269 B.n462 B.n461 10.6151
R1270 B.n462 B.n232 10.6151
R1271 B.n472 B.n232 10.6151
R1272 B.n473 B.n472 10.6151
R1273 B.n474 B.n473 10.6151
R1274 B.n474 B.n224 10.6151
R1275 B.n484 B.n224 10.6151
R1276 B.n485 B.n484 10.6151
R1277 B.n486 B.n485 10.6151
R1278 B.n486 B.n216 10.6151
R1279 B.n496 B.n216 10.6151
R1280 B.n497 B.n496 10.6151
R1281 B.n498 B.n497 10.6151
R1282 B.n498 B.n208 10.6151
R1283 B.n508 B.n208 10.6151
R1284 B.n509 B.n508 10.6151
R1285 B.n510 B.n509 10.6151
R1286 B.n510 B.n200 10.6151
R1287 B.n520 B.n200 10.6151
R1288 B.n521 B.n520 10.6151
R1289 B.n522 B.n521 10.6151
R1290 B.n522 B.n192 10.6151
R1291 B.n533 B.n192 10.6151
R1292 B.n534 B.n533 10.6151
R1293 B.n535 B.n534 10.6151
R1294 B.n535 B.n185 10.6151
R1295 B.n546 B.n185 10.6151
R1296 B.n547 B.n546 10.6151
R1297 B.n548 B.n547 10.6151
R1298 B.n548 B.n0 10.6151
R1299 B.n364 B.n363 10.6151
R1300 B.n363 B.n362 10.6151
R1301 B.n362 B.n361 10.6151
R1302 B.n361 B.n359 10.6151
R1303 B.n359 B.n356 10.6151
R1304 B.n356 B.n355 10.6151
R1305 B.n355 B.n352 10.6151
R1306 B.n350 B.n347 10.6151
R1307 B.n347 B.n346 10.6151
R1308 B.n346 B.n343 10.6151
R1309 B.n343 B.n342 10.6151
R1310 B.n342 B.n339 10.6151
R1311 B.n339 B.n338 10.6151
R1312 B.n338 B.n335 10.6151
R1313 B.n335 B.n334 10.6151
R1314 B.n334 B.n331 10.6151
R1315 B.n329 B.n326 10.6151
R1316 B.n326 B.n325 10.6151
R1317 B.n325 B.n322 10.6151
R1318 B.n322 B.n321 10.6151
R1319 B.n321 B.n318 10.6151
R1320 B.n318 B.n299 10.6151
R1321 B.n369 B.n299 10.6151
R1322 B.n371 B.n370 10.6151
R1323 B.n371 B.n291 10.6151
R1324 B.n381 B.n291 10.6151
R1325 B.n382 B.n381 10.6151
R1326 B.n383 B.n382 10.6151
R1327 B.n383 B.n282 10.6151
R1328 B.n393 B.n282 10.6151
R1329 B.n394 B.n393 10.6151
R1330 B.n395 B.n394 10.6151
R1331 B.n395 B.n275 10.6151
R1332 B.n405 B.n275 10.6151
R1333 B.n406 B.n405 10.6151
R1334 B.n407 B.n406 10.6151
R1335 B.n407 B.n267 10.6151
R1336 B.n417 B.n267 10.6151
R1337 B.n418 B.n417 10.6151
R1338 B.n419 B.n418 10.6151
R1339 B.n419 B.n259 10.6151
R1340 B.n429 B.n259 10.6151
R1341 B.n430 B.n429 10.6151
R1342 B.n431 B.n430 10.6151
R1343 B.n431 B.n252 10.6151
R1344 B.n442 B.n252 10.6151
R1345 B.n443 B.n442 10.6151
R1346 B.n444 B.n443 10.6151
R1347 B.n444 B.n244 10.6151
R1348 B.n454 B.n244 10.6151
R1349 B.n455 B.n454 10.6151
R1350 B.n456 B.n455 10.6151
R1351 B.n456 B.n236 10.6151
R1352 B.n466 B.n236 10.6151
R1353 B.n467 B.n466 10.6151
R1354 B.n468 B.n467 10.6151
R1355 B.n468 B.n228 10.6151
R1356 B.n478 B.n228 10.6151
R1357 B.n479 B.n478 10.6151
R1358 B.n480 B.n479 10.6151
R1359 B.n480 B.n220 10.6151
R1360 B.n490 B.n220 10.6151
R1361 B.n491 B.n490 10.6151
R1362 B.n492 B.n491 10.6151
R1363 B.n492 B.n212 10.6151
R1364 B.n502 B.n212 10.6151
R1365 B.n503 B.n502 10.6151
R1366 B.n504 B.n503 10.6151
R1367 B.n504 B.n204 10.6151
R1368 B.n514 B.n204 10.6151
R1369 B.n515 B.n514 10.6151
R1370 B.n516 B.n515 10.6151
R1371 B.n516 B.n196 10.6151
R1372 B.n526 B.n196 10.6151
R1373 B.n527 B.n526 10.6151
R1374 B.n528 B.n527 10.6151
R1375 B.n528 B.n189 10.6151
R1376 B.n539 B.n189 10.6151
R1377 B.n540 B.n539 10.6151
R1378 B.n542 B.n540 10.6151
R1379 B.n542 B.n541 10.6151
R1380 B.n541 B.n181 10.6151
R1381 B.n553 B.n181 10.6151
R1382 B.n554 B.n553 10.6151
R1383 B.n555 B.n554 10.6151
R1384 B.n556 B.n555 10.6151
R1385 B.n557 B.n556 10.6151
R1386 B.n560 B.n557 10.6151
R1387 B.n561 B.n560 10.6151
R1388 B.n562 B.n561 10.6151
R1389 B.n563 B.n562 10.6151
R1390 B.n565 B.n563 10.6151
R1391 B.n566 B.n565 10.6151
R1392 B.n567 B.n566 10.6151
R1393 B.n568 B.n567 10.6151
R1394 B.n570 B.n568 10.6151
R1395 B.n571 B.n570 10.6151
R1396 B.n572 B.n571 10.6151
R1397 B.n573 B.n572 10.6151
R1398 B.n575 B.n573 10.6151
R1399 B.n576 B.n575 10.6151
R1400 B.n577 B.n576 10.6151
R1401 B.n578 B.n577 10.6151
R1402 B.n580 B.n578 10.6151
R1403 B.n581 B.n580 10.6151
R1404 B.n582 B.n581 10.6151
R1405 B.n583 B.n582 10.6151
R1406 B.n585 B.n583 10.6151
R1407 B.n586 B.n585 10.6151
R1408 B.n587 B.n586 10.6151
R1409 B.n588 B.n587 10.6151
R1410 B.n590 B.n588 10.6151
R1411 B.n591 B.n590 10.6151
R1412 B.n592 B.n591 10.6151
R1413 B.n593 B.n592 10.6151
R1414 B.n595 B.n593 10.6151
R1415 B.n596 B.n595 10.6151
R1416 B.n597 B.n596 10.6151
R1417 B.n598 B.n597 10.6151
R1418 B.n600 B.n598 10.6151
R1419 B.n601 B.n600 10.6151
R1420 B.n602 B.n601 10.6151
R1421 B.n603 B.n602 10.6151
R1422 B.n605 B.n603 10.6151
R1423 B.n606 B.n605 10.6151
R1424 B.n607 B.n606 10.6151
R1425 B.n608 B.n607 10.6151
R1426 B.n610 B.n608 10.6151
R1427 B.n611 B.n610 10.6151
R1428 B.n612 B.n611 10.6151
R1429 B.n613 B.n612 10.6151
R1430 B.n615 B.n613 10.6151
R1431 B.n616 B.n615 10.6151
R1432 B.n617 B.n616 10.6151
R1433 B.n618 B.n617 10.6151
R1434 B.n620 B.n618 10.6151
R1435 B.n621 B.n620 10.6151
R1436 B.n622 B.n621 10.6151
R1437 B.n623 B.n622 10.6151
R1438 B.n625 B.n623 10.6151
R1439 B.n626 B.n625 10.6151
R1440 B.n627 B.n626 10.6151
R1441 B.n628 B.n627 10.6151
R1442 B.n630 B.n628 10.6151
R1443 B.n631 B.n630 10.6151
R1444 B.n632 B.n631 10.6151
R1445 B.n754 B.n1 10.6151
R1446 B.n754 B.n753 10.6151
R1447 B.n753 B.n752 10.6151
R1448 B.n752 B.n10 10.6151
R1449 B.n746 B.n10 10.6151
R1450 B.n746 B.n745 10.6151
R1451 B.n745 B.n744 10.6151
R1452 B.n744 B.n17 10.6151
R1453 B.n738 B.n17 10.6151
R1454 B.n738 B.n737 10.6151
R1455 B.n737 B.n736 10.6151
R1456 B.n736 B.n25 10.6151
R1457 B.n730 B.n25 10.6151
R1458 B.n730 B.n729 10.6151
R1459 B.n729 B.n728 10.6151
R1460 B.n728 B.n32 10.6151
R1461 B.n722 B.n32 10.6151
R1462 B.n722 B.n721 10.6151
R1463 B.n721 B.n720 10.6151
R1464 B.n720 B.n39 10.6151
R1465 B.n714 B.n39 10.6151
R1466 B.n714 B.n713 10.6151
R1467 B.n713 B.n712 10.6151
R1468 B.n712 B.n46 10.6151
R1469 B.n706 B.n46 10.6151
R1470 B.n706 B.n705 10.6151
R1471 B.n705 B.n704 10.6151
R1472 B.n704 B.n53 10.6151
R1473 B.n698 B.n53 10.6151
R1474 B.n698 B.n697 10.6151
R1475 B.n697 B.n696 10.6151
R1476 B.n696 B.n60 10.6151
R1477 B.n690 B.n60 10.6151
R1478 B.n690 B.n689 10.6151
R1479 B.n689 B.n688 10.6151
R1480 B.n688 B.n67 10.6151
R1481 B.n682 B.n67 10.6151
R1482 B.n682 B.n681 10.6151
R1483 B.n681 B.n680 10.6151
R1484 B.n680 B.n73 10.6151
R1485 B.n674 B.n73 10.6151
R1486 B.n674 B.n673 10.6151
R1487 B.n673 B.n672 10.6151
R1488 B.n672 B.n81 10.6151
R1489 B.n666 B.n81 10.6151
R1490 B.n666 B.n665 10.6151
R1491 B.n665 B.n664 10.6151
R1492 B.n664 B.n88 10.6151
R1493 B.n658 B.n88 10.6151
R1494 B.n658 B.n657 10.6151
R1495 B.n657 B.n656 10.6151
R1496 B.n656 B.n95 10.6151
R1497 B.n650 B.n95 10.6151
R1498 B.n650 B.n649 10.6151
R1499 B.n649 B.n648 10.6151
R1500 B.n648 B.n102 10.6151
R1501 B.n642 B.n102 10.6151
R1502 B.n642 B.n641 10.6151
R1503 B.n641 B.n640 10.6151
R1504 B.n640 B.n109 10.6151
R1505 B.n134 B.n133 10.6151
R1506 B.n137 B.n134 10.6151
R1507 B.n138 B.n137 10.6151
R1508 B.n141 B.n138 10.6151
R1509 B.n142 B.n141 10.6151
R1510 B.n145 B.n142 10.6151
R1511 B.n146 B.n145 10.6151
R1512 B.n150 B.n149 10.6151
R1513 B.n153 B.n150 10.6151
R1514 B.n154 B.n153 10.6151
R1515 B.n157 B.n154 10.6151
R1516 B.n158 B.n157 10.6151
R1517 B.n161 B.n158 10.6151
R1518 B.n162 B.n161 10.6151
R1519 B.n165 B.n162 10.6151
R1520 B.n166 B.n165 10.6151
R1521 B.n170 B.n169 10.6151
R1522 B.n173 B.n170 10.6151
R1523 B.n174 B.n173 10.6151
R1524 B.n177 B.n174 10.6151
R1525 B.n179 B.n177 10.6151
R1526 B.n180 B.n179 10.6151
R1527 B.n633 B.n180 10.6151
R1528 B.n352 B.n351 9.36635
R1529 B.n330 B.n329 9.36635
R1530 B.n146 B.n131 9.36635
R1531 B.n169 B.n128 9.36635
R1532 B.n762 B.n0 8.11757
R1533 B.n762 B.n1 8.11757
R1534 B.n351 B.n350 1.24928
R1535 B.n331 B.n330 1.24928
R1536 B.n149 B.n131 1.24928
R1537 B.n166 B.n128 1.24928
R1538 VN.n68 VN.n67 161.3
R1539 VN.n66 VN.n36 161.3
R1540 VN.n65 VN.n64 161.3
R1541 VN.n63 VN.n37 161.3
R1542 VN.n62 VN.n61 161.3
R1543 VN.n60 VN.n38 161.3
R1544 VN.n59 VN.n58 161.3
R1545 VN.n57 VN.n56 161.3
R1546 VN.n55 VN.n40 161.3
R1547 VN.n54 VN.n53 161.3
R1548 VN.n52 VN.n41 161.3
R1549 VN.n51 VN.n50 161.3
R1550 VN.n49 VN.n42 161.3
R1551 VN.n48 VN.n47 161.3
R1552 VN.n46 VN.n43 161.3
R1553 VN.n33 VN.n32 161.3
R1554 VN.n31 VN.n1 161.3
R1555 VN.n30 VN.n29 161.3
R1556 VN.n28 VN.n2 161.3
R1557 VN.n27 VN.n26 161.3
R1558 VN.n25 VN.n3 161.3
R1559 VN.n24 VN.n23 161.3
R1560 VN.n22 VN.n21 161.3
R1561 VN.n20 VN.n5 161.3
R1562 VN.n19 VN.n18 161.3
R1563 VN.n17 VN.n6 161.3
R1564 VN.n16 VN.n15 161.3
R1565 VN.n14 VN.n7 161.3
R1566 VN.n13 VN.n12 161.3
R1567 VN.n11 VN.n8 161.3
R1568 VN.n34 VN.n0 79.7913
R1569 VN.n69 VN.n35 79.7913
R1570 VN.n10 VN.n9 71.1565
R1571 VN.n45 VN.n44 71.1565
R1572 VN.n15 VN.n6 56.5193
R1573 VN.n50 VN.n41 56.5193
R1574 VN.n26 VN.n2 51.1773
R1575 VN.n61 VN.n37 51.1773
R1576 VN VN.n69 45.8465
R1577 VN.n45 VN.t7 37.0503
R1578 VN.n10 VN.t6 37.0503
R1579 VN.n30 VN.n2 29.8095
R1580 VN.n65 VN.n37 29.8095
R1581 VN.n13 VN.n8 24.4675
R1582 VN.n14 VN.n13 24.4675
R1583 VN.n15 VN.n14 24.4675
R1584 VN.n19 VN.n6 24.4675
R1585 VN.n20 VN.n19 24.4675
R1586 VN.n21 VN.n20 24.4675
R1587 VN.n25 VN.n24 24.4675
R1588 VN.n26 VN.n25 24.4675
R1589 VN.n31 VN.n30 24.4675
R1590 VN.n32 VN.n31 24.4675
R1591 VN.n50 VN.n49 24.4675
R1592 VN.n49 VN.n48 24.4675
R1593 VN.n48 VN.n43 24.4675
R1594 VN.n61 VN.n60 24.4675
R1595 VN.n60 VN.n59 24.4675
R1596 VN.n56 VN.n55 24.4675
R1597 VN.n55 VN.n54 24.4675
R1598 VN.n54 VN.n41 24.4675
R1599 VN.n67 VN.n66 24.4675
R1600 VN.n66 VN.n65 24.4675
R1601 VN.n24 VN.n4 21.0421
R1602 VN.n59 VN.n39 21.0421
R1603 VN.n32 VN.n0 10.2766
R1604 VN.n67 VN.n35 10.2766
R1605 VN.n9 VN.t5 4.87875
R1606 VN.n4 VN.t4 4.87875
R1607 VN.n0 VN.t2 4.87875
R1608 VN.n44 VN.t3 4.87875
R1609 VN.n39 VN.t1 4.87875
R1610 VN.n35 VN.t0 4.87875
R1611 VN.n46 VN.n45 4.39147
R1612 VN.n11 VN.n10 4.39147
R1613 VN.n9 VN.n8 3.42588
R1614 VN.n21 VN.n4 3.42588
R1615 VN.n44 VN.n43 3.42588
R1616 VN.n56 VN.n39 3.42588
R1617 VN.n69 VN.n68 0.354971
R1618 VN.n34 VN.n33 0.354971
R1619 VN VN.n34 0.26696
R1620 VN.n68 VN.n36 0.189894
R1621 VN.n64 VN.n36 0.189894
R1622 VN.n64 VN.n63 0.189894
R1623 VN.n63 VN.n62 0.189894
R1624 VN.n62 VN.n38 0.189894
R1625 VN.n58 VN.n38 0.189894
R1626 VN.n58 VN.n57 0.189894
R1627 VN.n57 VN.n40 0.189894
R1628 VN.n53 VN.n40 0.189894
R1629 VN.n53 VN.n52 0.189894
R1630 VN.n52 VN.n51 0.189894
R1631 VN.n51 VN.n42 0.189894
R1632 VN.n47 VN.n42 0.189894
R1633 VN.n47 VN.n46 0.189894
R1634 VN.n12 VN.n11 0.189894
R1635 VN.n12 VN.n7 0.189894
R1636 VN.n16 VN.n7 0.189894
R1637 VN.n17 VN.n16 0.189894
R1638 VN.n18 VN.n17 0.189894
R1639 VN.n18 VN.n5 0.189894
R1640 VN.n22 VN.n5 0.189894
R1641 VN.n23 VN.n22 0.189894
R1642 VN.n23 VN.n3 0.189894
R1643 VN.n27 VN.n3 0.189894
R1644 VN.n28 VN.n27 0.189894
R1645 VN.n29 VN.n28 0.189894
R1646 VN.n29 VN.n1 0.189894
R1647 VN.n33 VN.n1 0.189894
R1648 VDD2.n2 VDD2.n1 236.736
R1649 VDD2.n2 VDD2.n0 236.736
R1650 VDD2 VDD2.n5 236.732
R1651 VDD2.n4 VDD2.n3 235.221
R1652 VDD2.n4 VDD2.n2 38.4136
R1653 VDD2.n5 VDD2.t4 29.5527
R1654 VDD2.n5 VDD2.t0 29.5527
R1655 VDD2.n3 VDD2.t7 29.5527
R1656 VDD2.n3 VDD2.t6 29.5527
R1657 VDD2.n1 VDD2.t3 29.5527
R1658 VDD2.n1 VDD2.t5 29.5527
R1659 VDD2.n0 VDD2.t1 29.5527
R1660 VDD2.n0 VDD2.t2 29.5527
R1661 VDD2 VDD2.n4 1.62766
C0 VN VDD2 0.964559f
C1 VN VDD1 0.160619f
C2 VTAIL VDD2 5.02514f
C3 VTAIL VDD1 4.96596f
C4 VN VP 6.44652f
C5 VDD1 VDD2 2.14413f
C6 VP VTAIL 2.69f
C7 VP VDD2 0.605445f
C8 VP VDD1 1.40427f
C9 VN VTAIL 2.67589f
C10 VDD2 B 5.176694f
C11 VDD1 B 5.670357f
C12 VTAIL B 3.597411f
C13 VN B 17.5053f
C14 VP B 15.814066f
C15 VDD2.t1 B 0.016061f
C16 VDD2.t2 B 0.016061f
C17 VDD2.n0 B 0.043528f
C18 VDD2.t3 B 0.016061f
C19 VDD2.t5 B 0.016061f
C20 VDD2.n1 B 0.043528f
C21 VDD2.n2 B 3.31525f
C22 VDD2.t7 B 0.016061f
C23 VDD2.t6 B 0.016061f
C24 VDD2.n3 B 0.040047f
C25 VDD2.n4 B 2.63874f
C26 VDD2.t4 B 0.016061f
C27 VDD2.t0 B 0.016061f
C28 VDD2.n5 B 0.043517f
C29 VN.t2 B 0.097175f
C30 VN.n0 B 0.20761f
C31 VN.n1 B 0.031116f
C32 VN.n2 B 0.030352f
C33 VN.n3 B 0.031116f
C34 VN.t4 B 0.097175f
C35 VN.n4 B 0.093094f
C36 VN.n5 B 0.031116f
C37 VN.n6 B 0.045424f
C38 VN.n7 B 0.031116f
C39 VN.n8 B 0.03337f
C40 VN.t5 B 0.097175f
C41 VN.n9 B 0.188353f
C42 VN.t6 B 0.36727f
C43 VN.n10 B 0.241588f
C44 VN.n11 B 0.368156f
C45 VN.n12 B 0.031116f
C46 VN.n13 B 0.057992f
C47 VN.n14 B 0.057992f
C48 VN.n15 B 0.045424f
C49 VN.n16 B 0.031116f
C50 VN.n17 B 0.031116f
C51 VN.n18 B 0.031116f
C52 VN.n19 B 0.057992f
C53 VN.n20 B 0.057992f
C54 VN.n21 B 0.03337f
C55 VN.n22 B 0.031116f
C56 VN.n23 B 0.031116f
C57 VN.n24 B 0.053984f
C58 VN.n25 B 0.057992f
C59 VN.n26 B 0.056496f
C60 VN.n27 B 0.031116f
C61 VN.n28 B 0.031116f
C62 VN.n29 B 0.031116f
C63 VN.n30 B 0.061993f
C64 VN.n31 B 0.057992f
C65 VN.n32 B 0.041386f
C66 VN.n33 B 0.050221f
C67 VN.n34 B 0.080481f
C68 VN.t0 B 0.097175f
C69 VN.n35 B 0.20761f
C70 VN.n36 B 0.031116f
C71 VN.n37 B 0.030352f
C72 VN.n38 B 0.031116f
C73 VN.t1 B 0.097175f
C74 VN.n39 B 0.093094f
C75 VN.n40 B 0.031116f
C76 VN.n41 B 0.045424f
C77 VN.n42 B 0.031116f
C78 VN.n43 B 0.03337f
C79 VN.t7 B 0.36727f
C80 VN.t3 B 0.097175f
C81 VN.n44 B 0.188353f
C82 VN.n45 B 0.241588f
C83 VN.n46 B 0.368156f
C84 VN.n47 B 0.031116f
C85 VN.n48 B 0.057992f
C86 VN.n49 B 0.057992f
C87 VN.n50 B 0.045424f
C88 VN.n51 B 0.031116f
C89 VN.n52 B 0.031116f
C90 VN.n53 B 0.031116f
C91 VN.n54 B 0.057992f
C92 VN.n55 B 0.057992f
C93 VN.n56 B 0.03337f
C94 VN.n57 B 0.031116f
C95 VN.n58 B 0.031116f
C96 VN.n59 B 0.053984f
C97 VN.n60 B 0.057992f
C98 VN.n61 B 0.056496f
C99 VN.n62 B 0.031116f
C100 VN.n63 B 0.031116f
C101 VN.n64 B 0.031116f
C102 VN.n65 B 0.061993f
C103 VN.n66 B 0.057992f
C104 VN.n67 B 0.041386f
C105 VN.n68 B 0.050221f
C106 VN.n69 B 1.56696f
C107 VTAIL.t4 B 0.025814f
C108 VTAIL.t5 B 0.025814f
C109 VTAIL.n0 B 0.055624f
C110 VTAIL.n1 B 0.568436f
C111 VTAIL.t6 B 0.11409f
C112 VTAIL.n2 B 0.645043f
C113 VTAIL.t13 B 0.11409f
C114 VTAIL.n3 B 0.645043f
C115 VTAIL.t9 B 0.025814f
C116 VTAIL.t14 B 0.025814f
C117 VTAIL.n4 B 0.055624f
C118 VTAIL.n5 B 1.05228f
C119 VTAIL.t8 B 0.11409f
C120 VTAIL.n6 B 1.81725f
C121 VTAIL.t3 B 0.11409f
C122 VTAIL.n7 B 1.81725f
C123 VTAIL.t2 B 0.025814f
C124 VTAIL.t7 B 0.025814f
C125 VTAIL.n8 B 0.055624f
C126 VTAIL.n9 B 1.05228f
C127 VTAIL.t0 B 0.11409f
C128 VTAIL.n10 B 0.645043f
C129 VTAIL.t11 B 0.11409f
C130 VTAIL.n11 B 0.645043f
C131 VTAIL.t12 B 0.025814f
C132 VTAIL.t15 B 0.025814f
C133 VTAIL.n12 B 0.055624f
C134 VTAIL.n13 B 1.05228f
C135 VTAIL.t10 B 0.11409f
C136 VTAIL.n14 B 1.81725f
C137 VTAIL.t1 B 0.11409f
C138 VTAIL.n15 B 1.80811f
C139 VDD1.t1 B 0.015811f
C140 VDD1.t0 B 0.015811f
C141 VDD1.n0 B 0.043179f
C142 VDD1.t6 B 0.015811f
C143 VDD1.t3 B 0.015811f
C144 VDD1.n1 B 0.042852f
C145 VDD1.t4 B 0.015811f
C146 VDD1.t2 B 0.015811f
C147 VDD1.n2 B 0.042852f
C148 VDD1.n3 B 3.32573f
C149 VDD1.t7 B 0.015811f
C150 VDD1.t5 B 0.015811f
C151 VDD1.n4 B 0.039425f
C152 VDD1.n5 B 2.63487f
C153 VP.t2 B 0.097644f
C154 VP.n0 B 0.208613f
C155 VP.n1 B 0.031266f
C156 VP.n2 B 0.030498f
C157 VP.n3 B 0.031266f
C158 VP.t1 B 0.097644f
C159 VP.n4 B 0.093543f
C160 VP.n5 B 0.031266f
C161 VP.n6 B 0.045643f
C162 VP.n7 B 0.031266f
C163 VP.n8 B 0.033531f
C164 VP.n9 B 0.031266f
C165 VP.n10 B 0.030498f
C166 VP.n11 B 0.031266f
C167 VP.t7 B 0.097644f
C168 VP.n12 B 0.208613f
C169 VP.t5 B 0.097644f
C170 VP.n13 B 0.208613f
C171 VP.n14 B 0.031266f
C172 VP.n15 B 0.030498f
C173 VP.n16 B 0.031266f
C174 VP.t0 B 0.097644f
C175 VP.n17 B 0.093543f
C176 VP.n18 B 0.031266f
C177 VP.n19 B 0.045643f
C178 VP.n20 B 0.031266f
C179 VP.n21 B 0.033531f
C180 VP.t4 B 0.369044f
C181 VP.t3 B 0.097644f
C182 VP.n22 B 0.189263f
C183 VP.n23 B 0.242756f
C184 VP.n24 B 0.369935f
C185 VP.n25 B 0.031266f
C186 VP.n26 B 0.058273f
C187 VP.n27 B 0.058273f
C188 VP.n28 B 0.045643f
C189 VP.n29 B 0.031266f
C190 VP.n30 B 0.031266f
C191 VP.n31 B 0.031266f
C192 VP.n32 B 0.058273f
C193 VP.n33 B 0.058273f
C194 VP.n34 B 0.033531f
C195 VP.n35 B 0.031266f
C196 VP.n36 B 0.031266f
C197 VP.n37 B 0.054245f
C198 VP.n38 B 0.058273f
C199 VP.n39 B 0.056768f
C200 VP.n40 B 0.031266f
C201 VP.n41 B 0.031266f
C202 VP.n42 B 0.031266f
C203 VP.n43 B 0.062292f
C204 VP.n44 B 0.058273f
C205 VP.n45 B 0.041586f
C206 VP.n46 B 0.050463f
C207 VP.n47 B 1.56131f
C208 VP.n48 B 1.58592f
C209 VP.n49 B 0.050463f
C210 VP.n50 B 0.041586f
C211 VP.n51 B 0.058273f
C212 VP.n52 B 0.062292f
C213 VP.n53 B 0.031266f
C214 VP.n54 B 0.031266f
C215 VP.n55 B 0.031266f
C216 VP.n56 B 0.056768f
C217 VP.n57 B 0.058273f
C218 VP.t6 B 0.097644f
C219 VP.n58 B 0.093543f
C220 VP.n59 B 0.054245f
C221 VP.n60 B 0.031266f
C222 VP.n61 B 0.031266f
C223 VP.n62 B 0.031266f
C224 VP.n63 B 0.058273f
C225 VP.n64 B 0.058273f
C226 VP.n65 B 0.045643f
C227 VP.n66 B 0.031266f
C228 VP.n67 B 0.031266f
C229 VP.n68 B 0.031266f
C230 VP.n69 B 0.058273f
C231 VP.n70 B 0.058273f
C232 VP.n71 B 0.033531f
C233 VP.n72 B 0.031266f
C234 VP.n73 B 0.031266f
C235 VP.n74 B 0.054245f
C236 VP.n75 B 0.058273f
C237 VP.n76 B 0.056768f
C238 VP.n77 B 0.031266f
C239 VP.n78 B 0.031266f
C240 VP.n79 B 0.031266f
C241 VP.n80 B 0.062292f
C242 VP.n81 B 0.058273f
C243 VP.n82 B 0.041586f
C244 VP.n83 B 0.050463f
C245 VP.n84 B 0.08087f
.ends

