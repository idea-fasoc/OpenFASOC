* NGSPICE file created from diff_pair_sample_1463.ext - technology: sky130A

.subckt diff_pair_sample_1463 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=1.27
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=1.27
X2 VDD1.t3 VP.t1 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X3 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X4 VDD1.t2 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=1.27
X5 VDD1.t7 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=1.27
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=1.27
X7 VTAIL.t11 VP.t4 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=1.27
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=1.27
X9 VTAIL.t10 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X10 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X11 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=1.27
X12 VTAIL.t9 VP.t6 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X13 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=1.27
X14 VTAIL.t7 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X15 VDD1.t5 VP.t7 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X16 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=0.53955 ps=3.6 w=3.27 l=1.27
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0 ps=0 w=3.27 l=1.27
X18 VTAIL.t3 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2753 pd=7.32 as=0.53955 ps=3.6 w=3.27 l=1.27
X19 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.53955 pd=3.6 as=1.2753 ps=7.32 w=3.27 l=1.27
R0 VP.n11 VP.n10 161.3
R1 VP.n12 VP.n7 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n5 161.3
R5 VP.n32 VP.n0 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n29 VP.n28 161.3
R8 VP.n27 VP.n2 161.3
R9 VP.n26 VP.n25 161.3
R10 VP.n24 VP.n23 161.3
R11 VP.n22 VP.n4 161.3
R12 VP.n9 VP.t4 113.796
R13 VP.n21 VP.t0 93.1745
R14 VP.n33 VP.t2 93.1745
R15 VP.n18 VP.t3 93.1745
R16 VP.n19 VP.n18 80.6037
R17 VP.n34 VP.n33 80.6037
R18 VP.n21 VP.n20 80.6037
R19 VP.n3 VP.t7 62.0533
R20 VP.n1 VP.t5 62.0533
R21 VP.n6 VP.t6 62.0533
R22 VP.n8 VP.t1 62.0533
R23 VP.n9 VP.n8 42.5535
R24 VP.n27 VP.n26 40.4934
R25 VP.n28 VP.n27 40.4934
R26 VP.n13 VP.n12 40.4934
R27 VP.n12 VP.n11 40.4934
R28 VP.n22 VP.n21 38.7066
R29 VP.n33 VP.n32 38.7066
R30 VP.n18 VP.n17 38.7066
R31 VP.n20 VP.n19 38.2665
R32 VP.n23 VP.n22 30.7807
R33 VP.n32 VP.n31 30.7807
R34 VP.n17 VP.n16 30.7807
R35 VP.n10 VP.n9 29.0195
R36 VP.n26 VP.n3 14.6807
R37 VP.n28 VP.n1 14.6807
R38 VP.n13 VP.n6 14.6807
R39 VP.n11 VP.n8 14.6807
R40 VP.n23 VP.n3 9.7873
R41 VP.n31 VP.n1 9.7873
R42 VP.n16 VP.n6 9.7873
R43 VP.n19 VP.n5 0.285035
R44 VP.n20 VP.n4 0.285035
R45 VP.n34 VP.n0 0.285035
R46 VP.n10 VP.n7 0.189894
R47 VP.n14 VP.n7 0.189894
R48 VP.n15 VP.n14 0.189894
R49 VP.n15 VP.n5 0.189894
R50 VP.n24 VP.n4 0.189894
R51 VP.n25 VP.n24 0.189894
R52 VP.n25 VP.n2 0.189894
R53 VP.n29 VP.n2 0.189894
R54 VP.n30 VP.n29 0.189894
R55 VP.n30 VP.n0 0.189894
R56 VP VP.n34 0.146778
R57 VDD1 VDD1.n0 81.4061
R58 VDD1.n3 VDD1.n2 81.2925
R59 VDD1.n3 VDD1.n1 81.2925
R60 VDD1.n5 VDD1.n4 80.6582
R61 VDD1.n5 VDD1.n3 33.3242
R62 VDD1.n4 VDD1.t4 6.05555
R63 VDD1.n4 VDD1.t7 6.05555
R64 VDD1.n0 VDD1.t6 6.05555
R65 VDD1.n0 VDD1.t3 6.05555
R66 VDD1.n2 VDD1.t0 6.05555
R67 VDD1.n2 VDD1.t2 6.05555
R68 VDD1.n1 VDD1.t1 6.05555
R69 VDD1.n1 VDD1.t5 6.05555
R70 VDD1 VDD1.n5 0.631965
R71 VTAIL.n130 VTAIL.n120 289.615
R72 VTAIL.n12 VTAIL.n2 289.615
R73 VTAIL.n28 VTAIL.n18 289.615
R74 VTAIL.n46 VTAIL.n36 289.615
R75 VTAIL.n114 VTAIL.n104 289.615
R76 VTAIL.n96 VTAIL.n86 289.615
R77 VTAIL.n80 VTAIL.n70 289.615
R78 VTAIL.n62 VTAIL.n52 289.615
R79 VTAIL.n124 VTAIL.n123 185
R80 VTAIL.n129 VTAIL.n128 185
R81 VTAIL.n131 VTAIL.n130 185
R82 VTAIL.n6 VTAIL.n5 185
R83 VTAIL.n11 VTAIL.n10 185
R84 VTAIL.n13 VTAIL.n12 185
R85 VTAIL.n22 VTAIL.n21 185
R86 VTAIL.n27 VTAIL.n26 185
R87 VTAIL.n29 VTAIL.n28 185
R88 VTAIL.n40 VTAIL.n39 185
R89 VTAIL.n45 VTAIL.n44 185
R90 VTAIL.n47 VTAIL.n46 185
R91 VTAIL.n115 VTAIL.n114 185
R92 VTAIL.n113 VTAIL.n112 185
R93 VTAIL.n108 VTAIL.n107 185
R94 VTAIL.n97 VTAIL.n96 185
R95 VTAIL.n95 VTAIL.n94 185
R96 VTAIL.n90 VTAIL.n89 185
R97 VTAIL.n81 VTAIL.n80 185
R98 VTAIL.n79 VTAIL.n78 185
R99 VTAIL.n74 VTAIL.n73 185
R100 VTAIL.n63 VTAIL.n62 185
R101 VTAIL.n61 VTAIL.n60 185
R102 VTAIL.n56 VTAIL.n55 185
R103 VTAIL.n125 VTAIL.t4 148.606
R104 VTAIL.n7 VTAIL.t3 148.606
R105 VTAIL.n23 VTAIL.t13 148.606
R106 VTAIL.n41 VTAIL.t15 148.606
R107 VTAIL.n109 VTAIL.t12 148.606
R108 VTAIL.n91 VTAIL.t11 148.606
R109 VTAIL.n75 VTAIL.t5 148.606
R110 VTAIL.n57 VTAIL.t6 148.606
R111 VTAIL.n129 VTAIL.n123 104.615
R112 VTAIL.n130 VTAIL.n129 104.615
R113 VTAIL.n11 VTAIL.n5 104.615
R114 VTAIL.n12 VTAIL.n11 104.615
R115 VTAIL.n27 VTAIL.n21 104.615
R116 VTAIL.n28 VTAIL.n27 104.615
R117 VTAIL.n45 VTAIL.n39 104.615
R118 VTAIL.n46 VTAIL.n45 104.615
R119 VTAIL.n114 VTAIL.n113 104.615
R120 VTAIL.n113 VTAIL.n107 104.615
R121 VTAIL.n96 VTAIL.n95 104.615
R122 VTAIL.n95 VTAIL.n89 104.615
R123 VTAIL.n80 VTAIL.n79 104.615
R124 VTAIL.n79 VTAIL.n73 104.615
R125 VTAIL.n62 VTAIL.n61 104.615
R126 VTAIL.n61 VTAIL.n55 104.615
R127 VTAIL.n103 VTAIL.n102 63.9795
R128 VTAIL.n69 VTAIL.n68 63.9795
R129 VTAIL.n1 VTAIL.n0 63.9794
R130 VTAIL.n35 VTAIL.n34 63.9794
R131 VTAIL.t4 VTAIL.n123 52.3082
R132 VTAIL.t3 VTAIL.n5 52.3082
R133 VTAIL.t13 VTAIL.n21 52.3082
R134 VTAIL.t15 VTAIL.n39 52.3082
R135 VTAIL.t12 VTAIL.n107 52.3082
R136 VTAIL.t11 VTAIL.n89 52.3082
R137 VTAIL.t5 VTAIL.n73 52.3082
R138 VTAIL.t6 VTAIL.n55 52.3082
R139 VTAIL.n135 VTAIL.n134 35.0944
R140 VTAIL.n17 VTAIL.n16 35.0944
R141 VTAIL.n33 VTAIL.n32 35.0944
R142 VTAIL.n51 VTAIL.n50 35.0944
R143 VTAIL.n119 VTAIL.n118 35.0944
R144 VTAIL.n101 VTAIL.n100 35.0944
R145 VTAIL.n85 VTAIL.n84 35.0944
R146 VTAIL.n67 VTAIL.n66 35.0944
R147 VTAIL.n135 VTAIL.n119 16.5652
R148 VTAIL.n67 VTAIL.n51 16.5652
R149 VTAIL.n125 VTAIL.n124 15.5966
R150 VTAIL.n7 VTAIL.n6 15.5966
R151 VTAIL.n23 VTAIL.n22 15.5966
R152 VTAIL.n41 VTAIL.n40 15.5966
R153 VTAIL.n109 VTAIL.n108 15.5966
R154 VTAIL.n91 VTAIL.n90 15.5966
R155 VTAIL.n75 VTAIL.n74 15.5966
R156 VTAIL.n57 VTAIL.n56 15.5966
R157 VTAIL.n128 VTAIL.n127 12.8005
R158 VTAIL.n10 VTAIL.n9 12.8005
R159 VTAIL.n26 VTAIL.n25 12.8005
R160 VTAIL.n44 VTAIL.n43 12.8005
R161 VTAIL.n112 VTAIL.n111 12.8005
R162 VTAIL.n94 VTAIL.n93 12.8005
R163 VTAIL.n78 VTAIL.n77 12.8005
R164 VTAIL.n60 VTAIL.n59 12.8005
R165 VTAIL.n131 VTAIL.n122 12.0247
R166 VTAIL.n13 VTAIL.n4 12.0247
R167 VTAIL.n29 VTAIL.n20 12.0247
R168 VTAIL.n47 VTAIL.n38 12.0247
R169 VTAIL.n115 VTAIL.n106 12.0247
R170 VTAIL.n97 VTAIL.n88 12.0247
R171 VTAIL.n81 VTAIL.n72 12.0247
R172 VTAIL.n63 VTAIL.n54 12.0247
R173 VTAIL.n132 VTAIL.n120 11.249
R174 VTAIL.n14 VTAIL.n2 11.249
R175 VTAIL.n30 VTAIL.n18 11.249
R176 VTAIL.n48 VTAIL.n36 11.249
R177 VTAIL.n116 VTAIL.n104 11.249
R178 VTAIL.n98 VTAIL.n86 11.249
R179 VTAIL.n82 VTAIL.n70 11.249
R180 VTAIL.n64 VTAIL.n52 11.249
R181 VTAIL.n134 VTAIL.n133 9.45567
R182 VTAIL.n16 VTAIL.n15 9.45567
R183 VTAIL.n32 VTAIL.n31 9.45567
R184 VTAIL.n50 VTAIL.n49 9.45567
R185 VTAIL.n118 VTAIL.n117 9.45567
R186 VTAIL.n100 VTAIL.n99 9.45567
R187 VTAIL.n84 VTAIL.n83 9.45567
R188 VTAIL.n66 VTAIL.n65 9.45567
R189 VTAIL.n133 VTAIL.n132 9.3005
R190 VTAIL.n122 VTAIL.n121 9.3005
R191 VTAIL.n127 VTAIL.n126 9.3005
R192 VTAIL.n15 VTAIL.n14 9.3005
R193 VTAIL.n4 VTAIL.n3 9.3005
R194 VTAIL.n9 VTAIL.n8 9.3005
R195 VTAIL.n31 VTAIL.n30 9.3005
R196 VTAIL.n20 VTAIL.n19 9.3005
R197 VTAIL.n25 VTAIL.n24 9.3005
R198 VTAIL.n49 VTAIL.n48 9.3005
R199 VTAIL.n38 VTAIL.n37 9.3005
R200 VTAIL.n43 VTAIL.n42 9.3005
R201 VTAIL.n117 VTAIL.n116 9.3005
R202 VTAIL.n106 VTAIL.n105 9.3005
R203 VTAIL.n111 VTAIL.n110 9.3005
R204 VTAIL.n99 VTAIL.n98 9.3005
R205 VTAIL.n88 VTAIL.n87 9.3005
R206 VTAIL.n93 VTAIL.n92 9.3005
R207 VTAIL.n83 VTAIL.n82 9.3005
R208 VTAIL.n72 VTAIL.n71 9.3005
R209 VTAIL.n77 VTAIL.n76 9.3005
R210 VTAIL.n65 VTAIL.n64 9.3005
R211 VTAIL.n54 VTAIL.n53 9.3005
R212 VTAIL.n59 VTAIL.n58 9.3005
R213 VTAIL.n0 VTAIL.t2 6.05555
R214 VTAIL.n0 VTAIL.t7 6.05555
R215 VTAIL.n34 VTAIL.t8 6.05555
R216 VTAIL.n34 VTAIL.t10 6.05555
R217 VTAIL.n102 VTAIL.t14 6.05555
R218 VTAIL.n102 VTAIL.t9 6.05555
R219 VTAIL.n68 VTAIL.t0 6.05555
R220 VTAIL.n68 VTAIL.t1 6.05555
R221 VTAIL.n126 VTAIL.n125 4.46457
R222 VTAIL.n8 VTAIL.n7 4.46457
R223 VTAIL.n24 VTAIL.n23 4.46457
R224 VTAIL.n42 VTAIL.n41 4.46457
R225 VTAIL.n110 VTAIL.n109 4.46457
R226 VTAIL.n92 VTAIL.n91 4.46457
R227 VTAIL.n76 VTAIL.n75 4.46457
R228 VTAIL.n58 VTAIL.n57 4.46457
R229 VTAIL.n134 VTAIL.n120 2.71565
R230 VTAIL.n16 VTAIL.n2 2.71565
R231 VTAIL.n32 VTAIL.n18 2.71565
R232 VTAIL.n50 VTAIL.n36 2.71565
R233 VTAIL.n118 VTAIL.n104 2.71565
R234 VTAIL.n100 VTAIL.n86 2.71565
R235 VTAIL.n84 VTAIL.n70 2.71565
R236 VTAIL.n66 VTAIL.n52 2.71565
R237 VTAIL.n132 VTAIL.n131 1.93989
R238 VTAIL.n14 VTAIL.n13 1.93989
R239 VTAIL.n30 VTAIL.n29 1.93989
R240 VTAIL.n48 VTAIL.n47 1.93989
R241 VTAIL.n116 VTAIL.n115 1.93989
R242 VTAIL.n98 VTAIL.n97 1.93989
R243 VTAIL.n82 VTAIL.n81 1.93989
R244 VTAIL.n64 VTAIL.n63 1.93989
R245 VTAIL.n69 VTAIL.n67 1.37981
R246 VTAIL.n85 VTAIL.n69 1.37981
R247 VTAIL.n103 VTAIL.n101 1.37981
R248 VTAIL.n119 VTAIL.n103 1.37981
R249 VTAIL.n51 VTAIL.n35 1.37981
R250 VTAIL.n35 VTAIL.n33 1.37981
R251 VTAIL.n17 VTAIL.n1 1.37981
R252 VTAIL VTAIL.n135 1.32162
R253 VTAIL.n128 VTAIL.n122 1.16414
R254 VTAIL.n10 VTAIL.n4 1.16414
R255 VTAIL.n26 VTAIL.n20 1.16414
R256 VTAIL.n44 VTAIL.n38 1.16414
R257 VTAIL.n112 VTAIL.n106 1.16414
R258 VTAIL.n94 VTAIL.n88 1.16414
R259 VTAIL.n78 VTAIL.n72 1.16414
R260 VTAIL.n60 VTAIL.n54 1.16414
R261 VTAIL.n101 VTAIL.n85 0.470328
R262 VTAIL.n33 VTAIL.n17 0.470328
R263 VTAIL.n127 VTAIL.n124 0.388379
R264 VTAIL.n9 VTAIL.n6 0.388379
R265 VTAIL.n25 VTAIL.n22 0.388379
R266 VTAIL.n43 VTAIL.n40 0.388379
R267 VTAIL.n111 VTAIL.n108 0.388379
R268 VTAIL.n93 VTAIL.n90 0.388379
R269 VTAIL.n77 VTAIL.n74 0.388379
R270 VTAIL.n59 VTAIL.n56 0.388379
R271 VTAIL.n126 VTAIL.n121 0.155672
R272 VTAIL.n133 VTAIL.n121 0.155672
R273 VTAIL.n8 VTAIL.n3 0.155672
R274 VTAIL.n15 VTAIL.n3 0.155672
R275 VTAIL.n24 VTAIL.n19 0.155672
R276 VTAIL.n31 VTAIL.n19 0.155672
R277 VTAIL.n42 VTAIL.n37 0.155672
R278 VTAIL.n49 VTAIL.n37 0.155672
R279 VTAIL.n117 VTAIL.n105 0.155672
R280 VTAIL.n110 VTAIL.n105 0.155672
R281 VTAIL.n99 VTAIL.n87 0.155672
R282 VTAIL.n92 VTAIL.n87 0.155672
R283 VTAIL.n83 VTAIL.n71 0.155672
R284 VTAIL.n76 VTAIL.n71 0.155672
R285 VTAIL.n65 VTAIL.n53 0.155672
R286 VTAIL.n58 VTAIL.n53 0.155672
R287 VTAIL VTAIL.n1 0.0586897
R288 B.n467 B.n466 585
R289 B.n468 B.n467 585
R290 B.n162 B.n80 585
R291 B.n161 B.n160 585
R292 B.n159 B.n158 585
R293 B.n157 B.n156 585
R294 B.n155 B.n154 585
R295 B.n153 B.n152 585
R296 B.n151 B.n150 585
R297 B.n149 B.n148 585
R298 B.n147 B.n146 585
R299 B.n145 B.n144 585
R300 B.n143 B.n142 585
R301 B.n141 B.n140 585
R302 B.n139 B.n138 585
R303 B.n137 B.n136 585
R304 B.n135 B.n134 585
R305 B.n132 B.n131 585
R306 B.n130 B.n129 585
R307 B.n128 B.n127 585
R308 B.n126 B.n125 585
R309 B.n124 B.n123 585
R310 B.n122 B.n121 585
R311 B.n120 B.n119 585
R312 B.n118 B.n117 585
R313 B.n116 B.n115 585
R314 B.n114 B.n113 585
R315 B.n112 B.n111 585
R316 B.n110 B.n109 585
R317 B.n108 B.n107 585
R318 B.n106 B.n105 585
R319 B.n104 B.n103 585
R320 B.n102 B.n101 585
R321 B.n100 B.n99 585
R322 B.n98 B.n97 585
R323 B.n96 B.n95 585
R324 B.n94 B.n93 585
R325 B.n92 B.n91 585
R326 B.n90 B.n89 585
R327 B.n88 B.n87 585
R328 B.n60 B.n59 585
R329 B.n471 B.n470 585
R330 B.n465 B.n81 585
R331 B.n81 B.n57 585
R332 B.n464 B.n56 585
R333 B.n475 B.n56 585
R334 B.n463 B.n55 585
R335 B.n476 B.n55 585
R336 B.n462 B.n54 585
R337 B.n477 B.n54 585
R338 B.n461 B.n460 585
R339 B.n460 B.n50 585
R340 B.n459 B.n49 585
R341 B.n483 B.n49 585
R342 B.n458 B.n48 585
R343 B.n484 B.n48 585
R344 B.n457 B.n47 585
R345 B.n485 B.n47 585
R346 B.n456 B.n455 585
R347 B.n455 B.n43 585
R348 B.n454 B.n42 585
R349 B.n491 B.n42 585
R350 B.n453 B.n41 585
R351 B.n492 B.n41 585
R352 B.n452 B.n40 585
R353 B.n493 B.n40 585
R354 B.n451 B.n450 585
R355 B.n450 B.n36 585
R356 B.n449 B.n35 585
R357 B.n499 B.n35 585
R358 B.n448 B.n34 585
R359 B.n500 B.n34 585
R360 B.n447 B.n33 585
R361 B.n501 B.n33 585
R362 B.n446 B.n445 585
R363 B.n445 B.n29 585
R364 B.n444 B.n28 585
R365 B.n507 B.n28 585
R366 B.n443 B.n27 585
R367 B.n508 B.n27 585
R368 B.n442 B.n26 585
R369 B.n509 B.n26 585
R370 B.n441 B.n440 585
R371 B.n440 B.n22 585
R372 B.n439 B.n21 585
R373 B.n515 B.n21 585
R374 B.n438 B.n20 585
R375 B.n516 B.n20 585
R376 B.n437 B.n19 585
R377 B.n517 B.n19 585
R378 B.n436 B.n435 585
R379 B.n435 B.n15 585
R380 B.n434 B.n14 585
R381 B.n523 B.n14 585
R382 B.n433 B.n13 585
R383 B.n524 B.n13 585
R384 B.n432 B.n12 585
R385 B.n525 B.n12 585
R386 B.n431 B.n430 585
R387 B.n430 B.n429 585
R388 B.n428 B.n427 585
R389 B.n428 B.n8 585
R390 B.n426 B.n7 585
R391 B.n532 B.n7 585
R392 B.n425 B.n6 585
R393 B.n533 B.n6 585
R394 B.n424 B.n5 585
R395 B.n534 B.n5 585
R396 B.n423 B.n422 585
R397 B.n422 B.n4 585
R398 B.n421 B.n163 585
R399 B.n421 B.n420 585
R400 B.n411 B.n164 585
R401 B.n165 B.n164 585
R402 B.n413 B.n412 585
R403 B.n414 B.n413 585
R404 B.n410 B.n170 585
R405 B.n170 B.n169 585
R406 B.n409 B.n408 585
R407 B.n408 B.n407 585
R408 B.n172 B.n171 585
R409 B.n173 B.n172 585
R410 B.n400 B.n399 585
R411 B.n401 B.n400 585
R412 B.n398 B.n177 585
R413 B.n181 B.n177 585
R414 B.n397 B.n396 585
R415 B.n396 B.n395 585
R416 B.n179 B.n178 585
R417 B.n180 B.n179 585
R418 B.n388 B.n387 585
R419 B.n389 B.n388 585
R420 B.n386 B.n185 585
R421 B.n189 B.n185 585
R422 B.n385 B.n384 585
R423 B.n384 B.n383 585
R424 B.n187 B.n186 585
R425 B.n188 B.n187 585
R426 B.n376 B.n375 585
R427 B.n377 B.n376 585
R428 B.n374 B.n194 585
R429 B.n194 B.n193 585
R430 B.n373 B.n372 585
R431 B.n372 B.n371 585
R432 B.n196 B.n195 585
R433 B.n197 B.n196 585
R434 B.n364 B.n363 585
R435 B.n365 B.n364 585
R436 B.n362 B.n202 585
R437 B.n202 B.n201 585
R438 B.n361 B.n360 585
R439 B.n360 B.n359 585
R440 B.n204 B.n203 585
R441 B.n205 B.n204 585
R442 B.n352 B.n351 585
R443 B.n353 B.n352 585
R444 B.n350 B.n210 585
R445 B.n210 B.n209 585
R446 B.n349 B.n348 585
R447 B.n348 B.n347 585
R448 B.n212 B.n211 585
R449 B.n213 B.n212 585
R450 B.n340 B.n339 585
R451 B.n341 B.n340 585
R452 B.n338 B.n218 585
R453 B.n218 B.n217 585
R454 B.n337 B.n336 585
R455 B.n336 B.n335 585
R456 B.n220 B.n219 585
R457 B.n221 B.n220 585
R458 B.n331 B.n330 585
R459 B.n224 B.n223 585
R460 B.n327 B.n326 585
R461 B.n328 B.n327 585
R462 B.n325 B.n244 585
R463 B.n324 B.n323 585
R464 B.n322 B.n321 585
R465 B.n320 B.n319 585
R466 B.n318 B.n317 585
R467 B.n316 B.n315 585
R468 B.n314 B.n313 585
R469 B.n312 B.n311 585
R470 B.n310 B.n309 585
R471 B.n308 B.n307 585
R472 B.n306 B.n305 585
R473 B.n304 B.n303 585
R474 B.n302 B.n301 585
R475 B.n299 B.n298 585
R476 B.n297 B.n296 585
R477 B.n295 B.n294 585
R478 B.n293 B.n292 585
R479 B.n291 B.n290 585
R480 B.n289 B.n288 585
R481 B.n287 B.n286 585
R482 B.n285 B.n284 585
R483 B.n283 B.n282 585
R484 B.n281 B.n280 585
R485 B.n279 B.n278 585
R486 B.n277 B.n276 585
R487 B.n275 B.n274 585
R488 B.n273 B.n272 585
R489 B.n271 B.n270 585
R490 B.n269 B.n268 585
R491 B.n267 B.n266 585
R492 B.n265 B.n264 585
R493 B.n263 B.n262 585
R494 B.n261 B.n260 585
R495 B.n259 B.n258 585
R496 B.n257 B.n256 585
R497 B.n255 B.n254 585
R498 B.n253 B.n252 585
R499 B.n251 B.n250 585
R500 B.n332 B.n222 585
R501 B.n222 B.n221 585
R502 B.n334 B.n333 585
R503 B.n335 B.n334 585
R504 B.n216 B.n215 585
R505 B.n217 B.n216 585
R506 B.n343 B.n342 585
R507 B.n342 B.n341 585
R508 B.n344 B.n214 585
R509 B.n214 B.n213 585
R510 B.n346 B.n345 585
R511 B.n347 B.n346 585
R512 B.n208 B.n207 585
R513 B.n209 B.n208 585
R514 B.n355 B.n354 585
R515 B.n354 B.n353 585
R516 B.n356 B.n206 585
R517 B.n206 B.n205 585
R518 B.n358 B.n357 585
R519 B.n359 B.n358 585
R520 B.n200 B.n199 585
R521 B.n201 B.n200 585
R522 B.n367 B.n366 585
R523 B.n366 B.n365 585
R524 B.n368 B.n198 585
R525 B.n198 B.n197 585
R526 B.n370 B.n369 585
R527 B.n371 B.n370 585
R528 B.n192 B.n191 585
R529 B.n193 B.n192 585
R530 B.n379 B.n378 585
R531 B.n378 B.n377 585
R532 B.n380 B.n190 585
R533 B.n190 B.n188 585
R534 B.n382 B.n381 585
R535 B.n383 B.n382 585
R536 B.n184 B.n183 585
R537 B.n189 B.n184 585
R538 B.n391 B.n390 585
R539 B.n390 B.n389 585
R540 B.n392 B.n182 585
R541 B.n182 B.n180 585
R542 B.n394 B.n393 585
R543 B.n395 B.n394 585
R544 B.n176 B.n175 585
R545 B.n181 B.n176 585
R546 B.n403 B.n402 585
R547 B.n402 B.n401 585
R548 B.n404 B.n174 585
R549 B.n174 B.n173 585
R550 B.n406 B.n405 585
R551 B.n407 B.n406 585
R552 B.n168 B.n167 585
R553 B.n169 B.n168 585
R554 B.n416 B.n415 585
R555 B.n415 B.n414 585
R556 B.n417 B.n166 585
R557 B.n166 B.n165 585
R558 B.n419 B.n418 585
R559 B.n420 B.n419 585
R560 B.n3 B.n0 585
R561 B.n4 B.n3 585
R562 B.n531 B.n1 585
R563 B.n532 B.n531 585
R564 B.n530 B.n529 585
R565 B.n530 B.n8 585
R566 B.n528 B.n9 585
R567 B.n429 B.n9 585
R568 B.n527 B.n526 585
R569 B.n526 B.n525 585
R570 B.n11 B.n10 585
R571 B.n524 B.n11 585
R572 B.n522 B.n521 585
R573 B.n523 B.n522 585
R574 B.n520 B.n16 585
R575 B.n16 B.n15 585
R576 B.n519 B.n518 585
R577 B.n518 B.n517 585
R578 B.n18 B.n17 585
R579 B.n516 B.n18 585
R580 B.n514 B.n513 585
R581 B.n515 B.n514 585
R582 B.n512 B.n23 585
R583 B.n23 B.n22 585
R584 B.n511 B.n510 585
R585 B.n510 B.n509 585
R586 B.n25 B.n24 585
R587 B.n508 B.n25 585
R588 B.n506 B.n505 585
R589 B.n507 B.n506 585
R590 B.n504 B.n30 585
R591 B.n30 B.n29 585
R592 B.n503 B.n502 585
R593 B.n502 B.n501 585
R594 B.n32 B.n31 585
R595 B.n500 B.n32 585
R596 B.n498 B.n497 585
R597 B.n499 B.n498 585
R598 B.n496 B.n37 585
R599 B.n37 B.n36 585
R600 B.n495 B.n494 585
R601 B.n494 B.n493 585
R602 B.n39 B.n38 585
R603 B.n492 B.n39 585
R604 B.n490 B.n489 585
R605 B.n491 B.n490 585
R606 B.n488 B.n44 585
R607 B.n44 B.n43 585
R608 B.n487 B.n486 585
R609 B.n486 B.n485 585
R610 B.n46 B.n45 585
R611 B.n484 B.n46 585
R612 B.n482 B.n481 585
R613 B.n483 B.n482 585
R614 B.n480 B.n51 585
R615 B.n51 B.n50 585
R616 B.n479 B.n478 585
R617 B.n478 B.n477 585
R618 B.n53 B.n52 585
R619 B.n476 B.n53 585
R620 B.n474 B.n473 585
R621 B.n475 B.n474 585
R622 B.n472 B.n58 585
R623 B.n58 B.n57 585
R624 B.n535 B.n534 585
R625 B.n533 B.n2 585
R626 B.n470 B.n58 559.769
R627 B.n467 B.n81 559.769
R628 B.n250 B.n220 559.769
R629 B.n330 B.n222 559.769
R630 B.n84 B.t12 266.521
R631 B.n82 B.t19 266.521
R632 B.n247 B.t16 266.521
R633 B.n245 B.t8 266.521
R634 B.n468 B.n79 256.663
R635 B.n468 B.n78 256.663
R636 B.n468 B.n77 256.663
R637 B.n468 B.n76 256.663
R638 B.n468 B.n75 256.663
R639 B.n468 B.n74 256.663
R640 B.n468 B.n73 256.663
R641 B.n468 B.n72 256.663
R642 B.n468 B.n71 256.663
R643 B.n468 B.n70 256.663
R644 B.n468 B.n69 256.663
R645 B.n468 B.n68 256.663
R646 B.n468 B.n67 256.663
R647 B.n468 B.n66 256.663
R648 B.n468 B.n65 256.663
R649 B.n468 B.n64 256.663
R650 B.n468 B.n63 256.663
R651 B.n468 B.n62 256.663
R652 B.n468 B.n61 256.663
R653 B.n469 B.n468 256.663
R654 B.n329 B.n328 256.663
R655 B.n328 B.n225 256.663
R656 B.n328 B.n226 256.663
R657 B.n328 B.n227 256.663
R658 B.n328 B.n228 256.663
R659 B.n328 B.n229 256.663
R660 B.n328 B.n230 256.663
R661 B.n328 B.n231 256.663
R662 B.n328 B.n232 256.663
R663 B.n328 B.n233 256.663
R664 B.n328 B.n234 256.663
R665 B.n328 B.n235 256.663
R666 B.n328 B.n236 256.663
R667 B.n328 B.n237 256.663
R668 B.n328 B.n238 256.663
R669 B.n328 B.n239 256.663
R670 B.n328 B.n240 256.663
R671 B.n328 B.n241 256.663
R672 B.n328 B.n242 256.663
R673 B.n328 B.n243 256.663
R674 B.n537 B.n536 256.663
R675 B.n328 B.n221 171.212
R676 B.n468 B.n57 171.212
R677 B.n82 B.t20 164.567
R678 B.n247 B.t18 164.567
R679 B.n84 B.t14 164.567
R680 B.n245 B.t11 164.567
R681 B.n87 B.n60 163.367
R682 B.n91 B.n90 163.367
R683 B.n95 B.n94 163.367
R684 B.n99 B.n98 163.367
R685 B.n103 B.n102 163.367
R686 B.n107 B.n106 163.367
R687 B.n111 B.n110 163.367
R688 B.n115 B.n114 163.367
R689 B.n119 B.n118 163.367
R690 B.n123 B.n122 163.367
R691 B.n127 B.n126 163.367
R692 B.n131 B.n130 163.367
R693 B.n136 B.n135 163.367
R694 B.n140 B.n139 163.367
R695 B.n144 B.n143 163.367
R696 B.n148 B.n147 163.367
R697 B.n152 B.n151 163.367
R698 B.n156 B.n155 163.367
R699 B.n160 B.n159 163.367
R700 B.n467 B.n80 163.367
R701 B.n336 B.n220 163.367
R702 B.n336 B.n218 163.367
R703 B.n340 B.n218 163.367
R704 B.n340 B.n212 163.367
R705 B.n348 B.n212 163.367
R706 B.n348 B.n210 163.367
R707 B.n352 B.n210 163.367
R708 B.n352 B.n204 163.367
R709 B.n360 B.n204 163.367
R710 B.n360 B.n202 163.367
R711 B.n364 B.n202 163.367
R712 B.n364 B.n196 163.367
R713 B.n372 B.n196 163.367
R714 B.n372 B.n194 163.367
R715 B.n376 B.n194 163.367
R716 B.n376 B.n187 163.367
R717 B.n384 B.n187 163.367
R718 B.n384 B.n185 163.367
R719 B.n388 B.n185 163.367
R720 B.n388 B.n179 163.367
R721 B.n396 B.n179 163.367
R722 B.n396 B.n177 163.367
R723 B.n400 B.n177 163.367
R724 B.n400 B.n172 163.367
R725 B.n408 B.n172 163.367
R726 B.n408 B.n170 163.367
R727 B.n413 B.n170 163.367
R728 B.n413 B.n164 163.367
R729 B.n421 B.n164 163.367
R730 B.n422 B.n421 163.367
R731 B.n422 B.n5 163.367
R732 B.n6 B.n5 163.367
R733 B.n7 B.n6 163.367
R734 B.n428 B.n7 163.367
R735 B.n430 B.n428 163.367
R736 B.n430 B.n12 163.367
R737 B.n13 B.n12 163.367
R738 B.n14 B.n13 163.367
R739 B.n435 B.n14 163.367
R740 B.n435 B.n19 163.367
R741 B.n20 B.n19 163.367
R742 B.n21 B.n20 163.367
R743 B.n440 B.n21 163.367
R744 B.n440 B.n26 163.367
R745 B.n27 B.n26 163.367
R746 B.n28 B.n27 163.367
R747 B.n445 B.n28 163.367
R748 B.n445 B.n33 163.367
R749 B.n34 B.n33 163.367
R750 B.n35 B.n34 163.367
R751 B.n450 B.n35 163.367
R752 B.n450 B.n40 163.367
R753 B.n41 B.n40 163.367
R754 B.n42 B.n41 163.367
R755 B.n455 B.n42 163.367
R756 B.n455 B.n47 163.367
R757 B.n48 B.n47 163.367
R758 B.n49 B.n48 163.367
R759 B.n460 B.n49 163.367
R760 B.n460 B.n54 163.367
R761 B.n55 B.n54 163.367
R762 B.n56 B.n55 163.367
R763 B.n81 B.n56 163.367
R764 B.n327 B.n224 163.367
R765 B.n327 B.n244 163.367
R766 B.n323 B.n322 163.367
R767 B.n319 B.n318 163.367
R768 B.n315 B.n314 163.367
R769 B.n311 B.n310 163.367
R770 B.n307 B.n306 163.367
R771 B.n303 B.n302 163.367
R772 B.n298 B.n297 163.367
R773 B.n294 B.n293 163.367
R774 B.n290 B.n289 163.367
R775 B.n286 B.n285 163.367
R776 B.n282 B.n281 163.367
R777 B.n278 B.n277 163.367
R778 B.n274 B.n273 163.367
R779 B.n270 B.n269 163.367
R780 B.n266 B.n265 163.367
R781 B.n262 B.n261 163.367
R782 B.n258 B.n257 163.367
R783 B.n254 B.n253 163.367
R784 B.n334 B.n222 163.367
R785 B.n334 B.n216 163.367
R786 B.n342 B.n216 163.367
R787 B.n342 B.n214 163.367
R788 B.n346 B.n214 163.367
R789 B.n346 B.n208 163.367
R790 B.n354 B.n208 163.367
R791 B.n354 B.n206 163.367
R792 B.n358 B.n206 163.367
R793 B.n358 B.n200 163.367
R794 B.n366 B.n200 163.367
R795 B.n366 B.n198 163.367
R796 B.n370 B.n198 163.367
R797 B.n370 B.n192 163.367
R798 B.n378 B.n192 163.367
R799 B.n378 B.n190 163.367
R800 B.n382 B.n190 163.367
R801 B.n382 B.n184 163.367
R802 B.n390 B.n184 163.367
R803 B.n390 B.n182 163.367
R804 B.n394 B.n182 163.367
R805 B.n394 B.n176 163.367
R806 B.n402 B.n176 163.367
R807 B.n402 B.n174 163.367
R808 B.n406 B.n174 163.367
R809 B.n406 B.n168 163.367
R810 B.n415 B.n168 163.367
R811 B.n415 B.n166 163.367
R812 B.n419 B.n166 163.367
R813 B.n419 B.n3 163.367
R814 B.n535 B.n3 163.367
R815 B.n531 B.n2 163.367
R816 B.n531 B.n530 163.367
R817 B.n530 B.n9 163.367
R818 B.n526 B.n9 163.367
R819 B.n526 B.n11 163.367
R820 B.n522 B.n11 163.367
R821 B.n522 B.n16 163.367
R822 B.n518 B.n16 163.367
R823 B.n518 B.n18 163.367
R824 B.n514 B.n18 163.367
R825 B.n514 B.n23 163.367
R826 B.n510 B.n23 163.367
R827 B.n510 B.n25 163.367
R828 B.n506 B.n25 163.367
R829 B.n506 B.n30 163.367
R830 B.n502 B.n30 163.367
R831 B.n502 B.n32 163.367
R832 B.n498 B.n32 163.367
R833 B.n498 B.n37 163.367
R834 B.n494 B.n37 163.367
R835 B.n494 B.n39 163.367
R836 B.n490 B.n39 163.367
R837 B.n490 B.n44 163.367
R838 B.n486 B.n44 163.367
R839 B.n486 B.n46 163.367
R840 B.n482 B.n46 163.367
R841 B.n482 B.n51 163.367
R842 B.n478 B.n51 163.367
R843 B.n478 B.n53 163.367
R844 B.n474 B.n53 163.367
R845 B.n474 B.n58 163.367
R846 B.n83 B.t21 133.536
R847 B.n248 B.t17 133.536
R848 B.n85 B.t15 133.536
R849 B.n246 B.t10 133.536
R850 B.n335 B.n221 87.5371
R851 B.n335 B.n217 87.5371
R852 B.n341 B.n217 87.5371
R853 B.n341 B.n213 87.5371
R854 B.n347 B.n213 87.5371
R855 B.n353 B.n209 87.5371
R856 B.n353 B.n205 87.5371
R857 B.n359 B.n205 87.5371
R858 B.n359 B.n201 87.5371
R859 B.n365 B.n201 87.5371
R860 B.n365 B.n197 87.5371
R861 B.n371 B.n197 87.5371
R862 B.n377 B.n193 87.5371
R863 B.n377 B.n188 87.5371
R864 B.n383 B.n188 87.5371
R865 B.n383 B.n189 87.5371
R866 B.n389 B.n180 87.5371
R867 B.n395 B.n180 87.5371
R868 B.n395 B.n181 87.5371
R869 B.n401 B.n173 87.5371
R870 B.n407 B.n173 87.5371
R871 B.n407 B.n169 87.5371
R872 B.n414 B.n169 87.5371
R873 B.n420 B.n165 87.5371
R874 B.n420 B.n4 87.5371
R875 B.n534 B.n4 87.5371
R876 B.n534 B.n533 87.5371
R877 B.n533 B.n532 87.5371
R878 B.n532 B.n8 87.5371
R879 B.n429 B.n8 87.5371
R880 B.n525 B.n524 87.5371
R881 B.n524 B.n523 87.5371
R882 B.n523 B.n15 87.5371
R883 B.n517 B.n15 87.5371
R884 B.n516 B.n515 87.5371
R885 B.n515 B.n22 87.5371
R886 B.n509 B.n22 87.5371
R887 B.n508 B.n507 87.5371
R888 B.n507 B.n29 87.5371
R889 B.n501 B.n29 87.5371
R890 B.n501 B.n500 87.5371
R891 B.n499 B.n36 87.5371
R892 B.n493 B.n36 87.5371
R893 B.n493 B.n492 87.5371
R894 B.n492 B.n491 87.5371
R895 B.n491 B.n43 87.5371
R896 B.n485 B.n43 87.5371
R897 B.n485 B.n484 87.5371
R898 B.n483 B.n50 87.5371
R899 B.n477 B.n50 87.5371
R900 B.n477 B.n476 87.5371
R901 B.n476 B.n475 87.5371
R902 B.n475 B.n57 87.5371
R903 B.n389 B.t0 75.9514
R904 B.n509 B.t7 75.9514
R905 B.n181 B.t1 73.3767
R906 B.t2 B.n516 73.3767
R907 B.n470 B.n469 71.676
R908 B.n87 B.n61 71.676
R909 B.n91 B.n62 71.676
R910 B.n95 B.n63 71.676
R911 B.n99 B.n64 71.676
R912 B.n103 B.n65 71.676
R913 B.n107 B.n66 71.676
R914 B.n111 B.n67 71.676
R915 B.n115 B.n68 71.676
R916 B.n119 B.n69 71.676
R917 B.n123 B.n70 71.676
R918 B.n127 B.n71 71.676
R919 B.n131 B.n72 71.676
R920 B.n136 B.n73 71.676
R921 B.n140 B.n74 71.676
R922 B.n144 B.n75 71.676
R923 B.n148 B.n76 71.676
R924 B.n152 B.n77 71.676
R925 B.n156 B.n78 71.676
R926 B.n160 B.n79 71.676
R927 B.n80 B.n79 71.676
R928 B.n159 B.n78 71.676
R929 B.n155 B.n77 71.676
R930 B.n151 B.n76 71.676
R931 B.n147 B.n75 71.676
R932 B.n143 B.n74 71.676
R933 B.n139 B.n73 71.676
R934 B.n135 B.n72 71.676
R935 B.n130 B.n71 71.676
R936 B.n126 B.n70 71.676
R937 B.n122 B.n69 71.676
R938 B.n118 B.n68 71.676
R939 B.n114 B.n67 71.676
R940 B.n110 B.n66 71.676
R941 B.n106 B.n65 71.676
R942 B.n102 B.n64 71.676
R943 B.n98 B.n63 71.676
R944 B.n94 B.n62 71.676
R945 B.n90 B.n61 71.676
R946 B.n469 B.n60 71.676
R947 B.n330 B.n329 71.676
R948 B.n244 B.n225 71.676
R949 B.n322 B.n226 71.676
R950 B.n318 B.n227 71.676
R951 B.n314 B.n228 71.676
R952 B.n310 B.n229 71.676
R953 B.n306 B.n230 71.676
R954 B.n302 B.n231 71.676
R955 B.n297 B.n232 71.676
R956 B.n293 B.n233 71.676
R957 B.n289 B.n234 71.676
R958 B.n285 B.n235 71.676
R959 B.n281 B.n236 71.676
R960 B.n277 B.n237 71.676
R961 B.n273 B.n238 71.676
R962 B.n269 B.n239 71.676
R963 B.n265 B.n240 71.676
R964 B.n261 B.n241 71.676
R965 B.n257 B.n242 71.676
R966 B.n253 B.n243 71.676
R967 B.n329 B.n224 71.676
R968 B.n323 B.n225 71.676
R969 B.n319 B.n226 71.676
R970 B.n315 B.n227 71.676
R971 B.n311 B.n228 71.676
R972 B.n307 B.n229 71.676
R973 B.n303 B.n230 71.676
R974 B.n298 B.n231 71.676
R975 B.n294 B.n232 71.676
R976 B.n290 B.n233 71.676
R977 B.n286 B.n234 71.676
R978 B.n282 B.n235 71.676
R979 B.n278 B.n236 71.676
R980 B.n274 B.n237 71.676
R981 B.n270 B.n238 71.676
R982 B.n266 B.n239 71.676
R983 B.n262 B.n240 71.676
R984 B.n258 B.n241 71.676
R985 B.n254 B.n242 71.676
R986 B.n250 B.n243 71.676
R987 B.n536 B.n535 71.676
R988 B.n536 B.n2 71.676
R989 B.n86 B.n85 59.5399
R990 B.n133 B.n83 59.5399
R991 B.n249 B.n248 59.5399
R992 B.n300 B.n246 59.5399
R993 B.t6 B.n193 50.2053
R994 B.n500 B.t4 50.2053
R995 B.n414 B.t5 47.6307
R996 B.n525 B.t3 47.6307
R997 B.n347 B.t9 45.0561
R998 B.t13 B.n483 45.0561
R999 B.t9 B.n209 42.4815
R1000 B.n484 B.t13 42.4815
R1001 B.t5 B.n165 39.9069
R1002 B.n429 B.t3 39.9069
R1003 B.n371 B.t6 37.3323
R1004 B.t4 B.n499 37.3323
R1005 B.n332 B.n331 36.3712
R1006 B.n251 B.n219 36.3712
R1007 B.n472 B.n471 36.3712
R1008 B.n466 B.n465 36.3712
R1009 B.n85 B.n84 31.0308
R1010 B.n83 B.n82 31.0308
R1011 B.n248 B.n247 31.0308
R1012 B.n246 B.n245 31.0308
R1013 B B.n537 18.0485
R1014 B.n401 B.t1 14.1608
R1015 B.n517 B.t2 14.1608
R1016 B.n189 B.t0 11.5862
R1017 B.t7 B.n508 11.5862
R1018 B.n333 B.n332 10.6151
R1019 B.n333 B.n215 10.6151
R1020 B.n343 B.n215 10.6151
R1021 B.n344 B.n343 10.6151
R1022 B.n345 B.n344 10.6151
R1023 B.n345 B.n207 10.6151
R1024 B.n355 B.n207 10.6151
R1025 B.n356 B.n355 10.6151
R1026 B.n357 B.n356 10.6151
R1027 B.n357 B.n199 10.6151
R1028 B.n367 B.n199 10.6151
R1029 B.n368 B.n367 10.6151
R1030 B.n369 B.n368 10.6151
R1031 B.n369 B.n191 10.6151
R1032 B.n379 B.n191 10.6151
R1033 B.n380 B.n379 10.6151
R1034 B.n381 B.n380 10.6151
R1035 B.n381 B.n183 10.6151
R1036 B.n391 B.n183 10.6151
R1037 B.n392 B.n391 10.6151
R1038 B.n393 B.n392 10.6151
R1039 B.n393 B.n175 10.6151
R1040 B.n403 B.n175 10.6151
R1041 B.n404 B.n403 10.6151
R1042 B.n405 B.n404 10.6151
R1043 B.n405 B.n167 10.6151
R1044 B.n416 B.n167 10.6151
R1045 B.n417 B.n416 10.6151
R1046 B.n418 B.n417 10.6151
R1047 B.n418 B.n0 10.6151
R1048 B.n331 B.n223 10.6151
R1049 B.n326 B.n223 10.6151
R1050 B.n326 B.n325 10.6151
R1051 B.n325 B.n324 10.6151
R1052 B.n324 B.n321 10.6151
R1053 B.n321 B.n320 10.6151
R1054 B.n320 B.n317 10.6151
R1055 B.n317 B.n316 10.6151
R1056 B.n316 B.n313 10.6151
R1057 B.n313 B.n312 10.6151
R1058 B.n312 B.n309 10.6151
R1059 B.n309 B.n308 10.6151
R1060 B.n308 B.n305 10.6151
R1061 B.n305 B.n304 10.6151
R1062 B.n304 B.n301 10.6151
R1063 B.n299 B.n296 10.6151
R1064 B.n296 B.n295 10.6151
R1065 B.n295 B.n292 10.6151
R1066 B.n292 B.n291 10.6151
R1067 B.n291 B.n288 10.6151
R1068 B.n288 B.n287 10.6151
R1069 B.n287 B.n284 10.6151
R1070 B.n284 B.n283 10.6151
R1071 B.n280 B.n279 10.6151
R1072 B.n279 B.n276 10.6151
R1073 B.n276 B.n275 10.6151
R1074 B.n275 B.n272 10.6151
R1075 B.n272 B.n271 10.6151
R1076 B.n271 B.n268 10.6151
R1077 B.n268 B.n267 10.6151
R1078 B.n267 B.n264 10.6151
R1079 B.n264 B.n263 10.6151
R1080 B.n263 B.n260 10.6151
R1081 B.n260 B.n259 10.6151
R1082 B.n259 B.n256 10.6151
R1083 B.n256 B.n255 10.6151
R1084 B.n255 B.n252 10.6151
R1085 B.n252 B.n251 10.6151
R1086 B.n337 B.n219 10.6151
R1087 B.n338 B.n337 10.6151
R1088 B.n339 B.n338 10.6151
R1089 B.n339 B.n211 10.6151
R1090 B.n349 B.n211 10.6151
R1091 B.n350 B.n349 10.6151
R1092 B.n351 B.n350 10.6151
R1093 B.n351 B.n203 10.6151
R1094 B.n361 B.n203 10.6151
R1095 B.n362 B.n361 10.6151
R1096 B.n363 B.n362 10.6151
R1097 B.n363 B.n195 10.6151
R1098 B.n373 B.n195 10.6151
R1099 B.n374 B.n373 10.6151
R1100 B.n375 B.n374 10.6151
R1101 B.n375 B.n186 10.6151
R1102 B.n385 B.n186 10.6151
R1103 B.n386 B.n385 10.6151
R1104 B.n387 B.n386 10.6151
R1105 B.n387 B.n178 10.6151
R1106 B.n397 B.n178 10.6151
R1107 B.n398 B.n397 10.6151
R1108 B.n399 B.n398 10.6151
R1109 B.n399 B.n171 10.6151
R1110 B.n409 B.n171 10.6151
R1111 B.n410 B.n409 10.6151
R1112 B.n412 B.n410 10.6151
R1113 B.n412 B.n411 10.6151
R1114 B.n411 B.n163 10.6151
R1115 B.n423 B.n163 10.6151
R1116 B.n424 B.n423 10.6151
R1117 B.n425 B.n424 10.6151
R1118 B.n426 B.n425 10.6151
R1119 B.n427 B.n426 10.6151
R1120 B.n431 B.n427 10.6151
R1121 B.n432 B.n431 10.6151
R1122 B.n433 B.n432 10.6151
R1123 B.n434 B.n433 10.6151
R1124 B.n436 B.n434 10.6151
R1125 B.n437 B.n436 10.6151
R1126 B.n438 B.n437 10.6151
R1127 B.n439 B.n438 10.6151
R1128 B.n441 B.n439 10.6151
R1129 B.n442 B.n441 10.6151
R1130 B.n443 B.n442 10.6151
R1131 B.n444 B.n443 10.6151
R1132 B.n446 B.n444 10.6151
R1133 B.n447 B.n446 10.6151
R1134 B.n448 B.n447 10.6151
R1135 B.n449 B.n448 10.6151
R1136 B.n451 B.n449 10.6151
R1137 B.n452 B.n451 10.6151
R1138 B.n453 B.n452 10.6151
R1139 B.n454 B.n453 10.6151
R1140 B.n456 B.n454 10.6151
R1141 B.n457 B.n456 10.6151
R1142 B.n458 B.n457 10.6151
R1143 B.n459 B.n458 10.6151
R1144 B.n461 B.n459 10.6151
R1145 B.n462 B.n461 10.6151
R1146 B.n463 B.n462 10.6151
R1147 B.n464 B.n463 10.6151
R1148 B.n465 B.n464 10.6151
R1149 B.n529 B.n1 10.6151
R1150 B.n529 B.n528 10.6151
R1151 B.n528 B.n527 10.6151
R1152 B.n527 B.n10 10.6151
R1153 B.n521 B.n10 10.6151
R1154 B.n521 B.n520 10.6151
R1155 B.n520 B.n519 10.6151
R1156 B.n519 B.n17 10.6151
R1157 B.n513 B.n17 10.6151
R1158 B.n513 B.n512 10.6151
R1159 B.n512 B.n511 10.6151
R1160 B.n511 B.n24 10.6151
R1161 B.n505 B.n24 10.6151
R1162 B.n505 B.n504 10.6151
R1163 B.n504 B.n503 10.6151
R1164 B.n503 B.n31 10.6151
R1165 B.n497 B.n31 10.6151
R1166 B.n497 B.n496 10.6151
R1167 B.n496 B.n495 10.6151
R1168 B.n495 B.n38 10.6151
R1169 B.n489 B.n38 10.6151
R1170 B.n489 B.n488 10.6151
R1171 B.n488 B.n487 10.6151
R1172 B.n487 B.n45 10.6151
R1173 B.n481 B.n45 10.6151
R1174 B.n481 B.n480 10.6151
R1175 B.n480 B.n479 10.6151
R1176 B.n479 B.n52 10.6151
R1177 B.n473 B.n52 10.6151
R1178 B.n473 B.n472 10.6151
R1179 B.n471 B.n59 10.6151
R1180 B.n88 B.n59 10.6151
R1181 B.n89 B.n88 10.6151
R1182 B.n92 B.n89 10.6151
R1183 B.n93 B.n92 10.6151
R1184 B.n96 B.n93 10.6151
R1185 B.n97 B.n96 10.6151
R1186 B.n100 B.n97 10.6151
R1187 B.n101 B.n100 10.6151
R1188 B.n104 B.n101 10.6151
R1189 B.n105 B.n104 10.6151
R1190 B.n108 B.n105 10.6151
R1191 B.n109 B.n108 10.6151
R1192 B.n112 B.n109 10.6151
R1193 B.n113 B.n112 10.6151
R1194 B.n117 B.n116 10.6151
R1195 B.n120 B.n117 10.6151
R1196 B.n121 B.n120 10.6151
R1197 B.n124 B.n121 10.6151
R1198 B.n125 B.n124 10.6151
R1199 B.n128 B.n125 10.6151
R1200 B.n129 B.n128 10.6151
R1201 B.n132 B.n129 10.6151
R1202 B.n137 B.n134 10.6151
R1203 B.n138 B.n137 10.6151
R1204 B.n141 B.n138 10.6151
R1205 B.n142 B.n141 10.6151
R1206 B.n145 B.n142 10.6151
R1207 B.n146 B.n145 10.6151
R1208 B.n149 B.n146 10.6151
R1209 B.n150 B.n149 10.6151
R1210 B.n153 B.n150 10.6151
R1211 B.n154 B.n153 10.6151
R1212 B.n157 B.n154 10.6151
R1213 B.n158 B.n157 10.6151
R1214 B.n161 B.n158 10.6151
R1215 B.n162 B.n161 10.6151
R1216 B.n466 B.n162 10.6151
R1217 B.n537 B.n0 8.11757
R1218 B.n537 B.n1 8.11757
R1219 B.n300 B.n299 6.5566
R1220 B.n283 B.n249 6.5566
R1221 B.n116 B.n86 6.5566
R1222 B.n133 B.n132 6.5566
R1223 B.n301 B.n300 4.05904
R1224 B.n280 B.n249 4.05904
R1225 B.n113 B.n86 4.05904
R1226 B.n134 B.n133 4.05904
R1227 VN.n27 VN.n15 161.3
R1228 VN.n26 VN.n25 161.3
R1229 VN.n24 VN.n23 161.3
R1230 VN.n22 VN.n17 161.3
R1231 VN.n21 VN.n20 161.3
R1232 VN.n12 VN.n0 161.3
R1233 VN.n11 VN.n10 161.3
R1234 VN.n9 VN.n8 161.3
R1235 VN.n7 VN.n2 161.3
R1236 VN.n6 VN.n5 161.3
R1237 VN.n4 VN.t6 113.796
R1238 VN.n19 VN.t2 113.796
R1239 VN.n13 VN.t7 93.1745
R1240 VN.n28 VN.t3 93.1745
R1241 VN.n29 VN.n28 80.6037
R1242 VN.n14 VN.n13 80.6037
R1243 VN.n3 VN.t1 62.0533
R1244 VN.n1 VN.t4 62.0533
R1245 VN.n18 VN.t0 62.0533
R1246 VN.n16 VN.t5 62.0533
R1247 VN.n4 VN.n3 42.5535
R1248 VN.n19 VN.n18 42.5535
R1249 VN.n7 VN.n6 40.4934
R1250 VN.n8 VN.n7 40.4934
R1251 VN.n22 VN.n21 40.4934
R1252 VN.n23 VN.n22 40.4934
R1253 VN.n13 VN.n12 38.7066
R1254 VN.n28 VN.n27 38.7066
R1255 VN VN.n29 38.5521
R1256 VN.n12 VN.n11 30.7807
R1257 VN.n27 VN.n26 30.7807
R1258 VN.n20 VN.n19 29.0195
R1259 VN.n5 VN.n4 29.0195
R1260 VN.n6 VN.n3 14.6807
R1261 VN.n8 VN.n1 14.6807
R1262 VN.n21 VN.n18 14.6807
R1263 VN.n23 VN.n16 14.6807
R1264 VN.n11 VN.n1 9.7873
R1265 VN.n26 VN.n16 9.7873
R1266 VN.n29 VN.n15 0.285035
R1267 VN.n14 VN.n0 0.285035
R1268 VN.n25 VN.n15 0.189894
R1269 VN.n25 VN.n24 0.189894
R1270 VN.n24 VN.n17 0.189894
R1271 VN.n20 VN.n17 0.189894
R1272 VN.n5 VN.n2 0.189894
R1273 VN.n9 VN.n2 0.189894
R1274 VN.n10 VN.n9 0.189894
R1275 VN.n10 VN.n0 0.189894
R1276 VN VN.n14 0.146778
R1277 VDD2.n2 VDD2.n1 81.2925
R1278 VDD2.n2 VDD2.n0 81.2925
R1279 VDD2 VDD2.n5 81.2896
R1280 VDD2.n4 VDD2.n3 80.6583
R1281 VDD2.n4 VDD2.n2 32.7412
R1282 VDD2.n5 VDD2.t7 6.05555
R1283 VDD2.n5 VDD2.t5 6.05555
R1284 VDD2.n3 VDD2.t4 6.05555
R1285 VDD2.n3 VDD2.t2 6.05555
R1286 VDD2.n1 VDD2.t3 6.05555
R1287 VDD2.n1 VDD2.t0 6.05555
R1288 VDD2.n0 VDD2.t1 6.05555
R1289 VDD2.n0 VDD2.t6 6.05555
R1290 VDD2 VDD2.n4 0.748345
C0 VP VDD1 2.47938f
C1 VDD1 VDD2 1.11077f
C2 VP VTAIL 2.70978f
C3 VDD1 VN 0.153897f
C4 VTAIL VDD2 4.40671f
C5 VP VDD2 0.383261f
C6 VTAIL VN 2.69567f
C7 VP VN 4.42246f
C8 VN VDD2 2.25133f
C9 VTAIL VDD1 4.36121f
C10 VDD2 B 3.334462f
C11 VDD1 B 3.634264f
C12 VTAIL B 4.152266f
C13 VN B 9.612399f
C14 VP B 8.126328f
C15 VDD2.t1 B 0.064756f
C16 VDD2.t6 B 0.064756f
C17 VDD2.n0 B 0.491532f
C18 VDD2.t3 B 0.064756f
C19 VDD2.t0 B 0.064756f
C20 VDD2.n1 B 0.491532f
C21 VDD2.n2 B 1.95907f
C22 VDD2.t4 B 0.064756f
C23 VDD2.t2 B 0.064756f
C24 VDD2.n3 B 0.488687f
C25 VDD2.n4 B 1.78736f
C26 VDD2.t7 B 0.064756f
C27 VDD2.t5 B 0.064756f
C28 VDD2.n5 B 0.49151f
C29 VN.n0 B 0.050629f
C30 VN.t4 B 0.396567f
C31 VN.n1 B 0.182105f
C32 VN.n2 B 0.037942f
C33 VN.t1 B 0.396567f
C34 VN.n3 B 0.234406f
C35 VN.t6 B 0.518843f
C36 VN.n4 B 0.245534f
C37 VN.n5 B 0.201186f
C38 VN.n6 B 0.061444f
C39 VN.n7 B 0.030672f
C40 VN.n8 B 0.061444f
C41 VN.n9 B 0.037942f
C42 VN.n10 B 0.037942f
C43 VN.n11 B 0.055063f
C44 VN.n12 B 0.030665f
C45 VN.t7 B 0.470388f
C46 VN.n13 B 0.258703f
C47 VN.n14 B 0.035534f
C48 VN.n15 B 0.050629f
C49 VN.t5 B 0.396567f
C50 VN.n16 B 0.182105f
C51 VN.n17 B 0.037942f
C52 VN.t0 B 0.396567f
C53 VN.n18 B 0.234406f
C54 VN.t2 B 0.518843f
C55 VN.n19 B 0.245534f
C56 VN.n20 B 0.201186f
C57 VN.n21 B 0.061444f
C58 VN.n22 B 0.030672f
C59 VN.n23 B 0.061444f
C60 VN.n24 B 0.037942f
C61 VN.n25 B 0.037942f
C62 VN.n26 B 0.055063f
C63 VN.n27 B 0.030665f
C64 VN.t3 B 0.470388f
C65 VN.n28 B 0.258703f
C66 VN.n29 B 1.36912f
C67 VTAIL.t2 B 0.064156f
C68 VTAIL.t7 B 0.064156f
C69 VTAIL.n0 B 0.435993f
C70 VTAIL.n1 B 0.318893f
C71 VTAIL.n2 B 0.03473f
C72 VTAIL.n3 B 0.024828f
C73 VTAIL.n4 B 0.013341f
C74 VTAIL.n5 B 0.023651f
C75 VTAIL.n6 B 0.018388f
C76 VTAIL.t3 B 0.053515f
C77 VTAIL.n7 B 0.092923f
C78 VTAIL.n8 B 0.274333f
C79 VTAIL.n9 B 0.013341f
C80 VTAIL.n10 B 0.014126f
C81 VTAIL.n11 B 0.031534f
C82 VTAIL.n12 B 0.06797f
C83 VTAIL.n13 B 0.014126f
C84 VTAIL.n14 B 0.013341f
C85 VTAIL.n15 B 0.062476f
C86 VTAIL.n16 B 0.038152f
C87 VTAIL.n17 B 0.172014f
C88 VTAIL.n18 B 0.03473f
C89 VTAIL.n19 B 0.024828f
C90 VTAIL.n20 B 0.013341f
C91 VTAIL.n21 B 0.023651f
C92 VTAIL.n22 B 0.018388f
C93 VTAIL.t13 B 0.053515f
C94 VTAIL.n23 B 0.092923f
C95 VTAIL.n24 B 0.274333f
C96 VTAIL.n25 B 0.013341f
C97 VTAIL.n26 B 0.014126f
C98 VTAIL.n27 B 0.031534f
C99 VTAIL.n28 B 0.06797f
C100 VTAIL.n29 B 0.014126f
C101 VTAIL.n30 B 0.013341f
C102 VTAIL.n31 B 0.062476f
C103 VTAIL.n32 B 0.038152f
C104 VTAIL.n33 B 0.172014f
C105 VTAIL.t8 B 0.064156f
C106 VTAIL.t10 B 0.064156f
C107 VTAIL.n34 B 0.435993f
C108 VTAIL.n35 B 0.424584f
C109 VTAIL.n36 B 0.03473f
C110 VTAIL.n37 B 0.024828f
C111 VTAIL.n38 B 0.013341f
C112 VTAIL.n39 B 0.023651f
C113 VTAIL.n40 B 0.018388f
C114 VTAIL.t15 B 0.053515f
C115 VTAIL.n41 B 0.092923f
C116 VTAIL.n42 B 0.274333f
C117 VTAIL.n43 B 0.013341f
C118 VTAIL.n44 B 0.014126f
C119 VTAIL.n45 B 0.031534f
C120 VTAIL.n46 B 0.06797f
C121 VTAIL.n47 B 0.014126f
C122 VTAIL.n48 B 0.013341f
C123 VTAIL.n49 B 0.062476f
C124 VTAIL.n50 B 0.038152f
C125 VTAIL.n51 B 0.807548f
C126 VTAIL.n52 B 0.03473f
C127 VTAIL.n53 B 0.024828f
C128 VTAIL.n54 B 0.013341f
C129 VTAIL.n55 B 0.023651f
C130 VTAIL.n56 B 0.018388f
C131 VTAIL.t6 B 0.053515f
C132 VTAIL.n57 B 0.092923f
C133 VTAIL.n58 B 0.274333f
C134 VTAIL.n59 B 0.013341f
C135 VTAIL.n60 B 0.014126f
C136 VTAIL.n61 B 0.031534f
C137 VTAIL.n62 B 0.06797f
C138 VTAIL.n63 B 0.014126f
C139 VTAIL.n64 B 0.013341f
C140 VTAIL.n65 B 0.062476f
C141 VTAIL.n66 B 0.038152f
C142 VTAIL.n67 B 0.807548f
C143 VTAIL.t0 B 0.064156f
C144 VTAIL.t1 B 0.064156f
C145 VTAIL.n68 B 0.435996f
C146 VTAIL.n69 B 0.424581f
C147 VTAIL.n70 B 0.03473f
C148 VTAIL.n71 B 0.024828f
C149 VTAIL.n72 B 0.013341f
C150 VTAIL.n73 B 0.023651f
C151 VTAIL.n74 B 0.018388f
C152 VTAIL.t5 B 0.053515f
C153 VTAIL.n75 B 0.092923f
C154 VTAIL.n76 B 0.274333f
C155 VTAIL.n77 B 0.013341f
C156 VTAIL.n78 B 0.014126f
C157 VTAIL.n79 B 0.031534f
C158 VTAIL.n80 B 0.06797f
C159 VTAIL.n81 B 0.014126f
C160 VTAIL.n82 B 0.013341f
C161 VTAIL.n83 B 0.062476f
C162 VTAIL.n84 B 0.038152f
C163 VTAIL.n85 B 0.172014f
C164 VTAIL.n86 B 0.03473f
C165 VTAIL.n87 B 0.024828f
C166 VTAIL.n88 B 0.013341f
C167 VTAIL.n89 B 0.023651f
C168 VTAIL.n90 B 0.018388f
C169 VTAIL.t11 B 0.053515f
C170 VTAIL.n91 B 0.092923f
C171 VTAIL.n92 B 0.274333f
C172 VTAIL.n93 B 0.013341f
C173 VTAIL.n94 B 0.014126f
C174 VTAIL.n95 B 0.031534f
C175 VTAIL.n96 B 0.06797f
C176 VTAIL.n97 B 0.014126f
C177 VTAIL.n98 B 0.013341f
C178 VTAIL.n99 B 0.062476f
C179 VTAIL.n100 B 0.038152f
C180 VTAIL.n101 B 0.172014f
C181 VTAIL.t14 B 0.064156f
C182 VTAIL.t9 B 0.064156f
C183 VTAIL.n102 B 0.435996f
C184 VTAIL.n103 B 0.424581f
C185 VTAIL.n104 B 0.03473f
C186 VTAIL.n105 B 0.024828f
C187 VTAIL.n106 B 0.013341f
C188 VTAIL.n107 B 0.023651f
C189 VTAIL.n108 B 0.018388f
C190 VTAIL.t12 B 0.053515f
C191 VTAIL.n109 B 0.092923f
C192 VTAIL.n110 B 0.274333f
C193 VTAIL.n111 B 0.013341f
C194 VTAIL.n112 B 0.014126f
C195 VTAIL.n113 B 0.031534f
C196 VTAIL.n114 B 0.06797f
C197 VTAIL.n115 B 0.014126f
C198 VTAIL.n116 B 0.013341f
C199 VTAIL.n117 B 0.062476f
C200 VTAIL.n118 B 0.038152f
C201 VTAIL.n119 B 0.807548f
C202 VTAIL.n120 B 0.03473f
C203 VTAIL.n121 B 0.024828f
C204 VTAIL.n122 B 0.013341f
C205 VTAIL.n123 B 0.023651f
C206 VTAIL.n124 B 0.018388f
C207 VTAIL.t4 B 0.053515f
C208 VTAIL.n125 B 0.092923f
C209 VTAIL.n126 B 0.274333f
C210 VTAIL.n127 B 0.013341f
C211 VTAIL.n128 B 0.014126f
C212 VTAIL.n129 B 0.031534f
C213 VTAIL.n130 B 0.06797f
C214 VTAIL.n131 B 0.014126f
C215 VTAIL.n132 B 0.013341f
C216 VTAIL.n133 B 0.062476f
C217 VTAIL.n134 B 0.038152f
C218 VTAIL.n135 B 0.802892f
C219 VDD1.t6 B 0.065781f
C220 VDD1.t3 B 0.065781f
C221 VDD1.n0 B 0.499898f
C222 VDD1.t1 B 0.065781f
C223 VDD1.t5 B 0.065781f
C224 VDD1.n1 B 0.499306f
C225 VDD1.t0 B 0.065781f
C226 VDD1.t2 B 0.065781f
C227 VDD1.n2 B 0.499306f
C228 VDD1.n3 B 2.04418f
C229 VDD1.t4 B 0.065781f
C230 VDD1.t7 B 0.065781f
C231 VDD1.n4 B 0.496414f
C232 VDD1.n5 B 1.84598f
C233 VP.n0 B 0.052001f
C234 VP.t5 B 0.407315f
C235 VP.n1 B 0.187041f
C236 VP.n2 B 0.03897f
C237 VP.t7 B 0.407315f
C238 VP.n3 B 0.187041f
C239 VP.n4 B 0.052001f
C240 VP.n5 B 0.052001f
C241 VP.t3 B 0.483138f
C242 VP.t6 B 0.407315f
C243 VP.n6 B 0.187041f
C244 VP.n7 B 0.03897f
C245 VP.t1 B 0.407315f
C246 VP.n8 B 0.240759f
C247 VP.t4 B 0.532906f
C248 VP.n9 B 0.252189f
C249 VP.n10 B 0.206639f
C250 VP.n11 B 0.06311f
C251 VP.n12 B 0.031504f
C252 VP.n13 B 0.06311f
C253 VP.n14 B 0.03897f
C254 VP.n15 B 0.03897f
C255 VP.n16 B 0.056556f
C256 VP.n17 B 0.031496f
C257 VP.n18 B 0.265715f
C258 VP.n19 B 1.38399f
C259 VP.n20 B 1.4206f
C260 VP.t0 B 0.483138f
C261 VP.n21 B 0.265715f
C262 VP.n22 B 0.031496f
C263 VP.n23 B 0.056556f
C264 VP.n24 B 0.03897f
C265 VP.n25 B 0.03897f
C266 VP.n26 B 0.06311f
C267 VP.n27 B 0.031504f
C268 VP.n28 B 0.06311f
C269 VP.n29 B 0.03897f
C270 VP.n30 B 0.03897f
C271 VP.n31 B 0.056556f
C272 VP.n32 B 0.031496f
C273 VP.t2 B 0.483138f
C274 VP.n33 B 0.265715f
C275 VP.n34 B 0.036497f
.ends

