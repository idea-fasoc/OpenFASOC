* NGSPICE file created from diff_pair_sample_0056.ext - technology: sky130A

.subckt diff_pair_sample_0056 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=1.64
X1 VDD2.t3 VN.t0 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=1.64
X2 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=1.64
X3 VTAIL.t5 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=1.64
X4 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=1.64
X5 VTAIL.t4 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=1.64
X6 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=1.64
X7 VDD1.t0 VP.t3 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=1.64
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=1.64
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=1.64
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=1.64
X11 VTAIL.t7 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=1.64
R0 VP.n4 VP.n3 174.334
R1 VP.n12 VP.n11 174.334
R2 VP.n10 VP.n0 161.3
R3 VP.n9 VP.n8 161.3
R4 VP.n7 VP.n1 161.3
R5 VP.n6 VP.n5 161.3
R6 VP.n2 VP.t2 136.898
R7 VP.n2 VP.t0 136.569
R8 VP.n4 VP.t1 98.4578
R9 VP.n11 VP.t3 98.4578
R10 VP.n9 VP.n1 56.5617
R11 VP.n3 VP.n2 51.8858
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 11.5587
R15 VP.n11 VP.n10 11.5587
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VTAIL.n282 VTAIL.n252 289.615
R23 VTAIL.n30 VTAIL.n0 289.615
R24 VTAIL.n66 VTAIL.n36 289.615
R25 VTAIL.n102 VTAIL.n72 289.615
R26 VTAIL.n246 VTAIL.n216 289.615
R27 VTAIL.n210 VTAIL.n180 289.615
R28 VTAIL.n174 VTAIL.n144 289.615
R29 VTAIL.n138 VTAIL.n108 289.615
R30 VTAIL.n265 VTAIL.n264 185
R31 VTAIL.n267 VTAIL.n266 185
R32 VTAIL.n260 VTAIL.n259 185
R33 VTAIL.n273 VTAIL.n272 185
R34 VTAIL.n275 VTAIL.n274 185
R35 VTAIL.n256 VTAIL.n255 185
R36 VTAIL.n281 VTAIL.n280 185
R37 VTAIL.n283 VTAIL.n282 185
R38 VTAIL.n13 VTAIL.n12 185
R39 VTAIL.n15 VTAIL.n14 185
R40 VTAIL.n8 VTAIL.n7 185
R41 VTAIL.n21 VTAIL.n20 185
R42 VTAIL.n23 VTAIL.n22 185
R43 VTAIL.n4 VTAIL.n3 185
R44 VTAIL.n29 VTAIL.n28 185
R45 VTAIL.n31 VTAIL.n30 185
R46 VTAIL.n49 VTAIL.n48 185
R47 VTAIL.n51 VTAIL.n50 185
R48 VTAIL.n44 VTAIL.n43 185
R49 VTAIL.n57 VTAIL.n56 185
R50 VTAIL.n59 VTAIL.n58 185
R51 VTAIL.n40 VTAIL.n39 185
R52 VTAIL.n65 VTAIL.n64 185
R53 VTAIL.n67 VTAIL.n66 185
R54 VTAIL.n85 VTAIL.n84 185
R55 VTAIL.n87 VTAIL.n86 185
R56 VTAIL.n80 VTAIL.n79 185
R57 VTAIL.n93 VTAIL.n92 185
R58 VTAIL.n95 VTAIL.n94 185
R59 VTAIL.n76 VTAIL.n75 185
R60 VTAIL.n101 VTAIL.n100 185
R61 VTAIL.n103 VTAIL.n102 185
R62 VTAIL.n247 VTAIL.n246 185
R63 VTAIL.n245 VTAIL.n244 185
R64 VTAIL.n220 VTAIL.n219 185
R65 VTAIL.n239 VTAIL.n238 185
R66 VTAIL.n237 VTAIL.n236 185
R67 VTAIL.n224 VTAIL.n223 185
R68 VTAIL.n231 VTAIL.n230 185
R69 VTAIL.n229 VTAIL.n228 185
R70 VTAIL.n211 VTAIL.n210 185
R71 VTAIL.n209 VTAIL.n208 185
R72 VTAIL.n184 VTAIL.n183 185
R73 VTAIL.n203 VTAIL.n202 185
R74 VTAIL.n201 VTAIL.n200 185
R75 VTAIL.n188 VTAIL.n187 185
R76 VTAIL.n195 VTAIL.n194 185
R77 VTAIL.n193 VTAIL.n192 185
R78 VTAIL.n175 VTAIL.n174 185
R79 VTAIL.n173 VTAIL.n172 185
R80 VTAIL.n148 VTAIL.n147 185
R81 VTAIL.n167 VTAIL.n166 185
R82 VTAIL.n165 VTAIL.n164 185
R83 VTAIL.n152 VTAIL.n151 185
R84 VTAIL.n159 VTAIL.n158 185
R85 VTAIL.n157 VTAIL.n156 185
R86 VTAIL.n139 VTAIL.n138 185
R87 VTAIL.n137 VTAIL.n136 185
R88 VTAIL.n112 VTAIL.n111 185
R89 VTAIL.n131 VTAIL.n130 185
R90 VTAIL.n129 VTAIL.n128 185
R91 VTAIL.n116 VTAIL.n115 185
R92 VTAIL.n123 VTAIL.n122 185
R93 VTAIL.n121 VTAIL.n120 185
R94 VTAIL.n263 VTAIL.t6 147.659
R95 VTAIL.n11 VTAIL.t7 147.659
R96 VTAIL.n47 VTAIL.t2 147.659
R97 VTAIL.n83 VTAIL.t5 147.659
R98 VTAIL.n227 VTAIL.t3 147.659
R99 VTAIL.n191 VTAIL.t4 147.659
R100 VTAIL.n155 VTAIL.t0 147.659
R101 VTAIL.n119 VTAIL.t1 147.659
R102 VTAIL.n266 VTAIL.n265 104.615
R103 VTAIL.n266 VTAIL.n259 104.615
R104 VTAIL.n273 VTAIL.n259 104.615
R105 VTAIL.n274 VTAIL.n273 104.615
R106 VTAIL.n274 VTAIL.n255 104.615
R107 VTAIL.n281 VTAIL.n255 104.615
R108 VTAIL.n282 VTAIL.n281 104.615
R109 VTAIL.n14 VTAIL.n13 104.615
R110 VTAIL.n14 VTAIL.n7 104.615
R111 VTAIL.n21 VTAIL.n7 104.615
R112 VTAIL.n22 VTAIL.n21 104.615
R113 VTAIL.n22 VTAIL.n3 104.615
R114 VTAIL.n29 VTAIL.n3 104.615
R115 VTAIL.n30 VTAIL.n29 104.615
R116 VTAIL.n50 VTAIL.n49 104.615
R117 VTAIL.n50 VTAIL.n43 104.615
R118 VTAIL.n57 VTAIL.n43 104.615
R119 VTAIL.n58 VTAIL.n57 104.615
R120 VTAIL.n58 VTAIL.n39 104.615
R121 VTAIL.n65 VTAIL.n39 104.615
R122 VTAIL.n66 VTAIL.n65 104.615
R123 VTAIL.n86 VTAIL.n85 104.615
R124 VTAIL.n86 VTAIL.n79 104.615
R125 VTAIL.n93 VTAIL.n79 104.615
R126 VTAIL.n94 VTAIL.n93 104.615
R127 VTAIL.n94 VTAIL.n75 104.615
R128 VTAIL.n101 VTAIL.n75 104.615
R129 VTAIL.n102 VTAIL.n101 104.615
R130 VTAIL.n246 VTAIL.n245 104.615
R131 VTAIL.n245 VTAIL.n219 104.615
R132 VTAIL.n238 VTAIL.n219 104.615
R133 VTAIL.n238 VTAIL.n237 104.615
R134 VTAIL.n237 VTAIL.n223 104.615
R135 VTAIL.n230 VTAIL.n223 104.615
R136 VTAIL.n230 VTAIL.n229 104.615
R137 VTAIL.n210 VTAIL.n209 104.615
R138 VTAIL.n209 VTAIL.n183 104.615
R139 VTAIL.n202 VTAIL.n183 104.615
R140 VTAIL.n202 VTAIL.n201 104.615
R141 VTAIL.n201 VTAIL.n187 104.615
R142 VTAIL.n194 VTAIL.n187 104.615
R143 VTAIL.n194 VTAIL.n193 104.615
R144 VTAIL.n174 VTAIL.n173 104.615
R145 VTAIL.n173 VTAIL.n147 104.615
R146 VTAIL.n166 VTAIL.n147 104.615
R147 VTAIL.n166 VTAIL.n165 104.615
R148 VTAIL.n165 VTAIL.n151 104.615
R149 VTAIL.n158 VTAIL.n151 104.615
R150 VTAIL.n158 VTAIL.n157 104.615
R151 VTAIL.n138 VTAIL.n137 104.615
R152 VTAIL.n137 VTAIL.n111 104.615
R153 VTAIL.n130 VTAIL.n111 104.615
R154 VTAIL.n130 VTAIL.n129 104.615
R155 VTAIL.n129 VTAIL.n115 104.615
R156 VTAIL.n122 VTAIL.n115 104.615
R157 VTAIL.n122 VTAIL.n121 104.615
R158 VTAIL.n265 VTAIL.t6 52.3082
R159 VTAIL.n13 VTAIL.t7 52.3082
R160 VTAIL.n49 VTAIL.t2 52.3082
R161 VTAIL.n85 VTAIL.t5 52.3082
R162 VTAIL.n229 VTAIL.t3 52.3082
R163 VTAIL.n193 VTAIL.t4 52.3082
R164 VTAIL.n157 VTAIL.t0 52.3082
R165 VTAIL.n121 VTAIL.t1 52.3082
R166 VTAIL.n287 VTAIL.n286 31.7975
R167 VTAIL.n35 VTAIL.n34 31.7975
R168 VTAIL.n71 VTAIL.n70 31.7975
R169 VTAIL.n107 VTAIL.n106 31.7975
R170 VTAIL.n251 VTAIL.n250 31.7975
R171 VTAIL.n215 VTAIL.n214 31.7975
R172 VTAIL.n179 VTAIL.n178 31.7975
R173 VTAIL.n143 VTAIL.n142 31.7975
R174 VTAIL.n287 VTAIL.n251 19.841
R175 VTAIL.n143 VTAIL.n107 19.841
R176 VTAIL.n264 VTAIL.n263 15.6676
R177 VTAIL.n12 VTAIL.n11 15.6676
R178 VTAIL.n48 VTAIL.n47 15.6676
R179 VTAIL.n84 VTAIL.n83 15.6676
R180 VTAIL.n228 VTAIL.n227 15.6676
R181 VTAIL.n192 VTAIL.n191 15.6676
R182 VTAIL.n156 VTAIL.n155 15.6676
R183 VTAIL.n120 VTAIL.n119 15.6676
R184 VTAIL.n267 VTAIL.n262 12.8005
R185 VTAIL.n15 VTAIL.n10 12.8005
R186 VTAIL.n51 VTAIL.n46 12.8005
R187 VTAIL.n87 VTAIL.n82 12.8005
R188 VTAIL.n231 VTAIL.n226 12.8005
R189 VTAIL.n195 VTAIL.n190 12.8005
R190 VTAIL.n159 VTAIL.n154 12.8005
R191 VTAIL.n123 VTAIL.n118 12.8005
R192 VTAIL.n268 VTAIL.n260 12.0247
R193 VTAIL.n16 VTAIL.n8 12.0247
R194 VTAIL.n52 VTAIL.n44 12.0247
R195 VTAIL.n88 VTAIL.n80 12.0247
R196 VTAIL.n232 VTAIL.n224 12.0247
R197 VTAIL.n196 VTAIL.n188 12.0247
R198 VTAIL.n160 VTAIL.n152 12.0247
R199 VTAIL.n124 VTAIL.n116 12.0247
R200 VTAIL.n272 VTAIL.n271 11.249
R201 VTAIL.n20 VTAIL.n19 11.249
R202 VTAIL.n56 VTAIL.n55 11.249
R203 VTAIL.n92 VTAIL.n91 11.249
R204 VTAIL.n236 VTAIL.n235 11.249
R205 VTAIL.n200 VTAIL.n199 11.249
R206 VTAIL.n164 VTAIL.n163 11.249
R207 VTAIL.n128 VTAIL.n127 11.249
R208 VTAIL.n275 VTAIL.n258 10.4732
R209 VTAIL.n23 VTAIL.n6 10.4732
R210 VTAIL.n59 VTAIL.n42 10.4732
R211 VTAIL.n95 VTAIL.n78 10.4732
R212 VTAIL.n239 VTAIL.n222 10.4732
R213 VTAIL.n203 VTAIL.n186 10.4732
R214 VTAIL.n167 VTAIL.n150 10.4732
R215 VTAIL.n131 VTAIL.n114 10.4732
R216 VTAIL.n276 VTAIL.n256 9.69747
R217 VTAIL.n24 VTAIL.n4 9.69747
R218 VTAIL.n60 VTAIL.n40 9.69747
R219 VTAIL.n96 VTAIL.n76 9.69747
R220 VTAIL.n240 VTAIL.n220 9.69747
R221 VTAIL.n204 VTAIL.n184 9.69747
R222 VTAIL.n168 VTAIL.n148 9.69747
R223 VTAIL.n132 VTAIL.n112 9.69747
R224 VTAIL.n286 VTAIL.n285 9.45567
R225 VTAIL.n34 VTAIL.n33 9.45567
R226 VTAIL.n70 VTAIL.n69 9.45567
R227 VTAIL.n106 VTAIL.n105 9.45567
R228 VTAIL.n250 VTAIL.n249 9.45567
R229 VTAIL.n214 VTAIL.n213 9.45567
R230 VTAIL.n178 VTAIL.n177 9.45567
R231 VTAIL.n142 VTAIL.n141 9.45567
R232 VTAIL.n254 VTAIL.n253 9.3005
R233 VTAIL.n279 VTAIL.n278 9.3005
R234 VTAIL.n277 VTAIL.n276 9.3005
R235 VTAIL.n258 VTAIL.n257 9.3005
R236 VTAIL.n271 VTAIL.n270 9.3005
R237 VTAIL.n269 VTAIL.n268 9.3005
R238 VTAIL.n262 VTAIL.n261 9.3005
R239 VTAIL.n285 VTAIL.n284 9.3005
R240 VTAIL.n2 VTAIL.n1 9.3005
R241 VTAIL.n27 VTAIL.n26 9.3005
R242 VTAIL.n25 VTAIL.n24 9.3005
R243 VTAIL.n6 VTAIL.n5 9.3005
R244 VTAIL.n19 VTAIL.n18 9.3005
R245 VTAIL.n17 VTAIL.n16 9.3005
R246 VTAIL.n10 VTAIL.n9 9.3005
R247 VTAIL.n33 VTAIL.n32 9.3005
R248 VTAIL.n38 VTAIL.n37 9.3005
R249 VTAIL.n63 VTAIL.n62 9.3005
R250 VTAIL.n61 VTAIL.n60 9.3005
R251 VTAIL.n42 VTAIL.n41 9.3005
R252 VTAIL.n55 VTAIL.n54 9.3005
R253 VTAIL.n53 VTAIL.n52 9.3005
R254 VTAIL.n46 VTAIL.n45 9.3005
R255 VTAIL.n69 VTAIL.n68 9.3005
R256 VTAIL.n74 VTAIL.n73 9.3005
R257 VTAIL.n99 VTAIL.n98 9.3005
R258 VTAIL.n97 VTAIL.n96 9.3005
R259 VTAIL.n78 VTAIL.n77 9.3005
R260 VTAIL.n91 VTAIL.n90 9.3005
R261 VTAIL.n89 VTAIL.n88 9.3005
R262 VTAIL.n82 VTAIL.n81 9.3005
R263 VTAIL.n105 VTAIL.n104 9.3005
R264 VTAIL.n249 VTAIL.n248 9.3005
R265 VTAIL.n218 VTAIL.n217 9.3005
R266 VTAIL.n243 VTAIL.n242 9.3005
R267 VTAIL.n241 VTAIL.n240 9.3005
R268 VTAIL.n222 VTAIL.n221 9.3005
R269 VTAIL.n235 VTAIL.n234 9.3005
R270 VTAIL.n233 VTAIL.n232 9.3005
R271 VTAIL.n226 VTAIL.n225 9.3005
R272 VTAIL.n213 VTAIL.n212 9.3005
R273 VTAIL.n182 VTAIL.n181 9.3005
R274 VTAIL.n207 VTAIL.n206 9.3005
R275 VTAIL.n205 VTAIL.n204 9.3005
R276 VTAIL.n186 VTAIL.n185 9.3005
R277 VTAIL.n199 VTAIL.n198 9.3005
R278 VTAIL.n197 VTAIL.n196 9.3005
R279 VTAIL.n190 VTAIL.n189 9.3005
R280 VTAIL.n177 VTAIL.n176 9.3005
R281 VTAIL.n146 VTAIL.n145 9.3005
R282 VTAIL.n171 VTAIL.n170 9.3005
R283 VTAIL.n169 VTAIL.n168 9.3005
R284 VTAIL.n150 VTAIL.n149 9.3005
R285 VTAIL.n163 VTAIL.n162 9.3005
R286 VTAIL.n161 VTAIL.n160 9.3005
R287 VTAIL.n154 VTAIL.n153 9.3005
R288 VTAIL.n141 VTAIL.n140 9.3005
R289 VTAIL.n110 VTAIL.n109 9.3005
R290 VTAIL.n135 VTAIL.n134 9.3005
R291 VTAIL.n133 VTAIL.n132 9.3005
R292 VTAIL.n114 VTAIL.n113 9.3005
R293 VTAIL.n127 VTAIL.n126 9.3005
R294 VTAIL.n125 VTAIL.n124 9.3005
R295 VTAIL.n118 VTAIL.n117 9.3005
R296 VTAIL.n280 VTAIL.n279 8.92171
R297 VTAIL.n28 VTAIL.n27 8.92171
R298 VTAIL.n64 VTAIL.n63 8.92171
R299 VTAIL.n100 VTAIL.n99 8.92171
R300 VTAIL.n244 VTAIL.n243 8.92171
R301 VTAIL.n208 VTAIL.n207 8.92171
R302 VTAIL.n172 VTAIL.n171 8.92171
R303 VTAIL.n136 VTAIL.n135 8.92171
R304 VTAIL.n283 VTAIL.n254 8.14595
R305 VTAIL.n31 VTAIL.n2 8.14595
R306 VTAIL.n67 VTAIL.n38 8.14595
R307 VTAIL.n103 VTAIL.n74 8.14595
R308 VTAIL.n247 VTAIL.n218 8.14595
R309 VTAIL.n211 VTAIL.n182 8.14595
R310 VTAIL.n175 VTAIL.n146 8.14595
R311 VTAIL.n139 VTAIL.n110 8.14595
R312 VTAIL.n284 VTAIL.n252 7.3702
R313 VTAIL.n32 VTAIL.n0 7.3702
R314 VTAIL.n68 VTAIL.n36 7.3702
R315 VTAIL.n104 VTAIL.n72 7.3702
R316 VTAIL.n248 VTAIL.n216 7.3702
R317 VTAIL.n212 VTAIL.n180 7.3702
R318 VTAIL.n176 VTAIL.n144 7.3702
R319 VTAIL.n140 VTAIL.n108 7.3702
R320 VTAIL.n286 VTAIL.n252 6.59444
R321 VTAIL.n34 VTAIL.n0 6.59444
R322 VTAIL.n70 VTAIL.n36 6.59444
R323 VTAIL.n106 VTAIL.n72 6.59444
R324 VTAIL.n250 VTAIL.n216 6.59444
R325 VTAIL.n214 VTAIL.n180 6.59444
R326 VTAIL.n178 VTAIL.n144 6.59444
R327 VTAIL.n142 VTAIL.n108 6.59444
R328 VTAIL.n284 VTAIL.n283 5.81868
R329 VTAIL.n32 VTAIL.n31 5.81868
R330 VTAIL.n68 VTAIL.n67 5.81868
R331 VTAIL.n104 VTAIL.n103 5.81868
R332 VTAIL.n248 VTAIL.n247 5.81868
R333 VTAIL.n212 VTAIL.n211 5.81868
R334 VTAIL.n176 VTAIL.n175 5.81868
R335 VTAIL.n140 VTAIL.n139 5.81868
R336 VTAIL.n280 VTAIL.n254 5.04292
R337 VTAIL.n28 VTAIL.n2 5.04292
R338 VTAIL.n64 VTAIL.n38 5.04292
R339 VTAIL.n100 VTAIL.n74 5.04292
R340 VTAIL.n244 VTAIL.n218 5.04292
R341 VTAIL.n208 VTAIL.n182 5.04292
R342 VTAIL.n172 VTAIL.n146 5.04292
R343 VTAIL.n136 VTAIL.n110 5.04292
R344 VTAIL.n263 VTAIL.n261 4.38571
R345 VTAIL.n11 VTAIL.n9 4.38571
R346 VTAIL.n47 VTAIL.n45 4.38571
R347 VTAIL.n83 VTAIL.n81 4.38571
R348 VTAIL.n227 VTAIL.n225 4.38571
R349 VTAIL.n191 VTAIL.n189 4.38571
R350 VTAIL.n155 VTAIL.n153 4.38571
R351 VTAIL.n119 VTAIL.n117 4.38571
R352 VTAIL.n279 VTAIL.n256 4.26717
R353 VTAIL.n27 VTAIL.n4 4.26717
R354 VTAIL.n63 VTAIL.n40 4.26717
R355 VTAIL.n99 VTAIL.n76 4.26717
R356 VTAIL.n243 VTAIL.n220 4.26717
R357 VTAIL.n207 VTAIL.n184 4.26717
R358 VTAIL.n171 VTAIL.n148 4.26717
R359 VTAIL.n135 VTAIL.n112 4.26717
R360 VTAIL.n276 VTAIL.n275 3.49141
R361 VTAIL.n24 VTAIL.n23 3.49141
R362 VTAIL.n60 VTAIL.n59 3.49141
R363 VTAIL.n96 VTAIL.n95 3.49141
R364 VTAIL.n240 VTAIL.n239 3.49141
R365 VTAIL.n204 VTAIL.n203 3.49141
R366 VTAIL.n168 VTAIL.n167 3.49141
R367 VTAIL.n132 VTAIL.n131 3.49141
R368 VTAIL.n272 VTAIL.n258 2.71565
R369 VTAIL.n20 VTAIL.n6 2.71565
R370 VTAIL.n56 VTAIL.n42 2.71565
R371 VTAIL.n92 VTAIL.n78 2.71565
R372 VTAIL.n236 VTAIL.n222 2.71565
R373 VTAIL.n200 VTAIL.n186 2.71565
R374 VTAIL.n164 VTAIL.n150 2.71565
R375 VTAIL.n128 VTAIL.n114 2.71565
R376 VTAIL.n271 VTAIL.n260 1.93989
R377 VTAIL.n19 VTAIL.n8 1.93989
R378 VTAIL.n55 VTAIL.n44 1.93989
R379 VTAIL.n91 VTAIL.n80 1.93989
R380 VTAIL.n235 VTAIL.n224 1.93989
R381 VTAIL.n199 VTAIL.n188 1.93989
R382 VTAIL.n163 VTAIL.n152 1.93989
R383 VTAIL.n127 VTAIL.n116 1.93989
R384 VTAIL.n179 VTAIL.n143 1.69878
R385 VTAIL.n251 VTAIL.n215 1.69878
R386 VTAIL.n107 VTAIL.n71 1.69878
R387 VTAIL.n268 VTAIL.n267 1.16414
R388 VTAIL.n16 VTAIL.n15 1.16414
R389 VTAIL.n52 VTAIL.n51 1.16414
R390 VTAIL.n88 VTAIL.n87 1.16414
R391 VTAIL.n232 VTAIL.n231 1.16414
R392 VTAIL.n196 VTAIL.n195 1.16414
R393 VTAIL.n160 VTAIL.n159 1.16414
R394 VTAIL.n124 VTAIL.n123 1.16414
R395 VTAIL VTAIL.n35 0.907828
R396 VTAIL VTAIL.n287 0.791448
R397 VTAIL.n215 VTAIL.n179 0.470328
R398 VTAIL.n71 VTAIL.n35 0.470328
R399 VTAIL.n264 VTAIL.n262 0.388379
R400 VTAIL.n12 VTAIL.n10 0.388379
R401 VTAIL.n48 VTAIL.n46 0.388379
R402 VTAIL.n84 VTAIL.n82 0.388379
R403 VTAIL.n228 VTAIL.n226 0.388379
R404 VTAIL.n192 VTAIL.n190 0.388379
R405 VTAIL.n156 VTAIL.n154 0.388379
R406 VTAIL.n120 VTAIL.n118 0.388379
R407 VTAIL.n269 VTAIL.n261 0.155672
R408 VTAIL.n270 VTAIL.n269 0.155672
R409 VTAIL.n270 VTAIL.n257 0.155672
R410 VTAIL.n277 VTAIL.n257 0.155672
R411 VTAIL.n278 VTAIL.n277 0.155672
R412 VTAIL.n278 VTAIL.n253 0.155672
R413 VTAIL.n285 VTAIL.n253 0.155672
R414 VTAIL.n17 VTAIL.n9 0.155672
R415 VTAIL.n18 VTAIL.n17 0.155672
R416 VTAIL.n18 VTAIL.n5 0.155672
R417 VTAIL.n25 VTAIL.n5 0.155672
R418 VTAIL.n26 VTAIL.n25 0.155672
R419 VTAIL.n26 VTAIL.n1 0.155672
R420 VTAIL.n33 VTAIL.n1 0.155672
R421 VTAIL.n53 VTAIL.n45 0.155672
R422 VTAIL.n54 VTAIL.n53 0.155672
R423 VTAIL.n54 VTAIL.n41 0.155672
R424 VTAIL.n61 VTAIL.n41 0.155672
R425 VTAIL.n62 VTAIL.n61 0.155672
R426 VTAIL.n62 VTAIL.n37 0.155672
R427 VTAIL.n69 VTAIL.n37 0.155672
R428 VTAIL.n89 VTAIL.n81 0.155672
R429 VTAIL.n90 VTAIL.n89 0.155672
R430 VTAIL.n90 VTAIL.n77 0.155672
R431 VTAIL.n97 VTAIL.n77 0.155672
R432 VTAIL.n98 VTAIL.n97 0.155672
R433 VTAIL.n98 VTAIL.n73 0.155672
R434 VTAIL.n105 VTAIL.n73 0.155672
R435 VTAIL.n249 VTAIL.n217 0.155672
R436 VTAIL.n242 VTAIL.n217 0.155672
R437 VTAIL.n242 VTAIL.n241 0.155672
R438 VTAIL.n241 VTAIL.n221 0.155672
R439 VTAIL.n234 VTAIL.n221 0.155672
R440 VTAIL.n234 VTAIL.n233 0.155672
R441 VTAIL.n233 VTAIL.n225 0.155672
R442 VTAIL.n213 VTAIL.n181 0.155672
R443 VTAIL.n206 VTAIL.n181 0.155672
R444 VTAIL.n206 VTAIL.n205 0.155672
R445 VTAIL.n205 VTAIL.n185 0.155672
R446 VTAIL.n198 VTAIL.n185 0.155672
R447 VTAIL.n198 VTAIL.n197 0.155672
R448 VTAIL.n197 VTAIL.n189 0.155672
R449 VTAIL.n177 VTAIL.n145 0.155672
R450 VTAIL.n170 VTAIL.n145 0.155672
R451 VTAIL.n170 VTAIL.n169 0.155672
R452 VTAIL.n169 VTAIL.n149 0.155672
R453 VTAIL.n162 VTAIL.n149 0.155672
R454 VTAIL.n162 VTAIL.n161 0.155672
R455 VTAIL.n161 VTAIL.n153 0.155672
R456 VTAIL.n141 VTAIL.n109 0.155672
R457 VTAIL.n134 VTAIL.n109 0.155672
R458 VTAIL.n134 VTAIL.n133 0.155672
R459 VTAIL.n133 VTAIL.n113 0.155672
R460 VTAIL.n126 VTAIL.n113 0.155672
R461 VTAIL.n126 VTAIL.n125 0.155672
R462 VTAIL.n125 VTAIL.n117 0.155672
R463 VDD1 VDD1.n1 100.796
R464 VDD1 VDD1.n0 65.7443
R465 VDD1.n0 VDD1.t1 2.95572
R466 VDD1.n0 VDD1.t3 2.95572
R467 VDD1.n1 VDD1.t2 2.95572
R468 VDD1.n1 VDD1.t0 2.95572
R469 B.n525 B.n524 585
R470 B.n207 B.n80 585
R471 B.n206 B.n205 585
R472 B.n204 B.n203 585
R473 B.n202 B.n201 585
R474 B.n200 B.n199 585
R475 B.n198 B.n197 585
R476 B.n196 B.n195 585
R477 B.n194 B.n193 585
R478 B.n192 B.n191 585
R479 B.n190 B.n189 585
R480 B.n188 B.n187 585
R481 B.n186 B.n185 585
R482 B.n184 B.n183 585
R483 B.n182 B.n181 585
R484 B.n180 B.n179 585
R485 B.n178 B.n177 585
R486 B.n176 B.n175 585
R487 B.n174 B.n173 585
R488 B.n172 B.n171 585
R489 B.n170 B.n169 585
R490 B.n168 B.n167 585
R491 B.n166 B.n165 585
R492 B.n164 B.n163 585
R493 B.n162 B.n161 585
R494 B.n160 B.n159 585
R495 B.n158 B.n157 585
R496 B.n156 B.n155 585
R497 B.n154 B.n153 585
R498 B.n152 B.n151 585
R499 B.n150 B.n149 585
R500 B.n148 B.n147 585
R501 B.n146 B.n145 585
R502 B.n144 B.n143 585
R503 B.n142 B.n141 585
R504 B.n140 B.n139 585
R505 B.n138 B.n137 585
R506 B.n136 B.n135 585
R507 B.n134 B.n133 585
R508 B.n132 B.n131 585
R509 B.n130 B.n129 585
R510 B.n128 B.n127 585
R511 B.n126 B.n125 585
R512 B.n124 B.n123 585
R513 B.n122 B.n121 585
R514 B.n120 B.n119 585
R515 B.n118 B.n117 585
R516 B.n116 B.n115 585
R517 B.n114 B.n113 585
R518 B.n112 B.n111 585
R519 B.n110 B.n109 585
R520 B.n108 B.n107 585
R521 B.n106 B.n105 585
R522 B.n104 B.n103 585
R523 B.n102 B.n101 585
R524 B.n100 B.n99 585
R525 B.n98 B.n97 585
R526 B.n96 B.n95 585
R527 B.n94 B.n93 585
R528 B.n92 B.n91 585
R529 B.n90 B.n89 585
R530 B.n88 B.n87 585
R531 B.n523 B.n49 585
R532 B.n528 B.n49 585
R533 B.n522 B.n48 585
R534 B.n529 B.n48 585
R535 B.n521 B.n520 585
R536 B.n520 B.n44 585
R537 B.n519 B.n43 585
R538 B.n535 B.n43 585
R539 B.n518 B.n42 585
R540 B.n536 B.n42 585
R541 B.n517 B.n41 585
R542 B.n537 B.n41 585
R543 B.n516 B.n515 585
R544 B.n515 B.n40 585
R545 B.n514 B.n36 585
R546 B.n543 B.n36 585
R547 B.n513 B.n35 585
R548 B.n544 B.n35 585
R549 B.n512 B.n34 585
R550 B.n545 B.n34 585
R551 B.n511 B.n510 585
R552 B.n510 B.n30 585
R553 B.n509 B.n29 585
R554 B.n551 B.n29 585
R555 B.n508 B.n28 585
R556 B.n552 B.n28 585
R557 B.n507 B.n27 585
R558 B.n553 B.n27 585
R559 B.n506 B.n505 585
R560 B.n505 B.n23 585
R561 B.n504 B.n22 585
R562 B.n559 B.n22 585
R563 B.n503 B.n21 585
R564 B.n560 B.n21 585
R565 B.n502 B.n20 585
R566 B.n561 B.n20 585
R567 B.n501 B.n500 585
R568 B.n500 B.n16 585
R569 B.n499 B.n15 585
R570 B.n567 B.n15 585
R571 B.n498 B.n14 585
R572 B.n568 B.n14 585
R573 B.n497 B.n13 585
R574 B.t2 B.n13 585
R575 B.n496 B.n495 585
R576 B.n495 B.n12 585
R577 B.n494 B.n493 585
R578 B.n494 B.n8 585
R579 B.n492 B.n7 585
R580 B.n575 B.n7 585
R581 B.n491 B.n6 585
R582 B.n576 B.n6 585
R583 B.n490 B.n5 585
R584 B.n577 B.n5 585
R585 B.n489 B.n488 585
R586 B.n488 B.n4 585
R587 B.n487 B.n208 585
R588 B.n487 B.n486 585
R589 B.n478 B.n209 585
R590 B.n210 B.n209 585
R591 B.n480 B.n479 585
R592 B.t0 B.n480 585
R593 B.n477 B.n215 585
R594 B.n215 B.n214 585
R595 B.n476 B.n475 585
R596 B.n475 B.n474 585
R597 B.n217 B.n216 585
R598 B.n218 B.n217 585
R599 B.n467 B.n466 585
R600 B.n468 B.n467 585
R601 B.n465 B.n223 585
R602 B.n223 B.n222 585
R603 B.n464 B.n463 585
R604 B.n463 B.n462 585
R605 B.n225 B.n224 585
R606 B.n226 B.n225 585
R607 B.n455 B.n454 585
R608 B.n456 B.n455 585
R609 B.n453 B.n231 585
R610 B.n231 B.n230 585
R611 B.n452 B.n451 585
R612 B.n451 B.n450 585
R613 B.n233 B.n232 585
R614 B.n234 B.n233 585
R615 B.n443 B.n442 585
R616 B.n444 B.n443 585
R617 B.n441 B.n239 585
R618 B.n239 B.n238 585
R619 B.n440 B.n439 585
R620 B.n439 B.n438 585
R621 B.n241 B.n240 585
R622 B.n431 B.n241 585
R623 B.n430 B.n429 585
R624 B.n432 B.n430 585
R625 B.n428 B.n246 585
R626 B.n246 B.n245 585
R627 B.n427 B.n426 585
R628 B.n426 B.n425 585
R629 B.n248 B.n247 585
R630 B.n249 B.n248 585
R631 B.n418 B.n417 585
R632 B.n419 B.n418 585
R633 B.n416 B.n254 585
R634 B.n254 B.n253 585
R635 B.n411 B.n410 585
R636 B.n409 B.n287 585
R637 B.n408 B.n286 585
R638 B.n413 B.n286 585
R639 B.n407 B.n406 585
R640 B.n405 B.n404 585
R641 B.n403 B.n402 585
R642 B.n401 B.n400 585
R643 B.n399 B.n398 585
R644 B.n397 B.n396 585
R645 B.n395 B.n394 585
R646 B.n393 B.n392 585
R647 B.n391 B.n390 585
R648 B.n389 B.n388 585
R649 B.n387 B.n386 585
R650 B.n385 B.n384 585
R651 B.n383 B.n382 585
R652 B.n381 B.n380 585
R653 B.n379 B.n378 585
R654 B.n377 B.n376 585
R655 B.n375 B.n374 585
R656 B.n373 B.n372 585
R657 B.n371 B.n370 585
R658 B.n369 B.n368 585
R659 B.n367 B.n366 585
R660 B.n365 B.n364 585
R661 B.n363 B.n362 585
R662 B.n360 B.n359 585
R663 B.n358 B.n357 585
R664 B.n356 B.n355 585
R665 B.n354 B.n353 585
R666 B.n352 B.n351 585
R667 B.n350 B.n349 585
R668 B.n348 B.n347 585
R669 B.n346 B.n345 585
R670 B.n344 B.n343 585
R671 B.n342 B.n341 585
R672 B.n339 B.n338 585
R673 B.n337 B.n336 585
R674 B.n335 B.n334 585
R675 B.n333 B.n332 585
R676 B.n331 B.n330 585
R677 B.n329 B.n328 585
R678 B.n327 B.n326 585
R679 B.n325 B.n324 585
R680 B.n323 B.n322 585
R681 B.n321 B.n320 585
R682 B.n319 B.n318 585
R683 B.n317 B.n316 585
R684 B.n315 B.n314 585
R685 B.n313 B.n312 585
R686 B.n311 B.n310 585
R687 B.n309 B.n308 585
R688 B.n307 B.n306 585
R689 B.n305 B.n304 585
R690 B.n303 B.n302 585
R691 B.n301 B.n300 585
R692 B.n299 B.n298 585
R693 B.n297 B.n296 585
R694 B.n295 B.n294 585
R695 B.n293 B.n292 585
R696 B.n256 B.n255 585
R697 B.n415 B.n414 585
R698 B.n414 B.n413 585
R699 B.n252 B.n251 585
R700 B.n253 B.n252 585
R701 B.n421 B.n420 585
R702 B.n420 B.n419 585
R703 B.n422 B.n250 585
R704 B.n250 B.n249 585
R705 B.n424 B.n423 585
R706 B.n425 B.n424 585
R707 B.n244 B.n243 585
R708 B.n245 B.n244 585
R709 B.n434 B.n433 585
R710 B.n433 B.n432 585
R711 B.n435 B.n242 585
R712 B.n431 B.n242 585
R713 B.n437 B.n436 585
R714 B.n438 B.n437 585
R715 B.n237 B.n236 585
R716 B.n238 B.n237 585
R717 B.n446 B.n445 585
R718 B.n445 B.n444 585
R719 B.n447 B.n235 585
R720 B.n235 B.n234 585
R721 B.n449 B.n448 585
R722 B.n450 B.n449 585
R723 B.n229 B.n228 585
R724 B.n230 B.n229 585
R725 B.n458 B.n457 585
R726 B.n457 B.n456 585
R727 B.n459 B.n227 585
R728 B.n227 B.n226 585
R729 B.n461 B.n460 585
R730 B.n462 B.n461 585
R731 B.n221 B.n220 585
R732 B.n222 B.n221 585
R733 B.n470 B.n469 585
R734 B.n469 B.n468 585
R735 B.n471 B.n219 585
R736 B.n219 B.n218 585
R737 B.n473 B.n472 585
R738 B.n474 B.n473 585
R739 B.n213 B.n212 585
R740 B.n214 B.n213 585
R741 B.n482 B.n481 585
R742 B.n481 B.t0 585
R743 B.n483 B.n211 585
R744 B.n211 B.n210 585
R745 B.n485 B.n484 585
R746 B.n486 B.n485 585
R747 B.n3 B.n0 585
R748 B.n4 B.n3 585
R749 B.n574 B.n1 585
R750 B.n575 B.n574 585
R751 B.n573 B.n572 585
R752 B.n573 B.n8 585
R753 B.n571 B.n9 585
R754 B.n12 B.n9 585
R755 B.n570 B.n569 585
R756 B.n569 B.t2 585
R757 B.n11 B.n10 585
R758 B.n568 B.n11 585
R759 B.n566 B.n565 585
R760 B.n567 B.n566 585
R761 B.n564 B.n17 585
R762 B.n17 B.n16 585
R763 B.n563 B.n562 585
R764 B.n562 B.n561 585
R765 B.n19 B.n18 585
R766 B.n560 B.n19 585
R767 B.n558 B.n557 585
R768 B.n559 B.n558 585
R769 B.n556 B.n24 585
R770 B.n24 B.n23 585
R771 B.n555 B.n554 585
R772 B.n554 B.n553 585
R773 B.n26 B.n25 585
R774 B.n552 B.n26 585
R775 B.n550 B.n549 585
R776 B.n551 B.n550 585
R777 B.n548 B.n31 585
R778 B.n31 B.n30 585
R779 B.n547 B.n546 585
R780 B.n546 B.n545 585
R781 B.n33 B.n32 585
R782 B.n544 B.n33 585
R783 B.n542 B.n541 585
R784 B.n543 B.n542 585
R785 B.n540 B.n37 585
R786 B.n40 B.n37 585
R787 B.n539 B.n538 585
R788 B.n538 B.n537 585
R789 B.n39 B.n38 585
R790 B.n536 B.n39 585
R791 B.n534 B.n533 585
R792 B.n535 B.n534 585
R793 B.n532 B.n45 585
R794 B.n45 B.n44 585
R795 B.n531 B.n530 585
R796 B.n530 B.n529 585
R797 B.n47 B.n46 585
R798 B.n528 B.n47 585
R799 B.n578 B.n577 585
R800 B.n576 B.n2 585
R801 B.n87 B.n47 468.476
R802 B.n525 B.n49 468.476
R803 B.n414 B.n254 468.476
R804 B.n411 B.n252 468.476
R805 B.n84 B.t15 304.384
R806 B.n81 B.t4 304.384
R807 B.n290 B.t8 304.384
R808 B.n288 B.t12 304.384
R809 B.n527 B.n526 256.663
R810 B.n527 B.n79 256.663
R811 B.n527 B.n78 256.663
R812 B.n527 B.n77 256.663
R813 B.n527 B.n76 256.663
R814 B.n527 B.n75 256.663
R815 B.n527 B.n74 256.663
R816 B.n527 B.n73 256.663
R817 B.n527 B.n72 256.663
R818 B.n527 B.n71 256.663
R819 B.n527 B.n70 256.663
R820 B.n527 B.n69 256.663
R821 B.n527 B.n68 256.663
R822 B.n527 B.n67 256.663
R823 B.n527 B.n66 256.663
R824 B.n527 B.n65 256.663
R825 B.n527 B.n64 256.663
R826 B.n527 B.n63 256.663
R827 B.n527 B.n62 256.663
R828 B.n527 B.n61 256.663
R829 B.n527 B.n60 256.663
R830 B.n527 B.n59 256.663
R831 B.n527 B.n58 256.663
R832 B.n527 B.n57 256.663
R833 B.n527 B.n56 256.663
R834 B.n527 B.n55 256.663
R835 B.n527 B.n54 256.663
R836 B.n527 B.n53 256.663
R837 B.n527 B.n52 256.663
R838 B.n527 B.n51 256.663
R839 B.n527 B.n50 256.663
R840 B.n413 B.n412 256.663
R841 B.n413 B.n257 256.663
R842 B.n413 B.n258 256.663
R843 B.n413 B.n259 256.663
R844 B.n413 B.n260 256.663
R845 B.n413 B.n261 256.663
R846 B.n413 B.n262 256.663
R847 B.n413 B.n263 256.663
R848 B.n413 B.n264 256.663
R849 B.n413 B.n265 256.663
R850 B.n413 B.n266 256.663
R851 B.n413 B.n267 256.663
R852 B.n413 B.n268 256.663
R853 B.n413 B.n269 256.663
R854 B.n413 B.n270 256.663
R855 B.n413 B.n271 256.663
R856 B.n413 B.n272 256.663
R857 B.n413 B.n273 256.663
R858 B.n413 B.n274 256.663
R859 B.n413 B.n275 256.663
R860 B.n413 B.n276 256.663
R861 B.n413 B.n277 256.663
R862 B.n413 B.n278 256.663
R863 B.n413 B.n279 256.663
R864 B.n413 B.n280 256.663
R865 B.n413 B.n281 256.663
R866 B.n413 B.n282 256.663
R867 B.n413 B.n283 256.663
R868 B.n413 B.n284 256.663
R869 B.n413 B.n285 256.663
R870 B.n580 B.n579 256.663
R871 B.n81 B.t6 229.258
R872 B.n290 B.t11 229.258
R873 B.n84 B.t16 229.258
R874 B.n288 B.t14 229.258
R875 B.n82 B.t7 191.053
R876 B.n291 B.t10 191.053
R877 B.n85 B.t17 191.053
R878 B.n289 B.t13 191.053
R879 B.n91 B.n90 163.367
R880 B.n95 B.n94 163.367
R881 B.n99 B.n98 163.367
R882 B.n103 B.n102 163.367
R883 B.n107 B.n106 163.367
R884 B.n111 B.n110 163.367
R885 B.n115 B.n114 163.367
R886 B.n119 B.n118 163.367
R887 B.n123 B.n122 163.367
R888 B.n127 B.n126 163.367
R889 B.n131 B.n130 163.367
R890 B.n135 B.n134 163.367
R891 B.n139 B.n138 163.367
R892 B.n143 B.n142 163.367
R893 B.n147 B.n146 163.367
R894 B.n151 B.n150 163.367
R895 B.n155 B.n154 163.367
R896 B.n159 B.n158 163.367
R897 B.n163 B.n162 163.367
R898 B.n167 B.n166 163.367
R899 B.n171 B.n170 163.367
R900 B.n175 B.n174 163.367
R901 B.n179 B.n178 163.367
R902 B.n183 B.n182 163.367
R903 B.n187 B.n186 163.367
R904 B.n191 B.n190 163.367
R905 B.n195 B.n194 163.367
R906 B.n199 B.n198 163.367
R907 B.n203 B.n202 163.367
R908 B.n205 B.n80 163.367
R909 B.n418 B.n254 163.367
R910 B.n418 B.n248 163.367
R911 B.n426 B.n248 163.367
R912 B.n426 B.n246 163.367
R913 B.n430 B.n246 163.367
R914 B.n430 B.n241 163.367
R915 B.n439 B.n241 163.367
R916 B.n439 B.n239 163.367
R917 B.n443 B.n239 163.367
R918 B.n443 B.n233 163.367
R919 B.n451 B.n233 163.367
R920 B.n451 B.n231 163.367
R921 B.n455 B.n231 163.367
R922 B.n455 B.n225 163.367
R923 B.n463 B.n225 163.367
R924 B.n463 B.n223 163.367
R925 B.n467 B.n223 163.367
R926 B.n467 B.n217 163.367
R927 B.n475 B.n217 163.367
R928 B.n475 B.n215 163.367
R929 B.n480 B.n215 163.367
R930 B.n480 B.n209 163.367
R931 B.n487 B.n209 163.367
R932 B.n488 B.n487 163.367
R933 B.n488 B.n5 163.367
R934 B.n6 B.n5 163.367
R935 B.n7 B.n6 163.367
R936 B.n494 B.n7 163.367
R937 B.n495 B.n494 163.367
R938 B.n495 B.n13 163.367
R939 B.n14 B.n13 163.367
R940 B.n15 B.n14 163.367
R941 B.n500 B.n15 163.367
R942 B.n500 B.n20 163.367
R943 B.n21 B.n20 163.367
R944 B.n22 B.n21 163.367
R945 B.n505 B.n22 163.367
R946 B.n505 B.n27 163.367
R947 B.n28 B.n27 163.367
R948 B.n29 B.n28 163.367
R949 B.n510 B.n29 163.367
R950 B.n510 B.n34 163.367
R951 B.n35 B.n34 163.367
R952 B.n36 B.n35 163.367
R953 B.n515 B.n36 163.367
R954 B.n515 B.n41 163.367
R955 B.n42 B.n41 163.367
R956 B.n43 B.n42 163.367
R957 B.n520 B.n43 163.367
R958 B.n520 B.n48 163.367
R959 B.n49 B.n48 163.367
R960 B.n287 B.n286 163.367
R961 B.n406 B.n286 163.367
R962 B.n404 B.n403 163.367
R963 B.n400 B.n399 163.367
R964 B.n396 B.n395 163.367
R965 B.n392 B.n391 163.367
R966 B.n388 B.n387 163.367
R967 B.n384 B.n383 163.367
R968 B.n380 B.n379 163.367
R969 B.n376 B.n375 163.367
R970 B.n372 B.n371 163.367
R971 B.n368 B.n367 163.367
R972 B.n364 B.n363 163.367
R973 B.n359 B.n358 163.367
R974 B.n355 B.n354 163.367
R975 B.n351 B.n350 163.367
R976 B.n347 B.n346 163.367
R977 B.n343 B.n342 163.367
R978 B.n338 B.n337 163.367
R979 B.n334 B.n333 163.367
R980 B.n330 B.n329 163.367
R981 B.n326 B.n325 163.367
R982 B.n322 B.n321 163.367
R983 B.n318 B.n317 163.367
R984 B.n314 B.n313 163.367
R985 B.n310 B.n309 163.367
R986 B.n306 B.n305 163.367
R987 B.n302 B.n301 163.367
R988 B.n298 B.n297 163.367
R989 B.n294 B.n293 163.367
R990 B.n414 B.n256 163.367
R991 B.n420 B.n252 163.367
R992 B.n420 B.n250 163.367
R993 B.n424 B.n250 163.367
R994 B.n424 B.n244 163.367
R995 B.n433 B.n244 163.367
R996 B.n433 B.n242 163.367
R997 B.n437 B.n242 163.367
R998 B.n437 B.n237 163.367
R999 B.n445 B.n237 163.367
R1000 B.n445 B.n235 163.367
R1001 B.n449 B.n235 163.367
R1002 B.n449 B.n229 163.367
R1003 B.n457 B.n229 163.367
R1004 B.n457 B.n227 163.367
R1005 B.n461 B.n227 163.367
R1006 B.n461 B.n221 163.367
R1007 B.n469 B.n221 163.367
R1008 B.n469 B.n219 163.367
R1009 B.n473 B.n219 163.367
R1010 B.n473 B.n213 163.367
R1011 B.n481 B.n213 163.367
R1012 B.n481 B.n211 163.367
R1013 B.n485 B.n211 163.367
R1014 B.n485 B.n3 163.367
R1015 B.n578 B.n3 163.367
R1016 B.n574 B.n2 163.367
R1017 B.n574 B.n573 163.367
R1018 B.n573 B.n9 163.367
R1019 B.n569 B.n9 163.367
R1020 B.n569 B.n11 163.367
R1021 B.n566 B.n11 163.367
R1022 B.n566 B.n17 163.367
R1023 B.n562 B.n17 163.367
R1024 B.n562 B.n19 163.367
R1025 B.n558 B.n19 163.367
R1026 B.n558 B.n24 163.367
R1027 B.n554 B.n24 163.367
R1028 B.n554 B.n26 163.367
R1029 B.n550 B.n26 163.367
R1030 B.n550 B.n31 163.367
R1031 B.n546 B.n31 163.367
R1032 B.n546 B.n33 163.367
R1033 B.n542 B.n33 163.367
R1034 B.n542 B.n37 163.367
R1035 B.n538 B.n37 163.367
R1036 B.n538 B.n39 163.367
R1037 B.n534 B.n39 163.367
R1038 B.n534 B.n45 163.367
R1039 B.n530 B.n45 163.367
R1040 B.n530 B.n47 163.367
R1041 B.n413 B.n253 112.986
R1042 B.n528 B.n527 112.986
R1043 B.n87 B.n50 71.676
R1044 B.n91 B.n51 71.676
R1045 B.n95 B.n52 71.676
R1046 B.n99 B.n53 71.676
R1047 B.n103 B.n54 71.676
R1048 B.n107 B.n55 71.676
R1049 B.n111 B.n56 71.676
R1050 B.n115 B.n57 71.676
R1051 B.n119 B.n58 71.676
R1052 B.n123 B.n59 71.676
R1053 B.n127 B.n60 71.676
R1054 B.n131 B.n61 71.676
R1055 B.n135 B.n62 71.676
R1056 B.n139 B.n63 71.676
R1057 B.n143 B.n64 71.676
R1058 B.n147 B.n65 71.676
R1059 B.n151 B.n66 71.676
R1060 B.n155 B.n67 71.676
R1061 B.n159 B.n68 71.676
R1062 B.n163 B.n69 71.676
R1063 B.n167 B.n70 71.676
R1064 B.n171 B.n71 71.676
R1065 B.n175 B.n72 71.676
R1066 B.n179 B.n73 71.676
R1067 B.n183 B.n74 71.676
R1068 B.n187 B.n75 71.676
R1069 B.n191 B.n76 71.676
R1070 B.n195 B.n77 71.676
R1071 B.n199 B.n78 71.676
R1072 B.n203 B.n79 71.676
R1073 B.n526 B.n80 71.676
R1074 B.n526 B.n525 71.676
R1075 B.n205 B.n79 71.676
R1076 B.n202 B.n78 71.676
R1077 B.n198 B.n77 71.676
R1078 B.n194 B.n76 71.676
R1079 B.n190 B.n75 71.676
R1080 B.n186 B.n74 71.676
R1081 B.n182 B.n73 71.676
R1082 B.n178 B.n72 71.676
R1083 B.n174 B.n71 71.676
R1084 B.n170 B.n70 71.676
R1085 B.n166 B.n69 71.676
R1086 B.n162 B.n68 71.676
R1087 B.n158 B.n67 71.676
R1088 B.n154 B.n66 71.676
R1089 B.n150 B.n65 71.676
R1090 B.n146 B.n64 71.676
R1091 B.n142 B.n63 71.676
R1092 B.n138 B.n62 71.676
R1093 B.n134 B.n61 71.676
R1094 B.n130 B.n60 71.676
R1095 B.n126 B.n59 71.676
R1096 B.n122 B.n58 71.676
R1097 B.n118 B.n57 71.676
R1098 B.n114 B.n56 71.676
R1099 B.n110 B.n55 71.676
R1100 B.n106 B.n54 71.676
R1101 B.n102 B.n53 71.676
R1102 B.n98 B.n52 71.676
R1103 B.n94 B.n51 71.676
R1104 B.n90 B.n50 71.676
R1105 B.n412 B.n411 71.676
R1106 B.n406 B.n257 71.676
R1107 B.n403 B.n258 71.676
R1108 B.n399 B.n259 71.676
R1109 B.n395 B.n260 71.676
R1110 B.n391 B.n261 71.676
R1111 B.n387 B.n262 71.676
R1112 B.n383 B.n263 71.676
R1113 B.n379 B.n264 71.676
R1114 B.n375 B.n265 71.676
R1115 B.n371 B.n266 71.676
R1116 B.n367 B.n267 71.676
R1117 B.n363 B.n268 71.676
R1118 B.n358 B.n269 71.676
R1119 B.n354 B.n270 71.676
R1120 B.n350 B.n271 71.676
R1121 B.n346 B.n272 71.676
R1122 B.n342 B.n273 71.676
R1123 B.n337 B.n274 71.676
R1124 B.n333 B.n275 71.676
R1125 B.n329 B.n276 71.676
R1126 B.n325 B.n277 71.676
R1127 B.n321 B.n278 71.676
R1128 B.n317 B.n279 71.676
R1129 B.n313 B.n280 71.676
R1130 B.n309 B.n281 71.676
R1131 B.n305 B.n282 71.676
R1132 B.n301 B.n283 71.676
R1133 B.n297 B.n284 71.676
R1134 B.n293 B.n285 71.676
R1135 B.n412 B.n287 71.676
R1136 B.n404 B.n257 71.676
R1137 B.n400 B.n258 71.676
R1138 B.n396 B.n259 71.676
R1139 B.n392 B.n260 71.676
R1140 B.n388 B.n261 71.676
R1141 B.n384 B.n262 71.676
R1142 B.n380 B.n263 71.676
R1143 B.n376 B.n264 71.676
R1144 B.n372 B.n265 71.676
R1145 B.n368 B.n266 71.676
R1146 B.n364 B.n267 71.676
R1147 B.n359 B.n268 71.676
R1148 B.n355 B.n269 71.676
R1149 B.n351 B.n270 71.676
R1150 B.n347 B.n271 71.676
R1151 B.n343 B.n272 71.676
R1152 B.n338 B.n273 71.676
R1153 B.n334 B.n274 71.676
R1154 B.n330 B.n275 71.676
R1155 B.n326 B.n276 71.676
R1156 B.n322 B.n277 71.676
R1157 B.n318 B.n278 71.676
R1158 B.n314 B.n279 71.676
R1159 B.n310 B.n280 71.676
R1160 B.n306 B.n281 71.676
R1161 B.n302 B.n282 71.676
R1162 B.n298 B.n283 71.676
R1163 B.n294 B.n284 71.676
R1164 B.n285 B.n256 71.676
R1165 B.n579 B.n578 71.676
R1166 B.n579 B.n2 71.676
R1167 B.n419 B.n253 62.464
R1168 B.n419 B.n249 62.464
R1169 B.n425 B.n249 62.464
R1170 B.n425 B.n245 62.464
R1171 B.n432 B.n245 62.464
R1172 B.n432 B.n431 62.464
R1173 B.n438 B.n238 62.464
R1174 B.n444 B.n238 62.464
R1175 B.n444 B.n234 62.464
R1176 B.n450 B.n234 62.464
R1177 B.n450 B.n230 62.464
R1178 B.n456 B.n230 62.464
R1179 B.n456 B.n226 62.464
R1180 B.n462 B.n226 62.464
R1181 B.n468 B.n222 62.464
R1182 B.n468 B.n218 62.464
R1183 B.n474 B.n218 62.464
R1184 B.n474 B.n214 62.464
R1185 B.t0 B.n214 62.464
R1186 B.t0 B.n210 62.464
R1187 B.n486 B.n210 62.464
R1188 B.n486 B.n4 62.464
R1189 B.n577 B.n4 62.464
R1190 B.n577 B.n576 62.464
R1191 B.n576 B.n575 62.464
R1192 B.n575 B.n8 62.464
R1193 B.n12 B.n8 62.464
R1194 B.t2 B.n12 62.464
R1195 B.t2 B.n568 62.464
R1196 B.n568 B.n567 62.464
R1197 B.n567 B.n16 62.464
R1198 B.n561 B.n16 62.464
R1199 B.n561 B.n560 62.464
R1200 B.n559 B.n23 62.464
R1201 B.n553 B.n23 62.464
R1202 B.n553 B.n552 62.464
R1203 B.n552 B.n551 62.464
R1204 B.n551 B.n30 62.464
R1205 B.n545 B.n30 62.464
R1206 B.n545 B.n544 62.464
R1207 B.n544 B.n543 62.464
R1208 B.n537 B.n40 62.464
R1209 B.n537 B.n536 62.464
R1210 B.n536 B.n535 62.464
R1211 B.n535 B.n44 62.464
R1212 B.n529 B.n44 62.464
R1213 B.n529 B.n528 62.464
R1214 B.n86 B.n85 59.5399
R1215 B.n83 B.n82 59.5399
R1216 B.n340 B.n291 59.5399
R1217 B.n361 B.n289 59.5399
R1218 B.n438 B.t9 49.6038
R1219 B.t1 B.n222 49.6038
R1220 B.n560 B.t3 49.6038
R1221 B.n543 B.t5 49.6038
R1222 B.n85 B.n84 38.2066
R1223 B.n82 B.n81 38.2066
R1224 B.n291 B.n290 38.2066
R1225 B.n289 B.n288 38.2066
R1226 B.n410 B.n251 30.4395
R1227 B.n416 B.n415 30.4395
R1228 B.n524 B.n523 30.4395
R1229 B.n88 B.n46 30.4395
R1230 B B.n580 18.0485
R1231 B.n431 B.t9 12.8606
R1232 B.n462 B.t1 12.8606
R1233 B.t3 B.n559 12.8606
R1234 B.n40 B.t5 12.8606
R1235 B.n421 B.n251 10.6151
R1236 B.n422 B.n421 10.6151
R1237 B.n423 B.n422 10.6151
R1238 B.n423 B.n243 10.6151
R1239 B.n434 B.n243 10.6151
R1240 B.n435 B.n434 10.6151
R1241 B.n436 B.n435 10.6151
R1242 B.n436 B.n236 10.6151
R1243 B.n446 B.n236 10.6151
R1244 B.n447 B.n446 10.6151
R1245 B.n448 B.n447 10.6151
R1246 B.n448 B.n228 10.6151
R1247 B.n458 B.n228 10.6151
R1248 B.n459 B.n458 10.6151
R1249 B.n460 B.n459 10.6151
R1250 B.n460 B.n220 10.6151
R1251 B.n470 B.n220 10.6151
R1252 B.n471 B.n470 10.6151
R1253 B.n472 B.n471 10.6151
R1254 B.n472 B.n212 10.6151
R1255 B.n482 B.n212 10.6151
R1256 B.n483 B.n482 10.6151
R1257 B.n484 B.n483 10.6151
R1258 B.n484 B.n0 10.6151
R1259 B.n410 B.n409 10.6151
R1260 B.n409 B.n408 10.6151
R1261 B.n408 B.n407 10.6151
R1262 B.n407 B.n405 10.6151
R1263 B.n405 B.n402 10.6151
R1264 B.n402 B.n401 10.6151
R1265 B.n401 B.n398 10.6151
R1266 B.n398 B.n397 10.6151
R1267 B.n397 B.n394 10.6151
R1268 B.n394 B.n393 10.6151
R1269 B.n393 B.n390 10.6151
R1270 B.n390 B.n389 10.6151
R1271 B.n389 B.n386 10.6151
R1272 B.n386 B.n385 10.6151
R1273 B.n385 B.n382 10.6151
R1274 B.n382 B.n381 10.6151
R1275 B.n381 B.n378 10.6151
R1276 B.n378 B.n377 10.6151
R1277 B.n377 B.n374 10.6151
R1278 B.n374 B.n373 10.6151
R1279 B.n373 B.n370 10.6151
R1280 B.n370 B.n369 10.6151
R1281 B.n369 B.n366 10.6151
R1282 B.n366 B.n365 10.6151
R1283 B.n365 B.n362 10.6151
R1284 B.n360 B.n357 10.6151
R1285 B.n357 B.n356 10.6151
R1286 B.n356 B.n353 10.6151
R1287 B.n353 B.n352 10.6151
R1288 B.n352 B.n349 10.6151
R1289 B.n349 B.n348 10.6151
R1290 B.n348 B.n345 10.6151
R1291 B.n345 B.n344 10.6151
R1292 B.n344 B.n341 10.6151
R1293 B.n339 B.n336 10.6151
R1294 B.n336 B.n335 10.6151
R1295 B.n335 B.n332 10.6151
R1296 B.n332 B.n331 10.6151
R1297 B.n331 B.n328 10.6151
R1298 B.n328 B.n327 10.6151
R1299 B.n327 B.n324 10.6151
R1300 B.n324 B.n323 10.6151
R1301 B.n323 B.n320 10.6151
R1302 B.n320 B.n319 10.6151
R1303 B.n319 B.n316 10.6151
R1304 B.n316 B.n315 10.6151
R1305 B.n315 B.n312 10.6151
R1306 B.n312 B.n311 10.6151
R1307 B.n311 B.n308 10.6151
R1308 B.n308 B.n307 10.6151
R1309 B.n307 B.n304 10.6151
R1310 B.n304 B.n303 10.6151
R1311 B.n303 B.n300 10.6151
R1312 B.n300 B.n299 10.6151
R1313 B.n299 B.n296 10.6151
R1314 B.n296 B.n295 10.6151
R1315 B.n295 B.n292 10.6151
R1316 B.n292 B.n255 10.6151
R1317 B.n415 B.n255 10.6151
R1318 B.n417 B.n416 10.6151
R1319 B.n417 B.n247 10.6151
R1320 B.n427 B.n247 10.6151
R1321 B.n428 B.n427 10.6151
R1322 B.n429 B.n428 10.6151
R1323 B.n429 B.n240 10.6151
R1324 B.n440 B.n240 10.6151
R1325 B.n441 B.n440 10.6151
R1326 B.n442 B.n441 10.6151
R1327 B.n442 B.n232 10.6151
R1328 B.n452 B.n232 10.6151
R1329 B.n453 B.n452 10.6151
R1330 B.n454 B.n453 10.6151
R1331 B.n454 B.n224 10.6151
R1332 B.n464 B.n224 10.6151
R1333 B.n465 B.n464 10.6151
R1334 B.n466 B.n465 10.6151
R1335 B.n466 B.n216 10.6151
R1336 B.n476 B.n216 10.6151
R1337 B.n477 B.n476 10.6151
R1338 B.n479 B.n477 10.6151
R1339 B.n479 B.n478 10.6151
R1340 B.n478 B.n208 10.6151
R1341 B.n489 B.n208 10.6151
R1342 B.n490 B.n489 10.6151
R1343 B.n491 B.n490 10.6151
R1344 B.n492 B.n491 10.6151
R1345 B.n493 B.n492 10.6151
R1346 B.n496 B.n493 10.6151
R1347 B.n497 B.n496 10.6151
R1348 B.n498 B.n497 10.6151
R1349 B.n499 B.n498 10.6151
R1350 B.n501 B.n499 10.6151
R1351 B.n502 B.n501 10.6151
R1352 B.n503 B.n502 10.6151
R1353 B.n504 B.n503 10.6151
R1354 B.n506 B.n504 10.6151
R1355 B.n507 B.n506 10.6151
R1356 B.n508 B.n507 10.6151
R1357 B.n509 B.n508 10.6151
R1358 B.n511 B.n509 10.6151
R1359 B.n512 B.n511 10.6151
R1360 B.n513 B.n512 10.6151
R1361 B.n514 B.n513 10.6151
R1362 B.n516 B.n514 10.6151
R1363 B.n517 B.n516 10.6151
R1364 B.n518 B.n517 10.6151
R1365 B.n519 B.n518 10.6151
R1366 B.n521 B.n519 10.6151
R1367 B.n522 B.n521 10.6151
R1368 B.n523 B.n522 10.6151
R1369 B.n572 B.n1 10.6151
R1370 B.n572 B.n571 10.6151
R1371 B.n571 B.n570 10.6151
R1372 B.n570 B.n10 10.6151
R1373 B.n565 B.n10 10.6151
R1374 B.n565 B.n564 10.6151
R1375 B.n564 B.n563 10.6151
R1376 B.n563 B.n18 10.6151
R1377 B.n557 B.n18 10.6151
R1378 B.n557 B.n556 10.6151
R1379 B.n556 B.n555 10.6151
R1380 B.n555 B.n25 10.6151
R1381 B.n549 B.n25 10.6151
R1382 B.n549 B.n548 10.6151
R1383 B.n548 B.n547 10.6151
R1384 B.n547 B.n32 10.6151
R1385 B.n541 B.n32 10.6151
R1386 B.n541 B.n540 10.6151
R1387 B.n540 B.n539 10.6151
R1388 B.n539 B.n38 10.6151
R1389 B.n533 B.n38 10.6151
R1390 B.n533 B.n532 10.6151
R1391 B.n532 B.n531 10.6151
R1392 B.n531 B.n46 10.6151
R1393 B.n89 B.n88 10.6151
R1394 B.n92 B.n89 10.6151
R1395 B.n93 B.n92 10.6151
R1396 B.n96 B.n93 10.6151
R1397 B.n97 B.n96 10.6151
R1398 B.n100 B.n97 10.6151
R1399 B.n101 B.n100 10.6151
R1400 B.n104 B.n101 10.6151
R1401 B.n105 B.n104 10.6151
R1402 B.n108 B.n105 10.6151
R1403 B.n109 B.n108 10.6151
R1404 B.n112 B.n109 10.6151
R1405 B.n113 B.n112 10.6151
R1406 B.n116 B.n113 10.6151
R1407 B.n117 B.n116 10.6151
R1408 B.n120 B.n117 10.6151
R1409 B.n121 B.n120 10.6151
R1410 B.n124 B.n121 10.6151
R1411 B.n125 B.n124 10.6151
R1412 B.n128 B.n125 10.6151
R1413 B.n129 B.n128 10.6151
R1414 B.n132 B.n129 10.6151
R1415 B.n133 B.n132 10.6151
R1416 B.n136 B.n133 10.6151
R1417 B.n137 B.n136 10.6151
R1418 B.n141 B.n140 10.6151
R1419 B.n144 B.n141 10.6151
R1420 B.n145 B.n144 10.6151
R1421 B.n148 B.n145 10.6151
R1422 B.n149 B.n148 10.6151
R1423 B.n152 B.n149 10.6151
R1424 B.n153 B.n152 10.6151
R1425 B.n156 B.n153 10.6151
R1426 B.n157 B.n156 10.6151
R1427 B.n161 B.n160 10.6151
R1428 B.n164 B.n161 10.6151
R1429 B.n165 B.n164 10.6151
R1430 B.n168 B.n165 10.6151
R1431 B.n169 B.n168 10.6151
R1432 B.n172 B.n169 10.6151
R1433 B.n173 B.n172 10.6151
R1434 B.n176 B.n173 10.6151
R1435 B.n177 B.n176 10.6151
R1436 B.n180 B.n177 10.6151
R1437 B.n181 B.n180 10.6151
R1438 B.n184 B.n181 10.6151
R1439 B.n185 B.n184 10.6151
R1440 B.n188 B.n185 10.6151
R1441 B.n189 B.n188 10.6151
R1442 B.n192 B.n189 10.6151
R1443 B.n193 B.n192 10.6151
R1444 B.n196 B.n193 10.6151
R1445 B.n197 B.n196 10.6151
R1446 B.n200 B.n197 10.6151
R1447 B.n201 B.n200 10.6151
R1448 B.n204 B.n201 10.6151
R1449 B.n206 B.n204 10.6151
R1450 B.n207 B.n206 10.6151
R1451 B.n524 B.n207 10.6151
R1452 B.n362 B.n361 9.36635
R1453 B.n340 B.n339 9.36635
R1454 B.n137 B.n86 9.36635
R1455 B.n160 B.n83 9.36635
R1456 B.n580 B.n0 8.11757
R1457 B.n580 B.n1 8.11757
R1458 B.n361 B.n360 1.24928
R1459 B.n341 B.n340 1.24928
R1460 B.n140 B.n86 1.24928
R1461 B.n157 B.n83 1.24928
R1462 VN.n0 VN.t3 136.898
R1463 VN.n1 VN.t2 136.898
R1464 VN.n0 VN.t0 136.569
R1465 VN.n1 VN.t1 136.569
R1466 VN VN.n1 52.2664
R1467 VN VN.n0 12.5505
R1468 VDD2.n2 VDD2.n0 100.272
R1469 VDD2.n2 VDD2.n1 65.6861
R1470 VDD2.n1 VDD2.t2 2.95572
R1471 VDD2.n1 VDD2.t1 2.95572
R1472 VDD2.n0 VDD2.t0 2.95572
R1473 VDD2.n0 VDD2.t3 2.95572
R1474 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 2.59875f
C1 VDD1 VP 2.71308f
C2 VTAIL VP 2.61286f
C3 VDD2 VN 2.52849f
C4 VDD2 VP 0.333672f
C5 VDD1 VTAIL 3.93482f
C6 VDD2 VDD1 0.794225f
C7 VDD2 VTAIL 3.98259f
C8 VN VP 4.51089f
C9 VDD1 VN 0.148586f
C10 VDD2 B 2.812079f
C11 VDD1 B 6.04128f
C12 VTAIL B 6.185709f
C13 VN B 8.46262f
C14 VP B 6.42299f
C15 VDD2.t0 B 0.142642f
C16 VDD2.t3 B 0.142642f
C17 VDD2.n0 B 1.642f
C18 VDD2.t2 B 0.142642f
C19 VDD2.t1 B 0.142642f
C20 VDD2.n1 B 1.20469f
C21 VDD2.n2 B 2.92951f
C22 VN.t3 B 1.19455f
C23 VN.t0 B 1.19323f
C24 VN.n0 B 0.857502f
C25 VN.t2 B 1.19455f
C26 VN.t1 B 1.19323f
C27 VN.n1 B 2.02665f
C28 VDD1.t1 B 0.142653f
C29 VDD1.t3 B 0.142653f
C30 VDD1.n0 B 1.20512f
C31 VDD1.t2 B 0.142653f
C32 VDD1.t0 B 0.142653f
C33 VDD1.n1 B 1.66551f
C34 VTAIL.n0 B 0.025517f
C35 VTAIL.n1 B 0.017981f
C36 VTAIL.n2 B 0.009662f
C37 VTAIL.n3 B 0.022838f
C38 VTAIL.n4 B 0.010231f
C39 VTAIL.n5 B 0.017981f
C40 VTAIL.n6 B 0.009662f
C41 VTAIL.n7 B 0.022838f
C42 VTAIL.n8 B 0.010231f
C43 VTAIL.n9 B 0.485712f
C44 VTAIL.n10 B 0.009662f
C45 VTAIL.t7 B 0.037208f
C46 VTAIL.n11 B 0.079987f
C47 VTAIL.n12 B 0.013491f
C48 VTAIL.n13 B 0.017129f
C49 VTAIL.n14 B 0.022838f
C50 VTAIL.n15 B 0.010231f
C51 VTAIL.n16 B 0.009662f
C52 VTAIL.n17 B 0.017981f
C53 VTAIL.n18 B 0.017981f
C54 VTAIL.n19 B 0.009662f
C55 VTAIL.n20 B 0.010231f
C56 VTAIL.n21 B 0.022838f
C57 VTAIL.n22 B 0.022838f
C58 VTAIL.n23 B 0.010231f
C59 VTAIL.n24 B 0.009662f
C60 VTAIL.n25 B 0.017981f
C61 VTAIL.n26 B 0.017981f
C62 VTAIL.n27 B 0.009662f
C63 VTAIL.n28 B 0.010231f
C64 VTAIL.n29 B 0.022838f
C65 VTAIL.n30 B 0.049871f
C66 VTAIL.n31 B 0.010231f
C67 VTAIL.n32 B 0.009662f
C68 VTAIL.n33 B 0.041072f
C69 VTAIL.n34 B 0.027933f
C70 VTAIL.n35 B 0.094873f
C71 VTAIL.n36 B 0.025517f
C72 VTAIL.n37 B 0.017981f
C73 VTAIL.n38 B 0.009662f
C74 VTAIL.n39 B 0.022838f
C75 VTAIL.n40 B 0.010231f
C76 VTAIL.n41 B 0.017981f
C77 VTAIL.n42 B 0.009662f
C78 VTAIL.n43 B 0.022838f
C79 VTAIL.n44 B 0.010231f
C80 VTAIL.n45 B 0.485712f
C81 VTAIL.n46 B 0.009662f
C82 VTAIL.t2 B 0.037208f
C83 VTAIL.n47 B 0.079987f
C84 VTAIL.n48 B 0.013491f
C85 VTAIL.n49 B 0.017129f
C86 VTAIL.n50 B 0.022838f
C87 VTAIL.n51 B 0.010231f
C88 VTAIL.n52 B 0.009662f
C89 VTAIL.n53 B 0.017981f
C90 VTAIL.n54 B 0.017981f
C91 VTAIL.n55 B 0.009662f
C92 VTAIL.n56 B 0.010231f
C93 VTAIL.n57 B 0.022838f
C94 VTAIL.n58 B 0.022838f
C95 VTAIL.n59 B 0.010231f
C96 VTAIL.n60 B 0.009662f
C97 VTAIL.n61 B 0.017981f
C98 VTAIL.n62 B 0.017981f
C99 VTAIL.n63 B 0.009662f
C100 VTAIL.n64 B 0.010231f
C101 VTAIL.n65 B 0.022838f
C102 VTAIL.n66 B 0.049871f
C103 VTAIL.n67 B 0.010231f
C104 VTAIL.n68 B 0.009662f
C105 VTAIL.n69 B 0.041072f
C106 VTAIL.n70 B 0.027933f
C107 VTAIL.n71 B 0.140701f
C108 VTAIL.n72 B 0.025517f
C109 VTAIL.n73 B 0.017981f
C110 VTAIL.n74 B 0.009662f
C111 VTAIL.n75 B 0.022838f
C112 VTAIL.n76 B 0.010231f
C113 VTAIL.n77 B 0.017981f
C114 VTAIL.n78 B 0.009662f
C115 VTAIL.n79 B 0.022838f
C116 VTAIL.n80 B 0.010231f
C117 VTAIL.n81 B 0.485712f
C118 VTAIL.n82 B 0.009662f
C119 VTAIL.t5 B 0.037208f
C120 VTAIL.n83 B 0.079987f
C121 VTAIL.n84 B 0.013491f
C122 VTAIL.n85 B 0.017129f
C123 VTAIL.n86 B 0.022838f
C124 VTAIL.n87 B 0.010231f
C125 VTAIL.n88 B 0.009662f
C126 VTAIL.n89 B 0.017981f
C127 VTAIL.n90 B 0.017981f
C128 VTAIL.n91 B 0.009662f
C129 VTAIL.n92 B 0.010231f
C130 VTAIL.n93 B 0.022838f
C131 VTAIL.n94 B 0.022838f
C132 VTAIL.n95 B 0.010231f
C133 VTAIL.n96 B 0.009662f
C134 VTAIL.n97 B 0.017981f
C135 VTAIL.n98 B 0.017981f
C136 VTAIL.n99 B 0.009662f
C137 VTAIL.n100 B 0.010231f
C138 VTAIL.n101 B 0.022838f
C139 VTAIL.n102 B 0.049871f
C140 VTAIL.n103 B 0.010231f
C141 VTAIL.n104 B 0.009662f
C142 VTAIL.n105 B 0.041072f
C143 VTAIL.n106 B 0.027933f
C144 VTAIL.n107 B 0.790788f
C145 VTAIL.n108 B 0.025517f
C146 VTAIL.n109 B 0.017981f
C147 VTAIL.n110 B 0.009662f
C148 VTAIL.n111 B 0.022838f
C149 VTAIL.n112 B 0.010231f
C150 VTAIL.n113 B 0.017981f
C151 VTAIL.n114 B 0.009662f
C152 VTAIL.n115 B 0.022838f
C153 VTAIL.n116 B 0.010231f
C154 VTAIL.n117 B 0.485712f
C155 VTAIL.n118 B 0.009662f
C156 VTAIL.t1 B 0.037208f
C157 VTAIL.n119 B 0.079987f
C158 VTAIL.n120 B 0.013491f
C159 VTAIL.n121 B 0.017129f
C160 VTAIL.n122 B 0.022838f
C161 VTAIL.n123 B 0.010231f
C162 VTAIL.n124 B 0.009662f
C163 VTAIL.n125 B 0.017981f
C164 VTAIL.n126 B 0.017981f
C165 VTAIL.n127 B 0.009662f
C166 VTAIL.n128 B 0.010231f
C167 VTAIL.n129 B 0.022838f
C168 VTAIL.n130 B 0.022838f
C169 VTAIL.n131 B 0.010231f
C170 VTAIL.n132 B 0.009662f
C171 VTAIL.n133 B 0.017981f
C172 VTAIL.n134 B 0.017981f
C173 VTAIL.n135 B 0.009662f
C174 VTAIL.n136 B 0.010231f
C175 VTAIL.n137 B 0.022838f
C176 VTAIL.n138 B 0.049871f
C177 VTAIL.n139 B 0.010231f
C178 VTAIL.n140 B 0.009662f
C179 VTAIL.n141 B 0.041072f
C180 VTAIL.n142 B 0.027933f
C181 VTAIL.n143 B 0.790788f
C182 VTAIL.n144 B 0.025517f
C183 VTAIL.n145 B 0.017981f
C184 VTAIL.n146 B 0.009662f
C185 VTAIL.n147 B 0.022838f
C186 VTAIL.n148 B 0.010231f
C187 VTAIL.n149 B 0.017981f
C188 VTAIL.n150 B 0.009662f
C189 VTAIL.n151 B 0.022838f
C190 VTAIL.n152 B 0.010231f
C191 VTAIL.n153 B 0.485712f
C192 VTAIL.n154 B 0.009662f
C193 VTAIL.t0 B 0.037208f
C194 VTAIL.n155 B 0.079987f
C195 VTAIL.n156 B 0.013491f
C196 VTAIL.n157 B 0.017129f
C197 VTAIL.n158 B 0.022838f
C198 VTAIL.n159 B 0.010231f
C199 VTAIL.n160 B 0.009662f
C200 VTAIL.n161 B 0.017981f
C201 VTAIL.n162 B 0.017981f
C202 VTAIL.n163 B 0.009662f
C203 VTAIL.n164 B 0.010231f
C204 VTAIL.n165 B 0.022838f
C205 VTAIL.n166 B 0.022838f
C206 VTAIL.n167 B 0.010231f
C207 VTAIL.n168 B 0.009662f
C208 VTAIL.n169 B 0.017981f
C209 VTAIL.n170 B 0.017981f
C210 VTAIL.n171 B 0.009662f
C211 VTAIL.n172 B 0.010231f
C212 VTAIL.n173 B 0.022838f
C213 VTAIL.n174 B 0.049871f
C214 VTAIL.n175 B 0.010231f
C215 VTAIL.n176 B 0.009662f
C216 VTAIL.n177 B 0.041072f
C217 VTAIL.n178 B 0.027933f
C218 VTAIL.n179 B 0.140701f
C219 VTAIL.n180 B 0.025517f
C220 VTAIL.n181 B 0.017981f
C221 VTAIL.n182 B 0.009662f
C222 VTAIL.n183 B 0.022838f
C223 VTAIL.n184 B 0.010231f
C224 VTAIL.n185 B 0.017981f
C225 VTAIL.n186 B 0.009662f
C226 VTAIL.n187 B 0.022838f
C227 VTAIL.n188 B 0.010231f
C228 VTAIL.n189 B 0.485712f
C229 VTAIL.n190 B 0.009662f
C230 VTAIL.t4 B 0.037208f
C231 VTAIL.n191 B 0.079987f
C232 VTAIL.n192 B 0.013491f
C233 VTAIL.n193 B 0.017129f
C234 VTAIL.n194 B 0.022838f
C235 VTAIL.n195 B 0.010231f
C236 VTAIL.n196 B 0.009662f
C237 VTAIL.n197 B 0.017981f
C238 VTAIL.n198 B 0.017981f
C239 VTAIL.n199 B 0.009662f
C240 VTAIL.n200 B 0.010231f
C241 VTAIL.n201 B 0.022838f
C242 VTAIL.n202 B 0.022838f
C243 VTAIL.n203 B 0.010231f
C244 VTAIL.n204 B 0.009662f
C245 VTAIL.n205 B 0.017981f
C246 VTAIL.n206 B 0.017981f
C247 VTAIL.n207 B 0.009662f
C248 VTAIL.n208 B 0.010231f
C249 VTAIL.n209 B 0.022838f
C250 VTAIL.n210 B 0.049871f
C251 VTAIL.n211 B 0.010231f
C252 VTAIL.n212 B 0.009662f
C253 VTAIL.n213 B 0.041072f
C254 VTAIL.n214 B 0.027933f
C255 VTAIL.n215 B 0.140701f
C256 VTAIL.n216 B 0.025517f
C257 VTAIL.n217 B 0.017981f
C258 VTAIL.n218 B 0.009662f
C259 VTAIL.n219 B 0.022838f
C260 VTAIL.n220 B 0.010231f
C261 VTAIL.n221 B 0.017981f
C262 VTAIL.n222 B 0.009662f
C263 VTAIL.n223 B 0.022838f
C264 VTAIL.n224 B 0.010231f
C265 VTAIL.n225 B 0.485712f
C266 VTAIL.n226 B 0.009662f
C267 VTAIL.t3 B 0.037208f
C268 VTAIL.n227 B 0.079987f
C269 VTAIL.n228 B 0.013491f
C270 VTAIL.n229 B 0.017129f
C271 VTAIL.n230 B 0.022838f
C272 VTAIL.n231 B 0.010231f
C273 VTAIL.n232 B 0.009662f
C274 VTAIL.n233 B 0.017981f
C275 VTAIL.n234 B 0.017981f
C276 VTAIL.n235 B 0.009662f
C277 VTAIL.n236 B 0.010231f
C278 VTAIL.n237 B 0.022838f
C279 VTAIL.n238 B 0.022838f
C280 VTAIL.n239 B 0.010231f
C281 VTAIL.n240 B 0.009662f
C282 VTAIL.n241 B 0.017981f
C283 VTAIL.n242 B 0.017981f
C284 VTAIL.n243 B 0.009662f
C285 VTAIL.n244 B 0.010231f
C286 VTAIL.n245 B 0.022838f
C287 VTAIL.n246 B 0.049871f
C288 VTAIL.n247 B 0.010231f
C289 VTAIL.n248 B 0.009662f
C290 VTAIL.n249 B 0.041072f
C291 VTAIL.n250 B 0.027933f
C292 VTAIL.n251 B 0.790788f
C293 VTAIL.n252 B 0.025517f
C294 VTAIL.n253 B 0.017981f
C295 VTAIL.n254 B 0.009662f
C296 VTAIL.n255 B 0.022838f
C297 VTAIL.n256 B 0.010231f
C298 VTAIL.n257 B 0.017981f
C299 VTAIL.n258 B 0.009662f
C300 VTAIL.n259 B 0.022838f
C301 VTAIL.n260 B 0.010231f
C302 VTAIL.n261 B 0.485712f
C303 VTAIL.n262 B 0.009662f
C304 VTAIL.t6 B 0.037208f
C305 VTAIL.n263 B 0.079987f
C306 VTAIL.n264 B 0.013491f
C307 VTAIL.n265 B 0.017129f
C308 VTAIL.n266 B 0.022838f
C309 VTAIL.n267 B 0.010231f
C310 VTAIL.n268 B 0.009662f
C311 VTAIL.n269 B 0.017981f
C312 VTAIL.n270 B 0.017981f
C313 VTAIL.n271 B 0.009662f
C314 VTAIL.n272 B 0.010231f
C315 VTAIL.n273 B 0.022838f
C316 VTAIL.n274 B 0.022838f
C317 VTAIL.n275 B 0.010231f
C318 VTAIL.n276 B 0.009662f
C319 VTAIL.n277 B 0.017981f
C320 VTAIL.n278 B 0.017981f
C321 VTAIL.n279 B 0.009662f
C322 VTAIL.n280 B 0.010231f
C323 VTAIL.n281 B 0.022838f
C324 VTAIL.n282 B 0.049871f
C325 VTAIL.n283 B 0.010231f
C326 VTAIL.n284 B 0.009662f
C327 VTAIL.n285 B 0.041072f
C328 VTAIL.n286 B 0.027933f
C329 VTAIL.n287 B 0.738218f
C330 VP.n0 B 0.036448f
C331 VP.t3 B 1.06652f
C332 VP.n1 B 0.052983f
C333 VP.t2 B 1.22582f
C334 VP.t0 B 1.22445f
C335 VP.n2 B 2.05869f
C336 VP.n3 B 1.763f
C337 VP.t1 B 1.06652f
C338 VP.n4 B 0.493178f
C339 VP.n5 B 0.049905f
C340 VP.n6 B 0.036448f
C341 VP.n7 B 0.036448f
C342 VP.n8 B 0.036448f
C343 VP.n9 B 0.052983f
C344 VP.n10 B 0.049905f
C345 VP.n11 B 0.493178f
C346 VP.n12 B 0.03517f
.ends

