* NGSPICE file created from diff_pair_sample_0648.ext - technology: sky130A

.subckt diff_pair_sample_0648 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=0 ps=0 w=18.95 l=0.94
X1 VDD2.t3 VN.t0 VTAIL.t6 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=3.12675 pd=19.28 as=7.3905 ps=38.68 w=18.95 l=0.94
X2 VTAIL.t1 VP.t0 VDD1.t3 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=3.12675 ps=19.28 w=18.95 l=0.94
X3 VTAIL.t4 VN.t1 VDD2.t2 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=3.12675 ps=19.28 w=18.95 l=0.94
X4 VDD2.t1 VN.t2 VTAIL.t7 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=3.12675 pd=19.28 as=7.3905 ps=38.68 w=18.95 l=0.94
X5 VDD1.t2 VP.t1 VTAIL.t2 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=3.12675 pd=19.28 as=7.3905 ps=38.68 w=18.95 l=0.94
X6 VTAIL.t0 VP.t2 VDD1.t1 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=3.12675 ps=19.28 w=18.95 l=0.94
X7 B.t8 B.t6 B.t7 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=0 ps=0 w=18.95 l=0.94
X8 VDD1.t0 VP.t3 VTAIL.t3 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=3.12675 pd=19.28 as=7.3905 ps=38.68 w=18.95 l=0.94
X9 B.t5 B.t3 B.t4 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=0 ps=0 w=18.95 l=0.94
X10 B.t2 B.t0 B.t1 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=0 ps=0 w=18.95 l=0.94
X11 VTAIL.t5 VN.t3 VDD2.t0 w_n1732_n4758# sky130_fd_pr__pfet_01v8 ad=7.3905 pd=38.68 as=3.12675 ps=19.28 w=18.95 l=0.94
R0 B.n300 B.t9 688.346
R1 B.n135 B.t6 688.346
R2 B.n51 B.t3 688.346
R3 B.n44 B.t0 688.346
R4 B.n413 B.n412 585
R5 B.n411 B.n104 585
R6 B.n410 B.n409 585
R7 B.n408 B.n105 585
R8 B.n407 B.n406 585
R9 B.n405 B.n106 585
R10 B.n404 B.n403 585
R11 B.n402 B.n107 585
R12 B.n401 B.n400 585
R13 B.n399 B.n108 585
R14 B.n398 B.n397 585
R15 B.n396 B.n109 585
R16 B.n395 B.n394 585
R17 B.n393 B.n110 585
R18 B.n392 B.n391 585
R19 B.n390 B.n111 585
R20 B.n389 B.n388 585
R21 B.n387 B.n112 585
R22 B.n386 B.n385 585
R23 B.n384 B.n113 585
R24 B.n383 B.n382 585
R25 B.n381 B.n114 585
R26 B.n380 B.n379 585
R27 B.n378 B.n115 585
R28 B.n377 B.n376 585
R29 B.n375 B.n116 585
R30 B.n374 B.n373 585
R31 B.n372 B.n117 585
R32 B.n371 B.n370 585
R33 B.n369 B.n118 585
R34 B.n368 B.n367 585
R35 B.n366 B.n119 585
R36 B.n365 B.n364 585
R37 B.n363 B.n120 585
R38 B.n362 B.n361 585
R39 B.n360 B.n121 585
R40 B.n359 B.n358 585
R41 B.n357 B.n122 585
R42 B.n356 B.n355 585
R43 B.n354 B.n123 585
R44 B.n353 B.n352 585
R45 B.n351 B.n124 585
R46 B.n350 B.n349 585
R47 B.n348 B.n125 585
R48 B.n347 B.n346 585
R49 B.n345 B.n126 585
R50 B.n344 B.n343 585
R51 B.n342 B.n127 585
R52 B.n341 B.n340 585
R53 B.n339 B.n128 585
R54 B.n338 B.n337 585
R55 B.n336 B.n129 585
R56 B.n335 B.n334 585
R57 B.n333 B.n130 585
R58 B.n332 B.n331 585
R59 B.n330 B.n131 585
R60 B.n329 B.n328 585
R61 B.n327 B.n132 585
R62 B.n326 B.n325 585
R63 B.n324 B.n133 585
R64 B.n323 B.n322 585
R65 B.n321 B.n134 585
R66 B.n319 B.n318 585
R67 B.n317 B.n137 585
R68 B.n316 B.n315 585
R69 B.n314 B.n138 585
R70 B.n313 B.n312 585
R71 B.n311 B.n139 585
R72 B.n310 B.n309 585
R73 B.n308 B.n140 585
R74 B.n307 B.n306 585
R75 B.n305 B.n141 585
R76 B.n304 B.n303 585
R77 B.n299 B.n142 585
R78 B.n298 B.n297 585
R79 B.n296 B.n143 585
R80 B.n295 B.n294 585
R81 B.n293 B.n144 585
R82 B.n292 B.n291 585
R83 B.n290 B.n145 585
R84 B.n289 B.n288 585
R85 B.n287 B.n146 585
R86 B.n286 B.n285 585
R87 B.n284 B.n147 585
R88 B.n283 B.n282 585
R89 B.n281 B.n148 585
R90 B.n280 B.n279 585
R91 B.n278 B.n149 585
R92 B.n277 B.n276 585
R93 B.n275 B.n150 585
R94 B.n274 B.n273 585
R95 B.n272 B.n151 585
R96 B.n271 B.n270 585
R97 B.n269 B.n152 585
R98 B.n268 B.n267 585
R99 B.n266 B.n153 585
R100 B.n265 B.n264 585
R101 B.n263 B.n154 585
R102 B.n262 B.n261 585
R103 B.n260 B.n155 585
R104 B.n259 B.n258 585
R105 B.n257 B.n156 585
R106 B.n256 B.n255 585
R107 B.n254 B.n157 585
R108 B.n253 B.n252 585
R109 B.n251 B.n158 585
R110 B.n250 B.n249 585
R111 B.n248 B.n159 585
R112 B.n247 B.n246 585
R113 B.n245 B.n160 585
R114 B.n244 B.n243 585
R115 B.n242 B.n161 585
R116 B.n241 B.n240 585
R117 B.n239 B.n162 585
R118 B.n238 B.n237 585
R119 B.n236 B.n163 585
R120 B.n235 B.n234 585
R121 B.n233 B.n164 585
R122 B.n232 B.n231 585
R123 B.n230 B.n165 585
R124 B.n229 B.n228 585
R125 B.n227 B.n166 585
R126 B.n226 B.n225 585
R127 B.n224 B.n167 585
R128 B.n223 B.n222 585
R129 B.n221 B.n168 585
R130 B.n220 B.n219 585
R131 B.n218 B.n169 585
R132 B.n217 B.n216 585
R133 B.n215 B.n170 585
R134 B.n214 B.n213 585
R135 B.n212 B.n171 585
R136 B.n211 B.n210 585
R137 B.n209 B.n172 585
R138 B.n414 B.n103 585
R139 B.n416 B.n415 585
R140 B.n417 B.n102 585
R141 B.n419 B.n418 585
R142 B.n420 B.n101 585
R143 B.n422 B.n421 585
R144 B.n423 B.n100 585
R145 B.n425 B.n424 585
R146 B.n426 B.n99 585
R147 B.n428 B.n427 585
R148 B.n429 B.n98 585
R149 B.n431 B.n430 585
R150 B.n432 B.n97 585
R151 B.n434 B.n433 585
R152 B.n435 B.n96 585
R153 B.n437 B.n436 585
R154 B.n438 B.n95 585
R155 B.n440 B.n439 585
R156 B.n441 B.n94 585
R157 B.n443 B.n442 585
R158 B.n444 B.n93 585
R159 B.n446 B.n445 585
R160 B.n447 B.n92 585
R161 B.n449 B.n448 585
R162 B.n450 B.n91 585
R163 B.n452 B.n451 585
R164 B.n453 B.n90 585
R165 B.n455 B.n454 585
R166 B.n456 B.n89 585
R167 B.n458 B.n457 585
R168 B.n459 B.n88 585
R169 B.n461 B.n460 585
R170 B.n462 B.n87 585
R171 B.n464 B.n463 585
R172 B.n465 B.n86 585
R173 B.n467 B.n466 585
R174 B.n468 B.n85 585
R175 B.n470 B.n469 585
R176 B.n471 B.n84 585
R177 B.n473 B.n472 585
R178 B.n675 B.n674 585
R179 B.n673 B.n12 585
R180 B.n672 B.n671 585
R181 B.n670 B.n13 585
R182 B.n669 B.n668 585
R183 B.n667 B.n14 585
R184 B.n666 B.n665 585
R185 B.n664 B.n15 585
R186 B.n663 B.n662 585
R187 B.n661 B.n16 585
R188 B.n660 B.n659 585
R189 B.n658 B.n17 585
R190 B.n657 B.n656 585
R191 B.n655 B.n18 585
R192 B.n654 B.n653 585
R193 B.n652 B.n19 585
R194 B.n651 B.n650 585
R195 B.n649 B.n20 585
R196 B.n648 B.n647 585
R197 B.n646 B.n21 585
R198 B.n645 B.n644 585
R199 B.n643 B.n22 585
R200 B.n642 B.n641 585
R201 B.n640 B.n23 585
R202 B.n639 B.n638 585
R203 B.n637 B.n24 585
R204 B.n636 B.n635 585
R205 B.n634 B.n25 585
R206 B.n633 B.n632 585
R207 B.n631 B.n26 585
R208 B.n630 B.n629 585
R209 B.n628 B.n27 585
R210 B.n627 B.n626 585
R211 B.n625 B.n28 585
R212 B.n624 B.n623 585
R213 B.n622 B.n29 585
R214 B.n621 B.n620 585
R215 B.n619 B.n30 585
R216 B.n618 B.n617 585
R217 B.n616 B.n31 585
R218 B.n615 B.n614 585
R219 B.n613 B.n32 585
R220 B.n612 B.n611 585
R221 B.n610 B.n33 585
R222 B.n609 B.n608 585
R223 B.n607 B.n34 585
R224 B.n606 B.n605 585
R225 B.n604 B.n35 585
R226 B.n603 B.n602 585
R227 B.n601 B.n36 585
R228 B.n600 B.n599 585
R229 B.n598 B.n37 585
R230 B.n597 B.n596 585
R231 B.n595 B.n38 585
R232 B.n594 B.n593 585
R233 B.n592 B.n39 585
R234 B.n591 B.n590 585
R235 B.n589 B.n40 585
R236 B.n588 B.n587 585
R237 B.n586 B.n41 585
R238 B.n585 B.n584 585
R239 B.n583 B.n42 585
R240 B.n582 B.n581 585
R241 B.n580 B.n43 585
R242 B.n579 B.n578 585
R243 B.n577 B.n47 585
R244 B.n576 B.n575 585
R245 B.n574 B.n48 585
R246 B.n573 B.n572 585
R247 B.n571 B.n49 585
R248 B.n570 B.n569 585
R249 B.n568 B.n50 585
R250 B.n566 B.n565 585
R251 B.n564 B.n53 585
R252 B.n563 B.n562 585
R253 B.n561 B.n54 585
R254 B.n560 B.n559 585
R255 B.n558 B.n55 585
R256 B.n557 B.n556 585
R257 B.n555 B.n56 585
R258 B.n554 B.n553 585
R259 B.n552 B.n57 585
R260 B.n551 B.n550 585
R261 B.n549 B.n58 585
R262 B.n548 B.n547 585
R263 B.n546 B.n59 585
R264 B.n545 B.n544 585
R265 B.n543 B.n60 585
R266 B.n542 B.n541 585
R267 B.n540 B.n61 585
R268 B.n539 B.n538 585
R269 B.n537 B.n62 585
R270 B.n536 B.n535 585
R271 B.n534 B.n63 585
R272 B.n533 B.n532 585
R273 B.n531 B.n64 585
R274 B.n530 B.n529 585
R275 B.n528 B.n65 585
R276 B.n527 B.n526 585
R277 B.n525 B.n66 585
R278 B.n524 B.n523 585
R279 B.n522 B.n67 585
R280 B.n521 B.n520 585
R281 B.n519 B.n68 585
R282 B.n518 B.n517 585
R283 B.n516 B.n69 585
R284 B.n515 B.n514 585
R285 B.n513 B.n70 585
R286 B.n512 B.n511 585
R287 B.n510 B.n71 585
R288 B.n509 B.n508 585
R289 B.n507 B.n72 585
R290 B.n506 B.n505 585
R291 B.n504 B.n73 585
R292 B.n503 B.n502 585
R293 B.n501 B.n74 585
R294 B.n500 B.n499 585
R295 B.n498 B.n75 585
R296 B.n497 B.n496 585
R297 B.n495 B.n76 585
R298 B.n494 B.n493 585
R299 B.n492 B.n77 585
R300 B.n491 B.n490 585
R301 B.n489 B.n78 585
R302 B.n488 B.n487 585
R303 B.n486 B.n79 585
R304 B.n485 B.n484 585
R305 B.n483 B.n80 585
R306 B.n482 B.n481 585
R307 B.n480 B.n81 585
R308 B.n479 B.n478 585
R309 B.n477 B.n82 585
R310 B.n476 B.n475 585
R311 B.n474 B.n83 585
R312 B.n676 B.n11 585
R313 B.n678 B.n677 585
R314 B.n679 B.n10 585
R315 B.n681 B.n680 585
R316 B.n682 B.n9 585
R317 B.n684 B.n683 585
R318 B.n685 B.n8 585
R319 B.n687 B.n686 585
R320 B.n688 B.n7 585
R321 B.n690 B.n689 585
R322 B.n691 B.n6 585
R323 B.n693 B.n692 585
R324 B.n694 B.n5 585
R325 B.n696 B.n695 585
R326 B.n697 B.n4 585
R327 B.n699 B.n698 585
R328 B.n700 B.n3 585
R329 B.n702 B.n701 585
R330 B.n703 B.n0 585
R331 B.n2 B.n1 585
R332 B.n182 B.n181 585
R333 B.n184 B.n183 585
R334 B.n185 B.n180 585
R335 B.n187 B.n186 585
R336 B.n188 B.n179 585
R337 B.n190 B.n189 585
R338 B.n191 B.n178 585
R339 B.n193 B.n192 585
R340 B.n194 B.n177 585
R341 B.n196 B.n195 585
R342 B.n197 B.n176 585
R343 B.n199 B.n198 585
R344 B.n200 B.n175 585
R345 B.n202 B.n201 585
R346 B.n203 B.n174 585
R347 B.n205 B.n204 585
R348 B.n206 B.n173 585
R349 B.n208 B.n207 585
R350 B.n135 B.t7 525.549
R351 B.n51 B.t5 525.549
R352 B.n300 B.t10 525.549
R353 B.n44 B.t2 525.549
R354 B.n136 B.t8 500.92
R355 B.n52 B.t4 500.92
R356 B.n301 B.t11 500.918
R357 B.n45 B.t1 500.918
R358 B.n207 B.n172 444.452
R359 B.n414 B.n413 444.452
R360 B.n474 B.n473 444.452
R361 B.n674 B.n11 444.452
R362 B.n705 B.n704 256.663
R363 B.n704 B.n703 235.042
R364 B.n704 B.n2 235.042
R365 B.n211 B.n172 163.367
R366 B.n212 B.n211 163.367
R367 B.n213 B.n212 163.367
R368 B.n213 B.n170 163.367
R369 B.n217 B.n170 163.367
R370 B.n218 B.n217 163.367
R371 B.n219 B.n218 163.367
R372 B.n219 B.n168 163.367
R373 B.n223 B.n168 163.367
R374 B.n224 B.n223 163.367
R375 B.n225 B.n224 163.367
R376 B.n225 B.n166 163.367
R377 B.n229 B.n166 163.367
R378 B.n230 B.n229 163.367
R379 B.n231 B.n230 163.367
R380 B.n231 B.n164 163.367
R381 B.n235 B.n164 163.367
R382 B.n236 B.n235 163.367
R383 B.n237 B.n236 163.367
R384 B.n237 B.n162 163.367
R385 B.n241 B.n162 163.367
R386 B.n242 B.n241 163.367
R387 B.n243 B.n242 163.367
R388 B.n243 B.n160 163.367
R389 B.n247 B.n160 163.367
R390 B.n248 B.n247 163.367
R391 B.n249 B.n248 163.367
R392 B.n249 B.n158 163.367
R393 B.n253 B.n158 163.367
R394 B.n254 B.n253 163.367
R395 B.n255 B.n254 163.367
R396 B.n255 B.n156 163.367
R397 B.n259 B.n156 163.367
R398 B.n260 B.n259 163.367
R399 B.n261 B.n260 163.367
R400 B.n261 B.n154 163.367
R401 B.n265 B.n154 163.367
R402 B.n266 B.n265 163.367
R403 B.n267 B.n266 163.367
R404 B.n267 B.n152 163.367
R405 B.n271 B.n152 163.367
R406 B.n272 B.n271 163.367
R407 B.n273 B.n272 163.367
R408 B.n273 B.n150 163.367
R409 B.n277 B.n150 163.367
R410 B.n278 B.n277 163.367
R411 B.n279 B.n278 163.367
R412 B.n279 B.n148 163.367
R413 B.n283 B.n148 163.367
R414 B.n284 B.n283 163.367
R415 B.n285 B.n284 163.367
R416 B.n285 B.n146 163.367
R417 B.n289 B.n146 163.367
R418 B.n290 B.n289 163.367
R419 B.n291 B.n290 163.367
R420 B.n291 B.n144 163.367
R421 B.n295 B.n144 163.367
R422 B.n296 B.n295 163.367
R423 B.n297 B.n296 163.367
R424 B.n297 B.n142 163.367
R425 B.n304 B.n142 163.367
R426 B.n305 B.n304 163.367
R427 B.n306 B.n305 163.367
R428 B.n306 B.n140 163.367
R429 B.n310 B.n140 163.367
R430 B.n311 B.n310 163.367
R431 B.n312 B.n311 163.367
R432 B.n312 B.n138 163.367
R433 B.n316 B.n138 163.367
R434 B.n317 B.n316 163.367
R435 B.n318 B.n317 163.367
R436 B.n318 B.n134 163.367
R437 B.n323 B.n134 163.367
R438 B.n324 B.n323 163.367
R439 B.n325 B.n324 163.367
R440 B.n325 B.n132 163.367
R441 B.n329 B.n132 163.367
R442 B.n330 B.n329 163.367
R443 B.n331 B.n330 163.367
R444 B.n331 B.n130 163.367
R445 B.n335 B.n130 163.367
R446 B.n336 B.n335 163.367
R447 B.n337 B.n336 163.367
R448 B.n337 B.n128 163.367
R449 B.n341 B.n128 163.367
R450 B.n342 B.n341 163.367
R451 B.n343 B.n342 163.367
R452 B.n343 B.n126 163.367
R453 B.n347 B.n126 163.367
R454 B.n348 B.n347 163.367
R455 B.n349 B.n348 163.367
R456 B.n349 B.n124 163.367
R457 B.n353 B.n124 163.367
R458 B.n354 B.n353 163.367
R459 B.n355 B.n354 163.367
R460 B.n355 B.n122 163.367
R461 B.n359 B.n122 163.367
R462 B.n360 B.n359 163.367
R463 B.n361 B.n360 163.367
R464 B.n361 B.n120 163.367
R465 B.n365 B.n120 163.367
R466 B.n366 B.n365 163.367
R467 B.n367 B.n366 163.367
R468 B.n367 B.n118 163.367
R469 B.n371 B.n118 163.367
R470 B.n372 B.n371 163.367
R471 B.n373 B.n372 163.367
R472 B.n373 B.n116 163.367
R473 B.n377 B.n116 163.367
R474 B.n378 B.n377 163.367
R475 B.n379 B.n378 163.367
R476 B.n379 B.n114 163.367
R477 B.n383 B.n114 163.367
R478 B.n384 B.n383 163.367
R479 B.n385 B.n384 163.367
R480 B.n385 B.n112 163.367
R481 B.n389 B.n112 163.367
R482 B.n390 B.n389 163.367
R483 B.n391 B.n390 163.367
R484 B.n391 B.n110 163.367
R485 B.n395 B.n110 163.367
R486 B.n396 B.n395 163.367
R487 B.n397 B.n396 163.367
R488 B.n397 B.n108 163.367
R489 B.n401 B.n108 163.367
R490 B.n402 B.n401 163.367
R491 B.n403 B.n402 163.367
R492 B.n403 B.n106 163.367
R493 B.n407 B.n106 163.367
R494 B.n408 B.n407 163.367
R495 B.n409 B.n408 163.367
R496 B.n409 B.n104 163.367
R497 B.n413 B.n104 163.367
R498 B.n473 B.n84 163.367
R499 B.n469 B.n84 163.367
R500 B.n469 B.n468 163.367
R501 B.n468 B.n467 163.367
R502 B.n467 B.n86 163.367
R503 B.n463 B.n86 163.367
R504 B.n463 B.n462 163.367
R505 B.n462 B.n461 163.367
R506 B.n461 B.n88 163.367
R507 B.n457 B.n88 163.367
R508 B.n457 B.n456 163.367
R509 B.n456 B.n455 163.367
R510 B.n455 B.n90 163.367
R511 B.n451 B.n90 163.367
R512 B.n451 B.n450 163.367
R513 B.n450 B.n449 163.367
R514 B.n449 B.n92 163.367
R515 B.n445 B.n92 163.367
R516 B.n445 B.n444 163.367
R517 B.n444 B.n443 163.367
R518 B.n443 B.n94 163.367
R519 B.n439 B.n94 163.367
R520 B.n439 B.n438 163.367
R521 B.n438 B.n437 163.367
R522 B.n437 B.n96 163.367
R523 B.n433 B.n96 163.367
R524 B.n433 B.n432 163.367
R525 B.n432 B.n431 163.367
R526 B.n431 B.n98 163.367
R527 B.n427 B.n98 163.367
R528 B.n427 B.n426 163.367
R529 B.n426 B.n425 163.367
R530 B.n425 B.n100 163.367
R531 B.n421 B.n100 163.367
R532 B.n421 B.n420 163.367
R533 B.n420 B.n419 163.367
R534 B.n419 B.n102 163.367
R535 B.n415 B.n102 163.367
R536 B.n415 B.n414 163.367
R537 B.n674 B.n673 163.367
R538 B.n673 B.n672 163.367
R539 B.n672 B.n13 163.367
R540 B.n668 B.n13 163.367
R541 B.n668 B.n667 163.367
R542 B.n667 B.n666 163.367
R543 B.n666 B.n15 163.367
R544 B.n662 B.n15 163.367
R545 B.n662 B.n661 163.367
R546 B.n661 B.n660 163.367
R547 B.n660 B.n17 163.367
R548 B.n656 B.n17 163.367
R549 B.n656 B.n655 163.367
R550 B.n655 B.n654 163.367
R551 B.n654 B.n19 163.367
R552 B.n650 B.n19 163.367
R553 B.n650 B.n649 163.367
R554 B.n649 B.n648 163.367
R555 B.n648 B.n21 163.367
R556 B.n644 B.n21 163.367
R557 B.n644 B.n643 163.367
R558 B.n643 B.n642 163.367
R559 B.n642 B.n23 163.367
R560 B.n638 B.n23 163.367
R561 B.n638 B.n637 163.367
R562 B.n637 B.n636 163.367
R563 B.n636 B.n25 163.367
R564 B.n632 B.n25 163.367
R565 B.n632 B.n631 163.367
R566 B.n631 B.n630 163.367
R567 B.n630 B.n27 163.367
R568 B.n626 B.n27 163.367
R569 B.n626 B.n625 163.367
R570 B.n625 B.n624 163.367
R571 B.n624 B.n29 163.367
R572 B.n620 B.n29 163.367
R573 B.n620 B.n619 163.367
R574 B.n619 B.n618 163.367
R575 B.n618 B.n31 163.367
R576 B.n614 B.n31 163.367
R577 B.n614 B.n613 163.367
R578 B.n613 B.n612 163.367
R579 B.n612 B.n33 163.367
R580 B.n608 B.n33 163.367
R581 B.n608 B.n607 163.367
R582 B.n607 B.n606 163.367
R583 B.n606 B.n35 163.367
R584 B.n602 B.n35 163.367
R585 B.n602 B.n601 163.367
R586 B.n601 B.n600 163.367
R587 B.n600 B.n37 163.367
R588 B.n596 B.n37 163.367
R589 B.n596 B.n595 163.367
R590 B.n595 B.n594 163.367
R591 B.n594 B.n39 163.367
R592 B.n590 B.n39 163.367
R593 B.n590 B.n589 163.367
R594 B.n589 B.n588 163.367
R595 B.n588 B.n41 163.367
R596 B.n584 B.n41 163.367
R597 B.n584 B.n583 163.367
R598 B.n583 B.n582 163.367
R599 B.n582 B.n43 163.367
R600 B.n578 B.n43 163.367
R601 B.n578 B.n577 163.367
R602 B.n577 B.n576 163.367
R603 B.n576 B.n48 163.367
R604 B.n572 B.n48 163.367
R605 B.n572 B.n571 163.367
R606 B.n571 B.n570 163.367
R607 B.n570 B.n50 163.367
R608 B.n565 B.n50 163.367
R609 B.n565 B.n564 163.367
R610 B.n564 B.n563 163.367
R611 B.n563 B.n54 163.367
R612 B.n559 B.n54 163.367
R613 B.n559 B.n558 163.367
R614 B.n558 B.n557 163.367
R615 B.n557 B.n56 163.367
R616 B.n553 B.n56 163.367
R617 B.n553 B.n552 163.367
R618 B.n552 B.n551 163.367
R619 B.n551 B.n58 163.367
R620 B.n547 B.n58 163.367
R621 B.n547 B.n546 163.367
R622 B.n546 B.n545 163.367
R623 B.n545 B.n60 163.367
R624 B.n541 B.n60 163.367
R625 B.n541 B.n540 163.367
R626 B.n540 B.n539 163.367
R627 B.n539 B.n62 163.367
R628 B.n535 B.n62 163.367
R629 B.n535 B.n534 163.367
R630 B.n534 B.n533 163.367
R631 B.n533 B.n64 163.367
R632 B.n529 B.n64 163.367
R633 B.n529 B.n528 163.367
R634 B.n528 B.n527 163.367
R635 B.n527 B.n66 163.367
R636 B.n523 B.n66 163.367
R637 B.n523 B.n522 163.367
R638 B.n522 B.n521 163.367
R639 B.n521 B.n68 163.367
R640 B.n517 B.n68 163.367
R641 B.n517 B.n516 163.367
R642 B.n516 B.n515 163.367
R643 B.n515 B.n70 163.367
R644 B.n511 B.n70 163.367
R645 B.n511 B.n510 163.367
R646 B.n510 B.n509 163.367
R647 B.n509 B.n72 163.367
R648 B.n505 B.n72 163.367
R649 B.n505 B.n504 163.367
R650 B.n504 B.n503 163.367
R651 B.n503 B.n74 163.367
R652 B.n499 B.n74 163.367
R653 B.n499 B.n498 163.367
R654 B.n498 B.n497 163.367
R655 B.n497 B.n76 163.367
R656 B.n493 B.n76 163.367
R657 B.n493 B.n492 163.367
R658 B.n492 B.n491 163.367
R659 B.n491 B.n78 163.367
R660 B.n487 B.n78 163.367
R661 B.n487 B.n486 163.367
R662 B.n486 B.n485 163.367
R663 B.n485 B.n80 163.367
R664 B.n481 B.n80 163.367
R665 B.n481 B.n480 163.367
R666 B.n480 B.n479 163.367
R667 B.n479 B.n82 163.367
R668 B.n475 B.n82 163.367
R669 B.n475 B.n474 163.367
R670 B.n678 B.n11 163.367
R671 B.n679 B.n678 163.367
R672 B.n680 B.n679 163.367
R673 B.n680 B.n9 163.367
R674 B.n684 B.n9 163.367
R675 B.n685 B.n684 163.367
R676 B.n686 B.n685 163.367
R677 B.n686 B.n7 163.367
R678 B.n690 B.n7 163.367
R679 B.n691 B.n690 163.367
R680 B.n692 B.n691 163.367
R681 B.n692 B.n5 163.367
R682 B.n696 B.n5 163.367
R683 B.n697 B.n696 163.367
R684 B.n698 B.n697 163.367
R685 B.n698 B.n3 163.367
R686 B.n702 B.n3 163.367
R687 B.n703 B.n702 163.367
R688 B.n182 B.n2 163.367
R689 B.n183 B.n182 163.367
R690 B.n183 B.n180 163.367
R691 B.n187 B.n180 163.367
R692 B.n188 B.n187 163.367
R693 B.n189 B.n188 163.367
R694 B.n189 B.n178 163.367
R695 B.n193 B.n178 163.367
R696 B.n194 B.n193 163.367
R697 B.n195 B.n194 163.367
R698 B.n195 B.n176 163.367
R699 B.n199 B.n176 163.367
R700 B.n200 B.n199 163.367
R701 B.n201 B.n200 163.367
R702 B.n201 B.n174 163.367
R703 B.n205 B.n174 163.367
R704 B.n206 B.n205 163.367
R705 B.n207 B.n206 163.367
R706 B.n302 B.n301 59.5399
R707 B.n320 B.n136 59.5399
R708 B.n567 B.n52 59.5399
R709 B.n46 B.n45 59.5399
R710 B.n676 B.n675 28.8785
R711 B.n472 B.n83 28.8785
R712 B.n209 B.n208 28.8785
R713 B.n412 B.n103 28.8785
R714 B.n301 B.n300 24.6308
R715 B.n136 B.n135 24.6308
R716 B.n52 B.n51 24.6308
R717 B.n45 B.n44 24.6308
R718 B B.n705 18.0485
R719 B.n677 B.n676 10.6151
R720 B.n677 B.n10 10.6151
R721 B.n681 B.n10 10.6151
R722 B.n682 B.n681 10.6151
R723 B.n683 B.n682 10.6151
R724 B.n683 B.n8 10.6151
R725 B.n687 B.n8 10.6151
R726 B.n688 B.n687 10.6151
R727 B.n689 B.n688 10.6151
R728 B.n689 B.n6 10.6151
R729 B.n693 B.n6 10.6151
R730 B.n694 B.n693 10.6151
R731 B.n695 B.n694 10.6151
R732 B.n695 B.n4 10.6151
R733 B.n699 B.n4 10.6151
R734 B.n700 B.n699 10.6151
R735 B.n701 B.n700 10.6151
R736 B.n701 B.n0 10.6151
R737 B.n675 B.n12 10.6151
R738 B.n671 B.n12 10.6151
R739 B.n671 B.n670 10.6151
R740 B.n670 B.n669 10.6151
R741 B.n669 B.n14 10.6151
R742 B.n665 B.n14 10.6151
R743 B.n665 B.n664 10.6151
R744 B.n664 B.n663 10.6151
R745 B.n663 B.n16 10.6151
R746 B.n659 B.n16 10.6151
R747 B.n659 B.n658 10.6151
R748 B.n658 B.n657 10.6151
R749 B.n657 B.n18 10.6151
R750 B.n653 B.n18 10.6151
R751 B.n653 B.n652 10.6151
R752 B.n652 B.n651 10.6151
R753 B.n651 B.n20 10.6151
R754 B.n647 B.n20 10.6151
R755 B.n647 B.n646 10.6151
R756 B.n646 B.n645 10.6151
R757 B.n645 B.n22 10.6151
R758 B.n641 B.n22 10.6151
R759 B.n641 B.n640 10.6151
R760 B.n640 B.n639 10.6151
R761 B.n639 B.n24 10.6151
R762 B.n635 B.n24 10.6151
R763 B.n635 B.n634 10.6151
R764 B.n634 B.n633 10.6151
R765 B.n633 B.n26 10.6151
R766 B.n629 B.n26 10.6151
R767 B.n629 B.n628 10.6151
R768 B.n628 B.n627 10.6151
R769 B.n627 B.n28 10.6151
R770 B.n623 B.n28 10.6151
R771 B.n623 B.n622 10.6151
R772 B.n622 B.n621 10.6151
R773 B.n621 B.n30 10.6151
R774 B.n617 B.n30 10.6151
R775 B.n617 B.n616 10.6151
R776 B.n616 B.n615 10.6151
R777 B.n615 B.n32 10.6151
R778 B.n611 B.n32 10.6151
R779 B.n611 B.n610 10.6151
R780 B.n610 B.n609 10.6151
R781 B.n609 B.n34 10.6151
R782 B.n605 B.n34 10.6151
R783 B.n605 B.n604 10.6151
R784 B.n604 B.n603 10.6151
R785 B.n603 B.n36 10.6151
R786 B.n599 B.n36 10.6151
R787 B.n599 B.n598 10.6151
R788 B.n598 B.n597 10.6151
R789 B.n597 B.n38 10.6151
R790 B.n593 B.n38 10.6151
R791 B.n593 B.n592 10.6151
R792 B.n592 B.n591 10.6151
R793 B.n591 B.n40 10.6151
R794 B.n587 B.n40 10.6151
R795 B.n587 B.n586 10.6151
R796 B.n586 B.n585 10.6151
R797 B.n585 B.n42 10.6151
R798 B.n581 B.n580 10.6151
R799 B.n580 B.n579 10.6151
R800 B.n579 B.n47 10.6151
R801 B.n575 B.n47 10.6151
R802 B.n575 B.n574 10.6151
R803 B.n574 B.n573 10.6151
R804 B.n573 B.n49 10.6151
R805 B.n569 B.n49 10.6151
R806 B.n569 B.n568 10.6151
R807 B.n566 B.n53 10.6151
R808 B.n562 B.n53 10.6151
R809 B.n562 B.n561 10.6151
R810 B.n561 B.n560 10.6151
R811 B.n560 B.n55 10.6151
R812 B.n556 B.n55 10.6151
R813 B.n556 B.n555 10.6151
R814 B.n555 B.n554 10.6151
R815 B.n554 B.n57 10.6151
R816 B.n550 B.n57 10.6151
R817 B.n550 B.n549 10.6151
R818 B.n549 B.n548 10.6151
R819 B.n548 B.n59 10.6151
R820 B.n544 B.n59 10.6151
R821 B.n544 B.n543 10.6151
R822 B.n543 B.n542 10.6151
R823 B.n542 B.n61 10.6151
R824 B.n538 B.n61 10.6151
R825 B.n538 B.n537 10.6151
R826 B.n537 B.n536 10.6151
R827 B.n536 B.n63 10.6151
R828 B.n532 B.n63 10.6151
R829 B.n532 B.n531 10.6151
R830 B.n531 B.n530 10.6151
R831 B.n530 B.n65 10.6151
R832 B.n526 B.n65 10.6151
R833 B.n526 B.n525 10.6151
R834 B.n525 B.n524 10.6151
R835 B.n524 B.n67 10.6151
R836 B.n520 B.n67 10.6151
R837 B.n520 B.n519 10.6151
R838 B.n519 B.n518 10.6151
R839 B.n518 B.n69 10.6151
R840 B.n514 B.n69 10.6151
R841 B.n514 B.n513 10.6151
R842 B.n513 B.n512 10.6151
R843 B.n512 B.n71 10.6151
R844 B.n508 B.n71 10.6151
R845 B.n508 B.n507 10.6151
R846 B.n507 B.n506 10.6151
R847 B.n506 B.n73 10.6151
R848 B.n502 B.n73 10.6151
R849 B.n502 B.n501 10.6151
R850 B.n501 B.n500 10.6151
R851 B.n500 B.n75 10.6151
R852 B.n496 B.n75 10.6151
R853 B.n496 B.n495 10.6151
R854 B.n495 B.n494 10.6151
R855 B.n494 B.n77 10.6151
R856 B.n490 B.n77 10.6151
R857 B.n490 B.n489 10.6151
R858 B.n489 B.n488 10.6151
R859 B.n488 B.n79 10.6151
R860 B.n484 B.n79 10.6151
R861 B.n484 B.n483 10.6151
R862 B.n483 B.n482 10.6151
R863 B.n482 B.n81 10.6151
R864 B.n478 B.n81 10.6151
R865 B.n478 B.n477 10.6151
R866 B.n477 B.n476 10.6151
R867 B.n476 B.n83 10.6151
R868 B.n472 B.n471 10.6151
R869 B.n471 B.n470 10.6151
R870 B.n470 B.n85 10.6151
R871 B.n466 B.n85 10.6151
R872 B.n466 B.n465 10.6151
R873 B.n465 B.n464 10.6151
R874 B.n464 B.n87 10.6151
R875 B.n460 B.n87 10.6151
R876 B.n460 B.n459 10.6151
R877 B.n459 B.n458 10.6151
R878 B.n458 B.n89 10.6151
R879 B.n454 B.n89 10.6151
R880 B.n454 B.n453 10.6151
R881 B.n453 B.n452 10.6151
R882 B.n452 B.n91 10.6151
R883 B.n448 B.n91 10.6151
R884 B.n448 B.n447 10.6151
R885 B.n447 B.n446 10.6151
R886 B.n446 B.n93 10.6151
R887 B.n442 B.n93 10.6151
R888 B.n442 B.n441 10.6151
R889 B.n441 B.n440 10.6151
R890 B.n440 B.n95 10.6151
R891 B.n436 B.n95 10.6151
R892 B.n436 B.n435 10.6151
R893 B.n435 B.n434 10.6151
R894 B.n434 B.n97 10.6151
R895 B.n430 B.n97 10.6151
R896 B.n430 B.n429 10.6151
R897 B.n429 B.n428 10.6151
R898 B.n428 B.n99 10.6151
R899 B.n424 B.n99 10.6151
R900 B.n424 B.n423 10.6151
R901 B.n423 B.n422 10.6151
R902 B.n422 B.n101 10.6151
R903 B.n418 B.n101 10.6151
R904 B.n418 B.n417 10.6151
R905 B.n417 B.n416 10.6151
R906 B.n416 B.n103 10.6151
R907 B.n181 B.n1 10.6151
R908 B.n184 B.n181 10.6151
R909 B.n185 B.n184 10.6151
R910 B.n186 B.n185 10.6151
R911 B.n186 B.n179 10.6151
R912 B.n190 B.n179 10.6151
R913 B.n191 B.n190 10.6151
R914 B.n192 B.n191 10.6151
R915 B.n192 B.n177 10.6151
R916 B.n196 B.n177 10.6151
R917 B.n197 B.n196 10.6151
R918 B.n198 B.n197 10.6151
R919 B.n198 B.n175 10.6151
R920 B.n202 B.n175 10.6151
R921 B.n203 B.n202 10.6151
R922 B.n204 B.n203 10.6151
R923 B.n204 B.n173 10.6151
R924 B.n208 B.n173 10.6151
R925 B.n210 B.n209 10.6151
R926 B.n210 B.n171 10.6151
R927 B.n214 B.n171 10.6151
R928 B.n215 B.n214 10.6151
R929 B.n216 B.n215 10.6151
R930 B.n216 B.n169 10.6151
R931 B.n220 B.n169 10.6151
R932 B.n221 B.n220 10.6151
R933 B.n222 B.n221 10.6151
R934 B.n222 B.n167 10.6151
R935 B.n226 B.n167 10.6151
R936 B.n227 B.n226 10.6151
R937 B.n228 B.n227 10.6151
R938 B.n228 B.n165 10.6151
R939 B.n232 B.n165 10.6151
R940 B.n233 B.n232 10.6151
R941 B.n234 B.n233 10.6151
R942 B.n234 B.n163 10.6151
R943 B.n238 B.n163 10.6151
R944 B.n239 B.n238 10.6151
R945 B.n240 B.n239 10.6151
R946 B.n240 B.n161 10.6151
R947 B.n244 B.n161 10.6151
R948 B.n245 B.n244 10.6151
R949 B.n246 B.n245 10.6151
R950 B.n246 B.n159 10.6151
R951 B.n250 B.n159 10.6151
R952 B.n251 B.n250 10.6151
R953 B.n252 B.n251 10.6151
R954 B.n252 B.n157 10.6151
R955 B.n256 B.n157 10.6151
R956 B.n257 B.n256 10.6151
R957 B.n258 B.n257 10.6151
R958 B.n258 B.n155 10.6151
R959 B.n262 B.n155 10.6151
R960 B.n263 B.n262 10.6151
R961 B.n264 B.n263 10.6151
R962 B.n264 B.n153 10.6151
R963 B.n268 B.n153 10.6151
R964 B.n269 B.n268 10.6151
R965 B.n270 B.n269 10.6151
R966 B.n270 B.n151 10.6151
R967 B.n274 B.n151 10.6151
R968 B.n275 B.n274 10.6151
R969 B.n276 B.n275 10.6151
R970 B.n276 B.n149 10.6151
R971 B.n280 B.n149 10.6151
R972 B.n281 B.n280 10.6151
R973 B.n282 B.n281 10.6151
R974 B.n282 B.n147 10.6151
R975 B.n286 B.n147 10.6151
R976 B.n287 B.n286 10.6151
R977 B.n288 B.n287 10.6151
R978 B.n288 B.n145 10.6151
R979 B.n292 B.n145 10.6151
R980 B.n293 B.n292 10.6151
R981 B.n294 B.n293 10.6151
R982 B.n294 B.n143 10.6151
R983 B.n298 B.n143 10.6151
R984 B.n299 B.n298 10.6151
R985 B.n303 B.n299 10.6151
R986 B.n307 B.n141 10.6151
R987 B.n308 B.n307 10.6151
R988 B.n309 B.n308 10.6151
R989 B.n309 B.n139 10.6151
R990 B.n313 B.n139 10.6151
R991 B.n314 B.n313 10.6151
R992 B.n315 B.n314 10.6151
R993 B.n315 B.n137 10.6151
R994 B.n319 B.n137 10.6151
R995 B.n322 B.n321 10.6151
R996 B.n322 B.n133 10.6151
R997 B.n326 B.n133 10.6151
R998 B.n327 B.n326 10.6151
R999 B.n328 B.n327 10.6151
R1000 B.n328 B.n131 10.6151
R1001 B.n332 B.n131 10.6151
R1002 B.n333 B.n332 10.6151
R1003 B.n334 B.n333 10.6151
R1004 B.n334 B.n129 10.6151
R1005 B.n338 B.n129 10.6151
R1006 B.n339 B.n338 10.6151
R1007 B.n340 B.n339 10.6151
R1008 B.n340 B.n127 10.6151
R1009 B.n344 B.n127 10.6151
R1010 B.n345 B.n344 10.6151
R1011 B.n346 B.n345 10.6151
R1012 B.n346 B.n125 10.6151
R1013 B.n350 B.n125 10.6151
R1014 B.n351 B.n350 10.6151
R1015 B.n352 B.n351 10.6151
R1016 B.n352 B.n123 10.6151
R1017 B.n356 B.n123 10.6151
R1018 B.n357 B.n356 10.6151
R1019 B.n358 B.n357 10.6151
R1020 B.n358 B.n121 10.6151
R1021 B.n362 B.n121 10.6151
R1022 B.n363 B.n362 10.6151
R1023 B.n364 B.n363 10.6151
R1024 B.n364 B.n119 10.6151
R1025 B.n368 B.n119 10.6151
R1026 B.n369 B.n368 10.6151
R1027 B.n370 B.n369 10.6151
R1028 B.n370 B.n117 10.6151
R1029 B.n374 B.n117 10.6151
R1030 B.n375 B.n374 10.6151
R1031 B.n376 B.n375 10.6151
R1032 B.n376 B.n115 10.6151
R1033 B.n380 B.n115 10.6151
R1034 B.n381 B.n380 10.6151
R1035 B.n382 B.n381 10.6151
R1036 B.n382 B.n113 10.6151
R1037 B.n386 B.n113 10.6151
R1038 B.n387 B.n386 10.6151
R1039 B.n388 B.n387 10.6151
R1040 B.n388 B.n111 10.6151
R1041 B.n392 B.n111 10.6151
R1042 B.n393 B.n392 10.6151
R1043 B.n394 B.n393 10.6151
R1044 B.n394 B.n109 10.6151
R1045 B.n398 B.n109 10.6151
R1046 B.n399 B.n398 10.6151
R1047 B.n400 B.n399 10.6151
R1048 B.n400 B.n107 10.6151
R1049 B.n404 B.n107 10.6151
R1050 B.n405 B.n404 10.6151
R1051 B.n406 B.n405 10.6151
R1052 B.n406 B.n105 10.6151
R1053 B.n410 B.n105 10.6151
R1054 B.n411 B.n410 10.6151
R1055 B.n412 B.n411 10.6151
R1056 B.n46 B.n42 9.36635
R1057 B.n567 B.n566 9.36635
R1058 B.n303 B.n302 9.36635
R1059 B.n321 B.n320 9.36635
R1060 B.n705 B.n0 8.11757
R1061 B.n705 B.n1 8.11757
R1062 B.n581 B.n46 1.24928
R1063 B.n568 B.n567 1.24928
R1064 B.n302 B.n141 1.24928
R1065 B.n320 B.n319 1.24928
R1066 VN.n0 VN.t3 546.5
R1067 VN.n1 VN.t2 546.5
R1068 VN.n1 VN.t1 546.413
R1069 VN.n0 VN.t0 546.413
R1070 VN VN.n1 77.9857
R1071 VN VN.n0 31.2622
R1072 VTAIL.n842 VTAIL.n742 756.745
R1073 VTAIL.n100 VTAIL.n0 756.745
R1074 VTAIL.n206 VTAIL.n106 756.745
R1075 VTAIL.n312 VTAIL.n212 756.745
R1076 VTAIL.n736 VTAIL.n636 756.745
R1077 VTAIL.n630 VTAIL.n530 756.745
R1078 VTAIL.n524 VTAIL.n424 756.745
R1079 VTAIL.n418 VTAIL.n318 756.745
R1080 VTAIL.n777 VTAIL.n776 585
R1081 VTAIL.n774 VTAIL.n773 585
R1082 VTAIL.n783 VTAIL.n782 585
R1083 VTAIL.n785 VTAIL.n784 585
R1084 VTAIL.n770 VTAIL.n769 585
R1085 VTAIL.n791 VTAIL.n790 585
R1086 VTAIL.n793 VTAIL.n792 585
R1087 VTAIL.n766 VTAIL.n765 585
R1088 VTAIL.n799 VTAIL.n798 585
R1089 VTAIL.n801 VTAIL.n800 585
R1090 VTAIL.n762 VTAIL.n761 585
R1091 VTAIL.n807 VTAIL.n806 585
R1092 VTAIL.n809 VTAIL.n808 585
R1093 VTAIL.n758 VTAIL.n757 585
R1094 VTAIL.n815 VTAIL.n814 585
R1095 VTAIL.n818 VTAIL.n817 585
R1096 VTAIL.n816 VTAIL.n754 585
R1097 VTAIL.n823 VTAIL.n753 585
R1098 VTAIL.n825 VTAIL.n824 585
R1099 VTAIL.n827 VTAIL.n826 585
R1100 VTAIL.n750 VTAIL.n749 585
R1101 VTAIL.n833 VTAIL.n832 585
R1102 VTAIL.n835 VTAIL.n834 585
R1103 VTAIL.n746 VTAIL.n745 585
R1104 VTAIL.n841 VTAIL.n840 585
R1105 VTAIL.n843 VTAIL.n842 585
R1106 VTAIL.n35 VTAIL.n34 585
R1107 VTAIL.n32 VTAIL.n31 585
R1108 VTAIL.n41 VTAIL.n40 585
R1109 VTAIL.n43 VTAIL.n42 585
R1110 VTAIL.n28 VTAIL.n27 585
R1111 VTAIL.n49 VTAIL.n48 585
R1112 VTAIL.n51 VTAIL.n50 585
R1113 VTAIL.n24 VTAIL.n23 585
R1114 VTAIL.n57 VTAIL.n56 585
R1115 VTAIL.n59 VTAIL.n58 585
R1116 VTAIL.n20 VTAIL.n19 585
R1117 VTAIL.n65 VTAIL.n64 585
R1118 VTAIL.n67 VTAIL.n66 585
R1119 VTAIL.n16 VTAIL.n15 585
R1120 VTAIL.n73 VTAIL.n72 585
R1121 VTAIL.n76 VTAIL.n75 585
R1122 VTAIL.n74 VTAIL.n12 585
R1123 VTAIL.n81 VTAIL.n11 585
R1124 VTAIL.n83 VTAIL.n82 585
R1125 VTAIL.n85 VTAIL.n84 585
R1126 VTAIL.n8 VTAIL.n7 585
R1127 VTAIL.n91 VTAIL.n90 585
R1128 VTAIL.n93 VTAIL.n92 585
R1129 VTAIL.n4 VTAIL.n3 585
R1130 VTAIL.n99 VTAIL.n98 585
R1131 VTAIL.n101 VTAIL.n100 585
R1132 VTAIL.n141 VTAIL.n140 585
R1133 VTAIL.n138 VTAIL.n137 585
R1134 VTAIL.n147 VTAIL.n146 585
R1135 VTAIL.n149 VTAIL.n148 585
R1136 VTAIL.n134 VTAIL.n133 585
R1137 VTAIL.n155 VTAIL.n154 585
R1138 VTAIL.n157 VTAIL.n156 585
R1139 VTAIL.n130 VTAIL.n129 585
R1140 VTAIL.n163 VTAIL.n162 585
R1141 VTAIL.n165 VTAIL.n164 585
R1142 VTAIL.n126 VTAIL.n125 585
R1143 VTAIL.n171 VTAIL.n170 585
R1144 VTAIL.n173 VTAIL.n172 585
R1145 VTAIL.n122 VTAIL.n121 585
R1146 VTAIL.n179 VTAIL.n178 585
R1147 VTAIL.n182 VTAIL.n181 585
R1148 VTAIL.n180 VTAIL.n118 585
R1149 VTAIL.n187 VTAIL.n117 585
R1150 VTAIL.n189 VTAIL.n188 585
R1151 VTAIL.n191 VTAIL.n190 585
R1152 VTAIL.n114 VTAIL.n113 585
R1153 VTAIL.n197 VTAIL.n196 585
R1154 VTAIL.n199 VTAIL.n198 585
R1155 VTAIL.n110 VTAIL.n109 585
R1156 VTAIL.n205 VTAIL.n204 585
R1157 VTAIL.n207 VTAIL.n206 585
R1158 VTAIL.n247 VTAIL.n246 585
R1159 VTAIL.n244 VTAIL.n243 585
R1160 VTAIL.n253 VTAIL.n252 585
R1161 VTAIL.n255 VTAIL.n254 585
R1162 VTAIL.n240 VTAIL.n239 585
R1163 VTAIL.n261 VTAIL.n260 585
R1164 VTAIL.n263 VTAIL.n262 585
R1165 VTAIL.n236 VTAIL.n235 585
R1166 VTAIL.n269 VTAIL.n268 585
R1167 VTAIL.n271 VTAIL.n270 585
R1168 VTAIL.n232 VTAIL.n231 585
R1169 VTAIL.n277 VTAIL.n276 585
R1170 VTAIL.n279 VTAIL.n278 585
R1171 VTAIL.n228 VTAIL.n227 585
R1172 VTAIL.n285 VTAIL.n284 585
R1173 VTAIL.n288 VTAIL.n287 585
R1174 VTAIL.n286 VTAIL.n224 585
R1175 VTAIL.n293 VTAIL.n223 585
R1176 VTAIL.n295 VTAIL.n294 585
R1177 VTAIL.n297 VTAIL.n296 585
R1178 VTAIL.n220 VTAIL.n219 585
R1179 VTAIL.n303 VTAIL.n302 585
R1180 VTAIL.n305 VTAIL.n304 585
R1181 VTAIL.n216 VTAIL.n215 585
R1182 VTAIL.n311 VTAIL.n310 585
R1183 VTAIL.n313 VTAIL.n312 585
R1184 VTAIL.n737 VTAIL.n736 585
R1185 VTAIL.n735 VTAIL.n734 585
R1186 VTAIL.n640 VTAIL.n639 585
R1187 VTAIL.n729 VTAIL.n728 585
R1188 VTAIL.n727 VTAIL.n726 585
R1189 VTAIL.n644 VTAIL.n643 585
R1190 VTAIL.n721 VTAIL.n720 585
R1191 VTAIL.n719 VTAIL.n718 585
R1192 VTAIL.n717 VTAIL.n647 585
R1193 VTAIL.n651 VTAIL.n648 585
R1194 VTAIL.n712 VTAIL.n711 585
R1195 VTAIL.n710 VTAIL.n709 585
R1196 VTAIL.n653 VTAIL.n652 585
R1197 VTAIL.n704 VTAIL.n703 585
R1198 VTAIL.n702 VTAIL.n701 585
R1199 VTAIL.n657 VTAIL.n656 585
R1200 VTAIL.n696 VTAIL.n695 585
R1201 VTAIL.n694 VTAIL.n693 585
R1202 VTAIL.n661 VTAIL.n660 585
R1203 VTAIL.n688 VTAIL.n687 585
R1204 VTAIL.n686 VTAIL.n685 585
R1205 VTAIL.n665 VTAIL.n664 585
R1206 VTAIL.n680 VTAIL.n679 585
R1207 VTAIL.n678 VTAIL.n677 585
R1208 VTAIL.n669 VTAIL.n668 585
R1209 VTAIL.n672 VTAIL.n671 585
R1210 VTAIL.n631 VTAIL.n630 585
R1211 VTAIL.n629 VTAIL.n628 585
R1212 VTAIL.n534 VTAIL.n533 585
R1213 VTAIL.n623 VTAIL.n622 585
R1214 VTAIL.n621 VTAIL.n620 585
R1215 VTAIL.n538 VTAIL.n537 585
R1216 VTAIL.n615 VTAIL.n614 585
R1217 VTAIL.n613 VTAIL.n612 585
R1218 VTAIL.n611 VTAIL.n541 585
R1219 VTAIL.n545 VTAIL.n542 585
R1220 VTAIL.n606 VTAIL.n605 585
R1221 VTAIL.n604 VTAIL.n603 585
R1222 VTAIL.n547 VTAIL.n546 585
R1223 VTAIL.n598 VTAIL.n597 585
R1224 VTAIL.n596 VTAIL.n595 585
R1225 VTAIL.n551 VTAIL.n550 585
R1226 VTAIL.n590 VTAIL.n589 585
R1227 VTAIL.n588 VTAIL.n587 585
R1228 VTAIL.n555 VTAIL.n554 585
R1229 VTAIL.n582 VTAIL.n581 585
R1230 VTAIL.n580 VTAIL.n579 585
R1231 VTAIL.n559 VTAIL.n558 585
R1232 VTAIL.n574 VTAIL.n573 585
R1233 VTAIL.n572 VTAIL.n571 585
R1234 VTAIL.n563 VTAIL.n562 585
R1235 VTAIL.n566 VTAIL.n565 585
R1236 VTAIL.n525 VTAIL.n524 585
R1237 VTAIL.n523 VTAIL.n522 585
R1238 VTAIL.n428 VTAIL.n427 585
R1239 VTAIL.n517 VTAIL.n516 585
R1240 VTAIL.n515 VTAIL.n514 585
R1241 VTAIL.n432 VTAIL.n431 585
R1242 VTAIL.n509 VTAIL.n508 585
R1243 VTAIL.n507 VTAIL.n506 585
R1244 VTAIL.n505 VTAIL.n435 585
R1245 VTAIL.n439 VTAIL.n436 585
R1246 VTAIL.n500 VTAIL.n499 585
R1247 VTAIL.n498 VTAIL.n497 585
R1248 VTAIL.n441 VTAIL.n440 585
R1249 VTAIL.n492 VTAIL.n491 585
R1250 VTAIL.n490 VTAIL.n489 585
R1251 VTAIL.n445 VTAIL.n444 585
R1252 VTAIL.n484 VTAIL.n483 585
R1253 VTAIL.n482 VTAIL.n481 585
R1254 VTAIL.n449 VTAIL.n448 585
R1255 VTAIL.n476 VTAIL.n475 585
R1256 VTAIL.n474 VTAIL.n473 585
R1257 VTAIL.n453 VTAIL.n452 585
R1258 VTAIL.n468 VTAIL.n467 585
R1259 VTAIL.n466 VTAIL.n465 585
R1260 VTAIL.n457 VTAIL.n456 585
R1261 VTAIL.n460 VTAIL.n459 585
R1262 VTAIL.n419 VTAIL.n418 585
R1263 VTAIL.n417 VTAIL.n416 585
R1264 VTAIL.n322 VTAIL.n321 585
R1265 VTAIL.n411 VTAIL.n410 585
R1266 VTAIL.n409 VTAIL.n408 585
R1267 VTAIL.n326 VTAIL.n325 585
R1268 VTAIL.n403 VTAIL.n402 585
R1269 VTAIL.n401 VTAIL.n400 585
R1270 VTAIL.n399 VTAIL.n329 585
R1271 VTAIL.n333 VTAIL.n330 585
R1272 VTAIL.n394 VTAIL.n393 585
R1273 VTAIL.n392 VTAIL.n391 585
R1274 VTAIL.n335 VTAIL.n334 585
R1275 VTAIL.n386 VTAIL.n385 585
R1276 VTAIL.n384 VTAIL.n383 585
R1277 VTAIL.n339 VTAIL.n338 585
R1278 VTAIL.n378 VTAIL.n377 585
R1279 VTAIL.n376 VTAIL.n375 585
R1280 VTAIL.n343 VTAIL.n342 585
R1281 VTAIL.n370 VTAIL.n369 585
R1282 VTAIL.n368 VTAIL.n367 585
R1283 VTAIL.n347 VTAIL.n346 585
R1284 VTAIL.n362 VTAIL.n361 585
R1285 VTAIL.n360 VTAIL.n359 585
R1286 VTAIL.n351 VTAIL.n350 585
R1287 VTAIL.n354 VTAIL.n353 585
R1288 VTAIL.t2 VTAIL.n670 327.466
R1289 VTAIL.t0 VTAIL.n564 327.466
R1290 VTAIL.t7 VTAIL.n458 327.466
R1291 VTAIL.t4 VTAIL.n352 327.466
R1292 VTAIL.t6 VTAIL.n775 327.466
R1293 VTAIL.t5 VTAIL.n33 327.466
R1294 VTAIL.t3 VTAIL.n139 327.466
R1295 VTAIL.t1 VTAIL.n245 327.466
R1296 VTAIL.n776 VTAIL.n773 171.744
R1297 VTAIL.n783 VTAIL.n773 171.744
R1298 VTAIL.n784 VTAIL.n783 171.744
R1299 VTAIL.n784 VTAIL.n769 171.744
R1300 VTAIL.n791 VTAIL.n769 171.744
R1301 VTAIL.n792 VTAIL.n791 171.744
R1302 VTAIL.n792 VTAIL.n765 171.744
R1303 VTAIL.n799 VTAIL.n765 171.744
R1304 VTAIL.n800 VTAIL.n799 171.744
R1305 VTAIL.n800 VTAIL.n761 171.744
R1306 VTAIL.n807 VTAIL.n761 171.744
R1307 VTAIL.n808 VTAIL.n807 171.744
R1308 VTAIL.n808 VTAIL.n757 171.744
R1309 VTAIL.n815 VTAIL.n757 171.744
R1310 VTAIL.n817 VTAIL.n815 171.744
R1311 VTAIL.n817 VTAIL.n816 171.744
R1312 VTAIL.n816 VTAIL.n753 171.744
R1313 VTAIL.n825 VTAIL.n753 171.744
R1314 VTAIL.n826 VTAIL.n825 171.744
R1315 VTAIL.n826 VTAIL.n749 171.744
R1316 VTAIL.n833 VTAIL.n749 171.744
R1317 VTAIL.n834 VTAIL.n833 171.744
R1318 VTAIL.n834 VTAIL.n745 171.744
R1319 VTAIL.n841 VTAIL.n745 171.744
R1320 VTAIL.n842 VTAIL.n841 171.744
R1321 VTAIL.n34 VTAIL.n31 171.744
R1322 VTAIL.n41 VTAIL.n31 171.744
R1323 VTAIL.n42 VTAIL.n41 171.744
R1324 VTAIL.n42 VTAIL.n27 171.744
R1325 VTAIL.n49 VTAIL.n27 171.744
R1326 VTAIL.n50 VTAIL.n49 171.744
R1327 VTAIL.n50 VTAIL.n23 171.744
R1328 VTAIL.n57 VTAIL.n23 171.744
R1329 VTAIL.n58 VTAIL.n57 171.744
R1330 VTAIL.n58 VTAIL.n19 171.744
R1331 VTAIL.n65 VTAIL.n19 171.744
R1332 VTAIL.n66 VTAIL.n65 171.744
R1333 VTAIL.n66 VTAIL.n15 171.744
R1334 VTAIL.n73 VTAIL.n15 171.744
R1335 VTAIL.n75 VTAIL.n73 171.744
R1336 VTAIL.n75 VTAIL.n74 171.744
R1337 VTAIL.n74 VTAIL.n11 171.744
R1338 VTAIL.n83 VTAIL.n11 171.744
R1339 VTAIL.n84 VTAIL.n83 171.744
R1340 VTAIL.n84 VTAIL.n7 171.744
R1341 VTAIL.n91 VTAIL.n7 171.744
R1342 VTAIL.n92 VTAIL.n91 171.744
R1343 VTAIL.n92 VTAIL.n3 171.744
R1344 VTAIL.n99 VTAIL.n3 171.744
R1345 VTAIL.n100 VTAIL.n99 171.744
R1346 VTAIL.n140 VTAIL.n137 171.744
R1347 VTAIL.n147 VTAIL.n137 171.744
R1348 VTAIL.n148 VTAIL.n147 171.744
R1349 VTAIL.n148 VTAIL.n133 171.744
R1350 VTAIL.n155 VTAIL.n133 171.744
R1351 VTAIL.n156 VTAIL.n155 171.744
R1352 VTAIL.n156 VTAIL.n129 171.744
R1353 VTAIL.n163 VTAIL.n129 171.744
R1354 VTAIL.n164 VTAIL.n163 171.744
R1355 VTAIL.n164 VTAIL.n125 171.744
R1356 VTAIL.n171 VTAIL.n125 171.744
R1357 VTAIL.n172 VTAIL.n171 171.744
R1358 VTAIL.n172 VTAIL.n121 171.744
R1359 VTAIL.n179 VTAIL.n121 171.744
R1360 VTAIL.n181 VTAIL.n179 171.744
R1361 VTAIL.n181 VTAIL.n180 171.744
R1362 VTAIL.n180 VTAIL.n117 171.744
R1363 VTAIL.n189 VTAIL.n117 171.744
R1364 VTAIL.n190 VTAIL.n189 171.744
R1365 VTAIL.n190 VTAIL.n113 171.744
R1366 VTAIL.n197 VTAIL.n113 171.744
R1367 VTAIL.n198 VTAIL.n197 171.744
R1368 VTAIL.n198 VTAIL.n109 171.744
R1369 VTAIL.n205 VTAIL.n109 171.744
R1370 VTAIL.n206 VTAIL.n205 171.744
R1371 VTAIL.n246 VTAIL.n243 171.744
R1372 VTAIL.n253 VTAIL.n243 171.744
R1373 VTAIL.n254 VTAIL.n253 171.744
R1374 VTAIL.n254 VTAIL.n239 171.744
R1375 VTAIL.n261 VTAIL.n239 171.744
R1376 VTAIL.n262 VTAIL.n261 171.744
R1377 VTAIL.n262 VTAIL.n235 171.744
R1378 VTAIL.n269 VTAIL.n235 171.744
R1379 VTAIL.n270 VTAIL.n269 171.744
R1380 VTAIL.n270 VTAIL.n231 171.744
R1381 VTAIL.n277 VTAIL.n231 171.744
R1382 VTAIL.n278 VTAIL.n277 171.744
R1383 VTAIL.n278 VTAIL.n227 171.744
R1384 VTAIL.n285 VTAIL.n227 171.744
R1385 VTAIL.n287 VTAIL.n285 171.744
R1386 VTAIL.n287 VTAIL.n286 171.744
R1387 VTAIL.n286 VTAIL.n223 171.744
R1388 VTAIL.n295 VTAIL.n223 171.744
R1389 VTAIL.n296 VTAIL.n295 171.744
R1390 VTAIL.n296 VTAIL.n219 171.744
R1391 VTAIL.n303 VTAIL.n219 171.744
R1392 VTAIL.n304 VTAIL.n303 171.744
R1393 VTAIL.n304 VTAIL.n215 171.744
R1394 VTAIL.n311 VTAIL.n215 171.744
R1395 VTAIL.n312 VTAIL.n311 171.744
R1396 VTAIL.n736 VTAIL.n735 171.744
R1397 VTAIL.n735 VTAIL.n639 171.744
R1398 VTAIL.n728 VTAIL.n639 171.744
R1399 VTAIL.n728 VTAIL.n727 171.744
R1400 VTAIL.n727 VTAIL.n643 171.744
R1401 VTAIL.n720 VTAIL.n643 171.744
R1402 VTAIL.n720 VTAIL.n719 171.744
R1403 VTAIL.n719 VTAIL.n647 171.744
R1404 VTAIL.n651 VTAIL.n647 171.744
R1405 VTAIL.n711 VTAIL.n651 171.744
R1406 VTAIL.n711 VTAIL.n710 171.744
R1407 VTAIL.n710 VTAIL.n652 171.744
R1408 VTAIL.n703 VTAIL.n652 171.744
R1409 VTAIL.n703 VTAIL.n702 171.744
R1410 VTAIL.n702 VTAIL.n656 171.744
R1411 VTAIL.n695 VTAIL.n656 171.744
R1412 VTAIL.n695 VTAIL.n694 171.744
R1413 VTAIL.n694 VTAIL.n660 171.744
R1414 VTAIL.n687 VTAIL.n660 171.744
R1415 VTAIL.n687 VTAIL.n686 171.744
R1416 VTAIL.n686 VTAIL.n664 171.744
R1417 VTAIL.n679 VTAIL.n664 171.744
R1418 VTAIL.n679 VTAIL.n678 171.744
R1419 VTAIL.n678 VTAIL.n668 171.744
R1420 VTAIL.n671 VTAIL.n668 171.744
R1421 VTAIL.n630 VTAIL.n629 171.744
R1422 VTAIL.n629 VTAIL.n533 171.744
R1423 VTAIL.n622 VTAIL.n533 171.744
R1424 VTAIL.n622 VTAIL.n621 171.744
R1425 VTAIL.n621 VTAIL.n537 171.744
R1426 VTAIL.n614 VTAIL.n537 171.744
R1427 VTAIL.n614 VTAIL.n613 171.744
R1428 VTAIL.n613 VTAIL.n541 171.744
R1429 VTAIL.n545 VTAIL.n541 171.744
R1430 VTAIL.n605 VTAIL.n545 171.744
R1431 VTAIL.n605 VTAIL.n604 171.744
R1432 VTAIL.n604 VTAIL.n546 171.744
R1433 VTAIL.n597 VTAIL.n546 171.744
R1434 VTAIL.n597 VTAIL.n596 171.744
R1435 VTAIL.n596 VTAIL.n550 171.744
R1436 VTAIL.n589 VTAIL.n550 171.744
R1437 VTAIL.n589 VTAIL.n588 171.744
R1438 VTAIL.n588 VTAIL.n554 171.744
R1439 VTAIL.n581 VTAIL.n554 171.744
R1440 VTAIL.n581 VTAIL.n580 171.744
R1441 VTAIL.n580 VTAIL.n558 171.744
R1442 VTAIL.n573 VTAIL.n558 171.744
R1443 VTAIL.n573 VTAIL.n572 171.744
R1444 VTAIL.n572 VTAIL.n562 171.744
R1445 VTAIL.n565 VTAIL.n562 171.744
R1446 VTAIL.n524 VTAIL.n523 171.744
R1447 VTAIL.n523 VTAIL.n427 171.744
R1448 VTAIL.n516 VTAIL.n427 171.744
R1449 VTAIL.n516 VTAIL.n515 171.744
R1450 VTAIL.n515 VTAIL.n431 171.744
R1451 VTAIL.n508 VTAIL.n431 171.744
R1452 VTAIL.n508 VTAIL.n507 171.744
R1453 VTAIL.n507 VTAIL.n435 171.744
R1454 VTAIL.n439 VTAIL.n435 171.744
R1455 VTAIL.n499 VTAIL.n439 171.744
R1456 VTAIL.n499 VTAIL.n498 171.744
R1457 VTAIL.n498 VTAIL.n440 171.744
R1458 VTAIL.n491 VTAIL.n440 171.744
R1459 VTAIL.n491 VTAIL.n490 171.744
R1460 VTAIL.n490 VTAIL.n444 171.744
R1461 VTAIL.n483 VTAIL.n444 171.744
R1462 VTAIL.n483 VTAIL.n482 171.744
R1463 VTAIL.n482 VTAIL.n448 171.744
R1464 VTAIL.n475 VTAIL.n448 171.744
R1465 VTAIL.n475 VTAIL.n474 171.744
R1466 VTAIL.n474 VTAIL.n452 171.744
R1467 VTAIL.n467 VTAIL.n452 171.744
R1468 VTAIL.n467 VTAIL.n466 171.744
R1469 VTAIL.n466 VTAIL.n456 171.744
R1470 VTAIL.n459 VTAIL.n456 171.744
R1471 VTAIL.n418 VTAIL.n417 171.744
R1472 VTAIL.n417 VTAIL.n321 171.744
R1473 VTAIL.n410 VTAIL.n321 171.744
R1474 VTAIL.n410 VTAIL.n409 171.744
R1475 VTAIL.n409 VTAIL.n325 171.744
R1476 VTAIL.n402 VTAIL.n325 171.744
R1477 VTAIL.n402 VTAIL.n401 171.744
R1478 VTAIL.n401 VTAIL.n329 171.744
R1479 VTAIL.n333 VTAIL.n329 171.744
R1480 VTAIL.n393 VTAIL.n333 171.744
R1481 VTAIL.n393 VTAIL.n392 171.744
R1482 VTAIL.n392 VTAIL.n334 171.744
R1483 VTAIL.n385 VTAIL.n334 171.744
R1484 VTAIL.n385 VTAIL.n384 171.744
R1485 VTAIL.n384 VTAIL.n338 171.744
R1486 VTAIL.n377 VTAIL.n338 171.744
R1487 VTAIL.n377 VTAIL.n376 171.744
R1488 VTAIL.n376 VTAIL.n342 171.744
R1489 VTAIL.n369 VTAIL.n342 171.744
R1490 VTAIL.n369 VTAIL.n368 171.744
R1491 VTAIL.n368 VTAIL.n346 171.744
R1492 VTAIL.n361 VTAIL.n346 171.744
R1493 VTAIL.n361 VTAIL.n360 171.744
R1494 VTAIL.n360 VTAIL.n350 171.744
R1495 VTAIL.n353 VTAIL.n350 171.744
R1496 VTAIL.n776 VTAIL.t6 85.8723
R1497 VTAIL.n34 VTAIL.t5 85.8723
R1498 VTAIL.n140 VTAIL.t3 85.8723
R1499 VTAIL.n246 VTAIL.t1 85.8723
R1500 VTAIL.n671 VTAIL.t2 85.8723
R1501 VTAIL.n565 VTAIL.t0 85.8723
R1502 VTAIL.n459 VTAIL.t7 85.8723
R1503 VTAIL.n353 VTAIL.t4 85.8723
R1504 VTAIL.n847 VTAIL.n846 31.9914
R1505 VTAIL.n105 VTAIL.n104 31.9914
R1506 VTAIL.n211 VTAIL.n210 31.9914
R1507 VTAIL.n317 VTAIL.n316 31.9914
R1508 VTAIL.n741 VTAIL.n740 31.9914
R1509 VTAIL.n635 VTAIL.n634 31.9914
R1510 VTAIL.n529 VTAIL.n528 31.9914
R1511 VTAIL.n423 VTAIL.n422 31.9914
R1512 VTAIL.n847 VTAIL.n741 29.7979
R1513 VTAIL.n423 VTAIL.n317 29.7979
R1514 VTAIL.n777 VTAIL.n775 16.3895
R1515 VTAIL.n35 VTAIL.n33 16.3895
R1516 VTAIL.n141 VTAIL.n139 16.3895
R1517 VTAIL.n247 VTAIL.n245 16.3895
R1518 VTAIL.n672 VTAIL.n670 16.3895
R1519 VTAIL.n566 VTAIL.n564 16.3895
R1520 VTAIL.n460 VTAIL.n458 16.3895
R1521 VTAIL.n354 VTAIL.n352 16.3895
R1522 VTAIL.n824 VTAIL.n823 13.1884
R1523 VTAIL.n82 VTAIL.n81 13.1884
R1524 VTAIL.n188 VTAIL.n187 13.1884
R1525 VTAIL.n294 VTAIL.n293 13.1884
R1526 VTAIL.n718 VTAIL.n717 13.1884
R1527 VTAIL.n612 VTAIL.n611 13.1884
R1528 VTAIL.n506 VTAIL.n505 13.1884
R1529 VTAIL.n400 VTAIL.n399 13.1884
R1530 VTAIL.n778 VTAIL.n774 12.8005
R1531 VTAIL.n822 VTAIL.n754 12.8005
R1532 VTAIL.n827 VTAIL.n752 12.8005
R1533 VTAIL.n36 VTAIL.n32 12.8005
R1534 VTAIL.n80 VTAIL.n12 12.8005
R1535 VTAIL.n85 VTAIL.n10 12.8005
R1536 VTAIL.n142 VTAIL.n138 12.8005
R1537 VTAIL.n186 VTAIL.n118 12.8005
R1538 VTAIL.n191 VTAIL.n116 12.8005
R1539 VTAIL.n248 VTAIL.n244 12.8005
R1540 VTAIL.n292 VTAIL.n224 12.8005
R1541 VTAIL.n297 VTAIL.n222 12.8005
R1542 VTAIL.n721 VTAIL.n646 12.8005
R1543 VTAIL.n716 VTAIL.n648 12.8005
R1544 VTAIL.n673 VTAIL.n669 12.8005
R1545 VTAIL.n615 VTAIL.n540 12.8005
R1546 VTAIL.n610 VTAIL.n542 12.8005
R1547 VTAIL.n567 VTAIL.n563 12.8005
R1548 VTAIL.n509 VTAIL.n434 12.8005
R1549 VTAIL.n504 VTAIL.n436 12.8005
R1550 VTAIL.n461 VTAIL.n457 12.8005
R1551 VTAIL.n403 VTAIL.n328 12.8005
R1552 VTAIL.n398 VTAIL.n330 12.8005
R1553 VTAIL.n355 VTAIL.n351 12.8005
R1554 VTAIL.n782 VTAIL.n781 12.0247
R1555 VTAIL.n819 VTAIL.n818 12.0247
R1556 VTAIL.n828 VTAIL.n750 12.0247
R1557 VTAIL.n40 VTAIL.n39 12.0247
R1558 VTAIL.n77 VTAIL.n76 12.0247
R1559 VTAIL.n86 VTAIL.n8 12.0247
R1560 VTAIL.n146 VTAIL.n145 12.0247
R1561 VTAIL.n183 VTAIL.n182 12.0247
R1562 VTAIL.n192 VTAIL.n114 12.0247
R1563 VTAIL.n252 VTAIL.n251 12.0247
R1564 VTAIL.n289 VTAIL.n288 12.0247
R1565 VTAIL.n298 VTAIL.n220 12.0247
R1566 VTAIL.n722 VTAIL.n644 12.0247
R1567 VTAIL.n713 VTAIL.n712 12.0247
R1568 VTAIL.n677 VTAIL.n676 12.0247
R1569 VTAIL.n616 VTAIL.n538 12.0247
R1570 VTAIL.n607 VTAIL.n606 12.0247
R1571 VTAIL.n571 VTAIL.n570 12.0247
R1572 VTAIL.n510 VTAIL.n432 12.0247
R1573 VTAIL.n501 VTAIL.n500 12.0247
R1574 VTAIL.n465 VTAIL.n464 12.0247
R1575 VTAIL.n404 VTAIL.n326 12.0247
R1576 VTAIL.n395 VTAIL.n394 12.0247
R1577 VTAIL.n359 VTAIL.n358 12.0247
R1578 VTAIL.n785 VTAIL.n772 11.249
R1579 VTAIL.n814 VTAIL.n756 11.249
R1580 VTAIL.n832 VTAIL.n831 11.249
R1581 VTAIL.n43 VTAIL.n30 11.249
R1582 VTAIL.n72 VTAIL.n14 11.249
R1583 VTAIL.n90 VTAIL.n89 11.249
R1584 VTAIL.n149 VTAIL.n136 11.249
R1585 VTAIL.n178 VTAIL.n120 11.249
R1586 VTAIL.n196 VTAIL.n195 11.249
R1587 VTAIL.n255 VTAIL.n242 11.249
R1588 VTAIL.n284 VTAIL.n226 11.249
R1589 VTAIL.n302 VTAIL.n301 11.249
R1590 VTAIL.n726 VTAIL.n725 11.249
R1591 VTAIL.n709 VTAIL.n650 11.249
R1592 VTAIL.n680 VTAIL.n667 11.249
R1593 VTAIL.n620 VTAIL.n619 11.249
R1594 VTAIL.n603 VTAIL.n544 11.249
R1595 VTAIL.n574 VTAIL.n561 11.249
R1596 VTAIL.n514 VTAIL.n513 11.249
R1597 VTAIL.n497 VTAIL.n438 11.249
R1598 VTAIL.n468 VTAIL.n455 11.249
R1599 VTAIL.n408 VTAIL.n407 11.249
R1600 VTAIL.n391 VTAIL.n332 11.249
R1601 VTAIL.n362 VTAIL.n349 11.249
R1602 VTAIL.n786 VTAIL.n770 10.4732
R1603 VTAIL.n813 VTAIL.n758 10.4732
R1604 VTAIL.n835 VTAIL.n748 10.4732
R1605 VTAIL.n44 VTAIL.n28 10.4732
R1606 VTAIL.n71 VTAIL.n16 10.4732
R1607 VTAIL.n93 VTAIL.n6 10.4732
R1608 VTAIL.n150 VTAIL.n134 10.4732
R1609 VTAIL.n177 VTAIL.n122 10.4732
R1610 VTAIL.n199 VTAIL.n112 10.4732
R1611 VTAIL.n256 VTAIL.n240 10.4732
R1612 VTAIL.n283 VTAIL.n228 10.4732
R1613 VTAIL.n305 VTAIL.n218 10.4732
R1614 VTAIL.n729 VTAIL.n642 10.4732
R1615 VTAIL.n708 VTAIL.n653 10.4732
R1616 VTAIL.n681 VTAIL.n665 10.4732
R1617 VTAIL.n623 VTAIL.n536 10.4732
R1618 VTAIL.n602 VTAIL.n547 10.4732
R1619 VTAIL.n575 VTAIL.n559 10.4732
R1620 VTAIL.n517 VTAIL.n430 10.4732
R1621 VTAIL.n496 VTAIL.n441 10.4732
R1622 VTAIL.n469 VTAIL.n453 10.4732
R1623 VTAIL.n411 VTAIL.n324 10.4732
R1624 VTAIL.n390 VTAIL.n335 10.4732
R1625 VTAIL.n363 VTAIL.n347 10.4732
R1626 VTAIL.n790 VTAIL.n789 9.69747
R1627 VTAIL.n810 VTAIL.n809 9.69747
R1628 VTAIL.n836 VTAIL.n746 9.69747
R1629 VTAIL.n48 VTAIL.n47 9.69747
R1630 VTAIL.n68 VTAIL.n67 9.69747
R1631 VTAIL.n94 VTAIL.n4 9.69747
R1632 VTAIL.n154 VTAIL.n153 9.69747
R1633 VTAIL.n174 VTAIL.n173 9.69747
R1634 VTAIL.n200 VTAIL.n110 9.69747
R1635 VTAIL.n260 VTAIL.n259 9.69747
R1636 VTAIL.n280 VTAIL.n279 9.69747
R1637 VTAIL.n306 VTAIL.n216 9.69747
R1638 VTAIL.n730 VTAIL.n640 9.69747
R1639 VTAIL.n705 VTAIL.n704 9.69747
R1640 VTAIL.n685 VTAIL.n684 9.69747
R1641 VTAIL.n624 VTAIL.n534 9.69747
R1642 VTAIL.n599 VTAIL.n598 9.69747
R1643 VTAIL.n579 VTAIL.n578 9.69747
R1644 VTAIL.n518 VTAIL.n428 9.69747
R1645 VTAIL.n493 VTAIL.n492 9.69747
R1646 VTAIL.n473 VTAIL.n472 9.69747
R1647 VTAIL.n412 VTAIL.n322 9.69747
R1648 VTAIL.n387 VTAIL.n386 9.69747
R1649 VTAIL.n367 VTAIL.n366 9.69747
R1650 VTAIL.n846 VTAIL.n845 9.45567
R1651 VTAIL.n104 VTAIL.n103 9.45567
R1652 VTAIL.n210 VTAIL.n209 9.45567
R1653 VTAIL.n316 VTAIL.n315 9.45567
R1654 VTAIL.n740 VTAIL.n739 9.45567
R1655 VTAIL.n634 VTAIL.n633 9.45567
R1656 VTAIL.n528 VTAIL.n527 9.45567
R1657 VTAIL.n422 VTAIL.n421 9.45567
R1658 VTAIL.n744 VTAIL.n743 9.3005
R1659 VTAIL.n839 VTAIL.n838 9.3005
R1660 VTAIL.n837 VTAIL.n836 9.3005
R1661 VTAIL.n748 VTAIL.n747 9.3005
R1662 VTAIL.n831 VTAIL.n830 9.3005
R1663 VTAIL.n829 VTAIL.n828 9.3005
R1664 VTAIL.n752 VTAIL.n751 9.3005
R1665 VTAIL.n797 VTAIL.n796 9.3005
R1666 VTAIL.n795 VTAIL.n794 9.3005
R1667 VTAIL.n768 VTAIL.n767 9.3005
R1668 VTAIL.n789 VTAIL.n788 9.3005
R1669 VTAIL.n787 VTAIL.n786 9.3005
R1670 VTAIL.n772 VTAIL.n771 9.3005
R1671 VTAIL.n781 VTAIL.n780 9.3005
R1672 VTAIL.n779 VTAIL.n778 9.3005
R1673 VTAIL.n764 VTAIL.n763 9.3005
R1674 VTAIL.n803 VTAIL.n802 9.3005
R1675 VTAIL.n805 VTAIL.n804 9.3005
R1676 VTAIL.n760 VTAIL.n759 9.3005
R1677 VTAIL.n811 VTAIL.n810 9.3005
R1678 VTAIL.n813 VTAIL.n812 9.3005
R1679 VTAIL.n756 VTAIL.n755 9.3005
R1680 VTAIL.n820 VTAIL.n819 9.3005
R1681 VTAIL.n822 VTAIL.n821 9.3005
R1682 VTAIL.n845 VTAIL.n844 9.3005
R1683 VTAIL.n2 VTAIL.n1 9.3005
R1684 VTAIL.n97 VTAIL.n96 9.3005
R1685 VTAIL.n95 VTAIL.n94 9.3005
R1686 VTAIL.n6 VTAIL.n5 9.3005
R1687 VTAIL.n89 VTAIL.n88 9.3005
R1688 VTAIL.n87 VTAIL.n86 9.3005
R1689 VTAIL.n10 VTAIL.n9 9.3005
R1690 VTAIL.n55 VTAIL.n54 9.3005
R1691 VTAIL.n53 VTAIL.n52 9.3005
R1692 VTAIL.n26 VTAIL.n25 9.3005
R1693 VTAIL.n47 VTAIL.n46 9.3005
R1694 VTAIL.n45 VTAIL.n44 9.3005
R1695 VTAIL.n30 VTAIL.n29 9.3005
R1696 VTAIL.n39 VTAIL.n38 9.3005
R1697 VTAIL.n37 VTAIL.n36 9.3005
R1698 VTAIL.n22 VTAIL.n21 9.3005
R1699 VTAIL.n61 VTAIL.n60 9.3005
R1700 VTAIL.n63 VTAIL.n62 9.3005
R1701 VTAIL.n18 VTAIL.n17 9.3005
R1702 VTAIL.n69 VTAIL.n68 9.3005
R1703 VTAIL.n71 VTAIL.n70 9.3005
R1704 VTAIL.n14 VTAIL.n13 9.3005
R1705 VTAIL.n78 VTAIL.n77 9.3005
R1706 VTAIL.n80 VTAIL.n79 9.3005
R1707 VTAIL.n103 VTAIL.n102 9.3005
R1708 VTAIL.n108 VTAIL.n107 9.3005
R1709 VTAIL.n203 VTAIL.n202 9.3005
R1710 VTAIL.n201 VTAIL.n200 9.3005
R1711 VTAIL.n112 VTAIL.n111 9.3005
R1712 VTAIL.n195 VTAIL.n194 9.3005
R1713 VTAIL.n193 VTAIL.n192 9.3005
R1714 VTAIL.n116 VTAIL.n115 9.3005
R1715 VTAIL.n161 VTAIL.n160 9.3005
R1716 VTAIL.n159 VTAIL.n158 9.3005
R1717 VTAIL.n132 VTAIL.n131 9.3005
R1718 VTAIL.n153 VTAIL.n152 9.3005
R1719 VTAIL.n151 VTAIL.n150 9.3005
R1720 VTAIL.n136 VTAIL.n135 9.3005
R1721 VTAIL.n145 VTAIL.n144 9.3005
R1722 VTAIL.n143 VTAIL.n142 9.3005
R1723 VTAIL.n128 VTAIL.n127 9.3005
R1724 VTAIL.n167 VTAIL.n166 9.3005
R1725 VTAIL.n169 VTAIL.n168 9.3005
R1726 VTAIL.n124 VTAIL.n123 9.3005
R1727 VTAIL.n175 VTAIL.n174 9.3005
R1728 VTAIL.n177 VTAIL.n176 9.3005
R1729 VTAIL.n120 VTAIL.n119 9.3005
R1730 VTAIL.n184 VTAIL.n183 9.3005
R1731 VTAIL.n186 VTAIL.n185 9.3005
R1732 VTAIL.n209 VTAIL.n208 9.3005
R1733 VTAIL.n214 VTAIL.n213 9.3005
R1734 VTAIL.n309 VTAIL.n308 9.3005
R1735 VTAIL.n307 VTAIL.n306 9.3005
R1736 VTAIL.n218 VTAIL.n217 9.3005
R1737 VTAIL.n301 VTAIL.n300 9.3005
R1738 VTAIL.n299 VTAIL.n298 9.3005
R1739 VTAIL.n222 VTAIL.n221 9.3005
R1740 VTAIL.n267 VTAIL.n266 9.3005
R1741 VTAIL.n265 VTAIL.n264 9.3005
R1742 VTAIL.n238 VTAIL.n237 9.3005
R1743 VTAIL.n259 VTAIL.n258 9.3005
R1744 VTAIL.n257 VTAIL.n256 9.3005
R1745 VTAIL.n242 VTAIL.n241 9.3005
R1746 VTAIL.n251 VTAIL.n250 9.3005
R1747 VTAIL.n249 VTAIL.n248 9.3005
R1748 VTAIL.n234 VTAIL.n233 9.3005
R1749 VTAIL.n273 VTAIL.n272 9.3005
R1750 VTAIL.n275 VTAIL.n274 9.3005
R1751 VTAIL.n230 VTAIL.n229 9.3005
R1752 VTAIL.n281 VTAIL.n280 9.3005
R1753 VTAIL.n283 VTAIL.n282 9.3005
R1754 VTAIL.n226 VTAIL.n225 9.3005
R1755 VTAIL.n290 VTAIL.n289 9.3005
R1756 VTAIL.n292 VTAIL.n291 9.3005
R1757 VTAIL.n315 VTAIL.n314 9.3005
R1758 VTAIL.n698 VTAIL.n697 9.3005
R1759 VTAIL.n700 VTAIL.n699 9.3005
R1760 VTAIL.n655 VTAIL.n654 9.3005
R1761 VTAIL.n706 VTAIL.n705 9.3005
R1762 VTAIL.n708 VTAIL.n707 9.3005
R1763 VTAIL.n650 VTAIL.n649 9.3005
R1764 VTAIL.n714 VTAIL.n713 9.3005
R1765 VTAIL.n716 VTAIL.n715 9.3005
R1766 VTAIL.n739 VTAIL.n738 9.3005
R1767 VTAIL.n638 VTAIL.n637 9.3005
R1768 VTAIL.n733 VTAIL.n732 9.3005
R1769 VTAIL.n731 VTAIL.n730 9.3005
R1770 VTAIL.n642 VTAIL.n641 9.3005
R1771 VTAIL.n725 VTAIL.n724 9.3005
R1772 VTAIL.n723 VTAIL.n722 9.3005
R1773 VTAIL.n646 VTAIL.n645 9.3005
R1774 VTAIL.n659 VTAIL.n658 9.3005
R1775 VTAIL.n692 VTAIL.n691 9.3005
R1776 VTAIL.n690 VTAIL.n689 9.3005
R1777 VTAIL.n663 VTAIL.n662 9.3005
R1778 VTAIL.n684 VTAIL.n683 9.3005
R1779 VTAIL.n682 VTAIL.n681 9.3005
R1780 VTAIL.n667 VTAIL.n666 9.3005
R1781 VTAIL.n676 VTAIL.n675 9.3005
R1782 VTAIL.n674 VTAIL.n673 9.3005
R1783 VTAIL.n592 VTAIL.n591 9.3005
R1784 VTAIL.n594 VTAIL.n593 9.3005
R1785 VTAIL.n549 VTAIL.n548 9.3005
R1786 VTAIL.n600 VTAIL.n599 9.3005
R1787 VTAIL.n602 VTAIL.n601 9.3005
R1788 VTAIL.n544 VTAIL.n543 9.3005
R1789 VTAIL.n608 VTAIL.n607 9.3005
R1790 VTAIL.n610 VTAIL.n609 9.3005
R1791 VTAIL.n633 VTAIL.n632 9.3005
R1792 VTAIL.n532 VTAIL.n531 9.3005
R1793 VTAIL.n627 VTAIL.n626 9.3005
R1794 VTAIL.n625 VTAIL.n624 9.3005
R1795 VTAIL.n536 VTAIL.n535 9.3005
R1796 VTAIL.n619 VTAIL.n618 9.3005
R1797 VTAIL.n617 VTAIL.n616 9.3005
R1798 VTAIL.n540 VTAIL.n539 9.3005
R1799 VTAIL.n553 VTAIL.n552 9.3005
R1800 VTAIL.n586 VTAIL.n585 9.3005
R1801 VTAIL.n584 VTAIL.n583 9.3005
R1802 VTAIL.n557 VTAIL.n556 9.3005
R1803 VTAIL.n578 VTAIL.n577 9.3005
R1804 VTAIL.n576 VTAIL.n575 9.3005
R1805 VTAIL.n561 VTAIL.n560 9.3005
R1806 VTAIL.n570 VTAIL.n569 9.3005
R1807 VTAIL.n568 VTAIL.n567 9.3005
R1808 VTAIL.n486 VTAIL.n485 9.3005
R1809 VTAIL.n488 VTAIL.n487 9.3005
R1810 VTAIL.n443 VTAIL.n442 9.3005
R1811 VTAIL.n494 VTAIL.n493 9.3005
R1812 VTAIL.n496 VTAIL.n495 9.3005
R1813 VTAIL.n438 VTAIL.n437 9.3005
R1814 VTAIL.n502 VTAIL.n501 9.3005
R1815 VTAIL.n504 VTAIL.n503 9.3005
R1816 VTAIL.n527 VTAIL.n526 9.3005
R1817 VTAIL.n426 VTAIL.n425 9.3005
R1818 VTAIL.n521 VTAIL.n520 9.3005
R1819 VTAIL.n519 VTAIL.n518 9.3005
R1820 VTAIL.n430 VTAIL.n429 9.3005
R1821 VTAIL.n513 VTAIL.n512 9.3005
R1822 VTAIL.n511 VTAIL.n510 9.3005
R1823 VTAIL.n434 VTAIL.n433 9.3005
R1824 VTAIL.n447 VTAIL.n446 9.3005
R1825 VTAIL.n480 VTAIL.n479 9.3005
R1826 VTAIL.n478 VTAIL.n477 9.3005
R1827 VTAIL.n451 VTAIL.n450 9.3005
R1828 VTAIL.n472 VTAIL.n471 9.3005
R1829 VTAIL.n470 VTAIL.n469 9.3005
R1830 VTAIL.n455 VTAIL.n454 9.3005
R1831 VTAIL.n464 VTAIL.n463 9.3005
R1832 VTAIL.n462 VTAIL.n461 9.3005
R1833 VTAIL.n380 VTAIL.n379 9.3005
R1834 VTAIL.n382 VTAIL.n381 9.3005
R1835 VTAIL.n337 VTAIL.n336 9.3005
R1836 VTAIL.n388 VTAIL.n387 9.3005
R1837 VTAIL.n390 VTAIL.n389 9.3005
R1838 VTAIL.n332 VTAIL.n331 9.3005
R1839 VTAIL.n396 VTAIL.n395 9.3005
R1840 VTAIL.n398 VTAIL.n397 9.3005
R1841 VTAIL.n421 VTAIL.n420 9.3005
R1842 VTAIL.n320 VTAIL.n319 9.3005
R1843 VTAIL.n415 VTAIL.n414 9.3005
R1844 VTAIL.n413 VTAIL.n412 9.3005
R1845 VTAIL.n324 VTAIL.n323 9.3005
R1846 VTAIL.n407 VTAIL.n406 9.3005
R1847 VTAIL.n405 VTAIL.n404 9.3005
R1848 VTAIL.n328 VTAIL.n327 9.3005
R1849 VTAIL.n341 VTAIL.n340 9.3005
R1850 VTAIL.n374 VTAIL.n373 9.3005
R1851 VTAIL.n372 VTAIL.n371 9.3005
R1852 VTAIL.n345 VTAIL.n344 9.3005
R1853 VTAIL.n366 VTAIL.n365 9.3005
R1854 VTAIL.n364 VTAIL.n363 9.3005
R1855 VTAIL.n349 VTAIL.n348 9.3005
R1856 VTAIL.n358 VTAIL.n357 9.3005
R1857 VTAIL.n356 VTAIL.n355 9.3005
R1858 VTAIL.n793 VTAIL.n768 8.92171
R1859 VTAIL.n806 VTAIL.n760 8.92171
R1860 VTAIL.n840 VTAIL.n839 8.92171
R1861 VTAIL.n51 VTAIL.n26 8.92171
R1862 VTAIL.n64 VTAIL.n18 8.92171
R1863 VTAIL.n98 VTAIL.n97 8.92171
R1864 VTAIL.n157 VTAIL.n132 8.92171
R1865 VTAIL.n170 VTAIL.n124 8.92171
R1866 VTAIL.n204 VTAIL.n203 8.92171
R1867 VTAIL.n263 VTAIL.n238 8.92171
R1868 VTAIL.n276 VTAIL.n230 8.92171
R1869 VTAIL.n310 VTAIL.n309 8.92171
R1870 VTAIL.n734 VTAIL.n733 8.92171
R1871 VTAIL.n701 VTAIL.n655 8.92171
R1872 VTAIL.n688 VTAIL.n663 8.92171
R1873 VTAIL.n628 VTAIL.n627 8.92171
R1874 VTAIL.n595 VTAIL.n549 8.92171
R1875 VTAIL.n582 VTAIL.n557 8.92171
R1876 VTAIL.n522 VTAIL.n521 8.92171
R1877 VTAIL.n489 VTAIL.n443 8.92171
R1878 VTAIL.n476 VTAIL.n451 8.92171
R1879 VTAIL.n416 VTAIL.n415 8.92171
R1880 VTAIL.n383 VTAIL.n337 8.92171
R1881 VTAIL.n370 VTAIL.n345 8.92171
R1882 VTAIL.n794 VTAIL.n766 8.14595
R1883 VTAIL.n805 VTAIL.n762 8.14595
R1884 VTAIL.n843 VTAIL.n744 8.14595
R1885 VTAIL.n52 VTAIL.n24 8.14595
R1886 VTAIL.n63 VTAIL.n20 8.14595
R1887 VTAIL.n101 VTAIL.n2 8.14595
R1888 VTAIL.n158 VTAIL.n130 8.14595
R1889 VTAIL.n169 VTAIL.n126 8.14595
R1890 VTAIL.n207 VTAIL.n108 8.14595
R1891 VTAIL.n264 VTAIL.n236 8.14595
R1892 VTAIL.n275 VTAIL.n232 8.14595
R1893 VTAIL.n313 VTAIL.n214 8.14595
R1894 VTAIL.n737 VTAIL.n638 8.14595
R1895 VTAIL.n700 VTAIL.n657 8.14595
R1896 VTAIL.n689 VTAIL.n661 8.14595
R1897 VTAIL.n631 VTAIL.n532 8.14595
R1898 VTAIL.n594 VTAIL.n551 8.14595
R1899 VTAIL.n583 VTAIL.n555 8.14595
R1900 VTAIL.n525 VTAIL.n426 8.14595
R1901 VTAIL.n488 VTAIL.n445 8.14595
R1902 VTAIL.n477 VTAIL.n449 8.14595
R1903 VTAIL.n419 VTAIL.n320 8.14595
R1904 VTAIL.n382 VTAIL.n339 8.14595
R1905 VTAIL.n371 VTAIL.n343 8.14595
R1906 VTAIL.n798 VTAIL.n797 7.3702
R1907 VTAIL.n802 VTAIL.n801 7.3702
R1908 VTAIL.n844 VTAIL.n742 7.3702
R1909 VTAIL.n56 VTAIL.n55 7.3702
R1910 VTAIL.n60 VTAIL.n59 7.3702
R1911 VTAIL.n102 VTAIL.n0 7.3702
R1912 VTAIL.n162 VTAIL.n161 7.3702
R1913 VTAIL.n166 VTAIL.n165 7.3702
R1914 VTAIL.n208 VTAIL.n106 7.3702
R1915 VTAIL.n268 VTAIL.n267 7.3702
R1916 VTAIL.n272 VTAIL.n271 7.3702
R1917 VTAIL.n314 VTAIL.n212 7.3702
R1918 VTAIL.n738 VTAIL.n636 7.3702
R1919 VTAIL.n697 VTAIL.n696 7.3702
R1920 VTAIL.n693 VTAIL.n692 7.3702
R1921 VTAIL.n632 VTAIL.n530 7.3702
R1922 VTAIL.n591 VTAIL.n590 7.3702
R1923 VTAIL.n587 VTAIL.n586 7.3702
R1924 VTAIL.n526 VTAIL.n424 7.3702
R1925 VTAIL.n485 VTAIL.n484 7.3702
R1926 VTAIL.n481 VTAIL.n480 7.3702
R1927 VTAIL.n420 VTAIL.n318 7.3702
R1928 VTAIL.n379 VTAIL.n378 7.3702
R1929 VTAIL.n375 VTAIL.n374 7.3702
R1930 VTAIL.n798 VTAIL.n764 6.59444
R1931 VTAIL.n801 VTAIL.n764 6.59444
R1932 VTAIL.n846 VTAIL.n742 6.59444
R1933 VTAIL.n56 VTAIL.n22 6.59444
R1934 VTAIL.n59 VTAIL.n22 6.59444
R1935 VTAIL.n104 VTAIL.n0 6.59444
R1936 VTAIL.n162 VTAIL.n128 6.59444
R1937 VTAIL.n165 VTAIL.n128 6.59444
R1938 VTAIL.n210 VTAIL.n106 6.59444
R1939 VTAIL.n268 VTAIL.n234 6.59444
R1940 VTAIL.n271 VTAIL.n234 6.59444
R1941 VTAIL.n316 VTAIL.n212 6.59444
R1942 VTAIL.n740 VTAIL.n636 6.59444
R1943 VTAIL.n696 VTAIL.n659 6.59444
R1944 VTAIL.n693 VTAIL.n659 6.59444
R1945 VTAIL.n634 VTAIL.n530 6.59444
R1946 VTAIL.n590 VTAIL.n553 6.59444
R1947 VTAIL.n587 VTAIL.n553 6.59444
R1948 VTAIL.n528 VTAIL.n424 6.59444
R1949 VTAIL.n484 VTAIL.n447 6.59444
R1950 VTAIL.n481 VTAIL.n447 6.59444
R1951 VTAIL.n422 VTAIL.n318 6.59444
R1952 VTAIL.n378 VTAIL.n341 6.59444
R1953 VTAIL.n375 VTAIL.n341 6.59444
R1954 VTAIL.n797 VTAIL.n766 5.81868
R1955 VTAIL.n802 VTAIL.n762 5.81868
R1956 VTAIL.n844 VTAIL.n843 5.81868
R1957 VTAIL.n55 VTAIL.n24 5.81868
R1958 VTAIL.n60 VTAIL.n20 5.81868
R1959 VTAIL.n102 VTAIL.n101 5.81868
R1960 VTAIL.n161 VTAIL.n130 5.81868
R1961 VTAIL.n166 VTAIL.n126 5.81868
R1962 VTAIL.n208 VTAIL.n207 5.81868
R1963 VTAIL.n267 VTAIL.n236 5.81868
R1964 VTAIL.n272 VTAIL.n232 5.81868
R1965 VTAIL.n314 VTAIL.n313 5.81868
R1966 VTAIL.n738 VTAIL.n737 5.81868
R1967 VTAIL.n697 VTAIL.n657 5.81868
R1968 VTAIL.n692 VTAIL.n661 5.81868
R1969 VTAIL.n632 VTAIL.n631 5.81868
R1970 VTAIL.n591 VTAIL.n551 5.81868
R1971 VTAIL.n586 VTAIL.n555 5.81868
R1972 VTAIL.n526 VTAIL.n525 5.81868
R1973 VTAIL.n485 VTAIL.n445 5.81868
R1974 VTAIL.n480 VTAIL.n449 5.81868
R1975 VTAIL.n420 VTAIL.n419 5.81868
R1976 VTAIL.n379 VTAIL.n339 5.81868
R1977 VTAIL.n374 VTAIL.n343 5.81868
R1978 VTAIL.n794 VTAIL.n793 5.04292
R1979 VTAIL.n806 VTAIL.n805 5.04292
R1980 VTAIL.n840 VTAIL.n744 5.04292
R1981 VTAIL.n52 VTAIL.n51 5.04292
R1982 VTAIL.n64 VTAIL.n63 5.04292
R1983 VTAIL.n98 VTAIL.n2 5.04292
R1984 VTAIL.n158 VTAIL.n157 5.04292
R1985 VTAIL.n170 VTAIL.n169 5.04292
R1986 VTAIL.n204 VTAIL.n108 5.04292
R1987 VTAIL.n264 VTAIL.n263 5.04292
R1988 VTAIL.n276 VTAIL.n275 5.04292
R1989 VTAIL.n310 VTAIL.n214 5.04292
R1990 VTAIL.n734 VTAIL.n638 5.04292
R1991 VTAIL.n701 VTAIL.n700 5.04292
R1992 VTAIL.n689 VTAIL.n688 5.04292
R1993 VTAIL.n628 VTAIL.n532 5.04292
R1994 VTAIL.n595 VTAIL.n594 5.04292
R1995 VTAIL.n583 VTAIL.n582 5.04292
R1996 VTAIL.n522 VTAIL.n426 5.04292
R1997 VTAIL.n489 VTAIL.n488 5.04292
R1998 VTAIL.n477 VTAIL.n476 5.04292
R1999 VTAIL.n416 VTAIL.n320 5.04292
R2000 VTAIL.n383 VTAIL.n382 5.04292
R2001 VTAIL.n371 VTAIL.n370 5.04292
R2002 VTAIL.n790 VTAIL.n768 4.26717
R2003 VTAIL.n809 VTAIL.n760 4.26717
R2004 VTAIL.n839 VTAIL.n746 4.26717
R2005 VTAIL.n48 VTAIL.n26 4.26717
R2006 VTAIL.n67 VTAIL.n18 4.26717
R2007 VTAIL.n97 VTAIL.n4 4.26717
R2008 VTAIL.n154 VTAIL.n132 4.26717
R2009 VTAIL.n173 VTAIL.n124 4.26717
R2010 VTAIL.n203 VTAIL.n110 4.26717
R2011 VTAIL.n260 VTAIL.n238 4.26717
R2012 VTAIL.n279 VTAIL.n230 4.26717
R2013 VTAIL.n309 VTAIL.n216 4.26717
R2014 VTAIL.n733 VTAIL.n640 4.26717
R2015 VTAIL.n704 VTAIL.n655 4.26717
R2016 VTAIL.n685 VTAIL.n663 4.26717
R2017 VTAIL.n627 VTAIL.n534 4.26717
R2018 VTAIL.n598 VTAIL.n549 4.26717
R2019 VTAIL.n579 VTAIL.n557 4.26717
R2020 VTAIL.n521 VTAIL.n428 4.26717
R2021 VTAIL.n492 VTAIL.n443 4.26717
R2022 VTAIL.n473 VTAIL.n451 4.26717
R2023 VTAIL.n415 VTAIL.n322 4.26717
R2024 VTAIL.n386 VTAIL.n337 4.26717
R2025 VTAIL.n367 VTAIL.n345 4.26717
R2026 VTAIL.n779 VTAIL.n775 3.70982
R2027 VTAIL.n37 VTAIL.n33 3.70982
R2028 VTAIL.n143 VTAIL.n139 3.70982
R2029 VTAIL.n249 VTAIL.n245 3.70982
R2030 VTAIL.n674 VTAIL.n670 3.70982
R2031 VTAIL.n568 VTAIL.n564 3.70982
R2032 VTAIL.n462 VTAIL.n458 3.70982
R2033 VTAIL.n356 VTAIL.n352 3.70982
R2034 VTAIL.n789 VTAIL.n770 3.49141
R2035 VTAIL.n810 VTAIL.n758 3.49141
R2036 VTAIL.n836 VTAIL.n835 3.49141
R2037 VTAIL.n47 VTAIL.n28 3.49141
R2038 VTAIL.n68 VTAIL.n16 3.49141
R2039 VTAIL.n94 VTAIL.n93 3.49141
R2040 VTAIL.n153 VTAIL.n134 3.49141
R2041 VTAIL.n174 VTAIL.n122 3.49141
R2042 VTAIL.n200 VTAIL.n199 3.49141
R2043 VTAIL.n259 VTAIL.n240 3.49141
R2044 VTAIL.n280 VTAIL.n228 3.49141
R2045 VTAIL.n306 VTAIL.n305 3.49141
R2046 VTAIL.n730 VTAIL.n729 3.49141
R2047 VTAIL.n705 VTAIL.n653 3.49141
R2048 VTAIL.n684 VTAIL.n665 3.49141
R2049 VTAIL.n624 VTAIL.n623 3.49141
R2050 VTAIL.n599 VTAIL.n547 3.49141
R2051 VTAIL.n578 VTAIL.n559 3.49141
R2052 VTAIL.n518 VTAIL.n517 3.49141
R2053 VTAIL.n493 VTAIL.n441 3.49141
R2054 VTAIL.n472 VTAIL.n453 3.49141
R2055 VTAIL.n412 VTAIL.n411 3.49141
R2056 VTAIL.n387 VTAIL.n335 3.49141
R2057 VTAIL.n366 VTAIL.n347 3.49141
R2058 VTAIL.n786 VTAIL.n785 2.71565
R2059 VTAIL.n814 VTAIL.n813 2.71565
R2060 VTAIL.n832 VTAIL.n748 2.71565
R2061 VTAIL.n44 VTAIL.n43 2.71565
R2062 VTAIL.n72 VTAIL.n71 2.71565
R2063 VTAIL.n90 VTAIL.n6 2.71565
R2064 VTAIL.n150 VTAIL.n149 2.71565
R2065 VTAIL.n178 VTAIL.n177 2.71565
R2066 VTAIL.n196 VTAIL.n112 2.71565
R2067 VTAIL.n256 VTAIL.n255 2.71565
R2068 VTAIL.n284 VTAIL.n283 2.71565
R2069 VTAIL.n302 VTAIL.n218 2.71565
R2070 VTAIL.n726 VTAIL.n642 2.71565
R2071 VTAIL.n709 VTAIL.n708 2.71565
R2072 VTAIL.n681 VTAIL.n680 2.71565
R2073 VTAIL.n620 VTAIL.n536 2.71565
R2074 VTAIL.n603 VTAIL.n602 2.71565
R2075 VTAIL.n575 VTAIL.n574 2.71565
R2076 VTAIL.n514 VTAIL.n430 2.71565
R2077 VTAIL.n497 VTAIL.n496 2.71565
R2078 VTAIL.n469 VTAIL.n468 2.71565
R2079 VTAIL.n408 VTAIL.n324 2.71565
R2080 VTAIL.n391 VTAIL.n390 2.71565
R2081 VTAIL.n363 VTAIL.n362 2.71565
R2082 VTAIL.n782 VTAIL.n772 1.93989
R2083 VTAIL.n818 VTAIL.n756 1.93989
R2084 VTAIL.n831 VTAIL.n750 1.93989
R2085 VTAIL.n40 VTAIL.n30 1.93989
R2086 VTAIL.n76 VTAIL.n14 1.93989
R2087 VTAIL.n89 VTAIL.n8 1.93989
R2088 VTAIL.n146 VTAIL.n136 1.93989
R2089 VTAIL.n182 VTAIL.n120 1.93989
R2090 VTAIL.n195 VTAIL.n114 1.93989
R2091 VTAIL.n252 VTAIL.n242 1.93989
R2092 VTAIL.n288 VTAIL.n226 1.93989
R2093 VTAIL.n301 VTAIL.n220 1.93989
R2094 VTAIL.n725 VTAIL.n644 1.93989
R2095 VTAIL.n712 VTAIL.n650 1.93989
R2096 VTAIL.n677 VTAIL.n667 1.93989
R2097 VTAIL.n619 VTAIL.n538 1.93989
R2098 VTAIL.n606 VTAIL.n544 1.93989
R2099 VTAIL.n571 VTAIL.n561 1.93989
R2100 VTAIL.n513 VTAIL.n432 1.93989
R2101 VTAIL.n500 VTAIL.n438 1.93989
R2102 VTAIL.n465 VTAIL.n455 1.93989
R2103 VTAIL.n407 VTAIL.n326 1.93989
R2104 VTAIL.n394 VTAIL.n332 1.93989
R2105 VTAIL.n359 VTAIL.n349 1.93989
R2106 VTAIL.n781 VTAIL.n774 1.16414
R2107 VTAIL.n819 VTAIL.n754 1.16414
R2108 VTAIL.n828 VTAIL.n827 1.16414
R2109 VTAIL.n39 VTAIL.n32 1.16414
R2110 VTAIL.n77 VTAIL.n12 1.16414
R2111 VTAIL.n86 VTAIL.n85 1.16414
R2112 VTAIL.n145 VTAIL.n138 1.16414
R2113 VTAIL.n183 VTAIL.n118 1.16414
R2114 VTAIL.n192 VTAIL.n191 1.16414
R2115 VTAIL.n251 VTAIL.n244 1.16414
R2116 VTAIL.n289 VTAIL.n224 1.16414
R2117 VTAIL.n298 VTAIL.n297 1.16414
R2118 VTAIL.n722 VTAIL.n721 1.16414
R2119 VTAIL.n713 VTAIL.n648 1.16414
R2120 VTAIL.n676 VTAIL.n669 1.16414
R2121 VTAIL.n616 VTAIL.n615 1.16414
R2122 VTAIL.n607 VTAIL.n542 1.16414
R2123 VTAIL.n570 VTAIL.n563 1.16414
R2124 VTAIL.n510 VTAIL.n509 1.16414
R2125 VTAIL.n501 VTAIL.n436 1.16414
R2126 VTAIL.n464 VTAIL.n457 1.16414
R2127 VTAIL.n404 VTAIL.n403 1.16414
R2128 VTAIL.n395 VTAIL.n330 1.16414
R2129 VTAIL.n358 VTAIL.n351 1.16414
R2130 VTAIL.n529 VTAIL.n423 1.09533
R2131 VTAIL.n741 VTAIL.n635 1.09533
R2132 VTAIL.n317 VTAIL.n211 1.09533
R2133 VTAIL VTAIL.n105 0.606103
R2134 VTAIL VTAIL.n847 0.489724
R2135 VTAIL.n635 VTAIL.n529 0.470328
R2136 VTAIL.n211 VTAIL.n105 0.470328
R2137 VTAIL.n778 VTAIL.n777 0.388379
R2138 VTAIL.n823 VTAIL.n822 0.388379
R2139 VTAIL.n824 VTAIL.n752 0.388379
R2140 VTAIL.n36 VTAIL.n35 0.388379
R2141 VTAIL.n81 VTAIL.n80 0.388379
R2142 VTAIL.n82 VTAIL.n10 0.388379
R2143 VTAIL.n142 VTAIL.n141 0.388379
R2144 VTAIL.n187 VTAIL.n186 0.388379
R2145 VTAIL.n188 VTAIL.n116 0.388379
R2146 VTAIL.n248 VTAIL.n247 0.388379
R2147 VTAIL.n293 VTAIL.n292 0.388379
R2148 VTAIL.n294 VTAIL.n222 0.388379
R2149 VTAIL.n718 VTAIL.n646 0.388379
R2150 VTAIL.n717 VTAIL.n716 0.388379
R2151 VTAIL.n673 VTAIL.n672 0.388379
R2152 VTAIL.n612 VTAIL.n540 0.388379
R2153 VTAIL.n611 VTAIL.n610 0.388379
R2154 VTAIL.n567 VTAIL.n566 0.388379
R2155 VTAIL.n506 VTAIL.n434 0.388379
R2156 VTAIL.n505 VTAIL.n504 0.388379
R2157 VTAIL.n461 VTAIL.n460 0.388379
R2158 VTAIL.n400 VTAIL.n328 0.388379
R2159 VTAIL.n399 VTAIL.n398 0.388379
R2160 VTAIL.n355 VTAIL.n354 0.388379
R2161 VTAIL.n780 VTAIL.n779 0.155672
R2162 VTAIL.n780 VTAIL.n771 0.155672
R2163 VTAIL.n787 VTAIL.n771 0.155672
R2164 VTAIL.n788 VTAIL.n787 0.155672
R2165 VTAIL.n788 VTAIL.n767 0.155672
R2166 VTAIL.n795 VTAIL.n767 0.155672
R2167 VTAIL.n796 VTAIL.n795 0.155672
R2168 VTAIL.n796 VTAIL.n763 0.155672
R2169 VTAIL.n803 VTAIL.n763 0.155672
R2170 VTAIL.n804 VTAIL.n803 0.155672
R2171 VTAIL.n804 VTAIL.n759 0.155672
R2172 VTAIL.n811 VTAIL.n759 0.155672
R2173 VTAIL.n812 VTAIL.n811 0.155672
R2174 VTAIL.n812 VTAIL.n755 0.155672
R2175 VTAIL.n820 VTAIL.n755 0.155672
R2176 VTAIL.n821 VTAIL.n820 0.155672
R2177 VTAIL.n821 VTAIL.n751 0.155672
R2178 VTAIL.n829 VTAIL.n751 0.155672
R2179 VTAIL.n830 VTAIL.n829 0.155672
R2180 VTAIL.n830 VTAIL.n747 0.155672
R2181 VTAIL.n837 VTAIL.n747 0.155672
R2182 VTAIL.n838 VTAIL.n837 0.155672
R2183 VTAIL.n838 VTAIL.n743 0.155672
R2184 VTAIL.n845 VTAIL.n743 0.155672
R2185 VTAIL.n38 VTAIL.n37 0.155672
R2186 VTAIL.n38 VTAIL.n29 0.155672
R2187 VTAIL.n45 VTAIL.n29 0.155672
R2188 VTAIL.n46 VTAIL.n45 0.155672
R2189 VTAIL.n46 VTAIL.n25 0.155672
R2190 VTAIL.n53 VTAIL.n25 0.155672
R2191 VTAIL.n54 VTAIL.n53 0.155672
R2192 VTAIL.n54 VTAIL.n21 0.155672
R2193 VTAIL.n61 VTAIL.n21 0.155672
R2194 VTAIL.n62 VTAIL.n61 0.155672
R2195 VTAIL.n62 VTAIL.n17 0.155672
R2196 VTAIL.n69 VTAIL.n17 0.155672
R2197 VTAIL.n70 VTAIL.n69 0.155672
R2198 VTAIL.n70 VTAIL.n13 0.155672
R2199 VTAIL.n78 VTAIL.n13 0.155672
R2200 VTAIL.n79 VTAIL.n78 0.155672
R2201 VTAIL.n79 VTAIL.n9 0.155672
R2202 VTAIL.n87 VTAIL.n9 0.155672
R2203 VTAIL.n88 VTAIL.n87 0.155672
R2204 VTAIL.n88 VTAIL.n5 0.155672
R2205 VTAIL.n95 VTAIL.n5 0.155672
R2206 VTAIL.n96 VTAIL.n95 0.155672
R2207 VTAIL.n96 VTAIL.n1 0.155672
R2208 VTAIL.n103 VTAIL.n1 0.155672
R2209 VTAIL.n144 VTAIL.n143 0.155672
R2210 VTAIL.n144 VTAIL.n135 0.155672
R2211 VTAIL.n151 VTAIL.n135 0.155672
R2212 VTAIL.n152 VTAIL.n151 0.155672
R2213 VTAIL.n152 VTAIL.n131 0.155672
R2214 VTAIL.n159 VTAIL.n131 0.155672
R2215 VTAIL.n160 VTAIL.n159 0.155672
R2216 VTAIL.n160 VTAIL.n127 0.155672
R2217 VTAIL.n167 VTAIL.n127 0.155672
R2218 VTAIL.n168 VTAIL.n167 0.155672
R2219 VTAIL.n168 VTAIL.n123 0.155672
R2220 VTAIL.n175 VTAIL.n123 0.155672
R2221 VTAIL.n176 VTAIL.n175 0.155672
R2222 VTAIL.n176 VTAIL.n119 0.155672
R2223 VTAIL.n184 VTAIL.n119 0.155672
R2224 VTAIL.n185 VTAIL.n184 0.155672
R2225 VTAIL.n185 VTAIL.n115 0.155672
R2226 VTAIL.n193 VTAIL.n115 0.155672
R2227 VTAIL.n194 VTAIL.n193 0.155672
R2228 VTAIL.n194 VTAIL.n111 0.155672
R2229 VTAIL.n201 VTAIL.n111 0.155672
R2230 VTAIL.n202 VTAIL.n201 0.155672
R2231 VTAIL.n202 VTAIL.n107 0.155672
R2232 VTAIL.n209 VTAIL.n107 0.155672
R2233 VTAIL.n250 VTAIL.n249 0.155672
R2234 VTAIL.n250 VTAIL.n241 0.155672
R2235 VTAIL.n257 VTAIL.n241 0.155672
R2236 VTAIL.n258 VTAIL.n257 0.155672
R2237 VTAIL.n258 VTAIL.n237 0.155672
R2238 VTAIL.n265 VTAIL.n237 0.155672
R2239 VTAIL.n266 VTAIL.n265 0.155672
R2240 VTAIL.n266 VTAIL.n233 0.155672
R2241 VTAIL.n273 VTAIL.n233 0.155672
R2242 VTAIL.n274 VTAIL.n273 0.155672
R2243 VTAIL.n274 VTAIL.n229 0.155672
R2244 VTAIL.n281 VTAIL.n229 0.155672
R2245 VTAIL.n282 VTAIL.n281 0.155672
R2246 VTAIL.n282 VTAIL.n225 0.155672
R2247 VTAIL.n290 VTAIL.n225 0.155672
R2248 VTAIL.n291 VTAIL.n290 0.155672
R2249 VTAIL.n291 VTAIL.n221 0.155672
R2250 VTAIL.n299 VTAIL.n221 0.155672
R2251 VTAIL.n300 VTAIL.n299 0.155672
R2252 VTAIL.n300 VTAIL.n217 0.155672
R2253 VTAIL.n307 VTAIL.n217 0.155672
R2254 VTAIL.n308 VTAIL.n307 0.155672
R2255 VTAIL.n308 VTAIL.n213 0.155672
R2256 VTAIL.n315 VTAIL.n213 0.155672
R2257 VTAIL.n739 VTAIL.n637 0.155672
R2258 VTAIL.n732 VTAIL.n637 0.155672
R2259 VTAIL.n732 VTAIL.n731 0.155672
R2260 VTAIL.n731 VTAIL.n641 0.155672
R2261 VTAIL.n724 VTAIL.n641 0.155672
R2262 VTAIL.n724 VTAIL.n723 0.155672
R2263 VTAIL.n723 VTAIL.n645 0.155672
R2264 VTAIL.n715 VTAIL.n645 0.155672
R2265 VTAIL.n715 VTAIL.n714 0.155672
R2266 VTAIL.n714 VTAIL.n649 0.155672
R2267 VTAIL.n707 VTAIL.n649 0.155672
R2268 VTAIL.n707 VTAIL.n706 0.155672
R2269 VTAIL.n706 VTAIL.n654 0.155672
R2270 VTAIL.n699 VTAIL.n654 0.155672
R2271 VTAIL.n699 VTAIL.n698 0.155672
R2272 VTAIL.n698 VTAIL.n658 0.155672
R2273 VTAIL.n691 VTAIL.n658 0.155672
R2274 VTAIL.n691 VTAIL.n690 0.155672
R2275 VTAIL.n690 VTAIL.n662 0.155672
R2276 VTAIL.n683 VTAIL.n662 0.155672
R2277 VTAIL.n683 VTAIL.n682 0.155672
R2278 VTAIL.n682 VTAIL.n666 0.155672
R2279 VTAIL.n675 VTAIL.n666 0.155672
R2280 VTAIL.n675 VTAIL.n674 0.155672
R2281 VTAIL.n633 VTAIL.n531 0.155672
R2282 VTAIL.n626 VTAIL.n531 0.155672
R2283 VTAIL.n626 VTAIL.n625 0.155672
R2284 VTAIL.n625 VTAIL.n535 0.155672
R2285 VTAIL.n618 VTAIL.n535 0.155672
R2286 VTAIL.n618 VTAIL.n617 0.155672
R2287 VTAIL.n617 VTAIL.n539 0.155672
R2288 VTAIL.n609 VTAIL.n539 0.155672
R2289 VTAIL.n609 VTAIL.n608 0.155672
R2290 VTAIL.n608 VTAIL.n543 0.155672
R2291 VTAIL.n601 VTAIL.n543 0.155672
R2292 VTAIL.n601 VTAIL.n600 0.155672
R2293 VTAIL.n600 VTAIL.n548 0.155672
R2294 VTAIL.n593 VTAIL.n548 0.155672
R2295 VTAIL.n593 VTAIL.n592 0.155672
R2296 VTAIL.n592 VTAIL.n552 0.155672
R2297 VTAIL.n585 VTAIL.n552 0.155672
R2298 VTAIL.n585 VTAIL.n584 0.155672
R2299 VTAIL.n584 VTAIL.n556 0.155672
R2300 VTAIL.n577 VTAIL.n556 0.155672
R2301 VTAIL.n577 VTAIL.n576 0.155672
R2302 VTAIL.n576 VTAIL.n560 0.155672
R2303 VTAIL.n569 VTAIL.n560 0.155672
R2304 VTAIL.n569 VTAIL.n568 0.155672
R2305 VTAIL.n527 VTAIL.n425 0.155672
R2306 VTAIL.n520 VTAIL.n425 0.155672
R2307 VTAIL.n520 VTAIL.n519 0.155672
R2308 VTAIL.n519 VTAIL.n429 0.155672
R2309 VTAIL.n512 VTAIL.n429 0.155672
R2310 VTAIL.n512 VTAIL.n511 0.155672
R2311 VTAIL.n511 VTAIL.n433 0.155672
R2312 VTAIL.n503 VTAIL.n433 0.155672
R2313 VTAIL.n503 VTAIL.n502 0.155672
R2314 VTAIL.n502 VTAIL.n437 0.155672
R2315 VTAIL.n495 VTAIL.n437 0.155672
R2316 VTAIL.n495 VTAIL.n494 0.155672
R2317 VTAIL.n494 VTAIL.n442 0.155672
R2318 VTAIL.n487 VTAIL.n442 0.155672
R2319 VTAIL.n487 VTAIL.n486 0.155672
R2320 VTAIL.n486 VTAIL.n446 0.155672
R2321 VTAIL.n479 VTAIL.n446 0.155672
R2322 VTAIL.n479 VTAIL.n478 0.155672
R2323 VTAIL.n478 VTAIL.n450 0.155672
R2324 VTAIL.n471 VTAIL.n450 0.155672
R2325 VTAIL.n471 VTAIL.n470 0.155672
R2326 VTAIL.n470 VTAIL.n454 0.155672
R2327 VTAIL.n463 VTAIL.n454 0.155672
R2328 VTAIL.n463 VTAIL.n462 0.155672
R2329 VTAIL.n421 VTAIL.n319 0.155672
R2330 VTAIL.n414 VTAIL.n319 0.155672
R2331 VTAIL.n414 VTAIL.n413 0.155672
R2332 VTAIL.n413 VTAIL.n323 0.155672
R2333 VTAIL.n406 VTAIL.n323 0.155672
R2334 VTAIL.n406 VTAIL.n405 0.155672
R2335 VTAIL.n405 VTAIL.n327 0.155672
R2336 VTAIL.n397 VTAIL.n327 0.155672
R2337 VTAIL.n397 VTAIL.n396 0.155672
R2338 VTAIL.n396 VTAIL.n331 0.155672
R2339 VTAIL.n389 VTAIL.n331 0.155672
R2340 VTAIL.n389 VTAIL.n388 0.155672
R2341 VTAIL.n388 VTAIL.n336 0.155672
R2342 VTAIL.n381 VTAIL.n336 0.155672
R2343 VTAIL.n381 VTAIL.n380 0.155672
R2344 VTAIL.n380 VTAIL.n340 0.155672
R2345 VTAIL.n373 VTAIL.n340 0.155672
R2346 VTAIL.n373 VTAIL.n372 0.155672
R2347 VTAIL.n372 VTAIL.n344 0.155672
R2348 VTAIL.n365 VTAIL.n344 0.155672
R2349 VTAIL.n365 VTAIL.n364 0.155672
R2350 VTAIL.n364 VTAIL.n348 0.155672
R2351 VTAIL.n357 VTAIL.n348 0.155672
R2352 VTAIL.n357 VTAIL.n356 0.155672
R2353 VDD2.n2 VDD2.n0 111.526
R2354 VDD2.n2 VDD2.n1 68.1908
R2355 VDD2.n1 VDD2.t2 1.7158
R2356 VDD2.n1 VDD2.t1 1.7158
R2357 VDD2.n0 VDD2.t0 1.7158
R2358 VDD2.n0 VDD2.t3 1.7158
R2359 VDD2 VDD2.n2 0.0586897
R2360 VP.n0 VP.t2 546.5
R2361 VP.n0 VP.t1 546.413
R2362 VP.n2 VP.t0 527.894
R2363 VP.n3 VP.t3 527.894
R2364 VP.n4 VP.n3 80.6037
R2365 VP.n2 VP.n1 80.6037
R2366 VP.n1 VP.n0 77.7001
R2367 VP.n3 VP.n2 48.2005
R2368 VP.n4 VP.n1 0.380177
R2369 VP VP.n4 0.146778
R2370 VDD1 VDD1.n1 112.052
R2371 VDD1 VDD1.n0 68.249
R2372 VDD1.n0 VDD1.t1 1.7158
R2373 VDD1.n0 VDD1.t2 1.7158
R2374 VDD1.n1 VDD1.t3 1.7158
R2375 VDD1.n1 VDD1.t0 1.7158
C0 VTAIL VDD1 8.80317f
C1 w_n1732_n4758# VDD2 1.32535f
C2 VTAIL VDD2 8.846251f
C3 VN VDD1 0.14761f
C4 VTAIL w_n1732_n4758# 5.80555f
C5 VN VDD2 5.47532f
C6 VN w_n1732_n4758# 2.76146f
C7 VN VTAIL 4.84898f
C8 B VP 1.22925f
C9 B VDD1 1.15597f
C10 B VDD2 1.18112f
C11 VP VDD1 5.61618f
C12 VP VDD2 0.288787f
C13 w_n1732_n4758# B 9.15164f
C14 VTAIL B 5.94966f
C15 w_n1732_n4758# VP 2.97992f
C16 VTAIL VP 4.86309f
C17 VDD1 VDD2 0.624375f
C18 VN B 0.874456f
C19 VN VP 6.28443f
C20 w_n1732_n4758# VDD1 1.30591f
C21 VDD2 VSUBS 0.875712f
C22 VDD1 VSUBS 5.961699f
C23 VTAIL VSUBS 1.239598f
C24 VN VSUBS 6.08092f
C25 VP VSUBS 1.695114f
C26 B VSUBS 3.423459f
C27 w_n1732_n4758# VSUBS 0.100698p
C28 VDD1.t1 VSUBS 0.409777f
C29 VDD1.t2 VSUBS 0.409777f
C30 VDD1.n0 VSUBS 3.42358f
C31 VDD1.t3 VSUBS 0.409777f
C32 VDD1.t0 VSUBS 0.409777f
C33 VDD1.n1 VSUBS 4.37998f
C34 VP.t1 VSUBS 2.65301f
C35 VP.t2 VSUBS 2.65318f
C36 VP.n0 VSUBS 3.50164f
C37 VP.n1 VSUBS 3.67949f
C38 VP.t0 VSUBS 2.61975f
C39 VP.n2 VSUBS 0.981331f
C40 VP.t3 VSUBS 2.61975f
C41 VP.n3 VSUBS 0.981331f
C42 VP.n4 VSUBS 0.065953f
C43 VDD2.t0 VSUBS 0.409808f
C44 VDD2.t3 VSUBS 0.409808f
C45 VDD2.n0 VSUBS 4.35213f
C46 VDD2.t2 VSUBS 0.409808f
C47 VDD2.t1 VSUBS 0.409808f
C48 VDD2.n1 VSUBS 3.42328f
C49 VDD2.n2 VSUBS 4.78293f
C50 VTAIL.n0 VSUBS 0.024134f
C51 VTAIL.n1 VSUBS 0.021795f
C52 VTAIL.n2 VSUBS 0.011712f
C53 VTAIL.n3 VSUBS 0.027682f
C54 VTAIL.n4 VSUBS 0.012401f
C55 VTAIL.n5 VSUBS 0.021795f
C56 VTAIL.n6 VSUBS 0.011712f
C57 VTAIL.n7 VSUBS 0.027682f
C58 VTAIL.n8 VSUBS 0.012401f
C59 VTAIL.n9 VSUBS 0.021795f
C60 VTAIL.n10 VSUBS 0.011712f
C61 VTAIL.n11 VSUBS 0.027682f
C62 VTAIL.n12 VSUBS 0.012401f
C63 VTAIL.n13 VSUBS 0.021795f
C64 VTAIL.n14 VSUBS 0.011712f
C65 VTAIL.n15 VSUBS 0.027682f
C66 VTAIL.n16 VSUBS 0.012401f
C67 VTAIL.n17 VSUBS 0.021795f
C68 VTAIL.n18 VSUBS 0.011712f
C69 VTAIL.n19 VSUBS 0.027682f
C70 VTAIL.n20 VSUBS 0.012401f
C71 VTAIL.n21 VSUBS 0.021795f
C72 VTAIL.n22 VSUBS 0.011712f
C73 VTAIL.n23 VSUBS 0.027682f
C74 VTAIL.n24 VSUBS 0.012401f
C75 VTAIL.n25 VSUBS 0.021795f
C76 VTAIL.n26 VSUBS 0.011712f
C77 VTAIL.n27 VSUBS 0.027682f
C78 VTAIL.n28 VSUBS 0.012401f
C79 VTAIL.n29 VSUBS 0.021795f
C80 VTAIL.n30 VSUBS 0.011712f
C81 VTAIL.n31 VSUBS 0.027682f
C82 VTAIL.n32 VSUBS 0.012401f
C83 VTAIL.n33 VSUBS 0.17903f
C84 VTAIL.t5 VSUBS 0.059476f
C85 VTAIL.n34 VSUBS 0.020762f
C86 VTAIL.n35 VSUBS 0.01761f
C87 VTAIL.n36 VSUBS 0.011712f
C88 VTAIL.n37 VSUBS 1.78249f
C89 VTAIL.n38 VSUBS 0.021795f
C90 VTAIL.n39 VSUBS 0.011712f
C91 VTAIL.n40 VSUBS 0.012401f
C92 VTAIL.n41 VSUBS 0.027682f
C93 VTAIL.n42 VSUBS 0.027682f
C94 VTAIL.n43 VSUBS 0.012401f
C95 VTAIL.n44 VSUBS 0.011712f
C96 VTAIL.n45 VSUBS 0.021795f
C97 VTAIL.n46 VSUBS 0.021795f
C98 VTAIL.n47 VSUBS 0.011712f
C99 VTAIL.n48 VSUBS 0.012401f
C100 VTAIL.n49 VSUBS 0.027682f
C101 VTAIL.n50 VSUBS 0.027682f
C102 VTAIL.n51 VSUBS 0.012401f
C103 VTAIL.n52 VSUBS 0.011712f
C104 VTAIL.n53 VSUBS 0.021795f
C105 VTAIL.n54 VSUBS 0.021795f
C106 VTAIL.n55 VSUBS 0.011712f
C107 VTAIL.n56 VSUBS 0.012401f
C108 VTAIL.n57 VSUBS 0.027682f
C109 VTAIL.n58 VSUBS 0.027682f
C110 VTAIL.n59 VSUBS 0.012401f
C111 VTAIL.n60 VSUBS 0.011712f
C112 VTAIL.n61 VSUBS 0.021795f
C113 VTAIL.n62 VSUBS 0.021795f
C114 VTAIL.n63 VSUBS 0.011712f
C115 VTAIL.n64 VSUBS 0.012401f
C116 VTAIL.n65 VSUBS 0.027682f
C117 VTAIL.n66 VSUBS 0.027682f
C118 VTAIL.n67 VSUBS 0.012401f
C119 VTAIL.n68 VSUBS 0.011712f
C120 VTAIL.n69 VSUBS 0.021795f
C121 VTAIL.n70 VSUBS 0.021795f
C122 VTAIL.n71 VSUBS 0.011712f
C123 VTAIL.n72 VSUBS 0.012401f
C124 VTAIL.n73 VSUBS 0.027682f
C125 VTAIL.n74 VSUBS 0.027682f
C126 VTAIL.n75 VSUBS 0.027682f
C127 VTAIL.n76 VSUBS 0.012401f
C128 VTAIL.n77 VSUBS 0.011712f
C129 VTAIL.n78 VSUBS 0.021795f
C130 VTAIL.n79 VSUBS 0.021795f
C131 VTAIL.n80 VSUBS 0.011712f
C132 VTAIL.n81 VSUBS 0.012056f
C133 VTAIL.n82 VSUBS 0.012056f
C134 VTAIL.n83 VSUBS 0.027682f
C135 VTAIL.n84 VSUBS 0.027682f
C136 VTAIL.n85 VSUBS 0.012401f
C137 VTAIL.n86 VSUBS 0.011712f
C138 VTAIL.n87 VSUBS 0.021795f
C139 VTAIL.n88 VSUBS 0.021795f
C140 VTAIL.n89 VSUBS 0.011712f
C141 VTAIL.n90 VSUBS 0.012401f
C142 VTAIL.n91 VSUBS 0.027682f
C143 VTAIL.n92 VSUBS 0.027682f
C144 VTAIL.n93 VSUBS 0.012401f
C145 VTAIL.n94 VSUBS 0.011712f
C146 VTAIL.n95 VSUBS 0.021795f
C147 VTAIL.n96 VSUBS 0.021795f
C148 VTAIL.n97 VSUBS 0.011712f
C149 VTAIL.n98 VSUBS 0.012401f
C150 VTAIL.n99 VSUBS 0.027682f
C151 VTAIL.n100 VSUBS 0.06765f
C152 VTAIL.n101 VSUBS 0.012401f
C153 VTAIL.n102 VSUBS 0.011712f
C154 VTAIL.n103 VSUBS 0.050081f
C155 VTAIL.n104 VSUBS 0.034039f
C156 VTAIL.n105 VSUBS 0.093973f
C157 VTAIL.n106 VSUBS 0.024134f
C158 VTAIL.n107 VSUBS 0.021795f
C159 VTAIL.n108 VSUBS 0.011712f
C160 VTAIL.n109 VSUBS 0.027682f
C161 VTAIL.n110 VSUBS 0.012401f
C162 VTAIL.n111 VSUBS 0.021795f
C163 VTAIL.n112 VSUBS 0.011712f
C164 VTAIL.n113 VSUBS 0.027682f
C165 VTAIL.n114 VSUBS 0.012401f
C166 VTAIL.n115 VSUBS 0.021795f
C167 VTAIL.n116 VSUBS 0.011712f
C168 VTAIL.n117 VSUBS 0.027682f
C169 VTAIL.n118 VSUBS 0.012401f
C170 VTAIL.n119 VSUBS 0.021795f
C171 VTAIL.n120 VSUBS 0.011712f
C172 VTAIL.n121 VSUBS 0.027682f
C173 VTAIL.n122 VSUBS 0.012401f
C174 VTAIL.n123 VSUBS 0.021795f
C175 VTAIL.n124 VSUBS 0.011712f
C176 VTAIL.n125 VSUBS 0.027682f
C177 VTAIL.n126 VSUBS 0.012401f
C178 VTAIL.n127 VSUBS 0.021795f
C179 VTAIL.n128 VSUBS 0.011712f
C180 VTAIL.n129 VSUBS 0.027682f
C181 VTAIL.n130 VSUBS 0.012401f
C182 VTAIL.n131 VSUBS 0.021795f
C183 VTAIL.n132 VSUBS 0.011712f
C184 VTAIL.n133 VSUBS 0.027682f
C185 VTAIL.n134 VSUBS 0.012401f
C186 VTAIL.n135 VSUBS 0.021795f
C187 VTAIL.n136 VSUBS 0.011712f
C188 VTAIL.n137 VSUBS 0.027682f
C189 VTAIL.n138 VSUBS 0.012401f
C190 VTAIL.n139 VSUBS 0.17903f
C191 VTAIL.t3 VSUBS 0.059476f
C192 VTAIL.n140 VSUBS 0.020762f
C193 VTAIL.n141 VSUBS 0.01761f
C194 VTAIL.n142 VSUBS 0.011712f
C195 VTAIL.n143 VSUBS 1.78249f
C196 VTAIL.n144 VSUBS 0.021795f
C197 VTAIL.n145 VSUBS 0.011712f
C198 VTAIL.n146 VSUBS 0.012401f
C199 VTAIL.n147 VSUBS 0.027682f
C200 VTAIL.n148 VSUBS 0.027682f
C201 VTAIL.n149 VSUBS 0.012401f
C202 VTAIL.n150 VSUBS 0.011712f
C203 VTAIL.n151 VSUBS 0.021795f
C204 VTAIL.n152 VSUBS 0.021795f
C205 VTAIL.n153 VSUBS 0.011712f
C206 VTAIL.n154 VSUBS 0.012401f
C207 VTAIL.n155 VSUBS 0.027682f
C208 VTAIL.n156 VSUBS 0.027682f
C209 VTAIL.n157 VSUBS 0.012401f
C210 VTAIL.n158 VSUBS 0.011712f
C211 VTAIL.n159 VSUBS 0.021795f
C212 VTAIL.n160 VSUBS 0.021795f
C213 VTAIL.n161 VSUBS 0.011712f
C214 VTAIL.n162 VSUBS 0.012401f
C215 VTAIL.n163 VSUBS 0.027682f
C216 VTAIL.n164 VSUBS 0.027682f
C217 VTAIL.n165 VSUBS 0.012401f
C218 VTAIL.n166 VSUBS 0.011712f
C219 VTAIL.n167 VSUBS 0.021795f
C220 VTAIL.n168 VSUBS 0.021795f
C221 VTAIL.n169 VSUBS 0.011712f
C222 VTAIL.n170 VSUBS 0.012401f
C223 VTAIL.n171 VSUBS 0.027682f
C224 VTAIL.n172 VSUBS 0.027682f
C225 VTAIL.n173 VSUBS 0.012401f
C226 VTAIL.n174 VSUBS 0.011712f
C227 VTAIL.n175 VSUBS 0.021795f
C228 VTAIL.n176 VSUBS 0.021795f
C229 VTAIL.n177 VSUBS 0.011712f
C230 VTAIL.n178 VSUBS 0.012401f
C231 VTAIL.n179 VSUBS 0.027682f
C232 VTAIL.n180 VSUBS 0.027682f
C233 VTAIL.n181 VSUBS 0.027682f
C234 VTAIL.n182 VSUBS 0.012401f
C235 VTAIL.n183 VSUBS 0.011712f
C236 VTAIL.n184 VSUBS 0.021795f
C237 VTAIL.n185 VSUBS 0.021795f
C238 VTAIL.n186 VSUBS 0.011712f
C239 VTAIL.n187 VSUBS 0.012056f
C240 VTAIL.n188 VSUBS 0.012056f
C241 VTAIL.n189 VSUBS 0.027682f
C242 VTAIL.n190 VSUBS 0.027682f
C243 VTAIL.n191 VSUBS 0.012401f
C244 VTAIL.n192 VSUBS 0.011712f
C245 VTAIL.n193 VSUBS 0.021795f
C246 VTAIL.n194 VSUBS 0.021795f
C247 VTAIL.n195 VSUBS 0.011712f
C248 VTAIL.n196 VSUBS 0.012401f
C249 VTAIL.n197 VSUBS 0.027682f
C250 VTAIL.n198 VSUBS 0.027682f
C251 VTAIL.n199 VSUBS 0.012401f
C252 VTAIL.n200 VSUBS 0.011712f
C253 VTAIL.n201 VSUBS 0.021795f
C254 VTAIL.n202 VSUBS 0.021795f
C255 VTAIL.n203 VSUBS 0.011712f
C256 VTAIL.n204 VSUBS 0.012401f
C257 VTAIL.n205 VSUBS 0.027682f
C258 VTAIL.n206 VSUBS 0.06765f
C259 VTAIL.n207 VSUBS 0.012401f
C260 VTAIL.n208 VSUBS 0.011712f
C261 VTAIL.n209 VSUBS 0.050081f
C262 VTAIL.n210 VSUBS 0.034039f
C263 VTAIL.n211 VSUBS 0.12833f
C264 VTAIL.n212 VSUBS 0.024134f
C265 VTAIL.n213 VSUBS 0.021795f
C266 VTAIL.n214 VSUBS 0.011712f
C267 VTAIL.n215 VSUBS 0.027682f
C268 VTAIL.n216 VSUBS 0.012401f
C269 VTAIL.n217 VSUBS 0.021795f
C270 VTAIL.n218 VSUBS 0.011712f
C271 VTAIL.n219 VSUBS 0.027682f
C272 VTAIL.n220 VSUBS 0.012401f
C273 VTAIL.n221 VSUBS 0.021795f
C274 VTAIL.n222 VSUBS 0.011712f
C275 VTAIL.n223 VSUBS 0.027682f
C276 VTAIL.n224 VSUBS 0.012401f
C277 VTAIL.n225 VSUBS 0.021795f
C278 VTAIL.n226 VSUBS 0.011712f
C279 VTAIL.n227 VSUBS 0.027682f
C280 VTAIL.n228 VSUBS 0.012401f
C281 VTAIL.n229 VSUBS 0.021795f
C282 VTAIL.n230 VSUBS 0.011712f
C283 VTAIL.n231 VSUBS 0.027682f
C284 VTAIL.n232 VSUBS 0.012401f
C285 VTAIL.n233 VSUBS 0.021795f
C286 VTAIL.n234 VSUBS 0.011712f
C287 VTAIL.n235 VSUBS 0.027682f
C288 VTAIL.n236 VSUBS 0.012401f
C289 VTAIL.n237 VSUBS 0.021795f
C290 VTAIL.n238 VSUBS 0.011712f
C291 VTAIL.n239 VSUBS 0.027682f
C292 VTAIL.n240 VSUBS 0.012401f
C293 VTAIL.n241 VSUBS 0.021795f
C294 VTAIL.n242 VSUBS 0.011712f
C295 VTAIL.n243 VSUBS 0.027682f
C296 VTAIL.n244 VSUBS 0.012401f
C297 VTAIL.n245 VSUBS 0.17903f
C298 VTAIL.t1 VSUBS 0.059476f
C299 VTAIL.n246 VSUBS 0.020762f
C300 VTAIL.n247 VSUBS 0.01761f
C301 VTAIL.n248 VSUBS 0.011712f
C302 VTAIL.n249 VSUBS 1.78249f
C303 VTAIL.n250 VSUBS 0.021795f
C304 VTAIL.n251 VSUBS 0.011712f
C305 VTAIL.n252 VSUBS 0.012401f
C306 VTAIL.n253 VSUBS 0.027682f
C307 VTAIL.n254 VSUBS 0.027682f
C308 VTAIL.n255 VSUBS 0.012401f
C309 VTAIL.n256 VSUBS 0.011712f
C310 VTAIL.n257 VSUBS 0.021795f
C311 VTAIL.n258 VSUBS 0.021795f
C312 VTAIL.n259 VSUBS 0.011712f
C313 VTAIL.n260 VSUBS 0.012401f
C314 VTAIL.n261 VSUBS 0.027682f
C315 VTAIL.n262 VSUBS 0.027682f
C316 VTAIL.n263 VSUBS 0.012401f
C317 VTAIL.n264 VSUBS 0.011712f
C318 VTAIL.n265 VSUBS 0.021795f
C319 VTAIL.n266 VSUBS 0.021795f
C320 VTAIL.n267 VSUBS 0.011712f
C321 VTAIL.n268 VSUBS 0.012401f
C322 VTAIL.n269 VSUBS 0.027682f
C323 VTAIL.n270 VSUBS 0.027682f
C324 VTAIL.n271 VSUBS 0.012401f
C325 VTAIL.n272 VSUBS 0.011712f
C326 VTAIL.n273 VSUBS 0.021795f
C327 VTAIL.n274 VSUBS 0.021795f
C328 VTAIL.n275 VSUBS 0.011712f
C329 VTAIL.n276 VSUBS 0.012401f
C330 VTAIL.n277 VSUBS 0.027682f
C331 VTAIL.n278 VSUBS 0.027682f
C332 VTAIL.n279 VSUBS 0.012401f
C333 VTAIL.n280 VSUBS 0.011712f
C334 VTAIL.n281 VSUBS 0.021795f
C335 VTAIL.n282 VSUBS 0.021795f
C336 VTAIL.n283 VSUBS 0.011712f
C337 VTAIL.n284 VSUBS 0.012401f
C338 VTAIL.n285 VSUBS 0.027682f
C339 VTAIL.n286 VSUBS 0.027682f
C340 VTAIL.n287 VSUBS 0.027682f
C341 VTAIL.n288 VSUBS 0.012401f
C342 VTAIL.n289 VSUBS 0.011712f
C343 VTAIL.n290 VSUBS 0.021795f
C344 VTAIL.n291 VSUBS 0.021795f
C345 VTAIL.n292 VSUBS 0.011712f
C346 VTAIL.n293 VSUBS 0.012056f
C347 VTAIL.n294 VSUBS 0.012056f
C348 VTAIL.n295 VSUBS 0.027682f
C349 VTAIL.n296 VSUBS 0.027682f
C350 VTAIL.n297 VSUBS 0.012401f
C351 VTAIL.n298 VSUBS 0.011712f
C352 VTAIL.n299 VSUBS 0.021795f
C353 VTAIL.n300 VSUBS 0.021795f
C354 VTAIL.n301 VSUBS 0.011712f
C355 VTAIL.n302 VSUBS 0.012401f
C356 VTAIL.n303 VSUBS 0.027682f
C357 VTAIL.n304 VSUBS 0.027682f
C358 VTAIL.n305 VSUBS 0.012401f
C359 VTAIL.n306 VSUBS 0.011712f
C360 VTAIL.n307 VSUBS 0.021795f
C361 VTAIL.n308 VSUBS 0.021795f
C362 VTAIL.n309 VSUBS 0.011712f
C363 VTAIL.n310 VSUBS 0.012401f
C364 VTAIL.n311 VSUBS 0.027682f
C365 VTAIL.n312 VSUBS 0.06765f
C366 VTAIL.n313 VSUBS 0.012401f
C367 VTAIL.n314 VSUBS 0.011712f
C368 VTAIL.n315 VSUBS 0.050081f
C369 VTAIL.n316 VSUBS 0.034039f
C370 VTAIL.n317 VSUBS 1.61556f
C371 VTAIL.n318 VSUBS 0.024134f
C372 VTAIL.n319 VSUBS 0.021795f
C373 VTAIL.n320 VSUBS 0.011712f
C374 VTAIL.n321 VSUBS 0.027682f
C375 VTAIL.n322 VSUBS 0.012401f
C376 VTAIL.n323 VSUBS 0.021795f
C377 VTAIL.n324 VSUBS 0.011712f
C378 VTAIL.n325 VSUBS 0.027682f
C379 VTAIL.n326 VSUBS 0.012401f
C380 VTAIL.n327 VSUBS 0.021795f
C381 VTAIL.n328 VSUBS 0.011712f
C382 VTAIL.n329 VSUBS 0.027682f
C383 VTAIL.n330 VSUBS 0.012401f
C384 VTAIL.n331 VSUBS 0.021795f
C385 VTAIL.n332 VSUBS 0.011712f
C386 VTAIL.n333 VSUBS 0.027682f
C387 VTAIL.n334 VSUBS 0.027682f
C388 VTAIL.n335 VSUBS 0.012401f
C389 VTAIL.n336 VSUBS 0.021795f
C390 VTAIL.n337 VSUBS 0.011712f
C391 VTAIL.n338 VSUBS 0.027682f
C392 VTAIL.n339 VSUBS 0.012401f
C393 VTAIL.n340 VSUBS 0.021795f
C394 VTAIL.n341 VSUBS 0.011712f
C395 VTAIL.n342 VSUBS 0.027682f
C396 VTAIL.n343 VSUBS 0.012401f
C397 VTAIL.n344 VSUBS 0.021795f
C398 VTAIL.n345 VSUBS 0.011712f
C399 VTAIL.n346 VSUBS 0.027682f
C400 VTAIL.n347 VSUBS 0.012401f
C401 VTAIL.n348 VSUBS 0.021795f
C402 VTAIL.n349 VSUBS 0.011712f
C403 VTAIL.n350 VSUBS 0.027682f
C404 VTAIL.n351 VSUBS 0.012401f
C405 VTAIL.n352 VSUBS 0.17903f
C406 VTAIL.t4 VSUBS 0.059476f
C407 VTAIL.n353 VSUBS 0.020762f
C408 VTAIL.n354 VSUBS 0.01761f
C409 VTAIL.n355 VSUBS 0.011712f
C410 VTAIL.n356 VSUBS 1.78249f
C411 VTAIL.n357 VSUBS 0.021795f
C412 VTAIL.n358 VSUBS 0.011712f
C413 VTAIL.n359 VSUBS 0.012401f
C414 VTAIL.n360 VSUBS 0.027682f
C415 VTAIL.n361 VSUBS 0.027682f
C416 VTAIL.n362 VSUBS 0.012401f
C417 VTAIL.n363 VSUBS 0.011712f
C418 VTAIL.n364 VSUBS 0.021795f
C419 VTAIL.n365 VSUBS 0.021795f
C420 VTAIL.n366 VSUBS 0.011712f
C421 VTAIL.n367 VSUBS 0.012401f
C422 VTAIL.n368 VSUBS 0.027682f
C423 VTAIL.n369 VSUBS 0.027682f
C424 VTAIL.n370 VSUBS 0.012401f
C425 VTAIL.n371 VSUBS 0.011712f
C426 VTAIL.n372 VSUBS 0.021795f
C427 VTAIL.n373 VSUBS 0.021795f
C428 VTAIL.n374 VSUBS 0.011712f
C429 VTAIL.n375 VSUBS 0.012401f
C430 VTAIL.n376 VSUBS 0.027682f
C431 VTAIL.n377 VSUBS 0.027682f
C432 VTAIL.n378 VSUBS 0.012401f
C433 VTAIL.n379 VSUBS 0.011712f
C434 VTAIL.n380 VSUBS 0.021795f
C435 VTAIL.n381 VSUBS 0.021795f
C436 VTAIL.n382 VSUBS 0.011712f
C437 VTAIL.n383 VSUBS 0.012401f
C438 VTAIL.n384 VSUBS 0.027682f
C439 VTAIL.n385 VSUBS 0.027682f
C440 VTAIL.n386 VSUBS 0.012401f
C441 VTAIL.n387 VSUBS 0.011712f
C442 VTAIL.n388 VSUBS 0.021795f
C443 VTAIL.n389 VSUBS 0.021795f
C444 VTAIL.n390 VSUBS 0.011712f
C445 VTAIL.n391 VSUBS 0.012401f
C446 VTAIL.n392 VSUBS 0.027682f
C447 VTAIL.n393 VSUBS 0.027682f
C448 VTAIL.n394 VSUBS 0.012401f
C449 VTAIL.n395 VSUBS 0.011712f
C450 VTAIL.n396 VSUBS 0.021795f
C451 VTAIL.n397 VSUBS 0.021795f
C452 VTAIL.n398 VSUBS 0.011712f
C453 VTAIL.n399 VSUBS 0.012056f
C454 VTAIL.n400 VSUBS 0.012056f
C455 VTAIL.n401 VSUBS 0.027682f
C456 VTAIL.n402 VSUBS 0.027682f
C457 VTAIL.n403 VSUBS 0.012401f
C458 VTAIL.n404 VSUBS 0.011712f
C459 VTAIL.n405 VSUBS 0.021795f
C460 VTAIL.n406 VSUBS 0.021795f
C461 VTAIL.n407 VSUBS 0.011712f
C462 VTAIL.n408 VSUBS 0.012401f
C463 VTAIL.n409 VSUBS 0.027682f
C464 VTAIL.n410 VSUBS 0.027682f
C465 VTAIL.n411 VSUBS 0.012401f
C466 VTAIL.n412 VSUBS 0.011712f
C467 VTAIL.n413 VSUBS 0.021795f
C468 VTAIL.n414 VSUBS 0.021795f
C469 VTAIL.n415 VSUBS 0.011712f
C470 VTAIL.n416 VSUBS 0.012401f
C471 VTAIL.n417 VSUBS 0.027682f
C472 VTAIL.n418 VSUBS 0.06765f
C473 VTAIL.n419 VSUBS 0.012401f
C474 VTAIL.n420 VSUBS 0.011712f
C475 VTAIL.n421 VSUBS 0.050081f
C476 VTAIL.n422 VSUBS 0.034039f
C477 VTAIL.n423 VSUBS 1.61556f
C478 VTAIL.n424 VSUBS 0.024134f
C479 VTAIL.n425 VSUBS 0.021795f
C480 VTAIL.n426 VSUBS 0.011712f
C481 VTAIL.n427 VSUBS 0.027682f
C482 VTAIL.n428 VSUBS 0.012401f
C483 VTAIL.n429 VSUBS 0.021795f
C484 VTAIL.n430 VSUBS 0.011712f
C485 VTAIL.n431 VSUBS 0.027682f
C486 VTAIL.n432 VSUBS 0.012401f
C487 VTAIL.n433 VSUBS 0.021795f
C488 VTAIL.n434 VSUBS 0.011712f
C489 VTAIL.n435 VSUBS 0.027682f
C490 VTAIL.n436 VSUBS 0.012401f
C491 VTAIL.n437 VSUBS 0.021795f
C492 VTAIL.n438 VSUBS 0.011712f
C493 VTAIL.n439 VSUBS 0.027682f
C494 VTAIL.n440 VSUBS 0.027682f
C495 VTAIL.n441 VSUBS 0.012401f
C496 VTAIL.n442 VSUBS 0.021795f
C497 VTAIL.n443 VSUBS 0.011712f
C498 VTAIL.n444 VSUBS 0.027682f
C499 VTAIL.n445 VSUBS 0.012401f
C500 VTAIL.n446 VSUBS 0.021795f
C501 VTAIL.n447 VSUBS 0.011712f
C502 VTAIL.n448 VSUBS 0.027682f
C503 VTAIL.n449 VSUBS 0.012401f
C504 VTAIL.n450 VSUBS 0.021795f
C505 VTAIL.n451 VSUBS 0.011712f
C506 VTAIL.n452 VSUBS 0.027682f
C507 VTAIL.n453 VSUBS 0.012401f
C508 VTAIL.n454 VSUBS 0.021795f
C509 VTAIL.n455 VSUBS 0.011712f
C510 VTAIL.n456 VSUBS 0.027682f
C511 VTAIL.n457 VSUBS 0.012401f
C512 VTAIL.n458 VSUBS 0.17903f
C513 VTAIL.t7 VSUBS 0.059476f
C514 VTAIL.n459 VSUBS 0.020762f
C515 VTAIL.n460 VSUBS 0.01761f
C516 VTAIL.n461 VSUBS 0.011712f
C517 VTAIL.n462 VSUBS 1.78249f
C518 VTAIL.n463 VSUBS 0.021795f
C519 VTAIL.n464 VSUBS 0.011712f
C520 VTAIL.n465 VSUBS 0.012401f
C521 VTAIL.n466 VSUBS 0.027682f
C522 VTAIL.n467 VSUBS 0.027682f
C523 VTAIL.n468 VSUBS 0.012401f
C524 VTAIL.n469 VSUBS 0.011712f
C525 VTAIL.n470 VSUBS 0.021795f
C526 VTAIL.n471 VSUBS 0.021795f
C527 VTAIL.n472 VSUBS 0.011712f
C528 VTAIL.n473 VSUBS 0.012401f
C529 VTAIL.n474 VSUBS 0.027682f
C530 VTAIL.n475 VSUBS 0.027682f
C531 VTAIL.n476 VSUBS 0.012401f
C532 VTAIL.n477 VSUBS 0.011712f
C533 VTAIL.n478 VSUBS 0.021795f
C534 VTAIL.n479 VSUBS 0.021795f
C535 VTAIL.n480 VSUBS 0.011712f
C536 VTAIL.n481 VSUBS 0.012401f
C537 VTAIL.n482 VSUBS 0.027682f
C538 VTAIL.n483 VSUBS 0.027682f
C539 VTAIL.n484 VSUBS 0.012401f
C540 VTAIL.n485 VSUBS 0.011712f
C541 VTAIL.n486 VSUBS 0.021795f
C542 VTAIL.n487 VSUBS 0.021795f
C543 VTAIL.n488 VSUBS 0.011712f
C544 VTAIL.n489 VSUBS 0.012401f
C545 VTAIL.n490 VSUBS 0.027682f
C546 VTAIL.n491 VSUBS 0.027682f
C547 VTAIL.n492 VSUBS 0.012401f
C548 VTAIL.n493 VSUBS 0.011712f
C549 VTAIL.n494 VSUBS 0.021795f
C550 VTAIL.n495 VSUBS 0.021795f
C551 VTAIL.n496 VSUBS 0.011712f
C552 VTAIL.n497 VSUBS 0.012401f
C553 VTAIL.n498 VSUBS 0.027682f
C554 VTAIL.n499 VSUBS 0.027682f
C555 VTAIL.n500 VSUBS 0.012401f
C556 VTAIL.n501 VSUBS 0.011712f
C557 VTAIL.n502 VSUBS 0.021795f
C558 VTAIL.n503 VSUBS 0.021795f
C559 VTAIL.n504 VSUBS 0.011712f
C560 VTAIL.n505 VSUBS 0.012056f
C561 VTAIL.n506 VSUBS 0.012056f
C562 VTAIL.n507 VSUBS 0.027682f
C563 VTAIL.n508 VSUBS 0.027682f
C564 VTAIL.n509 VSUBS 0.012401f
C565 VTAIL.n510 VSUBS 0.011712f
C566 VTAIL.n511 VSUBS 0.021795f
C567 VTAIL.n512 VSUBS 0.021795f
C568 VTAIL.n513 VSUBS 0.011712f
C569 VTAIL.n514 VSUBS 0.012401f
C570 VTAIL.n515 VSUBS 0.027682f
C571 VTAIL.n516 VSUBS 0.027682f
C572 VTAIL.n517 VSUBS 0.012401f
C573 VTAIL.n518 VSUBS 0.011712f
C574 VTAIL.n519 VSUBS 0.021795f
C575 VTAIL.n520 VSUBS 0.021795f
C576 VTAIL.n521 VSUBS 0.011712f
C577 VTAIL.n522 VSUBS 0.012401f
C578 VTAIL.n523 VSUBS 0.027682f
C579 VTAIL.n524 VSUBS 0.06765f
C580 VTAIL.n525 VSUBS 0.012401f
C581 VTAIL.n526 VSUBS 0.011712f
C582 VTAIL.n527 VSUBS 0.050081f
C583 VTAIL.n528 VSUBS 0.034039f
C584 VTAIL.n529 VSUBS 0.12833f
C585 VTAIL.n530 VSUBS 0.024134f
C586 VTAIL.n531 VSUBS 0.021795f
C587 VTAIL.n532 VSUBS 0.011712f
C588 VTAIL.n533 VSUBS 0.027682f
C589 VTAIL.n534 VSUBS 0.012401f
C590 VTAIL.n535 VSUBS 0.021795f
C591 VTAIL.n536 VSUBS 0.011712f
C592 VTAIL.n537 VSUBS 0.027682f
C593 VTAIL.n538 VSUBS 0.012401f
C594 VTAIL.n539 VSUBS 0.021795f
C595 VTAIL.n540 VSUBS 0.011712f
C596 VTAIL.n541 VSUBS 0.027682f
C597 VTAIL.n542 VSUBS 0.012401f
C598 VTAIL.n543 VSUBS 0.021795f
C599 VTAIL.n544 VSUBS 0.011712f
C600 VTAIL.n545 VSUBS 0.027682f
C601 VTAIL.n546 VSUBS 0.027682f
C602 VTAIL.n547 VSUBS 0.012401f
C603 VTAIL.n548 VSUBS 0.021795f
C604 VTAIL.n549 VSUBS 0.011712f
C605 VTAIL.n550 VSUBS 0.027682f
C606 VTAIL.n551 VSUBS 0.012401f
C607 VTAIL.n552 VSUBS 0.021795f
C608 VTAIL.n553 VSUBS 0.011712f
C609 VTAIL.n554 VSUBS 0.027682f
C610 VTAIL.n555 VSUBS 0.012401f
C611 VTAIL.n556 VSUBS 0.021795f
C612 VTAIL.n557 VSUBS 0.011712f
C613 VTAIL.n558 VSUBS 0.027682f
C614 VTAIL.n559 VSUBS 0.012401f
C615 VTAIL.n560 VSUBS 0.021795f
C616 VTAIL.n561 VSUBS 0.011712f
C617 VTAIL.n562 VSUBS 0.027682f
C618 VTAIL.n563 VSUBS 0.012401f
C619 VTAIL.n564 VSUBS 0.17903f
C620 VTAIL.t0 VSUBS 0.059476f
C621 VTAIL.n565 VSUBS 0.020762f
C622 VTAIL.n566 VSUBS 0.01761f
C623 VTAIL.n567 VSUBS 0.011712f
C624 VTAIL.n568 VSUBS 1.78249f
C625 VTAIL.n569 VSUBS 0.021795f
C626 VTAIL.n570 VSUBS 0.011712f
C627 VTAIL.n571 VSUBS 0.012401f
C628 VTAIL.n572 VSUBS 0.027682f
C629 VTAIL.n573 VSUBS 0.027682f
C630 VTAIL.n574 VSUBS 0.012401f
C631 VTAIL.n575 VSUBS 0.011712f
C632 VTAIL.n576 VSUBS 0.021795f
C633 VTAIL.n577 VSUBS 0.021795f
C634 VTAIL.n578 VSUBS 0.011712f
C635 VTAIL.n579 VSUBS 0.012401f
C636 VTAIL.n580 VSUBS 0.027682f
C637 VTAIL.n581 VSUBS 0.027682f
C638 VTAIL.n582 VSUBS 0.012401f
C639 VTAIL.n583 VSUBS 0.011712f
C640 VTAIL.n584 VSUBS 0.021795f
C641 VTAIL.n585 VSUBS 0.021795f
C642 VTAIL.n586 VSUBS 0.011712f
C643 VTAIL.n587 VSUBS 0.012401f
C644 VTAIL.n588 VSUBS 0.027682f
C645 VTAIL.n589 VSUBS 0.027682f
C646 VTAIL.n590 VSUBS 0.012401f
C647 VTAIL.n591 VSUBS 0.011712f
C648 VTAIL.n592 VSUBS 0.021795f
C649 VTAIL.n593 VSUBS 0.021795f
C650 VTAIL.n594 VSUBS 0.011712f
C651 VTAIL.n595 VSUBS 0.012401f
C652 VTAIL.n596 VSUBS 0.027682f
C653 VTAIL.n597 VSUBS 0.027682f
C654 VTAIL.n598 VSUBS 0.012401f
C655 VTAIL.n599 VSUBS 0.011712f
C656 VTAIL.n600 VSUBS 0.021795f
C657 VTAIL.n601 VSUBS 0.021795f
C658 VTAIL.n602 VSUBS 0.011712f
C659 VTAIL.n603 VSUBS 0.012401f
C660 VTAIL.n604 VSUBS 0.027682f
C661 VTAIL.n605 VSUBS 0.027682f
C662 VTAIL.n606 VSUBS 0.012401f
C663 VTAIL.n607 VSUBS 0.011712f
C664 VTAIL.n608 VSUBS 0.021795f
C665 VTAIL.n609 VSUBS 0.021795f
C666 VTAIL.n610 VSUBS 0.011712f
C667 VTAIL.n611 VSUBS 0.012056f
C668 VTAIL.n612 VSUBS 0.012056f
C669 VTAIL.n613 VSUBS 0.027682f
C670 VTAIL.n614 VSUBS 0.027682f
C671 VTAIL.n615 VSUBS 0.012401f
C672 VTAIL.n616 VSUBS 0.011712f
C673 VTAIL.n617 VSUBS 0.021795f
C674 VTAIL.n618 VSUBS 0.021795f
C675 VTAIL.n619 VSUBS 0.011712f
C676 VTAIL.n620 VSUBS 0.012401f
C677 VTAIL.n621 VSUBS 0.027682f
C678 VTAIL.n622 VSUBS 0.027682f
C679 VTAIL.n623 VSUBS 0.012401f
C680 VTAIL.n624 VSUBS 0.011712f
C681 VTAIL.n625 VSUBS 0.021795f
C682 VTAIL.n626 VSUBS 0.021795f
C683 VTAIL.n627 VSUBS 0.011712f
C684 VTAIL.n628 VSUBS 0.012401f
C685 VTAIL.n629 VSUBS 0.027682f
C686 VTAIL.n630 VSUBS 0.06765f
C687 VTAIL.n631 VSUBS 0.012401f
C688 VTAIL.n632 VSUBS 0.011712f
C689 VTAIL.n633 VSUBS 0.050081f
C690 VTAIL.n634 VSUBS 0.034039f
C691 VTAIL.n635 VSUBS 0.12833f
C692 VTAIL.n636 VSUBS 0.024134f
C693 VTAIL.n637 VSUBS 0.021795f
C694 VTAIL.n638 VSUBS 0.011712f
C695 VTAIL.n639 VSUBS 0.027682f
C696 VTAIL.n640 VSUBS 0.012401f
C697 VTAIL.n641 VSUBS 0.021795f
C698 VTAIL.n642 VSUBS 0.011712f
C699 VTAIL.n643 VSUBS 0.027682f
C700 VTAIL.n644 VSUBS 0.012401f
C701 VTAIL.n645 VSUBS 0.021795f
C702 VTAIL.n646 VSUBS 0.011712f
C703 VTAIL.n647 VSUBS 0.027682f
C704 VTAIL.n648 VSUBS 0.012401f
C705 VTAIL.n649 VSUBS 0.021795f
C706 VTAIL.n650 VSUBS 0.011712f
C707 VTAIL.n651 VSUBS 0.027682f
C708 VTAIL.n652 VSUBS 0.027682f
C709 VTAIL.n653 VSUBS 0.012401f
C710 VTAIL.n654 VSUBS 0.021795f
C711 VTAIL.n655 VSUBS 0.011712f
C712 VTAIL.n656 VSUBS 0.027682f
C713 VTAIL.n657 VSUBS 0.012401f
C714 VTAIL.n658 VSUBS 0.021795f
C715 VTAIL.n659 VSUBS 0.011712f
C716 VTAIL.n660 VSUBS 0.027682f
C717 VTAIL.n661 VSUBS 0.012401f
C718 VTAIL.n662 VSUBS 0.021795f
C719 VTAIL.n663 VSUBS 0.011712f
C720 VTAIL.n664 VSUBS 0.027682f
C721 VTAIL.n665 VSUBS 0.012401f
C722 VTAIL.n666 VSUBS 0.021795f
C723 VTAIL.n667 VSUBS 0.011712f
C724 VTAIL.n668 VSUBS 0.027682f
C725 VTAIL.n669 VSUBS 0.012401f
C726 VTAIL.n670 VSUBS 0.17903f
C727 VTAIL.t2 VSUBS 0.059476f
C728 VTAIL.n671 VSUBS 0.020762f
C729 VTAIL.n672 VSUBS 0.01761f
C730 VTAIL.n673 VSUBS 0.011712f
C731 VTAIL.n674 VSUBS 1.78249f
C732 VTAIL.n675 VSUBS 0.021795f
C733 VTAIL.n676 VSUBS 0.011712f
C734 VTAIL.n677 VSUBS 0.012401f
C735 VTAIL.n678 VSUBS 0.027682f
C736 VTAIL.n679 VSUBS 0.027682f
C737 VTAIL.n680 VSUBS 0.012401f
C738 VTAIL.n681 VSUBS 0.011712f
C739 VTAIL.n682 VSUBS 0.021795f
C740 VTAIL.n683 VSUBS 0.021795f
C741 VTAIL.n684 VSUBS 0.011712f
C742 VTAIL.n685 VSUBS 0.012401f
C743 VTAIL.n686 VSUBS 0.027682f
C744 VTAIL.n687 VSUBS 0.027682f
C745 VTAIL.n688 VSUBS 0.012401f
C746 VTAIL.n689 VSUBS 0.011712f
C747 VTAIL.n690 VSUBS 0.021795f
C748 VTAIL.n691 VSUBS 0.021795f
C749 VTAIL.n692 VSUBS 0.011712f
C750 VTAIL.n693 VSUBS 0.012401f
C751 VTAIL.n694 VSUBS 0.027682f
C752 VTAIL.n695 VSUBS 0.027682f
C753 VTAIL.n696 VSUBS 0.012401f
C754 VTAIL.n697 VSUBS 0.011712f
C755 VTAIL.n698 VSUBS 0.021795f
C756 VTAIL.n699 VSUBS 0.021795f
C757 VTAIL.n700 VSUBS 0.011712f
C758 VTAIL.n701 VSUBS 0.012401f
C759 VTAIL.n702 VSUBS 0.027682f
C760 VTAIL.n703 VSUBS 0.027682f
C761 VTAIL.n704 VSUBS 0.012401f
C762 VTAIL.n705 VSUBS 0.011712f
C763 VTAIL.n706 VSUBS 0.021795f
C764 VTAIL.n707 VSUBS 0.021795f
C765 VTAIL.n708 VSUBS 0.011712f
C766 VTAIL.n709 VSUBS 0.012401f
C767 VTAIL.n710 VSUBS 0.027682f
C768 VTAIL.n711 VSUBS 0.027682f
C769 VTAIL.n712 VSUBS 0.012401f
C770 VTAIL.n713 VSUBS 0.011712f
C771 VTAIL.n714 VSUBS 0.021795f
C772 VTAIL.n715 VSUBS 0.021795f
C773 VTAIL.n716 VSUBS 0.011712f
C774 VTAIL.n717 VSUBS 0.012056f
C775 VTAIL.n718 VSUBS 0.012056f
C776 VTAIL.n719 VSUBS 0.027682f
C777 VTAIL.n720 VSUBS 0.027682f
C778 VTAIL.n721 VSUBS 0.012401f
C779 VTAIL.n722 VSUBS 0.011712f
C780 VTAIL.n723 VSUBS 0.021795f
C781 VTAIL.n724 VSUBS 0.021795f
C782 VTAIL.n725 VSUBS 0.011712f
C783 VTAIL.n726 VSUBS 0.012401f
C784 VTAIL.n727 VSUBS 0.027682f
C785 VTAIL.n728 VSUBS 0.027682f
C786 VTAIL.n729 VSUBS 0.012401f
C787 VTAIL.n730 VSUBS 0.011712f
C788 VTAIL.n731 VSUBS 0.021795f
C789 VTAIL.n732 VSUBS 0.021795f
C790 VTAIL.n733 VSUBS 0.011712f
C791 VTAIL.n734 VSUBS 0.012401f
C792 VTAIL.n735 VSUBS 0.027682f
C793 VTAIL.n736 VSUBS 0.06765f
C794 VTAIL.n737 VSUBS 0.012401f
C795 VTAIL.n738 VSUBS 0.011712f
C796 VTAIL.n739 VSUBS 0.050081f
C797 VTAIL.n740 VSUBS 0.034039f
C798 VTAIL.n741 VSUBS 1.61556f
C799 VTAIL.n742 VSUBS 0.024134f
C800 VTAIL.n743 VSUBS 0.021795f
C801 VTAIL.n744 VSUBS 0.011712f
C802 VTAIL.n745 VSUBS 0.027682f
C803 VTAIL.n746 VSUBS 0.012401f
C804 VTAIL.n747 VSUBS 0.021795f
C805 VTAIL.n748 VSUBS 0.011712f
C806 VTAIL.n749 VSUBS 0.027682f
C807 VTAIL.n750 VSUBS 0.012401f
C808 VTAIL.n751 VSUBS 0.021795f
C809 VTAIL.n752 VSUBS 0.011712f
C810 VTAIL.n753 VSUBS 0.027682f
C811 VTAIL.n754 VSUBS 0.012401f
C812 VTAIL.n755 VSUBS 0.021795f
C813 VTAIL.n756 VSUBS 0.011712f
C814 VTAIL.n757 VSUBS 0.027682f
C815 VTAIL.n758 VSUBS 0.012401f
C816 VTAIL.n759 VSUBS 0.021795f
C817 VTAIL.n760 VSUBS 0.011712f
C818 VTAIL.n761 VSUBS 0.027682f
C819 VTAIL.n762 VSUBS 0.012401f
C820 VTAIL.n763 VSUBS 0.021795f
C821 VTAIL.n764 VSUBS 0.011712f
C822 VTAIL.n765 VSUBS 0.027682f
C823 VTAIL.n766 VSUBS 0.012401f
C824 VTAIL.n767 VSUBS 0.021795f
C825 VTAIL.n768 VSUBS 0.011712f
C826 VTAIL.n769 VSUBS 0.027682f
C827 VTAIL.n770 VSUBS 0.012401f
C828 VTAIL.n771 VSUBS 0.021795f
C829 VTAIL.n772 VSUBS 0.011712f
C830 VTAIL.n773 VSUBS 0.027682f
C831 VTAIL.n774 VSUBS 0.012401f
C832 VTAIL.n775 VSUBS 0.17903f
C833 VTAIL.t6 VSUBS 0.059476f
C834 VTAIL.n776 VSUBS 0.020762f
C835 VTAIL.n777 VSUBS 0.01761f
C836 VTAIL.n778 VSUBS 0.011712f
C837 VTAIL.n779 VSUBS 1.78249f
C838 VTAIL.n780 VSUBS 0.021795f
C839 VTAIL.n781 VSUBS 0.011712f
C840 VTAIL.n782 VSUBS 0.012401f
C841 VTAIL.n783 VSUBS 0.027682f
C842 VTAIL.n784 VSUBS 0.027682f
C843 VTAIL.n785 VSUBS 0.012401f
C844 VTAIL.n786 VSUBS 0.011712f
C845 VTAIL.n787 VSUBS 0.021795f
C846 VTAIL.n788 VSUBS 0.021795f
C847 VTAIL.n789 VSUBS 0.011712f
C848 VTAIL.n790 VSUBS 0.012401f
C849 VTAIL.n791 VSUBS 0.027682f
C850 VTAIL.n792 VSUBS 0.027682f
C851 VTAIL.n793 VSUBS 0.012401f
C852 VTAIL.n794 VSUBS 0.011712f
C853 VTAIL.n795 VSUBS 0.021795f
C854 VTAIL.n796 VSUBS 0.021795f
C855 VTAIL.n797 VSUBS 0.011712f
C856 VTAIL.n798 VSUBS 0.012401f
C857 VTAIL.n799 VSUBS 0.027682f
C858 VTAIL.n800 VSUBS 0.027682f
C859 VTAIL.n801 VSUBS 0.012401f
C860 VTAIL.n802 VSUBS 0.011712f
C861 VTAIL.n803 VSUBS 0.021795f
C862 VTAIL.n804 VSUBS 0.021795f
C863 VTAIL.n805 VSUBS 0.011712f
C864 VTAIL.n806 VSUBS 0.012401f
C865 VTAIL.n807 VSUBS 0.027682f
C866 VTAIL.n808 VSUBS 0.027682f
C867 VTAIL.n809 VSUBS 0.012401f
C868 VTAIL.n810 VSUBS 0.011712f
C869 VTAIL.n811 VSUBS 0.021795f
C870 VTAIL.n812 VSUBS 0.021795f
C871 VTAIL.n813 VSUBS 0.011712f
C872 VTAIL.n814 VSUBS 0.012401f
C873 VTAIL.n815 VSUBS 0.027682f
C874 VTAIL.n816 VSUBS 0.027682f
C875 VTAIL.n817 VSUBS 0.027682f
C876 VTAIL.n818 VSUBS 0.012401f
C877 VTAIL.n819 VSUBS 0.011712f
C878 VTAIL.n820 VSUBS 0.021795f
C879 VTAIL.n821 VSUBS 0.021795f
C880 VTAIL.n822 VSUBS 0.011712f
C881 VTAIL.n823 VSUBS 0.012056f
C882 VTAIL.n824 VSUBS 0.012056f
C883 VTAIL.n825 VSUBS 0.027682f
C884 VTAIL.n826 VSUBS 0.027682f
C885 VTAIL.n827 VSUBS 0.012401f
C886 VTAIL.n828 VSUBS 0.011712f
C887 VTAIL.n829 VSUBS 0.021795f
C888 VTAIL.n830 VSUBS 0.021795f
C889 VTAIL.n831 VSUBS 0.011712f
C890 VTAIL.n832 VSUBS 0.012401f
C891 VTAIL.n833 VSUBS 0.027682f
C892 VTAIL.n834 VSUBS 0.027682f
C893 VTAIL.n835 VSUBS 0.012401f
C894 VTAIL.n836 VSUBS 0.011712f
C895 VTAIL.n837 VSUBS 0.021795f
C896 VTAIL.n838 VSUBS 0.021795f
C897 VTAIL.n839 VSUBS 0.011712f
C898 VTAIL.n840 VSUBS 0.012401f
C899 VTAIL.n841 VSUBS 0.027682f
C900 VTAIL.n842 VSUBS 0.06765f
C901 VTAIL.n843 VSUBS 0.012401f
C902 VTAIL.n844 VSUBS 0.011712f
C903 VTAIL.n845 VSUBS 0.050081f
C904 VTAIL.n846 VSUBS 0.034039f
C905 VTAIL.n847 VSUBS 1.57302f
C906 VN.t3 VSUBS 2.59004f
C907 VN.t0 VSUBS 2.58987f
C908 VN.n0 VSUBS 1.85216f
C909 VN.t2 VSUBS 2.59004f
C910 VN.t1 VSUBS 2.58987f
C911 VN.n1 VSUBS 3.43893f
C912 B.n0 VSUBS 0.00651f
C913 B.n1 VSUBS 0.00651f
C914 B.n2 VSUBS 0.009628f
C915 B.n3 VSUBS 0.007378f
C916 B.n4 VSUBS 0.007378f
C917 B.n5 VSUBS 0.007378f
C918 B.n6 VSUBS 0.007378f
C919 B.n7 VSUBS 0.007378f
C920 B.n8 VSUBS 0.007378f
C921 B.n9 VSUBS 0.007378f
C922 B.n10 VSUBS 0.007378f
C923 B.n11 VSUBS 0.015506f
C924 B.n12 VSUBS 0.007378f
C925 B.n13 VSUBS 0.007378f
C926 B.n14 VSUBS 0.007378f
C927 B.n15 VSUBS 0.007378f
C928 B.n16 VSUBS 0.007378f
C929 B.n17 VSUBS 0.007378f
C930 B.n18 VSUBS 0.007378f
C931 B.n19 VSUBS 0.007378f
C932 B.n20 VSUBS 0.007378f
C933 B.n21 VSUBS 0.007378f
C934 B.n22 VSUBS 0.007378f
C935 B.n23 VSUBS 0.007378f
C936 B.n24 VSUBS 0.007378f
C937 B.n25 VSUBS 0.007378f
C938 B.n26 VSUBS 0.007378f
C939 B.n27 VSUBS 0.007378f
C940 B.n28 VSUBS 0.007378f
C941 B.n29 VSUBS 0.007378f
C942 B.n30 VSUBS 0.007378f
C943 B.n31 VSUBS 0.007378f
C944 B.n32 VSUBS 0.007378f
C945 B.n33 VSUBS 0.007378f
C946 B.n34 VSUBS 0.007378f
C947 B.n35 VSUBS 0.007378f
C948 B.n36 VSUBS 0.007378f
C949 B.n37 VSUBS 0.007378f
C950 B.n38 VSUBS 0.007378f
C951 B.n39 VSUBS 0.007378f
C952 B.n40 VSUBS 0.007378f
C953 B.n41 VSUBS 0.007378f
C954 B.n42 VSUBS 0.006944f
C955 B.n43 VSUBS 0.007378f
C956 B.t1 VSUBS 0.39449f
C957 B.t2 VSUBS 0.410446f
C958 B.t0 VSUBS 0.768923f
C959 B.n44 VSUBS 0.515293f
C960 B.n45 VSUBS 0.351003f
C961 B.n46 VSUBS 0.017095f
C962 B.n47 VSUBS 0.007378f
C963 B.n48 VSUBS 0.007378f
C964 B.n49 VSUBS 0.007378f
C965 B.n50 VSUBS 0.007378f
C966 B.t4 VSUBS 0.394493f
C967 B.t5 VSUBS 0.41045f
C968 B.t3 VSUBS 0.768923f
C969 B.n51 VSUBS 0.515289f
C970 B.n52 VSUBS 0.350999f
C971 B.n53 VSUBS 0.007378f
C972 B.n54 VSUBS 0.007378f
C973 B.n55 VSUBS 0.007378f
C974 B.n56 VSUBS 0.007378f
C975 B.n57 VSUBS 0.007378f
C976 B.n58 VSUBS 0.007378f
C977 B.n59 VSUBS 0.007378f
C978 B.n60 VSUBS 0.007378f
C979 B.n61 VSUBS 0.007378f
C980 B.n62 VSUBS 0.007378f
C981 B.n63 VSUBS 0.007378f
C982 B.n64 VSUBS 0.007378f
C983 B.n65 VSUBS 0.007378f
C984 B.n66 VSUBS 0.007378f
C985 B.n67 VSUBS 0.007378f
C986 B.n68 VSUBS 0.007378f
C987 B.n69 VSUBS 0.007378f
C988 B.n70 VSUBS 0.007378f
C989 B.n71 VSUBS 0.007378f
C990 B.n72 VSUBS 0.007378f
C991 B.n73 VSUBS 0.007378f
C992 B.n74 VSUBS 0.007378f
C993 B.n75 VSUBS 0.007378f
C994 B.n76 VSUBS 0.007378f
C995 B.n77 VSUBS 0.007378f
C996 B.n78 VSUBS 0.007378f
C997 B.n79 VSUBS 0.007378f
C998 B.n80 VSUBS 0.007378f
C999 B.n81 VSUBS 0.007378f
C1000 B.n82 VSUBS 0.007378f
C1001 B.n83 VSUBS 0.016395f
C1002 B.n84 VSUBS 0.007378f
C1003 B.n85 VSUBS 0.007378f
C1004 B.n86 VSUBS 0.007378f
C1005 B.n87 VSUBS 0.007378f
C1006 B.n88 VSUBS 0.007378f
C1007 B.n89 VSUBS 0.007378f
C1008 B.n90 VSUBS 0.007378f
C1009 B.n91 VSUBS 0.007378f
C1010 B.n92 VSUBS 0.007378f
C1011 B.n93 VSUBS 0.007378f
C1012 B.n94 VSUBS 0.007378f
C1013 B.n95 VSUBS 0.007378f
C1014 B.n96 VSUBS 0.007378f
C1015 B.n97 VSUBS 0.007378f
C1016 B.n98 VSUBS 0.007378f
C1017 B.n99 VSUBS 0.007378f
C1018 B.n100 VSUBS 0.007378f
C1019 B.n101 VSUBS 0.007378f
C1020 B.n102 VSUBS 0.007378f
C1021 B.n103 VSUBS 0.016492f
C1022 B.n104 VSUBS 0.007378f
C1023 B.n105 VSUBS 0.007378f
C1024 B.n106 VSUBS 0.007378f
C1025 B.n107 VSUBS 0.007378f
C1026 B.n108 VSUBS 0.007378f
C1027 B.n109 VSUBS 0.007378f
C1028 B.n110 VSUBS 0.007378f
C1029 B.n111 VSUBS 0.007378f
C1030 B.n112 VSUBS 0.007378f
C1031 B.n113 VSUBS 0.007378f
C1032 B.n114 VSUBS 0.007378f
C1033 B.n115 VSUBS 0.007378f
C1034 B.n116 VSUBS 0.007378f
C1035 B.n117 VSUBS 0.007378f
C1036 B.n118 VSUBS 0.007378f
C1037 B.n119 VSUBS 0.007378f
C1038 B.n120 VSUBS 0.007378f
C1039 B.n121 VSUBS 0.007378f
C1040 B.n122 VSUBS 0.007378f
C1041 B.n123 VSUBS 0.007378f
C1042 B.n124 VSUBS 0.007378f
C1043 B.n125 VSUBS 0.007378f
C1044 B.n126 VSUBS 0.007378f
C1045 B.n127 VSUBS 0.007378f
C1046 B.n128 VSUBS 0.007378f
C1047 B.n129 VSUBS 0.007378f
C1048 B.n130 VSUBS 0.007378f
C1049 B.n131 VSUBS 0.007378f
C1050 B.n132 VSUBS 0.007378f
C1051 B.n133 VSUBS 0.007378f
C1052 B.n134 VSUBS 0.007378f
C1053 B.t8 VSUBS 0.394493f
C1054 B.t7 VSUBS 0.41045f
C1055 B.t6 VSUBS 0.768923f
C1056 B.n135 VSUBS 0.515289f
C1057 B.n136 VSUBS 0.350999f
C1058 B.n137 VSUBS 0.007378f
C1059 B.n138 VSUBS 0.007378f
C1060 B.n139 VSUBS 0.007378f
C1061 B.n140 VSUBS 0.007378f
C1062 B.n141 VSUBS 0.004123f
C1063 B.n142 VSUBS 0.007378f
C1064 B.n143 VSUBS 0.007378f
C1065 B.n144 VSUBS 0.007378f
C1066 B.n145 VSUBS 0.007378f
C1067 B.n146 VSUBS 0.007378f
C1068 B.n147 VSUBS 0.007378f
C1069 B.n148 VSUBS 0.007378f
C1070 B.n149 VSUBS 0.007378f
C1071 B.n150 VSUBS 0.007378f
C1072 B.n151 VSUBS 0.007378f
C1073 B.n152 VSUBS 0.007378f
C1074 B.n153 VSUBS 0.007378f
C1075 B.n154 VSUBS 0.007378f
C1076 B.n155 VSUBS 0.007378f
C1077 B.n156 VSUBS 0.007378f
C1078 B.n157 VSUBS 0.007378f
C1079 B.n158 VSUBS 0.007378f
C1080 B.n159 VSUBS 0.007378f
C1081 B.n160 VSUBS 0.007378f
C1082 B.n161 VSUBS 0.007378f
C1083 B.n162 VSUBS 0.007378f
C1084 B.n163 VSUBS 0.007378f
C1085 B.n164 VSUBS 0.007378f
C1086 B.n165 VSUBS 0.007378f
C1087 B.n166 VSUBS 0.007378f
C1088 B.n167 VSUBS 0.007378f
C1089 B.n168 VSUBS 0.007378f
C1090 B.n169 VSUBS 0.007378f
C1091 B.n170 VSUBS 0.007378f
C1092 B.n171 VSUBS 0.007378f
C1093 B.n172 VSUBS 0.016395f
C1094 B.n173 VSUBS 0.007378f
C1095 B.n174 VSUBS 0.007378f
C1096 B.n175 VSUBS 0.007378f
C1097 B.n176 VSUBS 0.007378f
C1098 B.n177 VSUBS 0.007378f
C1099 B.n178 VSUBS 0.007378f
C1100 B.n179 VSUBS 0.007378f
C1101 B.n180 VSUBS 0.007378f
C1102 B.n181 VSUBS 0.007378f
C1103 B.n182 VSUBS 0.007378f
C1104 B.n183 VSUBS 0.007378f
C1105 B.n184 VSUBS 0.007378f
C1106 B.n185 VSUBS 0.007378f
C1107 B.n186 VSUBS 0.007378f
C1108 B.n187 VSUBS 0.007378f
C1109 B.n188 VSUBS 0.007378f
C1110 B.n189 VSUBS 0.007378f
C1111 B.n190 VSUBS 0.007378f
C1112 B.n191 VSUBS 0.007378f
C1113 B.n192 VSUBS 0.007378f
C1114 B.n193 VSUBS 0.007378f
C1115 B.n194 VSUBS 0.007378f
C1116 B.n195 VSUBS 0.007378f
C1117 B.n196 VSUBS 0.007378f
C1118 B.n197 VSUBS 0.007378f
C1119 B.n198 VSUBS 0.007378f
C1120 B.n199 VSUBS 0.007378f
C1121 B.n200 VSUBS 0.007378f
C1122 B.n201 VSUBS 0.007378f
C1123 B.n202 VSUBS 0.007378f
C1124 B.n203 VSUBS 0.007378f
C1125 B.n204 VSUBS 0.007378f
C1126 B.n205 VSUBS 0.007378f
C1127 B.n206 VSUBS 0.007378f
C1128 B.n207 VSUBS 0.015506f
C1129 B.n208 VSUBS 0.015506f
C1130 B.n209 VSUBS 0.016395f
C1131 B.n210 VSUBS 0.007378f
C1132 B.n211 VSUBS 0.007378f
C1133 B.n212 VSUBS 0.007378f
C1134 B.n213 VSUBS 0.007378f
C1135 B.n214 VSUBS 0.007378f
C1136 B.n215 VSUBS 0.007378f
C1137 B.n216 VSUBS 0.007378f
C1138 B.n217 VSUBS 0.007378f
C1139 B.n218 VSUBS 0.007378f
C1140 B.n219 VSUBS 0.007378f
C1141 B.n220 VSUBS 0.007378f
C1142 B.n221 VSUBS 0.007378f
C1143 B.n222 VSUBS 0.007378f
C1144 B.n223 VSUBS 0.007378f
C1145 B.n224 VSUBS 0.007378f
C1146 B.n225 VSUBS 0.007378f
C1147 B.n226 VSUBS 0.007378f
C1148 B.n227 VSUBS 0.007378f
C1149 B.n228 VSUBS 0.007378f
C1150 B.n229 VSUBS 0.007378f
C1151 B.n230 VSUBS 0.007378f
C1152 B.n231 VSUBS 0.007378f
C1153 B.n232 VSUBS 0.007378f
C1154 B.n233 VSUBS 0.007378f
C1155 B.n234 VSUBS 0.007378f
C1156 B.n235 VSUBS 0.007378f
C1157 B.n236 VSUBS 0.007378f
C1158 B.n237 VSUBS 0.007378f
C1159 B.n238 VSUBS 0.007378f
C1160 B.n239 VSUBS 0.007378f
C1161 B.n240 VSUBS 0.007378f
C1162 B.n241 VSUBS 0.007378f
C1163 B.n242 VSUBS 0.007378f
C1164 B.n243 VSUBS 0.007378f
C1165 B.n244 VSUBS 0.007378f
C1166 B.n245 VSUBS 0.007378f
C1167 B.n246 VSUBS 0.007378f
C1168 B.n247 VSUBS 0.007378f
C1169 B.n248 VSUBS 0.007378f
C1170 B.n249 VSUBS 0.007378f
C1171 B.n250 VSUBS 0.007378f
C1172 B.n251 VSUBS 0.007378f
C1173 B.n252 VSUBS 0.007378f
C1174 B.n253 VSUBS 0.007378f
C1175 B.n254 VSUBS 0.007378f
C1176 B.n255 VSUBS 0.007378f
C1177 B.n256 VSUBS 0.007378f
C1178 B.n257 VSUBS 0.007378f
C1179 B.n258 VSUBS 0.007378f
C1180 B.n259 VSUBS 0.007378f
C1181 B.n260 VSUBS 0.007378f
C1182 B.n261 VSUBS 0.007378f
C1183 B.n262 VSUBS 0.007378f
C1184 B.n263 VSUBS 0.007378f
C1185 B.n264 VSUBS 0.007378f
C1186 B.n265 VSUBS 0.007378f
C1187 B.n266 VSUBS 0.007378f
C1188 B.n267 VSUBS 0.007378f
C1189 B.n268 VSUBS 0.007378f
C1190 B.n269 VSUBS 0.007378f
C1191 B.n270 VSUBS 0.007378f
C1192 B.n271 VSUBS 0.007378f
C1193 B.n272 VSUBS 0.007378f
C1194 B.n273 VSUBS 0.007378f
C1195 B.n274 VSUBS 0.007378f
C1196 B.n275 VSUBS 0.007378f
C1197 B.n276 VSUBS 0.007378f
C1198 B.n277 VSUBS 0.007378f
C1199 B.n278 VSUBS 0.007378f
C1200 B.n279 VSUBS 0.007378f
C1201 B.n280 VSUBS 0.007378f
C1202 B.n281 VSUBS 0.007378f
C1203 B.n282 VSUBS 0.007378f
C1204 B.n283 VSUBS 0.007378f
C1205 B.n284 VSUBS 0.007378f
C1206 B.n285 VSUBS 0.007378f
C1207 B.n286 VSUBS 0.007378f
C1208 B.n287 VSUBS 0.007378f
C1209 B.n288 VSUBS 0.007378f
C1210 B.n289 VSUBS 0.007378f
C1211 B.n290 VSUBS 0.007378f
C1212 B.n291 VSUBS 0.007378f
C1213 B.n292 VSUBS 0.007378f
C1214 B.n293 VSUBS 0.007378f
C1215 B.n294 VSUBS 0.007378f
C1216 B.n295 VSUBS 0.007378f
C1217 B.n296 VSUBS 0.007378f
C1218 B.n297 VSUBS 0.007378f
C1219 B.n298 VSUBS 0.007378f
C1220 B.n299 VSUBS 0.007378f
C1221 B.t11 VSUBS 0.39449f
C1222 B.t10 VSUBS 0.410446f
C1223 B.t9 VSUBS 0.768923f
C1224 B.n300 VSUBS 0.515293f
C1225 B.n301 VSUBS 0.351003f
C1226 B.n302 VSUBS 0.017095f
C1227 B.n303 VSUBS 0.006944f
C1228 B.n304 VSUBS 0.007378f
C1229 B.n305 VSUBS 0.007378f
C1230 B.n306 VSUBS 0.007378f
C1231 B.n307 VSUBS 0.007378f
C1232 B.n308 VSUBS 0.007378f
C1233 B.n309 VSUBS 0.007378f
C1234 B.n310 VSUBS 0.007378f
C1235 B.n311 VSUBS 0.007378f
C1236 B.n312 VSUBS 0.007378f
C1237 B.n313 VSUBS 0.007378f
C1238 B.n314 VSUBS 0.007378f
C1239 B.n315 VSUBS 0.007378f
C1240 B.n316 VSUBS 0.007378f
C1241 B.n317 VSUBS 0.007378f
C1242 B.n318 VSUBS 0.007378f
C1243 B.n319 VSUBS 0.004123f
C1244 B.n320 VSUBS 0.017095f
C1245 B.n321 VSUBS 0.006944f
C1246 B.n322 VSUBS 0.007378f
C1247 B.n323 VSUBS 0.007378f
C1248 B.n324 VSUBS 0.007378f
C1249 B.n325 VSUBS 0.007378f
C1250 B.n326 VSUBS 0.007378f
C1251 B.n327 VSUBS 0.007378f
C1252 B.n328 VSUBS 0.007378f
C1253 B.n329 VSUBS 0.007378f
C1254 B.n330 VSUBS 0.007378f
C1255 B.n331 VSUBS 0.007378f
C1256 B.n332 VSUBS 0.007378f
C1257 B.n333 VSUBS 0.007378f
C1258 B.n334 VSUBS 0.007378f
C1259 B.n335 VSUBS 0.007378f
C1260 B.n336 VSUBS 0.007378f
C1261 B.n337 VSUBS 0.007378f
C1262 B.n338 VSUBS 0.007378f
C1263 B.n339 VSUBS 0.007378f
C1264 B.n340 VSUBS 0.007378f
C1265 B.n341 VSUBS 0.007378f
C1266 B.n342 VSUBS 0.007378f
C1267 B.n343 VSUBS 0.007378f
C1268 B.n344 VSUBS 0.007378f
C1269 B.n345 VSUBS 0.007378f
C1270 B.n346 VSUBS 0.007378f
C1271 B.n347 VSUBS 0.007378f
C1272 B.n348 VSUBS 0.007378f
C1273 B.n349 VSUBS 0.007378f
C1274 B.n350 VSUBS 0.007378f
C1275 B.n351 VSUBS 0.007378f
C1276 B.n352 VSUBS 0.007378f
C1277 B.n353 VSUBS 0.007378f
C1278 B.n354 VSUBS 0.007378f
C1279 B.n355 VSUBS 0.007378f
C1280 B.n356 VSUBS 0.007378f
C1281 B.n357 VSUBS 0.007378f
C1282 B.n358 VSUBS 0.007378f
C1283 B.n359 VSUBS 0.007378f
C1284 B.n360 VSUBS 0.007378f
C1285 B.n361 VSUBS 0.007378f
C1286 B.n362 VSUBS 0.007378f
C1287 B.n363 VSUBS 0.007378f
C1288 B.n364 VSUBS 0.007378f
C1289 B.n365 VSUBS 0.007378f
C1290 B.n366 VSUBS 0.007378f
C1291 B.n367 VSUBS 0.007378f
C1292 B.n368 VSUBS 0.007378f
C1293 B.n369 VSUBS 0.007378f
C1294 B.n370 VSUBS 0.007378f
C1295 B.n371 VSUBS 0.007378f
C1296 B.n372 VSUBS 0.007378f
C1297 B.n373 VSUBS 0.007378f
C1298 B.n374 VSUBS 0.007378f
C1299 B.n375 VSUBS 0.007378f
C1300 B.n376 VSUBS 0.007378f
C1301 B.n377 VSUBS 0.007378f
C1302 B.n378 VSUBS 0.007378f
C1303 B.n379 VSUBS 0.007378f
C1304 B.n380 VSUBS 0.007378f
C1305 B.n381 VSUBS 0.007378f
C1306 B.n382 VSUBS 0.007378f
C1307 B.n383 VSUBS 0.007378f
C1308 B.n384 VSUBS 0.007378f
C1309 B.n385 VSUBS 0.007378f
C1310 B.n386 VSUBS 0.007378f
C1311 B.n387 VSUBS 0.007378f
C1312 B.n388 VSUBS 0.007378f
C1313 B.n389 VSUBS 0.007378f
C1314 B.n390 VSUBS 0.007378f
C1315 B.n391 VSUBS 0.007378f
C1316 B.n392 VSUBS 0.007378f
C1317 B.n393 VSUBS 0.007378f
C1318 B.n394 VSUBS 0.007378f
C1319 B.n395 VSUBS 0.007378f
C1320 B.n396 VSUBS 0.007378f
C1321 B.n397 VSUBS 0.007378f
C1322 B.n398 VSUBS 0.007378f
C1323 B.n399 VSUBS 0.007378f
C1324 B.n400 VSUBS 0.007378f
C1325 B.n401 VSUBS 0.007378f
C1326 B.n402 VSUBS 0.007378f
C1327 B.n403 VSUBS 0.007378f
C1328 B.n404 VSUBS 0.007378f
C1329 B.n405 VSUBS 0.007378f
C1330 B.n406 VSUBS 0.007378f
C1331 B.n407 VSUBS 0.007378f
C1332 B.n408 VSUBS 0.007378f
C1333 B.n409 VSUBS 0.007378f
C1334 B.n410 VSUBS 0.007378f
C1335 B.n411 VSUBS 0.007378f
C1336 B.n412 VSUBS 0.015409f
C1337 B.n413 VSUBS 0.016395f
C1338 B.n414 VSUBS 0.015506f
C1339 B.n415 VSUBS 0.007378f
C1340 B.n416 VSUBS 0.007378f
C1341 B.n417 VSUBS 0.007378f
C1342 B.n418 VSUBS 0.007378f
C1343 B.n419 VSUBS 0.007378f
C1344 B.n420 VSUBS 0.007378f
C1345 B.n421 VSUBS 0.007378f
C1346 B.n422 VSUBS 0.007378f
C1347 B.n423 VSUBS 0.007378f
C1348 B.n424 VSUBS 0.007378f
C1349 B.n425 VSUBS 0.007378f
C1350 B.n426 VSUBS 0.007378f
C1351 B.n427 VSUBS 0.007378f
C1352 B.n428 VSUBS 0.007378f
C1353 B.n429 VSUBS 0.007378f
C1354 B.n430 VSUBS 0.007378f
C1355 B.n431 VSUBS 0.007378f
C1356 B.n432 VSUBS 0.007378f
C1357 B.n433 VSUBS 0.007378f
C1358 B.n434 VSUBS 0.007378f
C1359 B.n435 VSUBS 0.007378f
C1360 B.n436 VSUBS 0.007378f
C1361 B.n437 VSUBS 0.007378f
C1362 B.n438 VSUBS 0.007378f
C1363 B.n439 VSUBS 0.007378f
C1364 B.n440 VSUBS 0.007378f
C1365 B.n441 VSUBS 0.007378f
C1366 B.n442 VSUBS 0.007378f
C1367 B.n443 VSUBS 0.007378f
C1368 B.n444 VSUBS 0.007378f
C1369 B.n445 VSUBS 0.007378f
C1370 B.n446 VSUBS 0.007378f
C1371 B.n447 VSUBS 0.007378f
C1372 B.n448 VSUBS 0.007378f
C1373 B.n449 VSUBS 0.007378f
C1374 B.n450 VSUBS 0.007378f
C1375 B.n451 VSUBS 0.007378f
C1376 B.n452 VSUBS 0.007378f
C1377 B.n453 VSUBS 0.007378f
C1378 B.n454 VSUBS 0.007378f
C1379 B.n455 VSUBS 0.007378f
C1380 B.n456 VSUBS 0.007378f
C1381 B.n457 VSUBS 0.007378f
C1382 B.n458 VSUBS 0.007378f
C1383 B.n459 VSUBS 0.007378f
C1384 B.n460 VSUBS 0.007378f
C1385 B.n461 VSUBS 0.007378f
C1386 B.n462 VSUBS 0.007378f
C1387 B.n463 VSUBS 0.007378f
C1388 B.n464 VSUBS 0.007378f
C1389 B.n465 VSUBS 0.007378f
C1390 B.n466 VSUBS 0.007378f
C1391 B.n467 VSUBS 0.007378f
C1392 B.n468 VSUBS 0.007378f
C1393 B.n469 VSUBS 0.007378f
C1394 B.n470 VSUBS 0.007378f
C1395 B.n471 VSUBS 0.007378f
C1396 B.n472 VSUBS 0.015506f
C1397 B.n473 VSUBS 0.015506f
C1398 B.n474 VSUBS 0.016395f
C1399 B.n475 VSUBS 0.007378f
C1400 B.n476 VSUBS 0.007378f
C1401 B.n477 VSUBS 0.007378f
C1402 B.n478 VSUBS 0.007378f
C1403 B.n479 VSUBS 0.007378f
C1404 B.n480 VSUBS 0.007378f
C1405 B.n481 VSUBS 0.007378f
C1406 B.n482 VSUBS 0.007378f
C1407 B.n483 VSUBS 0.007378f
C1408 B.n484 VSUBS 0.007378f
C1409 B.n485 VSUBS 0.007378f
C1410 B.n486 VSUBS 0.007378f
C1411 B.n487 VSUBS 0.007378f
C1412 B.n488 VSUBS 0.007378f
C1413 B.n489 VSUBS 0.007378f
C1414 B.n490 VSUBS 0.007378f
C1415 B.n491 VSUBS 0.007378f
C1416 B.n492 VSUBS 0.007378f
C1417 B.n493 VSUBS 0.007378f
C1418 B.n494 VSUBS 0.007378f
C1419 B.n495 VSUBS 0.007378f
C1420 B.n496 VSUBS 0.007378f
C1421 B.n497 VSUBS 0.007378f
C1422 B.n498 VSUBS 0.007378f
C1423 B.n499 VSUBS 0.007378f
C1424 B.n500 VSUBS 0.007378f
C1425 B.n501 VSUBS 0.007378f
C1426 B.n502 VSUBS 0.007378f
C1427 B.n503 VSUBS 0.007378f
C1428 B.n504 VSUBS 0.007378f
C1429 B.n505 VSUBS 0.007378f
C1430 B.n506 VSUBS 0.007378f
C1431 B.n507 VSUBS 0.007378f
C1432 B.n508 VSUBS 0.007378f
C1433 B.n509 VSUBS 0.007378f
C1434 B.n510 VSUBS 0.007378f
C1435 B.n511 VSUBS 0.007378f
C1436 B.n512 VSUBS 0.007378f
C1437 B.n513 VSUBS 0.007378f
C1438 B.n514 VSUBS 0.007378f
C1439 B.n515 VSUBS 0.007378f
C1440 B.n516 VSUBS 0.007378f
C1441 B.n517 VSUBS 0.007378f
C1442 B.n518 VSUBS 0.007378f
C1443 B.n519 VSUBS 0.007378f
C1444 B.n520 VSUBS 0.007378f
C1445 B.n521 VSUBS 0.007378f
C1446 B.n522 VSUBS 0.007378f
C1447 B.n523 VSUBS 0.007378f
C1448 B.n524 VSUBS 0.007378f
C1449 B.n525 VSUBS 0.007378f
C1450 B.n526 VSUBS 0.007378f
C1451 B.n527 VSUBS 0.007378f
C1452 B.n528 VSUBS 0.007378f
C1453 B.n529 VSUBS 0.007378f
C1454 B.n530 VSUBS 0.007378f
C1455 B.n531 VSUBS 0.007378f
C1456 B.n532 VSUBS 0.007378f
C1457 B.n533 VSUBS 0.007378f
C1458 B.n534 VSUBS 0.007378f
C1459 B.n535 VSUBS 0.007378f
C1460 B.n536 VSUBS 0.007378f
C1461 B.n537 VSUBS 0.007378f
C1462 B.n538 VSUBS 0.007378f
C1463 B.n539 VSUBS 0.007378f
C1464 B.n540 VSUBS 0.007378f
C1465 B.n541 VSUBS 0.007378f
C1466 B.n542 VSUBS 0.007378f
C1467 B.n543 VSUBS 0.007378f
C1468 B.n544 VSUBS 0.007378f
C1469 B.n545 VSUBS 0.007378f
C1470 B.n546 VSUBS 0.007378f
C1471 B.n547 VSUBS 0.007378f
C1472 B.n548 VSUBS 0.007378f
C1473 B.n549 VSUBS 0.007378f
C1474 B.n550 VSUBS 0.007378f
C1475 B.n551 VSUBS 0.007378f
C1476 B.n552 VSUBS 0.007378f
C1477 B.n553 VSUBS 0.007378f
C1478 B.n554 VSUBS 0.007378f
C1479 B.n555 VSUBS 0.007378f
C1480 B.n556 VSUBS 0.007378f
C1481 B.n557 VSUBS 0.007378f
C1482 B.n558 VSUBS 0.007378f
C1483 B.n559 VSUBS 0.007378f
C1484 B.n560 VSUBS 0.007378f
C1485 B.n561 VSUBS 0.007378f
C1486 B.n562 VSUBS 0.007378f
C1487 B.n563 VSUBS 0.007378f
C1488 B.n564 VSUBS 0.007378f
C1489 B.n565 VSUBS 0.007378f
C1490 B.n566 VSUBS 0.006944f
C1491 B.n567 VSUBS 0.017095f
C1492 B.n568 VSUBS 0.004123f
C1493 B.n569 VSUBS 0.007378f
C1494 B.n570 VSUBS 0.007378f
C1495 B.n571 VSUBS 0.007378f
C1496 B.n572 VSUBS 0.007378f
C1497 B.n573 VSUBS 0.007378f
C1498 B.n574 VSUBS 0.007378f
C1499 B.n575 VSUBS 0.007378f
C1500 B.n576 VSUBS 0.007378f
C1501 B.n577 VSUBS 0.007378f
C1502 B.n578 VSUBS 0.007378f
C1503 B.n579 VSUBS 0.007378f
C1504 B.n580 VSUBS 0.007378f
C1505 B.n581 VSUBS 0.004123f
C1506 B.n582 VSUBS 0.007378f
C1507 B.n583 VSUBS 0.007378f
C1508 B.n584 VSUBS 0.007378f
C1509 B.n585 VSUBS 0.007378f
C1510 B.n586 VSUBS 0.007378f
C1511 B.n587 VSUBS 0.007378f
C1512 B.n588 VSUBS 0.007378f
C1513 B.n589 VSUBS 0.007378f
C1514 B.n590 VSUBS 0.007378f
C1515 B.n591 VSUBS 0.007378f
C1516 B.n592 VSUBS 0.007378f
C1517 B.n593 VSUBS 0.007378f
C1518 B.n594 VSUBS 0.007378f
C1519 B.n595 VSUBS 0.007378f
C1520 B.n596 VSUBS 0.007378f
C1521 B.n597 VSUBS 0.007378f
C1522 B.n598 VSUBS 0.007378f
C1523 B.n599 VSUBS 0.007378f
C1524 B.n600 VSUBS 0.007378f
C1525 B.n601 VSUBS 0.007378f
C1526 B.n602 VSUBS 0.007378f
C1527 B.n603 VSUBS 0.007378f
C1528 B.n604 VSUBS 0.007378f
C1529 B.n605 VSUBS 0.007378f
C1530 B.n606 VSUBS 0.007378f
C1531 B.n607 VSUBS 0.007378f
C1532 B.n608 VSUBS 0.007378f
C1533 B.n609 VSUBS 0.007378f
C1534 B.n610 VSUBS 0.007378f
C1535 B.n611 VSUBS 0.007378f
C1536 B.n612 VSUBS 0.007378f
C1537 B.n613 VSUBS 0.007378f
C1538 B.n614 VSUBS 0.007378f
C1539 B.n615 VSUBS 0.007378f
C1540 B.n616 VSUBS 0.007378f
C1541 B.n617 VSUBS 0.007378f
C1542 B.n618 VSUBS 0.007378f
C1543 B.n619 VSUBS 0.007378f
C1544 B.n620 VSUBS 0.007378f
C1545 B.n621 VSUBS 0.007378f
C1546 B.n622 VSUBS 0.007378f
C1547 B.n623 VSUBS 0.007378f
C1548 B.n624 VSUBS 0.007378f
C1549 B.n625 VSUBS 0.007378f
C1550 B.n626 VSUBS 0.007378f
C1551 B.n627 VSUBS 0.007378f
C1552 B.n628 VSUBS 0.007378f
C1553 B.n629 VSUBS 0.007378f
C1554 B.n630 VSUBS 0.007378f
C1555 B.n631 VSUBS 0.007378f
C1556 B.n632 VSUBS 0.007378f
C1557 B.n633 VSUBS 0.007378f
C1558 B.n634 VSUBS 0.007378f
C1559 B.n635 VSUBS 0.007378f
C1560 B.n636 VSUBS 0.007378f
C1561 B.n637 VSUBS 0.007378f
C1562 B.n638 VSUBS 0.007378f
C1563 B.n639 VSUBS 0.007378f
C1564 B.n640 VSUBS 0.007378f
C1565 B.n641 VSUBS 0.007378f
C1566 B.n642 VSUBS 0.007378f
C1567 B.n643 VSUBS 0.007378f
C1568 B.n644 VSUBS 0.007378f
C1569 B.n645 VSUBS 0.007378f
C1570 B.n646 VSUBS 0.007378f
C1571 B.n647 VSUBS 0.007378f
C1572 B.n648 VSUBS 0.007378f
C1573 B.n649 VSUBS 0.007378f
C1574 B.n650 VSUBS 0.007378f
C1575 B.n651 VSUBS 0.007378f
C1576 B.n652 VSUBS 0.007378f
C1577 B.n653 VSUBS 0.007378f
C1578 B.n654 VSUBS 0.007378f
C1579 B.n655 VSUBS 0.007378f
C1580 B.n656 VSUBS 0.007378f
C1581 B.n657 VSUBS 0.007378f
C1582 B.n658 VSUBS 0.007378f
C1583 B.n659 VSUBS 0.007378f
C1584 B.n660 VSUBS 0.007378f
C1585 B.n661 VSUBS 0.007378f
C1586 B.n662 VSUBS 0.007378f
C1587 B.n663 VSUBS 0.007378f
C1588 B.n664 VSUBS 0.007378f
C1589 B.n665 VSUBS 0.007378f
C1590 B.n666 VSUBS 0.007378f
C1591 B.n667 VSUBS 0.007378f
C1592 B.n668 VSUBS 0.007378f
C1593 B.n669 VSUBS 0.007378f
C1594 B.n670 VSUBS 0.007378f
C1595 B.n671 VSUBS 0.007378f
C1596 B.n672 VSUBS 0.007378f
C1597 B.n673 VSUBS 0.007378f
C1598 B.n674 VSUBS 0.016395f
C1599 B.n675 VSUBS 0.016395f
C1600 B.n676 VSUBS 0.015506f
C1601 B.n677 VSUBS 0.007378f
C1602 B.n678 VSUBS 0.007378f
C1603 B.n679 VSUBS 0.007378f
C1604 B.n680 VSUBS 0.007378f
C1605 B.n681 VSUBS 0.007378f
C1606 B.n682 VSUBS 0.007378f
C1607 B.n683 VSUBS 0.007378f
C1608 B.n684 VSUBS 0.007378f
C1609 B.n685 VSUBS 0.007378f
C1610 B.n686 VSUBS 0.007378f
C1611 B.n687 VSUBS 0.007378f
C1612 B.n688 VSUBS 0.007378f
C1613 B.n689 VSUBS 0.007378f
C1614 B.n690 VSUBS 0.007378f
C1615 B.n691 VSUBS 0.007378f
C1616 B.n692 VSUBS 0.007378f
C1617 B.n693 VSUBS 0.007378f
C1618 B.n694 VSUBS 0.007378f
C1619 B.n695 VSUBS 0.007378f
C1620 B.n696 VSUBS 0.007378f
C1621 B.n697 VSUBS 0.007378f
C1622 B.n698 VSUBS 0.007378f
C1623 B.n699 VSUBS 0.007378f
C1624 B.n700 VSUBS 0.007378f
C1625 B.n701 VSUBS 0.007378f
C1626 B.n702 VSUBS 0.007378f
C1627 B.n703 VSUBS 0.009628f
C1628 B.n704 VSUBS 0.010257f
C1629 B.n705 VSUBS 0.020397f
.ends

