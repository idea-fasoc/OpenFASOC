* NGSPICE file created from diff_pair_sample_0663.ext - technology: sky130A

.subckt diff_pair_sample_0663 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0.81675 ps=5.28 w=4.95 l=2.42
X1 VDD1.t8 VP.t1 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0.81675 ps=5.28 w=4.95 l=2.42
X2 VDD1.t7 VP.t2 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X3 VDD1.t6 VP.t3 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=1.9305 ps=10.68 w=4.95 l=2.42
X4 VTAIL.t14 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X5 VDD2.t9 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X6 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=1.9305 ps=10.68 w=4.95 l=2.42
X7 VDD1.t4 VP.t5 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=1.9305 ps=10.68 w=4.95 l=2.42
X8 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X9 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.42
X10 VDD2.t6 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0.81675 ps=5.28 w=4.95 l=2.42
X11 VTAIL.t16 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X12 VDD2.t5 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=1.9305 ps=10.68 w=4.95 l=2.42
X13 VTAIL.t8 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X14 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.42
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.42
X16 VTAIL.t0 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X17 VTAIL.t17 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.42
X19 VTAIL.t18 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X20 VTAIL.t9 VN.t7 VDD2.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X21 VDD1.t0 VP.t9 VTAIL.t19 B.t3 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
X22 VDD2.t1 VN.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0.81675 ps=5.28 w=4.95 l=2.42
X23 VTAIL.t6 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.81675 pd=5.28 as=0.81675 ps=5.28 w=4.95 l=2.42
R0 VP.n23 VP.n22 161.3
R1 VP.n24 VP.n19 161.3
R2 VP.n26 VP.n25 161.3
R3 VP.n27 VP.n18 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n17 161.3
R6 VP.n33 VP.n32 161.3
R7 VP.n34 VP.n16 161.3
R8 VP.n36 VP.n35 161.3
R9 VP.n37 VP.n15 161.3
R10 VP.n39 VP.n38 161.3
R11 VP.n40 VP.n14 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n43 VP.n13 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n12 161.3
R16 VP.n83 VP.n0 161.3
R17 VP.n82 VP.n81 161.3
R18 VP.n80 VP.n1 161.3
R19 VP.n79 VP.n78 161.3
R20 VP.n77 VP.n2 161.3
R21 VP.n76 VP.n75 161.3
R22 VP.n74 VP.n3 161.3
R23 VP.n73 VP.n72 161.3
R24 VP.n71 VP.n4 161.3
R25 VP.n70 VP.n69 161.3
R26 VP.n68 VP.n5 161.3
R27 VP.n67 VP.n66 161.3
R28 VP.n64 VP.n6 161.3
R29 VP.n63 VP.n62 161.3
R30 VP.n61 VP.n7 161.3
R31 VP.n60 VP.n59 161.3
R32 VP.n58 VP.n8 161.3
R33 VP.n57 VP.n56 161.3
R34 VP.n55 VP.n9 161.3
R35 VP.n54 VP.n53 161.3
R36 VP.n52 VP.n10 161.3
R37 VP.n51 VP.n50 161.3
R38 VP.n49 VP.n11 98.5229
R39 VP.n85 VP.n84 98.5229
R40 VP.n48 VP.n47 98.5229
R41 VP.n20 VP.t1 83.6784
R42 VP.n53 VP.n9 52.6342
R43 VP.n63 VP.n7 52.6342
R44 VP.n72 VP.n71 52.6342
R45 VP.n78 VP.n1 52.6342
R46 VP.n41 VP.n13 52.6342
R47 VP.n35 VP.n34 52.6342
R48 VP.n26 VP.n19 52.6342
R49 VP.n76 VP.t7 49.296
R50 VP.n58 VP.t6 49.296
R51 VP.n11 VP.t0 49.296
R52 VP.n65 VP.t2 49.296
R53 VP.n84 VP.t5 49.296
R54 VP.n21 VP.t4 49.296
R55 VP.n39 VP.t8 49.296
R56 VP.n47 VP.t3 49.296
R57 VP.n28 VP.t9 49.296
R58 VP.n21 VP.n20 48.0049
R59 VP.n49 VP.n48 46.8064
R60 VP.n53 VP.n52 28.3526
R61 VP.n64 VP.n63 28.3526
R62 VP.n71 VP.n70 28.3526
R63 VP.n82 VP.n1 28.3526
R64 VP.n45 VP.n13 28.3526
R65 VP.n34 VP.n33 28.3526
R66 VP.n27 VP.n26 28.3526
R67 VP.n52 VP.n51 24.4675
R68 VP.n57 VP.n9 24.4675
R69 VP.n58 VP.n57 24.4675
R70 VP.n59 VP.n58 24.4675
R71 VP.n59 VP.n7 24.4675
R72 VP.n66 VP.n64 24.4675
R73 VP.n70 VP.n5 24.4675
R74 VP.n72 VP.n3 24.4675
R75 VP.n76 VP.n3 24.4675
R76 VP.n77 VP.n76 24.4675
R77 VP.n78 VP.n77 24.4675
R78 VP.n83 VP.n82 24.4675
R79 VP.n46 VP.n45 24.4675
R80 VP.n35 VP.n15 24.4675
R81 VP.n39 VP.n15 24.4675
R82 VP.n40 VP.n39 24.4675
R83 VP.n41 VP.n40 24.4675
R84 VP.n29 VP.n27 24.4675
R85 VP.n33 VP.n17 24.4675
R86 VP.n22 VP.n21 24.4675
R87 VP.n22 VP.n19 24.4675
R88 VP.n51 VP.n11 12.234
R89 VP.n66 VP.n65 12.234
R90 VP.n65 VP.n5 12.234
R91 VP.n84 VP.n83 12.234
R92 VP.n47 VP.n46 12.234
R93 VP.n29 VP.n28 12.234
R94 VP.n28 VP.n17 12.234
R95 VP.n23 VP.n20 6.69041
R96 VP.n48 VP.n12 0.278367
R97 VP.n50 VP.n49 0.278367
R98 VP.n85 VP.n0 0.278367
R99 VP.n24 VP.n23 0.189894
R100 VP.n25 VP.n24 0.189894
R101 VP.n25 VP.n18 0.189894
R102 VP.n30 VP.n18 0.189894
R103 VP.n31 VP.n30 0.189894
R104 VP.n32 VP.n31 0.189894
R105 VP.n32 VP.n16 0.189894
R106 VP.n36 VP.n16 0.189894
R107 VP.n37 VP.n36 0.189894
R108 VP.n38 VP.n37 0.189894
R109 VP.n38 VP.n14 0.189894
R110 VP.n42 VP.n14 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n44 VP.n43 0.189894
R113 VP.n44 VP.n12 0.189894
R114 VP.n50 VP.n10 0.189894
R115 VP.n54 VP.n10 0.189894
R116 VP.n55 VP.n54 0.189894
R117 VP.n56 VP.n55 0.189894
R118 VP.n56 VP.n8 0.189894
R119 VP.n60 VP.n8 0.189894
R120 VP.n61 VP.n60 0.189894
R121 VP.n62 VP.n61 0.189894
R122 VP.n62 VP.n6 0.189894
R123 VP.n67 VP.n6 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n69 VP.n68 0.189894
R126 VP.n69 VP.n4 0.189894
R127 VP.n73 VP.n4 0.189894
R128 VP.n74 VP.n73 0.189894
R129 VP.n75 VP.n74 0.189894
R130 VP.n75 VP.n2 0.189894
R131 VP.n79 VP.n2 0.189894
R132 VP.n80 VP.n79 0.189894
R133 VP.n81 VP.n80 0.189894
R134 VP.n81 VP.n0 0.189894
R135 VP VP.n85 0.153454
R136 VTAIL.n11 VTAIL.t7 57.47
R137 VTAIL.n17 VTAIL.t1 57.47
R138 VTAIL.n2 VTAIL.t15 57.47
R139 VTAIL.n16 VTAIL.t11 57.47
R140 VTAIL.n15 VTAIL.n14 53.4701
R141 VTAIL.n13 VTAIL.n12 53.4701
R142 VTAIL.n10 VTAIL.n9 53.4701
R143 VTAIL.n8 VTAIL.n7 53.4701
R144 VTAIL.n19 VTAIL.n18 53.4699
R145 VTAIL.n1 VTAIL.n0 53.4699
R146 VTAIL.n4 VTAIL.n3 53.4699
R147 VTAIL.n6 VTAIL.n5 53.4699
R148 VTAIL.n8 VTAIL.n6 21.3755
R149 VTAIL.n17 VTAIL.n16 19.0048
R150 VTAIL.n18 VTAIL.t3 4.0005
R151 VTAIL.n18 VTAIL.t0 4.0005
R152 VTAIL.n0 VTAIL.t5 4.0005
R153 VTAIL.n0 VTAIL.t6 4.0005
R154 VTAIL.n3 VTAIL.t12 4.0005
R155 VTAIL.n3 VTAIL.t17 4.0005
R156 VTAIL.n5 VTAIL.t10 4.0005
R157 VTAIL.n5 VTAIL.t16 4.0005
R158 VTAIL.n14 VTAIL.t19 4.0005
R159 VTAIL.n14 VTAIL.t18 4.0005
R160 VTAIL.n12 VTAIL.t13 4.0005
R161 VTAIL.n12 VTAIL.t14 4.0005
R162 VTAIL.n9 VTAIL.t4 4.0005
R163 VTAIL.n9 VTAIL.t9 4.0005
R164 VTAIL.n7 VTAIL.t2 4.0005
R165 VTAIL.n7 VTAIL.t8 4.0005
R166 VTAIL.n10 VTAIL.n8 2.37119
R167 VTAIL.n11 VTAIL.n10 2.37119
R168 VTAIL.n15 VTAIL.n13 2.37119
R169 VTAIL.n16 VTAIL.n15 2.37119
R170 VTAIL.n6 VTAIL.n4 2.37119
R171 VTAIL.n4 VTAIL.n2 2.37119
R172 VTAIL.n19 VTAIL.n17 2.37119
R173 VTAIL VTAIL.n1 1.83671
R174 VTAIL.n13 VTAIL.n11 1.65567
R175 VTAIL.n2 VTAIL.n1 1.65567
R176 VTAIL VTAIL.n19 0.534983
R177 VDD1.n1 VDD1.t8 76.5195
R178 VDD1.n3 VDD1.t9 76.5194
R179 VDD1.n5 VDD1.n4 71.8713
R180 VDD1.n1 VDD1.n0 70.1489
R181 VDD1.n7 VDD1.n6 70.1487
R182 VDD1.n3 VDD1.n2 70.1487
R183 VDD1.n7 VDD1.n5 41.0117
R184 VDD1.n6 VDD1.t1 4.0005
R185 VDD1.n6 VDD1.t6 4.0005
R186 VDD1.n0 VDD1.t5 4.0005
R187 VDD1.n0 VDD1.t0 4.0005
R188 VDD1.n4 VDD1.t2 4.0005
R189 VDD1.n4 VDD1.t4 4.0005
R190 VDD1.n2 VDD1.t3 4.0005
R191 VDD1.n2 VDD1.t7 4.0005
R192 VDD1 VDD1.n7 1.72033
R193 VDD1 VDD1.n1 0.651362
R194 VDD1.n5 VDD1.n3 0.537826
R195 B.n719 B.n718 585
R196 B.n720 B.n719 585
R197 B.n233 B.n130 585
R198 B.n232 B.n231 585
R199 B.n230 B.n229 585
R200 B.n228 B.n227 585
R201 B.n226 B.n225 585
R202 B.n224 B.n223 585
R203 B.n222 B.n221 585
R204 B.n220 B.n219 585
R205 B.n218 B.n217 585
R206 B.n216 B.n215 585
R207 B.n214 B.n213 585
R208 B.n212 B.n211 585
R209 B.n210 B.n209 585
R210 B.n208 B.n207 585
R211 B.n206 B.n205 585
R212 B.n204 B.n203 585
R213 B.n202 B.n201 585
R214 B.n200 B.n199 585
R215 B.n198 B.n197 585
R216 B.n196 B.n195 585
R217 B.n194 B.n193 585
R218 B.n192 B.n191 585
R219 B.n190 B.n189 585
R220 B.n188 B.n187 585
R221 B.n186 B.n185 585
R222 B.n184 B.n183 585
R223 B.n182 B.n181 585
R224 B.n180 B.n179 585
R225 B.n178 B.n177 585
R226 B.n175 B.n174 585
R227 B.n173 B.n172 585
R228 B.n171 B.n170 585
R229 B.n169 B.n168 585
R230 B.n167 B.n166 585
R231 B.n165 B.n164 585
R232 B.n163 B.n162 585
R233 B.n161 B.n160 585
R234 B.n159 B.n158 585
R235 B.n157 B.n156 585
R236 B.n155 B.n154 585
R237 B.n153 B.n152 585
R238 B.n151 B.n150 585
R239 B.n149 B.n148 585
R240 B.n147 B.n146 585
R241 B.n145 B.n144 585
R242 B.n143 B.n142 585
R243 B.n141 B.n140 585
R244 B.n139 B.n138 585
R245 B.n137 B.n136 585
R246 B.n103 B.n102 585
R247 B.n717 B.n104 585
R248 B.n721 B.n104 585
R249 B.n716 B.n715 585
R250 B.n715 B.n100 585
R251 B.n714 B.n99 585
R252 B.n727 B.n99 585
R253 B.n713 B.n98 585
R254 B.n728 B.n98 585
R255 B.n712 B.n97 585
R256 B.n729 B.n97 585
R257 B.n711 B.n710 585
R258 B.n710 B.n93 585
R259 B.n709 B.n92 585
R260 B.n735 B.n92 585
R261 B.n708 B.n91 585
R262 B.n736 B.n91 585
R263 B.n707 B.n90 585
R264 B.n737 B.n90 585
R265 B.n706 B.n705 585
R266 B.n705 B.n86 585
R267 B.n704 B.n85 585
R268 B.n743 B.n85 585
R269 B.n703 B.n84 585
R270 B.n744 B.n84 585
R271 B.n702 B.n83 585
R272 B.n745 B.n83 585
R273 B.n701 B.n700 585
R274 B.n700 B.n79 585
R275 B.n699 B.n78 585
R276 B.n751 B.n78 585
R277 B.n698 B.n77 585
R278 B.n752 B.n77 585
R279 B.n697 B.n76 585
R280 B.n753 B.n76 585
R281 B.n696 B.n695 585
R282 B.n695 B.n72 585
R283 B.n694 B.n71 585
R284 B.n759 B.n71 585
R285 B.n693 B.n70 585
R286 B.n760 B.n70 585
R287 B.n692 B.n69 585
R288 B.n761 B.n69 585
R289 B.n691 B.n690 585
R290 B.n690 B.n65 585
R291 B.n689 B.n64 585
R292 B.n767 B.n64 585
R293 B.n688 B.n63 585
R294 B.n768 B.n63 585
R295 B.n687 B.n62 585
R296 B.n769 B.n62 585
R297 B.n686 B.n685 585
R298 B.n685 B.n58 585
R299 B.n684 B.n57 585
R300 B.n775 B.n57 585
R301 B.n683 B.n56 585
R302 B.n776 B.n56 585
R303 B.n682 B.n55 585
R304 B.n777 B.n55 585
R305 B.n681 B.n680 585
R306 B.n680 B.n51 585
R307 B.n679 B.n50 585
R308 B.n783 B.n50 585
R309 B.n678 B.n49 585
R310 B.n784 B.n49 585
R311 B.n677 B.n48 585
R312 B.n785 B.n48 585
R313 B.n676 B.n675 585
R314 B.n675 B.n44 585
R315 B.n674 B.n43 585
R316 B.n791 B.n43 585
R317 B.n673 B.n42 585
R318 B.n792 B.n42 585
R319 B.n672 B.n41 585
R320 B.n793 B.n41 585
R321 B.n671 B.n670 585
R322 B.n670 B.n37 585
R323 B.n669 B.n36 585
R324 B.n799 B.n36 585
R325 B.n668 B.n35 585
R326 B.n800 B.n35 585
R327 B.n667 B.n34 585
R328 B.n801 B.n34 585
R329 B.n666 B.n665 585
R330 B.n665 B.n30 585
R331 B.n664 B.n29 585
R332 B.n807 B.n29 585
R333 B.n663 B.n28 585
R334 B.n808 B.n28 585
R335 B.n662 B.n27 585
R336 B.n809 B.n27 585
R337 B.n661 B.n660 585
R338 B.n660 B.n23 585
R339 B.n659 B.n22 585
R340 B.n815 B.n22 585
R341 B.n658 B.n21 585
R342 B.n816 B.n21 585
R343 B.n657 B.n20 585
R344 B.n817 B.n20 585
R345 B.n656 B.n655 585
R346 B.n655 B.n16 585
R347 B.n654 B.n15 585
R348 B.n823 B.n15 585
R349 B.n653 B.n14 585
R350 B.n824 B.n14 585
R351 B.n652 B.n13 585
R352 B.n825 B.n13 585
R353 B.n651 B.n650 585
R354 B.n650 B.n12 585
R355 B.n649 B.n648 585
R356 B.n649 B.n8 585
R357 B.n647 B.n7 585
R358 B.n832 B.n7 585
R359 B.n646 B.n6 585
R360 B.n833 B.n6 585
R361 B.n645 B.n5 585
R362 B.n834 B.n5 585
R363 B.n644 B.n643 585
R364 B.n643 B.n4 585
R365 B.n642 B.n234 585
R366 B.n642 B.n641 585
R367 B.n632 B.n235 585
R368 B.n236 B.n235 585
R369 B.n634 B.n633 585
R370 B.n635 B.n634 585
R371 B.n631 B.n241 585
R372 B.n241 B.n240 585
R373 B.n630 B.n629 585
R374 B.n629 B.n628 585
R375 B.n243 B.n242 585
R376 B.n244 B.n243 585
R377 B.n621 B.n620 585
R378 B.n622 B.n621 585
R379 B.n619 B.n249 585
R380 B.n249 B.n248 585
R381 B.n618 B.n617 585
R382 B.n617 B.n616 585
R383 B.n251 B.n250 585
R384 B.n252 B.n251 585
R385 B.n609 B.n608 585
R386 B.n610 B.n609 585
R387 B.n607 B.n257 585
R388 B.n257 B.n256 585
R389 B.n606 B.n605 585
R390 B.n605 B.n604 585
R391 B.n259 B.n258 585
R392 B.n260 B.n259 585
R393 B.n597 B.n596 585
R394 B.n598 B.n597 585
R395 B.n595 B.n265 585
R396 B.n265 B.n264 585
R397 B.n594 B.n593 585
R398 B.n593 B.n592 585
R399 B.n267 B.n266 585
R400 B.n268 B.n267 585
R401 B.n585 B.n584 585
R402 B.n586 B.n585 585
R403 B.n583 B.n273 585
R404 B.n273 B.n272 585
R405 B.n582 B.n581 585
R406 B.n581 B.n580 585
R407 B.n275 B.n274 585
R408 B.n276 B.n275 585
R409 B.n573 B.n572 585
R410 B.n574 B.n573 585
R411 B.n571 B.n281 585
R412 B.n281 B.n280 585
R413 B.n570 B.n569 585
R414 B.n569 B.n568 585
R415 B.n283 B.n282 585
R416 B.n284 B.n283 585
R417 B.n561 B.n560 585
R418 B.n562 B.n561 585
R419 B.n559 B.n289 585
R420 B.n289 B.n288 585
R421 B.n558 B.n557 585
R422 B.n557 B.n556 585
R423 B.n291 B.n290 585
R424 B.n292 B.n291 585
R425 B.n549 B.n548 585
R426 B.n550 B.n549 585
R427 B.n547 B.n297 585
R428 B.n297 B.n296 585
R429 B.n546 B.n545 585
R430 B.n545 B.n544 585
R431 B.n299 B.n298 585
R432 B.n300 B.n299 585
R433 B.n537 B.n536 585
R434 B.n538 B.n537 585
R435 B.n535 B.n305 585
R436 B.n305 B.n304 585
R437 B.n534 B.n533 585
R438 B.n533 B.n532 585
R439 B.n307 B.n306 585
R440 B.n308 B.n307 585
R441 B.n525 B.n524 585
R442 B.n526 B.n525 585
R443 B.n523 B.n313 585
R444 B.n313 B.n312 585
R445 B.n522 B.n521 585
R446 B.n521 B.n520 585
R447 B.n315 B.n314 585
R448 B.n316 B.n315 585
R449 B.n513 B.n512 585
R450 B.n514 B.n513 585
R451 B.n511 B.n321 585
R452 B.n321 B.n320 585
R453 B.n510 B.n509 585
R454 B.n509 B.n508 585
R455 B.n323 B.n322 585
R456 B.n324 B.n323 585
R457 B.n501 B.n500 585
R458 B.n502 B.n501 585
R459 B.n499 B.n328 585
R460 B.n332 B.n328 585
R461 B.n498 B.n497 585
R462 B.n497 B.n496 585
R463 B.n330 B.n329 585
R464 B.n331 B.n330 585
R465 B.n489 B.n488 585
R466 B.n490 B.n489 585
R467 B.n487 B.n337 585
R468 B.n337 B.n336 585
R469 B.n486 B.n485 585
R470 B.n485 B.n484 585
R471 B.n339 B.n338 585
R472 B.n340 B.n339 585
R473 B.n477 B.n476 585
R474 B.n478 B.n477 585
R475 B.n343 B.n342 585
R476 B.n377 B.n376 585
R477 B.n378 B.n374 585
R478 B.n374 B.n344 585
R479 B.n380 B.n379 585
R480 B.n382 B.n373 585
R481 B.n385 B.n384 585
R482 B.n386 B.n372 585
R483 B.n388 B.n387 585
R484 B.n390 B.n371 585
R485 B.n393 B.n392 585
R486 B.n394 B.n370 585
R487 B.n396 B.n395 585
R488 B.n398 B.n369 585
R489 B.n401 B.n400 585
R490 B.n402 B.n368 585
R491 B.n404 B.n403 585
R492 B.n406 B.n367 585
R493 B.n409 B.n408 585
R494 B.n410 B.n366 585
R495 B.n412 B.n411 585
R496 B.n414 B.n365 585
R497 B.n417 B.n416 585
R498 B.n418 B.n361 585
R499 B.n420 B.n419 585
R500 B.n422 B.n360 585
R501 B.n425 B.n424 585
R502 B.n426 B.n359 585
R503 B.n428 B.n427 585
R504 B.n430 B.n358 585
R505 B.n433 B.n432 585
R506 B.n435 B.n355 585
R507 B.n437 B.n436 585
R508 B.n439 B.n354 585
R509 B.n442 B.n441 585
R510 B.n443 B.n353 585
R511 B.n445 B.n444 585
R512 B.n447 B.n352 585
R513 B.n450 B.n449 585
R514 B.n451 B.n351 585
R515 B.n453 B.n452 585
R516 B.n455 B.n350 585
R517 B.n458 B.n457 585
R518 B.n459 B.n349 585
R519 B.n461 B.n460 585
R520 B.n463 B.n348 585
R521 B.n466 B.n465 585
R522 B.n467 B.n347 585
R523 B.n469 B.n468 585
R524 B.n471 B.n346 585
R525 B.n474 B.n473 585
R526 B.n475 B.n345 585
R527 B.n480 B.n479 585
R528 B.n479 B.n478 585
R529 B.n481 B.n341 585
R530 B.n341 B.n340 585
R531 B.n483 B.n482 585
R532 B.n484 B.n483 585
R533 B.n335 B.n334 585
R534 B.n336 B.n335 585
R535 B.n492 B.n491 585
R536 B.n491 B.n490 585
R537 B.n493 B.n333 585
R538 B.n333 B.n331 585
R539 B.n495 B.n494 585
R540 B.n496 B.n495 585
R541 B.n327 B.n326 585
R542 B.n332 B.n327 585
R543 B.n504 B.n503 585
R544 B.n503 B.n502 585
R545 B.n505 B.n325 585
R546 B.n325 B.n324 585
R547 B.n507 B.n506 585
R548 B.n508 B.n507 585
R549 B.n319 B.n318 585
R550 B.n320 B.n319 585
R551 B.n516 B.n515 585
R552 B.n515 B.n514 585
R553 B.n517 B.n317 585
R554 B.n317 B.n316 585
R555 B.n519 B.n518 585
R556 B.n520 B.n519 585
R557 B.n311 B.n310 585
R558 B.n312 B.n311 585
R559 B.n528 B.n527 585
R560 B.n527 B.n526 585
R561 B.n529 B.n309 585
R562 B.n309 B.n308 585
R563 B.n531 B.n530 585
R564 B.n532 B.n531 585
R565 B.n303 B.n302 585
R566 B.n304 B.n303 585
R567 B.n540 B.n539 585
R568 B.n539 B.n538 585
R569 B.n541 B.n301 585
R570 B.n301 B.n300 585
R571 B.n543 B.n542 585
R572 B.n544 B.n543 585
R573 B.n295 B.n294 585
R574 B.n296 B.n295 585
R575 B.n552 B.n551 585
R576 B.n551 B.n550 585
R577 B.n553 B.n293 585
R578 B.n293 B.n292 585
R579 B.n555 B.n554 585
R580 B.n556 B.n555 585
R581 B.n287 B.n286 585
R582 B.n288 B.n287 585
R583 B.n564 B.n563 585
R584 B.n563 B.n562 585
R585 B.n565 B.n285 585
R586 B.n285 B.n284 585
R587 B.n567 B.n566 585
R588 B.n568 B.n567 585
R589 B.n279 B.n278 585
R590 B.n280 B.n279 585
R591 B.n576 B.n575 585
R592 B.n575 B.n574 585
R593 B.n577 B.n277 585
R594 B.n277 B.n276 585
R595 B.n579 B.n578 585
R596 B.n580 B.n579 585
R597 B.n271 B.n270 585
R598 B.n272 B.n271 585
R599 B.n588 B.n587 585
R600 B.n587 B.n586 585
R601 B.n589 B.n269 585
R602 B.n269 B.n268 585
R603 B.n591 B.n590 585
R604 B.n592 B.n591 585
R605 B.n263 B.n262 585
R606 B.n264 B.n263 585
R607 B.n600 B.n599 585
R608 B.n599 B.n598 585
R609 B.n601 B.n261 585
R610 B.n261 B.n260 585
R611 B.n603 B.n602 585
R612 B.n604 B.n603 585
R613 B.n255 B.n254 585
R614 B.n256 B.n255 585
R615 B.n612 B.n611 585
R616 B.n611 B.n610 585
R617 B.n613 B.n253 585
R618 B.n253 B.n252 585
R619 B.n615 B.n614 585
R620 B.n616 B.n615 585
R621 B.n247 B.n246 585
R622 B.n248 B.n247 585
R623 B.n624 B.n623 585
R624 B.n623 B.n622 585
R625 B.n625 B.n245 585
R626 B.n245 B.n244 585
R627 B.n627 B.n626 585
R628 B.n628 B.n627 585
R629 B.n239 B.n238 585
R630 B.n240 B.n239 585
R631 B.n637 B.n636 585
R632 B.n636 B.n635 585
R633 B.n638 B.n237 585
R634 B.n237 B.n236 585
R635 B.n640 B.n639 585
R636 B.n641 B.n640 585
R637 B.n3 B.n0 585
R638 B.n4 B.n3 585
R639 B.n831 B.n1 585
R640 B.n832 B.n831 585
R641 B.n830 B.n829 585
R642 B.n830 B.n8 585
R643 B.n828 B.n9 585
R644 B.n12 B.n9 585
R645 B.n827 B.n826 585
R646 B.n826 B.n825 585
R647 B.n11 B.n10 585
R648 B.n824 B.n11 585
R649 B.n822 B.n821 585
R650 B.n823 B.n822 585
R651 B.n820 B.n17 585
R652 B.n17 B.n16 585
R653 B.n819 B.n818 585
R654 B.n818 B.n817 585
R655 B.n19 B.n18 585
R656 B.n816 B.n19 585
R657 B.n814 B.n813 585
R658 B.n815 B.n814 585
R659 B.n812 B.n24 585
R660 B.n24 B.n23 585
R661 B.n811 B.n810 585
R662 B.n810 B.n809 585
R663 B.n26 B.n25 585
R664 B.n808 B.n26 585
R665 B.n806 B.n805 585
R666 B.n807 B.n806 585
R667 B.n804 B.n31 585
R668 B.n31 B.n30 585
R669 B.n803 B.n802 585
R670 B.n802 B.n801 585
R671 B.n33 B.n32 585
R672 B.n800 B.n33 585
R673 B.n798 B.n797 585
R674 B.n799 B.n798 585
R675 B.n796 B.n38 585
R676 B.n38 B.n37 585
R677 B.n795 B.n794 585
R678 B.n794 B.n793 585
R679 B.n40 B.n39 585
R680 B.n792 B.n40 585
R681 B.n790 B.n789 585
R682 B.n791 B.n790 585
R683 B.n788 B.n45 585
R684 B.n45 B.n44 585
R685 B.n787 B.n786 585
R686 B.n786 B.n785 585
R687 B.n47 B.n46 585
R688 B.n784 B.n47 585
R689 B.n782 B.n781 585
R690 B.n783 B.n782 585
R691 B.n780 B.n52 585
R692 B.n52 B.n51 585
R693 B.n779 B.n778 585
R694 B.n778 B.n777 585
R695 B.n54 B.n53 585
R696 B.n776 B.n54 585
R697 B.n774 B.n773 585
R698 B.n775 B.n774 585
R699 B.n772 B.n59 585
R700 B.n59 B.n58 585
R701 B.n771 B.n770 585
R702 B.n770 B.n769 585
R703 B.n61 B.n60 585
R704 B.n768 B.n61 585
R705 B.n766 B.n765 585
R706 B.n767 B.n766 585
R707 B.n764 B.n66 585
R708 B.n66 B.n65 585
R709 B.n763 B.n762 585
R710 B.n762 B.n761 585
R711 B.n68 B.n67 585
R712 B.n760 B.n68 585
R713 B.n758 B.n757 585
R714 B.n759 B.n758 585
R715 B.n756 B.n73 585
R716 B.n73 B.n72 585
R717 B.n755 B.n754 585
R718 B.n754 B.n753 585
R719 B.n75 B.n74 585
R720 B.n752 B.n75 585
R721 B.n750 B.n749 585
R722 B.n751 B.n750 585
R723 B.n748 B.n80 585
R724 B.n80 B.n79 585
R725 B.n747 B.n746 585
R726 B.n746 B.n745 585
R727 B.n82 B.n81 585
R728 B.n744 B.n82 585
R729 B.n742 B.n741 585
R730 B.n743 B.n742 585
R731 B.n740 B.n87 585
R732 B.n87 B.n86 585
R733 B.n739 B.n738 585
R734 B.n738 B.n737 585
R735 B.n89 B.n88 585
R736 B.n736 B.n89 585
R737 B.n734 B.n733 585
R738 B.n735 B.n734 585
R739 B.n732 B.n94 585
R740 B.n94 B.n93 585
R741 B.n731 B.n730 585
R742 B.n730 B.n729 585
R743 B.n96 B.n95 585
R744 B.n728 B.n96 585
R745 B.n726 B.n725 585
R746 B.n727 B.n726 585
R747 B.n724 B.n101 585
R748 B.n101 B.n100 585
R749 B.n723 B.n722 585
R750 B.n722 B.n721 585
R751 B.n835 B.n834 585
R752 B.n833 B.n2 585
R753 B.n722 B.n103 550.159
R754 B.n719 B.n104 550.159
R755 B.n477 B.n345 550.159
R756 B.n479 B.n343 550.159
R757 B.n134 B.t10 257.053
R758 B.n131 B.t21 257.053
R759 B.n356 B.t14 257.053
R760 B.n362 B.t18 257.053
R761 B.n720 B.n129 256.663
R762 B.n720 B.n128 256.663
R763 B.n720 B.n127 256.663
R764 B.n720 B.n126 256.663
R765 B.n720 B.n125 256.663
R766 B.n720 B.n124 256.663
R767 B.n720 B.n123 256.663
R768 B.n720 B.n122 256.663
R769 B.n720 B.n121 256.663
R770 B.n720 B.n120 256.663
R771 B.n720 B.n119 256.663
R772 B.n720 B.n118 256.663
R773 B.n720 B.n117 256.663
R774 B.n720 B.n116 256.663
R775 B.n720 B.n115 256.663
R776 B.n720 B.n114 256.663
R777 B.n720 B.n113 256.663
R778 B.n720 B.n112 256.663
R779 B.n720 B.n111 256.663
R780 B.n720 B.n110 256.663
R781 B.n720 B.n109 256.663
R782 B.n720 B.n108 256.663
R783 B.n720 B.n107 256.663
R784 B.n720 B.n106 256.663
R785 B.n720 B.n105 256.663
R786 B.n375 B.n344 256.663
R787 B.n381 B.n344 256.663
R788 B.n383 B.n344 256.663
R789 B.n389 B.n344 256.663
R790 B.n391 B.n344 256.663
R791 B.n397 B.n344 256.663
R792 B.n399 B.n344 256.663
R793 B.n405 B.n344 256.663
R794 B.n407 B.n344 256.663
R795 B.n413 B.n344 256.663
R796 B.n415 B.n344 256.663
R797 B.n421 B.n344 256.663
R798 B.n423 B.n344 256.663
R799 B.n429 B.n344 256.663
R800 B.n431 B.n344 256.663
R801 B.n438 B.n344 256.663
R802 B.n440 B.n344 256.663
R803 B.n446 B.n344 256.663
R804 B.n448 B.n344 256.663
R805 B.n454 B.n344 256.663
R806 B.n456 B.n344 256.663
R807 B.n462 B.n344 256.663
R808 B.n464 B.n344 256.663
R809 B.n470 B.n344 256.663
R810 B.n472 B.n344 256.663
R811 B.n837 B.n836 256.663
R812 B.n138 B.n137 163.367
R813 B.n142 B.n141 163.367
R814 B.n146 B.n145 163.367
R815 B.n150 B.n149 163.367
R816 B.n154 B.n153 163.367
R817 B.n158 B.n157 163.367
R818 B.n162 B.n161 163.367
R819 B.n166 B.n165 163.367
R820 B.n170 B.n169 163.367
R821 B.n174 B.n173 163.367
R822 B.n179 B.n178 163.367
R823 B.n183 B.n182 163.367
R824 B.n187 B.n186 163.367
R825 B.n191 B.n190 163.367
R826 B.n195 B.n194 163.367
R827 B.n199 B.n198 163.367
R828 B.n203 B.n202 163.367
R829 B.n207 B.n206 163.367
R830 B.n211 B.n210 163.367
R831 B.n215 B.n214 163.367
R832 B.n219 B.n218 163.367
R833 B.n223 B.n222 163.367
R834 B.n227 B.n226 163.367
R835 B.n231 B.n230 163.367
R836 B.n719 B.n130 163.367
R837 B.n477 B.n339 163.367
R838 B.n485 B.n339 163.367
R839 B.n485 B.n337 163.367
R840 B.n489 B.n337 163.367
R841 B.n489 B.n330 163.367
R842 B.n497 B.n330 163.367
R843 B.n497 B.n328 163.367
R844 B.n501 B.n328 163.367
R845 B.n501 B.n323 163.367
R846 B.n509 B.n323 163.367
R847 B.n509 B.n321 163.367
R848 B.n513 B.n321 163.367
R849 B.n513 B.n315 163.367
R850 B.n521 B.n315 163.367
R851 B.n521 B.n313 163.367
R852 B.n525 B.n313 163.367
R853 B.n525 B.n307 163.367
R854 B.n533 B.n307 163.367
R855 B.n533 B.n305 163.367
R856 B.n537 B.n305 163.367
R857 B.n537 B.n299 163.367
R858 B.n545 B.n299 163.367
R859 B.n545 B.n297 163.367
R860 B.n549 B.n297 163.367
R861 B.n549 B.n291 163.367
R862 B.n557 B.n291 163.367
R863 B.n557 B.n289 163.367
R864 B.n561 B.n289 163.367
R865 B.n561 B.n283 163.367
R866 B.n569 B.n283 163.367
R867 B.n569 B.n281 163.367
R868 B.n573 B.n281 163.367
R869 B.n573 B.n275 163.367
R870 B.n581 B.n275 163.367
R871 B.n581 B.n273 163.367
R872 B.n585 B.n273 163.367
R873 B.n585 B.n267 163.367
R874 B.n593 B.n267 163.367
R875 B.n593 B.n265 163.367
R876 B.n597 B.n265 163.367
R877 B.n597 B.n259 163.367
R878 B.n605 B.n259 163.367
R879 B.n605 B.n257 163.367
R880 B.n609 B.n257 163.367
R881 B.n609 B.n251 163.367
R882 B.n617 B.n251 163.367
R883 B.n617 B.n249 163.367
R884 B.n621 B.n249 163.367
R885 B.n621 B.n243 163.367
R886 B.n629 B.n243 163.367
R887 B.n629 B.n241 163.367
R888 B.n634 B.n241 163.367
R889 B.n634 B.n235 163.367
R890 B.n642 B.n235 163.367
R891 B.n643 B.n642 163.367
R892 B.n643 B.n5 163.367
R893 B.n6 B.n5 163.367
R894 B.n7 B.n6 163.367
R895 B.n649 B.n7 163.367
R896 B.n650 B.n649 163.367
R897 B.n650 B.n13 163.367
R898 B.n14 B.n13 163.367
R899 B.n15 B.n14 163.367
R900 B.n655 B.n15 163.367
R901 B.n655 B.n20 163.367
R902 B.n21 B.n20 163.367
R903 B.n22 B.n21 163.367
R904 B.n660 B.n22 163.367
R905 B.n660 B.n27 163.367
R906 B.n28 B.n27 163.367
R907 B.n29 B.n28 163.367
R908 B.n665 B.n29 163.367
R909 B.n665 B.n34 163.367
R910 B.n35 B.n34 163.367
R911 B.n36 B.n35 163.367
R912 B.n670 B.n36 163.367
R913 B.n670 B.n41 163.367
R914 B.n42 B.n41 163.367
R915 B.n43 B.n42 163.367
R916 B.n675 B.n43 163.367
R917 B.n675 B.n48 163.367
R918 B.n49 B.n48 163.367
R919 B.n50 B.n49 163.367
R920 B.n680 B.n50 163.367
R921 B.n680 B.n55 163.367
R922 B.n56 B.n55 163.367
R923 B.n57 B.n56 163.367
R924 B.n685 B.n57 163.367
R925 B.n685 B.n62 163.367
R926 B.n63 B.n62 163.367
R927 B.n64 B.n63 163.367
R928 B.n690 B.n64 163.367
R929 B.n690 B.n69 163.367
R930 B.n70 B.n69 163.367
R931 B.n71 B.n70 163.367
R932 B.n695 B.n71 163.367
R933 B.n695 B.n76 163.367
R934 B.n77 B.n76 163.367
R935 B.n78 B.n77 163.367
R936 B.n700 B.n78 163.367
R937 B.n700 B.n83 163.367
R938 B.n84 B.n83 163.367
R939 B.n85 B.n84 163.367
R940 B.n705 B.n85 163.367
R941 B.n705 B.n90 163.367
R942 B.n91 B.n90 163.367
R943 B.n92 B.n91 163.367
R944 B.n710 B.n92 163.367
R945 B.n710 B.n97 163.367
R946 B.n98 B.n97 163.367
R947 B.n99 B.n98 163.367
R948 B.n715 B.n99 163.367
R949 B.n715 B.n104 163.367
R950 B.n376 B.n374 163.367
R951 B.n380 B.n374 163.367
R952 B.n384 B.n382 163.367
R953 B.n388 B.n372 163.367
R954 B.n392 B.n390 163.367
R955 B.n396 B.n370 163.367
R956 B.n400 B.n398 163.367
R957 B.n404 B.n368 163.367
R958 B.n408 B.n406 163.367
R959 B.n412 B.n366 163.367
R960 B.n416 B.n414 163.367
R961 B.n420 B.n361 163.367
R962 B.n424 B.n422 163.367
R963 B.n428 B.n359 163.367
R964 B.n432 B.n430 163.367
R965 B.n437 B.n355 163.367
R966 B.n441 B.n439 163.367
R967 B.n445 B.n353 163.367
R968 B.n449 B.n447 163.367
R969 B.n453 B.n351 163.367
R970 B.n457 B.n455 163.367
R971 B.n461 B.n349 163.367
R972 B.n465 B.n463 163.367
R973 B.n469 B.n347 163.367
R974 B.n473 B.n471 163.367
R975 B.n479 B.n341 163.367
R976 B.n483 B.n341 163.367
R977 B.n483 B.n335 163.367
R978 B.n491 B.n335 163.367
R979 B.n491 B.n333 163.367
R980 B.n495 B.n333 163.367
R981 B.n495 B.n327 163.367
R982 B.n503 B.n327 163.367
R983 B.n503 B.n325 163.367
R984 B.n507 B.n325 163.367
R985 B.n507 B.n319 163.367
R986 B.n515 B.n319 163.367
R987 B.n515 B.n317 163.367
R988 B.n519 B.n317 163.367
R989 B.n519 B.n311 163.367
R990 B.n527 B.n311 163.367
R991 B.n527 B.n309 163.367
R992 B.n531 B.n309 163.367
R993 B.n531 B.n303 163.367
R994 B.n539 B.n303 163.367
R995 B.n539 B.n301 163.367
R996 B.n543 B.n301 163.367
R997 B.n543 B.n295 163.367
R998 B.n551 B.n295 163.367
R999 B.n551 B.n293 163.367
R1000 B.n555 B.n293 163.367
R1001 B.n555 B.n287 163.367
R1002 B.n563 B.n287 163.367
R1003 B.n563 B.n285 163.367
R1004 B.n567 B.n285 163.367
R1005 B.n567 B.n279 163.367
R1006 B.n575 B.n279 163.367
R1007 B.n575 B.n277 163.367
R1008 B.n579 B.n277 163.367
R1009 B.n579 B.n271 163.367
R1010 B.n587 B.n271 163.367
R1011 B.n587 B.n269 163.367
R1012 B.n591 B.n269 163.367
R1013 B.n591 B.n263 163.367
R1014 B.n599 B.n263 163.367
R1015 B.n599 B.n261 163.367
R1016 B.n603 B.n261 163.367
R1017 B.n603 B.n255 163.367
R1018 B.n611 B.n255 163.367
R1019 B.n611 B.n253 163.367
R1020 B.n615 B.n253 163.367
R1021 B.n615 B.n247 163.367
R1022 B.n623 B.n247 163.367
R1023 B.n623 B.n245 163.367
R1024 B.n627 B.n245 163.367
R1025 B.n627 B.n239 163.367
R1026 B.n636 B.n239 163.367
R1027 B.n636 B.n237 163.367
R1028 B.n640 B.n237 163.367
R1029 B.n640 B.n3 163.367
R1030 B.n835 B.n3 163.367
R1031 B.n831 B.n2 163.367
R1032 B.n831 B.n830 163.367
R1033 B.n830 B.n9 163.367
R1034 B.n826 B.n9 163.367
R1035 B.n826 B.n11 163.367
R1036 B.n822 B.n11 163.367
R1037 B.n822 B.n17 163.367
R1038 B.n818 B.n17 163.367
R1039 B.n818 B.n19 163.367
R1040 B.n814 B.n19 163.367
R1041 B.n814 B.n24 163.367
R1042 B.n810 B.n24 163.367
R1043 B.n810 B.n26 163.367
R1044 B.n806 B.n26 163.367
R1045 B.n806 B.n31 163.367
R1046 B.n802 B.n31 163.367
R1047 B.n802 B.n33 163.367
R1048 B.n798 B.n33 163.367
R1049 B.n798 B.n38 163.367
R1050 B.n794 B.n38 163.367
R1051 B.n794 B.n40 163.367
R1052 B.n790 B.n40 163.367
R1053 B.n790 B.n45 163.367
R1054 B.n786 B.n45 163.367
R1055 B.n786 B.n47 163.367
R1056 B.n782 B.n47 163.367
R1057 B.n782 B.n52 163.367
R1058 B.n778 B.n52 163.367
R1059 B.n778 B.n54 163.367
R1060 B.n774 B.n54 163.367
R1061 B.n774 B.n59 163.367
R1062 B.n770 B.n59 163.367
R1063 B.n770 B.n61 163.367
R1064 B.n766 B.n61 163.367
R1065 B.n766 B.n66 163.367
R1066 B.n762 B.n66 163.367
R1067 B.n762 B.n68 163.367
R1068 B.n758 B.n68 163.367
R1069 B.n758 B.n73 163.367
R1070 B.n754 B.n73 163.367
R1071 B.n754 B.n75 163.367
R1072 B.n750 B.n75 163.367
R1073 B.n750 B.n80 163.367
R1074 B.n746 B.n80 163.367
R1075 B.n746 B.n82 163.367
R1076 B.n742 B.n82 163.367
R1077 B.n742 B.n87 163.367
R1078 B.n738 B.n87 163.367
R1079 B.n738 B.n89 163.367
R1080 B.n734 B.n89 163.367
R1081 B.n734 B.n94 163.367
R1082 B.n730 B.n94 163.367
R1083 B.n730 B.n96 163.367
R1084 B.n726 B.n96 163.367
R1085 B.n726 B.n101 163.367
R1086 B.n722 B.n101 163.367
R1087 B.n478 B.n344 143.082
R1088 B.n721 B.n720 143.082
R1089 B.n131 B.t22 127.246
R1090 B.n356 B.t17 127.246
R1091 B.n134 B.t12 127.242
R1092 B.n362 B.t20 127.242
R1093 B.n132 B.t23 73.9128
R1094 B.n357 B.t16 73.9128
R1095 B.n135 B.t13 73.9079
R1096 B.n363 B.t19 73.9079
R1097 B.n478 B.n340 73.1545
R1098 B.n484 B.n340 73.1545
R1099 B.n484 B.n336 73.1545
R1100 B.n490 B.n336 73.1545
R1101 B.n490 B.n331 73.1545
R1102 B.n496 B.n331 73.1545
R1103 B.n496 B.n332 73.1545
R1104 B.n502 B.n324 73.1545
R1105 B.n508 B.n324 73.1545
R1106 B.n508 B.n320 73.1545
R1107 B.n514 B.n320 73.1545
R1108 B.n514 B.n316 73.1545
R1109 B.n520 B.n316 73.1545
R1110 B.n520 B.n312 73.1545
R1111 B.n526 B.n312 73.1545
R1112 B.n526 B.n308 73.1545
R1113 B.n532 B.n308 73.1545
R1114 B.n538 B.n304 73.1545
R1115 B.n538 B.n300 73.1545
R1116 B.n544 B.n300 73.1545
R1117 B.n544 B.n296 73.1545
R1118 B.n550 B.n296 73.1545
R1119 B.n550 B.n292 73.1545
R1120 B.n556 B.n292 73.1545
R1121 B.n562 B.n288 73.1545
R1122 B.n562 B.n284 73.1545
R1123 B.n568 B.n284 73.1545
R1124 B.n568 B.n280 73.1545
R1125 B.n574 B.n280 73.1545
R1126 B.n574 B.n276 73.1545
R1127 B.n580 B.n276 73.1545
R1128 B.n586 B.n272 73.1545
R1129 B.n586 B.n268 73.1545
R1130 B.n592 B.n268 73.1545
R1131 B.n592 B.n264 73.1545
R1132 B.n598 B.n264 73.1545
R1133 B.n598 B.n260 73.1545
R1134 B.n604 B.n260 73.1545
R1135 B.n610 B.n256 73.1545
R1136 B.n610 B.n252 73.1545
R1137 B.n616 B.n252 73.1545
R1138 B.n616 B.n248 73.1545
R1139 B.n622 B.n248 73.1545
R1140 B.n622 B.n244 73.1545
R1141 B.n628 B.n244 73.1545
R1142 B.n635 B.n240 73.1545
R1143 B.n635 B.n236 73.1545
R1144 B.n641 B.n236 73.1545
R1145 B.n641 B.n4 73.1545
R1146 B.n834 B.n4 73.1545
R1147 B.n834 B.n833 73.1545
R1148 B.n833 B.n832 73.1545
R1149 B.n832 B.n8 73.1545
R1150 B.n12 B.n8 73.1545
R1151 B.n825 B.n12 73.1545
R1152 B.n825 B.n824 73.1545
R1153 B.n823 B.n16 73.1545
R1154 B.n817 B.n16 73.1545
R1155 B.n817 B.n816 73.1545
R1156 B.n816 B.n815 73.1545
R1157 B.n815 B.n23 73.1545
R1158 B.n809 B.n23 73.1545
R1159 B.n809 B.n808 73.1545
R1160 B.n807 B.n30 73.1545
R1161 B.n801 B.n30 73.1545
R1162 B.n801 B.n800 73.1545
R1163 B.n800 B.n799 73.1545
R1164 B.n799 B.n37 73.1545
R1165 B.n793 B.n37 73.1545
R1166 B.n793 B.n792 73.1545
R1167 B.n791 B.n44 73.1545
R1168 B.n785 B.n44 73.1545
R1169 B.n785 B.n784 73.1545
R1170 B.n784 B.n783 73.1545
R1171 B.n783 B.n51 73.1545
R1172 B.n777 B.n51 73.1545
R1173 B.n777 B.n776 73.1545
R1174 B.n775 B.n58 73.1545
R1175 B.n769 B.n58 73.1545
R1176 B.n769 B.n768 73.1545
R1177 B.n768 B.n767 73.1545
R1178 B.n767 B.n65 73.1545
R1179 B.n761 B.n65 73.1545
R1180 B.n761 B.n760 73.1545
R1181 B.n759 B.n72 73.1545
R1182 B.n753 B.n72 73.1545
R1183 B.n753 B.n752 73.1545
R1184 B.n752 B.n751 73.1545
R1185 B.n751 B.n79 73.1545
R1186 B.n745 B.n79 73.1545
R1187 B.n745 B.n744 73.1545
R1188 B.n744 B.n743 73.1545
R1189 B.n743 B.n86 73.1545
R1190 B.n737 B.n86 73.1545
R1191 B.n736 B.n735 73.1545
R1192 B.n735 B.n93 73.1545
R1193 B.n729 B.n93 73.1545
R1194 B.n729 B.n728 73.1545
R1195 B.n728 B.n727 73.1545
R1196 B.n727 B.n100 73.1545
R1197 B.n721 B.n100 73.1545
R1198 B.n105 B.n103 71.676
R1199 B.n138 B.n106 71.676
R1200 B.n142 B.n107 71.676
R1201 B.n146 B.n108 71.676
R1202 B.n150 B.n109 71.676
R1203 B.n154 B.n110 71.676
R1204 B.n158 B.n111 71.676
R1205 B.n162 B.n112 71.676
R1206 B.n166 B.n113 71.676
R1207 B.n170 B.n114 71.676
R1208 B.n174 B.n115 71.676
R1209 B.n179 B.n116 71.676
R1210 B.n183 B.n117 71.676
R1211 B.n187 B.n118 71.676
R1212 B.n191 B.n119 71.676
R1213 B.n195 B.n120 71.676
R1214 B.n199 B.n121 71.676
R1215 B.n203 B.n122 71.676
R1216 B.n207 B.n123 71.676
R1217 B.n211 B.n124 71.676
R1218 B.n215 B.n125 71.676
R1219 B.n219 B.n126 71.676
R1220 B.n223 B.n127 71.676
R1221 B.n227 B.n128 71.676
R1222 B.n231 B.n129 71.676
R1223 B.n130 B.n129 71.676
R1224 B.n230 B.n128 71.676
R1225 B.n226 B.n127 71.676
R1226 B.n222 B.n126 71.676
R1227 B.n218 B.n125 71.676
R1228 B.n214 B.n124 71.676
R1229 B.n210 B.n123 71.676
R1230 B.n206 B.n122 71.676
R1231 B.n202 B.n121 71.676
R1232 B.n198 B.n120 71.676
R1233 B.n194 B.n119 71.676
R1234 B.n190 B.n118 71.676
R1235 B.n186 B.n117 71.676
R1236 B.n182 B.n116 71.676
R1237 B.n178 B.n115 71.676
R1238 B.n173 B.n114 71.676
R1239 B.n169 B.n113 71.676
R1240 B.n165 B.n112 71.676
R1241 B.n161 B.n111 71.676
R1242 B.n157 B.n110 71.676
R1243 B.n153 B.n109 71.676
R1244 B.n149 B.n108 71.676
R1245 B.n145 B.n107 71.676
R1246 B.n141 B.n106 71.676
R1247 B.n137 B.n105 71.676
R1248 B.n375 B.n343 71.676
R1249 B.n381 B.n380 71.676
R1250 B.n384 B.n383 71.676
R1251 B.n389 B.n388 71.676
R1252 B.n392 B.n391 71.676
R1253 B.n397 B.n396 71.676
R1254 B.n400 B.n399 71.676
R1255 B.n405 B.n404 71.676
R1256 B.n408 B.n407 71.676
R1257 B.n413 B.n412 71.676
R1258 B.n416 B.n415 71.676
R1259 B.n421 B.n420 71.676
R1260 B.n424 B.n423 71.676
R1261 B.n429 B.n428 71.676
R1262 B.n432 B.n431 71.676
R1263 B.n438 B.n437 71.676
R1264 B.n441 B.n440 71.676
R1265 B.n446 B.n445 71.676
R1266 B.n449 B.n448 71.676
R1267 B.n454 B.n453 71.676
R1268 B.n457 B.n456 71.676
R1269 B.n462 B.n461 71.676
R1270 B.n465 B.n464 71.676
R1271 B.n470 B.n469 71.676
R1272 B.n473 B.n472 71.676
R1273 B.n376 B.n375 71.676
R1274 B.n382 B.n381 71.676
R1275 B.n383 B.n372 71.676
R1276 B.n390 B.n389 71.676
R1277 B.n391 B.n370 71.676
R1278 B.n398 B.n397 71.676
R1279 B.n399 B.n368 71.676
R1280 B.n406 B.n405 71.676
R1281 B.n407 B.n366 71.676
R1282 B.n414 B.n413 71.676
R1283 B.n415 B.n361 71.676
R1284 B.n422 B.n421 71.676
R1285 B.n423 B.n359 71.676
R1286 B.n430 B.n429 71.676
R1287 B.n431 B.n355 71.676
R1288 B.n439 B.n438 71.676
R1289 B.n440 B.n353 71.676
R1290 B.n447 B.n446 71.676
R1291 B.n448 B.n351 71.676
R1292 B.n455 B.n454 71.676
R1293 B.n456 B.n349 71.676
R1294 B.n463 B.n462 71.676
R1295 B.n464 B.n347 71.676
R1296 B.n471 B.n470 71.676
R1297 B.n472 B.n345 71.676
R1298 B.n836 B.n835 71.676
R1299 B.n836 B.n2 71.676
R1300 B.n628 B.t7 62.3966
R1301 B.t5 B.n823 62.3966
R1302 B.n176 B.n135 59.5399
R1303 B.n133 B.n132 59.5399
R1304 B.n434 B.n357 59.5399
R1305 B.n364 B.n363 59.5399
R1306 B.n502 B.t15 58.0934
R1307 B.n737 B.t11 58.0934
R1308 B.n604 B.t9 55.9418
R1309 B.t6 B.n807 55.9418
R1310 B.n135 B.n134 53.3338
R1311 B.n132 B.n131 53.3338
R1312 B.n357 B.n356 53.3338
R1313 B.n363 B.n362 53.3338
R1314 B.n580 B.t4 49.487
R1315 B.t3 B.n791 49.487
R1316 B.n556 B.t8 43.0323
R1317 B.t0 B.n775 43.0323
R1318 B.n532 B.t2 36.5775
R1319 B.t2 B.n304 36.5775
R1320 B.n760 B.t1 36.5775
R1321 B.t1 B.n759 36.5775
R1322 B.n480 B.n342 35.7468
R1323 B.n476 B.n475 35.7468
R1324 B.n723 B.n102 35.7468
R1325 B.n718 B.n717 35.7468
R1326 B.t8 B.n288 30.1227
R1327 B.n776 B.t0 30.1227
R1328 B.t4 B.n272 23.668
R1329 B.n792 B.t3 23.668
R1330 B B.n837 18.0485
R1331 B.t9 B.n256 17.2132
R1332 B.n808 B.t6 17.2132
R1333 B.n332 B.t15 15.0616
R1334 B.t11 B.n736 15.0616
R1335 B.t7 B.n240 10.7584
R1336 B.n824 B.t5 10.7584
R1337 B.n481 B.n480 10.6151
R1338 B.n482 B.n481 10.6151
R1339 B.n482 B.n334 10.6151
R1340 B.n492 B.n334 10.6151
R1341 B.n493 B.n492 10.6151
R1342 B.n494 B.n493 10.6151
R1343 B.n494 B.n326 10.6151
R1344 B.n504 B.n326 10.6151
R1345 B.n505 B.n504 10.6151
R1346 B.n506 B.n505 10.6151
R1347 B.n506 B.n318 10.6151
R1348 B.n516 B.n318 10.6151
R1349 B.n517 B.n516 10.6151
R1350 B.n518 B.n517 10.6151
R1351 B.n518 B.n310 10.6151
R1352 B.n528 B.n310 10.6151
R1353 B.n529 B.n528 10.6151
R1354 B.n530 B.n529 10.6151
R1355 B.n530 B.n302 10.6151
R1356 B.n540 B.n302 10.6151
R1357 B.n541 B.n540 10.6151
R1358 B.n542 B.n541 10.6151
R1359 B.n542 B.n294 10.6151
R1360 B.n552 B.n294 10.6151
R1361 B.n553 B.n552 10.6151
R1362 B.n554 B.n553 10.6151
R1363 B.n554 B.n286 10.6151
R1364 B.n564 B.n286 10.6151
R1365 B.n565 B.n564 10.6151
R1366 B.n566 B.n565 10.6151
R1367 B.n566 B.n278 10.6151
R1368 B.n576 B.n278 10.6151
R1369 B.n577 B.n576 10.6151
R1370 B.n578 B.n577 10.6151
R1371 B.n578 B.n270 10.6151
R1372 B.n588 B.n270 10.6151
R1373 B.n589 B.n588 10.6151
R1374 B.n590 B.n589 10.6151
R1375 B.n590 B.n262 10.6151
R1376 B.n600 B.n262 10.6151
R1377 B.n601 B.n600 10.6151
R1378 B.n602 B.n601 10.6151
R1379 B.n602 B.n254 10.6151
R1380 B.n612 B.n254 10.6151
R1381 B.n613 B.n612 10.6151
R1382 B.n614 B.n613 10.6151
R1383 B.n614 B.n246 10.6151
R1384 B.n624 B.n246 10.6151
R1385 B.n625 B.n624 10.6151
R1386 B.n626 B.n625 10.6151
R1387 B.n626 B.n238 10.6151
R1388 B.n637 B.n238 10.6151
R1389 B.n638 B.n637 10.6151
R1390 B.n639 B.n638 10.6151
R1391 B.n639 B.n0 10.6151
R1392 B.n377 B.n342 10.6151
R1393 B.n378 B.n377 10.6151
R1394 B.n379 B.n378 10.6151
R1395 B.n379 B.n373 10.6151
R1396 B.n385 B.n373 10.6151
R1397 B.n386 B.n385 10.6151
R1398 B.n387 B.n386 10.6151
R1399 B.n387 B.n371 10.6151
R1400 B.n393 B.n371 10.6151
R1401 B.n394 B.n393 10.6151
R1402 B.n395 B.n394 10.6151
R1403 B.n395 B.n369 10.6151
R1404 B.n401 B.n369 10.6151
R1405 B.n402 B.n401 10.6151
R1406 B.n403 B.n402 10.6151
R1407 B.n403 B.n367 10.6151
R1408 B.n409 B.n367 10.6151
R1409 B.n410 B.n409 10.6151
R1410 B.n411 B.n410 10.6151
R1411 B.n411 B.n365 10.6151
R1412 B.n418 B.n417 10.6151
R1413 B.n419 B.n418 10.6151
R1414 B.n419 B.n360 10.6151
R1415 B.n425 B.n360 10.6151
R1416 B.n426 B.n425 10.6151
R1417 B.n427 B.n426 10.6151
R1418 B.n427 B.n358 10.6151
R1419 B.n433 B.n358 10.6151
R1420 B.n436 B.n435 10.6151
R1421 B.n436 B.n354 10.6151
R1422 B.n442 B.n354 10.6151
R1423 B.n443 B.n442 10.6151
R1424 B.n444 B.n443 10.6151
R1425 B.n444 B.n352 10.6151
R1426 B.n450 B.n352 10.6151
R1427 B.n451 B.n450 10.6151
R1428 B.n452 B.n451 10.6151
R1429 B.n452 B.n350 10.6151
R1430 B.n458 B.n350 10.6151
R1431 B.n459 B.n458 10.6151
R1432 B.n460 B.n459 10.6151
R1433 B.n460 B.n348 10.6151
R1434 B.n466 B.n348 10.6151
R1435 B.n467 B.n466 10.6151
R1436 B.n468 B.n467 10.6151
R1437 B.n468 B.n346 10.6151
R1438 B.n474 B.n346 10.6151
R1439 B.n475 B.n474 10.6151
R1440 B.n476 B.n338 10.6151
R1441 B.n486 B.n338 10.6151
R1442 B.n487 B.n486 10.6151
R1443 B.n488 B.n487 10.6151
R1444 B.n488 B.n329 10.6151
R1445 B.n498 B.n329 10.6151
R1446 B.n499 B.n498 10.6151
R1447 B.n500 B.n499 10.6151
R1448 B.n500 B.n322 10.6151
R1449 B.n510 B.n322 10.6151
R1450 B.n511 B.n510 10.6151
R1451 B.n512 B.n511 10.6151
R1452 B.n512 B.n314 10.6151
R1453 B.n522 B.n314 10.6151
R1454 B.n523 B.n522 10.6151
R1455 B.n524 B.n523 10.6151
R1456 B.n524 B.n306 10.6151
R1457 B.n534 B.n306 10.6151
R1458 B.n535 B.n534 10.6151
R1459 B.n536 B.n535 10.6151
R1460 B.n536 B.n298 10.6151
R1461 B.n546 B.n298 10.6151
R1462 B.n547 B.n546 10.6151
R1463 B.n548 B.n547 10.6151
R1464 B.n548 B.n290 10.6151
R1465 B.n558 B.n290 10.6151
R1466 B.n559 B.n558 10.6151
R1467 B.n560 B.n559 10.6151
R1468 B.n560 B.n282 10.6151
R1469 B.n570 B.n282 10.6151
R1470 B.n571 B.n570 10.6151
R1471 B.n572 B.n571 10.6151
R1472 B.n572 B.n274 10.6151
R1473 B.n582 B.n274 10.6151
R1474 B.n583 B.n582 10.6151
R1475 B.n584 B.n583 10.6151
R1476 B.n584 B.n266 10.6151
R1477 B.n594 B.n266 10.6151
R1478 B.n595 B.n594 10.6151
R1479 B.n596 B.n595 10.6151
R1480 B.n596 B.n258 10.6151
R1481 B.n606 B.n258 10.6151
R1482 B.n607 B.n606 10.6151
R1483 B.n608 B.n607 10.6151
R1484 B.n608 B.n250 10.6151
R1485 B.n618 B.n250 10.6151
R1486 B.n619 B.n618 10.6151
R1487 B.n620 B.n619 10.6151
R1488 B.n620 B.n242 10.6151
R1489 B.n630 B.n242 10.6151
R1490 B.n631 B.n630 10.6151
R1491 B.n633 B.n631 10.6151
R1492 B.n633 B.n632 10.6151
R1493 B.n632 B.n234 10.6151
R1494 B.n644 B.n234 10.6151
R1495 B.n645 B.n644 10.6151
R1496 B.n646 B.n645 10.6151
R1497 B.n647 B.n646 10.6151
R1498 B.n648 B.n647 10.6151
R1499 B.n651 B.n648 10.6151
R1500 B.n652 B.n651 10.6151
R1501 B.n653 B.n652 10.6151
R1502 B.n654 B.n653 10.6151
R1503 B.n656 B.n654 10.6151
R1504 B.n657 B.n656 10.6151
R1505 B.n658 B.n657 10.6151
R1506 B.n659 B.n658 10.6151
R1507 B.n661 B.n659 10.6151
R1508 B.n662 B.n661 10.6151
R1509 B.n663 B.n662 10.6151
R1510 B.n664 B.n663 10.6151
R1511 B.n666 B.n664 10.6151
R1512 B.n667 B.n666 10.6151
R1513 B.n668 B.n667 10.6151
R1514 B.n669 B.n668 10.6151
R1515 B.n671 B.n669 10.6151
R1516 B.n672 B.n671 10.6151
R1517 B.n673 B.n672 10.6151
R1518 B.n674 B.n673 10.6151
R1519 B.n676 B.n674 10.6151
R1520 B.n677 B.n676 10.6151
R1521 B.n678 B.n677 10.6151
R1522 B.n679 B.n678 10.6151
R1523 B.n681 B.n679 10.6151
R1524 B.n682 B.n681 10.6151
R1525 B.n683 B.n682 10.6151
R1526 B.n684 B.n683 10.6151
R1527 B.n686 B.n684 10.6151
R1528 B.n687 B.n686 10.6151
R1529 B.n688 B.n687 10.6151
R1530 B.n689 B.n688 10.6151
R1531 B.n691 B.n689 10.6151
R1532 B.n692 B.n691 10.6151
R1533 B.n693 B.n692 10.6151
R1534 B.n694 B.n693 10.6151
R1535 B.n696 B.n694 10.6151
R1536 B.n697 B.n696 10.6151
R1537 B.n698 B.n697 10.6151
R1538 B.n699 B.n698 10.6151
R1539 B.n701 B.n699 10.6151
R1540 B.n702 B.n701 10.6151
R1541 B.n703 B.n702 10.6151
R1542 B.n704 B.n703 10.6151
R1543 B.n706 B.n704 10.6151
R1544 B.n707 B.n706 10.6151
R1545 B.n708 B.n707 10.6151
R1546 B.n709 B.n708 10.6151
R1547 B.n711 B.n709 10.6151
R1548 B.n712 B.n711 10.6151
R1549 B.n713 B.n712 10.6151
R1550 B.n714 B.n713 10.6151
R1551 B.n716 B.n714 10.6151
R1552 B.n717 B.n716 10.6151
R1553 B.n829 B.n1 10.6151
R1554 B.n829 B.n828 10.6151
R1555 B.n828 B.n827 10.6151
R1556 B.n827 B.n10 10.6151
R1557 B.n821 B.n10 10.6151
R1558 B.n821 B.n820 10.6151
R1559 B.n820 B.n819 10.6151
R1560 B.n819 B.n18 10.6151
R1561 B.n813 B.n18 10.6151
R1562 B.n813 B.n812 10.6151
R1563 B.n812 B.n811 10.6151
R1564 B.n811 B.n25 10.6151
R1565 B.n805 B.n25 10.6151
R1566 B.n805 B.n804 10.6151
R1567 B.n804 B.n803 10.6151
R1568 B.n803 B.n32 10.6151
R1569 B.n797 B.n32 10.6151
R1570 B.n797 B.n796 10.6151
R1571 B.n796 B.n795 10.6151
R1572 B.n795 B.n39 10.6151
R1573 B.n789 B.n39 10.6151
R1574 B.n789 B.n788 10.6151
R1575 B.n788 B.n787 10.6151
R1576 B.n787 B.n46 10.6151
R1577 B.n781 B.n46 10.6151
R1578 B.n781 B.n780 10.6151
R1579 B.n780 B.n779 10.6151
R1580 B.n779 B.n53 10.6151
R1581 B.n773 B.n53 10.6151
R1582 B.n773 B.n772 10.6151
R1583 B.n772 B.n771 10.6151
R1584 B.n771 B.n60 10.6151
R1585 B.n765 B.n60 10.6151
R1586 B.n765 B.n764 10.6151
R1587 B.n764 B.n763 10.6151
R1588 B.n763 B.n67 10.6151
R1589 B.n757 B.n67 10.6151
R1590 B.n757 B.n756 10.6151
R1591 B.n756 B.n755 10.6151
R1592 B.n755 B.n74 10.6151
R1593 B.n749 B.n74 10.6151
R1594 B.n749 B.n748 10.6151
R1595 B.n748 B.n747 10.6151
R1596 B.n747 B.n81 10.6151
R1597 B.n741 B.n81 10.6151
R1598 B.n741 B.n740 10.6151
R1599 B.n740 B.n739 10.6151
R1600 B.n739 B.n88 10.6151
R1601 B.n733 B.n88 10.6151
R1602 B.n733 B.n732 10.6151
R1603 B.n732 B.n731 10.6151
R1604 B.n731 B.n95 10.6151
R1605 B.n725 B.n95 10.6151
R1606 B.n725 B.n724 10.6151
R1607 B.n724 B.n723 10.6151
R1608 B.n136 B.n102 10.6151
R1609 B.n139 B.n136 10.6151
R1610 B.n140 B.n139 10.6151
R1611 B.n143 B.n140 10.6151
R1612 B.n144 B.n143 10.6151
R1613 B.n147 B.n144 10.6151
R1614 B.n148 B.n147 10.6151
R1615 B.n151 B.n148 10.6151
R1616 B.n152 B.n151 10.6151
R1617 B.n155 B.n152 10.6151
R1618 B.n156 B.n155 10.6151
R1619 B.n159 B.n156 10.6151
R1620 B.n160 B.n159 10.6151
R1621 B.n163 B.n160 10.6151
R1622 B.n164 B.n163 10.6151
R1623 B.n167 B.n164 10.6151
R1624 B.n168 B.n167 10.6151
R1625 B.n171 B.n168 10.6151
R1626 B.n172 B.n171 10.6151
R1627 B.n175 B.n172 10.6151
R1628 B.n180 B.n177 10.6151
R1629 B.n181 B.n180 10.6151
R1630 B.n184 B.n181 10.6151
R1631 B.n185 B.n184 10.6151
R1632 B.n188 B.n185 10.6151
R1633 B.n189 B.n188 10.6151
R1634 B.n192 B.n189 10.6151
R1635 B.n193 B.n192 10.6151
R1636 B.n197 B.n196 10.6151
R1637 B.n200 B.n197 10.6151
R1638 B.n201 B.n200 10.6151
R1639 B.n204 B.n201 10.6151
R1640 B.n205 B.n204 10.6151
R1641 B.n208 B.n205 10.6151
R1642 B.n209 B.n208 10.6151
R1643 B.n212 B.n209 10.6151
R1644 B.n213 B.n212 10.6151
R1645 B.n216 B.n213 10.6151
R1646 B.n217 B.n216 10.6151
R1647 B.n220 B.n217 10.6151
R1648 B.n221 B.n220 10.6151
R1649 B.n224 B.n221 10.6151
R1650 B.n225 B.n224 10.6151
R1651 B.n228 B.n225 10.6151
R1652 B.n229 B.n228 10.6151
R1653 B.n232 B.n229 10.6151
R1654 B.n233 B.n232 10.6151
R1655 B.n718 B.n233 10.6151
R1656 B.n837 B.n0 8.11757
R1657 B.n837 B.n1 8.11757
R1658 B.n417 B.n364 6.5566
R1659 B.n434 B.n433 6.5566
R1660 B.n177 B.n176 6.5566
R1661 B.n193 B.n133 6.5566
R1662 B.n365 B.n364 4.05904
R1663 B.n435 B.n434 4.05904
R1664 B.n176 B.n175 4.05904
R1665 B.n196 B.n133 4.05904
R1666 VN.n71 VN.n37 161.3
R1667 VN.n70 VN.n69 161.3
R1668 VN.n68 VN.n38 161.3
R1669 VN.n67 VN.n66 161.3
R1670 VN.n65 VN.n39 161.3
R1671 VN.n64 VN.n63 161.3
R1672 VN.n62 VN.n40 161.3
R1673 VN.n61 VN.n60 161.3
R1674 VN.n59 VN.n41 161.3
R1675 VN.n58 VN.n57 161.3
R1676 VN.n56 VN.n42 161.3
R1677 VN.n55 VN.n54 161.3
R1678 VN.n53 VN.n43 161.3
R1679 VN.n52 VN.n51 161.3
R1680 VN.n50 VN.n45 161.3
R1681 VN.n49 VN.n48 161.3
R1682 VN.n34 VN.n0 161.3
R1683 VN.n33 VN.n32 161.3
R1684 VN.n31 VN.n1 161.3
R1685 VN.n30 VN.n29 161.3
R1686 VN.n28 VN.n2 161.3
R1687 VN.n27 VN.n26 161.3
R1688 VN.n25 VN.n3 161.3
R1689 VN.n24 VN.n23 161.3
R1690 VN.n22 VN.n4 161.3
R1691 VN.n21 VN.n20 161.3
R1692 VN.n19 VN.n5 161.3
R1693 VN.n18 VN.n17 161.3
R1694 VN.n15 VN.n6 161.3
R1695 VN.n14 VN.n13 161.3
R1696 VN.n12 VN.n7 161.3
R1697 VN.n11 VN.n10 161.3
R1698 VN.n36 VN.n35 98.5229
R1699 VN.n73 VN.n72 98.5229
R1700 VN.n8 VN.t3 83.6784
R1701 VN.n46 VN.t4 83.6784
R1702 VN.n14 VN.n7 52.6342
R1703 VN.n23 VN.n22 52.6342
R1704 VN.n29 VN.n1 52.6342
R1705 VN.n52 VN.n45 52.6342
R1706 VN.n60 VN.n59 52.6342
R1707 VN.n66 VN.n38 52.6342
R1708 VN.n27 VN.t6 49.296
R1709 VN.n9 VN.t9 49.296
R1710 VN.n16 VN.t2 49.296
R1711 VN.n35 VN.t1 49.296
R1712 VN.n64 VN.t5 49.296
R1713 VN.n47 VN.t7 49.296
R1714 VN.n44 VN.t0 49.296
R1715 VN.n72 VN.t8 49.296
R1716 VN.n9 VN.n8 48.0049
R1717 VN.n47 VN.n46 48.0049
R1718 VN VN.n73 47.0853
R1719 VN.n15 VN.n14 28.3526
R1720 VN.n22 VN.n21 28.3526
R1721 VN.n33 VN.n1 28.3526
R1722 VN.n53 VN.n52 28.3526
R1723 VN.n59 VN.n58 28.3526
R1724 VN.n70 VN.n38 28.3526
R1725 VN.n10 VN.n9 24.4675
R1726 VN.n10 VN.n7 24.4675
R1727 VN.n17 VN.n15 24.4675
R1728 VN.n21 VN.n5 24.4675
R1729 VN.n23 VN.n3 24.4675
R1730 VN.n27 VN.n3 24.4675
R1731 VN.n28 VN.n27 24.4675
R1732 VN.n29 VN.n28 24.4675
R1733 VN.n34 VN.n33 24.4675
R1734 VN.n48 VN.n45 24.4675
R1735 VN.n48 VN.n47 24.4675
R1736 VN.n58 VN.n42 24.4675
R1737 VN.n54 VN.n53 24.4675
R1738 VN.n66 VN.n65 24.4675
R1739 VN.n65 VN.n64 24.4675
R1740 VN.n64 VN.n40 24.4675
R1741 VN.n60 VN.n40 24.4675
R1742 VN.n71 VN.n70 24.4675
R1743 VN.n17 VN.n16 12.234
R1744 VN.n16 VN.n5 12.234
R1745 VN.n35 VN.n34 12.234
R1746 VN.n44 VN.n42 12.234
R1747 VN.n54 VN.n44 12.234
R1748 VN.n72 VN.n71 12.234
R1749 VN.n49 VN.n46 6.69041
R1750 VN.n11 VN.n8 6.69041
R1751 VN.n73 VN.n37 0.278367
R1752 VN.n36 VN.n0 0.278367
R1753 VN.n69 VN.n37 0.189894
R1754 VN.n69 VN.n68 0.189894
R1755 VN.n68 VN.n67 0.189894
R1756 VN.n67 VN.n39 0.189894
R1757 VN.n63 VN.n39 0.189894
R1758 VN.n63 VN.n62 0.189894
R1759 VN.n62 VN.n61 0.189894
R1760 VN.n61 VN.n41 0.189894
R1761 VN.n57 VN.n41 0.189894
R1762 VN.n57 VN.n56 0.189894
R1763 VN.n56 VN.n55 0.189894
R1764 VN.n55 VN.n43 0.189894
R1765 VN.n51 VN.n43 0.189894
R1766 VN.n51 VN.n50 0.189894
R1767 VN.n50 VN.n49 0.189894
R1768 VN.n12 VN.n11 0.189894
R1769 VN.n13 VN.n12 0.189894
R1770 VN.n13 VN.n6 0.189894
R1771 VN.n18 VN.n6 0.189894
R1772 VN.n19 VN.n18 0.189894
R1773 VN.n20 VN.n19 0.189894
R1774 VN.n20 VN.n4 0.189894
R1775 VN.n24 VN.n4 0.189894
R1776 VN.n25 VN.n24 0.189894
R1777 VN.n26 VN.n25 0.189894
R1778 VN.n26 VN.n2 0.189894
R1779 VN.n30 VN.n2 0.189894
R1780 VN.n31 VN.n30 0.189894
R1781 VN.n32 VN.n31 0.189894
R1782 VN.n32 VN.n0 0.189894
R1783 VN VN.n36 0.153454
R1784 VDD2.n1 VDD2.t6 76.5194
R1785 VDD2.n4 VDD2.t1 74.1488
R1786 VDD2.n3 VDD2.n2 71.8713
R1787 VDD2 VDD2.n7 71.8686
R1788 VDD2.n6 VDD2.n5 70.1489
R1789 VDD2.n1 VDD2.n0 70.1487
R1790 VDD2.n4 VDD2.n3 39.2433
R1791 VDD2.n7 VDD2.t2 4.0005
R1792 VDD2.n7 VDD2.t5 4.0005
R1793 VDD2.n5 VDD2.t4 4.0005
R1794 VDD2.n5 VDD2.t9 4.0005
R1795 VDD2.n2 VDD2.t3 4.0005
R1796 VDD2.n2 VDD2.t8 4.0005
R1797 VDD2.n0 VDD2.t0 4.0005
R1798 VDD2.n0 VDD2.t7 4.0005
R1799 VDD2.n6 VDD2.n4 2.37119
R1800 VDD2 VDD2.n6 0.651362
R1801 VDD2.n3 VDD2.n1 0.537826
C0 VN VDD1 0.152945f
C1 VP VDD1 5.04202f
C2 VN VDD2 4.63765f
C3 VN VTAIL 5.71891f
C4 VP VDD2 0.564361f
C5 VP VTAIL 5.73309f
C6 VDD2 VDD1 2.05638f
C7 VTAIL VDD1 6.99975f
C8 VDD2 VTAIL 7.05104f
C9 VN VP 6.827721f
C10 VDD2 B 5.820929f
C11 VDD1 B 5.737153f
C12 VTAIL B 4.852513f
C13 VN B 16.5469f
C14 VP B 15.096876f
C15 VDD2.t6 B 1.09417f
C16 VDD2.t0 B 0.104502f
C17 VDD2.t7 B 0.104502f
C18 VDD2.n0 B 0.849781f
C19 VDD2.n1 B 0.93203f
C20 VDD2.t3 B 0.104502f
C21 VDD2.t8 B 0.104502f
C22 VDD2.n2 B 0.863588f
C23 VDD2.n3 B 2.54221f
C24 VDD2.t1 B 1.07921f
C25 VDD2.n4 B 2.65127f
C26 VDD2.t4 B 0.104502f
C27 VDD2.t9 B 0.104502f
C28 VDD2.n5 B 0.849784f
C29 VDD2.n6 B 0.472648f
C30 VDD2.t2 B 0.104502f
C31 VDD2.t5 B 0.104502f
C32 VDD2.n7 B 0.863551f
C33 VN.n0 B 0.033706f
C34 VN.t1 B 0.800464f
C35 VN.n1 B 0.026306f
C36 VN.n2 B 0.025566f
C37 VN.t6 B 0.800464f
C38 VN.n3 B 0.047648f
C39 VN.n4 B 0.025566f
C40 VN.n5 B 0.035886f
C41 VN.n6 B 0.025566f
C42 VN.n7 B 0.045634f
C43 VN.t3 B 0.990344f
C44 VN.n8 B 0.362658f
C45 VN.t9 B 0.800464f
C46 VN.n9 B 0.394143f
C47 VN.n10 B 0.047648f
C48 VN.n11 B 0.242498f
C49 VN.n12 B 0.025566f
C50 VN.n13 B 0.025566f
C51 VN.n14 B 0.026306f
C52 VN.n15 B 0.050356f
C53 VN.t2 B 0.800464f
C54 VN.n16 B 0.30961f
C55 VN.n17 B 0.035886f
C56 VN.n18 B 0.025566f
C57 VN.n19 B 0.025566f
C58 VN.n20 B 0.025566f
C59 VN.n21 B 0.050356f
C60 VN.n22 B 0.026306f
C61 VN.n23 B 0.045634f
C62 VN.n24 B 0.025566f
C63 VN.n25 B 0.025566f
C64 VN.n26 B 0.025566f
C65 VN.n27 B 0.333734f
C66 VN.n28 B 0.047648f
C67 VN.n29 B 0.045634f
C68 VN.n30 B 0.025566f
C69 VN.n31 B 0.025566f
C70 VN.n32 B 0.025566f
C71 VN.n33 B 0.050356f
C72 VN.n34 B 0.035886f
C73 VN.n35 B 0.392303f
C74 VN.n36 B 0.038741f
C75 VN.n37 B 0.033706f
C76 VN.t8 B 0.800464f
C77 VN.n38 B 0.026306f
C78 VN.n39 B 0.025566f
C79 VN.t5 B 0.800464f
C80 VN.n40 B 0.047648f
C81 VN.n41 B 0.025566f
C82 VN.n42 B 0.035886f
C83 VN.n43 B 0.025566f
C84 VN.t0 B 0.800464f
C85 VN.n44 B 0.30961f
C86 VN.n45 B 0.045634f
C87 VN.t4 B 0.990344f
C88 VN.n46 B 0.362658f
C89 VN.t7 B 0.800464f
C90 VN.n47 B 0.394143f
C91 VN.n48 B 0.047648f
C92 VN.n49 B 0.242498f
C93 VN.n50 B 0.025566f
C94 VN.n51 B 0.025566f
C95 VN.n52 B 0.026306f
C96 VN.n53 B 0.050356f
C97 VN.n54 B 0.035886f
C98 VN.n55 B 0.025566f
C99 VN.n56 B 0.025566f
C100 VN.n57 B 0.025566f
C101 VN.n58 B 0.050356f
C102 VN.n59 B 0.026306f
C103 VN.n60 B 0.045634f
C104 VN.n61 B 0.025566f
C105 VN.n62 B 0.025566f
C106 VN.n63 B 0.025566f
C107 VN.n64 B 0.333734f
C108 VN.n65 B 0.047648f
C109 VN.n66 B 0.045634f
C110 VN.n67 B 0.025566f
C111 VN.n68 B 0.025566f
C112 VN.n69 B 0.025566f
C113 VN.n70 B 0.050356f
C114 VN.n71 B 0.035886f
C115 VN.n72 B 0.392303f
C116 VN.n73 B 1.29984f
C117 VDD1.t8 B 1.11002f
C118 VDD1.t5 B 0.106015f
C119 VDD1.t0 B 0.106015f
C120 VDD1.n0 B 0.862094f
C121 VDD1.n1 B 0.954269f
C122 VDD1.t9 B 1.11002f
C123 VDD1.t3 B 0.106015f
C124 VDD1.t7 B 0.106015f
C125 VDD1.n2 B 0.862091f
C126 VDD1.n3 B 0.945531f
C127 VDD1.t2 B 0.106015f
C128 VDD1.t4 B 0.106015f
C129 VDD1.n4 B 0.876098f
C130 VDD1.n5 B 2.70318f
C131 VDD1.t1 B 0.106015f
C132 VDD1.t6 B 0.106015f
C133 VDD1.n6 B 0.86209f
C134 VDD1.n7 B 2.75945f
C135 VTAIL.t5 B 0.115335f
C136 VTAIL.t6 B 0.115335f
C137 VTAIL.n0 B 0.866454f
C138 VTAIL.n1 B 0.597632f
C139 VTAIL.t15 B 1.10683f
C140 VTAIL.n2 B 0.722586f
C141 VTAIL.t12 B 0.115335f
C142 VTAIL.t17 B 0.115335f
C143 VTAIL.n3 B 0.866454f
C144 VTAIL.n4 B 0.716391f
C145 VTAIL.t10 B 0.115335f
C146 VTAIL.t16 B 0.115335f
C147 VTAIL.n5 B 0.866454f
C148 VTAIL.n6 B 1.74756f
C149 VTAIL.t2 B 0.115335f
C150 VTAIL.t8 B 0.115335f
C151 VTAIL.n7 B 0.866458f
C152 VTAIL.n8 B 1.74756f
C153 VTAIL.t4 B 0.115335f
C154 VTAIL.t9 B 0.115335f
C155 VTAIL.n9 B 0.866458f
C156 VTAIL.n10 B 0.716386f
C157 VTAIL.t7 B 1.10684f
C158 VTAIL.n11 B 0.722579f
C159 VTAIL.t13 B 0.115335f
C160 VTAIL.t14 B 0.115335f
C161 VTAIL.n12 B 0.866458f
C162 VTAIL.n13 B 0.648407f
C163 VTAIL.t19 B 0.115335f
C164 VTAIL.t18 B 0.115335f
C165 VTAIL.n14 B 0.866458f
C166 VTAIL.n15 B 0.716386f
C167 VTAIL.t11 B 1.10683f
C168 VTAIL.n16 B 1.5965f
C169 VTAIL.t1 B 1.10683f
C170 VTAIL.n17 B 1.5965f
C171 VTAIL.t3 B 0.115335f
C172 VTAIL.t0 B 0.115335f
C173 VTAIL.n18 B 0.866454f
C174 VTAIL.n19 B 0.541938f
C175 VP.n0 B 0.034567f
C176 VP.t5 B 0.820913f
C177 VP.n1 B 0.026978f
C178 VP.n2 B 0.026219f
C179 VP.t7 B 0.820913f
C180 VP.n3 B 0.048865f
C181 VP.n4 B 0.026219f
C182 VP.n5 B 0.036803f
C183 VP.n6 B 0.026219f
C184 VP.n7 B 0.0468f
C185 VP.n8 B 0.026219f
C186 VP.t6 B 0.820913f
C187 VP.n9 B 0.0468f
C188 VP.n10 B 0.026219f
C189 VP.t0 B 0.820913f
C190 VP.n11 B 0.402325f
C191 VP.n12 B 0.034567f
C192 VP.t3 B 0.820913f
C193 VP.n13 B 0.026978f
C194 VP.n14 B 0.026219f
C195 VP.t8 B 0.820913f
C196 VP.n15 B 0.048865f
C197 VP.n16 B 0.026219f
C198 VP.n17 B 0.036803f
C199 VP.n18 B 0.026219f
C200 VP.n19 B 0.0468f
C201 VP.t1 B 1.01564f
C202 VP.n20 B 0.371923f
C203 VP.t4 B 0.820913f
C204 VP.n21 B 0.404212f
C205 VP.n22 B 0.048865f
C206 VP.n23 B 0.248693f
C207 VP.n24 B 0.026219f
C208 VP.n25 B 0.026219f
C209 VP.n26 B 0.026978f
C210 VP.n27 B 0.051642f
C211 VP.t9 B 0.820913f
C212 VP.n28 B 0.31752f
C213 VP.n29 B 0.036803f
C214 VP.n30 B 0.026219f
C215 VP.n31 B 0.026219f
C216 VP.n32 B 0.026219f
C217 VP.n33 B 0.051642f
C218 VP.n34 B 0.026978f
C219 VP.n35 B 0.0468f
C220 VP.n36 B 0.026219f
C221 VP.n37 B 0.026219f
C222 VP.n38 B 0.026219f
C223 VP.n39 B 0.34226f
C224 VP.n40 B 0.048865f
C225 VP.n41 B 0.0468f
C226 VP.n42 B 0.026219f
C227 VP.n43 B 0.026219f
C228 VP.n44 B 0.026219f
C229 VP.n45 B 0.051642f
C230 VP.n46 B 0.036803f
C231 VP.n47 B 0.402325f
C232 VP.n48 B 1.31881f
C233 VP.n49 B 1.33894f
C234 VP.n50 B 0.034567f
C235 VP.n51 B 0.036803f
C236 VP.n52 B 0.051642f
C237 VP.n53 B 0.026978f
C238 VP.n54 B 0.026219f
C239 VP.n55 B 0.026219f
C240 VP.n56 B 0.026219f
C241 VP.n57 B 0.048865f
C242 VP.n58 B 0.34226f
C243 VP.n59 B 0.048865f
C244 VP.n60 B 0.026219f
C245 VP.n61 B 0.026219f
C246 VP.n62 B 0.026219f
C247 VP.n63 B 0.026978f
C248 VP.n64 B 0.051642f
C249 VP.t2 B 0.820913f
C250 VP.n65 B 0.31752f
C251 VP.n66 B 0.036803f
C252 VP.n67 B 0.026219f
C253 VP.n68 B 0.026219f
C254 VP.n69 B 0.026219f
C255 VP.n70 B 0.051642f
C256 VP.n71 B 0.026978f
C257 VP.n72 B 0.0468f
C258 VP.n73 B 0.026219f
C259 VP.n74 B 0.026219f
C260 VP.n75 B 0.026219f
C261 VP.n76 B 0.34226f
C262 VP.n77 B 0.048865f
C263 VP.n78 B 0.0468f
C264 VP.n79 B 0.026219f
C265 VP.n80 B 0.026219f
C266 VP.n81 B 0.026219f
C267 VP.n82 B 0.051642f
C268 VP.n83 B 0.036803f
C269 VP.n84 B 0.402325f
C270 VP.n85 B 0.039731f
.ends

