* NGSPICE file created from diff_pair_sample_0885.ext - technology: sky130A

.subckt diff_pair_sample_0885 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=3.07065 ps=18.94 w=18.61 l=0.96
X1 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=0.96
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=0.96
X3 VTAIL.t9 VP.t1 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=3.07065 ps=18.94 w=18.61 l=0.96
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=0.96
X5 VDD1.t5 VP.t2 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=0.96
X6 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=0.96
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=0 ps=0 w=18.61 l=0.96
X8 VTAIL.t4 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=3.07065 ps=18.94 w=18.61 l=0.96
X9 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=3.07065 ps=18.94 w=18.61 l=0.96
X10 VDD1.t4 VP.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=0.96
X11 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=0.96
X12 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=0.96
X13 VDD1.t2 VP.t4 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=0.96
X14 VDD1.t1 VP.t5 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.07065 pd=18.94 as=7.2579 ps=38 w=18.61 l=0.96
X15 VDD2.t0 VN.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2579 pd=38 as=3.07065 ps=18.94 w=18.61 l=0.96
R0 VP.n5 VP.t3 527.299
R1 VP.n12 VP.t2 508.36
R2 VP.n19 VP.t4 508.36
R3 VP.n9 VP.t5 508.36
R4 VP.n1 VP.t1 467.19
R5 VP.n4 VP.t0 467.19
R6 VP.n20 VP.n19 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n8 VP.n3 161.3
R9 VP.n10 VP.n9 161.3
R10 VP.n18 VP.n0 161.3
R11 VP.n17 VP.n16 161.3
R12 VP.n15 VP.n14 161.3
R13 VP.n13 VP.n2 161.3
R14 VP.n12 VP.n11 161.3
R15 VP.n14 VP.n13 50.6917
R16 VP.n18 VP.n17 50.6917
R17 VP.n8 VP.n7 50.6917
R18 VP.n11 VP.n10 47.2997
R19 VP.n6 VP.n5 43.2502
R20 VP.n5 VP.n4 42.2819
R21 VP.n14 VP.n1 12.234
R22 VP.n17 VP.n1 12.234
R23 VP.n7 VP.n4 12.234
R24 VP.n13 VP.n12 8.76414
R25 VP.n19 VP.n18 8.76414
R26 VP.n9 VP.n8 8.76414
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VDD1 VDD1.t4 62.7841
R36 VDD1.n1 VDD1.t5 62.6705
R37 VDD1.n1 VDD1.n0 61.0504
R38 VDD1.n3 VDD1.n2 60.8278
R39 VDD1.n3 VDD1.n1 44.5117
R40 VDD1.n2 VDD1.t0 1.06444
R41 VDD1.n2 VDD1.t1 1.06444
R42 VDD1.n0 VDD1.t3 1.06444
R43 VDD1.n0 VDD1.t2 1.06444
R44 VDD1 VDD1.n3 0.220328
R45 VTAIL.n7 VTAIL.t3 45.2131
R46 VTAIL.n11 VTAIL.t1 45.213
R47 VTAIL.n2 VTAIL.t6 45.213
R48 VTAIL.n10 VTAIL.t5 45.213
R49 VTAIL.n9 VTAIL.n8 44.1492
R50 VTAIL.n6 VTAIL.n5 44.1492
R51 VTAIL.n1 VTAIL.n0 44.149
R52 VTAIL.n4 VTAIL.n3 44.149
R53 VTAIL.n6 VTAIL.n4 30.6341
R54 VTAIL.n11 VTAIL.n10 29.5221
R55 VTAIL.n7 VTAIL.n6 1.11257
R56 VTAIL.n10 VTAIL.n9 1.11257
R57 VTAIL.n4 VTAIL.n2 1.11257
R58 VTAIL.n0 VTAIL.t2 1.06444
R59 VTAIL.n0 VTAIL.t0 1.06444
R60 VTAIL.n3 VTAIL.t8 1.06444
R61 VTAIL.n3 VTAIL.t9 1.06444
R62 VTAIL.n8 VTAIL.t7 1.06444
R63 VTAIL.n8 VTAIL.t10 1.06444
R64 VTAIL.n5 VTAIL.t11 1.06444
R65 VTAIL.n5 VTAIL.t4 1.06444
R66 VTAIL.n9 VTAIL.n7 1.02636
R67 VTAIL.n2 VTAIL.n1 1.02636
R68 VTAIL VTAIL.n11 0.776362
R69 VTAIL VTAIL.n1 0.336707
R70 B.n115 B.t17 669.835
R71 B.n113 B.t13 669.835
R72 B.n488 B.t6 669.835
R73 B.n485 B.t10 669.835
R74 B.n855 B.n854 585
R75 B.n375 B.n111 585
R76 B.n374 B.n373 585
R77 B.n372 B.n371 585
R78 B.n370 B.n369 585
R79 B.n368 B.n367 585
R80 B.n366 B.n365 585
R81 B.n364 B.n363 585
R82 B.n362 B.n361 585
R83 B.n360 B.n359 585
R84 B.n358 B.n357 585
R85 B.n356 B.n355 585
R86 B.n354 B.n353 585
R87 B.n352 B.n351 585
R88 B.n350 B.n349 585
R89 B.n348 B.n347 585
R90 B.n346 B.n345 585
R91 B.n344 B.n343 585
R92 B.n342 B.n341 585
R93 B.n340 B.n339 585
R94 B.n338 B.n337 585
R95 B.n336 B.n335 585
R96 B.n334 B.n333 585
R97 B.n332 B.n331 585
R98 B.n330 B.n329 585
R99 B.n328 B.n327 585
R100 B.n326 B.n325 585
R101 B.n324 B.n323 585
R102 B.n322 B.n321 585
R103 B.n320 B.n319 585
R104 B.n318 B.n317 585
R105 B.n316 B.n315 585
R106 B.n314 B.n313 585
R107 B.n312 B.n311 585
R108 B.n310 B.n309 585
R109 B.n308 B.n307 585
R110 B.n306 B.n305 585
R111 B.n304 B.n303 585
R112 B.n302 B.n301 585
R113 B.n300 B.n299 585
R114 B.n298 B.n297 585
R115 B.n296 B.n295 585
R116 B.n294 B.n293 585
R117 B.n292 B.n291 585
R118 B.n290 B.n289 585
R119 B.n288 B.n287 585
R120 B.n286 B.n285 585
R121 B.n284 B.n283 585
R122 B.n282 B.n281 585
R123 B.n280 B.n279 585
R124 B.n278 B.n277 585
R125 B.n276 B.n275 585
R126 B.n274 B.n273 585
R127 B.n272 B.n271 585
R128 B.n270 B.n269 585
R129 B.n268 B.n267 585
R130 B.n266 B.n265 585
R131 B.n264 B.n263 585
R132 B.n262 B.n261 585
R133 B.n260 B.n259 585
R134 B.n258 B.n257 585
R135 B.n255 B.n254 585
R136 B.n253 B.n252 585
R137 B.n251 B.n250 585
R138 B.n249 B.n248 585
R139 B.n247 B.n246 585
R140 B.n245 B.n244 585
R141 B.n243 B.n242 585
R142 B.n241 B.n240 585
R143 B.n239 B.n238 585
R144 B.n237 B.n236 585
R145 B.n234 B.n233 585
R146 B.n232 B.n231 585
R147 B.n230 B.n229 585
R148 B.n228 B.n227 585
R149 B.n226 B.n225 585
R150 B.n224 B.n223 585
R151 B.n222 B.n221 585
R152 B.n220 B.n219 585
R153 B.n218 B.n217 585
R154 B.n216 B.n215 585
R155 B.n214 B.n213 585
R156 B.n212 B.n211 585
R157 B.n210 B.n209 585
R158 B.n208 B.n207 585
R159 B.n206 B.n205 585
R160 B.n204 B.n203 585
R161 B.n202 B.n201 585
R162 B.n200 B.n199 585
R163 B.n198 B.n197 585
R164 B.n196 B.n195 585
R165 B.n194 B.n193 585
R166 B.n192 B.n191 585
R167 B.n190 B.n189 585
R168 B.n188 B.n187 585
R169 B.n186 B.n185 585
R170 B.n184 B.n183 585
R171 B.n182 B.n181 585
R172 B.n180 B.n179 585
R173 B.n178 B.n177 585
R174 B.n176 B.n175 585
R175 B.n174 B.n173 585
R176 B.n172 B.n171 585
R177 B.n170 B.n169 585
R178 B.n168 B.n167 585
R179 B.n166 B.n165 585
R180 B.n164 B.n163 585
R181 B.n162 B.n161 585
R182 B.n160 B.n159 585
R183 B.n158 B.n157 585
R184 B.n156 B.n155 585
R185 B.n154 B.n153 585
R186 B.n152 B.n151 585
R187 B.n150 B.n149 585
R188 B.n148 B.n147 585
R189 B.n146 B.n145 585
R190 B.n144 B.n143 585
R191 B.n142 B.n141 585
R192 B.n140 B.n139 585
R193 B.n138 B.n137 585
R194 B.n136 B.n135 585
R195 B.n134 B.n133 585
R196 B.n132 B.n131 585
R197 B.n130 B.n129 585
R198 B.n128 B.n127 585
R199 B.n126 B.n125 585
R200 B.n124 B.n123 585
R201 B.n122 B.n121 585
R202 B.n120 B.n119 585
R203 B.n118 B.n117 585
R204 B.n46 B.n45 585
R205 B.n860 B.n859 585
R206 B.n853 B.n112 585
R207 B.n112 B.n43 585
R208 B.n852 B.n42 585
R209 B.n864 B.n42 585
R210 B.n851 B.n41 585
R211 B.n865 B.n41 585
R212 B.n850 B.n40 585
R213 B.n866 B.n40 585
R214 B.n849 B.n848 585
R215 B.n848 B.n36 585
R216 B.n847 B.n35 585
R217 B.n872 B.n35 585
R218 B.n846 B.n34 585
R219 B.n873 B.n34 585
R220 B.n845 B.n33 585
R221 B.n874 B.n33 585
R222 B.n844 B.n843 585
R223 B.n843 B.n29 585
R224 B.n842 B.n28 585
R225 B.n880 B.n28 585
R226 B.n841 B.n27 585
R227 B.n881 B.n27 585
R228 B.n840 B.n26 585
R229 B.n882 B.n26 585
R230 B.n839 B.n838 585
R231 B.n838 B.n25 585
R232 B.n837 B.n21 585
R233 B.n888 B.n21 585
R234 B.n836 B.n20 585
R235 B.n889 B.n20 585
R236 B.n835 B.n19 585
R237 B.n890 B.n19 585
R238 B.n834 B.n833 585
R239 B.n833 B.n18 585
R240 B.n832 B.n14 585
R241 B.n896 B.n14 585
R242 B.n831 B.n13 585
R243 B.n897 B.n13 585
R244 B.n830 B.n12 585
R245 B.n898 B.n12 585
R246 B.n829 B.n828 585
R247 B.n828 B.t2 585
R248 B.n827 B.n826 585
R249 B.n827 B.n8 585
R250 B.n825 B.n7 585
R251 B.n905 B.n7 585
R252 B.n824 B.n6 585
R253 B.n906 B.n6 585
R254 B.n823 B.n5 585
R255 B.n907 B.n5 585
R256 B.n822 B.n821 585
R257 B.n821 B.n4 585
R258 B.n820 B.n376 585
R259 B.n820 B.n819 585
R260 B.n810 B.n377 585
R261 B.t3 B.n377 585
R262 B.n812 B.n811 585
R263 B.n813 B.n812 585
R264 B.n809 B.n382 585
R265 B.n382 B.n381 585
R266 B.n808 B.n807 585
R267 B.n807 B.n806 585
R268 B.n384 B.n383 585
R269 B.n799 B.n384 585
R270 B.n798 B.n797 585
R271 B.n800 B.n798 585
R272 B.n796 B.n389 585
R273 B.n389 B.n388 585
R274 B.n795 B.n794 585
R275 B.n794 B.n793 585
R276 B.n391 B.n390 585
R277 B.n786 B.n391 585
R278 B.n785 B.n784 585
R279 B.n787 B.n785 585
R280 B.n783 B.n396 585
R281 B.n396 B.n395 585
R282 B.n782 B.n781 585
R283 B.n781 B.n780 585
R284 B.n398 B.n397 585
R285 B.n399 B.n398 585
R286 B.n773 B.n772 585
R287 B.n774 B.n773 585
R288 B.n771 B.n404 585
R289 B.n404 B.n403 585
R290 B.n770 B.n769 585
R291 B.n769 B.n768 585
R292 B.n406 B.n405 585
R293 B.n407 B.n406 585
R294 B.n761 B.n760 585
R295 B.n762 B.n761 585
R296 B.n759 B.n412 585
R297 B.n412 B.n411 585
R298 B.n758 B.n757 585
R299 B.n757 B.n756 585
R300 B.n414 B.n413 585
R301 B.n415 B.n414 585
R302 B.n752 B.n751 585
R303 B.n418 B.n417 585
R304 B.n748 B.n747 585
R305 B.n749 B.n748 585
R306 B.n746 B.n484 585
R307 B.n745 B.n744 585
R308 B.n743 B.n742 585
R309 B.n741 B.n740 585
R310 B.n739 B.n738 585
R311 B.n737 B.n736 585
R312 B.n735 B.n734 585
R313 B.n733 B.n732 585
R314 B.n731 B.n730 585
R315 B.n729 B.n728 585
R316 B.n727 B.n726 585
R317 B.n725 B.n724 585
R318 B.n723 B.n722 585
R319 B.n721 B.n720 585
R320 B.n719 B.n718 585
R321 B.n717 B.n716 585
R322 B.n715 B.n714 585
R323 B.n713 B.n712 585
R324 B.n711 B.n710 585
R325 B.n709 B.n708 585
R326 B.n707 B.n706 585
R327 B.n705 B.n704 585
R328 B.n703 B.n702 585
R329 B.n701 B.n700 585
R330 B.n699 B.n698 585
R331 B.n697 B.n696 585
R332 B.n695 B.n694 585
R333 B.n693 B.n692 585
R334 B.n691 B.n690 585
R335 B.n689 B.n688 585
R336 B.n687 B.n686 585
R337 B.n685 B.n684 585
R338 B.n683 B.n682 585
R339 B.n681 B.n680 585
R340 B.n679 B.n678 585
R341 B.n677 B.n676 585
R342 B.n675 B.n674 585
R343 B.n673 B.n672 585
R344 B.n671 B.n670 585
R345 B.n669 B.n668 585
R346 B.n667 B.n666 585
R347 B.n665 B.n664 585
R348 B.n663 B.n662 585
R349 B.n661 B.n660 585
R350 B.n659 B.n658 585
R351 B.n657 B.n656 585
R352 B.n655 B.n654 585
R353 B.n653 B.n652 585
R354 B.n651 B.n650 585
R355 B.n649 B.n648 585
R356 B.n647 B.n646 585
R357 B.n645 B.n644 585
R358 B.n643 B.n642 585
R359 B.n641 B.n640 585
R360 B.n639 B.n638 585
R361 B.n637 B.n636 585
R362 B.n635 B.n634 585
R363 B.n633 B.n632 585
R364 B.n631 B.n630 585
R365 B.n629 B.n628 585
R366 B.n627 B.n626 585
R367 B.n625 B.n624 585
R368 B.n623 B.n622 585
R369 B.n621 B.n620 585
R370 B.n619 B.n618 585
R371 B.n617 B.n616 585
R372 B.n615 B.n614 585
R373 B.n613 B.n612 585
R374 B.n611 B.n610 585
R375 B.n609 B.n608 585
R376 B.n607 B.n606 585
R377 B.n605 B.n604 585
R378 B.n603 B.n602 585
R379 B.n601 B.n600 585
R380 B.n599 B.n598 585
R381 B.n597 B.n596 585
R382 B.n595 B.n594 585
R383 B.n593 B.n592 585
R384 B.n591 B.n590 585
R385 B.n589 B.n588 585
R386 B.n587 B.n586 585
R387 B.n585 B.n584 585
R388 B.n583 B.n582 585
R389 B.n581 B.n580 585
R390 B.n579 B.n578 585
R391 B.n577 B.n576 585
R392 B.n575 B.n574 585
R393 B.n573 B.n572 585
R394 B.n571 B.n570 585
R395 B.n569 B.n568 585
R396 B.n567 B.n566 585
R397 B.n565 B.n564 585
R398 B.n563 B.n562 585
R399 B.n561 B.n560 585
R400 B.n559 B.n558 585
R401 B.n557 B.n556 585
R402 B.n555 B.n554 585
R403 B.n553 B.n552 585
R404 B.n551 B.n550 585
R405 B.n549 B.n548 585
R406 B.n547 B.n546 585
R407 B.n545 B.n544 585
R408 B.n543 B.n542 585
R409 B.n541 B.n540 585
R410 B.n539 B.n538 585
R411 B.n537 B.n536 585
R412 B.n535 B.n534 585
R413 B.n533 B.n532 585
R414 B.n531 B.n530 585
R415 B.n529 B.n528 585
R416 B.n527 B.n526 585
R417 B.n525 B.n524 585
R418 B.n523 B.n522 585
R419 B.n521 B.n520 585
R420 B.n519 B.n518 585
R421 B.n517 B.n516 585
R422 B.n515 B.n514 585
R423 B.n513 B.n512 585
R424 B.n511 B.n510 585
R425 B.n509 B.n508 585
R426 B.n507 B.n506 585
R427 B.n505 B.n504 585
R428 B.n503 B.n502 585
R429 B.n501 B.n500 585
R430 B.n499 B.n498 585
R431 B.n497 B.n496 585
R432 B.n495 B.n494 585
R433 B.n493 B.n492 585
R434 B.n491 B.n483 585
R435 B.n749 B.n483 585
R436 B.n753 B.n416 585
R437 B.n416 B.n415 585
R438 B.n755 B.n754 585
R439 B.n756 B.n755 585
R440 B.n410 B.n409 585
R441 B.n411 B.n410 585
R442 B.n764 B.n763 585
R443 B.n763 B.n762 585
R444 B.n765 B.n408 585
R445 B.n408 B.n407 585
R446 B.n767 B.n766 585
R447 B.n768 B.n767 585
R448 B.n402 B.n401 585
R449 B.n403 B.n402 585
R450 B.n776 B.n775 585
R451 B.n775 B.n774 585
R452 B.n777 B.n400 585
R453 B.n400 B.n399 585
R454 B.n779 B.n778 585
R455 B.n780 B.n779 585
R456 B.n394 B.n393 585
R457 B.n395 B.n394 585
R458 B.n789 B.n788 585
R459 B.n788 B.n787 585
R460 B.n790 B.n392 585
R461 B.n786 B.n392 585
R462 B.n792 B.n791 585
R463 B.n793 B.n792 585
R464 B.n387 B.n386 585
R465 B.n388 B.n387 585
R466 B.n802 B.n801 585
R467 B.n801 B.n800 585
R468 B.n803 B.n385 585
R469 B.n799 B.n385 585
R470 B.n805 B.n804 585
R471 B.n806 B.n805 585
R472 B.n380 B.n379 585
R473 B.n381 B.n380 585
R474 B.n815 B.n814 585
R475 B.n814 B.n813 585
R476 B.n816 B.n378 585
R477 B.n378 B.t3 585
R478 B.n818 B.n817 585
R479 B.n819 B.n818 585
R480 B.n3 B.n0 585
R481 B.n4 B.n3 585
R482 B.n904 B.n1 585
R483 B.n905 B.n904 585
R484 B.n903 B.n902 585
R485 B.n903 B.n8 585
R486 B.n901 B.n9 585
R487 B.t2 B.n9 585
R488 B.n900 B.n899 585
R489 B.n899 B.n898 585
R490 B.n11 B.n10 585
R491 B.n897 B.n11 585
R492 B.n895 B.n894 585
R493 B.n896 B.n895 585
R494 B.n893 B.n15 585
R495 B.n18 B.n15 585
R496 B.n892 B.n891 585
R497 B.n891 B.n890 585
R498 B.n17 B.n16 585
R499 B.n889 B.n17 585
R500 B.n887 B.n886 585
R501 B.n888 B.n887 585
R502 B.n885 B.n22 585
R503 B.n25 B.n22 585
R504 B.n884 B.n883 585
R505 B.n883 B.n882 585
R506 B.n24 B.n23 585
R507 B.n881 B.n24 585
R508 B.n879 B.n878 585
R509 B.n880 B.n879 585
R510 B.n877 B.n30 585
R511 B.n30 B.n29 585
R512 B.n876 B.n875 585
R513 B.n875 B.n874 585
R514 B.n32 B.n31 585
R515 B.n873 B.n32 585
R516 B.n871 B.n870 585
R517 B.n872 B.n871 585
R518 B.n869 B.n37 585
R519 B.n37 B.n36 585
R520 B.n868 B.n867 585
R521 B.n867 B.n866 585
R522 B.n39 B.n38 585
R523 B.n865 B.n39 585
R524 B.n863 B.n862 585
R525 B.n864 B.n863 585
R526 B.n861 B.n44 585
R527 B.n44 B.n43 585
R528 B.n908 B.n907 585
R529 B.n906 B.n2 585
R530 B.n859 B.n44 439.647
R531 B.n855 B.n112 439.647
R532 B.n483 B.n414 439.647
R533 B.n751 B.n416 439.647
R534 B.n857 B.n856 256.663
R535 B.n857 B.n110 256.663
R536 B.n857 B.n109 256.663
R537 B.n857 B.n108 256.663
R538 B.n857 B.n107 256.663
R539 B.n857 B.n106 256.663
R540 B.n857 B.n105 256.663
R541 B.n857 B.n104 256.663
R542 B.n857 B.n103 256.663
R543 B.n857 B.n102 256.663
R544 B.n857 B.n101 256.663
R545 B.n857 B.n100 256.663
R546 B.n857 B.n99 256.663
R547 B.n857 B.n98 256.663
R548 B.n857 B.n97 256.663
R549 B.n857 B.n96 256.663
R550 B.n857 B.n95 256.663
R551 B.n857 B.n94 256.663
R552 B.n857 B.n93 256.663
R553 B.n857 B.n92 256.663
R554 B.n857 B.n91 256.663
R555 B.n857 B.n90 256.663
R556 B.n857 B.n89 256.663
R557 B.n857 B.n88 256.663
R558 B.n857 B.n87 256.663
R559 B.n857 B.n86 256.663
R560 B.n857 B.n85 256.663
R561 B.n857 B.n84 256.663
R562 B.n857 B.n83 256.663
R563 B.n857 B.n82 256.663
R564 B.n857 B.n81 256.663
R565 B.n857 B.n80 256.663
R566 B.n857 B.n79 256.663
R567 B.n857 B.n78 256.663
R568 B.n857 B.n77 256.663
R569 B.n857 B.n76 256.663
R570 B.n857 B.n75 256.663
R571 B.n857 B.n74 256.663
R572 B.n857 B.n73 256.663
R573 B.n857 B.n72 256.663
R574 B.n857 B.n71 256.663
R575 B.n857 B.n70 256.663
R576 B.n857 B.n69 256.663
R577 B.n857 B.n68 256.663
R578 B.n857 B.n67 256.663
R579 B.n857 B.n66 256.663
R580 B.n857 B.n65 256.663
R581 B.n857 B.n64 256.663
R582 B.n857 B.n63 256.663
R583 B.n857 B.n62 256.663
R584 B.n857 B.n61 256.663
R585 B.n857 B.n60 256.663
R586 B.n857 B.n59 256.663
R587 B.n857 B.n58 256.663
R588 B.n857 B.n57 256.663
R589 B.n857 B.n56 256.663
R590 B.n857 B.n55 256.663
R591 B.n857 B.n54 256.663
R592 B.n857 B.n53 256.663
R593 B.n857 B.n52 256.663
R594 B.n857 B.n51 256.663
R595 B.n857 B.n50 256.663
R596 B.n857 B.n49 256.663
R597 B.n857 B.n48 256.663
R598 B.n857 B.n47 256.663
R599 B.n858 B.n857 256.663
R600 B.n750 B.n749 256.663
R601 B.n749 B.n419 256.663
R602 B.n749 B.n420 256.663
R603 B.n749 B.n421 256.663
R604 B.n749 B.n422 256.663
R605 B.n749 B.n423 256.663
R606 B.n749 B.n424 256.663
R607 B.n749 B.n425 256.663
R608 B.n749 B.n426 256.663
R609 B.n749 B.n427 256.663
R610 B.n749 B.n428 256.663
R611 B.n749 B.n429 256.663
R612 B.n749 B.n430 256.663
R613 B.n749 B.n431 256.663
R614 B.n749 B.n432 256.663
R615 B.n749 B.n433 256.663
R616 B.n749 B.n434 256.663
R617 B.n749 B.n435 256.663
R618 B.n749 B.n436 256.663
R619 B.n749 B.n437 256.663
R620 B.n749 B.n438 256.663
R621 B.n749 B.n439 256.663
R622 B.n749 B.n440 256.663
R623 B.n749 B.n441 256.663
R624 B.n749 B.n442 256.663
R625 B.n749 B.n443 256.663
R626 B.n749 B.n444 256.663
R627 B.n749 B.n445 256.663
R628 B.n749 B.n446 256.663
R629 B.n749 B.n447 256.663
R630 B.n749 B.n448 256.663
R631 B.n749 B.n449 256.663
R632 B.n749 B.n450 256.663
R633 B.n749 B.n451 256.663
R634 B.n749 B.n452 256.663
R635 B.n749 B.n453 256.663
R636 B.n749 B.n454 256.663
R637 B.n749 B.n455 256.663
R638 B.n749 B.n456 256.663
R639 B.n749 B.n457 256.663
R640 B.n749 B.n458 256.663
R641 B.n749 B.n459 256.663
R642 B.n749 B.n460 256.663
R643 B.n749 B.n461 256.663
R644 B.n749 B.n462 256.663
R645 B.n749 B.n463 256.663
R646 B.n749 B.n464 256.663
R647 B.n749 B.n465 256.663
R648 B.n749 B.n466 256.663
R649 B.n749 B.n467 256.663
R650 B.n749 B.n468 256.663
R651 B.n749 B.n469 256.663
R652 B.n749 B.n470 256.663
R653 B.n749 B.n471 256.663
R654 B.n749 B.n472 256.663
R655 B.n749 B.n473 256.663
R656 B.n749 B.n474 256.663
R657 B.n749 B.n475 256.663
R658 B.n749 B.n476 256.663
R659 B.n749 B.n477 256.663
R660 B.n749 B.n478 256.663
R661 B.n749 B.n479 256.663
R662 B.n749 B.n480 256.663
R663 B.n749 B.n481 256.663
R664 B.n749 B.n482 256.663
R665 B.n910 B.n909 256.663
R666 B.n117 B.n46 163.367
R667 B.n121 B.n120 163.367
R668 B.n125 B.n124 163.367
R669 B.n129 B.n128 163.367
R670 B.n133 B.n132 163.367
R671 B.n137 B.n136 163.367
R672 B.n141 B.n140 163.367
R673 B.n145 B.n144 163.367
R674 B.n149 B.n148 163.367
R675 B.n153 B.n152 163.367
R676 B.n157 B.n156 163.367
R677 B.n161 B.n160 163.367
R678 B.n165 B.n164 163.367
R679 B.n169 B.n168 163.367
R680 B.n173 B.n172 163.367
R681 B.n177 B.n176 163.367
R682 B.n181 B.n180 163.367
R683 B.n185 B.n184 163.367
R684 B.n189 B.n188 163.367
R685 B.n193 B.n192 163.367
R686 B.n197 B.n196 163.367
R687 B.n201 B.n200 163.367
R688 B.n205 B.n204 163.367
R689 B.n209 B.n208 163.367
R690 B.n213 B.n212 163.367
R691 B.n217 B.n216 163.367
R692 B.n221 B.n220 163.367
R693 B.n225 B.n224 163.367
R694 B.n229 B.n228 163.367
R695 B.n233 B.n232 163.367
R696 B.n238 B.n237 163.367
R697 B.n242 B.n241 163.367
R698 B.n246 B.n245 163.367
R699 B.n250 B.n249 163.367
R700 B.n254 B.n253 163.367
R701 B.n259 B.n258 163.367
R702 B.n263 B.n262 163.367
R703 B.n267 B.n266 163.367
R704 B.n271 B.n270 163.367
R705 B.n275 B.n274 163.367
R706 B.n279 B.n278 163.367
R707 B.n283 B.n282 163.367
R708 B.n287 B.n286 163.367
R709 B.n291 B.n290 163.367
R710 B.n295 B.n294 163.367
R711 B.n299 B.n298 163.367
R712 B.n303 B.n302 163.367
R713 B.n307 B.n306 163.367
R714 B.n311 B.n310 163.367
R715 B.n315 B.n314 163.367
R716 B.n319 B.n318 163.367
R717 B.n323 B.n322 163.367
R718 B.n327 B.n326 163.367
R719 B.n331 B.n330 163.367
R720 B.n335 B.n334 163.367
R721 B.n339 B.n338 163.367
R722 B.n343 B.n342 163.367
R723 B.n347 B.n346 163.367
R724 B.n351 B.n350 163.367
R725 B.n355 B.n354 163.367
R726 B.n359 B.n358 163.367
R727 B.n363 B.n362 163.367
R728 B.n367 B.n366 163.367
R729 B.n371 B.n370 163.367
R730 B.n373 B.n111 163.367
R731 B.n757 B.n414 163.367
R732 B.n757 B.n412 163.367
R733 B.n761 B.n412 163.367
R734 B.n761 B.n406 163.367
R735 B.n769 B.n406 163.367
R736 B.n769 B.n404 163.367
R737 B.n773 B.n404 163.367
R738 B.n773 B.n398 163.367
R739 B.n781 B.n398 163.367
R740 B.n781 B.n396 163.367
R741 B.n785 B.n396 163.367
R742 B.n785 B.n391 163.367
R743 B.n794 B.n391 163.367
R744 B.n794 B.n389 163.367
R745 B.n798 B.n389 163.367
R746 B.n798 B.n384 163.367
R747 B.n807 B.n384 163.367
R748 B.n807 B.n382 163.367
R749 B.n812 B.n382 163.367
R750 B.n812 B.n377 163.367
R751 B.n820 B.n377 163.367
R752 B.n821 B.n820 163.367
R753 B.n821 B.n5 163.367
R754 B.n6 B.n5 163.367
R755 B.n7 B.n6 163.367
R756 B.n827 B.n7 163.367
R757 B.n828 B.n827 163.367
R758 B.n828 B.n12 163.367
R759 B.n13 B.n12 163.367
R760 B.n14 B.n13 163.367
R761 B.n833 B.n14 163.367
R762 B.n833 B.n19 163.367
R763 B.n20 B.n19 163.367
R764 B.n21 B.n20 163.367
R765 B.n838 B.n21 163.367
R766 B.n838 B.n26 163.367
R767 B.n27 B.n26 163.367
R768 B.n28 B.n27 163.367
R769 B.n843 B.n28 163.367
R770 B.n843 B.n33 163.367
R771 B.n34 B.n33 163.367
R772 B.n35 B.n34 163.367
R773 B.n848 B.n35 163.367
R774 B.n848 B.n40 163.367
R775 B.n41 B.n40 163.367
R776 B.n42 B.n41 163.367
R777 B.n112 B.n42 163.367
R778 B.n748 B.n418 163.367
R779 B.n748 B.n484 163.367
R780 B.n744 B.n743 163.367
R781 B.n740 B.n739 163.367
R782 B.n736 B.n735 163.367
R783 B.n732 B.n731 163.367
R784 B.n728 B.n727 163.367
R785 B.n724 B.n723 163.367
R786 B.n720 B.n719 163.367
R787 B.n716 B.n715 163.367
R788 B.n712 B.n711 163.367
R789 B.n708 B.n707 163.367
R790 B.n704 B.n703 163.367
R791 B.n700 B.n699 163.367
R792 B.n696 B.n695 163.367
R793 B.n692 B.n691 163.367
R794 B.n688 B.n687 163.367
R795 B.n684 B.n683 163.367
R796 B.n680 B.n679 163.367
R797 B.n676 B.n675 163.367
R798 B.n672 B.n671 163.367
R799 B.n668 B.n667 163.367
R800 B.n664 B.n663 163.367
R801 B.n660 B.n659 163.367
R802 B.n656 B.n655 163.367
R803 B.n652 B.n651 163.367
R804 B.n648 B.n647 163.367
R805 B.n644 B.n643 163.367
R806 B.n640 B.n639 163.367
R807 B.n636 B.n635 163.367
R808 B.n632 B.n631 163.367
R809 B.n628 B.n627 163.367
R810 B.n624 B.n623 163.367
R811 B.n620 B.n619 163.367
R812 B.n616 B.n615 163.367
R813 B.n612 B.n611 163.367
R814 B.n608 B.n607 163.367
R815 B.n604 B.n603 163.367
R816 B.n600 B.n599 163.367
R817 B.n596 B.n595 163.367
R818 B.n592 B.n591 163.367
R819 B.n588 B.n587 163.367
R820 B.n584 B.n583 163.367
R821 B.n580 B.n579 163.367
R822 B.n576 B.n575 163.367
R823 B.n572 B.n571 163.367
R824 B.n568 B.n567 163.367
R825 B.n564 B.n563 163.367
R826 B.n560 B.n559 163.367
R827 B.n556 B.n555 163.367
R828 B.n552 B.n551 163.367
R829 B.n548 B.n547 163.367
R830 B.n544 B.n543 163.367
R831 B.n540 B.n539 163.367
R832 B.n536 B.n535 163.367
R833 B.n532 B.n531 163.367
R834 B.n528 B.n527 163.367
R835 B.n524 B.n523 163.367
R836 B.n520 B.n519 163.367
R837 B.n516 B.n515 163.367
R838 B.n512 B.n511 163.367
R839 B.n508 B.n507 163.367
R840 B.n504 B.n503 163.367
R841 B.n500 B.n499 163.367
R842 B.n496 B.n495 163.367
R843 B.n492 B.n483 163.367
R844 B.n755 B.n416 163.367
R845 B.n755 B.n410 163.367
R846 B.n763 B.n410 163.367
R847 B.n763 B.n408 163.367
R848 B.n767 B.n408 163.367
R849 B.n767 B.n402 163.367
R850 B.n775 B.n402 163.367
R851 B.n775 B.n400 163.367
R852 B.n779 B.n400 163.367
R853 B.n779 B.n394 163.367
R854 B.n788 B.n394 163.367
R855 B.n788 B.n392 163.367
R856 B.n792 B.n392 163.367
R857 B.n792 B.n387 163.367
R858 B.n801 B.n387 163.367
R859 B.n801 B.n385 163.367
R860 B.n805 B.n385 163.367
R861 B.n805 B.n380 163.367
R862 B.n814 B.n380 163.367
R863 B.n814 B.n378 163.367
R864 B.n818 B.n378 163.367
R865 B.n818 B.n3 163.367
R866 B.n908 B.n3 163.367
R867 B.n904 B.n2 163.367
R868 B.n904 B.n903 163.367
R869 B.n903 B.n9 163.367
R870 B.n899 B.n9 163.367
R871 B.n899 B.n11 163.367
R872 B.n895 B.n11 163.367
R873 B.n895 B.n15 163.367
R874 B.n891 B.n15 163.367
R875 B.n891 B.n17 163.367
R876 B.n887 B.n17 163.367
R877 B.n887 B.n22 163.367
R878 B.n883 B.n22 163.367
R879 B.n883 B.n24 163.367
R880 B.n879 B.n24 163.367
R881 B.n879 B.n30 163.367
R882 B.n875 B.n30 163.367
R883 B.n875 B.n32 163.367
R884 B.n871 B.n32 163.367
R885 B.n871 B.n37 163.367
R886 B.n867 B.n37 163.367
R887 B.n867 B.n39 163.367
R888 B.n863 B.n39 163.367
R889 B.n863 B.n44 163.367
R890 B.n113 B.t15 97.08
R891 B.n488 B.t9 97.08
R892 B.n115 B.t18 97.0553
R893 B.n485 B.t12 97.0553
R894 B.n114 B.t16 72.0618
R895 B.n489 B.t8 72.0618
R896 B.n116 B.t19 72.0371
R897 B.n486 B.t11 72.0371
R898 B.n859 B.n858 71.676
R899 B.n117 B.n47 71.676
R900 B.n121 B.n48 71.676
R901 B.n125 B.n49 71.676
R902 B.n129 B.n50 71.676
R903 B.n133 B.n51 71.676
R904 B.n137 B.n52 71.676
R905 B.n141 B.n53 71.676
R906 B.n145 B.n54 71.676
R907 B.n149 B.n55 71.676
R908 B.n153 B.n56 71.676
R909 B.n157 B.n57 71.676
R910 B.n161 B.n58 71.676
R911 B.n165 B.n59 71.676
R912 B.n169 B.n60 71.676
R913 B.n173 B.n61 71.676
R914 B.n177 B.n62 71.676
R915 B.n181 B.n63 71.676
R916 B.n185 B.n64 71.676
R917 B.n189 B.n65 71.676
R918 B.n193 B.n66 71.676
R919 B.n197 B.n67 71.676
R920 B.n201 B.n68 71.676
R921 B.n205 B.n69 71.676
R922 B.n209 B.n70 71.676
R923 B.n213 B.n71 71.676
R924 B.n217 B.n72 71.676
R925 B.n221 B.n73 71.676
R926 B.n225 B.n74 71.676
R927 B.n229 B.n75 71.676
R928 B.n233 B.n76 71.676
R929 B.n238 B.n77 71.676
R930 B.n242 B.n78 71.676
R931 B.n246 B.n79 71.676
R932 B.n250 B.n80 71.676
R933 B.n254 B.n81 71.676
R934 B.n259 B.n82 71.676
R935 B.n263 B.n83 71.676
R936 B.n267 B.n84 71.676
R937 B.n271 B.n85 71.676
R938 B.n275 B.n86 71.676
R939 B.n279 B.n87 71.676
R940 B.n283 B.n88 71.676
R941 B.n287 B.n89 71.676
R942 B.n291 B.n90 71.676
R943 B.n295 B.n91 71.676
R944 B.n299 B.n92 71.676
R945 B.n303 B.n93 71.676
R946 B.n307 B.n94 71.676
R947 B.n311 B.n95 71.676
R948 B.n315 B.n96 71.676
R949 B.n319 B.n97 71.676
R950 B.n323 B.n98 71.676
R951 B.n327 B.n99 71.676
R952 B.n331 B.n100 71.676
R953 B.n335 B.n101 71.676
R954 B.n339 B.n102 71.676
R955 B.n343 B.n103 71.676
R956 B.n347 B.n104 71.676
R957 B.n351 B.n105 71.676
R958 B.n355 B.n106 71.676
R959 B.n359 B.n107 71.676
R960 B.n363 B.n108 71.676
R961 B.n367 B.n109 71.676
R962 B.n371 B.n110 71.676
R963 B.n856 B.n111 71.676
R964 B.n856 B.n855 71.676
R965 B.n373 B.n110 71.676
R966 B.n370 B.n109 71.676
R967 B.n366 B.n108 71.676
R968 B.n362 B.n107 71.676
R969 B.n358 B.n106 71.676
R970 B.n354 B.n105 71.676
R971 B.n350 B.n104 71.676
R972 B.n346 B.n103 71.676
R973 B.n342 B.n102 71.676
R974 B.n338 B.n101 71.676
R975 B.n334 B.n100 71.676
R976 B.n330 B.n99 71.676
R977 B.n326 B.n98 71.676
R978 B.n322 B.n97 71.676
R979 B.n318 B.n96 71.676
R980 B.n314 B.n95 71.676
R981 B.n310 B.n94 71.676
R982 B.n306 B.n93 71.676
R983 B.n302 B.n92 71.676
R984 B.n298 B.n91 71.676
R985 B.n294 B.n90 71.676
R986 B.n290 B.n89 71.676
R987 B.n286 B.n88 71.676
R988 B.n282 B.n87 71.676
R989 B.n278 B.n86 71.676
R990 B.n274 B.n85 71.676
R991 B.n270 B.n84 71.676
R992 B.n266 B.n83 71.676
R993 B.n262 B.n82 71.676
R994 B.n258 B.n81 71.676
R995 B.n253 B.n80 71.676
R996 B.n249 B.n79 71.676
R997 B.n245 B.n78 71.676
R998 B.n241 B.n77 71.676
R999 B.n237 B.n76 71.676
R1000 B.n232 B.n75 71.676
R1001 B.n228 B.n74 71.676
R1002 B.n224 B.n73 71.676
R1003 B.n220 B.n72 71.676
R1004 B.n216 B.n71 71.676
R1005 B.n212 B.n70 71.676
R1006 B.n208 B.n69 71.676
R1007 B.n204 B.n68 71.676
R1008 B.n200 B.n67 71.676
R1009 B.n196 B.n66 71.676
R1010 B.n192 B.n65 71.676
R1011 B.n188 B.n64 71.676
R1012 B.n184 B.n63 71.676
R1013 B.n180 B.n62 71.676
R1014 B.n176 B.n61 71.676
R1015 B.n172 B.n60 71.676
R1016 B.n168 B.n59 71.676
R1017 B.n164 B.n58 71.676
R1018 B.n160 B.n57 71.676
R1019 B.n156 B.n56 71.676
R1020 B.n152 B.n55 71.676
R1021 B.n148 B.n54 71.676
R1022 B.n144 B.n53 71.676
R1023 B.n140 B.n52 71.676
R1024 B.n136 B.n51 71.676
R1025 B.n132 B.n50 71.676
R1026 B.n128 B.n49 71.676
R1027 B.n124 B.n48 71.676
R1028 B.n120 B.n47 71.676
R1029 B.n858 B.n46 71.676
R1030 B.n751 B.n750 71.676
R1031 B.n484 B.n419 71.676
R1032 B.n743 B.n420 71.676
R1033 B.n739 B.n421 71.676
R1034 B.n735 B.n422 71.676
R1035 B.n731 B.n423 71.676
R1036 B.n727 B.n424 71.676
R1037 B.n723 B.n425 71.676
R1038 B.n719 B.n426 71.676
R1039 B.n715 B.n427 71.676
R1040 B.n711 B.n428 71.676
R1041 B.n707 B.n429 71.676
R1042 B.n703 B.n430 71.676
R1043 B.n699 B.n431 71.676
R1044 B.n695 B.n432 71.676
R1045 B.n691 B.n433 71.676
R1046 B.n687 B.n434 71.676
R1047 B.n683 B.n435 71.676
R1048 B.n679 B.n436 71.676
R1049 B.n675 B.n437 71.676
R1050 B.n671 B.n438 71.676
R1051 B.n667 B.n439 71.676
R1052 B.n663 B.n440 71.676
R1053 B.n659 B.n441 71.676
R1054 B.n655 B.n442 71.676
R1055 B.n651 B.n443 71.676
R1056 B.n647 B.n444 71.676
R1057 B.n643 B.n445 71.676
R1058 B.n639 B.n446 71.676
R1059 B.n635 B.n447 71.676
R1060 B.n631 B.n448 71.676
R1061 B.n627 B.n449 71.676
R1062 B.n623 B.n450 71.676
R1063 B.n619 B.n451 71.676
R1064 B.n615 B.n452 71.676
R1065 B.n611 B.n453 71.676
R1066 B.n607 B.n454 71.676
R1067 B.n603 B.n455 71.676
R1068 B.n599 B.n456 71.676
R1069 B.n595 B.n457 71.676
R1070 B.n591 B.n458 71.676
R1071 B.n587 B.n459 71.676
R1072 B.n583 B.n460 71.676
R1073 B.n579 B.n461 71.676
R1074 B.n575 B.n462 71.676
R1075 B.n571 B.n463 71.676
R1076 B.n567 B.n464 71.676
R1077 B.n563 B.n465 71.676
R1078 B.n559 B.n466 71.676
R1079 B.n555 B.n467 71.676
R1080 B.n551 B.n468 71.676
R1081 B.n547 B.n469 71.676
R1082 B.n543 B.n470 71.676
R1083 B.n539 B.n471 71.676
R1084 B.n535 B.n472 71.676
R1085 B.n531 B.n473 71.676
R1086 B.n527 B.n474 71.676
R1087 B.n523 B.n475 71.676
R1088 B.n519 B.n476 71.676
R1089 B.n515 B.n477 71.676
R1090 B.n511 B.n478 71.676
R1091 B.n507 B.n479 71.676
R1092 B.n503 B.n480 71.676
R1093 B.n499 B.n481 71.676
R1094 B.n495 B.n482 71.676
R1095 B.n750 B.n418 71.676
R1096 B.n744 B.n419 71.676
R1097 B.n740 B.n420 71.676
R1098 B.n736 B.n421 71.676
R1099 B.n732 B.n422 71.676
R1100 B.n728 B.n423 71.676
R1101 B.n724 B.n424 71.676
R1102 B.n720 B.n425 71.676
R1103 B.n716 B.n426 71.676
R1104 B.n712 B.n427 71.676
R1105 B.n708 B.n428 71.676
R1106 B.n704 B.n429 71.676
R1107 B.n700 B.n430 71.676
R1108 B.n696 B.n431 71.676
R1109 B.n692 B.n432 71.676
R1110 B.n688 B.n433 71.676
R1111 B.n684 B.n434 71.676
R1112 B.n680 B.n435 71.676
R1113 B.n676 B.n436 71.676
R1114 B.n672 B.n437 71.676
R1115 B.n668 B.n438 71.676
R1116 B.n664 B.n439 71.676
R1117 B.n660 B.n440 71.676
R1118 B.n656 B.n441 71.676
R1119 B.n652 B.n442 71.676
R1120 B.n648 B.n443 71.676
R1121 B.n644 B.n444 71.676
R1122 B.n640 B.n445 71.676
R1123 B.n636 B.n446 71.676
R1124 B.n632 B.n447 71.676
R1125 B.n628 B.n448 71.676
R1126 B.n624 B.n449 71.676
R1127 B.n620 B.n450 71.676
R1128 B.n616 B.n451 71.676
R1129 B.n612 B.n452 71.676
R1130 B.n608 B.n453 71.676
R1131 B.n604 B.n454 71.676
R1132 B.n600 B.n455 71.676
R1133 B.n596 B.n456 71.676
R1134 B.n592 B.n457 71.676
R1135 B.n588 B.n458 71.676
R1136 B.n584 B.n459 71.676
R1137 B.n580 B.n460 71.676
R1138 B.n576 B.n461 71.676
R1139 B.n572 B.n462 71.676
R1140 B.n568 B.n463 71.676
R1141 B.n564 B.n464 71.676
R1142 B.n560 B.n465 71.676
R1143 B.n556 B.n466 71.676
R1144 B.n552 B.n467 71.676
R1145 B.n548 B.n468 71.676
R1146 B.n544 B.n469 71.676
R1147 B.n540 B.n470 71.676
R1148 B.n536 B.n471 71.676
R1149 B.n532 B.n472 71.676
R1150 B.n528 B.n473 71.676
R1151 B.n524 B.n474 71.676
R1152 B.n520 B.n475 71.676
R1153 B.n516 B.n476 71.676
R1154 B.n512 B.n477 71.676
R1155 B.n508 B.n478 71.676
R1156 B.n504 B.n479 71.676
R1157 B.n500 B.n480 71.676
R1158 B.n496 B.n481 71.676
R1159 B.n492 B.n482 71.676
R1160 B.n909 B.n908 71.676
R1161 B.n909 B.n2 71.676
R1162 B.n235 B.n116 59.5399
R1163 B.n256 B.n114 59.5399
R1164 B.n490 B.n489 59.5399
R1165 B.n487 B.n486 59.5399
R1166 B.n749 B.n415 50.1994
R1167 B.n857 B.n43 50.1994
R1168 B.n756 B.n415 31.3172
R1169 B.n756 B.n411 31.3172
R1170 B.n762 B.n411 31.3172
R1171 B.n762 B.n407 31.3172
R1172 B.n768 B.n407 31.3172
R1173 B.n774 B.n403 31.3172
R1174 B.n774 B.n399 31.3172
R1175 B.n780 B.n399 31.3172
R1176 B.n780 B.n395 31.3172
R1177 B.n787 B.n395 31.3172
R1178 B.n787 B.n786 31.3172
R1179 B.n793 B.n388 31.3172
R1180 B.n800 B.n388 31.3172
R1181 B.n800 B.n799 31.3172
R1182 B.n806 B.n381 31.3172
R1183 B.n813 B.n381 31.3172
R1184 B.n813 B.t3 31.3172
R1185 B.n819 B.t3 31.3172
R1186 B.n819 B.n4 31.3172
R1187 B.n907 B.n4 31.3172
R1188 B.n907 B.n906 31.3172
R1189 B.n906 B.n905 31.3172
R1190 B.n905 B.n8 31.3172
R1191 B.t2 B.n8 31.3172
R1192 B.n898 B.t2 31.3172
R1193 B.n898 B.n897 31.3172
R1194 B.n897 B.n896 31.3172
R1195 B.n890 B.n18 31.3172
R1196 B.n890 B.n889 31.3172
R1197 B.n889 B.n888 31.3172
R1198 B.n882 B.n25 31.3172
R1199 B.n882 B.n881 31.3172
R1200 B.n881 B.n880 31.3172
R1201 B.n880 B.n29 31.3172
R1202 B.n874 B.n29 31.3172
R1203 B.n874 B.n873 31.3172
R1204 B.n872 B.n36 31.3172
R1205 B.n866 B.n36 31.3172
R1206 B.n866 B.n865 31.3172
R1207 B.n865 B.n864 31.3172
R1208 B.n864 B.n43 31.3172
R1209 B.n753 B.n752 28.5664
R1210 B.n491 B.n413 28.5664
R1211 B.n861 B.n860 28.5664
R1212 B.n854 B.n853 28.5664
R1213 B.n116 B.n115 25.0187
R1214 B.n114 B.n113 25.0187
R1215 B.n489 B.n488 25.0187
R1216 B.n486 B.n485 25.0187
R1217 B.n806 B.t4 24.8697
R1218 B.n896 B.t0 24.8697
R1219 B.t7 B.n403 18.4221
R1220 B.n793 B.t5 18.4221
R1221 B.n888 B.t1 18.4221
R1222 B.n873 B.t14 18.4221
R1223 B B.n910 18.0485
R1224 B.n768 B.t7 12.8956
R1225 B.n786 B.t5 12.8956
R1226 B.n25 B.t1 12.8956
R1227 B.t14 B.n872 12.8956
R1228 B.n754 B.n753 10.6151
R1229 B.n754 B.n409 10.6151
R1230 B.n764 B.n409 10.6151
R1231 B.n765 B.n764 10.6151
R1232 B.n766 B.n765 10.6151
R1233 B.n766 B.n401 10.6151
R1234 B.n776 B.n401 10.6151
R1235 B.n777 B.n776 10.6151
R1236 B.n778 B.n777 10.6151
R1237 B.n778 B.n393 10.6151
R1238 B.n789 B.n393 10.6151
R1239 B.n790 B.n789 10.6151
R1240 B.n791 B.n790 10.6151
R1241 B.n791 B.n386 10.6151
R1242 B.n802 B.n386 10.6151
R1243 B.n803 B.n802 10.6151
R1244 B.n804 B.n803 10.6151
R1245 B.n804 B.n379 10.6151
R1246 B.n815 B.n379 10.6151
R1247 B.n816 B.n815 10.6151
R1248 B.n817 B.n816 10.6151
R1249 B.n817 B.n0 10.6151
R1250 B.n752 B.n417 10.6151
R1251 B.n747 B.n417 10.6151
R1252 B.n747 B.n746 10.6151
R1253 B.n746 B.n745 10.6151
R1254 B.n745 B.n742 10.6151
R1255 B.n742 B.n741 10.6151
R1256 B.n741 B.n738 10.6151
R1257 B.n738 B.n737 10.6151
R1258 B.n737 B.n734 10.6151
R1259 B.n734 B.n733 10.6151
R1260 B.n733 B.n730 10.6151
R1261 B.n730 B.n729 10.6151
R1262 B.n729 B.n726 10.6151
R1263 B.n726 B.n725 10.6151
R1264 B.n725 B.n722 10.6151
R1265 B.n722 B.n721 10.6151
R1266 B.n721 B.n718 10.6151
R1267 B.n718 B.n717 10.6151
R1268 B.n717 B.n714 10.6151
R1269 B.n714 B.n713 10.6151
R1270 B.n713 B.n710 10.6151
R1271 B.n710 B.n709 10.6151
R1272 B.n709 B.n706 10.6151
R1273 B.n706 B.n705 10.6151
R1274 B.n705 B.n702 10.6151
R1275 B.n702 B.n701 10.6151
R1276 B.n701 B.n698 10.6151
R1277 B.n698 B.n697 10.6151
R1278 B.n697 B.n694 10.6151
R1279 B.n694 B.n693 10.6151
R1280 B.n693 B.n690 10.6151
R1281 B.n690 B.n689 10.6151
R1282 B.n689 B.n686 10.6151
R1283 B.n686 B.n685 10.6151
R1284 B.n685 B.n682 10.6151
R1285 B.n682 B.n681 10.6151
R1286 B.n681 B.n678 10.6151
R1287 B.n678 B.n677 10.6151
R1288 B.n677 B.n674 10.6151
R1289 B.n674 B.n673 10.6151
R1290 B.n673 B.n670 10.6151
R1291 B.n670 B.n669 10.6151
R1292 B.n669 B.n666 10.6151
R1293 B.n666 B.n665 10.6151
R1294 B.n665 B.n662 10.6151
R1295 B.n662 B.n661 10.6151
R1296 B.n661 B.n658 10.6151
R1297 B.n658 B.n657 10.6151
R1298 B.n657 B.n654 10.6151
R1299 B.n654 B.n653 10.6151
R1300 B.n653 B.n650 10.6151
R1301 B.n650 B.n649 10.6151
R1302 B.n649 B.n646 10.6151
R1303 B.n646 B.n645 10.6151
R1304 B.n645 B.n642 10.6151
R1305 B.n642 B.n641 10.6151
R1306 B.n641 B.n638 10.6151
R1307 B.n638 B.n637 10.6151
R1308 B.n637 B.n634 10.6151
R1309 B.n634 B.n633 10.6151
R1310 B.n630 B.n629 10.6151
R1311 B.n629 B.n626 10.6151
R1312 B.n626 B.n625 10.6151
R1313 B.n625 B.n622 10.6151
R1314 B.n622 B.n621 10.6151
R1315 B.n621 B.n618 10.6151
R1316 B.n618 B.n617 10.6151
R1317 B.n617 B.n614 10.6151
R1318 B.n614 B.n613 10.6151
R1319 B.n610 B.n609 10.6151
R1320 B.n609 B.n606 10.6151
R1321 B.n606 B.n605 10.6151
R1322 B.n605 B.n602 10.6151
R1323 B.n602 B.n601 10.6151
R1324 B.n601 B.n598 10.6151
R1325 B.n598 B.n597 10.6151
R1326 B.n597 B.n594 10.6151
R1327 B.n594 B.n593 10.6151
R1328 B.n593 B.n590 10.6151
R1329 B.n590 B.n589 10.6151
R1330 B.n589 B.n586 10.6151
R1331 B.n586 B.n585 10.6151
R1332 B.n585 B.n582 10.6151
R1333 B.n582 B.n581 10.6151
R1334 B.n581 B.n578 10.6151
R1335 B.n578 B.n577 10.6151
R1336 B.n577 B.n574 10.6151
R1337 B.n574 B.n573 10.6151
R1338 B.n573 B.n570 10.6151
R1339 B.n570 B.n569 10.6151
R1340 B.n569 B.n566 10.6151
R1341 B.n566 B.n565 10.6151
R1342 B.n565 B.n562 10.6151
R1343 B.n562 B.n561 10.6151
R1344 B.n561 B.n558 10.6151
R1345 B.n558 B.n557 10.6151
R1346 B.n557 B.n554 10.6151
R1347 B.n554 B.n553 10.6151
R1348 B.n553 B.n550 10.6151
R1349 B.n550 B.n549 10.6151
R1350 B.n549 B.n546 10.6151
R1351 B.n546 B.n545 10.6151
R1352 B.n545 B.n542 10.6151
R1353 B.n542 B.n541 10.6151
R1354 B.n541 B.n538 10.6151
R1355 B.n538 B.n537 10.6151
R1356 B.n537 B.n534 10.6151
R1357 B.n534 B.n533 10.6151
R1358 B.n533 B.n530 10.6151
R1359 B.n530 B.n529 10.6151
R1360 B.n529 B.n526 10.6151
R1361 B.n526 B.n525 10.6151
R1362 B.n525 B.n522 10.6151
R1363 B.n522 B.n521 10.6151
R1364 B.n521 B.n518 10.6151
R1365 B.n518 B.n517 10.6151
R1366 B.n517 B.n514 10.6151
R1367 B.n514 B.n513 10.6151
R1368 B.n513 B.n510 10.6151
R1369 B.n510 B.n509 10.6151
R1370 B.n509 B.n506 10.6151
R1371 B.n506 B.n505 10.6151
R1372 B.n505 B.n502 10.6151
R1373 B.n502 B.n501 10.6151
R1374 B.n501 B.n498 10.6151
R1375 B.n498 B.n497 10.6151
R1376 B.n497 B.n494 10.6151
R1377 B.n494 B.n493 10.6151
R1378 B.n493 B.n491 10.6151
R1379 B.n758 B.n413 10.6151
R1380 B.n759 B.n758 10.6151
R1381 B.n760 B.n759 10.6151
R1382 B.n760 B.n405 10.6151
R1383 B.n770 B.n405 10.6151
R1384 B.n771 B.n770 10.6151
R1385 B.n772 B.n771 10.6151
R1386 B.n772 B.n397 10.6151
R1387 B.n782 B.n397 10.6151
R1388 B.n783 B.n782 10.6151
R1389 B.n784 B.n783 10.6151
R1390 B.n784 B.n390 10.6151
R1391 B.n795 B.n390 10.6151
R1392 B.n796 B.n795 10.6151
R1393 B.n797 B.n796 10.6151
R1394 B.n797 B.n383 10.6151
R1395 B.n808 B.n383 10.6151
R1396 B.n809 B.n808 10.6151
R1397 B.n811 B.n809 10.6151
R1398 B.n811 B.n810 10.6151
R1399 B.n810 B.n376 10.6151
R1400 B.n822 B.n376 10.6151
R1401 B.n823 B.n822 10.6151
R1402 B.n824 B.n823 10.6151
R1403 B.n825 B.n824 10.6151
R1404 B.n826 B.n825 10.6151
R1405 B.n829 B.n826 10.6151
R1406 B.n830 B.n829 10.6151
R1407 B.n831 B.n830 10.6151
R1408 B.n832 B.n831 10.6151
R1409 B.n834 B.n832 10.6151
R1410 B.n835 B.n834 10.6151
R1411 B.n836 B.n835 10.6151
R1412 B.n837 B.n836 10.6151
R1413 B.n839 B.n837 10.6151
R1414 B.n840 B.n839 10.6151
R1415 B.n841 B.n840 10.6151
R1416 B.n842 B.n841 10.6151
R1417 B.n844 B.n842 10.6151
R1418 B.n845 B.n844 10.6151
R1419 B.n846 B.n845 10.6151
R1420 B.n847 B.n846 10.6151
R1421 B.n849 B.n847 10.6151
R1422 B.n850 B.n849 10.6151
R1423 B.n851 B.n850 10.6151
R1424 B.n852 B.n851 10.6151
R1425 B.n853 B.n852 10.6151
R1426 B.n902 B.n1 10.6151
R1427 B.n902 B.n901 10.6151
R1428 B.n901 B.n900 10.6151
R1429 B.n900 B.n10 10.6151
R1430 B.n894 B.n10 10.6151
R1431 B.n894 B.n893 10.6151
R1432 B.n893 B.n892 10.6151
R1433 B.n892 B.n16 10.6151
R1434 B.n886 B.n16 10.6151
R1435 B.n886 B.n885 10.6151
R1436 B.n885 B.n884 10.6151
R1437 B.n884 B.n23 10.6151
R1438 B.n878 B.n23 10.6151
R1439 B.n878 B.n877 10.6151
R1440 B.n877 B.n876 10.6151
R1441 B.n876 B.n31 10.6151
R1442 B.n870 B.n31 10.6151
R1443 B.n870 B.n869 10.6151
R1444 B.n869 B.n868 10.6151
R1445 B.n868 B.n38 10.6151
R1446 B.n862 B.n38 10.6151
R1447 B.n862 B.n861 10.6151
R1448 B.n860 B.n45 10.6151
R1449 B.n118 B.n45 10.6151
R1450 B.n119 B.n118 10.6151
R1451 B.n122 B.n119 10.6151
R1452 B.n123 B.n122 10.6151
R1453 B.n126 B.n123 10.6151
R1454 B.n127 B.n126 10.6151
R1455 B.n130 B.n127 10.6151
R1456 B.n131 B.n130 10.6151
R1457 B.n134 B.n131 10.6151
R1458 B.n135 B.n134 10.6151
R1459 B.n138 B.n135 10.6151
R1460 B.n139 B.n138 10.6151
R1461 B.n142 B.n139 10.6151
R1462 B.n143 B.n142 10.6151
R1463 B.n146 B.n143 10.6151
R1464 B.n147 B.n146 10.6151
R1465 B.n150 B.n147 10.6151
R1466 B.n151 B.n150 10.6151
R1467 B.n154 B.n151 10.6151
R1468 B.n155 B.n154 10.6151
R1469 B.n158 B.n155 10.6151
R1470 B.n159 B.n158 10.6151
R1471 B.n162 B.n159 10.6151
R1472 B.n163 B.n162 10.6151
R1473 B.n166 B.n163 10.6151
R1474 B.n167 B.n166 10.6151
R1475 B.n170 B.n167 10.6151
R1476 B.n171 B.n170 10.6151
R1477 B.n174 B.n171 10.6151
R1478 B.n175 B.n174 10.6151
R1479 B.n178 B.n175 10.6151
R1480 B.n179 B.n178 10.6151
R1481 B.n182 B.n179 10.6151
R1482 B.n183 B.n182 10.6151
R1483 B.n186 B.n183 10.6151
R1484 B.n187 B.n186 10.6151
R1485 B.n190 B.n187 10.6151
R1486 B.n191 B.n190 10.6151
R1487 B.n194 B.n191 10.6151
R1488 B.n195 B.n194 10.6151
R1489 B.n198 B.n195 10.6151
R1490 B.n199 B.n198 10.6151
R1491 B.n202 B.n199 10.6151
R1492 B.n203 B.n202 10.6151
R1493 B.n206 B.n203 10.6151
R1494 B.n207 B.n206 10.6151
R1495 B.n210 B.n207 10.6151
R1496 B.n211 B.n210 10.6151
R1497 B.n214 B.n211 10.6151
R1498 B.n215 B.n214 10.6151
R1499 B.n218 B.n215 10.6151
R1500 B.n219 B.n218 10.6151
R1501 B.n222 B.n219 10.6151
R1502 B.n223 B.n222 10.6151
R1503 B.n226 B.n223 10.6151
R1504 B.n227 B.n226 10.6151
R1505 B.n230 B.n227 10.6151
R1506 B.n231 B.n230 10.6151
R1507 B.n234 B.n231 10.6151
R1508 B.n239 B.n236 10.6151
R1509 B.n240 B.n239 10.6151
R1510 B.n243 B.n240 10.6151
R1511 B.n244 B.n243 10.6151
R1512 B.n247 B.n244 10.6151
R1513 B.n248 B.n247 10.6151
R1514 B.n251 B.n248 10.6151
R1515 B.n252 B.n251 10.6151
R1516 B.n255 B.n252 10.6151
R1517 B.n260 B.n257 10.6151
R1518 B.n261 B.n260 10.6151
R1519 B.n264 B.n261 10.6151
R1520 B.n265 B.n264 10.6151
R1521 B.n268 B.n265 10.6151
R1522 B.n269 B.n268 10.6151
R1523 B.n272 B.n269 10.6151
R1524 B.n273 B.n272 10.6151
R1525 B.n276 B.n273 10.6151
R1526 B.n277 B.n276 10.6151
R1527 B.n280 B.n277 10.6151
R1528 B.n281 B.n280 10.6151
R1529 B.n284 B.n281 10.6151
R1530 B.n285 B.n284 10.6151
R1531 B.n288 B.n285 10.6151
R1532 B.n289 B.n288 10.6151
R1533 B.n292 B.n289 10.6151
R1534 B.n293 B.n292 10.6151
R1535 B.n296 B.n293 10.6151
R1536 B.n297 B.n296 10.6151
R1537 B.n300 B.n297 10.6151
R1538 B.n301 B.n300 10.6151
R1539 B.n304 B.n301 10.6151
R1540 B.n305 B.n304 10.6151
R1541 B.n308 B.n305 10.6151
R1542 B.n309 B.n308 10.6151
R1543 B.n312 B.n309 10.6151
R1544 B.n313 B.n312 10.6151
R1545 B.n316 B.n313 10.6151
R1546 B.n317 B.n316 10.6151
R1547 B.n320 B.n317 10.6151
R1548 B.n321 B.n320 10.6151
R1549 B.n324 B.n321 10.6151
R1550 B.n325 B.n324 10.6151
R1551 B.n328 B.n325 10.6151
R1552 B.n329 B.n328 10.6151
R1553 B.n332 B.n329 10.6151
R1554 B.n333 B.n332 10.6151
R1555 B.n336 B.n333 10.6151
R1556 B.n337 B.n336 10.6151
R1557 B.n340 B.n337 10.6151
R1558 B.n341 B.n340 10.6151
R1559 B.n344 B.n341 10.6151
R1560 B.n345 B.n344 10.6151
R1561 B.n348 B.n345 10.6151
R1562 B.n349 B.n348 10.6151
R1563 B.n352 B.n349 10.6151
R1564 B.n353 B.n352 10.6151
R1565 B.n356 B.n353 10.6151
R1566 B.n357 B.n356 10.6151
R1567 B.n360 B.n357 10.6151
R1568 B.n361 B.n360 10.6151
R1569 B.n364 B.n361 10.6151
R1570 B.n365 B.n364 10.6151
R1571 B.n368 B.n365 10.6151
R1572 B.n369 B.n368 10.6151
R1573 B.n372 B.n369 10.6151
R1574 B.n374 B.n372 10.6151
R1575 B.n375 B.n374 10.6151
R1576 B.n854 B.n375 10.6151
R1577 B.n633 B.n487 9.36635
R1578 B.n610 B.n490 9.36635
R1579 B.n235 B.n234 9.36635
R1580 B.n257 B.n256 9.36635
R1581 B.n910 B.n0 8.11757
R1582 B.n910 B.n1 8.11757
R1583 B.n799 B.t4 6.44806
R1584 B.n18 B.t0 6.44806
R1585 B.n630 B.n487 1.24928
R1586 B.n613 B.n490 1.24928
R1587 B.n236 B.n235 1.24928
R1588 B.n256 B.n255 1.24928
R1589 VN.n2 VN.t3 527.299
R1590 VN.n10 VN.t4 527.299
R1591 VN.n6 VN.t0 508.36
R1592 VN.n14 VN.t5 508.36
R1593 VN.n1 VN.t2 467.19
R1594 VN.n9 VN.t1 467.19
R1595 VN.n7 VN.n6 161.3
R1596 VN.n15 VN.n14 161.3
R1597 VN.n13 VN.n8 161.3
R1598 VN.n12 VN.n11 161.3
R1599 VN.n5 VN.n0 161.3
R1600 VN.n4 VN.n3 161.3
R1601 VN.n5 VN.n4 50.6917
R1602 VN.n13 VN.n12 50.6917
R1603 VN VN.n15 47.6804
R1604 VN.n11 VN.n10 43.2502
R1605 VN.n3 VN.n2 43.2502
R1606 VN.n2 VN.n1 42.2819
R1607 VN.n10 VN.n9 42.2819
R1608 VN.n4 VN.n1 12.234
R1609 VN.n12 VN.n9 12.234
R1610 VN.n6 VN.n5 8.76414
R1611 VN.n14 VN.n13 8.76414
R1612 VN.n15 VN.n8 0.189894
R1613 VN.n11 VN.n8 0.189894
R1614 VN.n3 VN.n0 0.189894
R1615 VN.n7 VN.n0 0.189894
R1616 VN VN.n7 0.0516364
R1617 VDD2.n1 VDD2.t2 62.6705
R1618 VDD2.n2 VDD2.t0 61.8919
R1619 VDD2.n1 VDD2.n0 61.0504
R1620 VDD2 VDD2.n3 61.0477
R1621 VDD2.n2 VDD2.n1 43.3726
R1622 VDD2.n3 VDD2.t4 1.06444
R1623 VDD2.n3 VDD2.t1 1.06444
R1624 VDD2.n0 VDD2.t3 1.06444
R1625 VDD2.n0 VDD2.t5 1.06444
R1626 VDD2 VDD2.n2 0.892741
C0 VTAIL VN 7.06685f
C1 VDD1 VN 0.148442f
C2 VDD2 VTAIL 12.7196f
C3 VDD2 VDD1 0.806882f
C4 VTAIL VDD1 12.6861f
C5 VP VN 6.55428f
C6 VDD2 VP 0.320412f
C7 VP VTAIL 7.08162f
C8 VDD2 VN 7.57481f
C9 VP VDD1 7.74053f
C10 VDD2 B 5.879022f
C11 VDD1 B 6.125343f
C12 VTAIL B 9.097461f
C13 VN B 9.118099f
C14 VP B 6.990656f
C15 VDD2.t2 B 3.84671f
C16 VDD2.t3 B 0.329508f
C17 VDD2.t5 B 0.329508f
C18 VDD2.n0 B 3.00668f
C19 VDD2.n1 B 2.34329f
C20 VDD2.t0 B 3.84282f
C21 VDD2.n2 B 2.56467f
C22 VDD2.t4 B 0.329508f
C23 VDD2.t1 B 0.329508f
C24 VDD2.n3 B 3.00665f
C25 VN.n0 B 0.040113f
C26 VN.t2 B 1.97238f
C27 VN.n1 B 0.74608f
C28 VN.t3 B 2.05886f
C29 VN.n2 B 0.757415f
C30 VN.n3 B 0.172934f
C31 VN.n4 B 0.054778f
C32 VN.n5 B 0.014355f
C33 VN.t0 B 2.03137f
C34 VN.n6 B 0.754612f
C35 VN.n7 B 0.031086f
C36 VN.n8 B 0.040113f
C37 VN.t1 B 1.97238f
C38 VN.n9 B 0.74608f
C39 VN.t4 B 2.05886f
C40 VN.n10 B 0.757415f
C41 VN.n11 B 0.172934f
C42 VN.n12 B 0.054778f
C43 VN.n13 B 0.014355f
C44 VN.t5 B 2.03137f
C45 VN.n14 B 0.754612f
C46 VN.n15 B 2.02982f
C47 VTAIL.t2 B 0.336332f
C48 VTAIL.t0 B 0.336332f
C49 VTAIL.n0 B 2.99749f
C50 VTAIL.n1 B 0.330239f
C51 VTAIL.t6 B 3.83055f
C52 VTAIL.n2 B 0.471631f
C53 VTAIL.t8 B 0.336332f
C54 VTAIL.t9 B 0.336332f
C55 VTAIL.n3 B 2.99749f
C56 VTAIL.n4 B 1.96864f
C57 VTAIL.t11 B 0.336332f
C58 VTAIL.t4 B 0.336332f
C59 VTAIL.n5 B 2.9975f
C60 VTAIL.n6 B 1.96864f
C61 VTAIL.t3 B 3.83057f
C62 VTAIL.n7 B 0.471609f
C63 VTAIL.t7 B 0.336332f
C64 VTAIL.t10 B 0.336332f
C65 VTAIL.n8 B 2.9975f
C66 VTAIL.n9 B 0.38741f
C67 VTAIL.t5 B 3.83055f
C68 VTAIL.n10 B 1.97091f
C69 VTAIL.t1 B 3.83055f
C70 VTAIL.n11 B 1.94613f
C71 VDD1.t4 B 3.85064f
C72 VDD1.t5 B 3.84996f
C73 VDD1.t3 B 0.329786f
C74 VDD1.t2 B 0.329786f
C75 VDD1.n0 B 3.00922f
C76 VDD1.n1 B 2.42185f
C77 VDD1.t0 B 0.329786f
C78 VDD1.t1 B 0.329786f
C79 VDD1.n2 B 3.00814f
C80 VDD1.n3 B 2.54338f
C81 VP.n0 B 0.040408f
C82 VP.t1 B 1.9869f
C83 VP.n1 B 0.71156f
C84 VP.n2 B 0.040408f
C85 VP.n3 B 0.040408f
C86 VP.t5 B 2.04633f
C87 VP.t0 B 1.9869f
C88 VP.n4 B 0.751572f
C89 VP.t3 B 2.07401f
C90 VP.n5 B 0.76299f
C91 VP.n6 B 0.174207f
C92 VP.n7 B 0.055181f
C93 VP.n8 B 0.01446f
C94 VP.n9 B 0.760168f
C95 VP.n10 B 2.01842f
C96 VP.n11 B 2.04913f
C97 VP.t2 B 2.04633f
C98 VP.n12 B 0.760168f
C99 VP.n13 B 0.01446f
C100 VP.n14 B 0.055181f
C101 VP.n15 B 0.040408f
C102 VP.n16 B 0.040408f
C103 VP.n17 B 0.055181f
C104 VP.n18 B 0.01446f
C105 VP.t4 B 2.04633f
C106 VP.n19 B 0.760168f
C107 VP.n20 B 0.031315f
.ends

