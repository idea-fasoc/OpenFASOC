* NGSPICE file created from diff_pair_sample_1178.ext - technology: sky130A

.subckt diff_pair_sample_1178 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=0 ps=0 w=17.9 l=1.8
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=0 ps=0 w=17.9 l=1.8
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=6.981 ps=36.58 w=17.9 l=1.8
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=0 ps=0 w=17.9 l=1.8
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=6.981 ps=36.58 w=17.9 l=1.8
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=6.981 ps=36.58 w=17.9 l=1.8
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=6.981 ps=36.58 w=17.9 l=1.8
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.981 pd=36.58 as=0 ps=0 w=17.9 l=1.8
R0 B.n815 B.n814 585
R1 B.n362 B.n105 585
R2 B.n361 B.n360 585
R3 B.n359 B.n358 585
R4 B.n357 B.n356 585
R5 B.n355 B.n354 585
R6 B.n353 B.n352 585
R7 B.n351 B.n350 585
R8 B.n349 B.n348 585
R9 B.n347 B.n346 585
R10 B.n345 B.n344 585
R11 B.n343 B.n342 585
R12 B.n341 B.n340 585
R13 B.n339 B.n338 585
R14 B.n337 B.n336 585
R15 B.n335 B.n334 585
R16 B.n333 B.n332 585
R17 B.n331 B.n330 585
R18 B.n329 B.n328 585
R19 B.n327 B.n326 585
R20 B.n325 B.n324 585
R21 B.n323 B.n322 585
R22 B.n321 B.n320 585
R23 B.n319 B.n318 585
R24 B.n317 B.n316 585
R25 B.n315 B.n314 585
R26 B.n313 B.n312 585
R27 B.n311 B.n310 585
R28 B.n309 B.n308 585
R29 B.n307 B.n306 585
R30 B.n305 B.n304 585
R31 B.n303 B.n302 585
R32 B.n301 B.n300 585
R33 B.n299 B.n298 585
R34 B.n297 B.n296 585
R35 B.n295 B.n294 585
R36 B.n293 B.n292 585
R37 B.n291 B.n290 585
R38 B.n289 B.n288 585
R39 B.n287 B.n286 585
R40 B.n285 B.n284 585
R41 B.n283 B.n282 585
R42 B.n281 B.n280 585
R43 B.n279 B.n278 585
R44 B.n277 B.n276 585
R45 B.n275 B.n274 585
R46 B.n273 B.n272 585
R47 B.n271 B.n270 585
R48 B.n269 B.n268 585
R49 B.n267 B.n266 585
R50 B.n265 B.n264 585
R51 B.n263 B.n262 585
R52 B.n261 B.n260 585
R53 B.n259 B.n258 585
R54 B.n257 B.n256 585
R55 B.n255 B.n254 585
R56 B.n253 B.n252 585
R57 B.n251 B.n250 585
R58 B.n249 B.n248 585
R59 B.n246 B.n245 585
R60 B.n244 B.n243 585
R61 B.n242 B.n241 585
R62 B.n240 B.n239 585
R63 B.n238 B.n237 585
R64 B.n236 B.n235 585
R65 B.n234 B.n233 585
R66 B.n232 B.n231 585
R67 B.n230 B.n229 585
R68 B.n228 B.n227 585
R69 B.n225 B.n224 585
R70 B.n223 B.n222 585
R71 B.n221 B.n220 585
R72 B.n219 B.n218 585
R73 B.n217 B.n216 585
R74 B.n215 B.n214 585
R75 B.n213 B.n212 585
R76 B.n211 B.n210 585
R77 B.n209 B.n208 585
R78 B.n207 B.n206 585
R79 B.n205 B.n204 585
R80 B.n203 B.n202 585
R81 B.n201 B.n200 585
R82 B.n199 B.n198 585
R83 B.n197 B.n196 585
R84 B.n195 B.n194 585
R85 B.n193 B.n192 585
R86 B.n191 B.n190 585
R87 B.n189 B.n188 585
R88 B.n187 B.n186 585
R89 B.n185 B.n184 585
R90 B.n183 B.n182 585
R91 B.n181 B.n180 585
R92 B.n179 B.n178 585
R93 B.n177 B.n176 585
R94 B.n175 B.n174 585
R95 B.n173 B.n172 585
R96 B.n171 B.n170 585
R97 B.n169 B.n168 585
R98 B.n167 B.n166 585
R99 B.n165 B.n164 585
R100 B.n163 B.n162 585
R101 B.n161 B.n160 585
R102 B.n159 B.n158 585
R103 B.n157 B.n156 585
R104 B.n155 B.n154 585
R105 B.n153 B.n152 585
R106 B.n151 B.n150 585
R107 B.n149 B.n148 585
R108 B.n147 B.n146 585
R109 B.n145 B.n144 585
R110 B.n143 B.n142 585
R111 B.n141 B.n140 585
R112 B.n139 B.n138 585
R113 B.n137 B.n136 585
R114 B.n135 B.n134 585
R115 B.n133 B.n132 585
R116 B.n131 B.n130 585
R117 B.n129 B.n128 585
R118 B.n127 B.n126 585
R119 B.n125 B.n124 585
R120 B.n123 B.n122 585
R121 B.n121 B.n120 585
R122 B.n119 B.n118 585
R123 B.n117 B.n116 585
R124 B.n115 B.n114 585
R125 B.n113 B.n112 585
R126 B.n111 B.n110 585
R127 B.n40 B.n39 585
R128 B.n813 B.n41 585
R129 B.n818 B.n41 585
R130 B.n812 B.n811 585
R131 B.n811 B.n37 585
R132 B.n810 B.n36 585
R133 B.n824 B.n36 585
R134 B.n809 B.n35 585
R135 B.n825 B.n35 585
R136 B.n808 B.n34 585
R137 B.n826 B.n34 585
R138 B.n807 B.n806 585
R139 B.n806 B.n30 585
R140 B.n805 B.n29 585
R141 B.n832 B.n29 585
R142 B.n804 B.n28 585
R143 B.n833 B.n28 585
R144 B.n803 B.n27 585
R145 B.n834 B.n27 585
R146 B.n802 B.n801 585
R147 B.n801 B.n23 585
R148 B.n800 B.n22 585
R149 B.n840 B.n22 585
R150 B.n799 B.n21 585
R151 B.n841 B.n21 585
R152 B.n798 B.n20 585
R153 B.n842 B.n20 585
R154 B.n797 B.n796 585
R155 B.n796 B.n16 585
R156 B.n795 B.n15 585
R157 B.n848 B.n15 585
R158 B.n794 B.n14 585
R159 B.n849 B.n14 585
R160 B.n793 B.n13 585
R161 B.n850 B.n13 585
R162 B.n792 B.n791 585
R163 B.n791 B.n12 585
R164 B.n790 B.n789 585
R165 B.n790 B.n8 585
R166 B.n788 B.n7 585
R167 B.n857 B.n7 585
R168 B.n787 B.n6 585
R169 B.n858 B.n6 585
R170 B.n786 B.n5 585
R171 B.n859 B.n5 585
R172 B.n785 B.n784 585
R173 B.n784 B.n4 585
R174 B.n783 B.n363 585
R175 B.n783 B.n782 585
R176 B.n773 B.n364 585
R177 B.n365 B.n364 585
R178 B.n775 B.n774 585
R179 B.n776 B.n775 585
R180 B.n772 B.n369 585
R181 B.n373 B.n369 585
R182 B.n771 B.n770 585
R183 B.n770 B.n769 585
R184 B.n371 B.n370 585
R185 B.n372 B.n371 585
R186 B.n762 B.n761 585
R187 B.n763 B.n762 585
R188 B.n760 B.n378 585
R189 B.n378 B.n377 585
R190 B.n759 B.n758 585
R191 B.n758 B.n757 585
R192 B.n380 B.n379 585
R193 B.n381 B.n380 585
R194 B.n750 B.n749 585
R195 B.n751 B.n750 585
R196 B.n748 B.n386 585
R197 B.n386 B.n385 585
R198 B.n747 B.n746 585
R199 B.n746 B.n745 585
R200 B.n388 B.n387 585
R201 B.n389 B.n388 585
R202 B.n738 B.n737 585
R203 B.n739 B.n738 585
R204 B.n736 B.n394 585
R205 B.n394 B.n393 585
R206 B.n735 B.n734 585
R207 B.n734 B.n733 585
R208 B.n396 B.n395 585
R209 B.n397 B.n396 585
R210 B.n726 B.n725 585
R211 B.n727 B.n726 585
R212 B.n400 B.n399 585
R213 B.n473 B.n472 585
R214 B.n474 B.n470 585
R215 B.n470 B.n401 585
R216 B.n476 B.n475 585
R217 B.n478 B.n469 585
R218 B.n481 B.n480 585
R219 B.n482 B.n468 585
R220 B.n484 B.n483 585
R221 B.n486 B.n467 585
R222 B.n489 B.n488 585
R223 B.n490 B.n466 585
R224 B.n492 B.n491 585
R225 B.n494 B.n465 585
R226 B.n497 B.n496 585
R227 B.n498 B.n464 585
R228 B.n500 B.n499 585
R229 B.n502 B.n463 585
R230 B.n505 B.n504 585
R231 B.n506 B.n462 585
R232 B.n508 B.n507 585
R233 B.n510 B.n461 585
R234 B.n513 B.n512 585
R235 B.n514 B.n460 585
R236 B.n516 B.n515 585
R237 B.n518 B.n459 585
R238 B.n521 B.n520 585
R239 B.n522 B.n458 585
R240 B.n524 B.n523 585
R241 B.n526 B.n457 585
R242 B.n529 B.n528 585
R243 B.n530 B.n456 585
R244 B.n532 B.n531 585
R245 B.n534 B.n455 585
R246 B.n537 B.n536 585
R247 B.n538 B.n454 585
R248 B.n540 B.n539 585
R249 B.n542 B.n453 585
R250 B.n545 B.n544 585
R251 B.n546 B.n452 585
R252 B.n548 B.n547 585
R253 B.n550 B.n451 585
R254 B.n553 B.n552 585
R255 B.n554 B.n450 585
R256 B.n556 B.n555 585
R257 B.n558 B.n449 585
R258 B.n561 B.n560 585
R259 B.n562 B.n448 585
R260 B.n564 B.n563 585
R261 B.n566 B.n447 585
R262 B.n569 B.n568 585
R263 B.n570 B.n446 585
R264 B.n572 B.n571 585
R265 B.n574 B.n445 585
R266 B.n577 B.n576 585
R267 B.n578 B.n444 585
R268 B.n580 B.n579 585
R269 B.n582 B.n443 585
R270 B.n585 B.n584 585
R271 B.n586 B.n440 585
R272 B.n589 B.n588 585
R273 B.n591 B.n439 585
R274 B.n594 B.n593 585
R275 B.n595 B.n438 585
R276 B.n597 B.n596 585
R277 B.n599 B.n437 585
R278 B.n602 B.n601 585
R279 B.n603 B.n436 585
R280 B.n605 B.n604 585
R281 B.n607 B.n435 585
R282 B.n610 B.n609 585
R283 B.n611 B.n431 585
R284 B.n613 B.n612 585
R285 B.n615 B.n430 585
R286 B.n618 B.n617 585
R287 B.n619 B.n429 585
R288 B.n621 B.n620 585
R289 B.n623 B.n428 585
R290 B.n626 B.n625 585
R291 B.n627 B.n427 585
R292 B.n629 B.n628 585
R293 B.n631 B.n426 585
R294 B.n634 B.n633 585
R295 B.n635 B.n425 585
R296 B.n637 B.n636 585
R297 B.n639 B.n424 585
R298 B.n642 B.n641 585
R299 B.n643 B.n423 585
R300 B.n645 B.n644 585
R301 B.n647 B.n422 585
R302 B.n650 B.n649 585
R303 B.n651 B.n421 585
R304 B.n653 B.n652 585
R305 B.n655 B.n420 585
R306 B.n658 B.n657 585
R307 B.n659 B.n419 585
R308 B.n661 B.n660 585
R309 B.n663 B.n418 585
R310 B.n666 B.n665 585
R311 B.n667 B.n417 585
R312 B.n669 B.n668 585
R313 B.n671 B.n416 585
R314 B.n674 B.n673 585
R315 B.n675 B.n415 585
R316 B.n677 B.n676 585
R317 B.n679 B.n414 585
R318 B.n682 B.n681 585
R319 B.n683 B.n413 585
R320 B.n685 B.n684 585
R321 B.n687 B.n412 585
R322 B.n690 B.n689 585
R323 B.n691 B.n411 585
R324 B.n693 B.n692 585
R325 B.n695 B.n410 585
R326 B.n698 B.n697 585
R327 B.n699 B.n409 585
R328 B.n701 B.n700 585
R329 B.n703 B.n408 585
R330 B.n706 B.n705 585
R331 B.n707 B.n407 585
R332 B.n709 B.n708 585
R333 B.n711 B.n406 585
R334 B.n714 B.n713 585
R335 B.n715 B.n405 585
R336 B.n717 B.n716 585
R337 B.n719 B.n404 585
R338 B.n720 B.n403 585
R339 B.n723 B.n722 585
R340 B.n724 B.n402 585
R341 B.n402 B.n401 585
R342 B.n729 B.n728 585
R343 B.n728 B.n727 585
R344 B.n730 B.n398 585
R345 B.n398 B.n397 585
R346 B.n732 B.n731 585
R347 B.n733 B.n732 585
R348 B.n392 B.n391 585
R349 B.n393 B.n392 585
R350 B.n741 B.n740 585
R351 B.n740 B.n739 585
R352 B.n742 B.n390 585
R353 B.n390 B.n389 585
R354 B.n744 B.n743 585
R355 B.n745 B.n744 585
R356 B.n384 B.n383 585
R357 B.n385 B.n384 585
R358 B.n753 B.n752 585
R359 B.n752 B.n751 585
R360 B.n754 B.n382 585
R361 B.n382 B.n381 585
R362 B.n756 B.n755 585
R363 B.n757 B.n756 585
R364 B.n376 B.n375 585
R365 B.n377 B.n376 585
R366 B.n765 B.n764 585
R367 B.n764 B.n763 585
R368 B.n766 B.n374 585
R369 B.n374 B.n372 585
R370 B.n768 B.n767 585
R371 B.n769 B.n768 585
R372 B.n368 B.n367 585
R373 B.n373 B.n368 585
R374 B.n778 B.n777 585
R375 B.n777 B.n776 585
R376 B.n779 B.n366 585
R377 B.n366 B.n365 585
R378 B.n781 B.n780 585
R379 B.n782 B.n781 585
R380 B.n3 B.n0 585
R381 B.n4 B.n3 585
R382 B.n856 B.n1 585
R383 B.n857 B.n856 585
R384 B.n855 B.n854 585
R385 B.n855 B.n8 585
R386 B.n853 B.n9 585
R387 B.n12 B.n9 585
R388 B.n852 B.n851 585
R389 B.n851 B.n850 585
R390 B.n11 B.n10 585
R391 B.n849 B.n11 585
R392 B.n847 B.n846 585
R393 B.n848 B.n847 585
R394 B.n845 B.n17 585
R395 B.n17 B.n16 585
R396 B.n844 B.n843 585
R397 B.n843 B.n842 585
R398 B.n19 B.n18 585
R399 B.n841 B.n19 585
R400 B.n839 B.n838 585
R401 B.n840 B.n839 585
R402 B.n837 B.n24 585
R403 B.n24 B.n23 585
R404 B.n836 B.n835 585
R405 B.n835 B.n834 585
R406 B.n26 B.n25 585
R407 B.n833 B.n26 585
R408 B.n831 B.n830 585
R409 B.n832 B.n831 585
R410 B.n829 B.n31 585
R411 B.n31 B.n30 585
R412 B.n828 B.n827 585
R413 B.n827 B.n826 585
R414 B.n33 B.n32 585
R415 B.n825 B.n33 585
R416 B.n823 B.n822 585
R417 B.n824 B.n823 585
R418 B.n821 B.n38 585
R419 B.n38 B.n37 585
R420 B.n820 B.n819 585
R421 B.n819 B.n818 585
R422 B.n860 B.n859 585
R423 B.n858 B.n2 585
R424 B.n819 B.n40 482.89
R425 B.n815 B.n41 482.89
R426 B.n726 B.n402 482.89
R427 B.n728 B.n400 482.89
R428 B.n108 B.t10 446.067
R429 B.n106 B.t2 446.067
R430 B.n432 B.t13 446.067
R431 B.n441 B.t6 446.067
R432 B.n817 B.n816 256.663
R433 B.n817 B.n104 256.663
R434 B.n817 B.n103 256.663
R435 B.n817 B.n102 256.663
R436 B.n817 B.n101 256.663
R437 B.n817 B.n100 256.663
R438 B.n817 B.n99 256.663
R439 B.n817 B.n98 256.663
R440 B.n817 B.n97 256.663
R441 B.n817 B.n96 256.663
R442 B.n817 B.n95 256.663
R443 B.n817 B.n94 256.663
R444 B.n817 B.n93 256.663
R445 B.n817 B.n92 256.663
R446 B.n817 B.n91 256.663
R447 B.n817 B.n90 256.663
R448 B.n817 B.n89 256.663
R449 B.n817 B.n88 256.663
R450 B.n817 B.n87 256.663
R451 B.n817 B.n86 256.663
R452 B.n817 B.n85 256.663
R453 B.n817 B.n84 256.663
R454 B.n817 B.n83 256.663
R455 B.n817 B.n82 256.663
R456 B.n817 B.n81 256.663
R457 B.n817 B.n80 256.663
R458 B.n817 B.n79 256.663
R459 B.n817 B.n78 256.663
R460 B.n817 B.n77 256.663
R461 B.n817 B.n76 256.663
R462 B.n817 B.n75 256.663
R463 B.n817 B.n74 256.663
R464 B.n817 B.n73 256.663
R465 B.n817 B.n72 256.663
R466 B.n817 B.n71 256.663
R467 B.n817 B.n70 256.663
R468 B.n817 B.n69 256.663
R469 B.n817 B.n68 256.663
R470 B.n817 B.n67 256.663
R471 B.n817 B.n66 256.663
R472 B.n817 B.n65 256.663
R473 B.n817 B.n64 256.663
R474 B.n817 B.n63 256.663
R475 B.n817 B.n62 256.663
R476 B.n817 B.n61 256.663
R477 B.n817 B.n60 256.663
R478 B.n817 B.n59 256.663
R479 B.n817 B.n58 256.663
R480 B.n817 B.n57 256.663
R481 B.n817 B.n56 256.663
R482 B.n817 B.n55 256.663
R483 B.n817 B.n54 256.663
R484 B.n817 B.n53 256.663
R485 B.n817 B.n52 256.663
R486 B.n817 B.n51 256.663
R487 B.n817 B.n50 256.663
R488 B.n817 B.n49 256.663
R489 B.n817 B.n48 256.663
R490 B.n817 B.n47 256.663
R491 B.n817 B.n46 256.663
R492 B.n817 B.n45 256.663
R493 B.n817 B.n44 256.663
R494 B.n817 B.n43 256.663
R495 B.n817 B.n42 256.663
R496 B.n471 B.n401 256.663
R497 B.n477 B.n401 256.663
R498 B.n479 B.n401 256.663
R499 B.n485 B.n401 256.663
R500 B.n487 B.n401 256.663
R501 B.n493 B.n401 256.663
R502 B.n495 B.n401 256.663
R503 B.n501 B.n401 256.663
R504 B.n503 B.n401 256.663
R505 B.n509 B.n401 256.663
R506 B.n511 B.n401 256.663
R507 B.n517 B.n401 256.663
R508 B.n519 B.n401 256.663
R509 B.n525 B.n401 256.663
R510 B.n527 B.n401 256.663
R511 B.n533 B.n401 256.663
R512 B.n535 B.n401 256.663
R513 B.n541 B.n401 256.663
R514 B.n543 B.n401 256.663
R515 B.n549 B.n401 256.663
R516 B.n551 B.n401 256.663
R517 B.n557 B.n401 256.663
R518 B.n559 B.n401 256.663
R519 B.n565 B.n401 256.663
R520 B.n567 B.n401 256.663
R521 B.n573 B.n401 256.663
R522 B.n575 B.n401 256.663
R523 B.n581 B.n401 256.663
R524 B.n583 B.n401 256.663
R525 B.n590 B.n401 256.663
R526 B.n592 B.n401 256.663
R527 B.n598 B.n401 256.663
R528 B.n600 B.n401 256.663
R529 B.n606 B.n401 256.663
R530 B.n608 B.n401 256.663
R531 B.n614 B.n401 256.663
R532 B.n616 B.n401 256.663
R533 B.n622 B.n401 256.663
R534 B.n624 B.n401 256.663
R535 B.n630 B.n401 256.663
R536 B.n632 B.n401 256.663
R537 B.n638 B.n401 256.663
R538 B.n640 B.n401 256.663
R539 B.n646 B.n401 256.663
R540 B.n648 B.n401 256.663
R541 B.n654 B.n401 256.663
R542 B.n656 B.n401 256.663
R543 B.n662 B.n401 256.663
R544 B.n664 B.n401 256.663
R545 B.n670 B.n401 256.663
R546 B.n672 B.n401 256.663
R547 B.n678 B.n401 256.663
R548 B.n680 B.n401 256.663
R549 B.n686 B.n401 256.663
R550 B.n688 B.n401 256.663
R551 B.n694 B.n401 256.663
R552 B.n696 B.n401 256.663
R553 B.n702 B.n401 256.663
R554 B.n704 B.n401 256.663
R555 B.n710 B.n401 256.663
R556 B.n712 B.n401 256.663
R557 B.n718 B.n401 256.663
R558 B.n721 B.n401 256.663
R559 B.n862 B.n861 256.663
R560 B.n112 B.n111 163.367
R561 B.n116 B.n115 163.367
R562 B.n120 B.n119 163.367
R563 B.n124 B.n123 163.367
R564 B.n128 B.n127 163.367
R565 B.n132 B.n131 163.367
R566 B.n136 B.n135 163.367
R567 B.n140 B.n139 163.367
R568 B.n144 B.n143 163.367
R569 B.n148 B.n147 163.367
R570 B.n152 B.n151 163.367
R571 B.n156 B.n155 163.367
R572 B.n160 B.n159 163.367
R573 B.n164 B.n163 163.367
R574 B.n168 B.n167 163.367
R575 B.n172 B.n171 163.367
R576 B.n176 B.n175 163.367
R577 B.n180 B.n179 163.367
R578 B.n184 B.n183 163.367
R579 B.n188 B.n187 163.367
R580 B.n192 B.n191 163.367
R581 B.n196 B.n195 163.367
R582 B.n200 B.n199 163.367
R583 B.n204 B.n203 163.367
R584 B.n208 B.n207 163.367
R585 B.n212 B.n211 163.367
R586 B.n216 B.n215 163.367
R587 B.n220 B.n219 163.367
R588 B.n224 B.n223 163.367
R589 B.n229 B.n228 163.367
R590 B.n233 B.n232 163.367
R591 B.n237 B.n236 163.367
R592 B.n241 B.n240 163.367
R593 B.n245 B.n244 163.367
R594 B.n250 B.n249 163.367
R595 B.n254 B.n253 163.367
R596 B.n258 B.n257 163.367
R597 B.n262 B.n261 163.367
R598 B.n266 B.n265 163.367
R599 B.n270 B.n269 163.367
R600 B.n274 B.n273 163.367
R601 B.n278 B.n277 163.367
R602 B.n282 B.n281 163.367
R603 B.n286 B.n285 163.367
R604 B.n290 B.n289 163.367
R605 B.n294 B.n293 163.367
R606 B.n298 B.n297 163.367
R607 B.n302 B.n301 163.367
R608 B.n306 B.n305 163.367
R609 B.n310 B.n309 163.367
R610 B.n314 B.n313 163.367
R611 B.n318 B.n317 163.367
R612 B.n322 B.n321 163.367
R613 B.n326 B.n325 163.367
R614 B.n330 B.n329 163.367
R615 B.n334 B.n333 163.367
R616 B.n338 B.n337 163.367
R617 B.n342 B.n341 163.367
R618 B.n346 B.n345 163.367
R619 B.n350 B.n349 163.367
R620 B.n354 B.n353 163.367
R621 B.n358 B.n357 163.367
R622 B.n360 B.n105 163.367
R623 B.n726 B.n396 163.367
R624 B.n734 B.n396 163.367
R625 B.n734 B.n394 163.367
R626 B.n738 B.n394 163.367
R627 B.n738 B.n388 163.367
R628 B.n746 B.n388 163.367
R629 B.n746 B.n386 163.367
R630 B.n750 B.n386 163.367
R631 B.n750 B.n380 163.367
R632 B.n758 B.n380 163.367
R633 B.n758 B.n378 163.367
R634 B.n762 B.n378 163.367
R635 B.n762 B.n371 163.367
R636 B.n770 B.n371 163.367
R637 B.n770 B.n369 163.367
R638 B.n775 B.n369 163.367
R639 B.n775 B.n364 163.367
R640 B.n783 B.n364 163.367
R641 B.n784 B.n783 163.367
R642 B.n784 B.n5 163.367
R643 B.n6 B.n5 163.367
R644 B.n7 B.n6 163.367
R645 B.n790 B.n7 163.367
R646 B.n791 B.n790 163.367
R647 B.n791 B.n13 163.367
R648 B.n14 B.n13 163.367
R649 B.n15 B.n14 163.367
R650 B.n796 B.n15 163.367
R651 B.n796 B.n20 163.367
R652 B.n21 B.n20 163.367
R653 B.n22 B.n21 163.367
R654 B.n801 B.n22 163.367
R655 B.n801 B.n27 163.367
R656 B.n28 B.n27 163.367
R657 B.n29 B.n28 163.367
R658 B.n806 B.n29 163.367
R659 B.n806 B.n34 163.367
R660 B.n35 B.n34 163.367
R661 B.n36 B.n35 163.367
R662 B.n811 B.n36 163.367
R663 B.n811 B.n41 163.367
R664 B.n472 B.n470 163.367
R665 B.n476 B.n470 163.367
R666 B.n480 B.n478 163.367
R667 B.n484 B.n468 163.367
R668 B.n488 B.n486 163.367
R669 B.n492 B.n466 163.367
R670 B.n496 B.n494 163.367
R671 B.n500 B.n464 163.367
R672 B.n504 B.n502 163.367
R673 B.n508 B.n462 163.367
R674 B.n512 B.n510 163.367
R675 B.n516 B.n460 163.367
R676 B.n520 B.n518 163.367
R677 B.n524 B.n458 163.367
R678 B.n528 B.n526 163.367
R679 B.n532 B.n456 163.367
R680 B.n536 B.n534 163.367
R681 B.n540 B.n454 163.367
R682 B.n544 B.n542 163.367
R683 B.n548 B.n452 163.367
R684 B.n552 B.n550 163.367
R685 B.n556 B.n450 163.367
R686 B.n560 B.n558 163.367
R687 B.n564 B.n448 163.367
R688 B.n568 B.n566 163.367
R689 B.n572 B.n446 163.367
R690 B.n576 B.n574 163.367
R691 B.n580 B.n444 163.367
R692 B.n584 B.n582 163.367
R693 B.n589 B.n440 163.367
R694 B.n593 B.n591 163.367
R695 B.n597 B.n438 163.367
R696 B.n601 B.n599 163.367
R697 B.n605 B.n436 163.367
R698 B.n609 B.n607 163.367
R699 B.n613 B.n431 163.367
R700 B.n617 B.n615 163.367
R701 B.n621 B.n429 163.367
R702 B.n625 B.n623 163.367
R703 B.n629 B.n427 163.367
R704 B.n633 B.n631 163.367
R705 B.n637 B.n425 163.367
R706 B.n641 B.n639 163.367
R707 B.n645 B.n423 163.367
R708 B.n649 B.n647 163.367
R709 B.n653 B.n421 163.367
R710 B.n657 B.n655 163.367
R711 B.n661 B.n419 163.367
R712 B.n665 B.n663 163.367
R713 B.n669 B.n417 163.367
R714 B.n673 B.n671 163.367
R715 B.n677 B.n415 163.367
R716 B.n681 B.n679 163.367
R717 B.n685 B.n413 163.367
R718 B.n689 B.n687 163.367
R719 B.n693 B.n411 163.367
R720 B.n697 B.n695 163.367
R721 B.n701 B.n409 163.367
R722 B.n705 B.n703 163.367
R723 B.n709 B.n407 163.367
R724 B.n713 B.n711 163.367
R725 B.n717 B.n405 163.367
R726 B.n720 B.n719 163.367
R727 B.n722 B.n402 163.367
R728 B.n728 B.n398 163.367
R729 B.n732 B.n398 163.367
R730 B.n732 B.n392 163.367
R731 B.n740 B.n392 163.367
R732 B.n740 B.n390 163.367
R733 B.n744 B.n390 163.367
R734 B.n744 B.n384 163.367
R735 B.n752 B.n384 163.367
R736 B.n752 B.n382 163.367
R737 B.n756 B.n382 163.367
R738 B.n756 B.n376 163.367
R739 B.n764 B.n376 163.367
R740 B.n764 B.n374 163.367
R741 B.n768 B.n374 163.367
R742 B.n768 B.n368 163.367
R743 B.n777 B.n368 163.367
R744 B.n777 B.n366 163.367
R745 B.n781 B.n366 163.367
R746 B.n781 B.n3 163.367
R747 B.n860 B.n3 163.367
R748 B.n856 B.n2 163.367
R749 B.n856 B.n855 163.367
R750 B.n855 B.n9 163.367
R751 B.n851 B.n9 163.367
R752 B.n851 B.n11 163.367
R753 B.n847 B.n11 163.367
R754 B.n847 B.n17 163.367
R755 B.n843 B.n17 163.367
R756 B.n843 B.n19 163.367
R757 B.n839 B.n19 163.367
R758 B.n839 B.n24 163.367
R759 B.n835 B.n24 163.367
R760 B.n835 B.n26 163.367
R761 B.n831 B.n26 163.367
R762 B.n831 B.n31 163.367
R763 B.n827 B.n31 163.367
R764 B.n827 B.n33 163.367
R765 B.n823 B.n33 163.367
R766 B.n823 B.n38 163.367
R767 B.n819 B.n38 163.367
R768 B.n106 B.t4 112.831
R769 B.n432 B.t15 112.831
R770 B.n108 B.t11 112.806
R771 B.n441 B.t9 112.806
R772 B.n42 B.n40 71.676
R773 B.n112 B.n43 71.676
R774 B.n116 B.n44 71.676
R775 B.n120 B.n45 71.676
R776 B.n124 B.n46 71.676
R777 B.n128 B.n47 71.676
R778 B.n132 B.n48 71.676
R779 B.n136 B.n49 71.676
R780 B.n140 B.n50 71.676
R781 B.n144 B.n51 71.676
R782 B.n148 B.n52 71.676
R783 B.n152 B.n53 71.676
R784 B.n156 B.n54 71.676
R785 B.n160 B.n55 71.676
R786 B.n164 B.n56 71.676
R787 B.n168 B.n57 71.676
R788 B.n172 B.n58 71.676
R789 B.n176 B.n59 71.676
R790 B.n180 B.n60 71.676
R791 B.n184 B.n61 71.676
R792 B.n188 B.n62 71.676
R793 B.n192 B.n63 71.676
R794 B.n196 B.n64 71.676
R795 B.n200 B.n65 71.676
R796 B.n204 B.n66 71.676
R797 B.n208 B.n67 71.676
R798 B.n212 B.n68 71.676
R799 B.n216 B.n69 71.676
R800 B.n220 B.n70 71.676
R801 B.n224 B.n71 71.676
R802 B.n229 B.n72 71.676
R803 B.n233 B.n73 71.676
R804 B.n237 B.n74 71.676
R805 B.n241 B.n75 71.676
R806 B.n245 B.n76 71.676
R807 B.n250 B.n77 71.676
R808 B.n254 B.n78 71.676
R809 B.n258 B.n79 71.676
R810 B.n262 B.n80 71.676
R811 B.n266 B.n81 71.676
R812 B.n270 B.n82 71.676
R813 B.n274 B.n83 71.676
R814 B.n278 B.n84 71.676
R815 B.n282 B.n85 71.676
R816 B.n286 B.n86 71.676
R817 B.n290 B.n87 71.676
R818 B.n294 B.n88 71.676
R819 B.n298 B.n89 71.676
R820 B.n302 B.n90 71.676
R821 B.n306 B.n91 71.676
R822 B.n310 B.n92 71.676
R823 B.n314 B.n93 71.676
R824 B.n318 B.n94 71.676
R825 B.n322 B.n95 71.676
R826 B.n326 B.n96 71.676
R827 B.n330 B.n97 71.676
R828 B.n334 B.n98 71.676
R829 B.n338 B.n99 71.676
R830 B.n342 B.n100 71.676
R831 B.n346 B.n101 71.676
R832 B.n350 B.n102 71.676
R833 B.n354 B.n103 71.676
R834 B.n358 B.n104 71.676
R835 B.n816 B.n105 71.676
R836 B.n816 B.n815 71.676
R837 B.n360 B.n104 71.676
R838 B.n357 B.n103 71.676
R839 B.n353 B.n102 71.676
R840 B.n349 B.n101 71.676
R841 B.n345 B.n100 71.676
R842 B.n341 B.n99 71.676
R843 B.n337 B.n98 71.676
R844 B.n333 B.n97 71.676
R845 B.n329 B.n96 71.676
R846 B.n325 B.n95 71.676
R847 B.n321 B.n94 71.676
R848 B.n317 B.n93 71.676
R849 B.n313 B.n92 71.676
R850 B.n309 B.n91 71.676
R851 B.n305 B.n90 71.676
R852 B.n301 B.n89 71.676
R853 B.n297 B.n88 71.676
R854 B.n293 B.n87 71.676
R855 B.n289 B.n86 71.676
R856 B.n285 B.n85 71.676
R857 B.n281 B.n84 71.676
R858 B.n277 B.n83 71.676
R859 B.n273 B.n82 71.676
R860 B.n269 B.n81 71.676
R861 B.n265 B.n80 71.676
R862 B.n261 B.n79 71.676
R863 B.n257 B.n78 71.676
R864 B.n253 B.n77 71.676
R865 B.n249 B.n76 71.676
R866 B.n244 B.n75 71.676
R867 B.n240 B.n74 71.676
R868 B.n236 B.n73 71.676
R869 B.n232 B.n72 71.676
R870 B.n228 B.n71 71.676
R871 B.n223 B.n70 71.676
R872 B.n219 B.n69 71.676
R873 B.n215 B.n68 71.676
R874 B.n211 B.n67 71.676
R875 B.n207 B.n66 71.676
R876 B.n203 B.n65 71.676
R877 B.n199 B.n64 71.676
R878 B.n195 B.n63 71.676
R879 B.n191 B.n62 71.676
R880 B.n187 B.n61 71.676
R881 B.n183 B.n60 71.676
R882 B.n179 B.n59 71.676
R883 B.n175 B.n58 71.676
R884 B.n171 B.n57 71.676
R885 B.n167 B.n56 71.676
R886 B.n163 B.n55 71.676
R887 B.n159 B.n54 71.676
R888 B.n155 B.n53 71.676
R889 B.n151 B.n52 71.676
R890 B.n147 B.n51 71.676
R891 B.n143 B.n50 71.676
R892 B.n139 B.n49 71.676
R893 B.n135 B.n48 71.676
R894 B.n131 B.n47 71.676
R895 B.n127 B.n46 71.676
R896 B.n123 B.n45 71.676
R897 B.n119 B.n44 71.676
R898 B.n115 B.n43 71.676
R899 B.n111 B.n42 71.676
R900 B.n471 B.n400 71.676
R901 B.n477 B.n476 71.676
R902 B.n480 B.n479 71.676
R903 B.n485 B.n484 71.676
R904 B.n488 B.n487 71.676
R905 B.n493 B.n492 71.676
R906 B.n496 B.n495 71.676
R907 B.n501 B.n500 71.676
R908 B.n504 B.n503 71.676
R909 B.n509 B.n508 71.676
R910 B.n512 B.n511 71.676
R911 B.n517 B.n516 71.676
R912 B.n520 B.n519 71.676
R913 B.n525 B.n524 71.676
R914 B.n528 B.n527 71.676
R915 B.n533 B.n532 71.676
R916 B.n536 B.n535 71.676
R917 B.n541 B.n540 71.676
R918 B.n544 B.n543 71.676
R919 B.n549 B.n548 71.676
R920 B.n552 B.n551 71.676
R921 B.n557 B.n556 71.676
R922 B.n560 B.n559 71.676
R923 B.n565 B.n564 71.676
R924 B.n568 B.n567 71.676
R925 B.n573 B.n572 71.676
R926 B.n576 B.n575 71.676
R927 B.n581 B.n580 71.676
R928 B.n584 B.n583 71.676
R929 B.n590 B.n589 71.676
R930 B.n593 B.n592 71.676
R931 B.n598 B.n597 71.676
R932 B.n601 B.n600 71.676
R933 B.n606 B.n605 71.676
R934 B.n609 B.n608 71.676
R935 B.n614 B.n613 71.676
R936 B.n617 B.n616 71.676
R937 B.n622 B.n621 71.676
R938 B.n625 B.n624 71.676
R939 B.n630 B.n629 71.676
R940 B.n633 B.n632 71.676
R941 B.n638 B.n637 71.676
R942 B.n641 B.n640 71.676
R943 B.n646 B.n645 71.676
R944 B.n649 B.n648 71.676
R945 B.n654 B.n653 71.676
R946 B.n657 B.n656 71.676
R947 B.n662 B.n661 71.676
R948 B.n665 B.n664 71.676
R949 B.n670 B.n669 71.676
R950 B.n673 B.n672 71.676
R951 B.n678 B.n677 71.676
R952 B.n681 B.n680 71.676
R953 B.n686 B.n685 71.676
R954 B.n689 B.n688 71.676
R955 B.n694 B.n693 71.676
R956 B.n697 B.n696 71.676
R957 B.n702 B.n701 71.676
R958 B.n705 B.n704 71.676
R959 B.n710 B.n709 71.676
R960 B.n713 B.n712 71.676
R961 B.n718 B.n717 71.676
R962 B.n721 B.n720 71.676
R963 B.n472 B.n471 71.676
R964 B.n478 B.n477 71.676
R965 B.n479 B.n468 71.676
R966 B.n486 B.n485 71.676
R967 B.n487 B.n466 71.676
R968 B.n494 B.n493 71.676
R969 B.n495 B.n464 71.676
R970 B.n502 B.n501 71.676
R971 B.n503 B.n462 71.676
R972 B.n510 B.n509 71.676
R973 B.n511 B.n460 71.676
R974 B.n518 B.n517 71.676
R975 B.n519 B.n458 71.676
R976 B.n526 B.n525 71.676
R977 B.n527 B.n456 71.676
R978 B.n534 B.n533 71.676
R979 B.n535 B.n454 71.676
R980 B.n542 B.n541 71.676
R981 B.n543 B.n452 71.676
R982 B.n550 B.n549 71.676
R983 B.n551 B.n450 71.676
R984 B.n558 B.n557 71.676
R985 B.n559 B.n448 71.676
R986 B.n566 B.n565 71.676
R987 B.n567 B.n446 71.676
R988 B.n574 B.n573 71.676
R989 B.n575 B.n444 71.676
R990 B.n582 B.n581 71.676
R991 B.n583 B.n440 71.676
R992 B.n591 B.n590 71.676
R993 B.n592 B.n438 71.676
R994 B.n599 B.n598 71.676
R995 B.n600 B.n436 71.676
R996 B.n607 B.n606 71.676
R997 B.n608 B.n431 71.676
R998 B.n615 B.n614 71.676
R999 B.n616 B.n429 71.676
R1000 B.n623 B.n622 71.676
R1001 B.n624 B.n427 71.676
R1002 B.n631 B.n630 71.676
R1003 B.n632 B.n425 71.676
R1004 B.n639 B.n638 71.676
R1005 B.n640 B.n423 71.676
R1006 B.n647 B.n646 71.676
R1007 B.n648 B.n421 71.676
R1008 B.n655 B.n654 71.676
R1009 B.n656 B.n419 71.676
R1010 B.n663 B.n662 71.676
R1011 B.n664 B.n417 71.676
R1012 B.n671 B.n670 71.676
R1013 B.n672 B.n415 71.676
R1014 B.n679 B.n678 71.676
R1015 B.n680 B.n413 71.676
R1016 B.n687 B.n686 71.676
R1017 B.n688 B.n411 71.676
R1018 B.n695 B.n694 71.676
R1019 B.n696 B.n409 71.676
R1020 B.n703 B.n702 71.676
R1021 B.n704 B.n407 71.676
R1022 B.n711 B.n710 71.676
R1023 B.n712 B.n405 71.676
R1024 B.n719 B.n718 71.676
R1025 B.n722 B.n721 71.676
R1026 B.n861 B.n860 71.676
R1027 B.n861 B.n2 71.676
R1028 B.n107 B.t5 71.5212
R1029 B.n433 B.t14 71.5212
R1030 B.n109 B.t12 71.4975
R1031 B.n442 B.t8 71.4975
R1032 B.n727 B.n401 63.1289
R1033 B.n818 B.n817 63.1289
R1034 B.n226 B.n109 59.5399
R1035 B.n247 B.n107 59.5399
R1036 B.n434 B.n433 59.5399
R1037 B.n587 B.n442 59.5399
R1038 B.n109 B.n108 41.3096
R1039 B.n107 B.n106 41.3096
R1040 B.n433 B.n432 41.3096
R1041 B.n442 B.n441 41.3096
R1042 B.n727 B.n397 32.2767
R1043 B.n733 B.n397 32.2767
R1044 B.n733 B.n393 32.2767
R1045 B.n739 B.n393 32.2767
R1046 B.n739 B.n389 32.2767
R1047 B.n745 B.n389 32.2767
R1048 B.n751 B.n385 32.2767
R1049 B.n751 B.n381 32.2767
R1050 B.n757 B.n381 32.2767
R1051 B.n757 B.n377 32.2767
R1052 B.n763 B.n377 32.2767
R1053 B.n763 B.n372 32.2767
R1054 B.n769 B.n372 32.2767
R1055 B.n769 B.n373 32.2767
R1056 B.n776 B.n365 32.2767
R1057 B.n782 B.n365 32.2767
R1058 B.n782 B.n4 32.2767
R1059 B.n859 B.n4 32.2767
R1060 B.n859 B.n858 32.2767
R1061 B.n858 B.n857 32.2767
R1062 B.n857 B.n8 32.2767
R1063 B.n12 B.n8 32.2767
R1064 B.n850 B.n12 32.2767
R1065 B.n849 B.n848 32.2767
R1066 B.n848 B.n16 32.2767
R1067 B.n842 B.n16 32.2767
R1068 B.n842 B.n841 32.2767
R1069 B.n841 B.n840 32.2767
R1070 B.n840 B.n23 32.2767
R1071 B.n834 B.n23 32.2767
R1072 B.n834 B.n833 32.2767
R1073 B.n832 B.n30 32.2767
R1074 B.n826 B.n30 32.2767
R1075 B.n826 B.n825 32.2767
R1076 B.n825 B.n824 32.2767
R1077 B.n824 B.n37 32.2767
R1078 B.n818 B.n37 32.2767
R1079 B.n729 B.n399 31.3761
R1080 B.n725 B.n724 31.3761
R1081 B.n814 B.n813 31.3761
R1082 B.n820 B.n39 31.3761
R1083 B.n373 B.t1 24.6823
R1084 B.t0 B.n849 24.6823
R1085 B.t7 B.n385 22.7837
R1086 B.n833 B.t3 22.7837
R1087 B B.n862 18.0485
R1088 B.n730 B.n729 10.6151
R1089 B.n731 B.n730 10.6151
R1090 B.n731 B.n391 10.6151
R1091 B.n741 B.n391 10.6151
R1092 B.n742 B.n741 10.6151
R1093 B.n743 B.n742 10.6151
R1094 B.n743 B.n383 10.6151
R1095 B.n753 B.n383 10.6151
R1096 B.n754 B.n753 10.6151
R1097 B.n755 B.n754 10.6151
R1098 B.n755 B.n375 10.6151
R1099 B.n765 B.n375 10.6151
R1100 B.n766 B.n765 10.6151
R1101 B.n767 B.n766 10.6151
R1102 B.n767 B.n367 10.6151
R1103 B.n778 B.n367 10.6151
R1104 B.n779 B.n778 10.6151
R1105 B.n780 B.n779 10.6151
R1106 B.n780 B.n0 10.6151
R1107 B.n473 B.n399 10.6151
R1108 B.n474 B.n473 10.6151
R1109 B.n475 B.n474 10.6151
R1110 B.n475 B.n469 10.6151
R1111 B.n481 B.n469 10.6151
R1112 B.n482 B.n481 10.6151
R1113 B.n483 B.n482 10.6151
R1114 B.n483 B.n467 10.6151
R1115 B.n489 B.n467 10.6151
R1116 B.n490 B.n489 10.6151
R1117 B.n491 B.n490 10.6151
R1118 B.n491 B.n465 10.6151
R1119 B.n497 B.n465 10.6151
R1120 B.n498 B.n497 10.6151
R1121 B.n499 B.n498 10.6151
R1122 B.n499 B.n463 10.6151
R1123 B.n505 B.n463 10.6151
R1124 B.n506 B.n505 10.6151
R1125 B.n507 B.n506 10.6151
R1126 B.n507 B.n461 10.6151
R1127 B.n513 B.n461 10.6151
R1128 B.n514 B.n513 10.6151
R1129 B.n515 B.n514 10.6151
R1130 B.n515 B.n459 10.6151
R1131 B.n521 B.n459 10.6151
R1132 B.n522 B.n521 10.6151
R1133 B.n523 B.n522 10.6151
R1134 B.n523 B.n457 10.6151
R1135 B.n529 B.n457 10.6151
R1136 B.n530 B.n529 10.6151
R1137 B.n531 B.n530 10.6151
R1138 B.n531 B.n455 10.6151
R1139 B.n537 B.n455 10.6151
R1140 B.n538 B.n537 10.6151
R1141 B.n539 B.n538 10.6151
R1142 B.n539 B.n453 10.6151
R1143 B.n545 B.n453 10.6151
R1144 B.n546 B.n545 10.6151
R1145 B.n547 B.n546 10.6151
R1146 B.n547 B.n451 10.6151
R1147 B.n553 B.n451 10.6151
R1148 B.n554 B.n553 10.6151
R1149 B.n555 B.n554 10.6151
R1150 B.n555 B.n449 10.6151
R1151 B.n561 B.n449 10.6151
R1152 B.n562 B.n561 10.6151
R1153 B.n563 B.n562 10.6151
R1154 B.n563 B.n447 10.6151
R1155 B.n569 B.n447 10.6151
R1156 B.n570 B.n569 10.6151
R1157 B.n571 B.n570 10.6151
R1158 B.n571 B.n445 10.6151
R1159 B.n577 B.n445 10.6151
R1160 B.n578 B.n577 10.6151
R1161 B.n579 B.n578 10.6151
R1162 B.n579 B.n443 10.6151
R1163 B.n585 B.n443 10.6151
R1164 B.n586 B.n585 10.6151
R1165 B.n588 B.n439 10.6151
R1166 B.n594 B.n439 10.6151
R1167 B.n595 B.n594 10.6151
R1168 B.n596 B.n595 10.6151
R1169 B.n596 B.n437 10.6151
R1170 B.n602 B.n437 10.6151
R1171 B.n603 B.n602 10.6151
R1172 B.n604 B.n603 10.6151
R1173 B.n604 B.n435 10.6151
R1174 B.n611 B.n610 10.6151
R1175 B.n612 B.n611 10.6151
R1176 B.n612 B.n430 10.6151
R1177 B.n618 B.n430 10.6151
R1178 B.n619 B.n618 10.6151
R1179 B.n620 B.n619 10.6151
R1180 B.n620 B.n428 10.6151
R1181 B.n626 B.n428 10.6151
R1182 B.n627 B.n626 10.6151
R1183 B.n628 B.n627 10.6151
R1184 B.n628 B.n426 10.6151
R1185 B.n634 B.n426 10.6151
R1186 B.n635 B.n634 10.6151
R1187 B.n636 B.n635 10.6151
R1188 B.n636 B.n424 10.6151
R1189 B.n642 B.n424 10.6151
R1190 B.n643 B.n642 10.6151
R1191 B.n644 B.n643 10.6151
R1192 B.n644 B.n422 10.6151
R1193 B.n650 B.n422 10.6151
R1194 B.n651 B.n650 10.6151
R1195 B.n652 B.n651 10.6151
R1196 B.n652 B.n420 10.6151
R1197 B.n658 B.n420 10.6151
R1198 B.n659 B.n658 10.6151
R1199 B.n660 B.n659 10.6151
R1200 B.n660 B.n418 10.6151
R1201 B.n666 B.n418 10.6151
R1202 B.n667 B.n666 10.6151
R1203 B.n668 B.n667 10.6151
R1204 B.n668 B.n416 10.6151
R1205 B.n674 B.n416 10.6151
R1206 B.n675 B.n674 10.6151
R1207 B.n676 B.n675 10.6151
R1208 B.n676 B.n414 10.6151
R1209 B.n682 B.n414 10.6151
R1210 B.n683 B.n682 10.6151
R1211 B.n684 B.n683 10.6151
R1212 B.n684 B.n412 10.6151
R1213 B.n690 B.n412 10.6151
R1214 B.n691 B.n690 10.6151
R1215 B.n692 B.n691 10.6151
R1216 B.n692 B.n410 10.6151
R1217 B.n698 B.n410 10.6151
R1218 B.n699 B.n698 10.6151
R1219 B.n700 B.n699 10.6151
R1220 B.n700 B.n408 10.6151
R1221 B.n706 B.n408 10.6151
R1222 B.n707 B.n706 10.6151
R1223 B.n708 B.n707 10.6151
R1224 B.n708 B.n406 10.6151
R1225 B.n714 B.n406 10.6151
R1226 B.n715 B.n714 10.6151
R1227 B.n716 B.n715 10.6151
R1228 B.n716 B.n404 10.6151
R1229 B.n404 B.n403 10.6151
R1230 B.n723 B.n403 10.6151
R1231 B.n724 B.n723 10.6151
R1232 B.n725 B.n395 10.6151
R1233 B.n735 B.n395 10.6151
R1234 B.n736 B.n735 10.6151
R1235 B.n737 B.n736 10.6151
R1236 B.n737 B.n387 10.6151
R1237 B.n747 B.n387 10.6151
R1238 B.n748 B.n747 10.6151
R1239 B.n749 B.n748 10.6151
R1240 B.n749 B.n379 10.6151
R1241 B.n759 B.n379 10.6151
R1242 B.n760 B.n759 10.6151
R1243 B.n761 B.n760 10.6151
R1244 B.n761 B.n370 10.6151
R1245 B.n771 B.n370 10.6151
R1246 B.n772 B.n771 10.6151
R1247 B.n774 B.n772 10.6151
R1248 B.n774 B.n773 10.6151
R1249 B.n773 B.n363 10.6151
R1250 B.n785 B.n363 10.6151
R1251 B.n786 B.n785 10.6151
R1252 B.n787 B.n786 10.6151
R1253 B.n788 B.n787 10.6151
R1254 B.n789 B.n788 10.6151
R1255 B.n792 B.n789 10.6151
R1256 B.n793 B.n792 10.6151
R1257 B.n794 B.n793 10.6151
R1258 B.n795 B.n794 10.6151
R1259 B.n797 B.n795 10.6151
R1260 B.n798 B.n797 10.6151
R1261 B.n799 B.n798 10.6151
R1262 B.n800 B.n799 10.6151
R1263 B.n802 B.n800 10.6151
R1264 B.n803 B.n802 10.6151
R1265 B.n804 B.n803 10.6151
R1266 B.n805 B.n804 10.6151
R1267 B.n807 B.n805 10.6151
R1268 B.n808 B.n807 10.6151
R1269 B.n809 B.n808 10.6151
R1270 B.n810 B.n809 10.6151
R1271 B.n812 B.n810 10.6151
R1272 B.n813 B.n812 10.6151
R1273 B.n854 B.n1 10.6151
R1274 B.n854 B.n853 10.6151
R1275 B.n853 B.n852 10.6151
R1276 B.n852 B.n10 10.6151
R1277 B.n846 B.n10 10.6151
R1278 B.n846 B.n845 10.6151
R1279 B.n845 B.n844 10.6151
R1280 B.n844 B.n18 10.6151
R1281 B.n838 B.n18 10.6151
R1282 B.n838 B.n837 10.6151
R1283 B.n837 B.n836 10.6151
R1284 B.n836 B.n25 10.6151
R1285 B.n830 B.n25 10.6151
R1286 B.n830 B.n829 10.6151
R1287 B.n829 B.n828 10.6151
R1288 B.n828 B.n32 10.6151
R1289 B.n822 B.n32 10.6151
R1290 B.n822 B.n821 10.6151
R1291 B.n821 B.n820 10.6151
R1292 B.n110 B.n39 10.6151
R1293 B.n113 B.n110 10.6151
R1294 B.n114 B.n113 10.6151
R1295 B.n117 B.n114 10.6151
R1296 B.n118 B.n117 10.6151
R1297 B.n121 B.n118 10.6151
R1298 B.n122 B.n121 10.6151
R1299 B.n125 B.n122 10.6151
R1300 B.n126 B.n125 10.6151
R1301 B.n129 B.n126 10.6151
R1302 B.n130 B.n129 10.6151
R1303 B.n133 B.n130 10.6151
R1304 B.n134 B.n133 10.6151
R1305 B.n137 B.n134 10.6151
R1306 B.n138 B.n137 10.6151
R1307 B.n141 B.n138 10.6151
R1308 B.n142 B.n141 10.6151
R1309 B.n145 B.n142 10.6151
R1310 B.n146 B.n145 10.6151
R1311 B.n149 B.n146 10.6151
R1312 B.n150 B.n149 10.6151
R1313 B.n153 B.n150 10.6151
R1314 B.n154 B.n153 10.6151
R1315 B.n157 B.n154 10.6151
R1316 B.n158 B.n157 10.6151
R1317 B.n161 B.n158 10.6151
R1318 B.n162 B.n161 10.6151
R1319 B.n165 B.n162 10.6151
R1320 B.n166 B.n165 10.6151
R1321 B.n169 B.n166 10.6151
R1322 B.n170 B.n169 10.6151
R1323 B.n173 B.n170 10.6151
R1324 B.n174 B.n173 10.6151
R1325 B.n177 B.n174 10.6151
R1326 B.n178 B.n177 10.6151
R1327 B.n181 B.n178 10.6151
R1328 B.n182 B.n181 10.6151
R1329 B.n185 B.n182 10.6151
R1330 B.n186 B.n185 10.6151
R1331 B.n189 B.n186 10.6151
R1332 B.n190 B.n189 10.6151
R1333 B.n193 B.n190 10.6151
R1334 B.n194 B.n193 10.6151
R1335 B.n197 B.n194 10.6151
R1336 B.n198 B.n197 10.6151
R1337 B.n201 B.n198 10.6151
R1338 B.n202 B.n201 10.6151
R1339 B.n205 B.n202 10.6151
R1340 B.n206 B.n205 10.6151
R1341 B.n209 B.n206 10.6151
R1342 B.n210 B.n209 10.6151
R1343 B.n213 B.n210 10.6151
R1344 B.n214 B.n213 10.6151
R1345 B.n217 B.n214 10.6151
R1346 B.n218 B.n217 10.6151
R1347 B.n221 B.n218 10.6151
R1348 B.n222 B.n221 10.6151
R1349 B.n225 B.n222 10.6151
R1350 B.n230 B.n227 10.6151
R1351 B.n231 B.n230 10.6151
R1352 B.n234 B.n231 10.6151
R1353 B.n235 B.n234 10.6151
R1354 B.n238 B.n235 10.6151
R1355 B.n239 B.n238 10.6151
R1356 B.n242 B.n239 10.6151
R1357 B.n243 B.n242 10.6151
R1358 B.n246 B.n243 10.6151
R1359 B.n251 B.n248 10.6151
R1360 B.n252 B.n251 10.6151
R1361 B.n255 B.n252 10.6151
R1362 B.n256 B.n255 10.6151
R1363 B.n259 B.n256 10.6151
R1364 B.n260 B.n259 10.6151
R1365 B.n263 B.n260 10.6151
R1366 B.n264 B.n263 10.6151
R1367 B.n267 B.n264 10.6151
R1368 B.n268 B.n267 10.6151
R1369 B.n271 B.n268 10.6151
R1370 B.n272 B.n271 10.6151
R1371 B.n275 B.n272 10.6151
R1372 B.n276 B.n275 10.6151
R1373 B.n279 B.n276 10.6151
R1374 B.n280 B.n279 10.6151
R1375 B.n283 B.n280 10.6151
R1376 B.n284 B.n283 10.6151
R1377 B.n287 B.n284 10.6151
R1378 B.n288 B.n287 10.6151
R1379 B.n291 B.n288 10.6151
R1380 B.n292 B.n291 10.6151
R1381 B.n295 B.n292 10.6151
R1382 B.n296 B.n295 10.6151
R1383 B.n299 B.n296 10.6151
R1384 B.n300 B.n299 10.6151
R1385 B.n303 B.n300 10.6151
R1386 B.n304 B.n303 10.6151
R1387 B.n307 B.n304 10.6151
R1388 B.n308 B.n307 10.6151
R1389 B.n311 B.n308 10.6151
R1390 B.n312 B.n311 10.6151
R1391 B.n315 B.n312 10.6151
R1392 B.n316 B.n315 10.6151
R1393 B.n319 B.n316 10.6151
R1394 B.n320 B.n319 10.6151
R1395 B.n323 B.n320 10.6151
R1396 B.n324 B.n323 10.6151
R1397 B.n327 B.n324 10.6151
R1398 B.n328 B.n327 10.6151
R1399 B.n331 B.n328 10.6151
R1400 B.n332 B.n331 10.6151
R1401 B.n335 B.n332 10.6151
R1402 B.n336 B.n335 10.6151
R1403 B.n339 B.n336 10.6151
R1404 B.n340 B.n339 10.6151
R1405 B.n343 B.n340 10.6151
R1406 B.n344 B.n343 10.6151
R1407 B.n347 B.n344 10.6151
R1408 B.n348 B.n347 10.6151
R1409 B.n351 B.n348 10.6151
R1410 B.n352 B.n351 10.6151
R1411 B.n355 B.n352 10.6151
R1412 B.n356 B.n355 10.6151
R1413 B.n359 B.n356 10.6151
R1414 B.n361 B.n359 10.6151
R1415 B.n362 B.n361 10.6151
R1416 B.n814 B.n362 10.6151
R1417 B.n745 B.t7 9.49349
R1418 B.t3 B.n832 9.49349
R1419 B.n587 B.n586 9.36635
R1420 B.n610 B.n434 9.36635
R1421 B.n226 B.n225 9.36635
R1422 B.n248 B.n247 9.36635
R1423 B.n862 B.n0 8.11757
R1424 B.n862 B.n1 8.11757
R1425 B.n776 B.t1 7.59489
R1426 B.n850 B.t0 7.59489
R1427 B.n588 B.n587 1.24928
R1428 B.n435 B.n434 1.24928
R1429 B.n227 B.n226 1.24928
R1430 B.n247 B.n246 1.24928
R1431 VP.n0 VP.t0 345.551
R1432 VP.n0 VP.t1 298.548
R1433 VP VP.n0 0.241678
R1434 VTAIL.n1 VTAIL.t1 45.4792
R1435 VTAIL.n3 VTAIL.t0 45.479
R1436 VTAIL.n0 VTAIL.t2 45.479
R1437 VTAIL.n2 VTAIL.t3 45.479
R1438 VTAIL.n1 VTAIL.n0 31.4703
R1439 VTAIL.n3 VTAIL.n2 29.6341
R1440 VTAIL.n2 VTAIL.n1 1.38843
R1441 VTAIL VTAIL.n0 0.987569
R1442 VTAIL VTAIL.n3 0.401362
R1443 VDD1 VDD1.t0 105.904
R1444 VDD1 VDD1.t1 62.675
R1445 VN VN.t0 345.743
R1446 VN VN.t1 298.788
R1447 VDD2.n0 VDD2.t0 104.921
R1448 VDD2.n0 VDD2.t1 62.1578
R1449 VDD2 VDD2.n0 0.517741
C0 VDD2 VDD1 0.581157f
C1 VDD1 VP 3.90996f
C2 VTAIL VN 3.11333f
C3 VDD2 VN 3.76197f
C4 VN VP 6.17117f
C5 VTAIL VDD2 6.74405f
C6 VTAIL VP 3.12783f
C7 VN VDD1 0.148089f
C8 VDD2 VP 0.300472f
C9 VTAIL VDD1 6.7018f
C10 VDD2 B 5.210653f
C11 VDD1 B 8.61442f
C12 VTAIL B 9.294222f
C13 VN B 11.485519f
C14 VP B 5.807191f
C15 VDD2.t0 B 3.94692f
C16 VDD2.t1 B 3.28277f
C17 VDD2.n0 B 3.17757f
C18 VN.t1 B 3.53393f
C19 VN.t0 B 3.94162f
C20 VDD1.t1 B 3.29312f
C21 VDD1.t0 B 3.99089f
C22 VTAIL.t2 B 3.13742f
C23 VTAIL.n0 B 1.79512f
C24 VTAIL.t1 B 3.13742f
C25 VTAIL.n1 B 1.82033f
C26 VTAIL.t3 B 3.13742f
C27 VTAIL.n2 B 1.70483f
C28 VTAIL.t0 B 3.13742f
C29 VTAIL.n3 B 1.64275f
C30 VP.t0 B 3.98378f
C31 VP.t1 B 3.57412f
C32 VP.n0 B 5.58528f
.ends

