* NGSPICE file created from diff_pair_sample_1532.ext - technology: sky130A

.subckt diff_pair_sample_1532 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=3.3618 ps=18.02 w=8.62 l=3.2
X1 VTAIL.t14 VP.t1 VDD1.t8 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X2 VDD1.t7 VP.t2 VTAIL.t11 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X3 VTAIL.t6 VN.t0 VDD2.t9 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X4 VDD2.t8 VN.t1 VTAIL.t4 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=1.4223 ps=8.95 w=8.62 l=3.2
X5 VDD1.t6 VP.t3 VTAIL.t10 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=1.4223 ps=8.95 w=8.62 l=3.2
X6 VDD2.t7 VN.t2 VTAIL.t3 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X7 VTAIL.t12 VP.t4 VDD1.t5 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X8 B.t11 B.t9 B.t10 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=0 ps=0 w=8.62 l=3.2
X9 B.t8 B.t6 B.t7 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=0 ps=0 w=8.62 l=3.2
X10 VDD2.t6 VN.t3 VTAIL.t1 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=3.3618 ps=18.02 w=8.62 l=3.2
X11 B.t5 B.t3 B.t4 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=0 ps=0 w=8.62 l=3.2
X12 VDD1.t4 VP.t5 VTAIL.t13 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X13 VTAIL.t15 VP.t6 VDD1.t3 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X14 VDD2.t5 VN.t4 VTAIL.t0 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=3.3618 ps=18.02 w=8.62 l=3.2
X15 VTAIL.t2 VN.t5 VDD2.t4 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X16 VDD2.t3 VN.t6 VTAIL.t5 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X17 VDD2.t2 VN.t7 VTAIL.t9 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=1.4223 ps=8.95 w=8.62 l=3.2
X18 VDD1.t2 VP.t7 VTAIL.t19 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=1.4223 ps=8.95 w=8.62 l=3.2
X19 VTAIL.t18 VP.t8 VDD1.t1 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X20 B.t2 B.t0 B.t1 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=3.3618 pd=18.02 as=0 ps=0 w=8.62 l=3.2
X21 VDD1.t0 VP.t9 VTAIL.t17 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=3.3618 ps=18.02 w=8.62 l=3.2
X22 VTAIL.t7 VN.t8 VDD2.t1 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
X23 VTAIL.t8 VN.t9 VDD2.t0 w_n5206_n2692# sky130_fd_pr__pfet_01v8 ad=1.4223 pd=8.95 as=1.4223 ps=8.95 w=8.62 l=3.2
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n109 VP.n108 161.3
R22 VP.n107 VP.n1 161.3
R23 VP.n106 VP.n105 161.3
R24 VP.n104 VP.n2 161.3
R25 VP.n103 VP.n102 161.3
R26 VP.n101 VP.n3 161.3
R27 VP.n100 VP.n99 161.3
R28 VP.n98 VP.n97 161.3
R29 VP.n96 VP.n5 161.3
R30 VP.n95 VP.n94 161.3
R31 VP.n93 VP.n6 161.3
R32 VP.n92 VP.n91 161.3
R33 VP.n90 VP.n7 161.3
R34 VP.n89 VP.n88 161.3
R35 VP.n87 VP.n86 161.3
R36 VP.n85 VP.n9 161.3
R37 VP.n84 VP.n83 161.3
R38 VP.n82 VP.n10 161.3
R39 VP.n81 VP.n80 161.3
R40 VP.n79 VP.n11 161.3
R41 VP.n78 VP.n77 161.3
R42 VP.n76 VP.n75 161.3
R43 VP.n74 VP.n13 161.3
R44 VP.n73 VP.n72 161.3
R45 VP.n71 VP.n14 161.3
R46 VP.n70 VP.n69 161.3
R47 VP.n68 VP.n15 161.3
R48 VP.n67 VP.n66 161.3
R49 VP.n30 VP.t7 98.0241
R50 VP.n65 VP.n16 74.9986
R51 VP.n110 VP.n0 74.9986
R52 VP.n64 VP.n17 74.9986
R53 VP.n16 VP.t3 64.9199
R54 VP.n12 VP.t8 64.9199
R55 VP.n8 VP.t5 64.9199
R56 VP.n4 VP.t4 64.9199
R57 VP.n0 VP.t9 64.9199
R58 VP.n17 VP.t0 64.9199
R59 VP.n21 VP.t1 64.9199
R60 VP.n25 VP.t2 64.9199
R61 VP.n29 VP.t6 64.9199
R62 VP.n30 VP.n29 60.6744
R63 VP.n65 VP.n64 53.9124
R64 VP.n69 VP.n14 44.9365
R65 VP.n106 VP.n2 44.9365
R66 VP.n60 VP.n19 44.9365
R67 VP.n80 VP.n10 42.0302
R68 VP.n95 VP.n6 42.0302
R69 VP.n49 VP.n23 42.0302
R70 VP.n34 VP.n27 42.0302
R71 VP.n84 VP.n10 39.1239
R72 VP.n91 VP.n6 39.1239
R73 VP.n45 VP.n23 39.1239
R74 VP.n38 VP.n27 39.1239
R75 VP.n73 VP.n14 36.2176
R76 VP.n102 VP.n2 36.2176
R77 VP.n56 VP.n19 36.2176
R78 VP.n68 VP.n67 24.5923
R79 VP.n69 VP.n68 24.5923
R80 VP.n74 VP.n73 24.5923
R81 VP.n75 VP.n74 24.5923
R82 VP.n79 VP.n78 24.5923
R83 VP.n80 VP.n79 24.5923
R84 VP.n85 VP.n84 24.5923
R85 VP.n86 VP.n85 24.5923
R86 VP.n90 VP.n89 24.5923
R87 VP.n91 VP.n90 24.5923
R88 VP.n96 VP.n95 24.5923
R89 VP.n97 VP.n96 24.5923
R90 VP.n101 VP.n100 24.5923
R91 VP.n102 VP.n101 24.5923
R92 VP.n107 VP.n106 24.5923
R93 VP.n108 VP.n107 24.5923
R94 VP.n61 VP.n60 24.5923
R95 VP.n62 VP.n61 24.5923
R96 VP.n50 VP.n49 24.5923
R97 VP.n51 VP.n50 24.5923
R98 VP.n55 VP.n54 24.5923
R99 VP.n56 VP.n55 24.5923
R100 VP.n39 VP.n38 24.5923
R101 VP.n40 VP.n39 24.5923
R102 VP.n44 VP.n43 24.5923
R103 VP.n45 VP.n44 24.5923
R104 VP.n33 VP.n32 24.5923
R105 VP.n34 VP.n33 24.5923
R106 VP.n67 VP.n16 15.2474
R107 VP.n108 VP.n0 15.2474
R108 VP.n62 VP.n17 15.2474
R109 VP.n78 VP.n12 13.7719
R110 VP.n97 VP.n4 13.7719
R111 VP.n51 VP.n21 13.7719
R112 VP.n32 VP.n29 13.7719
R113 VP.n86 VP.n8 12.2964
R114 VP.n89 VP.n8 12.2964
R115 VP.n40 VP.n25 12.2964
R116 VP.n43 VP.n25 12.2964
R117 VP.n75 VP.n12 10.8209
R118 VP.n100 VP.n4 10.8209
R119 VP.n54 VP.n21 10.8209
R120 VP.n31 VP.n30 4.12004
R121 VP.n64 VP.n63 0.354861
R122 VP.n66 VP.n65 0.354861
R123 VP.n110 VP.n109 0.354861
R124 VP VP.n110 0.267071
R125 VP.n31 VP.n28 0.189894
R126 VP.n35 VP.n28 0.189894
R127 VP.n36 VP.n35 0.189894
R128 VP.n37 VP.n36 0.189894
R129 VP.n37 VP.n26 0.189894
R130 VP.n41 VP.n26 0.189894
R131 VP.n42 VP.n41 0.189894
R132 VP.n42 VP.n24 0.189894
R133 VP.n46 VP.n24 0.189894
R134 VP.n47 VP.n46 0.189894
R135 VP.n48 VP.n47 0.189894
R136 VP.n48 VP.n22 0.189894
R137 VP.n52 VP.n22 0.189894
R138 VP.n53 VP.n52 0.189894
R139 VP.n53 VP.n20 0.189894
R140 VP.n57 VP.n20 0.189894
R141 VP.n58 VP.n57 0.189894
R142 VP.n59 VP.n58 0.189894
R143 VP.n59 VP.n18 0.189894
R144 VP.n63 VP.n18 0.189894
R145 VP.n66 VP.n15 0.189894
R146 VP.n70 VP.n15 0.189894
R147 VP.n71 VP.n70 0.189894
R148 VP.n72 VP.n71 0.189894
R149 VP.n72 VP.n13 0.189894
R150 VP.n76 VP.n13 0.189894
R151 VP.n77 VP.n76 0.189894
R152 VP.n77 VP.n11 0.189894
R153 VP.n81 VP.n11 0.189894
R154 VP.n82 VP.n81 0.189894
R155 VP.n83 VP.n82 0.189894
R156 VP.n83 VP.n9 0.189894
R157 VP.n87 VP.n9 0.189894
R158 VP.n88 VP.n87 0.189894
R159 VP.n88 VP.n7 0.189894
R160 VP.n92 VP.n7 0.189894
R161 VP.n93 VP.n92 0.189894
R162 VP.n94 VP.n93 0.189894
R163 VP.n94 VP.n5 0.189894
R164 VP.n98 VP.n5 0.189894
R165 VP.n99 VP.n98 0.189894
R166 VP.n99 VP.n3 0.189894
R167 VP.n103 VP.n3 0.189894
R168 VP.n104 VP.n103 0.189894
R169 VP.n105 VP.n104 0.189894
R170 VP.n105 VP.n1 0.189894
R171 VP.n109 VP.n1 0.189894
R172 VTAIL.n192 VTAIL.n152 756.745
R173 VTAIL.n42 VTAIL.n2 756.745
R174 VTAIL.n146 VTAIL.n106 756.745
R175 VTAIL.n96 VTAIL.n56 756.745
R176 VTAIL.n167 VTAIL.n166 585
R177 VTAIL.n164 VTAIL.n163 585
R178 VTAIL.n173 VTAIL.n172 585
R179 VTAIL.n175 VTAIL.n174 585
R180 VTAIL.n160 VTAIL.n159 585
R181 VTAIL.n181 VTAIL.n180 585
R182 VTAIL.n184 VTAIL.n183 585
R183 VTAIL.n182 VTAIL.n156 585
R184 VTAIL.n189 VTAIL.n155 585
R185 VTAIL.n191 VTAIL.n190 585
R186 VTAIL.n193 VTAIL.n192 585
R187 VTAIL.n17 VTAIL.n16 585
R188 VTAIL.n14 VTAIL.n13 585
R189 VTAIL.n23 VTAIL.n22 585
R190 VTAIL.n25 VTAIL.n24 585
R191 VTAIL.n10 VTAIL.n9 585
R192 VTAIL.n31 VTAIL.n30 585
R193 VTAIL.n34 VTAIL.n33 585
R194 VTAIL.n32 VTAIL.n6 585
R195 VTAIL.n39 VTAIL.n5 585
R196 VTAIL.n41 VTAIL.n40 585
R197 VTAIL.n43 VTAIL.n42 585
R198 VTAIL.n147 VTAIL.n146 585
R199 VTAIL.n145 VTAIL.n144 585
R200 VTAIL.n143 VTAIL.n109 585
R201 VTAIL.n113 VTAIL.n110 585
R202 VTAIL.n138 VTAIL.n137 585
R203 VTAIL.n136 VTAIL.n135 585
R204 VTAIL.n115 VTAIL.n114 585
R205 VTAIL.n130 VTAIL.n129 585
R206 VTAIL.n128 VTAIL.n127 585
R207 VTAIL.n119 VTAIL.n118 585
R208 VTAIL.n122 VTAIL.n121 585
R209 VTAIL.n97 VTAIL.n96 585
R210 VTAIL.n95 VTAIL.n94 585
R211 VTAIL.n93 VTAIL.n59 585
R212 VTAIL.n63 VTAIL.n60 585
R213 VTAIL.n88 VTAIL.n87 585
R214 VTAIL.n86 VTAIL.n85 585
R215 VTAIL.n65 VTAIL.n64 585
R216 VTAIL.n80 VTAIL.n79 585
R217 VTAIL.n78 VTAIL.n77 585
R218 VTAIL.n69 VTAIL.n68 585
R219 VTAIL.n72 VTAIL.n71 585
R220 VTAIL.t16 VTAIL.n120 329.039
R221 VTAIL.t0 VTAIL.n70 329.039
R222 VTAIL.t1 VTAIL.n165 329.038
R223 VTAIL.t17 VTAIL.n15 329.038
R224 VTAIL.n166 VTAIL.n163 171.744
R225 VTAIL.n173 VTAIL.n163 171.744
R226 VTAIL.n174 VTAIL.n173 171.744
R227 VTAIL.n174 VTAIL.n159 171.744
R228 VTAIL.n181 VTAIL.n159 171.744
R229 VTAIL.n183 VTAIL.n181 171.744
R230 VTAIL.n183 VTAIL.n182 171.744
R231 VTAIL.n182 VTAIL.n155 171.744
R232 VTAIL.n191 VTAIL.n155 171.744
R233 VTAIL.n192 VTAIL.n191 171.744
R234 VTAIL.n16 VTAIL.n13 171.744
R235 VTAIL.n23 VTAIL.n13 171.744
R236 VTAIL.n24 VTAIL.n23 171.744
R237 VTAIL.n24 VTAIL.n9 171.744
R238 VTAIL.n31 VTAIL.n9 171.744
R239 VTAIL.n33 VTAIL.n31 171.744
R240 VTAIL.n33 VTAIL.n32 171.744
R241 VTAIL.n32 VTAIL.n5 171.744
R242 VTAIL.n41 VTAIL.n5 171.744
R243 VTAIL.n42 VTAIL.n41 171.744
R244 VTAIL.n146 VTAIL.n145 171.744
R245 VTAIL.n145 VTAIL.n109 171.744
R246 VTAIL.n113 VTAIL.n109 171.744
R247 VTAIL.n137 VTAIL.n113 171.744
R248 VTAIL.n137 VTAIL.n136 171.744
R249 VTAIL.n136 VTAIL.n114 171.744
R250 VTAIL.n129 VTAIL.n114 171.744
R251 VTAIL.n129 VTAIL.n128 171.744
R252 VTAIL.n128 VTAIL.n118 171.744
R253 VTAIL.n121 VTAIL.n118 171.744
R254 VTAIL.n96 VTAIL.n95 171.744
R255 VTAIL.n95 VTAIL.n59 171.744
R256 VTAIL.n63 VTAIL.n59 171.744
R257 VTAIL.n87 VTAIL.n63 171.744
R258 VTAIL.n87 VTAIL.n86 171.744
R259 VTAIL.n86 VTAIL.n64 171.744
R260 VTAIL.n79 VTAIL.n64 171.744
R261 VTAIL.n79 VTAIL.n78 171.744
R262 VTAIL.n78 VTAIL.n68 171.744
R263 VTAIL.n71 VTAIL.n68 171.744
R264 VTAIL.n166 VTAIL.t1 85.8723
R265 VTAIL.n16 VTAIL.t17 85.8723
R266 VTAIL.n121 VTAIL.t16 85.8723
R267 VTAIL.n71 VTAIL.t0 85.8723
R268 VTAIL.n105 VTAIL.n104 65.5649
R269 VTAIL.n103 VTAIL.n102 65.5649
R270 VTAIL.n55 VTAIL.n54 65.5649
R271 VTAIL.n53 VTAIL.n52 65.5649
R272 VTAIL.n199 VTAIL.n198 65.5647
R273 VTAIL.n1 VTAIL.n0 65.5647
R274 VTAIL.n49 VTAIL.n48 65.5647
R275 VTAIL.n51 VTAIL.n50 65.5647
R276 VTAIL.n197 VTAIL.n196 34.1247
R277 VTAIL.n47 VTAIL.n46 34.1247
R278 VTAIL.n151 VTAIL.n150 34.1247
R279 VTAIL.n101 VTAIL.n100 34.1247
R280 VTAIL.n53 VTAIL.n51 25.8841
R281 VTAIL.n197 VTAIL.n151 22.841
R282 VTAIL.n190 VTAIL.n189 13.1884
R283 VTAIL.n40 VTAIL.n39 13.1884
R284 VTAIL.n144 VTAIL.n143 13.1884
R285 VTAIL.n94 VTAIL.n93 13.1884
R286 VTAIL.n188 VTAIL.n156 12.8005
R287 VTAIL.n193 VTAIL.n154 12.8005
R288 VTAIL.n38 VTAIL.n6 12.8005
R289 VTAIL.n43 VTAIL.n4 12.8005
R290 VTAIL.n147 VTAIL.n108 12.8005
R291 VTAIL.n142 VTAIL.n110 12.8005
R292 VTAIL.n97 VTAIL.n58 12.8005
R293 VTAIL.n92 VTAIL.n60 12.8005
R294 VTAIL.n185 VTAIL.n184 12.0247
R295 VTAIL.n194 VTAIL.n152 12.0247
R296 VTAIL.n35 VTAIL.n34 12.0247
R297 VTAIL.n44 VTAIL.n2 12.0247
R298 VTAIL.n148 VTAIL.n106 12.0247
R299 VTAIL.n139 VTAIL.n138 12.0247
R300 VTAIL.n98 VTAIL.n56 12.0247
R301 VTAIL.n89 VTAIL.n88 12.0247
R302 VTAIL.n180 VTAIL.n158 11.249
R303 VTAIL.n30 VTAIL.n8 11.249
R304 VTAIL.n135 VTAIL.n112 11.249
R305 VTAIL.n85 VTAIL.n62 11.249
R306 VTAIL.n167 VTAIL.n165 10.7239
R307 VTAIL.n17 VTAIL.n15 10.7239
R308 VTAIL.n122 VTAIL.n120 10.7239
R309 VTAIL.n72 VTAIL.n70 10.7239
R310 VTAIL.n179 VTAIL.n160 10.4732
R311 VTAIL.n29 VTAIL.n10 10.4732
R312 VTAIL.n134 VTAIL.n115 10.4732
R313 VTAIL.n84 VTAIL.n65 10.4732
R314 VTAIL.n176 VTAIL.n175 9.69747
R315 VTAIL.n26 VTAIL.n25 9.69747
R316 VTAIL.n131 VTAIL.n130 9.69747
R317 VTAIL.n81 VTAIL.n80 9.69747
R318 VTAIL.n196 VTAIL.n195 9.45567
R319 VTAIL.n46 VTAIL.n45 9.45567
R320 VTAIL.n150 VTAIL.n149 9.45567
R321 VTAIL.n100 VTAIL.n99 9.45567
R322 VTAIL.n195 VTAIL.n194 9.3005
R323 VTAIL.n154 VTAIL.n153 9.3005
R324 VTAIL.n169 VTAIL.n168 9.3005
R325 VTAIL.n171 VTAIL.n170 9.3005
R326 VTAIL.n162 VTAIL.n161 9.3005
R327 VTAIL.n177 VTAIL.n176 9.3005
R328 VTAIL.n179 VTAIL.n178 9.3005
R329 VTAIL.n158 VTAIL.n157 9.3005
R330 VTAIL.n186 VTAIL.n185 9.3005
R331 VTAIL.n188 VTAIL.n187 9.3005
R332 VTAIL.n45 VTAIL.n44 9.3005
R333 VTAIL.n4 VTAIL.n3 9.3005
R334 VTAIL.n19 VTAIL.n18 9.3005
R335 VTAIL.n21 VTAIL.n20 9.3005
R336 VTAIL.n12 VTAIL.n11 9.3005
R337 VTAIL.n27 VTAIL.n26 9.3005
R338 VTAIL.n29 VTAIL.n28 9.3005
R339 VTAIL.n8 VTAIL.n7 9.3005
R340 VTAIL.n36 VTAIL.n35 9.3005
R341 VTAIL.n38 VTAIL.n37 9.3005
R342 VTAIL.n124 VTAIL.n123 9.3005
R343 VTAIL.n126 VTAIL.n125 9.3005
R344 VTAIL.n117 VTAIL.n116 9.3005
R345 VTAIL.n132 VTAIL.n131 9.3005
R346 VTAIL.n134 VTAIL.n133 9.3005
R347 VTAIL.n112 VTAIL.n111 9.3005
R348 VTAIL.n140 VTAIL.n139 9.3005
R349 VTAIL.n142 VTAIL.n141 9.3005
R350 VTAIL.n149 VTAIL.n148 9.3005
R351 VTAIL.n108 VTAIL.n107 9.3005
R352 VTAIL.n74 VTAIL.n73 9.3005
R353 VTAIL.n76 VTAIL.n75 9.3005
R354 VTAIL.n67 VTAIL.n66 9.3005
R355 VTAIL.n82 VTAIL.n81 9.3005
R356 VTAIL.n84 VTAIL.n83 9.3005
R357 VTAIL.n62 VTAIL.n61 9.3005
R358 VTAIL.n90 VTAIL.n89 9.3005
R359 VTAIL.n92 VTAIL.n91 9.3005
R360 VTAIL.n99 VTAIL.n98 9.3005
R361 VTAIL.n58 VTAIL.n57 9.3005
R362 VTAIL.n172 VTAIL.n162 8.92171
R363 VTAIL.n22 VTAIL.n12 8.92171
R364 VTAIL.n127 VTAIL.n117 8.92171
R365 VTAIL.n77 VTAIL.n67 8.92171
R366 VTAIL.n171 VTAIL.n164 8.14595
R367 VTAIL.n21 VTAIL.n14 8.14595
R368 VTAIL.n126 VTAIL.n119 8.14595
R369 VTAIL.n76 VTAIL.n69 8.14595
R370 VTAIL.n168 VTAIL.n167 7.3702
R371 VTAIL.n18 VTAIL.n17 7.3702
R372 VTAIL.n123 VTAIL.n122 7.3702
R373 VTAIL.n73 VTAIL.n72 7.3702
R374 VTAIL.n168 VTAIL.n164 5.81868
R375 VTAIL.n18 VTAIL.n14 5.81868
R376 VTAIL.n123 VTAIL.n119 5.81868
R377 VTAIL.n73 VTAIL.n69 5.81868
R378 VTAIL.n172 VTAIL.n171 5.04292
R379 VTAIL.n22 VTAIL.n21 5.04292
R380 VTAIL.n127 VTAIL.n126 5.04292
R381 VTAIL.n77 VTAIL.n76 5.04292
R382 VTAIL.n175 VTAIL.n162 4.26717
R383 VTAIL.n25 VTAIL.n12 4.26717
R384 VTAIL.n130 VTAIL.n117 4.26717
R385 VTAIL.n80 VTAIL.n67 4.26717
R386 VTAIL.n198 VTAIL.t3 3.77138
R387 VTAIL.n198 VTAIL.t7 3.77138
R388 VTAIL.n0 VTAIL.t9 3.77138
R389 VTAIL.n0 VTAIL.t8 3.77138
R390 VTAIL.n48 VTAIL.t13 3.77138
R391 VTAIL.n48 VTAIL.t12 3.77138
R392 VTAIL.n50 VTAIL.t10 3.77138
R393 VTAIL.n50 VTAIL.t18 3.77138
R394 VTAIL.n104 VTAIL.t11 3.77138
R395 VTAIL.n104 VTAIL.t14 3.77138
R396 VTAIL.n102 VTAIL.t19 3.77138
R397 VTAIL.n102 VTAIL.t15 3.77138
R398 VTAIL.n54 VTAIL.t5 3.77138
R399 VTAIL.n54 VTAIL.t2 3.77138
R400 VTAIL.n52 VTAIL.t4 3.77138
R401 VTAIL.n52 VTAIL.t6 3.77138
R402 VTAIL.n176 VTAIL.n160 3.49141
R403 VTAIL.n26 VTAIL.n10 3.49141
R404 VTAIL.n131 VTAIL.n115 3.49141
R405 VTAIL.n81 VTAIL.n65 3.49141
R406 VTAIL.n55 VTAIL.n53 3.0436
R407 VTAIL.n101 VTAIL.n55 3.0436
R408 VTAIL.n105 VTAIL.n103 3.0436
R409 VTAIL.n151 VTAIL.n105 3.0436
R410 VTAIL.n51 VTAIL.n49 3.0436
R411 VTAIL.n49 VTAIL.n47 3.0436
R412 VTAIL.n199 VTAIL.n197 3.0436
R413 VTAIL.n180 VTAIL.n179 2.71565
R414 VTAIL.n30 VTAIL.n29 2.71565
R415 VTAIL.n135 VTAIL.n134 2.71565
R416 VTAIL.n85 VTAIL.n84 2.71565
R417 VTAIL.n169 VTAIL.n165 2.41285
R418 VTAIL.n19 VTAIL.n15 2.41285
R419 VTAIL.n124 VTAIL.n120 2.41285
R420 VTAIL.n74 VTAIL.n70 2.41285
R421 VTAIL VTAIL.n1 2.34102
R422 VTAIL.n103 VTAIL.n101 1.99188
R423 VTAIL.n47 VTAIL.n1 1.99188
R424 VTAIL.n184 VTAIL.n158 1.93989
R425 VTAIL.n196 VTAIL.n152 1.93989
R426 VTAIL.n34 VTAIL.n8 1.93989
R427 VTAIL.n46 VTAIL.n2 1.93989
R428 VTAIL.n150 VTAIL.n106 1.93989
R429 VTAIL.n138 VTAIL.n112 1.93989
R430 VTAIL.n100 VTAIL.n56 1.93989
R431 VTAIL.n88 VTAIL.n62 1.93989
R432 VTAIL.n185 VTAIL.n156 1.16414
R433 VTAIL.n194 VTAIL.n193 1.16414
R434 VTAIL.n35 VTAIL.n6 1.16414
R435 VTAIL.n44 VTAIL.n43 1.16414
R436 VTAIL.n148 VTAIL.n147 1.16414
R437 VTAIL.n139 VTAIL.n110 1.16414
R438 VTAIL.n98 VTAIL.n97 1.16414
R439 VTAIL.n89 VTAIL.n60 1.16414
R440 VTAIL VTAIL.n199 0.703086
R441 VTAIL.n189 VTAIL.n188 0.388379
R442 VTAIL.n190 VTAIL.n154 0.388379
R443 VTAIL.n39 VTAIL.n38 0.388379
R444 VTAIL.n40 VTAIL.n4 0.388379
R445 VTAIL.n144 VTAIL.n108 0.388379
R446 VTAIL.n143 VTAIL.n142 0.388379
R447 VTAIL.n94 VTAIL.n58 0.388379
R448 VTAIL.n93 VTAIL.n92 0.388379
R449 VTAIL.n170 VTAIL.n169 0.155672
R450 VTAIL.n170 VTAIL.n161 0.155672
R451 VTAIL.n177 VTAIL.n161 0.155672
R452 VTAIL.n178 VTAIL.n177 0.155672
R453 VTAIL.n178 VTAIL.n157 0.155672
R454 VTAIL.n186 VTAIL.n157 0.155672
R455 VTAIL.n187 VTAIL.n186 0.155672
R456 VTAIL.n187 VTAIL.n153 0.155672
R457 VTAIL.n195 VTAIL.n153 0.155672
R458 VTAIL.n20 VTAIL.n19 0.155672
R459 VTAIL.n20 VTAIL.n11 0.155672
R460 VTAIL.n27 VTAIL.n11 0.155672
R461 VTAIL.n28 VTAIL.n27 0.155672
R462 VTAIL.n28 VTAIL.n7 0.155672
R463 VTAIL.n36 VTAIL.n7 0.155672
R464 VTAIL.n37 VTAIL.n36 0.155672
R465 VTAIL.n37 VTAIL.n3 0.155672
R466 VTAIL.n45 VTAIL.n3 0.155672
R467 VTAIL.n149 VTAIL.n107 0.155672
R468 VTAIL.n141 VTAIL.n107 0.155672
R469 VTAIL.n141 VTAIL.n140 0.155672
R470 VTAIL.n140 VTAIL.n111 0.155672
R471 VTAIL.n133 VTAIL.n111 0.155672
R472 VTAIL.n133 VTAIL.n132 0.155672
R473 VTAIL.n132 VTAIL.n116 0.155672
R474 VTAIL.n125 VTAIL.n116 0.155672
R475 VTAIL.n125 VTAIL.n124 0.155672
R476 VTAIL.n99 VTAIL.n57 0.155672
R477 VTAIL.n91 VTAIL.n57 0.155672
R478 VTAIL.n91 VTAIL.n90 0.155672
R479 VTAIL.n90 VTAIL.n61 0.155672
R480 VTAIL.n83 VTAIL.n61 0.155672
R481 VTAIL.n83 VTAIL.n82 0.155672
R482 VTAIL.n82 VTAIL.n66 0.155672
R483 VTAIL.n75 VTAIL.n66 0.155672
R484 VTAIL.n75 VTAIL.n74 0.155672
R485 VDD1.n40 VDD1.n0 756.745
R486 VDD1.n87 VDD1.n47 756.745
R487 VDD1.n41 VDD1.n40 585
R488 VDD1.n39 VDD1.n38 585
R489 VDD1.n37 VDD1.n3 585
R490 VDD1.n7 VDD1.n4 585
R491 VDD1.n32 VDD1.n31 585
R492 VDD1.n30 VDD1.n29 585
R493 VDD1.n9 VDD1.n8 585
R494 VDD1.n24 VDD1.n23 585
R495 VDD1.n22 VDD1.n21 585
R496 VDD1.n13 VDD1.n12 585
R497 VDD1.n16 VDD1.n15 585
R498 VDD1.n62 VDD1.n61 585
R499 VDD1.n59 VDD1.n58 585
R500 VDD1.n68 VDD1.n67 585
R501 VDD1.n70 VDD1.n69 585
R502 VDD1.n55 VDD1.n54 585
R503 VDD1.n76 VDD1.n75 585
R504 VDD1.n79 VDD1.n78 585
R505 VDD1.n77 VDD1.n51 585
R506 VDD1.n84 VDD1.n50 585
R507 VDD1.n86 VDD1.n85 585
R508 VDD1.n88 VDD1.n87 585
R509 VDD1.t2 VDD1.n14 329.039
R510 VDD1.t6 VDD1.n60 329.038
R511 VDD1.n40 VDD1.n39 171.744
R512 VDD1.n39 VDD1.n3 171.744
R513 VDD1.n7 VDD1.n3 171.744
R514 VDD1.n31 VDD1.n7 171.744
R515 VDD1.n31 VDD1.n30 171.744
R516 VDD1.n30 VDD1.n8 171.744
R517 VDD1.n23 VDD1.n8 171.744
R518 VDD1.n23 VDD1.n22 171.744
R519 VDD1.n22 VDD1.n12 171.744
R520 VDD1.n15 VDD1.n12 171.744
R521 VDD1.n61 VDD1.n58 171.744
R522 VDD1.n68 VDD1.n58 171.744
R523 VDD1.n69 VDD1.n68 171.744
R524 VDD1.n69 VDD1.n54 171.744
R525 VDD1.n76 VDD1.n54 171.744
R526 VDD1.n78 VDD1.n76 171.744
R527 VDD1.n78 VDD1.n77 171.744
R528 VDD1.n77 VDD1.n50 171.744
R529 VDD1.n86 VDD1.n50 171.744
R530 VDD1.n87 VDD1.n86 171.744
R531 VDD1.n15 VDD1.t2 85.8723
R532 VDD1.n61 VDD1.t6 85.8723
R533 VDD1.n95 VDD1.n94 84.4705
R534 VDD1.n46 VDD1.n45 82.2437
R535 VDD1.n97 VDD1.n96 82.2435
R536 VDD1.n93 VDD1.n92 82.2435
R537 VDD1.n46 VDD1.n44 53.8466
R538 VDD1.n93 VDD1.n91 53.8466
R539 VDD1.n97 VDD1.n95 47.7056
R540 VDD1.n38 VDD1.n37 13.1884
R541 VDD1.n85 VDD1.n84 13.1884
R542 VDD1.n41 VDD1.n2 12.8005
R543 VDD1.n36 VDD1.n4 12.8005
R544 VDD1.n83 VDD1.n51 12.8005
R545 VDD1.n88 VDD1.n49 12.8005
R546 VDD1.n42 VDD1.n0 12.0247
R547 VDD1.n33 VDD1.n32 12.0247
R548 VDD1.n80 VDD1.n79 12.0247
R549 VDD1.n89 VDD1.n47 12.0247
R550 VDD1.n29 VDD1.n6 11.249
R551 VDD1.n75 VDD1.n53 11.249
R552 VDD1.n16 VDD1.n14 10.7239
R553 VDD1.n62 VDD1.n60 10.7239
R554 VDD1.n28 VDD1.n9 10.4732
R555 VDD1.n74 VDD1.n55 10.4732
R556 VDD1.n25 VDD1.n24 9.69747
R557 VDD1.n71 VDD1.n70 9.69747
R558 VDD1.n44 VDD1.n43 9.45567
R559 VDD1.n91 VDD1.n90 9.45567
R560 VDD1.n18 VDD1.n17 9.3005
R561 VDD1.n20 VDD1.n19 9.3005
R562 VDD1.n11 VDD1.n10 9.3005
R563 VDD1.n26 VDD1.n25 9.3005
R564 VDD1.n28 VDD1.n27 9.3005
R565 VDD1.n6 VDD1.n5 9.3005
R566 VDD1.n34 VDD1.n33 9.3005
R567 VDD1.n36 VDD1.n35 9.3005
R568 VDD1.n43 VDD1.n42 9.3005
R569 VDD1.n2 VDD1.n1 9.3005
R570 VDD1.n90 VDD1.n89 9.3005
R571 VDD1.n49 VDD1.n48 9.3005
R572 VDD1.n64 VDD1.n63 9.3005
R573 VDD1.n66 VDD1.n65 9.3005
R574 VDD1.n57 VDD1.n56 9.3005
R575 VDD1.n72 VDD1.n71 9.3005
R576 VDD1.n74 VDD1.n73 9.3005
R577 VDD1.n53 VDD1.n52 9.3005
R578 VDD1.n81 VDD1.n80 9.3005
R579 VDD1.n83 VDD1.n82 9.3005
R580 VDD1.n21 VDD1.n11 8.92171
R581 VDD1.n67 VDD1.n57 8.92171
R582 VDD1.n20 VDD1.n13 8.14595
R583 VDD1.n66 VDD1.n59 8.14595
R584 VDD1.n17 VDD1.n16 7.3702
R585 VDD1.n63 VDD1.n62 7.3702
R586 VDD1.n17 VDD1.n13 5.81868
R587 VDD1.n63 VDD1.n59 5.81868
R588 VDD1.n21 VDD1.n20 5.04292
R589 VDD1.n67 VDD1.n66 5.04292
R590 VDD1.n24 VDD1.n11 4.26717
R591 VDD1.n70 VDD1.n57 4.26717
R592 VDD1.n96 VDD1.t8 3.77138
R593 VDD1.n96 VDD1.t9 3.77138
R594 VDD1.n45 VDD1.t3 3.77138
R595 VDD1.n45 VDD1.t7 3.77138
R596 VDD1.n94 VDD1.t5 3.77138
R597 VDD1.n94 VDD1.t0 3.77138
R598 VDD1.n92 VDD1.t1 3.77138
R599 VDD1.n92 VDD1.t4 3.77138
R600 VDD1.n25 VDD1.n9 3.49141
R601 VDD1.n71 VDD1.n55 3.49141
R602 VDD1.n29 VDD1.n28 2.71565
R603 VDD1.n75 VDD1.n74 2.71565
R604 VDD1.n18 VDD1.n14 2.41285
R605 VDD1.n64 VDD1.n60 2.41285
R606 VDD1 VDD1.n97 2.22464
R607 VDD1.n44 VDD1.n0 1.93989
R608 VDD1.n32 VDD1.n6 1.93989
R609 VDD1.n79 VDD1.n53 1.93989
R610 VDD1.n91 VDD1.n47 1.93989
R611 VDD1.n42 VDD1.n41 1.16414
R612 VDD1.n33 VDD1.n4 1.16414
R613 VDD1.n80 VDD1.n51 1.16414
R614 VDD1.n89 VDD1.n88 1.16414
R615 VDD1 VDD1.n46 0.819465
R616 VDD1.n95 VDD1.n93 0.70593
R617 VDD1.n38 VDD1.n2 0.388379
R618 VDD1.n37 VDD1.n36 0.388379
R619 VDD1.n84 VDD1.n83 0.388379
R620 VDD1.n85 VDD1.n49 0.388379
R621 VDD1.n43 VDD1.n1 0.155672
R622 VDD1.n35 VDD1.n1 0.155672
R623 VDD1.n35 VDD1.n34 0.155672
R624 VDD1.n34 VDD1.n5 0.155672
R625 VDD1.n27 VDD1.n5 0.155672
R626 VDD1.n27 VDD1.n26 0.155672
R627 VDD1.n26 VDD1.n10 0.155672
R628 VDD1.n19 VDD1.n10 0.155672
R629 VDD1.n19 VDD1.n18 0.155672
R630 VDD1.n65 VDD1.n64 0.155672
R631 VDD1.n65 VDD1.n56 0.155672
R632 VDD1.n72 VDD1.n56 0.155672
R633 VDD1.n73 VDD1.n72 0.155672
R634 VDD1.n73 VDD1.n52 0.155672
R635 VDD1.n81 VDD1.n52 0.155672
R636 VDD1.n82 VDD1.n81 0.155672
R637 VDD1.n82 VDD1.n48 0.155672
R638 VDD1.n90 VDD1.n48 0.155672
R639 VN.n94 VN.n93 161.3
R640 VN.n92 VN.n49 161.3
R641 VN.n91 VN.n90 161.3
R642 VN.n89 VN.n50 161.3
R643 VN.n88 VN.n87 161.3
R644 VN.n86 VN.n51 161.3
R645 VN.n85 VN.n84 161.3
R646 VN.n83 VN.n82 161.3
R647 VN.n81 VN.n53 161.3
R648 VN.n80 VN.n79 161.3
R649 VN.n78 VN.n54 161.3
R650 VN.n77 VN.n76 161.3
R651 VN.n75 VN.n55 161.3
R652 VN.n74 VN.n73 161.3
R653 VN.n72 VN.n71 161.3
R654 VN.n70 VN.n57 161.3
R655 VN.n69 VN.n68 161.3
R656 VN.n67 VN.n58 161.3
R657 VN.n66 VN.n65 161.3
R658 VN.n64 VN.n59 161.3
R659 VN.n63 VN.n62 161.3
R660 VN.n46 VN.n45 161.3
R661 VN.n44 VN.n1 161.3
R662 VN.n43 VN.n42 161.3
R663 VN.n41 VN.n2 161.3
R664 VN.n40 VN.n39 161.3
R665 VN.n38 VN.n3 161.3
R666 VN.n37 VN.n36 161.3
R667 VN.n35 VN.n34 161.3
R668 VN.n33 VN.n5 161.3
R669 VN.n32 VN.n31 161.3
R670 VN.n30 VN.n6 161.3
R671 VN.n29 VN.n28 161.3
R672 VN.n27 VN.n7 161.3
R673 VN.n26 VN.n25 161.3
R674 VN.n24 VN.n23 161.3
R675 VN.n22 VN.n9 161.3
R676 VN.n21 VN.n20 161.3
R677 VN.n19 VN.n10 161.3
R678 VN.n18 VN.n17 161.3
R679 VN.n16 VN.n11 161.3
R680 VN.n15 VN.n14 161.3
R681 VN.n61 VN.t4 98.0243
R682 VN.n13 VN.t7 98.0243
R683 VN.n47 VN.n0 74.9986
R684 VN.n95 VN.n48 74.9986
R685 VN.n12 VN.t9 64.9199
R686 VN.n8 VN.t2 64.9199
R687 VN.n4 VN.t8 64.9199
R688 VN.n0 VN.t3 64.9199
R689 VN.n60 VN.t5 64.9199
R690 VN.n56 VN.t6 64.9199
R691 VN.n52 VN.t0 64.9199
R692 VN.n48 VN.t1 64.9199
R693 VN.n13 VN.n12 60.6744
R694 VN.n61 VN.n60 60.6744
R695 VN VN.n95 54.0777
R696 VN.n43 VN.n2 44.9365
R697 VN.n91 VN.n50 44.9365
R698 VN.n17 VN.n10 42.0302
R699 VN.n32 VN.n6 42.0302
R700 VN.n65 VN.n58 42.0302
R701 VN.n80 VN.n54 42.0302
R702 VN.n21 VN.n10 39.1239
R703 VN.n28 VN.n6 39.1239
R704 VN.n69 VN.n58 39.1239
R705 VN.n76 VN.n54 39.1239
R706 VN.n39 VN.n2 36.2176
R707 VN.n87 VN.n50 36.2176
R708 VN.n16 VN.n15 24.5923
R709 VN.n17 VN.n16 24.5923
R710 VN.n22 VN.n21 24.5923
R711 VN.n23 VN.n22 24.5923
R712 VN.n27 VN.n26 24.5923
R713 VN.n28 VN.n27 24.5923
R714 VN.n33 VN.n32 24.5923
R715 VN.n34 VN.n33 24.5923
R716 VN.n38 VN.n37 24.5923
R717 VN.n39 VN.n38 24.5923
R718 VN.n44 VN.n43 24.5923
R719 VN.n45 VN.n44 24.5923
R720 VN.n65 VN.n64 24.5923
R721 VN.n64 VN.n63 24.5923
R722 VN.n76 VN.n75 24.5923
R723 VN.n75 VN.n74 24.5923
R724 VN.n71 VN.n70 24.5923
R725 VN.n70 VN.n69 24.5923
R726 VN.n87 VN.n86 24.5923
R727 VN.n86 VN.n85 24.5923
R728 VN.n82 VN.n81 24.5923
R729 VN.n81 VN.n80 24.5923
R730 VN.n93 VN.n92 24.5923
R731 VN.n92 VN.n91 24.5923
R732 VN.n45 VN.n0 15.2474
R733 VN.n93 VN.n48 15.2474
R734 VN.n15 VN.n12 13.7719
R735 VN.n34 VN.n4 13.7719
R736 VN.n63 VN.n60 13.7719
R737 VN.n82 VN.n52 13.7719
R738 VN.n23 VN.n8 12.2964
R739 VN.n26 VN.n8 12.2964
R740 VN.n74 VN.n56 12.2964
R741 VN.n71 VN.n56 12.2964
R742 VN.n37 VN.n4 10.8209
R743 VN.n85 VN.n52 10.8209
R744 VN.n62 VN.n61 4.12006
R745 VN.n14 VN.n13 4.12006
R746 VN.n95 VN.n94 0.354861
R747 VN.n47 VN.n46 0.354861
R748 VN VN.n47 0.267071
R749 VN.n94 VN.n49 0.189894
R750 VN.n90 VN.n49 0.189894
R751 VN.n90 VN.n89 0.189894
R752 VN.n89 VN.n88 0.189894
R753 VN.n88 VN.n51 0.189894
R754 VN.n84 VN.n51 0.189894
R755 VN.n84 VN.n83 0.189894
R756 VN.n83 VN.n53 0.189894
R757 VN.n79 VN.n53 0.189894
R758 VN.n79 VN.n78 0.189894
R759 VN.n78 VN.n77 0.189894
R760 VN.n77 VN.n55 0.189894
R761 VN.n73 VN.n55 0.189894
R762 VN.n73 VN.n72 0.189894
R763 VN.n72 VN.n57 0.189894
R764 VN.n68 VN.n57 0.189894
R765 VN.n68 VN.n67 0.189894
R766 VN.n67 VN.n66 0.189894
R767 VN.n66 VN.n59 0.189894
R768 VN.n62 VN.n59 0.189894
R769 VN.n14 VN.n11 0.189894
R770 VN.n18 VN.n11 0.189894
R771 VN.n19 VN.n18 0.189894
R772 VN.n20 VN.n19 0.189894
R773 VN.n20 VN.n9 0.189894
R774 VN.n24 VN.n9 0.189894
R775 VN.n25 VN.n24 0.189894
R776 VN.n25 VN.n7 0.189894
R777 VN.n29 VN.n7 0.189894
R778 VN.n30 VN.n29 0.189894
R779 VN.n31 VN.n30 0.189894
R780 VN.n31 VN.n5 0.189894
R781 VN.n35 VN.n5 0.189894
R782 VN.n36 VN.n35 0.189894
R783 VN.n36 VN.n3 0.189894
R784 VN.n40 VN.n3 0.189894
R785 VN.n41 VN.n40 0.189894
R786 VN.n42 VN.n41 0.189894
R787 VN.n42 VN.n1 0.189894
R788 VN.n46 VN.n1 0.189894
R789 VDD2.n89 VDD2.n49 756.745
R790 VDD2.n40 VDD2.n0 756.745
R791 VDD2.n90 VDD2.n89 585
R792 VDD2.n88 VDD2.n87 585
R793 VDD2.n86 VDD2.n52 585
R794 VDD2.n56 VDD2.n53 585
R795 VDD2.n81 VDD2.n80 585
R796 VDD2.n79 VDD2.n78 585
R797 VDD2.n58 VDD2.n57 585
R798 VDD2.n73 VDD2.n72 585
R799 VDD2.n71 VDD2.n70 585
R800 VDD2.n62 VDD2.n61 585
R801 VDD2.n65 VDD2.n64 585
R802 VDD2.n15 VDD2.n14 585
R803 VDD2.n12 VDD2.n11 585
R804 VDD2.n21 VDD2.n20 585
R805 VDD2.n23 VDD2.n22 585
R806 VDD2.n8 VDD2.n7 585
R807 VDD2.n29 VDD2.n28 585
R808 VDD2.n32 VDD2.n31 585
R809 VDD2.n30 VDD2.n4 585
R810 VDD2.n37 VDD2.n3 585
R811 VDD2.n39 VDD2.n38 585
R812 VDD2.n41 VDD2.n40 585
R813 VDD2.t8 VDD2.n63 329.039
R814 VDD2.t2 VDD2.n13 329.038
R815 VDD2.n89 VDD2.n88 171.744
R816 VDD2.n88 VDD2.n52 171.744
R817 VDD2.n56 VDD2.n52 171.744
R818 VDD2.n80 VDD2.n56 171.744
R819 VDD2.n80 VDD2.n79 171.744
R820 VDD2.n79 VDD2.n57 171.744
R821 VDD2.n72 VDD2.n57 171.744
R822 VDD2.n72 VDD2.n71 171.744
R823 VDD2.n71 VDD2.n61 171.744
R824 VDD2.n64 VDD2.n61 171.744
R825 VDD2.n14 VDD2.n11 171.744
R826 VDD2.n21 VDD2.n11 171.744
R827 VDD2.n22 VDD2.n21 171.744
R828 VDD2.n22 VDD2.n7 171.744
R829 VDD2.n29 VDD2.n7 171.744
R830 VDD2.n31 VDD2.n29 171.744
R831 VDD2.n31 VDD2.n30 171.744
R832 VDD2.n30 VDD2.n3 171.744
R833 VDD2.n39 VDD2.n3 171.744
R834 VDD2.n40 VDD2.n39 171.744
R835 VDD2.n64 VDD2.t8 85.8723
R836 VDD2.n14 VDD2.t2 85.8723
R837 VDD2.n48 VDD2.n47 84.4705
R838 VDD2 VDD2.n97 84.4676
R839 VDD2.n96 VDD2.n95 82.2437
R840 VDD2.n46 VDD2.n45 82.2435
R841 VDD2.n46 VDD2.n44 53.8466
R842 VDD2.n94 VDD2.n93 50.8035
R843 VDD2.n94 VDD2.n48 45.6011
R844 VDD2.n87 VDD2.n86 13.1884
R845 VDD2.n38 VDD2.n37 13.1884
R846 VDD2.n90 VDD2.n51 12.8005
R847 VDD2.n85 VDD2.n53 12.8005
R848 VDD2.n36 VDD2.n4 12.8005
R849 VDD2.n41 VDD2.n2 12.8005
R850 VDD2.n91 VDD2.n49 12.0247
R851 VDD2.n82 VDD2.n81 12.0247
R852 VDD2.n33 VDD2.n32 12.0247
R853 VDD2.n42 VDD2.n0 12.0247
R854 VDD2.n78 VDD2.n55 11.249
R855 VDD2.n28 VDD2.n6 11.249
R856 VDD2.n65 VDD2.n63 10.7239
R857 VDD2.n15 VDD2.n13 10.7239
R858 VDD2.n77 VDD2.n58 10.4732
R859 VDD2.n27 VDD2.n8 10.4732
R860 VDD2.n74 VDD2.n73 9.69747
R861 VDD2.n24 VDD2.n23 9.69747
R862 VDD2.n93 VDD2.n92 9.45567
R863 VDD2.n44 VDD2.n43 9.45567
R864 VDD2.n67 VDD2.n66 9.3005
R865 VDD2.n69 VDD2.n68 9.3005
R866 VDD2.n60 VDD2.n59 9.3005
R867 VDD2.n75 VDD2.n74 9.3005
R868 VDD2.n77 VDD2.n76 9.3005
R869 VDD2.n55 VDD2.n54 9.3005
R870 VDD2.n83 VDD2.n82 9.3005
R871 VDD2.n85 VDD2.n84 9.3005
R872 VDD2.n92 VDD2.n91 9.3005
R873 VDD2.n51 VDD2.n50 9.3005
R874 VDD2.n43 VDD2.n42 9.3005
R875 VDD2.n2 VDD2.n1 9.3005
R876 VDD2.n17 VDD2.n16 9.3005
R877 VDD2.n19 VDD2.n18 9.3005
R878 VDD2.n10 VDD2.n9 9.3005
R879 VDD2.n25 VDD2.n24 9.3005
R880 VDD2.n27 VDD2.n26 9.3005
R881 VDD2.n6 VDD2.n5 9.3005
R882 VDD2.n34 VDD2.n33 9.3005
R883 VDD2.n36 VDD2.n35 9.3005
R884 VDD2.n70 VDD2.n60 8.92171
R885 VDD2.n20 VDD2.n10 8.92171
R886 VDD2.n69 VDD2.n62 8.14595
R887 VDD2.n19 VDD2.n12 8.14595
R888 VDD2.n66 VDD2.n65 7.3702
R889 VDD2.n16 VDD2.n15 7.3702
R890 VDD2.n66 VDD2.n62 5.81868
R891 VDD2.n16 VDD2.n12 5.81868
R892 VDD2.n70 VDD2.n69 5.04292
R893 VDD2.n20 VDD2.n19 5.04292
R894 VDD2.n73 VDD2.n60 4.26717
R895 VDD2.n23 VDD2.n10 4.26717
R896 VDD2.n97 VDD2.t4 3.77138
R897 VDD2.n97 VDD2.t5 3.77138
R898 VDD2.n95 VDD2.t9 3.77138
R899 VDD2.n95 VDD2.t3 3.77138
R900 VDD2.n47 VDD2.t1 3.77138
R901 VDD2.n47 VDD2.t6 3.77138
R902 VDD2.n45 VDD2.t0 3.77138
R903 VDD2.n45 VDD2.t7 3.77138
R904 VDD2.n74 VDD2.n58 3.49141
R905 VDD2.n24 VDD2.n8 3.49141
R906 VDD2.n96 VDD2.n94 3.0436
R907 VDD2.n78 VDD2.n77 2.71565
R908 VDD2.n28 VDD2.n27 2.71565
R909 VDD2.n67 VDD2.n63 2.41285
R910 VDD2.n17 VDD2.n13 2.41285
R911 VDD2.n93 VDD2.n49 1.93989
R912 VDD2.n81 VDD2.n55 1.93989
R913 VDD2.n32 VDD2.n6 1.93989
R914 VDD2.n44 VDD2.n0 1.93989
R915 VDD2.n91 VDD2.n90 1.16414
R916 VDD2.n82 VDD2.n53 1.16414
R917 VDD2.n33 VDD2.n4 1.16414
R918 VDD2.n42 VDD2.n41 1.16414
R919 VDD2 VDD2.n96 0.819465
R920 VDD2.n48 VDD2.n46 0.70593
R921 VDD2.n87 VDD2.n51 0.388379
R922 VDD2.n86 VDD2.n85 0.388379
R923 VDD2.n37 VDD2.n36 0.388379
R924 VDD2.n38 VDD2.n2 0.388379
R925 VDD2.n92 VDD2.n50 0.155672
R926 VDD2.n84 VDD2.n50 0.155672
R927 VDD2.n84 VDD2.n83 0.155672
R928 VDD2.n83 VDD2.n54 0.155672
R929 VDD2.n76 VDD2.n54 0.155672
R930 VDD2.n76 VDD2.n75 0.155672
R931 VDD2.n75 VDD2.n59 0.155672
R932 VDD2.n68 VDD2.n59 0.155672
R933 VDD2.n68 VDD2.n67 0.155672
R934 VDD2.n18 VDD2.n17 0.155672
R935 VDD2.n18 VDD2.n9 0.155672
R936 VDD2.n25 VDD2.n9 0.155672
R937 VDD2.n26 VDD2.n25 0.155672
R938 VDD2.n26 VDD2.n5 0.155672
R939 VDD2.n34 VDD2.n5 0.155672
R940 VDD2.n35 VDD2.n34 0.155672
R941 VDD2.n35 VDD2.n1 0.155672
R942 VDD2.n43 VDD2.n1 0.155672
R943 B.n438 B.n437 585
R944 B.n436 B.n149 585
R945 B.n435 B.n434 585
R946 B.n433 B.n150 585
R947 B.n432 B.n431 585
R948 B.n430 B.n151 585
R949 B.n429 B.n428 585
R950 B.n427 B.n152 585
R951 B.n426 B.n425 585
R952 B.n424 B.n153 585
R953 B.n423 B.n422 585
R954 B.n421 B.n154 585
R955 B.n420 B.n419 585
R956 B.n418 B.n155 585
R957 B.n417 B.n416 585
R958 B.n415 B.n156 585
R959 B.n414 B.n413 585
R960 B.n412 B.n157 585
R961 B.n411 B.n410 585
R962 B.n409 B.n158 585
R963 B.n408 B.n407 585
R964 B.n406 B.n159 585
R965 B.n405 B.n404 585
R966 B.n403 B.n160 585
R967 B.n402 B.n401 585
R968 B.n400 B.n161 585
R969 B.n399 B.n398 585
R970 B.n397 B.n162 585
R971 B.n396 B.n395 585
R972 B.n394 B.n163 585
R973 B.n393 B.n392 585
R974 B.n391 B.n164 585
R975 B.n390 B.n389 585
R976 B.n385 B.n165 585
R977 B.n384 B.n383 585
R978 B.n382 B.n166 585
R979 B.n381 B.n380 585
R980 B.n379 B.n167 585
R981 B.n378 B.n377 585
R982 B.n376 B.n168 585
R983 B.n375 B.n374 585
R984 B.n372 B.n169 585
R985 B.n371 B.n370 585
R986 B.n369 B.n172 585
R987 B.n368 B.n367 585
R988 B.n366 B.n173 585
R989 B.n365 B.n364 585
R990 B.n363 B.n174 585
R991 B.n362 B.n361 585
R992 B.n360 B.n175 585
R993 B.n359 B.n358 585
R994 B.n357 B.n176 585
R995 B.n356 B.n355 585
R996 B.n354 B.n177 585
R997 B.n353 B.n352 585
R998 B.n351 B.n178 585
R999 B.n350 B.n349 585
R1000 B.n348 B.n179 585
R1001 B.n347 B.n346 585
R1002 B.n345 B.n180 585
R1003 B.n344 B.n343 585
R1004 B.n342 B.n181 585
R1005 B.n341 B.n340 585
R1006 B.n339 B.n182 585
R1007 B.n338 B.n337 585
R1008 B.n336 B.n183 585
R1009 B.n335 B.n334 585
R1010 B.n333 B.n184 585
R1011 B.n332 B.n331 585
R1012 B.n330 B.n185 585
R1013 B.n329 B.n328 585
R1014 B.n327 B.n186 585
R1015 B.n326 B.n325 585
R1016 B.n439 B.n148 585
R1017 B.n441 B.n440 585
R1018 B.n442 B.n147 585
R1019 B.n444 B.n443 585
R1020 B.n445 B.n146 585
R1021 B.n447 B.n446 585
R1022 B.n448 B.n145 585
R1023 B.n450 B.n449 585
R1024 B.n451 B.n144 585
R1025 B.n453 B.n452 585
R1026 B.n454 B.n143 585
R1027 B.n456 B.n455 585
R1028 B.n457 B.n142 585
R1029 B.n459 B.n458 585
R1030 B.n460 B.n141 585
R1031 B.n462 B.n461 585
R1032 B.n463 B.n140 585
R1033 B.n465 B.n464 585
R1034 B.n466 B.n139 585
R1035 B.n468 B.n467 585
R1036 B.n469 B.n138 585
R1037 B.n471 B.n470 585
R1038 B.n472 B.n137 585
R1039 B.n474 B.n473 585
R1040 B.n475 B.n136 585
R1041 B.n477 B.n476 585
R1042 B.n478 B.n135 585
R1043 B.n480 B.n479 585
R1044 B.n481 B.n134 585
R1045 B.n483 B.n482 585
R1046 B.n484 B.n133 585
R1047 B.n486 B.n485 585
R1048 B.n487 B.n132 585
R1049 B.n489 B.n488 585
R1050 B.n490 B.n131 585
R1051 B.n492 B.n491 585
R1052 B.n493 B.n130 585
R1053 B.n495 B.n494 585
R1054 B.n496 B.n129 585
R1055 B.n498 B.n497 585
R1056 B.n499 B.n128 585
R1057 B.n501 B.n500 585
R1058 B.n502 B.n127 585
R1059 B.n504 B.n503 585
R1060 B.n505 B.n126 585
R1061 B.n507 B.n506 585
R1062 B.n508 B.n125 585
R1063 B.n510 B.n509 585
R1064 B.n511 B.n124 585
R1065 B.n513 B.n512 585
R1066 B.n514 B.n123 585
R1067 B.n516 B.n515 585
R1068 B.n517 B.n122 585
R1069 B.n519 B.n518 585
R1070 B.n520 B.n121 585
R1071 B.n522 B.n521 585
R1072 B.n523 B.n120 585
R1073 B.n525 B.n524 585
R1074 B.n526 B.n119 585
R1075 B.n528 B.n527 585
R1076 B.n529 B.n118 585
R1077 B.n531 B.n530 585
R1078 B.n532 B.n117 585
R1079 B.n534 B.n533 585
R1080 B.n535 B.n116 585
R1081 B.n537 B.n536 585
R1082 B.n538 B.n115 585
R1083 B.n540 B.n539 585
R1084 B.n541 B.n114 585
R1085 B.n543 B.n542 585
R1086 B.n544 B.n113 585
R1087 B.n546 B.n545 585
R1088 B.n547 B.n112 585
R1089 B.n549 B.n548 585
R1090 B.n550 B.n111 585
R1091 B.n552 B.n551 585
R1092 B.n553 B.n110 585
R1093 B.n555 B.n554 585
R1094 B.n556 B.n109 585
R1095 B.n558 B.n557 585
R1096 B.n559 B.n108 585
R1097 B.n561 B.n560 585
R1098 B.n562 B.n107 585
R1099 B.n564 B.n563 585
R1100 B.n565 B.n106 585
R1101 B.n567 B.n566 585
R1102 B.n568 B.n105 585
R1103 B.n570 B.n569 585
R1104 B.n571 B.n104 585
R1105 B.n573 B.n572 585
R1106 B.n574 B.n103 585
R1107 B.n576 B.n575 585
R1108 B.n577 B.n102 585
R1109 B.n579 B.n578 585
R1110 B.n580 B.n101 585
R1111 B.n582 B.n581 585
R1112 B.n583 B.n100 585
R1113 B.n585 B.n584 585
R1114 B.n586 B.n99 585
R1115 B.n588 B.n587 585
R1116 B.n589 B.n98 585
R1117 B.n591 B.n590 585
R1118 B.n592 B.n97 585
R1119 B.n594 B.n593 585
R1120 B.n595 B.n96 585
R1121 B.n597 B.n596 585
R1122 B.n598 B.n95 585
R1123 B.n600 B.n599 585
R1124 B.n601 B.n94 585
R1125 B.n603 B.n602 585
R1126 B.n604 B.n93 585
R1127 B.n606 B.n605 585
R1128 B.n607 B.n92 585
R1129 B.n609 B.n608 585
R1130 B.n610 B.n91 585
R1131 B.n612 B.n611 585
R1132 B.n613 B.n90 585
R1133 B.n615 B.n614 585
R1134 B.n616 B.n89 585
R1135 B.n618 B.n617 585
R1136 B.n619 B.n88 585
R1137 B.n621 B.n620 585
R1138 B.n622 B.n87 585
R1139 B.n624 B.n623 585
R1140 B.n625 B.n86 585
R1141 B.n627 B.n626 585
R1142 B.n628 B.n85 585
R1143 B.n630 B.n629 585
R1144 B.n631 B.n84 585
R1145 B.n633 B.n632 585
R1146 B.n634 B.n83 585
R1147 B.n636 B.n635 585
R1148 B.n637 B.n82 585
R1149 B.n639 B.n638 585
R1150 B.n640 B.n81 585
R1151 B.n642 B.n641 585
R1152 B.n643 B.n80 585
R1153 B.n645 B.n644 585
R1154 B.n646 B.n79 585
R1155 B.n648 B.n647 585
R1156 B.n649 B.n78 585
R1157 B.n651 B.n650 585
R1158 B.n762 B.n37 585
R1159 B.n761 B.n760 585
R1160 B.n759 B.n38 585
R1161 B.n758 B.n757 585
R1162 B.n756 B.n39 585
R1163 B.n755 B.n754 585
R1164 B.n753 B.n40 585
R1165 B.n752 B.n751 585
R1166 B.n750 B.n41 585
R1167 B.n749 B.n748 585
R1168 B.n747 B.n42 585
R1169 B.n746 B.n745 585
R1170 B.n744 B.n43 585
R1171 B.n743 B.n742 585
R1172 B.n741 B.n44 585
R1173 B.n740 B.n739 585
R1174 B.n738 B.n45 585
R1175 B.n737 B.n736 585
R1176 B.n735 B.n46 585
R1177 B.n734 B.n733 585
R1178 B.n732 B.n47 585
R1179 B.n731 B.n730 585
R1180 B.n729 B.n48 585
R1181 B.n728 B.n727 585
R1182 B.n726 B.n49 585
R1183 B.n725 B.n724 585
R1184 B.n723 B.n50 585
R1185 B.n722 B.n721 585
R1186 B.n720 B.n51 585
R1187 B.n719 B.n718 585
R1188 B.n717 B.n52 585
R1189 B.n716 B.n715 585
R1190 B.n713 B.n53 585
R1191 B.n712 B.n711 585
R1192 B.n710 B.n56 585
R1193 B.n709 B.n708 585
R1194 B.n707 B.n57 585
R1195 B.n706 B.n705 585
R1196 B.n704 B.n58 585
R1197 B.n703 B.n702 585
R1198 B.n701 B.n59 585
R1199 B.n699 B.n698 585
R1200 B.n697 B.n62 585
R1201 B.n696 B.n695 585
R1202 B.n694 B.n63 585
R1203 B.n693 B.n692 585
R1204 B.n691 B.n64 585
R1205 B.n690 B.n689 585
R1206 B.n688 B.n65 585
R1207 B.n687 B.n686 585
R1208 B.n685 B.n66 585
R1209 B.n684 B.n683 585
R1210 B.n682 B.n67 585
R1211 B.n681 B.n680 585
R1212 B.n679 B.n68 585
R1213 B.n678 B.n677 585
R1214 B.n676 B.n69 585
R1215 B.n675 B.n674 585
R1216 B.n673 B.n70 585
R1217 B.n672 B.n671 585
R1218 B.n670 B.n71 585
R1219 B.n669 B.n668 585
R1220 B.n667 B.n72 585
R1221 B.n666 B.n665 585
R1222 B.n664 B.n73 585
R1223 B.n663 B.n662 585
R1224 B.n661 B.n74 585
R1225 B.n660 B.n659 585
R1226 B.n658 B.n75 585
R1227 B.n657 B.n656 585
R1228 B.n655 B.n76 585
R1229 B.n654 B.n653 585
R1230 B.n652 B.n77 585
R1231 B.n764 B.n763 585
R1232 B.n765 B.n36 585
R1233 B.n767 B.n766 585
R1234 B.n768 B.n35 585
R1235 B.n770 B.n769 585
R1236 B.n771 B.n34 585
R1237 B.n773 B.n772 585
R1238 B.n774 B.n33 585
R1239 B.n776 B.n775 585
R1240 B.n777 B.n32 585
R1241 B.n779 B.n778 585
R1242 B.n780 B.n31 585
R1243 B.n782 B.n781 585
R1244 B.n783 B.n30 585
R1245 B.n785 B.n784 585
R1246 B.n786 B.n29 585
R1247 B.n788 B.n787 585
R1248 B.n789 B.n28 585
R1249 B.n791 B.n790 585
R1250 B.n792 B.n27 585
R1251 B.n794 B.n793 585
R1252 B.n795 B.n26 585
R1253 B.n797 B.n796 585
R1254 B.n798 B.n25 585
R1255 B.n800 B.n799 585
R1256 B.n801 B.n24 585
R1257 B.n803 B.n802 585
R1258 B.n804 B.n23 585
R1259 B.n806 B.n805 585
R1260 B.n807 B.n22 585
R1261 B.n809 B.n808 585
R1262 B.n810 B.n21 585
R1263 B.n812 B.n811 585
R1264 B.n813 B.n20 585
R1265 B.n815 B.n814 585
R1266 B.n816 B.n19 585
R1267 B.n818 B.n817 585
R1268 B.n819 B.n18 585
R1269 B.n821 B.n820 585
R1270 B.n822 B.n17 585
R1271 B.n824 B.n823 585
R1272 B.n825 B.n16 585
R1273 B.n827 B.n826 585
R1274 B.n828 B.n15 585
R1275 B.n830 B.n829 585
R1276 B.n831 B.n14 585
R1277 B.n833 B.n832 585
R1278 B.n834 B.n13 585
R1279 B.n836 B.n835 585
R1280 B.n837 B.n12 585
R1281 B.n839 B.n838 585
R1282 B.n840 B.n11 585
R1283 B.n842 B.n841 585
R1284 B.n843 B.n10 585
R1285 B.n845 B.n844 585
R1286 B.n846 B.n9 585
R1287 B.n848 B.n847 585
R1288 B.n849 B.n8 585
R1289 B.n851 B.n850 585
R1290 B.n852 B.n7 585
R1291 B.n854 B.n853 585
R1292 B.n855 B.n6 585
R1293 B.n857 B.n856 585
R1294 B.n858 B.n5 585
R1295 B.n860 B.n859 585
R1296 B.n861 B.n4 585
R1297 B.n863 B.n862 585
R1298 B.n864 B.n3 585
R1299 B.n866 B.n865 585
R1300 B.n867 B.n0 585
R1301 B.n2 B.n1 585
R1302 B.n222 B.n221 585
R1303 B.n224 B.n223 585
R1304 B.n225 B.n220 585
R1305 B.n227 B.n226 585
R1306 B.n228 B.n219 585
R1307 B.n230 B.n229 585
R1308 B.n231 B.n218 585
R1309 B.n233 B.n232 585
R1310 B.n234 B.n217 585
R1311 B.n236 B.n235 585
R1312 B.n237 B.n216 585
R1313 B.n239 B.n238 585
R1314 B.n240 B.n215 585
R1315 B.n242 B.n241 585
R1316 B.n243 B.n214 585
R1317 B.n245 B.n244 585
R1318 B.n246 B.n213 585
R1319 B.n248 B.n247 585
R1320 B.n249 B.n212 585
R1321 B.n251 B.n250 585
R1322 B.n252 B.n211 585
R1323 B.n254 B.n253 585
R1324 B.n255 B.n210 585
R1325 B.n257 B.n256 585
R1326 B.n258 B.n209 585
R1327 B.n260 B.n259 585
R1328 B.n261 B.n208 585
R1329 B.n263 B.n262 585
R1330 B.n264 B.n207 585
R1331 B.n266 B.n265 585
R1332 B.n267 B.n206 585
R1333 B.n269 B.n268 585
R1334 B.n270 B.n205 585
R1335 B.n272 B.n271 585
R1336 B.n273 B.n204 585
R1337 B.n275 B.n274 585
R1338 B.n276 B.n203 585
R1339 B.n278 B.n277 585
R1340 B.n279 B.n202 585
R1341 B.n281 B.n280 585
R1342 B.n282 B.n201 585
R1343 B.n284 B.n283 585
R1344 B.n285 B.n200 585
R1345 B.n287 B.n286 585
R1346 B.n288 B.n199 585
R1347 B.n290 B.n289 585
R1348 B.n291 B.n198 585
R1349 B.n293 B.n292 585
R1350 B.n294 B.n197 585
R1351 B.n296 B.n295 585
R1352 B.n297 B.n196 585
R1353 B.n299 B.n298 585
R1354 B.n300 B.n195 585
R1355 B.n302 B.n301 585
R1356 B.n303 B.n194 585
R1357 B.n305 B.n304 585
R1358 B.n306 B.n193 585
R1359 B.n308 B.n307 585
R1360 B.n309 B.n192 585
R1361 B.n311 B.n310 585
R1362 B.n312 B.n191 585
R1363 B.n314 B.n313 585
R1364 B.n315 B.n190 585
R1365 B.n317 B.n316 585
R1366 B.n318 B.n189 585
R1367 B.n320 B.n319 585
R1368 B.n321 B.n188 585
R1369 B.n323 B.n322 585
R1370 B.n324 B.n187 585
R1371 B.n326 B.n187 478.086
R1372 B.n439 B.n438 478.086
R1373 B.n650 B.n77 478.086
R1374 B.n764 B.n37 478.086
R1375 B.n386 B.t1 383.192
R1376 B.n60 B.t11 383.192
R1377 B.n170 B.t7 383.192
R1378 B.n54 B.t5 383.192
R1379 B.n387 B.t2 314.731
R1380 B.n61 B.t10 314.731
R1381 B.n171 B.t8 314.731
R1382 B.n55 B.t4 314.731
R1383 B.n170 B.t6 273.723
R1384 B.n386 B.t0 273.723
R1385 B.n60 B.t9 273.723
R1386 B.n54 B.t3 273.723
R1387 B.n869 B.n868 256.663
R1388 B.n868 B.n867 235.042
R1389 B.n868 B.n2 235.042
R1390 B.n327 B.n326 163.367
R1391 B.n328 B.n327 163.367
R1392 B.n328 B.n185 163.367
R1393 B.n332 B.n185 163.367
R1394 B.n333 B.n332 163.367
R1395 B.n334 B.n333 163.367
R1396 B.n334 B.n183 163.367
R1397 B.n338 B.n183 163.367
R1398 B.n339 B.n338 163.367
R1399 B.n340 B.n339 163.367
R1400 B.n340 B.n181 163.367
R1401 B.n344 B.n181 163.367
R1402 B.n345 B.n344 163.367
R1403 B.n346 B.n345 163.367
R1404 B.n346 B.n179 163.367
R1405 B.n350 B.n179 163.367
R1406 B.n351 B.n350 163.367
R1407 B.n352 B.n351 163.367
R1408 B.n352 B.n177 163.367
R1409 B.n356 B.n177 163.367
R1410 B.n357 B.n356 163.367
R1411 B.n358 B.n357 163.367
R1412 B.n358 B.n175 163.367
R1413 B.n362 B.n175 163.367
R1414 B.n363 B.n362 163.367
R1415 B.n364 B.n363 163.367
R1416 B.n364 B.n173 163.367
R1417 B.n368 B.n173 163.367
R1418 B.n369 B.n368 163.367
R1419 B.n370 B.n369 163.367
R1420 B.n370 B.n169 163.367
R1421 B.n375 B.n169 163.367
R1422 B.n376 B.n375 163.367
R1423 B.n377 B.n376 163.367
R1424 B.n377 B.n167 163.367
R1425 B.n381 B.n167 163.367
R1426 B.n382 B.n381 163.367
R1427 B.n383 B.n382 163.367
R1428 B.n383 B.n165 163.367
R1429 B.n390 B.n165 163.367
R1430 B.n391 B.n390 163.367
R1431 B.n392 B.n391 163.367
R1432 B.n392 B.n163 163.367
R1433 B.n396 B.n163 163.367
R1434 B.n397 B.n396 163.367
R1435 B.n398 B.n397 163.367
R1436 B.n398 B.n161 163.367
R1437 B.n402 B.n161 163.367
R1438 B.n403 B.n402 163.367
R1439 B.n404 B.n403 163.367
R1440 B.n404 B.n159 163.367
R1441 B.n408 B.n159 163.367
R1442 B.n409 B.n408 163.367
R1443 B.n410 B.n409 163.367
R1444 B.n410 B.n157 163.367
R1445 B.n414 B.n157 163.367
R1446 B.n415 B.n414 163.367
R1447 B.n416 B.n415 163.367
R1448 B.n416 B.n155 163.367
R1449 B.n420 B.n155 163.367
R1450 B.n421 B.n420 163.367
R1451 B.n422 B.n421 163.367
R1452 B.n422 B.n153 163.367
R1453 B.n426 B.n153 163.367
R1454 B.n427 B.n426 163.367
R1455 B.n428 B.n427 163.367
R1456 B.n428 B.n151 163.367
R1457 B.n432 B.n151 163.367
R1458 B.n433 B.n432 163.367
R1459 B.n434 B.n433 163.367
R1460 B.n434 B.n149 163.367
R1461 B.n438 B.n149 163.367
R1462 B.n650 B.n649 163.367
R1463 B.n649 B.n648 163.367
R1464 B.n648 B.n79 163.367
R1465 B.n644 B.n79 163.367
R1466 B.n644 B.n643 163.367
R1467 B.n643 B.n642 163.367
R1468 B.n642 B.n81 163.367
R1469 B.n638 B.n81 163.367
R1470 B.n638 B.n637 163.367
R1471 B.n637 B.n636 163.367
R1472 B.n636 B.n83 163.367
R1473 B.n632 B.n83 163.367
R1474 B.n632 B.n631 163.367
R1475 B.n631 B.n630 163.367
R1476 B.n630 B.n85 163.367
R1477 B.n626 B.n85 163.367
R1478 B.n626 B.n625 163.367
R1479 B.n625 B.n624 163.367
R1480 B.n624 B.n87 163.367
R1481 B.n620 B.n87 163.367
R1482 B.n620 B.n619 163.367
R1483 B.n619 B.n618 163.367
R1484 B.n618 B.n89 163.367
R1485 B.n614 B.n89 163.367
R1486 B.n614 B.n613 163.367
R1487 B.n613 B.n612 163.367
R1488 B.n612 B.n91 163.367
R1489 B.n608 B.n91 163.367
R1490 B.n608 B.n607 163.367
R1491 B.n607 B.n606 163.367
R1492 B.n606 B.n93 163.367
R1493 B.n602 B.n93 163.367
R1494 B.n602 B.n601 163.367
R1495 B.n601 B.n600 163.367
R1496 B.n600 B.n95 163.367
R1497 B.n596 B.n95 163.367
R1498 B.n596 B.n595 163.367
R1499 B.n595 B.n594 163.367
R1500 B.n594 B.n97 163.367
R1501 B.n590 B.n97 163.367
R1502 B.n590 B.n589 163.367
R1503 B.n589 B.n588 163.367
R1504 B.n588 B.n99 163.367
R1505 B.n584 B.n99 163.367
R1506 B.n584 B.n583 163.367
R1507 B.n583 B.n582 163.367
R1508 B.n582 B.n101 163.367
R1509 B.n578 B.n101 163.367
R1510 B.n578 B.n577 163.367
R1511 B.n577 B.n576 163.367
R1512 B.n576 B.n103 163.367
R1513 B.n572 B.n103 163.367
R1514 B.n572 B.n571 163.367
R1515 B.n571 B.n570 163.367
R1516 B.n570 B.n105 163.367
R1517 B.n566 B.n105 163.367
R1518 B.n566 B.n565 163.367
R1519 B.n565 B.n564 163.367
R1520 B.n564 B.n107 163.367
R1521 B.n560 B.n107 163.367
R1522 B.n560 B.n559 163.367
R1523 B.n559 B.n558 163.367
R1524 B.n558 B.n109 163.367
R1525 B.n554 B.n109 163.367
R1526 B.n554 B.n553 163.367
R1527 B.n553 B.n552 163.367
R1528 B.n552 B.n111 163.367
R1529 B.n548 B.n111 163.367
R1530 B.n548 B.n547 163.367
R1531 B.n547 B.n546 163.367
R1532 B.n546 B.n113 163.367
R1533 B.n542 B.n113 163.367
R1534 B.n542 B.n541 163.367
R1535 B.n541 B.n540 163.367
R1536 B.n540 B.n115 163.367
R1537 B.n536 B.n115 163.367
R1538 B.n536 B.n535 163.367
R1539 B.n535 B.n534 163.367
R1540 B.n534 B.n117 163.367
R1541 B.n530 B.n117 163.367
R1542 B.n530 B.n529 163.367
R1543 B.n529 B.n528 163.367
R1544 B.n528 B.n119 163.367
R1545 B.n524 B.n119 163.367
R1546 B.n524 B.n523 163.367
R1547 B.n523 B.n522 163.367
R1548 B.n522 B.n121 163.367
R1549 B.n518 B.n121 163.367
R1550 B.n518 B.n517 163.367
R1551 B.n517 B.n516 163.367
R1552 B.n516 B.n123 163.367
R1553 B.n512 B.n123 163.367
R1554 B.n512 B.n511 163.367
R1555 B.n511 B.n510 163.367
R1556 B.n510 B.n125 163.367
R1557 B.n506 B.n125 163.367
R1558 B.n506 B.n505 163.367
R1559 B.n505 B.n504 163.367
R1560 B.n504 B.n127 163.367
R1561 B.n500 B.n127 163.367
R1562 B.n500 B.n499 163.367
R1563 B.n499 B.n498 163.367
R1564 B.n498 B.n129 163.367
R1565 B.n494 B.n129 163.367
R1566 B.n494 B.n493 163.367
R1567 B.n493 B.n492 163.367
R1568 B.n492 B.n131 163.367
R1569 B.n488 B.n131 163.367
R1570 B.n488 B.n487 163.367
R1571 B.n487 B.n486 163.367
R1572 B.n486 B.n133 163.367
R1573 B.n482 B.n133 163.367
R1574 B.n482 B.n481 163.367
R1575 B.n481 B.n480 163.367
R1576 B.n480 B.n135 163.367
R1577 B.n476 B.n135 163.367
R1578 B.n476 B.n475 163.367
R1579 B.n475 B.n474 163.367
R1580 B.n474 B.n137 163.367
R1581 B.n470 B.n137 163.367
R1582 B.n470 B.n469 163.367
R1583 B.n469 B.n468 163.367
R1584 B.n468 B.n139 163.367
R1585 B.n464 B.n139 163.367
R1586 B.n464 B.n463 163.367
R1587 B.n463 B.n462 163.367
R1588 B.n462 B.n141 163.367
R1589 B.n458 B.n141 163.367
R1590 B.n458 B.n457 163.367
R1591 B.n457 B.n456 163.367
R1592 B.n456 B.n143 163.367
R1593 B.n452 B.n143 163.367
R1594 B.n452 B.n451 163.367
R1595 B.n451 B.n450 163.367
R1596 B.n450 B.n145 163.367
R1597 B.n446 B.n145 163.367
R1598 B.n446 B.n445 163.367
R1599 B.n445 B.n444 163.367
R1600 B.n444 B.n147 163.367
R1601 B.n440 B.n147 163.367
R1602 B.n440 B.n439 163.367
R1603 B.n760 B.n37 163.367
R1604 B.n760 B.n759 163.367
R1605 B.n759 B.n758 163.367
R1606 B.n758 B.n39 163.367
R1607 B.n754 B.n39 163.367
R1608 B.n754 B.n753 163.367
R1609 B.n753 B.n752 163.367
R1610 B.n752 B.n41 163.367
R1611 B.n748 B.n41 163.367
R1612 B.n748 B.n747 163.367
R1613 B.n747 B.n746 163.367
R1614 B.n746 B.n43 163.367
R1615 B.n742 B.n43 163.367
R1616 B.n742 B.n741 163.367
R1617 B.n741 B.n740 163.367
R1618 B.n740 B.n45 163.367
R1619 B.n736 B.n45 163.367
R1620 B.n736 B.n735 163.367
R1621 B.n735 B.n734 163.367
R1622 B.n734 B.n47 163.367
R1623 B.n730 B.n47 163.367
R1624 B.n730 B.n729 163.367
R1625 B.n729 B.n728 163.367
R1626 B.n728 B.n49 163.367
R1627 B.n724 B.n49 163.367
R1628 B.n724 B.n723 163.367
R1629 B.n723 B.n722 163.367
R1630 B.n722 B.n51 163.367
R1631 B.n718 B.n51 163.367
R1632 B.n718 B.n717 163.367
R1633 B.n717 B.n716 163.367
R1634 B.n716 B.n53 163.367
R1635 B.n711 B.n53 163.367
R1636 B.n711 B.n710 163.367
R1637 B.n710 B.n709 163.367
R1638 B.n709 B.n57 163.367
R1639 B.n705 B.n57 163.367
R1640 B.n705 B.n704 163.367
R1641 B.n704 B.n703 163.367
R1642 B.n703 B.n59 163.367
R1643 B.n698 B.n59 163.367
R1644 B.n698 B.n697 163.367
R1645 B.n697 B.n696 163.367
R1646 B.n696 B.n63 163.367
R1647 B.n692 B.n63 163.367
R1648 B.n692 B.n691 163.367
R1649 B.n691 B.n690 163.367
R1650 B.n690 B.n65 163.367
R1651 B.n686 B.n65 163.367
R1652 B.n686 B.n685 163.367
R1653 B.n685 B.n684 163.367
R1654 B.n684 B.n67 163.367
R1655 B.n680 B.n67 163.367
R1656 B.n680 B.n679 163.367
R1657 B.n679 B.n678 163.367
R1658 B.n678 B.n69 163.367
R1659 B.n674 B.n69 163.367
R1660 B.n674 B.n673 163.367
R1661 B.n673 B.n672 163.367
R1662 B.n672 B.n71 163.367
R1663 B.n668 B.n71 163.367
R1664 B.n668 B.n667 163.367
R1665 B.n667 B.n666 163.367
R1666 B.n666 B.n73 163.367
R1667 B.n662 B.n73 163.367
R1668 B.n662 B.n661 163.367
R1669 B.n661 B.n660 163.367
R1670 B.n660 B.n75 163.367
R1671 B.n656 B.n75 163.367
R1672 B.n656 B.n655 163.367
R1673 B.n655 B.n654 163.367
R1674 B.n654 B.n77 163.367
R1675 B.n765 B.n764 163.367
R1676 B.n766 B.n765 163.367
R1677 B.n766 B.n35 163.367
R1678 B.n770 B.n35 163.367
R1679 B.n771 B.n770 163.367
R1680 B.n772 B.n771 163.367
R1681 B.n772 B.n33 163.367
R1682 B.n776 B.n33 163.367
R1683 B.n777 B.n776 163.367
R1684 B.n778 B.n777 163.367
R1685 B.n778 B.n31 163.367
R1686 B.n782 B.n31 163.367
R1687 B.n783 B.n782 163.367
R1688 B.n784 B.n783 163.367
R1689 B.n784 B.n29 163.367
R1690 B.n788 B.n29 163.367
R1691 B.n789 B.n788 163.367
R1692 B.n790 B.n789 163.367
R1693 B.n790 B.n27 163.367
R1694 B.n794 B.n27 163.367
R1695 B.n795 B.n794 163.367
R1696 B.n796 B.n795 163.367
R1697 B.n796 B.n25 163.367
R1698 B.n800 B.n25 163.367
R1699 B.n801 B.n800 163.367
R1700 B.n802 B.n801 163.367
R1701 B.n802 B.n23 163.367
R1702 B.n806 B.n23 163.367
R1703 B.n807 B.n806 163.367
R1704 B.n808 B.n807 163.367
R1705 B.n808 B.n21 163.367
R1706 B.n812 B.n21 163.367
R1707 B.n813 B.n812 163.367
R1708 B.n814 B.n813 163.367
R1709 B.n814 B.n19 163.367
R1710 B.n818 B.n19 163.367
R1711 B.n819 B.n818 163.367
R1712 B.n820 B.n819 163.367
R1713 B.n820 B.n17 163.367
R1714 B.n824 B.n17 163.367
R1715 B.n825 B.n824 163.367
R1716 B.n826 B.n825 163.367
R1717 B.n826 B.n15 163.367
R1718 B.n830 B.n15 163.367
R1719 B.n831 B.n830 163.367
R1720 B.n832 B.n831 163.367
R1721 B.n832 B.n13 163.367
R1722 B.n836 B.n13 163.367
R1723 B.n837 B.n836 163.367
R1724 B.n838 B.n837 163.367
R1725 B.n838 B.n11 163.367
R1726 B.n842 B.n11 163.367
R1727 B.n843 B.n842 163.367
R1728 B.n844 B.n843 163.367
R1729 B.n844 B.n9 163.367
R1730 B.n848 B.n9 163.367
R1731 B.n849 B.n848 163.367
R1732 B.n850 B.n849 163.367
R1733 B.n850 B.n7 163.367
R1734 B.n854 B.n7 163.367
R1735 B.n855 B.n854 163.367
R1736 B.n856 B.n855 163.367
R1737 B.n856 B.n5 163.367
R1738 B.n860 B.n5 163.367
R1739 B.n861 B.n860 163.367
R1740 B.n862 B.n861 163.367
R1741 B.n862 B.n3 163.367
R1742 B.n866 B.n3 163.367
R1743 B.n867 B.n866 163.367
R1744 B.n221 B.n2 163.367
R1745 B.n224 B.n221 163.367
R1746 B.n225 B.n224 163.367
R1747 B.n226 B.n225 163.367
R1748 B.n226 B.n219 163.367
R1749 B.n230 B.n219 163.367
R1750 B.n231 B.n230 163.367
R1751 B.n232 B.n231 163.367
R1752 B.n232 B.n217 163.367
R1753 B.n236 B.n217 163.367
R1754 B.n237 B.n236 163.367
R1755 B.n238 B.n237 163.367
R1756 B.n238 B.n215 163.367
R1757 B.n242 B.n215 163.367
R1758 B.n243 B.n242 163.367
R1759 B.n244 B.n243 163.367
R1760 B.n244 B.n213 163.367
R1761 B.n248 B.n213 163.367
R1762 B.n249 B.n248 163.367
R1763 B.n250 B.n249 163.367
R1764 B.n250 B.n211 163.367
R1765 B.n254 B.n211 163.367
R1766 B.n255 B.n254 163.367
R1767 B.n256 B.n255 163.367
R1768 B.n256 B.n209 163.367
R1769 B.n260 B.n209 163.367
R1770 B.n261 B.n260 163.367
R1771 B.n262 B.n261 163.367
R1772 B.n262 B.n207 163.367
R1773 B.n266 B.n207 163.367
R1774 B.n267 B.n266 163.367
R1775 B.n268 B.n267 163.367
R1776 B.n268 B.n205 163.367
R1777 B.n272 B.n205 163.367
R1778 B.n273 B.n272 163.367
R1779 B.n274 B.n273 163.367
R1780 B.n274 B.n203 163.367
R1781 B.n278 B.n203 163.367
R1782 B.n279 B.n278 163.367
R1783 B.n280 B.n279 163.367
R1784 B.n280 B.n201 163.367
R1785 B.n284 B.n201 163.367
R1786 B.n285 B.n284 163.367
R1787 B.n286 B.n285 163.367
R1788 B.n286 B.n199 163.367
R1789 B.n290 B.n199 163.367
R1790 B.n291 B.n290 163.367
R1791 B.n292 B.n291 163.367
R1792 B.n292 B.n197 163.367
R1793 B.n296 B.n197 163.367
R1794 B.n297 B.n296 163.367
R1795 B.n298 B.n297 163.367
R1796 B.n298 B.n195 163.367
R1797 B.n302 B.n195 163.367
R1798 B.n303 B.n302 163.367
R1799 B.n304 B.n303 163.367
R1800 B.n304 B.n193 163.367
R1801 B.n308 B.n193 163.367
R1802 B.n309 B.n308 163.367
R1803 B.n310 B.n309 163.367
R1804 B.n310 B.n191 163.367
R1805 B.n314 B.n191 163.367
R1806 B.n315 B.n314 163.367
R1807 B.n316 B.n315 163.367
R1808 B.n316 B.n189 163.367
R1809 B.n320 B.n189 163.367
R1810 B.n321 B.n320 163.367
R1811 B.n322 B.n321 163.367
R1812 B.n322 B.n187 163.367
R1813 B.n171 B.n170 68.4611
R1814 B.n387 B.n386 68.4611
R1815 B.n61 B.n60 68.4611
R1816 B.n55 B.n54 68.4611
R1817 B.n373 B.n171 59.5399
R1818 B.n388 B.n387 59.5399
R1819 B.n700 B.n61 59.5399
R1820 B.n714 B.n55 59.5399
R1821 B.n763 B.n762 31.0639
R1822 B.n652 B.n651 31.0639
R1823 B.n437 B.n148 31.0639
R1824 B.n325 B.n324 31.0639
R1825 B B.n869 18.0485
R1826 B.n763 B.n36 10.6151
R1827 B.n767 B.n36 10.6151
R1828 B.n768 B.n767 10.6151
R1829 B.n769 B.n768 10.6151
R1830 B.n769 B.n34 10.6151
R1831 B.n773 B.n34 10.6151
R1832 B.n774 B.n773 10.6151
R1833 B.n775 B.n774 10.6151
R1834 B.n775 B.n32 10.6151
R1835 B.n779 B.n32 10.6151
R1836 B.n780 B.n779 10.6151
R1837 B.n781 B.n780 10.6151
R1838 B.n781 B.n30 10.6151
R1839 B.n785 B.n30 10.6151
R1840 B.n786 B.n785 10.6151
R1841 B.n787 B.n786 10.6151
R1842 B.n787 B.n28 10.6151
R1843 B.n791 B.n28 10.6151
R1844 B.n792 B.n791 10.6151
R1845 B.n793 B.n792 10.6151
R1846 B.n793 B.n26 10.6151
R1847 B.n797 B.n26 10.6151
R1848 B.n798 B.n797 10.6151
R1849 B.n799 B.n798 10.6151
R1850 B.n799 B.n24 10.6151
R1851 B.n803 B.n24 10.6151
R1852 B.n804 B.n803 10.6151
R1853 B.n805 B.n804 10.6151
R1854 B.n805 B.n22 10.6151
R1855 B.n809 B.n22 10.6151
R1856 B.n810 B.n809 10.6151
R1857 B.n811 B.n810 10.6151
R1858 B.n811 B.n20 10.6151
R1859 B.n815 B.n20 10.6151
R1860 B.n816 B.n815 10.6151
R1861 B.n817 B.n816 10.6151
R1862 B.n817 B.n18 10.6151
R1863 B.n821 B.n18 10.6151
R1864 B.n822 B.n821 10.6151
R1865 B.n823 B.n822 10.6151
R1866 B.n823 B.n16 10.6151
R1867 B.n827 B.n16 10.6151
R1868 B.n828 B.n827 10.6151
R1869 B.n829 B.n828 10.6151
R1870 B.n829 B.n14 10.6151
R1871 B.n833 B.n14 10.6151
R1872 B.n834 B.n833 10.6151
R1873 B.n835 B.n834 10.6151
R1874 B.n835 B.n12 10.6151
R1875 B.n839 B.n12 10.6151
R1876 B.n840 B.n839 10.6151
R1877 B.n841 B.n840 10.6151
R1878 B.n841 B.n10 10.6151
R1879 B.n845 B.n10 10.6151
R1880 B.n846 B.n845 10.6151
R1881 B.n847 B.n846 10.6151
R1882 B.n847 B.n8 10.6151
R1883 B.n851 B.n8 10.6151
R1884 B.n852 B.n851 10.6151
R1885 B.n853 B.n852 10.6151
R1886 B.n853 B.n6 10.6151
R1887 B.n857 B.n6 10.6151
R1888 B.n858 B.n857 10.6151
R1889 B.n859 B.n858 10.6151
R1890 B.n859 B.n4 10.6151
R1891 B.n863 B.n4 10.6151
R1892 B.n864 B.n863 10.6151
R1893 B.n865 B.n864 10.6151
R1894 B.n865 B.n0 10.6151
R1895 B.n762 B.n761 10.6151
R1896 B.n761 B.n38 10.6151
R1897 B.n757 B.n38 10.6151
R1898 B.n757 B.n756 10.6151
R1899 B.n756 B.n755 10.6151
R1900 B.n755 B.n40 10.6151
R1901 B.n751 B.n40 10.6151
R1902 B.n751 B.n750 10.6151
R1903 B.n750 B.n749 10.6151
R1904 B.n749 B.n42 10.6151
R1905 B.n745 B.n42 10.6151
R1906 B.n745 B.n744 10.6151
R1907 B.n744 B.n743 10.6151
R1908 B.n743 B.n44 10.6151
R1909 B.n739 B.n44 10.6151
R1910 B.n739 B.n738 10.6151
R1911 B.n738 B.n737 10.6151
R1912 B.n737 B.n46 10.6151
R1913 B.n733 B.n46 10.6151
R1914 B.n733 B.n732 10.6151
R1915 B.n732 B.n731 10.6151
R1916 B.n731 B.n48 10.6151
R1917 B.n727 B.n48 10.6151
R1918 B.n727 B.n726 10.6151
R1919 B.n726 B.n725 10.6151
R1920 B.n725 B.n50 10.6151
R1921 B.n721 B.n50 10.6151
R1922 B.n721 B.n720 10.6151
R1923 B.n720 B.n719 10.6151
R1924 B.n719 B.n52 10.6151
R1925 B.n715 B.n52 10.6151
R1926 B.n713 B.n712 10.6151
R1927 B.n712 B.n56 10.6151
R1928 B.n708 B.n56 10.6151
R1929 B.n708 B.n707 10.6151
R1930 B.n707 B.n706 10.6151
R1931 B.n706 B.n58 10.6151
R1932 B.n702 B.n58 10.6151
R1933 B.n702 B.n701 10.6151
R1934 B.n699 B.n62 10.6151
R1935 B.n695 B.n62 10.6151
R1936 B.n695 B.n694 10.6151
R1937 B.n694 B.n693 10.6151
R1938 B.n693 B.n64 10.6151
R1939 B.n689 B.n64 10.6151
R1940 B.n689 B.n688 10.6151
R1941 B.n688 B.n687 10.6151
R1942 B.n687 B.n66 10.6151
R1943 B.n683 B.n66 10.6151
R1944 B.n683 B.n682 10.6151
R1945 B.n682 B.n681 10.6151
R1946 B.n681 B.n68 10.6151
R1947 B.n677 B.n68 10.6151
R1948 B.n677 B.n676 10.6151
R1949 B.n676 B.n675 10.6151
R1950 B.n675 B.n70 10.6151
R1951 B.n671 B.n70 10.6151
R1952 B.n671 B.n670 10.6151
R1953 B.n670 B.n669 10.6151
R1954 B.n669 B.n72 10.6151
R1955 B.n665 B.n72 10.6151
R1956 B.n665 B.n664 10.6151
R1957 B.n664 B.n663 10.6151
R1958 B.n663 B.n74 10.6151
R1959 B.n659 B.n74 10.6151
R1960 B.n659 B.n658 10.6151
R1961 B.n658 B.n657 10.6151
R1962 B.n657 B.n76 10.6151
R1963 B.n653 B.n76 10.6151
R1964 B.n653 B.n652 10.6151
R1965 B.n651 B.n78 10.6151
R1966 B.n647 B.n78 10.6151
R1967 B.n647 B.n646 10.6151
R1968 B.n646 B.n645 10.6151
R1969 B.n645 B.n80 10.6151
R1970 B.n641 B.n80 10.6151
R1971 B.n641 B.n640 10.6151
R1972 B.n640 B.n639 10.6151
R1973 B.n639 B.n82 10.6151
R1974 B.n635 B.n82 10.6151
R1975 B.n635 B.n634 10.6151
R1976 B.n634 B.n633 10.6151
R1977 B.n633 B.n84 10.6151
R1978 B.n629 B.n84 10.6151
R1979 B.n629 B.n628 10.6151
R1980 B.n628 B.n627 10.6151
R1981 B.n627 B.n86 10.6151
R1982 B.n623 B.n86 10.6151
R1983 B.n623 B.n622 10.6151
R1984 B.n622 B.n621 10.6151
R1985 B.n621 B.n88 10.6151
R1986 B.n617 B.n88 10.6151
R1987 B.n617 B.n616 10.6151
R1988 B.n616 B.n615 10.6151
R1989 B.n615 B.n90 10.6151
R1990 B.n611 B.n90 10.6151
R1991 B.n611 B.n610 10.6151
R1992 B.n610 B.n609 10.6151
R1993 B.n609 B.n92 10.6151
R1994 B.n605 B.n92 10.6151
R1995 B.n605 B.n604 10.6151
R1996 B.n604 B.n603 10.6151
R1997 B.n603 B.n94 10.6151
R1998 B.n599 B.n94 10.6151
R1999 B.n599 B.n598 10.6151
R2000 B.n598 B.n597 10.6151
R2001 B.n597 B.n96 10.6151
R2002 B.n593 B.n96 10.6151
R2003 B.n593 B.n592 10.6151
R2004 B.n592 B.n591 10.6151
R2005 B.n591 B.n98 10.6151
R2006 B.n587 B.n98 10.6151
R2007 B.n587 B.n586 10.6151
R2008 B.n586 B.n585 10.6151
R2009 B.n585 B.n100 10.6151
R2010 B.n581 B.n100 10.6151
R2011 B.n581 B.n580 10.6151
R2012 B.n580 B.n579 10.6151
R2013 B.n579 B.n102 10.6151
R2014 B.n575 B.n102 10.6151
R2015 B.n575 B.n574 10.6151
R2016 B.n574 B.n573 10.6151
R2017 B.n573 B.n104 10.6151
R2018 B.n569 B.n104 10.6151
R2019 B.n569 B.n568 10.6151
R2020 B.n568 B.n567 10.6151
R2021 B.n567 B.n106 10.6151
R2022 B.n563 B.n106 10.6151
R2023 B.n563 B.n562 10.6151
R2024 B.n562 B.n561 10.6151
R2025 B.n561 B.n108 10.6151
R2026 B.n557 B.n108 10.6151
R2027 B.n557 B.n556 10.6151
R2028 B.n556 B.n555 10.6151
R2029 B.n555 B.n110 10.6151
R2030 B.n551 B.n110 10.6151
R2031 B.n551 B.n550 10.6151
R2032 B.n550 B.n549 10.6151
R2033 B.n549 B.n112 10.6151
R2034 B.n545 B.n112 10.6151
R2035 B.n545 B.n544 10.6151
R2036 B.n544 B.n543 10.6151
R2037 B.n543 B.n114 10.6151
R2038 B.n539 B.n114 10.6151
R2039 B.n539 B.n538 10.6151
R2040 B.n538 B.n537 10.6151
R2041 B.n537 B.n116 10.6151
R2042 B.n533 B.n116 10.6151
R2043 B.n533 B.n532 10.6151
R2044 B.n532 B.n531 10.6151
R2045 B.n531 B.n118 10.6151
R2046 B.n527 B.n118 10.6151
R2047 B.n527 B.n526 10.6151
R2048 B.n526 B.n525 10.6151
R2049 B.n525 B.n120 10.6151
R2050 B.n521 B.n120 10.6151
R2051 B.n521 B.n520 10.6151
R2052 B.n520 B.n519 10.6151
R2053 B.n519 B.n122 10.6151
R2054 B.n515 B.n122 10.6151
R2055 B.n515 B.n514 10.6151
R2056 B.n514 B.n513 10.6151
R2057 B.n513 B.n124 10.6151
R2058 B.n509 B.n124 10.6151
R2059 B.n509 B.n508 10.6151
R2060 B.n508 B.n507 10.6151
R2061 B.n507 B.n126 10.6151
R2062 B.n503 B.n126 10.6151
R2063 B.n503 B.n502 10.6151
R2064 B.n502 B.n501 10.6151
R2065 B.n501 B.n128 10.6151
R2066 B.n497 B.n128 10.6151
R2067 B.n497 B.n496 10.6151
R2068 B.n496 B.n495 10.6151
R2069 B.n495 B.n130 10.6151
R2070 B.n491 B.n130 10.6151
R2071 B.n491 B.n490 10.6151
R2072 B.n490 B.n489 10.6151
R2073 B.n489 B.n132 10.6151
R2074 B.n485 B.n132 10.6151
R2075 B.n485 B.n484 10.6151
R2076 B.n484 B.n483 10.6151
R2077 B.n483 B.n134 10.6151
R2078 B.n479 B.n134 10.6151
R2079 B.n479 B.n478 10.6151
R2080 B.n478 B.n477 10.6151
R2081 B.n477 B.n136 10.6151
R2082 B.n473 B.n136 10.6151
R2083 B.n473 B.n472 10.6151
R2084 B.n472 B.n471 10.6151
R2085 B.n471 B.n138 10.6151
R2086 B.n467 B.n138 10.6151
R2087 B.n467 B.n466 10.6151
R2088 B.n466 B.n465 10.6151
R2089 B.n465 B.n140 10.6151
R2090 B.n461 B.n140 10.6151
R2091 B.n461 B.n460 10.6151
R2092 B.n460 B.n459 10.6151
R2093 B.n459 B.n142 10.6151
R2094 B.n455 B.n142 10.6151
R2095 B.n455 B.n454 10.6151
R2096 B.n454 B.n453 10.6151
R2097 B.n453 B.n144 10.6151
R2098 B.n449 B.n144 10.6151
R2099 B.n449 B.n448 10.6151
R2100 B.n448 B.n447 10.6151
R2101 B.n447 B.n146 10.6151
R2102 B.n443 B.n146 10.6151
R2103 B.n443 B.n442 10.6151
R2104 B.n442 B.n441 10.6151
R2105 B.n441 B.n148 10.6151
R2106 B.n222 B.n1 10.6151
R2107 B.n223 B.n222 10.6151
R2108 B.n223 B.n220 10.6151
R2109 B.n227 B.n220 10.6151
R2110 B.n228 B.n227 10.6151
R2111 B.n229 B.n228 10.6151
R2112 B.n229 B.n218 10.6151
R2113 B.n233 B.n218 10.6151
R2114 B.n234 B.n233 10.6151
R2115 B.n235 B.n234 10.6151
R2116 B.n235 B.n216 10.6151
R2117 B.n239 B.n216 10.6151
R2118 B.n240 B.n239 10.6151
R2119 B.n241 B.n240 10.6151
R2120 B.n241 B.n214 10.6151
R2121 B.n245 B.n214 10.6151
R2122 B.n246 B.n245 10.6151
R2123 B.n247 B.n246 10.6151
R2124 B.n247 B.n212 10.6151
R2125 B.n251 B.n212 10.6151
R2126 B.n252 B.n251 10.6151
R2127 B.n253 B.n252 10.6151
R2128 B.n253 B.n210 10.6151
R2129 B.n257 B.n210 10.6151
R2130 B.n258 B.n257 10.6151
R2131 B.n259 B.n258 10.6151
R2132 B.n259 B.n208 10.6151
R2133 B.n263 B.n208 10.6151
R2134 B.n264 B.n263 10.6151
R2135 B.n265 B.n264 10.6151
R2136 B.n265 B.n206 10.6151
R2137 B.n269 B.n206 10.6151
R2138 B.n270 B.n269 10.6151
R2139 B.n271 B.n270 10.6151
R2140 B.n271 B.n204 10.6151
R2141 B.n275 B.n204 10.6151
R2142 B.n276 B.n275 10.6151
R2143 B.n277 B.n276 10.6151
R2144 B.n277 B.n202 10.6151
R2145 B.n281 B.n202 10.6151
R2146 B.n282 B.n281 10.6151
R2147 B.n283 B.n282 10.6151
R2148 B.n283 B.n200 10.6151
R2149 B.n287 B.n200 10.6151
R2150 B.n288 B.n287 10.6151
R2151 B.n289 B.n288 10.6151
R2152 B.n289 B.n198 10.6151
R2153 B.n293 B.n198 10.6151
R2154 B.n294 B.n293 10.6151
R2155 B.n295 B.n294 10.6151
R2156 B.n295 B.n196 10.6151
R2157 B.n299 B.n196 10.6151
R2158 B.n300 B.n299 10.6151
R2159 B.n301 B.n300 10.6151
R2160 B.n301 B.n194 10.6151
R2161 B.n305 B.n194 10.6151
R2162 B.n306 B.n305 10.6151
R2163 B.n307 B.n306 10.6151
R2164 B.n307 B.n192 10.6151
R2165 B.n311 B.n192 10.6151
R2166 B.n312 B.n311 10.6151
R2167 B.n313 B.n312 10.6151
R2168 B.n313 B.n190 10.6151
R2169 B.n317 B.n190 10.6151
R2170 B.n318 B.n317 10.6151
R2171 B.n319 B.n318 10.6151
R2172 B.n319 B.n188 10.6151
R2173 B.n323 B.n188 10.6151
R2174 B.n324 B.n323 10.6151
R2175 B.n325 B.n186 10.6151
R2176 B.n329 B.n186 10.6151
R2177 B.n330 B.n329 10.6151
R2178 B.n331 B.n330 10.6151
R2179 B.n331 B.n184 10.6151
R2180 B.n335 B.n184 10.6151
R2181 B.n336 B.n335 10.6151
R2182 B.n337 B.n336 10.6151
R2183 B.n337 B.n182 10.6151
R2184 B.n341 B.n182 10.6151
R2185 B.n342 B.n341 10.6151
R2186 B.n343 B.n342 10.6151
R2187 B.n343 B.n180 10.6151
R2188 B.n347 B.n180 10.6151
R2189 B.n348 B.n347 10.6151
R2190 B.n349 B.n348 10.6151
R2191 B.n349 B.n178 10.6151
R2192 B.n353 B.n178 10.6151
R2193 B.n354 B.n353 10.6151
R2194 B.n355 B.n354 10.6151
R2195 B.n355 B.n176 10.6151
R2196 B.n359 B.n176 10.6151
R2197 B.n360 B.n359 10.6151
R2198 B.n361 B.n360 10.6151
R2199 B.n361 B.n174 10.6151
R2200 B.n365 B.n174 10.6151
R2201 B.n366 B.n365 10.6151
R2202 B.n367 B.n366 10.6151
R2203 B.n367 B.n172 10.6151
R2204 B.n371 B.n172 10.6151
R2205 B.n372 B.n371 10.6151
R2206 B.n374 B.n168 10.6151
R2207 B.n378 B.n168 10.6151
R2208 B.n379 B.n378 10.6151
R2209 B.n380 B.n379 10.6151
R2210 B.n380 B.n166 10.6151
R2211 B.n384 B.n166 10.6151
R2212 B.n385 B.n384 10.6151
R2213 B.n389 B.n385 10.6151
R2214 B.n393 B.n164 10.6151
R2215 B.n394 B.n393 10.6151
R2216 B.n395 B.n394 10.6151
R2217 B.n395 B.n162 10.6151
R2218 B.n399 B.n162 10.6151
R2219 B.n400 B.n399 10.6151
R2220 B.n401 B.n400 10.6151
R2221 B.n401 B.n160 10.6151
R2222 B.n405 B.n160 10.6151
R2223 B.n406 B.n405 10.6151
R2224 B.n407 B.n406 10.6151
R2225 B.n407 B.n158 10.6151
R2226 B.n411 B.n158 10.6151
R2227 B.n412 B.n411 10.6151
R2228 B.n413 B.n412 10.6151
R2229 B.n413 B.n156 10.6151
R2230 B.n417 B.n156 10.6151
R2231 B.n418 B.n417 10.6151
R2232 B.n419 B.n418 10.6151
R2233 B.n419 B.n154 10.6151
R2234 B.n423 B.n154 10.6151
R2235 B.n424 B.n423 10.6151
R2236 B.n425 B.n424 10.6151
R2237 B.n425 B.n152 10.6151
R2238 B.n429 B.n152 10.6151
R2239 B.n430 B.n429 10.6151
R2240 B.n431 B.n430 10.6151
R2241 B.n431 B.n150 10.6151
R2242 B.n435 B.n150 10.6151
R2243 B.n436 B.n435 10.6151
R2244 B.n437 B.n436 10.6151
R2245 B.n869 B.n0 8.11757
R2246 B.n869 B.n1 8.11757
R2247 B.n714 B.n713 6.5566
R2248 B.n701 B.n700 6.5566
R2249 B.n374 B.n373 6.5566
R2250 B.n389 B.n388 6.5566
R2251 B.n715 B.n714 4.05904
R2252 B.n700 B.n699 4.05904
R2253 B.n373 B.n372 4.05904
R2254 B.n388 B.n164 4.05904
C0 VTAIL VDD1 9.21153f
C1 VDD1 w_n5206_n2692# 2.77881f
C2 VTAIL w_n5206_n2692# 2.82256f
C3 B VP 2.54674f
C4 VP VN 8.65149f
C5 B VN 1.40057f
C6 VDD2 VP 0.659908f
C7 VDD2 B 2.58526f
C8 VDD2 VN 8.11548f
C9 VDD1 VP 8.617249f
C10 VDD1 B 2.44398f
C11 VDD1 VN 0.15474f
C12 VTAIL VP 9.18591f
C13 w_n5206_n2692# VP 11.9318f
C14 VTAIL B 3.18184f
C15 w_n5206_n2692# B 10.6081f
C16 VTAIL VN 9.17171f
C17 w_n5206_n2692# VN 11.2521f
C18 VDD1 VDD2 2.56259f
C19 VTAIL VDD2 9.267691f
C20 VDD2 w_n5206_n2692# 2.95354f
C21 VDD2 VSUBS 2.345105f
C22 VDD1 VSUBS 2.128607f
C23 VTAIL VSUBS 1.342037f
C24 VN VSUBS 8.648041f
C25 VP VSUBS 4.887289f
C26 B VSUBS 5.826433f
C27 w_n5206_n2692# VSUBS 0.17361p
C28 B.n0 VSUBS 0.009005f
C29 B.n1 VSUBS 0.009005f
C30 B.n2 VSUBS 0.013318f
C31 B.n3 VSUBS 0.010206f
C32 B.n4 VSUBS 0.010206f
C33 B.n5 VSUBS 0.010206f
C34 B.n6 VSUBS 0.010206f
C35 B.n7 VSUBS 0.010206f
C36 B.n8 VSUBS 0.010206f
C37 B.n9 VSUBS 0.010206f
C38 B.n10 VSUBS 0.010206f
C39 B.n11 VSUBS 0.010206f
C40 B.n12 VSUBS 0.010206f
C41 B.n13 VSUBS 0.010206f
C42 B.n14 VSUBS 0.010206f
C43 B.n15 VSUBS 0.010206f
C44 B.n16 VSUBS 0.010206f
C45 B.n17 VSUBS 0.010206f
C46 B.n18 VSUBS 0.010206f
C47 B.n19 VSUBS 0.010206f
C48 B.n20 VSUBS 0.010206f
C49 B.n21 VSUBS 0.010206f
C50 B.n22 VSUBS 0.010206f
C51 B.n23 VSUBS 0.010206f
C52 B.n24 VSUBS 0.010206f
C53 B.n25 VSUBS 0.010206f
C54 B.n26 VSUBS 0.010206f
C55 B.n27 VSUBS 0.010206f
C56 B.n28 VSUBS 0.010206f
C57 B.n29 VSUBS 0.010206f
C58 B.n30 VSUBS 0.010206f
C59 B.n31 VSUBS 0.010206f
C60 B.n32 VSUBS 0.010206f
C61 B.n33 VSUBS 0.010206f
C62 B.n34 VSUBS 0.010206f
C63 B.n35 VSUBS 0.010206f
C64 B.n36 VSUBS 0.010206f
C65 B.n37 VSUBS 0.023654f
C66 B.n38 VSUBS 0.010206f
C67 B.n39 VSUBS 0.010206f
C68 B.n40 VSUBS 0.010206f
C69 B.n41 VSUBS 0.010206f
C70 B.n42 VSUBS 0.010206f
C71 B.n43 VSUBS 0.010206f
C72 B.n44 VSUBS 0.010206f
C73 B.n45 VSUBS 0.010206f
C74 B.n46 VSUBS 0.010206f
C75 B.n47 VSUBS 0.010206f
C76 B.n48 VSUBS 0.010206f
C77 B.n49 VSUBS 0.010206f
C78 B.n50 VSUBS 0.010206f
C79 B.n51 VSUBS 0.010206f
C80 B.n52 VSUBS 0.010206f
C81 B.n53 VSUBS 0.010206f
C82 B.t4 VSUBS 0.202499f
C83 B.t5 VSUBS 0.253099f
C84 B.t3 VSUBS 1.88938f
C85 B.n54 VSUBS 0.413297f
C86 B.n55 VSUBS 0.297779f
C87 B.n56 VSUBS 0.010206f
C88 B.n57 VSUBS 0.010206f
C89 B.n58 VSUBS 0.010206f
C90 B.n59 VSUBS 0.010206f
C91 B.t10 VSUBS 0.202502f
C92 B.t11 VSUBS 0.253102f
C93 B.t9 VSUBS 1.88938f
C94 B.n60 VSUBS 0.413294f
C95 B.n61 VSUBS 0.297776f
C96 B.n62 VSUBS 0.010206f
C97 B.n63 VSUBS 0.010206f
C98 B.n64 VSUBS 0.010206f
C99 B.n65 VSUBS 0.010206f
C100 B.n66 VSUBS 0.010206f
C101 B.n67 VSUBS 0.010206f
C102 B.n68 VSUBS 0.010206f
C103 B.n69 VSUBS 0.010206f
C104 B.n70 VSUBS 0.010206f
C105 B.n71 VSUBS 0.010206f
C106 B.n72 VSUBS 0.010206f
C107 B.n73 VSUBS 0.010206f
C108 B.n74 VSUBS 0.010206f
C109 B.n75 VSUBS 0.010206f
C110 B.n76 VSUBS 0.010206f
C111 B.n77 VSUBS 0.023654f
C112 B.n78 VSUBS 0.010206f
C113 B.n79 VSUBS 0.010206f
C114 B.n80 VSUBS 0.010206f
C115 B.n81 VSUBS 0.010206f
C116 B.n82 VSUBS 0.010206f
C117 B.n83 VSUBS 0.010206f
C118 B.n84 VSUBS 0.010206f
C119 B.n85 VSUBS 0.010206f
C120 B.n86 VSUBS 0.010206f
C121 B.n87 VSUBS 0.010206f
C122 B.n88 VSUBS 0.010206f
C123 B.n89 VSUBS 0.010206f
C124 B.n90 VSUBS 0.010206f
C125 B.n91 VSUBS 0.010206f
C126 B.n92 VSUBS 0.010206f
C127 B.n93 VSUBS 0.010206f
C128 B.n94 VSUBS 0.010206f
C129 B.n95 VSUBS 0.010206f
C130 B.n96 VSUBS 0.010206f
C131 B.n97 VSUBS 0.010206f
C132 B.n98 VSUBS 0.010206f
C133 B.n99 VSUBS 0.010206f
C134 B.n100 VSUBS 0.010206f
C135 B.n101 VSUBS 0.010206f
C136 B.n102 VSUBS 0.010206f
C137 B.n103 VSUBS 0.010206f
C138 B.n104 VSUBS 0.010206f
C139 B.n105 VSUBS 0.010206f
C140 B.n106 VSUBS 0.010206f
C141 B.n107 VSUBS 0.010206f
C142 B.n108 VSUBS 0.010206f
C143 B.n109 VSUBS 0.010206f
C144 B.n110 VSUBS 0.010206f
C145 B.n111 VSUBS 0.010206f
C146 B.n112 VSUBS 0.010206f
C147 B.n113 VSUBS 0.010206f
C148 B.n114 VSUBS 0.010206f
C149 B.n115 VSUBS 0.010206f
C150 B.n116 VSUBS 0.010206f
C151 B.n117 VSUBS 0.010206f
C152 B.n118 VSUBS 0.010206f
C153 B.n119 VSUBS 0.010206f
C154 B.n120 VSUBS 0.010206f
C155 B.n121 VSUBS 0.010206f
C156 B.n122 VSUBS 0.010206f
C157 B.n123 VSUBS 0.010206f
C158 B.n124 VSUBS 0.010206f
C159 B.n125 VSUBS 0.010206f
C160 B.n126 VSUBS 0.010206f
C161 B.n127 VSUBS 0.010206f
C162 B.n128 VSUBS 0.010206f
C163 B.n129 VSUBS 0.010206f
C164 B.n130 VSUBS 0.010206f
C165 B.n131 VSUBS 0.010206f
C166 B.n132 VSUBS 0.010206f
C167 B.n133 VSUBS 0.010206f
C168 B.n134 VSUBS 0.010206f
C169 B.n135 VSUBS 0.010206f
C170 B.n136 VSUBS 0.010206f
C171 B.n137 VSUBS 0.010206f
C172 B.n138 VSUBS 0.010206f
C173 B.n139 VSUBS 0.010206f
C174 B.n140 VSUBS 0.010206f
C175 B.n141 VSUBS 0.010206f
C176 B.n142 VSUBS 0.010206f
C177 B.n143 VSUBS 0.010206f
C178 B.n144 VSUBS 0.010206f
C179 B.n145 VSUBS 0.010206f
C180 B.n146 VSUBS 0.010206f
C181 B.n147 VSUBS 0.010206f
C182 B.n148 VSUBS 0.023839f
C183 B.n149 VSUBS 0.010206f
C184 B.n150 VSUBS 0.010206f
C185 B.n151 VSUBS 0.010206f
C186 B.n152 VSUBS 0.010206f
C187 B.n153 VSUBS 0.010206f
C188 B.n154 VSUBS 0.010206f
C189 B.n155 VSUBS 0.010206f
C190 B.n156 VSUBS 0.010206f
C191 B.n157 VSUBS 0.010206f
C192 B.n158 VSUBS 0.010206f
C193 B.n159 VSUBS 0.010206f
C194 B.n160 VSUBS 0.010206f
C195 B.n161 VSUBS 0.010206f
C196 B.n162 VSUBS 0.010206f
C197 B.n163 VSUBS 0.010206f
C198 B.n164 VSUBS 0.007054f
C199 B.n165 VSUBS 0.010206f
C200 B.n166 VSUBS 0.010206f
C201 B.n167 VSUBS 0.010206f
C202 B.n168 VSUBS 0.010206f
C203 B.n169 VSUBS 0.010206f
C204 B.t8 VSUBS 0.202499f
C205 B.t7 VSUBS 0.253099f
C206 B.t6 VSUBS 1.88938f
C207 B.n170 VSUBS 0.413297f
C208 B.n171 VSUBS 0.297779f
C209 B.n172 VSUBS 0.010206f
C210 B.n173 VSUBS 0.010206f
C211 B.n174 VSUBS 0.010206f
C212 B.n175 VSUBS 0.010206f
C213 B.n176 VSUBS 0.010206f
C214 B.n177 VSUBS 0.010206f
C215 B.n178 VSUBS 0.010206f
C216 B.n179 VSUBS 0.010206f
C217 B.n180 VSUBS 0.010206f
C218 B.n181 VSUBS 0.010206f
C219 B.n182 VSUBS 0.010206f
C220 B.n183 VSUBS 0.010206f
C221 B.n184 VSUBS 0.010206f
C222 B.n185 VSUBS 0.010206f
C223 B.n186 VSUBS 0.010206f
C224 B.n187 VSUBS 0.022572f
C225 B.n188 VSUBS 0.010206f
C226 B.n189 VSUBS 0.010206f
C227 B.n190 VSUBS 0.010206f
C228 B.n191 VSUBS 0.010206f
C229 B.n192 VSUBS 0.010206f
C230 B.n193 VSUBS 0.010206f
C231 B.n194 VSUBS 0.010206f
C232 B.n195 VSUBS 0.010206f
C233 B.n196 VSUBS 0.010206f
C234 B.n197 VSUBS 0.010206f
C235 B.n198 VSUBS 0.010206f
C236 B.n199 VSUBS 0.010206f
C237 B.n200 VSUBS 0.010206f
C238 B.n201 VSUBS 0.010206f
C239 B.n202 VSUBS 0.010206f
C240 B.n203 VSUBS 0.010206f
C241 B.n204 VSUBS 0.010206f
C242 B.n205 VSUBS 0.010206f
C243 B.n206 VSUBS 0.010206f
C244 B.n207 VSUBS 0.010206f
C245 B.n208 VSUBS 0.010206f
C246 B.n209 VSUBS 0.010206f
C247 B.n210 VSUBS 0.010206f
C248 B.n211 VSUBS 0.010206f
C249 B.n212 VSUBS 0.010206f
C250 B.n213 VSUBS 0.010206f
C251 B.n214 VSUBS 0.010206f
C252 B.n215 VSUBS 0.010206f
C253 B.n216 VSUBS 0.010206f
C254 B.n217 VSUBS 0.010206f
C255 B.n218 VSUBS 0.010206f
C256 B.n219 VSUBS 0.010206f
C257 B.n220 VSUBS 0.010206f
C258 B.n221 VSUBS 0.010206f
C259 B.n222 VSUBS 0.010206f
C260 B.n223 VSUBS 0.010206f
C261 B.n224 VSUBS 0.010206f
C262 B.n225 VSUBS 0.010206f
C263 B.n226 VSUBS 0.010206f
C264 B.n227 VSUBS 0.010206f
C265 B.n228 VSUBS 0.010206f
C266 B.n229 VSUBS 0.010206f
C267 B.n230 VSUBS 0.010206f
C268 B.n231 VSUBS 0.010206f
C269 B.n232 VSUBS 0.010206f
C270 B.n233 VSUBS 0.010206f
C271 B.n234 VSUBS 0.010206f
C272 B.n235 VSUBS 0.010206f
C273 B.n236 VSUBS 0.010206f
C274 B.n237 VSUBS 0.010206f
C275 B.n238 VSUBS 0.010206f
C276 B.n239 VSUBS 0.010206f
C277 B.n240 VSUBS 0.010206f
C278 B.n241 VSUBS 0.010206f
C279 B.n242 VSUBS 0.010206f
C280 B.n243 VSUBS 0.010206f
C281 B.n244 VSUBS 0.010206f
C282 B.n245 VSUBS 0.010206f
C283 B.n246 VSUBS 0.010206f
C284 B.n247 VSUBS 0.010206f
C285 B.n248 VSUBS 0.010206f
C286 B.n249 VSUBS 0.010206f
C287 B.n250 VSUBS 0.010206f
C288 B.n251 VSUBS 0.010206f
C289 B.n252 VSUBS 0.010206f
C290 B.n253 VSUBS 0.010206f
C291 B.n254 VSUBS 0.010206f
C292 B.n255 VSUBS 0.010206f
C293 B.n256 VSUBS 0.010206f
C294 B.n257 VSUBS 0.010206f
C295 B.n258 VSUBS 0.010206f
C296 B.n259 VSUBS 0.010206f
C297 B.n260 VSUBS 0.010206f
C298 B.n261 VSUBS 0.010206f
C299 B.n262 VSUBS 0.010206f
C300 B.n263 VSUBS 0.010206f
C301 B.n264 VSUBS 0.010206f
C302 B.n265 VSUBS 0.010206f
C303 B.n266 VSUBS 0.010206f
C304 B.n267 VSUBS 0.010206f
C305 B.n268 VSUBS 0.010206f
C306 B.n269 VSUBS 0.010206f
C307 B.n270 VSUBS 0.010206f
C308 B.n271 VSUBS 0.010206f
C309 B.n272 VSUBS 0.010206f
C310 B.n273 VSUBS 0.010206f
C311 B.n274 VSUBS 0.010206f
C312 B.n275 VSUBS 0.010206f
C313 B.n276 VSUBS 0.010206f
C314 B.n277 VSUBS 0.010206f
C315 B.n278 VSUBS 0.010206f
C316 B.n279 VSUBS 0.010206f
C317 B.n280 VSUBS 0.010206f
C318 B.n281 VSUBS 0.010206f
C319 B.n282 VSUBS 0.010206f
C320 B.n283 VSUBS 0.010206f
C321 B.n284 VSUBS 0.010206f
C322 B.n285 VSUBS 0.010206f
C323 B.n286 VSUBS 0.010206f
C324 B.n287 VSUBS 0.010206f
C325 B.n288 VSUBS 0.010206f
C326 B.n289 VSUBS 0.010206f
C327 B.n290 VSUBS 0.010206f
C328 B.n291 VSUBS 0.010206f
C329 B.n292 VSUBS 0.010206f
C330 B.n293 VSUBS 0.010206f
C331 B.n294 VSUBS 0.010206f
C332 B.n295 VSUBS 0.010206f
C333 B.n296 VSUBS 0.010206f
C334 B.n297 VSUBS 0.010206f
C335 B.n298 VSUBS 0.010206f
C336 B.n299 VSUBS 0.010206f
C337 B.n300 VSUBS 0.010206f
C338 B.n301 VSUBS 0.010206f
C339 B.n302 VSUBS 0.010206f
C340 B.n303 VSUBS 0.010206f
C341 B.n304 VSUBS 0.010206f
C342 B.n305 VSUBS 0.010206f
C343 B.n306 VSUBS 0.010206f
C344 B.n307 VSUBS 0.010206f
C345 B.n308 VSUBS 0.010206f
C346 B.n309 VSUBS 0.010206f
C347 B.n310 VSUBS 0.010206f
C348 B.n311 VSUBS 0.010206f
C349 B.n312 VSUBS 0.010206f
C350 B.n313 VSUBS 0.010206f
C351 B.n314 VSUBS 0.010206f
C352 B.n315 VSUBS 0.010206f
C353 B.n316 VSUBS 0.010206f
C354 B.n317 VSUBS 0.010206f
C355 B.n318 VSUBS 0.010206f
C356 B.n319 VSUBS 0.010206f
C357 B.n320 VSUBS 0.010206f
C358 B.n321 VSUBS 0.010206f
C359 B.n322 VSUBS 0.010206f
C360 B.n323 VSUBS 0.010206f
C361 B.n324 VSUBS 0.022572f
C362 B.n325 VSUBS 0.023654f
C363 B.n326 VSUBS 0.023654f
C364 B.n327 VSUBS 0.010206f
C365 B.n328 VSUBS 0.010206f
C366 B.n329 VSUBS 0.010206f
C367 B.n330 VSUBS 0.010206f
C368 B.n331 VSUBS 0.010206f
C369 B.n332 VSUBS 0.010206f
C370 B.n333 VSUBS 0.010206f
C371 B.n334 VSUBS 0.010206f
C372 B.n335 VSUBS 0.010206f
C373 B.n336 VSUBS 0.010206f
C374 B.n337 VSUBS 0.010206f
C375 B.n338 VSUBS 0.010206f
C376 B.n339 VSUBS 0.010206f
C377 B.n340 VSUBS 0.010206f
C378 B.n341 VSUBS 0.010206f
C379 B.n342 VSUBS 0.010206f
C380 B.n343 VSUBS 0.010206f
C381 B.n344 VSUBS 0.010206f
C382 B.n345 VSUBS 0.010206f
C383 B.n346 VSUBS 0.010206f
C384 B.n347 VSUBS 0.010206f
C385 B.n348 VSUBS 0.010206f
C386 B.n349 VSUBS 0.010206f
C387 B.n350 VSUBS 0.010206f
C388 B.n351 VSUBS 0.010206f
C389 B.n352 VSUBS 0.010206f
C390 B.n353 VSUBS 0.010206f
C391 B.n354 VSUBS 0.010206f
C392 B.n355 VSUBS 0.010206f
C393 B.n356 VSUBS 0.010206f
C394 B.n357 VSUBS 0.010206f
C395 B.n358 VSUBS 0.010206f
C396 B.n359 VSUBS 0.010206f
C397 B.n360 VSUBS 0.010206f
C398 B.n361 VSUBS 0.010206f
C399 B.n362 VSUBS 0.010206f
C400 B.n363 VSUBS 0.010206f
C401 B.n364 VSUBS 0.010206f
C402 B.n365 VSUBS 0.010206f
C403 B.n366 VSUBS 0.010206f
C404 B.n367 VSUBS 0.010206f
C405 B.n368 VSUBS 0.010206f
C406 B.n369 VSUBS 0.010206f
C407 B.n370 VSUBS 0.010206f
C408 B.n371 VSUBS 0.010206f
C409 B.n372 VSUBS 0.007054f
C410 B.n373 VSUBS 0.023645f
C411 B.n374 VSUBS 0.008255f
C412 B.n375 VSUBS 0.010206f
C413 B.n376 VSUBS 0.010206f
C414 B.n377 VSUBS 0.010206f
C415 B.n378 VSUBS 0.010206f
C416 B.n379 VSUBS 0.010206f
C417 B.n380 VSUBS 0.010206f
C418 B.n381 VSUBS 0.010206f
C419 B.n382 VSUBS 0.010206f
C420 B.n383 VSUBS 0.010206f
C421 B.n384 VSUBS 0.010206f
C422 B.n385 VSUBS 0.010206f
C423 B.t2 VSUBS 0.202502f
C424 B.t1 VSUBS 0.253102f
C425 B.t0 VSUBS 1.88938f
C426 B.n386 VSUBS 0.413294f
C427 B.n387 VSUBS 0.297776f
C428 B.n388 VSUBS 0.023645f
C429 B.n389 VSUBS 0.008255f
C430 B.n390 VSUBS 0.010206f
C431 B.n391 VSUBS 0.010206f
C432 B.n392 VSUBS 0.010206f
C433 B.n393 VSUBS 0.010206f
C434 B.n394 VSUBS 0.010206f
C435 B.n395 VSUBS 0.010206f
C436 B.n396 VSUBS 0.010206f
C437 B.n397 VSUBS 0.010206f
C438 B.n398 VSUBS 0.010206f
C439 B.n399 VSUBS 0.010206f
C440 B.n400 VSUBS 0.010206f
C441 B.n401 VSUBS 0.010206f
C442 B.n402 VSUBS 0.010206f
C443 B.n403 VSUBS 0.010206f
C444 B.n404 VSUBS 0.010206f
C445 B.n405 VSUBS 0.010206f
C446 B.n406 VSUBS 0.010206f
C447 B.n407 VSUBS 0.010206f
C448 B.n408 VSUBS 0.010206f
C449 B.n409 VSUBS 0.010206f
C450 B.n410 VSUBS 0.010206f
C451 B.n411 VSUBS 0.010206f
C452 B.n412 VSUBS 0.010206f
C453 B.n413 VSUBS 0.010206f
C454 B.n414 VSUBS 0.010206f
C455 B.n415 VSUBS 0.010206f
C456 B.n416 VSUBS 0.010206f
C457 B.n417 VSUBS 0.010206f
C458 B.n418 VSUBS 0.010206f
C459 B.n419 VSUBS 0.010206f
C460 B.n420 VSUBS 0.010206f
C461 B.n421 VSUBS 0.010206f
C462 B.n422 VSUBS 0.010206f
C463 B.n423 VSUBS 0.010206f
C464 B.n424 VSUBS 0.010206f
C465 B.n425 VSUBS 0.010206f
C466 B.n426 VSUBS 0.010206f
C467 B.n427 VSUBS 0.010206f
C468 B.n428 VSUBS 0.010206f
C469 B.n429 VSUBS 0.010206f
C470 B.n430 VSUBS 0.010206f
C471 B.n431 VSUBS 0.010206f
C472 B.n432 VSUBS 0.010206f
C473 B.n433 VSUBS 0.010206f
C474 B.n434 VSUBS 0.010206f
C475 B.n435 VSUBS 0.010206f
C476 B.n436 VSUBS 0.010206f
C477 B.n437 VSUBS 0.022386f
C478 B.n438 VSUBS 0.023654f
C479 B.n439 VSUBS 0.022572f
C480 B.n440 VSUBS 0.010206f
C481 B.n441 VSUBS 0.010206f
C482 B.n442 VSUBS 0.010206f
C483 B.n443 VSUBS 0.010206f
C484 B.n444 VSUBS 0.010206f
C485 B.n445 VSUBS 0.010206f
C486 B.n446 VSUBS 0.010206f
C487 B.n447 VSUBS 0.010206f
C488 B.n448 VSUBS 0.010206f
C489 B.n449 VSUBS 0.010206f
C490 B.n450 VSUBS 0.010206f
C491 B.n451 VSUBS 0.010206f
C492 B.n452 VSUBS 0.010206f
C493 B.n453 VSUBS 0.010206f
C494 B.n454 VSUBS 0.010206f
C495 B.n455 VSUBS 0.010206f
C496 B.n456 VSUBS 0.010206f
C497 B.n457 VSUBS 0.010206f
C498 B.n458 VSUBS 0.010206f
C499 B.n459 VSUBS 0.010206f
C500 B.n460 VSUBS 0.010206f
C501 B.n461 VSUBS 0.010206f
C502 B.n462 VSUBS 0.010206f
C503 B.n463 VSUBS 0.010206f
C504 B.n464 VSUBS 0.010206f
C505 B.n465 VSUBS 0.010206f
C506 B.n466 VSUBS 0.010206f
C507 B.n467 VSUBS 0.010206f
C508 B.n468 VSUBS 0.010206f
C509 B.n469 VSUBS 0.010206f
C510 B.n470 VSUBS 0.010206f
C511 B.n471 VSUBS 0.010206f
C512 B.n472 VSUBS 0.010206f
C513 B.n473 VSUBS 0.010206f
C514 B.n474 VSUBS 0.010206f
C515 B.n475 VSUBS 0.010206f
C516 B.n476 VSUBS 0.010206f
C517 B.n477 VSUBS 0.010206f
C518 B.n478 VSUBS 0.010206f
C519 B.n479 VSUBS 0.010206f
C520 B.n480 VSUBS 0.010206f
C521 B.n481 VSUBS 0.010206f
C522 B.n482 VSUBS 0.010206f
C523 B.n483 VSUBS 0.010206f
C524 B.n484 VSUBS 0.010206f
C525 B.n485 VSUBS 0.010206f
C526 B.n486 VSUBS 0.010206f
C527 B.n487 VSUBS 0.010206f
C528 B.n488 VSUBS 0.010206f
C529 B.n489 VSUBS 0.010206f
C530 B.n490 VSUBS 0.010206f
C531 B.n491 VSUBS 0.010206f
C532 B.n492 VSUBS 0.010206f
C533 B.n493 VSUBS 0.010206f
C534 B.n494 VSUBS 0.010206f
C535 B.n495 VSUBS 0.010206f
C536 B.n496 VSUBS 0.010206f
C537 B.n497 VSUBS 0.010206f
C538 B.n498 VSUBS 0.010206f
C539 B.n499 VSUBS 0.010206f
C540 B.n500 VSUBS 0.010206f
C541 B.n501 VSUBS 0.010206f
C542 B.n502 VSUBS 0.010206f
C543 B.n503 VSUBS 0.010206f
C544 B.n504 VSUBS 0.010206f
C545 B.n505 VSUBS 0.010206f
C546 B.n506 VSUBS 0.010206f
C547 B.n507 VSUBS 0.010206f
C548 B.n508 VSUBS 0.010206f
C549 B.n509 VSUBS 0.010206f
C550 B.n510 VSUBS 0.010206f
C551 B.n511 VSUBS 0.010206f
C552 B.n512 VSUBS 0.010206f
C553 B.n513 VSUBS 0.010206f
C554 B.n514 VSUBS 0.010206f
C555 B.n515 VSUBS 0.010206f
C556 B.n516 VSUBS 0.010206f
C557 B.n517 VSUBS 0.010206f
C558 B.n518 VSUBS 0.010206f
C559 B.n519 VSUBS 0.010206f
C560 B.n520 VSUBS 0.010206f
C561 B.n521 VSUBS 0.010206f
C562 B.n522 VSUBS 0.010206f
C563 B.n523 VSUBS 0.010206f
C564 B.n524 VSUBS 0.010206f
C565 B.n525 VSUBS 0.010206f
C566 B.n526 VSUBS 0.010206f
C567 B.n527 VSUBS 0.010206f
C568 B.n528 VSUBS 0.010206f
C569 B.n529 VSUBS 0.010206f
C570 B.n530 VSUBS 0.010206f
C571 B.n531 VSUBS 0.010206f
C572 B.n532 VSUBS 0.010206f
C573 B.n533 VSUBS 0.010206f
C574 B.n534 VSUBS 0.010206f
C575 B.n535 VSUBS 0.010206f
C576 B.n536 VSUBS 0.010206f
C577 B.n537 VSUBS 0.010206f
C578 B.n538 VSUBS 0.010206f
C579 B.n539 VSUBS 0.010206f
C580 B.n540 VSUBS 0.010206f
C581 B.n541 VSUBS 0.010206f
C582 B.n542 VSUBS 0.010206f
C583 B.n543 VSUBS 0.010206f
C584 B.n544 VSUBS 0.010206f
C585 B.n545 VSUBS 0.010206f
C586 B.n546 VSUBS 0.010206f
C587 B.n547 VSUBS 0.010206f
C588 B.n548 VSUBS 0.010206f
C589 B.n549 VSUBS 0.010206f
C590 B.n550 VSUBS 0.010206f
C591 B.n551 VSUBS 0.010206f
C592 B.n552 VSUBS 0.010206f
C593 B.n553 VSUBS 0.010206f
C594 B.n554 VSUBS 0.010206f
C595 B.n555 VSUBS 0.010206f
C596 B.n556 VSUBS 0.010206f
C597 B.n557 VSUBS 0.010206f
C598 B.n558 VSUBS 0.010206f
C599 B.n559 VSUBS 0.010206f
C600 B.n560 VSUBS 0.010206f
C601 B.n561 VSUBS 0.010206f
C602 B.n562 VSUBS 0.010206f
C603 B.n563 VSUBS 0.010206f
C604 B.n564 VSUBS 0.010206f
C605 B.n565 VSUBS 0.010206f
C606 B.n566 VSUBS 0.010206f
C607 B.n567 VSUBS 0.010206f
C608 B.n568 VSUBS 0.010206f
C609 B.n569 VSUBS 0.010206f
C610 B.n570 VSUBS 0.010206f
C611 B.n571 VSUBS 0.010206f
C612 B.n572 VSUBS 0.010206f
C613 B.n573 VSUBS 0.010206f
C614 B.n574 VSUBS 0.010206f
C615 B.n575 VSUBS 0.010206f
C616 B.n576 VSUBS 0.010206f
C617 B.n577 VSUBS 0.010206f
C618 B.n578 VSUBS 0.010206f
C619 B.n579 VSUBS 0.010206f
C620 B.n580 VSUBS 0.010206f
C621 B.n581 VSUBS 0.010206f
C622 B.n582 VSUBS 0.010206f
C623 B.n583 VSUBS 0.010206f
C624 B.n584 VSUBS 0.010206f
C625 B.n585 VSUBS 0.010206f
C626 B.n586 VSUBS 0.010206f
C627 B.n587 VSUBS 0.010206f
C628 B.n588 VSUBS 0.010206f
C629 B.n589 VSUBS 0.010206f
C630 B.n590 VSUBS 0.010206f
C631 B.n591 VSUBS 0.010206f
C632 B.n592 VSUBS 0.010206f
C633 B.n593 VSUBS 0.010206f
C634 B.n594 VSUBS 0.010206f
C635 B.n595 VSUBS 0.010206f
C636 B.n596 VSUBS 0.010206f
C637 B.n597 VSUBS 0.010206f
C638 B.n598 VSUBS 0.010206f
C639 B.n599 VSUBS 0.010206f
C640 B.n600 VSUBS 0.010206f
C641 B.n601 VSUBS 0.010206f
C642 B.n602 VSUBS 0.010206f
C643 B.n603 VSUBS 0.010206f
C644 B.n604 VSUBS 0.010206f
C645 B.n605 VSUBS 0.010206f
C646 B.n606 VSUBS 0.010206f
C647 B.n607 VSUBS 0.010206f
C648 B.n608 VSUBS 0.010206f
C649 B.n609 VSUBS 0.010206f
C650 B.n610 VSUBS 0.010206f
C651 B.n611 VSUBS 0.010206f
C652 B.n612 VSUBS 0.010206f
C653 B.n613 VSUBS 0.010206f
C654 B.n614 VSUBS 0.010206f
C655 B.n615 VSUBS 0.010206f
C656 B.n616 VSUBS 0.010206f
C657 B.n617 VSUBS 0.010206f
C658 B.n618 VSUBS 0.010206f
C659 B.n619 VSUBS 0.010206f
C660 B.n620 VSUBS 0.010206f
C661 B.n621 VSUBS 0.010206f
C662 B.n622 VSUBS 0.010206f
C663 B.n623 VSUBS 0.010206f
C664 B.n624 VSUBS 0.010206f
C665 B.n625 VSUBS 0.010206f
C666 B.n626 VSUBS 0.010206f
C667 B.n627 VSUBS 0.010206f
C668 B.n628 VSUBS 0.010206f
C669 B.n629 VSUBS 0.010206f
C670 B.n630 VSUBS 0.010206f
C671 B.n631 VSUBS 0.010206f
C672 B.n632 VSUBS 0.010206f
C673 B.n633 VSUBS 0.010206f
C674 B.n634 VSUBS 0.010206f
C675 B.n635 VSUBS 0.010206f
C676 B.n636 VSUBS 0.010206f
C677 B.n637 VSUBS 0.010206f
C678 B.n638 VSUBS 0.010206f
C679 B.n639 VSUBS 0.010206f
C680 B.n640 VSUBS 0.010206f
C681 B.n641 VSUBS 0.010206f
C682 B.n642 VSUBS 0.010206f
C683 B.n643 VSUBS 0.010206f
C684 B.n644 VSUBS 0.010206f
C685 B.n645 VSUBS 0.010206f
C686 B.n646 VSUBS 0.010206f
C687 B.n647 VSUBS 0.010206f
C688 B.n648 VSUBS 0.010206f
C689 B.n649 VSUBS 0.010206f
C690 B.n650 VSUBS 0.022572f
C691 B.n651 VSUBS 0.022572f
C692 B.n652 VSUBS 0.023654f
C693 B.n653 VSUBS 0.010206f
C694 B.n654 VSUBS 0.010206f
C695 B.n655 VSUBS 0.010206f
C696 B.n656 VSUBS 0.010206f
C697 B.n657 VSUBS 0.010206f
C698 B.n658 VSUBS 0.010206f
C699 B.n659 VSUBS 0.010206f
C700 B.n660 VSUBS 0.010206f
C701 B.n661 VSUBS 0.010206f
C702 B.n662 VSUBS 0.010206f
C703 B.n663 VSUBS 0.010206f
C704 B.n664 VSUBS 0.010206f
C705 B.n665 VSUBS 0.010206f
C706 B.n666 VSUBS 0.010206f
C707 B.n667 VSUBS 0.010206f
C708 B.n668 VSUBS 0.010206f
C709 B.n669 VSUBS 0.010206f
C710 B.n670 VSUBS 0.010206f
C711 B.n671 VSUBS 0.010206f
C712 B.n672 VSUBS 0.010206f
C713 B.n673 VSUBS 0.010206f
C714 B.n674 VSUBS 0.010206f
C715 B.n675 VSUBS 0.010206f
C716 B.n676 VSUBS 0.010206f
C717 B.n677 VSUBS 0.010206f
C718 B.n678 VSUBS 0.010206f
C719 B.n679 VSUBS 0.010206f
C720 B.n680 VSUBS 0.010206f
C721 B.n681 VSUBS 0.010206f
C722 B.n682 VSUBS 0.010206f
C723 B.n683 VSUBS 0.010206f
C724 B.n684 VSUBS 0.010206f
C725 B.n685 VSUBS 0.010206f
C726 B.n686 VSUBS 0.010206f
C727 B.n687 VSUBS 0.010206f
C728 B.n688 VSUBS 0.010206f
C729 B.n689 VSUBS 0.010206f
C730 B.n690 VSUBS 0.010206f
C731 B.n691 VSUBS 0.010206f
C732 B.n692 VSUBS 0.010206f
C733 B.n693 VSUBS 0.010206f
C734 B.n694 VSUBS 0.010206f
C735 B.n695 VSUBS 0.010206f
C736 B.n696 VSUBS 0.010206f
C737 B.n697 VSUBS 0.010206f
C738 B.n698 VSUBS 0.010206f
C739 B.n699 VSUBS 0.007054f
C740 B.n700 VSUBS 0.023645f
C741 B.n701 VSUBS 0.008255f
C742 B.n702 VSUBS 0.010206f
C743 B.n703 VSUBS 0.010206f
C744 B.n704 VSUBS 0.010206f
C745 B.n705 VSUBS 0.010206f
C746 B.n706 VSUBS 0.010206f
C747 B.n707 VSUBS 0.010206f
C748 B.n708 VSUBS 0.010206f
C749 B.n709 VSUBS 0.010206f
C750 B.n710 VSUBS 0.010206f
C751 B.n711 VSUBS 0.010206f
C752 B.n712 VSUBS 0.010206f
C753 B.n713 VSUBS 0.008255f
C754 B.n714 VSUBS 0.023645f
C755 B.n715 VSUBS 0.007054f
C756 B.n716 VSUBS 0.010206f
C757 B.n717 VSUBS 0.010206f
C758 B.n718 VSUBS 0.010206f
C759 B.n719 VSUBS 0.010206f
C760 B.n720 VSUBS 0.010206f
C761 B.n721 VSUBS 0.010206f
C762 B.n722 VSUBS 0.010206f
C763 B.n723 VSUBS 0.010206f
C764 B.n724 VSUBS 0.010206f
C765 B.n725 VSUBS 0.010206f
C766 B.n726 VSUBS 0.010206f
C767 B.n727 VSUBS 0.010206f
C768 B.n728 VSUBS 0.010206f
C769 B.n729 VSUBS 0.010206f
C770 B.n730 VSUBS 0.010206f
C771 B.n731 VSUBS 0.010206f
C772 B.n732 VSUBS 0.010206f
C773 B.n733 VSUBS 0.010206f
C774 B.n734 VSUBS 0.010206f
C775 B.n735 VSUBS 0.010206f
C776 B.n736 VSUBS 0.010206f
C777 B.n737 VSUBS 0.010206f
C778 B.n738 VSUBS 0.010206f
C779 B.n739 VSUBS 0.010206f
C780 B.n740 VSUBS 0.010206f
C781 B.n741 VSUBS 0.010206f
C782 B.n742 VSUBS 0.010206f
C783 B.n743 VSUBS 0.010206f
C784 B.n744 VSUBS 0.010206f
C785 B.n745 VSUBS 0.010206f
C786 B.n746 VSUBS 0.010206f
C787 B.n747 VSUBS 0.010206f
C788 B.n748 VSUBS 0.010206f
C789 B.n749 VSUBS 0.010206f
C790 B.n750 VSUBS 0.010206f
C791 B.n751 VSUBS 0.010206f
C792 B.n752 VSUBS 0.010206f
C793 B.n753 VSUBS 0.010206f
C794 B.n754 VSUBS 0.010206f
C795 B.n755 VSUBS 0.010206f
C796 B.n756 VSUBS 0.010206f
C797 B.n757 VSUBS 0.010206f
C798 B.n758 VSUBS 0.010206f
C799 B.n759 VSUBS 0.010206f
C800 B.n760 VSUBS 0.010206f
C801 B.n761 VSUBS 0.010206f
C802 B.n762 VSUBS 0.023654f
C803 B.n763 VSUBS 0.022572f
C804 B.n764 VSUBS 0.022572f
C805 B.n765 VSUBS 0.010206f
C806 B.n766 VSUBS 0.010206f
C807 B.n767 VSUBS 0.010206f
C808 B.n768 VSUBS 0.010206f
C809 B.n769 VSUBS 0.010206f
C810 B.n770 VSUBS 0.010206f
C811 B.n771 VSUBS 0.010206f
C812 B.n772 VSUBS 0.010206f
C813 B.n773 VSUBS 0.010206f
C814 B.n774 VSUBS 0.010206f
C815 B.n775 VSUBS 0.010206f
C816 B.n776 VSUBS 0.010206f
C817 B.n777 VSUBS 0.010206f
C818 B.n778 VSUBS 0.010206f
C819 B.n779 VSUBS 0.010206f
C820 B.n780 VSUBS 0.010206f
C821 B.n781 VSUBS 0.010206f
C822 B.n782 VSUBS 0.010206f
C823 B.n783 VSUBS 0.010206f
C824 B.n784 VSUBS 0.010206f
C825 B.n785 VSUBS 0.010206f
C826 B.n786 VSUBS 0.010206f
C827 B.n787 VSUBS 0.010206f
C828 B.n788 VSUBS 0.010206f
C829 B.n789 VSUBS 0.010206f
C830 B.n790 VSUBS 0.010206f
C831 B.n791 VSUBS 0.010206f
C832 B.n792 VSUBS 0.010206f
C833 B.n793 VSUBS 0.010206f
C834 B.n794 VSUBS 0.010206f
C835 B.n795 VSUBS 0.010206f
C836 B.n796 VSUBS 0.010206f
C837 B.n797 VSUBS 0.010206f
C838 B.n798 VSUBS 0.010206f
C839 B.n799 VSUBS 0.010206f
C840 B.n800 VSUBS 0.010206f
C841 B.n801 VSUBS 0.010206f
C842 B.n802 VSUBS 0.010206f
C843 B.n803 VSUBS 0.010206f
C844 B.n804 VSUBS 0.010206f
C845 B.n805 VSUBS 0.010206f
C846 B.n806 VSUBS 0.010206f
C847 B.n807 VSUBS 0.010206f
C848 B.n808 VSUBS 0.010206f
C849 B.n809 VSUBS 0.010206f
C850 B.n810 VSUBS 0.010206f
C851 B.n811 VSUBS 0.010206f
C852 B.n812 VSUBS 0.010206f
C853 B.n813 VSUBS 0.010206f
C854 B.n814 VSUBS 0.010206f
C855 B.n815 VSUBS 0.010206f
C856 B.n816 VSUBS 0.010206f
C857 B.n817 VSUBS 0.010206f
C858 B.n818 VSUBS 0.010206f
C859 B.n819 VSUBS 0.010206f
C860 B.n820 VSUBS 0.010206f
C861 B.n821 VSUBS 0.010206f
C862 B.n822 VSUBS 0.010206f
C863 B.n823 VSUBS 0.010206f
C864 B.n824 VSUBS 0.010206f
C865 B.n825 VSUBS 0.010206f
C866 B.n826 VSUBS 0.010206f
C867 B.n827 VSUBS 0.010206f
C868 B.n828 VSUBS 0.010206f
C869 B.n829 VSUBS 0.010206f
C870 B.n830 VSUBS 0.010206f
C871 B.n831 VSUBS 0.010206f
C872 B.n832 VSUBS 0.010206f
C873 B.n833 VSUBS 0.010206f
C874 B.n834 VSUBS 0.010206f
C875 B.n835 VSUBS 0.010206f
C876 B.n836 VSUBS 0.010206f
C877 B.n837 VSUBS 0.010206f
C878 B.n838 VSUBS 0.010206f
C879 B.n839 VSUBS 0.010206f
C880 B.n840 VSUBS 0.010206f
C881 B.n841 VSUBS 0.010206f
C882 B.n842 VSUBS 0.010206f
C883 B.n843 VSUBS 0.010206f
C884 B.n844 VSUBS 0.010206f
C885 B.n845 VSUBS 0.010206f
C886 B.n846 VSUBS 0.010206f
C887 B.n847 VSUBS 0.010206f
C888 B.n848 VSUBS 0.010206f
C889 B.n849 VSUBS 0.010206f
C890 B.n850 VSUBS 0.010206f
C891 B.n851 VSUBS 0.010206f
C892 B.n852 VSUBS 0.010206f
C893 B.n853 VSUBS 0.010206f
C894 B.n854 VSUBS 0.010206f
C895 B.n855 VSUBS 0.010206f
C896 B.n856 VSUBS 0.010206f
C897 B.n857 VSUBS 0.010206f
C898 B.n858 VSUBS 0.010206f
C899 B.n859 VSUBS 0.010206f
C900 B.n860 VSUBS 0.010206f
C901 B.n861 VSUBS 0.010206f
C902 B.n862 VSUBS 0.010206f
C903 B.n863 VSUBS 0.010206f
C904 B.n864 VSUBS 0.010206f
C905 B.n865 VSUBS 0.010206f
C906 B.n866 VSUBS 0.010206f
C907 B.n867 VSUBS 0.013318f
C908 B.n868 VSUBS 0.014187f
C909 B.n869 VSUBS 0.028212f
C910 VDD2.n0 VSUBS 0.034368f
C911 VDD2.n1 VSUBS 0.032662f
C912 VDD2.n2 VSUBS 0.017551f
C913 VDD2.n3 VSUBS 0.041485f
C914 VDD2.n4 VSUBS 0.018584f
C915 VDD2.n5 VSUBS 0.032662f
C916 VDD2.n6 VSUBS 0.017551f
C917 VDD2.n7 VSUBS 0.041485f
C918 VDD2.n8 VSUBS 0.018584f
C919 VDD2.n9 VSUBS 0.032662f
C920 VDD2.n10 VSUBS 0.017551f
C921 VDD2.n11 VSUBS 0.041485f
C922 VDD2.n12 VSUBS 0.018584f
C923 VDD2.n13 VSUBS 0.207387f
C924 VDD2.t2 VSUBS 0.089106f
C925 VDD2.n14 VSUBS 0.031113f
C926 VDD2.n15 VSUBS 0.031207f
C927 VDD2.n16 VSUBS 0.017551f
C928 VDD2.n17 VSUBS 1.12091f
C929 VDD2.n18 VSUBS 0.032662f
C930 VDD2.n19 VSUBS 0.017551f
C931 VDD2.n20 VSUBS 0.018584f
C932 VDD2.n21 VSUBS 0.041485f
C933 VDD2.n22 VSUBS 0.041485f
C934 VDD2.n23 VSUBS 0.018584f
C935 VDD2.n24 VSUBS 0.017551f
C936 VDD2.n25 VSUBS 0.032662f
C937 VDD2.n26 VSUBS 0.032662f
C938 VDD2.n27 VSUBS 0.017551f
C939 VDD2.n28 VSUBS 0.018584f
C940 VDD2.n29 VSUBS 0.041485f
C941 VDD2.n30 VSUBS 0.041485f
C942 VDD2.n31 VSUBS 0.041485f
C943 VDD2.n32 VSUBS 0.018584f
C944 VDD2.n33 VSUBS 0.017551f
C945 VDD2.n34 VSUBS 0.032662f
C946 VDD2.n35 VSUBS 0.032662f
C947 VDD2.n36 VSUBS 0.017551f
C948 VDD2.n37 VSUBS 0.018067f
C949 VDD2.n38 VSUBS 0.018067f
C950 VDD2.n39 VSUBS 0.041485f
C951 VDD2.n40 VSUBS 0.095248f
C952 VDD2.n41 VSUBS 0.018584f
C953 VDD2.n42 VSUBS 0.017551f
C954 VDD2.n43 VSUBS 0.079959f
C955 VDD2.n44 VSUBS 0.092121f
C956 VDD2.t0 VSUBS 0.222487f
C957 VDD2.t7 VSUBS 0.222487f
C958 VDD2.n45 VSUBS 1.63663f
C959 VDD2.n46 VSUBS 1.32298f
C960 VDD2.t1 VSUBS 0.222487f
C961 VDD2.t6 VSUBS 0.222487f
C962 VDD2.n47 VSUBS 1.66646f
C963 VDD2.n48 VSUBS 4.22545f
C964 VDD2.n49 VSUBS 0.034368f
C965 VDD2.n50 VSUBS 0.032662f
C966 VDD2.n51 VSUBS 0.017551f
C967 VDD2.n52 VSUBS 0.041485f
C968 VDD2.n53 VSUBS 0.018584f
C969 VDD2.n54 VSUBS 0.032662f
C970 VDD2.n55 VSUBS 0.017551f
C971 VDD2.n56 VSUBS 0.041485f
C972 VDD2.n57 VSUBS 0.041485f
C973 VDD2.n58 VSUBS 0.018584f
C974 VDD2.n59 VSUBS 0.032662f
C975 VDD2.n60 VSUBS 0.017551f
C976 VDD2.n61 VSUBS 0.041485f
C977 VDD2.n62 VSUBS 0.018584f
C978 VDD2.n63 VSUBS 0.207387f
C979 VDD2.t8 VSUBS 0.089106f
C980 VDD2.n64 VSUBS 0.031113f
C981 VDD2.n65 VSUBS 0.031207f
C982 VDD2.n66 VSUBS 0.017551f
C983 VDD2.n67 VSUBS 1.12091f
C984 VDD2.n68 VSUBS 0.032662f
C985 VDD2.n69 VSUBS 0.017551f
C986 VDD2.n70 VSUBS 0.018584f
C987 VDD2.n71 VSUBS 0.041485f
C988 VDD2.n72 VSUBS 0.041485f
C989 VDD2.n73 VSUBS 0.018584f
C990 VDD2.n74 VSUBS 0.017551f
C991 VDD2.n75 VSUBS 0.032662f
C992 VDD2.n76 VSUBS 0.032662f
C993 VDD2.n77 VSUBS 0.017551f
C994 VDD2.n78 VSUBS 0.018584f
C995 VDD2.n79 VSUBS 0.041485f
C996 VDD2.n80 VSUBS 0.041485f
C997 VDD2.n81 VSUBS 0.018584f
C998 VDD2.n82 VSUBS 0.017551f
C999 VDD2.n83 VSUBS 0.032662f
C1000 VDD2.n84 VSUBS 0.032662f
C1001 VDD2.n85 VSUBS 0.017551f
C1002 VDD2.n86 VSUBS 0.018067f
C1003 VDD2.n87 VSUBS 0.018067f
C1004 VDD2.n88 VSUBS 0.041485f
C1005 VDD2.n89 VSUBS 0.095248f
C1006 VDD2.n90 VSUBS 0.018584f
C1007 VDD2.n91 VSUBS 0.017551f
C1008 VDD2.n92 VSUBS 0.079959f
C1009 VDD2.n93 VSUBS 0.070322f
C1010 VDD2.n94 VSUBS 3.74315f
C1011 VDD2.t9 VSUBS 0.222487f
C1012 VDD2.t3 VSUBS 0.222487f
C1013 VDD2.n95 VSUBS 1.63664f
C1014 VDD2.n96 VSUBS 0.969929f
C1015 VDD2.t4 VSUBS 0.222487f
C1016 VDD2.t5 VSUBS 0.222487f
C1017 VDD2.n97 VSUBS 1.66641f
C1018 VN.t3 VSUBS 2.11365f
C1019 VN.n0 VSUBS 0.867932f
C1020 VN.n1 VSUBS 0.028442f
C1021 VN.n2 VSUBS 0.023715f
C1022 VN.n3 VSUBS 0.028442f
C1023 VN.t8 VSUBS 2.11365f
C1024 VN.n4 VSUBS 0.758928f
C1025 VN.n5 VSUBS 0.028442f
C1026 VN.n6 VSUBS 0.023053f
C1027 VN.n7 VSUBS 0.028442f
C1028 VN.t2 VSUBS 2.11365f
C1029 VN.n8 VSUBS 0.758928f
C1030 VN.n9 VSUBS 0.028442f
C1031 VN.n10 VSUBS 0.023053f
C1032 VN.n11 VSUBS 0.028442f
C1033 VN.t9 VSUBS 2.11365f
C1034 VN.n12 VSUBS 0.853381f
C1035 VN.t7 VSUBS 2.43719f
C1036 VN.n13 VSUBS 0.80974f
C1037 VN.n14 VSUBS 0.33035f
C1038 VN.n15 VSUBS 0.041287f
C1039 VN.n16 VSUBS 0.052743f
C1040 VN.n17 VSUBS 0.055768f
C1041 VN.n18 VSUBS 0.028442f
C1042 VN.n19 VSUBS 0.028442f
C1043 VN.n20 VSUBS 0.028442f
C1044 VN.n21 VSUBS 0.056612f
C1045 VN.n22 VSUBS 0.052743f
C1046 VN.n23 VSUBS 0.039724f
C1047 VN.n24 VSUBS 0.028442f
C1048 VN.n25 VSUBS 0.028442f
C1049 VN.n26 VSUBS 0.039724f
C1050 VN.n27 VSUBS 0.052743f
C1051 VN.n28 VSUBS 0.056612f
C1052 VN.n29 VSUBS 0.028442f
C1053 VN.n30 VSUBS 0.028442f
C1054 VN.n31 VSUBS 0.028442f
C1055 VN.n32 VSUBS 0.055768f
C1056 VN.n33 VSUBS 0.052743f
C1057 VN.n34 VSUBS 0.041287f
C1058 VN.n35 VSUBS 0.028442f
C1059 VN.n36 VSUBS 0.028442f
C1060 VN.n37 VSUBS 0.038162f
C1061 VN.n38 VSUBS 0.052743f
C1062 VN.n39 VSUBS 0.057089f
C1063 VN.n40 VSUBS 0.028442f
C1064 VN.n41 VSUBS 0.028442f
C1065 VN.n42 VSUBS 0.028442f
C1066 VN.n43 VSUBS 0.054629f
C1067 VN.n44 VSUBS 0.052743f
C1068 VN.n45 VSUBS 0.042849f
C1069 VN.n46 VSUBS 0.045898f
C1070 VN.n47 VSUBS 0.067048f
C1071 VN.t1 VSUBS 2.11365f
C1072 VN.n48 VSUBS 0.867932f
C1073 VN.n49 VSUBS 0.028442f
C1074 VN.n50 VSUBS 0.023715f
C1075 VN.n51 VSUBS 0.028442f
C1076 VN.t0 VSUBS 2.11365f
C1077 VN.n52 VSUBS 0.758928f
C1078 VN.n53 VSUBS 0.028442f
C1079 VN.n54 VSUBS 0.023053f
C1080 VN.n55 VSUBS 0.028442f
C1081 VN.t6 VSUBS 2.11365f
C1082 VN.n56 VSUBS 0.758928f
C1083 VN.n57 VSUBS 0.028442f
C1084 VN.n58 VSUBS 0.023053f
C1085 VN.n59 VSUBS 0.028442f
C1086 VN.t5 VSUBS 2.11365f
C1087 VN.n60 VSUBS 0.853381f
C1088 VN.t4 VSUBS 2.43719f
C1089 VN.n61 VSUBS 0.80974f
C1090 VN.n62 VSUBS 0.33035f
C1091 VN.n63 VSUBS 0.041287f
C1092 VN.n64 VSUBS 0.052743f
C1093 VN.n65 VSUBS 0.055768f
C1094 VN.n66 VSUBS 0.028442f
C1095 VN.n67 VSUBS 0.028442f
C1096 VN.n68 VSUBS 0.028442f
C1097 VN.n69 VSUBS 0.056612f
C1098 VN.n70 VSUBS 0.052743f
C1099 VN.n71 VSUBS 0.039724f
C1100 VN.n72 VSUBS 0.028442f
C1101 VN.n73 VSUBS 0.028442f
C1102 VN.n74 VSUBS 0.039724f
C1103 VN.n75 VSUBS 0.052743f
C1104 VN.n76 VSUBS 0.056612f
C1105 VN.n77 VSUBS 0.028442f
C1106 VN.n78 VSUBS 0.028442f
C1107 VN.n79 VSUBS 0.028442f
C1108 VN.n80 VSUBS 0.055768f
C1109 VN.n81 VSUBS 0.052743f
C1110 VN.n82 VSUBS 0.041287f
C1111 VN.n83 VSUBS 0.028442f
C1112 VN.n84 VSUBS 0.028442f
C1113 VN.n85 VSUBS 0.038162f
C1114 VN.n86 VSUBS 0.052743f
C1115 VN.n87 VSUBS 0.057089f
C1116 VN.n88 VSUBS 0.028442f
C1117 VN.n89 VSUBS 0.028442f
C1118 VN.n90 VSUBS 0.028442f
C1119 VN.n91 VSUBS 0.054629f
C1120 VN.n92 VSUBS 0.052743f
C1121 VN.n93 VSUBS 0.042849f
C1122 VN.n94 VSUBS 0.045898f
C1123 VN.n95 VSUBS 1.80872f
C1124 VDD1.n0 VSUBS 0.034206f
C1125 VDD1.n1 VSUBS 0.032509f
C1126 VDD1.n2 VSUBS 0.017469f
C1127 VDD1.n3 VSUBS 0.04129f
C1128 VDD1.n4 VSUBS 0.018496f
C1129 VDD1.n5 VSUBS 0.032509f
C1130 VDD1.n6 VSUBS 0.017469f
C1131 VDD1.n7 VSUBS 0.04129f
C1132 VDD1.n8 VSUBS 0.04129f
C1133 VDD1.n9 VSUBS 0.018496f
C1134 VDD1.n10 VSUBS 0.032509f
C1135 VDD1.n11 VSUBS 0.017469f
C1136 VDD1.n12 VSUBS 0.04129f
C1137 VDD1.n13 VSUBS 0.018496f
C1138 VDD1.n14 VSUBS 0.206414f
C1139 VDD1.t2 VSUBS 0.088688f
C1140 VDD1.n15 VSUBS 0.030968f
C1141 VDD1.n16 VSUBS 0.03106f
C1142 VDD1.n17 VSUBS 0.017469f
C1143 VDD1.n18 VSUBS 1.11566f
C1144 VDD1.n19 VSUBS 0.032509f
C1145 VDD1.n20 VSUBS 0.017469f
C1146 VDD1.n21 VSUBS 0.018496f
C1147 VDD1.n22 VSUBS 0.04129f
C1148 VDD1.n23 VSUBS 0.04129f
C1149 VDD1.n24 VSUBS 0.018496f
C1150 VDD1.n25 VSUBS 0.017469f
C1151 VDD1.n26 VSUBS 0.032509f
C1152 VDD1.n27 VSUBS 0.032509f
C1153 VDD1.n28 VSUBS 0.017469f
C1154 VDD1.n29 VSUBS 0.018496f
C1155 VDD1.n30 VSUBS 0.04129f
C1156 VDD1.n31 VSUBS 0.04129f
C1157 VDD1.n32 VSUBS 0.018496f
C1158 VDD1.n33 VSUBS 0.017469f
C1159 VDD1.n34 VSUBS 0.032509f
C1160 VDD1.n35 VSUBS 0.032509f
C1161 VDD1.n36 VSUBS 0.017469f
C1162 VDD1.n37 VSUBS 0.017983f
C1163 VDD1.n38 VSUBS 0.017983f
C1164 VDD1.n39 VSUBS 0.04129f
C1165 VDD1.n40 VSUBS 0.094802f
C1166 VDD1.n41 VSUBS 0.018496f
C1167 VDD1.n42 VSUBS 0.017469f
C1168 VDD1.n43 VSUBS 0.079584f
C1169 VDD1.n44 VSUBS 0.091689f
C1170 VDD1.t3 VSUBS 0.221443f
C1171 VDD1.t7 VSUBS 0.221443f
C1172 VDD1.n45 VSUBS 1.62896f
C1173 VDD1.n46 VSUBS 1.32759f
C1174 VDD1.n47 VSUBS 0.034206f
C1175 VDD1.n48 VSUBS 0.032509f
C1176 VDD1.n49 VSUBS 0.017469f
C1177 VDD1.n50 VSUBS 0.04129f
C1178 VDD1.n51 VSUBS 0.018496f
C1179 VDD1.n52 VSUBS 0.032509f
C1180 VDD1.n53 VSUBS 0.017469f
C1181 VDD1.n54 VSUBS 0.04129f
C1182 VDD1.n55 VSUBS 0.018496f
C1183 VDD1.n56 VSUBS 0.032509f
C1184 VDD1.n57 VSUBS 0.017469f
C1185 VDD1.n58 VSUBS 0.04129f
C1186 VDD1.n59 VSUBS 0.018496f
C1187 VDD1.n60 VSUBS 0.206414f
C1188 VDD1.t6 VSUBS 0.088688f
C1189 VDD1.n61 VSUBS 0.030968f
C1190 VDD1.n62 VSUBS 0.03106f
C1191 VDD1.n63 VSUBS 0.017469f
C1192 VDD1.n64 VSUBS 1.11566f
C1193 VDD1.n65 VSUBS 0.032509f
C1194 VDD1.n66 VSUBS 0.017469f
C1195 VDD1.n67 VSUBS 0.018496f
C1196 VDD1.n68 VSUBS 0.04129f
C1197 VDD1.n69 VSUBS 0.04129f
C1198 VDD1.n70 VSUBS 0.018496f
C1199 VDD1.n71 VSUBS 0.017469f
C1200 VDD1.n72 VSUBS 0.032509f
C1201 VDD1.n73 VSUBS 0.032509f
C1202 VDD1.n74 VSUBS 0.017469f
C1203 VDD1.n75 VSUBS 0.018496f
C1204 VDD1.n76 VSUBS 0.04129f
C1205 VDD1.n77 VSUBS 0.04129f
C1206 VDD1.n78 VSUBS 0.04129f
C1207 VDD1.n79 VSUBS 0.018496f
C1208 VDD1.n80 VSUBS 0.017469f
C1209 VDD1.n81 VSUBS 0.032509f
C1210 VDD1.n82 VSUBS 0.032509f
C1211 VDD1.n83 VSUBS 0.017469f
C1212 VDD1.n84 VSUBS 0.017983f
C1213 VDD1.n85 VSUBS 0.017983f
C1214 VDD1.n86 VSUBS 0.04129f
C1215 VDD1.n87 VSUBS 0.094802f
C1216 VDD1.n88 VSUBS 0.018496f
C1217 VDD1.n89 VSUBS 0.017469f
C1218 VDD1.n90 VSUBS 0.079584f
C1219 VDD1.n91 VSUBS 0.091689f
C1220 VDD1.t1 VSUBS 0.221443f
C1221 VDD1.t4 VSUBS 0.221443f
C1222 VDD1.n92 VSUBS 1.62895f
C1223 VDD1.n93 VSUBS 1.31678f
C1224 VDD1.t5 VSUBS 0.221443f
C1225 VDD1.t0 VSUBS 0.221443f
C1226 VDD1.n94 VSUBS 1.65865f
C1227 VDD1.n95 VSUBS 4.38592f
C1228 VDD1.t8 VSUBS 0.221443f
C1229 VDD1.t9 VSUBS 0.221443f
C1230 VDD1.n96 VSUBS 1.62895f
C1231 VDD1.n97 VSUBS 4.40714f
C1232 VTAIL.t9 VSUBS 0.213802f
C1233 VTAIL.t8 VSUBS 0.213802f
C1234 VTAIL.n0 VSUBS 1.43651f
C1235 VTAIL.n1 VSUBS 1.07315f
C1236 VTAIL.n2 VSUBS 0.033026f
C1237 VTAIL.n3 VSUBS 0.031387f
C1238 VTAIL.n4 VSUBS 0.016866f
C1239 VTAIL.n5 VSUBS 0.039865f
C1240 VTAIL.n6 VSUBS 0.017858f
C1241 VTAIL.n7 VSUBS 0.031387f
C1242 VTAIL.n8 VSUBS 0.016866f
C1243 VTAIL.n9 VSUBS 0.039865f
C1244 VTAIL.n10 VSUBS 0.017858f
C1245 VTAIL.n11 VSUBS 0.031387f
C1246 VTAIL.n12 VSUBS 0.016866f
C1247 VTAIL.n13 VSUBS 0.039865f
C1248 VTAIL.n14 VSUBS 0.017858f
C1249 VTAIL.n15 VSUBS 0.199291f
C1250 VTAIL.t17 VSUBS 0.085628f
C1251 VTAIL.n16 VSUBS 0.029899f
C1252 VTAIL.n17 VSUBS 0.029988f
C1253 VTAIL.n18 VSUBS 0.016866f
C1254 VTAIL.n19 VSUBS 1.07716f
C1255 VTAIL.n20 VSUBS 0.031387f
C1256 VTAIL.n21 VSUBS 0.016866f
C1257 VTAIL.n22 VSUBS 0.017858f
C1258 VTAIL.n23 VSUBS 0.039865f
C1259 VTAIL.n24 VSUBS 0.039865f
C1260 VTAIL.n25 VSUBS 0.017858f
C1261 VTAIL.n26 VSUBS 0.016866f
C1262 VTAIL.n27 VSUBS 0.031387f
C1263 VTAIL.n28 VSUBS 0.031387f
C1264 VTAIL.n29 VSUBS 0.016866f
C1265 VTAIL.n30 VSUBS 0.017858f
C1266 VTAIL.n31 VSUBS 0.039865f
C1267 VTAIL.n32 VSUBS 0.039865f
C1268 VTAIL.n33 VSUBS 0.039865f
C1269 VTAIL.n34 VSUBS 0.017858f
C1270 VTAIL.n35 VSUBS 0.016866f
C1271 VTAIL.n36 VSUBS 0.031387f
C1272 VTAIL.n37 VSUBS 0.031387f
C1273 VTAIL.n38 VSUBS 0.016866f
C1274 VTAIL.n39 VSUBS 0.017362f
C1275 VTAIL.n40 VSUBS 0.017362f
C1276 VTAIL.n41 VSUBS 0.039865f
C1277 VTAIL.n42 VSUBS 0.09153f
C1278 VTAIL.n43 VSUBS 0.017858f
C1279 VTAIL.n44 VSUBS 0.016866f
C1280 VTAIL.n45 VSUBS 0.076837f
C1281 VTAIL.n46 VSUBS 0.045937f
C1282 VTAIL.n47 VSUBS 0.538398f
C1283 VTAIL.t13 VSUBS 0.213802f
C1284 VTAIL.t12 VSUBS 0.213802f
C1285 VTAIL.n48 VSUBS 1.43651f
C1286 VTAIL.n49 VSUBS 1.25058f
C1287 VTAIL.t10 VSUBS 0.213802f
C1288 VTAIL.t18 VSUBS 0.213802f
C1289 VTAIL.n50 VSUBS 1.43651f
C1290 VTAIL.n51 VSUBS 2.73625f
C1291 VTAIL.t4 VSUBS 0.213802f
C1292 VTAIL.t6 VSUBS 0.213802f
C1293 VTAIL.n52 VSUBS 1.43652f
C1294 VTAIL.n53 VSUBS 2.73624f
C1295 VTAIL.t5 VSUBS 0.213802f
C1296 VTAIL.t2 VSUBS 0.213802f
C1297 VTAIL.n54 VSUBS 1.43652f
C1298 VTAIL.n55 VSUBS 1.25057f
C1299 VTAIL.n56 VSUBS 0.033026f
C1300 VTAIL.n57 VSUBS 0.031387f
C1301 VTAIL.n58 VSUBS 0.016866f
C1302 VTAIL.n59 VSUBS 0.039865f
C1303 VTAIL.n60 VSUBS 0.017858f
C1304 VTAIL.n61 VSUBS 0.031387f
C1305 VTAIL.n62 VSUBS 0.016866f
C1306 VTAIL.n63 VSUBS 0.039865f
C1307 VTAIL.n64 VSUBS 0.039865f
C1308 VTAIL.n65 VSUBS 0.017858f
C1309 VTAIL.n66 VSUBS 0.031387f
C1310 VTAIL.n67 VSUBS 0.016866f
C1311 VTAIL.n68 VSUBS 0.039865f
C1312 VTAIL.n69 VSUBS 0.017858f
C1313 VTAIL.n70 VSUBS 0.199291f
C1314 VTAIL.t0 VSUBS 0.085628f
C1315 VTAIL.n71 VSUBS 0.029899f
C1316 VTAIL.n72 VSUBS 0.029988f
C1317 VTAIL.n73 VSUBS 0.016866f
C1318 VTAIL.n74 VSUBS 1.07716f
C1319 VTAIL.n75 VSUBS 0.031387f
C1320 VTAIL.n76 VSUBS 0.016866f
C1321 VTAIL.n77 VSUBS 0.017858f
C1322 VTAIL.n78 VSUBS 0.039865f
C1323 VTAIL.n79 VSUBS 0.039865f
C1324 VTAIL.n80 VSUBS 0.017858f
C1325 VTAIL.n81 VSUBS 0.016866f
C1326 VTAIL.n82 VSUBS 0.031387f
C1327 VTAIL.n83 VSUBS 0.031387f
C1328 VTAIL.n84 VSUBS 0.016866f
C1329 VTAIL.n85 VSUBS 0.017858f
C1330 VTAIL.n86 VSUBS 0.039865f
C1331 VTAIL.n87 VSUBS 0.039865f
C1332 VTAIL.n88 VSUBS 0.017858f
C1333 VTAIL.n89 VSUBS 0.016866f
C1334 VTAIL.n90 VSUBS 0.031387f
C1335 VTAIL.n91 VSUBS 0.031387f
C1336 VTAIL.n92 VSUBS 0.016866f
C1337 VTAIL.n93 VSUBS 0.017362f
C1338 VTAIL.n94 VSUBS 0.017362f
C1339 VTAIL.n95 VSUBS 0.039865f
C1340 VTAIL.n96 VSUBS 0.09153f
C1341 VTAIL.n97 VSUBS 0.017858f
C1342 VTAIL.n98 VSUBS 0.016866f
C1343 VTAIL.n99 VSUBS 0.076837f
C1344 VTAIL.n100 VSUBS 0.045937f
C1345 VTAIL.n101 VSUBS 0.538398f
C1346 VTAIL.t19 VSUBS 0.213802f
C1347 VTAIL.t15 VSUBS 0.213802f
C1348 VTAIL.n102 VSUBS 1.43652f
C1349 VTAIL.n103 VSUBS 1.1442f
C1350 VTAIL.t11 VSUBS 0.213802f
C1351 VTAIL.t14 VSUBS 0.213802f
C1352 VTAIL.n104 VSUBS 1.43652f
C1353 VTAIL.n105 VSUBS 1.25057f
C1354 VTAIL.n106 VSUBS 0.033026f
C1355 VTAIL.n107 VSUBS 0.031387f
C1356 VTAIL.n108 VSUBS 0.016866f
C1357 VTAIL.n109 VSUBS 0.039865f
C1358 VTAIL.n110 VSUBS 0.017858f
C1359 VTAIL.n111 VSUBS 0.031387f
C1360 VTAIL.n112 VSUBS 0.016866f
C1361 VTAIL.n113 VSUBS 0.039865f
C1362 VTAIL.n114 VSUBS 0.039865f
C1363 VTAIL.n115 VSUBS 0.017858f
C1364 VTAIL.n116 VSUBS 0.031387f
C1365 VTAIL.n117 VSUBS 0.016866f
C1366 VTAIL.n118 VSUBS 0.039865f
C1367 VTAIL.n119 VSUBS 0.017858f
C1368 VTAIL.n120 VSUBS 0.199291f
C1369 VTAIL.t16 VSUBS 0.085628f
C1370 VTAIL.n121 VSUBS 0.029899f
C1371 VTAIL.n122 VSUBS 0.029988f
C1372 VTAIL.n123 VSUBS 0.016866f
C1373 VTAIL.n124 VSUBS 1.07716f
C1374 VTAIL.n125 VSUBS 0.031387f
C1375 VTAIL.n126 VSUBS 0.016866f
C1376 VTAIL.n127 VSUBS 0.017858f
C1377 VTAIL.n128 VSUBS 0.039865f
C1378 VTAIL.n129 VSUBS 0.039865f
C1379 VTAIL.n130 VSUBS 0.017858f
C1380 VTAIL.n131 VSUBS 0.016866f
C1381 VTAIL.n132 VSUBS 0.031387f
C1382 VTAIL.n133 VSUBS 0.031387f
C1383 VTAIL.n134 VSUBS 0.016866f
C1384 VTAIL.n135 VSUBS 0.017858f
C1385 VTAIL.n136 VSUBS 0.039865f
C1386 VTAIL.n137 VSUBS 0.039865f
C1387 VTAIL.n138 VSUBS 0.017858f
C1388 VTAIL.n139 VSUBS 0.016866f
C1389 VTAIL.n140 VSUBS 0.031387f
C1390 VTAIL.n141 VSUBS 0.031387f
C1391 VTAIL.n142 VSUBS 0.016866f
C1392 VTAIL.n143 VSUBS 0.017362f
C1393 VTAIL.n144 VSUBS 0.017362f
C1394 VTAIL.n145 VSUBS 0.039865f
C1395 VTAIL.n146 VSUBS 0.09153f
C1396 VTAIL.n147 VSUBS 0.017858f
C1397 VTAIL.n148 VSUBS 0.016866f
C1398 VTAIL.n149 VSUBS 0.076837f
C1399 VTAIL.n150 VSUBS 0.045937f
C1400 VTAIL.n151 VSUBS 1.82267f
C1401 VTAIL.n152 VSUBS 0.033026f
C1402 VTAIL.n153 VSUBS 0.031387f
C1403 VTAIL.n154 VSUBS 0.016866f
C1404 VTAIL.n155 VSUBS 0.039865f
C1405 VTAIL.n156 VSUBS 0.017858f
C1406 VTAIL.n157 VSUBS 0.031387f
C1407 VTAIL.n158 VSUBS 0.016866f
C1408 VTAIL.n159 VSUBS 0.039865f
C1409 VTAIL.n160 VSUBS 0.017858f
C1410 VTAIL.n161 VSUBS 0.031387f
C1411 VTAIL.n162 VSUBS 0.016866f
C1412 VTAIL.n163 VSUBS 0.039865f
C1413 VTAIL.n164 VSUBS 0.017858f
C1414 VTAIL.n165 VSUBS 0.199291f
C1415 VTAIL.t1 VSUBS 0.085628f
C1416 VTAIL.n166 VSUBS 0.029899f
C1417 VTAIL.n167 VSUBS 0.029988f
C1418 VTAIL.n168 VSUBS 0.016866f
C1419 VTAIL.n169 VSUBS 1.07716f
C1420 VTAIL.n170 VSUBS 0.031387f
C1421 VTAIL.n171 VSUBS 0.016866f
C1422 VTAIL.n172 VSUBS 0.017858f
C1423 VTAIL.n173 VSUBS 0.039865f
C1424 VTAIL.n174 VSUBS 0.039865f
C1425 VTAIL.n175 VSUBS 0.017858f
C1426 VTAIL.n176 VSUBS 0.016866f
C1427 VTAIL.n177 VSUBS 0.031387f
C1428 VTAIL.n178 VSUBS 0.031387f
C1429 VTAIL.n179 VSUBS 0.016866f
C1430 VTAIL.n180 VSUBS 0.017858f
C1431 VTAIL.n181 VSUBS 0.039865f
C1432 VTAIL.n182 VSUBS 0.039865f
C1433 VTAIL.n183 VSUBS 0.039865f
C1434 VTAIL.n184 VSUBS 0.017858f
C1435 VTAIL.n185 VSUBS 0.016866f
C1436 VTAIL.n186 VSUBS 0.031387f
C1437 VTAIL.n187 VSUBS 0.031387f
C1438 VTAIL.n188 VSUBS 0.016866f
C1439 VTAIL.n189 VSUBS 0.017362f
C1440 VTAIL.n190 VSUBS 0.017362f
C1441 VTAIL.n191 VSUBS 0.039865f
C1442 VTAIL.n192 VSUBS 0.09153f
C1443 VTAIL.n193 VSUBS 0.017858f
C1444 VTAIL.n194 VSUBS 0.016866f
C1445 VTAIL.n195 VSUBS 0.076837f
C1446 VTAIL.n196 VSUBS 0.045937f
C1447 VTAIL.n197 VSUBS 1.82267f
C1448 VTAIL.t3 VSUBS 0.213802f
C1449 VTAIL.t7 VSUBS 0.213802f
C1450 VTAIL.n198 VSUBS 1.43651f
C1451 VTAIL.n199 VSUBS 1.01387f
C1452 VP.t9 VSUBS 2.32013f
C1453 VP.n0 VSUBS 0.952721f
C1454 VP.n1 VSUBS 0.031221f
C1455 VP.n2 VSUBS 0.026031f
C1456 VP.n3 VSUBS 0.031221f
C1457 VP.t4 VSUBS 2.32013f
C1458 VP.n4 VSUBS 0.833068f
C1459 VP.n5 VSUBS 0.031221f
C1460 VP.n6 VSUBS 0.025306f
C1461 VP.n7 VSUBS 0.031221f
C1462 VP.t5 VSUBS 2.32013f
C1463 VP.n8 VSUBS 0.833068f
C1464 VP.n9 VSUBS 0.031221f
C1465 VP.n10 VSUBS 0.025306f
C1466 VP.n11 VSUBS 0.031221f
C1467 VP.t8 VSUBS 2.32013f
C1468 VP.n12 VSUBS 0.833068f
C1469 VP.n13 VSUBS 0.031221f
C1470 VP.n14 VSUBS 0.026031f
C1471 VP.n15 VSUBS 0.031221f
C1472 VP.t3 VSUBS 2.32013f
C1473 VP.n16 VSUBS 0.952721f
C1474 VP.t0 VSUBS 2.32013f
C1475 VP.n17 VSUBS 0.952721f
C1476 VP.n18 VSUBS 0.031221f
C1477 VP.n19 VSUBS 0.026031f
C1478 VP.n20 VSUBS 0.031221f
C1479 VP.t1 VSUBS 2.32013f
C1480 VP.n21 VSUBS 0.833068f
C1481 VP.n22 VSUBS 0.031221f
C1482 VP.n23 VSUBS 0.025306f
C1483 VP.n24 VSUBS 0.031221f
C1484 VP.t2 VSUBS 2.32013f
C1485 VP.n25 VSUBS 0.833068f
C1486 VP.n26 VSUBS 0.031221f
C1487 VP.n27 VSUBS 0.025306f
C1488 VP.n28 VSUBS 0.031221f
C1489 VP.t6 VSUBS 2.32013f
C1490 VP.n29 VSUBS 0.936749f
C1491 VP.t7 VSUBS 2.67528f
C1492 VP.n30 VSUBS 0.888845f
C1493 VP.n31 VSUBS 0.362622f
C1494 VP.n32 VSUBS 0.04532f
C1495 VP.n33 VSUBS 0.057896f
C1496 VP.n34 VSUBS 0.061216f
C1497 VP.n35 VSUBS 0.031221f
C1498 VP.n36 VSUBS 0.031221f
C1499 VP.n37 VSUBS 0.031221f
C1500 VP.n38 VSUBS 0.062142f
C1501 VP.n39 VSUBS 0.057896f
C1502 VP.n40 VSUBS 0.043605f
C1503 VP.n41 VSUBS 0.031221f
C1504 VP.n42 VSUBS 0.031221f
C1505 VP.n43 VSUBS 0.043605f
C1506 VP.n44 VSUBS 0.057896f
C1507 VP.n45 VSUBS 0.062142f
C1508 VP.n46 VSUBS 0.031221f
C1509 VP.n47 VSUBS 0.031221f
C1510 VP.n48 VSUBS 0.031221f
C1511 VP.n49 VSUBS 0.061216f
C1512 VP.n50 VSUBS 0.057896f
C1513 VP.n51 VSUBS 0.04532f
C1514 VP.n52 VSUBS 0.031221f
C1515 VP.n53 VSUBS 0.031221f
C1516 VP.n54 VSUBS 0.04189f
C1517 VP.n55 VSUBS 0.057896f
C1518 VP.n56 VSUBS 0.062666f
C1519 VP.n57 VSUBS 0.031221f
C1520 VP.n58 VSUBS 0.031221f
C1521 VP.n59 VSUBS 0.031221f
C1522 VP.n60 VSUBS 0.059966f
C1523 VP.n61 VSUBS 0.057896f
C1524 VP.n62 VSUBS 0.047035f
C1525 VP.n63 VSUBS 0.050382f
C1526 VP.n64 VSUBS 1.97296f
C1527 VP.n65 VSUBS 1.99384f
C1528 VP.n66 VSUBS 0.050382f
C1529 VP.n67 VSUBS 0.047035f
C1530 VP.n68 VSUBS 0.057896f
C1531 VP.n69 VSUBS 0.059966f
C1532 VP.n70 VSUBS 0.031221f
C1533 VP.n71 VSUBS 0.031221f
C1534 VP.n72 VSUBS 0.031221f
C1535 VP.n73 VSUBS 0.062666f
C1536 VP.n74 VSUBS 0.057896f
C1537 VP.n75 VSUBS 0.04189f
C1538 VP.n76 VSUBS 0.031221f
C1539 VP.n77 VSUBS 0.031221f
C1540 VP.n78 VSUBS 0.04532f
C1541 VP.n79 VSUBS 0.057896f
C1542 VP.n80 VSUBS 0.061216f
C1543 VP.n81 VSUBS 0.031221f
C1544 VP.n82 VSUBS 0.031221f
C1545 VP.n83 VSUBS 0.031221f
C1546 VP.n84 VSUBS 0.062142f
C1547 VP.n85 VSUBS 0.057896f
C1548 VP.n86 VSUBS 0.043605f
C1549 VP.n87 VSUBS 0.031221f
C1550 VP.n88 VSUBS 0.031221f
C1551 VP.n89 VSUBS 0.043605f
C1552 VP.n90 VSUBS 0.057896f
C1553 VP.n91 VSUBS 0.062142f
C1554 VP.n92 VSUBS 0.031221f
C1555 VP.n93 VSUBS 0.031221f
C1556 VP.n94 VSUBS 0.031221f
C1557 VP.n95 VSUBS 0.061216f
C1558 VP.n96 VSUBS 0.057896f
C1559 VP.n97 VSUBS 0.04532f
C1560 VP.n98 VSUBS 0.031221f
C1561 VP.n99 VSUBS 0.031221f
C1562 VP.n100 VSUBS 0.04189f
C1563 VP.n101 VSUBS 0.057896f
C1564 VP.n102 VSUBS 0.062666f
C1565 VP.n103 VSUBS 0.031221f
C1566 VP.n104 VSUBS 0.031221f
C1567 VP.n105 VSUBS 0.031221f
C1568 VP.n106 VSUBS 0.059966f
C1569 VP.n107 VSUBS 0.057896f
C1570 VP.n108 VSUBS 0.047035f
C1571 VP.n109 VSUBS 0.050382f
C1572 VP.n110 VSUBS 0.073598f
.ends

