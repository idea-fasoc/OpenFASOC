* NGSPICE file created from diff_pair_sample_0068.ext - technology: sky130A

.subckt diff_pair_sample_0068 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=2.61
X1 B.t11 B.t9 B.t10 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=2.61
X2 B.t8 B.t6 B.t7 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=2.61
X3 B.t5 B.t3 B.t4 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=2.61
X4 VTAIL.t10 VN.t1 VDD2.t4 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=2.61
X5 VDD1.t5 VP.t0 VTAIL.t11 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=2.61
X6 VDD2.t3 VN.t2 VTAIL.t7 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=2.61
X7 VTAIL.t5 VN.t3 VDD2.t2 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=2.61
X8 VTAIL.t2 VP.t1 VDD1.t4 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=2.61
X9 VDD1.t3 VP.t2 VTAIL.t0 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=2.61
X10 VTAIL.t4 VP.t3 VDD1.t2 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=2.8809 ps=17.79 w=17.46 l=2.61
X11 VDD2.t1 VN.t4 VTAIL.t8 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=2.61
X12 VDD1.t1 VP.t4 VTAIL.t3 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=2.61
X13 VDD2.t0 VN.t5 VTAIL.t6 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=2.8809 pd=17.79 as=6.8094 ps=35.7 w=17.46 l=2.61
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=2.8809 ps=17.79 w=17.46 l=2.61
X15 B.t2 B.t0 B.t1 w_n3322_n4460# sky130_fd_pr__pfet_01v8 ad=6.8094 pd=35.7 as=0 ps=0 w=17.46 l=2.61
R0 VN.n4 VN.t0 194.712
R1 VN.n20 VN.t2 194.712
R2 VN.n29 VN.n16 161.3
R3 VN.n28 VN.n27 161.3
R4 VN.n26 VN.n17 161.3
R5 VN.n25 VN.n24 161.3
R6 VN.n23 VN.n18 161.3
R7 VN.n22 VN.n21 161.3
R8 VN.n13 VN.n0 161.3
R9 VN.n12 VN.n11 161.3
R10 VN.n10 VN.n1 161.3
R11 VN.n9 VN.n8 161.3
R12 VN.n7 VN.n2 161.3
R13 VN.n6 VN.n5 161.3
R14 VN.n3 VN.t1 161.221
R15 VN.n14 VN.t5 161.221
R16 VN.n19 VN.t3 161.221
R17 VN.n30 VN.t4 161.221
R18 VN.n15 VN.n14 101.564
R19 VN.n31 VN.n30 101.564
R20 VN.n4 VN.n3 60.3423
R21 VN.n20 VN.n19 60.3423
R22 VN.n8 VN.n1 56.5617
R23 VN.n24 VN.n17 56.5617
R24 VN VN.n31 53.1421
R25 VN.n7 VN.n6 24.5923
R26 VN.n8 VN.n7 24.5923
R27 VN.n12 VN.n1 24.5923
R28 VN.n13 VN.n12 24.5923
R29 VN.n24 VN.n23 24.5923
R30 VN.n23 VN.n22 24.5923
R31 VN.n29 VN.n28 24.5923
R32 VN.n28 VN.n17 24.5923
R33 VN.n6 VN.n3 12.2964
R34 VN.n22 VN.n19 12.2964
R35 VN.n14 VN.n13 9.3454
R36 VN.n30 VN.n29 9.3454
R37 VN.n21 VN.n20 6.87456
R38 VN.n5 VN.n4 6.87456
R39 VN.n31 VN.n16 0.278335
R40 VN.n15 VN.n0 0.278335
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153485
R52 VTAIL.n394 VTAIL.n302 756.745
R53 VTAIL.n94 VTAIL.n2 756.745
R54 VTAIL.n296 VTAIL.n204 756.745
R55 VTAIL.n196 VTAIL.n104 756.745
R56 VTAIL.n335 VTAIL.n334 585
R57 VTAIL.n337 VTAIL.n336 585
R58 VTAIL.n330 VTAIL.n329 585
R59 VTAIL.n343 VTAIL.n342 585
R60 VTAIL.n345 VTAIL.n344 585
R61 VTAIL.n326 VTAIL.n325 585
R62 VTAIL.n351 VTAIL.n350 585
R63 VTAIL.n353 VTAIL.n352 585
R64 VTAIL.n322 VTAIL.n321 585
R65 VTAIL.n359 VTAIL.n358 585
R66 VTAIL.n361 VTAIL.n360 585
R67 VTAIL.n318 VTAIL.n317 585
R68 VTAIL.n367 VTAIL.n366 585
R69 VTAIL.n369 VTAIL.n368 585
R70 VTAIL.n314 VTAIL.n313 585
R71 VTAIL.n376 VTAIL.n375 585
R72 VTAIL.n377 VTAIL.n312 585
R73 VTAIL.n379 VTAIL.n378 585
R74 VTAIL.n310 VTAIL.n309 585
R75 VTAIL.n385 VTAIL.n384 585
R76 VTAIL.n387 VTAIL.n386 585
R77 VTAIL.n306 VTAIL.n305 585
R78 VTAIL.n393 VTAIL.n392 585
R79 VTAIL.n395 VTAIL.n394 585
R80 VTAIL.n35 VTAIL.n34 585
R81 VTAIL.n37 VTAIL.n36 585
R82 VTAIL.n30 VTAIL.n29 585
R83 VTAIL.n43 VTAIL.n42 585
R84 VTAIL.n45 VTAIL.n44 585
R85 VTAIL.n26 VTAIL.n25 585
R86 VTAIL.n51 VTAIL.n50 585
R87 VTAIL.n53 VTAIL.n52 585
R88 VTAIL.n22 VTAIL.n21 585
R89 VTAIL.n59 VTAIL.n58 585
R90 VTAIL.n61 VTAIL.n60 585
R91 VTAIL.n18 VTAIL.n17 585
R92 VTAIL.n67 VTAIL.n66 585
R93 VTAIL.n69 VTAIL.n68 585
R94 VTAIL.n14 VTAIL.n13 585
R95 VTAIL.n76 VTAIL.n75 585
R96 VTAIL.n77 VTAIL.n12 585
R97 VTAIL.n79 VTAIL.n78 585
R98 VTAIL.n10 VTAIL.n9 585
R99 VTAIL.n85 VTAIL.n84 585
R100 VTAIL.n87 VTAIL.n86 585
R101 VTAIL.n6 VTAIL.n5 585
R102 VTAIL.n93 VTAIL.n92 585
R103 VTAIL.n95 VTAIL.n94 585
R104 VTAIL.n297 VTAIL.n296 585
R105 VTAIL.n295 VTAIL.n294 585
R106 VTAIL.n208 VTAIL.n207 585
R107 VTAIL.n289 VTAIL.n288 585
R108 VTAIL.n287 VTAIL.n286 585
R109 VTAIL.n212 VTAIL.n211 585
R110 VTAIL.n216 VTAIL.n214 585
R111 VTAIL.n281 VTAIL.n280 585
R112 VTAIL.n279 VTAIL.n278 585
R113 VTAIL.n218 VTAIL.n217 585
R114 VTAIL.n273 VTAIL.n272 585
R115 VTAIL.n271 VTAIL.n270 585
R116 VTAIL.n222 VTAIL.n221 585
R117 VTAIL.n265 VTAIL.n264 585
R118 VTAIL.n263 VTAIL.n262 585
R119 VTAIL.n226 VTAIL.n225 585
R120 VTAIL.n257 VTAIL.n256 585
R121 VTAIL.n255 VTAIL.n254 585
R122 VTAIL.n230 VTAIL.n229 585
R123 VTAIL.n249 VTAIL.n248 585
R124 VTAIL.n247 VTAIL.n246 585
R125 VTAIL.n234 VTAIL.n233 585
R126 VTAIL.n241 VTAIL.n240 585
R127 VTAIL.n239 VTAIL.n238 585
R128 VTAIL.n197 VTAIL.n196 585
R129 VTAIL.n195 VTAIL.n194 585
R130 VTAIL.n108 VTAIL.n107 585
R131 VTAIL.n189 VTAIL.n188 585
R132 VTAIL.n187 VTAIL.n186 585
R133 VTAIL.n112 VTAIL.n111 585
R134 VTAIL.n116 VTAIL.n114 585
R135 VTAIL.n181 VTAIL.n180 585
R136 VTAIL.n179 VTAIL.n178 585
R137 VTAIL.n118 VTAIL.n117 585
R138 VTAIL.n173 VTAIL.n172 585
R139 VTAIL.n171 VTAIL.n170 585
R140 VTAIL.n122 VTAIL.n121 585
R141 VTAIL.n165 VTAIL.n164 585
R142 VTAIL.n163 VTAIL.n162 585
R143 VTAIL.n126 VTAIL.n125 585
R144 VTAIL.n157 VTAIL.n156 585
R145 VTAIL.n155 VTAIL.n154 585
R146 VTAIL.n130 VTAIL.n129 585
R147 VTAIL.n149 VTAIL.n148 585
R148 VTAIL.n147 VTAIL.n146 585
R149 VTAIL.n134 VTAIL.n133 585
R150 VTAIL.n141 VTAIL.n140 585
R151 VTAIL.n139 VTAIL.n138 585
R152 VTAIL.n333 VTAIL.t6 327.466
R153 VTAIL.n33 VTAIL.t11 327.466
R154 VTAIL.n237 VTAIL.t3 327.466
R155 VTAIL.n137 VTAIL.t7 327.466
R156 VTAIL.n336 VTAIL.n335 171.744
R157 VTAIL.n336 VTAIL.n329 171.744
R158 VTAIL.n343 VTAIL.n329 171.744
R159 VTAIL.n344 VTAIL.n343 171.744
R160 VTAIL.n344 VTAIL.n325 171.744
R161 VTAIL.n351 VTAIL.n325 171.744
R162 VTAIL.n352 VTAIL.n351 171.744
R163 VTAIL.n352 VTAIL.n321 171.744
R164 VTAIL.n359 VTAIL.n321 171.744
R165 VTAIL.n360 VTAIL.n359 171.744
R166 VTAIL.n360 VTAIL.n317 171.744
R167 VTAIL.n367 VTAIL.n317 171.744
R168 VTAIL.n368 VTAIL.n367 171.744
R169 VTAIL.n368 VTAIL.n313 171.744
R170 VTAIL.n376 VTAIL.n313 171.744
R171 VTAIL.n377 VTAIL.n376 171.744
R172 VTAIL.n378 VTAIL.n377 171.744
R173 VTAIL.n378 VTAIL.n309 171.744
R174 VTAIL.n385 VTAIL.n309 171.744
R175 VTAIL.n386 VTAIL.n385 171.744
R176 VTAIL.n386 VTAIL.n305 171.744
R177 VTAIL.n393 VTAIL.n305 171.744
R178 VTAIL.n394 VTAIL.n393 171.744
R179 VTAIL.n36 VTAIL.n35 171.744
R180 VTAIL.n36 VTAIL.n29 171.744
R181 VTAIL.n43 VTAIL.n29 171.744
R182 VTAIL.n44 VTAIL.n43 171.744
R183 VTAIL.n44 VTAIL.n25 171.744
R184 VTAIL.n51 VTAIL.n25 171.744
R185 VTAIL.n52 VTAIL.n51 171.744
R186 VTAIL.n52 VTAIL.n21 171.744
R187 VTAIL.n59 VTAIL.n21 171.744
R188 VTAIL.n60 VTAIL.n59 171.744
R189 VTAIL.n60 VTAIL.n17 171.744
R190 VTAIL.n67 VTAIL.n17 171.744
R191 VTAIL.n68 VTAIL.n67 171.744
R192 VTAIL.n68 VTAIL.n13 171.744
R193 VTAIL.n76 VTAIL.n13 171.744
R194 VTAIL.n77 VTAIL.n76 171.744
R195 VTAIL.n78 VTAIL.n77 171.744
R196 VTAIL.n78 VTAIL.n9 171.744
R197 VTAIL.n85 VTAIL.n9 171.744
R198 VTAIL.n86 VTAIL.n85 171.744
R199 VTAIL.n86 VTAIL.n5 171.744
R200 VTAIL.n93 VTAIL.n5 171.744
R201 VTAIL.n94 VTAIL.n93 171.744
R202 VTAIL.n296 VTAIL.n295 171.744
R203 VTAIL.n295 VTAIL.n207 171.744
R204 VTAIL.n288 VTAIL.n207 171.744
R205 VTAIL.n288 VTAIL.n287 171.744
R206 VTAIL.n287 VTAIL.n211 171.744
R207 VTAIL.n216 VTAIL.n211 171.744
R208 VTAIL.n280 VTAIL.n216 171.744
R209 VTAIL.n280 VTAIL.n279 171.744
R210 VTAIL.n279 VTAIL.n217 171.744
R211 VTAIL.n272 VTAIL.n217 171.744
R212 VTAIL.n272 VTAIL.n271 171.744
R213 VTAIL.n271 VTAIL.n221 171.744
R214 VTAIL.n264 VTAIL.n221 171.744
R215 VTAIL.n264 VTAIL.n263 171.744
R216 VTAIL.n263 VTAIL.n225 171.744
R217 VTAIL.n256 VTAIL.n225 171.744
R218 VTAIL.n256 VTAIL.n255 171.744
R219 VTAIL.n255 VTAIL.n229 171.744
R220 VTAIL.n248 VTAIL.n229 171.744
R221 VTAIL.n248 VTAIL.n247 171.744
R222 VTAIL.n247 VTAIL.n233 171.744
R223 VTAIL.n240 VTAIL.n233 171.744
R224 VTAIL.n240 VTAIL.n239 171.744
R225 VTAIL.n196 VTAIL.n195 171.744
R226 VTAIL.n195 VTAIL.n107 171.744
R227 VTAIL.n188 VTAIL.n107 171.744
R228 VTAIL.n188 VTAIL.n187 171.744
R229 VTAIL.n187 VTAIL.n111 171.744
R230 VTAIL.n116 VTAIL.n111 171.744
R231 VTAIL.n180 VTAIL.n116 171.744
R232 VTAIL.n180 VTAIL.n179 171.744
R233 VTAIL.n179 VTAIL.n117 171.744
R234 VTAIL.n172 VTAIL.n117 171.744
R235 VTAIL.n172 VTAIL.n171 171.744
R236 VTAIL.n171 VTAIL.n121 171.744
R237 VTAIL.n164 VTAIL.n121 171.744
R238 VTAIL.n164 VTAIL.n163 171.744
R239 VTAIL.n163 VTAIL.n125 171.744
R240 VTAIL.n156 VTAIL.n125 171.744
R241 VTAIL.n156 VTAIL.n155 171.744
R242 VTAIL.n155 VTAIL.n129 171.744
R243 VTAIL.n148 VTAIL.n129 171.744
R244 VTAIL.n148 VTAIL.n147 171.744
R245 VTAIL.n147 VTAIL.n133 171.744
R246 VTAIL.n140 VTAIL.n133 171.744
R247 VTAIL.n140 VTAIL.n139 171.744
R248 VTAIL.n335 VTAIL.t6 85.8723
R249 VTAIL.n35 VTAIL.t11 85.8723
R250 VTAIL.n239 VTAIL.t3 85.8723
R251 VTAIL.n139 VTAIL.t7 85.8723
R252 VTAIL.n203 VTAIL.n202 51.1798
R253 VTAIL.n103 VTAIL.n102 51.1798
R254 VTAIL.n1 VTAIL.n0 51.1796
R255 VTAIL.n101 VTAIL.n100 51.1796
R256 VTAIL.n103 VTAIL.n101 32.4876
R257 VTAIL.n399 VTAIL.n398 31.0217
R258 VTAIL.n99 VTAIL.n98 31.0217
R259 VTAIL.n301 VTAIL.n300 31.0217
R260 VTAIL.n201 VTAIL.n200 31.0217
R261 VTAIL.n399 VTAIL.n301 29.9531
R262 VTAIL.n334 VTAIL.n333 16.3895
R263 VTAIL.n34 VTAIL.n33 16.3895
R264 VTAIL.n238 VTAIL.n237 16.3895
R265 VTAIL.n138 VTAIL.n137 16.3895
R266 VTAIL.n379 VTAIL.n310 13.1884
R267 VTAIL.n79 VTAIL.n10 13.1884
R268 VTAIL.n214 VTAIL.n212 13.1884
R269 VTAIL.n114 VTAIL.n112 13.1884
R270 VTAIL.n337 VTAIL.n332 12.8005
R271 VTAIL.n380 VTAIL.n312 12.8005
R272 VTAIL.n384 VTAIL.n383 12.8005
R273 VTAIL.n37 VTAIL.n32 12.8005
R274 VTAIL.n80 VTAIL.n12 12.8005
R275 VTAIL.n84 VTAIL.n83 12.8005
R276 VTAIL.n286 VTAIL.n285 12.8005
R277 VTAIL.n282 VTAIL.n281 12.8005
R278 VTAIL.n241 VTAIL.n236 12.8005
R279 VTAIL.n186 VTAIL.n185 12.8005
R280 VTAIL.n182 VTAIL.n181 12.8005
R281 VTAIL.n141 VTAIL.n136 12.8005
R282 VTAIL.n338 VTAIL.n330 12.0247
R283 VTAIL.n375 VTAIL.n374 12.0247
R284 VTAIL.n387 VTAIL.n308 12.0247
R285 VTAIL.n38 VTAIL.n30 12.0247
R286 VTAIL.n75 VTAIL.n74 12.0247
R287 VTAIL.n87 VTAIL.n8 12.0247
R288 VTAIL.n289 VTAIL.n210 12.0247
R289 VTAIL.n278 VTAIL.n215 12.0247
R290 VTAIL.n242 VTAIL.n234 12.0247
R291 VTAIL.n189 VTAIL.n110 12.0247
R292 VTAIL.n178 VTAIL.n115 12.0247
R293 VTAIL.n142 VTAIL.n134 12.0247
R294 VTAIL.n342 VTAIL.n341 11.249
R295 VTAIL.n373 VTAIL.n314 11.249
R296 VTAIL.n388 VTAIL.n306 11.249
R297 VTAIL.n42 VTAIL.n41 11.249
R298 VTAIL.n73 VTAIL.n14 11.249
R299 VTAIL.n88 VTAIL.n6 11.249
R300 VTAIL.n290 VTAIL.n208 11.249
R301 VTAIL.n277 VTAIL.n218 11.249
R302 VTAIL.n246 VTAIL.n245 11.249
R303 VTAIL.n190 VTAIL.n108 11.249
R304 VTAIL.n177 VTAIL.n118 11.249
R305 VTAIL.n146 VTAIL.n145 11.249
R306 VTAIL.n345 VTAIL.n328 10.4732
R307 VTAIL.n370 VTAIL.n369 10.4732
R308 VTAIL.n392 VTAIL.n391 10.4732
R309 VTAIL.n45 VTAIL.n28 10.4732
R310 VTAIL.n70 VTAIL.n69 10.4732
R311 VTAIL.n92 VTAIL.n91 10.4732
R312 VTAIL.n294 VTAIL.n293 10.4732
R313 VTAIL.n274 VTAIL.n273 10.4732
R314 VTAIL.n249 VTAIL.n232 10.4732
R315 VTAIL.n194 VTAIL.n193 10.4732
R316 VTAIL.n174 VTAIL.n173 10.4732
R317 VTAIL.n149 VTAIL.n132 10.4732
R318 VTAIL.n346 VTAIL.n326 9.69747
R319 VTAIL.n366 VTAIL.n316 9.69747
R320 VTAIL.n395 VTAIL.n304 9.69747
R321 VTAIL.n46 VTAIL.n26 9.69747
R322 VTAIL.n66 VTAIL.n16 9.69747
R323 VTAIL.n95 VTAIL.n4 9.69747
R324 VTAIL.n297 VTAIL.n206 9.69747
R325 VTAIL.n270 VTAIL.n220 9.69747
R326 VTAIL.n250 VTAIL.n230 9.69747
R327 VTAIL.n197 VTAIL.n106 9.69747
R328 VTAIL.n170 VTAIL.n120 9.69747
R329 VTAIL.n150 VTAIL.n130 9.69747
R330 VTAIL.n398 VTAIL.n397 9.45567
R331 VTAIL.n98 VTAIL.n97 9.45567
R332 VTAIL.n300 VTAIL.n299 9.45567
R333 VTAIL.n200 VTAIL.n199 9.45567
R334 VTAIL.n397 VTAIL.n396 9.3005
R335 VTAIL.n304 VTAIL.n303 9.3005
R336 VTAIL.n391 VTAIL.n390 9.3005
R337 VTAIL.n389 VTAIL.n388 9.3005
R338 VTAIL.n308 VTAIL.n307 9.3005
R339 VTAIL.n383 VTAIL.n382 9.3005
R340 VTAIL.n355 VTAIL.n354 9.3005
R341 VTAIL.n324 VTAIL.n323 9.3005
R342 VTAIL.n349 VTAIL.n348 9.3005
R343 VTAIL.n347 VTAIL.n346 9.3005
R344 VTAIL.n328 VTAIL.n327 9.3005
R345 VTAIL.n341 VTAIL.n340 9.3005
R346 VTAIL.n339 VTAIL.n338 9.3005
R347 VTAIL.n332 VTAIL.n331 9.3005
R348 VTAIL.n357 VTAIL.n356 9.3005
R349 VTAIL.n320 VTAIL.n319 9.3005
R350 VTAIL.n363 VTAIL.n362 9.3005
R351 VTAIL.n365 VTAIL.n364 9.3005
R352 VTAIL.n316 VTAIL.n315 9.3005
R353 VTAIL.n371 VTAIL.n370 9.3005
R354 VTAIL.n373 VTAIL.n372 9.3005
R355 VTAIL.n374 VTAIL.n311 9.3005
R356 VTAIL.n381 VTAIL.n380 9.3005
R357 VTAIL.n97 VTAIL.n96 9.3005
R358 VTAIL.n4 VTAIL.n3 9.3005
R359 VTAIL.n91 VTAIL.n90 9.3005
R360 VTAIL.n89 VTAIL.n88 9.3005
R361 VTAIL.n8 VTAIL.n7 9.3005
R362 VTAIL.n83 VTAIL.n82 9.3005
R363 VTAIL.n55 VTAIL.n54 9.3005
R364 VTAIL.n24 VTAIL.n23 9.3005
R365 VTAIL.n49 VTAIL.n48 9.3005
R366 VTAIL.n47 VTAIL.n46 9.3005
R367 VTAIL.n28 VTAIL.n27 9.3005
R368 VTAIL.n41 VTAIL.n40 9.3005
R369 VTAIL.n39 VTAIL.n38 9.3005
R370 VTAIL.n32 VTAIL.n31 9.3005
R371 VTAIL.n57 VTAIL.n56 9.3005
R372 VTAIL.n20 VTAIL.n19 9.3005
R373 VTAIL.n63 VTAIL.n62 9.3005
R374 VTAIL.n65 VTAIL.n64 9.3005
R375 VTAIL.n16 VTAIL.n15 9.3005
R376 VTAIL.n71 VTAIL.n70 9.3005
R377 VTAIL.n73 VTAIL.n72 9.3005
R378 VTAIL.n74 VTAIL.n11 9.3005
R379 VTAIL.n81 VTAIL.n80 9.3005
R380 VTAIL.n224 VTAIL.n223 9.3005
R381 VTAIL.n267 VTAIL.n266 9.3005
R382 VTAIL.n269 VTAIL.n268 9.3005
R383 VTAIL.n220 VTAIL.n219 9.3005
R384 VTAIL.n275 VTAIL.n274 9.3005
R385 VTAIL.n277 VTAIL.n276 9.3005
R386 VTAIL.n215 VTAIL.n213 9.3005
R387 VTAIL.n283 VTAIL.n282 9.3005
R388 VTAIL.n299 VTAIL.n298 9.3005
R389 VTAIL.n206 VTAIL.n205 9.3005
R390 VTAIL.n293 VTAIL.n292 9.3005
R391 VTAIL.n291 VTAIL.n290 9.3005
R392 VTAIL.n210 VTAIL.n209 9.3005
R393 VTAIL.n285 VTAIL.n284 9.3005
R394 VTAIL.n261 VTAIL.n260 9.3005
R395 VTAIL.n259 VTAIL.n258 9.3005
R396 VTAIL.n228 VTAIL.n227 9.3005
R397 VTAIL.n253 VTAIL.n252 9.3005
R398 VTAIL.n251 VTAIL.n250 9.3005
R399 VTAIL.n232 VTAIL.n231 9.3005
R400 VTAIL.n245 VTAIL.n244 9.3005
R401 VTAIL.n243 VTAIL.n242 9.3005
R402 VTAIL.n236 VTAIL.n235 9.3005
R403 VTAIL.n124 VTAIL.n123 9.3005
R404 VTAIL.n167 VTAIL.n166 9.3005
R405 VTAIL.n169 VTAIL.n168 9.3005
R406 VTAIL.n120 VTAIL.n119 9.3005
R407 VTAIL.n175 VTAIL.n174 9.3005
R408 VTAIL.n177 VTAIL.n176 9.3005
R409 VTAIL.n115 VTAIL.n113 9.3005
R410 VTAIL.n183 VTAIL.n182 9.3005
R411 VTAIL.n199 VTAIL.n198 9.3005
R412 VTAIL.n106 VTAIL.n105 9.3005
R413 VTAIL.n193 VTAIL.n192 9.3005
R414 VTAIL.n191 VTAIL.n190 9.3005
R415 VTAIL.n110 VTAIL.n109 9.3005
R416 VTAIL.n185 VTAIL.n184 9.3005
R417 VTAIL.n161 VTAIL.n160 9.3005
R418 VTAIL.n159 VTAIL.n158 9.3005
R419 VTAIL.n128 VTAIL.n127 9.3005
R420 VTAIL.n153 VTAIL.n152 9.3005
R421 VTAIL.n151 VTAIL.n150 9.3005
R422 VTAIL.n132 VTAIL.n131 9.3005
R423 VTAIL.n145 VTAIL.n144 9.3005
R424 VTAIL.n143 VTAIL.n142 9.3005
R425 VTAIL.n136 VTAIL.n135 9.3005
R426 VTAIL.n350 VTAIL.n349 8.92171
R427 VTAIL.n365 VTAIL.n318 8.92171
R428 VTAIL.n396 VTAIL.n302 8.92171
R429 VTAIL.n50 VTAIL.n49 8.92171
R430 VTAIL.n65 VTAIL.n18 8.92171
R431 VTAIL.n96 VTAIL.n2 8.92171
R432 VTAIL.n298 VTAIL.n204 8.92171
R433 VTAIL.n269 VTAIL.n222 8.92171
R434 VTAIL.n254 VTAIL.n253 8.92171
R435 VTAIL.n198 VTAIL.n104 8.92171
R436 VTAIL.n169 VTAIL.n122 8.92171
R437 VTAIL.n154 VTAIL.n153 8.92171
R438 VTAIL.n353 VTAIL.n324 8.14595
R439 VTAIL.n362 VTAIL.n361 8.14595
R440 VTAIL.n53 VTAIL.n24 8.14595
R441 VTAIL.n62 VTAIL.n61 8.14595
R442 VTAIL.n266 VTAIL.n265 8.14595
R443 VTAIL.n257 VTAIL.n228 8.14595
R444 VTAIL.n166 VTAIL.n165 8.14595
R445 VTAIL.n157 VTAIL.n128 8.14595
R446 VTAIL.n354 VTAIL.n322 7.3702
R447 VTAIL.n358 VTAIL.n320 7.3702
R448 VTAIL.n54 VTAIL.n22 7.3702
R449 VTAIL.n58 VTAIL.n20 7.3702
R450 VTAIL.n262 VTAIL.n224 7.3702
R451 VTAIL.n258 VTAIL.n226 7.3702
R452 VTAIL.n162 VTAIL.n124 7.3702
R453 VTAIL.n158 VTAIL.n126 7.3702
R454 VTAIL.n357 VTAIL.n322 6.59444
R455 VTAIL.n358 VTAIL.n357 6.59444
R456 VTAIL.n57 VTAIL.n22 6.59444
R457 VTAIL.n58 VTAIL.n57 6.59444
R458 VTAIL.n262 VTAIL.n261 6.59444
R459 VTAIL.n261 VTAIL.n226 6.59444
R460 VTAIL.n162 VTAIL.n161 6.59444
R461 VTAIL.n161 VTAIL.n126 6.59444
R462 VTAIL.n354 VTAIL.n353 5.81868
R463 VTAIL.n361 VTAIL.n320 5.81868
R464 VTAIL.n54 VTAIL.n53 5.81868
R465 VTAIL.n61 VTAIL.n20 5.81868
R466 VTAIL.n265 VTAIL.n224 5.81868
R467 VTAIL.n258 VTAIL.n257 5.81868
R468 VTAIL.n165 VTAIL.n124 5.81868
R469 VTAIL.n158 VTAIL.n157 5.81868
R470 VTAIL.n350 VTAIL.n324 5.04292
R471 VTAIL.n362 VTAIL.n318 5.04292
R472 VTAIL.n398 VTAIL.n302 5.04292
R473 VTAIL.n50 VTAIL.n24 5.04292
R474 VTAIL.n62 VTAIL.n18 5.04292
R475 VTAIL.n98 VTAIL.n2 5.04292
R476 VTAIL.n300 VTAIL.n204 5.04292
R477 VTAIL.n266 VTAIL.n222 5.04292
R478 VTAIL.n254 VTAIL.n228 5.04292
R479 VTAIL.n200 VTAIL.n104 5.04292
R480 VTAIL.n166 VTAIL.n122 5.04292
R481 VTAIL.n154 VTAIL.n128 5.04292
R482 VTAIL.n349 VTAIL.n326 4.26717
R483 VTAIL.n366 VTAIL.n365 4.26717
R484 VTAIL.n396 VTAIL.n395 4.26717
R485 VTAIL.n49 VTAIL.n26 4.26717
R486 VTAIL.n66 VTAIL.n65 4.26717
R487 VTAIL.n96 VTAIL.n95 4.26717
R488 VTAIL.n298 VTAIL.n297 4.26717
R489 VTAIL.n270 VTAIL.n269 4.26717
R490 VTAIL.n253 VTAIL.n230 4.26717
R491 VTAIL.n198 VTAIL.n197 4.26717
R492 VTAIL.n170 VTAIL.n169 4.26717
R493 VTAIL.n153 VTAIL.n130 4.26717
R494 VTAIL.n333 VTAIL.n331 3.70982
R495 VTAIL.n33 VTAIL.n31 3.70982
R496 VTAIL.n237 VTAIL.n235 3.70982
R497 VTAIL.n137 VTAIL.n135 3.70982
R498 VTAIL.n346 VTAIL.n345 3.49141
R499 VTAIL.n369 VTAIL.n316 3.49141
R500 VTAIL.n392 VTAIL.n304 3.49141
R501 VTAIL.n46 VTAIL.n45 3.49141
R502 VTAIL.n69 VTAIL.n16 3.49141
R503 VTAIL.n92 VTAIL.n4 3.49141
R504 VTAIL.n294 VTAIL.n206 3.49141
R505 VTAIL.n273 VTAIL.n220 3.49141
R506 VTAIL.n250 VTAIL.n249 3.49141
R507 VTAIL.n194 VTAIL.n106 3.49141
R508 VTAIL.n173 VTAIL.n120 3.49141
R509 VTAIL.n150 VTAIL.n149 3.49141
R510 VTAIL.n342 VTAIL.n328 2.71565
R511 VTAIL.n370 VTAIL.n314 2.71565
R512 VTAIL.n391 VTAIL.n306 2.71565
R513 VTAIL.n42 VTAIL.n28 2.71565
R514 VTAIL.n70 VTAIL.n14 2.71565
R515 VTAIL.n91 VTAIL.n6 2.71565
R516 VTAIL.n293 VTAIL.n208 2.71565
R517 VTAIL.n274 VTAIL.n218 2.71565
R518 VTAIL.n246 VTAIL.n232 2.71565
R519 VTAIL.n193 VTAIL.n108 2.71565
R520 VTAIL.n174 VTAIL.n118 2.71565
R521 VTAIL.n146 VTAIL.n132 2.71565
R522 VTAIL.n201 VTAIL.n103 2.53498
R523 VTAIL.n301 VTAIL.n203 2.53498
R524 VTAIL.n101 VTAIL.n99 2.53498
R525 VTAIL.n341 VTAIL.n330 1.93989
R526 VTAIL.n375 VTAIL.n373 1.93989
R527 VTAIL.n388 VTAIL.n387 1.93989
R528 VTAIL.n41 VTAIL.n30 1.93989
R529 VTAIL.n75 VTAIL.n73 1.93989
R530 VTAIL.n88 VTAIL.n87 1.93989
R531 VTAIL.n290 VTAIL.n289 1.93989
R532 VTAIL.n278 VTAIL.n277 1.93989
R533 VTAIL.n245 VTAIL.n234 1.93989
R534 VTAIL.n190 VTAIL.n189 1.93989
R535 VTAIL.n178 VTAIL.n177 1.93989
R536 VTAIL.n145 VTAIL.n134 1.93989
R537 VTAIL.n0 VTAIL.t9 1.86218
R538 VTAIL.n0 VTAIL.t10 1.86218
R539 VTAIL.n100 VTAIL.t1 1.86218
R540 VTAIL.n100 VTAIL.t2 1.86218
R541 VTAIL.n202 VTAIL.t0 1.86218
R542 VTAIL.n202 VTAIL.t4 1.86218
R543 VTAIL.n102 VTAIL.t8 1.86218
R544 VTAIL.n102 VTAIL.t5 1.86218
R545 VTAIL VTAIL.n399 1.84317
R546 VTAIL.n203 VTAIL.n201 1.73757
R547 VTAIL.n99 VTAIL.n1 1.73757
R548 VTAIL.n338 VTAIL.n337 1.16414
R549 VTAIL.n374 VTAIL.n312 1.16414
R550 VTAIL.n384 VTAIL.n308 1.16414
R551 VTAIL.n38 VTAIL.n37 1.16414
R552 VTAIL.n74 VTAIL.n12 1.16414
R553 VTAIL.n84 VTAIL.n8 1.16414
R554 VTAIL.n286 VTAIL.n210 1.16414
R555 VTAIL.n281 VTAIL.n215 1.16414
R556 VTAIL.n242 VTAIL.n241 1.16414
R557 VTAIL.n186 VTAIL.n110 1.16414
R558 VTAIL.n181 VTAIL.n115 1.16414
R559 VTAIL.n142 VTAIL.n141 1.16414
R560 VTAIL VTAIL.n1 0.69231
R561 VTAIL.n334 VTAIL.n332 0.388379
R562 VTAIL.n380 VTAIL.n379 0.388379
R563 VTAIL.n383 VTAIL.n310 0.388379
R564 VTAIL.n34 VTAIL.n32 0.388379
R565 VTAIL.n80 VTAIL.n79 0.388379
R566 VTAIL.n83 VTAIL.n10 0.388379
R567 VTAIL.n285 VTAIL.n212 0.388379
R568 VTAIL.n282 VTAIL.n214 0.388379
R569 VTAIL.n238 VTAIL.n236 0.388379
R570 VTAIL.n185 VTAIL.n112 0.388379
R571 VTAIL.n182 VTAIL.n114 0.388379
R572 VTAIL.n138 VTAIL.n136 0.388379
R573 VTAIL.n339 VTAIL.n331 0.155672
R574 VTAIL.n340 VTAIL.n339 0.155672
R575 VTAIL.n340 VTAIL.n327 0.155672
R576 VTAIL.n347 VTAIL.n327 0.155672
R577 VTAIL.n348 VTAIL.n347 0.155672
R578 VTAIL.n348 VTAIL.n323 0.155672
R579 VTAIL.n355 VTAIL.n323 0.155672
R580 VTAIL.n356 VTAIL.n355 0.155672
R581 VTAIL.n356 VTAIL.n319 0.155672
R582 VTAIL.n363 VTAIL.n319 0.155672
R583 VTAIL.n364 VTAIL.n363 0.155672
R584 VTAIL.n364 VTAIL.n315 0.155672
R585 VTAIL.n371 VTAIL.n315 0.155672
R586 VTAIL.n372 VTAIL.n371 0.155672
R587 VTAIL.n372 VTAIL.n311 0.155672
R588 VTAIL.n381 VTAIL.n311 0.155672
R589 VTAIL.n382 VTAIL.n381 0.155672
R590 VTAIL.n382 VTAIL.n307 0.155672
R591 VTAIL.n389 VTAIL.n307 0.155672
R592 VTAIL.n390 VTAIL.n389 0.155672
R593 VTAIL.n390 VTAIL.n303 0.155672
R594 VTAIL.n397 VTAIL.n303 0.155672
R595 VTAIL.n39 VTAIL.n31 0.155672
R596 VTAIL.n40 VTAIL.n39 0.155672
R597 VTAIL.n40 VTAIL.n27 0.155672
R598 VTAIL.n47 VTAIL.n27 0.155672
R599 VTAIL.n48 VTAIL.n47 0.155672
R600 VTAIL.n48 VTAIL.n23 0.155672
R601 VTAIL.n55 VTAIL.n23 0.155672
R602 VTAIL.n56 VTAIL.n55 0.155672
R603 VTAIL.n56 VTAIL.n19 0.155672
R604 VTAIL.n63 VTAIL.n19 0.155672
R605 VTAIL.n64 VTAIL.n63 0.155672
R606 VTAIL.n64 VTAIL.n15 0.155672
R607 VTAIL.n71 VTAIL.n15 0.155672
R608 VTAIL.n72 VTAIL.n71 0.155672
R609 VTAIL.n72 VTAIL.n11 0.155672
R610 VTAIL.n81 VTAIL.n11 0.155672
R611 VTAIL.n82 VTAIL.n81 0.155672
R612 VTAIL.n82 VTAIL.n7 0.155672
R613 VTAIL.n89 VTAIL.n7 0.155672
R614 VTAIL.n90 VTAIL.n89 0.155672
R615 VTAIL.n90 VTAIL.n3 0.155672
R616 VTAIL.n97 VTAIL.n3 0.155672
R617 VTAIL.n299 VTAIL.n205 0.155672
R618 VTAIL.n292 VTAIL.n205 0.155672
R619 VTAIL.n292 VTAIL.n291 0.155672
R620 VTAIL.n291 VTAIL.n209 0.155672
R621 VTAIL.n284 VTAIL.n209 0.155672
R622 VTAIL.n284 VTAIL.n283 0.155672
R623 VTAIL.n283 VTAIL.n213 0.155672
R624 VTAIL.n276 VTAIL.n213 0.155672
R625 VTAIL.n276 VTAIL.n275 0.155672
R626 VTAIL.n275 VTAIL.n219 0.155672
R627 VTAIL.n268 VTAIL.n219 0.155672
R628 VTAIL.n268 VTAIL.n267 0.155672
R629 VTAIL.n267 VTAIL.n223 0.155672
R630 VTAIL.n260 VTAIL.n223 0.155672
R631 VTAIL.n260 VTAIL.n259 0.155672
R632 VTAIL.n259 VTAIL.n227 0.155672
R633 VTAIL.n252 VTAIL.n227 0.155672
R634 VTAIL.n252 VTAIL.n251 0.155672
R635 VTAIL.n251 VTAIL.n231 0.155672
R636 VTAIL.n244 VTAIL.n231 0.155672
R637 VTAIL.n244 VTAIL.n243 0.155672
R638 VTAIL.n243 VTAIL.n235 0.155672
R639 VTAIL.n199 VTAIL.n105 0.155672
R640 VTAIL.n192 VTAIL.n105 0.155672
R641 VTAIL.n192 VTAIL.n191 0.155672
R642 VTAIL.n191 VTAIL.n109 0.155672
R643 VTAIL.n184 VTAIL.n109 0.155672
R644 VTAIL.n184 VTAIL.n183 0.155672
R645 VTAIL.n183 VTAIL.n113 0.155672
R646 VTAIL.n176 VTAIL.n113 0.155672
R647 VTAIL.n176 VTAIL.n175 0.155672
R648 VTAIL.n175 VTAIL.n119 0.155672
R649 VTAIL.n168 VTAIL.n119 0.155672
R650 VTAIL.n168 VTAIL.n167 0.155672
R651 VTAIL.n167 VTAIL.n123 0.155672
R652 VTAIL.n160 VTAIL.n123 0.155672
R653 VTAIL.n160 VTAIL.n159 0.155672
R654 VTAIL.n159 VTAIL.n127 0.155672
R655 VTAIL.n152 VTAIL.n127 0.155672
R656 VTAIL.n152 VTAIL.n151 0.155672
R657 VTAIL.n151 VTAIL.n131 0.155672
R658 VTAIL.n144 VTAIL.n131 0.155672
R659 VTAIL.n144 VTAIL.n143 0.155672
R660 VTAIL.n143 VTAIL.n135 0.155672
R661 VDD2.n191 VDD2.n99 756.745
R662 VDD2.n92 VDD2.n0 756.745
R663 VDD2.n192 VDD2.n191 585
R664 VDD2.n190 VDD2.n189 585
R665 VDD2.n103 VDD2.n102 585
R666 VDD2.n184 VDD2.n183 585
R667 VDD2.n182 VDD2.n181 585
R668 VDD2.n107 VDD2.n106 585
R669 VDD2.n111 VDD2.n109 585
R670 VDD2.n176 VDD2.n175 585
R671 VDD2.n174 VDD2.n173 585
R672 VDD2.n113 VDD2.n112 585
R673 VDD2.n168 VDD2.n167 585
R674 VDD2.n166 VDD2.n165 585
R675 VDD2.n117 VDD2.n116 585
R676 VDD2.n160 VDD2.n159 585
R677 VDD2.n158 VDD2.n157 585
R678 VDD2.n121 VDD2.n120 585
R679 VDD2.n152 VDD2.n151 585
R680 VDD2.n150 VDD2.n149 585
R681 VDD2.n125 VDD2.n124 585
R682 VDD2.n144 VDD2.n143 585
R683 VDD2.n142 VDD2.n141 585
R684 VDD2.n129 VDD2.n128 585
R685 VDD2.n136 VDD2.n135 585
R686 VDD2.n134 VDD2.n133 585
R687 VDD2.n33 VDD2.n32 585
R688 VDD2.n35 VDD2.n34 585
R689 VDD2.n28 VDD2.n27 585
R690 VDD2.n41 VDD2.n40 585
R691 VDD2.n43 VDD2.n42 585
R692 VDD2.n24 VDD2.n23 585
R693 VDD2.n49 VDD2.n48 585
R694 VDD2.n51 VDD2.n50 585
R695 VDD2.n20 VDD2.n19 585
R696 VDD2.n57 VDD2.n56 585
R697 VDD2.n59 VDD2.n58 585
R698 VDD2.n16 VDD2.n15 585
R699 VDD2.n65 VDD2.n64 585
R700 VDD2.n67 VDD2.n66 585
R701 VDD2.n12 VDD2.n11 585
R702 VDD2.n74 VDD2.n73 585
R703 VDD2.n75 VDD2.n10 585
R704 VDD2.n77 VDD2.n76 585
R705 VDD2.n8 VDD2.n7 585
R706 VDD2.n83 VDD2.n82 585
R707 VDD2.n85 VDD2.n84 585
R708 VDD2.n4 VDD2.n3 585
R709 VDD2.n91 VDD2.n90 585
R710 VDD2.n93 VDD2.n92 585
R711 VDD2.n132 VDD2.t1 327.466
R712 VDD2.n31 VDD2.t5 327.466
R713 VDD2.n191 VDD2.n190 171.744
R714 VDD2.n190 VDD2.n102 171.744
R715 VDD2.n183 VDD2.n102 171.744
R716 VDD2.n183 VDD2.n182 171.744
R717 VDD2.n182 VDD2.n106 171.744
R718 VDD2.n111 VDD2.n106 171.744
R719 VDD2.n175 VDD2.n111 171.744
R720 VDD2.n175 VDD2.n174 171.744
R721 VDD2.n174 VDD2.n112 171.744
R722 VDD2.n167 VDD2.n112 171.744
R723 VDD2.n167 VDD2.n166 171.744
R724 VDD2.n166 VDD2.n116 171.744
R725 VDD2.n159 VDD2.n116 171.744
R726 VDD2.n159 VDD2.n158 171.744
R727 VDD2.n158 VDD2.n120 171.744
R728 VDD2.n151 VDD2.n120 171.744
R729 VDD2.n151 VDD2.n150 171.744
R730 VDD2.n150 VDD2.n124 171.744
R731 VDD2.n143 VDD2.n124 171.744
R732 VDD2.n143 VDD2.n142 171.744
R733 VDD2.n142 VDD2.n128 171.744
R734 VDD2.n135 VDD2.n128 171.744
R735 VDD2.n135 VDD2.n134 171.744
R736 VDD2.n34 VDD2.n33 171.744
R737 VDD2.n34 VDD2.n27 171.744
R738 VDD2.n41 VDD2.n27 171.744
R739 VDD2.n42 VDD2.n41 171.744
R740 VDD2.n42 VDD2.n23 171.744
R741 VDD2.n49 VDD2.n23 171.744
R742 VDD2.n50 VDD2.n49 171.744
R743 VDD2.n50 VDD2.n19 171.744
R744 VDD2.n57 VDD2.n19 171.744
R745 VDD2.n58 VDD2.n57 171.744
R746 VDD2.n58 VDD2.n15 171.744
R747 VDD2.n65 VDD2.n15 171.744
R748 VDD2.n66 VDD2.n65 171.744
R749 VDD2.n66 VDD2.n11 171.744
R750 VDD2.n74 VDD2.n11 171.744
R751 VDD2.n75 VDD2.n74 171.744
R752 VDD2.n76 VDD2.n75 171.744
R753 VDD2.n76 VDD2.n7 171.744
R754 VDD2.n83 VDD2.n7 171.744
R755 VDD2.n84 VDD2.n83 171.744
R756 VDD2.n84 VDD2.n3 171.744
R757 VDD2.n91 VDD2.n3 171.744
R758 VDD2.n92 VDD2.n91 171.744
R759 VDD2.n134 VDD2.t1 85.8723
R760 VDD2.n33 VDD2.t5 85.8723
R761 VDD2.n98 VDD2.n97 68.4367
R762 VDD2 VDD2.n197 68.4338
R763 VDD2.n98 VDD2.n96 49.546
R764 VDD2.n196 VDD2.n195 47.7005
R765 VDD2.n196 VDD2.n98 47.0041
R766 VDD2.n133 VDD2.n132 16.3895
R767 VDD2.n32 VDD2.n31 16.3895
R768 VDD2.n109 VDD2.n107 13.1884
R769 VDD2.n77 VDD2.n8 13.1884
R770 VDD2.n181 VDD2.n180 12.8005
R771 VDD2.n177 VDD2.n176 12.8005
R772 VDD2.n136 VDD2.n131 12.8005
R773 VDD2.n35 VDD2.n30 12.8005
R774 VDD2.n78 VDD2.n10 12.8005
R775 VDD2.n82 VDD2.n81 12.8005
R776 VDD2.n184 VDD2.n105 12.0247
R777 VDD2.n173 VDD2.n110 12.0247
R778 VDD2.n137 VDD2.n129 12.0247
R779 VDD2.n36 VDD2.n28 12.0247
R780 VDD2.n73 VDD2.n72 12.0247
R781 VDD2.n85 VDD2.n6 12.0247
R782 VDD2.n185 VDD2.n103 11.249
R783 VDD2.n172 VDD2.n113 11.249
R784 VDD2.n141 VDD2.n140 11.249
R785 VDD2.n40 VDD2.n39 11.249
R786 VDD2.n71 VDD2.n12 11.249
R787 VDD2.n86 VDD2.n4 11.249
R788 VDD2.n189 VDD2.n188 10.4732
R789 VDD2.n169 VDD2.n168 10.4732
R790 VDD2.n144 VDD2.n127 10.4732
R791 VDD2.n43 VDD2.n26 10.4732
R792 VDD2.n68 VDD2.n67 10.4732
R793 VDD2.n90 VDD2.n89 10.4732
R794 VDD2.n192 VDD2.n101 9.69747
R795 VDD2.n165 VDD2.n115 9.69747
R796 VDD2.n145 VDD2.n125 9.69747
R797 VDD2.n44 VDD2.n24 9.69747
R798 VDD2.n64 VDD2.n14 9.69747
R799 VDD2.n93 VDD2.n2 9.69747
R800 VDD2.n195 VDD2.n194 9.45567
R801 VDD2.n96 VDD2.n95 9.45567
R802 VDD2.n119 VDD2.n118 9.3005
R803 VDD2.n162 VDD2.n161 9.3005
R804 VDD2.n164 VDD2.n163 9.3005
R805 VDD2.n115 VDD2.n114 9.3005
R806 VDD2.n170 VDD2.n169 9.3005
R807 VDD2.n172 VDD2.n171 9.3005
R808 VDD2.n110 VDD2.n108 9.3005
R809 VDD2.n178 VDD2.n177 9.3005
R810 VDD2.n194 VDD2.n193 9.3005
R811 VDD2.n101 VDD2.n100 9.3005
R812 VDD2.n188 VDD2.n187 9.3005
R813 VDD2.n186 VDD2.n185 9.3005
R814 VDD2.n105 VDD2.n104 9.3005
R815 VDD2.n180 VDD2.n179 9.3005
R816 VDD2.n156 VDD2.n155 9.3005
R817 VDD2.n154 VDD2.n153 9.3005
R818 VDD2.n123 VDD2.n122 9.3005
R819 VDD2.n148 VDD2.n147 9.3005
R820 VDD2.n146 VDD2.n145 9.3005
R821 VDD2.n127 VDD2.n126 9.3005
R822 VDD2.n140 VDD2.n139 9.3005
R823 VDD2.n138 VDD2.n137 9.3005
R824 VDD2.n131 VDD2.n130 9.3005
R825 VDD2.n95 VDD2.n94 9.3005
R826 VDD2.n2 VDD2.n1 9.3005
R827 VDD2.n89 VDD2.n88 9.3005
R828 VDD2.n87 VDD2.n86 9.3005
R829 VDD2.n6 VDD2.n5 9.3005
R830 VDD2.n81 VDD2.n80 9.3005
R831 VDD2.n53 VDD2.n52 9.3005
R832 VDD2.n22 VDD2.n21 9.3005
R833 VDD2.n47 VDD2.n46 9.3005
R834 VDD2.n45 VDD2.n44 9.3005
R835 VDD2.n26 VDD2.n25 9.3005
R836 VDD2.n39 VDD2.n38 9.3005
R837 VDD2.n37 VDD2.n36 9.3005
R838 VDD2.n30 VDD2.n29 9.3005
R839 VDD2.n55 VDD2.n54 9.3005
R840 VDD2.n18 VDD2.n17 9.3005
R841 VDD2.n61 VDD2.n60 9.3005
R842 VDD2.n63 VDD2.n62 9.3005
R843 VDD2.n14 VDD2.n13 9.3005
R844 VDD2.n69 VDD2.n68 9.3005
R845 VDD2.n71 VDD2.n70 9.3005
R846 VDD2.n72 VDD2.n9 9.3005
R847 VDD2.n79 VDD2.n78 9.3005
R848 VDD2.n193 VDD2.n99 8.92171
R849 VDD2.n164 VDD2.n117 8.92171
R850 VDD2.n149 VDD2.n148 8.92171
R851 VDD2.n48 VDD2.n47 8.92171
R852 VDD2.n63 VDD2.n16 8.92171
R853 VDD2.n94 VDD2.n0 8.92171
R854 VDD2.n161 VDD2.n160 8.14595
R855 VDD2.n152 VDD2.n123 8.14595
R856 VDD2.n51 VDD2.n22 8.14595
R857 VDD2.n60 VDD2.n59 8.14595
R858 VDD2.n157 VDD2.n119 7.3702
R859 VDD2.n153 VDD2.n121 7.3702
R860 VDD2.n52 VDD2.n20 7.3702
R861 VDD2.n56 VDD2.n18 7.3702
R862 VDD2.n157 VDD2.n156 6.59444
R863 VDD2.n156 VDD2.n121 6.59444
R864 VDD2.n55 VDD2.n20 6.59444
R865 VDD2.n56 VDD2.n55 6.59444
R866 VDD2.n160 VDD2.n119 5.81868
R867 VDD2.n153 VDD2.n152 5.81868
R868 VDD2.n52 VDD2.n51 5.81868
R869 VDD2.n59 VDD2.n18 5.81868
R870 VDD2.n195 VDD2.n99 5.04292
R871 VDD2.n161 VDD2.n117 5.04292
R872 VDD2.n149 VDD2.n123 5.04292
R873 VDD2.n48 VDD2.n22 5.04292
R874 VDD2.n60 VDD2.n16 5.04292
R875 VDD2.n96 VDD2.n0 5.04292
R876 VDD2.n193 VDD2.n192 4.26717
R877 VDD2.n165 VDD2.n164 4.26717
R878 VDD2.n148 VDD2.n125 4.26717
R879 VDD2.n47 VDD2.n24 4.26717
R880 VDD2.n64 VDD2.n63 4.26717
R881 VDD2.n94 VDD2.n93 4.26717
R882 VDD2.n132 VDD2.n130 3.70982
R883 VDD2.n31 VDD2.n29 3.70982
R884 VDD2.n189 VDD2.n101 3.49141
R885 VDD2.n168 VDD2.n115 3.49141
R886 VDD2.n145 VDD2.n144 3.49141
R887 VDD2.n44 VDD2.n43 3.49141
R888 VDD2.n67 VDD2.n14 3.49141
R889 VDD2.n90 VDD2.n2 3.49141
R890 VDD2.n188 VDD2.n103 2.71565
R891 VDD2.n169 VDD2.n113 2.71565
R892 VDD2.n141 VDD2.n127 2.71565
R893 VDD2.n40 VDD2.n26 2.71565
R894 VDD2.n68 VDD2.n12 2.71565
R895 VDD2.n89 VDD2.n4 2.71565
R896 VDD2 VDD2.n196 1.95955
R897 VDD2.n185 VDD2.n184 1.93989
R898 VDD2.n173 VDD2.n172 1.93989
R899 VDD2.n140 VDD2.n129 1.93989
R900 VDD2.n39 VDD2.n28 1.93989
R901 VDD2.n73 VDD2.n71 1.93989
R902 VDD2.n86 VDD2.n85 1.93989
R903 VDD2.n197 VDD2.t2 1.86218
R904 VDD2.n197 VDD2.t3 1.86218
R905 VDD2.n97 VDD2.t4 1.86218
R906 VDD2.n97 VDD2.t0 1.86218
R907 VDD2.n181 VDD2.n105 1.16414
R908 VDD2.n176 VDD2.n110 1.16414
R909 VDD2.n137 VDD2.n136 1.16414
R910 VDD2.n36 VDD2.n35 1.16414
R911 VDD2.n72 VDD2.n10 1.16414
R912 VDD2.n82 VDD2.n6 1.16414
R913 VDD2.n180 VDD2.n107 0.388379
R914 VDD2.n177 VDD2.n109 0.388379
R915 VDD2.n133 VDD2.n131 0.388379
R916 VDD2.n32 VDD2.n30 0.388379
R917 VDD2.n78 VDD2.n77 0.388379
R918 VDD2.n81 VDD2.n8 0.388379
R919 VDD2.n194 VDD2.n100 0.155672
R920 VDD2.n187 VDD2.n100 0.155672
R921 VDD2.n187 VDD2.n186 0.155672
R922 VDD2.n186 VDD2.n104 0.155672
R923 VDD2.n179 VDD2.n104 0.155672
R924 VDD2.n179 VDD2.n178 0.155672
R925 VDD2.n178 VDD2.n108 0.155672
R926 VDD2.n171 VDD2.n108 0.155672
R927 VDD2.n171 VDD2.n170 0.155672
R928 VDD2.n170 VDD2.n114 0.155672
R929 VDD2.n163 VDD2.n114 0.155672
R930 VDD2.n163 VDD2.n162 0.155672
R931 VDD2.n162 VDD2.n118 0.155672
R932 VDD2.n155 VDD2.n118 0.155672
R933 VDD2.n155 VDD2.n154 0.155672
R934 VDD2.n154 VDD2.n122 0.155672
R935 VDD2.n147 VDD2.n122 0.155672
R936 VDD2.n147 VDD2.n146 0.155672
R937 VDD2.n146 VDD2.n126 0.155672
R938 VDD2.n139 VDD2.n126 0.155672
R939 VDD2.n139 VDD2.n138 0.155672
R940 VDD2.n138 VDD2.n130 0.155672
R941 VDD2.n37 VDD2.n29 0.155672
R942 VDD2.n38 VDD2.n37 0.155672
R943 VDD2.n38 VDD2.n25 0.155672
R944 VDD2.n45 VDD2.n25 0.155672
R945 VDD2.n46 VDD2.n45 0.155672
R946 VDD2.n46 VDD2.n21 0.155672
R947 VDD2.n53 VDD2.n21 0.155672
R948 VDD2.n54 VDD2.n53 0.155672
R949 VDD2.n54 VDD2.n17 0.155672
R950 VDD2.n61 VDD2.n17 0.155672
R951 VDD2.n62 VDD2.n61 0.155672
R952 VDD2.n62 VDD2.n13 0.155672
R953 VDD2.n69 VDD2.n13 0.155672
R954 VDD2.n70 VDD2.n69 0.155672
R955 VDD2.n70 VDD2.n9 0.155672
R956 VDD2.n79 VDD2.n9 0.155672
R957 VDD2.n80 VDD2.n79 0.155672
R958 VDD2.n80 VDD2.n5 0.155672
R959 VDD2.n87 VDD2.n5 0.155672
R960 VDD2.n88 VDD2.n87 0.155672
R961 VDD2.n88 VDD2.n1 0.155672
R962 VDD2.n95 VDD2.n1 0.155672
R963 B.n470 B.n133 585
R964 B.n469 B.n468 585
R965 B.n467 B.n134 585
R966 B.n466 B.n465 585
R967 B.n464 B.n135 585
R968 B.n463 B.n462 585
R969 B.n461 B.n136 585
R970 B.n460 B.n459 585
R971 B.n458 B.n137 585
R972 B.n457 B.n456 585
R973 B.n455 B.n138 585
R974 B.n454 B.n453 585
R975 B.n452 B.n139 585
R976 B.n451 B.n450 585
R977 B.n449 B.n140 585
R978 B.n448 B.n447 585
R979 B.n446 B.n141 585
R980 B.n445 B.n444 585
R981 B.n443 B.n142 585
R982 B.n442 B.n441 585
R983 B.n440 B.n143 585
R984 B.n439 B.n438 585
R985 B.n437 B.n144 585
R986 B.n436 B.n435 585
R987 B.n434 B.n145 585
R988 B.n433 B.n432 585
R989 B.n431 B.n146 585
R990 B.n430 B.n429 585
R991 B.n428 B.n147 585
R992 B.n427 B.n426 585
R993 B.n425 B.n148 585
R994 B.n424 B.n423 585
R995 B.n422 B.n149 585
R996 B.n421 B.n420 585
R997 B.n419 B.n150 585
R998 B.n418 B.n417 585
R999 B.n416 B.n151 585
R1000 B.n415 B.n414 585
R1001 B.n413 B.n152 585
R1002 B.n412 B.n411 585
R1003 B.n410 B.n153 585
R1004 B.n409 B.n408 585
R1005 B.n407 B.n154 585
R1006 B.n406 B.n405 585
R1007 B.n404 B.n155 585
R1008 B.n403 B.n402 585
R1009 B.n401 B.n156 585
R1010 B.n400 B.n399 585
R1011 B.n398 B.n157 585
R1012 B.n397 B.n396 585
R1013 B.n395 B.n158 585
R1014 B.n394 B.n393 585
R1015 B.n392 B.n159 585
R1016 B.n391 B.n390 585
R1017 B.n389 B.n160 585
R1018 B.n388 B.n387 585
R1019 B.n386 B.n161 585
R1020 B.n385 B.n384 585
R1021 B.n383 B.n382 585
R1022 B.n381 B.n165 585
R1023 B.n380 B.n379 585
R1024 B.n378 B.n166 585
R1025 B.n377 B.n376 585
R1026 B.n375 B.n167 585
R1027 B.n374 B.n373 585
R1028 B.n372 B.n168 585
R1029 B.n371 B.n370 585
R1030 B.n368 B.n169 585
R1031 B.n367 B.n366 585
R1032 B.n365 B.n172 585
R1033 B.n364 B.n363 585
R1034 B.n362 B.n173 585
R1035 B.n361 B.n360 585
R1036 B.n359 B.n174 585
R1037 B.n358 B.n357 585
R1038 B.n356 B.n175 585
R1039 B.n355 B.n354 585
R1040 B.n353 B.n176 585
R1041 B.n352 B.n351 585
R1042 B.n350 B.n177 585
R1043 B.n349 B.n348 585
R1044 B.n347 B.n178 585
R1045 B.n346 B.n345 585
R1046 B.n344 B.n179 585
R1047 B.n343 B.n342 585
R1048 B.n341 B.n180 585
R1049 B.n340 B.n339 585
R1050 B.n338 B.n181 585
R1051 B.n337 B.n336 585
R1052 B.n335 B.n182 585
R1053 B.n334 B.n333 585
R1054 B.n332 B.n183 585
R1055 B.n331 B.n330 585
R1056 B.n329 B.n184 585
R1057 B.n328 B.n327 585
R1058 B.n326 B.n185 585
R1059 B.n325 B.n324 585
R1060 B.n323 B.n186 585
R1061 B.n322 B.n321 585
R1062 B.n320 B.n187 585
R1063 B.n319 B.n318 585
R1064 B.n317 B.n188 585
R1065 B.n316 B.n315 585
R1066 B.n314 B.n189 585
R1067 B.n313 B.n312 585
R1068 B.n311 B.n190 585
R1069 B.n310 B.n309 585
R1070 B.n308 B.n191 585
R1071 B.n307 B.n306 585
R1072 B.n305 B.n192 585
R1073 B.n304 B.n303 585
R1074 B.n302 B.n193 585
R1075 B.n301 B.n300 585
R1076 B.n299 B.n194 585
R1077 B.n298 B.n297 585
R1078 B.n296 B.n195 585
R1079 B.n295 B.n294 585
R1080 B.n293 B.n196 585
R1081 B.n292 B.n291 585
R1082 B.n290 B.n197 585
R1083 B.n289 B.n288 585
R1084 B.n287 B.n198 585
R1085 B.n286 B.n285 585
R1086 B.n284 B.n199 585
R1087 B.n283 B.n282 585
R1088 B.n472 B.n471 585
R1089 B.n473 B.n132 585
R1090 B.n475 B.n474 585
R1091 B.n476 B.n131 585
R1092 B.n478 B.n477 585
R1093 B.n479 B.n130 585
R1094 B.n481 B.n480 585
R1095 B.n482 B.n129 585
R1096 B.n484 B.n483 585
R1097 B.n485 B.n128 585
R1098 B.n487 B.n486 585
R1099 B.n488 B.n127 585
R1100 B.n490 B.n489 585
R1101 B.n491 B.n126 585
R1102 B.n493 B.n492 585
R1103 B.n494 B.n125 585
R1104 B.n496 B.n495 585
R1105 B.n497 B.n124 585
R1106 B.n499 B.n498 585
R1107 B.n500 B.n123 585
R1108 B.n502 B.n501 585
R1109 B.n503 B.n122 585
R1110 B.n505 B.n504 585
R1111 B.n506 B.n121 585
R1112 B.n508 B.n507 585
R1113 B.n509 B.n120 585
R1114 B.n511 B.n510 585
R1115 B.n512 B.n119 585
R1116 B.n514 B.n513 585
R1117 B.n515 B.n118 585
R1118 B.n517 B.n516 585
R1119 B.n518 B.n117 585
R1120 B.n520 B.n519 585
R1121 B.n521 B.n116 585
R1122 B.n523 B.n522 585
R1123 B.n524 B.n115 585
R1124 B.n526 B.n525 585
R1125 B.n527 B.n114 585
R1126 B.n529 B.n528 585
R1127 B.n530 B.n113 585
R1128 B.n532 B.n531 585
R1129 B.n533 B.n112 585
R1130 B.n535 B.n534 585
R1131 B.n536 B.n111 585
R1132 B.n538 B.n537 585
R1133 B.n539 B.n110 585
R1134 B.n541 B.n540 585
R1135 B.n542 B.n109 585
R1136 B.n544 B.n543 585
R1137 B.n545 B.n108 585
R1138 B.n547 B.n546 585
R1139 B.n548 B.n107 585
R1140 B.n550 B.n549 585
R1141 B.n551 B.n106 585
R1142 B.n553 B.n552 585
R1143 B.n554 B.n105 585
R1144 B.n556 B.n555 585
R1145 B.n557 B.n104 585
R1146 B.n559 B.n558 585
R1147 B.n560 B.n103 585
R1148 B.n562 B.n561 585
R1149 B.n563 B.n102 585
R1150 B.n565 B.n564 585
R1151 B.n566 B.n101 585
R1152 B.n568 B.n567 585
R1153 B.n569 B.n100 585
R1154 B.n571 B.n570 585
R1155 B.n572 B.n99 585
R1156 B.n574 B.n573 585
R1157 B.n575 B.n98 585
R1158 B.n577 B.n576 585
R1159 B.n578 B.n97 585
R1160 B.n580 B.n579 585
R1161 B.n581 B.n96 585
R1162 B.n583 B.n582 585
R1163 B.n584 B.n95 585
R1164 B.n586 B.n585 585
R1165 B.n587 B.n94 585
R1166 B.n589 B.n588 585
R1167 B.n590 B.n93 585
R1168 B.n592 B.n591 585
R1169 B.n593 B.n92 585
R1170 B.n595 B.n594 585
R1171 B.n596 B.n91 585
R1172 B.n598 B.n597 585
R1173 B.n599 B.n90 585
R1174 B.n788 B.n23 585
R1175 B.n787 B.n786 585
R1176 B.n785 B.n24 585
R1177 B.n784 B.n783 585
R1178 B.n782 B.n25 585
R1179 B.n781 B.n780 585
R1180 B.n779 B.n26 585
R1181 B.n778 B.n777 585
R1182 B.n776 B.n27 585
R1183 B.n775 B.n774 585
R1184 B.n773 B.n28 585
R1185 B.n772 B.n771 585
R1186 B.n770 B.n29 585
R1187 B.n769 B.n768 585
R1188 B.n767 B.n30 585
R1189 B.n766 B.n765 585
R1190 B.n764 B.n31 585
R1191 B.n763 B.n762 585
R1192 B.n761 B.n32 585
R1193 B.n760 B.n759 585
R1194 B.n758 B.n33 585
R1195 B.n757 B.n756 585
R1196 B.n755 B.n34 585
R1197 B.n754 B.n753 585
R1198 B.n752 B.n35 585
R1199 B.n751 B.n750 585
R1200 B.n749 B.n36 585
R1201 B.n748 B.n747 585
R1202 B.n746 B.n37 585
R1203 B.n745 B.n744 585
R1204 B.n743 B.n38 585
R1205 B.n742 B.n741 585
R1206 B.n740 B.n39 585
R1207 B.n739 B.n738 585
R1208 B.n737 B.n40 585
R1209 B.n736 B.n735 585
R1210 B.n734 B.n41 585
R1211 B.n733 B.n732 585
R1212 B.n731 B.n42 585
R1213 B.n730 B.n729 585
R1214 B.n728 B.n43 585
R1215 B.n727 B.n726 585
R1216 B.n725 B.n44 585
R1217 B.n724 B.n723 585
R1218 B.n722 B.n45 585
R1219 B.n721 B.n720 585
R1220 B.n719 B.n46 585
R1221 B.n718 B.n717 585
R1222 B.n716 B.n47 585
R1223 B.n715 B.n714 585
R1224 B.n713 B.n48 585
R1225 B.n712 B.n711 585
R1226 B.n710 B.n49 585
R1227 B.n709 B.n708 585
R1228 B.n707 B.n50 585
R1229 B.n706 B.n705 585
R1230 B.n704 B.n51 585
R1231 B.n703 B.n702 585
R1232 B.n701 B.n700 585
R1233 B.n699 B.n55 585
R1234 B.n698 B.n697 585
R1235 B.n696 B.n56 585
R1236 B.n695 B.n694 585
R1237 B.n693 B.n57 585
R1238 B.n692 B.n691 585
R1239 B.n690 B.n58 585
R1240 B.n689 B.n688 585
R1241 B.n686 B.n59 585
R1242 B.n685 B.n684 585
R1243 B.n683 B.n62 585
R1244 B.n682 B.n681 585
R1245 B.n680 B.n63 585
R1246 B.n679 B.n678 585
R1247 B.n677 B.n64 585
R1248 B.n676 B.n675 585
R1249 B.n674 B.n65 585
R1250 B.n673 B.n672 585
R1251 B.n671 B.n66 585
R1252 B.n670 B.n669 585
R1253 B.n668 B.n67 585
R1254 B.n667 B.n666 585
R1255 B.n665 B.n68 585
R1256 B.n664 B.n663 585
R1257 B.n662 B.n69 585
R1258 B.n661 B.n660 585
R1259 B.n659 B.n70 585
R1260 B.n658 B.n657 585
R1261 B.n656 B.n71 585
R1262 B.n655 B.n654 585
R1263 B.n653 B.n72 585
R1264 B.n652 B.n651 585
R1265 B.n650 B.n73 585
R1266 B.n649 B.n648 585
R1267 B.n647 B.n74 585
R1268 B.n646 B.n645 585
R1269 B.n644 B.n75 585
R1270 B.n643 B.n642 585
R1271 B.n641 B.n76 585
R1272 B.n640 B.n639 585
R1273 B.n638 B.n77 585
R1274 B.n637 B.n636 585
R1275 B.n635 B.n78 585
R1276 B.n634 B.n633 585
R1277 B.n632 B.n79 585
R1278 B.n631 B.n630 585
R1279 B.n629 B.n80 585
R1280 B.n628 B.n627 585
R1281 B.n626 B.n81 585
R1282 B.n625 B.n624 585
R1283 B.n623 B.n82 585
R1284 B.n622 B.n621 585
R1285 B.n620 B.n83 585
R1286 B.n619 B.n618 585
R1287 B.n617 B.n84 585
R1288 B.n616 B.n615 585
R1289 B.n614 B.n85 585
R1290 B.n613 B.n612 585
R1291 B.n611 B.n86 585
R1292 B.n610 B.n609 585
R1293 B.n608 B.n87 585
R1294 B.n607 B.n606 585
R1295 B.n605 B.n88 585
R1296 B.n604 B.n603 585
R1297 B.n602 B.n89 585
R1298 B.n601 B.n600 585
R1299 B.n790 B.n789 585
R1300 B.n791 B.n22 585
R1301 B.n793 B.n792 585
R1302 B.n794 B.n21 585
R1303 B.n796 B.n795 585
R1304 B.n797 B.n20 585
R1305 B.n799 B.n798 585
R1306 B.n800 B.n19 585
R1307 B.n802 B.n801 585
R1308 B.n803 B.n18 585
R1309 B.n805 B.n804 585
R1310 B.n806 B.n17 585
R1311 B.n808 B.n807 585
R1312 B.n809 B.n16 585
R1313 B.n811 B.n810 585
R1314 B.n812 B.n15 585
R1315 B.n814 B.n813 585
R1316 B.n815 B.n14 585
R1317 B.n817 B.n816 585
R1318 B.n818 B.n13 585
R1319 B.n820 B.n819 585
R1320 B.n821 B.n12 585
R1321 B.n823 B.n822 585
R1322 B.n824 B.n11 585
R1323 B.n826 B.n825 585
R1324 B.n827 B.n10 585
R1325 B.n829 B.n828 585
R1326 B.n830 B.n9 585
R1327 B.n832 B.n831 585
R1328 B.n833 B.n8 585
R1329 B.n835 B.n834 585
R1330 B.n836 B.n7 585
R1331 B.n838 B.n837 585
R1332 B.n839 B.n6 585
R1333 B.n841 B.n840 585
R1334 B.n842 B.n5 585
R1335 B.n844 B.n843 585
R1336 B.n845 B.n4 585
R1337 B.n847 B.n846 585
R1338 B.n848 B.n3 585
R1339 B.n850 B.n849 585
R1340 B.n851 B.n0 585
R1341 B.n2 B.n1 585
R1342 B.n221 B.n220 585
R1343 B.n223 B.n222 585
R1344 B.n224 B.n219 585
R1345 B.n226 B.n225 585
R1346 B.n227 B.n218 585
R1347 B.n229 B.n228 585
R1348 B.n230 B.n217 585
R1349 B.n232 B.n231 585
R1350 B.n233 B.n216 585
R1351 B.n235 B.n234 585
R1352 B.n236 B.n215 585
R1353 B.n238 B.n237 585
R1354 B.n239 B.n214 585
R1355 B.n241 B.n240 585
R1356 B.n242 B.n213 585
R1357 B.n244 B.n243 585
R1358 B.n245 B.n212 585
R1359 B.n247 B.n246 585
R1360 B.n248 B.n211 585
R1361 B.n250 B.n249 585
R1362 B.n251 B.n210 585
R1363 B.n253 B.n252 585
R1364 B.n254 B.n209 585
R1365 B.n256 B.n255 585
R1366 B.n257 B.n208 585
R1367 B.n259 B.n258 585
R1368 B.n260 B.n207 585
R1369 B.n262 B.n261 585
R1370 B.n263 B.n206 585
R1371 B.n265 B.n264 585
R1372 B.n266 B.n205 585
R1373 B.n268 B.n267 585
R1374 B.n269 B.n204 585
R1375 B.n271 B.n270 585
R1376 B.n272 B.n203 585
R1377 B.n274 B.n273 585
R1378 B.n275 B.n202 585
R1379 B.n277 B.n276 585
R1380 B.n278 B.n201 585
R1381 B.n280 B.n279 585
R1382 B.n281 B.n200 585
R1383 B.n162 B.t1 530.919
R1384 B.n60 B.t11 530.919
R1385 B.n170 B.t4 530.919
R1386 B.n52 B.t8 530.919
R1387 B.n282 B.n281 526.135
R1388 B.n472 B.n133 526.135
R1389 B.n600 B.n599 526.135
R1390 B.n790 B.n23 526.135
R1391 B.n163 B.t2 473.901
R1392 B.n61 B.t10 473.901
R1393 B.n171 B.t5 473.901
R1394 B.n53 B.t7 473.901
R1395 B.n170 B.t3 369.283
R1396 B.n162 B.t0 369.283
R1397 B.n60 B.t9 369.283
R1398 B.n52 B.t6 369.283
R1399 B.n853 B.n852 256.663
R1400 B.n852 B.n851 235.042
R1401 B.n852 B.n2 235.042
R1402 B.n282 B.n199 163.367
R1403 B.n286 B.n199 163.367
R1404 B.n287 B.n286 163.367
R1405 B.n288 B.n287 163.367
R1406 B.n288 B.n197 163.367
R1407 B.n292 B.n197 163.367
R1408 B.n293 B.n292 163.367
R1409 B.n294 B.n293 163.367
R1410 B.n294 B.n195 163.367
R1411 B.n298 B.n195 163.367
R1412 B.n299 B.n298 163.367
R1413 B.n300 B.n299 163.367
R1414 B.n300 B.n193 163.367
R1415 B.n304 B.n193 163.367
R1416 B.n305 B.n304 163.367
R1417 B.n306 B.n305 163.367
R1418 B.n306 B.n191 163.367
R1419 B.n310 B.n191 163.367
R1420 B.n311 B.n310 163.367
R1421 B.n312 B.n311 163.367
R1422 B.n312 B.n189 163.367
R1423 B.n316 B.n189 163.367
R1424 B.n317 B.n316 163.367
R1425 B.n318 B.n317 163.367
R1426 B.n318 B.n187 163.367
R1427 B.n322 B.n187 163.367
R1428 B.n323 B.n322 163.367
R1429 B.n324 B.n323 163.367
R1430 B.n324 B.n185 163.367
R1431 B.n328 B.n185 163.367
R1432 B.n329 B.n328 163.367
R1433 B.n330 B.n329 163.367
R1434 B.n330 B.n183 163.367
R1435 B.n334 B.n183 163.367
R1436 B.n335 B.n334 163.367
R1437 B.n336 B.n335 163.367
R1438 B.n336 B.n181 163.367
R1439 B.n340 B.n181 163.367
R1440 B.n341 B.n340 163.367
R1441 B.n342 B.n341 163.367
R1442 B.n342 B.n179 163.367
R1443 B.n346 B.n179 163.367
R1444 B.n347 B.n346 163.367
R1445 B.n348 B.n347 163.367
R1446 B.n348 B.n177 163.367
R1447 B.n352 B.n177 163.367
R1448 B.n353 B.n352 163.367
R1449 B.n354 B.n353 163.367
R1450 B.n354 B.n175 163.367
R1451 B.n358 B.n175 163.367
R1452 B.n359 B.n358 163.367
R1453 B.n360 B.n359 163.367
R1454 B.n360 B.n173 163.367
R1455 B.n364 B.n173 163.367
R1456 B.n365 B.n364 163.367
R1457 B.n366 B.n365 163.367
R1458 B.n366 B.n169 163.367
R1459 B.n371 B.n169 163.367
R1460 B.n372 B.n371 163.367
R1461 B.n373 B.n372 163.367
R1462 B.n373 B.n167 163.367
R1463 B.n377 B.n167 163.367
R1464 B.n378 B.n377 163.367
R1465 B.n379 B.n378 163.367
R1466 B.n379 B.n165 163.367
R1467 B.n383 B.n165 163.367
R1468 B.n384 B.n383 163.367
R1469 B.n384 B.n161 163.367
R1470 B.n388 B.n161 163.367
R1471 B.n389 B.n388 163.367
R1472 B.n390 B.n389 163.367
R1473 B.n390 B.n159 163.367
R1474 B.n394 B.n159 163.367
R1475 B.n395 B.n394 163.367
R1476 B.n396 B.n395 163.367
R1477 B.n396 B.n157 163.367
R1478 B.n400 B.n157 163.367
R1479 B.n401 B.n400 163.367
R1480 B.n402 B.n401 163.367
R1481 B.n402 B.n155 163.367
R1482 B.n406 B.n155 163.367
R1483 B.n407 B.n406 163.367
R1484 B.n408 B.n407 163.367
R1485 B.n408 B.n153 163.367
R1486 B.n412 B.n153 163.367
R1487 B.n413 B.n412 163.367
R1488 B.n414 B.n413 163.367
R1489 B.n414 B.n151 163.367
R1490 B.n418 B.n151 163.367
R1491 B.n419 B.n418 163.367
R1492 B.n420 B.n419 163.367
R1493 B.n420 B.n149 163.367
R1494 B.n424 B.n149 163.367
R1495 B.n425 B.n424 163.367
R1496 B.n426 B.n425 163.367
R1497 B.n426 B.n147 163.367
R1498 B.n430 B.n147 163.367
R1499 B.n431 B.n430 163.367
R1500 B.n432 B.n431 163.367
R1501 B.n432 B.n145 163.367
R1502 B.n436 B.n145 163.367
R1503 B.n437 B.n436 163.367
R1504 B.n438 B.n437 163.367
R1505 B.n438 B.n143 163.367
R1506 B.n442 B.n143 163.367
R1507 B.n443 B.n442 163.367
R1508 B.n444 B.n443 163.367
R1509 B.n444 B.n141 163.367
R1510 B.n448 B.n141 163.367
R1511 B.n449 B.n448 163.367
R1512 B.n450 B.n449 163.367
R1513 B.n450 B.n139 163.367
R1514 B.n454 B.n139 163.367
R1515 B.n455 B.n454 163.367
R1516 B.n456 B.n455 163.367
R1517 B.n456 B.n137 163.367
R1518 B.n460 B.n137 163.367
R1519 B.n461 B.n460 163.367
R1520 B.n462 B.n461 163.367
R1521 B.n462 B.n135 163.367
R1522 B.n466 B.n135 163.367
R1523 B.n467 B.n466 163.367
R1524 B.n468 B.n467 163.367
R1525 B.n468 B.n133 163.367
R1526 B.n599 B.n598 163.367
R1527 B.n598 B.n91 163.367
R1528 B.n594 B.n91 163.367
R1529 B.n594 B.n593 163.367
R1530 B.n593 B.n592 163.367
R1531 B.n592 B.n93 163.367
R1532 B.n588 B.n93 163.367
R1533 B.n588 B.n587 163.367
R1534 B.n587 B.n586 163.367
R1535 B.n586 B.n95 163.367
R1536 B.n582 B.n95 163.367
R1537 B.n582 B.n581 163.367
R1538 B.n581 B.n580 163.367
R1539 B.n580 B.n97 163.367
R1540 B.n576 B.n97 163.367
R1541 B.n576 B.n575 163.367
R1542 B.n575 B.n574 163.367
R1543 B.n574 B.n99 163.367
R1544 B.n570 B.n99 163.367
R1545 B.n570 B.n569 163.367
R1546 B.n569 B.n568 163.367
R1547 B.n568 B.n101 163.367
R1548 B.n564 B.n101 163.367
R1549 B.n564 B.n563 163.367
R1550 B.n563 B.n562 163.367
R1551 B.n562 B.n103 163.367
R1552 B.n558 B.n103 163.367
R1553 B.n558 B.n557 163.367
R1554 B.n557 B.n556 163.367
R1555 B.n556 B.n105 163.367
R1556 B.n552 B.n105 163.367
R1557 B.n552 B.n551 163.367
R1558 B.n551 B.n550 163.367
R1559 B.n550 B.n107 163.367
R1560 B.n546 B.n107 163.367
R1561 B.n546 B.n545 163.367
R1562 B.n545 B.n544 163.367
R1563 B.n544 B.n109 163.367
R1564 B.n540 B.n109 163.367
R1565 B.n540 B.n539 163.367
R1566 B.n539 B.n538 163.367
R1567 B.n538 B.n111 163.367
R1568 B.n534 B.n111 163.367
R1569 B.n534 B.n533 163.367
R1570 B.n533 B.n532 163.367
R1571 B.n532 B.n113 163.367
R1572 B.n528 B.n113 163.367
R1573 B.n528 B.n527 163.367
R1574 B.n527 B.n526 163.367
R1575 B.n526 B.n115 163.367
R1576 B.n522 B.n115 163.367
R1577 B.n522 B.n521 163.367
R1578 B.n521 B.n520 163.367
R1579 B.n520 B.n117 163.367
R1580 B.n516 B.n117 163.367
R1581 B.n516 B.n515 163.367
R1582 B.n515 B.n514 163.367
R1583 B.n514 B.n119 163.367
R1584 B.n510 B.n119 163.367
R1585 B.n510 B.n509 163.367
R1586 B.n509 B.n508 163.367
R1587 B.n508 B.n121 163.367
R1588 B.n504 B.n121 163.367
R1589 B.n504 B.n503 163.367
R1590 B.n503 B.n502 163.367
R1591 B.n502 B.n123 163.367
R1592 B.n498 B.n123 163.367
R1593 B.n498 B.n497 163.367
R1594 B.n497 B.n496 163.367
R1595 B.n496 B.n125 163.367
R1596 B.n492 B.n125 163.367
R1597 B.n492 B.n491 163.367
R1598 B.n491 B.n490 163.367
R1599 B.n490 B.n127 163.367
R1600 B.n486 B.n127 163.367
R1601 B.n486 B.n485 163.367
R1602 B.n485 B.n484 163.367
R1603 B.n484 B.n129 163.367
R1604 B.n480 B.n129 163.367
R1605 B.n480 B.n479 163.367
R1606 B.n479 B.n478 163.367
R1607 B.n478 B.n131 163.367
R1608 B.n474 B.n131 163.367
R1609 B.n474 B.n473 163.367
R1610 B.n473 B.n472 163.367
R1611 B.n786 B.n23 163.367
R1612 B.n786 B.n785 163.367
R1613 B.n785 B.n784 163.367
R1614 B.n784 B.n25 163.367
R1615 B.n780 B.n25 163.367
R1616 B.n780 B.n779 163.367
R1617 B.n779 B.n778 163.367
R1618 B.n778 B.n27 163.367
R1619 B.n774 B.n27 163.367
R1620 B.n774 B.n773 163.367
R1621 B.n773 B.n772 163.367
R1622 B.n772 B.n29 163.367
R1623 B.n768 B.n29 163.367
R1624 B.n768 B.n767 163.367
R1625 B.n767 B.n766 163.367
R1626 B.n766 B.n31 163.367
R1627 B.n762 B.n31 163.367
R1628 B.n762 B.n761 163.367
R1629 B.n761 B.n760 163.367
R1630 B.n760 B.n33 163.367
R1631 B.n756 B.n33 163.367
R1632 B.n756 B.n755 163.367
R1633 B.n755 B.n754 163.367
R1634 B.n754 B.n35 163.367
R1635 B.n750 B.n35 163.367
R1636 B.n750 B.n749 163.367
R1637 B.n749 B.n748 163.367
R1638 B.n748 B.n37 163.367
R1639 B.n744 B.n37 163.367
R1640 B.n744 B.n743 163.367
R1641 B.n743 B.n742 163.367
R1642 B.n742 B.n39 163.367
R1643 B.n738 B.n39 163.367
R1644 B.n738 B.n737 163.367
R1645 B.n737 B.n736 163.367
R1646 B.n736 B.n41 163.367
R1647 B.n732 B.n41 163.367
R1648 B.n732 B.n731 163.367
R1649 B.n731 B.n730 163.367
R1650 B.n730 B.n43 163.367
R1651 B.n726 B.n43 163.367
R1652 B.n726 B.n725 163.367
R1653 B.n725 B.n724 163.367
R1654 B.n724 B.n45 163.367
R1655 B.n720 B.n45 163.367
R1656 B.n720 B.n719 163.367
R1657 B.n719 B.n718 163.367
R1658 B.n718 B.n47 163.367
R1659 B.n714 B.n47 163.367
R1660 B.n714 B.n713 163.367
R1661 B.n713 B.n712 163.367
R1662 B.n712 B.n49 163.367
R1663 B.n708 B.n49 163.367
R1664 B.n708 B.n707 163.367
R1665 B.n707 B.n706 163.367
R1666 B.n706 B.n51 163.367
R1667 B.n702 B.n51 163.367
R1668 B.n702 B.n701 163.367
R1669 B.n701 B.n55 163.367
R1670 B.n697 B.n55 163.367
R1671 B.n697 B.n696 163.367
R1672 B.n696 B.n695 163.367
R1673 B.n695 B.n57 163.367
R1674 B.n691 B.n57 163.367
R1675 B.n691 B.n690 163.367
R1676 B.n690 B.n689 163.367
R1677 B.n689 B.n59 163.367
R1678 B.n684 B.n59 163.367
R1679 B.n684 B.n683 163.367
R1680 B.n683 B.n682 163.367
R1681 B.n682 B.n63 163.367
R1682 B.n678 B.n63 163.367
R1683 B.n678 B.n677 163.367
R1684 B.n677 B.n676 163.367
R1685 B.n676 B.n65 163.367
R1686 B.n672 B.n65 163.367
R1687 B.n672 B.n671 163.367
R1688 B.n671 B.n670 163.367
R1689 B.n670 B.n67 163.367
R1690 B.n666 B.n67 163.367
R1691 B.n666 B.n665 163.367
R1692 B.n665 B.n664 163.367
R1693 B.n664 B.n69 163.367
R1694 B.n660 B.n69 163.367
R1695 B.n660 B.n659 163.367
R1696 B.n659 B.n658 163.367
R1697 B.n658 B.n71 163.367
R1698 B.n654 B.n71 163.367
R1699 B.n654 B.n653 163.367
R1700 B.n653 B.n652 163.367
R1701 B.n652 B.n73 163.367
R1702 B.n648 B.n73 163.367
R1703 B.n648 B.n647 163.367
R1704 B.n647 B.n646 163.367
R1705 B.n646 B.n75 163.367
R1706 B.n642 B.n75 163.367
R1707 B.n642 B.n641 163.367
R1708 B.n641 B.n640 163.367
R1709 B.n640 B.n77 163.367
R1710 B.n636 B.n77 163.367
R1711 B.n636 B.n635 163.367
R1712 B.n635 B.n634 163.367
R1713 B.n634 B.n79 163.367
R1714 B.n630 B.n79 163.367
R1715 B.n630 B.n629 163.367
R1716 B.n629 B.n628 163.367
R1717 B.n628 B.n81 163.367
R1718 B.n624 B.n81 163.367
R1719 B.n624 B.n623 163.367
R1720 B.n623 B.n622 163.367
R1721 B.n622 B.n83 163.367
R1722 B.n618 B.n83 163.367
R1723 B.n618 B.n617 163.367
R1724 B.n617 B.n616 163.367
R1725 B.n616 B.n85 163.367
R1726 B.n612 B.n85 163.367
R1727 B.n612 B.n611 163.367
R1728 B.n611 B.n610 163.367
R1729 B.n610 B.n87 163.367
R1730 B.n606 B.n87 163.367
R1731 B.n606 B.n605 163.367
R1732 B.n605 B.n604 163.367
R1733 B.n604 B.n89 163.367
R1734 B.n600 B.n89 163.367
R1735 B.n791 B.n790 163.367
R1736 B.n792 B.n791 163.367
R1737 B.n792 B.n21 163.367
R1738 B.n796 B.n21 163.367
R1739 B.n797 B.n796 163.367
R1740 B.n798 B.n797 163.367
R1741 B.n798 B.n19 163.367
R1742 B.n802 B.n19 163.367
R1743 B.n803 B.n802 163.367
R1744 B.n804 B.n803 163.367
R1745 B.n804 B.n17 163.367
R1746 B.n808 B.n17 163.367
R1747 B.n809 B.n808 163.367
R1748 B.n810 B.n809 163.367
R1749 B.n810 B.n15 163.367
R1750 B.n814 B.n15 163.367
R1751 B.n815 B.n814 163.367
R1752 B.n816 B.n815 163.367
R1753 B.n816 B.n13 163.367
R1754 B.n820 B.n13 163.367
R1755 B.n821 B.n820 163.367
R1756 B.n822 B.n821 163.367
R1757 B.n822 B.n11 163.367
R1758 B.n826 B.n11 163.367
R1759 B.n827 B.n826 163.367
R1760 B.n828 B.n827 163.367
R1761 B.n828 B.n9 163.367
R1762 B.n832 B.n9 163.367
R1763 B.n833 B.n832 163.367
R1764 B.n834 B.n833 163.367
R1765 B.n834 B.n7 163.367
R1766 B.n838 B.n7 163.367
R1767 B.n839 B.n838 163.367
R1768 B.n840 B.n839 163.367
R1769 B.n840 B.n5 163.367
R1770 B.n844 B.n5 163.367
R1771 B.n845 B.n844 163.367
R1772 B.n846 B.n845 163.367
R1773 B.n846 B.n3 163.367
R1774 B.n850 B.n3 163.367
R1775 B.n851 B.n850 163.367
R1776 B.n221 B.n2 163.367
R1777 B.n222 B.n221 163.367
R1778 B.n222 B.n219 163.367
R1779 B.n226 B.n219 163.367
R1780 B.n227 B.n226 163.367
R1781 B.n228 B.n227 163.367
R1782 B.n228 B.n217 163.367
R1783 B.n232 B.n217 163.367
R1784 B.n233 B.n232 163.367
R1785 B.n234 B.n233 163.367
R1786 B.n234 B.n215 163.367
R1787 B.n238 B.n215 163.367
R1788 B.n239 B.n238 163.367
R1789 B.n240 B.n239 163.367
R1790 B.n240 B.n213 163.367
R1791 B.n244 B.n213 163.367
R1792 B.n245 B.n244 163.367
R1793 B.n246 B.n245 163.367
R1794 B.n246 B.n211 163.367
R1795 B.n250 B.n211 163.367
R1796 B.n251 B.n250 163.367
R1797 B.n252 B.n251 163.367
R1798 B.n252 B.n209 163.367
R1799 B.n256 B.n209 163.367
R1800 B.n257 B.n256 163.367
R1801 B.n258 B.n257 163.367
R1802 B.n258 B.n207 163.367
R1803 B.n262 B.n207 163.367
R1804 B.n263 B.n262 163.367
R1805 B.n264 B.n263 163.367
R1806 B.n264 B.n205 163.367
R1807 B.n268 B.n205 163.367
R1808 B.n269 B.n268 163.367
R1809 B.n270 B.n269 163.367
R1810 B.n270 B.n203 163.367
R1811 B.n274 B.n203 163.367
R1812 B.n275 B.n274 163.367
R1813 B.n276 B.n275 163.367
R1814 B.n276 B.n201 163.367
R1815 B.n280 B.n201 163.367
R1816 B.n281 B.n280 163.367
R1817 B.n369 B.n171 59.5399
R1818 B.n164 B.n163 59.5399
R1819 B.n687 B.n61 59.5399
R1820 B.n54 B.n53 59.5399
R1821 B.n171 B.n170 57.0187
R1822 B.n163 B.n162 57.0187
R1823 B.n61 B.n60 57.0187
R1824 B.n53 B.n52 57.0187
R1825 B.n789 B.n788 34.1859
R1826 B.n601 B.n90 34.1859
R1827 B.n471 B.n470 34.1859
R1828 B.n283 B.n200 34.1859
R1829 B B.n853 18.0485
R1830 B.n789 B.n22 10.6151
R1831 B.n793 B.n22 10.6151
R1832 B.n794 B.n793 10.6151
R1833 B.n795 B.n794 10.6151
R1834 B.n795 B.n20 10.6151
R1835 B.n799 B.n20 10.6151
R1836 B.n800 B.n799 10.6151
R1837 B.n801 B.n800 10.6151
R1838 B.n801 B.n18 10.6151
R1839 B.n805 B.n18 10.6151
R1840 B.n806 B.n805 10.6151
R1841 B.n807 B.n806 10.6151
R1842 B.n807 B.n16 10.6151
R1843 B.n811 B.n16 10.6151
R1844 B.n812 B.n811 10.6151
R1845 B.n813 B.n812 10.6151
R1846 B.n813 B.n14 10.6151
R1847 B.n817 B.n14 10.6151
R1848 B.n818 B.n817 10.6151
R1849 B.n819 B.n818 10.6151
R1850 B.n819 B.n12 10.6151
R1851 B.n823 B.n12 10.6151
R1852 B.n824 B.n823 10.6151
R1853 B.n825 B.n824 10.6151
R1854 B.n825 B.n10 10.6151
R1855 B.n829 B.n10 10.6151
R1856 B.n830 B.n829 10.6151
R1857 B.n831 B.n830 10.6151
R1858 B.n831 B.n8 10.6151
R1859 B.n835 B.n8 10.6151
R1860 B.n836 B.n835 10.6151
R1861 B.n837 B.n836 10.6151
R1862 B.n837 B.n6 10.6151
R1863 B.n841 B.n6 10.6151
R1864 B.n842 B.n841 10.6151
R1865 B.n843 B.n842 10.6151
R1866 B.n843 B.n4 10.6151
R1867 B.n847 B.n4 10.6151
R1868 B.n848 B.n847 10.6151
R1869 B.n849 B.n848 10.6151
R1870 B.n849 B.n0 10.6151
R1871 B.n788 B.n787 10.6151
R1872 B.n787 B.n24 10.6151
R1873 B.n783 B.n24 10.6151
R1874 B.n783 B.n782 10.6151
R1875 B.n782 B.n781 10.6151
R1876 B.n781 B.n26 10.6151
R1877 B.n777 B.n26 10.6151
R1878 B.n777 B.n776 10.6151
R1879 B.n776 B.n775 10.6151
R1880 B.n775 B.n28 10.6151
R1881 B.n771 B.n28 10.6151
R1882 B.n771 B.n770 10.6151
R1883 B.n770 B.n769 10.6151
R1884 B.n769 B.n30 10.6151
R1885 B.n765 B.n30 10.6151
R1886 B.n765 B.n764 10.6151
R1887 B.n764 B.n763 10.6151
R1888 B.n763 B.n32 10.6151
R1889 B.n759 B.n32 10.6151
R1890 B.n759 B.n758 10.6151
R1891 B.n758 B.n757 10.6151
R1892 B.n757 B.n34 10.6151
R1893 B.n753 B.n34 10.6151
R1894 B.n753 B.n752 10.6151
R1895 B.n752 B.n751 10.6151
R1896 B.n751 B.n36 10.6151
R1897 B.n747 B.n36 10.6151
R1898 B.n747 B.n746 10.6151
R1899 B.n746 B.n745 10.6151
R1900 B.n745 B.n38 10.6151
R1901 B.n741 B.n38 10.6151
R1902 B.n741 B.n740 10.6151
R1903 B.n740 B.n739 10.6151
R1904 B.n739 B.n40 10.6151
R1905 B.n735 B.n40 10.6151
R1906 B.n735 B.n734 10.6151
R1907 B.n734 B.n733 10.6151
R1908 B.n733 B.n42 10.6151
R1909 B.n729 B.n42 10.6151
R1910 B.n729 B.n728 10.6151
R1911 B.n728 B.n727 10.6151
R1912 B.n727 B.n44 10.6151
R1913 B.n723 B.n44 10.6151
R1914 B.n723 B.n722 10.6151
R1915 B.n722 B.n721 10.6151
R1916 B.n721 B.n46 10.6151
R1917 B.n717 B.n46 10.6151
R1918 B.n717 B.n716 10.6151
R1919 B.n716 B.n715 10.6151
R1920 B.n715 B.n48 10.6151
R1921 B.n711 B.n48 10.6151
R1922 B.n711 B.n710 10.6151
R1923 B.n710 B.n709 10.6151
R1924 B.n709 B.n50 10.6151
R1925 B.n705 B.n50 10.6151
R1926 B.n705 B.n704 10.6151
R1927 B.n704 B.n703 10.6151
R1928 B.n700 B.n699 10.6151
R1929 B.n699 B.n698 10.6151
R1930 B.n698 B.n56 10.6151
R1931 B.n694 B.n56 10.6151
R1932 B.n694 B.n693 10.6151
R1933 B.n693 B.n692 10.6151
R1934 B.n692 B.n58 10.6151
R1935 B.n688 B.n58 10.6151
R1936 B.n686 B.n685 10.6151
R1937 B.n685 B.n62 10.6151
R1938 B.n681 B.n62 10.6151
R1939 B.n681 B.n680 10.6151
R1940 B.n680 B.n679 10.6151
R1941 B.n679 B.n64 10.6151
R1942 B.n675 B.n64 10.6151
R1943 B.n675 B.n674 10.6151
R1944 B.n674 B.n673 10.6151
R1945 B.n673 B.n66 10.6151
R1946 B.n669 B.n66 10.6151
R1947 B.n669 B.n668 10.6151
R1948 B.n668 B.n667 10.6151
R1949 B.n667 B.n68 10.6151
R1950 B.n663 B.n68 10.6151
R1951 B.n663 B.n662 10.6151
R1952 B.n662 B.n661 10.6151
R1953 B.n661 B.n70 10.6151
R1954 B.n657 B.n70 10.6151
R1955 B.n657 B.n656 10.6151
R1956 B.n656 B.n655 10.6151
R1957 B.n655 B.n72 10.6151
R1958 B.n651 B.n72 10.6151
R1959 B.n651 B.n650 10.6151
R1960 B.n650 B.n649 10.6151
R1961 B.n649 B.n74 10.6151
R1962 B.n645 B.n74 10.6151
R1963 B.n645 B.n644 10.6151
R1964 B.n644 B.n643 10.6151
R1965 B.n643 B.n76 10.6151
R1966 B.n639 B.n76 10.6151
R1967 B.n639 B.n638 10.6151
R1968 B.n638 B.n637 10.6151
R1969 B.n637 B.n78 10.6151
R1970 B.n633 B.n78 10.6151
R1971 B.n633 B.n632 10.6151
R1972 B.n632 B.n631 10.6151
R1973 B.n631 B.n80 10.6151
R1974 B.n627 B.n80 10.6151
R1975 B.n627 B.n626 10.6151
R1976 B.n626 B.n625 10.6151
R1977 B.n625 B.n82 10.6151
R1978 B.n621 B.n82 10.6151
R1979 B.n621 B.n620 10.6151
R1980 B.n620 B.n619 10.6151
R1981 B.n619 B.n84 10.6151
R1982 B.n615 B.n84 10.6151
R1983 B.n615 B.n614 10.6151
R1984 B.n614 B.n613 10.6151
R1985 B.n613 B.n86 10.6151
R1986 B.n609 B.n86 10.6151
R1987 B.n609 B.n608 10.6151
R1988 B.n608 B.n607 10.6151
R1989 B.n607 B.n88 10.6151
R1990 B.n603 B.n88 10.6151
R1991 B.n603 B.n602 10.6151
R1992 B.n602 B.n601 10.6151
R1993 B.n597 B.n90 10.6151
R1994 B.n597 B.n596 10.6151
R1995 B.n596 B.n595 10.6151
R1996 B.n595 B.n92 10.6151
R1997 B.n591 B.n92 10.6151
R1998 B.n591 B.n590 10.6151
R1999 B.n590 B.n589 10.6151
R2000 B.n589 B.n94 10.6151
R2001 B.n585 B.n94 10.6151
R2002 B.n585 B.n584 10.6151
R2003 B.n584 B.n583 10.6151
R2004 B.n583 B.n96 10.6151
R2005 B.n579 B.n96 10.6151
R2006 B.n579 B.n578 10.6151
R2007 B.n578 B.n577 10.6151
R2008 B.n577 B.n98 10.6151
R2009 B.n573 B.n98 10.6151
R2010 B.n573 B.n572 10.6151
R2011 B.n572 B.n571 10.6151
R2012 B.n571 B.n100 10.6151
R2013 B.n567 B.n100 10.6151
R2014 B.n567 B.n566 10.6151
R2015 B.n566 B.n565 10.6151
R2016 B.n565 B.n102 10.6151
R2017 B.n561 B.n102 10.6151
R2018 B.n561 B.n560 10.6151
R2019 B.n560 B.n559 10.6151
R2020 B.n559 B.n104 10.6151
R2021 B.n555 B.n104 10.6151
R2022 B.n555 B.n554 10.6151
R2023 B.n554 B.n553 10.6151
R2024 B.n553 B.n106 10.6151
R2025 B.n549 B.n106 10.6151
R2026 B.n549 B.n548 10.6151
R2027 B.n548 B.n547 10.6151
R2028 B.n547 B.n108 10.6151
R2029 B.n543 B.n108 10.6151
R2030 B.n543 B.n542 10.6151
R2031 B.n542 B.n541 10.6151
R2032 B.n541 B.n110 10.6151
R2033 B.n537 B.n110 10.6151
R2034 B.n537 B.n536 10.6151
R2035 B.n536 B.n535 10.6151
R2036 B.n535 B.n112 10.6151
R2037 B.n531 B.n112 10.6151
R2038 B.n531 B.n530 10.6151
R2039 B.n530 B.n529 10.6151
R2040 B.n529 B.n114 10.6151
R2041 B.n525 B.n114 10.6151
R2042 B.n525 B.n524 10.6151
R2043 B.n524 B.n523 10.6151
R2044 B.n523 B.n116 10.6151
R2045 B.n519 B.n116 10.6151
R2046 B.n519 B.n518 10.6151
R2047 B.n518 B.n517 10.6151
R2048 B.n517 B.n118 10.6151
R2049 B.n513 B.n118 10.6151
R2050 B.n513 B.n512 10.6151
R2051 B.n512 B.n511 10.6151
R2052 B.n511 B.n120 10.6151
R2053 B.n507 B.n120 10.6151
R2054 B.n507 B.n506 10.6151
R2055 B.n506 B.n505 10.6151
R2056 B.n505 B.n122 10.6151
R2057 B.n501 B.n122 10.6151
R2058 B.n501 B.n500 10.6151
R2059 B.n500 B.n499 10.6151
R2060 B.n499 B.n124 10.6151
R2061 B.n495 B.n124 10.6151
R2062 B.n495 B.n494 10.6151
R2063 B.n494 B.n493 10.6151
R2064 B.n493 B.n126 10.6151
R2065 B.n489 B.n126 10.6151
R2066 B.n489 B.n488 10.6151
R2067 B.n488 B.n487 10.6151
R2068 B.n487 B.n128 10.6151
R2069 B.n483 B.n128 10.6151
R2070 B.n483 B.n482 10.6151
R2071 B.n482 B.n481 10.6151
R2072 B.n481 B.n130 10.6151
R2073 B.n477 B.n130 10.6151
R2074 B.n477 B.n476 10.6151
R2075 B.n476 B.n475 10.6151
R2076 B.n475 B.n132 10.6151
R2077 B.n471 B.n132 10.6151
R2078 B.n220 B.n1 10.6151
R2079 B.n223 B.n220 10.6151
R2080 B.n224 B.n223 10.6151
R2081 B.n225 B.n224 10.6151
R2082 B.n225 B.n218 10.6151
R2083 B.n229 B.n218 10.6151
R2084 B.n230 B.n229 10.6151
R2085 B.n231 B.n230 10.6151
R2086 B.n231 B.n216 10.6151
R2087 B.n235 B.n216 10.6151
R2088 B.n236 B.n235 10.6151
R2089 B.n237 B.n236 10.6151
R2090 B.n237 B.n214 10.6151
R2091 B.n241 B.n214 10.6151
R2092 B.n242 B.n241 10.6151
R2093 B.n243 B.n242 10.6151
R2094 B.n243 B.n212 10.6151
R2095 B.n247 B.n212 10.6151
R2096 B.n248 B.n247 10.6151
R2097 B.n249 B.n248 10.6151
R2098 B.n249 B.n210 10.6151
R2099 B.n253 B.n210 10.6151
R2100 B.n254 B.n253 10.6151
R2101 B.n255 B.n254 10.6151
R2102 B.n255 B.n208 10.6151
R2103 B.n259 B.n208 10.6151
R2104 B.n260 B.n259 10.6151
R2105 B.n261 B.n260 10.6151
R2106 B.n261 B.n206 10.6151
R2107 B.n265 B.n206 10.6151
R2108 B.n266 B.n265 10.6151
R2109 B.n267 B.n266 10.6151
R2110 B.n267 B.n204 10.6151
R2111 B.n271 B.n204 10.6151
R2112 B.n272 B.n271 10.6151
R2113 B.n273 B.n272 10.6151
R2114 B.n273 B.n202 10.6151
R2115 B.n277 B.n202 10.6151
R2116 B.n278 B.n277 10.6151
R2117 B.n279 B.n278 10.6151
R2118 B.n279 B.n200 10.6151
R2119 B.n284 B.n283 10.6151
R2120 B.n285 B.n284 10.6151
R2121 B.n285 B.n198 10.6151
R2122 B.n289 B.n198 10.6151
R2123 B.n290 B.n289 10.6151
R2124 B.n291 B.n290 10.6151
R2125 B.n291 B.n196 10.6151
R2126 B.n295 B.n196 10.6151
R2127 B.n296 B.n295 10.6151
R2128 B.n297 B.n296 10.6151
R2129 B.n297 B.n194 10.6151
R2130 B.n301 B.n194 10.6151
R2131 B.n302 B.n301 10.6151
R2132 B.n303 B.n302 10.6151
R2133 B.n303 B.n192 10.6151
R2134 B.n307 B.n192 10.6151
R2135 B.n308 B.n307 10.6151
R2136 B.n309 B.n308 10.6151
R2137 B.n309 B.n190 10.6151
R2138 B.n313 B.n190 10.6151
R2139 B.n314 B.n313 10.6151
R2140 B.n315 B.n314 10.6151
R2141 B.n315 B.n188 10.6151
R2142 B.n319 B.n188 10.6151
R2143 B.n320 B.n319 10.6151
R2144 B.n321 B.n320 10.6151
R2145 B.n321 B.n186 10.6151
R2146 B.n325 B.n186 10.6151
R2147 B.n326 B.n325 10.6151
R2148 B.n327 B.n326 10.6151
R2149 B.n327 B.n184 10.6151
R2150 B.n331 B.n184 10.6151
R2151 B.n332 B.n331 10.6151
R2152 B.n333 B.n332 10.6151
R2153 B.n333 B.n182 10.6151
R2154 B.n337 B.n182 10.6151
R2155 B.n338 B.n337 10.6151
R2156 B.n339 B.n338 10.6151
R2157 B.n339 B.n180 10.6151
R2158 B.n343 B.n180 10.6151
R2159 B.n344 B.n343 10.6151
R2160 B.n345 B.n344 10.6151
R2161 B.n345 B.n178 10.6151
R2162 B.n349 B.n178 10.6151
R2163 B.n350 B.n349 10.6151
R2164 B.n351 B.n350 10.6151
R2165 B.n351 B.n176 10.6151
R2166 B.n355 B.n176 10.6151
R2167 B.n356 B.n355 10.6151
R2168 B.n357 B.n356 10.6151
R2169 B.n357 B.n174 10.6151
R2170 B.n361 B.n174 10.6151
R2171 B.n362 B.n361 10.6151
R2172 B.n363 B.n362 10.6151
R2173 B.n363 B.n172 10.6151
R2174 B.n367 B.n172 10.6151
R2175 B.n368 B.n367 10.6151
R2176 B.n370 B.n168 10.6151
R2177 B.n374 B.n168 10.6151
R2178 B.n375 B.n374 10.6151
R2179 B.n376 B.n375 10.6151
R2180 B.n376 B.n166 10.6151
R2181 B.n380 B.n166 10.6151
R2182 B.n381 B.n380 10.6151
R2183 B.n382 B.n381 10.6151
R2184 B.n386 B.n385 10.6151
R2185 B.n387 B.n386 10.6151
R2186 B.n387 B.n160 10.6151
R2187 B.n391 B.n160 10.6151
R2188 B.n392 B.n391 10.6151
R2189 B.n393 B.n392 10.6151
R2190 B.n393 B.n158 10.6151
R2191 B.n397 B.n158 10.6151
R2192 B.n398 B.n397 10.6151
R2193 B.n399 B.n398 10.6151
R2194 B.n399 B.n156 10.6151
R2195 B.n403 B.n156 10.6151
R2196 B.n404 B.n403 10.6151
R2197 B.n405 B.n404 10.6151
R2198 B.n405 B.n154 10.6151
R2199 B.n409 B.n154 10.6151
R2200 B.n410 B.n409 10.6151
R2201 B.n411 B.n410 10.6151
R2202 B.n411 B.n152 10.6151
R2203 B.n415 B.n152 10.6151
R2204 B.n416 B.n415 10.6151
R2205 B.n417 B.n416 10.6151
R2206 B.n417 B.n150 10.6151
R2207 B.n421 B.n150 10.6151
R2208 B.n422 B.n421 10.6151
R2209 B.n423 B.n422 10.6151
R2210 B.n423 B.n148 10.6151
R2211 B.n427 B.n148 10.6151
R2212 B.n428 B.n427 10.6151
R2213 B.n429 B.n428 10.6151
R2214 B.n429 B.n146 10.6151
R2215 B.n433 B.n146 10.6151
R2216 B.n434 B.n433 10.6151
R2217 B.n435 B.n434 10.6151
R2218 B.n435 B.n144 10.6151
R2219 B.n439 B.n144 10.6151
R2220 B.n440 B.n439 10.6151
R2221 B.n441 B.n440 10.6151
R2222 B.n441 B.n142 10.6151
R2223 B.n445 B.n142 10.6151
R2224 B.n446 B.n445 10.6151
R2225 B.n447 B.n446 10.6151
R2226 B.n447 B.n140 10.6151
R2227 B.n451 B.n140 10.6151
R2228 B.n452 B.n451 10.6151
R2229 B.n453 B.n452 10.6151
R2230 B.n453 B.n138 10.6151
R2231 B.n457 B.n138 10.6151
R2232 B.n458 B.n457 10.6151
R2233 B.n459 B.n458 10.6151
R2234 B.n459 B.n136 10.6151
R2235 B.n463 B.n136 10.6151
R2236 B.n464 B.n463 10.6151
R2237 B.n465 B.n464 10.6151
R2238 B.n465 B.n134 10.6151
R2239 B.n469 B.n134 10.6151
R2240 B.n470 B.n469 10.6151
R2241 B.n853 B.n0 8.11757
R2242 B.n853 B.n1 8.11757
R2243 B.n700 B.n54 6.5566
R2244 B.n688 B.n687 6.5566
R2245 B.n370 B.n369 6.5566
R2246 B.n382 B.n164 6.5566
R2247 B.n703 B.n54 4.05904
R2248 B.n687 B.n686 4.05904
R2249 B.n369 B.n368 4.05904
R2250 B.n385 B.n164 4.05904
R2251 VP.n11 VP.t2 194.712
R2252 VP.n13 VP.n12 161.3
R2253 VP.n14 VP.n9 161.3
R2254 VP.n16 VP.n15 161.3
R2255 VP.n17 VP.n8 161.3
R2256 VP.n19 VP.n18 161.3
R2257 VP.n20 VP.n7 161.3
R2258 VP.n42 VP.n0 161.3
R2259 VP.n41 VP.n40 161.3
R2260 VP.n39 VP.n1 161.3
R2261 VP.n38 VP.n37 161.3
R2262 VP.n36 VP.n2 161.3
R2263 VP.n35 VP.n34 161.3
R2264 VP.n33 VP.n32 161.3
R2265 VP.n31 VP.n4 161.3
R2266 VP.n30 VP.n29 161.3
R2267 VP.n28 VP.n5 161.3
R2268 VP.n27 VP.n26 161.3
R2269 VP.n25 VP.n6 161.3
R2270 VP.n24 VP.t5 161.221
R2271 VP.n3 VP.t1 161.221
R2272 VP.n43 VP.t0 161.221
R2273 VP.n21 VP.t4 161.221
R2274 VP.n10 VP.t3 161.221
R2275 VP.n24 VP.n23 101.564
R2276 VP.n44 VP.n43 101.564
R2277 VP.n22 VP.n21 101.564
R2278 VP.n11 VP.n10 60.3423
R2279 VP.n30 VP.n5 56.5617
R2280 VP.n37 VP.n1 56.5617
R2281 VP.n15 VP.n8 56.5617
R2282 VP.n23 VP.n22 52.8633
R2283 VP.n26 VP.n25 24.5923
R2284 VP.n26 VP.n5 24.5923
R2285 VP.n31 VP.n30 24.5923
R2286 VP.n32 VP.n31 24.5923
R2287 VP.n36 VP.n35 24.5923
R2288 VP.n37 VP.n36 24.5923
R2289 VP.n41 VP.n1 24.5923
R2290 VP.n42 VP.n41 24.5923
R2291 VP.n19 VP.n8 24.5923
R2292 VP.n20 VP.n19 24.5923
R2293 VP.n14 VP.n13 24.5923
R2294 VP.n15 VP.n14 24.5923
R2295 VP.n32 VP.n3 12.2964
R2296 VP.n35 VP.n3 12.2964
R2297 VP.n13 VP.n10 12.2964
R2298 VP.n25 VP.n24 9.3454
R2299 VP.n43 VP.n42 9.3454
R2300 VP.n21 VP.n20 9.3454
R2301 VP.n12 VP.n11 6.87456
R2302 VP.n22 VP.n7 0.278335
R2303 VP.n23 VP.n6 0.278335
R2304 VP.n44 VP.n0 0.278335
R2305 VP.n12 VP.n9 0.189894
R2306 VP.n16 VP.n9 0.189894
R2307 VP.n17 VP.n16 0.189894
R2308 VP.n18 VP.n17 0.189894
R2309 VP.n18 VP.n7 0.189894
R2310 VP.n27 VP.n6 0.189894
R2311 VP.n28 VP.n27 0.189894
R2312 VP.n29 VP.n28 0.189894
R2313 VP.n29 VP.n4 0.189894
R2314 VP.n33 VP.n4 0.189894
R2315 VP.n34 VP.n33 0.189894
R2316 VP.n34 VP.n2 0.189894
R2317 VP.n38 VP.n2 0.189894
R2318 VP.n39 VP.n38 0.189894
R2319 VP.n40 VP.n39 0.189894
R2320 VP.n40 VP.n0 0.189894
R2321 VP VP.n44 0.153485
R2322 VDD1.n92 VDD1.n0 756.745
R2323 VDD1.n189 VDD1.n97 756.745
R2324 VDD1.n93 VDD1.n92 585
R2325 VDD1.n91 VDD1.n90 585
R2326 VDD1.n4 VDD1.n3 585
R2327 VDD1.n85 VDD1.n84 585
R2328 VDD1.n83 VDD1.n82 585
R2329 VDD1.n8 VDD1.n7 585
R2330 VDD1.n12 VDD1.n10 585
R2331 VDD1.n77 VDD1.n76 585
R2332 VDD1.n75 VDD1.n74 585
R2333 VDD1.n14 VDD1.n13 585
R2334 VDD1.n69 VDD1.n68 585
R2335 VDD1.n67 VDD1.n66 585
R2336 VDD1.n18 VDD1.n17 585
R2337 VDD1.n61 VDD1.n60 585
R2338 VDD1.n59 VDD1.n58 585
R2339 VDD1.n22 VDD1.n21 585
R2340 VDD1.n53 VDD1.n52 585
R2341 VDD1.n51 VDD1.n50 585
R2342 VDD1.n26 VDD1.n25 585
R2343 VDD1.n45 VDD1.n44 585
R2344 VDD1.n43 VDD1.n42 585
R2345 VDD1.n30 VDD1.n29 585
R2346 VDD1.n37 VDD1.n36 585
R2347 VDD1.n35 VDD1.n34 585
R2348 VDD1.n130 VDD1.n129 585
R2349 VDD1.n132 VDD1.n131 585
R2350 VDD1.n125 VDD1.n124 585
R2351 VDD1.n138 VDD1.n137 585
R2352 VDD1.n140 VDD1.n139 585
R2353 VDD1.n121 VDD1.n120 585
R2354 VDD1.n146 VDD1.n145 585
R2355 VDD1.n148 VDD1.n147 585
R2356 VDD1.n117 VDD1.n116 585
R2357 VDD1.n154 VDD1.n153 585
R2358 VDD1.n156 VDD1.n155 585
R2359 VDD1.n113 VDD1.n112 585
R2360 VDD1.n162 VDD1.n161 585
R2361 VDD1.n164 VDD1.n163 585
R2362 VDD1.n109 VDD1.n108 585
R2363 VDD1.n171 VDD1.n170 585
R2364 VDD1.n172 VDD1.n107 585
R2365 VDD1.n174 VDD1.n173 585
R2366 VDD1.n105 VDD1.n104 585
R2367 VDD1.n180 VDD1.n179 585
R2368 VDD1.n182 VDD1.n181 585
R2369 VDD1.n101 VDD1.n100 585
R2370 VDD1.n188 VDD1.n187 585
R2371 VDD1.n190 VDD1.n189 585
R2372 VDD1.n33 VDD1.t3 327.466
R2373 VDD1.n128 VDD1.t0 327.466
R2374 VDD1.n92 VDD1.n91 171.744
R2375 VDD1.n91 VDD1.n3 171.744
R2376 VDD1.n84 VDD1.n3 171.744
R2377 VDD1.n84 VDD1.n83 171.744
R2378 VDD1.n83 VDD1.n7 171.744
R2379 VDD1.n12 VDD1.n7 171.744
R2380 VDD1.n76 VDD1.n12 171.744
R2381 VDD1.n76 VDD1.n75 171.744
R2382 VDD1.n75 VDD1.n13 171.744
R2383 VDD1.n68 VDD1.n13 171.744
R2384 VDD1.n68 VDD1.n67 171.744
R2385 VDD1.n67 VDD1.n17 171.744
R2386 VDD1.n60 VDD1.n17 171.744
R2387 VDD1.n60 VDD1.n59 171.744
R2388 VDD1.n59 VDD1.n21 171.744
R2389 VDD1.n52 VDD1.n21 171.744
R2390 VDD1.n52 VDD1.n51 171.744
R2391 VDD1.n51 VDD1.n25 171.744
R2392 VDD1.n44 VDD1.n25 171.744
R2393 VDD1.n44 VDD1.n43 171.744
R2394 VDD1.n43 VDD1.n29 171.744
R2395 VDD1.n36 VDD1.n29 171.744
R2396 VDD1.n36 VDD1.n35 171.744
R2397 VDD1.n131 VDD1.n130 171.744
R2398 VDD1.n131 VDD1.n124 171.744
R2399 VDD1.n138 VDD1.n124 171.744
R2400 VDD1.n139 VDD1.n138 171.744
R2401 VDD1.n139 VDD1.n120 171.744
R2402 VDD1.n146 VDD1.n120 171.744
R2403 VDD1.n147 VDD1.n146 171.744
R2404 VDD1.n147 VDD1.n116 171.744
R2405 VDD1.n154 VDD1.n116 171.744
R2406 VDD1.n155 VDD1.n154 171.744
R2407 VDD1.n155 VDD1.n112 171.744
R2408 VDD1.n162 VDD1.n112 171.744
R2409 VDD1.n163 VDD1.n162 171.744
R2410 VDD1.n163 VDD1.n108 171.744
R2411 VDD1.n171 VDD1.n108 171.744
R2412 VDD1.n172 VDD1.n171 171.744
R2413 VDD1.n173 VDD1.n172 171.744
R2414 VDD1.n173 VDD1.n104 171.744
R2415 VDD1.n180 VDD1.n104 171.744
R2416 VDD1.n181 VDD1.n180 171.744
R2417 VDD1.n181 VDD1.n100 171.744
R2418 VDD1.n188 VDD1.n100 171.744
R2419 VDD1.n189 VDD1.n188 171.744
R2420 VDD1.n35 VDD1.t3 85.8723
R2421 VDD1.n130 VDD1.t0 85.8723
R2422 VDD1.n195 VDD1.n194 68.4367
R2423 VDD1.n197 VDD1.n196 67.8584
R2424 VDD1 VDD1.n96 49.6595
R2425 VDD1.n195 VDD1.n193 49.546
R2426 VDD1.n197 VDD1.n195 48.8543
R2427 VDD1.n34 VDD1.n33 16.3895
R2428 VDD1.n129 VDD1.n128 16.3895
R2429 VDD1.n10 VDD1.n8 13.1884
R2430 VDD1.n174 VDD1.n105 13.1884
R2431 VDD1.n82 VDD1.n81 12.8005
R2432 VDD1.n78 VDD1.n77 12.8005
R2433 VDD1.n37 VDD1.n32 12.8005
R2434 VDD1.n132 VDD1.n127 12.8005
R2435 VDD1.n175 VDD1.n107 12.8005
R2436 VDD1.n179 VDD1.n178 12.8005
R2437 VDD1.n85 VDD1.n6 12.0247
R2438 VDD1.n74 VDD1.n11 12.0247
R2439 VDD1.n38 VDD1.n30 12.0247
R2440 VDD1.n133 VDD1.n125 12.0247
R2441 VDD1.n170 VDD1.n169 12.0247
R2442 VDD1.n182 VDD1.n103 12.0247
R2443 VDD1.n86 VDD1.n4 11.249
R2444 VDD1.n73 VDD1.n14 11.249
R2445 VDD1.n42 VDD1.n41 11.249
R2446 VDD1.n137 VDD1.n136 11.249
R2447 VDD1.n168 VDD1.n109 11.249
R2448 VDD1.n183 VDD1.n101 11.249
R2449 VDD1.n90 VDD1.n89 10.4732
R2450 VDD1.n70 VDD1.n69 10.4732
R2451 VDD1.n45 VDD1.n28 10.4732
R2452 VDD1.n140 VDD1.n123 10.4732
R2453 VDD1.n165 VDD1.n164 10.4732
R2454 VDD1.n187 VDD1.n186 10.4732
R2455 VDD1.n93 VDD1.n2 9.69747
R2456 VDD1.n66 VDD1.n16 9.69747
R2457 VDD1.n46 VDD1.n26 9.69747
R2458 VDD1.n141 VDD1.n121 9.69747
R2459 VDD1.n161 VDD1.n111 9.69747
R2460 VDD1.n190 VDD1.n99 9.69747
R2461 VDD1.n96 VDD1.n95 9.45567
R2462 VDD1.n193 VDD1.n192 9.45567
R2463 VDD1.n20 VDD1.n19 9.3005
R2464 VDD1.n63 VDD1.n62 9.3005
R2465 VDD1.n65 VDD1.n64 9.3005
R2466 VDD1.n16 VDD1.n15 9.3005
R2467 VDD1.n71 VDD1.n70 9.3005
R2468 VDD1.n73 VDD1.n72 9.3005
R2469 VDD1.n11 VDD1.n9 9.3005
R2470 VDD1.n79 VDD1.n78 9.3005
R2471 VDD1.n95 VDD1.n94 9.3005
R2472 VDD1.n2 VDD1.n1 9.3005
R2473 VDD1.n89 VDD1.n88 9.3005
R2474 VDD1.n87 VDD1.n86 9.3005
R2475 VDD1.n6 VDD1.n5 9.3005
R2476 VDD1.n81 VDD1.n80 9.3005
R2477 VDD1.n57 VDD1.n56 9.3005
R2478 VDD1.n55 VDD1.n54 9.3005
R2479 VDD1.n24 VDD1.n23 9.3005
R2480 VDD1.n49 VDD1.n48 9.3005
R2481 VDD1.n47 VDD1.n46 9.3005
R2482 VDD1.n28 VDD1.n27 9.3005
R2483 VDD1.n41 VDD1.n40 9.3005
R2484 VDD1.n39 VDD1.n38 9.3005
R2485 VDD1.n32 VDD1.n31 9.3005
R2486 VDD1.n192 VDD1.n191 9.3005
R2487 VDD1.n99 VDD1.n98 9.3005
R2488 VDD1.n186 VDD1.n185 9.3005
R2489 VDD1.n184 VDD1.n183 9.3005
R2490 VDD1.n103 VDD1.n102 9.3005
R2491 VDD1.n178 VDD1.n177 9.3005
R2492 VDD1.n150 VDD1.n149 9.3005
R2493 VDD1.n119 VDD1.n118 9.3005
R2494 VDD1.n144 VDD1.n143 9.3005
R2495 VDD1.n142 VDD1.n141 9.3005
R2496 VDD1.n123 VDD1.n122 9.3005
R2497 VDD1.n136 VDD1.n135 9.3005
R2498 VDD1.n134 VDD1.n133 9.3005
R2499 VDD1.n127 VDD1.n126 9.3005
R2500 VDD1.n152 VDD1.n151 9.3005
R2501 VDD1.n115 VDD1.n114 9.3005
R2502 VDD1.n158 VDD1.n157 9.3005
R2503 VDD1.n160 VDD1.n159 9.3005
R2504 VDD1.n111 VDD1.n110 9.3005
R2505 VDD1.n166 VDD1.n165 9.3005
R2506 VDD1.n168 VDD1.n167 9.3005
R2507 VDD1.n169 VDD1.n106 9.3005
R2508 VDD1.n176 VDD1.n175 9.3005
R2509 VDD1.n94 VDD1.n0 8.92171
R2510 VDD1.n65 VDD1.n18 8.92171
R2511 VDD1.n50 VDD1.n49 8.92171
R2512 VDD1.n145 VDD1.n144 8.92171
R2513 VDD1.n160 VDD1.n113 8.92171
R2514 VDD1.n191 VDD1.n97 8.92171
R2515 VDD1.n62 VDD1.n61 8.14595
R2516 VDD1.n53 VDD1.n24 8.14595
R2517 VDD1.n148 VDD1.n119 8.14595
R2518 VDD1.n157 VDD1.n156 8.14595
R2519 VDD1.n58 VDD1.n20 7.3702
R2520 VDD1.n54 VDD1.n22 7.3702
R2521 VDD1.n149 VDD1.n117 7.3702
R2522 VDD1.n153 VDD1.n115 7.3702
R2523 VDD1.n58 VDD1.n57 6.59444
R2524 VDD1.n57 VDD1.n22 6.59444
R2525 VDD1.n152 VDD1.n117 6.59444
R2526 VDD1.n153 VDD1.n152 6.59444
R2527 VDD1.n61 VDD1.n20 5.81868
R2528 VDD1.n54 VDD1.n53 5.81868
R2529 VDD1.n149 VDD1.n148 5.81868
R2530 VDD1.n156 VDD1.n115 5.81868
R2531 VDD1.n96 VDD1.n0 5.04292
R2532 VDD1.n62 VDD1.n18 5.04292
R2533 VDD1.n50 VDD1.n24 5.04292
R2534 VDD1.n145 VDD1.n119 5.04292
R2535 VDD1.n157 VDD1.n113 5.04292
R2536 VDD1.n193 VDD1.n97 5.04292
R2537 VDD1.n94 VDD1.n93 4.26717
R2538 VDD1.n66 VDD1.n65 4.26717
R2539 VDD1.n49 VDD1.n26 4.26717
R2540 VDD1.n144 VDD1.n121 4.26717
R2541 VDD1.n161 VDD1.n160 4.26717
R2542 VDD1.n191 VDD1.n190 4.26717
R2543 VDD1.n33 VDD1.n31 3.70982
R2544 VDD1.n128 VDD1.n126 3.70982
R2545 VDD1.n90 VDD1.n2 3.49141
R2546 VDD1.n69 VDD1.n16 3.49141
R2547 VDD1.n46 VDD1.n45 3.49141
R2548 VDD1.n141 VDD1.n140 3.49141
R2549 VDD1.n164 VDD1.n111 3.49141
R2550 VDD1.n187 VDD1.n99 3.49141
R2551 VDD1.n89 VDD1.n4 2.71565
R2552 VDD1.n70 VDD1.n14 2.71565
R2553 VDD1.n42 VDD1.n28 2.71565
R2554 VDD1.n137 VDD1.n123 2.71565
R2555 VDD1.n165 VDD1.n109 2.71565
R2556 VDD1.n186 VDD1.n101 2.71565
R2557 VDD1.n86 VDD1.n85 1.93989
R2558 VDD1.n74 VDD1.n73 1.93989
R2559 VDD1.n41 VDD1.n30 1.93989
R2560 VDD1.n136 VDD1.n125 1.93989
R2561 VDD1.n170 VDD1.n168 1.93989
R2562 VDD1.n183 VDD1.n182 1.93989
R2563 VDD1.n196 VDD1.t2 1.86218
R2564 VDD1.n196 VDD1.t1 1.86218
R2565 VDD1.n194 VDD1.t4 1.86218
R2566 VDD1.n194 VDD1.t5 1.86218
R2567 VDD1.n82 VDD1.n6 1.16414
R2568 VDD1.n77 VDD1.n11 1.16414
R2569 VDD1.n38 VDD1.n37 1.16414
R2570 VDD1.n133 VDD1.n132 1.16414
R2571 VDD1.n169 VDD1.n107 1.16414
R2572 VDD1.n179 VDD1.n103 1.16414
R2573 VDD1 VDD1.n197 0.575931
R2574 VDD1.n81 VDD1.n8 0.388379
R2575 VDD1.n78 VDD1.n10 0.388379
R2576 VDD1.n34 VDD1.n32 0.388379
R2577 VDD1.n129 VDD1.n127 0.388379
R2578 VDD1.n175 VDD1.n174 0.388379
R2579 VDD1.n178 VDD1.n105 0.388379
R2580 VDD1.n95 VDD1.n1 0.155672
R2581 VDD1.n88 VDD1.n1 0.155672
R2582 VDD1.n88 VDD1.n87 0.155672
R2583 VDD1.n87 VDD1.n5 0.155672
R2584 VDD1.n80 VDD1.n5 0.155672
R2585 VDD1.n80 VDD1.n79 0.155672
R2586 VDD1.n79 VDD1.n9 0.155672
R2587 VDD1.n72 VDD1.n9 0.155672
R2588 VDD1.n72 VDD1.n71 0.155672
R2589 VDD1.n71 VDD1.n15 0.155672
R2590 VDD1.n64 VDD1.n15 0.155672
R2591 VDD1.n64 VDD1.n63 0.155672
R2592 VDD1.n63 VDD1.n19 0.155672
R2593 VDD1.n56 VDD1.n19 0.155672
R2594 VDD1.n56 VDD1.n55 0.155672
R2595 VDD1.n55 VDD1.n23 0.155672
R2596 VDD1.n48 VDD1.n23 0.155672
R2597 VDD1.n48 VDD1.n47 0.155672
R2598 VDD1.n47 VDD1.n27 0.155672
R2599 VDD1.n40 VDD1.n27 0.155672
R2600 VDD1.n40 VDD1.n39 0.155672
R2601 VDD1.n39 VDD1.n31 0.155672
R2602 VDD1.n134 VDD1.n126 0.155672
R2603 VDD1.n135 VDD1.n134 0.155672
R2604 VDD1.n135 VDD1.n122 0.155672
R2605 VDD1.n142 VDD1.n122 0.155672
R2606 VDD1.n143 VDD1.n142 0.155672
R2607 VDD1.n143 VDD1.n118 0.155672
R2608 VDD1.n150 VDD1.n118 0.155672
R2609 VDD1.n151 VDD1.n150 0.155672
R2610 VDD1.n151 VDD1.n114 0.155672
R2611 VDD1.n158 VDD1.n114 0.155672
R2612 VDD1.n159 VDD1.n158 0.155672
R2613 VDD1.n159 VDD1.n110 0.155672
R2614 VDD1.n166 VDD1.n110 0.155672
R2615 VDD1.n167 VDD1.n166 0.155672
R2616 VDD1.n167 VDD1.n106 0.155672
R2617 VDD1.n176 VDD1.n106 0.155672
R2618 VDD1.n177 VDD1.n176 0.155672
R2619 VDD1.n177 VDD1.n102 0.155672
R2620 VDD1.n184 VDD1.n102 0.155672
R2621 VDD1.n185 VDD1.n184 0.155672
R2622 VDD1.n185 VDD1.n98 0.155672
R2623 VDD1.n192 VDD1.n98 0.155672
C0 w_n3322_n4460# B 11.220799f
C1 VDD2 VDD1 1.41209f
C2 VP VDD2 0.460018f
C3 VN VDD1 0.151167f
C4 VP VN 7.94168f
C5 VTAIL VDD1 9.708529f
C6 VP VTAIL 9.54427f
C7 VDD2 w_n3322_n4460# 2.7597f
C8 VN w_n3322_n4460# 6.38461f
C9 w_n3322_n4460# VTAIL 3.73945f
C10 VP VDD1 9.91963f
C11 w_n3322_n4460# VDD1 2.67434f
C12 VP w_n3322_n4460# 6.81412f
C13 VDD2 B 2.60125f
C14 VN B 1.23715f
C15 B VTAIL 4.92251f
C16 B VDD1 2.52692f
C17 VN VDD2 9.61492f
C18 VP B 1.95432f
C19 VDD2 VTAIL 9.75817f
C20 VN VTAIL 9.529901f
C21 VDD2 VSUBS 2.07863f
C22 VDD1 VSUBS 1.983235f
C23 VTAIL VSUBS 1.385587f
C24 VN VSUBS 6.06306f
C25 VP VSUBS 3.140201f
C26 B VSUBS 5.109948f
C27 w_n3322_n4460# VSUBS 0.181262p
C28 VDD1.n0 VSUBS 0.028444f
C29 VDD1.n1 VSUBS 0.027032f
C30 VDD1.n2 VSUBS 0.014526f
C31 VDD1.n3 VSUBS 0.034334f
C32 VDD1.n4 VSUBS 0.015381f
C33 VDD1.n5 VSUBS 0.027032f
C34 VDD1.n6 VSUBS 0.014526f
C35 VDD1.n7 VSUBS 0.034334f
C36 VDD1.n8 VSUBS 0.014953f
C37 VDD1.n9 VSUBS 0.027032f
C38 VDD1.n10 VSUBS 0.014953f
C39 VDD1.n11 VSUBS 0.014526f
C40 VDD1.n12 VSUBS 0.034334f
C41 VDD1.n13 VSUBS 0.034334f
C42 VDD1.n14 VSUBS 0.015381f
C43 VDD1.n15 VSUBS 0.027032f
C44 VDD1.n16 VSUBS 0.014526f
C45 VDD1.n17 VSUBS 0.034334f
C46 VDD1.n18 VSUBS 0.015381f
C47 VDD1.n19 VSUBS 0.027032f
C48 VDD1.n20 VSUBS 0.014526f
C49 VDD1.n21 VSUBS 0.034334f
C50 VDD1.n22 VSUBS 0.015381f
C51 VDD1.n23 VSUBS 0.027032f
C52 VDD1.n24 VSUBS 0.014526f
C53 VDD1.n25 VSUBS 0.034334f
C54 VDD1.n26 VSUBS 0.015381f
C55 VDD1.n27 VSUBS 0.027032f
C56 VDD1.n28 VSUBS 0.014526f
C57 VDD1.n29 VSUBS 0.034334f
C58 VDD1.n30 VSUBS 0.015381f
C59 VDD1.n31 VSUBS 2.02796f
C60 VDD1.n32 VSUBS 0.014526f
C61 VDD1.t3 VSUBS 0.073668f
C62 VDD1.n33 VSUBS 0.210169f
C63 VDD1.n34 VSUBS 0.021842f
C64 VDD1.n35 VSUBS 0.025751f
C65 VDD1.n36 VSUBS 0.034334f
C66 VDD1.n37 VSUBS 0.015381f
C67 VDD1.n38 VSUBS 0.014526f
C68 VDD1.n39 VSUBS 0.027032f
C69 VDD1.n40 VSUBS 0.027032f
C70 VDD1.n41 VSUBS 0.014526f
C71 VDD1.n42 VSUBS 0.015381f
C72 VDD1.n43 VSUBS 0.034334f
C73 VDD1.n44 VSUBS 0.034334f
C74 VDD1.n45 VSUBS 0.015381f
C75 VDD1.n46 VSUBS 0.014526f
C76 VDD1.n47 VSUBS 0.027032f
C77 VDD1.n48 VSUBS 0.027032f
C78 VDD1.n49 VSUBS 0.014526f
C79 VDD1.n50 VSUBS 0.015381f
C80 VDD1.n51 VSUBS 0.034334f
C81 VDD1.n52 VSUBS 0.034334f
C82 VDD1.n53 VSUBS 0.015381f
C83 VDD1.n54 VSUBS 0.014526f
C84 VDD1.n55 VSUBS 0.027032f
C85 VDD1.n56 VSUBS 0.027032f
C86 VDD1.n57 VSUBS 0.014526f
C87 VDD1.n58 VSUBS 0.015381f
C88 VDD1.n59 VSUBS 0.034334f
C89 VDD1.n60 VSUBS 0.034334f
C90 VDD1.n61 VSUBS 0.015381f
C91 VDD1.n62 VSUBS 0.014526f
C92 VDD1.n63 VSUBS 0.027032f
C93 VDD1.n64 VSUBS 0.027032f
C94 VDD1.n65 VSUBS 0.014526f
C95 VDD1.n66 VSUBS 0.015381f
C96 VDD1.n67 VSUBS 0.034334f
C97 VDD1.n68 VSUBS 0.034334f
C98 VDD1.n69 VSUBS 0.015381f
C99 VDD1.n70 VSUBS 0.014526f
C100 VDD1.n71 VSUBS 0.027032f
C101 VDD1.n72 VSUBS 0.027032f
C102 VDD1.n73 VSUBS 0.014526f
C103 VDD1.n74 VSUBS 0.015381f
C104 VDD1.n75 VSUBS 0.034334f
C105 VDD1.n76 VSUBS 0.034334f
C106 VDD1.n77 VSUBS 0.015381f
C107 VDD1.n78 VSUBS 0.014526f
C108 VDD1.n79 VSUBS 0.027032f
C109 VDD1.n80 VSUBS 0.027032f
C110 VDD1.n81 VSUBS 0.014526f
C111 VDD1.n82 VSUBS 0.015381f
C112 VDD1.n83 VSUBS 0.034334f
C113 VDD1.n84 VSUBS 0.034334f
C114 VDD1.n85 VSUBS 0.015381f
C115 VDD1.n86 VSUBS 0.014526f
C116 VDD1.n87 VSUBS 0.027032f
C117 VDD1.n88 VSUBS 0.027032f
C118 VDD1.n89 VSUBS 0.014526f
C119 VDD1.n90 VSUBS 0.015381f
C120 VDD1.n91 VSUBS 0.034334f
C121 VDD1.n92 VSUBS 0.078831f
C122 VDD1.n93 VSUBS 0.015381f
C123 VDD1.n94 VSUBS 0.014526f
C124 VDD1.n95 VSUBS 0.060268f
C125 VDD1.n96 VSUBS 0.066803f
C126 VDD1.n97 VSUBS 0.028444f
C127 VDD1.n98 VSUBS 0.027032f
C128 VDD1.n99 VSUBS 0.014526f
C129 VDD1.n100 VSUBS 0.034334f
C130 VDD1.n101 VSUBS 0.015381f
C131 VDD1.n102 VSUBS 0.027032f
C132 VDD1.n103 VSUBS 0.014526f
C133 VDD1.n104 VSUBS 0.034334f
C134 VDD1.n105 VSUBS 0.014953f
C135 VDD1.n106 VSUBS 0.027032f
C136 VDD1.n107 VSUBS 0.015381f
C137 VDD1.n108 VSUBS 0.034334f
C138 VDD1.n109 VSUBS 0.015381f
C139 VDD1.n110 VSUBS 0.027032f
C140 VDD1.n111 VSUBS 0.014526f
C141 VDD1.n112 VSUBS 0.034334f
C142 VDD1.n113 VSUBS 0.015381f
C143 VDD1.n114 VSUBS 0.027032f
C144 VDD1.n115 VSUBS 0.014526f
C145 VDD1.n116 VSUBS 0.034334f
C146 VDD1.n117 VSUBS 0.015381f
C147 VDD1.n118 VSUBS 0.027032f
C148 VDD1.n119 VSUBS 0.014526f
C149 VDD1.n120 VSUBS 0.034334f
C150 VDD1.n121 VSUBS 0.015381f
C151 VDD1.n122 VSUBS 0.027032f
C152 VDD1.n123 VSUBS 0.014526f
C153 VDD1.n124 VSUBS 0.034334f
C154 VDD1.n125 VSUBS 0.015381f
C155 VDD1.n126 VSUBS 2.02796f
C156 VDD1.n127 VSUBS 0.014526f
C157 VDD1.t0 VSUBS 0.073668f
C158 VDD1.n128 VSUBS 0.210169f
C159 VDD1.n129 VSUBS 0.021842f
C160 VDD1.n130 VSUBS 0.025751f
C161 VDD1.n131 VSUBS 0.034334f
C162 VDD1.n132 VSUBS 0.015381f
C163 VDD1.n133 VSUBS 0.014526f
C164 VDD1.n134 VSUBS 0.027032f
C165 VDD1.n135 VSUBS 0.027032f
C166 VDD1.n136 VSUBS 0.014526f
C167 VDD1.n137 VSUBS 0.015381f
C168 VDD1.n138 VSUBS 0.034334f
C169 VDD1.n139 VSUBS 0.034334f
C170 VDD1.n140 VSUBS 0.015381f
C171 VDD1.n141 VSUBS 0.014526f
C172 VDD1.n142 VSUBS 0.027032f
C173 VDD1.n143 VSUBS 0.027032f
C174 VDD1.n144 VSUBS 0.014526f
C175 VDD1.n145 VSUBS 0.015381f
C176 VDD1.n146 VSUBS 0.034334f
C177 VDD1.n147 VSUBS 0.034334f
C178 VDD1.n148 VSUBS 0.015381f
C179 VDD1.n149 VSUBS 0.014526f
C180 VDD1.n150 VSUBS 0.027032f
C181 VDD1.n151 VSUBS 0.027032f
C182 VDD1.n152 VSUBS 0.014526f
C183 VDD1.n153 VSUBS 0.015381f
C184 VDD1.n154 VSUBS 0.034334f
C185 VDD1.n155 VSUBS 0.034334f
C186 VDD1.n156 VSUBS 0.015381f
C187 VDD1.n157 VSUBS 0.014526f
C188 VDD1.n158 VSUBS 0.027032f
C189 VDD1.n159 VSUBS 0.027032f
C190 VDD1.n160 VSUBS 0.014526f
C191 VDD1.n161 VSUBS 0.015381f
C192 VDD1.n162 VSUBS 0.034334f
C193 VDD1.n163 VSUBS 0.034334f
C194 VDD1.n164 VSUBS 0.015381f
C195 VDD1.n165 VSUBS 0.014526f
C196 VDD1.n166 VSUBS 0.027032f
C197 VDD1.n167 VSUBS 0.027032f
C198 VDD1.n168 VSUBS 0.014526f
C199 VDD1.n169 VSUBS 0.014526f
C200 VDD1.n170 VSUBS 0.015381f
C201 VDD1.n171 VSUBS 0.034334f
C202 VDD1.n172 VSUBS 0.034334f
C203 VDD1.n173 VSUBS 0.034334f
C204 VDD1.n174 VSUBS 0.014953f
C205 VDD1.n175 VSUBS 0.014526f
C206 VDD1.n176 VSUBS 0.027032f
C207 VDD1.n177 VSUBS 0.027032f
C208 VDD1.n178 VSUBS 0.014526f
C209 VDD1.n179 VSUBS 0.015381f
C210 VDD1.n180 VSUBS 0.034334f
C211 VDD1.n181 VSUBS 0.034334f
C212 VDD1.n182 VSUBS 0.015381f
C213 VDD1.n183 VSUBS 0.014526f
C214 VDD1.n184 VSUBS 0.027032f
C215 VDD1.n185 VSUBS 0.027032f
C216 VDD1.n186 VSUBS 0.014526f
C217 VDD1.n187 VSUBS 0.015381f
C218 VDD1.n188 VSUBS 0.034334f
C219 VDD1.n189 VSUBS 0.078831f
C220 VDD1.n190 VSUBS 0.015381f
C221 VDD1.n191 VSUBS 0.014526f
C222 VDD1.n192 VSUBS 0.060268f
C223 VDD1.n193 VSUBS 0.065959f
C224 VDD1.t4 VSUBS 0.372976f
C225 VDD1.t5 VSUBS 0.372976f
C226 VDD1.n194 VSUBS 3.08722f
C227 VDD1.n195 VSUBS 3.71862f
C228 VDD1.t2 VSUBS 0.372976f
C229 VDD1.t1 VSUBS 0.372976f
C230 VDD1.n196 VSUBS 3.08029f
C231 VDD1.n197 VSUBS 3.78184f
C232 VP.n0 VSUBS 0.036985f
C233 VP.t0 VSUBS 3.51445f
C234 VP.n1 VSUBS 0.04311f
C235 VP.n2 VSUBS 0.028055f
C236 VP.t1 VSUBS 3.51445f
C237 VP.n3 VSUBS 1.21997f
C238 VP.n4 VSUBS 0.028055f
C239 VP.n5 VSUBS 0.04311f
C240 VP.n6 VSUBS 0.036985f
C241 VP.t5 VSUBS 3.51445f
C242 VP.n7 VSUBS 0.036985f
C243 VP.t4 VSUBS 3.51445f
C244 VP.n8 VSUBS 0.04311f
C245 VP.n9 VSUBS 0.028055f
C246 VP.t3 VSUBS 3.51445f
C247 VP.n10 VSUBS 1.30049f
C248 VP.t2 VSUBS 3.75405f
C249 VP.n11 VSUBS 1.26975f
C250 VP.n12 VSUBS 0.271409f
C251 VP.n13 VSUBS 0.039183f
C252 VP.n14 VSUBS 0.052025f
C253 VP.n15 VSUBS 0.038453f
C254 VP.n16 VSUBS 0.028055f
C255 VP.n17 VSUBS 0.028055f
C256 VP.n18 VSUBS 0.028055f
C257 VP.n19 VSUBS 0.052025f
C258 VP.n20 VSUBS 0.036101f
C259 VP.n21 VSUBS 1.31281f
C260 VP.n22 VSUBS 1.69294f
C261 VP.n23 VSUBS 1.71207f
C262 VP.n24 VSUBS 1.31281f
C263 VP.n25 VSUBS 0.036101f
C264 VP.n26 VSUBS 0.052025f
C265 VP.n27 VSUBS 0.028055f
C266 VP.n28 VSUBS 0.028055f
C267 VP.n29 VSUBS 0.028055f
C268 VP.n30 VSUBS 0.038453f
C269 VP.n31 VSUBS 0.052025f
C270 VP.n32 VSUBS 0.039183f
C271 VP.n33 VSUBS 0.028055f
C272 VP.n34 VSUBS 0.028055f
C273 VP.n35 VSUBS 0.039183f
C274 VP.n36 VSUBS 0.052025f
C275 VP.n37 VSUBS 0.038453f
C276 VP.n38 VSUBS 0.028055f
C277 VP.n39 VSUBS 0.028055f
C278 VP.n40 VSUBS 0.028055f
C279 VP.n41 VSUBS 0.052025f
C280 VP.n42 VSUBS 0.036101f
C281 VP.n43 VSUBS 1.31281f
C282 VP.n44 VSUBS 0.046205f
C283 B.n0 VSUBS 0.006343f
C284 B.n1 VSUBS 0.006343f
C285 B.n2 VSUBS 0.00938f
C286 B.n3 VSUBS 0.007188f
C287 B.n4 VSUBS 0.007188f
C288 B.n5 VSUBS 0.007188f
C289 B.n6 VSUBS 0.007188f
C290 B.n7 VSUBS 0.007188f
C291 B.n8 VSUBS 0.007188f
C292 B.n9 VSUBS 0.007188f
C293 B.n10 VSUBS 0.007188f
C294 B.n11 VSUBS 0.007188f
C295 B.n12 VSUBS 0.007188f
C296 B.n13 VSUBS 0.007188f
C297 B.n14 VSUBS 0.007188f
C298 B.n15 VSUBS 0.007188f
C299 B.n16 VSUBS 0.007188f
C300 B.n17 VSUBS 0.007188f
C301 B.n18 VSUBS 0.007188f
C302 B.n19 VSUBS 0.007188f
C303 B.n20 VSUBS 0.007188f
C304 B.n21 VSUBS 0.007188f
C305 B.n22 VSUBS 0.007188f
C306 B.n23 VSUBS 0.017881f
C307 B.n24 VSUBS 0.007188f
C308 B.n25 VSUBS 0.007188f
C309 B.n26 VSUBS 0.007188f
C310 B.n27 VSUBS 0.007188f
C311 B.n28 VSUBS 0.007188f
C312 B.n29 VSUBS 0.007188f
C313 B.n30 VSUBS 0.007188f
C314 B.n31 VSUBS 0.007188f
C315 B.n32 VSUBS 0.007188f
C316 B.n33 VSUBS 0.007188f
C317 B.n34 VSUBS 0.007188f
C318 B.n35 VSUBS 0.007188f
C319 B.n36 VSUBS 0.007188f
C320 B.n37 VSUBS 0.007188f
C321 B.n38 VSUBS 0.007188f
C322 B.n39 VSUBS 0.007188f
C323 B.n40 VSUBS 0.007188f
C324 B.n41 VSUBS 0.007188f
C325 B.n42 VSUBS 0.007188f
C326 B.n43 VSUBS 0.007188f
C327 B.n44 VSUBS 0.007188f
C328 B.n45 VSUBS 0.007188f
C329 B.n46 VSUBS 0.007188f
C330 B.n47 VSUBS 0.007188f
C331 B.n48 VSUBS 0.007188f
C332 B.n49 VSUBS 0.007188f
C333 B.n50 VSUBS 0.007188f
C334 B.n51 VSUBS 0.007188f
C335 B.t7 VSUBS 0.347059f
C336 B.t8 VSUBS 0.381507f
C337 B.t6 VSUBS 2.08068f
C338 B.n52 VSUBS 0.586145f
C339 B.n53 VSUBS 0.331007f
C340 B.n54 VSUBS 0.016654f
C341 B.n55 VSUBS 0.007188f
C342 B.n56 VSUBS 0.007188f
C343 B.n57 VSUBS 0.007188f
C344 B.n58 VSUBS 0.007188f
C345 B.n59 VSUBS 0.007188f
C346 B.t10 VSUBS 0.347063f
C347 B.t11 VSUBS 0.38151f
C348 B.t9 VSUBS 2.08068f
C349 B.n60 VSUBS 0.586141f
C350 B.n61 VSUBS 0.331003f
C351 B.n62 VSUBS 0.007188f
C352 B.n63 VSUBS 0.007188f
C353 B.n64 VSUBS 0.007188f
C354 B.n65 VSUBS 0.007188f
C355 B.n66 VSUBS 0.007188f
C356 B.n67 VSUBS 0.007188f
C357 B.n68 VSUBS 0.007188f
C358 B.n69 VSUBS 0.007188f
C359 B.n70 VSUBS 0.007188f
C360 B.n71 VSUBS 0.007188f
C361 B.n72 VSUBS 0.007188f
C362 B.n73 VSUBS 0.007188f
C363 B.n74 VSUBS 0.007188f
C364 B.n75 VSUBS 0.007188f
C365 B.n76 VSUBS 0.007188f
C366 B.n77 VSUBS 0.007188f
C367 B.n78 VSUBS 0.007188f
C368 B.n79 VSUBS 0.007188f
C369 B.n80 VSUBS 0.007188f
C370 B.n81 VSUBS 0.007188f
C371 B.n82 VSUBS 0.007188f
C372 B.n83 VSUBS 0.007188f
C373 B.n84 VSUBS 0.007188f
C374 B.n85 VSUBS 0.007188f
C375 B.n86 VSUBS 0.007188f
C376 B.n87 VSUBS 0.007188f
C377 B.n88 VSUBS 0.007188f
C378 B.n89 VSUBS 0.007188f
C379 B.n90 VSUBS 0.016792f
C380 B.n91 VSUBS 0.007188f
C381 B.n92 VSUBS 0.007188f
C382 B.n93 VSUBS 0.007188f
C383 B.n94 VSUBS 0.007188f
C384 B.n95 VSUBS 0.007188f
C385 B.n96 VSUBS 0.007188f
C386 B.n97 VSUBS 0.007188f
C387 B.n98 VSUBS 0.007188f
C388 B.n99 VSUBS 0.007188f
C389 B.n100 VSUBS 0.007188f
C390 B.n101 VSUBS 0.007188f
C391 B.n102 VSUBS 0.007188f
C392 B.n103 VSUBS 0.007188f
C393 B.n104 VSUBS 0.007188f
C394 B.n105 VSUBS 0.007188f
C395 B.n106 VSUBS 0.007188f
C396 B.n107 VSUBS 0.007188f
C397 B.n108 VSUBS 0.007188f
C398 B.n109 VSUBS 0.007188f
C399 B.n110 VSUBS 0.007188f
C400 B.n111 VSUBS 0.007188f
C401 B.n112 VSUBS 0.007188f
C402 B.n113 VSUBS 0.007188f
C403 B.n114 VSUBS 0.007188f
C404 B.n115 VSUBS 0.007188f
C405 B.n116 VSUBS 0.007188f
C406 B.n117 VSUBS 0.007188f
C407 B.n118 VSUBS 0.007188f
C408 B.n119 VSUBS 0.007188f
C409 B.n120 VSUBS 0.007188f
C410 B.n121 VSUBS 0.007188f
C411 B.n122 VSUBS 0.007188f
C412 B.n123 VSUBS 0.007188f
C413 B.n124 VSUBS 0.007188f
C414 B.n125 VSUBS 0.007188f
C415 B.n126 VSUBS 0.007188f
C416 B.n127 VSUBS 0.007188f
C417 B.n128 VSUBS 0.007188f
C418 B.n129 VSUBS 0.007188f
C419 B.n130 VSUBS 0.007188f
C420 B.n131 VSUBS 0.007188f
C421 B.n132 VSUBS 0.007188f
C422 B.n133 VSUBS 0.017881f
C423 B.n134 VSUBS 0.007188f
C424 B.n135 VSUBS 0.007188f
C425 B.n136 VSUBS 0.007188f
C426 B.n137 VSUBS 0.007188f
C427 B.n138 VSUBS 0.007188f
C428 B.n139 VSUBS 0.007188f
C429 B.n140 VSUBS 0.007188f
C430 B.n141 VSUBS 0.007188f
C431 B.n142 VSUBS 0.007188f
C432 B.n143 VSUBS 0.007188f
C433 B.n144 VSUBS 0.007188f
C434 B.n145 VSUBS 0.007188f
C435 B.n146 VSUBS 0.007188f
C436 B.n147 VSUBS 0.007188f
C437 B.n148 VSUBS 0.007188f
C438 B.n149 VSUBS 0.007188f
C439 B.n150 VSUBS 0.007188f
C440 B.n151 VSUBS 0.007188f
C441 B.n152 VSUBS 0.007188f
C442 B.n153 VSUBS 0.007188f
C443 B.n154 VSUBS 0.007188f
C444 B.n155 VSUBS 0.007188f
C445 B.n156 VSUBS 0.007188f
C446 B.n157 VSUBS 0.007188f
C447 B.n158 VSUBS 0.007188f
C448 B.n159 VSUBS 0.007188f
C449 B.n160 VSUBS 0.007188f
C450 B.n161 VSUBS 0.007188f
C451 B.t2 VSUBS 0.347063f
C452 B.t1 VSUBS 0.38151f
C453 B.t0 VSUBS 2.08068f
C454 B.n162 VSUBS 0.586141f
C455 B.n163 VSUBS 0.331003f
C456 B.n164 VSUBS 0.016654f
C457 B.n165 VSUBS 0.007188f
C458 B.n166 VSUBS 0.007188f
C459 B.n167 VSUBS 0.007188f
C460 B.n168 VSUBS 0.007188f
C461 B.n169 VSUBS 0.007188f
C462 B.t5 VSUBS 0.347059f
C463 B.t4 VSUBS 0.381507f
C464 B.t3 VSUBS 2.08068f
C465 B.n170 VSUBS 0.586145f
C466 B.n171 VSUBS 0.331007f
C467 B.n172 VSUBS 0.007188f
C468 B.n173 VSUBS 0.007188f
C469 B.n174 VSUBS 0.007188f
C470 B.n175 VSUBS 0.007188f
C471 B.n176 VSUBS 0.007188f
C472 B.n177 VSUBS 0.007188f
C473 B.n178 VSUBS 0.007188f
C474 B.n179 VSUBS 0.007188f
C475 B.n180 VSUBS 0.007188f
C476 B.n181 VSUBS 0.007188f
C477 B.n182 VSUBS 0.007188f
C478 B.n183 VSUBS 0.007188f
C479 B.n184 VSUBS 0.007188f
C480 B.n185 VSUBS 0.007188f
C481 B.n186 VSUBS 0.007188f
C482 B.n187 VSUBS 0.007188f
C483 B.n188 VSUBS 0.007188f
C484 B.n189 VSUBS 0.007188f
C485 B.n190 VSUBS 0.007188f
C486 B.n191 VSUBS 0.007188f
C487 B.n192 VSUBS 0.007188f
C488 B.n193 VSUBS 0.007188f
C489 B.n194 VSUBS 0.007188f
C490 B.n195 VSUBS 0.007188f
C491 B.n196 VSUBS 0.007188f
C492 B.n197 VSUBS 0.007188f
C493 B.n198 VSUBS 0.007188f
C494 B.n199 VSUBS 0.007188f
C495 B.n200 VSUBS 0.016792f
C496 B.n201 VSUBS 0.007188f
C497 B.n202 VSUBS 0.007188f
C498 B.n203 VSUBS 0.007188f
C499 B.n204 VSUBS 0.007188f
C500 B.n205 VSUBS 0.007188f
C501 B.n206 VSUBS 0.007188f
C502 B.n207 VSUBS 0.007188f
C503 B.n208 VSUBS 0.007188f
C504 B.n209 VSUBS 0.007188f
C505 B.n210 VSUBS 0.007188f
C506 B.n211 VSUBS 0.007188f
C507 B.n212 VSUBS 0.007188f
C508 B.n213 VSUBS 0.007188f
C509 B.n214 VSUBS 0.007188f
C510 B.n215 VSUBS 0.007188f
C511 B.n216 VSUBS 0.007188f
C512 B.n217 VSUBS 0.007188f
C513 B.n218 VSUBS 0.007188f
C514 B.n219 VSUBS 0.007188f
C515 B.n220 VSUBS 0.007188f
C516 B.n221 VSUBS 0.007188f
C517 B.n222 VSUBS 0.007188f
C518 B.n223 VSUBS 0.007188f
C519 B.n224 VSUBS 0.007188f
C520 B.n225 VSUBS 0.007188f
C521 B.n226 VSUBS 0.007188f
C522 B.n227 VSUBS 0.007188f
C523 B.n228 VSUBS 0.007188f
C524 B.n229 VSUBS 0.007188f
C525 B.n230 VSUBS 0.007188f
C526 B.n231 VSUBS 0.007188f
C527 B.n232 VSUBS 0.007188f
C528 B.n233 VSUBS 0.007188f
C529 B.n234 VSUBS 0.007188f
C530 B.n235 VSUBS 0.007188f
C531 B.n236 VSUBS 0.007188f
C532 B.n237 VSUBS 0.007188f
C533 B.n238 VSUBS 0.007188f
C534 B.n239 VSUBS 0.007188f
C535 B.n240 VSUBS 0.007188f
C536 B.n241 VSUBS 0.007188f
C537 B.n242 VSUBS 0.007188f
C538 B.n243 VSUBS 0.007188f
C539 B.n244 VSUBS 0.007188f
C540 B.n245 VSUBS 0.007188f
C541 B.n246 VSUBS 0.007188f
C542 B.n247 VSUBS 0.007188f
C543 B.n248 VSUBS 0.007188f
C544 B.n249 VSUBS 0.007188f
C545 B.n250 VSUBS 0.007188f
C546 B.n251 VSUBS 0.007188f
C547 B.n252 VSUBS 0.007188f
C548 B.n253 VSUBS 0.007188f
C549 B.n254 VSUBS 0.007188f
C550 B.n255 VSUBS 0.007188f
C551 B.n256 VSUBS 0.007188f
C552 B.n257 VSUBS 0.007188f
C553 B.n258 VSUBS 0.007188f
C554 B.n259 VSUBS 0.007188f
C555 B.n260 VSUBS 0.007188f
C556 B.n261 VSUBS 0.007188f
C557 B.n262 VSUBS 0.007188f
C558 B.n263 VSUBS 0.007188f
C559 B.n264 VSUBS 0.007188f
C560 B.n265 VSUBS 0.007188f
C561 B.n266 VSUBS 0.007188f
C562 B.n267 VSUBS 0.007188f
C563 B.n268 VSUBS 0.007188f
C564 B.n269 VSUBS 0.007188f
C565 B.n270 VSUBS 0.007188f
C566 B.n271 VSUBS 0.007188f
C567 B.n272 VSUBS 0.007188f
C568 B.n273 VSUBS 0.007188f
C569 B.n274 VSUBS 0.007188f
C570 B.n275 VSUBS 0.007188f
C571 B.n276 VSUBS 0.007188f
C572 B.n277 VSUBS 0.007188f
C573 B.n278 VSUBS 0.007188f
C574 B.n279 VSUBS 0.007188f
C575 B.n280 VSUBS 0.007188f
C576 B.n281 VSUBS 0.016792f
C577 B.n282 VSUBS 0.017881f
C578 B.n283 VSUBS 0.017881f
C579 B.n284 VSUBS 0.007188f
C580 B.n285 VSUBS 0.007188f
C581 B.n286 VSUBS 0.007188f
C582 B.n287 VSUBS 0.007188f
C583 B.n288 VSUBS 0.007188f
C584 B.n289 VSUBS 0.007188f
C585 B.n290 VSUBS 0.007188f
C586 B.n291 VSUBS 0.007188f
C587 B.n292 VSUBS 0.007188f
C588 B.n293 VSUBS 0.007188f
C589 B.n294 VSUBS 0.007188f
C590 B.n295 VSUBS 0.007188f
C591 B.n296 VSUBS 0.007188f
C592 B.n297 VSUBS 0.007188f
C593 B.n298 VSUBS 0.007188f
C594 B.n299 VSUBS 0.007188f
C595 B.n300 VSUBS 0.007188f
C596 B.n301 VSUBS 0.007188f
C597 B.n302 VSUBS 0.007188f
C598 B.n303 VSUBS 0.007188f
C599 B.n304 VSUBS 0.007188f
C600 B.n305 VSUBS 0.007188f
C601 B.n306 VSUBS 0.007188f
C602 B.n307 VSUBS 0.007188f
C603 B.n308 VSUBS 0.007188f
C604 B.n309 VSUBS 0.007188f
C605 B.n310 VSUBS 0.007188f
C606 B.n311 VSUBS 0.007188f
C607 B.n312 VSUBS 0.007188f
C608 B.n313 VSUBS 0.007188f
C609 B.n314 VSUBS 0.007188f
C610 B.n315 VSUBS 0.007188f
C611 B.n316 VSUBS 0.007188f
C612 B.n317 VSUBS 0.007188f
C613 B.n318 VSUBS 0.007188f
C614 B.n319 VSUBS 0.007188f
C615 B.n320 VSUBS 0.007188f
C616 B.n321 VSUBS 0.007188f
C617 B.n322 VSUBS 0.007188f
C618 B.n323 VSUBS 0.007188f
C619 B.n324 VSUBS 0.007188f
C620 B.n325 VSUBS 0.007188f
C621 B.n326 VSUBS 0.007188f
C622 B.n327 VSUBS 0.007188f
C623 B.n328 VSUBS 0.007188f
C624 B.n329 VSUBS 0.007188f
C625 B.n330 VSUBS 0.007188f
C626 B.n331 VSUBS 0.007188f
C627 B.n332 VSUBS 0.007188f
C628 B.n333 VSUBS 0.007188f
C629 B.n334 VSUBS 0.007188f
C630 B.n335 VSUBS 0.007188f
C631 B.n336 VSUBS 0.007188f
C632 B.n337 VSUBS 0.007188f
C633 B.n338 VSUBS 0.007188f
C634 B.n339 VSUBS 0.007188f
C635 B.n340 VSUBS 0.007188f
C636 B.n341 VSUBS 0.007188f
C637 B.n342 VSUBS 0.007188f
C638 B.n343 VSUBS 0.007188f
C639 B.n344 VSUBS 0.007188f
C640 B.n345 VSUBS 0.007188f
C641 B.n346 VSUBS 0.007188f
C642 B.n347 VSUBS 0.007188f
C643 B.n348 VSUBS 0.007188f
C644 B.n349 VSUBS 0.007188f
C645 B.n350 VSUBS 0.007188f
C646 B.n351 VSUBS 0.007188f
C647 B.n352 VSUBS 0.007188f
C648 B.n353 VSUBS 0.007188f
C649 B.n354 VSUBS 0.007188f
C650 B.n355 VSUBS 0.007188f
C651 B.n356 VSUBS 0.007188f
C652 B.n357 VSUBS 0.007188f
C653 B.n358 VSUBS 0.007188f
C654 B.n359 VSUBS 0.007188f
C655 B.n360 VSUBS 0.007188f
C656 B.n361 VSUBS 0.007188f
C657 B.n362 VSUBS 0.007188f
C658 B.n363 VSUBS 0.007188f
C659 B.n364 VSUBS 0.007188f
C660 B.n365 VSUBS 0.007188f
C661 B.n366 VSUBS 0.007188f
C662 B.n367 VSUBS 0.007188f
C663 B.n368 VSUBS 0.004968f
C664 B.n369 VSUBS 0.016654f
C665 B.n370 VSUBS 0.005814f
C666 B.n371 VSUBS 0.007188f
C667 B.n372 VSUBS 0.007188f
C668 B.n373 VSUBS 0.007188f
C669 B.n374 VSUBS 0.007188f
C670 B.n375 VSUBS 0.007188f
C671 B.n376 VSUBS 0.007188f
C672 B.n377 VSUBS 0.007188f
C673 B.n378 VSUBS 0.007188f
C674 B.n379 VSUBS 0.007188f
C675 B.n380 VSUBS 0.007188f
C676 B.n381 VSUBS 0.007188f
C677 B.n382 VSUBS 0.005814f
C678 B.n383 VSUBS 0.007188f
C679 B.n384 VSUBS 0.007188f
C680 B.n385 VSUBS 0.004968f
C681 B.n386 VSUBS 0.007188f
C682 B.n387 VSUBS 0.007188f
C683 B.n388 VSUBS 0.007188f
C684 B.n389 VSUBS 0.007188f
C685 B.n390 VSUBS 0.007188f
C686 B.n391 VSUBS 0.007188f
C687 B.n392 VSUBS 0.007188f
C688 B.n393 VSUBS 0.007188f
C689 B.n394 VSUBS 0.007188f
C690 B.n395 VSUBS 0.007188f
C691 B.n396 VSUBS 0.007188f
C692 B.n397 VSUBS 0.007188f
C693 B.n398 VSUBS 0.007188f
C694 B.n399 VSUBS 0.007188f
C695 B.n400 VSUBS 0.007188f
C696 B.n401 VSUBS 0.007188f
C697 B.n402 VSUBS 0.007188f
C698 B.n403 VSUBS 0.007188f
C699 B.n404 VSUBS 0.007188f
C700 B.n405 VSUBS 0.007188f
C701 B.n406 VSUBS 0.007188f
C702 B.n407 VSUBS 0.007188f
C703 B.n408 VSUBS 0.007188f
C704 B.n409 VSUBS 0.007188f
C705 B.n410 VSUBS 0.007188f
C706 B.n411 VSUBS 0.007188f
C707 B.n412 VSUBS 0.007188f
C708 B.n413 VSUBS 0.007188f
C709 B.n414 VSUBS 0.007188f
C710 B.n415 VSUBS 0.007188f
C711 B.n416 VSUBS 0.007188f
C712 B.n417 VSUBS 0.007188f
C713 B.n418 VSUBS 0.007188f
C714 B.n419 VSUBS 0.007188f
C715 B.n420 VSUBS 0.007188f
C716 B.n421 VSUBS 0.007188f
C717 B.n422 VSUBS 0.007188f
C718 B.n423 VSUBS 0.007188f
C719 B.n424 VSUBS 0.007188f
C720 B.n425 VSUBS 0.007188f
C721 B.n426 VSUBS 0.007188f
C722 B.n427 VSUBS 0.007188f
C723 B.n428 VSUBS 0.007188f
C724 B.n429 VSUBS 0.007188f
C725 B.n430 VSUBS 0.007188f
C726 B.n431 VSUBS 0.007188f
C727 B.n432 VSUBS 0.007188f
C728 B.n433 VSUBS 0.007188f
C729 B.n434 VSUBS 0.007188f
C730 B.n435 VSUBS 0.007188f
C731 B.n436 VSUBS 0.007188f
C732 B.n437 VSUBS 0.007188f
C733 B.n438 VSUBS 0.007188f
C734 B.n439 VSUBS 0.007188f
C735 B.n440 VSUBS 0.007188f
C736 B.n441 VSUBS 0.007188f
C737 B.n442 VSUBS 0.007188f
C738 B.n443 VSUBS 0.007188f
C739 B.n444 VSUBS 0.007188f
C740 B.n445 VSUBS 0.007188f
C741 B.n446 VSUBS 0.007188f
C742 B.n447 VSUBS 0.007188f
C743 B.n448 VSUBS 0.007188f
C744 B.n449 VSUBS 0.007188f
C745 B.n450 VSUBS 0.007188f
C746 B.n451 VSUBS 0.007188f
C747 B.n452 VSUBS 0.007188f
C748 B.n453 VSUBS 0.007188f
C749 B.n454 VSUBS 0.007188f
C750 B.n455 VSUBS 0.007188f
C751 B.n456 VSUBS 0.007188f
C752 B.n457 VSUBS 0.007188f
C753 B.n458 VSUBS 0.007188f
C754 B.n459 VSUBS 0.007188f
C755 B.n460 VSUBS 0.007188f
C756 B.n461 VSUBS 0.007188f
C757 B.n462 VSUBS 0.007188f
C758 B.n463 VSUBS 0.007188f
C759 B.n464 VSUBS 0.007188f
C760 B.n465 VSUBS 0.007188f
C761 B.n466 VSUBS 0.007188f
C762 B.n467 VSUBS 0.007188f
C763 B.n468 VSUBS 0.007188f
C764 B.n469 VSUBS 0.007188f
C765 B.n470 VSUBS 0.017069f
C766 B.n471 VSUBS 0.017604f
C767 B.n472 VSUBS 0.016792f
C768 B.n473 VSUBS 0.007188f
C769 B.n474 VSUBS 0.007188f
C770 B.n475 VSUBS 0.007188f
C771 B.n476 VSUBS 0.007188f
C772 B.n477 VSUBS 0.007188f
C773 B.n478 VSUBS 0.007188f
C774 B.n479 VSUBS 0.007188f
C775 B.n480 VSUBS 0.007188f
C776 B.n481 VSUBS 0.007188f
C777 B.n482 VSUBS 0.007188f
C778 B.n483 VSUBS 0.007188f
C779 B.n484 VSUBS 0.007188f
C780 B.n485 VSUBS 0.007188f
C781 B.n486 VSUBS 0.007188f
C782 B.n487 VSUBS 0.007188f
C783 B.n488 VSUBS 0.007188f
C784 B.n489 VSUBS 0.007188f
C785 B.n490 VSUBS 0.007188f
C786 B.n491 VSUBS 0.007188f
C787 B.n492 VSUBS 0.007188f
C788 B.n493 VSUBS 0.007188f
C789 B.n494 VSUBS 0.007188f
C790 B.n495 VSUBS 0.007188f
C791 B.n496 VSUBS 0.007188f
C792 B.n497 VSUBS 0.007188f
C793 B.n498 VSUBS 0.007188f
C794 B.n499 VSUBS 0.007188f
C795 B.n500 VSUBS 0.007188f
C796 B.n501 VSUBS 0.007188f
C797 B.n502 VSUBS 0.007188f
C798 B.n503 VSUBS 0.007188f
C799 B.n504 VSUBS 0.007188f
C800 B.n505 VSUBS 0.007188f
C801 B.n506 VSUBS 0.007188f
C802 B.n507 VSUBS 0.007188f
C803 B.n508 VSUBS 0.007188f
C804 B.n509 VSUBS 0.007188f
C805 B.n510 VSUBS 0.007188f
C806 B.n511 VSUBS 0.007188f
C807 B.n512 VSUBS 0.007188f
C808 B.n513 VSUBS 0.007188f
C809 B.n514 VSUBS 0.007188f
C810 B.n515 VSUBS 0.007188f
C811 B.n516 VSUBS 0.007188f
C812 B.n517 VSUBS 0.007188f
C813 B.n518 VSUBS 0.007188f
C814 B.n519 VSUBS 0.007188f
C815 B.n520 VSUBS 0.007188f
C816 B.n521 VSUBS 0.007188f
C817 B.n522 VSUBS 0.007188f
C818 B.n523 VSUBS 0.007188f
C819 B.n524 VSUBS 0.007188f
C820 B.n525 VSUBS 0.007188f
C821 B.n526 VSUBS 0.007188f
C822 B.n527 VSUBS 0.007188f
C823 B.n528 VSUBS 0.007188f
C824 B.n529 VSUBS 0.007188f
C825 B.n530 VSUBS 0.007188f
C826 B.n531 VSUBS 0.007188f
C827 B.n532 VSUBS 0.007188f
C828 B.n533 VSUBS 0.007188f
C829 B.n534 VSUBS 0.007188f
C830 B.n535 VSUBS 0.007188f
C831 B.n536 VSUBS 0.007188f
C832 B.n537 VSUBS 0.007188f
C833 B.n538 VSUBS 0.007188f
C834 B.n539 VSUBS 0.007188f
C835 B.n540 VSUBS 0.007188f
C836 B.n541 VSUBS 0.007188f
C837 B.n542 VSUBS 0.007188f
C838 B.n543 VSUBS 0.007188f
C839 B.n544 VSUBS 0.007188f
C840 B.n545 VSUBS 0.007188f
C841 B.n546 VSUBS 0.007188f
C842 B.n547 VSUBS 0.007188f
C843 B.n548 VSUBS 0.007188f
C844 B.n549 VSUBS 0.007188f
C845 B.n550 VSUBS 0.007188f
C846 B.n551 VSUBS 0.007188f
C847 B.n552 VSUBS 0.007188f
C848 B.n553 VSUBS 0.007188f
C849 B.n554 VSUBS 0.007188f
C850 B.n555 VSUBS 0.007188f
C851 B.n556 VSUBS 0.007188f
C852 B.n557 VSUBS 0.007188f
C853 B.n558 VSUBS 0.007188f
C854 B.n559 VSUBS 0.007188f
C855 B.n560 VSUBS 0.007188f
C856 B.n561 VSUBS 0.007188f
C857 B.n562 VSUBS 0.007188f
C858 B.n563 VSUBS 0.007188f
C859 B.n564 VSUBS 0.007188f
C860 B.n565 VSUBS 0.007188f
C861 B.n566 VSUBS 0.007188f
C862 B.n567 VSUBS 0.007188f
C863 B.n568 VSUBS 0.007188f
C864 B.n569 VSUBS 0.007188f
C865 B.n570 VSUBS 0.007188f
C866 B.n571 VSUBS 0.007188f
C867 B.n572 VSUBS 0.007188f
C868 B.n573 VSUBS 0.007188f
C869 B.n574 VSUBS 0.007188f
C870 B.n575 VSUBS 0.007188f
C871 B.n576 VSUBS 0.007188f
C872 B.n577 VSUBS 0.007188f
C873 B.n578 VSUBS 0.007188f
C874 B.n579 VSUBS 0.007188f
C875 B.n580 VSUBS 0.007188f
C876 B.n581 VSUBS 0.007188f
C877 B.n582 VSUBS 0.007188f
C878 B.n583 VSUBS 0.007188f
C879 B.n584 VSUBS 0.007188f
C880 B.n585 VSUBS 0.007188f
C881 B.n586 VSUBS 0.007188f
C882 B.n587 VSUBS 0.007188f
C883 B.n588 VSUBS 0.007188f
C884 B.n589 VSUBS 0.007188f
C885 B.n590 VSUBS 0.007188f
C886 B.n591 VSUBS 0.007188f
C887 B.n592 VSUBS 0.007188f
C888 B.n593 VSUBS 0.007188f
C889 B.n594 VSUBS 0.007188f
C890 B.n595 VSUBS 0.007188f
C891 B.n596 VSUBS 0.007188f
C892 B.n597 VSUBS 0.007188f
C893 B.n598 VSUBS 0.007188f
C894 B.n599 VSUBS 0.016792f
C895 B.n600 VSUBS 0.017881f
C896 B.n601 VSUBS 0.017881f
C897 B.n602 VSUBS 0.007188f
C898 B.n603 VSUBS 0.007188f
C899 B.n604 VSUBS 0.007188f
C900 B.n605 VSUBS 0.007188f
C901 B.n606 VSUBS 0.007188f
C902 B.n607 VSUBS 0.007188f
C903 B.n608 VSUBS 0.007188f
C904 B.n609 VSUBS 0.007188f
C905 B.n610 VSUBS 0.007188f
C906 B.n611 VSUBS 0.007188f
C907 B.n612 VSUBS 0.007188f
C908 B.n613 VSUBS 0.007188f
C909 B.n614 VSUBS 0.007188f
C910 B.n615 VSUBS 0.007188f
C911 B.n616 VSUBS 0.007188f
C912 B.n617 VSUBS 0.007188f
C913 B.n618 VSUBS 0.007188f
C914 B.n619 VSUBS 0.007188f
C915 B.n620 VSUBS 0.007188f
C916 B.n621 VSUBS 0.007188f
C917 B.n622 VSUBS 0.007188f
C918 B.n623 VSUBS 0.007188f
C919 B.n624 VSUBS 0.007188f
C920 B.n625 VSUBS 0.007188f
C921 B.n626 VSUBS 0.007188f
C922 B.n627 VSUBS 0.007188f
C923 B.n628 VSUBS 0.007188f
C924 B.n629 VSUBS 0.007188f
C925 B.n630 VSUBS 0.007188f
C926 B.n631 VSUBS 0.007188f
C927 B.n632 VSUBS 0.007188f
C928 B.n633 VSUBS 0.007188f
C929 B.n634 VSUBS 0.007188f
C930 B.n635 VSUBS 0.007188f
C931 B.n636 VSUBS 0.007188f
C932 B.n637 VSUBS 0.007188f
C933 B.n638 VSUBS 0.007188f
C934 B.n639 VSUBS 0.007188f
C935 B.n640 VSUBS 0.007188f
C936 B.n641 VSUBS 0.007188f
C937 B.n642 VSUBS 0.007188f
C938 B.n643 VSUBS 0.007188f
C939 B.n644 VSUBS 0.007188f
C940 B.n645 VSUBS 0.007188f
C941 B.n646 VSUBS 0.007188f
C942 B.n647 VSUBS 0.007188f
C943 B.n648 VSUBS 0.007188f
C944 B.n649 VSUBS 0.007188f
C945 B.n650 VSUBS 0.007188f
C946 B.n651 VSUBS 0.007188f
C947 B.n652 VSUBS 0.007188f
C948 B.n653 VSUBS 0.007188f
C949 B.n654 VSUBS 0.007188f
C950 B.n655 VSUBS 0.007188f
C951 B.n656 VSUBS 0.007188f
C952 B.n657 VSUBS 0.007188f
C953 B.n658 VSUBS 0.007188f
C954 B.n659 VSUBS 0.007188f
C955 B.n660 VSUBS 0.007188f
C956 B.n661 VSUBS 0.007188f
C957 B.n662 VSUBS 0.007188f
C958 B.n663 VSUBS 0.007188f
C959 B.n664 VSUBS 0.007188f
C960 B.n665 VSUBS 0.007188f
C961 B.n666 VSUBS 0.007188f
C962 B.n667 VSUBS 0.007188f
C963 B.n668 VSUBS 0.007188f
C964 B.n669 VSUBS 0.007188f
C965 B.n670 VSUBS 0.007188f
C966 B.n671 VSUBS 0.007188f
C967 B.n672 VSUBS 0.007188f
C968 B.n673 VSUBS 0.007188f
C969 B.n674 VSUBS 0.007188f
C970 B.n675 VSUBS 0.007188f
C971 B.n676 VSUBS 0.007188f
C972 B.n677 VSUBS 0.007188f
C973 B.n678 VSUBS 0.007188f
C974 B.n679 VSUBS 0.007188f
C975 B.n680 VSUBS 0.007188f
C976 B.n681 VSUBS 0.007188f
C977 B.n682 VSUBS 0.007188f
C978 B.n683 VSUBS 0.007188f
C979 B.n684 VSUBS 0.007188f
C980 B.n685 VSUBS 0.007188f
C981 B.n686 VSUBS 0.004968f
C982 B.n687 VSUBS 0.016654f
C983 B.n688 VSUBS 0.005814f
C984 B.n689 VSUBS 0.007188f
C985 B.n690 VSUBS 0.007188f
C986 B.n691 VSUBS 0.007188f
C987 B.n692 VSUBS 0.007188f
C988 B.n693 VSUBS 0.007188f
C989 B.n694 VSUBS 0.007188f
C990 B.n695 VSUBS 0.007188f
C991 B.n696 VSUBS 0.007188f
C992 B.n697 VSUBS 0.007188f
C993 B.n698 VSUBS 0.007188f
C994 B.n699 VSUBS 0.007188f
C995 B.n700 VSUBS 0.005814f
C996 B.n701 VSUBS 0.007188f
C997 B.n702 VSUBS 0.007188f
C998 B.n703 VSUBS 0.004968f
C999 B.n704 VSUBS 0.007188f
C1000 B.n705 VSUBS 0.007188f
C1001 B.n706 VSUBS 0.007188f
C1002 B.n707 VSUBS 0.007188f
C1003 B.n708 VSUBS 0.007188f
C1004 B.n709 VSUBS 0.007188f
C1005 B.n710 VSUBS 0.007188f
C1006 B.n711 VSUBS 0.007188f
C1007 B.n712 VSUBS 0.007188f
C1008 B.n713 VSUBS 0.007188f
C1009 B.n714 VSUBS 0.007188f
C1010 B.n715 VSUBS 0.007188f
C1011 B.n716 VSUBS 0.007188f
C1012 B.n717 VSUBS 0.007188f
C1013 B.n718 VSUBS 0.007188f
C1014 B.n719 VSUBS 0.007188f
C1015 B.n720 VSUBS 0.007188f
C1016 B.n721 VSUBS 0.007188f
C1017 B.n722 VSUBS 0.007188f
C1018 B.n723 VSUBS 0.007188f
C1019 B.n724 VSUBS 0.007188f
C1020 B.n725 VSUBS 0.007188f
C1021 B.n726 VSUBS 0.007188f
C1022 B.n727 VSUBS 0.007188f
C1023 B.n728 VSUBS 0.007188f
C1024 B.n729 VSUBS 0.007188f
C1025 B.n730 VSUBS 0.007188f
C1026 B.n731 VSUBS 0.007188f
C1027 B.n732 VSUBS 0.007188f
C1028 B.n733 VSUBS 0.007188f
C1029 B.n734 VSUBS 0.007188f
C1030 B.n735 VSUBS 0.007188f
C1031 B.n736 VSUBS 0.007188f
C1032 B.n737 VSUBS 0.007188f
C1033 B.n738 VSUBS 0.007188f
C1034 B.n739 VSUBS 0.007188f
C1035 B.n740 VSUBS 0.007188f
C1036 B.n741 VSUBS 0.007188f
C1037 B.n742 VSUBS 0.007188f
C1038 B.n743 VSUBS 0.007188f
C1039 B.n744 VSUBS 0.007188f
C1040 B.n745 VSUBS 0.007188f
C1041 B.n746 VSUBS 0.007188f
C1042 B.n747 VSUBS 0.007188f
C1043 B.n748 VSUBS 0.007188f
C1044 B.n749 VSUBS 0.007188f
C1045 B.n750 VSUBS 0.007188f
C1046 B.n751 VSUBS 0.007188f
C1047 B.n752 VSUBS 0.007188f
C1048 B.n753 VSUBS 0.007188f
C1049 B.n754 VSUBS 0.007188f
C1050 B.n755 VSUBS 0.007188f
C1051 B.n756 VSUBS 0.007188f
C1052 B.n757 VSUBS 0.007188f
C1053 B.n758 VSUBS 0.007188f
C1054 B.n759 VSUBS 0.007188f
C1055 B.n760 VSUBS 0.007188f
C1056 B.n761 VSUBS 0.007188f
C1057 B.n762 VSUBS 0.007188f
C1058 B.n763 VSUBS 0.007188f
C1059 B.n764 VSUBS 0.007188f
C1060 B.n765 VSUBS 0.007188f
C1061 B.n766 VSUBS 0.007188f
C1062 B.n767 VSUBS 0.007188f
C1063 B.n768 VSUBS 0.007188f
C1064 B.n769 VSUBS 0.007188f
C1065 B.n770 VSUBS 0.007188f
C1066 B.n771 VSUBS 0.007188f
C1067 B.n772 VSUBS 0.007188f
C1068 B.n773 VSUBS 0.007188f
C1069 B.n774 VSUBS 0.007188f
C1070 B.n775 VSUBS 0.007188f
C1071 B.n776 VSUBS 0.007188f
C1072 B.n777 VSUBS 0.007188f
C1073 B.n778 VSUBS 0.007188f
C1074 B.n779 VSUBS 0.007188f
C1075 B.n780 VSUBS 0.007188f
C1076 B.n781 VSUBS 0.007188f
C1077 B.n782 VSUBS 0.007188f
C1078 B.n783 VSUBS 0.007188f
C1079 B.n784 VSUBS 0.007188f
C1080 B.n785 VSUBS 0.007188f
C1081 B.n786 VSUBS 0.007188f
C1082 B.n787 VSUBS 0.007188f
C1083 B.n788 VSUBS 0.017881f
C1084 B.n789 VSUBS 0.016792f
C1085 B.n790 VSUBS 0.016792f
C1086 B.n791 VSUBS 0.007188f
C1087 B.n792 VSUBS 0.007188f
C1088 B.n793 VSUBS 0.007188f
C1089 B.n794 VSUBS 0.007188f
C1090 B.n795 VSUBS 0.007188f
C1091 B.n796 VSUBS 0.007188f
C1092 B.n797 VSUBS 0.007188f
C1093 B.n798 VSUBS 0.007188f
C1094 B.n799 VSUBS 0.007188f
C1095 B.n800 VSUBS 0.007188f
C1096 B.n801 VSUBS 0.007188f
C1097 B.n802 VSUBS 0.007188f
C1098 B.n803 VSUBS 0.007188f
C1099 B.n804 VSUBS 0.007188f
C1100 B.n805 VSUBS 0.007188f
C1101 B.n806 VSUBS 0.007188f
C1102 B.n807 VSUBS 0.007188f
C1103 B.n808 VSUBS 0.007188f
C1104 B.n809 VSUBS 0.007188f
C1105 B.n810 VSUBS 0.007188f
C1106 B.n811 VSUBS 0.007188f
C1107 B.n812 VSUBS 0.007188f
C1108 B.n813 VSUBS 0.007188f
C1109 B.n814 VSUBS 0.007188f
C1110 B.n815 VSUBS 0.007188f
C1111 B.n816 VSUBS 0.007188f
C1112 B.n817 VSUBS 0.007188f
C1113 B.n818 VSUBS 0.007188f
C1114 B.n819 VSUBS 0.007188f
C1115 B.n820 VSUBS 0.007188f
C1116 B.n821 VSUBS 0.007188f
C1117 B.n822 VSUBS 0.007188f
C1118 B.n823 VSUBS 0.007188f
C1119 B.n824 VSUBS 0.007188f
C1120 B.n825 VSUBS 0.007188f
C1121 B.n826 VSUBS 0.007188f
C1122 B.n827 VSUBS 0.007188f
C1123 B.n828 VSUBS 0.007188f
C1124 B.n829 VSUBS 0.007188f
C1125 B.n830 VSUBS 0.007188f
C1126 B.n831 VSUBS 0.007188f
C1127 B.n832 VSUBS 0.007188f
C1128 B.n833 VSUBS 0.007188f
C1129 B.n834 VSUBS 0.007188f
C1130 B.n835 VSUBS 0.007188f
C1131 B.n836 VSUBS 0.007188f
C1132 B.n837 VSUBS 0.007188f
C1133 B.n838 VSUBS 0.007188f
C1134 B.n839 VSUBS 0.007188f
C1135 B.n840 VSUBS 0.007188f
C1136 B.n841 VSUBS 0.007188f
C1137 B.n842 VSUBS 0.007188f
C1138 B.n843 VSUBS 0.007188f
C1139 B.n844 VSUBS 0.007188f
C1140 B.n845 VSUBS 0.007188f
C1141 B.n846 VSUBS 0.007188f
C1142 B.n847 VSUBS 0.007188f
C1143 B.n848 VSUBS 0.007188f
C1144 B.n849 VSUBS 0.007188f
C1145 B.n850 VSUBS 0.007188f
C1146 B.n851 VSUBS 0.00938f
C1147 B.n852 VSUBS 0.009992f
C1148 B.n853 VSUBS 0.019871f
C1149 VDD2.n0 VSUBS 0.028559f
C1150 VDD2.n1 VSUBS 0.027142f
C1151 VDD2.n2 VSUBS 0.014585f
C1152 VDD2.n3 VSUBS 0.034473f
C1153 VDD2.n4 VSUBS 0.015443f
C1154 VDD2.n5 VSUBS 0.027142f
C1155 VDD2.n6 VSUBS 0.014585f
C1156 VDD2.n7 VSUBS 0.034473f
C1157 VDD2.n8 VSUBS 0.015014f
C1158 VDD2.n9 VSUBS 0.027142f
C1159 VDD2.n10 VSUBS 0.015443f
C1160 VDD2.n11 VSUBS 0.034473f
C1161 VDD2.n12 VSUBS 0.015443f
C1162 VDD2.n13 VSUBS 0.027142f
C1163 VDD2.n14 VSUBS 0.014585f
C1164 VDD2.n15 VSUBS 0.034473f
C1165 VDD2.n16 VSUBS 0.015443f
C1166 VDD2.n17 VSUBS 0.027142f
C1167 VDD2.n18 VSUBS 0.014585f
C1168 VDD2.n19 VSUBS 0.034473f
C1169 VDD2.n20 VSUBS 0.015443f
C1170 VDD2.n21 VSUBS 0.027142f
C1171 VDD2.n22 VSUBS 0.014585f
C1172 VDD2.n23 VSUBS 0.034473f
C1173 VDD2.n24 VSUBS 0.015443f
C1174 VDD2.n25 VSUBS 0.027142f
C1175 VDD2.n26 VSUBS 0.014585f
C1176 VDD2.n27 VSUBS 0.034473f
C1177 VDD2.n28 VSUBS 0.015443f
C1178 VDD2.n29 VSUBS 2.03615f
C1179 VDD2.n30 VSUBS 0.014585f
C1180 VDD2.t5 VSUBS 0.073966f
C1181 VDD2.n31 VSUBS 0.211018f
C1182 VDD2.n32 VSUBS 0.02193f
C1183 VDD2.n33 VSUBS 0.025855f
C1184 VDD2.n34 VSUBS 0.034473f
C1185 VDD2.n35 VSUBS 0.015443f
C1186 VDD2.n36 VSUBS 0.014585f
C1187 VDD2.n37 VSUBS 0.027142f
C1188 VDD2.n38 VSUBS 0.027142f
C1189 VDD2.n39 VSUBS 0.014585f
C1190 VDD2.n40 VSUBS 0.015443f
C1191 VDD2.n41 VSUBS 0.034473f
C1192 VDD2.n42 VSUBS 0.034473f
C1193 VDD2.n43 VSUBS 0.015443f
C1194 VDD2.n44 VSUBS 0.014585f
C1195 VDD2.n45 VSUBS 0.027142f
C1196 VDD2.n46 VSUBS 0.027142f
C1197 VDD2.n47 VSUBS 0.014585f
C1198 VDD2.n48 VSUBS 0.015443f
C1199 VDD2.n49 VSUBS 0.034473f
C1200 VDD2.n50 VSUBS 0.034473f
C1201 VDD2.n51 VSUBS 0.015443f
C1202 VDD2.n52 VSUBS 0.014585f
C1203 VDD2.n53 VSUBS 0.027142f
C1204 VDD2.n54 VSUBS 0.027142f
C1205 VDD2.n55 VSUBS 0.014585f
C1206 VDD2.n56 VSUBS 0.015443f
C1207 VDD2.n57 VSUBS 0.034473f
C1208 VDD2.n58 VSUBS 0.034473f
C1209 VDD2.n59 VSUBS 0.015443f
C1210 VDD2.n60 VSUBS 0.014585f
C1211 VDD2.n61 VSUBS 0.027142f
C1212 VDD2.n62 VSUBS 0.027142f
C1213 VDD2.n63 VSUBS 0.014585f
C1214 VDD2.n64 VSUBS 0.015443f
C1215 VDD2.n65 VSUBS 0.034473f
C1216 VDD2.n66 VSUBS 0.034473f
C1217 VDD2.n67 VSUBS 0.015443f
C1218 VDD2.n68 VSUBS 0.014585f
C1219 VDD2.n69 VSUBS 0.027142f
C1220 VDD2.n70 VSUBS 0.027142f
C1221 VDD2.n71 VSUBS 0.014585f
C1222 VDD2.n72 VSUBS 0.014585f
C1223 VDD2.n73 VSUBS 0.015443f
C1224 VDD2.n74 VSUBS 0.034473f
C1225 VDD2.n75 VSUBS 0.034473f
C1226 VDD2.n76 VSUBS 0.034473f
C1227 VDD2.n77 VSUBS 0.015014f
C1228 VDD2.n78 VSUBS 0.014585f
C1229 VDD2.n79 VSUBS 0.027142f
C1230 VDD2.n80 VSUBS 0.027142f
C1231 VDD2.n81 VSUBS 0.014585f
C1232 VDD2.n82 VSUBS 0.015443f
C1233 VDD2.n83 VSUBS 0.034473f
C1234 VDD2.n84 VSUBS 0.034473f
C1235 VDD2.n85 VSUBS 0.015443f
C1236 VDD2.n86 VSUBS 0.014585f
C1237 VDD2.n87 VSUBS 0.027142f
C1238 VDD2.n88 VSUBS 0.027142f
C1239 VDD2.n89 VSUBS 0.014585f
C1240 VDD2.n90 VSUBS 0.015443f
C1241 VDD2.n91 VSUBS 0.034473f
C1242 VDD2.n92 VSUBS 0.07915f
C1243 VDD2.n93 VSUBS 0.015443f
C1244 VDD2.n94 VSUBS 0.014585f
C1245 VDD2.n95 VSUBS 0.060512f
C1246 VDD2.n96 VSUBS 0.066226f
C1247 VDD2.t4 VSUBS 0.374484f
C1248 VDD2.t0 VSUBS 0.374484f
C1249 VDD2.n97 VSUBS 3.0997f
C1250 VDD2.n98 VSUBS 3.59462f
C1251 VDD2.n99 VSUBS 0.028559f
C1252 VDD2.n100 VSUBS 0.027142f
C1253 VDD2.n101 VSUBS 0.014585f
C1254 VDD2.n102 VSUBS 0.034473f
C1255 VDD2.n103 VSUBS 0.015443f
C1256 VDD2.n104 VSUBS 0.027142f
C1257 VDD2.n105 VSUBS 0.014585f
C1258 VDD2.n106 VSUBS 0.034473f
C1259 VDD2.n107 VSUBS 0.015014f
C1260 VDD2.n108 VSUBS 0.027142f
C1261 VDD2.n109 VSUBS 0.015014f
C1262 VDD2.n110 VSUBS 0.014585f
C1263 VDD2.n111 VSUBS 0.034473f
C1264 VDD2.n112 VSUBS 0.034473f
C1265 VDD2.n113 VSUBS 0.015443f
C1266 VDD2.n114 VSUBS 0.027142f
C1267 VDD2.n115 VSUBS 0.014585f
C1268 VDD2.n116 VSUBS 0.034473f
C1269 VDD2.n117 VSUBS 0.015443f
C1270 VDD2.n118 VSUBS 0.027142f
C1271 VDD2.n119 VSUBS 0.014585f
C1272 VDD2.n120 VSUBS 0.034473f
C1273 VDD2.n121 VSUBS 0.015443f
C1274 VDD2.n122 VSUBS 0.027142f
C1275 VDD2.n123 VSUBS 0.014585f
C1276 VDD2.n124 VSUBS 0.034473f
C1277 VDD2.n125 VSUBS 0.015443f
C1278 VDD2.n126 VSUBS 0.027142f
C1279 VDD2.n127 VSUBS 0.014585f
C1280 VDD2.n128 VSUBS 0.034473f
C1281 VDD2.n129 VSUBS 0.015443f
C1282 VDD2.n130 VSUBS 2.03615f
C1283 VDD2.n131 VSUBS 0.014585f
C1284 VDD2.t1 VSUBS 0.073966f
C1285 VDD2.n132 VSUBS 0.211018f
C1286 VDD2.n133 VSUBS 0.02193f
C1287 VDD2.n134 VSUBS 0.025855f
C1288 VDD2.n135 VSUBS 0.034473f
C1289 VDD2.n136 VSUBS 0.015443f
C1290 VDD2.n137 VSUBS 0.014585f
C1291 VDD2.n138 VSUBS 0.027142f
C1292 VDD2.n139 VSUBS 0.027142f
C1293 VDD2.n140 VSUBS 0.014585f
C1294 VDD2.n141 VSUBS 0.015443f
C1295 VDD2.n142 VSUBS 0.034473f
C1296 VDD2.n143 VSUBS 0.034473f
C1297 VDD2.n144 VSUBS 0.015443f
C1298 VDD2.n145 VSUBS 0.014585f
C1299 VDD2.n146 VSUBS 0.027142f
C1300 VDD2.n147 VSUBS 0.027142f
C1301 VDD2.n148 VSUBS 0.014585f
C1302 VDD2.n149 VSUBS 0.015443f
C1303 VDD2.n150 VSUBS 0.034473f
C1304 VDD2.n151 VSUBS 0.034473f
C1305 VDD2.n152 VSUBS 0.015443f
C1306 VDD2.n153 VSUBS 0.014585f
C1307 VDD2.n154 VSUBS 0.027142f
C1308 VDD2.n155 VSUBS 0.027142f
C1309 VDD2.n156 VSUBS 0.014585f
C1310 VDD2.n157 VSUBS 0.015443f
C1311 VDD2.n158 VSUBS 0.034473f
C1312 VDD2.n159 VSUBS 0.034473f
C1313 VDD2.n160 VSUBS 0.015443f
C1314 VDD2.n161 VSUBS 0.014585f
C1315 VDD2.n162 VSUBS 0.027142f
C1316 VDD2.n163 VSUBS 0.027142f
C1317 VDD2.n164 VSUBS 0.014585f
C1318 VDD2.n165 VSUBS 0.015443f
C1319 VDD2.n166 VSUBS 0.034473f
C1320 VDD2.n167 VSUBS 0.034473f
C1321 VDD2.n168 VSUBS 0.015443f
C1322 VDD2.n169 VSUBS 0.014585f
C1323 VDD2.n170 VSUBS 0.027142f
C1324 VDD2.n171 VSUBS 0.027142f
C1325 VDD2.n172 VSUBS 0.014585f
C1326 VDD2.n173 VSUBS 0.015443f
C1327 VDD2.n174 VSUBS 0.034473f
C1328 VDD2.n175 VSUBS 0.034473f
C1329 VDD2.n176 VSUBS 0.015443f
C1330 VDD2.n177 VSUBS 0.014585f
C1331 VDD2.n178 VSUBS 0.027142f
C1332 VDD2.n179 VSUBS 0.027142f
C1333 VDD2.n180 VSUBS 0.014585f
C1334 VDD2.n181 VSUBS 0.015443f
C1335 VDD2.n182 VSUBS 0.034473f
C1336 VDD2.n183 VSUBS 0.034473f
C1337 VDD2.n184 VSUBS 0.015443f
C1338 VDD2.n185 VSUBS 0.014585f
C1339 VDD2.n186 VSUBS 0.027142f
C1340 VDD2.n187 VSUBS 0.027142f
C1341 VDD2.n188 VSUBS 0.014585f
C1342 VDD2.n189 VSUBS 0.015443f
C1343 VDD2.n190 VSUBS 0.034473f
C1344 VDD2.n191 VSUBS 0.07915f
C1345 VDD2.n192 VSUBS 0.015443f
C1346 VDD2.n193 VSUBS 0.014585f
C1347 VDD2.n194 VSUBS 0.060512f
C1348 VDD2.n195 VSUBS 0.058302f
C1349 VDD2.n196 VSUBS 3.23573f
C1350 VDD2.t2 VSUBS 0.374484f
C1351 VDD2.t3 VSUBS 0.374484f
C1352 VDD2.n197 VSUBS 3.09966f
C1353 VTAIL.t9 VSUBS 0.380989f
C1354 VTAIL.t10 VSUBS 0.380989f
C1355 VTAIL.n0 VSUBS 2.96928f
C1356 VTAIL.n1 VSUBS 0.90473f
C1357 VTAIL.n2 VSUBS 0.029055f
C1358 VTAIL.n3 VSUBS 0.027613f
C1359 VTAIL.n4 VSUBS 0.014838f
C1360 VTAIL.n5 VSUBS 0.035072f
C1361 VTAIL.n6 VSUBS 0.015711f
C1362 VTAIL.n7 VSUBS 0.027613f
C1363 VTAIL.n8 VSUBS 0.014838f
C1364 VTAIL.n9 VSUBS 0.035072f
C1365 VTAIL.n10 VSUBS 0.015275f
C1366 VTAIL.n11 VSUBS 0.027613f
C1367 VTAIL.n12 VSUBS 0.015711f
C1368 VTAIL.n13 VSUBS 0.035072f
C1369 VTAIL.n14 VSUBS 0.015711f
C1370 VTAIL.n15 VSUBS 0.027613f
C1371 VTAIL.n16 VSUBS 0.014838f
C1372 VTAIL.n17 VSUBS 0.035072f
C1373 VTAIL.n18 VSUBS 0.015711f
C1374 VTAIL.n19 VSUBS 0.027613f
C1375 VTAIL.n20 VSUBS 0.014838f
C1376 VTAIL.n21 VSUBS 0.035072f
C1377 VTAIL.n22 VSUBS 0.015711f
C1378 VTAIL.n23 VSUBS 0.027613f
C1379 VTAIL.n24 VSUBS 0.014838f
C1380 VTAIL.n25 VSUBS 0.035072f
C1381 VTAIL.n26 VSUBS 0.015711f
C1382 VTAIL.n27 VSUBS 0.027613f
C1383 VTAIL.n28 VSUBS 0.014838f
C1384 VTAIL.n29 VSUBS 0.035072f
C1385 VTAIL.n30 VSUBS 0.015711f
C1386 VTAIL.n31 VSUBS 2.07153f
C1387 VTAIL.n32 VSUBS 0.014838f
C1388 VTAIL.t11 VSUBS 0.075251f
C1389 VTAIL.n33 VSUBS 0.214684f
C1390 VTAIL.n34 VSUBS 0.022311f
C1391 VTAIL.n35 VSUBS 0.026304f
C1392 VTAIL.n36 VSUBS 0.035072f
C1393 VTAIL.n37 VSUBS 0.015711f
C1394 VTAIL.n38 VSUBS 0.014838f
C1395 VTAIL.n39 VSUBS 0.027613f
C1396 VTAIL.n40 VSUBS 0.027613f
C1397 VTAIL.n41 VSUBS 0.014838f
C1398 VTAIL.n42 VSUBS 0.015711f
C1399 VTAIL.n43 VSUBS 0.035072f
C1400 VTAIL.n44 VSUBS 0.035072f
C1401 VTAIL.n45 VSUBS 0.015711f
C1402 VTAIL.n46 VSUBS 0.014838f
C1403 VTAIL.n47 VSUBS 0.027613f
C1404 VTAIL.n48 VSUBS 0.027613f
C1405 VTAIL.n49 VSUBS 0.014838f
C1406 VTAIL.n50 VSUBS 0.015711f
C1407 VTAIL.n51 VSUBS 0.035072f
C1408 VTAIL.n52 VSUBS 0.035072f
C1409 VTAIL.n53 VSUBS 0.015711f
C1410 VTAIL.n54 VSUBS 0.014838f
C1411 VTAIL.n55 VSUBS 0.027613f
C1412 VTAIL.n56 VSUBS 0.027613f
C1413 VTAIL.n57 VSUBS 0.014838f
C1414 VTAIL.n58 VSUBS 0.015711f
C1415 VTAIL.n59 VSUBS 0.035072f
C1416 VTAIL.n60 VSUBS 0.035072f
C1417 VTAIL.n61 VSUBS 0.015711f
C1418 VTAIL.n62 VSUBS 0.014838f
C1419 VTAIL.n63 VSUBS 0.027613f
C1420 VTAIL.n64 VSUBS 0.027613f
C1421 VTAIL.n65 VSUBS 0.014838f
C1422 VTAIL.n66 VSUBS 0.015711f
C1423 VTAIL.n67 VSUBS 0.035072f
C1424 VTAIL.n68 VSUBS 0.035072f
C1425 VTAIL.n69 VSUBS 0.015711f
C1426 VTAIL.n70 VSUBS 0.014838f
C1427 VTAIL.n71 VSUBS 0.027613f
C1428 VTAIL.n72 VSUBS 0.027613f
C1429 VTAIL.n73 VSUBS 0.014838f
C1430 VTAIL.n74 VSUBS 0.014838f
C1431 VTAIL.n75 VSUBS 0.015711f
C1432 VTAIL.n76 VSUBS 0.035072f
C1433 VTAIL.n77 VSUBS 0.035072f
C1434 VTAIL.n78 VSUBS 0.035072f
C1435 VTAIL.n79 VSUBS 0.015275f
C1436 VTAIL.n80 VSUBS 0.014838f
C1437 VTAIL.n81 VSUBS 0.027613f
C1438 VTAIL.n82 VSUBS 0.027613f
C1439 VTAIL.n83 VSUBS 0.014838f
C1440 VTAIL.n84 VSUBS 0.015711f
C1441 VTAIL.n85 VSUBS 0.035072f
C1442 VTAIL.n86 VSUBS 0.035072f
C1443 VTAIL.n87 VSUBS 0.015711f
C1444 VTAIL.n88 VSUBS 0.014838f
C1445 VTAIL.n89 VSUBS 0.027613f
C1446 VTAIL.n90 VSUBS 0.027613f
C1447 VTAIL.n91 VSUBS 0.014838f
C1448 VTAIL.n92 VSUBS 0.015711f
C1449 VTAIL.n93 VSUBS 0.035072f
C1450 VTAIL.n94 VSUBS 0.080525f
C1451 VTAIL.n95 VSUBS 0.015711f
C1452 VTAIL.n96 VSUBS 0.014838f
C1453 VTAIL.n97 VSUBS 0.061563f
C1454 VTAIL.n98 VSUBS 0.04023f
C1455 VTAIL.n99 VSUBS 0.402371f
C1456 VTAIL.t1 VSUBS 0.380989f
C1457 VTAIL.t2 VSUBS 0.380989f
C1458 VTAIL.n100 VSUBS 2.96928f
C1459 VTAIL.n101 VSUBS 3.07947f
C1460 VTAIL.t8 VSUBS 0.380989f
C1461 VTAIL.t5 VSUBS 0.380989f
C1462 VTAIL.n102 VSUBS 2.9693f
C1463 VTAIL.n103 VSUBS 3.07945f
C1464 VTAIL.n104 VSUBS 0.029055f
C1465 VTAIL.n105 VSUBS 0.027613f
C1466 VTAIL.n106 VSUBS 0.014838f
C1467 VTAIL.n107 VSUBS 0.035072f
C1468 VTAIL.n108 VSUBS 0.015711f
C1469 VTAIL.n109 VSUBS 0.027613f
C1470 VTAIL.n110 VSUBS 0.014838f
C1471 VTAIL.n111 VSUBS 0.035072f
C1472 VTAIL.n112 VSUBS 0.015275f
C1473 VTAIL.n113 VSUBS 0.027613f
C1474 VTAIL.n114 VSUBS 0.015275f
C1475 VTAIL.n115 VSUBS 0.014838f
C1476 VTAIL.n116 VSUBS 0.035072f
C1477 VTAIL.n117 VSUBS 0.035072f
C1478 VTAIL.n118 VSUBS 0.015711f
C1479 VTAIL.n119 VSUBS 0.027613f
C1480 VTAIL.n120 VSUBS 0.014838f
C1481 VTAIL.n121 VSUBS 0.035072f
C1482 VTAIL.n122 VSUBS 0.015711f
C1483 VTAIL.n123 VSUBS 0.027613f
C1484 VTAIL.n124 VSUBS 0.014838f
C1485 VTAIL.n125 VSUBS 0.035072f
C1486 VTAIL.n126 VSUBS 0.015711f
C1487 VTAIL.n127 VSUBS 0.027613f
C1488 VTAIL.n128 VSUBS 0.014838f
C1489 VTAIL.n129 VSUBS 0.035072f
C1490 VTAIL.n130 VSUBS 0.015711f
C1491 VTAIL.n131 VSUBS 0.027613f
C1492 VTAIL.n132 VSUBS 0.014838f
C1493 VTAIL.n133 VSUBS 0.035072f
C1494 VTAIL.n134 VSUBS 0.015711f
C1495 VTAIL.n135 VSUBS 2.07153f
C1496 VTAIL.n136 VSUBS 0.014838f
C1497 VTAIL.t7 VSUBS 0.075251f
C1498 VTAIL.n137 VSUBS 0.214684f
C1499 VTAIL.n138 VSUBS 0.022311f
C1500 VTAIL.n139 VSUBS 0.026304f
C1501 VTAIL.n140 VSUBS 0.035072f
C1502 VTAIL.n141 VSUBS 0.015711f
C1503 VTAIL.n142 VSUBS 0.014838f
C1504 VTAIL.n143 VSUBS 0.027613f
C1505 VTAIL.n144 VSUBS 0.027613f
C1506 VTAIL.n145 VSUBS 0.014838f
C1507 VTAIL.n146 VSUBS 0.015711f
C1508 VTAIL.n147 VSUBS 0.035072f
C1509 VTAIL.n148 VSUBS 0.035072f
C1510 VTAIL.n149 VSUBS 0.015711f
C1511 VTAIL.n150 VSUBS 0.014838f
C1512 VTAIL.n151 VSUBS 0.027613f
C1513 VTAIL.n152 VSUBS 0.027613f
C1514 VTAIL.n153 VSUBS 0.014838f
C1515 VTAIL.n154 VSUBS 0.015711f
C1516 VTAIL.n155 VSUBS 0.035072f
C1517 VTAIL.n156 VSUBS 0.035072f
C1518 VTAIL.n157 VSUBS 0.015711f
C1519 VTAIL.n158 VSUBS 0.014838f
C1520 VTAIL.n159 VSUBS 0.027613f
C1521 VTAIL.n160 VSUBS 0.027613f
C1522 VTAIL.n161 VSUBS 0.014838f
C1523 VTAIL.n162 VSUBS 0.015711f
C1524 VTAIL.n163 VSUBS 0.035072f
C1525 VTAIL.n164 VSUBS 0.035072f
C1526 VTAIL.n165 VSUBS 0.015711f
C1527 VTAIL.n166 VSUBS 0.014838f
C1528 VTAIL.n167 VSUBS 0.027613f
C1529 VTAIL.n168 VSUBS 0.027613f
C1530 VTAIL.n169 VSUBS 0.014838f
C1531 VTAIL.n170 VSUBS 0.015711f
C1532 VTAIL.n171 VSUBS 0.035072f
C1533 VTAIL.n172 VSUBS 0.035072f
C1534 VTAIL.n173 VSUBS 0.015711f
C1535 VTAIL.n174 VSUBS 0.014838f
C1536 VTAIL.n175 VSUBS 0.027613f
C1537 VTAIL.n176 VSUBS 0.027613f
C1538 VTAIL.n177 VSUBS 0.014838f
C1539 VTAIL.n178 VSUBS 0.015711f
C1540 VTAIL.n179 VSUBS 0.035072f
C1541 VTAIL.n180 VSUBS 0.035072f
C1542 VTAIL.n181 VSUBS 0.015711f
C1543 VTAIL.n182 VSUBS 0.014838f
C1544 VTAIL.n183 VSUBS 0.027613f
C1545 VTAIL.n184 VSUBS 0.027613f
C1546 VTAIL.n185 VSUBS 0.014838f
C1547 VTAIL.n186 VSUBS 0.015711f
C1548 VTAIL.n187 VSUBS 0.035072f
C1549 VTAIL.n188 VSUBS 0.035072f
C1550 VTAIL.n189 VSUBS 0.015711f
C1551 VTAIL.n190 VSUBS 0.014838f
C1552 VTAIL.n191 VSUBS 0.027613f
C1553 VTAIL.n192 VSUBS 0.027613f
C1554 VTAIL.n193 VSUBS 0.014838f
C1555 VTAIL.n194 VSUBS 0.015711f
C1556 VTAIL.n195 VSUBS 0.035072f
C1557 VTAIL.n196 VSUBS 0.080525f
C1558 VTAIL.n197 VSUBS 0.015711f
C1559 VTAIL.n198 VSUBS 0.014838f
C1560 VTAIL.n199 VSUBS 0.061563f
C1561 VTAIL.n200 VSUBS 0.04023f
C1562 VTAIL.n201 VSUBS 0.402371f
C1563 VTAIL.t0 VSUBS 0.380989f
C1564 VTAIL.t4 VSUBS 0.380989f
C1565 VTAIL.n202 VSUBS 2.9693f
C1566 VTAIL.n203 VSUBS 1.06866f
C1567 VTAIL.n204 VSUBS 0.029055f
C1568 VTAIL.n205 VSUBS 0.027613f
C1569 VTAIL.n206 VSUBS 0.014838f
C1570 VTAIL.n207 VSUBS 0.035072f
C1571 VTAIL.n208 VSUBS 0.015711f
C1572 VTAIL.n209 VSUBS 0.027613f
C1573 VTAIL.n210 VSUBS 0.014838f
C1574 VTAIL.n211 VSUBS 0.035072f
C1575 VTAIL.n212 VSUBS 0.015275f
C1576 VTAIL.n213 VSUBS 0.027613f
C1577 VTAIL.n214 VSUBS 0.015275f
C1578 VTAIL.n215 VSUBS 0.014838f
C1579 VTAIL.n216 VSUBS 0.035072f
C1580 VTAIL.n217 VSUBS 0.035072f
C1581 VTAIL.n218 VSUBS 0.015711f
C1582 VTAIL.n219 VSUBS 0.027613f
C1583 VTAIL.n220 VSUBS 0.014838f
C1584 VTAIL.n221 VSUBS 0.035072f
C1585 VTAIL.n222 VSUBS 0.015711f
C1586 VTAIL.n223 VSUBS 0.027613f
C1587 VTAIL.n224 VSUBS 0.014838f
C1588 VTAIL.n225 VSUBS 0.035072f
C1589 VTAIL.n226 VSUBS 0.015711f
C1590 VTAIL.n227 VSUBS 0.027613f
C1591 VTAIL.n228 VSUBS 0.014838f
C1592 VTAIL.n229 VSUBS 0.035072f
C1593 VTAIL.n230 VSUBS 0.015711f
C1594 VTAIL.n231 VSUBS 0.027613f
C1595 VTAIL.n232 VSUBS 0.014838f
C1596 VTAIL.n233 VSUBS 0.035072f
C1597 VTAIL.n234 VSUBS 0.015711f
C1598 VTAIL.n235 VSUBS 2.07153f
C1599 VTAIL.n236 VSUBS 0.014838f
C1600 VTAIL.t3 VSUBS 0.075251f
C1601 VTAIL.n237 VSUBS 0.214684f
C1602 VTAIL.n238 VSUBS 0.022311f
C1603 VTAIL.n239 VSUBS 0.026304f
C1604 VTAIL.n240 VSUBS 0.035072f
C1605 VTAIL.n241 VSUBS 0.015711f
C1606 VTAIL.n242 VSUBS 0.014838f
C1607 VTAIL.n243 VSUBS 0.027613f
C1608 VTAIL.n244 VSUBS 0.027613f
C1609 VTAIL.n245 VSUBS 0.014838f
C1610 VTAIL.n246 VSUBS 0.015711f
C1611 VTAIL.n247 VSUBS 0.035072f
C1612 VTAIL.n248 VSUBS 0.035072f
C1613 VTAIL.n249 VSUBS 0.015711f
C1614 VTAIL.n250 VSUBS 0.014838f
C1615 VTAIL.n251 VSUBS 0.027613f
C1616 VTAIL.n252 VSUBS 0.027613f
C1617 VTAIL.n253 VSUBS 0.014838f
C1618 VTAIL.n254 VSUBS 0.015711f
C1619 VTAIL.n255 VSUBS 0.035072f
C1620 VTAIL.n256 VSUBS 0.035072f
C1621 VTAIL.n257 VSUBS 0.015711f
C1622 VTAIL.n258 VSUBS 0.014838f
C1623 VTAIL.n259 VSUBS 0.027613f
C1624 VTAIL.n260 VSUBS 0.027613f
C1625 VTAIL.n261 VSUBS 0.014838f
C1626 VTAIL.n262 VSUBS 0.015711f
C1627 VTAIL.n263 VSUBS 0.035072f
C1628 VTAIL.n264 VSUBS 0.035072f
C1629 VTAIL.n265 VSUBS 0.015711f
C1630 VTAIL.n266 VSUBS 0.014838f
C1631 VTAIL.n267 VSUBS 0.027613f
C1632 VTAIL.n268 VSUBS 0.027613f
C1633 VTAIL.n269 VSUBS 0.014838f
C1634 VTAIL.n270 VSUBS 0.015711f
C1635 VTAIL.n271 VSUBS 0.035072f
C1636 VTAIL.n272 VSUBS 0.035072f
C1637 VTAIL.n273 VSUBS 0.015711f
C1638 VTAIL.n274 VSUBS 0.014838f
C1639 VTAIL.n275 VSUBS 0.027613f
C1640 VTAIL.n276 VSUBS 0.027613f
C1641 VTAIL.n277 VSUBS 0.014838f
C1642 VTAIL.n278 VSUBS 0.015711f
C1643 VTAIL.n279 VSUBS 0.035072f
C1644 VTAIL.n280 VSUBS 0.035072f
C1645 VTAIL.n281 VSUBS 0.015711f
C1646 VTAIL.n282 VSUBS 0.014838f
C1647 VTAIL.n283 VSUBS 0.027613f
C1648 VTAIL.n284 VSUBS 0.027613f
C1649 VTAIL.n285 VSUBS 0.014838f
C1650 VTAIL.n286 VSUBS 0.015711f
C1651 VTAIL.n287 VSUBS 0.035072f
C1652 VTAIL.n288 VSUBS 0.035072f
C1653 VTAIL.n289 VSUBS 0.015711f
C1654 VTAIL.n290 VSUBS 0.014838f
C1655 VTAIL.n291 VSUBS 0.027613f
C1656 VTAIL.n292 VSUBS 0.027613f
C1657 VTAIL.n293 VSUBS 0.014838f
C1658 VTAIL.n294 VSUBS 0.015711f
C1659 VTAIL.n295 VSUBS 0.035072f
C1660 VTAIL.n296 VSUBS 0.080525f
C1661 VTAIL.n297 VSUBS 0.015711f
C1662 VTAIL.n298 VSUBS 0.014838f
C1663 VTAIL.n299 VSUBS 0.061563f
C1664 VTAIL.n300 VSUBS 0.04023f
C1665 VTAIL.n301 VSUBS 2.18765f
C1666 VTAIL.n302 VSUBS 0.029055f
C1667 VTAIL.n303 VSUBS 0.027613f
C1668 VTAIL.n304 VSUBS 0.014838f
C1669 VTAIL.n305 VSUBS 0.035072f
C1670 VTAIL.n306 VSUBS 0.015711f
C1671 VTAIL.n307 VSUBS 0.027613f
C1672 VTAIL.n308 VSUBS 0.014838f
C1673 VTAIL.n309 VSUBS 0.035072f
C1674 VTAIL.n310 VSUBS 0.015275f
C1675 VTAIL.n311 VSUBS 0.027613f
C1676 VTAIL.n312 VSUBS 0.015711f
C1677 VTAIL.n313 VSUBS 0.035072f
C1678 VTAIL.n314 VSUBS 0.015711f
C1679 VTAIL.n315 VSUBS 0.027613f
C1680 VTAIL.n316 VSUBS 0.014838f
C1681 VTAIL.n317 VSUBS 0.035072f
C1682 VTAIL.n318 VSUBS 0.015711f
C1683 VTAIL.n319 VSUBS 0.027613f
C1684 VTAIL.n320 VSUBS 0.014838f
C1685 VTAIL.n321 VSUBS 0.035072f
C1686 VTAIL.n322 VSUBS 0.015711f
C1687 VTAIL.n323 VSUBS 0.027613f
C1688 VTAIL.n324 VSUBS 0.014838f
C1689 VTAIL.n325 VSUBS 0.035072f
C1690 VTAIL.n326 VSUBS 0.015711f
C1691 VTAIL.n327 VSUBS 0.027613f
C1692 VTAIL.n328 VSUBS 0.014838f
C1693 VTAIL.n329 VSUBS 0.035072f
C1694 VTAIL.n330 VSUBS 0.015711f
C1695 VTAIL.n331 VSUBS 2.07153f
C1696 VTAIL.n332 VSUBS 0.014838f
C1697 VTAIL.t6 VSUBS 0.075251f
C1698 VTAIL.n333 VSUBS 0.214684f
C1699 VTAIL.n334 VSUBS 0.022311f
C1700 VTAIL.n335 VSUBS 0.026304f
C1701 VTAIL.n336 VSUBS 0.035072f
C1702 VTAIL.n337 VSUBS 0.015711f
C1703 VTAIL.n338 VSUBS 0.014838f
C1704 VTAIL.n339 VSUBS 0.027613f
C1705 VTAIL.n340 VSUBS 0.027613f
C1706 VTAIL.n341 VSUBS 0.014838f
C1707 VTAIL.n342 VSUBS 0.015711f
C1708 VTAIL.n343 VSUBS 0.035072f
C1709 VTAIL.n344 VSUBS 0.035072f
C1710 VTAIL.n345 VSUBS 0.015711f
C1711 VTAIL.n346 VSUBS 0.014838f
C1712 VTAIL.n347 VSUBS 0.027613f
C1713 VTAIL.n348 VSUBS 0.027613f
C1714 VTAIL.n349 VSUBS 0.014838f
C1715 VTAIL.n350 VSUBS 0.015711f
C1716 VTAIL.n351 VSUBS 0.035072f
C1717 VTAIL.n352 VSUBS 0.035072f
C1718 VTAIL.n353 VSUBS 0.015711f
C1719 VTAIL.n354 VSUBS 0.014838f
C1720 VTAIL.n355 VSUBS 0.027613f
C1721 VTAIL.n356 VSUBS 0.027613f
C1722 VTAIL.n357 VSUBS 0.014838f
C1723 VTAIL.n358 VSUBS 0.015711f
C1724 VTAIL.n359 VSUBS 0.035072f
C1725 VTAIL.n360 VSUBS 0.035072f
C1726 VTAIL.n361 VSUBS 0.015711f
C1727 VTAIL.n362 VSUBS 0.014838f
C1728 VTAIL.n363 VSUBS 0.027613f
C1729 VTAIL.n364 VSUBS 0.027613f
C1730 VTAIL.n365 VSUBS 0.014838f
C1731 VTAIL.n366 VSUBS 0.015711f
C1732 VTAIL.n367 VSUBS 0.035072f
C1733 VTAIL.n368 VSUBS 0.035072f
C1734 VTAIL.n369 VSUBS 0.015711f
C1735 VTAIL.n370 VSUBS 0.014838f
C1736 VTAIL.n371 VSUBS 0.027613f
C1737 VTAIL.n372 VSUBS 0.027613f
C1738 VTAIL.n373 VSUBS 0.014838f
C1739 VTAIL.n374 VSUBS 0.014838f
C1740 VTAIL.n375 VSUBS 0.015711f
C1741 VTAIL.n376 VSUBS 0.035072f
C1742 VTAIL.n377 VSUBS 0.035072f
C1743 VTAIL.n378 VSUBS 0.035072f
C1744 VTAIL.n379 VSUBS 0.015275f
C1745 VTAIL.n380 VSUBS 0.014838f
C1746 VTAIL.n381 VSUBS 0.027613f
C1747 VTAIL.n382 VSUBS 0.027613f
C1748 VTAIL.n383 VSUBS 0.014838f
C1749 VTAIL.n384 VSUBS 0.015711f
C1750 VTAIL.n385 VSUBS 0.035072f
C1751 VTAIL.n386 VSUBS 0.035072f
C1752 VTAIL.n387 VSUBS 0.015711f
C1753 VTAIL.n388 VSUBS 0.014838f
C1754 VTAIL.n389 VSUBS 0.027613f
C1755 VTAIL.n390 VSUBS 0.027613f
C1756 VTAIL.n391 VSUBS 0.014838f
C1757 VTAIL.n392 VSUBS 0.015711f
C1758 VTAIL.n393 VSUBS 0.035072f
C1759 VTAIL.n394 VSUBS 0.080525f
C1760 VTAIL.n395 VSUBS 0.015711f
C1761 VTAIL.n396 VSUBS 0.014838f
C1762 VTAIL.n397 VSUBS 0.061563f
C1763 VTAIL.n398 VSUBS 0.04023f
C1764 VTAIL.n399 VSUBS 2.12609f
C1765 VN.n0 VSUBS 0.036184f
C1766 VN.t5 VSUBS 3.43833f
C1767 VN.n1 VSUBS 0.042176f
C1768 VN.n2 VSUBS 0.027447f
C1769 VN.t1 VSUBS 3.43833f
C1770 VN.n3 VSUBS 1.27233f
C1771 VN.t0 VSUBS 3.67274f
C1772 VN.n4 VSUBS 1.24225f
C1773 VN.n5 VSUBS 0.26553f
C1774 VN.n6 VSUBS 0.038334f
C1775 VN.n7 VSUBS 0.050898f
C1776 VN.n8 VSUBS 0.03762f
C1777 VN.n9 VSUBS 0.027447f
C1778 VN.n10 VSUBS 0.027447f
C1779 VN.n11 VSUBS 0.027447f
C1780 VN.n12 VSUBS 0.050898f
C1781 VN.n13 VSUBS 0.035319f
C1782 VN.n14 VSUBS 1.28438f
C1783 VN.n15 VSUBS 0.045204f
C1784 VN.n16 VSUBS 0.036184f
C1785 VN.t4 VSUBS 3.43833f
C1786 VN.n17 VSUBS 0.042176f
C1787 VN.n18 VSUBS 0.027447f
C1788 VN.t3 VSUBS 3.43833f
C1789 VN.n19 VSUBS 1.27233f
C1790 VN.t2 VSUBS 3.67274f
C1791 VN.n20 VSUBS 1.24225f
C1792 VN.n21 VSUBS 0.26553f
C1793 VN.n22 VSUBS 0.038334f
C1794 VN.n23 VSUBS 0.050898f
C1795 VN.n24 VSUBS 0.03762f
C1796 VN.n25 VSUBS 0.027447f
C1797 VN.n26 VSUBS 0.027447f
C1798 VN.n27 VSUBS 0.027447f
C1799 VN.n28 VSUBS 0.050898f
C1800 VN.n29 VSUBS 0.035319f
C1801 VN.n30 VSUBS 1.28438f
C1802 VN.n31 VSUBS 1.67089f
.ends

