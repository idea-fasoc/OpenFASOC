* NGSPICE file created from diff_pair_sample_1656.ext - technology: sky130A

.subckt diff_pair_sample_1656 VTAIL VN VP B VDD2 VDD1
X0 B.t13 B.t11 B.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=0 ps=0 w=10.05 l=3.87
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t14 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=3.9195 ps=20.88 w=10.05 l=3.87
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t15 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=3.9195 ps=20.88 w=10.05 l=3.87
X3 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=0 ps=0 w=10.05 l=3.87
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t14 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=3.9195 ps=20.88 w=10.05 l=3.87
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t15 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=3.9195 ps=20.88 w=10.05 l=3.87
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=0 ps=0 w=10.05 l=3.87
X7 B.t3 B.t0 B.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.9195 pd=20.88 as=0 ps=0 w=10.05 l=3.87
R0 B.n683 B.n682 585
R1 B.n684 B.n683 585
R2 B.n268 B.n103 585
R3 B.n267 B.n266 585
R4 B.n265 B.n264 585
R5 B.n263 B.n262 585
R6 B.n261 B.n260 585
R7 B.n259 B.n258 585
R8 B.n257 B.n256 585
R9 B.n255 B.n254 585
R10 B.n253 B.n252 585
R11 B.n251 B.n250 585
R12 B.n249 B.n248 585
R13 B.n247 B.n246 585
R14 B.n245 B.n244 585
R15 B.n243 B.n242 585
R16 B.n241 B.n240 585
R17 B.n239 B.n238 585
R18 B.n237 B.n236 585
R19 B.n235 B.n234 585
R20 B.n233 B.n232 585
R21 B.n231 B.n230 585
R22 B.n229 B.n228 585
R23 B.n227 B.n226 585
R24 B.n225 B.n224 585
R25 B.n223 B.n222 585
R26 B.n221 B.n220 585
R27 B.n219 B.n218 585
R28 B.n217 B.n216 585
R29 B.n215 B.n214 585
R30 B.n213 B.n212 585
R31 B.n211 B.n210 585
R32 B.n209 B.n208 585
R33 B.n207 B.n206 585
R34 B.n205 B.n204 585
R35 B.n203 B.n202 585
R36 B.n201 B.n200 585
R37 B.n198 B.n197 585
R38 B.n196 B.n195 585
R39 B.n194 B.n193 585
R40 B.n192 B.n191 585
R41 B.n190 B.n189 585
R42 B.n188 B.n187 585
R43 B.n186 B.n185 585
R44 B.n184 B.n183 585
R45 B.n182 B.n181 585
R46 B.n180 B.n179 585
R47 B.n178 B.n177 585
R48 B.n176 B.n175 585
R49 B.n174 B.n173 585
R50 B.n172 B.n171 585
R51 B.n170 B.n169 585
R52 B.n168 B.n167 585
R53 B.n166 B.n165 585
R54 B.n164 B.n163 585
R55 B.n162 B.n161 585
R56 B.n160 B.n159 585
R57 B.n158 B.n157 585
R58 B.n156 B.n155 585
R59 B.n154 B.n153 585
R60 B.n152 B.n151 585
R61 B.n150 B.n149 585
R62 B.n148 B.n147 585
R63 B.n146 B.n145 585
R64 B.n144 B.n143 585
R65 B.n142 B.n141 585
R66 B.n140 B.n139 585
R67 B.n138 B.n137 585
R68 B.n136 B.n135 585
R69 B.n134 B.n133 585
R70 B.n132 B.n131 585
R71 B.n130 B.n129 585
R72 B.n128 B.n127 585
R73 B.n126 B.n125 585
R74 B.n124 B.n123 585
R75 B.n122 B.n121 585
R76 B.n120 B.n119 585
R77 B.n118 B.n117 585
R78 B.n116 B.n115 585
R79 B.n114 B.n113 585
R80 B.n112 B.n111 585
R81 B.n110 B.n109 585
R82 B.n681 B.n62 585
R83 B.n685 B.n62 585
R84 B.n680 B.n61 585
R85 B.n686 B.n61 585
R86 B.n679 B.n678 585
R87 B.n678 B.n57 585
R88 B.n677 B.n56 585
R89 B.n692 B.n56 585
R90 B.n676 B.n55 585
R91 B.n693 B.n55 585
R92 B.n675 B.n54 585
R93 B.n694 B.n54 585
R94 B.n674 B.n673 585
R95 B.n673 B.n50 585
R96 B.n672 B.n49 585
R97 B.n700 B.n49 585
R98 B.n671 B.n48 585
R99 B.n701 B.n48 585
R100 B.n670 B.n47 585
R101 B.n702 B.n47 585
R102 B.n669 B.n668 585
R103 B.n668 B.n43 585
R104 B.n667 B.n42 585
R105 B.n708 B.n42 585
R106 B.n666 B.n41 585
R107 B.n709 B.n41 585
R108 B.n665 B.n40 585
R109 B.n710 B.n40 585
R110 B.n664 B.n663 585
R111 B.n663 B.n36 585
R112 B.n662 B.n35 585
R113 B.n716 B.n35 585
R114 B.n661 B.n34 585
R115 B.n717 B.n34 585
R116 B.n660 B.n33 585
R117 B.n718 B.n33 585
R118 B.n659 B.n658 585
R119 B.n658 B.n29 585
R120 B.n657 B.n28 585
R121 B.n724 B.n28 585
R122 B.n656 B.n27 585
R123 B.n725 B.n27 585
R124 B.n655 B.n26 585
R125 B.n726 B.n26 585
R126 B.n654 B.n653 585
R127 B.n653 B.n22 585
R128 B.n652 B.n21 585
R129 B.n732 B.n21 585
R130 B.n651 B.n20 585
R131 B.n733 B.n20 585
R132 B.n650 B.n19 585
R133 B.n734 B.n19 585
R134 B.n649 B.n648 585
R135 B.n648 B.n15 585
R136 B.n647 B.n14 585
R137 B.n740 B.n14 585
R138 B.n646 B.n13 585
R139 B.n741 B.n13 585
R140 B.n645 B.n12 585
R141 B.n742 B.n12 585
R142 B.n644 B.n643 585
R143 B.n643 B.n8 585
R144 B.n642 B.n7 585
R145 B.n748 B.n7 585
R146 B.n641 B.n6 585
R147 B.n749 B.n6 585
R148 B.n640 B.n5 585
R149 B.n750 B.n5 585
R150 B.n639 B.n638 585
R151 B.n638 B.n4 585
R152 B.n637 B.n269 585
R153 B.n637 B.n636 585
R154 B.n627 B.n270 585
R155 B.n271 B.n270 585
R156 B.n629 B.n628 585
R157 B.n630 B.n629 585
R158 B.n626 B.n276 585
R159 B.n276 B.n275 585
R160 B.n625 B.n624 585
R161 B.n624 B.n623 585
R162 B.n278 B.n277 585
R163 B.n279 B.n278 585
R164 B.n616 B.n615 585
R165 B.n617 B.n616 585
R166 B.n614 B.n284 585
R167 B.n284 B.n283 585
R168 B.n613 B.n612 585
R169 B.n612 B.n611 585
R170 B.n286 B.n285 585
R171 B.n287 B.n286 585
R172 B.n604 B.n603 585
R173 B.n605 B.n604 585
R174 B.n602 B.n292 585
R175 B.n292 B.n291 585
R176 B.n601 B.n600 585
R177 B.n600 B.n599 585
R178 B.n294 B.n293 585
R179 B.n295 B.n294 585
R180 B.n592 B.n591 585
R181 B.n593 B.n592 585
R182 B.n590 B.n300 585
R183 B.n300 B.n299 585
R184 B.n589 B.n588 585
R185 B.n588 B.n587 585
R186 B.n302 B.n301 585
R187 B.n303 B.n302 585
R188 B.n580 B.n579 585
R189 B.n581 B.n580 585
R190 B.n578 B.n308 585
R191 B.n308 B.n307 585
R192 B.n577 B.n576 585
R193 B.n576 B.n575 585
R194 B.n310 B.n309 585
R195 B.n311 B.n310 585
R196 B.n568 B.n567 585
R197 B.n569 B.n568 585
R198 B.n566 B.n316 585
R199 B.n316 B.n315 585
R200 B.n565 B.n564 585
R201 B.n564 B.n563 585
R202 B.n318 B.n317 585
R203 B.n319 B.n318 585
R204 B.n556 B.n555 585
R205 B.n557 B.n556 585
R206 B.n554 B.n324 585
R207 B.n324 B.n323 585
R208 B.n553 B.n552 585
R209 B.n552 B.n551 585
R210 B.n326 B.n325 585
R211 B.n327 B.n326 585
R212 B.n544 B.n543 585
R213 B.n545 B.n544 585
R214 B.n542 B.n332 585
R215 B.n332 B.n331 585
R216 B.n536 B.n535 585
R217 B.n534 B.n374 585
R218 B.n533 B.n373 585
R219 B.n538 B.n373 585
R220 B.n532 B.n531 585
R221 B.n530 B.n529 585
R222 B.n528 B.n527 585
R223 B.n526 B.n525 585
R224 B.n524 B.n523 585
R225 B.n522 B.n521 585
R226 B.n520 B.n519 585
R227 B.n518 B.n517 585
R228 B.n516 B.n515 585
R229 B.n514 B.n513 585
R230 B.n512 B.n511 585
R231 B.n510 B.n509 585
R232 B.n508 B.n507 585
R233 B.n506 B.n505 585
R234 B.n504 B.n503 585
R235 B.n502 B.n501 585
R236 B.n500 B.n499 585
R237 B.n498 B.n497 585
R238 B.n496 B.n495 585
R239 B.n494 B.n493 585
R240 B.n492 B.n491 585
R241 B.n490 B.n489 585
R242 B.n488 B.n487 585
R243 B.n486 B.n485 585
R244 B.n484 B.n483 585
R245 B.n482 B.n481 585
R246 B.n480 B.n479 585
R247 B.n478 B.n477 585
R248 B.n476 B.n475 585
R249 B.n474 B.n473 585
R250 B.n472 B.n471 585
R251 B.n470 B.n469 585
R252 B.n468 B.n467 585
R253 B.n465 B.n464 585
R254 B.n463 B.n462 585
R255 B.n461 B.n460 585
R256 B.n459 B.n458 585
R257 B.n457 B.n456 585
R258 B.n455 B.n454 585
R259 B.n453 B.n452 585
R260 B.n451 B.n450 585
R261 B.n449 B.n448 585
R262 B.n447 B.n446 585
R263 B.n445 B.n444 585
R264 B.n443 B.n442 585
R265 B.n441 B.n440 585
R266 B.n439 B.n438 585
R267 B.n437 B.n436 585
R268 B.n435 B.n434 585
R269 B.n433 B.n432 585
R270 B.n431 B.n430 585
R271 B.n429 B.n428 585
R272 B.n427 B.n426 585
R273 B.n425 B.n424 585
R274 B.n423 B.n422 585
R275 B.n421 B.n420 585
R276 B.n419 B.n418 585
R277 B.n417 B.n416 585
R278 B.n415 B.n414 585
R279 B.n413 B.n412 585
R280 B.n411 B.n410 585
R281 B.n409 B.n408 585
R282 B.n407 B.n406 585
R283 B.n405 B.n404 585
R284 B.n403 B.n402 585
R285 B.n401 B.n400 585
R286 B.n399 B.n398 585
R287 B.n397 B.n396 585
R288 B.n395 B.n394 585
R289 B.n393 B.n392 585
R290 B.n391 B.n390 585
R291 B.n389 B.n388 585
R292 B.n387 B.n386 585
R293 B.n385 B.n384 585
R294 B.n383 B.n382 585
R295 B.n381 B.n380 585
R296 B.n334 B.n333 585
R297 B.n541 B.n540 585
R298 B.n330 B.n329 585
R299 B.n331 B.n330 585
R300 B.n547 B.n546 585
R301 B.n546 B.n545 585
R302 B.n548 B.n328 585
R303 B.n328 B.n327 585
R304 B.n550 B.n549 585
R305 B.n551 B.n550 585
R306 B.n322 B.n321 585
R307 B.n323 B.n322 585
R308 B.n559 B.n558 585
R309 B.n558 B.n557 585
R310 B.n560 B.n320 585
R311 B.n320 B.n319 585
R312 B.n562 B.n561 585
R313 B.n563 B.n562 585
R314 B.n314 B.n313 585
R315 B.n315 B.n314 585
R316 B.n571 B.n570 585
R317 B.n570 B.n569 585
R318 B.n572 B.n312 585
R319 B.n312 B.n311 585
R320 B.n574 B.n573 585
R321 B.n575 B.n574 585
R322 B.n306 B.n305 585
R323 B.n307 B.n306 585
R324 B.n583 B.n582 585
R325 B.n582 B.n581 585
R326 B.n584 B.n304 585
R327 B.n304 B.n303 585
R328 B.n586 B.n585 585
R329 B.n587 B.n586 585
R330 B.n298 B.n297 585
R331 B.n299 B.n298 585
R332 B.n595 B.n594 585
R333 B.n594 B.n593 585
R334 B.n596 B.n296 585
R335 B.n296 B.n295 585
R336 B.n598 B.n597 585
R337 B.n599 B.n598 585
R338 B.n290 B.n289 585
R339 B.n291 B.n290 585
R340 B.n607 B.n606 585
R341 B.n606 B.n605 585
R342 B.n608 B.n288 585
R343 B.n288 B.n287 585
R344 B.n610 B.n609 585
R345 B.n611 B.n610 585
R346 B.n282 B.n281 585
R347 B.n283 B.n282 585
R348 B.n619 B.n618 585
R349 B.n618 B.n617 585
R350 B.n620 B.n280 585
R351 B.n280 B.n279 585
R352 B.n622 B.n621 585
R353 B.n623 B.n622 585
R354 B.n274 B.n273 585
R355 B.n275 B.n274 585
R356 B.n632 B.n631 585
R357 B.n631 B.n630 585
R358 B.n633 B.n272 585
R359 B.n272 B.n271 585
R360 B.n635 B.n634 585
R361 B.n636 B.n635 585
R362 B.n2 B.n0 585
R363 B.n4 B.n2 585
R364 B.n3 B.n1 585
R365 B.n749 B.n3 585
R366 B.n747 B.n746 585
R367 B.n748 B.n747 585
R368 B.n745 B.n9 585
R369 B.n9 B.n8 585
R370 B.n744 B.n743 585
R371 B.n743 B.n742 585
R372 B.n11 B.n10 585
R373 B.n741 B.n11 585
R374 B.n739 B.n738 585
R375 B.n740 B.n739 585
R376 B.n737 B.n16 585
R377 B.n16 B.n15 585
R378 B.n736 B.n735 585
R379 B.n735 B.n734 585
R380 B.n18 B.n17 585
R381 B.n733 B.n18 585
R382 B.n731 B.n730 585
R383 B.n732 B.n731 585
R384 B.n729 B.n23 585
R385 B.n23 B.n22 585
R386 B.n728 B.n727 585
R387 B.n727 B.n726 585
R388 B.n25 B.n24 585
R389 B.n725 B.n25 585
R390 B.n723 B.n722 585
R391 B.n724 B.n723 585
R392 B.n721 B.n30 585
R393 B.n30 B.n29 585
R394 B.n720 B.n719 585
R395 B.n719 B.n718 585
R396 B.n32 B.n31 585
R397 B.n717 B.n32 585
R398 B.n715 B.n714 585
R399 B.n716 B.n715 585
R400 B.n713 B.n37 585
R401 B.n37 B.n36 585
R402 B.n712 B.n711 585
R403 B.n711 B.n710 585
R404 B.n39 B.n38 585
R405 B.n709 B.n39 585
R406 B.n707 B.n706 585
R407 B.n708 B.n707 585
R408 B.n705 B.n44 585
R409 B.n44 B.n43 585
R410 B.n704 B.n703 585
R411 B.n703 B.n702 585
R412 B.n46 B.n45 585
R413 B.n701 B.n46 585
R414 B.n699 B.n698 585
R415 B.n700 B.n699 585
R416 B.n697 B.n51 585
R417 B.n51 B.n50 585
R418 B.n696 B.n695 585
R419 B.n695 B.n694 585
R420 B.n53 B.n52 585
R421 B.n693 B.n53 585
R422 B.n691 B.n690 585
R423 B.n692 B.n691 585
R424 B.n689 B.n58 585
R425 B.n58 B.n57 585
R426 B.n688 B.n687 585
R427 B.n687 B.n686 585
R428 B.n60 B.n59 585
R429 B.n685 B.n60 585
R430 B.n752 B.n751 585
R431 B.n751 B.n750 585
R432 B.n536 B.n330 497.305
R433 B.n109 B.n60 497.305
R434 B.n540 B.n332 497.305
R435 B.n683 B.n62 497.305
R436 B.n377 B.t3 330.072
R437 B.n104 B.t6 330.072
R438 B.n375 B.t13 330.072
R439 B.n106 B.t9 330.072
R440 B.n377 B.t0 271.983
R441 B.n375 B.t11 271.983
R442 B.n106 B.t8 271.983
R443 B.n104 B.t4 271.983
R444 B.n684 B.n102 256.663
R445 B.n684 B.n101 256.663
R446 B.n684 B.n100 256.663
R447 B.n684 B.n99 256.663
R448 B.n684 B.n98 256.663
R449 B.n684 B.n97 256.663
R450 B.n684 B.n96 256.663
R451 B.n684 B.n95 256.663
R452 B.n684 B.n94 256.663
R453 B.n684 B.n93 256.663
R454 B.n684 B.n92 256.663
R455 B.n684 B.n91 256.663
R456 B.n684 B.n90 256.663
R457 B.n684 B.n89 256.663
R458 B.n684 B.n88 256.663
R459 B.n684 B.n87 256.663
R460 B.n684 B.n86 256.663
R461 B.n684 B.n85 256.663
R462 B.n684 B.n84 256.663
R463 B.n684 B.n83 256.663
R464 B.n684 B.n82 256.663
R465 B.n684 B.n81 256.663
R466 B.n684 B.n80 256.663
R467 B.n684 B.n79 256.663
R468 B.n684 B.n78 256.663
R469 B.n684 B.n77 256.663
R470 B.n684 B.n76 256.663
R471 B.n684 B.n75 256.663
R472 B.n684 B.n74 256.663
R473 B.n684 B.n73 256.663
R474 B.n684 B.n72 256.663
R475 B.n684 B.n71 256.663
R476 B.n684 B.n70 256.663
R477 B.n684 B.n69 256.663
R478 B.n684 B.n68 256.663
R479 B.n684 B.n67 256.663
R480 B.n684 B.n66 256.663
R481 B.n684 B.n65 256.663
R482 B.n684 B.n64 256.663
R483 B.n684 B.n63 256.663
R484 B.n538 B.n537 256.663
R485 B.n538 B.n335 256.663
R486 B.n538 B.n336 256.663
R487 B.n538 B.n337 256.663
R488 B.n538 B.n338 256.663
R489 B.n538 B.n339 256.663
R490 B.n538 B.n340 256.663
R491 B.n538 B.n341 256.663
R492 B.n538 B.n342 256.663
R493 B.n538 B.n343 256.663
R494 B.n538 B.n344 256.663
R495 B.n538 B.n345 256.663
R496 B.n538 B.n346 256.663
R497 B.n538 B.n347 256.663
R498 B.n538 B.n348 256.663
R499 B.n538 B.n349 256.663
R500 B.n538 B.n350 256.663
R501 B.n538 B.n351 256.663
R502 B.n538 B.n352 256.663
R503 B.n538 B.n353 256.663
R504 B.n538 B.n354 256.663
R505 B.n538 B.n355 256.663
R506 B.n538 B.n356 256.663
R507 B.n538 B.n357 256.663
R508 B.n538 B.n358 256.663
R509 B.n538 B.n359 256.663
R510 B.n538 B.n360 256.663
R511 B.n538 B.n361 256.663
R512 B.n538 B.n362 256.663
R513 B.n538 B.n363 256.663
R514 B.n538 B.n364 256.663
R515 B.n538 B.n365 256.663
R516 B.n538 B.n366 256.663
R517 B.n538 B.n367 256.663
R518 B.n538 B.n368 256.663
R519 B.n538 B.n369 256.663
R520 B.n538 B.n370 256.663
R521 B.n538 B.n371 256.663
R522 B.n538 B.n372 256.663
R523 B.n539 B.n538 256.663
R524 B.n378 B.t2 248.617
R525 B.n105 B.t7 248.617
R526 B.n376 B.t12 248.617
R527 B.n107 B.t10 248.617
R528 B.n546 B.n330 163.367
R529 B.n546 B.n328 163.367
R530 B.n550 B.n328 163.367
R531 B.n550 B.n322 163.367
R532 B.n558 B.n322 163.367
R533 B.n558 B.n320 163.367
R534 B.n562 B.n320 163.367
R535 B.n562 B.n314 163.367
R536 B.n570 B.n314 163.367
R537 B.n570 B.n312 163.367
R538 B.n574 B.n312 163.367
R539 B.n574 B.n306 163.367
R540 B.n582 B.n306 163.367
R541 B.n582 B.n304 163.367
R542 B.n586 B.n304 163.367
R543 B.n586 B.n298 163.367
R544 B.n594 B.n298 163.367
R545 B.n594 B.n296 163.367
R546 B.n598 B.n296 163.367
R547 B.n598 B.n290 163.367
R548 B.n606 B.n290 163.367
R549 B.n606 B.n288 163.367
R550 B.n610 B.n288 163.367
R551 B.n610 B.n282 163.367
R552 B.n618 B.n282 163.367
R553 B.n618 B.n280 163.367
R554 B.n622 B.n280 163.367
R555 B.n622 B.n274 163.367
R556 B.n631 B.n274 163.367
R557 B.n631 B.n272 163.367
R558 B.n635 B.n272 163.367
R559 B.n635 B.n2 163.367
R560 B.n751 B.n2 163.367
R561 B.n751 B.n3 163.367
R562 B.n747 B.n3 163.367
R563 B.n747 B.n9 163.367
R564 B.n743 B.n9 163.367
R565 B.n743 B.n11 163.367
R566 B.n739 B.n11 163.367
R567 B.n739 B.n16 163.367
R568 B.n735 B.n16 163.367
R569 B.n735 B.n18 163.367
R570 B.n731 B.n18 163.367
R571 B.n731 B.n23 163.367
R572 B.n727 B.n23 163.367
R573 B.n727 B.n25 163.367
R574 B.n723 B.n25 163.367
R575 B.n723 B.n30 163.367
R576 B.n719 B.n30 163.367
R577 B.n719 B.n32 163.367
R578 B.n715 B.n32 163.367
R579 B.n715 B.n37 163.367
R580 B.n711 B.n37 163.367
R581 B.n711 B.n39 163.367
R582 B.n707 B.n39 163.367
R583 B.n707 B.n44 163.367
R584 B.n703 B.n44 163.367
R585 B.n703 B.n46 163.367
R586 B.n699 B.n46 163.367
R587 B.n699 B.n51 163.367
R588 B.n695 B.n51 163.367
R589 B.n695 B.n53 163.367
R590 B.n691 B.n53 163.367
R591 B.n691 B.n58 163.367
R592 B.n687 B.n58 163.367
R593 B.n687 B.n60 163.367
R594 B.n374 B.n373 163.367
R595 B.n531 B.n373 163.367
R596 B.n529 B.n528 163.367
R597 B.n525 B.n524 163.367
R598 B.n521 B.n520 163.367
R599 B.n517 B.n516 163.367
R600 B.n513 B.n512 163.367
R601 B.n509 B.n508 163.367
R602 B.n505 B.n504 163.367
R603 B.n501 B.n500 163.367
R604 B.n497 B.n496 163.367
R605 B.n493 B.n492 163.367
R606 B.n489 B.n488 163.367
R607 B.n485 B.n484 163.367
R608 B.n481 B.n480 163.367
R609 B.n477 B.n476 163.367
R610 B.n473 B.n472 163.367
R611 B.n469 B.n468 163.367
R612 B.n464 B.n463 163.367
R613 B.n460 B.n459 163.367
R614 B.n456 B.n455 163.367
R615 B.n452 B.n451 163.367
R616 B.n448 B.n447 163.367
R617 B.n444 B.n443 163.367
R618 B.n440 B.n439 163.367
R619 B.n436 B.n435 163.367
R620 B.n432 B.n431 163.367
R621 B.n428 B.n427 163.367
R622 B.n424 B.n423 163.367
R623 B.n420 B.n419 163.367
R624 B.n416 B.n415 163.367
R625 B.n412 B.n411 163.367
R626 B.n408 B.n407 163.367
R627 B.n404 B.n403 163.367
R628 B.n400 B.n399 163.367
R629 B.n396 B.n395 163.367
R630 B.n392 B.n391 163.367
R631 B.n388 B.n387 163.367
R632 B.n384 B.n383 163.367
R633 B.n380 B.n334 163.367
R634 B.n544 B.n332 163.367
R635 B.n544 B.n326 163.367
R636 B.n552 B.n326 163.367
R637 B.n552 B.n324 163.367
R638 B.n556 B.n324 163.367
R639 B.n556 B.n318 163.367
R640 B.n564 B.n318 163.367
R641 B.n564 B.n316 163.367
R642 B.n568 B.n316 163.367
R643 B.n568 B.n310 163.367
R644 B.n576 B.n310 163.367
R645 B.n576 B.n308 163.367
R646 B.n580 B.n308 163.367
R647 B.n580 B.n302 163.367
R648 B.n588 B.n302 163.367
R649 B.n588 B.n300 163.367
R650 B.n592 B.n300 163.367
R651 B.n592 B.n294 163.367
R652 B.n600 B.n294 163.367
R653 B.n600 B.n292 163.367
R654 B.n604 B.n292 163.367
R655 B.n604 B.n286 163.367
R656 B.n612 B.n286 163.367
R657 B.n612 B.n284 163.367
R658 B.n616 B.n284 163.367
R659 B.n616 B.n278 163.367
R660 B.n624 B.n278 163.367
R661 B.n624 B.n276 163.367
R662 B.n629 B.n276 163.367
R663 B.n629 B.n270 163.367
R664 B.n637 B.n270 163.367
R665 B.n638 B.n637 163.367
R666 B.n638 B.n5 163.367
R667 B.n6 B.n5 163.367
R668 B.n7 B.n6 163.367
R669 B.n643 B.n7 163.367
R670 B.n643 B.n12 163.367
R671 B.n13 B.n12 163.367
R672 B.n14 B.n13 163.367
R673 B.n648 B.n14 163.367
R674 B.n648 B.n19 163.367
R675 B.n20 B.n19 163.367
R676 B.n21 B.n20 163.367
R677 B.n653 B.n21 163.367
R678 B.n653 B.n26 163.367
R679 B.n27 B.n26 163.367
R680 B.n28 B.n27 163.367
R681 B.n658 B.n28 163.367
R682 B.n658 B.n33 163.367
R683 B.n34 B.n33 163.367
R684 B.n35 B.n34 163.367
R685 B.n663 B.n35 163.367
R686 B.n663 B.n40 163.367
R687 B.n41 B.n40 163.367
R688 B.n42 B.n41 163.367
R689 B.n668 B.n42 163.367
R690 B.n668 B.n47 163.367
R691 B.n48 B.n47 163.367
R692 B.n49 B.n48 163.367
R693 B.n673 B.n49 163.367
R694 B.n673 B.n54 163.367
R695 B.n55 B.n54 163.367
R696 B.n56 B.n55 163.367
R697 B.n678 B.n56 163.367
R698 B.n678 B.n61 163.367
R699 B.n62 B.n61 163.367
R700 B.n113 B.n112 163.367
R701 B.n117 B.n116 163.367
R702 B.n121 B.n120 163.367
R703 B.n125 B.n124 163.367
R704 B.n129 B.n128 163.367
R705 B.n133 B.n132 163.367
R706 B.n137 B.n136 163.367
R707 B.n141 B.n140 163.367
R708 B.n145 B.n144 163.367
R709 B.n149 B.n148 163.367
R710 B.n153 B.n152 163.367
R711 B.n157 B.n156 163.367
R712 B.n161 B.n160 163.367
R713 B.n165 B.n164 163.367
R714 B.n169 B.n168 163.367
R715 B.n173 B.n172 163.367
R716 B.n177 B.n176 163.367
R717 B.n181 B.n180 163.367
R718 B.n185 B.n184 163.367
R719 B.n189 B.n188 163.367
R720 B.n193 B.n192 163.367
R721 B.n197 B.n196 163.367
R722 B.n202 B.n201 163.367
R723 B.n206 B.n205 163.367
R724 B.n210 B.n209 163.367
R725 B.n214 B.n213 163.367
R726 B.n218 B.n217 163.367
R727 B.n222 B.n221 163.367
R728 B.n226 B.n225 163.367
R729 B.n230 B.n229 163.367
R730 B.n234 B.n233 163.367
R731 B.n238 B.n237 163.367
R732 B.n242 B.n241 163.367
R733 B.n246 B.n245 163.367
R734 B.n250 B.n249 163.367
R735 B.n254 B.n253 163.367
R736 B.n258 B.n257 163.367
R737 B.n262 B.n261 163.367
R738 B.n266 B.n265 163.367
R739 B.n683 B.n103 163.367
R740 B.n378 B.n377 81.455
R741 B.n376 B.n375 81.455
R742 B.n107 B.n106 81.455
R743 B.n105 B.n104 81.455
R744 B.n538 B.n331 79.6742
R745 B.n685 B.n684 79.6742
R746 B.n537 B.n536 71.676
R747 B.n531 B.n335 71.676
R748 B.n528 B.n336 71.676
R749 B.n524 B.n337 71.676
R750 B.n520 B.n338 71.676
R751 B.n516 B.n339 71.676
R752 B.n512 B.n340 71.676
R753 B.n508 B.n341 71.676
R754 B.n504 B.n342 71.676
R755 B.n500 B.n343 71.676
R756 B.n496 B.n344 71.676
R757 B.n492 B.n345 71.676
R758 B.n488 B.n346 71.676
R759 B.n484 B.n347 71.676
R760 B.n480 B.n348 71.676
R761 B.n476 B.n349 71.676
R762 B.n472 B.n350 71.676
R763 B.n468 B.n351 71.676
R764 B.n463 B.n352 71.676
R765 B.n459 B.n353 71.676
R766 B.n455 B.n354 71.676
R767 B.n451 B.n355 71.676
R768 B.n447 B.n356 71.676
R769 B.n443 B.n357 71.676
R770 B.n439 B.n358 71.676
R771 B.n435 B.n359 71.676
R772 B.n431 B.n360 71.676
R773 B.n427 B.n361 71.676
R774 B.n423 B.n362 71.676
R775 B.n419 B.n363 71.676
R776 B.n415 B.n364 71.676
R777 B.n411 B.n365 71.676
R778 B.n407 B.n366 71.676
R779 B.n403 B.n367 71.676
R780 B.n399 B.n368 71.676
R781 B.n395 B.n369 71.676
R782 B.n391 B.n370 71.676
R783 B.n387 B.n371 71.676
R784 B.n383 B.n372 71.676
R785 B.n539 B.n334 71.676
R786 B.n109 B.n63 71.676
R787 B.n113 B.n64 71.676
R788 B.n117 B.n65 71.676
R789 B.n121 B.n66 71.676
R790 B.n125 B.n67 71.676
R791 B.n129 B.n68 71.676
R792 B.n133 B.n69 71.676
R793 B.n137 B.n70 71.676
R794 B.n141 B.n71 71.676
R795 B.n145 B.n72 71.676
R796 B.n149 B.n73 71.676
R797 B.n153 B.n74 71.676
R798 B.n157 B.n75 71.676
R799 B.n161 B.n76 71.676
R800 B.n165 B.n77 71.676
R801 B.n169 B.n78 71.676
R802 B.n173 B.n79 71.676
R803 B.n177 B.n80 71.676
R804 B.n181 B.n81 71.676
R805 B.n185 B.n82 71.676
R806 B.n189 B.n83 71.676
R807 B.n193 B.n84 71.676
R808 B.n197 B.n85 71.676
R809 B.n202 B.n86 71.676
R810 B.n206 B.n87 71.676
R811 B.n210 B.n88 71.676
R812 B.n214 B.n89 71.676
R813 B.n218 B.n90 71.676
R814 B.n222 B.n91 71.676
R815 B.n226 B.n92 71.676
R816 B.n230 B.n93 71.676
R817 B.n234 B.n94 71.676
R818 B.n238 B.n95 71.676
R819 B.n242 B.n96 71.676
R820 B.n246 B.n97 71.676
R821 B.n250 B.n98 71.676
R822 B.n254 B.n99 71.676
R823 B.n258 B.n100 71.676
R824 B.n262 B.n101 71.676
R825 B.n266 B.n102 71.676
R826 B.n103 B.n102 71.676
R827 B.n265 B.n101 71.676
R828 B.n261 B.n100 71.676
R829 B.n257 B.n99 71.676
R830 B.n253 B.n98 71.676
R831 B.n249 B.n97 71.676
R832 B.n245 B.n96 71.676
R833 B.n241 B.n95 71.676
R834 B.n237 B.n94 71.676
R835 B.n233 B.n93 71.676
R836 B.n229 B.n92 71.676
R837 B.n225 B.n91 71.676
R838 B.n221 B.n90 71.676
R839 B.n217 B.n89 71.676
R840 B.n213 B.n88 71.676
R841 B.n209 B.n87 71.676
R842 B.n205 B.n86 71.676
R843 B.n201 B.n85 71.676
R844 B.n196 B.n84 71.676
R845 B.n192 B.n83 71.676
R846 B.n188 B.n82 71.676
R847 B.n184 B.n81 71.676
R848 B.n180 B.n80 71.676
R849 B.n176 B.n79 71.676
R850 B.n172 B.n78 71.676
R851 B.n168 B.n77 71.676
R852 B.n164 B.n76 71.676
R853 B.n160 B.n75 71.676
R854 B.n156 B.n74 71.676
R855 B.n152 B.n73 71.676
R856 B.n148 B.n72 71.676
R857 B.n144 B.n71 71.676
R858 B.n140 B.n70 71.676
R859 B.n136 B.n69 71.676
R860 B.n132 B.n68 71.676
R861 B.n128 B.n67 71.676
R862 B.n124 B.n66 71.676
R863 B.n120 B.n65 71.676
R864 B.n116 B.n64 71.676
R865 B.n112 B.n63 71.676
R866 B.n537 B.n374 71.676
R867 B.n529 B.n335 71.676
R868 B.n525 B.n336 71.676
R869 B.n521 B.n337 71.676
R870 B.n517 B.n338 71.676
R871 B.n513 B.n339 71.676
R872 B.n509 B.n340 71.676
R873 B.n505 B.n341 71.676
R874 B.n501 B.n342 71.676
R875 B.n497 B.n343 71.676
R876 B.n493 B.n344 71.676
R877 B.n489 B.n345 71.676
R878 B.n485 B.n346 71.676
R879 B.n481 B.n347 71.676
R880 B.n477 B.n348 71.676
R881 B.n473 B.n349 71.676
R882 B.n469 B.n350 71.676
R883 B.n464 B.n351 71.676
R884 B.n460 B.n352 71.676
R885 B.n456 B.n353 71.676
R886 B.n452 B.n354 71.676
R887 B.n448 B.n355 71.676
R888 B.n444 B.n356 71.676
R889 B.n440 B.n357 71.676
R890 B.n436 B.n358 71.676
R891 B.n432 B.n359 71.676
R892 B.n428 B.n360 71.676
R893 B.n424 B.n361 71.676
R894 B.n420 B.n362 71.676
R895 B.n416 B.n363 71.676
R896 B.n412 B.n364 71.676
R897 B.n408 B.n365 71.676
R898 B.n404 B.n366 71.676
R899 B.n400 B.n367 71.676
R900 B.n396 B.n368 71.676
R901 B.n392 B.n369 71.676
R902 B.n388 B.n370 71.676
R903 B.n384 B.n371 71.676
R904 B.n380 B.n372 71.676
R905 B.n540 B.n539 71.676
R906 B.n379 B.n378 59.5399
R907 B.n466 B.n376 59.5399
R908 B.n108 B.n107 59.5399
R909 B.n199 B.n105 59.5399
R910 B.n545 B.n331 48.8096
R911 B.n545 B.n327 48.8096
R912 B.n551 B.n327 48.8096
R913 B.n551 B.n323 48.8096
R914 B.n557 B.n323 48.8096
R915 B.n557 B.n319 48.8096
R916 B.n563 B.n319 48.8096
R917 B.n563 B.n315 48.8096
R918 B.n569 B.n315 48.8096
R919 B.n575 B.n311 48.8096
R920 B.n575 B.n307 48.8096
R921 B.n581 B.n307 48.8096
R922 B.n581 B.n303 48.8096
R923 B.n587 B.n303 48.8096
R924 B.n587 B.n299 48.8096
R925 B.n593 B.n299 48.8096
R926 B.n593 B.n295 48.8096
R927 B.n599 B.n295 48.8096
R928 B.n599 B.n291 48.8096
R929 B.n605 B.n291 48.8096
R930 B.n605 B.n287 48.8096
R931 B.n611 B.n287 48.8096
R932 B.n611 B.n283 48.8096
R933 B.n617 B.n283 48.8096
R934 B.n623 B.n279 48.8096
R935 B.n623 B.n275 48.8096
R936 B.n630 B.n275 48.8096
R937 B.n630 B.n271 48.8096
R938 B.n636 B.n271 48.8096
R939 B.n636 B.n4 48.8096
R940 B.n750 B.n4 48.8096
R941 B.n750 B.n749 48.8096
R942 B.n749 B.n748 48.8096
R943 B.n748 B.n8 48.8096
R944 B.n742 B.n8 48.8096
R945 B.n742 B.n741 48.8096
R946 B.n741 B.n740 48.8096
R947 B.n740 B.n15 48.8096
R948 B.n734 B.n733 48.8096
R949 B.n733 B.n732 48.8096
R950 B.n732 B.n22 48.8096
R951 B.n726 B.n22 48.8096
R952 B.n726 B.n725 48.8096
R953 B.n725 B.n724 48.8096
R954 B.n724 B.n29 48.8096
R955 B.n718 B.n29 48.8096
R956 B.n718 B.n717 48.8096
R957 B.n717 B.n716 48.8096
R958 B.n716 B.n36 48.8096
R959 B.n710 B.n36 48.8096
R960 B.n710 B.n709 48.8096
R961 B.n709 B.n708 48.8096
R962 B.n708 B.n43 48.8096
R963 B.n702 B.n701 48.8096
R964 B.n701 B.n700 48.8096
R965 B.n700 B.n50 48.8096
R966 B.n694 B.n50 48.8096
R967 B.n694 B.n693 48.8096
R968 B.n693 B.n692 48.8096
R969 B.n692 B.n57 48.8096
R970 B.n686 B.n57 48.8096
R971 B.n686 B.n685 48.8096
R972 B.t14 B.n279 38.0429
R973 B.t15 B.n15 38.0429
R974 B.n110 B.n59 32.3127
R975 B.n682 B.n681 32.3127
R976 B.n542 B.n541 32.3127
R977 B.n535 B.n329 32.3127
R978 B.n569 B.t1 32.3007
R979 B.n702 B.t5 32.3007
R980 B B.n752 18.0485
R981 B.t1 B.n311 16.5095
R982 B.t5 B.n43 16.5095
R983 B.n617 B.t14 10.7672
R984 B.n734 B.t15 10.7672
R985 B.n111 B.n110 10.6151
R986 B.n114 B.n111 10.6151
R987 B.n115 B.n114 10.6151
R988 B.n118 B.n115 10.6151
R989 B.n119 B.n118 10.6151
R990 B.n122 B.n119 10.6151
R991 B.n123 B.n122 10.6151
R992 B.n126 B.n123 10.6151
R993 B.n127 B.n126 10.6151
R994 B.n130 B.n127 10.6151
R995 B.n131 B.n130 10.6151
R996 B.n134 B.n131 10.6151
R997 B.n135 B.n134 10.6151
R998 B.n138 B.n135 10.6151
R999 B.n139 B.n138 10.6151
R1000 B.n142 B.n139 10.6151
R1001 B.n143 B.n142 10.6151
R1002 B.n146 B.n143 10.6151
R1003 B.n147 B.n146 10.6151
R1004 B.n150 B.n147 10.6151
R1005 B.n151 B.n150 10.6151
R1006 B.n154 B.n151 10.6151
R1007 B.n155 B.n154 10.6151
R1008 B.n158 B.n155 10.6151
R1009 B.n159 B.n158 10.6151
R1010 B.n162 B.n159 10.6151
R1011 B.n163 B.n162 10.6151
R1012 B.n166 B.n163 10.6151
R1013 B.n167 B.n166 10.6151
R1014 B.n170 B.n167 10.6151
R1015 B.n171 B.n170 10.6151
R1016 B.n174 B.n171 10.6151
R1017 B.n175 B.n174 10.6151
R1018 B.n178 B.n175 10.6151
R1019 B.n179 B.n178 10.6151
R1020 B.n183 B.n182 10.6151
R1021 B.n186 B.n183 10.6151
R1022 B.n187 B.n186 10.6151
R1023 B.n190 B.n187 10.6151
R1024 B.n191 B.n190 10.6151
R1025 B.n194 B.n191 10.6151
R1026 B.n195 B.n194 10.6151
R1027 B.n198 B.n195 10.6151
R1028 B.n203 B.n200 10.6151
R1029 B.n204 B.n203 10.6151
R1030 B.n207 B.n204 10.6151
R1031 B.n208 B.n207 10.6151
R1032 B.n211 B.n208 10.6151
R1033 B.n212 B.n211 10.6151
R1034 B.n215 B.n212 10.6151
R1035 B.n216 B.n215 10.6151
R1036 B.n219 B.n216 10.6151
R1037 B.n220 B.n219 10.6151
R1038 B.n223 B.n220 10.6151
R1039 B.n224 B.n223 10.6151
R1040 B.n227 B.n224 10.6151
R1041 B.n228 B.n227 10.6151
R1042 B.n231 B.n228 10.6151
R1043 B.n232 B.n231 10.6151
R1044 B.n235 B.n232 10.6151
R1045 B.n236 B.n235 10.6151
R1046 B.n239 B.n236 10.6151
R1047 B.n240 B.n239 10.6151
R1048 B.n243 B.n240 10.6151
R1049 B.n244 B.n243 10.6151
R1050 B.n247 B.n244 10.6151
R1051 B.n248 B.n247 10.6151
R1052 B.n251 B.n248 10.6151
R1053 B.n252 B.n251 10.6151
R1054 B.n255 B.n252 10.6151
R1055 B.n256 B.n255 10.6151
R1056 B.n259 B.n256 10.6151
R1057 B.n260 B.n259 10.6151
R1058 B.n263 B.n260 10.6151
R1059 B.n264 B.n263 10.6151
R1060 B.n267 B.n264 10.6151
R1061 B.n268 B.n267 10.6151
R1062 B.n682 B.n268 10.6151
R1063 B.n543 B.n542 10.6151
R1064 B.n543 B.n325 10.6151
R1065 B.n553 B.n325 10.6151
R1066 B.n554 B.n553 10.6151
R1067 B.n555 B.n554 10.6151
R1068 B.n555 B.n317 10.6151
R1069 B.n565 B.n317 10.6151
R1070 B.n566 B.n565 10.6151
R1071 B.n567 B.n566 10.6151
R1072 B.n567 B.n309 10.6151
R1073 B.n577 B.n309 10.6151
R1074 B.n578 B.n577 10.6151
R1075 B.n579 B.n578 10.6151
R1076 B.n579 B.n301 10.6151
R1077 B.n589 B.n301 10.6151
R1078 B.n590 B.n589 10.6151
R1079 B.n591 B.n590 10.6151
R1080 B.n591 B.n293 10.6151
R1081 B.n601 B.n293 10.6151
R1082 B.n602 B.n601 10.6151
R1083 B.n603 B.n602 10.6151
R1084 B.n603 B.n285 10.6151
R1085 B.n613 B.n285 10.6151
R1086 B.n614 B.n613 10.6151
R1087 B.n615 B.n614 10.6151
R1088 B.n615 B.n277 10.6151
R1089 B.n625 B.n277 10.6151
R1090 B.n626 B.n625 10.6151
R1091 B.n628 B.n626 10.6151
R1092 B.n628 B.n627 10.6151
R1093 B.n627 B.n269 10.6151
R1094 B.n639 B.n269 10.6151
R1095 B.n640 B.n639 10.6151
R1096 B.n641 B.n640 10.6151
R1097 B.n642 B.n641 10.6151
R1098 B.n644 B.n642 10.6151
R1099 B.n645 B.n644 10.6151
R1100 B.n646 B.n645 10.6151
R1101 B.n647 B.n646 10.6151
R1102 B.n649 B.n647 10.6151
R1103 B.n650 B.n649 10.6151
R1104 B.n651 B.n650 10.6151
R1105 B.n652 B.n651 10.6151
R1106 B.n654 B.n652 10.6151
R1107 B.n655 B.n654 10.6151
R1108 B.n656 B.n655 10.6151
R1109 B.n657 B.n656 10.6151
R1110 B.n659 B.n657 10.6151
R1111 B.n660 B.n659 10.6151
R1112 B.n661 B.n660 10.6151
R1113 B.n662 B.n661 10.6151
R1114 B.n664 B.n662 10.6151
R1115 B.n665 B.n664 10.6151
R1116 B.n666 B.n665 10.6151
R1117 B.n667 B.n666 10.6151
R1118 B.n669 B.n667 10.6151
R1119 B.n670 B.n669 10.6151
R1120 B.n671 B.n670 10.6151
R1121 B.n672 B.n671 10.6151
R1122 B.n674 B.n672 10.6151
R1123 B.n675 B.n674 10.6151
R1124 B.n676 B.n675 10.6151
R1125 B.n677 B.n676 10.6151
R1126 B.n679 B.n677 10.6151
R1127 B.n680 B.n679 10.6151
R1128 B.n681 B.n680 10.6151
R1129 B.n535 B.n534 10.6151
R1130 B.n534 B.n533 10.6151
R1131 B.n533 B.n532 10.6151
R1132 B.n532 B.n530 10.6151
R1133 B.n530 B.n527 10.6151
R1134 B.n527 B.n526 10.6151
R1135 B.n526 B.n523 10.6151
R1136 B.n523 B.n522 10.6151
R1137 B.n522 B.n519 10.6151
R1138 B.n519 B.n518 10.6151
R1139 B.n518 B.n515 10.6151
R1140 B.n515 B.n514 10.6151
R1141 B.n514 B.n511 10.6151
R1142 B.n511 B.n510 10.6151
R1143 B.n510 B.n507 10.6151
R1144 B.n507 B.n506 10.6151
R1145 B.n506 B.n503 10.6151
R1146 B.n503 B.n502 10.6151
R1147 B.n502 B.n499 10.6151
R1148 B.n499 B.n498 10.6151
R1149 B.n498 B.n495 10.6151
R1150 B.n495 B.n494 10.6151
R1151 B.n494 B.n491 10.6151
R1152 B.n491 B.n490 10.6151
R1153 B.n490 B.n487 10.6151
R1154 B.n487 B.n486 10.6151
R1155 B.n486 B.n483 10.6151
R1156 B.n483 B.n482 10.6151
R1157 B.n482 B.n479 10.6151
R1158 B.n479 B.n478 10.6151
R1159 B.n478 B.n475 10.6151
R1160 B.n475 B.n474 10.6151
R1161 B.n474 B.n471 10.6151
R1162 B.n471 B.n470 10.6151
R1163 B.n470 B.n467 10.6151
R1164 B.n465 B.n462 10.6151
R1165 B.n462 B.n461 10.6151
R1166 B.n461 B.n458 10.6151
R1167 B.n458 B.n457 10.6151
R1168 B.n457 B.n454 10.6151
R1169 B.n454 B.n453 10.6151
R1170 B.n453 B.n450 10.6151
R1171 B.n450 B.n449 10.6151
R1172 B.n446 B.n445 10.6151
R1173 B.n445 B.n442 10.6151
R1174 B.n442 B.n441 10.6151
R1175 B.n441 B.n438 10.6151
R1176 B.n438 B.n437 10.6151
R1177 B.n437 B.n434 10.6151
R1178 B.n434 B.n433 10.6151
R1179 B.n433 B.n430 10.6151
R1180 B.n430 B.n429 10.6151
R1181 B.n429 B.n426 10.6151
R1182 B.n426 B.n425 10.6151
R1183 B.n425 B.n422 10.6151
R1184 B.n422 B.n421 10.6151
R1185 B.n421 B.n418 10.6151
R1186 B.n418 B.n417 10.6151
R1187 B.n417 B.n414 10.6151
R1188 B.n414 B.n413 10.6151
R1189 B.n413 B.n410 10.6151
R1190 B.n410 B.n409 10.6151
R1191 B.n409 B.n406 10.6151
R1192 B.n406 B.n405 10.6151
R1193 B.n405 B.n402 10.6151
R1194 B.n402 B.n401 10.6151
R1195 B.n401 B.n398 10.6151
R1196 B.n398 B.n397 10.6151
R1197 B.n397 B.n394 10.6151
R1198 B.n394 B.n393 10.6151
R1199 B.n393 B.n390 10.6151
R1200 B.n390 B.n389 10.6151
R1201 B.n389 B.n386 10.6151
R1202 B.n386 B.n385 10.6151
R1203 B.n385 B.n382 10.6151
R1204 B.n382 B.n381 10.6151
R1205 B.n381 B.n333 10.6151
R1206 B.n541 B.n333 10.6151
R1207 B.n547 B.n329 10.6151
R1208 B.n548 B.n547 10.6151
R1209 B.n549 B.n548 10.6151
R1210 B.n549 B.n321 10.6151
R1211 B.n559 B.n321 10.6151
R1212 B.n560 B.n559 10.6151
R1213 B.n561 B.n560 10.6151
R1214 B.n561 B.n313 10.6151
R1215 B.n571 B.n313 10.6151
R1216 B.n572 B.n571 10.6151
R1217 B.n573 B.n572 10.6151
R1218 B.n573 B.n305 10.6151
R1219 B.n583 B.n305 10.6151
R1220 B.n584 B.n583 10.6151
R1221 B.n585 B.n584 10.6151
R1222 B.n585 B.n297 10.6151
R1223 B.n595 B.n297 10.6151
R1224 B.n596 B.n595 10.6151
R1225 B.n597 B.n596 10.6151
R1226 B.n597 B.n289 10.6151
R1227 B.n607 B.n289 10.6151
R1228 B.n608 B.n607 10.6151
R1229 B.n609 B.n608 10.6151
R1230 B.n609 B.n281 10.6151
R1231 B.n619 B.n281 10.6151
R1232 B.n620 B.n619 10.6151
R1233 B.n621 B.n620 10.6151
R1234 B.n621 B.n273 10.6151
R1235 B.n632 B.n273 10.6151
R1236 B.n633 B.n632 10.6151
R1237 B.n634 B.n633 10.6151
R1238 B.n634 B.n0 10.6151
R1239 B.n746 B.n1 10.6151
R1240 B.n746 B.n745 10.6151
R1241 B.n745 B.n744 10.6151
R1242 B.n744 B.n10 10.6151
R1243 B.n738 B.n10 10.6151
R1244 B.n738 B.n737 10.6151
R1245 B.n737 B.n736 10.6151
R1246 B.n736 B.n17 10.6151
R1247 B.n730 B.n17 10.6151
R1248 B.n730 B.n729 10.6151
R1249 B.n729 B.n728 10.6151
R1250 B.n728 B.n24 10.6151
R1251 B.n722 B.n24 10.6151
R1252 B.n722 B.n721 10.6151
R1253 B.n721 B.n720 10.6151
R1254 B.n720 B.n31 10.6151
R1255 B.n714 B.n31 10.6151
R1256 B.n714 B.n713 10.6151
R1257 B.n713 B.n712 10.6151
R1258 B.n712 B.n38 10.6151
R1259 B.n706 B.n38 10.6151
R1260 B.n706 B.n705 10.6151
R1261 B.n705 B.n704 10.6151
R1262 B.n704 B.n45 10.6151
R1263 B.n698 B.n45 10.6151
R1264 B.n698 B.n697 10.6151
R1265 B.n697 B.n696 10.6151
R1266 B.n696 B.n52 10.6151
R1267 B.n690 B.n52 10.6151
R1268 B.n690 B.n689 10.6151
R1269 B.n689 B.n688 10.6151
R1270 B.n688 B.n59 10.6151
R1271 B.n182 B.n108 6.5566
R1272 B.n199 B.n198 6.5566
R1273 B.n466 B.n465 6.5566
R1274 B.n449 B.n379 6.5566
R1275 B.n179 B.n108 4.05904
R1276 B.n200 B.n199 4.05904
R1277 B.n467 B.n466 4.05904
R1278 B.n446 B.n379 4.05904
R1279 B.n752 B.n0 2.81026
R1280 B.n752 B.n1 2.81026
R1281 VP.n0 VP.t1 144.169
R1282 VP.n0 VP.t0 97.6229
R1283 VP VP.n0 0.621237
R1284 VTAIL.n210 VTAIL.n162 289.615
R1285 VTAIL.n48 VTAIL.n0 289.615
R1286 VTAIL.n156 VTAIL.n108 289.615
R1287 VTAIL.n102 VTAIL.n54 289.615
R1288 VTAIL.n178 VTAIL.n177 185
R1289 VTAIL.n183 VTAIL.n182 185
R1290 VTAIL.n185 VTAIL.n184 185
R1291 VTAIL.n174 VTAIL.n173 185
R1292 VTAIL.n191 VTAIL.n190 185
R1293 VTAIL.n193 VTAIL.n192 185
R1294 VTAIL.n170 VTAIL.n169 185
R1295 VTAIL.n200 VTAIL.n199 185
R1296 VTAIL.n201 VTAIL.n168 185
R1297 VTAIL.n203 VTAIL.n202 185
R1298 VTAIL.n166 VTAIL.n165 185
R1299 VTAIL.n209 VTAIL.n208 185
R1300 VTAIL.n211 VTAIL.n210 185
R1301 VTAIL.n16 VTAIL.n15 185
R1302 VTAIL.n21 VTAIL.n20 185
R1303 VTAIL.n23 VTAIL.n22 185
R1304 VTAIL.n12 VTAIL.n11 185
R1305 VTAIL.n29 VTAIL.n28 185
R1306 VTAIL.n31 VTAIL.n30 185
R1307 VTAIL.n8 VTAIL.n7 185
R1308 VTAIL.n38 VTAIL.n37 185
R1309 VTAIL.n39 VTAIL.n6 185
R1310 VTAIL.n41 VTAIL.n40 185
R1311 VTAIL.n4 VTAIL.n3 185
R1312 VTAIL.n47 VTAIL.n46 185
R1313 VTAIL.n49 VTAIL.n48 185
R1314 VTAIL.n157 VTAIL.n156 185
R1315 VTAIL.n155 VTAIL.n154 185
R1316 VTAIL.n112 VTAIL.n111 185
R1317 VTAIL.n149 VTAIL.n148 185
R1318 VTAIL.n147 VTAIL.n114 185
R1319 VTAIL.n146 VTAIL.n145 185
R1320 VTAIL.n117 VTAIL.n115 185
R1321 VTAIL.n140 VTAIL.n139 185
R1322 VTAIL.n138 VTAIL.n137 185
R1323 VTAIL.n121 VTAIL.n120 185
R1324 VTAIL.n132 VTAIL.n131 185
R1325 VTAIL.n130 VTAIL.n129 185
R1326 VTAIL.n125 VTAIL.n124 185
R1327 VTAIL.n103 VTAIL.n102 185
R1328 VTAIL.n101 VTAIL.n100 185
R1329 VTAIL.n58 VTAIL.n57 185
R1330 VTAIL.n95 VTAIL.n94 185
R1331 VTAIL.n93 VTAIL.n60 185
R1332 VTAIL.n92 VTAIL.n91 185
R1333 VTAIL.n63 VTAIL.n61 185
R1334 VTAIL.n86 VTAIL.n85 185
R1335 VTAIL.n84 VTAIL.n83 185
R1336 VTAIL.n67 VTAIL.n66 185
R1337 VTAIL.n78 VTAIL.n77 185
R1338 VTAIL.n76 VTAIL.n75 185
R1339 VTAIL.n71 VTAIL.n70 185
R1340 VTAIL.n179 VTAIL.t1 149.524
R1341 VTAIL.n17 VTAIL.t2 149.524
R1342 VTAIL.n126 VTAIL.t3 149.524
R1343 VTAIL.n72 VTAIL.t0 149.524
R1344 VTAIL.n183 VTAIL.n177 104.615
R1345 VTAIL.n184 VTAIL.n183 104.615
R1346 VTAIL.n184 VTAIL.n173 104.615
R1347 VTAIL.n191 VTAIL.n173 104.615
R1348 VTAIL.n192 VTAIL.n191 104.615
R1349 VTAIL.n192 VTAIL.n169 104.615
R1350 VTAIL.n200 VTAIL.n169 104.615
R1351 VTAIL.n201 VTAIL.n200 104.615
R1352 VTAIL.n202 VTAIL.n201 104.615
R1353 VTAIL.n202 VTAIL.n165 104.615
R1354 VTAIL.n209 VTAIL.n165 104.615
R1355 VTAIL.n210 VTAIL.n209 104.615
R1356 VTAIL.n21 VTAIL.n15 104.615
R1357 VTAIL.n22 VTAIL.n21 104.615
R1358 VTAIL.n22 VTAIL.n11 104.615
R1359 VTAIL.n29 VTAIL.n11 104.615
R1360 VTAIL.n30 VTAIL.n29 104.615
R1361 VTAIL.n30 VTAIL.n7 104.615
R1362 VTAIL.n38 VTAIL.n7 104.615
R1363 VTAIL.n39 VTAIL.n38 104.615
R1364 VTAIL.n40 VTAIL.n39 104.615
R1365 VTAIL.n40 VTAIL.n3 104.615
R1366 VTAIL.n47 VTAIL.n3 104.615
R1367 VTAIL.n48 VTAIL.n47 104.615
R1368 VTAIL.n156 VTAIL.n155 104.615
R1369 VTAIL.n155 VTAIL.n111 104.615
R1370 VTAIL.n148 VTAIL.n111 104.615
R1371 VTAIL.n148 VTAIL.n147 104.615
R1372 VTAIL.n147 VTAIL.n146 104.615
R1373 VTAIL.n146 VTAIL.n115 104.615
R1374 VTAIL.n139 VTAIL.n115 104.615
R1375 VTAIL.n139 VTAIL.n138 104.615
R1376 VTAIL.n138 VTAIL.n120 104.615
R1377 VTAIL.n131 VTAIL.n120 104.615
R1378 VTAIL.n131 VTAIL.n130 104.615
R1379 VTAIL.n130 VTAIL.n124 104.615
R1380 VTAIL.n102 VTAIL.n101 104.615
R1381 VTAIL.n101 VTAIL.n57 104.615
R1382 VTAIL.n94 VTAIL.n57 104.615
R1383 VTAIL.n94 VTAIL.n93 104.615
R1384 VTAIL.n93 VTAIL.n92 104.615
R1385 VTAIL.n92 VTAIL.n61 104.615
R1386 VTAIL.n85 VTAIL.n61 104.615
R1387 VTAIL.n85 VTAIL.n84 104.615
R1388 VTAIL.n84 VTAIL.n66 104.615
R1389 VTAIL.n77 VTAIL.n66 104.615
R1390 VTAIL.n77 VTAIL.n76 104.615
R1391 VTAIL.n76 VTAIL.n70 104.615
R1392 VTAIL.t1 VTAIL.n177 52.3082
R1393 VTAIL.t2 VTAIL.n15 52.3082
R1394 VTAIL.t3 VTAIL.n124 52.3082
R1395 VTAIL.t0 VTAIL.n70 52.3082
R1396 VTAIL.n215 VTAIL.n214 33.9308
R1397 VTAIL.n53 VTAIL.n52 33.9308
R1398 VTAIL.n161 VTAIL.n160 33.9308
R1399 VTAIL.n107 VTAIL.n106 33.9308
R1400 VTAIL.n107 VTAIL.n53 28.2721
R1401 VTAIL.n215 VTAIL.n161 24.6514
R1402 VTAIL.n203 VTAIL.n168 13.1884
R1403 VTAIL.n41 VTAIL.n6 13.1884
R1404 VTAIL.n149 VTAIL.n114 13.1884
R1405 VTAIL.n95 VTAIL.n60 13.1884
R1406 VTAIL.n199 VTAIL.n198 12.8005
R1407 VTAIL.n204 VTAIL.n166 12.8005
R1408 VTAIL.n37 VTAIL.n36 12.8005
R1409 VTAIL.n42 VTAIL.n4 12.8005
R1410 VTAIL.n150 VTAIL.n112 12.8005
R1411 VTAIL.n145 VTAIL.n116 12.8005
R1412 VTAIL.n96 VTAIL.n58 12.8005
R1413 VTAIL.n91 VTAIL.n62 12.8005
R1414 VTAIL.n197 VTAIL.n170 12.0247
R1415 VTAIL.n208 VTAIL.n207 12.0247
R1416 VTAIL.n35 VTAIL.n8 12.0247
R1417 VTAIL.n46 VTAIL.n45 12.0247
R1418 VTAIL.n154 VTAIL.n153 12.0247
R1419 VTAIL.n144 VTAIL.n117 12.0247
R1420 VTAIL.n100 VTAIL.n99 12.0247
R1421 VTAIL.n90 VTAIL.n63 12.0247
R1422 VTAIL.n194 VTAIL.n193 11.249
R1423 VTAIL.n211 VTAIL.n164 11.249
R1424 VTAIL.n32 VTAIL.n31 11.249
R1425 VTAIL.n49 VTAIL.n2 11.249
R1426 VTAIL.n157 VTAIL.n110 11.249
R1427 VTAIL.n141 VTAIL.n140 11.249
R1428 VTAIL.n103 VTAIL.n56 11.249
R1429 VTAIL.n87 VTAIL.n86 11.249
R1430 VTAIL.n190 VTAIL.n172 10.4732
R1431 VTAIL.n212 VTAIL.n162 10.4732
R1432 VTAIL.n28 VTAIL.n10 10.4732
R1433 VTAIL.n50 VTAIL.n0 10.4732
R1434 VTAIL.n158 VTAIL.n108 10.4732
R1435 VTAIL.n137 VTAIL.n119 10.4732
R1436 VTAIL.n104 VTAIL.n54 10.4732
R1437 VTAIL.n83 VTAIL.n65 10.4732
R1438 VTAIL.n179 VTAIL.n178 10.2747
R1439 VTAIL.n17 VTAIL.n16 10.2747
R1440 VTAIL.n126 VTAIL.n125 10.2747
R1441 VTAIL.n72 VTAIL.n71 10.2747
R1442 VTAIL.n189 VTAIL.n174 9.69747
R1443 VTAIL.n27 VTAIL.n12 9.69747
R1444 VTAIL.n136 VTAIL.n121 9.69747
R1445 VTAIL.n82 VTAIL.n67 9.69747
R1446 VTAIL.n214 VTAIL.n213 9.45567
R1447 VTAIL.n52 VTAIL.n51 9.45567
R1448 VTAIL.n160 VTAIL.n159 9.45567
R1449 VTAIL.n106 VTAIL.n105 9.45567
R1450 VTAIL.n213 VTAIL.n212 9.3005
R1451 VTAIL.n164 VTAIL.n163 9.3005
R1452 VTAIL.n207 VTAIL.n206 9.3005
R1453 VTAIL.n205 VTAIL.n204 9.3005
R1454 VTAIL.n181 VTAIL.n180 9.3005
R1455 VTAIL.n176 VTAIL.n175 9.3005
R1456 VTAIL.n187 VTAIL.n186 9.3005
R1457 VTAIL.n189 VTAIL.n188 9.3005
R1458 VTAIL.n172 VTAIL.n171 9.3005
R1459 VTAIL.n195 VTAIL.n194 9.3005
R1460 VTAIL.n197 VTAIL.n196 9.3005
R1461 VTAIL.n198 VTAIL.n167 9.3005
R1462 VTAIL.n51 VTAIL.n50 9.3005
R1463 VTAIL.n2 VTAIL.n1 9.3005
R1464 VTAIL.n45 VTAIL.n44 9.3005
R1465 VTAIL.n43 VTAIL.n42 9.3005
R1466 VTAIL.n19 VTAIL.n18 9.3005
R1467 VTAIL.n14 VTAIL.n13 9.3005
R1468 VTAIL.n25 VTAIL.n24 9.3005
R1469 VTAIL.n27 VTAIL.n26 9.3005
R1470 VTAIL.n10 VTAIL.n9 9.3005
R1471 VTAIL.n33 VTAIL.n32 9.3005
R1472 VTAIL.n35 VTAIL.n34 9.3005
R1473 VTAIL.n36 VTAIL.n5 9.3005
R1474 VTAIL.n128 VTAIL.n127 9.3005
R1475 VTAIL.n123 VTAIL.n122 9.3005
R1476 VTAIL.n134 VTAIL.n133 9.3005
R1477 VTAIL.n136 VTAIL.n135 9.3005
R1478 VTAIL.n119 VTAIL.n118 9.3005
R1479 VTAIL.n142 VTAIL.n141 9.3005
R1480 VTAIL.n144 VTAIL.n143 9.3005
R1481 VTAIL.n116 VTAIL.n113 9.3005
R1482 VTAIL.n159 VTAIL.n158 9.3005
R1483 VTAIL.n110 VTAIL.n109 9.3005
R1484 VTAIL.n153 VTAIL.n152 9.3005
R1485 VTAIL.n151 VTAIL.n150 9.3005
R1486 VTAIL.n74 VTAIL.n73 9.3005
R1487 VTAIL.n69 VTAIL.n68 9.3005
R1488 VTAIL.n80 VTAIL.n79 9.3005
R1489 VTAIL.n82 VTAIL.n81 9.3005
R1490 VTAIL.n65 VTAIL.n64 9.3005
R1491 VTAIL.n88 VTAIL.n87 9.3005
R1492 VTAIL.n90 VTAIL.n89 9.3005
R1493 VTAIL.n62 VTAIL.n59 9.3005
R1494 VTAIL.n105 VTAIL.n104 9.3005
R1495 VTAIL.n56 VTAIL.n55 9.3005
R1496 VTAIL.n99 VTAIL.n98 9.3005
R1497 VTAIL.n97 VTAIL.n96 9.3005
R1498 VTAIL.n186 VTAIL.n185 8.92171
R1499 VTAIL.n24 VTAIL.n23 8.92171
R1500 VTAIL.n133 VTAIL.n132 8.92171
R1501 VTAIL.n79 VTAIL.n78 8.92171
R1502 VTAIL.n182 VTAIL.n176 8.14595
R1503 VTAIL.n20 VTAIL.n14 8.14595
R1504 VTAIL.n129 VTAIL.n123 8.14595
R1505 VTAIL.n75 VTAIL.n69 8.14595
R1506 VTAIL.n181 VTAIL.n178 7.3702
R1507 VTAIL.n19 VTAIL.n16 7.3702
R1508 VTAIL.n128 VTAIL.n125 7.3702
R1509 VTAIL.n74 VTAIL.n71 7.3702
R1510 VTAIL.n182 VTAIL.n181 5.81868
R1511 VTAIL.n20 VTAIL.n19 5.81868
R1512 VTAIL.n129 VTAIL.n128 5.81868
R1513 VTAIL.n75 VTAIL.n74 5.81868
R1514 VTAIL.n185 VTAIL.n176 5.04292
R1515 VTAIL.n23 VTAIL.n14 5.04292
R1516 VTAIL.n132 VTAIL.n123 5.04292
R1517 VTAIL.n78 VTAIL.n69 5.04292
R1518 VTAIL.n186 VTAIL.n174 4.26717
R1519 VTAIL.n24 VTAIL.n12 4.26717
R1520 VTAIL.n133 VTAIL.n121 4.26717
R1521 VTAIL.n79 VTAIL.n67 4.26717
R1522 VTAIL.n190 VTAIL.n189 3.49141
R1523 VTAIL.n214 VTAIL.n162 3.49141
R1524 VTAIL.n28 VTAIL.n27 3.49141
R1525 VTAIL.n52 VTAIL.n0 3.49141
R1526 VTAIL.n160 VTAIL.n108 3.49141
R1527 VTAIL.n137 VTAIL.n136 3.49141
R1528 VTAIL.n106 VTAIL.n54 3.49141
R1529 VTAIL.n83 VTAIL.n82 3.49141
R1530 VTAIL.n180 VTAIL.n179 2.84303
R1531 VTAIL.n18 VTAIL.n17 2.84303
R1532 VTAIL.n127 VTAIL.n126 2.84303
R1533 VTAIL.n73 VTAIL.n72 2.84303
R1534 VTAIL.n193 VTAIL.n172 2.71565
R1535 VTAIL.n212 VTAIL.n211 2.71565
R1536 VTAIL.n31 VTAIL.n10 2.71565
R1537 VTAIL.n50 VTAIL.n49 2.71565
R1538 VTAIL.n158 VTAIL.n157 2.71565
R1539 VTAIL.n140 VTAIL.n119 2.71565
R1540 VTAIL.n104 VTAIL.n103 2.71565
R1541 VTAIL.n86 VTAIL.n65 2.71565
R1542 VTAIL.n161 VTAIL.n107 2.28067
R1543 VTAIL.n194 VTAIL.n170 1.93989
R1544 VTAIL.n208 VTAIL.n164 1.93989
R1545 VTAIL.n32 VTAIL.n8 1.93989
R1546 VTAIL.n46 VTAIL.n2 1.93989
R1547 VTAIL.n154 VTAIL.n110 1.93989
R1548 VTAIL.n141 VTAIL.n117 1.93989
R1549 VTAIL.n100 VTAIL.n56 1.93989
R1550 VTAIL.n87 VTAIL.n63 1.93989
R1551 VTAIL VTAIL.n53 1.43369
R1552 VTAIL.n199 VTAIL.n197 1.16414
R1553 VTAIL.n207 VTAIL.n166 1.16414
R1554 VTAIL.n37 VTAIL.n35 1.16414
R1555 VTAIL.n45 VTAIL.n4 1.16414
R1556 VTAIL.n153 VTAIL.n112 1.16414
R1557 VTAIL.n145 VTAIL.n144 1.16414
R1558 VTAIL.n99 VTAIL.n58 1.16414
R1559 VTAIL.n91 VTAIL.n90 1.16414
R1560 VTAIL VTAIL.n215 0.847483
R1561 VTAIL.n198 VTAIL.n168 0.388379
R1562 VTAIL.n204 VTAIL.n203 0.388379
R1563 VTAIL.n36 VTAIL.n6 0.388379
R1564 VTAIL.n42 VTAIL.n41 0.388379
R1565 VTAIL.n150 VTAIL.n149 0.388379
R1566 VTAIL.n116 VTAIL.n114 0.388379
R1567 VTAIL.n96 VTAIL.n95 0.388379
R1568 VTAIL.n62 VTAIL.n60 0.388379
R1569 VTAIL.n180 VTAIL.n175 0.155672
R1570 VTAIL.n187 VTAIL.n175 0.155672
R1571 VTAIL.n188 VTAIL.n187 0.155672
R1572 VTAIL.n188 VTAIL.n171 0.155672
R1573 VTAIL.n195 VTAIL.n171 0.155672
R1574 VTAIL.n196 VTAIL.n195 0.155672
R1575 VTAIL.n196 VTAIL.n167 0.155672
R1576 VTAIL.n205 VTAIL.n167 0.155672
R1577 VTAIL.n206 VTAIL.n205 0.155672
R1578 VTAIL.n206 VTAIL.n163 0.155672
R1579 VTAIL.n213 VTAIL.n163 0.155672
R1580 VTAIL.n18 VTAIL.n13 0.155672
R1581 VTAIL.n25 VTAIL.n13 0.155672
R1582 VTAIL.n26 VTAIL.n25 0.155672
R1583 VTAIL.n26 VTAIL.n9 0.155672
R1584 VTAIL.n33 VTAIL.n9 0.155672
R1585 VTAIL.n34 VTAIL.n33 0.155672
R1586 VTAIL.n34 VTAIL.n5 0.155672
R1587 VTAIL.n43 VTAIL.n5 0.155672
R1588 VTAIL.n44 VTAIL.n43 0.155672
R1589 VTAIL.n44 VTAIL.n1 0.155672
R1590 VTAIL.n51 VTAIL.n1 0.155672
R1591 VTAIL.n159 VTAIL.n109 0.155672
R1592 VTAIL.n152 VTAIL.n109 0.155672
R1593 VTAIL.n152 VTAIL.n151 0.155672
R1594 VTAIL.n151 VTAIL.n113 0.155672
R1595 VTAIL.n143 VTAIL.n113 0.155672
R1596 VTAIL.n143 VTAIL.n142 0.155672
R1597 VTAIL.n142 VTAIL.n118 0.155672
R1598 VTAIL.n135 VTAIL.n118 0.155672
R1599 VTAIL.n135 VTAIL.n134 0.155672
R1600 VTAIL.n134 VTAIL.n122 0.155672
R1601 VTAIL.n127 VTAIL.n122 0.155672
R1602 VTAIL.n105 VTAIL.n55 0.155672
R1603 VTAIL.n98 VTAIL.n55 0.155672
R1604 VTAIL.n98 VTAIL.n97 0.155672
R1605 VTAIL.n97 VTAIL.n59 0.155672
R1606 VTAIL.n89 VTAIL.n59 0.155672
R1607 VTAIL.n89 VTAIL.n88 0.155672
R1608 VTAIL.n88 VTAIL.n64 0.155672
R1609 VTAIL.n81 VTAIL.n64 0.155672
R1610 VTAIL.n81 VTAIL.n80 0.155672
R1611 VTAIL.n80 VTAIL.n68 0.155672
R1612 VTAIL.n73 VTAIL.n68 0.155672
R1613 VDD1.n48 VDD1.n0 289.615
R1614 VDD1.n101 VDD1.n53 289.615
R1615 VDD1.n49 VDD1.n48 185
R1616 VDD1.n47 VDD1.n46 185
R1617 VDD1.n4 VDD1.n3 185
R1618 VDD1.n41 VDD1.n40 185
R1619 VDD1.n39 VDD1.n6 185
R1620 VDD1.n38 VDD1.n37 185
R1621 VDD1.n9 VDD1.n7 185
R1622 VDD1.n32 VDD1.n31 185
R1623 VDD1.n30 VDD1.n29 185
R1624 VDD1.n13 VDD1.n12 185
R1625 VDD1.n24 VDD1.n23 185
R1626 VDD1.n22 VDD1.n21 185
R1627 VDD1.n17 VDD1.n16 185
R1628 VDD1.n69 VDD1.n68 185
R1629 VDD1.n74 VDD1.n73 185
R1630 VDD1.n76 VDD1.n75 185
R1631 VDD1.n65 VDD1.n64 185
R1632 VDD1.n82 VDD1.n81 185
R1633 VDD1.n84 VDD1.n83 185
R1634 VDD1.n61 VDD1.n60 185
R1635 VDD1.n91 VDD1.n90 185
R1636 VDD1.n92 VDD1.n59 185
R1637 VDD1.n94 VDD1.n93 185
R1638 VDD1.n57 VDD1.n56 185
R1639 VDD1.n100 VDD1.n99 185
R1640 VDD1.n102 VDD1.n101 185
R1641 VDD1.n18 VDD1.t0 149.524
R1642 VDD1.n70 VDD1.t1 149.524
R1643 VDD1.n48 VDD1.n47 104.615
R1644 VDD1.n47 VDD1.n3 104.615
R1645 VDD1.n40 VDD1.n3 104.615
R1646 VDD1.n40 VDD1.n39 104.615
R1647 VDD1.n39 VDD1.n38 104.615
R1648 VDD1.n38 VDD1.n7 104.615
R1649 VDD1.n31 VDD1.n7 104.615
R1650 VDD1.n31 VDD1.n30 104.615
R1651 VDD1.n30 VDD1.n12 104.615
R1652 VDD1.n23 VDD1.n12 104.615
R1653 VDD1.n23 VDD1.n22 104.615
R1654 VDD1.n22 VDD1.n16 104.615
R1655 VDD1.n74 VDD1.n68 104.615
R1656 VDD1.n75 VDD1.n74 104.615
R1657 VDD1.n75 VDD1.n64 104.615
R1658 VDD1.n82 VDD1.n64 104.615
R1659 VDD1.n83 VDD1.n82 104.615
R1660 VDD1.n83 VDD1.n60 104.615
R1661 VDD1.n91 VDD1.n60 104.615
R1662 VDD1.n92 VDD1.n91 104.615
R1663 VDD1.n93 VDD1.n92 104.615
R1664 VDD1.n93 VDD1.n56 104.615
R1665 VDD1.n100 VDD1.n56 104.615
R1666 VDD1.n101 VDD1.n100 104.615
R1667 VDD1 VDD1.n105 91.6042
R1668 VDD1.t0 VDD1.n16 52.3082
R1669 VDD1.t1 VDD1.n68 52.3082
R1670 VDD1 VDD1.n52 51.573
R1671 VDD1.n41 VDD1.n6 13.1884
R1672 VDD1.n94 VDD1.n59 13.1884
R1673 VDD1.n42 VDD1.n4 12.8005
R1674 VDD1.n37 VDD1.n8 12.8005
R1675 VDD1.n90 VDD1.n89 12.8005
R1676 VDD1.n95 VDD1.n57 12.8005
R1677 VDD1.n46 VDD1.n45 12.0247
R1678 VDD1.n36 VDD1.n9 12.0247
R1679 VDD1.n88 VDD1.n61 12.0247
R1680 VDD1.n99 VDD1.n98 12.0247
R1681 VDD1.n49 VDD1.n2 11.249
R1682 VDD1.n33 VDD1.n32 11.249
R1683 VDD1.n85 VDD1.n84 11.249
R1684 VDD1.n102 VDD1.n55 11.249
R1685 VDD1.n50 VDD1.n0 10.4732
R1686 VDD1.n29 VDD1.n11 10.4732
R1687 VDD1.n81 VDD1.n63 10.4732
R1688 VDD1.n103 VDD1.n53 10.4732
R1689 VDD1.n18 VDD1.n17 10.2747
R1690 VDD1.n70 VDD1.n69 10.2747
R1691 VDD1.n28 VDD1.n13 9.69747
R1692 VDD1.n80 VDD1.n65 9.69747
R1693 VDD1.n52 VDD1.n51 9.45567
R1694 VDD1.n105 VDD1.n104 9.45567
R1695 VDD1.n20 VDD1.n19 9.3005
R1696 VDD1.n15 VDD1.n14 9.3005
R1697 VDD1.n26 VDD1.n25 9.3005
R1698 VDD1.n28 VDD1.n27 9.3005
R1699 VDD1.n11 VDD1.n10 9.3005
R1700 VDD1.n34 VDD1.n33 9.3005
R1701 VDD1.n36 VDD1.n35 9.3005
R1702 VDD1.n8 VDD1.n5 9.3005
R1703 VDD1.n51 VDD1.n50 9.3005
R1704 VDD1.n2 VDD1.n1 9.3005
R1705 VDD1.n45 VDD1.n44 9.3005
R1706 VDD1.n43 VDD1.n42 9.3005
R1707 VDD1.n104 VDD1.n103 9.3005
R1708 VDD1.n55 VDD1.n54 9.3005
R1709 VDD1.n98 VDD1.n97 9.3005
R1710 VDD1.n96 VDD1.n95 9.3005
R1711 VDD1.n72 VDD1.n71 9.3005
R1712 VDD1.n67 VDD1.n66 9.3005
R1713 VDD1.n78 VDD1.n77 9.3005
R1714 VDD1.n80 VDD1.n79 9.3005
R1715 VDD1.n63 VDD1.n62 9.3005
R1716 VDD1.n86 VDD1.n85 9.3005
R1717 VDD1.n88 VDD1.n87 9.3005
R1718 VDD1.n89 VDD1.n58 9.3005
R1719 VDD1.n25 VDD1.n24 8.92171
R1720 VDD1.n77 VDD1.n76 8.92171
R1721 VDD1.n21 VDD1.n15 8.14595
R1722 VDD1.n73 VDD1.n67 8.14595
R1723 VDD1.n20 VDD1.n17 7.3702
R1724 VDD1.n72 VDD1.n69 7.3702
R1725 VDD1.n21 VDD1.n20 5.81868
R1726 VDD1.n73 VDD1.n72 5.81868
R1727 VDD1.n24 VDD1.n15 5.04292
R1728 VDD1.n76 VDD1.n67 5.04292
R1729 VDD1.n25 VDD1.n13 4.26717
R1730 VDD1.n77 VDD1.n65 4.26717
R1731 VDD1.n52 VDD1.n0 3.49141
R1732 VDD1.n29 VDD1.n28 3.49141
R1733 VDD1.n81 VDD1.n80 3.49141
R1734 VDD1.n105 VDD1.n53 3.49141
R1735 VDD1.n19 VDD1.n18 2.84303
R1736 VDD1.n71 VDD1.n70 2.84303
R1737 VDD1.n50 VDD1.n49 2.71565
R1738 VDD1.n32 VDD1.n11 2.71565
R1739 VDD1.n84 VDD1.n63 2.71565
R1740 VDD1.n103 VDD1.n102 2.71565
R1741 VDD1.n46 VDD1.n2 1.93989
R1742 VDD1.n33 VDD1.n9 1.93989
R1743 VDD1.n85 VDD1.n61 1.93989
R1744 VDD1.n99 VDD1.n55 1.93989
R1745 VDD1.n45 VDD1.n4 1.16414
R1746 VDD1.n37 VDD1.n36 1.16414
R1747 VDD1.n90 VDD1.n88 1.16414
R1748 VDD1.n98 VDD1.n57 1.16414
R1749 VDD1.n42 VDD1.n41 0.388379
R1750 VDD1.n8 VDD1.n6 0.388379
R1751 VDD1.n89 VDD1.n59 0.388379
R1752 VDD1.n95 VDD1.n94 0.388379
R1753 VDD1.n51 VDD1.n1 0.155672
R1754 VDD1.n44 VDD1.n1 0.155672
R1755 VDD1.n44 VDD1.n43 0.155672
R1756 VDD1.n43 VDD1.n5 0.155672
R1757 VDD1.n35 VDD1.n5 0.155672
R1758 VDD1.n35 VDD1.n34 0.155672
R1759 VDD1.n34 VDD1.n10 0.155672
R1760 VDD1.n27 VDD1.n10 0.155672
R1761 VDD1.n27 VDD1.n26 0.155672
R1762 VDD1.n26 VDD1.n14 0.155672
R1763 VDD1.n19 VDD1.n14 0.155672
R1764 VDD1.n71 VDD1.n66 0.155672
R1765 VDD1.n78 VDD1.n66 0.155672
R1766 VDD1.n79 VDD1.n78 0.155672
R1767 VDD1.n79 VDD1.n62 0.155672
R1768 VDD1.n86 VDD1.n62 0.155672
R1769 VDD1.n87 VDD1.n86 0.155672
R1770 VDD1.n87 VDD1.n58 0.155672
R1771 VDD1.n96 VDD1.n58 0.155672
R1772 VDD1.n97 VDD1.n96 0.155672
R1773 VDD1.n97 VDD1.n54 0.155672
R1774 VDD1.n104 VDD1.n54 0.155672
R1775 VN VN.t0 143.982
R1776 VN VN.t1 98.2436
R1777 VDD2.n101 VDD2.n53 289.615
R1778 VDD2.n48 VDD2.n0 289.615
R1779 VDD2.n102 VDD2.n101 185
R1780 VDD2.n100 VDD2.n99 185
R1781 VDD2.n57 VDD2.n56 185
R1782 VDD2.n94 VDD2.n93 185
R1783 VDD2.n92 VDD2.n59 185
R1784 VDD2.n91 VDD2.n90 185
R1785 VDD2.n62 VDD2.n60 185
R1786 VDD2.n85 VDD2.n84 185
R1787 VDD2.n83 VDD2.n82 185
R1788 VDD2.n66 VDD2.n65 185
R1789 VDD2.n77 VDD2.n76 185
R1790 VDD2.n75 VDD2.n74 185
R1791 VDD2.n70 VDD2.n69 185
R1792 VDD2.n16 VDD2.n15 185
R1793 VDD2.n21 VDD2.n20 185
R1794 VDD2.n23 VDD2.n22 185
R1795 VDD2.n12 VDD2.n11 185
R1796 VDD2.n29 VDD2.n28 185
R1797 VDD2.n31 VDD2.n30 185
R1798 VDD2.n8 VDD2.n7 185
R1799 VDD2.n38 VDD2.n37 185
R1800 VDD2.n39 VDD2.n6 185
R1801 VDD2.n41 VDD2.n40 185
R1802 VDD2.n4 VDD2.n3 185
R1803 VDD2.n47 VDD2.n46 185
R1804 VDD2.n49 VDD2.n48 185
R1805 VDD2.n71 VDD2.t1 149.524
R1806 VDD2.n17 VDD2.t0 149.524
R1807 VDD2.n101 VDD2.n100 104.615
R1808 VDD2.n100 VDD2.n56 104.615
R1809 VDD2.n93 VDD2.n56 104.615
R1810 VDD2.n93 VDD2.n92 104.615
R1811 VDD2.n92 VDD2.n91 104.615
R1812 VDD2.n91 VDD2.n60 104.615
R1813 VDD2.n84 VDD2.n60 104.615
R1814 VDD2.n84 VDD2.n83 104.615
R1815 VDD2.n83 VDD2.n65 104.615
R1816 VDD2.n76 VDD2.n65 104.615
R1817 VDD2.n76 VDD2.n75 104.615
R1818 VDD2.n75 VDD2.n69 104.615
R1819 VDD2.n21 VDD2.n15 104.615
R1820 VDD2.n22 VDD2.n21 104.615
R1821 VDD2.n22 VDD2.n11 104.615
R1822 VDD2.n29 VDD2.n11 104.615
R1823 VDD2.n30 VDD2.n29 104.615
R1824 VDD2.n30 VDD2.n7 104.615
R1825 VDD2.n38 VDD2.n7 104.615
R1826 VDD2.n39 VDD2.n38 104.615
R1827 VDD2.n40 VDD2.n39 104.615
R1828 VDD2.n40 VDD2.n3 104.615
R1829 VDD2.n47 VDD2.n3 104.615
R1830 VDD2.n48 VDD2.n47 104.615
R1831 VDD2.n106 VDD2.n52 90.1742
R1832 VDD2.t1 VDD2.n69 52.3082
R1833 VDD2.t0 VDD2.n15 52.3082
R1834 VDD2.n106 VDD2.n105 50.6096
R1835 VDD2.n94 VDD2.n59 13.1884
R1836 VDD2.n41 VDD2.n6 13.1884
R1837 VDD2.n95 VDD2.n57 12.8005
R1838 VDD2.n90 VDD2.n61 12.8005
R1839 VDD2.n37 VDD2.n36 12.8005
R1840 VDD2.n42 VDD2.n4 12.8005
R1841 VDD2.n99 VDD2.n98 12.0247
R1842 VDD2.n89 VDD2.n62 12.0247
R1843 VDD2.n35 VDD2.n8 12.0247
R1844 VDD2.n46 VDD2.n45 12.0247
R1845 VDD2.n102 VDD2.n55 11.249
R1846 VDD2.n86 VDD2.n85 11.249
R1847 VDD2.n32 VDD2.n31 11.249
R1848 VDD2.n49 VDD2.n2 11.249
R1849 VDD2.n103 VDD2.n53 10.4732
R1850 VDD2.n82 VDD2.n64 10.4732
R1851 VDD2.n28 VDD2.n10 10.4732
R1852 VDD2.n50 VDD2.n0 10.4732
R1853 VDD2.n71 VDD2.n70 10.2747
R1854 VDD2.n17 VDD2.n16 10.2747
R1855 VDD2.n81 VDD2.n66 9.69747
R1856 VDD2.n27 VDD2.n12 9.69747
R1857 VDD2.n105 VDD2.n104 9.45567
R1858 VDD2.n52 VDD2.n51 9.45567
R1859 VDD2.n73 VDD2.n72 9.3005
R1860 VDD2.n68 VDD2.n67 9.3005
R1861 VDD2.n79 VDD2.n78 9.3005
R1862 VDD2.n81 VDD2.n80 9.3005
R1863 VDD2.n64 VDD2.n63 9.3005
R1864 VDD2.n87 VDD2.n86 9.3005
R1865 VDD2.n89 VDD2.n88 9.3005
R1866 VDD2.n61 VDD2.n58 9.3005
R1867 VDD2.n104 VDD2.n103 9.3005
R1868 VDD2.n55 VDD2.n54 9.3005
R1869 VDD2.n98 VDD2.n97 9.3005
R1870 VDD2.n96 VDD2.n95 9.3005
R1871 VDD2.n51 VDD2.n50 9.3005
R1872 VDD2.n2 VDD2.n1 9.3005
R1873 VDD2.n45 VDD2.n44 9.3005
R1874 VDD2.n43 VDD2.n42 9.3005
R1875 VDD2.n19 VDD2.n18 9.3005
R1876 VDD2.n14 VDD2.n13 9.3005
R1877 VDD2.n25 VDD2.n24 9.3005
R1878 VDD2.n27 VDD2.n26 9.3005
R1879 VDD2.n10 VDD2.n9 9.3005
R1880 VDD2.n33 VDD2.n32 9.3005
R1881 VDD2.n35 VDD2.n34 9.3005
R1882 VDD2.n36 VDD2.n5 9.3005
R1883 VDD2.n78 VDD2.n77 8.92171
R1884 VDD2.n24 VDD2.n23 8.92171
R1885 VDD2.n74 VDD2.n68 8.14595
R1886 VDD2.n20 VDD2.n14 8.14595
R1887 VDD2.n73 VDD2.n70 7.3702
R1888 VDD2.n19 VDD2.n16 7.3702
R1889 VDD2.n74 VDD2.n73 5.81868
R1890 VDD2.n20 VDD2.n19 5.81868
R1891 VDD2.n77 VDD2.n68 5.04292
R1892 VDD2.n23 VDD2.n14 5.04292
R1893 VDD2.n78 VDD2.n66 4.26717
R1894 VDD2.n24 VDD2.n12 4.26717
R1895 VDD2.n105 VDD2.n53 3.49141
R1896 VDD2.n82 VDD2.n81 3.49141
R1897 VDD2.n28 VDD2.n27 3.49141
R1898 VDD2.n52 VDD2.n0 3.49141
R1899 VDD2.n72 VDD2.n71 2.84303
R1900 VDD2.n18 VDD2.n17 2.84303
R1901 VDD2.n103 VDD2.n102 2.71565
R1902 VDD2.n85 VDD2.n64 2.71565
R1903 VDD2.n31 VDD2.n10 2.71565
R1904 VDD2.n50 VDD2.n49 2.71565
R1905 VDD2.n99 VDD2.n55 1.93989
R1906 VDD2.n86 VDD2.n62 1.93989
R1907 VDD2.n32 VDD2.n8 1.93989
R1908 VDD2.n46 VDD2.n2 1.93989
R1909 VDD2.n98 VDD2.n57 1.16414
R1910 VDD2.n90 VDD2.n89 1.16414
R1911 VDD2.n37 VDD2.n35 1.16414
R1912 VDD2.n45 VDD2.n4 1.16414
R1913 VDD2 VDD2.n106 0.963862
R1914 VDD2.n95 VDD2.n94 0.388379
R1915 VDD2.n61 VDD2.n59 0.388379
R1916 VDD2.n36 VDD2.n6 0.388379
R1917 VDD2.n42 VDD2.n41 0.388379
R1918 VDD2.n104 VDD2.n54 0.155672
R1919 VDD2.n97 VDD2.n54 0.155672
R1920 VDD2.n97 VDD2.n96 0.155672
R1921 VDD2.n96 VDD2.n58 0.155672
R1922 VDD2.n88 VDD2.n58 0.155672
R1923 VDD2.n88 VDD2.n87 0.155672
R1924 VDD2.n87 VDD2.n63 0.155672
R1925 VDD2.n80 VDD2.n63 0.155672
R1926 VDD2.n80 VDD2.n79 0.155672
R1927 VDD2.n79 VDD2.n67 0.155672
R1928 VDD2.n72 VDD2.n67 0.155672
R1929 VDD2.n18 VDD2.n13 0.155672
R1930 VDD2.n25 VDD2.n13 0.155672
R1931 VDD2.n26 VDD2.n25 0.155672
R1932 VDD2.n26 VDD2.n9 0.155672
R1933 VDD2.n33 VDD2.n9 0.155672
R1934 VDD2.n34 VDD2.n33 0.155672
R1935 VDD2.n34 VDD2.n5 0.155672
R1936 VDD2.n43 VDD2.n5 0.155672
R1937 VDD2.n44 VDD2.n43 0.155672
R1938 VDD2.n44 VDD2.n1 0.155672
R1939 VDD2.n51 VDD2.n1 0.155672
C0 VDD2 VTAIL 4.9071f
C1 VP VDD1 2.72823f
C2 VN VDD1 0.148706f
C3 VDD2 VP 0.385802f
C4 VDD2 VN 2.49243f
C5 VTAIL VP 2.34533f
C6 VN VTAIL 2.3306f
C7 VN VP 5.69169f
C8 VDD2 VDD1 0.816701f
C9 VTAIL VDD1 4.84668f
C10 VDD2 B 4.5436f
C11 VDD1 B 7.39947f
C12 VTAIL B 7.152942f
C13 VN B 11.58884f
C14 VP B 7.84969f
C15 VDD2.n0 B 0.028704f
C16 VDD2.n1 B 0.02072f
C17 VDD2.n2 B 0.011134f
C18 VDD2.n3 B 0.026317f
C19 VDD2.n4 B 0.011789f
C20 VDD2.n5 B 0.02072f
C21 VDD2.n6 B 0.011461f
C22 VDD2.n7 B 0.026317f
C23 VDD2.n8 B 0.011789f
C24 VDD2.n9 B 0.02072f
C25 VDD2.n10 B 0.011134f
C26 VDD2.n11 B 0.026317f
C27 VDD2.n12 B 0.011789f
C28 VDD2.n13 B 0.02072f
C29 VDD2.n14 B 0.011134f
C30 VDD2.n15 B 0.019737f
C31 VDD2.n16 B 0.018604f
C32 VDD2.t0 B 0.044231f
C33 VDD2.n17 B 0.133879f
C34 VDD2.n18 B 0.865567f
C35 VDD2.n19 B 0.011134f
C36 VDD2.n20 B 0.011789f
C37 VDD2.n21 B 0.026317f
C38 VDD2.n22 B 0.026317f
C39 VDD2.n23 B 0.011789f
C40 VDD2.n24 B 0.011134f
C41 VDD2.n25 B 0.02072f
C42 VDD2.n26 B 0.02072f
C43 VDD2.n27 B 0.011134f
C44 VDD2.n28 B 0.011789f
C45 VDD2.n29 B 0.026317f
C46 VDD2.n30 B 0.026317f
C47 VDD2.n31 B 0.011789f
C48 VDD2.n32 B 0.011134f
C49 VDD2.n33 B 0.02072f
C50 VDD2.n34 B 0.02072f
C51 VDD2.n35 B 0.011134f
C52 VDD2.n36 B 0.011134f
C53 VDD2.n37 B 0.011789f
C54 VDD2.n38 B 0.026317f
C55 VDD2.n39 B 0.026317f
C56 VDD2.n40 B 0.026317f
C57 VDD2.n41 B 0.011461f
C58 VDD2.n42 B 0.011134f
C59 VDD2.n43 B 0.02072f
C60 VDD2.n44 B 0.02072f
C61 VDD2.n45 B 0.011134f
C62 VDD2.n46 B 0.011789f
C63 VDD2.n47 B 0.026317f
C64 VDD2.n48 B 0.05623f
C65 VDD2.n49 B 0.011789f
C66 VDD2.n50 B 0.011134f
C67 VDD2.n51 B 0.05044f
C68 VDD2.n52 B 0.610016f
C69 VDD2.n53 B 0.028704f
C70 VDD2.n54 B 0.02072f
C71 VDD2.n55 B 0.011134f
C72 VDD2.n56 B 0.026317f
C73 VDD2.n57 B 0.011789f
C74 VDD2.n58 B 0.02072f
C75 VDD2.n59 B 0.011461f
C76 VDD2.n60 B 0.026317f
C77 VDD2.n61 B 0.011134f
C78 VDD2.n62 B 0.011789f
C79 VDD2.n63 B 0.02072f
C80 VDD2.n64 B 0.011134f
C81 VDD2.n65 B 0.026317f
C82 VDD2.n66 B 0.011789f
C83 VDD2.n67 B 0.02072f
C84 VDD2.n68 B 0.011134f
C85 VDD2.n69 B 0.019737f
C86 VDD2.n70 B 0.018604f
C87 VDD2.t1 B 0.044231f
C88 VDD2.n71 B 0.133879f
C89 VDD2.n72 B 0.865567f
C90 VDD2.n73 B 0.011134f
C91 VDD2.n74 B 0.011789f
C92 VDD2.n75 B 0.026317f
C93 VDD2.n76 B 0.026317f
C94 VDD2.n77 B 0.011789f
C95 VDD2.n78 B 0.011134f
C96 VDD2.n79 B 0.02072f
C97 VDD2.n80 B 0.02072f
C98 VDD2.n81 B 0.011134f
C99 VDD2.n82 B 0.011789f
C100 VDD2.n83 B 0.026317f
C101 VDD2.n84 B 0.026317f
C102 VDD2.n85 B 0.011789f
C103 VDD2.n86 B 0.011134f
C104 VDD2.n87 B 0.02072f
C105 VDD2.n88 B 0.02072f
C106 VDD2.n89 B 0.011134f
C107 VDD2.n90 B 0.011789f
C108 VDD2.n91 B 0.026317f
C109 VDD2.n92 B 0.026317f
C110 VDD2.n93 B 0.026317f
C111 VDD2.n94 B 0.011461f
C112 VDD2.n95 B 0.011134f
C113 VDD2.n96 B 0.02072f
C114 VDD2.n97 B 0.02072f
C115 VDD2.n98 B 0.011134f
C116 VDD2.n99 B 0.011789f
C117 VDD2.n100 B 0.026317f
C118 VDD2.n101 B 0.05623f
C119 VDD2.n102 B 0.011789f
C120 VDD2.n103 B 0.011134f
C121 VDD2.n104 B 0.05044f
C122 VDD2.n105 B 0.04575f
C123 VDD2.n106 B 2.58148f
C124 VN.t1 B 3.04457f
C125 VN.t0 B 3.74205f
C126 VDD1.n0 B 0.028794f
C127 VDD1.n1 B 0.020785f
C128 VDD1.n2 B 0.011169f
C129 VDD1.n3 B 0.026399f
C130 VDD1.n4 B 0.011826f
C131 VDD1.n5 B 0.020785f
C132 VDD1.n6 B 0.011497f
C133 VDD1.n7 B 0.026399f
C134 VDD1.n8 B 0.011169f
C135 VDD1.n9 B 0.011826f
C136 VDD1.n10 B 0.020785f
C137 VDD1.n11 B 0.011169f
C138 VDD1.n12 B 0.026399f
C139 VDD1.n13 B 0.011826f
C140 VDD1.n14 B 0.020785f
C141 VDD1.n15 B 0.011169f
C142 VDD1.n16 B 0.019799f
C143 VDD1.n17 B 0.018662f
C144 VDD1.t0 B 0.04437f
C145 VDD1.n18 B 0.1343f
C146 VDD1.n19 B 0.868285f
C147 VDD1.n20 B 0.011169f
C148 VDD1.n21 B 0.011826f
C149 VDD1.n22 B 0.026399f
C150 VDD1.n23 B 0.026399f
C151 VDD1.n24 B 0.011826f
C152 VDD1.n25 B 0.011169f
C153 VDD1.n26 B 0.020785f
C154 VDD1.n27 B 0.020785f
C155 VDD1.n28 B 0.011169f
C156 VDD1.n29 B 0.011826f
C157 VDD1.n30 B 0.026399f
C158 VDD1.n31 B 0.026399f
C159 VDD1.n32 B 0.011826f
C160 VDD1.n33 B 0.011169f
C161 VDD1.n34 B 0.020785f
C162 VDD1.n35 B 0.020785f
C163 VDD1.n36 B 0.011169f
C164 VDD1.n37 B 0.011826f
C165 VDD1.n38 B 0.026399f
C166 VDD1.n39 B 0.026399f
C167 VDD1.n40 B 0.026399f
C168 VDD1.n41 B 0.011497f
C169 VDD1.n42 B 0.011169f
C170 VDD1.n43 B 0.020785f
C171 VDD1.n44 B 0.020785f
C172 VDD1.n45 B 0.011169f
C173 VDD1.n46 B 0.011826f
C174 VDD1.n47 B 0.026399f
C175 VDD1.n48 B 0.056406f
C176 VDD1.n49 B 0.011826f
C177 VDD1.n50 B 0.011169f
C178 VDD1.n51 B 0.050599f
C179 VDD1.n52 B 0.047874f
C180 VDD1.n53 B 0.028794f
C181 VDD1.n54 B 0.020785f
C182 VDD1.n55 B 0.011169f
C183 VDD1.n56 B 0.026399f
C184 VDD1.n57 B 0.011826f
C185 VDD1.n58 B 0.020785f
C186 VDD1.n59 B 0.011497f
C187 VDD1.n60 B 0.026399f
C188 VDD1.n61 B 0.011826f
C189 VDD1.n62 B 0.020785f
C190 VDD1.n63 B 0.011169f
C191 VDD1.n64 B 0.026399f
C192 VDD1.n65 B 0.011826f
C193 VDD1.n66 B 0.020785f
C194 VDD1.n67 B 0.011169f
C195 VDD1.n68 B 0.019799f
C196 VDD1.n69 B 0.018662f
C197 VDD1.t1 B 0.04437f
C198 VDD1.n70 B 0.1343f
C199 VDD1.n71 B 0.868285f
C200 VDD1.n72 B 0.011169f
C201 VDD1.n73 B 0.011826f
C202 VDD1.n74 B 0.026399f
C203 VDD1.n75 B 0.026399f
C204 VDD1.n76 B 0.011826f
C205 VDD1.n77 B 0.011169f
C206 VDD1.n78 B 0.020785f
C207 VDD1.n79 B 0.020785f
C208 VDD1.n80 B 0.011169f
C209 VDD1.n81 B 0.011826f
C210 VDD1.n82 B 0.026399f
C211 VDD1.n83 B 0.026399f
C212 VDD1.n84 B 0.011826f
C213 VDD1.n85 B 0.011169f
C214 VDD1.n86 B 0.020785f
C215 VDD1.n87 B 0.020785f
C216 VDD1.n88 B 0.011169f
C217 VDD1.n89 B 0.011169f
C218 VDD1.n90 B 0.011826f
C219 VDD1.n91 B 0.026399f
C220 VDD1.n92 B 0.026399f
C221 VDD1.n93 B 0.026399f
C222 VDD1.n94 B 0.011497f
C223 VDD1.n95 B 0.011169f
C224 VDD1.n96 B 0.020785f
C225 VDD1.n97 B 0.020785f
C226 VDD1.n98 B 0.011169f
C227 VDD1.n99 B 0.011826f
C228 VDD1.n100 B 0.026399f
C229 VDD1.n101 B 0.056406f
C230 VDD1.n102 B 0.011826f
C231 VDD1.n103 B 0.011169f
C232 VDD1.n104 B 0.050599f
C233 VDD1.n105 B 0.659949f
C234 VTAIL.n0 B 0.03006f
C235 VTAIL.n1 B 0.021698f
C236 VTAIL.n2 B 0.01166f
C237 VTAIL.n3 B 0.027559f
C238 VTAIL.n4 B 0.012346f
C239 VTAIL.n5 B 0.021698f
C240 VTAIL.n6 B 0.012003f
C241 VTAIL.n7 B 0.027559f
C242 VTAIL.n8 B 0.012346f
C243 VTAIL.n9 B 0.021698f
C244 VTAIL.n10 B 0.01166f
C245 VTAIL.n11 B 0.027559f
C246 VTAIL.n12 B 0.012346f
C247 VTAIL.n13 B 0.021698f
C248 VTAIL.n14 B 0.01166f
C249 VTAIL.n15 B 0.020669f
C250 VTAIL.n16 B 0.019482f
C251 VTAIL.t2 B 0.04632f
C252 VTAIL.n17 B 0.140201f
C253 VTAIL.n18 B 0.906437f
C254 VTAIL.n19 B 0.01166f
C255 VTAIL.n20 B 0.012346f
C256 VTAIL.n21 B 0.027559f
C257 VTAIL.n22 B 0.027559f
C258 VTAIL.n23 B 0.012346f
C259 VTAIL.n24 B 0.01166f
C260 VTAIL.n25 B 0.021698f
C261 VTAIL.n26 B 0.021698f
C262 VTAIL.n27 B 0.01166f
C263 VTAIL.n28 B 0.012346f
C264 VTAIL.n29 B 0.027559f
C265 VTAIL.n30 B 0.027559f
C266 VTAIL.n31 B 0.012346f
C267 VTAIL.n32 B 0.01166f
C268 VTAIL.n33 B 0.021698f
C269 VTAIL.n34 B 0.021698f
C270 VTAIL.n35 B 0.01166f
C271 VTAIL.n36 B 0.01166f
C272 VTAIL.n37 B 0.012346f
C273 VTAIL.n38 B 0.027559f
C274 VTAIL.n39 B 0.027559f
C275 VTAIL.n40 B 0.027559f
C276 VTAIL.n41 B 0.012003f
C277 VTAIL.n42 B 0.01166f
C278 VTAIL.n43 B 0.021698f
C279 VTAIL.n44 B 0.021698f
C280 VTAIL.n45 B 0.01166f
C281 VTAIL.n46 B 0.012346f
C282 VTAIL.n47 B 0.027559f
C283 VTAIL.n48 B 0.058884f
C284 VTAIL.n49 B 0.012346f
C285 VTAIL.n50 B 0.01166f
C286 VTAIL.n51 B 0.052822f
C287 VTAIL.n52 B 0.032948f
C288 VTAIL.n53 B 1.52702f
C289 VTAIL.n54 B 0.03006f
C290 VTAIL.n55 B 0.021698f
C291 VTAIL.n56 B 0.01166f
C292 VTAIL.n57 B 0.027559f
C293 VTAIL.n58 B 0.012346f
C294 VTAIL.n59 B 0.021698f
C295 VTAIL.n60 B 0.012003f
C296 VTAIL.n61 B 0.027559f
C297 VTAIL.n62 B 0.01166f
C298 VTAIL.n63 B 0.012346f
C299 VTAIL.n64 B 0.021698f
C300 VTAIL.n65 B 0.01166f
C301 VTAIL.n66 B 0.027559f
C302 VTAIL.n67 B 0.012346f
C303 VTAIL.n68 B 0.021698f
C304 VTAIL.n69 B 0.01166f
C305 VTAIL.n70 B 0.020669f
C306 VTAIL.n71 B 0.019482f
C307 VTAIL.t0 B 0.04632f
C308 VTAIL.n72 B 0.140201f
C309 VTAIL.n73 B 0.906437f
C310 VTAIL.n74 B 0.01166f
C311 VTAIL.n75 B 0.012346f
C312 VTAIL.n76 B 0.027559f
C313 VTAIL.n77 B 0.027559f
C314 VTAIL.n78 B 0.012346f
C315 VTAIL.n79 B 0.01166f
C316 VTAIL.n80 B 0.021698f
C317 VTAIL.n81 B 0.021698f
C318 VTAIL.n82 B 0.01166f
C319 VTAIL.n83 B 0.012346f
C320 VTAIL.n84 B 0.027559f
C321 VTAIL.n85 B 0.027559f
C322 VTAIL.n86 B 0.012346f
C323 VTAIL.n87 B 0.01166f
C324 VTAIL.n88 B 0.021698f
C325 VTAIL.n89 B 0.021698f
C326 VTAIL.n90 B 0.01166f
C327 VTAIL.n91 B 0.012346f
C328 VTAIL.n92 B 0.027559f
C329 VTAIL.n93 B 0.027559f
C330 VTAIL.n94 B 0.027559f
C331 VTAIL.n95 B 0.012003f
C332 VTAIL.n96 B 0.01166f
C333 VTAIL.n97 B 0.021698f
C334 VTAIL.n98 B 0.021698f
C335 VTAIL.n99 B 0.01166f
C336 VTAIL.n100 B 0.012346f
C337 VTAIL.n101 B 0.027559f
C338 VTAIL.n102 B 0.058884f
C339 VTAIL.n103 B 0.012346f
C340 VTAIL.n104 B 0.01166f
C341 VTAIL.n105 B 0.052822f
C342 VTAIL.n106 B 0.032948f
C343 VTAIL.n107 B 1.58624f
C344 VTAIL.n108 B 0.03006f
C345 VTAIL.n109 B 0.021698f
C346 VTAIL.n110 B 0.01166f
C347 VTAIL.n111 B 0.027559f
C348 VTAIL.n112 B 0.012346f
C349 VTAIL.n113 B 0.021698f
C350 VTAIL.n114 B 0.012003f
C351 VTAIL.n115 B 0.027559f
C352 VTAIL.n116 B 0.01166f
C353 VTAIL.n117 B 0.012346f
C354 VTAIL.n118 B 0.021698f
C355 VTAIL.n119 B 0.01166f
C356 VTAIL.n120 B 0.027559f
C357 VTAIL.n121 B 0.012346f
C358 VTAIL.n122 B 0.021698f
C359 VTAIL.n123 B 0.01166f
C360 VTAIL.n124 B 0.020669f
C361 VTAIL.n125 B 0.019482f
C362 VTAIL.t3 B 0.04632f
C363 VTAIL.n126 B 0.140201f
C364 VTAIL.n127 B 0.906437f
C365 VTAIL.n128 B 0.01166f
C366 VTAIL.n129 B 0.012346f
C367 VTAIL.n130 B 0.027559f
C368 VTAIL.n131 B 0.027559f
C369 VTAIL.n132 B 0.012346f
C370 VTAIL.n133 B 0.01166f
C371 VTAIL.n134 B 0.021698f
C372 VTAIL.n135 B 0.021698f
C373 VTAIL.n136 B 0.01166f
C374 VTAIL.n137 B 0.012346f
C375 VTAIL.n138 B 0.027559f
C376 VTAIL.n139 B 0.027559f
C377 VTAIL.n140 B 0.012346f
C378 VTAIL.n141 B 0.01166f
C379 VTAIL.n142 B 0.021698f
C380 VTAIL.n143 B 0.021698f
C381 VTAIL.n144 B 0.01166f
C382 VTAIL.n145 B 0.012346f
C383 VTAIL.n146 B 0.027559f
C384 VTAIL.n147 B 0.027559f
C385 VTAIL.n148 B 0.027559f
C386 VTAIL.n149 B 0.012003f
C387 VTAIL.n150 B 0.01166f
C388 VTAIL.n151 B 0.021698f
C389 VTAIL.n152 B 0.021698f
C390 VTAIL.n153 B 0.01166f
C391 VTAIL.n154 B 0.012346f
C392 VTAIL.n155 B 0.027559f
C393 VTAIL.n156 B 0.058884f
C394 VTAIL.n157 B 0.012346f
C395 VTAIL.n158 B 0.01166f
C396 VTAIL.n159 B 0.052822f
C397 VTAIL.n160 B 0.032948f
C398 VTAIL.n161 B 1.33309f
C399 VTAIL.n162 B 0.03006f
C400 VTAIL.n163 B 0.021698f
C401 VTAIL.n164 B 0.01166f
C402 VTAIL.n165 B 0.027559f
C403 VTAIL.n166 B 0.012346f
C404 VTAIL.n167 B 0.021698f
C405 VTAIL.n168 B 0.012003f
C406 VTAIL.n169 B 0.027559f
C407 VTAIL.n170 B 0.012346f
C408 VTAIL.n171 B 0.021698f
C409 VTAIL.n172 B 0.01166f
C410 VTAIL.n173 B 0.027559f
C411 VTAIL.n174 B 0.012346f
C412 VTAIL.n175 B 0.021698f
C413 VTAIL.n176 B 0.01166f
C414 VTAIL.n177 B 0.020669f
C415 VTAIL.n178 B 0.019482f
C416 VTAIL.t1 B 0.04632f
C417 VTAIL.n179 B 0.140201f
C418 VTAIL.n180 B 0.906437f
C419 VTAIL.n181 B 0.01166f
C420 VTAIL.n182 B 0.012346f
C421 VTAIL.n183 B 0.027559f
C422 VTAIL.n184 B 0.027559f
C423 VTAIL.n185 B 0.012346f
C424 VTAIL.n186 B 0.01166f
C425 VTAIL.n187 B 0.021698f
C426 VTAIL.n188 B 0.021698f
C427 VTAIL.n189 B 0.01166f
C428 VTAIL.n190 B 0.012346f
C429 VTAIL.n191 B 0.027559f
C430 VTAIL.n192 B 0.027559f
C431 VTAIL.n193 B 0.012346f
C432 VTAIL.n194 B 0.01166f
C433 VTAIL.n195 B 0.021698f
C434 VTAIL.n196 B 0.021698f
C435 VTAIL.n197 B 0.01166f
C436 VTAIL.n198 B 0.01166f
C437 VTAIL.n199 B 0.012346f
C438 VTAIL.n200 B 0.027559f
C439 VTAIL.n201 B 0.027559f
C440 VTAIL.n202 B 0.027559f
C441 VTAIL.n203 B 0.012003f
C442 VTAIL.n204 B 0.01166f
C443 VTAIL.n205 B 0.021698f
C444 VTAIL.n206 B 0.021698f
C445 VTAIL.n207 B 0.01166f
C446 VTAIL.n208 B 0.012346f
C447 VTAIL.n209 B 0.027559f
C448 VTAIL.n210 B 0.058884f
C449 VTAIL.n211 B 0.012346f
C450 VTAIL.n212 B 0.01166f
C451 VTAIL.n213 B 0.052822f
C452 VTAIL.n214 B 0.032948f
C453 VTAIL.n215 B 1.23289f
C454 VP.t1 B 3.82795f
C455 VP.t0 B 3.10692f
C456 VP.n0 B 3.65429f
.ends

