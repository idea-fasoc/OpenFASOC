* NGSPICE file created from diff_pair_sample_1245.ext - technology: sky130A

.subckt diff_pair_sample_1245 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=2.4816 ps=15.37 w=15.04 l=2.53
X1 VTAIL.t13 VP.t1 VDD1.t8 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X2 VDD1.t7 VP.t2 VTAIL.t14 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X3 B.t11 B.t9 B.t10 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=0 ps=0 w=15.04 l=2.53
X4 VTAIL.t18 VN.t0 VDD2.t9 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X5 VDD2.t8 VN.t1 VTAIL.t19 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X6 VTAIL.t2 VN.t2 VDD2.t7 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X7 VTAIL.t15 VP.t3 VDD1.t6 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X8 VTAIL.t16 VP.t4 VDD1.t5 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X9 VDD2.t6 VN.t3 VTAIL.t6 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=2.4816 ps=15.37 w=15.04 l=2.53
X10 VDD2.t5 VN.t4 VTAIL.t5 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=5.8656 ps=30.86 w=15.04 l=2.53
X11 VDD1.t4 VP.t5 VTAIL.t17 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X12 VDD2.t4 VN.t5 VTAIL.t4 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=5.8656 ps=30.86 w=15.04 l=2.53
X13 B.t8 B.t6 B.t7 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=0 ps=0 w=15.04 l=2.53
X14 VDD1.t3 VP.t6 VTAIL.t8 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=5.8656 ps=30.86 w=15.04 l=2.53
X15 VDD1.t2 VP.t7 VTAIL.t9 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=5.8656 ps=30.86 w=15.04 l=2.53
X16 VDD2.t3 VN.t6 VTAIL.t3 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=2.4816 ps=15.37 w=15.04 l=2.53
X17 B.t5 B.t3 B.t4 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=0 ps=0 w=15.04 l=2.53
X18 VTAIL.t1 VN.t7 VDD2.t2 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X19 VTAIL.t7 VN.t8 VDD2.t1 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X20 VTAIL.t10 VP.t8 VDD1.t1 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
X21 VDD1.t0 VP.t9 VTAIL.t11 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=2.4816 ps=15.37 w=15.04 l=2.53
X22 B.t2 B.t0 B.t1 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=5.8656 pd=30.86 as=0 ps=0 w=15.04 l=2.53
X23 VDD2.t0 VN.t9 VTAIL.t0 w_n4402_n3976# sky130_fd_pr__pfet_01v8 ad=2.4816 pd=15.37 as=2.4816 ps=15.37 w=15.04 l=2.53
R0 VP.n23 VP.t9 177.169
R1 VP.n25 VP.n24 161.3
R2 VP.n26 VP.n21 161.3
R3 VP.n28 VP.n27 161.3
R4 VP.n29 VP.n20 161.3
R5 VP.n31 VP.n30 161.3
R6 VP.n32 VP.n19 161.3
R7 VP.n34 VP.n33 161.3
R8 VP.n35 VP.n18 161.3
R9 VP.n37 VP.n36 161.3
R10 VP.n38 VP.n17 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n43 VP.n15 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n14 161.3
R16 VP.n48 VP.n47 161.3
R17 VP.n49 VP.n13 161.3
R18 VP.n88 VP.n0 161.3
R19 VP.n87 VP.n86 161.3
R20 VP.n85 VP.n1 161.3
R21 VP.n84 VP.n83 161.3
R22 VP.n82 VP.n2 161.3
R23 VP.n81 VP.n80 161.3
R24 VP.n79 VP.n78 161.3
R25 VP.n77 VP.n4 161.3
R26 VP.n76 VP.n75 161.3
R27 VP.n74 VP.n5 161.3
R28 VP.n73 VP.n72 161.3
R29 VP.n71 VP.n6 161.3
R30 VP.n70 VP.n69 161.3
R31 VP.n68 VP.n7 161.3
R32 VP.n67 VP.n66 161.3
R33 VP.n65 VP.n8 161.3
R34 VP.n64 VP.n63 161.3
R35 VP.n62 VP.n61 161.3
R36 VP.n60 VP.n10 161.3
R37 VP.n59 VP.n58 161.3
R38 VP.n57 VP.n11 161.3
R39 VP.n56 VP.n55 161.3
R40 VP.n54 VP.n12 161.3
R41 VP.n71 VP.t5 143.267
R42 VP.n53 VP.t0 143.267
R43 VP.n9 VP.t8 143.267
R44 VP.n3 VP.t3 143.267
R45 VP.n89 VP.t7 143.267
R46 VP.n32 VP.t2 143.267
R47 VP.n50 VP.t6 143.267
R48 VP.n16 VP.t4 143.267
R49 VP.n22 VP.t1 143.267
R50 VP.n53 VP.n52 100.088
R51 VP.n90 VP.n89 100.088
R52 VP.n51 VP.n50 100.088
R53 VP.n59 VP.n11 56.5617
R54 VP.n83 VP.n1 56.5617
R55 VP.n44 VP.n14 56.5617
R56 VP.n52 VP.n51 55.0527
R57 VP.n23 VP.n22 55.0245
R58 VP.n66 VP.n7 47.3584
R59 VP.n76 VP.n5 47.3584
R60 VP.n37 VP.n18 47.3584
R61 VP.n27 VP.n20 47.3584
R62 VP.n66 VP.n65 33.7956
R63 VP.n77 VP.n76 33.7956
R64 VP.n38 VP.n37 33.7956
R65 VP.n27 VP.n26 33.7956
R66 VP.n55 VP.n54 24.5923
R67 VP.n55 VP.n11 24.5923
R68 VP.n60 VP.n59 24.5923
R69 VP.n61 VP.n60 24.5923
R70 VP.n65 VP.n64 24.5923
R71 VP.n70 VP.n7 24.5923
R72 VP.n71 VP.n70 24.5923
R73 VP.n72 VP.n71 24.5923
R74 VP.n72 VP.n5 24.5923
R75 VP.n78 VP.n77 24.5923
R76 VP.n82 VP.n81 24.5923
R77 VP.n83 VP.n82 24.5923
R78 VP.n87 VP.n1 24.5923
R79 VP.n88 VP.n87 24.5923
R80 VP.n48 VP.n14 24.5923
R81 VP.n49 VP.n48 24.5923
R82 VP.n39 VP.n38 24.5923
R83 VP.n43 VP.n42 24.5923
R84 VP.n44 VP.n43 24.5923
R85 VP.n31 VP.n20 24.5923
R86 VP.n32 VP.n31 24.5923
R87 VP.n33 VP.n32 24.5923
R88 VP.n33 VP.n18 24.5923
R89 VP.n26 VP.n25 24.5923
R90 VP.n64 VP.n9 17.7066
R91 VP.n78 VP.n3 17.7066
R92 VP.n39 VP.n16 17.7066
R93 VP.n25 VP.n22 17.7066
R94 VP.n54 VP.n53 10.8209
R95 VP.n89 VP.n88 10.8209
R96 VP.n50 VP.n49 10.8209
R97 VP.n61 VP.n9 6.88621
R98 VP.n81 VP.n3 6.88621
R99 VP.n42 VP.n16 6.88621
R100 VP.n24 VP.n23 6.78213
R101 VP.n51 VP.n13 0.278335
R102 VP.n52 VP.n12 0.278335
R103 VP.n90 VP.n0 0.278335
R104 VP.n24 VP.n21 0.189894
R105 VP.n28 VP.n21 0.189894
R106 VP.n29 VP.n28 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n30 VP.n19 0.189894
R109 VP.n34 VP.n19 0.189894
R110 VP.n35 VP.n34 0.189894
R111 VP.n36 VP.n35 0.189894
R112 VP.n36 VP.n17 0.189894
R113 VP.n40 VP.n17 0.189894
R114 VP.n41 VP.n40 0.189894
R115 VP.n41 VP.n15 0.189894
R116 VP.n45 VP.n15 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n13 0.189894
R120 VP.n56 VP.n12 0.189894
R121 VP.n57 VP.n56 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n58 VP.n10 0.189894
R124 VP.n62 VP.n10 0.189894
R125 VP.n63 VP.n62 0.189894
R126 VP.n63 VP.n8 0.189894
R127 VP.n67 VP.n8 0.189894
R128 VP.n68 VP.n67 0.189894
R129 VP.n69 VP.n68 0.189894
R130 VP.n69 VP.n6 0.189894
R131 VP.n73 VP.n6 0.189894
R132 VP.n74 VP.n73 0.189894
R133 VP.n75 VP.n74 0.189894
R134 VP.n75 VP.n4 0.189894
R135 VP.n79 VP.n4 0.189894
R136 VP.n80 VP.n79 0.189894
R137 VP.n80 VP.n2 0.189894
R138 VP.n84 VP.n2 0.189894
R139 VP.n85 VP.n84 0.189894
R140 VP.n86 VP.n85 0.189894
R141 VP.n86 VP.n0 0.189894
R142 VP VP.n90 0.153485
R143 VTAIL.n11 VTAIL.t4 56.7634
R144 VTAIL.n17 VTAIL.t5 56.7631
R145 VTAIL.n2 VTAIL.t9 56.7631
R146 VTAIL.n16 VTAIL.t8 56.7631
R147 VTAIL.n15 VTAIL.n14 54.6021
R148 VTAIL.n13 VTAIL.n12 54.6021
R149 VTAIL.n10 VTAIL.n9 54.6021
R150 VTAIL.n8 VTAIL.n7 54.6021
R151 VTAIL.n19 VTAIL.n18 54.6019
R152 VTAIL.n1 VTAIL.n0 54.6019
R153 VTAIL.n4 VTAIL.n3 54.6019
R154 VTAIL.n6 VTAIL.n5 54.6019
R155 VTAIL.n8 VTAIL.n6 30.2634
R156 VTAIL.n17 VTAIL.n16 27.7979
R157 VTAIL.n10 VTAIL.n8 2.46602
R158 VTAIL.n11 VTAIL.n10 2.46602
R159 VTAIL.n15 VTAIL.n13 2.46602
R160 VTAIL.n16 VTAIL.n15 2.46602
R161 VTAIL.n6 VTAIL.n4 2.46602
R162 VTAIL.n4 VTAIL.n2 2.46602
R163 VTAIL.n19 VTAIL.n17 2.46602
R164 VTAIL.n18 VTAIL.t19 2.16174
R165 VTAIL.n18 VTAIL.t1 2.16174
R166 VTAIL.n0 VTAIL.t3 2.16174
R167 VTAIL.n0 VTAIL.t2 2.16174
R168 VTAIL.n3 VTAIL.t17 2.16174
R169 VTAIL.n3 VTAIL.t15 2.16174
R170 VTAIL.n5 VTAIL.t12 2.16174
R171 VTAIL.n5 VTAIL.t10 2.16174
R172 VTAIL.n14 VTAIL.t14 2.16174
R173 VTAIL.n14 VTAIL.t16 2.16174
R174 VTAIL.n12 VTAIL.t11 2.16174
R175 VTAIL.n12 VTAIL.t13 2.16174
R176 VTAIL.n9 VTAIL.t0 2.16174
R177 VTAIL.n9 VTAIL.t7 2.16174
R178 VTAIL.n7 VTAIL.t6 2.16174
R179 VTAIL.n7 VTAIL.t18 2.16174
R180 VTAIL VTAIL.n1 1.90783
R181 VTAIL.n13 VTAIL.n11 1.70309
R182 VTAIL.n2 VTAIL.n1 1.70309
R183 VTAIL VTAIL.n19 0.55869
R184 VDD1.n1 VDD1.t0 75.9077
R185 VDD1.n3 VDD1.t9 75.9074
R186 VDD1.n5 VDD1.n4 73.0745
R187 VDD1.n1 VDD1.n0 71.2809
R188 VDD1.n7 VDD1.n6 71.2807
R189 VDD1.n3 VDD1.n2 71.2807
R190 VDD1.n7 VDD1.n5 50.2078
R191 VDD1.n6 VDD1.t5 2.16174
R192 VDD1.n6 VDD1.t3 2.16174
R193 VDD1.n0 VDD1.t8 2.16174
R194 VDD1.n0 VDD1.t7 2.16174
R195 VDD1.n4 VDD1.t6 2.16174
R196 VDD1.n4 VDD1.t2 2.16174
R197 VDD1.n2 VDD1.t1 2.16174
R198 VDD1.n2 VDD1.t4 2.16174
R199 VDD1 VDD1.n7 1.79145
R200 VDD1 VDD1.n1 0.675069
R201 VDD1.n5 VDD1.n3 0.561533
R202 B.n492 B.n491 585
R203 B.n490 B.n151 585
R204 B.n489 B.n488 585
R205 B.n487 B.n152 585
R206 B.n486 B.n485 585
R207 B.n484 B.n153 585
R208 B.n483 B.n482 585
R209 B.n481 B.n154 585
R210 B.n480 B.n479 585
R211 B.n478 B.n155 585
R212 B.n477 B.n476 585
R213 B.n475 B.n156 585
R214 B.n474 B.n473 585
R215 B.n472 B.n157 585
R216 B.n471 B.n470 585
R217 B.n469 B.n158 585
R218 B.n468 B.n467 585
R219 B.n466 B.n159 585
R220 B.n465 B.n464 585
R221 B.n463 B.n160 585
R222 B.n462 B.n461 585
R223 B.n460 B.n161 585
R224 B.n459 B.n458 585
R225 B.n457 B.n162 585
R226 B.n456 B.n455 585
R227 B.n454 B.n163 585
R228 B.n453 B.n452 585
R229 B.n451 B.n164 585
R230 B.n450 B.n449 585
R231 B.n448 B.n165 585
R232 B.n447 B.n446 585
R233 B.n445 B.n166 585
R234 B.n444 B.n443 585
R235 B.n442 B.n167 585
R236 B.n441 B.n440 585
R237 B.n439 B.n168 585
R238 B.n438 B.n437 585
R239 B.n436 B.n169 585
R240 B.n435 B.n434 585
R241 B.n433 B.n170 585
R242 B.n432 B.n431 585
R243 B.n430 B.n171 585
R244 B.n429 B.n428 585
R245 B.n427 B.n172 585
R246 B.n426 B.n425 585
R247 B.n424 B.n173 585
R248 B.n423 B.n422 585
R249 B.n421 B.n174 585
R250 B.n420 B.n419 585
R251 B.n418 B.n175 585
R252 B.n417 B.n416 585
R253 B.n414 B.n176 585
R254 B.n413 B.n412 585
R255 B.n411 B.n179 585
R256 B.n410 B.n409 585
R257 B.n408 B.n180 585
R258 B.n407 B.n406 585
R259 B.n405 B.n181 585
R260 B.n404 B.n403 585
R261 B.n402 B.n182 585
R262 B.n400 B.n399 585
R263 B.n398 B.n185 585
R264 B.n397 B.n396 585
R265 B.n395 B.n186 585
R266 B.n394 B.n393 585
R267 B.n392 B.n187 585
R268 B.n391 B.n390 585
R269 B.n389 B.n188 585
R270 B.n388 B.n387 585
R271 B.n386 B.n189 585
R272 B.n385 B.n384 585
R273 B.n383 B.n190 585
R274 B.n382 B.n381 585
R275 B.n380 B.n191 585
R276 B.n379 B.n378 585
R277 B.n377 B.n192 585
R278 B.n376 B.n375 585
R279 B.n374 B.n193 585
R280 B.n373 B.n372 585
R281 B.n371 B.n194 585
R282 B.n370 B.n369 585
R283 B.n368 B.n195 585
R284 B.n367 B.n366 585
R285 B.n365 B.n196 585
R286 B.n364 B.n363 585
R287 B.n362 B.n197 585
R288 B.n361 B.n360 585
R289 B.n359 B.n198 585
R290 B.n358 B.n357 585
R291 B.n356 B.n199 585
R292 B.n355 B.n354 585
R293 B.n353 B.n200 585
R294 B.n352 B.n351 585
R295 B.n350 B.n201 585
R296 B.n349 B.n348 585
R297 B.n347 B.n202 585
R298 B.n346 B.n345 585
R299 B.n344 B.n203 585
R300 B.n343 B.n342 585
R301 B.n341 B.n204 585
R302 B.n340 B.n339 585
R303 B.n338 B.n205 585
R304 B.n337 B.n336 585
R305 B.n335 B.n206 585
R306 B.n334 B.n333 585
R307 B.n332 B.n207 585
R308 B.n331 B.n330 585
R309 B.n329 B.n208 585
R310 B.n328 B.n327 585
R311 B.n326 B.n209 585
R312 B.n325 B.n324 585
R313 B.n493 B.n150 585
R314 B.n495 B.n494 585
R315 B.n496 B.n149 585
R316 B.n498 B.n497 585
R317 B.n499 B.n148 585
R318 B.n501 B.n500 585
R319 B.n502 B.n147 585
R320 B.n504 B.n503 585
R321 B.n505 B.n146 585
R322 B.n507 B.n506 585
R323 B.n508 B.n145 585
R324 B.n510 B.n509 585
R325 B.n511 B.n144 585
R326 B.n513 B.n512 585
R327 B.n514 B.n143 585
R328 B.n516 B.n515 585
R329 B.n517 B.n142 585
R330 B.n519 B.n518 585
R331 B.n520 B.n141 585
R332 B.n522 B.n521 585
R333 B.n523 B.n140 585
R334 B.n525 B.n524 585
R335 B.n526 B.n139 585
R336 B.n528 B.n527 585
R337 B.n529 B.n138 585
R338 B.n531 B.n530 585
R339 B.n532 B.n137 585
R340 B.n534 B.n533 585
R341 B.n535 B.n136 585
R342 B.n537 B.n536 585
R343 B.n538 B.n135 585
R344 B.n540 B.n539 585
R345 B.n541 B.n134 585
R346 B.n543 B.n542 585
R347 B.n544 B.n133 585
R348 B.n546 B.n545 585
R349 B.n547 B.n132 585
R350 B.n549 B.n548 585
R351 B.n550 B.n131 585
R352 B.n552 B.n551 585
R353 B.n553 B.n130 585
R354 B.n555 B.n554 585
R355 B.n556 B.n129 585
R356 B.n558 B.n557 585
R357 B.n559 B.n128 585
R358 B.n561 B.n560 585
R359 B.n562 B.n127 585
R360 B.n564 B.n563 585
R361 B.n565 B.n126 585
R362 B.n567 B.n566 585
R363 B.n568 B.n125 585
R364 B.n570 B.n569 585
R365 B.n571 B.n124 585
R366 B.n573 B.n572 585
R367 B.n574 B.n123 585
R368 B.n576 B.n575 585
R369 B.n577 B.n122 585
R370 B.n579 B.n578 585
R371 B.n580 B.n121 585
R372 B.n582 B.n581 585
R373 B.n583 B.n120 585
R374 B.n585 B.n584 585
R375 B.n586 B.n119 585
R376 B.n588 B.n587 585
R377 B.n589 B.n118 585
R378 B.n591 B.n590 585
R379 B.n592 B.n117 585
R380 B.n594 B.n593 585
R381 B.n595 B.n116 585
R382 B.n597 B.n596 585
R383 B.n598 B.n115 585
R384 B.n600 B.n599 585
R385 B.n601 B.n114 585
R386 B.n603 B.n602 585
R387 B.n604 B.n113 585
R388 B.n606 B.n605 585
R389 B.n607 B.n112 585
R390 B.n609 B.n608 585
R391 B.n610 B.n111 585
R392 B.n612 B.n611 585
R393 B.n613 B.n110 585
R394 B.n615 B.n614 585
R395 B.n616 B.n109 585
R396 B.n618 B.n617 585
R397 B.n619 B.n108 585
R398 B.n621 B.n620 585
R399 B.n622 B.n107 585
R400 B.n624 B.n623 585
R401 B.n625 B.n106 585
R402 B.n627 B.n626 585
R403 B.n628 B.n105 585
R404 B.n630 B.n629 585
R405 B.n631 B.n104 585
R406 B.n633 B.n632 585
R407 B.n634 B.n103 585
R408 B.n636 B.n635 585
R409 B.n637 B.n102 585
R410 B.n639 B.n638 585
R411 B.n640 B.n101 585
R412 B.n642 B.n641 585
R413 B.n643 B.n100 585
R414 B.n645 B.n644 585
R415 B.n646 B.n99 585
R416 B.n648 B.n647 585
R417 B.n649 B.n98 585
R418 B.n651 B.n650 585
R419 B.n652 B.n97 585
R420 B.n654 B.n653 585
R421 B.n655 B.n96 585
R422 B.n657 B.n656 585
R423 B.n658 B.n95 585
R424 B.n660 B.n659 585
R425 B.n661 B.n94 585
R426 B.n663 B.n662 585
R427 B.n664 B.n93 585
R428 B.n666 B.n665 585
R429 B.n667 B.n92 585
R430 B.n669 B.n668 585
R431 B.n836 B.n31 585
R432 B.n835 B.n834 585
R433 B.n833 B.n32 585
R434 B.n832 B.n831 585
R435 B.n830 B.n33 585
R436 B.n829 B.n828 585
R437 B.n827 B.n34 585
R438 B.n826 B.n825 585
R439 B.n824 B.n35 585
R440 B.n823 B.n822 585
R441 B.n821 B.n36 585
R442 B.n820 B.n819 585
R443 B.n818 B.n37 585
R444 B.n817 B.n816 585
R445 B.n815 B.n38 585
R446 B.n814 B.n813 585
R447 B.n812 B.n39 585
R448 B.n811 B.n810 585
R449 B.n809 B.n40 585
R450 B.n808 B.n807 585
R451 B.n806 B.n41 585
R452 B.n805 B.n804 585
R453 B.n803 B.n42 585
R454 B.n802 B.n801 585
R455 B.n800 B.n43 585
R456 B.n799 B.n798 585
R457 B.n797 B.n44 585
R458 B.n796 B.n795 585
R459 B.n794 B.n45 585
R460 B.n793 B.n792 585
R461 B.n791 B.n46 585
R462 B.n790 B.n789 585
R463 B.n788 B.n47 585
R464 B.n787 B.n786 585
R465 B.n785 B.n48 585
R466 B.n784 B.n783 585
R467 B.n782 B.n49 585
R468 B.n781 B.n780 585
R469 B.n779 B.n50 585
R470 B.n778 B.n777 585
R471 B.n776 B.n51 585
R472 B.n775 B.n774 585
R473 B.n773 B.n52 585
R474 B.n772 B.n771 585
R475 B.n770 B.n53 585
R476 B.n769 B.n768 585
R477 B.n767 B.n54 585
R478 B.n766 B.n765 585
R479 B.n764 B.n55 585
R480 B.n763 B.n762 585
R481 B.n761 B.n56 585
R482 B.n760 B.n759 585
R483 B.n758 B.n57 585
R484 B.n757 B.n756 585
R485 B.n755 B.n61 585
R486 B.n754 B.n753 585
R487 B.n752 B.n62 585
R488 B.n751 B.n750 585
R489 B.n749 B.n63 585
R490 B.n748 B.n747 585
R491 B.n745 B.n64 585
R492 B.n744 B.n743 585
R493 B.n742 B.n67 585
R494 B.n741 B.n740 585
R495 B.n739 B.n68 585
R496 B.n738 B.n737 585
R497 B.n736 B.n69 585
R498 B.n735 B.n734 585
R499 B.n733 B.n70 585
R500 B.n732 B.n731 585
R501 B.n730 B.n71 585
R502 B.n729 B.n728 585
R503 B.n727 B.n72 585
R504 B.n726 B.n725 585
R505 B.n724 B.n73 585
R506 B.n723 B.n722 585
R507 B.n721 B.n74 585
R508 B.n720 B.n719 585
R509 B.n718 B.n75 585
R510 B.n717 B.n716 585
R511 B.n715 B.n76 585
R512 B.n714 B.n713 585
R513 B.n712 B.n77 585
R514 B.n711 B.n710 585
R515 B.n709 B.n78 585
R516 B.n708 B.n707 585
R517 B.n706 B.n79 585
R518 B.n705 B.n704 585
R519 B.n703 B.n80 585
R520 B.n702 B.n701 585
R521 B.n700 B.n81 585
R522 B.n699 B.n698 585
R523 B.n697 B.n82 585
R524 B.n696 B.n695 585
R525 B.n694 B.n83 585
R526 B.n693 B.n692 585
R527 B.n691 B.n84 585
R528 B.n690 B.n689 585
R529 B.n688 B.n85 585
R530 B.n687 B.n686 585
R531 B.n685 B.n86 585
R532 B.n684 B.n683 585
R533 B.n682 B.n87 585
R534 B.n681 B.n680 585
R535 B.n679 B.n88 585
R536 B.n678 B.n677 585
R537 B.n676 B.n89 585
R538 B.n675 B.n674 585
R539 B.n673 B.n90 585
R540 B.n672 B.n671 585
R541 B.n670 B.n91 585
R542 B.n838 B.n837 585
R543 B.n839 B.n30 585
R544 B.n841 B.n840 585
R545 B.n842 B.n29 585
R546 B.n844 B.n843 585
R547 B.n845 B.n28 585
R548 B.n847 B.n846 585
R549 B.n848 B.n27 585
R550 B.n850 B.n849 585
R551 B.n851 B.n26 585
R552 B.n853 B.n852 585
R553 B.n854 B.n25 585
R554 B.n856 B.n855 585
R555 B.n857 B.n24 585
R556 B.n859 B.n858 585
R557 B.n860 B.n23 585
R558 B.n862 B.n861 585
R559 B.n863 B.n22 585
R560 B.n865 B.n864 585
R561 B.n866 B.n21 585
R562 B.n868 B.n867 585
R563 B.n869 B.n20 585
R564 B.n871 B.n870 585
R565 B.n872 B.n19 585
R566 B.n874 B.n873 585
R567 B.n875 B.n18 585
R568 B.n877 B.n876 585
R569 B.n878 B.n17 585
R570 B.n880 B.n879 585
R571 B.n881 B.n16 585
R572 B.n883 B.n882 585
R573 B.n884 B.n15 585
R574 B.n886 B.n885 585
R575 B.n887 B.n14 585
R576 B.n889 B.n888 585
R577 B.n890 B.n13 585
R578 B.n892 B.n891 585
R579 B.n893 B.n12 585
R580 B.n895 B.n894 585
R581 B.n896 B.n11 585
R582 B.n898 B.n897 585
R583 B.n899 B.n10 585
R584 B.n901 B.n900 585
R585 B.n902 B.n9 585
R586 B.n904 B.n903 585
R587 B.n905 B.n8 585
R588 B.n907 B.n906 585
R589 B.n908 B.n7 585
R590 B.n910 B.n909 585
R591 B.n911 B.n6 585
R592 B.n913 B.n912 585
R593 B.n914 B.n5 585
R594 B.n916 B.n915 585
R595 B.n917 B.n4 585
R596 B.n919 B.n918 585
R597 B.n920 B.n3 585
R598 B.n922 B.n921 585
R599 B.n923 B.n0 585
R600 B.n2 B.n1 585
R601 B.n239 B.n238 585
R602 B.n241 B.n240 585
R603 B.n242 B.n237 585
R604 B.n244 B.n243 585
R605 B.n245 B.n236 585
R606 B.n247 B.n246 585
R607 B.n248 B.n235 585
R608 B.n250 B.n249 585
R609 B.n251 B.n234 585
R610 B.n253 B.n252 585
R611 B.n254 B.n233 585
R612 B.n256 B.n255 585
R613 B.n257 B.n232 585
R614 B.n259 B.n258 585
R615 B.n260 B.n231 585
R616 B.n262 B.n261 585
R617 B.n263 B.n230 585
R618 B.n265 B.n264 585
R619 B.n266 B.n229 585
R620 B.n268 B.n267 585
R621 B.n269 B.n228 585
R622 B.n271 B.n270 585
R623 B.n272 B.n227 585
R624 B.n274 B.n273 585
R625 B.n275 B.n226 585
R626 B.n277 B.n276 585
R627 B.n278 B.n225 585
R628 B.n280 B.n279 585
R629 B.n281 B.n224 585
R630 B.n283 B.n282 585
R631 B.n284 B.n223 585
R632 B.n286 B.n285 585
R633 B.n287 B.n222 585
R634 B.n289 B.n288 585
R635 B.n290 B.n221 585
R636 B.n292 B.n291 585
R637 B.n293 B.n220 585
R638 B.n295 B.n294 585
R639 B.n296 B.n219 585
R640 B.n298 B.n297 585
R641 B.n299 B.n218 585
R642 B.n301 B.n300 585
R643 B.n302 B.n217 585
R644 B.n304 B.n303 585
R645 B.n305 B.n216 585
R646 B.n307 B.n306 585
R647 B.n308 B.n215 585
R648 B.n310 B.n309 585
R649 B.n311 B.n214 585
R650 B.n313 B.n312 585
R651 B.n314 B.n213 585
R652 B.n316 B.n315 585
R653 B.n317 B.n212 585
R654 B.n319 B.n318 585
R655 B.n320 B.n211 585
R656 B.n322 B.n321 585
R657 B.n323 B.n210 585
R658 B.n325 B.n210 487.695
R659 B.n491 B.n150 487.695
R660 B.n670 B.n669 487.695
R661 B.n838 B.n31 487.695
R662 B.n183 B.t9 351.205
R663 B.n177 B.t3 351.205
R664 B.n65 B.t6 351.205
R665 B.n58 B.t0 351.205
R666 B.n925 B.n924 256.663
R667 B.n924 B.n923 235.042
R668 B.n924 B.n2 235.042
R669 B.n177 B.t4 163.573
R670 B.n65 B.t8 163.573
R671 B.n183 B.t10 163.554
R672 B.n58 B.t2 163.554
R673 B.n326 B.n325 163.367
R674 B.n327 B.n326 163.367
R675 B.n327 B.n208 163.367
R676 B.n331 B.n208 163.367
R677 B.n332 B.n331 163.367
R678 B.n333 B.n332 163.367
R679 B.n333 B.n206 163.367
R680 B.n337 B.n206 163.367
R681 B.n338 B.n337 163.367
R682 B.n339 B.n338 163.367
R683 B.n339 B.n204 163.367
R684 B.n343 B.n204 163.367
R685 B.n344 B.n343 163.367
R686 B.n345 B.n344 163.367
R687 B.n345 B.n202 163.367
R688 B.n349 B.n202 163.367
R689 B.n350 B.n349 163.367
R690 B.n351 B.n350 163.367
R691 B.n351 B.n200 163.367
R692 B.n355 B.n200 163.367
R693 B.n356 B.n355 163.367
R694 B.n357 B.n356 163.367
R695 B.n357 B.n198 163.367
R696 B.n361 B.n198 163.367
R697 B.n362 B.n361 163.367
R698 B.n363 B.n362 163.367
R699 B.n363 B.n196 163.367
R700 B.n367 B.n196 163.367
R701 B.n368 B.n367 163.367
R702 B.n369 B.n368 163.367
R703 B.n369 B.n194 163.367
R704 B.n373 B.n194 163.367
R705 B.n374 B.n373 163.367
R706 B.n375 B.n374 163.367
R707 B.n375 B.n192 163.367
R708 B.n379 B.n192 163.367
R709 B.n380 B.n379 163.367
R710 B.n381 B.n380 163.367
R711 B.n381 B.n190 163.367
R712 B.n385 B.n190 163.367
R713 B.n386 B.n385 163.367
R714 B.n387 B.n386 163.367
R715 B.n387 B.n188 163.367
R716 B.n391 B.n188 163.367
R717 B.n392 B.n391 163.367
R718 B.n393 B.n392 163.367
R719 B.n393 B.n186 163.367
R720 B.n397 B.n186 163.367
R721 B.n398 B.n397 163.367
R722 B.n399 B.n398 163.367
R723 B.n399 B.n182 163.367
R724 B.n404 B.n182 163.367
R725 B.n405 B.n404 163.367
R726 B.n406 B.n405 163.367
R727 B.n406 B.n180 163.367
R728 B.n410 B.n180 163.367
R729 B.n411 B.n410 163.367
R730 B.n412 B.n411 163.367
R731 B.n412 B.n176 163.367
R732 B.n417 B.n176 163.367
R733 B.n418 B.n417 163.367
R734 B.n419 B.n418 163.367
R735 B.n419 B.n174 163.367
R736 B.n423 B.n174 163.367
R737 B.n424 B.n423 163.367
R738 B.n425 B.n424 163.367
R739 B.n425 B.n172 163.367
R740 B.n429 B.n172 163.367
R741 B.n430 B.n429 163.367
R742 B.n431 B.n430 163.367
R743 B.n431 B.n170 163.367
R744 B.n435 B.n170 163.367
R745 B.n436 B.n435 163.367
R746 B.n437 B.n436 163.367
R747 B.n437 B.n168 163.367
R748 B.n441 B.n168 163.367
R749 B.n442 B.n441 163.367
R750 B.n443 B.n442 163.367
R751 B.n443 B.n166 163.367
R752 B.n447 B.n166 163.367
R753 B.n448 B.n447 163.367
R754 B.n449 B.n448 163.367
R755 B.n449 B.n164 163.367
R756 B.n453 B.n164 163.367
R757 B.n454 B.n453 163.367
R758 B.n455 B.n454 163.367
R759 B.n455 B.n162 163.367
R760 B.n459 B.n162 163.367
R761 B.n460 B.n459 163.367
R762 B.n461 B.n460 163.367
R763 B.n461 B.n160 163.367
R764 B.n465 B.n160 163.367
R765 B.n466 B.n465 163.367
R766 B.n467 B.n466 163.367
R767 B.n467 B.n158 163.367
R768 B.n471 B.n158 163.367
R769 B.n472 B.n471 163.367
R770 B.n473 B.n472 163.367
R771 B.n473 B.n156 163.367
R772 B.n477 B.n156 163.367
R773 B.n478 B.n477 163.367
R774 B.n479 B.n478 163.367
R775 B.n479 B.n154 163.367
R776 B.n483 B.n154 163.367
R777 B.n484 B.n483 163.367
R778 B.n485 B.n484 163.367
R779 B.n485 B.n152 163.367
R780 B.n489 B.n152 163.367
R781 B.n490 B.n489 163.367
R782 B.n491 B.n490 163.367
R783 B.n669 B.n92 163.367
R784 B.n665 B.n92 163.367
R785 B.n665 B.n664 163.367
R786 B.n664 B.n663 163.367
R787 B.n663 B.n94 163.367
R788 B.n659 B.n94 163.367
R789 B.n659 B.n658 163.367
R790 B.n658 B.n657 163.367
R791 B.n657 B.n96 163.367
R792 B.n653 B.n96 163.367
R793 B.n653 B.n652 163.367
R794 B.n652 B.n651 163.367
R795 B.n651 B.n98 163.367
R796 B.n647 B.n98 163.367
R797 B.n647 B.n646 163.367
R798 B.n646 B.n645 163.367
R799 B.n645 B.n100 163.367
R800 B.n641 B.n100 163.367
R801 B.n641 B.n640 163.367
R802 B.n640 B.n639 163.367
R803 B.n639 B.n102 163.367
R804 B.n635 B.n102 163.367
R805 B.n635 B.n634 163.367
R806 B.n634 B.n633 163.367
R807 B.n633 B.n104 163.367
R808 B.n629 B.n104 163.367
R809 B.n629 B.n628 163.367
R810 B.n628 B.n627 163.367
R811 B.n627 B.n106 163.367
R812 B.n623 B.n106 163.367
R813 B.n623 B.n622 163.367
R814 B.n622 B.n621 163.367
R815 B.n621 B.n108 163.367
R816 B.n617 B.n108 163.367
R817 B.n617 B.n616 163.367
R818 B.n616 B.n615 163.367
R819 B.n615 B.n110 163.367
R820 B.n611 B.n110 163.367
R821 B.n611 B.n610 163.367
R822 B.n610 B.n609 163.367
R823 B.n609 B.n112 163.367
R824 B.n605 B.n112 163.367
R825 B.n605 B.n604 163.367
R826 B.n604 B.n603 163.367
R827 B.n603 B.n114 163.367
R828 B.n599 B.n114 163.367
R829 B.n599 B.n598 163.367
R830 B.n598 B.n597 163.367
R831 B.n597 B.n116 163.367
R832 B.n593 B.n116 163.367
R833 B.n593 B.n592 163.367
R834 B.n592 B.n591 163.367
R835 B.n591 B.n118 163.367
R836 B.n587 B.n118 163.367
R837 B.n587 B.n586 163.367
R838 B.n586 B.n585 163.367
R839 B.n585 B.n120 163.367
R840 B.n581 B.n120 163.367
R841 B.n581 B.n580 163.367
R842 B.n580 B.n579 163.367
R843 B.n579 B.n122 163.367
R844 B.n575 B.n122 163.367
R845 B.n575 B.n574 163.367
R846 B.n574 B.n573 163.367
R847 B.n573 B.n124 163.367
R848 B.n569 B.n124 163.367
R849 B.n569 B.n568 163.367
R850 B.n568 B.n567 163.367
R851 B.n567 B.n126 163.367
R852 B.n563 B.n126 163.367
R853 B.n563 B.n562 163.367
R854 B.n562 B.n561 163.367
R855 B.n561 B.n128 163.367
R856 B.n557 B.n128 163.367
R857 B.n557 B.n556 163.367
R858 B.n556 B.n555 163.367
R859 B.n555 B.n130 163.367
R860 B.n551 B.n130 163.367
R861 B.n551 B.n550 163.367
R862 B.n550 B.n549 163.367
R863 B.n549 B.n132 163.367
R864 B.n545 B.n132 163.367
R865 B.n545 B.n544 163.367
R866 B.n544 B.n543 163.367
R867 B.n543 B.n134 163.367
R868 B.n539 B.n134 163.367
R869 B.n539 B.n538 163.367
R870 B.n538 B.n537 163.367
R871 B.n537 B.n136 163.367
R872 B.n533 B.n136 163.367
R873 B.n533 B.n532 163.367
R874 B.n532 B.n531 163.367
R875 B.n531 B.n138 163.367
R876 B.n527 B.n138 163.367
R877 B.n527 B.n526 163.367
R878 B.n526 B.n525 163.367
R879 B.n525 B.n140 163.367
R880 B.n521 B.n140 163.367
R881 B.n521 B.n520 163.367
R882 B.n520 B.n519 163.367
R883 B.n519 B.n142 163.367
R884 B.n515 B.n142 163.367
R885 B.n515 B.n514 163.367
R886 B.n514 B.n513 163.367
R887 B.n513 B.n144 163.367
R888 B.n509 B.n144 163.367
R889 B.n509 B.n508 163.367
R890 B.n508 B.n507 163.367
R891 B.n507 B.n146 163.367
R892 B.n503 B.n146 163.367
R893 B.n503 B.n502 163.367
R894 B.n502 B.n501 163.367
R895 B.n501 B.n148 163.367
R896 B.n497 B.n148 163.367
R897 B.n497 B.n496 163.367
R898 B.n496 B.n495 163.367
R899 B.n495 B.n150 163.367
R900 B.n834 B.n31 163.367
R901 B.n834 B.n833 163.367
R902 B.n833 B.n832 163.367
R903 B.n832 B.n33 163.367
R904 B.n828 B.n33 163.367
R905 B.n828 B.n827 163.367
R906 B.n827 B.n826 163.367
R907 B.n826 B.n35 163.367
R908 B.n822 B.n35 163.367
R909 B.n822 B.n821 163.367
R910 B.n821 B.n820 163.367
R911 B.n820 B.n37 163.367
R912 B.n816 B.n37 163.367
R913 B.n816 B.n815 163.367
R914 B.n815 B.n814 163.367
R915 B.n814 B.n39 163.367
R916 B.n810 B.n39 163.367
R917 B.n810 B.n809 163.367
R918 B.n809 B.n808 163.367
R919 B.n808 B.n41 163.367
R920 B.n804 B.n41 163.367
R921 B.n804 B.n803 163.367
R922 B.n803 B.n802 163.367
R923 B.n802 B.n43 163.367
R924 B.n798 B.n43 163.367
R925 B.n798 B.n797 163.367
R926 B.n797 B.n796 163.367
R927 B.n796 B.n45 163.367
R928 B.n792 B.n45 163.367
R929 B.n792 B.n791 163.367
R930 B.n791 B.n790 163.367
R931 B.n790 B.n47 163.367
R932 B.n786 B.n47 163.367
R933 B.n786 B.n785 163.367
R934 B.n785 B.n784 163.367
R935 B.n784 B.n49 163.367
R936 B.n780 B.n49 163.367
R937 B.n780 B.n779 163.367
R938 B.n779 B.n778 163.367
R939 B.n778 B.n51 163.367
R940 B.n774 B.n51 163.367
R941 B.n774 B.n773 163.367
R942 B.n773 B.n772 163.367
R943 B.n772 B.n53 163.367
R944 B.n768 B.n53 163.367
R945 B.n768 B.n767 163.367
R946 B.n767 B.n766 163.367
R947 B.n766 B.n55 163.367
R948 B.n762 B.n55 163.367
R949 B.n762 B.n761 163.367
R950 B.n761 B.n760 163.367
R951 B.n760 B.n57 163.367
R952 B.n756 B.n57 163.367
R953 B.n756 B.n755 163.367
R954 B.n755 B.n754 163.367
R955 B.n754 B.n62 163.367
R956 B.n750 B.n62 163.367
R957 B.n750 B.n749 163.367
R958 B.n749 B.n748 163.367
R959 B.n748 B.n64 163.367
R960 B.n743 B.n64 163.367
R961 B.n743 B.n742 163.367
R962 B.n742 B.n741 163.367
R963 B.n741 B.n68 163.367
R964 B.n737 B.n68 163.367
R965 B.n737 B.n736 163.367
R966 B.n736 B.n735 163.367
R967 B.n735 B.n70 163.367
R968 B.n731 B.n70 163.367
R969 B.n731 B.n730 163.367
R970 B.n730 B.n729 163.367
R971 B.n729 B.n72 163.367
R972 B.n725 B.n72 163.367
R973 B.n725 B.n724 163.367
R974 B.n724 B.n723 163.367
R975 B.n723 B.n74 163.367
R976 B.n719 B.n74 163.367
R977 B.n719 B.n718 163.367
R978 B.n718 B.n717 163.367
R979 B.n717 B.n76 163.367
R980 B.n713 B.n76 163.367
R981 B.n713 B.n712 163.367
R982 B.n712 B.n711 163.367
R983 B.n711 B.n78 163.367
R984 B.n707 B.n78 163.367
R985 B.n707 B.n706 163.367
R986 B.n706 B.n705 163.367
R987 B.n705 B.n80 163.367
R988 B.n701 B.n80 163.367
R989 B.n701 B.n700 163.367
R990 B.n700 B.n699 163.367
R991 B.n699 B.n82 163.367
R992 B.n695 B.n82 163.367
R993 B.n695 B.n694 163.367
R994 B.n694 B.n693 163.367
R995 B.n693 B.n84 163.367
R996 B.n689 B.n84 163.367
R997 B.n689 B.n688 163.367
R998 B.n688 B.n687 163.367
R999 B.n687 B.n86 163.367
R1000 B.n683 B.n86 163.367
R1001 B.n683 B.n682 163.367
R1002 B.n682 B.n681 163.367
R1003 B.n681 B.n88 163.367
R1004 B.n677 B.n88 163.367
R1005 B.n677 B.n676 163.367
R1006 B.n676 B.n675 163.367
R1007 B.n675 B.n90 163.367
R1008 B.n671 B.n90 163.367
R1009 B.n671 B.n670 163.367
R1010 B.n839 B.n838 163.367
R1011 B.n840 B.n839 163.367
R1012 B.n840 B.n29 163.367
R1013 B.n844 B.n29 163.367
R1014 B.n845 B.n844 163.367
R1015 B.n846 B.n845 163.367
R1016 B.n846 B.n27 163.367
R1017 B.n850 B.n27 163.367
R1018 B.n851 B.n850 163.367
R1019 B.n852 B.n851 163.367
R1020 B.n852 B.n25 163.367
R1021 B.n856 B.n25 163.367
R1022 B.n857 B.n856 163.367
R1023 B.n858 B.n857 163.367
R1024 B.n858 B.n23 163.367
R1025 B.n862 B.n23 163.367
R1026 B.n863 B.n862 163.367
R1027 B.n864 B.n863 163.367
R1028 B.n864 B.n21 163.367
R1029 B.n868 B.n21 163.367
R1030 B.n869 B.n868 163.367
R1031 B.n870 B.n869 163.367
R1032 B.n870 B.n19 163.367
R1033 B.n874 B.n19 163.367
R1034 B.n875 B.n874 163.367
R1035 B.n876 B.n875 163.367
R1036 B.n876 B.n17 163.367
R1037 B.n880 B.n17 163.367
R1038 B.n881 B.n880 163.367
R1039 B.n882 B.n881 163.367
R1040 B.n882 B.n15 163.367
R1041 B.n886 B.n15 163.367
R1042 B.n887 B.n886 163.367
R1043 B.n888 B.n887 163.367
R1044 B.n888 B.n13 163.367
R1045 B.n892 B.n13 163.367
R1046 B.n893 B.n892 163.367
R1047 B.n894 B.n893 163.367
R1048 B.n894 B.n11 163.367
R1049 B.n898 B.n11 163.367
R1050 B.n899 B.n898 163.367
R1051 B.n900 B.n899 163.367
R1052 B.n900 B.n9 163.367
R1053 B.n904 B.n9 163.367
R1054 B.n905 B.n904 163.367
R1055 B.n906 B.n905 163.367
R1056 B.n906 B.n7 163.367
R1057 B.n910 B.n7 163.367
R1058 B.n911 B.n910 163.367
R1059 B.n912 B.n911 163.367
R1060 B.n912 B.n5 163.367
R1061 B.n916 B.n5 163.367
R1062 B.n917 B.n916 163.367
R1063 B.n918 B.n917 163.367
R1064 B.n918 B.n3 163.367
R1065 B.n922 B.n3 163.367
R1066 B.n923 B.n922 163.367
R1067 B.n238 B.n2 163.367
R1068 B.n241 B.n238 163.367
R1069 B.n242 B.n241 163.367
R1070 B.n243 B.n242 163.367
R1071 B.n243 B.n236 163.367
R1072 B.n247 B.n236 163.367
R1073 B.n248 B.n247 163.367
R1074 B.n249 B.n248 163.367
R1075 B.n249 B.n234 163.367
R1076 B.n253 B.n234 163.367
R1077 B.n254 B.n253 163.367
R1078 B.n255 B.n254 163.367
R1079 B.n255 B.n232 163.367
R1080 B.n259 B.n232 163.367
R1081 B.n260 B.n259 163.367
R1082 B.n261 B.n260 163.367
R1083 B.n261 B.n230 163.367
R1084 B.n265 B.n230 163.367
R1085 B.n266 B.n265 163.367
R1086 B.n267 B.n266 163.367
R1087 B.n267 B.n228 163.367
R1088 B.n271 B.n228 163.367
R1089 B.n272 B.n271 163.367
R1090 B.n273 B.n272 163.367
R1091 B.n273 B.n226 163.367
R1092 B.n277 B.n226 163.367
R1093 B.n278 B.n277 163.367
R1094 B.n279 B.n278 163.367
R1095 B.n279 B.n224 163.367
R1096 B.n283 B.n224 163.367
R1097 B.n284 B.n283 163.367
R1098 B.n285 B.n284 163.367
R1099 B.n285 B.n222 163.367
R1100 B.n289 B.n222 163.367
R1101 B.n290 B.n289 163.367
R1102 B.n291 B.n290 163.367
R1103 B.n291 B.n220 163.367
R1104 B.n295 B.n220 163.367
R1105 B.n296 B.n295 163.367
R1106 B.n297 B.n296 163.367
R1107 B.n297 B.n218 163.367
R1108 B.n301 B.n218 163.367
R1109 B.n302 B.n301 163.367
R1110 B.n303 B.n302 163.367
R1111 B.n303 B.n216 163.367
R1112 B.n307 B.n216 163.367
R1113 B.n308 B.n307 163.367
R1114 B.n309 B.n308 163.367
R1115 B.n309 B.n214 163.367
R1116 B.n313 B.n214 163.367
R1117 B.n314 B.n313 163.367
R1118 B.n315 B.n314 163.367
R1119 B.n315 B.n212 163.367
R1120 B.n319 B.n212 163.367
R1121 B.n320 B.n319 163.367
R1122 B.n321 B.n320 163.367
R1123 B.n321 B.n210 163.367
R1124 B.n178 B.t5 108.108
R1125 B.n66 B.t7 108.108
R1126 B.n184 B.t11 108.088
R1127 B.n59 B.t1 108.088
R1128 B.n401 B.n184 59.5399
R1129 B.n415 B.n178 59.5399
R1130 B.n746 B.n66 59.5399
R1131 B.n60 B.n59 59.5399
R1132 B.n184 B.n183 55.4672
R1133 B.n178 B.n177 55.4672
R1134 B.n66 B.n65 55.4672
R1135 B.n59 B.n58 55.4672
R1136 B.n837 B.n836 31.6883
R1137 B.n668 B.n91 31.6883
R1138 B.n493 B.n492 31.6883
R1139 B.n324 B.n323 31.6883
R1140 B B.n925 18.0485
R1141 B.n837 B.n30 10.6151
R1142 B.n841 B.n30 10.6151
R1143 B.n842 B.n841 10.6151
R1144 B.n843 B.n842 10.6151
R1145 B.n843 B.n28 10.6151
R1146 B.n847 B.n28 10.6151
R1147 B.n848 B.n847 10.6151
R1148 B.n849 B.n848 10.6151
R1149 B.n849 B.n26 10.6151
R1150 B.n853 B.n26 10.6151
R1151 B.n854 B.n853 10.6151
R1152 B.n855 B.n854 10.6151
R1153 B.n855 B.n24 10.6151
R1154 B.n859 B.n24 10.6151
R1155 B.n860 B.n859 10.6151
R1156 B.n861 B.n860 10.6151
R1157 B.n861 B.n22 10.6151
R1158 B.n865 B.n22 10.6151
R1159 B.n866 B.n865 10.6151
R1160 B.n867 B.n866 10.6151
R1161 B.n867 B.n20 10.6151
R1162 B.n871 B.n20 10.6151
R1163 B.n872 B.n871 10.6151
R1164 B.n873 B.n872 10.6151
R1165 B.n873 B.n18 10.6151
R1166 B.n877 B.n18 10.6151
R1167 B.n878 B.n877 10.6151
R1168 B.n879 B.n878 10.6151
R1169 B.n879 B.n16 10.6151
R1170 B.n883 B.n16 10.6151
R1171 B.n884 B.n883 10.6151
R1172 B.n885 B.n884 10.6151
R1173 B.n885 B.n14 10.6151
R1174 B.n889 B.n14 10.6151
R1175 B.n890 B.n889 10.6151
R1176 B.n891 B.n890 10.6151
R1177 B.n891 B.n12 10.6151
R1178 B.n895 B.n12 10.6151
R1179 B.n896 B.n895 10.6151
R1180 B.n897 B.n896 10.6151
R1181 B.n897 B.n10 10.6151
R1182 B.n901 B.n10 10.6151
R1183 B.n902 B.n901 10.6151
R1184 B.n903 B.n902 10.6151
R1185 B.n903 B.n8 10.6151
R1186 B.n907 B.n8 10.6151
R1187 B.n908 B.n907 10.6151
R1188 B.n909 B.n908 10.6151
R1189 B.n909 B.n6 10.6151
R1190 B.n913 B.n6 10.6151
R1191 B.n914 B.n913 10.6151
R1192 B.n915 B.n914 10.6151
R1193 B.n915 B.n4 10.6151
R1194 B.n919 B.n4 10.6151
R1195 B.n920 B.n919 10.6151
R1196 B.n921 B.n920 10.6151
R1197 B.n921 B.n0 10.6151
R1198 B.n836 B.n835 10.6151
R1199 B.n835 B.n32 10.6151
R1200 B.n831 B.n32 10.6151
R1201 B.n831 B.n830 10.6151
R1202 B.n830 B.n829 10.6151
R1203 B.n829 B.n34 10.6151
R1204 B.n825 B.n34 10.6151
R1205 B.n825 B.n824 10.6151
R1206 B.n824 B.n823 10.6151
R1207 B.n823 B.n36 10.6151
R1208 B.n819 B.n36 10.6151
R1209 B.n819 B.n818 10.6151
R1210 B.n818 B.n817 10.6151
R1211 B.n817 B.n38 10.6151
R1212 B.n813 B.n38 10.6151
R1213 B.n813 B.n812 10.6151
R1214 B.n812 B.n811 10.6151
R1215 B.n811 B.n40 10.6151
R1216 B.n807 B.n40 10.6151
R1217 B.n807 B.n806 10.6151
R1218 B.n806 B.n805 10.6151
R1219 B.n805 B.n42 10.6151
R1220 B.n801 B.n42 10.6151
R1221 B.n801 B.n800 10.6151
R1222 B.n800 B.n799 10.6151
R1223 B.n799 B.n44 10.6151
R1224 B.n795 B.n44 10.6151
R1225 B.n795 B.n794 10.6151
R1226 B.n794 B.n793 10.6151
R1227 B.n793 B.n46 10.6151
R1228 B.n789 B.n46 10.6151
R1229 B.n789 B.n788 10.6151
R1230 B.n788 B.n787 10.6151
R1231 B.n787 B.n48 10.6151
R1232 B.n783 B.n48 10.6151
R1233 B.n783 B.n782 10.6151
R1234 B.n782 B.n781 10.6151
R1235 B.n781 B.n50 10.6151
R1236 B.n777 B.n50 10.6151
R1237 B.n777 B.n776 10.6151
R1238 B.n776 B.n775 10.6151
R1239 B.n775 B.n52 10.6151
R1240 B.n771 B.n52 10.6151
R1241 B.n771 B.n770 10.6151
R1242 B.n770 B.n769 10.6151
R1243 B.n769 B.n54 10.6151
R1244 B.n765 B.n54 10.6151
R1245 B.n765 B.n764 10.6151
R1246 B.n764 B.n763 10.6151
R1247 B.n763 B.n56 10.6151
R1248 B.n759 B.n758 10.6151
R1249 B.n758 B.n757 10.6151
R1250 B.n757 B.n61 10.6151
R1251 B.n753 B.n61 10.6151
R1252 B.n753 B.n752 10.6151
R1253 B.n752 B.n751 10.6151
R1254 B.n751 B.n63 10.6151
R1255 B.n747 B.n63 10.6151
R1256 B.n745 B.n744 10.6151
R1257 B.n744 B.n67 10.6151
R1258 B.n740 B.n67 10.6151
R1259 B.n740 B.n739 10.6151
R1260 B.n739 B.n738 10.6151
R1261 B.n738 B.n69 10.6151
R1262 B.n734 B.n69 10.6151
R1263 B.n734 B.n733 10.6151
R1264 B.n733 B.n732 10.6151
R1265 B.n732 B.n71 10.6151
R1266 B.n728 B.n71 10.6151
R1267 B.n728 B.n727 10.6151
R1268 B.n727 B.n726 10.6151
R1269 B.n726 B.n73 10.6151
R1270 B.n722 B.n73 10.6151
R1271 B.n722 B.n721 10.6151
R1272 B.n721 B.n720 10.6151
R1273 B.n720 B.n75 10.6151
R1274 B.n716 B.n75 10.6151
R1275 B.n716 B.n715 10.6151
R1276 B.n715 B.n714 10.6151
R1277 B.n714 B.n77 10.6151
R1278 B.n710 B.n77 10.6151
R1279 B.n710 B.n709 10.6151
R1280 B.n709 B.n708 10.6151
R1281 B.n708 B.n79 10.6151
R1282 B.n704 B.n79 10.6151
R1283 B.n704 B.n703 10.6151
R1284 B.n703 B.n702 10.6151
R1285 B.n702 B.n81 10.6151
R1286 B.n698 B.n81 10.6151
R1287 B.n698 B.n697 10.6151
R1288 B.n697 B.n696 10.6151
R1289 B.n696 B.n83 10.6151
R1290 B.n692 B.n83 10.6151
R1291 B.n692 B.n691 10.6151
R1292 B.n691 B.n690 10.6151
R1293 B.n690 B.n85 10.6151
R1294 B.n686 B.n85 10.6151
R1295 B.n686 B.n685 10.6151
R1296 B.n685 B.n684 10.6151
R1297 B.n684 B.n87 10.6151
R1298 B.n680 B.n87 10.6151
R1299 B.n680 B.n679 10.6151
R1300 B.n679 B.n678 10.6151
R1301 B.n678 B.n89 10.6151
R1302 B.n674 B.n89 10.6151
R1303 B.n674 B.n673 10.6151
R1304 B.n673 B.n672 10.6151
R1305 B.n672 B.n91 10.6151
R1306 B.n668 B.n667 10.6151
R1307 B.n667 B.n666 10.6151
R1308 B.n666 B.n93 10.6151
R1309 B.n662 B.n93 10.6151
R1310 B.n662 B.n661 10.6151
R1311 B.n661 B.n660 10.6151
R1312 B.n660 B.n95 10.6151
R1313 B.n656 B.n95 10.6151
R1314 B.n656 B.n655 10.6151
R1315 B.n655 B.n654 10.6151
R1316 B.n654 B.n97 10.6151
R1317 B.n650 B.n97 10.6151
R1318 B.n650 B.n649 10.6151
R1319 B.n649 B.n648 10.6151
R1320 B.n648 B.n99 10.6151
R1321 B.n644 B.n99 10.6151
R1322 B.n644 B.n643 10.6151
R1323 B.n643 B.n642 10.6151
R1324 B.n642 B.n101 10.6151
R1325 B.n638 B.n101 10.6151
R1326 B.n638 B.n637 10.6151
R1327 B.n637 B.n636 10.6151
R1328 B.n636 B.n103 10.6151
R1329 B.n632 B.n103 10.6151
R1330 B.n632 B.n631 10.6151
R1331 B.n631 B.n630 10.6151
R1332 B.n630 B.n105 10.6151
R1333 B.n626 B.n105 10.6151
R1334 B.n626 B.n625 10.6151
R1335 B.n625 B.n624 10.6151
R1336 B.n624 B.n107 10.6151
R1337 B.n620 B.n107 10.6151
R1338 B.n620 B.n619 10.6151
R1339 B.n619 B.n618 10.6151
R1340 B.n618 B.n109 10.6151
R1341 B.n614 B.n109 10.6151
R1342 B.n614 B.n613 10.6151
R1343 B.n613 B.n612 10.6151
R1344 B.n612 B.n111 10.6151
R1345 B.n608 B.n111 10.6151
R1346 B.n608 B.n607 10.6151
R1347 B.n607 B.n606 10.6151
R1348 B.n606 B.n113 10.6151
R1349 B.n602 B.n113 10.6151
R1350 B.n602 B.n601 10.6151
R1351 B.n601 B.n600 10.6151
R1352 B.n600 B.n115 10.6151
R1353 B.n596 B.n115 10.6151
R1354 B.n596 B.n595 10.6151
R1355 B.n595 B.n594 10.6151
R1356 B.n594 B.n117 10.6151
R1357 B.n590 B.n117 10.6151
R1358 B.n590 B.n589 10.6151
R1359 B.n589 B.n588 10.6151
R1360 B.n588 B.n119 10.6151
R1361 B.n584 B.n119 10.6151
R1362 B.n584 B.n583 10.6151
R1363 B.n583 B.n582 10.6151
R1364 B.n582 B.n121 10.6151
R1365 B.n578 B.n121 10.6151
R1366 B.n578 B.n577 10.6151
R1367 B.n577 B.n576 10.6151
R1368 B.n576 B.n123 10.6151
R1369 B.n572 B.n123 10.6151
R1370 B.n572 B.n571 10.6151
R1371 B.n571 B.n570 10.6151
R1372 B.n570 B.n125 10.6151
R1373 B.n566 B.n125 10.6151
R1374 B.n566 B.n565 10.6151
R1375 B.n565 B.n564 10.6151
R1376 B.n564 B.n127 10.6151
R1377 B.n560 B.n127 10.6151
R1378 B.n560 B.n559 10.6151
R1379 B.n559 B.n558 10.6151
R1380 B.n558 B.n129 10.6151
R1381 B.n554 B.n129 10.6151
R1382 B.n554 B.n553 10.6151
R1383 B.n553 B.n552 10.6151
R1384 B.n552 B.n131 10.6151
R1385 B.n548 B.n131 10.6151
R1386 B.n548 B.n547 10.6151
R1387 B.n547 B.n546 10.6151
R1388 B.n546 B.n133 10.6151
R1389 B.n542 B.n133 10.6151
R1390 B.n542 B.n541 10.6151
R1391 B.n541 B.n540 10.6151
R1392 B.n540 B.n135 10.6151
R1393 B.n536 B.n135 10.6151
R1394 B.n536 B.n535 10.6151
R1395 B.n535 B.n534 10.6151
R1396 B.n534 B.n137 10.6151
R1397 B.n530 B.n137 10.6151
R1398 B.n530 B.n529 10.6151
R1399 B.n529 B.n528 10.6151
R1400 B.n528 B.n139 10.6151
R1401 B.n524 B.n139 10.6151
R1402 B.n524 B.n523 10.6151
R1403 B.n523 B.n522 10.6151
R1404 B.n522 B.n141 10.6151
R1405 B.n518 B.n141 10.6151
R1406 B.n518 B.n517 10.6151
R1407 B.n517 B.n516 10.6151
R1408 B.n516 B.n143 10.6151
R1409 B.n512 B.n143 10.6151
R1410 B.n512 B.n511 10.6151
R1411 B.n511 B.n510 10.6151
R1412 B.n510 B.n145 10.6151
R1413 B.n506 B.n145 10.6151
R1414 B.n506 B.n505 10.6151
R1415 B.n505 B.n504 10.6151
R1416 B.n504 B.n147 10.6151
R1417 B.n500 B.n147 10.6151
R1418 B.n500 B.n499 10.6151
R1419 B.n499 B.n498 10.6151
R1420 B.n498 B.n149 10.6151
R1421 B.n494 B.n149 10.6151
R1422 B.n494 B.n493 10.6151
R1423 B.n239 B.n1 10.6151
R1424 B.n240 B.n239 10.6151
R1425 B.n240 B.n237 10.6151
R1426 B.n244 B.n237 10.6151
R1427 B.n245 B.n244 10.6151
R1428 B.n246 B.n245 10.6151
R1429 B.n246 B.n235 10.6151
R1430 B.n250 B.n235 10.6151
R1431 B.n251 B.n250 10.6151
R1432 B.n252 B.n251 10.6151
R1433 B.n252 B.n233 10.6151
R1434 B.n256 B.n233 10.6151
R1435 B.n257 B.n256 10.6151
R1436 B.n258 B.n257 10.6151
R1437 B.n258 B.n231 10.6151
R1438 B.n262 B.n231 10.6151
R1439 B.n263 B.n262 10.6151
R1440 B.n264 B.n263 10.6151
R1441 B.n264 B.n229 10.6151
R1442 B.n268 B.n229 10.6151
R1443 B.n269 B.n268 10.6151
R1444 B.n270 B.n269 10.6151
R1445 B.n270 B.n227 10.6151
R1446 B.n274 B.n227 10.6151
R1447 B.n275 B.n274 10.6151
R1448 B.n276 B.n275 10.6151
R1449 B.n276 B.n225 10.6151
R1450 B.n280 B.n225 10.6151
R1451 B.n281 B.n280 10.6151
R1452 B.n282 B.n281 10.6151
R1453 B.n282 B.n223 10.6151
R1454 B.n286 B.n223 10.6151
R1455 B.n287 B.n286 10.6151
R1456 B.n288 B.n287 10.6151
R1457 B.n288 B.n221 10.6151
R1458 B.n292 B.n221 10.6151
R1459 B.n293 B.n292 10.6151
R1460 B.n294 B.n293 10.6151
R1461 B.n294 B.n219 10.6151
R1462 B.n298 B.n219 10.6151
R1463 B.n299 B.n298 10.6151
R1464 B.n300 B.n299 10.6151
R1465 B.n300 B.n217 10.6151
R1466 B.n304 B.n217 10.6151
R1467 B.n305 B.n304 10.6151
R1468 B.n306 B.n305 10.6151
R1469 B.n306 B.n215 10.6151
R1470 B.n310 B.n215 10.6151
R1471 B.n311 B.n310 10.6151
R1472 B.n312 B.n311 10.6151
R1473 B.n312 B.n213 10.6151
R1474 B.n316 B.n213 10.6151
R1475 B.n317 B.n316 10.6151
R1476 B.n318 B.n317 10.6151
R1477 B.n318 B.n211 10.6151
R1478 B.n322 B.n211 10.6151
R1479 B.n323 B.n322 10.6151
R1480 B.n324 B.n209 10.6151
R1481 B.n328 B.n209 10.6151
R1482 B.n329 B.n328 10.6151
R1483 B.n330 B.n329 10.6151
R1484 B.n330 B.n207 10.6151
R1485 B.n334 B.n207 10.6151
R1486 B.n335 B.n334 10.6151
R1487 B.n336 B.n335 10.6151
R1488 B.n336 B.n205 10.6151
R1489 B.n340 B.n205 10.6151
R1490 B.n341 B.n340 10.6151
R1491 B.n342 B.n341 10.6151
R1492 B.n342 B.n203 10.6151
R1493 B.n346 B.n203 10.6151
R1494 B.n347 B.n346 10.6151
R1495 B.n348 B.n347 10.6151
R1496 B.n348 B.n201 10.6151
R1497 B.n352 B.n201 10.6151
R1498 B.n353 B.n352 10.6151
R1499 B.n354 B.n353 10.6151
R1500 B.n354 B.n199 10.6151
R1501 B.n358 B.n199 10.6151
R1502 B.n359 B.n358 10.6151
R1503 B.n360 B.n359 10.6151
R1504 B.n360 B.n197 10.6151
R1505 B.n364 B.n197 10.6151
R1506 B.n365 B.n364 10.6151
R1507 B.n366 B.n365 10.6151
R1508 B.n366 B.n195 10.6151
R1509 B.n370 B.n195 10.6151
R1510 B.n371 B.n370 10.6151
R1511 B.n372 B.n371 10.6151
R1512 B.n372 B.n193 10.6151
R1513 B.n376 B.n193 10.6151
R1514 B.n377 B.n376 10.6151
R1515 B.n378 B.n377 10.6151
R1516 B.n378 B.n191 10.6151
R1517 B.n382 B.n191 10.6151
R1518 B.n383 B.n382 10.6151
R1519 B.n384 B.n383 10.6151
R1520 B.n384 B.n189 10.6151
R1521 B.n388 B.n189 10.6151
R1522 B.n389 B.n388 10.6151
R1523 B.n390 B.n389 10.6151
R1524 B.n390 B.n187 10.6151
R1525 B.n394 B.n187 10.6151
R1526 B.n395 B.n394 10.6151
R1527 B.n396 B.n395 10.6151
R1528 B.n396 B.n185 10.6151
R1529 B.n400 B.n185 10.6151
R1530 B.n403 B.n402 10.6151
R1531 B.n403 B.n181 10.6151
R1532 B.n407 B.n181 10.6151
R1533 B.n408 B.n407 10.6151
R1534 B.n409 B.n408 10.6151
R1535 B.n409 B.n179 10.6151
R1536 B.n413 B.n179 10.6151
R1537 B.n414 B.n413 10.6151
R1538 B.n416 B.n175 10.6151
R1539 B.n420 B.n175 10.6151
R1540 B.n421 B.n420 10.6151
R1541 B.n422 B.n421 10.6151
R1542 B.n422 B.n173 10.6151
R1543 B.n426 B.n173 10.6151
R1544 B.n427 B.n426 10.6151
R1545 B.n428 B.n427 10.6151
R1546 B.n428 B.n171 10.6151
R1547 B.n432 B.n171 10.6151
R1548 B.n433 B.n432 10.6151
R1549 B.n434 B.n433 10.6151
R1550 B.n434 B.n169 10.6151
R1551 B.n438 B.n169 10.6151
R1552 B.n439 B.n438 10.6151
R1553 B.n440 B.n439 10.6151
R1554 B.n440 B.n167 10.6151
R1555 B.n444 B.n167 10.6151
R1556 B.n445 B.n444 10.6151
R1557 B.n446 B.n445 10.6151
R1558 B.n446 B.n165 10.6151
R1559 B.n450 B.n165 10.6151
R1560 B.n451 B.n450 10.6151
R1561 B.n452 B.n451 10.6151
R1562 B.n452 B.n163 10.6151
R1563 B.n456 B.n163 10.6151
R1564 B.n457 B.n456 10.6151
R1565 B.n458 B.n457 10.6151
R1566 B.n458 B.n161 10.6151
R1567 B.n462 B.n161 10.6151
R1568 B.n463 B.n462 10.6151
R1569 B.n464 B.n463 10.6151
R1570 B.n464 B.n159 10.6151
R1571 B.n468 B.n159 10.6151
R1572 B.n469 B.n468 10.6151
R1573 B.n470 B.n469 10.6151
R1574 B.n470 B.n157 10.6151
R1575 B.n474 B.n157 10.6151
R1576 B.n475 B.n474 10.6151
R1577 B.n476 B.n475 10.6151
R1578 B.n476 B.n155 10.6151
R1579 B.n480 B.n155 10.6151
R1580 B.n481 B.n480 10.6151
R1581 B.n482 B.n481 10.6151
R1582 B.n482 B.n153 10.6151
R1583 B.n486 B.n153 10.6151
R1584 B.n487 B.n486 10.6151
R1585 B.n488 B.n487 10.6151
R1586 B.n488 B.n151 10.6151
R1587 B.n492 B.n151 10.6151
R1588 B.n925 B.n0 8.11757
R1589 B.n925 B.n1 8.11757
R1590 B.n759 B.n60 6.5566
R1591 B.n747 B.n746 6.5566
R1592 B.n402 B.n401 6.5566
R1593 B.n415 B.n414 6.5566
R1594 B.n60 B.n56 4.05904
R1595 B.n746 B.n745 4.05904
R1596 B.n401 B.n400 4.05904
R1597 B.n416 B.n415 4.05904
R1598 VN.n10 VN.t6 177.169
R1599 VN.n49 VN.t5 177.169
R1600 VN.n75 VN.n39 161.3
R1601 VN.n74 VN.n73 161.3
R1602 VN.n72 VN.n40 161.3
R1603 VN.n71 VN.n70 161.3
R1604 VN.n69 VN.n41 161.3
R1605 VN.n68 VN.n67 161.3
R1606 VN.n66 VN.n65 161.3
R1607 VN.n64 VN.n43 161.3
R1608 VN.n63 VN.n62 161.3
R1609 VN.n61 VN.n44 161.3
R1610 VN.n60 VN.n59 161.3
R1611 VN.n58 VN.n45 161.3
R1612 VN.n57 VN.n56 161.3
R1613 VN.n55 VN.n46 161.3
R1614 VN.n54 VN.n53 161.3
R1615 VN.n52 VN.n47 161.3
R1616 VN.n51 VN.n50 161.3
R1617 VN.n36 VN.n0 161.3
R1618 VN.n35 VN.n34 161.3
R1619 VN.n33 VN.n1 161.3
R1620 VN.n32 VN.n31 161.3
R1621 VN.n30 VN.n2 161.3
R1622 VN.n29 VN.n28 161.3
R1623 VN.n27 VN.n26 161.3
R1624 VN.n25 VN.n4 161.3
R1625 VN.n24 VN.n23 161.3
R1626 VN.n22 VN.n5 161.3
R1627 VN.n21 VN.n20 161.3
R1628 VN.n19 VN.n6 161.3
R1629 VN.n18 VN.n17 161.3
R1630 VN.n16 VN.n7 161.3
R1631 VN.n15 VN.n14 161.3
R1632 VN.n13 VN.n8 161.3
R1633 VN.n12 VN.n11 161.3
R1634 VN.n19 VN.t1 143.267
R1635 VN.n9 VN.t2 143.267
R1636 VN.n3 VN.t7 143.267
R1637 VN.n37 VN.t4 143.267
R1638 VN.n58 VN.t9 143.267
R1639 VN.n48 VN.t8 143.267
R1640 VN.n42 VN.t0 143.267
R1641 VN.n76 VN.t3 143.267
R1642 VN.n38 VN.n37 100.088
R1643 VN.n77 VN.n76 100.088
R1644 VN.n31 VN.n1 56.5617
R1645 VN.n70 VN.n40 56.5617
R1646 VN VN.n77 55.3315
R1647 VN.n10 VN.n9 55.0245
R1648 VN.n49 VN.n48 55.0245
R1649 VN.n14 VN.n7 47.3584
R1650 VN.n24 VN.n5 47.3584
R1651 VN.n53 VN.n46 47.3584
R1652 VN.n63 VN.n44 47.3584
R1653 VN.n14 VN.n13 33.7956
R1654 VN.n25 VN.n24 33.7956
R1655 VN.n53 VN.n52 33.7956
R1656 VN.n64 VN.n63 33.7956
R1657 VN.n13 VN.n12 24.5923
R1658 VN.n18 VN.n7 24.5923
R1659 VN.n19 VN.n18 24.5923
R1660 VN.n20 VN.n19 24.5923
R1661 VN.n20 VN.n5 24.5923
R1662 VN.n26 VN.n25 24.5923
R1663 VN.n30 VN.n29 24.5923
R1664 VN.n31 VN.n30 24.5923
R1665 VN.n35 VN.n1 24.5923
R1666 VN.n36 VN.n35 24.5923
R1667 VN.n52 VN.n51 24.5923
R1668 VN.n59 VN.n44 24.5923
R1669 VN.n59 VN.n58 24.5923
R1670 VN.n58 VN.n57 24.5923
R1671 VN.n57 VN.n46 24.5923
R1672 VN.n70 VN.n69 24.5923
R1673 VN.n69 VN.n68 24.5923
R1674 VN.n65 VN.n64 24.5923
R1675 VN.n75 VN.n74 24.5923
R1676 VN.n74 VN.n40 24.5923
R1677 VN.n12 VN.n9 17.7066
R1678 VN.n26 VN.n3 17.7066
R1679 VN.n51 VN.n48 17.7066
R1680 VN.n65 VN.n42 17.7066
R1681 VN.n37 VN.n36 10.8209
R1682 VN.n76 VN.n75 10.8209
R1683 VN.n29 VN.n3 6.88621
R1684 VN.n68 VN.n42 6.88621
R1685 VN.n50 VN.n49 6.78213
R1686 VN.n11 VN.n10 6.78213
R1687 VN.n77 VN.n39 0.278335
R1688 VN.n38 VN.n0 0.278335
R1689 VN.n73 VN.n39 0.189894
R1690 VN.n73 VN.n72 0.189894
R1691 VN.n72 VN.n71 0.189894
R1692 VN.n71 VN.n41 0.189894
R1693 VN.n67 VN.n41 0.189894
R1694 VN.n67 VN.n66 0.189894
R1695 VN.n66 VN.n43 0.189894
R1696 VN.n62 VN.n43 0.189894
R1697 VN.n62 VN.n61 0.189894
R1698 VN.n61 VN.n60 0.189894
R1699 VN.n60 VN.n45 0.189894
R1700 VN.n56 VN.n45 0.189894
R1701 VN.n56 VN.n55 0.189894
R1702 VN.n55 VN.n54 0.189894
R1703 VN.n54 VN.n47 0.189894
R1704 VN.n50 VN.n47 0.189894
R1705 VN.n11 VN.n8 0.189894
R1706 VN.n15 VN.n8 0.189894
R1707 VN.n16 VN.n15 0.189894
R1708 VN.n17 VN.n16 0.189894
R1709 VN.n17 VN.n6 0.189894
R1710 VN.n21 VN.n6 0.189894
R1711 VN.n22 VN.n21 0.189894
R1712 VN.n23 VN.n22 0.189894
R1713 VN.n23 VN.n4 0.189894
R1714 VN.n27 VN.n4 0.189894
R1715 VN.n28 VN.n27 0.189894
R1716 VN.n28 VN.n2 0.189894
R1717 VN.n32 VN.n2 0.189894
R1718 VN.n33 VN.n32 0.189894
R1719 VN.n34 VN.n33 0.189894
R1720 VN.n34 VN.n0 0.189894
R1721 VN VN.n38 0.153485
R1722 VDD2.n1 VDD2.t3 75.9074
R1723 VDD2.n4 VDD2.t6 73.4422
R1724 VDD2.n3 VDD2.n2 73.0745
R1725 VDD2 VDD2.n7 73.0717
R1726 VDD2.n6 VDD2.n5 71.2809
R1727 VDD2.n1 VDD2.n0 71.2807
R1728 VDD2.n4 VDD2.n3 48.392
R1729 VDD2.n6 VDD2.n4 2.46602
R1730 VDD2.n7 VDD2.t1 2.16174
R1731 VDD2.n7 VDD2.t4 2.16174
R1732 VDD2.n5 VDD2.t9 2.16174
R1733 VDD2.n5 VDD2.t0 2.16174
R1734 VDD2.n2 VDD2.t2 2.16174
R1735 VDD2.n2 VDD2.t5 2.16174
R1736 VDD2.n0 VDD2.t7 2.16174
R1737 VDD2.n0 VDD2.t8 2.16174
R1738 VDD2 VDD2.n6 0.675069
R1739 VDD2.n3 VDD2.n1 0.561533
C0 VDD2 VN 13.1673f
C1 VTAIL w_n4402_n3976# 3.62611f
C2 VDD1 w_n4402_n3976# 2.9736f
C3 VP VTAIL 13.658501f
C4 VP VDD1 13.584599f
C5 VP w_n4402_n3976# 10.008901f
C6 VTAIL B 4.3796f
C7 VTAIL VN 13.644199f
C8 VDD1 B 2.69251f
C9 VDD1 VN 0.153514f
C10 VDD2 VTAIL 11.8517f
C11 VDD2 VDD1 2.12906f
C12 B w_n4402_n3976# 11.2817f
C13 VN w_n4402_n3976# 9.43599f
C14 VDD2 w_n4402_n3976# 3.11352f
C15 VP B 2.26794f
C16 VP VN 8.850901f
C17 VP VDD2 0.575213f
C18 VTAIL VDD1 11.802f
C19 B VN 1.30496f
C20 VDD2 B 2.8077f
C21 VDD2 VSUBS 2.21171f
C22 VDD1 VSUBS 2.012365f
C23 VTAIL VSUBS 1.383721f
C24 VN VSUBS 7.66886f
C25 VP VSUBS 4.258379f
C26 B VSUBS 5.538363f
C27 w_n4402_n3976# VSUBS 0.214624p
C28 VDD2.t3 VSUBS 3.6707f
C29 VDD2.t7 VSUBS 0.344764f
C30 VDD2.t8 VSUBS 0.344764f
C31 VDD2.n0 VSUBS 2.80132f
C32 VDD2.n1 VSUBS 1.70307f
C33 VDD2.t2 VSUBS 0.344764f
C34 VDD2.t5 VSUBS 0.344764f
C35 VDD2.n2 VSUBS 2.82497f
C36 VDD2.n3 VSUBS 3.85697f
C37 VDD2.t6 VSUBS 3.64163f
C38 VDD2.n4 VSUBS 4.20112f
C39 VDD2.t9 VSUBS 0.344764f
C40 VDD2.t0 VSUBS 0.344764f
C41 VDD2.n5 VSUBS 2.80133f
C42 VDD2.n6 VSUBS 0.846479f
C43 VDD2.t1 VSUBS 0.344764f
C44 VDD2.t4 VSUBS 0.344764f
C45 VDD2.n7 VSUBS 2.82491f
C46 VN.n0 VSUBS 0.035505f
C47 VN.t4 VSUBS 2.8083f
C48 VN.n1 VSUBS 0.036169f
C49 VN.n2 VSUBS 0.026932f
C50 VN.t7 VSUBS 2.8083f
C51 VN.n3 VSUBS 0.981974f
C52 VN.n4 VSUBS 0.026932f
C53 VN.n5 VSUBS 0.050654f
C54 VN.n6 VSUBS 0.026932f
C55 VN.t1 VSUBS 2.8083f
C56 VN.n7 VSUBS 0.050654f
C57 VN.n8 VSUBS 0.026932f
C58 VN.t2 VSUBS 2.8083f
C59 VN.n9 VSUBS 1.06379f
C60 VN.t6 VSUBS 3.02748f
C61 VN.n10 VSUBS 1.03151f
C62 VN.n11 VSUBS 0.258398f
C63 VN.n12 VSUBS 0.043039f
C64 VN.n13 VSUBS 0.054106f
C65 VN.n14 VSUBS 0.023483f
C66 VN.n15 VSUBS 0.026932f
C67 VN.n16 VSUBS 0.026932f
C68 VN.n17 VSUBS 0.026932f
C69 VN.n18 VSUBS 0.049943f
C70 VN.n19 VSUBS 1.00726f
C71 VN.n20 VSUBS 0.049943f
C72 VN.n21 VSUBS 0.026932f
C73 VN.n22 VSUBS 0.026932f
C74 VN.n23 VSUBS 0.026932f
C75 VN.n24 VSUBS 0.023483f
C76 VN.n25 VSUBS 0.054106f
C77 VN.n26 VSUBS 0.043039f
C78 VN.n27 VSUBS 0.026932f
C79 VN.n28 VSUBS 0.026932f
C80 VN.n29 VSUBS 0.032191f
C81 VN.n30 VSUBS 0.049943f
C82 VN.n31 VSUBS 0.04213f
C83 VN.n32 VSUBS 0.026932f
C84 VN.n33 VSUBS 0.026932f
C85 VN.n34 VSUBS 0.026932f
C86 VN.n35 VSUBS 0.049943f
C87 VN.n36 VSUBS 0.036136f
C88 VN.n37 VSUBS 1.07041f
C89 VN.n38 VSUBS 0.042677f
C90 VN.n39 VSUBS 0.035505f
C91 VN.t3 VSUBS 2.8083f
C92 VN.n40 VSUBS 0.036169f
C93 VN.n41 VSUBS 0.026932f
C94 VN.t0 VSUBS 2.8083f
C95 VN.n42 VSUBS 0.981974f
C96 VN.n43 VSUBS 0.026932f
C97 VN.n44 VSUBS 0.050654f
C98 VN.n45 VSUBS 0.026932f
C99 VN.t9 VSUBS 2.8083f
C100 VN.n46 VSUBS 0.050654f
C101 VN.n47 VSUBS 0.026932f
C102 VN.t8 VSUBS 2.8083f
C103 VN.n48 VSUBS 1.06379f
C104 VN.t5 VSUBS 3.02748f
C105 VN.n49 VSUBS 1.03151f
C106 VN.n50 VSUBS 0.258398f
C107 VN.n51 VSUBS 0.043039f
C108 VN.n52 VSUBS 0.054106f
C109 VN.n53 VSUBS 0.023483f
C110 VN.n54 VSUBS 0.026932f
C111 VN.n55 VSUBS 0.026932f
C112 VN.n56 VSUBS 0.026932f
C113 VN.n57 VSUBS 0.049943f
C114 VN.n58 VSUBS 1.00726f
C115 VN.n59 VSUBS 0.049943f
C116 VN.n60 VSUBS 0.026932f
C117 VN.n61 VSUBS 0.026932f
C118 VN.n62 VSUBS 0.026932f
C119 VN.n63 VSUBS 0.023483f
C120 VN.n64 VSUBS 0.054106f
C121 VN.n65 VSUBS 0.043039f
C122 VN.n66 VSUBS 0.026932f
C123 VN.n67 VSUBS 0.026932f
C124 VN.n68 VSUBS 0.032191f
C125 VN.n69 VSUBS 0.049943f
C126 VN.n70 VSUBS 0.04213f
C127 VN.n71 VSUBS 0.026932f
C128 VN.n72 VSUBS 0.026932f
C129 VN.n73 VSUBS 0.026932f
C130 VN.n74 VSUBS 0.049943f
C131 VN.n75 VSUBS 0.036136f
C132 VN.n76 VSUBS 1.07041f
C133 VN.n77 VSUBS 1.73403f
C134 B.n0 VSUBS 0.007672f
C135 B.n1 VSUBS 0.007672f
C136 B.n2 VSUBS 0.011346f
C137 B.n3 VSUBS 0.008695f
C138 B.n4 VSUBS 0.008695f
C139 B.n5 VSUBS 0.008695f
C140 B.n6 VSUBS 0.008695f
C141 B.n7 VSUBS 0.008695f
C142 B.n8 VSUBS 0.008695f
C143 B.n9 VSUBS 0.008695f
C144 B.n10 VSUBS 0.008695f
C145 B.n11 VSUBS 0.008695f
C146 B.n12 VSUBS 0.008695f
C147 B.n13 VSUBS 0.008695f
C148 B.n14 VSUBS 0.008695f
C149 B.n15 VSUBS 0.008695f
C150 B.n16 VSUBS 0.008695f
C151 B.n17 VSUBS 0.008695f
C152 B.n18 VSUBS 0.008695f
C153 B.n19 VSUBS 0.008695f
C154 B.n20 VSUBS 0.008695f
C155 B.n21 VSUBS 0.008695f
C156 B.n22 VSUBS 0.008695f
C157 B.n23 VSUBS 0.008695f
C158 B.n24 VSUBS 0.008695f
C159 B.n25 VSUBS 0.008695f
C160 B.n26 VSUBS 0.008695f
C161 B.n27 VSUBS 0.008695f
C162 B.n28 VSUBS 0.008695f
C163 B.n29 VSUBS 0.008695f
C164 B.n30 VSUBS 0.008695f
C165 B.n31 VSUBS 0.020657f
C166 B.n32 VSUBS 0.008695f
C167 B.n33 VSUBS 0.008695f
C168 B.n34 VSUBS 0.008695f
C169 B.n35 VSUBS 0.008695f
C170 B.n36 VSUBS 0.008695f
C171 B.n37 VSUBS 0.008695f
C172 B.n38 VSUBS 0.008695f
C173 B.n39 VSUBS 0.008695f
C174 B.n40 VSUBS 0.008695f
C175 B.n41 VSUBS 0.008695f
C176 B.n42 VSUBS 0.008695f
C177 B.n43 VSUBS 0.008695f
C178 B.n44 VSUBS 0.008695f
C179 B.n45 VSUBS 0.008695f
C180 B.n46 VSUBS 0.008695f
C181 B.n47 VSUBS 0.008695f
C182 B.n48 VSUBS 0.008695f
C183 B.n49 VSUBS 0.008695f
C184 B.n50 VSUBS 0.008695f
C185 B.n51 VSUBS 0.008695f
C186 B.n52 VSUBS 0.008695f
C187 B.n53 VSUBS 0.008695f
C188 B.n54 VSUBS 0.008695f
C189 B.n55 VSUBS 0.008695f
C190 B.n56 VSUBS 0.006009f
C191 B.n57 VSUBS 0.008695f
C192 B.t1 VSUBS 0.622f
C193 B.t2 VSUBS 0.647999f
C194 B.t0 VSUBS 2.11768f
C195 B.n58 VSUBS 0.342507f
C196 B.n59 VSUBS 0.089064f
C197 B.n60 VSUBS 0.020144f
C198 B.n61 VSUBS 0.008695f
C199 B.n62 VSUBS 0.008695f
C200 B.n63 VSUBS 0.008695f
C201 B.n64 VSUBS 0.008695f
C202 B.t7 VSUBS 0.621982f
C203 B.t8 VSUBS 0.647984f
C204 B.t6 VSUBS 2.11768f
C205 B.n65 VSUBS 0.342522f
C206 B.n66 VSUBS 0.089082f
C207 B.n67 VSUBS 0.008695f
C208 B.n68 VSUBS 0.008695f
C209 B.n69 VSUBS 0.008695f
C210 B.n70 VSUBS 0.008695f
C211 B.n71 VSUBS 0.008695f
C212 B.n72 VSUBS 0.008695f
C213 B.n73 VSUBS 0.008695f
C214 B.n74 VSUBS 0.008695f
C215 B.n75 VSUBS 0.008695f
C216 B.n76 VSUBS 0.008695f
C217 B.n77 VSUBS 0.008695f
C218 B.n78 VSUBS 0.008695f
C219 B.n79 VSUBS 0.008695f
C220 B.n80 VSUBS 0.008695f
C221 B.n81 VSUBS 0.008695f
C222 B.n82 VSUBS 0.008695f
C223 B.n83 VSUBS 0.008695f
C224 B.n84 VSUBS 0.008695f
C225 B.n85 VSUBS 0.008695f
C226 B.n86 VSUBS 0.008695f
C227 B.n87 VSUBS 0.008695f
C228 B.n88 VSUBS 0.008695f
C229 B.n89 VSUBS 0.008695f
C230 B.n90 VSUBS 0.008695f
C231 B.n91 VSUBS 0.020657f
C232 B.n92 VSUBS 0.008695f
C233 B.n93 VSUBS 0.008695f
C234 B.n94 VSUBS 0.008695f
C235 B.n95 VSUBS 0.008695f
C236 B.n96 VSUBS 0.008695f
C237 B.n97 VSUBS 0.008695f
C238 B.n98 VSUBS 0.008695f
C239 B.n99 VSUBS 0.008695f
C240 B.n100 VSUBS 0.008695f
C241 B.n101 VSUBS 0.008695f
C242 B.n102 VSUBS 0.008695f
C243 B.n103 VSUBS 0.008695f
C244 B.n104 VSUBS 0.008695f
C245 B.n105 VSUBS 0.008695f
C246 B.n106 VSUBS 0.008695f
C247 B.n107 VSUBS 0.008695f
C248 B.n108 VSUBS 0.008695f
C249 B.n109 VSUBS 0.008695f
C250 B.n110 VSUBS 0.008695f
C251 B.n111 VSUBS 0.008695f
C252 B.n112 VSUBS 0.008695f
C253 B.n113 VSUBS 0.008695f
C254 B.n114 VSUBS 0.008695f
C255 B.n115 VSUBS 0.008695f
C256 B.n116 VSUBS 0.008695f
C257 B.n117 VSUBS 0.008695f
C258 B.n118 VSUBS 0.008695f
C259 B.n119 VSUBS 0.008695f
C260 B.n120 VSUBS 0.008695f
C261 B.n121 VSUBS 0.008695f
C262 B.n122 VSUBS 0.008695f
C263 B.n123 VSUBS 0.008695f
C264 B.n124 VSUBS 0.008695f
C265 B.n125 VSUBS 0.008695f
C266 B.n126 VSUBS 0.008695f
C267 B.n127 VSUBS 0.008695f
C268 B.n128 VSUBS 0.008695f
C269 B.n129 VSUBS 0.008695f
C270 B.n130 VSUBS 0.008695f
C271 B.n131 VSUBS 0.008695f
C272 B.n132 VSUBS 0.008695f
C273 B.n133 VSUBS 0.008695f
C274 B.n134 VSUBS 0.008695f
C275 B.n135 VSUBS 0.008695f
C276 B.n136 VSUBS 0.008695f
C277 B.n137 VSUBS 0.008695f
C278 B.n138 VSUBS 0.008695f
C279 B.n139 VSUBS 0.008695f
C280 B.n140 VSUBS 0.008695f
C281 B.n141 VSUBS 0.008695f
C282 B.n142 VSUBS 0.008695f
C283 B.n143 VSUBS 0.008695f
C284 B.n144 VSUBS 0.008695f
C285 B.n145 VSUBS 0.008695f
C286 B.n146 VSUBS 0.008695f
C287 B.n147 VSUBS 0.008695f
C288 B.n148 VSUBS 0.008695f
C289 B.n149 VSUBS 0.008695f
C290 B.n150 VSUBS 0.019236f
C291 B.n151 VSUBS 0.008695f
C292 B.n152 VSUBS 0.008695f
C293 B.n153 VSUBS 0.008695f
C294 B.n154 VSUBS 0.008695f
C295 B.n155 VSUBS 0.008695f
C296 B.n156 VSUBS 0.008695f
C297 B.n157 VSUBS 0.008695f
C298 B.n158 VSUBS 0.008695f
C299 B.n159 VSUBS 0.008695f
C300 B.n160 VSUBS 0.008695f
C301 B.n161 VSUBS 0.008695f
C302 B.n162 VSUBS 0.008695f
C303 B.n163 VSUBS 0.008695f
C304 B.n164 VSUBS 0.008695f
C305 B.n165 VSUBS 0.008695f
C306 B.n166 VSUBS 0.008695f
C307 B.n167 VSUBS 0.008695f
C308 B.n168 VSUBS 0.008695f
C309 B.n169 VSUBS 0.008695f
C310 B.n170 VSUBS 0.008695f
C311 B.n171 VSUBS 0.008695f
C312 B.n172 VSUBS 0.008695f
C313 B.n173 VSUBS 0.008695f
C314 B.n174 VSUBS 0.008695f
C315 B.n175 VSUBS 0.008695f
C316 B.n176 VSUBS 0.008695f
C317 B.t5 VSUBS 0.621982f
C318 B.t4 VSUBS 0.647984f
C319 B.t3 VSUBS 2.11768f
C320 B.n177 VSUBS 0.342522f
C321 B.n178 VSUBS 0.089082f
C322 B.n179 VSUBS 0.008695f
C323 B.n180 VSUBS 0.008695f
C324 B.n181 VSUBS 0.008695f
C325 B.n182 VSUBS 0.008695f
C326 B.t11 VSUBS 0.622f
C327 B.t10 VSUBS 0.647999f
C328 B.t9 VSUBS 2.11768f
C329 B.n183 VSUBS 0.342507f
C330 B.n184 VSUBS 0.089064f
C331 B.n185 VSUBS 0.008695f
C332 B.n186 VSUBS 0.008695f
C333 B.n187 VSUBS 0.008695f
C334 B.n188 VSUBS 0.008695f
C335 B.n189 VSUBS 0.008695f
C336 B.n190 VSUBS 0.008695f
C337 B.n191 VSUBS 0.008695f
C338 B.n192 VSUBS 0.008695f
C339 B.n193 VSUBS 0.008695f
C340 B.n194 VSUBS 0.008695f
C341 B.n195 VSUBS 0.008695f
C342 B.n196 VSUBS 0.008695f
C343 B.n197 VSUBS 0.008695f
C344 B.n198 VSUBS 0.008695f
C345 B.n199 VSUBS 0.008695f
C346 B.n200 VSUBS 0.008695f
C347 B.n201 VSUBS 0.008695f
C348 B.n202 VSUBS 0.008695f
C349 B.n203 VSUBS 0.008695f
C350 B.n204 VSUBS 0.008695f
C351 B.n205 VSUBS 0.008695f
C352 B.n206 VSUBS 0.008695f
C353 B.n207 VSUBS 0.008695f
C354 B.n208 VSUBS 0.008695f
C355 B.n209 VSUBS 0.008695f
C356 B.n210 VSUBS 0.019236f
C357 B.n211 VSUBS 0.008695f
C358 B.n212 VSUBS 0.008695f
C359 B.n213 VSUBS 0.008695f
C360 B.n214 VSUBS 0.008695f
C361 B.n215 VSUBS 0.008695f
C362 B.n216 VSUBS 0.008695f
C363 B.n217 VSUBS 0.008695f
C364 B.n218 VSUBS 0.008695f
C365 B.n219 VSUBS 0.008695f
C366 B.n220 VSUBS 0.008695f
C367 B.n221 VSUBS 0.008695f
C368 B.n222 VSUBS 0.008695f
C369 B.n223 VSUBS 0.008695f
C370 B.n224 VSUBS 0.008695f
C371 B.n225 VSUBS 0.008695f
C372 B.n226 VSUBS 0.008695f
C373 B.n227 VSUBS 0.008695f
C374 B.n228 VSUBS 0.008695f
C375 B.n229 VSUBS 0.008695f
C376 B.n230 VSUBS 0.008695f
C377 B.n231 VSUBS 0.008695f
C378 B.n232 VSUBS 0.008695f
C379 B.n233 VSUBS 0.008695f
C380 B.n234 VSUBS 0.008695f
C381 B.n235 VSUBS 0.008695f
C382 B.n236 VSUBS 0.008695f
C383 B.n237 VSUBS 0.008695f
C384 B.n238 VSUBS 0.008695f
C385 B.n239 VSUBS 0.008695f
C386 B.n240 VSUBS 0.008695f
C387 B.n241 VSUBS 0.008695f
C388 B.n242 VSUBS 0.008695f
C389 B.n243 VSUBS 0.008695f
C390 B.n244 VSUBS 0.008695f
C391 B.n245 VSUBS 0.008695f
C392 B.n246 VSUBS 0.008695f
C393 B.n247 VSUBS 0.008695f
C394 B.n248 VSUBS 0.008695f
C395 B.n249 VSUBS 0.008695f
C396 B.n250 VSUBS 0.008695f
C397 B.n251 VSUBS 0.008695f
C398 B.n252 VSUBS 0.008695f
C399 B.n253 VSUBS 0.008695f
C400 B.n254 VSUBS 0.008695f
C401 B.n255 VSUBS 0.008695f
C402 B.n256 VSUBS 0.008695f
C403 B.n257 VSUBS 0.008695f
C404 B.n258 VSUBS 0.008695f
C405 B.n259 VSUBS 0.008695f
C406 B.n260 VSUBS 0.008695f
C407 B.n261 VSUBS 0.008695f
C408 B.n262 VSUBS 0.008695f
C409 B.n263 VSUBS 0.008695f
C410 B.n264 VSUBS 0.008695f
C411 B.n265 VSUBS 0.008695f
C412 B.n266 VSUBS 0.008695f
C413 B.n267 VSUBS 0.008695f
C414 B.n268 VSUBS 0.008695f
C415 B.n269 VSUBS 0.008695f
C416 B.n270 VSUBS 0.008695f
C417 B.n271 VSUBS 0.008695f
C418 B.n272 VSUBS 0.008695f
C419 B.n273 VSUBS 0.008695f
C420 B.n274 VSUBS 0.008695f
C421 B.n275 VSUBS 0.008695f
C422 B.n276 VSUBS 0.008695f
C423 B.n277 VSUBS 0.008695f
C424 B.n278 VSUBS 0.008695f
C425 B.n279 VSUBS 0.008695f
C426 B.n280 VSUBS 0.008695f
C427 B.n281 VSUBS 0.008695f
C428 B.n282 VSUBS 0.008695f
C429 B.n283 VSUBS 0.008695f
C430 B.n284 VSUBS 0.008695f
C431 B.n285 VSUBS 0.008695f
C432 B.n286 VSUBS 0.008695f
C433 B.n287 VSUBS 0.008695f
C434 B.n288 VSUBS 0.008695f
C435 B.n289 VSUBS 0.008695f
C436 B.n290 VSUBS 0.008695f
C437 B.n291 VSUBS 0.008695f
C438 B.n292 VSUBS 0.008695f
C439 B.n293 VSUBS 0.008695f
C440 B.n294 VSUBS 0.008695f
C441 B.n295 VSUBS 0.008695f
C442 B.n296 VSUBS 0.008695f
C443 B.n297 VSUBS 0.008695f
C444 B.n298 VSUBS 0.008695f
C445 B.n299 VSUBS 0.008695f
C446 B.n300 VSUBS 0.008695f
C447 B.n301 VSUBS 0.008695f
C448 B.n302 VSUBS 0.008695f
C449 B.n303 VSUBS 0.008695f
C450 B.n304 VSUBS 0.008695f
C451 B.n305 VSUBS 0.008695f
C452 B.n306 VSUBS 0.008695f
C453 B.n307 VSUBS 0.008695f
C454 B.n308 VSUBS 0.008695f
C455 B.n309 VSUBS 0.008695f
C456 B.n310 VSUBS 0.008695f
C457 B.n311 VSUBS 0.008695f
C458 B.n312 VSUBS 0.008695f
C459 B.n313 VSUBS 0.008695f
C460 B.n314 VSUBS 0.008695f
C461 B.n315 VSUBS 0.008695f
C462 B.n316 VSUBS 0.008695f
C463 B.n317 VSUBS 0.008695f
C464 B.n318 VSUBS 0.008695f
C465 B.n319 VSUBS 0.008695f
C466 B.n320 VSUBS 0.008695f
C467 B.n321 VSUBS 0.008695f
C468 B.n322 VSUBS 0.008695f
C469 B.n323 VSUBS 0.019236f
C470 B.n324 VSUBS 0.020657f
C471 B.n325 VSUBS 0.020657f
C472 B.n326 VSUBS 0.008695f
C473 B.n327 VSUBS 0.008695f
C474 B.n328 VSUBS 0.008695f
C475 B.n329 VSUBS 0.008695f
C476 B.n330 VSUBS 0.008695f
C477 B.n331 VSUBS 0.008695f
C478 B.n332 VSUBS 0.008695f
C479 B.n333 VSUBS 0.008695f
C480 B.n334 VSUBS 0.008695f
C481 B.n335 VSUBS 0.008695f
C482 B.n336 VSUBS 0.008695f
C483 B.n337 VSUBS 0.008695f
C484 B.n338 VSUBS 0.008695f
C485 B.n339 VSUBS 0.008695f
C486 B.n340 VSUBS 0.008695f
C487 B.n341 VSUBS 0.008695f
C488 B.n342 VSUBS 0.008695f
C489 B.n343 VSUBS 0.008695f
C490 B.n344 VSUBS 0.008695f
C491 B.n345 VSUBS 0.008695f
C492 B.n346 VSUBS 0.008695f
C493 B.n347 VSUBS 0.008695f
C494 B.n348 VSUBS 0.008695f
C495 B.n349 VSUBS 0.008695f
C496 B.n350 VSUBS 0.008695f
C497 B.n351 VSUBS 0.008695f
C498 B.n352 VSUBS 0.008695f
C499 B.n353 VSUBS 0.008695f
C500 B.n354 VSUBS 0.008695f
C501 B.n355 VSUBS 0.008695f
C502 B.n356 VSUBS 0.008695f
C503 B.n357 VSUBS 0.008695f
C504 B.n358 VSUBS 0.008695f
C505 B.n359 VSUBS 0.008695f
C506 B.n360 VSUBS 0.008695f
C507 B.n361 VSUBS 0.008695f
C508 B.n362 VSUBS 0.008695f
C509 B.n363 VSUBS 0.008695f
C510 B.n364 VSUBS 0.008695f
C511 B.n365 VSUBS 0.008695f
C512 B.n366 VSUBS 0.008695f
C513 B.n367 VSUBS 0.008695f
C514 B.n368 VSUBS 0.008695f
C515 B.n369 VSUBS 0.008695f
C516 B.n370 VSUBS 0.008695f
C517 B.n371 VSUBS 0.008695f
C518 B.n372 VSUBS 0.008695f
C519 B.n373 VSUBS 0.008695f
C520 B.n374 VSUBS 0.008695f
C521 B.n375 VSUBS 0.008695f
C522 B.n376 VSUBS 0.008695f
C523 B.n377 VSUBS 0.008695f
C524 B.n378 VSUBS 0.008695f
C525 B.n379 VSUBS 0.008695f
C526 B.n380 VSUBS 0.008695f
C527 B.n381 VSUBS 0.008695f
C528 B.n382 VSUBS 0.008695f
C529 B.n383 VSUBS 0.008695f
C530 B.n384 VSUBS 0.008695f
C531 B.n385 VSUBS 0.008695f
C532 B.n386 VSUBS 0.008695f
C533 B.n387 VSUBS 0.008695f
C534 B.n388 VSUBS 0.008695f
C535 B.n389 VSUBS 0.008695f
C536 B.n390 VSUBS 0.008695f
C537 B.n391 VSUBS 0.008695f
C538 B.n392 VSUBS 0.008695f
C539 B.n393 VSUBS 0.008695f
C540 B.n394 VSUBS 0.008695f
C541 B.n395 VSUBS 0.008695f
C542 B.n396 VSUBS 0.008695f
C543 B.n397 VSUBS 0.008695f
C544 B.n398 VSUBS 0.008695f
C545 B.n399 VSUBS 0.008695f
C546 B.n400 VSUBS 0.006009f
C547 B.n401 VSUBS 0.020144f
C548 B.n402 VSUBS 0.007032f
C549 B.n403 VSUBS 0.008695f
C550 B.n404 VSUBS 0.008695f
C551 B.n405 VSUBS 0.008695f
C552 B.n406 VSUBS 0.008695f
C553 B.n407 VSUBS 0.008695f
C554 B.n408 VSUBS 0.008695f
C555 B.n409 VSUBS 0.008695f
C556 B.n410 VSUBS 0.008695f
C557 B.n411 VSUBS 0.008695f
C558 B.n412 VSUBS 0.008695f
C559 B.n413 VSUBS 0.008695f
C560 B.n414 VSUBS 0.007032f
C561 B.n415 VSUBS 0.020144f
C562 B.n416 VSUBS 0.006009f
C563 B.n417 VSUBS 0.008695f
C564 B.n418 VSUBS 0.008695f
C565 B.n419 VSUBS 0.008695f
C566 B.n420 VSUBS 0.008695f
C567 B.n421 VSUBS 0.008695f
C568 B.n422 VSUBS 0.008695f
C569 B.n423 VSUBS 0.008695f
C570 B.n424 VSUBS 0.008695f
C571 B.n425 VSUBS 0.008695f
C572 B.n426 VSUBS 0.008695f
C573 B.n427 VSUBS 0.008695f
C574 B.n428 VSUBS 0.008695f
C575 B.n429 VSUBS 0.008695f
C576 B.n430 VSUBS 0.008695f
C577 B.n431 VSUBS 0.008695f
C578 B.n432 VSUBS 0.008695f
C579 B.n433 VSUBS 0.008695f
C580 B.n434 VSUBS 0.008695f
C581 B.n435 VSUBS 0.008695f
C582 B.n436 VSUBS 0.008695f
C583 B.n437 VSUBS 0.008695f
C584 B.n438 VSUBS 0.008695f
C585 B.n439 VSUBS 0.008695f
C586 B.n440 VSUBS 0.008695f
C587 B.n441 VSUBS 0.008695f
C588 B.n442 VSUBS 0.008695f
C589 B.n443 VSUBS 0.008695f
C590 B.n444 VSUBS 0.008695f
C591 B.n445 VSUBS 0.008695f
C592 B.n446 VSUBS 0.008695f
C593 B.n447 VSUBS 0.008695f
C594 B.n448 VSUBS 0.008695f
C595 B.n449 VSUBS 0.008695f
C596 B.n450 VSUBS 0.008695f
C597 B.n451 VSUBS 0.008695f
C598 B.n452 VSUBS 0.008695f
C599 B.n453 VSUBS 0.008695f
C600 B.n454 VSUBS 0.008695f
C601 B.n455 VSUBS 0.008695f
C602 B.n456 VSUBS 0.008695f
C603 B.n457 VSUBS 0.008695f
C604 B.n458 VSUBS 0.008695f
C605 B.n459 VSUBS 0.008695f
C606 B.n460 VSUBS 0.008695f
C607 B.n461 VSUBS 0.008695f
C608 B.n462 VSUBS 0.008695f
C609 B.n463 VSUBS 0.008695f
C610 B.n464 VSUBS 0.008695f
C611 B.n465 VSUBS 0.008695f
C612 B.n466 VSUBS 0.008695f
C613 B.n467 VSUBS 0.008695f
C614 B.n468 VSUBS 0.008695f
C615 B.n469 VSUBS 0.008695f
C616 B.n470 VSUBS 0.008695f
C617 B.n471 VSUBS 0.008695f
C618 B.n472 VSUBS 0.008695f
C619 B.n473 VSUBS 0.008695f
C620 B.n474 VSUBS 0.008695f
C621 B.n475 VSUBS 0.008695f
C622 B.n476 VSUBS 0.008695f
C623 B.n477 VSUBS 0.008695f
C624 B.n478 VSUBS 0.008695f
C625 B.n479 VSUBS 0.008695f
C626 B.n480 VSUBS 0.008695f
C627 B.n481 VSUBS 0.008695f
C628 B.n482 VSUBS 0.008695f
C629 B.n483 VSUBS 0.008695f
C630 B.n484 VSUBS 0.008695f
C631 B.n485 VSUBS 0.008695f
C632 B.n486 VSUBS 0.008695f
C633 B.n487 VSUBS 0.008695f
C634 B.n488 VSUBS 0.008695f
C635 B.n489 VSUBS 0.008695f
C636 B.n490 VSUBS 0.008695f
C637 B.n491 VSUBS 0.020657f
C638 B.n492 VSUBS 0.019598f
C639 B.n493 VSUBS 0.020295f
C640 B.n494 VSUBS 0.008695f
C641 B.n495 VSUBS 0.008695f
C642 B.n496 VSUBS 0.008695f
C643 B.n497 VSUBS 0.008695f
C644 B.n498 VSUBS 0.008695f
C645 B.n499 VSUBS 0.008695f
C646 B.n500 VSUBS 0.008695f
C647 B.n501 VSUBS 0.008695f
C648 B.n502 VSUBS 0.008695f
C649 B.n503 VSUBS 0.008695f
C650 B.n504 VSUBS 0.008695f
C651 B.n505 VSUBS 0.008695f
C652 B.n506 VSUBS 0.008695f
C653 B.n507 VSUBS 0.008695f
C654 B.n508 VSUBS 0.008695f
C655 B.n509 VSUBS 0.008695f
C656 B.n510 VSUBS 0.008695f
C657 B.n511 VSUBS 0.008695f
C658 B.n512 VSUBS 0.008695f
C659 B.n513 VSUBS 0.008695f
C660 B.n514 VSUBS 0.008695f
C661 B.n515 VSUBS 0.008695f
C662 B.n516 VSUBS 0.008695f
C663 B.n517 VSUBS 0.008695f
C664 B.n518 VSUBS 0.008695f
C665 B.n519 VSUBS 0.008695f
C666 B.n520 VSUBS 0.008695f
C667 B.n521 VSUBS 0.008695f
C668 B.n522 VSUBS 0.008695f
C669 B.n523 VSUBS 0.008695f
C670 B.n524 VSUBS 0.008695f
C671 B.n525 VSUBS 0.008695f
C672 B.n526 VSUBS 0.008695f
C673 B.n527 VSUBS 0.008695f
C674 B.n528 VSUBS 0.008695f
C675 B.n529 VSUBS 0.008695f
C676 B.n530 VSUBS 0.008695f
C677 B.n531 VSUBS 0.008695f
C678 B.n532 VSUBS 0.008695f
C679 B.n533 VSUBS 0.008695f
C680 B.n534 VSUBS 0.008695f
C681 B.n535 VSUBS 0.008695f
C682 B.n536 VSUBS 0.008695f
C683 B.n537 VSUBS 0.008695f
C684 B.n538 VSUBS 0.008695f
C685 B.n539 VSUBS 0.008695f
C686 B.n540 VSUBS 0.008695f
C687 B.n541 VSUBS 0.008695f
C688 B.n542 VSUBS 0.008695f
C689 B.n543 VSUBS 0.008695f
C690 B.n544 VSUBS 0.008695f
C691 B.n545 VSUBS 0.008695f
C692 B.n546 VSUBS 0.008695f
C693 B.n547 VSUBS 0.008695f
C694 B.n548 VSUBS 0.008695f
C695 B.n549 VSUBS 0.008695f
C696 B.n550 VSUBS 0.008695f
C697 B.n551 VSUBS 0.008695f
C698 B.n552 VSUBS 0.008695f
C699 B.n553 VSUBS 0.008695f
C700 B.n554 VSUBS 0.008695f
C701 B.n555 VSUBS 0.008695f
C702 B.n556 VSUBS 0.008695f
C703 B.n557 VSUBS 0.008695f
C704 B.n558 VSUBS 0.008695f
C705 B.n559 VSUBS 0.008695f
C706 B.n560 VSUBS 0.008695f
C707 B.n561 VSUBS 0.008695f
C708 B.n562 VSUBS 0.008695f
C709 B.n563 VSUBS 0.008695f
C710 B.n564 VSUBS 0.008695f
C711 B.n565 VSUBS 0.008695f
C712 B.n566 VSUBS 0.008695f
C713 B.n567 VSUBS 0.008695f
C714 B.n568 VSUBS 0.008695f
C715 B.n569 VSUBS 0.008695f
C716 B.n570 VSUBS 0.008695f
C717 B.n571 VSUBS 0.008695f
C718 B.n572 VSUBS 0.008695f
C719 B.n573 VSUBS 0.008695f
C720 B.n574 VSUBS 0.008695f
C721 B.n575 VSUBS 0.008695f
C722 B.n576 VSUBS 0.008695f
C723 B.n577 VSUBS 0.008695f
C724 B.n578 VSUBS 0.008695f
C725 B.n579 VSUBS 0.008695f
C726 B.n580 VSUBS 0.008695f
C727 B.n581 VSUBS 0.008695f
C728 B.n582 VSUBS 0.008695f
C729 B.n583 VSUBS 0.008695f
C730 B.n584 VSUBS 0.008695f
C731 B.n585 VSUBS 0.008695f
C732 B.n586 VSUBS 0.008695f
C733 B.n587 VSUBS 0.008695f
C734 B.n588 VSUBS 0.008695f
C735 B.n589 VSUBS 0.008695f
C736 B.n590 VSUBS 0.008695f
C737 B.n591 VSUBS 0.008695f
C738 B.n592 VSUBS 0.008695f
C739 B.n593 VSUBS 0.008695f
C740 B.n594 VSUBS 0.008695f
C741 B.n595 VSUBS 0.008695f
C742 B.n596 VSUBS 0.008695f
C743 B.n597 VSUBS 0.008695f
C744 B.n598 VSUBS 0.008695f
C745 B.n599 VSUBS 0.008695f
C746 B.n600 VSUBS 0.008695f
C747 B.n601 VSUBS 0.008695f
C748 B.n602 VSUBS 0.008695f
C749 B.n603 VSUBS 0.008695f
C750 B.n604 VSUBS 0.008695f
C751 B.n605 VSUBS 0.008695f
C752 B.n606 VSUBS 0.008695f
C753 B.n607 VSUBS 0.008695f
C754 B.n608 VSUBS 0.008695f
C755 B.n609 VSUBS 0.008695f
C756 B.n610 VSUBS 0.008695f
C757 B.n611 VSUBS 0.008695f
C758 B.n612 VSUBS 0.008695f
C759 B.n613 VSUBS 0.008695f
C760 B.n614 VSUBS 0.008695f
C761 B.n615 VSUBS 0.008695f
C762 B.n616 VSUBS 0.008695f
C763 B.n617 VSUBS 0.008695f
C764 B.n618 VSUBS 0.008695f
C765 B.n619 VSUBS 0.008695f
C766 B.n620 VSUBS 0.008695f
C767 B.n621 VSUBS 0.008695f
C768 B.n622 VSUBS 0.008695f
C769 B.n623 VSUBS 0.008695f
C770 B.n624 VSUBS 0.008695f
C771 B.n625 VSUBS 0.008695f
C772 B.n626 VSUBS 0.008695f
C773 B.n627 VSUBS 0.008695f
C774 B.n628 VSUBS 0.008695f
C775 B.n629 VSUBS 0.008695f
C776 B.n630 VSUBS 0.008695f
C777 B.n631 VSUBS 0.008695f
C778 B.n632 VSUBS 0.008695f
C779 B.n633 VSUBS 0.008695f
C780 B.n634 VSUBS 0.008695f
C781 B.n635 VSUBS 0.008695f
C782 B.n636 VSUBS 0.008695f
C783 B.n637 VSUBS 0.008695f
C784 B.n638 VSUBS 0.008695f
C785 B.n639 VSUBS 0.008695f
C786 B.n640 VSUBS 0.008695f
C787 B.n641 VSUBS 0.008695f
C788 B.n642 VSUBS 0.008695f
C789 B.n643 VSUBS 0.008695f
C790 B.n644 VSUBS 0.008695f
C791 B.n645 VSUBS 0.008695f
C792 B.n646 VSUBS 0.008695f
C793 B.n647 VSUBS 0.008695f
C794 B.n648 VSUBS 0.008695f
C795 B.n649 VSUBS 0.008695f
C796 B.n650 VSUBS 0.008695f
C797 B.n651 VSUBS 0.008695f
C798 B.n652 VSUBS 0.008695f
C799 B.n653 VSUBS 0.008695f
C800 B.n654 VSUBS 0.008695f
C801 B.n655 VSUBS 0.008695f
C802 B.n656 VSUBS 0.008695f
C803 B.n657 VSUBS 0.008695f
C804 B.n658 VSUBS 0.008695f
C805 B.n659 VSUBS 0.008695f
C806 B.n660 VSUBS 0.008695f
C807 B.n661 VSUBS 0.008695f
C808 B.n662 VSUBS 0.008695f
C809 B.n663 VSUBS 0.008695f
C810 B.n664 VSUBS 0.008695f
C811 B.n665 VSUBS 0.008695f
C812 B.n666 VSUBS 0.008695f
C813 B.n667 VSUBS 0.008695f
C814 B.n668 VSUBS 0.019236f
C815 B.n669 VSUBS 0.019236f
C816 B.n670 VSUBS 0.020657f
C817 B.n671 VSUBS 0.008695f
C818 B.n672 VSUBS 0.008695f
C819 B.n673 VSUBS 0.008695f
C820 B.n674 VSUBS 0.008695f
C821 B.n675 VSUBS 0.008695f
C822 B.n676 VSUBS 0.008695f
C823 B.n677 VSUBS 0.008695f
C824 B.n678 VSUBS 0.008695f
C825 B.n679 VSUBS 0.008695f
C826 B.n680 VSUBS 0.008695f
C827 B.n681 VSUBS 0.008695f
C828 B.n682 VSUBS 0.008695f
C829 B.n683 VSUBS 0.008695f
C830 B.n684 VSUBS 0.008695f
C831 B.n685 VSUBS 0.008695f
C832 B.n686 VSUBS 0.008695f
C833 B.n687 VSUBS 0.008695f
C834 B.n688 VSUBS 0.008695f
C835 B.n689 VSUBS 0.008695f
C836 B.n690 VSUBS 0.008695f
C837 B.n691 VSUBS 0.008695f
C838 B.n692 VSUBS 0.008695f
C839 B.n693 VSUBS 0.008695f
C840 B.n694 VSUBS 0.008695f
C841 B.n695 VSUBS 0.008695f
C842 B.n696 VSUBS 0.008695f
C843 B.n697 VSUBS 0.008695f
C844 B.n698 VSUBS 0.008695f
C845 B.n699 VSUBS 0.008695f
C846 B.n700 VSUBS 0.008695f
C847 B.n701 VSUBS 0.008695f
C848 B.n702 VSUBS 0.008695f
C849 B.n703 VSUBS 0.008695f
C850 B.n704 VSUBS 0.008695f
C851 B.n705 VSUBS 0.008695f
C852 B.n706 VSUBS 0.008695f
C853 B.n707 VSUBS 0.008695f
C854 B.n708 VSUBS 0.008695f
C855 B.n709 VSUBS 0.008695f
C856 B.n710 VSUBS 0.008695f
C857 B.n711 VSUBS 0.008695f
C858 B.n712 VSUBS 0.008695f
C859 B.n713 VSUBS 0.008695f
C860 B.n714 VSUBS 0.008695f
C861 B.n715 VSUBS 0.008695f
C862 B.n716 VSUBS 0.008695f
C863 B.n717 VSUBS 0.008695f
C864 B.n718 VSUBS 0.008695f
C865 B.n719 VSUBS 0.008695f
C866 B.n720 VSUBS 0.008695f
C867 B.n721 VSUBS 0.008695f
C868 B.n722 VSUBS 0.008695f
C869 B.n723 VSUBS 0.008695f
C870 B.n724 VSUBS 0.008695f
C871 B.n725 VSUBS 0.008695f
C872 B.n726 VSUBS 0.008695f
C873 B.n727 VSUBS 0.008695f
C874 B.n728 VSUBS 0.008695f
C875 B.n729 VSUBS 0.008695f
C876 B.n730 VSUBS 0.008695f
C877 B.n731 VSUBS 0.008695f
C878 B.n732 VSUBS 0.008695f
C879 B.n733 VSUBS 0.008695f
C880 B.n734 VSUBS 0.008695f
C881 B.n735 VSUBS 0.008695f
C882 B.n736 VSUBS 0.008695f
C883 B.n737 VSUBS 0.008695f
C884 B.n738 VSUBS 0.008695f
C885 B.n739 VSUBS 0.008695f
C886 B.n740 VSUBS 0.008695f
C887 B.n741 VSUBS 0.008695f
C888 B.n742 VSUBS 0.008695f
C889 B.n743 VSUBS 0.008695f
C890 B.n744 VSUBS 0.008695f
C891 B.n745 VSUBS 0.006009f
C892 B.n746 VSUBS 0.020144f
C893 B.n747 VSUBS 0.007032f
C894 B.n748 VSUBS 0.008695f
C895 B.n749 VSUBS 0.008695f
C896 B.n750 VSUBS 0.008695f
C897 B.n751 VSUBS 0.008695f
C898 B.n752 VSUBS 0.008695f
C899 B.n753 VSUBS 0.008695f
C900 B.n754 VSUBS 0.008695f
C901 B.n755 VSUBS 0.008695f
C902 B.n756 VSUBS 0.008695f
C903 B.n757 VSUBS 0.008695f
C904 B.n758 VSUBS 0.008695f
C905 B.n759 VSUBS 0.007032f
C906 B.n760 VSUBS 0.008695f
C907 B.n761 VSUBS 0.008695f
C908 B.n762 VSUBS 0.008695f
C909 B.n763 VSUBS 0.008695f
C910 B.n764 VSUBS 0.008695f
C911 B.n765 VSUBS 0.008695f
C912 B.n766 VSUBS 0.008695f
C913 B.n767 VSUBS 0.008695f
C914 B.n768 VSUBS 0.008695f
C915 B.n769 VSUBS 0.008695f
C916 B.n770 VSUBS 0.008695f
C917 B.n771 VSUBS 0.008695f
C918 B.n772 VSUBS 0.008695f
C919 B.n773 VSUBS 0.008695f
C920 B.n774 VSUBS 0.008695f
C921 B.n775 VSUBS 0.008695f
C922 B.n776 VSUBS 0.008695f
C923 B.n777 VSUBS 0.008695f
C924 B.n778 VSUBS 0.008695f
C925 B.n779 VSUBS 0.008695f
C926 B.n780 VSUBS 0.008695f
C927 B.n781 VSUBS 0.008695f
C928 B.n782 VSUBS 0.008695f
C929 B.n783 VSUBS 0.008695f
C930 B.n784 VSUBS 0.008695f
C931 B.n785 VSUBS 0.008695f
C932 B.n786 VSUBS 0.008695f
C933 B.n787 VSUBS 0.008695f
C934 B.n788 VSUBS 0.008695f
C935 B.n789 VSUBS 0.008695f
C936 B.n790 VSUBS 0.008695f
C937 B.n791 VSUBS 0.008695f
C938 B.n792 VSUBS 0.008695f
C939 B.n793 VSUBS 0.008695f
C940 B.n794 VSUBS 0.008695f
C941 B.n795 VSUBS 0.008695f
C942 B.n796 VSUBS 0.008695f
C943 B.n797 VSUBS 0.008695f
C944 B.n798 VSUBS 0.008695f
C945 B.n799 VSUBS 0.008695f
C946 B.n800 VSUBS 0.008695f
C947 B.n801 VSUBS 0.008695f
C948 B.n802 VSUBS 0.008695f
C949 B.n803 VSUBS 0.008695f
C950 B.n804 VSUBS 0.008695f
C951 B.n805 VSUBS 0.008695f
C952 B.n806 VSUBS 0.008695f
C953 B.n807 VSUBS 0.008695f
C954 B.n808 VSUBS 0.008695f
C955 B.n809 VSUBS 0.008695f
C956 B.n810 VSUBS 0.008695f
C957 B.n811 VSUBS 0.008695f
C958 B.n812 VSUBS 0.008695f
C959 B.n813 VSUBS 0.008695f
C960 B.n814 VSUBS 0.008695f
C961 B.n815 VSUBS 0.008695f
C962 B.n816 VSUBS 0.008695f
C963 B.n817 VSUBS 0.008695f
C964 B.n818 VSUBS 0.008695f
C965 B.n819 VSUBS 0.008695f
C966 B.n820 VSUBS 0.008695f
C967 B.n821 VSUBS 0.008695f
C968 B.n822 VSUBS 0.008695f
C969 B.n823 VSUBS 0.008695f
C970 B.n824 VSUBS 0.008695f
C971 B.n825 VSUBS 0.008695f
C972 B.n826 VSUBS 0.008695f
C973 B.n827 VSUBS 0.008695f
C974 B.n828 VSUBS 0.008695f
C975 B.n829 VSUBS 0.008695f
C976 B.n830 VSUBS 0.008695f
C977 B.n831 VSUBS 0.008695f
C978 B.n832 VSUBS 0.008695f
C979 B.n833 VSUBS 0.008695f
C980 B.n834 VSUBS 0.008695f
C981 B.n835 VSUBS 0.008695f
C982 B.n836 VSUBS 0.020657f
C983 B.n837 VSUBS 0.019236f
C984 B.n838 VSUBS 0.019236f
C985 B.n839 VSUBS 0.008695f
C986 B.n840 VSUBS 0.008695f
C987 B.n841 VSUBS 0.008695f
C988 B.n842 VSUBS 0.008695f
C989 B.n843 VSUBS 0.008695f
C990 B.n844 VSUBS 0.008695f
C991 B.n845 VSUBS 0.008695f
C992 B.n846 VSUBS 0.008695f
C993 B.n847 VSUBS 0.008695f
C994 B.n848 VSUBS 0.008695f
C995 B.n849 VSUBS 0.008695f
C996 B.n850 VSUBS 0.008695f
C997 B.n851 VSUBS 0.008695f
C998 B.n852 VSUBS 0.008695f
C999 B.n853 VSUBS 0.008695f
C1000 B.n854 VSUBS 0.008695f
C1001 B.n855 VSUBS 0.008695f
C1002 B.n856 VSUBS 0.008695f
C1003 B.n857 VSUBS 0.008695f
C1004 B.n858 VSUBS 0.008695f
C1005 B.n859 VSUBS 0.008695f
C1006 B.n860 VSUBS 0.008695f
C1007 B.n861 VSUBS 0.008695f
C1008 B.n862 VSUBS 0.008695f
C1009 B.n863 VSUBS 0.008695f
C1010 B.n864 VSUBS 0.008695f
C1011 B.n865 VSUBS 0.008695f
C1012 B.n866 VSUBS 0.008695f
C1013 B.n867 VSUBS 0.008695f
C1014 B.n868 VSUBS 0.008695f
C1015 B.n869 VSUBS 0.008695f
C1016 B.n870 VSUBS 0.008695f
C1017 B.n871 VSUBS 0.008695f
C1018 B.n872 VSUBS 0.008695f
C1019 B.n873 VSUBS 0.008695f
C1020 B.n874 VSUBS 0.008695f
C1021 B.n875 VSUBS 0.008695f
C1022 B.n876 VSUBS 0.008695f
C1023 B.n877 VSUBS 0.008695f
C1024 B.n878 VSUBS 0.008695f
C1025 B.n879 VSUBS 0.008695f
C1026 B.n880 VSUBS 0.008695f
C1027 B.n881 VSUBS 0.008695f
C1028 B.n882 VSUBS 0.008695f
C1029 B.n883 VSUBS 0.008695f
C1030 B.n884 VSUBS 0.008695f
C1031 B.n885 VSUBS 0.008695f
C1032 B.n886 VSUBS 0.008695f
C1033 B.n887 VSUBS 0.008695f
C1034 B.n888 VSUBS 0.008695f
C1035 B.n889 VSUBS 0.008695f
C1036 B.n890 VSUBS 0.008695f
C1037 B.n891 VSUBS 0.008695f
C1038 B.n892 VSUBS 0.008695f
C1039 B.n893 VSUBS 0.008695f
C1040 B.n894 VSUBS 0.008695f
C1041 B.n895 VSUBS 0.008695f
C1042 B.n896 VSUBS 0.008695f
C1043 B.n897 VSUBS 0.008695f
C1044 B.n898 VSUBS 0.008695f
C1045 B.n899 VSUBS 0.008695f
C1046 B.n900 VSUBS 0.008695f
C1047 B.n901 VSUBS 0.008695f
C1048 B.n902 VSUBS 0.008695f
C1049 B.n903 VSUBS 0.008695f
C1050 B.n904 VSUBS 0.008695f
C1051 B.n905 VSUBS 0.008695f
C1052 B.n906 VSUBS 0.008695f
C1053 B.n907 VSUBS 0.008695f
C1054 B.n908 VSUBS 0.008695f
C1055 B.n909 VSUBS 0.008695f
C1056 B.n910 VSUBS 0.008695f
C1057 B.n911 VSUBS 0.008695f
C1058 B.n912 VSUBS 0.008695f
C1059 B.n913 VSUBS 0.008695f
C1060 B.n914 VSUBS 0.008695f
C1061 B.n915 VSUBS 0.008695f
C1062 B.n916 VSUBS 0.008695f
C1063 B.n917 VSUBS 0.008695f
C1064 B.n918 VSUBS 0.008695f
C1065 B.n919 VSUBS 0.008695f
C1066 B.n920 VSUBS 0.008695f
C1067 B.n921 VSUBS 0.008695f
C1068 B.n922 VSUBS 0.008695f
C1069 B.n923 VSUBS 0.011346f
C1070 B.n924 VSUBS 0.012086f
C1071 B.n925 VSUBS 0.024035f
C1072 VDD1.t0 VSUBS 3.66992f
C1073 VDD1.t8 VSUBS 0.34469f
C1074 VDD1.t7 VSUBS 0.34469f
C1075 VDD1.n0 VSUBS 2.80072f
C1076 VDD1.n1 VSUBS 1.71211f
C1077 VDD1.t9 VSUBS 3.66991f
C1078 VDD1.t1 VSUBS 0.34469f
C1079 VDD1.t4 VSUBS 0.34469f
C1080 VDD1.n2 VSUBS 2.80072f
C1081 VDD1.n3 VSUBS 1.70271f
C1082 VDD1.t6 VSUBS 0.34469f
C1083 VDD1.t2 VSUBS 0.34469f
C1084 VDD1.n4 VSUBS 2.82436f
C1085 VDD1.n5 VSUBS 4.00127f
C1086 VDD1.t5 VSUBS 0.34469f
C1087 VDD1.t3 VSUBS 0.34469f
C1088 VDD1.n6 VSUBS 2.80071f
C1089 VDD1.n7 VSUBS 4.22964f
C1090 VTAIL.t3 VSUBS 0.332447f
C1091 VTAIL.t2 VSUBS 0.332447f
C1092 VTAIL.n0 VSUBS 2.53998f
C1093 VTAIL.n1 VSUBS 0.981819f
C1094 VTAIL.t9 VSUBS 3.32808f
C1095 VTAIL.n2 VSUBS 1.1507f
C1096 VTAIL.t17 VSUBS 0.332447f
C1097 VTAIL.t15 VSUBS 0.332447f
C1098 VTAIL.n3 VSUBS 2.53998f
C1099 VTAIL.n4 VSUBS 1.10089f
C1100 VTAIL.t12 VSUBS 0.332447f
C1101 VTAIL.t10 VSUBS 0.332447f
C1102 VTAIL.n5 VSUBS 2.53998f
C1103 VTAIL.n6 VSUBS 2.87168f
C1104 VTAIL.t6 VSUBS 0.332447f
C1105 VTAIL.t18 VSUBS 0.332447f
C1106 VTAIL.n7 VSUBS 2.53999f
C1107 VTAIL.n8 VSUBS 2.87167f
C1108 VTAIL.t0 VSUBS 0.332447f
C1109 VTAIL.t7 VSUBS 0.332447f
C1110 VTAIL.n9 VSUBS 2.53999f
C1111 VTAIL.n10 VSUBS 1.10089f
C1112 VTAIL.t4 VSUBS 3.32809f
C1113 VTAIL.n11 VSUBS 1.1507f
C1114 VTAIL.t11 VSUBS 0.332447f
C1115 VTAIL.t13 VSUBS 0.332447f
C1116 VTAIL.n12 VSUBS 2.53999f
C1117 VTAIL.n13 VSUBS 1.03212f
C1118 VTAIL.t14 VSUBS 0.332447f
C1119 VTAIL.t16 VSUBS 0.332447f
C1120 VTAIL.n14 VSUBS 2.53999f
C1121 VTAIL.n15 VSUBS 1.10089f
C1122 VTAIL.t8 VSUBS 3.32808f
C1123 VTAIL.n16 VSUBS 2.76803f
C1124 VTAIL.t5 VSUBS 3.32808f
C1125 VTAIL.n17 VSUBS 2.76803f
C1126 VTAIL.t19 VSUBS 0.332447f
C1127 VTAIL.t1 VSUBS 0.332447f
C1128 VTAIL.n18 VSUBS 2.53998f
C1129 VTAIL.n19 VSUBS 0.928983f
C1130 VP.n0 VSUBS 0.038214f
C1131 VP.t7 VSUBS 3.02255f
C1132 VP.n1 VSUBS 0.038929f
C1133 VP.n2 VSUBS 0.028987f
C1134 VP.t3 VSUBS 3.02255f
C1135 VP.n3 VSUBS 1.05689f
C1136 VP.n4 VSUBS 0.028987f
C1137 VP.n5 VSUBS 0.054519f
C1138 VP.n6 VSUBS 0.028987f
C1139 VP.t5 VSUBS 3.02255f
C1140 VP.n7 VSUBS 0.054519f
C1141 VP.n8 VSUBS 0.028987f
C1142 VP.t8 VSUBS 3.02255f
C1143 VP.n9 VSUBS 1.05689f
C1144 VP.n10 VSUBS 0.028987f
C1145 VP.n11 VSUBS 0.038929f
C1146 VP.n12 VSUBS 0.038214f
C1147 VP.t0 VSUBS 3.02255f
C1148 VP.n13 VSUBS 0.038214f
C1149 VP.t6 VSUBS 3.02255f
C1150 VP.n14 VSUBS 0.038929f
C1151 VP.n15 VSUBS 0.028987f
C1152 VP.t4 VSUBS 3.02255f
C1153 VP.n16 VSUBS 1.05689f
C1154 VP.n17 VSUBS 0.028987f
C1155 VP.n18 VSUBS 0.054519f
C1156 VP.n19 VSUBS 0.028987f
C1157 VP.t2 VSUBS 3.02255f
C1158 VP.n20 VSUBS 0.054519f
C1159 VP.n21 VSUBS 0.028987f
C1160 VP.t1 VSUBS 3.02255f
C1161 VP.n22 VSUBS 1.14495f
C1162 VP.t9 VSUBS 3.25845f
C1163 VP.n23 VSUBS 1.1102f
C1164 VP.n24 VSUBS 0.278111f
C1165 VP.n25 VSUBS 0.046323f
C1166 VP.n26 VSUBS 0.058234f
C1167 VP.n27 VSUBS 0.025274f
C1168 VP.n28 VSUBS 0.028987f
C1169 VP.n29 VSUBS 0.028987f
C1170 VP.n30 VSUBS 0.028987f
C1171 VP.n31 VSUBS 0.053753f
C1172 VP.n32 VSUBS 1.08411f
C1173 VP.n33 VSUBS 0.053753f
C1174 VP.n34 VSUBS 0.028987f
C1175 VP.n35 VSUBS 0.028987f
C1176 VP.n36 VSUBS 0.028987f
C1177 VP.n37 VSUBS 0.025274f
C1178 VP.n38 VSUBS 0.058234f
C1179 VP.n39 VSUBS 0.046323f
C1180 VP.n40 VSUBS 0.028987f
C1181 VP.n41 VSUBS 0.028987f
C1182 VP.n42 VSUBS 0.034647f
C1183 VP.n43 VSUBS 0.053753f
C1184 VP.n44 VSUBS 0.045345f
C1185 VP.n45 VSUBS 0.028987f
C1186 VP.n46 VSUBS 0.028987f
C1187 VP.n47 VSUBS 0.028987f
C1188 VP.n48 VSUBS 0.053753f
C1189 VP.n49 VSUBS 0.038893f
C1190 VP.n50 VSUBS 1.15207f
C1191 VP.n51 VSUBS 1.85098f
C1192 VP.n52 VSUBS 1.86996f
C1193 VP.n53 VSUBS 1.15207f
C1194 VP.n54 VSUBS 0.038893f
C1195 VP.n55 VSUBS 0.053753f
C1196 VP.n56 VSUBS 0.028987f
C1197 VP.n57 VSUBS 0.028987f
C1198 VP.n58 VSUBS 0.028987f
C1199 VP.n59 VSUBS 0.045345f
C1200 VP.n60 VSUBS 0.053753f
C1201 VP.n61 VSUBS 0.034647f
C1202 VP.n62 VSUBS 0.028987f
C1203 VP.n63 VSUBS 0.028987f
C1204 VP.n64 VSUBS 0.046323f
C1205 VP.n65 VSUBS 0.058234f
C1206 VP.n66 VSUBS 0.025274f
C1207 VP.n67 VSUBS 0.028987f
C1208 VP.n68 VSUBS 0.028987f
C1209 VP.n69 VSUBS 0.028987f
C1210 VP.n70 VSUBS 0.053753f
C1211 VP.n71 VSUBS 1.08411f
C1212 VP.n72 VSUBS 0.053753f
C1213 VP.n73 VSUBS 0.028987f
C1214 VP.n74 VSUBS 0.028987f
C1215 VP.n75 VSUBS 0.028987f
C1216 VP.n76 VSUBS 0.025274f
C1217 VP.n77 VSUBS 0.058234f
C1218 VP.n78 VSUBS 0.046323f
C1219 VP.n79 VSUBS 0.028987f
C1220 VP.n80 VSUBS 0.028987f
C1221 VP.n81 VSUBS 0.034647f
C1222 VP.n82 VSUBS 0.053753f
C1223 VP.n83 VSUBS 0.045345f
C1224 VP.n84 VSUBS 0.028987f
C1225 VP.n85 VSUBS 0.028987f
C1226 VP.n86 VSUBS 0.028987f
C1227 VP.n87 VSUBS 0.053753f
C1228 VP.n88 VSUBS 0.038893f
C1229 VP.n89 VSUBS 1.15207f
C1230 VP.n90 VSUBS 0.045933f
.ends

