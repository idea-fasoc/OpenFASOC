* NGSPICE file created from diff_pair_sample_1440.ext - technology: sky130A

.subckt diff_pair_sample_1440 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=0 ps=0 w=16.05 l=3.91
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=6.2595 ps=32.88 w=16.05 l=3.91
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=0 ps=0 w=16.05 l=3.91
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=0 ps=0 w=16.05 l=3.91
X4 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=6.2595 ps=32.88 w=16.05 l=3.91
X5 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=6.2595 ps=32.88 w=16.05 l=3.91
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=0 ps=0 w=16.05 l=3.91
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2595 pd=32.88 as=6.2595 ps=32.88 w=16.05 l=3.91
R0 B.n863 B.n862 585
R1 B.n864 B.n863 585
R2 B.n358 B.n121 585
R3 B.n357 B.n356 585
R4 B.n355 B.n354 585
R5 B.n353 B.n352 585
R6 B.n351 B.n350 585
R7 B.n349 B.n348 585
R8 B.n347 B.n346 585
R9 B.n345 B.n344 585
R10 B.n343 B.n342 585
R11 B.n341 B.n340 585
R12 B.n339 B.n338 585
R13 B.n337 B.n336 585
R14 B.n335 B.n334 585
R15 B.n333 B.n332 585
R16 B.n331 B.n330 585
R17 B.n329 B.n328 585
R18 B.n327 B.n326 585
R19 B.n325 B.n324 585
R20 B.n323 B.n322 585
R21 B.n321 B.n320 585
R22 B.n319 B.n318 585
R23 B.n317 B.n316 585
R24 B.n315 B.n314 585
R25 B.n313 B.n312 585
R26 B.n311 B.n310 585
R27 B.n309 B.n308 585
R28 B.n307 B.n306 585
R29 B.n305 B.n304 585
R30 B.n303 B.n302 585
R31 B.n301 B.n300 585
R32 B.n299 B.n298 585
R33 B.n297 B.n296 585
R34 B.n295 B.n294 585
R35 B.n293 B.n292 585
R36 B.n291 B.n290 585
R37 B.n289 B.n288 585
R38 B.n287 B.n286 585
R39 B.n285 B.n284 585
R40 B.n283 B.n282 585
R41 B.n281 B.n280 585
R42 B.n279 B.n278 585
R43 B.n277 B.n276 585
R44 B.n275 B.n274 585
R45 B.n273 B.n272 585
R46 B.n271 B.n270 585
R47 B.n269 B.n268 585
R48 B.n267 B.n266 585
R49 B.n265 B.n264 585
R50 B.n263 B.n262 585
R51 B.n261 B.n260 585
R52 B.n259 B.n258 585
R53 B.n257 B.n256 585
R54 B.n255 B.n254 585
R55 B.n252 B.n251 585
R56 B.n250 B.n249 585
R57 B.n248 B.n247 585
R58 B.n246 B.n245 585
R59 B.n244 B.n243 585
R60 B.n242 B.n241 585
R61 B.n240 B.n239 585
R62 B.n238 B.n237 585
R63 B.n236 B.n235 585
R64 B.n234 B.n233 585
R65 B.n232 B.n231 585
R66 B.n230 B.n229 585
R67 B.n228 B.n227 585
R68 B.n226 B.n225 585
R69 B.n224 B.n223 585
R70 B.n222 B.n221 585
R71 B.n220 B.n219 585
R72 B.n218 B.n217 585
R73 B.n216 B.n215 585
R74 B.n214 B.n213 585
R75 B.n212 B.n211 585
R76 B.n210 B.n209 585
R77 B.n208 B.n207 585
R78 B.n206 B.n205 585
R79 B.n204 B.n203 585
R80 B.n202 B.n201 585
R81 B.n200 B.n199 585
R82 B.n198 B.n197 585
R83 B.n196 B.n195 585
R84 B.n194 B.n193 585
R85 B.n192 B.n191 585
R86 B.n190 B.n189 585
R87 B.n188 B.n187 585
R88 B.n186 B.n185 585
R89 B.n184 B.n183 585
R90 B.n182 B.n181 585
R91 B.n180 B.n179 585
R92 B.n178 B.n177 585
R93 B.n176 B.n175 585
R94 B.n174 B.n173 585
R95 B.n172 B.n171 585
R96 B.n170 B.n169 585
R97 B.n168 B.n167 585
R98 B.n166 B.n165 585
R99 B.n164 B.n163 585
R100 B.n162 B.n161 585
R101 B.n160 B.n159 585
R102 B.n158 B.n157 585
R103 B.n156 B.n155 585
R104 B.n154 B.n153 585
R105 B.n152 B.n151 585
R106 B.n150 B.n149 585
R107 B.n148 B.n147 585
R108 B.n146 B.n145 585
R109 B.n144 B.n143 585
R110 B.n142 B.n141 585
R111 B.n140 B.n139 585
R112 B.n138 B.n137 585
R113 B.n136 B.n135 585
R114 B.n134 B.n133 585
R115 B.n132 B.n131 585
R116 B.n130 B.n129 585
R117 B.n128 B.n127 585
R118 B.n861 B.n62 585
R119 B.n865 B.n62 585
R120 B.n860 B.n61 585
R121 B.n866 B.n61 585
R122 B.n859 B.n858 585
R123 B.n858 B.n57 585
R124 B.n857 B.n56 585
R125 B.n872 B.n56 585
R126 B.n856 B.n55 585
R127 B.n873 B.n55 585
R128 B.n855 B.n54 585
R129 B.n874 B.n54 585
R130 B.n854 B.n853 585
R131 B.n853 B.n50 585
R132 B.n852 B.n49 585
R133 B.n880 B.n49 585
R134 B.n851 B.n48 585
R135 B.n881 B.n48 585
R136 B.n850 B.n47 585
R137 B.n882 B.n47 585
R138 B.n849 B.n848 585
R139 B.n848 B.n43 585
R140 B.n847 B.n42 585
R141 B.n888 B.n42 585
R142 B.n846 B.n41 585
R143 B.n889 B.n41 585
R144 B.n845 B.n40 585
R145 B.n890 B.n40 585
R146 B.n844 B.n843 585
R147 B.n843 B.n36 585
R148 B.n842 B.n35 585
R149 B.n896 B.n35 585
R150 B.n841 B.n34 585
R151 B.n897 B.n34 585
R152 B.n840 B.n33 585
R153 B.n898 B.n33 585
R154 B.n839 B.n838 585
R155 B.n838 B.n29 585
R156 B.n837 B.n28 585
R157 B.n904 B.n28 585
R158 B.n836 B.n27 585
R159 B.n905 B.n27 585
R160 B.n835 B.n26 585
R161 B.n906 B.n26 585
R162 B.n834 B.n833 585
R163 B.n833 B.n22 585
R164 B.n832 B.n21 585
R165 B.n912 B.n21 585
R166 B.n831 B.n20 585
R167 B.n913 B.n20 585
R168 B.n830 B.n19 585
R169 B.n914 B.n19 585
R170 B.n829 B.n828 585
R171 B.n828 B.n15 585
R172 B.n827 B.n14 585
R173 B.n920 B.n14 585
R174 B.n826 B.n13 585
R175 B.n921 B.n13 585
R176 B.n825 B.n12 585
R177 B.n922 B.n12 585
R178 B.n824 B.n823 585
R179 B.n823 B.n8 585
R180 B.n822 B.n7 585
R181 B.n928 B.n7 585
R182 B.n821 B.n6 585
R183 B.n929 B.n6 585
R184 B.n820 B.n5 585
R185 B.n930 B.n5 585
R186 B.n819 B.n818 585
R187 B.n818 B.n4 585
R188 B.n817 B.n359 585
R189 B.n817 B.n816 585
R190 B.n807 B.n360 585
R191 B.n361 B.n360 585
R192 B.n809 B.n808 585
R193 B.n810 B.n809 585
R194 B.n806 B.n366 585
R195 B.n366 B.n365 585
R196 B.n805 B.n804 585
R197 B.n804 B.n803 585
R198 B.n368 B.n367 585
R199 B.n369 B.n368 585
R200 B.n796 B.n795 585
R201 B.n797 B.n796 585
R202 B.n794 B.n374 585
R203 B.n374 B.n373 585
R204 B.n793 B.n792 585
R205 B.n792 B.n791 585
R206 B.n376 B.n375 585
R207 B.n377 B.n376 585
R208 B.n784 B.n783 585
R209 B.n785 B.n784 585
R210 B.n782 B.n382 585
R211 B.n382 B.n381 585
R212 B.n781 B.n780 585
R213 B.n780 B.n779 585
R214 B.n384 B.n383 585
R215 B.n385 B.n384 585
R216 B.n772 B.n771 585
R217 B.n773 B.n772 585
R218 B.n770 B.n390 585
R219 B.n390 B.n389 585
R220 B.n769 B.n768 585
R221 B.n768 B.n767 585
R222 B.n392 B.n391 585
R223 B.n393 B.n392 585
R224 B.n760 B.n759 585
R225 B.n761 B.n760 585
R226 B.n758 B.n398 585
R227 B.n398 B.n397 585
R228 B.n757 B.n756 585
R229 B.n756 B.n755 585
R230 B.n400 B.n399 585
R231 B.n401 B.n400 585
R232 B.n748 B.n747 585
R233 B.n749 B.n748 585
R234 B.n746 B.n406 585
R235 B.n406 B.n405 585
R236 B.n745 B.n744 585
R237 B.n744 B.n743 585
R238 B.n408 B.n407 585
R239 B.n409 B.n408 585
R240 B.n736 B.n735 585
R241 B.n737 B.n736 585
R242 B.n734 B.n414 585
R243 B.n414 B.n413 585
R244 B.n733 B.n732 585
R245 B.n732 B.n731 585
R246 B.n416 B.n415 585
R247 B.n417 B.n416 585
R248 B.n724 B.n723 585
R249 B.n725 B.n724 585
R250 B.n722 B.n422 585
R251 B.n422 B.n421 585
R252 B.n716 B.n715 585
R253 B.n714 B.n482 585
R254 B.n713 B.n481 585
R255 B.n718 B.n481 585
R256 B.n712 B.n711 585
R257 B.n710 B.n709 585
R258 B.n708 B.n707 585
R259 B.n706 B.n705 585
R260 B.n704 B.n703 585
R261 B.n702 B.n701 585
R262 B.n700 B.n699 585
R263 B.n698 B.n697 585
R264 B.n696 B.n695 585
R265 B.n694 B.n693 585
R266 B.n692 B.n691 585
R267 B.n690 B.n689 585
R268 B.n688 B.n687 585
R269 B.n686 B.n685 585
R270 B.n684 B.n683 585
R271 B.n682 B.n681 585
R272 B.n680 B.n679 585
R273 B.n678 B.n677 585
R274 B.n676 B.n675 585
R275 B.n674 B.n673 585
R276 B.n672 B.n671 585
R277 B.n670 B.n669 585
R278 B.n668 B.n667 585
R279 B.n666 B.n665 585
R280 B.n664 B.n663 585
R281 B.n662 B.n661 585
R282 B.n660 B.n659 585
R283 B.n658 B.n657 585
R284 B.n656 B.n655 585
R285 B.n654 B.n653 585
R286 B.n652 B.n651 585
R287 B.n650 B.n649 585
R288 B.n648 B.n647 585
R289 B.n646 B.n645 585
R290 B.n644 B.n643 585
R291 B.n642 B.n641 585
R292 B.n640 B.n639 585
R293 B.n638 B.n637 585
R294 B.n636 B.n635 585
R295 B.n634 B.n633 585
R296 B.n632 B.n631 585
R297 B.n630 B.n629 585
R298 B.n628 B.n627 585
R299 B.n626 B.n625 585
R300 B.n624 B.n623 585
R301 B.n622 B.n621 585
R302 B.n620 B.n619 585
R303 B.n618 B.n617 585
R304 B.n616 B.n615 585
R305 B.n614 B.n613 585
R306 B.n612 B.n611 585
R307 B.n609 B.n608 585
R308 B.n607 B.n606 585
R309 B.n605 B.n604 585
R310 B.n603 B.n602 585
R311 B.n601 B.n600 585
R312 B.n599 B.n598 585
R313 B.n597 B.n596 585
R314 B.n595 B.n594 585
R315 B.n593 B.n592 585
R316 B.n591 B.n590 585
R317 B.n589 B.n588 585
R318 B.n587 B.n586 585
R319 B.n585 B.n584 585
R320 B.n583 B.n582 585
R321 B.n581 B.n580 585
R322 B.n579 B.n578 585
R323 B.n577 B.n576 585
R324 B.n575 B.n574 585
R325 B.n573 B.n572 585
R326 B.n571 B.n570 585
R327 B.n569 B.n568 585
R328 B.n567 B.n566 585
R329 B.n565 B.n564 585
R330 B.n563 B.n562 585
R331 B.n561 B.n560 585
R332 B.n559 B.n558 585
R333 B.n557 B.n556 585
R334 B.n555 B.n554 585
R335 B.n553 B.n552 585
R336 B.n551 B.n550 585
R337 B.n549 B.n548 585
R338 B.n547 B.n546 585
R339 B.n545 B.n544 585
R340 B.n543 B.n542 585
R341 B.n541 B.n540 585
R342 B.n539 B.n538 585
R343 B.n537 B.n536 585
R344 B.n535 B.n534 585
R345 B.n533 B.n532 585
R346 B.n531 B.n530 585
R347 B.n529 B.n528 585
R348 B.n527 B.n526 585
R349 B.n525 B.n524 585
R350 B.n523 B.n522 585
R351 B.n521 B.n520 585
R352 B.n519 B.n518 585
R353 B.n517 B.n516 585
R354 B.n515 B.n514 585
R355 B.n513 B.n512 585
R356 B.n511 B.n510 585
R357 B.n509 B.n508 585
R358 B.n507 B.n506 585
R359 B.n505 B.n504 585
R360 B.n503 B.n502 585
R361 B.n501 B.n500 585
R362 B.n499 B.n498 585
R363 B.n497 B.n496 585
R364 B.n495 B.n494 585
R365 B.n493 B.n492 585
R366 B.n491 B.n490 585
R367 B.n489 B.n488 585
R368 B.n424 B.n423 585
R369 B.n721 B.n720 585
R370 B.n420 B.n419 585
R371 B.n421 B.n420 585
R372 B.n727 B.n726 585
R373 B.n726 B.n725 585
R374 B.n728 B.n418 585
R375 B.n418 B.n417 585
R376 B.n730 B.n729 585
R377 B.n731 B.n730 585
R378 B.n412 B.n411 585
R379 B.n413 B.n412 585
R380 B.n739 B.n738 585
R381 B.n738 B.n737 585
R382 B.n740 B.n410 585
R383 B.n410 B.n409 585
R384 B.n742 B.n741 585
R385 B.n743 B.n742 585
R386 B.n404 B.n403 585
R387 B.n405 B.n404 585
R388 B.n751 B.n750 585
R389 B.n750 B.n749 585
R390 B.n752 B.n402 585
R391 B.n402 B.n401 585
R392 B.n754 B.n753 585
R393 B.n755 B.n754 585
R394 B.n396 B.n395 585
R395 B.n397 B.n396 585
R396 B.n763 B.n762 585
R397 B.n762 B.n761 585
R398 B.n764 B.n394 585
R399 B.n394 B.n393 585
R400 B.n766 B.n765 585
R401 B.n767 B.n766 585
R402 B.n388 B.n387 585
R403 B.n389 B.n388 585
R404 B.n775 B.n774 585
R405 B.n774 B.n773 585
R406 B.n776 B.n386 585
R407 B.n386 B.n385 585
R408 B.n778 B.n777 585
R409 B.n779 B.n778 585
R410 B.n380 B.n379 585
R411 B.n381 B.n380 585
R412 B.n787 B.n786 585
R413 B.n786 B.n785 585
R414 B.n788 B.n378 585
R415 B.n378 B.n377 585
R416 B.n790 B.n789 585
R417 B.n791 B.n790 585
R418 B.n372 B.n371 585
R419 B.n373 B.n372 585
R420 B.n799 B.n798 585
R421 B.n798 B.n797 585
R422 B.n800 B.n370 585
R423 B.n370 B.n369 585
R424 B.n802 B.n801 585
R425 B.n803 B.n802 585
R426 B.n364 B.n363 585
R427 B.n365 B.n364 585
R428 B.n812 B.n811 585
R429 B.n811 B.n810 585
R430 B.n813 B.n362 585
R431 B.n362 B.n361 585
R432 B.n815 B.n814 585
R433 B.n816 B.n815 585
R434 B.n2 B.n0 585
R435 B.n4 B.n2 585
R436 B.n3 B.n1 585
R437 B.n929 B.n3 585
R438 B.n927 B.n926 585
R439 B.n928 B.n927 585
R440 B.n925 B.n9 585
R441 B.n9 B.n8 585
R442 B.n924 B.n923 585
R443 B.n923 B.n922 585
R444 B.n11 B.n10 585
R445 B.n921 B.n11 585
R446 B.n919 B.n918 585
R447 B.n920 B.n919 585
R448 B.n917 B.n16 585
R449 B.n16 B.n15 585
R450 B.n916 B.n915 585
R451 B.n915 B.n914 585
R452 B.n18 B.n17 585
R453 B.n913 B.n18 585
R454 B.n911 B.n910 585
R455 B.n912 B.n911 585
R456 B.n909 B.n23 585
R457 B.n23 B.n22 585
R458 B.n908 B.n907 585
R459 B.n907 B.n906 585
R460 B.n25 B.n24 585
R461 B.n905 B.n25 585
R462 B.n903 B.n902 585
R463 B.n904 B.n903 585
R464 B.n901 B.n30 585
R465 B.n30 B.n29 585
R466 B.n900 B.n899 585
R467 B.n899 B.n898 585
R468 B.n32 B.n31 585
R469 B.n897 B.n32 585
R470 B.n895 B.n894 585
R471 B.n896 B.n895 585
R472 B.n893 B.n37 585
R473 B.n37 B.n36 585
R474 B.n892 B.n891 585
R475 B.n891 B.n890 585
R476 B.n39 B.n38 585
R477 B.n889 B.n39 585
R478 B.n887 B.n886 585
R479 B.n888 B.n887 585
R480 B.n885 B.n44 585
R481 B.n44 B.n43 585
R482 B.n884 B.n883 585
R483 B.n883 B.n882 585
R484 B.n46 B.n45 585
R485 B.n881 B.n46 585
R486 B.n879 B.n878 585
R487 B.n880 B.n879 585
R488 B.n877 B.n51 585
R489 B.n51 B.n50 585
R490 B.n876 B.n875 585
R491 B.n875 B.n874 585
R492 B.n53 B.n52 585
R493 B.n873 B.n53 585
R494 B.n871 B.n870 585
R495 B.n872 B.n871 585
R496 B.n869 B.n58 585
R497 B.n58 B.n57 585
R498 B.n868 B.n867 585
R499 B.n867 B.n866 585
R500 B.n60 B.n59 585
R501 B.n865 B.n60 585
R502 B.n932 B.n931 585
R503 B.n931 B.n930 585
R504 B.n716 B.n420 478.086
R505 B.n127 B.n60 478.086
R506 B.n720 B.n422 478.086
R507 B.n863 B.n62 478.086
R508 B.n485 B.t5 433.932
R509 B.n483 B.t8 433.932
R510 B.n124 B.t11 433.932
R511 B.n122 B.t14 433.932
R512 B.n486 B.t4 351.7
R513 B.n123 B.t15 351.7
R514 B.n484 B.t7 351.7
R515 B.n125 B.t12 351.7
R516 B.n485 B.t2 308.353
R517 B.n483 B.t6 308.353
R518 B.n124 B.t9 308.353
R519 B.n122 B.t13 308.353
R520 B.n864 B.n120 256.663
R521 B.n864 B.n119 256.663
R522 B.n864 B.n118 256.663
R523 B.n864 B.n117 256.663
R524 B.n864 B.n116 256.663
R525 B.n864 B.n115 256.663
R526 B.n864 B.n114 256.663
R527 B.n864 B.n113 256.663
R528 B.n864 B.n112 256.663
R529 B.n864 B.n111 256.663
R530 B.n864 B.n110 256.663
R531 B.n864 B.n109 256.663
R532 B.n864 B.n108 256.663
R533 B.n864 B.n107 256.663
R534 B.n864 B.n106 256.663
R535 B.n864 B.n105 256.663
R536 B.n864 B.n104 256.663
R537 B.n864 B.n103 256.663
R538 B.n864 B.n102 256.663
R539 B.n864 B.n101 256.663
R540 B.n864 B.n100 256.663
R541 B.n864 B.n99 256.663
R542 B.n864 B.n98 256.663
R543 B.n864 B.n97 256.663
R544 B.n864 B.n96 256.663
R545 B.n864 B.n95 256.663
R546 B.n864 B.n94 256.663
R547 B.n864 B.n93 256.663
R548 B.n864 B.n92 256.663
R549 B.n864 B.n91 256.663
R550 B.n864 B.n90 256.663
R551 B.n864 B.n89 256.663
R552 B.n864 B.n88 256.663
R553 B.n864 B.n87 256.663
R554 B.n864 B.n86 256.663
R555 B.n864 B.n85 256.663
R556 B.n864 B.n84 256.663
R557 B.n864 B.n83 256.663
R558 B.n864 B.n82 256.663
R559 B.n864 B.n81 256.663
R560 B.n864 B.n80 256.663
R561 B.n864 B.n79 256.663
R562 B.n864 B.n78 256.663
R563 B.n864 B.n77 256.663
R564 B.n864 B.n76 256.663
R565 B.n864 B.n75 256.663
R566 B.n864 B.n74 256.663
R567 B.n864 B.n73 256.663
R568 B.n864 B.n72 256.663
R569 B.n864 B.n71 256.663
R570 B.n864 B.n70 256.663
R571 B.n864 B.n69 256.663
R572 B.n864 B.n68 256.663
R573 B.n864 B.n67 256.663
R574 B.n864 B.n66 256.663
R575 B.n864 B.n65 256.663
R576 B.n864 B.n64 256.663
R577 B.n864 B.n63 256.663
R578 B.n718 B.n717 256.663
R579 B.n718 B.n425 256.663
R580 B.n718 B.n426 256.663
R581 B.n718 B.n427 256.663
R582 B.n718 B.n428 256.663
R583 B.n718 B.n429 256.663
R584 B.n718 B.n430 256.663
R585 B.n718 B.n431 256.663
R586 B.n718 B.n432 256.663
R587 B.n718 B.n433 256.663
R588 B.n718 B.n434 256.663
R589 B.n718 B.n435 256.663
R590 B.n718 B.n436 256.663
R591 B.n718 B.n437 256.663
R592 B.n718 B.n438 256.663
R593 B.n718 B.n439 256.663
R594 B.n718 B.n440 256.663
R595 B.n718 B.n441 256.663
R596 B.n718 B.n442 256.663
R597 B.n718 B.n443 256.663
R598 B.n718 B.n444 256.663
R599 B.n718 B.n445 256.663
R600 B.n718 B.n446 256.663
R601 B.n718 B.n447 256.663
R602 B.n718 B.n448 256.663
R603 B.n718 B.n449 256.663
R604 B.n718 B.n450 256.663
R605 B.n718 B.n451 256.663
R606 B.n718 B.n452 256.663
R607 B.n718 B.n453 256.663
R608 B.n718 B.n454 256.663
R609 B.n718 B.n455 256.663
R610 B.n718 B.n456 256.663
R611 B.n718 B.n457 256.663
R612 B.n718 B.n458 256.663
R613 B.n718 B.n459 256.663
R614 B.n718 B.n460 256.663
R615 B.n718 B.n461 256.663
R616 B.n718 B.n462 256.663
R617 B.n718 B.n463 256.663
R618 B.n718 B.n464 256.663
R619 B.n718 B.n465 256.663
R620 B.n718 B.n466 256.663
R621 B.n718 B.n467 256.663
R622 B.n718 B.n468 256.663
R623 B.n718 B.n469 256.663
R624 B.n718 B.n470 256.663
R625 B.n718 B.n471 256.663
R626 B.n718 B.n472 256.663
R627 B.n718 B.n473 256.663
R628 B.n718 B.n474 256.663
R629 B.n718 B.n475 256.663
R630 B.n718 B.n476 256.663
R631 B.n718 B.n477 256.663
R632 B.n718 B.n478 256.663
R633 B.n718 B.n479 256.663
R634 B.n718 B.n480 256.663
R635 B.n719 B.n718 256.663
R636 B.n726 B.n420 163.367
R637 B.n726 B.n418 163.367
R638 B.n730 B.n418 163.367
R639 B.n730 B.n412 163.367
R640 B.n738 B.n412 163.367
R641 B.n738 B.n410 163.367
R642 B.n742 B.n410 163.367
R643 B.n742 B.n404 163.367
R644 B.n750 B.n404 163.367
R645 B.n750 B.n402 163.367
R646 B.n754 B.n402 163.367
R647 B.n754 B.n396 163.367
R648 B.n762 B.n396 163.367
R649 B.n762 B.n394 163.367
R650 B.n766 B.n394 163.367
R651 B.n766 B.n388 163.367
R652 B.n774 B.n388 163.367
R653 B.n774 B.n386 163.367
R654 B.n778 B.n386 163.367
R655 B.n778 B.n380 163.367
R656 B.n786 B.n380 163.367
R657 B.n786 B.n378 163.367
R658 B.n790 B.n378 163.367
R659 B.n790 B.n372 163.367
R660 B.n798 B.n372 163.367
R661 B.n798 B.n370 163.367
R662 B.n802 B.n370 163.367
R663 B.n802 B.n364 163.367
R664 B.n811 B.n364 163.367
R665 B.n811 B.n362 163.367
R666 B.n815 B.n362 163.367
R667 B.n815 B.n2 163.367
R668 B.n931 B.n2 163.367
R669 B.n931 B.n3 163.367
R670 B.n927 B.n3 163.367
R671 B.n927 B.n9 163.367
R672 B.n923 B.n9 163.367
R673 B.n923 B.n11 163.367
R674 B.n919 B.n11 163.367
R675 B.n919 B.n16 163.367
R676 B.n915 B.n16 163.367
R677 B.n915 B.n18 163.367
R678 B.n911 B.n18 163.367
R679 B.n911 B.n23 163.367
R680 B.n907 B.n23 163.367
R681 B.n907 B.n25 163.367
R682 B.n903 B.n25 163.367
R683 B.n903 B.n30 163.367
R684 B.n899 B.n30 163.367
R685 B.n899 B.n32 163.367
R686 B.n895 B.n32 163.367
R687 B.n895 B.n37 163.367
R688 B.n891 B.n37 163.367
R689 B.n891 B.n39 163.367
R690 B.n887 B.n39 163.367
R691 B.n887 B.n44 163.367
R692 B.n883 B.n44 163.367
R693 B.n883 B.n46 163.367
R694 B.n879 B.n46 163.367
R695 B.n879 B.n51 163.367
R696 B.n875 B.n51 163.367
R697 B.n875 B.n53 163.367
R698 B.n871 B.n53 163.367
R699 B.n871 B.n58 163.367
R700 B.n867 B.n58 163.367
R701 B.n867 B.n60 163.367
R702 B.n482 B.n481 163.367
R703 B.n711 B.n481 163.367
R704 B.n709 B.n708 163.367
R705 B.n705 B.n704 163.367
R706 B.n701 B.n700 163.367
R707 B.n697 B.n696 163.367
R708 B.n693 B.n692 163.367
R709 B.n689 B.n688 163.367
R710 B.n685 B.n684 163.367
R711 B.n681 B.n680 163.367
R712 B.n677 B.n676 163.367
R713 B.n673 B.n672 163.367
R714 B.n669 B.n668 163.367
R715 B.n665 B.n664 163.367
R716 B.n661 B.n660 163.367
R717 B.n657 B.n656 163.367
R718 B.n653 B.n652 163.367
R719 B.n649 B.n648 163.367
R720 B.n645 B.n644 163.367
R721 B.n641 B.n640 163.367
R722 B.n637 B.n636 163.367
R723 B.n633 B.n632 163.367
R724 B.n629 B.n628 163.367
R725 B.n625 B.n624 163.367
R726 B.n621 B.n620 163.367
R727 B.n617 B.n616 163.367
R728 B.n613 B.n612 163.367
R729 B.n608 B.n607 163.367
R730 B.n604 B.n603 163.367
R731 B.n600 B.n599 163.367
R732 B.n596 B.n595 163.367
R733 B.n592 B.n591 163.367
R734 B.n588 B.n587 163.367
R735 B.n584 B.n583 163.367
R736 B.n580 B.n579 163.367
R737 B.n576 B.n575 163.367
R738 B.n572 B.n571 163.367
R739 B.n568 B.n567 163.367
R740 B.n564 B.n563 163.367
R741 B.n560 B.n559 163.367
R742 B.n556 B.n555 163.367
R743 B.n552 B.n551 163.367
R744 B.n548 B.n547 163.367
R745 B.n544 B.n543 163.367
R746 B.n540 B.n539 163.367
R747 B.n536 B.n535 163.367
R748 B.n532 B.n531 163.367
R749 B.n528 B.n527 163.367
R750 B.n524 B.n523 163.367
R751 B.n520 B.n519 163.367
R752 B.n516 B.n515 163.367
R753 B.n512 B.n511 163.367
R754 B.n508 B.n507 163.367
R755 B.n504 B.n503 163.367
R756 B.n500 B.n499 163.367
R757 B.n496 B.n495 163.367
R758 B.n492 B.n491 163.367
R759 B.n488 B.n424 163.367
R760 B.n724 B.n422 163.367
R761 B.n724 B.n416 163.367
R762 B.n732 B.n416 163.367
R763 B.n732 B.n414 163.367
R764 B.n736 B.n414 163.367
R765 B.n736 B.n408 163.367
R766 B.n744 B.n408 163.367
R767 B.n744 B.n406 163.367
R768 B.n748 B.n406 163.367
R769 B.n748 B.n400 163.367
R770 B.n756 B.n400 163.367
R771 B.n756 B.n398 163.367
R772 B.n760 B.n398 163.367
R773 B.n760 B.n392 163.367
R774 B.n768 B.n392 163.367
R775 B.n768 B.n390 163.367
R776 B.n772 B.n390 163.367
R777 B.n772 B.n384 163.367
R778 B.n780 B.n384 163.367
R779 B.n780 B.n382 163.367
R780 B.n784 B.n382 163.367
R781 B.n784 B.n376 163.367
R782 B.n792 B.n376 163.367
R783 B.n792 B.n374 163.367
R784 B.n796 B.n374 163.367
R785 B.n796 B.n368 163.367
R786 B.n804 B.n368 163.367
R787 B.n804 B.n366 163.367
R788 B.n809 B.n366 163.367
R789 B.n809 B.n360 163.367
R790 B.n817 B.n360 163.367
R791 B.n818 B.n817 163.367
R792 B.n818 B.n5 163.367
R793 B.n6 B.n5 163.367
R794 B.n7 B.n6 163.367
R795 B.n823 B.n7 163.367
R796 B.n823 B.n12 163.367
R797 B.n13 B.n12 163.367
R798 B.n14 B.n13 163.367
R799 B.n828 B.n14 163.367
R800 B.n828 B.n19 163.367
R801 B.n20 B.n19 163.367
R802 B.n21 B.n20 163.367
R803 B.n833 B.n21 163.367
R804 B.n833 B.n26 163.367
R805 B.n27 B.n26 163.367
R806 B.n28 B.n27 163.367
R807 B.n838 B.n28 163.367
R808 B.n838 B.n33 163.367
R809 B.n34 B.n33 163.367
R810 B.n35 B.n34 163.367
R811 B.n843 B.n35 163.367
R812 B.n843 B.n40 163.367
R813 B.n41 B.n40 163.367
R814 B.n42 B.n41 163.367
R815 B.n848 B.n42 163.367
R816 B.n848 B.n47 163.367
R817 B.n48 B.n47 163.367
R818 B.n49 B.n48 163.367
R819 B.n853 B.n49 163.367
R820 B.n853 B.n54 163.367
R821 B.n55 B.n54 163.367
R822 B.n56 B.n55 163.367
R823 B.n858 B.n56 163.367
R824 B.n858 B.n61 163.367
R825 B.n62 B.n61 163.367
R826 B.n131 B.n130 163.367
R827 B.n135 B.n134 163.367
R828 B.n139 B.n138 163.367
R829 B.n143 B.n142 163.367
R830 B.n147 B.n146 163.367
R831 B.n151 B.n150 163.367
R832 B.n155 B.n154 163.367
R833 B.n159 B.n158 163.367
R834 B.n163 B.n162 163.367
R835 B.n167 B.n166 163.367
R836 B.n171 B.n170 163.367
R837 B.n175 B.n174 163.367
R838 B.n179 B.n178 163.367
R839 B.n183 B.n182 163.367
R840 B.n187 B.n186 163.367
R841 B.n191 B.n190 163.367
R842 B.n195 B.n194 163.367
R843 B.n199 B.n198 163.367
R844 B.n203 B.n202 163.367
R845 B.n207 B.n206 163.367
R846 B.n211 B.n210 163.367
R847 B.n215 B.n214 163.367
R848 B.n219 B.n218 163.367
R849 B.n223 B.n222 163.367
R850 B.n227 B.n226 163.367
R851 B.n231 B.n230 163.367
R852 B.n235 B.n234 163.367
R853 B.n239 B.n238 163.367
R854 B.n243 B.n242 163.367
R855 B.n247 B.n246 163.367
R856 B.n251 B.n250 163.367
R857 B.n256 B.n255 163.367
R858 B.n260 B.n259 163.367
R859 B.n264 B.n263 163.367
R860 B.n268 B.n267 163.367
R861 B.n272 B.n271 163.367
R862 B.n276 B.n275 163.367
R863 B.n280 B.n279 163.367
R864 B.n284 B.n283 163.367
R865 B.n288 B.n287 163.367
R866 B.n292 B.n291 163.367
R867 B.n296 B.n295 163.367
R868 B.n300 B.n299 163.367
R869 B.n304 B.n303 163.367
R870 B.n308 B.n307 163.367
R871 B.n312 B.n311 163.367
R872 B.n316 B.n315 163.367
R873 B.n320 B.n319 163.367
R874 B.n324 B.n323 163.367
R875 B.n328 B.n327 163.367
R876 B.n332 B.n331 163.367
R877 B.n336 B.n335 163.367
R878 B.n340 B.n339 163.367
R879 B.n344 B.n343 163.367
R880 B.n348 B.n347 163.367
R881 B.n352 B.n351 163.367
R882 B.n356 B.n355 163.367
R883 B.n863 B.n121 163.367
R884 B.n486 B.n485 82.2308
R885 B.n484 B.n483 82.2308
R886 B.n125 B.n124 82.2308
R887 B.n123 B.n122 82.2308
R888 B.n717 B.n716 71.676
R889 B.n711 B.n425 71.676
R890 B.n708 B.n426 71.676
R891 B.n704 B.n427 71.676
R892 B.n700 B.n428 71.676
R893 B.n696 B.n429 71.676
R894 B.n692 B.n430 71.676
R895 B.n688 B.n431 71.676
R896 B.n684 B.n432 71.676
R897 B.n680 B.n433 71.676
R898 B.n676 B.n434 71.676
R899 B.n672 B.n435 71.676
R900 B.n668 B.n436 71.676
R901 B.n664 B.n437 71.676
R902 B.n660 B.n438 71.676
R903 B.n656 B.n439 71.676
R904 B.n652 B.n440 71.676
R905 B.n648 B.n441 71.676
R906 B.n644 B.n442 71.676
R907 B.n640 B.n443 71.676
R908 B.n636 B.n444 71.676
R909 B.n632 B.n445 71.676
R910 B.n628 B.n446 71.676
R911 B.n624 B.n447 71.676
R912 B.n620 B.n448 71.676
R913 B.n616 B.n449 71.676
R914 B.n612 B.n450 71.676
R915 B.n607 B.n451 71.676
R916 B.n603 B.n452 71.676
R917 B.n599 B.n453 71.676
R918 B.n595 B.n454 71.676
R919 B.n591 B.n455 71.676
R920 B.n587 B.n456 71.676
R921 B.n583 B.n457 71.676
R922 B.n579 B.n458 71.676
R923 B.n575 B.n459 71.676
R924 B.n571 B.n460 71.676
R925 B.n567 B.n461 71.676
R926 B.n563 B.n462 71.676
R927 B.n559 B.n463 71.676
R928 B.n555 B.n464 71.676
R929 B.n551 B.n465 71.676
R930 B.n547 B.n466 71.676
R931 B.n543 B.n467 71.676
R932 B.n539 B.n468 71.676
R933 B.n535 B.n469 71.676
R934 B.n531 B.n470 71.676
R935 B.n527 B.n471 71.676
R936 B.n523 B.n472 71.676
R937 B.n519 B.n473 71.676
R938 B.n515 B.n474 71.676
R939 B.n511 B.n475 71.676
R940 B.n507 B.n476 71.676
R941 B.n503 B.n477 71.676
R942 B.n499 B.n478 71.676
R943 B.n495 B.n479 71.676
R944 B.n491 B.n480 71.676
R945 B.n719 B.n424 71.676
R946 B.n127 B.n63 71.676
R947 B.n131 B.n64 71.676
R948 B.n135 B.n65 71.676
R949 B.n139 B.n66 71.676
R950 B.n143 B.n67 71.676
R951 B.n147 B.n68 71.676
R952 B.n151 B.n69 71.676
R953 B.n155 B.n70 71.676
R954 B.n159 B.n71 71.676
R955 B.n163 B.n72 71.676
R956 B.n167 B.n73 71.676
R957 B.n171 B.n74 71.676
R958 B.n175 B.n75 71.676
R959 B.n179 B.n76 71.676
R960 B.n183 B.n77 71.676
R961 B.n187 B.n78 71.676
R962 B.n191 B.n79 71.676
R963 B.n195 B.n80 71.676
R964 B.n199 B.n81 71.676
R965 B.n203 B.n82 71.676
R966 B.n207 B.n83 71.676
R967 B.n211 B.n84 71.676
R968 B.n215 B.n85 71.676
R969 B.n219 B.n86 71.676
R970 B.n223 B.n87 71.676
R971 B.n227 B.n88 71.676
R972 B.n231 B.n89 71.676
R973 B.n235 B.n90 71.676
R974 B.n239 B.n91 71.676
R975 B.n243 B.n92 71.676
R976 B.n247 B.n93 71.676
R977 B.n251 B.n94 71.676
R978 B.n256 B.n95 71.676
R979 B.n260 B.n96 71.676
R980 B.n264 B.n97 71.676
R981 B.n268 B.n98 71.676
R982 B.n272 B.n99 71.676
R983 B.n276 B.n100 71.676
R984 B.n280 B.n101 71.676
R985 B.n284 B.n102 71.676
R986 B.n288 B.n103 71.676
R987 B.n292 B.n104 71.676
R988 B.n296 B.n105 71.676
R989 B.n300 B.n106 71.676
R990 B.n304 B.n107 71.676
R991 B.n308 B.n108 71.676
R992 B.n312 B.n109 71.676
R993 B.n316 B.n110 71.676
R994 B.n320 B.n111 71.676
R995 B.n324 B.n112 71.676
R996 B.n328 B.n113 71.676
R997 B.n332 B.n114 71.676
R998 B.n336 B.n115 71.676
R999 B.n340 B.n116 71.676
R1000 B.n344 B.n117 71.676
R1001 B.n348 B.n118 71.676
R1002 B.n352 B.n119 71.676
R1003 B.n356 B.n120 71.676
R1004 B.n121 B.n120 71.676
R1005 B.n355 B.n119 71.676
R1006 B.n351 B.n118 71.676
R1007 B.n347 B.n117 71.676
R1008 B.n343 B.n116 71.676
R1009 B.n339 B.n115 71.676
R1010 B.n335 B.n114 71.676
R1011 B.n331 B.n113 71.676
R1012 B.n327 B.n112 71.676
R1013 B.n323 B.n111 71.676
R1014 B.n319 B.n110 71.676
R1015 B.n315 B.n109 71.676
R1016 B.n311 B.n108 71.676
R1017 B.n307 B.n107 71.676
R1018 B.n303 B.n106 71.676
R1019 B.n299 B.n105 71.676
R1020 B.n295 B.n104 71.676
R1021 B.n291 B.n103 71.676
R1022 B.n287 B.n102 71.676
R1023 B.n283 B.n101 71.676
R1024 B.n279 B.n100 71.676
R1025 B.n275 B.n99 71.676
R1026 B.n271 B.n98 71.676
R1027 B.n267 B.n97 71.676
R1028 B.n263 B.n96 71.676
R1029 B.n259 B.n95 71.676
R1030 B.n255 B.n94 71.676
R1031 B.n250 B.n93 71.676
R1032 B.n246 B.n92 71.676
R1033 B.n242 B.n91 71.676
R1034 B.n238 B.n90 71.676
R1035 B.n234 B.n89 71.676
R1036 B.n230 B.n88 71.676
R1037 B.n226 B.n87 71.676
R1038 B.n222 B.n86 71.676
R1039 B.n218 B.n85 71.676
R1040 B.n214 B.n84 71.676
R1041 B.n210 B.n83 71.676
R1042 B.n206 B.n82 71.676
R1043 B.n202 B.n81 71.676
R1044 B.n198 B.n80 71.676
R1045 B.n194 B.n79 71.676
R1046 B.n190 B.n78 71.676
R1047 B.n186 B.n77 71.676
R1048 B.n182 B.n76 71.676
R1049 B.n178 B.n75 71.676
R1050 B.n174 B.n74 71.676
R1051 B.n170 B.n73 71.676
R1052 B.n166 B.n72 71.676
R1053 B.n162 B.n71 71.676
R1054 B.n158 B.n70 71.676
R1055 B.n154 B.n69 71.676
R1056 B.n150 B.n68 71.676
R1057 B.n146 B.n67 71.676
R1058 B.n142 B.n66 71.676
R1059 B.n138 B.n65 71.676
R1060 B.n134 B.n64 71.676
R1061 B.n130 B.n63 71.676
R1062 B.n717 B.n482 71.676
R1063 B.n709 B.n425 71.676
R1064 B.n705 B.n426 71.676
R1065 B.n701 B.n427 71.676
R1066 B.n697 B.n428 71.676
R1067 B.n693 B.n429 71.676
R1068 B.n689 B.n430 71.676
R1069 B.n685 B.n431 71.676
R1070 B.n681 B.n432 71.676
R1071 B.n677 B.n433 71.676
R1072 B.n673 B.n434 71.676
R1073 B.n669 B.n435 71.676
R1074 B.n665 B.n436 71.676
R1075 B.n661 B.n437 71.676
R1076 B.n657 B.n438 71.676
R1077 B.n653 B.n439 71.676
R1078 B.n649 B.n440 71.676
R1079 B.n645 B.n441 71.676
R1080 B.n641 B.n442 71.676
R1081 B.n637 B.n443 71.676
R1082 B.n633 B.n444 71.676
R1083 B.n629 B.n445 71.676
R1084 B.n625 B.n446 71.676
R1085 B.n621 B.n447 71.676
R1086 B.n617 B.n448 71.676
R1087 B.n613 B.n449 71.676
R1088 B.n608 B.n450 71.676
R1089 B.n604 B.n451 71.676
R1090 B.n600 B.n452 71.676
R1091 B.n596 B.n453 71.676
R1092 B.n592 B.n454 71.676
R1093 B.n588 B.n455 71.676
R1094 B.n584 B.n456 71.676
R1095 B.n580 B.n457 71.676
R1096 B.n576 B.n458 71.676
R1097 B.n572 B.n459 71.676
R1098 B.n568 B.n460 71.676
R1099 B.n564 B.n461 71.676
R1100 B.n560 B.n462 71.676
R1101 B.n556 B.n463 71.676
R1102 B.n552 B.n464 71.676
R1103 B.n548 B.n465 71.676
R1104 B.n544 B.n466 71.676
R1105 B.n540 B.n467 71.676
R1106 B.n536 B.n468 71.676
R1107 B.n532 B.n469 71.676
R1108 B.n528 B.n470 71.676
R1109 B.n524 B.n471 71.676
R1110 B.n520 B.n472 71.676
R1111 B.n516 B.n473 71.676
R1112 B.n512 B.n474 71.676
R1113 B.n508 B.n475 71.676
R1114 B.n504 B.n476 71.676
R1115 B.n500 B.n477 71.676
R1116 B.n496 B.n478 71.676
R1117 B.n492 B.n479 71.676
R1118 B.n488 B.n480 71.676
R1119 B.n720 B.n719 71.676
R1120 B.n718 B.n421 65.5105
R1121 B.n865 B.n864 65.5105
R1122 B.n487 B.n486 59.5399
R1123 B.n610 B.n484 59.5399
R1124 B.n126 B.n125 59.5399
R1125 B.n253 B.n123 59.5399
R1126 B.n725 B.n421 35.0767
R1127 B.n725 B.n417 35.0767
R1128 B.n731 B.n417 35.0767
R1129 B.n731 B.n413 35.0767
R1130 B.n737 B.n413 35.0767
R1131 B.n737 B.n409 35.0767
R1132 B.n743 B.n409 35.0767
R1133 B.n743 B.n405 35.0767
R1134 B.n749 B.n405 35.0767
R1135 B.n755 B.n401 35.0767
R1136 B.n755 B.n397 35.0767
R1137 B.n761 B.n397 35.0767
R1138 B.n761 B.n393 35.0767
R1139 B.n767 B.n393 35.0767
R1140 B.n767 B.n389 35.0767
R1141 B.n773 B.n389 35.0767
R1142 B.n773 B.n385 35.0767
R1143 B.n779 B.n385 35.0767
R1144 B.n779 B.n381 35.0767
R1145 B.n785 B.n381 35.0767
R1146 B.n785 B.n377 35.0767
R1147 B.n791 B.n377 35.0767
R1148 B.n791 B.n373 35.0767
R1149 B.n797 B.n373 35.0767
R1150 B.n803 B.n369 35.0767
R1151 B.n803 B.n365 35.0767
R1152 B.n810 B.n365 35.0767
R1153 B.n810 B.n361 35.0767
R1154 B.n816 B.n361 35.0767
R1155 B.n816 B.n4 35.0767
R1156 B.n930 B.n4 35.0767
R1157 B.n930 B.n929 35.0767
R1158 B.n929 B.n928 35.0767
R1159 B.n928 B.n8 35.0767
R1160 B.n922 B.n8 35.0767
R1161 B.n922 B.n921 35.0767
R1162 B.n921 B.n920 35.0767
R1163 B.n920 B.n15 35.0767
R1164 B.n914 B.n913 35.0767
R1165 B.n913 B.n912 35.0767
R1166 B.n912 B.n22 35.0767
R1167 B.n906 B.n22 35.0767
R1168 B.n906 B.n905 35.0767
R1169 B.n905 B.n904 35.0767
R1170 B.n904 B.n29 35.0767
R1171 B.n898 B.n29 35.0767
R1172 B.n898 B.n897 35.0767
R1173 B.n897 B.n896 35.0767
R1174 B.n896 B.n36 35.0767
R1175 B.n890 B.n36 35.0767
R1176 B.n890 B.n889 35.0767
R1177 B.n889 B.n888 35.0767
R1178 B.n888 B.n43 35.0767
R1179 B.n882 B.n881 35.0767
R1180 B.n881 B.n880 35.0767
R1181 B.n880 B.n50 35.0767
R1182 B.n874 B.n50 35.0767
R1183 B.n874 B.n873 35.0767
R1184 B.n873 B.n872 35.0767
R1185 B.n872 B.n57 35.0767
R1186 B.n866 B.n57 35.0767
R1187 B.n866 B.n865 35.0767
R1188 B.n128 B.n59 31.0639
R1189 B.n862 B.n861 31.0639
R1190 B.n722 B.n721 31.0639
R1191 B.n715 B.n419 31.0639
R1192 B.t0 B.n369 29.4026
R1193 B.t1 B.n15 29.4026
R1194 B.t3 B.n401 18.0544
R1195 B.t10 B.n43 18.0544
R1196 B B.n932 18.0485
R1197 B.n749 B.t3 17.0228
R1198 B.n882 B.t10 17.0228
R1199 B.n129 B.n128 10.6151
R1200 B.n132 B.n129 10.6151
R1201 B.n133 B.n132 10.6151
R1202 B.n136 B.n133 10.6151
R1203 B.n137 B.n136 10.6151
R1204 B.n140 B.n137 10.6151
R1205 B.n141 B.n140 10.6151
R1206 B.n144 B.n141 10.6151
R1207 B.n145 B.n144 10.6151
R1208 B.n148 B.n145 10.6151
R1209 B.n149 B.n148 10.6151
R1210 B.n152 B.n149 10.6151
R1211 B.n153 B.n152 10.6151
R1212 B.n156 B.n153 10.6151
R1213 B.n157 B.n156 10.6151
R1214 B.n160 B.n157 10.6151
R1215 B.n161 B.n160 10.6151
R1216 B.n164 B.n161 10.6151
R1217 B.n165 B.n164 10.6151
R1218 B.n168 B.n165 10.6151
R1219 B.n169 B.n168 10.6151
R1220 B.n172 B.n169 10.6151
R1221 B.n173 B.n172 10.6151
R1222 B.n176 B.n173 10.6151
R1223 B.n177 B.n176 10.6151
R1224 B.n180 B.n177 10.6151
R1225 B.n181 B.n180 10.6151
R1226 B.n184 B.n181 10.6151
R1227 B.n185 B.n184 10.6151
R1228 B.n188 B.n185 10.6151
R1229 B.n189 B.n188 10.6151
R1230 B.n192 B.n189 10.6151
R1231 B.n193 B.n192 10.6151
R1232 B.n196 B.n193 10.6151
R1233 B.n197 B.n196 10.6151
R1234 B.n200 B.n197 10.6151
R1235 B.n201 B.n200 10.6151
R1236 B.n204 B.n201 10.6151
R1237 B.n205 B.n204 10.6151
R1238 B.n208 B.n205 10.6151
R1239 B.n209 B.n208 10.6151
R1240 B.n212 B.n209 10.6151
R1241 B.n213 B.n212 10.6151
R1242 B.n216 B.n213 10.6151
R1243 B.n217 B.n216 10.6151
R1244 B.n220 B.n217 10.6151
R1245 B.n221 B.n220 10.6151
R1246 B.n224 B.n221 10.6151
R1247 B.n225 B.n224 10.6151
R1248 B.n228 B.n225 10.6151
R1249 B.n229 B.n228 10.6151
R1250 B.n232 B.n229 10.6151
R1251 B.n233 B.n232 10.6151
R1252 B.n237 B.n236 10.6151
R1253 B.n240 B.n237 10.6151
R1254 B.n241 B.n240 10.6151
R1255 B.n244 B.n241 10.6151
R1256 B.n245 B.n244 10.6151
R1257 B.n248 B.n245 10.6151
R1258 B.n249 B.n248 10.6151
R1259 B.n252 B.n249 10.6151
R1260 B.n257 B.n254 10.6151
R1261 B.n258 B.n257 10.6151
R1262 B.n261 B.n258 10.6151
R1263 B.n262 B.n261 10.6151
R1264 B.n265 B.n262 10.6151
R1265 B.n266 B.n265 10.6151
R1266 B.n269 B.n266 10.6151
R1267 B.n270 B.n269 10.6151
R1268 B.n273 B.n270 10.6151
R1269 B.n274 B.n273 10.6151
R1270 B.n277 B.n274 10.6151
R1271 B.n278 B.n277 10.6151
R1272 B.n281 B.n278 10.6151
R1273 B.n282 B.n281 10.6151
R1274 B.n285 B.n282 10.6151
R1275 B.n286 B.n285 10.6151
R1276 B.n289 B.n286 10.6151
R1277 B.n290 B.n289 10.6151
R1278 B.n293 B.n290 10.6151
R1279 B.n294 B.n293 10.6151
R1280 B.n297 B.n294 10.6151
R1281 B.n298 B.n297 10.6151
R1282 B.n301 B.n298 10.6151
R1283 B.n302 B.n301 10.6151
R1284 B.n305 B.n302 10.6151
R1285 B.n306 B.n305 10.6151
R1286 B.n309 B.n306 10.6151
R1287 B.n310 B.n309 10.6151
R1288 B.n313 B.n310 10.6151
R1289 B.n314 B.n313 10.6151
R1290 B.n317 B.n314 10.6151
R1291 B.n318 B.n317 10.6151
R1292 B.n321 B.n318 10.6151
R1293 B.n322 B.n321 10.6151
R1294 B.n325 B.n322 10.6151
R1295 B.n326 B.n325 10.6151
R1296 B.n329 B.n326 10.6151
R1297 B.n330 B.n329 10.6151
R1298 B.n333 B.n330 10.6151
R1299 B.n334 B.n333 10.6151
R1300 B.n337 B.n334 10.6151
R1301 B.n338 B.n337 10.6151
R1302 B.n341 B.n338 10.6151
R1303 B.n342 B.n341 10.6151
R1304 B.n345 B.n342 10.6151
R1305 B.n346 B.n345 10.6151
R1306 B.n349 B.n346 10.6151
R1307 B.n350 B.n349 10.6151
R1308 B.n353 B.n350 10.6151
R1309 B.n354 B.n353 10.6151
R1310 B.n357 B.n354 10.6151
R1311 B.n358 B.n357 10.6151
R1312 B.n862 B.n358 10.6151
R1313 B.n723 B.n722 10.6151
R1314 B.n723 B.n415 10.6151
R1315 B.n733 B.n415 10.6151
R1316 B.n734 B.n733 10.6151
R1317 B.n735 B.n734 10.6151
R1318 B.n735 B.n407 10.6151
R1319 B.n745 B.n407 10.6151
R1320 B.n746 B.n745 10.6151
R1321 B.n747 B.n746 10.6151
R1322 B.n747 B.n399 10.6151
R1323 B.n757 B.n399 10.6151
R1324 B.n758 B.n757 10.6151
R1325 B.n759 B.n758 10.6151
R1326 B.n759 B.n391 10.6151
R1327 B.n769 B.n391 10.6151
R1328 B.n770 B.n769 10.6151
R1329 B.n771 B.n770 10.6151
R1330 B.n771 B.n383 10.6151
R1331 B.n781 B.n383 10.6151
R1332 B.n782 B.n781 10.6151
R1333 B.n783 B.n782 10.6151
R1334 B.n783 B.n375 10.6151
R1335 B.n793 B.n375 10.6151
R1336 B.n794 B.n793 10.6151
R1337 B.n795 B.n794 10.6151
R1338 B.n795 B.n367 10.6151
R1339 B.n805 B.n367 10.6151
R1340 B.n806 B.n805 10.6151
R1341 B.n808 B.n806 10.6151
R1342 B.n808 B.n807 10.6151
R1343 B.n807 B.n359 10.6151
R1344 B.n819 B.n359 10.6151
R1345 B.n820 B.n819 10.6151
R1346 B.n821 B.n820 10.6151
R1347 B.n822 B.n821 10.6151
R1348 B.n824 B.n822 10.6151
R1349 B.n825 B.n824 10.6151
R1350 B.n826 B.n825 10.6151
R1351 B.n827 B.n826 10.6151
R1352 B.n829 B.n827 10.6151
R1353 B.n830 B.n829 10.6151
R1354 B.n831 B.n830 10.6151
R1355 B.n832 B.n831 10.6151
R1356 B.n834 B.n832 10.6151
R1357 B.n835 B.n834 10.6151
R1358 B.n836 B.n835 10.6151
R1359 B.n837 B.n836 10.6151
R1360 B.n839 B.n837 10.6151
R1361 B.n840 B.n839 10.6151
R1362 B.n841 B.n840 10.6151
R1363 B.n842 B.n841 10.6151
R1364 B.n844 B.n842 10.6151
R1365 B.n845 B.n844 10.6151
R1366 B.n846 B.n845 10.6151
R1367 B.n847 B.n846 10.6151
R1368 B.n849 B.n847 10.6151
R1369 B.n850 B.n849 10.6151
R1370 B.n851 B.n850 10.6151
R1371 B.n852 B.n851 10.6151
R1372 B.n854 B.n852 10.6151
R1373 B.n855 B.n854 10.6151
R1374 B.n856 B.n855 10.6151
R1375 B.n857 B.n856 10.6151
R1376 B.n859 B.n857 10.6151
R1377 B.n860 B.n859 10.6151
R1378 B.n861 B.n860 10.6151
R1379 B.n715 B.n714 10.6151
R1380 B.n714 B.n713 10.6151
R1381 B.n713 B.n712 10.6151
R1382 B.n712 B.n710 10.6151
R1383 B.n710 B.n707 10.6151
R1384 B.n707 B.n706 10.6151
R1385 B.n706 B.n703 10.6151
R1386 B.n703 B.n702 10.6151
R1387 B.n702 B.n699 10.6151
R1388 B.n699 B.n698 10.6151
R1389 B.n698 B.n695 10.6151
R1390 B.n695 B.n694 10.6151
R1391 B.n694 B.n691 10.6151
R1392 B.n691 B.n690 10.6151
R1393 B.n690 B.n687 10.6151
R1394 B.n687 B.n686 10.6151
R1395 B.n686 B.n683 10.6151
R1396 B.n683 B.n682 10.6151
R1397 B.n682 B.n679 10.6151
R1398 B.n679 B.n678 10.6151
R1399 B.n678 B.n675 10.6151
R1400 B.n675 B.n674 10.6151
R1401 B.n674 B.n671 10.6151
R1402 B.n671 B.n670 10.6151
R1403 B.n670 B.n667 10.6151
R1404 B.n667 B.n666 10.6151
R1405 B.n666 B.n663 10.6151
R1406 B.n663 B.n662 10.6151
R1407 B.n662 B.n659 10.6151
R1408 B.n659 B.n658 10.6151
R1409 B.n658 B.n655 10.6151
R1410 B.n655 B.n654 10.6151
R1411 B.n654 B.n651 10.6151
R1412 B.n651 B.n650 10.6151
R1413 B.n650 B.n647 10.6151
R1414 B.n647 B.n646 10.6151
R1415 B.n646 B.n643 10.6151
R1416 B.n643 B.n642 10.6151
R1417 B.n642 B.n639 10.6151
R1418 B.n639 B.n638 10.6151
R1419 B.n638 B.n635 10.6151
R1420 B.n635 B.n634 10.6151
R1421 B.n634 B.n631 10.6151
R1422 B.n631 B.n630 10.6151
R1423 B.n630 B.n627 10.6151
R1424 B.n627 B.n626 10.6151
R1425 B.n626 B.n623 10.6151
R1426 B.n623 B.n622 10.6151
R1427 B.n622 B.n619 10.6151
R1428 B.n619 B.n618 10.6151
R1429 B.n618 B.n615 10.6151
R1430 B.n615 B.n614 10.6151
R1431 B.n614 B.n611 10.6151
R1432 B.n609 B.n606 10.6151
R1433 B.n606 B.n605 10.6151
R1434 B.n605 B.n602 10.6151
R1435 B.n602 B.n601 10.6151
R1436 B.n601 B.n598 10.6151
R1437 B.n598 B.n597 10.6151
R1438 B.n597 B.n594 10.6151
R1439 B.n594 B.n593 10.6151
R1440 B.n590 B.n589 10.6151
R1441 B.n589 B.n586 10.6151
R1442 B.n586 B.n585 10.6151
R1443 B.n585 B.n582 10.6151
R1444 B.n582 B.n581 10.6151
R1445 B.n581 B.n578 10.6151
R1446 B.n578 B.n577 10.6151
R1447 B.n577 B.n574 10.6151
R1448 B.n574 B.n573 10.6151
R1449 B.n573 B.n570 10.6151
R1450 B.n570 B.n569 10.6151
R1451 B.n569 B.n566 10.6151
R1452 B.n566 B.n565 10.6151
R1453 B.n565 B.n562 10.6151
R1454 B.n562 B.n561 10.6151
R1455 B.n561 B.n558 10.6151
R1456 B.n558 B.n557 10.6151
R1457 B.n557 B.n554 10.6151
R1458 B.n554 B.n553 10.6151
R1459 B.n553 B.n550 10.6151
R1460 B.n550 B.n549 10.6151
R1461 B.n549 B.n546 10.6151
R1462 B.n546 B.n545 10.6151
R1463 B.n545 B.n542 10.6151
R1464 B.n542 B.n541 10.6151
R1465 B.n541 B.n538 10.6151
R1466 B.n538 B.n537 10.6151
R1467 B.n537 B.n534 10.6151
R1468 B.n534 B.n533 10.6151
R1469 B.n533 B.n530 10.6151
R1470 B.n530 B.n529 10.6151
R1471 B.n529 B.n526 10.6151
R1472 B.n526 B.n525 10.6151
R1473 B.n525 B.n522 10.6151
R1474 B.n522 B.n521 10.6151
R1475 B.n521 B.n518 10.6151
R1476 B.n518 B.n517 10.6151
R1477 B.n517 B.n514 10.6151
R1478 B.n514 B.n513 10.6151
R1479 B.n513 B.n510 10.6151
R1480 B.n510 B.n509 10.6151
R1481 B.n509 B.n506 10.6151
R1482 B.n506 B.n505 10.6151
R1483 B.n505 B.n502 10.6151
R1484 B.n502 B.n501 10.6151
R1485 B.n501 B.n498 10.6151
R1486 B.n498 B.n497 10.6151
R1487 B.n497 B.n494 10.6151
R1488 B.n494 B.n493 10.6151
R1489 B.n493 B.n490 10.6151
R1490 B.n490 B.n489 10.6151
R1491 B.n489 B.n423 10.6151
R1492 B.n721 B.n423 10.6151
R1493 B.n727 B.n419 10.6151
R1494 B.n728 B.n727 10.6151
R1495 B.n729 B.n728 10.6151
R1496 B.n729 B.n411 10.6151
R1497 B.n739 B.n411 10.6151
R1498 B.n740 B.n739 10.6151
R1499 B.n741 B.n740 10.6151
R1500 B.n741 B.n403 10.6151
R1501 B.n751 B.n403 10.6151
R1502 B.n752 B.n751 10.6151
R1503 B.n753 B.n752 10.6151
R1504 B.n753 B.n395 10.6151
R1505 B.n763 B.n395 10.6151
R1506 B.n764 B.n763 10.6151
R1507 B.n765 B.n764 10.6151
R1508 B.n765 B.n387 10.6151
R1509 B.n775 B.n387 10.6151
R1510 B.n776 B.n775 10.6151
R1511 B.n777 B.n776 10.6151
R1512 B.n777 B.n379 10.6151
R1513 B.n787 B.n379 10.6151
R1514 B.n788 B.n787 10.6151
R1515 B.n789 B.n788 10.6151
R1516 B.n789 B.n371 10.6151
R1517 B.n799 B.n371 10.6151
R1518 B.n800 B.n799 10.6151
R1519 B.n801 B.n800 10.6151
R1520 B.n801 B.n363 10.6151
R1521 B.n812 B.n363 10.6151
R1522 B.n813 B.n812 10.6151
R1523 B.n814 B.n813 10.6151
R1524 B.n814 B.n0 10.6151
R1525 B.n926 B.n1 10.6151
R1526 B.n926 B.n925 10.6151
R1527 B.n925 B.n924 10.6151
R1528 B.n924 B.n10 10.6151
R1529 B.n918 B.n10 10.6151
R1530 B.n918 B.n917 10.6151
R1531 B.n917 B.n916 10.6151
R1532 B.n916 B.n17 10.6151
R1533 B.n910 B.n17 10.6151
R1534 B.n910 B.n909 10.6151
R1535 B.n909 B.n908 10.6151
R1536 B.n908 B.n24 10.6151
R1537 B.n902 B.n24 10.6151
R1538 B.n902 B.n901 10.6151
R1539 B.n901 B.n900 10.6151
R1540 B.n900 B.n31 10.6151
R1541 B.n894 B.n31 10.6151
R1542 B.n894 B.n893 10.6151
R1543 B.n893 B.n892 10.6151
R1544 B.n892 B.n38 10.6151
R1545 B.n886 B.n38 10.6151
R1546 B.n886 B.n885 10.6151
R1547 B.n885 B.n884 10.6151
R1548 B.n884 B.n45 10.6151
R1549 B.n878 B.n45 10.6151
R1550 B.n878 B.n877 10.6151
R1551 B.n877 B.n876 10.6151
R1552 B.n876 B.n52 10.6151
R1553 B.n870 B.n52 10.6151
R1554 B.n870 B.n869 10.6151
R1555 B.n869 B.n868 10.6151
R1556 B.n868 B.n59 10.6151
R1557 B.n236 B.n126 6.5566
R1558 B.n253 B.n252 6.5566
R1559 B.n610 B.n609 6.5566
R1560 B.n593 B.n487 6.5566
R1561 B.n797 B.t0 5.67459
R1562 B.n914 B.t1 5.67459
R1563 B.n233 B.n126 4.05904
R1564 B.n254 B.n253 4.05904
R1565 B.n611 B.n610 4.05904
R1566 B.n590 B.n487 4.05904
R1567 B.n932 B.n0 2.81026
R1568 B.n932 B.n1 2.81026
R1569 VN VN.t1 184.976
R1570 VN VN.t0 134.585
R1571 VTAIL.n354 VTAIL.n270 289.615
R1572 VTAIL.n84 VTAIL.n0 289.615
R1573 VTAIL.n264 VTAIL.n180 289.615
R1574 VTAIL.n174 VTAIL.n90 289.615
R1575 VTAIL.n298 VTAIL.n297 185
R1576 VTAIL.n303 VTAIL.n302 185
R1577 VTAIL.n305 VTAIL.n304 185
R1578 VTAIL.n294 VTAIL.n293 185
R1579 VTAIL.n311 VTAIL.n310 185
R1580 VTAIL.n313 VTAIL.n312 185
R1581 VTAIL.n290 VTAIL.n289 185
R1582 VTAIL.n319 VTAIL.n318 185
R1583 VTAIL.n321 VTAIL.n320 185
R1584 VTAIL.n286 VTAIL.n285 185
R1585 VTAIL.n327 VTAIL.n326 185
R1586 VTAIL.n329 VTAIL.n328 185
R1587 VTAIL.n282 VTAIL.n281 185
R1588 VTAIL.n335 VTAIL.n334 185
R1589 VTAIL.n337 VTAIL.n336 185
R1590 VTAIL.n278 VTAIL.n277 185
R1591 VTAIL.n344 VTAIL.n343 185
R1592 VTAIL.n345 VTAIL.n276 185
R1593 VTAIL.n347 VTAIL.n346 185
R1594 VTAIL.n274 VTAIL.n273 185
R1595 VTAIL.n353 VTAIL.n352 185
R1596 VTAIL.n355 VTAIL.n354 185
R1597 VTAIL.n28 VTAIL.n27 185
R1598 VTAIL.n33 VTAIL.n32 185
R1599 VTAIL.n35 VTAIL.n34 185
R1600 VTAIL.n24 VTAIL.n23 185
R1601 VTAIL.n41 VTAIL.n40 185
R1602 VTAIL.n43 VTAIL.n42 185
R1603 VTAIL.n20 VTAIL.n19 185
R1604 VTAIL.n49 VTAIL.n48 185
R1605 VTAIL.n51 VTAIL.n50 185
R1606 VTAIL.n16 VTAIL.n15 185
R1607 VTAIL.n57 VTAIL.n56 185
R1608 VTAIL.n59 VTAIL.n58 185
R1609 VTAIL.n12 VTAIL.n11 185
R1610 VTAIL.n65 VTAIL.n64 185
R1611 VTAIL.n67 VTAIL.n66 185
R1612 VTAIL.n8 VTAIL.n7 185
R1613 VTAIL.n74 VTAIL.n73 185
R1614 VTAIL.n75 VTAIL.n6 185
R1615 VTAIL.n77 VTAIL.n76 185
R1616 VTAIL.n4 VTAIL.n3 185
R1617 VTAIL.n83 VTAIL.n82 185
R1618 VTAIL.n85 VTAIL.n84 185
R1619 VTAIL.n265 VTAIL.n264 185
R1620 VTAIL.n263 VTAIL.n262 185
R1621 VTAIL.n184 VTAIL.n183 185
R1622 VTAIL.n257 VTAIL.n256 185
R1623 VTAIL.n255 VTAIL.n186 185
R1624 VTAIL.n254 VTAIL.n253 185
R1625 VTAIL.n189 VTAIL.n187 185
R1626 VTAIL.n248 VTAIL.n247 185
R1627 VTAIL.n246 VTAIL.n245 185
R1628 VTAIL.n193 VTAIL.n192 185
R1629 VTAIL.n240 VTAIL.n239 185
R1630 VTAIL.n238 VTAIL.n237 185
R1631 VTAIL.n197 VTAIL.n196 185
R1632 VTAIL.n232 VTAIL.n231 185
R1633 VTAIL.n230 VTAIL.n229 185
R1634 VTAIL.n201 VTAIL.n200 185
R1635 VTAIL.n224 VTAIL.n223 185
R1636 VTAIL.n222 VTAIL.n221 185
R1637 VTAIL.n205 VTAIL.n204 185
R1638 VTAIL.n216 VTAIL.n215 185
R1639 VTAIL.n214 VTAIL.n213 185
R1640 VTAIL.n209 VTAIL.n208 185
R1641 VTAIL.n175 VTAIL.n174 185
R1642 VTAIL.n173 VTAIL.n172 185
R1643 VTAIL.n94 VTAIL.n93 185
R1644 VTAIL.n167 VTAIL.n166 185
R1645 VTAIL.n165 VTAIL.n96 185
R1646 VTAIL.n164 VTAIL.n163 185
R1647 VTAIL.n99 VTAIL.n97 185
R1648 VTAIL.n158 VTAIL.n157 185
R1649 VTAIL.n156 VTAIL.n155 185
R1650 VTAIL.n103 VTAIL.n102 185
R1651 VTAIL.n150 VTAIL.n149 185
R1652 VTAIL.n148 VTAIL.n147 185
R1653 VTAIL.n107 VTAIL.n106 185
R1654 VTAIL.n142 VTAIL.n141 185
R1655 VTAIL.n140 VTAIL.n139 185
R1656 VTAIL.n111 VTAIL.n110 185
R1657 VTAIL.n134 VTAIL.n133 185
R1658 VTAIL.n132 VTAIL.n131 185
R1659 VTAIL.n115 VTAIL.n114 185
R1660 VTAIL.n126 VTAIL.n125 185
R1661 VTAIL.n124 VTAIL.n123 185
R1662 VTAIL.n119 VTAIL.n118 185
R1663 VTAIL.n299 VTAIL.t3 147.659
R1664 VTAIL.n29 VTAIL.t0 147.659
R1665 VTAIL.n210 VTAIL.t1 147.659
R1666 VTAIL.n120 VTAIL.t2 147.659
R1667 VTAIL.n303 VTAIL.n297 104.615
R1668 VTAIL.n304 VTAIL.n303 104.615
R1669 VTAIL.n304 VTAIL.n293 104.615
R1670 VTAIL.n311 VTAIL.n293 104.615
R1671 VTAIL.n312 VTAIL.n311 104.615
R1672 VTAIL.n312 VTAIL.n289 104.615
R1673 VTAIL.n319 VTAIL.n289 104.615
R1674 VTAIL.n320 VTAIL.n319 104.615
R1675 VTAIL.n320 VTAIL.n285 104.615
R1676 VTAIL.n327 VTAIL.n285 104.615
R1677 VTAIL.n328 VTAIL.n327 104.615
R1678 VTAIL.n328 VTAIL.n281 104.615
R1679 VTAIL.n335 VTAIL.n281 104.615
R1680 VTAIL.n336 VTAIL.n335 104.615
R1681 VTAIL.n336 VTAIL.n277 104.615
R1682 VTAIL.n344 VTAIL.n277 104.615
R1683 VTAIL.n345 VTAIL.n344 104.615
R1684 VTAIL.n346 VTAIL.n345 104.615
R1685 VTAIL.n346 VTAIL.n273 104.615
R1686 VTAIL.n353 VTAIL.n273 104.615
R1687 VTAIL.n354 VTAIL.n353 104.615
R1688 VTAIL.n33 VTAIL.n27 104.615
R1689 VTAIL.n34 VTAIL.n33 104.615
R1690 VTAIL.n34 VTAIL.n23 104.615
R1691 VTAIL.n41 VTAIL.n23 104.615
R1692 VTAIL.n42 VTAIL.n41 104.615
R1693 VTAIL.n42 VTAIL.n19 104.615
R1694 VTAIL.n49 VTAIL.n19 104.615
R1695 VTAIL.n50 VTAIL.n49 104.615
R1696 VTAIL.n50 VTAIL.n15 104.615
R1697 VTAIL.n57 VTAIL.n15 104.615
R1698 VTAIL.n58 VTAIL.n57 104.615
R1699 VTAIL.n58 VTAIL.n11 104.615
R1700 VTAIL.n65 VTAIL.n11 104.615
R1701 VTAIL.n66 VTAIL.n65 104.615
R1702 VTAIL.n66 VTAIL.n7 104.615
R1703 VTAIL.n74 VTAIL.n7 104.615
R1704 VTAIL.n75 VTAIL.n74 104.615
R1705 VTAIL.n76 VTAIL.n75 104.615
R1706 VTAIL.n76 VTAIL.n3 104.615
R1707 VTAIL.n83 VTAIL.n3 104.615
R1708 VTAIL.n84 VTAIL.n83 104.615
R1709 VTAIL.n264 VTAIL.n263 104.615
R1710 VTAIL.n263 VTAIL.n183 104.615
R1711 VTAIL.n256 VTAIL.n183 104.615
R1712 VTAIL.n256 VTAIL.n255 104.615
R1713 VTAIL.n255 VTAIL.n254 104.615
R1714 VTAIL.n254 VTAIL.n187 104.615
R1715 VTAIL.n247 VTAIL.n187 104.615
R1716 VTAIL.n247 VTAIL.n246 104.615
R1717 VTAIL.n246 VTAIL.n192 104.615
R1718 VTAIL.n239 VTAIL.n192 104.615
R1719 VTAIL.n239 VTAIL.n238 104.615
R1720 VTAIL.n238 VTAIL.n196 104.615
R1721 VTAIL.n231 VTAIL.n196 104.615
R1722 VTAIL.n231 VTAIL.n230 104.615
R1723 VTAIL.n230 VTAIL.n200 104.615
R1724 VTAIL.n223 VTAIL.n200 104.615
R1725 VTAIL.n223 VTAIL.n222 104.615
R1726 VTAIL.n222 VTAIL.n204 104.615
R1727 VTAIL.n215 VTAIL.n204 104.615
R1728 VTAIL.n215 VTAIL.n214 104.615
R1729 VTAIL.n214 VTAIL.n208 104.615
R1730 VTAIL.n174 VTAIL.n173 104.615
R1731 VTAIL.n173 VTAIL.n93 104.615
R1732 VTAIL.n166 VTAIL.n93 104.615
R1733 VTAIL.n166 VTAIL.n165 104.615
R1734 VTAIL.n165 VTAIL.n164 104.615
R1735 VTAIL.n164 VTAIL.n97 104.615
R1736 VTAIL.n157 VTAIL.n97 104.615
R1737 VTAIL.n157 VTAIL.n156 104.615
R1738 VTAIL.n156 VTAIL.n102 104.615
R1739 VTAIL.n149 VTAIL.n102 104.615
R1740 VTAIL.n149 VTAIL.n148 104.615
R1741 VTAIL.n148 VTAIL.n106 104.615
R1742 VTAIL.n141 VTAIL.n106 104.615
R1743 VTAIL.n141 VTAIL.n140 104.615
R1744 VTAIL.n140 VTAIL.n110 104.615
R1745 VTAIL.n133 VTAIL.n110 104.615
R1746 VTAIL.n133 VTAIL.n132 104.615
R1747 VTAIL.n132 VTAIL.n114 104.615
R1748 VTAIL.n125 VTAIL.n114 104.615
R1749 VTAIL.n125 VTAIL.n124 104.615
R1750 VTAIL.n124 VTAIL.n118 104.615
R1751 VTAIL.t3 VTAIL.n297 52.3082
R1752 VTAIL.t0 VTAIL.n27 52.3082
R1753 VTAIL.t1 VTAIL.n208 52.3082
R1754 VTAIL.t2 VTAIL.n118 52.3082
R1755 VTAIL.n179 VTAIL.n89 33.5134
R1756 VTAIL.n359 VTAIL.n358 31.6035
R1757 VTAIL.n89 VTAIL.n88 31.6035
R1758 VTAIL.n269 VTAIL.n268 31.6035
R1759 VTAIL.n179 VTAIL.n178 31.6035
R1760 VTAIL.n359 VTAIL.n269 29.8583
R1761 VTAIL.n299 VTAIL.n298 15.6677
R1762 VTAIL.n29 VTAIL.n28 15.6677
R1763 VTAIL.n210 VTAIL.n209 15.6677
R1764 VTAIL.n120 VTAIL.n119 15.6677
R1765 VTAIL.n347 VTAIL.n276 13.1884
R1766 VTAIL.n77 VTAIL.n6 13.1884
R1767 VTAIL.n257 VTAIL.n186 13.1884
R1768 VTAIL.n167 VTAIL.n96 13.1884
R1769 VTAIL.n302 VTAIL.n301 12.8005
R1770 VTAIL.n343 VTAIL.n342 12.8005
R1771 VTAIL.n348 VTAIL.n274 12.8005
R1772 VTAIL.n32 VTAIL.n31 12.8005
R1773 VTAIL.n73 VTAIL.n72 12.8005
R1774 VTAIL.n78 VTAIL.n4 12.8005
R1775 VTAIL.n258 VTAIL.n184 12.8005
R1776 VTAIL.n253 VTAIL.n188 12.8005
R1777 VTAIL.n213 VTAIL.n212 12.8005
R1778 VTAIL.n168 VTAIL.n94 12.8005
R1779 VTAIL.n163 VTAIL.n98 12.8005
R1780 VTAIL.n123 VTAIL.n122 12.8005
R1781 VTAIL.n305 VTAIL.n296 12.0247
R1782 VTAIL.n341 VTAIL.n278 12.0247
R1783 VTAIL.n352 VTAIL.n351 12.0247
R1784 VTAIL.n35 VTAIL.n26 12.0247
R1785 VTAIL.n71 VTAIL.n8 12.0247
R1786 VTAIL.n82 VTAIL.n81 12.0247
R1787 VTAIL.n262 VTAIL.n261 12.0247
R1788 VTAIL.n252 VTAIL.n189 12.0247
R1789 VTAIL.n216 VTAIL.n207 12.0247
R1790 VTAIL.n172 VTAIL.n171 12.0247
R1791 VTAIL.n162 VTAIL.n99 12.0247
R1792 VTAIL.n126 VTAIL.n117 12.0247
R1793 VTAIL.n306 VTAIL.n294 11.249
R1794 VTAIL.n338 VTAIL.n337 11.249
R1795 VTAIL.n355 VTAIL.n272 11.249
R1796 VTAIL.n36 VTAIL.n24 11.249
R1797 VTAIL.n68 VTAIL.n67 11.249
R1798 VTAIL.n85 VTAIL.n2 11.249
R1799 VTAIL.n265 VTAIL.n182 11.249
R1800 VTAIL.n249 VTAIL.n248 11.249
R1801 VTAIL.n217 VTAIL.n205 11.249
R1802 VTAIL.n175 VTAIL.n92 11.249
R1803 VTAIL.n159 VTAIL.n158 11.249
R1804 VTAIL.n127 VTAIL.n115 11.249
R1805 VTAIL.n310 VTAIL.n309 10.4732
R1806 VTAIL.n334 VTAIL.n280 10.4732
R1807 VTAIL.n356 VTAIL.n270 10.4732
R1808 VTAIL.n40 VTAIL.n39 10.4732
R1809 VTAIL.n64 VTAIL.n10 10.4732
R1810 VTAIL.n86 VTAIL.n0 10.4732
R1811 VTAIL.n266 VTAIL.n180 10.4732
R1812 VTAIL.n245 VTAIL.n191 10.4732
R1813 VTAIL.n221 VTAIL.n220 10.4732
R1814 VTAIL.n176 VTAIL.n90 10.4732
R1815 VTAIL.n155 VTAIL.n101 10.4732
R1816 VTAIL.n131 VTAIL.n130 10.4732
R1817 VTAIL.n313 VTAIL.n292 9.69747
R1818 VTAIL.n333 VTAIL.n282 9.69747
R1819 VTAIL.n43 VTAIL.n22 9.69747
R1820 VTAIL.n63 VTAIL.n12 9.69747
R1821 VTAIL.n244 VTAIL.n193 9.69747
R1822 VTAIL.n224 VTAIL.n203 9.69747
R1823 VTAIL.n154 VTAIL.n103 9.69747
R1824 VTAIL.n134 VTAIL.n113 9.69747
R1825 VTAIL.n358 VTAIL.n357 9.45567
R1826 VTAIL.n88 VTAIL.n87 9.45567
R1827 VTAIL.n268 VTAIL.n267 9.45567
R1828 VTAIL.n178 VTAIL.n177 9.45567
R1829 VTAIL.n357 VTAIL.n356 9.3005
R1830 VTAIL.n272 VTAIL.n271 9.3005
R1831 VTAIL.n351 VTAIL.n350 9.3005
R1832 VTAIL.n349 VTAIL.n348 9.3005
R1833 VTAIL.n288 VTAIL.n287 9.3005
R1834 VTAIL.n317 VTAIL.n316 9.3005
R1835 VTAIL.n315 VTAIL.n314 9.3005
R1836 VTAIL.n292 VTAIL.n291 9.3005
R1837 VTAIL.n309 VTAIL.n308 9.3005
R1838 VTAIL.n307 VTAIL.n306 9.3005
R1839 VTAIL.n296 VTAIL.n295 9.3005
R1840 VTAIL.n301 VTAIL.n300 9.3005
R1841 VTAIL.n323 VTAIL.n322 9.3005
R1842 VTAIL.n325 VTAIL.n324 9.3005
R1843 VTAIL.n284 VTAIL.n283 9.3005
R1844 VTAIL.n331 VTAIL.n330 9.3005
R1845 VTAIL.n333 VTAIL.n332 9.3005
R1846 VTAIL.n280 VTAIL.n279 9.3005
R1847 VTAIL.n339 VTAIL.n338 9.3005
R1848 VTAIL.n341 VTAIL.n340 9.3005
R1849 VTAIL.n342 VTAIL.n275 9.3005
R1850 VTAIL.n87 VTAIL.n86 9.3005
R1851 VTAIL.n2 VTAIL.n1 9.3005
R1852 VTAIL.n81 VTAIL.n80 9.3005
R1853 VTAIL.n79 VTAIL.n78 9.3005
R1854 VTAIL.n18 VTAIL.n17 9.3005
R1855 VTAIL.n47 VTAIL.n46 9.3005
R1856 VTAIL.n45 VTAIL.n44 9.3005
R1857 VTAIL.n22 VTAIL.n21 9.3005
R1858 VTAIL.n39 VTAIL.n38 9.3005
R1859 VTAIL.n37 VTAIL.n36 9.3005
R1860 VTAIL.n26 VTAIL.n25 9.3005
R1861 VTAIL.n31 VTAIL.n30 9.3005
R1862 VTAIL.n53 VTAIL.n52 9.3005
R1863 VTAIL.n55 VTAIL.n54 9.3005
R1864 VTAIL.n14 VTAIL.n13 9.3005
R1865 VTAIL.n61 VTAIL.n60 9.3005
R1866 VTAIL.n63 VTAIL.n62 9.3005
R1867 VTAIL.n10 VTAIL.n9 9.3005
R1868 VTAIL.n69 VTAIL.n68 9.3005
R1869 VTAIL.n71 VTAIL.n70 9.3005
R1870 VTAIL.n72 VTAIL.n5 9.3005
R1871 VTAIL.n236 VTAIL.n235 9.3005
R1872 VTAIL.n195 VTAIL.n194 9.3005
R1873 VTAIL.n242 VTAIL.n241 9.3005
R1874 VTAIL.n244 VTAIL.n243 9.3005
R1875 VTAIL.n191 VTAIL.n190 9.3005
R1876 VTAIL.n250 VTAIL.n249 9.3005
R1877 VTAIL.n252 VTAIL.n251 9.3005
R1878 VTAIL.n188 VTAIL.n185 9.3005
R1879 VTAIL.n267 VTAIL.n266 9.3005
R1880 VTAIL.n182 VTAIL.n181 9.3005
R1881 VTAIL.n261 VTAIL.n260 9.3005
R1882 VTAIL.n259 VTAIL.n258 9.3005
R1883 VTAIL.n234 VTAIL.n233 9.3005
R1884 VTAIL.n199 VTAIL.n198 9.3005
R1885 VTAIL.n228 VTAIL.n227 9.3005
R1886 VTAIL.n226 VTAIL.n225 9.3005
R1887 VTAIL.n203 VTAIL.n202 9.3005
R1888 VTAIL.n220 VTAIL.n219 9.3005
R1889 VTAIL.n218 VTAIL.n217 9.3005
R1890 VTAIL.n207 VTAIL.n206 9.3005
R1891 VTAIL.n212 VTAIL.n211 9.3005
R1892 VTAIL.n146 VTAIL.n145 9.3005
R1893 VTAIL.n105 VTAIL.n104 9.3005
R1894 VTAIL.n152 VTAIL.n151 9.3005
R1895 VTAIL.n154 VTAIL.n153 9.3005
R1896 VTAIL.n101 VTAIL.n100 9.3005
R1897 VTAIL.n160 VTAIL.n159 9.3005
R1898 VTAIL.n162 VTAIL.n161 9.3005
R1899 VTAIL.n98 VTAIL.n95 9.3005
R1900 VTAIL.n177 VTAIL.n176 9.3005
R1901 VTAIL.n92 VTAIL.n91 9.3005
R1902 VTAIL.n171 VTAIL.n170 9.3005
R1903 VTAIL.n169 VTAIL.n168 9.3005
R1904 VTAIL.n144 VTAIL.n143 9.3005
R1905 VTAIL.n109 VTAIL.n108 9.3005
R1906 VTAIL.n138 VTAIL.n137 9.3005
R1907 VTAIL.n136 VTAIL.n135 9.3005
R1908 VTAIL.n113 VTAIL.n112 9.3005
R1909 VTAIL.n130 VTAIL.n129 9.3005
R1910 VTAIL.n128 VTAIL.n127 9.3005
R1911 VTAIL.n117 VTAIL.n116 9.3005
R1912 VTAIL.n122 VTAIL.n121 9.3005
R1913 VTAIL.n314 VTAIL.n290 8.92171
R1914 VTAIL.n330 VTAIL.n329 8.92171
R1915 VTAIL.n44 VTAIL.n20 8.92171
R1916 VTAIL.n60 VTAIL.n59 8.92171
R1917 VTAIL.n241 VTAIL.n240 8.92171
R1918 VTAIL.n225 VTAIL.n201 8.92171
R1919 VTAIL.n151 VTAIL.n150 8.92171
R1920 VTAIL.n135 VTAIL.n111 8.92171
R1921 VTAIL.n318 VTAIL.n317 8.14595
R1922 VTAIL.n326 VTAIL.n284 8.14595
R1923 VTAIL.n48 VTAIL.n47 8.14595
R1924 VTAIL.n56 VTAIL.n14 8.14595
R1925 VTAIL.n237 VTAIL.n195 8.14595
R1926 VTAIL.n229 VTAIL.n228 8.14595
R1927 VTAIL.n147 VTAIL.n105 8.14595
R1928 VTAIL.n139 VTAIL.n138 8.14595
R1929 VTAIL.n321 VTAIL.n288 7.3702
R1930 VTAIL.n325 VTAIL.n286 7.3702
R1931 VTAIL.n51 VTAIL.n18 7.3702
R1932 VTAIL.n55 VTAIL.n16 7.3702
R1933 VTAIL.n236 VTAIL.n197 7.3702
R1934 VTAIL.n232 VTAIL.n199 7.3702
R1935 VTAIL.n146 VTAIL.n107 7.3702
R1936 VTAIL.n142 VTAIL.n109 7.3702
R1937 VTAIL.n322 VTAIL.n321 6.59444
R1938 VTAIL.n322 VTAIL.n286 6.59444
R1939 VTAIL.n52 VTAIL.n51 6.59444
R1940 VTAIL.n52 VTAIL.n16 6.59444
R1941 VTAIL.n233 VTAIL.n197 6.59444
R1942 VTAIL.n233 VTAIL.n232 6.59444
R1943 VTAIL.n143 VTAIL.n107 6.59444
R1944 VTAIL.n143 VTAIL.n142 6.59444
R1945 VTAIL.n318 VTAIL.n288 5.81868
R1946 VTAIL.n326 VTAIL.n325 5.81868
R1947 VTAIL.n48 VTAIL.n18 5.81868
R1948 VTAIL.n56 VTAIL.n55 5.81868
R1949 VTAIL.n237 VTAIL.n236 5.81868
R1950 VTAIL.n229 VTAIL.n199 5.81868
R1951 VTAIL.n147 VTAIL.n146 5.81868
R1952 VTAIL.n139 VTAIL.n109 5.81868
R1953 VTAIL.n317 VTAIL.n290 5.04292
R1954 VTAIL.n329 VTAIL.n284 5.04292
R1955 VTAIL.n47 VTAIL.n20 5.04292
R1956 VTAIL.n59 VTAIL.n14 5.04292
R1957 VTAIL.n240 VTAIL.n195 5.04292
R1958 VTAIL.n228 VTAIL.n201 5.04292
R1959 VTAIL.n150 VTAIL.n105 5.04292
R1960 VTAIL.n138 VTAIL.n111 5.04292
R1961 VTAIL.n300 VTAIL.n299 4.38563
R1962 VTAIL.n30 VTAIL.n29 4.38563
R1963 VTAIL.n211 VTAIL.n210 4.38563
R1964 VTAIL.n121 VTAIL.n120 4.38563
R1965 VTAIL.n314 VTAIL.n313 4.26717
R1966 VTAIL.n330 VTAIL.n282 4.26717
R1967 VTAIL.n44 VTAIL.n43 4.26717
R1968 VTAIL.n60 VTAIL.n12 4.26717
R1969 VTAIL.n241 VTAIL.n193 4.26717
R1970 VTAIL.n225 VTAIL.n224 4.26717
R1971 VTAIL.n151 VTAIL.n103 4.26717
R1972 VTAIL.n135 VTAIL.n134 4.26717
R1973 VTAIL.n310 VTAIL.n292 3.49141
R1974 VTAIL.n334 VTAIL.n333 3.49141
R1975 VTAIL.n358 VTAIL.n270 3.49141
R1976 VTAIL.n40 VTAIL.n22 3.49141
R1977 VTAIL.n64 VTAIL.n63 3.49141
R1978 VTAIL.n88 VTAIL.n0 3.49141
R1979 VTAIL.n268 VTAIL.n180 3.49141
R1980 VTAIL.n245 VTAIL.n244 3.49141
R1981 VTAIL.n221 VTAIL.n203 3.49141
R1982 VTAIL.n178 VTAIL.n90 3.49141
R1983 VTAIL.n155 VTAIL.n154 3.49141
R1984 VTAIL.n131 VTAIL.n113 3.49141
R1985 VTAIL.n309 VTAIL.n294 2.71565
R1986 VTAIL.n337 VTAIL.n280 2.71565
R1987 VTAIL.n356 VTAIL.n355 2.71565
R1988 VTAIL.n39 VTAIL.n24 2.71565
R1989 VTAIL.n67 VTAIL.n10 2.71565
R1990 VTAIL.n86 VTAIL.n85 2.71565
R1991 VTAIL.n266 VTAIL.n265 2.71565
R1992 VTAIL.n248 VTAIL.n191 2.71565
R1993 VTAIL.n220 VTAIL.n205 2.71565
R1994 VTAIL.n176 VTAIL.n175 2.71565
R1995 VTAIL.n158 VTAIL.n101 2.71565
R1996 VTAIL.n130 VTAIL.n115 2.71565
R1997 VTAIL.n269 VTAIL.n179 2.29791
R1998 VTAIL.n306 VTAIL.n305 1.93989
R1999 VTAIL.n338 VTAIL.n278 1.93989
R2000 VTAIL.n352 VTAIL.n272 1.93989
R2001 VTAIL.n36 VTAIL.n35 1.93989
R2002 VTAIL.n68 VTAIL.n8 1.93989
R2003 VTAIL.n82 VTAIL.n2 1.93989
R2004 VTAIL.n262 VTAIL.n182 1.93989
R2005 VTAIL.n249 VTAIL.n189 1.93989
R2006 VTAIL.n217 VTAIL.n216 1.93989
R2007 VTAIL.n172 VTAIL.n92 1.93989
R2008 VTAIL.n159 VTAIL.n99 1.93989
R2009 VTAIL.n127 VTAIL.n126 1.93989
R2010 VTAIL VTAIL.n89 1.44231
R2011 VTAIL.n302 VTAIL.n296 1.16414
R2012 VTAIL.n343 VTAIL.n341 1.16414
R2013 VTAIL.n351 VTAIL.n274 1.16414
R2014 VTAIL.n32 VTAIL.n26 1.16414
R2015 VTAIL.n73 VTAIL.n71 1.16414
R2016 VTAIL.n81 VTAIL.n4 1.16414
R2017 VTAIL.n261 VTAIL.n184 1.16414
R2018 VTAIL.n253 VTAIL.n252 1.16414
R2019 VTAIL.n213 VTAIL.n207 1.16414
R2020 VTAIL.n171 VTAIL.n94 1.16414
R2021 VTAIL.n163 VTAIL.n162 1.16414
R2022 VTAIL.n123 VTAIL.n117 1.16414
R2023 VTAIL VTAIL.n359 0.856103
R2024 VTAIL.n301 VTAIL.n298 0.388379
R2025 VTAIL.n342 VTAIL.n276 0.388379
R2026 VTAIL.n348 VTAIL.n347 0.388379
R2027 VTAIL.n31 VTAIL.n28 0.388379
R2028 VTAIL.n72 VTAIL.n6 0.388379
R2029 VTAIL.n78 VTAIL.n77 0.388379
R2030 VTAIL.n258 VTAIL.n257 0.388379
R2031 VTAIL.n188 VTAIL.n186 0.388379
R2032 VTAIL.n212 VTAIL.n209 0.388379
R2033 VTAIL.n168 VTAIL.n167 0.388379
R2034 VTAIL.n98 VTAIL.n96 0.388379
R2035 VTAIL.n122 VTAIL.n119 0.388379
R2036 VTAIL.n300 VTAIL.n295 0.155672
R2037 VTAIL.n307 VTAIL.n295 0.155672
R2038 VTAIL.n308 VTAIL.n307 0.155672
R2039 VTAIL.n308 VTAIL.n291 0.155672
R2040 VTAIL.n315 VTAIL.n291 0.155672
R2041 VTAIL.n316 VTAIL.n315 0.155672
R2042 VTAIL.n316 VTAIL.n287 0.155672
R2043 VTAIL.n323 VTAIL.n287 0.155672
R2044 VTAIL.n324 VTAIL.n323 0.155672
R2045 VTAIL.n324 VTAIL.n283 0.155672
R2046 VTAIL.n331 VTAIL.n283 0.155672
R2047 VTAIL.n332 VTAIL.n331 0.155672
R2048 VTAIL.n332 VTAIL.n279 0.155672
R2049 VTAIL.n339 VTAIL.n279 0.155672
R2050 VTAIL.n340 VTAIL.n339 0.155672
R2051 VTAIL.n340 VTAIL.n275 0.155672
R2052 VTAIL.n349 VTAIL.n275 0.155672
R2053 VTAIL.n350 VTAIL.n349 0.155672
R2054 VTAIL.n350 VTAIL.n271 0.155672
R2055 VTAIL.n357 VTAIL.n271 0.155672
R2056 VTAIL.n30 VTAIL.n25 0.155672
R2057 VTAIL.n37 VTAIL.n25 0.155672
R2058 VTAIL.n38 VTAIL.n37 0.155672
R2059 VTAIL.n38 VTAIL.n21 0.155672
R2060 VTAIL.n45 VTAIL.n21 0.155672
R2061 VTAIL.n46 VTAIL.n45 0.155672
R2062 VTAIL.n46 VTAIL.n17 0.155672
R2063 VTAIL.n53 VTAIL.n17 0.155672
R2064 VTAIL.n54 VTAIL.n53 0.155672
R2065 VTAIL.n54 VTAIL.n13 0.155672
R2066 VTAIL.n61 VTAIL.n13 0.155672
R2067 VTAIL.n62 VTAIL.n61 0.155672
R2068 VTAIL.n62 VTAIL.n9 0.155672
R2069 VTAIL.n69 VTAIL.n9 0.155672
R2070 VTAIL.n70 VTAIL.n69 0.155672
R2071 VTAIL.n70 VTAIL.n5 0.155672
R2072 VTAIL.n79 VTAIL.n5 0.155672
R2073 VTAIL.n80 VTAIL.n79 0.155672
R2074 VTAIL.n80 VTAIL.n1 0.155672
R2075 VTAIL.n87 VTAIL.n1 0.155672
R2076 VTAIL.n267 VTAIL.n181 0.155672
R2077 VTAIL.n260 VTAIL.n181 0.155672
R2078 VTAIL.n260 VTAIL.n259 0.155672
R2079 VTAIL.n259 VTAIL.n185 0.155672
R2080 VTAIL.n251 VTAIL.n185 0.155672
R2081 VTAIL.n251 VTAIL.n250 0.155672
R2082 VTAIL.n250 VTAIL.n190 0.155672
R2083 VTAIL.n243 VTAIL.n190 0.155672
R2084 VTAIL.n243 VTAIL.n242 0.155672
R2085 VTAIL.n242 VTAIL.n194 0.155672
R2086 VTAIL.n235 VTAIL.n194 0.155672
R2087 VTAIL.n235 VTAIL.n234 0.155672
R2088 VTAIL.n234 VTAIL.n198 0.155672
R2089 VTAIL.n227 VTAIL.n198 0.155672
R2090 VTAIL.n227 VTAIL.n226 0.155672
R2091 VTAIL.n226 VTAIL.n202 0.155672
R2092 VTAIL.n219 VTAIL.n202 0.155672
R2093 VTAIL.n219 VTAIL.n218 0.155672
R2094 VTAIL.n218 VTAIL.n206 0.155672
R2095 VTAIL.n211 VTAIL.n206 0.155672
R2096 VTAIL.n177 VTAIL.n91 0.155672
R2097 VTAIL.n170 VTAIL.n91 0.155672
R2098 VTAIL.n170 VTAIL.n169 0.155672
R2099 VTAIL.n169 VTAIL.n95 0.155672
R2100 VTAIL.n161 VTAIL.n95 0.155672
R2101 VTAIL.n161 VTAIL.n160 0.155672
R2102 VTAIL.n160 VTAIL.n100 0.155672
R2103 VTAIL.n153 VTAIL.n100 0.155672
R2104 VTAIL.n153 VTAIL.n152 0.155672
R2105 VTAIL.n152 VTAIL.n104 0.155672
R2106 VTAIL.n145 VTAIL.n104 0.155672
R2107 VTAIL.n145 VTAIL.n144 0.155672
R2108 VTAIL.n144 VTAIL.n108 0.155672
R2109 VTAIL.n137 VTAIL.n108 0.155672
R2110 VTAIL.n137 VTAIL.n136 0.155672
R2111 VTAIL.n136 VTAIL.n112 0.155672
R2112 VTAIL.n129 VTAIL.n112 0.155672
R2113 VTAIL.n129 VTAIL.n128 0.155672
R2114 VTAIL.n128 VTAIL.n116 0.155672
R2115 VTAIL.n121 VTAIL.n116 0.155672
R2116 VDD2.n173 VDD2.n89 289.615
R2117 VDD2.n84 VDD2.n0 289.615
R2118 VDD2.n174 VDD2.n173 185
R2119 VDD2.n172 VDD2.n171 185
R2120 VDD2.n93 VDD2.n92 185
R2121 VDD2.n166 VDD2.n165 185
R2122 VDD2.n164 VDD2.n95 185
R2123 VDD2.n163 VDD2.n162 185
R2124 VDD2.n98 VDD2.n96 185
R2125 VDD2.n157 VDD2.n156 185
R2126 VDD2.n155 VDD2.n154 185
R2127 VDD2.n102 VDD2.n101 185
R2128 VDD2.n149 VDD2.n148 185
R2129 VDD2.n147 VDD2.n146 185
R2130 VDD2.n106 VDD2.n105 185
R2131 VDD2.n141 VDD2.n140 185
R2132 VDD2.n139 VDD2.n138 185
R2133 VDD2.n110 VDD2.n109 185
R2134 VDD2.n133 VDD2.n132 185
R2135 VDD2.n131 VDD2.n130 185
R2136 VDD2.n114 VDD2.n113 185
R2137 VDD2.n125 VDD2.n124 185
R2138 VDD2.n123 VDD2.n122 185
R2139 VDD2.n118 VDD2.n117 185
R2140 VDD2.n28 VDD2.n27 185
R2141 VDD2.n33 VDD2.n32 185
R2142 VDD2.n35 VDD2.n34 185
R2143 VDD2.n24 VDD2.n23 185
R2144 VDD2.n41 VDD2.n40 185
R2145 VDD2.n43 VDD2.n42 185
R2146 VDD2.n20 VDD2.n19 185
R2147 VDD2.n49 VDD2.n48 185
R2148 VDD2.n51 VDD2.n50 185
R2149 VDD2.n16 VDD2.n15 185
R2150 VDD2.n57 VDD2.n56 185
R2151 VDD2.n59 VDD2.n58 185
R2152 VDD2.n12 VDD2.n11 185
R2153 VDD2.n65 VDD2.n64 185
R2154 VDD2.n67 VDD2.n66 185
R2155 VDD2.n8 VDD2.n7 185
R2156 VDD2.n74 VDD2.n73 185
R2157 VDD2.n75 VDD2.n6 185
R2158 VDD2.n77 VDD2.n76 185
R2159 VDD2.n4 VDD2.n3 185
R2160 VDD2.n83 VDD2.n82 185
R2161 VDD2.n85 VDD2.n84 185
R2162 VDD2.n119 VDD2.t0 147.659
R2163 VDD2.n29 VDD2.t1 147.659
R2164 VDD2.n173 VDD2.n172 104.615
R2165 VDD2.n172 VDD2.n92 104.615
R2166 VDD2.n165 VDD2.n92 104.615
R2167 VDD2.n165 VDD2.n164 104.615
R2168 VDD2.n164 VDD2.n163 104.615
R2169 VDD2.n163 VDD2.n96 104.615
R2170 VDD2.n156 VDD2.n96 104.615
R2171 VDD2.n156 VDD2.n155 104.615
R2172 VDD2.n155 VDD2.n101 104.615
R2173 VDD2.n148 VDD2.n101 104.615
R2174 VDD2.n148 VDD2.n147 104.615
R2175 VDD2.n147 VDD2.n105 104.615
R2176 VDD2.n140 VDD2.n105 104.615
R2177 VDD2.n140 VDD2.n139 104.615
R2178 VDD2.n139 VDD2.n109 104.615
R2179 VDD2.n132 VDD2.n109 104.615
R2180 VDD2.n132 VDD2.n131 104.615
R2181 VDD2.n131 VDD2.n113 104.615
R2182 VDD2.n124 VDD2.n113 104.615
R2183 VDD2.n124 VDD2.n123 104.615
R2184 VDD2.n123 VDD2.n117 104.615
R2185 VDD2.n33 VDD2.n27 104.615
R2186 VDD2.n34 VDD2.n33 104.615
R2187 VDD2.n34 VDD2.n23 104.615
R2188 VDD2.n41 VDD2.n23 104.615
R2189 VDD2.n42 VDD2.n41 104.615
R2190 VDD2.n42 VDD2.n19 104.615
R2191 VDD2.n49 VDD2.n19 104.615
R2192 VDD2.n50 VDD2.n49 104.615
R2193 VDD2.n50 VDD2.n15 104.615
R2194 VDD2.n57 VDD2.n15 104.615
R2195 VDD2.n58 VDD2.n57 104.615
R2196 VDD2.n58 VDD2.n11 104.615
R2197 VDD2.n65 VDD2.n11 104.615
R2198 VDD2.n66 VDD2.n65 104.615
R2199 VDD2.n66 VDD2.n7 104.615
R2200 VDD2.n74 VDD2.n7 104.615
R2201 VDD2.n75 VDD2.n74 104.615
R2202 VDD2.n76 VDD2.n75 104.615
R2203 VDD2.n76 VDD2.n3 104.615
R2204 VDD2.n83 VDD2.n3 104.615
R2205 VDD2.n84 VDD2.n83 104.615
R2206 VDD2.n178 VDD2.n88 93.0883
R2207 VDD2.t0 VDD2.n117 52.3082
R2208 VDD2.t1 VDD2.n27 52.3082
R2209 VDD2.n178 VDD2.n177 48.2823
R2210 VDD2.n119 VDD2.n118 15.6677
R2211 VDD2.n29 VDD2.n28 15.6677
R2212 VDD2.n166 VDD2.n95 13.1884
R2213 VDD2.n77 VDD2.n6 13.1884
R2214 VDD2.n167 VDD2.n93 12.8005
R2215 VDD2.n162 VDD2.n97 12.8005
R2216 VDD2.n122 VDD2.n121 12.8005
R2217 VDD2.n32 VDD2.n31 12.8005
R2218 VDD2.n73 VDD2.n72 12.8005
R2219 VDD2.n78 VDD2.n4 12.8005
R2220 VDD2.n171 VDD2.n170 12.0247
R2221 VDD2.n161 VDD2.n98 12.0247
R2222 VDD2.n125 VDD2.n116 12.0247
R2223 VDD2.n35 VDD2.n26 12.0247
R2224 VDD2.n71 VDD2.n8 12.0247
R2225 VDD2.n82 VDD2.n81 12.0247
R2226 VDD2.n174 VDD2.n91 11.249
R2227 VDD2.n158 VDD2.n157 11.249
R2228 VDD2.n126 VDD2.n114 11.249
R2229 VDD2.n36 VDD2.n24 11.249
R2230 VDD2.n68 VDD2.n67 11.249
R2231 VDD2.n85 VDD2.n2 11.249
R2232 VDD2.n175 VDD2.n89 10.4732
R2233 VDD2.n154 VDD2.n100 10.4732
R2234 VDD2.n130 VDD2.n129 10.4732
R2235 VDD2.n40 VDD2.n39 10.4732
R2236 VDD2.n64 VDD2.n10 10.4732
R2237 VDD2.n86 VDD2.n0 10.4732
R2238 VDD2.n153 VDD2.n102 9.69747
R2239 VDD2.n133 VDD2.n112 9.69747
R2240 VDD2.n43 VDD2.n22 9.69747
R2241 VDD2.n63 VDD2.n12 9.69747
R2242 VDD2.n177 VDD2.n176 9.45567
R2243 VDD2.n88 VDD2.n87 9.45567
R2244 VDD2.n145 VDD2.n144 9.3005
R2245 VDD2.n104 VDD2.n103 9.3005
R2246 VDD2.n151 VDD2.n150 9.3005
R2247 VDD2.n153 VDD2.n152 9.3005
R2248 VDD2.n100 VDD2.n99 9.3005
R2249 VDD2.n159 VDD2.n158 9.3005
R2250 VDD2.n161 VDD2.n160 9.3005
R2251 VDD2.n97 VDD2.n94 9.3005
R2252 VDD2.n176 VDD2.n175 9.3005
R2253 VDD2.n91 VDD2.n90 9.3005
R2254 VDD2.n170 VDD2.n169 9.3005
R2255 VDD2.n168 VDD2.n167 9.3005
R2256 VDD2.n143 VDD2.n142 9.3005
R2257 VDD2.n108 VDD2.n107 9.3005
R2258 VDD2.n137 VDD2.n136 9.3005
R2259 VDD2.n135 VDD2.n134 9.3005
R2260 VDD2.n112 VDD2.n111 9.3005
R2261 VDD2.n129 VDD2.n128 9.3005
R2262 VDD2.n127 VDD2.n126 9.3005
R2263 VDD2.n116 VDD2.n115 9.3005
R2264 VDD2.n121 VDD2.n120 9.3005
R2265 VDD2.n87 VDD2.n86 9.3005
R2266 VDD2.n2 VDD2.n1 9.3005
R2267 VDD2.n81 VDD2.n80 9.3005
R2268 VDD2.n79 VDD2.n78 9.3005
R2269 VDD2.n18 VDD2.n17 9.3005
R2270 VDD2.n47 VDD2.n46 9.3005
R2271 VDD2.n45 VDD2.n44 9.3005
R2272 VDD2.n22 VDD2.n21 9.3005
R2273 VDD2.n39 VDD2.n38 9.3005
R2274 VDD2.n37 VDD2.n36 9.3005
R2275 VDD2.n26 VDD2.n25 9.3005
R2276 VDD2.n31 VDD2.n30 9.3005
R2277 VDD2.n53 VDD2.n52 9.3005
R2278 VDD2.n55 VDD2.n54 9.3005
R2279 VDD2.n14 VDD2.n13 9.3005
R2280 VDD2.n61 VDD2.n60 9.3005
R2281 VDD2.n63 VDD2.n62 9.3005
R2282 VDD2.n10 VDD2.n9 9.3005
R2283 VDD2.n69 VDD2.n68 9.3005
R2284 VDD2.n71 VDD2.n70 9.3005
R2285 VDD2.n72 VDD2.n5 9.3005
R2286 VDD2.n150 VDD2.n149 8.92171
R2287 VDD2.n134 VDD2.n110 8.92171
R2288 VDD2.n44 VDD2.n20 8.92171
R2289 VDD2.n60 VDD2.n59 8.92171
R2290 VDD2.n146 VDD2.n104 8.14595
R2291 VDD2.n138 VDD2.n137 8.14595
R2292 VDD2.n48 VDD2.n47 8.14595
R2293 VDD2.n56 VDD2.n14 8.14595
R2294 VDD2.n145 VDD2.n106 7.3702
R2295 VDD2.n141 VDD2.n108 7.3702
R2296 VDD2.n51 VDD2.n18 7.3702
R2297 VDD2.n55 VDD2.n16 7.3702
R2298 VDD2.n142 VDD2.n106 6.59444
R2299 VDD2.n142 VDD2.n141 6.59444
R2300 VDD2.n52 VDD2.n51 6.59444
R2301 VDD2.n52 VDD2.n16 6.59444
R2302 VDD2.n146 VDD2.n145 5.81868
R2303 VDD2.n138 VDD2.n108 5.81868
R2304 VDD2.n48 VDD2.n18 5.81868
R2305 VDD2.n56 VDD2.n55 5.81868
R2306 VDD2.n149 VDD2.n104 5.04292
R2307 VDD2.n137 VDD2.n110 5.04292
R2308 VDD2.n47 VDD2.n20 5.04292
R2309 VDD2.n59 VDD2.n14 5.04292
R2310 VDD2.n120 VDD2.n119 4.38563
R2311 VDD2.n30 VDD2.n29 4.38563
R2312 VDD2.n150 VDD2.n102 4.26717
R2313 VDD2.n134 VDD2.n133 4.26717
R2314 VDD2.n44 VDD2.n43 4.26717
R2315 VDD2.n60 VDD2.n12 4.26717
R2316 VDD2.n177 VDD2.n89 3.49141
R2317 VDD2.n154 VDD2.n153 3.49141
R2318 VDD2.n130 VDD2.n112 3.49141
R2319 VDD2.n40 VDD2.n22 3.49141
R2320 VDD2.n64 VDD2.n63 3.49141
R2321 VDD2.n88 VDD2.n0 3.49141
R2322 VDD2.n175 VDD2.n174 2.71565
R2323 VDD2.n157 VDD2.n100 2.71565
R2324 VDD2.n129 VDD2.n114 2.71565
R2325 VDD2.n39 VDD2.n24 2.71565
R2326 VDD2.n67 VDD2.n10 2.71565
R2327 VDD2.n86 VDD2.n85 2.71565
R2328 VDD2.n171 VDD2.n91 1.93989
R2329 VDD2.n158 VDD2.n98 1.93989
R2330 VDD2.n126 VDD2.n125 1.93989
R2331 VDD2.n36 VDD2.n35 1.93989
R2332 VDD2.n68 VDD2.n8 1.93989
R2333 VDD2.n82 VDD2.n2 1.93989
R2334 VDD2.n170 VDD2.n93 1.16414
R2335 VDD2.n162 VDD2.n161 1.16414
R2336 VDD2.n122 VDD2.n116 1.16414
R2337 VDD2.n32 VDD2.n26 1.16414
R2338 VDD2.n73 VDD2.n71 1.16414
R2339 VDD2.n81 VDD2.n4 1.16414
R2340 VDD2 VDD2.n178 0.972483
R2341 VDD2.n167 VDD2.n166 0.388379
R2342 VDD2.n97 VDD2.n95 0.388379
R2343 VDD2.n121 VDD2.n118 0.388379
R2344 VDD2.n31 VDD2.n28 0.388379
R2345 VDD2.n72 VDD2.n6 0.388379
R2346 VDD2.n78 VDD2.n77 0.388379
R2347 VDD2.n176 VDD2.n90 0.155672
R2348 VDD2.n169 VDD2.n90 0.155672
R2349 VDD2.n169 VDD2.n168 0.155672
R2350 VDD2.n168 VDD2.n94 0.155672
R2351 VDD2.n160 VDD2.n94 0.155672
R2352 VDD2.n160 VDD2.n159 0.155672
R2353 VDD2.n159 VDD2.n99 0.155672
R2354 VDD2.n152 VDD2.n99 0.155672
R2355 VDD2.n152 VDD2.n151 0.155672
R2356 VDD2.n151 VDD2.n103 0.155672
R2357 VDD2.n144 VDD2.n103 0.155672
R2358 VDD2.n144 VDD2.n143 0.155672
R2359 VDD2.n143 VDD2.n107 0.155672
R2360 VDD2.n136 VDD2.n107 0.155672
R2361 VDD2.n136 VDD2.n135 0.155672
R2362 VDD2.n135 VDD2.n111 0.155672
R2363 VDD2.n128 VDD2.n111 0.155672
R2364 VDD2.n128 VDD2.n127 0.155672
R2365 VDD2.n127 VDD2.n115 0.155672
R2366 VDD2.n120 VDD2.n115 0.155672
R2367 VDD2.n30 VDD2.n25 0.155672
R2368 VDD2.n37 VDD2.n25 0.155672
R2369 VDD2.n38 VDD2.n37 0.155672
R2370 VDD2.n38 VDD2.n21 0.155672
R2371 VDD2.n45 VDD2.n21 0.155672
R2372 VDD2.n46 VDD2.n45 0.155672
R2373 VDD2.n46 VDD2.n17 0.155672
R2374 VDD2.n53 VDD2.n17 0.155672
R2375 VDD2.n54 VDD2.n53 0.155672
R2376 VDD2.n54 VDD2.n13 0.155672
R2377 VDD2.n61 VDD2.n13 0.155672
R2378 VDD2.n62 VDD2.n61 0.155672
R2379 VDD2.n62 VDD2.n9 0.155672
R2380 VDD2.n69 VDD2.n9 0.155672
R2381 VDD2.n70 VDD2.n69 0.155672
R2382 VDD2.n70 VDD2.n5 0.155672
R2383 VDD2.n79 VDD2.n5 0.155672
R2384 VDD2.n80 VDD2.n79 0.155672
R2385 VDD2.n80 VDD2.n1 0.155672
R2386 VDD2.n87 VDD2.n1 0.155672
R2387 VP.n0 VP.t1 185.163
R2388 VP.n0 VP.t0 133.964
R2389 VP VP.n0 0.621237
R2390 VDD1.n84 VDD1.n0 289.615
R2391 VDD1.n173 VDD1.n89 289.615
R2392 VDD1.n85 VDD1.n84 185
R2393 VDD1.n83 VDD1.n82 185
R2394 VDD1.n4 VDD1.n3 185
R2395 VDD1.n77 VDD1.n76 185
R2396 VDD1.n75 VDD1.n6 185
R2397 VDD1.n74 VDD1.n73 185
R2398 VDD1.n9 VDD1.n7 185
R2399 VDD1.n68 VDD1.n67 185
R2400 VDD1.n66 VDD1.n65 185
R2401 VDD1.n13 VDD1.n12 185
R2402 VDD1.n60 VDD1.n59 185
R2403 VDD1.n58 VDD1.n57 185
R2404 VDD1.n17 VDD1.n16 185
R2405 VDD1.n52 VDD1.n51 185
R2406 VDD1.n50 VDD1.n49 185
R2407 VDD1.n21 VDD1.n20 185
R2408 VDD1.n44 VDD1.n43 185
R2409 VDD1.n42 VDD1.n41 185
R2410 VDD1.n25 VDD1.n24 185
R2411 VDD1.n36 VDD1.n35 185
R2412 VDD1.n34 VDD1.n33 185
R2413 VDD1.n29 VDD1.n28 185
R2414 VDD1.n117 VDD1.n116 185
R2415 VDD1.n122 VDD1.n121 185
R2416 VDD1.n124 VDD1.n123 185
R2417 VDD1.n113 VDD1.n112 185
R2418 VDD1.n130 VDD1.n129 185
R2419 VDD1.n132 VDD1.n131 185
R2420 VDD1.n109 VDD1.n108 185
R2421 VDD1.n138 VDD1.n137 185
R2422 VDD1.n140 VDD1.n139 185
R2423 VDD1.n105 VDD1.n104 185
R2424 VDD1.n146 VDD1.n145 185
R2425 VDD1.n148 VDD1.n147 185
R2426 VDD1.n101 VDD1.n100 185
R2427 VDD1.n154 VDD1.n153 185
R2428 VDD1.n156 VDD1.n155 185
R2429 VDD1.n97 VDD1.n96 185
R2430 VDD1.n163 VDD1.n162 185
R2431 VDD1.n164 VDD1.n95 185
R2432 VDD1.n166 VDD1.n165 185
R2433 VDD1.n93 VDD1.n92 185
R2434 VDD1.n172 VDD1.n171 185
R2435 VDD1.n174 VDD1.n173 185
R2436 VDD1.n30 VDD1.t0 147.659
R2437 VDD1.n118 VDD1.t1 147.659
R2438 VDD1.n84 VDD1.n83 104.615
R2439 VDD1.n83 VDD1.n3 104.615
R2440 VDD1.n76 VDD1.n3 104.615
R2441 VDD1.n76 VDD1.n75 104.615
R2442 VDD1.n75 VDD1.n74 104.615
R2443 VDD1.n74 VDD1.n7 104.615
R2444 VDD1.n67 VDD1.n7 104.615
R2445 VDD1.n67 VDD1.n66 104.615
R2446 VDD1.n66 VDD1.n12 104.615
R2447 VDD1.n59 VDD1.n12 104.615
R2448 VDD1.n59 VDD1.n58 104.615
R2449 VDD1.n58 VDD1.n16 104.615
R2450 VDD1.n51 VDD1.n16 104.615
R2451 VDD1.n51 VDD1.n50 104.615
R2452 VDD1.n50 VDD1.n20 104.615
R2453 VDD1.n43 VDD1.n20 104.615
R2454 VDD1.n43 VDD1.n42 104.615
R2455 VDD1.n42 VDD1.n24 104.615
R2456 VDD1.n35 VDD1.n24 104.615
R2457 VDD1.n35 VDD1.n34 104.615
R2458 VDD1.n34 VDD1.n28 104.615
R2459 VDD1.n122 VDD1.n116 104.615
R2460 VDD1.n123 VDD1.n122 104.615
R2461 VDD1.n123 VDD1.n112 104.615
R2462 VDD1.n130 VDD1.n112 104.615
R2463 VDD1.n131 VDD1.n130 104.615
R2464 VDD1.n131 VDD1.n108 104.615
R2465 VDD1.n138 VDD1.n108 104.615
R2466 VDD1.n139 VDD1.n138 104.615
R2467 VDD1.n139 VDD1.n104 104.615
R2468 VDD1.n146 VDD1.n104 104.615
R2469 VDD1.n147 VDD1.n146 104.615
R2470 VDD1.n147 VDD1.n100 104.615
R2471 VDD1.n154 VDD1.n100 104.615
R2472 VDD1.n155 VDD1.n154 104.615
R2473 VDD1.n155 VDD1.n96 104.615
R2474 VDD1.n163 VDD1.n96 104.615
R2475 VDD1.n164 VDD1.n163 104.615
R2476 VDD1.n165 VDD1.n164 104.615
R2477 VDD1.n165 VDD1.n92 104.615
R2478 VDD1.n172 VDD1.n92 104.615
R2479 VDD1.n173 VDD1.n172 104.615
R2480 VDD1 VDD1.n177 94.5269
R2481 VDD1.t0 VDD1.n28 52.3082
R2482 VDD1.t1 VDD1.n116 52.3082
R2483 VDD1 VDD1.n88 49.2543
R2484 VDD1.n30 VDD1.n29 15.6677
R2485 VDD1.n118 VDD1.n117 15.6677
R2486 VDD1.n77 VDD1.n6 13.1884
R2487 VDD1.n166 VDD1.n95 13.1884
R2488 VDD1.n78 VDD1.n4 12.8005
R2489 VDD1.n73 VDD1.n8 12.8005
R2490 VDD1.n33 VDD1.n32 12.8005
R2491 VDD1.n121 VDD1.n120 12.8005
R2492 VDD1.n162 VDD1.n161 12.8005
R2493 VDD1.n167 VDD1.n93 12.8005
R2494 VDD1.n82 VDD1.n81 12.0247
R2495 VDD1.n72 VDD1.n9 12.0247
R2496 VDD1.n36 VDD1.n27 12.0247
R2497 VDD1.n124 VDD1.n115 12.0247
R2498 VDD1.n160 VDD1.n97 12.0247
R2499 VDD1.n171 VDD1.n170 12.0247
R2500 VDD1.n85 VDD1.n2 11.249
R2501 VDD1.n69 VDD1.n68 11.249
R2502 VDD1.n37 VDD1.n25 11.249
R2503 VDD1.n125 VDD1.n113 11.249
R2504 VDD1.n157 VDD1.n156 11.249
R2505 VDD1.n174 VDD1.n91 11.249
R2506 VDD1.n86 VDD1.n0 10.4732
R2507 VDD1.n65 VDD1.n11 10.4732
R2508 VDD1.n41 VDD1.n40 10.4732
R2509 VDD1.n129 VDD1.n128 10.4732
R2510 VDD1.n153 VDD1.n99 10.4732
R2511 VDD1.n175 VDD1.n89 10.4732
R2512 VDD1.n64 VDD1.n13 9.69747
R2513 VDD1.n44 VDD1.n23 9.69747
R2514 VDD1.n132 VDD1.n111 9.69747
R2515 VDD1.n152 VDD1.n101 9.69747
R2516 VDD1.n88 VDD1.n87 9.45567
R2517 VDD1.n177 VDD1.n176 9.45567
R2518 VDD1.n56 VDD1.n55 9.3005
R2519 VDD1.n15 VDD1.n14 9.3005
R2520 VDD1.n62 VDD1.n61 9.3005
R2521 VDD1.n64 VDD1.n63 9.3005
R2522 VDD1.n11 VDD1.n10 9.3005
R2523 VDD1.n70 VDD1.n69 9.3005
R2524 VDD1.n72 VDD1.n71 9.3005
R2525 VDD1.n8 VDD1.n5 9.3005
R2526 VDD1.n87 VDD1.n86 9.3005
R2527 VDD1.n2 VDD1.n1 9.3005
R2528 VDD1.n81 VDD1.n80 9.3005
R2529 VDD1.n79 VDD1.n78 9.3005
R2530 VDD1.n54 VDD1.n53 9.3005
R2531 VDD1.n19 VDD1.n18 9.3005
R2532 VDD1.n48 VDD1.n47 9.3005
R2533 VDD1.n46 VDD1.n45 9.3005
R2534 VDD1.n23 VDD1.n22 9.3005
R2535 VDD1.n40 VDD1.n39 9.3005
R2536 VDD1.n38 VDD1.n37 9.3005
R2537 VDD1.n27 VDD1.n26 9.3005
R2538 VDD1.n32 VDD1.n31 9.3005
R2539 VDD1.n176 VDD1.n175 9.3005
R2540 VDD1.n91 VDD1.n90 9.3005
R2541 VDD1.n170 VDD1.n169 9.3005
R2542 VDD1.n168 VDD1.n167 9.3005
R2543 VDD1.n107 VDD1.n106 9.3005
R2544 VDD1.n136 VDD1.n135 9.3005
R2545 VDD1.n134 VDD1.n133 9.3005
R2546 VDD1.n111 VDD1.n110 9.3005
R2547 VDD1.n128 VDD1.n127 9.3005
R2548 VDD1.n126 VDD1.n125 9.3005
R2549 VDD1.n115 VDD1.n114 9.3005
R2550 VDD1.n120 VDD1.n119 9.3005
R2551 VDD1.n142 VDD1.n141 9.3005
R2552 VDD1.n144 VDD1.n143 9.3005
R2553 VDD1.n103 VDD1.n102 9.3005
R2554 VDD1.n150 VDD1.n149 9.3005
R2555 VDD1.n152 VDD1.n151 9.3005
R2556 VDD1.n99 VDD1.n98 9.3005
R2557 VDD1.n158 VDD1.n157 9.3005
R2558 VDD1.n160 VDD1.n159 9.3005
R2559 VDD1.n161 VDD1.n94 9.3005
R2560 VDD1.n61 VDD1.n60 8.92171
R2561 VDD1.n45 VDD1.n21 8.92171
R2562 VDD1.n133 VDD1.n109 8.92171
R2563 VDD1.n149 VDD1.n148 8.92171
R2564 VDD1.n57 VDD1.n15 8.14595
R2565 VDD1.n49 VDD1.n48 8.14595
R2566 VDD1.n137 VDD1.n136 8.14595
R2567 VDD1.n145 VDD1.n103 8.14595
R2568 VDD1.n56 VDD1.n17 7.3702
R2569 VDD1.n52 VDD1.n19 7.3702
R2570 VDD1.n140 VDD1.n107 7.3702
R2571 VDD1.n144 VDD1.n105 7.3702
R2572 VDD1.n53 VDD1.n17 6.59444
R2573 VDD1.n53 VDD1.n52 6.59444
R2574 VDD1.n141 VDD1.n140 6.59444
R2575 VDD1.n141 VDD1.n105 6.59444
R2576 VDD1.n57 VDD1.n56 5.81868
R2577 VDD1.n49 VDD1.n19 5.81868
R2578 VDD1.n137 VDD1.n107 5.81868
R2579 VDD1.n145 VDD1.n144 5.81868
R2580 VDD1.n60 VDD1.n15 5.04292
R2581 VDD1.n48 VDD1.n21 5.04292
R2582 VDD1.n136 VDD1.n109 5.04292
R2583 VDD1.n148 VDD1.n103 5.04292
R2584 VDD1.n31 VDD1.n30 4.38563
R2585 VDD1.n119 VDD1.n118 4.38563
R2586 VDD1.n61 VDD1.n13 4.26717
R2587 VDD1.n45 VDD1.n44 4.26717
R2588 VDD1.n133 VDD1.n132 4.26717
R2589 VDD1.n149 VDD1.n101 4.26717
R2590 VDD1.n88 VDD1.n0 3.49141
R2591 VDD1.n65 VDD1.n64 3.49141
R2592 VDD1.n41 VDD1.n23 3.49141
R2593 VDD1.n129 VDD1.n111 3.49141
R2594 VDD1.n153 VDD1.n152 3.49141
R2595 VDD1.n177 VDD1.n89 3.49141
R2596 VDD1.n86 VDD1.n85 2.71565
R2597 VDD1.n68 VDD1.n11 2.71565
R2598 VDD1.n40 VDD1.n25 2.71565
R2599 VDD1.n128 VDD1.n113 2.71565
R2600 VDD1.n156 VDD1.n99 2.71565
R2601 VDD1.n175 VDD1.n174 2.71565
R2602 VDD1.n82 VDD1.n2 1.93989
R2603 VDD1.n69 VDD1.n9 1.93989
R2604 VDD1.n37 VDD1.n36 1.93989
R2605 VDD1.n125 VDD1.n124 1.93989
R2606 VDD1.n157 VDD1.n97 1.93989
R2607 VDD1.n171 VDD1.n91 1.93989
R2608 VDD1.n81 VDD1.n4 1.16414
R2609 VDD1.n73 VDD1.n72 1.16414
R2610 VDD1.n33 VDD1.n27 1.16414
R2611 VDD1.n121 VDD1.n115 1.16414
R2612 VDD1.n162 VDD1.n160 1.16414
R2613 VDD1.n170 VDD1.n93 1.16414
R2614 VDD1.n78 VDD1.n77 0.388379
R2615 VDD1.n8 VDD1.n6 0.388379
R2616 VDD1.n32 VDD1.n29 0.388379
R2617 VDD1.n120 VDD1.n117 0.388379
R2618 VDD1.n161 VDD1.n95 0.388379
R2619 VDD1.n167 VDD1.n166 0.388379
R2620 VDD1.n87 VDD1.n1 0.155672
R2621 VDD1.n80 VDD1.n1 0.155672
R2622 VDD1.n80 VDD1.n79 0.155672
R2623 VDD1.n79 VDD1.n5 0.155672
R2624 VDD1.n71 VDD1.n5 0.155672
R2625 VDD1.n71 VDD1.n70 0.155672
R2626 VDD1.n70 VDD1.n10 0.155672
R2627 VDD1.n63 VDD1.n10 0.155672
R2628 VDD1.n63 VDD1.n62 0.155672
R2629 VDD1.n62 VDD1.n14 0.155672
R2630 VDD1.n55 VDD1.n14 0.155672
R2631 VDD1.n55 VDD1.n54 0.155672
R2632 VDD1.n54 VDD1.n18 0.155672
R2633 VDD1.n47 VDD1.n18 0.155672
R2634 VDD1.n47 VDD1.n46 0.155672
R2635 VDD1.n46 VDD1.n22 0.155672
R2636 VDD1.n39 VDD1.n22 0.155672
R2637 VDD1.n39 VDD1.n38 0.155672
R2638 VDD1.n38 VDD1.n26 0.155672
R2639 VDD1.n31 VDD1.n26 0.155672
R2640 VDD1.n119 VDD1.n114 0.155672
R2641 VDD1.n126 VDD1.n114 0.155672
R2642 VDD1.n127 VDD1.n126 0.155672
R2643 VDD1.n127 VDD1.n110 0.155672
R2644 VDD1.n134 VDD1.n110 0.155672
R2645 VDD1.n135 VDD1.n134 0.155672
R2646 VDD1.n135 VDD1.n106 0.155672
R2647 VDD1.n142 VDD1.n106 0.155672
R2648 VDD1.n143 VDD1.n142 0.155672
R2649 VDD1.n143 VDD1.n102 0.155672
R2650 VDD1.n150 VDD1.n102 0.155672
R2651 VDD1.n151 VDD1.n150 0.155672
R2652 VDD1.n151 VDD1.n98 0.155672
R2653 VDD1.n158 VDD1.n98 0.155672
R2654 VDD1.n159 VDD1.n158 0.155672
R2655 VDD1.n159 VDD1.n94 0.155672
R2656 VDD1.n168 VDD1.n94 0.155672
R2657 VDD1.n169 VDD1.n168 0.155672
R2658 VDD1.n169 VDD1.n90 0.155672
R2659 VDD1.n176 VDD1.n90 0.155672
C0 VP VN 6.82094f
C1 VP VTAIL 3.39827f
C2 VN VTAIL 3.38312f
C3 VDD2 VP 0.387456f
C4 VDD2 VN 3.83227f
C5 VDD2 VTAIL 6.40607f
C6 VDD1 VP 4.06936f
C7 VDD1 VN 0.148724f
C8 VDD1 VTAIL 6.34626f
C9 VDD1 VDD2 0.822234f
C10 VDD2 B 5.627538f
C11 VDD1 B 8.91048f
C12 VTAIL B 9.65037f
C13 VN B 12.935f
C14 VP B 8.294754f
C15 VDD1.n0 B 0.026559f
C16 VDD1.n1 B 0.020362f
C17 VDD1.n2 B 0.010941f
C18 VDD1.n3 B 0.025862f
C19 VDD1.n4 B 0.011585f
C20 VDD1.n5 B 0.020362f
C21 VDD1.n6 B 0.011263f
C22 VDD1.n7 B 0.025862f
C23 VDD1.n8 B 0.010941f
C24 VDD1.n9 B 0.011585f
C25 VDD1.n10 B 0.020362f
C26 VDD1.n11 B 0.010941f
C27 VDD1.n12 B 0.025862f
C28 VDD1.n13 B 0.011585f
C29 VDD1.n14 B 0.020362f
C30 VDD1.n15 B 0.010941f
C31 VDD1.n16 B 0.025862f
C32 VDD1.n17 B 0.011585f
C33 VDD1.n18 B 0.020362f
C34 VDD1.n19 B 0.010941f
C35 VDD1.n20 B 0.025862f
C36 VDD1.n21 B 0.011585f
C37 VDD1.n22 B 0.020362f
C38 VDD1.n23 B 0.010941f
C39 VDD1.n24 B 0.025862f
C40 VDD1.n25 B 0.011585f
C41 VDD1.n26 B 0.020362f
C42 VDD1.n27 B 0.010941f
C43 VDD1.n28 B 0.019396f
C44 VDD1.n29 B 0.015277f
C45 VDD1.t0 B 0.042716f
C46 VDD1.n30 B 0.138164f
C47 VDD1.n31 B 1.42274f
C48 VDD1.n32 B 0.010941f
C49 VDD1.n33 B 0.011585f
C50 VDD1.n34 B 0.025862f
C51 VDD1.n35 B 0.025862f
C52 VDD1.n36 B 0.011585f
C53 VDD1.n37 B 0.010941f
C54 VDD1.n38 B 0.020362f
C55 VDD1.n39 B 0.020362f
C56 VDD1.n40 B 0.010941f
C57 VDD1.n41 B 0.011585f
C58 VDD1.n42 B 0.025862f
C59 VDD1.n43 B 0.025862f
C60 VDD1.n44 B 0.011585f
C61 VDD1.n45 B 0.010941f
C62 VDD1.n46 B 0.020362f
C63 VDD1.n47 B 0.020362f
C64 VDD1.n48 B 0.010941f
C65 VDD1.n49 B 0.011585f
C66 VDD1.n50 B 0.025862f
C67 VDD1.n51 B 0.025862f
C68 VDD1.n52 B 0.011585f
C69 VDD1.n53 B 0.010941f
C70 VDD1.n54 B 0.020362f
C71 VDD1.n55 B 0.020362f
C72 VDD1.n56 B 0.010941f
C73 VDD1.n57 B 0.011585f
C74 VDD1.n58 B 0.025862f
C75 VDD1.n59 B 0.025862f
C76 VDD1.n60 B 0.011585f
C77 VDD1.n61 B 0.010941f
C78 VDD1.n62 B 0.020362f
C79 VDD1.n63 B 0.020362f
C80 VDD1.n64 B 0.010941f
C81 VDD1.n65 B 0.011585f
C82 VDD1.n66 B 0.025862f
C83 VDD1.n67 B 0.025862f
C84 VDD1.n68 B 0.011585f
C85 VDD1.n69 B 0.010941f
C86 VDD1.n70 B 0.020362f
C87 VDD1.n71 B 0.020362f
C88 VDD1.n72 B 0.010941f
C89 VDD1.n73 B 0.011585f
C90 VDD1.n74 B 0.025862f
C91 VDD1.n75 B 0.025862f
C92 VDD1.n76 B 0.025862f
C93 VDD1.n77 B 0.011263f
C94 VDD1.n78 B 0.010941f
C95 VDD1.n79 B 0.020362f
C96 VDD1.n80 B 0.020362f
C97 VDD1.n81 B 0.010941f
C98 VDD1.n82 B 0.011585f
C99 VDD1.n83 B 0.025862f
C100 VDD1.n84 B 0.052342f
C101 VDD1.n85 B 0.011585f
C102 VDD1.n86 B 0.010941f
C103 VDD1.n87 B 0.04623f
C104 VDD1.n88 B 0.044976f
C105 VDD1.n89 B 0.026559f
C106 VDD1.n90 B 0.020362f
C107 VDD1.n91 B 0.010941f
C108 VDD1.n92 B 0.025862f
C109 VDD1.n93 B 0.011585f
C110 VDD1.n94 B 0.020362f
C111 VDD1.n95 B 0.011263f
C112 VDD1.n96 B 0.025862f
C113 VDD1.n97 B 0.011585f
C114 VDD1.n98 B 0.020362f
C115 VDD1.n99 B 0.010941f
C116 VDD1.n100 B 0.025862f
C117 VDD1.n101 B 0.011585f
C118 VDD1.n102 B 0.020362f
C119 VDD1.n103 B 0.010941f
C120 VDD1.n104 B 0.025862f
C121 VDD1.n105 B 0.011585f
C122 VDD1.n106 B 0.020362f
C123 VDD1.n107 B 0.010941f
C124 VDD1.n108 B 0.025862f
C125 VDD1.n109 B 0.011585f
C126 VDD1.n110 B 0.020362f
C127 VDD1.n111 B 0.010941f
C128 VDD1.n112 B 0.025862f
C129 VDD1.n113 B 0.011585f
C130 VDD1.n114 B 0.020362f
C131 VDD1.n115 B 0.010941f
C132 VDD1.n116 B 0.019396f
C133 VDD1.n117 B 0.015277f
C134 VDD1.t1 B 0.042716f
C135 VDD1.n118 B 0.138164f
C136 VDD1.n119 B 1.42274f
C137 VDD1.n120 B 0.010941f
C138 VDD1.n121 B 0.011585f
C139 VDD1.n122 B 0.025862f
C140 VDD1.n123 B 0.025862f
C141 VDD1.n124 B 0.011585f
C142 VDD1.n125 B 0.010941f
C143 VDD1.n126 B 0.020362f
C144 VDD1.n127 B 0.020362f
C145 VDD1.n128 B 0.010941f
C146 VDD1.n129 B 0.011585f
C147 VDD1.n130 B 0.025862f
C148 VDD1.n131 B 0.025862f
C149 VDD1.n132 B 0.011585f
C150 VDD1.n133 B 0.010941f
C151 VDD1.n134 B 0.020362f
C152 VDD1.n135 B 0.020362f
C153 VDD1.n136 B 0.010941f
C154 VDD1.n137 B 0.011585f
C155 VDD1.n138 B 0.025862f
C156 VDD1.n139 B 0.025862f
C157 VDD1.n140 B 0.011585f
C158 VDD1.n141 B 0.010941f
C159 VDD1.n142 B 0.020362f
C160 VDD1.n143 B 0.020362f
C161 VDD1.n144 B 0.010941f
C162 VDD1.n145 B 0.011585f
C163 VDD1.n146 B 0.025862f
C164 VDD1.n147 B 0.025862f
C165 VDD1.n148 B 0.011585f
C166 VDD1.n149 B 0.010941f
C167 VDD1.n150 B 0.020362f
C168 VDD1.n151 B 0.020362f
C169 VDD1.n152 B 0.010941f
C170 VDD1.n153 B 0.011585f
C171 VDD1.n154 B 0.025862f
C172 VDD1.n155 B 0.025862f
C173 VDD1.n156 B 0.011585f
C174 VDD1.n157 B 0.010941f
C175 VDD1.n158 B 0.020362f
C176 VDD1.n159 B 0.020362f
C177 VDD1.n160 B 0.010941f
C178 VDD1.n161 B 0.010941f
C179 VDD1.n162 B 0.011585f
C180 VDD1.n163 B 0.025862f
C181 VDD1.n164 B 0.025862f
C182 VDD1.n165 B 0.025862f
C183 VDD1.n166 B 0.011263f
C184 VDD1.n167 B 0.010941f
C185 VDD1.n168 B 0.020362f
C186 VDD1.n169 B 0.020362f
C187 VDD1.n170 B 0.010941f
C188 VDD1.n171 B 0.011585f
C189 VDD1.n172 B 0.025862f
C190 VDD1.n173 B 0.052342f
C191 VDD1.n174 B 0.011585f
C192 VDD1.n175 B 0.010941f
C193 VDD1.n176 B 0.04623f
C194 VDD1.n177 B 0.850242f
C195 VP.t1 B 5.18135f
C196 VP.t0 B 4.43209f
C197 VP.n0 B 4.58403f
C198 VDD2.n0 B 0.026238f
C199 VDD2.n1 B 0.020116f
C200 VDD2.n2 B 0.010809f
C201 VDD2.n3 B 0.025549f
C202 VDD2.n4 B 0.011445f
C203 VDD2.n5 B 0.020116f
C204 VDD2.n6 B 0.011127f
C205 VDD2.n7 B 0.025549f
C206 VDD2.n8 B 0.011445f
C207 VDD2.n9 B 0.020116f
C208 VDD2.n10 B 0.010809f
C209 VDD2.n11 B 0.025549f
C210 VDD2.n12 B 0.011445f
C211 VDD2.n13 B 0.020116f
C212 VDD2.n14 B 0.010809f
C213 VDD2.n15 B 0.025549f
C214 VDD2.n16 B 0.011445f
C215 VDD2.n17 B 0.020116f
C216 VDD2.n18 B 0.010809f
C217 VDD2.n19 B 0.025549f
C218 VDD2.n20 B 0.011445f
C219 VDD2.n21 B 0.020116f
C220 VDD2.n22 B 0.010809f
C221 VDD2.n23 B 0.025549f
C222 VDD2.n24 B 0.011445f
C223 VDD2.n25 B 0.020116f
C224 VDD2.n26 B 0.010809f
C225 VDD2.n27 B 0.019162f
C226 VDD2.n28 B 0.015093f
C227 VDD2.t1 B 0.0422f
C228 VDD2.n29 B 0.136494f
C229 VDD2.n30 B 1.40555f
C230 VDD2.n31 B 0.010809f
C231 VDD2.n32 B 0.011445f
C232 VDD2.n33 B 0.025549f
C233 VDD2.n34 B 0.025549f
C234 VDD2.n35 B 0.011445f
C235 VDD2.n36 B 0.010809f
C236 VDD2.n37 B 0.020116f
C237 VDD2.n38 B 0.020116f
C238 VDD2.n39 B 0.010809f
C239 VDD2.n40 B 0.011445f
C240 VDD2.n41 B 0.025549f
C241 VDD2.n42 B 0.025549f
C242 VDD2.n43 B 0.011445f
C243 VDD2.n44 B 0.010809f
C244 VDD2.n45 B 0.020116f
C245 VDD2.n46 B 0.020116f
C246 VDD2.n47 B 0.010809f
C247 VDD2.n48 B 0.011445f
C248 VDD2.n49 B 0.025549f
C249 VDD2.n50 B 0.025549f
C250 VDD2.n51 B 0.011445f
C251 VDD2.n52 B 0.010809f
C252 VDD2.n53 B 0.020116f
C253 VDD2.n54 B 0.020116f
C254 VDD2.n55 B 0.010809f
C255 VDD2.n56 B 0.011445f
C256 VDD2.n57 B 0.025549f
C257 VDD2.n58 B 0.025549f
C258 VDD2.n59 B 0.011445f
C259 VDD2.n60 B 0.010809f
C260 VDD2.n61 B 0.020116f
C261 VDD2.n62 B 0.020116f
C262 VDD2.n63 B 0.010809f
C263 VDD2.n64 B 0.011445f
C264 VDD2.n65 B 0.025549f
C265 VDD2.n66 B 0.025549f
C266 VDD2.n67 B 0.011445f
C267 VDD2.n68 B 0.010809f
C268 VDD2.n69 B 0.020116f
C269 VDD2.n70 B 0.020116f
C270 VDD2.n71 B 0.010809f
C271 VDD2.n72 B 0.010809f
C272 VDD2.n73 B 0.011445f
C273 VDD2.n74 B 0.025549f
C274 VDD2.n75 B 0.025549f
C275 VDD2.n76 B 0.025549f
C276 VDD2.n77 B 0.011127f
C277 VDD2.n78 B 0.010809f
C278 VDD2.n79 B 0.020116f
C279 VDD2.n80 B 0.020116f
C280 VDD2.n81 B 0.010809f
C281 VDD2.n82 B 0.011445f
C282 VDD2.n83 B 0.025549f
C283 VDD2.n84 B 0.051709f
C284 VDD2.n85 B 0.011445f
C285 VDD2.n86 B 0.010809f
C286 VDD2.n87 B 0.045672f
C287 VDD2.n88 B 0.787471f
C288 VDD2.n89 B 0.026238f
C289 VDD2.n90 B 0.020116f
C290 VDD2.n91 B 0.010809f
C291 VDD2.n92 B 0.025549f
C292 VDD2.n93 B 0.011445f
C293 VDD2.n94 B 0.020116f
C294 VDD2.n95 B 0.011127f
C295 VDD2.n96 B 0.025549f
C296 VDD2.n97 B 0.010809f
C297 VDD2.n98 B 0.011445f
C298 VDD2.n99 B 0.020116f
C299 VDD2.n100 B 0.010809f
C300 VDD2.n101 B 0.025549f
C301 VDD2.n102 B 0.011445f
C302 VDD2.n103 B 0.020116f
C303 VDD2.n104 B 0.010809f
C304 VDD2.n105 B 0.025549f
C305 VDD2.n106 B 0.011445f
C306 VDD2.n107 B 0.020116f
C307 VDD2.n108 B 0.010809f
C308 VDD2.n109 B 0.025549f
C309 VDD2.n110 B 0.011445f
C310 VDD2.n111 B 0.020116f
C311 VDD2.n112 B 0.010809f
C312 VDD2.n113 B 0.025549f
C313 VDD2.n114 B 0.011445f
C314 VDD2.n115 B 0.020116f
C315 VDD2.n116 B 0.010809f
C316 VDD2.n117 B 0.019162f
C317 VDD2.n118 B 0.015093f
C318 VDD2.t0 B 0.0422f
C319 VDD2.n119 B 0.136494f
C320 VDD2.n120 B 1.40555f
C321 VDD2.n121 B 0.010809f
C322 VDD2.n122 B 0.011445f
C323 VDD2.n123 B 0.025549f
C324 VDD2.n124 B 0.025549f
C325 VDD2.n125 B 0.011445f
C326 VDD2.n126 B 0.010809f
C327 VDD2.n127 B 0.020116f
C328 VDD2.n128 B 0.020116f
C329 VDD2.n129 B 0.010809f
C330 VDD2.n130 B 0.011445f
C331 VDD2.n131 B 0.025549f
C332 VDD2.n132 B 0.025549f
C333 VDD2.n133 B 0.011445f
C334 VDD2.n134 B 0.010809f
C335 VDD2.n135 B 0.020116f
C336 VDD2.n136 B 0.020116f
C337 VDD2.n137 B 0.010809f
C338 VDD2.n138 B 0.011445f
C339 VDD2.n139 B 0.025549f
C340 VDD2.n140 B 0.025549f
C341 VDD2.n141 B 0.011445f
C342 VDD2.n142 B 0.010809f
C343 VDD2.n143 B 0.020116f
C344 VDD2.n144 B 0.020116f
C345 VDD2.n145 B 0.010809f
C346 VDD2.n146 B 0.011445f
C347 VDD2.n147 B 0.025549f
C348 VDD2.n148 B 0.025549f
C349 VDD2.n149 B 0.011445f
C350 VDD2.n150 B 0.010809f
C351 VDD2.n151 B 0.020116f
C352 VDD2.n152 B 0.020116f
C353 VDD2.n153 B 0.010809f
C354 VDD2.n154 B 0.011445f
C355 VDD2.n155 B 0.025549f
C356 VDD2.n156 B 0.025549f
C357 VDD2.n157 B 0.011445f
C358 VDD2.n158 B 0.010809f
C359 VDD2.n159 B 0.020116f
C360 VDD2.n160 B 0.020116f
C361 VDD2.n161 B 0.010809f
C362 VDD2.n162 B 0.011445f
C363 VDD2.n163 B 0.025549f
C364 VDD2.n164 B 0.025549f
C365 VDD2.n165 B 0.025549f
C366 VDD2.n166 B 0.011127f
C367 VDD2.n167 B 0.010809f
C368 VDD2.n168 B 0.020116f
C369 VDD2.n169 B 0.020116f
C370 VDD2.n170 B 0.010809f
C371 VDD2.n171 B 0.011445f
C372 VDD2.n172 B 0.025549f
C373 VDD2.n173 B 0.051709f
C374 VDD2.n174 B 0.011445f
C375 VDD2.n175 B 0.010809f
C376 VDD2.n176 B 0.045672f
C377 VDD2.n177 B 0.042434f
C378 VDD2.n178 B 2.98409f
C379 VTAIL.n0 B 0.026529f
C380 VTAIL.n1 B 0.020338f
C381 VTAIL.n2 B 0.010929f
C382 VTAIL.n3 B 0.025832f
C383 VTAIL.n4 B 0.011572f
C384 VTAIL.n5 B 0.020338f
C385 VTAIL.n6 B 0.01125f
C386 VTAIL.n7 B 0.025832f
C387 VTAIL.n8 B 0.011572f
C388 VTAIL.n9 B 0.020338f
C389 VTAIL.n10 B 0.010929f
C390 VTAIL.n11 B 0.025832f
C391 VTAIL.n12 B 0.011572f
C392 VTAIL.n13 B 0.020338f
C393 VTAIL.n14 B 0.010929f
C394 VTAIL.n15 B 0.025832f
C395 VTAIL.n16 B 0.011572f
C396 VTAIL.n17 B 0.020338f
C397 VTAIL.n18 B 0.010929f
C398 VTAIL.n19 B 0.025832f
C399 VTAIL.n20 B 0.011572f
C400 VTAIL.n21 B 0.020338f
C401 VTAIL.n22 B 0.010929f
C402 VTAIL.n23 B 0.025832f
C403 VTAIL.n24 B 0.011572f
C404 VTAIL.n25 B 0.020338f
C405 VTAIL.n26 B 0.010929f
C406 VTAIL.n27 B 0.019374f
C407 VTAIL.n28 B 0.01526f
C408 VTAIL.t0 B 0.042667f
C409 VTAIL.n29 B 0.138005f
C410 VTAIL.n30 B 1.42111f
C411 VTAIL.n31 B 0.010929f
C412 VTAIL.n32 B 0.011572f
C413 VTAIL.n33 B 0.025832f
C414 VTAIL.n34 B 0.025832f
C415 VTAIL.n35 B 0.011572f
C416 VTAIL.n36 B 0.010929f
C417 VTAIL.n37 B 0.020338f
C418 VTAIL.n38 B 0.020338f
C419 VTAIL.n39 B 0.010929f
C420 VTAIL.n40 B 0.011572f
C421 VTAIL.n41 B 0.025832f
C422 VTAIL.n42 B 0.025832f
C423 VTAIL.n43 B 0.011572f
C424 VTAIL.n44 B 0.010929f
C425 VTAIL.n45 B 0.020338f
C426 VTAIL.n46 B 0.020338f
C427 VTAIL.n47 B 0.010929f
C428 VTAIL.n48 B 0.011572f
C429 VTAIL.n49 B 0.025832f
C430 VTAIL.n50 B 0.025832f
C431 VTAIL.n51 B 0.011572f
C432 VTAIL.n52 B 0.010929f
C433 VTAIL.n53 B 0.020338f
C434 VTAIL.n54 B 0.020338f
C435 VTAIL.n55 B 0.010929f
C436 VTAIL.n56 B 0.011572f
C437 VTAIL.n57 B 0.025832f
C438 VTAIL.n58 B 0.025832f
C439 VTAIL.n59 B 0.011572f
C440 VTAIL.n60 B 0.010929f
C441 VTAIL.n61 B 0.020338f
C442 VTAIL.n62 B 0.020338f
C443 VTAIL.n63 B 0.010929f
C444 VTAIL.n64 B 0.011572f
C445 VTAIL.n65 B 0.025832f
C446 VTAIL.n66 B 0.025832f
C447 VTAIL.n67 B 0.011572f
C448 VTAIL.n68 B 0.010929f
C449 VTAIL.n69 B 0.020338f
C450 VTAIL.n70 B 0.020338f
C451 VTAIL.n71 B 0.010929f
C452 VTAIL.n72 B 0.010929f
C453 VTAIL.n73 B 0.011572f
C454 VTAIL.n74 B 0.025832f
C455 VTAIL.n75 B 0.025832f
C456 VTAIL.n76 B 0.025832f
C457 VTAIL.n77 B 0.01125f
C458 VTAIL.n78 B 0.010929f
C459 VTAIL.n79 B 0.020338f
C460 VTAIL.n80 B 0.020338f
C461 VTAIL.n81 B 0.010929f
C462 VTAIL.n82 B 0.011572f
C463 VTAIL.n83 B 0.025832f
C464 VTAIL.n84 B 0.052282f
C465 VTAIL.n85 B 0.011572f
C466 VTAIL.n86 B 0.010929f
C467 VTAIL.n87 B 0.046178f
C468 VTAIL.n88 B 0.028854f
C469 VTAIL.n89 B 1.77349f
C470 VTAIL.n90 B 0.026529f
C471 VTAIL.n91 B 0.020338f
C472 VTAIL.n92 B 0.010929f
C473 VTAIL.n93 B 0.025832f
C474 VTAIL.n94 B 0.011572f
C475 VTAIL.n95 B 0.020338f
C476 VTAIL.n96 B 0.01125f
C477 VTAIL.n97 B 0.025832f
C478 VTAIL.n98 B 0.010929f
C479 VTAIL.n99 B 0.011572f
C480 VTAIL.n100 B 0.020338f
C481 VTAIL.n101 B 0.010929f
C482 VTAIL.n102 B 0.025832f
C483 VTAIL.n103 B 0.011572f
C484 VTAIL.n104 B 0.020338f
C485 VTAIL.n105 B 0.010929f
C486 VTAIL.n106 B 0.025832f
C487 VTAIL.n107 B 0.011572f
C488 VTAIL.n108 B 0.020338f
C489 VTAIL.n109 B 0.010929f
C490 VTAIL.n110 B 0.025832f
C491 VTAIL.n111 B 0.011572f
C492 VTAIL.n112 B 0.020338f
C493 VTAIL.n113 B 0.010929f
C494 VTAIL.n114 B 0.025832f
C495 VTAIL.n115 B 0.011572f
C496 VTAIL.n116 B 0.020338f
C497 VTAIL.n117 B 0.010929f
C498 VTAIL.n118 B 0.019374f
C499 VTAIL.n119 B 0.01526f
C500 VTAIL.t2 B 0.042667f
C501 VTAIL.n120 B 0.138005f
C502 VTAIL.n121 B 1.42111f
C503 VTAIL.n122 B 0.010929f
C504 VTAIL.n123 B 0.011572f
C505 VTAIL.n124 B 0.025832f
C506 VTAIL.n125 B 0.025832f
C507 VTAIL.n126 B 0.011572f
C508 VTAIL.n127 B 0.010929f
C509 VTAIL.n128 B 0.020338f
C510 VTAIL.n129 B 0.020338f
C511 VTAIL.n130 B 0.010929f
C512 VTAIL.n131 B 0.011572f
C513 VTAIL.n132 B 0.025832f
C514 VTAIL.n133 B 0.025832f
C515 VTAIL.n134 B 0.011572f
C516 VTAIL.n135 B 0.010929f
C517 VTAIL.n136 B 0.020338f
C518 VTAIL.n137 B 0.020338f
C519 VTAIL.n138 B 0.010929f
C520 VTAIL.n139 B 0.011572f
C521 VTAIL.n140 B 0.025832f
C522 VTAIL.n141 B 0.025832f
C523 VTAIL.n142 B 0.011572f
C524 VTAIL.n143 B 0.010929f
C525 VTAIL.n144 B 0.020338f
C526 VTAIL.n145 B 0.020338f
C527 VTAIL.n146 B 0.010929f
C528 VTAIL.n147 B 0.011572f
C529 VTAIL.n148 B 0.025832f
C530 VTAIL.n149 B 0.025832f
C531 VTAIL.n150 B 0.011572f
C532 VTAIL.n151 B 0.010929f
C533 VTAIL.n152 B 0.020338f
C534 VTAIL.n153 B 0.020338f
C535 VTAIL.n154 B 0.010929f
C536 VTAIL.n155 B 0.011572f
C537 VTAIL.n156 B 0.025832f
C538 VTAIL.n157 B 0.025832f
C539 VTAIL.n158 B 0.011572f
C540 VTAIL.n159 B 0.010929f
C541 VTAIL.n160 B 0.020338f
C542 VTAIL.n161 B 0.020338f
C543 VTAIL.n162 B 0.010929f
C544 VTAIL.n163 B 0.011572f
C545 VTAIL.n164 B 0.025832f
C546 VTAIL.n165 B 0.025832f
C547 VTAIL.n166 B 0.025832f
C548 VTAIL.n167 B 0.01125f
C549 VTAIL.n168 B 0.010929f
C550 VTAIL.n169 B 0.020338f
C551 VTAIL.n170 B 0.020338f
C552 VTAIL.n171 B 0.010929f
C553 VTAIL.n172 B 0.011572f
C554 VTAIL.n173 B 0.025832f
C555 VTAIL.n174 B 0.052282f
C556 VTAIL.n175 B 0.011572f
C557 VTAIL.n176 B 0.010929f
C558 VTAIL.n177 B 0.046178f
C559 VTAIL.n178 B 0.028854f
C560 VTAIL.n179 B 1.82957f
C561 VTAIL.n180 B 0.026529f
C562 VTAIL.n181 B 0.020338f
C563 VTAIL.n182 B 0.010929f
C564 VTAIL.n183 B 0.025832f
C565 VTAIL.n184 B 0.011572f
C566 VTAIL.n185 B 0.020338f
C567 VTAIL.n186 B 0.01125f
C568 VTAIL.n187 B 0.025832f
C569 VTAIL.n188 B 0.010929f
C570 VTAIL.n189 B 0.011572f
C571 VTAIL.n190 B 0.020338f
C572 VTAIL.n191 B 0.010929f
C573 VTAIL.n192 B 0.025832f
C574 VTAIL.n193 B 0.011572f
C575 VTAIL.n194 B 0.020338f
C576 VTAIL.n195 B 0.010929f
C577 VTAIL.n196 B 0.025832f
C578 VTAIL.n197 B 0.011572f
C579 VTAIL.n198 B 0.020338f
C580 VTAIL.n199 B 0.010929f
C581 VTAIL.n200 B 0.025832f
C582 VTAIL.n201 B 0.011572f
C583 VTAIL.n202 B 0.020338f
C584 VTAIL.n203 B 0.010929f
C585 VTAIL.n204 B 0.025832f
C586 VTAIL.n205 B 0.011572f
C587 VTAIL.n206 B 0.020338f
C588 VTAIL.n207 B 0.010929f
C589 VTAIL.n208 B 0.019374f
C590 VTAIL.n209 B 0.01526f
C591 VTAIL.t1 B 0.042667f
C592 VTAIL.n210 B 0.138005f
C593 VTAIL.n211 B 1.42111f
C594 VTAIL.n212 B 0.010929f
C595 VTAIL.n213 B 0.011572f
C596 VTAIL.n214 B 0.025832f
C597 VTAIL.n215 B 0.025832f
C598 VTAIL.n216 B 0.011572f
C599 VTAIL.n217 B 0.010929f
C600 VTAIL.n218 B 0.020338f
C601 VTAIL.n219 B 0.020338f
C602 VTAIL.n220 B 0.010929f
C603 VTAIL.n221 B 0.011572f
C604 VTAIL.n222 B 0.025832f
C605 VTAIL.n223 B 0.025832f
C606 VTAIL.n224 B 0.011572f
C607 VTAIL.n225 B 0.010929f
C608 VTAIL.n226 B 0.020338f
C609 VTAIL.n227 B 0.020338f
C610 VTAIL.n228 B 0.010929f
C611 VTAIL.n229 B 0.011572f
C612 VTAIL.n230 B 0.025832f
C613 VTAIL.n231 B 0.025832f
C614 VTAIL.n232 B 0.011572f
C615 VTAIL.n233 B 0.010929f
C616 VTAIL.n234 B 0.020338f
C617 VTAIL.n235 B 0.020338f
C618 VTAIL.n236 B 0.010929f
C619 VTAIL.n237 B 0.011572f
C620 VTAIL.n238 B 0.025832f
C621 VTAIL.n239 B 0.025832f
C622 VTAIL.n240 B 0.011572f
C623 VTAIL.n241 B 0.010929f
C624 VTAIL.n242 B 0.020338f
C625 VTAIL.n243 B 0.020338f
C626 VTAIL.n244 B 0.010929f
C627 VTAIL.n245 B 0.011572f
C628 VTAIL.n246 B 0.025832f
C629 VTAIL.n247 B 0.025832f
C630 VTAIL.n248 B 0.011572f
C631 VTAIL.n249 B 0.010929f
C632 VTAIL.n250 B 0.020338f
C633 VTAIL.n251 B 0.020338f
C634 VTAIL.n252 B 0.010929f
C635 VTAIL.n253 B 0.011572f
C636 VTAIL.n254 B 0.025832f
C637 VTAIL.n255 B 0.025832f
C638 VTAIL.n256 B 0.025832f
C639 VTAIL.n257 B 0.01125f
C640 VTAIL.n258 B 0.010929f
C641 VTAIL.n259 B 0.020338f
C642 VTAIL.n260 B 0.020338f
C643 VTAIL.n261 B 0.010929f
C644 VTAIL.n262 B 0.011572f
C645 VTAIL.n263 B 0.025832f
C646 VTAIL.n264 B 0.052282f
C647 VTAIL.n265 B 0.011572f
C648 VTAIL.n266 B 0.010929f
C649 VTAIL.n267 B 0.046178f
C650 VTAIL.n268 B 0.028854f
C651 VTAIL.n269 B 1.59002f
C652 VTAIL.n270 B 0.026529f
C653 VTAIL.n271 B 0.020338f
C654 VTAIL.n272 B 0.010929f
C655 VTAIL.n273 B 0.025832f
C656 VTAIL.n274 B 0.011572f
C657 VTAIL.n275 B 0.020338f
C658 VTAIL.n276 B 0.01125f
C659 VTAIL.n277 B 0.025832f
C660 VTAIL.n278 B 0.011572f
C661 VTAIL.n279 B 0.020338f
C662 VTAIL.n280 B 0.010929f
C663 VTAIL.n281 B 0.025832f
C664 VTAIL.n282 B 0.011572f
C665 VTAIL.n283 B 0.020338f
C666 VTAIL.n284 B 0.010929f
C667 VTAIL.n285 B 0.025832f
C668 VTAIL.n286 B 0.011572f
C669 VTAIL.n287 B 0.020338f
C670 VTAIL.n288 B 0.010929f
C671 VTAIL.n289 B 0.025832f
C672 VTAIL.n290 B 0.011572f
C673 VTAIL.n291 B 0.020338f
C674 VTAIL.n292 B 0.010929f
C675 VTAIL.n293 B 0.025832f
C676 VTAIL.n294 B 0.011572f
C677 VTAIL.n295 B 0.020338f
C678 VTAIL.n296 B 0.010929f
C679 VTAIL.n297 B 0.019374f
C680 VTAIL.n298 B 0.01526f
C681 VTAIL.t3 B 0.042667f
C682 VTAIL.n299 B 0.138005f
C683 VTAIL.n300 B 1.42111f
C684 VTAIL.n301 B 0.010929f
C685 VTAIL.n302 B 0.011572f
C686 VTAIL.n303 B 0.025832f
C687 VTAIL.n304 B 0.025832f
C688 VTAIL.n305 B 0.011572f
C689 VTAIL.n306 B 0.010929f
C690 VTAIL.n307 B 0.020338f
C691 VTAIL.n308 B 0.020338f
C692 VTAIL.n309 B 0.010929f
C693 VTAIL.n310 B 0.011572f
C694 VTAIL.n311 B 0.025832f
C695 VTAIL.n312 B 0.025832f
C696 VTAIL.n313 B 0.011572f
C697 VTAIL.n314 B 0.010929f
C698 VTAIL.n315 B 0.020338f
C699 VTAIL.n316 B 0.020338f
C700 VTAIL.n317 B 0.010929f
C701 VTAIL.n318 B 0.011572f
C702 VTAIL.n319 B 0.025832f
C703 VTAIL.n320 B 0.025832f
C704 VTAIL.n321 B 0.011572f
C705 VTAIL.n322 B 0.010929f
C706 VTAIL.n323 B 0.020338f
C707 VTAIL.n324 B 0.020338f
C708 VTAIL.n325 B 0.010929f
C709 VTAIL.n326 B 0.011572f
C710 VTAIL.n327 B 0.025832f
C711 VTAIL.n328 B 0.025832f
C712 VTAIL.n329 B 0.011572f
C713 VTAIL.n330 B 0.010929f
C714 VTAIL.n331 B 0.020338f
C715 VTAIL.n332 B 0.020338f
C716 VTAIL.n333 B 0.010929f
C717 VTAIL.n334 B 0.011572f
C718 VTAIL.n335 B 0.025832f
C719 VTAIL.n336 B 0.025832f
C720 VTAIL.n337 B 0.011572f
C721 VTAIL.n338 B 0.010929f
C722 VTAIL.n339 B 0.020338f
C723 VTAIL.n340 B 0.020338f
C724 VTAIL.n341 B 0.010929f
C725 VTAIL.n342 B 0.010929f
C726 VTAIL.n343 B 0.011572f
C727 VTAIL.n344 B 0.025832f
C728 VTAIL.n345 B 0.025832f
C729 VTAIL.n346 B 0.025832f
C730 VTAIL.n347 B 0.01125f
C731 VTAIL.n348 B 0.010929f
C732 VTAIL.n349 B 0.020338f
C733 VTAIL.n350 B 0.020338f
C734 VTAIL.n351 B 0.010929f
C735 VTAIL.n352 B 0.011572f
C736 VTAIL.n353 B 0.025832f
C737 VTAIL.n354 B 0.052282f
C738 VTAIL.n355 B 0.011572f
C739 VTAIL.n356 B 0.010929f
C740 VTAIL.n357 B 0.046178f
C741 VTAIL.n358 B 0.028854f
C742 VTAIL.n359 B 1.49554f
C743 VN.t0 B 4.33534f
C744 VN.t1 B 5.05902f
.ends

