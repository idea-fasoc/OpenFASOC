* NGSPICE file created from diff_pair_sample_1742.ext - technology: sky130A

.subckt diff_pair_sample_1742 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0.3663 ps=2.55 w=2.22 l=3.43
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.8658 ps=5.22 w=2.22 l=3.43
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0 ps=0 w=2.22 l=3.43
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0 ps=0 w=2.22 l=3.43
X4 VTAIL.t6 VP.t2 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.3663 ps=2.55 w=2.22 l=3.43
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0 ps=0 w=2.22 l=3.43
X6 VDD1.t2 VP.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0.3663 ps=2.55 w=2.22 l=3.43
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0 ps=0 w=2.22 l=3.43
X8 VTAIL.t2 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.3663 ps=2.55 w=2.22 l=3.43
X9 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.8658 ps=5.22 w=2.22 l=3.43
X10 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.8658 ps=5.22 w=2.22 l=3.43
X11 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0.3663 ps=2.55 w=2.22 l=3.43
X12 VDD1.t1 VP.t4 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.8658 ps=5.22 w=2.22 l=3.43
X13 VTAIL.t9 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.3663 ps=2.55 w=2.22 l=3.43
X14 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8658 pd=5.22 as=0.3663 ps=2.55 w=2.22 l=3.43
X15 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3663 pd=2.55 as=0.3663 ps=2.55 w=2.22 l=3.43
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n27 VP.n8 77.2324
R23 VP.n51 VP.n0 77.2324
R24 VP.n26 VP.n9 77.2324
R25 VP.n35 VP.n6 52.0954
R26 VP.n43 VP.n2 52.0954
R27 VP.n18 VP.n11 52.0954
R28 VP.n14 VP.n13 50.0561
R29 VP.n14 VP.t0 49.3621
R30 VP.n27 VP.n26 44.6355
R31 VP.n31 VP.n6 28.7258
R32 VP.n47 VP.n2 28.7258
R33 VP.n22 VP.n11 28.7258
R34 VP.n30 VP.n29 24.3439
R35 VP.n31 VP.n30 24.3439
R36 VP.n36 VP.n35 24.3439
R37 VP.n37 VP.n36 24.3439
R38 VP.n37 VP.n4 24.3439
R39 VP.n41 VP.n4 24.3439
R40 VP.n42 VP.n41 24.3439
R41 VP.n43 VP.n42 24.3439
R42 VP.n48 VP.n47 24.3439
R43 VP.n49 VP.n48 24.3439
R44 VP.n23 VP.n22 24.3439
R45 VP.n24 VP.n23 24.3439
R46 VP.n16 VP.n13 24.3439
R47 VP.n17 VP.n16 24.3439
R48 VP.n18 VP.n17 24.3439
R49 VP.n4 VP.t2 15.5988
R50 VP.n8 VP.t3 15.5988
R51 VP.n0 VP.t1 15.5988
R52 VP.n13 VP.t5 15.5988
R53 VP.n9 VP.t4 15.5988
R54 VP.n29 VP.n8 12.6591
R55 VP.n49 VP.n0 12.6591
R56 VP.n24 VP.n9 12.6591
R57 VP.n15 VP.n14 3.07272
R58 VP.n26 VP.n25 0.355081
R59 VP.n28 VP.n27 0.355081
R60 VP.n51 VP.n50 0.355081
R61 VP VP.n51 0.26685
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n10 VTAIL.t8 86.4835
R83 VTAIL.n11 VTAIL.t4 86.4835
R84 VTAIL.n2 VTAIL.t10 86.4835
R85 VTAIL.n7 VTAIL.t5 86.4834
R86 VTAIL.n9 VTAIL.n8 77.5647
R87 VTAIL.n6 VTAIL.n5 77.5647
R88 VTAIL.n1 VTAIL.n0 77.5644
R89 VTAIL.n4 VTAIL.n3 77.5644
R90 VTAIL.n6 VTAIL.n4 20.7634
R91 VTAIL.n11 VTAIL.n10 17.5221
R92 VTAIL.n0 VTAIL.t1 8.91942
R93 VTAIL.n0 VTAIL.t0 8.91942
R94 VTAIL.n3 VTAIL.t11 8.91942
R95 VTAIL.n3 VTAIL.t6 8.91942
R96 VTAIL.n8 VTAIL.t7 8.91942
R97 VTAIL.n8 VTAIL.t9 8.91942
R98 VTAIL.n5 VTAIL.t3 8.91942
R99 VTAIL.n5 VTAIL.t2 8.91942
R100 VTAIL.n7 VTAIL.n6 3.24188
R101 VTAIL.n10 VTAIL.n9 3.24188
R102 VTAIL.n4 VTAIL.n2 3.24188
R103 VTAIL VTAIL.n11 2.37334
R104 VTAIL.n9 VTAIL.n7 2.09102
R105 VTAIL.n2 VTAIL.n1 2.09102
R106 VTAIL VTAIL.n1 0.869035
R107 VDD1 VDD1.t5 105.651
R108 VDD1.n1 VDD1.t2 105.537
R109 VDD1.n1 VDD1.n0 94.9982
R110 VDD1.n3 VDD1.n2 94.2434
R111 VDD1.n3 VDD1.n1 38.3673
R112 VDD1.n2 VDD1.t0 8.91942
R113 VDD1.n2 VDD1.t1 8.91942
R114 VDD1.n0 VDD1.t3 8.91942
R115 VDD1.n0 VDD1.t4 8.91942
R116 VDD1 VDD1.n3 0.752655
R117 B.n607 B.n606 585
R118 B.n608 B.n607 585
R119 B.n186 B.n115 585
R120 B.n185 B.n184 585
R121 B.n183 B.n182 585
R122 B.n181 B.n180 585
R123 B.n179 B.n178 585
R124 B.n177 B.n176 585
R125 B.n175 B.n174 585
R126 B.n173 B.n172 585
R127 B.n171 B.n170 585
R128 B.n169 B.n168 585
R129 B.n167 B.n166 585
R130 B.n165 B.n164 585
R131 B.n163 B.n162 585
R132 B.n161 B.n160 585
R133 B.n159 B.n158 585
R134 B.n157 B.n156 585
R135 B.n155 B.n154 585
R136 B.n153 B.n152 585
R137 B.n151 B.n150 585
R138 B.n149 B.n148 585
R139 B.n147 B.n146 585
R140 B.n144 B.n143 585
R141 B.n142 B.n141 585
R142 B.n140 B.n139 585
R143 B.n138 B.n137 585
R144 B.n136 B.n135 585
R145 B.n134 B.n133 585
R146 B.n132 B.n131 585
R147 B.n130 B.n129 585
R148 B.n128 B.n127 585
R149 B.n126 B.n125 585
R150 B.n124 B.n123 585
R151 B.n122 B.n121 585
R152 B.n96 B.n95 585
R153 B.n605 B.n97 585
R154 B.n609 B.n97 585
R155 B.n604 B.n603 585
R156 B.n603 B.n93 585
R157 B.n602 B.n92 585
R158 B.n615 B.n92 585
R159 B.n601 B.n91 585
R160 B.n616 B.n91 585
R161 B.n600 B.n90 585
R162 B.n617 B.n90 585
R163 B.n599 B.n598 585
R164 B.n598 B.n86 585
R165 B.n597 B.n85 585
R166 B.n623 B.n85 585
R167 B.n596 B.n84 585
R168 B.n624 B.n84 585
R169 B.n595 B.n83 585
R170 B.n625 B.n83 585
R171 B.n594 B.n593 585
R172 B.n593 B.n79 585
R173 B.n592 B.n78 585
R174 B.n631 B.n78 585
R175 B.n591 B.n77 585
R176 B.n632 B.n77 585
R177 B.n590 B.n76 585
R178 B.n633 B.n76 585
R179 B.n589 B.n588 585
R180 B.n588 B.n72 585
R181 B.n587 B.n71 585
R182 B.n639 B.n71 585
R183 B.n586 B.n70 585
R184 B.n640 B.n70 585
R185 B.n585 B.n69 585
R186 B.n641 B.n69 585
R187 B.n584 B.n583 585
R188 B.n583 B.n65 585
R189 B.n582 B.n64 585
R190 B.n647 B.n64 585
R191 B.n581 B.n63 585
R192 B.n648 B.n63 585
R193 B.n580 B.n62 585
R194 B.n649 B.n62 585
R195 B.n579 B.n578 585
R196 B.n578 B.n58 585
R197 B.n577 B.n57 585
R198 B.n655 B.n57 585
R199 B.n576 B.n56 585
R200 B.n656 B.n56 585
R201 B.n575 B.n55 585
R202 B.n657 B.n55 585
R203 B.n574 B.n573 585
R204 B.n573 B.n51 585
R205 B.n572 B.n50 585
R206 B.n663 B.n50 585
R207 B.n571 B.n49 585
R208 B.n664 B.n49 585
R209 B.n570 B.n48 585
R210 B.n665 B.n48 585
R211 B.n569 B.n568 585
R212 B.n568 B.n44 585
R213 B.n567 B.n43 585
R214 B.n671 B.n43 585
R215 B.n566 B.n42 585
R216 B.n672 B.n42 585
R217 B.n565 B.n41 585
R218 B.n673 B.n41 585
R219 B.n564 B.n563 585
R220 B.n563 B.n37 585
R221 B.n562 B.n36 585
R222 B.n679 B.n36 585
R223 B.n561 B.n35 585
R224 B.n680 B.n35 585
R225 B.n560 B.n34 585
R226 B.n681 B.n34 585
R227 B.n559 B.n558 585
R228 B.n558 B.n30 585
R229 B.n557 B.n29 585
R230 B.n687 B.n29 585
R231 B.n556 B.n28 585
R232 B.n688 B.n28 585
R233 B.n555 B.n27 585
R234 B.n689 B.n27 585
R235 B.n554 B.n553 585
R236 B.n553 B.n23 585
R237 B.n552 B.n22 585
R238 B.n695 B.n22 585
R239 B.n551 B.n21 585
R240 B.n696 B.n21 585
R241 B.n550 B.n20 585
R242 B.n697 B.n20 585
R243 B.n549 B.n548 585
R244 B.n548 B.n19 585
R245 B.n547 B.n15 585
R246 B.n703 B.n15 585
R247 B.n546 B.n14 585
R248 B.n704 B.n14 585
R249 B.n545 B.n13 585
R250 B.n705 B.n13 585
R251 B.n544 B.n543 585
R252 B.n543 B.n12 585
R253 B.n542 B.n541 585
R254 B.n542 B.n8 585
R255 B.n540 B.n7 585
R256 B.n712 B.n7 585
R257 B.n539 B.n6 585
R258 B.n713 B.n6 585
R259 B.n538 B.n5 585
R260 B.n714 B.n5 585
R261 B.n537 B.n536 585
R262 B.n536 B.n4 585
R263 B.n535 B.n187 585
R264 B.n535 B.n534 585
R265 B.n525 B.n188 585
R266 B.n189 B.n188 585
R267 B.n527 B.n526 585
R268 B.n528 B.n527 585
R269 B.n524 B.n194 585
R270 B.n194 B.n193 585
R271 B.n523 B.n522 585
R272 B.n522 B.n521 585
R273 B.n196 B.n195 585
R274 B.n514 B.n196 585
R275 B.n513 B.n512 585
R276 B.n515 B.n513 585
R277 B.n511 B.n201 585
R278 B.n201 B.n200 585
R279 B.n510 B.n509 585
R280 B.n509 B.n508 585
R281 B.n203 B.n202 585
R282 B.n204 B.n203 585
R283 B.n501 B.n500 585
R284 B.n502 B.n501 585
R285 B.n499 B.n209 585
R286 B.n209 B.n208 585
R287 B.n498 B.n497 585
R288 B.n497 B.n496 585
R289 B.n211 B.n210 585
R290 B.n212 B.n211 585
R291 B.n489 B.n488 585
R292 B.n490 B.n489 585
R293 B.n487 B.n217 585
R294 B.n217 B.n216 585
R295 B.n486 B.n485 585
R296 B.n485 B.n484 585
R297 B.n219 B.n218 585
R298 B.n220 B.n219 585
R299 B.n477 B.n476 585
R300 B.n478 B.n477 585
R301 B.n475 B.n225 585
R302 B.n225 B.n224 585
R303 B.n474 B.n473 585
R304 B.n473 B.n472 585
R305 B.n227 B.n226 585
R306 B.n228 B.n227 585
R307 B.n465 B.n464 585
R308 B.n466 B.n465 585
R309 B.n463 B.n233 585
R310 B.n233 B.n232 585
R311 B.n462 B.n461 585
R312 B.n461 B.n460 585
R313 B.n235 B.n234 585
R314 B.n236 B.n235 585
R315 B.n453 B.n452 585
R316 B.n454 B.n453 585
R317 B.n451 B.n240 585
R318 B.n244 B.n240 585
R319 B.n450 B.n449 585
R320 B.n449 B.n448 585
R321 B.n242 B.n241 585
R322 B.n243 B.n242 585
R323 B.n441 B.n440 585
R324 B.n442 B.n441 585
R325 B.n439 B.n249 585
R326 B.n249 B.n248 585
R327 B.n438 B.n437 585
R328 B.n437 B.n436 585
R329 B.n251 B.n250 585
R330 B.n252 B.n251 585
R331 B.n429 B.n428 585
R332 B.n430 B.n429 585
R333 B.n427 B.n257 585
R334 B.n257 B.n256 585
R335 B.n426 B.n425 585
R336 B.n425 B.n424 585
R337 B.n259 B.n258 585
R338 B.n260 B.n259 585
R339 B.n417 B.n416 585
R340 B.n418 B.n417 585
R341 B.n415 B.n265 585
R342 B.n265 B.n264 585
R343 B.n414 B.n413 585
R344 B.n413 B.n412 585
R345 B.n267 B.n266 585
R346 B.n268 B.n267 585
R347 B.n405 B.n404 585
R348 B.n406 B.n405 585
R349 B.n403 B.n273 585
R350 B.n273 B.n272 585
R351 B.n402 B.n401 585
R352 B.n401 B.n400 585
R353 B.n275 B.n274 585
R354 B.n276 B.n275 585
R355 B.n393 B.n392 585
R356 B.n394 B.n393 585
R357 B.n391 B.n281 585
R358 B.n281 B.n280 585
R359 B.n390 B.n389 585
R360 B.n389 B.n388 585
R361 B.n283 B.n282 585
R362 B.n284 B.n283 585
R363 B.n381 B.n380 585
R364 B.n382 B.n381 585
R365 B.n287 B.n286 585
R366 B.n313 B.n312 585
R367 B.n314 B.n310 585
R368 B.n310 B.n288 585
R369 B.n316 B.n315 585
R370 B.n318 B.n309 585
R371 B.n321 B.n320 585
R372 B.n322 B.n308 585
R373 B.n324 B.n323 585
R374 B.n326 B.n307 585
R375 B.n329 B.n328 585
R376 B.n330 B.n306 585
R377 B.n332 B.n331 585
R378 B.n334 B.n305 585
R379 B.n337 B.n336 585
R380 B.n338 B.n301 585
R381 B.n340 B.n339 585
R382 B.n342 B.n300 585
R383 B.n345 B.n344 585
R384 B.n346 B.n299 585
R385 B.n348 B.n347 585
R386 B.n350 B.n298 585
R387 B.n353 B.n352 585
R388 B.n355 B.n295 585
R389 B.n357 B.n356 585
R390 B.n359 B.n294 585
R391 B.n362 B.n361 585
R392 B.n363 B.n293 585
R393 B.n365 B.n364 585
R394 B.n367 B.n292 585
R395 B.n370 B.n369 585
R396 B.n371 B.n291 585
R397 B.n373 B.n372 585
R398 B.n375 B.n290 585
R399 B.n378 B.n377 585
R400 B.n379 B.n289 585
R401 B.n384 B.n383 585
R402 B.n383 B.n382 585
R403 B.n385 B.n285 585
R404 B.n285 B.n284 585
R405 B.n387 B.n386 585
R406 B.n388 B.n387 585
R407 B.n279 B.n278 585
R408 B.n280 B.n279 585
R409 B.n396 B.n395 585
R410 B.n395 B.n394 585
R411 B.n397 B.n277 585
R412 B.n277 B.n276 585
R413 B.n399 B.n398 585
R414 B.n400 B.n399 585
R415 B.n271 B.n270 585
R416 B.n272 B.n271 585
R417 B.n408 B.n407 585
R418 B.n407 B.n406 585
R419 B.n409 B.n269 585
R420 B.n269 B.n268 585
R421 B.n411 B.n410 585
R422 B.n412 B.n411 585
R423 B.n263 B.n262 585
R424 B.n264 B.n263 585
R425 B.n420 B.n419 585
R426 B.n419 B.n418 585
R427 B.n421 B.n261 585
R428 B.n261 B.n260 585
R429 B.n423 B.n422 585
R430 B.n424 B.n423 585
R431 B.n255 B.n254 585
R432 B.n256 B.n255 585
R433 B.n432 B.n431 585
R434 B.n431 B.n430 585
R435 B.n433 B.n253 585
R436 B.n253 B.n252 585
R437 B.n435 B.n434 585
R438 B.n436 B.n435 585
R439 B.n247 B.n246 585
R440 B.n248 B.n247 585
R441 B.n444 B.n443 585
R442 B.n443 B.n442 585
R443 B.n445 B.n245 585
R444 B.n245 B.n243 585
R445 B.n447 B.n446 585
R446 B.n448 B.n447 585
R447 B.n239 B.n238 585
R448 B.n244 B.n239 585
R449 B.n456 B.n455 585
R450 B.n455 B.n454 585
R451 B.n457 B.n237 585
R452 B.n237 B.n236 585
R453 B.n459 B.n458 585
R454 B.n460 B.n459 585
R455 B.n231 B.n230 585
R456 B.n232 B.n231 585
R457 B.n468 B.n467 585
R458 B.n467 B.n466 585
R459 B.n469 B.n229 585
R460 B.n229 B.n228 585
R461 B.n471 B.n470 585
R462 B.n472 B.n471 585
R463 B.n223 B.n222 585
R464 B.n224 B.n223 585
R465 B.n480 B.n479 585
R466 B.n479 B.n478 585
R467 B.n481 B.n221 585
R468 B.n221 B.n220 585
R469 B.n483 B.n482 585
R470 B.n484 B.n483 585
R471 B.n215 B.n214 585
R472 B.n216 B.n215 585
R473 B.n492 B.n491 585
R474 B.n491 B.n490 585
R475 B.n493 B.n213 585
R476 B.n213 B.n212 585
R477 B.n495 B.n494 585
R478 B.n496 B.n495 585
R479 B.n207 B.n206 585
R480 B.n208 B.n207 585
R481 B.n504 B.n503 585
R482 B.n503 B.n502 585
R483 B.n505 B.n205 585
R484 B.n205 B.n204 585
R485 B.n507 B.n506 585
R486 B.n508 B.n507 585
R487 B.n199 B.n198 585
R488 B.n200 B.n199 585
R489 B.n517 B.n516 585
R490 B.n516 B.n515 585
R491 B.n518 B.n197 585
R492 B.n514 B.n197 585
R493 B.n520 B.n519 585
R494 B.n521 B.n520 585
R495 B.n192 B.n191 585
R496 B.n193 B.n192 585
R497 B.n530 B.n529 585
R498 B.n529 B.n528 585
R499 B.n531 B.n190 585
R500 B.n190 B.n189 585
R501 B.n533 B.n532 585
R502 B.n534 B.n533 585
R503 B.n3 B.n0 585
R504 B.n4 B.n3 585
R505 B.n711 B.n1 585
R506 B.n712 B.n711 585
R507 B.n710 B.n709 585
R508 B.n710 B.n8 585
R509 B.n708 B.n9 585
R510 B.n12 B.n9 585
R511 B.n707 B.n706 585
R512 B.n706 B.n705 585
R513 B.n11 B.n10 585
R514 B.n704 B.n11 585
R515 B.n702 B.n701 585
R516 B.n703 B.n702 585
R517 B.n700 B.n16 585
R518 B.n19 B.n16 585
R519 B.n699 B.n698 585
R520 B.n698 B.n697 585
R521 B.n18 B.n17 585
R522 B.n696 B.n18 585
R523 B.n694 B.n693 585
R524 B.n695 B.n694 585
R525 B.n692 B.n24 585
R526 B.n24 B.n23 585
R527 B.n691 B.n690 585
R528 B.n690 B.n689 585
R529 B.n26 B.n25 585
R530 B.n688 B.n26 585
R531 B.n686 B.n685 585
R532 B.n687 B.n686 585
R533 B.n684 B.n31 585
R534 B.n31 B.n30 585
R535 B.n683 B.n682 585
R536 B.n682 B.n681 585
R537 B.n33 B.n32 585
R538 B.n680 B.n33 585
R539 B.n678 B.n677 585
R540 B.n679 B.n678 585
R541 B.n676 B.n38 585
R542 B.n38 B.n37 585
R543 B.n675 B.n674 585
R544 B.n674 B.n673 585
R545 B.n40 B.n39 585
R546 B.n672 B.n40 585
R547 B.n670 B.n669 585
R548 B.n671 B.n670 585
R549 B.n668 B.n45 585
R550 B.n45 B.n44 585
R551 B.n667 B.n666 585
R552 B.n666 B.n665 585
R553 B.n47 B.n46 585
R554 B.n664 B.n47 585
R555 B.n662 B.n661 585
R556 B.n663 B.n662 585
R557 B.n660 B.n52 585
R558 B.n52 B.n51 585
R559 B.n659 B.n658 585
R560 B.n658 B.n657 585
R561 B.n54 B.n53 585
R562 B.n656 B.n54 585
R563 B.n654 B.n653 585
R564 B.n655 B.n654 585
R565 B.n652 B.n59 585
R566 B.n59 B.n58 585
R567 B.n651 B.n650 585
R568 B.n650 B.n649 585
R569 B.n61 B.n60 585
R570 B.n648 B.n61 585
R571 B.n646 B.n645 585
R572 B.n647 B.n646 585
R573 B.n644 B.n66 585
R574 B.n66 B.n65 585
R575 B.n643 B.n642 585
R576 B.n642 B.n641 585
R577 B.n68 B.n67 585
R578 B.n640 B.n68 585
R579 B.n638 B.n637 585
R580 B.n639 B.n638 585
R581 B.n636 B.n73 585
R582 B.n73 B.n72 585
R583 B.n635 B.n634 585
R584 B.n634 B.n633 585
R585 B.n75 B.n74 585
R586 B.n632 B.n75 585
R587 B.n630 B.n629 585
R588 B.n631 B.n630 585
R589 B.n628 B.n80 585
R590 B.n80 B.n79 585
R591 B.n627 B.n626 585
R592 B.n626 B.n625 585
R593 B.n82 B.n81 585
R594 B.n624 B.n82 585
R595 B.n622 B.n621 585
R596 B.n623 B.n622 585
R597 B.n620 B.n87 585
R598 B.n87 B.n86 585
R599 B.n619 B.n618 585
R600 B.n618 B.n617 585
R601 B.n89 B.n88 585
R602 B.n616 B.n89 585
R603 B.n614 B.n613 585
R604 B.n615 B.n614 585
R605 B.n612 B.n94 585
R606 B.n94 B.n93 585
R607 B.n611 B.n610 585
R608 B.n610 B.n609 585
R609 B.n715 B.n714 585
R610 B.n713 B.n2 585
R611 B.n610 B.n96 497.305
R612 B.n607 B.n97 497.305
R613 B.n381 B.n289 497.305
R614 B.n383 B.n287 497.305
R615 B.n608 B.n114 256.663
R616 B.n608 B.n113 256.663
R617 B.n608 B.n112 256.663
R618 B.n608 B.n111 256.663
R619 B.n608 B.n110 256.663
R620 B.n608 B.n109 256.663
R621 B.n608 B.n108 256.663
R622 B.n608 B.n107 256.663
R623 B.n608 B.n106 256.663
R624 B.n608 B.n105 256.663
R625 B.n608 B.n104 256.663
R626 B.n608 B.n103 256.663
R627 B.n608 B.n102 256.663
R628 B.n608 B.n101 256.663
R629 B.n608 B.n100 256.663
R630 B.n608 B.n99 256.663
R631 B.n608 B.n98 256.663
R632 B.n311 B.n288 256.663
R633 B.n317 B.n288 256.663
R634 B.n319 B.n288 256.663
R635 B.n325 B.n288 256.663
R636 B.n327 B.n288 256.663
R637 B.n333 B.n288 256.663
R638 B.n335 B.n288 256.663
R639 B.n341 B.n288 256.663
R640 B.n343 B.n288 256.663
R641 B.n349 B.n288 256.663
R642 B.n351 B.n288 256.663
R643 B.n358 B.n288 256.663
R644 B.n360 B.n288 256.663
R645 B.n366 B.n288 256.663
R646 B.n368 B.n288 256.663
R647 B.n374 B.n288 256.663
R648 B.n376 B.n288 256.663
R649 B.n717 B.n716 256.663
R650 B.n119 B.t14 224.629
R651 B.n116 B.t10 224.629
R652 B.n296 B.t17 224.629
R653 B.n302 B.t6 224.629
R654 B.n382 B.n288 165.845
R655 B.n609 B.n608 165.845
R656 B.n123 B.n122 163.367
R657 B.n127 B.n126 163.367
R658 B.n131 B.n130 163.367
R659 B.n135 B.n134 163.367
R660 B.n139 B.n138 163.367
R661 B.n143 B.n142 163.367
R662 B.n148 B.n147 163.367
R663 B.n152 B.n151 163.367
R664 B.n156 B.n155 163.367
R665 B.n160 B.n159 163.367
R666 B.n164 B.n163 163.367
R667 B.n168 B.n167 163.367
R668 B.n172 B.n171 163.367
R669 B.n176 B.n175 163.367
R670 B.n180 B.n179 163.367
R671 B.n184 B.n183 163.367
R672 B.n607 B.n115 163.367
R673 B.n381 B.n283 163.367
R674 B.n389 B.n283 163.367
R675 B.n389 B.n281 163.367
R676 B.n393 B.n281 163.367
R677 B.n393 B.n275 163.367
R678 B.n401 B.n275 163.367
R679 B.n401 B.n273 163.367
R680 B.n405 B.n273 163.367
R681 B.n405 B.n267 163.367
R682 B.n413 B.n267 163.367
R683 B.n413 B.n265 163.367
R684 B.n417 B.n265 163.367
R685 B.n417 B.n259 163.367
R686 B.n425 B.n259 163.367
R687 B.n425 B.n257 163.367
R688 B.n429 B.n257 163.367
R689 B.n429 B.n251 163.367
R690 B.n437 B.n251 163.367
R691 B.n437 B.n249 163.367
R692 B.n441 B.n249 163.367
R693 B.n441 B.n242 163.367
R694 B.n449 B.n242 163.367
R695 B.n449 B.n240 163.367
R696 B.n453 B.n240 163.367
R697 B.n453 B.n235 163.367
R698 B.n461 B.n235 163.367
R699 B.n461 B.n233 163.367
R700 B.n465 B.n233 163.367
R701 B.n465 B.n227 163.367
R702 B.n473 B.n227 163.367
R703 B.n473 B.n225 163.367
R704 B.n477 B.n225 163.367
R705 B.n477 B.n219 163.367
R706 B.n485 B.n219 163.367
R707 B.n485 B.n217 163.367
R708 B.n489 B.n217 163.367
R709 B.n489 B.n211 163.367
R710 B.n497 B.n211 163.367
R711 B.n497 B.n209 163.367
R712 B.n501 B.n209 163.367
R713 B.n501 B.n203 163.367
R714 B.n509 B.n203 163.367
R715 B.n509 B.n201 163.367
R716 B.n513 B.n201 163.367
R717 B.n513 B.n196 163.367
R718 B.n522 B.n196 163.367
R719 B.n522 B.n194 163.367
R720 B.n527 B.n194 163.367
R721 B.n527 B.n188 163.367
R722 B.n535 B.n188 163.367
R723 B.n536 B.n535 163.367
R724 B.n536 B.n5 163.367
R725 B.n6 B.n5 163.367
R726 B.n7 B.n6 163.367
R727 B.n542 B.n7 163.367
R728 B.n543 B.n542 163.367
R729 B.n543 B.n13 163.367
R730 B.n14 B.n13 163.367
R731 B.n15 B.n14 163.367
R732 B.n548 B.n15 163.367
R733 B.n548 B.n20 163.367
R734 B.n21 B.n20 163.367
R735 B.n22 B.n21 163.367
R736 B.n553 B.n22 163.367
R737 B.n553 B.n27 163.367
R738 B.n28 B.n27 163.367
R739 B.n29 B.n28 163.367
R740 B.n558 B.n29 163.367
R741 B.n558 B.n34 163.367
R742 B.n35 B.n34 163.367
R743 B.n36 B.n35 163.367
R744 B.n563 B.n36 163.367
R745 B.n563 B.n41 163.367
R746 B.n42 B.n41 163.367
R747 B.n43 B.n42 163.367
R748 B.n568 B.n43 163.367
R749 B.n568 B.n48 163.367
R750 B.n49 B.n48 163.367
R751 B.n50 B.n49 163.367
R752 B.n573 B.n50 163.367
R753 B.n573 B.n55 163.367
R754 B.n56 B.n55 163.367
R755 B.n57 B.n56 163.367
R756 B.n578 B.n57 163.367
R757 B.n578 B.n62 163.367
R758 B.n63 B.n62 163.367
R759 B.n64 B.n63 163.367
R760 B.n583 B.n64 163.367
R761 B.n583 B.n69 163.367
R762 B.n70 B.n69 163.367
R763 B.n71 B.n70 163.367
R764 B.n588 B.n71 163.367
R765 B.n588 B.n76 163.367
R766 B.n77 B.n76 163.367
R767 B.n78 B.n77 163.367
R768 B.n593 B.n78 163.367
R769 B.n593 B.n83 163.367
R770 B.n84 B.n83 163.367
R771 B.n85 B.n84 163.367
R772 B.n598 B.n85 163.367
R773 B.n598 B.n90 163.367
R774 B.n91 B.n90 163.367
R775 B.n92 B.n91 163.367
R776 B.n603 B.n92 163.367
R777 B.n603 B.n97 163.367
R778 B.n312 B.n310 163.367
R779 B.n316 B.n310 163.367
R780 B.n320 B.n318 163.367
R781 B.n324 B.n308 163.367
R782 B.n328 B.n326 163.367
R783 B.n332 B.n306 163.367
R784 B.n336 B.n334 163.367
R785 B.n340 B.n301 163.367
R786 B.n344 B.n342 163.367
R787 B.n348 B.n299 163.367
R788 B.n352 B.n350 163.367
R789 B.n357 B.n295 163.367
R790 B.n361 B.n359 163.367
R791 B.n365 B.n293 163.367
R792 B.n369 B.n367 163.367
R793 B.n373 B.n291 163.367
R794 B.n377 B.n375 163.367
R795 B.n383 B.n285 163.367
R796 B.n387 B.n285 163.367
R797 B.n387 B.n279 163.367
R798 B.n395 B.n279 163.367
R799 B.n395 B.n277 163.367
R800 B.n399 B.n277 163.367
R801 B.n399 B.n271 163.367
R802 B.n407 B.n271 163.367
R803 B.n407 B.n269 163.367
R804 B.n411 B.n269 163.367
R805 B.n411 B.n263 163.367
R806 B.n419 B.n263 163.367
R807 B.n419 B.n261 163.367
R808 B.n423 B.n261 163.367
R809 B.n423 B.n255 163.367
R810 B.n431 B.n255 163.367
R811 B.n431 B.n253 163.367
R812 B.n435 B.n253 163.367
R813 B.n435 B.n247 163.367
R814 B.n443 B.n247 163.367
R815 B.n443 B.n245 163.367
R816 B.n447 B.n245 163.367
R817 B.n447 B.n239 163.367
R818 B.n455 B.n239 163.367
R819 B.n455 B.n237 163.367
R820 B.n459 B.n237 163.367
R821 B.n459 B.n231 163.367
R822 B.n467 B.n231 163.367
R823 B.n467 B.n229 163.367
R824 B.n471 B.n229 163.367
R825 B.n471 B.n223 163.367
R826 B.n479 B.n223 163.367
R827 B.n479 B.n221 163.367
R828 B.n483 B.n221 163.367
R829 B.n483 B.n215 163.367
R830 B.n491 B.n215 163.367
R831 B.n491 B.n213 163.367
R832 B.n495 B.n213 163.367
R833 B.n495 B.n207 163.367
R834 B.n503 B.n207 163.367
R835 B.n503 B.n205 163.367
R836 B.n507 B.n205 163.367
R837 B.n507 B.n199 163.367
R838 B.n516 B.n199 163.367
R839 B.n516 B.n197 163.367
R840 B.n520 B.n197 163.367
R841 B.n520 B.n192 163.367
R842 B.n529 B.n192 163.367
R843 B.n529 B.n190 163.367
R844 B.n533 B.n190 163.367
R845 B.n533 B.n3 163.367
R846 B.n715 B.n3 163.367
R847 B.n711 B.n2 163.367
R848 B.n711 B.n710 163.367
R849 B.n710 B.n9 163.367
R850 B.n706 B.n9 163.367
R851 B.n706 B.n11 163.367
R852 B.n702 B.n11 163.367
R853 B.n702 B.n16 163.367
R854 B.n698 B.n16 163.367
R855 B.n698 B.n18 163.367
R856 B.n694 B.n18 163.367
R857 B.n694 B.n24 163.367
R858 B.n690 B.n24 163.367
R859 B.n690 B.n26 163.367
R860 B.n686 B.n26 163.367
R861 B.n686 B.n31 163.367
R862 B.n682 B.n31 163.367
R863 B.n682 B.n33 163.367
R864 B.n678 B.n33 163.367
R865 B.n678 B.n38 163.367
R866 B.n674 B.n38 163.367
R867 B.n674 B.n40 163.367
R868 B.n670 B.n40 163.367
R869 B.n670 B.n45 163.367
R870 B.n666 B.n45 163.367
R871 B.n666 B.n47 163.367
R872 B.n662 B.n47 163.367
R873 B.n662 B.n52 163.367
R874 B.n658 B.n52 163.367
R875 B.n658 B.n54 163.367
R876 B.n654 B.n54 163.367
R877 B.n654 B.n59 163.367
R878 B.n650 B.n59 163.367
R879 B.n650 B.n61 163.367
R880 B.n646 B.n61 163.367
R881 B.n646 B.n66 163.367
R882 B.n642 B.n66 163.367
R883 B.n642 B.n68 163.367
R884 B.n638 B.n68 163.367
R885 B.n638 B.n73 163.367
R886 B.n634 B.n73 163.367
R887 B.n634 B.n75 163.367
R888 B.n630 B.n75 163.367
R889 B.n630 B.n80 163.367
R890 B.n626 B.n80 163.367
R891 B.n626 B.n82 163.367
R892 B.n622 B.n82 163.367
R893 B.n622 B.n87 163.367
R894 B.n618 B.n87 163.367
R895 B.n618 B.n89 163.367
R896 B.n614 B.n89 163.367
R897 B.n614 B.n94 163.367
R898 B.n610 B.n94 163.367
R899 B.n116 B.t12 158.935
R900 B.n296 B.t19 158.935
R901 B.n119 B.t15 158.935
R902 B.n302 B.t9 158.935
R903 B.n382 B.n284 99.8004
R904 B.n388 B.n284 99.8004
R905 B.n388 B.n280 99.8004
R906 B.n394 B.n280 99.8004
R907 B.n394 B.n276 99.8004
R908 B.n400 B.n276 99.8004
R909 B.n400 B.n272 99.8004
R910 B.n406 B.n272 99.8004
R911 B.n412 B.n268 99.8004
R912 B.n412 B.n264 99.8004
R913 B.n418 B.n264 99.8004
R914 B.n418 B.n260 99.8004
R915 B.n424 B.n260 99.8004
R916 B.n424 B.n256 99.8004
R917 B.n430 B.n256 99.8004
R918 B.n430 B.n252 99.8004
R919 B.n436 B.n252 99.8004
R920 B.n436 B.n248 99.8004
R921 B.n442 B.n248 99.8004
R922 B.n442 B.n243 99.8004
R923 B.n448 B.n243 99.8004
R924 B.n448 B.n244 99.8004
R925 B.n454 B.n236 99.8004
R926 B.n460 B.n236 99.8004
R927 B.n460 B.n232 99.8004
R928 B.n466 B.n232 99.8004
R929 B.n466 B.n228 99.8004
R930 B.n472 B.n228 99.8004
R931 B.n472 B.n224 99.8004
R932 B.n478 B.n224 99.8004
R933 B.n478 B.n220 99.8004
R934 B.n484 B.n220 99.8004
R935 B.n490 B.n216 99.8004
R936 B.n490 B.n212 99.8004
R937 B.n496 B.n212 99.8004
R938 B.n496 B.n208 99.8004
R939 B.n502 B.n208 99.8004
R940 B.n502 B.n204 99.8004
R941 B.n508 B.n204 99.8004
R942 B.n508 B.n200 99.8004
R943 B.n515 B.n200 99.8004
R944 B.n515 B.n514 99.8004
R945 B.n521 B.n193 99.8004
R946 B.n528 B.n193 99.8004
R947 B.n528 B.n189 99.8004
R948 B.n534 B.n189 99.8004
R949 B.n534 B.n4 99.8004
R950 B.n714 B.n4 99.8004
R951 B.n714 B.n713 99.8004
R952 B.n713 B.n712 99.8004
R953 B.n712 B.n8 99.8004
R954 B.n12 B.n8 99.8004
R955 B.n705 B.n12 99.8004
R956 B.n705 B.n704 99.8004
R957 B.n704 B.n703 99.8004
R958 B.n697 B.n19 99.8004
R959 B.n697 B.n696 99.8004
R960 B.n696 B.n695 99.8004
R961 B.n695 B.n23 99.8004
R962 B.n689 B.n23 99.8004
R963 B.n689 B.n688 99.8004
R964 B.n688 B.n687 99.8004
R965 B.n687 B.n30 99.8004
R966 B.n681 B.n30 99.8004
R967 B.n681 B.n680 99.8004
R968 B.n679 B.n37 99.8004
R969 B.n673 B.n37 99.8004
R970 B.n673 B.n672 99.8004
R971 B.n672 B.n671 99.8004
R972 B.n671 B.n44 99.8004
R973 B.n665 B.n44 99.8004
R974 B.n665 B.n664 99.8004
R975 B.n664 B.n663 99.8004
R976 B.n663 B.n51 99.8004
R977 B.n657 B.n51 99.8004
R978 B.n656 B.n655 99.8004
R979 B.n655 B.n58 99.8004
R980 B.n649 B.n58 99.8004
R981 B.n649 B.n648 99.8004
R982 B.n648 B.n647 99.8004
R983 B.n647 B.n65 99.8004
R984 B.n641 B.n65 99.8004
R985 B.n641 B.n640 99.8004
R986 B.n640 B.n639 99.8004
R987 B.n639 B.n72 99.8004
R988 B.n633 B.n72 99.8004
R989 B.n633 B.n632 99.8004
R990 B.n632 B.n631 99.8004
R991 B.n631 B.n79 99.8004
R992 B.n625 B.n624 99.8004
R993 B.n624 B.n623 99.8004
R994 B.n623 B.n86 99.8004
R995 B.n617 B.n86 99.8004
R996 B.n617 B.n616 99.8004
R997 B.n616 B.n615 99.8004
R998 B.n615 B.n93 99.8004
R999 B.n609 B.n93 99.8004
R1000 B.n406 B.t7 98.3327
R1001 B.n625 B.t11 98.3327
R1002 B.n117 B.t13 86.0146
R1003 B.n297 B.t18 86.0146
R1004 B.n120 B.t16 86.0143
R1005 B.n303 B.t8 86.0143
R1006 B.n454 B.t3 74.8504
R1007 B.n657 B.t4 74.8504
R1008 B.n120 B.n119 72.9217
R1009 B.n117 B.n116 72.9217
R1010 B.n297 B.n296 72.9217
R1011 B.n303 B.n302 72.9217
R1012 B.n98 B.n96 71.676
R1013 B.n123 B.n99 71.676
R1014 B.n127 B.n100 71.676
R1015 B.n131 B.n101 71.676
R1016 B.n135 B.n102 71.676
R1017 B.n139 B.n103 71.676
R1018 B.n143 B.n104 71.676
R1019 B.n148 B.n105 71.676
R1020 B.n152 B.n106 71.676
R1021 B.n156 B.n107 71.676
R1022 B.n160 B.n108 71.676
R1023 B.n164 B.n109 71.676
R1024 B.n168 B.n110 71.676
R1025 B.n172 B.n111 71.676
R1026 B.n176 B.n112 71.676
R1027 B.n180 B.n113 71.676
R1028 B.n184 B.n114 71.676
R1029 B.n115 B.n114 71.676
R1030 B.n183 B.n113 71.676
R1031 B.n179 B.n112 71.676
R1032 B.n175 B.n111 71.676
R1033 B.n171 B.n110 71.676
R1034 B.n167 B.n109 71.676
R1035 B.n163 B.n108 71.676
R1036 B.n159 B.n107 71.676
R1037 B.n155 B.n106 71.676
R1038 B.n151 B.n105 71.676
R1039 B.n147 B.n104 71.676
R1040 B.n142 B.n103 71.676
R1041 B.n138 B.n102 71.676
R1042 B.n134 B.n101 71.676
R1043 B.n130 B.n100 71.676
R1044 B.n126 B.n99 71.676
R1045 B.n122 B.n98 71.676
R1046 B.n311 B.n287 71.676
R1047 B.n317 B.n316 71.676
R1048 B.n320 B.n319 71.676
R1049 B.n325 B.n324 71.676
R1050 B.n328 B.n327 71.676
R1051 B.n333 B.n332 71.676
R1052 B.n336 B.n335 71.676
R1053 B.n341 B.n340 71.676
R1054 B.n344 B.n343 71.676
R1055 B.n349 B.n348 71.676
R1056 B.n352 B.n351 71.676
R1057 B.n358 B.n357 71.676
R1058 B.n361 B.n360 71.676
R1059 B.n366 B.n365 71.676
R1060 B.n369 B.n368 71.676
R1061 B.n374 B.n373 71.676
R1062 B.n377 B.n376 71.676
R1063 B.n312 B.n311 71.676
R1064 B.n318 B.n317 71.676
R1065 B.n319 B.n308 71.676
R1066 B.n326 B.n325 71.676
R1067 B.n327 B.n306 71.676
R1068 B.n334 B.n333 71.676
R1069 B.n335 B.n301 71.676
R1070 B.n342 B.n341 71.676
R1071 B.n343 B.n299 71.676
R1072 B.n350 B.n349 71.676
R1073 B.n351 B.n295 71.676
R1074 B.n359 B.n358 71.676
R1075 B.n360 B.n293 71.676
R1076 B.n367 B.n366 71.676
R1077 B.n368 B.n291 71.676
R1078 B.n375 B.n374 71.676
R1079 B.n376 B.n289 71.676
R1080 B.n716 B.n715 71.676
R1081 B.n716 B.n2 71.676
R1082 B.t2 B.n216 68.9798
R1083 B.n680 B.t0 68.9798
R1084 B.n521 B.t5 63.1092
R1085 B.n703 B.t1 63.1092
R1086 B.n145 B.n120 59.5399
R1087 B.n118 B.n117 59.5399
R1088 B.n354 B.n297 59.5399
R1089 B.n304 B.n303 59.5399
R1090 B.n514 B.t5 36.6916
R1091 B.n19 B.t1 36.6916
R1092 B.n384 B.n286 32.3127
R1093 B.n380 B.n379 32.3127
R1094 B.n606 B.n605 32.3127
R1095 B.n611 B.n95 32.3127
R1096 B.n484 B.t2 30.821
R1097 B.t0 B.n679 30.821
R1098 B.n244 B.t3 24.9505
R1099 B.t4 B.n656 24.9505
R1100 B B.n717 18.0485
R1101 B.n385 B.n384 10.6151
R1102 B.n386 B.n385 10.6151
R1103 B.n386 B.n278 10.6151
R1104 B.n396 B.n278 10.6151
R1105 B.n397 B.n396 10.6151
R1106 B.n398 B.n397 10.6151
R1107 B.n398 B.n270 10.6151
R1108 B.n408 B.n270 10.6151
R1109 B.n409 B.n408 10.6151
R1110 B.n410 B.n409 10.6151
R1111 B.n410 B.n262 10.6151
R1112 B.n420 B.n262 10.6151
R1113 B.n421 B.n420 10.6151
R1114 B.n422 B.n421 10.6151
R1115 B.n422 B.n254 10.6151
R1116 B.n432 B.n254 10.6151
R1117 B.n433 B.n432 10.6151
R1118 B.n434 B.n433 10.6151
R1119 B.n434 B.n246 10.6151
R1120 B.n444 B.n246 10.6151
R1121 B.n445 B.n444 10.6151
R1122 B.n446 B.n445 10.6151
R1123 B.n446 B.n238 10.6151
R1124 B.n456 B.n238 10.6151
R1125 B.n457 B.n456 10.6151
R1126 B.n458 B.n457 10.6151
R1127 B.n458 B.n230 10.6151
R1128 B.n468 B.n230 10.6151
R1129 B.n469 B.n468 10.6151
R1130 B.n470 B.n469 10.6151
R1131 B.n470 B.n222 10.6151
R1132 B.n480 B.n222 10.6151
R1133 B.n481 B.n480 10.6151
R1134 B.n482 B.n481 10.6151
R1135 B.n482 B.n214 10.6151
R1136 B.n492 B.n214 10.6151
R1137 B.n493 B.n492 10.6151
R1138 B.n494 B.n493 10.6151
R1139 B.n494 B.n206 10.6151
R1140 B.n504 B.n206 10.6151
R1141 B.n505 B.n504 10.6151
R1142 B.n506 B.n505 10.6151
R1143 B.n506 B.n198 10.6151
R1144 B.n517 B.n198 10.6151
R1145 B.n518 B.n517 10.6151
R1146 B.n519 B.n518 10.6151
R1147 B.n519 B.n191 10.6151
R1148 B.n530 B.n191 10.6151
R1149 B.n531 B.n530 10.6151
R1150 B.n532 B.n531 10.6151
R1151 B.n532 B.n0 10.6151
R1152 B.n313 B.n286 10.6151
R1153 B.n314 B.n313 10.6151
R1154 B.n315 B.n314 10.6151
R1155 B.n315 B.n309 10.6151
R1156 B.n321 B.n309 10.6151
R1157 B.n322 B.n321 10.6151
R1158 B.n323 B.n322 10.6151
R1159 B.n323 B.n307 10.6151
R1160 B.n329 B.n307 10.6151
R1161 B.n330 B.n329 10.6151
R1162 B.n331 B.n330 10.6151
R1163 B.n331 B.n305 10.6151
R1164 B.n338 B.n337 10.6151
R1165 B.n339 B.n338 10.6151
R1166 B.n339 B.n300 10.6151
R1167 B.n345 B.n300 10.6151
R1168 B.n346 B.n345 10.6151
R1169 B.n347 B.n346 10.6151
R1170 B.n347 B.n298 10.6151
R1171 B.n353 B.n298 10.6151
R1172 B.n356 B.n355 10.6151
R1173 B.n356 B.n294 10.6151
R1174 B.n362 B.n294 10.6151
R1175 B.n363 B.n362 10.6151
R1176 B.n364 B.n363 10.6151
R1177 B.n364 B.n292 10.6151
R1178 B.n370 B.n292 10.6151
R1179 B.n371 B.n370 10.6151
R1180 B.n372 B.n371 10.6151
R1181 B.n372 B.n290 10.6151
R1182 B.n378 B.n290 10.6151
R1183 B.n379 B.n378 10.6151
R1184 B.n380 B.n282 10.6151
R1185 B.n390 B.n282 10.6151
R1186 B.n391 B.n390 10.6151
R1187 B.n392 B.n391 10.6151
R1188 B.n392 B.n274 10.6151
R1189 B.n402 B.n274 10.6151
R1190 B.n403 B.n402 10.6151
R1191 B.n404 B.n403 10.6151
R1192 B.n404 B.n266 10.6151
R1193 B.n414 B.n266 10.6151
R1194 B.n415 B.n414 10.6151
R1195 B.n416 B.n415 10.6151
R1196 B.n416 B.n258 10.6151
R1197 B.n426 B.n258 10.6151
R1198 B.n427 B.n426 10.6151
R1199 B.n428 B.n427 10.6151
R1200 B.n428 B.n250 10.6151
R1201 B.n438 B.n250 10.6151
R1202 B.n439 B.n438 10.6151
R1203 B.n440 B.n439 10.6151
R1204 B.n440 B.n241 10.6151
R1205 B.n450 B.n241 10.6151
R1206 B.n451 B.n450 10.6151
R1207 B.n452 B.n451 10.6151
R1208 B.n452 B.n234 10.6151
R1209 B.n462 B.n234 10.6151
R1210 B.n463 B.n462 10.6151
R1211 B.n464 B.n463 10.6151
R1212 B.n464 B.n226 10.6151
R1213 B.n474 B.n226 10.6151
R1214 B.n475 B.n474 10.6151
R1215 B.n476 B.n475 10.6151
R1216 B.n476 B.n218 10.6151
R1217 B.n486 B.n218 10.6151
R1218 B.n487 B.n486 10.6151
R1219 B.n488 B.n487 10.6151
R1220 B.n488 B.n210 10.6151
R1221 B.n498 B.n210 10.6151
R1222 B.n499 B.n498 10.6151
R1223 B.n500 B.n499 10.6151
R1224 B.n500 B.n202 10.6151
R1225 B.n510 B.n202 10.6151
R1226 B.n511 B.n510 10.6151
R1227 B.n512 B.n511 10.6151
R1228 B.n512 B.n195 10.6151
R1229 B.n523 B.n195 10.6151
R1230 B.n524 B.n523 10.6151
R1231 B.n526 B.n524 10.6151
R1232 B.n526 B.n525 10.6151
R1233 B.n525 B.n187 10.6151
R1234 B.n537 B.n187 10.6151
R1235 B.n538 B.n537 10.6151
R1236 B.n539 B.n538 10.6151
R1237 B.n540 B.n539 10.6151
R1238 B.n541 B.n540 10.6151
R1239 B.n544 B.n541 10.6151
R1240 B.n545 B.n544 10.6151
R1241 B.n546 B.n545 10.6151
R1242 B.n547 B.n546 10.6151
R1243 B.n549 B.n547 10.6151
R1244 B.n550 B.n549 10.6151
R1245 B.n551 B.n550 10.6151
R1246 B.n552 B.n551 10.6151
R1247 B.n554 B.n552 10.6151
R1248 B.n555 B.n554 10.6151
R1249 B.n556 B.n555 10.6151
R1250 B.n557 B.n556 10.6151
R1251 B.n559 B.n557 10.6151
R1252 B.n560 B.n559 10.6151
R1253 B.n561 B.n560 10.6151
R1254 B.n562 B.n561 10.6151
R1255 B.n564 B.n562 10.6151
R1256 B.n565 B.n564 10.6151
R1257 B.n566 B.n565 10.6151
R1258 B.n567 B.n566 10.6151
R1259 B.n569 B.n567 10.6151
R1260 B.n570 B.n569 10.6151
R1261 B.n571 B.n570 10.6151
R1262 B.n572 B.n571 10.6151
R1263 B.n574 B.n572 10.6151
R1264 B.n575 B.n574 10.6151
R1265 B.n576 B.n575 10.6151
R1266 B.n577 B.n576 10.6151
R1267 B.n579 B.n577 10.6151
R1268 B.n580 B.n579 10.6151
R1269 B.n581 B.n580 10.6151
R1270 B.n582 B.n581 10.6151
R1271 B.n584 B.n582 10.6151
R1272 B.n585 B.n584 10.6151
R1273 B.n586 B.n585 10.6151
R1274 B.n587 B.n586 10.6151
R1275 B.n589 B.n587 10.6151
R1276 B.n590 B.n589 10.6151
R1277 B.n591 B.n590 10.6151
R1278 B.n592 B.n591 10.6151
R1279 B.n594 B.n592 10.6151
R1280 B.n595 B.n594 10.6151
R1281 B.n596 B.n595 10.6151
R1282 B.n597 B.n596 10.6151
R1283 B.n599 B.n597 10.6151
R1284 B.n600 B.n599 10.6151
R1285 B.n601 B.n600 10.6151
R1286 B.n602 B.n601 10.6151
R1287 B.n604 B.n602 10.6151
R1288 B.n605 B.n604 10.6151
R1289 B.n709 B.n1 10.6151
R1290 B.n709 B.n708 10.6151
R1291 B.n708 B.n707 10.6151
R1292 B.n707 B.n10 10.6151
R1293 B.n701 B.n10 10.6151
R1294 B.n701 B.n700 10.6151
R1295 B.n700 B.n699 10.6151
R1296 B.n699 B.n17 10.6151
R1297 B.n693 B.n17 10.6151
R1298 B.n693 B.n692 10.6151
R1299 B.n692 B.n691 10.6151
R1300 B.n691 B.n25 10.6151
R1301 B.n685 B.n25 10.6151
R1302 B.n685 B.n684 10.6151
R1303 B.n684 B.n683 10.6151
R1304 B.n683 B.n32 10.6151
R1305 B.n677 B.n32 10.6151
R1306 B.n677 B.n676 10.6151
R1307 B.n676 B.n675 10.6151
R1308 B.n675 B.n39 10.6151
R1309 B.n669 B.n39 10.6151
R1310 B.n669 B.n668 10.6151
R1311 B.n668 B.n667 10.6151
R1312 B.n667 B.n46 10.6151
R1313 B.n661 B.n46 10.6151
R1314 B.n661 B.n660 10.6151
R1315 B.n660 B.n659 10.6151
R1316 B.n659 B.n53 10.6151
R1317 B.n653 B.n53 10.6151
R1318 B.n653 B.n652 10.6151
R1319 B.n652 B.n651 10.6151
R1320 B.n651 B.n60 10.6151
R1321 B.n645 B.n60 10.6151
R1322 B.n645 B.n644 10.6151
R1323 B.n644 B.n643 10.6151
R1324 B.n643 B.n67 10.6151
R1325 B.n637 B.n67 10.6151
R1326 B.n637 B.n636 10.6151
R1327 B.n636 B.n635 10.6151
R1328 B.n635 B.n74 10.6151
R1329 B.n629 B.n74 10.6151
R1330 B.n629 B.n628 10.6151
R1331 B.n628 B.n627 10.6151
R1332 B.n627 B.n81 10.6151
R1333 B.n621 B.n81 10.6151
R1334 B.n621 B.n620 10.6151
R1335 B.n620 B.n619 10.6151
R1336 B.n619 B.n88 10.6151
R1337 B.n613 B.n88 10.6151
R1338 B.n613 B.n612 10.6151
R1339 B.n612 B.n611 10.6151
R1340 B.n121 B.n95 10.6151
R1341 B.n124 B.n121 10.6151
R1342 B.n125 B.n124 10.6151
R1343 B.n128 B.n125 10.6151
R1344 B.n129 B.n128 10.6151
R1345 B.n132 B.n129 10.6151
R1346 B.n133 B.n132 10.6151
R1347 B.n136 B.n133 10.6151
R1348 B.n137 B.n136 10.6151
R1349 B.n140 B.n137 10.6151
R1350 B.n141 B.n140 10.6151
R1351 B.n144 B.n141 10.6151
R1352 B.n149 B.n146 10.6151
R1353 B.n150 B.n149 10.6151
R1354 B.n153 B.n150 10.6151
R1355 B.n154 B.n153 10.6151
R1356 B.n157 B.n154 10.6151
R1357 B.n158 B.n157 10.6151
R1358 B.n161 B.n158 10.6151
R1359 B.n162 B.n161 10.6151
R1360 B.n166 B.n165 10.6151
R1361 B.n169 B.n166 10.6151
R1362 B.n170 B.n169 10.6151
R1363 B.n173 B.n170 10.6151
R1364 B.n174 B.n173 10.6151
R1365 B.n177 B.n174 10.6151
R1366 B.n178 B.n177 10.6151
R1367 B.n181 B.n178 10.6151
R1368 B.n182 B.n181 10.6151
R1369 B.n185 B.n182 10.6151
R1370 B.n186 B.n185 10.6151
R1371 B.n606 B.n186 10.6151
R1372 B.n717 B.n0 8.11757
R1373 B.n717 B.n1 8.11757
R1374 B.n337 B.n304 6.5566
R1375 B.n354 B.n353 6.5566
R1376 B.n146 B.n145 6.5566
R1377 B.n162 B.n118 6.5566
R1378 B.n305 B.n304 4.05904
R1379 B.n355 B.n354 4.05904
R1380 B.n145 B.n144 4.05904
R1381 B.n165 B.n118 4.05904
R1382 B.t7 B.n268 1.46815
R1383 B.t11 B.n79 1.46815
R1384 VN.n34 VN.n33 161.3
R1385 VN.n32 VN.n19 161.3
R1386 VN.n31 VN.n30 161.3
R1387 VN.n29 VN.n20 161.3
R1388 VN.n28 VN.n27 161.3
R1389 VN.n26 VN.n21 161.3
R1390 VN.n25 VN.n24 161.3
R1391 VN.n16 VN.n15 161.3
R1392 VN.n14 VN.n1 161.3
R1393 VN.n13 VN.n12 161.3
R1394 VN.n11 VN.n2 161.3
R1395 VN.n10 VN.n9 161.3
R1396 VN.n8 VN.n3 161.3
R1397 VN.n7 VN.n6 161.3
R1398 VN.n17 VN.n0 77.2324
R1399 VN.n35 VN.n18 77.2324
R1400 VN.n9 VN.n2 52.0954
R1401 VN.n27 VN.n20 52.0954
R1402 VN.n5 VN.n4 50.0561
R1403 VN.n23 VN.n22 50.0561
R1404 VN.n5 VN.t3 49.3623
R1405 VN.n23 VN.t2 49.3623
R1406 VN VN.n35 44.8009
R1407 VN.n13 VN.n2 28.7258
R1408 VN.n31 VN.n20 28.7258
R1409 VN.n7 VN.n4 24.3439
R1410 VN.n8 VN.n7 24.3439
R1411 VN.n9 VN.n8 24.3439
R1412 VN.n14 VN.n13 24.3439
R1413 VN.n15 VN.n14 24.3439
R1414 VN.n27 VN.n26 24.3439
R1415 VN.n26 VN.n25 24.3439
R1416 VN.n25 VN.n22 24.3439
R1417 VN.n33 VN.n32 24.3439
R1418 VN.n32 VN.n31 24.3439
R1419 VN.n4 VN.t5 15.5988
R1420 VN.n0 VN.t1 15.5988
R1421 VN.n22 VN.t0 15.5988
R1422 VN.n18 VN.t4 15.5988
R1423 VN.n15 VN.n0 12.6591
R1424 VN.n33 VN.n18 12.6591
R1425 VN.n6 VN.n5 3.07273
R1426 VN.n24 VN.n23 3.07273
R1427 VN.n35 VN.n34 0.355081
R1428 VN.n17 VN.n16 0.355081
R1429 VN VN.n17 0.26685
R1430 VN.n34 VN.n19 0.189894
R1431 VN.n30 VN.n19 0.189894
R1432 VN.n30 VN.n29 0.189894
R1433 VN.n29 VN.n28 0.189894
R1434 VN.n28 VN.n21 0.189894
R1435 VN.n24 VN.n21 0.189894
R1436 VN.n6 VN.n3 0.189894
R1437 VN.n10 VN.n3 0.189894
R1438 VN.n11 VN.n10 0.189894
R1439 VN.n12 VN.n11 0.189894
R1440 VN.n12 VN.n1 0.189894
R1441 VN.n16 VN.n1 0.189894
R1442 VDD2.n1 VDD2.t2 105.537
R1443 VDD2.n2 VDD2.t1 103.162
R1444 VDD2.n1 VDD2.n0 94.9982
R1445 VDD2 VDD2.n3 94.9955
R1446 VDD2.n2 VDD2.n1 36.1636
R1447 VDD2.n3 VDD2.t5 8.91942
R1448 VDD2.n3 VDD2.t3 8.91942
R1449 VDD2.n0 VDD2.t0 8.91942
R1450 VDD2.n0 VDD2.t4 8.91942
R1451 VDD2 VDD2.n2 2.48972
C0 VN VP 5.93566f
C1 VP VTAIL 2.75737f
C2 VDD1 VDD2 1.72996f
C3 VP VDD2 0.534891f
C4 VN VTAIL 2.74324f
C5 VP VDD1 2.00668f
C6 VN VDD2 1.63242f
C7 VDD2 VTAIL 4.83293f
C8 VN VDD1 0.157606f
C9 VDD1 VTAIL 4.77411f
C10 VDD2 B 4.699908f
C11 VDD1 B 5.230542f
C12 VTAIL B 3.910561f
C13 VN B 14.371289f
C14 VP B 13.103121f
C15 VDD2.t2 B 0.266065f
C16 VDD2.t0 B 0.029515f
C17 VDD2.t4 B 0.029515f
C18 VDD2.n0 B 0.203809f
C19 VDD2.n1 B 1.75218f
C20 VDD2.t1 B 0.259761f
C21 VDD2.n2 B 1.47749f
C22 VDD2.t5 B 0.029515f
C23 VDD2.t3 B 0.029515f
C24 VDD2.n3 B 0.203793f
C25 VN.t1 B 0.429912f
C26 VN.n0 B 0.28483f
C27 VN.n1 B 0.023705f
C28 VN.n2 B 0.024003f
C29 VN.n3 B 0.023705f
C30 VN.t5 B 0.429912f
C31 VN.n4 B 0.285077f
C32 VN.t3 B 0.68254f
C33 VN.n5 B 0.289696f
C34 VN.n6 B 0.289754f
C35 VN.n7 B 0.044403f
C36 VN.n8 B 0.044403f
C37 VN.n9 B 0.042768f
C38 VN.n10 B 0.023705f
C39 VN.n11 B 0.023705f
C40 VN.n12 B 0.023705f
C41 VN.n13 B 0.047145f
C42 VN.n14 B 0.044403f
C43 VN.n15 B 0.033879f
C44 VN.n16 B 0.038266f
C45 VN.n17 B 0.060572f
C46 VN.t4 B 0.429912f
C47 VN.n18 B 0.28483f
C48 VN.n19 B 0.023705f
C49 VN.n20 B 0.024003f
C50 VN.n21 B 0.023705f
C51 VN.t0 B 0.429912f
C52 VN.n22 B 0.285077f
C53 VN.t2 B 0.68254f
C54 VN.n23 B 0.289696f
C55 VN.n24 B 0.289754f
C56 VN.n25 B 0.044403f
C57 VN.n26 B 0.044403f
C58 VN.n27 B 0.042768f
C59 VN.n28 B 0.023705f
C60 VN.n29 B 0.023705f
C61 VN.n30 B 0.023705f
C62 VN.n31 B 0.047145f
C63 VN.n32 B 0.044403f
C64 VN.n33 B 0.033879f
C65 VN.n34 B 0.038266f
C66 VN.n35 B 1.1544f
C67 VDD1.t5 B 0.372719f
C68 VDD1.t2 B 0.372108f
C69 VDD1.t3 B 0.041278f
C70 VDD1.t4 B 0.041278f
C71 VDD1.n0 B 0.285039f
C72 VDD1.n1 B 2.57704f
C73 VDD1.t0 B 0.041278f
C74 VDD1.t1 B 0.041278f
C75 VDD1.n2 B 0.281186f
C76 VDD1.n3 B 2.11033f
C77 VTAIL.t1 B 0.06184f
C78 VTAIL.t0 B 0.06184f
C79 VTAIL.n0 B 0.367462f
C80 VTAIL.n1 B 0.598843f
C81 VTAIL.t10 B 0.487204f
C82 VTAIL.n2 B 0.917274f
C83 VTAIL.t11 B 0.06184f
C84 VTAIL.t6 B 0.06184f
C85 VTAIL.n3 B 0.367462f
C86 VTAIL.n4 B 2.06347f
C87 VTAIL.t3 B 0.06184f
C88 VTAIL.t2 B 0.06184f
C89 VTAIL.n5 B 0.367463f
C90 VTAIL.n6 B 2.06346f
C91 VTAIL.t5 B 0.487207f
C92 VTAIL.n7 B 0.917272f
C93 VTAIL.t7 B 0.06184f
C94 VTAIL.t9 B 0.06184f
C95 VTAIL.n8 B 0.367463f
C96 VTAIL.n9 B 0.86836f
C97 VTAIL.t8 B 0.487204f
C98 VTAIL.n10 B 1.74421f
C99 VTAIL.t4 B 0.487204f
C100 VTAIL.n11 B 1.64555f
C101 VP.t1 B 0.536971f
C102 VP.n0 B 0.35576f
C103 VP.n1 B 0.029609f
C104 VP.n2 B 0.02998f
C105 VP.n3 B 0.029609f
C106 VP.t2 B 0.536971f
C107 VP.n4 B 0.266074f
C108 VP.n5 B 0.029609f
C109 VP.n6 B 0.02998f
C110 VP.n7 B 0.029609f
C111 VP.t3 B 0.536971f
C112 VP.n8 B 0.35576f
C113 VP.t4 B 0.536971f
C114 VP.n9 B 0.35576f
C115 VP.n10 B 0.029609f
C116 VP.n11 B 0.02998f
C117 VP.n12 B 0.029609f
C118 VP.t5 B 0.536971f
C119 VP.n13 B 0.356069f
C120 VP.t0 B 0.852509f
C121 VP.n14 B 0.361838f
C122 VP.n15 B 0.361911f
C123 VP.n16 B 0.05546f
C124 VP.n17 B 0.05546f
C125 VP.n18 B 0.053418f
C126 VP.n19 B 0.029609f
C127 VP.n20 B 0.029609f
C128 VP.n21 B 0.029609f
C129 VP.n22 B 0.058885f
C130 VP.n23 B 0.05546f
C131 VP.n24 B 0.042316f
C132 VP.n25 B 0.047796f
C133 VP.n26 B 1.42926f
C134 VP.n27 B 1.45304f
C135 VP.n28 B 0.047796f
C136 VP.n29 B 0.042316f
C137 VP.n30 B 0.05546f
C138 VP.n31 B 0.058885f
C139 VP.n32 B 0.029609f
C140 VP.n33 B 0.029609f
C141 VP.n34 B 0.029609f
C142 VP.n35 B 0.053418f
C143 VP.n36 B 0.05546f
C144 VP.n37 B 0.05546f
C145 VP.n38 B 0.029609f
C146 VP.n39 B 0.029609f
C147 VP.n40 B 0.029609f
C148 VP.n41 B 0.05546f
C149 VP.n42 B 0.05546f
C150 VP.n43 B 0.053418f
C151 VP.n44 B 0.029609f
C152 VP.n45 B 0.029609f
C153 VP.n46 B 0.029609f
C154 VP.n47 B 0.058885f
C155 VP.n48 B 0.05546f
C156 VP.n49 B 0.042316f
C157 VP.n50 B 0.047796f
C158 VP.n51 B 0.075656f
.ends

