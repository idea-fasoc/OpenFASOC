* NGSPICE file created from diff_pair_sample_0340.ext - technology: sky130A

.subckt diff_pair_sample_0340 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=1.10055 ps=7 w=6.67 l=1.73
X1 VDD1.t9 VP.t0 VTAIL.t2 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X2 VTAIL.t17 VN.t1 VDD2.t8 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X3 B.t11 B.t9 B.t10 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=0 ps=0 w=6.67 l=1.73
X4 VDD2.t7 VN.t2 VTAIL.t19 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X5 VTAIL.t14 VN.t3 VDD2.t6 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X6 VDD1.t8 VP.t1 VTAIL.t0 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=1.10055 ps=7 w=6.67 l=1.73
X7 VTAIL.t1 VP.t2 VDD1.t7 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X8 VTAIL.t7 VP.t3 VDD1.t6 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X9 VTAIL.t15 VN.t4 VDD2.t5 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X10 VTAIL.t4 VP.t4 VDD1.t5 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X11 B.t8 B.t6 B.t7 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=0 ps=0 w=6.67 l=1.73
X12 VDD1.t4 VP.t5 VTAIL.t3 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X13 VDD2.t4 VN.t5 VTAIL.t11 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=2.6013 ps=14.12 w=6.67 l=1.73
X14 VDD2.t3 VN.t6 VTAIL.t12 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X15 VDD1.t3 VP.t6 VTAIL.t8 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=1.10055 ps=7 w=6.67 l=1.73
X16 VDD1.t2 VP.t7 VTAIL.t6 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=2.6013 ps=14.12 w=6.67 l=1.73
X17 B.t5 B.t3 B.t4 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=0 ps=0 w=6.67 l=1.73
X18 VTAIL.t10 VN.t7 VDD2.t2 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X19 B.t2 B.t0 B.t1 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=0 ps=0 w=6.67 l=1.73
X20 VTAIL.t5 VP.t8 VDD1.t1 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=1.10055 ps=7 w=6.67 l=1.73
X21 VDD2.t1 VN.t8 VTAIL.t16 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=2.6013 pd=14.12 as=1.10055 ps=7 w=6.67 l=1.73
X22 VDD2.t0 VN.t9 VTAIL.t13 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=2.6013 ps=14.12 w=6.67 l=1.73
X23 VDD1.t0 VP.t9 VTAIL.t9 w_n3442_n2302# sky130_fd_pr__pfet_01v8 ad=1.10055 pd=7 as=2.6013 ps=14.12 w=6.67 l=1.73
R0 VN.n30 VN.n29 179.895
R1 VN.n61 VN.n60 179.895
R2 VN.n59 VN.n31 161.3
R3 VN.n58 VN.n57 161.3
R4 VN.n56 VN.n32 161.3
R5 VN.n55 VN.n54 161.3
R6 VN.n52 VN.n33 161.3
R7 VN.n51 VN.n50 161.3
R8 VN.n49 VN.n34 161.3
R9 VN.n48 VN.n47 161.3
R10 VN.n46 VN.n35 161.3
R11 VN.n45 VN.n44 161.3
R12 VN.n43 VN.n36 161.3
R13 VN.n42 VN.n41 161.3
R14 VN.n40 VN.n37 161.3
R15 VN.n28 VN.n0 161.3
R16 VN.n27 VN.n26 161.3
R17 VN.n25 VN.n1 161.3
R18 VN.n24 VN.n23 161.3
R19 VN.n21 VN.n2 161.3
R20 VN.n20 VN.n19 161.3
R21 VN.n18 VN.n3 161.3
R22 VN.n17 VN.n16 161.3
R23 VN.n15 VN.n4 161.3
R24 VN.n14 VN.n13 161.3
R25 VN.n12 VN.n5 161.3
R26 VN.n11 VN.n10 161.3
R27 VN.n9 VN.n6 161.3
R28 VN.n7 VN.t8 123.969
R29 VN.n38 VN.t5 123.969
R30 VN.n15 VN.t6 92.9178
R31 VN.n8 VN.t7 92.9178
R32 VN.n22 VN.t1 92.9178
R33 VN.n29 VN.t9 92.9178
R34 VN.n46 VN.t2 92.9178
R35 VN.n39 VN.t4 92.9178
R36 VN.n53 VN.t3 92.9178
R37 VN.n60 VN.t0 92.9178
R38 VN.n8 VN.n7 64.8059
R39 VN.n39 VN.n38 64.8059
R40 VN.n27 VN.n1 49.2348
R41 VN.n58 VN.n32 49.2348
R42 VN VN.n61 44.6463
R43 VN.n10 VN.n5 43.4072
R44 VN.n20 VN.n3 43.4072
R45 VN.n41 VN.n36 43.4072
R46 VN.n51 VN.n34 43.4072
R47 VN.n14 VN.n5 37.5796
R48 VN.n16 VN.n3 37.5796
R49 VN.n45 VN.n36 37.5796
R50 VN.n47 VN.n34 37.5796
R51 VN.n23 VN.n1 31.752
R52 VN.n54 VN.n32 31.752
R53 VN.n10 VN.n9 24.4675
R54 VN.n15 VN.n14 24.4675
R55 VN.n16 VN.n15 24.4675
R56 VN.n21 VN.n20 24.4675
R57 VN.n28 VN.n27 24.4675
R58 VN.n41 VN.n40 24.4675
R59 VN.n47 VN.n46 24.4675
R60 VN.n46 VN.n45 24.4675
R61 VN.n52 VN.n51 24.4675
R62 VN.n59 VN.n58 24.4675
R63 VN.n23 VN.n22 21.5315
R64 VN.n54 VN.n53 21.5315
R65 VN.n38 VN.n37 18.3181
R66 VN.n7 VN.n6 18.3181
R67 VN.n29 VN.n28 5.87258
R68 VN.n60 VN.n59 5.87258
R69 VN.n9 VN.n8 2.93654
R70 VN.n22 VN.n21 2.93654
R71 VN.n40 VN.n39 2.93654
R72 VN.n53 VN.n52 2.93654
R73 VN.n61 VN.n31 0.189894
R74 VN.n57 VN.n31 0.189894
R75 VN.n57 VN.n56 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n33 0.189894
R78 VN.n50 VN.n33 0.189894
R79 VN.n50 VN.n49 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n35 0.189894
R82 VN.n44 VN.n35 0.189894
R83 VN.n44 VN.n43 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n37 0.189894
R86 VN.n11 VN.n6 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n13 VN.n12 0.189894
R89 VN.n13 VN.n4 0.189894
R90 VN.n17 VN.n4 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n19 VN.n18 0.189894
R93 VN.n19 VN.n2 0.189894
R94 VN.n24 VN.n2 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n26 VN.n25 0.189894
R97 VN.n26 VN.n0 0.189894
R98 VN.n30 VN.n0 0.189894
R99 VN VN.n30 0.0516364
R100 VTAIL.n152 VTAIL.n122 756.745
R101 VTAIL.n32 VTAIL.n2 756.745
R102 VTAIL.n116 VTAIL.n86 756.745
R103 VTAIL.n76 VTAIL.n46 756.745
R104 VTAIL.n135 VTAIL.n134 585
R105 VTAIL.n137 VTAIL.n136 585
R106 VTAIL.n130 VTAIL.n129 585
R107 VTAIL.n143 VTAIL.n142 585
R108 VTAIL.n145 VTAIL.n144 585
R109 VTAIL.n126 VTAIL.n125 585
R110 VTAIL.n151 VTAIL.n150 585
R111 VTAIL.n153 VTAIL.n152 585
R112 VTAIL.n15 VTAIL.n14 585
R113 VTAIL.n17 VTAIL.n16 585
R114 VTAIL.n10 VTAIL.n9 585
R115 VTAIL.n23 VTAIL.n22 585
R116 VTAIL.n25 VTAIL.n24 585
R117 VTAIL.n6 VTAIL.n5 585
R118 VTAIL.n31 VTAIL.n30 585
R119 VTAIL.n33 VTAIL.n32 585
R120 VTAIL.n117 VTAIL.n116 585
R121 VTAIL.n115 VTAIL.n114 585
R122 VTAIL.n90 VTAIL.n89 585
R123 VTAIL.n109 VTAIL.n108 585
R124 VTAIL.n107 VTAIL.n106 585
R125 VTAIL.n94 VTAIL.n93 585
R126 VTAIL.n101 VTAIL.n100 585
R127 VTAIL.n99 VTAIL.n98 585
R128 VTAIL.n77 VTAIL.n76 585
R129 VTAIL.n75 VTAIL.n74 585
R130 VTAIL.n50 VTAIL.n49 585
R131 VTAIL.n69 VTAIL.n68 585
R132 VTAIL.n67 VTAIL.n66 585
R133 VTAIL.n54 VTAIL.n53 585
R134 VTAIL.n61 VTAIL.n60 585
R135 VTAIL.n59 VTAIL.n58 585
R136 VTAIL.n133 VTAIL.t13 327.514
R137 VTAIL.n13 VTAIL.t6 327.514
R138 VTAIL.n97 VTAIL.t9 327.514
R139 VTAIL.n57 VTAIL.t11 327.514
R140 VTAIL.n136 VTAIL.n135 171.744
R141 VTAIL.n136 VTAIL.n129 171.744
R142 VTAIL.n143 VTAIL.n129 171.744
R143 VTAIL.n144 VTAIL.n143 171.744
R144 VTAIL.n144 VTAIL.n125 171.744
R145 VTAIL.n151 VTAIL.n125 171.744
R146 VTAIL.n152 VTAIL.n151 171.744
R147 VTAIL.n16 VTAIL.n15 171.744
R148 VTAIL.n16 VTAIL.n9 171.744
R149 VTAIL.n23 VTAIL.n9 171.744
R150 VTAIL.n24 VTAIL.n23 171.744
R151 VTAIL.n24 VTAIL.n5 171.744
R152 VTAIL.n31 VTAIL.n5 171.744
R153 VTAIL.n32 VTAIL.n31 171.744
R154 VTAIL.n116 VTAIL.n115 171.744
R155 VTAIL.n115 VTAIL.n89 171.744
R156 VTAIL.n108 VTAIL.n89 171.744
R157 VTAIL.n108 VTAIL.n107 171.744
R158 VTAIL.n107 VTAIL.n93 171.744
R159 VTAIL.n100 VTAIL.n93 171.744
R160 VTAIL.n100 VTAIL.n99 171.744
R161 VTAIL.n76 VTAIL.n75 171.744
R162 VTAIL.n75 VTAIL.n49 171.744
R163 VTAIL.n68 VTAIL.n49 171.744
R164 VTAIL.n68 VTAIL.n67 171.744
R165 VTAIL.n67 VTAIL.n53 171.744
R166 VTAIL.n60 VTAIL.n53 171.744
R167 VTAIL.n60 VTAIL.n59 171.744
R168 VTAIL.n135 VTAIL.t13 85.8723
R169 VTAIL.n15 VTAIL.t6 85.8723
R170 VTAIL.n99 VTAIL.t9 85.8723
R171 VTAIL.n59 VTAIL.t11 85.8723
R172 VTAIL.n85 VTAIL.n84 70.7505
R173 VTAIL.n83 VTAIL.n82 70.7505
R174 VTAIL.n45 VTAIL.n44 70.7505
R175 VTAIL.n43 VTAIL.n42 70.7505
R176 VTAIL.n159 VTAIL.n158 70.7503
R177 VTAIL.n1 VTAIL.n0 70.7503
R178 VTAIL.n39 VTAIL.n38 70.7503
R179 VTAIL.n41 VTAIL.n40 70.7503
R180 VTAIL.n157 VTAIL.n156 31.2157
R181 VTAIL.n37 VTAIL.n36 31.2157
R182 VTAIL.n121 VTAIL.n120 31.2157
R183 VTAIL.n81 VTAIL.n80 31.2157
R184 VTAIL.n43 VTAIL.n41 21.6686
R185 VTAIL.n157 VTAIL.n121 19.8927
R186 VTAIL.n134 VTAIL.n133 16.3884
R187 VTAIL.n14 VTAIL.n13 16.3884
R188 VTAIL.n98 VTAIL.n97 16.3884
R189 VTAIL.n58 VTAIL.n57 16.3884
R190 VTAIL.n137 VTAIL.n132 12.8005
R191 VTAIL.n17 VTAIL.n12 12.8005
R192 VTAIL.n101 VTAIL.n96 12.8005
R193 VTAIL.n61 VTAIL.n56 12.8005
R194 VTAIL.n138 VTAIL.n130 12.0247
R195 VTAIL.n18 VTAIL.n10 12.0247
R196 VTAIL.n102 VTAIL.n94 12.0247
R197 VTAIL.n62 VTAIL.n54 12.0247
R198 VTAIL.n142 VTAIL.n141 11.249
R199 VTAIL.n22 VTAIL.n21 11.249
R200 VTAIL.n106 VTAIL.n105 11.249
R201 VTAIL.n66 VTAIL.n65 11.249
R202 VTAIL.n145 VTAIL.n128 10.4732
R203 VTAIL.n25 VTAIL.n8 10.4732
R204 VTAIL.n109 VTAIL.n92 10.4732
R205 VTAIL.n69 VTAIL.n52 10.4732
R206 VTAIL.n146 VTAIL.n126 9.69747
R207 VTAIL.n26 VTAIL.n6 9.69747
R208 VTAIL.n110 VTAIL.n90 9.69747
R209 VTAIL.n70 VTAIL.n50 9.69747
R210 VTAIL.n156 VTAIL.n155 9.45567
R211 VTAIL.n36 VTAIL.n35 9.45567
R212 VTAIL.n120 VTAIL.n119 9.45567
R213 VTAIL.n80 VTAIL.n79 9.45567
R214 VTAIL.n124 VTAIL.n123 9.3005
R215 VTAIL.n149 VTAIL.n148 9.3005
R216 VTAIL.n147 VTAIL.n146 9.3005
R217 VTAIL.n128 VTAIL.n127 9.3005
R218 VTAIL.n141 VTAIL.n140 9.3005
R219 VTAIL.n139 VTAIL.n138 9.3005
R220 VTAIL.n132 VTAIL.n131 9.3005
R221 VTAIL.n155 VTAIL.n154 9.3005
R222 VTAIL.n4 VTAIL.n3 9.3005
R223 VTAIL.n29 VTAIL.n28 9.3005
R224 VTAIL.n27 VTAIL.n26 9.3005
R225 VTAIL.n8 VTAIL.n7 9.3005
R226 VTAIL.n21 VTAIL.n20 9.3005
R227 VTAIL.n19 VTAIL.n18 9.3005
R228 VTAIL.n12 VTAIL.n11 9.3005
R229 VTAIL.n35 VTAIL.n34 9.3005
R230 VTAIL.n119 VTAIL.n118 9.3005
R231 VTAIL.n88 VTAIL.n87 9.3005
R232 VTAIL.n113 VTAIL.n112 9.3005
R233 VTAIL.n111 VTAIL.n110 9.3005
R234 VTAIL.n92 VTAIL.n91 9.3005
R235 VTAIL.n105 VTAIL.n104 9.3005
R236 VTAIL.n103 VTAIL.n102 9.3005
R237 VTAIL.n96 VTAIL.n95 9.3005
R238 VTAIL.n79 VTAIL.n78 9.3005
R239 VTAIL.n48 VTAIL.n47 9.3005
R240 VTAIL.n73 VTAIL.n72 9.3005
R241 VTAIL.n71 VTAIL.n70 9.3005
R242 VTAIL.n52 VTAIL.n51 9.3005
R243 VTAIL.n65 VTAIL.n64 9.3005
R244 VTAIL.n63 VTAIL.n62 9.3005
R245 VTAIL.n56 VTAIL.n55 9.3005
R246 VTAIL.n150 VTAIL.n149 8.92171
R247 VTAIL.n30 VTAIL.n29 8.92171
R248 VTAIL.n114 VTAIL.n113 8.92171
R249 VTAIL.n74 VTAIL.n73 8.92171
R250 VTAIL.n153 VTAIL.n124 8.14595
R251 VTAIL.n33 VTAIL.n4 8.14595
R252 VTAIL.n117 VTAIL.n88 8.14595
R253 VTAIL.n77 VTAIL.n48 8.14595
R254 VTAIL.n154 VTAIL.n122 7.3702
R255 VTAIL.n34 VTAIL.n2 7.3702
R256 VTAIL.n118 VTAIL.n86 7.3702
R257 VTAIL.n78 VTAIL.n46 7.3702
R258 VTAIL.n156 VTAIL.n122 6.59444
R259 VTAIL.n36 VTAIL.n2 6.59444
R260 VTAIL.n120 VTAIL.n86 6.59444
R261 VTAIL.n80 VTAIL.n46 6.59444
R262 VTAIL.n154 VTAIL.n153 5.81868
R263 VTAIL.n34 VTAIL.n33 5.81868
R264 VTAIL.n118 VTAIL.n117 5.81868
R265 VTAIL.n78 VTAIL.n77 5.81868
R266 VTAIL.n150 VTAIL.n124 5.04292
R267 VTAIL.n30 VTAIL.n4 5.04292
R268 VTAIL.n114 VTAIL.n88 5.04292
R269 VTAIL.n74 VTAIL.n48 5.04292
R270 VTAIL.n158 VTAIL.t12 4.87381
R271 VTAIL.n158 VTAIL.t17 4.87381
R272 VTAIL.n0 VTAIL.t16 4.87381
R273 VTAIL.n0 VTAIL.t10 4.87381
R274 VTAIL.n38 VTAIL.t2 4.87381
R275 VTAIL.n38 VTAIL.t1 4.87381
R276 VTAIL.n40 VTAIL.t0 4.87381
R277 VTAIL.n40 VTAIL.t5 4.87381
R278 VTAIL.n84 VTAIL.t3 4.87381
R279 VTAIL.n84 VTAIL.t7 4.87381
R280 VTAIL.n82 VTAIL.t8 4.87381
R281 VTAIL.n82 VTAIL.t4 4.87381
R282 VTAIL.n44 VTAIL.t19 4.87381
R283 VTAIL.n44 VTAIL.t15 4.87381
R284 VTAIL.n42 VTAIL.t18 4.87381
R285 VTAIL.n42 VTAIL.t14 4.87381
R286 VTAIL.n149 VTAIL.n126 4.26717
R287 VTAIL.n29 VTAIL.n6 4.26717
R288 VTAIL.n113 VTAIL.n90 4.26717
R289 VTAIL.n73 VTAIL.n50 4.26717
R290 VTAIL.n133 VTAIL.n131 3.71088
R291 VTAIL.n13 VTAIL.n11 3.71088
R292 VTAIL.n97 VTAIL.n95 3.71088
R293 VTAIL.n57 VTAIL.n55 3.71088
R294 VTAIL.n146 VTAIL.n145 3.49141
R295 VTAIL.n26 VTAIL.n25 3.49141
R296 VTAIL.n110 VTAIL.n109 3.49141
R297 VTAIL.n70 VTAIL.n69 3.49141
R298 VTAIL.n142 VTAIL.n128 2.71565
R299 VTAIL.n22 VTAIL.n8 2.71565
R300 VTAIL.n106 VTAIL.n92 2.71565
R301 VTAIL.n66 VTAIL.n52 2.71565
R302 VTAIL.n141 VTAIL.n130 1.93989
R303 VTAIL.n21 VTAIL.n10 1.93989
R304 VTAIL.n105 VTAIL.n94 1.93989
R305 VTAIL.n65 VTAIL.n54 1.93989
R306 VTAIL.n45 VTAIL.n43 1.77636
R307 VTAIL.n81 VTAIL.n45 1.77636
R308 VTAIL.n85 VTAIL.n83 1.77636
R309 VTAIL.n121 VTAIL.n85 1.77636
R310 VTAIL.n41 VTAIL.n39 1.77636
R311 VTAIL.n39 VTAIL.n37 1.77636
R312 VTAIL.n159 VTAIL.n157 1.77636
R313 VTAIL VTAIL.n1 1.39059
R314 VTAIL.n83 VTAIL.n81 1.35826
R315 VTAIL.n37 VTAIL.n1 1.35826
R316 VTAIL.n138 VTAIL.n137 1.16414
R317 VTAIL.n18 VTAIL.n17 1.16414
R318 VTAIL.n102 VTAIL.n101 1.16414
R319 VTAIL.n62 VTAIL.n61 1.16414
R320 VTAIL.n134 VTAIL.n132 0.388379
R321 VTAIL.n14 VTAIL.n12 0.388379
R322 VTAIL.n98 VTAIL.n96 0.388379
R323 VTAIL.n58 VTAIL.n56 0.388379
R324 VTAIL VTAIL.n159 0.386276
R325 VTAIL.n139 VTAIL.n131 0.155672
R326 VTAIL.n140 VTAIL.n139 0.155672
R327 VTAIL.n140 VTAIL.n127 0.155672
R328 VTAIL.n147 VTAIL.n127 0.155672
R329 VTAIL.n148 VTAIL.n147 0.155672
R330 VTAIL.n148 VTAIL.n123 0.155672
R331 VTAIL.n155 VTAIL.n123 0.155672
R332 VTAIL.n19 VTAIL.n11 0.155672
R333 VTAIL.n20 VTAIL.n19 0.155672
R334 VTAIL.n20 VTAIL.n7 0.155672
R335 VTAIL.n27 VTAIL.n7 0.155672
R336 VTAIL.n28 VTAIL.n27 0.155672
R337 VTAIL.n28 VTAIL.n3 0.155672
R338 VTAIL.n35 VTAIL.n3 0.155672
R339 VTAIL.n119 VTAIL.n87 0.155672
R340 VTAIL.n112 VTAIL.n87 0.155672
R341 VTAIL.n112 VTAIL.n111 0.155672
R342 VTAIL.n111 VTAIL.n91 0.155672
R343 VTAIL.n104 VTAIL.n91 0.155672
R344 VTAIL.n104 VTAIL.n103 0.155672
R345 VTAIL.n103 VTAIL.n95 0.155672
R346 VTAIL.n79 VTAIL.n47 0.155672
R347 VTAIL.n72 VTAIL.n47 0.155672
R348 VTAIL.n72 VTAIL.n71 0.155672
R349 VTAIL.n71 VTAIL.n51 0.155672
R350 VTAIL.n64 VTAIL.n51 0.155672
R351 VTAIL.n64 VTAIL.n63 0.155672
R352 VTAIL.n63 VTAIL.n55 0.155672
R353 VDD2.n69 VDD2.n39 756.745
R354 VDD2.n30 VDD2.n0 756.745
R355 VDD2.n70 VDD2.n69 585
R356 VDD2.n68 VDD2.n67 585
R357 VDD2.n43 VDD2.n42 585
R358 VDD2.n62 VDD2.n61 585
R359 VDD2.n60 VDD2.n59 585
R360 VDD2.n47 VDD2.n46 585
R361 VDD2.n54 VDD2.n53 585
R362 VDD2.n52 VDD2.n51 585
R363 VDD2.n13 VDD2.n12 585
R364 VDD2.n15 VDD2.n14 585
R365 VDD2.n8 VDD2.n7 585
R366 VDD2.n21 VDD2.n20 585
R367 VDD2.n23 VDD2.n22 585
R368 VDD2.n4 VDD2.n3 585
R369 VDD2.n29 VDD2.n28 585
R370 VDD2.n31 VDD2.n30 585
R371 VDD2.n50 VDD2.t9 327.514
R372 VDD2.n11 VDD2.t1 327.514
R373 VDD2.n69 VDD2.n68 171.744
R374 VDD2.n68 VDD2.n42 171.744
R375 VDD2.n61 VDD2.n42 171.744
R376 VDD2.n61 VDD2.n60 171.744
R377 VDD2.n60 VDD2.n46 171.744
R378 VDD2.n53 VDD2.n46 171.744
R379 VDD2.n53 VDD2.n52 171.744
R380 VDD2.n14 VDD2.n13 171.744
R381 VDD2.n14 VDD2.n7 171.744
R382 VDD2.n21 VDD2.n7 171.744
R383 VDD2.n22 VDD2.n21 171.744
R384 VDD2.n22 VDD2.n3 171.744
R385 VDD2.n29 VDD2.n3 171.744
R386 VDD2.n30 VDD2.n29 171.744
R387 VDD2.n38 VDD2.n37 88.7057
R388 VDD2 VDD2.n77 88.7028
R389 VDD2.n76 VDD2.n75 87.4293
R390 VDD2.n36 VDD2.n35 87.4291
R391 VDD2.n52 VDD2.t9 85.8723
R392 VDD2.n13 VDD2.t1 85.8723
R393 VDD2.n36 VDD2.n34 49.6703
R394 VDD2.n74 VDD2.n73 47.8944
R395 VDD2.n74 VDD2.n38 37.9006
R396 VDD2.n12 VDD2.n11 16.3884
R397 VDD2.n51 VDD2.n50 16.3884
R398 VDD2.n54 VDD2.n49 12.8005
R399 VDD2.n15 VDD2.n10 12.8005
R400 VDD2.n55 VDD2.n47 12.0247
R401 VDD2.n16 VDD2.n8 12.0247
R402 VDD2.n59 VDD2.n58 11.249
R403 VDD2.n20 VDD2.n19 11.249
R404 VDD2.n62 VDD2.n45 10.4732
R405 VDD2.n23 VDD2.n6 10.4732
R406 VDD2.n63 VDD2.n43 9.69747
R407 VDD2.n24 VDD2.n4 9.69747
R408 VDD2.n73 VDD2.n72 9.45567
R409 VDD2.n34 VDD2.n33 9.45567
R410 VDD2.n72 VDD2.n71 9.3005
R411 VDD2.n41 VDD2.n40 9.3005
R412 VDD2.n66 VDD2.n65 9.3005
R413 VDD2.n64 VDD2.n63 9.3005
R414 VDD2.n45 VDD2.n44 9.3005
R415 VDD2.n58 VDD2.n57 9.3005
R416 VDD2.n56 VDD2.n55 9.3005
R417 VDD2.n49 VDD2.n48 9.3005
R418 VDD2.n2 VDD2.n1 9.3005
R419 VDD2.n27 VDD2.n26 9.3005
R420 VDD2.n25 VDD2.n24 9.3005
R421 VDD2.n6 VDD2.n5 9.3005
R422 VDD2.n19 VDD2.n18 9.3005
R423 VDD2.n17 VDD2.n16 9.3005
R424 VDD2.n10 VDD2.n9 9.3005
R425 VDD2.n33 VDD2.n32 9.3005
R426 VDD2.n67 VDD2.n66 8.92171
R427 VDD2.n28 VDD2.n27 8.92171
R428 VDD2.n70 VDD2.n41 8.14595
R429 VDD2.n31 VDD2.n2 8.14595
R430 VDD2.n71 VDD2.n39 7.3702
R431 VDD2.n32 VDD2.n0 7.3702
R432 VDD2.n73 VDD2.n39 6.59444
R433 VDD2.n34 VDD2.n0 6.59444
R434 VDD2.n71 VDD2.n70 5.81868
R435 VDD2.n32 VDD2.n31 5.81868
R436 VDD2.n67 VDD2.n41 5.04292
R437 VDD2.n28 VDD2.n2 5.04292
R438 VDD2.n77 VDD2.t5 4.87381
R439 VDD2.n77 VDD2.t4 4.87381
R440 VDD2.n75 VDD2.t6 4.87381
R441 VDD2.n75 VDD2.t7 4.87381
R442 VDD2.n37 VDD2.t8 4.87381
R443 VDD2.n37 VDD2.t0 4.87381
R444 VDD2.n35 VDD2.t2 4.87381
R445 VDD2.n35 VDD2.t3 4.87381
R446 VDD2.n66 VDD2.n43 4.26717
R447 VDD2.n27 VDD2.n4 4.26717
R448 VDD2.n50 VDD2.n48 3.71088
R449 VDD2.n11 VDD2.n9 3.71088
R450 VDD2.n63 VDD2.n62 3.49141
R451 VDD2.n24 VDD2.n23 3.49141
R452 VDD2.n59 VDD2.n45 2.71565
R453 VDD2.n20 VDD2.n6 2.71565
R454 VDD2.n58 VDD2.n47 1.93989
R455 VDD2.n19 VDD2.n8 1.93989
R456 VDD2.n76 VDD2.n74 1.77636
R457 VDD2.n55 VDD2.n54 1.16414
R458 VDD2.n16 VDD2.n15 1.16414
R459 VDD2 VDD2.n76 0.502655
R460 VDD2.n38 VDD2.n36 0.389119
R461 VDD2.n51 VDD2.n49 0.388379
R462 VDD2.n12 VDD2.n10 0.388379
R463 VDD2.n72 VDD2.n40 0.155672
R464 VDD2.n65 VDD2.n40 0.155672
R465 VDD2.n65 VDD2.n64 0.155672
R466 VDD2.n64 VDD2.n44 0.155672
R467 VDD2.n57 VDD2.n44 0.155672
R468 VDD2.n57 VDD2.n56 0.155672
R469 VDD2.n56 VDD2.n48 0.155672
R470 VDD2.n17 VDD2.n9 0.155672
R471 VDD2.n18 VDD2.n17 0.155672
R472 VDD2.n18 VDD2.n5 0.155672
R473 VDD2.n25 VDD2.n5 0.155672
R474 VDD2.n26 VDD2.n25 0.155672
R475 VDD2.n26 VDD2.n1 0.155672
R476 VDD2.n33 VDD2.n1 0.155672
R477 VP.n41 VP.n40 179.895
R478 VP.n70 VP.n69 179.895
R479 VP.n39 VP.n38 179.895
R480 VP.n18 VP.n15 161.3
R481 VP.n20 VP.n19 161.3
R482 VP.n21 VP.n14 161.3
R483 VP.n23 VP.n22 161.3
R484 VP.n24 VP.n13 161.3
R485 VP.n26 VP.n25 161.3
R486 VP.n27 VP.n12 161.3
R487 VP.n29 VP.n28 161.3
R488 VP.n30 VP.n11 161.3
R489 VP.n33 VP.n32 161.3
R490 VP.n34 VP.n10 161.3
R491 VP.n36 VP.n35 161.3
R492 VP.n37 VP.n9 161.3
R493 VP.n68 VP.n0 161.3
R494 VP.n67 VP.n66 161.3
R495 VP.n65 VP.n1 161.3
R496 VP.n64 VP.n63 161.3
R497 VP.n61 VP.n2 161.3
R498 VP.n60 VP.n59 161.3
R499 VP.n58 VP.n3 161.3
R500 VP.n57 VP.n56 161.3
R501 VP.n55 VP.n4 161.3
R502 VP.n54 VP.n53 161.3
R503 VP.n52 VP.n5 161.3
R504 VP.n51 VP.n50 161.3
R505 VP.n49 VP.n6 161.3
R506 VP.n47 VP.n46 161.3
R507 VP.n45 VP.n7 161.3
R508 VP.n44 VP.n43 161.3
R509 VP.n42 VP.n8 161.3
R510 VP.n16 VP.t6 123.969
R511 VP.n55 VP.t0 92.9178
R512 VP.n41 VP.t1 92.9178
R513 VP.n48 VP.t8 92.9178
R514 VP.n62 VP.t2 92.9178
R515 VP.n69 VP.t7 92.9178
R516 VP.n24 VP.t5 92.9178
R517 VP.n38 VP.t9 92.9178
R518 VP.n31 VP.t3 92.9178
R519 VP.n17 VP.t4 92.9178
R520 VP.n17 VP.n16 64.8059
R521 VP.n43 VP.n7 49.2348
R522 VP.n67 VP.n1 49.2348
R523 VP.n36 VP.n10 49.2348
R524 VP.n40 VP.n39 44.2656
R525 VP.n50 VP.n5 43.4072
R526 VP.n60 VP.n3 43.4072
R527 VP.n29 VP.n12 43.4072
R528 VP.n19 VP.n14 43.4072
R529 VP.n54 VP.n5 37.5796
R530 VP.n56 VP.n3 37.5796
R531 VP.n25 VP.n12 37.5796
R532 VP.n23 VP.n14 37.5796
R533 VP.n47 VP.n7 31.752
R534 VP.n63 VP.n1 31.752
R535 VP.n32 VP.n10 31.752
R536 VP.n43 VP.n42 24.4675
R537 VP.n50 VP.n49 24.4675
R538 VP.n55 VP.n54 24.4675
R539 VP.n56 VP.n55 24.4675
R540 VP.n61 VP.n60 24.4675
R541 VP.n68 VP.n67 24.4675
R542 VP.n37 VP.n36 24.4675
R543 VP.n30 VP.n29 24.4675
R544 VP.n24 VP.n23 24.4675
R545 VP.n25 VP.n24 24.4675
R546 VP.n19 VP.n18 24.4675
R547 VP.n48 VP.n47 21.5315
R548 VP.n63 VP.n62 21.5315
R549 VP.n32 VP.n31 21.5315
R550 VP.n16 VP.n15 18.3181
R551 VP.n42 VP.n41 5.87258
R552 VP.n69 VP.n68 5.87258
R553 VP.n38 VP.n37 5.87258
R554 VP.n49 VP.n48 2.93654
R555 VP.n62 VP.n61 2.93654
R556 VP.n31 VP.n30 2.93654
R557 VP.n18 VP.n17 2.93654
R558 VP.n20 VP.n15 0.189894
R559 VP.n21 VP.n20 0.189894
R560 VP.n22 VP.n21 0.189894
R561 VP.n22 VP.n13 0.189894
R562 VP.n26 VP.n13 0.189894
R563 VP.n27 VP.n26 0.189894
R564 VP.n28 VP.n27 0.189894
R565 VP.n28 VP.n11 0.189894
R566 VP.n33 VP.n11 0.189894
R567 VP.n34 VP.n33 0.189894
R568 VP.n35 VP.n34 0.189894
R569 VP.n35 VP.n9 0.189894
R570 VP.n39 VP.n9 0.189894
R571 VP.n40 VP.n8 0.189894
R572 VP.n44 VP.n8 0.189894
R573 VP.n45 VP.n44 0.189894
R574 VP.n46 VP.n45 0.189894
R575 VP.n46 VP.n6 0.189894
R576 VP.n51 VP.n6 0.189894
R577 VP.n52 VP.n51 0.189894
R578 VP.n53 VP.n52 0.189894
R579 VP.n53 VP.n4 0.189894
R580 VP.n57 VP.n4 0.189894
R581 VP.n58 VP.n57 0.189894
R582 VP.n59 VP.n58 0.189894
R583 VP.n59 VP.n2 0.189894
R584 VP.n64 VP.n2 0.189894
R585 VP.n65 VP.n64 0.189894
R586 VP.n66 VP.n65 0.189894
R587 VP.n66 VP.n0 0.189894
R588 VP.n70 VP.n0 0.189894
R589 VP VP.n70 0.0516364
R590 VDD1.n30 VDD1.n0 756.745
R591 VDD1.n67 VDD1.n37 756.745
R592 VDD1.n31 VDD1.n30 585
R593 VDD1.n29 VDD1.n28 585
R594 VDD1.n4 VDD1.n3 585
R595 VDD1.n23 VDD1.n22 585
R596 VDD1.n21 VDD1.n20 585
R597 VDD1.n8 VDD1.n7 585
R598 VDD1.n15 VDD1.n14 585
R599 VDD1.n13 VDD1.n12 585
R600 VDD1.n50 VDD1.n49 585
R601 VDD1.n52 VDD1.n51 585
R602 VDD1.n45 VDD1.n44 585
R603 VDD1.n58 VDD1.n57 585
R604 VDD1.n60 VDD1.n59 585
R605 VDD1.n41 VDD1.n40 585
R606 VDD1.n66 VDD1.n65 585
R607 VDD1.n68 VDD1.n67 585
R608 VDD1.n11 VDD1.t3 327.514
R609 VDD1.n48 VDD1.t8 327.514
R610 VDD1.n30 VDD1.n29 171.744
R611 VDD1.n29 VDD1.n3 171.744
R612 VDD1.n22 VDD1.n3 171.744
R613 VDD1.n22 VDD1.n21 171.744
R614 VDD1.n21 VDD1.n7 171.744
R615 VDD1.n14 VDD1.n7 171.744
R616 VDD1.n14 VDD1.n13 171.744
R617 VDD1.n51 VDD1.n50 171.744
R618 VDD1.n51 VDD1.n44 171.744
R619 VDD1.n58 VDD1.n44 171.744
R620 VDD1.n59 VDD1.n58 171.744
R621 VDD1.n59 VDD1.n40 171.744
R622 VDD1.n66 VDD1.n40 171.744
R623 VDD1.n67 VDD1.n66 171.744
R624 VDD1.n75 VDD1.n74 88.7057
R625 VDD1.n36 VDD1.n35 87.4293
R626 VDD1.n77 VDD1.n76 87.4291
R627 VDD1.n73 VDD1.n72 87.4291
R628 VDD1.n13 VDD1.t3 85.8723
R629 VDD1.n50 VDD1.t8 85.8723
R630 VDD1.n36 VDD1.n34 49.6703
R631 VDD1.n73 VDD1.n71 49.6703
R632 VDD1.n77 VDD1.n75 39.3716
R633 VDD1.n49 VDD1.n48 16.3884
R634 VDD1.n12 VDD1.n11 16.3884
R635 VDD1.n15 VDD1.n10 12.8005
R636 VDD1.n52 VDD1.n47 12.8005
R637 VDD1.n16 VDD1.n8 12.0247
R638 VDD1.n53 VDD1.n45 12.0247
R639 VDD1.n20 VDD1.n19 11.249
R640 VDD1.n57 VDD1.n56 11.249
R641 VDD1.n23 VDD1.n6 10.4732
R642 VDD1.n60 VDD1.n43 10.4732
R643 VDD1.n24 VDD1.n4 9.69747
R644 VDD1.n61 VDD1.n41 9.69747
R645 VDD1.n34 VDD1.n33 9.45567
R646 VDD1.n71 VDD1.n70 9.45567
R647 VDD1.n33 VDD1.n32 9.3005
R648 VDD1.n2 VDD1.n1 9.3005
R649 VDD1.n27 VDD1.n26 9.3005
R650 VDD1.n25 VDD1.n24 9.3005
R651 VDD1.n6 VDD1.n5 9.3005
R652 VDD1.n19 VDD1.n18 9.3005
R653 VDD1.n17 VDD1.n16 9.3005
R654 VDD1.n10 VDD1.n9 9.3005
R655 VDD1.n39 VDD1.n38 9.3005
R656 VDD1.n64 VDD1.n63 9.3005
R657 VDD1.n62 VDD1.n61 9.3005
R658 VDD1.n43 VDD1.n42 9.3005
R659 VDD1.n56 VDD1.n55 9.3005
R660 VDD1.n54 VDD1.n53 9.3005
R661 VDD1.n47 VDD1.n46 9.3005
R662 VDD1.n70 VDD1.n69 9.3005
R663 VDD1.n28 VDD1.n27 8.92171
R664 VDD1.n65 VDD1.n64 8.92171
R665 VDD1.n31 VDD1.n2 8.14595
R666 VDD1.n68 VDD1.n39 8.14595
R667 VDD1.n32 VDD1.n0 7.3702
R668 VDD1.n69 VDD1.n37 7.3702
R669 VDD1.n34 VDD1.n0 6.59444
R670 VDD1.n71 VDD1.n37 6.59444
R671 VDD1.n32 VDD1.n31 5.81868
R672 VDD1.n69 VDD1.n68 5.81868
R673 VDD1.n28 VDD1.n2 5.04292
R674 VDD1.n65 VDD1.n39 5.04292
R675 VDD1.n76 VDD1.t6 4.87381
R676 VDD1.n76 VDD1.t0 4.87381
R677 VDD1.n35 VDD1.t5 4.87381
R678 VDD1.n35 VDD1.t4 4.87381
R679 VDD1.n74 VDD1.t7 4.87381
R680 VDD1.n74 VDD1.t2 4.87381
R681 VDD1.n72 VDD1.t1 4.87381
R682 VDD1.n72 VDD1.t9 4.87381
R683 VDD1.n27 VDD1.n4 4.26717
R684 VDD1.n64 VDD1.n41 4.26717
R685 VDD1.n11 VDD1.n9 3.71088
R686 VDD1.n48 VDD1.n46 3.71088
R687 VDD1.n24 VDD1.n23 3.49141
R688 VDD1.n61 VDD1.n60 3.49141
R689 VDD1.n20 VDD1.n6 2.71565
R690 VDD1.n57 VDD1.n43 2.71565
R691 VDD1.n19 VDD1.n8 1.93989
R692 VDD1.n56 VDD1.n45 1.93989
R693 VDD1 VDD1.n77 1.27421
R694 VDD1.n16 VDD1.n15 1.16414
R695 VDD1.n53 VDD1.n52 1.16414
R696 VDD1 VDD1.n36 0.502655
R697 VDD1.n75 VDD1.n73 0.389119
R698 VDD1.n12 VDD1.n10 0.388379
R699 VDD1.n49 VDD1.n47 0.388379
R700 VDD1.n33 VDD1.n1 0.155672
R701 VDD1.n26 VDD1.n1 0.155672
R702 VDD1.n26 VDD1.n25 0.155672
R703 VDD1.n25 VDD1.n5 0.155672
R704 VDD1.n18 VDD1.n5 0.155672
R705 VDD1.n18 VDD1.n17 0.155672
R706 VDD1.n17 VDD1.n9 0.155672
R707 VDD1.n54 VDD1.n46 0.155672
R708 VDD1.n55 VDD1.n54 0.155672
R709 VDD1.n55 VDD1.n42 0.155672
R710 VDD1.n62 VDD1.n42 0.155672
R711 VDD1.n63 VDD1.n62 0.155672
R712 VDD1.n63 VDD1.n38 0.155672
R713 VDD1.n70 VDD1.n38 0.155672
R714 B.n317 B.n316 585
R715 B.n315 B.n104 585
R716 B.n314 B.n313 585
R717 B.n312 B.n105 585
R718 B.n311 B.n310 585
R719 B.n309 B.n106 585
R720 B.n308 B.n307 585
R721 B.n306 B.n107 585
R722 B.n305 B.n304 585
R723 B.n303 B.n108 585
R724 B.n302 B.n301 585
R725 B.n300 B.n109 585
R726 B.n299 B.n298 585
R727 B.n297 B.n110 585
R728 B.n296 B.n295 585
R729 B.n294 B.n111 585
R730 B.n293 B.n292 585
R731 B.n291 B.n112 585
R732 B.n290 B.n289 585
R733 B.n288 B.n113 585
R734 B.n287 B.n286 585
R735 B.n285 B.n114 585
R736 B.n284 B.n283 585
R737 B.n282 B.n115 585
R738 B.n281 B.n280 585
R739 B.n279 B.n116 585
R740 B.n278 B.n277 585
R741 B.n273 B.n117 585
R742 B.n272 B.n271 585
R743 B.n270 B.n118 585
R744 B.n269 B.n268 585
R745 B.n267 B.n119 585
R746 B.n266 B.n265 585
R747 B.n264 B.n120 585
R748 B.n263 B.n262 585
R749 B.n260 B.n121 585
R750 B.n259 B.n258 585
R751 B.n257 B.n124 585
R752 B.n256 B.n255 585
R753 B.n254 B.n125 585
R754 B.n253 B.n252 585
R755 B.n251 B.n126 585
R756 B.n250 B.n249 585
R757 B.n248 B.n127 585
R758 B.n247 B.n246 585
R759 B.n245 B.n128 585
R760 B.n244 B.n243 585
R761 B.n242 B.n129 585
R762 B.n241 B.n240 585
R763 B.n239 B.n130 585
R764 B.n238 B.n237 585
R765 B.n236 B.n131 585
R766 B.n235 B.n234 585
R767 B.n233 B.n132 585
R768 B.n232 B.n231 585
R769 B.n230 B.n133 585
R770 B.n229 B.n228 585
R771 B.n227 B.n134 585
R772 B.n226 B.n225 585
R773 B.n224 B.n135 585
R774 B.n223 B.n222 585
R775 B.n318 B.n103 585
R776 B.n320 B.n319 585
R777 B.n321 B.n102 585
R778 B.n323 B.n322 585
R779 B.n324 B.n101 585
R780 B.n326 B.n325 585
R781 B.n327 B.n100 585
R782 B.n329 B.n328 585
R783 B.n330 B.n99 585
R784 B.n332 B.n331 585
R785 B.n333 B.n98 585
R786 B.n335 B.n334 585
R787 B.n336 B.n97 585
R788 B.n338 B.n337 585
R789 B.n339 B.n96 585
R790 B.n341 B.n340 585
R791 B.n342 B.n95 585
R792 B.n344 B.n343 585
R793 B.n345 B.n94 585
R794 B.n347 B.n346 585
R795 B.n348 B.n93 585
R796 B.n350 B.n349 585
R797 B.n351 B.n92 585
R798 B.n353 B.n352 585
R799 B.n354 B.n91 585
R800 B.n356 B.n355 585
R801 B.n357 B.n90 585
R802 B.n359 B.n358 585
R803 B.n360 B.n89 585
R804 B.n362 B.n361 585
R805 B.n363 B.n88 585
R806 B.n365 B.n364 585
R807 B.n366 B.n87 585
R808 B.n368 B.n367 585
R809 B.n369 B.n86 585
R810 B.n371 B.n370 585
R811 B.n372 B.n85 585
R812 B.n374 B.n373 585
R813 B.n375 B.n84 585
R814 B.n377 B.n376 585
R815 B.n378 B.n83 585
R816 B.n380 B.n379 585
R817 B.n381 B.n82 585
R818 B.n383 B.n382 585
R819 B.n384 B.n81 585
R820 B.n386 B.n385 585
R821 B.n387 B.n80 585
R822 B.n389 B.n388 585
R823 B.n390 B.n79 585
R824 B.n392 B.n391 585
R825 B.n393 B.n78 585
R826 B.n395 B.n394 585
R827 B.n396 B.n77 585
R828 B.n398 B.n397 585
R829 B.n399 B.n76 585
R830 B.n401 B.n400 585
R831 B.n402 B.n75 585
R832 B.n404 B.n403 585
R833 B.n405 B.n74 585
R834 B.n407 B.n406 585
R835 B.n408 B.n73 585
R836 B.n410 B.n409 585
R837 B.n411 B.n72 585
R838 B.n413 B.n412 585
R839 B.n414 B.n71 585
R840 B.n416 B.n415 585
R841 B.n417 B.n70 585
R842 B.n419 B.n418 585
R843 B.n420 B.n69 585
R844 B.n422 B.n421 585
R845 B.n423 B.n68 585
R846 B.n425 B.n424 585
R847 B.n426 B.n67 585
R848 B.n428 B.n427 585
R849 B.n429 B.n66 585
R850 B.n431 B.n430 585
R851 B.n432 B.n65 585
R852 B.n434 B.n433 585
R853 B.n435 B.n64 585
R854 B.n437 B.n436 585
R855 B.n438 B.n63 585
R856 B.n440 B.n439 585
R857 B.n441 B.n62 585
R858 B.n443 B.n442 585
R859 B.n444 B.n61 585
R860 B.n446 B.n445 585
R861 B.n447 B.n60 585
R862 B.n449 B.n448 585
R863 B.n450 B.n59 585
R864 B.n452 B.n451 585
R865 B.n545 B.n24 585
R866 B.n544 B.n543 585
R867 B.n542 B.n25 585
R868 B.n541 B.n540 585
R869 B.n539 B.n26 585
R870 B.n538 B.n537 585
R871 B.n536 B.n27 585
R872 B.n535 B.n534 585
R873 B.n533 B.n28 585
R874 B.n532 B.n531 585
R875 B.n530 B.n29 585
R876 B.n529 B.n528 585
R877 B.n527 B.n30 585
R878 B.n526 B.n525 585
R879 B.n524 B.n31 585
R880 B.n523 B.n522 585
R881 B.n521 B.n32 585
R882 B.n520 B.n519 585
R883 B.n518 B.n33 585
R884 B.n517 B.n516 585
R885 B.n515 B.n34 585
R886 B.n514 B.n513 585
R887 B.n512 B.n35 585
R888 B.n511 B.n510 585
R889 B.n509 B.n36 585
R890 B.n508 B.n507 585
R891 B.n505 B.n37 585
R892 B.n504 B.n503 585
R893 B.n502 B.n40 585
R894 B.n501 B.n500 585
R895 B.n499 B.n41 585
R896 B.n498 B.n497 585
R897 B.n496 B.n42 585
R898 B.n495 B.n494 585
R899 B.n493 B.n43 585
R900 B.n491 B.n490 585
R901 B.n489 B.n46 585
R902 B.n488 B.n487 585
R903 B.n486 B.n47 585
R904 B.n485 B.n484 585
R905 B.n483 B.n48 585
R906 B.n482 B.n481 585
R907 B.n480 B.n49 585
R908 B.n479 B.n478 585
R909 B.n477 B.n50 585
R910 B.n476 B.n475 585
R911 B.n474 B.n51 585
R912 B.n473 B.n472 585
R913 B.n471 B.n52 585
R914 B.n470 B.n469 585
R915 B.n468 B.n53 585
R916 B.n467 B.n466 585
R917 B.n465 B.n54 585
R918 B.n464 B.n463 585
R919 B.n462 B.n55 585
R920 B.n461 B.n460 585
R921 B.n459 B.n56 585
R922 B.n458 B.n457 585
R923 B.n456 B.n57 585
R924 B.n455 B.n454 585
R925 B.n453 B.n58 585
R926 B.n547 B.n546 585
R927 B.n548 B.n23 585
R928 B.n550 B.n549 585
R929 B.n551 B.n22 585
R930 B.n553 B.n552 585
R931 B.n554 B.n21 585
R932 B.n556 B.n555 585
R933 B.n557 B.n20 585
R934 B.n559 B.n558 585
R935 B.n560 B.n19 585
R936 B.n562 B.n561 585
R937 B.n563 B.n18 585
R938 B.n565 B.n564 585
R939 B.n566 B.n17 585
R940 B.n568 B.n567 585
R941 B.n569 B.n16 585
R942 B.n571 B.n570 585
R943 B.n572 B.n15 585
R944 B.n574 B.n573 585
R945 B.n575 B.n14 585
R946 B.n577 B.n576 585
R947 B.n578 B.n13 585
R948 B.n580 B.n579 585
R949 B.n581 B.n12 585
R950 B.n583 B.n582 585
R951 B.n584 B.n11 585
R952 B.n586 B.n585 585
R953 B.n587 B.n10 585
R954 B.n589 B.n588 585
R955 B.n590 B.n9 585
R956 B.n592 B.n591 585
R957 B.n593 B.n8 585
R958 B.n595 B.n594 585
R959 B.n596 B.n7 585
R960 B.n598 B.n597 585
R961 B.n599 B.n6 585
R962 B.n601 B.n600 585
R963 B.n602 B.n5 585
R964 B.n604 B.n603 585
R965 B.n605 B.n4 585
R966 B.n607 B.n606 585
R967 B.n608 B.n3 585
R968 B.n610 B.n609 585
R969 B.n611 B.n0 585
R970 B.n2 B.n1 585
R971 B.n158 B.n157 585
R972 B.n160 B.n159 585
R973 B.n161 B.n156 585
R974 B.n163 B.n162 585
R975 B.n164 B.n155 585
R976 B.n166 B.n165 585
R977 B.n167 B.n154 585
R978 B.n169 B.n168 585
R979 B.n170 B.n153 585
R980 B.n172 B.n171 585
R981 B.n173 B.n152 585
R982 B.n175 B.n174 585
R983 B.n176 B.n151 585
R984 B.n178 B.n177 585
R985 B.n179 B.n150 585
R986 B.n181 B.n180 585
R987 B.n182 B.n149 585
R988 B.n184 B.n183 585
R989 B.n185 B.n148 585
R990 B.n187 B.n186 585
R991 B.n188 B.n147 585
R992 B.n190 B.n189 585
R993 B.n191 B.n146 585
R994 B.n193 B.n192 585
R995 B.n194 B.n145 585
R996 B.n196 B.n195 585
R997 B.n197 B.n144 585
R998 B.n199 B.n198 585
R999 B.n200 B.n143 585
R1000 B.n202 B.n201 585
R1001 B.n203 B.n142 585
R1002 B.n205 B.n204 585
R1003 B.n206 B.n141 585
R1004 B.n208 B.n207 585
R1005 B.n209 B.n140 585
R1006 B.n211 B.n210 585
R1007 B.n212 B.n139 585
R1008 B.n214 B.n213 585
R1009 B.n215 B.n138 585
R1010 B.n217 B.n216 585
R1011 B.n218 B.n137 585
R1012 B.n220 B.n219 585
R1013 B.n221 B.n136 585
R1014 B.n222 B.n221 530.939
R1015 B.n316 B.n103 530.939
R1016 B.n453 B.n452 530.939
R1017 B.n546 B.n545 530.939
R1018 B.n274 B.t1 319.945
R1019 B.n44 B.t11 319.945
R1020 B.n122 B.t7 319.945
R1021 B.n38 B.t5 319.945
R1022 B.n122 B.t6 299.123
R1023 B.n274 B.t0 299.123
R1024 B.n44 B.t9 299.123
R1025 B.n38 B.t3 299.123
R1026 B.n275 B.t2 279.993
R1027 B.n45 B.t10 279.993
R1028 B.n123 B.t8 279.993
R1029 B.n39 B.t4 279.993
R1030 B.n613 B.n612 256.663
R1031 B.n612 B.n611 235.042
R1032 B.n612 B.n2 235.042
R1033 B.n222 B.n135 163.367
R1034 B.n226 B.n135 163.367
R1035 B.n227 B.n226 163.367
R1036 B.n228 B.n227 163.367
R1037 B.n228 B.n133 163.367
R1038 B.n232 B.n133 163.367
R1039 B.n233 B.n232 163.367
R1040 B.n234 B.n233 163.367
R1041 B.n234 B.n131 163.367
R1042 B.n238 B.n131 163.367
R1043 B.n239 B.n238 163.367
R1044 B.n240 B.n239 163.367
R1045 B.n240 B.n129 163.367
R1046 B.n244 B.n129 163.367
R1047 B.n245 B.n244 163.367
R1048 B.n246 B.n245 163.367
R1049 B.n246 B.n127 163.367
R1050 B.n250 B.n127 163.367
R1051 B.n251 B.n250 163.367
R1052 B.n252 B.n251 163.367
R1053 B.n252 B.n125 163.367
R1054 B.n256 B.n125 163.367
R1055 B.n257 B.n256 163.367
R1056 B.n258 B.n257 163.367
R1057 B.n258 B.n121 163.367
R1058 B.n263 B.n121 163.367
R1059 B.n264 B.n263 163.367
R1060 B.n265 B.n264 163.367
R1061 B.n265 B.n119 163.367
R1062 B.n269 B.n119 163.367
R1063 B.n270 B.n269 163.367
R1064 B.n271 B.n270 163.367
R1065 B.n271 B.n117 163.367
R1066 B.n278 B.n117 163.367
R1067 B.n279 B.n278 163.367
R1068 B.n280 B.n279 163.367
R1069 B.n280 B.n115 163.367
R1070 B.n284 B.n115 163.367
R1071 B.n285 B.n284 163.367
R1072 B.n286 B.n285 163.367
R1073 B.n286 B.n113 163.367
R1074 B.n290 B.n113 163.367
R1075 B.n291 B.n290 163.367
R1076 B.n292 B.n291 163.367
R1077 B.n292 B.n111 163.367
R1078 B.n296 B.n111 163.367
R1079 B.n297 B.n296 163.367
R1080 B.n298 B.n297 163.367
R1081 B.n298 B.n109 163.367
R1082 B.n302 B.n109 163.367
R1083 B.n303 B.n302 163.367
R1084 B.n304 B.n303 163.367
R1085 B.n304 B.n107 163.367
R1086 B.n308 B.n107 163.367
R1087 B.n309 B.n308 163.367
R1088 B.n310 B.n309 163.367
R1089 B.n310 B.n105 163.367
R1090 B.n314 B.n105 163.367
R1091 B.n315 B.n314 163.367
R1092 B.n316 B.n315 163.367
R1093 B.n452 B.n59 163.367
R1094 B.n448 B.n59 163.367
R1095 B.n448 B.n447 163.367
R1096 B.n447 B.n446 163.367
R1097 B.n446 B.n61 163.367
R1098 B.n442 B.n61 163.367
R1099 B.n442 B.n441 163.367
R1100 B.n441 B.n440 163.367
R1101 B.n440 B.n63 163.367
R1102 B.n436 B.n63 163.367
R1103 B.n436 B.n435 163.367
R1104 B.n435 B.n434 163.367
R1105 B.n434 B.n65 163.367
R1106 B.n430 B.n65 163.367
R1107 B.n430 B.n429 163.367
R1108 B.n429 B.n428 163.367
R1109 B.n428 B.n67 163.367
R1110 B.n424 B.n67 163.367
R1111 B.n424 B.n423 163.367
R1112 B.n423 B.n422 163.367
R1113 B.n422 B.n69 163.367
R1114 B.n418 B.n69 163.367
R1115 B.n418 B.n417 163.367
R1116 B.n417 B.n416 163.367
R1117 B.n416 B.n71 163.367
R1118 B.n412 B.n71 163.367
R1119 B.n412 B.n411 163.367
R1120 B.n411 B.n410 163.367
R1121 B.n410 B.n73 163.367
R1122 B.n406 B.n73 163.367
R1123 B.n406 B.n405 163.367
R1124 B.n405 B.n404 163.367
R1125 B.n404 B.n75 163.367
R1126 B.n400 B.n75 163.367
R1127 B.n400 B.n399 163.367
R1128 B.n399 B.n398 163.367
R1129 B.n398 B.n77 163.367
R1130 B.n394 B.n77 163.367
R1131 B.n394 B.n393 163.367
R1132 B.n393 B.n392 163.367
R1133 B.n392 B.n79 163.367
R1134 B.n388 B.n79 163.367
R1135 B.n388 B.n387 163.367
R1136 B.n387 B.n386 163.367
R1137 B.n386 B.n81 163.367
R1138 B.n382 B.n81 163.367
R1139 B.n382 B.n381 163.367
R1140 B.n381 B.n380 163.367
R1141 B.n380 B.n83 163.367
R1142 B.n376 B.n83 163.367
R1143 B.n376 B.n375 163.367
R1144 B.n375 B.n374 163.367
R1145 B.n374 B.n85 163.367
R1146 B.n370 B.n85 163.367
R1147 B.n370 B.n369 163.367
R1148 B.n369 B.n368 163.367
R1149 B.n368 B.n87 163.367
R1150 B.n364 B.n87 163.367
R1151 B.n364 B.n363 163.367
R1152 B.n363 B.n362 163.367
R1153 B.n362 B.n89 163.367
R1154 B.n358 B.n89 163.367
R1155 B.n358 B.n357 163.367
R1156 B.n357 B.n356 163.367
R1157 B.n356 B.n91 163.367
R1158 B.n352 B.n91 163.367
R1159 B.n352 B.n351 163.367
R1160 B.n351 B.n350 163.367
R1161 B.n350 B.n93 163.367
R1162 B.n346 B.n93 163.367
R1163 B.n346 B.n345 163.367
R1164 B.n345 B.n344 163.367
R1165 B.n344 B.n95 163.367
R1166 B.n340 B.n95 163.367
R1167 B.n340 B.n339 163.367
R1168 B.n339 B.n338 163.367
R1169 B.n338 B.n97 163.367
R1170 B.n334 B.n97 163.367
R1171 B.n334 B.n333 163.367
R1172 B.n333 B.n332 163.367
R1173 B.n332 B.n99 163.367
R1174 B.n328 B.n99 163.367
R1175 B.n328 B.n327 163.367
R1176 B.n327 B.n326 163.367
R1177 B.n326 B.n101 163.367
R1178 B.n322 B.n101 163.367
R1179 B.n322 B.n321 163.367
R1180 B.n321 B.n320 163.367
R1181 B.n320 B.n103 163.367
R1182 B.n545 B.n544 163.367
R1183 B.n544 B.n25 163.367
R1184 B.n540 B.n25 163.367
R1185 B.n540 B.n539 163.367
R1186 B.n539 B.n538 163.367
R1187 B.n538 B.n27 163.367
R1188 B.n534 B.n27 163.367
R1189 B.n534 B.n533 163.367
R1190 B.n533 B.n532 163.367
R1191 B.n532 B.n29 163.367
R1192 B.n528 B.n29 163.367
R1193 B.n528 B.n527 163.367
R1194 B.n527 B.n526 163.367
R1195 B.n526 B.n31 163.367
R1196 B.n522 B.n31 163.367
R1197 B.n522 B.n521 163.367
R1198 B.n521 B.n520 163.367
R1199 B.n520 B.n33 163.367
R1200 B.n516 B.n33 163.367
R1201 B.n516 B.n515 163.367
R1202 B.n515 B.n514 163.367
R1203 B.n514 B.n35 163.367
R1204 B.n510 B.n35 163.367
R1205 B.n510 B.n509 163.367
R1206 B.n509 B.n508 163.367
R1207 B.n508 B.n37 163.367
R1208 B.n503 B.n37 163.367
R1209 B.n503 B.n502 163.367
R1210 B.n502 B.n501 163.367
R1211 B.n501 B.n41 163.367
R1212 B.n497 B.n41 163.367
R1213 B.n497 B.n496 163.367
R1214 B.n496 B.n495 163.367
R1215 B.n495 B.n43 163.367
R1216 B.n490 B.n43 163.367
R1217 B.n490 B.n489 163.367
R1218 B.n489 B.n488 163.367
R1219 B.n488 B.n47 163.367
R1220 B.n484 B.n47 163.367
R1221 B.n484 B.n483 163.367
R1222 B.n483 B.n482 163.367
R1223 B.n482 B.n49 163.367
R1224 B.n478 B.n49 163.367
R1225 B.n478 B.n477 163.367
R1226 B.n477 B.n476 163.367
R1227 B.n476 B.n51 163.367
R1228 B.n472 B.n51 163.367
R1229 B.n472 B.n471 163.367
R1230 B.n471 B.n470 163.367
R1231 B.n470 B.n53 163.367
R1232 B.n466 B.n53 163.367
R1233 B.n466 B.n465 163.367
R1234 B.n465 B.n464 163.367
R1235 B.n464 B.n55 163.367
R1236 B.n460 B.n55 163.367
R1237 B.n460 B.n459 163.367
R1238 B.n459 B.n458 163.367
R1239 B.n458 B.n57 163.367
R1240 B.n454 B.n57 163.367
R1241 B.n454 B.n453 163.367
R1242 B.n546 B.n23 163.367
R1243 B.n550 B.n23 163.367
R1244 B.n551 B.n550 163.367
R1245 B.n552 B.n551 163.367
R1246 B.n552 B.n21 163.367
R1247 B.n556 B.n21 163.367
R1248 B.n557 B.n556 163.367
R1249 B.n558 B.n557 163.367
R1250 B.n558 B.n19 163.367
R1251 B.n562 B.n19 163.367
R1252 B.n563 B.n562 163.367
R1253 B.n564 B.n563 163.367
R1254 B.n564 B.n17 163.367
R1255 B.n568 B.n17 163.367
R1256 B.n569 B.n568 163.367
R1257 B.n570 B.n569 163.367
R1258 B.n570 B.n15 163.367
R1259 B.n574 B.n15 163.367
R1260 B.n575 B.n574 163.367
R1261 B.n576 B.n575 163.367
R1262 B.n576 B.n13 163.367
R1263 B.n580 B.n13 163.367
R1264 B.n581 B.n580 163.367
R1265 B.n582 B.n581 163.367
R1266 B.n582 B.n11 163.367
R1267 B.n586 B.n11 163.367
R1268 B.n587 B.n586 163.367
R1269 B.n588 B.n587 163.367
R1270 B.n588 B.n9 163.367
R1271 B.n592 B.n9 163.367
R1272 B.n593 B.n592 163.367
R1273 B.n594 B.n593 163.367
R1274 B.n594 B.n7 163.367
R1275 B.n598 B.n7 163.367
R1276 B.n599 B.n598 163.367
R1277 B.n600 B.n599 163.367
R1278 B.n600 B.n5 163.367
R1279 B.n604 B.n5 163.367
R1280 B.n605 B.n604 163.367
R1281 B.n606 B.n605 163.367
R1282 B.n606 B.n3 163.367
R1283 B.n610 B.n3 163.367
R1284 B.n611 B.n610 163.367
R1285 B.n157 B.n2 163.367
R1286 B.n160 B.n157 163.367
R1287 B.n161 B.n160 163.367
R1288 B.n162 B.n161 163.367
R1289 B.n162 B.n155 163.367
R1290 B.n166 B.n155 163.367
R1291 B.n167 B.n166 163.367
R1292 B.n168 B.n167 163.367
R1293 B.n168 B.n153 163.367
R1294 B.n172 B.n153 163.367
R1295 B.n173 B.n172 163.367
R1296 B.n174 B.n173 163.367
R1297 B.n174 B.n151 163.367
R1298 B.n178 B.n151 163.367
R1299 B.n179 B.n178 163.367
R1300 B.n180 B.n179 163.367
R1301 B.n180 B.n149 163.367
R1302 B.n184 B.n149 163.367
R1303 B.n185 B.n184 163.367
R1304 B.n186 B.n185 163.367
R1305 B.n186 B.n147 163.367
R1306 B.n190 B.n147 163.367
R1307 B.n191 B.n190 163.367
R1308 B.n192 B.n191 163.367
R1309 B.n192 B.n145 163.367
R1310 B.n196 B.n145 163.367
R1311 B.n197 B.n196 163.367
R1312 B.n198 B.n197 163.367
R1313 B.n198 B.n143 163.367
R1314 B.n202 B.n143 163.367
R1315 B.n203 B.n202 163.367
R1316 B.n204 B.n203 163.367
R1317 B.n204 B.n141 163.367
R1318 B.n208 B.n141 163.367
R1319 B.n209 B.n208 163.367
R1320 B.n210 B.n209 163.367
R1321 B.n210 B.n139 163.367
R1322 B.n214 B.n139 163.367
R1323 B.n215 B.n214 163.367
R1324 B.n216 B.n215 163.367
R1325 B.n216 B.n137 163.367
R1326 B.n220 B.n137 163.367
R1327 B.n221 B.n220 163.367
R1328 B.n261 B.n123 59.5399
R1329 B.n276 B.n275 59.5399
R1330 B.n492 B.n45 59.5399
R1331 B.n506 B.n39 59.5399
R1332 B.n123 B.n122 39.952
R1333 B.n275 B.n274 39.952
R1334 B.n45 B.n44 39.952
R1335 B.n39 B.n38 39.952
R1336 B.n547 B.n24 34.4981
R1337 B.n451 B.n58 34.4981
R1338 B.n318 B.n317 34.4981
R1339 B.n223 B.n136 34.4981
R1340 B B.n613 18.0485
R1341 B.n548 B.n547 10.6151
R1342 B.n549 B.n548 10.6151
R1343 B.n549 B.n22 10.6151
R1344 B.n553 B.n22 10.6151
R1345 B.n554 B.n553 10.6151
R1346 B.n555 B.n554 10.6151
R1347 B.n555 B.n20 10.6151
R1348 B.n559 B.n20 10.6151
R1349 B.n560 B.n559 10.6151
R1350 B.n561 B.n560 10.6151
R1351 B.n561 B.n18 10.6151
R1352 B.n565 B.n18 10.6151
R1353 B.n566 B.n565 10.6151
R1354 B.n567 B.n566 10.6151
R1355 B.n567 B.n16 10.6151
R1356 B.n571 B.n16 10.6151
R1357 B.n572 B.n571 10.6151
R1358 B.n573 B.n572 10.6151
R1359 B.n573 B.n14 10.6151
R1360 B.n577 B.n14 10.6151
R1361 B.n578 B.n577 10.6151
R1362 B.n579 B.n578 10.6151
R1363 B.n579 B.n12 10.6151
R1364 B.n583 B.n12 10.6151
R1365 B.n584 B.n583 10.6151
R1366 B.n585 B.n584 10.6151
R1367 B.n585 B.n10 10.6151
R1368 B.n589 B.n10 10.6151
R1369 B.n590 B.n589 10.6151
R1370 B.n591 B.n590 10.6151
R1371 B.n591 B.n8 10.6151
R1372 B.n595 B.n8 10.6151
R1373 B.n596 B.n595 10.6151
R1374 B.n597 B.n596 10.6151
R1375 B.n597 B.n6 10.6151
R1376 B.n601 B.n6 10.6151
R1377 B.n602 B.n601 10.6151
R1378 B.n603 B.n602 10.6151
R1379 B.n603 B.n4 10.6151
R1380 B.n607 B.n4 10.6151
R1381 B.n608 B.n607 10.6151
R1382 B.n609 B.n608 10.6151
R1383 B.n609 B.n0 10.6151
R1384 B.n543 B.n24 10.6151
R1385 B.n543 B.n542 10.6151
R1386 B.n542 B.n541 10.6151
R1387 B.n541 B.n26 10.6151
R1388 B.n537 B.n26 10.6151
R1389 B.n537 B.n536 10.6151
R1390 B.n536 B.n535 10.6151
R1391 B.n535 B.n28 10.6151
R1392 B.n531 B.n28 10.6151
R1393 B.n531 B.n530 10.6151
R1394 B.n530 B.n529 10.6151
R1395 B.n529 B.n30 10.6151
R1396 B.n525 B.n30 10.6151
R1397 B.n525 B.n524 10.6151
R1398 B.n524 B.n523 10.6151
R1399 B.n523 B.n32 10.6151
R1400 B.n519 B.n32 10.6151
R1401 B.n519 B.n518 10.6151
R1402 B.n518 B.n517 10.6151
R1403 B.n517 B.n34 10.6151
R1404 B.n513 B.n34 10.6151
R1405 B.n513 B.n512 10.6151
R1406 B.n512 B.n511 10.6151
R1407 B.n511 B.n36 10.6151
R1408 B.n507 B.n36 10.6151
R1409 B.n505 B.n504 10.6151
R1410 B.n504 B.n40 10.6151
R1411 B.n500 B.n40 10.6151
R1412 B.n500 B.n499 10.6151
R1413 B.n499 B.n498 10.6151
R1414 B.n498 B.n42 10.6151
R1415 B.n494 B.n42 10.6151
R1416 B.n494 B.n493 10.6151
R1417 B.n491 B.n46 10.6151
R1418 B.n487 B.n46 10.6151
R1419 B.n487 B.n486 10.6151
R1420 B.n486 B.n485 10.6151
R1421 B.n485 B.n48 10.6151
R1422 B.n481 B.n48 10.6151
R1423 B.n481 B.n480 10.6151
R1424 B.n480 B.n479 10.6151
R1425 B.n479 B.n50 10.6151
R1426 B.n475 B.n50 10.6151
R1427 B.n475 B.n474 10.6151
R1428 B.n474 B.n473 10.6151
R1429 B.n473 B.n52 10.6151
R1430 B.n469 B.n52 10.6151
R1431 B.n469 B.n468 10.6151
R1432 B.n468 B.n467 10.6151
R1433 B.n467 B.n54 10.6151
R1434 B.n463 B.n54 10.6151
R1435 B.n463 B.n462 10.6151
R1436 B.n462 B.n461 10.6151
R1437 B.n461 B.n56 10.6151
R1438 B.n457 B.n56 10.6151
R1439 B.n457 B.n456 10.6151
R1440 B.n456 B.n455 10.6151
R1441 B.n455 B.n58 10.6151
R1442 B.n451 B.n450 10.6151
R1443 B.n450 B.n449 10.6151
R1444 B.n449 B.n60 10.6151
R1445 B.n445 B.n60 10.6151
R1446 B.n445 B.n444 10.6151
R1447 B.n444 B.n443 10.6151
R1448 B.n443 B.n62 10.6151
R1449 B.n439 B.n62 10.6151
R1450 B.n439 B.n438 10.6151
R1451 B.n438 B.n437 10.6151
R1452 B.n437 B.n64 10.6151
R1453 B.n433 B.n64 10.6151
R1454 B.n433 B.n432 10.6151
R1455 B.n432 B.n431 10.6151
R1456 B.n431 B.n66 10.6151
R1457 B.n427 B.n66 10.6151
R1458 B.n427 B.n426 10.6151
R1459 B.n426 B.n425 10.6151
R1460 B.n425 B.n68 10.6151
R1461 B.n421 B.n68 10.6151
R1462 B.n421 B.n420 10.6151
R1463 B.n420 B.n419 10.6151
R1464 B.n419 B.n70 10.6151
R1465 B.n415 B.n70 10.6151
R1466 B.n415 B.n414 10.6151
R1467 B.n414 B.n413 10.6151
R1468 B.n413 B.n72 10.6151
R1469 B.n409 B.n72 10.6151
R1470 B.n409 B.n408 10.6151
R1471 B.n408 B.n407 10.6151
R1472 B.n407 B.n74 10.6151
R1473 B.n403 B.n74 10.6151
R1474 B.n403 B.n402 10.6151
R1475 B.n402 B.n401 10.6151
R1476 B.n401 B.n76 10.6151
R1477 B.n397 B.n76 10.6151
R1478 B.n397 B.n396 10.6151
R1479 B.n396 B.n395 10.6151
R1480 B.n395 B.n78 10.6151
R1481 B.n391 B.n78 10.6151
R1482 B.n391 B.n390 10.6151
R1483 B.n390 B.n389 10.6151
R1484 B.n389 B.n80 10.6151
R1485 B.n385 B.n80 10.6151
R1486 B.n385 B.n384 10.6151
R1487 B.n384 B.n383 10.6151
R1488 B.n383 B.n82 10.6151
R1489 B.n379 B.n82 10.6151
R1490 B.n379 B.n378 10.6151
R1491 B.n378 B.n377 10.6151
R1492 B.n377 B.n84 10.6151
R1493 B.n373 B.n84 10.6151
R1494 B.n373 B.n372 10.6151
R1495 B.n372 B.n371 10.6151
R1496 B.n371 B.n86 10.6151
R1497 B.n367 B.n86 10.6151
R1498 B.n367 B.n366 10.6151
R1499 B.n366 B.n365 10.6151
R1500 B.n365 B.n88 10.6151
R1501 B.n361 B.n88 10.6151
R1502 B.n361 B.n360 10.6151
R1503 B.n360 B.n359 10.6151
R1504 B.n359 B.n90 10.6151
R1505 B.n355 B.n90 10.6151
R1506 B.n355 B.n354 10.6151
R1507 B.n354 B.n353 10.6151
R1508 B.n353 B.n92 10.6151
R1509 B.n349 B.n92 10.6151
R1510 B.n349 B.n348 10.6151
R1511 B.n348 B.n347 10.6151
R1512 B.n347 B.n94 10.6151
R1513 B.n343 B.n94 10.6151
R1514 B.n343 B.n342 10.6151
R1515 B.n342 B.n341 10.6151
R1516 B.n341 B.n96 10.6151
R1517 B.n337 B.n96 10.6151
R1518 B.n337 B.n336 10.6151
R1519 B.n336 B.n335 10.6151
R1520 B.n335 B.n98 10.6151
R1521 B.n331 B.n98 10.6151
R1522 B.n331 B.n330 10.6151
R1523 B.n330 B.n329 10.6151
R1524 B.n329 B.n100 10.6151
R1525 B.n325 B.n100 10.6151
R1526 B.n325 B.n324 10.6151
R1527 B.n324 B.n323 10.6151
R1528 B.n323 B.n102 10.6151
R1529 B.n319 B.n102 10.6151
R1530 B.n319 B.n318 10.6151
R1531 B.n158 B.n1 10.6151
R1532 B.n159 B.n158 10.6151
R1533 B.n159 B.n156 10.6151
R1534 B.n163 B.n156 10.6151
R1535 B.n164 B.n163 10.6151
R1536 B.n165 B.n164 10.6151
R1537 B.n165 B.n154 10.6151
R1538 B.n169 B.n154 10.6151
R1539 B.n170 B.n169 10.6151
R1540 B.n171 B.n170 10.6151
R1541 B.n171 B.n152 10.6151
R1542 B.n175 B.n152 10.6151
R1543 B.n176 B.n175 10.6151
R1544 B.n177 B.n176 10.6151
R1545 B.n177 B.n150 10.6151
R1546 B.n181 B.n150 10.6151
R1547 B.n182 B.n181 10.6151
R1548 B.n183 B.n182 10.6151
R1549 B.n183 B.n148 10.6151
R1550 B.n187 B.n148 10.6151
R1551 B.n188 B.n187 10.6151
R1552 B.n189 B.n188 10.6151
R1553 B.n189 B.n146 10.6151
R1554 B.n193 B.n146 10.6151
R1555 B.n194 B.n193 10.6151
R1556 B.n195 B.n194 10.6151
R1557 B.n195 B.n144 10.6151
R1558 B.n199 B.n144 10.6151
R1559 B.n200 B.n199 10.6151
R1560 B.n201 B.n200 10.6151
R1561 B.n201 B.n142 10.6151
R1562 B.n205 B.n142 10.6151
R1563 B.n206 B.n205 10.6151
R1564 B.n207 B.n206 10.6151
R1565 B.n207 B.n140 10.6151
R1566 B.n211 B.n140 10.6151
R1567 B.n212 B.n211 10.6151
R1568 B.n213 B.n212 10.6151
R1569 B.n213 B.n138 10.6151
R1570 B.n217 B.n138 10.6151
R1571 B.n218 B.n217 10.6151
R1572 B.n219 B.n218 10.6151
R1573 B.n219 B.n136 10.6151
R1574 B.n224 B.n223 10.6151
R1575 B.n225 B.n224 10.6151
R1576 B.n225 B.n134 10.6151
R1577 B.n229 B.n134 10.6151
R1578 B.n230 B.n229 10.6151
R1579 B.n231 B.n230 10.6151
R1580 B.n231 B.n132 10.6151
R1581 B.n235 B.n132 10.6151
R1582 B.n236 B.n235 10.6151
R1583 B.n237 B.n236 10.6151
R1584 B.n237 B.n130 10.6151
R1585 B.n241 B.n130 10.6151
R1586 B.n242 B.n241 10.6151
R1587 B.n243 B.n242 10.6151
R1588 B.n243 B.n128 10.6151
R1589 B.n247 B.n128 10.6151
R1590 B.n248 B.n247 10.6151
R1591 B.n249 B.n248 10.6151
R1592 B.n249 B.n126 10.6151
R1593 B.n253 B.n126 10.6151
R1594 B.n254 B.n253 10.6151
R1595 B.n255 B.n254 10.6151
R1596 B.n255 B.n124 10.6151
R1597 B.n259 B.n124 10.6151
R1598 B.n260 B.n259 10.6151
R1599 B.n262 B.n120 10.6151
R1600 B.n266 B.n120 10.6151
R1601 B.n267 B.n266 10.6151
R1602 B.n268 B.n267 10.6151
R1603 B.n268 B.n118 10.6151
R1604 B.n272 B.n118 10.6151
R1605 B.n273 B.n272 10.6151
R1606 B.n277 B.n273 10.6151
R1607 B.n281 B.n116 10.6151
R1608 B.n282 B.n281 10.6151
R1609 B.n283 B.n282 10.6151
R1610 B.n283 B.n114 10.6151
R1611 B.n287 B.n114 10.6151
R1612 B.n288 B.n287 10.6151
R1613 B.n289 B.n288 10.6151
R1614 B.n289 B.n112 10.6151
R1615 B.n293 B.n112 10.6151
R1616 B.n294 B.n293 10.6151
R1617 B.n295 B.n294 10.6151
R1618 B.n295 B.n110 10.6151
R1619 B.n299 B.n110 10.6151
R1620 B.n300 B.n299 10.6151
R1621 B.n301 B.n300 10.6151
R1622 B.n301 B.n108 10.6151
R1623 B.n305 B.n108 10.6151
R1624 B.n306 B.n305 10.6151
R1625 B.n307 B.n306 10.6151
R1626 B.n307 B.n106 10.6151
R1627 B.n311 B.n106 10.6151
R1628 B.n312 B.n311 10.6151
R1629 B.n313 B.n312 10.6151
R1630 B.n313 B.n104 10.6151
R1631 B.n317 B.n104 10.6151
R1632 B.n613 B.n0 8.11757
R1633 B.n613 B.n1 8.11757
R1634 B.n506 B.n505 6.5566
R1635 B.n493 B.n492 6.5566
R1636 B.n262 B.n261 6.5566
R1637 B.n277 B.n276 6.5566
R1638 B.n507 B.n506 4.05904
R1639 B.n492 B.n491 4.05904
R1640 B.n261 B.n260 4.05904
R1641 B.n276 B.n116 4.05904
C0 VP w_n3442_n2302# 7.44673f
C1 VP VDD1 5.91518f
C2 VTAIL B 2.22351f
C3 VN VP 6.12771f
C4 VDD2 B 1.80898f
C5 VTAIL w_n3442_n2302# 2.32217f
C6 VTAIL VDD1 7.58682f
C7 VDD2 w_n3442_n2302# 2.17349f
C8 VDD2 VDD1 1.60599f
C9 VN VTAIL 6.23244f
C10 VN VDD2 5.59719f
C11 B w_n3442_n2302# 7.59291f
C12 VTAIL VP 6.2467f
C13 B VDD1 1.72494f
C14 VDD2 VP 0.471865f
C15 VDD1 w_n3442_n2302# 2.07505f
C16 VN B 0.99803f
C17 VN w_n3442_n2302# 7.001279f
C18 VN VDD1 0.151126f
C19 VTAIL VDD2 7.63247f
C20 VP B 1.74227f
C21 VDD2 VSUBS 1.562983f
C22 VDD1 VSUBS 1.425833f
C23 VTAIL VSUBS 0.597792f
C24 VN VSUBS 5.95088f
C25 VP VSUBS 2.756588f
C26 B VSUBS 3.834599f
C27 w_n3442_n2302# VSUBS 98.6753f
C28 B.n0 VSUBS 0.006762f
C29 B.n1 VSUBS 0.006762f
C30 B.n2 VSUBS 0.01f
C31 B.n3 VSUBS 0.007663f
C32 B.n4 VSUBS 0.007663f
C33 B.n5 VSUBS 0.007663f
C34 B.n6 VSUBS 0.007663f
C35 B.n7 VSUBS 0.007663f
C36 B.n8 VSUBS 0.007663f
C37 B.n9 VSUBS 0.007663f
C38 B.n10 VSUBS 0.007663f
C39 B.n11 VSUBS 0.007663f
C40 B.n12 VSUBS 0.007663f
C41 B.n13 VSUBS 0.007663f
C42 B.n14 VSUBS 0.007663f
C43 B.n15 VSUBS 0.007663f
C44 B.n16 VSUBS 0.007663f
C45 B.n17 VSUBS 0.007663f
C46 B.n18 VSUBS 0.007663f
C47 B.n19 VSUBS 0.007663f
C48 B.n20 VSUBS 0.007663f
C49 B.n21 VSUBS 0.007663f
C50 B.n22 VSUBS 0.007663f
C51 B.n23 VSUBS 0.007663f
C52 B.n24 VSUBS 0.018815f
C53 B.n25 VSUBS 0.007663f
C54 B.n26 VSUBS 0.007663f
C55 B.n27 VSUBS 0.007663f
C56 B.n28 VSUBS 0.007663f
C57 B.n29 VSUBS 0.007663f
C58 B.n30 VSUBS 0.007663f
C59 B.n31 VSUBS 0.007663f
C60 B.n32 VSUBS 0.007663f
C61 B.n33 VSUBS 0.007663f
C62 B.n34 VSUBS 0.007663f
C63 B.n35 VSUBS 0.007663f
C64 B.n36 VSUBS 0.007663f
C65 B.n37 VSUBS 0.007663f
C66 B.t4 VSUBS 0.111052f
C67 B.t5 VSUBS 0.132259f
C68 B.t3 VSUBS 0.580478f
C69 B.n38 VSUBS 0.227177f
C70 B.n39 VSUBS 0.180761f
C71 B.n40 VSUBS 0.007663f
C72 B.n41 VSUBS 0.007663f
C73 B.n42 VSUBS 0.007663f
C74 B.n43 VSUBS 0.007663f
C75 B.t10 VSUBS 0.111054f
C76 B.t11 VSUBS 0.132261f
C77 B.t9 VSUBS 0.580478f
C78 B.n44 VSUBS 0.227175f
C79 B.n45 VSUBS 0.180759f
C80 B.n46 VSUBS 0.007663f
C81 B.n47 VSUBS 0.007663f
C82 B.n48 VSUBS 0.007663f
C83 B.n49 VSUBS 0.007663f
C84 B.n50 VSUBS 0.007663f
C85 B.n51 VSUBS 0.007663f
C86 B.n52 VSUBS 0.007663f
C87 B.n53 VSUBS 0.007663f
C88 B.n54 VSUBS 0.007663f
C89 B.n55 VSUBS 0.007663f
C90 B.n56 VSUBS 0.007663f
C91 B.n57 VSUBS 0.007663f
C92 B.n58 VSUBS 0.018815f
C93 B.n59 VSUBS 0.007663f
C94 B.n60 VSUBS 0.007663f
C95 B.n61 VSUBS 0.007663f
C96 B.n62 VSUBS 0.007663f
C97 B.n63 VSUBS 0.007663f
C98 B.n64 VSUBS 0.007663f
C99 B.n65 VSUBS 0.007663f
C100 B.n66 VSUBS 0.007663f
C101 B.n67 VSUBS 0.007663f
C102 B.n68 VSUBS 0.007663f
C103 B.n69 VSUBS 0.007663f
C104 B.n70 VSUBS 0.007663f
C105 B.n71 VSUBS 0.007663f
C106 B.n72 VSUBS 0.007663f
C107 B.n73 VSUBS 0.007663f
C108 B.n74 VSUBS 0.007663f
C109 B.n75 VSUBS 0.007663f
C110 B.n76 VSUBS 0.007663f
C111 B.n77 VSUBS 0.007663f
C112 B.n78 VSUBS 0.007663f
C113 B.n79 VSUBS 0.007663f
C114 B.n80 VSUBS 0.007663f
C115 B.n81 VSUBS 0.007663f
C116 B.n82 VSUBS 0.007663f
C117 B.n83 VSUBS 0.007663f
C118 B.n84 VSUBS 0.007663f
C119 B.n85 VSUBS 0.007663f
C120 B.n86 VSUBS 0.007663f
C121 B.n87 VSUBS 0.007663f
C122 B.n88 VSUBS 0.007663f
C123 B.n89 VSUBS 0.007663f
C124 B.n90 VSUBS 0.007663f
C125 B.n91 VSUBS 0.007663f
C126 B.n92 VSUBS 0.007663f
C127 B.n93 VSUBS 0.007663f
C128 B.n94 VSUBS 0.007663f
C129 B.n95 VSUBS 0.007663f
C130 B.n96 VSUBS 0.007663f
C131 B.n97 VSUBS 0.007663f
C132 B.n98 VSUBS 0.007663f
C133 B.n99 VSUBS 0.007663f
C134 B.n100 VSUBS 0.007663f
C135 B.n101 VSUBS 0.007663f
C136 B.n102 VSUBS 0.007663f
C137 B.n103 VSUBS 0.018376f
C138 B.n104 VSUBS 0.007663f
C139 B.n105 VSUBS 0.007663f
C140 B.n106 VSUBS 0.007663f
C141 B.n107 VSUBS 0.007663f
C142 B.n108 VSUBS 0.007663f
C143 B.n109 VSUBS 0.007663f
C144 B.n110 VSUBS 0.007663f
C145 B.n111 VSUBS 0.007663f
C146 B.n112 VSUBS 0.007663f
C147 B.n113 VSUBS 0.007663f
C148 B.n114 VSUBS 0.007663f
C149 B.n115 VSUBS 0.007663f
C150 B.n116 VSUBS 0.005297f
C151 B.n117 VSUBS 0.007663f
C152 B.n118 VSUBS 0.007663f
C153 B.n119 VSUBS 0.007663f
C154 B.n120 VSUBS 0.007663f
C155 B.n121 VSUBS 0.007663f
C156 B.t8 VSUBS 0.111052f
C157 B.t7 VSUBS 0.132259f
C158 B.t6 VSUBS 0.580478f
C159 B.n122 VSUBS 0.227177f
C160 B.n123 VSUBS 0.180761f
C161 B.n124 VSUBS 0.007663f
C162 B.n125 VSUBS 0.007663f
C163 B.n126 VSUBS 0.007663f
C164 B.n127 VSUBS 0.007663f
C165 B.n128 VSUBS 0.007663f
C166 B.n129 VSUBS 0.007663f
C167 B.n130 VSUBS 0.007663f
C168 B.n131 VSUBS 0.007663f
C169 B.n132 VSUBS 0.007663f
C170 B.n133 VSUBS 0.007663f
C171 B.n134 VSUBS 0.007663f
C172 B.n135 VSUBS 0.007663f
C173 B.n136 VSUBS 0.018376f
C174 B.n137 VSUBS 0.007663f
C175 B.n138 VSUBS 0.007663f
C176 B.n139 VSUBS 0.007663f
C177 B.n140 VSUBS 0.007663f
C178 B.n141 VSUBS 0.007663f
C179 B.n142 VSUBS 0.007663f
C180 B.n143 VSUBS 0.007663f
C181 B.n144 VSUBS 0.007663f
C182 B.n145 VSUBS 0.007663f
C183 B.n146 VSUBS 0.007663f
C184 B.n147 VSUBS 0.007663f
C185 B.n148 VSUBS 0.007663f
C186 B.n149 VSUBS 0.007663f
C187 B.n150 VSUBS 0.007663f
C188 B.n151 VSUBS 0.007663f
C189 B.n152 VSUBS 0.007663f
C190 B.n153 VSUBS 0.007663f
C191 B.n154 VSUBS 0.007663f
C192 B.n155 VSUBS 0.007663f
C193 B.n156 VSUBS 0.007663f
C194 B.n157 VSUBS 0.007663f
C195 B.n158 VSUBS 0.007663f
C196 B.n159 VSUBS 0.007663f
C197 B.n160 VSUBS 0.007663f
C198 B.n161 VSUBS 0.007663f
C199 B.n162 VSUBS 0.007663f
C200 B.n163 VSUBS 0.007663f
C201 B.n164 VSUBS 0.007663f
C202 B.n165 VSUBS 0.007663f
C203 B.n166 VSUBS 0.007663f
C204 B.n167 VSUBS 0.007663f
C205 B.n168 VSUBS 0.007663f
C206 B.n169 VSUBS 0.007663f
C207 B.n170 VSUBS 0.007663f
C208 B.n171 VSUBS 0.007663f
C209 B.n172 VSUBS 0.007663f
C210 B.n173 VSUBS 0.007663f
C211 B.n174 VSUBS 0.007663f
C212 B.n175 VSUBS 0.007663f
C213 B.n176 VSUBS 0.007663f
C214 B.n177 VSUBS 0.007663f
C215 B.n178 VSUBS 0.007663f
C216 B.n179 VSUBS 0.007663f
C217 B.n180 VSUBS 0.007663f
C218 B.n181 VSUBS 0.007663f
C219 B.n182 VSUBS 0.007663f
C220 B.n183 VSUBS 0.007663f
C221 B.n184 VSUBS 0.007663f
C222 B.n185 VSUBS 0.007663f
C223 B.n186 VSUBS 0.007663f
C224 B.n187 VSUBS 0.007663f
C225 B.n188 VSUBS 0.007663f
C226 B.n189 VSUBS 0.007663f
C227 B.n190 VSUBS 0.007663f
C228 B.n191 VSUBS 0.007663f
C229 B.n192 VSUBS 0.007663f
C230 B.n193 VSUBS 0.007663f
C231 B.n194 VSUBS 0.007663f
C232 B.n195 VSUBS 0.007663f
C233 B.n196 VSUBS 0.007663f
C234 B.n197 VSUBS 0.007663f
C235 B.n198 VSUBS 0.007663f
C236 B.n199 VSUBS 0.007663f
C237 B.n200 VSUBS 0.007663f
C238 B.n201 VSUBS 0.007663f
C239 B.n202 VSUBS 0.007663f
C240 B.n203 VSUBS 0.007663f
C241 B.n204 VSUBS 0.007663f
C242 B.n205 VSUBS 0.007663f
C243 B.n206 VSUBS 0.007663f
C244 B.n207 VSUBS 0.007663f
C245 B.n208 VSUBS 0.007663f
C246 B.n209 VSUBS 0.007663f
C247 B.n210 VSUBS 0.007663f
C248 B.n211 VSUBS 0.007663f
C249 B.n212 VSUBS 0.007663f
C250 B.n213 VSUBS 0.007663f
C251 B.n214 VSUBS 0.007663f
C252 B.n215 VSUBS 0.007663f
C253 B.n216 VSUBS 0.007663f
C254 B.n217 VSUBS 0.007663f
C255 B.n218 VSUBS 0.007663f
C256 B.n219 VSUBS 0.007663f
C257 B.n220 VSUBS 0.007663f
C258 B.n221 VSUBS 0.018376f
C259 B.n222 VSUBS 0.018815f
C260 B.n223 VSUBS 0.018815f
C261 B.n224 VSUBS 0.007663f
C262 B.n225 VSUBS 0.007663f
C263 B.n226 VSUBS 0.007663f
C264 B.n227 VSUBS 0.007663f
C265 B.n228 VSUBS 0.007663f
C266 B.n229 VSUBS 0.007663f
C267 B.n230 VSUBS 0.007663f
C268 B.n231 VSUBS 0.007663f
C269 B.n232 VSUBS 0.007663f
C270 B.n233 VSUBS 0.007663f
C271 B.n234 VSUBS 0.007663f
C272 B.n235 VSUBS 0.007663f
C273 B.n236 VSUBS 0.007663f
C274 B.n237 VSUBS 0.007663f
C275 B.n238 VSUBS 0.007663f
C276 B.n239 VSUBS 0.007663f
C277 B.n240 VSUBS 0.007663f
C278 B.n241 VSUBS 0.007663f
C279 B.n242 VSUBS 0.007663f
C280 B.n243 VSUBS 0.007663f
C281 B.n244 VSUBS 0.007663f
C282 B.n245 VSUBS 0.007663f
C283 B.n246 VSUBS 0.007663f
C284 B.n247 VSUBS 0.007663f
C285 B.n248 VSUBS 0.007663f
C286 B.n249 VSUBS 0.007663f
C287 B.n250 VSUBS 0.007663f
C288 B.n251 VSUBS 0.007663f
C289 B.n252 VSUBS 0.007663f
C290 B.n253 VSUBS 0.007663f
C291 B.n254 VSUBS 0.007663f
C292 B.n255 VSUBS 0.007663f
C293 B.n256 VSUBS 0.007663f
C294 B.n257 VSUBS 0.007663f
C295 B.n258 VSUBS 0.007663f
C296 B.n259 VSUBS 0.007663f
C297 B.n260 VSUBS 0.005297f
C298 B.n261 VSUBS 0.017756f
C299 B.n262 VSUBS 0.006198f
C300 B.n263 VSUBS 0.007663f
C301 B.n264 VSUBS 0.007663f
C302 B.n265 VSUBS 0.007663f
C303 B.n266 VSUBS 0.007663f
C304 B.n267 VSUBS 0.007663f
C305 B.n268 VSUBS 0.007663f
C306 B.n269 VSUBS 0.007663f
C307 B.n270 VSUBS 0.007663f
C308 B.n271 VSUBS 0.007663f
C309 B.n272 VSUBS 0.007663f
C310 B.n273 VSUBS 0.007663f
C311 B.t2 VSUBS 0.111054f
C312 B.t1 VSUBS 0.132261f
C313 B.t0 VSUBS 0.580478f
C314 B.n274 VSUBS 0.227175f
C315 B.n275 VSUBS 0.180759f
C316 B.n276 VSUBS 0.017756f
C317 B.n277 VSUBS 0.006198f
C318 B.n278 VSUBS 0.007663f
C319 B.n279 VSUBS 0.007663f
C320 B.n280 VSUBS 0.007663f
C321 B.n281 VSUBS 0.007663f
C322 B.n282 VSUBS 0.007663f
C323 B.n283 VSUBS 0.007663f
C324 B.n284 VSUBS 0.007663f
C325 B.n285 VSUBS 0.007663f
C326 B.n286 VSUBS 0.007663f
C327 B.n287 VSUBS 0.007663f
C328 B.n288 VSUBS 0.007663f
C329 B.n289 VSUBS 0.007663f
C330 B.n290 VSUBS 0.007663f
C331 B.n291 VSUBS 0.007663f
C332 B.n292 VSUBS 0.007663f
C333 B.n293 VSUBS 0.007663f
C334 B.n294 VSUBS 0.007663f
C335 B.n295 VSUBS 0.007663f
C336 B.n296 VSUBS 0.007663f
C337 B.n297 VSUBS 0.007663f
C338 B.n298 VSUBS 0.007663f
C339 B.n299 VSUBS 0.007663f
C340 B.n300 VSUBS 0.007663f
C341 B.n301 VSUBS 0.007663f
C342 B.n302 VSUBS 0.007663f
C343 B.n303 VSUBS 0.007663f
C344 B.n304 VSUBS 0.007663f
C345 B.n305 VSUBS 0.007663f
C346 B.n306 VSUBS 0.007663f
C347 B.n307 VSUBS 0.007663f
C348 B.n308 VSUBS 0.007663f
C349 B.n309 VSUBS 0.007663f
C350 B.n310 VSUBS 0.007663f
C351 B.n311 VSUBS 0.007663f
C352 B.n312 VSUBS 0.007663f
C353 B.n313 VSUBS 0.007663f
C354 B.n314 VSUBS 0.007663f
C355 B.n315 VSUBS 0.007663f
C356 B.n316 VSUBS 0.018815f
C357 B.n317 VSUBS 0.017958f
C358 B.n318 VSUBS 0.019233f
C359 B.n319 VSUBS 0.007663f
C360 B.n320 VSUBS 0.007663f
C361 B.n321 VSUBS 0.007663f
C362 B.n322 VSUBS 0.007663f
C363 B.n323 VSUBS 0.007663f
C364 B.n324 VSUBS 0.007663f
C365 B.n325 VSUBS 0.007663f
C366 B.n326 VSUBS 0.007663f
C367 B.n327 VSUBS 0.007663f
C368 B.n328 VSUBS 0.007663f
C369 B.n329 VSUBS 0.007663f
C370 B.n330 VSUBS 0.007663f
C371 B.n331 VSUBS 0.007663f
C372 B.n332 VSUBS 0.007663f
C373 B.n333 VSUBS 0.007663f
C374 B.n334 VSUBS 0.007663f
C375 B.n335 VSUBS 0.007663f
C376 B.n336 VSUBS 0.007663f
C377 B.n337 VSUBS 0.007663f
C378 B.n338 VSUBS 0.007663f
C379 B.n339 VSUBS 0.007663f
C380 B.n340 VSUBS 0.007663f
C381 B.n341 VSUBS 0.007663f
C382 B.n342 VSUBS 0.007663f
C383 B.n343 VSUBS 0.007663f
C384 B.n344 VSUBS 0.007663f
C385 B.n345 VSUBS 0.007663f
C386 B.n346 VSUBS 0.007663f
C387 B.n347 VSUBS 0.007663f
C388 B.n348 VSUBS 0.007663f
C389 B.n349 VSUBS 0.007663f
C390 B.n350 VSUBS 0.007663f
C391 B.n351 VSUBS 0.007663f
C392 B.n352 VSUBS 0.007663f
C393 B.n353 VSUBS 0.007663f
C394 B.n354 VSUBS 0.007663f
C395 B.n355 VSUBS 0.007663f
C396 B.n356 VSUBS 0.007663f
C397 B.n357 VSUBS 0.007663f
C398 B.n358 VSUBS 0.007663f
C399 B.n359 VSUBS 0.007663f
C400 B.n360 VSUBS 0.007663f
C401 B.n361 VSUBS 0.007663f
C402 B.n362 VSUBS 0.007663f
C403 B.n363 VSUBS 0.007663f
C404 B.n364 VSUBS 0.007663f
C405 B.n365 VSUBS 0.007663f
C406 B.n366 VSUBS 0.007663f
C407 B.n367 VSUBS 0.007663f
C408 B.n368 VSUBS 0.007663f
C409 B.n369 VSUBS 0.007663f
C410 B.n370 VSUBS 0.007663f
C411 B.n371 VSUBS 0.007663f
C412 B.n372 VSUBS 0.007663f
C413 B.n373 VSUBS 0.007663f
C414 B.n374 VSUBS 0.007663f
C415 B.n375 VSUBS 0.007663f
C416 B.n376 VSUBS 0.007663f
C417 B.n377 VSUBS 0.007663f
C418 B.n378 VSUBS 0.007663f
C419 B.n379 VSUBS 0.007663f
C420 B.n380 VSUBS 0.007663f
C421 B.n381 VSUBS 0.007663f
C422 B.n382 VSUBS 0.007663f
C423 B.n383 VSUBS 0.007663f
C424 B.n384 VSUBS 0.007663f
C425 B.n385 VSUBS 0.007663f
C426 B.n386 VSUBS 0.007663f
C427 B.n387 VSUBS 0.007663f
C428 B.n388 VSUBS 0.007663f
C429 B.n389 VSUBS 0.007663f
C430 B.n390 VSUBS 0.007663f
C431 B.n391 VSUBS 0.007663f
C432 B.n392 VSUBS 0.007663f
C433 B.n393 VSUBS 0.007663f
C434 B.n394 VSUBS 0.007663f
C435 B.n395 VSUBS 0.007663f
C436 B.n396 VSUBS 0.007663f
C437 B.n397 VSUBS 0.007663f
C438 B.n398 VSUBS 0.007663f
C439 B.n399 VSUBS 0.007663f
C440 B.n400 VSUBS 0.007663f
C441 B.n401 VSUBS 0.007663f
C442 B.n402 VSUBS 0.007663f
C443 B.n403 VSUBS 0.007663f
C444 B.n404 VSUBS 0.007663f
C445 B.n405 VSUBS 0.007663f
C446 B.n406 VSUBS 0.007663f
C447 B.n407 VSUBS 0.007663f
C448 B.n408 VSUBS 0.007663f
C449 B.n409 VSUBS 0.007663f
C450 B.n410 VSUBS 0.007663f
C451 B.n411 VSUBS 0.007663f
C452 B.n412 VSUBS 0.007663f
C453 B.n413 VSUBS 0.007663f
C454 B.n414 VSUBS 0.007663f
C455 B.n415 VSUBS 0.007663f
C456 B.n416 VSUBS 0.007663f
C457 B.n417 VSUBS 0.007663f
C458 B.n418 VSUBS 0.007663f
C459 B.n419 VSUBS 0.007663f
C460 B.n420 VSUBS 0.007663f
C461 B.n421 VSUBS 0.007663f
C462 B.n422 VSUBS 0.007663f
C463 B.n423 VSUBS 0.007663f
C464 B.n424 VSUBS 0.007663f
C465 B.n425 VSUBS 0.007663f
C466 B.n426 VSUBS 0.007663f
C467 B.n427 VSUBS 0.007663f
C468 B.n428 VSUBS 0.007663f
C469 B.n429 VSUBS 0.007663f
C470 B.n430 VSUBS 0.007663f
C471 B.n431 VSUBS 0.007663f
C472 B.n432 VSUBS 0.007663f
C473 B.n433 VSUBS 0.007663f
C474 B.n434 VSUBS 0.007663f
C475 B.n435 VSUBS 0.007663f
C476 B.n436 VSUBS 0.007663f
C477 B.n437 VSUBS 0.007663f
C478 B.n438 VSUBS 0.007663f
C479 B.n439 VSUBS 0.007663f
C480 B.n440 VSUBS 0.007663f
C481 B.n441 VSUBS 0.007663f
C482 B.n442 VSUBS 0.007663f
C483 B.n443 VSUBS 0.007663f
C484 B.n444 VSUBS 0.007663f
C485 B.n445 VSUBS 0.007663f
C486 B.n446 VSUBS 0.007663f
C487 B.n447 VSUBS 0.007663f
C488 B.n448 VSUBS 0.007663f
C489 B.n449 VSUBS 0.007663f
C490 B.n450 VSUBS 0.007663f
C491 B.n451 VSUBS 0.018376f
C492 B.n452 VSUBS 0.018376f
C493 B.n453 VSUBS 0.018815f
C494 B.n454 VSUBS 0.007663f
C495 B.n455 VSUBS 0.007663f
C496 B.n456 VSUBS 0.007663f
C497 B.n457 VSUBS 0.007663f
C498 B.n458 VSUBS 0.007663f
C499 B.n459 VSUBS 0.007663f
C500 B.n460 VSUBS 0.007663f
C501 B.n461 VSUBS 0.007663f
C502 B.n462 VSUBS 0.007663f
C503 B.n463 VSUBS 0.007663f
C504 B.n464 VSUBS 0.007663f
C505 B.n465 VSUBS 0.007663f
C506 B.n466 VSUBS 0.007663f
C507 B.n467 VSUBS 0.007663f
C508 B.n468 VSUBS 0.007663f
C509 B.n469 VSUBS 0.007663f
C510 B.n470 VSUBS 0.007663f
C511 B.n471 VSUBS 0.007663f
C512 B.n472 VSUBS 0.007663f
C513 B.n473 VSUBS 0.007663f
C514 B.n474 VSUBS 0.007663f
C515 B.n475 VSUBS 0.007663f
C516 B.n476 VSUBS 0.007663f
C517 B.n477 VSUBS 0.007663f
C518 B.n478 VSUBS 0.007663f
C519 B.n479 VSUBS 0.007663f
C520 B.n480 VSUBS 0.007663f
C521 B.n481 VSUBS 0.007663f
C522 B.n482 VSUBS 0.007663f
C523 B.n483 VSUBS 0.007663f
C524 B.n484 VSUBS 0.007663f
C525 B.n485 VSUBS 0.007663f
C526 B.n486 VSUBS 0.007663f
C527 B.n487 VSUBS 0.007663f
C528 B.n488 VSUBS 0.007663f
C529 B.n489 VSUBS 0.007663f
C530 B.n490 VSUBS 0.007663f
C531 B.n491 VSUBS 0.005297f
C532 B.n492 VSUBS 0.017756f
C533 B.n493 VSUBS 0.006198f
C534 B.n494 VSUBS 0.007663f
C535 B.n495 VSUBS 0.007663f
C536 B.n496 VSUBS 0.007663f
C537 B.n497 VSUBS 0.007663f
C538 B.n498 VSUBS 0.007663f
C539 B.n499 VSUBS 0.007663f
C540 B.n500 VSUBS 0.007663f
C541 B.n501 VSUBS 0.007663f
C542 B.n502 VSUBS 0.007663f
C543 B.n503 VSUBS 0.007663f
C544 B.n504 VSUBS 0.007663f
C545 B.n505 VSUBS 0.006198f
C546 B.n506 VSUBS 0.017756f
C547 B.n507 VSUBS 0.005297f
C548 B.n508 VSUBS 0.007663f
C549 B.n509 VSUBS 0.007663f
C550 B.n510 VSUBS 0.007663f
C551 B.n511 VSUBS 0.007663f
C552 B.n512 VSUBS 0.007663f
C553 B.n513 VSUBS 0.007663f
C554 B.n514 VSUBS 0.007663f
C555 B.n515 VSUBS 0.007663f
C556 B.n516 VSUBS 0.007663f
C557 B.n517 VSUBS 0.007663f
C558 B.n518 VSUBS 0.007663f
C559 B.n519 VSUBS 0.007663f
C560 B.n520 VSUBS 0.007663f
C561 B.n521 VSUBS 0.007663f
C562 B.n522 VSUBS 0.007663f
C563 B.n523 VSUBS 0.007663f
C564 B.n524 VSUBS 0.007663f
C565 B.n525 VSUBS 0.007663f
C566 B.n526 VSUBS 0.007663f
C567 B.n527 VSUBS 0.007663f
C568 B.n528 VSUBS 0.007663f
C569 B.n529 VSUBS 0.007663f
C570 B.n530 VSUBS 0.007663f
C571 B.n531 VSUBS 0.007663f
C572 B.n532 VSUBS 0.007663f
C573 B.n533 VSUBS 0.007663f
C574 B.n534 VSUBS 0.007663f
C575 B.n535 VSUBS 0.007663f
C576 B.n536 VSUBS 0.007663f
C577 B.n537 VSUBS 0.007663f
C578 B.n538 VSUBS 0.007663f
C579 B.n539 VSUBS 0.007663f
C580 B.n540 VSUBS 0.007663f
C581 B.n541 VSUBS 0.007663f
C582 B.n542 VSUBS 0.007663f
C583 B.n543 VSUBS 0.007663f
C584 B.n544 VSUBS 0.007663f
C585 B.n545 VSUBS 0.018815f
C586 B.n546 VSUBS 0.018376f
C587 B.n547 VSUBS 0.018376f
C588 B.n548 VSUBS 0.007663f
C589 B.n549 VSUBS 0.007663f
C590 B.n550 VSUBS 0.007663f
C591 B.n551 VSUBS 0.007663f
C592 B.n552 VSUBS 0.007663f
C593 B.n553 VSUBS 0.007663f
C594 B.n554 VSUBS 0.007663f
C595 B.n555 VSUBS 0.007663f
C596 B.n556 VSUBS 0.007663f
C597 B.n557 VSUBS 0.007663f
C598 B.n558 VSUBS 0.007663f
C599 B.n559 VSUBS 0.007663f
C600 B.n560 VSUBS 0.007663f
C601 B.n561 VSUBS 0.007663f
C602 B.n562 VSUBS 0.007663f
C603 B.n563 VSUBS 0.007663f
C604 B.n564 VSUBS 0.007663f
C605 B.n565 VSUBS 0.007663f
C606 B.n566 VSUBS 0.007663f
C607 B.n567 VSUBS 0.007663f
C608 B.n568 VSUBS 0.007663f
C609 B.n569 VSUBS 0.007663f
C610 B.n570 VSUBS 0.007663f
C611 B.n571 VSUBS 0.007663f
C612 B.n572 VSUBS 0.007663f
C613 B.n573 VSUBS 0.007663f
C614 B.n574 VSUBS 0.007663f
C615 B.n575 VSUBS 0.007663f
C616 B.n576 VSUBS 0.007663f
C617 B.n577 VSUBS 0.007663f
C618 B.n578 VSUBS 0.007663f
C619 B.n579 VSUBS 0.007663f
C620 B.n580 VSUBS 0.007663f
C621 B.n581 VSUBS 0.007663f
C622 B.n582 VSUBS 0.007663f
C623 B.n583 VSUBS 0.007663f
C624 B.n584 VSUBS 0.007663f
C625 B.n585 VSUBS 0.007663f
C626 B.n586 VSUBS 0.007663f
C627 B.n587 VSUBS 0.007663f
C628 B.n588 VSUBS 0.007663f
C629 B.n589 VSUBS 0.007663f
C630 B.n590 VSUBS 0.007663f
C631 B.n591 VSUBS 0.007663f
C632 B.n592 VSUBS 0.007663f
C633 B.n593 VSUBS 0.007663f
C634 B.n594 VSUBS 0.007663f
C635 B.n595 VSUBS 0.007663f
C636 B.n596 VSUBS 0.007663f
C637 B.n597 VSUBS 0.007663f
C638 B.n598 VSUBS 0.007663f
C639 B.n599 VSUBS 0.007663f
C640 B.n600 VSUBS 0.007663f
C641 B.n601 VSUBS 0.007663f
C642 B.n602 VSUBS 0.007663f
C643 B.n603 VSUBS 0.007663f
C644 B.n604 VSUBS 0.007663f
C645 B.n605 VSUBS 0.007663f
C646 B.n606 VSUBS 0.007663f
C647 B.n607 VSUBS 0.007663f
C648 B.n608 VSUBS 0.007663f
C649 B.n609 VSUBS 0.007663f
C650 B.n610 VSUBS 0.007663f
C651 B.n611 VSUBS 0.01f
C652 B.n612 VSUBS 0.010653f
C653 B.n613 VSUBS 0.021184f
C654 VDD1.n0 VSUBS 0.028913f
C655 VDD1.n1 VSUBS 0.026517f
C656 VDD1.n2 VSUBS 0.014249f
C657 VDD1.n3 VSUBS 0.033679f
C658 VDD1.n4 VSUBS 0.015087f
C659 VDD1.n5 VSUBS 0.026517f
C660 VDD1.n6 VSUBS 0.014249f
C661 VDD1.n7 VSUBS 0.033679f
C662 VDD1.n8 VSUBS 0.015087f
C663 VDD1.n9 VSUBS 0.689518f
C664 VDD1.n10 VSUBS 0.014249f
C665 VDD1.t3 VSUBS 0.071996f
C666 VDD1.n11 VSUBS 0.122196f
C667 VDD1.n12 VSUBS 0.021421f
C668 VDD1.n13 VSUBS 0.025259f
C669 VDD1.n14 VSUBS 0.033679f
C670 VDD1.n15 VSUBS 0.015087f
C671 VDD1.n16 VSUBS 0.014249f
C672 VDD1.n17 VSUBS 0.026517f
C673 VDD1.n18 VSUBS 0.026517f
C674 VDD1.n19 VSUBS 0.014249f
C675 VDD1.n20 VSUBS 0.015087f
C676 VDD1.n21 VSUBS 0.033679f
C677 VDD1.n22 VSUBS 0.033679f
C678 VDD1.n23 VSUBS 0.015087f
C679 VDD1.n24 VSUBS 0.014249f
C680 VDD1.n25 VSUBS 0.026517f
C681 VDD1.n26 VSUBS 0.026517f
C682 VDD1.n27 VSUBS 0.014249f
C683 VDD1.n28 VSUBS 0.015087f
C684 VDD1.n29 VSUBS 0.033679f
C685 VDD1.n30 VSUBS 0.080773f
C686 VDD1.n31 VSUBS 0.015087f
C687 VDD1.n32 VSUBS 0.014249f
C688 VDD1.n33 VSUBS 0.05948f
C689 VDD1.n34 VSUBS 0.066067f
C690 VDD1.t5 VSUBS 0.139764f
C691 VDD1.t4 VSUBS 0.139764f
C692 VDD1.n35 VSUBS 0.950881f
C693 VDD1.n36 VSUBS 0.835651f
C694 VDD1.n37 VSUBS 0.028913f
C695 VDD1.n38 VSUBS 0.026517f
C696 VDD1.n39 VSUBS 0.014249f
C697 VDD1.n40 VSUBS 0.033679f
C698 VDD1.n41 VSUBS 0.015087f
C699 VDD1.n42 VSUBS 0.026517f
C700 VDD1.n43 VSUBS 0.014249f
C701 VDD1.n44 VSUBS 0.033679f
C702 VDD1.n45 VSUBS 0.015087f
C703 VDD1.n46 VSUBS 0.689518f
C704 VDD1.n47 VSUBS 0.014249f
C705 VDD1.t8 VSUBS 0.071996f
C706 VDD1.n48 VSUBS 0.122196f
C707 VDD1.n49 VSUBS 0.021421f
C708 VDD1.n50 VSUBS 0.025259f
C709 VDD1.n51 VSUBS 0.033679f
C710 VDD1.n52 VSUBS 0.015087f
C711 VDD1.n53 VSUBS 0.014249f
C712 VDD1.n54 VSUBS 0.026517f
C713 VDD1.n55 VSUBS 0.026517f
C714 VDD1.n56 VSUBS 0.014249f
C715 VDD1.n57 VSUBS 0.015087f
C716 VDD1.n58 VSUBS 0.033679f
C717 VDD1.n59 VSUBS 0.033679f
C718 VDD1.n60 VSUBS 0.015087f
C719 VDD1.n61 VSUBS 0.014249f
C720 VDD1.n62 VSUBS 0.026517f
C721 VDD1.n63 VSUBS 0.026517f
C722 VDD1.n64 VSUBS 0.014249f
C723 VDD1.n65 VSUBS 0.015087f
C724 VDD1.n66 VSUBS 0.033679f
C725 VDD1.n67 VSUBS 0.080773f
C726 VDD1.n68 VSUBS 0.015087f
C727 VDD1.n69 VSUBS 0.014249f
C728 VDD1.n70 VSUBS 0.05948f
C729 VDD1.n71 VSUBS 0.066067f
C730 VDD1.t1 VSUBS 0.139764f
C731 VDD1.t9 VSUBS 0.139764f
C732 VDD1.n72 VSUBS 0.950876f
C733 VDD1.n73 VSUBS 0.827536f
C734 VDD1.t7 VSUBS 0.139764f
C735 VDD1.t2 VSUBS 0.139764f
C736 VDD1.n74 VSUBS 0.961215f
C737 VDD1.n75 VSUBS 2.58848f
C738 VDD1.t6 VSUBS 0.139764f
C739 VDD1.t0 VSUBS 0.139764f
C740 VDD1.n76 VSUBS 0.950876f
C741 VDD1.n77 VSUBS 2.77184f
C742 VP.n0 VSUBS 0.041954f
C743 VP.t7 VSUBS 1.2889f
C744 VP.n1 VSUBS 0.038493f
C745 VP.n2 VSUBS 0.041954f
C746 VP.t2 VSUBS 1.2889f
C747 VP.n3 VSUBS 0.034403f
C748 VP.n4 VSUBS 0.041954f
C749 VP.t0 VSUBS 1.2889f
C750 VP.n5 VSUBS 0.034403f
C751 VP.n6 VSUBS 0.041954f
C752 VP.t8 VSUBS 1.2889f
C753 VP.n7 VSUBS 0.038493f
C754 VP.n8 VSUBS 0.041954f
C755 VP.t1 VSUBS 1.2889f
C756 VP.n9 VSUBS 0.041954f
C757 VP.t9 VSUBS 1.2889f
C758 VP.n10 VSUBS 0.038493f
C759 VP.n11 VSUBS 0.041954f
C760 VP.t3 VSUBS 1.2889f
C761 VP.n12 VSUBS 0.034403f
C762 VP.n13 VSUBS 0.041954f
C763 VP.t5 VSUBS 1.2889f
C764 VP.n14 VSUBS 0.034403f
C765 VP.n15 VSUBS 0.270266f
C766 VP.t4 VSUBS 1.2889f
C767 VP.t6 VSUBS 1.4572f
C768 VP.n16 VSUBS 0.591549f
C769 VP.n17 VSUBS 0.565545f
C770 VP.n18 VSUBS 0.04422f
C771 VP.n19 VSUBS 0.081894f
C772 VP.n20 VSUBS 0.041954f
C773 VP.n21 VSUBS 0.041954f
C774 VP.n22 VSUBS 0.041954f
C775 VP.n23 VSUBS 0.084384f
C776 VP.n24 VSUBS 0.530424f
C777 VP.n25 VSUBS 0.084384f
C778 VP.n26 VSUBS 0.041954f
C779 VP.n27 VSUBS 0.041954f
C780 VP.n28 VSUBS 0.041954f
C781 VP.n29 VSUBS 0.081894f
C782 VP.n30 VSUBS 0.04422f
C783 VP.n31 VSUBS 0.490836f
C784 VP.n32 VSUBS 0.079756f
C785 VP.n33 VSUBS 0.041954f
C786 VP.n34 VSUBS 0.041954f
C787 VP.n35 VSUBS 0.041954f
C788 VP.n36 VSUBS 0.077799f
C789 VP.n37 VSUBS 0.048853f
C790 VP.n38 VSUBS 0.585174f
C791 VP.n39 VSUBS 1.89823f
C792 VP.n40 VSUBS 1.9323f
C793 VP.n41 VSUBS 0.585174f
C794 VP.n42 VSUBS 0.048853f
C795 VP.n43 VSUBS 0.077799f
C796 VP.n44 VSUBS 0.041954f
C797 VP.n45 VSUBS 0.041954f
C798 VP.n46 VSUBS 0.041954f
C799 VP.n47 VSUBS 0.079756f
C800 VP.n48 VSUBS 0.490836f
C801 VP.n49 VSUBS 0.04422f
C802 VP.n50 VSUBS 0.081894f
C803 VP.n51 VSUBS 0.041954f
C804 VP.n52 VSUBS 0.041954f
C805 VP.n53 VSUBS 0.041954f
C806 VP.n54 VSUBS 0.084384f
C807 VP.n55 VSUBS 0.530424f
C808 VP.n56 VSUBS 0.084384f
C809 VP.n57 VSUBS 0.041954f
C810 VP.n58 VSUBS 0.041954f
C811 VP.n59 VSUBS 0.041954f
C812 VP.n60 VSUBS 0.081894f
C813 VP.n61 VSUBS 0.04422f
C814 VP.n62 VSUBS 0.490836f
C815 VP.n63 VSUBS 0.079756f
C816 VP.n64 VSUBS 0.041954f
C817 VP.n65 VSUBS 0.041954f
C818 VP.n66 VSUBS 0.041954f
C819 VP.n67 VSUBS 0.077799f
C820 VP.n68 VSUBS 0.048853f
C821 VP.n69 VSUBS 0.585174f
C822 VP.n70 VSUBS 0.043388f
C823 VDD2.n0 VSUBS 0.028722f
C824 VDD2.n1 VSUBS 0.026342f
C825 VDD2.n2 VSUBS 0.014155f
C826 VDD2.n3 VSUBS 0.033457f
C827 VDD2.n4 VSUBS 0.014988f
C828 VDD2.n5 VSUBS 0.026342f
C829 VDD2.n6 VSUBS 0.014155f
C830 VDD2.n7 VSUBS 0.033457f
C831 VDD2.n8 VSUBS 0.014988f
C832 VDD2.n9 VSUBS 0.684978f
C833 VDD2.n10 VSUBS 0.014155f
C834 VDD2.t1 VSUBS 0.071522f
C835 VDD2.n11 VSUBS 0.121392f
C836 VDD2.n12 VSUBS 0.02128f
C837 VDD2.n13 VSUBS 0.025093f
C838 VDD2.n14 VSUBS 0.033457f
C839 VDD2.n15 VSUBS 0.014988f
C840 VDD2.n16 VSUBS 0.014155f
C841 VDD2.n17 VSUBS 0.026342f
C842 VDD2.n18 VSUBS 0.026342f
C843 VDD2.n19 VSUBS 0.014155f
C844 VDD2.n20 VSUBS 0.014988f
C845 VDD2.n21 VSUBS 0.033457f
C846 VDD2.n22 VSUBS 0.033457f
C847 VDD2.n23 VSUBS 0.014988f
C848 VDD2.n24 VSUBS 0.014155f
C849 VDD2.n25 VSUBS 0.026342f
C850 VDD2.n26 VSUBS 0.026342f
C851 VDD2.n27 VSUBS 0.014155f
C852 VDD2.n28 VSUBS 0.014988f
C853 VDD2.n29 VSUBS 0.033457f
C854 VDD2.n30 VSUBS 0.080241f
C855 VDD2.n31 VSUBS 0.014988f
C856 VDD2.n32 VSUBS 0.014155f
C857 VDD2.n33 VSUBS 0.059089f
C858 VDD2.n34 VSUBS 0.065632f
C859 VDD2.t2 VSUBS 0.138844f
C860 VDD2.t3 VSUBS 0.138844f
C861 VDD2.n35 VSUBS 0.944616f
C862 VDD2.n36 VSUBS 0.822088f
C863 VDD2.t8 VSUBS 0.138844f
C864 VDD2.t0 VSUBS 0.138844f
C865 VDD2.n37 VSUBS 0.954887f
C866 VDD2.n38 VSUBS 2.46738f
C867 VDD2.n39 VSUBS 0.028722f
C868 VDD2.n40 VSUBS 0.026342f
C869 VDD2.n41 VSUBS 0.014155f
C870 VDD2.n42 VSUBS 0.033457f
C871 VDD2.n43 VSUBS 0.014988f
C872 VDD2.n44 VSUBS 0.026342f
C873 VDD2.n45 VSUBS 0.014155f
C874 VDD2.n46 VSUBS 0.033457f
C875 VDD2.n47 VSUBS 0.014988f
C876 VDD2.n48 VSUBS 0.684978f
C877 VDD2.n49 VSUBS 0.014155f
C878 VDD2.t9 VSUBS 0.071522f
C879 VDD2.n50 VSUBS 0.121392f
C880 VDD2.n51 VSUBS 0.02128f
C881 VDD2.n52 VSUBS 0.025093f
C882 VDD2.n53 VSUBS 0.033457f
C883 VDD2.n54 VSUBS 0.014988f
C884 VDD2.n55 VSUBS 0.014155f
C885 VDD2.n56 VSUBS 0.026342f
C886 VDD2.n57 VSUBS 0.026342f
C887 VDD2.n58 VSUBS 0.014155f
C888 VDD2.n59 VSUBS 0.014988f
C889 VDD2.n60 VSUBS 0.033457f
C890 VDD2.n61 VSUBS 0.033457f
C891 VDD2.n62 VSUBS 0.014988f
C892 VDD2.n63 VSUBS 0.014155f
C893 VDD2.n64 VSUBS 0.026342f
C894 VDD2.n65 VSUBS 0.026342f
C895 VDD2.n66 VSUBS 0.014155f
C896 VDD2.n67 VSUBS 0.014988f
C897 VDD2.n68 VSUBS 0.033457f
C898 VDD2.n69 VSUBS 0.080241f
C899 VDD2.n70 VSUBS 0.014988f
C900 VDD2.n71 VSUBS 0.014155f
C901 VDD2.n72 VSUBS 0.059089f
C902 VDD2.n73 VSUBS 0.058466f
C903 VDD2.n74 VSUBS 2.2478f
C904 VDD2.t6 VSUBS 0.138844f
C905 VDD2.t7 VSUBS 0.138844f
C906 VDD2.n75 VSUBS 0.944621f
C907 VDD2.n76 VSUBS 0.636887f
C908 VDD2.t5 VSUBS 0.138844f
C909 VDD2.t4 VSUBS 0.138844f
C910 VDD2.n77 VSUBS 0.954854f
C911 VTAIL.t16 VSUBS 0.164309f
C912 VTAIL.t10 VSUBS 0.164309f
C913 VTAIL.n0 VSUBS 0.99553f
C914 VTAIL.n1 VSUBS 0.880865f
C915 VTAIL.n2 VSUBS 0.03399f
C916 VTAIL.n3 VSUBS 0.031173f
C917 VTAIL.n4 VSUBS 0.016751f
C918 VTAIL.n5 VSUBS 0.039594f
C919 VTAIL.n6 VSUBS 0.017737f
C920 VTAIL.n7 VSUBS 0.031173f
C921 VTAIL.n8 VSUBS 0.016751f
C922 VTAIL.n9 VSUBS 0.039594f
C923 VTAIL.n10 VSUBS 0.017737f
C924 VTAIL.n11 VSUBS 0.81061f
C925 VTAIL.n12 VSUBS 0.016751f
C926 VTAIL.t6 VSUBS 0.08464f
C927 VTAIL.n13 VSUBS 0.143656f
C928 VTAIL.n14 VSUBS 0.025183f
C929 VTAIL.n15 VSUBS 0.029695f
C930 VTAIL.n16 VSUBS 0.039594f
C931 VTAIL.n17 VSUBS 0.017737f
C932 VTAIL.n18 VSUBS 0.016751f
C933 VTAIL.n19 VSUBS 0.031173f
C934 VTAIL.n20 VSUBS 0.031173f
C935 VTAIL.n21 VSUBS 0.016751f
C936 VTAIL.n22 VSUBS 0.017737f
C937 VTAIL.n23 VSUBS 0.039594f
C938 VTAIL.n24 VSUBS 0.039594f
C939 VTAIL.n25 VSUBS 0.017737f
C940 VTAIL.n26 VSUBS 0.016751f
C941 VTAIL.n27 VSUBS 0.031173f
C942 VTAIL.n28 VSUBS 0.031173f
C943 VTAIL.n29 VSUBS 0.016751f
C944 VTAIL.n30 VSUBS 0.017737f
C945 VTAIL.n31 VSUBS 0.039594f
C946 VTAIL.n32 VSUBS 0.094958f
C947 VTAIL.n33 VSUBS 0.017737f
C948 VTAIL.n34 VSUBS 0.016751f
C949 VTAIL.n35 VSUBS 0.069926f
C950 VTAIL.n36 VSUBS 0.047647f
C951 VTAIL.n37 VSUBS 0.340187f
C952 VTAIL.t2 VSUBS 0.164309f
C953 VTAIL.t1 VSUBS 0.164309f
C954 VTAIL.n38 VSUBS 0.99553f
C955 VTAIL.n39 VSUBS 0.961612f
C956 VTAIL.t0 VSUBS 0.164309f
C957 VTAIL.t5 VSUBS 0.164309f
C958 VTAIL.n40 VSUBS 0.99553f
C959 VTAIL.n41 VSUBS 2.14102f
C960 VTAIL.t18 VSUBS 0.164309f
C961 VTAIL.t14 VSUBS 0.164309f
C962 VTAIL.n42 VSUBS 0.995537f
C963 VTAIL.n43 VSUBS 2.14101f
C964 VTAIL.t19 VSUBS 0.164309f
C965 VTAIL.t15 VSUBS 0.164309f
C966 VTAIL.n44 VSUBS 0.995537f
C967 VTAIL.n45 VSUBS 0.961605f
C968 VTAIL.n46 VSUBS 0.03399f
C969 VTAIL.n47 VSUBS 0.031173f
C970 VTAIL.n48 VSUBS 0.016751f
C971 VTAIL.n49 VSUBS 0.039594f
C972 VTAIL.n50 VSUBS 0.017737f
C973 VTAIL.n51 VSUBS 0.031173f
C974 VTAIL.n52 VSUBS 0.016751f
C975 VTAIL.n53 VSUBS 0.039594f
C976 VTAIL.n54 VSUBS 0.017737f
C977 VTAIL.n55 VSUBS 0.81061f
C978 VTAIL.n56 VSUBS 0.016751f
C979 VTAIL.t11 VSUBS 0.08464f
C980 VTAIL.n57 VSUBS 0.143656f
C981 VTAIL.n58 VSUBS 0.025183f
C982 VTAIL.n59 VSUBS 0.029695f
C983 VTAIL.n60 VSUBS 0.039594f
C984 VTAIL.n61 VSUBS 0.017737f
C985 VTAIL.n62 VSUBS 0.016751f
C986 VTAIL.n63 VSUBS 0.031173f
C987 VTAIL.n64 VSUBS 0.031173f
C988 VTAIL.n65 VSUBS 0.016751f
C989 VTAIL.n66 VSUBS 0.017737f
C990 VTAIL.n67 VSUBS 0.039594f
C991 VTAIL.n68 VSUBS 0.039594f
C992 VTAIL.n69 VSUBS 0.017737f
C993 VTAIL.n70 VSUBS 0.016751f
C994 VTAIL.n71 VSUBS 0.031173f
C995 VTAIL.n72 VSUBS 0.031173f
C996 VTAIL.n73 VSUBS 0.016751f
C997 VTAIL.n74 VSUBS 0.017737f
C998 VTAIL.n75 VSUBS 0.039594f
C999 VTAIL.n76 VSUBS 0.094958f
C1000 VTAIL.n77 VSUBS 0.017737f
C1001 VTAIL.n78 VSUBS 0.016751f
C1002 VTAIL.n79 VSUBS 0.069926f
C1003 VTAIL.n80 VSUBS 0.047647f
C1004 VTAIL.n81 VSUBS 0.340187f
C1005 VTAIL.t8 VSUBS 0.164309f
C1006 VTAIL.t4 VSUBS 0.164309f
C1007 VTAIL.n82 VSUBS 0.995537f
C1008 VTAIL.n83 VSUBS 0.919608f
C1009 VTAIL.t3 VSUBS 0.164309f
C1010 VTAIL.t7 VSUBS 0.164309f
C1011 VTAIL.n84 VSUBS 0.995537f
C1012 VTAIL.n85 VSUBS 0.961605f
C1013 VTAIL.n86 VSUBS 0.03399f
C1014 VTAIL.n87 VSUBS 0.031173f
C1015 VTAIL.n88 VSUBS 0.016751f
C1016 VTAIL.n89 VSUBS 0.039594f
C1017 VTAIL.n90 VSUBS 0.017737f
C1018 VTAIL.n91 VSUBS 0.031173f
C1019 VTAIL.n92 VSUBS 0.016751f
C1020 VTAIL.n93 VSUBS 0.039594f
C1021 VTAIL.n94 VSUBS 0.017737f
C1022 VTAIL.n95 VSUBS 0.81061f
C1023 VTAIL.n96 VSUBS 0.016751f
C1024 VTAIL.t9 VSUBS 0.08464f
C1025 VTAIL.n97 VSUBS 0.143656f
C1026 VTAIL.n98 VSUBS 0.025183f
C1027 VTAIL.n99 VSUBS 0.029695f
C1028 VTAIL.n100 VSUBS 0.039594f
C1029 VTAIL.n101 VSUBS 0.017737f
C1030 VTAIL.n102 VSUBS 0.016751f
C1031 VTAIL.n103 VSUBS 0.031173f
C1032 VTAIL.n104 VSUBS 0.031173f
C1033 VTAIL.n105 VSUBS 0.016751f
C1034 VTAIL.n106 VSUBS 0.017737f
C1035 VTAIL.n107 VSUBS 0.039594f
C1036 VTAIL.n108 VSUBS 0.039594f
C1037 VTAIL.n109 VSUBS 0.017737f
C1038 VTAIL.n110 VSUBS 0.016751f
C1039 VTAIL.n111 VSUBS 0.031173f
C1040 VTAIL.n112 VSUBS 0.031173f
C1041 VTAIL.n113 VSUBS 0.016751f
C1042 VTAIL.n114 VSUBS 0.017737f
C1043 VTAIL.n115 VSUBS 0.039594f
C1044 VTAIL.n116 VSUBS 0.094958f
C1045 VTAIL.n117 VSUBS 0.017737f
C1046 VTAIL.n118 VSUBS 0.016751f
C1047 VTAIL.n119 VSUBS 0.069926f
C1048 VTAIL.n120 VSUBS 0.047647f
C1049 VTAIL.n121 VSUBS 1.38321f
C1050 VTAIL.n122 VSUBS 0.03399f
C1051 VTAIL.n123 VSUBS 0.031173f
C1052 VTAIL.n124 VSUBS 0.016751f
C1053 VTAIL.n125 VSUBS 0.039594f
C1054 VTAIL.n126 VSUBS 0.017737f
C1055 VTAIL.n127 VSUBS 0.031173f
C1056 VTAIL.n128 VSUBS 0.016751f
C1057 VTAIL.n129 VSUBS 0.039594f
C1058 VTAIL.n130 VSUBS 0.017737f
C1059 VTAIL.n131 VSUBS 0.81061f
C1060 VTAIL.n132 VSUBS 0.016751f
C1061 VTAIL.t13 VSUBS 0.08464f
C1062 VTAIL.n133 VSUBS 0.143656f
C1063 VTAIL.n134 VSUBS 0.025183f
C1064 VTAIL.n135 VSUBS 0.029695f
C1065 VTAIL.n136 VSUBS 0.039594f
C1066 VTAIL.n137 VSUBS 0.017737f
C1067 VTAIL.n138 VSUBS 0.016751f
C1068 VTAIL.n139 VSUBS 0.031173f
C1069 VTAIL.n140 VSUBS 0.031173f
C1070 VTAIL.n141 VSUBS 0.016751f
C1071 VTAIL.n142 VSUBS 0.017737f
C1072 VTAIL.n143 VSUBS 0.039594f
C1073 VTAIL.n144 VSUBS 0.039594f
C1074 VTAIL.n145 VSUBS 0.017737f
C1075 VTAIL.n146 VSUBS 0.016751f
C1076 VTAIL.n147 VSUBS 0.031173f
C1077 VTAIL.n148 VSUBS 0.031173f
C1078 VTAIL.n149 VSUBS 0.016751f
C1079 VTAIL.n150 VSUBS 0.017737f
C1080 VTAIL.n151 VSUBS 0.039594f
C1081 VTAIL.n152 VSUBS 0.094958f
C1082 VTAIL.n153 VSUBS 0.017737f
C1083 VTAIL.n154 VSUBS 0.016751f
C1084 VTAIL.n155 VSUBS 0.069926f
C1085 VTAIL.n156 VSUBS 0.047647f
C1086 VTAIL.n157 VSUBS 1.38321f
C1087 VTAIL.t12 VSUBS 0.164309f
C1088 VTAIL.t17 VSUBS 0.164309f
C1089 VTAIL.n158 VSUBS 0.99553f
C1090 VTAIL.n159 VSUBS 0.821982f
C1091 VN.n0 VSUBS 0.040713f
C1092 VN.t9 VSUBS 1.25077f
C1093 VN.n1 VSUBS 0.037355f
C1094 VN.n2 VSUBS 0.040713f
C1095 VN.t1 VSUBS 1.25077f
C1096 VN.n3 VSUBS 0.033386f
C1097 VN.n4 VSUBS 0.040713f
C1098 VN.t6 VSUBS 1.25077f
C1099 VN.n5 VSUBS 0.033386f
C1100 VN.n6 VSUBS 0.262272f
C1101 VN.t7 VSUBS 1.25077f
C1102 VN.t8 VSUBS 1.4141f
C1103 VN.n7 VSUBS 0.574051f
C1104 VN.n8 VSUBS 0.548816f
C1105 VN.n9 VSUBS 0.042912f
C1106 VN.n10 VSUBS 0.079471f
C1107 VN.n11 VSUBS 0.040713f
C1108 VN.n12 VSUBS 0.040713f
C1109 VN.n13 VSUBS 0.040713f
C1110 VN.n14 VSUBS 0.081888f
C1111 VN.n15 VSUBS 0.514734f
C1112 VN.n16 VSUBS 0.081888f
C1113 VN.n17 VSUBS 0.040713f
C1114 VN.n18 VSUBS 0.040713f
C1115 VN.n19 VSUBS 0.040713f
C1116 VN.n20 VSUBS 0.079471f
C1117 VN.n21 VSUBS 0.042912f
C1118 VN.n22 VSUBS 0.476318f
C1119 VN.n23 VSUBS 0.077397f
C1120 VN.n24 VSUBS 0.040713f
C1121 VN.n25 VSUBS 0.040713f
C1122 VN.n26 VSUBS 0.040713f
C1123 VN.n27 VSUBS 0.075498f
C1124 VN.n28 VSUBS 0.047408f
C1125 VN.n29 VSUBS 0.567865f
C1126 VN.n30 VSUBS 0.042105f
C1127 VN.n31 VSUBS 0.040713f
C1128 VN.t0 VSUBS 1.25077f
C1129 VN.n32 VSUBS 0.037355f
C1130 VN.n33 VSUBS 0.040713f
C1131 VN.t3 VSUBS 1.25077f
C1132 VN.n34 VSUBS 0.033386f
C1133 VN.n35 VSUBS 0.040713f
C1134 VN.t2 VSUBS 1.25077f
C1135 VN.n36 VSUBS 0.033386f
C1136 VN.n37 VSUBS 0.262272f
C1137 VN.t4 VSUBS 1.25077f
C1138 VN.t5 VSUBS 1.4141f
C1139 VN.n38 VSUBS 0.574051f
C1140 VN.n39 VSUBS 0.548816f
C1141 VN.n40 VSUBS 0.042912f
C1142 VN.n41 VSUBS 0.079471f
C1143 VN.n42 VSUBS 0.040713f
C1144 VN.n43 VSUBS 0.040713f
C1145 VN.n44 VSUBS 0.040713f
C1146 VN.n45 VSUBS 0.081888f
C1147 VN.n46 VSUBS 0.514734f
C1148 VN.n47 VSUBS 0.081888f
C1149 VN.n48 VSUBS 0.040713f
C1150 VN.n49 VSUBS 0.040713f
C1151 VN.n50 VSUBS 0.040713f
C1152 VN.n51 VSUBS 0.079471f
C1153 VN.n52 VSUBS 0.042912f
C1154 VN.n53 VSUBS 0.476318f
C1155 VN.n54 VSUBS 0.077397f
C1156 VN.n55 VSUBS 0.040713f
C1157 VN.n56 VSUBS 0.040713f
C1158 VN.n57 VSUBS 0.040713f
C1159 VN.n58 VSUBS 0.075498f
C1160 VN.n59 VSUBS 0.047408f
C1161 VN.n60 VSUBS 0.567865f
C1162 VN.n61 VSUBS 1.86872f
.ends

