* NGSPICE file created from diff_pair_sample_1173.ext - technology: sky130A

.subckt diff_pair_sample_1173 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=0 ps=0 w=11.59 l=3.26
X1 B.t8 B.t6 B.t7 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=0 ps=0 w=11.59 l=3.26
X2 VTAIL.t19 VN.t0 VDD2.t9 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X3 B.t5 B.t3 B.t4 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=0 ps=0 w=11.59 l=3.26
X4 VTAIL.t18 VN.t1 VDD2.t1 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X5 VDD2.t6 VN.t2 VTAIL.t17 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=1.91235 ps=11.92 w=11.59 l=3.26
X6 VDD2.t7 VN.t3 VTAIL.t16 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=4.5201 ps=23.96 w=11.59 l=3.26
X7 VTAIL.t15 VN.t4 VDD2.t4 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X8 VDD2.t3 VN.t5 VTAIL.t14 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=1.91235 ps=11.92 w=11.59 l=3.26
X9 VDD1.t9 VP.t0 VTAIL.t6 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=4.5201 ps=23.96 w=11.59 l=3.26
X10 VDD1.t8 VP.t1 VTAIL.t3 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X11 VDD1.t7 VP.t2 VTAIL.t9 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=4.5201 ps=23.96 w=11.59 l=3.26
X12 VTAIL.t13 VN.t6 VDD2.t2 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X13 VDD1.t6 VP.t3 VTAIL.t2 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=1.91235 ps=11.92 w=11.59 l=3.26
X14 VDD1.t5 VP.t4 VTAIL.t4 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=1.91235 ps=11.92 w=11.59 l=3.26
X15 VDD2.t8 VN.t7 VTAIL.t12 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=4.5201 ps=23.96 w=11.59 l=3.26
X16 VDD1.t4 VP.t5 VTAIL.t1 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X17 VDD2.t5 VN.t8 VTAIL.t11 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X18 VTAIL.t8 VP.t6 VDD1.t3 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X19 VDD2.t0 VN.t9 VTAIL.t10 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X20 VTAIL.t0 VP.t7 VDD1.t2 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X21 VTAIL.t5 VP.t8 VDD1.t1 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X22 VTAIL.t7 VP.t9 VDD1.t0 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=1.91235 pd=11.92 as=1.91235 ps=11.92 w=11.59 l=3.26
X23 B.t2 B.t0 B.t1 w_n5278_n3286# sky130_fd_pr__pfet_01v8 ad=4.5201 pd=23.96 as=0 ps=0 w=11.59 l=3.26
R0 B.n485 B.n484 585
R1 B.n483 B.n160 585
R2 B.n482 B.n481 585
R3 B.n480 B.n161 585
R4 B.n479 B.n478 585
R5 B.n477 B.n162 585
R6 B.n476 B.n475 585
R7 B.n474 B.n163 585
R8 B.n473 B.n472 585
R9 B.n471 B.n164 585
R10 B.n470 B.n469 585
R11 B.n468 B.n165 585
R12 B.n467 B.n466 585
R13 B.n465 B.n166 585
R14 B.n464 B.n463 585
R15 B.n462 B.n167 585
R16 B.n461 B.n460 585
R17 B.n459 B.n168 585
R18 B.n458 B.n457 585
R19 B.n456 B.n169 585
R20 B.n455 B.n454 585
R21 B.n453 B.n170 585
R22 B.n452 B.n451 585
R23 B.n450 B.n171 585
R24 B.n449 B.n448 585
R25 B.n447 B.n172 585
R26 B.n446 B.n445 585
R27 B.n444 B.n173 585
R28 B.n443 B.n442 585
R29 B.n441 B.n174 585
R30 B.n440 B.n439 585
R31 B.n438 B.n175 585
R32 B.n437 B.n436 585
R33 B.n435 B.n176 585
R34 B.n434 B.n433 585
R35 B.n432 B.n177 585
R36 B.n431 B.n430 585
R37 B.n429 B.n178 585
R38 B.n428 B.n427 585
R39 B.n426 B.n179 585
R40 B.n425 B.n424 585
R41 B.n420 B.n180 585
R42 B.n419 B.n418 585
R43 B.n417 B.n181 585
R44 B.n416 B.n415 585
R45 B.n414 B.n182 585
R46 B.n413 B.n412 585
R47 B.n411 B.n183 585
R48 B.n410 B.n409 585
R49 B.n408 B.n184 585
R50 B.n406 B.n405 585
R51 B.n404 B.n187 585
R52 B.n403 B.n402 585
R53 B.n401 B.n188 585
R54 B.n400 B.n399 585
R55 B.n398 B.n189 585
R56 B.n397 B.n396 585
R57 B.n395 B.n190 585
R58 B.n394 B.n393 585
R59 B.n392 B.n191 585
R60 B.n391 B.n390 585
R61 B.n389 B.n192 585
R62 B.n388 B.n387 585
R63 B.n386 B.n193 585
R64 B.n385 B.n384 585
R65 B.n383 B.n194 585
R66 B.n382 B.n381 585
R67 B.n380 B.n195 585
R68 B.n379 B.n378 585
R69 B.n377 B.n196 585
R70 B.n376 B.n375 585
R71 B.n374 B.n197 585
R72 B.n373 B.n372 585
R73 B.n371 B.n198 585
R74 B.n370 B.n369 585
R75 B.n368 B.n199 585
R76 B.n367 B.n366 585
R77 B.n365 B.n200 585
R78 B.n364 B.n363 585
R79 B.n362 B.n201 585
R80 B.n361 B.n360 585
R81 B.n359 B.n202 585
R82 B.n358 B.n357 585
R83 B.n356 B.n203 585
R84 B.n355 B.n354 585
R85 B.n353 B.n204 585
R86 B.n352 B.n351 585
R87 B.n350 B.n205 585
R88 B.n349 B.n348 585
R89 B.n347 B.n206 585
R90 B.n486 B.n159 585
R91 B.n488 B.n487 585
R92 B.n489 B.n158 585
R93 B.n491 B.n490 585
R94 B.n492 B.n157 585
R95 B.n494 B.n493 585
R96 B.n495 B.n156 585
R97 B.n497 B.n496 585
R98 B.n498 B.n155 585
R99 B.n500 B.n499 585
R100 B.n501 B.n154 585
R101 B.n503 B.n502 585
R102 B.n504 B.n153 585
R103 B.n506 B.n505 585
R104 B.n507 B.n152 585
R105 B.n509 B.n508 585
R106 B.n510 B.n151 585
R107 B.n512 B.n511 585
R108 B.n513 B.n150 585
R109 B.n515 B.n514 585
R110 B.n516 B.n149 585
R111 B.n518 B.n517 585
R112 B.n519 B.n148 585
R113 B.n521 B.n520 585
R114 B.n522 B.n147 585
R115 B.n524 B.n523 585
R116 B.n525 B.n146 585
R117 B.n527 B.n526 585
R118 B.n528 B.n145 585
R119 B.n530 B.n529 585
R120 B.n531 B.n144 585
R121 B.n533 B.n532 585
R122 B.n534 B.n143 585
R123 B.n536 B.n535 585
R124 B.n537 B.n142 585
R125 B.n539 B.n538 585
R126 B.n540 B.n141 585
R127 B.n542 B.n541 585
R128 B.n543 B.n140 585
R129 B.n545 B.n544 585
R130 B.n546 B.n139 585
R131 B.n548 B.n547 585
R132 B.n549 B.n138 585
R133 B.n551 B.n550 585
R134 B.n552 B.n137 585
R135 B.n554 B.n553 585
R136 B.n555 B.n136 585
R137 B.n557 B.n556 585
R138 B.n558 B.n135 585
R139 B.n560 B.n559 585
R140 B.n561 B.n134 585
R141 B.n563 B.n562 585
R142 B.n564 B.n133 585
R143 B.n566 B.n565 585
R144 B.n567 B.n132 585
R145 B.n569 B.n568 585
R146 B.n570 B.n131 585
R147 B.n572 B.n571 585
R148 B.n573 B.n130 585
R149 B.n575 B.n574 585
R150 B.n576 B.n129 585
R151 B.n578 B.n577 585
R152 B.n579 B.n128 585
R153 B.n581 B.n580 585
R154 B.n582 B.n127 585
R155 B.n584 B.n583 585
R156 B.n585 B.n126 585
R157 B.n587 B.n586 585
R158 B.n588 B.n125 585
R159 B.n590 B.n589 585
R160 B.n591 B.n124 585
R161 B.n593 B.n592 585
R162 B.n594 B.n123 585
R163 B.n596 B.n595 585
R164 B.n597 B.n122 585
R165 B.n599 B.n598 585
R166 B.n600 B.n121 585
R167 B.n602 B.n601 585
R168 B.n603 B.n120 585
R169 B.n605 B.n604 585
R170 B.n606 B.n119 585
R171 B.n608 B.n607 585
R172 B.n609 B.n118 585
R173 B.n611 B.n610 585
R174 B.n612 B.n117 585
R175 B.n614 B.n613 585
R176 B.n615 B.n116 585
R177 B.n617 B.n616 585
R178 B.n618 B.n115 585
R179 B.n620 B.n619 585
R180 B.n621 B.n114 585
R181 B.n623 B.n622 585
R182 B.n624 B.n113 585
R183 B.n626 B.n625 585
R184 B.n627 B.n112 585
R185 B.n629 B.n628 585
R186 B.n630 B.n111 585
R187 B.n632 B.n631 585
R188 B.n633 B.n110 585
R189 B.n635 B.n634 585
R190 B.n636 B.n109 585
R191 B.n638 B.n637 585
R192 B.n639 B.n108 585
R193 B.n641 B.n640 585
R194 B.n642 B.n107 585
R195 B.n644 B.n643 585
R196 B.n645 B.n106 585
R197 B.n647 B.n646 585
R198 B.n648 B.n105 585
R199 B.n650 B.n649 585
R200 B.n651 B.n104 585
R201 B.n653 B.n652 585
R202 B.n654 B.n103 585
R203 B.n656 B.n655 585
R204 B.n657 B.n102 585
R205 B.n659 B.n658 585
R206 B.n660 B.n101 585
R207 B.n662 B.n661 585
R208 B.n663 B.n100 585
R209 B.n665 B.n664 585
R210 B.n666 B.n99 585
R211 B.n668 B.n667 585
R212 B.n669 B.n98 585
R213 B.n671 B.n670 585
R214 B.n672 B.n97 585
R215 B.n674 B.n673 585
R216 B.n675 B.n96 585
R217 B.n677 B.n676 585
R218 B.n678 B.n95 585
R219 B.n680 B.n679 585
R220 B.n681 B.n94 585
R221 B.n683 B.n682 585
R222 B.n684 B.n93 585
R223 B.n686 B.n685 585
R224 B.n687 B.n92 585
R225 B.n689 B.n688 585
R226 B.n690 B.n91 585
R227 B.n692 B.n691 585
R228 B.n693 B.n90 585
R229 B.n695 B.n694 585
R230 B.n696 B.n89 585
R231 B.n698 B.n697 585
R232 B.n699 B.n88 585
R233 B.n701 B.n700 585
R234 B.n837 B.n836 585
R235 B.n835 B.n38 585
R236 B.n834 B.n833 585
R237 B.n832 B.n39 585
R238 B.n831 B.n830 585
R239 B.n829 B.n40 585
R240 B.n828 B.n827 585
R241 B.n826 B.n41 585
R242 B.n825 B.n824 585
R243 B.n823 B.n42 585
R244 B.n822 B.n821 585
R245 B.n820 B.n43 585
R246 B.n819 B.n818 585
R247 B.n817 B.n44 585
R248 B.n816 B.n815 585
R249 B.n814 B.n45 585
R250 B.n813 B.n812 585
R251 B.n811 B.n46 585
R252 B.n810 B.n809 585
R253 B.n808 B.n47 585
R254 B.n807 B.n806 585
R255 B.n805 B.n48 585
R256 B.n804 B.n803 585
R257 B.n802 B.n49 585
R258 B.n801 B.n800 585
R259 B.n799 B.n50 585
R260 B.n798 B.n797 585
R261 B.n796 B.n51 585
R262 B.n795 B.n794 585
R263 B.n793 B.n52 585
R264 B.n792 B.n791 585
R265 B.n790 B.n53 585
R266 B.n789 B.n788 585
R267 B.n787 B.n54 585
R268 B.n786 B.n785 585
R269 B.n784 B.n55 585
R270 B.n783 B.n782 585
R271 B.n781 B.n56 585
R272 B.n780 B.n779 585
R273 B.n778 B.n57 585
R274 B.n776 B.n775 585
R275 B.n774 B.n60 585
R276 B.n773 B.n772 585
R277 B.n771 B.n61 585
R278 B.n770 B.n769 585
R279 B.n768 B.n62 585
R280 B.n767 B.n766 585
R281 B.n765 B.n63 585
R282 B.n764 B.n763 585
R283 B.n762 B.n64 585
R284 B.n761 B.n760 585
R285 B.n759 B.n65 585
R286 B.n758 B.n757 585
R287 B.n756 B.n69 585
R288 B.n755 B.n754 585
R289 B.n753 B.n70 585
R290 B.n752 B.n751 585
R291 B.n750 B.n71 585
R292 B.n749 B.n748 585
R293 B.n747 B.n72 585
R294 B.n746 B.n745 585
R295 B.n744 B.n73 585
R296 B.n743 B.n742 585
R297 B.n741 B.n74 585
R298 B.n740 B.n739 585
R299 B.n738 B.n75 585
R300 B.n737 B.n736 585
R301 B.n735 B.n76 585
R302 B.n734 B.n733 585
R303 B.n732 B.n77 585
R304 B.n731 B.n730 585
R305 B.n729 B.n78 585
R306 B.n728 B.n727 585
R307 B.n726 B.n79 585
R308 B.n725 B.n724 585
R309 B.n723 B.n80 585
R310 B.n722 B.n721 585
R311 B.n720 B.n81 585
R312 B.n719 B.n718 585
R313 B.n717 B.n82 585
R314 B.n716 B.n715 585
R315 B.n714 B.n83 585
R316 B.n713 B.n712 585
R317 B.n711 B.n84 585
R318 B.n710 B.n709 585
R319 B.n708 B.n85 585
R320 B.n707 B.n706 585
R321 B.n705 B.n86 585
R322 B.n704 B.n703 585
R323 B.n702 B.n87 585
R324 B.n838 B.n37 585
R325 B.n840 B.n839 585
R326 B.n841 B.n36 585
R327 B.n843 B.n842 585
R328 B.n844 B.n35 585
R329 B.n846 B.n845 585
R330 B.n847 B.n34 585
R331 B.n849 B.n848 585
R332 B.n850 B.n33 585
R333 B.n852 B.n851 585
R334 B.n853 B.n32 585
R335 B.n855 B.n854 585
R336 B.n856 B.n31 585
R337 B.n858 B.n857 585
R338 B.n859 B.n30 585
R339 B.n861 B.n860 585
R340 B.n862 B.n29 585
R341 B.n864 B.n863 585
R342 B.n865 B.n28 585
R343 B.n867 B.n866 585
R344 B.n868 B.n27 585
R345 B.n870 B.n869 585
R346 B.n871 B.n26 585
R347 B.n873 B.n872 585
R348 B.n874 B.n25 585
R349 B.n876 B.n875 585
R350 B.n877 B.n24 585
R351 B.n879 B.n878 585
R352 B.n880 B.n23 585
R353 B.n882 B.n881 585
R354 B.n883 B.n22 585
R355 B.n885 B.n884 585
R356 B.n886 B.n21 585
R357 B.n888 B.n887 585
R358 B.n889 B.n20 585
R359 B.n891 B.n890 585
R360 B.n892 B.n19 585
R361 B.n894 B.n893 585
R362 B.n895 B.n18 585
R363 B.n897 B.n896 585
R364 B.n898 B.n17 585
R365 B.n900 B.n899 585
R366 B.n901 B.n16 585
R367 B.n903 B.n902 585
R368 B.n904 B.n15 585
R369 B.n906 B.n905 585
R370 B.n907 B.n14 585
R371 B.n909 B.n908 585
R372 B.n910 B.n13 585
R373 B.n912 B.n911 585
R374 B.n913 B.n12 585
R375 B.n915 B.n914 585
R376 B.n916 B.n11 585
R377 B.n918 B.n917 585
R378 B.n919 B.n10 585
R379 B.n921 B.n920 585
R380 B.n922 B.n9 585
R381 B.n924 B.n923 585
R382 B.n925 B.n8 585
R383 B.n927 B.n926 585
R384 B.n928 B.n7 585
R385 B.n930 B.n929 585
R386 B.n931 B.n6 585
R387 B.n933 B.n932 585
R388 B.n934 B.n5 585
R389 B.n936 B.n935 585
R390 B.n937 B.n4 585
R391 B.n939 B.n938 585
R392 B.n940 B.n3 585
R393 B.n942 B.n941 585
R394 B.n943 B.n0 585
R395 B.n2 B.n1 585
R396 B.n242 B.n241 585
R397 B.n244 B.n243 585
R398 B.n245 B.n240 585
R399 B.n247 B.n246 585
R400 B.n248 B.n239 585
R401 B.n250 B.n249 585
R402 B.n251 B.n238 585
R403 B.n253 B.n252 585
R404 B.n254 B.n237 585
R405 B.n256 B.n255 585
R406 B.n257 B.n236 585
R407 B.n259 B.n258 585
R408 B.n260 B.n235 585
R409 B.n262 B.n261 585
R410 B.n263 B.n234 585
R411 B.n265 B.n264 585
R412 B.n266 B.n233 585
R413 B.n268 B.n267 585
R414 B.n269 B.n232 585
R415 B.n271 B.n270 585
R416 B.n272 B.n231 585
R417 B.n274 B.n273 585
R418 B.n275 B.n230 585
R419 B.n277 B.n276 585
R420 B.n278 B.n229 585
R421 B.n280 B.n279 585
R422 B.n281 B.n228 585
R423 B.n283 B.n282 585
R424 B.n284 B.n227 585
R425 B.n286 B.n285 585
R426 B.n287 B.n226 585
R427 B.n289 B.n288 585
R428 B.n290 B.n225 585
R429 B.n292 B.n291 585
R430 B.n293 B.n224 585
R431 B.n295 B.n294 585
R432 B.n296 B.n223 585
R433 B.n298 B.n297 585
R434 B.n299 B.n222 585
R435 B.n301 B.n300 585
R436 B.n302 B.n221 585
R437 B.n304 B.n303 585
R438 B.n305 B.n220 585
R439 B.n307 B.n306 585
R440 B.n308 B.n219 585
R441 B.n310 B.n309 585
R442 B.n311 B.n218 585
R443 B.n313 B.n312 585
R444 B.n314 B.n217 585
R445 B.n316 B.n315 585
R446 B.n317 B.n216 585
R447 B.n319 B.n318 585
R448 B.n320 B.n215 585
R449 B.n322 B.n321 585
R450 B.n323 B.n214 585
R451 B.n325 B.n324 585
R452 B.n326 B.n213 585
R453 B.n328 B.n327 585
R454 B.n329 B.n212 585
R455 B.n331 B.n330 585
R456 B.n332 B.n211 585
R457 B.n334 B.n333 585
R458 B.n335 B.n210 585
R459 B.n337 B.n336 585
R460 B.n338 B.n209 585
R461 B.n340 B.n339 585
R462 B.n341 B.n208 585
R463 B.n343 B.n342 585
R464 B.n344 B.n207 585
R465 B.n346 B.n345 585
R466 B.n345 B.n206 526.135
R467 B.n486 B.n485 526.135
R468 B.n702 B.n701 526.135
R469 B.n836 B.n37 526.135
R470 B.n185 B.t9 294.546
R471 B.n421 B.t3 294.546
R472 B.n66 B.t0 294.546
R473 B.n58 B.t6 294.546
R474 B.n945 B.n944 256.663
R475 B.n944 B.n943 235.042
R476 B.n944 B.n2 235.042
R477 B.n421 B.t4 177.409
R478 B.n66 B.t2 177.409
R479 B.n185 B.t10 177.394
R480 B.n58 B.t8 177.394
R481 B.n349 B.n206 163.367
R482 B.n350 B.n349 163.367
R483 B.n351 B.n350 163.367
R484 B.n351 B.n204 163.367
R485 B.n355 B.n204 163.367
R486 B.n356 B.n355 163.367
R487 B.n357 B.n356 163.367
R488 B.n357 B.n202 163.367
R489 B.n361 B.n202 163.367
R490 B.n362 B.n361 163.367
R491 B.n363 B.n362 163.367
R492 B.n363 B.n200 163.367
R493 B.n367 B.n200 163.367
R494 B.n368 B.n367 163.367
R495 B.n369 B.n368 163.367
R496 B.n369 B.n198 163.367
R497 B.n373 B.n198 163.367
R498 B.n374 B.n373 163.367
R499 B.n375 B.n374 163.367
R500 B.n375 B.n196 163.367
R501 B.n379 B.n196 163.367
R502 B.n380 B.n379 163.367
R503 B.n381 B.n380 163.367
R504 B.n381 B.n194 163.367
R505 B.n385 B.n194 163.367
R506 B.n386 B.n385 163.367
R507 B.n387 B.n386 163.367
R508 B.n387 B.n192 163.367
R509 B.n391 B.n192 163.367
R510 B.n392 B.n391 163.367
R511 B.n393 B.n392 163.367
R512 B.n393 B.n190 163.367
R513 B.n397 B.n190 163.367
R514 B.n398 B.n397 163.367
R515 B.n399 B.n398 163.367
R516 B.n399 B.n188 163.367
R517 B.n403 B.n188 163.367
R518 B.n404 B.n403 163.367
R519 B.n405 B.n404 163.367
R520 B.n405 B.n184 163.367
R521 B.n410 B.n184 163.367
R522 B.n411 B.n410 163.367
R523 B.n412 B.n411 163.367
R524 B.n412 B.n182 163.367
R525 B.n416 B.n182 163.367
R526 B.n417 B.n416 163.367
R527 B.n418 B.n417 163.367
R528 B.n418 B.n180 163.367
R529 B.n425 B.n180 163.367
R530 B.n426 B.n425 163.367
R531 B.n427 B.n426 163.367
R532 B.n427 B.n178 163.367
R533 B.n431 B.n178 163.367
R534 B.n432 B.n431 163.367
R535 B.n433 B.n432 163.367
R536 B.n433 B.n176 163.367
R537 B.n437 B.n176 163.367
R538 B.n438 B.n437 163.367
R539 B.n439 B.n438 163.367
R540 B.n439 B.n174 163.367
R541 B.n443 B.n174 163.367
R542 B.n444 B.n443 163.367
R543 B.n445 B.n444 163.367
R544 B.n445 B.n172 163.367
R545 B.n449 B.n172 163.367
R546 B.n450 B.n449 163.367
R547 B.n451 B.n450 163.367
R548 B.n451 B.n170 163.367
R549 B.n455 B.n170 163.367
R550 B.n456 B.n455 163.367
R551 B.n457 B.n456 163.367
R552 B.n457 B.n168 163.367
R553 B.n461 B.n168 163.367
R554 B.n462 B.n461 163.367
R555 B.n463 B.n462 163.367
R556 B.n463 B.n166 163.367
R557 B.n467 B.n166 163.367
R558 B.n468 B.n467 163.367
R559 B.n469 B.n468 163.367
R560 B.n469 B.n164 163.367
R561 B.n473 B.n164 163.367
R562 B.n474 B.n473 163.367
R563 B.n475 B.n474 163.367
R564 B.n475 B.n162 163.367
R565 B.n479 B.n162 163.367
R566 B.n480 B.n479 163.367
R567 B.n481 B.n480 163.367
R568 B.n481 B.n160 163.367
R569 B.n485 B.n160 163.367
R570 B.n701 B.n88 163.367
R571 B.n697 B.n88 163.367
R572 B.n697 B.n696 163.367
R573 B.n696 B.n695 163.367
R574 B.n695 B.n90 163.367
R575 B.n691 B.n90 163.367
R576 B.n691 B.n690 163.367
R577 B.n690 B.n689 163.367
R578 B.n689 B.n92 163.367
R579 B.n685 B.n92 163.367
R580 B.n685 B.n684 163.367
R581 B.n684 B.n683 163.367
R582 B.n683 B.n94 163.367
R583 B.n679 B.n94 163.367
R584 B.n679 B.n678 163.367
R585 B.n678 B.n677 163.367
R586 B.n677 B.n96 163.367
R587 B.n673 B.n96 163.367
R588 B.n673 B.n672 163.367
R589 B.n672 B.n671 163.367
R590 B.n671 B.n98 163.367
R591 B.n667 B.n98 163.367
R592 B.n667 B.n666 163.367
R593 B.n666 B.n665 163.367
R594 B.n665 B.n100 163.367
R595 B.n661 B.n100 163.367
R596 B.n661 B.n660 163.367
R597 B.n660 B.n659 163.367
R598 B.n659 B.n102 163.367
R599 B.n655 B.n102 163.367
R600 B.n655 B.n654 163.367
R601 B.n654 B.n653 163.367
R602 B.n653 B.n104 163.367
R603 B.n649 B.n104 163.367
R604 B.n649 B.n648 163.367
R605 B.n648 B.n647 163.367
R606 B.n647 B.n106 163.367
R607 B.n643 B.n106 163.367
R608 B.n643 B.n642 163.367
R609 B.n642 B.n641 163.367
R610 B.n641 B.n108 163.367
R611 B.n637 B.n108 163.367
R612 B.n637 B.n636 163.367
R613 B.n636 B.n635 163.367
R614 B.n635 B.n110 163.367
R615 B.n631 B.n110 163.367
R616 B.n631 B.n630 163.367
R617 B.n630 B.n629 163.367
R618 B.n629 B.n112 163.367
R619 B.n625 B.n112 163.367
R620 B.n625 B.n624 163.367
R621 B.n624 B.n623 163.367
R622 B.n623 B.n114 163.367
R623 B.n619 B.n114 163.367
R624 B.n619 B.n618 163.367
R625 B.n618 B.n617 163.367
R626 B.n617 B.n116 163.367
R627 B.n613 B.n116 163.367
R628 B.n613 B.n612 163.367
R629 B.n612 B.n611 163.367
R630 B.n611 B.n118 163.367
R631 B.n607 B.n118 163.367
R632 B.n607 B.n606 163.367
R633 B.n606 B.n605 163.367
R634 B.n605 B.n120 163.367
R635 B.n601 B.n120 163.367
R636 B.n601 B.n600 163.367
R637 B.n600 B.n599 163.367
R638 B.n599 B.n122 163.367
R639 B.n595 B.n122 163.367
R640 B.n595 B.n594 163.367
R641 B.n594 B.n593 163.367
R642 B.n593 B.n124 163.367
R643 B.n589 B.n124 163.367
R644 B.n589 B.n588 163.367
R645 B.n588 B.n587 163.367
R646 B.n587 B.n126 163.367
R647 B.n583 B.n126 163.367
R648 B.n583 B.n582 163.367
R649 B.n582 B.n581 163.367
R650 B.n581 B.n128 163.367
R651 B.n577 B.n128 163.367
R652 B.n577 B.n576 163.367
R653 B.n576 B.n575 163.367
R654 B.n575 B.n130 163.367
R655 B.n571 B.n130 163.367
R656 B.n571 B.n570 163.367
R657 B.n570 B.n569 163.367
R658 B.n569 B.n132 163.367
R659 B.n565 B.n132 163.367
R660 B.n565 B.n564 163.367
R661 B.n564 B.n563 163.367
R662 B.n563 B.n134 163.367
R663 B.n559 B.n134 163.367
R664 B.n559 B.n558 163.367
R665 B.n558 B.n557 163.367
R666 B.n557 B.n136 163.367
R667 B.n553 B.n136 163.367
R668 B.n553 B.n552 163.367
R669 B.n552 B.n551 163.367
R670 B.n551 B.n138 163.367
R671 B.n547 B.n138 163.367
R672 B.n547 B.n546 163.367
R673 B.n546 B.n545 163.367
R674 B.n545 B.n140 163.367
R675 B.n541 B.n140 163.367
R676 B.n541 B.n540 163.367
R677 B.n540 B.n539 163.367
R678 B.n539 B.n142 163.367
R679 B.n535 B.n142 163.367
R680 B.n535 B.n534 163.367
R681 B.n534 B.n533 163.367
R682 B.n533 B.n144 163.367
R683 B.n529 B.n144 163.367
R684 B.n529 B.n528 163.367
R685 B.n528 B.n527 163.367
R686 B.n527 B.n146 163.367
R687 B.n523 B.n146 163.367
R688 B.n523 B.n522 163.367
R689 B.n522 B.n521 163.367
R690 B.n521 B.n148 163.367
R691 B.n517 B.n148 163.367
R692 B.n517 B.n516 163.367
R693 B.n516 B.n515 163.367
R694 B.n515 B.n150 163.367
R695 B.n511 B.n150 163.367
R696 B.n511 B.n510 163.367
R697 B.n510 B.n509 163.367
R698 B.n509 B.n152 163.367
R699 B.n505 B.n152 163.367
R700 B.n505 B.n504 163.367
R701 B.n504 B.n503 163.367
R702 B.n503 B.n154 163.367
R703 B.n499 B.n154 163.367
R704 B.n499 B.n498 163.367
R705 B.n498 B.n497 163.367
R706 B.n497 B.n156 163.367
R707 B.n493 B.n156 163.367
R708 B.n493 B.n492 163.367
R709 B.n492 B.n491 163.367
R710 B.n491 B.n158 163.367
R711 B.n487 B.n158 163.367
R712 B.n487 B.n486 163.367
R713 B.n836 B.n835 163.367
R714 B.n835 B.n834 163.367
R715 B.n834 B.n39 163.367
R716 B.n830 B.n39 163.367
R717 B.n830 B.n829 163.367
R718 B.n829 B.n828 163.367
R719 B.n828 B.n41 163.367
R720 B.n824 B.n41 163.367
R721 B.n824 B.n823 163.367
R722 B.n823 B.n822 163.367
R723 B.n822 B.n43 163.367
R724 B.n818 B.n43 163.367
R725 B.n818 B.n817 163.367
R726 B.n817 B.n816 163.367
R727 B.n816 B.n45 163.367
R728 B.n812 B.n45 163.367
R729 B.n812 B.n811 163.367
R730 B.n811 B.n810 163.367
R731 B.n810 B.n47 163.367
R732 B.n806 B.n47 163.367
R733 B.n806 B.n805 163.367
R734 B.n805 B.n804 163.367
R735 B.n804 B.n49 163.367
R736 B.n800 B.n49 163.367
R737 B.n800 B.n799 163.367
R738 B.n799 B.n798 163.367
R739 B.n798 B.n51 163.367
R740 B.n794 B.n51 163.367
R741 B.n794 B.n793 163.367
R742 B.n793 B.n792 163.367
R743 B.n792 B.n53 163.367
R744 B.n788 B.n53 163.367
R745 B.n788 B.n787 163.367
R746 B.n787 B.n786 163.367
R747 B.n786 B.n55 163.367
R748 B.n782 B.n55 163.367
R749 B.n782 B.n781 163.367
R750 B.n781 B.n780 163.367
R751 B.n780 B.n57 163.367
R752 B.n775 B.n57 163.367
R753 B.n775 B.n774 163.367
R754 B.n774 B.n773 163.367
R755 B.n773 B.n61 163.367
R756 B.n769 B.n61 163.367
R757 B.n769 B.n768 163.367
R758 B.n768 B.n767 163.367
R759 B.n767 B.n63 163.367
R760 B.n763 B.n63 163.367
R761 B.n763 B.n762 163.367
R762 B.n762 B.n761 163.367
R763 B.n761 B.n65 163.367
R764 B.n757 B.n65 163.367
R765 B.n757 B.n756 163.367
R766 B.n756 B.n755 163.367
R767 B.n755 B.n70 163.367
R768 B.n751 B.n70 163.367
R769 B.n751 B.n750 163.367
R770 B.n750 B.n749 163.367
R771 B.n749 B.n72 163.367
R772 B.n745 B.n72 163.367
R773 B.n745 B.n744 163.367
R774 B.n744 B.n743 163.367
R775 B.n743 B.n74 163.367
R776 B.n739 B.n74 163.367
R777 B.n739 B.n738 163.367
R778 B.n738 B.n737 163.367
R779 B.n737 B.n76 163.367
R780 B.n733 B.n76 163.367
R781 B.n733 B.n732 163.367
R782 B.n732 B.n731 163.367
R783 B.n731 B.n78 163.367
R784 B.n727 B.n78 163.367
R785 B.n727 B.n726 163.367
R786 B.n726 B.n725 163.367
R787 B.n725 B.n80 163.367
R788 B.n721 B.n80 163.367
R789 B.n721 B.n720 163.367
R790 B.n720 B.n719 163.367
R791 B.n719 B.n82 163.367
R792 B.n715 B.n82 163.367
R793 B.n715 B.n714 163.367
R794 B.n714 B.n713 163.367
R795 B.n713 B.n84 163.367
R796 B.n709 B.n84 163.367
R797 B.n709 B.n708 163.367
R798 B.n708 B.n707 163.367
R799 B.n707 B.n86 163.367
R800 B.n703 B.n86 163.367
R801 B.n703 B.n702 163.367
R802 B.n840 B.n37 163.367
R803 B.n841 B.n840 163.367
R804 B.n842 B.n841 163.367
R805 B.n842 B.n35 163.367
R806 B.n846 B.n35 163.367
R807 B.n847 B.n846 163.367
R808 B.n848 B.n847 163.367
R809 B.n848 B.n33 163.367
R810 B.n852 B.n33 163.367
R811 B.n853 B.n852 163.367
R812 B.n854 B.n853 163.367
R813 B.n854 B.n31 163.367
R814 B.n858 B.n31 163.367
R815 B.n859 B.n858 163.367
R816 B.n860 B.n859 163.367
R817 B.n860 B.n29 163.367
R818 B.n864 B.n29 163.367
R819 B.n865 B.n864 163.367
R820 B.n866 B.n865 163.367
R821 B.n866 B.n27 163.367
R822 B.n870 B.n27 163.367
R823 B.n871 B.n870 163.367
R824 B.n872 B.n871 163.367
R825 B.n872 B.n25 163.367
R826 B.n876 B.n25 163.367
R827 B.n877 B.n876 163.367
R828 B.n878 B.n877 163.367
R829 B.n878 B.n23 163.367
R830 B.n882 B.n23 163.367
R831 B.n883 B.n882 163.367
R832 B.n884 B.n883 163.367
R833 B.n884 B.n21 163.367
R834 B.n888 B.n21 163.367
R835 B.n889 B.n888 163.367
R836 B.n890 B.n889 163.367
R837 B.n890 B.n19 163.367
R838 B.n894 B.n19 163.367
R839 B.n895 B.n894 163.367
R840 B.n896 B.n895 163.367
R841 B.n896 B.n17 163.367
R842 B.n900 B.n17 163.367
R843 B.n901 B.n900 163.367
R844 B.n902 B.n901 163.367
R845 B.n902 B.n15 163.367
R846 B.n906 B.n15 163.367
R847 B.n907 B.n906 163.367
R848 B.n908 B.n907 163.367
R849 B.n908 B.n13 163.367
R850 B.n912 B.n13 163.367
R851 B.n913 B.n912 163.367
R852 B.n914 B.n913 163.367
R853 B.n914 B.n11 163.367
R854 B.n918 B.n11 163.367
R855 B.n919 B.n918 163.367
R856 B.n920 B.n919 163.367
R857 B.n920 B.n9 163.367
R858 B.n924 B.n9 163.367
R859 B.n925 B.n924 163.367
R860 B.n926 B.n925 163.367
R861 B.n926 B.n7 163.367
R862 B.n930 B.n7 163.367
R863 B.n931 B.n930 163.367
R864 B.n932 B.n931 163.367
R865 B.n932 B.n5 163.367
R866 B.n936 B.n5 163.367
R867 B.n937 B.n936 163.367
R868 B.n938 B.n937 163.367
R869 B.n938 B.n3 163.367
R870 B.n942 B.n3 163.367
R871 B.n943 B.n942 163.367
R872 B.n242 B.n2 163.367
R873 B.n243 B.n242 163.367
R874 B.n243 B.n240 163.367
R875 B.n247 B.n240 163.367
R876 B.n248 B.n247 163.367
R877 B.n249 B.n248 163.367
R878 B.n249 B.n238 163.367
R879 B.n253 B.n238 163.367
R880 B.n254 B.n253 163.367
R881 B.n255 B.n254 163.367
R882 B.n255 B.n236 163.367
R883 B.n259 B.n236 163.367
R884 B.n260 B.n259 163.367
R885 B.n261 B.n260 163.367
R886 B.n261 B.n234 163.367
R887 B.n265 B.n234 163.367
R888 B.n266 B.n265 163.367
R889 B.n267 B.n266 163.367
R890 B.n267 B.n232 163.367
R891 B.n271 B.n232 163.367
R892 B.n272 B.n271 163.367
R893 B.n273 B.n272 163.367
R894 B.n273 B.n230 163.367
R895 B.n277 B.n230 163.367
R896 B.n278 B.n277 163.367
R897 B.n279 B.n278 163.367
R898 B.n279 B.n228 163.367
R899 B.n283 B.n228 163.367
R900 B.n284 B.n283 163.367
R901 B.n285 B.n284 163.367
R902 B.n285 B.n226 163.367
R903 B.n289 B.n226 163.367
R904 B.n290 B.n289 163.367
R905 B.n291 B.n290 163.367
R906 B.n291 B.n224 163.367
R907 B.n295 B.n224 163.367
R908 B.n296 B.n295 163.367
R909 B.n297 B.n296 163.367
R910 B.n297 B.n222 163.367
R911 B.n301 B.n222 163.367
R912 B.n302 B.n301 163.367
R913 B.n303 B.n302 163.367
R914 B.n303 B.n220 163.367
R915 B.n307 B.n220 163.367
R916 B.n308 B.n307 163.367
R917 B.n309 B.n308 163.367
R918 B.n309 B.n218 163.367
R919 B.n313 B.n218 163.367
R920 B.n314 B.n313 163.367
R921 B.n315 B.n314 163.367
R922 B.n315 B.n216 163.367
R923 B.n319 B.n216 163.367
R924 B.n320 B.n319 163.367
R925 B.n321 B.n320 163.367
R926 B.n321 B.n214 163.367
R927 B.n325 B.n214 163.367
R928 B.n326 B.n325 163.367
R929 B.n327 B.n326 163.367
R930 B.n327 B.n212 163.367
R931 B.n331 B.n212 163.367
R932 B.n332 B.n331 163.367
R933 B.n333 B.n332 163.367
R934 B.n333 B.n210 163.367
R935 B.n337 B.n210 163.367
R936 B.n338 B.n337 163.367
R937 B.n339 B.n338 163.367
R938 B.n339 B.n208 163.367
R939 B.n343 B.n208 163.367
R940 B.n344 B.n343 163.367
R941 B.n345 B.n344 163.367
R942 B.n422 B.t5 107.784
R943 B.n67 B.t1 107.784
R944 B.n186 B.t11 107.77
R945 B.n59 B.t7 107.77
R946 B.n186 B.n185 69.6247
R947 B.n422 B.n421 69.6247
R948 B.n67 B.n66 69.6247
R949 B.n59 B.n58 69.6247
R950 B.n407 B.n186 59.5399
R951 B.n423 B.n422 59.5399
R952 B.n68 B.n67 59.5399
R953 B.n777 B.n59 59.5399
R954 B.n838 B.n837 34.1859
R955 B.n700 B.n87 34.1859
R956 B.n484 B.n159 34.1859
R957 B.n347 B.n346 34.1859
R958 B B.n945 18.0485
R959 B.n839 B.n838 10.6151
R960 B.n839 B.n36 10.6151
R961 B.n843 B.n36 10.6151
R962 B.n844 B.n843 10.6151
R963 B.n845 B.n844 10.6151
R964 B.n845 B.n34 10.6151
R965 B.n849 B.n34 10.6151
R966 B.n850 B.n849 10.6151
R967 B.n851 B.n850 10.6151
R968 B.n851 B.n32 10.6151
R969 B.n855 B.n32 10.6151
R970 B.n856 B.n855 10.6151
R971 B.n857 B.n856 10.6151
R972 B.n857 B.n30 10.6151
R973 B.n861 B.n30 10.6151
R974 B.n862 B.n861 10.6151
R975 B.n863 B.n862 10.6151
R976 B.n863 B.n28 10.6151
R977 B.n867 B.n28 10.6151
R978 B.n868 B.n867 10.6151
R979 B.n869 B.n868 10.6151
R980 B.n869 B.n26 10.6151
R981 B.n873 B.n26 10.6151
R982 B.n874 B.n873 10.6151
R983 B.n875 B.n874 10.6151
R984 B.n875 B.n24 10.6151
R985 B.n879 B.n24 10.6151
R986 B.n880 B.n879 10.6151
R987 B.n881 B.n880 10.6151
R988 B.n881 B.n22 10.6151
R989 B.n885 B.n22 10.6151
R990 B.n886 B.n885 10.6151
R991 B.n887 B.n886 10.6151
R992 B.n887 B.n20 10.6151
R993 B.n891 B.n20 10.6151
R994 B.n892 B.n891 10.6151
R995 B.n893 B.n892 10.6151
R996 B.n893 B.n18 10.6151
R997 B.n897 B.n18 10.6151
R998 B.n898 B.n897 10.6151
R999 B.n899 B.n898 10.6151
R1000 B.n899 B.n16 10.6151
R1001 B.n903 B.n16 10.6151
R1002 B.n904 B.n903 10.6151
R1003 B.n905 B.n904 10.6151
R1004 B.n905 B.n14 10.6151
R1005 B.n909 B.n14 10.6151
R1006 B.n910 B.n909 10.6151
R1007 B.n911 B.n910 10.6151
R1008 B.n911 B.n12 10.6151
R1009 B.n915 B.n12 10.6151
R1010 B.n916 B.n915 10.6151
R1011 B.n917 B.n916 10.6151
R1012 B.n917 B.n10 10.6151
R1013 B.n921 B.n10 10.6151
R1014 B.n922 B.n921 10.6151
R1015 B.n923 B.n922 10.6151
R1016 B.n923 B.n8 10.6151
R1017 B.n927 B.n8 10.6151
R1018 B.n928 B.n927 10.6151
R1019 B.n929 B.n928 10.6151
R1020 B.n929 B.n6 10.6151
R1021 B.n933 B.n6 10.6151
R1022 B.n934 B.n933 10.6151
R1023 B.n935 B.n934 10.6151
R1024 B.n935 B.n4 10.6151
R1025 B.n939 B.n4 10.6151
R1026 B.n940 B.n939 10.6151
R1027 B.n941 B.n940 10.6151
R1028 B.n941 B.n0 10.6151
R1029 B.n837 B.n38 10.6151
R1030 B.n833 B.n38 10.6151
R1031 B.n833 B.n832 10.6151
R1032 B.n832 B.n831 10.6151
R1033 B.n831 B.n40 10.6151
R1034 B.n827 B.n40 10.6151
R1035 B.n827 B.n826 10.6151
R1036 B.n826 B.n825 10.6151
R1037 B.n825 B.n42 10.6151
R1038 B.n821 B.n42 10.6151
R1039 B.n821 B.n820 10.6151
R1040 B.n820 B.n819 10.6151
R1041 B.n819 B.n44 10.6151
R1042 B.n815 B.n44 10.6151
R1043 B.n815 B.n814 10.6151
R1044 B.n814 B.n813 10.6151
R1045 B.n813 B.n46 10.6151
R1046 B.n809 B.n46 10.6151
R1047 B.n809 B.n808 10.6151
R1048 B.n808 B.n807 10.6151
R1049 B.n807 B.n48 10.6151
R1050 B.n803 B.n48 10.6151
R1051 B.n803 B.n802 10.6151
R1052 B.n802 B.n801 10.6151
R1053 B.n801 B.n50 10.6151
R1054 B.n797 B.n50 10.6151
R1055 B.n797 B.n796 10.6151
R1056 B.n796 B.n795 10.6151
R1057 B.n795 B.n52 10.6151
R1058 B.n791 B.n52 10.6151
R1059 B.n791 B.n790 10.6151
R1060 B.n790 B.n789 10.6151
R1061 B.n789 B.n54 10.6151
R1062 B.n785 B.n54 10.6151
R1063 B.n785 B.n784 10.6151
R1064 B.n784 B.n783 10.6151
R1065 B.n783 B.n56 10.6151
R1066 B.n779 B.n56 10.6151
R1067 B.n779 B.n778 10.6151
R1068 B.n776 B.n60 10.6151
R1069 B.n772 B.n60 10.6151
R1070 B.n772 B.n771 10.6151
R1071 B.n771 B.n770 10.6151
R1072 B.n770 B.n62 10.6151
R1073 B.n766 B.n62 10.6151
R1074 B.n766 B.n765 10.6151
R1075 B.n765 B.n764 10.6151
R1076 B.n764 B.n64 10.6151
R1077 B.n760 B.n759 10.6151
R1078 B.n759 B.n758 10.6151
R1079 B.n758 B.n69 10.6151
R1080 B.n754 B.n69 10.6151
R1081 B.n754 B.n753 10.6151
R1082 B.n753 B.n752 10.6151
R1083 B.n752 B.n71 10.6151
R1084 B.n748 B.n71 10.6151
R1085 B.n748 B.n747 10.6151
R1086 B.n747 B.n746 10.6151
R1087 B.n746 B.n73 10.6151
R1088 B.n742 B.n73 10.6151
R1089 B.n742 B.n741 10.6151
R1090 B.n741 B.n740 10.6151
R1091 B.n740 B.n75 10.6151
R1092 B.n736 B.n75 10.6151
R1093 B.n736 B.n735 10.6151
R1094 B.n735 B.n734 10.6151
R1095 B.n734 B.n77 10.6151
R1096 B.n730 B.n77 10.6151
R1097 B.n730 B.n729 10.6151
R1098 B.n729 B.n728 10.6151
R1099 B.n728 B.n79 10.6151
R1100 B.n724 B.n79 10.6151
R1101 B.n724 B.n723 10.6151
R1102 B.n723 B.n722 10.6151
R1103 B.n722 B.n81 10.6151
R1104 B.n718 B.n81 10.6151
R1105 B.n718 B.n717 10.6151
R1106 B.n717 B.n716 10.6151
R1107 B.n716 B.n83 10.6151
R1108 B.n712 B.n83 10.6151
R1109 B.n712 B.n711 10.6151
R1110 B.n711 B.n710 10.6151
R1111 B.n710 B.n85 10.6151
R1112 B.n706 B.n85 10.6151
R1113 B.n706 B.n705 10.6151
R1114 B.n705 B.n704 10.6151
R1115 B.n704 B.n87 10.6151
R1116 B.n700 B.n699 10.6151
R1117 B.n699 B.n698 10.6151
R1118 B.n698 B.n89 10.6151
R1119 B.n694 B.n89 10.6151
R1120 B.n694 B.n693 10.6151
R1121 B.n693 B.n692 10.6151
R1122 B.n692 B.n91 10.6151
R1123 B.n688 B.n91 10.6151
R1124 B.n688 B.n687 10.6151
R1125 B.n687 B.n686 10.6151
R1126 B.n686 B.n93 10.6151
R1127 B.n682 B.n93 10.6151
R1128 B.n682 B.n681 10.6151
R1129 B.n681 B.n680 10.6151
R1130 B.n680 B.n95 10.6151
R1131 B.n676 B.n95 10.6151
R1132 B.n676 B.n675 10.6151
R1133 B.n675 B.n674 10.6151
R1134 B.n674 B.n97 10.6151
R1135 B.n670 B.n97 10.6151
R1136 B.n670 B.n669 10.6151
R1137 B.n669 B.n668 10.6151
R1138 B.n668 B.n99 10.6151
R1139 B.n664 B.n99 10.6151
R1140 B.n664 B.n663 10.6151
R1141 B.n663 B.n662 10.6151
R1142 B.n662 B.n101 10.6151
R1143 B.n658 B.n101 10.6151
R1144 B.n658 B.n657 10.6151
R1145 B.n657 B.n656 10.6151
R1146 B.n656 B.n103 10.6151
R1147 B.n652 B.n103 10.6151
R1148 B.n652 B.n651 10.6151
R1149 B.n651 B.n650 10.6151
R1150 B.n650 B.n105 10.6151
R1151 B.n646 B.n105 10.6151
R1152 B.n646 B.n645 10.6151
R1153 B.n645 B.n644 10.6151
R1154 B.n644 B.n107 10.6151
R1155 B.n640 B.n107 10.6151
R1156 B.n640 B.n639 10.6151
R1157 B.n639 B.n638 10.6151
R1158 B.n638 B.n109 10.6151
R1159 B.n634 B.n109 10.6151
R1160 B.n634 B.n633 10.6151
R1161 B.n633 B.n632 10.6151
R1162 B.n632 B.n111 10.6151
R1163 B.n628 B.n111 10.6151
R1164 B.n628 B.n627 10.6151
R1165 B.n627 B.n626 10.6151
R1166 B.n626 B.n113 10.6151
R1167 B.n622 B.n113 10.6151
R1168 B.n622 B.n621 10.6151
R1169 B.n621 B.n620 10.6151
R1170 B.n620 B.n115 10.6151
R1171 B.n616 B.n115 10.6151
R1172 B.n616 B.n615 10.6151
R1173 B.n615 B.n614 10.6151
R1174 B.n614 B.n117 10.6151
R1175 B.n610 B.n117 10.6151
R1176 B.n610 B.n609 10.6151
R1177 B.n609 B.n608 10.6151
R1178 B.n608 B.n119 10.6151
R1179 B.n604 B.n119 10.6151
R1180 B.n604 B.n603 10.6151
R1181 B.n603 B.n602 10.6151
R1182 B.n602 B.n121 10.6151
R1183 B.n598 B.n121 10.6151
R1184 B.n598 B.n597 10.6151
R1185 B.n597 B.n596 10.6151
R1186 B.n596 B.n123 10.6151
R1187 B.n592 B.n123 10.6151
R1188 B.n592 B.n591 10.6151
R1189 B.n591 B.n590 10.6151
R1190 B.n590 B.n125 10.6151
R1191 B.n586 B.n125 10.6151
R1192 B.n586 B.n585 10.6151
R1193 B.n585 B.n584 10.6151
R1194 B.n584 B.n127 10.6151
R1195 B.n580 B.n127 10.6151
R1196 B.n580 B.n579 10.6151
R1197 B.n579 B.n578 10.6151
R1198 B.n578 B.n129 10.6151
R1199 B.n574 B.n129 10.6151
R1200 B.n574 B.n573 10.6151
R1201 B.n573 B.n572 10.6151
R1202 B.n572 B.n131 10.6151
R1203 B.n568 B.n131 10.6151
R1204 B.n568 B.n567 10.6151
R1205 B.n567 B.n566 10.6151
R1206 B.n566 B.n133 10.6151
R1207 B.n562 B.n133 10.6151
R1208 B.n562 B.n561 10.6151
R1209 B.n561 B.n560 10.6151
R1210 B.n560 B.n135 10.6151
R1211 B.n556 B.n135 10.6151
R1212 B.n556 B.n555 10.6151
R1213 B.n555 B.n554 10.6151
R1214 B.n554 B.n137 10.6151
R1215 B.n550 B.n137 10.6151
R1216 B.n550 B.n549 10.6151
R1217 B.n549 B.n548 10.6151
R1218 B.n548 B.n139 10.6151
R1219 B.n544 B.n139 10.6151
R1220 B.n544 B.n543 10.6151
R1221 B.n543 B.n542 10.6151
R1222 B.n542 B.n141 10.6151
R1223 B.n538 B.n141 10.6151
R1224 B.n538 B.n537 10.6151
R1225 B.n537 B.n536 10.6151
R1226 B.n536 B.n143 10.6151
R1227 B.n532 B.n143 10.6151
R1228 B.n532 B.n531 10.6151
R1229 B.n531 B.n530 10.6151
R1230 B.n530 B.n145 10.6151
R1231 B.n526 B.n145 10.6151
R1232 B.n526 B.n525 10.6151
R1233 B.n525 B.n524 10.6151
R1234 B.n524 B.n147 10.6151
R1235 B.n520 B.n147 10.6151
R1236 B.n520 B.n519 10.6151
R1237 B.n519 B.n518 10.6151
R1238 B.n518 B.n149 10.6151
R1239 B.n514 B.n149 10.6151
R1240 B.n514 B.n513 10.6151
R1241 B.n513 B.n512 10.6151
R1242 B.n512 B.n151 10.6151
R1243 B.n508 B.n151 10.6151
R1244 B.n508 B.n507 10.6151
R1245 B.n507 B.n506 10.6151
R1246 B.n506 B.n153 10.6151
R1247 B.n502 B.n153 10.6151
R1248 B.n502 B.n501 10.6151
R1249 B.n501 B.n500 10.6151
R1250 B.n500 B.n155 10.6151
R1251 B.n496 B.n155 10.6151
R1252 B.n496 B.n495 10.6151
R1253 B.n495 B.n494 10.6151
R1254 B.n494 B.n157 10.6151
R1255 B.n490 B.n157 10.6151
R1256 B.n490 B.n489 10.6151
R1257 B.n489 B.n488 10.6151
R1258 B.n488 B.n159 10.6151
R1259 B.n241 B.n1 10.6151
R1260 B.n244 B.n241 10.6151
R1261 B.n245 B.n244 10.6151
R1262 B.n246 B.n245 10.6151
R1263 B.n246 B.n239 10.6151
R1264 B.n250 B.n239 10.6151
R1265 B.n251 B.n250 10.6151
R1266 B.n252 B.n251 10.6151
R1267 B.n252 B.n237 10.6151
R1268 B.n256 B.n237 10.6151
R1269 B.n257 B.n256 10.6151
R1270 B.n258 B.n257 10.6151
R1271 B.n258 B.n235 10.6151
R1272 B.n262 B.n235 10.6151
R1273 B.n263 B.n262 10.6151
R1274 B.n264 B.n263 10.6151
R1275 B.n264 B.n233 10.6151
R1276 B.n268 B.n233 10.6151
R1277 B.n269 B.n268 10.6151
R1278 B.n270 B.n269 10.6151
R1279 B.n270 B.n231 10.6151
R1280 B.n274 B.n231 10.6151
R1281 B.n275 B.n274 10.6151
R1282 B.n276 B.n275 10.6151
R1283 B.n276 B.n229 10.6151
R1284 B.n280 B.n229 10.6151
R1285 B.n281 B.n280 10.6151
R1286 B.n282 B.n281 10.6151
R1287 B.n282 B.n227 10.6151
R1288 B.n286 B.n227 10.6151
R1289 B.n287 B.n286 10.6151
R1290 B.n288 B.n287 10.6151
R1291 B.n288 B.n225 10.6151
R1292 B.n292 B.n225 10.6151
R1293 B.n293 B.n292 10.6151
R1294 B.n294 B.n293 10.6151
R1295 B.n294 B.n223 10.6151
R1296 B.n298 B.n223 10.6151
R1297 B.n299 B.n298 10.6151
R1298 B.n300 B.n299 10.6151
R1299 B.n300 B.n221 10.6151
R1300 B.n304 B.n221 10.6151
R1301 B.n305 B.n304 10.6151
R1302 B.n306 B.n305 10.6151
R1303 B.n306 B.n219 10.6151
R1304 B.n310 B.n219 10.6151
R1305 B.n311 B.n310 10.6151
R1306 B.n312 B.n311 10.6151
R1307 B.n312 B.n217 10.6151
R1308 B.n316 B.n217 10.6151
R1309 B.n317 B.n316 10.6151
R1310 B.n318 B.n317 10.6151
R1311 B.n318 B.n215 10.6151
R1312 B.n322 B.n215 10.6151
R1313 B.n323 B.n322 10.6151
R1314 B.n324 B.n323 10.6151
R1315 B.n324 B.n213 10.6151
R1316 B.n328 B.n213 10.6151
R1317 B.n329 B.n328 10.6151
R1318 B.n330 B.n329 10.6151
R1319 B.n330 B.n211 10.6151
R1320 B.n334 B.n211 10.6151
R1321 B.n335 B.n334 10.6151
R1322 B.n336 B.n335 10.6151
R1323 B.n336 B.n209 10.6151
R1324 B.n340 B.n209 10.6151
R1325 B.n341 B.n340 10.6151
R1326 B.n342 B.n341 10.6151
R1327 B.n342 B.n207 10.6151
R1328 B.n346 B.n207 10.6151
R1329 B.n348 B.n347 10.6151
R1330 B.n348 B.n205 10.6151
R1331 B.n352 B.n205 10.6151
R1332 B.n353 B.n352 10.6151
R1333 B.n354 B.n353 10.6151
R1334 B.n354 B.n203 10.6151
R1335 B.n358 B.n203 10.6151
R1336 B.n359 B.n358 10.6151
R1337 B.n360 B.n359 10.6151
R1338 B.n360 B.n201 10.6151
R1339 B.n364 B.n201 10.6151
R1340 B.n365 B.n364 10.6151
R1341 B.n366 B.n365 10.6151
R1342 B.n366 B.n199 10.6151
R1343 B.n370 B.n199 10.6151
R1344 B.n371 B.n370 10.6151
R1345 B.n372 B.n371 10.6151
R1346 B.n372 B.n197 10.6151
R1347 B.n376 B.n197 10.6151
R1348 B.n377 B.n376 10.6151
R1349 B.n378 B.n377 10.6151
R1350 B.n378 B.n195 10.6151
R1351 B.n382 B.n195 10.6151
R1352 B.n383 B.n382 10.6151
R1353 B.n384 B.n383 10.6151
R1354 B.n384 B.n193 10.6151
R1355 B.n388 B.n193 10.6151
R1356 B.n389 B.n388 10.6151
R1357 B.n390 B.n389 10.6151
R1358 B.n390 B.n191 10.6151
R1359 B.n394 B.n191 10.6151
R1360 B.n395 B.n394 10.6151
R1361 B.n396 B.n395 10.6151
R1362 B.n396 B.n189 10.6151
R1363 B.n400 B.n189 10.6151
R1364 B.n401 B.n400 10.6151
R1365 B.n402 B.n401 10.6151
R1366 B.n402 B.n187 10.6151
R1367 B.n406 B.n187 10.6151
R1368 B.n409 B.n408 10.6151
R1369 B.n409 B.n183 10.6151
R1370 B.n413 B.n183 10.6151
R1371 B.n414 B.n413 10.6151
R1372 B.n415 B.n414 10.6151
R1373 B.n415 B.n181 10.6151
R1374 B.n419 B.n181 10.6151
R1375 B.n420 B.n419 10.6151
R1376 B.n424 B.n420 10.6151
R1377 B.n428 B.n179 10.6151
R1378 B.n429 B.n428 10.6151
R1379 B.n430 B.n429 10.6151
R1380 B.n430 B.n177 10.6151
R1381 B.n434 B.n177 10.6151
R1382 B.n435 B.n434 10.6151
R1383 B.n436 B.n435 10.6151
R1384 B.n436 B.n175 10.6151
R1385 B.n440 B.n175 10.6151
R1386 B.n441 B.n440 10.6151
R1387 B.n442 B.n441 10.6151
R1388 B.n442 B.n173 10.6151
R1389 B.n446 B.n173 10.6151
R1390 B.n447 B.n446 10.6151
R1391 B.n448 B.n447 10.6151
R1392 B.n448 B.n171 10.6151
R1393 B.n452 B.n171 10.6151
R1394 B.n453 B.n452 10.6151
R1395 B.n454 B.n453 10.6151
R1396 B.n454 B.n169 10.6151
R1397 B.n458 B.n169 10.6151
R1398 B.n459 B.n458 10.6151
R1399 B.n460 B.n459 10.6151
R1400 B.n460 B.n167 10.6151
R1401 B.n464 B.n167 10.6151
R1402 B.n465 B.n464 10.6151
R1403 B.n466 B.n465 10.6151
R1404 B.n466 B.n165 10.6151
R1405 B.n470 B.n165 10.6151
R1406 B.n471 B.n470 10.6151
R1407 B.n472 B.n471 10.6151
R1408 B.n472 B.n163 10.6151
R1409 B.n476 B.n163 10.6151
R1410 B.n477 B.n476 10.6151
R1411 B.n478 B.n477 10.6151
R1412 B.n478 B.n161 10.6151
R1413 B.n482 B.n161 10.6151
R1414 B.n483 B.n482 10.6151
R1415 B.n484 B.n483 10.6151
R1416 B.n778 B.n777 9.36635
R1417 B.n760 B.n68 9.36635
R1418 B.n407 B.n406 9.36635
R1419 B.n423 B.n179 9.36635
R1420 B.n945 B.n0 8.11757
R1421 B.n945 B.n1 8.11757
R1422 B.n777 B.n776 1.24928
R1423 B.n68 B.n64 1.24928
R1424 B.n408 B.n407 1.24928
R1425 B.n424 B.n423 1.24928
R1426 VN.n96 VN.n95 161.3
R1427 VN.n94 VN.n50 161.3
R1428 VN.n93 VN.n92 161.3
R1429 VN.n91 VN.n51 161.3
R1430 VN.n90 VN.n89 161.3
R1431 VN.n88 VN.n52 161.3
R1432 VN.n87 VN.n86 161.3
R1433 VN.n85 VN.n84 161.3
R1434 VN.n83 VN.n54 161.3
R1435 VN.n82 VN.n81 161.3
R1436 VN.n80 VN.n55 161.3
R1437 VN.n79 VN.n78 161.3
R1438 VN.n77 VN.n56 161.3
R1439 VN.n76 VN.n75 161.3
R1440 VN.n74 VN.n57 161.3
R1441 VN.n73 VN.n72 161.3
R1442 VN.n71 VN.n58 161.3
R1443 VN.n70 VN.n69 161.3
R1444 VN.n68 VN.n59 161.3
R1445 VN.n67 VN.n66 161.3
R1446 VN.n65 VN.n60 161.3
R1447 VN.n64 VN.n63 161.3
R1448 VN.n47 VN.n46 161.3
R1449 VN.n45 VN.n1 161.3
R1450 VN.n44 VN.n43 161.3
R1451 VN.n42 VN.n2 161.3
R1452 VN.n41 VN.n40 161.3
R1453 VN.n39 VN.n3 161.3
R1454 VN.n38 VN.n37 161.3
R1455 VN.n36 VN.n35 161.3
R1456 VN.n34 VN.n5 161.3
R1457 VN.n33 VN.n32 161.3
R1458 VN.n31 VN.n6 161.3
R1459 VN.n30 VN.n29 161.3
R1460 VN.n28 VN.n7 161.3
R1461 VN.n27 VN.n26 161.3
R1462 VN.n25 VN.n8 161.3
R1463 VN.n24 VN.n23 161.3
R1464 VN.n22 VN.n9 161.3
R1465 VN.n21 VN.n20 161.3
R1466 VN.n19 VN.n10 161.3
R1467 VN.n18 VN.n17 161.3
R1468 VN.n16 VN.n11 161.3
R1469 VN.n15 VN.n14 161.3
R1470 VN.n62 VN.t3 117.587
R1471 VN.n13 VN.t2 117.587
R1472 VN.n8 VN.t9 85.6812
R1473 VN.n12 VN.t0 85.6812
R1474 VN.n4 VN.t1 85.6812
R1475 VN.n0 VN.t7 85.6812
R1476 VN.n57 VN.t8 85.6812
R1477 VN.n61 VN.t6 85.6812
R1478 VN.n53 VN.t4 85.6812
R1479 VN.n49 VN.t5 85.6812
R1480 VN.n48 VN.n0 81.2593
R1481 VN.n97 VN.n49 81.2593
R1482 VN.n13 VN.n12 70.1236
R1483 VN.n62 VN.n61 70.1236
R1484 VN VN.n97 56.57
R1485 VN.n21 VN.n10 56.5193
R1486 VN.n29 VN.n6 56.5193
R1487 VN.n70 VN.n59 56.5193
R1488 VN.n78 VN.n55 56.5193
R1489 VN.n40 VN.n2 51.663
R1490 VN.n89 VN.n51 51.663
R1491 VN.n44 VN.n2 29.3238
R1492 VN.n93 VN.n51 29.3238
R1493 VN.n16 VN.n15 24.4675
R1494 VN.n17 VN.n16 24.4675
R1495 VN.n17 VN.n10 24.4675
R1496 VN.n22 VN.n21 24.4675
R1497 VN.n23 VN.n22 24.4675
R1498 VN.n23 VN.n8 24.4675
R1499 VN.n27 VN.n8 24.4675
R1500 VN.n28 VN.n27 24.4675
R1501 VN.n29 VN.n28 24.4675
R1502 VN.n33 VN.n6 24.4675
R1503 VN.n34 VN.n33 24.4675
R1504 VN.n35 VN.n34 24.4675
R1505 VN.n39 VN.n38 24.4675
R1506 VN.n40 VN.n39 24.4675
R1507 VN.n45 VN.n44 24.4675
R1508 VN.n46 VN.n45 24.4675
R1509 VN.n66 VN.n59 24.4675
R1510 VN.n66 VN.n65 24.4675
R1511 VN.n65 VN.n64 24.4675
R1512 VN.n78 VN.n77 24.4675
R1513 VN.n77 VN.n76 24.4675
R1514 VN.n76 VN.n57 24.4675
R1515 VN.n72 VN.n57 24.4675
R1516 VN.n72 VN.n71 24.4675
R1517 VN.n71 VN.n70 24.4675
R1518 VN.n89 VN.n88 24.4675
R1519 VN.n88 VN.n87 24.4675
R1520 VN.n84 VN.n83 24.4675
R1521 VN.n83 VN.n82 24.4675
R1522 VN.n82 VN.n55 24.4675
R1523 VN.n95 VN.n94 24.4675
R1524 VN.n94 VN.n93 24.4675
R1525 VN.n38 VN.n4 20.0634
R1526 VN.n87 VN.n53 20.0634
R1527 VN.n46 VN.n0 8.80862
R1528 VN.n95 VN.n49 8.80862
R1529 VN.n63 VN.n62 4.46393
R1530 VN.n14 VN.n13 4.46393
R1531 VN.n15 VN.n12 4.40456
R1532 VN.n35 VN.n4 4.40456
R1533 VN.n64 VN.n61 4.40456
R1534 VN.n84 VN.n53 4.40456
R1535 VN.n97 VN.n96 0.354971
R1536 VN.n48 VN.n47 0.354971
R1537 VN VN.n48 0.26696
R1538 VN.n96 VN.n50 0.189894
R1539 VN.n92 VN.n50 0.189894
R1540 VN.n92 VN.n91 0.189894
R1541 VN.n91 VN.n90 0.189894
R1542 VN.n90 VN.n52 0.189894
R1543 VN.n86 VN.n52 0.189894
R1544 VN.n86 VN.n85 0.189894
R1545 VN.n85 VN.n54 0.189894
R1546 VN.n81 VN.n54 0.189894
R1547 VN.n81 VN.n80 0.189894
R1548 VN.n80 VN.n79 0.189894
R1549 VN.n79 VN.n56 0.189894
R1550 VN.n75 VN.n56 0.189894
R1551 VN.n75 VN.n74 0.189894
R1552 VN.n74 VN.n73 0.189894
R1553 VN.n73 VN.n58 0.189894
R1554 VN.n69 VN.n58 0.189894
R1555 VN.n69 VN.n68 0.189894
R1556 VN.n68 VN.n67 0.189894
R1557 VN.n67 VN.n60 0.189894
R1558 VN.n63 VN.n60 0.189894
R1559 VN.n14 VN.n11 0.189894
R1560 VN.n18 VN.n11 0.189894
R1561 VN.n19 VN.n18 0.189894
R1562 VN.n20 VN.n19 0.189894
R1563 VN.n20 VN.n9 0.189894
R1564 VN.n24 VN.n9 0.189894
R1565 VN.n25 VN.n24 0.189894
R1566 VN.n26 VN.n25 0.189894
R1567 VN.n26 VN.n7 0.189894
R1568 VN.n30 VN.n7 0.189894
R1569 VN.n31 VN.n30 0.189894
R1570 VN.n32 VN.n31 0.189894
R1571 VN.n32 VN.n5 0.189894
R1572 VN.n36 VN.n5 0.189894
R1573 VN.n37 VN.n36 0.189894
R1574 VN.n37 VN.n3 0.189894
R1575 VN.n41 VN.n3 0.189894
R1576 VN.n42 VN.n41 0.189894
R1577 VN.n43 VN.n42 0.189894
R1578 VN.n43 VN.n1 0.189894
R1579 VN.n47 VN.n1 0.189894
R1580 VDD2.n1 VDD2.t6 83.4184
R1581 VDD2.n4 VDD2.t3 80.3245
R1582 VDD2.n3 VDD2.n2 79.7847
R1583 VDD2 VDD2.n7 79.7817
R1584 VDD2.n6 VDD2.n5 77.52
R1585 VDD2.n1 VDD2.n0 77.5189
R1586 VDD2.n4 VDD2.n3 48.4071
R1587 VDD2.n6 VDD2.n4 3.09533
R1588 VDD2.n7 VDD2.t2 2.80507
R1589 VDD2.n7 VDD2.t7 2.80507
R1590 VDD2.n5 VDD2.t4 2.80507
R1591 VDD2.n5 VDD2.t5 2.80507
R1592 VDD2.n2 VDD2.t1 2.80507
R1593 VDD2.n2 VDD2.t8 2.80507
R1594 VDD2.n0 VDD2.t9 2.80507
R1595 VDD2.n0 VDD2.t0 2.80507
R1596 VDD2 VDD2.n6 0.832397
R1597 VDD2.n3 VDD2.n1 0.718861
R1598 VTAIL.n11 VTAIL.t16 63.6457
R1599 VTAIL.n17 VTAIL.t12 63.6447
R1600 VTAIL.n2 VTAIL.t6 63.6447
R1601 VTAIL.n16 VTAIL.t9 63.6446
R1602 VTAIL.n15 VTAIL.n14 60.8412
R1603 VTAIL.n13 VTAIL.n12 60.8412
R1604 VTAIL.n10 VTAIL.n9 60.8412
R1605 VTAIL.n8 VTAIL.n7 60.8412
R1606 VTAIL.n19 VTAIL.n18 60.8401
R1607 VTAIL.n1 VTAIL.n0 60.8401
R1608 VTAIL.n4 VTAIL.n3 60.8401
R1609 VTAIL.n6 VTAIL.n5 60.8401
R1610 VTAIL.n8 VTAIL.n6 28.5479
R1611 VTAIL.n17 VTAIL.n16 25.4531
R1612 VTAIL.n10 VTAIL.n8 3.09533
R1613 VTAIL.n11 VTAIL.n10 3.09533
R1614 VTAIL.n15 VTAIL.n13 3.09533
R1615 VTAIL.n16 VTAIL.n15 3.09533
R1616 VTAIL.n6 VTAIL.n4 3.09533
R1617 VTAIL.n4 VTAIL.n2 3.09533
R1618 VTAIL.n19 VTAIL.n17 3.09533
R1619 VTAIL.n18 VTAIL.t10 2.80507
R1620 VTAIL.n18 VTAIL.t18 2.80507
R1621 VTAIL.n0 VTAIL.t17 2.80507
R1622 VTAIL.n0 VTAIL.t19 2.80507
R1623 VTAIL.n3 VTAIL.t3 2.80507
R1624 VTAIL.n3 VTAIL.t7 2.80507
R1625 VTAIL.n5 VTAIL.t2 2.80507
R1626 VTAIL.n5 VTAIL.t5 2.80507
R1627 VTAIL.n14 VTAIL.t1 2.80507
R1628 VTAIL.n14 VTAIL.t8 2.80507
R1629 VTAIL.n12 VTAIL.t4 2.80507
R1630 VTAIL.n12 VTAIL.t0 2.80507
R1631 VTAIL.n9 VTAIL.t11 2.80507
R1632 VTAIL.n9 VTAIL.t13 2.80507
R1633 VTAIL.n7 VTAIL.t14 2.80507
R1634 VTAIL.n7 VTAIL.t15 2.80507
R1635 VTAIL VTAIL.n1 2.37981
R1636 VTAIL.n13 VTAIL.n11 2.01774
R1637 VTAIL.n2 VTAIL.n1 2.01774
R1638 VTAIL VTAIL.n19 0.716017
R1639 VP.n32 VP.n31 161.3
R1640 VP.n33 VP.n28 161.3
R1641 VP.n35 VP.n34 161.3
R1642 VP.n36 VP.n27 161.3
R1643 VP.n38 VP.n37 161.3
R1644 VP.n39 VP.n26 161.3
R1645 VP.n41 VP.n40 161.3
R1646 VP.n42 VP.n25 161.3
R1647 VP.n44 VP.n43 161.3
R1648 VP.n45 VP.n24 161.3
R1649 VP.n47 VP.n46 161.3
R1650 VP.n48 VP.n23 161.3
R1651 VP.n50 VP.n49 161.3
R1652 VP.n51 VP.n22 161.3
R1653 VP.n53 VP.n52 161.3
R1654 VP.n55 VP.n54 161.3
R1655 VP.n56 VP.n20 161.3
R1656 VP.n58 VP.n57 161.3
R1657 VP.n59 VP.n19 161.3
R1658 VP.n61 VP.n60 161.3
R1659 VP.n62 VP.n18 161.3
R1660 VP.n64 VP.n63 161.3
R1661 VP.n111 VP.n110 161.3
R1662 VP.n109 VP.n1 161.3
R1663 VP.n108 VP.n107 161.3
R1664 VP.n106 VP.n2 161.3
R1665 VP.n105 VP.n104 161.3
R1666 VP.n103 VP.n3 161.3
R1667 VP.n102 VP.n101 161.3
R1668 VP.n100 VP.n99 161.3
R1669 VP.n98 VP.n5 161.3
R1670 VP.n97 VP.n96 161.3
R1671 VP.n95 VP.n6 161.3
R1672 VP.n94 VP.n93 161.3
R1673 VP.n92 VP.n7 161.3
R1674 VP.n91 VP.n90 161.3
R1675 VP.n89 VP.n8 161.3
R1676 VP.n88 VP.n87 161.3
R1677 VP.n86 VP.n9 161.3
R1678 VP.n85 VP.n84 161.3
R1679 VP.n83 VP.n10 161.3
R1680 VP.n82 VP.n81 161.3
R1681 VP.n80 VP.n11 161.3
R1682 VP.n79 VP.n78 161.3
R1683 VP.n77 VP.n76 161.3
R1684 VP.n75 VP.n13 161.3
R1685 VP.n74 VP.n73 161.3
R1686 VP.n72 VP.n14 161.3
R1687 VP.n71 VP.n70 161.3
R1688 VP.n69 VP.n15 161.3
R1689 VP.n68 VP.n67 161.3
R1690 VP.n30 VP.t4 117.587
R1691 VP.n8 VP.t1 85.6812
R1692 VP.n16 VP.t3 85.6812
R1693 VP.n12 VP.t8 85.6812
R1694 VP.n4 VP.t9 85.6812
R1695 VP.n0 VP.t0 85.6812
R1696 VP.n25 VP.t5 85.6812
R1697 VP.n17 VP.t2 85.6812
R1698 VP.n21 VP.t6 85.6812
R1699 VP.n29 VP.t7 85.6812
R1700 VP.n66 VP.n16 81.2593
R1701 VP.n112 VP.n0 81.2593
R1702 VP.n65 VP.n17 81.2593
R1703 VP.n30 VP.n29 70.1236
R1704 VP.n85 VP.n10 56.5193
R1705 VP.n93 VP.n6 56.5193
R1706 VP.n46 VP.n23 56.5193
R1707 VP.n38 VP.n27 56.5193
R1708 VP.n66 VP.n65 56.4046
R1709 VP.n74 VP.n14 51.663
R1710 VP.n104 VP.n2 51.663
R1711 VP.n57 VP.n19 51.663
R1712 VP.n70 VP.n14 29.3238
R1713 VP.n108 VP.n2 29.3238
R1714 VP.n61 VP.n19 29.3238
R1715 VP.n69 VP.n68 24.4675
R1716 VP.n70 VP.n69 24.4675
R1717 VP.n75 VP.n74 24.4675
R1718 VP.n76 VP.n75 24.4675
R1719 VP.n80 VP.n79 24.4675
R1720 VP.n81 VP.n80 24.4675
R1721 VP.n81 VP.n10 24.4675
R1722 VP.n86 VP.n85 24.4675
R1723 VP.n87 VP.n86 24.4675
R1724 VP.n87 VP.n8 24.4675
R1725 VP.n91 VP.n8 24.4675
R1726 VP.n92 VP.n91 24.4675
R1727 VP.n93 VP.n92 24.4675
R1728 VP.n97 VP.n6 24.4675
R1729 VP.n98 VP.n97 24.4675
R1730 VP.n99 VP.n98 24.4675
R1731 VP.n103 VP.n102 24.4675
R1732 VP.n104 VP.n103 24.4675
R1733 VP.n109 VP.n108 24.4675
R1734 VP.n110 VP.n109 24.4675
R1735 VP.n62 VP.n61 24.4675
R1736 VP.n63 VP.n62 24.4675
R1737 VP.n50 VP.n23 24.4675
R1738 VP.n51 VP.n50 24.4675
R1739 VP.n52 VP.n51 24.4675
R1740 VP.n56 VP.n55 24.4675
R1741 VP.n57 VP.n56 24.4675
R1742 VP.n39 VP.n38 24.4675
R1743 VP.n40 VP.n39 24.4675
R1744 VP.n40 VP.n25 24.4675
R1745 VP.n44 VP.n25 24.4675
R1746 VP.n45 VP.n44 24.4675
R1747 VP.n46 VP.n45 24.4675
R1748 VP.n33 VP.n32 24.4675
R1749 VP.n34 VP.n33 24.4675
R1750 VP.n34 VP.n27 24.4675
R1751 VP.n76 VP.n12 20.0634
R1752 VP.n102 VP.n4 20.0634
R1753 VP.n55 VP.n21 20.0634
R1754 VP.n68 VP.n16 8.80862
R1755 VP.n110 VP.n0 8.80862
R1756 VP.n63 VP.n17 8.80862
R1757 VP.n31 VP.n30 4.46391
R1758 VP.n79 VP.n12 4.40456
R1759 VP.n99 VP.n4 4.40456
R1760 VP.n52 VP.n21 4.40456
R1761 VP.n32 VP.n29 4.40456
R1762 VP.n65 VP.n64 0.354971
R1763 VP.n67 VP.n66 0.354971
R1764 VP.n112 VP.n111 0.354971
R1765 VP VP.n112 0.26696
R1766 VP.n31 VP.n28 0.189894
R1767 VP.n35 VP.n28 0.189894
R1768 VP.n36 VP.n35 0.189894
R1769 VP.n37 VP.n36 0.189894
R1770 VP.n37 VP.n26 0.189894
R1771 VP.n41 VP.n26 0.189894
R1772 VP.n42 VP.n41 0.189894
R1773 VP.n43 VP.n42 0.189894
R1774 VP.n43 VP.n24 0.189894
R1775 VP.n47 VP.n24 0.189894
R1776 VP.n48 VP.n47 0.189894
R1777 VP.n49 VP.n48 0.189894
R1778 VP.n49 VP.n22 0.189894
R1779 VP.n53 VP.n22 0.189894
R1780 VP.n54 VP.n53 0.189894
R1781 VP.n54 VP.n20 0.189894
R1782 VP.n58 VP.n20 0.189894
R1783 VP.n59 VP.n58 0.189894
R1784 VP.n60 VP.n59 0.189894
R1785 VP.n60 VP.n18 0.189894
R1786 VP.n64 VP.n18 0.189894
R1787 VP.n67 VP.n15 0.189894
R1788 VP.n71 VP.n15 0.189894
R1789 VP.n72 VP.n71 0.189894
R1790 VP.n73 VP.n72 0.189894
R1791 VP.n73 VP.n13 0.189894
R1792 VP.n77 VP.n13 0.189894
R1793 VP.n78 VP.n77 0.189894
R1794 VP.n78 VP.n11 0.189894
R1795 VP.n82 VP.n11 0.189894
R1796 VP.n83 VP.n82 0.189894
R1797 VP.n84 VP.n83 0.189894
R1798 VP.n84 VP.n9 0.189894
R1799 VP.n88 VP.n9 0.189894
R1800 VP.n89 VP.n88 0.189894
R1801 VP.n90 VP.n89 0.189894
R1802 VP.n90 VP.n7 0.189894
R1803 VP.n94 VP.n7 0.189894
R1804 VP.n95 VP.n94 0.189894
R1805 VP.n96 VP.n95 0.189894
R1806 VP.n96 VP.n5 0.189894
R1807 VP.n100 VP.n5 0.189894
R1808 VP.n101 VP.n100 0.189894
R1809 VP.n101 VP.n3 0.189894
R1810 VP.n105 VP.n3 0.189894
R1811 VP.n106 VP.n105 0.189894
R1812 VP.n107 VP.n106 0.189894
R1813 VP.n107 VP.n1 0.189894
R1814 VP.n111 VP.n1 0.189894
R1815 VDD1.n1 VDD1.t5 83.4193
R1816 VDD1.n3 VDD1.t6 83.4184
R1817 VDD1.n5 VDD1.n4 79.7847
R1818 VDD1.n1 VDD1.n0 77.52
R1819 VDD1.n3 VDD1.n2 77.5189
R1820 VDD1.n7 VDD1.n6 77.5188
R1821 VDD1.n7 VDD1.n5 50.5375
R1822 VDD1.n6 VDD1.t3 2.80507
R1823 VDD1.n6 VDD1.t7 2.80507
R1824 VDD1.n0 VDD1.t2 2.80507
R1825 VDD1.n0 VDD1.t4 2.80507
R1826 VDD1.n4 VDD1.t0 2.80507
R1827 VDD1.n4 VDD1.t9 2.80507
R1828 VDD1.n2 VDD1.t1 2.80507
R1829 VDD1.n2 VDD1.t8 2.80507
R1830 VDD1 VDD1.n7 2.26343
R1831 VDD1 VDD1.n1 0.832397
R1832 VDD1.n5 VDD1.n3 0.718861
C0 VTAIL w_n5278_n3286# 3.25154f
C1 VDD2 VTAIL 10.5426f
C2 B VDD1 2.70486f
C3 VDD2 w_n5278_n3286# 3.19051f
C4 VP VDD1 11.257401f
C5 B VTAIL 3.89386f
C6 VP VTAIL 11.7072f
C7 B w_n5278_n3286# 11.5415f
C8 VDD2 B 2.84847f
C9 VP w_n5278_n3286# 12.181901f
C10 VDD2 VP 0.667831f
C11 VN VDD1 0.154942f
C12 VN VTAIL 11.693f
C13 B VP 2.60903f
C14 VN w_n5278_n3286# 11.492701f
C15 VDD2 VN 10.7483f
C16 VTAIL VDD1 10.4865f
C17 B VN 1.44645f
C18 VDD1 w_n5278_n3286# 3.01266f
C19 VDD2 VDD1 2.60476f
C20 VP VN 9.30119f
C21 VDD2 VSUBS 2.37975f
C22 VDD1 VSUBS 2.222678f
C23 VTAIL VSUBS 1.44887f
C24 VN VSUBS 8.77483f
C25 VP VSUBS 5.066479f
C26 B VSUBS 6.15068f
C27 w_n5278_n3286# VSUBS 0.213632p
C28 VDD1.t5 VSUBS 2.93974f
C29 VDD1.t2 VSUBS 0.283388f
C30 VDD1.t4 VSUBS 0.283388f
C31 VDD1.n0 VSUBS 2.22587f
C32 VDD1.n1 VSUBS 1.87021f
C33 VDD1.t6 VSUBS 2.93974f
C34 VDD1.t1 VSUBS 0.283388f
C35 VDD1.t8 VSUBS 0.283388f
C36 VDD1.n2 VSUBS 2.22587f
C37 VDD1.n3 VSUBS 1.85989f
C38 VDD1.t0 VSUBS 0.283388f
C39 VDD1.t9 VSUBS 0.283388f
C40 VDD1.n4 VSUBS 2.25701f
C41 VDD1.n5 VSUBS 4.45813f
C42 VDD1.t3 VSUBS 0.283388f
C43 VDD1.t7 VSUBS 0.283388f
C44 VDD1.n6 VSUBS 2.22586f
C45 VDD1.n7 VSUBS 4.52202f
C46 VP.t0 VSUBS 2.84379f
C47 VP.n0 VSUBS 1.09955f
C48 VP.n1 VSUBS 0.027652f
C49 VP.n2 VSUBS 0.027439f
C50 VP.n3 VSUBS 0.027652f
C51 VP.t9 VSUBS 2.84379f
C52 VP.n4 VSUBS 1.00144f
C53 VP.n5 VSUBS 0.027652f
C54 VP.n6 VSUBS 0.036902f
C55 VP.n7 VSUBS 0.027652f
C56 VP.t1 VSUBS 2.84379f
C57 VP.n8 VSUBS 1.02754f
C58 VP.n9 VSUBS 0.027652f
C59 VP.n10 VSUBS 0.036902f
C60 VP.n11 VSUBS 0.027652f
C61 VP.t8 VSUBS 2.84379f
C62 VP.n12 VSUBS 1.00144f
C63 VP.n13 VSUBS 0.027652f
C64 VP.n14 VSUBS 0.027439f
C65 VP.n15 VSUBS 0.027652f
C66 VP.t3 VSUBS 2.84379f
C67 VP.n16 VSUBS 1.09955f
C68 VP.t2 VSUBS 2.84379f
C69 VP.n17 VSUBS 1.09955f
C70 VP.n18 VSUBS 0.027652f
C71 VP.n19 VSUBS 0.027439f
C72 VP.n20 VSUBS 0.027652f
C73 VP.t6 VSUBS 2.84379f
C74 VP.n21 VSUBS 1.00144f
C75 VP.n22 VSUBS 0.027652f
C76 VP.n23 VSUBS 0.036902f
C77 VP.n24 VSUBS 0.027652f
C78 VP.t5 VSUBS 2.84379f
C79 VP.n25 VSUBS 1.02754f
C80 VP.n26 VSUBS 0.027652f
C81 VP.n27 VSUBS 0.036902f
C82 VP.n28 VSUBS 0.027652f
C83 VP.t7 VSUBS 2.84379f
C84 VP.n29 VSUBS 1.08626f
C85 VP.t4 VSUBS 3.16733f
C86 VP.n30 VSUBS 1.04268f
C87 VP.n31 VSUBS 0.325733f
C88 VP.n32 VSUBS 0.030673f
C89 VP.n33 VSUBS 0.051537f
C90 VP.n34 VSUBS 0.051537f
C91 VP.n35 VSUBS 0.027652f
C92 VP.n36 VSUBS 0.027652f
C93 VP.n37 VSUBS 0.027652f
C94 VP.n38 VSUBS 0.043837f
C95 VP.n39 VSUBS 0.051537f
C96 VP.n40 VSUBS 0.051537f
C97 VP.n41 VSUBS 0.027652f
C98 VP.n42 VSUBS 0.027652f
C99 VP.n43 VSUBS 0.027652f
C100 VP.n44 VSUBS 0.051537f
C101 VP.n45 VSUBS 0.051537f
C102 VP.n46 VSUBS 0.043837f
C103 VP.n47 VSUBS 0.027652f
C104 VP.n48 VSUBS 0.027652f
C105 VP.n49 VSUBS 0.027652f
C106 VP.n50 VSUBS 0.051537f
C107 VP.n51 VSUBS 0.051537f
C108 VP.n52 VSUBS 0.030673f
C109 VP.n53 VSUBS 0.027652f
C110 VP.n54 VSUBS 0.027652f
C111 VP.n55 VSUBS 0.046957f
C112 VP.n56 VSUBS 0.051537f
C113 VP.n57 VSUBS 0.049929f
C114 VP.n58 VSUBS 0.027652f
C115 VP.n59 VSUBS 0.027652f
C116 VP.n60 VSUBS 0.027652f
C117 VP.n61 VSUBS 0.054908f
C118 VP.n62 VSUBS 0.051537f
C119 VP.n63 VSUBS 0.035253f
C120 VP.n64 VSUBS 0.04463f
C121 VP.n65 VSUBS 1.86515f
C122 VP.n66 VSUBS 1.88277f
C123 VP.n67 VSUBS 0.04463f
C124 VP.n68 VSUBS 0.035253f
C125 VP.n69 VSUBS 0.051537f
C126 VP.n70 VSUBS 0.054908f
C127 VP.n71 VSUBS 0.027652f
C128 VP.n72 VSUBS 0.027652f
C129 VP.n73 VSUBS 0.027652f
C130 VP.n74 VSUBS 0.049929f
C131 VP.n75 VSUBS 0.051537f
C132 VP.n76 VSUBS 0.046957f
C133 VP.n77 VSUBS 0.027652f
C134 VP.n78 VSUBS 0.027652f
C135 VP.n79 VSUBS 0.030673f
C136 VP.n80 VSUBS 0.051537f
C137 VP.n81 VSUBS 0.051537f
C138 VP.n82 VSUBS 0.027652f
C139 VP.n83 VSUBS 0.027652f
C140 VP.n84 VSUBS 0.027652f
C141 VP.n85 VSUBS 0.043837f
C142 VP.n86 VSUBS 0.051537f
C143 VP.n87 VSUBS 0.051537f
C144 VP.n88 VSUBS 0.027652f
C145 VP.n89 VSUBS 0.027652f
C146 VP.n90 VSUBS 0.027652f
C147 VP.n91 VSUBS 0.051537f
C148 VP.n92 VSUBS 0.051537f
C149 VP.n93 VSUBS 0.043837f
C150 VP.n94 VSUBS 0.027652f
C151 VP.n95 VSUBS 0.027652f
C152 VP.n96 VSUBS 0.027652f
C153 VP.n97 VSUBS 0.051537f
C154 VP.n98 VSUBS 0.051537f
C155 VP.n99 VSUBS 0.030673f
C156 VP.n100 VSUBS 0.027652f
C157 VP.n101 VSUBS 0.027652f
C158 VP.n102 VSUBS 0.046957f
C159 VP.n103 VSUBS 0.051537f
C160 VP.n104 VSUBS 0.049929f
C161 VP.n105 VSUBS 0.027652f
C162 VP.n106 VSUBS 0.027652f
C163 VP.n107 VSUBS 0.027652f
C164 VP.n108 VSUBS 0.054908f
C165 VP.n109 VSUBS 0.051537f
C166 VP.n110 VSUBS 0.035253f
C167 VP.n111 VSUBS 0.04463f
C168 VP.n112 VSUBS 0.072167f
C169 VTAIL.t17 VSUBS 0.272396f
C170 VTAIL.t19 VSUBS 0.272396f
C171 VTAIL.n0 VSUBS 1.99633f
C172 VTAIL.n1 VSUBS 1.05216f
C173 VTAIL.t6 VSUBS 2.63052f
C174 VTAIL.n2 VSUBS 1.22943f
C175 VTAIL.t3 VSUBS 0.272396f
C176 VTAIL.t7 VSUBS 0.272396f
C177 VTAIL.n3 VSUBS 1.99633f
C178 VTAIL.n4 VSUBS 1.224f
C179 VTAIL.t2 VSUBS 0.272396f
C180 VTAIL.t5 VSUBS 0.272396f
C181 VTAIL.n5 VSUBS 1.99633f
C182 VTAIL.n6 VSUBS 2.88211f
C183 VTAIL.t14 VSUBS 0.272396f
C184 VTAIL.t15 VSUBS 0.272396f
C185 VTAIL.n7 VSUBS 1.99633f
C186 VTAIL.n8 VSUBS 2.8821f
C187 VTAIL.t11 VSUBS 0.272396f
C188 VTAIL.t13 VSUBS 0.272396f
C189 VTAIL.n9 VSUBS 1.99633f
C190 VTAIL.n10 VSUBS 1.224f
C191 VTAIL.t16 VSUBS 2.63053f
C192 VTAIL.n11 VSUBS 1.22943f
C193 VTAIL.t4 VSUBS 0.272396f
C194 VTAIL.t0 VSUBS 0.272396f
C195 VTAIL.n12 VSUBS 1.99633f
C196 VTAIL.n13 VSUBS 1.12073f
C197 VTAIL.t1 VSUBS 0.272396f
C198 VTAIL.t8 VSUBS 0.272396f
C199 VTAIL.n14 VSUBS 1.99633f
C200 VTAIL.n15 VSUBS 1.224f
C201 VTAIL.t9 VSUBS 2.63051f
C202 VTAIL.n16 VSUBS 2.69423f
C203 VTAIL.t12 VSUBS 2.63052f
C204 VTAIL.n17 VSUBS 2.69422f
C205 VTAIL.t10 VSUBS 0.272396f
C206 VTAIL.t18 VSUBS 0.272396f
C207 VTAIL.n18 VSUBS 1.99633f
C208 VTAIL.n19 VSUBS 0.995979f
C209 VDD2.t6 VSUBS 2.92153f
C210 VDD2.t9 VSUBS 0.281633f
C211 VDD2.t0 VSUBS 0.281633f
C212 VDD2.n0 VSUBS 2.21208f
C213 VDD2.n1 VSUBS 1.84837f
C214 VDD2.t1 VSUBS 0.281633f
C215 VDD2.t8 VSUBS 0.281633f
C216 VDD2.n2 VSUBS 2.24303f
C217 VDD2.n3 VSUBS 4.25492f
C218 VDD2.t3 VSUBS 2.88595f
C219 VDD2.n4 VSUBS 4.42603f
C220 VDD2.t4 VSUBS 0.281633f
C221 VDD2.t5 VSUBS 0.281633f
C222 VDD2.n5 VSUBS 2.21208f
C223 VDD2.n6 VSUBS 0.935017f
C224 VDD2.t2 VSUBS 0.281633f
C225 VDD2.t7 VSUBS 0.281633f
C226 VDD2.n7 VSUBS 2.24297f
C227 VN.t7 VSUBS 2.60616f
C228 VN.n0 VSUBS 1.00767f
C229 VN.n1 VSUBS 0.025342f
C230 VN.n2 VSUBS 0.025146f
C231 VN.n3 VSUBS 0.025342f
C232 VN.t1 VSUBS 2.60616f
C233 VN.n4 VSUBS 0.917764f
C234 VN.n5 VSUBS 0.025342f
C235 VN.n6 VSUBS 0.033819f
C236 VN.n7 VSUBS 0.025342f
C237 VN.t9 VSUBS 2.60616f
C238 VN.n8 VSUBS 0.941677f
C239 VN.n9 VSUBS 0.025342f
C240 VN.n10 VSUBS 0.033819f
C241 VN.n11 VSUBS 0.025342f
C242 VN.t0 VSUBS 2.60616f
C243 VN.n12 VSUBS 0.995497f
C244 VN.t2 VSUBS 2.90267f
C245 VN.n13 VSUBS 0.955557f
C246 VN.n14 VSUBS 0.298515f
C247 VN.n15 VSUBS 0.02811f
C248 VN.n16 VSUBS 0.04723f
C249 VN.n17 VSUBS 0.04723f
C250 VN.n18 VSUBS 0.025342f
C251 VN.n19 VSUBS 0.025342f
C252 VN.n20 VSUBS 0.025342f
C253 VN.n21 VSUBS 0.040174f
C254 VN.n22 VSUBS 0.04723f
C255 VN.n23 VSUBS 0.04723f
C256 VN.n24 VSUBS 0.025342f
C257 VN.n25 VSUBS 0.025342f
C258 VN.n26 VSUBS 0.025342f
C259 VN.n27 VSUBS 0.04723f
C260 VN.n28 VSUBS 0.04723f
C261 VN.n29 VSUBS 0.040174f
C262 VN.n30 VSUBS 0.025342f
C263 VN.n31 VSUBS 0.025342f
C264 VN.n32 VSUBS 0.025342f
C265 VN.n33 VSUBS 0.04723f
C266 VN.n34 VSUBS 0.04723f
C267 VN.n35 VSUBS 0.02811f
C268 VN.n36 VSUBS 0.025342f
C269 VN.n37 VSUBS 0.025342f
C270 VN.n38 VSUBS 0.043033f
C271 VN.n39 VSUBS 0.04723f
C272 VN.n40 VSUBS 0.045757f
C273 VN.n41 VSUBS 0.025342f
C274 VN.n42 VSUBS 0.025342f
C275 VN.n43 VSUBS 0.025342f
C276 VN.n44 VSUBS 0.05032f
C277 VN.n45 VSUBS 0.04723f
C278 VN.n46 VSUBS 0.032307f
C279 VN.n47 VSUBS 0.040901f
C280 VN.n48 VSUBS 0.066137f
C281 VN.t5 VSUBS 2.60616f
C282 VN.n49 VSUBS 1.00767f
C283 VN.n50 VSUBS 0.025342f
C284 VN.n51 VSUBS 0.025146f
C285 VN.n52 VSUBS 0.025342f
C286 VN.t4 VSUBS 2.60616f
C287 VN.n53 VSUBS 0.917764f
C288 VN.n54 VSUBS 0.025342f
C289 VN.n55 VSUBS 0.033819f
C290 VN.n56 VSUBS 0.025342f
C291 VN.t8 VSUBS 2.60616f
C292 VN.n57 VSUBS 0.941677f
C293 VN.n58 VSUBS 0.025342f
C294 VN.n59 VSUBS 0.033819f
C295 VN.n60 VSUBS 0.025342f
C296 VN.t6 VSUBS 2.60616f
C297 VN.n61 VSUBS 0.995497f
C298 VN.t3 VSUBS 2.90267f
C299 VN.n62 VSUBS 0.955557f
C300 VN.n63 VSUBS 0.298515f
C301 VN.n64 VSUBS 0.02811f
C302 VN.n65 VSUBS 0.04723f
C303 VN.n66 VSUBS 0.04723f
C304 VN.n67 VSUBS 0.025342f
C305 VN.n68 VSUBS 0.025342f
C306 VN.n69 VSUBS 0.025342f
C307 VN.n70 VSUBS 0.040174f
C308 VN.n71 VSUBS 0.04723f
C309 VN.n72 VSUBS 0.04723f
C310 VN.n73 VSUBS 0.025342f
C311 VN.n74 VSUBS 0.025342f
C312 VN.n75 VSUBS 0.025342f
C313 VN.n76 VSUBS 0.04723f
C314 VN.n77 VSUBS 0.04723f
C315 VN.n78 VSUBS 0.040174f
C316 VN.n79 VSUBS 0.025342f
C317 VN.n80 VSUBS 0.025342f
C318 VN.n81 VSUBS 0.025342f
C319 VN.n82 VSUBS 0.04723f
C320 VN.n83 VSUBS 0.04723f
C321 VN.n84 VSUBS 0.02811f
C322 VN.n85 VSUBS 0.025342f
C323 VN.n86 VSUBS 0.025342f
C324 VN.n87 VSUBS 0.043033f
C325 VN.n88 VSUBS 0.04723f
C326 VN.n89 VSUBS 0.045757f
C327 VN.n90 VSUBS 0.025342f
C328 VN.n91 VSUBS 0.025342f
C329 VN.n92 VSUBS 0.025342f
C330 VN.n93 VSUBS 0.05032f
C331 VN.n94 VSUBS 0.04723f
C332 VN.n95 VSUBS 0.032307f
C333 VN.n96 VSUBS 0.040901f
C334 VN.n97 VSUBS 1.71927f
C335 B.n0 VSUBS 0.008033f
C336 B.n1 VSUBS 0.008033f
C337 B.n2 VSUBS 0.01188f
C338 B.n3 VSUBS 0.009104f
C339 B.n4 VSUBS 0.009104f
C340 B.n5 VSUBS 0.009104f
C341 B.n6 VSUBS 0.009104f
C342 B.n7 VSUBS 0.009104f
C343 B.n8 VSUBS 0.009104f
C344 B.n9 VSUBS 0.009104f
C345 B.n10 VSUBS 0.009104f
C346 B.n11 VSUBS 0.009104f
C347 B.n12 VSUBS 0.009104f
C348 B.n13 VSUBS 0.009104f
C349 B.n14 VSUBS 0.009104f
C350 B.n15 VSUBS 0.009104f
C351 B.n16 VSUBS 0.009104f
C352 B.n17 VSUBS 0.009104f
C353 B.n18 VSUBS 0.009104f
C354 B.n19 VSUBS 0.009104f
C355 B.n20 VSUBS 0.009104f
C356 B.n21 VSUBS 0.009104f
C357 B.n22 VSUBS 0.009104f
C358 B.n23 VSUBS 0.009104f
C359 B.n24 VSUBS 0.009104f
C360 B.n25 VSUBS 0.009104f
C361 B.n26 VSUBS 0.009104f
C362 B.n27 VSUBS 0.009104f
C363 B.n28 VSUBS 0.009104f
C364 B.n29 VSUBS 0.009104f
C365 B.n30 VSUBS 0.009104f
C366 B.n31 VSUBS 0.009104f
C367 B.n32 VSUBS 0.009104f
C368 B.n33 VSUBS 0.009104f
C369 B.n34 VSUBS 0.009104f
C370 B.n35 VSUBS 0.009104f
C371 B.n36 VSUBS 0.009104f
C372 B.n37 VSUBS 0.021667f
C373 B.n38 VSUBS 0.009104f
C374 B.n39 VSUBS 0.009104f
C375 B.n40 VSUBS 0.009104f
C376 B.n41 VSUBS 0.009104f
C377 B.n42 VSUBS 0.009104f
C378 B.n43 VSUBS 0.009104f
C379 B.n44 VSUBS 0.009104f
C380 B.n45 VSUBS 0.009104f
C381 B.n46 VSUBS 0.009104f
C382 B.n47 VSUBS 0.009104f
C383 B.n48 VSUBS 0.009104f
C384 B.n49 VSUBS 0.009104f
C385 B.n50 VSUBS 0.009104f
C386 B.n51 VSUBS 0.009104f
C387 B.n52 VSUBS 0.009104f
C388 B.n53 VSUBS 0.009104f
C389 B.n54 VSUBS 0.009104f
C390 B.n55 VSUBS 0.009104f
C391 B.n56 VSUBS 0.009104f
C392 B.n57 VSUBS 0.009104f
C393 B.t7 VSUBS 0.489322f
C394 B.t8 VSUBS 0.522261f
C395 B.t6 VSUBS 2.27548f
C396 B.n58 VSUBS 0.28876f
C397 B.n59 VSUBS 0.096909f
C398 B.n60 VSUBS 0.009104f
C399 B.n61 VSUBS 0.009104f
C400 B.n62 VSUBS 0.009104f
C401 B.n63 VSUBS 0.009104f
C402 B.n64 VSUBS 0.005087f
C403 B.n65 VSUBS 0.009104f
C404 B.t1 VSUBS 0.489313f
C405 B.t2 VSUBS 0.522253f
C406 B.t0 VSUBS 2.27548f
C407 B.n66 VSUBS 0.288768f
C408 B.n67 VSUBS 0.096918f
C409 B.n68 VSUBS 0.021092f
C410 B.n69 VSUBS 0.009104f
C411 B.n70 VSUBS 0.009104f
C412 B.n71 VSUBS 0.009104f
C413 B.n72 VSUBS 0.009104f
C414 B.n73 VSUBS 0.009104f
C415 B.n74 VSUBS 0.009104f
C416 B.n75 VSUBS 0.009104f
C417 B.n76 VSUBS 0.009104f
C418 B.n77 VSUBS 0.009104f
C419 B.n78 VSUBS 0.009104f
C420 B.n79 VSUBS 0.009104f
C421 B.n80 VSUBS 0.009104f
C422 B.n81 VSUBS 0.009104f
C423 B.n82 VSUBS 0.009104f
C424 B.n83 VSUBS 0.009104f
C425 B.n84 VSUBS 0.009104f
C426 B.n85 VSUBS 0.009104f
C427 B.n86 VSUBS 0.009104f
C428 B.n87 VSUBS 0.022244f
C429 B.n88 VSUBS 0.009104f
C430 B.n89 VSUBS 0.009104f
C431 B.n90 VSUBS 0.009104f
C432 B.n91 VSUBS 0.009104f
C433 B.n92 VSUBS 0.009104f
C434 B.n93 VSUBS 0.009104f
C435 B.n94 VSUBS 0.009104f
C436 B.n95 VSUBS 0.009104f
C437 B.n96 VSUBS 0.009104f
C438 B.n97 VSUBS 0.009104f
C439 B.n98 VSUBS 0.009104f
C440 B.n99 VSUBS 0.009104f
C441 B.n100 VSUBS 0.009104f
C442 B.n101 VSUBS 0.009104f
C443 B.n102 VSUBS 0.009104f
C444 B.n103 VSUBS 0.009104f
C445 B.n104 VSUBS 0.009104f
C446 B.n105 VSUBS 0.009104f
C447 B.n106 VSUBS 0.009104f
C448 B.n107 VSUBS 0.009104f
C449 B.n108 VSUBS 0.009104f
C450 B.n109 VSUBS 0.009104f
C451 B.n110 VSUBS 0.009104f
C452 B.n111 VSUBS 0.009104f
C453 B.n112 VSUBS 0.009104f
C454 B.n113 VSUBS 0.009104f
C455 B.n114 VSUBS 0.009104f
C456 B.n115 VSUBS 0.009104f
C457 B.n116 VSUBS 0.009104f
C458 B.n117 VSUBS 0.009104f
C459 B.n118 VSUBS 0.009104f
C460 B.n119 VSUBS 0.009104f
C461 B.n120 VSUBS 0.009104f
C462 B.n121 VSUBS 0.009104f
C463 B.n122 VSUBS 0.009104f
C464 B.n123 VSUBS 0.009104f
C465 B.n124 VSUBS 0.009104f
C466 B.n125 VSUBS 0.009104f
C467 B.n126 VSUBS 0.009104f
C468 B.n127 VSUBS 0.009104f
C469 B.n128 VSUBS 0.009104f
C470 B.n129 VSUBS 0.009104f
C471 B.n130 VSUBS 0.009104f
C472 B.n131 VSUBS 0.009104f
C473 B.n132 VSUBS 0.009104f
C474 B.n133 VSUBS 0.009104f
C475 B.n134 VSUBS 0.009104f
C476 B.n135 VSUBS 0.009104f
C477 B.n136 VSUBS 0.009104f
C478 B.n137 VSUBS 0.009104f
C479 B.n138 VSUBS 0.009104f
C480 B.n139 VSUBS 0.009104f
C481 B.n140 VSUBS 0.009104f
C482 B.n141 VSUBS 0.009104f
C483 B.n142 VSUBS 0.009104f
C484 B.n143 VSUBS 0.009104f
C485 B.n144 VSUBS 0.009104f
C486 B.n145 VSUBS 0.009104f
C487 B.n146 VSUBS 0.009104f
C488 B.n147 VSUBS 0.009104f
C489 B.n148 VSUBS 0.009104f
C490 B.n149 VSUBS 0.009104f
C491 B.n150 VSUBS 0.009104f
C492 B.n151 VSUBS 0.009104f
C493 B.n152 VSUBS 0.009104f
C494 B.n153 VSUBS 0.009104f
C495 B.n154 VSUBS 0.009104f
C496 B.n155 VSUBS 0.009104f
C497 B.n156 VSUBS 0.009104f
C498 B.n157 VSUBS 0.009104f
C499 B.n158 VSUBS 0.009104f
C500 B.n159 VSUBS 0.022695f
C501 B.n160 VSUBS 0.009104f
C502 B.n161 VSUBS 0.009104f
C503 B.n162 VSUBS 0.009104f
C504 B.n163 VSUBS 0.009104f
C505 B.n164 VSUBS 0.009104f
C506 B.n165 VSUBS 0.009104f
C507 B.n166 VSUBS 0.009104f
C508 B.n167 VSUBS 0.009104f
C509 B.n168 VSUBS 0.009104f
C510 B.n169 VSUBS 0.009104f
C511 B.n170 VSUBS 0.009104f
C512 B.n171 VSUBS 0.009104f
C513 B.n172 VSUBS 0.009104f
C514 B.n173 VSUBS 0.009104f
C515 B.n174 VSUBS 0.009104f
C516 B.n175 VSUBS 0.009104f
C517 B.n176 VSUBS 0.009104f
C518 B.n177 VSUBS 0.009104f
C519 B.n178 VSUBS 0.009104f
C520 B.n179 VSUBS 0.008568f
C521 B.n180 VSUBS 0.009104f
C522 B.n181 VSUBS 0.009104f
C523 B.n182 VSUBS 0.009104f
C524 B.n183 VSUBS 0.009104f
C525 B.n184 VSUBS 0.009104f
C526 B.t11 VSUBS 0.489322f
C527 B.t10 VSUBS 0.522261f
C528 B.t9 VSUBS 2.27548f
C529 B.n185 VSUBS 0.28876f
C530 B.n186 VSUBS 0.096909f
C531 B.n187 VSUBS 0.009104f
C532 B.n188 VSUBS 0.009104f
C533 B.n189 VSUBS 0.009104f
C534 B.n190 VSUBS 0.009104f
C535 B.n191 VSUBS 0.009104f
C536 B.n192 VSUBS 0.009104f
C537 B.n193 VSUBS 0.009104f
C538 B.n194 VSUBS 0.009104f
C539 B.n195 VSUBS 0.009104f
C540 B.n196 VSUBS 0.009104f
C541 B.n197 VSUBS 0.009104f
C542 B.n198 VSUBS 0.009104f
C543 B.n199 VSUBS 0.009104f
C544 B.n200 VSUBS 0.009104f
C545 B.n201 VSUBS 0.009104f
C546 B.n202 VSUBS 0.009104f
C547 B.n203 VSUBS 0.009104f
C548 B.n204 VSUBS 0.009104f
C549 B.n205 VSUBS 0.009104f
C550 B.n206 VSUBS 0.022244f
C551 B.n207 VSUBS 0.009104f
C552 B.n208 VSUBS 0.009104f
C553 B.n209 VSUBS 0.009104f
C554 B.n210 VSUBS 0.009104f
C555 B.n211 VSUBS 0.009104f
C556 B.n212 VSUBS 0.009104f
C557 B.n213 VSUBS 0.009104f
C558 B.n214 VSUBS 0.009104f
C559 B.n215 VSUBS 0.009104f
C560 B.n216 VSUBS 0.009104f
C561 B.n217 VSUBS 0.009104f
C562 B.n218 VSUBS 0.009104f
C563 B.n219 VSUBS 0.009104f
C564 B.n220 VSUBS 0.009104f
C565 B.n221 VSUBS 0.009104f
C566 B.n222 VSUBS 0.009104f
C567 B.n223 VSUBS 0.009104f
C568 B.n224 VSUBS 0.009104f
C569 B.n225 VSUBS 0.009104f
C570 B.n226 VSUBS 0.009104f
C571 B.n227 VSUBS 0.009104f
C572 B.n228 VSUBS 0.009104f
C573 B.n229 VSUBS 0.009104f
C574 B.n230 VSUBS 0.009104f
C575 B.n231 VSUBS 0.009104f
C576 B.n232 VSUBS 0.009104f
C577 B.n233 VSUBS 0.009104f
C578 B.n234 VSUBS 0.009104f
C579 B.n235 VSUBS 0.009104f
C580 B.n236 VSUBS 0.009104f
C581 B.n237 VSUBS 0.009104f
C582 B.n238 VSUBS 0.009104f
C583 B.n239 VSUBS 0.009104f
C584 B.n240 VSUBS 0.009104f
C585 B.n241 VSUBS 0.009104f
C586 B.n242 VSUBS 0.009104f
C587 B.n243 VSUBS 0.009104f
C588 B.n244 VSUBS 0.009104f
C589 B.n245 VSUBS 0.009104f
C590 B.n246 VSUBS 0.009104f
C591 B.n247 VSUBS 0.009104f
C592 B.n248 VSUBS 0.009104f
C593 B.n249 VSUBS 0.009104f
C594 B.n250 VSUBS 0.009104f
C595 B.n251 VSUBS 0.009104f
C596 B.n252 VSUBS 0.009104f
C597 B.n253 VSUBS 0.009104f
C598 B.n254 VSUBS 0.009104f
C599 B.n255 VSUBS 0.009104f
C600 B.n256 VSUBS 0.009104f
C601 B.n257 VSUBS 0.009104f
C602 B.n258 VSUBS 0.009104f
C603 B.n259 VSUBS 0.009104f
C604 B.n260 VSUBS 0.009104f
C605 B.n261 VSUBS 0.009104f
C606 B.n262 VSUBS 0.009104f
C607 B.n263 VSUBS 0.009104f
C608 B.n264 VSUBS 0.009104f
C609 B.n265 VSUBS 0.009104f
C610 B.n266 VSUBS 0.009104f
C611 B.n267 VSUBS 0.009104f
C612 B.n268 VSUBS 0.009104f
C613 B.n269 VSUBS 0.009104f
C614 B.n270 VSUBS 0.009104f
C615 B.n271 VSUBS 0.009104f
C616 B.n272 VSUBS 0.009104f
C617 B.n273 VSUBS 0.009104f
C618 B.n274 VSUBS 0.009104f
C619 B.n275 VSUBS 0.009104f
C620 B.n276 VSUBS 0.009104f
C621 B.n277 VSUBS 0.009104f
C622 B.n278 VSUBS 0.009104f
C623 B.n279 VSUBS 0.009104f
C624 B.n280 VSUBS 0.009104f
C625 B.n281 VSUBS 0.009104f
C626 B.n282 VSUBS 0.009104f
C627 B.n283 VSUBS 0.009104f
C628 B.n284 VSUBS 0.009104f
C629 B.n285 VSUBS 0.009104f
C630 B.n286 VSUBS 0.009104f
C631 B.n287 VSUBS 0.009104f
C632 B.n288 VSUBS 0.009104f
C633 B.n289 VSUBS 0.009104f
C634 B.n290 VSUBS 0.009104f
C635 B.n291 VSUBS 0.009104f
C636 B.n292 VSUBS 0.009104f
C637 B.n293 VSUBS 0.009104f
C638 B.n294 VSUBS 0.009104f
C639 B.n295 VSUBS 0.009104f
C640 B.n296 VSUBS 0.009104f
C641 B.n297 VSUBS 0.009104f
C642 B.n298 VSUBS 0.009104f
C643 B.n299 VSUBS 0.009104f
C644 B.n300 VSUBS 0.009104f
C645 B.n301 VSUBS 0.009104f
C646 B.n302 VSUBS 0.009104f
C647 B.n303 VSUBS 0.009104f
C648 B.n304 VSUBS 0.009104f
C649 B.n305 VSUBS 0.009104f
C650 B.n306 VSUBS 0.009104f
C651 B.n307 VSUBS 0.009104f
C652 B.n308 VSUBS 0.009104f
C653 B.n309 VSUBS 0.009104f
C654 B.n310 VSUBS 0.009104f
C655 B.n311 VSUBS 0.009104f
C656 B.n312 VSUBS 0.009104f
C657 B.n313 VSUBS 0.009104f
C658 B.n314 VSUBS 0.009104f
C659 B.n315 VSUBS 0.009104f
C660 B.n316 VSUBS 0.009104f
C661 B.n317 VSUBS 0.009104f
C662 B.n318 VSUBS 0.009104f
C663 B.n319 VSUBS 0.009104f
C664 B.n320 VSUBS 0.009104f
C665 B.n321 VSUBS 0.009104f
C666 B.n322 VSUBS 0.009104f
C667 B.n323 VSUBS 0.009104f
C668 B.n324 VSUBS 0.009104f
C669 B.n325 VSUBS 0.009104f
C670 B.n326 VSUBS 0.009104f
C671 B.n327 VSUBS 0.009104f
C672 B.n328 VSUBS 0.009104f
C673 B.n329 VSUBS 0.009104f
C674 B.n330 VSUBS 0.009104f
C675 B.n331 VSUBS 0.009104f
C676 B.n332 VSUBS 0.009104f
C677 B.n333 VSUBS 0.009104f
C678 B.n334 VSUBS 0.009104f
C679 B.n335 VSUBS 0.009104f
C680 B.n336 VSUBS 0.009104f
C681 B.n337 VSUBS 0.009104f
C682 B.n338 VSUBS 0.009104f
C683 B.n339 VSUBS 0.009104f
C684 B.n340 VSUBS 0.009104f
C685 B.n341 VSUBS 0.009104f
C686 B.n342 VSUBS 0.009104f
C687 B.n343 VSUBS 0.009104f
C688 B.n344 VSUBS 0.009104f
C689 B.n345 VSUBS 0.021667f
C690 B.n346 VSUBS 0.021667f
C691 B.n347 VSUBS 0.022244f
C692 B.n348 VSUBS 0.009104f
C693 B.n349 VSUBS 0.009104f
C694 B.n350 VSUBS 0.009104f
C695 B.n351 VSUBS 0.009104f
C696 B.n352 VSUBS 0.009104f
C697 B.n353 VSUBS 0.009104f
C698 B.n354 VSUBS 0.009104f
C699 B.n355 VSUBS 0.009104f
C700 B.n356 VSUBS 0.009104f
C701 B.n357 VSUBS 0.009104f
C702 B.n358 VSUBS 0.009104f
C703 B.n359 VSUBS 0.009104f
C704 B.n360 VSUBS 0.009104f
C705 B.n361 VSUBS 0.009104f
C706 B.n362 VSUBS 0.009104f
C707 B.n363 VSUBS 0.009104f
C708 B.n364 VSUBS 0.009104f
C709 B.n365 VSUBS 0.009104f
C710 B.n366 VSUBS 0.009104f
C711 B.n367 VSUBS 0.009104f
C712 B.n368 VSUBS 0.009104f
C713 B.n369 VSUBS 0.009104f
C714 B.n370 VSUBS 0.009104f
C715 B.n371 VSUBS 0.009104f
C716 B.n372 VSUBS 0.009104f
C717 B.n373 VSUBS 0.009104f
C718 B.n374 VSUBS 0.009104f
C719 B.n375 VSUBS 0.009104f
C720 B.n376 VSUBS 0.009104f
C721 B.n377 VSUBS 0.009104f
C722 B.n378 VSUBS 0.009104f
C723 B.n379 VSUBS 0.009104f
C724 B.n380 VSUBS 0.009104f
C725 B.n381 VSUBS 0.009104f
C726 B.n382 VSUBS 0.009104f
C727 B.n383 VSUBS 0.009104f
C728 B.n384 VSUBS 0.009104f
C729 B.n385 VSUBS 0.009104f
C730 B.n386 VSUBS 0.009104f
C731 B.n387 VSUBS 0.009104f
C732 B.n388 VSUBS 0.009104f
C733 B.n389 VSUBS 0.009104f
C734 B.n390 VSUBS 0.009104f
C735 B.n391 VSUBS 0.009104f
C736 B.n392 VSUBS 0.009104f
C737 B.n393 VSUBS 0.009104f
C738 B.n394 VSUBS 0.009104f
C739 B.n395 VSUBS 0.009104f
C740 B.n396 VSUBS 0.009104f
C741 B.n397 VSUBS 0.009104f
C742 B.n398 VSUBS 0.009104f
C743 B.n399 VSUBS 0.009104f
C744 B.n400 VSUBS 0.009104f
C745 B.n401 VSUBS 0.009104f
C746 B.n402 VSUBS 0.009104f
C747 B.n403 VSUBS 0.009104f
C748 B.n404 VSUBS 0.009104f
C749 B.n405 VSUBS 0.009104f
C750 B.n406 VSUBS 0.008568f
C751 B.n407 VSUBS 0.021092f
C752 B.n408 VSUBS 0.005087f
C753 B.n409 VSUBS 0.009104f
C754 B.n410 VSUBS 0.009104f
C755 B.n411 VSUBS 0.009104f
C756 B.n412 VSUBS 0.009104f
C757 B.n413 VSUBS 0.009104f
C758 B.n414 VSUBS 0.009104f
C759 B.n415 VSUBS 0.009104f
C760 B.n416 VSUBS 0.009104f
C761 B.n417 VSUBS 0.009104f
C762 B.n418 VSUBS 0.009104f
C763 B.n419 VSUBS 0.009104f
C764 B.n420 VSUBS 0.009104f
C765 B.t5 VSUBS 0.489313f
C766 B.t4 VSUBS 0.522253f
C767 B.t3 VSUBS 2.27548f
C768 B.n421 VSUBS 0.288768f
C769 B.n422 VSUBS 0.096918f
C770 B.n423 VSUBS 0.021092f
C771 B.n424 VSUBS 0.005087f
C772 B.n425 VSUBS 0.009104f
C773 B.n426 VSUBS 0.009104f
C774 B.n427 VSUBS 0.009104f
C775 B.n428 VSUBS 0.009104f
C776 B.n429 VSUBS 0.009104f
C777 B.n430 VSUBS 0.009104f
C778 B.n431 VSUBS 0.009104f
C779 B.n432 VSUBS 0.009104f
C780 B.n433 VSUBS 0.009104f
C781 B.n434 VSUBS 0.009104f
C782 B.n435 VSUBS 0.009104f
C783 B.n436 VSUBS 0.009104f
C784 B.n437 VSUBS 0.009104f
C785 B.n438 VSUBS 0.009104f
C786 B.n439 VSUBS 0.009104f
C787 B.n440 VSUBS 0.009104f
C788 B.n441 VSUBS 0.009104f
C789 B.n442 VSUBS 0.009104f
C790 B.n443 VSUBS 0.009104f
C791 B.n444 VSUBS 0.009104f
C792 B.n445 VSUBS 0.009104f
C793 B.n446 VSUBS 0.009104f
C794 B.n447 VSUBS 0.009104f
C795 B.n448 VSUBS 0.009104f
C796 B.n449 VSUBS 0.009104f
C797 B.n450 VSUBS 0.009104f
C798 B.n451 VSUBS 0.009104f
C799 B.n452 VSUBS 0.009104f
C800 B.n453 VSUBS 0.009104f
C801 B.n454 VSUBS 0.009104f
C802 B.n455 VSUBS 0.009104f
C803 B.n456 VSUBS 0.009104f
C804 B.n457 VSUBS 0.009104f
C805 B.n458 VSUBS 0.009104f
C806 B.n459 VSUBS 0.009104f
C807 B.n460 VSUBS 0.009104f
C808 B.n461 VSUBS 0.009104f
C809 B.n462 VSUBS 0.009104f
C810 B.n463 VSUBS 0.009104f
C811 B.n464 VSUBS 0.009104f
C812 B.n465 VSUBS 0.009104f
C813 B.n466 VSUBS 0.009104f
C814 B.n467 VSUBS 0.009104f
C815 B.n468 VSUBS 0.009104f
C816 B.n469 VSUBS 0.009104f
C817 B.n470 VSUBS 0.009104f
C818 B.n471 VSUBS 0.009104f
C819 B.n472 VSUBS 0.009104f
C820 B.n473 VSUBS 0.009104f
C821 B.n474 VSUBS 0.009104f
C822 B.n475 VSUBS 0.009104f
C823 B.n476 VSUBS 0.009104f
C824 B.n477 VSUBS 0.009104f
C825 B.n478 VSUBS 0.009104f
C826 B.n479 VSUBS 0.009104f
C827 B.n480 VSUBS 0.009104f
C828 B.n481 VSUBS 0.009104f
C829 B.n482 VSUBS 0.009104f
C830 B.n483 VSUBS 0.009104f
C831 B.n484 VSUBS 0.021216f
C832 B.n485 VSUBS 0.022244f
C833 B.n486 VSUBS 0.021667f
C834 B.n487 VSUBS 0.009104f
C835 B.n488 VSUBS 0.009104f
C836 B.n489 VSUBS 0.009104f
C837 B.n490 VSUBS 0.009104f
C838 B.n491 VSUBS 0.009104f
C839 B.n492 VSUBS 0.009104f
C840 B.n493 VSUBS 0.009104f
C841 B.n494 VSUBS 0.009104f
C842 B.n495 VSUBS 0.009104f
C843 B.n496 VSUBS 0.009104f
C844 B.n497 VSUBS 0.009104f
C845 B.n498 VSUBS 0.009104f
C846 B.n499 VSUBS 0.009104f
C847 B.n500 VSUBS 0.009104f
C848 B.n501 VSUBS 0.009104f
C849 B.n502 VSUBS 0.009104f
C850 B.n503 VSUBS 0.009104f
C851 B.n504 VSUBS 0.009104f
C852 B.n505 VSUBS 0.009104f
C853 B.n506 VSUBS 0.009104f
C854 B.n507 VSUBS 0.009104f
C855 B.n508 VSUBS 0.009104f
C856 B.n509 VSUBS 0.009104f
C857 B.n510 VSUBS 0.009104f
C858 B.n511 VSUBS 0.009104f
C859 B.n512 VSUBS 0.009104f
C860 B.n513 VSUBS 0.009104f
C861 B.n514 VSUBS 0.009104f
C862 B.n515 VSUBS 0.009104f
C863 B.n516 VSUBS 0.009104f
C864 B.n517 VSUBS 0.009104f
C865 B.n518 VSUBS 0.009104f
C866 B.n519 VSUBS 0.009104f
C867 B.n520 VSUBS 0.009104f
C868 B.n521 VSUBS 0.009104f
C869 B.n522 VSUBS 0.009104f
C870 B.n523 VSUBS 0.009104f
C871 B.n524 VSUBS 0.009104f
C872 B.n525 VSUBS 0.009104f
C873 B.n526 VSUBS 0.009104f
C874 B.n527 VSUBS 0.009104f
C875 B.n528 VSUBS 0.009104f
C876 B.n529 VSUBS 0.009104f
C877 B.n530 VSUBS 0.009104f
C878 B.n531 VSUBS 0.009104f
C879 B.n532 VSUBS 0.009104f
C880 B.n533 VSUBS 0.009104f
C881 B.n534 VSUBS 0.009104f
C882 B.n535 VSUBS 0.009104f
C883 B.n536 VSUBS 0.009104f
C884 B.n537 VSUBS 0.009104f
C885 B.n538 VSUBS 0.009104f
C886 B.n539 VSUBS 0.009104f
C887 B.n540 VSUBS 0.009104f
C888 B.n541 VSUBS 0.009104f
C889 B.n542 VSUBS 0.009104f
C890 B.n543 VSUBS 0.009104f
C891 B.n544 VSUBS 0.009104f
C892 B.n545 VSUBS 0.009104f
C893 B.n546 VSUBS 0.009104f
C894 B.n547 VSUBS 0.009104f
C895 B.n548 VSUBS 0.009104f
C896 B.n549 VSUBS 0.009104f
C897 B.n550 VSUBS 0.009104f
C898 B.n551 VSUBS 0.009104f
C899 B.n552 VSUBS 0.009104f
C900 B.n553 VSUBS 0.009104f
C901 B.n554 VSUBS 0.009104f
C902 B.n555 VSUBS 0.009104f
C903 B.n556 VSUBS 0.009104f
C904 B.n557 VSUBS 0.009104f
C905 B.n558 VSUBS 0.009104f
C906 B.n559 VSUBS 0.009104f
C907 B.n560 VSUBS 0.009104f
C908 B.n561 VSUBS 0.009104f
C909 B.n562 VSUBS 0.009104f
C910 B.n563 VSUBS 0.009104f
C911 B.n564 VSUBS 0.009104f
C912 B.n565 VSUBS 0.009104f
C913 B.n566 VSUBS 0.009104f
C914 B.n567 VSUBS 0.009104f
C915 B.n568 VSUBS 0.009104f
C916 B.n569 VSUBS 0.009104f
C917 B.n570 VSUBS 0.009104f
C918 B.n571 VSUBS 0.009104f
C919 B.n572 VSUBS 0.009104f
C920 B.n573 VSUBS 0.009104f
C921 B.n574 VSUBS 0.009104f
C922 B.n575 VSUBS 0.009104f
C923 B.n576 VSUBS 0.009104f
C924 B.n577 VSUBS 0.009104f
C925 B.n578 VSUBS 0.009104f
C926 B.n579 VSUBS 0.009104f
C927 B.n580 VSUBS 0.009104f
C928 B.n581 VSUBS 0.009104f
C929 B.n582 VSUBS 0.009104f
C930 B.n583 VSUBS 0.009104f
C931 B.n584 VSUBS 0.009104f
C932 B.n585 VSUBS 0.009104f
C933 B.n586 VSUBS 0.009104f
C934 B.n587 VSUBS 0.009104f
C935 B.n588 VSUBS 0.009104f
C936 B.n589 VSUBS 0.009104f
C937 B.n590 VSUBS 0.009104f
C938 B.n591 VSUBS 0.009104f
C939 B.n592 VSUBS 0.009104f
C940 B.n593 VSUBS 0.009104f
C941 B.n594 VSUBS 0.009104f
C942 B.n595 VSUBS 0.009104f
C943 B.n596 VSUBS 0.009104f
C944 B.n597 VSUBS 0.009104f
C945 B.n598 VSUBS 0.009104f
C946 B.n599 VSUBS 0.009104f
C947 B.n600 VSUBS 0.009104f
C948 B.n601 VSUBS 0.009104f
C949 B.n602 VSUBS 0.009104f
C950 B.n603 VSUBS 0.009104f
C951 B.n604 VSUBS 0.009104f
C952 B.n605 VSUBS 0.009104f
C953 B.n606 VSUBS 0.009104f
C954 B.n607 VSUBS 0.009104f
C955 B.n608 VSUBS 0.009104f
C956 B.n609 VSUBS 0.009104f
C957 B.n610 VSUBS 0.009104f
C958 B.n611 VSUBS 0.009104f
C959 B.n612 VSUBS 0.009104f
C960 B.n613 VSUBS 0.009104f
C961 B.n614 VSUBS 0.009104f
C962 B.n615 VSUBS 0.009104f
C963 B.n616 VSUBS 0.009104f
C964 B.n617 VSUBS 0.009104f
C965 B.n618 VSUBS 0.009104f
C966 B.n619 VSUBS 0.009104f
C967 B.n620 VSUBS 0.009104f
C968 B.n621 VSUBS 0.009104f
C969 B.n622 VSUBS 0.009104f
C970 B.n623 VSUBS 0.009104f
C971 B.n624 VSUBS 0.009104f
C972 B.n625 VSUBS 0.009104f
C973 B.n626 VSUBS 0.009104f
C974 B.n627 VSUBS 0.009104f
C975 B.n628 VSUBS 0.009104f
C976 B.n629 VSUBS 0.009104f
C977 B.n630 VSUBS 0.009104f
C978 B.n631 VSUBS 0.009104f
C979 B.n632 VSUBS 0.009104f
C980 B.n633 VSUBS 0.009104f
C981 B.n634 VSUBS 0.009104f
C982 B.n635 VSUBS 0.009104f
C983 B.n636 VSUBS 0.009104f
C984 B.n637 VSUBS 0.009104f
C985 B.n638 VSUBS 0.009104f
C986 B.n639 VSUBS 0.009104f
C987 B.n640 VSUBS 0.009104f
C988 B.n641 VSUBS 0.009104f
C989 B.n642 VSUBS 0.009104f
C990 B.n643 VSUBS 0.009104f
C991 B.n644 VSUBS 0.009104f
C992 B.n645 VSUBS 0.009104f
C993 B.n646 VSUBS 0.009104f
C994 B.n647 VSUBS 0.009104f
C995 B.n648 VSUBS 0.009104f
C996 B.n649 VSUBS 0.009104f
C997 B.n650 VSUBS 0.009104f
C998 B.n651 VSUBS 0.009104f
C999 B.n652 VSUBS 0.009104f
C1000 B.n653 VSUBS 0.009104f
C1001 B.n654 VSUBS 0.009104f
C1002 B.n655 VSUBS 0.009104f
C1003 B.n656 VSUBS 0.009104f
C1004 B.n657 VSUBS 0.009104f
C1005 B.n658 VSUBS 0.009104f
C1006 B.n659 VSUBS 0.009104f
C1007 B.n660 VSUBS 0.009104f
C1008 B.n661 VSUBS 0.009104f
C1009 B.n662 VSUBS 0.009104f
C1010 B.n663 VSUBS 0.009104f
C1011 B.n664 VSUBS 0.009104f
C1012 B.n665 VSUBS 0.009104f
C1013 B.n666 VSUBS 0.009104f
C1014 B.n667 VSUBS 0.009104f
C1015 B.n668 VSUBS 0.009104f
C1016 B.n669 VSUBS 0.009104f
C1017 B.n670 VSUBS 0.009104f
C1018 B.n671 VSUBS 0.009104f
C1019 B.n672 VSUBS 0.009104f
C1020 B.n673 VSUBS 0.009104f
C1021 B.n674 VSUBS 0.009104f
C1022 B.n675 VSUBS 0.009104f
C1023 B.n676 VSUBS 0.009104f
C1024 B.n677 VSUBS 0.009104f
C1025 B.n678 VSUBS 0.009104f
C1026 B.n679 VSUBS 0.009104f
C1027 B.n680 VSUBS 0.009104f
C1028 B.n681 VSUBS 0.009104f
C1029 B.n682 VSUBS 0.009104f
C1030 B.n683 VSUBS 0.009104f
C1031 B.n684 VSUBS 0.009104f
C1032 B.n685 VSUBS 0.009104f
C1033 B.n686 VSUBS 0.009104f
C1034 B.n687 VSUBS 0.009104f
C1035 B.n688 VSUBS 0.009104f
C1036 B.n689 VSUBS 0.009104f
C1037 B.n690 VSUBS 0.009104f
C1038 B.n691 VSUBS 0.009104f
C1039 B.n692 VSUBS 0.009104f
C1040 B.n693 VSUBS 0.009104f
C1041 B.n694 VSUBS 0.009104f
C1042 B.n695 VSUBS 0.009104f
C1043 B.n696 VSUBS 0.009104f
C1044 B.n697 VSUBS 0.009104f
C1045 B.n698 VSUBS 0.009104f
C1046 B.n699 VSUBS 0.009104f
C1047 B.n700 VSUBS 0.021667f
C1048 B.n701 VSUBS 0.021667f
C1049 B.n702 VSUBS 0.022244f
C1050 B.n703 VSUBS 0.009104f
C1051 B.n704 VSUBS 0.009104f
C1052 B.n705 VSUBS 0.009104f
C1053 B.n706 VSUBS 0.009104f
C1054 B.n707 VSUBS 0.009104f
C1055 B.n708 VSUBS 0.009104f
C1056 B.n709 VSUBS 0.009104f
C1057 B.n710 VSUBS 0.009104f
C1058 B.n711 VSUBS 0.009104f
C1059 B.n712 VSUBS 0.009104f
C1060 B.n713 VSUBS 0.009104f
C1061 B.n714 VSUBS 0.009104f
C1062 B.n715 VSUBS 0.009104f
C1063 B.n716 VSUBS 0.009104f
C1064 B.n717 VSUBS 0.009104f
C1065 B.n718 VSUBS 0.009104f
C1066 B.n719 VSUBS 0.009104f
C1067 B.n720 VSUBS 0.009104f
C1068 B.n721 VSUBS 0.009104f
C1069 B.n722 VSUBS 0.009104f
C1070 B.n723 VSUBS 0.009104f
C1071 B.n724 VSUBS 0.009104f
C1072 B.n725 VSUBS 0.009104f
C1073 B.n726 VSUBS 0.009104f
C1074 B.n727 VSUBS 0.009104f
C1075 B.n728 VSUBS 0.009104f
C1076 B.n729 VSUBS 0.009104f
C1077 B.n730 VSUBS 0.009104f
C1078 B.n731 VSUBS 0.009104f
C1079 B.n732 VSUBS 0.009104f
C1080 B.n733 VSUBS 0.009104f
C1081 B.n734 VSUBS 0.009104f
C1082 B.n735 VSUBS 0.009104f
C1083 B.n736 VSUBS 0.009104f
C1084 B.n737 VSUBS 0.009104f
C1085 B.n738 VSUBS 0.009104f
C1086 B.n739 VSUBS 0.009104f
C1087 B.n740 VSUBS 0.009104f
C1088 B.n741 VSUBS 0.009104f
C1089 B.n742 VSUBS 0.009104f
C1090 B.n743 VSUBS 0.009104f
C1091 B.n744 VSUBS 0.009104f
C1092 B.n745 VSUBS 0.009104f
C1093 B.n746 VSUBS 0.009104f
C1094 B.n747 VSUBS 0.009104f
C1095 B.n748 VSUBS 0.009104f
C1096 B.n749 VSUBS 0.009104f
C1097 B.n750 VSUBS 0.009104f
C1098 B.n751 VSUBS 0.009104f
C1099 B.n752 VSUBS 0.009104f
C1100 B.n753 VSUBS 0.009104f
C1101 B.n754 VSUBS 0.009104f
C1102 B.n755 VSUBS 0.009104f
C1103 B.n756 VSUBS 0.009104f
C1104 B.n757 VSUBS 0.009104f
C1105 B.n758 VSUBS 0.009104f
C1106 B.n759 VSUBS 0.009104f
C1107 B.n760 VSUBS 0.008568f
C1108 B.n761 VSUBS 0.009104f
C1109 B.n762 VSUBS 0.009104f
C1110 B.n763 VSUBS 0.009104f
C1111 B.n764 VSUBS 0.009104f
C1112 B.n765 VSUBS 0.009104f
C1113 B.n766 VSUBS 0.009104f
C1114 B.n767 VSUBS 0.009104f
C1115 B.n768 VSUBS 0.009104f
C1116 B.n769 VSUBS 0.009104f
C1117 B.n770 VSUBS 0.009104f
C1118 B.n771 VSUBS 0.009104f
C1119 B.n772 VSUBS 0.009104f
C1120 B.n773 VSUBS 0.009104f
C1121 B.n774 VSUBS 0.009104f
C1122 B.n775 VSUBS 0.009104f
C1123 B.n776 VSUBS 0.005087f
C1124 B.n777 VSUBS 0.021092f
C1125 B.n778 VSUBS 0.008568f
C1126 B.n779 VSUBS 0.009104f
C1127 B.n780 VSUBS 0.009104f
C1128 B.n781 VSUBS 0.009104f
C1129 B.n782 VSUBS 0.009104f
C1130 B.n783 VSUBS 0.009104f
C1131 B.n784 VSUBS 0.009104f
C1132 B.n785 VSUBS 0.009104f
C1133 B.n786 VSUBS 0.009104f
C1134 B.n787 VSUBS 0.009104f
C1135 B.n788 VSUBS 0.009104f
C1136 B.n789 VSUBS 0.009104f
C1137 B.n790 VSUBS 0.009104f
C1138 B.n791 VSUBS 0.009104f
C1139 B.n792 VSUBS 0.009104f
C1140 B.n793 VSUBS 0.009104f
C1141 B.n794 VSUBS 0.009104f
C1142 B.n795 VSUBS 0.009104f
C1143 B.n796 VSUBS 0.009104f
C1144 B.n797 VSUBS 0.009104f
C1145 B.n798 VSUBS 0.009104f
C1146 B.n799 VSUBS 0.009104f
C1147 B.n800 VSUBS 0.009104f
C1148 B.n801 VSUBS 0.009104f
C1149 B.n802 VSUBS 0.009104f
C1150 B.n803 VSUBS 0.009104f
C1151 B.n804 VSUBS 0.009104f
C1152 B.n805 VSUBS 0.009104f
C1153 B.n806 VSUBS 0.009104f
C1154 B.n807 VSUBS 0.009104f
C1155 B.n808 VSUBS 0.009104f
C1156 B.n809 VSUBS 0.009104f
C1157 B.n810 VSUBS 0.009104f
C1158 B.n811 VSUBS 0.009104f
C1159 B.n812 VSUBS 0.009104f
C1160 B.n813 VSUBS 0.009104f
C1161 B.n814 VSUBS 0.009104f
C1162 B.n815 VSUBS 0.009104f
C1163 B.n816 VSUBS 0.009104f
C1164 B.n817 VSUBS 0.009104f
C1165 B.n818 VSUBS 0.009104f
C1166 B.n819 VSUBS 0.009104f
C1167 B.n820 VSUBS 0.009104f
C1168 B.n821 VSUBS 0.009104f
C1169 B.n822 VSUBS 0.009104f
C1170 B.n823 VSUBS 0.009104f
C1171 B.n824 VSUBS 0.009104f
C1172 B.n825 VSUBS 0.009104f
C1173 B.n826 VSUBS 0.009104f
C1174 B.n827 VSUBS 0.009104f
C1175 B.n828 VSUBS 0.009104f
C1176 B.n829 VSUBS 0.009104f
C1177 B.n830 VSUBS 0.009104f
C1178 B.n831 VSUBS 0.009104f
C1179 B.n832 VSUBS 0.009104f
C1180 B.n833 VSUBS 0.009104f
C1181 B.n834 VSUBS 0.009104f
C1182 B.n835 VSUBS 0.009104f
C1183 B.n836 VSUBS 0.022244f
C1184 B.n837 VSUBS 0.022244f
C1185 B.n838 VSUBS 0.021667f
C1186 B.n839 VSUBS 0.009104f
C1187 B.n840 VSUBS 0.009104f
C1188 B.n841 VSUBS 0.009104f
C1189 B.n842 VSUBS 0.009104f
C1190 B.n843 VSUBS 0.009104f
C1191 B.n844 VSUBS 0.009104f
C1192 B.n845 VSUBS 0.009104f
C1193 B.n846 VSUBS 0.009104f
C1194 B.n847 VSUBS 0.009104f
C1195 B.n848 VSUBS 0.009104f
C1196 B.n849 VSUBS 0.009104f
C1197 B.n850 VSUBS 0.009104f
C1198 B.n851 VSUBS 0.009104f
C1199 B.n852 VSUBS 0.009104f
C1200 B.n853 VSUBS 0.009104f
C1201 B.n854 VSUBS 0.009104f
C1202 B.n855 VSUBS 0.009104f
C1203 B.n856 VSUBS 0.009104f
C1204 B.n857 VSUBS 0.009104f
C1205 B.n858 VSUBS 0.009104f
C1206 B.n859 VSUBS 0.009104f
C1207 B.n860 VSUBS 0.009104f
C1208 B.n861 VSUBS 0.009104f
C1209 B.n862 VSUBS 0.009104f
C1210 B.n863 VSUBS 0.009104f
C1211 B.n864 VSUBS 0.009104f
C1212 B.n865 VSUBS 0.009104f
C1213 B.n866 VSUBS 0.009104f
C1214 B.n867 VSUBS 0.009104f
C1215 B.n868 VSUBS 0.009104f
C1216 B.n869 VSUBS 0.009104f
C1217 B.n870 VSUBS 0.009104f
C1218 B.n871 VSUBS 0.009104f
C1219 B.n872 VSUBS 0.009104f
C1220 B.n873 VSUBS 0.009104f
C1221 B.n874 VSUBS 0.009104f
C1222 B.n875 VSUBS 0.009104f
C1223 B.n876 VSUBS 0.009104f
C1224 B.n877 VSUBS 0.009104f
C1225 B.n878 VSUBS 0.009104f
C1226 B.n879 VSUBS 0.009104f
C1227 B.n880 VSUBS 0.009104f
C1228 B.n881 VSUBS 0.009104f
C1229 B.n882 VSUBS 0.009104f
C1230 B.n883 VSUBS 0.009104f
C1231 B.n884 VSUBS 0.009104f
C1232 B.n885 VSUBS 0.009104f
C1233 B.n886 VSUBS 0.009104f
C1234 B.n887 VSUBS 0.009104f
C1235 B.n888 VSUBS 0.009104f
C1236 B.n889 VSUBS 0.009104f
C1237 B.n890 VSUBS 0.009104f
C1238 B.n891 VSUBS 0.009104f
C1239 B.n892 VSUBS 0.009104f
C1240 B.n893 VSUBS 0.009104f
C1241 B.n894 VSUBS 0.009104f
C1242 B.n895 VSUBS 0.009104f
C1243 B.n896 VSUBS 0.009104f
C1244 B.n897 VSUBS 0.009104f
C1245 B.n898 VSUBS 0.009104f
C1246 B.n899 VSUBS 0.009104f
C1247 B.n900 VSUBS 0.009104f
C1248 B.n901 VSUBS 0.009104f
C1249 B.n902 VSUBS 0.009104f
C1250 B.n903 VSUBS 0.009104f
C1251 B.n904 VSUBS 0.009104f
C1252 B.n905 VSUBS 0.009104f
C1253 B.n906 VSUBS 0.009104f
C1254 B.n907 VSUBS 0.009104f
C1255 B.n908 VSUBS 0.009104f
C1256 B.n909 VSUBS 0.009104f
C1257 B.n910 VSUBS 0.009104f
C1258 B.n911 VSUBS 0.009104f
C1259 B.n912 VSUBS 0.009104f
C1260 B.n913 VSUBS 0.009104f
C1261 B.n914 VSUBS 0.009104f
C1262 B.n915 VSUBS 0.009104f
C1263 B.n916 VSUBS 0.009104f
C1264 B.n917 VSUBS 0.009104f
C1265 B.n918 VSUBS 0.009104f
C1266 B.n919 VSUBS 0.009104f
C1267 B.n920 VSUBS 0.009104f
C1268 B.n921 VSUBS 0.009104f
C1269 B.n922 VSUBS 0.009104f
C1270 B.n923 VSUBS 0.009104f
C1271 B.n924 VSUBS 0.009104f
C1272 B.n925 VSUBS 0.009104f
C1273 B.n926 VSUBS 0.009104f
C1274 B.n927 VSUBS 0.009104f
C1275 B.n928 VSUBS 0.009104f
C1276 B.n929 VSUBS 0.009104f
C1277 B.n930 VSUBS 0.009104f
C1278 B.n931 VSUBS 0.009104f
C1279 B.n932 VSUBS 0.009104f
C1280 B.n933 VSUBS 0.009104f
C1281 B.n934 VSUBS 0.009104f
C1282 B.n935 VSUBS 0.009104f
C1283 B.n936 VSUBS 0.009104f
C1284 B.n937 VSUBS 0.009104f
C1285 B.n938 VSUBS 0.009104f
C1286 B.n939 VSUBS 0.009104f
C1287 B.n940 VSUBS 0.009104f
C1288 B.n941 VSUBS 0.009104f
C1289 B.n942 VSUBS 0.009104f
C1290 B.n943 VSUBS 0.01188f
C1291 B.n944 VSUBS 0.012655f
C1292 B.n945 VSUBS 0.025165f
.ends

