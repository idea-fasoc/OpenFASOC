* NGSPICE file created from diff_pair_sample_1497.ext - technology: sky130A

.subckt diff_pair_sample_1497 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X1 VTAIL.t14 VP.t1 VDD1.t0 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X2 VTAIL.t16 VN.t0 VDD2.t9 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X3 VDD1.t3 VP.t2 VTAIL.t13 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=0.34
X4 VDD1.t7 VP.t3 VTAIL.t12 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=0.34
X5 VTAIL.t11 VP.t4 VDD1.t8 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X6 VDD1.t4 VP.t5 VTAIL.t10 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X7 VDD1.t9 VP.t6 VTAIL.t9 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=0.34
X8 VDD2.t8 VN.t1 VTAIL.t17 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=0.34
X9 B.t11 B.t9 B.t10 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=0.34
X10 VDD2.t7 VN.t2 VTAIL.t18 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=0.34
X11 VDD1.t6 VP.t7 VTAIL.t8 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=0.34
X12 B.t8 B.t6 B.t7 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=0.34
X13 VDD2.t6 VN.t3 VTAIL.t0 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X14 VTAIL.t19 VN.t4 VDD2.t5 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X15 VTAIL.t7 VP.t8 VDD1.t1 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X16 VTAIL.t3 VN.t5 VDD2.t4 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X17 VDD2.t3 VN.t6 VTAIL.t1 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=0.34
X18 VTAIL.t2 VN.t7 VDD2.t2 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X19 VDD1.t2 VP.t9 VTAIL.t6 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
X20 B.t5 B.t3 B.t4 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=0.34
X21 VDD2.t1 VN.t8 VTAIL.t5 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=0.34
X22 B.t2 B.t0 B.t1 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=0.34
X23 VDD2.t0 VN.t9 VTAIL.t4 w_n1774_n2726# sky130_fd_pr__pfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=0.34
R0 VP.n4 VP.t7 775.037
R1 VP.n16 VP.t2 764.134
R2 VP.n10 VP.t3 764.134
R3 VP.n8 VP.t6 764.134
R4 VP.n1 VP.t4 739.303
R5 VP.n14 VP.t5 739.303
R6 VP.n15 VP.t0 739.303
R7 VP.n7 VP.t8 739.303
R8 VP.n6 VP.t9 739.303
R9 VP.n5 VP.t1 739.303
R10 VP.n17 VP.n16 161.3
R11 VP.n6 VP.n3 161.3
R12 VP.n7 VP.n2 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n15 VP.n0 161.3
R15 VP.n14 VP.n13 161.3
R16 VP.n12 VP.n1 161.3
R17 VP.n11 VP.n10 161.3
R18 VP.n4 VP.n3 75.4397
R19 VP.n14 VP.n1 48.2005
R20 VP.n15 VP.n14 48.2005
R21 VP.n7 VP.n6 48.2005
R22 VP.n6 VP.n5 48.2005
R23 VP.n11 VP.n9 38.5194
R24 VP.n10 VP.n1 23.3702
R25 VP.n16 VP.n15 23.3702
R26 VP.n8 VP.n7 23.3702
R27 VP.n5 VP.n4 10.8906
R28 VP.n3 VP.n2 0.189894
R29 VP.n9 VP.n2 0.189894
R30 VP.n12 VP.n11 0.189894
R31 VP.n13 VP.n12 0.189894
R32 VP.n13 VP.n0 0.189894
R33 VP.n17 VP.n0 0.189894
R34 VP VP.n17 0.0516364
R35 VDD1.n42 VDD1.n0 756.745
R36 VDD1.n91 VDD1.n49 756.745
R37 VDD1.n43 VDD1.n42 585
R38 VDD1.n41 VDD1.n40 585
R39 VDD1.n4 VDD1.n3 585
R40 VDD1.n35 VDD1.n34 585
R41 VDD1.n33 VDD1.n32 585
R42 VDD1.n8 VDD1.n7 585
R43 VDD1.n27 VDD1.n26 585
R44 VDD1.n25 VDD1.n24 585
R45 VDD1.n12 VDD1.n11 585
R46 VDD1.n19 VDD1.n18 585
R47 VDD1.n17 VDD1.n16 585
R48 VDD1.n66 VDD1.n65 585
R49 VDD1.n68 VDD1.n67 585
R50 VDD1.n61 VDD1.n60 585
R51 VDD1.n74 VDD1.n73 585
R52 VDD1.n76 VDD1.n75 585
R53 VDD1.n57 VDD1.n56 585
R54 VDD1.n82 VDD1.n81 585
R55 VDD1.n84 VDD1.n83 585
R56 VDD1.n53 VDD1.n52 585
R57 VDD1.n90 VDD1.n89 585
R58 VDD1.n92 VDD1.n91 585
R59 VDD1.n15 VDD1.t6 327.469
R60 VDD1.n64 VDD1.t7 327.469
R61 VDD1.n42 VDD1.n41 171.744
R62 VDD1.n41 VDD1.n3 171.744
R63 VDD1.n34 VDD1.n3 171.744
R64 VDD1.n34 VDD1.n33 171.744
R65 VDD1.n33 VDD1.n7 171.744
R66 VDD1.n26 VDD1.n7 171.744
R67 VDD1.n26 VDD1.n25 171.744
R68 VDD1.n25 VDD1.n11 171.744
R69 VDD1.n18 VDD1.n11 171.744
R70 VDD1.n18 VDD1.n17 171.744
R71 VDD1.n67 VDD1.n66 171.744
R72 VDD1.n67 VDD1.n60 171.744
R73 VDD1.n74 VDD1.n60 171.744
R74 VDD1.n75 VDD1.n74 171.744
R75 VDD1.n75 VDD1.n56 171.744
R76 VDD1.n82 VDD1.n56 171.744
R77 VDD1.n83 VDD1.n82 171.744
R78 VDD1.n83 VDD1.n52 171.744
R79 VDD1.n90 VDD1.n52 171.744
R80 VDD1.n91 VDD1.n90 171.744
R81 VDD1.n17 VDD1.t6 85.8723
R82 VDD1.n66 VDD1.t7 85.8723
R83 VDD1.n99 VDD1.n98 79.3391
R84 VDD1.n101 VDD1.n100 78.9615
R85 VDD1.n48 VDD1.n47 78.9615
R86 VDD1.n97 VDD1.n96 78.9613
R87 VDD1.n48 VDD1.n46 47.6963
R88 VDD1.n97 VDD1.n95 47.6963
R89 VDD1.n101 VDD1.n99 34.9082
R90 VDD1.n16 VDD1.n15 16.3894
R91 VDD1.n65 VDD1.n64 16.3894
R92 VDD1.n19 VDD1.n14 12.8005
R93 VDD1.n68 VDD1.n63 12.8005
R94 VDD1.n20 VDD1.n12 12.0247
R95 VDD1.n69 VDD1.n61 12.0247
R96 VDD1.n24 VDD1.n23 11.249
R97 VDD1.n73 VDD1.n72 11.249
R98 VDD1.n27 VDD1.n10 10.4732
R99 VDD1.n76 VDD1.n59 10.4732
R100 VDD1.n28 VDD1.n8 9.69747
R101 VDD1.n77 VDD1.n57 9.69747
R102 VDD1.n46 VDD1.n45 9.45567
R103 VDD1.n95 VDD1.n94 9.45567
R104 VDD1.n2 VDD1.n1 9.3005
R105 VDD1.n45 VDD1.n44 9.3005
R106 VDD1.n39 VDD1.n38 9.3005
R107 VDD1.n37 VDD1.n36 9.3005
R108 VDD1.n6 VDD1.n5 9.3005
R109 VDD1.n31 VDD1.n30 9.3005
R110 VDD1.n29 VDD1.n28 9.3005
R111 VDD1.n10 VDD1.n9 9.3005
R112 VDD1.n23 VDD1.n22 9.3005
R113 VDD1.n21 VDD1.n20 9.3005
R114 VDD1.n14 VDD1.n13 9.3005
R115 VDD1.n88 VDD1.n87 9.3005
R116 VDD1.n51 VDD1.n50 9.3005
R117 VDD1.n94 VDD1.n93 9.3005
R118 VDD1.n55 VDD1.n54 9.3005
R119 VDD1.n80 VDD1.n79 9.3005
R120 VDD1.n78 VDD1.n77 9.3005
R121 VDD1.n59 VDD1.n58 9.3005
R122 VDD1.n72 VDD1.n71 9.3005
R123 VDD1.n70 VDD1.n69 9.3005
R124 VDD1.n63 VDD1.n62 9.3005
R125 VDD1.n86 VDD1.n85 9.3005
R126 VDD1.n46 VDD1.n0 8.92171
R127 VDD1.n32 VDD1.n31 8.92171
R128 VDD1.n81 VDD1.n80 8.92171
R129 VDD1.n95 VDD1.n49 8.92171
R130 VDD1.n44 VDD1.n43 8.14595
R131 VDD1.n35 VDD1.n6 8.14595
R132 VDD1.n84 VDD1.n55 8.14595
R133 VDD1.n93 VDD1.n92 8.14595
R134 VDD1.n40 VDD1.n2 7.3702
R135 VDD1.n36 VDD1.n4 7.3702
R136 VDD1.n85 VDD1.n53 7.3702
R137 VDD1.n89 VDD1.n51 7.3702
R138 VDD1.n40 VDD1.n39 6.59444
R139 VDD1.n39 VDD1.n4 6.59444
R140 VDD1.n88 VDD1.n53 6.59444
R141 VDD1.n89 VDD1.n88 6.59444
R142 VDD1.n43 VDD1.n2 5.81868
R143 VDD1.n36 VDD1.n35 5.81868
R144 VDD1.n85 VDD1.n84 5.81868
R145 VDD1.n92 VDD1.n51 5.81868
R146 VDD1.n44 VDD1.n0 5.04292
R147 VDD1.n32 VDD1.n6 5.04292
R148 VDD1.n81 VDD1.n55 5.04292
R149 VDD1.n93 VDD1.n49 5.04292
R150 VDD1.n31 VDD1.n8 4.26717
R151 VDD1.n80 VDD1.n57 4.26717
R152 VDD1.n15 VDD1.n13 3.70987
R153 VDD1.n64 VDD1.n62 3.70987
R154 VDD1.n100 VDD1.t1 3.69845
R155 VDD1.n100 VDD1.t9 3.69845
R156 VDD1.n47 VDD1.t0 3.69845
R157 VDD1.n47 VDD1.t2 3.69845
R158 VDD1.n98 VDD1.t5 3.69845
R159 VDD1.n98 VDD1.t3 3.69845
R160 VDD1.n96 VDD1.t8 3.69845
R161 VDD1.n96 VDD1.t4 3.69845
R162 VDD1.n28 VDD1.n27 3.49141
R163 VDD1.n77 VDD1.n76 3.49141
R164 VDD1.n24 VDD1.n10 2.71565
R165 VDD1.n73 VDD1.n59 2.71565
R166 VDD1.n23 VDD1.n12 1.93989
R167 VDD1.n72 VDD1.n61 1.93989
R168 VDD1.n20 VDD1.n19 1.16414
R169 VDD1.n69 VDD1.n68 1.16414
R170 VDD1.n16 VDD1.n14 0.388379
R171 VDD1.n65 VDD1.n63 0.388379
R172 VDD1 VDD1.n101 0.3755
R173 VDD1 VDD1.n48 0.203086
R174 VDD1.n45 VDD1.n1 0.155672
R175 VDD1.n38 VDD1.n1 0.155672
R176 VDD1.n38 VDD1.n37 0.155672
R177 VDD1.n37 VDD1.n5 0.155672
R178 VDD1.n30 VDD1.n5 0.155672
R179 VDD1.n30 VDD1.n29 0.155672
R180 VDD1.n29 VDD1.n9 0.155672
R181 VDD1.n22 VDD1.n9 0.155672
R182 VDD1.n22 VDD1.n21 0.155672
R183 VDD1.n21 VDD1.n13 0.155672
R184 VDD1.n70 VDD1.n62 0.155672
R185 VDD1.n71 VDD1.n70 0.155672
R186 VDD1.n71 VDD1.n58 0.155672
R187 VDD1.n78 VDD1.n58 0.155672
R188 VDD1.n79 VDD1.n78 0.155672
R189 VDD1.n79 VDD1.n54 0.155672
R190 VDD1.n86 VDD1.n54 0.155672
R191 VDD1.n87 VDD1.n86 0.155672
R192 VDD1.n87 VDD1.n50 0.155672
R193 VDD1.n94 VDD1.n50 0.155672
R194 VDD1.n99 VDD1.n97 0.0895505
R195 VTAIL.n200 VTAIL.n158 756.745
R196 VTAIL.n44 VTAIL.n2 756.745
R197 VTAIL.n152 VTAIL.n110 756.745
R198 VTAIL.n100 VTAIL.n58 756.745
R199 VTAIL.n175 VTAIL.n174 585
R200 VTAIL.n177 VTAIL.n176 585
R201 VTAIL.n170 VTAIL.n169 585
R202 VTAIL.n183 VTAIL.n182 585
R203 VTAIL.n185 VTAIL.n184 585
R204 VTAIL.n166 VTAIL.n165 585
R205 VTAIL.n191 VTAIL.n190 585
R206 VTAIL.n193 VTAIL.n192 585
R207 VTAIL.n162 VTAIL.n161 585
R208 VTAIL.n199 VTAIL.n198 585
R209 VTAIL.n201 VTAIL.n200 585
R210 VTAIL.n19 VTAIL.n18 585
R211 VTAIL.n21 VTAIL.n20 585
R212 VTAIL.n14 VTAIL.n13 585
R213 VTAIL.n27 VTAIL.n26 585
R214 VTAIL.n29 VTAIL.n28 585
R215 VTAIL.n10 VTAIL.n9 585
R216 VTAIL.n35 VTAIL.n34 585
R217 VTAIL.n37 VTAIL.n36 585
R218 VTAIL.n6 VTAIL.n5 585
R219 VTAIL.n43 VTAIL.n42 585
R220 VTAIL.n45 VTAIL.n44 585
R221 VTAIL.n153 VTAIL.n152 585
R222 VTAIL.n151 VTAIL.n150 585
R223 VTAIL.n114 VTAIL.n113 585
R224 VTAIL.n145 VTAIL.n144 585
R225 VTAIL.n143 VTAIL.n142 585
R226 VTAIL.n118 VTAIL.n117 585
R227 VTAIL.n137 VTAIL.n136 585
R228 VTAIL.n135 VTAIL.n134 585
R229 VTAIL.n122 VTAIL.n121 585
R230 VTAIL.n129 VTAIL.n128 585
R231 VTAIL.n127 VTAIL.n126 585
R232 VTAIL.n101 VTAIL.n100 585
R233 VTAIL.n99 VTAIL.n98 585
R234 VTAIL.n62 VTAIL.n61 585
R235 VTAIL.n93 VTAIL.n92 585
R236 VTAIL.n91 VTAIL.n90 585
R237 VTAIL.n66 VTAIL.n65 585
R238 VTAIL.n85 VTAIL.n84 585
R239 VTAIL.n83 VTAIL.n82 585
R240 VTAIL.n70 VTAIL.n69 585
R241 VTAIL.n77 VTAIL.n76 585
R242 VTAIL.n75 VTAIL.n74 585
R243 VTAIL.n173 VTAIL.t1 327.469
R244 VTAIL.n17 VTAIL.t13 327.469
R245 VTAIL.n125 VTAIL.t9 327.469
R246 VTAIL.n73 VTAIL.t18 327.469
R247 VTAIL.n176 VTAIL.n175 171.744
R248 VTAIL.n176 VTAIL.n169 171.744
R249 VTAIL.n183 VTAIL.n169 171.744
R250 VTAIL.n184 VTAIL.n183 171.744
R251 VTAIL.n184 VTAIL.n165 171.744
R252 VTAIL.n191 VTAIL.n165 171.744
R253 VTAIL.n192 VTAIL.n191 171.744
R254 VTAIL.n192 VTAIL.n161 171.744
R255 VTAIL.n199 VTAIL.n161 171.744
R256 VTAIL.n200 VTAIL.n199 171.744
R257 VTAIL.n20 VTAIL.n19 171.744
R258 VTAIL.n20 VTAIL.n13 171.744
R259 VTAIL.n27 VTAIL.n13 171.744
R260 VTAIL.n28 VTAIL.n27 171.744
R261 VTAIL.n28 VTAIL.n9 171.744
R262 VTAIL.n35 VTAIL.n9 171.744
R263 VTAIL.n36 VTAIL.n35 171.744
R264 VTAIL.n36 VTAIL.n5 171.744
R265 VTAIL.n43 VTAIL.n5 171.744
R266 VTAIL.n44 VTAIL.n43 171.744
R267 VTAIL.n152 VTAIL.n151 171.744
R268 VTAIL.n151 VTAIL.n113 171.744
R269 VTAIL.n144 VTAIL.n113 171.744
R270 VTAIL.n144 VTAIL.n143 171.744
R271 VTAIL.n143 VTAIL.n117 171.744
R272 VTAIL.n136 VTAIL.n117 171.744
R273 VTAIL.n136 VTAIL.n135 171.744
R274 VTAIL.n135 VTAIL.n121 171.744
R275 VTAIL.n128 VTAIL.n121 171.744
R276 VTAIL.n128 VTAIL.n127 171.744
R277 VTAIL.n100 VTAIL.n99 171.744
R278 VTAIL.n99 VTAIL.n61 171.744
R279 VTAIL.n92 VTAIL.n61 171.744
R280 VTAIL.n92 VTAIL.n91 171.744
R281 VTAIL.n91 VTAIL.n65 171.744
R282 VTAIL.n84 VTAIL.n65 171.744
R283 VTAIL.n84 VTAIL.n83 171.744
R284 VTAIL.n83 VTAIL.n69 171.744
R285 VTAIL.n76 VTAIL.n69 171.744
R286 VTAIL.n76 VTAIL.n75 171.744
R287 VTAIL.n175 VTAIL.t1 85.8723
R288 VTAIL.n19 VTAIL.t13 85.8723
R289 VTAIL.n127 VTAIL.t9 85.8723
R290 VTAIL.n75 VTAIL.t18 85.8723
R291 VTAIL.n109 VTAIL.n108 62.2827
R292 VTAIL.n107 VTAIL.n106 62.2827
R293 VTAIL.n57 VTAIL.n56 62.2827
R294 VTAIL.n55 VTAIL.n54 62.2827
R295 VTAIL.n207 VTAIL.n206 62.2825
R296 VTAIL.n1 VTAIL.n0 62.2825
R297 VTAIL.n51 VTAIL.n50 62.2825
R298 VTAIL.n53 VTAIL.n52 62.2825
R299 VTAIL.n205 VTAIL.n204 30.4399
R300 VTAIL.n49 VTAIL.n48 30.4399
R301 VTAIL.n157 VTAIL.n156 30.4399
R302 VTAIL.n105 VTAIL.n104 30.4399
R303 VTAIL.n55 VTAIL.n53 21.0996
R304 VTAIL.n205 VTAIL.n157 20.5221
R305 VTAIL.n174 VTAIL.n173 16.3894
R306 VTAIL.n18 VTAIL.n17 16.3894
R307 VTAIL.n126 VTAIL.n125 16.3894
R308 VTAIL.n74 VTAIL.n73 16.3894
R309 VTAIL.n177 VTAIL.n172 12.8005
R310 VTAIL.n21 VTAIL.n16 12.8005
R311 VTAIL.n129 VTAIL.n124 12.8005
R312 VTAIL.n77 VTAIL.n72 12.8005
R313 VTAIL.n178 VTAIL.n170 12.0247
R314 VTAIL.n22 VTAIL.n14 12.0247
R315 VTAIL.n130 VTAIL.n122 12.0247
R316 VTAIL.n78 VTAIL.n70 12.0247
R317 VTAIL.n182 VTAIL.n181 11.249
R318 VTAIL.n26 VTAIL.n25 11.249
R319 VTAIL.n134 VTAIL.n133 11.249
R320 VTAIL.n82 VTAIL.n81 11.249
R321 VTAIL.n185 VTAIL.n168 10.4732
R322 VTAIL.n29 VTAIL.n12 10.4732
R323 VTAIL.n137 VTAIL.n120 10.4732
R324 VTAIL.n85 VTAIL.n68 10.4732
R325 VTAIL.n186 VTAIL.n166 9.69747
R326 VTAIL.n30 VTAIL.n10 9.69747
R327 VTAIL.n138 VTAIL.n118 9.69747
R328 VTAIL.n86 VTAIL.n66 9.69747
R329 VTAIL.n204 VTAIL.n203 9.45567
R330 VTAIL.n48 VTAIL.n47 9.45567
R331 VTAIL.n156 VTAIL.n155 9.45567
R332 VTAIL.n104 VTAIL.n103 9.45567
R333 VTAIL.n197 VTAIL.n196 9.3005
R334 VTAIL.n160 VTAIL.n159 9.3005
R335 VTAIL.n203 VTAIL.n202 9.3005
R336 VTAIL.n164 VTAIL.n163 9.3005
R337 VTAIL.n189 VTAIL.n188 9.3005
R338 VTAIL.n187 VTAIL.n186 9.3005
R339 VTAIL.n168 VTAIL.n167 9.3005
R340 VTAIL.n181 VTAIL.n180 9.3005
R341 VTAIL.n179 VTAIL.n178 9.3005
R342 VTAIL.n172 VTAIL.n171 9.3005
R343 VTAIL.n195 VTAIL.n194 9.3005
R344 VTAIL.n41 VTAIL.n40 9.3005
R345 VTAIL.n4 VTAIL.n3 9.3005
R346 VTAIL.n47 VTAIL.n46 9.3005
R347 VTAIL.n8 VTAIL.n7 9.3005
R348 VTAIL.n33 VTAIL.n32 9.3005
R349 VTAIL.n31 VTAIL.n30 9.3005
R350 VTAIL.n12 VTAIL.n11 9.3005
R351 VTAIL.n25 VTAIL.n24 9.3005
R352 VTAIL.n23 VTAIL.n22 9.3005
R353 VTAIL.n16 VTAIL.n15 9.3005
R354 VTAIL.n39 VTAIL.n38 9.3005
R355 VTAIL.n112 VTAIL.n111 9.3005
R356 VTAIL.n149 VTAIL.n148 9.3005
R357 VTAIL.n147 VTAIL.n146 9.3005
R358 VTAIL.n116 VTAIL.n115 9.3005
R359 VTAIL.n141 VTAIL.n140 9.3005
R360 VTAIL.n139 VTAIL.n138 9.3005
R361 VTAIL.n120 VTAIL.n119 9.3005
R362 VTAIL.n133 VTAIL.n132 9.3005
R363 VTAIL.n131 VTAIL.n130 9.3005
R364 VTAIL.n124 VTAIL.n123 9.3005
R365 VTAIL.n155 VTAIL.n154 9.3005
R366 VTAIL.n60 VTAIL.n59 9.3005
R367 VTAIL.n103 VTAIL.n102 9.3005
R368 VTAIL.n97 VTAIL.n96 9.3005
R369 VTAIL.n95 VTAIL.n94 9.3005
R370 VTAIL.n64 VTAIL.n63 9.3005
R371 VTAIL.n89 VTAIL.n88 9.3005
R372 VTAIL.n87 VTAIL.n86 9.3005
R373 VTAIL.n68 VTAIL.n67 9.3005
R374 VTAIL.n81 VTAIL.n80 9.3005
R375 VTAIL.n79 VTAIL.n78 9.3005
R376 VTAIL.n72 VTAIL.n71 9.3005
R377 VTAIL.n190 VTAIL.n189 8.92171
R378 VTAIL.n204 VTAIL.n158 8.92171
R379 VTAIL.n34 VTAIL.n33 8.92171
R380 VTAIL.n48 VTAIL.n2 8.92171
R381 VTAIL.n156 VTAIL.n110 8.92171
R382 VTAIL.n142 VTAIL.n141 8.92171
R383 VTAIL.n104 VTAIL.n58 8.92171
R384 VTAIL.n90 VTAIL.n89 8.92171
R385 VTAIL.n193 VTAIL.n164 8.14595
R386 VTAIL.n202 VTAIL.n201 8.14595
R387 VTAIL.n37 VTAIL.n8 8.14595
R388 VTAIL.n46 VTAIL.n45 8.14595
R389 VTAIL.n154 VTAIL.n153 8.14595
R390 VTAIL.n145 VTAIL.n116 8.14595
R391 VTAIL.n102 VTAIL.n101 8.14595
R392 VTAIL.n93 VTAIL.n64 8.14595
R393 VTAIL.n194 VTAIL.n162 7.3702
R394 VTAIL.n198 VTAIL.n160 7.3702
R395 VTAIL.n38 VTAIL.n6 7.3702
R396 VTAIL.n42 VTAIL.n4 7.3702
R397 VTAIL.n150 VTAIL.n112 7.3702
R398 VTAIL.n146 VTAIL.n114 7.3702
R399 VTAIL.n98 VTAIL.n60 7.3702
R400 VTAIL.n94 VTAIL.n62 7.3702
R401 VTAIL.n197 VTAIL.n162 6.59444
R402 VTAIL.n198 VTAIL.n197 6.59444
R403 VTAIL.n41 VTAIL.n6 6.59444
R404 VTAIL.n42 VTAIL.n41 6.59444
R405 VTAIL.n150 VTAIL.n149 6.59444
R406 VTAIL.n149 VTAIL.n114 6.59444
R407 VTAIL.n98 VTAIL.n97 6.59444
R408 VTAIL.n97 VTAIL.n62 6.59444
R409 VTAIL.n194 VTAIL.n193 5.81868
R410 VTAIL.n201 VTAIL.n160 5.81868
R411 VTAIL.n38 VTAIL.n37 5.81868
R412 VTAIL.n45 VTAIL.n4 5.81868
R413 VTAIL.n153 VTAIL.n112 5.81868
R414 VTAIL.n146 VTAIL.n145 5.81868
R415 VTAIL.n101 VTAIL.n60 5.81868
R416 VTAIL.n94 VTAIL.n93 5.81868
R417 VTAIL.n190 VTAIL.n164 5.04292
R418 VTAIL.n202 VTAIL.n158 5.04292
R419 VTAIL.n34 VTAIL.n8 5.04292
R420 VTAIL.n46 VTAIL.n2 5.04292
R421 VTAIL.n154 VTAIL.n110 5.04292
R422 VTAIL.n142 VTAIL.n116 5.04292
R423 VTAIL.n102 VTAIL.n58 5.04292
R424 VTAIL.n90 VTAIL.n64 5.04292
R425 VTAIL.n189 VTAIL.n166 4.26717
R426 VTAIL.n33 VTAIL.n10 4.26717
R427 VTAIL.n141 VTAIL.n118 4.26717
R428 VTAIL.n89 VTAIL.n66 4.26717
R429 VTAIL.n125 VTAIL.n123 3.70987
R430 VTAIL.n73 VTAIL.n71 3.70987
R431 VTAIL.n173 VTAIL.n171 3.70987
R432 VTAIL.n17 VTAIL.n15 3.70987
R433 VTAIL.n206 VTAIL.t0 3.69845
R434 VTAIL.n206 VTAIL.t2 3.69845
R435 VTAIL.n0 VTAIL.t5 3.69845
R436 VTAIL.n0 VTAIL.t19 3.69845
R437 VTAIL.n50 VTAIL.t10 3.69845
R438 VTAIL.n50 VTAIL.t15 3.69845
R439 VTAIL.n52 VTAIL.t12 3.69845
R440 VTAIL.n52 VTAIL.t11 3.69845
R441 VTAIL.n108 VTAIL.t6 3.69845
R442 VTAIL.n108 VTAIL.t7 3.69845
R443 VTAIL.n106 VTAIL.t8 3.69845
R444 VTAIL.n106 VTAIL.t14 3.69845
R445 VTAIL.n56 VTAIL.t4 3.69845
R446 VTAIL.n56 VTAIL.t16 3.69845
R447 VTAIL.n54 VTAIL.t17 3.69845
R448 VTAIL.n54 VTAIL.t3 3.69845
R449 VTAIL.n186 VTAIL.n185 3.49141
R450 VTAIL.n30 VTAIL.n29 3.49141
R451 VTAIL.n138 VTAIL.n137 3.49141
R452 VTAIL.n86 VTAIL.n85 3.49141
R453 VTAIL.n182 VTAIL.n168 2.71565
R454 VTAIL.n26 VTAIL.n12 2.71565
R455 VTAIL.n134 VTAIL.n120 2.71565
R456 VTAIL.n82 VTAIL.n68 2.71565
R457 VTAIL.n181 VTAIL.n170 1.93989
R458 VTAIL.n25 VTAIL.n14 1.93989
R459 VTAIL.n133 VTAIL.n122 1.93989
R460 VTAIL.n81 VTAIL.n70 1.93989
R461 VTAIL.n178 VTAIL.n177 1.16414
R462 VTAIL.n22 VTAIL.n21 1.16414
R463 VTAIL.n130 VTAIL.n129 1.16414
R464 VTAIL.n78 VTAIL.n77 1.16414
R465 VTAIL.n107 VTAIL.n105 0.759121
R466 VTAIL.n49 VTAIL.n1 0.759121
R467 VTAIL.n57 VTAIL.n55 0.578086
R468 VTAIL.n105 VTAIL.n57 0.578086
R469 VTAIL.n109 VTAIL.n107 0.578086
R470 VTAIL.n157 VTAIL.n109 0.578086
R471 VTAIL.n53 VTAIL.n51 0.578086
R472 VTAIL.n51 VTAIL.n49 0.578086
R473 VTAIL.n207 VTAIL.n205 0.578086
R474 VTAIL VTAIL.n1 0.491879
R475 VTAIL.n174 VTAIL.n172 0.388379
R476 VTAIL.n18 VTAIL.n16 0.388379
R477 VTAIL.n126 VTAIL.n124 0.388379
R478 VTAIL.n74 VTAIL.n72 0.388379
R479 VTAIL.n179 VTAIL.n171 0.155672
R480 VTAIL.n180 VTAIL.n179 0.155672
R481 VTAIL.n180 VTAIL.n167 0.155672
R482 VTAIL.n187 VTAIL.n167 0.155672
R483 VTAIL.n188 VTAIL.n187 0.155672
R484 VTAIL.n188 VTAIL.n163 0.155672
R485 VTAIL.n195 VTAIL.n163 0.155672
R486 VTAIL.n196 VTAIL.n195 0.155672
R487 VTAIL.n196 VTAIL.n159 0.155672
R488 VTAIL.n203 VTAIL.n159 0.155672
R489 VTAIL.n23 VTAIL.n15 0.155672
R490 VTAIL.n24 VTAIL.n23 0.155672
R491 VTAIL.n24 VTAIL.n11 0.155672
R492 VTAIL.n31 VTAIL.n11 0.155672
R493 VTAIL.n32 VTAIL.n31 0.155672
R494 VTAIL.n32 VTAIL.n7 0.155672
R495 VTAIL.n39 VTAIL.n7 0.155672
R496 VTAIL.n40 VTAIL.n39 0.155672
R497 VTAIL.n40 VTAIL.n3 0.155672
R498 VTAIL.n47 VTAIL.n3 0.155672
R499 VTAIL.n155 VTAIL.n111 0.155672
R500 VTAIL.n148 VTAIL.n111 0.155672
R501 VTAIL.n148 VTAIL.n147 0.155672
R502 VTAIL.n147 VTAIL.n115 0.155672
R503 VTAIL.n140 VTAIL.n115 0.155672
R504 VTAIL.n140 VTAIL.n139 0.155672
R505 VTAIL.n139 VTAIL.n119 0.155672
R506 VTAIL.n132 VTAIL.n119 0.155672
R507 VTAIL.n132 VTAIL.n131 0.155672
R508 VTAIL.n131 VTAIL.n123 0.155672
R509 VTAIL.n103 VTAIL.n59 0.155672
R510 VTAIL.n96 VTAIL.n59 0.155672
R511 VTAIL.n96 VTAIL.n95 0.155672
R512 VTAIL.n95 VTAIL.n63 0.155672
R513 VTAIL.n88 VTAIL.n63 0.155672
R514 VTAIL.n88 VTAIL.n87 0.155672
R515 VTAIL.n87 VTAIL.n67 0.155672
R516 VTAIL.n80 VTAIL.n67 0.155672
R517 VTAIL.n80 VTAIL.n79 0.155672
R518 VTAIL.n79 VTAIL.n71 0.155672
R519 VTAIL VTAIL.n207 0.0867069
R520 VN.n2 VN.t8 775.037
R521 VN.n10 VN.t2 775.037
R522 VN.n6 VN.t6 764.134
R523 VN.n14 VN.t1 764.134
R524 VN.n1 VN.t4 739.303
R525 VN.n4 VN.t3 739.303
R526 VN.n5 VN.t7 739.303
R527 VN.n9 VN.t0 739.303
R528 VN.n12 VN.t9 739.303
R529 VN.n13 VN.t5 739.303
R530 VN.n7 VN.n6 161.3
R531 VN.n15 VN.n14 161.3
R532 VN.n13 VN.n8 161.3
R533 VN.n12 VN.n11 161.3
R534 VN.n5 VN.n0 161.3
R535 VN.n4 VN.n3 161.3
R536 VN.n11 VN.n10 75.4397
R537 VN.n3 VN.n2 75.4397
R538 VN.n4 VN.n1 48.2005
R539 VN.n5 VN.n4 48.2005
R540 VN.n12 VN.n9 48.2005
R541 VN.n13 VN.n12 48.2005
R542 VN VN.n15 38.9001
R543 VN.n6 VN.n5 23.3702
R544 VN.n14 VN.n13 23.3702
R545 VN.n10 VN.n9 10.8906
R546 VN.n2 VN.n1 10.8906
R547 VN.n15 VN.n8 0.189894
R548 VN.n11 VN.n8 0.189894
R549 VN.n3 VN.n0 0.189894
R550 VN.n7 VN.n0 0.189894
R551 VN VN.n7 0.0516364
R552 VDD2.n93 VDD2.n51 756.745
R553 VDD2.n42 VDD2.n0 756.745
R554 VDD2.n94 VDD2.n93 585
R555 VDD2.n92 VDD2.n91 585
R556 VDD2.n55 VDD2.n54 585
R557 VDD2.n86 VDD2.n85 585
R558 VDD2.n84 VDD2.n83 585
R559 VDD2.n59 VDD2.n58 585
R560 VDD2.n78 VDD2.n77 585
R561 VDD2.n76 VDD2.n75 585
R562 VDD2.n63 VDD2.n62 585
R563 VDD2.n70 VDD2.n69 585
R564 VDD2.n68 VDD2.n67 585
R565 VDD2.n17 VDD2.n16 585
R566 VDD2.n19 VDD2.n18 585
R567 VDD2.n12 VDD2.n11 585
R568 VDD2.n25 VDD2.n24 585
R569 VDD2.n27 VDD2.n26 585
R570 VDD2.n8 VDD2.n7 585
R571 VDD2.n33 VDD2.n32 585
R572 VDD2.n35 VDD2.n34 585
R573 VDD2.n4 VDD2.n3 585
R574 VDD2.n41 VDD2.n40 585
R575 VDD2.n43 VDD2.n42 585
R576 VDD2.n66 VDD2.t8 327.469
R577 VDD2.n15 VDD2.t1 327.469
R578 VDD2.n93 VDD2.n92 171.744
R579 VDD2.n92 VDD2.n54 171.744
R580 VDD2.n85 VDD2.n54 171.744
R581 VDD2.n85 VDD2.n84 171.744
R582 VDD2.n84 VDD2.n58 171.744
R583 VDD2.n77 VDD2.n58 171.744
R584 VDD2.n77 VDD2.n76 171.744
R585 VDD2.n76 VDD2.n62 171.744
R586 VDD2.n69 VDD2.n62 171.744
R587 VDD2.n69 VDD2.n68 171.744
R588 VDD2.n18 VDD2.n17 171.744
R589 VDD2.n18 VDD2.n11 171.744
R590 VDD2.n25 VDD2.n11 171.744
R591 VDD2.n26 VDD2.n25 171.744
R592 VDD2.n26 VDD2.n7 171.744
R593 VDD2.n33 VDD2.n7 171.744
R594 VDD2.n34 VDD2.n33 171.744
R595 VDD2.n34 VDD2.n3 171.744
R596 VDD2.n41 VDD2.n3 171.744
R597 VDD2.n42 VDD2.n41 171.744
R598 VDD2.n68 VDD2.t8 85.8723
R599 VDD2.n17 VDD2.t1 85.8723
R600 VDD2.n50 VDD2.n49 79.3391
R601 VDD2 VDD2.n101 79.3365
R602 VDD2.n100 VDD2.n99 78.9615
R603 VDD2.n48 VDD2.n47 78.9613
R604 VDD2.n48 VDD2.n46 47.6963
R605 VDD2.n98 VDD2.n97 47.1187
R606 VDD2.n98 VDD2.n50 34.0364
R607 VDD2.n67 VDD2.n66 16.3894
R608 VDD2.n16 VDD2.n15 16.3894
R609 VDD2.n70 VDD2.n65 12.8005
R610 VDD2.n19 VDD2.n14 12.8005
R611 VDD2.n71 VDD2.n63 12.0247
R612 VDD2.n20 VDD2.n12 12.0247
R613 VDD2.n75 VDD2.n74 11.249
R614 VDD2.n24 VDD2.n23 11.249
R615 VDD2.n78 VDD2.n61 10.4732
R616 VDD2.n27 VDD2.n10 10.4732
R617 VDD2.n79 VDD2.n59 9.69747
R618 VDD2.n28 VDD2.n8 9.69747
R619 VDD2.n97 VDD2.n96 9.45567
R620 VDD2.n46 VDD2.n45 9.45567
R621 VDD2.n53 VDD2.n52 9.3005
R622 VDD2.n96 VDD2.n95 9.3005
R623 VDD2.n90 VDD2.n89 9.3005
R624 VDD2.n88 VDD2.n87 9.3005
R625 VDD2.n57 VDD2.n56 9.3005
R626 VDD2.n82 VDD2.n81 9.3005
R627 VDD2.n80 VDD2.n79 9.3005
R628 VDD2.n61 VDD2.n60 9.3005
R629 VDD2.n74 VDD2.n73 9.3005
R630 VDD2.n72 VDD2.n71 9.3005
R631 VDD2.n65 VDD2.n64 9.3005
R632 VDD2.n39 VDD2.n38 9.3005
R633 VDD2.n2 VDD2.n1 9.3005
R634 VDD2.n45 VDD2.n44 9.3005
R635 VDD2.n6 VDD2.n5 9.3005
R636 VDD2.n31 VDD2.n30 9.3005
R637 VDD2.n29 VDD2.n28 9.3005
R638 VDD2.n10 VDD2.n9 9.3005
R639 VDD2.n23 VDD2.n22 9.3005
R640 VDD2.n21 VDD2.n20 9.3005
R641 VDD2.n14 VDD2.n13 9.3005
R642 VDD2.n37 VDD2.n36 9.3005
R643 VDD2.n97 VDD2.n51 8.92171
R644 VDD2.n83 VDD2.n82 8.92171
R645 VDD2.n32 VDD2.n31 8.92171
R646 VDD2.n46 VDD2.n0 8.92171
R647 VDD2.n95 VDD2.n94 8.14595
R648 VDD2.n86 VDD2.n57 8.14595
R649 VDD2.n35 VDD2.n6 8.14595
R650 VDD2.n44 VDD2.n43 8.14595
R651 VDD2.n91 VDD2.n53 7.3702
R652 VDD2.n87 VDD2.n55 7.3702
R653 VDD2.n36 VDD2.n4 7.3702
R654 VDD2.n40 VDD2.n2 7.3702
R655 VDD2.n91 VDD2.n90 6.59444
R656 VDD2.n90 VDD2.n55 6.59444
R657 VDD2.n39 VDD2.n4 6.59444
R658 VDD2.n40 VDD2.n39 6.59444
R659 VDD2.n94 VDD2.n53 5.81868
R660 VDD2.n87 VDD2.n86 5.81868
R661 VDD2.n36 VDD2.n35 5.81868
R662 VDD2.n43 VDD2.n2 5.81868
R663 VDD2.n95 VDD2.n51 5.04292
R664 VDD2.n83 VDD2.n57 5.04292
R665 VDD2.n32 VDD2.n6 5.04292
R666 VDD2.n44 VDD2.n0 5.04292
R667 VDD2.n82 VDD2.n59 4.26717
R668 VDD2.n31 VDD2.n8 4.26717
R669 VDD2.n66 VDD2.n64 3.70987
R670 VDD2.n15 VDD2.n13 3.70987
R671 VDD2.n101 VDD2.t9 3.69845
R672 VDD2.n101 VDD2.t7 3.69845
R673 VDD2.n99 VDD2.t4 3.69845
R674 VDD2.n99 VDD2.t0 3.69845
R675 VDD2.n49 VDD2.t2 3.69845
R676 VDD2.n49 VDD2.t3 3.69845
R677 VDD2.n47 VDD2.t5 3.69845
R678 VDD2.n47 VDD2.t6 3.69845
R679 VDD2.n79 VDD2.n78 3.49141
R680 VDD2.n28 VDD2.n27 3.49141
R681 VDD2.n75 VDD2.n61 2.71565
R682 VDD2.n24 VDD2.n10 2.71565
R683 VDD2.n74 VDD2.n63 1.93989
R684 VDD2.n23 VDD2.n12 1.93989
R685 VDD2.n71 VDD2.n70 1.16414
R686 VDD2.n20 VDD2.n19 1.16414
R687 VDD2.n100 VDD2.n98 0.578086
R688 VDD2.n67 VDD2.n65 0.388379
R689 VDD2.n16 VDD2.n14 0.388379
R690 VDD2 VDD2.n100 0.203086
R691 VDD2.n96 VDD2.n52 0.155672
R692 VDD2.n89 VDD2.n52 0.155672
R693 VDD2.n89 VDD2.n88 0.155672
R694 VDD2.n88 VDD2.n56 0.155672
R695 VDD2.n81 VDD2.n56 0.155672
R696 VDD2.n81 VDD2.n80 0.155672
R697 VDD2.n80 VDD2.n60 0.155672
R698 VDD2.n73 VDD2.n60 0.155672
R699 VDD2.n73 VDD2.n72 0.155672
R700 VDD2.n72 VDD2.n64 0.155672
R701 VDD2.n21 VDD2.n13 0.155672
R702 VDD2.n22 VDD2.n21 0.155672
R703 VDD2.n22 VDD2.n9 0.155672
R704 VDD2.n29 VDD2.n9 0.155672
R705 VDD2.n30 VDD2.n29 0.155672
R706 VDD2.n30 VDD2.n5 0.155672
R707 VDD2.n37 VDD2.n5 0.155672
R708 VDD2.n38 VDD2.n37 0.155672
R709 VDD2.n38 VDD2.n1 0.155672
R710 VDD2.n45 VDD2.n1 0.155672
R711 VDD2.n50 VDD2.n48 0.0895505
R712 B.n90 B.t0 835.135
R713 B.n98 B.t3 835.135
R714 B.n28 B.t9 835.135
R715 B.n36 B.t6 835.135
R716 B.n328 B.n53 585
R717 B.n330 B.n329 585
R718 B.n331 B.n52 585
R719 B.n333 B.n332 585
R720 B.n334 B.n51 585
R721 B.n336 B.n335 585
R722 B.n337 B.n50 585
R723 B.n339 B.n338 585
R724 B.n340 B.n49 585
R725 B.n342 B.n341 585
R726 B.n343 B.n48 585
R727 B.n345 B.n344 585
R728 B.n346 B.n47 585
R729 B.n348 B.n347 585
R730 B.n349 B.n46 585
R731 B.n351 B.n350 585
R732 B.n352 B.n45 585
R733 B.n354 B.n353 585
R734 B.n355 B.n44 585
R735 B.n357 B.n356 585
R736 B.n358 B.n43 585
R737 B.n360 B.n359 585
R738 B.n361 B.n42 585
R739 B.n363 B.n362 585
R740 B.n364 B.n41 585
R741 B.n366 B.n365 585
R742 B.n367 B.n40 585
R743 B.n369 B.n368 585
R744 B.n370 B.n39 585
R745 B.n372 B.n371 585
R746 B.n373 B.n38 585
R747 B.n375 B.n374 585
R748 B.n377 B.n35 585
R749 B.n379 B.n378 585
R750 B.n380 B.n34 585
R751 B.n382 B.n381 585
R752 B.n383 B.n33 585
R753 B.n385 B.n384 585
R754 B.n386 B.n32 585
R755 B.n388 B.n387 585
R756 B.n389 B.n31 585
R757 B.n391 B.n390 585
R758 B.n393 B.n392 585
R759 B.n394 B.n27 585
R760 B.n396 B.n395 585
R761 B.n397 B.n26 585
R762 B.n399 B.n398 585
R763 B.n400 B.n25 585
R764 B.n402 B.n401 585
R765 B.n403 B.n24 585
R766 B.n405 B.n404 585
R767 B.n406 B.n23 585
R768 B.n408 B.n407 585
R769 B.n409 B.n22 585
R770 B.n411 B.n410 585
R771 B.n412 B.n21 585
R772 B.n414 B.n413 585
R773 B.n415 B.n20 585
R774 B.n417 B.n416 585
R775 B.n418 B.n19 585
R776 B.n420 B.n419 585
R777 B.n421 B.n18 585
R778 B.n423 B.n422 585
R779 B.n424 B.n17 585
R780 B.n426 B.n425 585
R781 B.n427 B.n16 585
R782 B.n429 B.n428 585
R783 B.n430 B.n15 585
R784 B.n432 B.n431 585
R785 B.n433 B.n14 585
R786 B.n435 B.n434 585
R787 B.n436 B.n13 585
R788 B.n438 B.n437 585
R789 B.n439 B.n12 585
R790 B.n327 B.n326 585
R791 B.n325 B.n54 585
R792 B.n324 B.n323 585
R793 B.n322 B.n55 585
R794 B.n321 B.n320 585
R795 B.n319 B.n56 585
R796 B.n318 B.n317 585
R797 B.n316 B.n57 585
R798 B.n315 B.n314 585
R799 B.n313 B.n58 585
R800 B.n312 B.n311 585
R801 B.n310 B.n59 585
R802 B.n309 B.n308 585
R803 B.n307 B.n60 585
R804 B.n306 B.n305 585
R805 B.n304 B.n61 585
R806 B.n303 B.n302 585
R807 B.n301 B.n62 585
R808 B.n300 B.n299 585
R809 B.n298 B.n63 585
R810 B.n297 B.n296 585
R811 B.n295 B.n64 585
R812 B.n294 B.n293 585
R813 B.n292 B.n65 585
R814 B.n291 B.n290 585
R815 B.n289 B.n66 585
R816 B.n288 B.n287 585
R817 B.n286 B.n67 585
R818 B.n285 B.n284 585
R819 B.n283 B.n68 585
R820 B.n282 B.n281 585
R821 B.n280 B.n69 585
R822 B.n279 B.n278 585
R823 B.n277 B.n70 585
R824 B.n276 B.n275 585
R825 B.n274 B.n71 585
R826 B.n273 B.n272 585
R827 B.n271 B.n72 585
R828 B.n270 B.n269 585
R829 B.n268 B.n73 585
R830 B.n267 B.n266 585
R831 B.n154 B.n115 585
R832 B.n156 B.n155 585
R833 B.n157 B.n114 585
R834 B.n159 B.n158 585
R835 B.n160 B.n113 585
R836 B.n162 B.n161 585
R837 B.n163 B.n112 585
R838 B.n165 B.n164 585
R839 B.n166 B.n111 585
R840 B.n168 B.n167 585
R841 B.n169 B.n110 585
R842 B.n171 B.n170 585
R843 B.n172 B.n109 585
R844 B.n174 B.n173 585
R845 B.n175 B.n108 585
R846 B.n177 B.n176 585
R847 B.n178 B.n107 585
R848 B.n180 B.n179 585
R849 B.n181 B.n106 585
R850 B.n183 B.n182 585
R851 B.n184 B.n105 585
R852 B.n186 B.n185 585
R853 B.n187 B.n104 585
R854 B.n189 B.n188 585
R855 B.n190 B.n103 585
R856 B.n192 B.n191 585
R857 B.n193 B.n102 585
R858 B.n195 B.n194 585
R859 B.n196 B.n101 585
R860 B.n198 B.n197 585
R861 B.n199 B.n100 585
R862 B.n201 B.n200 585
R863 B.n203 B.n97 585
R864 B.n205 B.n204 585
R865 B.n206 B.n96 585
R866 B.n208 B.n207 585
R867 B.n209 B.n95 585
R868 B.n211 B.n210 585
R869 B.n212 B.n94 585
R870 B.n214 B.n213 585
R871 B.n215 B.n93 585
R872 B.n217 B.n216 585
R873 B.n219 B.n218 585
R874 B.n220 B.n89 585
R875 B.n222 B.n221 585
R876 B.n223 B.n88 585
R877 B.n225 B.n224 585
R878 B.n226 B.n87 585
R879 B.n228 B.n227 585
R880 B.n229 B.n86 585
R881 B.n231 B.n230 585
R882 B.n232 B.n85 585
R883 B.n234 B.n233 585
R884 B.n235 B.n84 585
R885 B.n237 B.n236 585
R886 B.n238 B.n83 585
R887 B.n240 B.n239 585
R888 B.n241 B.n82 585
R889 B.n243 B.n242 585
R890 B.n244 B.n81 585
R891 B.n246 B.n245 585
R892 B.n247 B.n80 585
R893 B.n249 B.n248 585
R894 B.n250 B.n79 585
R895 B.n252 B.n251 585
R896 B.n253 B.n78 585
R897 B.n255 B.n254 585
R898 B.n256 B.n77 585
R899 B.n258 B.n257 585
R900 B.n259 B.n76 585
R901 B.n261 B.n260 585
R902 B.n262 B.n75 585
R903 B.n264 B.n263 585
R904 B.n265 B.n74 585
R905 B.n153 B.n152 585
R906 B.n151 B.n116 585
R907 B.n150 B.n149 585
R908 B.n148 B.n117 585
R909 B.n147 B.n146 585
R910 B.n145 B.n118 585
R911 B.n144 B.n143 585
R912 B.n142 B.n119 585
R913 B.n141 B.n140 585
R914 B.n139 B.n120 585
R915 B.n138 B.n137 585
R916 B.n136 B.n121 585
R917 B.n135 B.n134 585
R918 B.n133 B.n122 585
R919 B.n132 B.n131 585
R920 B.n130 B.n123 585
R921 B.n129 B.n128 585
R922 B.n127 B.n124 585
R923 B.n126 B.n125 585
R924 B.n2 B.n0 585
R925 B.n469 B.n1 585
R926 B.n468 B.n467 585
R927 B.n466 B.n3 585
R928 B.n465 B.n464 585
R929 B.n463 B.n4 585
R930 B.n462 B.n461 585
R931 B.n460 B.n5 585
R932 B.n459 B.n458 585
R933 B.n457 B.n6 585
R934 B.n456 B.n455 585
R935 B.n454 B.n7 585
R936 B.n453 B.n452 585
R937 B.n451 B.n8 585
R938 B.n450 B.n449 585
R939 B.n448 B.n9 585
R940 B.n447 B.n446 585
R941 B.n445 B.n10 585
R942 B.n444 B.n443 585
R943 B.n442 B.n11 585
R944 B.n441 B.n440 585
R945 B.n471 B.n470 585
R946 B.n152 B.n115 482.89
R947 B.n440 B.n439 482.89
R948 B.n266 B.n265 482.89
R949 B.n326 B.n53 482.89
R950 B.n90 B.t2 331.022
R951 B.n36 B.t7 331.022
R952 B.n98 B.t5 331.022
R953 B.n28 B.t10 331.022
R954 B.n91 B.t1 318.027
R955 B.n37 B.t8 318.027
R956 B.n99 B.t4 318.027
R957 B.n29 B.t11 318.027
R958 B.n152 B.n151 163.367
R959 B.n151 B.n150 163.367
R960 B.n150 B.n117 163.367
R961 B.n146 B.n117 163.367
R962 B.n146 B.n145 163.367
R963 B.n145 B.n144 163.367
R964 B.n144 B.n119 163.367
R965 B.n140 B.n119 163.367
R966 B.n140 B.n139 163.367
R967 B.n139 B.n138 163.367
R968 B.n138 B.n121 163.367
R969 B.n134 B.n121 163.367
R970 B.n134 B.n133 163.367
R971 B.n133 B.n132 163.367
R972 B.n132 B.n123 163.367
R973 B.n128 B.n123 163.367
R974 B.n128 B.n127 163.367
R975 B.n127 B.n126 163.367
R976 B.n126 B.n2 163.367
R977 B.n470 B.n2 163.367
R978 B.n470 B.n469 163.367
R979 B.n469 B.n468 163.367
R980 B.n468 B.n3 163.367
R981 B.n464 B.n3 163.367
R982 B.n464 B.n463 163.367
R983 B.n463 B.n462 163.367
R984 B.n462 B.n5 163.367
R985 B.n458 B.n5 163.367
R986 B.n458 B.n457 163.367
R987 B.n457 B.n456 163.367
R988 B.n456 B.n7 163.367
R989 B.n452 B.n7 163.367
R990 B.n452 B.n451 163.367
R991 B.n451 B.n450 163.367
R992 B.n450 B.n9 163.367
R993 B.n446 B.n9 163.367
R994 B.n446 B.n445 163.367
R995 B.n445 B.n444 163.367
R996 B.n444 B.n11 163.367
R997 B.n440 B.n11 163.367
R998 B.n156 B.n115 163.367
R999 B.n157 B.n156 163.367
R1000 B.n158 B.n157 163.367
R1001 B.n158 B.n113 163.367
R1002 B.n162 B.n113 163.367
R1003 B.n163 B.n162 163.367
R1004 B.n164 B.n163 163.367
R1005 B.n164 B.n111 163.367
R1006 B.n168 B.n111 163.367
R1007 B.n169 B.n168 163.367
R1008 B.n170 B.n169 163.367
R1009 B.n170 B.n109 163.367
R1010 B.n174 B.n109 163.367
R1011 B.n175 B.n174 163.367
R1012 B.n176 B.n175 163.367
R1013 B.n176 B.n107 163.367
R1014 B.n180 B.n107 163.367
R1015 B.n181 B.n180 163.367
R1016 B.n182 B.n181 163.367
R1017 B.n182 B.n105 163.367
R1018 B.n186 B.n105 163.367
R1019 B.n187 B.n186 163.367
R1020 B.n188 B.n187 163.367
R1021 B.n188 B.n103 163.367
R1022 B.n192 B.n103 163.367
R1023 B.n193 B.n192 163.367
R1024 B.n194 B.n193 163.367
R1025 B.n194 B.n101 163.367
R1026 B.n198 B.n101 163.367
R1027 B.n199 B.n198 163.367
R1028 B.n200 B.n199 163.367
R1029 B.n200 B.n97 163.367
R1030 B.n205 B.n97 163.367
R1031 B.n206 B.n205 163.367
R1032 B.n207 B.n206 163.367
R1033 B.n207 B.n95 163.367
R1034 B.n211 B.n95 163.367
R1035 B.n212 B.n211 163.367
R1036 B.n213 B.n212 163.367
R1037 B.n213 B.n93 163.367
R1038 B.n217 B.n93 163.367
R1039 B.n218 B.n217 163.367
R1040 B.n218 B.n89 163.367
R1041 B.n222 B.n89 163.367
R1042 B.n223 B.n222 163.367
R1043 B.n224 B.n223 163.367
R1044 B.n224 B.n87 163.367
R1045 B.n228 B.n87 163.367
R1046 B.n229 B.n228 163.367
R1047 B.n230 B.n229 163.367
R1048 B.n230 B.n85 163.367
R1049 B.n234 B.n85 163.367
R1050 B.n235 B.n234 163.367
R1051 B.n236 B.n235 163.367
R1052 B.n236 B.n83 163.367
R1053 B.n240 B.n83 163.367
R1054 B.n241 B.n240 163.367
R1055 B.n242 B.n241 163.367
R1056 B.n242 B.n81 163.367
R1057 B.n246 B.n81 163.367
R1058 B.n247 B.n246 163.367
R1059 B.n248 B.n247 163.367
R1060 B.n248 B.n79 163.367
R1061 B.n252 B.n79 163.367
R1062 B.n253 B.n252 163.367
R1063 B.n254 B.n253 163.367
R1064 B.n254 B.n77 163.367
R1065 B.n258 B.n77 163.367
R1066 B.n259 B.n258 163.367
R1067 B.n260 B.n259 163.367
R1068 B.n260 B.n75 163.367
R1069 B.n264 B.n75 163.367
R1070 B.n265 B.n264 163.367
R1071 B.n266 B.n73 163.367
R1072 B.n270 B.n73 163.367
R1073 B.n271 B.n270 163.367
R1074 B.n272 B.n271 163.367
R1075 B.n272 B.n71 163.367
R1076 B.n276 B.n71 163.367
R1077 B.n277 B.n276 163.367
R1078 B.n278 B.n277 163.367
R1079 B.n278 B.n69 163.367
R1080 B.n282 B.n69 163.367
R1081 B.n283 B.n282 163.367
R1082 B.n284 B.n283 163.367
R1083 B.n284 B.n67 163.367
R1084 B.n288 B.n67 163.367
R1085 B.n289 B.n288 163.367
R1086 B.n290 B.n289 163.367
R1087 B.n290 B.n65 163.367
R1088 B.n294 B.n65 163.367
R1089 B.n295 B.n294 163.367
R1090 B.n296 B.n295 163.367
R1091 B.n296 B.n63 163.367
R1092 B.n300 B.n63 163.367
R1093 B.n301 B.n300 163.367
R1094 B.n302 B.n301 163.367
R1095 B.n302 B.n61 163.367
R1096 B.n306 B.n61 163.367
R1097 B.n307 B.n306 163.367
R1098 B.n308 B.n307 163.367
R1099 B.n308 B.n59 163.367
R1100 B.n312 B.n59 163.367
R1101 B.n313 B.n312 163.367
R1102 B.n314 B.n313 163.367
R1103 B.n314 B.n57 163.367
R1104 B.n318 B.n57 163.367
R1105 B.n319 B.n318 163.367
R1106 B.n320 B.n319 163.367
R1107 B.n320 B.n55 163.367
R1108 B.n324 B.n55 163.367
R1109 B.n325 B.n324 163.367
R1110 B.n326 B.n325 163.367
R1111 B.n439 B.n438 163.367
R1112 B.n438 B.n13 163.367
R1113 B.n434 B.n13 163.367
R1114 B.n434 B.n433 163.367
R1115 B.n433 B.n432 163.367
R1116 B.n432 B.n15 163.367
R1117 B.n428 B.n15 163.367
R1118 B.n428 B.n427 163.367
R1119 B.n427 B.n426 163.367
R1120 B.n426 B.n17 163.367
R1121 B.n422 B.n17 163.367
R1122 B.n422 B.n421 163.367
R1123 B.n421 B.n420 163.367
R1124 B.n420 B.n19 163.367
R1125 B.n416 B.n19 163.367
R1126 B.n416 B.n415 163.367
R1127 B.n415 B.n414 163.367
R1128 B.n414 B.n21 163.367
R1129 B.n410 B.n21 163.367
R1130 B.n410 B.n409 163.367
R1131 B.n409 B.n408 163.367
R1132 B.n408 B.n23 163.367
R1133 B.n404 B.n23 163.367
R1134 B.n404 B.n403 163.367
R1135 B.n403 B.n402 163.367
R1136 B.n402 B.n25 163.367
R1137 B.n398 B.n25 163.367
R1138 B.n398 B.n397 163.367
R1139 B.n397 B.n396 163.367
R1140 B.n396 B.n27 163.367
R1141 B.n392 B.n27 163.367
R1142 B.n392 B.n391 163.367
R1143 B.n391 B.n31 163.367
R1144 B.n387 B.n31 163.367
R1145 B.n387 B.n386 163.367
R1146 B.n386 B.n385 163.367
R1147 B.n385 B.n33 163.367
R1148 B.n381 B.n33 163.367
R1149 B.n381 B.n380 163.367
R1150 B.n380 B.n379 163.367
R1151 B.n379 B.n35 163.367
R1152 B.n374 B.n35 163.367
R1153 B.n374 B.n373 163.367
R1154 B.n373 B.n372 163.367
R1155 B.n372 B.n39 163.367
R1156 B.n368 B.n39 163.367
R1157 B.n368 B.n367 163.367
R1158 B.n367 B.n366 163.367
R1159 B.n366 B.n41 163.367
R1160 B.n362 B.n41 163.367
R1161 B.n362 B.n361 163.367
R1162 B.n361 B.n360 163.367
R1163 B.n360 B.n43 163.367
R1164 B.n356 B.n43 163.367
R1165 B.n356 B.n355 163.367
R1166 B.n355 B.n354 163.367
R1167 B.n354 B.n45 163.367
R1168 B.n350 B.n45 163.367
R1169 B.n350 B.n349 163.367
R1170 B.n349 B.n348 163.367
R1171 B.n348 B.n47 163.367
R1172 B.n344 B.n47 163.367
R1173 B.n344 B.n343 163.367
R1174 B.n343 B.n342 163.367
R1175 B.n342 B.n49 163.367
R1176 B.n338 B.n49 163.367
R1177 B.n338 B.n337 163.367
R1178 B.n337 B.n336 163.367
R1179 B.n336 B.n51 163.367
R1180 B.n332 B.n51 163.367
R1181 B.n332 B.n331 163.367
R1182 B.n331 B.n330 163.367
R1183 B.n330 B.n53 163.367
R1184 B.n92 B.n91 59.5399
R1185 B.n202 B.n99 59.5399
R1186 B.n30 B.n29 59.5399
R1187 B.n376 B.n37 59.5399
R1188 B.n441 B.n12 31.3761
R1189 B.n328 B.n327 31.3761
R1190 B.n267 B.n74 31.3761
R1191 B.n154 B.n153 31.3761
R1192 B B.n471 18.0485
R1193 B.n91 B.n90 12.9944
R1194 B.n99 B.n98 12.9944
R1195 B.n29 B.n28 12.9944
R1196 B.n37 B.n36 12.9944
R1197 B.n437 B.n12 10.6151
R1198 B.n437 B.n436 10.6151
R1199 B.n436 B.n435 10.6151
R1200 B.n435 B.n14 10.6151
R1201 B.n431 B.n14 10.6151
R1202 B.n431 B.n430 10.6151
R1203 B.n430 B.n429 10.6151
R1204 B.n429 B.n16 10.6151
R1205 B.n425 B.n16 10.6151
R1206 B.n425 B.n424 10.6151
R1207 B.n424 B.n423 10.6151
R1208 B.n423 B.n18 10.6151
R1209 B.n419 B.n18 10.6151
R1210 B.n419 B.n418 10.6151
R1211 B.n418 B.n417 10.6151
R1212 B.n417 B.n20 10.6151
R1213 B.n413 B.n20 10.6151
R1214 B.n413 B.n412 10.6151
R1215 B.n412 B.n411 10.6151
R1216 B.n411 B.n22 10.6151
R1217 B.n407 B.n22 10.6151
R1218 B.n407 B.n406 10.6151
R1219 B.n406 B.n405 10.6151
R1220 B.n405 B.n24 10.6151
R1221 B.n401 B.n24 10.6151
R1222 B.n401 B.n400 10.6151
R1223 B.n400 B.n399 10.6151
R1224 B.n399 B.n26 10.6151
R1225 B.n395 B.n26 10.6151
R1226 B.n395 B.n394 10.6151
R1227 B.n394 B.n393 10.6151
R1228 B.n390 B.n389 10.6151
R1229 B.n389 B.n388 10.6151
R1230 B.n388 B.n32 10.6151
R1231 B.n384 B.n32 10.6151
R1232 B.n384 B.n383 10.6151
R1233 B.n383 B.n382 10.6151
R1234 B.n382 B.n34 10.6151
R1235 B.n378 B.n34 10.6151
R1236 B.n378 B.n377 10.6151
R1237 B.n375 B.n38 10.6151
R1238 B.n371 B.n38 10.6151
R1239 B.n371 B.n370 10.6151
R1240 B.n370 B.n369 10.6151
R1241 B.n369 B.n40 10.6151
R1242 B.n365 B.n40 10.6151
R1243 B.n365 B.n364 10.6151
R1244 B.n364 B.n363 10.6151
R1245 B.n363 B.n42 10.6151
R1246 B.n359 B.n42 10.6151
R1247 B.n359 B.n358 10.6151
R1248 B.n358 B.n357 10.6151
R1249 B.n357 B.n44 10.6151
R1250 B.n353 B.n44 10.6151
R1251 B.n353 B.n352 10.6151
R1252 B.n352 B.n351 10.6151
R1253 B.n351 B.n46 10.6151
R1254 B.n347 B.n46 10.6151
R1255 B.n347 B.n346 10.6151
R1256 B.n346 B.n345 10.6151
R1257 B.n345 B.n48 10.6151
R1258 B.n341 B.n48 10.6151
R1259 B.n341 B.n340 10.6151
R1260 B.n340 B.n339 10.6151
R1261 B.n339 B.n50 10.6151
R1262 B.n335 B.n50 10.6151
R1263 B.n335 B.n334 10.6151
R1264 B.n334 B.n333 10.6151
R1265 B.n333 B.n52 10.6151
R1266 B.n329 B.n52 10.6151
R1267 B.n329 B.n328 10.6151
R1268 B.n268 B.n267 10.6151
R1269 B.n269 B.n268 10.6151
R1270 B.n269 B.n72 10.6151
R1271 B.n273 B.n72 10.6151
R1272 B.n274 B.n273 10.6151
R1273 B.n275 B.n274 10.6151
R1274 B.n275 B.n70 10.6151
R1275 B.n279 B.n70 10.6151
R1276 B.n280 B.n279 10.6151
R1277 B.n281 B.n280 10.6151
R1278 B.n281 B.n68 10.6151
R1279 B.n285 B.n68 10.6151
R1280 B.n286 B.n285 10.6151
R1281 B.n287 B.n286 10.6151
R1282 B.n287 B.n66 10.6151
R1283 B.n291 B.n66 10.6151
R1284 B.n292 B.n291 10.6151
R1285 B.n293 B.n292 10.6151
R1286 B.n293 B.n64 10.6151
R1287 B.n297 B.n64 10.6151
R1288 B.n298 B.n297 10.6151
R1289 B.n299 B.n298 10.6151
R1290 B.n299 B.n62 10.6151
R1291 B.n303 B.n62 10.6151
R1292 B.n304 B.n303 10.6151
R1293 B.n305 B.n304 10.6151
R1294 B.n305 B.n60 10.6151
R1295 B.n309 B.n60 10.6151
R1296 B.n310 B.n309 10.6151
R1297 B.n311 B.n310 10.6151
R1298 B.n311 B.n58 10.6151
R1299 B.n315 B.n58 10.6151
R1300 B.n316 B.n315 10.6151
R1301 B.n317 B.n316 10.6151
R1302 B.n317 B.n56 10.6151
R1303 B.n321 B.n56 10.6151
R1304 B.n322 B.n321 10.6151
R1305 B.n323 B.n322 10.6151
R1306 B.n323 B.n54 10.6151
R1307 B.n327 B.n54 10.6151
R1308 B.n155 B.n154 10.6151
R1309 B.n155 B.n114 10.6151
R1310 B.n159 B.n114 10.6151
R1311 B.n160 B.n159 10.6151
R1312 B.n161 B.n160 10.6151
R1313 B.n161 B.n112 10.6151
R1314 B.n165 B.n112 10.6151
R1315 B.n166 B.n165 10.6151
R1316 B.n167 B.n166 10.6151
R1317 B.n167 B.n110 10.6151
R1318 B.n171 B.n110 10.6151
R1319 B.n172 B.n171 10.6151
R1320 B.n173 B.n172 10.6151
R1321 B.n173 B.n108 10.6151
R1322 B.n177 B.n108 10.6151
R1323 B.n178 B.n177 10.6151
R1324 B.n179 B.n178 10.6151
R1325 B.n179 B.n106 10.6151
R1326 B.n183 B.n106 10.6151
R1327 B.n184 B.n183 10.6151
R1328 B.n185 B.n184 10.6151
R1329 B.n185 B.n104 10.6151
R1330 B.n189 B.n104 10.6151
R1331 B.n190 B.n189 10.6151
R1332 B.n191 B.n190 10.6151
R1333 B.n191 B.n102 10.6151
R1334 B.n195 B.n102 10.6151
R1335 B.n196 B.n195 10.6151
R1336 B.n197 B.n196 10.6151
R1337 B.n197 B.n100 10.6151
R1338 B.n201 B.n100 10.6151
R1339 B.n204 B.n203 10.6151
R1340 B.n204 B.n96 10.6151
R1341 B.n208 B.n96 10.6151
R1342 B.n209 B.n208 10.6151
R1343 B.n210 B.n209 10.6151
R1344 B.n210 B.n94 10.6151
R1345 B.n214 B.n94 10.6151
R1346 B.n215 B.n214 10.6151
R1347 B.n216 B.n215 10.6151
R1348 B.n220 B.n219 10.6151
R1349 B.n221 B.n220 10.6151
R1350 B.n221 B.n88 10.6151
R1351 B.n225 B.n88 10.6151
R1352 B.n226 B.n225 10.6151
R1353 B.n227 B.n226 10.6151
R1354 B.n227 B.n86 10.6151
R1355 B.n231 B.n86 10.6151
R1356 B.n232 B.n231 10.6151
R1357 B.n233 B.n232 10.6151
R1358 B.n233 B.n84 10.6151
R1359 B.n237 B.n84 10.6151
R1360 B.n238 B.n237 10.6151
R1361 B.n239 B.n238 10.6151
R1362 B.n239 B.n82 10.6151
R1363 B.n243 B.n82 10.6151
R1364 B.n244 B.n243 10.6151
R1365 B.n245 B.n244 10.6151
R1366 B.n245 B.n80 10.6151
R1367 B.n249 B.n80 10.6151
R1368 B.n250 B.n249 10.6151
R1369 B.n251 B.n250 10.6151
R1370 B.n251 B.n78 10.6151
R1371 B.n255 B.n78 10.6151
R1372 B.n256 B.n255 10.6151
R1373 B.n257 B.n256 10.6151
R1374 B.n257 B.n76 10.6151
R1375 B.n261 B.n76 10.6151
R1376 B.n262 B.n261 10.6151
R1377 B.n263 B.n262 10.6151
R1378 B.n263 B.n74 10.6151
R1379 B.n153 B.n116 10.6151
R1380 B.n149 B.n116 10.6151
R1381 B.n149 B.n148 10.6151
R1382 B.n148 B.n147 10.6151
R1383 B.n147 B.n118 10.6151
R1384 B.n143 B.n118 10.6151
R1385 B.n143 B.n142 10.6151
R1386 B.n142 B.n141 10.6151
R1387 B.n141 B.n120 10.6151
R1388 B.n137 B.n120 10.6151
R1389 B.n137 B.n136 10.6151
R1390 B.n136 B.n135 10.6151
R1391 B.n135 B.n122 10.6151
R1392 B.n131 B.n122 10.6151
R1393 B.n131 B.n130 10.6151
R1394 B.n130 B.n129 10.6151
R1395 B.n129 B.n124 10.6151
R1396 B.n125 B.n124 10.6151
R1397 B.n125 B.n0 10.6151
R1398 B.n467 B.n1 10.6151
R1399 B.n467 B.n466 10.6151
R1400 B.n466 B.n465 10.6151
R1401 B.n465 B.n4 10.6151
R1402 B.n461 B.n4 10.6151
R1403 B.n461 B.n460 10.6151
R1404 B.n460 B.n459 10.6151
R1405 B.n459 B.n6 10.6151
R1406 B.n455 B.n6 10.6151
R1407 B.n455 B.n454 10.6151
R1408 B.n454 B.n453 10.6151
R1409 B.n453 B.n8 10.6151
R1410 B.n449 B.n8 10.6151
R1411 B.n449 B.n448 10.6151
R1412 B.n448 B.n447 10.6151
R1413 B.n447 B.n10 10.6151
R1414 B.n443 B.n10 10.6151
R1415 B.n443 B.n442 10.6151
R1416 B.n442 B.n441 10.6151
R1417 B.n393 B.n30 9.36635
R1418 B.n376 B.n375 9.36635
R1419 B.n202 B.n201 9.36635
R1420 B.n219 B.n92 9.36635
R1421 B.n471 B.n0 2.81026
R1422 B.n471 B.n1 2.81026
R1423 B.n390 B.n30 1.24928
R1424 B.n377 B.n376 1.24928
R1425 B.n203 B.n202 1.24928
R1426 B.n216 B.n92 1.24928
C0 w_n1774_n2726# VDD1 1.632f
C1 VP VN 4.46933f
C2 B VN 0.666911f
C3 VTAIL VDD2 15.0762f
C4 B VP 1.0311f
C5 VDD1 VN 0.148017f
C6 w_n1774_n2726# VDD2 1.65812f
C7 VDD1 VP 3.41732f
C8 B VDD1 1.31676f
C9 w_n1774_n2726# VTAIL 2.51547f
C10 VDD2 VN 3.27405f
C11 VP VDD2 0.29511f
C12 B VDD2 1.34728f
C13 VTAIL VN 3.03991f
C14 VTAIL VP 3.05448f
C15 B VTAIL 1.94694f
C16 VDD1 VDD2 0.747969f
C17 w_n1774_n2726# VN 3.04142f
C18 w_n1774_n2726# VP 3.26541f
C19 B w_n1774_n2726# 5.85315f
C20 VDD1 VTAIL 15.043799f
C21 VDD2 VSUBS 1.287449f
C22 VDD1 VSUBS 0.927349f
C23 VTAIL VSUBS 0.532772f
C24 VN VSUBS 4.35535f
C25 VP VSUBS 1.259441f
C26 B VSUBS 2.282908f
C27 w_n1774_n2726# VSUBS 59.883102f
C28 B.n0 VSUBS 0.00388f
C29 B.n1 VSUBS 0.00388f
C30 B.n2 VSUBS 0.006136f
C31 B.n3 VSUBS 0.006136f
C32 B.n4 VSUBS 0.006136f
C33 B.n5 VSUBS 0.006136f
C34 B.n6 VSUBS 0.006136f
C35 B.n7 VSUBS 0.006136f
C36 B.n8 VSUBS 0.006136f
C37 B.n9 VSUBS 0.006136f
C38 B.n10 VSUBS 0.006136f
C39 B.n11 VSUBS 0.006136f
C40 B.n12 VSUBS 0.014327f
C41 B.n13 VSUBS 0.006136f
C42 B.n14 VSUBS 0.006136f
C43 B.n15 VSUBS 0.006136f
C44 B.n16 VSUBS 0.006136f
C45 B.n17 VSUBS 0.006136f
C46 B.n18 VSUBS 0.006136f
C47 B.n19 VSUBS 0.006136f
C48 B.n20 VSUBS 0.006136f
C49 B.n21 VSUBS 0.006136f
C50 B.n22 VSUBS 0.006136f
C51 B.n23 VSUBS 0.006136f
C52 B.n24 VSUBS 0.006136f
C53 B.n25 VSUBS 0.006136f
C54 B.n26 VSUBS 0.006136f
C55 B.n27 VSUBS 0.006136f
C56 B.t11 VSUBS 0.125028f
C57 B.t10 VSUBS 0.131388f
C58 B.t9 VSUBS 0.105052f
C59 B.n28 VSUBS 0.191813f
C60 B.n29 VSUBS 0.170766f
C61 B.n30 VSUBS 0.014217f
C62 B.n31 VSUBS 0.006136f
C63 B.n32 VSUBS 0.006136f
C64 B.n33 VSUBS 0.006136f
C65 B.n34 VSUBS 0.006136f
C66 B.n35 VSUBS 0.006136f
C67 B.t8 VSUBS 0.12503f
C68 B.t7 VSUBS 0.13139f
C69 B.t6 VSUBS 0.105052f
C70 B.n36 VSUBS 0.191811f
C71 B.n37 VSUBS 0.170764f
C72 B.n38 VSUBS 0.006136f
C73 B.n39 VSUBS 0.006136f
C74 B.n40 VSUBS 0.006136f
C75 B.n41 VSUBS 0.006136f
C76 B.n42 VSUBS 0.006136f
C77 B.n43 VSUBS 0.006136f
C78 B.n44 VSUBS 0.006136f
C79 B.n45 VSUBS 0.006136f
C80 B.n46 VSUBS 0.006136f
C81 B.n47 VSUBS 0.006136f
C82 B.n48 VSUBS 0.006136f
C83 B.n49 VSUBS 0.006136f
C84 B.n50 VSUBS 0.006136f
C85 B.n51 VSUBS 0.006136f
C86 B.n52 VSUBS 0.006136f
C87 B.n53 VSUBS 0.014327f
C88 B.n54 VSUBS 0.006136f
C89 B.n55 VSUBS 0.006136f
C90 B.n56 VSUBS 0.006136f
C91 B.n57 VSUBS 0.006136f
C92 B.n58 VSUBS 0.006136f
C93 B.n59 VSUBS 0.006136f
C94 B.n60 VSUBS 0.006136f
C95 B.n61 VSUBS 0.006136f
C96 B.n62 VSUBS 0.006136f
C97 B.n63 VSUBS 0.006136f
C98 B.n64 VSUBS 0.006136f
C99 B.n65 VSUBS 0.006136f
C100 B.n66 VSUBS 0.006136f
C101 B.n67 VSUBS 0.006136f
C102 B.n68 VSUBS 0.006136f
C103 B.n69 VSUBS 0.006136f
C104 B.n70 VSUBS 0.006136f
C105 B.n71 VSUBS 0.006136f
C106 B.n72 VSUBS 0.006136f
C107 B.n73 VSUBS 0.006136f
C108 B.n74 VSUBS 0.014327f
C109 B.n75 VSUBS 0.006136f
C110 B.n76 VSUBS 0.006136f
C111 B.n77 VSUBS 0.006136f
C112 B.n78 VSUBS 0.006136f
C113 B.n79 VSUBS 0.006136f
C114 B.n80 VSUBS 0.006136f
C115 B.n81 VSUBS 0.006136f
C116 B.n82 VSUBS 0.006136f
C117 B.n83 VSUBS 0.006136f
C118 B.n84 VSUBS 0.006136f
C119 B.n85 VSUBS 0.006136f
C120 B.n86 VSUBS 0.006136f
C121 B.n87 VSUBS 0.006136f
C122 B.n88 VSUBS 0.006136f
C123 B.n89 VSUBS 0.006136f
C124 B.t1 VSUBS 0.12503f
C125 B.t2 VSUBS 0.13139f
C126 B.t0 VSUBS 0.105052f
C127 B.n90 VSUBS 0.191811f
C128 B.n91 VSUBS 0.170764f
C129 B.n92 VSUBS 0.014217f
C130 B.n93 VSUBS 0.006136f
C131 B.n94 VSUBS 0.006136f
C132 B.n95 VSUBS 0.006136f
C133 B.n96 VSUBS 0.006136f
C134 B.n97 VSUBS 0.006136f
C135 B.t4 VSUBS 0.125028f
C136 B.t5 VSUBS 0.131388f
C137 B.t3 VSUBS 0.105052f
C138 B.n98 VSUBS 0.191813f
C139 B.n99 VSUBS 0.170766f
C140 B.n100 VSUBS 0.006136f
C141 B.n101 VSUBS 0.006136f
C142 B.n102 VSUBS 0.006136f
C143 B.n103 VSUBS 0.006136f
C144 B.n104 VSUBS 0.006136f
C145 B.n105 VSUBS 0.006136f
C146 B.n106 VSUBS 0.006136f
C147 B.n107 VSUBS 0.006136f
C148 B.n108 VSUBS 0.006136f
C149 B.n109 VSUBS 0.006136f
C150 B.n110 VSUBS 0.006136f
C151 B.n111 VSUBS 0.006136f
C152 B.n112 VSUBS 0.006136f
C153 B.n113 VSUBS 0.006136f
C154 B.n114 VSUBS 0.006136f
C155 B.n115 VSUBS 0.014327f
C156 B.n116 VSUBS 0.006136f
C157 B.n117 VSUBS 0.006136f
C158 B.n118 VSUBS 0.006136f
C159 B.n119 VSUBS 0.006136f
C160 B.n120 VSUBS 0.006136f
C161 B.n121 VSUBS 0.006136f
C162 B.n122 VSUBS 0.006136f
C163 B.n123 VSUBS 0.006136f
C164 B.n124 VSUBS 0.006136f
C165 B.n125 VSUBS 0.006136f
C166 B.n126 VSUBS 0.006136f
C167 B.n127 VSUBS 0.006136f
C168 B.n128 VSUBS 0.006136f
C169 B.n129 VSUBS 0.006136f
C170 B.n130 VSUBS 0.006136f
C171 B.n131 VSUBS 0.006136f
C172 B.n132 VSUBS 0.006136f
C173 B.n133 VSUBS 0.006136f
C174 B.n134 VSUBS 0.006136f
C175 B.n135 VSUBS 0.006136f
C176 B.n136 VSUBS 0.006136f
C177 B.n137 VSUBS 0.006136f
C178 B.n138 VSUBS 0.006136f
C179 B.n139 VSUBS 0.006136f
C180 B.n140 VSUBS 0.006136f
C181 B.n141 VSUBS 0.006136f
C182 B.n142 VSUBS 0.006136f
C183 B.n143 VSUBS 0.006136f
C184 B.n144 VSUBS 0.006136f
C185 B.n145 VSUBS 0.006136f
C186 B.n146 VSUBS 0.006136f
C187 B.n147 VSUBS 0.006136f
C188 B.n148 VSUBS 0.006136f
C189 B.n149 VSUBS 0.006136f
C190 B.n150 VSUBS 0.006136f
C191 B.n151 VSUBS 0.006136f
C192 B.n152 VSUBS 0.013646f
C193 B.n153 VSUBS 0.013646f
C194 B.n154 VSUBS 0.014327f
C195 B.n155 VSUBS 0.006136f
C196 B.n156 VSUBS 0.006136f
C197 B.n157 VSUBS 0.006136f
C198 B.n158 VSUBS 0.006136f
C199 B.n159 VSUBS 0.006136f
C200 B.n160 VSUBS 0.006136f
C201 B.n161 VSUBS 0.006136f
C202 B.n162 VSUBS 0.006136f
C203 B.n163 VSUBS 0.006136f
C204 B.n164 VSUBS 0.006136f
C205 B.n165 VSUBS 0.006136f
C206 B.n166 VSUBS 0.006136f
C207 B.n167 VSUBS 0.006136f
C208 B.n168 VSUBS 0.006136f
C209 B.n169 VSUBS 0.006136f
C210 B.n170 VSUBS 0.006136f
C211 B.n171 VSUBS 0.006136f
C212 B.n172 VSUBS 0.006136f
C213 B.n173 VSUBS 0.006136f
C214 B.n174 VSUBS 0.006136f
C215 B.n175 VSUBS 0.006136f
C216 B.n176 VSUBS 0.006136f
C217 B.n177 VSUBS 0.006136f
C218 B.n178 VSUBS 0.006136f
C219 B.n179 VSUBS 0.006136f
C220 B.n180 VSUBS 0.006136f
C221 B.n181 VSUBS 0.006136f
C222 B.n182 VSUBS 0.006136f
C223 B.n183 VSUBS 0.006136f
C224 B.n184 VSUBS 0.006136f
C225 B.n185 VSUBS 0.006136f
C226 B.n186 VSUBS 0.006136f
C227 B.n187 VSUBS 0.006136f
C228 B.n188 VSUBS 0.006136f
C229 B.n189 VSUBS 0.006136f
C230 B.n190 VSUBS 0.006136f
C231 B.n191 VSUBS 0.006136f
C232 B.n192 VSUBS 0.006136f
C233 B.n193 VSUBS 0.006136f
C234 B.n194 VSUBS 0.006136f
C235 B.n195 VSUBS 0.006136f
C236 B.n196 VSUBS 0.006136f
C237 B.n197 VSUBS 0.006136f
C238 B.n198 VSUBS 0.006136f
C239 B.n199 VSUBS 0.006136f
C240 B.n200 VSUBS 0.006136f
C241 B.n201 VSUBS 0.005775f
C242 B.n202 VSUBS 0.014217f
C243 B.n203 VSUBS 0.003429f
C244 B.n204 VSUBS 0.006136f
C245 B.n205 VSUBS 0.006136f
C246 B.n206 VSUBS 0.006136f
C247 B.n207 VSUBS 0.006136f
C248 B.n208 VSUBS 0.006136f
C249 B.n209 VSUBS 0.006136f
C250 B.n210 VSUBS 0.006136f
C251 B.n211 VSUBS 0.006136f
C252 B.n212 VSUBS 0.006136f
C253 B.n213 VSUBS 0.006136f
C254 B.n214 VSUBS 0.006136f
C255 B.n215 VSUBS 0.006136f
C256 B.n216 VSUBS 0.003429f
C257 B.n217 VSUBS 0.006136f
C258 B.n218 VSUBS 0.006136f
C259 B.n219 VSUBS 0.005775f
C260 B.n220 VSUBS 0.006136f
C261 B.n221 VSUBS 0.006136f
C262 B.n222 VSUBS 0.006136f
C263 B.n223 VSUBS 0.006136f
C264 B.n224 VSUBS 0.006136f
C265 B.n225 VSUBS 0.006136f
C266 B.n226 VSUBS 0.006136f
C267 B.n227 VSUBS 0.006136f
C268 B.n228 VSUBS 0.006136f
C269 B.n229 VSUBS 0.006136f
C270 B.n230 VSUBS 0.006136f
C271 B.n231 VSUBS 0.006136f
C272 B.n232 VSUBS 0.006136f
C273 B.n233 VSUBS 0.006136f
C274 B.n234 VSUBS 0.006136f
C275 B.n235 VSUBS 0.006136f
C276 B.n236 VSUBS 0.006136f
C277 B.n237 VSUBS 0.006136f
C278 B.n238 VSUBS 0.006136f
C279 B.n239 VSUBS 0.006136f
C280 B.n240 VSUBS 0.006136f
C281 B.n241 VSUBS 0.006136f
C282 B.n242 VSUBS 0.006136f
C283 B.n243 VSUBS 0.006136f
C284 B.n244 VSUBS 0.006136f
C285 B.n245 VSUBS 0.006136f
C286 B.n246 VSUBS 0.006136f
C287 B.n247 VSUBS 0.006136f
C288 B.n248 VSUBS 0.006136f
C289 B.n249 VSUBS 0.006136f
C290 B.n250 VSUBS 0.006136f
C291 B.n251 VSUBS 0.006136f
C292 B.n252 VSUBS 0.006136f
C293 B.n253 VSUBS 0.006136f
C294 B.n254 VSUBS 0.006136f
C295 B.n255 VSUBS 0.006136f
C296 B.n256 VSUBS 0.006136f
C297 B.n257 VSUBS 0.006136f
C298 B.n258 VSUBS 0.006136f
C299 B.n259 VSUBS 0.006136f
C300 B.n260 VSUBS 0.006136f
C301 B.n261 VSUBS 0.006136f
C302 B.n262 VSUBS 0.006136f
C303 B.n263 VSUBS 0.006136f
C304 B.n264 VSUBS 0.006136f
C305 B.n265 VSUBS 0.014327f
C306 B.n266 VSUBS 0.013646f
C307 B.n267 VSUBS 0.013646f
C308 B.n268 VSUBS 0.006136f
C309 B.n269 VSUBS 0.006136f
C310 B.n270 VSUBS 0.006136f
C311 B.n271 VSUBS 0.006136f
C312 B.n272 VSUBS 0.006136f
C313 B.n273 VSUBS 0.006136f
C314 B.n274 VSUBS 0.006136f
C315 B.n275 VSUBS 0.006136f
C316 B.n276 VSUBS 0.006136f
C317 B.n277 VSUBS 0.006136f
C318 B.n278 VSUBS 0.006136f
C319 B.n279 VSUBS 0.006136f
C320 B.n280 VSUBS 0.006136f
C321 B.n281 VSUBS 0.006136f
C322 B.n282 VSUBS 0.006136f
C323 B.n283 VSUBS 0.006136f
C324 B.n284 VSUBS 0.006136f
C325 B.n285 VSUBS 0.006136f
C326 B.n286 VSUBS 0.006136f
C327 B.n287 VSUBS 0.006136f
C328 B.n288 VSUBS 0.006136f
C329 B.n289 VSUBS 0.006136f
C330 B.n290 VSUBS 0.006136f
C331 B.n291 VSUBS 0.006136f
C332 B.n292 VSUBS 0.006136f
C333 B.n293 VSUBS 0.006136f
C334 B.n294 VSUBS 0.006136f
C335 B.n295 VSUBS 0.006136f
C336 B.n296 VSUBS 0.006136f
C337 B.n297 VSUBS 0.006136f
C338 B.n298 VSUBS 0.006136f
C339 B.n299 VSUBS 0.006136f
C340 B.n300 VSUBS 0.006136f
C341 B.n301 VSUBS 0.006136f
C342 B.n302 VSUBS 0.006136f
C343 B.n303 VSUBS 0.006136f
C344 B.n304 VSUBS 0.006136f
C345 B.n305 VSUBS 0.006136f
C346 B.n306 VSUBS 0.006136f
C347 B.n307 VSUBS 0.006136f
C348 B.n308 VSUBS 0.006136f
C349 B.n309 VSUBS 0.006136f
C350 B.n310 VSUBS 0.006136f
C351 B.n311 VSUBS 0.006136f
C352 B.n312 VSUBS 0.006136f
C353 B.n313 VSUBS 0.006136f
C354 B.n314 VSUBS 0.006136f
C355 B.n315 VSUBS 0.006136f
C356 B.n316 VSUBS 0.006136f
C357 B.n317 VSUBS 0.006136f
C358 B.n318 VSUBS 0.006136f
C359 B.n319 VSUBS 0.006136f
C360 B.n320 VSUBS 0.006136f
C361 B.n321 VSUBS 0.006136f
C362 B.n322 VSUBS 0.006136f
C363 B.n323 VSUBS 0.006136f
C364 B.n324 VSUBS 0.006136f
C365 B.n325 VSUBS 0.006136f
C366 B.n326 VSUBS 0.013646f
C367 B.n327 VSUBS 0.014401f
C368 B.n328 VSUBS 0.013573f
C369 B.n329 VSUBS 0.006136f
C370 B.n330 VSUBS 0.006136f
C371 B.n331 VSUBS 0.006136f
C372 B.n332 VSUBS 0.006136f
C373 B.n333 VSUBS 0.006136f
C374 B.n334 VSUBS 0.006136f
C375 B.n335 VSUBS 0.006136f
C376 B.n336 VSUBS 0.006136f
C377 B.n337 VSUBS 0.006136f
C378 B.n338 VSUBS 0.006136f
C379 B.n339 VSUBS 0.006136f
C380 B.n340 VSUBS 0.006136f
C381 B.n341 VSUBS 0.006136f
C382 B.n342 VSUBS 0.006136f
C383 B.n343 VSUBS 0.006136f
C384 B.n344 VSUBS 0.006136f
C385 B.n345 VSUBS 0.006136f
C386 B.n346 VSUBS 0.006136f
C387 B.n347 VSUBS 0.006136f
C388 B.n348 VSUBS 0.006136f
C389 B.n349 VSUBS 0.006136f
C390 B.n350 VSUBS 0.006136f
C391 B.n351 VSUBS 0.006136f
C392 B.n352 VSUBS 0.006136f
C393 B.n353 VSUBS 0.006136f
C394 B.n354 VSUBS 0.006136f
C395 B.n355 VSUBS 0.006136f
C396 B.n356 VSUBS 0.006136f
C397 B.n357 VSUBS 0.006136f
C398 B.n358 VSUBS 0.006136f
C399 B.n359 VSUBS 0.006136f
C400 B.n360 VSUBS 0.006136f
C401 B.n361 VSUBS 0.006136f
C402 B.n362 VSUBS 0.006136f
C403 B.n363 VSUBS 0.006136f
C404 B.n364 VSUBS 0.006136f
C405 B.n365 VSUBS 0.006136f
C406 B.n366 VSUBS 0.006136f
C407 B.n367 VSUBS 0.006136f
C408 B.n368 VSUBS 0.006136f
C409 B.n369 VSUBS 0.006136f
C410 B.n370 VSUBS 0.006136f
C411 B.n371 VSUBS 0.006136f
C412 B.n372 VSUBS 0.006136f
C413 B.n373 VSUBS 0.006136f
C414 B.n374 VSUBS 0.006136f
C415 B.n375 VSUBS 0.005775f
C416 B.n376 VSUBS 0.014217f
C417 B.n377 VSUBS 0.003429f
C418 B.n378 VSUBS 0.006136f
C419 B.n379 VSUBS 0.006136f
C420 B.n380 VSUBS 0.006136f
C421 B.n381 VSUBS 0.006136f
C422 B.n382 VSUBS 0.006136f
C423 B.n383 VSUBS 0.006136f
C424 B.n384 VSUBS 0.006136f
C425 B.n385 VSUBS 0.006136f
C426 B.n386 VSUBS 0.006136f
C427 B.n387 VSUBS 0.006136f
C428 B.n388 VSUBS 0.006136f
C429 B.n389 VSUBS 0.006136f
C430 B.n390 VSUBS 0.003429f
C431 B.n391 VSUBS 0.006136f
C432 B.n392 VSUBS 0.006136f
C433 B.n393 VSUBS 0.005775f
C434 B.n394 VSUBS 0.006136f
C435 B.n395 VSUBS 0.006136f
C436 B.n396 VSUBS 0.006136f
C437 B.n397 VSUBS 0.006136f
C438 B.n398 VSUBS 0.006136f
C439 B.n399 VSUBS 0.006136f
C440 B.n400 VSUBS 0.006136f
C441 B.n401 VSUBS 0.006136f
C442 B.n402 VSUBS 0.006136f
C443 B.n403 VSUBS 0.006136f
C444 B.n404 VSUBS 0.006136f
C445 B.n405 VSUBS 0.006136f
C446 B.n406 VSUBS 0.006136f
C447 B.n407 VSUBS 0.006136f
C448 B.n408 VSUBS 0.006136f
C449 B.n409 VSUBS 0.006136f
C450 B.n410 VSUBS 0.006136f
C451 B.n411 VSUBS 0.006136f
C452 B.n412 VSUBS 0.006136f
C453 B.n413 VSUBS 0.006136f
C454 B.n414 VSUBS 0.006136f
C455 B.n415 VSUBS 0.006136f
C456 B.n416 VSUBS 0.006136f
C457 B.n417 VSUBS 0.006136f
C458 B.n418 VSUBS 0.006136f
C459 B.n419 VSUBS 0.006136f
C460 B.n420 VSUBS 0.006136f
C461 B.n421 VSUBS 0.006136f
C462 B.n422 VSUBS 0.006136f
C463 B.n423 VSUBS 0.006136f
C464 B.n424 VSUBS 0.006136f
C465 B.n425 VSUBS 0.006136f
C466 B.n426 VSUBS 0.006136f
C467 B.n427 VSUBS 0.006136f
C468 B.n428 VSUBS 0.006136f
C469 B.n429 VSUBS 0.006136f
C470 B.n430 VSUBS 0.006136f
C471 B.n431 VSUBS 0.006136f
C472 B.n432 VSUBS 0.006136f
C473 B.n433 VSUBS 0.006136f
C474 B.n434 VSUBS 0.006136f
C475 B.n435 VSUBS 0.006136f
C476 B.n436 VSUBS 0.006136f
C477 B.n437 VSUBS 0.006136f
C478 B.n438 VSUBS 0.006136f
C479 B.n439 VSUBS 0.014327f
C480 B.n440 VSUBS 0.013646f
C481 B.n441 VSUBS 0.013646f
C482 B.n442 VSUBS 0.006136f
C483 B.n443 VSUBS 0.006136f
C484 B.n444 VSUBS 0.006136f
C485 B.n445 VSUBS 0.006136f
C486 B.n446 VSUBS 0.006136f
C487 B.n447 VSUBS 0.006136f
C488 B.n448 VSUBS 0.006136f
C489 B.n449 VSUBS 0.006136f
C490 B.n450 VSUBS 0.006136f
C491 B.n451 VSUBS 0.006136f
C492 B.n452 VSUBS 0.006136f
C493 B.n453 VSUBS 0.006136f
C494 B.n454 VSUBS 0.006136f
C495 B.n455 VSUBS 0.006136f
C496 B.n456 VSUBS 0.006136f
C497 B.n457 VSUBS 0.006136f
C498 B.n458 VSUBS 0.006136f
C499 B.n459 VSUBS 0.006136f
C500 B.n460 VSUBS 0.006136f
C501 B.n461 VSUBS 0.006136f
C502 B.n462 VSUBS 0.006136f
C503 B.n463 VSUBS 0.006136f
C504 B.n464 VSUBS 0.006136f
C505 B.n465 VSUBS 0.006136f
C506 B.n466 VSUBS 0.006136f
C507 B.n467 VSUBS 0.006136f
C508 B.n468 VSUBS 0.006136f
C509 B.n469 VSUBS 0.006136f
C510 B.n470 VSUBS 0.006136f
C511 B.n471 VSUBS 0.013894f
C512 VDD2.n0 VSUBS 0.032359f
C513 VDD2.n1 VSUBS 0.028782f
C514 VDD2.n2 VSUBS 0.015466f
C515 VDD2.n3 VSUBS 0.036556f
C516 VDD2.n4 VSUBS 0.016376f
C517 VDD2.n5 VSUBS 0.028782f
C518 VDD2.n6 VSUBS 0.015466f
C519 VDD2.n7 VSUBS 0.036556f
C520 VDD2.n8 VSUBS 0.016376f
C521 VDD2.n9 VSUBS 0.028782f
C522 VDD2.n10 VSUBS 0.015466f
C523 VDD2.n11 VSUBS 0.036556f
C524 VDD2.n12 VSUBS 0.016376f
C525 VDD2.n13 VSUBS 1.02615f
C526 VDD2.n14 VSUBS 0.015466f
C527 VDD2.t1 VSUBS 0.07793f
C528 VDD2.n15 VSUBS 0.150282f
C529 VDD2.n16 VSUBS 0.023255f
C530 VDD2.n17 VSUBS 0.027417f
C531 VDD2.n18 VSUBS 0.036556f
C532 VDD2.n19 VSUBS 0.016376f
C533 VDD2.n20 VSUBS 0.015466f
C534 VDD2.n21 VSUBS 0.028782f
C535 VDD2.n22 VSUBS 0.028782f
C536 VDD2.n23 VSUBS 0.015466f
C537 VDD2.n24 VSUBS 0.016376f
C538 VDD2.n25 VSUBS 0.036556f
C539 VDD2.n26 VSUBS 0.036556f
C540 VDD2.n27 VSUBS 0.016376f
C541 VDD2.n28 VSUBS 0.015466f
C542 VDD2.n29 VSUBS 0.028782f
C543 VDD2.n30 VSUBS 0.028782f
C544 VDD2.n31 VSUBS 0.015466f
C545 VDD2.n32 VSUBS 0.016376f
C546 VDD2.n33 VSUBS 0.036556f
C547 VDD2.n34 VSUBS 0.036556f
C548 VDD2.n35 VSUBS 0.016376f
C549 VDD2.n36 VSUBS 0.015466f
C550 VDD2.n37 VSUBS 0.028782f
C551 VDD2.n38 VSUBS 0.028782f
C552 VDD2.n39 VSUBS 0.015466f
C553 VDD2.n40 VSUBS 0.016376f
C554 VDD2.n41 VSUBS 0.036556f
C555 VDD2.n42 VSUBS 0.090998f
C556 VDD2.n43 VSUBS 0.016376f
C557 VDD2.n44 VSUBS 0.015466f
C558 VDD2.n45 VSUBS 0.062989f
C559 VDD2.n46 VSUBS 0.06696f
C560 VDD2.t5 VSUBS 0.199923f
C561 VDD2.t6 VSUBS 0.199923f
C562 VDD2.n47 VSUBS 1.45137f
C563 VDD2.n48 VSUBS 0.699156f
C564 VDD2.t2 VSUBS 0.199923f
C565 VDD2.t3 VSUBS 0.199923f
C566 VDD2.n49 VSUBS 1.45435f
C567 VDD2.n50 VSUBS 2.03211f
C568 VDD2.n51 VSUBS 0.032359f
C569 VDD2.n52 VSUBS 0.028782f
C570 VDD2.n53 VSUBS 0.015466f
C571 VDD2.n54 VSUBS 0.036556f
C572 VDD2.n55 VSUBS 0.016376f
C573 VDD2.n56 VSUBS 0.028782f
C574 VDD2.n57 VSUBS 0.015466f
C575 VDD2.n58 VSUBS 0.036556f
C576 VDD2.n59 VSUBS 0.016376f
C577 VDD2.n60 VSUBS 0.028782f
C578 VDD2.n61 VSUBS 0.015466f
C579 VDD2.n62 VSUBS 0.036556f
C580 VDD2.n63 VSUBS 0.016376f
C581 VDD2.n64 VSUBS 1.02615f
C582 VDD2.n65 VSUBS 0.015466f
C583 VDD2.t8 VSUBS 0.07793f
C584 VDD2.n66 VSUBS 0.150282f
C585 VDD2.n67 VSUBS 0.023255f
C586 VDD2.n68 VSUBS 0.027417f
C587 VDD2.n69 VSUBS 0.036556f
C588 VDD2.n70 VSUBS 0.016376f
C589 VDD2.n71 VSUBS 0.015466f
C590 VDD2.n72 VSUBS 0.028782f
C591 VDD2.n73 VSUBS 0.028782f
C592 VDD2.n74 VSUBS 0.015466f
C593 VDD2.n75 VSUBS 0.016376f
C594 VDD2.n76 VSUBS 0.036556f
C595 VDD2.n77 VSUBS 0.036556f
C596 VDD2.n78 VSUBS 0.016376f
C597 VDD2.n79 VSUBS 0.015466f
C598 VDD2.n80 VSUBS 0.028782f
C599 VDD2.n81 VSUBS 0.028782f
C600 VDD2.n82 VSUBS 0.015466f
C601 VDD2.n83 VSUBS 0.016376f
C602 VDD2.n84 VSUBS 0.036556f
C603 VDD2.n85 VSUBS 0.036556f
C604 VDD2.n86 VSUBS 0.016376f
C605 VDD2.n87 VSUBS 0.015466f
C606 VDD2.n88 VSUBS 0.028782f
C607 VDD2.n89 VSUBS 0.028782f
C608 VDD2.n90 VSUBS 0.015466f
C609 VDD2.n91 VSUBS 0.016376f
C610 VDD2.n92 VSUBS 0.036556f
C611 VDD2.n93 VSUBS 0.090998f
C612 VDD2.n94 VSUBS 0.016376f
C613 VDD2.n95 VSUBS 0.015466f
C614 VDD2.n96 VSUBS 0.062989f
C615 VDD2.n97 VSUBS 0.065665f
C616 VDD2.n98 VSUBS 2.02745f
C617 VDD2.t4 VSUBS 0.199923f
C618 VDD2.t0 VSUBS 0.199923f
C619 VDD2.n99 VSUBS 1.45137f
C620 VDD2.n100 VSUBS 0.596516f
C621 VDD2.t9 VSUBS 0.199923f
C622 VDD2.t7 VSUBS 0.199923f
C623 VDD2.n101 VSUBS 1.45432f
C624 VN.n0 VSUBS 0.066787f
C625 VN.t4 VSUBS 0.572948f
C626 VN.n1 VSUBS 0.25699f
C627 VN.t8 VSUBS 0.584332f
C628 VN.n2 VSUBS 0.24651f
C629 VN.n3 VSUBS 0.221281f
C630 VN.t3 VSUBS 0.572948f
C631 VN.n4 VSUBS 0.26399f
C632 VN.t7 VSUBS 0.572948f
C633 VN.n5 VSUBS 0.25699f
C634 VN.t6 VSUBS 0.58082f
C635 VN.n6 VSUBS 0.24953f
C636 VN.n7 VSUBS 0.051757f
C637 VN.n8 VSUBS 0.066787f
C638 VN.t1 VSUBS 0.58082f
C639 VN.t0 VSUBS 0.572948f
C640 VN.n9 VSUBS 0.25699f
C641 VN.t9 VSUBS 0.572948f
C642 VN.t2 VSUBS 0.584332f
C643 VN.n10 VSUBS 0.24651f
C644 VN.n11 VSUBS 0.221281f
C645 VN.n12 VSUBS 0.26399f
C646 VN.t5 VSUBS 0.572948f
C647 VN.n13 VSUBS 0.25699f
C648 VN.n14 VSUBS 0.24953f
C649 VN.n15 VSUBS 2.41991f
C650 VTAIL.t5 VSUBS 0.224577f
C651 VTAIL.t19 VSUBS 0.224577f
C652 VTAIL.n0 VSUBS 1.47431f
C653 VTAIL.n1 VSUBS 0.831118f
C654 VTAIL.n2 VSUBS 0.036349f
C655 VTAIL.n3 VSUBS 0.032331f
C656 VTAIL.n4 VSUBS 0.017373f
C657 VTAIL.n5 VSUBS 0.041064f
C658 VTAIL.n6 VSUBS 0.018395f
C659 VTAIL.n7 VSUBS 0.032331f
C660 VTAIL.n8 VSUBS 0.017373f
C661 VTAIL.n9 VSUBS 0.041064f
C662 VTAIL.n10 VSUBS 0.018395f
C663 VTAIL.n11 VSUBS 0.032331f
C664 VTAIL.n12 VSUBS 0.017373f
C665 VTAIL.n13 VSUBS 0.041064f
C666 VTAIL.n14 VSUBS 0.018395f
C667 VTAIL.n15 VSUBS 1.15269f
C668 VTAIL.n16 VSUBS 0.017373f
C669 VTAIL.t13 VSUBS 0.08754f
C670 VTAIL.n17 VSUBS 0.168815f
C671 VTAIL.n18 VSUBS 0.026123f
C672 VTAIL.n19 VSUBS 0.030798f
C673 VTAIL.n20 VSUBS 0.041064f
C674 VTAIL.n21 VSUBS 0.018395f
C675 VTAIL.n22 VSUBS 0.017373f
C676 VTAIL.n23 VSUBS 0.032331f
C677 VTAIL.n24 VSUBS 0.032331f
C678 VTAIL.n25 VSUBS 0.017373f
C679 VTAIL.n26 VSUBS 0.018395f
C680 VTAIL.n27 VSUBS 0.041064f
C681 VTAIL.n28 VSUBS 0.041064f
C682 VTAIL.n29 VSUBS 0.018395f
C683 VTAIL.n30 VSUBS 0.017373f
C684 VTAIL.n31 VSUBS 0.032331f
C685 VTAIL.n32 VSUBS 0.032331f
C686 VTAIL.n33 VSUBS 0.017373f
C687 VTAIL.n34 VSUBS 0.018395f
C688 VTAIL.n35 VSUBS 0.041064f
C689 VTAIL.n36 VSUBS 0.041064f
C690 VTAIL.n37 VSUBS 0.018395f
C691 VTAIL.n38 VSUBS 0.017373f
C692 VTAIL.n39 VSUBS 0.032331f
C693 VTAIL.n40 VSUBS 0.032331f
C694 VTAIL.n41 VSUBS 0.017373f
C695 VTAIL.n42 VSUBS 0.018395f
C696 VTAIL.n43 VSUBS 0.041064f
C697 VTAIL.n44 VSUBS 0.10222f
C698 VTAIL.n45 VSUBS 0.018395f
C699 VTAIL.n46 VSUBS 0.017373f
C700 VTAIL.n47 VSUBS 0.070757f
C701 VTAIL.n48 VSUBS 0.051405f
C702 VTAIL.n49 VSUBS 0.164577f
C703 VTAIL.t10 VSUBS 0.224577f
C704 VTAIL.t15 VSUBS 0.224577f
C705 VTAIL.n50 VSUBS 1.47431f
C706 VTAIL.n51 VSUBS 0.821239f
C707 VTAIL.t12 VSUBS 0.224577f
C708 VTAIL.t11 VSUBS 0.224577f
C709 VTAIL.n52 VSUBS 1.47431f
C710 VTAIL.n53 VSUBS 2.11002f
C711 VTAIL.t17 VSUBS 0.224577f
C712 VTAIL.t3 VSUBS 0.224577f
C713 VTAIL.n54 VSUBS 1.47432f
C714 VTAIL.n55 VSUBS 2.11f
C715 VTAIL.t4 VSUBS 0.224577f
C716 VTAIL.t16 VSUBS 0.224577f
C717 VTAIL.n56 VSUBS 1.47432f
C718 VTAIL.n57 VSUBS 0.821228f
C719 VTAIL.n58 VSUBS 0.036349f
C720 VTAIL.n59 VSUBS 0.032331f
C721 VTAIL.n60 VSUBS 0.017373f
C722 VTAIL.n61 VSUBS 0.041064f
C723 VTAIL.n62 VSUBS 0.018395f
C724 VTAIL.n63 VSUBS 0.032331f
C725 VTAIL.n64 VSUBS 0.017373f
C726 VTAIL.n65 VSUBS 0.041064f
C727 VTAIL.n66 VSUBS 0.018395f
C728 VTAIL.n67 VSUBS 0.032331f
C729 VTAIL.n68 VSUBS 0.017373f
C730 VTAIL.n69 VSUBS 0.041064f
C731 VTAIL.n70 VSUBS 0.018395f
C732 VTAIL.n71 VSUBS 1.15269f
C733 VTAIL.n72 VSUBS 0.017373f
C734 VTAIL.t18 VSUBS 0.08754f
C735 VTAIL.n73 VSUBS 0.168815f
C736 VTAIL.n74 VSUBS 0.026123f
C737 VTAIL.n75 VSUBS 0.030798f
C738 VTAIL.n76 VSUBS 0.041064f
C739 VTAIL.n77 VSUBS 0.018395f
C740 VTAIL.n78 VSUBS 0.017373f
C741 VTAIL.n79 VSUBS 0.032331f
C742 VTAIL.n80 VSUBS 0.032331f
C743 VTAIL.n81 VSUBS 0.017373f
C744 VTAIL.n82 VSUBS 0.018395f
C745 VTAIL.n83 VSUBS 0.041064f
C746 VTAIL.n84 VSUBS 0.041064f
C747 VTAIL.n85 VSUBS 0.018395f
C748 VTAIL.n86 VSUBS 0.017373f
C749 VTAIL.n87 VSUBS 0.032331f
C750 VTAIL.n88 VSUBS 0.032331f
C751 VTAIL.n89 VSUBS 0.017373f
C752 VTAIL.n90 VSUBS 0.018395f
C753 VTAIL.n91 VSUBS 0.041064f
C754 VTAIL.n92 VSUBS 0.041064f
C755 VTAIL.n93 VSUBS 0.018395f
C756 VTAIL.n94 VSUBS 0.017373f
C757 VTAIL.n95 VSUBS 0.032331f
C758 VTAIL.n96 VSUBS 0.032331f
C759 VTAIL.n97 VSUBS 0.017373f
C760 VTAIL.n98 VSUBS 0.018395f
C761 VTAIL.n99 VSUBS 0.041064f
C762 VTAIL.n100 VSUBS 0.10222f
C763 VTAIL.n101 VSUBS 0.018395f
C764 VTAIL.n102 VSUBS 0.017373f
C765 VTAIL.n103 VSUBS 0.070757f
C766 VTAIL.n104 VSUBS 0.051405f
C767 VTAIL.n105 VSUBS 0.164577f
C768 VTAIL.t8 VSUBS 0.224577f
C769 VTAIL.t14 VSUBS 0.224577f
C770 VTAIL.n106 VSUBS 1.47432f
C771 VTAIL.n107 VSUBS 0.840088f
C772 VTAIL.t6 VSUBS 0.224577f
C773 VTAIL.t7 VSUBS 0.224577f
C774 VTAIL.n108 VSUBS 1.47432f
C775 VTAIL.n109 VSUBS 0.821228f
C776 VTAIL.n110 VSUBS 0.036349f
C777 VTAIL.n111 VSUBS 0.032331f
C778 VTAIL.n112 VSUBS 0.017373f
C779 VTAIL.n113 VSUBS 0.041064f
C780 VTAIL.n114 VSUBS 0.018395f
C781 VTAIL.n115 VSUBS 0.032331f
C782 VTAIL.n116 VSUBS 0.017373f
C783 VTAIL.n117 VSUBS 0.041064f
C784 VTAIL.n118 VSUBS 0.018395f
C785 VTAIL.n119 VSUBS 0.032331f
C786 VTAIL.n120 VSUBS 0.017373f
C787 VTAIL.n121 VSUBS 0.041064f
C788 VTAIL.n122 VSUBS 0.018395f
C789 VTAIL.n123 VSUBS 1.15269f
C790 VTAIL.n124 VSUBS 0.017373f
C791 VTAIL.t9 VSUBS 0.08754f
C792 VTAIL.n125 VSUBS 0.168814f
C793 VTAIL.n126 VSUBS 0.026123f
C794 VTAIL.n127 VSUBS 0.030798f
C795 VTAIL.n128 VSUBS 0.041064f
C796 VTAIL.n129 VSUBS 0.018395f
C797 VTAIL.n130 VSUBS 0.017373f
C798 VTAIL.n131 VSUBS 0.032331f
C799 VTAIL.n132 VSUBS 0.032331f
C800 VTAIL.n133 VSUBS 0.017373f
C801 VTAIL.n134 VSUBS 0.018395f
C802 VTAIL.n135 VSUBS 0.041064f
C803 VTAIL.n136 VSUBS 0.041064f
C804 VTAIL.n137 VSUBS 0.018395f
C805 VTAIL.n138 VSUBS 0.017373f
C806 VTAIL.n139 VSUBS 0.032331f
C807 VTAIL.n140 VSUBS 0.032331f
C808 VTAIL.n141 VSUBS 0.017373f
C809 VTAIL.n142 VSUBS 0.018395f
C810 VTAIL.n143 VSUBS 0.041064f
C811 VTAIL.n144 VSUBS 0.041064f
C812 VTAIL.n145 VSUBS 0.018395f
C813 VTAIL.n146 VSUBS 0.017373f
C814 VTAIL.n147 VSUBS 0.032331f
C815 VTAIL.n148 VSUBS 0.032331f
C816 VTAIL.n149 VSUBS 0.017373f
C817 VTAIL.n150 VSUBS 0.018395f
C818 VTAIL.n151 VSUBS 0.041064f
C819 VTAIL.n152 VSUBS 0.10222f
C820 VTAIL.n153 VSUBS 0.018395f
C821 VTAIL.n154 VSUBS 0.017373f
C822 VTAIL.n155 VSUBS 0.070757f
C823 VTAIL.n156 VSUBS 0.051405f
C824 VTAIL.n157 VSUBS 1.37432f
C825 VTAIL.n158 VSUBS 0.036349f
C826 VTAIL.n159 VSUBS 0.032331f
C827 VTAIL.n160 VSUBS 0.017373f
C828 VTAIL.n161 VSUBS 0.041064f
C829 VTAIL.n162 VSUBS 0.018395f
C830 VTAIL.n163 VSUBS 0.032331f
C831 VTAIL.n164 VSUBS 0.017373f
C832 VTAIL.n165 VSUBS 0.041064f
C833 VTAIL.n166 VSUBS 0.018395f
C834 VTAIL.n167 VSUBS 0.032331f
C835 VTAIL.n168 VSUBS 0.017373f
C836 VTAIL.n169 VSUBS 0.041064f
C837 VTAIL.n170 VSUBS 0.018395f
C838 VTAIL.n171 VSUBS 1.15269f
C839 VTAIL.n172 VSUBS 0.017373f
C840 VTAIL.t1 VSUBS 0.08754f
C841 VTAIL.n173 VSUBS 0.168815f
C842 VTAIL.n174 VSUBS 0.026123f
C843 VTAIL.n175 VSUBS 0.030798f
C844 VTAIL.n176 VSUBS 0.041064f
C845 VTAIL.n177 VSUBS 0.018395f
C846 VTAIL.n178 VSUBS 0.017373f
C847 VTAIL.n179 VSUBS 0.032331f
C848 VTAIL.n180 VSUBS 0.032331f
C849 VTAIL.n181 VSUBS 0.017373f
C850 VTAIL.n182 VSUBS 0.018395f
C851 VTAIL.n183 VSUBS 0.041064f
C852 VTAIL.n184 VSUBS 0.041064f
C853 VTAIL.n185 VSUBS 0.018395f
C854 VTAIL.n186 VSUBS 0.017373f
C855 VTAIL.n187 VSUBS 0.032331f
C856 VTAIL.n188 VSUBS 0.032331f
C857 VTAIL.n189 VSUBS 0.017373f
C858 VTAIL.n190 VSUBS 0.018395f
C859 VTAIL.n191 VSUBS 0.041064f
C860 VTAIL.n192 VSUBS 0.041064f
C861 VTAIL.n193 VSUBS 0.018395f
C862 VTAIL.n194 VSUBS 0.017373f
C863 VTAIL.n195 VSUBS 0.032331f
C864 VTAIL.n196 VSUBS 0.032331f
C865 VTAIL.n197 VSUBS 0.017373f
C866 VTAIL.n198 VSUBS 0.018395f
C867 VTAIL.n199 VSUBS 0.041064f
C868 VTAIL.n200 VSUBS 0.10222f
C869 VTAIL.n201 VSUBS 0.018395f
C870 VTAIL.n202 VSUBS 0.017373f
C871 VTAIL.n203 VSUBS 0.070757f
C872 VTAIL.n204 VSUBS 0.051405f
C873 VTAIL.n205 VSUBS 1.37432f
C874 VTAIL.t0 VSUBS 0.224577f
C875 VTAIL.t2 VSUBS 0.224577f
C876 VTAIL.n206 VSUBS 1.47431f
C877 VTAIL.n207 VSUBS 0.770048f
C878 VDD1.n0 VSUBS 0.032173f
C879 VDD1.n1 VSUBS 0.028617f
C880 VDD1.n2 VSUBS 0.015377f
C881 VDD1.n3 VSUBS 0.036346f
C882 VDD1.n4 VSUBS 0.016282f
C883 VDD1.n5 VSUBS 0.028617f
C884 VDD1.n6 VSUBS 0.015377f
C885 VDD1.n7 VSUBS 0.036346f
C886 VDD1.n8 VSUBS 0.016282f
C887 VDD1.n9 VSUBS 0.028617f
C888 VDD1.n10 VSUBS 0.015377f
C889 VDD1.n11 VSUBS 0.036346f
C890 VDD1.n12 VSUBS 0.016282f
C891 VDD1.n13 VSUBS 1.02025f
C892 VDD1.n14 VSUBS 0.015377f
C893 VDD1.t6 VSUBS 0.077482f
C894 VDD1.n15 VSUBS 0.149419f
C895 VDD1.n16 VSUBS 0.023122f
C896 VDD1.n17 VSUBS 0.02726f
C897 VDD1.n18 VSUBS 0.036346f
C898 VDD1.n19 VSUBS 0.016282f
C899 VDD1.n20 VSUBS 0.015377f
C900 VDD1.n21 VSUBS 0.028617f
C901 VDD1.n22 VSUBS 0.028617f
C902 VDD1.n23 VSUBS 0.015377f
C903 VDD1.n24 VSUBS 0.016282f
C904 VDD1.n25 VSUBS 0.036346f
C905 VDD1.n26 VSUBS 0.036346f
C906 VDD1.n27 VSUBS 0.016282f
C907 VDD1.n28 VSUBS 0.015377f
C908 VDD1.n29 VSUBS 0.028617f
C909 VDD1.n30 VSUBS 0.028617f
C910 VDD1.n31 VSUBS 0.015377f
C911 VDD1.n32 VSUBS 0.016282f
C912 VDD1.n33 VSUBS 0.036346f
C913 VDD1.n34 VSUBS 0.036346f
C914 VDD1.n35 VSUBS 0.016282f
C915 VDD1.n36 VSUBS 0.015377f
C916 VDD1.n37 VSUBS 0.028617f
C917 VDD1.n38 VSUBS 0.028617f
C918 VDD1.n39 VSUBS 0.015377f
C919 VDD1.n40 VSUBS 0.016282f
C920 VDD1.n41 VSUBS 0.036346f
C921 VDD1.n42 VSUBS 0.090476f
C922 VDD1.n43 VSUBS 0.016282f
C923 VDD1.n44 VSUBS 0.015377f
C924 VDD1.n45 VSUBS 0.062628f
C925 VDD1.n46 VSUBS 0.066576f
C926 VDD1.t0 VSUBS 0.198775f
C927 VDD1.t2 VSUBS 0.198775f
C928 VDD1.n47 VSUBS 1.44304f
C929 VDD1.n48 VSUBS 0.698151f
C930 VDD1.n49 VSUBS 0.032173f
C931 VDD1.n50 VSUBS 0.028617f
C932 VDD1.n51 VSUBS 0.015377f
C933 VDD1.n52 VSUBS 0.036346f
C934 VDD1.n53 VSUBS 0.016282f
C935 VDD1.n54 VSUBS 0.028617f
C936 VDD1.n55 VSUBS 0.015377f
C937 VDD1.n56 VSUBS 0.036346f
C938 VDD1.n57 VSUBS 0.016282f
C939 VDD1.n58 VSUBS 0.028617f
C940 VDD1.n59 VSUBS 0.015377f
C941 VDD1.n60 VSUBS 0.036346f
C942 VDD1.n61 VSUBS 0.016282f
C943 VDD1.n62 VSUBS 1.02025f
C944 VDD1.n63 VSUBS 0.015377f
C945 VDD1.t7 VSUBS 0.077482f
C946 VDD1.n64 VSUBS 0.149419f
C947 VDD1.n65 VSUBS 0.023122f
C948 VDD1.n66 VSUBS 0.02726f
C949 VDD1.n67 VSUBS 0.036346f
C950 VDD1.n68 VSUBS 0.016282f
C951 VDD1.n69 VSUBS 0.015377f
C952 VDD1.n70 VSUBS 0.028617f
C953 VDD1.n71 VSUBS 0.028617f
C954 VDD1.n72 VSUBS 0.015377f
C955 VDD1.n73 VSUBS 0.016282f
C956 VDD1.n74 VSUBS 0.036346f
C957 VDD1.n75 VSUBS 0.036346f
C958 VDD1.n76 VSUBS 0.016282f
C959 VDD1.n77 VSUBS 0.015377f
C960 VDD1.n78 VSUBS 0.028617f
C961 VDD1.n79 VSUBS 0.028617f
C962 VDD1.n80 VSUBS 0.015377f
C963 VDD1.n81 VSUBS 0.016282f
C964 VDD1.n82 VSUBS 0.036346f
C965 VDD1.n83 VSUBS 0.036346f
C966 VDD1.n84 VSUBS 0.016282f
C967 VDD1.n85 VSUBS 0.015377f
C968 VDD1.n86 VSUBS 0.028617f
C969 VDD1.n87 VSUBS 0.028617f
C970 VDD1.n88 VSUBS 0.015377f
C971 VDD1.n89 VSUBS 0.016282f
C972 VDD1.n90 VSUBS 0.036346f
C973 VDD1.n91 VSUBS 0.090476f
C974 VDD1.n92 VSUBS 0.016282f
C975 VDD1.n93 VSUBS 0.015377f
C976 VDD1.n94 VSUBS 0.062628f
C977 VDD1.n95 VSUBS 0.066576f
C978 VDD1.t8 VSUBS 0.198775f
C979 VDD1.t4 VSUBS 0.198775f
C980 VDD1.n96 VSUBS 1.44303f
C981 VDD1.n97 VSUBS 0.69514f
C982 VDD1.t5 VSUBS 0.198775f
C983 VDD1.t3 VSUBS 0.198775f
C984 VDD1.n98 VSUBS 1.44599f
C985 VDD1.n99 VSUBS 2.09824f
C986 VDD1.t1 VSUBS 0.198775f
C987 VDD1.t9 VSUBS 0.198775f
C988 VDD1.n100 VSUBS 1.44304f
C989 VDD1.n101 VSUBS 2.55787f
C990 VP.n0 VSUBS 0.069681f
C991 VP.t4 VSUBS 0.597774f
C992 VP.n1 VSUBS 0.268125f
C993 VP.n2 VSUBS 0.069681f
C994 VP.t8 VSUBS 0.597774f
C995 VP.t9 VSUBS 0.597774f
C996 VP.n3 VSUBS 0.230869f
C997 VP.t1 VSUBS 0.597774f
C998 VP.t7 VSUBS 0.609651f
C999 VP.n4 VSUBS 0.257192f
C1000 VP.n5 VSUBS 0.268125f
C1001 VP.n6 VSUBS 0.275429f
C1002 VP.n7 VSUBS 0.268125f
C1003 VP.t6 VSUBS 0.605987f
C1004 VP.n8 VSUBS 0.260342f
C1005 VP.n9 VSUBS 2.47876f
C1006 VP.t3 VSUBS 0.605987f
C1007 VP.n10 VSUBS 0.260342f
C1008 VP.n11 VSUBS 2.54379f
C1009 VP.n12 VSUBS 0.069681f
C1010 VP.n13 VSUBS 0.069681f
C1011 VP.t5 VSUBS 0.597774f
C1012 VP.n14 VSUBS 0.275429f
C1013 VP.t0 VSUBS 0.597774f
C1014 VP.n15 VSUBS 0.268125f
C1015 VP.t2 VSUBS 0.605987f
C1016 VP.n16 VSUBS 0.260342f
C1017 VP.n17 VSUBS 0.054f
.ends

