* NGSPICE file created from diff_pair_sample_0482.ext - technology: sky130A

.subckt diff_pair_sample_0482 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0.89595 ps=5.76 w=5.43 l=1.4
X1 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0.89595 ps=5.76 w=5.43 l=1.4
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0 ps=0 w=5.43 l=1.4
X3 VTAIL.t4 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=0.89595 ps=5.76 w=5.43 l=1.4
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0 ps=0 w=5.43 l=1.4
X5 VTAIL.t10 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=0.89595 ps=5.76 w=5.43 l=1.4
X6 VDD2.t3 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=2.1177 ps=11.64 w=5.43 l=1.4
X7 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0.89595 ps=5.76 w=5.43 l=1.4
X8 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0 ps=0 w=5.43 l=1.4
X9 VDD1.t3 VP.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=2.1177 ps=11.64 w=5.43 l=1.4
X10 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=2.1177 ps=11.64 w=5.43 l=1.4
X11 VTAIL.t7 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=0.89595 ps=5.76 w=5.43 l=1.4
X12 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=0.89595 ps=5.76 w=5.43 l=1.4
X13 VDD1.t1 VP.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.89595 pd=5.76 as=2.1177 ps=11.64 w=5.43 l=1.4
X14 VDD1.t0 VP.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0.89595 ps=5.76 w=5.43 l=1.4
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1177 pd=11.64 as=0 ps=0 w=5.43 l=1.4
R0 VP.n15 VP.n14 174.512
R1 VP.n27 VP.n26 174.512
R2 VP.n13 VP.n12 174.512
R3 VP.n8 VP.n5 161.3
R4 VP.n10 VP.n9 161.3
R5 VP.n11 VP.n4 161.3
R6 VP.n25 VP.n0 161.3
R7 VP.n24 VP.n23 161.3
R8 VP.n22 VP.n1 161.3
R9 VP.n21 VP.n20 161.3
R10 VP.n19 VP.n2 161.3
R11 VP.n18 VP.n17 161.3
R12 VP.n16 VP.n3 161.3
R13 VP.n7 VP.t0 128.267
R14 VP.n20 VP.t3 93.4741
R15 VP.n14 VP.t5 93.4741
R16 VP.n26 VP.t4 93.4741
R17 VP.n6 VP.t1 93.4741
R18 VP.n12 VP.t2 93.4741
R19 VP.n19 VP.n18 53.6055
R20 VP.n24 VP.n1 53.6055
R21 VP.n10 VP.n5 53.6055
R22 VP.n7 VP.n6 41.8065
R23 VP.n15 VP.n13 38.9134
R24 VP.n18 VP.n3 27.3813
R25 VP.n25 VP.n24 27.3813
R26 VP.n11 VP.n10 27.3813
R27 VP.n20 VP.n19 24.4675
R28 VP.n20 VP.n1 24.4675
R29 VP.n6 VP.n5 24.4675
R30 VP.n8 VP.n7 17.6362
R31 VP.n14 VP.n3 11.2553
R32 VP.n26 VP.n25 11.2553
R33 VP.n12 VP.n11 11.2553
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n4 0.189894
R36 VP.n13 VP.n4 0.189894
R37 VP.n16 VP.n15 0.189894
R38 VP.n17 VP.n16 0.189894
R39 VP.n17 VP.n2 0.189894
R40 VP.n21 VP.n2 0.189894
R41 VP.n22 VP.n21 0.189894
R42 VP.n23 VP.n22 0.189894
R43 VP.n23 VP.n0 0.189894
R44 VP.n27 VP.n0 0.189894
R45 VP VP.n27 0.0516364
R46 VTAIL.n114 VTAIL.n92 289.615
R47 VTAIL.n24 VTAIL.n2 289.615
R48 VTAIL.n86 VTAIL.n64 289.615
R49 VTAIL.n56 VTAIL.n34 289.615
R50 VTAIL.n100 VTAIL.n99 185
R51 VTAIL.n105 VTAIL.n104 185
R52 VTAIL.n107 VTAIL.n106 185
R53 VTAIL.n96 VTAIL.n95 185
R54 VTAIL.n113 VTAIL.n112 185
R55 VTAIL.n115 VTAIL.n114 185
R56 VTAIL.n10 VTAIL.n9 185
R57 VTAIL.n15 VTAIL.n14 185
R58 VTAIL.n17 VTAIL.n16 185
R59 VTAIL.n6 VTAIL.n5 185
R60 VTAIL.n23 VTAIL.n22 185
R61 VTAIL.n25 VTAIL.n24 185
R62 VTAIL.n87 VTAIL.n86 185
R63 VTAIL.n85 VTAIL.n84 185
R64 VTAIL.n68 VTAIL.n67 185
R65 VTAIL.n79 VTAIL.n78 185
R66 VTAIL.n77 VTAIL.n76 185
R67 VTAIL.n72 VTAIL.n71 185
R68 VTAIL.n57 VTAIL.n56 185
R69 VTAIL.n55 VTAIL.n54 185
R70 VTAIL.n38 VTAIL.n37 185
R71 VTAIL.n49 VTAIL.n48 185
R72 VTAIL.n47 VTAIL.n46 185
R73 VTAIL.n42 VTAIL.n41 185
R74 VTAIL.n101 VTAIL.t5 147.672
R75 VTAIL.n11 VTAIL.t11 147.672
R76 VTAIL.n73 VTAIL.t9 147.672
R77 VTAIL.n43 VTAIL.t0 147.672
R78 VTAIL.n105 VTAIL.n99 104.615
R79 VTAIL.n106 VTAIL.n105 104.615
R80 VTAIL.n106 VTAIL.n95 104.615
R81 VTAIL.n113 VTAIL.n95 104.615
R82 VTAIL.n114 VTAIL.n113 104.615
R83 VTAIL.n15 VTAIL.n9 104.615
R84 VTAIL.n16 VTAIL.n15 104.615
R85 VTAIL.n16 VTAIL.n5 104.615
R86 VTAIL.n23 VTAIL.n5 104.615
R87 VTAIL.n24 VTAIL.n23 104.615
R88 VTAIL.n86 VTAIL.n85 104.615
R89 VTAIL.n85 VTAIL.n67 104.615
R90 VTAIL.n78 VTAIL.n67 104.615
R91 VTAIL.n78 VTAIL.n77 104.615
R92 VTAIL.n77 VTAIL.n71 104.615
R93 VTAIL.n56 VTAIL.n55 104.615
R94 VTAIL.n55 VTAIL.n37 104.615
R95 VTAIL.n48 VTAIL.n37 104.615
R96 VTAIL.n48 VTAIL.n47 104.615
R97 VTAIL.n47 VTAIL.n41 104.615
R98 VTAIL.n63 VTAIL.n62 54.8856
R99 VTAIL.n33 VTAIL.n32 54.8856
R100 VTAIL.n1 VTAIL.n0 54.8854
R101 VTAIL.n31 VTAIL.n30 54.8854
R102 VTAIL.t5 VTAIL.n99 52.3082
R103 VTAIL.t11 VTAIL.n9 52.3082
R104 VTAIL.t9 VTAIL.n71 52.3082
R105 VTAIL.t0 VTAIL.n41 52.3082
R106 VTAIL.n119 VTAIL.n118 35.0944
R107 VTAIL.n29 VTAIL.n28 35.0944
R108 VTAIL.n91 VTAIL.n90 35.0944
R109 VTAIL.n61 VTAIL.n60 35.0944
R110 VTAIL.n33 VTAIL.n31 20.0307
R111 VTAIL.n119 VTAIL.n91 18.5393
R112 VTAIL.n101 VTAIL.n100 15.6666
R113 VTAIL.n11 VTAIL.n10 15.6666
R114 VTAIL.n73 VTAIL.n72 15.6666
R115 VTAIL.n43 VTAIL.n42 15.6666
R116 VTAIL.n104 VTAIL.n103 12.8005
R117 VTAIL.n14 VTAIL.n13 12.8005
R118 VTAIL.n76 VTAIL.n75 12.8005
R119 VTAIL.n46 VTAIL.n45 12.8005
R120 VTAIL.n107 VTAIL.n98 12.0247
R121 VTAIL.n17 VTAIL.n8 12.0247
R122 VTAIL.n79 VTAIL.n70 12.0247
R123 VTAIL.n49 VTAIL.n40 12.0247
R124 VTAIL.n108 VTAIL.n96 11.249
R125 VTAIL.n18 VTAIL.n6 11.249
R126 VTAIL.n80 VTAIL.n68 11.249
R127 VTAIL.n50 VTAIL.n38 11.249
R128 VTAIL.n112 VTAIL.n111 10.4732
R129 VTAIL.n22 VTAIL.n21 10.4732
R130 VTAIL.n84 VTAIL.n83 10.4732
R131 VTAIL.n54 VTAIL.n53 10.4732
R132 VTAIL.n115 VTAIL.n94 9.69747
R133 VTAIL.n25 VTAIL.n4 9.69747
R134 VTAIL.n87 VTAIL.n66 9.69747
R135 VTAIL.n57 VTAIL.n36 9.69747
R136 VTAIL.n118 VTAIL.n117 9.45567
R137 VTAIL.n28 VTAIL.n27 9.45567
R138 VTAIL.n90 VTAIL.n89 9.45567
R139 VTAIL.n60 VTAIL.n59 9.45567
R140 VTAIL.n117 VTAIL.n116 9.3005
R141 VTAIL.n94 VTAIL.n93 9.3005
R142 VTAIL.n111 VTAIL.n110 9.3005
R143 VTAIL.n109 VTAIL.n108 9.3005
R144 VTAIL.n98 VTAIL.n97 9.3005
R145 VTAIL.n103 VTAIL.n102 9.3005
R146 VTAIL.n27 VTAIL.n26 9.3005
R147 VTAIL.n4 VTAIL.n3 9.3005
R148 VTAIL.n21 VTAIL.n20 9.3005
R149 VTAIL.n19 VTAIL.n18 9.3005
R150 VTAIL.n8 VTAIL.n7 9.3005
R151 VTAIL.n13 VTAIL.n12 9.3005
R152 VTAIL.n89 VTAIL.n88 9.3005
R153 VTAIL.n66 VTAIL.n65 9.3005
R154 VTAIL.n83 VTAIL.n82 9.3005
R155 VTAIL.n81 VTAIL.n80 9.3005
R156 VTAIL.n70 VTAIL.n69 9.3005
R157 VTAIL.n75 VTAIL.n74 9.3005
R158 VTAIL.n59 VTAIL.n58 9.3005
R159 VTAIL.n36 VTAIL.n35 9.3005
R160 VTAIL.n53 VTAIL.n52 9.3005
R161 VTAIL.n51 VTAIL.n50 9.3005
R162 VTAIL.n40 VTAIL.n39 9.3005
R163 VTAIL.n45 VTAIL.n44 9.3005
R164 VTAIL.n116 VTAIL.n92 8.92171
R165 VTAIL.n26 VTAIL.n2 8.92171
R166 VTAIL.n88 VTAIL.n64 8.92171
R167 VTAIL.n58 VTAIL.n34 8.92171
R168 VTAIL.n118 VTAIL.n92 5.04292
R169 VTAIL.n28 VTAIL.n2 5.04292
R170 VTAIL.n90 VTAIL.n64 5.04292
R171 VTAIL.n60 VTAIL.n34 5.04292
R172 VTAIL.n102 VTAIL.n101 4.38687
R173 VTAIL.n12 VTAIL.n11 4.38687
R174 VTAIL.n74 VTAIL.n73 4.38687
R175 VTAIL.n44 VTAIL.n43 4.38687
R176 VTAIL.n116 VTAIL.n115 4.26717
R177 VTAIL.n26 VTAIL.n25 4.26717
R178 VTAIL.n88 VTAIL.n87 4.26717
R179 VTAIL.n58 VTAIL.n57 4.26717
R180 VTAIL.n0 VTAIL.t1 3.64691
R181 VTAIL.n0 VTAIL.t4 3.64691
R182 VTAIL.n30 VTAIL.t6 3.64691
R183 VTAIL.n30 VTAIL.t7 3.64691
R184 VTAIL.n62 VTAIL.t8 3.64691
R185 VTAIL.n62 VTAIL.t10 3.64691
R186 VTAIL.n32 VTAIL.t2 3.64691
R187 VTAIL.n32 VTAIL.t3 3.64691
R188 VTAIL.n112 VTAIL.n94 3.49141
R189 VTAIL.n22 VTAIL.n4 3.49141
R190 VTAIL.n84 VTAIL.n66 3.49141
R191 VTAIL.n54 VTAIL.n36 3.49141
R192 VTAIL.n111 VTAIL.n96 2.71565
R193 VTAIL.n21 VTAIL.n6 2.71565
R194 VTAIL.n83 VTAIL.n68 2.71565
R195 VTAIL.n53 VTAIL.n38 2.71565
R196 VTAIL.n108 VTAIL.n107 1.93989
R197 VTAIL.n18 VTAIL.n17 1.93989
R198 VTAIL.n80 VTAIL.n79 1.93989
R199 VTAIL.n50 VTAIL.n49 1.93989
R200 VTAIL.n61 VTAIL.n33 1.49188
R201 VTAIL.n91 VTAIL.n63 1.49188
R202 VTAIL.n31 VTAIL.n29 1.49188
R203 VTAIL.n63 VTAIL.n61 1.21602
R204 VTAIL.n29 VTAIL.n1 1.21602
R205 VTAIL.n104 VTAIL.n98 1.16414
R206 VTAIL.n14 VTAIL.n8 1.16414
R207 VTAIL.n76 VTAIL.n70 1.16414
R208 VTAIL.n46 VTAIL.n40 1.16414
R209 VTAIL VTAIL.n119 1.06084
R210 VTAIL VTAIL.n1 0.431534
R211 VTAIL.n103 VTAIL.n100 0.388379
R212 VTAIL.n13 VTAIL.n10 0.388379
R213 VTAIL.n75 VTAIL.n72 0.388379
R214 VTAIL.n45 VTAIL.n42 0.388379
R215 VTAIL.n102 VTAIL.n97 0.155672
R216 VTAIL.n109 VTAIL.n97 0.155672
R217 VTAIL.n110 VTAIL.n109 0.155672
R218 VTAIL.n110 VTAIL.n93 0.155672
R219 VTAIL.n117 VTAIL.n93 0.155672
R220 VTAIL.n12 VTAIL.n7 0.155672
R221 VTAIL.n19 VTAIL.n7 0.155672
R222 VTAIL.n20 VTAIL.n19 0.155672
R223 VTAIL.n20 VTAIL.n3 0.155672
R224 VTAIL.n27 VTAIL.n3 0.155672
R225 VTAIL.n89 VTAIL.n65 0.155672
R226 VTAIL.n82 VTAIL.n65 0.155672
R227 VTAIL.n82 VTAIL.n81 0.155672
R228 VTAIL.n81 VTAIL.n69 0.155672
R229 VTAIL.n74 VTAIL.n69 0.155672
R230 VTAIL.n59 VTAIL.n35 0.155672
R231 VTAIL.n52 VTAIL.n35 0.155672
R232 VTAIL.n52 VTAIL.n51 0.155672
R233 VTAIL.n51 VTAIL.n39 0.155672
R234 VTAIL.n44 VTAIL.n39 0.155672
R235 VDD1.n22 VDD1.n0 289.615
R236 VDD1.n49 VDD1.n27 289.615
R237 VDD1.n23 VDD1.n22 185
R238 VDD1.n21 VDD1.n20 185
R239 VDD1.n4 VDD1.n3 185
R240 VDD1.n15 VDD1.n14 185
R241 VDD1.n13 VDD1.n12 185
R242 VDD1.n8 VDD1.n7 185
R243 VDD1.n35 VDD1.n34 185
R244 VDD1.n40 VDD1.n39 185
R245 VDD1.n42 VDD1.n41 185
R246 VDD1.n31 VDD1.n30 185
R247 VDD1.n48 VDD1.n47 185
R248 VDD1.n50 VDD1.n49 185
R249 VDD1.n9 VDD1.t5 147.672
R250 VDD1.n36 VDD1.t0 147.672
R251 VDD1.n22 VDD1.n21 104.615
R252 VDD1.n21 VDD1.n3 104.615
R253 VDD1.n14 VDD1.n3 104.615
R254 VDD1.n14 VDD1.n13 104.615
R255 VDD1.n13 VDD1.n7 104.615
R256 VDD1.n40 VDD1.n34 104.615
R257 VDD1.n41 VDD1.n40 104.615
R258 VDD1.n41 VDD1.n30 104.615
R259 VDD1.n48 VDD1.n30 104.615
R260 VDD1.n49 VDD1.n48 104.615
R261 VDD1.n55 VDD1.n54 71.8817
R262 VDD1.n57 VDD1.n56 71.5642
R263 VDD1 VDD1.n26 52.95
R264 VDD1.n55 VDD1.n53 52.8364
R265 VDD1.t5 VDD1.n7 52.3082
R266 VDD1.t0 VDD1.n34 52.3082
R267 VDD1.n57 VDD1.n55 34.572
R268 VDD1.n9 VDD1.n8 15.6666
R269 VDD1.n36 VDD1.n35 15.6666
R270 VDD1.n12 VDD1.n11 12.8005
R271 VDD1.n39 VDD1.n38 12.8005
R272 VDD1.n15 VDD1.n6 12.0247
R273 VDD1.n42 VDD1.n33 12.0247
R274 VDD1.n16 VDD1.n4 11.249
R275 VDD1.n43 VDD1.n31 11.249
R276 VDD1.n20 VDD1.n19 10.4732
R277 VDD1.n47 VDD1.n46 10.4732
R278 VDD1.n23 VDD1.n2 9.69747
R279 VDD1.n50 VDD1.n29 9.69747
R280 VDD1.n26 VDD1.n25 9.45567
R281 VDD1.n53 VDD1.n52 9.45567
R282 VDD1.n25 VDD1.n24 9.3005
R283 VDD1.n2 VDD1.n1 9.3005
R284 VDD1.n19 VDD1.n18 9.3005
R285 VDD1.n17 VDD1.n16 9.3005
R286 VDD1.n6 VDD1.n5 9.3005
R287 VDD1.n11 VDD1.n10 9.3005
R288 VDD1.n52 VDD1.n51 9.3005
R289 VDD1.n29 VDD1.n28 9.3005
R290 VDD1.n46 VDD1.n45 9.3005
R291 VDD1.n44 VDD1.n43 9.3005
R292 VDD1.n33 VDD1.n32 9.3005
R293 VDD1.n38 VDD1.n37 9.3005
R294 VDD1.n24 VDD1.n0 8.92171
R295 VDD1.n51 VDD1.n27 8.92171
R296 VDD1.n26 VDD1.n0 5.04292
R297 VDD1.n53 VDD1.n27 5.04292
R298 VDD1.n10 VDD1.n9 4.38687
R299 VDD1.n37 VDD1.n36 4.38687
R300 VDD1.n24 VDD1.n23 4.26717
R301 VDD1.n51 VDD1.n50 4.26717
R302 VDD1.n56 VDD1.t4 3.64691
R303 VDD1.n56 VDD1.t3 3.64691
R304 VDD1.n54 VDD1.t2 3.64691
R305 VDD1.n54 VDD1.t1 3.64691
R306 VDD1.n20 VDD1.n2 3.49141
R307 VDD1.n47 VDD1.n29 3.49141
R308 VDD1.n19 VDD1.n4 2.71565
R309 VDD1.n46 VDD1.n31 2.71565
R310 VDD1.n16 VDD1.n15 1.93989
R311 VDD1.n43 VDD1.n42 1.93989
R312 VDD1.n12 VDD1.n6 1.16414
R313 VDD1.n39 VDD1.n33 1.16414
R314 VDD1.n11 VDD1.n8 0.388379
R315 VDD1.n38 VDD1.n35 0.388379
R316 VDD1 VDD1.n57 0.315155
R317 VDD1.n25 VDD1.n1 0.155672
R318 VDD1.n18 VDD1.n1 0.155672
R319 VDD1.n18 VDD1.n17 0.155672
R320 VDD1.n17 VDD1.n5 0.155672
R321 VDD1.n10 VDD1.n5 0.155672
R322 VDD1.n37 VDD1.n32 0.155672
R323 VDD1.n44 VDD1.n32 0.155672
R324 VDD1.n45 VDD1.n44 0.155672
R325 VDD1.n45 VDD1.n28 0.155672
R326 VDD1.n52 VDD1.n28 0.155672
R327 B.n509 B.n508 585
R328 B.n190 B.n81 585
R329 B.n189 B.n188 585
R330 B.n187 B.n186 585
R331 B.n185 B.n184 585
R332 B.n183 B.n182 585
R333 B.n181 B.n180 585
R334 B.n179 B.n178 585
R335 B.n177 B.n176 585
R336 B.n175 B.n174 585
R337 B.n173 B.n172 585
R338 B.n171 B.n170 585
R339 B.n169 B.n168 585
R340 B.n167 B.n166 585
R341 B.n165 B.n164 585
R342 B.n163 B.n162 585
R343 B.n161 B.n160 585
R344 B.n159 B.n158 585
R345 B.n157 B.n156 585
R346 B.n155 B.n154 585
R347 B.n153 B.n152 585
R348 B.n151 B.n150 585
R349 B.n149 B.n148 585
R350 B.n147 B.n146 585
R351 B.n145 B.n144 585
R352 B.n143 B.n142 585
R353 B.n141 B.n140 585
R354 B.n139 B.n138 585
R355 B.n137 B.n136 585
R356 B.n135 B.n134 585
R357 B.n133 B.n132 585
R358 B.n131 B.n130 585
R359 B.n129 B.n128 585
R360 B.n127 B.n126 585
R361 B.n125 B.n124 585
R362 B.n123 B.n122 585
R363 B.n121 B.n120 585
R364 B.n119 B.n118 585
R365 B.n117 B.n116 585
R366 B.n115 B.n114 585
R367 B.n113 B.n112 585
R368 B.n111 B.n110 585
R369 B.n109 B.n108 585
R370 B.n107 B.n106 585
R371 B.n105 B.n104 585
R372 B.n103 B.n102 585
R373 B.n101 B.n100 585
R374 B.n99 B.n98 585
R375 B.n97 B.n96 585
R376 B.n95 B.n94 585
R377 B.n93 B.n92 585
R378 B.n91 B.n90 585
R379 B.n89 B.n88 585
R380 B.n53 B.n52 585
R381 B.n507 B.n54 585
R382 B.n512 B.n54 585
R383 B.n506 B.n505 585
R384 B.n505 B.n50 585
R385 B.n504 B.n49 585
R386 B.n518 B.n49 585
R387 B.n503 B.n48 585
R388 B.n519 B.n48 585
R389 B.n502 B.n47 585
R390 B.n520 B.n47 585
R391 B.n501 B.n500 585
R392 B.n500 B.n46 585
R393 B.n499 B.n42 585
R394 B.n526 B.n42 585
R395 B.n498 B.n41 585
R396 B.n527 B.n41 585
R397 B.n497 B.n40 585
R398 B.n528 B.n40 585
R399 B.n496 B.n495 585
R400 B.n495 B.n36 585
R401 B.n494 B.n35 585
R402 B.n534 B.n35 585
R403 B.n493 B.n34 585
R404 B.n535 B.n34 585
R405 B.n492 B.n33 585
R406 B.n536 B.n33 585
R407 B.n491 B.n490 585
R408 B.n490 B.n29 585
R409 B.n489 B.n28 585
R410 B.n542 B.n28 585
R411 B.n488 B.n27 585
R412 B.n543 B.n27 585
R413 B.n487 B.n26 585
R414 B.n544 B.n26 585
R415 B.n486 B.n485 585
R416 B.n485 B.n22 585
R417 B.n484 B.n21 585
R418 B.n550 B.n21 585
R419 B.n483 B.n20 585
R420 B.n551 B.n20 585
R421 B.n482 B.n19 585
R422 B.n552 B.n19 585
R423 B.n481 B.n480 585
R424 B.n480 B.n15 585
R425 B.n479 B.n14 585
R426 B.n558 B.n14 585
R427 B.n478 B.n13 585
R428 B.n559 B.n13 585
R429 B.n477 B.n12 585
R430 B.n560 B.n12 585
R431 B.n476 B.n475 585
R432 B.n475 B.n474 585
R433 B.n473 B.n472 585
R434 B.n473 B.n8 585
R435 B.n471 B.n7 585
R436 B.n567 B.n7 585
R437 B.n470 B.n6 585
R438 B.n568 B.n6 585
R439 B.n469 B.n5 585
R440 B.n569 B.n5 585
R441 B.n468 B.n467 585
R442 B.n467 B.n4 585
R443 B.n466 B.n191 585
R444 B.n466 B.n465 585
R445 B.n456 B.n192 585
R446 B.n193 B.n192 585
R447 B.n458 B.n457 585
R448 B.n459 B.n458 585
R449 B.n455 B.n198 585
R450 B.n198 B.n197 585
R451 B.n454 B.n453 585
R452 B.n453 B.n452 585
R453 B.n200 B.n199 585
R454 B.n201 B.n200 585
R455 B.n445 B.n444 585
R456 B.n446 B.n445 585
R457 B.n443 B.n205 585
R458 B.n209 B.n205 585
R459 B.n442 B.n441 585
R460 B.n441 B.n440 585
R461 B.n207 B.n206 585
R462 B.n208 B.n207 585
R463 B.n433 B.n432 585
R464 B.n434 B.n433 585
R465 B.n431 B.n214 585
R466 B.n214 B.n213 585
R467 B.n430 B.n429 585
R468 B.n429 B.n428 585
R469 B.n216 B.n215 585
R470 B.n217 B.n216 585
R471 B.n421 B.n420 585
R472 B.n422 B.n421 585
R473 B.n419 B.n222 585
R474 B.n222 B.n221 585
R475 B.n418 B.n417 585
R476 B.n417 B.n416 585
R477 B.n224 B.n223 585
R478 B.n225 B.n224 585
R479 B.n409 B.n408 585
R480 B.n410 B.n409 585
R481 B.n407 B.n230 585
R482 B.n230 B.n229 585
R483 B.n406 B.n405 585
R484 B.n405 B.n404 585
R485 B.n232 B.n231 585
R486 B.n397 B.n232 585
R487 B.n396 B.n395 585
R488 B.n398 B.n396 585
R489 B.n394 B.n237 585
R490 B.n237 B.n236 585
R491 B.n393 B.n392 585
R492 B.n392 B.n391 585
R493 B.n239 B.n238 585
R494 B.n240 B.n239 585
R495 B.n384 B.n383 585
R496 B.n385 B.n384 585
R497 B.n243 B.n242 585
R498 B.n276 B.n274 585
R499 B.n277 B.n273 585
R500 B.n277 B.n244 585
R501 B.n280 B.n279 585
R502 B.n281 B.n272 585
R503 B.n283 B.n282 585
R504 B.n285 B.n271 585
R505 B.n288 B.n287 585
R506 B.n289 B.n270 585
R507 B.n291 B.n290 585
R508 B.n293 B.n269 585
R509 B.n296 B.n295 585
R510 B.n297 B.n268 585
R511 B.n299 B.n298 585
R512 B.n301 B.n267 585
R513 B.n304 B.n303 585
R514 B.n305 B.n266 585
R515 B.n307 B.n306 585
R516 B.n309 B.n265 585
R517 B.n312 B.n311 585
R518 B.n313 B.n264 585
R519 B.n318 B.n317 585
R520 B.n320 B.n263 585
R521 B.n323 B.n322 585
R522 B.n324 B.n262 585
R523 B.n326 B.n325 585
R524 B.n328 B.n261 585
R525 B.n331 B.n330 585
R526 B.n332 B.n260 585
R527 B.n334 B.n333 585
R528 B.n336 B.n259 585
R529 B.n339 B.n338 585
R530 B.n341 B.n256 585
R531 B.n343 B.n342 585
R532 B.n345 B.n255 585
R533 B.n348 B.n347 585
R534 B.n349 B.n254 585
R535 B.n351 B.n350 585
R536 B.n353 B.n253 585
R537 B.n356 B.n355 585
R538 B.n357 B.n252 585
R539 B.n359 B.n358 585
R540 B.n361 B.n251 585
R541 B.n364 B.n363 585
R542 B.n365 B.n250 585
R543 B.n367 B.n366 585
R544 B.n369 B.n249 585
R545 B.n372 B.n371 585
R546 B.n373 B.n248 585
R547 B.n375 B.n374 585
R548 B.n377 B.n247 585
R549 B.n378 B.n246 585
R550 B.n381 B.n380 585
R551 B.n382 B.n245 585
R552 B.n245 B.n244 585
R553 B.n387 B.n386 585
R554 B.n386 B.n385 585
R555 B.n388 B.n241 585
R556 B.n241 B.n240 585
R557 B.n390 B.n389 585
R558 B.n391 B.n390 585
R559 B.n235 B.n234 585
R560 B.n236 B.n235 585
R561 B.n400 B.n399 585
R562 B.n399 B.n398 585
R563 B.n401 B.n233 585
R564 B.n397 B.n233 585
R565 B.n403 B.n402 585
R566 B.n404 B.n403 585
R567 B.n228 B.n227 585
R568 B.n229 B.n228 585
R569 B.n412 B.n411 585
R570 B.n411 B.n410 585
R571 B.n413 B.n226 585
R572 B.n226 B.n225 585
R573 B.n415 B.n414 585
R574 B.n416 B.n415 585
R575 B.n220 B.n219 585
R576 B.n221 B.n220 585
R577 B.n424 B.n423 585
R578 B.n423 B.n422 585
R579 B.n425 B.n218 585
R580 B.n218 B.n217 585
R581 B.n427 B.n426 585
R582 B.n428 B.n427 585
R583 B.n212 B.n211 585
R584 B.n213 B.n212 585
R585 B.n436 B.n435 585
R586 B.n435 B.n434 585
R587 B.n437 B.n210 585
R588 B.n210 B.n208 585
R589 B.n439 B.n438 585
R590 B.n440 B.n439 585
R591 B.n204 B.n203 585
R592 B.n209 B.n204 585
R593 B.n448 B.n447 585
R594 B.n447 B.n446 585
R595 B.n449 B.n202 585
R596 B.n202 B.n201 585
R597 B.n451 B.n450 585
R598 B.n452 B.n451 585
R599 B.n196 B.n195 585
R600 B.n197 B.n196 585
R601 B.n461 B.n460 585
R602 B.n460 B.n459 585
R603 B.n462 B.n194 585
R604 B.n194 B.n193 585
R605 B.n464 B.n463 585
R606 B.n465 B.n464 585
R607 B.n3 B.n0 585
R608 B.n4 B.n3 585
R609 B.n566 B.n1 585
R610 B.n567 B.n566 585
R611 B.n565 B.n564 585
R612 B.n565 B.n8 585
R613 B.n563 B.n9 585
R614 B.n474 B.n9 585
R615 B.n562 B.n561 585
R616 B.n561 B.n560 585
R617 B.n11 B.n10 585
R618 B.n559 B.n11 585
R619 B.n557 B.n556 585
R620 B.n558 B.n557 585
R621 B.n555 B.n16 585
R622 B.n16 B.n15 585
R623 B.n554 B.n553 585
R624 B.n553 B.n552 585
R625 B.n18 B.n17 585
R626 B.n551 B.n18 585
R627 B.n549 B.n548 585
R628 B.n550 B.n549 585
R629 B.n547 B.n23 585
R630 B.n23 B.n22 585
R631 B.n546 B.n545 585
R632 B.n545 B.n544 585
R633 B.n25 B.n24 585
R634 B.n543 B.n25 585
R635 B.n541 B.n540 585
R636 B.n542 B.n541 585
R637 B.n539 B.n30 585
R638 B.n30 B.n29 585
R639 B.n538 B.n537 585
R640 B.n537 B.n536 585
R641 B.n32 B.n31 585
R642 B.n535 B.n32 585
R643 B.n533 B.n532 585
R644 B.n534 B.n533 585
R645 B.n531 B.n37 585
R646 B.n37 B.n36 585
R647 B.n530 B.n529 585
R648 B.n529 B.n528 585
R649 B.n39 B.n38 585
R650 B.n527 B.n39 585
R651 B.n525 B.n524 585
R652 B.n526 B.n525 585
R653 B.n523 B.n43 585
R654 B.n46 B.n43 585
R655 B.n522 B.n521 585
R656 B.n521 B.n520 585
R657 B.n45 B.n44 585
R658 B.n519 B.n45 585
R659 B.n517 B.n516 585
R660 B.n518 B.n517 585
R661 B.n515 B.n51 585
R662 B.n51 B.n50 585
R663 B.n514 B.n513 585
R664 B.n513 B.n512 585
R665 B.n570 B.n569 585
R666 B.n568 B.n2 585
R667 B.n513 B.n53 506.916
R668 B.n509 B.n54 506.916
R669 B.n384 B.n245 506.916
R670 B.n386 B.n243 506.916
R671 B.n85 B.t13 298.521
R672 B.n82 B.t17 298.521
R673 B.n257 B.t10 298.521
R674 B.n314 B.t6 298.521
R675 B.n511 B.n510 256.663
R676 B.n511 B.n80 256.663
R677 B.n511 B.n79 256.663
R678 B.n511 B.n78 256.663
R679 B.n511 B.n77 256.663
R680 B.n511 B.n76 256.663
R681 B.n511 B.n75 256.663
R682 B.n511 B.n74 256.663
R683 B.n511 B.n73 256.663
R684 B.n511 B.n72 256.663
R685 B.n511 B.n71 256.663
R686 B.n511 B.n70 256.663
R687 B.n511 B.n69 256.663
R688 B.n511 B.n68 256.663
R689 B.n511 B.n67 256.663
R690 B.n511 B.n66 256.663
R691 B.n511 B.n65 256.663
R692 B.n511 B.n64 256.663
R693 B.n511 B.n63 256.663
R694 B.n511 B.n62 256.663
R695 B.n511 B.n61 256.663
R696 B.n511 B.n60 256.663
R697 B.n511 B.n59 256.663
R698 B.n511 B.n58 256.663
R699 B.n511 B.n57 256.663
R700 B.n511 B.n56 256.663
R701 B.n511 B.n55 256.663
R702 B.n275 B.n244 256.663
R703 B.n278 B.n244 256.663
R704 B.n284 B.n244 256.663
R705 B.n286 B.n244 256.663
R706 B.n292 B.n244 256.663
R707 B.n294 B.n244 256.663
R708 B.n300 B.n244 256.663
R709 B.n302 B.n244 256.663
R710 B.n308 B.n244 256.663
R711 B.n310 B.n244 256.663
R712 B.n319 B.n244 256.663
R713 B.n321 B.n244 256.663
R714 B.n327 B.n244 256.663
R715 B.n329 B.n244 256.663
R716 B.n335 B.n244 256.663
R717 B.n337 B.n244 256.663
R718 B.n344 B.n244 256.663
R719 B.n346 B.n244 256.663
R720 B.n352 B.n244 256.663
R721 B.n354 B.n244 256.663
R722 B.n360 B.n244 256.663
R723 B.n362 B.n244 256.663
R724 B.n368 B.n244 256.663
R725 B.n370 B.n244 256.663
R726 B.n376 B.n244 256.663
R727 B.n379 B.n244 256.663
R728 B.n572 B.n571 256.663
R729 B.n82 B.t18 203.035
R730 B.n257 B.t12 203.035
R731 B.n85 B.t15 203.035
R732 B.n314 B.t9 203.035
R733 B.n83 B.t19 169.482
R734 B.n258 B.t11 169.482
R735 B.n86 B.t16 169.482
R736 B.n315 B.t8 169.482
R737 B.n90 B.n89 163.367
R738 B.n94 B.n93 163.367
R739 B.n98 B.n97 163.367
R740 B.n102 B.n101 163.367
R741 B.n106 B.n105 163.367
R742 B.n110 B.n109 163.367
R743 B.n114 B.n113 163.367
R744 B.n118 B.n117 163.367
R745 B.n122 B.n121 163.367
R746 B.n126 B.n125 163.367
R747 B.n130 B.n129 163.367
R748 B.n134 B.n133 163.367
R749 B.n138 B.n137 163.367
R750 B.n142 B.n141 163.367
R751 B.n146 B.n145 163.367
R752 B.n150 B.n149 163.367
R753 B.n154 B.n153 163.367
R754 B.n158 B.n157 163.367
R755 B.n162 B.n161 163.367
R756 B.n166 B.n165 163.367
R757 B.n170 B.n169 163.367
R758 B.n174 B.n173 163.367
R759 B.n178 B.n177 163.367
R760 B.n182 B.n181 163.367
R761 B.n186 B.n185 163.367
R762 B.n188 B.n81 163.367
R763 B.n384 B.n239 163.367
R764 B.n392 B.n239 163.367
R765 B.n392 B.n237 163.367
R766 B.n396 B.n237 163.367
R767 B.n396 B.n232 163.367
R768 B.n405 B.n232 163.367
R769 B.n405 B.n230 163.367
R770 B.n409 B.n230 163.367
R771 B.n409 B.n224 163.367
R772 B.n417 B.n224 163.367
R773 B.n417 B.n222 163.367
R774 B.n421 B.n222 163.367
R775 B.n421 B.n216 163.367
R776 B.n429 B.n216 163.367
R777 B.n429 B.n214 163.367
R778 B.n433 B.n214 163.367
R779 B.n433 B.n207 163.367
R780 B.n441 B.n207 163.367
R781 B.n441 B.n205 163.367
R782 B.n445 B.n205 163.367
R783 B.n445 B.n200 163.367
R784 B.n453 B.n200 163.367
R785 B.n453 B.n198 163.367
R786 B.n458 B.n198 163.367
R787 B.n458 B.n192 163.367
R788 B.n466 B.n192 163.367
R789 B.n467 B.n466 163.367
R790 B.n467 B.n5 163.367
R791 B.n6 B.n5 163.367
R792 B.n7 B.n6 163.367
R793 B.n473 B.n7 163.367
R794 B.n475 B.n473 163.367
R795 B.n475 B.n12 163.367
R796 B.n13 B.n12 163.367
R797 B.n14 B.n13 163.367
R798 B.n480 B.n14 163.367
R799 B.n480 B.n19 163.367
R800 B.n20 B.n19 163.367
R801 B.n21 B.n20 163.367
R802 B.n485 B.n21 163.367
R803 B.n485 B.n26 163.367
R804 B.n27 B.n26 163.367
R805 B.n28 B.n27 163.367
R806 B.n490 B.n28 163.367
R807 B.n490 B.n33 163.367
R808 B.n34 B.n33 163.367
R809 B.n35 B.n34 163.367
R810 B.n495 B.n35 163.367
R811 B.n495 B.n40 163.367
R812 B.n41 B.n40 163.367
R813 B.n42 B.n41 163.367
R814 B.n500 B.n42 163.367
R815 B.n500 B.n47 163.367
R816 B.n48 B.n47 163.367
R817 B.n49 B.n48 163.367
R818 B.n505 B.n49 163.367
R819 B.n505 B.n54 163.367
R820 B.n277 B.n276 163.367
R821 B.n279 B.n277 163.367
R822 B.n283 B.n272 163.367
R823 B.n287 B.n285 163.367
R824 B.n291 B.n270 163.367
R825 B.n295 B.n293 163.367
R826 B.n299 B.n268 163.367
R827 B.n303 B.n301 163.367
R828 B.n307 B.n266 163.367
R829 B.n311 B.n309 163.367
R830 B.n318 B.n264 163.367
R831 B.n322 B.n320 163.367
R832 B.n326 B.n262 163.367
R833 B.n330 B.n328 163.367
R834 B.n334 B.n260 163.367
R835 B.n338 B.n336 163.367
R836 B.n343 B.n256 163.367
R837 B.n347 B.n345 163.367
R838 B.n351 B.n254 163.367
R839 B.n355 B.n353 163.367
R840 B.n359 B.n252 163.367
R841 B.n363 B.n361 163.367
R842 B.n367 B.n250 163.367
R843 B.n371 B.n369 163.367
R844 B.n375 B.n248 163.367
R845 B.n378 B.n377 163.367
R846 B.n380 B.n245 163.367
R847 B.n386 B.n241 163.367
R848 B.n390 B.n241 163.367
R849 B.n390 B.n235 163.367
R850 B.n399 B.n235 163.367
R851 B.n399 B.n233 163.367
R852 B.n403 B.n233 163.367
R853 B.n403 B.n228 163.367
R854 B.n411 B.n228 163.367
R855 B.n411 B.n226 163.367
R856 B.n415 B.n226 163.367
R857 B.n415 B.n220 163.367
R858 B.n423 B.n220 163.367
R859 B.n423 B.n218 163.367
R860 B.n427 B.n218 163.367
R861 B.n427 B.n212 163.367
R862 B.n435 B.n212 163.367
R863 B.n435 B.n210 163.367
R864 B.n439 B.n210 163.367
R865 B.n439 B.n204 163.367
R866 B.n447 B.n204 163.367
R867 B.n447 B.n202 163.367
R868 B.n451 B.n202 163.367
R869 B.n451 B.n196 163.367
R870 B.n460 B.n196 163.367
R871 B.n460 B.n194 163.367
R872 B.n464 B.n194 163.367
R873 B.n464 B.n3 163.367
R874 B.n570 B.n3 163.367
R875 B.n566 B.n2 163.367
R876 B.n566 B.n565 163.367
R877 B.n565 B.n9 163.367
R878 B.n561 B.n9 163.367
R879 B.n561 B.n11 163.367
R880 B.n557 B.n11 163.367
R881 B.n557 B.n16 163.367
R882 B.n553 B.n16 163.367
R883 B.n553 B.n18 163.367
R884 B.n549 B.n18 163.367
R885 B.n549 B.n23 163.367
R886 B.n545 B.n23 163.367
R887 B.n545 B.n25 163.367
R888 B.n541 B.n25 163.367
R889 B.n541 B.n30 163.367
R890 B.n537 B.n30 163.367
R891 B.n537 B.n32 163.367
R892 B.n533 B.n32 163.367
R893 B.n533 B.n37 163.367
R894 B.n529 B.n37 163.367
R895 B.n529 B.n39 163.367
R896 B.n525 B.n39 163.367
R897 B.n525 B.n43 163.367
R898 B.n521 B.n43 163.367
R899 B.n521 B.n45 163.367
R900 B.n517 B.n45 163.367
R901 B.n517 B.n51 163.367
R902 B.n513 B.n51 163.367
R903 B.n385 B.n244 124.335
R904 B.n512 B.n511 124.335
R905 B.n55 B.n53 71.676
R906 B.n90 B.n56 71.676
R907 B.n94 B.n57 71.676
R908 B.n98 B.n58 71.676
R909 B.n102 B.n59 71.676
R910 B.n106 B.n60 71.676
R911 B.n110 B.n61 71.676
R912 B.n114 B.n62 71.676
R913 B.n118 B.n63 71.676
R914 B.n122 B.n64 71.676
R915 B.n126 B.n65 71.676
R916 B.n130 B.n66 71.676
R917 B.n134 B.n67 71.676
R918 B.n138 B.n68 71.676
R919 B.n142 B.n69 71.676
R920 B.n146 B.n70 71.676
R921 B.n150 B.n71 71.676
R922 B.n154 B.n72 71.676
R923 B.n158 B.n73 71.676
R924 B.n162 B.n74 71.676
R925 B.n166 B.n75 71.676
R926 B.n170 B.n76 71.676
R927 B.n174 B.n77 71.676
R928 B.n178 B.n78 71.676
R929 B.n182 B.n79 71.676
R930 B.n186 B.n80 71.676
R931 B.n510 B.n81 71.676
R932 B.n510 B.n509 71.676
R933 B.n188 B.n80 71.676
R934 B.n185 B.n79 71.676
R935 B.n181 B.n78 71.676
R936 B.n177 B.n77 71.676
R937 B.n173 B.n76 71.676
R938 B.n169 B.n75 71.676
R939 B.n165 B.n74 71.676
R940 B.n161 B.n73 71.676
R941 B.n157 B.n72 71.676
R942 B.n153 B.n71 71.676
R943 B.n149 B.n70 71.676
R944 B.n145 B.n69 71.676
R945 B.n141 B.n68 71.676
R946 B.n137 B.n67 71.676
R947 B.n133 B.n66 71.676
R948 B.n129 B.n65 71.676
R949 B.n125 B.n64 71.676
R950 B.n121 B.n63 71.676
R951 B.n117 B.n62 71.676
R952 B.n113 B.n61 71.676
R953 B.n109 B.n60 71.676
R954 B.n105 B.n59 71.676
R955 B.n101 B.n58 71.676
R956 B.n97 B.n57 71.676
R957 B.n93 B.n56 71.676
R958 B.n89 B.n55 71.676
R959 B.n275 B.n243 71.676
R960 B.n279 B.n278 71.676
R961 B.n284 B.n283 71.676
R962 B.n287 B.n286 71.676
R963 B.n292 B.n291 71.676
R964 B.n295 B.n294 71.676
R965 B.n300 B.n299 71.676
R966 B.n303 B.n302 71.676
R967 B.n308 B.n307 71.676
R968 B.n311 B.n310 71.676
R969 B.n319 B.n318 71.676
R970 B.n322 B.n321 71.676
R971 B.n327 B.n326 71.676
R972 B.n330 B.n329 71.676
R973 B.n335 B.n334 71.676
R974 B.n338 B.n337 71.676
R975 B.n344 B.n343 71.676
R976 B.n347 B.n346 71.676
R977 B.n352 B.n351 71.676
R978 B.n355 B.n354 71.676
R979 B.n360 B.n359 71.676
R980 B.n363 B.n362 71.676
R981 B.n368 B.n367 71.676
R982 B.n371 B.n370 71.676
R983 B.n376 B.n375 71.676
R984 B.n379 B.n378 71.676
R985 B.n276 B.n275 71.676
R986 B.n278 B.n272 71.676
R987 B.n285 B.n284 71.676
R988 B.n286 B.n270 71.676
R989 B.n293 B.n292 71.676
R990 B.n294 B.n268 71.676
R991 B.n301 B.n300 71.676
R992 B.n302 B.n266 71.676
R993 B.n309 B.n308 71.676
R994 B.n310 B.n264 71.676
R995 B.n320 B.n319 71.676
R996 B.n321 B.n262 71.676
R997 B.n328 B.n327 71.676
R998 B.n329 B.n260 71.676
R999 B.n336 B.n335 71.676
R1000 B.n337 B.n256 71.676
R1001 B.n345 B.n344 71.676
R1002 B.n346 B.n254 71.676
R1003 B.n353 B.n352 71.676
R1004 B.n354 B.n252 71.676
R1005 B.n361 B.n360 71.676
R1006 B.n362 B.n250 71.676
R1007 B.n369 B.n368 71.676
R1008 B.n370 B.n248 71.676
R1009 B.n377 B.n376 71.676
R1010 B.n380 B.n379 71.676
R1011 B.n571 B.n570 71.676
R1012 B.n571 B.n2 71.676
R1013 B.n385 B.n240 69.8744
R1014 B.n391 B.n240 69.8744
R1015 B.n391 B.n236 69.8744
R1016 B.n398 B.n236 69.8744
R1017 B.n398 B.n397 69.8744
R1018 B.n404 B.n229 69.8744
R1019 B.n410 B.n229 69.8744
R1020 B.n410 B.n225 69.8744
R1021 B.n416 B.n225 69.8744
R1022 B.n416 B.n221 69.8744
R1023 B.n422 B.n221 69.8744
R1024 B.n422 B.n217 69.8744
R1025 B.n428 B.n217 69.8744
R1026 B.n434 B.n213 69.8744
R1027 B.n434 B.n208 69.8744
R1028 B.n440 B.n208 69.8744
R1029 B.n440 B.n209 69.8744
R1030 B.n446 B.n201 69.8744
R1031 B.n452 B.n201 69.8744
R1032 B.n452 B.n197 69.8744
R1033 B.n459 B.n197 69.8744
R1034 B.n465 B.n193 69.8744
R1035 B.n465 B.n4 69.8744
R1036 B.n569 B.n4 69.8744
R1037 B.n569 B.n568 69.8744
R1038 B.n568 B.n567 69.8744
R1039 B.n567 B.n8 69.8744
R1040 B.n474 B.n8 69.8744
R1041 B.n560 B.n559 69.8744
R1042 B.n559 B.n558 69.8744
R1043 B.n558 B.n15 69.8744
R1044 B.n552 B.n15 69.8744
R1045 B.n551 B.n550 69.8744
R1046 B.n550 B.n22 69.8744
R1047 B.n544 B.n22 69.8744
R1048 B.n544 B.n543 69.8744
R1049 B.n542 B.n29 69.8744
R1050 B.n536 B.n29 69.8744
R1051 B.n536 B.n535 69.8744
R1052 B.n535 B.n534 69.8744
R1053 B.n534 B.n36 69.8744
R1054 B.n528 B.n36 69.8744
R1055 B.n528 B.n527 69.8744
R1056 B.n527 B.n526 69.8744
R1057 B.n520 B.n46 69.8744
R1058 B.n520 B.n519 69.8744
R1059 B.n519 B.n518 69.8744
R1060 B.n518 B.n50 69.8744
R1061 B.n512 B.n50 69.8744
R1062 B.n397 B.t7 61.6539
R1063 B.n46 B.t14 61.6539
R1064 B.n87 B.n86 59.5399
R1065 B.n84 B.n83 59.5399
R1066 B.n340 B.n258 59.5399
R1067 B.n316 B.n315 59.5399
R1068 B.t2 B.n213 57.5437
R1069 B.n543 B.t5 57.5437
R1070 B.n446 B.t3 51.3784
R1071 B.n552 B.t4 51.3784
R1072 B.t0 B.n193 45.213
R1073 B.n474 B.t1 45.213
R1074 B.n86 B.n85 33.552
R1075 B.n83 B.n82 33.552
R1076 B.n258 B.n257 33.552
R1077 B.n315 B.n314 33.552
R1078 B.n387 B.n242 32.9371
R1079 B.n383 B.n382 32.9371
R1080 B.n508 B.n507 32.9371
R1081 B.n514 B.n52 32.9371
R1082 B.n459 B.t0 24.6619
R1083 B.n560 B.t1 24.6619
R1084 B.n209 B.t3 18.4965
R1085 B.t4 B.n551 18.4965
R1086 B B.n572 18.0485
R1087 B.n428 B.t2 12.3312
R1088 B.t5 B.n542 12.3312
R1089 B.n388 B.n387 10.6151
R1090 B.n389 B.n388 10.6151
R1091 B.n389 B.n234 10.6151
R1092 B.n400 B.n234 10.6151
R1093 B.n401 B.n400 10.6151
R1094 B.n402 B.n401 10.6151
R1095 B.n402 B.n227 10.6151
R1096 B.n412 B.n227 10.6151
R1097 B.n413 B.n412 10.6151
R1098 B.n414 B.n413 10.6151
R1099 B.n414 B.n219 10.6151
R1100 B.n424 B.n219 10.6151
R1101 B.n425 B.n424 10.6151
R1102 B.n426 B.n425 10.6151
R1103 B.n426 B.n211 10.6151
R1104 B.n436 B.n211 10.6151
R1105 B.n437 B.n436 10.6151
R1106 B.n438 B.n437 10.6151
R1107 B.n438 B.n203 10.6151
R1108 B.n448 B.n203 10.6151
R1109 B.n449 B.n448 10.6151
R1110 B.n450 B.n449 10.6151
R1111 B.n450 B.n195 10.6151
R1112 B.n461 B.n195 10.6151
R1113 B.n462 B.n461 10.6151
R1114 B.n463 B.n462 10.6151
R1115 B.n463 B.n0 10.6151
R1116 B.n274 B.n242 10.6151
R1117 B.n274 B.n273 10.6151
R1118 B.n280 B.n273 10.6151
R1119 B.n281 B.n280 10.6151
R1120 B.n282 B.n281 10.6151
R1121 B.n282 B.n271 10.6151
R1122 B.n288 B.n271 10.6151
R1123 B.n289 B.n288 10.6151
R1124 B.n290 B.n289 10.6151
R1125 B.n290 B.n269 10.6151
R1126 B.n296 B.n269 10.6151
R1127 B.n297 B.n296 10.6151
R1128 B.n298 B.n297 10.6151
R1129 B.n298 B.n267 10.6151
R1130 B.n304 B.n267 10.6151
R1131 B.n305 B.n304 10.6151
R1132 B.n306 B.n305 10.6151
R1133 B.n306 B.n265 10.6151
R1134 B.n312 B.n265 10.6151
R1135 B.n313 B.n312 10.6151
R1136 B.n317 B.n313 10.6151
R1137 B.n323 B.n263 10.6151
R1138 B.n324 B.n323 10.6151
R1139 B.n325 B.n324 10.6151
R1140 B.n325 B.n261 10.6151
R1141 B.n331 B.n261 10.6151
R1142 B.n332 B.n331 10.6151
R1143 B.n333 B.n332 10.6151
R1144 B.n333 B.n259 10.6151
R1145 B.n339 B.n259 10.6151
R1146 B.n342 B.n341 10.6151
R1147 B.n342 B.n255 10.6151
R1148 B.n348 B.n255 10.6151
R1149 B.n349 B.n348 10.6151
R1150 B.n350 B.n349 10.6151
R1151 B.n350 B.n253 10.6151
R1152 B.n356 B.n253 10.6151
R1153 B.n357 B.n356 10.6151
R1154 B.n358 B.n357 10.6151
R1155 B.n358 B.n251 10.6151
R1156 B.n364 B.n251 10.6151
R1157 B.n365 B.n364 10.6151
R1158 B.n366 B.n365 10.6151
R1159 B.n366 B.n249 10.6151
R1160 B.n372 B.n249 10.6151
R1161 B.n373 B.n372 10.6151
R1162 B.n374 B.n373 10.6151
R1163 B.n374 B.n247 10.6151
R1164 B.n247 B.n246 10.6151
R1165 B.n381 B.n246 10.6151
R1166 B.n382 B.n381 10.6151
R1167 B.n383 B.n238 10.6151
R1168 B.n393 B.n238 10.6151
R1169 B.n394 B.n393 10.6151
R1170 B.n395 B.n394 10.6151
R1171 B.n395 B.n231 10.6151
R1172 B.n406 B.n231 10.6151
R1173 B.n407 B.n406 10.6151
R1174 B.n408 B.n407 10.6151
R1175 B.n408 B.n223 10.6151
R1176 B.n418 B.n223 10.6151
R1177 B.n419 B.n418 10.6151
R1178 B.n420 B.n419 10.6151
R1179 B.n420 B.n215 10.6151
R1180 B.n430 B.n215 10.6151
R1181 B.n431 B.n430 10.6151
R1182 B.n432 B.n431 10.6151
R1183 B.n432 B.n206 10.6151
R1184 B.n442 B.n206 10.6151
R1185 B.n443 B.n442 10.6151
R1186 B.n444 B.n443 10.6151
R1187 B.n444 B.n199 10.6151
R1188 B.n454 B.n199 10.6151
R1189 B.n455 B.n454 10.6151
R1190 B.n457 B.n455 10.6151
R1191 B.n457 B.n456 10.6151
R1192 B.n456 B.n191 10.6151
R1193 B.n468 B.n191 10.6151
R1194 B.n469 B.n468 10.6151
R1195 B.n470 B.n469 10.6151
R1196 B.n471 B.n470 10.6151
R1197 B.n472 B.n471 10.6151
R1198 B.n476 B.n472 10.6151
R1199 B.n477 B.n476 10.6151
R1200 B.n478 B.n477 10.6151
R1201 B.n479 B.n478 10.6151
R1202 B.n481 B.n479 10.6151
R1203 B.n482 B.n481 10.6151
R1204 B.n483 B.n482 10.6151
R1205 B.n484 B.n483 10.6151
R1206 B.n486 B.n484 10.6151
R1207 B.n487 B.n486 10.6151
R1208 B.n488 B.n487 10.6151
R1209 B.n489 B.n488 10.6151
R1210 B.n491 B.n489 10.6151
R1211 B.n492 B.n491 10.6151
R1212 B.n493 B.n492 10.6151
R1213 B.n494 B.n493 10.6151
R1214 B.n496 B.n494 10.6151
R1215 B.n497 B.n496 10.6151
R1216 B.n498 B.n497 10.6151
R1217 B.n499 B.n498 10.6151
R1218 B.n501 B.n499 10.6151
R1219 B.n502 B.n501 10.6151
R1220 B.n503 B.n502 10.6151
R1221 B.n504 B.n503 10.6151
R1222 B.n506 B.n504 10.6151
R1223 B.n507 B.n506 10.6151
R1224 B.n564 B.n1 10.6151
R1225 B.n564 B.n563 10.6151
R1226 B.n563 B.n562 10.6151
R1227 B.n562 B.n10 10.6151
R1228 B.n556 B.n10 10.6151
R1229 B.n556 B.n555 10.6151
R1230 B.n555 B.n554 10.6151
R1231 B.n554 B.n17 10.6151
R1232 B.n548 B.n17 10.6151
R1233 B.n548 B.n547 10.6151
R1234 B.n547 B.n546 10.6151
R1235 B.n546 B.n24 10.6151
R1236 B.n540 B.n24 10.6151
R1237 B.n540 B.n539 10.6151
R1238 B.n539 B.n538 10.6151
R1239 B.n538 B.n31 10.6151
R1240 B.n532 B.n31 10.6151
R1241 B.n532 B.n531 10.6151
R1242 B.n531 B.n530 10.6151
R1243 B.n530 B.n38 10.6151
R1244 B.n524 B.n38 10.6151
R1245 B.n524 B.n523 10.6151
R1246 B.n523 B.n522 10.6151
R1247 B.n522 B.n44 10.6151
R1248 B.n516 B.n44 10.6151
R1249 B.n516 B.n515 10.6151
R1250 B.n515 B.n514 10.6151
R1251 B.n88 B.n52 10.6151
R1252 B.n91 B.n88 10.6151
R1253 B.n92 B.n91 10.6151
R1254 B.n95 B.n92 10.6151
R1255 B.n96 B.n95 10.6151
R1256 B.n99 B.n96 10.6151
R1257 B.n100 B.n99 10.6151
R1258 B.n103 B.n100 10.6151
R1259 B.n104 B.n103 10.6151
R1260 B.n107 B.n104 10.6151
R1261 B.n108 B.n107 10.6151
R1262 B.n111 B.n108 10.6151
R1263 B.n112 B.n111 10.6151
R1264 B.n115 B.n112 10.6151
R1265 B.n116 B.n115 10.6151
R1266 B.n119 B.n116 10.6151
R1267 B.n120 B.n119 10.6151
R1268 B.n123 B.n120 10.6151
R1269 B.n124 B.n123 10.6151
R1270 B.n127 B.n124 10.6151
R1271 B.n128 B.n127 10.6151
R1272 B.n132 B.n131 10.6151
R1273 B.n135 B.n132 10.6151
R1274 B.n136 B.n135 10.6151
R1275 B.n139 B.n136 10.6151
R1276 B.n140 B.n139 10.6151
R1277 B.n143 B.n140 10.6151
R1278 B.n144 B.n143 10.6151
R1279 B.n147 B.n144 10.6151
R1280 B.n148 B.n147 10.6151
R1281 B.n152 B.n151 10.6151
R1282 B.n155 B.n152 10.6151
R1283 B.n156 B.n155 10.6151
R1284 B.n159 B.n156 10.6151
R1285 B.n160 B.n159 10.6151
R1286 B.n163 B.n160 10.6151
R1287 B.n164 B.n163 10.6151
R1288 B.n167 B.n164 10.6151
R1289 B.n168 B.n167 10.6151
R1290 B.n171 B.n168 10.6151
R1291 B.n172 B.n171 10.6151
R1292 B.n175 B.n172 10.6151
R1293 B.n176 B.n175 10.6151
R1294 B.n179 B.n176 10.6151
R1295 B.n180 B.n179 10.6151
R1296 B.n183 B.n180 10.6151
R1297 B.n184 B.n183 10.6151
R1298 B.n187 B.n184 10.6151
R1299 B.n189 B.n187 10.6151
R1300 B.n190 B.n189 10.6151
R1301 B.n508 B.n190 10.6151
R1302 B.n317 B.n316 9.36635
R1303 B.n341 B.n340 9.36635
R1304 B.n128 B.n87 9.36635
R1305 B.n151 B.n84 9.36635
R1306 B.n404 B.t7 8.22096
R1307 B.n526 B.t14 8.22096
R1308 B.n572 B.n0 8.11757
R1309 B.n572 B.n1 8.11757
R1310 B.n316 B.n263 1.24928
R1311 B.n340 B.n339 1.24928
R1312 B.n131 B.n87 1.24928
R1313 B.n148 B.n84 1.24928
R1314 VN.n9 VN.n8 174.512
R1315 VN.n19 VN.n18 174.512
R1316 VN.n17 VN.n10 161.3
R1317 VN.n16 VN.n15 161.3
R1318 VN.n14 VN.n11 161.3
R1319 VN.n7 VN.n0 161.3
R1320 VN.n6 VN.n5 161.3
R1321 VN.n4 VN.n1 161.3
R1322 VN.n3 VN.t3 128.267
R1323 VN.n13 VN.t4 128.267
R1324 VN.n2 VN.t1 93.4741
R1325 VN.n8 VN.t2 93.4741
R1326 VN.n12 VN.t5 93.4741
R1327 VN.n18 VN.t0 93.4741
R1328 VN.n6 VN.n1 53.6055
R1329 VN.n16 VN.n11 53.6055
R1330 VN.n3 VN.n2 41.8065
R1331 VN.n13 VN.n12 41.8065
R1332 VN VN.n19 39.2941
R1333 VN.n7 VN.n6 27.3813
R1334 VN.n17 VN.n16 27.3813
R1335 VN.n2 VN.n1 24.4675
R1336 VN.n12 VN.n11 24.4675
R1337 VN.n14 VN.n13 17.6362
R1338 VN.n4 VN.n3 17.6362
R1339 VN.n8 VN.n7 11.2553
R1340 VN.n18 VN.n17 11.2553
R1341 VN.n19 VN.n10 0.189894
R1342 VN.n15 VN.n10 0.189894
R1343 VN.n15 VN.n14 0.189894
R1344 VN.n5 VN.n4 0.189894
R1345 VN.n5 VN.n0 0.189894
R1346 VN.n9 VN.n0 0.189894
R1347 VN VN.n9 0.0516364
R1348 VDD2.n51 VDD2.n29 289.615
R1349 VDD2.n22 VDD2.n0 289.615
R1350 VDD2.n52 VDD2.n51 185
R1351 VDD2.n50 VDD2.n49 185
R1352 VDD2.n33 VDD2.n32 185
R1353 VDD2.n44 VDD2.n43 185
R1354 VDD2.n42 VDD2.n41 185
R1355 VDD2.n37 VDD2.n36 185
R1356 VDD2.n8 VDD2.n7 185
R1357 VDD2.n13 VDD2.n12 185
R1358 VDD2.n15 VDD2.n14 185
R1359 VDD2.n4 VDD2.n3 185
R1360 VDD2.n21 VDD2.n20 185
R1361 VDD2.n23 VDD2.n22 185
R1362 VDD2.n38 VDD2.t5 147.672
R1363 VDD2.n9 VDD2.t2 147.672
R1364 VDD2.n51 VDD2.n50 104.615
R1365 VDD2.n50 VDD2.n32 104.615
R1366 VDD2.n43 VDD2.n32 104.615
R1367 VDD2.n43 VDD2.n42 104.615
R1368 VDD2.n42 VDD2.n36 104.615
R1369 VDD2.n13 VDD2.n7 104.615
R1370 VDD2.n14 VDD2.n13 104.615
R1371 VDD2.n14 VDD2.n3 104.615
R1372 VDD2.n21 VDD2.n3 104.615
R1373 VDD2.n22 VDD2.n21 104.615
R1374 VDD2.n28 VDD2.n27 71.8817
R1375 VDD2 VDD2.n57 71.8788
R1376 VDD2.n28 VDD2.n26 52.8364
R1377 VDD2.t5 VDD2.n36 52.3082
R1378 VDD2.t2 VDD2.n7 52.3082
R1379 VDD2.n56 VDD2.n55 51.7732
R1380 VDD2.n56 VDD2.n28 33.2433
R1381 VDD2.n38 VDD2.n37 15.6666
R1382 VDD2.n9 VDD2.n8 15.6666
R1383 VDD2.n41 VDD2.n40 12.8005
R1384 VDD2.n12 VDD2.n11 12.8005
R1385 VDD2.n44 VDD2.n35 12.0247
R1386 VDD2.n15 VDD2.n6 12.0247
R1387 VDD2.n45 VDD2.n33 11.249
R1388 VDD2.n16 VDD2.n4 11.249
R1389 VDD2.n49 VDD2.n48 10.4732
R1390 VDD2.n20 VDD2.n19 10.4732
R1391 VDD2.n52 VDD2.n31 9.69747
R1392 VDD2.n23 VDD2.n2 9.69747
R1393 VDD2.n55 VDD2.n54 9.45567
R1394 VDD2.n26 VDD2.n25 9.45567
R1395 VDD2.n54 VDD2.n53 9.3005
R1396 VDD2.n31 VDD2.n30 9.3005
R1397 VDD2.n48 VDD2.n47 9.3005
R1398 VDD2.n46 VDD2.n45 9.3005
R1399 VDD2.n35 VDD2.n34 9.3005
R1400 VDD2.n40 VDD2.n39 9.3005
R1401 VDD2.n25 VDD2.n24 9.3005
R1402 VDD2.n2 VDD2.n1 9.3005
R1403 VDD2.n19 VDD2.n18 9.3005
R1404 VDD2.n17 VDD2.n16 9.3005
R1405 VDD2.n6 VDD2.n5 9.3005
R1406 VDD2.n11 VDD2.n10 9.3005
R1407 VDD2.n53 VDD2.n29 8.92171
R1408 VDD2.n24 VDD2.n0 8.92171
R1409 VDD2.n55 VDD2.n29 5.04292
R1410 VDD2.n26 VDD2.n0 5.04292
R1411 VDD2.n39 VDD2.n38 4.38687
R1412 VDD2.n10 VDD2.n9 4.38687
R1413 VDD2.n53 VDD2.n52 4.26717
R1414 VDD2.n24 VDD2.n23 4.26717
R1415 VDD2.n57 VDD2.t0 3.64691
R1416 VDD2.n57 VDD2.t1 3.64691
R1417 VDD2.n27 VDD2.t4 3.64691
R1418 VDD2.n27 VDD2.t3 3.64691
R1419 VDD2.n49 VDD2.n31 3.49141
R1420 VDD2.n20 VDD2.n2 3.49141
R1421 VDD2.n48 VDD2.n33 2.71565
R1422 VDD2.n19 VDD2.n4 2.71565
R1423 VDD2.n45 VDD2.n44 1.93989
R1424 VDD2.n16 VDD2.n15 1.93989
R1425 VDD2 VDD2.n56 1.17722
R1426 VDD2.n41 VDD2.n35 1.16414
R1427 VDD2.n12 VDD2.n6 1.16414
R1428 VDD2.n40 VDD2.n37 0.388379
R1429 VDD2.n11 VDD2.n8 0.388379
R1430 VDD2.n54 VDD2.n30 0.155672
R1431 VDD2.n47 VDD2.n30 0.155672
R1432 VDD2.n47 VDD2.n46 0.155672
R1433 VDD2.n46 VDD2.n34 0.155672
R1434 VDD2.n39 VDD2.n34 0.155672
R1435 VDD2.n10 VDD2.n5 0.155672
R1436 VDD2.n17 VDD2.n5 0.155672
R1437 VDD2.n18 VDD2.n17 0.155672
R1438 VDD2.n18 VDD2.n1 0.155672
R1439 VDD2.n25 VDD2.n1 0.155672
C0 VDD2 VN 2.8002f
C1 VDD1 VDD2 0.968262f
C2 VTAIL VP 3.0525f
C3 VTAIL VN 3.03824f
C4 VTAIL VDD1 4.98686f
C5 VTAIL VDD2 5.03028f
C6 VP VN 4.5444f
C7 VDD1 VP 3.005f
C8 VDD2 VP 0.359807f
C9 VDD1 VN 0.149102f
C10 VDD2 B 3.851791f
C11 VDD1 B 3.926753f
C12 VTAIL B 4.238941f
C13 VN B 8.76787f
C14 VP B 7.319204f
C15 VDD2.n0 B 0.032682f
C16 VDD2.n1 B 0.022085f
C17 VDD2.n2 B 0.011868f
C18 VDD2.n3 B 0.028051f
C19 VDD2.n4 B 0.012566f
C20 VDD2.n5 B 0.022085f
C21 VDD2.n6 B 0.011868f
C22 VDD2.n7 B 0.021038f
C23 VDD2.n8 B 0.016566f
C24 VDD2.t2 B 0.045889f
C25 VDD2.n9 B 0.091773f
C26 VDD2.n10 B 0.46717f
C27 VDD2.n11 B 0.011868f
C28 VDD2.n12 B 0.012566f
C29 VDD2.n13 B 0.028051f
C30 VDD2.n14 B 0.028051f
C31 VDD2.n15 B 0.012566f
C32 VDD2.n16 B 0.011868f
C33 VDD2.n17 B 0.022085f
C34 VDD2.n18 B 0.022085f
C35 VDD2.n19 B 0.011868f
C36 VDD2.n20 B 0.012566f
C37 VDD2.n21 B 0.028051f
C38 VDD2.n22 B 0.063624f
C39 VDD2.n23 B 0.012566f
C40 VDD2.n24 B 0.011868f
C41 VDD2.n25 B 0.055574f
C42 VDD2.n26 B 0.053689f
C43 VDD2.t4 B 0.094766f
C44 VDD2.t3 B 0.094766f
C45 VDD2.n27 B 0.782161f
C46 VDD2.n28 B 1.55787f
C47 VDD2.n29 B 0.032682f
C48 VDD2.n30 B 0.022085f
C49 VDD2.n31 B 0.011868f
C50 VDD2.n32 B 0.028051f
C51 VDD2.n33 B 0.012566f
C52 VDD2.n34 B 0.022085f
C53 VDD2.n35 B 0.011868f
C54 VDD2.n36 B 0.021038f
C55 VDD2.n37 B 0.016566f
C56 VDD2.t5 B 0.045889f
C57 VDD2.n38 B 0.091773f
C58 VDD2.n39 B 0.46717f
C59 VDD2.n40 B 0.011868f
C60 VDD2.n41 B 0.012566f
C61 VDD2.n42 B 0.028051f
C62 VDD2.n43 B 0.028051f
C63 VDD2.n44 B 0.012566f
C64 VDD2.n45 B 0.011868f
C65 VDD2.n46 B 0.022085f
C66 VDD2.n47 B 0.022085f
C67 VDD2.n48 B 0.011868f
C68 VDD2.n49 B 0.012566f
C69 VDD2.n50 B 0.028051f
C70 VDD2.n51 B 0.063624f
C71 VDD2.n52 B 0.012566f
C72 VDD2.n53 B 0.011868f
C73 VDD2.n54 B 0.055574f
C74 VDD2.n55 B 0.051249f
C75 VDD2.n56 B 1.51672f
C76 VDD2.t0 B 0.094766f
C77 VDD2.t1 B 0.094766f
C78 VDD2.n57 B 0.78214f
C79 VN.n0 B 0.035918f
C80 VN.t2 B 0.718231f
C81 VN.n1 B 0.063349f
C82 VN.t3 B 0.832271f
C83 VN.t1 B 0.718231f
C84 VN.n2 B 0.369648f
C85 VN.n3 B 0.354089f
C86 VN.n4 B 0.225333f
C87 VN.n5 B 0.035918f
C88 VN.n6 B 0.03843f
C89 VN.n7 B 0.05219f
C90 VN.n8 B 0.357934f
C91 VN.n9 B 0.033554f
C92 VN.n10 B 0.035918f
C93 VN.t0 B 0.718231f
C94 VN.n11 B 0.063349f
C95 VN.t4 B 0.832271f
C96 VN.t5 B 0.718231f
C97 VN.n12 B 0.369648f
C98 VN.n13 B 0.354089f
C99 VN.n14 B 0.225333f
C100 VN.n15 B 0.035918f
C101 VN.n16 B 0.03843f
C102 VN.n17 B 0.05219f
C103 VN.n18 B 0.357934f
C104 VN.n19 B 1.33032f
C105 VDD1.n0 B 0.033173f
C106 VDD1.n1 B 0.022417f
C107 VDD1.n2 B 0.012046f
C108 VDD1.n3 B 0.028472f
C109 VDD1.n4 B 0.012755f
C110 VDD1.n5 B 0.022417f
C111 VDD1.n6 B 0.012046f
C112 VDD1.n7 B 0.021354f
C113 VDD1.n8 B 0.016815f
C114 VDD1.t5 B 0.046579f
C115 VDD1.n9 B 0.093152f
C116 VDD1.n10 B 0.47419f
C117 VDD1.n11 B 0.012046f
C118 VDD1.n12 B 0.012755f
C119 VDD1.n13 B 0.028472f
C120 VDD1.n14 B 0.028472f
C121 VDD1.n15 B 0.012755f
C122 VDD1.n16 B 0.012046f
C123 VDD1.n17 B 0.022417f
C124 VDD1.n18 B 0.022417f
C125 VDD1.n19 B 0.012046f
C126 VDD1.n20 B 0.012755f
C127 VDD1.n21 B 0.028472f
C128 VDD1.n22 B 0.06458f
C129 VDD1.n23 B 0.012755f
C130 VDD1.n24 B 0.012046f
C131 VDD1.n25 B 0.056409f
C132 VDD1.n26 B 0.054925f
C133 VDD1.n27 B 0.033173f
C134 VDD1.n28 B 0.022417f
C135 VDD1.n29 B 0.012046f
C136 VDD1.n30 B 0.028472f
C137 VDD1.n31 B 0.012755f
C138 VDD1.n32 B 0.022417f
C139 VDD1.n33 B 0.012046f
C140 VDD1.n34 B 0.021354f
C141 VDD1.n35 B 0.016815f
C142 VDD1.t0 B 0.046579f
C143 VDD1.n36 B 0.093152f
C144 VDD1.n37 B 0.47419f
C145 VDD1.n38 B 0.012046f
C146 VDD1.n39 B 0.012755f
C147 VDD1.n40 B 0.028472f
C148 VDD1.n41 B 0.028472f
C149 VDD1.n42 B 0.012755f
C150 VDD1.n43 B 0.012046f
C151 VDD1.n44 B 0.022417f
C152 VDD1.n45 B 0.022417f
C153 VDD1.n46 B 0.012046f
C154 VDD1.n47 B 0.012755f
C155 VDD1.n48 B 0.028472f
C156 VDD1.n49 B 0.06458f
C157 VDD1.n50 B 0.012755f
C158 VDD1.n51 B 0.012046f
C159 VDD1.n52 B 0.056409f
C160 VDD1.n53 B 0.054495f
C161 VDD1.t2 B 0.09619f
C162 VDD1.t1 B 0.09619f
C163 VDD1.n54 B 0.793913f
C164 VDD1.n55 B 1.66147f
C165 VDD1.t4 B 0.09619f
C166 VDD1.t3 B 0.09619f
C167 VDD1.n56 B 0.792495f
C168 VDD1.n57 B 1.73062f
C169 VTAIL.t1 B 0.112357f
C170 VTAIL.t4 B 0.112357f
C171 VTAIL.n0 B 0.863378f
C172 VTAIL.n1 B 0.375674f
C173 VTAIL.n2 B 0.038748f
C174 VTAIL.n3 B 0.026185f
C175 VTAIL.n4 B 0.01407f
C176 VTAIL.n5 B 0.033257f
C177 VTAIL.n6 B 0.014898f
C178 VTAIL.n7 B 0.026185f
C179 VTAIL.n8 B 0.01407f
C180 VTAIL.n9 B 0.024943f
C181 VTAIL.n10 B 0.019641f
C182 VTAIL.t11 B 0.054407f
C183 VTAIL.n11 B 0.108808f
C184 VTAIL.n12 B 0.553886f
C185 VTAIL.n13 B 0.01407f
C186 VTAIL.n14 B 0.014898f
C187 VTAIL.n15 B 0.033257f
C188 VTAIL.n16 B 0.033257f
C189 VTAIL.n17 B 0.014898f
C190 VTAIL.n18 B 0.01407f
C191 VTAIL.n19 B 0.026185f
C192 VTAIL.n20 B 0.026185f
C193 VTAIL.n21 B 0.01407f
C194 VTAIL.n22 B 0.014898f
C195 VTAIL.n23 B 0.033257f
C196 VTAIL.n24 B 0.075433f
C197 VTAIL.n25 B 0.014898f
C198 VTAIL.n26 B 0.01407f
C199 VTAIL.n27 B 0.06589f
C200 VTAIL.n28 B 0.04272f
C201 VTAIL.n29 B 0.253786f
C202 VTAIL.t6 B 0.112357f
C203 VTAIL.t7 B 0.112357f
C204 VTAIL.n30 B 0.863378f
C205 VTAIL.n31 B 1.36488f
C206 VTAIL.t2 B 0.112357f
C207 VTAIL.t3 B 0.112357f
C208 VTAIL.n32 B 0.863383f
C209 VTAIL.n33 B 1.36488f
C210 VTAIL.n34 B 0.038748f
C211 VTAIL.n35 B 0.026185f
C212 VTAIL.n36 B 0.01407f
C213 VTAIL.n37 B 0.033257f
C214 VTAIL.n38 B 0.014898f
C215 VTAIL.n39 B 0.026185f
C216 VTAIL.n40 B 0.01407f
C217 VTAIL.n41 B 0.024943f
C218 VTAIL.n42 B 0.019641f
C219 VTAIL.t0 B 0.054407f
C220 VTAIL.n43 B 0.108808f
C221 VTAIL.n44 B 0.553886f
C222 VTAIL.n45 B 0.01407f
C223 VTAIL.n46 B 0.014898f
C224 VTAIL.n47 B 0.033257f
C225 VTAIL.n48 B 0.033257f
C226 VTAIL.n49 B 0.014898f
C227 VTAIL.n50 B 0.01407f
C228 VTAIL.n51 B 0.026185f
C229 VTAIL.n52 B 0.026185f
C230 VTAIL.n53 B 0.01407f
C231 VTAIL.n54 B 0.014898f
C232 VTAIL.n55 B 0.033257f
C233 VTAIL.n56 B 0.075433f
C234 VTAIL.n57 B 0.014898f
C235 VTAIL.n58 B 0.01407f
C236 VTAIL.n59 B 0.06589f
C237 VTAIL.n60 B 0.04272f
C238 VTAIL.n61 B 0.253786f
C239 VTAIL.t8 B 0.112357f
C240 VTAIL.t10 B 0.112357f
C241 VTAIL.n62 B 0.863383f
C242 VTAIL.n63 B 0.465133f
C243 VTAIL.n64 B 0.038748f
C244 VTAIL.n65 B 0.026185f
C245 VTAIL.n66 B 0.01407f
C246 VTAIL.n67 B 0.033257f
C247 VTAIL.n68 B 0.014898f
C248 VTAIL.n69 B 0.026185f
C249 VTAIL.n70 B 0.01407f
C250 VTAIL.n71 B 0.024943f
C251 VTAIL.n72 B 0.019641f
C252 VTAIL.t9 B 0.054407f
C253 VTAIL.n73 B 0.108808f
C254 VTAIL.n74 B 0.553886f
C255 VTAIL.n75 B 0.01407f
C256 VTAIL.n76 B 0.014898f
C257 VTAIL.n77 B 0.033257f
C258 VTAIL.n78 B 0.033257f
C259 VTAIL.n79 B 0.014898f
C260 VTAIL.n80 B 0.01407f
C261 VTAIL.n81 B 0.026185f
C262 VTAIL.n82 B 0.026185f
C263 VTAIL.n83 B 0.01407f
C264 VTAIL.n84 B 0.014898f
C265 VTAIL.n85 B 0.033257f
C266 VTAIL.n86 B 0.075433f
C267 VTAIL.n87 B 0.014898f
C268 VTAIL.n88 B 0.01407f
C269 VTAIL.n89 B 0.06589f
C270 VTAIL.n90 B 0.04272f
C271 VTAIL.n91 B 1.0277f
C272 VTAIL.n92 B 0.038748f
C273 VTAIL.n93 B 0.026185f
C274 VTAIL.n94 B 0.01407f
C275 VTAIL.n95 B 0.033257f
C276 VTAIL.n96 B 0.014898f
C277 VTAIL.n97 B 0.026185f
C278 VTAIL.n98 B 0.01407f
C279 VTAIL.n99 B 0.024943f
C280 VTAIL.n100 B 0.019641f
C281 VTAIL.t5 B 0.054407f
C282 VTAIL.n101 B 0.108808f
C283 VTAIL.n102 B 0.553886f
C284 VTAIL.n103 B 0.01407f
C285 VTAIL.n104 B 0.014898f
C286 VTAIL.n105 B 0.033257f
C287 VTAIL.n106 B 0.033257f
C288 VTAIL.n107 B 0.014898f
C289 VTAIL.n108 B 0.01407f
C290 VTAIL.n109 B 0.026185f
C291 VTAIL.n110 B 0.026185f
C292 VTAIL.n111 B 0.01407f
C293 VTAIL.n112 B 0.014898f
C294 VTAIL.n113 B 0.033257f
C295 VTAIL.n114 B 0.075433f
C296 VTAIL.n115 B 0.014898f
C297 VTAIL.n116 B 0.01407f
C298 VTAIL.n117 B 0.06589f
C299 VTAIL.n118 B 0.04272f
C300 VTAIL.n119 B 0.99133f
C301 VP.n0 B 0.037146f
C302 VP.t4 B 0.742792f
C303 VP.n1 B 0.065515f
C304 VP.n2 B 0.037146f
C305 VP.t3 B 0.742792f
C306 VP.n3 B 0.053975f
C307 VP.n4 B 0.037146f
C308 VP.t2 B 0.742792f
C309 VP.n5 B 0.065515f
C310 VP.t0 B 0.860732f
C311 VP.t1 B 0.742792f
C312 VP.n6 B 0.382288f
C313 VP.n7 B 0.366198f
C314 VP.n8 B 0.233038f
C315 VP.n9 B 0.037146f
C316 VP.n10 B 0.039744f
C317 VP.n11 B 0.053975f
C318 VP.n12 B 0.370174f
C319 VP.n13 B 1.3513f
C320 VP.t5 B 0.742792f
C321 VP.n14 B 0.370174f
C322 VP.n15 B 1.38562f
C323 VP.n16 B 0.037146f
C324 VP.n17 B 0.037146f
C325 VP.n18 B 0.039744f
C326 VP.n19 B 0.065515f
C327 VP.n20 B 0.333022f
C328 VP.n21 B 0.037146f
C329 VP.n22 B 0.037146f
C330 VP.n23 B 0.037146f
C331 VP.n24 B 0.039744f
C332 VP.n25 B 0.053975f
C333 VP.n26 B 0.370174f
C334 VP.n27 B 0.034701f
.ends

