* NGSPICE file created from diff_pair_sample_0080.ext - technology: sky130A

.subckt diff_pair_sample_0080 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=5.0661 ps=26.76 w=12.99 l=1.66
X1 VDD2.t1 VN.t0 VTAIL.t1 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=5.0661 ps=26.76 w=12.99 l=1.66
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=5.0661 ps=26.76 w=12.99 l=1.66
X3 VDD2.t0 VN.t1 VTAIL.t0 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=5.0661 ps=26.76 w=12.99 l=1.66
X4 B.t11 B.t9 B.t10 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=0 ps=0 w=12.99 l=1.66
X5 B.t8 B.t6 B.t7 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=0 ps=0 w=12.99 l=1.66
X6 B.t5 B.t3 B.t4 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=0 ps=0 w=12.99 l=1.66
X7 B.t2 B.t0 B.t1 w_n1766_n3566# sky130_fd_pr__pfet_01v8 ad=5.0661 pd=26.76 as=0 ps=0 w=12.99 l=1.66
R0 VP.n0 VP.t0 290.365
R1 VP.n0 VP.t1 247.452
R2 VP VP.n0 0.241678
R3 VTAIL.n1 VTAIL.t0 61.0424
R4 VTAIL.n3 VTAIL.t1 61.0412
R5 VTAIL.n0 VTAIL.t2 61.0412
R6 VTAIL.n2 VTAIL.t3 61.0412
R7 VTAIL.n1 VTAIL.n0 26.9962
R8 VTAIL.n3 VTAIL.n2 25.2807
R9 VTAIL.n2 VTAIL.n1 1.32809
R10 VTAIL VTAIL.n0 0.957397
R11 VTAIL VTAIL.n3 0.37119
R12 VDD1 VDD1.t0 116.963
R13 VDD1 VDD1.t1 78.2081
R14 VN VN.t1 290.555
R15 VN VN.t0 247.692
R16 VDD2.n0 VDD2.t1 116.008
R17 VDD2.n0 VDD2.t0 77.721
R18 VDD2 VDD2.n0 0.487569
R19 B.n391 B.n66 585
R20 B.n393 B.n392 585
R21 B.n394 B.n65 585
R22 B.n396 B.n395 585
R23 B.n397 B.n64 585
R24 B.n399 B.n398 585
R25 B.n400 B.n63 585
R26 B.n402 B.n401 585
R27 B.n403 B.n62 585
R28 B.n405 B.n404 585
R29 B.n406 B.n61 585
R30 B.n408 B.n407 585
R31 B.n409 B.n60 585
R32 B.n411 B.n410 585
R33 B.n412 B.n59 585
R34 B.n414 B.n413 585
R35 B.n415 B.n58 585
R36 B.n417 B.n416 585
R37 B.n418 B.n57 585
R38 B.n420 B.n419 585
R39 B.n421 B.n56 585
R40 B.n423 B.n422 585
R41 B.n424 B.n55 585
R42 B.n426 B.n425 585
R43 B.n427 B.n54 585
R44 B.n429 B.n428 585
R45 B.n430 B.n53 585
R46 B.n432 B.n431 585
R47 B.n433 B.n52 585
R48 B.n435 B.n434 585
R49 B.n436 B.n51 585
R50 B.n438 B.n437 585
R51 B.n439 B.n50 585
R52 B.n441 B.n440 585
R53 B.n442 B.n49 585
R54 B.n444 B.n443 585
R55 B.n445 B.n48 585
R56 B.n447 B.n446 585
R57 B.n448 B.n47 585
R58 B.n450 B.n449 585
R59 B.n451 B.n46 585
R60 B.n453 B.n452 585
R61 B.n454 B.n45 585
R62 B.n456 B.n455 585
R63 B.n457 B.n42 585
R64 B.n460 B.n459 585
R65 B.n461 B.n41 585
R66 B.n463 B.n462 585
R67 B.n464 B.n40 585
R68 B.n466 B.n465 585
R69 B.n467 B.n39 585
R70 B.n469 B.n468 585
R71 B.n470 B.n35 585
R72 B.n472 B.n471 585
R73 B.n473 B.n34 585
R74 B.n475 B.n474 585
R75 B.n476 B.n33 585
R76 B.n478 B.n477 585
R77 B.n479 B.n32 585
R78 B.n481 B.n480 585
R79 B.n482 B.n31 585
R80 B.n484 B.n483 585
R81 B.n485 B.n30 585
R82 B.n487 B.n486 585
R83 B.n488 B.n29 585
R84 B.n490 B.n489 585
R85 B.n491 B.n28 585
R86 B.n493 B.n492 585
R87 B.n494 B.n27 585
R88 B.n496 B.n495 585
R89 B.n497 B.n26 585
R90 B.n499 B.n498 585
R91 B.n500 B.n25 585
R92 B.n502 B.n501 585
R93 B.n503 B.n24 585
R94 B.n505 B.n504 585
R95 B.n506 B.n23 585
R96 B.n508 B.n507 585
R97 B.n509 B.n22 585
R98 B.n511 B.n510 585
R99 B.n512 B.n21 585
R100 B.n514 B.n513 585
R101 B.n515 B.n20 585
R102 B.n517 B.n516 585
R103 B.n518 B.n19 585
R104 B.n520 B.n519 585
R105 B.n521 B.n18 585
R106 B.n523 B.n522 585
R107 B.n524 B.n17 585
R108 B.n526 B.n525 585
R109 B.n527 B.n16 585
R110 B.n529 B.n528 585
R111 B.n530 B.n15 585
R112 B.n532 B.n531 585
R113 B.n533 B.n14 585
R114 B.n535 B.n534 585
R115 B.n536 B.n13 585
R116 B.n538 B.n537 585
R117 B.n539 B.n12 585
R118 B.n390 B.n389 585
R119 B.n388 B.n67 585
R120 B.n387 B.n386 585
R121 B.n385 B.n68 585
R122 B.n384 B.n383 585
R123 B.n382 B.n69 585
R124 B.n381 B.n380 585
R125 B.n379 B.n70 585
R126 B.n378 B.n377 585
R127 B.n376 B.n71 585
R128 B.n375 B.n374 585
R129 B.n373 B.n72 585
R130 B.n372 B.n371 585
R131 B.n370 B.n73 585
R132 B.n369 B.n368 585
R133 B.n367 B.n74 585
R134 B.n366 B.n365 585
R135 B.n364 B.n75 585
R136 B.n363 B.n362 585
R137 B.n361 B.n76 585
R138 B.n360 B.n359 585
R139 B.n358 B.n77 585
R140 B.n357 B.n356 585
R141 B.n355 B.n78 585
R142 B.n354 B.n353 585
R143 B.n352 B.n79 585
R144 B.n351 B.n350 585
R145 B.n349 B.n80 585
R146 B.n348 B.n347 585
R147 B.n346 B.n81 585
R148 B.n345 B.n344 585
R149 B.n343 B.n82 585
R150 B.n342 B.n341 585
R151 B.n340 B.n83 585
R152 B.n339 B.n338 585
R153 B.n337 B.n84 585
R154 B.n336 B.n335 585
R155 B.n334 B.n85 585
R156 B.n333 B.n332 585
R157 B.n331 B.n86 585
R158 B.n330 B.n329 585
R159 B.n177 B.n138 585
R160 B.n179 B.n178 585
R161 B.n180 B.n137 585
R162 B.n182 B.n181 585
R163 B.n183 B.n136 585
R164 B.n185 B.n184 585
R165 B.n186 B.n135 585
R166 B.n188 B.n187 585
R167 B.n189 B.n134 585
R168 B.n191 B.n190 585
R169 B.n192 B.n133 585
R170 B.n194 B.n193 585
R171 B.n195 B.n132 585
R172 B.n197 B.n196 585
R173 B.n198 B.n131 585
R174 B.n200 B.n199 585
R175 B.n201 B.n130 585
R176 B.n203 B.n202 585
R177 B.n204 B.n129 585
R178 B.n206 B.n205 585
R179 B.n207 B.n128 585
R180 B.n209 B.n208 585
R181 B.n210 B.n127 585
R182 B.n212 B.n211 585
R183 B.n213 B.n126 585
R184 B.n215 B.n214 585
R185 B.n216 B.n125 585
R186 B.n218 B.n217 585
R187 B.n219 B.n124 585
R188 B.n221 B.n220 585
R189 B.n222 B.n123 585
R190 B.n224 B.n223 585
R191 B.n225 B.n122 585
R192 B.n227 B.n226 585
R193 B.n228 B.n121 585
R194 B.n230 B.n229 585
R195 B.n231 B.n120 585
R196 B.n233 B.n232 585
R197 B.n234 B.n119 585
R198 B.n236 B.n235 585
R199 B.n237 B.n118 585
R200 B.n239 B.n238 585
R201 B.n240 B.n117 585
R202 B.n242 B.n241 585
R203 B.n243 B.n114 585
R204 B.n246 B.n245 585
R205 B.n247 B.n113 585
R206 B.n249 B.n248 585
R207 B.n250 B.n112 585
R208 B.n252 B.n251 585
R209 B.n253 B.n111 585
R210 B.n255 B.n254 585
R211 B.n256 B.n110 585
R212 B.n261 B.n260 585
R213 B.n262 B.n109 585
R214 B.n264 B.n263 585
R215 B.n265 B.n108 585
R216 B.n267 B.n266 585
R217 B.n268 B.n107 585
R218 B.n270 B.n269 585
R219 B.n271 B.n106 585
R220 B.n273 B.n272 585
R221 B.n274 B.n105 585
R222 B.n276 B.n275 585
R223 B.n277 B.n104 585
R224 B.n279 B.n278 585
R225 B.n280 B.n103 585
R226 B.n282 B.n281 585
R227 B.n283 B.n102 585
R228 B.n285 B.n284 585
R229 B.n286 B.n101 585
R230 B.n288 B.n287 585
R231 B.n289 B.n100 585
R232 B.n291 B.n290 585
R233 B.n292 B.n99 585
R234 B.n294 B.n293 585
R235 B.n295 B.n98 585
R236 B.n297 B.n296 585
R237 B.n298 B.n97 585
R238 B.n300 B.n299 585
R239 B.n301 B.n96 585
R240 B.n303 B.n302 585
R241 B.n304 B.n95 585
R242 B.n306 B.n305 585
R243 B.n307 B.n94 585
R244 B.n309 B.n308 585
R245 B.n310 B.n93 585
R246 B.n312 B.n311 585
R247 B.n313 B.n92 585
R248 B.n315 B.n314 585
R249 B.n316 B.n91 585
R250 B.n318 B.n317 585
R251 B.n319 B.n90 585
R252 B.n321 B.n320 585
R253 B.n322 B.n89 585
R254 B.n324 B.n323 585
R255 B.n325 B.n88 585
R256 B.n327 B.n326 585
R257 B.n328 B.n87 585
R258 B.n176 B.n175 585
R259 B.n174 B.n139 585
R260 B.n173 B.n172 585
R261 B.n171 B.n140 585
R262 B.n170 B.n169 585
R263 B.n168 B.n141 585
R264 B.n167 B.n166 585
R265 B.n165 B.n142 585
R266 B.n164 B.n163 585
R267 B.n162 B.n143 585
R268 B.n161 B.n160 585
R269 B.n159 B.n144 585
R270 B.n158 B.n157 585
R271 B.n156 B.n145 585
R272 B.n155 B.n154 585
R273 B.n153 B.n146 585
R274 B.n152 B.n151 585
R275 B.n150 B.n147 585
R276 B.n149 B.n148 585
R277 B.n2 B.n0 585
R278 B.n569 B.n1 585
R279 B.n568 B.n567 585
R280 B.n566 B.n3 585
R281 B.n565 B.n564 585
R282 B.n563 B.n4 585
R283 B.n562 B.n561 585
R284 B.n560 B.n5 585
R285 B.n559 B.n558 585
R286 B.n557 B.n6 585
R287 B.n556 B.n555 585
R288 B.n554 B.n7 585
R289 B.n553 B.n552 585
R290 B.n551 B.n8 585
R291 B.n550 B.n549 585
R292 B.n548 B.n9 585
R293 B.n547 B.n546 585
R294 B.n545 B.n10 585
R295 B.n544 B.n543 585
R296 B.n542 B.n11 585
R297 B.n541 B.n540 585
R298 B.n571 B.n570 585
R299 B.n175 B.n138 439.647
R300 B.n540 B.n539 439.647
R301 B.n329 B.n328 439.647
R302 B.n389 B.n66 439.647
R303 B.n257 B.t3 394.579
R304 B.n115 B.t9 394.579
R305 B.n36 B.t0 394.579
R306 B.n43 B.t6 394.579
R307 B.n175 B.n174 163.367
R308 B.n174 B.n173 163.367
R309 B.n173 B.n140 163.367
R310 B.n169 B.n140 163.367
R311 B.n169 B.n168 163.367
R312 B.n168 B.n167 163.367
R313 B.n167 B.n142 163.367
R314 B.n163 B.n142 163.367
R315 B.n163 B.n162 163.367
R316 B.n162 B.n161 163.367
R317 B.n161 B.n144 163.367
R318 B.n157 B.n144 163.367
R319 B.n157 B.n156 163.367
R320 B.n156 B.n155 163.367
R321 B.n155 B.n146 163.367
R322 B.n151 B.n146 163.367
R323 B.n151 B.n150 163.367
R324 B.n150 B.n149 163.367
R325 B.n149 B.n2 163.367
R326 B.n570 B.n2 163.367
R327 B.n570 B.n569 163.367
R328 B.n569 B.n568 163.367
R329 B.n568 B.n3 163.367
R330 B.n564 B.n3 163.367
R331 B.n564 B.n563 163.367
R332 B.n563 B.n562 163.367
R333 B.n562 B.n5 163.367
R334 B.n558 B.n5 163.367
R335 B.n558 B.n557 163.367
R336 B.n557 B.n556 163.367
R337 B.n556 B.n7 163.367
R338 B.n552 B.n7 163.367
R339 B.n552 B.n551 163.367
R340 B.n551 B.n550 163.367
R341 B.n550 B.n9 163.367
R342 B.n546 B.n9 163.367
R343 B.n546 B.n545 163.367
R344 B.n545 B.n544 163.367
R345 B.n544 B.n11 163.367
R346 B.n540 B.n11 163.367
R347 B.n179 B.n138 163.367
R348 B.n180 B.n179 163.367
R349 B.n181 B.n180 163.367
R350 B.n181 B.n136 163.367
R351 B.n185 B.n136 163.367
R352 B.n186 B.n185 163.367
R353 B.n187 B.n186 163.367
R354 B.n187 B.n134 163.367
R355 B.n191 B.n134 163.367
R356 B.n192 B.n191 163.367
R357 B.n193 B.n192 163.367
R358 B.n193 B.n132 163.367
R359 B.n197 B.n132 163.367
R360 B.n198 B.n197 163.367
R361 B.n199 B.n198 163.367
R362 B.n199 B.n130 163.367
R363 B.n203 B.n130 163.367
R364 B.n204 B.n203 163.367
R365 B.n205 B.n204 163.367
R366 B.n205 B.n128 163.367
R367 B.n209 B.n128 163.367
R368 B.n210 B.n209 163.367
R369 B.n211 B.n210 163.367
R370 B.n211 B.n126 163.367
R371 B.n215 B.n126 163.367
R372 B.n216 B.n215 163.367
R373 B.n217 B.n216 163.367
R374 B.n217 B.n124 163.367
R375 B.n221 B.n124 163.367
R376 B.n222 B.n221 163.367
R377 B.n223 B.n222 163.367
R378 B.n223 B.n122 163.367
R379 B.n227 B.n122 163.367
R380 B.n228 B.n227 163.367
R381 B.n229 B.n228 163.367
R382 B.n229 B.n120 163.367
R383 B.n233 B.n120 163.367
R384 B.n234 B.n233 163.367
R385 B.n235 B.n234 163.367
R386 B.n235 B.n118 163.367
R387 B.n239 B.n118 163.367
R388 B.n240 B.n239 163.367
R389 B.n241 B.n240 163.367
R390 B.n241 B.n114 163.367
R391 B.n246 B.n114 163.367
R392 B.n247 B.n246 163.367
R393 B.n248 B.n247 163.367
R394 B.n248 B.n112 163.367
R395 B.n252 B.n112 163.367
R396 B.n253 B.n252 163.367
R397 B.n254 B.n253 163.367
R398 B.n254 B.n110 163.367
R399 B.n261 B.n110 163.367
R400 B.n262 B.n261 163.367
R401 B.n263 B.n262 163.367
R402 B.n263 B.n108 163.367
R403 B.n267 B.n108 163.367
R404 B.n268 B.n267 163.367
R405 B.n269 B.n268 163.367
R406 B.n269 B.n106 163.367
R407 B.n273 B.n106 163.367
R408 B.n274 B.n273 163.367
R409 B.n275 B.n274 163.367
R410 B.n275 B.n104 163.367
R411 B.n279 B.n104 163.367
R412 B.n280 B.n279 163.367
R413 B.n281 B.n280 163.367
R414 B.n281 B.n102 163.367
R415 B.n285 B.n102 163.367
R416 B.n286 B.n285 163.367
R417 B.n287 B.n286 163.367
R418 B.n287 B.n100 163.367
R419 B.n291 B.n100 163.367
R420 B.n292 B.n291 163.367
R421 B.n293 B.n292 163.367
R422 B.n293 B.n98 163.367
R423 B.n297 B.n98 163.367
R424 B.n298 B.n297 163.367
R425 B.n299 B.n298 163.367
R426 B.n299 B.n96 163.367
R427 B.n303 B.n96 163.367
R428 B.n304 B.n303 163.367
R429 B.n305 B.n304 163.367
R430 B.n305 B.n94 163.367
R431 B.n309 B.n94 163.367
R432 B.n310 B.n309 163.367
R433 B.n311 B.n310 163.367
R434 B.n311 B.n92 163.367
R435 B.n315 B.n92 163.367
R436 B.n316 B.n315 163.367
R437 B.n317 B.n316 163.367
R438 B.n317 B.n90 163.367
R439 B.n321 B.n90 163.367
R440 B.n322 B.n321 163.367
R441 B.n323 B.n322 163.367
R442 B.n323 B.n88 163.367
R443 B.n327 B.n88 163.367
R444 B.n328 B.n327 163.367
R445 B.n329 B.n86 163.367
R446 B.n333 B.n86 163.367
R447 B.n334 B.n333 163.367
R448 B.n335 B.n334 163.367
R449 B.n335 B.n84 163.367
R450 B.n339 B.n84 163.367
R451 B.n340 B.n339 163.367
R452 B.n341 B.n340 163.367
R453 B.n341 B.n82 163.367
R454 B.n345 B.n82 163.367
R455 B.n346 B.n345 163.367
R456 B.n347 B.n346 163.367
R457 B.n347 B.n80 163.367
R458 B.n351 B.n80 163.367
R459 B.n352 B.n351 163.367
R460 B.n353 B.n352 163.367
R461 B.n353 B.n78 163.367
R462 B.n357 B.n78 163.367
R463 B.n358 B.n357 163.367
R464 B.n359 B.n358 163.367
R465 B.n359 B.n76 163.367
R466 B.n363 B.n76 163.367
R467 B.n364 B.n363 163.367
R468 B.n365 B.n364 163.367
R469 B.n365 B.n74 163.367
R470 B.n369 B.n74 163.367
R471 B.n370 B.n369 163.367
R472 B.n371 B.n370 163.367
R473 B.n371 B.n72 163.367
R474 B.n375 B.n72 163.367
R475 B.n376 B.n375 163.367
R476 B.n377 B.n376 163.367
R477 B.n377 B.n70 163.367
R478 B.n381 B.n70 163.367
R479 B.n382 B.n381 163.367
R480 B.n383 B.n382 163.367
R481 B.n383 B.n68 163.367
R482 B.n387 B.n68 163.367
R483 B.n388 B.n387 163.367
R484 B.n389 B.n388 163.367
R485 B.n539 B.n538 163.367
R486 B.n538 B.n13 163.367
R487 B.n534 B.n13 163.367
R488 B.n534 B.n533 163.367
R489 B.n533 B.n532 163.367
R490 B.n532 B.n15 163.367
R491 B.n528 B.n15 163.367
R492 B.n528 B.n527 163.367
R493 B.n527 B.n526 163.367
R494 B.n526 B.n17 163.367
R495 B.n522 B.n17 163.367
R496 B.n522 B.n521 163.367
R497 B.n521 B.n520 163.367
R498 B.n520 B.n19 163.367
R499 B.n516 B.n19 163.367
R500 B.n516 B.n515 163.367
R501 B.n515 B.n514 163.367
R502 B.n514 B.n21 163.367
R503 B.n510 B.n21 163.367
R504 B.n510 B.n509 163.367
R505 B.n509 B.n508 163.367
R506 B.n508 B.n23 163.367
R507 B.n504 B.n23 163.367
R508 B.n504 B.n503 163.367
R509 B.n503 B.n502 163.367
R510 B.n502 B.n25 163.367
R511 B.n498 B.n25 163.367
R512 B.n498 B.n497 163.367
R513 B.n497 B.n496 163.367
R514 B.n496 B.n27 163.367
R515 B.n492 B.n27 163.367
R516 B.n492 B.n491 163.367
R517 B.n491 B.n490 163.367
R518 B.n490 B.n29 163.367
R519 B.n486 B.n29 163.367
R520 B.n486 B.n485 163.367
R521 B.n485 B.n484 163.367
R522 B.n484 B.n31 163.367
R523 B.n480 B.n31 163.367
R524 B.n480 B.n479 163.367
R525 B.n479 B.n478 163.367
R526 B.n478 B.n33 163.367
R527 B.n474 B.n33 163.367
R528 B.n474 B.n473 163.367
R529 B.n473 B.n472 163.367
R530 B.n472 B.n35 163.367
R531 B.n468 B.n35 163.367
R532 B.n468 B.n467 163.367
R533 B.n467 B.n466 163.367
R534 B.n466 B.n40 163.367
R535 B.n462 B.n40 163.367
R536 B.n462 B.n461 163.367
R537 B.n461 B.n460 163.367
R538 B.n460 B.n42 163.367
R539 B.n455 B.n42 163.367
R540 B.n455 B.n454 163.367
R541 B.n454 B.n453 163.367
R542 B.n453 B.n46 163.367
R543 B.n449 B.n46 163.367
R544 B.n449 B.n448 163.367
R545 B.n448 B.n447 163.367
R546 B.n447 B.n48 163.367
R547 B.n443 B.n48 163.367
R548 B.n443 B.n442 163.367
R549 B.n442 B.n441 163.367
R550 B.n441 B.n50 163.367
R551 B.n437 B.n50 163.367
R552 B.n437 B.n436 163.367
R553 B.n436 B.n435 163.367
R554 B.n435 B.n52 163.367
R555 B.n431 B.n52 163.367
R556 B.n431 B.n430 163.367
R557 B.n430 B.n429 163.367
R558 B.n429 B.n54 163.367
R559 B.n425 B.n54 163.367
R560 B.n425 B.n424 163.367
R561 B.n424 B.n423 163.367
R562 B.n423 B.n56 163.367
R563 B.n419 B.n56 163.367
R564 B.n419 B.n418 163.367
R565 B.n418 B.n417 163.367
R566 B.n417 B.n58 163.367
R567 B.n413 B.n58 163.367
R568 B.n413 B.n412 163.367
R569 B.n412 B.n411 163.367
R570 B.n411 B.n60 163.367
R571 B.n407 B.n60 163.367
R572 B.n407 B.n406 163.367
R573 B.n406 B.n405 163.367
R574 B.n405 B.n62 163.367
R575 B.n401 B.n62 163.367
R576 B.n401 B.n400 163.367
R577 B.n400 B.n399 163.367
R578 B.n399 B.n64 163.367
R579 B.n395 B.n64 163.367
R580 B.n395 B.n394 163.367
R581 B.n394 B.n393 163.367
R582 B.n393 B.n66 163.367
R583 B.n257 B.t5 146.847
R584 B.n43 B.t7 146.847
R585 B.n115 B.t11 146.832
R586 B.n36 B.t1 146.832
R587 B.n258 B.t4 108.254
R588 B.n44 B.t8 108.254
R589 B.n116 B.t10 108.237
R590 B.n37 B.t2 108.237
R591 B.n259 B.n258 59.5399
R592 B.n244 B.n116 59.5399
R593 B.n38 B.n37 59.5399
R594 B.n458 B.n44 59.5399
R595 B.n258 B.n257 38.5944
R596 B.n116 B.n115 38.5944
R597 B.n37 B.n36 38.5944
R598 B.n44 B.n43 38.5944
R599 B.n541 B.n12 28.5664
R600 B.n330 B.n87 28.5664
R601 B.n177 B.n176 28.5664
R602 B.n391 B.n390 28.5664
R603 B B.n571 18.0485
R604 B.n537 B.n12 10.6151
R605 B.n537 B.n536 10.6151
R606 B.n536 B.n535 10.6151
R607 B.n535 B.n14 10.6151
R608 B.n531 B.n14 10.6151
R609 B.n531 B.n530 10.6151
R610 B.n530 B.n529 10.6151
R611 B.n529 B.n16 10.6151
R612 B.n525 B.n16 10.6151
R613 B.n525 B.n524 10.6151
R614 B.n524 B.n523 10.6151
R615 B.n523 B.n18 10.6151
R616 B.n519 B.n18 10.6151
R617 B.n519 B.n518 10.6151
R618 B.n518 B.n517 10.6151
R619 B.n517 B.n20 10.6151
R620 B.n513 B.n20 10.6151
R621 B.n513 B.n512 10.6151
R622 B.n512 B.n511 10.6151
R623 B.n511 B.n22 10.6151
R624 B.n507 B.n22 10.6151
R625 B.n507 B.n506 10.6151
R626 B.n506 B.n505 10.6151
R627 B.n505 B.n24 10.6151
R628 B.n501 B.n24 10.6151
R629 B.n501 B.n500 10.6151
R630 B.n500 B.n499 10.6151
R631 B.n499 B.n26 10.6151
R632 B.n495 B.n26 10.6151
R633 B.n495 B.n494 10.6151
R634 B.n494 B.n493 10.6151
R635 B.n493 B.n28 10.6151
R636 B.n489 B.n28 10.6151
R637 B.n489 B.n488 10.6151
R638 B.n488 B.n487 10.6151
R639 B.n487 B.n30 10.6151
R640 B.n483 B.n30 10.6151
R641 B.n483 B.n482 10.6151
R642 B.n482 B.n481 10.6151
R643 B.n481 B.n32 10.6151
R644 B.n477 B.n32 10.6151
R645 B.n477 B.n476 10.6151
R646 B.n476 B.n475 10.6151
R647 B.n475 B.n34 10.6151
R648 B.n471 B.n470 10.6151
R649 B.n470 B.n469 10.6151
R650 B.n469 B.n39 10.6151
R651 B.n465 B.n39 10.6151
R652 B.n465 B.n464 10.6151
R653 B.n464 B.n463 10.6151
R654 B.n463 B.n41 10.6151
R655 B.n459 B.n41 10.6151
R656 B.n457 B.n456 10.6151
R657 B.n456 B.n45 10.6151
R658 B.n452 B.n45 10.6151
R659 B.n452 B.n451 10.6151
R660 B.n451 B.n450 10.6151
R661 B.n450 B.n47 10.6151
R662 B.n446 B.n47 10.6151
R663 B.n446 B.n445 10.6151
R664 B.n445 B.n444 10.6151
R665 B.n444 B.n49 10.6151
R666 B.n440 B.n49 10.6151
R667 B.n440 B.n439 10.6151
R668 B.n439 B.n438 10.6151
R669 B.n438 B.n51 10.6151
R670 B.n434 B.n51 10.6151
R671 B.n434 B.n433 10.6151
R672 B.n433 B.n432 10.6151
R673 B.n432 B.n53 10.6151
R674 B.n428 B.n53 10.6151
R675 B.n428 B.n427 10.6151
R676 B.n427 B.n426 10.6151
R677 B.n426 B.n55 10.6151
R678 B.n422 B.n55 10.6151
R679 B.n422 B.n421 10.6151
R680 B.n421 B.n420 10.6151
R681 B.n420 B.n57 10.6151
R682 B.n416 B.n57 10.6151
R683 B.n416 B.n415 10.6151
R684 B.n415 B.n414 10.6151
R685 B.n414 B.n59 10.6151
R686 B.n410 B.n59 10.6151
R687 B.n410 B.n409 10.6151
R688 B.n409 B.n408 10.6151
R689 B.n408 B.n61 10.6151
R690 B.n404 B.n61 10.6151
R691 B.n404 B.n403 10.6151
R692 B.n403 B.n402 10.6151
R693 B.n402 B.n63 10.6151
R694 B.n398 B.n63 10.6151
R695 B.n398 B.n397 10.6151
R696 B.n397 B.n396 10.6151
R697 B.n396 B.n65 10.6151
R698 B.n392 B.n65 10.6151
R699 B.n392 B.n391 10.6151
R700 B.n331 B.n330 10.6151
R701 B.n332 B.n331 10.6151
R702 B.n332 B.n85 10.6151
R703 B.n336 B.n85 10.6151
R704 B.n337 B.n336 10.6151
R705 B.n338 B.n337 10.6151
R706 B.n338 B.n83 10.6151
R707 B.n342 B.n83 10.6151
R708 B.n343 B.n342 10.6151
R709 B.n344 B.n343 10.6151
R710 B.n344 B.n81 10.6151
R711 B.n348 B.n81 10.6151
R712 B.n349 B.n348 10.6151
R713 B.n350 B.n349 10.6151
R714 B.n350 B.n79 10.6151
R715 B.n354 B.n79 10.6151
R716 B.n355 B.n354 10.6151
R717 B.n356 B.n355 10.6151
R718 B.n356 B.n77 10.6151
R719 B.n360 B.n77 10.6151
R720 B.n361 B.n360 10.6151
R721 B.n362 B.n361 10.6151
R722 B.n362 B.n75 10.6151
R723 B.n366 B.n75 10.6151
R724 B.n367 B.n366 10.6151
R725 B.n368 B.n367 10.6151
R726 B.n368 B.n73 10.6151
R727 B.n372 B.n73 10.6151
R728 B.n373 B.n372 10.6151
R729 B.n374 B.n373 10.6151
R730 B.n374 B.n71 10.6151
R731 B.n378 B.n71 10.6151
R732 B.n379 B.n378 10.6151
R733 B.n380 B.n379 10.6151
R734 B.n380 B.n69 10.6151
R735 B.n384 B.n69 10.6151
R736 B.n385 B.n384 10.6151
R737 B.n386 B.n385 10.6151
R738 B.n386 B.n67 10.6151
R739 B.n390 B.n67 10.6151
R740 B.n178 B.n177 10.6151
R741 B.n178 B.n137 10.6151
R742 B.n182 B.n137 10.6151
R743 B.n183 B.n182 10.6151
R744 B.n184 B.n183 10.6151
R745 B.n184 B.n135 10.6151
R746 B.n188 B.n135 10.6151
R747 B.n189 B.n188 10.6151
R748 B.n190 B.n189 10.6151
R749 B.n190 B.n133 10.6151
R750 B.n194 B.n133 10.6151
R751 B.n195 B.n194 10.6151
R752 B.n196 B.n195 10.6151
R753 B.n196 B.n131 10.6151
R754 B.n200 B.n131 10.6151
R755 B.n201 B.n200 10.6151
R756 B.n202 B.n201 10.6151
R757 B.n202 B.n129 10.6151
R758 B.n206 B.n129 10.6151
R759 B.n207 B.n206 10.6151
R760 B.n208 B.n207 10.6151
R761 B.n208 B.n127 10.6151
R762 B.n212 B.n127 10.6151
R763 B.n213 B.n212 10.6151
R764 B.n214 B.n213 10.6151
R765 B.n214 B.n125 10.6151
R766 B.n218 B.n125 10.6151
R767 B.n219 B.n218 10.6151
R768 B.n220 B.n219 10.6151
R769 B.n220 B.n123 10.6151
R770 B.n224 B.n123 10.6151
R771 B.n225 B.n224 10.6151
R772 B.n226 B.n225 10.6151
R773 B.n226 B.n121 10.6151
R774 B.n230 B.n121 10.6151
R775 B.n231 B.n230 10.6151
R776 B.n232 B.n231 10.6151
R777 B.n232 B.n119 10.6151
R778 B.n236 B.n119 10.6151
R779 B.n237 B.n236 10.6151
R780 B.n238 B.n237 10.6151
R781 B.n238 B.n117 10.6151
R782 B.n242 B.n117 10.6151
R783 B.n243 B.n242 10.6151
R784 B.n245 B.n113 10.6151
R785 B.n249 B.n113 10.6151
R786 B.n250 B.n249 10.6151
R787 B.n251 B.n250 10.6151
R788 B.n251 B.n111 10.6151
R789 B.n255 B.n111 10.6151
R790 B.n256 B.n255 10.6151
R791 B.n260 B.n256 10.6151
R792 B.n264 B.n109 10.6151
R793 B.n265 B.n264 10.6151
R794 B.n266 B.n265 10.6151
R795 B.n266 B.n107 10.6151
R796 B.n270 B.n107 10.6151
R797 B.n271 B.n270 10.6151
R798 B.n272 B.n271 10.6151
R799 B.n272 B.n105 10.6151
R800 B.n276 B.n105 10.6151
R801 B.n277 B.n276 10.6151
R802 B.n278 B.n277 10.6151
R803 B.n278 B.n103 10.6151
R804 B.n282 B.n103 10.6151
R805 B.n283 B.n282 10.6151
R806 B.n284 B.n283 10.6151
R807 B.n284 B.n101 10.6151
R808 B.n288 B.n101 10.6151
R809 B.n289 B.n288 10.6151
R810 B.n290 B.n289 10.6151
R811 B.n290 B.n99 10.6151
R812 B.n294 B.n99 10.6151
R813 B.n295 B.n294 10.6151
R814 B.n296 B.n295 10.6151
R815 B.n296 B.n97 10.6151
R816 B.n300 B.n97 10.6151
R817 B.n301 B.n300 10.6151
R818 B.n302 B.n301 10.6151
R819 B.n302 B.n95 10.6151
R820 B.n306 B.n95 10.6151
R821 B.n307 B.n306 10.6151
R822 B.n308 B.n307 10.6151
R823 B.n308 B.n93 10.6151
R824 B.n312 B.n93 10.6151
R825 B.n313 B.n312 10.6151
R826 B.n314 B.n313 10.6151
R827 B.n314 B.n91 10.6151
R828 B.n318 B.n91 10.6151
R829 B.n319 B.n318 10.6151
R830 B.n320 B.n319 10.6151
R831 B.n320 B.n89 10.6151
R832 B.n324 B.n89 10.6151
R833 B.n325 B.n324 10.6151
R834 B.n326 B.n325 10.6151
R835 B.n326 B.n87 10.6151
R836 B.n176 B.n139 10.6151
R837 B.n172 B.n139 10.6151
R838 B.n172 B.n171 10.6151
R839 B.n171 B.n170 10.6151
R840 B.n170 B.n141 10.6151
R841 B.n166 B.n141 10.6151
R842 B.n166 B.n165 10.6151
R843 B.n165 B.n164 10.6151
R844 B.n164 B.n143 10.6151
R845 B.n160 B.n143 10.6151
R846 B.n160 B.n159 10.6151
R847 B.n159 B.n158 10.6151
R848 B.n158 B.n145 10.6151
R849 B.n154 B.n145 10.6151
R850 B.n154 B.n153 10.6151
R851 B.n153 B.n152 10.6151
R852 B.n152 B.n147 10.6151
R853 B.n148 B.n147 10.6151
R854 B.n148 B.n0 10.6151
R855 B.n567 B.n1 10.6151
R856 B.n567 B.n566 10.6151
R857 B.n566 B.n565 10.6151
R858 B.n565 B.n4 10.6151
R859 B.n561 B.n4 10.6151
R860 B.n561 B.n560 10.6151
R861 B.n560 B.n559 10.6151
R862 B.n559 B.n6 10.6151
R863 B.n555 B.n6 10.6151
R864 B.n555 B.n554 10.6151
R865 B.n554 B.n553 10.6151
R866 B.n553 B.n8 10.6151
R867 B.n549 B.n8 10.6151
R868 B.n549 B.n548 10.6151
R869 B.n548 B.n547 10.6151
R870 B.n547 B.n10 10.6151
R871 B.n543 B.n10 10.6151
R872 B.n543 B.n542 10.6151
R873 B.n542 B.n541 10.6151
R874 B.n471 B.n38 6.5566
R875 B.n459 B.n458 6.5566
R876 B.n245 B.n244 6.5566
R877 B.n260 B.n259 6.5566
R878 B.n38 B.n34 4.05904
R879 B.n458 B.n457 4.05904
R880 B.n244 B.n243 4.05904
R881 B.n259 B.n109 4.05904
R882 B.n571 B.n0 2.81026
R883 B.n571 B.n1 2.81026
C0 VN w_n1766_n3566# 2.38439f
C1 VN B 0.902659f
C2 B w_n1766_n3566# 8.07058f
C3 VN VDD2 2.74819f
C4 VDD2 w_n1766_n3566# 1.76122f
C5 VDD2 B 1.67055f
C6 VDD1 VTAIL 5.3243f
C7 VDD1 VP 2.89087f
C8 VP VTAIL 2.32208f
C9 VN VDD1 0.147691f
C10 VDD1 w_n1766_n3566# 1.74661f
C11 VDD1 B 1.64877f
C12 VN VTAIL 2.30766f
C13 VN VP 5.20106f
C14 VTAIL w_n1766_n3566# 2.93284f
C15 VTAIL B 3.4417f
C16 VP w_n1766_n3566# 2.60732f
C17 VP B 1.26539f
C18 VDD1 VDD2 0.564383f
C19 VDD2 VTAIL 5.36692f
C20 VDD2 VP 0.293785f
C21 VDD2 VSUBS 0.846586f
C22 VDD1 VSUBS 4.304294f
C23 VTAIL VSUBS 0.935259f
C24 VN VSUBS 7.93584f
C25 VP VSUBS 1.450027f
C26 B VSUBS 3.281236f
C27 w_n1766_n3566# VSUBS 77.4144f
C28 B.n0 VSUBS 0.004089f
C29 B.n1 VSUBS 0.004089f
C30 B.n2 VSUBS 0.006466f
C31 B.n3 VSUBS 0.006466f
C32 B.n4 VSUBS 0.006466f
C33 B.n5 VSUBS 0.006466f
C34 B.n6 VSUBS 0.006466f
C35 B.n7 VSUBS 0.006466f
C36 B.n8 VSUBS 0.006466f
C37 B.n9 VSUBS 0.006466f
C38 B.n10 VSUBS 0.006466f
C39 B.n11 VSUBS 0.006466f
C40 B.n12 VSUBS 0.014299f
C41 B.n13 VSUBS 0.006466f
C42 B.n14 VSUBS 0.006466f
C43 B.n15 VSUBS 0.006466f
C44 B.n16 VSUBS 0.006466f
C45 B.n17 VSUBS 0.006466f
C46 B.n18 VSUBS 0.006466f
C47 B.n19 VSUBS 0.006466f
C48 B.n20 VSUBS 0.006466f
C49 B.n21 VSUBS 0.006466f
C50 B.n22 VSUBS 0.006466f
C51 B.n23 VSUBS 0.006466f
C52 B.n24 VSUBS 0.006466f
C53 B.n25 VSUBS 0.006466f
C54 B.n26 VSUBS 0.006466f
C55 B.n27 VSUBS 0.006466f
C56 B.n28 VSUBS 0.006466f
C57 B.n29 VSUBS 0.006466f
C58 B.n30 VSUBS 0.006466f
C59 B.n31 VSUBS 0.006466f
C60 B.n32 VSUBS 0.006466f
C61 B.n33 VSUBS 0.006466f
C62 B.n34 VSUBS 0.004469f
C63 B.n35 VSUBS 0.006466f
C64 B.t2 VSUBS 0.39424f
C65 B.t1 VSUBS 0.408322f
C66 B.t0 VSUBS 0.87332f
C67 B.n36 VSUBS 0.186716f
C68 B.n37 VSUBS 0.062799f
C69 B.n38 VSUBS 0.014982f
C70 B.n39 VSUBS 0.006466f
C71 B.n40 VSUBS 0.006466f
C72 B.n41 VSUBS 0.006466f
C73 B.n42 VSUBS 0.006466f
C74 B.t8 VSUBS 0.394231f
C75 B.t7 VSUBS 0.408314f
C76 B.t6 VSUBS 0.87332f
C77 B.n43 VSUBS 0.186724f
C78 B.n44 VSUBS 0.062808f
C79 B.n45 VSUBS 0.006466f
C80 B.n46 VSUBS 0.006466f
C81 B.n47 VSUBS 0.006466f
C82 B.n48 VSUBS 0.006466f
C83 B.n49 VSUBS 0.006466f
C84 B.n50 VSUBS 0.006466f
C85 B.n51 VSUBS 0.006466f
C86 B.n52 VSUBS 0.006466f
C87 B.n53 VSUBS 0.006466f
C88 B.n54 VSUBS 0.006466f
C89 B.n55 VSUBS 0.006466f
C90 B.n56 VSUBS 0.006466f
C91 B.n57 VSUBS 0.006466f
C92 B.n58 VSUBS 0.006466f
C93 B.n59 VSUBS 0.006466f
C94 B.n60 VSUBS 0.006466f
C95 B.n61 VSUBS 0.006466f
C96 B.n62 VSUBS 0.006466f
C97 B.n63 VSUBS 0.006466f
C98 B.n64 VSUBS 0.006466f
C99 B.n65 VSUBS 0.006466f
C100 B.n66 VSUBS 0.014299f
C101 B.n67 VSUBS 0.006466f
C102 B.n68 VSUBS 0.006466f
C103 B.n69 VSUBS 0.006466f
C104 B.n70 VSUBS 0.006466f
C105 B.n71 VSUBS 0.006466f
C106 B.n72 VSUBS 0.006466f
C107 B.n73 VSUBS 0.006466f
C108 B.n74 VSUBS 0.006466f
C109 B.n75 VSUBS 0.006466f
C110 B.n76 VSUBS 0.006466f
C111 B.n77 VSUBS 0.006466f
C112 B.n78 VSUBS 0.006466f
C113 B.n79 VSUBS 0.006466f
C114 B.n80 VSUBS 0.006466f
C115 B.n81 VSUBS 0.006466f
C116 B.n82 VSUBS 0.006466f
C117 B.n83 VSUBS 0.006466f
C118 B.n84 VSUBS 0.006466f
C119 B.n85 VSUBS 0.006466f
C120 B.n86 VSUBS 0.006466f
C121 B.n87 VSUBS 0.014299f
C122 B.n88 VSUBS 0.006466f
C123 B.n89 VSUBS 0.006466f
C124 B.n90 VSUBS 0.006466f
C125 B.n91 VSUBS 0.006466f
C126 B.n92 VSUBS 0.006466f
C127 B.n93 VSUBS 0.006466f
C128 B.n94 VSUBS 0.006466f
C129 B.n95 VSUBS 0.006466f
C130 B.n96 VSUBS 0.006466f
C131 B.n97 VSUBS 0.006466f
C132 B.n98 VSUBS 0.006466f
C133 B.n99 VSUBS 0.006466f
C134 B.n100 VSUBS 0.006466f
C135 B.n101 VSUBS 0.006466f
C136 B.n102 VSUBS 0.006466f
C137 B.n103 VSUBS 0.006466f
C138 B.n104 VSUBS 0.006466f
C139 B.n105 VSUBS 0.006466f
C140 B.n106 VSUBS 0.006466f
C141 B.n107 VSUBS 0.006466f
C142 B.n108 VSUBS 0.006466f
C143 B.n109 VSUBS 0.004469f
C144 B.n110 VSUBS 0.006466f
C145 B.n111 VSUBS 0.006466f
C146 B.n112 VSUBS 0.006466f
C147 B.n113 VSUBS 0.006466f
C148 B.n114 VSUBS 0.006466f
C149 B.t10 VSUBS 0.39424f
C150 B.t11 VSUBS 0.408322f
C151 B.t9 VSUBS 0.87332f
C152 B.n115 VSUBS 0.186716f
C153 B.n116 VSUBS 0.062799f
C154 B.n117 VSUBS 0.006466f
C155 B.n118 VSUBS 0.006466f
C156 B.n119 VSUBS 0.006466f
C157 B.n120 VSUBS 0.006466f
C158 B.n121 VSUBS 0.006466f
C159 B.n122 VSUBS 0.006466f
C160 B.n123 VSUBS 0.006466f
C161 B.n124 VSUBS 0.006466f
C162 B.n125 VSUBS 0.006466f
C163 B.n126 VSUBS 0.006466f
C164 B.n127 VSUBS 0.006466f
C165 B.n128 VSUBS 0.006466f
C166 B.n129 VSUBS 0.006466f
C167 B.n130 VSUBS 0.006466f
C168 B.n131 VSUBS 0.006466f
C169 B.n132 VSUBS 0.006466f
C170 B.n133 VSUBS 0.006466f
C171 B.n134 VSUBS 0.006466f
C172 B.n135 VSUBS 0.006466f
C173 B.n136 VSUBS 0.006466f
C174 B.n137 VSUBS 0.006466f
C175 B.n138 VSUBS 0.014299f
C176 B.n139 VSUBS 0.006466f
C177 B.n140 VSUBS 0.006466f
C178 B.n141 VSUBS 0.006466f
C179 B.n142 VSUBS 0.006466f
C180 B.n143 VSUBS 0.006466f
C181 B.n144 VSUBS 0.006466f
C182 B.n145 VSUBS 0.006466f
C183 B.n146 VSUBS 0.006466f
C184 B.n147 VSUBS 0.006466f
C185 B.n148 VSUBS 0.006466f
C186 B.n149 VSUBS 0.006466f
C187 B.n150 VSUBS 0.006466f
C188 B.n151 VSUBS 0.006466f
C189 B.n152 VSUBS 0.006466f
C190 B.n153 VSUBS 0.006466f
C191 B.n154 VSUBS 0.006466f
C192 B.n155 VSUBS 0.006466f
C193 B.n156 VSUBS 0.006466f
C194 B.n157 VSUBS 0.006466f
C195 B.n158 VSUBS 0.006466f
C196 B.n159 VSUBS 0.006466f
C197 B.n160 VSUBS 0.006466f
C198 B.n161 VSUBS 0.006466f
C199 B.n162 VSUBS 0.006466f
C200 B.n163 VSUBS 0.006466f
C201 B.n164 VSUBS 0.006466f
C202 B.n165 VSUBS 0.006466f
C203 B.n166 VSUBS 0.006466f
C204 B.n167 VSUBS 0.006466f
C205 B.n168 VSUBS 0.006466f
C206 B.n169 VSUBS 0.006466f
C207 B.n170 VSUBS 0.006466f
C208 B.n171 VSUBS 0.006466f
C209 B.n172 VSUBS 0.006466f
C210 B.n173 VSUBS 0.006466f
C211 B.n174 VSUBS 0.006466f
C212 B.n175 VSUBS 0.013468f
C213 B.n176 VSUBS 0.013468f
C214 B.n177 VSUBS 0.014299f
C215 B.n178 VSUBS 0.006466f
C216 B.n179 VSUBS 0.006466f
C217 B.n180 VSUBS 0.006466f
C218 B.n181 VSUBS 0.006466f
C219 B.n182 VSUBS 0.006466f
C220 B.n183 VSUBS 0.006466f
C221 B.n184 VSUBS 0.006466f
C222 B.n185 VSUBS 0.006466f
C223 B.n186 VSUBS 0.006466f
C224 B.n187 VSUBS 0.006466f
C225 B.n188 VSUBS 0.006466f
C226 B.n189 VSUBS 0.006466f
C227 B.n190 VSUBS 0.006466f
C228 B.n191 VSUBS 0.006466f
C229 B.n192 VSUBS 0.006466f
C230 B.n193 VSUBS 0.006466f
C231 B.n194 VSUBS 0.006466f
C232 B.n195 VSUBS 0.006466f
C233 B.n196 VSUBS 0.006466f
C234 B.n197 VSUBS 0.006466f
C235 B.n198 VSUBS 0.006466f
C236 B.n199 VSUBS 0.006466f
C237 B.n200 VSUBS 0.006466f
C238 B.n201 VSUBS 0.006466f
C239 B.n202 VSUBS 0.006466f
C240 B.n203 VSUBS 0.006466f
C241 B.n204 VSUBS 0.006466f
C242 B.n205 VSUBS 0.006466f
C243 B.n206 VSUBS 0.006466f
C244 B.n207 VSUBS 0.006466f
C245 B.n208 VSUBS 0.006466f
C246 B.n209 VSUBS 0.006466f
C247 B.n210 VSUBS 0.006466f
C248 B.n211 VSUBS 0.006466f
C249 B.n212 VSUBS 0.006466f
C250 B.n213 VSUBS 0.006466f
C251 B.n214 VSUBS 0.006466f
C252 B.n215 VSUBS 0.006466f
C253 B.n216 VSUBS 0.006466f
C254 B.n217 VSUBS 0.006466f
C255 B.n218 VSUBS 0.006466f
C256 B.n219 VSUBS 0.006466f
C257 B.n220 VSUBS 0.006466f
C258 B.n221 VSUBS 0.006466f
C259 B.n222 VSUBS 0.006466f
C260 B.n223 VSUBS 0.006466f
C261 B.n224 VSUBS 0.006466f
C262 B.n225 VSUBS 0.006466f
C263 B.n226 VSUBS 0.006466f
C264 B.n227 VSUBS 0.006466f
C265 B.n228 VSUBS 0.006466f
C266 B.n229 VSUBS 0.006466f
C267 B.n230 VSUBS 0.006466f
C268 B.n231 VSUBS 0.006466f
C269 B.n232 VSUBS 0.006466f
C270 B.n233 VSUBS 0.006466f
C271 B.n234 VSUBS 0.006466f
C272 B.n235 VSUBS 0.006466f
C273 B.n236 VSUBS 0.006466f
C274 B.n237 VSUBS 0.006466f
C275 B.n238 VSUBS 0.006466f
C276 B.n239 VSUBS 0.006466f
C277 B.n240 VSUBS 0.006466f
C278 B.n241 VSUBS 0.006466f
C279 B.n242 VSUBS 0.006466f
C280 B.n243 VSUBS 0.004469f
C281 B.n244 VSUBS 0.014982f
C282 B.n245 VSUBS 0.00523f
C283 B.n246 VSUBS 0.006466f
C284 B.n247 VSUBS 0.006466f
C285 B.n248 VSUBS 0.006466f
C286 B.n249 VSUBS 0.006466f
C287 B.n250 VSUBS 0.006466f
C288 B.n251 VSUBS 0.006466f
C289 B.n252 VSUBS 0.006466f
C290 B.n253 VSUBS 0.006466f
C291 B.n254 VSUBS 0.006466f
C292 B.n255 VSUBS 0.006466f
C293 B.n256 VSUBS 0.006466f
C294 B.t4 VSUBS 0.394231f
C295 B.t5 VSUBS 0.408314f
C296 B.t3 VSUBS 0.87332f
C297 B.n257 VSUBS 0.186724f
C298 B.n258 VSUBS 0.062808f
C299 B.n259 VSUBS 0.014982f
C300 B.n260 VSUBS 0.00523f
C301 B.n261 VSUBS 0.006466f
C302 B.n262 VSUBS 0.006466f
C303 B.n263 VSUBS 0.006466f
C304 B.n264 VSUBS 0.006466f
C305 B.n265 VSUBS 0.006466f
C306 B.n266 VSUBS 0.006466f
C307 B.n267 VSUBS 0.006466f
C308 B.n268 VSUBS 0.006466f
C309 B.n269 VSUBS 0.006466f
C310 B.n270 VSUBS 0.006466f
C311 B.n271 VSUBS 0.006466f
C312 B.n272 VSUBS 0.006466f
C313 B.n273 VSUBS 0.006466f
C314 B.n274 VSUBS 0.006466f
C315 B.n275 VSUBS 0.006466f
C316 B.n276 VSUBS 0.006466f
C317 B.n277 VSUBS 0.006466f
C318 B.n278 VSUBS 0.006466f
C319 B.n279 VSUBS 0.006466f
C320 B.n280 VSUBS 0.006466f
C321 B.n281 VSUBS 0.006466f
C322 B.n282 VSUBS 0.006466f
C323 B.n283 VSUBS 0.006466f
C324 B.n284 VSUBS 0.006466f
C325 B.n285 VSUBS 0.006466f
C326 B.n286 VSUBS 0.006466f
C327 B.n287 VSUBS 0.006466f
C328 B.n288 VSUBS 0.006466f
C329 B.n289 VSUBS 0.006466f
C330 B.n290 VSUBS 0.006466f
C331 B.n291 VSUBS 0.006466f
C332 B.n292 VSUBS 0.006466f
C333 B.n293 VSUBS 0.006466f
C334 B.n294 VSUBS 0.006466f
C335 B.n295 VSUBS 0.006466f
C336 B.n296 VSUBS 0.006466f
C337 B.n297 VSUBS 0.006466f
C338 B.n298 VSUBS 0.006466f
C339 B.n299 VSUBS 0.006466f
C340 B.n300 VSUBS 0.006466f
C341 B.n301 VSUBS 0.006466f
C342 B.n302 VSUBS 0.006466f
C343 B.n303 VSUBS 0.006466f
C344 B.n304 VSUBS 0.006466f
C345 B.n305 VSUBS 0.006466f
C346 B.n306 VSUBS 0.006466f
C347 B.n307 VSUBS 0.006466f
C348 B.n308 VSUBS 0.006466f
C349 B.n309 VSUBS 0.006466f
C350 B.n310 VSUBS 0.006466f
C351 B.n311 VSUBS 0.006466f
C352 B.n312 VSUBS 0.006466f
C353 B.n313 VSUBS 0.006466f
C354 B.n314 VSUBS 0.006466f
C355 B.n315 VSUBS 0.006466f
C356 B.n316 VSUBS 0.006466f
C357 B.n317 VSUBS 0.006466f
C358 B.n318 VSUBS 0.006466f
C359 B.n319 VSUBS 0.006466f
C360 B.n320 VSUBS 0.006466f
C361 B.n321 VSUBS 0.006466f
C362 B.n322 VSUBS 0.006466f
C363 B.n323 VSUBS 0.006466f
C364 B.n324 VSUBS 0.006466f
C365 B.n325 VSUBS 0.006466f
C366 B.n326 VSUBS 0.006466f
C367 B.n327 VSUBS 0.006466f
C368 B.n328 VSUBS 0.014299f
C369 B.n329 VSUBS 0.013468f
C370 B.n330 VSUBS 0.013468f
C371 B.n331 VSUBS 0.006466f
C372 B.n332 VSUBS 0.006466f
C373 B.n333 VSUBS 0.006466f
C374 B.n334 VSUBS 0.006466f
C375 B.n335 VSUBS 0.006466f
C376 B.n336 VSUBS 0.006466f
C377 B.n337 VSUBS 0.006466f
C378 B.n338 VSUBS 0.006466f
C379 B.n339 VSUBS 0.006466f
C380 B.n340 VSUBS 0.006466f
C381 B.n341 VSUBS 0.006466f
C382 B.n342 VSUBS 0.006466f
C383 B.n343 VSUBS 0.006466f
C384 B.n344 VSUBS 0.006466f
C385 B.n345 VSUBS 0.006466f
C386 B.n346 VSUBS 0.006466f
C387 B.n347 VSUBS 0.006466f
C388 B.n348 VSUBS 0.006466f
C389 B.n349 VSUBS 0.006466f
C390 B.n350 VSUBS 0.006466f
C391 B.n351 VSUBS 0.006466f
C392 B.n352 VSUBS 0.006466f
C393 B.n353 VSUBS 0.006466f
C394 B.n354 VSUBS 0.006466f
C395 B.n355 VSUBS 0.006466f
C396 B.n356 VSUBS 0.006466f
C397 B.n357 VSUBS 0.006466f
C398 B.n358 VSUBS 0.006466f
C399 B.n359 VSUBS 0.006466f
C400 B.n360 VSUBS 0.006466f
C401 B.n361 VSUBS 0.006466f
C402 B.n362 VSUBS 0.006466f
C403 B.n363 VSUBS 0.006466f
C404 B.n364 VSUBS 0.006466f
C405 B.n365 VSUBS 0.006466f
C406 B.n366 VSUBS 0.006466f
C407 B.n367 VSUBS 0.006466f
C408 B.n368 VSUBS 0.006466f
C409 B.n369 VSUBS 0.006466f
C410 B.n370 VSUBS 0.006466f
C411 B.n371 VSUBS 0.006466f
C412 B.n372 VSUBS 0.006466f
C413 B.n373 VSUBS 0.006466f
C414 B.n374 VSUBS 0.006466f
C415 B.n375 VSUBS 0.006466f
C416 B.n376 VSUBS 0.006466f
C417 B.n377 VSUBS 0.006466f
C418 B.n378 VSUBS 0.006466f
C419 B.n379 VSUBS 0.006466f
C420 B.n380 VSUBS 0.006466f
C421 B.n381 VSUBS 0.006466f
C422 B.n382 VSUBS 0.006466f
C423 B.n383 VSUBS 0.006466f
C424 B.n384 VSUBS 0.006466f
C425 B.n385 VSUBS 0.006466f
C426 B.n386 VSUBS 0.006466f
C427 B.n387 VSUBS 0.006466f
C428 B.n388 VSUBS 0.006466f
C429 B.n389 VSUBS 0.013468f
C430 B.n390 VSUBS 0.014342f
C431 B.n391 VSUBS 0.013425f
C432 B.n392 VSUBS 0.006466f
C433 B.n393 VSUBS 0.006466f
C434 B.n394 VSUBS 0.006466f
C435 B.n395 VSUBS 0.006466f
C436 B.n396 VSUBS 0.006466f
C437 B.n397 VSUBS 0.006466f
C438 B.n398 VSUBS 0.006466f
C439 B.n399 VSUBS 0.006466f
C440 B.n400 VSUBS 0.006466f
C441 B.n401 VSUBS 0.006466f
C442 B.n402 VSUBS 0.006466f
C443 B.n403 VSUBS 0.006466f
C444 B.n404 VSUBS 0.006466f
C445 B.n405 VSUBS 0.006466f
C446 B.n406 VSUBS 0.006466f
C447 B.n407 VSUBS 0.006466f
C448 B.n408 VSUBS 0.006466f
C449 B.n409 VSUBS 0.006466f
C450 B.n410 VSUBS 0.006466f
C451 B.n411 VSUBS 0.006466f
C452 B.n412 VSUBS 0.006466f
C453 B.n413 VSUBS 0.006466f
C454 B.n414 VSUBS 0.006466f
C455 B.n415 VSUBS 0.006466f
C456 B.n416 VSUBS 0.006466f
C457 B.n417 VSUBS 0.006466f
C458 B.n418 VSUBS 0.006466f
C459 B.n419 VSUBS 0.006466f
C460 B.n420 VSUBS 0.006466f
C461 B.n421 VSUBS 0.006466f
C462 B.n422 VSUBS 0.006466f
C463 B.n423 VSUBS 0.006466f
C464 B.n424 VSUBS 0.006466f
C465 B.n425 VSUBS 0.006466f
C466 B.n426 VSUBS 0.006466f
C467 B.n427 VSUBS 0.006466f
C468 B.n428 VSUBS 0.006466f
C469 B.n429 VSUBS 0.006466f
C470 B.n430 VSUBS 0.006466f
C471 B.n431 VSUBS 0.006466f
C472 B.n432 VSUBS 0.006466f
C473 B.n433 VSUBS 0.006466f
C474 B.n434 VSUBS 0.006466f
C475 B.n435 VSUBS 0.006466f
C476 B.n436 VSUBS 0.006466f
C477 B.n437 VSUBS 0.006466f
C478 B.n438 VSUBS 0.006466f
C479 B.n439 VSUBS 0.006466f
C480 B.n440 VSUBS 0.006466f
C481 B.n441 VSUBS 0.006466f
C482 B.n442 VSUBS 0.006466f
C483 B.n443 VSUBS 0.006466f
C484 B.n444 VSUBS 0.006466f
C485 B.n445 VSUBS 0.006466f
C486 B.n446 VSUBS 0.006466f
C487 B.n447 VSUBS 0.006466f
C488 B.n448 VSUBS 0.006466f
C489 B.n449 VSUBS 0.006466f
C490 B.n450 VSUBS 0.006466f
C491 B.n451 VSUBS 0.006466f
C492 B.n452 VSUBS 0.006466f
C493 B.n453 VSUBS 0.006466f
C494 B.n454 VSUBS 0.006466f
C495 B.n455 VSUBS 0.006466f
C496 B.n456 VSUBS 0.006466f
C497 B.n457 VSUBS 0.004469f
C498 B.n458 VSUBS 0.014982f
C499 B.n459 VSUBS 0.00523f
C500 B.n460 VSUBS 0.006466f
C501 B.n461 VSUBS 0.006466f
C502 B.n462 VSUBS 0.006466f
C503 B.n463 VSUBS 0.006466f
C504 B.n464 VSUBS 0.006466f
C505 B.n465 VSUBS 0.006466f
C506 B.n466 VSUBS 0.006466f
C507 B.n467 VSUBS 0.006466f
C508 B.n468 VSUBS 0.006466f
C509 B.n469 VSUBS 0.006466f
C510 B.n470 VSUBS 0.006466f
C511 B.n471 VSUBS 0.00523f
C512 B.n472 VSUBS 0.006466f
C513 B.n473 VSUBS 0.006466f
C514 B.n474 VSUBS 0.006466f
C515 B.n475 VSUBS 0.006466f
C516 B.n476 VSUBS 0.006466f
C517 B.n477 VSUBS 0.006466f
C518 B.n478 VSUBS 0.006466f
C519 B.n479 VSUBS 0.006466f
C520 B.n480 VSUBS 0.006466f
C521 B.n481 VSUBS 0.006466f
C522 B.n482 VSUBS 0.006466f
C523 B.n483 VSUBS 0.006466f
C524 B.n484 VSUBS 0.006466f
C525 B.n485 VSUBS 0.006466f
C526 B.n486 VSUBS 0.006466f
C527 B.n487 VSUBS 0.006466f
C528 B.n488 VSUBS 0.006466f
C529 B.n489 VSUBS 0.006466f
C530 B.n490 VSUBS 0.006466f
C531 B.n491 VSUBS 0.006466f
C532 B.n492 VSUBS 0.006466f
C533 B.n493 VSUBS 0.006466f
C534 B.n494 VSUBS 0.006466f
C535 B.n495 VSUBS 0.006466f
C536 B.n496 VSUBS 0.006466f
C537 B.n497 VSUBS 0.006466f
C538 B.n498 VSUBS 0.006466f
C539 B.n499 VSUBS 0.006466f
C540 B.n500 VSUBS 0.006466f
C541 B.n501 VSUBS 0.006466f
C542 B.n502 VSUBS 0.006466f
C543 B.n503 VSUBS 0.006466f
C544 B.n504 VSUBS 0.006466f
C545 B.n505 VSUBS 0.006466f
C546 B.n506 VSUBS 0.006466f
C547 B.n507 VSUBS 0.006466f
C548 B.n508 VSUBS 0.006466f
C549 B.n509 VSUBS 0.006466f
C550 B.n510 VSUBS 0.006466f
C551 B.n511 VSUBS 0.006466f
C552 B.n512 VSUBS 0.006466f
C553 B.n513 VSUBS 0.006466f
C554 B.n514 VSUBS 0.006466f
C555 B.n515 VSUBS 0.006466f
C556 B.n516 VSUBS 0.006466f
C557 B.n517 VSUBS 0.006466f
C558 B.n518 VSUBS 0.006466f
C559 B.n519 VSUBS 0.006466f
C560 B.n520 VSUBS 0.006466f
C561 B.n521 VSUBS 0.006466f
C562 B.n522 VSUBS 0.006466f
C563 B.n523 VSUBS 0.006466f
C564 B.n524 VSUBS 0.006466f
C565 B.n525 VSUBS 0.006466f
C566 B.n526 VSUBS 0.006466f
C567 B.n527 VSUBS 0.006466f
C568 B.n528 VSUBS 0.006466f
C569 B.n529 VSUBS 0.006466f
C570 B.n530 VSUBS 0.006466f
C571 B.n531 VSUBS 0.006466f
C572 B.n532 VSUBS 0.006466f
C573 B.n533 VSUBS 0.006466f
C574 B.n534 VSUBS 0.006466f
C575 B.n535 VSUBS 0.006466f
C576 B.n536 VSUBS 0.006466f
C577 B.n537 VSUBS 0.006466f
C578 B.n538 VSUBS 0.006466f
C579 B.n539 VSUBS 0.014299f
C580 B.n540 VSUBS 0.013468f
C581 B.n541 VSUBS 0.013468f
C582 B.n542 VSUBS 0.006466f
C583 B.n543 VSUBS 0.006466f
C584 B.n544 VSUBS 0.006466f
C585 B.n545 VSUBS 0.006466f
C586 B.n546 VSUBS 0.006466f
C587 B.n547 VSUBS 0.006466f
C588 B.n548 VSUBS 0.006466f
C589 B.n549 VSUBS 0.006466f
C590 B.n550 VSUBS 0.006466f
C591 B.n551 VSUBS 0.006466f
C592 B.n552 VSUBS 0.006466f
C593 B.n553 VSUBS 0.006466f
C594 B.n554 VSUBS 0.006466f
C595 B.n555 VSUBS 0.006466f
C596 B.n556 VSUBS 0.006466f
C597 B.n557 VSUBS 0.006466f
C598 B.n558 VSUBS 0.006466f
C599 B.n559 VSUBS 0.006466f
C600 B.n560 VSUBS 0.006466f
C601 B.n561 VSUBS 0.006466f
C602 B.n562 VSUBS 0.006466f
C603 B.n563 VSUBS 0.006466f
C604 B.n564 VSUBS 0.006466f
C605 B.n565 VSUBS 0.006466f
C606 B.n566 VSUBS 0.006466f
C607 B.n567 VSUBS 0.006466f
C608 B.n568 VSUBS 0.006466f
C609 B.n569 VSUBS 0.006466f
C610 B.n570 VSUBS 0.006466f
C611 B.n571 VSUBS 0.014642f
C612 VDD2.t1 VSUBS 2.6739f
C613 VDD2.t0 VSUBS 2.14689f
C614 VDD2.n0 VSUBS 3.19149f
C615 VN.t0 VSUBS 3.13734f
C616 VN.t1 VSUBS 3.60092f
C617 VDD1.t1 VSUBS 2.15659f
C618 VDD1.t0 VSUBS 2.71094f
C619 VTAIL.t2 VSUBS 2.88235f
C620 VTAIL.n0 VSUBS 2.56247f
C621 VTAIL.t0 VSUBS 2.88238f
C622 VTAIL.n1 VSUBS 2.59655f
C623 VTAIL.t3 VSUBS 2.88235f
C624 VTAIL.n2 VSUBS 2.43872f
C625 VTAIL.t1 VSUBS 2.88235f
C626 VTAIL.n3 VSUBS 2.35067f
C627 VP.t0 VSUBS 3.73012f
C628 VP.t1 VSUBS 3.25339f
C629 VP.n0 VSUBS 5.94596f
.ends

