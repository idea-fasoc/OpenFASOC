* NGSPICE file created from diff_pair_sample_1660.ext - technology: sky130A

.subckt diff_pair_sample_1660 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=0.47
X1 VTAIL.t4 VP.t0 VDD1.t5 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=0.47
X2 VDD2.t4 VN.t1 VTAIL.t6 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=0.47
X3 VTAIL.t8 VN.t2 VDD2.t3 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=0.47
X4 VDD2.t2 VN.t3 VTAIL.t9 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=0.47
X5 VTAIL.t0 VP.t1 VDD1.t4 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=0.47
X6 B.t11 B.t9 B.t10 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=0.47
X7 VDD1.t3 VP.t2 VTAIL.t11 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=0.47
X8 B.t8 B.t6 B.t7 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=0.47
X9 VDD1.t2 VP.t3 VTAIL.t2 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=0.47
X10 VTAIL.t5 VN.t4 VDD2.t1 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=0.47
X11 B.t5 B.t3 B.t4 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=0.47
X12 VDD1.t1 VP.t4 VTAIL.t1 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=0.47
X13 VDD2.t0 VN.t5 VTAIL.t10 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=0.47
X14 VDD1.t0 VP.t5 VTAIL.t3 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=0.47
X15 B.t2 B.t0 B.t1 w_n1610_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=0.47
R0 VN.n0 VN.t5 604.673
R1 VN.n4 VN.t3 604.673
R2 VN.n2 VN.t1 587.381
R3 VN.n6 VN.t0 587.381
R4 VN.n1 VN.t2 577.888
R5 VN.n5 VN.t4 577.888
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 72.2473
R9 VN.n3 VN.n0 72.2473
R10 VN VN.n7 39.0327
R11 VN.n2 VN.n1 38.7066
R12 VN.n6 VN.n5 38.7066
R13 VN.n5 VN.n4 17.2717
R14 VN.n1 VN.n0 17.2717
R15 VN VN.n3 0.0516364
R16 VTAIL.n7 VTAIL.t9 65.0987
R17 VTAIL.n11 VTAIL.t6 65.0986
R18 VTAIL.n2 VTAIL.t2 65.0986
R19 VTAIL.n10 VTAIL.t11 65.0986
R20 VTAIL.n9 VTAIL.n8 61.7234
R21 VTAIL.n6 VTAIL.n5 61.7234
R22 VTAIL.n1 VTAIL.n0 61.7232
R23 VTAIL.n4 VTAIL.n3 61.7232
R24 VTAIL.n6 VTAIL.n4 22.0479
R25 VTAIL.n11 VTAIL.n10 21.3583
R26 VTAIL.n0 VTAIL.t10 3.37589
R27 VTAIL.n0 VTAIL.t8 3.37589
R28 VTAIL.n3 VTAIL.t1 3.37589
R29 VTAIL.n3 VTAIL.t0 3.37589
R30 VTAIL.n8 VTAIL.t3 3.37589
R31 VTAIL.n8 VTAIL.t4 3.37589
R32 VTAIL.n5 VTAIL.t7 3.37589
R33 VTAIL.n5 VTAIL.t5 3.37589
R34 VTAIL.n9 VTAIL.n7 0.815155
R35 VTAIL.n2 VTAIL.n1 0.815155
R36 VTAIL.n7 VTAIL.n6 0.690155
R37 VTAIL.n10 VTAIL.n9 0.690155
R38 VTAIL.n4 VTAIL.n2 0.690155
R39 VTAIL VTAIL.n11 0.459552
R40 VTAIL VTAIL.n1 0.231103
R41 VDD2.n1 VDD2.t0 82.2393
R42 VDD2.n2 VDD2.t5 81.7775
R43 VDD2.n1 VDD2.n0 78.519
R44 VDD2 VDD2.n3 78.5162
R45 VDD2.n2 VDD2.n1 34.2584
R46 VDD2.n3 VDD2.t1 3.37589
R47 VDD2.n3 VDD2.t2 3.37589
R48 VDD2.n0 VDD2.t3 3.37589
R49 VDD2.n0 VDD2.t4 3.37589
R50 VDD2 VDD2.n2 0.575931
R51 VP.n1 VP.t5 604.673
R52 VP.n8 VP.t3 587.381
R53 VP.n6 VP.t4 587.381
R54 VP.n3 VP.t2 587.381
R55 VP.n7 VP.t1 577.888
R56 VP.n2 VP.t0 577.888
R57 VP.n9 VP.n8 161.3
R58 VP.n4 VP.n3 161.3
R59 VP.n7 VP.n0 161.3
R60 VP.n6 VP.n5 161.3
R61 VP.n4 VP.n1 72.2473
R62 VP.n7 VP.n6 38.7066
R63 VP.n8 VP.n7 38.7066
R64 VP.n3 VP.n2 38.7066
R65 VP.n5 VP.n4 38.652
R66 VP.n2 VP.n1 17.2717
R67 VP.n5 VP.n0 0.189894
R68 VP.n9 VP.n0 0.189894
R69 VP VP.n9 0.0516364
R70 VDD1 VDD1.t0 82.353
R71 VDD1.n1 VDD1.t1 82.2393
R72 VDD1.n1 VDD1.n0 78.519
R73 VDD1.n3 VDD1.n2 78.402
R74 VDD1.n3 VDD1.n1 35.1862
R75 VDD1.n2 VDD1.t5 3.37589
R76 VDD1.n2 VDD1.t3 3.37589
R77 VDD1.n0 VDD1.t4 3.37589
R78 VDD1.n0 VDD1.t2 3.37589
R79 VDD1 VDD1.n3 0.114724
R80 B.n98 B.t9 700.971
R81 B.n90 B.t3 700.971
R82 B.n36 B.t6 700.971
R83 B.n28 B.t0 700.971
R84 B.n268 B.n267 585
R85 B.n266 B.n73 585
R86 B.n265 B.n264 585
R87 B.n263 B.n74 585
R88 B.n262 B.n261 585
R89 B.n260 B.n75 585
R90 B.n259 B.n258 585
R91 B.n257 B.n76 585
R92 B.n256 B.n255 585
R93 B.n254 B.n77 585
R94 B.n253 B.n252 585
R95 B.n251 B.n78 585
R96 B.n250 B.n249 585
R97 B.n248 B.n79 585
R98 B.n247 B.n246 585
R99 B.n245 B.n80 585
R100 B.n244 B.n243 585
R101 B.n242 B.n81 585
R102 B.n241 B.n240 585
R103 B.n239 B.n82 585
R104 B.n238 B.n237 585
R105 B.n236 B.n83 585
R106 B.n235 B.n234 585
R107 B.n233 B.n84 585
R108 B.n232 B.n231 585
R109 B.n230 B.n85 585
R110 B.n229 B.n228 585
R111 B.n227 B.n86 585
R112 B.n226 B.n225 585
R113 B.n224 B.n87 585
R114 B.n223 B.n222 585
R115 B.n221 B.n88 585
R116 B.n220 B.n219 585
R117 B.n218 B.n89 585
R118 B.n217 B.n216 585
R119 B.n215 B.n214 585
R120 B.n213 B.n93 585
R121 B.n212 B.n211 585
R122 B.n210 B.n94 585
R123 B.n209 B.n208 585
R124 B.n207 B.n95 585
R125 B.n206 B.n205 585
R126 B.n204 B.n96 585
R127 B.n203 B.n202 585
R128 B.n200 B.n97 585
R129 B.n199 B.n198 585
R130 B.n197 B.n100 585
R131 B.n196 B.n195 585
R132 B.n194 B.n101 585
R133 B.n193 B.n192 585
R134 B.n191 B.n102 585
R135 B.n190 B.n189 585
R136 B.n188 B.n103 585
R137 B.n187 B.n186 585
R138 B.n185 B.n104 585
R139 B.n184 B.n183 585
R140 B.n182 B.n105 585
R141 B.n181 B.n180 585
R142 B.n179 B.n106 585
R143 B.n178 B.n177 585
R144 B.n176 B.n107 585
R145 B.n175 B.n174 585
R146 B.n173 B.n108 585
R147 B.n172 B.n171 585
R148 B.n170 B.n109 585
R149 B.n169 B.n168 585
R150 B.n167 B.n110 585
R151 B.n166 B.n165 585
R152 B.n164 B.n111 585
R153 B.n163 B.n162 585
R154 B.n161 B.n112 585
R155 B.n160 B.n159 585
R156 B.n158 B.n113 585
R157 B.n157 B.n156 585
R158 B.n155 B.n114 585
R159 B.n154 B.n153 585
R160 B.n152 B.n115 585
R161 B.n151 B.n150 585
R162 B.n149 B.n116 585
R163 B.n269 B.n72 585
R164 B.n271 B.n270 585
R165 B.n272 B.n71 585
R166 B.n274 B.n273 585
R167 B.n275 B.n70 585
R168 B.n277 B.n276 585
R169 B.n278 B.n69 585
R170 B.n280 B.n279 585
R171 B.n281 B.n68 585
R172 B.n283 B.n282 585
R173 B.n284 B.n67 585
R174 B.n286 B.n285 585
R175 B.n287 B.n66 585
R176 B.n289 B.n288 585
R177 B.n290 B.n65 585
R178 B.n292 B.n291 585
R179 B.n293 B.n64 585
R180 B.n295 B.n294 585
R181 B.n296 B.n63 585
R182 B.n298 B.n297 585
R183 B.n299 B.n62 585
R184 B.n301 B.n300 585
R185 B.n302 B.n61 585
R186 B.n304 B.n303 585
R187 B.n305 B.n60 585
R188 B.n307 B.n306 585
R189 B.n308 B.n59 585
R190 B.n310 B.n309 585
R191 B.n311 B.n58 585
R192 B.n313 B.n312 585
R193 B.n314 B.n57 585
R194 B.n316 B.n315 585
R195 B.n317 B.n56 585
R196 B.n319 B.n318 585
R197 B.n320 B.n55 585
R198 B.n322 B.n321 585
R199 B.n442 B.n441 585
R200 B.n440 B.n11 585
R201 B.n439 B.n438 585
R202 B.n437 B.n12 585
R203 B.n436 B.n435 585
R204 B.n434 B.n13 585
R205 B.n433 B.n432 585
R206 B.n431 B.n14 585
R207 B.n430 B.n429 585
R208 B.n428 B.n15 585
R209 B.n427 B.n426 585
R210 B.n425 B.n16 585
R211 B.n424 B.n423 585
R212 B.n422 B.n17 585
R213 B.n421 B.n420 585
R214 B.n419 B.n18 585
R215 B.n418 B.n417 585
R216 B.n416 B.n19 585
R217 B.n415 B.n414 585
R218 B.n413 B.n20 585
R219 B.n412 B.n411 585
R220 B.n410 B.n21 585
R221 B.n409 B.n408 585
R222 B.n407 B.n22 585
R223 B.n406 B.n405 585
R224 B.n404 B.n23 585
R225 B.n403 B.n402 585
R226 B.n401 B.n24 585
R227 B.n400 B.n399 585
R228 B.n398 B.n25 585
R229 B.n397 B.n396 585
R230 B.n395 B.n26 585
R231 B.n394 B.n393 585
R232 B.n392 B.n27 585
R233 B.n391 B.n390 585
R234 B.n389 B.n388 585
R235 B.n387 B.n31 585
R236 B.n386 B.n385 585
R237 B.n384 B.n32 585
R238 B.n383 B.n382 585
R239 B.n381 B.n33 585
R240 B.n380 B.n379 585
R241 B.n378 B.n34 585
R242 B.n377 B.n376 585
R243 B.n374 B.n35 585
R244 B.n373 B.n372 585
R245 B.n371 B.n38 585
R246 B.n370 B.n369 585
R247 B.n368 B.n39 585
R248 B.n367 B.n366 585
R249 B.n365 B.n40 585
R250 B.n364 B.n363 585
R251 B.n362 B.n41 585
R252 B.n361 B.n360 585
R253 B.n359 B.n42 585
R254 B.n358 B.n357 585
R255 B.n356 B.n43 585
R256 B.n355 B.n354 585
R257 B.n353 B.n44 585
R258 B.n352 B.n351 585
R259 B.n350 B.n45 585
R260 B.n349 B.n348 585
R261 B.n347 B.n46 585
R262 B.n346 B.n345 585
R263 B.n344 B.n47 585
R264 B.n343 B.n342 585
R265 B.n341 B.n48 585
R266 B.n340 B.n339 585
R267 B.n338 B.n49 585
R268 B.n337 B.n336 585
R269 B.n335 B.n50 585
R270 B.n334 B.n333 585
R271 B.n332 B.n51 585
R272 B.n331 B.n330 585
R273 B.n329 B.n52 585
R274 B.n328 B.n327 585
R275 B.n326 B.n53 585
R276 B.n325 B.n324 585
R277 B.n323 B.n54 585
R278 B.n443 B.n10 585
R279 B.n445 B.n444 585
R280 B.n446 B.n9 585
R281 B.n448 B.n447 585
R282 B.n449 B.n8 585
R283 B.n451 B.n450 585
R284 B.n452 B.n7 585
R285 B.n454 B.n453 585
R286 B.n455 B.n6 585
R287 B.n457 B.n456 585
R288 B.n458 B.n5 585
R289 B.n460 B.n459 585
R290 B.n461 B.n4 585
R291 B.n463 B.n462 585
R292 B.n464 B.n3 585
R293 B.n466 B.n465 585
R294 B.n467 B.n0 585
R295 B.n2 B.n1 585
R296 B.n125 B.n124 585
R297 B.n127 B.n126 585
R298 B.n128 B.n123 585
R299 B.n130 B.n129 585
R300 B.n131 B.n122 585
R301 B.n133 B.n132 585
R302 B.n134 B.n121 585
R303 B.n136 B.n135 585
R304 B.n137 B.n120 585
R305 B.n139 B.n138 585
R306 B.n140 B.n119 585
R307 B.n142 B.n141 585
R308 B.n143 B.n118 585
R309 B.n145 B.n144 585
R310 B.n146 B.n117 585
R311 B.n148 B.n147 585
R312 B.n149 B.n148 492.5
R313 B.n269 B.n268 492.5
R314 B.n323 B.n322 492.5
R315 B.n443 B.n442 492.5
R316 B.n469 B.n468 256.663
R317 B.n468 B.n467 235.042
R318 B.n468 B.n2 235.042
R319 B.n150 B.n149 163.367
R320 B.n150 B.n115 163.367
R321 B.n154 B.n115 163.367
R322 B.n155 B.n154 163.367
R323 B.n156 B.n155 163.367
R324 B.n156 B.n113 163.367
R325 B.n160 B.n113 163.367
R326 B.n161 B.n160 163.367
R327 B.n162 B.n161 163.367
R328 B.n162 B.n111 163.367
R329 B.n166 B.n111 163.367
R330 B.n167 B.n166 163.367
R331 B.n168 B.n167 163.367
R332 B.n168 B.n109 163.367
R333 B.n172 B.n109 163.367
R334 B.n173 B.n172 163.367
R335 B.n174 B.n173 163.367
R336 B.n174 B.n107 163.367
R337 B.n178 B.n107 163.367
R338 B.n179 B.n178 163.367
R339 B.n180 B.n179 163.367
R340 B.n180 B.n105 163.367
R341 B.n184 B.n105 163.367
R342 B.n185 B.n184 163.367
R343 B.n186 B.n185 163.367
R344 B.n186 B.n103 163.367
R345 B.n190 B.n103 163.367
R346 B.n191 B.n190 163.367
R347 B.n192 B.n191 163.367
R348 B.n192 B.n101 163.367
R349 B.n196 B.n101 163.367
R350 B.n197 B.n196 163.367
R351 B.n198 B.n197 163.367
R352 B.n198 B.n97 163.367
R353 B.n203 B.n97 163.367
R354 B.n204 B.n203 163.367
R355 B.n205 B.n204 163.367
R356 B.n205 B.n95 163.367
R357 B.n209 B.n95 163.367
R358 B.n210 B.n209 163.367
R359 B.n211 B.n210 163.367
R360 B.n211 B.n93 163.367
R361 B.n215 B.n93 163.367
R362 B.n216 B.n215 163.367
R363 B.n216 B.n89 163.367
R364 B.n220 B.n89 163.367
R365 B.n221 B.n220 163.367
R366 B.n222 B.n221 163.367
R367 B.n222 B.n87 163.367
R368 B.n226 B.n87 163.367
R369 B.n227 B.n226 163.367
R370 B.n228 B.n227 163.367
R371 B.n228 B.n85 163.367
R372 B.n232 B.n85 163.367
R373 B.n233 B.n232 163.367
R374 B.n234 B.n233 163.367
R375 B.n234 B.n83 163.367
R376 B.n238 B.n83 163.367
R377 B.n239 B.n238 163.367
R378 B.n240 B.n239 163.367
R379 B.n240 B.n81 163.367
R380 B.n244 B.n81 163.367
R381 B.n245 B.n244 163.367
R382 B.n246 B.n245 163.367
R383 B.n246 B.n79 163.367
R384 B.n250 B.n79 163.367
R385 B.n251 B.n250 163.367
R386 B.n252 B.n251 163.367
R387 B.n252 B.n77 163.367
R388 B.n256 B.n77 163.367
R389 B.n257 B.n256 163.367
R390 B.n258 B.n257 163.367
R391 B.n258 B.n75 163.367
R392 B.n262 B.n75 163.367
R393 B.n263 B.n262 163.367
R394 B.n264 B.n263 163.367
R395 B.n264 B.n73 163.367
R396 B.n268 B.n73 163.367
R397 B.n322 B.n55 163.367
R398 B.n318 B.n55 163.367
R399 B.n318 B.n317 163.367
R400 B.n317 B.n316 163.367
R401 B.n316 B.n57 163.367
R402 B.n312 B.n57 163.367
R403 B.n312 B.n311 163.367
R404 B.n311 B.n310 163.367
R405 B.n310 B.n59 163.367
R406 B.n306 B.n59 163.367
R407 B.n306 B.n305 163.367
R408 B.n305 B.n304 163.367
R409 B.n304 B.n61 163.367
R410 B.n300 B.n61 163.367
R411 B.n300 B.n299 163.367
R412 B.n299 B.n298 163.367
R413 B.n298 B.n63 163.367
R414 B.n294 B.n63 163.367
R415 B.n294 B.n293 163.367
R416 B.n293 B.n292 163.367
R417 B.n292 B.n65 163.367
R418 B.n288 B.n65 163.367
R419 B.n288 B.n287 163.367
R420 B.n287 B.n286 163.367
R421 B.n286 B.n67 163.367
R422 B.n282 B.n67 163.367
R423 B.n282 B.n281 163.367
R424 B.n281 B.n280 163.367
R425 B.n280 B.n69 163.367
R426 B.n276 B.n69 163.367
R427 B.n276 B.n275 163.367
R428 B.n275 B.n274 163.367
R429 B.n274 B.n71 163.367
R430 B.n270 B.n71 163.367
R431 B.n270 B.n269 163.367
R432 B.n442 B.n11 163.367
R433 B.n438 B.n11 163.367
R434 B.n438 B.n437 163.367
R435 B.n437 B.n436 163.367
R436 B.n436 B.n13 163.367
R437 B.n432 B.n13 163.367
R438 B.n432 B.n431 163.367
R439 B.n431 B.n430 163.367
R440 B.n430 B.n15 163.367
R441 B.n426 B.n15 163.367
R442 B.n426 B.n425 163.367
R443 B.n425 B.n424 163.367
R444 B.n424 B.n17 163.367
R445 B.n420 B.n17 163.367
R446 B.n420 B.n419 163.367
R447 B.n419 B.n418 163.367
R448 B.n418 B.n19 163.367
R449 B.n414 B.n19 163.367
R450 B.n414 B.n413 163.367
R451 B.n413 B.n412 163.367
R452 B.n412 B.n21 163.367
R453 B.n408 B.n21 163.367
R454 B.n408 B.n407 163.367
R455 B.n407 B.n406 163.367
R456 B.n406 B.n23 163.367
R457 B.n402 B.n23 163.367
R458 B.n402 B.n401 163.367
R459 B.n401 B.n400 163.367
R460 B.n400 B.n25 163.367
R461 B.n396 B.n25 163.367
R462 B.n396 B.n395 163.367
R463 B.n395 B.n394 163.367
R464 B.n394 B.n27 163.367
R465 B.n390 B.n27 163.367
R466 B.n390 B.n389 163.367
R467 B.n389 B.n31 163.367
R468 B.n385 B.n31 163.367
R469 B.n385 B.n384 163.367
R470 B.n384 B.n383 163.367
R471 B.n383 B.n33 163.367
R472 B.n379 B.n33 163.367
R473 B.n379 B.n378 163.367
R474 B.n378 B.n377 163.367
R475 B.n377 B.n35 163.367
R476 B.n372 B.n35 163.367
R477 B.n372 B.n371 163.367
R478 B.n371 B.n370 163.367
R479 B.n370 B.n39 163.367
R480 B.n366 B.n39 163.367
R481 B.n366 B.n365 163.367
R482 B.n365 B.n364 163.367
R483 B.n364 B.n41 163.367
R484 B.n360 B.n41 163.367
R485 B.n360 B.n359 163.367
R486 B.n359 B.n358 163.367
R487 B.n358 B.n43 163.367
R488 B.n354 B.n43 163.367
R489 B.n354 B.n353 163.367
R490 B.n353 B.n352 163.367
R491 B.n352 B.n45 163.367
R492 B.n348 B.n45 163.367
R493 B.n348 B.n347 163.367
R494 B.n347 B.n346 163.367
R495 B.n346 B.n47 163.367
R496 B.n342 B.n47 163.367
R497 B.n342 B.n341 163.367
R498 B.n341 B.n340 163.367
R499 B.n340 B.n49 163.367
R500 B.n336 B.n49 163.367
R501 B.n336 B.n335 163.367
R502 B.n335 B.n334 163.367
R503 B.n334 B.n51 163.367
R504 B.n330 B.n51 163.367
R505 B.n330 B.n329 163.367
R506 B.n329 B.n328 163.367
R507 B.n328 B.n53 163.367
R508 B.n324 B.n53 163.367
R509 B.n324 B.n323 163.367
R510 B.n444 B.n443 163.367
R511 B.n444 B.n9 163.367
R512 B.n448 B.n9 163.367
R513 B.n449 B.n448 163.367
R514 B.n450 B.n449 163.367
R515 B.n450 B.n7 163.367
R516 B.n454 B.n7 163.367
R517 B.n455 B.n454 163.367
R518 B.n456 B.n455 163.367
R519 B.n456 B.n5 163.367
R520 B.n460 B.n5 163.367
R521 B.n461 B.n460 163.367
R522 B.n462 B.n461 163.367
R523 B.n462 B.n3 163.367
R524 B.n466 B.n3 163.367
R525 B.n467 B.n466 163.367
R526 B.n125 B.n2 163.367
R527 B.n126 B.n125 163.367
R528 B.n126 B.n123 163.367
R529 B.n130 B.n123 163.367
R530 B.n131 B.n130 163.367
R531 B.n132 B.n131 163.367
R532 B.n132 B.n121 163.367
R533 B.n136 B.n121 163.367
R534 B.n137 B.n136 163.367
R535 B.n138 B.n137 163.367
R536 B.n138 B.n119 163.367
R537 B.n142 B.n119 163.367
R538 B.n143 B.n142 163.367
R539 B.n144 B.n143 163.367
R540 B.n144 B.n117 163.367
R541 B.n148 B.n117 163.367
R542 B.n90 B.t4 125.463
R543 B.n36 B.t8 125.463
R544 B.n98 B.t10 125.453
R545 B.n28 B.t2 125.453
R546 B.n91 B.t5 109.948
R547 B.n37 B.t7 109.948
R548 B.n99 B.t11 109.938
R549 B.n29 B.t1 109.938
R550 B.n201 B.n99 59.5399
R551 B.n92 B.n91 59.5399
R552 B.n375 B.n37 59.5399
R553 B.n30 B.n29 59.5399
R554 B.n441 B.n10 32.0005
R555 B.n321 B.n54 32.0005
R556 B.n267 B.n72 32.0005
R557 B.n147 B.n116 32.0005
R558 B B.n469 18.0485
R559 B.n99 B.n98 15.5157
R560 B.n91 B.n90 15.5157
R561 B.n37 B.n36 15.5157
R562 B.n29 B.n28 15.5157
R563 B.n445 B.n10 10.6151
R564 B.n446 B.n445 10.6151
R565 B.n447 B.n446 10.6151
R566 B.n447 B.n8 10.6151
R567 B.n451 B.n8 10.6151
R568 B.n452 B.n451 10.6151
R569 B.n453 B.n452 10.6151
R570 B.n453 B.n6 10.6151
R571 B.n457 B.n6 10.6151
R572 B.n458 B.n457 10.6151
R573 B.n459 B.n458 10.6151
R574 B.n459 B.n4 10.6151
R575 B.n463 B.n4 10.6151
R576 B.n464 B.n463 10.6151
R577 B.n465 B.n464 10.6151
R578 B.n465 B.n0 10.6151
R579 B.n441 B.n440 10.6151
R580 B.n440 B.n439 10.6151
R581 B.n439 B.n12 10.6151
R582 B.n435 B.n12 10.6151
R583 B.n435 B.n434 10.6151
R584 B.n434 B.n433 10.6151
R585 B.n433 B.n14 10.6151
R586 B.n429 B.n14 10.6151
R587 B.n429 B.n428 10.6151
R588 B.n428 B.n427 10.6151
R589 B.n427 B.n16 10.6151
R590 B.n423 B.n16 10.6151
R591 B.n423 B.n422 10.6151
R592 B.n422 B.n421 10.6151
R593 B.n421 B.n18 10.6151
R594 B.n417 B.n18 10.6151
R595 B.n417 B.n416 10.6151
R596 B.n416 B.n415 10.6151
R597 B.n415 B.n20 10.6151
R598 B.n411 B.n20 10.6151
R599 B.n411 B.n410 10.6151
R600 B.n410 B.n409 10.6151
R601 B.n409 B.n22 10.6151
R602 B.n405 B.n22 10.6151
R603 B.n405 B.n404 10.6151
R604 B.n404 B.n403 10.6151
R605 B.n403 B.n24 10.6151
R606 B.n399 B.n24 10.6151
R607 B.n399 B.n398 10.6151
R608 B.n398 B.n397 10.6151
R609 B.n397 B.n26 10.6151
R610 B.n393 B.n26 10.6151
R611 B.n393 B.n392 10.6151
R612 B.n392 B.n391 10.6151
R613 B.n388 B.n387 10.6151
R614 B.n387 B.n386 10.6151
R615 B.n386 B.n32 10.6151
R616 B.n382 B.n32 10.6151
R617 B.n382 B.n381 10.6151
R618 B.n381 B.n380 10.6151
R619 B.n380 B.n34 10.6151
R620 B.n376 B.n34 10.6151
R621 B.n374 B.n373 10.6151
R622 B.n373 B.n38 10.6151
R623 B.n369 B.n38 10.6151
R624 B.n369 B.n368 10.6151
R625 B.n368 B.n367 10.6151
R626 B.n367 B.n40 10.6151
R627 B.n363 B.n40 10.6151
R628 B.n363 B.n362 10.6151
R629 B.n362 B.n361 10.6151
R630 B.n361 B.n42 10.6151
R631 B.n357 B.n42 10.6151
R632 B.n357 B.n356 10.6151
R633 B.n356 B.n355 10.6151
R634 B.n355 B.n44 10.6151
R635 B.n351 B.n44 10.6151
R636 B.n351 B.n350 10.6151
R637 B.n350 B.n349 10.6151
R638 B.n349 B.n46 10.6151
R639 B.n345 B.n46 10.6151
R640 B.n345 B.n344 10.6151
R641 B.n344 B.n343 10.6151
R642 B.n343 B.n48 10.6151
R643 B.n339 B.n48 10.6151
R644 B.n339 B.n338 10.6151
R645 B.n338 B.n337 10.6151
R646 B.n337 B.n50 10.6151
R647 B.n333 B.n50 10.6151
R648 B.n333 B.n332 10.6151
R649 B.n332 B.n331 10.6151
R650 B.n331 B.n52 10.6151
R651 B.n327 B.n52 10.6151
R652 B.n327 B.n326 10.6151
R653 B.n326 B.n325 10.6151
R654 B.n325 B.n54 10.6151
R655 B.n321 B.n320 10.6151
R656 B.n320 B.n319 10.6151
R657 B.n319 B.n56 10.6151
R658 B.n315 B.n56 10.6151
R659 B.n315 B.n314 10.6151
R660 B.n314 B.n313 10.6151
R661 B.n313 B.n58 10.6151
R662 B.n309 B.n58 10.6151
R663 B.n309 B.n308 10.6151
R664 B.n308 B.n307 10.6151
R665 B.n307 B.n60 10.6151
R666 B.n303 B.n60 10.6151
R667 B.n303 B.n302 10.6151
R668 B.n302 B.n301 10.6151
R669 B.n301 B.n62 10.6151
R670 B.n297 B.n62 10.6151
R671 B.n297 B.n296 10.6151
R672 B.n296 B.n295 10.6151
R673 B.n295 B.n64 10.6151
R674 B.n291 B.n64 10.6151
R675 B.n291 B.n290 10.6151
R676 B.n290 B.n289 10.6151
R677 B.n289 B.n66 10.6151
R678 B.n285 B.n66 10.6151
R679 B.n285 B.n284 10.6151
R680 B.n284 B.n283 10.6151
R681 B.n283 B.n68 10.6151
R682 B.n279 B.n68 10.6151
R683 B.n279 B.n278 10.6151
R684 B.n278 B.n277 10.6151
R685 B.n277 B.n70 10.6151
R686 B.n273 B.n70 10.6151
R687 B.n273 B.n272 10.6151
R688 B.n272 B.n271 10.6151
R689 B.n271 B.n72 10.6151
R690 B.n124 B.n1 10.6151
R691 B.n127 B.n124 10.6151
R692 B.n128 B.n127 10.6151
R693 B.n129 B.n128 10.6151
R694 B.n129 B.n122 10.6151
R695 B.n133 B.n122 10.6151
R696 B.n134 B.n133 10.6151
R697 B.n135 B.n134 10.6151
R698 B.n135 B.n120 10.6151
R699 B.n139 B.n120 10.6151
R700 B.n140 B.n139 10.6151
R701 B.n141 B.n140 10.6151
R702 B.n141 B.n118 10.6151
R703 B.n145 B.n118 10.6151
R704 B.n146 B.n145 10.6151
R705 B.n147 B.n146 10.6151
R706 B.n151 B.n116 10.6151
R707 B.n152 B.n151 10.6151
R708 B.n153 B.n152 10.6151
R709 B.n153 B.n114 10.6151
R710 B.n157 B.n114 10.6151
R711 B.n158 B.n157 10.6151
R712 B.n159 B.n158 10.6151
R713 B.n159 B.n112 10.6151
R714 B.n163 B.n112 10.6151
R715 B.n164 B.n163 10.6151
R716 B.n165 B.n164 10.6151
R717 B.n165 B.n110 10.6151
R718 B.n169 B.n110 10.6151
R719 B.n170 B.n169 10.6151
R720 B.n171 B.n170 10.6151
R721 B.n171 B.n108 10.6151
R722 B.n175 B.n108 10.6151
R723 B.n176 B.n175 10.6151
R724 B.n177 B.n176 10.6151
R725 B.n177 B.n106 10.6151
R726 B.n181 B.n106 10.6151
R727 B.n182 B.n181 10.6151
R728 B.n183 B.n182 10.6151
R729 B.n183 B.n104 10.6151
R730 B.n187 B.n104 10.6151
R731 B.n188 B.n187 10.6151
R732 B.n189 B.n188 10.6151
R733 B.n189 B.n102 10.6151
R734 B.n193 B.n102 10.6151
R735 B.n194 B.n193 10.6151
R736 B.n195 B.n194 10.6151
R737 B.n195 B.n100 10.6151
R738 B.n199 B.n100 10.6151
R739 B.n200 B.n199 10.6151
R740 B.n202 B.n96 10.6151
R741 B.n206 B.n96 10.6151
R742 B.n207 B.n206 10.6151
R743 B.n208 B.n207 10.6151
R744 B.n208 B.n94 10.6151
R745 B.n212 B.n94 10.6151
R746 B.n213 B.n212 10.6151
R747 B.n214 B.n213 10.6151
R748 B.n218 B.n217 10.6151
R749 B.n219 B.n218 10.6151
R750 B.n219 B.n88 10.6151
R751 B.n223 B.n88 10.6151
R752 B.n224 B.n223 10.6151
R753 B.n225 B.n224 10.6151
R754 B.n225 B.n86 10.6151
R755 B.n229 B.n86 10.6151
R756 B.n230 B.n229 10.6151
R757 B.n231 B.n230 10.6151
R758 B.n231 B.n84 10.6151
R759 B.n235 B.n84 10.6151
R760 B.n236 B.n235 10.6151
R761 B.n237 B.n236 10.6151
R762 B.n237 B.n82 10.6151
R763 B.n241 B.n82 10.6151
R764 B.n242 B.n241 10.6151
R765 B.n243 B.n242 10.6151
R766 B.n243 B.n80 10.6151
R767 B.n247 B.n80 10.6151
R768 B.n248 B.n247 10.6151
R769 B.n249 B.n248 10.6151
R770 B.n249 B.n78 10.6151
R771 B.n253 B.n78 10.6151
R772 B.n254 B.n253 10.6151
R773 B.n255 B.n254 10.6151
R774 B.n255 B.n76 10.6151
R775 B.n259 B.n76 10.6151
R776 B.n260 B.n259 10.6151
R777 B.n261 B.n260 10.6151
R778 B.n261 B.n74 10.6151
R779 B.n265 B.n74 10.6151
R780 B.n266 B.n265 10.6151
R781 B.n267 B.n266 10.6151
R782 B.n469 B.n0 8.11757
R783 B.n469 B.n1 8.11757
R784 B.n388 B.n30 6.5566
R785 B.n376 B.n375 6.5566
R786 B.n202 B.n201 6.5566
R787 B.n214 B.n92 6.5566
R788 B.n391 B.n30 4.05904
R789 B.n375 B.n374 4.05904
R790 B.n201 B.n200 4.05904
R791 B.n217 B.n92 4.05904
C0 VN B 0.686436f
C1 VDD2 VN 2.88302f
C2 VDD1 VTAIL 9.65638f
C3 VDD2 B 1.34188f
C4 VDD1 VP 3.00907f
C5 VDD1 w_n1610_n2894# 1.5682f
C6 VN VTAIL 2.59033f
C7 VP VN 4.41433f
C8 B VTAIL 2.14664f
C9 VDD2 VTAIL 9.68941f
C10 w_n1610_n2894# VN 2.48112f
C11 VP B 1.01333f
C12 VP VDD2 0.277784f
C13 w_n1610_n2894# B 6.07307f
C14 w_n1610_n2894# VDD2 1.58529f
C15 VDD1 VN 0.147758f
C16 VDD1 B 1.31818f
C17 VP VTAIL 2.6049f
C18 VDD1 VDD2 0.627839f
C19 w_n1610_n2894# VTAIL 2.57203f
C20 VP w_n1610_n2894# 2.68333f
C21 VDD2 VSUBS 1.210604f
C22 VDD1 VSUBS 1.468469f
C23 VTAIL VSUBS 0.605105f
C24 VN VSUBS 4.211451f
C25 VP VSUBS 1.217411f
C26 B VSUBS 2.316619f
C27 w_n1610_n2894# VSUBS 57.5929f
C28 B.n0 VSUBS 0.006943f
C29 B.n1 VSUBS 0.006943f
C30 B.n2 VSUBS 0.010269f
C31 B.n3 VSUBS 0.007869f
C32 B.n4 VSUBS 0.007869f
C33 B.n5 VSUBS 0.007869f
C34 B.n6 VSUBS 0.007869f
C35 B.n7 VSUBS 0.007869f
C36 B.n8 VSUBS 0.007869f
C37 B.n9 VSUBS 0.007869f
C38 B.n10 VSUBS 0.017648f
C39 B.n11 VSUBS 0.007869f
C40 B.n12 VSUBS 0.007869f
C41 B.n13 VSUBS 0.007869f
C42 B.n14 VSUBS 0.007869f
C43 B.n15 VSUBS 0.007869f
C44 B.n16 VSUBS 0.007869f
C45 B.n17 VSUBS 0.007869f
C46 B.n18 VSUBS 0.007869f
C47 B.n19 VSUBS 0.007869f
C48 B.n20 VSUBS 0.007869f
C49 B.n21 VSUBS 0.007869f
C50 B.n22 VSUBS 0.007869f
C51 B.n23 VSUBS 0.007869f
C52 B.n24 VSUBS 0.007869f
C53 B.n25 VSUBS 0.007869f
C54 B.n26 VSUBS 0.007869f
C55 B.n27 VSUBS 0.007869f
C56 B.t1 VSUBS 0.343523f
C57 B.t2 VSUBS 0.350861f
C58 B.t0 VSUBS 0.207093f
C59 B.n28 VSUBS 0.113997f
C60 B.n29 VSUBS 0.070557f
C61 B.n30 VSUBS 0.018232f
C62 B.n31 VSUBS 0.007869f
C63 B.n32 VSUBS 0.007869f
C64 B.n33 VSUBS 0.007869f
C65 B.n34 VSUBS 0.007869f
C66 B.n35 VSUBS 0.007869f
C67 B.t7 VSUBS 0.343519f
C68 B.t8 VSUBS 0.350857f
C69 B.t6 VSUBS 0.207093f
C70 B.n36 VSUBS 0.114002f
C71 B.n37 VSUBS 0.070561f
C72 B.n38 VSUBS 0.007869f
C73 B.n39 VSUBS 0.007869f
C74 B.n40 VSUBS 0.007869f
C75 B.n41 VSUBS 0.007869f
C76 B.n42 VSUBS 0.007869f
C77 B.n43 VSUBS 0.007869f
C78 B.n44 VSUBS 0.007869f
C79 B.n45 VSUBS 0.007869f
C80 B.n46 VSUBS 0.007869f
C81 B.n47 VSUBS 0.007869f
C82 B.n48 VSUBS 0.007869f
C83 B.n49 VSUBS 0.007869f
C84 B.n50 VSUBS 0.007869f
C85 B.n51 VSUBS 0.007869f
C86 B.n52 VSUBS 0.007869f
C87 B.n53 VSUBS 0.007869f
C88 B.n54 VSUBS 0.018689f
C89 B.n55 VSUBS 0.007869f
C90 B.n56 VSUBS 0.007869f
C91 B.n57 VSUBS 0.007869f
C92 B.n58 VSUBS 0.007869f
C93 B.n59 VSUBS 0.007869f
C94 B.n60 VSUBS 0.007869f
C95 B.n61 VSUBS 0.007869f
C96 B.n62 VSUBS 0.007869f
C97 B.n63 VSUBS 0.007869f
C98 B.n64 VSUBS 0.007869f
C99 B.n65 VSUBS 0.007869f
C100 B.n66 VSUBS 0.007869f
C101 B.n67 VSUBS 0.007869f
C102 B.n68 VSUBS 0.007869f
C103 B.n69 VSUBS 0.007869f
C104 B.n70 VSUBS 0.007869f
C105 B.n71 VSUBS 0.007869f
C106 B.n72 VSUBS 0.018597f
C107 B.n73 VSUBS 0.007869f
C108 B.n74 VSUBS 0.007869f
C109 B.n75 VSUBS 0.007869f
C110 B.n76 VSUBS 0.007869f
C111 B.n77 VSUBS 0.007869f
C112 B.n78 VSUBS 0.007869f
C113 B.n79 VSUBS 0.007869f
C114 B.n80 VSUBS 0.007869f
C115 B.n81 VSUBS 0.007869f
C116 B.n82 VSUBS 0.007869f
C117 B.n83 VSUBS 0.007869f
C118 B.n84 VSUBS 0.007869f
C119 B.n85 VSUBS 0.007869f
C120 B.n86 VSUBS 0.007869f
C121 B.n87 VSUBS 0.007869f
C122 B.n88 VSUBS 0.007869f
C123 B.n89 VSUBS 0.007869f
C124 B.t5 VSUBS 0.343519f
C125 B.t4 VSUBS 0.350857f
C126 B.t3 VSUBS 0.207093f
C127 B.n90 VSUBS 0.114002f
C128 B.n91 VSUBS 0.070561f
C129 B.n92 VSUBS 0.018232f
C130 B.n93 VSUBS 0.007869f
C131 B.n94 VSUBS 0.007869f
C132 B.n95 VSUBS 0.007869f
C133 B.n96 VSUBS 0.007869f
C134 B.n97 VSUBS 0.007869f
C135 B.t11 VSUBS 0.343523f
C136 B.t10 VSUBS 0.350861f
C137 B.t9 VSUBS 0.207093f
C138 B.n98 VSUBS 0.113997f
C139 B.n99 VSUBS 0.070557f
C140 B.n100 VSUBS 0.007869f
C141 B.n101 VSUBS 0.007869f
C142 B.n102 VSUBS 0.007869f
C143 B.n103 VSUBS 0.007869f
C144 B.n104 VSUBS 0.007869f
C145 B.n105 VSUBS 0.007869f
C146 B.n106 VSUBS 0.007869f
C147 B.n107 VSUBS 0.007869f
C148 B.n108 VSUBS 0.007869f
C149 B.n109 VSUBS 0.007869f
C150 B.n110 VSUBS 0.007869f
C151 B.n111 VSUBS 0.007869f
C152 B.n112 VSUBS 0.007869f
C153 B.n113 VSUBS 0.007869f
C154 B.n114 VSUBS 0.007869f
C155 B.n115 VSUBS 0.007869f
C156 B.n116 VSUBS 0.018689f
C157 B.n117 VSUBS 0.007869f
C158 B.n118 VSUBS 0.007869f
C159 B.n119 VSUBS 0.007869f
C160 B.n120 VSUBS 0.007869f
C161 B.n121 VSUBS 0.007869f
C162 B.n122 VSUBS 0.007869f
C163 B.n123 VSUBS 0.007869f
C164 B.n124 VSUBS 0.007869f
C165 B.n125 VSUBS 0.007869f
C166 B.n126 VSUBS 0.007869f
C167 B.n127 VSUBS 0.007869f
C168 B.n128 VSUBS 0.007869f
C169 B.n129 VSUBS 0.007869f
C170 B.n130 VSUBS 0.007869f
C171 B.n131 VSUBS 0.007869f
C172 B.n132 VSUBS 0.007869f
C173 B.n133 VSUBS 0.007869f
C174 B.n134 VSUBS 0.007869f
C175 B.n135 VSUBS 0.007869f
C176 B.n136 VSUBS 0.007869f
C177 B.n137 VSUBS 0.007869f
C178 B.n138 VSUBS 0.007869f
C179 B.n139 VSUBS 0.007869f
C180 B.n140 VSUBS 0.007869f
C181 B.n141 VSUBS 0.007869f
C182 B.n142 VSUBS 0.007869f
C183 B.n143 VSUBS 0.007869f
C184 B.n144 VSUBS 0.007869f
C185 B.n145 VSUBS 0.007869f
C186 B.n146 VSUBS 0.007869f
C187 B.n147 VSUBS 0.017648f
C188 B.n148 VSUBS 0.017648f
C189 B.n149 VSUBS 0.018689f
C190 B.n150 VSUBS 0.007869f
C191 B.n151 VSUBS 0.007869f
C192 B.n152 VSUBS 0.007869f
C193 B.n153 VSUBS 0.007869f
C194 B.n154 VSUBS 0.007869f
C195 B.n155 VSUBS 0.007869f
C196 B.n156 VSUBS 0.007869f
C197 B.n157 VSUBS 0.007869f
C198 B.n158 VSUBS 0.007869f
C199 B.n159 VSUBS 0.007869f
C200 B.n160 VSUBS 0.007869f
C201 B.n161 VSUBS 0.007869f
C202 B.n162 VSUBS 0.007869f
C203 B.n163 VSUBS 0.007869f
C204 B.n164 VSUBS 0.007869f
C205 B.n165 VSUBS 0.007869f
C206 B.n166 VSUBS 0.007869f
C207 B.n167 VSUBS 0.007869f
C208 B.n168 VSUBS 0.007869f
C209 B.n169 VSUBS 0.007869f
C210 B.n170 VSUBS 0.007869f
C211 B.n171 VSUBS 0.007869f
C212 B.n172 VSUBS 0.007869f
C213 B.n173 VSUBS 0.007869f
C214 B.n174 VSUBS 0.007869f
C215 B.n175 VSUBS 0.007869f
C216 B.n176 VSUBS 0.007869f
C217 B.n177 VSUBS 0.007869f
C218 B.n178 VSUBS 0.007869f
C219 B.n179 VSUBS 0.007869f
C220 B.n180 VSUBS 0.007869f
C221 B.n181 VSUBS 0.007869f
C222 B.n182 VSUBS 0.007869f
C223 B.n183 VSUBS 0.007869f
C224 B.n184 VSUBS 0.007869f
C225 B.n185 VSUBS 0.007869f
C226 B.n186 VSUBS 0.007869f
C227 B.n187 VSUBS 0.007869f
C228 B.n188 VSUBS 0.007869f
C229 B.n189 VSUBS 0.007869f
C230 B.n190 VSUBS 0.007869f
C231 B.n191 VSUBS 0.007869f
C232 B.n192 VSUBS 0.007869f
C233 B.n193 VSUBS 0.007869f
C234 B.n194 VSUBS 0.007869f
C235 B.n195 VSUBS 0.007869f
C236 B.n196 VSUBS 0.007869f
C237 B.n197 VSUBS 0.007869f
C238 B.n198 VSUBS 0.007869f
C239 B.n199 VSUBS 0.007869f
C240 B.n200 VSUBS 0.005439f
C241 B.n201 VSUBS 0.018232f
C242 B.n202 VSUBS 0.006365f
C243 B.n203 VSUBS 0.007869f
C244 B.n204 VSUBS 0.007869f
C245 B.n205 VSUBS 0.007869f
C246 B.n206 VSUBS 0.007869f
C247 B.n207 VSUBS 0.007869f
C248 B.n208 VSUBS 0.007869f
C249 B.n209 VSUBS 0.007869f
C250 B.n210 VSUBS 0.007869f
C251 B.n211 VSUBS 0.007869f
C252 B.n212 VSUBS 0.007869f
C253 B.n213 VSUBS 0.007869f
C254 B.n214 VSUBS 0.006365f
C255 B.n215 VSUBS 0.007869f
C256 B.n216 VSUBS 0.007869f
C257 B.n217 VSUBS 0.005439f
C258 B.n218 VSUBS 0.007869f
C259 B.n219 VSUBS 0.007869f
C260 B.n220 VSUBS 0.007869f
C261 B.n221 VSUBS 0.007869f
C262 B.n222 VSUBS 0.007869f
C263 B.n223 VSUBS 0.007869f
C264 B.n224 VSUBS 0.007869f
C265 B.n225 VSUBS 0.007869f
C266 B.n226 VSUBS 0.007869f
C267 B.n227 VSUBS 0.007869f
C268 B.n228 VSUBS 0.007869f
C269 B.n229 VSUBS 0.007869f
C270 B.n230 VSUBS 0.007869f
C271 B.n231 VSUBS 0.007869f
C272 B.n232 VSUBS 0.007869f
C273 B.n233 VSUBS 0.007869f
C274 B.n234 VSUBS 0.007869f
C275 B.n235 VSUBS 0.007869f
C276 B.n236 VSUBS 0.007869f
C277 B.n237 VSUBS 0.007869f
C278 B.n238 VSUBS 0.007869f
C279 B.n239 VSUBS 0.007869f
C280 B.n240 VSUBS 0.007869f
C281 B.n241 VSUBS 0.007869f
C282 B.n242 VSUBS 0.007869f
C283 B.n243 VSUBS 0.007869f
C284 B.n244 VSUBS 0.007869f
C285 B.n245 VSUBS 0.007869f
C286 B.n246 VSUBS 0.007869f
C287 B.n247 VSUBS 0.007869f
C288 B.n248 VSUBS 0.007869f
C289 B.n249 VSUBS 0.007869f
C290 B.n250 VSUBS 0.007869f
C291 B.n251 VSUBS 0.007869f
C292 B.n252 VSUBS 0.007869f
C293 B.n253 VSUBS 0.007869f
C294 B.n254 VSUBS 0.007869f
C295 B.n255 VSUBS 0.007869f
C296 B.n256 VSUBS 0.007869f
C297 B.n257 VSUBS 0.007869f
C298 B.n258 VSUBS 0.007869f
C299 B.n259 VSUBS 0.007869f
C300 B.n260 VSUBS 0.007869f
C301 B.n261 VSUBS 0.007869f
C302 B.n262 VSUBS 0.007869f
C303 B.n263 VSUBS 0.007869f
C304 B.n264 VSUBS 0.007869f
C305 B.n265 VSUBS 0.007869f
C306 B.n266 VSUBS 0.007869f
C307 B.n267 VSUBS 0.01774f
C308 B.n268 VSUBS 0.018689f
C309 B.n269 VSUBS 0.017648f
C310 B.n270 VSUBS 0.007869f
C311 B.n271 VSUBS 0.007869f
C312 B.n272 VSUBS 0.007869f
C313 B.n273 VSUBS 0.007869f
C314 B.n274 VSUBS 0.007869f
C315 B.n275 VSUBS 0.007869f
C316 B.n276 VSUBS 0.007869f
C317 B.n277 VSUBS 0.007869f
C318 B.n278 VSUBS 0.007869f
C319 B.n279 VSUBS 0.007869f
C320 B.n280 VSUBS 0.007869f
C321 B.n281 VSUBS 0.007869f
C322 B.n282 VSUBS 0.007869f
C323 B.n283 VSUBS 0.007869f
C324 B.n284 VSUBS 0.007869f
C325 B.n285 VSUBS 0.007869f
C326 B.n286 VSUBS 0.007869f
C327 B.n287 VSUBS 0.007869f
C328 B.n288 VSUBS 0.007869f
C329 B.n289 VSUBS 0.007869f
C330 B.n290 VSUBS 0.007869f
C331 B.n291 VSUBS 0.007869f
C332 B.n292 VSUBS 0.007869f
C333 B.n293 VSUBS 0.007869f
C334 B.n294 VSUBS 0.007869f
C335 B.n295 VSUBS 0.007869f
C336 B.n296 VSUBS 0.007869f
C337 B.n297 VSUBS 0.007869f
C338 B.n298 VSUBS 0.007869f
C339 B.n299 VSUBS 0.007869f
C340 B.n300 VSUBS 0.007869f
C341 B.n301 VSUBS 0.007869f
C342 B.n302 VSUBS 0.007869f
C343 B.n303 VSUBS 0.007869f
C344 B.n304 VSUBS 0.007869f
C345 B.n305 VSUBS 0.007869f
C346 B.n306 VSUBS 0.007869f
C347 B.n307 VSUBS 0.007869f
C348 B.n308 VSUBS 0.007869f
C349 B.n309 VSUBS 0.007869f
C350 B.n310 VSUBS 0.007869f
C351 B.n311 VSUBS 0.007869f
C352 B.n312 VSUBS 0.007869f
C353 B.n313 VSUBS 0.007869f
C354 B.n314 VSUBS 0.007869f
C355 B.n315 VSUBS 0.007869f
C356 B.n316 VSUBS 0.007869f
C357 B.n317 VSUBS 0.007869f
C358 B.n318 VSUBS 0.007869f
C359 B.n319 VSUBS 0.007869f
C360 B.n320 VSUBS 0.007869f
C361 B.n321 VSUBS 0.017648f
C362 B.n322 VSUBS 0.017648f
C363 B.n323 VSUBS 0.018689f
C364 B.n324 VSUBS 0.007869f
C365 B.n325 VSUBS 0.007869f
C366 B.n326 VSUBS 0.007869f
C367 B.n327 VSUBS 0.007869f
C368 B.n328 VSUBS 0.007869f
C369 B.n329 VSUBS 0.007869f
C370 B.n330 VSUBS 0.007869f
C371 B.n331 VSUBS 0.007869f
C372 B.n332 VSUBS 0.007869f
C373 B.n333 VSUBS 0.007869f
C374 B.n334 VSUBS 0.007869f
C375 B.n335 VSUBS 0.007869f
C376 B.n336 VSUBS 0.007869f
C377 B.n337 VSUBS 0.007869f
C378 B.n338 VSUBS 0.007869f
C379 B.n339 VSUBS 0.007869f
C380 B.n340 VSUBS 0.007869f
C381 B.n341 VSUBS 0.007869f
C382 B.n342 VSUBS 0.007869f
C383 B.n343 VSUBS 0.007869f
C384 B.n344 VSUBS 0.007869f
C385 B.n345 VSUBS 0.007869f
C386 B.n346 VSUBS 0.007869f
C387 B.n347 VSUBS 0.007869f
C388 B.n348 VSUBS 0.007869f
C389 B.n349 VSUBS 0.007869f
C390 B.n350 VSUBS 0.007869f
C391 B.n351 VSUBS 0.007869f
C392 B.n352 VSUBS 0.007869f
C393 B.n353 VSUBS 0.007869f
C394 B.n354 VSUBS 0.007869f
C395 B.n355 VSUBS 0.007869f
C396 B.n356 VSUBS 0.007869f
C397 B.n357 VSUBS 0.007869f
C398 B.n358 VSUBS 0.007869f
C399 B.n359 VSUBS 0.007869f
C400 B.n360 VSUBS 0.007869f
C401 B.n361 VSUBS 0.007869f
C402 B.n362 VSUBS 0.007869f
C403 B.n363 VSUBS 0.007869f
C404 B.n364 VSUBS 0.007869f
C405 B.n365 VSUBS 0.007869f
C406 B.n366 VSUBS 0.007869f
C407 B.n367 VSUBS 0.007869f
C408 B.n368 VSUBS 0.007869f
C409 B.n369 VSUBS 0.007869f
C410 B.n370 VSUBS 0.007869f
C411 B.n371 VSUBS 0.007869f
C412 B.n372 VSUBS 0.007869f
C413 B.n373 VSUBS 0.007869f
C414 B.n374 VSUBS 0.005439f
C415 B.n375 VSUBS 0.018232f
C416 B.n376 VSUBS 0.006365f
C417 B.n377 VSUBS 0.007869f
C418 B.n378 VSUBS 0.007869f
C419 B.n379 VSUBS 0.007869f
C420 B.n380 VSUBS 0.007869f
C421 B.n381 VSUBS 0.007869f
C422 B.n382 VSUBS 0.007869f
C423 B.n383 VSUBS 0.007869f
C424 B.n384 VSUBS 0.007869f
C425 B.n385 VSUBS 0.007869f
C426 B.n386 VSUBS 0.007869f
C427 B.n387 VSUBS 0.007869f
C428 B.n388 VSUBS 0.006365f
C429 B.n389 VSUBS 0.007869f
C430 B.n390 VSUBS 0.007869f
C431 B.n391 VSUBS 0.005439f
C432 B.n392 VSUBS 0.007869f
C433 B.n393 VSUBS 0.007869f
C434 B.n394 VSUBS 0.007869f
C435 B.n395 VSUBS 0.007869f
C436 B.n396 VSUBS 0.007869f
C437 B.n397 VSUBS 0.007869f
C438 B.n398 VSUBS 0.007869f
C439 B.n399 VSUBS 0.007869f
C440 B.n400 VSUBS 0.007869f
C441 B.n401 VSUBS 0.007869f
C442 B.n402 VSUBS 0.007869f
C443 B.n403 VSUBS 0.007869f
C444 B.n404 VSUBS 0.007869f
C445 B.n405 VSUBS 0.007869f
C446 B.n406 VSUBS 0.007869f
C447 B.n407 VSUBS 0.007869f
C448 B.n408 VSUBS 0.007869f
C449 B.n409 VSUBS 0.007869f
C450 B.n410 VSUBS 0.007869f
C451 B.n411 VSUBS 0.007869f
C452 B.n412 VSUBS 0.007869f
C453 B.n413 VSUBS 0.007869f
C454 B.n414 VSUBS 0.007869f
C455 B.n415 VSUBS 0.007869f
C456 B.n416 VSUBS 0.007869f
C457 B.n417 VSUBS 0.007869f
C458 B.n418 VSUBS 0.007869f
C459 B.n419 VSUBS 0.007869f
C460 B.n420 VSUBS 0.007869f
C461 B.n421 VSUBS 0.007869f
C462 B.n422 VSUBS 0.007869f
C463 B.n423 VSUBS 0.007869f
C464 B.n424 VSUBS 0.007869f
C465 B.n425 VSUBS 0.007869f
C466 B.n426 VSUBS 0.007869f
C467 B.n427 VSUBS 0.007869f
C468 B.n428 VSUBS 0.007869f
C469 B.n429 VSUBS 0.007869f
C470 B.n430 VSUBS 0.007869f
C471 B.n431 VSUBS 0.007869f
C472 B.n432 VSUBS 0.007869f
C473 B.n433 VSUBS 0.007869f
C474 B.n434 VSUBS 0.007869f
C475 B.n435 VSUBS 0.007869f
C476 B.n436 VSUBS 0.007869f
C477 B.n437 VSUBS 0.007869f
C478 B.n438 VSUBS 0.007869f
C479 B.n439 VSUBS 0.007869f
C480 B.n440 VSUBS 0.007869f
C481 B.n441 VSUBS 0.018689f
C482 B.n442 VSUBS 0.018689f
C483 B.n443 VSUBS 0.017648f
C484 B.n444 VSUBS 0.007869f
C485 B.n445 VSUBS 0.007869f
C486 B.n446 VSUBS 0.007869f
C487 B.n447 VSUBS 0.007869f
C488 B.n448 VSUBS 0.007869f
C489 B.n449 VSUBS 0.007869f
C490 B.n450 VSUBS 0.007869f
C491 B.n451 VSUBS 0.007869f
C492 B.n452 VSUBS 0.007869f
C493 B.n453 VSUBS 0.007869f
C494 B.n454 VSUBS 0.007869f
C495 B.n455 VSUBS 0.007869f
C496 B.n456 VSUBS 0.007869f
C497 B.n457 VSUBS 0.007869f
C498 B.n458 VSUBS 0.007869f
C499 B.n459 VSUBS 0.007869f
C500 B.n460 VSUBS 0.007869f
C501 B.n461 VSUBS 0.007869f
C502 B.n462 VSUBS 0.007869f
C503 B.n463 VSUBS 0.007869f
C504 B.n464 VSUBS 0.007869f
C505 B.n465 VSUBS 0.007869f
C506 B.n466 VSUBS 0.007869f
C507 B.n467 VSUBS 0.010269f
C508 B.n468 VSUBS 0.010939f
C509 B.n469 VSUBS 0.021753f
C510 VDD1.t0 VSUBS 1.88677f
C511 VDD1.t1 VSUBS 1.88593f
C512 VDD1.t4 VSUBS 0.191145f
C513 VDD1.t2 VSUBS 0.191145f
C514 VDD1.n0 VSUBS 1.43504f
C515 VDD1.n1 VSUBS 2.41036f
C516 VDD1.t5 VSUBS 0.191145f
C517 VDD1.t3 VSUBS 0.191145f
C518 VDD1.n2 VSUBS 1.43425f
C519 VDD1.n3 VSUBS 2.25334f
C520 VP.n0 VSUBS 0.067481f
C521 VP.t4 VSUBS 0.880665f
C522 VP.t5 VSUBS 0.891126f
C523 VP.n1 VSUBS 0.355781f
C524 VP.t0 VSUBS 0.874908f
C525 VP.n2 VSUBS 0.377093f
C526 VP.t2 VSUBS 0.880665f
C527 VP.n3 VSUBS 0.36572f
C528 VP.n4 VSUBS 2.57333f
C529 VP.n5 VSUBS 2.47793f
C530 VP.n6 VSUBS 0.36572f
C531 VP.t1 VSUBS 0.874908f
C532 VP.n7 VSUBS 0.377093f
C533 VP.t3 VSUBS 0.880665f
C534 VP.n8 VSUBS 0.36572f
C535 VP.n9 VSUBS 0.052295f
C536 VDD2.t0 VSUBS 1.88485f
C537 VDD2.t3 VSUBS 0.191036f
C538 VDD2.t4 VSUBS 0.191036f
C539 VDD2.n0 VSUBS 1.43422f
C540 VDD2.n1 VSUBS 2.33752f
C541 VDD2.t5 VSUBS 1.88166f
C542 VDD2.n2 VSUBS 2.28509f
C543 VDD2.t1 VSUBS 0.191036f
C544 VDD2.t2 VSUBS 0.191036f
C545 VDD2.n3 VSUBS 1.43419f
C546 VTAIL.t10 VSUBS 0.238318f
C547 VTAIL.t8 VSUBS 0.238318f
C548 VTAIL.n0 VSUBS 1.63874f
C549 VTAIL.n1 VSUBS 0.771491f
C550 VTAIL.t2 VSUBS 2.18238f
C551 VTAIL.n2 VSUBS 0.924131f
C552 VTAIL.t1 VSUBS 0.238318f
C553 VTAIL.t0 VSUBS 0.238318f
C554 VTAIL.n3 VSUBS 1.63874f
C555 VTAIL.n4 VSUBS 2.13792f
C556 VTAIL.t7 VSUBS 0.238318f
C557 VTAIL.t5 VSUBS 0.238318f
C558 VTAIL.n5 VSUBS 1.63874f
C559 VTAIL.n6 VSUBS 2.13791f
C560 VTAIL.t9 VSUBS 2.18239f
C561 VTAIL.n7 VSUBS 0.924116f
C562 VTAIL.t3 VSUBS 0.238318f
C563 VTAIL.t4 VSUBS 0.238318f
C564 VTAIL.n8 VSUBS 1.63874f
C565 VTAIL.n9 VSUBS 0.817807f
C566 VTAIL.t11 VSUBS 2.18238f
C567 VTAIL.n10 VSUBS 2.17464f
C568 VTAIL.t6 VSUBS 2.18238f
C569 VTAIL.n11 VSUBS 2.15137f
C570 VN.t5 VSUBS 0.863625f
C571 VN.n0 VSUBS 0.344801f
C572 VN.t2 VSUBS 0.847908f
C573 VN.n1 VSUBS 0.365456f
C574 VN.t1 VSUBS 0.853487f
C575 VN.n2 VSUBS 0.354433f
C576 VN.n3 VSUBS 0.203955f
C577 VN.t3 VSUBS 0.863625f
C578 VN.n4 VSUBS 0.344801f
C579 VN.t0 VSUBS 0.853487f
C580 VN.t4 VSUBS 0.847908f
C581 VN.n5 VSUBS 0.365456f
C582 VN.n6 VSUBS 0.354433f
C583 VN.n7 VSUBS 2.53708f
.ends

