* NGSPICE file created from diff_pair_sample_1488.ext - technology: sky130A

.subckt diff_pair_sample_1488 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=0 ps=0 w=13.74 l=1.91
X1 VDD2.t7 VN.t0 VTAIL.t7 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X2 VDD1.t7 VP.t0 VTAIL.t4 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X3 VDD2.t6 VN.t1 VTAIL.t10 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X4 VTAIL.t8 VN.t2 VDD2.t5 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=2.2671 ps=14.07 w=13.74 l=1.91
X5 VTAIL.t9 VN.t3 VDD2.t4 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=2.2671 ps=14.07 w=13.74 l=1.91
X6 VDD1.t6 VP.t1 VTAIL.t0 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=5.3586 ps=28.26 w=13.74 l=1.91
X7 VTAIL.t6 VP.t2 VDD1.t5 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X8 B.t8 B.t6 B.t7 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=0 ps=0 w=13.74 l=1.91
X9 VDD2.t3 VN.t4 VTAIL.t11 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=5.3586 ps=28.26 w=13.74 l=1.91
X10 VTAIL.t3 VP.t3 VDD1.t4 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X11 VTAIL.t14 VN.t5 VDD2.t2 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X12 VDD1.t3 VP.t4 VTAIL.t5 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=5.3586 ps=28.26 w=13.74 l=1.91
X13 VTAIL.t13 VN.t6 VDD2.t1 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X14 VDD2.t0 VN.t7 VTAIL.t12 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=5.3586 ps=28.26 w=13.74 l=1.91
X15 VDD1.t2 VP.t5 VTAIL.t2 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=2.2671 pd=14.07 as=2.2671 ps=14.07 w=13.74 l=1.91
X16 VTAIL.t15 VP.t6 VDD1.t1 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=2.2671 ps=14.07 w=13.74 l=1.91
X17 B.t5 B.t3 B.t4 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=0 ps=0 w=13.74 l=1.91
X18 VTAIL.t1 VP.t7 VDD1.t0 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=2.2671 ps=14.07 w=13.74 l=1.91
X19 B.t2 B.t0 B.t1 w_n3210_n3716# sky130_fd_pr__pfet_01v8 ad=5.3586 pd=28.26 as=0 ps=0 w=13.74 l=1.91
R0 B.n537 B.n78 585
R1 B.n539 B.n538 585
R2 B.n540 B.n77 585
R3 B.n542 B.n541 585
R4 B.n543 B.n76 585
R5 B.n545 B.n544 585
R6 B.n546 B.n75 585
R7 B.n548 B.n547 585
R8 B.n549 B.n74 585
R9 B.n551 B.n550 585
R10 B.n552 B.n73 585
R11 B.n554 B.n553 585
R12 B.n555 B.n72 585
R13 B.n557 B.n556 585
R14 B.n558 B.n71 585
R15 B.n560 B.n559 585
R16 B.n561 B.n70 585
R17 B.n563 B.n562 585
R18 B.n564 B.n69 585
R19 B.n566 B.n565 585
R20 B.n567 B.n68 585
R21 B.n569 B.n568 585
R22 B.n570 B.n67 585
R23 B.n572 B.n571 585
R24 B.n573 B.n66 585
R25 B.n575 B.n574 585
R26 B.n576 B.n65 585
R27 B.n578 B.n577 585
R28 B.n579 B.n64 585
R29 B.n581 B.n580 585
R30 B.n582 B.n63 585
R31 B.n584 B.n583 585
R32 B.n585 B.n62 585
R33 B.n587 B.n586 585
R34 B.n588 B.n61 585
R35 B.n590 B.n589 585
R36 B.n591 B.n60 585
R37 B.n593 B.n592 585
R38 B.n594 B.n59 585
R39 B.n596 B.n595 585
R40 B.n597 B.n58 585
R41 B.n599 B.n598 585
R42 B.n600 B.n57 585
R43 B.n602 B.n601 585
R44 B.n603 B.n56 585
R45 B.n605 B.n604 585
R46 B.n606 B.n53 585
R47 B.n609 B.n608 585
R48 B.n610 B.n52 585
R49 B.n612 B.n611 585
R50 B.n613 B.n51 585
R51 B.n615 B.n614 585
R52 B.n616 B.n50 585
R53 B.n618 B.n617 585
R54 B.n619 B.n49 585
R55 B.n621 B.n620 585
R56 B.n623 B.n622 585
R57 B.n624 B.n45 585
R58 B.n626 B.n625 585
R59 B.n627 B.n44 585
R60 B.n629 B.n628 585
R61 B.n630 B.n43 585
R62 B.n632 B.n631 585
R63 B.n633 B.n42 585
R64 B.n635 B.n634 585
R65 B.n636 B.n41 585
R66 B.n638 B.n637 585
R67 B.n639 B.n40 585
R68 B.n641 B.n640 585
R69 B.n642 B.n39 585
R70 B.n644 B.n643 585
R71 B.n645 B.n38 585
R72 B.n647 B.n646 585
R73 B.n648 B.n37 585
R74 B.n650 B.n649 585
R75 B.n651 B.n36 585
R76 B.n653 B.n652 585
R77 B.n654 B.n35 585
R78 B.n656 B.n655 585
R79 B.n657 B.n34 585
R80 B.n659 B.n658 585
R81 B.n660 B.n33 585
R82 B.n662 B.n661 585
R83 B.n663 B.n32 585
R84 B.n665 B.n664 585
R85 B.n666 B.n31 585
R86 B.n668 B.n667 585
R87 B.n669 B.n30 585
R88 B.n671 B.n670 585
R89 B.n672 B.n29 585
R90 B.n674 B.n673 585
R91 B.n675 B.n28 585
R92 B.n677 B.n676 585
R93 B.n678 B.n27 585
R94 B.n680 B.n679 585
R95 B.n681 B.n26 585
R96 B.n683 B.n682 585
R97 B.n684 B.n25 585
R98 B.n686 B.n685 585
R99 B.n687 B.n24 585
R100 B.n689 B.n688 585
R101 B.n690 B.n23 585
R102 B.n692 B.n691 585
R103 B.n536 B.n535 585
R104 B.n534 B.n79 585
R105 B.n533 B.n532 585
R106 B.n531 B.n80 585
R107 B.n530 B.n529 585
R108 B.n528 B.n81 585
R109 B.n527 B.n526 585
R110 B.n525 B.n82 585
R111 B.n524 B.n523 585
R112 B.n522 B.n83 585
R113 B.n521 B.n520 585
R114 B.n519 B.n84 585
R115 B.n518 B.n517 585
R116 B.n516 B.n85 585
R117 B.n515 B.n514 585
R118 B.n513 B.n86 585
R119 B.n512 B.n511 585
R120 B.n510 B.n87 585
R121 B.n509 B.n508 585
R122 B.n507 B.n88 585
R123 B.n506 B.n505 585
R124 B.n504 B.n89 585
R125 B.n503 B.n502 585
R126 B.n501 B.n90 585
R127 B.n500 B.n499 585
R128 B.n498 B.n91 585
R129 B.n497 B.n496 585
R130 B.n495 B.n92 585
R131 B.n494 B.n493 585
R132 B.n492 B.n93 585
R133 B.n491 B.n490 585
R134 B.n489 B.n94 585
R135 B.n488 B.n487 585
R136 B.n486 B.n95 585
R137 B.n485 B.n484 585
R138 B.n483 B.n96 585
R139 B.n482 B.n481 585
R140 B.n480 B.n97 585
R141 B.n479 B.n478 585
R142 B.n477 B.n98 585
R143 B.n476 B.n475 585
R144 B.n474 B.n99 585
R145 B.n473 B.n472 585
R146 B.n471 B.n100 585
R147 B.n470 B.n469 585
R148 B.n468 B.n101 585
R149 B.n467 B.n466 585
R150 B.n465 B.n102 585
R151 B.n464 B.n463 585
R152 B.n462 B.n103 585
R153 B.n461 B.n460 585
R154 B.n459 B.n104 585
R155 B.n458 B.n457 585
R156 B.n456 B.n105 585
R157 B.n455 B.n454 585
R158 B.n453 B.n106 585
R159 B.n452 B.n451 585
R160 B.n450 B.n107 585
R161 B.n449 B.n448 585
R162 B.n447 B.n108 585
R163 B.n446 B.n445 585
R164 B.n444 B.n109 585
R165 B.n443 B.n442 585
R166 B.n441 B.n110 585
R167 B.n440 B.n439 585
R168 B.n438 B.n111 585
R169 B.n437 B.n436 585
R170 B.n435 B.n112 585
R171 B.n434 B.n433 585
R172 B.n432 B.n113 585
R173 B.n431 B.n430 585
R174 B.n429 B.n114 585
R175 B.n428 B.n427 585
R176 B.n426 B.n115 585
R177 B.n425 B.n424 585
R178 B.n423 B.n116 585
R179 B.n422 B.n421 585
R180 B.n420 B.n117 585
R181 B.n419 B.n418 585
R182 B.n417 B.n118 585
R183 B.n416 B.n415 585
R184 B.n414 B.n119 585
R185 B.n413 B.n412 585
R186 B.n257 B.n256 585
R187 B.n258 B.n175 585
R188 B.n260 B.n259 585
R189 B.n261 B.n174 585
R190 B.n263 B.n262 585
R191 B.n264 B.n173 585
R192 B.n266 B.n265 585
R193 B.n267 B.n172 585
R194 B.n269 B.n268 585
R195 B.n270 B.n171 585
R196 B.n272 B.n271 585
R197 B.n273 B.n170 585
R198 B.n275 B.n274 585
R199 B.n276 B.n169 585
R200 B.n278 B.n277 585
R201 B.n279 B.n168 585
R202 B.n281 B.n280 585
R203 B.n282 B.n167 585
R204 B.n284 B.n283 585
R205 B.n285 B.n166 585
R206 B.n287 B.n286 585
R207 B.n288 B.n165 585
R208 B.n290 B.n289 585
R209 B.n291 B.n164 585
R210 B.n293 B.n292 585
R211 B.n294 B.n163 585
R212 B.n296 B.n295 585
R213 B.n297 B.n162 585
R214 B.n299 B.n298 585
R215 B.n300 B.n161 585
R216 B.n302 B.n301 585
R217 B.n303 B.n160 585
R218 B.n305 B.n304 585
R219 B.n306 B.n159 585
R220 B.n308 B.n307 585
R221 B.n309 B.n158 585
R222 B.n311 B.n310 585
R223 B.n312 B.n157 585
R224 B.n314 B.n313 585
R225 B.n315 B.n156 585
R226 B.n317 B.n316 585
R227 B.n318 B.n155 585
R228 B.n320 B.n319 585
R229 B.n321 B.n154 585
R230 B.n323 B.n322 585
R231 B.n324 B.n153 585
R232 B.n326 B.n325 585
R233 B.n328 B.n327 585
R234 B.n329 B.n149 585
R235 B.n331 B.n330 585
R236 B.n332 B.n148 585
R237 B.n334 B.n333 585
R238 B.n335 B.n147 585
R239 B.n337 B.n336 585
R240 B.n338 B.n146 585
R241 B.n340 B.n339 585
R242 B.n342 B.n143 585
R243 B.n344 B.n343 585
R244 B.n345 B.n142 585
R245 B.n347 B.n346 585
R246 B.n348 B.n141 585
R247 B.n350 B.n349 585
R248 B.n351 B.n140 585
R249 B.n353 B.n352 585
R250 B.n354 B.n139 585
R251 B.n356 B.n355 585
R252 B.n357 B.n138 585
R253 B.n359 B.n358 585
R254 B.n360 B.n137 585
R255 B.n362 B.n361 585
R256 B.n363 B.n136 585
R257 B.n365 B.n364 585
R258 B.n366 B.n135 585
R259 B.n368 B.n367 585
R260 B.n369 B.n134 585
R261 B.n371 B.n370 585
R262 B.n372 B.n133 585
R263 B.n374 B.n373 585
R264 B.n375 B.n132 585
R265 B.n377 B.n376 585
R266 B.n378 B.n131 585
R267 B.n380 B.n379 585
R268 B.n381 B.n130 585
R269 B.n383 B.n382 585
R270 B.n384 B.n129 585
R271 B.n386 B.n385 585
R272 B.n387 B.n128 585
R273 B.n389 B.n388 585
R274 B.n390 B.n127 585
R275 B.n392 B.n391 585
R276 B.n393 B.n126 585
R277 B.n395 B.n394 585
R278 B.n396 B.n125 585
R279 B.n398 B.n397 585
R280 B.n399 B.n124 585
R281 B.n401 B.n400 585
R282 B.n402 B.n123 585
R283 B.n404 B.n403 585
R284 B.n405 B.n122 585
R285 B.n407 B.n406 585
R286 B.n408 B.n121 585
R287 B.n410 B.n409 585
R288 B.n411 B.n120 585
R289 B.n255 B.n176 585
R290 B.n254 B.n253 585
R291 B.n252 B.n177 585
R292 B.n251 B.n250 585
R293 B.n249 B.n178 585
R294 B.n248 B.n247 585
R295 B.n246 B.n179 585
R296 B.n245 B.n244 585
R297 B.n243 B.n180 585
R298 B.n242 B.n241 585
R299 B.n240 B.n181 585
R300 B.n239 B.n238 585
R301 B.n237 B.n182 585
R302 B.n236 B.n235 585
R303 B.n234 B.n183 585
R304 B.n233 B.n232 585
R305 B.n231 B.n184 585
R306 B.n230 B.n229 585
R307 B.n228 B.n185 585
R308 B.n227 B.n226 585
R309 B.n225 B.n186 585
R310 B.n224 B.n223 585
R311 B.n222 B.n187 585
R312 B.n221 B.n220 585
R313 B.n219 B.n188 585
R314 B.n218 B.n217 585
R315 B.n216 B.n189 585
R316 B.n215 B.n214 585
R317 B.n213 B.n190 585
R318 B.n212 B.n211 585
R319 B.n210 B.n191 585
R320 B.n209 B.n208 585
R321 B.n207 B.n192 585
R322 B.n206 B.n205 585
R323 B.n204 B.n193 585
R324 B.n203 B.n202 585
R325 B.n201 B.n194 585
R326 B.n200 B.n199 585
R327 B.n198 B.n195 585
R328 B.n197 B.n196 585
R329 B.n2 B.n0 585
R330 B.n753 B.n1 585
R331 B.n752 B.n751 585
R332 B.n750 B.n3 585
R333 B.n749 B.n748 585
R334 B.n747 B.n4 585
R335 B.n746 B.n745 585
R336 B.n744 B.n5 585
R337 B.n743 B.n742 585
R338 B.n741 B.n6 585
R339 B.n740 B.n739 585
R340 B.n738 B.n7 585
R341 B.n737 B.n736 585
R342 B.n735 B.n8 585
R343 B.n734 B.n733 585
R344 B.n732 B.n9 585
R345 B.n731 B.n730 585
R346 B.n729 B.n10 585
R347 B.n728 B.n727 585
R348 B.n726 B.n11 585
R349 B.n725 B.n724 585
R350 B.n723 B.n12 585
R351 B.n722 B.n721 585
R352 B.n720 B.n13 585
R353 B.n719 B.n718 585
R354 B.n717 B.n14 585
R355 B.n716 B.n715 585
R356 B.n714 B.n15 585
R357 B.n713 B.n712 585
R358 B.n711 B.n16 585
R359 B.n710 B.n709 585
R360 B.n708 B.n17 585
R361 B.n707 B.n706 585
R362 B.n705 B.n18 585
R363 B.n704 B.n703 585
R364 B.n702 B.n19 585
R365 B.n701 B.n700 585
R366 B.n699 B.n20 585
R367 B.n698 B.n697 585
R368 B.n696 B.n21 585
R369 B.n695 B.n694 585
R370 B.n693 B.n22 585
R371 B.n755 B.n754 585
R372 B.n256 B.n255 511.721
R373 B.n693 B.n692 511.721
R374 B.n412 B.n411 511.721
R375 B.n537 B.n536 511.721
R376 B.n144 B.t0 380.067
R377 B.n150 B.t9 380.067
R378 B.n46 B.t6 380.067
R379 B.n54 B.t3 380.067
R380 B.n255 B.n254 163.367
R381 B.n254 B.n177 163.367
R382 B.n250 B.n177 163.367
R383 B.n250 B.n249 163.367
R384 B.n249 B.n248 163.367
R385 B.n248 B.n179 163.367
R386 B.n244 B.n179 163.367
R387 B.n244 B.n243 163.367
R388 B.n243 B.n242 163.367
R389 B.n242 B.n181 163.367
R390 B.n238 B.n181 163.367
R391 B.n238 B.n237 163.367
R392 B.n237 B.n236 163.367
R393 B.n236 B.n183 163.367
R394 B.n232 B.n183 163.367
R395 B.n232 B.n231 163.367
R396 B.n231 B.n230 163.367
R397 B.n230 B.n185 163.367
R398 B.n226 B.n185 163.367
R399 B.n226 B.n225 163.367
R400 B.n225 B.n224 163.367
R401 B.n224 B.n187 163.367
R402 B.n220 B.n187 163.367
R403 B.n220 B.n219 163.367
R404 B.n219 B.n218 163.367
R405 B.n218 B.n189 163.367
R406 B.n214 B.n189 163.367
R407 B.n214 B.n213 163.367
R408 B.n213 B.n212 163.367
R409 B.n212 B.n191 163.367
R410 B.n208 B.n191 163.367
R411 B.n208 B.n207 163.367
R412 B.n207 B.n206 163.367
R413 B.n206 B.n193 163.367
R414 B.n202 B.n193 163.367
R415 B.n202 B.n201 163.367
R416 B.n201 B.n200 163.367
R417 B.n200 B.n195 163.367
R418 B.n196 B.n195 163.367
R419 B.n196 B.n2 163.367
R420 B.n754 B.n2 163.367
R421 B.n754 B.n753 163.367
R422 B.n753 B.n752 163.367
R423 B.n752 B.n3 163.367
R424 B.n748 B.n3 163.367
R425 B.n748 B.n747 163.367
R426 B.n747 B.n746 163.367
R427 B.n746 B.n5 163.367
R428 B.n742 B.n5 163.367
R429 B.n742 B.n741 163.367
R430 B.n741 B.n740 163.367
R431 B.n740 B.n7 163.367
R432 B.n736 B.n7 163.367
R433 B.n736 B.n735 163.367
R434 B.n735 B.n734 163.367
R435 B.n734 B.n9 163.367
R436 B.n730 B.n9 163.367
R437 B.n730 B.n729 163.367
R438 B.n729 B.n728 163.367
R439 B.n728 B.n11 163.367
R440 B.n724 B.n11 163.367
R441 B.n724 B.n723 163.367
R442 B.n723 B.n722 163.367
R443 B.n722 B.n13 163.367
R444 B.n718 B.n13 163.367
R445 B.n718 B.n717 163.367
R446 B.n717 B.n716 163.367
R447 B.n716 B.n15 163.367
R448 B.n712 B.n15 163.367
R449 B.n712 B.n711 163.367
R450 B.n711 B.n710 163.367
R451 B.n710 B.n17 163.367
R452 B.n706 B.n17 163.367
R453 B.n706 B.n705 163.367
R454 B.n705 B.n704 163.367
R455 B.n704 B.n19 163.367
R456 B.n700 B.n19 163.367
R457 B.n700 B.n699 163.367
R458 B.n699 B.n698 163.367
R459 B.n698 B.n21 163.367
R460 B.n694 B.n21 163.367
R461 B.n694 B.n693 163.367
R462 B.n256 B.n175 163.367
R463 B.n260 B.n175 163.367
R464 B.n261 B.n260 163.367
R465 B.n262 B.n261 163.367
R466 B.n262 B.n173 163.367
R467 B.n266 B.n173 163.367
R468 B.n267 B.n266 163.367
R469 B.n268 B.n267 163.367
R470 B.n268 B.n171 163.367
R471 B.n272 B.n171 163.367
R472 B.n273 B.n272 163.367
R473 B.n274 B.n273 163.367
R474 B.n274 B.n169 163.367
R475 B.n278 B.n169 163.367
R476 B.n279 B.n278 163.367
R477 B.n280 B.n279 163.367
R478 B.n280 B.n167 163.367
R479 B.n284 B.n167 163.367
R480 B.n285 B.n284 163.367
R481 B.n286 B.n285 163.367
R482 B.n286 B.n165 163.367
R483 B.n290 B.n165 163.367
R484 B.n291 B.n290 163.367
R485 B.n292 B.n291 163.367
R486 B.n292 B.n163 163.367
R487 B.n296 B.n163 163.367
R488 B.n297 B.n296 163.367
R489 B.n298 B.n297 163.367
R490 B.n298 B.n161 163.367
R491 B.n302 B.n161 163.367
R492 B.n303 B.n302 163.367
R493 B.n304 B.n303 163.367
R494 B.n304 B.n159 163.367
R495 B.n308 B.n159 163.367
R496 B.n309 B.n308 163.367
R497 B.n310 B.n309 163.367
R498 B.n310 B.n157 163.367
R499 B.n314 B.n157 163.367
R500 B.n315 B.n314 163.367
R501 B.n316 B.n315 163.367
R502 B.n316 B.n155 163.367
R503 B.n320 B.n155 163.367
R504 B.n321 B.n320 163.367
R505 B.n322 B.n321 163.367
R506 B.n322 B.n153 163.367
R507 B.n326 B.n153 163.367
R508 B.n327 B.n326 163.367
R509 B.n327 B.n149 163.367
R510 B.n331 B.n149 163.367
R511 B.n332 B.n331 163.367
R512 B.n333 B.n332 163.367
R513 B.n333 B.n147 163.367
R514 B.n337 B.n147 163.367
R515 B.n338 B.n337 163.367
R516 B.n339 B.n338 163.367
R517 B.n339 B.n143 163.367
R518 B.n344 B.n143 163.367
R519 B.n345 B.n344 163.367
R520 B.n346 B.n345 163.367
R521 B.n346 B.n141 163.367
R522 B.n350 B.n141 163.367
R523 B.n351 B.n350 163.367
R524 B.n352 B.n351 163.367
R525 B.n352 B.n139 163.367
R526 B.n356 B.n139 163.367
R527 B.n357 B.n356 163.367
R528 B.n358 B.n357 163.367
R529 B.n358 B.n137 163.367
R530 B.n362 B.n137 163.367
R531 B.n363 B.n362 163.367
R532 B.n364 B.n363 163.367
R533 B.n364 B.n135 163.367
R534 B.n368 B.n135 163.367
R535 B.n369 B.n368 163.367
R536 B.n370 B.n369 163.367
R537 B.n370 B.n133 163.367
R538 B.n374 B.n133 163.367
R539 B.n375 B.n374 163.367
R540 B.n376 B.n375 163.367
R541 B.n376 B.n131 163.367
R542 B.n380 B.n131 163.367
R543 B.n381 B.n380 163.367
R544 B.n382 B.n381 163.367
R545 B.n382 B.n129 163.367
R546 B.n386 B.n129 163.367
R547 B.n387 B.n386 163.367
R548 B.n388 B.n387 163.367
R549 B.n388 B.n127 163.367
R550 B.n392 B.n127 163.367
R551 B.n393 B.n392 163.367
R552 B.n394 B.n393 163.367
R553 B.n394 B.n125 163.367
R554 B.n398 B.n125 163.367
R555 B.n399 B.n398 163.367
R556 B.n400 B.n399 163.367
R557 B.n400 B.n123 163.367
R558 B.n404 B.n123 163.367
R559 B.n405 B.n404 163.367
R560 B.n406 B.n405 163.367
R561 B.n406 B.n121 163.367
R562 B.n410 B.n121 163.367
R563 B.n411 B.n410 163.367
R564 B.n412 B.n119 163.367
R565 B.n416 B.n119 163.367
R566 B.n417 B.n416 163.367
R567 B.n418 B.n417 163.367
R568 B.n418 B.n117 163.367
R569 B.n422 B.n117 163.367
R570 B.n423 B.n422 163.367
R571 B.n424 B.n423 163.367
R572 B.n424 B.n115 163.367
R573 B.n428 B.n115 163.367
R574 B.n429 B.n428 163.367
R575 B.n430 B.n429 163.367
R576 B.n430 B.n113 163.367
R577 B.n434 B.n113 163.367
R578 B.n435 B.n434 163.367
R579 B.n436 B.n435 163.367
R580 B.n436 B.n111 163.367
R581 B.n440 B.n111 163.367
R582 B.n441 B.n440 163.367
R583 B.n442 B.n441 163.367
R584 B.n442 B.n109 163.367
R585 B.n446 B.n109 163.367
R586 B.n447 B.n446 163.367
R587 B.n448 B.n447 163.367
R588 B.n448 B.n107 163.367
R589 B.n452 B.n107 163.367
R590 B.n453 B.n452 163.367
R591 B.n454 B.n453 163.367
R592 B.n454 B.n105 163.367
R593 B.n458 B.n105 163.367
R594 B.n459 B.n458 163.367
R595 B.n460 B.n459 163.367
R596 B.n460 B.n103 163.367
R597 B.n464 B.n103 163.367
R598 B.n465 B.n464 163.367
R599 B.n466 B.n465 163.367
R600 B.n466 B.n101 163.367
R601 B.n470 B.n101 163.367
R602 B.n471 B.n470 163.367
R603 B.n472 B.n471 163.367
R604 B.n472 B.n99 163.367
R605 B.n476 B.n99 163.367
R606 B.n477 B.n476 163.367
R607 B.n478 B.n477 163.367
R608 B.n478 B.n97 163.367
R609 B.n482 B.n97 163.367
R610 B.n483 B.n482 163.367
R611 B.n484 B.n483 163.367
R612 B.n484 B.n95 163.367
R613 B.n488 B.n95 163.367
R614 B.n489 B.n488 163.367
R615 B.n490 B.n489 163.367
R616 B.n490 B.n93 163.367
R617 B.n494 B.n93 163.367
R618 B.n495 B.n494 163.367
R619 B.n496 B.n495 163.367
R620 B.n496 B.n91 163.367
R621 B.n500 B.n91 163.367
R622 B.n501 B.n500 163.367
R623 B.n502 B.n501 163.367
R624 B.n502 B.n89 163.367
R625 B.n506 B.n89 163.367
R626 B.n507 B.n506 163.367
R627 B.n508 B.n507 163.367
R628 B.n508 B.n87 163.367
R629 B.n512 B.n87 163.367
R630 B.n513 B.n512 163.367
R631 B.n514 B.n513 163.367
R632 B.n514 B.n85 163.367
R633 B.n518 B.n85 163.367
R634 B.n519 B.n518 163.367
R635 B.n520 B.n519 163.367
R636 B.n520 B.n83 163.367
R637 B.n524 B.n83 163.367
R638 B.n525 B.n524 163.367
R639 B.n526 B.n525 163.367
R640 B.n526 B.n81 163.367
R641 B.n530 B.n81 163.367
R642 B.n531 B.n530 163.367
R643 B.n532 B.n531 163.367
R644 B.n532 B.n79 163.367
R645 B.n536 B.n79 163.367
R646 B.n692 B.n23 163.367
R647 B.n688 B.n23 163.367
R648 B.n688 B.n687 163.367
R649 B.n687 B.n686 163.367
R650 B.n686 B.n25 163.367
R651 B.n682 B.n25 163.367
R652 B.n682 B.n681 163.367
R653 B.n681 B.n680 163.367
R654 B.n680 B.n27 163.367
R655 B.n676 B.n27 163.367
R656 B.n676 B.n675 163.367
R657 B.n675 B.n674 163.367
R658 B.n674 B.n29 163.367
R659 B.n670 B.n29 163.367
R660 B.n670 B.n669 163.367
R661 B.n669 B.n668 163.367
R662 B.n668 B.n31 163.367
R663 B.n664 B.n31 163.367
R664 B.n664 B.n663 163.367
R665 B.n663 B.n662 163.367
R666 B.n662 B.n33 163.367
R667 B.n658 B.n33 163.367
R668 B.n658 B.n657 163.367
R669 B.n657 B.n656 163.367
R670 B.n656 B.n35 163.367
R671 B.n652 B.n35 163.367
R672 B.n652 B.n651 163.367
R673 B.n651 B.n650 163.367
R674 B.n650 B.n37 163.367
R675 B.n646 B.n37 163.367
R676 B.n646 B.n645 163.367
R677 B.n645 B.n644 163.367
R678 B.n644 B.n39 163.367
R679 B.n640 B.n39 163.367
R680 B.n640 B.n639 163.367
R681 B.n639 B.n638 163.367
R682 B.n638 B.n41 163.367
R683 B.n634 B.n41 163.367
R684 B.n634 B.n633 163.367
R685 B.n633 B.n632 163.367
R686 B.n632 B.n43 163.367
R687 B.n628 B.n43 163.367
R688 B.n628 B.n627 163.367
R689 B.n627 B.n626 163.367
R690 B.n626 B.n45 163.367
R691 B.n622 B.n45 163.367
R692 B.n622 B.n621 163.367
R693 B.n621 B.n49 163.367
R694 B.n617 B.n49 163.367
R695 B.n617 B.n616 163.367
R696 B.n616 B.n615 163.367
R697 B.n615 B.n51 163.367
R698 B.n611 B.n51 163.367
R699 B.n611 B.n610 163.367
R700 B.n610 B.n609 163.367
R701 B.n609 B.n53 163.367
R702 B.n604 B.n53 163.367
R703 B.n604 B.n603 163.367
R704 B.n603 B.n602 163.367
R705 B.n602 B.n57 163.367
R706 B.n598 B.n57 163.367
R707 B.n598 B.n597 163.367
R708 B.n597 B.n596 163.367
R709 B.n596 B.n59 163.367
R710 B.n592 B.n59 163.367
R711 B.n592 B.n591 163.367
R712 B.n591 B.n590 163.367
R713 B.n590 B.n61 163.367
R714 B.n586 B.n61 163.367
R715 B.n586 B.n585 163.367
R716 B.n585 B.n584 163.367
R717 B.n584 B.n63 163.367
R718 B.n580 B.n63 163.367
R719 B.n580 B.n579 163.367
R720 B.n579 B.n578 163.367
R721 B.n578 B.n65 163.367
R722 B.n574 B.n65 163.367
R723 B.n574 B.n573 163.367
R724 B.n573 B.n572 163.367
R725 B.n572 B.n67 163.367
R726 B.n568 B.n67 163.367
R727 B.n568 B.n567 163.367
R728 B.n567 B.n566 163.367
R729 B.n566 B.n69 163.367
R730 B.n562 B.n69 163.367
R731 B.n562 B.n561 163.367
R732 B.n561 B.n560 163.367
R733 B.n560 B.n71 163.367
R734 B.n556 B.n71 163.367
R735 B.n556 B.n555 163.367
R736 B.n555 B.n554 163.367
R737 B.n554 B.n73 163.367
R738 B.n550 B.n73 163.367
R739 B.n550 B.n549 163.367
R740 B.n549 B.n548 163.367
R741 B.n548 B.n75 163.367
R742 B.n544 B.n75 163.367
R743 B.n544 B.n543 163.367
R744 B.n543 B.n542 163.367
R745 B.n542 B.n77 163.367
R746 B.n538 B.n77 163.367
R747 B.n538 B.n537 163.367
R748 B.n144 B.t2 152.917
R749 B.n54 B.t4 152.917
R750 B.n150 B.t11 152.899
R751 B.n46 B.t7 152.899
R752 B.n145 B.t1 109.475
R753 B.n55 B.t5 109.475
R754 B.n151 B.t10 109.457
R755 B.n47 B.t8 109.457
R756 B.n341 B.n145 59.5399
R757 B.n152 B.n151 59.5399
R758 B.n48 B.n47 59.5399
R759 B.n607 B.n55 59.5399
R760 B.n145 B.n144 43.4429
R761 B.n151 B.n150 43.4429
R762 B.n47 B.n46 43.4429
R763 B.n55 B.n54 43.4429
R764 B.n691 B.n22 33.2493
R765 B.n535 B.n78 33.2493
R766 B.n413 B.n120 33.2493
R767 B.n257 B.n176 33.2493
R768 B B.n755 18.0485
R769 B.n691 B.n690 10.6151
R770 B.n690 B.n689 10.6151
R771 B.n689 B.n24 10.6151
R772 B.n685 B.n24 10.6151
R773 B.n685 B.n684 10.6151
R774 B.n684 B.n683 10.6151
R775 B.n683 B.n26 10.6151
R776 B.n679 B.n26 10.6151
R777 B.n679 B.n678 10.6151
R778 B.n678 B.n677 10.6151
R779 B.n677 B.n28 10.6151
R780 B.n673 B.n28 10.6151
R781 B.n673 B.n672 10.6151
R782 B.n672 B.n671 10.6151
R783 B.n671 B.n30 10.6151
R784 B.n667 B.n30 10.6151
R785 B.n667 B.n666 10.6151
R786 B.n666 B.n665 10.6151
R787 B.n665 B.n32 10.6151
R788 B.n661 B.n32 10.6151
R789 B.n661 B.n660 10.6151
R790 B.n660 B.n659 10.6151
R791 B.n659 B.n34 10.6151
R792 B.n655 B.n34 10.6151
R793 B.n655 B.n654 10.6151
R794 B.n654 B.n653 10.6151
R795 B.n653 B.n36 10.6151
R796 B.n649 B.n36 10.6151
R797 B.n649 B.n648 10.6151
R798 B.n648 B.n647 10.6151
R799 B.n647 B.n38 10.6151
R800 B.n643 B.n38 10.6151
R801 B.n643 B.n642 10.6151
R802 B.n642 B.n641 10.6151
R803 B.n641 B.n40 10.6151
R804 B.n637 B.n40 10.6151
R805 B.n637 B.n636 10.6151
R806 B.n636 B.n635 10.6151
R807 B.n635 B.n42 10.6151
R808 B.n631 B.n42 10.6151
R809 B.n631 B.n630 10.6151
R810 B.n630 B.n629 10.6151
R811 B.n629 B.n44 10.6151
R812 B.n625 B.n44 10.6151
R813 B.n625 B.n624 10.6151
R814 B.n624 B.n623 10.6151
R815 B.n620 B.n619 10.6151
R816 B.n619 B.n618 10.6151
R817 B.n618 B.n50 10.6151
R818 B.n614 B.n50 10.6151
R819 B.n614 B.n613 10.6151
R820 B.n613 B.n612 10.6151
R821 B.n612 B.n52 10.6151
R822 B.n608 B.n52 10.6151
R823 B.n606 B.n605 10.6151
R824 B.n605 B.n56 10.6151
R825 B.n601 B.n56 10.6151
R826 B.n601 B.n600 10.6151
R827 B.n600 B.n599 10.6151
R828 B.n599 B.n58 10.6151
R829 B.n595 B.n58 10.6151
R830 B.n595 B.n594 10.6151
R831 B.n594 B.n593 10.6151
R832 B.n593 B.n60 10.6151
R833 B.n589 B.n60 10.6151
R834 B.n589 B.n588 10.6151
R835 B.n588 B.n587 10.6151
R836 B.n587 B.n62 10.6151
R837 B.n583 B.n62 10.6151
R838 B.n583 B.n582 10.6151
R839 B.n582 B.n581 10.6151
R840 B.n581 B.n64 10.6151
R841 B.n577 B.n64 10.6151
R842 B.n577 B.n576 10.6151
R843 B.n576 B.n575 10.6151
R844 B.n575 B.n66 10.6151
R845 B.n571 B.n66 10.6151
R846 B.n571 B.n570 10.6151
R847 B.n570 B.n569 10.6151
R848 B.n569 B.n68 10.6151
R849 B.n565 B.n68 10.6151
R850 B.n565 B.n564 10.6151
R851 B.n564 B.n563 10.6151
R852 B.n563 B.n70 10.6151
R853 B.n559 B.n70 10.6151
R854 B.n559 B.n558 10.6151
R855 B.n558 B.n557 10.6151
R856 B.n557 B.n72 10.6151
R857 B.n553 B.n72 10.6151
R858 B.n553 B.n552 10.6151
R859 B.n552 B.n551 10.6151
R860 B.n551 B.n74 10.6151
R861 B.n547 B.n74 10.6151
R862 B.n547 B.n546 10.6151
R863 B.n546 B.n545 10.6151
R864 B.n545 B.n76 10.6151
R865 B.n541 B.n76 10.6151
R866 B.n541 B.n540 10.6151
R867 B.n540 B.n539 10.6151
R868 B.n539 B.n78 10.6151
R869 B.n414 B.n413 10.6151
R870 B.n415 B.n414 10.6151
R871 B.n415 B.n118 10.6151
R872 B.n419 B.n118 10.6151
R873 B.n420 B.n419 10.6151
R874 B.n421 B.n420 10.6151
R875 B.n421 B.n116 10.6151
R876 B.n425 B.n116 10.6151
R877 B.n426 B.n425 10.6151
R878 B.n427 B.n426 10.6151
R879 B.n427 B.n114 10.6151
R880 B.n431 B.n114 10.6151
R881 B.n432 B.n431 10.6151
R882 B.n433 B.n432 10.6151
R883 B.n433 B.n112 10.6151
R884 B.n437 B.n112 10.6151
R885 B.n438 B.n437 10.6151
R886 B.n439 B.n438 10.6151
R887 B.n439 B.n110 10.6151
R888 B.n443 B.n110 10.6151
R889 B.n444 B.n443 10.6151
R890 B.n445 B.n444 10.6151
R891 B.n445 B.n108 10.6151
R892 B.n449 B.n108 10.6151
R893 B.n450 B.n449 10.6151
R894 B.n451 B.n450 10.6151
R895 B.n451 B.n106 10.6151
R896 B.n455 B.n106 10.6151
R897 B.n456 B.n455 10.6151
R898 B.n457 B.n456 10.6151
R899 B.n457 B.n104 10.6151
R900 B.n461 B.n104 10.6151
R901 B.n462 B.n461 10.6151
R902 B.n463 B.n462 10.6151
R903 B.n463 B.n102 10.6151
R904 B.n467 B.n102 10.6151
R905 B.n468 B.n467 10.6151
R906 B.n469 B.n468 10.6151
R907 B.n469 B.n100 10.6151
R908 B.n473 B.n100 10.6151
R909 B.n474 B.n473 10.6151
R910 B.n475 B.n474 10.6151
R911 B.n475 B.n98 10.6151
R912 B.n479 B.n98 10.6151
R913 B.n480 B.n479 10.6151
R914 B.n481 B.n480 10.6151
R915 B.n481 B.n96 10.6151
R916 B.n485 B.n96 10.6151
R917 B.n486 B.n485 10.6151
R918 B.n487 B.n486 10.6151
R919 B.n487 B.n94 10.6151
R920 B.n491 B.n94 10.6151
R921 B.n492 B.n491 10.6151
R922 B.n493 B.n492 10.6151
R923 B.n493 B.n92 10.6151
R924 B.n497 B.n92 10.6151
R925 B.n498 B.n497 10.6151
R926 B.n499 B.n498 10.6151
R927 B.n499 B.n90 10.6151
R928 B.n503 B.n90 10.6151
R929 B.n504 B.n503 10.6151
R930 B.n505 B.n504 10.6151
R931 B.n505 B.n88 10.6151
R932 B.n509 B.n88 10.6151
R933 B.n510 B.n509 10.6151
R934 B.n511 B.n510 10.6151
R935 B.n511 B.n86 10.6151
R936 B.n515 B.n86 10.6151
R937 B.n516 B.n515 10.6151
R938 B.n517 B.n516 10.6151
R939 B.n517 B.n84 10.6151
R940 B.n521 B.n84 10.6151
R941 B.n522 B.n521 10.6151
R942 B.n523 B.n522 10.6151
R943 B.n523 B.n82 10.6151
R944 B.n527 B.n82 10.6151
R945 B.n528 B.n527 10.6151
R946 B.n529 B.n528 10.6151
R947 B.n529 B.n80 10.6151
R948 B.n533 B.n80 10.6151
R949 B.n534 B.n533 10.6151
R950 B.n535 B.n534 10.6151
R951 B.n258 B.n257 10.6151
R952 B.n259 B.n258 10.6151
R953 B.n259 B.n174 10.6151
R954 B.n263 B.n174 10.6151
R955 B.n264 B.n263 10.6151
R956 B.n265 B.n264 10.6151
R957 B.n265 B.n172 10.6151
R958 B.n269 B.n172 10.6151
R959 B.n270 B.n269 10.6151
R960 B.n271 B.n270 10.6151
R961 B.n271 B.n170 10.6151
R962 B.n275 B.n170 10.6151
R963 B.n276 B.n275 10.6151
R964 B.n277 B.n276 10.6151
R965 B.n277 B.n168 10.6151
R966 B.n281 B.n168 10.6151
R967 B.n282 B.n281 10.6151
R968 B.n283 B.n282 10.6151
R969 B.n283 B.n166 10.6151
R970 B.n287 B.n166 10.6151
R971 B.n288 B.n287 10.6151
R972 B.n289 B.n288 10.6151
R973 B.n289 B.n164 10.6151
R974 B.n293 B.n164 10.6151
R975 B.n294 B.n293 10.6151
R976 B.n295 B.n294 10.6151
R977 B.n295 B.n162 10.6151
R978 B.n299 B.n162 10.6151
R979 B.n300 B.n299 10.6151
R980 B.n301 B.n300 10.6151
R981 B.n301 B.n160 10.6151
R982 B.n305 B.n160 10.6151
R983 B.n306 B.n305 10.6151
R984 B.n307 B.n306 10.6151
R985 B.n307 B.n158 10.6151
R986 B.n311 B.n158 10.6151
R987 B.n312 B.n311 10.6151
R988 B.n313 B.n312 10.6151
R989 B.n313 B.n156 10.6151
R990 B.n317 B.n156 10.6151
R991 B.n318 B.n317 10.6151
R992 B.n319 B.n318 10.6151
R993 B.n319 B.n154 10.6151
R994 B.n323 B.n154 10.6151
R995 B.n324 B.n323 10.6151
R996 B.n325 B.n324 10.6151
R997 B.n329 B.n328 10.6151
R998 B.n330 B.n329 10.6151
R999 B.n330 B.n148 10.6151
R1000 B.n334 B.n148 10.6151
R1001 B.n335 B.n334 10.6151
R1002 B.n336 B.n335 10.6151
R1003 B.n336 B.n146 10.6151
R1004 B.n340 B.n146 10.6151
R1005 B.n343 B.n342 10.6151
R1006 B.n343 B.n142 10.6151
R1007 B.n347 B.n142 10.6151
R1008 B.n348 B.n347 10.6151
R1009 B.n349 B.n348 10.6151
R1010 B.n349 B.n140 10.6151
R1011 B.n353 B.n140 10.6151
R1012 B.n354 B.n353 10.6151
R1013 B.n355 B.n354 10.6151
R1014 B.n355 B.n138 10.6151
R1015 B.n359 B.n138 10.6151
R1016 B.n360 B.n359 10.6151
R1017 B.n361 B.n360 10.6151
R1018 B.n361 B.n136 10.6151
R1019 B.n365 B.n136 10.6151
R1020 B.n366 B.n365 10.6151
R1021 B.n367 B.n366 10.6151
R1022 B.n367 B.n134 10.6151
R1023 B.n371 B.n134 10.6151
R1024 B.n372 B.n371 10.6151
R1025 B.n373 B.n372 10.6151
R1026 B.n373 B.n132 10.6151
R1027 B.n377 B.n132 10.6151
R1028 B.n378 B.n377 10.6151
R1029 B.n379 B.n378 10.6151
R1030 B.n379 B.n130 10.6151
R1031 B.n383 B.n130 10.6151
R1032 B.n384 B.n383 10.6151
R1033 B.n385 B.n384 10.6151
R1034 B.n385 B.n128 10.6151
R1035 B.n389 B.n128 10.6151
R1036 B.n390 B.n389 10.6151
R1037 B.n391 B.n390 10.6151
R1038 B.n391 B.n126 10.6151
R1039 B.n395 B.n126 10.6151
R1040 B.n396 B.n395 10.6151
R1041 B.n397 B.n396 10.6151
R1042 B.n397 B.n124 10.6151
R1043 B.n401 B.n124 10.6151
R1044 B.n402 B.n401 10.6151
R1045 B.n403 B.n402 10.6151
R1046 B.n403 B.n122 10.6151
R1047 B.n407 B.n122 10.6151
R1048 B.n408 B.n407 10.6151
R1049 B.n409 B.n408 10.6151
R1050 B.n409 B.n120 10.6151
R1051 B.n253 B.n176 10.6151
R1052 B.n253 B.n252 10.6151
R1053 B.n252 B.n251 10.6151
R1054 B.n251 B.n178 10.6151
R1055 B.n247 B.n178 10.6151
R1056 B.n247 B.n246 10.6151
R1057 B.n246 B.n245 10.6151
R1058 B.n245 B.n180 10.6151
R1059 B.n241 B.n180 10.6151
R1060 B.n241 B.n240 10.6151
R1061 B.n240 B.n239 10.6151
R1062 B.n239 B.n182 10.6151
R1063 B.n235 B.n182 10.6151
R1064 B.n235 B.n234 10.6151
R1065 B.n234 B.n233 10.6151
R1066 B.n233 B.n184 10.6151
R1067 B.n229 B.n184 10.6151
R1068 B.n229 B.n228 10.6151
R1069 B.n228 B.n227 10.6151
R1070 B.n227 B.n186 10.6151
R1071 B.n223 B.n186 10.6151
R1072 B.n223 B.n222 10.6151
R1073 B.n222 B.n221 10.6151
R1074 B.n221 B.n188 10.6151
R1075 B.n217 B.n188 10.6151
R1076 B.n217 B.n216 10.6151
R1077 B.n216 B.n215 10.6151
R1078 B.n215 B.n190 10.6151
R1079 B.n211 B.n190 10.6151
R1080 B.n211 B.n210 10.6151
R1081 B.n210 B.n209 10.6151
R1082 B.n209 B.n192 10.6151
R1083 B.n205 B.n192 10.6151
R1084 B.n205 B.n204 10.6151
R1085 B.n204 B.n203 10.6151
R1086 B.n203 B.n194 10.6151
R1087 B.n199 B.n194 10.6151
R1088 B.n199 B.n198 10.6151
R1089 B.n198 B.n197 10.6151
R1090 B.n197 B.n0 10.6151
R1091 B.n751 B.n1 10.6151
R1092 B.n751 B.n750 10.6151
R1093 B.n750 B.n749 10.6151
R1094 B.n749 B.n4 10.6151
R1095 B.n745 B.n4 10.6151
R1096 B.n745 B.n744 10.6151
R1097 B.n744 B.n743 10.6151
R1098 B.n743 B.n6 10.6151
R1099 B.n739 B.n6 10.6151
R1100 B.n739 B.n738 10.6151
R1101 B.n738 B.n737 10.6151
R1102 B.n737 B.n8 10.6151
R1103 B.n733 B.n8 10.6151
R1104 B.n733 B.n732 10.6151
R1105 B.n732 B.n731 10.6151
R1106 B.n731 B.n10 10.6151
R1107 B.n727 B.n10 10.6151
R1108 B.n727 B.n726 10.6151
R1109 B.n726 B.n725 10.6151
R1110 B.n725 B.n12 10.6151
R1111 B.n721 B.n12 10.6151
R1112 B.n721 B.n720 10.6151
R1113 B.n720 B.n719 10.6151
R1114 B.n719 B.n14 10.6151
R1115 B.n715 B.n14 10.6151
R1116 B.n715 B.n714 10.6151
R1117 B.n714 B.n713 10.6151
R1118 B.n713 B.n16 10.6151
R1119 B.n709 B.n16 10.6151
R1120 B.n709 B.n708 10.6151
R1121 B.n708 B.n707 10.6151
R1122 B.n707 B.n18 10.6151
R1123 B.n703 B.n18 10.6151
R1124 B.n703 B.n702 10.6151
R1125 B.n702 B.n701 10.6151
R1126 B.n701 B.n20 10.6151
R1127 B.n697 B.n20 10.6151
R1128 B.n697 B.n696 10.6151
R1129 B.n696 B.n695 10.6151
R1130 B.n695 B.n22 10.6151
R1131 B.n620 B.n48 6.5566
R1132 B.n608 B.n607 6.5566
R1133 B.n328 B.n152 6.5566
R1134 B.n341 B.n340 6.5566
R1135 B.n623 B.n48 4.05904
R1136 B.n607 B.n606 4.05904
R1137 B.n325 B.n152 4.05904
R1138 B.n342 B.n341 4.05904
R1139 B.n755 B.n0 2.81026
R1140 B.n755 B.n1 2.81026
R1141 VN.n5 VN.t2 203.144
R1142 VN.n28 VN.t4 203.144
R1143 VN.n6 VN.t1 173.369
R1144 VN.n14 VN.t6 173.369
R1145 VN.n21 VN.t7 173.369
R1146 VN.n29 VN.t5 173.369
R1147 VN.n37 VN.t0 173.369
R1148 VN.n44 VN.t3 173.369
R1149 VN.n43 VN.n23 161.3
R1150 VN.n42 VN.n41 161.3
R1151 VN.n40 VN.n24 161.3
R1152 VN.n39 VN.n38 161.3
R1153 VN.n36 VN.n25 161.3
R1154 VN.n35 VN.n34 161.3
R1155 VN.n33 VN.n26 161.3
R1156 VN.n32 VN.n31 161.3
R1157 VN.n30 VN.n27 161.3
R1158 VN.n20 VN.n0 161.3
R1159 VN.n19 VN.n18 161.3
R1160 VN.n17 VN.n1 161.3
R1161 VN.n16 VN.n15 161.3
R1162 VN.n13 VN.n2 161.3
R1163 VN.n12 VN.n11 161.3
R1164 VN.n10 VN.n3 161.3
R1165 VN.n9 VN.n8 161.3
R1166 VN.n7 VN.n4 161.3
R1167 VN.n22 VN.n21 93.0789
R1168 VN.n45 VN.n44 93.0789
R1169 VN.n6 VN.n5 63.4148
R1170 VN.n29 VN.n28 63.4148
R1171 VN.n19 VN.n1 56.4773
R1172 VN.n42 VN.n24 56.4773
R1173 VN VN.n45 49.233
R1174 VN.n8 VN.n3 40.4106
R1175 VN.n12 VN.n3 40.4106
R1176 VN.n31 VN.n26 40.4106
R1177 VN.n35 VN.n26 40.4106
R1178 VN.n8 VN.n7 24.3439
R1179 VN.n13 VN.n12 24.3439
R1180 VN.n15 VN.n1 24.3439
R1181 VN.n20 VN.n19 24.3439
R1182 VN.n31 VN.n30 24.3439
R1183 VN.n38 VN.n24 24.3439
R1184 VN.n36 VN.n35 24.3439
R1185 VN.n43 VN.n42 24.3439
R1186 VN.n15 VN.n14 18.5015
R1187 VN.n38 VN.n37 18.5015
R1188 VN.n21 VN.n20 17.5278
R1189 VN.n44 VN.n43 17.5278
R1190 VN.n28 VN.n27 13.6639
R1191 VN.n5 VN.n4 13.6639
R1192 VN.n7 VN.n6 5.84292
R1193 VN.n14 VN.n13 5.84292
R1194 VN.n30 VN.n29 5.84292
R1195 VN.n37 VN.n36 5.84292
R1196 VN.n45 VN.n23 0.278398
R1197 VN.n22 VN.n0 0.278398
R1198 VN.n41 VN.n23 0.189894
R1199 VN.n41 VN.n40 0.189894
R1200 VN.n40 VN.n39 0.189894
R1201 VN.n39 VN.n25 0.189894
R1202 VN.n34 VN.n25 0.189894
R1203 VN.n34 VN.n33 0.189894
R1204 VN.n33 VN.n32 0.189894
R1205 VN.n32 VN.n27 0.189894
R1206 VN.n9 VN.n4 0.189894
R1207 VN.n10 VN.n9 0.189894
R1208 VN.n11 VN.n10 0.189894
R1209 VN.n11 VN.n2 0.189894
R1210 VN.n16 VN.n2 0.189894
R1211 VN.n17 VN.n16 0.189894
R1212 VN.n18 VN.n17 0.189894
R1213 VN.n18 VN.n0 0.189894
R1214 VN VN.n22 0.153422
R1215 VTAIL.n11 VTAIL.t1 60.8209
R1216 VTAIL.n10 VTAIL.t11 60.8209
R1217 VTAIL.n7 VTAIL.t9 60.8209
R1218 VTAIL.n15 VTAIL.t12 60.8207
R1219 VTAIL.n2 VTAIL.t8 60.8207
R1220 VTAIL.n3 VTAIL.t0 60.8207
R1221 VTAIL.n6 VTAIL.t15 60.8207
R1222 VTAIL.n14 VTAIL.t5 60.8207
R1223 VTAIL.n13 VTAIL.n12 58.4551
R1224 VTAIL.n9 VTAIL.n8 58.4551
R1225 VTAIL.n1 VTAIL.n0 58.4549
R1226 VTAIL.n5 VTAIL.n4 58.4549
R1227 VTAIL.n15 VTAIL.n14 26.1427
R1228 VTAIL.n7 VTAIL.n6 26.1427
R1229 VTAIL.n0 VTAIL.t10 2.36622
R1230 VTAIL.n0 VTAIL.t13 2.36622
R1231 VTAIL.n4 VTAIL.t2 2.36622
R1232 VTAIL.n4 VTAIL.t6 2.36622
R1233 VTAIL.n12 VTAIL.t4 2.36622
R1234 VTAIL.n12 VTAIL.t3 2.36622
R1235 VTAIL.n8 VTAIL.t7 2.36622
R1236 VTAIL.n8 VTAIL.t14 2.36622
R1237 VTAIL.n9 VTAIL.n7 1.93153
R1238 VTAIL.n10 VTAIL.n9 1.93153
R1239 VTAIL.n13 VTAIL.n11 1.93153
R1240 VTAIL.n14 VTAIL.n13 1.93153
R1241 VTAIL.n6 VTAIL.n5 1.93153
R1242 VTAIL.n5 VTAIL.n3 1.93153
R1243 VTAIL.n2 VTAIL.n1 1.93153
R1244 VTAIL VTAIL.n15 1.87334
R1245 VTAIL.n11 VTAIL.n10 0.470328
R1246 VTAIL.n3 VTAIL.n2 0.470328
R1247 VTAIL VTAIL.n1 0.0586897
R1248 VDD2.n2 VDD2.n1 76.0439
R1249 VDD2.n2 VDD2.n0 76.0439
R1250 VDD2 VDD2.n5 76.0411
R1251 VDD2.n4 VDD2.n3 75.1339
R1252 VDD2.n4 VDD2.n2 44.2498
R1253 VDD2.n5 VDD2.t2 2.36622
R1254 VDD2.n5 VDD2.t3 2.36622
R1255 VDD2.n3 VDD2.t4 2.36622
R1256 VDD2.n3 VDD2.t7 2.36622
R1257 VDD2.n1 VDD2.t1 2.36622
R1258 VDD2.n1 VDD2.t0 2.36622
R1259 VDD2.n0 VDD2.t5 2.36622
R1260 VDD2.n0 VDD2.t6 2.36622
R1261 VDD2 VDD2.n4 1.02421
R1262 VP.n12 VP.t7 203.144
R1263 VP.n31 VP.t6 173.369
R1264 VP.n38 VP.t5 173.369
R1265 VP.n46 VP.t2 173.369
R1266 VP.n53 VP.t1 173.369
R1267 VP.n28 VP.t4 173.369
R1268 VP.n21 VP.t3 173.369
R1269 VP.n13 VP.t0 173.369
R1270 VP.n14 VP.n11 161.3
R1271 VP.n16 VP.n15 161.3
R1272 VP.n17 VP.n10 161.3
R1273 VP.n19 VP.n18 161.3
R1274 VP.n20 VP.n9 161.3
R1275 VP.n23 VP.n22 161.3
R1276 VP.n24 VP.n8 161.3
R1277 VP.n26 VP.n25 161.3
R1278 VP.n27 VP.n7 161.3
R1279 VP.n52 VP.n0 161.3
R1280 VP.n51 VP.n50 161.3
R1281 VP.n49 VP.n1 161.3
R1282 VP.n48 VP.n47 161.3
R1283 VP.n45 VP.n2 161.3
R1284 VP.n44 VP.n43 161.3
R1285 VP.n42 VP.n3 161.3
R1286 VP.n41 VP.n40 161.3
R1287 VP.n39 VP.n4 161.3
R1288 VP.n37 VP.n36 161.3
R1289 VP.n35 VP.n5 161.3
R1290 VP.n34 VP.n33 161.3
R1291 VP.n32 VP.n6 161.3
R1292 VP.n31 VP.n30 93.0789
R1293 VP.n54 VP.n53 93.0789
R1294 VP.n29 VP.n28 93.0789
R1295 VP.n13 VP.n12 63.4148
R1296 VP.n33 VP.n5 56.4773
R1297 VP.n51 VP.n1 56.4773
R1298 VP.n26 VP.n8 56.4773
R1299 VP.n30 VP.n29 48.9541
R1300 VP.n40 VP.n3 40.4106
R1301 VP.n44 VP.n3 40.4106
R1302 VP.n19 VP.n10 40.4106
R1303 VP.n15 VP.n10 40.4106
R1304 VP.n33 VP.n32 24.3439
R1305 VP.n37 VP.n5 24.3439
R1306 VP.n40 VP.n39 24.3439
R1307 VP.n45 VP.n44 24.3439
R1308 VP.n47 VP.n1 24.3439
R1309 VP.n52 VP.n51 24.3439
R1310 VP.n27 VP.n26 24.3439
R1311 VP.n20 VP.n19 24.3439
R1312 VP.n22 VP.n8 24.3439
R1313 VP.n15 VP.n14 24.3439
R1314 VP.n38 VP.n37 18.5015
R1315 VP.n47 VP.n46 18.5015
R1316 VP.n22 VP.n21 18.5015
R1317 VP.n32 VP.n31 17.5278
R1318 VP.n53 VP.n52 17.5278
R1319 VP.n28 VP.n27 17.5278
R1320 VP.n12 VP.n11 13.6639
R1321 VP.n39 VP.n38 5.84292
R1322 VP.n46 VP.n45 5.84292
R1323 VP.n21 VP.n20 5.84292
R1324 VP.n14 VP.n13 5.84292
R1325 VP.n29 VP.n7 0.278398
R1326 VP.n30 VP.n6 0.278398
R1327 VP.n54 VP.n0 0.278398
R1328 VP.n16 VP.n11 0.189894
R1329 VP.n17 VP.n16 0.189894
R1330 VP.n18 VP.n17 0.189894
R1331 VP.n18 VP.n9 0.189894
R1332 VP.n23 VP.n9 0.189894
R1333 VP.n24 VP.n23 0.189894
R1334 VP.n25 VP.n24 0.189894
R1335 VP.n25 VP.n7 0.189894
R1336 VP.n34 VP.n6 0.189894
R1337 VP.n35 VP.n34 0.189894
R1338 VP.n36 VP.n35 0.189894
R1339 VP.n36 VP.n4 0.189894
R1340 VP.n41 VP.n4 0.189894
R1341 VP.n42 VP.n41 0.189894
R1342 VP.n43 VP.n42 0.189894
R1343 VP.n43 VP.n2 0.189894
R1344 VP.n48 VP.n2 0.189894
R1345 VP.n49 VP.n48 0.189894
R1346 VP.n50 VP.n49 0.189894
R1347 VP.n50 VP.n0 0.189894
R1348 VP VP.n54 0.153422
R1349 VDD1 VDD1.n0 76.1576
R1350 VDD1.n3 VDD1.n2 76.0439
R1351 VDD1.n3 VDD1.n1 76.0439
R1352 VDD1.n5 VDD1.n4 75.1338
R1353 VDD1.n5 VDD1.n3 44.8328
R1354 VDD1.n4 VDD1.t4 2.36622
R1355 VDD1.n4 VDD1.t3 2.36622
R1356 VDD1.n0 VDD1.t0 2.36622
R1357 VDD1.n0 VDD1.t7 2.36622
R1358 VDD1.n2 VDD1.t5 2.36622
R1359 VDD1.n2 VDD1.t6 2.36622
R1360 VDD1.n1 VDD1.t1 2.36622
R1361 VDD1.n1 VDD1.t2 2.36622
R1362 VDD1 VDD1.n5 0.907828
C0 VTAIL w_n3210_n3716# 4.56454f
C1 VTAIL VP 9.341089f
C2 VTAIL VDD2 8.885731f
C3 VTAIL VDD1 8.83594f
C4 VN w_n3210_n3716# 6.39198f
C5 VN VP 7.15046f
C6 VN VDD2 9.21538f
C7 w_n3210_n3716# B 9.54684f
C8 B VP 1.77331f
C9 VN VDD1 0.15023f
C10 B VDD2 1.56102f
C11 VDD1 B 1.4867f
C12 w_n3210_n3716# VP 6.80667f
C13 VTAIL VN 9.326981f
C14 w_n3210_n3716# VDD2 1.86394f
C15 VDD2 VP 0.445997f
C16 VDD1 w_n3210_n3716# 1.77818f
C17 VDD1 VP 9.510099f
C18 VTAIL B 5.18427f
C19 VDD1 VDD2 1.41895f
C20 VN B 1.08183f
C21 VDD2 VSUBS 1.645649f
C22 VDD1 VSUBS 2.167873f
C23 VTAIL VSUBS 1.298309f
C24 VN VSUBS 5.95717f
C25 VP VSUBS 2.946007f
C26 B VSUBS 4.377921f
C27 w_n3210_n3716# VSUBS 0.146492p
C28 VDD1.t0 VSUBS 0.268962f
C29 VDD1.t7 VSUBS 0.268962f
C30 VDD1.n0 VSUBS 2.17671f
C31 VDD1.t1 VSUBS 0.268962f
C32 VDD1.t2 VSUBS 0.268962f
C33 VDD1.n1 VSUBS 2.17557f
C34 VDD1.t5 VSUBS 0.268962f
C35 VDD1.t6 VSUBS 0.268962f
C36 VDD1.n2 VSUBS 2.17557f
C37 VDD1.n3 VSUBS 3.5087f
C38 VDD1.t4 VSUBS 0.268962f
C39 VDD1.t3 VSUBS 0.268962f
C40 VDD1.n4 VSUBS 2.16728f
C41 VDD1.n5 VSUBS 3.09898f
C42 VP.n0 VSUBS 0.044697f
C43 VP.t1 VSUBS 2.43279f
C44 VP.n1 VSUBS 0.048753f
C45 VP.n2 VSUBS 0.033901f
C46 VP.t2 VSUBS 2.43279f
C47 VP.n3 VSUBS 0.027433f
C48 VP.n4 VSUBS 0.033901f
C49 VP.t5 VSUBS 2.43279f
C50 VP.n5 VSUBS 0.048753f
C51 VP.n6 VSUBS 0.044697f
C52 VP.t6 VSUBS 2.43279f
C53 VP.n7 VSUBS 0.044697f
C54 VP.t4 VSUBS 2.43279f
C55 VP.n8 VSUBS 0.048753f
C56 VP.n9 VSUBS 0.033901f
C57 VP.t3 VSUBS 2.43279f
C58 VP.n10 VSUBS 0.027433f
C59 VP.n11 VSUBS 0.250782f
C60 VP.t0 VSUBS 2.43279f
C61 VP.t7 VSUBS 2.58239f
C62 VP.n12 VSUBS 0.953755f
C63 VP.n13 VSUBS 0.933459f
C64 VP.n14 VSUBS 0.039672f
C65 VP.n15 VSUBS 0.067737f
C66 VP.n16 VSUBS 0.033901f
C67 VP.n17 VSUBS 0.033901f
C68 VP.n18 VSUBS 0.033901f
C69 VP.n19 VSUBS 0.067737f
C70 VP.n20 VSUBS 0.039672f
C71 VP.n21 VSUBS 0.862445f
C72 VP.n22 VSUBS 0.055975f
C73 VP.n23 VSUBS 0.033901f
C74 VP.n24 VSUBS 0.033901f
C75 VP.n25 VSUBS 0.033901f
C76 VP.n26 VSUBS 0.050656f
C77 VP.n27 VSUBS 0.054721f
C78 VP.n28 VSUBS 0.95807f
C79 VP.n29 VSUBS 1.81396f
C80 VP.n30 VSUBS 1.83878f
C81 VP.n31 VSUBS 0.95807f
C82 VP.n32 VSUBS 0.054721f
C83 VP.n33 VSUBS 0.050656f
C84 VP.n34 VSUBS 0.033901f
C85 VP.n35 VSUBS 0.033901f
C86 VP.n36 VSUBS 0.033901f
C87 VP.n37 VSUBS 0.055975f
C88 VP.n38 VSUBS 0.862445f
C89 VP.n39 VSUBS 0.039672f
C90 VP.n40 VSUBS 0.067737f
C91 VP.n41 VSUBS 0.033901f
C92 VP.n42 VSUBS 0.033901f
C93 VP.n43 VSUBS 0.033901f
C94 VP.n44 VSUBS 0.067737f
C95 VP.n45 VSUBS 0.039672f
C96 VP.n46 VSUBS 0.862445f
C97 VP.n47 VSUBS 0.055975f
C98 VP.n48 VSUBS 0.033901f
C99 VP.n49 VSUBS 0.033901f
C100 VP.n50 VSUBS 0.033901f
C101 VP.n51 VSUBS 0.050656f
C102 VP.n52 VSUBS 0.054721f
C103 VP.n53 VSUBS 0.95807f
C104 VP.n54 VSUBS 0.042587f
C105 VDD2.t5 VSUBS 0.267359f
C106 VDD2.t6 VSUBS 0.267359f
C107 VDD2.n0 VSUBS 2.16261f
C108 VDD2.t1 VSUBS 0.267359f
C109 VDD2.t0 VSUBS 0.267359f
C110 VDD2.n1 VSUBS 2.16261f
C111 VDD2.n2 VSUBS 3.43617f
C112 VDD2.t4 VSUBS 0.267359f
C113 VDD2.t7 VSUBS 0.267359f
C114 VDD2.n3 VSUBS 2.15437f
C115 VDD2.n4 VSUBS 3.05041f
C116 VDD2.t2 VSUBS 0.267359f
C117 VDD2.t3 VSUBS 0.267359f
C118 VDD2.n5 VSUBS 2.16257f
C119 VTAIL.t10 VSUBS 0.261347f
C120 VTAIL.t13 VSUBS 0.261347f
C121 VTAIL.n0 VSUBS 1.98109f
C122 VTAIL.n1 VSUBS 0.688476f
C123 VTAIL.t8 VSUBS 2.59924f
C124 VTAIL.n2 VSUBS 0.81502f
C125 VTAIL.t0 VSUBS 2.59924f
C126 VTAIL.n3 VSUBS 0.81502f
C127 VTAIL.t2 VSUBS 0.261347f
C128 VTAIL.t6 VSUBS 0.261347f
C129 VTAIL.n4 VSUBS 1.98109f
C130 VTAIL.n5 VSUBS 0.833732f
C131 VTAIL.t15 VSUBS 2.59924f
C132 VTAIL.n6 VSUBS 2.17399f
C133 VTAIL.t9 VSUBS 2.59924f
C134 VTAIL.n7 VSUBS 2.17398f
C135 VTAIL.t7 VSUBS 0.261347f
C136 VTAIL.t14 VSUBS 0.261347f
C137 VTAIL.n8 VSUBS 1.98109f
C138 VTAIL.n9 VSUBS 0.833729f
C139 VTAIL.t11 VSUBS 2.59924f
C140 VTAIL.n10 VSUBS 0.815016f
C141 VTAIL.t1 VSUBS 2.59924f
C142 VTAIL.n11 VSUBS 0.815016f
C143 VTAIL.t4 VSUBS 0.261347f
C144 VTAIL.t3 VSUBS 0.261347f
C145 VTAIL.n12 VSUBS 1.98109f
C146 VTAIL.n13 VSUBS 0.833729f
C147 VTAIL.t5 VSUBS 2.59924f
C148 VTAIL.n14 VSUBS 2.17399f
C149 VTAIL.t12 VSUBS 2.59924f
C150 VTAIL.n15 VSUBS 2.16947f
C151 VN.n0 VSUBS 0.04368f
C152 VN.t7 VSUBS 2.37742f
C153 VN.n1 VSUBS 0.047643f
C154 VN.n2 VSUBS 0.033129f
C155 VN.t6 VSUBS 2.37742f
C156 VN.n3 VSUBS 0.026809f
C157 VN.n4 VSUBS 0.245074f
C158 VN.t1 VSUBS 2.37742f
C159 VN.t2 VSUBS 2.52361f
C160 VN.n5 VSUBS 0.932046f
C161 VN.n6 VSUBS 0.912213f
C162 VN.n7 VSUBS 0.038769f
C163 VN.n8 VSUBS 0.066196f
C164 VN.n9 VSUBS 0.033129f
C165 VN.n10 VSUBS 0.033129f
C166 VN.n11 VSUBS 0.033129f
C167 VN.n12 VSUBS 0.066196f
C168 VN.n13 VSUBS 0.038769f
C169 VN.n14 VSUBS 0.842814f
C170 VN.n15 VSUBS 0.054701f
C171 VN.n16 VSUBS 0.033129f
C172 VN.n17 VSUBS 0.033129f
C173 VN.n18 VSUBS 0.033129f
C174 VN.n19 VSUBS 0.049503f
C175 VN.n20 VSUBS 0.053475f
C176 VN.n21 VSUBS 0.936263f
C177 VN.n22 VSUBS 0.041618f
C178 VN.n23 VSUBS 0.04368f
C179 VN.t3 VSUBS 2.37742f
C180 VN.n24 VSUBS 0.047643f
C181 VN.n25 VSUBS 0.033129f
C182 VN.t0 VSUBS 2.37742f
C183 VN.n26 VSUBS 0.026809f
C184 VN.n27 VSUBS 0.245074f
C185 VN.t5 VSUBS 2.37742f
C186 VN.t4 VSUBS 2.52361f
C187 VN.n28 VSUBS 0.932046f
C188 VN.n29 VSUBS 0.912213f
C189 VN.n30 VSUBS 0.038769f
C190 VN.n31 VSUBS 0.066196f
C191 VN.n32 VSUBS 0.033129f
C192 VN.n33 VSUBS 0.033129f
C193 VN.n34 VSUBS 0.033129f
C194 VN.n35 VSUBS 0.066196f
C195 VN.n36 VSUBS 0.038769f
C196 VN.n37 VSUBS 0.842814f
C197 VN.n38 VSUBS 0.054701f
C198 VN.n39 VSUBS 0.033129f
C199 VN.n40 VSUBS 0.033129f
C200 VN.n41 VSUBS 0.033129f
C201 VN.n42 VSUBS 0.049503f
C202 VN.n43 VSUBS 0.053475f
C203 VN.n44 VSUBS 0.936263f
C204 VN.n45 VSUBS 1.79054f
C205 B.n0 VSUBS 0.004357f
C206 B.n1 VSUBS 0.004357f
C207 B.n2 VSUBS 0.00689f
C208 B.n3 VSUBS 0.00689f
C209 B.n4 VSUBS 0.00689f
C210 B.n5 VSUBS 0.00689f
C211 B.n6 VSUBS 0.00689f
C212 B.n7 VSUBS 0.00689f
C213 B.n8 VSUBS 0.00689f
C214 B.n9 VSUBS 0.00689f
C215 B.n10 VSUBS 0.00689f
C216 B.n11 VSUBS 0.00689f
C217 B.n12 VSUBS 0.00689f
C218 B.n13 VSUBS 0.00689f
C219 B.n14 VSUBS 0.00689f
C220 B.n15 VSUBS 0.00689f
C221 B.n16 VSUBS 0.00689f
C222 B.n17 VSUBS 0.00689f
C223 B.n18 VSUBS 0.00689f
C224 B.n19 VSUBS 0.00689f
C225 B.n20 VSUBS 0.00689f
C226 B.n21 VSUBS 0.00689f
C227 B.n22 VSUBS 0.015913f
C228 B.n23 VSUBS 0.00689f
C229 B.n24 VSUBS 0.00689f
C230 B.n25 VSUBS 0.00689f
C231 B.n26 VSUBS 0.00689f
C232 B.n27 VSUBS 0.00689f
C233 B.n28 VSUBS 0.00689f
C234 B.n29 VSUBS 0.00689f
C235 B.n30 VSUBS 0.00689f
C236 B.n31 VSUBS 0.00689f
C237 B.n32 VSUBS 0.00689f
C238 B.n33 VSUBS 0.00689f
C239 B.n34 VSUBS 0.00689f
C240 B.n35 VSUBS 0.00689f
C241 B.n36 VSUBS 0.00689f
C242 B.n37 VSUBS 0.00689f
C243 B.n38 VSUBS 0.00689f
C244 B.n39 VSUBS 0.00689f
C245 B.n40 VSUBS 0.00689f
C246 B.n41 VSUBS 0.00689f
C247 B.n42 VSUBS 0.00689f
C248 B.n43 VSUBS 0.00689f
C249 B.n44 VSUBS 0.00689f
C250 B.n45 VSUBS 0.00689f
C251 B.t8 VSUBS 0.44671f
C252 B.t7 VSUBS 0.463227f
C253 B.t6 VSUBS 1.14031f
C254 B.n46 VSUBS 0.222014f
C255 B.n47 VSUBS 0.067961f
C256 B.n48 VSUBS 0.015963f
C257 B.n49 VSUBS 0.00689f
C258 B.n50 VSUBS 0.00689f
C259 B.n51 VSUBS 0.00689f
C260 B.n52 VSUBS 0.00689f
C261 B.n53 VSUBS 0.00689f
C262 B.t5 VSUBS 0.446699f
C263 B.t4 VSUBS 0.463217f
C264 B.t3 VSUBS 1.14031f
C265 B.n54 VSUBS 0.222024f
C266 B.n55 VSUBS 0.067972f
C267 B.n56 VSUBS 0.00689f
C268 B.n57 VSUBS 0.00689f
C269 B.n58 VSUBS 0.00689f
C270 B.n59 VSUBS 0.00689f
C271 B.n60 VSUBS 0.00689f
C272 B.n61 VSUBS 0.00689f
C273 B.n62 VSUBS 0.00689f
C274 B.n63 VSUBS 0.00689f
C275 B.n64 VSUBS 0.00689f
C276 B.n65 VSUBS 0.00689f
C277 B.n66 VSUBS 0.00689f
C278 B.n67 VSUBS 0.00689f
C279 B.n68 VSUBS 0.00689f
C280 B.n69 VSUBS 0.00689f
C281 B.n70 VSUBS 0.00689f
C282 B.n71 VSUBS 0.00689f
C283 B.n72 VSUBS 0.00689f
C284 B.n73 VSUBS 0.00689f
C285 B.n74 VSUBS 0.00689f
C286 B.n75 VSUBS 0.00689f
C287 B.n76 VSUBS 0.00689f
C288 B.n77 VSUBS 0.00689f
C289 B.n78 VSUBS 0.015913f
C290 B.n79 VSUBS 0.00689f
C291 B.n80 VSUBS 0.00689f
C292 B.n81 VSUBS 0.00689f
C293 B.n82 VSUBS 0.00689f
C294 B.n83 VSUBS 0.00689f
C295 B.n84 VSUBS 0.00689f
C296 B.n85 VSUBS 0.00689f
C297 B.n86 VSUBS 0.00689f
C298 B.n87 VSUBS 0.00689f
C299 B.n88 VSUBS 0.00689f
C300 B.n89 VSUBS 0.00689f
C301 B.n90 VSUBS 0.00689f
C302 B.n91 VSUBS 0.00689f
C303 B.n92 VSUBS 0.00689f
C304 B.n93 VSUBS 0.00689f
C305 B.n94 VSUBS 0.00689f
C306 B.n95 VSUBS 0.00689f
C307 B.n96 VSUBS 0.00689f
C308 B.n97 VSUBS 0.00689f
C309 B.n98 VSUBS 0.00689f
C310 B.n99 VSUBS 0.00689f
C311 B.n100 VSUBS 0.00689f
C312 B.n101 VSUBS 0.00689f
C313 B.n102 VSUBS 0.00689f
C314 B.n103 VSUBS 0.00689f
C315 B.n104 VSUBS 0.00689f
C316 B.n105 VSUBS 0.00689f
C317 B.n106 VSUBS 0.00689f
C318 B.n107 VSUBS 0.00689f
C319 B.n108 VSUBS 0.00689f
C320 B.n109 VSUBS 0.00689f
C321 B.n110 VSUBS 0.00689f
C322 B.n111 VSUBS 0.00689f
C323 B.n112 VSUBS 0.00689f
C324 B.n113 VSUBS 0.00689f
C325 B.n114 VSUBS 0.00689f
C326 B.n115 VSUBS 0.00689f
C327 B.n116 VSUBS 0.00689f
C328 B.n117 VSUBS 0.00689f
C329 B.n118 VSUBS 0.00689f
C330 B.n119 VSUBS 0.00689f
C331 B.n120 VSUBS 0.016712f
C332 B.n121 VSUBS 0.00689f
C333 B.n122 VSUBS 0.00689f
C334 B.n123 VSUBS 0.00689f
C335 B.n124 VSUBS 0.00689f
C336 B.n125 VSUBS 0.00689f
C337 B.n126 VSUBS 0.00689f
C338 B.n127 VSUBS 0.00689f
C339 B.n128 VSUBS 0.00689f
C340 B.n129 VSUBS 0.00689f
C341 B.n130 VSUBS 0.00689f
C342 B.n131 VSUBS 0.00689f
C343 B.n132 VSUBS 0.00689f
C344 B.n133 VSUBS 0.00689f
C345 B.n134 VSUBS 0.00689f
C346 B.n135 VSUBS 0.00689f
C347 B.n136 VSUBS 0.00689f
C348 B.n137 VSUBS 0.00689f
C349 B.n138 VSUBS 0.00689f
C350 B.n139 VSUBS 0.00689f
C351 B.n140 VSUBS 0.00689f
C352 B.n141 VSUBS 0.00689f
C353 B.n142 VSUBS 0.00689f
C354 B.n143 VSUBS 0.00689f
C355 B.t1 VSUBS 0.446699f
C356 B.t2 VSUBS 0.463217f
C357 B.t0 VSUBS 1.14031f
C358 B.n144 VSUBS 0.222024f
C359 B.n145 VSUBS 0.067972f
C360 B.n146 VSUBS 0.00689f
C361 B.n147 VSUBS 0.00689f
C362 B.n148 VSUBS 0.00689f
C363 B.n149 VSUBS 0.00689f
C364 B.t10 VSUBS 0.44671f
C365 B.t11 VSUBS 0.463227f
C366 B.t9 VSUBS 1.14031f
C367 B.n150 VSUBS 0.222014f
C368 B.n151 VSUBS 0.067961f
C369 B.n152 VSUBS 0.015963f
C370 B.n153 VSUBS 0.00689f
C371 B.n154 VSUBS 0.00689f
C372 B.n155 VSUBS 0.00689f
C373 B.n156 VSUBS 0.00689f
C374 B.n157 VSUBS 0.00689f
C375 B.n158 VSUBS 0.00689f
C376 B.n159 VSUBS 0.00689f
C377 B.n160 VSUBS 0.00689f
C378 B.n161 VSUBS 0.00689f
C379 B.n162 VSUBS 0.00689f
C380 B.n163 VSUBS 0.00689f
C381 B.n164 VSUBS 0.00689f
C382 B.n165 VSUBS 0.00689f
C383 B.n166 VSUBS 0.00689f
C384 B.n167 VSUBS 0.00689f
C385 B.n168 VSUBS 0.00689f
C386 B.n169 VSUBS 0.00689f
C387 B.n170 VSUBS 0.00689f
C388 B.n171 VSUBS 0.00689f
C389 B.n172 VSUBS 0.00689f
C390 B.n173 VSUBS 0.00689f
C391 B.n174 VSUBS 0.00689f
C392 B.n175 VSUBS 0.00689f
C393 B.n176 VSUBS 0.015913f
C394 B.n177 VSUBS 0.00689f
C395 B.n178 VSUBS 0.00689f
C396 B.n179 VSUBS 0.00689f
C397 B.n180 VSUBS 0.00689f
C398 B.n181 VSUBS 0.00689f
C399 B.n182 VSUBS 0.00689f
C400 B.n183 VSUBS 0.00689f
C401 B.n184 VSUBS 0.00689f
C402 B.n185 VSUBS 0.00689f
C403 B.n186 VSUBS 0.00689f
C404 B.n187 VSUBS 0.00689f
C405 B.n188 VSUBS 0.00689f
C406 B.n189 VSUBS 0.00689f
C407 B.n190 VSUBS 0.00689f
C408 B.n191 VSUBS 0.00689f
C409 B.n192 VSUBS 0.00689f
C410 B.n193 VSUBS 0.00689f
C411 B.n194 VSUBS 0.00689f
C412 B.n195 VSUBS 0.00689f
C413 B.n196 VSUBS 0.00689f
C414 B.n197 VSUBS 0.00689f
C415 B.n198 VSUBS 0.00689f
C416 B.n199 VSUBS 0.00689f
C417 B.n200 VSUBS 0.00689f
C418 B.n201 VSUBS 0.00689f
C419 B.n202 VSUBS 0.00689f
C420 B.n203 VSUBS 0.00689f
C421 B.n204 VSUBS 0.00689f
C422 B.n205 VSUBS 0.00689f
C423 B.n206 VSUBS 0.00689f
C424 B.n207 VSUBS 0.00689f
C425 B.n208 VSUBS 0.00689f
C426 B.n209 VSUBS 0.00689f
C427 B.n210 VSUBS 0.00689f
C428 B.n211 VSUBS 0.00689f
C429 B.n212 VSUBS 0.00689f
C430 B.n213 VSUBS 0.00689f
C431 B.n214 VSUBS 0.00689f
C432 B.n215 VSUBS 0.00689f
C433 B.n216 VSUBS 0.00689f
C434 B.n217 VSUBS 0.00689f
C435 B.n218 VSUBS 0.00689f
C436 B.n219 VSUBS 0.00689f
C437 B.n220 VSUBS 0.00689f
C438 B.n221 VSUBS 0.00689f
C439 B.n222 VSUBS 0.00689f
C440 B.n223 VSUBS 0.00689f
C441 B.n224 VSUBS 0.00689f
C442 B.n225 VSUBS 0.00689f
C443 B.n226 VSUBS 0.00689f
C444 B.n227 VSUBS 0.00689f
C445 B.n228 VSUBS 0.00689f
C446 B.n229 VSUBS 0.00689f
C447 B.n230 VSUBS 0.00689f
C448 B.n231 VSUBS 0.00689f
C449 B.n232 VSUBS 0.00689f
C450 B.n233 VSUBS 0.00689f
C451 B.n234 VSUBS 0.00689f
C452 B.n235 VSUBS 0.00689f
C453 B.n236 VSUBS 0.00689f
C454 B.n237 VSUBS 0.00689f
C455 B.n238 VSUBS 0.00689f
C456 B.n239 VSUBS 0.00689f
C457 B.n240 VSUBS 0.00689f
C458 B.n241 VSUBS 0.00689f
C459 B.n242 VSUBS 0.00689f
C460 B.n243 VSUBS 0.00689f
C461 B.n244 VSUBS 0.00689f
C462 B.n245 VSUBS 0.00689f
C463 B.n246 VSUBS 0.00689f
C464 B.n247 VSUBS 0.00689f
C465 B.n248 VSUBS 0.00689f
C466 B.n249 VSUBS 0.00689f
C467 B.n250 VSUBS 0.00689f
C468 B.n251 VSUBS 0.00689f
C469 B.n252 VSUBS 0.00689f
C470 B.n253 VSUBS 0.00689f
C471 B.n254 VSUBS 0.00689f
C472 B.n255 VSUBS 0.015913f
C473 B.n256 VSUBS 0.016712f
C474 B.n257 VSUBS 0.016712f
C475 B.n258 VSUBS 0.00689f
C476 B.n259 VSUBS 0.00689f
C477 B.n260 VSUBS 0.00689f
C478 B.n261 VSUBS 0.00689f
C479 B.n262 VSUBS 0.00689f
C480 B.n263 VSUBS 0.00689f
C481 B.n264 VSUBS 0.00689f
C482 B.n265 VSUBS 0.00689f
C483 B.n266 VSUBS 0.00689f
C484 B.n267 VSUBS 0.00689f
C485 B.n268 VSUBS 0.00689f
C486 B.n269 VSUBS 0.00689f
C487 B.n270 VSUBS 0.00689f
C488 B.n271 VSUBS 0.00689f
C489 B.n272 VSUBS 0.00689f
C490 B.n273 VSUBS 0.00689f
C491 B.n274 VSUBS 0.00689f
C492 B.n275 VSUBS 0.00689f
C493 B.n276 VSUBS 0.00689f
C494 B.n277 VSUBS 0.00689f
C495 B.n278 VSUBS 0.00689f
C496 B.n279 VSUBS 0.00689f
C497 B.n280 VSUBS 0.00689f
C498 B.n281 VSUBS 0.00689f
C499 B.n282 VSUBS 0.00689f
C500 B.n283 VSUBS 0.00689f
C501 B.n284 VSUBS 0.00689f
C502 B.n285 VSUBS 0.00689f
C503 B.n286 VSUBS 0.00689f
C504 B.n287 VSUBS 0.00689f
C505 B.n288 VSUBS 0.00689f
C506 B.n289 VSUBS 0.00689f
C507 B.n290 VSUBS 0.00689f
C508 B.n291 VSUBS 0.00689f
C509 B.n292 VSUBS 0.00689f
C510 B.n293 VSUBS 0.00689f
C511 B.n294 VSUBS 0.00689f
C512 B.n295 VSUBS 0.00689f
C513 B.n296 VSUBS 0.00689f
C514 B.n297 VSUBS 0.00689f
C515 B.n298 VSUBS 0.00689f
C516 B.n299 VSUBS 0.00689f
C517 B.n300 VSUBS 0.00689f
C518 B.n301 VSUBS 0.00689f
C519 B.n302 VSUBS 0.00689f
C520 B.n303 VSUBS 0.00689f
C521 B.n304 VSUBS 0.00689f
C522 B.n305 VSUBS 0.00689f
C523 B.n306 VSUBS 0.00689f
C524 B.n307 VSUBS 0.00689f
C525 B.n308 VSUBS 0.00689f
C526 B.n309 VSUBS 0.00689f
C527 B.n310 VSUBS 0.00689f
C528 B.n311 VSUBS 0.00689f
C529 B.n312 VSUBS 0.00689f
C530 B.n313 VSUBS 0.00689f
C531 B.n314 VSUBS 0.00689f
C532 B.n315 VSUBS 0.00689f
C533 B.n316 VSUBS 0.00689f
C534 B.n317 VSUBS 0.00689f
C535 B.n318 VSUBS 0.00689f
C536 B.n319 VSUBS 0.00689f
C537 B.n320 VSUBS 0.00689f
C538 B.n321 VSUBS 0.00689f
C539 B.n322 VSUBS 0.00689f
C540 B.n323 VSUBS 0.00689f
C541 B.n324 VSUBS 0.00689f
C542 B.n325 VSUBS 0.004762f
C543 B.n326 VSUBS 0.00689f
C544 B.n327 VSUBS 0.00689f
C545 B.n328 VSUBS 0.005573f
C546 B.n329 VSUBS 0.00689f
C547 B.n330 VSUBS 0.00689f
C548 B.n331 VSUBS 0.00689f
C549 B.n332 VSUBS 0.00689f
C550 B.n333 VSUBS 0.00689f
C551 B.n334 VSUBS 0.00689f
C552 B.n335 VSUBS 0.00689f
C553 B.n336 VSUBS 0.00689f
C554 B.n337 VSUBS 0.00689f
C555 B.n338 VSUBS 0.00689f
C556 B.n339 VSUBS 0.00689f
C557 B.n340 VSUBS 0.005573f
C558 B.n341 VSUBS 0.015963f
C559 B.n342 VSUBS 0.004762f
C560 B.n343 VSUBS 0.00689f
C561 B.n344 VSUBS 0.00689f
C562 B.n345 VSUBS 0.00689f
C563 B.n346 VSUBS 0.00689f
C564 B.n347 VSUBS 0.00689f
C565 B.n348 VSUBS 0.00689f
C566 B.n349 VSUBS 0.00689f
C567 B.n350 VSUBS 0.00689f
C568 B.n351 VSUBS 0.00689f
C569 B.n352 VSUBS 0.00689f
C570 B.n353 VSUBS 0.00689f
C571 B.n354 VSUBS 0.00689f
C572 B.n355 VSUBS 0.00689f
C573 B.n356 VSUBS 0.00689f
C574 B.n357 VSUBS 0.00689f
C575 B.n358 VSUBS 0.00689f
C576 B.n359 VSUBS 0.00689f
C577 B.n360 VSUBS 0.00689f
C578 B.n361 VSUBS 0.00689f
C579 B.n362 VSUBS 0.00689f
C580 B.n363 VSUBS 0.00689f
C581 B.n364 VSUBS 0.00689f
C582 B.n365 VSUBS 0.00689f
C583 B.n366 VSUBS 0.00689f
C584 B.n367 VSUBS 0.00689f
C585 B.n368 VSUBS 0.00689f
C586 B.n369 VSUBS 0.00689f
C587 B.n370 VSUBS 0.00689f
C588 B.n371 VSUBS 0.00689f
C589 B.n372 VSUBS 0.00689f
C590 B.n373 VSUBS 0.00689f
C591 B.n374 VSUBS 0.00689f
C592 B.n375 VSUBS 0.00689f
C593 B.n376 VSUBS 0.00689f
C594 B.n377 VSUBS 0.00689f
C595 B.n378 VSUBS 0.00689f
C596 B.n379 VSUBS 0.00689f
C597 B.n380 VSUBS 0.00689f
C598 B.n381 VSUBS 0.00689f
C599 B.n382 VSUBS 0.00689f
C600 B.n383 VSUBS 0.00689f
C601 B.n384 VSUBS 0.00689f
C602 B.n385 VSUBS 0.00689f
C603 B.n386 VSUBS 0.00689f
C604 B.n387 VSUBS 0.00689f
C605 B.n388 VSUBS 0.00689f
C606 B.n389 VSUBS 0.00689f
C607 B.n390 VSUBS 0.00689f
C608 B.n391 VSUBS 0.00689f
C609 B.n392 VSUBS 0.00689f
C610 B.n393 VSUBS 0.00689f
C611 B.n394 VSUBS 0.00689f
C612 B.n395 VSUBS 0.00689f
C613 B.n396 VSUBS 0.00689f
C614 B.n397 VSUBS 0.00689f
C615 B.n398 VSUBS 0.00689f
C616 B.n399 VSUBS 0.00689f
C617 B.n400 VSUBS 0.00689f
C618 B.n401 VSUBS 0.00689f
C619 B.n402 VSUBS 0.00689f
C620 B.n403 VSUBS 0.00689f
C621 B.n404 VSUBS 0.00689f
C622 B.n405 VSUBS 0.00689f
C623 B.n406 VSUBS 0.00689f
C624 B.n407 VSUBS 0.00689f
C625 B.n408 VSUBS 0.00689f
C626 B.n409 VSUBS 0.00689f
C627 B.n410 VSUBS 0.00689f
C628 B.n411 VSUBS 0.016712f
C629 B.n412 VSUBS 0.015913f
C630 B.n413 VSUBS 0.015913f
C631 B.n414 VSUBS 0.00689f
C632 B.n415 VSUBS 0.00689f
C633 B.n416 VSUBS 0.00689f
C634 B.n417 VSUBS 0.00689f
C635 B.n418 VSUBS 0.00689f
C636 B.n419 VSUBS 0.00689f
C637 B.n420 VSUBS 0.00689f
C638 B.n421 VSUBS 0.00689f
C639 B.n422 VSUBS 0.00689f
C640 B.n423 VSUBS 0.00689f
C641 B.n424 VSUBS 0.00689f
C642 B.n425 VSUBS 0.00689f
C643 B.n426 VSUBS 0.00689f
C644 B.n427 VSUBS 0.00689f
C645 B.n428 VSUBS 0.00689f
C646 B.n429 VSUBS 0.00689f
C647 B.n430 VSUBS 0.00689f
C648 B.n431 VSUBS 0.00689f
C649 B.n432 VSUBS 0.00689f
C650 B.n433 VSUBS 0.00689f
C651 B.n434 VSUBS 0.00689f
C652 B.n435 VSUBS 0.00689f
C653 B.n436 VSUBS 0.00689f
C654 B.n437 VSUBS 0.00689f
C655 B.n438 VSUBS 0.00689f
C656 B.n439 VSUBS 0.00689f
C657 B.n440 VSUBS 0.00689f
C658 B.n441 VSUBS 0.00689f
C659 B.n442 VSUBS 0.00689f
C660 B.n443 VSUBS 0.00689f
C661 B.n444 VSUBS 0.00689f
C662 B.n445 VSUBS 0.00689f
C663 B.n446 VSUBS 0.00689f
C664 B.n447 VSUBS 0.00689f
C665 B.n448 VSUBS 0.00689f
C666 B.n449 VSUBS 0.00689f
C667 B.n450 VSUBS 0.00689f
C668 B.n451 VSUBS 0.00689f
C669 B.n452 VSUBS 0.00689f
C670 B.n453 VSUBS 0.00689f
C671 B.n454 VSUBS 0.00689f
C672 B.n455 VSUBS 0.00689f
C673 B.n456 VSUBS 0.00689f
C674 B.n457 VSUBS 0.00689f
C675 B.n458 VSUBS 0.00689f
C676 B.n459 VSUBS 0.00689f
C677 B.n460 VSUBS 0.00689f
C678 B.n461 VSUBS 0.00689f
C679 B.n462 VSUBS 0.00689f
C680 B.n463 VSUBS 0.00689f
C681 B.n464 VSUBS 0.00689f
C682 B.n465 VSUBS 0.00689f
C683 B.n466 VSUBS 0.00689f
C684 B.n467 VSUBS 0.00689f
C685 B.n468 VSUBS 0.00689f
C686 B.n469 VSUBS 0.00689f
C687 B.n470 VSUBS 0.00689f
C688 B.n471 VSUBS 0.00689f
C689 B.n472 VSUBS 0.00689f
C690 B.n473 VSUBS 0.00689f
C691 B.n474 VSUBS 0.00689f
C692 B.n475 VSUBS 0.00689f
C693 B.n476 VSUBS 0.00689f
C694 B.n477 VSUBS 0.00689f
C695 B.n478 VSUBS 0.00689f
C696 B.n479 VSUBS 0.00689f
C697 B.n480 VSUBS 0.00689f
C698 B.n481 VSUBS 0.00689f
C699 B.n482 VSUBS 0.00689f
C700 B.n483 VSUBS 0.00689f
C701 B.n484 VSUBS 0.00689f
C702 B.n485 VSUBS 0.00689f
C703 B.n486 VSUBS 0.00689f
C704 B.n487 VSUBS 0.00689f
C705 B.n488 VSUBS 0.00689f
C706 B.n489 VSUBS 0.00689f
C707 B.n490 VSUBS 0.00689f
C708 B.n491 VSUBS 0.00689f
C709 B.n492 VSUBS 0.00689f
C710 B.n493 VSUBS 0.00689f
C711 B.n494 VSUBS 0.00689f
C712 B.n495 VSUBS 0.00689f
C713 B.n496 VSUBS 0.00689f
C714 B.n497 VSUBS 0.00689f
C715 B.n498 VSUBS 0.00689f
C716 B.n499 VSUBS 0.00689f
C717 B.n500 VSUBS 0.00689f
C718 B.n501 VSUBS 0.00689f
C719 B.n502 VSUBS 0.00689f
C720 B.n503 VSUBS 0.00689f
C721 B.n504 VSUBS 0.00689f
C722 B.n505 VSUBS 0.00689f
C723 B.n506 VSUBS 0.00689f
C724 B.n507 VSUBS 0.00689f
C725 B.n508 VSUBS 0.00689f
C726 B.n509 VSUBS 0.00689f
C727 B.n510 VSUBS 0.00689f
C728 B.n511 VSUBS 0.00689f
C729 B.n512 VSUBS 0.00689f
C730 B.n513 VSUBS 0.00689f
C731 B.n514 VSUBS 0.00689f
C732 B.n515 VSUBS 0.00689f
C733 B.n516 VSUBS 0.00689f
C734 B.n517 VSUBS 0.00689f
C735 B.n518 VSUBS 0.00689f
C736 B.n519 VSUBS 0.00689f
C737 B.n520 VSUBS 0.00689f
C738 B.n521 VSUBS 0.00689f
C739 B.n522 VSUBS 0.00689f
C740 B.n523 VSUBS 0.00689f
C741 B.n524 VSUBS 0.00689f
C742 B.n525 VSUBS 0.00689f
C743 B.n526 VSUBS 0.00689f
C744 B.n527 VSUBS 0.00689f
C745 B.n528 VSUBS 0.00689f
C746 B.n529 VSUBS 0.00689f
C747 B.n530 VSUBS 0.00689f
C748 B.n531 VSUBS 0.00689f
C749 B.n532 VSUBS 0.00689f
C750 B.n533 VSUBS 0.00689f
C751 B.n534 VSUBS 0.00689f
C752 B.n535 VSUBS 0.016712f
C753 B.n536 VSUBS 0.015913f
C754 B.n537 VSUBS 0.016712f
C755 B.n538 VSUBS 0.00689f
C756 B.n539 VSUBS 0.00689f
C757 B.n540 VSUBS 0.00689f
C758 B.n541 VSUBS 0.00689f
C759 B.n542 VSUBS 0.00689f
C760 B.n543 VSUBS 0.00689f
C761 B.n544 VSUBS 0.00689f
C762 B.n545 VSUBS 0.00689f
C763 B.n546 VSUBS 0.00689f
C764 B.n547 VSUBS 0.00689f
C765 B.n548 VSUBS 0.00689f
C766 B.n549 VSUBS 0.00689f
C767 B.n550 VSUBS 0.00689f
C768 B.n551 VSUBS 0.00689f
C769 B.n552 VSUBS 0.00689f
C770 B.n553 VSUBS 0.00689f
C771 B.n554 VSUBS 0.00689f
C772 B.n555 VSUBS 0.00689f
C773 B.n556 VSUBS 0.00689f
C774 B.n557 VSUBS 0.00689f
C775 B.n558 VSUBS 0.00689f
C776 B.n559 VSUBS 0.00689f
C777 B.n560 VSUBS 0.00689f
C778 B.n561 VSUBS 0.00689f
C779 B.n562 VSUBS 0.00689f
C780 B.n563 VSUBS 0.00689f
C781 B.n564 VSUBS 0.00689f
C782 B.n565 VSUBS 0.00689f
C783 B.n566 VSUBS 0.00689f
C784 B.n567 VSUBS 0.00689f
C785 B.n568 VSUBS 0.00689f
C786 B.n569 VSUBS 0.00689f
C787 B.n570 VSUBS 0.00689f
C788 B.n571 VSUBS 0.00689f
C789 B.n572 VSUBS 0.00689f
C790 B.n573 VSUBS 0.00689f
C791 B.n574 VSUBS 0.00689f
C792 B.n575 VSUBS 0.00689f
C793 B.n576 VSUBS 0.00689f
C794 B.n577 VSUBS 0.00689f
C795 B.n578 VSUBS 0.00689f
C796 B.n579 VSUBS 0.00689f
C797 B.n580 VSUBS 0.00689f
C798 B.n581 VSUBS 0.00689f
C799 B.n582 VSUBS 0.00689f
C800 B.n583 VSUBS 0.00689f
C801 B.n584 VSUBS 0.00689f
C802 B.n585 VSUBS 0.00689f
C803 B.n586 VSUBS 0.00689f
C804 B.n587 VSUBS 0.00689f
C805 B.n588 VSUBS 0.00689f
C806 B.n589 VSUBS 0.00689f
C807 B.n590 VSUBS 0.00689f
C808 B.n591 VSUBS 0.00689f
C809 B.n592 VSUBS 0.00689f
C810 B.n593 VSUBS 0.00689f
C811 B.n594 VSUBS 0.00689f
C812 B.n595 VSUBS 0.00689f
C813 B.n596 VSUBS 0.00689f
C814 B.n597 VSUBS 0.00689f
C815 B.n598 VSUBS 0.00689f
C816 B.n599 VSUBS 0.00689f
C817 B.n600 VSUBS 0.00689f
C818 B.n601 VSUBS 0.00689f
C819 B.n602 VSUBS 0.00689f
C820 B.n603 VSUBS 0.00689f
C821 B.n604 VSUBS 0.00689f
C822 B.n605 VSUBS 0.00689f
C823 B.n606 VSUBS 0.004762f
C824 B.n607 VSUBS 0.015963f
C825 B.n608 VSUBS 0.005573f
C826 B.n609 VSUBS 0.00689f
C827 B.n610 VSUBS 0.00689f
C828 B.n611 VSUBS 0.00689f
C829 B.n612 VSUBS 0.00689f
C830 B.n613 VSUBS 0.00689f
C831 B.n614 VSUBS 0.00689f
C832 B.n615 VSUBS 0.00689f
C833 B.n616 VSUBS 0.00689f
C834 B.n617 VSUBS 0.00689f
C835 B.n618 VSUBS 0.00689f
C836 B.n619 VSUBS 0.00689f
C837 B.n620 VSUBS 0.005573f
C838 B.n621 VSUBS 0.00689f
C839 B.n622 VSUBS 0.00689f
C840 B.n623 VSUBS 0.004762f
C841 B.n624 VSUBS 0.00689f
C842 B.n625 VSUBS 0.00689f
C843 B.n626 VSUBS 0.00689f
C844 B.n627 VSUBS 0.00689f
C845 B.n628 VSUBS 0.00689f
C846 B.n629 VSUBS 0.00689f
C847 B.n630 VSUBS 0.00689f
C848 B.n631 VSUBS 0.00689f
C849 B.n632 VSUBS 0.00689f
C850 B.n633 VSUBS 0.00689f
C851 B.n634 VSUBS 0.00689f
C852 B.n635 VSUBS 0.00689f
C853 B.n636 VSUBS 0.00689f
C854 B.n637 VSUBS 0.00689f
C855 B.n638 VSUBS 0.00689f
C856 B.n639 VSUBS 0.00689f
C857 B.n640 VSUBS 0.00689f
C858 B.n641 VSUBS 0.00689f
C859 B.n642 VSUBS 0.00689f
C860 B.n643 VSUBS 0.00689f
C861 B.n644 VSUBS 0.00689f
C862 B.n645 VSUBS 0.00689f
C863 B.n646 VSUBS 0.00689f
C864 B.n647 VSUBS 0.00689f
C865 B.n648 VSUBS 0.00689f
C866 B.n649 VSUBS 0.00689f
C867 B.n650 VSUBS 0.00689f
C868 B.n651 VSUBS 0.00689f
C869 B.n652 VSUBS 0.00689f
C870 B.n653 VSUBS 0.00689f
C871 B.n654 VSUBS 0.00689f
C872 B.n655 VSUBS 0.00689f
C873 B.n656 VSUBS 0.00689f
C874 B.n657 VSUBS 0.00689f
C875 B.n658 VSUBS 0.00689f
C876 B.n659 VSUBS 0.00689f
C877 B.n660 VSUBS 0.00689f
C878 B.n661 VSUBS 0.00689f
C879 B.n662 VSUBS 0.00689f
C880 B.n663 VSUBS 0.00689f
C881 B.n664 VSUBS 0.00689f
C882 B.n665 VSUBS 0.00689f
C883 B.n666 VSUBS 0.00689f
C884 B.n667 VSUBS 0.00689f
C885 B.n668 VSUBS 0.00689f
C886 B.n669 VSUBS 0.00689f
C887 B.n670 VSUBS 0.00689f
C888 B.n671 VSUBS 0.00689f
C889 B.n672 VSUBS 0.00689f
C890 B.n673 VSUBS 0.00689f
C891 B.n674 VSUBS 0.00689f
C892 B.n675 VSUBS 0.00689f
C893 B.n676 VSUBS 0.00689f
C894 B.n677 VSUBS 0.00689f
C895 B.n678 VSUBS 0.00689f
C896 B.n679 VSUBS 0.00689f
C897 B.n680 VSUBS 0.00689f
C898 B.n681 VSUBS 0.00689f
C899 B.n682 VSUBS 0.00689f
C900 B.n683 VSUBS 0.00689f
C901 B.n684 VSUBS 0.00689f
C902 B.n685 VSUBS 0.00689f
C903 B.n686 VSUBS 0.00689f
C904 B.n687 VSUBS 0.00689f
C905 B.n688 VSUBS 0.00689f
C906 B.n689 VSUBS 0.00689f
C907 B.n690 VSUBS 0.00689f
C908 B.n691 VSUBS 0.016712f
C909 B.n692 VSUBS 0.016712f
C910 B.n693 VSUBS 0.015913f
C911 B.n694 VSUBS 0.00689f
C912 B.n695 VSUBS 0.00689f
C913 B.n696 VSUBS 0.00689f
C914 B.n697 VSUBS 0.00689f
C915 B.n698 VSUBS 0.00689f
C916 B.n699 VSUBS 0.00689f
C917 B.n700 VSUBS 0.00689f
C918 B.n701 VSUBS 0.00689f
C919 B.n702 VSUBS 0.00689f
C920 B.n703 VSUBS 0.00689f
C921 B.n704 VSUBS 0.00689f
C922 B.n705 VSUBS 0.00689f
C923 B.n706 VSUBS 0.00689f
C924 B.n707 VSUBS 0.00689f
C925 B.n708 VSUBS 0.00689f
C926 B.n709 VSUBS 0.00689f
C927 B.n710 VSUBS 0.00689f
C928 B.n711 VSUBS 0.00689f
C929 B.n712 VSUBS 0.00689f
C930 B.n713 VSUBS 0.00689f
C931 B.n714 VSUBS 0.00689f
C932 B.n715 VSUBS 0.00689f
C933 B.n716 VSUBS 0.00689f
C934 B.n717 VSUBS 0.00689f
C935 B.n718 VSUBS 0.00689f
C936 B.n719 VSUBS 0.00689f
C937 B.n720 VSUBS 0.00689f
C938 B.n721 VSUBS 0.00689f
C939 B.n722 VSUBS 0.00689f
C940 B.n723 VSUBS 0.00689f
C941 B.n724 VSUBS 0.00689f
C942 B.n725 VSUBS 0.00689f
C943 B.n726 VSUBS 0.00689f
C944 B.n727 VSUBS 0.00689f
C945 B.n728 VSUBS 0.00689f
C946 B.n729 VSUBS 0.00689f
C947 B.n730 VSUBS 0.00689f
C948 B.n731 VSUBS 0.00689f
C949 B.n732 VSUBS 0.00689f
C950 B.n733 VSUBS 0.00689f
C951 B.n734 VSUBS 0.00689f
C952 B.n735 VSUBS 0.00689f
C953 B.n736 VSUBS 0.00689f
C954 B.n737 VSUBS 0.00689f
C955 B.n738 VSUBS 0.00689f
C956 B.n739 VSUBS 0.00689f
C957 B.n740 VSUBS 0.00689f
C958 B.n741 VSUBS 0.00689f
C959 B.n742 VSUBS 0.00689f
C960 B.n743 VSUBS 0.00689f
C961 B.n744 VSUBS 0.00689f
C962 B.n745 VSUBS 0.00689f
C963 B.n746 VSUBS 0.00689f
C964 B.n747 VSUBS 0.00689f
C965 B.n748 VSUBS 0.00689f
C966 B.n749 VSUBS 0.00689f
C967 B.n750 VSUBS 0.00689f
C968 B.n751 VSUBS 0.00689f
C969 B.n752 VSUBS 0.00689f
C970 B.n753 VSUBS 0.00689f
C971 B.n754 VSUBS 0.00689f
C972 B.n755 VSUBS 0.015601f
.ends

