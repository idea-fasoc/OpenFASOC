* NGSPICE file created from diff_pair_sample_0940.ext - technology: sky130A

.subckt diff_pair_sample_0940 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=2.6202 ps=16.21 w=15.88 l=1.67
X1 VDD1.t3 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6202 pd=16.21 as=6.1932 ps=32.54 w=15.88 l=1.67
X2 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=2.6202 ps=16.21 w=15.88 l=1.67
X3 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6202 pd=16.21 as=6.1932 ps=32.54 w=15.88 l=1.67
X4 VTAIL.t5 VP.t2 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=2.6202 ps=16.21 w=15.88 l=1.67
X5 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=0 ps=0 w=15.88 l=1.67
X6 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6202 pd=16.21 as=6.1932 ps=32.54 w=15.88 l=1.67
X7 VDD1.t2 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6202 pd=16.21 as=6.1932 ps=32.54 w=15.88 l=1.67
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=0 ps=0 w=15.88 l=1.67
X9 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=2.6202 ps=16.21 w=15.88 l=1.67
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=0 ps=0 w=15.88 l=1.67
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1932 pd=32.54 as=0 ps=0 w=15.88 l=1.67
R0 VP.n2 VP.t2 263.668
R1 VP.n2 VP.t1 263.252
R2 VP.n9 VP.t3 229.167
R3 VP.n3 VP.t0 229.167
R4 VP.n8 VP.n0 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n1 161.3
R7 VP.n4 VP.n3 86.2628
R8 VP.n10 VP.n9 86.2628
R9 VP.n4 VP.n2 55.9727
R10 VP.n7 VP.n1 40.4106
R11 VP.n8 VP.n7 40.4106
R12 VP.n3 VP.n1 24.3439
R13 VP.n9 VP.n8 24.3439
R14 VP.n5 VP.n4 0.278398
R15 VP.n10 VP.n0 0.278398
R16 VP.n6 VP.n5 0.189894
R17 VP.n6 VP.n0 0.189894
R18 VP VP.n10 0.153422
R19 VDD1 VDD1.n1 107.013
R20 VDD1 VDD1.n0 63.9693
R21 VDD1.n0 VDD1.t0 1.24735
R22 VDD1.n0 VDD1.t3 1.24735
R23 VDD1.n1 VDD1.t1 1.24735
R24 VDD1.n1 VDD1.t2 1.24735
R25 VTAIL.n5 VTAIL.t5 48.4793
R26 VTAIL.n4 VTAIL.t1 48.4793
R27 VTAIL.n3 VTAIL.t3 48.4793
R28 VTAIL.n7 VTAIL.t0 48.4792
R29 VTAIL.n0 VTAIL.t2 48.4792
R30 VTAIL.n1 VTAIL.t4 48.4792
R31 VTAIL.n2 VTAIL.t7 48.4792
R32 VTAIL.n6 VTAIL.t6 48.4792
R33 VTAIL.n7 VTAIL.n6 27.7807
R34 VTAIL.n3 VTAIL.n2 27.7807
R35 VTAIL.n4 VTAIL.n3 1.72464
R36 VTAIL.n6 VTAIL.n5 1.72464
R37 VTAIL.n2 VTAIL.n1 1.72464
R38 VTAIL VTAIL.n0 0.920759
R39 VTAIL VTAIL.n7 0.804379
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 B.n796 B.n795 585
R43 B.n342 B.n107 585
R44 B.n341 B.n340 585
R45 B.n339 B.n338 585
R46 B.n337 B.n336 585
R47 B.n335 B.n334 585
R48 B.n333 B.n332 585
R49 B.n331 B.n330 585
R50 B.n329 B.n328 585
R51 B.n327 B.n326 585
R52 B.n325 B.n324 585
R53 B.n323 B.n322 585
R54 B.n321 B.n320 585
R55 B.n319 B.n318 585
R56 B.n317 B.n316 585
R57 B.n315 B.n314 585
R58 B.n313 B.n312 585
R59 B.n311 B.n310 585
R60 B.n309 B.n308 585
R61 B.n307 B.n306 585
R62 B.n305 B.n304 585
R63 B.n303 B.n302 585
R64 B.n301 B.n300 585
R65 B.n299 B.n298 585
R66 B.n297 B.n296 585
R67 B.n295 B.n294 585
R68 B.n293 B.n292 585
R69 B.n291 B.n290 585
R70 B.n289 B.n288 585
R71 B.n287 B.n286 585
R72 B.n285 B.n284 585
R73 B.n283 B.n282 585
R74 B.n281 B.n280 585
R75 B.n279 B.n278 585
R76 B.n277 B.n276 585
R77 B.n275 B.n274 585
R78 B.n273 B.n272 585
R79 B.n271 B.n270 585
R80 B.n269 B.n268 585
R81 B.n267 B.n266 585
R82 B.n265 B.n264 585
R83 B.n263 B.n262 585
R84 B.n261 B.n260 585
R85 B.n259 B.n258 585
R86 B.n257 B.n256 585
R87 B.n255 B.n254 585
R88 B.n253 B.n252 585
R89 B.n251 B.n250 585
R90 B.n249 B.n248 585
R91 B.n247 B.n246 585
R92 B.n245 B.n244 585
R93 B.n243 B.n242 585
R94 B.n241 B.n240 585
R95 B.n238 B.n237 585
R96 B.n236 B.n235 585
R97 B.n234 B.n233 585
R98 B.n232 B.n231 585
R99 B.n230 B.n229 585
R100 B.n228 B.n227 585
R101 B.n226 B.n225 585
R102 B.n224 B.n223 585
R103 B.n222 B.n221 585
R104 B.n220 B.n219 585
R105 B.n217 B.n216 585
R106 B.n215 B.n214 585
R107 B.n213 B.n212 585
R108 B.n211 B.n210 585
R109 B.n209 B.n208 585
R110 B.n207 B.n206 585
R111 B.n205 B.n204 585
R112 B.n203 B.n202 585
R113 B.n201 B.n200 585
R114 B.n199 B.n198 585
R115 B.n197 B.n196 585
R116 B.n195 B.n194 585
R117 B.n193 B.n192 585
R118 B.n191 B.n190 585
R119 B.n189 B.n188 585
R120 B.n187 B.n186 585
R121 B.n185 B.n184 585
R122 B.n183 B.n182 585
R123 B.n181 B.n180 585
R124 B.n179 B.n178 585
R125 B.n177 B.n176 585
R126 B.n175 B.n174 585
R127 B.n173 B.n172 585
R128 B.n171 B.n170 585
R129 B.n169 B.n168 585
R130 B.n167 B.n166 585
R131 B.n165 B.n164 585
R132 B.n163 B.n162 585
R133 B.n161 B.n160 585
R134 B.n159 B.n158 585
R135 B.n157 B.n156 585
R136 B.n155 B.n154 585
R137 B.n153 B.n152 585
R138 B.n151 B.n150 585
R139 B.n149 B.n148 585
R140 B.n147 B.n146 585
R141 B.n145 B.n144 585
R142 B.n143 B.n142 585
R143 B.n141 B.n140 585
R144 B.n139 B.n138 585
R145 B.n137 B.n136 585
R146 B.n135 B.n134 585
R147 B.n133 B.n132 585
R148 B.n131 B.n130 585
R149 B.n129 B.n128 585
R150 B.n127 B.n126 585
R151 B.n125 B.n124 585
R152 B.n123 B.n122 585
R153 B.n121 B.n120 585
R154 B.n119 B.n118 585
R155 B.n117 B.n116 585
R156 B.n115 B.n114 585
R157 B.n113 B.n112 585
R158 B.n794 B.n49 585
R159 B.n799 B.n49 585
R160 B.n793 B.n48 585
R161 B.n800 B.n48 585
R162 B.n792 B.n791 585
R163 B.n791 B.n44 585
R164 B.n790 B.n43 585
R165 B.n806 B.n43 585
R166 B.n789 B.n42 585
R167 B.n807 B.n42 585
R168 B.n788 B.n41 585
R169 B.n808 B.n41 585
R170 B.n787 B.n786 585
R171 B.n786 B.n37 585
R172 B.n785 B.n36 585
R173 B.n814 B.n36 585
R174 B.n784 B.n35 585
R175 B.n815 B.n35 585
R176 B.n783 B.n34 585
R177 B.n816 B.n34 585
R178 B.n782 B.n781 585
R179 B.n781 B.n30 585
R180 B.n780 B.n29 585
R181 B.n822 B.n29 585
R182 B.n779 B.n28 585
R183 B.n823 B.n28 585
R184 B.n778 B.n27 585
R185 B.n824 B.n27 585
R186 B.n777 B.n776 585
R187 B.n776 B.n23 585
R188 B.n775 B.n22 585
R189 B.n830 B.n22 585
R190 B.n774 B.n21 585
R191 B.n831 B.n21 585
R192 B.n773 B.n20 585
R193 B.n832 B.n20 585
R194 B.n772 B.n771 585
R195 B.n771 B.n16 585
R196 B.n770 B.n15 585
R197 B.n838 B.n15 585
R198 B.n769 B.n14 585
R199 B.n839 B.n14 585
R200 B.n768 B.n13 585
R201 B.n840 B.n13 585
R202 B.n767 B.n766 585
R203 B.n766 B.n12 585
R204 B.n765 B.n764 585
R205 B.n765 B.n8 585
R206 B.n763 B.n7 585
R207 B.n847 B.n7 585
R208 B.n762 B.n6 585
R209 B.n848 B.n6 585
R210 B.n761 B.n5 585
R211 B.n849 B.n5 585
R212 B.n760 B.n759 585
R213 B.n759 B.n4 585
R214 B.n758 B.n343 585
R215 B.n758 B.n757 585
R216 B.n748 B.n344 585
R217 B.n345 B.n344 585
R218 B.n750 B.n749 585
R219 B.n751 B.n750 585
R220 B.n747 B.n349 585
R221 B.n353 B.n349 585
R222 B.n746 B.n745 585
R223 B.n745 B.n744 585
R224 B.n351 B.n350 585
R225 B.n352 B.n351 585
R226 B.n737 B.n736 585
R227 B.n738 B.n737 585
R228 B.n735 B.n358 585
R229 B.n358 B.n357 585
R230 B.n734 B.n733 585
R231 B.n733 B.n732 585
R232 B.n360 B.n359 585
R233 B.n361 B.n360 585
R234 B.n725 B.n724 585
R235 B.n726 B.n725 585
R236 B.n723 B.n366 585
R237 B.n366 B.n365 585
R238 B.n722 B.n721 585
R239 B.n721 B.n720 585
R240 B.n368 B.n367 585
R241 B.n369 B.n368 585
R242 B.n713 B.n712 585
R243 B.n714 B.n713 585
R244 B.n711 B.n374 585
R245 B.n374 B.n373 585
R246 B.n710 B.n709 585
R247 B.n709 B.n708 585
R248 B.n376 B.n375 585
R249 B.n377 B.n376 585
R250 B.n701 B.n700 585
R251 B.n702 B.n701 585
R252 B.n699 B.n382 585
R253 B.n382 B.n381 585
R254 B.n698 B.n697 585
R255 B.n697 B.n696 585
R256 B.n384 B.n383 585
R257 B.n385 B.n384 585
R258 B.n689 B.n688 585
R259 B.n690 B.n689 585
R260 B.n687 B.n390 585
R261 B.n390 B.n389 585
R262 B.n682 B.n681 585
R263 B.n680 B.n450 585
R264 B.n679 B.n449 585
R265 B.n684 B.n449 585
R266 B.n678 B.n677 585
R267 B.n676 B.n675 585
R268 B.n674 B.n673 585
R269 B.n672 B.n671 585
R270 B.n670 B.n669 585
R271 B.n668 B.n667 585
R272 B.n666 B.n665 585
R273 B.n664 B.n663 585
R274 B.n662 B.n661 585
R275 B.n660 B.n659 585
R276 B.n658 B.n657 585
R277 B.n656 B.n655 585
R278 B.n654 B.n653 585
R279 B.n652 B.n651 585
R280 B.n650 B.n649 585
R281 B.n648 B.n647 585
R282 B.n646 B.n645 585
R283 B.n644 B.n643 585
R284 B.n642 B.n641 585
R285 B.n640 B.n639 585
R286 B.n638 B.n637 585
R287 B.n636 B.n635 585
R288 B.n634 B.n633 585
R289 B.n632 B.n631 585
R290 B.n630 B.n629 585
R291 B.n628 B.n627 585
R292 B.n626 B.n625 585
R293 B.n624 B.n623 585
R294 B.n622 B.n621 585
R295 B.n620 B.n619 585
R296 B.n618 B.n617 585
R297 B.n616 B.n615 585
R298 B.n614 B.n613 585
R299 B.n612 B.n611 585
R300 B.n610 B.n609 585
R301 B.n608 B.n607 585
R302 B.n606 B.n605 585
R303 B.n604 B.n603 585
R304 B.n602 B.n601 585
R305 B.n600 B.n599 585
R306 B.n598 B.n597 585
R307 B.n596 B.n595 585
R308 B.n594 B.n593 585
R309 B.n592 B.n591 585
R310 B.n590 B.n589 585
R311 B.n588 B.n587 585
R312 B.n586 B.n585 585
R313 B.n584 B.n583 585
R314 B.n582 B.n581 585
R315 B.n580 B.n579 585
R316 B.n578 B.n577 585
R317 B.n576 B.n575 585
R318 B.n574 B.n573 585
R319 B.n572 B.n571 585
R320 B.n570 B.n569 585
R321 B.n568 B.n567 585
R322 B.n566 B.n565 585
R323 B.n564 B.n563 585
R324 B.n562 B.n561 585
R325 B.n560 B.n559 585
R326 B.n558 B.n557 585
R327 B.n556 B.n555 585
R328 B.n554 B.n553 585
R329 B.n552 B.n551 585
R330 B.n550 B.n549 585
R331 B.n548 B.n547 585
R332 B.n546 B.n545 585
R333 B.n544 B.n543 585
R334 B.n542 B.n541 585
R335 B.n540 B.n539 585
R336 B.n538 B.n537 585
R337 B.n536 B.n535 585
R338 B.n534 B.n533 585
R339 B.n532 B.n531 585
R340 B.n530 B.n529 585
R341 B.n528 B.n527 585
R342 B.n526 B.n525 585
R343 B.n524 B.n523 585
R344 B.n522 B.n521 585
R345 B.n520 B.n519 585
R346 B.n518 B.n517 585
R347 B.n516 B.n515 585
R348 B.n514 B.n513 585
R349 B.n512 B.n511 585
R350 B.n510 B.n509 585
R351 B.n508 B.n507 585
R352 B.n506 B.n505 585
R353 B.n504 B.n503 585
R354 B.n502 B.n501 585
R355 B.n500 B.n499 585
R356 B.n498 B.n497 585
R357 B.n496 B.n495 585
R358 B.n494 B.n493 585
R359 B.n492 B.n491 585
R360 B.n490 B.n489 585
R361 B.n488 B.n487 585
R362 B.n486 B.n485 585
R363 B.n484 B.n483 585
R364 B.n482 B.n481 585
R365 B.n480 B.n479 585
R366 B.n478 B.n477 585
R367 B.n476 B.n475 585
R368 B.n474 B.n473 585
R369 B.n472 B.n471 585
R370 B.n470 B.n469 585
R371 B.n468 B.n467 585
R372 B.n466 B.n465 585
R373 B.n464 B.n463 585
R374 B.n462 B.n461 585
R375 B.n460 B.n459 585
R376 B.n458 B.n457 585
R377 B.n392 B.n391 585
R378 B.n686 B.n685 585
R379 B.n685 B.n684 585
R380 B.n388 B.n387 585
R381 B.n389 B.n388 585
R382 B.n692 B.n691 585
R383 B.n691 B.n690 585
R384 B.n693 B.n386 585
R385 B.n386 B.n385 585
R386 B.n695 B.n694 585
R387 B.n696 B.n695 585
R388 B.n380 B.n379 585
R389 B.n381 B.n380 585
R390 B.n704 B.n703 585
R391 B.n703 B.n702 585
R392 B.n705 B.n378 585
R393 B.n378 B.n377 585
R394 B.n707 B.n706 585
R395 B.n708 B.n707 585
R396 B.n372 B.n371 585
R397 B.n373 B.n372 585
R398 B.n716 B.n715 585
R399 B.n715 B.n714 585
R400 B.n717 B.n370 585
R401 B.n370 B.n369 585
R402 B.n719 B.n718 585
R403 B.n720 B.n719 585
R404 B.n364 B.n363 585
R405 B.n365 B.n364 585
R406 B.n728 B.n727 585
R407 B.n727 B.n726 585
R408 B.n729 B.n362 585
R409 B.n362 B.n361 585
R410 B.n731 B.n730 585
R411 B.n732 B.n731 585
R412 B.n356 B.n355 585
R413 B.n357 B.n356 585
R414 B.n740 B.n739 585
R415 B.n739 B.n738 585
R416 B.n741 B.n354 585
R417 B.n354 B.n352 585
R418 B.n743 B.n742 585
R419 B.n744 B.n743 585
R420 B.n348 B.n347 585
R421 B.n353 B.n348 585
R422 B.n753 B.n752 585
R423 B.n752 B.n751 585
R424 B.n754 B.n346 585
R425 B.n346 B.n345 585
R426 B.n756 B.n755 585
R427 B.n757 B.n756 585
R428 B.n3 B.n0 585
R429 B.n4 B.n3 585
R430 B.n846 B.n1 585
R431 B.n847 B.n846 585
R432 B.n845 B.n844 585
R433 B.n845 B.n8 585
R434 B.n843 B.n9 585
R435 B.n12 B.n9 585
R436 B.n842 B.n841 585
R437 B.n841 B.n840 585
R438 B.n11 B.n10 585
R439 B.n839 B.n11 585
R440 B.n837 B.n836 585
R441 B.n838 B.n837 585
R442 B.n835 B.n17 585
R443 B.n17 B.n16 585
R444 B.n834 B.n833 585
R445 B.n833 B.n832 585
R446 B.n19 B.n18 585
R447 B.n831 B.n19 585
R448 B.n829 B.n828 585
R449 B.n830 B.n829 585
R450 B.n827 B.n24 585
R451 B.n24 B.n23 585
R452 B.n826 B.n825 585
R453 B.n825 B.n824 585
R454 B.n26 B.n25 585
R455 B.n823 B.n26 585
R456 B.n821 B.n820 585
R457 B.n822 B.n821 585
R458 B.n819 B.n31 585
R459 B.n31 B.n30 585
R460 B.n818 B.n817 585
R461 B.n817 B.n816 585
R462 B.n33 B.n32 585
R463 B.n815 B.n33 585
R464 B.n813 B.n812 585
R465 B.n814 B.n813 585
R466 B.n811 B.n38 585
R467 B.n38 B.n37 585
R468 B.n810 B.n809 585
R469 B.n809 B.n808 585
R470 B.n40 B.n39 585
R471 B.n807 B.n40 585
R472 B.n805 B.n804 585
R473 B.n806 B.n805 585
R474 B.n803 B.n45 585
R475 B.n45 B.n44 585
R476 B.n802 B.n801 585
R477 B.n801 B.n800 585
R478 B.n47 B.n46 585
R479 B.n799 B.n47 585
R480 B.n850 B.n849 585
R481 B.n848 B.n2 585
R482 B.n112 B.n47 511.721
R483 B.n796 B.n49 511.721
R484 B.n685 B.n390 511.721
R485 B.n682 B.n388 511.721
R486 B.n108 B.t4 435.834
R487 B.n454 B.t12 435.834
R488 B.n110 B.t15 435.394
R489 B.n451 B.t8 435.394
R490 B.n798 B.n797 256.663
R491 B.n798 B.n106 256.663
R492 B.n798 B.n105 256.663
R493 B.n798 B.n104 256.663
R494 B.n798 B.n103 256.663
R495 B.n798 B.n102 256.663
R496 B.n798 B.n101 256.663
R497 B.n798 B.n100 256.663
R498 B.n798 B.n99 256.663
R499 B.n798 B.n98 256.663
R500 B.n798 B.n97 256.663
R501 B.n798 B.n96 256.663
R502 B.n798 B.n95 256.663
R503 B.n798 B.n94 256.663
R504 B.n798 B.n93 256.663
R505 B.n798 B.n92 256.663
R506 B.n798 B.n91 256.663
R507 B.n798 B.n90 256.663
R508 B.n798 B.n89 256.663
R509 B.n798 B.n88 256.663
R510 B.n798 B.n87 256.663
R511 B.n798 B.n86 256.663
R512 B.n798 B.n85 256.663
R513 B.n798 B.n84 256.663
R514 B.n798 B.n83 256.663
R515 B.n798 B.n82 256.663
R516 B.n798 B.n81 256.663
R517 B.n798 B.n80 256.663
R518 B.n798 B.n79 256.663
R519 B.n798 B.n78 256.663
R520 B.n798 B.n77 256.663
R521 B.n798 B.n76 256.663
R522 B.n798 B.n75 256.663
R523 B.n798 B.n74 256.663
R524 B.n798 B.n73 256.663
R525 B.n798 B.n72 256.663
R526 B.n798 B.n71 256.663
R527 B.n798 B.n70 256.663
R528 B.n798 B.n69 256.663
R529 B.n798 B.n68 256.663
R530 B.n798 B.n67 256.663
R531 B.n798 B.n66 256.663
R532 B.n798 B.n65 256.663
R533 B.n798 B.n64 256.663
R534 B.n798 B.n63 256.663
R535 B.n798 B.n62 256.663
R536 B.n798 B.n61 256.663
R537 B.n798 B.n60 256.663
R538 B.n798 B.n59 256.663
R539 B.n798 B.n58 256.663
R540 B.n798 B.n57 256.663
R541 B.n798 B.n56 256.663
R542 B.n798 B.n55 256.663
R543 B.n798 B.n54 256.663
R544 B.n798 B.n53 256.663
R545 B.n798 B.n52 256.663
R546 B.n798 B.n51 256.663
R547 B.n798 B.n50 256.663
R548 B.n684 B.n683 256.663
R549 B.n684 B.n393 256.663
R550 B.n684 B.n394 256.663
R551 B.n684 B.n395 256.663
R552 B.n684 B.n396 256.663
R553 B.n684 B.n397 256.663
R554 B.n684 B.n398 256.663
R555 B.n684 B.n399 256.663
R556 B.n684 B.n400 256.663
R557 B.n684 B.n401 256.663
R558 B.n684 B.n402 256.663
R559 B.n684 B.n403 256.663
R560 B.n684 B.n404 256.663
R561 B.n684 B.n405 256.663
R562 B.n684 B.n406 256.663
R563 B.n684 B.n407 256.663
R564 B.n684 B.n408 256.663
R565 B.n684 B.n409 256.663
R566 B.n684 B.n410 256.663
R567 B.n684 B.n411 256.663
R568 B.n684 B.n412 256.663
R569 B.n684 B.n413 256.663
R570 B.n684 B.n414 256.663
R571 B.n684 B.n415 256.663
R572 B.n684 B.n416 256.663
R573 B.n684 B.n417 256.663
R574 B.n684 B.n418 256.663
R575 B.n684 B.n419 256.663
R576 B.n684 B.n420 256.663
R577 B.n684 B.n421 256.663
R578 B.n684 B.n422 256.663
R579 B.n684 B.n423 256.663
R580 B.n684 B.n424 256.663
R581 B.n684 B.n425 256.663
R582 B.n684 B.n426 256.663
R583 B.n684 B.n427 256.663
R584 B.n684 B.n428 256.663
R585 B.n684 B.n429 256.663
R586 B.n684 B.n430 256.663
R587 B.n684 B.n431 256.663
R588 B.n684 B.n432 256.663
R589 B.n684 B.n433 256.663
R590 B.n684 B.n434 256.663
R591 B.n684 B.n435 256.663
R592 B.n684 B.n436 256.663
R593 B.n684 B.n437 256.663
R594 B.n684 B.n438 256.663
R595 B.n684 B.n439 256.663
R596 B.n684 B.n440 256.663
R597 B.n684 B.n441 256.663
R598 B.n684 B.n442 256.663
R599 B.n684 B.n443 256.663
R600 B.n684 B.n444 256.663
R601 B.n684 B.n445 256.663
R602 B.n684 B.n446 256.663
R603 B.n684 B.n447 256.663
R604 B.n684 B.n448 256.663
R605 B.n852 B.n851 256.663
R606 B.n116 B.n115 163.367
R607 B.n120 B.n119 163.367
R608 B.n124 B.n123 163.367
R609 B.n128 B.n127 163.367
R610 B.n132 B.n131 163.367
R611 B.n136 B.n135 163.367
R612 B.n140 B.n139 163.367
R613 B.n144 B.n143 163.367
R614 B.n148 B.n147 163.367
R615 B.n152 B.n151 163.367
R616 B.n156 B.n155 163.367
R617 B.n160 B.n159 163.367
R618 B.n164 B.n163 163.367
R619 B.n168 B.n167 163.367
R620 B.n172 B.n171 163.367
R621 B.n176 B.n175 163.367
R622 B.n180 B.n179 163.367
R623 B.n184 B.n183 163.367
R624 B.n188 B.n187 163.367
R625 B.n192 B.n191 163.367
R626 B.n196 B.n195 163.367
R627 B.n200 B.n199 163.367
R628 B.n204 B.n203 163.367
R629 B.n208 B.n207 163.367
R630 B.n212 B.n211 163.367
R631 B.n216 B.n215 163.367
R632 B.n221 B.n220 163.367
R633 B.n225 B.n224 163.367
R634 B.n229 B.n228 163.367
R635 B.n233 B.n232 163.367
R636 B.n237 B.n236 163.367
R637 B.n242 B.n241 163.367
R638 B.n246 B.n245 163.367
R639 B.n250 B.n249 163.367
R640 B.n254 B.n253 163.367
R641 B.n258 B.n257 163.367
R642 B.n262 B.n261 163.367
R643 B.n266 B.n265 163.367
R644 B.n270 B.n269 163.367
R645 B.n274 B.n273 163.367
R646 B.n278 B.n277 163.367
R647 B.n282 B.n281 163.367
R648 B.n286 B.n285 163.367
R649 B.n290 B.n289 163.367
R650 B.n294 B.n293 163.367
R651 B.n298 B.n297 163.367
R652 B.n302 B.n301 163.367
R653 B.n306 B.n305 163.367
R654 B.n310 B.n309 163.367
R655 B.n314 B.n313 163.367
R656 B.n318 B.n317 163.367
R657 B.n322 B.n321 163.367
R658 B.n326 B.n325 163.367
R659 B.n330 B.n329 163.367
R660 B.n334 B.n333 163.367
R661 B.n338 B.n337 163.367
R662 B.n340 B.n107 163.367
R663 B.n689 B.n390 163.367
R664 B.n689 B.n384 163.367
R665 B.n697 B.n384 163.367
R666 B.n697 B.n382 163.367
R667 B.n701 B.n382 163.367
R668 B.n701 B.n376 163.367
R669 B.n709 B.n376 163.367
R670 B.n709 B.n374 163.367
R671 B.n713 B.n374 163.367
R672 B.n713 B.n368 163.367
R673 B.n721 B.n368 163.367
R674 B.n721 B.n366 163.367
R675 B.n725 B.n366 163.367
R676 B.n725 B.n360 163.367
R677 B.n733 B.n360 163.367
R678 B.n733 B.n358 163.367
R679 B.n737 B.n358 163.367
R680 B.n737 B.n351 163.367
R681 B.n745 B.n351 163.367
R682 B.n745 B.n349 163.367
R683 B.n750 B.n349 163.367
R684 B.n750 B.n344 163.367
R685 B.n758 B.n344 163.367
R686 B.n759 B.n758 163.367
R687 B.n759 B.n5 163.367
R688 B.n6 B.n5 163.367
R689 B.n7 B.n6 163.367
R690 B.n765 B.n7 163.367
R691 B.n766 B.n765 163.367
R692 B.n766 B.n13 163.367
R693 B.n14 B.n13 163.367
R694 B.n15 B.n14 163.367
R695 B.n771 B.n15 163.367
R696 B.n771 B.n20 163.367
R697 B.n21 B.n20 163.367
R698 B.n22 B.n21 163.367
R699 B.n776 B.n22 163.367
R700 B.n776 B.n27 163.367
R701 B.n28 B.n27 163.367
R702 B.n29 B.n28 163.367
R703 B.n781 B.n29 163.367
R704 B.n781 B.n34 163.367
R705 B.n35 B.n34 163.367
R706 B.n36 B.n35 163.367
R707 B.n786 B.n36 163.367
R708 B.n786 B.n41 163.367
R709 B.n42 B.n41 163.367
R710 B.n43 B.n42 163.367
R711 B.n791 B.n43 163.367
R712 B.n791 B.n48 163.367
R713 B.n49 B.n48 163.367
R714 B.n450 B.n449 163.367
R715 B.n677 B.n449 163.367
R716 B.n675 B.n674 163.367
R717 B.n671 B.n670 163.367
R718 B.n667 B.n666 163.367
R719 B.n663 B.n662 163.367
R720 B.n659 B.n658 163.367
R721 B.n655 B.n654 163.367
R722 B.n651 B.n650 163.367
R723 B.n647 B.n646 163.367
R724 B.n643 B.n642 163.367
R725 B.n639 B.n638 163.367
R726 B.n635 B.n634 163.367
R727 B.n631 B.n630 163.367
R728 B.n627 B.n626 163.367
R729 B.n623 B.n622 163.367
R730 B.n619 B.n618 163.367
R731 B.n615 B.n614 163.367
R732 B.n611 B.n610 163.367
R733 B.n607 B.n606 163.367
R734 B.n603 B.n602 163.367
R735 B.n599 B.n598 163.367
R736 B.n595 B.n594 163.367
R737 B.n591 B.n590 163.367
R738 B.n587 B.n586 163.367
R739 B.n583 B.n582 163.367
R740 B.n579 B.n578 163.367
R741 B.n575 B.n574 163.367
R742 B.n571 B.n570 163.367
R743 B.n567 B.n566 163.367
R744 B.n563 B.n562 163.367
R745 B.n559 B.n558 163.367
R746 B.n555 B.n554 163.367
R747 B.n551 B.n550 163.367
R748 B.n547 B.n546 163.367
R749 B.n543 B.n542 163.367
R750 B.n539 B.n538 163.367
R751 B.n535 B.n534 163.367
R752 B.n531 B.n530 163.367
R753 B.n527 B.n526 163.367
R754 B.n523 B.n522 163.367
R755 B.n519 B.n518 163.367
R756 B.n515 B.n514 163.367
R757 B.n511 B.n510 163.367
R758 B.n507 B.n506 163.367
R759 B.n503 B.n502 163.367
R760 B.n499 B.n498 163.367
R761 B.n495 B.n494 163.367
R762 B.n491 B.n490 163.367
R763 B.n487 B.n486 163.367
R764 B.n483 B.n482 163.367
R765 B.n479 B.n478 163.367
R766 B.n475 B.n474 163.367
R767 B.n471 B.n470 163.367
R768 B.n467 B.n466 163.367
R769 B.n463 B.n462 163.367
R770 B.n459 B.n458 163.367
R771 B.n685 B.n392 163.367
R772 B.n691 B.n388 163.367
R773 B.n691 B.n386 163.367
R774 B.n695 B.n386 163.367
R775 B.n695 B.n380 163.367
R776 B.n703 B.n380 163.367
R777 B.n703 B.n378 163.367
R778 B.n707 B.n378 163.367
R779 B.n707 B.n372 163.367
R780 B.n715 B.n372 163.367
R781 B.n715 B.n370 163.367
R782 B.n719 B.n370 163.367
R783 B.n719 B.n364 163.367
R784 B.n727 B.n364 163.367
R785 B.n727 B.n362 163.367
R786 B.n731 B.n362 163.367
R787 B.n731 B.n356 163.367
R788 B.n739 B.n356 163.367
R789 B.n739 B.n354 163.367
R790 B.n743 B.n354 163.367
R791 B.n743 B.n348 163.367
R792 B.n752 B.n348 163.367
R793 B.n752 B.n346 163.367
R794 B.n756 B.n346 163.367
R795 B.n756 B.n3 163.367
R796 B.n850 B.n3 163.367
R797 B.n846 B.n2 163.367
R798 B.n846 B.n845 163.367
R799 B.n845 B.n9 163.367
R800 B.n841 B.n9 163.367
R801 B.n841 B.n11 163.367
R802 B.n837 B.n11 163.367
R803 B.n837 B.n17 163.367
R804 B.n833 B.n17 163.367
R805 B.n833 B.n19 163.367
R806 B.n829 B.n19 163.367
R807 B.n829 B.n24 163.367
R808 B.n825 B.n24 163.367
R809 B.n825 B.n26 163.367
R810 B.n821 B.n26 163.367
R811 B.n821 B.n31 163.367
R812 B.n817 B.n31 163.367
R813 B.n817 B.n33 163.367
R814 B.n813 B.n33 163.367
R815 B.n813 B.n38 163.367
R816 B.n809 B.n38 163.367
R817 B.n809 B.n40 163.367
R818 B.n805 B.n40 163.367
R819 B.n805 B.n45 163.367
R820 B.n801 B.n45 163.367
R821 B.n801 B.n47 163.367
R822 B.n108 B.t6 111.028
R823 B.n454 B.t14 111.028
R824 B.n110 B.t16 111.007
R825 B.n451 B.t11 111.007
R826 B.n684 B.n389 73.3165
R827 B.n799 B.n798 73.3165
R828 B.n109 B.t7 72.2407
R829 B.n455 B.t13 72.2407
R830 B.n111 B.t17 72.22
R831 B.n452 B.t10 72.22
R832 B.n112 B.n50 71.676
R833 B.n116 B.n51 71.676
R834 B.n120 B.n52 71.676
R835 B.n124 B.n53 71.676
R836 B.n128 B.n54 71.676
R837 B.n132 B.n55 71.676
R838 B.n136 B.n56 71.676
R839 B.n140 B.n57 71.676
R840 B.n144 B.n58 71.676
R841 B.n148 B.n59 71.676
R842 B.n152 B.n60 71.676
R843 B.n156 B.n61 71.676
R844 B.n160 B.n62 71.676
R845 B.n164 B.n63 71.676
R846 B.n168 B.n64 71.676
R847 B.n172 B.n65 71.676
R848 B.n176 B.n66 71.676
R849 B.n180 B.n67 71.676
R850 B.n184 B.n68 71.676
R851 B.n188 B.n69 71.676
R852 B.n192 B.n70 71.676
R853 B.n196 B.n71 71.676
R854 B.n200 B.n72 71.676
R855 B.n204 B.n73 71.676
R856 B.n208 B.n74 71.676
R857 B.n212 B.n75 71.676
R858 B.n216 B.n76 71.676
R859 B.n221 B.n77 71.676
R860 B.n225 B.n78 71.676
R861 B.n229 B.n79 71.676
R862 B.n233 B.n80 71.676
R863 B.n237 B.n81 71.676
R864 B.n242 B.n82 71.676
R865 B.n246 B.n83 71.676
R866 B.n250 B.n84 71.676
R867 B.n254 B.n85 71.676
R868 B.n258 B.n86 71.676
R869 B.n262 B.n87 71.676
R870 B.n266 B.n88 71.676
R871 B.n270 B.n89 71.676
R872 B.n274 B.n90 71.676
R873 B.n278 B.n91 71.676
R874 B.n282 B.n92 71.676
R875 B.n286 B.n93 71.676
R876 B.n290 B.n94 71.676
R877 B.n294 B.n95 71.676
R878 B.n298 B.n96 71.676
R879 B.n302 B.n97 71.676
R880 B.n306 B.n98 71.676
R881 B.n310 B.n99 71.676
R882 B.n314 B.n100 71.676
R883 B.n318 B.n101 71.676
R884 B.n322 B.n102 71.676
R885 B.n326 B.n103 71.676
R886 B.n330 B.n104 71.676
R887 B.n334 B.n105 71.676
R888 B.n338 B.n106 71.676
R889 B.n797 B.n107 71.676
R890 B.n797 B.n796 71.676
R891 B.n340 B.n106 71.676
R892 B.n337 B.n105 71.676
R893 B.n333 B.n104 71.676
R894 B.n329 B.n103 71.676
R895 B.n325 B.n102 71.676
R896 B.n321 B.n101 71.676
R897 B.n317 B.n100 71.676
R898 B.n313 B.n99 71.676
R899 B.n309 B.n98 71.676
R900 B.n305 B.n97 71.676
R901 B.n301 B.n96 71.676
R902 B.n297 B.n95 71.676
R903 B.n293 B.n94 71.676
R904 B.n289 B.n93 71.676
R905 B.n285 B.n92 71.676
R906 B.n281 B.n91 71.676
R907 B.n277 B.n90 71.676
R908 B.n273 B.n89 71.676
R909 B.n269 B.n88 71.676
R910 B.n265 B.n87 71.676
R911 B.n261 B.n86 71.676
R912 B.n257 B.n85 71.676
R913 B.n253 B.n84 71.676
R914 B.n249 B.n83 71.676
R915 B.n245 B.n82 71.676
R916 B.n241 B.n81 71.676
R917 B.n236 B.n80 71.676
R918 B.n232 B.n79 71.676
R919 B.n228 B.n78 71.676
R920 B.n224 B.n77 71.676
R921 B.n220 B.n76 71.676
R922 B.n215 B.n75 71.676
R923 B.n211 B.n74 71.676
R924 B.n207 B.n73 71.676
R925 B.n203 B.n72 71.676
R926 B.n199 B.n71 71.676
R927 B.n195 B.n70 71.676
R928 B.n191 B.n69 71.676
R929 B.n187 B.n68 71.676
R930 B.n183 B.n67 71.676
R931 B.n179 B.n66 71.676
R932 B.n175 B.n65 71.676
R933 B.n171 B.n64 71.676
R934 B.n167 B.n63 71.676
R935 B.n163 B.n62 71.676
R936 B.n159 B.n61 71.676
R937 B.n155 B.n60 71.676
R938 B.n151 B.n59 71.676
R939 B.n147 B.n58 71.676
R940 B.n143 B.n57 71.676
R941 B.n139 B.n56 71.676
R942 B.n135 B.n55 71.676
R943 B.n131 B.n54 71.676
R944 B.n127 B.n53 71.676
R945 B.n123 B.n52 71.676
R946 B.n119 B.n51 71.676
R947 B.n115 B.n50 71.676
R948 B.n683 B.n682 71.676
R949 B.n677 B.n393 71.676
R950 B.n674 B.n394 71.676
R951 B.n670 B.n395 71.676
R952 B.n666 B.n396 71.676
R953 B.n662 B.n397 71.676
R954 B.n658 B.n398 71.676
R955 B.n654 B.n399 71.676
R956 B.n650 B.n400 71.676
R957 B.n646 B.n401 71.676
R958 B.n642 B.n402 71.676
R959 B.n638 B.n403 71.676
R960 B.n634 B.n404 71.676
R961 B.n630 B.n405 71.676
R962 B.n626 B.n406 71.676
R963 B.n622 B.n407 71.676
R964 B.n618 B.n408 71.676
R965 B.n614 B.n409 71.676
R966 B.n610 B.n410 71.676
R967 B.n606 B.n411 71.676
R968 B.n602 B.n412 71.676
R969 B.n598 B.n413 71.676
R970 B.n594 B.n414 71.676
R971 B.n590 B.n415 71.676
R972 B.n586 B.n416 71.676
R973 B.n582 B.n417 71.676
R974 B.n578 B.n418 71.676
R975 B.n574 B.n419 71.676
R976 B.n570 B.n420 71.676
R977 B.n566 B.n421 71.676
R978 B.n562 B.n422 71.676
R979 B.n558 B.n423 71.676
R980 B.n554 B.n424 71.676
R981 B.n550 B.n425 71.676
R982 B.n546 B.n426 71.676
R983 B.n542 B.n427 71.676
R984 B.n538 B.n428 71.676
R985 B.n534 B.n429 71.676
R986 B.n530 B.n430 71.676
R987 B.n526 B.n431 71.676
R988 B.n522 B.n432 71.676
R989 B.n518 B.n433 71.676
R990 B.n514 B.n434 71.676
R991 B.n510 B.n435 71.676
R992 B.n506 B.n436 71.676
R993 B.n502 B.n437 71.676
R994 B.n498 B.n438 71.676
R995 B.n494 B.n439 71.676
R996 B.n490 B.n440 71.676
R997 B.n486 B.n441 71.676
R998 B.n482 B.n442 71.676
R999 B.n478 B.n443 71.676
R1000 B.n474 B.n444 71.676
R1001 B.n470 B.n445 71.676
R1002 B.n466 B.n446 71.676
R1003 B.n462 B.n447 71.676
R1004 B.n458 B.n448 71.676
R1005 B.n683 B.n450 71.676
R1006 B.n675 B.n393 71.676
R1007 B.n671 B.n394 71.676
R1008 B.n667 B.n395 71.676
R1009 B.n663 B.n396 71.676
R1010 B.n659 B.n397 71.676
R1011 B.n655 B.n398 71.676
R1012 B.n651 B.n399 71.676
R1013 B.n647 B.n400 71.676
R1014 B.n643 B.n401 71.676
R1015 B.n639 B.n402 71.676
R1016 B.n635 B.n403 71.676
R1017 B.n631 B.n404 71.676
R1018 B.n627 B.n405 71.676
R1019 B.n623 B.n406 71.676
R1020 B.n619 B.n407 71.676
R1021 B.n615 B.n408 71.676
R1022 B.n611 B.n409 71.676
R1023 B.n607 B.n410 71.676
R1024 B.n603 B.n411 71.676
R1025 B.n599 B.n412 71.676
R1026 B.n595 B.n413 71.676
R1027 B.n591 B.n414 71.676
R1028 B.n587 B.n415 71.676
R1029 B.n583 B.n416 71.676
R1030 B.n579 B.n417 71.676
R1031 B.n575 B.n418 71.676
R1032 B.n571 B.n419 71.676
R1033 B.n567 B.n420 71.676
R1034 B.n563 B.n421 71.676
R1035 B.n559 B.n422 71.676
R1036 B.n555 B.n423 71.676
R1037 B.n551 B.n424 71.676
R1038 B.n547 B.n425 71.676
R1039 B.n543 B.n426 71.676
R1040 B.n539 B.n427 71.676
R1041 B.n535 B.n428 71.676
R1042 B.n531 B.n429 71.676
R1043 B.n527 B.n430 71.676
R1044 B.n523 B.n431 71.676
R1045 B.n519 B.n432 71.676
R1046 B.n515 B.n433 71.676
R1047 B.n511 B.n434 71.676
R1048 B.n507 B.n435 71.676
R1049 B.n503 B.n436 71.676
R1050 B.n499 B.n437 71.676
R1051 B.n495 B.n438 71.676
R1052 B.n491 B.n439 71.676
R1053 B.n487 B.n440 71.676
R1054 B.n483 B.n441 71.676
R1055 B.n479 B.n442 71.676
R1056 B.n475 B.n443 71.676
R1057 B.n471 B.n444 71.676
R1058 B.n467 B.n445 71.676
R1059 B.n463 B.n446 71.676
R1060 B.n459 B.n447 71.676
R1061 B.n448 B.n392 71.676
R1062 B.n851 B.n850 71.676
R1063 B.n851 B.n2 71.676
R1064 B.n218 B.n111 59.5399
R1065 B.n239 B.n109 59.5399
R1066 B.n456 B.n455 59.5399
R1067 B.n453 B.n452 59.5399
R1068 B.n111 B.n110 38.7884
R1069 B.n109 B.n108 38.7884
R1070 B.n455 B.n454 38.7884
R1071 B.n452 B.n451 38.7884
R1072 B.n690 B.n389 35.3586
R1073 B.n690 B.n385 35.3586
R1074 B.n696 B.n385 35.3586
R1075 B.n696 B.n381 35.3586
R1076 B.n702 B.n381 35.3586
R1077 B.n708 B.n377 35.3586
R1078 B.n708 B.n373 35.3586
R1079 B.n714 B.n373 35.3586
R1080 B.n714 B.n369 35.3586
R1081 B.n720 B.n369 35.3586
R1082 B.n720 B.n365 35.3586
R1083 B.n726 B.n365 35.3586
R1084 B.n726 B.n361 35.3586
R1085 B.n732 B.n361 35.3586
R1086 B.n738 B.n357 35.3586
R1087 B.n738 B.n352 35.3586
R1088 B.n744 B.n352 35.3586
R1089 B.n744 B.n353 35.3586
R1090 B.n751 B.n345 35.3586
R1091 B.n757 B.n345 35.3586
R1092 B.n757 B.n4 35.3586
R1093 B.n849 B.n4 35.3586
R1094 B.n849 B.n848 35.3586
R1095 B.n848 B.n847 35.3586
R1096 B.n847 B.n8 35.3586
R1097 B.n12 B.n8 35.3586
R1098 B.n840 B.n12 35.3586
R1099 B.n839 B.n838 35.3586
R1100 B.n838 B.n16 35.3586
R1101 B.n832 B.n16 35.3586
R1102 B.n832 B.n831 35.3586
R1103 B.n830 B.n23 35.3586
R1104 B.n824 B.n23 35.3586
R1105 B.n824 B.n823 35.3586
R1106 B.n823 B.n822 35.3586
R1107 B.n822 B.n30 35.3586
R1108 B.n816 B.n30 35.3586
R1109 B.n816 B.n815 35.3586
R1110 B.n815 B.n814 35.3586
R1111 B.n814 B.n37 35.3586
R1112 B.n808 B.n807 35.3586
R1113 B.n807 B.n806 35.3586
R1114 B.n806 B.n44 35.3586
R1115 B.n800 B.n44 35.3586
R1116 B.n800 B.n799 35.3586
R1117 B.n702 B.t9 34.8386
R1118 B.n808 B.t5 34.8386
R1119 B.n353 B.t1 33.7987
R1120 B.t2 B.n839 33.7987
R1121 B.n681 B.n387 33.2493
R1122 B.n687 B.n686 33.2493
R1123 B.n795 B.n794 33.2493
R1124 B.n113 B.n46 33.2493
R1125 B.t3 B.n357 32.7587
R1126 B.n831 B.t0 32.7587
R1127 B B.n852 18.0485
R1128 B.n692 B.n387 10.6151
R1129 B.n693 B.n692 10.6151
R1130 B.n694 B.n693 10.6151
R1131 B.n694 B.n379 10.6151
R1132 B.n704 B.n379 10.6151
R1133 B.n705 B.n704 10.6151
R1134 B.n706 B.n705 10.6151
R1135 B.n706 B.n371 10.6151
R1136 B.n716 B.n371 10.6151
R1137 B.n717 B.n716 10.6151
R1138 B.n718 B.n717 10.6151
R1139 B.n718 B.n363 10.6151
R1140 B.n728 B.n363 10.6151
R1141 B.n729 B.n728 10.6151
R1142 B.n730 B.n729 10.6151
R1143 B.n730 B.n355 10.6151
R1144 B.n740 B.n355 10.6151
R1145 B.n741 B.n740 10.6151
R1146 B.n742 B.n741 10.6151
R1147 B.n742 B.n347 10.6151
R1148 B.n753 B.n347 10.6151
R1149 B.n754 B.n753 10.6151
R1150 B.n755 B.n754 10.6151
R1151 B.n755 B.n0 10.6151
R1152 B.n681 B.n680 10.6151
R1153 B.n680 B.n679 10.6151
R1154 B.n679 B.n678 10.6151
R1155 B.n678 B.n676 10.6151
R1156 B.n676 B.n673 10.6151
R1157 B.n673 B.n672 10.6151
R1158 B.n672 B.n669 10.6151
R1159 B.n669 B.n668 10.6151
R1160 B.n668 B.n665 10.6151
R1161 B.n665 B.n664 10.6151
R1162 B.n664 B.n661 10.6151
R1163 B.n661 B.n660 10.6151
R1164 B.n660 B.n657 10.6151
R1165 B.n657 B.n656 10.6151
R1166 B.n656 B.n653 10.6151
R1167 B.n653 B.n652 10.6151
R1168 B.n652 B.n649 10.6151
R1169 B.n649 B.n648 10.6151
R1170 B.n648 B.n645 10.6151
R1171 B.n645 B.n644 10.6151
R1172 B.n644 B.n641 10.6151
R1173 B.n641 B.n640 10.6151
R1174 B.n640 B.n637 10.6151
R1175 B.n637 B.n636 10.6151
R1176 B.n636 B.n633 10.6151
R1177 B.n633 B.n632 10.6151
R1178 B.n632 B.n629 10.6151
R1179 B.n629 B.n628 10.6151
R1180 B.n628 B.n625 10.6151
R1181 B.n625 B.n624 10.6151
R1182 B.n624 B.n621 10.6151
R1183 B.n621 B.n620 10.6151
R1184 B.n620 B.n617 10.6151
R1185 B.n617 B.n616 10.6151
R1186 B.n616 B.n613 10.6151
R1187 B.n613 B.n612 10.6151
R1188 B.n612 B.n609 10.6151
R1189 B.n609 B.n608 10.6151
R1190 B.n608 B.n605 10.6151
R1191 B.n605 B.n604 10.6151
R1192 B.n604 B.n601 10.6151
R1193 B.n601 B.n600 10.6151
R1194 B.n600 B.n597 10.6151
R1195 B.n597 B.n596 10.6151
R1196 B.n596 B.n593 10.6151
R1197 B.n593 B.n592 10.6151
R1198 B.n592 B.n589 10.6151
R1199 B.n589 B.n588 10.6151
R1200 B.n588 B.n585 10.6151
R1201 B.n585 B.n584 10.6151
R1202 B.n584 B.n581 10.6151
R1203 B.n581 B.n580 10.6151
R1204 B.n577 B.n576 10.6151
R1205 B.n576 B.n573 10.6151
R1206 B.n573 B.n572 10.6151
R1207 B.n572 B.n569 10.6151
R1208 B.n569 B.n568 10.6151
R1209 B.n568 B.n565 10.6151
R1210 B.n565 B.n564 10.6151
R1211 B.n564 B.n561 10.6151
R1212 B.n561 B.n560 10.6151
R1213 B.n557 B.n556 10.6151
R1214 B.n556 B.n553 10.6151
R1215 B.n553 B.n552 10.6151
R1216 B.n552 B.n549 10.6151
R1217 B.n549 B.n548 10.6151
R1218 B.n548 B.n545 10.6151
R1219 B.n545 B.n544 10.6151
R1220 B.n544 B.n541 10.6151
R1221 B.n541 B.n540 10.6151
R1222 B.n540 B.n537 10.6151
R1223 B.n537 B.n536 10.6151
R1224 B.n536 B.n533 10.6151
R1225 B.n533 B.n532 10.6151
R1226 B.n532 B.n529 10.6151
R1227 B.n529 B.n528 10.6151
R1228 B.n528 B.n525 10.6151
R1229 B.n525 B.n524 10.6151
R1230 B.n524 B.n521 10.6151
R1231 B.n521 B.n520 10.6151
R1232 B.n520 B.n517 10.6151
R1233 B.n517 B.n516 10.6151
R1234 B.n516 B.n513 10.6151
R1235 B.n513 B.n512 10.6151
R1236 B.n512 B.n509 10.6151
R1237 B.n509 B.n508 10.6151
R1238 B.n508 B.n505 10.6151
R1239 B.n505 B.n504 10.6151
R1240 B.n504 B.n501 10.6151
R1241 B.n501 B.n500 10.6151
R1242 B.n500 B.n497 10.6151
R1243 B.n497 B.n496 10.6151
R1244 B.n496 B.n493 10.6151
R1245 B.n493 B.n492 10.6151
R1246 B.n492 B.n489 10.6151
R1247 B.n489 B.n488 10.6151
R1248 B.n488 B.n485 10.6151
R1249 B.n485 B.n484 10.6151
R1250 B.n484 B.n481 10.6151
R1251 B.n481 B.n480 10.6151
R1252 B.n480 B.n477 10.6151
R1253 B.n477 B.n476 10.6151
R1254 B.n476 B.n473 10.6151
R1255 B.n473 B.n472 10.6151
R1256 B.n472 B.n469 10.6151
R1257 B.n469 B.n468 10.6151
R1258 B.n468 B.n465 10.6151
R1259 B.n465 B.n464 10.6151
R1260 B.n464 B.n461 10.6151
R1261 B.n461 B.n460 10.6151
R1262 B.n460 B.n457 10.6151
R1263 B.n457 B.n391 10.6151
R1264 B.n686 B.n391 10.6151
R1265 B.n688 B.n687 10.6151
R1266 B.n688 B.n383 10.6151
R1267 B.n698 B.n383 10.6151
R1268 B.n699 B.n698 10.6151
R1269 B.n700 B.n699 10.6151
R1270 B.n700 B.n375 10.6151
R1271 B.n710 B.n375 10.6151
R1272 B.n711 B.n710 10.6151
R1273 B.n712 B.n711 10.6151
R1274 B.n712 B.n367 10.6151
R1275 B.n722 B.n367 10.6151
R1276 B.n723 B.n722 10.6151
R1277 B.n724 B.n723 10.6151
R1278 B.n724 B.n359 10.6151
R1279 B.n734 B.n359 10.6151
R1280 B.n735 B.n734 10.6151
R1281 B.n736 B.n735 10.6151
R1282 B.n736 B.n350 10.6151
R1283 B.n746 B.n350 10.6151
R1284 B.n747 B.n746 10.6151
R1285 B.n749 B.n747 10.6151
R1286 B.n749 B.n748 10.6151
R1287 B.n748 B.n343 10.6151
R1288 B.n760 B.n343 10.6151
R1289 B.n761 B.n760 10.6151
R1290 B.n762 B.n761 10.6151
R1291 B.n763 B.n762 10.6151
R1292 B.n764 B.n763 10.6151
R1293 B.n767 B.n764 10.6151
R1294 B.n768 B.n767 10.6151
R1295 B.n769 B.n768 10.6151
R1296 B.n770 B.n769 10.6151
R1297 B.n772 B.n770 10.6151
R1298 B.n773 B.n772 10.6151
R1299 B.n774 B.n773 10.6151
R1300 B.n775 B.n774 10.6151
R1301 B.n777 B.n775 10.6151
R1302 B.n778 B.n777 10.6151
R1303 B.n779 B.n778 10.6151
R1304 B.n780 B.n779 10.6151
R1305 B.n782 B.n780 10.6151
R1306 B.n783 B.n782 10.6151
R1307 B.n784 B.n783 10.6151
R1308 B.n785 B.n784 10.6151
R1309 B.n787 B.n785 10.6151
R1310 B.n788 B.n787 10.6151
R1311 B.n789 B.n788 10.6151
R1312 B.n790 B.n789 10.6151
R1313 B.n792 B.n790 10.6151
R1314 B.n793 B.n792 10.6151
R1315 B.n794 B.n793 10.6151
R1316 B.n844 B.n1 10.6151
R1317 B.n844 B.n843 10.6151
R1318 B.n843 B.n842 10.6151
R1319 B.n842 B.n10 10.6151
R1320 B.n836 B.n10 10.6151
R1321 B.n836 B.n835 10.6151
R1322 B.n835 B.n834 10.6151
R1323 B.n834 B.n18 10.6151
R1324 B.n828 B.n18 10.6151
R1325 B.n828 B.n827 10.6151
R1326 B.n827 B.n826 10.6151
R1327 B.n826 B.n25 10.6151
R1328 B.n820 B.n25 10.6151
R1329 B.n820 B.n819 10.6151
R1330 B.n819 B.n818 10.6151
R1331 B.n818 B.n32 10.6151
R1332 B.n812 B.n32 10.6151
R1333 B.n812 B.n811 10.6151
R1334 B.n811 B.n810 10.6151
R1335 B.n810 B.n39 10.6151
R1336 B.n804 B.n39 10.6151
R1337 B.n804 B.n803 10.6151
R1338 B.n803 B.n802 10.6151
R1339 B.n802 B.n46 10.6151
R1340 B.n114 B.n113 10.6151
R1341 B.n117 B.n114 10.6151
R1342 B.n118 B.n117 10.6151
R1343 B.n121 B.n118 10.6151
R1344 B.n122 B.n121 10.6151
R1345 B.n125 B.n122 10.6151
R1346 B.n126 B.n125 10.6151
R1347 B.n129 B.n126 10.6151
R1348 B.n130 B.n129 10.6151
R1349 B.n133 B.n130 10.6151
R1350 B.n134 B.n133 10.6151
R1351 B.n137 B.n134 10.6151
R1352 B.n138 B.n137 10.6151
R1353 B.n141 B.n138 10.6151
R1354 B.n142 B.n141 10.6151
R1355 B.n145 B.n142 10.6151
R1356 B.n146 B.n145 10.6151
R1357 B.n149 B.n146 10.6151
R1358 B.n150 B.n149 10.6151
R1359 B.n153 B.n150 10.6151
R1360 B.n154 B.n153 10.6151
R1361 B.n157 B.n154 10.6151
R1362 B.n158 B.n157 10.6151
R1363 B.n161 B.n158 10.6151
R1364 B.n162 B.n161 10.6151
R1365 B.n165 B.n162 10.6151
R1366 B.n166 B.n165 10.6151
R1367 B.n169 B.n166 10.6151
R1368 B.n170 B.n169 10.6151
R1369 B.n173 B.n170 10.6151
R1370 B.n174 B.n173 10.6151
R1371 B.n177 B.n174 10.6151
R1372 B.n178 B.n177 10.6151
R1373 B.n181 B.n178 10.6151
R1374 B.n182 B.n181 10.6151
R1375 B.n185 B.n182 10.6151
R1376 B.n186 B.n185 10.6151
R1377 B.n189 B.n186 10.6151
R1378 B.n190 B.n189 10.6151
R1379 B.n193 B.n190 10.6151
R1380 B.n194 B.n193 10.6151
R1381 B.n197 B.n194 10.6151
R1382 B.n198 B.n197 10.6151
R1383 B.n201 B.n198 10.6151
R1384 B.n202 B.n201 10.6151
R1385 B.n205 B.n202 10.6151
R1386 B.n206 B.n205 10.6151
R1387 B.n209 B.n206 10.6151
R1388 B.n210 B.n209 10.6151
R1389 B.n213 B.n210 10.6151
R1390 B.n214 B.n213 10.6151
R1391 B.n217 B.n214 10.6151
R1392 B.n222 B.n219 10.6151
R1393 B.n223 B.n222 10.6151
R1394 B.n226 B.n223 10.6151
R1395 B.n227 B.n226 10.6151
R1396 B.n230 B.n227 10.6151
R1397 B.n231 B.n230 10.6151
R1398 B.n234 B.n231 10.6151
R1399 B.n235 B.n234 10.6151
R1400 B.n238 B.n235 10.6151
R1401 B.n243 B.n240 10.6151
R1402 B.n244 B.n243 10.6151
R1403 B.n247 B.n244 10.6151
R1404 B.n248 B.n247 10.6151
R1405 B.n251 B.n248 10.6151
R1406 B.n252 B.n251 10.6151
R1407 B.n255 B.n252 10.6151
R1408 B.n256 B.n255 10.6151
R1409 B.n259 B.n256 10.6151
R1410 B.n260 B.n259 10.6151
R1411 B.n263 B.n260 10.6151
R1412 B.n264 B.n263 10.6151
R1413 B.n267 B.n264 10.6151
R1414 B.n268 B.n267 10.6151
R1415 B.n271 B.n268 10.6151
R1416 B.n272 B.n271 10.6151
R1417 B.n275 B.n272 10.6151
R1418 B.n276 B.n275 10.6151
R1419 B.n279 B.n276 10.6151
R1420 B.n280 B.n279 10.6151
R1421 B.n283 B.n280 10.6151
R1422 B.n284 B.n283 10.6151
R1423 B.n287 B.n284 10.6151
R1424 B.n288 B.n287 10.6151
R1425 B.n291 B.n288 10.6151
R1426 B.n292 B.n291 10.6151
R1427 B.n295 B.n292 10.6151
R1428 B.n296 B.n295 10.6151
R1429 B.n299 B.n296 10.6151
R1430 B.n300 B.n299 10.6151
R1431 B.n303 B.n300 10.6151
R1432 B.n304 B.n303 10.6151
R1433 B.n307 B.n304 10.6151
R1434 B.n308 B.n307 10.6151
R1435 B.n311 B.n308 10.6151
R1436 B.n312 B.n311 10.6151
R1437 B.n315 B.n312 10.6151
R1438 B.n316 B.n315 10.6151
R1439 B.n319 B.n316 10.6151
R1440 B.n320 B.n319 10.6151
R1441 B.n323 B.n320 10.6151
R1442 B.n324 B.n323 10.6151
R1443 B.n327 B.n324 10.6151
R1444 B.n328 B.n327 10.6151
R1445 B.n331 B.n328 10.6151
R1446 B.n332 B.n331 10.6151
R1447 B.n335 B.n332 10.6151
R1448 B.n336 B.n335 10.6151
R1449 B.n339 B.n336 10.6151
R1450 B.n341 B.n339 10.6151
R1451 B.n342 B.n341 10.6151
R1452 B.n795 B.n342 10.6151
R1453 B.n580 B.n453 9.52245
R1454 B.n557 B.n456 9.52245
R1455 B.n218 B.n217 9.52245
R1456 B.n240 B.n239 9.52245
R1457 B.n852 B.n0 8.11757
R1458 B.n852 B.n1 8.11757
R1459 B.n732 B.t3 2.60036
R1460 B.t0 B.n830 2.60036
R1461 B.n751 B.t1 1.56041
R1462 B.n840 B.t2 1.56041
R1463 B.n577 B.n453 1.09318
R1464 B.n560 B.n456 1.09318
R1465 B.n219 B.n218 1.09318
R1466 B.n239 B.n238 1.09318
R1467 B.t9 B.n377 0.520472
R1468 B.t5 B.n37 0.520472
R1469 VN.n0 VN.t3 263.668
R1470 VN.n1 VN.t2 263.668
R1471 VN.n0 VN.t1 263.252
R1472 VN.n1 VN.t0 263.252
R1473 VN VN.n1 56.2516
R1474 VN VN.n0 9.65694
R1475 VDD2.n2 VDD2.n0 106.487
R1476 VDD2.n2 VDD2.n1 63.9112
R1477 VDD2.n1 VDD2.t3 1.24735
R1478 VDD2.n1 VDD2.t1 1.24735
R1479 VDD2.n0 VDD2.t0 1.24735
R1480 VDD2.n0 VDD2.t2 1.24735
R1481 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.14765f
C1 VP VTAIL 5.24131f
C2 VDD2 VTAIL 6.6152f
C3 VP VDD1 5.79877f
C4 VDD1 VDD2 0.799535f
C5 VP VN 6.24642f
C6 VN VDD2 5.6123f
C7 VDD1 VTAIL 6.56723f
C8 VP VDD2 0.33462f
C9 VN VTAIL 5.22721f
C10 VDD2 B 3.542446f
C11 VDD1 B 7.80692f
C12 VTAIL B 11.771826f
C13 VN B 9.45593f
C14 VP B 7.247967f
C15 VDD2.t0 B 0.332998f
C16 VDD2.t2 B 0.332998f
C17 VDD2.n0 B 3.7598f
C18 VDD2.t3 B 0.332998f
C19 VDD2.t1 B 0.332998f
C20 VDD2.n1 B 3.0213f
C21 VDD2.n2 B 3.93377f
C22 VN.t3 B 2.47498f
C23 VN.t1 B 2.47341f
C24 VN.n0 B 1.75094f
C25 VN.t2 B 2.47498f
C26 VN.t0 B 2.47341f
C27 VN.n1 B 3.23221f
C28 VTAIL.t2 B 2.17136f
C29 VTAIL.n0 B 0.266567f
C30 VTAIL.t4 B 2.17136f
C31 VTAIL.n1 B 0.306211f
C32 VTAIL.t7 B 2.17136f
C33 VTAIL.n2 B 1.25107f
C34 VTAIL.t3 B 2.17137f
C35 VTAIL.n3 B 1.25106f
C36 VTAIL.t1 B 2.17137f
C37 VTAIL.n4 B 0.306197f
C38 VTAIL.t5 B 2.17137f
C39 VTAIL.n5 B 0.306197f
C40 VTAIL.t6 B 2.17136f
C41 VTAIL.n6 B 1.25107f
C42 VTAIL.t0 B 2.17136f
C43 VTAIL.n7 B 1.20569f
C44 VDD1.t0 B 0.33576f
C45 VDD1.t3 B 0.33576f
C46 VDD1.n0 B 3.0467f
C47 VDD1.t1 B 0.33576f
C48 VDD1.t2 B 0.33576f
C49 VDD1.n1 B 3.81792f
C50 VP.n0 B 0.043166f
C51 VP.t3 B 2.38107f
C52 VP.n1 B 0.065416f
C53 VP.t1 B 2.5092f
C54 VP.t2 B 2.5108f
C55 VP.n2 B 3.26268f
C56 VP.t0 B 2.38107f
C57 VP.n3 B 0.934604f
C58 VP.n4 B 1.9417f
C59 VP.n5 B 0.043166f
C60 VP.n6 B 0.032739f
C61 VP.n7 B 0.026493f
C62 VP.n8 B 0.065416f
C63 VP.n9 B 0.934604f
C64 VP.n10 B 0.033937f
.ends

