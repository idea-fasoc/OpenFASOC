* NGSPICE file created from diff_pair_sample_0361.ext - technology: sky130A

.subckt diff_pair_sample_0361 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=0 ps=0 w=12.33 l=2.78
X1 VTAIL.t6 VP.t0 VDD1.t1 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=2.03445 ps=12.66 w=12.33 l=2.78
X2 VDD2.t3 VN.t0 VTAIL.t0 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=2.03445 pd=12.66 as=4.8087 ps=25.44 w=12.33 l=2.78
X3 B.t8 B.t6 B.t7 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=0 ps=0 w=12.33 l=2.78
X4 VDD2.t2 VN.t1 VTAIL.t1 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=2.03445 pd=12.66 as=4.8087 ps=25.44 w=12.33 l=2.78
X5 VTAIL.t7 VN.t2 VDD2.t1 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=2.03445 ps=12.66 w=12.33 l=2.78
X6 VTAIL.t5 VP.t1 VDD1.t2 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=2.03445 ps=12.66 w=12.33 l=2.78
X7 B.t5 B.t3 B.t4 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=0 ps=0 w=12.33 l=2.78
X8 B.t2 B.t0 B.t1 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=0 ps=0 w=12.33 l=2.78
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=4.8087 pd=25.44 as=2.03445 ps=12.66 w=12.33 l=2.78
X10 VDD1.t3 VP.t2 VTAIL.t4 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=2.03445 pd=12.66 as=4.8087 ps=25.44 w=12.33 l=2.78
X11 VDD1.t0 VP.t3 VTAIL.t3 w_n2836_n3434# sky130_fd_pr__pfet_01v8 ad=2.03445 pd=12.66 as=4.8087 ps=25.44 w=12.33 l=2.78
R0 B.n370 B.n107 585
R1 B.n369 B.n368 585
R2 B.n367 B.n108 585
R3 B.n366 B.n365 585
R4 B.n364 B.n109 585
R5 B.n363 B.n362 585
R6 B.n361 B.n110 585
R7 B.n360 B.n359 585
R8 B.n358 B.n111 585
R9 B.n357 B.n356 585
R10 B.n355 B.n112 585
R11 B.n354 B.n353 585
R12 B.n352 B.n113 585
R13 B.n351 B.n350 585
R14 B.n349 B.n114 585
R15 B.n348 B.n347 585
R16 B.n346 B.n115 585
R17 B.n345 B.n344 585
R18 B.n343 B.n116 585
R19 B.n342 B.n341 585
R20 B.n340 B.n117 585
R21 B.n339 B.n338 585
R22 B.n337 B.n118 585
R23 B.n336 B.n335 585
R24 B.n334 B.n119 585
R25 B.n333 B.n332 585
R26 B.n331 B.n120 585
R27 B.n330 B.n329 585
R28 B.n328 B.n121 585
R29 B.n327 B.n326 585
R30 B.n325 B.n122 585
R31 B.n324 B.n323 585
R32 B.n322 B.n123 585
R33 B.n321 B.n320 585
R34 B.n319 B.n124 585
R35 B.n318 B.n317 585
R36 B.n316 B.n125 585
R37 B.n315 B.n314 585
R38 B.n313 B.n126 585
R39 B.n312 B.n311 585
R40 B.n310 B.n127 585
R41 B.n309 B.n308 585
R42 B.n307 B.n128 585
R43 B.n306 B.n305 585
R44 B.n301 B.n129 585
R45 B.n300 B.n299 585
R46 B.n298 B.n130 585
R47 B.n297 B.n296 585
R48 B.n295 B.n131 585
R49 B.n294 B.n293 585
R50 B.n292 B.n132 585
R51 B.n291 B.n290 585
R52 B.n288 B.n133 585
R53 B.n287 B.n286 585
R54 B.n285 B.n136 585
R55 B.n284 B.n283 585
R56 B.n282 B.n137 585
R57 B.n281 B.n280 585
R58 B.n279 B.n138 585
R59 B.n278 B.n277 585
R60 B.n276 B.n139 585
R61 B.n275 B.n274 585
R62 B.n273 B.n140 585
R63 B.n272 B.n271 585
R64 B.n270 B.n141 585
R65 B.n269 B.n268 585
R66 B.n267 B.n142 585
R67 B.n266 B.n265 585
R68 B.n264 B.n143 585
R69 B.n263 B.n262 585
R70 B.n261 B.n144 585
R71 B.n260 B.n259 585
R72 B.n258 B.n145 585
R73 B.n257 B.n256 585
R74 B.n255 B.n146 585
R75 B.n254 B.n253 585
R76 B.n252 B.n147 585
R77 B.n251 B.n250 585
R78 B.n249 B.n148 585
R79 B.n248 B.n247 585
R80 B.n246 B.n149 585
R81 B.n245 B.n244 585
R82 B.n243 B.n150 585
R83 B.n242 B.n241 585
R84 B.n240 B.n151 585
R85 B.n239 B.n238 585
R86 B.n237 B.n152 585
R87 B.n236 B.n235 585
R88 B.n234 B.n153 585
R89 B.n233 B.n232 585
R90 B.n231 B.n154 585
R91 B.n230 B.n229 585
R92 B.n228 B.n155 585
R93 B.n227 B.n226 585
R94 B.n225 B.n156 585
R95 B.n372 B.n371 585
R96 B.n373 B.n106 585
R97 B.n375 B.n374 585
R98 B.n376 B.n105 585
R99 B.n378 B.n377 585
R100 B.n379 B.n104 585
R101 B.n381 B.n380 585
R102 B.n382 B.n103 585
R103 B.n384 B.n383 585
R104 B.n385 B.n102 585
R105 B.n387 B.n386 585
R106 B.n388 B.n101 585
R107 B.n390 B.n389 585
R108 B.n391 B.n100 585
R109 B.n393 B.n392 585
R110 B.n394 B.n99 585
R111 B.n396 B.n395 585
R112 B.n397 B.n98 585
R113 B.n399 B.n398 585
R114 B.n400 B.n97 585
R115 B.n402 B.n401 585
R116 B.n403 B.n96 585
R117 B.n405 B.n404 585
R118 B.n406 B.n95 585
R119 B.n408 B.n407 585
R120 B.n409 B.n94 585
R121 B.n411 B.n410 585
R122 B.n412 B.n93 585
R123 B.n414 B.n413 585
R124 B.n415 B.n92 585
R125 B.n417 B.n416 585
R126 B.n418 B.n91 585
R127 B.n420 B.n419 585
R128 B.n421 B.n90 585
R129 B.n423 B.n422 585
R130 B.n424 B.n89 585
R131 B.n426 B.n425 585
R132 B.n427 B.n88 585
R133 B.n429 B.n428 585
R134 B.n430 B.n87 585
R135 B.n432 B.n431 585
R136 B.n433 B.n86 585
R137 B.n435 B.n434 585
R138 B.n436 B.n85 585
R139 B.n438 B.n437 585
R140 B.n439 B.n84 585
R141 B.n441 B.n440 585
R142 B.n442 B.n83 585
R143 B.n444 B.n443 585
R144 B.n445 B.n82 585
R145 B.n447 B.n446 585
R146 B.n448 B.n81 585
R147 B.n450 B.n449 585
R148 B.n451 B.n80 585
R149 B.n453 B.n452 585
R150 B.n454 B.n79 585
R151 B.n456 B.n455 585
R152 B.n457 B.n78 585
R153 B.n459 B.n458 585
R154 B.n460 B.n77 585
R155 B.n462 B.n461 585
R156 B.n463 B.n76 585
R157 B.n465 B.n464 585
R158 B.n466 B.n75 585
R159 B.n468 B.n467 585
R160 B.n469 B.n74 585
R161 B.n471 B.n470 585
R162 B.n472 B.n73 585
R163 B.n474 B.n473 585
R164 B.n475 B.n72 585
R165 B.n477 B.n476 585
R166 B.n478 B.n71 585
R167 B.n623 B.n622 585
R168 B.n621 B.n20 585
R169 B.n620 B.n619 585
R170 B.n618 B.n21 585
R171 B.n617 B.n616 585
R172 B.n615 B.n22 585
R173 B.n614 B.n613 585
R174 B.n612 B.n23 585
R175 B.n611 B.n610 585
R176 B.n609 B.n24 585
R177 B.n608 B.n607 585
R178 B.n606 B.n25 585
R179 B.n605 B.n604 585
R180 B.n603 B.n26 585
R181 B.n602 B.n601 585
R182 B.n600 B.n27 585
R183 B.n599 B.n598 585
R184 B.n597 B.n28 585
R185 B.n596 B.n595 585
R186 B.n594 B.n29 585
R187 B.n593 B.n592 585
R188 B.n591 B.n30 585
R189 B.n590 B.n589 585
R190 B.n588 B.n31 585
R191 B.n587 B.n586 585
R192 B.n585 B.n32 585
R193 B.n584 B.n583 585
R194 B.n582 B.n33 585
R195 B.n581 B.n580 585
R196 B.n579 B.n34 585
R197 B.n578 B.n577 585
R198 B.n576 B.n35 585
R199 B.n575 B.n574 585
R200 B.n573 B.n36 585
R201 B.n572 B.n571 585
R202 B.n570 B.n37 585
R203 B.n569 B.n568 585
R204 B.n567 B.n38 585
R205 B.n566 B.n565 585
R206 B.n564 B.n39 585
R207 B.n563 B.n562 585
R208 B.n561 B.n40 585
R209 B.n560 B.n559 585
R210 B.n557 B.n41 585
R211 B.n556 B.n555 585
R212 B.n554 B.n44 585
R213 B.n553 B.n552 585
R214 B.n551 B.n45 585
R215 B.n550 B.n549 585
R216 B.n548 B.n46 585
R217 B.n547 B.n546 585
R218 B.n545 B.n47 585
R219 B.n543 B.n542 585
R220 B.n541 B.n50 585
R221 B.n540 B.n539 585
R222 B.n538 B.n51 585
R223 B.n537 B.n536 585
R224 B.n535 B.n52 585
R225 B.n534 B.n533 585
R226 B.n532 B.n53 585
R227 B.n531 B.n530 585
R228 B.n529 B.n54 585
R229 B.n528 B.n527 585
R230 B.n526 B.n55 585
R231 B.n525 B.n524 585
R232 B.n523 B.n56 585
R233 B.n522 B.n521 585
R234 B.n520 B.n57 585
R235 B.n519 B.n518 585
R236 B.n517 B.n58 585
R237 B.n516 B.n515 585
R238 B.n514 B.n59 585
R239 B.n513 B.n512 585
R240 B.n511 B.n60 585
R241 B.n510 B.n509 585
R242 B.n508 B.n61 585
R243 B.n507 B.n506 585
R244 B.n505 B.n62 585
R245 B.n504 B.n503 585
R246 B.n502 B.n63 585
R247 B.n501 B.n500 585
R248 B.n499 B.n64 585
R249 B.n498 B.n497 585
R250 B.n496 B.n65 585
R251 B.n495 B.n494 585
R252 B.n493 B.n66 585
R253 B.n492 B.n491 585
R254 B.n490 B.n67 585
R255 B.n489 B.n488 585
R256 B.n487 B.n68 585
R257 B.n486 B.n485 585
R258 B.n484 B.n69 585
R259 B.n483 B.n482 585
R260 B.n481 B.n70 585
R261 B.n480 B.n479 585
R262 B.n624 B.n19 585
R263 B.n626 B.n625 585
R264 B.n627 B.n18 585
R265 B.n629 B.n628 585
R266 B.n630 B.n17 585
R267 B.n632 B.n631 585
R268 B.n633 B.n16 585
R269 B.n635 B.n634 585
R270 B.n636 B.n15 585
R271 B.n638 B.n637 585
R272 B.n639 B.n14 585
R273 B.n641 B.n640 585
R274 B.n642 B.n13 585
R275 B.n644 B.n643 585
R276 B.n645 B.n12 585
R277 B.n647 B.n646 585
R278 B.n648 B.n11 585
R279 B.n650 B.n649 585
R280 B.n651 B.n10 585
R281 B.n653 B.n652 585
R282 B.n654 B.n9 585
R283 B.n656 B.n655 585
R284 B.n657 B.n8 585
R285 B.n659 B.n658 585
R286 B.n660 B.n7 585
R287 B.n662 B.n661 585
R288 B.n663 B.n6 585
R289 B.n665 B.n664 585
R290 B.n666 B.n5 585
R291 B.n668 B.n667 585
R292 B.n669 B.n4 585
R293 B.n671 B.n670 585
R294 B.n672 B.n3 585
R295 B.n674 B.n673 585
R296 B.n675 B.n0 585
R297 B.n2 B.n1 585
R298 B.n174 B.n173 585
R299 B.n176 B.n175 585
R300 B.n177 B.n172 585
R301 B.n179 B.n178 585
R302 B.n180 B.n171 585
R303 B.n182 B.n181 585
R304 B.n183 B.n170 585
R305 B.n185 B.n184 585
R306 B.n186 B.n169 585
R307 B.n188 B.n187 585
R308 B.n189 B.n168 585
R309 B.n191 B.n190 585
R310 B.n192 B.n167 585
R311 B.n194 B.n193 585
R312 B.n195 B.n166 585
R313 B.n197 B.n196 585
R314 B.n198 B.n165 585
R315 B.n200 B.n199 585
R316 B.n201 B.n164 585
R317 B.n203 B.n202 585
R318 B.n204 B.n163 585
R319 B.n206 B.n205 585
R320 B.n207 B.n162 585
R321 B.n209 B.n208 585
R322 B.n210 B.n161 585
R323 B.n212 B.n211 585
R324 B.n213 B.n160 585
R325 B.n215 B.n214 585
R326 B.n216 B.n159 585
R327 B.n218 B.n217 585
R328 B.n219 B.n158 585
R329 B.n221 B.n220 585
R330 B.n222 B.n157 585
R331 B.n224 B.n223 585
R332 B.n225 B.n224 487.695
R333 B.n372 B.n107 487.695
R334 B.n480 B.n71 487.695
R335 B.n622 B.n19 487.695
R336 B.n134 B.t9 315.193
R337 B.n302 B.t3 315.193
R338 B.n48 B.t0 315.193
R339 B.n42 B.t6 315.193
R340 B.n677 B.n676 256.663
R341 B.n676 B.n675 235.042
R342 B.n676 B.n2 235.042
R343 B.n302 B.t4 169.091
R344 B.n48 B.t2 169.091
R345 B.n134 B.t10 169.077
R346 B.n42 B.t8 169.077
R347 B.n226 B.n225 163.367
R348 B.n226 B.n155 163.367
R349 B.n230 B.n155 163.367
R350 B.n231 B.n230 163.367
R351 B.n232 B.n231 163.367
R352 B.n232 B.n153 163.367
R353 B.n236 B.n153 163.367
R354 B.n237 B.n236 163.367
R355 B.n238 B.n237 163.367
R356 B.n238 B.n151 163.367
R357 B.n242 B.n151 163.367
R358 B.n243 B.n242 163.367
R359 B.n244 B.n243 163.367
R360 B.n244 B.n149 163.367
R361 B.n248 B.n149 163.367
R362 B.n249 B.n248 163.367
R363 B.n250 B.n249 163.367
R364 B.n250 B.n147 163.367
R365 B.n254 B.n147 163.367
R366 B.n255 B.n254 163.367
R367 B.n256 B.n255 163.367
R368 B.n256 B.n145 163.367
R369 B.n260 B.n145 163.367
R370 B.n261 B.n260 163.367
R371 B.n262 B.n261 163.367
R372 B.n262 B.n143 163.367
R373 B.n266 B.n143 163.367
R374 B.n267 B.n266 163.367
R375 B.n268 B.n267 163.367
R376 B.n268 B.n141 163.367
R377 B.n272 B.n141 163.367
R378 B.n273 B.n272 163.367
R379 B.n274 B.n273 163.367
R380 B.n274 B.n139 163.367
R381 B.n278 B.n139 163.367
R382 B.n279 B.n278 163.367
R383 B.n280 B.n279 163.367
R384 B.n280 B.n137 163.367
R385 B.n284 B.n137 163.367
R386 B.n285 B.n284 163.367
R387 B.n286 B.n285 163.367
R388 B.n286 B.n133 163.367
R389 B.n291 B.n133 163.367
R390 B.n292 B.n291 163.367
R391 B.n293 B.n292 163.367
R392 B.n293 B.n131 163.367
R393 B.n297 B.n131 163.367
R394 B.n298 B.n297 163.367
R395 B.n299 B.n298 163.367
R396 B.n299 B.n129 163.367
R397 B.n306 B.n129 163.367
R398 B.n307 B.n306 163.367
R399 B.n308 B.n307 163.367
R400 B.n308 B.n127 163.367
R401 B.n312 B.n127 163.367
R402 B.n313 B.n312 163.367
R403 B.n314 B.n313 163.367
R404 B.n314 B.n125 163.367
R405 B.n318 B.n125 163.367
R406 B.n319 B.n318 163.367
R407 B.n320 B.n319 163.367
R408 B.n320 B.n123 163.367
R409 B.n324 B.n123 163.367
R410 B.n325 B.n324 163.367
R411 B.n326 B.n325 163.367
R412 B.n326 B.n121 163.367
R413 B.n330 B.n121 163.367
R414 B.n331 B.n330 163.367
R415 B.n332 B.n331 163.367
R416 B.n332 B.n119 163.367
R417 B.n336 B.n119 163.367
R418 B.n337 B.n336 163.367
R419 B.n338 B.n337 163.367
R420 B.n338 B.n117 163.367
R421 B.n342 B.n117 163.367
R422 B.n343 B.n342 163.367
R423 B.n344 B.n343 163.367
R424 B.n344 B.n115 163.367
R425 B.n348 B.n115 163.367
R426 B.n349 B.n348 163.367
R427 B.n350 B.n349 163.367
R428 B.n350 B.n113 163.367
R429 B.n354 B.n113 163.367
R430 B.n355 B.n354 163.367
R431 B.n356 B.n355 163.367
R432 B.n356 B.n111 163.367
R433 B.n360 B.n111 163.367
R434 B.n361 B.n360 163.367
R435 B.n362 B.n361 163.367
R436 B.n362 B.n109 163.367
R437 B.n366 B.n109 163.367
R438 B.n367 B.n366 163.367
R439 B.n368 B.n367 163.367
R440 B.n368 B.n107 163.367
R441 B.n476 B.n71 163.367
R442 B.n476 B.n475 163.367
R443 B.n475 B.n474 163.367
R444 B.n474 B.n73 163.367
R445 B.n470 B.n73 163.367
R446 B.n470 B.n469 163.367
R447 B.n469 B.n468 163.367
R448 B.n468 B.n75 163.367
R449 B.n464 B.n75 163.367
R450 B.n464 B.n463 163.367
R451 B.n463 B.n462 163.367
R452 B.n462 B.n77 163.367
R453 B.n458 B.n77 163.367
R454 B.n458 B.n457 163.367
R455 B.n457 B.n456 163.367
R456 B.n456 B.n79 163.367
R457 B.n452 B.n79 163.367
R458 B.n452 B.n451 163.367
R459 B.n451 B.n450 163.367
R460 B.n450 B.n81 163.367
R461 B.n446 B.n81 163.367
R462 B.n446 B.n445 163.367
R463 B.n445 B.n444 163.367
R464 B.n444 B.n83 163.367
R465 B.n440 B.n83 163.367
R466 B.n440 B.n439 163.367
R467 B.n439 B.n438 163.367
R468 B.n438 B.n85 163.367
R469 B.n434 B.n85 163.367
R470 B.n434 B.n433 163.367
R471 B.n433 B.n432 163.367
R472 B.n432 B.n87 163.367
R473 B.n428 B.n87 163.367
R474 B.n428 B.n427 163.367
R475 B.n427 B.n426 163.367
R476 B.n426 B.n89 163.367
R477 B.n422 B.n89 163.367
R478 B.n422 B.n421 163.367
R479 B.n421 B.n420 163.367
R480 B.n420 B.n91 163.367
R481 B.n416 B.n91 163.367
R482 B.n416 B.n415 163.367
R483 B.n415 B.n414 163.367
R484 B.n414 B.n93 163.367
R485 B.n410 B.n93 163.367
R486 B.n410 B.n409 163.367
R487 B.n409 B.n408 163.367
R488 B.n408 B.n95 163.367
R489 B.n404 B.n95 163.367
R490 B.n404 B.n403 163.367
R491 B.n403 B.n402 163.367
R492 B.n402 B.n97 163.367
R493 B.n398 B.n97 163.367
R494 B.n398 B.n397 163.367
R495 B.n397 B.n396 163.367
R496 B.n396 B.n99 163.367
R497 B.n392 B.n99 163.367
R498 B.n392 B.n391 163.367
R499 B.n391 B.n390 163.367
R500 B.n390 B.n101 163.367
R501 B.n386 B.n101 163.367
R502 B.n386 B.n385 163.367
R503 B.n385 B.n384 163.367
R504 B.n384 B.n103 163.367
R505 B.n380 B.n103 163.367
R506 B.n380 B.n379 163.367
R507 B.n379 B.n378 163.367
R508 B.n378 B.n105 163.367
R509 B.n374 B.n105 163.367
R510 B.n374 B.n373 163.367
R511 B.n373 B.n372 163.367
R512 B.n622 B.n621 163.367
R513 B.n621 B.n620 163.367
R514 B.n620 B.n21 163.367
R515 B.n616 B.n21 163.367
R516 B.n616 B.n615 163.367
R517 B.n615 B.n614 163.367
R518 B.n614 B.n23 163.367
R519 B.n610 B.n23 163.367
R520 B.n610 B.n609 163.367
R521 B.n609 B.n608 163.367
R522 B.n608 B.n25 163.367
R523 B.n604 B.n25 163.367
R524 B.n604 B.n603 163.367
R525 B.n603 B.n602 163.367
R526 B.n602 B.n27 163.367
R527 B.n598 B.n27 163.367
R528 B.n598 B.n597 163.367
R529 B.n597 B.n596 163.367
R530 B.n596 B.n29 163.367
R531 B.n592 B.n29 163.367
R532 B.n592 B.n591 163.367
R533 B.n591 B.n590 163.367
R534 B.n590 B.n31 163.367
R535 B.n586 B.n31 163.367
R536 B.n586 B.n585 163.367
R537 B.n585 B.n584 163.367
R538 B.n584 B.n33 163.367
R539 B.n580 B.n33 163.367
R540 B.n580 B.n579 163.367
R541 B.n579 B.n578 163.367
R542 B.n578 B.n35 163.367
R543 B.n574 B.n35 163.367
R544 B.n574 B.n573 163.367
R545 B.n573 B.n572 163.367
R546 B.n572 B.n37 163.367
R547 B.n568 B.n37 163.367
R548 B.n568 B.n567 163.367
R549 B.n567 B.n566 163.367
R550 B.n566 B.n39 163.367
R551 B.n562 B.n39 163.367
R552 B.n562 B.n561 163.367
R553 B.n561 B.n560 163.367
R554 B.n560 B.n41 163.367
R555 B.n555 B.n41 163.367
R556 B.n555 B.n554 163.367
R557 B.n554 B.n553 163.367
R558 B.n553 B.n45 163.367
R559 B.n549 B.n45 163.367
R560 B.n549 B.n548 163.367
R561 B.n548 B.n547 163.367
R562 B.n547 B.n47 163.367
R563 B.n542 B.n47 163.367
R564 B.n542 B.n541 163.367
R565 B.n541 B.n540 163.367
R566 B.n540 B.n51 163.367
R567 B.n536 B.n51 163.367
R568 B.n536 B.n535 163.367
R569 B.n535 B.n534 163.367
R570 B.n534 B.n53 163.367
R571 B.n530 B.n53 163.367
R572 B.n530 B.n529 163.367
R573 B.n529 B.n528 163.367
R574 B.n528 B.n55 163.367
R575 B.n524 B.n55 163.367
R576 B.n524 B.n523 163.367
R577 B.n523 B.n522 163.367
R578 B.n522 B.n57 163.367
R579 B.n518 B.n57 163.367
R580 B.n518 B.n517 163.367
R581 B.n517 B.n516 163.367
R582 B.n516 B.n59 163.367
R583 B.n512 B.n59 163.367
R584 B.n512 B.n511 163.367
R585 B.n511 B.n510 163.367
R586 B.n510 B.n61 163.367
R587 B.n506 B.n61 163.367
R588 B.n506 B.n505 163.367
R589 B.n505 B.n504 163.367
R590 B.n504 B.n63 163.367
R591 B.n500 B.n63 163.367
R592 B.n500 B.n499 163.367
R593 B.n499 B.n498 163.367
R594 B.n498 B.n65 163.367
R595 B.n494 B.n65 163.367
R596 B.n494 B.n493 163.367
R597 B.n493 B.n492 163.367
R598 B.n492 B.n67 163.367
R599 B.n488 B.n67 163.367
R600 B.n488 B.n487 163.367
R601 B.n487 B.n486 163.367
R602 B.n486 B.n69 163.367
R603 B.n482 B.n69 163.367
R604 B.n482 B.n481 163.367
R605 B.n481 B.n480 163.367
R606 B.n626 B.n19 163.367
R607 B.n627 B.n626 163.367
R608 B.n628 B.n627 163.367
R609 B.n628 B.n17 163.367
R610 B.n632 B.n17 163.367
R611 B.n633 B.n632 163.367
R612 B.n634 B.n633 163.367
R613 B.n634 B.n15 163.367
R614 B.n638 B.n15 163.367
R615 B.n639 B.n638 163.367
R616 B.n640 B.n639 163.367
R617 B.n640 B.n13 163.367
R618 B.n644 B.n13 163.367
R619 B.n645 B.n644 163.367
R620 B.n646 B.n645 163.367
R621 B.n646 B.n11 163.367
R622 B.n650 B.n11 163.367
R623 B.n651 B.n650 163.367
R624 B.n652 B.n651 163.367
R625 B.n652 B.n9 163.367
R626 B.n656 B.n9 163.367
R627 B.n657 B.n656 163.367
R628 B.n658 B.n657 163.367
R629 B.n658 B.n7 163.367
R630 B.n662 B.n7 163.367
R631 B.n663 B.n662 163.367
R632 B.n664 B.n663 163.367
R633 B.n664 B.n5 163.367
R634 B.n668 B.n5 163.367
R635 B.n669 B.n668 163.367
R636 B.n670 B.n669 163.367
R637 B.n670 B.n3 163.367
R638 B.n674 B.n3 163.367
R639 B.n675 B.n674 163.367
R640 B.n173 B.n2 163.367
R641 B.n176 B.n173 163.367
R642 B.n177 B.n176 163.367
R643 B.n178 B.n177 163.367
R644 B.n178 B.n171 163.367
R645 B.n182 B.n171 163.367
R646 B.n183 B.n182 163.367
R647 B.n184 B.n183 163.367
R648 B.n184 B.n169 163.367
R649 B.n188 B.n169 163.367
R650 B.n189 B.n188 163.367
R651 B.n190 B.n189 163.367
R652 B.n190 B.n167 163.367
R653 B.n194 B.n167 163.367
R654 B.n195 B.n194 163.367
R655 B.n196 B.n195 163.367
R656 B.n196 B.n165 163.367
R657 B.n200 B.n165 163.367
R658 B.n201 B.n200 163.367
R659 B.n202 B.n201 163.367
R660 B.n202 B.n163 163.367
R661 B.n206 B.n163 163.367
R662 B.n207 B.n206 163.367
R663 B.n208 B.n207 163.367
R664 B.n208 B.n161 163.367
R665 B.n212 B.n161 163.367
R666 B.n213 B.n212 163.367
R667 B.n214 B.n213 163.367
R668 B.n214 B.n159 163.367
R669 B.n218 B.n159 163.367
R670 B.n219 B.n218 163.367
R671 B.n220 B.n219 163.367
R672 B.n220 B.n157 163.367
R673 B.n224 B.n157 163.367
R674 B.n303 B.t5 108.776
R675 B.n49 B.t1 108.776
R676 B.n135 B.t11 108.761
R677 B.n43 B.t7 108.761
R678 B.n135 B.n134 60.3157
R679 B.n303 B.n302 60.3157
R680 B.n49 B.n48 60.3157
R681 B.n43 B.n42 60.3157
R682 B.n289 B.n135 59.5399
R683 B.n304 B.n303 59.5399
R684 B.n544 B.n49 59.5399
R685 B.n558 B.n43 59.5399
R686 B.n624 B.n623 31.6883
R687 B.n479 B.n478 31.6883
R688 B.n371 B.n370 31.6883
R689 B.n223 B.n156 31.6883
R690 B B.n677 18.0485
R691 B.n625 B.n624 10.6151
R692 B.n625 B.n18 10.6151
R693 B.n629 B.n18 10.6151
R694 B.n630 B.n629 10.6151
R695 B.n631 B.n630 10.6151
R696 B.n631 B.n16 10.6151
R697 B.n635 B.n16 10.6151
R698 B.n636 B.n635 10.6151
R699 B.n637 B.n636 10.6151
R700 B.n637 B.n14 10.6151
R701 B.n641 B.n14 10.6151
R702 B.n642 B.n641 10.6151
R703 B.n643 B.n642 10.6151
R704 B.n643 B.n12 10.6151
R705 B.n647 B.n12 10.6151
R706 B.n648 B.n647 10.6151
R707 B.n649 B.n648 10.6151
R708 B.n649 B.n10 10.6151
R709 B.n653 B.n10 10.6151
R710 B.n654 B.n653 10.6151
R711 B.n655 B.n654 10.6151
R712 B.n655 B.n8 10.6151
R713 B.n659 B.n8 10.6151
R714 B.n660 B.n659 10.6151
R715 B.n661 B.n660 10.6151
R716 B.n661 B.n6 10.6151
R717 B.n665 B.n6 10.6151
R718 B.n666 B.n665 10.6151
R719 B.n667 B.n666 10.6151
R720 B.n667 B.n4 10.6151
R721 B.n671 B.n4 10.6151
R722 B.n672 B.n671 10.6151
R723 B.n673 B.n672 10.6151
R724 B.n673 B.n0 10.6151
R725 B.n623 B.n20 10.6151
R726 B.n619 B.n20 10.6151
R727 B.n619 B.n618 10.6151
R728 B.n618 B.n617 10.6151
R729 B.n617 B.n22 10.6151
R730 B.n613 B.n22 10.6151
R731 B.n613 B.n612 10.6151
R732 B.n612 B.n611 10.6151
R733 B.n611 B.n24 10.6151
R734 B.n607 B.n24 10.6151
R735 B.n607 B.n606 10.6151
R736 B.n606 B.n605 10.6151
R737 B.n605 B.n26 10.6151
R738 B.n601 B.n26 10.6151
R739 B.n601 B.n600 10.6151
R740 B.n600 B.n599 10.6151
R741 B.n599 B.n28 10.6151
R742 B.n595 B.n28 10.6151
R743 B.n595 B.n594 10.6151
R744 B.n594 B.n593 10.6151
R745 B.n593 B.n30 10.6151
R746 B.n589 B.n30 10.6151
R747 B.n589 B.n588 10.6151
R748 B.n588 B.n587 10.6151
R749 B.n587 B.n32 10.6151
R750 B.n583 B.n32 10.6151
R751 B.n583 B.n582 10.6151
R752 B.n582 B.n581 10.6151
R753 B.n581 B.n34 10.6151
R754 B.n577 B.n34 10.6151
R755 B.n577 B.n576 10.6151
R756 B.n576 B.n575 10.6151
R757 B.n575 B.n36 10.6151
R758 B.n571 B.n36 10.6151
R759 B.n571 B.n570 10.6151
R760 B.n570 B.n569 10.6151
R761 B.n569 B.n38 10.6151
R762 B.n565 B.n38 10.6151
R763 B.n565 B.n564 10.6151
R764 B.n564 B.n563 10.6151
R765 B.n563 B.n40 10.6151
R766 B.n559 B.n40 10.6151
R767 B.n557 B.n556 10.6151
R768 B.n556 B.n44 10.6151
R769 B.n552 B.n44 10.6151
R770 B.n552 B.n551 10.6151
R771 B.n551 B.n550 10.6151
R772 B.n550 B.n46 10.6151
R773 B.n546 B.n46 10.6151
R774 B.n546 B.n545 10.6151
R775 B.n543 B.n50 10.6151
R776 B.n539 B.n50 10.6151
R777 B.n539 B.n538 10.6151
R778 B.n538 B.n537 10.6151
R779 B.n537 B.n52 10.6151
R780 B.n533 B.n52 10.6151
R781 B.n533 B.n532 10.6151
R782 B.n532 B.n531 10.6151
R783 B.n531 B.n54 10.6151
R784 B.n527 B.n54 10.6151
R785 B.n527 B.n526 10.6151
R786 B.n526 B.n525 10.6151
R787 B.n525 B.n56 10.6151
R788 B.n521 B.n56 10.6151
R789 B.n521 B.n520 10.6151
R790 B.n520 B.n519 10.6151
R791 B.n519 B.n58 10.6151
R792 B.n515 B.n58 10.6151
R793 B.n515 B.n514 10.6151
R794 B.n514 B.n513 10.6151
R795 B.n513 B.n60 10.6151
R796 B.n509 B.n60 10.6151
R797 B.n509 B.n508 10.6151
R798 B.n508 B.n507 10.6151
R799 B.n507 B.n62 10.6151
R800 B.n503 B.n62 10.6151
R801 B.n503 B.n502 10.6151
R802 B.n502 B.n501 10.6151
R803 B.n501 B.n64 10.6151
R804 B.n497 B.n64 10.6151
R805 B.n497 B.n496 10.6151
R806 B.n496 B.n495 10.6151
R807 B.n495 B.n66 10.6151
R808 B.n491 B.n66 10.6151
R809 B.n491 B.n490 10.6151
R810 B.n490 B.n489 10.6151
R811 B.n489 B.n68 10.6151
R812 B.n485 B.n68 10.6151
R813 B.n485 B.n484 10.6151
R814 B.n484 B.n483 10.6151
R815 B.n483 B.n70 10.6151
R816 B.n479 B.n70 10.6151
R817 B.n478 B.n477 10.6151
R818 B.n477 B.n72 10.6151
R819 B.n473 B.n72 10.6151
R820 B.n473 B.n472 10.6151
R821 B.n472 B.n471 10.6151
R822 B.n471 B.n74 10.6151
R823 B.n467 B.n74 10.6151
R824 B.n467 B.n466 10.6151
R825 B.n466 B.n465 10.6151
R826 B.n465 B.n76 10.6151
R827 B.n461 B.n76 10.6151
R828 B.n461 B.n460 10.6151
R829 B.n460 B.n459 10.6151
R830 B.n459 B.n78 10.6151
R831 B.n455 B.n78 10.6151
R832 B.n455 B.n454 10.6151
R833 B.n454 B.n453 10.6151
R834 B.n453 B.n80 10.6151
R835 B.n449 B.n80 10.6151
R836 B.n449 B.n448 10.6151
R837 B.n448 B.n447 10.6151
R838 B.n447 B.n82 10.6151
R839 B.n443 B.n82 10.6151
R840 B.n443 B.n442 10.6151
R841 B.n442 B.n441 10.6151
R842 B.n441 B.n84 10.6151
R843 B.n437 B.n84 10.6151
R844 B.n437 B.n436 10.6151
R845 B.n436 B.n435 10.6151
R846 B.n435 B.n86 10.6151
R847 B.n431 B.n86 10.6151
R848 B.n431 B.n430 10.6151
R849 B.n430 B.n429 10.6151
R850 B.n429 B.n88 10.6151
R851 B.n425 B.n88 10.6151
R852 B.n425 B.n424 10.6151
R853 B.n424 B.n423 10.6151
R854 B.n423 B.n90 10.6151
R855 B.n419 B.n90 10.6151
R856 B.n419 B.n418 10.6151
R857 B.n418 B.n417 10.6151
R858 B.n417 B.n92 10.6151
R859 B.n413 B.n92 10.6151
R860 B.n413 B.n412 10.6151
R861 B.n412 B.n411 10.6151
R862 B.n411 B.n94 10.6151
R863 B.n407 B.n94 10.6151
R864 B.n407 B.n406 10.6151
R865 B.n406 B.n405 10.6151
R866 B.n405 B.n96 10.6151
R867 B.n401 B.n96 10.6151
R868 B.n401 B.n400 10.6151
R869 B.n400 B.n399 10.6151
R870 B.n399 B.n98 10.6151
R871 B.n395 B.n98 10.6151
R872 B.n395 B.n394 10.6151
R873 B.n394 B.n393 10.6151
R874 B.n393 B.n100 10.6151
R875 B.n389 B.n100 10.6151
R876 B.n389 B.n388 10.6151
R877 B.n388 B.n387 10.6151
R878 B.n387 B.n102 10.6151
R879 B.n383 B.n102 10.6151
R880 B.n383 B.n382 10.6151
R881 B.n382 B.n381 10.6151
R882 B.n381 B.n104 10.6151
R883 B.n377 B.n104 10.6151
R884 B.n377 B.n376 10.6151
R885 B.n376 B.n375 10.6151
R886 B.n375 B.n106 10.6151
R887 B.n371 B.n106 10.6151
R888 B.n174 B.n1 10.6151
R889 B.n175 B.n174 10.6151
R890 B.n175 B.n172 10.6151
R891 B.n179 B.n172 10.6151
R892 B.n180 B.n179 10.6151
R893 B.n181 B.n180 10.6151
R894 B.n181 B.n170 10.6151
R895 B.n185 B.n170 10.6151
R896 B.n186 B.n185 10.6151
R897 B.n187 B.n186 10.6151
R898 B.n187 B.n168 10.6151
R899 B.n191 B.n168 10.6151
R900 B.n192 B.n191 10.6151
R901 B.n193 B.n192 10.6151
R902 B.n193 B.n166 10.6151
R903 B.n197 B.n166 10.6151
R904 B.n198 B.n197 10.6151
R905 B.n199 B.n198 10.6151
R906 B.n199 B.n164 10.6151
R907 B.n203 B.n164 10.6151
R908 B.n204 B.n203 10.6151
R909 B.n205 B.n204 10.6151
R910 B.n205 B.n162 10.6151
R911 B.n209 B.n162 10.6151
R912 B.n210 B.n209 10.6151
R913 B.n211 B.n210 10.6151
R914 B.n211 B.n160 10.6151
R915 B.n215 B.n160 10.6151
R916 B.n216 B.n215 10.6151
R917 B.n217 B.n216 10.6151
R918 B.n217 B.n158 10.6151
R919 B.n221 B.n158 10.6151
R920 B.n222 B.n221 10.6151
R921 B.n223 B.n222 10.6151
R922 B.n227 B.n156 10.6151
R923 B.n228 B.n227 10.6151
R924 B.n229 B.n228 10.6151
R925 B.n229 B.n154 10.6151
R926 B.n233 B.n154 10.6151
R927 B.n234 B.n233 10.6151
R928 B.n235 B.n234 10.6151
R929 B.n235 B.n152 10.6151
R930 B.n239 B.n152 10.6151
R931 B.n240 B.n239 10.6151
R932 B.n241 B.n240 10.6151
R933 B.n241 B.n150 10.6151
R934 B.n245 B.n150 10.6151
R935 B.n246 B.n245 10.6151
R936 B.n247 B.n246 10.6151
R937 B.n247 B.n148 10.6151
R938 B.n251 B.n148 10.6151
R939 B.n252 B.n251 10.6151
R940 B.n253 B.n252 10.6151
R941 B.n253 B.n146 10.6151
R942 B.n257 B.n146 10.6151
R943 B.n258 B.n257 10.6151
R944 B.n259 B.n258 10.6151
R945 B.n259 B.n144 10.6151
R946 B.n263 B.n144 10.6151
R947 B.n264 B.n263 10.6151
R948 B.n265 B.n264 10.6151
R949 B.n265 B.n142 10.6151
R950 B.n269 B.n142 10.6151
R951 B.n270 B.n269 10.6151
R952 B.n271 B.n270 10.6151
R953 B.n271 B.n140 10.6151
R954 B.n275 B.n140 10.6151
R955 B.n276 B.n275 10.6151
R956 B.n277 B.n276 10.6151
R957 B.n277 B.n138 10.6151
R958 B.n281 B.n138 10.6151
R959 B.n282 B.n281 10.6151
R960 B.n283 B.n282 10.6151
R961 B.n283 B.n136 10.6151
R962 B.n287 B.n136 10.6151
R963 B.n288 B.n287 10.6151
R964 B.n290 B.n132 10.6151
R965 B.n294 B.n132 10.6151
R966 B.n295 B.n294 10.6151
R967 B.n296 B.n295 10.6151
R968 B.n296 B.n130 10.6151
R969 B.n300 B.n130 10.6151
R970 B.n301 B.n300 10.6151
R971 B.n305 B.n301 10.6151
R972 B.n309 B.n128 10.6151
R973 B.n310 B.n309 10.6151
R974 B.n311 B.n310 10.6151
R975 B.n311 B.n126 10.6151
R976 B.n315 B.n126 10.6151
R977 B.n316 B.n315 10.6151
R978 B.n317 B.n316 10.6151
R979 B.n317 B.n124 10.6151
R980 B.n321 B.n124 10.6151
R981 B.n322 B.n321 10.6151
R982 B.n323 B.n322 10.6151
R983 B.n323 B.n122 10.6151
R984 B.n327 B.n122 10.6151
R985 B.n328 B.n327 10.6151
R986 B.n329 B.n328 10.6151
R987 B.n329 B.n120 10.6151
R988 B.n333 B.n120 10.6151
R989 B.n334 B.n333 10.6151
R990 B.n335 B.n334 10.6151
R991 B.n335 B.n118 10.6151
R992 B.n339 B.n118 10.6151
R993 B.n340 B.n339 10.6151
R994 B.n341 B.n340 10.6151
R995 B.n341 B.n116 10.6151
R996 B.n345 B.n116 10.6151
R997 B.n346 B.n345 10.6151
R998 B.n347 B.n346 10.6151
R999 B.n347 B.n114 10.6151
R1000 B.n351 B.n114 10.6151
R1001 B.n352 B.n351 10.6151
R1002 B.n353 B.n352 10.6151
R1003 B.n353 B.n112 10.6151
R1004 B.n357 B.n112 10.6151
R1005 B.n358 B.n357 10.6151
R1006 B.n359 B.n358 10.6151
R1007 B.n359 B.n110 10.6151
R1008 B.n363 B.n110 10.6151
R1009 B.n364 B.n363 10.6151
R1010 B.n365 B.n364 10.6151
R1011 B.n365 B.n108 10.6151
R1012 B.n369 B.n108 10.6151
R1013 B.n370 B.n369 10.6151
R1014 B.n677 B.n0 8.11757
R1015 B.n677 B.n1 8.11757
R1016 B.n558 B.n557 6.5566
R1017 B.n545 B.n544 6.5566
R1018 B.n290 B.n289 6.5566
R1019 B.n305 B.n304 6.5566
R1020 B.n559 B.n558 4.05904
R1021 B.n544 B.n543 4.05904
R1022 B.n289 B.n288 4.05904
R1023 B.n304 B.n128 4.05904
R1024 VP.n16 VP.n0 161.3
R1025 VP.n15 VP.n14 161.3
R1026 VP.n13 VP.n1 161.3
R1027 VP.n12 VP.n11 161.3
R1028 VP.n10 VP.n2 161.3
R1029 VP.n9 VP.n8 161.3
R1030 VP.n7 VP.n3 161.3
R1031 VP.n4 VP.t1 141.666
R1032 VP.n4 VP.t2 140.78
R1033 VP.n6 VP.n5 108.066
R1034 VP.n18 VP.n17 108.066
R1035 VP.n5 VP.t0 106.891
R1036 VP.n17 VP.t3 106.891
R1037 VP.n6 VP.n4 50.6101
R1038 VP.n11 VP.n10 40.4934
R1039 VP.n11 VP.n1 40.4934
R1040 VP.n9 VP.n3 24.4675
R1041 VP.n10 VP.n9 24.4675
R1042 VP.n15 VP.n1 24.4675
R1043 VP.n16 VP.n15 24.4675
R1044 VP.n5 VP.n3 2.69187
R1045 VP.n17 VP.n16 2.69187
R1046 VP.n7 VP.n6 0.278367
R1047 VP.n18 VP.n0 0.278367
R1048 VP.n8 VP.n7 0.189894
R1049 VP.n8 VP.n2 0.189894
R1050 VP.n12 VP.n2 0.189894
R1051 VP.n13 VP.n12 0.189894
R1052 VP.n14 VP.n13 0.189894
R1053 VP.n14 VP.n0 0.189894
R1054 VP VP.n18 0.153454
R1055 VDD1 VDD1.n1 120.007
R1056 VDD1 VDD1.n0 77.1531
R1057 VDD1.n0 VDD1.t2 2.63675
R1058 VDD1.n0 VDD1.t3 2.63675
R1059 VDD1.n1 VDD1.t1 2.63675
R1060 VDD1.n1 VDD1.t0 2.63675
R1061 VTAIL.n5 VTAIL.t5 63.0536
R1062 VTAIL.n4 VTAIL.t0 63.0536
R1063 VTAIL.n3 VTAIL.t7 63.0536
R1064 VTAIL.n7 VTAIL.t1 63.0525
R1065 VTAIL.n0 VTAIL.t2 63.0525
R1066 VTAIL.n1 VTAIL.t3 63.0525
R1067 VTAIL.n2 VTAIL.t6 63.0525
R1068 VTAIL.n6 VTAIL.t4 63.0524
R1069 VTAIL.n7 VTAIL.n6 25.6772
R1070 VTAIL.n3 VTAIL.n2 25.6772
R1071 VTAIL.n4 VTAIL.n3 2.68153
R1072 VTAIL.n6 VTAIL.n5 2.68153
R1073 VTAIL.n2 VTAIL.n1 2.68153
R1074 VTAIL VTAIL.n0 1.39921
R1075 VTAIL VTAIL.n7 1.28283
R1076 VTAIL.n5 VTAIL.n4 0.470328
R1077 VTAIL.n1 VTAIL.n0 0.470328
R1078 VN.n0 VN.t3 141.666
R1079 VN.n1 VN.t0 141.666
R1080 VN.n0 VN.t1 140.78
R1081 VN.n1 VN.t2 140.78
R1082 VN VN.n1 50.889
R1083 VN VN.n0 3.53673
R1084 VDD2.n2 VDD2.n0 119.484
R1085 VDD2.n2 VDD2.n1 77.0949
R1086 VDD2.n1 VDD2.t1 2.63675
R1087 VDD2.n1 VDD2.t3 2.63675
R1088 VDD2.n0 VDD2.t0 2.63675
R1089 VDD2.n0 VDD2.t2 2.63675
R1090 VDD2 VDD2.n2 0.0586897
C0 VP VDD1 5.18948f
C1 VN VDD2 4.93367f
C2 w_n2836_n3434# VDD1 1.49383f
C3 VP B 1.75333f
C4 B w_n2836_n3434# 9.55997f
C5 VDD1 VTAIL 5.51629f
C6 VP VN 6.38251f
C7 B VTAIL 5.1355f
C8 w_n2836_n3434# VN 4.84619f
C9 VP VDD2 0.405596f
C10 VN VTAIL 4.85012f
C11 w_n2836_n3434# VDD2 1.55394f
C12 VTAIL VDD2 5.57171f
C13 B VDD1 1.30171f
C14 VP w_n2836_n3434# 5.21123f
C15 VN VDD1 0.149f
C16 VP VTAIL 4.86423f
C17 B VN 1.14674f
C18 w_n2836_n3434# VTAIL 4.053f
C19 VDD1 VDD2 1.06458f
C20 B VDD2 1.35685f
C21 VDD2 VSUBS 0.987778f
C22 VDD1 VSUBS 5.86716f
C23 VTAIL VSUBS 1.251528f
C24 VN VSUBS 5.5445f
C25 VP VSUBS 2.382852f
C26 B VSUBS 4.459679f
C27 w_n2836_n3434# VSUBS 0.119827p
C28 VDD2.t0 VSUBS 0.261764f
C29 VDD2.t2 VSUBS 0.261764f
C30 VDD2.n0 VSUBS 2.77617f
C31 VDD2.t1 VSUBS 0.261764f
C32 VDD2.t3 VSUBS 0.261764f
C33 VDD2.n1 VSUBS 2.07746f
C34 VDD2.n2 VSUBS 4.36144f
C35 VN.t3 VSUBS 3.25591f
C36 VN.t1 VSUBS 3.24828f
C37 VN.n0 VSUBS 2.05518f
C38 VN.t0 VSUBS 3.25591f
C39 VN.t2 VSUBS 3.24828f
C40 VN.n1 VSUBS 3.84981f
C41 VTAIL.t2 VSUBS 2.26731f
C42 VTAIL.n0 VSUBS 0.742902f
C43 VTAIL.t3 VSUBS 2.26731f
C44 VTAIL.n1 VSUBS 0.841234f
C45 VTAIL.t6 VSUBS 2.26731f
C46 VTAIL.n2 VSUBS 2.14914f
C47 VTAIL.t7 VSUBS 2.26732f
C48 VTAIL.n3 VSUBS 2.14914f
C49 VTAIL.t0 VSUBS 2.26732f
C50 VTAIL.n4 VSUBS 0.841231f
C51 VTAIL.t5 VSUBS 2.26732f
C52 VTAIL.n5 VSUBS 0.841231f
C53 VTAIL.t4 VSUBS 2.26731f
C54 VTAIL.n6 VSUBS 2.14915f
C55 VTAIL.t1 VSUBS 2.26731f
C56 VTAIL.n7 VSUBS 2.04188f
C57 VDD1.t2 VSUBS 0.264253f
C58 VDD1.t3 VSUBS 0.264253f
C59 VDD1.n0 VSUBS 2.09777f
C60 VDD1.t1 VSUBS 0.264253f
C61 VDD1.t0 VSUBS 0.264253f
C62 VDD1.n1 VSUBS 2.82742f
C63 VP.n0 VSUBS 0.043058f
C64 VP.t3 VSUBS 3.05246f
C65 VP.n1 VSUBS 0.06491f
C66 VP.n2 VSUBS 0.032659f
C67 VP.n3 VSUBS 0.034121f
C68 VP.t2 VSUBS 3.36366f
C69 VP.t1 VSUBS 3.37156f
C70 VP.n4 VSUBS 3.96929f
C71 VP.t0 VSUBS 3.05246f
C72 VP.n5 VSUBS 1.18022f
C73 VP.n6 VSUBS 1.83427f
C74 VP.n7 VSUBS 0.043058f
C75 VP.n8 VSUBS 0.032659f
C76 VP.n9 VSUBS 0.060868f
C77 VP.n10 VSUBS 0.06491f
C78 VP.n11 VSUBS 0.026402f
C79 VP.n12 VSUBS 0.032659f
C80 VP.n13 VSUBS 0.032659f
C81 VP.n14 VSUBS 0.032659f
C82 VP.n15 VSUBS 0.060868f
C83 VP.n16 VSUBS 0.034121f
C84 VP.n17 VSUBS 1.18022f
C85 VP.n18 VSUBS 0.060784f
C86 B.n0 VSUBS 0.005798f
C87 B.n1 VSUBS 0.005798f
C88 B.n2 VSUBS 0.008575f
C89 B.n3 VSUBS 0.006571f
C90 B.n4 VSUBS 0.006571f
C91 B.n5 VSUBS 0.006571f
C92 B.n6 VSUBS 0.006571f
C93 B.n7 VSUBS 0.006571f
C94 B.n8 VSUBS 0.006571f
C95 B.n9 VSUBS 0.006571f
C96 B.n10 VSUBS 0.006571f
C97 B.n11 VSUBS 0.006571f
C98 B.n12 VSUBS 0.006571f
C99 B.n13 VSUBS 0.006571f
C100 B.n14 VSUBS 0.006571f
C101 B.n15 VSUBS 0.006571f
C102 B.n16 VSUBS 0.006571f
C103 B.n17 VSUBS 0.006571f
C104 B.n18 VSUBS 0.006571f
C105 B.n19 VSUBS 0.014578f
C106 B.n20 VSUBS 0.006571f
C107 B.n21 VSUBS 0.006571f
C108 B.n22 VSUBS 0.006571f
C109 B.n23 VSUBS 0.006571f
C110 B.n24 VSUBS 0.006571f
C111 B.n25 VSUBS 0.006571f
C112 B.n26 VSUBS 0.006571f
C113 B.n27 VSUBS 0.006571f
C114 B.n28 VSUBS 0.006571f
C115 B.n29 VSUBS 0.006571f
C116 B.n30 VSUBS 0.006571f
C117 B.n31 VSUBS 0.006571f
C118 B.n32 VSUBS 0.006571f
C119 B.n33 VSUBS 0.006571f
C120 B.n34 VSUBS 0.006571f
C121 B.n35 VSUBS 0.006571f
C122 B.n36 VSUBS 0.006571f
C123 B.n37 VSUBS 0.006571f
C124 B.n38 VSUBS 0.006571f
C125 B.n39 VSUBS 0.006571f
C126 B.n40 VSUBS 0.006571f
C127 B.n41 VSUBS 0.006571f
C128 B.t7 VSUBS 0.378295f
C129 B.t8 VSUBS 0.399255f
C130 B.t6 VSUBS 1.46983f
C131 B.n42 VSUBS 0.213156f
C132 B.n43 VSUBS 0.068128f
C133 B.n44 VSUBS 0.006571f
C134 B.n45 VSUBS 0.006571f
C135 B.n46 VSUBS 0.006571f
C136 B.n47 VSUBS 0.006571f
C137 B.t1 VSUBS 0.378287f
C138 B.t2 VSUBS 0.399248f
C139 B.t0 VSUBS 1.46983f
C140 B.n48 VSUBS 0.213163f
C141 B.n49 VSUBS 0.068135f
C142 B.n50 VSUBS 0.006571f
C143 B.n51 VSUBS 0.006571f
C144 B.n52 VSUBS 0.006571f
C145 B.n53 VSUBS 0.006571f
C146 B.n54 VSUBS 0.006571f
C147 B.n55 VSUBS 0.006571f
C148 B.n56 VSUBS 0.006571f
C149 B.n57 VSUBS 0.006571f
C150 B.n58 VSUBS 0.006571f
C151 B.n59 VSUBS 0.006571f
C152 B.n60 VSUBS 0.006571f
C153 B.n61 VSUBS 0.006571f
C154 B.n62 VSUBS 0.006571f
C155 B.n63 VSUBS 0.006571f
C156 B.n64 VSUBS 0.006571f
C157 B.n65 VSUBS 0.006571f
C158 B.n66 VSUBS 0.006571f
C159 B.n67 VSUBS 0.006571f
C160 B.n68 VSUBS 0.006571f
C161 B.n69 VSUBS 0.006571f
C162 B.n70 VSUBS 0.006571f
C163 B.n71 VSUBS 0.014578f
C164 B.n72 VSUBS 0.006571f
C165 B.n73 VSUBS 0.006571f
C166 B.n74 VSUBS 0.006571f
C167 B.n75 VSUBS 0.006571f
C168 B.n76 VSUBS 0.006571f
C169 B.n77 VSUBS 0.006571f
C170 B.n78 VSUBS 0.006571f
C171 B.n79 VSUBS 0.006571f
C172 B.n80 VSUBS 0.006571f
C173 B.n81 VSUBS 0.006571f
C174 B.n82 VSUBS 0.006571f
C175 B.n83 VSUBS 0.006571f
C176 B.n84 VSUBS 0.006571f
C177 B.n85 VSUBS 0.006571f
C178 B.n86 VSUBS 0.006571f
C179 B.n87 VSUBS 0.006571f
C180 B.n88 VSUBS 0.006571f
C181 B.n89 VSUBS 0.006571f
C182 B.n90 VSUBS 0.006571f
C183 B.n91 VSUBS 0.006571f
C184 B.n92 VSUBS 0.006571f
C185 B.n93 VSUBS 0.006571f
C186 B.n94 VSUBS 0.006571f
C187 B.n95 VSUBS 0.006571f
C188 B.n96 VSUBS 0.006571f
C189 B.n97 VSUBS 0.006571f
C190 B.n98 VSUBS 0.006571f
C191 B.n99 VSUBS 0.006571f
C192 B.n100 VSUBS 0.006571f
C193 B.n101 VSUBS 0.006571f
C194 B.n102 VSUBS 0.006571f
C195 B.n103 VSUBS 0.006571f
C196 B.n104 VSUBS 0.006571f
C197 B.n105 VSUBS 0.006571f
C198 B.n106 VSUBS 0.006571f
C199 B.n107 VSUBS 0.015573f
C200 B.n108 VSUBS 0.006571f
C201 B.n109 VSUBS 0.006571f
C202 B.n110 VSUBS 0.006571f
C203 B.n111 VSUBS 0.006571f
C204 B.n112 VSUBS 0.006571f
C205 B.n113 VSUBS 0.006571f
C206 B.n114 VSUBS 0.006571f
C207 B.n115 VSUBS 0.006571f
C208 B.n116 VSUBS 0.006571f
C209 B.n117 VSUBS 0.006571f
C210 B.n118 VSUBS 0.006571f
C211 B.n119 VSUBS 0.006571f
C212 B.n120 VSUBS 0.006571f
C213 B.n121 VSUBS 0.006571f
C214 B.n122 VSUBS 0.006571f
C215 B.n123 VSUBS 0.006571f
C216 B.n124 VSUBS 0.006571f
C217 B.n125 VSUBS 0.006571f
C218 B.n126 VSUBS 0.006571f
C219 B.n127 VSUBS 0.006571f
C220 B.n128 VSUBS 0.004542f
C221 B.n129 VSUBS 0.006571f
C222 B.n130 VSUBS 0.006571f
C223 B.n131 VSUBS 0.006571f
C224 B.n132 VSUBS 0.006571f
C225 B.n133 VSUBS 0.006571f
C226 B.t11 VSUBS 0.378295f
C227 B.t10 VSUBS 0.399255f
C228 B.t9 VSUBS 1.46983f
C229 B.n134 VSUBS 0.213156f
C230 B.n135 VSUBS 0.068128f
C231 B.n136 VSUBS 0.006571f
C232 B.n137 VSUBS 0.006571f
C233 B.n138 VSUBS 0.006571f
C234 B.n139 VSUBS 0.006571f
C235 B.n140 VSUBS 0.006571f
C236 B.n141 VSUBS 0.006571f
C237 B.n142 VSUBS 0.006571f
C238 B.n143 VSUBS 0.006571f
C239 B.n144 VSUBS 0.006571f
C240 B.n145 VSUBS 0.006571f
C241 B.n146 VSUBS 0.006571f
C242 B.n147 VSUBS 0.006571f
C243 B.n148 VSUBS 0.006571f
C244 B.n149 VSUBS 0.006571f
C245 B.n150 VSUBS 0.006571f
C246 B.n151 VSUBS 0.006571f
C247 B.n152 VSUBS 0.006571f
C248 B.n153 VSUBS 0.006571f
C249 B.n154 VSUBS 0.006571f
C250 B.n155 VSUBS 0.006571f
C251 B.n156 VSUBS 0.015573f
C252 B.n157 VSUBS 0.006571f
C253 B.n158 VSUBS 0.006571f
C254 B.n159 VSUBS 0.006571f
C255 B.n160 VSUBS 0.006571f
C256 B.n161 VSUBS 0.006571f
C257 B.n162 VSUBS 0.006571f
C258 B.n163 VSUBS 0.006571f
C259 B.n164 VSUBS 0.006571f
C260 B.n165 VSUBS 0.006571f
C261 B.n166 VSUBS 0.006571f
C262 B.n167 VSUBS 0.006571f
C263 B.n168 VSUBS 0.006571f
C264 B.n169 VSUBS 0.006571f
C265 B.n170 VSUBS 0.006571f
C266 B.n171 VSUBS 0.006571f
C267 B.n172 VSUBS 0.006571f
C268 B.n173 VSUBS 0.006571f
C269 B.n174 VSUBS 0.006571f
C270 B.n175 VSUBS 0.006571f
C271 B.n176 VSUBS 0.006571f
C272 B.n177 VSUBS 0.006571f
C273 B.n178 VSUBS 0.006571f
C274 B.n179 VSUBS 0.006571f
C275 B.n180 VSUBS 0.006571f
C276 B.n181 VSUBS 0.006571f
C277 B.n182 VSUBS 0.006571f
C278 B.n183 VSUBS 0.006571f
C279 B.n184 VSUBS 0.006571f
C280 B.n185 VSUBS 0.006571f
C281 B.n186 VSUBS 0.006571f
C282 B.n187 VSUBS 0.006571f
C283 B.n188 VSUBS 0.006571f
C284 B.n189 VSUBS 0.006571f
C285 B.n190 VSUBS 0.006571f
C286 B.n191 VSUBS 0.006571f
C287 B.n192 VSUBS 0.006571f
C288 B.n193 VSUBS 0.006571f
C289 B.n194 VSUBS 0.006571f
C290 B.n195 VSUBS 0.006571f
C291 B.n196 VSUBS 0.006571f
C292 B.n197 VSUBS 0.006571f
C293 B.n198 VSUBS 0.006571f
C294 B.n199 VSUBS 0.006571f
C295 B.n200 VSUBS 0.006571f
C296 B.n201 VSUBS 0.006571f
C297 B.n202 VSUBS 0.006571f
C298 B.n203 VSUBS 0.006571f
C299 B.n204 VSUBS 0.006571f
C300 B.n205 VSUBS 0.006571f
C301 B.n206 VSUBS 0.006571f
C302 B.n207 VSUBS 0.006571f
C303 B.n208 VSUBS 0.006571f
C304 B.n209 VSUBS 0.006571f
C305 B.n210 VSUBS 0.006571f
C306 B.n211 VSUBS 0.006571f
C307 B.n212 VSUBS 0.006571f
C308 B.n213 VSUBS 0.006571f
C309 B.n214 VSUBS 0.006571f
C310 B.n215 VSUBS 0.006571f
C311 B.n216 VSUBS 0.006571f
C312 B.n217 VSUBS 0.006571f
C313 B.n218 VSUBS 0.006571f
C314 B.n219 VSUBS 0.006571f
C315 B.n220 VSUBS 0.006571f
C316 B.n221 VSUBS 0.006571f
C317 B.n222 VSUBS 0.006571f
C318 B.n223 VSUBS 0.014578f
C319 B.n224 VSUBS 0.014578f
C320 B.n225 VSUBS 0.015573f
C321 B.n226 VSUBS 0.006571f
C322 B.n227 VSUBS 0.006571f
C323 B.n228 VSUBS 0.006571f
C324 B.n229 VSUBS 0.006571f
C325 B.n230 VSUBS 0.006571f
C326 B.n231 VSUBS 0.006571f
C327 B.n232 VSUBS 0.006571f
C328 B.n233 VSUBS 0.006571f
C329 B.n234 VSUBS 0.006571f
C330 B.n235 VSUBS 0.006571f
C331 B.n236 VSUBS 0.006571f
C332 B.n237 VSUBS 0.006571f
C333 B.n238 VSUBS 0.006571f
C334 B.n239 VSUBS 0.006571f
C335 B.n240 VSUBS 0.006571f
C336 B.n241 VSUBS 0.006571f
C337 B.n242 VSUBS 0.006571f
C338 B.n243 VSUBS 0.006571f
C339 B.n244 VSUBS 0.006571f
C340 B.n245 VSUBS 0.006571f
C341 B.n246 VSUBS 0.006571f
C342 B.n247 VSUBS 0.006571f
C343 B.n248 VSUBS 0.006571f
C344 B.n249 VSUBS 0.006571f
C345 B.n250 VSUBS 0.006571f
C346 B.n251 VSUBS 0.006571f
C347 B.n252 VSUBS 0.006571f
C348 B.n253 VSUBS 0.006571f
C349 B.n254 VSUBS 0.006571f
C350 B.n255 VSUBS 0.006571f
C351 B.n256 VSUBS 0.006571f
C352 B.n257 VSUBS 0.006571f
C353 B.n258 VSUBS 0.006571f
C354 B.n259 VSUBS 0.006571f
C355 B.n260 VSUBS 0.006571f
C356 B.n261 VSUBS 0.006571f
C357 B.n262 VSUBS 0.006571f
C358 B.n263 VSUBS 0.006571f
C359 B.n264 VSUBS 0.006571f
C360 B.n265 VSUBS 0.006571f
C361 B.n266 VSUBS 0.006571f
C362 B.n267 VSUBS 0.006571f
C363 B.n268 VSUBS 0.006571f
C364 B.n269 VSUBS 0.006571f
C365 B.n270 VSUBS 0.006571f
C366 B.n271 VSUBS 0.006571f
C367 B.n272 VSUBS 0.006571f
C368 B.n273 VSUBS 0.006571f
C369 B.n274 VSUBS 0.006571f
C370 B.n275 VSUBS 0.006571f
C371 B.n276 VSUBS 0.006571f
C372 B.n277 VSUBS 0.006571f
C373 B.n278 VSUBS 0.006571f
C374 B.n279 VSUBS 0.006571f
C375 B.n280 VSUBS 0.006571f
C376 B.n281 VSUBS 0.006571f
C377 B.n282 VSUBS 0.006571f
C378 B.n283 VSUBS 0.006571f
C379 B.n284 VSUBS 0.006571f
C380 B.n285 VSUBS 0.006571f
C381 B.n286 VSUBS 0.006571f
C382 B.n287 VSUBS 0.006571f
C383 B.n288 VSUBS 0.004542f
C384 B.n289 VSUBS 0.015225f
C385 B.n290 VSUBS 0.005315f
C386 B.n291 VSUBS 0.006571f
C387 B.n292 VSUBS 0.006571f
C388 B.n293 VSUBS 0.006571f
C389 B.n294 VSUBS 0.006571f
C390 B.n295 VSUBS 0.006571f
C391 B.n296 VSUBS 0.006571f
C392 B.n297 VSUBS 0.006571f
C393 B.n298 VSUBS 0.006571f
C394 B.n299 VSUBS 0.006571f
C395 B.n300 VSUBS 0.006571f
C396 B.n301 VSUBS 0.006571f
C397 B.t5 VSUBS 0.378287f
C398 B.t4 VSUBS 0.399248f
C399 B.t3 VSUBS 1.46983f
C400 B.n302 VSUBS 0.213163f
C401 B.n303 VSUBS 0.068135f
C402 B.n304 VSUBS 0.015225f
C403 B.n305 VSUBS 0.005315f
C404 B.n306 VSUBS 0.006571f
C405 B.n307 VSUBS 0.006571f
C406 B.n308 VSUBS 0.006571f
C407 B.n309 VSUBS 0.006571f
C408 B.n310 VSUBS 0.006571f
C409 B.n311 VSUBS 0.006571f
C410 B.n312 VSUBS 0.006571f
C411 B.n313 VSUBS 0.006571f
C412 B.n314 VSUBS 0.006571f
C413 B.n315 VSUBS 0.006571f
C414 B.n316 VSUBS 0.006571f
C415 B.n317 VSUBS 0.006571f
C416 B.n318 VSUBS 0.006571f
C417 B.n319 VSUBS 0.006571f
C418 B.n320 VSUBS 0.006571f
C419 B.n321 VSUBS 0.006571f
C420 B.n322 VSUBS 0.006571f
C421 B.n323 VSUBS 0.006571f
C422 B.n324 VSUBS 0.006571f
C423 B.n325 VSUBS 0.006571f
C424 B.n326 VSUBS 0.006571f
C425 B.n327 VSUBS 0.006571f
C426 B.n328 VSUBS 0.006571f
C427 B.n329 VSUBS 0.006571f
C428 B.n330 VSUBS 0.006571f
C429 B.n331 VSUBS 0.006571f
C430 B.n332 VSUBS 0.006571f
C431 B.n333 VSUBS 0.006571f
C432 B.n334 VSUBS 0.006571f
C433 B.n335 VSUBS 0.006571f
C434 B.n336 VSUBS 0.006571f
C435 B.n337 VSUBS 0.006571f
C436 B.n338 VSUBS 0.006571f
C437 B.n339 VSUBS 0.006571f
C438 B.n340 VSUBS 0.006571f
C439 B.n341 VSUBS 0.006571f
C440 B.n342 VSUBS 0.006571f
C441 B.n343 VSUBS 0.006571f
C442 B.n344 VSUBS 0.006571f
C443 B.n345 VSUBS 0.006571f
C444 B.n346 VSUBS 0.006571f
C445 B.n347 VSUBS 0.006571f
C446 B.n348 VSUBS 0.006571f
C447 B.n349 VSUBS 0.006571f
C448 B.n350 VSUBS 0.006571f
C449 B.n351 VSUBS 0.006571f
C450 B.n352 VSUBS 0.006571f
C451 B.n353 VSUBS 0.006571f
C452 B.n354 VSUBS 0.006571f
C453 B.n355 VSUBS 0.006571f
C454 B.n356 VSUBS 0.006571f
C455 B.n357 VSUBS 0.006571f
C456 B.n358 VSUBS 0.006571f
C457 B.n359 VSUBS 0.006571f
C458 B.n360 VSUBS 0.006571f
C459 B.n361 VSUBS 0.006571f
C460 B.n362 VSUBS 0.006571f
C461 B.n363 VSUBS 0.006571f
C462 B.n364 VSUBS 0.006571f
C463 B.n365 VSUBS 0.006571f
C464 B.n366 VSUBS 0.006571f
C465 B.n367 VSUBS 0.006571f
C466 B.n368 VSUBS 0.006571f
C467 B.n369 VSUBS 0.006571f
C468 B.n370 VSUBS 0.014773f
C469 B.n371 VSUBS 0.015378f
C470 B.n372 VSUBS 0.014578f
C471 B.n373 VSUBS 0.006571f
C472 B.n374 VSUBS 0.006571f
C473 B.n375 VSUBS 0.006571f
C474 B.n376 VSUBS 0.006571f
C475 B.n377 VSUBS 0.006571f
C476 B.n378 VSUBS 0.006571f
C477 B.n379 VSUBS 0.006571f
C478 B.n380 VSUBS 0.006571f
C479 B.n381 VSUBS 0.006571f
C480 B.n382 VSUBS 0.006571f
C481 B.n383 VSUBS 0.006571f
C482 B.n384 VSUBS 0.006571f
C483 B.n385 VSUBS 0.006571f
C484 B.n386 VSUBS 0.006571f
C485 B.n387 VSUBS 0.006571f
C486 B.n388 VSUBS 0.006571f
C487 B.n389 VSUBS 0.006571f
C488 B.n390 VSUBS 0.006571f
C489 B.n391 VSUBS 0.006571f
C490 B.n392 VSUBS 0.006571f
C491 B.n393 VSUBS 0.006571f
C492 B.n394 VSUBS 0.006571f
C493 B.n395 VSUBS 0.006571f
C494 B.n396 VSUBS 0.006571f
C495 B.n397 VSUBS 0.006571f
C496 B.n398 VSUBS 0.006571f
C497 B.n399 VSUBS 0.006571f
C498 B.n400 VSUBS 0.006571f
C499 B.n401 VSUBS 0.006571f
C500 B.n402 VSUBS 0.006571f
C501 B.n403 VSUBS 0.006571f
C502 B.n404 VSUBS 0.006571f
C503 B.n405 VSUBS 0.006571f
C504 B.n406 VSUBS 0.006571f
C505 B.n407 VSUBS 0.006571f
C506 B.n408 VSUBS 0.006571f
C507 B.n409 VSUBS 0.006571f
C508 B.n410 VSUBS 0.006571f
C509 B.n411 VSUBS 0.006571f
C510 B.n412 VSUBS 0.006571f
C511 B.n413 VSUBS 0.006571f
C512 B.n414 VSUBS 0.006571f
C513 B.n415 VSUBS 0.006571f
C514 B.n416 VSUBS 0.006571f
C515 B.n417 VSUBS 0.006571f
C516 B.n418 VSUBS 0.006571f
C517 B.n419 VSUBS 0.006571f
C518 B.n420 VSUBS 0.006571f
C519 B.n421 VSUBS 0.006571f
C520 B.n422 VSUBS 0.006571f
C521 B.n423 VSUBS 0.006571f
C522 B.n424 VSUBS 0.006571f
C523 B.n425 VSUBS 0.006571f
C524 B.n426 VSUBS 0.006571f
C525 B.n427 VSUBS 0.006571f
C526 B.n428 VSUBS 0.006571f
C527 B.n429 VSUBS 0.006571f
C528 B.n430 VSUBS 0.006571f
C529 B.n431 VSUBS 0.006571f
C530 B.n432 VSUBS 0.006571f
C531 B.n433 VSUBS 0.006571f
C532 B.n434 VSUBS 0.006571f
C533 B.n435 VSUBS 0.006571f
C534 B.n436 VSUBS 0.006571f
C535 B.n437 VSUBS 0.006571f
C536 B.n438 VSUBS 0.006571f
C537 B.n439 VSUBS 0.006571f
C538 B.n440 VSUBS 0.006571f
C539 B.n441 VSUBS 0.006571f
C540 B.n442 VSUBS 0.006571f
C541 B.n443 VSUBS 0.006571f
C542 B.n444 VSUBS 0.006571f
C543 B.n445 VSUBS 0.006571f
C544 B.n446 VSUBS 0.006571f
C545 B.n447 VSUBS 0.006571f
C546 B.n448 VSUBS 0.006571f
C547 B.n449 VSUBS 0.006571f
C548 B.n450 VSUBS 0.006571f
C549 B.n451 VSUBS 0.006571f
C550 B.n452 VSUBS 0.006571f
C551 B.n453 VSUBS 0.006571f
C552 B.n454 VSUBS 0.006571f
C553 B.n455 VSUBS 0.006571f
C554 B.n456 VSUBS 0.006571f
C555 B.n457 VSUBS 0.006571f
C556 B.n458 VSUBS 0.006571f
C557 B.n459 VSUBS 0.006571f
C558 B.n460 VSUBS 0.006571f
C559 B.n461 VSUBS 0.006571f
C560 B.n462 VSUBS 0.006571f
C561 B.n463 VSUBS 0.006571f
C562 B.n464 VSUBS 0.006571f
C563 B.n465 VSUBS 0.006571f
C564 B.n466 VSUBS 0.006571f
C565 B.n467 VSUBS 0.006571f
C566 B.n468 VSUBS 0.006571f
C567 B.n469 VSUBS 0.006571f
C568 B.n470 VSUBS 0.006571f
C569 B.n471 VSUBS 0.006571f
C570 B.n472 VSUBS 0.006571f
C571 B.n473 VSUBS 0.006571f
C572 B.n474 VSUBS 0.006571f
C573 B.n475 VSUBS 0.006571f
C574 B.n476 VSUBS 0.006571f
C575 B.n477 VSUBS 0.006571f
C576 B.n478 VSUBS 0.014578f
C577 B.n479 VSUBS 0.015573f
C578 B.n480 VSUBS 0.015573f
C579 B.n481 VSUBS 0.006571f
C580 B.n482 VSUBS 0.006571f
C581 B.n483 VSUBS 0.006571f
C582 B.n484 VSUBS 0.006571f
C583 B.n485 VSUBS 0.006571f
C584 B.n486 VSUBS 0.006571f
C585 B.n487 VSUBS 0.006571f
C586 B.n488 VSUBS 0.006571f
C587 B.n489 VSUBS 0.006571f
C588 B.n490 VSUBS 0.006571f
C589 B.n491 VSUBS 0.006571f
C590 B.n492 VSUBS 0.006571f
C591 B.n493 VSUBS 0.006571f
C592 B.n494 VSUBS 0.006571f
C593 B.n495 VSUBS 0.006571f
C594 B.n496 VSUBS 0.006571f
C595 B.n497 VSUBS 0.006571f
C596 B.n498 VSUBS 0.006571f
C597 B.n499 VSUBS 0.006571f
C598 B.n500 VSUBS 0.006571f
C599 B.n501 VSUBS 0.006571f
C600 B.n502 VSUBS 0.006571f
C601 B.n503 VSUBS 0.006571f
C602 B.n504 VSUBS 0.006571f
C603 B.n505 VSUBS 0.006571f
C604 B.n506 VSUBS 0.006571f
C605 B.n507 VSUBS 0.006571f
C606 B.n508 VSUBS 0.006571f
C607 B.n509 VSUBS 0.006571f
C608 B.n510 VSUBS 0.006571f
C609 B.n511 VSUBS 0.006571f
C610 B.n512 VSUBS 0.006571f
C611 B.n513 VSUBS 0.006571f
C612 B.n514 VSUBS 0.006571f
C613 B.n515 VSUBS 0.006571f
C614 B.n516 VSUBS 0.006571f
C615 B.n517 VSUBS 0.006571f
C616 B.n518 VSUBS 0.006571f
C617 B.n519 VSUBS 0.006571f
C618 B.n520 VSUBS 0.006571f
C619 B.n521 VSUBS 0.006571f
C620 B.n522 VSUBS 0.006571f
C621 B.n523 VSUBS 0.006571f
C622 B.n524 VSUBS 0.006571f
C623 B.n525 VSUBS 0.006571f
C624 B.n526 VSUBS 0.006571f
C625 B.n527 VSUBS 0.006571f
C626 B.n528 VSUBS 0.006571f
C627 B.n529 VSUBS 0.006571f
C628 B.n530 VSUBS 0.006571f
C629 B.n531 VSUBS 0.006571f
C630 B.n532 VSUBS 0.006571f
C631 B.n533 VSUBS 0.006571f
C632 B.n534 VSUBS 0.006571f
C633 B.n535 VSUBS 0.006571f
C634 B.n536 VSUBS 0.006571f
C635 B.n537 VSUBS 0.006571f
C636 B.n538 VSUBS 0.006571f
C637 B.n539 VSUBS 0.006571f
C638 B.n540 VSUBS 0.006571f
C639 B.n541 VSUBS 0.006571f
C640 B.n542 VSUBS 0.006571f
C641 B.n543 VSUBS 0.004542f
C642 B.n544 VSUBS 0.015225f
C643 B.n545 VSUBS 0.005315f
C644 B.n546 VSUBS 0.006571f
C645 B.n547 VSUBS 0.006571f
C646 B.n548 VSUBS 0.006571f
C647 B.n549 VSUBS 0.006571f
C648 B.n550 VSUBS 0.006571f
C649 B.n551 VSUBS 0.006571f
C650 B.n552 VSUBS 0.006571f
C651 B.n553 VSUBS 0.006571f
C652 B.n554 VSUBS 0.006571f
C653 B.n555 VSUBS 0.006571f
C654 B.n556 VSUBS 0.006571f
C655 B.n557 VSUBS 0.005315f
C656 B.n558 VSUBS 0.015225f
C657 B.n559 VSUBS 0.004542f
C658 B.n560 VSUBS 0.006571f
C659 B.n561 VSUBS 0.006571f
C660 B.n562 VSUBS 0.006571f
C661 B.n563 VSUBS 0.006571f
C662 B.n564 VSUBS 0.006571f
C663 B.n565 VSUBS 0.006571f
C664 B.n566 VSUBS 0.006571f
C665 B.n567 VSUBS 0.006571f
C666 B.n568 VSUBS 0.006571f
C667 B.n569 VSUBS 0.006571f
C668 B.n570 VSUBS 0.006571f
C669 B.n571 VSUBS 0.006571f
C670 B.n572 VSUBS 0.006571f
C671 B.n573 VSUBS 0.006571f
C672 B.n574 VSUBS 0.006571f
C673 B.n575 VSUBS 0.006571f
C674 B.n576 VSUBS 0.006571f
C675 B.n577 VSUBS 0.006571f
C676 B.n578 VSUBS 0.006571f
C677 B.n579 VSUBS 0.006571f
C678 B.n580 VSUBS 0.006571f
C679 B.n581 VSUBS 0.006571f
C680 B.n582 VSUBS 0.006571f
C681 B.n583 VSUBS 0.006571f
C682 B.n584 VSUBS 0.006571f
C683 B.n585 VSUBS 0.006571f
C684 B.n586 VSUBS 0.006571f
C685 B.n587 VSUBS 0.006571f
C686 B.n588 VSUBS 0.006571f
C687 B.n589 VSUBS 0.006571f
C688 B.n590 VSUBS 0.006571f
C689 B.n591 VSUBS 0.006571f
C690 B.n592 VSUBS 0.006571f
C691 B.n593 VSUBS 0.006571f
C692 B.n594 VSUBS 0.006571f
C693 B.n595 VSUBS 0.006571f
C694 B.n596 VSUBS 0.006571f
C695 B.n597 VSUBS 0.006571f
C696 B.n598 VSUBS 0.006571f
C697 B.n599 VSUBS 0.006571f
C698 B.n600 VSUBS 0.006571f
C699 B.n601 VSUBS 0.006571f
C700 B.n602 VSUBS 0.006571f
C701 B.n603 VSUBS 0.006571f
C702 B.n604 VSUBS 0.006571f
C703 B.n605 VSUBS 0.006571f
C704 B.n606 VSUBS 0.006571f
C705 B.n607 VSUBS 0.006571f
C706 B.n608 VSUBS 0.006571f
C707 B.n609 VSUBS 0.006571f
C708 B.n610 VSUBS 0.006571f
C709 B.n611 VSUBS 0.006571f
C710 B.n612 VSUBS 0.006571f
C711 B.n613 VSUBS 0.006571f
C712 B.n614 VSUBS 0.006571f
C713 B.n615 VSUBS 0.006571f
C714 B.n616 VSUBS 0.006571f
C715 B.n617 VSUBS 0.006571f
C716 B.n618 VSUBS 0.006571f
C717 B.n619 VSUBS 0.006571f
C718 B.n620 VSUBS 0.006571f
C719 B.n621 VSUBS 0.006571f
C720 B.n622 VSUBS 0.015573f
C721 B.n623 VSUBS 0.015573f
C722 B.n624 VSUBS 0.014578f
C723 B.n625 VSUBS 0.006571f
C724 B.n626 VSUBS 0.006571f
C725 B.n627 VSUBS 0.006571f
C726 B.n628 VSUBS 0.006571f
C727 B.n629 VSUBS 0.006571f
C728 B.n630 VSUBS 0.006571f
C729 B.n631 VSUBS 0.006571f
C730 B.n632 VSUBS 0.006571f
C731 B.n633 VSUBS 0.006571f
C732 B.n634 VSUBS 0.006571f
C733 B.n635 VSUBS 0.006571f
C734 B.n636 VSUBS 0.006571f
C735 B.n637 VSUBS 0.006571f
C736 B.n638 VSUBS 0.006571f
C737 B.n639 VSUBS 0.006571f
C738 B.n640 VSUBS 0.006571f
C739 B.n641 VSUBS 0.006571f
C740 B.n642 VSUBS 0.006571f
C741 B.n643 VSUBS 0.006571f
C742 B.n644 VSUBS 0.006571f
C743 B.n645 VSUBS 0.006571f
C744 B.n646 VSUBS 0.006571f
C745 B.n647 VSUBS 0.006571f
C746 B.n648 VSUBS 0.006571f
C747 B.n649 VSUBS 0.006571f
C748 B.n650 VSUBS 0.006571f
C749 B.n651 VSUBS 0.006571f
C750 B.n652 VSUBS 0.006571f
C751 B.n653 VSUBS 0.006571f
C752 B.n654 VSUBS 0.006571f
C753 B.n655 VSUBS 0.006571f
C754 B.n656 VSUBS 0.006571f
C755 B.n657 VSUBS 0.006571f
C756 B.n658 VSUBS 0.006571f
C757 B.n659 VSUBS 0.006571f
C758 B.n660 VSUBS 0.006571f
C759 B.n661 VSUBS 0.006571f
C760 B.n662 VSUBS 0.006571f
C761 B.n663 VSUBS 0.006571f
C762 B.n664 VSUBS 0.006571f
C763 B.n665 VSUBS 0.006571f
C764 B.n666 VSUBS 0.006571f
C765 B.n667 VSUBS 0.006571f
C766 B.n668 VSUBS 0.006571f
C767 B.n669 VSUBS 0.006571f
C768 B.n670 VSUBS 0.006571f
C769 B.n671 VSUBS 0.006571f
C770 B.n672 VSUBS 0.006571f
C771 B.n673 VSUBS 0.006571f
C772 B.n674 VSUBS 0.006571f
C773 B.n675 VSUBS 0.008575f
C774 B.n676 VSUBS 0.009135f
C775 B.n677 VSUBS 0.018166f
.ends

