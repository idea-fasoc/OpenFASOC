* NGSPICE file created from diff_pair_sample_1531.ext - technology: sky130A

.subckt diff_pair_sample_1531 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t4 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=2.04
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=2.04
X2 B.t11 B.t9 B.t10 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=2.04
X3 VDD1.t4 VP.t1 VTAIL.t3 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=2.04
X4 VDD2.t0 VN.t1 VTAIL.t10 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=2.04
X5 VDD2.t5 VN.t2 VTAIL.t9 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=2.04
X6 B.t8 B.t6 B.t7 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=2.04
X7 VTAIL.t4 VP.t2 VDD1.t3 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=2.04
X8 VDD2.t1 VN.t3 VTAIL.t8 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=2.04
X9 VTAIL.t7 VN.t4 VDD2.t3 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=2.04
X10 VDD1.t2 VP.t3 VTAIL.t1 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0.6765 ps=4.43 w=4.1 l=2.04
X11 B.t5 B.t3 B.t4 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=2.04
X12 B.t2 B.t0 B.t1 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=1.599 pd=8.98 as=0 ps=0 w=4.1 l=2.04
X13 VDD1.t1 VP.t4 VTAIL.t0 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=2.04
X14 VDD2.t2 VN.t5 VTAIL.t6 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=1.599 ps=8.98 w=4.1 l=2.04
X15 VTAIL.t2 VP.t5 VDD1.t0 w_n2866_n1788# sky130_fd_pr__pfet_01v8 ad=0.6765 pd=4.43 as=0.6765 ps=4.43 w=4.1 l=2.04
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n11 VN.n10 92.7103
R9 VN.n23 VN.n22 92.7103
R10 VN.n2 VN.t2 82.34
R11 VN.n14 VN.t3 82.34
R12 VN.n8 VN.n1 56.5617
R13 VN.n20 VN.n13 56.5617
R14 VN.n3 VN.t0 48.4368
R15 VN.n10 VN.t5 48.4368
R16 VN.n15 VN.t4 48.4368
R17 VN.n22 VN.t1 48.4368
R18 VN.n15 VN.n14 45.9982
R19 VN.n3 VN.n2 45.9982
R20 VN VN.n23 40.7823
R21 VN.n4 VN.n3 24.5923
R22 VN.n4 VN.n1 24.5923
R23 VN.n9 VN.n8 24.5923
R24 VN.n16 VN.n13 24.5923
R25 VN.n16 VN.n15 24.5923
R26 VN.n21 VN.n20 24.5923
R27 VN.n10 VN.n9 18.1985
R28 VN.n22 VN.n21 18.1985
R29 VN.n17 VN.n14 9.12552
R30 VN.n5 VN.n2 9.12552
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VDD2.n1 VDD2.t5 115.853
R41 VDD2.n2 VDD2.t0 114.376
R42 VDD2.n1 VDD2.n0 106.903
R43 VDD2 VDD2.n3 106.9
R44 VDD2.n2 VDD2.n1 33.8899
R45 VDD2.n3 VDD2.t3 7.92855
R46 VDD2.n3 VDD2.t1 7.92855
R47 VDD2.n0 VDD2.t4 7.92855
R48 VDD2.n0 VDD2.t2 7.92855
R49 VDD2 VDD2.n2 1.59102
R50 VTAIL.n7 VTAIL.t8 97.6965
R51 VTAIL.n11 VTAIL.t6 97.6963
R52 VTAIL.n2 VTAIL.t0 97.6963
R53 VTAIL.n10 VTAIL.t3 97.6963
R54 VTAIL.n9 VTAIL.n8 89.7684
R55 VTAIL.n6 VTAIL.n5 89.7684
R56 VTAIL.n1 VTAIL.n0 89.7682
R57 VTAIL.n4 VTAIL.n3 89.7682
R58 VTAIL.n6 VTAIL.n4 19.9876
R59 VTAIL.n11 VTAIL.n10 17.9445
R60 VTAIL.n0 VTAIL.t9 7.92855
R61 VTAIL.n0 VTAIL.t11 7.92855
R62 VTAIL.n3 VTAIL.t5 7.92855
R63 VTAIL.n3 VTAIL.t2 7.92855
R64 VTAIL.n8 VTAIL.t1 7.92855
R65 VTAIL.n8 VTAIL.t4 7.92855
R66 VTAIL.n5 VTAIL.t10 7.92855
R67 VTAIL.n5 VTAIL.t7 7.92855
R68 VTAIL.n7 VTAIL.n6 2.0436
R69 VTAIL.n10 VTAIL.n9 2.0436
R70 VTAIL.n4 VTAIL.n2 2.0436
R71 VTAIL.n9 VTAIL.n7 1.49188
R72 VTAIL.n2 VTAIL.n1 1.49188
R73 VTAIL VTAIL.n11 1.47464
R74 VTAIL VTAIL.n1 0.569465
R75 VP.n10 VP.n9 161.3
R76 VP.n11 VP.n6 161.3
R77 VP.n13 VP.n12 161.3
R78 VP.n14 VP.n5 161.3
R79 VP.n31 VP.n0 161.3
R80 VP.n30 VP.n29 161.3
R81 VP.n28 VP.n1 161.3
R82 VP.n27 VP.n26 161.3
R83 VP.n25 VP.n2 161.3
R84 VP.n24 VP.n23 161.3
R85 VP.n22 VP.n3 161.3
R86 VP.n21 VP.n20 161.3
R87 VP.n19 VP.n4 161.3
R88 VP.n18 VP.n17 92.7103
R89 VP.n33 VP.n32 92.7103
R90 VP.n16 VP.n15 92.7103
R91 VP.n7 VP.t3 82.34
R92 VP.n20 VP.n3 56.5617
R93 VP.n30 VP.n1 56.5617
R94 VP.n13 VP.n6 56.5617
R95 VP.n25 VP.t5 48.4368
R96 VP.n18 VP.t0 48.4368
R97 VP.n32 VP.t4 48.4368
R98 VP.n8 VP.t2 48.4368
R99 VP.n15 VP.t1 48.4368
R100 VP.n8 VP.n7 45.9982
R101 VP.n17 VP.n16 40.5034
R102 VP.n20 VP.n19 24.5923
R103 VP.n24 VP.n3 24.5923
R104 VP.n25 VP.n24 24.5923
R105 VP.n26 VP.n25 24.5923
R106 VP.n26 VP.n1 24.5923
R107 VP.n31 VP.n30 24.5923
R108 VP.n14 VP.n13 24.5923
R109 VP.n9 VP.n8 24.5923
R110 VP.n9 VP.n6 24.5923
R111 VP.n19 VP.n18 18.1985
R112 VP.n32 VP.n31 18.1985
R113 VP.n15 VP.n14 18.1985
R114 VP.n10 VP.n7 9.12552
R115 VP.n16 VP.n5 0.278335
R116 VP.n17 VP.n4 0.278335
R117 VP.n33 VP.n0 0.278335
R118 VP.n11 VP.n10 0.189894
R119 VP.n12 VP.n11 0.189894
R120 VP.n12 VP.n5 0.189894
R121 VP.n21 VP.n4 0.189894
R122 VP.n22 VP.n21 0.189894
R123 VP.n23 VP.n22 0.189894
R124 VP.n23 VP.n2 0.189894
R125 VP.n27 VP.n2 0.189894
R126 VP.n28 VP.n27 0.189894
R127 VP.n29 VP.n28 0.189894
R128 VP.n29 VP.n0 0.189894
R129 VP VP.n33 0.153485
R130 VDD1 VDD1.t2 115.966
R131 VDD1.n1 VDD1.t5 115.853
R132 VDD1.n1 VDD1.n0 106.903
R133 VDD1.n3 VDD1.n2 106.448
R134 VDD1.n3 VDD1.n1 35.4944
R135 VDD1.n2 VDD1.t3 7.92855
R136 VDD1.n2 VDD1.t4 7.92855
R137 VDD1.n0 VDD1.t0 7.92855
R138 VDD1.n0 VDD1.t1 7.92855
R139 VDD1 VDD1.n3 0.453086
R140 B.n362 B.n47 585
R141 B.n364 B.n363 585
R142 B.n365 B.n46 585
R143 B.n367 B.n366 585
R144 B.n368 B.n45 585
R145 B.n370 B.n369 585
R146 B.n371 B.n44 585
R147 B.n373 B.n372 585
R148 B.n374 B.n43 585
R149 B.n376 B.n375 585
R150 B.n377 B.n42 585
R151 B.n379 B.n378 585
R152 B.n380 B.n41 585
R153 B.n382 B.n381 585
R154 B.n383 B.n40 585
R155 B.n385 B.n384 585
R156 B.n386 B.n39 585
R157 B.n388 B.n387 585
R158 B.n390 B.n389 585
R159 B.n391 B.n35 585
R160 B.n393 B.n392 585
R161 B.n394 B.n34 585
R162 B.n396 B.n395 585
R163 B.n397 B.n33 585
R164 B.n399 B.n398 585
R165 B.n400 B.n32 585
R166 B.n402 B.n401 585
R167 B.n403 B.n29 585
R168 B.n406 B.n405 585
R169 B.n407 B.n28 585
R170 B.n409 B.n408 585
R171 B.n410 B.n27 585
R172 B.n412 B.n411 585
R173 B.n413 B.n26 585
R174 B.n415 B.n414 585
R175 B.n416 B.n25 585
R176 B.n418 B.n417 585
R177 B.n419 B.n24 585
R178 B.n421 B.n420 585
R179 B.n422 B.n23 585
R180 B.n424 B.n423 585
R181 B.n425 B.n22 585
R182 B.n427 B.n426 585
R183 B.n428 B.n21 585
R184 B.n430 B.n429 585
R185 B.n431 B.n20 585
R186 B.n361 B.n360 585
R187 B.n359 B.n48 585
R188 B.n358 B.n357 585
R189 B.n356 B.n49 585
R190 B.n355 B.n354 585
R191 B.n353 B.n50 585
R192 B.n352 B.n351 585
R193 B.n350 B.n51 585
R194 B.n349 B.n348 585
R195 B.n347 B.n52 585
R196 B.n346 B.n345 585
R197 B.n344 B.n53 585
R198 B.n343 B.n342 585
R199 B.n341 B.n54 585
R200 B.n340 B.n339 585
R201 B.n338 B.n55 585
R202 B.n337 B.n336 585
R203 B.n335 B.n56 585
R204 B.n334 B.n333 585
R205 B.n332 B.n57 585
R206 B.n331 B.n330 585
R207 B.n329 B.n58 585
R208 B.n328 B.n327 585
R209 B.n326 B.n59 585
R210 B.n325 B.n324 585
R211 B.n323 B.n60 585
R212 B.n322 B.n321 585
R213 B.n320 B.n61 585
R214 B.n319 B.n318 585
R215 B.n317 B.n62 585
R216 B.n316 B.n315 585
R217 B.n314 B.n63 585
R218 B.n313 B.n312 585
R219 B.n311 B.n64 585
R220 B.n310 B.n309 585
R221 B.n308 B.n65 585
R222 B.n307 B.n306 585
R223 B.n305 B.n66 585
R224 B.n304 B.n303 585
R225 B.n302 B.n67 585
R226 B.n301 B.n300 585
R227 B.n299 B.n68 585
R228 B.n298 B.n297 585
R229 B.n296 B.n69 585
R230 B.n295 B.n294 585
R231 B.n293 B.n70 585
R232 B.n292 B.n291 585
R233 B.n290 B.n71 585
R234 B.n289 B.n288 585
R235 B.n287 B.n72 585
R236 B.n286 B.n285 585
R237 B.n284 B.n73 585
R238 B.n283 B.n282 585
R239 B.n281 B.n74 585
R240 B.n280 B.n279 585
R241 B.n278 B.n75 585
R242 B.n277 B.n276 585
R243 B.n275 B.n76 585
R244 B.n274 B.n273 585
R245 B.n272 B.n77 585
R246 B.n271 B.n270 585
R247 B.n269 B.n78 585
R248 B.n268 B.n267 585
R249 B.n266 B.n79 585
R250 B.n265 B.n264 585
R251 B.n263 B.n80 585
R252 B.n262 B.n261 585
R253 B.n260 B.n81 585
R254 B.n259 B.n258 585
R255 B.n257 B.n82 585
R256 B.n256 B.n255 585
R257 B.n254 B.n83 585
R258 B.n253 B.n252 585
R259 B.n182 B.n111 585
R260 B.n184 B.n183 585
R261 B.n185 B.n110 585
R262 B.n187 B.n186 585
R263 B.n188 B.n109 585
R264 B.n190 B.n189 585
R265 B.n191 B.n108 585
R266 B.n193 B.n192 585
R267 B.n194 B.n107 585
R268 B.n196 B.n195 585
R269 B.n197 B.n106 585
R270 B.n199 B.n198 585
R271 B.n200 B.n105 585
R272 B.n202 B.n201 585
R273 B.n203 B.n104 585
R274 B.n205 B.n204 585
R275 B.n206 B.n103 585
R276 B.n208 B.n207 585
R277 B.n210 B.n209 585
R278 B.n211 B.n99 585
R279 B.n213 B.n212 585
R280 B.n214 B.n98 585
R281 B.n216 B.n215 585
R282 B.n217 B.n97 585
R283 B.n219 B.n218 585
R284 B.n220 B.n96 585
R285 B.n222 B.n221 585
R286 B.n223 B.n93 585
R287 B.n226 B.n225 585
R288 B.n227 B.n92 585
R289 B.n229 B.n228 585
R290 B.n230 B.n91 585
R291 B.n232 B.n231 585
R292 B.n233 B.n90 585
R293 B.n235 B.n234 585
R294 B.n236 B.n89 585
R295 B.n238 B.n237 585
R296 B.n239 B.n88 585
R297 B.n241 B.n240 585
R298 B.n242 B.n87 585
R299 B.n244 B.n243 585
R300 B.n245 B.n86 585
R301 B.n247 B.n246 585
R302 B.n248 B.n85 585
R303 B.n250 B.n249 585
R304 B.n251 B.n84 585
R305 B.n181 B.n180 585
R306 B.n179 B.n112 585
R307 B.n178 B.n177 585
R308 B.n176 B.n113 585
R309 B.n175 B.n174 585
R310 B.n173 B.n114 585
R311 B.n172 B.n171 585
R312 B.n170 B.n115 585
R313 B.n169 B.n168 585
R314 B.n167 B.n116 585
R315 B.n166 B.n165 585
R316 B.n164 B.n117 585
R317 B.n163 B.n162 585
R318 B.n161 B.n118 585
R319 B.n160 B.n159 585
R320 B.n158 B.n119 585
R321 B.n157 B.n156 585
R322 B.n155 B.n120 585
R323 B.n154 B.n153 585
R324 B.n152 B.n121 585
R325 B.n151 B.n150 585
R326 B.n149 B.n122 585
R327 B.n148 B.n147 585
R328 B.n146 B.n123 585
R329 B.n145 B.n144 585
R330 B.n143 B.n124 585
R331 B.n142 B.n141 585
R332 B.n140 B.n125 585
R333 B.n139 B.n138 585
R334 B.n137 B.n126 585
R335 B.n136 B.n135 585
R336 B.n134 B.n127 585
R337 B.n133 B.n132 585
R338 B.n131 B.n128 585
R339 B.n130 B.n129 585
R340 B.n2 B.n0 585
R341 B.n485 B.n1 585
R342 B.n484 B.n483 585
R343 B.n482 B.n3 585
R344 B.n481 B.n480 585
R345 B.n479 B.n4 585
R346 B.n478 B.n477 585
R347 B.n476 B.n5 585
R348 B.n475 B.n474 585
R349 B.n473 B.n6 585
R350 B.n472 B.n471 585
R351 B.n470 B.n7 585
R352 B.n469 B.n468 585
R353 B.n467 B.n8 585
R354 B.n466 B.n465 585
R355 B.n464 B.n9 585
R356 B.n463 B.n462 585
R357 B.n461 B.n10 585
R358 B.n460 B.n459 585
R359 B.n458 B.n11 585
R360 B.n457 B.n456 585
R361 B.n455 B.n12 585
R362 B.n454 B.n453 585
R363 B.n452 B.n13 585
R364 B.n451 B.n450 585
R365 B.n449 B.n14 585
R366 B.n448 B.n447 585
R367 B.n446 B.n15 585
R368 B.n445 B.n444 585
R369 B.n443 B.n16 585
R370 B.n442 B.n441 585
R371 B.n440 B.n17 585
R372 B.n439 B.n438 585
R373 B.n437 B.n18 585
R374 B.n436 B.n435 585
R375 B.n434 B.n19 585
R376 B.n433 B.n432 585
R377 B.n487 B.n486 585
R378 B.n180 B.n111 526.135
R379 B.n432 B.n431 526.135
R380 B.n252 B.n251 526.135
R381 B.n360 B.n47 526.135
R382 B.n94 B.t9 255.446
R383 B.n100 B.t0 255.446
R384 B.n30 B.t6 255.446
R385 B.n36 B.t3 255.446
R386 B.n94 B.t11 165.404
R387 B.n36 B.t4 165.404
R388 B.n100 B.t2 165.4
R389 B.n30 B.t7 165.4
R390 B.n180 B.n179 163.367
R391 B.n179 B.n178 163.367
R392 B.n178 B.n113 163.367
R393 B.n174 B.n113 163.367
R394 B.n174 B.n173 163.367
R395 B.n173 B.n172 163.367
R396 B.n172 B.n115 163.367
R397 B.n168 B.n115 163.367
R398 B.n168 B.n167 163.367
R399 B.n167 B.n166 163.367
R400 B.n166 B.n117 163.367
R401 B.n162 B.n117 163.367
R402 B.n162 B.n161 163.367
R403 B.n161 B.n160 163.367
R404 B.n160 B.n119 163.367
R405 B.n156 B.n119 163.367
R406 B.n156 B.n155 163.367
R407 B.n155 B.n154 163.367
R408 B.n154 B.n121 163.367
R409 B.n150 B.n121 163.367
R410 B.n150 B.n149 163.367
R411 B.n149 B.n148 163.367
R412 B.n148 B.n123 163.367
R413 B.n144 B.n123 163.367
R414 B.n144 B.n143 163.367
R415 B.n143 B.n142 163.367
R416 B.n142 B.n125 163.367
R417 B.n138 B.n125 163.367
R418 B.n138 B.n137 163.367
R419 B.n137 B.n136 163.367
R420 B.n136 B.n127 163.367
R421 B.n132 B.n127 163.367
R422 B.n132 B.n131 163.367
R423 B.n131 B.n130 163.367
R424 B.n130 B.n2 163.367
R425 B.n486 B.n2 163.367
R426 B.n486 B.n485 163.367
R427 B.n485 B.n484 163.367
R428 B.n484 B.n3 163.367
R429 B.n480 B.n3 163.367
R430 B.n480 B.n479 163.367
R431 B.n479 B.n478 163.367
R432 B.n478 B.n5 163.367
R433 B.n474 B.n5 163.367
R434 B.n474 B.n473 163.367
R435 B.n473 B.n472 163.367
R436 B.n472 B.n7 163.367
R437 B.n468 B.n7 163.367
R438 B.n468 B.n467 163.367
R439 B.n467 B.n466 163.367
R440 B.n466 B.n9 163.367
R441 B.n462 B.n9 163.367
R442 B.n462 B.n461 163.367
R443 B.n461 B.n460 163.367
R444 B.n460 B.n11 163.367
R445 B.n456 B.n11 163.367
R446 B.n456 B.n455 163.367
R447 B.n455 B.n454 163.367
R448 B.n454 B.n13 163.367
R449 B.n450 B.n13 163.367
R450 B.n450 B.n449 163.367
R451 B.n449 B.n448 163.367
R452 B.n448 B.n15 163.367
R453 B.n444 B.n15 163.367
R454 B.n444 B.n443 163.367
R455 B.n443 B.n442 163.367
R456 B.n442 B.n17 163.367
R457 B.n438 B.n17 163.367
R458 B.n438 B.n437 163.367
R459 B.n437 B.n436 163.367
R460 B.n436 B.n19 163.367
R461 B.n432 B.n19 163.367
R462 B.n184 B.n111 163.367
R463 B.n185 B.n184 163.367
R464 B.n186 B.n185 163.367
R465 B.n186 B.n109 163.367
R466 B.n190 B.n109 163.367
R467 B.n191 B.n190 163.367
R468 B.n192 B.n191 163.367
R469 B.n192 B.n107 163.367
R470 B.n196 B.n107 163.367
R471 B.n197 B.n196 163.367
R472 B.n198 B.n197 163.367
R473 B.n198 B.n105 163.367
R474 B.n202 B.n105 163.367
R475 B.n203 B.n202 163.367
R476 B.n204 B.n203 163.367
R477 B.n204 B.n103 163.367
R478 B.n208 B.n103 163.367
R479 B.n209 B.n208 163.367
R480 B.n209 B.n99 163.367
R481 B.n213 B.n99 163.367
R482 B.n214 B.n213 163.367
R483 B.n215 B.n214 163.367
R484 B.n215 B.n97 163.367
R485 B.n219 B.n97 163.367
R486 B.n220 B.n219 163.367
R487 B.n221 B.n220 163.367
R488 B.n221 B.n93 163.367
R489 B.n226 B.n93 163.367
R490 B.n227 B.n226 163.367
R491 B.n228 B.n227 163.367
R492 B.n228 B.n91 163.367
R493 B.n232 B.n91 163.367
R494 B.n233 B.n232 163.367
R495 B.n234 B.n233 163.367
R496 B.n234 B.n89 163.367
R497 B.n238 B.n89 163.367
R498 B.n239 B.n238 163.367
R499 B.n240 B.n239 163.367
R500 B.n240 B.n87 163.367
R501 B.n244 B.n87 163.367
R502 B.n245 B.n244 163.367
R503 B.n246 B.n245 163.367
R504 B.n246 B.n85 163.367
R505 B.n250 B.n85 163.367
R506 B.n251 B.n250 163.367
R507 B.n252 B.n83 163.367
R508 B.n256 B.n83 163.367
R509 B.n257 B.n256 163.367
R510 B.n258 B.n257 163.367
R511 B.n258 B.n81 163.367
R512 B.n262 B.n81 163.367
R513 B.n263 B.n262 163.367
R514 B.n264 B.n263 163.367
R515 B.n264 B.n79 163.367
R516 B.n268 B.n79 163.367
R517 B.n269 B.n268 163.367
R518 B.n270 B.n269 163.367
R519 B.n270 B.n77 163.367
R520 B.n274 B.n77 163.367
R521 B.n275 B.n274 163.367
R522 B.n276 B.n275 163.367
R523 B.n276 B.n75 163.367
R524 B.n280 B.n75 163.367
R525 B.n281 B.n280 163.367
R526 B.n282 B.n281 163.367
R527 B.n282 B.n73 163.367
R528 B.n286 B.n73 163.367
R529 B.n287 B.n286 163.367
R530 B.n288 B.n287 163.367
R531 B.n288 B.n71 163.367
R532 B.n292 B.n71 163.367
R533 B.n293 B.n292 163.367
R534 B.n294 B.n293 163.367
R535 B.n294 B.n69 163.367
R536 B.n298 B.n69 163.367
R537 B.n299 B.n298 163.367
R538 B.n300 B.n299 163.367
R539 B.n300 B.n67 163.367
R540 B.n304 B.n67 163.367
R541 B.n305 B.n304 163.367
R542 B.n306 B.n305 163.367
R543 B.n306 B.n65 163.367
R544 B.n310 B.n65 163.367
R545 B.n311 B.n310 163.367
R546 B.n312 B.n311 163.367
R547 B.n312 B.n63 163.367
R548 B.n316 B.n63 163.367
R549 B.n317 B.n316 163.367
R550 B.n318 B.n317 163.367
R551 B.n318 B.n61 163.367
R552 B.n322 B.n61 163.367
R553 B.n323 B.n322 163.367
R554 B.n324 B.n323 163.367
R555 B.n324 B.n59 163.367
R556 B.n328 B.n59 163.367
R557 B.n329 B.n328 163.367
R558 B.n330 B.n329 163.367
R559 B.n330 B.n57 163.367
R560 B.n334 B.n57 163.367
R561 B.n335 B.n334 163.367
R562 B.n336 B.n335 163.367
R563 B.n336 B.n55 163.367
R564 B.n340 B.n55 163.367
R565 B.n341 B.n340 163.367
R566 B.n342 B.n341 163.367
R567 B.n342 B.n53 163.367
R568 B.n346 B.n53 163.367
R569 B.n347 B.n346 163.367
R570 B.n348 B.n347 163.367
R571 B.n348 B.n51 163.367
R572 B.n352 B.n51 163.367
R573 B.n353 B.n352 163.367
R574 B.n354 B.n353 163.367
R575 B.n354 B.n49 163.367
R576 B.n358 B.n49 163.367
R577 B.n359 B.n358 163.367
R578 B.n360 B.n359 163.367
R579 B.n431 B.n430 163.367
R580 B.n430 B.n21 163.367
R581 B.n426 B.n21 163.367
R582 B.n426 B.n425 163.367
R583 B.n425 B.n424 163.367
R584 B.n424 B.n23 163.367
R585 B.n420 B.n23 163.367
R586 B.n420 B.n419 163.367
R587 B.n419 B.n418 163.367
R588 B.n418 B.n25 163.367
R589 B.n414 B.n25 163.367
R590 B.n414 B.n413 163.367
R591 B.n413 B.n412 163.367
R592 B.n412 B.n27 163.367
R593 B.n408 B.n27 163.367
R594 B.n408 B.n407 163.367
R595 B.n407 B.n406 163.367
R596 B.n406 B.n29 163.367
R597 B.n401 B.n29 163.367
R598 B.n401 B.n400 163.367
R599 B.n400 B.n399 163.367
R600 B.n399 B.n33 163.367
R601 B.n395 B.n33 163.367
R602 B.n395 B.n394 163.367
R603 B.n394 B.n393 163.367
R604 B.n393 B.n35 163.367
R605 B.n389 B.n35 163.367
R606 B.n389 B.n388 163.367
R607 B.n388 B.n39 163.367
R608 B.n384 B.n39 163.367
R609 B.n384 B.n383 163.367
R610 B.n383 B.n382 163.367
R611 B.n382 B.n41 163.367
R612 B.n378 B.n41 163.367
R613 B.n378 B.n377 163.367
R614 B.n377 B.n376 163.367
R615 B.n376 B.n43 163.367
R616 B.n372 B.n43 163.367
R617 B.n372 B.n371 163.367
R618 B.n371 B.n370 163.367
R619 B.n370 B.n45 163.367
R620 B.n366 B.n45 163.367
R621 B.n366 B.n365 163.367
R622 B.n365 B.n364 163.367
R623 B.n364 B.n47 163.367
R624 B.n95 B.t10 119.441
R625 B.n37 B.t5 119.441
R626 B.n101 B.t1 119.436
R627 B.n31 B.t8 119.436
R628 B.n224 B.n95 59.5399
R629 B.n102 B.n101 59.5399
R630 B.n404 B.n31 59.5399
R631 B.n38 B.n37 59.5399
R632 B.n95 B.n94 45.9641
R633 B.n101 B.n100 45.9641
R634 B.n31 B.n30 45.9641
R635 B.n37 B.n36 45.9641
R636 B.n433 B.n20 34.1859
R637 B.n362 B.n361 34.1859
R638 B.n253 B.n84 34.1859
R639 B.n182 B.n181 34.1859
R640 B B.n487 18.0485
R641 B.n429 B.n20 10.6151
R642 B.n429 B.n428 10.6151
R643 B.n428 B.n427 10.6151
R644 B.n427 B.n22 10.6151
R645 B.n423 B.n22 10.6151
R646 B.n423 B.n422 10.6151
R647 B.n422 B.n421 10.6151
R648 B.n421 B.n24 10.6151
R649 B.n417 B.n24 10.6151
R650 B.n417 B.n416 10.6151
R651 B.n416 B.n415 10.6151
R652 B.n415 B.n26 10.6151
R653 B.n411 B.n26 10.6151
R654 B.n411 B.n410 10.6151
R655 B.n410 B.n409 10.6151
R656 B.n409 B.n28 10.6151
R657 B.n405 B.n28 10.6151
R658 B.n403 B.n402 10.6151
R659 B.n402 B.n32 10.6151
R660 B.n398 B.n32 10.6151
R661 B.n398 B.n397 10.6151
R662 B.n397 B.n396 10.6151
R663 B.n396 B.n34 10.6151
R664 B.n392 B.n34 10.6151
R665 B.n392 B.n391 10.6151
R666 B.n391 B.n390 10.6151
R667 B.n387 B.n386 10.6151
R668 B.n386 B.n385 10.6151
R669 B.n385 B.n40 10.6151
R670 B.n381 B.n40 10.6151
R671 B.n381 B.n380 10.6151
R672 B.n380 B.n379 10.6151
R673 B.n379 B.n42 10.6151
R674 B.n375 B.n42 10.6151
R675 B.n375 B.n374 10.6151
R676 B.n374 B.n373 10.6151
R677 B.n373 B.n44 10.6151
R678 B.n369 B.n44 10.6151
R679 B.n369 B.n368 10.6151
R680 B.n368 B.n367 10.6151
R681 B.n367 B.n46 10.6151
R682 B.n363 B.n46 10.6151
R683 B.n363 B.n362 10.6151
R684 B.n254 B.n253 10.6151
R685 B.n255 B.n254 10.6151
R686 B.n255 B.n82 10.6151
R687 B.n259 B.n82 10.6151
R688 B.n260 B.n259 10.6151
R689 B.n261 B.n260 10.6151
R690 B.n261 B.n80 10.6151
R691 B.n265 B.n80 10.6151
R692 B.n266 B.n265 10.6151
R693 B.n267 B.n266 10.6151
R694 B.n267 B.n78 10.6151
R695 B.n271 B.n78 10.6151
R696 B.n272 B.n271 10.6151
R697 B.n273 B.n272 10.6151
R698 B.n273 B.n76 10.6151
R699 B.n277 B.n76 10.6151
R700 B.n278 B.n277 10.6151
R701 B.n279 B.n278 10.6151
R702 B.n279 B.n74 10.6151
R703 B.n283 B.n74 10.6151
R704 B.n284 B.n283 10.6151
R705 B.n285 B.n284 10.6151
R706 B.n285 B.n72 10.6151
R707 B.n289 B.n72 10.6151
R708 B.n290 B.n289 10.6151
R709 B.n291 B.n290 10.6151
R710 B.n291 B.n70 10.6151
R711 B.n295 B.n70 10.6151
R712 B.n296 B.n295 10.6151
R713 B.n297 B.n296 10.6151
R714 B.n297 B.n68 10.6151
R715 B.n301 B.n68 10.6151
R716 B.n302 B.n301 10.6151
R717 B.n303 B.n302 10.6151
R718 B.n303 B.n66 10.6151
R719 B.n307 B.n66 10.6151
R720 B.n308 B.n307 10.6151
R721 B.n309 B.n308 10.6151
R722 B.n309 B.n64 10.6151
R723 B.n313 B.n64 10.6151
R724 B.n314 B.n313 10.6151
R725 B.n315 B.n314 10.6151
R726 B.n315 B.n62 10.6151
R727 B.n319 B.n62 10.6151
R728 B.n320 B.n319 10.6151
R729 B.n321 B.n320 10.6151
R730 B.n321 B.n60 10.6151
R731 B.n325 B.n60 10.6151
R732 B.n326 B.n325 10.6151
R733 B.n327 B.n326 10.6151
R734 B.n327 B.n58 10.6151
R735 B.n331 B.n58 10.6151
R736 B.n332 B.n331 10.6151
R737 B.n333 B.n332 10.6151
R738 B.n333 B.n56 10.6151
R739 B.n337 B.n56 10.6151
R740 B.n338 B.n337 10.6151
R741 B.n339 B.n338 10.6151
R742 B.n339 B.n54 10.6151
R743 B.n343 B.n54 10.6151
R744 B.n344 B.n343 10.6151
R745 B.n345 B.n344 10.6151
R746 B.n345 B.n52 10.6151
R747 B.n349 B.n52 10.6151
R748 B.n350 B.n349 10.6151
R749 B.n351 B.n350 10.6151
R750 B.n351 B.n50 10.6151
R751 B.n355 B.n50 10.6151
R752 B.n356 B.n355 10.6151
R753 B.n357 B.n356 10.6151
R754 B.n357 B.n48 10.6151
R755 B.n361 B.n48 10.6151
R756 B.n183 B.n182 10.6151
R757 B.n183 B.n110 10.6151
R758 B.n187 B.n110 10.6151
R759 B.n188 B.n187 10.6151
R760 B.n189 B.n188 10.6151
R761 B.n189 B.n108 10.6151
R762 B.n193 B.n108 10.6151
R763 B.n194 B.n193 10.6151
R764 B.n195 B.n194 10.6151
R765 B.n195 B.n106 10.6151
R766 B.n199 B.n106 10.6151
R767 B.n200 B.n199 10.6151
R768 B.n201 B.n200 10.6151
R769 B.n201 B.n104 10.6151
R770 B.n205 B.n104 10.6151
R771 B.n206 B.n205 10.6151
R772 B.n207 B.n206 10.6151
R773 B.n211 B.n210 10.6151
R774 B.n212 B.n211 10.6151
R775 B.n212 B.n98 10.6151
R776 B.n216 B.n98 10.6151
R777 B.n217 B.n216 10.6151
R778 B.n218 B.n217 10.6151
R779 B.n218 B.n96 10.6151
R780 B.n222 B.n96 10.6151
R781 B.n223 B.n222 10.6151
R782 B.n225 B.n92 10.6151
R783 B.n229 B.n92 10.6151
R784 B.n230 B.n229 10.6151
R785 B.n231 B.n230 10.6151
R786 B.n231 B.n90 10.6151
R787 B.n235 B.n90 10.6151
R788 B.n236 B.n235 10.6151
R789 B.n237 B.n236 10.6151
R790 B.n237 B.n88 10.6151
R791 B.n241 B.n88 10.6151
R792 B.n242 B.n241 10.6151
R793 B.n243 B.n242 10.6151
R794 B.n243 B.n86 10.6151
R795 B.n247 B.n86 10.6151
R796 B.n248 B.n247 10.6151
R797 B.n249 B.n248 10.6151
R798 B.n249 B.n84 10.6151
R799 B.n181 B.n112 10.6151
R800 B.n177 B.n112 10.6151
R801 B.n177 B.n176 10.6151
R802 B.n176 B.n175 10.6151
R803 B.n175 B.n114 10.6151
R804 B.n171 B.n114 10.6151
R805 B.n171 B.n170 10.6151
R806 B.n170 B.n169 10.6151
R807 B.n169 B.n116 10.6151
R808 B.n165 B.n116 10.6151
R809 B.n165 B.n164 10.6151
R810 B.n164 B.n163 10.6151
R811 B.n163 B.n118 10.6151
R812 B.n159 B.n118 10.6151
R813 B.n159 B.n158 10.6151
R814 B.n158 B.n157 10.6151
R815 B.n157 B.n120 10.6151
R816 B.n153 B.n120 10.6151
R817 B.n153 B.n152 10.6151
R818 B.n152 B.n151 10.6151
R819 B.n151 B.n122 10.6151
R820 B.n147 B.n122 10.6151
R821 B.n147 B.n146 10.6151
R822 B.n146 B.n145 10.6151
R823 B.n145 B.n124 10.6151
R824 B.n141 B.n124 10.6151
R825 B.n141 B.n140 10.6151
R826 B.n140 B.n139 10.6151
R827 B.n139 B.n126 10.6151
R828 B.n135 B.n126 10.6151
R829 B.n135 B.n134 10.6151
R830 B.n134 B.n133 10.6151
R831 B.n133 B.n128 10.6151
R832 B.n129 B.n128 10.6151
R833 B.n129 B.n0 10.6151
R834 B.n483 B.n1 10.6151
R835 B.n483 B.n482 10.6151
R836 B.n482 B.n481 10.6151
R837 B.n481 B.n4 10.6151
R838 B.n477 B.n4 10.6151
R839 B.n477 B.n476 10.6151
R840 B.n476 B.n475 10.6151
R841 B.n475 B.n6 10.6151
R842 B.n471 B.n6 10.6151
R843 B.n471 B.n470 10.6151
R844 B.n470 B.n469 10.6151
R845 B.n469 B.n8 10.6151
R846 B.n465 B.n8 10.6151
R847 B.n465 B.n464 10.6151
R848 B.n464 B.n463 10.6151
R849 B.n463 B.n10 10.6151
R850 B.n459 B.n10 10.6151
R851 B.n459 B.n458 10.6151
R852 B.n458 B.n457 10.6151
R853 B.n457 B.n12 10.6151
R854 B.n453 B.n12 10.6151
R855 B.n453 B.n452 10.6151
R856 B.n452 B.n451 10.6151
R857 B.n451 B.n14 10.6151
R858 B.n447 B.n14 10.6151
R859 B.n447 B.n446 10.6151
R860 B.n446 B.n445 10.6151
R861 B.n445 B.n16 10.6151
R862 B.n441 B.n16 10.6151
R863 B.n441 B.n440 10.6151
R864 B.n440 B.n439 10.6151
R865 B.n439 B.n18 10.6151
R866 B.n435 B.n18 10.6151
R867 B.n435 B.n434 10.6151
R868 B.n434 B.n433 10.6151
R869 B.n405 B.n404 9.36635
R870 B.n387 B.n38 9.36635
R871 B.n207 B.n102 9.36635
R872 B.n225 B.n224 9.36635
R873 B.n487 B.n0 2.81026
R874 B.n487 B.n1 2.81026
R875 B.n404 B.n403 1.24928
R876 B.n390 B.n38 1.24928
R877 B.n210 B.n102 1.24928
R878 B.n224 B.n223 1.24928
C0 VTAIL B 1.72988f
C1 w_n2866_n1788# VN 5.14418f
C2 VTAIL VP 2.94926f
C3 w_n2866_n1788# B 6.69856f
C4 w_n2866_n1788# VP 5.51239f
C5 VDD2 VTAIL 4.61451f
C6 VDD2 w_n2866_n1788# 1.66675f
C7 VN B 0.971674f
C8 VP VN 4.92298f
C9 VP B 1.58471f
C10 VDD2 VN 2.42765f
C11 VDD2 B 1.38983f
C12 VDD2 VP 0.415231f
C13 VTAIL VDD1 4.56585f
C14 VDD1 w_n2866_n1788# 1.59989f
C15 VTAIL w_n2866_n1788# 1.79251f
C16 VDD1 VN 0.154603f
C17 VDD1 B 1.32905f
C18 VDD1 VP 2.686f
C19 VDD2 VDD1 1.1971f
C20 VTAIL VN 2.93508f
C21 VDD2 VSUBS 1.217214f
C22 VDD1 VSUBS 1.637051f
C23 VTAIL VSUBS 0.522749f
C24 VN VSUBS 5.0021f
C25 VP VSUBS 2.036148f
C26 B VSUBS 3.226239f
C27 w_n2866_n1788# VSUBS 64.485f
C28 B.n0 VSUBS 0.004431f
C29 B.n1 VSUBS 0.004431f
C30 B.n2 VSUBS 0.007007f
C31 B.n3 VSUBS 0.007007f
C32 B.n4 VSUBS 0.007007f
C33 B.n5 VSUBS 0.007007f
C34 B.n6 VSUBS 0.007007f
C35 B.n7 VSUBS 0.007007f
C36 B.n8 VSUBS 0.007007f
C37 B.n9 VSUBS 0.007007f
C38 B.n10 VSUBS 0.007007f
C39 B.n11 VSUBS 0.007007f
C40 B.n12 VSUBS 0.007007f
C41 B.n13 VSUBS 0.007007f
C42 B.n14 VSUBS 0.007007f
C43 B.n15 VSUBS 0.007007f
C44 B.n16 VSUBS 0.007007f
C45 B.n17 VSUBS 0.007007f
C46 B.n18 VSUBS 0.007007f
C47 B.n19 VSUBS 0.007007f
C48 B.n20 VSUBS 0.01716f
C49 B.n21 VSUBS 0.007007f
C50 B.n22 VSUBS 0.007007f
C51 B.n23 VSUBS 0.007007f
C52 B.n24 VSUBS 0.007007f
C53 B.n25 VSUBS 0.007007f
C54 B.n26 VSUBS 0.007007f
C55 B.n27 VSUBS 0.007007f
C56 B.n28 VSUBS 0.007007f
C57 B.n29 VSUBS 0.007007f
C58 B.t8 VSUBS 0.108793f
C59 B.t7 VSUBS 0.124439f
C60 B.t6 VSUBS 0.398519f
C61 B.n30 VSUBS 0.087684f
C62 B.n31 VSUBS 0.066296f
C63 B.n32 VSUBS 0.007007f
C64 B.n33 VSUBS 0.007007f
C65 B.n34 VSUBS 0.007007f
C66 B.n35 VSUBS 0.007007f
C67 B.t5 VSUBS 0.108793f
C68 B.t4 VSUBS 0.124438f
C69 B.t3 VSUBS 0.398519f
C70 B.n36 VSUBS 0.087684f
C71 B.n37 VSUBS 0.066296f
C72 B.n38 VSUBS 0.016234f
C73 B.n39 VSUBS 0.007007f
C74 B.n40 VSUBS 0.007007f
C75 B.n41 VSUBS 0.007007f
C76 B.n42 VSUBS 0.007007f
C77 B.n43 VSUBS 0.007007f
C78 B.n44 VSUBS 0.007007f
C79 B.n45 VSUBS 0.007007f
C80 B.n46 VSUBS 0.007007f
C81 B.n47 VSUBS 0.01716f
C82 B.n48 VSUBS 0.007007f
C83 B.n49 VSUBS 0.007007f
C84 B.n50 VSUBS 0.007007f
C85 B.n51 VSUBS 0.007007f
C86 B.n52 VSUBS 0.007007f
C87 B.n53 VSUBS 0.007007f
C88 B.n54 VSUBS 0.007007f
C89 B.n55 VSUBS 0.007007f
C90 B.n56 VSUBS 0.007007f
C91 B.n57 VSUBS 0.007007f
C92 B.n58 VSUBS 0.007007f
C93 B.n59 VSUBS 0.007007f
C94 B.n60 VSUBS 0.007007f
C95 B.n61 VSUBS 0.007007f
C96 B.n62 VSUBS 0.007007f
C97 B.n63 VSUBS 0.007007f
C98 B.n64 VSUBS 0.007007f
C99 B.n65 VSUBS 0.007007f
C100 B.n66 VSUBS 0.007007f
C101 B.n67 VSUBS 0.007007f
C102 B.n68 VSUBS 0.007007f
C103 B.n69 VSUBS 0.007007f
C104 B.n70 VSUBS 0.007007f
C105 B.n71 VSUBS 0.007007f
C106 B.n72 VSUBS 0.007007f
C107 B.n73 VSUBS 0.007007f
C108 B.n74 VSUBS 0.007007f
C109 B.n75 VSUBS 0.007007f
C110 B.n76 VSUBS 0.007007f
C111 B.n77 VSUBS 0.007007f
C112 B.n78 VSUBS 0.007007f
C113 B.n79 VSUBS 0.007007f
C114 B.n80 VSUBS 0.007007f
C115 B.n81 VSUBS 0.007007f
C116 B.n82 VSUBS 0.007007f
C117 B.n83 VSUBS 0.007007f
C118 B.n84 VSUBS 0.01716f
C119 B.n85 VSUBS 0.007007f
C120 B.n86 VSUBS 0.007007f
C121 B.n87 VSUBS 0.007007f
C122 B.n88 VSUBS 0.007007f
C123 B.n89 VSUBS 0.007007f
C124 B.n90 VSUBS 0.007007f
C125 B.n91 VSUBS 0.007007f
C126 B.n92 VSUBS 0.007007f
C127 B.n93 VSUBS 0.007007f
C128 B.t10 VSUBS 0.108793f
C129 B.t11 VSUBS 0.124438f
C130 B.t9 VSUBS 0.398519f
C131 B.n94 VSUBS 0.087684f
C132 B.n95 VSUBS 0.066296f
C133 B.n96 VSUBS 0.007007f
C134 B.n97 VSUBS 0.007007f
C135 B.n98 VSUBS 0.007007f
C136 B.n99 VSUBS 0.007007f
C137 B.t1 VSUBS 0.108793f
C138 B.t2 VSUBS 0.124439f
C139 B.t0 VSUBS 0.398519f
C140 B.n100 VSUBS 0.087684f
C141 B.n101 VSUBS 0.066296f
C142 B.n102 VSUBS 0.016234f
C143 B.n103 VSUBS 0.007007f
C144 B.n104 VSUBS 0.007007f
C145 B.n105 VSUBS 0.007007f
C146 B.n106 VSUBS 0.007007f
C147 B.n107 VSUBS 0.007007f
C148 B.n108 VSUBS 0.007007f
C149 B.n109 VSUBS 0.007007f
C150 B.n110 VSUBS 0.007007f
C151 B.n111 VSUBS 0.01716f
C152 B.n112 VSUBS 0.007007f
C153 B.n113 VSUBS 0.007007f
C154 B.n114 VSUBS 0.007007f
C155 B.n115 VSUBS 0.007007f
C156 B.n116 VSUBS 0.007007f
C157 B.n117 VSUBS 0.007007f
C158 B.n118 VSUBS 0.007007f
C159 B.n119 VSUBS 0.007007f
C160 B.n120 VSUBS 0.007007f
C161 B.n121 VSUBS 0.007007f
C162 B.n122 VSUBS 0.007007f
C163 B.n123 VSUBS 0.007007f
C164 B.n124 VSUBS 0.007007f
C165 B.n125 VSUBS 0.007007f
C166 B.n126 VSUBS 0.007007f
C167 B.n127 VSUBS 0.007007f
C168 B.n128 VSUBS 0.007007f
C169 B.n129 VSUBS 0.007007f
C170 B.n130 VSUBS 0.007007f
C171 B.n131 VSUBS 0.007007f
C172 B.n132 VSUBS 0.007007f
C173 B.n133 VSUBS 0.007007f
C174 B.n134 VSUBS 0.007007f
C175 B.n135 VSUBS 0.007007f
C176 B.n136 VSUBS 0.007007f
C177 B.n137 VSUBS 0.007007f
C178 B.n138 VSUBS 0.007007f
C179 B.n139 VSUBS 0.007007f
C180 B.n140 VSUBS 0.007007f
C181 B.n141 VSUBS 0.007007f
C182 B.n142 VSUBS 0.007007f
C183 B.n143 VSUBS 0.007007f
C184 B.n144 VSUBS 0.007007f
C185 B.n145 VSUBS 0.007007f
C186 B.n146 VSUBS 0.007007f
C187 B.n147 VSUBS 0.007007f
C188 B.n148 VSUBS 0.007007f
C189 B.n149 VSUBS 0.007007f
C190 B.n150 VSUBS 0.007007f
C191 B.n151 VSUBS 0.007007f
C192 B.n152 VSUBS 0.007007f
C193 B.n153 VSUBS 0.007007f
C194 B.n154 VSUBS 0.007007f
C195 B.n155 VSUBS 0.007007f
C196 B.n156 VSUBS 0.007007f
C197 B.n157 VSUBS 0.007007f
C198 B.n158 VSUBS 0.007007f
C199 B.n159 VSUBS 0.007007f
C200 B.n160 VSUBS 0.007007f
C201 B.n161 VSUBS 0.007007f
C202 B.n162 VSUBS 0.007007f
C203 B.n163 VSUBS 0.007007f
C204 B.n164 VSUBS 0.007007f
C205 B.n165 VSUBS 0.007007f
C206 B.n166 VSUBS 0.007007f
C207 B.n167 VSUBS 0.007007f
C208 B.n168 VSUBS 0.007007f
C209 B.n169 VSUBS 0.007007f
C210 B.n170 VSUBS 0.007007f
C211 B.n171 VSUBS 0.007007f
C212 B.n172 VSUBS 0.007007f
C213 B.n173 VSUBS 0.007007f
C214 B.n174 VSUBS 0.007007f
C215 B.n175 VSUBS 0.007007f
C216 B.n176 VSUBS 0.007007f
C217 B.n177 VSUBS 0.007007f
C218 B.n178 VSUBS 0.007007f
C219 B.n179 VSUBS 0.007007f
C220 B.n180 VSUBS 0.016639f
C221 B.n181 VSUBS 0.016639f
C222 B.n182 VSUBS 0.01716f
C223 B.n183 VSUBS 0.007007f
C224 B.n184 VSUBS 0.007007f
C225 B.n185 VSUBS 0.007007f
C226 B.n186 VSUBS 0.007007f
C227 B.n187 VSUBS 0.007007f
C228 B.n188 VSUBS 0.007007f
C229 B.n189 VSUBS 0.007007f
C230 B.n190 VSUBS 0.007007f
C231 B.n191 VSUBS 0.007007f
C232 B.n192 VSUBS 0.007007f
C233 B.n193 VSUBS 0.007007f
C234 B.n194 VSUBS 0.007007f
C235 B.n195 VSUBS 0.007007f
C236 B.n196 VSUBS 0.007007f
C237 B.n197 VSUBS 0.007007f
C238 B.n198 VSUBS 0.007007f
C239 B.n199 VSUBS 0.007007f
C240 B.n200 VSUBS 0.007007f
C241 B.n201 VSUBS 0.007007f
C242 B.n202 VSUBS 0.007007f
C243 B.n203 VSUBS 0.007007f
C244 B.n204 VSUBS 0.007007f
C245 B.n205 VSUBS 0.007007f
C246 B.n206 VSUBS 0.007007f
C247 B.n207 VSUBS 0.006595f
C248 B.n208 VSUBS 0.007007f
C249 B.n209 VSUBS 0.007007f
C250 B.n210 VSUBS 0.003916f
C251 B.n211 VSUBS 0.007007f
C252 B.n212 VSUBS 0.007007f
C253 B.n213 VSUBS 0.007007f
C254 B.n214 VSUBS 0.007007f
C255 B.n215 VSUBS 0.007007f
C256 B.n216 VSUBS 0.007007f
C257 B.n217 VSUBS 0.007007f
C258 B.n218 VSUBS 0.007007f
C259 B.n219 VSUBS 0.007007f
C260 B.n220 VSUBS 0.007007f
C261 B.n221 VSUBS 0.007007f
C262 B.n222 VSUBS 0.007007f
C263 B.n223 VSUBS 0.003916f
C264 B.n224 VSUBS 0.016234f
C265 B.n225 VSUBS 0.006595f
C266 B.n226 VSUBS 0.007007f
C267 B.n227 VSUBS 0.007007f
C268 B.n228 VSUBS 0.007007f
C269 B.n229 VSUBS 0.007007f
C270 B.n230 VSUBS 0.007007f
C271 B.n231 VSUBS 0.007007f
C272 B.n232 VSUBS 0.007007f
C273 B.n233 VSUBS 0.007007f
C274 B.n234 VSUBS 0.007007f
C275 B.n235 VSUBS 0.007007f
C276 B.n236 VSUBS 0.007007f
C277 B.n237 VSUBS 0.007007f
C278 B.n238 VSUBS 0.007007f
C279 B.n239 VSUBS 0.007007f
C280 B.n240 VSUBS 0.007007f
C281 B.n241 VSUBS 0.007007f
C282 B.n242 VSUBS 0.007007f
C283 B.n243 VSUBS 0.007007f
C284 B.n244 VSUBS 0.007007f
C285 B.n245 VSUBS 0.007007f
C286 B.n246 VSUBS 0.007007f
C287 B.n247 VSUBS 0.007007f
C288 B.n248 VSUBS 0.007007f
C289 B.n249 VSUBS 0.007007f
C290 B.n250 VSUBS 0.007007f
C291 B.n251 VSUBS 0.01716f
C292 B.n252 VSUBS 0.016639f
C293 B.n253 VSUBS 0.016639f
C294 B.n254 VSUBS 0.007007f
C295 B.n255 VSUBS 0.007007f
C296 B.n256 VSUBS 0.007007f
C297 B.n257 VSUBS 0.007007f
C298 B.n258 VSUBS 0.007007f
C299 B.n259 VSUBS 0.007007f
C300 B.n260 VSUBS 0.007007f
C301 B.n261 VSUBS 0.007007f
C302 B.n262 VSUBS 0.007007f
C303 B.n263 VSUBS 0.007007f
C304 B.n264 VSUBS 0.007007f
C305 B.n265 VSUBS 0.007007f
C306 B.n266 VSUBS 0.007007f
C307 B.n267 VSUBS 0.007007f
C308 B.n268 VSUBS 0.007007f
C309 B.n269 VSUBS 0.007007f
C310 B.n270 VSUBS 0.007007f
C311 B.n271 VSUBS 0.007007f
C312 B.n272 VSUBS 0.007007f
C313 B.n273 VSUBS 0.007007f
C314 B.n274 VSUBS 0.007007f
C315 B.n275 VSUBS 0.007007f
C316 B.n276 VSUBS 0.007007f
C317 B.n277 VSUBS 0.007007f
C318 B.n278 VSUBS 0.007007f
C319 B.n279 VSUBS 0.007007f
C320 B.n280 VSUBS 0.007007f
C321 B.n281 VSUBS 0.007007f
C322 B.n282 VSUBS 0.007007f
C323 B.n283 VSUBS 0.007007f
C324 B.n284 VSUBS 0.007007f
C325 B.n285 VSUBS 0.007007f
C326 B.n286 VSUBS 0.007007f
C327 B.n287 VSUBS 0.007007f
C328 B.n288 VSUBS 0.007007f
C329 B.n289 VSUBS 0.007007f
C330 B.n290 VSUBS 0.007007f
C331 B.n291 VSUBS 0.007007f
C332 B.n292 VSUBS 0.007007f
C333 B.n293 VSUBS 0.007007f
C334 B.n294 VSUBS 0.007007f
C335 B.n295 VSUBS 0.007007f
C336 B.n296 VSUBS 0.007007f
C337 B.n297 VSUBS 0.007007f
C338 B.n298 VSUBS 0.007007f
C339 B.n299 VSUBS 0.007007f
C340 B.n300 VSUBS 0.007007f
C341 B.n301 VSUBS 0.007007f
C342 B.n302 VSUBS 0.007007f
C343 B.n303 VSUBS 0.007007f
C344 B.n304 VSUBS 0.007007f
C345 B.n305 VSUBS 0.007007f
C346 B.n306 VSUBS 0.007007f
C347 B.n307 VSUBS 0.007007f
C348 B.n308 VSUBS 0.007007f
C349 B.n309 VSUBS 0.007007f
C350 B.n310 VSUBS 0.007007f
C351 B.n311 VSUBS 0.007007f
C352 B.n312 VSUBS 0.007007f
C353 B.n313 VSUBS 0.007007f
C354 B.n314 VSUBS 0.007007f
C355 B.n315 VSUBS 0.007007f
C356 B.n316 VSUBS 0.007007f
C357 B.n317 VSUBS 0.007007f
C358 B.n318 VSUBS 0.007007f
C359 B.n319 VSUBS 0.007007f
C360 B.n320 VSUBS 0.007007f
C361 B.n321 VSUBS 0.007007f
C362 B.n322 VSUBS 0.007007f
C363 B.n323 VSUBS 0.007007f
C364 B.n324 VSUBS 0.007007f
C365 B.n325 VSUBS 0.007007f
C366 B.n326 VSUBS 0.007007f
C367 B.n327 VSUBS 0.007007f
C368 B.n328 VSUBS 0.007007f
C369 B.n329 VSUBS 0.007007f
C370 B.n330 VSUBS 0.007007f
C371 B.n331 VSUBS 0.007007f
C372 B.n332 VSUBS 0.007007f
C373 B.n333 VSUBS 0.007007f
C374 B.n334 VSUBS 0.007007f
C375 B.n335 VSUBS 0.007007f
C376 B.n336 VSUBS 0.007007f
C377 B.n337 VSUBS 0.007007f
C378 B.n338 VSUBS 0.007007f
C379 B.n339 VSUBS 0.007007f
C380 B.n340 VSUBS 0.007007f
C381 B.n341 VSUBS 0.007007f
C382 B.n342 VSUBS 0.007007f
C383 B.n343 VSUBS 0.007007f
C384 B.n344 VSUBS 0.007007f
C385 B.n345 VSUBS 0.007007f
C386 B.n346 VSUBS 0.007007f
C387 B.n347 VSUBS 0.007007f
C388 B.n348 VSUBS 0.007007f
C389 B.n349 VSUBS 0.007007f
C390 B.n350 VSUBS 0.007007f
C391 B.n351 VSUBS 0.007007f
C392 B.n352 VSUBS 0.007007f
C393 B.n353 VSUBS 0.007007f
C394 B.n354 VSUBS 0.007007f
C395 B.n355 VSUBS 0.007007f
C396 B.n356 VSUBS 0.007007f
C397 B.n357 VSUBS 0.007007f
C398 B.n358 VSUBS 0.007007f
C399 B.n359 VSUBS 0.007007f
C400 B.n360 VSUBS 0.016639f
C401 B.n361 VSUBS 0.01743f
C402 B.n362 VSUBS 0.016369f
C403 B.n363 VSUBS 0.007007f
C404 B.n364 VSUBS 0.007007f
C405 B.n365 VSUBS 0.007007f
C406 B.n366 VSUBS 0.007007f
C407 B.n367 VSUBS 0.007007f
C408 B.n368 VSUBS 0.007007f
C409 B.n369 VSUBS 0.007007f
C410 B.n370 VSUBS 0.007007f
C411 B.n371 VSUBS 0.007007f
C412 B.n372 VSUBS 0.007007f
C413 B.n373 VSUBS 0.007007f
C414 B.n374 VSUBS 0.007007f
C415 B.n375 VSUBS 0.007007f
C416 B.n376 VSUBS 0.007007f
C417 B.n377 VSUBS 0.007007f
C418 B.n378 VSUBS 0.007007f
C419 B.n379 VSUBS 0.007007f
C420 B.n380 VSUBS 0.007007f
C421 B.n381 VSUBS 0.007007f
C422 B.n382 VSUBS 0.007007f
C423 B.n383 VSUBS 0.007007f
C424 B.n384 VSUBS 0.007007f
C425 B.n385 VSUBS 0.007007f
C426 B.n386 VSUBS 0.007007f
C427 B.n387 VSUBS 0.006595f
C428 B.n388 VSUBS 0.007007f
C429 B.n389 VSUBS 0.007007f
C430 B.n390 VSUBS 0.003916f
C431 B.n391 VSUBS 0.007007f
C432 B.n392 VSUBS 0.007007f
C433 B.n393 VSUBS 0.007007f
C434 B.n394 VSUBS 0.007007f
C435 B.n395 VSUBS 0.007007f
C436 B.n396 VSUBS 0.007007f
C437 B.n397 VSUBS 0.007007f
C438 B.n398 VSUBS 0.007007f
C439 B.n399 VSUBS 0.007007f
C440 B.n400 VSUBS 0.007007f
C441 B.n401 VSUBS 0.007007f
C442 B.n402 VSUBS 0.007007f
C443 B.n403 VSUBS 0.003916f
C444 B.n404 VSUBS 0.016234f
C445 B.n405 VSUBS 0.006595f
C446 B.n406 VSUBS 0.007007f
C447 B.n407 VSUBS 0.007007f
C448 B.n408 VSUBS 0.007007f
C449 B.n409 VSUBS 0.007007f
C450 B.n410 VSUBS 0.007007f
C451 B.n411 VSUBS 0.007007f
C452 B.n412 VSUBS 0.007007f
C453 B.n413 VSUBS 0.007007f
C454 B.n414 VSUBS 0.007007f
C455 B.n415 VSUBS 0.007007f
C456 B.n416 VSUBS 0.007007f
C457 B.n417 VSUBS 0.007007f
C458 B.n418 VSUBS 0.007007f
C459 B.n419 VSUBS 0.007007f
C460 B.n420 VSUBS 0.007007f
C461 B.n421 VSUBS 0.007007f
C462 B.n422 VSUBS 0.007007f
C463 B.n423 VSUBS 0.007007f
C464 B.n424 VSUBS 0.007007f
C465 B.n425 VSUBS 0.007007f
C466 B.n426 VSUBS 0.007007f
C467 B.n427 VSUBS 0.007007f
C468 B.n428 VSUBS 0.007007f
C469 B.n429 VSUBS 0.007007f
C470 B.n430 VSUBS 0.007007f
C471 B.n431 VSUBS 0.01716f
C472 B.n432 VSUBS 0.016639f
C473 B.n433 VSUBS 0.016639f
C474 B.n434 VSUBS 0.007007f
C475 B.n435 VSUBS 0.007007f
C476 B.n436 VSUBS 0.007007f
C477 B.n437 VSUBS 0.007007f
C478 B.n438 VSUBS 0.007007f
C479 B.n439 VSUBS 0.007007f
C480 B.n440 VSUBS 0.007007f
C481 B.n441 VSUBS 0.007007f
C482 B.n442 VSUBS 0.007007f
C483 B.n443 VSUBS 0.007007f
C484 B.n444 VSUBS 0.007007f
C485 B.n445 VSUBS 0.007007f
C486 B.n446 VSUBS 0.007007f
C487 B.n447 VSUBS 0.007007f
C488 B.n448 VSUBS 0.007007f
C489 B.n449 VSUBS 0.007007f
C490 B.n450 VSUBS 0.007007f
C491 B.n451 VSUBS 0.007007f
C492 B.n452 VSUBS 0.007007f
C493 B.n453 VSUBS 0.007007f
C494 B.n454 VSUBS 0.007007f
C495 B.n455 VSUBS 0.007007f
C496 B.n456 VSUBS 0.007007f
C497 B.n457 VSUBS 0.007007f
C498 B.n458 VSUBS 0.007007f
C499 B.n459 VSUBS 0.007007f
C500 B.n460 VSUBS 0.007007f
C501 B.n461 VSUBS 0.007007f
C502 B.n462 VSUBS 0.007007f
C503 B.n463 VSUBS 0.007007f
C504 B.n464 VSUBS 0.007007f
C505 B.n465 VSUBS 0.007007f
C506 B.n466 VSUBS 0.007007f
C507 B.n467 VSUBS 0.007007f
C508 B.n468 VSUBS 0.007007f
C509 B.n469 VSUBS 0.007007f
C510 B.n470 VSUBS 0.007007f
C511 B.n471 VSUBS 0.007007f
C512 B.n472 VSUBS 0.007007f
C513 B.n473 VSUBS 0.007007f
C514 B.n474 VSUBS 0.007007f
C515 B.n475 VSUBS 0.007007f
C516 B.n476 VSUBS 0.007007f
C517 B.n477 VSUBS 0.007007f
C518 B.n478 VSUBS 0.007007f
C519 B.n479 VSUBS 0.007007f
C520 B.n480 VSUBS 0.007007f
C521 B.n481 VSUBS 0.007007f
C522 B.n482 VSUBS 0.007007f
C523 B.n483 VSUBS 0.007007f
C524 B.n484 VSUBS 0.007007f
C525 B.n485 VSUBS 0.007007f
C526 B.n486 VSUBS 0.007007f
C527 B.n487 VSUBS 0.015866f
C528 VDD1.t2 VSUBS 0.601109f
C529 VDD1.t5 VSUBS 0.600534f
C530 VDD1.t0 VSUBS 0.073505f
C531 VDD1.t1 VSUBS 0.073505f
C532 VDD1.n0 VSUBS 0.434937f
C533 VDD1.n1 VSUBS 2.34017f
C534 VDD1.t3 VSUBS 0.073505f
C535 VDD1.t4 VSUBS 0.073505f
C536 VDD1.n2 VSUBS 0.432732f
C537 VDD1.n3 VSUBS 1.96523f
C538 VP.n0 VSUBS 0.064829f
C539 VP.t4 VSUBS 1.05896f
C540 VP.n1 VSUBS 0.062641f
C541 VP.n2 VSUBS 0.049176f
C542 VP.t5 VSUBS 1.05896f
C543 VP.n3 VSUBS 0.062641f
C544 VP.n4 VSUBS 0.064829f
C545 VP.t0 VSUBS 1.05896f
C546 VP.n5 VSUBS 0.064829f
C547 VP.t1 VSUBS 1.05896f
C548 VP.n6 VSUBS 0.062641f
C549 VP.t3 VSUBS 1.34074f
C550 VP.n7 VSUBS 0.527812f
C551 VP.t2 VSUBS 1.05896f
C552 VP.n8 VSUBS 0.573576f
C553 VP.n9 VSUBS 0.091192f
C554 VP.n10 VSUBS 0.411311f
C555 VP.n11 VSUBS 0.049176f
C556 VP.n12 VSUBS 0.049176f
C557 VP.n13 VSUBS 0.080328f
C558 VP.n14 VSUBS 0.079487f
C559 VP.n15 VSUBS 0.577166f
C560 VP.n16 VSUBS 1.95277f
C561 VP.n17 VSUBS 1.99654f
C562 VP.n18 VSUBS 0.577166f
C563 VP.n19 VSUBS 0.079487f
C564 VP.n20 VSUBS 0.080328f
C565 VP.n21 VSUBS 0.049176f
C566 VP.n22 VSUBS 0.049176f
C567 VP.n23 VSUBS 0.049176f
C568 VP.n24 VSUBS 0.091192f
C569 VP.n25 VSUBS 0.475415f
C570 VP.n26 VSUBS 0.091192f
C571 VP.n27 VSUBS 0.049176f
C572 VP.n28 VSUBS 0.049176f
C573 VP.n29 VSUBS 0.049176f
C574 VP.n30 VSUBS 0.080328f
C575 VP.n31 VSUBS 0.079487f
C576 VP.n32 VSUBS 0.577166f
C577 VP.n33 VSUBS 0.062365f
C578 VTAIL.t9 VSUBS 0.09193f
C579 VTAIL.t11 VSUBS 0.09193f
C580 VTAIL.n0 VSUBS 0.466819f
C581 VTAIL.n1 VSUBS 0.629911f
C582 VTAIL.t0 VSUBS 0.666768f
C583 VTAIL.n2 VSUBS 0.815455f
C584 VTAIL.t5 VSUBS 0.09193f
C585 VTAIL.t2 VSUBS 0.09193f
C586 VTAIL.n3 VSUBS 0.466819f
C587 VTAIL.n4 VSUBS 1.7105f
C588 VTAIL.t10 VSUBS 0.09193f
C589 VTAIL.t7 VSUBS 0.09193f
C590 VTAIL.n5 VSUBS 0.466822f
C591 VTAIL.n6 VSUBS 1.71049f
C592 VTAIL.t8 VSUBS 0.666771f
C593 VTAIL.n7 VSUBS 0.815452f
C594 VTAIL.t1 VSUBS 0.09193f
C595 VTAIL.t4 VSUBS 0.09193f
C596 VTAIL.n8 VSUBS 0.466822f
C597 VTAIL.n9 VSUBS 0.764684f
C598 VTAIL.t3 VSUBS 0.666768f
C599 VTAIL.n10 VSUBS 1.57447f
C600 VTAIL.t6 VSUBS 0.666768f
C601 VTAIL.n11 VSUBS 1.52245f
C602 VDD2.t5 VSUBS 0.582541f
C603 VDD2.t4 VSUBS 0.071303f
C604 VDD2.t2 VSUBS 0.071303f
C605 VDD2.n0 VSUBS 0.421906f
C606 VDD2.n1 VSUBS 2.17953f
C607 VDD2.t0 VSUBS 0.576598f
C608 VDD2.n2 VSUBS 1.88903f
C609 VDD2.t3 VSUBS 0.071303f
C610 VDD2.t1 VSUBS 0.071303f
C611 VDD2.n3 VSUBS 0.421886f
C612 VN.n0 VSUBS 0.061726f
C613 VN.t5 VSUBS 1.00827f
C614 VN.n1 VSUBS 0.059643f
C615 VN.t2 VSUBS 1.27657f
C616 VN.n2 VSUBS 0.502549f
C617 VN.t0 VSUBS 1.00827f
C618 VN.n3 VSUBS 0.546123f
C619 VN.n4 VSUBS 0.086827f
C620 VN.n5 VSUBS 0.391624f
C621 VN.n6 VSUBS 0.046822f
C622 VN.n7 VSUBS 0.046822f
C623 VN.n8 VSUBS 0.076483f
C624 VN.n9 VSUBS 0.075682f
C625 VN.n10 VSUBS 0.549541f
C626 VN.n11 VSUBS 0.05938f
C627 VN.n12 VSUBS 0.061726f
C628 VN.t1 VSUBS 1.00827f
C629 VN.n13 VSUBS 0.059643f
C630 VN.t3 VSUBS 1.27657f
C631 VN.n14 VSUBS 0.502549f
C632 VN.t4 VSUBS 1.00827f
C633 VN.n15 VSUBS 0.546123f
C634 VN.n16 VSUBS 0.086827f
C635 VN.n17 VSUBS 0.391624f
C636 VN.n18 VSUBS 0.046822f
C637 VN.n19 VSUBS 0.046822f
C638 VN.n20 VSUBS 0.076483f
C639 VN.n21 VSUBS 0.075682f
C640 VN.n22 VSUBS 0.549541f
C641 VN.n23 VSUBS 1.8854f
.ends

