* NGSPICE file created from diff_pair_sample_1654.ext - technology: sky130A

.subckt diff_pair_sample_1654 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=2.52
X1 VTAIL.t9 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=2.52
X3 VTAIL.t15 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X4 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=2.52
X5 VDD2.t6 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X6 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X7 VTAIL.t5 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=2.52
X8 VTAIL.t7 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X9 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=2.52
X10 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=2.52
X11 VDD1.t4 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X12 VDD2.t1 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=2.52
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=2.52
X14 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X15 VTAIL.t11 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=2.52
X16 VDD1.t2 VP.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=1.44705 ps=9.1 w=8.77 l=2.52
X17 VDD1.t1 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=1.44705 pd=9.1 as=3.4203 ps=18.32 w=8.77 l=2.52
X18 VTAIL.t8 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=1.44705 ps=9.1 w=8.77 l=2.52
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.4203 pd=18.32 as=0 ps=0 w=8.77 l=2.52
R0 VP.n19 VP.n18 161.3
R1 VP.n20 VP.n15 161.3
R2 VP.n22 VP.n21 161.3
R3 VP.n23 VP.n14 161.3
R4 VP.n25 VP.n24 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n28 VP.n12 161.3
R7 VP.n30 VP.n29 161.3
R8 VP.n31 VP.n11 161.3
R9 VP.n33 VP.n32 161.3
R10 VP.n34 VP.n10 161.3
R11 VP.n64 VP.n0 161.3
R12 VP.n63 VP.n62 161.3
R13 VP.n61 VP.n1 161.3
R14 VP.n60 VP.n59 161.3
R15 VP.n58 VP.n2 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n53 VP.n4 161.3
R19 VP.n52 VP.n51 161.3
R20 VP.n50 VP.n5 161.3
R21 VP.n49 VP.n48 161.3
R22 VP.n46 VP.n6 161.3
R23 VP.n45 VP.n44 161.3
R24 VP.n43 VP.n7 161.3
R25 VP.n42 VP.n41 161.3
R26 VP.n40 VP.n8 161.3
R27 VP.n39 VP.n38 161.3
R28 VP.n16 VP.t4 118.445
R29 VP.n37 VP.n9 97.2996
R30 VP.n66 VP.n65 97.2996
R31 VP.n36 VP.n35 97.2996
R32 VP.n9 VP.t7 83.8723
R33 VP.n47 VP.t5 83.8723
R34 VP.n3 VP.t1 83.8723
R35 VP.n65 VP.t6 83.8723
R36 VP.n35 VP.t0 83.8723
R37 VP.n13 VP.t2 83.8723
R38 VP.n17 VP.t3 83.8723
R39 VP.n41 VP.n7 55.0624
R40 VP.n59 VP.n1 55.0624
R41 VP.n29 VP.n11 55.0624
R42 VP.n17 VP.n16 51.8291
R43 VP.n37 VP.n36 48.1284
R44 VP.n52 VP.n5 40.4934
R45 VP.n53 VP.n52 40.4934
R46 VP.n23 VP.n22 40.4934
R47 VP.n22 VP.n15 40.4934
R48 VP.n41 VP.n40 25.9244
R49 VP.n63 VP.n1 25.9244
R50 VP.n33 VP.n11 25.9244
R51 VP.n40 VP.n39 24.4675
R52 VP.n45 VP.n7 24.4675
R53 VP.n46 VP.n45 24.4675
R54 VP.n48 VP.n5 24.4675
R55 VP.n54 VP.n53 24.4675
R56 VP.n58 VP.n57 24.4675
R57 VP.n59 VP.n58 24.4675
R58 VP.n64 VP.n63 24.4675
R59 VP.n34 VP.n33 24.4675
R60 VP.n24 VP.n23 24.4675
R61 VP.n28 VP.n27 24.4675
R62 VP.n29 VP.n28 24.4675
R63 VP.n18 VP.n15 24.4675
R64 VP.n48 VP.n47 20.7975
R65 VP.n54 VP.n3 20.7975
R66 VP.n24 VP.n13 20.7975
R67 VP.n18 VP.n17 20.7975
R68 VP.n39 VP.n9 13.4574
R69 VP.n65 VP.n64 13.4574
R70 VP.n35 VP.n34 13.4574
R71 VP.n19 VP.n16 6.62497
R72 VP.n47 VP.n46 3.67055
R73 VP.n57 VP.n3 3.67055
R74 VP.n27 VP.n13 3.67055
R75 VP.n36 VP.n10 0.278367
R76 VP.n38 VP.n37 0.278367
R77 VP.n66 VP.n0 0.278367
R78 VP.n20 VP.n19 0.189894
R79 VP.n21 VP.n20 0.189894
R80 VP.n21 VP.n14 0.189894
R81 VP.n25 VP.n14 0.189894
R82 VP.n26 VP.n25 0.189894
R83 VP.n26 VP.n12 0.189894
R84 VP.n30 VP.n12 0.189894
R85 VP.n31 VP.n30 0.189894
R86 VP.n32 VP.n31 0.189894
R87 VP.n32 VP.n10 0.189894
R88 VP.n38 VP.n8 0.189894
R89 VP.n42 VP.n8 0.189894
R90 VP.n43 VP.n42 0.189894
R91 VP.n44 VP.n43 0.189894
R92 VP.n44 VP.n6 0.189894
R93 VP.n49 VP.n6 0.189894
R94 VP.n50 VP.n49 0.189894
R95 VP.n51 VP.n50 0.189894
R96 VP.n51 VP.n4 0.189894
R97 VP.n55 VP.n4 0.189894
R98 VP.n56 VP.n55 0.189894
R99 VP.n56 VP.n2 0.189894
R100 VP.n60 VP.n2 0.189894
R101 VP.n61 VP.n60 0.189894
R102 VP.n62 VP.n61 0.189894
R103 VP.n62 VP.n0 0.189894
R104 VP VP.n66 0.153454
R105 VTAIL.n386 VTAIL.n344 289.615
R106 VTAIL.n44 VTAIL.n2 289.615
R107 VTAIL.n92 VTAIL.n50 289.615
R108 VTAIL.n142 VTAIL.n100 289.615
R109 VTAIL.n338 VTAIL.n296 289.615
R110 VTAIL.n288 VTAIL.n246 289.615
R111 VTAIL.n240 VTAIL.n198 289.615
R112 VTAIL.n190 VTAIL.n148 289.615
R113 VTAIL.n361 VTAIL.n360 185
R114 VTAIL.n363 VTAIL.n362 185
R115 VTAIL.n356 VTAIL.n355 185
R116 VTAIL.n369 VTAIL.n368 185
R117 VTAIL.n371 VTAIL.n370 185
R118 VTAIL.n352 VTAIL.n351 185
R119 VTAIL.n377 VTAIL.n376 185
R120 VTAIL.n379 VTAIL.n378 185
R121 VTAIL.n348 VTAIL.n347 185
R122 VTAIL.n385 VTAIL.n384 185
R123 VTAIL.n387 VTAIL.n386 185
R124 VTAIL.n19 VTAIL.n18 185
R125 VTAIL.n21 VTAIL.n20 185
R126 VTAIL.n14 VTAIL.n13 185
R127 VTAIL.n27 VTAIL.n26 185
R128 VTAIL.n29 VTAIL.n28 185
R129 VTAIL.n10 VTAIL.n9 185
R130 VTAIL.n35 VTAIL.n34 185
R131 VTAIL.n37 VTAIL.n36 185
R132 VTAIL.n6 VTAIL.n5 185
R133 VTAIL.n43 VTAIL.n42 185
R134 VTAIL.n45 VTAIL.n44 185
R135 VTAIL.n67 VTAIL.n66 185
R136 VTAIL.n69 VTAIL.n68 185
R137 VTAIL.n62 VTAIL.n61 185
R138 VTAIL.n75 VTAIL.n74 185
R139 VTAIL.n77 VTAIL.n76 185
R140 VTAIL.n58 VTAIL.n57 185
R141 VTAIL.n83 VTAIL.n82 185
R142 VTAIL.n85 VTAIL.n84 185
R143 VTAIL.n54 VTAIL.n53 185
R144 VTAIL.n91 VTAIL.n90 185
R145 VTAIL.n93 VTAIL.n92 185
R146 VTAIL.n117 VTAIL.n116 185
R147 VTAIL.n119 VTAIL.n118 185
R148 VTAIL.n112 VTAIL.n111 185
R149 VTAIL.n125 VTAIL.n124 185
R150 VTAIL.n127 VTAIL.n126 185
R151 VTAIL.n108 VTAIL.n107 185
R152 VTAIL.n133 VTAIL.n132 185
R153 VTAIL.n135 VTAIL.n134 185
R154 VTAIL.n104 VTAIL.n103 185
R155 VTAIL.n141 VTAIL.n140 185
R156 VTAIL.n143 VTAIL.n142 185
R157 VTAIL.n339 VTAIL.n338 185
R158 VTAIL.n337 VTAIL.n336 185
R159 VTAIL.n300 VTAIL.n299 185
R160 VTAIL.n331 VTAIL.n330 185
R161 VTAIL.n329 VTAIL.n328 185
R162 VTAIL.n304 VTAIL.n303 185
R163 VTAIL.n323 VTAIL.n322 185
R164 VTAIL.n321 VTAIL.n320 185
R165 VTAIL.n308 VTAIL.n307 185
R166 VTAIL.n315 VTAIL.n314 185
R167 VTAIL.n313 VTAIL.n312 185
R168 VTAIL.n289 VTAIL.n288 185
R169 VTAIL.n287 VTAIL.n286 185
R170 VTAIL.n250 VTAIL.n249 185
R171 VTAIL.n281 VTAIL.n280 185
R172 VTAIL.n279 VTAIL.n278 185
R173 VTAIL.n254 VTAIL.n253 185
R174 VTAIL.n273 VTAIL.n272 185
R175 VTAIL.n271 VTAIL.n270 185
R176 VTAIL.n258 VTAIL.n257 185
R177 VTAIL.n265 VTAIL.n264 185
R178 VTAIL.n263 VTAIL.n262 185
R179 VTAIL.n241 VTAIL.n240 185
R180 VTAIL.n239 VTAIL.n238 185
R181 VTAIL.n202 VTAIL.n201 185
R182 VTAIL.n233 VTAIL.n232 185
R183 VTAIL.n231 VTAIL.n230 185
R184 VTAIL.n206 VTAIL.n205 185
R185 VTAIL.n225 VTAIL.n224 185
R186 VTAIL.n223 VTAIL.n222 185
R187 VTAIL.n210 VTAIL.n209 185
R188 VTAIL.n217 VTAIL.n216 185
R189 VTAIL.n215 VTAIL.n214 185
R190 VTAIL.n191 VTAIL.n190 185
R191 VTAIL.n189 VTAIL.n188 185
R192 VTAIL.n152 VTAIL.n151 185
R193 VTAIL.n183 VTAIL.n182 185
R194 VTAIL.n181 VTAIL.n180 185
R195 VTAIL.n156 VTAIL.n155 185
R196 VTAIL.n175 VTAIL.n174 185
R197 VTAIL.n173 VTAIL.n172 185
R198 VTAIL.n160 VTAIL.n159 185
R199 VTAIL.n167 VTAIL.n166 185
R200 VTAIL.n165 VTAIL.n164 185
R201 VTAIL.n261 VTAIL.t11 147.659
R202 VTAIL.n213 VTAIL.t6 147.659
R203 VTAIL.n163 VTAIL.t3 147.659
R204 VTAIL.n359 VTAIL.t0 147.659
R205 VTAIL.n17 VTAIL.t5 147.659
R206 VTAIL.n65 VTAIL.t13 147.659
R207 VTAIL.n115 VTAIL.t8 147.659
R208 VTAIL.n311 VTAIL.t14 147.659
R209 VTAIL.n362 VTAIL.n361 104.615
R210 VTAIL.n362 VTAIL.n355 104.615
R211 VTAIL.n369 VTAIL.n355 104.615
R212 VTAIL.n370 VTAIL.n369 104.615
R213 VTAIL.n370 VTAIL.n351 104.615
R214 VTAIL.n377 VTAIL.n351 104.615
R215 VTAIL.n378 VTAIL.n377 104.615
R216 VTAIL.n378 VTAIL.n347 104.615
R217 VTAIL.n385 VTAIL.n347 104.615
R218 VTAIL.n386 VTAIL.n385 104.615
R219 VTAIL.n20 VTAIL.n19 104.615
R220 VTAIL.n20 VTAIL.n13 104.615
R221 VTAIL.n27 VTAIL.n13 104.615
R222 VTAIL.n28 VTAIL.n27 104.615
R223 VTAIL.n28 VTAIL.n9 104.615
R224 VTAIL.n35 VTAIL.n9 104.615
R225 VTAIL.n36 VTAIL.n35 104.615
R226 VTAIL.n36 VTAIL.n5 104.615
R227 VTAIL.n43 VTAIL.n5 104.615
R228 VTAIL.n44 VTAIL.n43 104.615
R229 VTAIL.n68 VTAIL.n67 104.615
R230 VTAIL.n68 VTAIL.n61 104.615
R231 VTAIL.n75 VTAIL.n61 104.615
R232 VTAIL.n76 VTAIL.n75 104.615
R233 VTAIL.n76 VTAIL.n57 104.615
R234 VTAIL.n83 VTAIL.n57 104.615
R235 VTAIL.n84 VTAIL.n83 104.615
R236 VTAIL.n84 VTAIL.n53 104.615
R237 VTAIL.n91 VTAIL.n53 104.615
R238 VTAIL.n92 VTAIL.n91 104.615
R239 VTAIL.n118 VTAIL.n117 104.615
R240 VTAIL.n118 VTAIL.n111 104.615
R241 VTAIL.n125 VTAIL.n111 104.615
R242 VTAIL.n126 VTAIL.n125 104.615
R243 VTAIL.n126 VTAIL.n107 104.615
R244 VTAIL.n133 VTAIL.n107 104.615
R245 VTAIL.n134 VTAIL.n133 104.615
R246 VTAIL.n134 VTAIL.n103 104.615
R247 VTAIL.n141 VTAIL.n103 104.615
R248 VTAIL.n142 VTAIL.n141 104.615
R249 VTAIL.n338 VTAIL.n337 104.615
R250 VTAIL.n337 VTAIL.n299 104.615
R251 VTAIL.n330 VTAIL.n299 104.615
R252 VTAIL.n330 VTAIL.n329 104.615
R253 VTAIL.n329 VTAIL.n303 104.615
R254 VTAIL.n322 VTAIL.n303 104.615
R255 VTAIL.n322 VTAIL.n321 104.615
R256 VTAIL.n321 VTAIL.n307 104.615
R257 VTAIL.n314 VTAIL.n307 104.615
R258 VTAIL.n314 VTAIL.n313 104.615
R259 VTAIL.n288 VTAIL.n287 104.615
R260 VTAIL.n287 VTAIL.n249 104.615
R261 VTAIL.n280 VTAIL.n249 104.615
R262 VTAIL.n280 VTAIL.n279 104.615
R263 VTAIL.n279 VTAIL.n253 104.615
R264 VTAIL.n272 VTAIL.n253 104.615
R265 VTAIL.n272 VTAIL.n271 104.615
R266 VTAIL.n271 VTAIL.n257 104.615
R267 VTAIL.n264 VTAIL.n257 104.615
R268 VTAIL.n264 VTAIL.n263 104.615
R269 VTAIL.n240 VTAIL.n239 104.615
R270 VTAIL.n239 VTAIL.n201 104.615
R271 VTAIL.n232 VTAIL.n201 104.615
R272 VTAIL.n232 VTAIL.n231 104.615
R273 VTAIL.n231 VTAIL.n205 104.615
R274 VTAIL.n224 VTAIL.n205 104.615
R275 VTAIL.n224 VTAIL.n223 104.615
R276 VTAIL.n223 VTAIL.n209 104.615
R277 VTAIL.n216 VTAIL.n209 104.615
R278 VTAIL.n216 VTAIL.n215 104.615
R279 VTAIL.n190 VTAIL.n189 104.615
R280 VTAIL.n189 VTAIL.n151 104.615
R281 VTAIL.n182 VTAIL.n151 104.615
R282 VTAIL.n182 VTAIL.n181 104.615
R283 VTAIL.n181 VTAIL.n155 104.615
R284 VTAIL.n174 VTAIL.n155 104.615
R285 VTAIL.n174 VTAIL.n173 104.615
R286 VTAIL.n173 VTAIL.n159 104.615
R287 VTAIL.n166 VTAIL.n159 104.615
R288 VTAIL.n166 VTAIL.n165 104.615
R289 VTAIL.n361 VTAIL.t0 52.3082
R290 VTAIL.n19 VTAIL.t5 52.3082
R291 VTAIL.n67 VTAIL.t13 52.3082
R292 VTAIL.n117 VTAIL.t8 52.3082
R293 VTAIL.n313 VTAIL.t14 52.3082
R294 VTAIL.n263 VTAIL.t11 52.3082
R295 VTAIL.n215 VTAIL.t6 52.3082
R296 VTAIL.n165 VTAIL.t3 52.3082
R297 VTAIL.n295 VTAIL.n294 45.126
R298 VTAIL.n197 VTAIL.n196 45.126
R299 VTAIL.n1 VTAIL.n0 45.1259
R300 VTAIL.n99 VTAIL.n98 45.1259
R301 VTAIL.n391 VTAIL.n390 30.052
R302 VTAIL.n49 VTAIL.n48 30.052
R303 VTAIL.n97 VTAIL.n96 30.052
R304 VTAIL.n147 VTAIL.n146 30.052
R305 VTAIL.n343 VTAIL.n342 30.052
R306 VTAIL.n293 VTAIL.n292 30.052
R307 VTAIL.n245 VTAIL.n244 30.052
R308 VTAIL.n195 VTAIL.n194 30.052
R309 VTAIL.n391 VTAIL.n343 22.3841
R310 VTAIL.n195 VTAIL.n147 22.3841
R311 VTAIL.n360 VTAIL.n359 15.6677
R312 VTAIL.n18 VTAIL.n17 15.6677
R313 VTAIL.n66 VTAIL.n65 15.6677
R314 VTAIL.n116 VTAIL.n115 15.6677
R315 VTAIL.n312 VTAIL.n311 15.6677
R316 VTAIL.n262 VTAIL.n261 15.6677
R317 VTAIL.n214 VTAIL.n213 15.6677
R318 VTAIL.n164 VTAIL.n163 15.6677
R319 VTAIL.n363 VTAIL.n358 12.8005
R320 VTAIL.n21 VTAIL.n16 12.8005
R321 VTAIL.n69 VTAIL.n64 12.8005
R322 VTAIL.n119 VTAIL.n114 12.8005
R323 VTAIL.n315 VTAIL.n310 12.8005
R324 VTAIL.n265 VTAIL.n260 12.8005
R325 VTAIL.n217 VTAIL.n212 12.8005
R326 VTAIL.n167 VTAIL.n162 12.8005
R327 VTAIL.n364 VTAIL.n356 12.0247
R328 VTAIL.n22 VTAIL.n14 12.0247
R329 VTAIL.n70 VTAIL.n62 12.0247
R330 VTAIL.n120 VTAIL.n112 12.0247
R331 VTAIL.n316 VTAIL.n308 12.0247
R332 VTAIL.n266 VTAIL.n258 12.0247
R333 VTAIL.n218 VTAIL.n210 12.0247
R334 VTAIL.n168 VTAIL.n160 12.0247
R335 VTAIL.n368 VTAIL.n367 11.249
R336 VTAIL.n26 VTAIL.n25 11.249
R337 VTAIL.n74 VTAIL.n73 11.249
R338 VTAIL.n124 VTAIL.n123 11.249
R339 VTAIL.n320 VTAIL.n319 11.249
R340 VTAIL.n270 VTAIL.n269 11.249
R341 VTAIL.n222 VTAIL.n221 11.249
R342 VTAIL.n172 VTAIL.n171 11.249
R343 VTAIL.n371 VTAIL.n354 10.4732
R344 VTAIL.n29 VTAIL.n12 10.4732
R345 VTAIL.n77 VTAIL.n60 10.4732
R346 VTAIL.n127 VTAIL.n110 10.4732
R347 VTAIL.n323 VTAIL.n306 10.4732
R348 VTAIL.n273 VTAIL.n256 10.4732
R349 VTAIL.n225 VTAIL.n208 10.4732
R350 VTAIL.n175 VTAIL.n158 10.4732
R351 VTAIL.n372 VTAIL.n352 9.69747
R352 VTAIL.n30 VTAIL.n10 9.69747
R353 VTAIL.n78 VTAIL.n58 9.69747
R354 VTAIL.n128 VTAIL.n108 9.69747
R355 VTAIL.n324 VTAIL.n304 9.69747
R356 VTAIL.n274 VTAIL.n254 9.69747
R357 VTAIL.n226 VTAIL.n206 9.69747
R358 VTAIL.n176 VTAIL.n156 9.69747
R359 VTAIL.n390 VTAIL.n389 9.45567
R360 VTAIL.n48 VTAIL.n47 9.45567
R361 VTAIL.n96 VTAIL.n95 9.45567
R362 VTAIL.n146 VTAIL.n145 9.45567
R363 VTAIL.n342 VTAIL.n341 9.45567
R364 VTAIL.n292 VTAIL.n291 9.45567
R365 VTAIL.n244 VTAIL.n243 9.45567
R366 VTAIL.n194 VTAIL.n193 9.45567
R367 VTAIL.n383 VTAIL.n382 9.3005
R368 VTAIL.n346 VTAIL.n345 9.3005
R369 VTAIL.n389 VTAIL.n388 9.3005
R370 VTAIL.n350 VTAIL.n349 9.3005
R371 VTAIL.n375 VTAIL.n374 9.3005
R372 VTAIL.n373 VTAIL.n372 9.3005
R373 VTAIL.n354 VTAIL.n353 9.3005
R374 VTAIL.n367 VTAIL.n366 9.3005
R375 VTAIL.n365 VTAIL.n364 9.3005
R376 VTAIL.n358 VTAIL.n357 9.3005
R377 VTAIL.n381 VTAIL.n380 9.3005
R378 VTAIL.n41 VTAIL.n40 9.3005
R379 VTAIL.n4 VTAIL.n3 9.3005
R380 VTAIL.n47 VTAIL.n46 9.3005
R381 VTAIL.n8 VTAIL.n7 9.3005
R382 VTAIL.n33 VTAIL.n32 9.3005
R383 VTAIL.n31 VTAIL.n30 9.3005
R384 VTAIL.n12 VTAIL.n11 9.3005
R385 VTAIL.n25 VTAIL.n24 9.3005
R386 VTAIL.n23 VTAIL.n22 9.3005
R387 VTAIL.n16 VTAIL.n15 9.3005
R388 VTAIL.n39 VTAIL.n38 9.3005
R389 VTAIL.n89 VTAIL.n88 9.3005
R390 VTAIL.n52 VTAIL.n51 9.3005
R391 VTAIL.n95 VTAIL.n94 9.3005
R392 VTAIL.n56 VTAIL.n55 9.3005
R393 VTAIL.n81 VTAIL.n80 9.3005
R394 VTAIL.n79 VTAIL.n78 9.3005
R395 VTAIL.n60 VTAIL.n59 9.3005
R396 VTAIL.n73 VTAIL.n72 9.3005
R397 VTAIL.n71 VTAIL.n70 9.3005
R398 VTAIL.n64 VTAIL.n63 9.3005
R399 VTAIL.n87 VTAIL.n86 9.3005
R400 VTAIL.n139 VTAIL.n138 9.3005
R401 VTAIL.n102 VTAIL.n101 9.3005
R402 VTAIL.n145 VTAIL.n144 9.3005
R403 VTAIL.n106 VTAIL.n105 9.3005
R404 VTAIL.n131 VTAIL.n130 9.3005
R405 VTAIL.n129 VTAIL.n128 9.3005
R406 VTAIL.n110 VTAIL.n109 9.3005
R407 VTAIL.n123 VTAIL.n122 9.3005
R408 VTAIL.n121 VTAIL.n120 9.3005
R409 VTAIL.n114 VTAIL.n113 9.3005
R410 VTAIL.n137 VTAIL.n136 9.3005
R411 VTAIL.n298 VTAIL.n297 9.3005
R412 VTAIL.n335 VTAIL.n334 9.3005
R413 VTAIL.n333 VTAIL.n332 9.3005
R414 VTAIL.n302 VTAIL.n301 9.3005
R415 VTAIL.n327 VTAIL.n326 9.3005
R416 VTAIL.n325 VTAIL.n324 9.3005
R417 VTAIL.n306 VTAIL.n305 9.3005
R418 VTAIL.n319 VTAIL.n318 9.3005
R419 VTAIL.n317 VTAIL.n316 9.3005
R420 VTAIL.n310 VTAIL.n309 9.3005
R421 VTAIL.n341 VTAIL.n340 9.3005
R422 VTAIL.n248 VTAIL.n247 9.3005
R423 VTAIL.n291 VTAIL.n290 9.3005
R424 VTAIL.n285 VTAIL.n284 9.3005
R425 VTAIL.n283 VTAIL.n282 9.3005
R426 VTAIL.n252 VTAIL.n251 9.3005
R427 VTAIL.n277 VTAIL.n276 9.3005
R428 VTAIL.n275 VTAIL.n274 9.3005
R429 VTAIL.n256 VTAIL.n255 9.3005
R430 VTAIL.n269 VTAIL.n268 9.3005
R431 VTAIL.n267 VTAIL.n266 9.3005
R432 VTAIL.n260 VTAIL.n259 9.3005
R433 VTAIL.n200 VTAIL.n199 9.3005
R434 VTAIL.n243 VTAIL.n242 9.3005
R435 VTAIL.n237 VTAIL.n236 9.3005
R436 VTAIL.n235 VTAIL.n234 9.3005
R437 VTAIL.n204 VTAIL.n203 9.3005
R438 VTAIL.n229 VTAIL.n228 9.3005
R439 VTAIL.n227 VTAIL.n226 9.3005
R440 VTAIL.n208 VTAIL.n207 9.3005
R441 VTAIL.n221 VTAIL.n220 9.3005
R442 VTAIL.n219 VTAIL.n218 9.3005
R443 VTAIL.n212 VTAIL.n211 9.3005
R444 VTAIL.n150 VTAIL.n149 9.3005
R445 VTAIL.n193 VTAIL.n192 9.3005
R446 VTAIL.n187 VTAIL.n186 9.3005
R447 VTAIL.n185 VTAIL.n184 9.3005
R448 VTAIL.n154 VTAIL.n153 9.3005
R449 VTAIL.n179 VTAIL.n178 9.3005
R450 VTAIL.n177 VTAIL.n176 9.3005
R451 VTAIL.n158 VTAIL.n157 9.3005
R452 VTAIL.n171 VTAIL.n170 9.3005
R453 VTAIL.n169 VTAIL.n168 9.3005
R454 VTAIL.n162 VTAIL.n161 9.3005
R455 VTAIL.n376 VTAIL.n375 8.92171
R456 VTAIL.n390 VTAIL.n344 8.92171
R457 VTAIL.n34 VTAIL.n33 8.92171
R458 VTAIL.n48 VTAIL.n2 8.92171
R459 VTAIL.n82 VTAIL.n81 8.92171
R460 VTAIL.n96 VTAIL.n50 8.92171
R461 VTAIL.n132 VTAIL.n131 8.92171
R462 VTAIL.n146 VTAIL.n100 8.92171
R463 VTAIL.n342 VTAIL.n296 8.92171
R464 VTAIL.n328 VTAIL.n327 8.92171
R465 VTAIL.n292 VTAIL.n246 8.92171
R466 VTAIL.n278 VTAIL.n277 8.92171
R467 VTAIL.n244 VTAIL.n198 8.92171
R468 VTAIL.n230 VTAIL.n229 8.92171
R469 VTAIL.n194 VTAIL.n148 8.92171
R470 VTAIL.n180 VTAIL.n179 8.92171
R471 VTAIL.n379 VTAIL.n350 8.14595
R472 VTAIL.n388 VTAIL.n387 8.14595
R473 VTAIL.n37 VTAIL.n8 8.14595
R474 VTAIL.n46 VTAIL.n45 8.14595
R475 VTAIL.n85 VTAIL.n56 8.14595
R476 VTAIL.n94 VTAIL.n93 8.14595
R477 VTAIL.n135 VTAIL.n106 8.14595
R478 VTAIL.n144 VTAIL.n143 8.14595
R479 VTAIL.n340 VTAIL.n339 8.14595
R480 VTAIL.n331 VTAIL.n302 8.14595
R481 VTAIL.n290 VTAIL.n289 8.14595
R482 VTAIL.n281 VTAIL.n252 8.14595
R483 VTAIL.n242 VTAIL.n241 8.14595
R484 VTAIL.n233 VTAIL.n204 8.14595
R485 VTAIL.n192 VTAIL.n191 8.14595
R486 VTAIL.n183 VTAIL.n154 8.14595
R487 VTAIL.n380 VTAIL.n348 7.3702
R488 VTAIL.n384 VTAIL.n346 7.3702
R489 VTAIL.n38 VTAIL.n6 7.3702
R490 VTAIL.n42 VTAIL.n4 7.3702
R491 VTAIL.n86 VTAIL.n54 7.3702
R492 VTAIL.n90 VTAIL.n52 7.3702
R493 VTAIL.n136 VTAIL.n104 7.3702
R494 VTAIL.n140 VTAIL.n102 7.3702
R495 VTAIL.n336 VTAIL.n298 7.3702
R496 VTAIL.n332 VTAIL.n300 7.3702
R497 VTAIL.n286 VTAIL.n248 7.3702
R498 VTAIL.n282 VTAIL.n250 7.3702
R499 VTAIL.n238 VTAIL.n200 7.3702
R500 VTAIL.n234 VTAIL.n202 7.3702
R501 VTAIL.n188 VTAIL.n150 7.3702
R502 VTAIL.n184 VTAIL.n152 7.3702
R503 VTAIL.n383 VTAIL.n348 6.59444
R504 VTAIL.n384 VTAIL.n383 6.59444
R505 VTAIL.n41 VTAIL.n6 6.59444
R506 VTAIL.n42 VTAIL.n41 6.59444
R507 VTAIL.n89 VTAIL.n54 6.59444
R508 VTAIL.n90 VTAIL.n89 6.59444
R509 VTAIL.n139 VTAIL.n104 6.59444
R510 VTAIL.n140 VTAIL.n139 6.59444
R511 VTAIL.n336 VTAIL.n335 6.59444
R512 VTAIL.n335 VTAIL.n300 6.59444
R513 VTAIL.n286 VTAIL.n285 6.59444
R514 VTAIL.n285 VTAIL.n250 6.59444
R515 VTAIL.n238 VTAIL.n237 6.59444
R516 VTAIL.n237 VTAIL.n202 6.59444
R517 VTAIL.n188 VTAIL.n187 6.59444
R518 VTAIL.n187 VTAIL.n152 6.59444
R519 VTAIL.n380 VTAIL.n379 5.81868
R520 VTAIL.n387 VTAIL.n346 5.81868
R521 VTAIL.n38 VTAIL.n37 5.81868
R522 VTAIL.n45 VTAIL.n4 5.81868
R523 VTAIL.n86 VTAIL.n85 5.81868
R524 VTAIL.n93 VTAIL.n52 5.81868
R525 VTAIL.n136 VTAIL.n135 5.81868
R526 VTAIL.n143 VTAIL.n102 5.81868
R527 VTAIL.n339 VTAIL.n298 5.81868
R528 VTAIL.n332 VTAIL.n331 5.81868
R529 VTAIL.n289 VTAIL.n248 5.81868
R530 VTAIL.n282 VTAIL.n281 5.81868
R531 VTAIL.n241 VTAIL.n200 5.81868
R532 VTAIL.n234 VTAIL.n233 5.81868
R533 VTAIL.n191 VTAIL.n150 5.81868
R534 VTAIL.n184 VTAIL.n183 5.81868
R535 VTAIL.n376 VTAIL.n350 5.04292
R536 VTAIL.n388 VTAIL.n344 5.04292
R537 VTAIL.n34 VTAIL.n8 5.04292
R538 VTAIL.n46 VTAIL.n2 5.04292
R539 VTAIL.n82 VTAIL.n56 5.04292
R540 VTAIL.n94 VTAIL.n50 5.04292
R541 VTAIL.n132 VTAIL.n106 5.04292
R542 VTAIL.n144 VTAIL.n100 5.04292
R543 VTAIL.n340 VTAIL.n296 5.04292
R544 VTAIL.n328 VTAIL.n302 5.04292
R545 VTAIL.n290 VTAIL.n246 5.04292
R546 VTAIL.n278 VTAIL.n252 5.04292
R547 VTAIL.n242 VTAIL.n198 5.04292
R548 VTAIL.n230 VTAIL.n204 5.04292
R549 VTAIL.n192 VTAIL.n148 5.04292
R550 VTAIL.n180 VTAIL.n154 5.04292
R551 VTAIL.n359 VTAIL.n357 4.38563
R552 VTAIL.n17 VTAIL.n15 4.38563
R553 VTAIL.n65 VTAIL.n63 4.38563
R554 VTAIL.n115 VTAIL.n113 4.38563
R555 VTAIL.n311 VTAIL.n309 4.38563
R556 VTAIL.n261 VTAIL.n259 4.38563
R557 VTAIL.n213 VTAIL.n211 4.38563
R558 VTAIL.n163 VTAIL.n161 4.38563
R559 VTAIL.n375 VTAIL.n352 4.26717
R560 VTAIL.n33 VTAIL.n10 4.26717
R561 VTAIL.n81 VTAIL.n58 4.26717
R562 VTAIL.n131 VTAIL.n108 4.26717
R563 VTAIL.n327 VTAIL.n304 4.26717
R564 VTAIL.n277 VTAIL.n254 4.26717
R565 VTAIL.n229 VTAIL.n206 4.26717
R566 VTAIL.n179 VTAIL.n156 4.26717
R567 VTAIL.n372 VTAIL.n371 3.49141
R568 VTAIL.n30 VTAIL.n29 3.49141
R569 VTAIL.n78 VTAIL.n77 3.49141
R570 VTAIL.n128 VTAIL.n127 3.49141
R571 VTAIL.n324 VTAIL.n323 3.49141
R572 VTAIL.n274 VTAIL.n273 3.49141
R573 VTAIL.n226 VTAIL.n225 3.49141
R574 VTAIL.n176 VTAIL.n175 3.49141
R575 VTAIL.n368 VTAIL.n354 2.71565
R576 VTAIL.n26 VTAIL.n12 2.71565
R577 VTAIL.n74 VTAIL.n60 2.71565
R578 VTAIL.n124 VTAIL.n110 2.71565
R579 VTAIL.n320 VTAIL.n306 2.71565
R580 VTAIL.n270 VTAIL.n256 2.71565
R581 VTAIL.n222 VTAIL.n208 2.71565
R582 VTAIL.n172 VTAIL.n158 2.71565
R583 VTAIL.n197 VTAIL.n195 2.4574
R584 VTAIL.n245 VTAIL.n197 2.4574
R585 VTAIL.n295 VTAIL.n293 2.4574
R586 VTAIL.n343 VTAIL.n295 2.4574
R587 VTAIL.n147 VTAIL.n99 2.4574
R588 VTAIL.n99 VTAIL.n97 2.4574
R589 VTAIL.n49 VTAIL.n1 2.4574
R590 VTAIL VTAIL.n391 2.39921
R591 VTAIL.n0 VTAIL.t4 2.2582
R592 VTAIL.n0 VTAIL.t2 2.2582
R593 VTAIL.n98 VTAIL.t10 2.2582
R594 VTAIL.n98 VTAIL.t9 2.2582
R595 VTAIL.n294 VTAIL.t12 2.2582
R596 VTAIL.n294 VTAIL.t15 2.2582
R597 VTAIL.n196 VTAIL.t1 2.2582
R598 VTAIL.n196 VTAIL.t7 2.2582
R599 VTAIL.n367 VTAIL.n356 1.93989
R600 VTAIL.n25 VTAIL.n14 1.93989
R601 VTAIL.n73 VTAIL.n62 1.93989
R602 VTAIL.n123 VTAIL.n112 1.93989
R603 VTAIL.n319 VTAIL.n308 1.93989
R604 VTAIL.n269 VTAIL.n258 1.93989
R605 VTAIL.n221 VTAIL.n210 1.93989
R606 VTAIL.n171 VTAIL.n160 1.93989
R607 VTAIL.n364 VTAIL.n363 1.16414
R608 VTAIL.n22 VTAIL.n21 1.16414
R609 VTAIL.n70 VTAIL.n69 1.16414
R610 VTAIL.n120 VTAIL.n119 1.16414
R611 VTAIL.n316 VTAIL.n315 1.16414
R612 VTAIL.n266 VTAIL.n265 1.16414
R613 VTAIL.n218 VTAIL.n217 1.16414
R614 VTAIL.n168 VTAIL.n167 1.16414
R615 VTAIL.n293 VTAIL.n245 0.470328
R616 VTAIL.n97 VTAIL.n49 0.470328
R617 VTAIL.n360 VTAIL.n358 0.388379
R618 VTAIL.n18 VTAIL.n16 0.388379
R619 VTAIL.n66 VTAIL.n64 0.388379
R620 VTAIL.n116 VTAIL.n114 0.388379
R621 VTAIL.n312 VTAIL.n310 0.388379
R622 VTAIL.n262 VTAIL.n260 0.388379
R623 VTAIL.n214 VTAIL.n212 0.388379
R624 VTAIL.n164 VTAIL.n162 0.388379
R625 VTAIL.n365 VTAIL.n357 0.155672
R626 VTAIL.n366 VTAIL.n365 0.155672
R627 VTAIL.n366 VTAIL.n353 0.155672
R628 VTAIL.n373 VTAIL.n353 0.155672
R629 VTAIL.n374 VTAIL.n373 0.155672
R630 VTAIL.n374 VTAIL.n349 0.155672
R631 VTAIL.n381 VTAIL.n349 0.155672
R632 VTAIL.n382 VTAIL.n381 0.155672
R633 VTAIL.n382 VTAIL.n345 0.155672
R634 VTAIL.n389 VTAIL.n345 0.155672
R635 VTAIL.n23 VTAIL.n15 0.155672
R636 VTAIL.n24 VTAIL.n23 0.155672
R637 VTAIL.n24 VTAIL.n11 0.155672
R638 VTAIL.n31 VTAIL.n11 0.155672
R639 VTAIL.n32 VTAIL.n31 0.155672
R640 VTAIL.n32 VTAIL.n7 0.155672
R641 VTAIL.n39 VTAIL.n7 0.155672
R642 VTAIL.n40 VTAIL.n39 0.155672
R643 VTAIL.n40 VTAIL.n3 0.155672
R644 VTAIL.n47 VTAIL.n3 0.155672
R645 VTAIL.n71 VTAIL.n63 0.155672
R646 VTAIL.n72 VTAIL.n71 0.155672
R647 VTAIL.n72 VTAIL.n59 0.155672
R648 VTAIL.n79 VTAIL.n59 0.155672
R649 VTAIL.n80 VTAIL.n79 0.155672
R650 VTAIL.n80 VTAIL.n55 0.155672
R651 VTAIL.n87 VTAIL.n55 0.155672
R652 VTAIL.n88 VTAIL.n87 0.155672
R653 VTAIL.n88 VTAIL.n51 0.155672
R654 VTAIL.n95 VTAIL.n51 0.155672
R655 VTAIL.n121 VTAIL.n113 0.155672
R656 VTAIL.n122 VTAIL.n121 0.155672
R657 VTAIL.n122 VTAIL.n109 0.155672
R658 VTAIL.n129 VTAIL.n109 0.155672
R659 VTAIL.n130 VTAIL.n129 0.155672
R660 VTAIL.n130 VTAIL.n105 0.155672
R661 VTAIL.n137 VTAIL.n105 0.155672
R662 VTAIL.n138 VTAIL.n137 0.155672
R663 VTAIL.n138 VTAIL.n101 0.155672
R664 VTAIL.n145 VTAIL.n101 0.155672
R665 VTAIL.n341 VTAIL.n297 0.155672
R666 VTAIL.n334 VTAIL.n297 0.155672
R667 VTAIL.n334 VTAIL.n333 0.155672
R668 VTAIL.n333 VTAIL.n301 0.155672
R669 VTAIL.n326 VTAIL.n301 0.155672
R670 VTAIL.n326 VTAIL.n325 0.155672
R671 VTAIL.n325 VTAIL.n305 0.155672
R672 VTAIL.n318 VTAIL.n305 0.155672
R673 VTAIL.n318 VTAIL.n317 0.155672
R674 VTAIL.n317 VTAIL.n309 0.155672
R675 VTAIL.n291 VTAIL.n247 0.155672
R676 VTAIL.n284 VTAIL.n247 0.155672
R677 VTAIL.n284 VTAIL.n283 0.155672
R678 VTAIL.n283 VTAIL.n251 0.155672
R679 VTAIL.n276 VTAIL.n251 0.155672
R680 VTAIL.n276 VTAIL.n275 0.155672
R681 VTAIL.n275 VTAIL.n255 0.155672
R682 VTAIL.n268 VTAIL.n255 0.155672
R683 VTAIL.n268 VTAIL.n267 0.155672
R684 VTAIL.n267 VTAIL.n259 0.155672
R685 VTAIL.n243 VTAIL.n199 0.155672
R686 VTAIL.n236 VTAIL.n199 0.155672
R687 VTAIL.n236 VTAIL.n235 0.155672
R688 VTAIL.n235 VTAIL.n203 0.155672
R689 VTAIL.n228 VTAIL.n203 0.155672
R690 VTAIL.n228 VTAIL.n227 0.155672
R691 VTAIL.n227 VTAIL.n207 0.155672
R692 VTAIL.n220 VTAIL.n207 0.155672
R693 VTAIL.n220 VTAIL.n219 0.155672
R694 VTAIL.n219 VTAIL.n211 0.155672
R695 VTAIL.n193 VTAIL.n149 0.155672
R696 VTAIL.n186 VTAIL.n149 0.155672
R697 VTAIL.n186 VTAIL.n185 0.155672
R698 VTAIL.n185 VTAIL.n153 0.155672
R699 VTAIL.n178 VTAIL.n153 0.155672
R700 VTAIL.n178 VTAIL.n177 0.155672
R701 VTAIL.n177 VTAIL.n157 0.155672
R702 VTAIL.n170 VTAIL.n157 0.155672
R703 VTAIL.n170 VTAIL.n169 0.155672
R704 VTAIL.n169 VTAIL.n161 0.155672
R705 VTAIL VTAIL.n1 0.0586897
R706 VDD1 VDD1.n0 63.0914
R707 VDD1.n3 VDD1.n2 62.9777
R708 VDD1.n3 VDD1.n1 62.9777
R709 VDD1.n5 VDD1.n4 61.8048
R710 VDD1.n5 VDD1.n3 42.9147
R711 VDD1.n4 VDD1.t5 2.2582
R712 VDD1.n4 VDD1.t7 2.2582
R713 VDD1.n0 VDD1.t3 2.2582
R714 VDD1.n0 VDD1.t4 2.2582
R715 VDD1.n2 VDD1.t6 2.2582
R716 VDD1.n2 VDD1.t1 2.2582
R717 VDD1.n1 VDD1.t0 2.2582
R718 VDD1.n1 VDD1.t2 2.2582
R719 VDD1 VDD1.n5 1.17076
R720 B.n637 B.n636 585
R721 B.n639 B.n134 585
R722 B.n642 B.n641 585
R723 B.n643 B.n133 585
R724 B.n645 B.n644 585
R725 B.n647 B.n132 585
R726 B.n650 B.n649 585
R727 B.n651 B.n131 585
R728 B.n653 B.n652 585
R729 B.n655 B.n130 585
R730 B.n658 B.n657 585
R731 B.n659 B.n129 585
R732 B.n661 B.n660 585
R733 B.n663 B.n128 585
R734 B.n666 B.n665 585
R735 B.n667 B.n127 585
R736 B.n669 B.n668 585
R737 B.n671 B.n126 585
R738 B.n674 B.n673 585
R739 B.n675 B.n125 585
R740 B.n677 B.n676 585
R741 B.n679 B.n124 585
R742 B.n682 B.n681 585
R743 B.n683 B.n123 585
R744 B.n685 B.n684 585
R745 B.n687 B.n122 585
R746 B.n690 B.n689 585
R747 B.n691 B.n121 585
R748 B.n693 B.n692 585
R749 B.n695 B.n120 585
R750 B.n697 B.n696 585
R751 B.n699 B.n698 585
R752 B.n702 B.n701 585
R753 B.n703 B.n115 585
R754 B.n705 B.n704 585
R755 B.n707 B.n114 585
R756 B.n710 B.n709 585
R757 B.n711 B.n113 585
R758 B.n713 B.n712 585
R759 B.n715 B.n112 585
R760 B.n718 B.n717 585
R761 B.n719 B.n109 585
R762 B.n722 B.n721 585
R763 B.n724 B.n108 585
R764 B.n727 B.n726 585
R765 B.n728 B.n107 585
R766 B.n730 B.n729 585
R767 B.n732 B.n106 585
R768 B.n735 B.n734 585
R769 B.n736 B.n105 585
R770 B.n738 B.n737 585
R771 B.n740 B.n104 585
R772 B.n743 B.n742 585
R773 B.n744 B.n103 585
R774 B.n746 B.n745 585
R775 B.n748 B.n102 585
R776 B.n751 B.n750 585
R777 B.n752 B.n101 585
R778 B.n754 B.n753 585
R779 B.n756 B.n100 585
R780 B.n759 B.n758 585
R781 B.n760 B.n99 585
R782 B.n762 B.n761 585
R783 B.n764 B.n98 585
R784 B.n767 B.n766 585
R785 B.n768 B.n97 585
R786 B.n770 B.n769 585
R787 B.n772 B.n96 585
R788 B.n775 B.n774 585
R789 B.n776 B.n95 585
R790 B.n778 B.n777 585
R791 B.n780 B.n94 585
R792 B.n783 B.n782 585
R793 B.n784 B.n93 585
R794 B.n635 B.n91 585
R795 B.n787 B.n91 585
R796 B.n634 B.n90 585
R797 B.n788 B.n90 585
R798 B.n633 B.n89 585
R799 B.n789 B.n89 585
R800 B.n632 B.n631 585
R801 B.n631 B.n85 585
R802 B.n630 B.n84 585
R803 B.n795 B.n84 585
R804 B.n629 B.n83 585
R805 B.n796 B.n83 585
R806 B.n628 B.n82 585
R807 B.n797 B.n82 585
R808 B.n627 B.n626 585
R809 B.n626 B.n81 585
R810 B.n625 B.n77 585
R811 B.n803 B.n77 585
R812 B.n624 B.n76 585
R813 B.n804 B.n76 585
R814 B.n623 B.n75 585
R815 B.n805 B.n75 585
R816 B.n622 B.n621 585
R817 B.n621 B.n71 585
R818 B.n620 B.n70 585
R819 B.n811 B.n70 585
R820 B.n619 B.n69 585
R821 B.n812 B.n69 585
R822 B.n618 B.n68 585
R823 B.n813 B.n68 585
R824 B.n617 B.n616 585
R825 B.n616 B.n64 585
R826 B.n615 B.n63 585
R827 B.n819 B.n63 585
R828 B.n614 B.n62 585
R829 B.n820 B.n62 585
R830 B.n613 B.n61 585
R831 B.n821 B.n61 585
R832 B.n612 B.n611 585
R833 B.n611 B.n60 585
R834 B.n610 B.n56 585
R835 B.n827 B.n56 585
R836 B.n609 B.n55 585
R837 B.n828 B.n55 585
R838 B.n608 B.n54 585
R839 B.n829 B.n54 585
R840 B.n607 B.n606 585
R841 B.n606 B.n50 585
R842 B.n605 B.n49 585
R843 B.n835 B.n49 585
R844 B.n604 B.n48 585
R845 B.n836 B.n48 585
R846 B.n603 B.n47 585
R847 B.n837 B.n47 585
R848 B.n602 B.n601 585
R849 B.n601 B.n46 585
R850 B.n600 B.n42 585
R851 B.n843 B.n42 585
R852 B.n599 B.n41 585
R853 B.n844 B.n41 585
R854 B.n598 B.n40 585
R855 B.n845 B.n40 585
R856 B.n597 B.n596 585
R857 B.n596 B.n36 585
R858 B.n595 B.n35 585
R859 B.n851 B.n35 585
R860 B.n594 B.n34 585
R861 B.n852 B.n34 585
R862 B.n593 B.n33 585
R863 B.n853 B.n33 585
R864 B.n592 B.n591 585
R865 B.n591 B.n32 585
R866 B.n590 B.n28 585
R867 B.n859 B.n28 585
R868 B.n589 B.n27 585
R869 B.n860 B.n27 585
R870 B.n588 B.n26 585
R871 B.n861 B.n26 585
R872 B.n587 B.n586 585
R873 B.n586 B.n22 585
R874 B.n585 B.n21 585
R875 B.n867 B.n21 585
R876 B.n584 B.n20 585
R877 B.n868 B.n20 585
R878 B.n583 B.n19 585
R879 B.n869 B.n19 585
R880 B.n582 B.n581 585
R881 B.n581 B.n15 585
R882 B.n580 B.n14 585
R883 B.n875 B.n14 585
R884 B.n579 B.n13 585
R885 B.n876 B.n13 585
R886 B.n578 B.n12 585
R887 B.n877 B.n12 585
R888 B.n577 B.n576 585
R889 B.n576 B.n8 585
R890 B.n575 B.n7 585
R891 B.n883 B.n7 585
R892 B.n574 B.n6 585
R893 B.n884 B.n6 585
R894 B.n573 B.n5 585
R895 B.n885 B.n5 585
R896 B.n572 B.n571 585
R897 B.n571 B.n4 585
R898 B.n570 B.n135 585
R899 B.n570 B.n569 585
R900 B.n560 B.n136 585
R901 B.n137 B.n136 585
R902 B.n562 B.n561 585
R903 B.n563 B.n562 585
R904 B.n559 B.n142 585
R905 B.n142 B.n141 585
R906 B.n558 B.n557 585
R907 B.n557 B.n556 585
R908 B.n144 B.n143 585
R909 B.n145 B.n144 585
R910 B.n549 B.n548 585
R911 B.n550 B.n549 585
R912 B.n547 B.n150 585
R913 B.n150 B.n149 585
R914 B.n546 B.n545 585
R915 B.n545 B.n544 585
R916 B.n152 B.n151 585
R917 B.n153 B.n152 585
R918 B.n537 B.n536 585
R919 B.n538 B.n537 585
R920 B.n535 B.n158 585
R921 B.n158 B.n157 585
R922 B.n534 B.n533 585
R923 B.n533 B.n532 585
R924 B.n160 B.n159 585
R925 B.n525 B.n160 585
R926 B.n524 B.n523 585
R927 B.n526 B.n524 585
R928 B.n522 B.n165 585
R929 B.n165 B.n164 585
R930 B.n521 B.n520 585
R931 B.n520 B.n519 585
R932 B.n167 B.n166 585
R933 B.n168 B.n167 585
R934 B.n512 B.n511 585
R935 B.n513 B.n512 585
R936 B.n510 B.n173 585
R937 B.n173 B.n172 585
R938 B.n509 B.n508 585
R939 B.n508 B.n507 585
R940 B.n175 B.n174 585
R941 B.n500 B.n175 585
R942 B.n499 B.n498 585
R943 B.n501 B.n499 585
R944 B.n497 B.n180 585
R945 B.n180 B.n179 585
R946 B.n496 B.n495 585
R947 B.n495 B.n494 585
R948 B.n182 B.n181 585
R949 B.n183 B.n182 585
R950 B.n487 B.n486 585
R951 B.n488 B.n487 585
R952 B.n485 B.n188 585
R953 B.n188 B.n187 585
R954 B.n484 B.n483 585
R955 B.n483 B.n482 585
R956 B.n190 B.n189 585
R957 B.n475 B.n190 585
R958 B.n474 B.n473 585
R959 B.n476 B.n474 585
R960 B.n472 B.n195 585
R961 B.n195 B.n194 585
R962 B.n471 B.n470 585
R963 B.n470 B.n469 585
R964 B.n197 B.n196 585
R965 B.n198 B.n197 585
R966 B.n462 B.n461 585
R967 B.n463 B.n462 585
R968 B.n460 B.n203 585
R969 B.n203 B.n202 585
R970 B.n459 B.n458 585
R971 B.n458 B.n457 585
R972 B.n205 B.n204 585
R973 B.n206 B.n205 585
R974 B.n450 B.n449 585
R975 B.n451 B.n450 585
R976 B.n448 B.n211 585
R977 B.n211 B.n210 585
R978 B.n447 B.n446 585
R979 B.n446 B.n445 585
R980 B.n213 B.n212 585
R981 B.n438 B.n213 585
R982 B.n437 B.n436 585
R983 B.n439 B.n437 585
R984 B.n435 B.n218 585
R985 B.n218 B.n217 585
R986 B.n434 B.n433 585
R987 B.n433 B.n432 585
R988 B.n220 B.n219 585
R989 B.n221 B.n220 585
R990 B.n425 B.n424 585
R991 B.n426 B.n425 585
R992 B.n423 B.n226 585
R993 B.n226 B.n225 585
R994 B.n422 B.n421 585
R995 B.n421 B.n420 585
R996 B.n417 B.n230 585
R997 B.n416 B.n415 585
R998 B.n413 B.n231 585
R999 B.n413 B.n229 585
R1000 B.n412 B.n411 585
R1001 B.n410 B.n409 585
R1002 B.n408 B.n233 585
R1003 B.n406 B.n405 585
R1004 B.n404 B.n234 585
R1005 B.n403 B.n402 585
R1006 B.n400 B.n235 585
R1007 B.n398 B.n397 585
R1008 B.n396 B.n236 585
R1009 B.n395 B.n394 585
R1010 B.n392 B.n237 585
R1011 B.n390 B.n389 585
R1012 B.n388 B.n238 585
R1013 B.n387 B.n386 585
R1014 B.n384 B.n239 585
R1015 B.n382 B.n381 585
R1016 B.n380 B.n240 585
R1017 B.n379 B.n378 585
R1018 B.n376 B.n241 585
R1019 B.n374 B.n373 585
R1020 B.n372 B.n242 585
R1021 B.n371 B.n370 585
R1022 B.n368 B.n243 585
R1023 B.n366 B.n365 585
R1024 B.n364 B.n244 585
R1025 B.n363 B.n362 585
R1026 B.n360 B.n245 585
R1027 B.n358 B.n357 585
R1028 B.n356 B.n246 585
R1029 B.n354 B.n353 585
R1030 B.n351 B.n249 585
R1031 B.n349 B.n348 585
R1032 B.n347 B.n250 585
R1033 B.n346 B.n345 585
R1034 B.n343 B.n251 585
R1035 B.n341 B.n340 585
R1036 B.n339 B.n252 585
R1037 B.n338 B.n337 585
R1038 B.n335 B.n253 585
R1039 B.n333 B.n332 585
R1040 B.n331 B.n254 585
R1041 B.n330 B.n329 585
R1042 B.n327 B.n258 585
R1043 B.n325 B.n324 585
R1044 B.n323 B.n259 585
R1045 B.n322 B.n321 585
R1046 B.n319 B.n260 585
R1047 B.n317 B.n316 585
R1048 B.n315 B.n261 585
R1049 B.n314 B.n313 585
R1050 B.n311 B.n262 585
R1051 B.n309 B.n308 585
R1052 B.n307 B.n263 585
R1053 B.n306 B.n305 585
R1054 B.n303 B.n264 585
R1055 B.n301 B.n300 585
R1056 B.n299 B.n265 585
R1057 B.n298 B.n297 585
R1058 B.n295 B.n266 585
R1059 B.n293 B.n292 585
R1060 B.n291 B.n267 585
R1061 B.n290 B.n289 585
R1062 B.n287 B.n268 585
R1063 B.n285 B.n284 585
R1064 B.n283 B.n269 585
R1065 B.n282 B.n281 585
R1066 B.n279 B.n270 585
R1067 B.n277 B.n276 585
R1068 B.n275 B.n271 585
R1069 B.n274 B.n273 585
R1070 B.n228 B.n227 585
R1071 B.n229 B.n228 585
R1072 B.n419 B.n418 585
R1073 B.n420 B.n419 585
R1074 B.n224 B.n223 585
R1075 B.n225 B.n224 585
R1076 B.n428 B.n427 585
R1077 B.n427 B.n426 585
R1078 B.n429 B.n222 585
R1079 B.n222 B.n221 585
R1080 B.n431 B.n430 585
R1081 B.n432 B.n431 585
R1082 B.n216 B.n215 585
R1083 B.n217 B.n216 585
R1084 B.n441 B.n440 585
R1085 B.n440 B.n439 585
R1086 B.n442 B.n214 585
R1087 B.n438 B.n214 585
R1088 B.n444 B.n443 585
R1089 B.n445 B.n444 585
R1090 B.n209 B.n208 585
R1091 B.n210 B.n209 585
R1092 B.n453 B.n452 585
R1093 B.n452 B.n451 585
R1094 B.n454 B.n207 585
R1095 B.n207 B.n206 585
R1096 B.n456 B.n455 585
R1097 B.n457 B.n456 585
R1098 B.n201 B.n200 585
R1099 B.n202 B.n201 585
R1100 B.n465 B.n464 585
R1101 B.n464 B.n463 585
R1102 B.n466 B.n199 585
R1103 B.n199 B.n198 585
R1104 B.n468 B.n467 585
R1105 B.n469 B.n468 585
R1106 B.n193 B.n192 585
R1107 B.n194 B.n193 585
R1108 B.n478 B.n477 585
R1109 B.n477 B.n476 585
R1110 B.n479 B.n191 585
R1111 B.n475 B.n191 585
R1112 B.n481 B.n480 585
R1113 B.n482 B.n481 585
R1114 B.n186 B.n185 585
R1115 B.n187 B.n186 585
R1116 B.n490 B.n489 585
R1117 B.n489 B.n488 585
R1118 B.n491 B.n184 585
R1119 B.n184 B.n183 585
R1120 B.n493 B.n492 585
R1121 B.n494 B.n493 585
R1122 B.n178 B.n177 585
R1123 B.n179 B.n178 585
R1124 B.n503 B.n502 585
R1125 B.n502 B.n501 585
R1126 B.n504 B.n176 585
R1127 B.n500 B.n176 585
R1128 B.n506 B.n505 585
R1129 B.n507 B.n506 585
R1130 B.n171 B.n170 585
R1131 B.n172 B.n171 585
R1132 B.n515 B.n514 585
R1133 B.n514 B.n513 585
R1134 B.n516 B.n169 585
R1135 B.n169 B.n168 585
R1136 B.n518 B.n517 585
R1137 B.n519 B.n518 585
R1138 B.n163 B.n162 585
R1139 B.n164 B.n163 585
R1140 B.n528 B.n527 585
R1141 B.n527 B.n526 585
R1142 B.n529 B.n161 585
R1143 B.n525 B.n161 585
R1144 B.n531 B.n530 585
R1145 B.n532 B.n531 585
R1146 B.n156 B.n155 585
R1147 B.n157 B.n156 585
R1148 B.n540 B.n539 585
R1149 B.n539 B.n538 585
R1150 B.n541 B.n154 585
R1151 B.n154 B.n153 585
R1152 B.n543 B.n542 585
R1153 B.n544 B.n543 585
R1154 B.n148 B.n147 585
R1155 B.n149 B.n148 585
R1156 B.n552 B.n551 585
R1157 B.n551 B.n550 585
R1158 B.n553 B.n146 585
R1159 B.n146 B.n145 585
R1160 B.n555 B.n554 585
R1161 B.n556 B.n555 585
R1162 B.n140 B.n139 585
R1163 B.n141 B.n140 585
R1164 B.n565 B.n564 585
R1165 B.n564 B.n563 585
R1166 B.n566 B.n138 585
R1167 B.n138 B.n137 585
R1168 B.n568 B.n567 585
R1169 B.n569 B.n568 585
R1170 B.n2 B.n0 585
R1171 B.n4 B.n2 585
R1172 B.n3 B.n1 585
R1173 B.n884 B.n3 585
R1174 B.n882 B.n881 585
R1175 B.n883 B.n882 585
R1176 B.n880 B.n9 585
R1177 B.n9 B.n8 585
R1178 B.n879 B.n878 585
R1179 B.n878 B.n877 585
R1180 B.n11 B.n10 585
R1181 B.n876 B.n11 585
R1182 B.n874 B.n873 585
R1183 B.n875 B.n874 585
R1184 B.n872 B.n16 585
R1185 B.n16 B.n15 585
R1186 B.n871 B.n870 585
R1187 B.n870 B.n869 585
R1188 B.n18 B.n17 585
R1189 B.n868 B.n18 585
R1190 B.n866 B.n865 585
R1191 B.n867 B.n866 585
R1192 B.n864 B.n23 585
R1193 B.n23 B.n22 585
R1194 B.n863 B.n862 585
R1195 B.n862 B.n861 585
R1196 B.n25 B.n24 585
R1197 B.n860 B.n25 585
R1198 B.n858 B.n857 585
R1199 B.n859 B.n858 585
R1200 B.n856 B.n29 585
R1201 B.n32 B.n29 585
R1202 B.n855 B.n854 585
R1203 B.n854 B.n853 585
R1204 B.n31 B.n30 585
R1205 B.n852 B.n31 585
R1206 B.n850 B.n849 585
R1207 B.n851 B.n850 585
R1208 B.n848 B.n37 585
R1209 B.n37 B.n36 585
R1210 B.n847 B.n846 585
R1211 B.n846 B.n845 585
R1212 B.n39 B.n38 585
R1213 B.n844 B.n39 585
R1214 B.n842 B.n841 585
R1215 B.n843 B.n842 585
R1216 B.n840 B.n43 585
R1217 B.n46 B.n43 585
R1218 B.n839 B.n838 585
R1219 B.n838 B.n837 585
R1220 B.n45 B.n44 585
R1221 B.n836 B.n45 585
R1222 B.n834 B.n833 585
R1223 B.n835 B.n834 585
R1224 B.n832 B.n51 585
R1225 B.n51 B.n50 585
R1226 B.n831 B.n830 585
R1227 B.n830 B.n829 585
R1228 B.n53 B.n52 585
R1229 B.n828 B.n53 585
R1230 B.n826 B.n825 585
R1231 B.n827 B.n826 585
R1232 B.n824 B.n57 585
R1233 B.n60 B.n57 585
R1234 B.n823 B.n822 585
R1235 B.n822 B.n821 585
R1236 B.n59 B.n58 585
R1237 B.n820 B.n59 585
R1238 B.n818 B.n817 585
R1239 B.n819 B.n818 585
R1240 B.n816 B.n65 585
R1241 B.n65 B.n64 585
R1242 B.n815 B.n814 585
R1243 B.n814 B.n813 585
R1244 B.n67 B.n66 585
R1245 B.n812 B.n67 585
R1246 B.n810 B.n809 585
R1247 B.n811 B.n810 585
R1248 B.n808 B.n72 585
R1249 B.n72 B.n71 585
R1250 B.n807 B.n806 585
R1251 B.n806 B.n805 585
R1252 B.n74 B.n73 585
R1253 B.n804 B.n74 585
R1254 B.n802 B.n801 585
R1255 B.n803 B.n802 585
R1256 B.n800 B.n78 585
R1257 B.n81 B.n78 585
R1258 B.n799 B.n798 585
R1259 B.n798 B.n797 585
R1260 B.n80 B.n79 585
R1261 B.n796 B.n80 585
R1262 B.n794 B.n793 585
R1263 B.n795 B.n794 585
R1264 B.n792 B.n86 585
R1265 B.n86 B.n85 585
R1266 B.n791 B.n790 585
R1267 B.n790 B.n789 585
R1268 B.n88 B.n87 585
R1269 B.n788 B.n88 585
R1270 B.n786 B.n785 585
R1271 B.n787 B.n786 585
R1272 B.n887 B.n886 585
R1273 B.n886 B.n885 585
R1274 B.n419 B.n230 487.695
R1275 B.n786 B.n93 487.695
R1276 B.n421 B.n228 487.695
R1277 B.n637 B.n91 487.695
R1278 B.n255 B.t8 291.795
R1279 B.n247 B.t12 291.795
R1280 B.n110 B.t19 291.795
R1281 B.n116 B.t15 291.795
R1282 B.n255 B.t11 282.019
R1283 B.n116 B.t17 282.019
R1284 B.n247 B.t14 282.019
R1285 B.n110 B.t20 282.019
R1286 B.n638 B.n92 256.663
R1287 B.n640 B.n92 256.663
R1288 B.n646 B.n92 256.663
R1289 B.n648 B.n92 256.663
R1290 B.n654 B.n92 256.663
R1291 B.n656 B.n92 256.663
R1292 B.n662 B.n92 256.663
R1293 B.n664 B.n92 256.663
R1294 B.n670 B.n92 256.663
R1295 B.n672 B.n92 256.663
R1296 B.n678 B.n92 256.663
R1297 B.n680 B.n92 256.663
R1298 B.n686 B.n92 256.663
R1299 B.n688 B.n92 256.663
R1300 B.n694 B.n92 256.663
R1301 B.n119 B.n92 256.663
R1302 B.n700 B.n92 256.663
R1303 B.n706 B.n92 256.663
R1304 B.n708 B.n92 256.663
R1305 B.n714 B.n92 256.663
R1306 B.n716 B.n92 256.663
R1307 B.n723 B.n92 256.663
R1308 B.n725 B.n92 256.663
R1309 B.n731 B.n92 256.663
R1310 B.n733 B.n92 256.663
R1311 B.n739 B.n92 256.663
R1312 B.n741 B.n92 256.663
R1313 B.n747 B.n92 256.663
R1314 B.n749 B.n92 256.663
R1315 B.n755 B.n92 256.663
R1316 B.n757 B.n92 256.663
R1317 B.n763 B.n92 256.663
R1318 B.n765 B.n92 256.663
R1319 B.n771 B.n92 256.663
R1320 B.n773 B.n92 256.663
R1321 B.n779 B.n92 256.663
R1322 B.n781 B.n92 256.663
R1323 B.n414 B.n229 256.663
R1324 B.n232 B.n229 256.663
R1325 B.n407 B.n229 256.663
R1326 B.n401 B.n229 256.663
R1327 B.n399 B.n229 256.663
R1328 B.n393 B.n229 256.663
R1329 B.n391 B.n229 256.663
R1330 B.n385 B.n229 256.663
R1331 B.n383 B.n229 256.663
R1332 B.n377 B.n229 256.663
R1333 B.n375 B.n229 256.663
R1334 B.n369 B.n229 256.663
R1335 B.n367 B.n229 256.663
R1336 B.n361 B.n229 256.663
R1337 B.n359 B.n229 256.663
R1338 B.n352 B.n229 256.663
R1339 B.n350 B.n229 256.663
R1340 B.n344 B.n229 256.663
R1341 B.n342 B.n229 256.663
R1342 B.n336 B.n229 256.663
R1343 B.n334 B.n229 256.663
R1344 B.n328 B.n229 256.663
R1345 B.n326 B.n229 256.663
R1346 B.n320 B.n229 256.663
R1347 B.n318 B.n229 256.663
R1348 B.n312 B.n229 256.663
R1349 B.n310 B.n229 256.663
R1350 B.n304 B.n229 256.663
R1351 B.n302 B.n229 256.663
R1352 B.n296 B.n229 256.663
R1353 B.n294 B.n229 256.663
R1354 B.n288 B.n229 256.663
R1355 B.n286 B.n229 256.663
R1356 B.n280 B.n229 256.663
R1357 B.n278 B.n229 256.663
R1358 B.n272 B.n229 256.663
R1359 B.n256 B.t10 226.745
R1360 B.n117 B.t18 226.745
R1361 B.n248 B.t13 226.745
R1362 B.n111 B.t21 226.745
R1363 B.n419 B.n224 163.367
R1364 B.n427 B.n224 163.367
R1365 B.n427 B.n222 163.367
R1366 B.n431 B.n222 163.367
R1367 B.n431 B.n216 163.367
R1368 B.n440 B.n216 163.367
R1369 B.n440 B.n214 163.367
R1370 B.n444 B.n214 163.367
R1371 B.n444 B.n209 163.367
R1372 B.n452 B.n209 163.367
R1373 B.n452 B.n207 163.367
R1374 B.n456 B.n207 163.367
R1375 B.n456 B.n201 163.367
R1376 B.n464 B.n201 163.367
R1377 B.n464 B.n199 163.367
R1378 B.n468 B.n199 163.367
R1379 B.n468 B.n193 163.367
R1380 B.n477 B.n193 163.367
R1381 B.n477 B.n191 163.367
R1382 B.n481 B.n191 163.367
R1383 B.n481 B.n186 163.367
R1384 B.n489 B.n186 163.367
R1385 B.n489 B.n184 163.367
R1386 B.n493 B.n184 163.367
R1387 B.n493 B.n178 163.367
R1388 B.n502 B.n178 163.367
R1389 B.n502 B.n176 163.367
R1390 B.n506 B.n176 163.367
R1391 B.n506 B.n171 163.367
R1392 B.n514 B.n171 163.367
R1393 B.n514 B.n169 163.367
R1394 B.n518 B.n169 163.367
R1395 B.n518 B.n163 163.367
R1396 B.n527 B.n163 163.367
R1397 B.n527 B.n161 163.367
R1398 B.n531 B.n161 163.367
R1399 B.n531 B.n156 163.367
R1400 B.n539 B.n156 163.367
R1401 B.n539 B.n154 163.367
R1402 B.n543 B.n154 163.367
R1403 B.n543 B.n148 163.367
R1404 B.n551 B.n148 163.367
R1405 B.n551 B.n146 163.367
R1406 B.n555 B.n146 163.367
R1407 B.n555 B.n140 163.367
R1408 B.n564 B.n140 163.367
R1409 B.n564 B.n138 163.367
R1410 B.n568 B.n138 163.367
R1411 B.n568 B.n2 163.367
R1412 B.n886 B.n2 163.367
R1413 B.n886 B.n3 163.367
R1414 B.n882 B.n3 163.367
R1415 B.n882 B.n9 163.367
R1416 B.n878 B.n9 163.367
R1417 B.n878 B.n11 163.367
R1418 B.n874 B.n11 163.367
R1419 B.n874 B.n16 163.367
R1420 B.n870 B.n16 163.367
R1421 B.n870 B.n18 163.367
R1422 B.n866 B.n18 163.367
R1423 B.n866 B.n23 163.367
R1424 B.n862 B.n23 163.367
R1425 B.n862 B.n25 163.367
R1426 B.n858 B.n25 163.367
R1427 B.n858 B.n29 163.367
R1428 B.n854 B.n29 163.367
R1429 B.n854 B.n31 163.367
R1430 B.n850 B.n31 163.367
R1431 B.n850 B.n37 163.367
R1432 B.n846 B.n37 163.367
R1433 B.n846 B.n39 163.367
R1434 B.n842 B.n39 163.367
R1435 B.n842 B.n43 163.367
R1436 B.n838 B.n43 163.367
R1437 B.n838 B.n45 163.367
R1438 B.n834 B.n45 163.367
R1439 B.n834 B.n51 163.367
R1440 B.n830 B.n51 163.367
R1441 B.n830 B.n53 163.367
R1442 B.n826 B.n53 163.367
R1443 B.n826 B.n57 163.367
R1444 B.n822 B.n57 163.367
R1445 B.n822 B.n59 163.367
R1446 B.n818 B.n59 163.367
R1447 B.n818 B.n65 163.367
R1448 B.n814 B.n65 163.367
R1449 B.n814 B.n67 163.367
R1450 B.n810 B.n67 163.367
R1451 B.n810 B.n72 163.367
R1452 B.n806 B.n72 163.367
R1453 B.n806 B.n74 163.367
R1454 B.n802 B.n74 163.367
R1455 B.n802 B.n78 163.367
R1456 B.n798 B.n78 163.367
R1457 B.n798 B.n80 163.367
R1458 B.n794 B.n80 163.367
R1459 B.n794 B.n86 163.367
R1460 B.n790 B.n86 163.367
R1461 B.n790 B.n88 163.367
R1462 B.n786 B.n88 163.367
R1463 B.n415 B.n413 163.367
R1464 B.n413 B.n412 163.367
R1465 B.n409 B.n408 163.367
R1466 B.n406 B.n234 163.367
R1467 B.n402 B.n400 163.367
R1468 B.n398 B.n236 163.367
R1469 B.n394 B.n392 163.367
R1470 B.n390 B.n238 163.367
R1471 B.n386 B.n384 163.367
R1472 B.n382 B.n240 163.367
R1473 B.n378 B.n376 163.367
R1474 B.n374 B.n242 163.367
R1475 B.n370 B.n368 163.367
R1476 B.n366 B.n244 163.367
R1477 B.n362 B.n360 163.367
R1478 B.n358 B.n246 163.367
R1479 B.n353 B.n351 163.367
R1480 B.n349 B.n250 163.367
R1481 B.n345 B.n343 163.367
R1482 B.n341 B.n252 163.367
R1483 B.n337 B.n335 163.367
R1484 B.n333 B.n254 163.367
R1485 B.n329 B.n327 163.367
R1486 B.n325 B.n259 163.367
R1487 B.n321 B.n319 163.367
R1488 B.n317 B.n261 163.367
R1489 B.n313 B.n311 163.367
R1490 B.n309 B.n263 163.367
R1491 B.n305 B.n303 163.367
R1492 B.n301 B.n265 163.367
R1493 B.n297 B.n295 163.367
R1494 B.n293 B.n267 163.367
R1495 B.n289 B.n287 163.367
R1496 B.n285 B.n269 163.367
R1497 B.n281 B.n279 163.367
R1498 B.n277 B.n271 163.367
R1499 B.n273 B.n228 163.367
R1500 B.n421 B.n226 163.367
R1501 B.n425 B.n226 163.367
R1502 B.n425 B.n220 163.367
R1503 B.n433 B.n220 163.367
R1504 B.n433 B.n218 163.367
R1505 B.n437 B.n218 163.367
R1506 B.n437 B.n213 163.367
R1507 B.n446 B.n213 163.367
R1508 B.n446 B.n211 163.367
R1509 B.n450 B.n211 163.367
R1510 B.n450 B.n205 163.367
R1511 B.n458 B.n205 163.367
R1512 B.n458 B.n203 163.367
R1513 B.n462 B.n203 163.367
R1514 B.n462 B.n197 163.367
R1515 B.n470 B.n197 163.367
R1516 B.n470 B.n195 163.367
R1517 B.n474 B.n195 163.367
R1518 B.n474 B.n190 163.367
R1519 B.n483 B.n190 163.367
R1520 B.n483 B.n188 163.367
R1521 B.n487 B.n188 163.367
R1522 B.n487 B.n182 163.367
R1523 B.n495 B.n182 163.367
R1524 B.n495 B.n180 163.367
R1525 B.n499 B.n180 163.367
R1526 B.n499 B.n175 163.367
R1527 B.n508 B.n175 163.367
R1528 B.n508 B.n173 163.367
R1529 B.n512 B.n173 163.367
R1530 B.n512 B.n167 163.367
R1531 B.n520 B.n167 163.367
R1532 B.n520 B.n165 163.367
R1533 B.n524 B.n165 163.367
R1534 B.n524 B.n160 163.367
R1535 B.n533 B.n160 163.367
R1536 B.n533 B.n158 163.367
R1537 B.n537 B.n158 163.367
R1538 B.n537 B.n152 163.367
R1539 B.n545 B.n152 163.367
R1540 B.n545 B.n150 163.367
R1541 B.n549 B.n150 163.367
R1542 B.n549 B.n144 163.367
R1543 B.n557 B.n144 163.367
R1544 B.n557 B.n142 163.367
R1545 B.n562 B.n142 163.367
R1546 B.n562 B.n136 163.367
R1547 B.n570 B.n136 163.367
R1548 B.n571 B.n570 163.367
R1549 B.n571 B.n5 163.367
R1550 B.n6 B.n5 163.367
R1551 B.n7 B.n6 163.367
R1552 B.n576 B.n7 163.367
R1553 B.n576 B.n12 163.367
R1554 B.n13 B.n12 163.367
R1555 B.n14 B.n13 163.367
R1556 B.n581 B.n14 163.367
R1557 B.n581 B.n19 163.367
R1558 B.n20 B.n19 163.367
R1559 B.n21 B.n20 163.367
R1560 B.n586 B.n21 163.367
R1561 B.n586 B.n26 163.367
R1562 B.n27 B.n26 163.367
R1563 B.n28 B.n27 163.367
R1564 B.n591 B.n28 163.367
R1565 B.n591 B.n33 163.367
R1566 B.n34 B.n33 163.367
R1567 B.n35 B.n34 163.367
R1568 B.n596 B.n35 163.367
R1569 B.n596 B.n40 163.367
R1570 B.n41 B.n40 163.367
R1571 B.n42 B.n41 163.367
R1572 B.n601 B.n42 163.367
R1573 B.n601 B.n47 163.367
R1574 B.n48 B.n47 163.367
R1575 B.n49 B.n48 163.367
R1576 B.n606 B.n49 163.367
R1577 B.n606 B.n54 163.367
R1578 B.n55 B.n54 163.367
R1579 B.n56 B.n55 163.367
R1580 B.n611 B.n56 163.367
R1581 B.n611 B.n61 163.367
R1582 B.n62 B.n61 163.367
R1583 B.n63 B.n62 163.367
R1584 B.n616 B.n63 163.367
R1585 B.n616 B.n68 163.367
R1586 B.n69 B.n68 163.367
R1587 B.n70 B.n69 163.367
R1588 B.n621 B.n70 163.367
R1589 B.n621 B.n75 163.367
R1590 B.n76 B.n75 163.367
R1591 B.n77 B.n76 163.367
R1592 B.n626 B.n77 163.367
R1593 B.n626 B.n82 163.367
R1594 B.n83 B.n82 163.367
R1595 B.n84 B.n83 163.367
R1596 B.n631 B.n84 163.367
R1597 B.n631 B.n89 163.367
R1598 B.n90 B.n89 163.367
R1599 B.n91 B.n90 163.367
R1600 B.n782 B.n780 163.367
R1601 B.n778 B.n95 163.367
R1602 B.n774 B.n772 163.367
R1603 B.n770 B.n97 163.367
R1604 B.n766 B.n764 163.367
R1605 B.n762 B.n99 163.367
R1606 B.n758 B.n756 163.367
R1607 B.n754 B.n101 163.367
R1608 B.n750 B.n748 163.367
R1609 B.n746 B.n103 163.367
R1610 B.n742 B.n740 163.367
R1611 B.n738 B.n105 163.367
R1612 B.n734 B.n732 163.367
R1613 B.n730 B.n107 163.367
R1614 B.n726 B.n724 163.367
R1615 B.n722 B.n109 163.367
R1616 B.n717 B.n715 163.367
R1617 B.n713 B.n113 163.367
R1618 B.n709 B.n707 163.367
R1619 B.n705 B.n115 163.367
R1620 B.n701 B.n699 163.367
R1621 B.n696 B.n695 163.367
R1622 B.n693 B.n121 163.367
R1623 B.n689 B.n687 163.367
R1624 B.n685 B.n123 163.367
R1625 B.n681 B.n679 163.367
R1626 B.n677 B.n125 163.367
R1627 B.n673 B.n671 163.367
R1628 B.n669 B.n127 163.367
R1629 B.n665 B.n663 163.367
R1630 B.n661 B.n129 163.367
R1631 B.n657 B.n655 163.367
R1632 B.n653 B.n131 163.367
R1633 B.n649 B.n647 163.367
R1634 B.n645 B.n133 163.367
R1635 B.n641 B.n639 163.367
R1636 B.n420 B.n229 97.9001
R1637 B.n787 B.n92 97.9001
R1638 B.n414 B.n230 71.676
R1639 B.n412 B.n232 71.676
R1640 B.n408 B.n407 71.676
R1641 B.n401 B.n234 71.676
R1642 B.n400 B.n399 71.676
R1643 B.n393 B.n236 71.676
R1644 B.n392 B.n391 71.676
R1645 B.n385 B.n238 71.676
R1646 B.n384 B.n383 71.676
R1647 B.n377 B.n240 71.676
R1648 B.n376 B.n375 71.676
R1649 B.n369 B.n242 71.676
R1650 B.n368 B.n367 71.676
R1651 B.n361 B.n244 71.676
R1652 B.n360 B.n359 71.676
R1653 B.n352 B.n246 71.676
R1654 B.n351 B.n350 71.676
R1655 B.n344 B.n250 71.676
R1656 B.n343 B.n342 71.676
R1657 B.n336 B.n252 71.676
R1658 B.n335 B.n334 71.676
R1659 B.n328 B.n254 71.676
R1660 B.n327 B.n326 71.676
R1661 B.n320 B.n259 71.676
R1662 B.n319 B.n318 71.676
R1663 B.n312 B.n261 71.676
R1664 B.n311 B.n310 71.676
R1665 B.n304 B.n263 71.676
R1666 B.n303 B.n302 71.676
R1667 B.n296 B.n265 71.676
R1668 B.n295 B.n294 71.676
R1669 B.n288 B.n267 71.676
R1670 B.n287 B.n286 71.676
R1671 B.n280 B.n269 71.676
R1672 B.n279 B.n278 71.676
R1673 B.n272 B.n271 71.676
R1674 B.n781 B.n93 71.676
R1675 B.n780 B.n779 71.676
R1676 B.n773 B.n95 71.676
R1677 B.n772 B.n771 71.676
R1678 B.n765 B.n97 71.676
R1679 B.n764 B.n763 71.676
R1680 B.n757 B.n99 71.676
R1681 B.n756 B.n755 71.676
R1682 B.n749 B.n101 71.676
R1683 B.n748 B.n747 71.676
R1684 B.n741 B.n103 71.676
R1685 B.n740 B.n739 71.676
R1686 B.n733 B.n105 71.676
R1687 B.n732 B.n731 71.676
R1688 B.n725 B.n107 71.676
R1689 B.n724 B.n723 71.676
R1690 B.n716 B.n109 71.676
R1691 B.n715 B.n714 71.676
R1692 B.n708 B.n113 71.676
R1693 B.n707 B.n706 71.676
R1694 B.n700 B.n115 71.676
R1695 B.n699 B.n119 71.676
R1696 B.n695 B.n694 71.676
R1697 B.n688 B.n121 71.676
R1698 B.n687 B.n686 71.676
R1699 B.n680 B.n123 71.676
R1700 B.n679 B.n678 71.676
R1701 B.n672 B.n125 71.676
R1702 B.n671 B.n670 71.676
R1703 B.n664 B.n127 71.676
R1704 B.n663 B.n662 71.676
R1705 B.n656 B.n129 71.676
R1706 B.n655 B.n654 71.676
R1707 B.n648 B.n131 71.676
R1708 B.n647 B.n646 71.676
R1709 B.n640 B.n133 71.676
R1710 B.n639 B.n638 71.676
R1711 B.n638 B.n637 71.676
R1712 B.n641 B.n640 71.676
R1713 B.n646 B.n645 71.676
R1714 B.n649 B.n648 71.676
R1715 B.n654 B.n653 71.676
R1716 B.n657 B.n656 71.676
R1717 B.n662 B.n661 71.676
R1718 B.n665 B.n664 71.676
R1719 B.n670 B.n669 71.676
R1720 B.n673 B.n672 71.676
R1721 B.n678 B.n677 71.676
R1722 B.n681 B.n680 71.676
R1723 B.n686 B.n685 71.676
R1724 B.n689 B.n688 71.676
R1725 B.n694 B.n693 71.676
R1726 B.n696 B.n119 71.676
R1727 B.n701 B.n700 71.676
R1728 B.n706 B.n705 71.676
R1729 B.n709 B.n708 71.676
R1730 B.n714 B.n713 71.676
R1731 B.n717 B.n716 71.676
R1732 B.n723 B.n722 71.676
R1733 B.n726 B.n725 71.676
R1734 B.n731 B.n730 71.676
R1735 B.n734 B.n733 71.676
R1736 B.n739 B.n738 71.676
R1737 B.n742 B.n741 71.676
R1738 B.n747 B.n746 71.676
R1739 B.n750 B.n749 71.676
R1740 B.n755 B.n754 71.676
R1741 B.n758 B.n757 71.676
R1742 B.n763 B.n762 71.676
R1743 B.n766 B.n765 71.676
R1744 B.n771 B.n770 71.676
R1745 B.n774 B.n773 71.676
R1746 B.n779 B.n778 71.676
R1747 B.n782 B.n781 71.676
R1748 B.n415 B.n414 71.676
R1749 B.n409 B.n232 71.676
R1750 B.n407 B.n406 71.676
R1751 B.n402 B.n401 71.676
R1752 B.n399 B.n398 71.676
R1753 B.n394 B.n393 71.676
R1754 B.n391 B.n390 71.676
R1755 B.n386 B.n385 71.676
R1756 B.n383 B.n382 71.676
R1757 B.n378 B.n377 71.676
R1758 B.n375 B.n374 71.676
R1759 B.n370 B.n369 71.676
R1760 B.n367 B.n366 71.676
R1761 B.n362 B.n361 71.676
R1762 B.n359 B.n358 71.676
R1763 B.n353 B.n352 71.676
R1764 B.n350 B.n349 71.676
R1765 B.n345 B.n344 71.676
R1766 B.n342 B.n341 71.676
R1767 B.n337 B.n336 71.676
R1768 B.n334 B.n333 71.676
R1769 B.n329 B.n328 71.676
R1770 B.n326 B.n325 71.676
R1771 B.n321 B.n320 71.676
R1772 B.n318 B.n317 71.676
R1773 B.n313 B.n312 71.676
R1774 B.n310 B.n309 71.676
R1775 B.n305 B.n304 71.676
R1776 B.n302 B.n301 71.676
R1777 B.n297 B.n296 71.676
R1778 B.n294 B.n293 71.676
R1779 B.n289 B.n288 71.676
R1780 B.n286 B.n285 71.676
R1781 B.n281 B.n280 71.676
R1782 B.n278 B.n277 71.676
R1783 B.n273 B.n272 71.676
R1784 B.n257 B.n256 59.5399
R1785 B.n355 B.n248 59.5399
R1786 B.n720 B.n111 59.5399
R1787 B.n118 B.n117 59.5399
R1788 B.n256 B.n255 55.2732
R1789 B.n248 B.n247 55.2732
R1790 B.n111 B.n110 55.2732
R1791 B.n117 B.n116 55.2732
R1792 B.n420 B.n225 53.2579
R1793 B.n426 B.n225 53.2579
R1794 B.n426 B.n221 53.2579
R1795 B.n432 B.n221 53.2579
R1796 B.n432 B.n217 53.2579
R1797 B.n439 B.n217 53.2579
R1798 B.n439 B.n438 53.2579
R1799 B.n445 B.n210 53.2579
R1800 B.n451 B.n210 53.2579
R1801 B.n451 B.n206 53.2579
R1802 B.n457 B.n206 53.2579
R1803 B.n457 B.n202 53.2579
R1804 B.n463 B.n202 53.2579
R1805 B.n463 B.n198 53.2579
R1806 B.n469 B.n198 53.2579
R1807 B.n469 B.n194 53.2579
R1808 B.n476 B.n194 53.2579
R1809 B.n476 B.n475 53.2579
R1810 B.n482 B.n187 53.2579
R1811 B.n488 B.n187 53.2579
R1812 B.n488 B.n183 53.2579
R1813 B.n494 B.n183 53.2579
R1814 B.n494 B.n179 53.2579
R1815 B.n501 B.n179 53.2579
R1816 B.n501 B.n500 53.2579
R1817 B.n507 B.n172 53.2579
R1818 B.n513 B.n172 53.2579
R1819 B.n513 B.n168 53.2579
R1820 B.n519 B.n168 53.2579
R1821 B.n519 B.n164 53.2579
R1822 B.n526 B.n164 53.2579
R1823 B.n526 B.n525 53.2579
R1824 B.n532 B.n157 53.2579
R1825 B.n538 B.n157 53.2579
R1826 B.n538 B.n153 53.2579
R1827 B.n544 B.n153 53.2579
R1828 B.n544 B.n149 53.2579
R1829 B.n550 B.n149 53.2579
R1830 B.n550 B.n145 53.2579
R1831 B.n556 B.n145 53.2579
R1832 B.n563 B.n141 53.2579
R1833 B.n563 B.n137 53.2579
R1834 B.n569 B.n137 53.2579
R1835 B.n569 B.n4 53.2579
R1836 B.n885 B.n4 53.2579
R1837 B.n885 B.n884 53.2579
R1838 B.n884 B.n883 53.2579
R1839 B.n883 B.n8 53.2579
R1840 B.n877 B.n8 53.2579
R1841 B.n877 B.n876 53.2579
R1842 B.n875 B.n15 53.2579
R1843 B.n869 B.n15 53.2579
R1844 B.n869 B.n868 53.2579
R1845 B.n868 B.n867 53.2579
R1846 B.n867 B.n22 53.2579
R1847 B.n861 B.n22 53.2579
R1848 B.n861 B.n860 53.2579
R1849 B.n860 B.n859 53.2579
R1850 B.n853 B.n32 53.2579
R1851 B.n853 B.n852 53.2579
R1852 B.n852 B.n851 53.2579
R1853 B.n851 B.n36 53.2579
R1854 B.n845 B.n36 53.2579
R1855 B.n845 B.n844 53.2579
R1856 B.n844 B.n843 53.2579
R1857 B.n837 B.n46 53.2579
R1858 B.n837 B.n836 53.2579
R1859 B.n836 B.n835 53.2579
R1860 B.n835 B.n50 53.2579
R1861 B.n829 B.n50 53.2579
R1862 B.n829 B.n828 53.2579
R1863 B.n828 B.n827 53.2579
R1864 B.n821 B.n60 53.2579
R1865 B.n821 B.n820 53.2579
R1866 B.n820 B.n819 53.2579
R1867 B.n819 B.n64 53.2579
R1868 B.n813 B.n64 53.2579
R1869 B.n813 B.n812 53.2579
R1870 B.n812 B.n811 53.2579
R1871 B.n811 B.n71 53.2579
R1872 B.n805 B.n71 53.2579
R1873 B.n805 B.n804 53.2579
R1874 B.n804 B.n803 53.2579
R1875 B.n797 B.n81 53.2579
R1876 B.n797 B.n796 53.2579
R1877 B.n796 B.n795 53.2579
R1878 B.n795 B.n85 53.2579
R1879 B.n789 B.n85 53.2579
R1880 B.n789 B.n788 53.2579
R1881 B.n788 B.n787 53.2579
R1882 B.n482 B.t3 50.1251
R1883 B.n827 B.t0 50.1251
R1884 B.n525 B.t7 43.8595
R1885 B.n32 B.t4 43.8595
R1886 B.t6 B.n141 42.2931
R1887 B.n876 B.t5 42.2931
R1888 B.n785 B.n784 31.6883
R1889 B.n636 B.n635 31.6883
R1890 B.n422 B.n227 31.6883
R1891 B.n418 B.n417 31.6883
R1892 B.n507 B.t1 29.762
R1893 B.n843 B.t2 29.762
R1894 B.n445 B.t9 28.1956
R1895 B.n803 B.t16 28.1956
R1896 B.n438 B.t9 25.0628
R1897 B.n81 B.t16 25.0628
R1898 B.n500 B.t1 23.4964
R1899 B.n46 B.t2 23.4964
R1900 B B.n887 18.0485
R1901 B.n556 B.t6 10.9653
R1902 B.t5 B.n875 10.9653
R1903 B.n784 B.n783 10.6151
R1904 B.n783 B.n94 10.6151
R1905 B.n777 B.n94 10.6151
R1906 B.n777 B.n776 10.6151
R1907 B.n776 B.n775 10.6151
R1908 B.n775 B.n96 10.6151
R1909 B.n769 B.n96 10.6151
R1910 B.n769 B.n768 10.6151
R1911 B.n768 B.n767 10.6151
R1912 B.n767 B.n98 10.6151
R1913 B.n761 B.n98 10.6151
R1914 B.n761 B.n760 10.6151
R1915 B.n760 B.n759 10.6151
R1916 B.n759 B.n100 10.6151
R1917 B.n753 B.n100 10.6151
R1918 B.n753 B.n752 10.6151
R1919 B.n752 B.n751 10.6151
R1920 B.n751 B.n102 10.6151
R1921 B.n745 B.n102 10.6151
R1922 B.n745 B.n744 10.6151
R1923 B.n744 B.n743 10.6151
R1924 B.n743 B.n104 10.6151
R1925 B.n737 B.n104 10.6151
R1926 B.n737 B.n736 10.6151
R1927 B.n736 B.n735 10.6151
R1928 B.n735 B.n106 10.6151
R1929 B.n729 B.n106 10.6151
R1930 B.n729 B.n728 10.6151
R1931 B.n728 B.n727 10.6151
R1932 B.n727 B.n108 10.6151
R1933 B.n721 B.n108 10.6151
R1934 B.n719 B.n718 10.6151
R1935 B.n718 B.n112 10.6151
R1936 B.n712 B.n112 10.6151
R1937 B.n712 B.n711 10.6151
R1938 B.n711 B.n710 10.6151
R1939 B.n710 B.n114 10.6151
R1940 B.n704 B.n114 10.6151
R1941 B.n704 B.n703 10.6151
R1942 B.n703 B.n702 10.6151
R1943 B.n698 B.n697 10.6151
R1944 B.n697 B.n120 10.6151
R1945 B.n692 B.n120 10.6151
R1946 B.n692 B.n691 10.6151
R1947 B.n691 B.n690 10.6151
R1948 B.n690 B.n122 10.6151
R1949 B.n684 B.n122 10.6151
R1950 B.n684 B.n683 10.6151
R1951 B.n683 B.n682 10.6151
R1952 B.n682 B.n124 10.6151
R1953 B.n676 B.n124 10.6151
R1954 B.n676 B.n675 10.6151
R1955 B.n675 B.n674 10.6151
R1956 B.n674 B.n126 10.6151
R1957 B.n668 B.n126 10.6151
R1958 B.n668 B.n667 10.6151
R1959 B.n667 B.n666 10.6151
R1960 B.n666 B.n128 10.6151
R1961 B.n660 B.n128 10.6151
R1962 B.n660 B.n659 10.6151
R1963 B.n659 B.n658 10.6151
R1964 B.n658 B.n130 10.6151
R1965 B.n652 B.n130 10.6151
R1966 B.n652 B.n651 10.6151
R1967 B.n651 B.n650 10.6151
R1968 B.n650 B.n132 10.6151
R1969 B.n644 B.n132 10.6151
R1970 B.n644 B.n643 10.6151
R1971 B.n643 B.n642 10.6151
R1972 B.n642 B.n134 10.6151
R1973 B.n636 B.n134 10.6151
R1974 B.n423 B.n422 10.6151
R1975 B.n424 B.n423 10.6151
R1976 B.n424 B.n219 10.6151
R1977 B.n434 B.n219 10.6151
R1978 B.n435 B.n434 10.6151
R1979 B.n436 B.n435 10.6151
R1980 B.n436 B.n212 10.6151
R1981 B.n447 B.n212 10.6151
R1982 B.n448 B.n447 10.6151
R1983 B.n449 B.n448 10.6151
R1984 B.n449 B.n204 10.6151
R1985 B.n459 B.n204 10.6151
R1986 B.n460 B.n459 10.6151
R1987 B.n461 B.n460 10.6151
R1988 B.n461 B.n196 10.6151
R1989 B.n471 B.n196 10.6151
R1990 B.n472 B.n471 10.6151
R1991 B.n473 B.n472 10.6151
R1992 B.n473 B.n189 10.6151
R1993 B.n484 B.n189 10.6151
R1994 B.n485 B.n484 10.6151
R1995 B.n486 B.n485 10.6151
R1996 B.n486 B.n181 10.6151
R1997 B.n496 B.n181 10.6151
R1998 B.n497 B.n496 10.6151
R1999 B.n498 B.n497 10.6151
R2000 B.n498 B.n174 10.6151
R2001 B.n509 B.n174 10.6151
R2002 B.n510 B.n509 10.6151
R2003 B.n511 B.n510 10.6151
R2004 B.n511 B.n166 10.6151
R2005 B.n521 B.n166 10.6151
R2006 B.n522 B.n521 10.6151
R2007 B.n523 B.n522 10.6151
R2008 B.n523 B.n159 10.6151
R2009 B.n534 B.n159 10.6151
R2010 B.n535 B.n534 10.6151
R2011 B.n536 B.n535 10.6151
R2012 B.n536 B.n151 10.6151
R2013 B.n546 B.n151 10.6151
R2014 B.n547 B.n546 10.6151
R2015 B.n548 B.n547 10.6151
R2016 B.n548 B.n143 10.6151
R2017 B.n558 B.n143 10.6151
R2018 B.n559 B.n558 10.6151
R2019 B.n561 B.n559 10.6151
R2020 B.n561 B.n560 10.6151
R2021 B.n560 B.n135 10.6151
R2022 B.n572 B.n135 10.6151
R2023 B.n573 B.n572 10.6151
R2024 B.n574 B.n573 10.6151
R2025 B.n575 B.n574 10.6151
R2026 B.n577 B.n575 10.6151
R2027 B.n578 B.n577 10.6151
R2028 B.n579 B.n578 10.6151
R2029 B.n580 B.n579 10.6151
R2030 B.n582 B.n580 10.6151
R2031 B.n583 B.n582 10.6151
R2032 B.n584 B.n583 10.6151
R2033 B.n585 B.n584 10.6151
R2034 B.n587 B.n585 10.6151
R2035 B.n588 B.n587 10.6151
R2036 B.n589 B.n588 10.6151
R2037 B.n590 B.n589 10.6151
R2038 B.n592 B.n590 10.6151
R2039 B.n593 B.n592 10.6151
R2040 B.n594 B.n593 10.6151
R2041 B.n595 B.n594 10.6151
R2042 B.n597 B.n595 10.6151
R2043 B.n598 B.n597 10.6151
R2044 B.n599 B.n598 10.6151
R2045 B.n600 B.n599 10.6151
R2046 B.n602 B.n600 10.6151
R2047 B.n603 B.n602 10.6151
R2048 B.n604 B.n603 10.6151
R2049 B.n605 B.n604 10.6151
R2050 B.n607 B.n605 10.6151
R2051 B.n608 B.n607 10.6151
R2052 B.n609 B.n608 10.6151
R2053 B.n610 B.n609 10.6151
R2054 B.n612 B.n610 10.6151
R2055 B.n613 B.n612 10.6151
R2056 B.n614 B.n613 10.6151
R2057 B.n615 B.n614 10.6151
R2058 B.n617 B.n615 10.6151
R2059 B.n618 B.n617 10.6151
R2060 B.n619 B.n618 10.6151
R2061 B.n620 B.n619 10.6151
R2062 B.n622 B.n620 10.6151
R2063 B.n623 B.n622 10.6151
R2064 B.n624 B.n623 10.6151
R2065 B.n625 B.n624 10.6151
R2066 B.n627 B.n625 10.6151
R2067 B.n628 B.n627 10.6151
R2068 B.n629 B.n628 10.6151
R2069 B.n630 B.n629 10.6151
R2070 B.n632 B.n630 10.6151
R2071 B.n633 B.n632 10.6151
R2072 B.n634 B.n633 10.6151
R2073 B.n635 B.n634 10.6151
R2074 B.n417 B.n416 10.6151
R2075 B.n416 B.n231 10.6151
R2076 B.n411 B.n231 10.6151
R2077 B.n411 B.n410 10.6151
R2078 B.n410 B.n233 10.6151
R2079 B.n405 B.n233 10.6151
R2080 B.n405 B.n404 10.6151
R2081 B.n404 B.n403 10.6151
R2082 B.n403 B.n235 10.6151
R2083 B.n397 B.n235 10.6151
R2084 B.n397 B.n396 10.6151
R2085 B.n396 B.n395 10.6151
R2086 B.n395 B.n237 10.6151
R2087 B.n389 B.n237 10.6151
R2088 B.n389 B.n388 10.6151
R2089 B.n388 B.n387 10.6151
R2090 B.n387 B.n239 10.6151
R2091 B.n381 B.n239 10.6151
R2092 B.n381 B.n380 10.6151
R2093 B.n380 B.n379 10.6151
R2094 B.n379 B.n241 10.6151
R2095 B.n373 B.n241 10.6151
R2096 B.n373 B.n372 10.6151
R2097 B.n372 B.n371 10.6151
R2098 B.n371 B.n243 10.6151
R2099 B.n365 B.n243 10.6151
R2100 B.n365 B.n364 10.6151
R2101 B.n364 B.n363 10.6151
R2102 B.n363 B.n245 10.6151
R2103 B.n357 B.n245 10.6151
R2104 B.n357 B.n356 10.6151
R2105 B.n354 B.n249 10.6151
R2106 B.n348 B.n249 10.6151
R2107 B.n348 B.n347 10.6151
R2108 B.n347 B.n346 10.6151
R2109 B.n346 B.n251 10.6151
R2110 B.n340 B.n251 10.6151
R2111 B.n340 B.n339 10.6151
R2112 B.n339 B.n338 10.6151
R2113 B.n338 B.n253 10.6151
R2114 B.n332 B.n331 10.6151
R2115 B.n331 B.n330 10.6151
R2116 B.n330 B.n258 10.6151
R2117 B.n324 B.n258 10.6151
R2118 B.n324 B.n323 10.6151
R2119 B.n323 B.n322 10.6151
R2120 B.n322 B.n260 10.6151
R2121 B.n316 B.n260 10.6151
R2122 B.n316 B.n315 10.6151
R2123 B.n315 B.n314 10.6151
R2124 B.n314 B.n262 10.6151
R2125 B.n308 B.n262 10.6151
R2126 B.n308 B.n307 10.6151
R2127 B.n307 B.n306 10.6151
R2128 B.n306 B.n264 10.6151
R2129 B.n300 B.n264 10.6151
R2130 B.n300 B.n299 10.6151
R2131 B.n299 B.n298 10.6151
R2132 B.n298 B.n266 10.6151
R2133 B.n292 B.n266 10.6151
R2134 B.n292 B.n291 10.6151
R2135 B.n291 B.n290 10.6151
R2136 B.n290 B.n268 10.6151
R2137 B.n284 B.n268 10.6151
R2138 B.n284 B.n283 10.6151
R2139 B.n283 B.n282 10.6151
R2140 B.n282 B.n270 10.6151
R2141 B.n276 B.n270 10.6151
R2142 B.n276 B.n275 10.6151
R2143 B.n275 B.n274 10.6151
R2144 B.n274 B.n227 10.6151
R2145 B.n418 B.n223 10.6151
R2146 B.n428 B.n223 10.6151
R2147 B.n429 B.n428 10.6151
R2148 B.n430 B.n429 10.6151
R2149 B.n430 B.n215 10.6151
R2150 B.n441 B.n215 10.6151
R2151 B.n442 B.n441 10.6151
R2152 B.n443 B.n442 10.6151
R2153 B.n443 B.n208 10.6151
R2154 B.n453 B.n208 10.6151
R2155 B.n454 B.n453 10.6151
R2156 B.n455 B.n454 10.6151
R2157 B.n455 B.n200 10.6151
R2158 B.n465 B.n200 10.6151
R2159 B.n466 B.n465 10.6151
R2160 B.n467 B.n466 10.6151
R2161 B.n467 B.n192 10.6151
R2162 B.n478 B.n192 10.6151
R2163 B.n479 B.n478 10.6151
R2164 B.n480 B.n479 10.6151
R2165 B.n480 B.n185 10.6151
R2166 B.n490 B.n185 10.6151
R2167 B.n491 B.n490 10.6151
R2168 B.n492 B.n491 10.6151
R2169 B.n492 B.n177 10.6151
R2170 B.n503 B.n177 10.6151
R2171 B.n504 B.n503 10.6151
R2172 B.n505 B.n504 10.6151
R2173 B.n505 B.n170 10.6151
R2174 B.n515 B.n170 10.6151
R2175 B.n516 B.n515 10.6151
R2176 B.n517 B.n516 10.6151
R2177 B.n517 B.n162 10.6151
R2178 B.n528 B.n162 10.6151
R2179 B.n529 B.n528 10.6151
R2180 B.n530 B.n529 10.6151
R2181 B.n530 B.n155 10.6151
R2182 B.n540 B.n155 10.6151
R2183 B.n541 B.n540 10.6151
R2184 B.n542 B.n541 10.6151
R2185 B.n542 B.n147 10.6151
R2186 B.n552 B.n147 10.6151
R2187 B.n553 B.n552 10.6151
R2188 B.n554 B.n553 10.6151
R2189 B.n554 B.n139 10.6151
R2190 B.n565 B.n139 10.6151
R2191 B.n566 B.n565 10.6151
R2192 B.n567 B.n566 10.6151
R2193 B.n567 B.n0 10.6151
R2194 B.n881 B.n1 10.6151
R2195 B.n881 B.n880 10.6151
R2196 B.n880 B.n879 10.6151
R2197 B.n879 B.n10 10.6151
R2198 B.n873 B.n10 10.6151
R2199 B.n873 B.n872 10.6151
R2200 B.n872 B.n871 10.6151
R2201 B.n871 B.n17 10.6151
R2202 B.n865 B.n17 10.6151
R2203 B.n865 B.n864 10.6151
R2204 B.n864 B.n863 10.6151
R2205 B.n863 B.n24 10.6151
R2206 B.n857 B.n24 10.6151
R2207 B.n857 B.n856 10.6151
R2208 B.n856 B.n855 10.6151
R2209 B.n855 B.n30 10.6151
R2210 B.n849 B.n30 10.6151
R2211 B.n849 B.n848 10.6151
R2212 B.n848 B.n847 10.6151
R2213 B.n847 B.n38 10.6151
R2214 B.n841 B.n38 10.6151
R2215 B.n841 B.n840 10.6151
R2216 B.n840 B.n839 10.6151
R2217 B.n839 B.n44 10.6151
R2218 B.n833 B.n44 10.6151
R2219 B.n833 B.n832 10.6151
R2220 B.n832 B.n831 10.6151
R2221 B.n831 B.n52 10.6151
R2222 B.n825 B.n52 10.6151
R2223 B.n825 B.n824 10.6151
R2224 B.n824 B.n823 10.6151
R2225 B.n823 B.n58 10.6151
R2226 B.n817 B.n58 10.6151
R2227 B.n817 B.n816 10.6151
R2228 B.n816 B.n815 10.6151
R2229 B.n815 B.n66 10.6151
R2230 B.n809 B.n66 10.6151
R2231 B.n809 B.n808 10.6151
R2232 B.n808 B.n807 10.6151
R2233 B.n807 B.n73 10.6151
R2234 B.n801 B.n73 10.6151
R2235 B.n801 B.n800 10.6151
R2236 B.n800 B.n799 10.6151
R2237 B.n799 B.n79 10.6151
R2238 B.n793 B.n79 10.6151
R2239 B.n793 B.n792 10.6151
R2240 B.n792 B.n791 10.6151
R2241 B.n791 B.n87 10.6151
R2242 B.n785 B.n87 10.6151
R2243 B.n532 B.t7 9.39886
R2244 B.n859 B.t4 9.39886
R2245 B.n721 B.n720 9.36635
R2246 B.n698 B.n118 9.36635
R2247 B.n356 B.n355 9.36635
R2248 B.n332 B.n257 9.36635
R2249 B.n475 B.t3 3.13329
R2250 B.n60 B.t0 3.13329
R2251 B.n887 B.n0 2.81026
R2252 B.n887 B.n1 2.81026
R2253 B.n720 B.n719 1.24928
R2254 B.n702 B.n118 1.24928
R2255 B.n355 B.n354 1.24928
R2256 B.n257 B.n253 1.24928
R2257 VN.n51 VN.n27 161.3
R2258 VN.n50 VN.n49 161.3
R2259 VN.n48 VN.n28 161.3
R2260 VN.n47 VN.n46 161.3
R2261 VN.n45 VN.n29 161.3
R2262 VN.n44 VN.n43 161.3
R2263 VN.n42 VN.n41 161.3
R2264 VN.n40 VN.n31 161.3
R2265 VN.n39 VN.n38 161.3
R2266 VN.n37 VN.n32 161.3
R2267 VN.n36 VN.n35 161.3
R2268 VN.n24 VN.n0 161.3
R2269 VN.n23 VN.n22 161.3
R2270 VN.n21 VN.n1 161.3
R2271 VN.n20 VN.n19 161.3
R2272 VN.n18 VN.n2 161.3
R2273 VN.n17 VN.n16 161.3
R2274 VN.n15 VN.n14 161.3
R2275 VN.n13 VN.n4 161.3
R2276 VN.n12 VN.n11 161.3
R2277 VN.n10 VN.n5 161.3
R2278 VN.n9 VN.n8 161.3
R2279 VN.n6 VN.t3 118.445
R2280 VN.n33 VN.t6 118.445
R2281 VN.n26 VN.n25 97.2996
R2282 VN.n53 VN.n52 97.2996
R2283 VN.n7 VN.t7 83.8723
R2284 VN.n3 VN.t2 83.8723
R2285 VN.n25 VN.t5 83.8723
R2286 VN.n34 VN.t4 83.8723
R2287 VN.n30 VN.t1 83.8723
R2288 VN.n52 VN.t0 83.8723
R2289 VN.n19 VN.n1 55.0624
R2290 VN.n46 VN.n28 55.0624
R2291 VN.n7 VN.n6 51.8291
R2292 VN.n34 VN.n33 51.8291
R2293 VN VN.n53 48.4072
R2294 VN.n12 VN.n5 40.4934
R2295 VN.n13 VN.n12 40.4934
R2296 VN.n39 VN.n32 40.4934
R2297 VN.n40 VN.n39 40.4934
R2298 VN.n23 VN.n1 25.9244
R2299 VN.n50 VN.n28 25.9244
R2300 VN.n8 VN.n5 24.4675
R2301 VN.n14 VN.n13 24.4675
R2302 VN.n18 VN.n17 24.4675
R2303 VN.n19 VN.n18 24.4675
R2304 VN.n24 VN.n23 24.4675
R2305 VN.n35 VN.n32 24.4675
R2306 VN.n46 VN.n45 24.4675
R2307 VN.n45 VN.n44 24.4675
R2308 VN.n41 VN.n40 24.4675
R2309 VN.n51 VN.n50 24.4675
R2310 VN.n8 VN.n7 20.7975
R2311 VN.n14 VN.n3 20.7975
R2312 VN.n35 VN.n34 20.7975
R2313 VN.n41 VN.n30 20.7975
R2314 VN.n25 VN.n24 13.4574
R2315 VN.n52 VN.n51 13.4574
R2316 VN.n36 VN.n33 6.62497
R2317 VN.n9 VN.n6 6.62497
R2318 VN.n17 VN.n3 3.67055
R2319 VN.n44 VN.n30 3.67055
R2320 VN.n53 VN.n27 0.278367
R2321 VN.n26 VN.n0 0.278367
R2322 VN.n49 VN.n27 0.189894
R2323 VN.n49 VN.n48 0.189894
R2324 VN.n48 VN.n47 0.189894
R2325 VN.n47 VN.n29 0.189894
R2326 VN.n43 VN.n29 0.189894
R2327 VN.n43 VN.n42 0.189894
R2328 VN.n42 VN.n31 0.189894
R2329 VN.n38 VN.n31 0.189894
R2330 VN.n38 VN.n37 0.189894
R2331 VN.n37 VN.n36 0.189894
R2332 VN.n10 VN.n9 0.189894
R2333 VN.n11 VN.n10 0.189894
R2334 VN.n11 VN.n4 0.189894
R2335 VN.n15 VN.n4 0.189894
R2336 VN.n16 VN.n15 0.189894
R2337 VN.n16 VN.n2 0.189894
R2338 VN.n20 VN.n2 0.189894
R2339 VN.n21 VN.n20 0.189894
R2340 VN.n22 VN.n21 0.189894
R2341 VN.n22 VN.n0 0.189894
R2342 VN VN.n26 0.153454
R2343 VDD2.n2 VDD2.n1 62.9777
R2344 VDD2.n2 VDD2.n0 62.9777
R2345 VDD2 VDD2.n5 62.9751
R2346 VDD2.n4 VDD2.n3 61.8048
R2347 VDD2.n4 VDD2.n2 42.3317
R2348 VDD2.n5 VDD2.t3 2.2582
R2349 VDD2.n5 VDD2.t1 2.2582
R2350 VDD2.n3 VDD2.t7 2.2582
R2351 VDD2.n3 VDD2.t6 2.2582
R2352 VDD2.n1 VDD2.t5 2.2582
R2353 VDD2.n1 VDD2.t2 2.2582
R2354 VDD2.n0 VDD2.t4 2.2582
R2355 VDD2.n0 VDD2.t0 2.2582
R2356 VDD2 VDD2.n4 1.28714
C0 VP VN 6.96432f
C1 VDD2 VN 6.42999f
C2 VP VTAIL 6.96298f
C3 VDD2 VTAIL 7.0141f
C4 VDD1 VN 0.151616f
C5 VDD1 VTAIL 6.96022f
C6 VN VTAIL 6.94887f
C7 VDD2 VP 0.51119f
C8 VDD1 VP 6.78821f
C9 VDD1 VDD2 1.73595f
C10 VDD2 B 5.023541f
C11 VDD1 B 5.459256f
C12 VTAIL B 8.498678f
C13 VN B 14.931411f
C14 VP B 13.554389f
C15 VDD2.t4 B 0.167731f
C16 VDD2.t0 B 0.167731f
C17 VDD2.n0 B 1.46215f
C18 VDD2.t5 B 0.167731f
C19 VDD2.t2 B 0.167731f
C20 VDD2.n1 B 1.46215f
C21 VDD2.n2 B 2.94506f
C22 VDD2.t7 B 0.167731f
C23 VDD2.t6 B 0.167731f
C24 VDD2.n3 B 1.45288f
C25 VDD2.n4 B 2.59412f
C26 VDD2.t3 B 0.167731f
C27 VDD2.t1 B 0.167731f
C28 VDD2.n5 B 1.46212f
C29 VN.n0 B 0.030968f
C30 VN.t5 B 1.3995f
C31 VN.n1 B 0.026785f
C32 VN.n2 B 0.023489f
C33 VN.t2 B 1.3995f
C34 VN.n3 B 0.506541f
C35 VN.n4 B 0.023489f
C36 VN.n5 B 0.046684f
C37 VN.t3 B 1.58963f
C38 VN.n6 B 0.551803f
C39 VN.t7 B 1.3995f
C40 VN.n7 B 0.581621f
C41 VN.n8 B 0.040534f
C42 VN.n9 B 0.225063f
C43 VN.n10 B 0.023489f
C44 VN.n11 B 0.023489f
C45 VN.n12 B 0.018988f
C46 VN.n13 B 0.046684f
C47 VN.n14 B 0.040534f
C48 VN.n15 B 0.023489f
C49 VN.n16 B 0.023489f
C50 VN.n17 B 0.025405f
C51 VN.n18 B 0.043777f
C52 VN.n19 B 0.040653f
C53 VN.n20 B 0.023489f
C54 VN.n21 B 0.023489f
C55 VN.n22 B 0.023489f
C56 VN.n23 B 0.044918f
C57 VN.n24 B 0.03405f
C58 VN.n25 B 0.587504f
C59 VN.n26 B 0.035439f
C60 VN.n27 B 0.030968f
C61 VN.t0 B 1.3995f
C62 VN.n28 B 0.026785f
C63 VN.n29 B 0.023489f
C64 VN.t1 B 1.3995f
C65 VN.n30 B 0.506541f
C66 VN.n31 B 0.023489f
C67 VN.n32 B 0.046684f
C68 VN.t6 B 1.58963f
C69 VN.n33 B 0.551803f
C70 VN.t4 B 1.3995f
C71 VN.n34 B 0.581621f
C72 VN.n35 B 0.040534f
C73 VN.n36 B 0.225063f
C74 VN.n37 B 0.023489f
C75 VN.n38 B 0.023489f
C76 VN.n39 B 0.018988f
C77 VN.n40 B 0.046684f
C78 VN.n41 B 0.040534f
C79 VN.n42 B 0.023489f
C80 VN.n43 B 0.023489f
C81 VN.n44 B 0.025405f
C82 VN.n45 B 0.043777f
C83 VN.n46 B 0.040653f
C84 VN.n47 B 0.023489f
C85 VN.n48 B 0.023489f
C86 VN.n49 B 0.023489f
C87 VN.n50 B 0.044918f
C88 VN.n51 B 0.03405f
C89 VN.n52 B 0.587504f
C90 VN.n53 B 1.24538f
C91 VDD1.t3 B 0.171593f
C92 VDD1.t4 B 0.171593f
C93 VDD1.n0 B 1.4969f
C94 VDD1.t0 B 0.171593f
C95 VDD1.t2 B 0.171593f
C96 VDD1.n1 B 1.49582f
C97 VDD1.t6 B 0.171593f
C98 VDD1.t1 B 0.171593f
C99 VDD1.n2 B 1.49582f
C100 VDD1.n3 B 3.0646f
C101 VDD1.t5 B 0.171593f
C102 VDD1.t7 B 0.171593f
C103 VDD1.n4 B 1.48633f
C104 VDD1.n5 B 2.68429f
C105 VTAIL.t4 B 0.14556f
C106 VTAIL.t2 B 0.14556f
C107 VTAIL.n0 B 1.19665f
C108 VTAIL.n1 B 0.38349f
C109 VTAIL.n2 B 0.030231f
C110 VTAIL.n3 B 0.021003f
C111 VTAIL.n4 B 0.011286f
C112 VTAIL.n5 B 0.026677f
C113 VTAIL.n6 B 0.01195f
C114 VTAIL.n7 B 0.021003f
C115 VTAIL.n8 B 0.011286f
C116 VTAIL.n9 B 0.026677f
C117 VTAIL.n10 B 0.01195f
C118 VTAIL.n11 B 0.021003f
C119 VTAIL.n12 B 0.011286f
C120 VTAIL.n13 B 0.026677f
C121 VTAIL.n14 B 0.01195f
C122 VTAIL.n15 B 0.766789f
C123 VTAIL.n16 B 0.011286f
C124 VTAIL.t5 B 0.043547f
C125 VTAIL.n17 B 0.1042f
C126 VTAIL.n18 B 0.015759f
C127 VTAIL.n19 B 0.020007f
C128 VTAIL.n20 B 0.026677f
C129 VTAIL.n21 B 0.01195f
C130 VTAIL.n22 B 0.011286f
C131 VTAIL.n23 B 0.021003f
C132 VTAIL.n24 B 0.021003f
C133 VTAIL.n25 B 0.011286f
C134 VTAIL.n26 B 0.01195f
C135 VTAIL.n27 B 0.026677f
C136 VTAIL.n28 B 0.026677f
C137 VTAIL.n29 B 0.01195f
C138 VTAIL.n30 B 0.011286f
C139 VTAIL.n31 B 0.021003f
C140 VTAIL.n32 B 0.021003f
C141 VTAIL.n33 B 0.011286f
C142 VTAIL.n34 B 0.01195f
C143 VTAIL.n35 B 0.026677f
C144 VTAIL.n36 B 0.026677f
C145 VTAIL.n37 B 0.01195f
C146 VTAIL.n38 B 0.011286f
C147 VTAIL.n39 B 0.021003f
C148 VTAIL.n40 B 0.021003f
C149 VTAIL.n41 B 0.011286f
C150 VTAIL.n42 B 0.01195f
C151 VTAIL.n43 B 0.026677f
C152 VTAIL.n44 B 0.059004f
C153 VTAIL.n45 B 0.01195f
C154 VTAIL.n46 B 0.011286f
C155 VTAIL.n47 B 0.045392f
C156 VTAIL.n48 B 0.033043f
C157 VTAIL.n49 B 0.214234f
C158 VTAIL.n50 B 0.030231f
C159 VTAIL.n51 B 0.021003f
C160 VTAIL.n52 B 0.011286f
C161 VTAIL.n53 B 0.026677f
C162 VTAIL.n54 B 0.01195f
C163 VTAIL.n55 B 0.021003f
C164 VTAIL.n56 B 0.011286f
C165 VTAIL.n57 B 0.026677f
C166 VTAIL.n58 B 0.01195f
C167 VTAIL.n59 B 0.021003f
C168 VTAIL.n60 B 0.011286f
C169 VTAIL.n61 B 0.026677f
C170 VTAIL.n62 B 0.01195f
C171 VTAIL.n63 B 0.766789f
C172 VTAIL.n64 B 0.011286f
C173 VTAIL.t13 B 0.043547f
C174 VTAIL.n65 B 0.1042f
C175 VTAIL.n66 B 0.015759f
C176 VTAIL.n67 B 0.020007f
C177 VTAIL.n68 B 0.026677f
C178 VTAIL.n69 B 0.01195f
C179 VTAIL.n70 B 0.011286f
C180 VTAIL.n71 B 0.021003f
C181 VTAIL.n72 B 0.021003f
C182 VTAIL.n73 B 0.011286f
C183 VTAIL.n74 B 0.01195f
C184 VTAIL.n75 B 0.026677f
C185 VTAIL.n76 B 0.026677f
C186 VTAIL.n77 B 0.01195f
C187 VTAIL.n78 B 0.011286f
C188 VTAIL.n79 B 0.021003f
C189 VTAIL.n80 B 0.021003f
C190 VTAIL.n81 B 0.011286f
C191 VTAIL.n82 B 0.01195f
C192 VTAIL.n83 B 0.026677f
C193 VTAIL.n84 B 0.026677f
C194 VTAIL.n85 B 0.01195f
C195 VTAIL.n86 B 0.011286f
C196 VTAIL.n87 B 0.021003f
C197 VTAIL.n88 B 0.021003f
C198 VTAIL.n89 B 0.011286f
C199 VTAIL.n90 B 0.01195f
C200 VTAIL.n91 B 0.026677f
C201 VTAIL.n92 B 0.059004f
C202 VTAIL.n93 B 0.01195f
C203 VTAIL.n94 B 0.011286f
C204 VTAIL.n95 B 0.045392f
C205 VTAIL.n96 B 0.033043f
C206 VTAIL.n97 B 0.214234f
C207 VTAIL.t10 B 0.14556f
C208 VTAIL.t9 B 0.14556f
C209 VTAIL.n98 B 1.19665f
C210 VTAIL.n99 B 0.545829f
C211 VTAIL.n100 B 0.030231f
C212 VTAIL.n101 B 0.021003f
C213 VTAIL.n102 B 0.011286f
C214 VTAIL.n103 B 0.026677f
C215 VTAIL.n104 B 0.01195f
C216 VTAIL.n105 B 0.021003f
C217 VTAIL.n106 B 0.011286f
C218 VTAIL.n107 B 0.026677f
C219 VTAIL.n108 B 0.01195f
C220 VTAIL.n109 B 0.021003f
C221 VTAIL.n110 B 0.011286f
C222 VTAIL.n111 B 0.026677f
C223 VTAIL.n112 B 0.01195f
C224 VTAIL.n113 B 0.766789f
C225 VTAIL.n114 B 0.011286f
C226 VTAIL.t8 B 0.043547f
C227 VTAIL.n115 B 0.1042f
C228 VTAIL.n116 B 0.015759f
C229 VTAIL.n117 B 0.020007f
C230 VTAIL.n118 B 0.026677f
C231 VTAIL.n119 B 0.01195f
C232 VTAIL.n120 B 0.011286f
C233 VTAIL.n121 B 0.021003f
C234 VTAIL.n122 B 0.021003f
C235 VTAIL.n123 B 0.011286f
C236 VTAIL.n124 B 0.01195f
C237 VTAIL.n125 B 0.026677f
C238 VTAIL.n126 B 0.026677f
C239 VTAIL.n127 B 0.01195f
C240 VTAIL.n128 B 0.011286f
C241 VTAIL.n129 B 0.021003f
C242 VTAIL.n130 B 0.021003f
C243 VTAIL.n131 B 0.011286f
C244 VTAIL.n132 B 0.01195f
C245 VTAIL.n133 B 0.026677f
C246 VTAIL.n134 B 0.026677f
C247 VTAIL.n135 B 0.01195f
C248 VTAIL.n136 B 0.011286f
C249 VTAIL.n137 B 0.021003f
C250 VTAIL.n138 B 0.021003f
C251 VTAIL.n139 B 0.011286f
C252 VTAIL.n140 B 0.01195f
C253 VTAIL.n141 B 0.026677f
C254 VTAIL.n142 B 0.059004f
C255 VTAIL.n143 B 0.01195f
C256 VTAIL.n144 B 0.011286f
C257 VTAIL.n145 B 0.045392f
C258 VTAIL.n146 B 0.033043f
C259 VTAIL.n147 B 1.14569f
C260 VTAIL.n148 B 0.030231f
C261 VTAIL.n149 B 0.021003f
C262 VTAIL.n150 B 0.011286f
C263 VTAIL.n151 B 0.026677f
C264 VTAIL.n152 B 0.01195f
C265 VTAIL.n153 B 0.021003f
C266 VTAIL.n154 B 0.011286f
C267 VTAIL.n155 B 0.026677f
C268 VTAIL.n156 B 0.01195f
C269 VTAIL.n157 B 0.021003f
C270 VTAIL.n158 B 0.011286f
C271 VTAIL.n159 B 0.026677f
C272 VTAIL.n160 B 0.01195f
C273 VTAIL.n161 B 0.766789f
C274 VTAIL.n162 B 0.011286f
C275 VTAIL.t3 B 0.043547f
C276 VTAIL.n163 B 0.1042f
C277 VTAIL.n164 B 0.015759f
C278 VTAIL.n165 B 0.020007f
C279 VTAIL.n166 B 0.026677f
C280 VTAIL.n167 B 0.01195f
C281 VTAIL.n168 B 0.011286f
C282 VTAIL.n169 B 0.021003f
C283 VTAIL.n170 B 0.021003f
C284 VTAIL.n171 B 0.011286f
C285 VTAIL.n172 B 0.01195f
C286 VTAIL.n173 B 0.026677f
C287 VTAIL.n174 B 0.026677f
C288 VTAIL.n175 B 0.01195f
C289 VTAIL.n176 B 0.011286f
C290 VTAIL.n177 B 0.021003f
C291 VTAIL.n178 B 0.021003f
C292 VTAIL.n179 B 0.011286f
C293 VTAIL.n180 B 0.01195f
C294 VTAIL.n181 B 0.026677f
C295 VTAIL.n182 B 0.026677f
C296 VTAIL.n183 B 0.01195f
C297 VTAIL.n184 B 0.011286f
C298 VTAIL.n185 B 0.021003f
C299 VTAIL.n186 B 0.021003f
C300 VTAIL.n187 B 0.011286f
C301 VTAIL.n188 B 0.01195f
C302 VTAIL.n189 B 0.026677f
C303 VTAIL.n190 B 0.059004f
C304 VTAIL.n191 B 0.01195f
C305 VTAIL.n192 B 0.011286f
C306 VTAIL.n193 B 0.045392f
C307 VTAIL.n194 B 0.033043f
C308 VTAIL.n195 B 1.14569f
C309 VTAIL.t1 B 0.14556f
C310 VTAIL.t7 B 0.14556f
C311 VTAIL.n196 B 1.19666f
C312 VTAIL.n197 B 0.545821f
C313 VTAIL.n198 B 0.030231f
C314 VTAIL.n199 B 0.021003f
C315 VTAIL.n200 B 0.011286f
C316 VTAIL.n201 B 0.026677f
C317 VTAIL.n202 B 0.01195f
C318 VTAIL.n203 B 0.021003f
C319 VTAIL.n204 B 0.011286f
C320 VTAIL.n205 B 0.026677f
C321 VTAIL.n206 B 0.01195f
C322 VTAIL.n207 B 0.021003f
C323 VTAIL.n208 B 0.011286f
C324 VTAIL.n209 B 0.026677f
C325 VTAIL.n210 B 0.01195f
C326 VTAIL.n211 B 0.766789f
C327 VTAIL.n212 B 0.011286f
C328 VTAIL.t6 B 0.043547f
C329 VTAIL.n213 B 0.1042f
C330 VTAIL.n214 B 0.015759f
C331 VTAIL.n215 B 0.020007f
C332 VTAIL.n216 B 0.026677f
C333 VTAIL.n217 B 0.01195f
C334 VTAIL.n218 B 0.011286f
C335 VTAIL.n219 B 0.021003f
C336 VTAIL.n220 B 0.021003f
C337 VTAIL.n221 B 0.011286f
C338 VTAIL.n222 B 0.01195f
C339 VTAIL.n223 B 0.026677f
C340 VTAIL.n224 B 0.026677f
C341 VTAIL.n225 B 0.01195f
C342 VTAIL.n226 B 0.011286f
C343 VTAIL.n227 B 0.021003f
C344 VTAIL.n228 B 0.021003f
C345 VTAIL.n229 B 0.011286f
C346 VTAIL.n230 B 0.01195f
C347 VTAIL.n231 B 0.026677f
C348 VTAIL.n232 B 0.026677f
C349 VTAIL.n233 B 0.01195f
C350 VTAIL.n234 B 0.011286f
C351 VTAIL.n235 B 0.021003f
C352 VTAIL.n236 B 0.021003f
C353 VTAIL.n237 B 0.011286f
C354 VTAIL.n238 B 0.01195f
C355 VTAIL.n239 B 0.026677f
C356 VTAIL.n240 B 0.059004f
C357 VTAIL.n241 B 0.01195f
C358 VTAIL.n242 B 0.011286f
C359 VTAIL.n243 B 0.045392f
C360 VTAIL.n244 B 0.033043f
C361 VTAIL.n245 B 0.214234f
C362 VTAIL.n246 B 0.030231f
C363 VTAIL.n247 B 0.021003f
C364 VTAIL.n248 B 0.011286f
C365 VTAIL.n249 B 0.026677f
C366 VTAIL.n250 B 0.01195f
C367 VTAIL.n251 B 0.021003f
C368 VTAIL.n252 B 0.011286f
C369 VTAIL.n253 B 0.026677f
C370 VTAIL.n254 B 0.01195f
C371 VTAIL.n255 B 0.021003f
C372 VTAIL.n256 B 0.011286f
C373 VTAIL.n257 B 0.026677f
C374 VTAIL.n258 B 0.01195f
C375 VTAIL.n259 B 0.766789f
C376 VTAIL.n260 B 0.011286f
C377 VTAIL.t11 B 0.043547f
C378 VTAIL.n261 B 0.1042f
C379 VTAIL.n262 B 0.015759f
C380 VTAIL.n263 B 0.020007f
C381 VTAIL.n264 B 0.026677f
C382 VTAIL.n265 B 0.01195f
C383 VTAIL.n266 B 0.011286f
C384 VTAIL.n267 B 0.021003f
C385 VTAIL.n268 B 0.021003f
C386 VTAIL.n269 B 0.011286f
C387 VTAIL.n270 B 0.01195f
C388 VTAIL.n271 B 0.026677f
C389 VTAIL.n272 B 0.026677f
C390 VTAIL.n273 B 0.01195f
C391 VTAIL.n274 B 0.011286f
C392 VTAIL.n275 B 0.021003f
C393 VTAIL.n276 B 0.021003f
C394 VTAIL.n277 B 0.011286f
C395 VTAIL.n278 B 0.01195f
C396 VTAIL.n279 B 0.026677f
C397 VTAIL.n280 B 0.026677f
C398 VTAIL.n281 B 0.01195f
C399 VTAIL.n282 B 0.011286f
C400 VTAIL.n283 B 0.021003f
C401 VTAIL.n284 B 0.021003f
C402 VTAIL.n285 B 0.011286f
C403 VTAIL.n286 B 0.01195f
C404 VTAIL.n287 B 0.026677f
C405 VTAIL.n288 B 0.059004f
C406 VTAIL.n289 B 0.01195f
C407 VTAIL.n290 B 0.011286f
C408 VTAIL.n291 B 0.045392f
C409 VTAIL.n292 B 0.033043f
C410 VTAIL.n293 B 0.214234f
C411 VTAIL.t12 B 0.14556f
C412 VTAIL.t15 B 0.14556f
C413 VTAIL.n294 B 1.19666f
C414 VTAIL.n295 B 0.545821f
C415 VTAIL.n296 B 0.030231f
C416 VTAIL.n297 B 0.021003f
C417 VTAIL.n298 B 0.011286f
C418 VTAIL.n299 B 0.026677f
C419 VTAIL.n300 B 0.01195f
C420 VTAIL.n301 B 0.021003f
C421 VTAIL.n302 B 0.011286f
C422 VTAIL.n303 B 0.026677f
C423 VTAIL.n304 B 0.01195f
C424 VTAIL.n305 B 0.021003f
C425 VTAIL.n306 B 0.011286f
C426 VTAIL.n307 B 0.026677f
C427 VTAIL.n308 B 0.01195f
C428 VTAIL.n309 B 0.766789f
C429 VTAIL.n310 B 0.011286f
C430 VTAIL.t14 B 0.043547f
C431 VTAIL.n311 B 0.1042f
C432 VTAIL.n312 B 0.015759f
C433 VTAIL.n313 B 0.020007f
C434 VTAIL.n314 B 0.026677f
C435 VTAIL.n315 B 0.01195f
C436 VTAIL.n316 B 0.011286f
C437 VTAIL.n317 B 0.021003f
C438 VTAIL.n318 B 0.021003f
C439 VTAIL.n319 B 0.011286f
C440 VTAIL.n320 B 0.01195f
C441 VTAIL.n321 B 0.026677f
C442 VTAIL.n322 B 0.026677f
C443 VTAIL.n323 B 0.01195f
C444 VTAIL.n324 B 0.011286f
C445 VTAIL.n325 B 0.021003f
C446 VTAIL.n326 B 0.021003f
C447 VTAIL.n327 B 0.011286f
C448 VTAIL.n328 B 0.01195f
C449 VTAIL.n329 B 0.026677f
C450 VTAIL.n330 B 0.026677f
C451 VTAIL.n331 B 0.01195f
C452 VTAIL.n332 B 0.011286f
C453 VTAIL.n333 B 0.021003f
C454 VTAIL.n334 B 0.021003f
C455 VTAIL.n335 B 0.011286f
C456 VTAIL.n336 B 0.01195f
C457 VTAIL.n337 B 0.026677f
C458 VTAIL.n338 B 0.059004f
C459 VTAIL.n339 B 0.01195f
C460 VTAIL.n340 B 0.011286f
C461 VTAIL.n341 B 0.045392f
C462 VTAIL.n342 B 0.033043f
C463 VTAIL.n343 B 1.14569f
C464 VTAIL.n344 B 0.030231f
C465 VTAIL.n345 B 0.021003f
C466 VTAIL.n346 B 0.011286f
C467 VTAIL.n347 B 0.026677f
C468 VTAIL.n348 B 0.01195f
C469 VTAIL.n349 B 0.021003f
C470 VTAIL.n350 B 0.011286f
C471 VTAIL.n351 B 0.026677f
C472 VTAIL.n352 B 0.01195f
C473 VTAIL.n353 B 0.021003f
C474 VTAIL.n354 B 0.011286f
C475 VTAIL.n355 B 0.026677f
C476 VTAIL.n356 B 0.01195f
C477 VTAIL.n357 B 0.766789f
C478 VTAIL.n358 B 0.011286f
C479 VTAIL.t0 B 0.043547f
C480 VTAIL.n359 B 0.1042f
C481 VTAIL.n360 B 0.015759f
C482 VTAIL.n361 B 0.020007f
C483 VTAIL.n362 B 0.026677f
C484 VTAIL.n363 B 0.01195f
C485 VTAIL.n364 B 0.011286f
C486 VTAIL.n365 B 0.021003f
C487 VTAIL.n366 B 0.021003f
C488 VTAIL.n367 B 0.011286f
C489 VTAIL.n368 B 0.01195f
C490 VTAIL.n369 B 0.026677f
C491 VTAIL.n370 B 0.026677f
C492 VTAIL.n371 B 0.01195f
C493 VTAIL.n372 B 0.011286f
C494 VTAIL.n373 B 0.021003f
C495 VTAIL.n374 B 0.021003f
C496 VTAIL.n375 B 0.011286f
C497 VTAIL.n376 B 0.01195f
C498 VTAIL.n377 B 0.026677f
C499 VTAIL.n378 B 0.026677f
C500 VTAIL.n379 B 0.01195f
C501 VTAIL.n380 B 0.011286f
C502 VTAIL.n381 B 0.021003f
C503 VTAIL.n382 B 0.021003f
C504 VTAIL.n383 B 0.011286f
C505 VTAIL.n384 B 0.01195f
C506 VTAIL.n385 B 0.026677f
C507 VTAIL.n386 B 0.059004f
C508 VTAIL.n387 B 0.01195f
C509 VTAIL.n388 B 0.011286f
C510 VTAIL.n389 B 0.045392f
C511 VTAIL.n390 B 0.033043f
C512 VTAIL.n391 B 1.14175f
C513 VP.n0 B 0.031782f
C514 VP.t6 B 1.4363f
C515 VP.n1 B 0.02749f
C516 VP.n2 B 0.024107f
C517 VP.t1 B 1.4363f
C518 VP.n3 B 0.519863f
C519 VP.n4 B 0.024107f
C520 VP.n5 B 0.047911f
C521 VP.n6 B 0.024107f
C522 VP.t5 B 1.4363f
C523 VP.n7 B 0.041722f
C524 VP.n8 B 0.024107f
C525 VP.t7 B 1.4363f
C526 VP.n9 B 0.602955f
C527 VP.n10 B 0.031782f
C528 VP.t0 B 1.4363f
C529 VP.n11 B 0.02749f
C530 VP.n12 B 0.024107f
C531 VP.t2 B 1.4363f
C532 VP.n13 B 0.519863f
C533 VP.n14 B 0.024107f
C534 VP.n15 B 0.047911f
C535 VP.t4 B 1.63144f
C536 VP.n16 B 0.566315f
C537 VP.t3 B 1.4363f
C538 VP.n17 B 0.596918f
C539 VP.n18 B 0.0416f
C540 VP.n19 B 0.230983f
C541 VP.n20 B 0.024107f
C542 VP.n21 B 0.024107f
C543 VP.n22 B 0.019488f
C544 VP.n23 B 0.047911f
C545 VP.n24 B 0.0416f
C546 VP.n25 B 0.024107f
C547 VP.n26 B 0.024107f
C548 VP.n27 B 0.026073f
C549 VP.n28 B 0.044928f
C550 VP.n29 B 0.041722f
C551 VP.n30 B 0.024107f
C552 VP.n31 B 0.024107f
C553 VP.n32 B 0.024107f
C554 VP.n33 B 0.046099f
C555 VP.n34 B 0.034946f
C556 VP.n35 B 0.602955f
C557 VP.n36 B 1.26511f
C558 VP.n37 B 1.28311f
C559 VP.n38 B 0.031782f
C560 VP.n39 B 0.034946f
C561 VP.n40 B 0.046099f
C562 VP.n41 B 0.02749f
C563 VP.n42 B 0.024107f
C564 VP.n43 B 0.024107f
C565 VP.n44 B 0.024107f
C566 VP.n45 B 0.044928f
C567 VP.n46 B 0.026073f
C568 VP.n47 B 0.519863f
C569 VP.n48 B 0.0416f
C570 VP.n49 B 0.024107f
C571 VP.n50 B 0.024107f
C572 VP.n51 B 0.024107f
C573 VP.n52 B 0.019488f
C574 VP.n53 B 0.047911f
C575 VP.n54 B 0.0416f
C576 VP.n55 B 0.024107f
C577 VP.n56 B 0.024107f
C578 VP.n57 B 0.026073f
C579 VP.n58 B 0.044928f
C580 VP.n59 B 0.041722f
C581 VP.n60 B 0.024107f
C582 VP.n61 B 0.024107f
C583 VP.n62 B 0.024107f
C584 VP.n63 B 0.046099f
C585 VP.n64 B 0.034946f
C586 VP.n65 B 0.602955f
C587 VP.n66 B 0.036371f
.ends

