* NGSPICE file created from diff_pair_sample_1604.ext - technology: sky130A

.subckt diff_pair_sample_1604 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=7.5348 ps=39.42 w=19.32 l=0.9
X1 VTAIL.t9 VP.t1 VDD1.t8 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X2 VTAIL.t10 VP.t2 VDD1.t7 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X3 VDD1.t6 VP.t3 VTAIL.t15 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X4 VDD1.t5 VP.t4 VTAIL.t17 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=3.1878 ps=19.65 w=19.32 l=0.9
X5 VDD1.t4 VP.t5 VTAIL.t8 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=3.1878 ps=19.65 w=19.32 l=0.9
X6 VDD1.t3 VP.t6 VTAIL.t16 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X7 B.t11 B.t9 B.t10 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=0 ps=0 w=19.32 l=0.9
X8 VDD1.t2 VP.t7 VTAIL.t14 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=7.5348 ps=39.42 w=19.32 l=0.9
X9 VDD2.t9 VN.t0 VTAIL.t5 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=7.5348 ps=39.42 w=19.32 l=0.9
X10 VDD2.t8 VN.t1 VTAIL.t2 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X11 VDD2.t7 VN.t2 VTAIL.t18 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=3.1878 ps=19.65 w=19.32 l=0.9
X12 VTAIL.t13 VP.t8 VDD1.t1 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X13 VTAIL.t4 VN.t3 VDD2.t6 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X14 B.t8 B.t6 B.t7 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=0 ps=0 w=19.32 l=0.9
X15 VTAIL.t12 VP.t9 VDD1.t0 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X16 VDD2.t5 VN.t4 VTAIL.t0 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=3.1878 ps=19.65 w=19.32 l=0.9
X17 VDD2.t4 VN.t5 VTAIL.t19 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X18 VTAIL.t3 VN.t6 VDD2.t3 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X19 VTAIL.t7 VN.t7 VDD2.t2 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X20 VTAIL.t6 VN.t8 VDD2.t1 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=3.1878 ps=19.65 w=19.32 l=0.9
X21 B.t5 B.t3 B.t4 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=0 ps=0 w=19.32 l=0.9
X22 B.t2 B.t0 B.t1 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=7.5348 pd=39.42 as=0 ps=0 w=19.32 l=0.9
X23 VDD2.t0 VN.t9 VTAIL.t1 w_n2446_n4832# sky130_fd_pr__pfet_01v8 ad=3.1878 pd=19.65 as=7.5348 ps=39.42 w=19.32 l=0.9
R0 VP.n10 VP.t5 576.934
R1 VP.n5 VP.t4 560.995
R2 VP.n41 VP.t0 560.995
R3 VP.n23 VP.t7 560.995
R4 VP.n34 VP.t3 517.347
R5 VP.n29 VP.t1 517.347
R6 VP.n1 VP.t2 517.347
R7 VP.n16 VP.t6 517.347
R8 VP.n7 VP.t9 517.347
R9 VP.n11 VP.t8 517.347
R10 VP.n42 VP.n41 161.3
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n9 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n8 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n40 VP.n0 161.3
R20 VP.n39 VP.n38 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n25 VP.n5 161.3
R29 VP.n28 VP.n27 55.593
R30 VP.n40 VP.n39 55.593
R31 VP.n22 VP.n21 55.593
R32 VP.n30 VP.n3 51.7179
R33 VP.n36 VP.n35 51.7179
R34 VP.n18 VP.n17 51.7179
R35 VP.n12 VP.n9 51.7179
R36 VP.n25 VP.n24 49.3906
R37 VP.n13 VP.n10 43.7549
R38 VP.n11 VP.n10 43.7503
R39 VP.n34 VP.n3 29.4362
R40 VP.n35 VP.n34 29.4362
R41 VP.n17 VP.n16 29.4362
R42 VP.n16 VP.n9 29.4362
R43 VP.n29 VP.n28 13.2801
R44 VP.n39 VP.n1 13.2801
R45 VP.n21 VP.n7 13.2801
R46 VP.n30 VP.n29 11.3127
R47 VP.n36 VP.n1 11.3127
R48 VP.n18 VP.n7 11.3127
R49 VP.n12 VP.n11 11.3127
R50 VP.n27 VP.n5 1.46111
R51 VP.n41 VP.n40 1.46111
R52 VP.n23 VP.n22 1.46111
R53 VP.n14 VP.n13 0.189894
R54 VP.n15 VP.n14 0.189894
R55 VP.n15 VP.n8 0.189894
R56 VP.n19 VP.n8 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n37 VP.n2 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n38 VP.n0 0.189894
R69 VP.n42 VP.n0 0.189894
R70 VP VP.n42 0.0516364
R71 VTAIL.n11 VTAIL.t5 53.2476
R72 VTAIL.n17 VTAIL.t1 53.2473
R73 VTAIL.n2 VTAIL.t11 53.2473
R74 VTAIL.n16 VTAIL.t14 53.2473
R75 VTAIL.n15 VTAIL.n14 51.5651
R76 VTAIL.n13 VTAIL.n12 51.5651
R77 VTAIL.n10 VTAIL.n9 51.5651
R78 VTAIL.n8 VTAIL.n7 51.5651
R79 VTAIL.n19 VTAIL.n18 51.5651
R80 VTAIL.n1 VTAIL.n0 51.5651
R81 VTAIL.n4 VTAIL.n3 51.5651
R82 VTAIL.n6 VTAIL.n5 51.5651
R83 VTAIL.n8 VTAIL.n6 31.1427
R84 VTAIL.n17 VTAIL.n16 30.0824
R85 VTAIL.n18 VTAIL.t19 1.68295
R86 VTAIL.n18 VTAIL.t3 1.68295
R87 VTAIL.n0 VTAIL.t18 1.68295
R88 VTAIL.n0 VTAIL.t4 1.68295
R89 VTAIL.n3 VTAIL.t15 1.68295
R90 VTAIL.n3 VTAIL.t10 1.68295
R91 VTAIL.n5 VTAIL.t17 1.68295
R92 VTAIL.n5 VTAIL.t9 1.68295
R93 VTAIL.n14 VTAIL.t16 1.68295
R94 VTAIL.n14 VTAIL.t12 1.68295
R95 VTAIL.n12 VTAIL.t8 1.68295
R96 VTAIL.n12 VTAIL.t13 1.68295
R97 VTAIL.n9 VTAIL.t2 1.68295
R98 VTAIL.n9 VTAIL.t7 1.68295
R99 VTAIL.n7 VTAIL.t0 1.68295
R100 VTAIL.n7 VTAIL.t6 1.68295
R101 VTAIL.n10 VTAIL.n8 1.06084
R102 VTAIL.n11 VTAIL.n10 1.06084
R103 VTAIL.n15 VTAIL.n13 1.06084
R104 VTAIL.n16 VTAIL.n15 1.06084
R105 VTAIL.n6 VTAIL.n4 1.06084
R106 VTAIL.n4 VTAIL.n2 1.06084
R107 VTAIL.n19 VTAIL.n17 1.06084
R108 VTAIL.n13 VTAIL.n11 1.0005
R109 VTAIL.n2 VTAIL.n1 1.0005
R110 VTAIL VTAIL.n1 0.853948
R111 VTAIL VTAIL.n19 0.207397
R112 VDD1.n1 VDD1.t4 70.9867
R113 VDD1.n3 VDD1.t5 70.9864
R114 VDD1.n5 VDD1.n4 68.9838
R115 VDD1.n1 VDD1.n0 68.2439
R116 VDD1.n3 VDD1.n2 68.2438
R117 VDD1.n7 VDD1.n6 68.2437
R118 VDD1.n7 VDD1.n5 46.5203
R119 VDD1.n6 VDD1.t0 1.68295
R120 VDD1.n6 VDD1.t2 1.68295
R121 VDD1.n0 VDD1.t1 1.68295
R122 VDD1.n0 VDD1.t3 1.68295
R123 VDD1.n4 VDD1.t7 1.68295
R124 VDD1.n4 VDD1.t9 1.68295
R125 VDD1.n2 VDD1.t8 1.68295
R126 VDD1.n2 VDD1.t6 1.68295
R127 VDD1 VDD1.n7 0.737569
R128 VDD1 VDD1.n1 0.323776
R129 VDD1.n5 VDD1.n3 0.21024
R130 B.n153 B.t0 719.543
R131 B.n159 B.t6 719.543
R132 B.n50 B.t9 719.543
R133 B.n57 B.t3 719.543
R134 B.n549 B.n548 585
R135 B.n550 B.n89 585
R136 B.n552 B.n551 585
R137 B.n553 B.n88 585
R138 B.n555 B.n554 585
R139 B.n556 B.n87 585
R140 B.n558 B.n557 585
R141 B.n559 B.n86 585
R142 B.n561 B.n560 585
R143 B.n562 B.n85 585
R144 B.n564 B.n563 585
R145 B.n565 B.n84 585
R146 B.n567 B.n566 585
R147 B.n568 B.n83 585
R148 B.n570 B.n569 585
R149 B.n571 B.n82 585
R150 B.n573 B.n572 585
R151 B.n574 B.n81 585
R152 B.n576 B.n575 585
R153 B.n577 B.n80 585
R154 B.n579 B.n578 585
R155 B.n580 B.n79 585
R156 B.n582 B.n581 585
R157 B.n583 B.n78 585
R158 B.n585 B.n584 585
R159 B.n586 B.n77 585
R160 B.n588 B.n587 585
R161 B.n589 B.n76 585
R162 B.n591 B.n590 585
R163 B.n592 B.n75 585
R164 B.n594 B.n593 585
R165 B.n595 B.n74 585
R166 B.n597 B.n596 585
R167 B.n598 B.n73 585
R168 B.n600 B.n599 585
R169 B.n601 B.n72 585
R170 B.n603 B.n602 585
R171 B.n604 B.n71 585
R172 B.n606 B.n605 585
R173 B.n607 B.n70 585
R174 B.n609 B.n608 585
R175 B.n610 B.n69 585
R176 B.n612 B.n611 585
R177 B.n613 B.n68 585
R178 B.n615 B.n614 585
R179 B.n616 B.n67 585
R180 B.n618 B.n617 585
R181 B.n619 B.n66 585
R182 B.n621 B.n620 585
R183 B.n622 B.n65 585
R184 B.n624 B.n623 585
R185 B.n625 B.n64 585
R186 B.n627 B.n626 585
R187 B.n628 B.n63 585
R188 B.n630 B.n629 585
R189 B.n631 B.n62 585
R190 B.n633 B.n632 585
R191 B.n634 B.n61 585
R192 B.n636 B.n635 585
R193 B.n637 B.n60 585
R194 B.n639 B.n638 585
R195 B.n640 B.n59 585
R196 B.n642 B.n641 585
R197 B.n644 B.n56 585
R198 B.n646 B.n645 585
R199 B.n647 B.n55 585
R200 B.n649 B.n648 585
R201 B.n650 B.n54 585
R202 B.n652 B.n651 585
R203 B.n653 B.n53 585
R204 B.n655 B.n654 585
R205 B.n656 B.n49 585
R206 B.n658 B.n657 585
R207 B.n659 B.n48 585
R208 B.n661 B.n660 585
R209 B.n662 B.n47 585
R210 B.n664 B.n663 585
R211 B.n665 B.n46 585
R212 B.n667 B.n666 585
R213 B.n668 B.n45 585
R214 B.n670 B.n669 585
R215 B.n671 B.n44 585
R216 B.n673 B.n672 585
R217 B.n674 B.n43 585
R218 B.n676 B.n675 585
R219 B.n677 B.n42 585
R220 B.n679 B.n678 585
R221 B.n680 B.n41 585
R222 B.n682 B.n681 585
R223 B.n683 B.n40 585
R224 B.n685 B.n684 585
R225 B.n686 B.n39 585
R226 B.n688 B.n687 585
R227 B.n689 B.n38 585
R228 B.n691 B.n690 585
R229 B.n692 B.n37 585
R230 B.n694 B.n693 585
R231 B.n695 B.n36 585
R232 B.n697 B.n696 585
R233 B.n698 B.n35 585
R234 B.n700 B.n699 585
R235 B.n701 B.n34 585
R236 B.n703 B.n702 585
R237 B.n704 B.n33 585
R238 B.n706 B.n705 585
R239 B.n707 B.n32 585
R240 B.n709 B.n708 585
R241 B.n710 B.n31 585
R242 B.n712 B.n711 585
R243 B.n713 B.n30 585
R244 B.n715 B.n714 585
R245 B.n716 B.n29 585
R246 B.n718 B.n717 585
R247 B.n719 B.n28 585
R248 B.n721 B.n720 585
R249 B.n722 B.n27 585
R250 B.n724 B.n723 585
R251 B.n725 B.n26 585
R252 B.n727 B.n726 585
R253 B.n728 B.n25 585
R254 B.n730 B.n729 585
R255 B.n731 B.n24 585
R256 B.n733 B.n732 585
R257 B.n734 B.n23 585
R258 B.n736 B.n735 585
R259 B.n737 B.n22 585
R260 B.n739 B.n738 585
R261 B.n740 B.n21 585
R262 B.n742 B.n741 585
R263 B.n743 B.n20 585
R264 B.n745 B.n744 585
R265 B.n746 B.n19 585
R266 B.n748 B.n747 585
R267 B.n749 B.n18 585
R268 B.n751 B.n750 585
R269 B.n752 B.n17 585
R270 B.n547 B.n90 585
R271 B.n546 B.n545 585
R272 B.n544 B.n91 585
R273 B.n543 B.n542 585
R274 B.n541 B.n92 585
R275 B.n540 B.n539 585
R276 B.n538 B.n93 585
R277 B.n537 B.n536 585
R278 B.n535 B.n94 585
R279 B.n534 B.n533 585
R280 B.n532 B.n95 585
R281 B.n531 B.n530 585
R282 B.n529 B.n96 585
R283 B.n528 B.n527 585
R284 B.n526 B.n97 585
R285 B.n525 B.n524 585
R286 B.n523 B.n98 585
R287 B.n522 B.n521 585
R288 B.n520 B.n99 585
R289 B.n519 B.n518 585
R290 B.n517 B.n100 585
R291 B.n516 B.n515 585
R292 B.n514 B.n101 585
R293 B.n513 B.n512 585
R294 B.n511 B.n102 585
R295 B.n510 B.n509 585
R296 B.n508 B.n103 585
R297 B.n507 B.n506 585
R298 B.n505 B.n104 585
R299 B.n504 B.n503 585
R300 B.n502 B.n105 585
R301 B.n501 B.n500 585
R302 B.n499 B.n106 585
R303 B.n498 B.n497 585
R304 B.n496 B.n107 585
R305 B.n495 B.n494 585
R306 B.n493 B.n108 585
R307 B.n492 B.n491 585
R308 B.n490 B.n109 585
R309 B.n489 B.n488 585
R310 B.n487 B.n110 585
R311 B.n486 B.n485 585
R312 B.n484 B.n111 585
R313 B.n483 B.n482 585
R314 B.n481 B.n112 585
R315 B.n480 B.n479 585
R316 B.n478 B.n113 585
R317 B.n477 B.n476 585
R318 B.n475 B.n114 585
R319 B.n474 B.n473 585
R320 B.n472 B.n115 585
R321 B.n471 B.n470 585
R322 B.n469 B.n116 585
R323 B.n468 B.n467 585
R324 B.n466 B.n117 585
R325 B.n465 B.n464 585
R326 B.n463 B.n118 585
R327 B.n462 B.n461 585
R328 B.n460 B.n119 585
R329 B.n459 B.n458 585
R330 B.n457 B.n120 585
R331 B.n252 B.n251 585
R332 B.n253 B.n192 585
R333 B.n255 B.n254 585
R334 B.n256 B.n191 585
R335 B.n258 B.n257 585
R336 B.n259 B.n190 585
R337 B.n261 B.n260 585
R338 B.n262 B.n189 585
R339 B.n264 B.n263 585
R340 B.n265 B.n188 585
R341 B.n267 B.n266 585
R342 B.n268 B.n187 585
R343 B.n270 B.n269 585
R344 B.n271 B.n186 585
R345 B.n273 B.n272 585
R346 B.n274 B.n185 585
R347 B.n276 B.n275 585
R348 B.n277 B.n184 585
R349 B.n279 B.n278 585
R350 B.n280 B.n183 585
R351 B.n282 B.n281 585
R352 B.n283 B.n182 585
R353 B.n285 B.n284 585
R354 B.n286 B.n181 585
R355 B.n288 B.n287 585
R356 B.n289 B.n180 585
R357 B.n291 B.n290 585
R358 B.n292 B.n179 585
R359 B.n294 B.n293 585
R360 B.n295 B.n178 585
R361 B.n297 B.n296 585
R362 B.n298 B.n177 585
R363 B.n300 B.n299 585
R364 B.n301 B.n176 585
R365 B.n303 B.n302 585
R366 B.n304 B.n175 585
R367 B.n306 B.n305 585
R368 B.n307 B.n174 585
R369 B.n309 B.n308 585
R370 B.n310 B.n173 585
R371 B.n312 B.n311 585
R372 B.n313 B.n172 585
R373 B.n315 B.n314 585
R374 B.n316 B.n171 585
R375 B.n318 B.n317 585
R376 B.n319 B.n170 585
R377 B.n321 B.n320 585
R378 B.n322 B.n169 585
R379 B.n324 B.n323 585
R380 B.n325 B.n168 585
R381 B.n327 B.n326 585
R382 B.n328 B.n167 585
R383 B.n330 B.n329 585
R384 B.n331 B.n166 585
R385 B.n333 B.n332 585
R386 B.n334 B.n165 585
R387 B.n336 B.n335 585
R388 B.n337 B.n164 585
R389 B.n339 B.n338 585
R390 B.n340 B.n163 585
R391 B.n342 B.n341 585
R392 B.n343 B.n162 585
R393 B.n345 B.n344 585
R394 B.n347 B.n346 585
R395 B.n348 B.n158 585
R396 B.n350 B.n349 585
R397 B.n351 B.n157 585
R398 B.n353 B.n352 585
R399 B.n354 B.n156 585
R400 B.n356 B.n355 585
R401 B.n357 B.n155 585
R402 B.n359 B.n358 585
R403 B.n360 B.n152 585
R404 B.n363 B.n362 585
R405 B.n364 B.n151 585
R406 B.n366 B.n365 585
R407 B.n367 B.n150 585
R408 B.n369 B.n368 585
R409 B.n370 B.n149 585
R410 B.n372 B.n371 585
R411 B.n373 B.n148 585
R412 B.n375 B.n374 585
R413 B.n376 B.n147 585
R414 B.n378 B.n377 585
R415 B.n379 B.n146 585
R416 B.n381 B.n380 585
R417 B.n382 B.n145 585
R418 B.n384 B.n383 585
R419 B.n385 B.n144 585
R420 B.n387 B.n386 585
R421 B.n388 B.n143 585
R422 B.n390 B.n389 585
R423 B.n391 B.n142 585
R424 B.n393 B.n392 585
R425 B.n394 B.n141 585
R426 B.n396 B.n395 585
R427 B.n397 B.n140 585
R428 B.n399 B.n398 585
R429 B.n400 B.n139 585
R430 B.n402 B.n401 585
R431 B.n403 B.n138 585
R432 B.n405 B.n404 585
R433 B.n406 B.n137 585
R434 B.n408 B.n407 585
R435 B.n409 B.n136 585
R436 B.n411 B.n410 585
R437 B.n412 B.n135 585
R438 B.n414 B.n413 585
R439 B.n415 B.n134 585
R440 B.n417 B.n416 585
R441 B.n418 B.n133 585
R442 B.n420 B.n419 585
R443 B.n421 B.n132 585
R444 B.n423 B.n422 585
R445 B.n424 B.n131 585
R446 B.n426 B.n425 585
R447 B.n427 B.n130 585
R448 B.n429 B.n428 585
R449 B.n430 B.n129 585
R450 B.n432 B.n431 585
R451 B.n433 B.n128 585
R452 B.n435 B.n434 585
R453 B.n436 B.n127 585
R454 B.n438 B.n437 585
R455 B.n439 B.n126 585
R456 B.n441 B.n440 585
R457 B.n442 B.n125 585
R458 B.n444 B.n443 585
R459 B.n445 B.n124 585
R460 B.n447 B.n446 585
R461 B.n448 B.n123 585
R462 B.n450 B.n449 585
R463 B.n451 B.n122 585
R464 B.n453 B.n452 585
R465 B.n454 B.n121 585
R466 B.n456 B.n455 585
R467 B.n250 B.n193 585
R468 B.n249 B.n248 585
R469 B.n247 B.n194 585
R470 B.n246 B.n245 585
R471 B.n244 B.n195 585
R472 B.n243 B.n242 585
R473 B.n241 B.n196 585
R474 B.n240 B.n239 585
R475 B.n238 B.n197 585
R476 B.n237 B.n236 585
R477 B.n235 B.n198 585
R478 B.n234 B.n233 585
R479 B.n232 B.n199 585
R480 B.n231 B.n230 585
R481 B.n229 B.n200 585
R482 B.n228 B.n227 585
R483 B.n226 B.n201 585
R484 B.n225 B.n224 585
R485 B.n223 B.n202 585
R486 B.n222 B.n221 585
R487 B.n220 B.n203 585
R488 B.n219 B.n218 585
R489 B.n217 B.n204 585
R490 B.n216 B.n215 585
R491 B.n214 B.n205 585
R492 B.n213 B.n212 585
R493 B.n211 B.n206 585
R494 B.n210 B.n209 585
R495 B.n208 B.n207 585
R496 B.n2 B.n0 585
R497 B.n797 B.n1 585
R498 B.n796 B.n795 585
R499 B.n794 B.n3 585
R500 B.n793 B.n792 585
R501 B.n791 B.n4 585
R502 B.n790 B.n789 585
R503 B.n788 B.n5 585
R504 B.n787 B.n786 585
R505 B.n785 B.n6 585
R506 B.n784 B.n783 585
R507 B.n782 B.n7 585
R508 B.n781 B.n780 585
R509 B.n779 B.n8 585
R510 B.n778 B.n777 585
R511 B.n776 B.n9 585
R512 B.n775 B.n774 585
R513 B.n773 B.n10 585
R514 B.n772 B.n771 585
R515 B.n770 B.n11 585
R516 B.n769 B.n768 585
R517 B.n767 B.n12 585
R518 B.n766 B.n765 585
R519 B.n764 B.n13 585
R520 B.n763 B.n762 585
R521 B.n761 B.n14 585
R522 B.n760 B.n759 585
R523 B.n758 B.n15 585
R524 B.n757 B.n756 585
R525 B.n755 B.n16 585
R526 B.n754 B.n753 585
R527 B.n799 B.n798 585
R528 B.n251 B.n250 458.866
R529 B.n754 B.n17 458.866
R530 B.n455 B.n120 458.866
R531 B.n549 B.n90 458.866
R532 B.n250 B.n249 163.367
R533 B.n249 B.n194 163.367
R534 B.n245 B.n194 163.367
R535 B.n245 B.n244 163.367
R536 B.n244 B.n243 163.367
R537 B.n243 B.n196 163.367
R538 B.n239 B.n196 163.367
R539 B.n239 B.n238 163.367
R540 B.n238 B.n237 163.367
R541 B.n237 B.n198 163.367
R542 B.n233 B.n198 163.367
R543 B.n233 B.n232 163.367
R544 B.n232 B.n231 163.367
R545 B.n231 B.n200 163.367
R546 B.n227 B.n200 163.367
R547 B.n227 B.n226 163.367
R548 B.n226 B.n225 163.367
R549 B.n225 B.n202 163.367
R550 B.n221 B.n202 163.367
R551 B.n221 B.n220 163.367
R552 B.n220 B.n219 163.367
R553 B.n219 B.n204 163.367
R554 B.n215 B.n204 163.367
R555 B.n215 B.n214 163.367
R556 B.n214 B.n213 163.367
R557 B.n213 B.n206 163.367
R558 B.n209 B.n206 163.367
R559 B.n209 B.n208 163.367
R560 B.n208 B.n2 163.367
R561 B.n798 B.n2 163.367
R562 B.n798 B.n797 163.367
R563 B.n797 B.n796 163.367
R564 B.n796 B.n3 163.367
R565 B.n792 B.n3 163.367
R566 B.n792 B.n791 163.367
R567 B.n791 B.n790 163.367
R568 B.n790 B.n5 163.367
R569 B.n786 B.n5 163.367
R570 B.n786 B.n785 163.367
R571 B.n785 B.n784 163.367
R572 B.n784 B.n7 163.367
R573 B.n780 B.n7 163.367
R574 B.n780 B.n779 163.367
R575 B.n779 B.n778 163.367
R576 B.n778 B.n9 163.367
R577 B.n774 B.n9 163.367
R578 B.n774 B.n773 163.367
R579 B.n773 B.n772 163.367
R580 B.n772 B.n11 163.367
R581 B.n768 B.n11 163.367
R582 B.n768 B.n767 163.367
R583 B.n767 B.n766 163.367
R584 B.n766 B.n13 163.367
R585 B.n762 B.n13 163.367
R586 B.n762 B.n761 163.367
R587 B.n761 B.n760 163.367
R588 B.n760 B.n15 163.367
R589 B.n756 B.n15 163.367
R590 B.n756 B.n755 163.367
R591 B.n755 B.n754 163.367
R592 B.n251 B.n192 163.367
R593 B.n255 B.n192 163.367
R594 B.n256 B.n255 163.367
R595 B.n257 B.n256 163.367
R596 B.n257 B.n190 163.367
R597 B.n261 B.n190 163.367
R598 B.n262 B.n261 163.367
R599 B.n263 B.n262 163.367
R600 B.n263 B.n188 163.367
R601 B.n267 B.n188 163.367
R602 B.n268 B.n267 163.367
R603 B.n269 B.n268 163.367
R604 B.n269 B.n186 163.367
R605 B.n273 B.n186 163.367
R606 B.n274 B.n273 163.367
R607 B.n275 B.n274 163.367
R608 B.n275 B.n184 163.367
R609 B.n279 B.n184 163.367
R610 B.n280 B.n279 163.367
R611 B.n281 B.n280 163.367
R612 B.n281 B.n182 163.367
R613 B.n285 B.n182 163.367
R614 B.n286 B.n285 163.367
R615 B.n287 B.n286 163.367
R616 B.n287 B.n180 163.367
R617 B.n291 B.n180 163.367
R618 B.n292 B.n291 163.367
R619 B.n293 B.n292 163.367
R620 B.n293 B.n178 163.367
R621 B.n297 B.n178 163.367
R622 B.n298 B.n297 163.367
R623 B.n299 B.n298 163.367
R624 B.n299 B.n176 163.367
R625 B.n303 B.n176 163.367
R626 B.n304 B.n303 163.367
R627 B.n305 B.n304 163.367
R628 B.n305 B.n174 163.367
R629 B.n309 B.n174 163.367
R630 B.n310 B.n309 163.367
R631 B.n311 B.n310 163.367
R632 B.n311 B.n172 163.367
R633 B.n315 B.n172 163.367
R634 B.n316 B.n315 163.367
R635 B.n317 B.n316 163.367
R636 B.n317 B.n170 163.367
R637 B.n321 B.n170 163.367
R638 B.n322 B.n321 163.367
R639 B.n323 B.n322 163.367
R640 B.n323 B.n168 163.367
R641 B.n327 B.n168 163.367
R642 B.n328 B.n327 163.367
R643 B.n329 B.n328 163.367
R644 B.n329 B.n166 163.367
R645 B.n333 B.n166 163.367
R646 B.n334 B.n333 163.367
R647 B.n335 B.n334 163.367
R648 B.n335 B.n164 163.367
R649 B.n339 B.n164 163.367
R650 B.n340 B.n339 163.367
R651 B.n341 B.n340 163.367
R652 B.n341 B.n162 163.367
R653 B.n345 B.n162 163.367
R654 B.n346 B.n345 163.367
R655 B.n346 B.n158 163.367
R656 B.n350 B.n158 163.367
R657 B.n351 B.n350 163.367
R658 B.n352 B.n351 163.367
R659 B.n352 B.n156 163.367
R660 B.n356 B.n156 163.367
R661 B.n357 B.n356 163.367
R662 B.n358 B.n357 163.367
R663 B.n358 B.n152 163.367
R664 B.n363 B.n152 163.367
R665 B.n364 B.n363 163.367
R666 B.n365 B.n364 163.367
R667 B.n365 B.n150 163.367
R668 B.n369 B.n150 163.367
R669 B.n370 B.n369 163.367
R670 B.n371 B.n370 163.367
R671 B.n371 B.n148 163.367
R672 B.n375 B.n148 163.367
R673 B.n376 B.n375 163.367
R674 B.n377 B.n376 163.367
R675 B.n377 B.n146 163.367
R676 B.n381 B.n146 163.367
R677 B.n382 B.n381 163.367
R678 B.n383 B.n382 163.367
R679 B.n383 B.n144 163.367
R680 B.n387 B.n144 163.367
R681 B.n388 B.n387 163.367
R682 B.n389 B.n388 163.367
R683 B.n389 B.n142 163.367
R684 B.n393 B.n142 163.367
R685 B.n394 B.n393 163.367
R686 B.n395 B.n394 163.367
R687 B.n395 B.n140 163.367
R688 B.n399 B.n140 163.367
R689 B.n400 B.n399 163.367
R690 B.n401 B.n400 163.367
R691 B.n401 B.n138 163.367
R692 B.n405 B.n138 163.367
R693 B.n406 B.n405 163.367
R694 B.n407 B.n406 163.367
R695 B.n407 B.n136 163.367
R696 B.n411 B.n136 163.367
R697 B.n412 B.n411 163.367
R698 B.n413 B.n412 163.367
R699 B.n413 B.n134 163.367
R700 B.n417 B.n134 163.367
R701 B.n418 B.n417 163.367
R702 B.n419 B.n418 163.367
R703 B.n419 B.n132 163.367
R704 B.n423 B.n132 163.367
R705 B.n424 B.n423 163.367
R706 B.n425 B.n424 163.367
R707 B.n425 B.n130 163.367
R708 B.n429 B.n130 163.367
R709 B.n430 B.n429 163.367
R710 B.n431 B.n430 163.367
R711 B.n431 B.n128 163.367
R712 B.n435 B.n128 163.367
R713 B.n436 B.n435 163.367
R714 B.n437 B.n436 163.367
R715 B.n437 B.n126 163.367
R716 B.n441 B.n126 163.367
R717 B.n442 B.n441 163.367
R718 B.n443 B.n442 163.367
R719 B.n443 B.n124 163.367
R720 B.n447 B.n124 163.367
R721 B.n448 B.n447 163.367
R722 B.n449 B.n448 163.367
R723 B.n449 B.n122 163.367
R724 B.n453 B.n122 163.367
R725 B.n454 B.n453 163.367
R726 B.n455 B.n454 163.367
R727 B.n459 B.n120 163.367
R728 B.n460 B.n459 163.367
R729 B.n461 B.n460 163.367
R730 B.n461 B.n118 163.367
R731 B.n465 B.n118 163.367
R732 B.n466 B.n465 163.367
R733 B.n467 B.n466 163.367
R734 B.n467 B.n116 163.367
R735 B.n471 B.n116 163.367
R736 B.n472 B.n471 163.367
R737 B.n473 B.n472 163.367
R738 B.n473 B.n114 163.367
R739 B.n477 B.n114 163.367
R740 B.n478 B.n477 163.367
R741 B.n479 B.n478 163.367
R742 B.n479 B.n112 163.367
R743 B.n483 B.n112 163.367
R744 B.n484 B.n483 163.367
R745 B.n485 B.n484 163.367
R746 B.n485 B.n110 163.367
R747 B.n489 B.n110 163.367
R748 B.n490 B.n489 163.367
R749 B.n491 B.n490 163.367
R750 B.n491 B.n108 163.367
R751 B.n495 B.n108 163.367
R752 B.n496 B.n495 163.367
R753 B.n497 B.n496 163.367
R754 B.n497 B.n106 163.367
R755 B.n501 B.n106 163.367
R756 B.n502 B.n501 163.367
R757 B.n503 B.n502 163.367
R758 B.n503 B.n104 163.367
R759 B.n507 B.n104 163.367
R760 B.n508 B.n507 163.367
R761 B.n509 B.n508 163.367
R762 B.n509 B.n102 163.367
R763 B.n513 B.n102 163.367
R764 B.n514 B.n513 163.367
R765 B.n515 B.n514 163.367
R766 B.n515 B.n100 163.367
R767 B.n519 B.n100 163.367
R768 B.n520 B.n519 163.367
R769 B.n521 B.n520 163.367
R770 B.n521 B.n98 163.367
R771 B.n525 B.n98 163.367
R772 B.n526 B.n525 163.367
R773 B.n527 B.n526 163.367
R774 B.n527 B.n96 163.367
R775 B.n531 B.n96 163.367
R776 B.n532 B.n531 163.367
R777 B.n533 B.n532 163.367
R778 B.n533 B.n94 163.367
R779 B.n537 B.n94 163.367
R780 B.n538 B.n537 163.367
R781 B.n539 B.n538 163.367
R782 B.n539 B.n92 163.367
R783 B.n543 B.n92 163.367
R784 B.n544 B.n543 163.367
R785 B.n545 B.n544 163.367
R786 B.n545 B.n90 163.367
R787 B.n750 B.n17 163.367
R788 B.n750 B.n749 163.367
R789 B.n749 B.n748 163.367
R790 B.n748 B.n19 163.367
R791 B.n744 B.n19 163.367
R792 B.n744 B.n743 163.367
R793 B.n743 B.n742 163.367
R794 B.n742 B.n21 163.367
R795 B.n738 B.n21 163.367
R796 B.n738 B.n737 163.367
R797 B.n737 B.n736 163.367
R798 B.n736 B.n23 163.367
R799 B.n732 B.n23 163.367
R800 B.n732 B.n731 163.367
R801 B.n731 B.n730 163.367
R802 B.n730 B.n25 163.367
R803 B.n726 B.n25 163.367
R804 B.n726 B.n725 163.367
R805 B.n725 B.n724 163.367
R806 B.n724 B.n27 163.367
R807 B.n720 B.n27 163.367
R808 B.n720 B.n719 163.367
R809 B.n719 B.n718 163.367
R810 B.n718 B.n29 163.367
R811 B.n714 B.n29 163.367
R812 B.n714 B.n713 163.367
R813 B.n713 B.n712 163.367
R814 B.n712 B.n31 163.367
R815 B.n708 B.n31 163.367
R816 B.n708 B.n707 163.367
R817 B.n707 B.n706 163.367
R818 B.n706 B.n33 163.367
R819 B.n702 B.n33 163.367
R820 B.n702 B.n701 163.367
R821 B.n701 B.n700 163.367
R822 B.n700 B.n35 163.367
R823 B.n696 B.n35 163.367
R824 B.n696 B.n695 163.367
R825 B.n695 B.n694 163.367
R826 B.n694 B.n37 163.367
R827 B.n690 B.n37 163.367
R828 B.n690 B.n689 163.367
R829 B.n689 B.n688 163.367
R830 B.n688 B.n39 163.367
R831 B.n684 B.n39 163.367
R832 B.n684 B.n683 163.367
R833 B.n683 B.n682 163.367
R834 B.n682 B.n41 163.367
R835 B.n678 B.n41 163.367
R836 B.n678 B.n677 163.367
R837 B.n677 B.n676 163.367
R838 B.n676 B.n43 163.367
R839 B.n672 B.n43 163.367
R840 B.n672 B.n671 163.367
R841 B.n671 B.n670 163.367
R842 B.n670 B.n45 163.367
R843 B.n666 B.n45 163.367
R844 B.n666 B.n665 163.367
R845 B.n665 B.n664 163.367
R846 B.n664 B.n47 163.367
R847 B.n660 B.n47 163.367
R848 B.n660 B.n659 163.367
R849 B.n659 B.n658 163.367
R850 B.n658 B.n49 163.367
R851 B.n654 B.n49 163.367
R852 B.n654 B.n653 163.367
R853 B.n653 B.n652 163.367
R854 B.n652 B.n54 163.367
R855 B.n648 B.n54 163.367
R856 B.n648 B.n647 163.367
R857 B.n647 B.n646 163.367
R858 B.n646 B.n56 163.367
R859 B.n641 B.n56 163.367
R860 B.n641 B.n640 163.367
R861 B.n640 B.n639 163.367
R862 B.n639 B.n60 163.367
R863 B.n635 B.n60 163.367
R864 B.n635 B.n634 163.367
R865 B.n634 B.n633 163.367
R866 B.n633 B.n62 163.367
R867 B.n629 B.n62 163.367
R868 B.n629 B.n628 163.367
R869 B.n628 B.n627 163.367
R870 B.n627 B.n64 163.367
R871 B.n623 B.n64 163.367
R872 B.n623 B.n622 163.367
R873 B.n622 B.n621 163.367
R874 B.n621 B.n66 163.367
R875 B.n617 B.n66 163.367
R876 B.n617 B.n616 163.367
R877 B.n616 B.n615 163.367
R878 B.n615 B.n68 163.367
R879 B.n611 B.n68 163.367
R880 B.n611 B.n610 163.367
R881 B.n610 B.n609 163.367
R882 B.n609 B.n70 163.367
R883 B.n605 B.n70 163.367
R884 B.n605 B.n604 163.367
R885 B.n604 B.n603 163.367
R886 B.n603 B.n72 163.367
R887 B.n599 B.n72 163.367
R888 B.n599 B.n598 163.367
R889 B.n598 B.n597 163.367
R890 B.n597 B.n74 163.367
R891 B.n593 B.n74 163.367
R892 B.n593 B.n592 163.367
R893 B.n592 B.n591 163.367
R894 B.n591 B.n76 163.367
R895 B.n587 B.n76 163.367
R896 B.n587 B.n586 163.367
R897 B.n586 B.n585 163.367
R898 B.n585 B.n78 163.367
R899 B.n581 B.n78 163.367
R900 B.n581 B.n580 163.367
R901 B.n580 B.n579 163.367
R902 B.n579 B.n80 163.367
R903 B.n575 B.n80 163.367
R904 B.n575 B.n574 163.367
R905 B.n574 B.n573 163.367
R906 B.n573 B.n82 163.367
R907 B.n569 B.n82 163.367
R908 B.n569 B.n568 163.367
R909 B.n568 B.n567 163.367
R910 B.n567 B.n84 163.367
R911 B.n563 B.n84 163.367
R912 B.n563 B.n562 163.367
R913 B.n562 B.n561 163.367
R914 B.n561 B.n86 163.367
R915 B.n557 B.n86 163.367
R916 B.n557 B.n556 163.367
R917 B.n556 B.n555 163.367
R918 B.n555 B.n88 163.367
R919 B.n551 B.n88 163.367
R920 B.n551 B.n550 163.367
R921 B.n550 B.n549 163.367
R922 B.n153 B.t2 135.368
R923 B.n57 B.t4 135.368
R924 B.n159 B.t8 135.343
R925 B.n50 B.t10 135.343
R926 B.n154 B.t1 111.513
R927 B.n58 B.t5 111.513
R928 B.n160 B.t7 111.487
R929 B.n51 B.t11 111.487
R930 B.n361 B.n154 59.5399
R931 B.n161 B.n160 59.5399
R932 B.n52 B.n51 59.5399
R933 B.n643 B.n58 59.5399
R934 B.n753 B.n752 29.8151
R935 B.n457 B.n456 29.8151
R936 B.n252 B.n193 29.8151
R937 B.n548 B.n547 29.8151
R938 B.n154 B.n153 23.855
R939 B.n160 B.n159 23.855
R940 B.n51 B.n50 23.855
R941 B.n58 B.n57 23.855
R942 B B.n799 18.0485
R943 B.n752 B.n751 10.6151
R944 B.n751 B.n18 10.6151
R945 B.n747 B.n18 10.6151
R946 B.n747 B.n746 10.6151
R947 B.n746 B.n745 10.6151
R948 B.n745 B.n20 10.6151
R949 B.n741 B.n20 10.6151
R950 B.n741 B.n740 10.6151
R951 B.n740 B.n739 10.6151
R952 B.n739 B.n22 10.6151
R953 B.n735 B.n22 10.6151
R954 B.n735 B.n734 10.6151
R955 B.n734 B.n733 10.6151
R956 B.n733 B.n24 10.6151
R957 B.n729 B.n24 10.6151
R958 B.n729 B.n728 10.6151
R959 B.n728 B.n727 10.6151
R960 B.n727 B.n26 10.6151
R961 B.n723 B.n26 10.6151
R962 B.n723 B.n722 10.6151
R963 B.n722 B.n721 10.6151
R964 B.n721 B.n28 10.6151
R965 B.n717 B.n28 10.6151
R966 B.n717 B.n716 10.6151
R967 B.n716 B.n715 10.6151
R968 B.n715 B.n30 10.6151
R969 B.n711 B.n30 10.6151
R970 B.n711 B.n710 10.6151
R971 B.n710 B.n709 10.6151
R972 B.n709 B.n32 10.6151
R973 B.n705 B.n32 10.6151
R974 B.n705 B.n704 10.6151
R975 B.n704 B.n703 10.6151
R976 B.n703 B.n34 10.6151
R977 B.n699 B.n34 10.6151
R978 B.n699 B.n698 10.6151
R979 B.n698 B.n697 10.6151
R980 B.n697 B.n36 10.6151
R981 B.n693 B.n36 10.6151
R982 B.n693 B.n692 10.6151
R983 B.n692 B.n691 10.6151
R984 B.n691 B.n38 10.6151
R985 B.n687 B.n38 10.6151
R986 B.n687 B.n686 10.6151
R987 B.n686 B.n685 10.6151
R988 B.n685 B.n40 10.6151
R989 B.n681 B.n40 10.6151
R990 B.n681 B.n680 10.6151
R991 B.n680 B.n679 10.6151
R992 B.n679 B.n42 10.6151
R993 B.n675 B.n42 10.6151
R994 B.n675 B.n674 10.6151
R995 B.n674 B.n673 10.6151
R996 B.n673 B.n44 10.6151
R997 B.n669 B.n44 10.6151
R998 B.n669 B.n668 10.6151
R999 B.n668 B.n667 10.6151
R1000 B.n667 B.n46 10.6151
R1001 B.n663 B.n46 10.6151
R1002 B.n663 B.n662 10.6151
R1003 B.n662 B.n661 10.6151
R1004 B.n661 B.n48 10.6151
R1005 B.n657 B.n656 10.6151
R1006 B.n656 B.n655 10.6151
R1007 B.n655 B.n53 10.6151
R1008 B.n651 B.n53 10.6151
R1009 B.n651 B.n650 10.6151
R1010 B.n650 B.n649 10.6151
R1011 B.n649 B.n55 10.6151
R1012 B.n645 B.n55 10.6151
R1013 B.n645 B.n644 10.6151
R1014 B.n642 B.n59 10.6151
R1015 B.n638 B.n59 10.6151
R1016 B.n638 B.n637 10.6151
R1017 B.n637 B.n636 10.6151
R1018 B.n636 B.n61 10.6151
R1019 B.n632 B.n61 10.6151
R1020 B.n632 B.n631 10.6151
R1021 B.n631 B.n630 10.6151
R1022 B.n630 B.n63 10.6151
R1023 B.n626 B.n63 10.6151
R1024 B.n626 B.n625 10.6151
R1025 B.n625 B.n624 10.6151
R1026 B.n624 B.n65 10.6151
R1027 B.n620 B.n65 10.6151
R1028 B.n620 B.n619 10.6151
R1029 B.n619 B.n618 10.6151
R1030 B.n618 B.n67 10.6151
R1031 B.n614 B.n67 10.6151
R1032 B.n614 B.n613 10.6151
R1033 B.n613 B.n612 10.6151
R1034 B.n612 B.n69 10.6151
R1035 B.n608 B.n69 10.6151
R1036 B.n608 B.n607 10.6151
R1037 B.n607 B.n606 10.6151
R1038 B.n606 B.n71 10.6151
R1039 B.n602 B.n71 10.6151
R1040 B.n602 B.n601 10.6151
R1041 B.n601 B.n600 10.6151
R1042 B.n600 B.n73 10.6151
R1043 B.n596 B.n73 10.6151
R1044 B.n596 B.n595 10.6151
R1045 B.n595 B.n594 10.6151
R1046 B.n594 B.n75 10.6151
R1047 B.n590 B.n75 10.6151
R1048 B.n590 B.n589 10.6151
R1049 B.n589 B.n588 10.6151
R1050 B.n588 B.n77 10.6151
R1051 B.n584 B.n77 10.6151
R1052 B.n584 B.n583 10.6151
R1053 B.n583 B.n582 10.6151
R1054 B.n582 B.n79 10.6151
R1055 B.n578 B.n79 10.6151
R1056 B.n578 B.n577 10.6151
R1057 B.n577 B.n576 10.6151
R1058 B.n576 B.n81 10.6151
R1059 B.n572 B.n81 10.6151
R1060 B.n572 B.n571 10.6151
R1061 B.n571 B.n570 10.6151
R1062 B.n570 B.n83 10.6151
R1063 B.n566 B.n83 10.6151
R1064 B.n566 B.n565 10.6151
R1065 B.n565 B.n564 10.6151
R1066 B.n564 B.n85 10.6151
R1067 B.n560 B.n85 10.6151
R1068 B.n560 B.n559 10.6151
R1069 B.n559 B.n558 10.6151
R1070 B.n558 B.n87 10.6151
R1071 B.n554 B.n87 10.6151
R1072 B.n554 B.n553 10.6151
R1073 B.n553 B.n552 10.6151
R1074 B.n552 B.n89 10.6151
R1075 B.n548 B.n89 10.6151
R1076 B.n458 B.n457 10.6151
R1077 B.n458 B.n119 10.6151
R1078 B.n462 B.n119 10.6151
R1079 B.n463 B.n462 10.6151
R1080 B.n464 B.n463 10.6151
R1081 B.n464 B.n117 10.6151
R1082 B.n468 B.n117 10.6151
R1083 B.n469 B.n468 10.6151
R1084 B.n470 B.n469 10.6151
R1085 B.n470 B.n115 10.6151
R1086 B.n474 B.n115 10.6151
R1087 B.n475 B.n474 10.6151
R1088 B.n476 B.n475 10.6151
R1089 B.n476 B.n113 10.6151
R1090 B.n480 B.n113 10.6151
R1091 B.n481 B.n480 10.6151
R1092 B.n482 B.n481 10.6151
R1093 B.n482 B.n111 10.6151
R1094 B.n486 B.n111 10.6151
R1095 B.n487 B.n486 10.6151
R1096 B.n488 B.n487 10.6151
R1097 B.n488 B.n109 10.6151
R1098 B.n492 B.n109 10.6151
R1099 B.n493 B.n492 10.6151
R1100 B.n494 B.n493 10.6151
R1101 B.n494 B.n107 10.6151
R1102 B.n498 B.n107 10.6151
R1103 B.n499 B.n498 10.6151
R1104 B.n500 B.n499 10.6151
R1105 B.n500 B.n105 10.6151
R1106 B.n504 B.n105 10.6151
R1107 B.n505 B.n504 10.6151
R1108 B.n506 B.n505 10.6151
R1109 B.n506 B.n103 10.6151
R1110 B.n510 B.n103 10.6151
R1111 B.n511 B.n510 10.6151
R1112 B.n512 B.n511 10.6151
R1113 B.n512 B.n101 10.6151
R1114 B.n516 B.n101 10.6151
R1115 B.n517 B.n516 10.6151
R1116 B.n518 B.n517 10.6151
R1117 B.n518 B.n99 10.6151
R1118 B.n522 B.n99 10.6151
R1119 B.n523 B.n522 10.6151
R1120 B.n524 B.n523 10.6151
R1121 B.n524 B.n97 10.6151
R1122 B.n528 B.n97 10.6151
R1123 B.n529 B.n528 10.6151
R1124 B.n530 B.n529 10.6151
R1125 B.n530 B.n95 10.6151
R1126 B.n534 B.n95 10.6151
R1127 B.n535 B.n534 10.6151
R1128 B.n536 B.n535 10.6151
R1129 B.n536 B.n93 10.6151
R1130 B.n540 B.n93 10.6151
R1131 B.n541 B.n540 10.6151
R1132 B.n542 B.n541 10.6151
R1133 B.n542 B.n91 10.6151
R1134 B.n546 B.n91 10.6151
R1135 B.n547 B.n546 10.6151
R1136 B.n253 B.n252 10.6151
R1137 B.n254 B.n253 10.6151
R1138 B.n254 B.n191 10.6151
R1139 B.n258 B.n191 10.6151
R1140 B.n259 B.n258 10.6151
R1141 B.n260 B.n259 10.6151
R1142 B.n260 B.n189 10.6151
R1143 B.n264 B.n189 10.6151
R1144 B.n265 B.n264 10.6151
R1145 B.n266 B.n265 10.6151
R1146 B.n266 B.n187 10.6151
R1147 B.n270 B.n187 10.6151
R1148 B.n271 B.n270 10.6151
R1149 B.n272 B.n271 10.6151
R1150 B.n272 B.n185 10.6151
R1151 B.n276 B.n185 10.6151
R1152 B.n277 B.n276 10.6151
R1153 B.n278 B.n277 10.6151
R1154 B.n278 B.n183 10.6151
R1155 B.n282 B.n183 10.6151
R1156 B.n283 B.n282 10.6151
R1157 B.n284 B.n283 10.6151
R1158 B.n284 B.n181 10.6151
R1159 B.n288 B.n181 10.6151
R1160 B.n289 B.n288 10.6151
R1161 B.n290 B.n289 10.6151
R1162 B.n290 B.n179 10.6151
R1163 B.n294 B.n179 10.6151
R1164 B.n295 B.n294 10.6151
R1165 B.n296 B.n295 10.6151
R1166 B.n296 B.n177 10.6151
R1167 B.n300 B.n177 10.6151
R1168 B.n301 B.n300 10.6151
R1169 B.n302 B.n301 10.6151
R1170 B.n302 B.n175 10.6151
R1171 B.n306 B.n175 10.6151
R1172 B.n307 B.n306 10.6151
R1173 B.n308 B.n307 10.6151
R1174 B.n308 B.n173 10.6151
R1175 B.n312 B.n173 10.6151
R1176 B.n313 B.n312 10.6151
R1177 B.n314 B.n313 10.6151
R1178 B.n314 B.n171 10.6151
R1179 B.n318 B.n171 10.6151
R1180 B.n319 B.n318 10.6151
R1181 B.n320 B.n319 10.6151
R1182 B.n320 B.n169 10.6151
R1183 B.n324 B.n169 10.6151
R1184 B.n325 B.n324 10.6151
R1185 B.n326 B.n325 10.6151
R1186 B.n326 B.n167 10.6151
R1187 B.n330 B.n167 10.6151
R1188 B.n331 B.n330 10.6151
R1189 B.n332 B.n331 10.6151
R1190 B.n332 B.n165 10.6151
R1191 B.n336 B.n165 10.6151
R1192 B.n337 B.n336 10.6151
R1193 B.n338 B.n337 10.6151
R1194 B.n338 B.n163 10.6151
R1195 B.n342 B.n163 10.6151
R1196 B.n343 B.n342 10.6151
R1197 B.n344 B.n343 10.6151
R1198 B.n348 B.n347 10.6151
R1199 B.n349 B.n348 10.6151
R1200 B.n349 B.n157 10.6151
R1201 B.n353 B.n157 10.6151
R1202 B.n354 B.n353 10.6151
R1203 B.n355 B.n354 10.6151
R1204 B.n355 B.n155 10.6151
R1205 B.n359 B.n155 10.6151
R1206 B.n360 B.n359 10.6151
R1207 B.n362 B.n151 10.6151
R1208 B.n366 B.n151 10.6151
R1209 B.n367 B.n366 10.6151
R1210 B.n368 B.n367 10.6151
R1211 B.n368 B.n149 10.6151
R1212 B.n372 B.n149 10.6151
R1213 B.n373 B.n372 10.6151
R1214 B.n374 B.n373 10.6151
R1215 B.n374 B.n147 10.6151
R1216 B.n378 B.n147 10.6151
R1217 B.n379 B.n378 10.6151
R1218 B.n380 B.n379 10.6151
R1219 B.n380 B.n145 10.6151
R1220 B.n384 B.n145 10.6151
R1221 B.n385 B.n384 10.6151
R1222 B.n386 B.n385 10.6151
R1223 B.n386 B.n143 10.6151
R1224 B.n390 B.n143 10.6151
R1225 B.n391 B.n390 10.6151
R1226 B.n392 B.n391 10.6151
R1227 B.n392 B.n141 10.6151
R1228 B.n396 B.n141 10.6151
R1229 B.n397 B.n396 10.6151
R1230 B.n398 B.n397 10.6151
R1231 B.n398 B.n139 10.6151
R1232 B.n402 B.n139 10.6151
R1233 B.n403 B.n402 10.6151
R1234 B.n404 B.n403 10.6151
R1235 B.n404 B.n137 10.6151
R1236 B.n408 B.n137 10.6151
R1237 B.n409 B.n408 10.6151
R1238 B.n410 B.n409 10.6151
R1239 B.n410 B.n135 10.6151
R1240 B.n414 B.n135 10.6151
R1241 B.n415 B.n414 10.6151
R1242 B.n416 B.n415 10.6151
R1243 B.n416 B.n133 10.6151
R1244 B.n420 B.n133 10.6151
R1245 B.n421 B.n420 10.6151
R1246 B.n422 B.n421 10.6151
R1247 B.n422 B.n131 10.6151
R1248 B.n426 B.n131 10.6151
R1249 B.n427 B.n426 10.6151
R1250 B.n428 B.n427 10.6151
R1251 B.n428 B.n129 10.6151
R1252 B.n432 B.n129 10.6151
R1253 B.n433 B.n432 10.6151
R1254 B.n434 B.n433 10.6151
R1255 B.n434 B.n127 10.6151
R1256 B.n438 B.n127 10.6151
R1257 B.n439 B.n438 10.6151
R1258 B.n440 B.n439 10.6151
R1259 B.n440 B.n125 10.6151
R1260 B.n444 B.n125 10.6151
R1261 B.n445 B.n444 10.6151
R1262 B.n446 B.n445 10.6151
R1263 B.n446 B.n123 10.6151
R1264 B.n450 B.n123 10.6151
R1265 B.n451 B.n450 10.6151
R1266 B.n452 B.n451 10.6151
R1267 B.n452 B.n121 10.6151
R1268 B.n456 B.n121 10.6151
R1269 B.n248 B.n193 10.6151
R1270 B.n248 B.n247 10.6151
R1271 B.n247 B.n246 10.6151
R1272 B.n246 B.n195 10.6151
R1273 B.n242 B.n195 10.6151
R1274 B.n242 B.n241 10.6151
R1275 B.n241 B.n240 10.6151
R1276 B.n240 B.n197 10.6151
R1277 B.n236 B.n197 10.6151
R1278 B.n236 B.n235 10.6151
R1279 B.n235 B.n234 10.6151
R1280 B.n234 B.n199 10.6151
R1281 B.n230 B.n199 10.6151
R1282 B.n230 B.n229 10.6151
R1283 B.n229 B.n228 10.6151
R1284 B.n228 B.n201 10.6151
R1285 B.n224 B.n201 10.6151
R1286 B.n224 B.n223 10.6151
R1287 B.n223 B.n222 10.6151
R1288 B.n222 B.n203 10.6151
R1289 B.n218 B.n203 10.6151
R1290 B.n218 B.n217 10.6151
R1291 B.n217 B.n216 10.6151
R1292 B.n216 B.n205 10.6151
R1293 B.n212 B.n205 10.6151
R1294 B.n212 B.n211 10.6151
R1295 B.n211 B.n210 10.6151
R1296 B.n210 B.n207 10.6151
R1297 B.n207 B.n0 10.6151
R1298 B.n795 B.n1 10.6151
R1299 B.n795 B.n794 10.6151
R1300 B.n794 B.n793 10.6151
R1301 B.n793 B.n4 10.6151
R1302 B.n789 B.n4 10.6151
R1303 B.n789 B.n788 10.6151
R1304 B.n788 B.n787 10.6151
R1305 B.n787 B.n6 10.6151
R1306 B.n783 B.n6 10.6151
R1307 B.n783 B.n782 10.6151
R1308 B.n782 B.n781 10.6151
R1309 B.n781 B.n8 10.6151
R1310 B.n777 B.n8 10.6151
R1311 B.n777 B.n776 10.6151
R1312 B.n776 B.n775 10.6151
R1313 B.n775 B.n10 10.6151
R1314 B.n771 B.n10 10.6151
R1315 B.n771 B.n770 10.6151
R1316 B.n770 B.n769 10.6151
R1317 B.n769 B.n12 10.6151
R1318 B.n765 B.n12 10.6151
R1319 B.n765 B.n764 10.6151
R1320 B.n764 B.n763 10.6151
R1321 B.n763 B.n14 10.6151
R1322 B.n759 B.n14 10.6151
R1323 B.n759 B.n758 10.6151
R1324 B.n758 B.n757 10.6151
R1325 B.n757 B.n16 10.6151
R1326 B.n753 B.n16 10.6151
R1327 B.n52 B.n48 9.36635
R1328 B.n643 B.n642 9.36635
R1329 B.n344 B.n161 9.36635
R1330 B.n362 B.n361 9.36635
R1331 B.n799 B.n0 2.81026
R1332 B.n799 B.n1 2.81026
R1333 B.n657 B.n52 1.24928
R1334 B.n644 B.n643 1.24928
R1335 B.n347 B.n161 1.24928
R1336 B.n361 B.n360 1.24928
R1337 VN.n4 VN.t2 576.934
R1338 VN.n23 VN.t0 576.934
R1339 VN.n17 VN.t9 560.995
R1340 VN.n36 VN.t4 560.995
R1341 VN.n10 VN.t5 517.347
R1342 VN.n5 VN.t3 517.347
R1343 VN.n1 VN.t6 517.347
R1344 VN.n29 VN.t1 517.347
R1345 VN.n24 VN.t7 517.347
R1346 VN.n20 VN.t8 517.347
R1347 VN.n18 VN.n17 161.3
R1348 VN.n37 VN.n36 161.3
R1349 VN.n35 VN.n19 161.3
R1350 VN.n34 VN.n33 161.3
R1351 VN.n32 VN.n31 161.3
R1352 VN.n30 VN.n21 161.3
R1353 VN.n29 VN.n28 161.3
R1354 VN.n27 VN.n22 161.3
R1355 VN.n26 VN.n25 161.3
R1356 VN.n16 VN.n0 161.3
R1357 VN.n15 VN.n14 161.3
R1358 VN.n13 VN.n12 161.3
R1359 VN.n11 VN.n2 161.3
R1360 VN.n10 VN.n9 161.3
R1361 VN.n8 VN.n3 161.3
R1362 VN.n7 VN.n6 161.3
R1363 VN.n16 VN.n15 55.593
R1364 VN.n35 VN.n34 55.593
R1365 VN.n6 VN.n3 51.7179
R1366 VN.n12 VN.n11 51.7179
R1367 VN.n25 VN.n22 51.7179
R1368 VN.n31 VN.n30 51.7179
R1369 VN VN.n37 49.7713
R1370 VN.n26 VN.n23 43.7549
R1371 VN.n7 VN.n4 43.7549
R1372 VN.n5 VN.n4 43.7503
R1373 VN.n24 VN.n23 43.7503
R1374 VN.n10 VN.n3 29.4362
R1375 VN.n11 VN.n10 29.4362
R1376 VN.n29 VN.n22 29.4362
R1377 VN.n30 VN.n29 29.4362
R1378 VN.n15 VN.n1 13.2801
R1379 VN.n34 VN.n20 13.2801
R1380 VN.n6 VN.n5 11.3127
R1381 VN.n12 VN.n1 11.3127
R1382 VN.n25 VN.n24 11.3127
R1383 VN.n31 VN.n20 11.3127
R1384 VN.n17 VN.n16 1.46111
R1385 VN.n36 VN.n35 1.46111
R1386 VN.n37 VN.n19 0.189894
R1387 VN.n33 VN.n19 0.189894
R1388 VN.n33 VN.n32 0.189894
R1389 VN.n32 VN.n21 0.189894
R1390 VN.n28 VN.n21 0.189894
R1391 VN.n28 VN.n27 0.189894
R1392 VN.n27 VN.n26 0.189894
R1393 VN.n8 VN.n7 0.189894
R1394 VN.n9 VN.n8 0.189894
R1395 VN.n9 VN.n2 0.189894
R1396 VN.n13 VN.n2 0.189894
R1397 VN.n14 VN.n13 0.189894
R1398 VN.n14 VN.n0 0.189894
R1399 VN.n18 VN.n0 0.189894
R1400 VN VN.n18 0.0516364
R1401 VDD2.n1 VDD2.t7 70.9864
R1402 VDD2.n4 VDD2.t5 69.9263
R1403 VDD2.n3 VDD2.n2 68.9838
R1404 VDD2 VDD2.n7 68.9808
R1405 VDD2.n6 VDD2.n5 68.2439
R1406 VDD2.n1 VDD2.n0 68.2438
R1407 VDD2.n4 VDD2.n3 45.4071
R1408 VDD2.n7 VDD2.t2 1.68295
R1409 VDD2.n7 VDD2.t9 1.68295
R1410 VDD2.n5 VDD2.t1 1.68295
R1411 VDD2.n5 VDD2.t8 1.68295
R1412 VDD2.n2 VDD2.t3 1.68295
R1413 VDD2.n2 VDD2.t0 1.68295
R1414 VDD2.n0 VDD2.t6 1.68295
R1415 VDD2.n0 VDD2.t4 1.68295
R1416 VDD2.n6 VDD2.n4 1.06084
R1417 VDD2 VDD2.n6 0.323776
R1418 VDD2.n3 VDD2.n1 0.21024
C0 VP w_n2446_n4832# 5.1587f
C1 w_n2446_n4832# VTAIL 4.14024f
C2 VP VDD2 0.368374f
C3 VDD2 VTAIL 18.9768f
C4 VDD1 B 2.33021f
C5 w_n2446_n4832# VN 4.84549f
C6 VDD2 VN 11.9282f
C7 B w_n2446_n4832# 9.74157f
C8 VDD1 w_n2446_n4832# 2.66202f
C9 B VDD2 2.38217f
C10 VDD1 VDD2 1.09999f
C11 VP VTAIL 11.5886f
C12 VP VN 7.24479f
C13 VDD2 w_n2446_n4832# 2.71716f
C14 VTAIL VN 11.5737f
C15 B VP 1.45553f
C16 VDD1 VP 12.139999f
C17 B VTAIL 4.21805f
C18 VDD1 VTAIL 18.944199f
C19 B VN 0.938226f
C20 VDD1 VN 0.149814f
C21 VDD2 VSUBS 1.794566f
C22 VDD1 VSUBS 1.469084f
C23 VTAIL VSUBS 1.06517f
C24 VN VSUBS 5.66412f
C25 VP VSUBS 2.343568f
C26 B VSUBS 3.879079f
C27 w_n2446_n4832# VSUBS 0.144382p
C28 VDD2.t7 VSUBS 4.54928f
C29 VDD2.t6 VSUBS 0.417918f
C30 VDD2.t4 VSUBS 0.417918f
C31 VDD2.n0 VSUBS 3.49985f
C32 VDD2.n1 VSUBS 1.40266f
C33 VDD2.t3 VSUBS 0.417918f
C34 VDD2.t0 VSUBS 0.417918f
C35 VDD2.n2 VSUBS 3.50754f
C36 VDD2.n3 VSUBS 3.01686f
C37 VDD2.t5 VSUBS 4.53805f
C38 VDD2.n4 VSUBS 3.66487f
C39 VDD2.t1 VSUBS 0.417918f
C40 VDD2.t8 VSUBS 0.417918f
C41 VDD2.n5 VSUBS 3.49985f
C42 VDD2.n6 VSUBS 0.668401f
C43 VDD2.t2 VSUBS 0.417918f
C44 VDD2.t9 VSUBS 0.417918f
C45 VDD2.n7 VSUBS 3.50748f
C46 VN.n0 VSUBS 0.043973f
C47 VN.t6 VSUBS 2.1058f
C48 VN.n1 VSUBS 0.754513f
C49 VN.n2 VSUBS 0.043973f
C50 VN.t5 VSUBS 2.1058f
C51 VN.n3 VSUBS 0.043533f
C52 VN.t2 VSUBS 2.18853f
C53 VN.n4 VSUBS 0.809413f
C54 VN.t3 VSUBS 2.1058f
C55 VN.n5 VSUBS 0.794154f
C56 VN.n6 VSUBS 0.057272f
C57 VN.n7 VSUBS 0.183671f
C58 VN.n8 VSUBS 0.043973f
C59 VN.n9 VSUBS 0.043973f
C60 VN.n10 VSUBS 0.8064f
C61 VN.n11 VSUBS 0.043533f
C62 VN.n12 VSUBS 0.057272f
C63 VN.n13 VSUBS 0.043973f
C64 VN.n14 VSUBS 0.043973f
C65 VN.n15 VSUBS 0.05674f
C66 VN.n16 VSUBS 0.013668f
C67 VN.t9 VSUBS 2.16606f
C68 VN.n17 VSUBS 0.800221f
C69 VN.n18 VSUBS 0.034077f
C70 VN.n19 VSUBS 0.043973f
C71 VN.t8 VSUBS 2.1058f
C72 VN.n20 VSUBS 0.754513f
C73 VN.n21 VSUBS 0.043973f
C74 VN.t1 VSUBS 2.1058f
C75 VN.n22 VSUBS 0.043533f
C76 VN.t0 VSUBS 2.18853f
C77 VN.n23 VSUBS 0.809413f
C78 VN.t7 VSUBS 2.1058f
C79 VN.n24 VSUBS 0.794154f
C80 VN.n25 VSUBS 0.057272f
C81 VN.n26 VSUBS 0.183671f
C82 VN.n27 VSUBS 0.043973f
C83 VN.n28 VSUBS 0.043973f
C84 VN.n29 VSUBS 0.8064f
C85 VN.n30 VSUBS 0.043533f
C86 VN.n31 VSUBS 0.057272f
C87 VN.n32 VSUBS 0.043973f
C88 VN.n33 VSUBS 0.043973f
C89 VN.n34 VSUBS 0.05674f
C90 VN.n35 VSUBS 0.013668f
C91 VN.t4 VSUBS 2.16606f
C92 VN.n36 VSUBS 0.800221f
C93 VN.n37 VSUBS 2.37542f
C94 B.n0 VSUBS 0.005491f
C95 B.n1 VSUBS 0.005491f
C96 B.n2 VSUBS 0.008684f
C97 B.n3 VSUBS 0.008684f
C98 B.n4 VSUBS 0.008684f
C99 B.n5 VSUBS 0.008684f
C100 B.n6 VSUBS 0.008684f
C101 B.n7 VSUBS 0.008684f
C102 B.n8 VSUBS 0.008684f
C103 B.n9 VSUBS 0.008684f
C104 B.n10 VSUBS 0.008684f
C105 B.n11 VSUBS 0.008684f
C106 B.n12 VSUBS 0.008684f
C107 B.n13 VSUBS 0.008684f
C108 B.n14 VSUBS 0.008684f
C109 B.n15 VSUBS 0.008684f
C110 B.n16 VSUBS 0.008684f
C111 B.n17 VSUBS 0.01958f
C112 B.n18 VSUBS 0.008684f
C113 B.n19 VSUBS 0.008684f
C114 B.n20 VSUBS 0.008684f
C115 B.n21 VSUBS 0.008684f
C116 B.n22 VSUBS 0.008684f
C117 B.n23 VSUBS 0.008684f
C118 B.n24 VSUBS 0.008684f
C119 B.n25 VSUBS 0.008684f
C120 B.n26 VSUBS 0.008684f
C121 B.n27 VSUBS 0.008684f
C122 B.n28 VSUBS 0.008684f
C123 B.n29 VSUBS 0.008684f
C124 B.n30 VSUBS 0.008684f
C125 B.n31 VSUBS 0.008684f
C126 B.n32 VSUBS 0.008684f
C127 B.n33 VSUBS 0.008684f
C128 B.n34 VSUBS 0.008684f
C129 B.n35 VSUBS 0.008684f
C130 B.n36 VSUBS 0.008684f
C131 B.n37 VSUBS 0.008684f
C132 B.n38 VSUBS 0.008684f
C133 B.n39 VSUBS 0.008684f
C134 B.n40 VSUBS 0.008684f
C135 B.n41 VSUBS 0.008684f
C136 B.n42 VSUBS 0.008684f
C137 B.n43 VSUBS 0.008684f
C138 B.n44 VSUBS 0.008684f
C139 B.n45 VSUBS 0.008684f
C140 B.n46 VSUBS 0.008684f
C141 B.n47 VSUBS 0.008684f
C142 B.n48 VSUBS 0.008173f
C143 B.n49 VSUBS 0.008684f
C144 B.t11 VSUBS 0.813017f
C145 B.t10 VSUBS 0.825067f
C146 B.t9 VSUBS 0.879781f
C147 B.n50 VSUBS 0.279127f
C148 B.n51 VSUBS 0.080752f
C149 B.n52 VSUBS 0.020119f
C150 B.n53 VSUBS 0.008684f
C151 B.n54 VSUBS 0.008684f
C152 B.n55 VSUBS 0.008684f
C153 B.n56 VSUBS 0.008684f
C154 B.t5 VSUBS 0.812984f
C155 B.t4 VSUBS 0.825038f
C156 B.t3 VSUBS 0.879781f
C157 B.n57 VSUBS 0.279156f
C158 B.n58 VSUBS 0.080785f
C159 B.n59 VSUBS 0.008684f
C160 B.n60 VSUBS 0.008684f
C161 B.n61 VSUBS 0.008684f
C162 B.n62 VSUBS 0.008684f
C163 B.n63 VSUBS 0.008684f
C164 B.n64 VSUBS 0.008684f
C165 B.n65 VSUBS 0.008684f
C166 B.n66 VSUBS 0.008684f
C167 B.n67 VSUBS 0.008684f
C168 B.n68 VSUBS 0.008684f
C169 B.n69 VSUBS 0.008684f
C170 B.n70 VSUBS 0.008684f
C171 B.n71 VSUBS 0.008684f
C172 B.n72 VSUBS 0.008684f
C173 B.n73 VSUBS 0.008684f
C174 B.n74 VSUBS 0.008684f
C175 B.n75 VSUBS 0.008684f
C176 B.n76 VSUBS 0.008684f
C177 B.n77 VSUBS 0.008684f
C178 B.n78 VSUBS 0.008684f
C179 B.n79 VSUBS 0.008684f
C180 B.n80 VSUBS 0.008684f
C181 B.n81 VSUBS 0.008684f
C182 B.n82 VSUBS 0.008684f
C183 B.n83 VSUBS 0.008684f
C184 B.n84 VSUBS 0.008684f
C185 B.n85 VSUBS 0.008684f
C186 B.n86 VSUBS 0.008684f
C187 B.n87 VSUBS 0.008684f
C188 B.n88 VSUBS 0.008684f
C189 B.n89 VSUBS 0.008684f
C190 B.n90 VSUBS 0.01873f
C191 B.n91 VSUBS 0.008684f
C192 B.n92 VSUBS 0.008684f
C193 B.n93 VSUBS 0.008684f
C194 B.n94 VSUBS 0.008684f
C195 B.n95 VSUBS 0.008684f
C196 B.n96 VSUBS 0.008684f
C197 B.n97 VSUBS 0.008684f
C198 B.n98 VSUBS 0.008684f
C199 B.n99 VSUBS 0.008684f
C200 B.n100 VSUBS 0.008684f
C201 B.n101 VSUBS 0.008684f
C202 B.n102 VSUBS 0.008684f
C203 B.n103 VSUBS 0.008684f
C204 B.n104 VSUBS 0.008684f
C205 B.n105 VSUBS 0.008684f
C206 B.n106 VSUBS 0.008684f
C207 B.n107 VSUBS 0.008684f
C208 B.n108 VSUBS 0.008684f
C209 B.n109 VSUBS 0.008684f
C210 B.n110 VSUBS 0.008684f
C211 B.n111 VSUBS 0.008684f
C212 B.n112 VSUBS 0.008684f
C213 B.n113 VSUBS 0.008684f
C214 B.n114 VSUBS 0.008684f
C215 B.n115 VSUBS 0.008684f
C216 B.n116 VSUBS 0.008684f
C217 B.n117 VSUBS 0.008684f
C218 B.n118 VSUBS 0.008684f
C219 B.n119 VSUBS 0.008684f
C220 B.n120 VSUBS 0.01873f
C221 B.n121 VSUBS 0.008684f
C222 B.n122 VSUBS 0.008684f
C223 B.n123 VSUBS 0.008684f
C224 B.n124 VSUBS 0.008684f
C225 B.n125 VSUBS 0.008684f
C226 B.n126 VSUBS 0.008684f
C227 B.n127 VSUBS 0.008684f
C228 B.n128 VSUBS 0.008684f
C229 B.n129 VSUBS 0.008684f
C230 B.n130 VSUBS 0.008684f
C231 B.n131 VSUBS 0.008684f
C232 B.n132 VSUBS 0.008684f
C233 B.n133 VSUBS 0.008684f
C234 B.n134 VSUBS 0.008684f
C235 B.n135 VSUBS 0.008684f
C236 B.n136 VSUBS 0.008684f
C237 B.n137 VSUBS 0.008684f
C238 B.n138 VSUBS 0.008684f
C239 B.n139 VSUBS 0.008684f
C240 B.n140 VSUBS 0.008684f
C241 B.n141 VSUBS 0.008684f
C242 B.n142 VSUBS 0.008684f
C243 B.n143 VSUBS 0.008684f
C244 B.n144 VSUBS 0.008684f
C245 B.n145 VSUBS 0.008684f
C246 B.n146 VSUBS 0.008684f
C247 B.n147 VSUBS 0.008684f
C248 B.n148 VSUBS 0.008684f
C249 B.n149 VSUBS 0.008684f
C250 B.n150 VSUBS 0.008684f
C251 B.n151 VSUBS 0.008684f
C252 B.n152 VSUBS 0.008684f
C253 B.t1 VSUBS 0.812984f
C254 B.t2 VSUBS 0.825038f
C255 B.t0 VSUBS 0.879781f
C256 B.n153 VSUBS 0.279156f
C257 B.n154 VSUBS 0.080785f
C258 B.n155 VSUBS 0.008684f
C259 B.n156 VSUBS 0.008684f
C260 B.n157 VSUBS 0.008684f
C261 B.n158 VSUBS 0.008684f
C262 B.t7 VSUBS 0.813017f
C263 B.t8 VSUBS 0.825067f
C264 B.t6 VSUBS 0.879781f
C265 B.n159 VSUBS 0.279127f
C266 B.n160 VSUBS 0.080752f
C267 B.n161 VSUBS 0.020119f
C268 B.n162 VSUBS 0.008684f
C269 B.n163 VSUBS 0.008684f
C270 B.n164 VSUBS 0.008684f
C271 B.n165 VSUBS 0.008684f
C272 B.n166 VSUBS 0.008684f
C273 B.n167 VSUBS 0.008684f
C274 B.n168 VSUBS 0.008684f
C275 B.n169 VSUBS 0.008684f
C276 B.n170 VSUBS 0.008684f
C277 B.n171 VSUBS 0.008684f
C278 B.n172 VSUBS 0.008684f
C279 B.n173 VSUBS 0.008684f
C280 B.n174 VSUBS 0.008684f
C281 B.n175 VSUBS 0.008684f
C282 B.n176 VSUBS 0.008684f
C283 B.n177 VSUBS 0.008684f
C284 B.n178 VSUBS 0.008684f
C285 B.n179 VSUBS 0.008684f
C286 B.n180 VSUBS 0.008684f
C287 B.n181 VSUBS 0.008684f
C288 B.n182 VSUBS 0.008684f
C289 B.n183 VSUBS 0.008684f
C290 B.n184 VSUBS 0.008684f
C291 B.n185 VSUBS 0.008684f
C292 B.n186 VSUBS 0.008684f
C293 B.n187 VSUBS 0.008684f
C294 B.n188 VSUBS 0.008684f
C295 B.n189 VSUBS 0.008684f
C296 B.n190 VSUBS 0.008684f
C297 B.n191 VSUBS 0.008684f
C298 B.n192 VSUBS 0.008684f
C299 B.n193 VSUBS 0.01873f
C300 B.n194 VSUBS 0.008684f
C301 B.n195 VSUBS 0.008684f
C302 B.n196 VSUBS 0.008684f
C303 B.n197 VSUBS 0.008684f
C304 B.n198 VSUBS 0.008684f
C305 B.n199 VSUBS 0.008684f
C306 B.n200 VSUBS 0.008684f
C307 B.n201 VSUBS 0.008684f
C308 B.n202 VSUBS 0.008684f
C309 B.n203 VSUBS 0.008684f
C310 B.n204 VSUBS 0.008684f
C311 B.n205 VSUBS 0.008684f
C312 B.n206 VSUBS 0.008684f
C313 B.n207 VSUBS 0.008684f
C314 B.n208 VSUBS 0.008684f
C315 B.n209 VSUBS 0.008684f
C316 B.n210 VSUBS 0.008684f
C317 B.n211 VSUBS 0.008684f
C318 B.n212 VSUBS 0.008684f
C319 B.n213 VSUBS 0.008684f
C320 B.n214 VSUBS 0.008684f
C321 B.n215 VSUBS 0.008684f
C322 B.n216 VSUBS 0.008684f
C323 B.n217 VSUBS 0.008684f
C324 B.n218 VSUBS 0.008684f
C325 B.n219 VSUBS 0.008684f
C326 B.n220 VSUBS 0.008684f
C327 B.n221 VSUBS 0.008684f
C328 B.n222 VSUBS 0.008684f
C329 B.n223 VSUBS 0.008684f
C330 B.n224 VSUBS 0.008684f
C331 B.n225 VSUBS 0.008684f
C332 B.n226 VSUBS 0.008684f
C333 B.n227 VSUBS 0.008684f
C334 B.n228 VSUBS 0.008684f
C335 B.n229 VSUBS 0.008684f
C336 B.n230 VSUBS 0.008684f
C337 B.n231 VSUBS 0.008684f
C338 B.n232 VSUBS 0.008684f
C339 B.n233 VSUBS 0.008684f
C340 B.n234 VSUBS 0.008684f
C341 B.n235 VSUBS 0.008684f
C342 B.n236 VSUBS 0.008684f
C343 B.n237 VSUBS 0.008684f
C344 B.n238 VSUBS 0.008684f
C345 B.n239 VSUBS 0.008684f
C346 B.n240 VSUBS 0.008684f
C347 B.n241 VSUBS 0.008684f
C348 B.n242 VSUBS 0.008684f
C349 B.n243 VSUBS 0.008684f
C350 B.n244 VSUBS 0.008684f
C351 B.n245 VSUBS 0.008684f
C352 B.n246 VSUBS 0.008684f
C353 B.n247 VSUBS 0.008684f
C354 B.n248 VSUBS 0.008684f
C355 B.n249 VSUBS 0.008684f
C356 B.n250 VSUBS 0.01873f
C357 B.n251 VSUBS 0.01958f
C358 B.n252 VSUBS 0.01958f
C359 B.n253 VSUBS 0.008684f
C360 B.n254 VSUBS 0.008684f
C361 B.n255 VSUBS 0.008684f
C362 B.n256 VSUBS 0.008684f
C363 B.n257 VSUBS 0.008684f
C364 B.n258 VSUBS 0.008684f
C365 B.n259 VSUBS 0.008684f
C366 B.n260 VSUBS 0.008684f
C367 B.n261 VSUBS 0.008684f
C368 B.n262 VSUBS 0.008684f
C369 B.n263 VSUBS 0.008684f
C370 B.n264 VSUBS 0.008684f
C371 B.n265 VSUBS 0.008684f
C372 B.n266 VSUBS 0.008684f
C373 B.n267 VSUBS 0.008684f
C374 B.n268 VSUBS 0.008684f
C375 B.n269 VSUBS 0.008684f
C376 B.n270 VSUBS 0.008684f
C377 B.n271 VSUBS 0.008684f
C378 B.n272 VSUBS 0.008684f
C379 B.n273 VSUBS 0.008684f
C380 B.n274 VSUBS 0.008684f
C381 B.n275 VSUBS 0.008684f
C382 B.n276 VSUBS 0.008684f
C383 B.n277 VSUBS 0.008684f
C384 B.n278 VSUBS 0.008684f
C385 B.n279 VSUBS 0.008684f
C386 B.n280 VSUBS 0.008684f
C387 B.n281 VSUBS 0.008684f
C388 B.n282 VSUBS 0.008684f
C389 B.n283 VSUBS 0.008684f
C390 B.n284 VSUBS 0.008684f
C391 B.n285 VSUBS 0.008684f
C392 B.n286 VSUBS 0.008684f
C393 B.n287 VSUBS 0.008684f
C394 B.n288 VSUBS 0.008684f
C395 B.n289 VSUBS 0.008684f
C396 B.n290 VSUBS 0.008684f
C397 B.n291 VSUBS 0.008684f
C398 B.n292 VSUBS 0.008684f
C399 B.n293 VSUBS 0.008684f
C400 B.n294 VSUBS 0.008684f
C401 B.n295 VSUBS 0.008684f
C402 B.n296 VSUBS 0.008684f
C403 B.n297 VSUBS 0.008684f
C404 B.n298 VSUBS 0.008684f
C405 B.n299 VSUBS 0.008684f
C406 B.n300 VSUBS 0.008684f
C407 B.n301 VSUBS 0.008684f
C408 B.n302 VSUBS 0.008684f
C409 B.n303 VSUBS 0.008684f
C410 B.n304 VSUBS 0.008684f
C411 B.n305 VSUBS 0.008684f
C412 B.n306 VSUBS 0.008684f
C413 B.n307 VSUBS 0.008684f
C414 B.n308 VSUBS 0.008684f
C415 B.n309 VSUBS 0.008684f
C416 B.n310 VSUBS 0.008684f
C417 B.n311 VSUBS 0.008684f
C418 B.n312 VSUBS 0.008684f
C419 B.n313 VSUBS 0.008684f
C420 B.n314 VSUBS 0.008684f
C421 B.n315 VSUBS 0.008684f
C422 B.n316 VSUBS 0.008684f
C423 B.n317 VSUBS 0.008684f
C424 B.n318 VSUBS 0.008684f
C425 B.n319 VSUBS 0.008684f
C426 B.n320 VSUBS 0.008684f
C427 B.n321 VSUBS 0.008684f
C428 B.n322 VSUBS 0.008684f
C429 B.n323 VSUBS 0.008684f
C430 B.n324 VSUBS 0.008684f
C431 B.n325 VSUBS 0.008684f
C432 B.n326 VSUBS 0.008684f
C433 B.n327 VSUBS 0.008684f
C434 B.n328 VSUBS 0.008684f
C435 B.n329 VSUBS 0.008684f
C436 B.n330 VSUBS 0.008684f
C437 B.n331 VSUBS 0.008684f
C438 B.n332 VSUBS 0.008684f
C439 B.n333 VSUBS 0.008684f
C440 B.n334 VSUBS 0.008684f
C441 B.n335 VSUBS 0.008684f
C442 B.n336 VSUBS 0.008684f
C443 B.n337 VSUBS 0.008684f
C444 B.n338 VSUBS 0.008684f
C445 B.n339 VSUBS 0.008684f
C446 B.n340 VSUBS 0.008684f
C447 B.n341 VSUBS 0.008684f
C448 B.n342 VSUBS 0.008684f
C449 B.n343 VSUBS 0.008684f
C450 B.n344 VSUBS 0.008173f
C451 B.n345 VSUBS 0.008684f
C452 B.n346 VSUBS 0.008684f
C453 B.n347 VSUBS 0.004853f
C454 B.n348 VSUBS 0.008684f
C455 B.n349 VSUBS 0.008684f
C456 B.n350 VSUBS 0.008684f
C457 B.n351 VSUBS 0.008684f
C458 B.n352 VSUBS 0.008684f
C459 B.n353 VSUBS 0.008684f
C460 B.n354 VSUBS 0.008684f
C461 B.n355 VSUBS 0.008684f
C462 B.n356 VSUBS 0.008684f
C463 B.n357 VSUBS 0.008684f
C464 B.n358 VSUBS 0.008684f
C465 B.n359 VSUBS 0.008684f
C466 B.n360 VSUBS 0.004853f
C467 B.n361 VSUBS 0.020119f
C468 B.n362 VSUBS 0.008173f
C469 B.n363 VSUBS 0.008684f
C470 B.n364 VSUBS 0.008684f
C471 B.n365 VSUBS 0.008684f
C472 B.n366 VSUBS 0.008684f
C473 B.n367 VSUBS 0.008684f
C474 B.n368 VSUBS 0.008684f
C475 B.n369 VSUBS 0.008684f
C476 B.n370 VSUBS 0.008684f
C477 B.n371 VSUBS 0.008684f
C478 B.n372 VSUBS 0.008684f
C479 B.n373 VSUBS 0.008684f
C480 B.n374 VSUBS 0.008684f
C481 B.n375 VSUBS 0.008684f
C482 B.n376 VSUBS 0.008684f
C483 B.n377 VSUBS 0.008684f
C484 B.n378 VSUBS 0.008684f
C485 B.n379 VSUBS 0.008684f
C486 B.n380 VSUBS 0.008684f
C487 B.n381 VSUBS 0.008684f
C488 B.n382 VSUBS 0.008684f
C489 B.n383 VSUBS 0.008684f
C490 B.n384 VSUBS 0.008684f
C491 B.n385 VSUBS 0.008684f
C492 B.n386 VSUBS 0.008684f
C493 B.n387 VSUBS 0.008684f
C494 B.n388 VSUBS 0.008684f
C495 B.n389 VSUBS 0.008684f
C496 B.n390 VSUBS 0.008684f
C497 B.n391 VSUBS 0.008684f
C498 B.n392 VSUBS 0.008684f
C499 B.n393 VSUBS 0.008684f
C500 B.n394 VSUBS 0.008684f
C501 B.n395 VSUBS 0.008684f
C502 B.n396 VSUBS 0.008684f
C503 B.n397 VSUBS 0.008684f
C504 B.n398 VSUBS 0.008684f
C505 B.n399 VSUBS 0.008684f
C506 B.n400 VSUBS 0.008684f
C507 B.n401 VSUBS 0.008684f
C508 B.n402 VSUBS 0.008684f
C509 B.n403 VSUBS 0.008684f
C510 B.n404 VSUBS 0.008684f
C511 B.n405 VSUBS 0.008684f
C512 B.n406 VSUBS 0.008684f
C513 B.n407 VSUBS 0.008684f
C514 B.n408 VSUBS 0.008684f
C515 B.n409 VSUBS 0.008684f
C516 B.n410 VSUBS 0.008684f
C517 B.n411 VSUBS 0.008684f
C518 B.n412 VSUBS 0.008684f
C519 B.n413 VSUBS 0.008684f
C520 B.n414 VSUBS 0.008684f
C521 B.n415 VSUBS 0.008684f
C522 B.n416 VSUBS 0.008684f
C523 B.n417 VSUBS 0.008684f
C524 B.n418 VSUBS 0.008684f
C525 B.n419 VSUBS 0.008684f
C526 B.n420 VSUBS 0.008684f
C527 B.n421 VSUBS 0.008684f
C528 B.n422 VSUBS 0.008684f
C529 B.n423 VSUBS 0.008684f
C530 B.n424 VSUBS 0.008684f
C531 B.n425 VSUBS 0.008684f
C532 B.n426 VSUBS 0.008684f
C533 B.n427 VSUBS 0.008684f
C534 B.n428 VSUBS 0.008684f
C535 B.n429 VSUBS 0.008684f
C536 B.n430 VSUBS 0.008684f
C537 B.n431 VSUBS 0.008684f
C538 B.n432 VSUBS 0.008684f
C539 B.n433 VSUBS 0.008684f
C540 B.n434 VSUBS 0.008684f
C541 B.n435 VSUBS 0.008684f
C542 B.n436 VSUBS 0.008684f
C543 B.n437 VSUBS 0.008684f
C544 B.n438 VSUBS 0.008684f
C545 B.n439 VSUBS 0.008684f
C546 B.n440 VSUBS 0.008684f
C547 B.n441 VSUBS 0.008684f
C548 B.n442 VSUBS 0.008684f
C549 B.n443 VSUBS 0.008684f
C550 B.n444 VSUBS 0.008684f
C551 B.n445 VSUBS 0.008684f
C552 B.n446 VSUBS 0.008684f
C553 B.n447 VSUBS 0.008684f
C554 B.n448 VSUBS 0.008684f
C555 B.n449 VSUBS 0.008684f
C556 B.n450 VSUBS 0.008684f
C557 B.n451 VSUBS 0.008684f
C558 B.n452 VSUBS 0.008684f
C559 B.n453 VSUBS 0.008684f
C560 B.n454 VSUBS 0.008684f
C561 B.n455 VSUBS 0.01958f
C562 B.n456 VSUBS 0.01958f
C563 B.n457 VSUBS 0.01873f
C564 B.n458 VSUBS 0.008684f
C565 B.n459 VSUBS 0.008684f
C566 B.n460 VSUBS 0.008684f
C567 B.n461 VSUBS 0.008684f
C568 B.n462 VSUBS 0.008684f
C569 B.n463 VSUBS 0.008684f
C570 B.n464 VSUBS 0.008684f
C571 B.n465 VSUBS 0.008684f
C572 B.n466 VSUBS 0.008684f
C573 B.n467 VSUBS 0.008684f
C574 B.n468 VSUBS 0.008684f
C575 B.n469 VSUBS 0.008684f
C576 B.n470 VSUBS 0.008684f
C577 B.n471 VSUBS 0.008684f
C578 B.n472 VSUBS 0.008684f
C579 B.n473 VSUBS 0.008684f
C580 B.n474 VSUBS 0.008684f
C581 B.n475 VSUBS 0.008684f
C582 B.n476 VSUBS 0.008684f
C583 B.n477 VSUBS 0.008684f
C584 B.n478 VSUBS 0.008684f
C585 B.n479 VSUBS 0.008684f
C586 B.n480 VSUBS 0.008684f
C587 B.n481 VSUBS 0.008684f
C588 B.n482 VSUBS 0.008684f
C589 B.n483 VSUBS 0.008684f
C590 B.n484 VSUBS 0.008684f
C591 B.n485 VSUBS 0.008684f
C592 B.n486 VSUBS 0.008684f
C593 B.n487 VSUBS 0.008684f
C594 B.n488 VSUBS 0.008684f
C595 B.n489 VSUBS 0.008684f
C596 B.n490 VSUBS 0.008684f
C597 B.n491 VSUBS 0.008684f
C598 B.n492 VSUBS 0.008684f
C599 B.n493 VSUBS 0.008684f
C600 B.n494 VSUBS 0.008684f
C601 B.n495 VSUBS 0.008684f
C602 B.n496 VSUBS 0.008684f
C603 B.n497 VSUBS 0.008684f
C604 B.n498 VSUBS 0.008684f
C605 B.n499 VSUBS 0.008684f
C606 B.n500 VSUBS 0.008684f
C607 B.n501 VSUBS 0.008684f
C608 B.n502 VSUBS 0.008684f
C609 B.n503 VSUBS 0.008684f
C610 B.n504 VSUBS 0.008684f
C611 B.n505 VSUBS 0.008684f
C612 B.n506 VSUBS 0.008684f
C613 B.n507 VSUBS 0.008684f
C614 B.n508 VSUBS 0.008684f
C615 B.n509 VSUBS 0.008684f
C616 B.n510 VSUBS 0.008684f
C617 B.n511 VSUBS 0.008684f
C618 B.n512 VSUBS 0.008684f
C619 B.n513 VSUBS 0.008684f
C620 B.n514 VSUBS 0.008684f
C621 B.n515 VSUBS 0.008684f
C622 B.n516 VSUBS 0.008684f
C623 B.n517 VSUBS 0.008684f
C624 B.n518 VSUBS 0.008684f
C625 B.n519 VSUBS 0.008684f
C626 B.n520 VSUBS 0.008684f
C627 B.n521 VSUBS 0.008684f
C628 B.n522 VSUBS 0.008684f
C629 B.n523 VSUBS 0.008684f
C630 B.n524 VSUBS 0.008684f
C631 B.n525 VSUBS 0.008684f
C632 B.n526 VSUBS 0.008684f
C633 B.n527 VSUBS 0.008684f
C634 B.n528 VSUBS 0.008684f
C635 B.n529 VSUBS 0.008684f
C636 B.n530 VSUBS 0.008684f
C637 B.n531 VSUBS 0.008684f
C638 B.n532 VSUBS 0.008684f
C639 B.n533 VSUBS 0.008684f
C640 B.n534 VSUBS 0.008684f
C641 B.n535 VSUBS 0.008684f
C642 B.n536 VSUBS 0.008684f
C643 B.n537 VSUBS 0.008684f
C644 B.n538 VSUBS 0.008684f
C645 B.n539 VSUBS 0.008684f
C646 B.n540 VSUBS 0.008684f
C647 B.n541 VSUBS 0.008684f
C648 B.n542 VSUBS 0.008684f
C649 B.n543 VSUBS 0.008684f
C650 B.n544 VSUBS 0.008684f
C651 B.n545 VSUBS 0.008684f
C652 B.n546 VSUBS 0.008684f
C653 B.n547 VSUBS 0.019854f
C654 B.n548 VSUBS 0.018456f
C655 B.n549 VSUBS 0.01958f
C656 B.n550 VSUBS 0.008684f
C657 B.n551 VSUBS 0.008684f
C658 B.n552 VSUBS 0.008684f
C659 B.n553 VSUBS 0.008684f
C660 B.n554 VSUBS 0.008684f
C661 B.n555 VSUBS 0.008684f
C662 B.n556 VSUBS 0.008684f
C663 B.n557 VSUBS 0.008684f
C664 B.n558 VSUBS 0.008684f
C665 B.n559 VSUBS 0.008684f
C666 B.n560 VSUBS 0.008684f
C667 B.n561 VSUBS 0.008684f
C668 B.n562 VSUBS 0.008684f
C669 B.n563 VSUBS 0.008684f
C670 B.n564 VSUBS 0.008684f
C671 B.n565 VSUBS 0.008684f
C672 B.n566 VSUBS 0.008684f
C673 B.n567 VSUBS 0.008684f
C674 B.n568 VSUBS 0.008684f
C675 B.n569 VSUBS 0.008684f
C676 B.n570 VSUBS 0.008684f
C677 B.n571 VSUBS 0.008684f
C678 B.n572 VSUBS 0.008684f
C679 B.n573 VSUBS 0.008684f
C680 B.n574 VSUBS 0.008684f
C681 B.n575 VSUBS 0.008684f
C682 B.n576 VSUBS 0.008684f
C683 B.n577 VSUBS 0.008684f
C684 B.n578 VSUBS 0.008684f
C685 B.n579 VSUBS 0.008684f
C686 B.n580 VSUBS 0.008684f
C687 B.n581 VSUBS 0.008684f
C688 B.n582 VSUBS 0.008684f
C689 B.n583 VSUBS 0.008684f
C690 B.n584 VSUBS 0.008684f
C691 B.n585 VSUBS 0.008684f
C692 B.n586 VSUBS 0.008684f
C693 B.n587 VSUBS 0.008684f
C694 B.n588 VSUBS 0.008684f
C695 B.n589 VSUBS 0.008684f
C696 B.n590 VSUBS 0.008684f
C697 B.n591 VSUBS 0.008684f
C698 B.n592 VSUBS 0.008684f
C699 B.n593 VSUBS 0.008684f
C700 B.n594 VSUBS 0.008684f
C701 B.n595 VSUBS 0.008684f
C702 B.n596 VSUBS 0.008684f
C703 B.n597 VSUBS 0.008684f
C704 B.n598 VSUBS 0.008684f
C705 B.n599 VSUBS 0.008684f
C706 B.n600 VSUBS 0.008684f
C707 B.n601 VSUBS 0.008684f
C708 B.n602 VSUBS 0.008684f
C709 B.n603 VSUBS 0.008684f
C710 B.n604 VSUBS 0.008684f
C711 B.n605 VSUBS 0.008684f
C712 B.n606 VSUBS 0.008684f
C713 B.n607 VSUBS 0.008684f
C714 B.n608 VSUBS 0.008684f
C715 B.n609 VSUBS 0.008684f
C716 B.n610 VSUBS 0.008684f
C717 B.n611 VSUBS 0.008684f
C718 B.n612 VSUBS 0.008684f
C719 B.n613 VSUBS 0.008684f
C720 B.n614 VSUBS 0.008684f
C721 B.n615 VSUBS 0.008684f
C722 B.n616 VSUBS 0.008684f
C723 B.n617 VSUBS 0.008684f
C724 B.n618 VSUBS 0.008684f
C725 B.n619 VSUBS 0.008684f
C726 B.n620 VSUBS 0.008684f
C727 B.n621 VSUBS 0.008684f
C728 B.n622 VSUBS 0.008684f
C729 B.n623 VSUBS 0.008684f
C730 B.n624 VSUBS 0.008684f
C731 B.n625 VSUBS 0.008684f
C732 B.n626 VSUBS 0.008684f
C733 B.n627 VSUBS 0.008684f
C734 B.n628 VSUBS 0.008684f
C735 B.n629 VSUBS 0.008684f
C736 B.n630 VSUBS 0.008684f
C737 B.n631 VSUBS 0.008684f
C738 B.n632 VSUBS 0.008684f
C739 B.n633 VSUBS 0.008684f
C740 B.n634 VSUBS 0.008684f
C741 B.n635 VSUBS 0.008684f
C742 B.n636 VSUBS 0.008684f
C743 B.n637 VSUBS 0.008684f
C744 B.n638 VSUBS 0.008684f
C745 B.n639 VSUBS 0.008684f
C746 B.n640 VSUBS 0.008684f
C747 B.n641 VSUBS 0.008684f
C748 B.n642 VSUBS 0.008173f
C749 B.n643 VSUBS 0.020119f
C750 B.n644 VSUBS 0.004853f
C751 B.n645 VSUBS 0.008684f
C752 B.n646 VSUBS 0.008684f
C753 B.n647 VSUBS 0.008684f
C754 B.n648 VSUBS 0.008684f
C755 B.n649 VSUBS 0.008684f
C756 B.n650 VSUBS 0.008684f
C757 B.n651 VSUBS 0.008684f
C758 B.n652 VSUBS 0.008684f
C759 B.n653 VSUBS 0.008684f
C760 B.n654 VSUBS 0.008684f
C761 B.n655 VSUBS 0.008684f
C762 B.n656 VSUBS 0.008684f
C763 B.n657 VSUBS 0.004853f
C764 B.n658 VSUBS 0.008684f
C765 B.n659 VSUBS 0.008684f
C766 B.n660 VSUBS 0.008684f
C767 B.n661 VSUBS 0.008684f
C768 B.n662 VSUBS 0.008684f
C769 B.n663 VSUBS 0.008684f
C770 B.n664 VSUBS 0.008684f
C771 B.n665 VSUBS 0.008684f
C772 B.n666 VSUBS 0.008684f
C773 B.n667 VSUBS 0.008684f
C774 B.n668 VSUBS 0.008684f
C775 B.n669 VSUBS 0.008684f
C776 B.n670 VSUBS 0.008684f
C777 B.n671 VSUBS 0.008684f
C778 B.n672 VSUBS 0.008684f
C779 B.n673 VSUBS 0.008684f
C780 B.n674 VSUBS 0.008684f
C781 B.n675 VSUBS 0.008684f
C782 B.n676 VSUBS 0.008684f
C783 B.n677 VSUBS 0.008684f
C784 B.n678 VSUBS 0.008684f
C785 B.n679 VSUBS 0.008684f
C786 B.n680 VSUBS 0.008684f
C787 B.n681 VSUBS 0.008684f
C788 B.n682 VSUBS 0.008684f
C789 B.n683 VSUBS 0.008684f
C790 B.n684 VSUBS 0.008684f
C791 B.n685 VSUBS 0.008684f
C792 B.n686 VSUBS 0.008684f
C793 B.n687 VSUBS 0.008684f
C794 B.n688 VSUBS 0.008684f
C795 B.n689 VSUBS 0.008684f
C796 B.n690 VSUBS 0.008684f
C797 B.n691 VSUBS 0.008684f
C798 B.n692 VSUBS 0.008684f
C799 B.n693 VSUBS 0.008684f
C800 B.n694 VSUBS 0.008684f
C801 B.n695 VSUBS 0.008684f
C802 B.n696 VSUBS 0.008684f
C803 B.n697 VSUBS 0.008684f
C804 B.n698 VSUBS 0.008684f
C805 B.n699 VSUBS 0.008684f
C806 B.n700 VSUBS 0.008684f
C807 B.n701 VSUBS 0.008684f
C808 B.n702 VSUBS 0.008684f
C809 B.n703 VSUBS 0.008684f
C810 B.n704 VSUBS 0.008684f
C811 B.n705 VSUBS 0.008684f
C812 B.n706 VSUBS 0.008684f
C813 B.n707 VSUBS 0.008684f
C814 B.n708 VSUBS 0.008684f
C815 B.n709 VSUBS 0.008684f
C816 B.n710 VSUBS 0.008684f
C817 B.n711 VSUBS 0.008684f
C818 B.n712 VSUBS 0.008684f
C819 B.n713 VSUBS 0.008684f
C820 B.n714 VSUBS 0.008684f
C821 B.n715 VSUBS 0.008684f
C822 B.n716 VSUBS 0.008684f
C823 B.n717 VSUBS 0.008684f
C824 B.n718 VSUBS 0.008684f
C825 B.n719 VSUBS 0.008684f
C826 B.n720 VSUBS 0.008684f
C827 B.n721 VSUBS 0.008684f
C828 B.n722 VSUBS 0.008684f
C829 B.n723 VSUBS 0.008684f
C830 B.n724 VSUBS 0.008684f
C831 B.n725 VSUBS 0.008684f
C832 B.n726 VSUBS 0.008684f
C833 B.n727 VSUBS 0.008684f
C834 B.n728 VSUBS 0.008684f
C835 B.n729 VSUBS 0.008684f
C836 B.n730 VSUBS 0.008684f
C837 B.n731 VSUBS 0.008684f
C838 B.n732 VSUBS 0.008684f
C839 B.n733 VSUBS 0.008684f
C840 B.n734 VSUBS 0.008684f
C841 B.n735 VSUBS 0.008684f
C842 B.n736 VSUBS 0.008684f
C843 B.n737 VSUBS 0.008684f
C844 B.n738 VSUBS 0.008684f
C845 B.n739 VSUBS 0.008684f
C846 B.n740 VSUBS 0.008684f
C847 B.n741 VSUBS 0.008684f
C848 B.n742 VSUBS 0.008684f
C849 B.n743 VSUBS 0.008684f
C850 B.n744 VSUBS 0.008684f
C851 B.n745 VSUBS 0.008684f
C852 B.n746 VSUBS 0.008684f
C853 B.n747 VSUBS 0.008684f
C854 B.n748 VSUBS 0.008684f
C855 B.n749 VSUBS 0.008684f
C856 B.n750 VSUBS 0.008684f
C857 B.n751 VSUBS 0.008684f
C858 B.n752 VSUBS 0.01958f
C859 B.n753 VSUBS 0.01873f
C860 B.n754 VSUBS 0.01873f
C861 B.n755 VSUBS 0.008684f
C862 B.n756 VSUBS 0.008684f
C863 B.n757 VSUBS 0.008684f
C864 B.n758 VSUBS 0.008684f
C865 B.n759 VSUBS 0.008684f
C866 B.n760 VSUBS 0.008684f
C867 B.n761 VSUBS 0.008684f
C868 B.n762 VSUBS 0.008684f
C869 B.n763 VSUBS 0.008684f
C870 B.n764 VSUBS 0.008684f
C871 B.n765 VSUBS 0.008684f
C872 B.n766 VSUBS 0.008684f
C873 B.n767 VSUBS 0.008684f
C874 B.n768 VSUBS 0.008684f
C875 B.n769 VSUBS 0.008684f
C876 B.n770 VSUBS 0.008684f
C877 B.n771 VSUBS 0.008684f
C878 B.n772 VSUBS 0.008684f
C879 B.n773 VSUBS 0.008684f
C880 B.n774 VSUBS 0.008684f
C881 B.n775 VSUBS 0.008684f
C882 B.n776 VSUBS 0.008684f
C883 B.n777 VSUBS 0.008684f
C884 B.n778 VSUBS 0.008684f
C885 B.n779 VSUBS 0.008684f
C886 B.n780 VSUBS 0.008684f
C887 B.n781 VSUBS 0.008684f
C888 B.n782 VSUBS 0.008684f
C889 B.n783 VSUBS 0.008684f
C890 B.n784 VSUBS 0.008684f
C891 B.n785 VSUBS 0.008684f
C892 B.n786 VSUBS 0.008684f
C893 B.n787 VSUBS 0.008684f
C894 B.n788 VSUBS 0.008684f
C895 B.n789 VSUBS 0.008684f
C896 B.n790 VSUBS 0.008684f
C897 B.n791 VSUBS 0.008684f
C898 B.n792 VSUBS 0.008684f
C899 B.n793 VSUBS 0.008684f
C900 B.n794 VSUBS 0.008684f
C901 B.n795 VSUBS 0.008684f
C902 B.n796 VSUBS 0.008684f
C903 B.n797 VSUBS 0.008684f
C904 B.n798 VSUBS 0.008684f
C905 B.n799 VSUBS 0.019663f
C906 VDD1.t4 VSUBS 4.53655f
C907 VDD1.t1 VSUBS 0.416748f
C908 VDD1.t3 VSUBS 0.416748f
C909 VDD1.n0 VSUBS 3.49005f
C910 VDD1.n1 VSUBS 1.4057f
C911 VDD1.t5 VSUBS 4.53654f
C912 VDD1.t8 VSUBS 0.416748f
C913 VDD1.t6 VSUBS 0.416748f
C914 VDD1.n2 VSUBS 3.49005f
C915 VDD1.n3 VSUBS 1.39874f
C916 VDD1.t7 VSUBS 0.416748f
C917 VDD1.t9 VSUBS 0.416748f
C918 VDD1.n4 VSUBS 3.49772f
C919 VDD1.n5 VSUBS 3.09998f
C920 VDD1.t0 VSUBS 0.416748f
C921 VDD1.t2 VSUBS 0.416748f
C922 VDD1.n6 VSUBS 3.49003f
C923 VDD1.n7 VSUBS 3.6274f
C924 VTAIL.t18 VSUBS 0.419564f
C925 VTAIL.t4 VSUBS 0.419564f
C926 VTAIL.n0 VSUBS 3.33791f
C927 VTAIL.n1 VSUBS 0.85101f
C928 VTAIL.t11 VSUBS 4.3538f
C929 VTAIL.n2 VSUBS 0.997706f
C930 VTAIL.t15 VSUBS 0.419564f
C931 VTAIL.t10 VSUBS 0.419564f
C932 VTAIL.n3 VSUBS 3.33791f
C933 VTAIL.n4 VSUBS 0.874674f
C934 VTAIL.t17 VSUBS 0.419564f
C935 VTAIL.t9 VSUBS 0.419564f
C936 VTAIL.n5 VSUBS 3.33791f
C937 VTAIL.n6 VSUBS 2.8167f
C938 VTAIL.t0 VSUBS 0.419564f
C939 VTAIL.t6 VSUBS 0.419564f
C940 VTAIL.n7 VSUBS 3.33791f
C941 VTAIL.n8 VSUBS 2.8167f
C942 VTAIL.t2 VSUBS 0.419564f
C943 VTAIL.t7 VSUBS 0.419564f
C944 VTAIL.n9 VSUBS 3.33791f
C945 VTAIL.n10 VSUBS 0.874675f
C946 VTAIL.t5 VSUBS 4.3538f
C947 VTAIL.n11 VSUBS 0.997698f
C948 VTAIL.t8 VSUBS 0.419564f
C949 VTAIL.t13 VSUBS 0.419564f
C950 VTAIL.n12 VSUBS 3.33791f
C951 VTAIL.n13 VSUBS 0.869331f
C952 VTAIL.t16 VSUBS 0.419564f
C953 VTAIL.t12 VSUBS 0.419564f
C954 VTAIL.n14 VSUBS 3.33791f
C955 VTAIL.n15 VSUBS 0.874675f
C956 VTAIL.t14 VSUBS 4.3538f
C957 VTAIL.n16 VSUBS 2.85118f
C958 VTAIL.t1 VSUBS 4.3538f
C959 VTAIL.n17 VSUBS 2.85118f
C960 VTAIL.t19 VSUBS 0.419564f
C961 VTAIL.t3 VSUBS 0.419564f
C962 VTAIL.n18 VSUBS 3.33791f
C963 VTAIL.n19 VSUBS 0.7991f
C964 VP.n0 VSUBS 0.044794f
C965 VP.t2 VSUBS 2.14513f
C966 VP.n1 VSUBS 0.768604f
C967 VP.n2 VSUBS 0.044794f
C968 VP.t3 VSUBS 2.14513f
C969 VP.n3 VSUBS 0.044346f
C970 VP.n4 VSUBS 0.044794f
C971 VP.t1 VSUBS 2.14513f
C972 VP.t4 VSUBS 2.20651f
C973 VP.n5 VSUBS 0.815165f
C974 VP.n6 VSUBS 0.044794f
C975 VP.t7 VSUBS 2.20651f
C976 VP.t9 VSUBS 2.14513f
C977 VP.n7 VSUBS 0.768604f
C978 VP.n8 VSUBS 0.044794f
C979 VP.t6 VSUBS 2.14513f
C980 VP.n9 VSUBS 0.044346f
C981 VP.t5 VSUBS 2.22941f
C982 VP.n10 VSUBS 0.824529f
C983 VP.t8 VSUBS 2.14513f
C984 VP.n11 VSUBS 0.808985f
C985 VP.n12 VSUBS 0.058341f
C986 VP.n13 VSUBS 0.187101f
C987 VP.n14 VSUBS 0.044794f
C988 VP.n15 VSUBS 0.044794f
C989 VP.n16 VSUBS 0.82146f
C990 VP.n17 VSUBS 0.044346f
C991 VP.n18 VSUBS 0.058341f
C992 VP.n19 VSUBS 0.044794f
C993 VP.n20 VSUBS 0.044794f
C994 VP.n21 VSUBS 0.0578f
C995 VP.n22 VSUBS 0.013923f
C996 VP.n23 VSUBS 0.815165f
C997 VP.n24 VSUBS 2.39064f
C998 VP.n25 VSUBS 2.42334f
C999 VP.n26 VSUBS 0.044794f
C1000 VP.n27 VSUBS 0.013923f
C1001 VP.n28 VSUBS 0.0578f
C1002 VP.n29 VSUBS 0.768604f
C1003 VP.n30 VSUBS 0.058341f
C1004 VP.n31 VSUBS 0.044794f
C1005 VP.n32 VSUBS 0.044794f
C1006 VP.n33 VSUBS 0.044794f
C1007 VP.n34 VSUBS 0.82146f
C1008 VP.n35 VSUBS 0.044346f
C1009 VP.n36 VSUBS 0.058341f
C1010 VP.n37 VSUBS 0.044794f
C1011 VP.n38 VSUBS 0.044794f
C1012 VP.n39 VSUBS 0.0578f
C1013 VP.n40 VSUBS 0.013923f
C1014 VP.t0 VSUBS 2.20651f
C1015 VP.n41 VSUBS 0.815165f
C1016 VP.n42 VSUBS 0.034714f
.ends

