* NGSPICE file created from diff_pair_sample_0938.ext - technology: sky130A

.subckt diff_pair_sample_0938 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=6.4623 ps=33.92 w=16.57 l=0.36
X1 VTAIL.t2 VN.t0 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=2.73405 ps=16.9 w=16.57 l=0.36
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=0.36
X3 VDD1.t4 VP.t1 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=6.4623 ps=33.92 w=16.57 l=0.36
X4 VDD1.t3 VP.t2 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=2.73405 ps=16.9 w=16.57 l=0.36
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=0.36
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=0.36
X7 VDD2.t4 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=2.73405 ps=16.9 w=16.57 l=0.36
X8 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=2.73405 ps=16.9 w=16.57 l=0.36
X9 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=6.4623 ps=33.92 w=16.57 l=0.36
X10 VTAIL.t9 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=2.73405 ps=16.9 w=16.57 l=0.36
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=0 ps=0 w=16.57 l=0.36
X12 VTAIL.t11 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=2.73405 ps=16.9 w=16.57 l=0.36
X13 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=6.4623 ps=33.92 w=16.57 l=0.36
X14 VDD1.t0 VP.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=6.4623 pd=33.92 as=2.73405 ps=16.9 w=16.57 l=0.36
X15 VTAIL.t1 VN.t5 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.73405 pd=16.9 as=2.73405 ps=16.9 w=16.57 l=0.36
R0 VP.n1 VP.t2 1240.95
R1 VP.n8 VP.t1 1220.52
R2 VP.n6 VP.t5 1220.52
R3 VP.n3 VP.t0 1220.52
R4 VP.n7 VP.t4 1219.06
R5 VP.n2 VP.t3 1219.06
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n7 VP.n0 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n4 VP.n1 70.6808
R11 VP.n7 VP.n6 46.7399
R12 VP.n8 VP.n7 46.7399
R13 VP.n3 VP.n2 46.7399
R14 VP.n5 VP.n4 43.3679
R15 VP.n2 VP.n1 20.4028
R16 VP.n5 VP.n0 0.189894
R17 VP.n9 VP.n0 0.189894
R18 VP VP.n9 0.0516364
R19 VTAIL.n7 VTAIL.t4 47.787
R20 VTAIL.n11 VTAIL.t0 47.7868
R21 VTAIL.n2 VTAIL.t6 47.7868
R22 VTAIL.n10 VTAIL.t7 47.7868
R23 VTAIL.n9 VTAIL.n8 46.5921
R24 VTAIL.n6 VTAIL.n5 46.5921
R25 VTAIL.n1 VTAIL.n0 46.5918
R26 VTAIL.n4 VTAIL.n3 46.5918
R27 VTAIL.n6 VTAIL.n4 27.841
R28 VTAIL.n11 VTAIL.n10 27.2462
R29 VTAIL.n0 VTAIL.t3 1.19543
R30 VTAIL.n0 VTAIL.t2 1.19543
R31 VTAIL.n3 VTAIL.t10 1.19543
R32 VTAIL.n3 VTAIL.t11 1.19543
R33 VTAIL.n8 VTAIL.t8 1.19543
R34 VTAIL.n8 VTAIL.t9 1.19543
R35 VTAIL.n5 VTAIL.t5 1.19543
R36 VTAIL.n5 VTAIL.t1 1.19543
R37 VTAIL.n9 VTAIL.n7 0.767741
R38 VTAIL.n2 VTAIL.n1 0.767741
R39 VTAIL.n7 VTAIL.n6 0.595328
R40 VTAIL.n10 VTAIL.n9 0.595328
R41 VTAIL.n4 VTAIL.n2 0.595328
R42 VTAIL VTAIL.n11 0.388431
R43 VTAIL VTAIL.n1 0.207397
R44 VDD1 VDD1.t3 64.9701
R45 VDD1.n1 VDD1.t0 64.8563
R46 VDD1.n1 VDD1.n0 63.364
R47 VDD1.n3 VDD1.n2 63.2707
R48 VDD1.n3 VDD1.n1 40.8134
R49 VDD1.n2 VDD1.t2 1.19543
R50 VDD1.n2 VDD1.t5 1.19543
R51 VDD1.n0 VDD1.t1 1.19543
R52 VDD1.n0 VDD1.t4 1.19543
R53 VDD1 VDD1.n3 0.0910172
R54 B.n392 B.t14 1320.36
R55 B.n401 B.t10 1320.36
R56 B.n96 B.t17 1320.36
R57 B.n94 B.t6 1320.36
R58 B.n740 B.n739 585
R59 B.n334 B.n93 585
R60 B.n333 B.n332 585
R61 B.n331 B.n330 585
R62 B.n329 B.n328 585
R63 B.n327 B.n326 585
R64 B.n325 B.n324 585
R65 B.n323 B.n322 585
R66 B.n321 B.n320 585
R67 B.n319 B.n318 585
R68 B.n317 B.n316 585
R69 B.n315 B.n314 585
R70 B.n313 B.n312 585
R71 B.n311 B.n310 585
R72 B.n309 B.n308 585
R73 B.n307 B.n306 585
R74 B.n305 B.n304 585
R75 B.n303 B.n302 585
R76 B.n301 B.n300 585
R77 B.n299 B.n298 585
R78 B.n297 B.n296 585
R79 B.n295 B.n294 585
R80 B.n293 B.n292 585
R81 B.n291 B.n290 585
R82 B.n289 B.n288 585
R83 B.n287 B.n286 585
R84 B.n285 B.n284 585
R85 B.n283 B.n282 585
R86 B.n281 B.n280 585
R87 B.n279 B.n278 585
R88 B.n277 B.n276 585
R89 B.n275 B.n274 585
R90 B.n273 B.n272 585
R91 B.n271 B.n270 585
R92 B.n269 B.n268 585
R93 B.n267 B.n266 585
R94 B.n265 B.n264 585
R95 B.n263 B.n262 585
R96 B.n261 B.n260 585
R97 B.n259 B.n258 585
R98 B.n257 B.n256 585
R99 B.n255 B.n254 585
R100 B.n253 B.n252 585
R101 B.n251 B.n250 585
R102 B.n249 B.n248 585
R103 B.n247 B.n246 585
R104 B.n245 B.n244 585
R105 B.n243 B.n242 585
R106 B.n241 B.n240 585
R107 B.n239 B.n238 585
R108 B.n237 B.n236 585
R109 B.n235 B.n234 585
R110 B.n233 B.n232 585
R111 B.n231 B.n230 585
R112 B.n229 B.n228 585
R113 B.n226 B.n225 585
R114 B.n224 B.n223 585
R115 B.n222 B.n221 585
R116 B.n220 B.n219 585
R117 B.n218 B.n217 585
R118 B.n216 B.n215 585
R119 B.n214 B.n213 585
R120 B.n212 B.n211 585
R121 B.n210 B.n209 585
R122 B.n208 B.n207 585
R123 B.n205 B.n204 585
R124 B.n203 B.n202 585
R125 B.n201 B.n200 585
R126 B.n199 B.n198 585
R127 B.n197 B.n196 585
R128 B.n195 B.n194 585
R129 B.n193 B.n192 585
R130 B.n191 B.n190 585
R131 B.n189 B.n188 585
R132 B.n187 B.n186 585
R133 B.n185 B.n184 585
R134 B.n183 B.n182 585
R135 B.n181 B.n180 585
R136 B.n179 B.n178 585
R137 B.n177 B.n176 585
R138 B.n175 B.n174 585
R139 B.n173 B.n172 585
R140 B.n171 B.n170 585
R141 B.n169 B.n168 585
R142 B.n167 B.n166 585
R143 B.n165 B.n164 585
R144 B.n163 B.n162 585
R145 B.n161 B.n160 585
R146 B.n159 B.n158 585
R147 B.n157 B.n156 585
R148 B.n155 B.n154 585
R149 B.n153 B.n152 585
R150 B.n151 B.n150 585
R151 B.n149 B.n148 585
R152 B.n147 B.n146 585
R153 B.n145 B.n144 585
R154 B.n143 B.n142 585
R155 B.n141 B.n140 585
R156 B.n139 B.n138 585
R157 B.n137 B.n136 585
R158 B.n135 B.n134 585
R159 B.n133 B.n132 585
R160 B.n131 B.n130 585
R161 B.n129 B.n128 585
R162 B.n127 B.n126 585
R163 B.n125 B.n124 585
R164 B.n123 B.n122 585
R165 B.n121 B.n120 585
R166 B.n119 B.n118 585
R167 B.n117 B.n116 585
R168 B.n115 B.n114 585
R169 B.n113 B.n112 585
R170 B.n111 B.n110 585
R171 B.n109 B.n108 585
R172 B.n107 B.n106 585
R173 B.n105 B.n104 585
R174 B.n103 B.n102 585
R175 B.n101 B.n100 585
R176 B.n99 B.n98 585
R177 B.n32 B.n31 585
R178 B.n738 B.n33 585
R179 B.n743 B.n33 585
R180 B.n737 B.n736 585
R181 B.n736 B.n29 585
R182 B.n735 B.n28 585
R183 B.n749 B.n28 585
R184 B.n734 B.n27 585
R185 B.n750 B.n27 585
R186 B.n733 B.n26 585
R187 B.n751 B.n26 585
R188 B.n732 B.n731 585
R189 B.n731 B.n22 585
R190 B.n730 B.n21 585
R191 B.n757 B.n21 585
R192 B.n729 B.n20 585
R193 B.n758 B.n20 585
R194 B.n728 B.n19 585
R195 B.n759 B.n19 585
R196 B.n727 B.n726 585
R197 B.n726 B.n18 585
R198 B.n725 B.n14 585
R199 B.n765 B.n14 585
R200 B.n724 B.n13 585
R201 B.n766 B.n13 585
R202 B.n723 B.n12 585
R203 B.n767 B.n12 585
R204 B.n722 B.n721 585
R205 B.n721 B.n11 585
R206 B.n720 B.n7 585
R207 B.n773 B.n7 585
R208 B.n719 B.n6 585
R209 B.n774 B.n6 585
R210 B.n718 B.n5 585
R211 B.n775 B.n5 585
R212 B.n717 B.n716 585
R213 B.n716 B.n4 585
R214 B.n715 B.n335 585
R215 B.n715 B.n714 585
R216 B.n704 B.n336 585
R217 B.n707 B.n336 585
R218 B.n706 B.n705 585
R219 B.n708 B.n706 585
R220 B.n703 B.n340 585
R221 B.n343 B.n340 585
R222 B.n702 B.n701 585
R223 B.n701 B.n700 585
R224 B.n342 B.n341 585
R225 B.n693 B.n342 585
R226 B.n692 B.n691 585
R227 B.n694 B.n692 585
R228 B.n690 B.n348 585
R229 B.n348 B.n347 585
R230 B.n689 B.n688 585
R231 B.n688 B.n687 585
R232 B.n350 B.n349 585
R233 B.n351 B.n350 585
R234 B.n680 B.n679 585
R235 B.n681 B.n680 585
R236 B.n678 B.n356 585
R237 B.n356 B.n355 585
R238 B.n677 B.n676 585
R239 B.n676 B.n675 585
R240 B.n358 B.n357 585
R241 B.n359 B.n358 585
R242 B.n668 B.n667 585
R243 B.n669 B.n668 585
R244 B.n362 B.n361 585
R245 B.n431 B.n430 585
R246 B.n432 B.n428 585
R247 B.n428 B.n363 585
R248 B.n434 B.n433 585
R249 B.n436 B.n427 585
R250 B.n439 B.n438 585
R251 B.n440 B.n426 585
R252 B.n442 B.n441 585
R253 B.n444 B.n425 585
R254 B.n447 B.n446 585
R255 B.n448 B.n424 585
R256 B.n450 B.n449 585
R257 B.n452 B.n423 585
R258 B.n455 B.n454 585
R259 B.n456 B.n422 585
R260 B.n458 B.n457 585
R261 B.n460 B.n421 585
R262 B.n463 B.n462 585
R263 B.n464 B.n420 585
R264 B.n466 B.n465 585
R265 B.n468 B.n419 585
R266 B.n471 B.n470 585
R267 B.n472 B.n418 585
R268 B.n474 B.n473 585
R269 B.n476 B.n417 585
R270 B.n479 B.n478 585
R271 B.n480 B.n416 585
R272 B.n482 B.n481 585
R273 B.n484 B.n415 585
R274 B.n487 B.n486 585
R275 B.n488 B.n414 585
R276 B.n490 B.n489 585
R277 B.n492 B.n413 585
R278 B.n495 B.n494 585
R279 B.n496 B.n412 585
R280 B.n498 B.n497 585
R281 B.n500 B.n411 585
R282 B.n503 B.n502 585
R283 B.n504 B.n410 585
R284 B.n506 B.n505 585
R285 B.n508 B.n409 585
R286 B.n511 B.n510 585
R287 B.n512 B.n408 585
R288 B.n514 B.n513 585
R289 B.n516 B.n407 585
R290 B.n519 B.n518 585
R291 B.n520 B.n406 585
R292 B.n522 B.n521 585
R293 B.n524 B.n405 585
R294 B.n527 B.n526 585
R295 B.n528 B.n404 585
R296 B.n530 B.n529 585
R297 B.n532 B.n403 585
R298 B.n535 B.n534 585
R299 B.n536 B.n400 585
R300 B.n539 B.n538 585
R301 B.n541 B.n399 585
R302 B.n544 B.n543 585
R303 B.n545 B.n398 585
R304 B.n547 B.n546 585
R305 B.n549 B.n397 585
R306 B.n552 B.n551 585
R307 B.n553 B.n396 585
R308 B.n555 B.n554 585
R309 B.n557 B.n395 585
R310 B.n560 B.n559 585
R311 B.n561 B.n391 585
R312 B.n563 B.n562 585
R313 B.n565 B.n390 585
R314 B.n568 B.n567 585
R315 B.n569 B.n389 585
R316 B.n571 B.n570 585
R317 B.n573 B.n388 585
R318 B.n576 B.n575 585
R319 B.n577 B.n387 585
R320 B.n579 B.n578 585
R321 B.n581 B.n386 585
R322 B.n584 B.n583 585
R323 B.n585 B.n385 585
R324 B.n587 B.n586 585
R325 B.n589 B.n384 585
R326 B.n592 B.n591 585
R327 B.n593 B.n383 585
R328 B.n595 B.n594 585
R329 B.n597 B.n382 585
R330 B.n600 B.n599 585
R331 B.n601 B.n381 585
R332 B.n603 B.n602 585
R333 B.n605 B.n380 585
R334 B.n608 B.n607 585
R335 B.n609 B.n379 585
R336 B.n611 B.n610 585
R337 B.n613 B.n378 585
R338 B.n616 B.n615 585
R339 B.n617 B.n377 585
R340 B.n619 B.n618 585
R341 B.n621 B.n376 585
R342 B.n624 B.n623 585
R343 B.n625 B.n375 585
R344 B.n627 B.n626 585
R345 B.n629 B.n374 585
R346 B.n632 B.n631 585
R347 B.n633 B.n373 585
R348 B.n635 B.n634 585
R349 B.n637 B.n372 585
R350 B.n640 B.n639 585
R351 B.n641 B.n371 585
R352 B.n643 B.n642 585
R353 B.n645 B.n370 585
R354 B.n648 B.n647 585
R355 B.n649 B.n369 585
R356 B.n651 B.n650 585
R357 B.n653 B.n368 585
R358 B.n656 B.n655 585
R359 B.n657 B.n367 585
R360 B.n659 B.n658 585
R361 B.n661 B.n366 585
R362 B.n662 B.n365 585
R363 B.n665 B.n664 585
R364 B.n666 B.n364 585
R365 B.n364 B.n363 585
R366 B.n671 B.n670 585
R367 B.n670 B.n669 585
R368 B.n672 B.n360 585
R369 B.n360 B.n359 585
R370 B.n674 B.n673 585
R371 B.n675 B.n674 585
R372 B.n354 B.n353 585
R373 B.n355 B.n354 585
R374 B.n683 B.n682 585
R375 B.n682 B.n681 585
R376 B.n684 B.n352 585
R377 B.n352 B.n351 585
R378 B.n686 B.n685 585
R379 B.n687 B.n686 585
R380 B.n346 B.n345 585
R381 B.n347 B.n346 585
R382 B.n696 B.n695 585
R383 B.n695 B.n694 585
R384 B.n697 B.n344 585
R385 B.n693 B.n344 585
R386 B.n699 B.n698 585
R387 B.n700 B.n699 585
R388 B.n339 B.n338 585
R389 B.n343 B.n339 585
R390 B.n710 B.n709 585
R391 B.n709 B.n708 585
R392 B.n711 B.n337 585
R393 B.n707 B.n337 585
R394 B.n713 B.n712 585
R395 B.n714 B.n713 585
R396 B.n2 B.n0 585
R397 B.n4 B.n2 585
R398 B.n3 B.n1 585
R399 B.n774 B.n3 585
R400 B.n772 B.n771 585
R401 B.n773 B.n772 585
R402 B.n770 B.n8 585
R403 B.n11 B.n8 585
R404 B.n769 B.n768 585
R405 B.n768 B.n767 585
R406 B.n10 B.n9 585
R407 B.n766 B.n10 585
R408 B.n764 B.n763 585
R409 B.n765 B.n764 585
R410 B.n762 B.n15 585
R411 B.n18 B.n15 585
R412 B.n761 B.n760 585
R413 B.n760 B.n759 585
R414 B.n17 B.n16 585
R415 B.n758 B.n17 585
R416 B.n756 B.n755 585
R417 B.n757 B.n756 585
R418 B.n754 B.n23 585
R419 B.n23 B.n22 585
R420 B.n753 B.n752 585
R421 B.n752 B.n751 585
R422 B.n25 B.n24 585
R423 B.n750 B.n25 585
R424 B.n748 B.n747 585
R425 B.n749 B.n748 585
R426 B.n746 B.n30 585
R427 B.n30 B.n29 585
R428 B.n745 B.n744 585
R429 B.n744 B.n743 585
R430 B.n777 B.n776 585
R431 B.n776 B.n775 585
R432 B.n670 B.n362 511.721
R433 B.n744 B.n32 511.721
R434 B.n668 B.n364 511.721
R435 B.n740 B.n33 511.721
R436 B.n742 B.n741 256.663
R437 B.n742 B.n92 256.663
R438 B.n742 B.n91 256.663
R439 B.n742 B.n90 256.663
R440 B.n742 B.n89 256.663
R441 B.n742 B.n88 256.663
R442 B.n742 B.n87 256.663
R443 B.n742 B.n86 256.663
R444 B.n742 B.n85 256.663
R445 B.n742 B.n84 256.663
R446 B.n742 B.n83 256.663
R447 B.n742 B.n82 256.663
R448 B.n742 B.n81 256.663
R449 B.n742 B.n80 256.663
R450 B.n742 B.n79 256.663
R451 B.n742 B.n78 256.663
R452 B.n742 B.n77 256.663
R453 B.n742 B.n76 256.663
R454 B.n742 B.n75 256.663
R455 B.n742 B.n74 256.663
R456 B.n742 B.n73 256.663
R457 B.n742 B.n72 256.663
R458 B.n742 B.n71 256.663
R459 B.n742 B.n70 256.663
R460 B.n742 B.n69 256.663
R461 B.n742 B.n68 256.663
R462 B.n742 B.n67 256.663
R463 B.n742 B.n66 256.663
R464 B.n742 B.n65 256.663
R465 B.n742 B.n64 256.663
R466 B.n742 B.n63 256.663
R467 B.n742 B.n62 256.663
R468 B.n742 B.n61 256.663
R469 B.n742 B.n60 256.663
R470 B.n742 B.n59 256.663
R471 B.n742 B.n58 256.663
R472 B.n742 B.n57 256.663
R473 B.n742 B.n56 256.663
R474 B.n742 B.n55 256.663
R475 B.n742 B.n54 256.663
R476 B.n742 B.n53 256.663
R477 B.n742 B.n52 256.663
R478 B.n742 B.n51 256.663
R479 B.n742 B.n50 256.663
R480 B.n742 B.n49 256.663
R481 B.n742 B.n48 256.663
R482 B.n742 B.n47 256.663
R483 B.n742 B.n46 256.663
R484 B.n742 B.n45 256.663
R485 B.n742 B.n44 256.663
R486 B.n742 B.n43 256.663
R487 B.n742 B.n42 256.663
R488 B.n742 B.n41 256.663
R489 B.n742 B.n40 256.663
R490 B.n742 B.n39 256.663
R491 B.n742 B.n38 256.663
R492 B.n742 B.n37 256.663
R493 B.n742 B.n36 256.663
R494 B.n742 B.n35 256.663
R495 B.n742 B.n34 256.663
R496 B.n429 B.n363 256.663
R497 B.n435 B.n363 256.663
R498 B.n437 B.n363 256.663
R499 B.n443 B.n363 256.663
R500 B.n445 B.n363 256.663
R501 B.n451 B.n363 256.663
R502 B.n453 B.n363 256.663
R503 B.n459 B.n363 256.663
R504 B.n461 B.n363 256.663
R505 B.n467 B.n363 256.663
R506 B.n469 B.n363 256.663
R507 B.n475 B.n363 256.663
R508 B.n477 B.n363 256.663
R509 B.n483 B.n363 256.663
R510 B.n485 B.n363 256.663
R511 B.n491 B.n363 256.663
R512 B.n493 B.n363 256.663
R513 B.n499 B.n363 256.663
R514 B.n501 B.n363 256.663
R515 B.n507 B.n363 256.663
R516 B.n509 B.n363 256.663
R517 B.n515 B.n363 256.663
R518 B.n517 B.n363 256.663
R519 B.n523 B.n363 256.663
R520 B.n525 B.n363 256.663
R521 B.n531 B.n363 256.663
R522 B.n533 B.n363 256.663
R523 B.n540 B.n363 256.663
R524 B.n542 B.n363 256.663
R525 B.n548 B.n363 256.663
R526 B.n550 B.n363 256.663
R527 B.n556 B.n363 256.663
R528 B.n558 B.n363 256.663
R529 B.n564 B.n363 256.663
R530 B.n566 B.n363 256.663
R531 B.n572 B.n363 256.663
R532 B.n574 B.n363 256.663
R533 B.n580 B.n363 256.663
R534 B.n582 B.n363 256.663
R535 B.n588 B.n363 256.663
R536 B.n590 B.n363 256.663
R537 B.n596 B.n363 256.663
R538 B.n598 B.n363 256.663
R539 B.n604 B.n363 256.663
R540 B.n606 B.n363 256.663
R541 B.n612 B.n363 256.663
R542 B.n614 B.n363 256.663
R543 B.n620 B.n363 256.663
R544 B.n622 B.n363 256.663
R545 B.n628 B.n363 256.663
R546 B.n630 B.n363 256.663
R547 B.n636 B.n363 256.663
R548 B.n638 B.n363 256.663
R549 B.n644 B.n363 256.663
R550 B.n646 B.n363 256.663
R551 B.n652 B.n363 256.663
R552 B.n654 B.n363 256.663
R553 B.n660 B.n363 256.663
R554 B.n663 B.n363 256.663
R555 B.n670 B.n360 163.367
R556 B.n674 B.n360 163.367
R557 B.n674 B.n354 163.367
R558 B.n682 B.n354 163.367
R559 B.n682 B.n352 163.367
R560 B.n686 B.n352 163.367
R561 B.n686 B.n346 163.367
R562 B.n695 B.n346 163.367
R563 B.n695 B.n344 163.367
R564 B.n699 B.n344 163.367
R565 B.n699 B.n339 163.367
R566 B.n709 B.n339 163.367
R567 B.n709 B.n337 163.367
R568 B.n713 B.n337 163.367
R569 B.n713 B.n2 163.367
R570 B.n776 B.n2 163.367
R571 B.n776 B.n3 163.367
R572 B.n772 B.n3 163.367
R573 B.n772 B.n8 163.367
R574 B.n768 B.n8 163.367
R575 B.n768 B.n10 163.367
R576 B.n764 B.n10 163.367
R577 B.n764 B.n15 163.367
R578 B.n760 B.n15 163.367
R579 B.n760 B.n17 163.367
R580 B.n756 B.n17 163.367
R581 B.n756 B.n23 163.367
R582 B.n752 B.n23 163.367
R583 B.n752 B.n25 163.367
R584 B.n748 B.n25 163.367
R585 B.n748 B.n30 163.367
R586 B.n744 B.n30 163.367
R587 B.n430 B.n428 163.367
R588 B.n434 B.n428 163.367
R589 B.n438 B.n436 163.367
R590 B.n442 B.n426 163.367
R591 B.n446 B.n444 163.367
R592 B.n450 B.n424 163.367
R593 B.n454 B.n452 163.367
R594 B.n458 B.n422 163.367
R595 B.n462 B.n460 163.367
R596 B.n466 B.n420 163.367
R597 B.n470 B.n468 163.367
R598 B.n474 B.n418 163.367
R599 B.n478 B.n476 163.367
R600 B.n482 B.n416 163.367
R601 B.n486 B.n484 163.367
R602 B.n490 B.n414 163.367
R603 B.n494 B.n492 163.367
R604 B.n498 B.n412 163.367
R605 B.n502 B.n500 163.367
R606 B.n506 B.n410 163.367
R607 B.n510 B.n508 163.367
R608 B.n514 B.n408 163.367
R609 B.n518 B.n516 163.367
R610 B.n522 B.n406 163.367
R611 B.n526 B.n524 163.367
R612 B.n530 B.n404 163.367
R613 B.n534 B.n532 163.367
R614 B.n539 B.n400 163.367
R615 B.n543 B.n541 163.367
R616 B.n547 B.n398 163.367
R617 B.n551 B.n549 163.367
R618 B.n555 B.n396 163.367
R619 B.n559 B.n557 163.367
R620 B.n563 B.n391 163.367
R621 B.n567 B.n565 163.367
R622 B.n571 B.n389 163.367
R623 B.n575 B.n573 163.367
R624 B.n579 B.n387 163.367
R625 B.n583 B.n581 163.367
R626 B.n587 B.n385 163.367
R627 B.n591 B.n589 163.367
R628 B.n595 B.n383 163.367
R629 B.n599 B.n597 163.367
R630 B.n603 B.n381 163.367
R631 B.n607 B.n605 163.367
R632 B.n611 B.n379 163.367
R633 B.n615 B.n613 163.367
R634 B.n619 B.n377 163.367
R635 B.n623 B.n621 163.367
R636 B.n627 B.n375 163.367
R637 B.n631 B.n629 163.367
R638 B.n635 B.n373 163.367
R639 B.n639 B.n637 163.367
R640 B.n643 B.n371 163.367
R641 B.n647 B.n645 163.367
R642 B.n651 B.n369 163.367
R643 B.n655 B.n653 163.367
R644 B.n659 B.n367 163.367
R645 B.n662 B.n661 163.367
R646 B.n664 B.n364 163.367
R647 B.n668 B.n358 163.367
R648 B.n676 B.n358 163.367
R649 B.n676 B.n356 163.367
R650 B.n680 B.n356 163.367
R651 B.n680 B.n350 163.367
R652 B.n688 B.n350 163.367
R653 B.n688 B.n348 163.367
R654 B.n692 B.n348 163.367
R655 B.n692 B.n342 163.367
R656 B.n701 B.n342 163.367
R657 B.n701 B.n340 163.367
R658 B.n706 B.n340 163.367
R659 B.n706 B.n336 163.367
R660 B.n715 B.n336 163.367
R661 B.n716 B.n715 163.367
R662 B.n716 B.n5 163.367
R663 B.n6 B.n5 163.367
R664 B.n7 B.n6 163.367
R665 B.n721 B.n7 163.367
R666 B.n721 B.n12 163.367
R667 B.n13 B.n12 163.367
R668 B.n14 B.n13 163.367
R669 B.n726 B.n14 163.367
R670 B.n726 B.n19 163.367
R671 B.n20 B.n19 163.367
R672 B.n21 B.n20 163.367
R673 B.n731 B.n21 163.367
R674 B.n731 B.n26 163.367
R675 B.n27 B.n26 163.367
R676 B.n28 B.n27 163.367
R677 B.n736 B.n28 163.367
R678 B.n736 B.n33 163.367
R679 B.n100 B.n99 163.367
R680 B.n104 B.n103 163.367
R681 B.n108 B.n107 163.367
R682 B.n112 B.n111 163.367
R683 B.n116 B.n115 163.367
R684 B.n120 B.n119 163.367
R685 B.n124 B.n123 163.367
R686 B.n128 B.n127 163.367
R687 B.n132 B.n131 163.367
R688 B.n136 B.n135 163.367
R689 B.n140 B.n139 163.367
R690 B.n144 B.n143 163.367
R691 B.n148 B.n147 163.367
R692 B.n152 B.n151 163.367
R693 B.n156 B.n155 163.367
R694 B.n160 B.n159 163.367
R695 B.n164 B.n163 163.367
R696 B.n168 B.n167 163.367
R697 B.n172 B.n171 163.367
R698 B.n176 B.n175 163.367
R699 B.n180 B.n179 163.367
R700 B.n184 B.n183 163.367
R701 B.n188 B.n187 163.367
R702 B.n192 B.n191 163.367
R703 B.n196 B.n195 163.367
R704 B.n200 B.n199 163.367
R705 B.n204 B.n203 163.367
R706 B.n209 B.n208 163.367
R707 B.n213 B.n212 163.367
R708 B.n217 B.n216 163.367
R709 B.n221 B.n220 163.367
R710 B.n225 B.n224 163.367
R711 B.n230 B.n229 163.367
R712 B.n234 B.n233 163.367
R713 B.n238 B.n237 163.367
R714 B.n242 B.n241 163.367
R715 B.n246 B.n245 163.367
R716 B.n250 B.n249 163.367
R717 B.n254 B.n253 163.367
R718 B.n258 B.n257 163.367
R719 B.n262 B.n261 163.367
R720 B.n266 B.n265 163.367
R721 B.n270 B.n269 163.367
R722 B.n274 B.n273 163.367
R723 B.n278 B.n277 163.367
R724 B.n282 B.n281 163.367
R725 B.n286 B.n285 163.367
R726 B.n290 B.n289 163.367
R727 B.n294 B.n293 163.367
R728 B.n298 B.n297 163.367
R729 B.n302 B.n301 163.367
R730 B.n306 B.n305 163.367
R731 B.n310 B.n309 163.367
R732 B.n314 B.n313 163.367
R733 B.n318 B.n317 163.367
R734 B.n322 B.n321 163.367
R735 B.n326 B.n325 163.367
R736 B.n330 B.n329 163.367
R737 B.n332 B.n93 163.367
R738 B.n392 B.t16 85.5716
R739 B.n94 B.t8 85.5716
R740 B.n401 B.t13 85.5499
R741 B.n96 B.t18 85.5499
R742 B.n393 B.t15 72.1898
R743 B.n95 B.t9 72.1898
R744 B.n402 B.t12 72.1681
R745 B.n97 B.t19 72.1681
R746 B.n429 B.n362 71.676
R747 B.n435 B.n434 71.676
R748 B.n438 B.n437 71.676
R749 B.n443 B.n442 71.676
R750 B.n446 B.n445 71.676
R751 B.n451 B.n450 71.676
R752 B.n454 B.n453 71.676
R753 B.n459 B.n458 71.676
R754 B.n462 B.n461 71.676
R755 B.n467 B.n466 71.676
R756 B.n470 B.n469 71.676
R757 B.n475 B.n474 71.676
R758 B.n478 B.n477 71.676
R759 B.n483 B.n482 71.676
R760 B.n486 B.n485 71.676
R761 B.n491 B.n490 71.676
R762 B.n494 B.n493 71.676
R763 B.n499 B.n498 71.676
R764 B.n502 B.n501 71.676
R765 B.n507 B.n506 71.676
R766 B.n510 B.n509 71.676
R767 B.n515 B.n514 71.676
R768 B.n518 B.n517 71.676
R769 B.n523 B.n522 71.676
R770 B.n526 B.n525 71.676
R771 B.n531 B.n530 71.676
R772 B.n534 B.n533 71.676
R773 B.n540 B.n539 71.676
R774 B.n543 B.n542 71.676
R775 B.n548 B.n547 71.676
R776 B.n551 B.n550 71.676
R777 B.n556 B.n555 71.676
R778 B.n559 B.n558 71.676
R779 B.n564 B.n563 71.676
R780 B.n567 B.n566 71.676
R781 B.n572 B.n571 71.676
R782 B.n575 B.n574 71.676
R783 B.n580 B.n579 71.676
R784 B.n583 B.n582 71.676
R785 B.n588 B.n587 71.676
R786 B.n591 B.n590 71.676
R787 B.n596 B.n595 71.676
R788 B.n599 B.n598 71.676
R789 B.n604 B.n603 71.676
R790 B.n607 B.n606 71.676
R791 B.n612 B.n611 71.676
R792 B.n615 B.n614 71.676
R793 B.n620 B.n619 71.676
R794 B.n623 B.n622 71.676
R795 B.n628 B.n627 71.676
R796 B.n631 B.n630 71.676
R797 B.n636 B.n635 71.676
R798 B.n639 B.n638 71.676
R799 B.n644 B.n643 71.676
R800 B.n647 B.n646 71.676
R801 B.n652 B.n651 71.676
R802 B.n655 B.n654 71.676
R803 B.n660 B.n659 71.676
R804 B.n663 B.n662 71.676
R805 B.n34 B.n32 71.676
R806 B.n100 B.n35 71.676
R807 B.n104 B.n36 71.676
R808 B.n108 B.n37 71.676
R809 B.n112 B.n38 71.676
R810 B.n116 B.n39 71.676
R811 B.n120 B.n40 71.676
R812 B.n124 B.n41 71.676
R813 B.n128 B.n42 71.676
R814 B.n132 B.n43 71.676
R815 B.n136 B.n44 71.676
R816 B.n140 B.n45 71.676
R817 B.n144 B.n46 71.676
R818 B.n148 B.n47 71.676
R819 B.n152 B.n48 71.676
R820 B.n156 B.n49 71.676
R821 B.n160 B.n50 71.676
R822 B.n164 B.n51 71.676
R823 B.n168 B.n52 71.676
R824 B.n172 B.n53 71.676
R825 B.n176 B.n54 71.676
R826 B.n180 B.n55 71.676
R827 B.n184 B.n56 71.676
R828 B.n188 B.n57 71.676
R829 B.n192 B.n58 71.676
R830 B.n196 B.n59 71.676
R831 B.n200 B.n60 71.676
R832 B.n204 B.n61 71.676
R833 B.n209 B.n62 71.676
R834 B.n213 B.n63 71.676
R835 B.n217 B.n64 71.676
R836 B.n221 B.n65 71.676
R837 B.n225 B.n66 71.676
R838 B.n230 B.n67 71.676
R839 B.n234 B.n68 71.676
R840 B.n238 B.n69 71.676
R841 B.n242 B.n70 71.676
R842 B.n246 B.n71 71.676
R843 B.n250 B.n72 71.676
R844 B.n254 B.n73 71.676
R845 B.n258 B.n74 71.676
R846 B.n262 B.n75 71.676
R847 B.n266 B.n76 71.676
R848 B.n270 B.n77 71.676
R849 B.n274 B.n78 71.676
R850 B.n278 B.n79 71.676
R851 B.n282 B.n80 71.676
R852 B.n286 B.n81 71.676
R853 B.n290 B.n82 71.676
R854 B.n294 B.n83 71.676
R855 B.n298 B.n84 71.676
R856 B.n302 B.n85 71.676
R857 B.n306 B.n86 71.676
R858 B.n310 B.n87 71.676
R859 B.n314 B.n88 71.676
R860 B.n318 B.n89 71.676
R861 B.n322 B.n90 71.676
R862 B.n326 B.n91 71.676
R863 B.n330 B.n92 71.676
R864 B.n741 B.n93 71.676
R865 B.n741 B.n740 71.676
R866 B.n332 B.n92 71.676
R867 B.n329 B.n91 71.676
R868 B.n325 B.n90 71.676
R869 B.n321 B.n89 71.676
R870 B.n317 B.n88 71.676
R871 B.n313 B.n87 71.676
R872 B.n309 B.n86 71.676
R873 B.n305 B.n85 71.676
R874 B.n301 B.n84 71.676
R875 B.n297 B.n83 71.676
R876 B.n293 B.n82 71.676
R877 B.n289 B.n81 71.676
R878 B.n285 B.n80 71.676
R879 B.n281 B.n79 71.676
R880 B.n277 B.n78 71.676
R881 B.n273 B.n77 71.676
R882 B.n269 B.n76 71.676
R883 B.n265 B.n75 71.676
R884 B.n261 B.n74 71.676
R885 B.n257 B.n73 71.676
R886 B.n253 B.n72 71.676
R887 B.n249 B.n71 71.676
R888 B.n245 B.n70 71.676
R889 B.n241 B.n69 71.676
R890 B.n237 B.n68 71.676
R891 B.n233 B.n67 71.676
R892 B.n229 B.n66 71.676
R893 B.n224 B.n65 71.676
R894 B.n220 B.n64 71.676
R895 B.n216 B.n63 71.676
R896 B.n212 B.n62 71.676
R897 B.n208 B.n61 71.676
R898 B.n203 B.n60 71.676
R899 B.n199 B.n59 71.676
R900 B.n195 B.n58 71.676
R901 B.n191 B.n57 71.676
R902 B.n187 B.n56 71.676
R903 B.n183 B.n55 71.676
R904 B.n179 B.n54 71.676
R905 B.n175 B.n53 71.676
R906 B.n171 B.n52 71.676
R907 B.n167 B.n51 71.676
R908 B.n163 B.n50 71.676
R909 B.n159 B.n49 71.676
R910 B.n155 B.n48 71.676
R911 B.n151 B.n47 71.676
R912 B.n147 B.n46 71.676
R913 B.n143 B.n45 71.676
R914 B.n139 B.n44 71.676
R915 B.n135 B.n43 71.676
R916 B.n131 B.n42 71.676
R917 B.n127 B.n41 71.676
R918 B.n123 B.n40 71.676
R919 B.n119 B.n39 71.676
R920 B.n115 B.n38 71.676
R921 B.n111 B.n37 71.676
R922 B.n107 B.n36 71.676
R923 B.n103 B.n35 71.676
R924 B.n99 B.n34 71.676
R925 B.n430 B.n429 71.676
R926 B.n436 B.n435 71.676
R927 B.n437 B.n426 71.676
R928 B.n444 B.n443 71.676
R929 B.n445 B.n424 71.676
R930 B.n452 B.n451 71.676
R931 B.n453 B.n422 71.676
R932 B.n460 B.n459 71.676
R933 B.n461 B.n420 71.676
R934 B.n468 B.n467 71.676
R935 B.n469 B.n418 71.676
R936 B.n476 B.n475 71.676
R937 B.n477 B.n416 71.676
R938 B.n484 B.n483 71.676
R939 B.n485 B.n414 71.676
R940 B.n492 B.n491 71.676
R941 B.n493 B.n412 71.676
R942 B.n500 B.n499 71.676
R943 B.n501 B.n410 71.676
R944 B.n508 B.n507 71.676
R945 B.n509 B.n408 71.676
R946 B.n516 B.n515 71.676
R947 B.n517 B.n406 71.676
R948 B.n524 B.n523 71.676
R949 B.n525 B.n404 71.676
R950 B.n532 B.n531 71.676
R951 B.n533 B.n400 71.676
R952 B.n541 B.n540 71.676
R953 B.n542 B.n398 71.676
R954 B.n549 B.n548 71.676
R955 B.n550 B.n396 71.676
R956 B.n557 B.n556 71.676
R957 B.n558 B.n391 71.676
R958 B.n565 B.n564 71.676
R959 B.n566 B.n389 71.676
R960 B.n573 B.n572 71.676
R961 B.n574 B.n387 71.676
R962 B.n581 B.n580 71.676
R963 B.n582 B.n385 71.676
R964 B.n589 B.n588 71.676
R965 B.n590 B.n383 71.676
R966 B.n597 B.n596 71.676
R967 B.n598 B.n381 71.676
R968 B.n605 B.n604 71.676
R969 B.n606 B.n379 71.676
R970 B.n613 B.n612 71.676
R971 B.n614 B.n377 71.676
R972 B.n621 B.n620 71.676
R973 B.n622 B.n375 71.676
R974 B.n629 B.n628 71.676
R975 B.n630 B.n373 71.676
R976 B.n637 B.n636 71.676
R977 B.n638 B.n371 71.676
R978 B.n645 B.n644 71.676
R979 B.n646 B.n369 71.676
R980 B.n653 B.n652 71.676
R981 B.n654 B.n367 71.676
R982 B.n661 B.n660 71.676
R983 B.n664 B.n663 71.676
R984 B.n669 B.n363 69.9936
R985 B.n743 B.n742 69.9936
R986 B.n394 B.n393 59.5399
R987 B.n537 B.n402 59.5399
R988 B.n206 B.n97 59.5399
R989 B.n227 B.n95 59.5399
R990 B.n669 B.n359 34.2417
R991 B.n675 B.n359 34.2417
R992 B.n675 B.n355 34.2417
R993 B.n681 B.n355 34.2417
R994 B.n687 B.n351 34.2417
R995 B.n687 B.n347 34.2417
R996 B.n694 B.n347 34.2417
R997 B.n694 B.n693 34.2417
R998 B.n700 B.n343 34.2417
R999 B.n708 B.n707 34.2417
R1000 B.n714 B.n4 34.2417
R1001 B.n775 B.n4 34.2417
R1002 B.n775 B.n774 34.2417
R1003 B.n774 B.n773 34.2417
R1004 B.n767 B.n11 34.2417
R1005 B.n766 B.n765 34.2417
R1006 B.n759 B.n18 34.2417
R1007 B.n759 B.n758 34.2417
R1008 B.n758 B.n757 34.2417
R1009 B.n757 B.n22 34.2417
R1010 B.n751 B.n750 34.2417
R1011 B.n750 B.n749 34.2417
R1012 B.n749 B.n29 34.2417
R1013 B.n743 B.n29 34.2417
R1014 B.n745 B.n31 33.2493
R1015 B.n739 B.n738 33.2493
R1016 B.n667 B.n666 33.2493
R1017 B.n671 B.n361 33.2493
R1018 B.t11 B.n351 31.2205
R1019 B.t7 B.n22 31.2205
R1020 B.n700 B.t5 23.1637
R1021 B.n765 B.t0 23.1637
R1022 B.n708 B.t1 22.1566
R1023 B.n767 B.t2 22.1566
R1024 B.n714 B.t4 21.1495
R1025 B.n773 B.t3 21.1495
R1026 B B.n777 18.0485
R1027 B.n393 B.n392 13.3823
R1028 B.n402 B.n401 13.3823
R1029 B.n97 B.n96 13.3823
R1030 B.n95 B.n94 13.3823
R1031 B.n707 B.t4 13.0927
R1032 B.n11 B.t3 13.0927
R1033 B.n343 B.t1 12.0856
R1034 B.t2 B.n766 12.0856
R1035 B.n693 B.t5 11.0785
R1036 B.n18 B.t0 11.0785
R1037 B.n98 B.n31 10.6151
R1038 B.n101 B.n98 10.6151
R1039 B.n102 B.n101 10.6151
R1040 B.n105 B.n102 10.6151
R1041 B.n106 B.n105 10.6151
R1042 B.n109 B.n106 10.6151
R1043 B.n110 B.n109 10.6151
R1044 B.n113 B.n110 10.6151
R1045 B.n114 B.n113 10.6151
R1046 B.n117 B.n114 10.6151
R1047 B.n118 B.n117 10.6151
R1048 B.n121 B.n118 10.6151
R1049 B.n122 B.n121 10.6151
R1050 B.n125 B.n122 10.6151
R1051 B.n126 B.n125 10.6151
R1052 B.n129 B.n126 10.6151
R1053 B.n130 B.n129 10.6151
R1054 B.n133 B.n130 10.6151
R1055 B.n134 B.n133 10.6151
R1056 B.n137 B.n134 10.6151
R1057 B.n138 B.n137 10.6151
R1058 B.n141 B.n138 10.6151
R1059 B.n142 B.n141 10.6151
R1060 B.n145 B.n142 10.6151
R1061 B.n146 B.n145 10.6151
R1062 B.n149 B.n146 10.6151
R1063 B.n150 B.n149 10.6151
R1064 B.n153 B.n150 10.6151
R1065 B.n154 B.n153 10.6151
R1066 B.n157 B.n154 10.6151
R1067 B.n158 B.n157 10.6151
R1068 B.n161 B.n158 10.6151
R1069 B.n162 B.n161 10.6151
R1070 B.n165 B.n162 10.6151
R1071 B.n166 B.n165 10.6151
R1072 B.n169 B.n166 10.6151
R1073 B.n170 B.n169 10.6151
R1074 B.n173 B.n170 10.6151
R1075 B.n174 B.n173 10.6151
R1076 B.n177 B.n174 10.6151
R1077 B.n178 B.n177 10.6151
R1078 B.n181 B.n178 10.6151
R1079 B.n182 B.n181 10.6151
R1080 B.n185 B.n182 10.6151
R1081 B.n186 B.n185 10.6151
R1082 B.n189 B.n186 10.6151
R1083 B.n190 B.n189 10.6151
R1084 B.n193 B.n190 10.6151
R1085 B.n194 B.n193 10.6151
R1086 B.n197 B.n194 10.6151
R1087 B.n198 B.n197 10.6151
R1088 B.n201 B.n198 10.6151
R1089 B.n202 B.n201 10.6151
R1090 B.n205 B.n202 10.6151
R1091 B.n210 B.n207 10.6151
R1092 B.n211 B.n210 10.6151
R1093 B.n214 B.n211 10.6151
R1094 B.n215 B.n214 10.6151
R1095 B.n218 B.n215 10.6151
R1096 B.n219 B.n218 10.6151
R1097 B.n222 B.n219 10.6151
R1098 B.n223 B.n222 10.6151
R1099 B.n226 B.n223 10.6151
R1100 B.n231 B.n228 10.6151
R1101 B.n232 B.n231 10.6151
R1102 B.n235 B.n232 10.6151
R1103 B.n236 B.n235 10.6151
R1104 B.n239 B.n236 10.6151
R1105 B.n240 B.n239 10.6151
R1106 B.n243 B.n240 10.6151
R1107 B.n244 B.n243 10.6151
R1108 B.n247 B.n244 10.6151
R1109 B.n248 B.n247 10.6151
R1110 B.n251 B.n248 10.6151
R1111 B.n252 B.n251 10.6151
R1112 B.n255 B.n252 10.6151
R1113 B.n256 B.n255 10.6151
R1114 B.n259 B.n256 10.6151
R1115 B.n260 B.n259 10.6151
R1116 B.n263 B.n260 10.6151
R1117 B.n264 B.n263 10.6151
R1118 B.n267 B.n264 10.6151
R1119 B.n268 B.n267 10.6151
R1120 B.n271 B.n268 10.6151
R1121 B.n272 B.n271 10.6151
R1122 B.n275 B.n272 10.6151
R1123 B.n276 B.n275 10.6151
R1124 B.n279 B.n276 10.6151
R1125 B.n280 B.n279 10.6151
R1126 B.n283 B.n280 10.6151
R1127 B.n284 B.n283 10.6151
R1128 B.n287 B.n284 10.6151
R1129 B.n288 B.n287 10.6151
R1130 B.n291 B.n288 10.6151
R1131 B.n292 B.n291 10.6151
R1132 B.n295 B.n292 10.6151
R1133 B.n296 B.n295 10.6151
R1134 B.n299 B.n296 10.6151
R1135 B.n300 B.n299 10.6151
R1136 B.n303 B.n300 10.6151
R1137 B.n304 B.n303 10.6151
R1138 B.n307 B.n304 10.6151
R1139 B.n308 B.n307 10.6151
R1140 B.n311 B.n308 10.6151
R1141 B.n312 B.n311 10.6151
R1142 B.n315 B.n312 10.6151
R1143 B.n316 B.n315 10.6151
R1144 B.n319 B.n316 10.6151
R1145 B.n320 B.n319 10.6151
R1146 B.n323 B.n320 10.6151
R1147 B.n324 B.n323 10.6151
R1148 B.n327 B.n324 10.6151
R1149 B.n328 B.n327 10.6151
R1150 B.n331 B.n328 10.6151
R1151 B.n333 B.n331 10.6151
R1152 B.n334 B.n333 10.6151
R1153 B.n739 B.n334 10.6151
R1154 B.n667 B.n357 10.6151
R1155 B.n677 B.n357 10.6151
R1156 B.n678 B.n677 10.6151
R1157 B.n679 B.n678 10.6151
R1158 B.n679 B.n349 10.6151
R1159 B.n689 B.n349 10.6151
R1160 B.n690 B.n689 10.6151
R1161 B.n691 B.n690 10.6151
R1162 B.n691 B.n341 10.6151
R1163 B.n702 B.n341 10.6151
R1164 B.n703 B.n702 10.6151
R1165 B.n705 B.n703 10.6151
R1166 B.n705 B.n704 10.6151
R1167 B.n704 B.n335 10.6151
R1168 B.n717 B.n335 10.6151
R1169 B.n718 B.n717 10.6151
R1170 B.n719 B.n718 10.6151
R1171 B.n720 B.n719 10.6151
R1172 B.n722 B.n720 10.6151
R1173 B.n723 B.n722 10.6151
R1174 B.n724 B.n723 10.6151
R1175 B.n725 B.n724 10.6151
R1176 B.n727 B.n725 10.6151
R1177 B.n728 B.n727 10.6151
R1178 B.n729 B.n728 10.6151
R1179 B.n730 B.n729 10.6151
R1180 B.n732 B.n730 10.6151
R1181 B.n733 B.n732 10.6151
R1182 B.n734 B.n733 10.6151
R1183 B.n735 B.n734 10.6151
R1184 B.n737 B.n735 10.6151
R1185 B.n738 B.n737 10.6151
R1186 B.n431 B.n361 10.6151
R1187 B.n432 B.n431 10.6151
R1188 B.n433 B.n432 10.6151
R1189 B.n433 B.n427 10.6151
R1190 B.n439 B.n427 10.6151
R1191 B.n440 B.n439 10.6151
R1192 B.n441 B.n440 10.6151
R1193 B.n441 B.n425 10.6151
R1194 B.n447 B.n425 10.6151
R1195 B.n448 B.n447 10.6151
R1196 B.n449 B.n448 10.6151
R1197 B.n449 B.n423 10.6151
R1198 B.n455 B.n423 10.6151
R1199 B.n456 B.n455 10.6151
R1200 B.n457 B.n456 10.6151
R1201 B.n457 B.n421 10.6151
R1202 B.n463 B.n421 10.6151
R1203 B.n464 B.n463 10.6151
R1204 B.n465 B.n464 10.6151
R1205 B.n465 B.n419 10.6151
R1206 B.n471 B.n419 10.6151
R1207 B.n472 B.n471 10.6151
R1208 B.n473 B.n472 10.6151
R1209 B.n473 B.n417 10.6151
R1210 B.n479 B.n417 10.6151
R1211 B.n480 B.n479 10.6151
R1212 B.n481 B.n480 10.6151
R1213 B.n481 B.n415 10.6151
R1214 B.n487 B.n415 10.6151
R1215 B.n488 B.n487 10.6151
R1216 B.n489 B.n488 10.6151
R1217 B.n489 B.n413 10.6151
R1218 B.n495 B.n413 10.6151
R1219 B.n496 B.n495 10.6151
R1220 B.n497 B.n496 10.6151
R1221 B.n497 B.n411 10.6151
R1222 B.n503 B.n411 10.6151
R1223 B.n504 B.n503 10.6151
R1224 B.n505 B.n504 10.6151
R1225 B.n505 B.n409 10.6151
R1226 B.n511 B.n409 10.6151
R1227 B.n512 B.n511 10.6151
R1228 B.n513 B.n512 10.6151
R1229 B.n513 B.n407 10.6151
R1230 B.n519 B.n407 10.6151
R1231 B.n520 B.n519 10.6151
R1232 B.n521 B.n520 10.6151
R1233 B.n521 B.n405 10.6151
R1234 B.n527 B.n405 10.6151
R1235 B.n528 B.n527 10.6151
R1236 B.n529 B.n528 10.6151
R1237 B.n529 B.n403 10.6151
R1238 B.n535 B.n403 10.6151
R1239 B.n536 B.n535 10.6151
R1240 B.n538 B.n399 10.6151
R1241 B.n544 B.n399 10.6151
R1242 B.n545 B.n544 10.6151
R1243 B.n546 B.n545 10.6151
R1244 B.n546 B.n397 10.6151
R1245 B.n552 B.n397 10.6151
R1246 B.n553 B.n552 10.6151
R1247 B.n554 B.n553 10.6151
R1248 B.n554 B.n395 10.6151
R1249 B.n561 B.n560 10.6151
R1250 B.n562 B.n561 10.6151
R1251 B.n562 B.n390 10.6151
R1252 B.n568 B.n390 10.6151
R1253 B.n569 B.n568 10.6151
R1254 B.n570 B.n569 10.6151
R1255 B.n570 B.n388 10.6151
R1256 B.n576 B.n388 10.6151
R1257 B.n577 B.n576 10.6151
R1258 B.n578 B.n577 10.6151
R1259 B.n578 B.n386 10.6151
R1260 B.n584 B.n386 10.6151
R1261 B.n585 B.n584 10.6151
R1262 B.n586 B.n585 10.6151
R1263 B.n586 B.n384 10.6151
R1264 B.n592 B.n384 10.6151
R1265 B.n593 B.n592 10.6151
R1266 B.n594 B.n593 10.6151
R1267 B.n594 B.n382 10.6151
R1268 B.n600 B.n382 10.6151
R1269 B.n601 B.n600 10.6151
R1270 B.n602 B.n601 10.6151
R1271 B.n602 B.n380 10.6151
R1272 B.n608 B.n380 10.6151
R1273 B.n609 B.n608 10.6151
R1274 B.n610 B.n609 10.6151
R1275 B.n610 B.n378 10.6151
R1276 B.n616 B.n378 10.6151
R1277 B.n617 B.n616 10.6151
R1278 B.n618 B.n617 10.6151
R1279 B.n618 B.n376 10.6151
R1280 B.n624 B.n376 10.6151
R1281 B.n625 B.n624 10.6151
R1282 B.n626 B.n625 10.6151
R1283 B.n626 B.n374 10.6151
R1284 B.n632 B.n374 10.6151
R1285 B.n633 B.n632 10.6151
R1286 B.n634 B.n633 10.6151
R1287 B.n634 B.n372 10.6151
R1288 B.n640 B.n372 10.6151
R1289 B.n641 B.n640 10.6151
R1290 B.n642 B.n641 10.6151
R1291 B.n642 B.n370 10.6151
R1292 B.n648 B.n370 10.6151
R1293 B.n649 B.n648 10.6151
R1294 B.n650 B.n649 10.6151
R1295 B.n650 B.n368 10.6151
R1296 B.n656 B.n368 10.6151
R1297 B.n657 B.n656 10.6151
R1298 B.n658 B.n657 10.6151
R1299 B.n658 B.n366 10.6151
R1300 B.n366 B.n365 10.6151
R1301 B.n665 B.n365 10.6151
R1302 B.n666 B.n665 10.6151
R1303 B.n672 B.n671 10.6151
R1304 B.n673 B.n672 10.6151
R1305 B.n673 B.n353 10.6151
R1306 B.n683 B.n353 10.6151
R1307 B.n684 B.n683 10.6151
R1308 B.n685 B.n684 10.6151
R1309 B.n685 B.n345 10.6151
R1310 B.n696 B.n345 10.6151
R1311 B.n697 B.n696 10.6151
R1312 B.n698 B.n697 10.6151
R1313 B.n698 B.n338 10.6151
R1314 B.n710 B.n338 10.6151
R1315 B.n711 B.n710 10.6151
R1316 B.n712 B.n711 10.6151
R1317 B.n712 B.n0 10.6151
R1318 B.n771 B.n1 10.6151
R1319 B.n771 B.n770 10.6151
R1320 B.n770 B.n769 10.6151
R1321 B.n769 B.n9 10.6151
R1322 B.n763 B.n9 10.6151
R1323 B.n763 B.n762 10.6151
R1324 B.n762 B.n761 10.6151
R1325 B.n761 B.n16 10.6151
R1326 B.n755 B.n16 10.6151
R1327 B.n755 B.n754 10.6151
R1328 B.n754 B.n753 10.6151
R1329 B.n753 B.n24 10.6151
R1330 B.n747 B.n24 10.6151
R1331 B.n747 B.n746 10.6151
R1332 B.n746 B.n745 10.6151
R1333 B.n206 B.n205 9.36635
R1334 B.n228 B.n227 9.36635
R1335 B.n537 B.n536 9.36635
R1336 B.n560 B.n394 9.36635
R1337 B.n681 B.t11 3.02179
R1338 B.n751 B.t7 3.02179
R1339 B.n777 B.n0 2.81026
R1340 B.n777 B.n1 2.81026
R1341 B.n207 B.n206 1.24928
R1342 B.n227 B.n226 1.24928
R1343 B.n538 B.n537 1.24928
R1344 B.n395 B.n394 1.24928
R1345 VN.n0 VN.t2 1240.95
R1346 VN.n4 VN.t3 1240.95
R1347 VN.n2 VN.t4 1220.52
R1348 VN.n6 VN.t1 1220.52
R1349 VN.n1 VN.t0 1219.06
R1350 VN.n5 VN.t5 1219.06
R1351 VN.n3 VN.n2 161.3
R1352 VN.n7 VN.n6 161.3
R1353 VN.n7 VN.n4 70.6808
R1354 VN.n3 VN.n0 70.6808
R1355 VN.n2 VN.n1 46.7399
R1356 VN.n6 VN.n5 46.7399
R1357 VN VN.n7 43.7486
R1358 VN.n5 VN.n4 20.4028
R1359 VN.n1 VN.n0 20.4028
R1360 VN VN.n3 0.0516364
R1361 VDD2.n1 VDD2.t3 64.8563
R1362 VDD2.n2 VDD2.t4 64.4658
R1363 VDD2.n1 VDD2.n0 63.364
R1364 VDD2 VDD2.n3 63.3612
R1365 VDD2.n2 VDD2.n1 39.933
R1366 VDD2.n3 VDD2.t0 1.19543
R1367 VDD2.n3 VDD2.t2 1.19543
R1368 VDD2.n0 VDD2.t5 1.19543
R1369 VDD2.n0 VDD2.t1 1.19543
R1370 VDD2 VDD2.n2 0.50481
C0 VDD2 VP 0.269819f
C1 VP VN 5.59803f
C2 VP VDD1 4.16132f
C3 VDD2 VN 4.04606f
C4 VP VTAIL 3.43245f
C5 VDD2 VDD1 0.59273f
C6 VDD1 VN 0.147704f
C7 VDD2 VTAIL 17.2808f
C8 VTAIL VN 3.41748f
C9 VDD1 VTAIL 17.253698f
C10 VDD2 B 5.061409f
C11 VDD1 B 5.272329f
C12 VTAIL B 7.668437f
C13 VN B 7.57942f
C14 VP B 5.047208f
C15 VDD2.t3 B 4.06514f
C16 VDD2.t5 B 0.349838f
C17 VDD2.t1 B 0.349838f
C18 VDD2.n0 B 3.17959f
C19 VDD2.n1 B 2.36408f
C20 VDD2.t4 B 4.06313f
C21 VDD2.n2 B 2.71099f
C22 VDD2.t0 B 0.349838f
C23 VDD2.t2 B 0.349838f
C24 VDD2.n3 B 3.17956f
C25 VN.t2 B 0.943084f
C26 VN.n0 B 0.357927f
C27 VN.t0 B 0.936679f
C28 VN.n1 B 0.374171f
C29 VN.t4 B 0.937099f
C30 VN.n2 B 0.363519f
C31 VN.n3 B 0.161299f
C32 VN.t3 B 0.943084f
C33 VN.n4 B 0.357927f
C34 VN.t1 B 0.937099f
C35 VN.t5 B 0.936679f
C36 VN.n5 B 0.374171f
C37 VN.n6 B 0.363519f
C38 VN.n7 B 2.56196f
C39 VDD1.t3 B 4.08504f
C40 VDD1.t0 B 4.08439f
C41 VDD1.t1 B 0.351494f
C42 VDD1.t4 B 0.351494f
C43 VDD1.n0 B 3.19465f
C44 VDD1.n1 B 2.45056f
C45 VDD1.t2 B 0.351494f
C46 VDD1.t5 B 0.351494f
C47 VDD1.n2 B 3.1942f
C48 VDD1.n3 B 2.69289f
C49 VTAIL.t3 B 0.354546f
C50 VTAIL.t2 B 0.354546f
C51 VTAIL.n0 B 3.14485f
C52 VTAIL.n1 B 0.345793f
C53 VTAIL.t6 B 4.01784f
C54 VTAIL.n2 B 0.473591f
C55 VTAIL.t10 B 0.354546f
C56 VTAIL.t11 B 0.354546f
C57 VTAIL.n3 B 3.14485f
C58 VTAIL.n4 B 2.03058f
C59 VTAIL.t5 B 0.354546f
C60 VTAIL.t1 B 0.354546f
C61 VTAIL.n5 B 3.14485f
C62 VTAIL.n6 B 2.03058f
C63 VTAIL.t4 B 4.01784f
C64 VTAIL.n7 B 0.473587f
C65 VTAIL.t8 B 0.354546f
C66 VTAIL.t9 B 0.354546f
C67 VTAIL.n8 B 3.14485f
C68 VTAIL.n9 B 0.379634f
C69 VTAIL.t7 B 4.01784f
C70 VTAIL.n10 B 2.07264f
C71 VTAIL.t0 B 4.01784f
C72 VTAIL.n11 B 2.05458f
C73 VP.n0 B 0.056507f
C74 VP.t5 B 0.957242f
C75 VP.t2 B 0.963355f
C76 VP.n1 B 0.36562f
C77 VP.t3 B 0.956812f
C78 VP.n2 B 0.382214f
C79 VP.t0 B 0.957242f
C80 VP.n3 B 0.371332f
C81 VP.n4 B 2.58f
C82 VP.n5 B 2.50587f
C83 VP.n6 B 0.371332f
C84 VP.t4 B 0.956812f
C85 VP.n7 B 0.382214f
C86 VP.t1 B 0.957242f
C87 VP.n8 B 0.371332f
C88 VP.n9 B 0.043791f
.ends

