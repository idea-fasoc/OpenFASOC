* NGSPICE file created from diff_pair_sample_1432.ext - technology: sky130A

.subckt diff_pair_sample_1432 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=0 ps=0 w=19.85 l=2.15
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=7.7415 ps=40.48 w=19.85 l=2.15
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=7.7415 ps=40.48 w=19.85 l=2.15
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=7.7415 ps=40.48 w=19.85 l=2.15
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=0 ps=0 w=19.85 l=2.15
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=0 ps=0 w=19.85 l=2.15
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=7.7415 ps=40.48 w=19.85 l=2.15
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.7415 pd=40.48 as=0 ps=0 w=19.85 l=2.15
R0 B.n611 B.n119 585
R1 B.n119 B.n44 585
R2 B.n613 B.n612 585
R3 B.n615 B.n118 585
R4 B.n618 B.n617 585
R5 B.n619 B.n117 585
R6 B.n621 B.n620 585
R7 B.n623 B.n116 585
R8 B.n626 B.n625 585
R9 B.n627 B.n115 585
R10 B.n629 B.n628 585
R11 B.n631 B.n114 585
R12 B.n634 B.n633 585
R13 B.n635 B.n113 585
R14 B.n637 B.n636 585
R15 B.n639 B.n112 585
R16 B.n642 B.n641 585
R17 B.n643 B.n111 585
R18 B.n645 B.n644 585
R19 B.n647 B.n110 585
R20 B.n650 B.n649 585
R21 B.n651 B.n109 585
R22 B.n653 B.n652 585
R23 B.n655 B.n108 585
R24 B.n658 B.n657 585
R25 B.n659 B.n107 585
R26 B.n661 B.n660 585
R27 B.n663 B.n106 585
R28 B.n666 B.n665 585
R29 B.n667 B.n105 585
R30 B.n669 B.n668 585
R31 B.n671 B.n104 585
R32 B.n674 B.n673 585
R33 B.n675 B.n103 585
R34 B.n677 B.n676 585
R35 B.n679 B.n102 585
R36 B.n682 B.n681 585
R37 B.n683 B.n101 585
R38 B.n685 B.n684 585
R39 B.n687 B.n100 585
R40 B.n690 B.n689 585
R41 B.n691 B.n99 585
R42 B.n693 B.n692 585
R43 B.n695 B.n98 585
R44 B.n698 B.n697 585
R45 B.n699 B.n97 585
R46 B.n701 B.n700 585
R47 B.n703 B.n96 585
R48 B.n706 B.n705 585
R49 B.n707 B.n95 585
R50 B.n709 B.n708 585
R51 B.n711 B.n94 585
R52 B.n714 B.n713 585
R53 B.n715 B.n93 585
R54 B.n717 B.n716 585
R55 B.n719 B.n92 585
R56 B.n722 B.n721 585
R57 B.n723 B.n91 585
R58 B.n725 B.n724 585
R59 B.n727 B.n90 585
R60 B.n730 B.n729 585
R61 B.n731 B.n89 585
R62 B.n733 B.n732 585
R63 B.n735 B.n88 585
R64 B.n737 B.n736 585
R65 B.n739 B.n738 585
R66 B.n742 B.n741 585
R67 B.n743 B.n83 585
R68 B.n745 B.n744 585
R69 B.n747 B.n82 585
R70 B.n750 B.n749 585
R71 B.n751 B.n81 585
R72 B.n753 B.n752 585
R73 B.n755 B.n80 585
R74 B.n758 B.n757 585
R75 B.n760 B.n77 585
R76 B.n762 B.n761 585
R77 B.n764 B.n76 585
R78 B.n767 B.n766 585
R79 B.n768 B.n75 585
R80 B.n770 B.n769 585
R81 B.n772 B.n74 585
R82 B.n775 B.n774 585
R83 B.n776 B.n73 585
R84 B.n778 B.n777 585
R85 B.n780 B.n72 585
R86 B.n783 B.n782 585
R87 B.n784 B.n71 585
R88 B.n786 B.n785 585
R89 B.n788 B.n70 585
R90 B.n791 B.n790 585
R91 B.n792 B.n69 585
R92 B.n794 B.n793 585
R93 B.n796 B.n68 585
R94 B.n799 B.n798 585
R95 B.n800 B.n67 585
R96 B.n802 B.n801 585
R97 B.n804 B.n66 585
R98 B.n807 B.n806 585
R99 B.n808 B.n65 585
R100 B.n810 B.n809 585
R101 B.n812 B.n64 585
R102 B.n815 B.n814 585
R103 B.n816 B.n63 585
R104 B.n818 B.n817 585
R105 B.n820 B.n62 585
R106 B.n823 B.n822 585
R107 B.n824 B.n61 585
R108 B.n826 B.n825 585
R109 B.n828 B.n60 585
R110 B.n831 B.n830 585
R111 B.n832 B.n59 585
R112 B.n834 B.n833 585
R113 B.n836 B.n58 585
R114 B.n839 B.n838 585
R115 B.n840 B.n57 585
R116 B.n842 B.n841 585
R117 B.n844 B.n56 585
R118 B.n847 B.n846 585
R119 B.n848 B.n55 585
R120 B.n850 B.n849 585
R121 B.n852 B.n54 585
R122 B.n855 B.n854 585
R123 B.n856 B.n53 585
R124 B.n858 B.n857 585
R125 B.n860 B.n52 585
R126 B.n863 B.n862 585
R127 B.n864 B.n51 585
R128 B.n866 B.n865 585
R129 B.n868 B.n50 585
R130 B.n871 B.n870 585
R131 B.n872 B.n49 585
R132 B.n874 B.n873 585
R133 B.n876 B.n48 585
R134 B.n879 B.n878 585
R135 B.n880 B.n47 585
R136 B.n882 B.n881 585
R137 B.n884 B.n46 585
R138 B.n887 B.n886 585
R139 B.n888 B.n45 585
R140 B.n610 B.n43 585
R141 B.n891 B.n43 585
R142 B.n609 B.n42 585
R143 B.n892 B.n42 585
R144 B.n608 B.n41 585
R145 B.n893 B.n41 585
R146 B.n607 B.n606 585
R147 B.n606 B.n37 585
R148 B.n605 B.n36 585
R149 B.n899 B.n36 585
R150 B.n604 B.n35 585
R151 B.n900 B.n35 585
R152 B.n603 B.n34 585
R153 B.n901 B.n34 585
R154 B.n602 B.n601 585
R155 B.n601 B.n30 585
R156 B.n600 B.n29 585
R157 B.n907 B.n29 585
R158 B.n599 B.n28 585
R159 B.n908 B.n28 585
R160 B.n598 B.n27 585
R161 B.n909 B.n27 585
R162 B.n597 B.n596 585
R163 B.n596 B.n23 585
R164 B.n595 B.n22 585
R165 B.n915 B.n22 585
R166 B.n594 B.n21 585
R167 B.n916 B.n21 585
R168 B.n593 B.n20 585
R169 B.n917 B.n20 585
R170 B.n592 B.n591 585
R171 B.n591 B.n16 585
R172 B.n590 B.n15 585
R173 B.n923 B.n15 585
R174 B.n589 B.n14 585
R175 B.n924 B.n14 585
R176 B.n588 B.n13 585
R177 B.n925 B.n13 585
R178 B.n587 B.n586 585
R179 B.n586 B.n12 585
R180 B.n585 B.n584 585
R181 B.n585 B.n8 585
R182 B.n583 B.n7 585
R183 B.n932 B.n7 585
R184 B.n582 B.n6 585
R185 B.n933 B.n6 585
R186 B.n581 B.n5 585
R187 B.n934 B.n5 585
R188 B.n580 B.n579 585
R189 B.n579 B.n4 585
R190 B.n578 B.n120 585
R191 B.n578 B.n577 585
R192 B.n568 B.n121 585
R193 B.n122 B.n121 585
R194 B.n570 B.n569 585
R195 B.n571 B.n570 585
R196 B.n567 B.n126 585
R197 B.n130 B.n126 585
R198 B.n566 B.n565 585
R199 B.n565 B.n564 585
R200 B.n128 B.n127 585
R201 B.n129 B.n128 585
R202 B.n557 B.n556 585
R203 B.n558 B.n557 585
R204 B.n555 B.n135 585
R205 B.n135 B.n134 585
R206 B.n554 B.n553 585
R207 B.n553 B.n552 585
R208 B.n137 B.n136 585
R209 B.n138 B.n137 585
R210 B.n545 B.n544 585
R211 B.n546 B.n545 585
R212 B.n543 B.n143 585
R213 B.n143 B.n142 585
R214 B.n542 B.n541 585
R215 B.n541 B.n540 585
R216 B.n145 B.n144 585
R217 B.n146 B.n145 585
R218 B.n533 B.n532 585
R219 B.n534 B.n533 585
R220 B.n531 B.n151 585
R221 B.n151 B.n150 585
R222 B.n530 B.n529 585
R223 B.n529 B.n528 585
R224 B.n153 B.n152 585
R225 B.n154 B.n153 585
R226 B.n521 B.n520 585
R227 B.n522 B.n521 585
R228 B.n519 B.n159 585
R229 B.n159 B.n158 585
R230 B.n518 B.n517 585
R231 B.n517 B.n516 585
R232 B.n513 B.n163 585
R233 B.n512 B.n511 585
R234 B.n509 B.n164 585
R235 B.n509 B.n162 585
R236 B.n508 B.n507 585
R237 B.n506 B.n505 585
R238 B.n504 B.n166 585
R239 B.n502 B.n501 585
R240 B.n500 B.n167 585
R241 B.n499 B.n498 585
R242 B.n496 B.n168 585
R243 B.n494 B.n493 585
R244 B.n492 B.n169 585
R245 B.n491 B.n490 585
R246 B.n488 B.n170 585
R247 B.n486 B.n485 585
R248 B.n484 B.n171 585
R249 B.n483 B.n482 585
R250 B.n480 B.n172 585
R251 B.n478 B.n477 585
R252 B.n476 B.n173 585
R253 B.n475 B.n474 585
R254 B.n472 B.n174 585
R255 B.n470 B.n469 585
R256 B.n468 B.n175 585
R257 B.n467 B.n466 585
R258 B.n464 B.n176 585
R259 B.n462 B.n461 585
R260 B.n460 B.n177 585
R261 B.n459 B.n458 585
R262 B.n456 B.n178 585
R263 B.n454 B.n453 585
R264 B.n452 B.n179 585
R265 B.n451 B.n450 585
R266 B.n448 B.n180 585
R267 B.n446 B.n445 585
R268 B.n444 B.n181 585
R269 B.n443 B.n442 585
R270 B.n440 B.n182 585
R271 B.n438 B.n437 585
R272 B.n436 B.n183 585
R273 B.n435 B.n434 585
R274 B.n432 B.n184 585
R275 B.n430 B.n429 585
R276 B.n428 B.n185 585
R277 B.n427 B.n426 585
R278 B.n424 B.n186 585
R279 B.n422 B.n421 585
R280 B.n420 B.n187 585
R281 B.n419 B.n418 585
R282 B.n416 B.n188 585
R283 B.n414 B.n413 585
R284 B.n412 B.n189 585
R285 B.n411 B.n410 585
R286 B.n408 B.n190 585
R287 B.n406 B.n405 585
R288 B.n404 B.n191 585
R289 B.n403 B.n402 585
R290 B.n400 B.n192 585
R291 B.n398 B.n397 585
R292 B.n396 B.n193 585
R293 B.n395 B.n394 585
R294 B.n392 B.n194 585
R295 B.n390 B.n389 585
R296 B.n388 B.n195 585
R297 B.n387 B.n386 585
R298 B.n384 B.n383 585
R299 B.n382 B.n381 585
R300 B.n380 B.n200 585
R301 B.n378 B.n377 585
R302 B.n376 B.n201 585
R303 B.n375 B.n374 585
R304 B.n372 B.n202 585
R305 B.n370 B.n369 585
R306 B.n368 B.n203 585
R307 B.n366 B.n365 585
R308 B.n363 B.n206 585
R309 B.n361 B.n360 585
R310 B.n359 B.n207 585
R311 B.n358 B.n357 585
R312 B.n355 B.n208 585
R313 B.n353 B.n352 585
R314 B.n351 B.n209 585
R315 B.n350 B.n349 585
R316 B.n347 B.n210 585
R317 B.n345 B.n344 585
R318 B.n343 B.n211 585
R319 B.n342 B.n341 585
R320 B.n339 B.n212 585
R321 B.n337 B.n336 585
R322 B.n335 B.n213 585
R323 B.n334 B.n333 585
R324 B.n331 B.n214 585
R325 B.n329 B.n328 585
R326 B.n327 B.n215 585
R327 B.n326 B.n325 585
R328 B.n323 B.n216 585
R329 B.n321 B.n320 585
R330 B.n319 B.n217 585
R331 B.n318 B.n317 585
R332 B.n315 B.n218 585
R333 B.n313 B.n312 585
R334 B.n311 B.n219 585
R335 B.n310 B.n309 585
R336 B.n307 B.n220 585
R337 B.n305 B.n304 585
R338 B.n303 B.n221 585
R339 B.n302 B.n301 585
R340 B.n299 B.n222 585
R341 B.n297 B.n296 585
R342 B.n295 B.n223 585
R343 B.n294 B.n293 585
R344 B.n291 B.n224 585
R345 B.n289 B.n288 585
R346 B.n287 B.n225 585
R347 B.n286 B.n285 585
R348 B.n283 B.n226 585
R349 B.n281 B.n280 585
R350 B.n279 B.n227 585
R351 B.n278 B.n277 585
R352 B.n275 B.n228 585
R353 B.n273 B.n272 585
R354 B.n271 B.n229 585
R355 B.n270 B.n269 585
R356 B.n267 B.n230 585
R357 B.n265 B.n264 585
R358 B.n263 B.n231 585
R359 B.n262 B.n261 585
R360 B.n259 B.n232 585
R361 B.n257 B.n256 585
R362 B.n255 B.n233 585
R363 B.n254 B.n253 585
R364 B.n251 B.n234 585
R365 B.n249 B.n248 585
R366 B.n247 B.n235 585
R367 B.n246 B.n245 585
R368 B.n243 B.n236 585
R369 B.n241 B.n240 585
R370 B.n239 B.n238 585
R371 B.n161 B.n160 585
R372 B.n515 B.n514 585
R373 B.n516 B.n515 585
R374 B.n157 B.n156 585
R375 B.n158 B.n157 585
R376 B.n524 B.n523 585
R377 B.n523 B.n522 585
R378 B.n525 B.n155 585
R379 B.n155 B.n154 585
R380 B.n527 B.n526 585
R381 B.n528 B.n527 585
R382 B.n149 B.n148 585
R383 B.n150 B.n149 585
R384 B.n536 B.n535 585
R385 B.n535 B.n534 585
R386 B.n537 B.n147 585
R387 B.n147 B.n146 585
R388 B.n539 B.n538 585
R389 B.n540 B.n539 585
R390 B.n141 B.n140 585
R391 B.n142 B.n141 585
R392 B.n548 B.n547 585
R393 B.n547 B.n546 585
R394 B.n549 B.n139 585
R395 B.n139 B.n138 585
R396 B.n551 B.n550 585
R397 B.n552 B.n551 585
R398 B.n133 B.n132 585
R399 B.n134 B.n133 585
R400 B.n560 B.n559 585
R401 B.n559 B.n558 585
R402 B.n561 B.n131 585
R403 B.n131 B.n129 585
R404 B.n563 B.n562 585
R405 B.n564 B.n563 585
R406 B.n125 B.n124 585
R407 B.n130 B.n125 585
R408 B.n573 B.n572 585
R409 B.n572 B.n571 585
R410 B.n574 B.n123 585
R411 B.n123 B.n122 585
R412 B.n576 B.n575 585
R413 B.n577 B.n576 585
R414 B.n3 B.n0 585
R415 B.n4 B.n3 585
R416 B.n931 B.n1 585
R417 B.n932 B.n931 585
R418 B.n930 B.n929 585
R419 B.n930 B.n8 585
R420 B.n928 B.n9 585
R421 B.n12 B.n9 585
R422 B.n927 B.n926 585
R423 B.n926 B.n925 585
R424 B.n11 B.n10 585
R425 B.n924 B.n11 585
R426 B.n922 B.n921 585
R427 B.n923 B.n922 585
R428 B.n920 B.n17 585
R429 B.n17 B.n16 585
R430 B.n919 B.n918 585
R431 B.n918 B.n917 585
R432 B.n19 B.n18 585
R433 B.n916 B.n19 585
R434 B.n914 B.n913 585
R435 B.n915 B.n914 585
R436 B.n912 B.n24 585
R437 B.n24 B.n23 585
R438 B.n911 B.n910 585
R439 B.n910 B.n909 585
R440 B.n26 B.n25 585
R441 B.n908 B.n26 585
R442 B.n906 B.n905 585
R443 B.n907 B.n906 585
R444 B.n904 B.n31 585
R445 B.n31 B.n30 585
R446 B.n903 B.n902 585
R447 B.n902 B.n901 585
R448 B.n33 B.n32 585
R449 B.n900 B.n33 585
R450 B.n898 B.n897 585
R451 B.n899 B.n898 585
R452 B.n896 B.n38 585
R453 B.n38 B.n37 585
R454 B.n895 B.n894 585
R455 B.n894 B.n893 585
R456 B.n40 B.n39 585
R457 B.n892 B.n40 585
R458 B.n890 B.n889 585
R459 B.n891 B.n890 585
R460 B.n935 B.n934 585
R461 B.n933 B.n2 585
R462 B.n890 B.n45 530.939
R463 B.n119 B.n43 530.939
R464 B.n517 B.n161 530.939
R465 B.n515 B.n163 530.939
R466 B.n78 B.t9 429.755
R467 B.n84 B.t13 429.755
R468 B.n204 B.t6 429.755
R469 B.n196 B.t2 429.755
R470 B.n614 B.n44 256.663
R471 B.n616 B.n44 256.663
R472 B.n622 B.n44 256.663
R473 B.n624 B.n44 256.663
R474 B.n630 B.n44 256.663
R475 B.n632 B.n44 256.663
R476 B.n638 B.n44 256.663
R477 B.n640 B.n44 256.663
R478 B.n646 B.n44 256.663
R479 B.n648 B.n44 256.663
R480 B.n654 B.n44 256.663
R481 B.n656 B.n44 256.663
R482 B.n662 B.n44 256.663
R483 B.n664 B.n44 256.663
R484 B.n670 B.n44 256.663
R485 B.n672 B.n44 256.663
R486 B.n678 B.n44 256.663
R487 B.n680 B.n44 256.663
R488 B.n686 B.n44 256.663
R489 B.n688 B.n44 256.663
R490 B.n694 B.n44 256.663
R491 B.n696 B.n44 256.663
R492 B.n702 B.n44 256.663
R493 B.n704 B.n44 256.663
R494 B.n710 B.n44 256.663
R495 B.n712 B.n44 256.663
R496 B.n718 B.n44 256.663
R497 B.n720 B.n44 256.663
R498 B.n726 B.n44 256.663
R499 B.n728 B.n44 256.663
R500 B.n734 B.n44 256.663
R501 B.n87 B.n44 256.663
R502 B.n740 B.n44 256.663
R503 B.n746 B.n44 256.663
R504 B.n748 B.n44 256.663
R505 B.n754 B.n44 256.663
R506 B.n756 B.n44 256.663
R507 B.n763 B.n44 256.663
R508 B.n765 B.n44 256.663
R509 B.n771 B.n44 256.663
R510 B.n773 B.n44 256.663
R511 B.n779 B.n44 256.663
R512 B.n781 B.n44 256.663
R513 B.n787 B.n44 256.663
R514 B.n789 B.n44 256.663
R515 B.n795 B.n44 256.663
R516 B.n797 B.n44 256.663
R517 B.n803 B.n44 256.663
R518 B.n805 B.n44 256.663
R519 B.n811 B.n44 256.663
R520 B.n813 B.n44 256.663
R521 B.n819 B.n44 256.663
R522 B.n821 B.n44 256.663
R523 B.n827 B.n44 256.663
R524 B.n829 B.n44 256.663
R525 B.n835 B.n44 256.663
R526 B.n837 B.n44 256.663
R527 B.n843 B.n44 256.663
R528 B.n845 B.n44 256.663
R529 B.n851 B.n44 256.663
R530 B.n853 B.n44 256.663
R531 B.n859 B.n44 256.663
R532 B.n861 B.n44 256.663
R533 B.n867 B.n44 256.663
R534 B.n869 B.n44 256.663
R535 B.n875 B.n44 256.663
R536 B.n877 B.n44 256.663
R537 B.n883 B.n44 256.663
R538 B.n885 B.n44 256.663
R539 B.n510 B.n162 256.663
R540 B.n165 B.n162 256.663
R541 B.n503 B.n162 256.663
R542 B.n497 B.n162 256.663
R543 B.n495 B.n162 256.663
R544 B.n489 B.n162 256.663
R545 B.n487 B.n162 256.663
R546 B.n481 B.n162 256.663
R547 B.n479 B.n162 256.663
R548 B.n473 B.n162 256.663
R549 B.n471 B.n162 256.663
R550 B.n465 B.n162 256.663
R551 B.n463 B.n162 256.663
R552 B.n457 B.n162 256.663
R553 B.n455 B.n162 256.663
R554 B.n449 B.n162 256.663
R555 B.n447 B.n162 256.663
R556 B.n441 B.n162 256.663
R557 B.n439 B.n162 256.663
R558 B.n433 B.n162 256.663
R559 B.n431 B.n162 256.663
R560 B.n425 B.n162 256.663
R561 B.n423 B.n162 256.663
R562 B.n417 B.n162 256.663
R563 B.n415 B.n162 256.663
R564 B.n409 B.n162 256.663
R565 B.n407 B.n162 256.663
R566 B.n401 B.n162 256.663
R567 B.n399 B.n162 256.663
R568 B.n393 B.n162 256.663
R569 B.n391 B.n162 256.663
R570 B.n385 B.n162 256.663
R571 B.n199 B.n162 256.663
R572 B.n379 B.n162 256.663
R573 B.n373 B.n162 256.663
R574 B.n371 B.n162 256.663
R575 B.n364 B.n162 256.663
R576 B.n362 B.n162 256.663
R577 B.n356 B.n162 256.663
R578 B.n354 B.n162 256.663
R579 B.n348 B.n162 256.663
R580 B.n346 B.n162 256.663
R581 B.n340 B.n162 256.663
R582 B.n338 B.n162 256.663
R583 B.n332 B.n162 256.663
R584 B.n330 B.n162 256.663
R585 B.n324 B.n162 256.663
R586 B.n322 B.n162 256.663
R587 B.n316 B.n162 256.663
R588 B.n314 B.n162 256.663
R589 B.n308 B.n162 256.663
R590 B.n306 B.n162 256.663
R591 B.n300 B.n162 256.663
R592 B.n298 B.n162 256.663
R593 B.n292 B.n162 256.663
R594 B.n290 B.n162 256.663
R595 B.n284 B.n162 256.663
R596 B.n282 B.n162 256.663
R597 B.n276 B.n162 256.663
R598 B.n274 B.n162 256.663
R599 B.n268 B.n162 256.663
R600 B.n266 B.n162 256.663
R601 B.n260 B.n162 256.663
R602 B.n258 B.n162 256.663
R603 B.n252 B.n162 256.663
R604 B.n250 B.n162 256.663
R605 B.n244 B.n162 256.663
R606 B.n242 B.n162 256.663
R607 B.n237 B.n162 256.663
R608 B.n937 B.n936 256.663
R609 B.n886 B.n884 163.367
R610 B.n882 B.n47 163.367
R611 B.n878 B.n876 163.367
R612 B.n874 B.n49 163.367
R613 B.n870 B.n868 163.367
R614 B.n866 B.n51 163.367
R615 B.n862 B.n860 163.367
R616 B.n858 B.n53 163.367
R617 B.n854 B.n852 163.367
R618 B.n850 B.n55 163.367
R619 B.n846 B.n844 163.367
R620 B.n842 B.n57 163.367
R621 B.n838 B.n836 163.367
R622 B.n834 B.n59 163.367
R623 B.n830 B.n828 163.367
R624 B.n826 B.n61 163.367
R625 B.n822 B.n820 163.367
R626 B.n818 B.n63 163.367
R627 B.n814 B.n812 163.367
R628 B.n810 B.n65 163.367
R629 B.n806 B.n804 163.367
R630 B.n802 B.n67 163.367
R631 B.n798 B.n796 163.367
R632 B.n794 B.n69 163.367
R633 B.n790 B.n788 163.367
R634 B.n786 B.n71 163.367
R635 B.n782 B.n780 163.367
R636 B.n778 B.n73 163.367
R637 B.n774 B.n772 163.367
R638 B.n770 B.n75 163.367
R639 B.n766 B.n764 163.367
R640 B.n762 B.n77 163.367
R641 B.n757 B.n755 163.367
R642 B.n753 B.n81 163.367
R643 B.n749 B.n747 163.367
R644 B.n745 B.n83 163.367
R645 B.n741 B.n739 163.367
R646 B.n736 B.n735 163.367
R647 B.n733 B.n89 163.367
R648 B.n729 B.n727 163.367
R649 B.n725 B.n91 163.367
R650 B.n721 B.n719 163.367
R651 B.n717 B.n93 163.367
R652 B.n713 B.n711 163.367
R653 B.n709 B.n95 163.367
R654 B.n705 B.n703 163.367
R655 B.n701 B.n97 163.367
R656 B.n697 B.n695 163.367
R657 B.n693 B.n99 163.367
R658 B.n689 B.n687 163.367
R659 B.n685 B.n101 163.367
R660 B.n681 B.n679 163.367
R661 B.n677 B.n103 163.367
R662 B.n673 B.n671 163.367
R663 B.n669 B.n105 163.367
R664 B.n665 B.n663 163.367
R665 B.n661 B.n107 163.367
R666 B.n657 B.n655 163.367
R667 B.n653 B.n109 163.367
R668 B.n649 B.n647 163.367
R669 B.n645 B.n111 163.367
R670 B.n641 B.n639 163.367
R671 B.n637 B.n113 163.367
R672 B.n633 B.n631 163.367
R673 B.n629 B.n115 163.367
R674 B.n625 B.n623 163.367
R675 B.n621 B.n117 163.367
R676 B.n617 B.n615 163.367
R677 B.n613 B.n119 163.367
R678 B.n517 B.n159 163.367
R679 B.n521 B.n159 163.367
R680 B.n521 B.n153 163.367
R681 B.n529 B.n153 163.367
R682 B.n529 B.n151 163.367
R683 B.n533 B.n151 163.367
R684 B.n533 B.n145 163.367
R685 B.n541 B.n145 163.367
R686 B.n541 B.n143 163.367
R687 B.n545 B.n143 163.367
R688 B.n545 B.n137 163.367
R689 B.n553 B.n137 163.367
R690 B.n553 B.n135 163.367
R691 B.n557 B.n135 163.367
R692 B.n557 B.n128 163.367
R693 B.n565 B.n128 163.367
R694 B.n565 B.n126 163.367
R695 B.n570 B.n126 163.367
R696 B.n570 B.n121 163.367
R697 B.n578 B.n121 163.367
R698 B.n579 B.n578 163.367
R699 B.n579 B.n5 163.367
R700 B.n6 B.n5 163.367
R701 B.n7 B.n6 163.367
R702 B.n585 B.n7 163.367
R703 B.n586 B.n585 163.367
R704 B.n586 B.n13 163.367
R705 B.n14 B.n13 163.367
R706 B.n15 B.n14 163.367
R707 B.n591 B.n15 163.367
R708 B.n591 B.n20 163.367
R709 B.n21 B.n20 163.367
R710 B.n22 B.n21 163.367
R711 B.n596 B.n22 163.367
R712 B.n596 B.n27 163.367
R713 B.n28 B.n27 163.367
R714 B.n29 B.n28 163.367
R715 B.n601 B.n29 163.367
R716 B.n601 B.n34 163.367
R717 B.n35 B.n34 163.367
R718 B.n36 B.n35 163.367
R719 B.n606 B.n36 163.367
R720 B.n606 B.n41 163.367
R721 B.n42 B.n41 163.367
R722 B.n43 B.n42 163.367
R723 B.n511 B.n509 163.367
R724 B.n509 B.n508 163.367
R725 B.n505 B.n504 163.367
R726 B.n502 B.n167 163.367
R727 B.n498 B.n496 163.367
R728 B.n494 B.n169 163.367
R729 B.n490 B.n488 163.367
R730 B.n486 B.n171 163.367
R731 B.n482 B.n480 163.367
R732 B.n478 B.n173 163.367
R733 B.n474 B.n472 163.367
R734 B.n470 B.n175 163.367
R735 B.n466 B.n464 163.367
R736 B.n462 B.n177 163.367
R737 B.n458 B.n456 163.367
R738 B.n454 B.n179 163.367
R739 B.n450 B.n448 163.367
R740 B.n446 B.n181 163.367
R741 B.n442 B.n440 163.367
R742 B.n438 B.n183 163.367
R743 B.n434 B.n432 163.367
R744 B.n430 B.n185 163.367
R745 B.n426 B.n424 163.367
R746 B.n422 B.n187 163.367
R747 B.n418 B.n416 163.367
R748 B.n414 B.n189 163.367
R749 B.n410 B.n408 163.367
R750 B.n406 B.n191 163.367
R751 B.n402 B.n400 163.367
R752 B.n398 B.n193 163.367
R753 B.n394 B.n392 163.367
R754 B.n390 B.n195 163.367
R755 B.n386 B.n384 163.367
R756 B.n381 B.n380 163.367
R757 B.n378 B.n201 163.367
R758 B.n374 B.n372 163.367
R759 B.n370 B.n203 163.367
R760 B.n365 B.n363 163.367
R761 B.n361 B.n207 163.367
R762 B.n357 B.n355 163.367
R763 B.n353 B.n209 163.367
R764 B.n349 B.n347 163.367
R765 B.n345 B.n211 163.367
R766 B.n341 B.n339 163.367
R767 B.n337 B.n213 163.367
R768 B.n333 B.n331 163.367
R769 B.n329 B.n215 163.367
R770 B.n325 B.n323 163.367
R771 B.n321 B.n217 163.367
R772 B.n317 B.n315 163.367
R773 B.n313 B.n219 163.367
R774 B.n309 B.n307 163.367
R775 B.n305 B.n221 163.367
R776 B.n301 B.n299 163.367
R777 B.n297 B.n223 163.367
R778 B.n293 B.n291 163.367
R779 B.n289 B.n225 163.367
R780 B.n285 B.n283 163.367
R781 B.n281 B.n227 163.367
R782 B.n277 B.n275 163.367
R783 B.n273 B.n229 163.367
R784 B.n269 B.n267 163.367
R785 B.n265 B.n231 163.367
R786 B.n261 B.n259 163.367
R787 B.n257 B.n233 163.367
R788 B.n253 B.n251 163.367
R789 B.n249 B.n235 163.367
R790 B.n245 B.n243 163.367
R791 B.n241 B.n238 163.367
R792 B.n515 B.n157 163.367
R793 B.n523 B.n157 163.367
R794 B.n523 B.n155 163.367
R795 B.n527 B.n155 163.367
R796 B.n527 B.n149 163.367
R797 B.n535 B.n149 163.367
R798 B.n535 B.n147 163.367
R799 B.n539 B.n147 163.367
R800 B.n539 B.n141 163.367
R801 B.n547 B.n141 163.367
R802 B.n547 B.n139 163.367
R803 B.n551 B.n139 163.367
R804 B.n551 B.n133 163.367
R805 B.n559 B.n133 163.367
R806 B.n559 B.n131 163.367
R807 B.n563 B.n131 163.367
R808 B.n563 B.n125 163.367
R809 B.n572 B.n125 163.367
R810 B.n572 B.n123 163.367
R811 B.n576 B.n123 163.367
R812 B.n576 B.n3 163.367
R813 B.n935 B.n3 163.367
R814 B.n931 B.n2 163.367
R815 B.n931 B.n930 163.367
R816 B.n930 B.n9 163.367
R817 B.n926 B.n9 163.367
R818 B.n926 B.n11 163.367
R819 B.n922 B.n11 163.367
R820 B.n922 B.n17 163.367
R821 B.n918 B.n17 163.367
R822 B.n918 B.n19 163.367
R823 B.n914 B.n19 163.367
R824 B.n914 B.n24 163.367
R825 B.n910 B.n24 163.367
R826 B.n910 B.n26 163.367
R827 B.n906 B.n26 163.367
R828 B.n906 B.n31 163.367
R829 B.n902 B.n31 163.367
R830 B.n902 B.n33 163.367
R831 B.n898 B.n33 163.367
R832 B.n898 B.n38 163.367
R833 B.n894 B.n38 163.367
R834 B.n894 B.n40 163.367
R835 B.n890 B.n40 163.367
R836 B.n84 B.t14 117.767
R837 B.n204 B.t8 117.767
R838 B.n78 B.t11 117.74
R839 B.n196 B.t5 117.74
R840 B.n885 B.n45 71.676
R841 B.n884 B.n883 71.676
R842 B.n877 B.n47 71.676
R843 B.n876 B.n875 71.676
R844 B.n869 B.n49 71.676
R845 B.n868 B.n867 71.676
R846 B.n861 B.n51 71.676
R847 B.n860 B.n859 71.676
R848 B.n853 B.n53 71.676
R849 B.n852 B.n851 71.676
R850 B.n845 B.n55 71.676
R851 B.n844 B.n843 71.676
R852 B.n837 B.n57 71.676
R853 B.n836 B.n835 71.676
R854 B.n829 B.n59 71.676
R855 B.n828 B.n827 71.676
R856 B.n821 B.n61 71.676
R857 B.n820 B.n819 71.676
R858 B.n813 B.n63 71.676
R859 B.n812 B.n811 71.676
R860 B.n805 B.n65 71.676
R861 B.n804 B.n803 71.676
R862 B.n797 B.n67 71.676
R863 B.n796 B.n795 71.676
R864 B.n789 B.n69 71.676
R865 B.n788 B.n787 71.676
R866 B.n781 B.n71 71.676
R867 B.n780 B.n779 71.676
R868 B.n773 B.n73 71.676
R869 B.n772 B.n771 71.676
R870 B.n765 B.n75 71.676
R871 B.n764 B.n763 71.676
R872 B.n756 B.n77 71.676
R873 B.n755 B.n754 71.676
R874 B.n748 B.n81 71.676
R875 B.n747 B.n746 71.676
R876 B.n740 B.n83 71.676
R877 B.n739 B.n87 71.676
R878 B.n735 B.n734 71.676
R879 B.n728 B.n89 71.676
R880 B.n727 B.n726 71.676
R881 B.n720 B.n91 71.676
R882 B.n719 B.n718 71.676
R883 B.n712 B.n93 71.676
R884 B.n711 B.n710 71.676
R885 B.n704 B.n95 71.676
R886 B.n703 B.n702 71.676
R887 B.n696 B.n97 71.676
R888 B.n695 B.n694 71.676
R889 B.n688 B.n99 71.676
R890 B.n687 B.n686 71.676
R891 B.n680 B.n101 71.676
R892 B.n679 B.n678 71.676
R893 B.n672 B.n103 71.676
R894 B.n671 B.n670 71.676
R895 B.n664 B.n105 71.676
R896 B.n663 B.n662 71.676
R897 B.n656 B.n107 71.676
R898 B.n655 B.n654 71.676
R899 B.n648 B.n109 71.676
R900 B.n647 B.n646 71.676
R901 B.n640 B.n111 71.676
R902 B.n639 B.n638 71.676
R903 B.n632 B.n113 71.676
R904 B.n631 B.n630 71.676
R905 B.n624 B.n115 71.676
R906 B.n623 B.n622 71.676
R907 B.n616 B.n117 71.676
R908 B.n615 B.n614 71.676
R909 B.n614 B.n613 71.676
R910 B.n617 B.n616 71.676
R911 B.n622 B.n621 71.676
R912 B.n625 B.n624 71.676
R913 B.n630 B.n629 71.676
R914 B.n633 B.n632 71.676
R915 B.n638 B.n637 71.676
R916 B.n641 B.n640 71.676
R917 B.n646 B.n645 71.676
R918 B.n649 B.n648 71.676
R919 B.n654 B.n653 71.676
R920 B.n657 B.n656 71.676
R921 B.n662 B.n661 71.676
R922 B.n665 B.n664 71.676
R923 B.n670 B.n669 71.676
R924 B.n673 B.n672 71.676
R925 B.n678 B.n677 71.676
R926 B.n681 B.n680 71.676
R927 B.n686 B.n685 71.676
R928 B.n689 B.n688 71.676
R929 B.n694 B.n693 71.676
R930 B.n697 B.n696 71.676
R931 B.n702 B.n701 71.676
R932 B.n705 B.n704 71.676
R933 B.n710 B.n709 71.676
R934 B.n713 B.n712 71.676
R935 B.n718 B.n717 71.676
R936 B.n721 B.n720 71.676
R937 B.n726 B.n725 71.676
R938 B.n729 B.n728 71.676
R939 B.n734 B.n733 71.676
R940 B.n736 B.n87 71.676
R941 B.n741 B.n740 71.676
R942 B.n746 B.n745 71.676
R943 B.n749 B.n748 71.676
R944 B.n754 B.n753 71.676
R945 B.n757 B.n756 71.676
R946 B.n763 B.n762 71.676
R947 B.n766 B.n765 71.676
R948 B.n771 B.n770 71.676
R949 B.n774 B.n773 71.676
R950 B.n779 B.n778 71.676
R951 B.n782 B.n781 71.676
R952 B.n787 B.n786 71.676
R953 B.n790 B.n789 71.676
R954 B.n795 B.n794 71.676
R955 B.n798 B.n797 71.676
R956 B.n803 B.n802 71.676
R957 B.n806 B.n805 71.676
R958 B.n811 B.n810 71.676
R959 B.n814 B.n813 71.676
R960 B.n819 B.n818 71.676
R961 B.n822 B.n821 71.676
R962 B.n827 B.n826 71.676
R963 B.n830 B.n829 71.676
R964 B.n835 B.n834 71.676
R965 B.n838 B.n837 71.676
R966 B.n843 B.n842 71.676
R967 B.n846 B.n845 71.676
R968 B.n851 B.n850 71.676
R969 B.n854 B.n853 71.676
R970 B.n859 B.n858 71.676
R971 B.n862 B.n861 71.676
R972 B.n867 B.n866 71.676
R973 B.n870 B.n869 71.676
R974 B.n875 B.n874 71.676
R975 B.n878 B.n877 71.676
R976 B.n883 B.n882 71.676
R977 B.n886 B.n885 71.676
R978 B.n510 B.n163 71.676
R979 B.n508 B.n165 71.676
R980 B.n504 B.n503 71.676
R981 B.n497 B.n167 71.676
R982 B.n496 B.n495 71.676
R983 B.n489 B.n169 71.676
R984 B.n488 B.n487 71.676
R985 B.n481 B.n171 71.676
R986 B.n480 B.n479 71.676
R987 B.n473 B.n173 71.676
R988 B.n472 B.n471 71.676
R989 B.n465 B.n175 71.676
R990 B.n464 B.n463 71.676
R991 B.n457 B.n177 71.676
R992 B.n456 B.n455 71.676
R993 B.n449 B.n179 71.676
R994 B.n448 B.n447 71.676
R995 B.n441 B.n181 71.676
R996 B.n440 B.n439 71.676
R997 B.n433 B.n183 71.676
R998 B.n432 B.n431 71.676
R999 B.n425 B.n185 71.676
R1000 B.n424 B.n423 71.676
R1001 B.n417 B.n187 71.676
R1002 B.n416 B.n415 71.676
R1003 B.n409 B.n189 71.676
R1004 B.n408 B.n407 71.676
R1005 B.n401 B.n191 71.676
R1006 B.n400 B.n399 71.676
R1007 B.n393 B.n193 71.676
R1008 B.n392 B.n391 71.676
R1009 B.n385 B.n195 71.676
R1010 B.n384 B.n199 71.676
R1011 B.n380 B.n379 71.676
R1012 B.n373 B.n201 71.676
R1013 B.n372 B.n371 71.676
R1014 B.n364 B.n203 71.676
R1015 B.n363 B.n362 71.676
R1016 B.n356 B.n207 71.676
R1017 B.n355 B.n354 71.676
R1018 B.n348 B.n209 71.676
R1019 B.n347 B.n346 71.676
R1020 B.n340 B.n211 71.676
R1021 B.n339 B.n338 71.676
R1022 B.n332 B.n213 71.676
R1023 B.n331 B.n330 71.676
R1024 B.n324 B.n215 71.676
R1025 B.n323 B.n322 71.676
R1026 B.n316 B.n217 71.676
R1027 B.n315 B.n314 71.676
R1028 B.n308 B.n219 71.676
R1029 B.n307 B.n306 71.676
R1030 B.n300 B.n221 71.676
R1031 B.n299 B.n298 71.676
R1032 B.n292 B.n223 71.676
R1033 B.n291 B.n290 71.676
R1034 B.n284 B.n225 71.676
R1035 B.n283 B.n282 71.676
R1036 B.n276 B.n227 71.676
R1037 B.n275 B.n274 71.676
R1038 B.n268 B.n229 71.676
R1039 B.n267 B.n266 71.676
R1040 B.n260 B.n231 71.676
R1041 B.n259 B.n258 71.676
R1042 B.n252 B.n233 71.676
R1043 B.n251 B.n250 71.676
R1044 B.n244 B.n235 71.676
R1045 B.n243 B.n242 71.676
R1046 B.n238 B.n237 71.676
R1047 B.n511 B.n510 71.676
R1048 B.n505 B.n165 71.676
R1049 B.n503 B.n502 71.676
R1050 B.n498 B.n497 71.676
R1051 B.n495 B.n494 71.676
R1052 B.n490 B.n489 71.676
R1053 B.n487 B.n486 71.676
R1054 B.n482 B.n481 71.676
R1055 B.n479 B.n478 71.676
R1056 B.n474 B.n473 71.676
R1057 B.n471 B.n470 71.676
R1058 B.n466 B.n465 71.676
R1059 B.n463 B.n462 71.676
R1060 B.n458 B.n457 71.676
R1061 B.n455 B.n454 71.676
R1062 B.n450 B.n449 71.676
R1063 B.n447 B.n446 71.676
R1064 B.n442 B.n441 71.676
R1065 B.n439 B.n438 71.676
R1066 B.n434 B.n433 71.676
R1067 B.n431 B.n430 71.676
R1068 B.n426 B.n425 71.676
R1069 B.n423 B.n422 71.676
R1070 B.n418 B.n417 71.676
R1071 B.n415 B.n414 71.676
R1072 B.n410 B.n409 71.676
R1073 B.n407 B.n406 71.676
R1074 B.n402 B.n401 71.676
R1075 B.n399 B.n398 71.676
R1076 B.n394 B.n393 71.676
R1077 B.n391 B.n390 71.676
R1078 B.n386 B.n385 71.676
R1079 B.n381 B.n199 71.676
R1080 B.n379 B.n378 71.676
R1081 B.n374 B.n373 71.676
R1082 B.n371 B.n370 71.676
R1083 B.n365 B.n364 71.676
R1084 B.n362 B.n361 71.676
R1085 B.n357 B.n356 71.676
R1086 B.n354 B.n353 71.676
R1087 B.n349 B.n348 71.676
R1088 B.n346 B.n345 71.676
R1089 B.n341 B.n340 71.676
R1090 B.n338 B.n337 71.676
R1091 B.n333 B.n332 71.676
R1092 B.n330 B.n329 71.676
R1093 B.n325 B.n324 71.676
R1094 B.n322 B.n321 71.676
R1095 B.n317 B.n316 71.676
R1096 B.n314 B.n313 71.676
R1097 B.n309 B.n308 71.676
R1098 B.n306 B.n305 71.676
R1099 B.n301 B.n300 71.676
R1100 B.n298 B.n297 71.676
R1101 B.n293 B.n292 71.676
R1102 B.n290 B.n289 71.676
R1103 B.n285 B.n284 71.676
R1104 B.n282 B.n281 71.676
R1105 B.n277 B.n276 71.676
R1106 B.n274 B.n273 71.676
R1107 B.n269 B.n268 71.676
R1108 B.n266 B.n265 71.676
R1109 B.n261 B.n260 71.676
R1110 B.n258 B.n257 71.676
R1111 B.n253 B.n252 71.676
R1112 B.n250 B.n249 71.676
R1113 B.n245 B.n244 71.676
R1114 B.n242 B.n241 71.676
R1115 B.n237 B.n161 71.676
R1116 B.n936 B.n935 71.676
R1117 B.n936 B.n2 71.676
R1118 B.n85 B.t15 69.6701
R1119 B.n205 B.t7 69.6701
R1120 B.n79 B.t12 69.6434
R1121 B.n197 B.t4 69.6434
R1122 B.n516 B.n162 59.9806
R1123 B.n891 B.n44 59.9806
R1124 B.n759 B.n79 59.5399
R1125 B.n86 B.n85 59.5399
R1126 B.n367 B.n205 59.5399
R1127 B.n198 B.n197 59.5399
R1128 B.n79 B.n78 48.0975
R1129 B.n85 B.n84 48.0975
R1130 B.n205 B.n204 48.0975
R1131 B.n197 B.n196 48.0975
R1132 B.n514 B.n513 34.4981
R1133 B.n518 B.n160 34.4981
R1134 B.n611 B.n610 34.4981
R1135 B.n889 B.n888 34.4981
R1136 B.n516 B.n158 29.7716
R1137 B.n522 B.n158 29.7716
R1138 B.n522 B.n154 29.7716
R1139 B.n528 B.n154 29.7716
R1140 B.n528 B.n150 29.7716
R1141 B.n534 B.n150 29.7716
R1142 B.n540 B.n146 29.7716
R1143 B.n540 B.n142 29.7716
R1144 B.n546 B.n142 29.7716
R1145 B.n546 B.n138 29.7716
R1146 B.n552 B.n138 29.7716
R1147 B.n552 B.n134 29.7716
R1148 B.n558 B.n134 29.7716
R1149 B.n558 B.n129 29.7716
R1150 B.n564 B.n129 29.7716
R1151 B.n564 B.n130 29.7716
R1152 B.n571 B.n122 29.7716
R1153 B.n577 B.n122 29.7716
R1154 B.n577 B.n4 29.7716
R1155 B.n934 B.n4 29.7716
R1156 B.n934 B.n933 29.7716
R1157 B.n933 B.n932 29.7716
R1158 B.n932 B.n8 29.7716
R1159 B.n12 B.n8 29.7716
R1160 B.n925 B.n12 29.7716
R1161 B.n924 B.n923 29.7716
R1162 B.n923 B.n16 29.7716
R1163 B.n917 B.n16 29.7716
R1164 B.n917 B.n916 29.7716
R1165 B.n916 B.n915 29.7716
R1166 B.n915 B.n23 29.7716
R1167 B.n909 B.n23 29.7716
R1168 B.n909 B.n908 29.7716
R1169 B.n908 B.n907 29.7716
R1170 B.n907 B.n30 29.7716
R1171 B.n901 B.n900 29.7716
R1172 B.n900 B.n899 29.7716
R1173 B.n899 B.n37 29.7716
R1174 B.n893 B.n37 29.7716
R1175 B.n893 B.n892 29.7716
R1176 B.n892 B.n891 29.7716
R1177 B.n534 B.t3 22.3289
R1178 B.n571 B.t0 22.3289
R1179 B.n925 B.t1 22.3289
R1180 B.n901 B.t10 22.3289
R1181 B B.n937 18.0485
R1182 B.n514 B.n156 10.6151
R1183 B.n524 B.n156 10.6151
R1184 B.n525 B.n524 10.6151
R1185 B.n526 B.n525 10.6151
R1186 B.n526 B.n148 10.6151
R1187 B.n536 B.n148 10.6151
R1188 B.n537 B.n536 10.6151
R1189 B.n538 B.n537 10.6151
R1190 B.n538 B.n140 10.6151
R1191 B.n548 B.n140 10.6151
R1192 B.n549 B.n548 10.6151
R1193 B.n550 B.n549 10.6151
R1194 B.n550 B.n132 10.6151
R1195 B.n560 B.n132 10.6151
R1196 B.n561 B.n560 10.6151
R1197 B.n562 B.n561 10.6151
R1198 B.n562 B.n124 10.6151
R1199 B.n573 B.n124 10.6151
R1200 B.n574 B.n573 10.6151
R1201 B.n575 B.n574 10.6151
R1202 B.n575 B.n0 10.6151
R1203 B.n513 B.n512 10.6151
R1204 B.n512 B.n164 10.6151
R1205 B.n507 B.n164 10.6151
R1206 B.n507 B.n506 10.6151
R1207 B.n506 B.n166 10.6151
R1208 B.n501 B.n166 10.6151
R1209 B.n501 B.n500 10.6151
R1210 B.n500 B.n499 10.6151
R1211 B.n499 B.n168 10.6151
R1212 B.n493 B.n168 10.6151
R1213 B.n493 B.n492 10.6151
R1214 B.n492 B.n491 10.6151
R1215 B.n491 B.n170 10.6151
R1216 B.n485 B.n170 10.6151
R1217 B.n485 B.n484 10.6151
R1218 B.n484 B.n483 10.6151
R1219 B.n483 B.n172 10.6151
R1220 B.n477 B.n172 10.6151
R1221 B.n477 B.n476 10.6151
R1222 B.n476 B.n475 10.6151
R1223 B.n475 B.n174 10.6151
R1224 B.n469 B.n174 10.6151
R1225 B.n469 B.n468 10.6151
R1226 B.n468 B.n467 10.6151
R1227 B.n467 B.n176 10.6151
R1228 B.n461 B.n176 10.6151
R1229 B.n461 B.n460 10.6151
R1230 B.n460 B.n459 10.6151
R1231 B.n459 B.n178 10.6151
R1232 B.n453 B.n178 10.6151
R1233 B.n453 B.n452 10.6151
R1234 B.n452 B.n451 10.6151
R1235 B.n451 B.n180 10.6151
R1236 B.n445 B.n180 10.6151
R1237 B.n445 B.n444 10.6151
R1238 B.n444 B.n443 10.6151
R1239 B.n443 B.n182 10.6151
R1240 B.n437 B.n182 10.6151
R1241 B.n437 B.n436 10.6151
R1242 B.n436 B.n435 10.6151
R1243 B.n435 B.n184 10.6151
R1244 B.n429 B.n184 10.6151
R1245 B.n429 B.n428 10.6151
R1246 B.n428 B.n427 10.6151
R1247 B.n427 B.n186 10.6151
R1248 B.n421 B.n186 10.6151
R1249 B.n421 B.n420 10.6151
R1250 B.n420 B.n419 10.6151
R1251 B.n419 B.n188 10.6151
R1252 B.n413 B.n188 10.6151
R1253 B.n413 B.n412 10.6151
R1254 B.n412 B.n411 10.6151
R1255 B.n411 B.n190 10.6151
R1256 B.n405 B.n190 10.6151
R1257 B.n405 B.n404 10.6151
R1258 B.n404 B.n403 10.6151
R1259 B.n403 B.n192 10.6151
R1260 B.n397 B.n192 10.6151
R1261 B.n397 B.n396 10.6151
R1262 B.n396 B.n395 10.6151
R1263 B.n395 B.n194 10.6151
R1264 B.n389 B.n194 10.6151
R1265 B.n389 B.n388 10.6151
R1266 B.n388 B.n387 10.6151
R1267 B.n383 B.n382 10.6151
R1268 B.n382 B.n200 10.6151
R1269 B.n377 B.n200 10.6151
R1270 B.n377 B.n376 10.6151
R1271 B.n376 B.n375 10.6151
R1272 B.n375 B.n202 10.6151
R1273 B.n369 B.n202 10.6151
R1274 B.n369 B.n368 10.6151
R1275 B.n366 B.n206 10.6151
R1276 B.n360 B.n206 10.6151
R1277 B.n360 B.n359 10.6151
R1278 B.n359 B.n358 10.6151
R1279 B.n358 B.n208 10.6151
R1280 B.n352 B.n208 10.6151
R1281 B.n352 B.n351 10.6151
R1282 B.n351 B.n350 10.6151
R1283 B.n350 B.n210 10.6151
R1284 B.n344 B.n210 10.6151
R1285 B.n344 B.n343 10.6151
R1286 B.n343 B.n342 10.6151
R1287 B.n342 B.n212 10.6151
R1288 B.n336 B.n212 10.6151
R1289 B.n336 B.n335 10.6151
R1290 B.n335 B.n334 10.6151
R1291 B.n334 B.n214 10.6151
R1292 B.n328 B.n214 10.6151
R1293 B.n328 B.n327 10.6151
R1294 B.n327 B.n326 10.6151
R1295 B.n326 B.n216 10.6151
R1296 B.n320 B.n216 10.6151
R1297 B.n320 B.n319 10.6151
R1298 B.n319 B.n318 10.6151
R1299 B.n318 B.n218 10.6151
R1300 B.n312 B.n218 10.6151
R1301 B.n312 B.n311 10.6151
R1302 B.n311 B.n310 10.6151
R1303 B.n310 B.n220 10.6151
R1304 B.n304 B.n220 10.6151
R1305 B.n304 B.n303 10.6151
R1306 B.n303 B.n302 10.6151
R1307 B.n302 B.n222 10.6151
R1308 B.n296 B.n222 10.6151
R1309 B.n296 B.n295 10.6151
R1310 B.n295 B.n294 10.6151
R1311 B.n294 B.n224 10.6151
R1312 B.n288 B.n224 10.6151
R1313 B.n288 B.n287 10.6151
R1314 B.n287 B.n286 10.6151
R1315 B.n286 B.n226 10.6151
R1316 B.n280 B.n226 10.6151
R1317 B.n280 B.n279 10.6151
R1318 B.n279 B.n278 10.6151
R1319 B.n278 B.n228 10.6151
R1320 B.n272 B.n228 10.6151
R1321 B.n272 B.n271 10.6151
R1322 B.n271 B.n270 10.6151
R1323 B.n270 B.n230 10.6151
R1324 B.n264 B.n230 10.6151
R1325 B.n264 B.n263 10.6151
R1326 B.n263 B.n262 10.6151
R1327 B.n262 B.n232 10.6151
R1328 B.n256 B.n232 10.6151
R1329 B.n256 B.n255 10.6151
R1330 B.n255 B.n254 10.6151
R1331 B.n254 B.n234 10.6151
R1332 B.n248 B.n234 10.6151
R1333 B.n248 B.n247 10.6151
R1334 B.n247 B.n246 10.6151
R1335 B.n246 B.n236 10.6151
R1336 B.n240 B.n236 10.6151
R1337 B.n240 B.n239 10.6151
R1338 B.n239 B.n160 10.6151
R1339 B.n519 B.n518 10.6151
R1340 B.n520 B.n519 10.6151
R1341 B.n520 B.n152 10.6151
R1342 B.n530 B.n152 10.6151
R1343 B.n531 B.n530 10.6151
R1344 B.n532 B.n531 10.6151
R1345 B.n532 B.n144 10.6151
R1346 B.n542 B.n144 10.6151
R1347 B.n543 B.n542 10.6151
R1348 B.n544 B.n543 10.6151
R1349 B.n544 B.n136 10.6151
R1350 B.n554 B.n136 10.6151
R1351 B.n555 B.n554 10.6151
R1352 B.n556 B.n555 10.6151
R1353 B.n556 B.n127 10.6151
R1354 B.n566 B.n127 10.6151
R1355 B.n567 B.n566 10.6151
R1356 B.n569 B.n567 10.6151
R1357 B.n569 B.n568 10.6151
R1358 B.n568 B.n120 10.6151
R1359 B.n580 B.n120 10.6151
R1360 B.n581 B.n580 10.6151
R1361 B.n582 B.n581 10.6151
R1362 B.n583 B.n582 10.6151
R1363 B.n584 B.n583 10.6151
R1364 B.n587 B.n584 10.6151
R1365 B.n588 B.n587 10.6151
R1366 B.n589 B.n588 10.6151
R1367 B.n590 B.n589 10.6151
R1368 B.n592 B.n590 10.6151
R1369 B.n593 B.n592 10.6151
R1370 B.n594 B.n593 10.6151
R1371 B.n595 B.n594 10.6151
R1372 B.n597 B.n595 10.6151
R1373 B.n598 B.n597 10.6151
R1374 B.n599 B.n598 10.6151
R1375 B.n600 B.n599 10.6151
R1376 B.n602 B.n600 10.6151
R1377 B.n603 B.n602 10.6151
R1378 B.n604 B.n603 10.6151
R1379 B.n605 B.n604 10.6151
R1380 B.n607 B.n605 10.6151
R1381 B.n608 B.n607 10.6151
R1382 B.n609 B.n608 10.6151
R1383 B.n610 B.n609 10.6151
R1384 B.n929 B.n1 10.6151
R1385 B.n929 B.n928 10.6151
R1386 B.n928 B.n927 10.6151
R1387 B.n927 B.n10 10.6151
R1388 B.n921 B.n10 10.6151
R1389 B.n921 B.n920 10.6151
R1390 B.n920 B.n919 10.6151
R1391 B.n919 B.n18 10.6151
R1392 B.n913 B.n18 10.6151
R1393 B.n913 B.n912 10.6151
R1394 B.n912 B.n911 10.6151
R1395 B.n911 B.n25 10.6151
R1396 B.n905 B.n25 10.6151
R1397 B.n905 B.n904 10.6151
R1398 B.n904 B.n903 10.6151
R1399 B.n903 B.n32 10.6151
R1400 B.n897 B.n32 10.6151
R1401 B.n897 B.n896 10.6151
R1402 B.n896 B.n895 10.6151
R1403 B.n895 B.n39 10.6151
R1404 B.n889 B.n39 10.6151
R1405 B.n888 B.n887 10.6151
R1406 B.n887 B.n46 10.6151
R1407 B.n881 B.n46 10.6151
R1408 B.n881 B.n880 10.6151
R1409 B.n880 B.n879 10.6151
R1410 B.n879 B.n48 10.6151
R1411 B.n873 B.n48 10.6151
R1412 B.n873 B.n872 10.6151
R1413 B.n872 B.n871 10.6151
R1414 B.n871 B.n50 10.6151
R1415 B.n865 B.n50 10.6151
R1416 B.n865 B.n864 10.6151
R1417 B.n864 B.n863 10.6151
R1418 B.n863 B.n52 10.6151
R1419 B.n857 B.n52 10.6151
R1420 B.n857 B.n856 10.6151
R1421 B.n856 B.n855 10.6151
R1422 B.n855 B.n54 10.6151
R1423 B.n849 B.n54 10.6151
R1424 B.n849 B.n848 10.6151
R1425 B.n848 B.n847 10.6151
R1426 B.n847 B.n56 10.6151
R1427 B.n841 B.n56 10.6151
R1428 B.n841 B.n840 10.6151
R1429 B.n840 B.n839 10.6151
R1430 B.n839 B.n58 10.6151
R1431 B.n833 B.n58 10.6151
R1432 B.n833 B.n832 10.6151
R1433 B.n832 B.n831 10.6151
R1434 B.n831 B.n60 10.6151
R1435 B.n825 B.n60 10.6151
R1436 B.n825 B.n824 10.6151
R1437 B.n824 B.n823 10.6151
R1438 B.n823 B.n62 10.6151
R1439 B.n817 B.n62 10.6151
R1440 B.n817 B.n816 10.6151
R1441 B.n816 B.n815 10.6151
R1442 B.n815 B.n64 10.6151
R1443 B.n809 B.n64 10.6151
R1444 B.n809 B.n808 10.6151
R1445 B.n808 B.n807 10.6151
R1446 B.n807 B.n66 10.6151
R1447 B.n801 B.n66 10.6151
R1448 B.n801 B.n800 10.6151
R1449 B.n800 B.n799 10.6151
R1450 B.n799 B.n68 10.6151
R1451 B.n793 B.n68 10.6151
R1452 B.n793 B.n792 10.6151
R1453 B.n792 B.n791 10.6151
R1454 B.n791 B.n70 10.6151
R1455 B.n785 B.n70 10.6151
R1456 B.n785 B.n784 10.6151
R1457 B.n784 B.n783 10.6151
R1458 B.n783 B.n72 10.6151
R1459 B.n777 B.n72 10.6151
R1460 B.n777 B.n776 10.6151
R1461 B.n776 B.n775 10.6151
R1462 B.n775 B.n74 10.6151
R1463 B.n769 B.n74 10.6151
R1464 B.n769 B.n768 10.6151
R1465 B.n768 B.n767 10.6151
R1466 B.n767 B.n76 10.6151
R1467 B.n761 B.n76 10.6151
R1468 B.n761 B.n760 10.6151
R1469 B.n758 B.n80 10.6151
R1470 B.n752 B.n80 10.6151
R1471 B.n752 B.n751 10.6151
R1472 B.n751 B.n750 10.6151
R1473 B.n750 B.n82 10.6151
R1474 B.n744 B.n82 10.6151
R1475 B.n744 B.n743 10.6151
R1476 B.n743 B.n742 10.6151
R1477 B.n738 B.n737 10.6151
R1478 B.n737 B.n88 10.6151
R1479 B.n732 B.n88 10.6151
R1480 B.n732 B.n731 10.6151
R1481 B.n731 B.n730 10.6151
R1482 B.n730 B.n90 10.6151
R1483 B.n724 B.n90 10.6151
R1484 B.n724 B.n723 10.6151
R1485 B.n723 B.n722 10.6151
R1486 B.n722 B.n92 10.6151
R1487 B.n716 B.n92 10.6151
R1488 B.n716 B.n715 10.6151
R1489 B.n715 B.n714 10.6151
R1490 B.n714 B.n94 10.6151
R1491 B.n708 B.n94 10.6151
R1492 B.n708 B.n707 10.6151
R1493 B.n707 B.n706 10.6151
R1494 B.n706 B.n96 10.6151
R1495 B.n700 B.n96 10.6151
R1496 B.n700 B.n699 10.6151
R1497 B.n699 B.n698 10.6151
R1498 B.n698 B.n98 10.6151
R1499 B.n692 B.n98 10.6151
R1500 B.n692 B.n691 10.6151
R1501 B.n691 B.n690 10.6151
R1502 B.n690 B.n100 10.6151
R1503 B.n684 B.n100 10.6151
R1504 B.n684 B.n683 10.6151
R1505 B.n683 B.n682 10.6151
R1506 B.n682 B.n102 10.6151
R1507 B.n676 B.n102 10.6151
R1508 B.n676 B.n675 10.6151
R1509 B.n675 B.n674 10.6151
R1510 B.n674 B.n104 10.6151
R1511 B.n668 B.n104 10.6151
R1512 B.n668 B.n667 10.6151
R1513 B.n667 B.n666 10.6151
R1514 B.n666 B.n106 10.6151
R1515 B.n660 B.n106 10.6151
R1516 B.n660 B.n659 10.6151
R1517 B.n659 B.n658 10.6151
R1518 B.n658 B.n108 10.6151
R1519 B.n652 B.n108 10.6151
R1520 B.n652 B.n651 10.6151
R1521 B.n651 B.n650 10.6151
R1522 B.n650 B.n110 10.6151
R1523 B.n644 B.n110 10.6151
R1524 B.n644 B.n643 10.6151
R1525 B.n643 B.n642 10.6151
R1526 B.n642 B.n112 10.6151
R1527 B.n636 B.n112 10.6151
R1528 B.n636 B.n635 10.6151
R1529 B.n635 B.n634 10.6151
R1530 B.n634 B.n114 10.6151
R1531 B.n628 B.n114 10.6151
R1532 B.n628 B.n627 10.6151
R1533 B.n627 B.n626 10.6151
R1534 B.n626 B.n116 10.6151
R1535 B.n620 B.n116 10.6151
R1536 B.n620 B.n619 10.6151
R1537 B.n619 B.n618 10.6151
R1538 B.n618 B.n118 10.6151
R1539 B.n612 B.n118 10.6151
R1540 B.n612 B.n611 10.6151
R1541 B.n937 B.n0 8.11757
R1542 B.n937 B.n1 8.11757
R1543 B.t3 B.n146 7.44329
R1544 B.n130 B.t0 7.44329
R1545 B.t1 B.n924 7.44329
R1546 B.t10 B.n30 7.44329
R1547 B.n383 B.n198 6.5566
R1548 B.n368 B.n367 6.5566
R1549 B.n759 B.n758 6.5566
R1550 B.n742 B.n86 6.5566
R1551 B.n387 B.n198 4.05904
R1552 B.n367 B.n366 4.05904
R1553 B.n760 B.n759 4.05904
R1554 B.n738 B.n86 4.05904
R1555 VN VN.t1 321.183
R1556 VN VN.t0 272.012
R1557 VTAIL.n1 VTAIL.t3 47.8205
R1558 VTAIL.n3 VTAIL.t2 47.8203
R1559 VTAIL.n0 VTAIL.t0 47.8203
R1560 VTAIL.n2 VTAIL.t1 47.8203
R1561 VTAIL.n1 VTAIL.n0 33.7548
R1562 VTAIL.n3 VTAIL.n2 31.6169
R1563 VTAIL.n2 VTAIL.n1 1.53929
R1564 VTAIL VTAIL.n0 1.063
R1565 VTAIL VTAIL.n3 0.476793
R1566 VDD2.n0 VDD2.t1 109.546
R1567 VDD2.n0 VDD2.t0 64.4991
R1568 VDD2 VDD2.n0 0.593172
R1569 VP.n0 VP.t0 321.086
R1570 VP.n0 VP.t1 271.675
R1571 VP VP.n0 0.336784
R1572 VDD1 VDD1.t0 110.606
R1573 VDD1 VDD1.t1 65.0918
C0 VDD1 VDD2 0.622057f
C1 VTAIL VN 3.56921f
C2 VDD1 VTAIL 7.17381f
C3 VDD1 VN 0.147916f
C4 VP VDD2 0.31491f
C5 VP VTAIL 3.58369f
C6 VTAIL VDD2 7.21868f
C7 VP VN 6.70186f
C8 VN VDD2 4.29494f
C9 VDD1 VP 4.45756f
C10 VDD2 B 5.683325f
C11 VDD1 B 9.32608f
C12 VTAIL B 10.284379f
C13 VN B 12.26303f
C14 VP B 6.382174f
C15 VDD1.t1 B 3.69073f
C16 VDD1.t0 B 4.45f
C17 VP.t0 B 4.70046f
C18 VP.t1 B 4.21169f
C19 VP.n0 B 5.821681f
C20 VDD2.t1 B 4.36521f
C21 VDD2.t0 B 3.64841f
C22 VDD2.n0 B 3.37962f
C23 VTAIL.t0 B 3.51111f
C24 VTAIL.n0 B 1.92609f
C25 VTAIL.t3 B 3.51111f
C26 VTAIL.n1 B 1.95598f
C27 VTAIL.t1 B 3.51111f
C28 VTAIL.n2 B 1.8218f
C29 VTAIL.t2 B 3.51111f
C30 VTAIL.n3 B 1.75512f
C31 VN.t0 B 4.14332f
C32 VN.t1 B 4.62475f
.ends

