* NGSPICE file created from diff_pair_sample_1602.ext - technology: sky130A

.subckt diff_pair_sample_1602 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0 ps=0 w=3.62 l=1.42
X1 VDD1.t5 VP.t0 VTAIL.t10 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0.5973 ps=3.95 w=3.62 l=1.42
X2 VTAIL.t7 VP.t1 VDD1.t4 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=0.5973 ps=3.95 w=3.62 l=1.42
X3 VTAIL.t4 VN.t0 VDD2.t5 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=0.5973 ps=3.95 w=3.62 l=1.42
X4 VDD2.t4 VN.t1 VTAIL.t11 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0.5973 ps=3.95 w=3.62 l=1.42
X5 VDD2.t3 VN.t2 VTAIL.t0 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=1.4118 ps=8.02 w=3.62 l=1.42
X6 VDD2.t2 VN.t3 VTAIL.t1 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=1.4118 ps=8.02 w=3.62 l=1.42
X7 VDD1.t3 VP.t2 VTAIL.t6 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=1.4118 ps=8.02 w=3.62 l=1.42
X8 VTAIL.t5 VP.t3 VDD1.t2 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=0.5973 ps=3.95 w=3.62 l=1.42
X9 VTAIL.t3 VN.t4 VDD2.t1 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=0.5973 ps=3.95 w=3.62 l=1.42
X10 VDD1.t1 VP.t4 VTAIL.t8 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0.5973 ps=3.95 w=3.62 l=1.42
X11 B.t8 B.t6 B.t7 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0 ps=0 w=3.62 l=1.42
X12 VDD1.t0 VP.t5 VTAIL.t9 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=0.5973 pd=3.95 as=1.4118 ps=8.02 w=3.62 l=1.42
X13 B.t5 B.t3 B.t4 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0 ps=0 w=3.62 l=1.42
X14 B.t2 B.t0 B.t1 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0 ps=0 w=3.62 l=1.42
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n2370_n1692# sky130_fd_pr__pfet_01v8 ad=1.4118 pd=8.02 as=0.5973 ps=3.95 w=3.62 l=1.42
R0 B.n219 B.n72 585
R1 B.n218 B.n217 585
R2 B.n216 B.n73 585
R3 B.n215 B.n214 585
R4 B.n213 B.n74 585
R5 B.n212 B.n211 585
R6 B.n210 B.n75 585
R7 B.n209 B.n208 585
R8 B.n207 B.n76 585
R9 B.n206 B.n205 585
R10 B.n204 B.n77 585
R11 B.n203 B.n202 585
R12 B.n201 B.n78 585
R13 B.n200 B.n199 585
R14 B.n198 B.n79 585
R15 B.n197 B.n196 585
R16 B.n195 B.n80 585
R17 B.n193 B.n192 585
R18 B.n191 B.n83 585
R19 B.n190 B.n189 585
R20 B.n188 B.n84 585
R21 B.n187 B.n186 585
R22 B.n185 B.n85 585
R23 B.n184 B.n183 585
R24 B.n182 B.n86 585
R25 B.n181 B.n180 585
R26 B.n179 B.n87 585
R27 B.n178 B.n177 585
R28 B.n173 B.n88 585
R29 B.n172 B.n171 585
R30 B.n170 B.n89 585
R31 B.n169 B.n168 585
R32 B.n167 B.n90 585
R33 B.n166 B.n165 585
R34 B.n164 B.n91 585
R35 B.n163 B.n162 585
R36 B.n161 B.n92 585
R37 B.n160 B.n159 585
R38 B.n158 B.n93 585
R39 B.n157 B.n156 585
R40 B.n155 B.n94 585
R41 B.n154 B.n153 585
R42 B.n152 B.n95 585
R43 B.n151 B.n150 585
R44 B.n221 B.n220 585
R45 B.n222 B.n71 585
R46 B.n224 B.n223 585
R47 B.n225 B.n70 585
R48 B.n227 B.n226 585
R49 B.n228 B.n69 585
R50 B.n230 B.n229 585
R51 B.n231 B.n68 585
R52 B.n233 B.n232 585
R53 B.n234 B.n67 585
R54 B.n236 B.n235 585
R55 B.n237 B.n66 585
R56 B.n239 B.n238 585
R57 B.n240 B.n65 585
R58 B.n242 B.n241 585
R59 B.n243 B.n64 585
R60 B.n245 B.n244 585
R61 B.n246 B.n63 585
R62 B.n248 B.n247 585
R63 B.n249 B.n62 585
R64 B.n251 B.n250 585
R65 B.n252 B.n61 585
R66 B.n254 B.n253 585
R67 B.n255 B.n60 585
R68 B.n257 B.n256 585
R69 B.n258 B.n59 585
R70 B.n260 B.n259 585
R71 B.n261 B.n58 585
R72 B.n263 B.n262 585
R73 B.n264 B.n57 585
R74 B.n266 B.n265 585
R75 B.n267 B.n56 585
R76 B.n269 B.n268 585
R77 B.n270 B.n55 585
R78 B.n272 B.n271 585
R79 B.n273 B.n54 585
R80 B.n275 B.n274 585
R81 B.n276 B.n53 585
R82 B.n278 B.n277 585
R83 B.n279 B.n52 585
R84 B.n281 B.n280 585
R85 B.n282 B.n51 585
R86 B.n284 B.n283 585
R87 B.n285 B.n50 585
R88 B.n287 B.n286 585
R89 B.n288 B.n49 585
R90 B.n290 B.n289 585
R91 B.n291 B.n48 585
R92 B.n293 B.n292 585
R93 B.n294 B.n47 585
R94 B.n296 B.n295 585
R95 B.n297 B.n46 585
R96 B.n299 B.n298 585
R97 B.n300 B.n45 585
R98 B.n302 B.n301 585
R99 B.n303 B.n44 585
R100 B.n305 B.n304 585
R101 B.n306 B.n43 585
R102 B.n373 B.n16 585
R103 B.n372 B.n371 585
R104 B.n370 B.n17 585
R105 B.n369 B.n368 585
R106 B.n367 B.n18 585
R107 B.n366 B.n365 585
R108 B.n364 B.n19 585
R109 B.n363 B.n362 585
R110 B.n361 B.n20 585
R111 B.n360 B.n359 585
R112 B.n358 B.n21 585
R113 B.n357 B.n356 585
R114 B.n355 B.n22 585
R115 B.n354 B.n353 585
R116 B.n352 B.n23 585
R117 B.n351 B.n350 585
R118 B.n349 B.n24 585
R119 B.n348 B.n347 585
R120 B.n346 B.n25 585
R121 B.n345 B.n344 585
R122 B.n343 B.n29 585
R123 B.n342 B.n341 585
R124 B.n340 B.n30 585
R125 B.n339 B.n338 585
R126 B.n337 B.n31 585
R127 B.n336 B.n335 585
R128 B.n334 B.n32 585
R129 B.n332 B.n331 585
R130 B.n330 B.n35 585
R131 B.n329 B.n328 585
R132 B.n327 B.n36 585
R133 B.n326 B.n325 585
R134 B.n324 B.n37 585
R135 B.n323 B.n322 585
R136 B.n321 B.n38 585
R137 B.n320 B.n319 585
R138 B.n318 B.n39 585
R139 B.n317 B.n316 585
R140 B.n315 B.n40 585
R141 B.n314 B.n313 585
R142 B.n312 B.n41 585
R143 B.n311 B.n310 585
R144 B.n309 B.n42 585
R145 B.n308 B.n307 585
R146 B.n375 B.n374 585
R147 B.n376 B.n15 585
R148 B.n378 B.n377 585
R149 B.n379 B.n14 585
R150 B.n381 B.n380 585
R151 B.n382 B.n13 585
R152 B.n384 B.n383 585
R153 B.n385 B.n12 585
R154 B.n387 B.n386 585
R155 B.n388 B.n11 585
R156 B.n390 B.n389 585
R157 B.n391 B.n10 585
R158 B.n393 B.n392 585
R159 B.n394 B.n9 585
R160 B.n396 B.n395 585
R161 B.n397 B.n8 585
R162 B.n399 B.n398 585
R163 B.n400 B.n7 585
R164 B.n402 B.n401 585
R165 B.n403 B.n6 585
R166 B.n405 B.n404 585
R167 B.n406 B.n5 585
R168 B.n408 B.n407 585
R169 B.n409 B.n4 585
R170 B.n411 B.n410 585
R171 B.n412 B.n3 585
R172 B.n414 B.n413 585
R173 B.n415 B.n0 585
R174 B.n2 B.n1 585
R175 B.n110 B.n109 585
R176 B.n112 B.n111 585
R177 B.n113 B.n108 585
R178 B.n115 B.n114 585
R179 B.n116 B.n107 585
R180 B.n118 B.n117 585
R181 B.n119 B.n106 585
R182 B.n121 B.n120 585
R183 B.n122 B.n105 585
R184 B.n124 B.n123 585
R185 B.n125 B.n104 585
R186 B.n127 B.n126 585
R187 B.n128 B.n103 585
R188 B.n130 B.n129 585
R189 B.n131 B.n102 585
R190 B.n133 B.n132 585
R191 B.n134 B.n101 585
R192 B.n136 B.n135 585
R193 B.n137 B.n100 585
R194 B.n139 B.n138 585
R195 B.n140 B.n99 585
R196 B.n142 B.n141 585
R197 B.n143 B.n98 585
R198 B.n145 B.n144 585
R199 B.n146 B.n97 585
R200 B.n148 B.n147 585
R201 B.n149 B.n96 585
R202 B.n151 B.n96 492.5
R203 B.n221 B.n72 492.5
R204 B.n307 B.n306 492.5
R205 B.n374 B.n373 492.5
R206 B.n174 B.t0 266.567
R207 B.n81 B.t3 266.567
R208 B.n33 B.t6 266.567
R209 B.n26 B.t9 266.567
R210 B.n417 B.n416 256.663
R211 B.n416 B.n415 235.042
R212 B.n416 B.n2 235.042
R213 B.n81 B.t4 164.254
R214 B.n33 B.t8 164.254
R215 B.n174 B.t1 164.251
R216 B.n26 B.t11 164.251
R217 B.n152 B.n151 163.367
R218 B.n153 B.n152 163.367
R219 B.n153 B.n94 163.367
R220 B.n157 B.n94 163.367
R221 B.n158 B.n157 163.367
R222 B.n159 B.n158 163.367
R223 B.n159 B.n92 163.367
R224 B.n163 B.n92 163.367
R225 B.n164 B.n163 163.367
R226 B.n165 B.n164 163.367
R227 B.n165 B.n90 163.367
R228 B.n169 B.n90 163.367
R229 B.n170 B.n169 163.367
R230 B.n171 B.n170 163.367
R231 B.n171 B.n88 163.367
R232 B.n178 B.n88 163.367
R233 B.n179 B.n178 163.367
R234 B.n180 B.n179 163.367
R235 B.n180 B.n86 163.367
R236 B.n184 B.n86 163.367
R237 B.n185 B.n184 163.367
R238 B.n186 B.n185 163.367
R239 B.n186 B.n84 163.367
R240 B.n190 B.n84 163.367
R241 B.n191 B.n190 163.367
R242 B.n192 B.n191 163.367
R243 B.n192 B.n80 163.367
R244 B.n197 B.n80 163.367
R245 B.n198 B.n197 163.367
R246 B.n199 B.n198 163.367
R247 B.n199 B.n78 163.367
R248 B.n203 B.n78 163.367
R249 B.n204 B.n203 163.367
R250 B.n205 B.n204 163.367
R251 B.n205 B.n76 163.367
R252 B.n209 B.n76 163.367
R253 B.n210 B.n209 163.367
R254 B.n211 B.n210 163.367
R255 B.n211 B.n74 163.367
R256 B.n215 B.n74 163.367
R257 B.n216 B.n215 163.367
R258 B.n217 B.n216 163.367
R259 B.n217 B.n72 163.367
R260 B.n306 B.n305 163.367
R261 B.n305 B.n44 163.367
R262 B.n301 B.n44 163.367
R263 B.n301 B.n300 163.367
R264 B.n300 B.n299 163.367
R265 B.n299 B.n46 163.367
R266 B.n295 B.n46 163.367
R267 B.n295 B.n294 163.367
R268 B.n294 B.n293 163.367
R269 B.n293 B.n48 163.367
R270 B.n289 B.n48 163.367
R271 B.n289 B.n288 163.367
R272 B.n288 B.n287 163.367
R273 B.n287 B.n50 163.367
R274 B.n283 B.n50 163.367
R275 B.n283 B.n282 163.367
R276 B.n282 B.n281 163.367
R277 B.n281 B.n52 163.367
R278 B.n277 B.n52 163.367
R279 B.n277 B.n276 163.367
R280 B.n276 B.n275 163.367
R281 B.n275 B.n54 163.367
R282 B.n271 B.n54 163.367
R283 B.n271 B.n270 163.367
R284 B.n270 B.n269 163.367
R285 B.n269 B.n56 163.367
R286 B.n265 B.n56 163.367
R287 B.n265 B.n264 163.367
R288 B.n264 B.n263 163.367
R289 B.n263 B.n58 163.367
R290 B.n259 B.n58 163.367
R291 B.n259 B.n258 163.367
R292 B.n258 B.n257 163.367
R293 B.n257 B.n60 163.367
R294 B.n253 B.n60 163.367
R295 B.n253 B.n252 163.367
R296 B.n252 B.n251 163.367
R297 B.n251 B.n62 163.367
R298 B.n247 B.n62 163.367
R299 B.n247 B.n246 163.367
R300 B.n246 B.n245 163.367
R301 B.n245 B.n64 163.367
R302 B.n241 B.n64 163.367
R303 B.n241 B.n240 163.367
R304 B.n240 B.n239 163.367
R305 B.n239 B.n66 163.367
R306 B.n235 B.n66 163.367
R307 B.n235 B.n234 163.367
R308 B.n234 B.n233 163.367
R309 B.n233 B.n68 163.367
R310 B.n229 B.n68 163.367
R311 B.n229 B.n228 163.367
R312 B.n228 B.n227 163.367
R313 B.n227 B.n70 163.367
R314 B.n223 B.n70 163.367
R315 B.n223 B.n222 163.367
R316 B.n222 B.n221 163.367
R317 B.n373 B.n372 163.367
R318 B.n372 B.n17 163.367
R319 B.n368 B.n17 163.367
R320 B.n368 B.n367 163.367
R321 B.n367 B.n366 163.367
R322 B.n366 B.n19 163.367
R323 B.n362 B.n19 163.367
R324 B.n362 B.n361 163.367
R325 B.n361 B.n360 163.367
R326 B.n360 B.n21 163.367
R327 B.n356 B.n21 163.367
R328 B.n356 B.n355 163.367
R329 B.n355 B.n354 163.367
R330 B.n354 B.n23 163.367
R331 B.n350 B.n23 163.367
R332 B.n350 B.n349 163.367
R333 B.n349 B.n348 163.367
R334 B.n348 B.n25 163.367
R335 B.n344 B.n25 163.367
R336 B.n344 B.n343 163.367
R337 B.n343 B.n342 163.367
R338 B.n342 B.n30 163.367
R339 B.n338 B.n30 163.367
R340 B.n338 B.n337 163.367
R341 B.n337 B.n336 163.367
R342 B.n336 B.n32 163.367
R343 B.n331 B.n32 163.367
R344 B.n331 B.n330 163.367
R345 B.n330 B.n329 163.367
R346 B.n329 B.n36 163.367
R347 B.n325 B.n36 163.367
R348 B.n325 B.n324 163.367
R349 B.n324 B.n323 163.367
R350 B.n323 B.n38 163.367
R351 B.n319 B.n38 163.367
R352 B.n319 B.n318 163.367
R353 B.n318 B.n317 163.367
R354 B.n317 B.n40 163.367
R355 B.n313 B.n40 163.367
R356 B.n313 B.n312 163.367
R357 B.n312 B.n311 163.367
R358 B.n311 B.n42 163.367
R359 B.n307 B.n42 163.367
R360 B.n374 B.n15 163.367
R361 B.n378 B.n15 163.367
R362 B.n379 B.n378 163.367
R363 B.n380 B.n379 163.367
R364 B.n380 B.n13 163.367
R365 B.n384 B.n13 163.367
R366 B.n385 B.n384 163.367
R367 B.n386 B.n385 163.367
R368 B.n386 B.n11 163.367
R369 B.n390 B.n11 163.367
R370 B.n391 B.n390 163.367
R371 B.n392 B.n391 163.367
R372 B.n392 B.n9 163.367
R373 B.n396 B.n9 163.367
R374 B.n397 B.n396 163.367
R375 B.n398 B.n397 163.367
R376 B.n398 B.n7 163.367
R377 B.n402 B.n7 163.367
R378 B.n403 B.n402 163.367
R379 B.n404 B.n403 163.367
R380 B.n404 B.n5 163.367
R381 B.n408 B.n5 163.367
R382 B.n409 B.n408 163.367
R383 B.n410 B.n409 163.367
R384 B.n410 B.n3 163.367
R385 B.n414 B.n3 163.367
R386 B.n415 B.n414 163.367
R387 B.n110 B.n2 163.367
R388 B.n111 B.n110 163.367
R389 B.n111 B.n108 163.367
R390 B.n115 B.n108 163.367
R391 B.n116 B.n115 163.367
R392 B.n117 B.n116 163.367
R393 B.n117 B.n106 163.367
R394 B.n121 B.n106 163.367
R395 B.n122 B.n121 163.367
R396 B.n123 B.n122 163.367
R397 B.n123 B.n104 163.367
R398 B.n127 B.n104 163.367
R399 B.n128 B.n127 163.367
R400 B.n129 B.n128 163.367
R401 B.n129 B.n102 163.367
R402 B.n133 B.n102 163.367
R403 B.n134 B.n133 163.367
R404 B.n135 B.n134 163.367
R405 B.n135 B.n100 163.367
R406 B.n139 B.n100 163.367
R407 B.n140 B.n139 163.367
R408 B.n141 B.n140 163.367
R409 B.n141 B.n98 163.367
R410 B.n145 B.n98 163.367
R411 B.n146 B.n145 163.367
R412 B.n147 B.n146 163.367
R413 B.n147 B.n96 163.367
R414 B.n82 B.t5 130.315
R415 B.n34 B.t7 130.315
R416 B.n175 B.t2 130.311
R417 B.n27 B.t10 130.311
R418 B.n176 B.n175 59.5399
R419 B.n194 B.n82 59.5399
R420 B.n333 B.n34 59.5399
R421 B.n28 B.n27 59.5399
R422 B.n175 B.n174 33.9399
R423 B.n82 B.n81 33.9399
R424 B.n34 B.n33 33.9399
R425 B.n27 B.n26 33.9399
R426 B.n375 B.n16 32.0005
R427 B.n308 B.n43 32.0005
R428 B.n220 B.n219 32.0005
R429 B.n150 B.n149 32.0005
R430 B B.n417 18.0485
R431 B.n376 B.n375 10.6151
R432 B.n377 B.n376 10.6151
R433 B.n377 B.n14 10.6151
R434 B.n381 B.n14 10.6151
R435 B.n382 B.n381 10.6151
R436 B.n383 B.n382 10.6151
R437 B.n383 B.n12 10.6151
R438 B.n387 B.n12 10.6151
R439 B.n388 B.n387 10.6151
R440 B.n389 B.n388 10.6151
R441 B.n389 B.n10 10.6151
R442 B.n393 B.n10 10.6151
R443 B.n394 B.n393 10.6151
R444 B.n395 B.n394 10.6151
R445 B.n395 B.n8 10.6151
R446 B.n399 B.n8 10.6151
R447 B.n400 B.n399 10.6151
R448 B.n401 B.n400 10.6151
R449 B.n401 B.n6 10.6151
R450 B.n405 B.n6 10.6151
R451 B.n406 B.n405 10.6151
R452 B.n407 B.n406 10.6151
R453 B.n407 B.n4 10.6151
R454 B.n411 B.n4 10.6151
R455 B.n412 B.n411 10.6151
R456 B.n413 B.n412 10.6151
R457 B.n413 B.n0 10.6151
R458 B.n371 B.n16 10.6151
R459 B.n371 B.n370 10.6151
R460 B.n370 B.n369 10.6151
R461 B.n369 B.n18 10.6151
R462 B.n365 B.n18 10.6151
R463 B.n365 B.n364 10.6151
R464 B.n364 B.n363 10.6151
R465 B.n363 B.n20 10.6151
R466 B.n359 B.n20 10.6151
R467 B.n359 B.n358 10.6151
R468 B.n358 B.n357 10.6151
R469 B.n357 B.n22 10.6151
R470 B.n353 B.n22 10.6151
R471 B.n353 B.n352 10.6151
R472 B.n352 B.n351 10.6151
R473 B.n351 B.n24 10.6151
R474 B.n347 B.n346 10.6151
R475 B.n346 B.n345 10.6151
R476 B.n345 B.n29 10.6151
R477 B.n341 B.n29 10.6151
R478 B.n341 B.n340 10.6151
R479 B.n340 B.n339 10.6151
R480 B.n339 B.n31 10.6151
R481 B.n335 B.n31 10.6151
R482 B.n335 B.n334 10.6151
R483 B.n332 B.n35 10.6151
R484 B.n328 B.n35 10.6151
R485 B.n328 B.n327 10.6151
R486 B.n327 B.n326 10.6151
R487 B.n326 B.n37 10.6151
R488 B.n322 B.n37 10.6151
R489 B.n322 B.n321 10.6151
R490 B.n321 B.n320 10.6151
R491 B.n320 B.n39 10.6151
R492 B.n316 B.n39 10.6151
R493 B.n316 B.n315 10.6151
R494 B.n315 B.n314 10.6151
R495 B.n314 B.n41 10.6151
R496 B.n310 B.n41 10.6151
R497 B.n310 B.n309 10.6151
R498 B.n309 B.n308 10.6151
R499 B.n304 B.n43 10.6151
R500 B.n304 B.n303 10.6151
R501 B.n303 B.n302 10.6151
R502 B.n302 B.n45 10.6151
R503 B.n298 B.n45 10.6151
R504 B.n298 B.n297 10.6151
R505 B.n297 B.n296 10.6151
R506 B.n296 B.n47 10.6151
R507 B.n292 B.n47 10.6151
R508 B.n292 B.n291 10.6151
R509 B.n291 B.n290 10.6151
R510 B.n290 B.n49 10.6151
R511 B.n286 B.n49 10.6151
R512 B.n286 B.n285 10.6151
R513 B.n285 B.n284 10.6151
R514 B.n284 B.n51 10.6151
R515 B.n280 B.n51 10.6151
R516 B.n280 B.n279 10.6151
R517 B.n279 B.n278 10.6151
R518 B.n278 B.n53 10.6151
R519 B.n274 B.n53 10.6151
R520 B.n274 B.n273 10.6151
R521 B.n273 B.n272 10.6151
R522 B.n272 B.n55 10.6151
R523 B.n268 B.n55 10.6151
R524 B.n268 B.n267 10.6151
R525 B.n267 B.n266 10.6151
R526 B.n266 B.n57 10.6151
R527 B.n262 B.n57 10.6151
R528 B.n262 B.n261 10.6151
R529 B.n261 B.n260 10.6151
R530 B.n260 B.n59 10.6151
R531 B.n256 B.n59 10.6151
R532 B.n256 B.n255 10.6151
R533 B.n255 B.n254 10.6151
R534 B.n254 B.n61 10.6151
R535 B.n250 B.n61 10.6151
R536 B.n250 B.n249 10.6151
R537 B.n249 B.n248 10.6151
R538 B.n248 B.n63 10.6151
R539 B.n244 B.n63 10.6151
R540 B.n244 B.n243 10.6151
R541 B.n243 B.n242 10.6151
R542 B.n242 B.n65 10.6151
R543 B.n238 B.n65 10.6151
R544 B.n238 B.n237 10.6151
R545 B.n237 B.n236 10.6151
R546 B.n236 B.n67 10.6151
R547 B.n232 B.n67 10.6151
R548 B.n232 B.n231 10.6151
R549 B.n231 B.n230 10.6151
R550 B.n230 B.n69 10.6151
R551 B.n226 B.n69 10.6151
R552 B.n226 B.n225 10.6151
R553 B.n225 B.n224 10.6151
R554 B.n224 B.n71 10.6151
R555 B.n220 B.n71 10.6151
R556 B.n109 B.n1 10.6151
R557 B.n112 B.n109 10.6151
R558 B.n113 B.n112 10.6151
R559 B.n114 B.n113 10.6151
R560 B.n114 B.n107 10.6151
R561 B.n118 B.n107 10.6151
R562 B.n119 B.n118 10.6151
R563 B.n120 B.n119 10.6151
R564 B.n120 B.n105 10.6151
R565 B.n124 B.n105 10.6151
R566 B.n125 B.n124 10.6151
R567 B.n126 B.n125 10.6151
R568 B.n126 B.n103 10.6151
R569 B.n130 B.n103 10.6151
R570 B.n131 B.n130 10.6151
R571 B.n132 B.n131 10.6151
R572 B.n132 B.n101 10.6151
R573 B.n136 B.n101 10.6151
R574 B.n137 B.n136 10.6151
R575 B.n138 B.n137 10.6151
R576 B.n138 B.n99 10.6151
R577 B.n142 B.n99 10.6151
R578 B.n143 B.n142 10.6151
R579 B.n144 B.n143 10.6151
R580 B.n144 B.n97 10.6151
R581 B.n148 B.n97 10.6151
R582 B.n149 B.n148 10.6151
R583 B.n150 B.n95 10.6151
R584 B.n154 B.n95 10.6151
R585 B.n155 B.n154 10.6151
R586 B.n156 B.n155 10.6151
R587 B.n156 B.n93 10.6151
R588 B.n160 B.n93 10.6151
R589 B.n161 B.n160 10.6151
R590 B.n162 B.n161 10.6151
R591 B.n162 B.n91 10.6151
R592 B.n166 B.n91 10.6151
R593 B.n167 B.n166 10.6151
R594 B.n168 B.n167 10.6151
R595 B.n168 B.n89 10.6151
R596 B.n172 B.n89 10.6151
R597 B.n173 B.n172 10.6151
R598 B.n177 B.n173 10.6151
R599 B.n181 B.n87 10.6151
R600 B.n182 B.n181 10.6151
R601 B.n183 B.n182 10.6151
R602 B.n183 B.n85 10.6151
R603 B.n187 B.n85 10.6151
R604 B.n188 B.n187 10.6151
R605 B.n189 B.n188 10.6151
R606 B.n189 B.n83 10.6151
R607 B.n193 B.n83 10.6151
R608 B.n196 B.n195 10.6151
R609 B.n196 B.n79 10.6151
R610 B.n200 B.n79 10.6151
R611 B.n201 B.n200 10.6151
R612 B.n202 B.n201 10.6151
R613 B.n202 B.n77 10.6151
R614 B.n206 B.n77 10.6151
R615 B.n207 B.n206 10.6151
R616 B.n208 B.n207 10.6151
R617 B.n208 B.n75 10.6151
R618 B.n212 B.n75 10.6151
R619 B.n213 B.n212 10.6151
R620 B.n214 B.n213 10.6151
R621 B.n214 B.n73 10.6151
R622 B.n218 B.n73 10.6151
R623 B.n219 B.n218 10.6151
R624 B.n28 B.n24 9.36635
R625 B.n333 B.n332 9.36635
R626 B.n177 B.n176 9.36635
R627 B.n195 B.n194 9.36635
R628 B.n417 B.n0 8.11757
R629 B.n417 B.n1 8.11757
R630 B.n347 B.n28 1.24928
R631 B.n334 B.n333 1.24928
R632 B.n176 B.n87 1.24928
R633 B.n194 B.n193 1.24928
R634 VP.n15 VP.n14 173.596
R635 VP.n27 VP.n26 173.596
R636 VP.n13 VP.n12 173.596
R637 VP.n8 VP.n5 161.3
R638 VP.n10 VP.n9 161.3
R639 VP.n11 VP.n4 161.3
R640 VP.n25 VP.n0 161.3
R641 VP.n24 VP.n23 161.3
R642 VP.n22 VP.n1 161.3
R643 VP.n21 VP.n20 161.3
R644 VP.n19 VP.n2 161.3
R645 VP.n18 VP.n17 161.3
R646 VP.n16 VP.n3 161.3
R647 VP.n7 VP.t4 96.9427
R648 VP.n20 VP.t1 61.4385
R649 VP.n14 VP.t0 61.4385
R650 VP.n26 VP.t5 61.4385
R651 VP.n6 VP.t3 61.4385
R652 VP.n12 VP.t2 61.4385
R653 VP.n19 VP.n18 52.6866
R654 VP.n24 VP.n1 52.6866
R655 VP.n10 VP.n5 52.6866
R656 VP.n7 VP.n6 41.915
R657 VP.n15 VP.n13 37.6407
R658 VP.n18 VP.n3 28.4674
R659 VP.n25 VP.n24 28.4674
R660 VP.n11 VP.n10 28.4674
R661 VP.n20 VP.n19 24.5923
R662 VP.n20 VP.n1 24.5923
R663 VP.n6 VP.n5 24.5923
R664 VP.n8 VP.n7 17.507
R665 VP.n14 VP.n3 12.2964
R666 VP.n26 VP.n25 12.2964
R667 VP.n12 VP.n11 12.2964
R668 VP.n9 VP.n8 0.189894
R669 VP.n9 VP.n4 0.189894
R670 VP.n13 VP.n4 0.189894
R671 VP.n16 VP.n15 0.189894
R672 VP.n17 VP.n16 0.189894
R673 VP.n17 VP.n2 0.189894
R674 VP.n21 VP.n2 0.189894
R675 VP.n22 VP.n21 0.189894
R676 VP.n23 VP.n22 0.189894
R677 VP.n23 VP.n0 0.189894
R678 VP.n27 VP.n0 0.189894
R679 VP VP.n27 0.0516364
R680 VTAIL.n7 VTAIL.t1 114.924
R681 VTAIL.n11 VTAIL.t0 114.924
R682 VTAIL.n2 VTAIL.t9 114.924
R683 VTAIL.n10 VTAIL.t6 114.924
R684 VTAIL.n9 VTAIL.n8 105.945
R685 VTAIL.n6 VTAIL.n5 105.945
R686 VTAIL.n1 VTAIL.n0 105.945
R687 VTAIL.n4 VTAIL.n3 105.945
R688 VTAIL.n6 VTAIL.n4 18.5048
R689 VTAIL.n11 VTAIL.n10 16.9962
R690 VTAIL.n0 VTAIL.t2 8.97978
R691 VTAIL.n0 VTAIL.t3 8.97978
R692 VTAIL.n3 VTAIL.t10 8.97978
R693 VTAIL.n3 VTAIL.t7 8.97978
R694 VTAIL.n8 VTAIL.t8 8.97978
R695 VTAIL.n8 VTAIL.t5 8.97978
R696 VTAIL.n5 VTAIL.t11 8.97978
R697 VTAIL.n5 VTAIL.t4 8.97978
R698 VTAIL.n7 VTAIL.n6 1.50912
R699 VTAIL.n10 VTAIL.n9 1.50912
R700 VTAIL.n4 VTAIL.n2 1.50912
R701 VTAIL.n9 VTAIL.n7 1.22464
R702 VTAIL.n2 VTAIL.n1 1.22464
R703 VTAIL VTAIL.n11 1.07378
R704 VTAIL VTAIL.n1 0.435845
R705 VDD1 VDD1.t1 132.792
R706 VDD1.n1 VDD1.t5 132.679
R707 VDD1.n1 VDD1.n0 122.945
R708 VDD1.n3 VDD1.n2 122.624
R709 VDD1.n3 VDD1.n1 33.0763
R710 VDD1.n2 VDD1.t2 8.97978
R711 VDD1.n2 VDD1.t3 8.97978
R712 VDD1.n0 VDD1.t4 8.97978
R713 VDD1.n0 VDD1.t0 8.97978
R714 VDD1 VDD1.n3 0.319466
R715 VN.n9 VN.n8 173.596
R716 VN.n19 VN.n18 173.596
R717 VN.n17 VN.n10 161.3
R718 VN.n16 VN.n15 161.3
R719 VN.n14 VN.n11 161.3
R720 VN.n7 VN.n0 161.3
R721 VN.n6 VN.n5 161.3
R722 VN.n4 VN.n1 161.3
R723 VN.n3 VN.t5 96.9427
R724 VN.n13 VN.t3 96.9427
R725 VN.n2 VN.t4 61.4385
R726 VN.n8 VN.t2 61.4385
R727 VN.n12 VN.t0 61.4385
R728 VN.n18 VN.t1 61.4385
R729 VN.n6 VN.n1 52.6866
R730 VN.n16 VN.n11 52.6866
R731 VN.n3 VN.n2 41.915
R732 VN.n13 VN.n12 41.915
R733 VN VN.n19 38.0213
R734 VN.n7 VN.n6 28.4674
R735 VN.n17 VN.n16 28.4674
R736 VN.n2 VN.n1 24.5923
R737 VN.n12 VN.n11 24.5923
R738 VN.n14 VN.n13 17.507
R739 VN.n4 VN.n3 17.507
R740 VN.n8 VN.n7 12.2964
R741 VN.n18 VN.n17 12.2964
R742 VN.n19 VN.n10 0.189894
R743 VN.n15 VN.n10 0.189894
R744 VN.n15 VN.n14 0.189894
R745 VN.n5 VN.n4 0.189894
R746 VN.n5 VN.n0 0.189894
R747 VN.n9 VN.n0 0.189894
R748 VN VN.n9 0.0516364
R749 VDD2.n1 VDD2.t0 132.679
R750 VDD2.n2 VDD2.t4 131.602
R751 VDD2.n1 VDD2.n0 122.945
R752 VDD2 VDD2.n3 122.942
R753 VDD2.n2 VDD2.n1 31.739
R754 VDD2.n3 VDD2.t5 8.97978
R755 VDD2.n3 VDD2.t2 8.97978
R756 VDD2.n0 VDD2.t1 8.97978
R757 VDD2.n0 VDD2.t3 8.97978
R758 VDD2 VDD2.n2 1.19016
C0 VP VN 4.22998f
C1 VDD2 VN 1.99549f
C2 VTAIL B 1.43564f
C3 VDD2 VP 0.362796f
C4 VTAIL w_n2370_n1692# 1.64594f
C5 VDD1 VN 0.154001f
C6 w_n2370_n1692# B 5.70315f
C7 VDD1 VP 2.20218f
C8 VDD1 VDD2 0.975325f
C9 VTAIL VN 2.33555f
C10 VTAIL VP 2.34975f
C11 VTAIL VDD2 4.17866f
C12 VN B 0.825169f
C13 VN w_n2370_n1692# 4.0344f
C14 VP B 1.32504f
C15 VDD2 B 1.181f
C16 VTAIL VDD1 4.13439f
C17 VP w_n2370_n1692# 4.33612f
C18 VDD2 w_n2370_n1692# 1.44406f
C19 VDD1 B 1.13495f
C20 VDD1 w_n2370_n1692# 1.39743f
C21 VDD2 VSUBS 0.869712f
C22 VDD1 VSUBS 1.382645f
C23 VTAIL VSUBS 0.448269f
C24 VN VSUBS 4.09279f
C25 VP VSUBS 1.560276f
C26 B VSUBS 2.62106f
C27 w_n2370_n1692# VSUBS 50.5948f
C28 VDD2.t0 VSUBS 0.344897f
C29 VDD2.t1 VSUBS 0.043554f
C30 VDD2.t3 VSUBS 0.043554f
C31 VDD2.n0 VSUBS 0.246464f
C32 VDD2.n1 VSUBS 1.30522f
C33 VDD2.t4 VSUBS 0.342557f
C34 VDD2.n2 VSUBS 1.16368f
C35 VDD2.t5 VSUBS 0.043554f
C36 VDD2.t2 VSUBS 0.043554f
C37 VDD2.n3 VSUBS 0.246454f
C38 VN.n0 VSUBS 0.046118f
C39 VN.t2 VSUBS 0.603186f
C40 VN.n1 VSUBS 0.081919f
C41 VN.t5 VSUBS 0.762735f
C42 VN.t4 VSUBS 0.603186f
C43 VN.n2 VSUBS 0.368649f
C44 VN.n3 VSUBS 0.338775f
C45 VN.n4 VSUBS 0.290686f
C46 VN.n5 VSUBS 0.046118f
C47 VN.n6 VSUBS 0.047332f
C48 VN.n7 VSUBS 0.069239f
C49 VN.n8 VSUBS 0.356474f
C50 VN.n9 VSUBS 0.042814f
C51 VN.n10 VSUBS 0.046118f
C52 VN.t1 VSUBS 0.603186f
C53 VN.n11 VSUBS 0.081919f
C54 VN.t3 VSUBS 0.762735f
C55 VN.t0 VSUBS 0.603186f
C56 VN.n12 VSUBS 0.368649f
C57 VN.n13 VSUBS 0.338775f
C58 VN.n14 VSUBS 0.290686f
C59 VN.n15 VSUBS 0.046118f
C60 VN.n16 VSUBS 0.047332f
C61 VN.n17 VSUBS 0.069239f
C62 VN.n18 VSUBS 0.356474f
C63 VN.n19 VSUBS 1.61158f
C64 VDD1.t1 VSUBS 0.510944f
C65 VDD1.t5 VSUBS 0.51051f
C66 VDD1.t4 VSUBS 0.064468f
C67 VDD1.t0 VSUBS 0.064468f
C68 VDD1.n0 VSUBS 0.364812f
C69 VDD1.n1 VSUBS 2.0115f
C70 VDD1.t2 VSUBS 0.064468f
C71 VDD1.t3 VSUBS 0.064468f
C72 VDD1.n2 VSUBS 0.363632f
C73 VDD1.n3 VSUBS 1.74007f
C74 VTAIL.t2 VSUBS 0.080271f
C75 VTAIL.t3 VSUBS 0.080271f
C76 VTAIL.n0 VSUBS 0.393405f
C77 VTAIL.n1 VSUBS 0.553692f
C78 VTAIL.t9 VSUBS 0.570754f
C79 VTAIL.n2 VSUBS 0.692306f
C80 VTAIL.t10 VSUBS 0.080271f
C81 VTAIL.t7 VSUBS 0.080271f
C82 VTAIL.n3 VSUBS 0.393405f
C83 VTAIL.n4 VSUBS 1.4762f
C84 VTAIL.t11 VSUBS 0.080271f
C85 VTAIL.t4 VSUBS 0.080271f
C86 VTAIL.n5 VSUBS 0.393407f
C87 VTAIL.n6 VSUBS 1.47619f
C88 VTAIL.t1 VSUBS 0.570757f
C89 VTAIL.n7 VSUBS 0.692304f
C90 VTAIL.t8 VSUBS 0.080271f
C91 VTAIL.t5 VSUBS 0.080271f
C92 VTAIL.n8 VSUBS 0.393407f
C93 VTAIL.n9 VSUBS 0.650733f
C94 VTAIL.t6 VSUBS 0.570754f
C95 VTAIL.n10 VSUBS 1.38136f
C96 VTAIL.t0 VSUBS 0.570754f
C97 VTAIL.n11 VSUBS 1.342f
C98 VP.n0 VSUBS 0.057453f
C99 VP.t5 VSUBS 0.751441f
C100 VP.n1 VSUBS 0.102053f
C101 VP.n2 VSUBS 0.057453f
C102 VP.t1 VSUBS 0.751441f
C103 VP.n3 VSUBS 0.086257f
C104 VP.n4 VSUBS 0.057453f
C105 VP.t2 VSUBS 0.751441f
C106 VP.n5 VSUBS 0.102053f
C107 VP.t4 VSUBS 0.950206f
C108 VP.t3 VSUBS 0.751441f
C109 VP.n6 VSUBS 0.459259f
C110 VP.n7 VSUBS 0.422041f
C111 VP.n8 VSUBS 0.362133f
C112 VP.n9 VSUBS 0.057453f
C113 VP.n10 VSUBS 0.058965f
C114 VP.n11 VSUBS 0.086257f
C115 VP.n12 VSUBS 0.444091f
C116 VP.n13 VSUBS 1.96969f
C117 VP.t0 VSUBS 0.751441f
C118 VP.n14 VSUBS 0.444091f
C119 VP.n15 VSUBS 2.02472f
C120 VP.n16 VSUBS 0.057453f
C121 VP.n17 VSUBS 0.057453f
C122 VP.n18 VSUBS 0.058965f
C123 VP.n19 VSUBS 0.102053f
C124 VP.n20 VSUBS 0.382425f
C125 VP.n21 VSUBS 0.057453f
C126 VP.n22 VSUBS 0.057453f
C127 VP.n23 VSUBS 0.057453f
C128 VP.n24 VSUBS 0.058965f
C129 VP.n25 VSUBS 0.086257f
C130 VP.n26 VSUBS 0.444091f
C131 VP.n27 VSUBS 0.053337f
C132 B.n0 VSUBS 0.006546f
C133 B.n1 VSUBS 0.006546f
C134 B.n2 VSUBS 0.009681f
C135 B.n3 VSUBS 0.007419f
C136 B.n4 VSUBS 0.007419f
C137 B.n5 VSUBS 0.007419f
C138 B.n6 VSUBS 0.007419f
C139 B.n7 VSUBS 0.007419f
C140 B.n8 VSUBS 0.007419f
C141 B.n9 VSUBS 0.007419f
C142 B.n10 VSUBS 0.007419f
C143 B.n11 VSUBS 0.007419f
C144 B.n12 VSUBS 0.007419f
C145 B.n13 VSUBS 0.007419f
C146 B.n14 VSUBS 0.007419f
C147 B.n15 VSUBS 0.007419f
C148 B.n16 VSUBS 0.017881f
C149 B.n17 VSUBS 0.007419f
C150 B.n18 VSUBS 0.007419f
C151 B.n19 VSUBS 0.007419f
C152 B.n20 VSUBS 0.007419f
C153 B.n21 VSUBS 0.007419f
C154 B.n22 VSUBS 0.007419f
C155 B.n23 VSUBS 0.007419f
C156 B.n24 VSUBS 0.006982f
C157 B.n25 VSUBS 0.007419f
C158 B.t10 VSUBS 0.097672f
C159 B.t11 VSUBS 0.109244f
C160 B.t9 VSUBS 0.256525f
C161 B.n26 VSUBS 0.082632f
C162 B.n27 VSUBS 0.066588f
C163 B.n28 VSUBS 0.017188f
C164 B.n29 VSUBS 0.007419f
C165 B.n30 VSUBS 0.007419f
C166 B.n31 VSUBS 0.007419f
C167 B.n32 VSUBS 0.007419f
C168 B.t7 VSUBS 0.097672f
C169 B.t8 VSUBS 0.109244f
C170 B.t6 VSUBS 0.256525f
C171 B.n33 VSUBS 0.082632f
C172 B.n34 VSUBS 0.066588f
C173 B.n35 VSUBS 0.007419f
C174 B.n36 VSUBS 0.007419f
C175 B.n37 VSUBS 0.007419f
C176 B.n38 VSUBS 0.007419f
C177 B.n39 VSUBS 0.007419f
C178 B.n40 VSUBS 0.007419f
C179 B.n41 VSUBS 0.007419f
C180 B.n42 VSUBS 0.007419f
C181 B.n43 VSUBS 0.016375f
C182 B.n44 VSUBS 0.007419f
C183 B.n45 VSUBS 0.007419f
C184 B.n46 VSUBS 0.007419f
C185 B.n47 VSUBS 0.007419f
C186 B.n48 VSUBS 0.007419f
C187 B.n49 VSUBS 0.007419f
C188 B.n50 VSUBS 0.007419f
C189 B.n51 VSUBS 0.007419f
C190 B.n52 VSUBS 0.007419f
C191 B.n53 VSUBS 0.007419f
C192 B.n54 VSUBS 0.007419f
C193 B.n55 VSUBS 0.007419f
C194 B.n56 VSUBS 0.007419f
C195 B.n57 VSUBS 0.007419f
C196 B.n58 VSUBS 0.007419f
C197 B.n59 VSUBS 0.007419f
C198 B.n60 VSUBS 0.007419f
C199 B.n61 VSUBS 0.007419f
C200 B.n62 VSUBS 0.007419f
C201 B.n63 VSUBS 0.007419f
C202 B.n64 VSUBS 0.007419f
C203 B.n65 VSUBS 0.007419f
C204 B.n66 VSUBS 0.007419f
C205 B.n67 VSUBS 0.007419f
C206 B.n68 VSUBS 0.007419f
C207 B.n69 VSUBS 0.007419f
C208 B.n70 VSUBS 0.007419f
C209 B.n71 VSUBS 0.007419f
C210 B.n72 VSUBS 0.017881f
C211 B.n73 VSUBS 0.007419f
C212 B.n74 VSUBS 0.007419f
C213 B.n75 VSUBS 0.007419f
C214 B.n76 VSUBS 0.007419f
C215 B.n77 VSUBS 0.007419f
C216 B.n78 VSUBS 0.007419f
C217 B.n79 VSUBS 0.007419f
C218 B.n80 VSUBS 0.007419f
C219 B.t5 VSUBS 0.097672f
C220 B.t4 VSUBS 0.109244f
C221 B.t3 VSUBS 0.256525f
C222 B.n81 VSUBS 0.082632f
C223 B.n82 VSUBS 0.066588f
C224 B.n83 VSUBS 0.007419f
C225 B.n84 VSUBS 0.007419f
C226 B.n85 VSUBS 0.007419f
C227 B.n86 VSUBS 0.007419f
C228 B.n87 VSUBS 0.004146f
C229 B.n88 VSUBS 0.007419f
C230 B.n89 VSUBS 0.007419f
C231 B.n90 VSUBS 0.007419f
C232 B.n91 VSUBS 0.007419f
C233 B.n92 VSUBS 0.007419f
C234 B.n93 VSUBS 0.007419f
C235 B.n94 VSUBS 0.007419f
C236 B.n95 VSUBS 0.007419f
C237 B.n96 VSUBS 0.016375f
C238 B.n97 VSUBS 0.007419f
C239 B.n98 VSUBS 0.007419f
C240 B.n99 VSUBS 0.007419f
C241 B.n100 VSUBS 0.007419f
C242 B.n101 VSUBS 0.007419f
C243 B.n102 VSUBS 0.007419f
C244 B.n103 VSUBS 0.007419f
C245 B.n104 VSUBS 0.007419f
C246 B.n105 VSUBS 0.007419f
C247 B.n106 VSUBS 0.007419f
C248 B.n107 VSUBS 0.007419f
C249 B.n108 VSUBS 0.007419f
C250 B.n109 VSUBS 0.007419f
C251 B.n110 VSUBS 0.007419f
C252 B.n111 VSUBS 0.007419f
C253 B.n112 VSUBS 0.007419f
C254 B.n113 VSUBS 0.007419f
C255 B.n114 VSUBS 0.007419f
C256 B.n115 VSUBS 0.007419f
C257 B.n116 VSUBS 0.007419f
C258 B.n117 VSUBS 0.007419f
C259 B.n118 VSUBS 0.007419f
C260 B.n119 VSUBS 0.007419f
C261 B.n120 VSUBS 0.007419f
C262 B.n121 VSUBS 0.007419f
C263 B.n122 VSUBS 0.007419f
C264 B.n123 VSUBS 0.007419f
C265 B.n124 VSUBS 0.007419f
C266 B.n125 VSUBS 0.007419f
C267 B.n126 VSUBS 0.007419f
C268 B.n127 VSUBS 0.007419f
C269 B.n128 VSUBS 0.007419f
C270 B.n129 VSUBS 0.007419f
C271 B.n130 VSUBS 0.007419f
C272 B.n131 VSUBS 0.007419f
C273 B.n132 VSUBS 0.007419f
C274 B.n133 VSUBS 0.007419f
C275 B.n134 VSUBS 0.007419f
C276 B.n135 VSUBS 0.007419f
C277 B.n136 VSUBS 0.007419f
C278 B.n137 VSUBS 0.007419f
C279 B.n138 VSUBS 0.007419f
C280 B.n139 VSUBS 0.007419f
C281 B.n140 VSUBS 0.007419f
C282 B.n141 VSUBS 0.007419f
C283 B.n142 VSUBS 0.007419f
C284 B.n143 VSUBS 0.007419f
C285 B.n144 VSUBS 0.007419f
C286 B.n145 VSUBS 0.007419f
C287 B.n146 VSUBS 0.007419f
C288 B.n147 VSUBS 0.007419f
C289 B.n148 VSUBS 0.007419f
C290 B.n149 VSUBS 0.016375f
C291 B.n150 VSUBS 0.017881f
C292 B.n151 VSUBS 0.017881f
C293 B.n152 VSUBS 0.007419f
C294 B.n153 VSUBS 0.007419f
C295 B.n154 VSUBS 0.007419f
C296 B.n155 VSUBS 0.007419f
C297 B.n156 VSUBS 0.007419f
C298 B.n157 VSUBS 0.007419f
C299 B.n158 VSUBS 0.007419f
C300 B.n159 VSUBS 0.007419f
C301 B.n160 VSUBS 0.007419f
C302 B.n161 VSUBS 0.007419f
C303 B.n162 VSUBS 0.007419f
C304 B.n163 VSUBS 0.007419f
C305 B.n164 VSUBS 0.007419f
C306 B.n165 VSUBS 0.007419f
C307 B.n166 VSUBS 0.007419f
C308 B.n167 VSUBS 0.007419f
C309 B.n168 VSUBS 0.007419f
C310 B.n169 VSUBS 0.007419f
C311 B.n170 VSUBS 0.007419f
C312 B.n171 VSUBS 0.007419f
C313 B.n172 VSUBS 0.007419f
C314 B.n173 VSUBS 0.007419f
C315 B.t2 VSUBS 0.097672f
C316 B.t1 VSUBS 0.109244f
C317 B.t0 VSUBS 0.256525f
C318 B.n174 VSUBS 0.082632f
C319 B.n175 VSUBS 0.066588f
C320 B.n176 VSUBS 0.017188f
C321 B.n177 VSUBS 0.006982f
C322 B.n178 VSUBS 0.007419f
C323 B.n179 VSUBS 0.007419f
C324 B.n180 VSUBS 0.007419f
C325 B.n181 VSUBS 0.007419f
C326 B.n182 VSUBS 0.007419f
C327 B.n183 VSUBS 0.007419f
C328 B.n184 VSUBS 0.007419f
C329 B.n185 VSUBS 0.007419f
C330 B.n186 VSUBS 0.007419f
C331 B.n187 VSUBS 0.007419f
C332 B.n188 VSUBS 0.007419f
C333 B.n189 VSUBS 0.007419f
C334 B.n190 VSUBS 0.007419f
C335 B.n191 VSUBS 0.007419f
C336 B.n192 VSUBS 0.007419f
C337 B.n193 VSUBS 0.004146f
C338 B.n194 VSUBS 0.017188f
C339 B.n195 VSUBS 0.006982f
C340 B.n196 VSUBS 0.007419f
C341 B.n197 VSUBS 0.007419f
C342 B.n198 VSUBS 0.007419f
C343 B.n199 VSUBS 0.007419f
C344 B.n200 VSUBS 0.007419f
C345 B.n201 VSUBS 0.007419f
C346 B.n202 VSUBS 0.007419f
C347 B.n203 VSUBS 0.007419f
C348 B.n204 VSUBS 0.007419f
C349 B.n205 VSUBS 0.007419f
C350 B.n206 VSUBS 0.007419f
C351 B.n207 VSUBS 0.007419f
C352 B.n208 VSUBS 0.007419f
C353 B.n209 VSUBS 0.007419f
C354 B.n210 VSUBS 0.007419f
C355 B.n211 VSUBS 0.007419f
C356 B.n212 VSUBS 0.007419f
C357 B.n213 VSUBS 0.007419f
C358 B.n214 VSUBS 0.007419f
C359 B.n215 VSUBS 0.007419f
C360 B.n216 VSUBS 0.007419f
C361 B.n217 VSUBS 0.007419f
C362 B.n218 VSUBS 0.007419f
C363 B.n219 VSUBS 0.016986f
C364 B.n220 VSUBS 0.01727f
C365 B.n221 VSUBS 0.016375f
C366 B.n222 VSUBS 0.007419f
C367 B.n223 VSUBS 0.007419f
C368 B.n224 VSUBS 0.007419f
C369 B.n225 VSUBS 0.007419f
C370 B.n226 VSUBS 0.007419f
C371 B.n227 VSUBS 0.007419f
C372 B.n228 VSUBS 0.007419f
C373 B.n229 VSUBS 0.007419f
C374 B.n230 VSUBS 0.007419f
C375 B.n231 VSUBS 0.007419f
C376 B.n232 VSUBS 0.007419f
C377 B.n233 VSUBS 0.007419f
C378 B.n234 VSUBS 0.007419f
C379 B.n235 VSUBS 0.007419f
C380 B.n236 VSUBS 0.007419f
C381 B.n237 VSUBS 0.007419f
C382 B.n238 VSUBS 0.007419f
C383 B.n239 VSUBS 0.007419f
C384 B.n240 VSUBS 0.007419f
C385 B.n241 VSUBS 0.007419f
C386 B.n242 VSUBS 0.007419f
C387 B.n243 VSUBS 0.007419f
C388 B.n244 VSUBS 0.007419f
C389 B.n245 VSUBS 0.007419f
C390 B.n246 VSUBS 0.007419f
C391 B.n247 VSUBS 0.007419f
C392 B.n248 VSUBS 0.007419f
C393 B.n249 VSUBS 0.007419f
C394 B.n250 VSUBS 0.007419f
C395 B.n251 VSUBS 0.007419f
C396 B.n252 VSUBS 0.007419f
C397 B.n253 VSUBS 0.007419f
C398 B.n254 VSUBS 0.007419f
C399 B.n255 VSUBS 0.007419f
C400 B.n256 VSUBS 0.007419f
C401 B.n257 VSUBS 0.007419f
C402 B.n258 VSUBS 0.007419f
C403 B.n259 VSUBS 0.007419f
C404 B.n260 VSUBS 0.007419f
C405 B.n261 VSUBS 0.007419f
C406 B.n262 VSUBS 0.007419f
C407 B.n263 VSUBS 0.007419f
C408 B.n264 VSUBS 0.007419f
C409 B.n265 VSUBS 0.007419f
C410 B.n266 VSUBS 0.007419f
C411 B.n267 VSUBS 0.007419f
C412 B.n268 VSUBS 0.007419f
C413 B.n269 VSUBS 0.007419f
C414 B.n270 VSUBS 0.007419f
C415 B.n271 VSUBS 0.007419f
C416 B.n272 VSUBS 0.007419f
C417 B.n273 VSUBS 0.007419f
C418 B.n274 VSUBS 0.007419f
C419 B.n275 VSUBS 0.007419f
C420 B.n276 VSUBS 0.007419f
C421 B.n277 VSUBS 0.007419f
C422 B.n278 VSUBS 0.007419f
C423 B.n279 VSUBS 0.007419f
C424 B.n280 VSUBS 0.007419f
C425 B.n281 VSUBS 0.007419f
C426 B.n282 VSUBS 0.007419f
C427 B.n283 VSUBS 0.007419f
C428 B.n284 VSUBS 0.007419f
C429 B.n285 VSUBS 0.007419f
C430 B.n286 VSUBS 0.007419f
C431 B.n287 VSUBS 0.007419f
C432 B.n288 VSUBS 0.007419f
C433 B.n289 VSUBS 0.007419f
C434 B.n290 VSUBS 0.007419f
C435 B.n291 VSUBS 0.007419f
C436 B.n292 VSUBS 0.007419f
C437 B.n293 VSUBS 0.007419f
C438 B.n294 VSUBS 0.007419f
C439 B.n295 VSUBS 0.007419f
C440 B.n296 VSUBS 0.007419f
C441 B.n297 VSUBS 0.007419f
C442 B.n298 VSUBS 0.007419f
C443 B.n299 VSUBS 0.007419f
C444 B.n300 VSUBS 0.007419f
C445 B.n301 VSUBS 0.007419f
C446 B.n302 VSUBS 0.007419f
C447 B.n303 VSUBS 0.007419f
C448 B.n304 VSUBS 0.007419f
C449 B.n305 VSUBS 0.007419f
C450 B.n306 VSUBS 0.016375f
C451 B.n307 VSUBS 0.017881f
C452 B.n308 VSUBS 0.017881f
C453 B.n309 VSUBS 0.007419f
C454 B.n310 VSUBS 0.007419f
C455 B.n311 VSUBS 0.007419f
C456 B.n312 VSUBS 0.007419f
C457 B.n313 VSUBS 0.007419f
C458 B.n314 VSUBS 0.007419f
C459 B.n315 VSUBS 0.007419f
C460 B.n316 VSUBS 0.007419f
C461 B.n317 VSUBS 0.007419f
C462 B.n318 VSUBS 0.007419f
C463 B.n319 VSUBS 0.007419f
C464 B.n320 VSUBS 0.007419f
C465 B.n321 VSUBS 0.007419f
C466 B.n322 VSUBS 0.007419f
C467 B.n323 VSUBS 0.007419f
C468 B.n324 VSUBS 0.007419f
C469 B.n325 VSUBS 0.007419f
C470 B.n326 VSUBS 0.007419f
C471 B.n327 VSUBS 0.007419f
C472 B.n328 VSUBS 0.007419f
C473 B.n329 VSUBS 0.007419f
C474 B.n330 VSUBS 0.007419f
C475 B.n331 VSUBS 0.007419f
C476 B.n332 VSUBS 0.006982f
C477 B.n333 VSUBS 0.017188f
C478 B.n334 VSUBS 0.004146f
C479 B.n335 VSUBS 0.007419f
C480 B.n336 VSUBS 0.007419f
C481 B.n337 VSUBS 0.007419f
C482 B.n338 VSUBS 0.007419f
C483 B.n339 VSUBS 0.007419f
C484 B.n340 VSUBS 0.007419f
C485 B.n341 VSUBS 0.007419f
C486 B.n342 VSUBS 0.007419f
C487 B.n343 VSUBS 0.007419f
C488 B.n344 VSUBS 0.007419f
C489 B.n345 VSUBS 0.007419f
C490 B.n346 VSUBS 0.007419f
C491 B.n347 VSUBS 0.004146f
C492 B.n348 VSUBS 0.007419f
C493 B.n349 VSUBS 0.007419f
C494 B.n350 VSUBS 0.007419f
C495 B.n351 VSUBS 0.007419f
C496 B.n352 VSUBS 0.007419f
C497 B.n353 VSUBS 0.007419f
C498 B.n354 VSUBS 0.007419f
C499 B.n355 VSUBS 0.007419f
C500 B.n356 VSUBS 0.007419f
C501 B.n357 VSUBS 0.007419f
C502 B.n358 VSUBS 0.007419f
C503 B.n359 VSUBS 0.007419f
C504 B.n360 VSUBS 0.007419f
C505 B.n361 VSUBS 0.007419f
C506 B.n362 VSUBS 0.007419f
C507 B.n363 VSUBS 0.007419f
C508 B.n364 VSUBS 0.007419f
C509 B.n365 VSUBS 0.007419f
C510 B.n366 VSUBS 0.007419f
C511 B.n367 VSUBS 0.007419f
C512 B.n368 VSUBS 0.007419f
C513 B.n369 VSUBS 0.007419f
C514 B.n370 VSUBS 0.007419f
C515 B.n371 VSUBS 0.007419f
C516 B.n372 VSUBS 0.007419f
C517 B.n373 VSUBS 0.017881f
C518 B.n374 VSUBS 0.016375f
C519 B.n375 VSUBS 0.016375f
C520 B.n376 VSUBS 0.007419f
C521 B.n377 VSUBS 0.007419f
C522 B.n378 VSUBS 0.007419f
C523 B.n379 VSUBS 0.007419f
C524 B.n380 VSUBS 0.007419f
C525 B.n381 VSUBS 0.007419f
C526 B.n382 VSUBS 0.007419f
C527 B.n383 VSUBS 0.007419f
C528 B.n384 VSUBS 0.007419f
C529 B.n385 VSUBS 0.007419f
C530 B.n386 VSUBS 0.007419f
C531 B.n387 VSUBS 0.007419f
C532 B.n388 VSUBS 0.007419f
C533 B.n389 VSUBS 0.007419f
C534 B.n390 VSUBS 0.007419f
C535 B.n391 VSUBS 0.007419f
C536 B.n392 VSUBS 0.007419f
C537 B.n393 VSUBS 0.007419f
C538 B.n394 VSUBS 0.007419f
C539 B.n395 VSUBS 0.007419f
C540 B.n396 VSUBS 0.007419f
C541 B.n397 VSUBS 0.007419f
C542 B.n398 VSUBS 0.007419f
C543 B.n399 VSUBS 0.007419f
C544 B.n400 VSUBS 0.007419f
C545 B.n401 VSUBS 0.007419f
C546 B.n402 VSUBS 0.007419f
C547 B.n403 VSUBS 0.007419f
C548 B.n404 VSUBS 0.007419f
C549 B.n405 VSUBS 0.007419f
C550 B.n406 VSUBS 0.007419f
C551 B.n407 VSUBS 0.007419f
C552 B.n408 VSUBS 0.007419f
C553 B.n409 VSUBS 0.007419f
C554 B.n410 VSUBS 0.007419f
C555 B.n411 VSUBS 0.007419f
C556 B.n412 VSUBS 0.007419f
C557 B.n413 VSUBS 0.007419f
C558 B.n414 VSUBS 0.007419f
C559 B.n415 VSUBS 0.009681f
C560 B.n416 VSUBS 0.010313f
C561 B.n417 VSUBS 0.020507f
.ends

