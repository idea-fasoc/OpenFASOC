* NGSPICE file created from diff_pair_sample_1442.ext - technology: sky130A

.subckt diff_pair_sample_1442 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=0 ps=0 w=18.41 l=0.64
X1 VDD1.t7 VP.t0 VTAIL.t11 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=7.1799 ps=37.6 w=18.41 l=0.64
X2 VDD2.t7 VN.t0 VTAIL.t2 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X3 B.t8 B.t6 B.t7 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=0 ps=0 w=18.41 l=0.64
X4 VDD1.t6 VP.t1 VTAIL.t8 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X5 VTAIL.t3 VN.t1 VDD2.t6 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=3.03765 ps=18.74 w=18.41 l=0.64
X6 VTAIL.t12 VP.t2 VDD1.t5 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=3.03765 ps=18.74 w=18.41 l=0.64
X7 VDD2.t5 VN.t2 VTAIL.t4 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=7.1799 ps=37.6 w=18.41 l=0.64
X8 VDD2.t4 VN.t3 VTAIL.t1 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=7.1799 ps=37.6 w=18.41 l=0.64
X9 B.t5 B.t3 B.t4 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=0 ps=0 w=18.41 l=0.64
X10 VTAIL.t0 VN.t4 VDD2.t3 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=3.03765 ps=18.74 w=18.41 l=0.64
X11 VDD1.t4 VP.t3 VTAIL.t13 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X12 VTAIL.t9 VP.t4 VDD1.t3 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X13 B.t2 B.t0 B.t1 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=0 ps=0 w=18.41 l=0.64
X14 VTAIL.t7 VN.t5 VDD2.t2 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X15 VTAIL.t6 VN.t6 VDD2.t1 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X16 VTAIL.t15 VP.t5 VDD1.t2 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
X17 VTAIL.t14 VP.t6 VDD1.t1 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=7.1799 pd=37.6 as=3.03765 ps=18.74 w=18.41 l=0.64
X18 VDD1.t0 VP.t7 VTAIL.t10 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=7.1799 ps=37.6 w=18.41 l=0.64
X19 VDD2.t0 VN.t7 VTAIL.t5 w_n1940_n4650# sky130_fd_pr__pfet_01v8 ad=3.03765 pd=18.74 as=3.03765 ps=18.74 w=18.41 l=0.64
R0 B.n142 B.t0 897.024
R1 B.n320 B.t6 897.024
R2 B.n50 B.t9 897.024
R3 B.n44 B.t3 897.024
R4 B.n415 B.n106 585
R5 B.n414 B.n413 585
R6 B.n412 B.n107 585
R7 B.n411 B.n410 585
R8 B.n409 B.n108 585
R9 B.n408 B.n407 585
R10 B.n406 B.n109 585
R11 B.n405 B.n404 585
R12 B.n403 B.n110 585
R13 B.n402 B.n401 585
R14 B.n400 B.n111 585
R15 B.n399 B.n398 585
R16 B.n397 B.n112 585
R17 B.n396 B.n395 585
R18 B.n394 B.n113 585
R19 B.n393 B.n392 585
R20 B.n391 B.n114 585
R21 B.n390 B.n389 585
R22 B.n388 B.n115 585
R23 B.n387 B.n386 585
R24 B.n385 B.n116 585
R25 B.n384 B.n383 585
R26 B.n382 B.n117 585
R27 B.n381 B.n380 585
R28 B.n379 B.n118 585
R29 B.n378 B.n377 585
R30 B.n376 B.n119 585
R31 B.n375 B.n374 585
R32 B.n373 B.n120 585
R33 B.n372 B.n371 585
R34 B.n370 B.n121 585
R35 B.n369 B.n368 585
R36 B.n367 B.n122 585
R37 B.n366 B.n365 585
R38 B.n364 B.n123 585
R39 B.n363 B.n362 585
R40 B.n361 B.n124 585
R41 B.n360 B.n359 585
R42 B.n358 B.n125 585
R43 B.n357 B.n356 585
R44 B.n355 B.n126 585
R45 B.n354 B.n353 585
R46 B.n352 B.n127 585
R47 B.n351 B.n350 585
R48 B.n349 B.n128 585
R49 B.n348 B.n347 585
R50 B.n346 B.n129 585
R51 B.n345 B.n344 585
R52 B.n343 B.n130 585
R53 B.n342 B.n341 585
R54 B.n340 B.n131 585
R55 B.n339 B.n338 585
R56 B.n337 B.n132 585
R57 B.n336 B.n335 585
R58 B.n334 B.n133 585
R59 B.n333 B.n332 585
R60 B.n331 B.n134 585
R61 B.n330 B.n329 585
R62 B.n328 B.n135 585
R63 B.n327 B.n326 585
R64 B.n325 B.n136 585
R65 B.n324 B.n323 585
R66 B.n319 B.n137 585
R67 B.n318 B.n317 585
R68 B.n316 B.n138 585
R69 B.n315 B.n314 585
R70 B.n313 B.n139 585
R71 B.n312 B.n311 585
R72 B.n310 B.n140 585
R73 B.n309 B.n308 585
R74 B.n306 B.n141 585
R75 B.n305 B.n304 585
R76 B.n303 B.n144 585
R77 B.n302 B.n301 585
R78 B.n300 B.n145 585
R79 B.n299 B.n298 585
R80 B.n297 B.n146 585
R81 B.n296 B.n295 585
R82 B.n294 B.n147 585
R83 B.n293 B.n292 585
R84 B.n291 B.n148 585
R85 B.n290 B.n289 585
R86 B.n288 B.n149 585
R87 B.n287 B.n286 585
R88 B.n285 B.n150 585
R89 B.n284 B.n283 585
R90 B.n282 B.n151 585
R91 B.n281 B.n280 585
R92 B.n279 B.n152 585
R93 B.n278 B.n277 585
R94 B.n276 B.n153 585
R95 B.n275 B.n274 585
R96 B.n273 B.n154 585
R97 B.n272 B.n271 585
R98 B.n270 B.n155 585
R99 B.n269 B.n268 585
R100 B.n267 B.n156 585
R101 B.n266 B.n265 585
R102 B.n264 B.n157 585
R103 B.n263 B.n262 585
R104 B.n261 B.n158 585
R105 B.n260 B.n259 585
R106 B.n258 B.n159 585
R107 B.n257 B.n256 585
R108 B.n255 B.n160 585
R109 B.n254 B.n253 585
R110 B.n252 B.n161 585
R111 B.n251 B.n250 585
R112 B.n249 B.n162 585
R113 B.n248 B.n247 585
R114 B.n246 B.n163 585
R115 B.n245 B.n244 585
R116 B.n243 B.n164 585
R117 B.n242 B.n241 585
R118 B.n240 B.n165 585
R119 B.n239 B.n238 585
R120 B.n237 B.n166 585
R121 B.n236 B.n235 585
R122 B.n234 B.n167 585
R123 B.n233 B.n232 585
R124 B.n231 B.n168 585
R125 B.n230 B.n229 585
R126 B.n228 B.n169 585
R127 B.n227 B.n226 585
R128 B.n225 B.n170 585
R129 B.n224 B.n223 585
R130 B.n222 B.n171 585
R131 B.n221 B.n220 585
R132 B.n219 B.n172 585
R133 B.n218 B.n217 585
R134 B.n216 B.n173 585
R135 B.n417 B.n416 585
R136 B.n418 B.n105 585
R137 B.n420 B.n419 585
R138 B.n421 B.n104 585
R139 B.n423 B.n422 585
R140 B.n424 B.n103 585
R141 B.n426 B.n425 585
R142 B.n427 B.n102 585
R143 B.n429 B.n428 585
R144 B.n430 B.n101 585
R145 B.n432 B.n431 585
R146 B.n433 B.n100 585
R147 B.n435 B.n434 585
R148 B.n436 B.n99 585
R149 B.n438 B.n437 585
R150 B.n439 B.n98 585
R151 B.n441 B.n440 585
R152 B.n442 B.n97 585
R153 B.n444 B.n443 585
R154 B.n445 B.n96 585
R155 B.n447 B.n446 585
R156 B.n448 B.n95 585
R157 B.n450 B.n449 585
R158 B.n451 B.n94 585
R159 B.n453 B.n452 585
R160 B.n454 B.n93 585
R161 B.n456 B.n455 585
R162 B.n457 B.n92 585
R163 B.n459 B.n458 585
R164 B.n460 B.n91 585
R165 B.n462 B.n461 585
R166 B.n463 B.n90 585
R167 B.n465 B.n464 585
R168 B.n466 B.n89 585
R169 B.n468 B.n467 585
R170 B.n469 B.n88 585
R171 B.n471 B.n470 585
R172 B.n472 B.n87 585
R173 B.n474 B.n473 585
R174 B.n475 B.n86 585
R175 B.n477 B.n476 585
R176 B.n478 B.n85 585
R177 B.n480 B.n479 585
R178 B.n481 B.n84 585
R179 B.n483 B.n482 585
R180 B.n484 B.n83 585
R181 B.n682 B.n13 585
R182 B.n681 B.n680 585
R183 B.n679 B.n14 585
R184 B.n678 B.n677 585
R185 B.n676 B.n15 585
R186 B.n675 B.n674 585
R187 B.n673 B.n16 585
R188 B.n672 B.n671 585
R189 B.n670 B.n17 585
R190 B.n669 B.n668 585
R191 B.n667 B.n18 585
R192 B.n666 B.n665 585
R193 B.n664 B.n19 585
R194 B.n663 B.n662 585
R195 B.n661 B.n20 585
R196 B.n660 B.n659 585
R197 B.n658 B.n21 585
R198 B.n657 B.n656 585
R199 B.n655 B.n22 585
R200 B.n654 B.n653 585
R201 B.n652 B.n23 585
R202 B.n651 B.n650 585
R203 B.n649 B.n24 585
R204 B.n648 B.n647 585
R205 B.n646 B.n25 585
R206 B.n645 B.n644 585
R207 B.n643 B.n26 585
R208 B.n642 B.n641 585
R209 B.n640 B.n27 585
R210 B.n639 B.n638 585
R211 B.n637 B.n28 585
R212 B.n636 B.n635 585
R213 B.n634 B.n29 585
R214 B.n633 B.n632 585
R215 B.n631 B.n30 585
R216 B.n630 B.n629 585
R217 B.n628 B.n31 585
R218 B.n627 B.n626 585
R219 B.n625 B.n32 585
R220 B.n624 B.n623 585
R221 B.n622 B.n33 585
R222 B.n621 B.n620 585
R223 B.n619 B.n34 585
R224 B.n618 B.n617 585
R225 B.n616 B.n35 585
R226 B.n615 B.n614 585
R227 B.n613 B.n36 585
R228 B.n612 B.n611 585
R229 B.n610 B.n37 585
R230 B.n609 B.n608 585
R231 B.n607 B.n38 585
R232 B.n606 B.n605 585
R233 B.n604 B.n39 585
R234 B.n603 B.n602 585
R235 B.n601 B.n40 585
R236 B.n600 B.n599 585
R237 B.n598 B.n41 585
R238 B.n597 B.n596 585
R239 B.n595 B.n42 585
R240 B.n594 B.n593 585
R241 B.n592 B.n43 585
R242 B.n590 B.n589 585
R243 B.n588 B.n46 585
R244 B.n587 B.n586 585
R245 B.n585 B.n47 585
R246 B.n584 B.n583 585
R247 B.n582 B.n48 585
R248 B.n581 B.n580 585
R249 B.n579 B.n49 585
R250 B.n578 B.n577 585
R251 B.n576 B.n575 585
R252 B.n574 B.n53 585
R253 B.n573 B.n572 585
R254 B.n571 B.n54 585
R255 B.n570 B.n569 585
R256 B.n568 B.n55 585
R257 B.n567 B.n566 585
R258 B.n565 B.n56 585
R259 B.n564 B.n563 585
R260 B.n562 B.n57 585
R261 B.n561 B.n560 585
R262 B.n559 B.n58 585
R263 B.n558 B.n557 585
R264 B.n556 B.n59 585
R265 B.n555 B.n554 585
R266 B.n553 B.n60 585
R267 B.n552 B.n551 585
R268 B.n550 B.n61 585
R269 B.n549 B.n548 585
R270 B.n547 B.n62 585
R271 B.n546 B.n545 585
R272 B.n544 B.n63 585
R273 B.n543 B.n542 585
R274 B.n541 B.n64 585
R275 B.n540 B.n539 585
R276 B.n538 B.n65 585
R277 B.n537 B.n536 585
R278 B.n535 B.n66 585
R279 B.n534 B.n533 585
R280 B.n532 B.n67 585
R281 B.n531 B.n530 585
R282 B.n529 B.n68 585
R283 B.n528 B.n527 585
R284 B.n526 B.n69 585
R285 B.n525 B.n524 585
R286 B.n523 B.n70 585
R287 B.n522 B.n521 585
R288 B.n520 B.n71 585
R289 B.n519 B.n518 585
R290 B.n517 B.n72 585
R291 B.n516 B.n515 585
R292 B.n514 B.n73 585
R293 B.n513 B.n512 585
R294 B.n511 B.n74 585
R295 B.n510 B.n509 585
R296 B.n508 B.n75 585
R297 B.n507 B.n506 585
R298 B.n505 B.n76 585
R299 B.n504 B.n503 585
R300 B.n502 B.n77 585
R301 B.n501 B.n500 585
R302 B.n499 B.n78 585
R303 B.n498 B.n497 585
R304 B.n496 B.n79 585
R305 B.n495 B.n494 585
R306 B.n493 B.n80 585
R307 B.n492 B.n491 585
R308 B.n490 B.n81 585
R309 B.n489 B.n488 585
R310 B.n487 B.n82 585
R311 B.n486 B.n485 585
R312 B.n684 B.n683 585
R313 B.n685 B.n12 585
R314 B.n687 B.n686 585
R315 B.n688 B.n11 585
R316 B.n690 B.n689 585
R317 B.n691 B.n10 585
R318 B.n693 B.n692 585
R319 B.n694 B.n9 585
R320 B.n696 B.n695 585
R321 B.n697 B.n8 585
R322 B.n699 B.n698 585
R323 B.n700 B.n7 585
R324 B.n702 B.n701 585
R325 B.n703 B.n6 585
R326 B.n705 B.n704 585
R327 B.n706 B.n5 585
R328 B.n708 B.n707 585
R329 B.n709 B.n4 585
R330 B.n711 B.n710 585
R331 B.n712 B.n3 585
R332 B.n714 B.n713 585
R333 B.n715 B.n0 585
R334 B.n2 B.n1 585
R335 B.n185 B.n184 585
R336 B.n186 B.n183 585
R337 B.n188 B.n187 585
R338 B.n189 B.n182 585
R339 B.n191 B.n190 585
R340 B.n192 B.n181 585
R341 B.n194 B.n193 585
R342 B.n195 B.n180 585
R343 B.n197 B.n196 585
R344 B.n198 B.n179 585
R345 B.n200 B.n199 585
R346 B.n201 B.n178 585
R347 B.n203 B.n202 585
R348 B.n204 B.n177 585
R349 B.n206 B.n205 585
R350 B.n207 B.n176 585
R351 B.n209 B.n208 585
R352 B.n210 B.n175 585
R353 B.n212 B.n211 585
R354 B.n213 B.n174 585
R355 B.n215 B.n214 585
R356 B.n214 B.n173 439.647
R357 B.n416 B.n415 439.647
R358 B.n486 B.n83 439.647
R359 B.n684 B.n13 439.647
R360 B.n717 B.n716 256.663
R361 B.n716 B.n715 235.042
R362 B.n716 B.n2 235.042
R363 B.n218 B.n173 163.367
R364 B.n219 B.n218 163.367
R365 B.n220 B.n219 163.367
R366 B.n220 B.n171 163.367
R367 B.n224 B.n171 163.367
R368 B.n225 B.n224 163.367
R369 B.n226 B.n225 163.367
R370 B.n226 B.n169 163.367
R371 B.n230 B.n169 163.367
R372 B.n231 B.n230 163.367
R373 B.n232 B.n231 163.367
R374 B.n232 B.n167 163.367
R375 B.n236 B.n167 163.367
R376 B.n237 B.n236 163.367
R377 B.n238 B.n237 163.367
R378 B.n238 B.n165 163.367
R379 B.n242 B.n165 163.367
R380 B.n243 B.n242 163.367
R381 B.n244 B.n243 163.367
R382 B.n244 B.n163 163.367
R383 B.n248 B.n163 163.367
R384 B.n249 B.n248 163.367
R385 B.n250 B.n249 163.367
R386 B.n250 B.n161 163.367
R387 B.n254 B.n161 163.367
R388 B.n255 B.n254 163.367
R389 B.n256 B.n255 163.367
R390 B.n256 B.n159 163.367
R391 B.n260 B.n159 163.367
R392 B.n261 B.n260 163.367
R393 B.n262 B.n261 163.367
R394 B.n262 B.n157 163.367
R395 B.n266 B.n157 163.367
R396 B.n267 B.n266 163.367
R397 B.n268 B.n267 163.367
R398 B.n268 B.n155 163.367
R399 B.n272 B.n155 163.367
R400 B.n273 B.n272 163.367
R401 B.n274 B.n273 163.367
R402 B.n274 B.n153 163.367
R403 B.n278 B.n153 163.367
R404 B.n279 B.n278 163.367
R405 B.n280 B.n279 163.367
R406 B.n280 B.n151 163.367
R407 B.n284 B.n151 163.367
R408 B.n285 B.n284 163.367
R409 B.n286 B.n285 163.367
R410 B.n286 B.n149 163.367
R411 B.n290 B.n149 163.367
R412 B.n291 B.n290 163.367
R413 B.n292 B.n291 163.367
R414 B.n292 B.n147 163.367
R415 B.n296 B.n147 163.367
R416 B.n297 B.n296 163.367
R417 B.n298 B.n297 163.367
R418 B.n298 B.n145 163.367
R419 B.n302 B.n145 163.367
R420 B.n303 B.n302 163.367
R421 B.n304 B.n303 163.367
R422 B.n304 B.n141 163.367
R423 B.n309 B.n141 163.367
R424 B.n310 B.n309 163.367
R425 B.n311 B.n310 163.367
R426 B.n311 B.n139 163.367
R427 B.n315 B.n139 163.367
R428 B.n316 B.n315 163.367
R429 B.n317 B.n316 163.367
R430 B.n317 B.n137 163.367
R431 B.n324 B.n137 163.367
R432 B.n325 B.n324 163.367
R433 B.n326 B.n325 163.367
R434 B.n326 B.n135 163.367
R435 B.n330 B.n135 163.367
R436 B.n331 B.n330 163.367
R437 B.n332 B.n331 163.367
R438 B.n332 B.n133 163.367
R439 B.n336 B.n133 163.367
R440 B.n337 B.n336 163.367
R441 B.n338 B.n337 163.367
R442 B.n338 B.n131 163.367
R443 B.n342 B.n131 163.367
R444 B.n343 B.n342 163.367
R445 B.n344 B.n343 163.367
R446 B.n344 B.n129 163.367
R447 B.n348 B.n129 163.367
R448 B.n349 B.n348 163.367
R449 B.n350 B.n349 163.367
R450 B.n350 B.n127 163.367
R451 B.n354 B.n127 163.367
R452 B.n355 B.n354 163.367
R453 B.n356 B.n355 163.367
R454 B.n356 B.n125 163.367
R455 B.n360 B.n125 163.367
R456 B.n361 B.n360 163.367
R457 B.n362 B.n361 163.367
R458 B.n362 B.n123 163.367
R459 B.n366 B.n123 163.367
R460 B.n367 B.n366 163.367
R461 B.n368 B.n367 163.367
R462 B.n368 B.n121 163.367
R463 B.n372 B.n121 163.367
R464 B.n373 B.n372 163.367
R465 B.n374 B.n373 163.367
R466 B.n374 B.n119 163.367
R467 B.n378 B.n119 163.367
R468 B.n379 B.n378 163.367
R469 B.n380 B.n379 163.367
R470 B.n380 B.n117 163.367
R471 B.n384 B.n117 163.367
R472 B.n385 B.n384 163.367
R473 B.n386 B.n385 163.367
R474 B.n386 B.n115 163.367
R475 B.n390 B.n115 163.367
R476 B.n391 B.n390 163.367
R477 B.n392 B.n391 163.367
R478 B.n392 B.n113 163.367
R479 B.n396 B.n113 163.367
R480 B.n397 B.n396 163.367
R481 B.n398 B.n397 163.367
R482 B.n398 B.n111 163.367
R483 B.n402 B.n111 163.367
R484 B.n403 B.n402 163.367
R485 B.n404 B.n403 163.367
R486 B.n404 B.n109 163.367
R487 B.n408 B.n109 163.367
R488 B.n409 B.n408 163.367
R489 B.n410 B.n409 163.367
R490 B.n410 B.n107 163.367
R491 B.n414 B.n107 163.367
R492 B.n415 B.n414 163.367
R493 B.n482 B.n83 163.367
R494 B.n482 B.n481 163.367
R495 B.n481 B.n480 163.367
R496 B.n480 B.n85 163.367
R497 B.n476 B.n85 163.367
R498 B.n476 B.n475 163.367
R499 B.n475 B.n474 163.367
R500 B.n474 B.n87 163.367
R501 B.n470 B.n87 163.367
R502 B.n470 B.n469 163.367
R503 B.n469 B.n468 163.367
R504 B.n468 B.n89 163.367
R505 B.n464 B.n89 163.367
R506 B.n464 B.n463 163.367
R507 B.n463 B.n462 163.367
R508 B.n462 B.n91 163.367
R509 B.n458 B.n91 163.367
R510 B.n458 B.n457 163.367
R511 B.n457 B.n456 163.367
R512 B.n456 B.n93 163.367
R513 B.n452 B.n93 163.367
R514 B.n452 B.n451 163.367
R515 B.n451 B.n450 163.367
R516 B.n450 B.n95 163.367
R517 B.n446 B.n95 163.367
R518 B.n446 B.n445 163.367
R519 B.n445 B.n444 163.367
R520 B.n444 B.n97 163.367
R521 B.n440 B.n97 163.367
R522 B.n440 B.n439 163.367
R523 B.n439 B.n438 163.367
R524 B.n438 B.n99 163.367
R525 B.n434 B.n99 163.367
R526 B.n434 B.n433 163.367
R527 B.n433 B.n432 163.367
R528 B.n432 B.n101 163.367
R529 B.n428 B.n101 163.367
R530 B.n428 B.n427 163.367
R531 B.n427 B.n426 163.367
R532 B.n426 B.n103 163.367
R533 B.n422 B.n103 163.367
R534 B.n422 B.n421 163.367
R535 B.n421 B.n420 163.367
R536 B.n420 B.n105 163.367
R537 B.n416 B.n105 163.367
R538 B.n680 B.n13 163.367
R539 B.n680 B.n679 163.367
R540 B.n679 B.n678 163.367
R541 B.n678 B.n15 163.367
R542 B.n674 B.n15 163.367
R543 B.n674 B.n673 163.367
R544 B.n673 B.n672 163.367
R545 B.n672 B.n17 163.367
R546 B.n668 B.n17 163.367
R547 B.n668 B.n667 163.367
R548 B.n667 B.n666 163.367
R549 B.n666 B.n19 163.367
R550 B.n662 B.n19 163.367
R551 B.n662 B.n661 163.367
R552 B.n661 B.n660 163.367
R553 B.n660 B.n21 163.367
R554 B.n656 B.n21 163.367
R555 B.n656 B.n655 163.367
R556 B.n655 B.n654 163.367
R557 B.n654 B.n23 163.367
R558 B.n650 B.n23 163.367
R559 B.n650 B.n649 163.367
R560 B.n649 B.n648 163.367
R561 B.n648 B.n25 163.367
R562 B.n644 B.n25 163.367
R563 B.n644 B.n643 163.367
R564 B.n643 B.n642 163.367
R565 B.n642 B.n27 163.367
R566 B.n638 B.n27 163.367
R567 B.n638 B.n637 163.367
R568 B.n637 B.n636 163.367
R569 B.n636 B.n29 163.367
R570 B.n632 B.n29 163.367
R571 B.n632 B.n631 163.367
R572 B.n631 B.n630 163.367
R573 B.n630 B.n31 163.367
R574 B.n626 B.n31 163.367
R575 B.n626 B.n625 163.367
R576 B.n625 B.n624 163.367
R577 B.n624 B.n33 163.367
R578 B.n620 B.n33 163.367
R579 B.n620 B.n619 163.367
R580 B.n619 B.n618 163.367
R581 B.n618 B.n35 163.367
R582 B.n614 B.n35 163.367
R583 B.n614 B.n613 163.367
R584 B.n613 B.n612 163.367
R585 B.n612 B.n37 163.367
R586 B.n608 B.n37 163.367
R587 B.n608 B.n607 163.367
R588 B.n607 B.n606 163.367
R589 B.n606 B.n39 163.367
R590 B.n602 B.n39 163.367
R591 B.n602 B.n601 163.367
R592 B.n601 B.n600 163.367
R593 B.n600 B.n41 163.367
R594 B.n596 B.n41 163.367
R595 B.n596 B.n595 163.367
R596 B.n595 B.n594 163.367
R597 B.n594 B.n43 163.367
R598 B.n589 B.n43 163.367
R599 B.n589 B.n588 163.367
R600 B.n588 B.n587 163.367
R601 B.n587 B.n47 163.367
R602 B.n583 B.n47 163.367
R603 B.n583 B.n582 163.367
R604 B.n582 B.n581 163.367
R605 B.n581 B.n49 163.367
R606 B.n577 B.n49 163.367
R607 B.n577 B.n576 163.367
R608 B.n576 B.n53 163.367
R609 B.n572 B.n53 163.367
R610 B.n572 B.n571 163.367
R611 B.n571 B.n570 163.367
R612 B.n570 B.n55 163.367
R613 B.n566 B.n55 163.367
R614 B.n566 B.n565 163.367
R615 B.n565 B.n564 163.367
R616 B.n564 B.n57 163.367
R617 B.n560 B.n57 163.367
R618 B.n560 B.n559 163.367
R619 B.n559 B.n558 163.367
R620 B.n558 B.n59 163.367
R621 B.n554 B.n59 163.367
R622 B.n554 B.n553 163.367
R623 B.n553 B.n552 163.367
R624 B.n552 B.n61 163.367
R625 B.n548 B.n61 163.367
R626 B.n548 B.n547 163.367
R627 B.n547 B.n546 163.367
R628 B.n546 B.n63 163.367
R629 B.n542 B.n63 163.367
R630 B.n542 B.n541 163.367
R631 B.n541 B.n540 163.367
R632 B.n540 B.n65 163.367
R633 B.n536 B.n65 163.367
R634 B.n536 B.n535 163.367
R635 B.n535 B.n534 163.367
R636 B.n534 B.n67 163.367
R637 B.n530 B.n67 163.367
R638 B.n530 B.n529 163.367
R639 B.n529 B.n528 163.367
R640 B.n528 B.n69 163.367
R641 B.n524 B.n69 163.367
R642 B.n524 B.n523 163.367
R643 B.n523 B.n522 163.367
R644 B.n522 B.n71 163.367
R645 B.n518 B.n71 163.367
R646 B.n518 B.n517 163.367
R647 B.n517 B.n516 163.367
R648 B.n516 B.n73 163.367
R649 B.n512 B.n73 163.367
R650 B.n512 B.n511 163.367
R651 B.n511 B.n510 163.367
R652 B.n510 B.n75 163.367
R653 B.n506 B.n75 163.367
R654 B.n506 B.n505 163.367
R655 B.n505 B.n504 163.367
R656 B.n504 B.n77 163.367
R657 B.n500 B.n77 163.367
R658 B.n500 B.n499 163.367
R659 B.n499 B.n498 163.367
R660 B.n498 B.n79 163.367
R661 B.n494 B.n79 163.367
R662 B.n494 B.n493 163.367
R663 B.n493 B.n492 163.367
R664 B.n492 B.n81 163.367
R665 B.n488 B.n81 163.367
R666 B.n488 B.n487 163.367
R667 B.n487 B.n486 163.367
R668 B.n685 B.n684 163.367
R669 B.n686 B.n685 163.367
R670 B.n686 B.n11 163.367
R671 B.n690 B.n11 163.367
R672 B.n691 B.n690 163.367
R673 B.n692 B.n691 163.367
R674 B.n692 B.n9 163.367
R675 B.n696 B.n9 163.367
R676 B.n697 B.n696 163.367
R677 B.n698 B.n697 163.367
R678 B.n698 B.n7 163.367
R679 B.n702 B.n7 163.367
R680 B.n703 B.n702 163.367
R681 B.n704 B.n703 163.367
R682 B.n704 B.n5 163.367
R683 B.n708 B.n5 163.367
R684 B.n709 B.n708 163.367
R685 B.n710 B.n709 163.367
R686 B.n710 B.n3 163.367
R687 B.n714 B.n3 163.367
R688 B.n715 B.n714 163.367
R689 B.n184 B.n2 163.367
R690 B.n184 B.n183 163.367
R691 B.n188 B.n183 163.367
R692 B.n189 B.n188 163.367
R693 B.n190 B.n189 163.367
R694 B.n190 B.n181 163.367
R695 B.n194 B.n181 163.367
R696 B.n195 B.n194 163.367
R697 B.n196 B.n195 163.367
R698 B.n196 B.n179 163.367
R699 B.n200 B.n179 163.367
R700 B.n201 B.n200 163.367
R701 B.n202 B.n201 163.367
R702 B.n202 B.n177 163.367
R703 B.n206 B.n177 163.367
R704 B.n207 B.n206 163.367
R705 B.n208 B.n207 163.367
R706 B.n208 B.n175 163.367
R707 B.n212 B.n175 163.367
R708 B.n213 B.n212 163.367
R709 B.n214 B.n213 163.367
R710 B.n320 B.t7 125.947
R711 B.n50 B.t11 125.947
R712 B.n142 B.t1 125.922
R713 B.n44 B.t5 125.922
R714 B.n321 B.t8 107.135
R715 B.n51 B.t10 107.135
R716 B.n143 B.t2 107.111
R717 B.n45 B.t4 107.111
R718 B.n307 B.n143 59.5399
R719 B.n322 B.n321 59.5399
R720 B.n52 B.n51 59.5399
R721 B.n591 B.n45 59.5399
R722 B.n417 B.n106 28.5664
R723 B.n683 B.n682 28.5664
R724 B.n485 B.n484 28.5664
R725 B.n216 B.n215 28.5664
R726 B.n143 B.n142 18.8126
R727 B.n321 B.n320 18.8126
R728 B.n51 B.n50 18.8126
R729 B.n45 B.n44 18.8126
R730 B B.n717 18.0485
R731 B.n683 B.n12 10.6151
R732 B.n687 B.n12 10.6151
R733 B.n688 B.n687 10.6151
R734 B.n689 B.n688 10.6151
R735 B.n689 B.n10 10.6151
R736 B.n693 B.n10 10.6151
R737 B.n694 B.n693 10.6151
R738 B.n695 B.n694 10.6151
R739 B.n695 B.n8 10.6151
R740 B.n699 B.n8 10.6151
R741 B.n700 B.n699 10.6151
R742 B.n701 B.n700 10.6151
R743 B.n701 B.n6 10.6151
R744 B.n705 B.n6 10.6151
R745 B.n706 B.n705 10.6151
R746 B.n707 B.n706 10.6151
R747 B.n707 B.n4 10.6151
R748 B.n711 B.n4 10.6151
R749 B.n712 B.n711 10.6151
R750 B.n713 B.n712 10.6151
R751 B.n713 B.n0 10.6151
R752 B.n682 B.n681 10.6151
R753 B.n681 B.n14 10.6151
R754 B.n677 B.n14 10.6151
R755 B.n677 B.n676 10.6151
R756 B.n676 B.n675 10.6151
R757 B.n675 B.n16 10.6151
R758 B.n671 B.n16 10.6151
R759 B.n671 B.n670 10.6151
R760 B.n670 B.n669 10.6151
R761 B.n669 B.n18 10.6151
R762 B.n665 B.n18 10.6151
R763 B.n665 B.n664 10.6151
R764 B.n664 B.n663 10.6151
R765 B.n663 B.n20 10.6151
R766 B.n659 B.n20 10.6151
R767 B.n659 B.n658 10.6151
R768 B.n658 B.n657 10.6151
R769 B.n657 B.n22 10.6151
R770 B.n653 B.n22 10.6151
R771 B.n653 B.n652 10.6151
R772 B.n652 B.n651 10.6151
R773 B.n651 B.n24 10.6151
R774 B.n647 B.n24 10.6151
R775 B.n647 B.n646 10.6151
R776 B.n646 B.n645 10.6151
R777 B.n645 B.n26 10.6151
R778 B.n641 B.n26 10.6151
R779 B.n641 B.n640 10.6151
R780 B.n640 B.n639 10.6151
R781 B.n639 B.n28 10.6151
R782 B.n635 B.n28 10.6151
R783 B.n635 B.n634 10.6151
R784 B.n634 B.n633 10.6151
R785 B.n633 B.n30 10.6151
R786 B.n629 B.n30 10.6151
R787 B.n629 B.n628 10.6151
R788 B.n628 B.n627 10.6151
R789 B.n627 B.n32 10.6151
R790 B.n623 B.n32 10.6151
R791 B.n623 B.n622 10.6151
R792 B.n622 B.n621 10.6151
R793 B.n621 B.n34 10.6151
R794 B.n617 B.n34 10.6151
R795 B.n617 B.n616 10.6151
R796 B.n616 B.n615 10.6151
R797 B.n615 B.n36 10.6151
R798 B.n611 B.n36 10.6151
R799 B.n611 B.n610 10.6151
R800 B.n610 B.n609 10.6151
R801 B.n609 B.n38 10.6151
R802 B.n605 B.n38 10.6151
R803 B.n605 B.n604 10.6151
R804 B.n604 B.n603 10.6151
R805 B.n603 B.n40 10.6151
R806 B.n599 B.n40 10.6151
R807 B.n599 B.n598 10.6151
R808 B.n598 B.n597 10.6151
R809 B.n597 B.n42 10.6151
R810 B.n593 B.n42 10.6151
R811 B.n593 B.n592 10.6151
R812 B.n590 B.n46 10.6151
R813 B.n586 B.n46 10.6151
R814 B.n586 B.n585 10.6151
R815 B.n585 B.n584 10.6151
R816 B.n584 B.n48 10.6151
R817 B.n580 B.n48 10.6151
R818 B.n580 B.n579 10.6151
R819 B.n579 B.n578 10.6151
R820 B.n575 B.n574 10.6151
R821 B.n574 B.n573 10.6151
R822 B.n573 B.n54 10.6151
R823 B.n569 B.n54 10.6151
R824 B.n569 B.n568 10.6151
R825 B.n568 B.n567 10.6151
R826 B.n567 B.n56 10.6151
R827 B.n563 B.n56 10.6151
R828 B.n563 B.n562 10.6151
R829 B.n562 B.n561 10.6151
R830 B.n561 B.n58 10.6151
R831 B.n557 B.n58 10.6151
R832 B.n557 B.n556 10.6151
R833 B.n556 B.n555 10.6151
R834 B.n555 B.n60 10.6151
R835 B.n551 B.n60 10.6151
R836 B.n551 B.n550 10.6151
R837 B.n550 B.n549 10.6151
R838 B.n549 B.n62 10.6151
R839 B.n545 B.n62 10.6151
R840 B.n545 B.n544 10.6151
R841 B.n544 B.n543 10.6151
R842 B.n543 B.n64 10.6151
R843 B.n539 B.n64 10.6151
R844 B.n539 B.n538 10.6151
R845 B.n538 B.n537 10.6151
R846 B.n537 B.n66 10.6151
R847 B.n533 B.n66 10.6151
R848 B.n533 B.n532 10.6151
R849 B.n532 B.n531 10.6151
R850 B.n531 B.n68 10.6151
R851 B.n527 B.n68 10.6151
R852 B.n527 B.n526 10.6151
R853 B.n526 B.n525 10.6151
R854 B.n525 B.n70 10.6151
R855 B.n521 B.n70 10.6151
R856 B.n521 B.n520 10.6151
R857 B.n520 B.n519 10.6151
R858 B.n519 B.n72 10.6151
R859 B.n515 B.n72 10.6151
R860 B.n515 B.n514 10.6151
R861 B.n514 B.n513 10.6151
R862 B.n513 B.n74 10.6151
R863 B.n509 B.n74 10.6151
R864 B.n509 B.n508 10.6151
R865 B.n508 B.n507 10.6151
R866 B.n507 B.n76 10.6151
R867 B.n503 B.n76 10.6151
R868 B.n503 B.n502 10.6151
R869 B.n502 B.n501 10.6151
R870 B.n501 B.n78 10.6151
R871 B.n497 B.n78 10.6151
R872 B.n497 B.n496 10.6151
R873 B.n496 B.n495 10.6151
R874 B.n495 B.n80 10.6151
R875 B.n491 B.n80 10.6151
R876 B.n491 B.n490 10.6151
R877 B.n490 B.n489 10.6151
R878 B.n489 B.n82 10.6151
R879 B.n485 B.n82 10.6151
R880 B.n484 B.n483 10.6151
R881 B.n483 B.n84 10.6151
R882 B.n479 B.n84 10.6151
R883 B.n479 B.n478 10.6151
R884 B.n478 B.n477 10.6151
R885 B.n477 B.n86 10.6151
R886 B.n473 B.n86 10.6151
R887 B.n473 B.n472 10.6151
R888 B.n472 B.n471 10.6151
R889 B.n471 B.n88 10.6151
R890 B.n467 B.n88 10.6151
R891 B.n467 B.n466 10.6151
R892 B.n466 B.n465 10.6151
R893 B.n465 B.n90 10.6151
R894 B.n461 B.n90 10.6151
R895 B.n461 B.n460 10.6151
R896 B.n460 B.n459 10.6151
R897 B.n459 B.n92 10.6151
R898 B.n455 B.n92 10.6151
R899 B.n455 B.n454 10.6151
R900 B.n454 B.n453 10.6151
R901 B.n453 B.n94 10.6151
R902 B.n449 B.n94 10.6151
R903 B.n449 B.n448 10.6151
R904 B.n448 B.n447 10.6151
R905 B.n447 B.n96 10.6151
R906 B.n443 B.n96 10.6151
R907 B.n443 B.n442 10.6151
R908 B.n442 B.n441 10.6151
R909 B.n441 B.n98 10.6151
R910 B.n437 B.n98 10.6151
R911 B.n437 B.n436 10.6151
R912 B.n436 B.n435 10.6151
R913 B.n435 B.n100 10.6151
R914 B.n431 B.n100 10.6151
R915 B.n431 B.n430 10.6151
R916 B.n430 B.n429 10.6151
R917 B.n429 B.n102 10.6151
R918 B.n425 B.n102 10.6151
R919 B.n425 B.n424 10.6151
R920 B.n424 B.n423 10.6151
R921 B.n423 B.n104 10.6151
R922 B.n419 B.n104 10.6151
R923 B.n419 B.n418 10.6151
R924 B.n418 B.n417 10.6151
R925 B.n185 B.n1 10.6151
R926 B.n186 B.n185 10.6151
R927 B.n187 B.n186 10.6151
R928 B.n187 B.n182 10.6151
R929 B.n191 B.n182 10.6151
R930 B.n192 B.n191 10.6151
R931 B.n193 B.n192 10.6151
R932 B.n193 B.n180 10.6151
R933 B.n197 B.n180 10.6151
R934 B.n198 B.n197 10.6151
R935 B.n199 B.n198 10.6151
R936 B.n199 B.n178 10.6151
R937 B.n203 B.n178 10.6151
R938 B.n204 B.n203 10.6151
R939 B.n205 B.n204 10.6151
R940 B.n205 B.n176 10.6151
R941 B.n209 B.n176 10.6151
R942 B.n210 B.n209 10.6151
R943 B.n211 B.n210 10.6151
R944 B.n211 B.n174 10.6151
R945 B.n215 B.n174 10.6151
R946 B.n217 B.n216 10.6151
R947 B.n217 B.n172 10.6151
R948 B.n221 B.n172 10.6151
R949 B.n222 B.n221 10.6151
R950 B.n223 B.n222 10.6151
R951 B.n223 B.n170 10.6151
R952 B.n227 B.n170 10.6151
R953 B.n228 B.n227 10.6151
R954 B.n229 B.n228 10.6151
R955 B.n229 B.n168 10.6151
R956 B.n233 B.n168 10.6151
R957 B.n234 B.n233 10.6151
R958 B.n235 B.n234 10.6151
R959 B.n235 B.n166 10.6151
R960 B.n239 B.n166 10.6151
R961 B.n240 B.n239 10.6151
R962 B.n241 B.n240 10.6151
R963 B.n241 B.n164 10.6151
R964 B.n245 B.n164 10.6151
R965 B.n246 B.n245 10.6151
R966 B.n247 B.n246 10.6151
R967 B.n247 B.n162 10.6151
R968 B.n251 B.n162 10.6151
R969 B.n252 B.n251 10.6151
R970 B.n253 B.n252 10.6151
R971 B.n253 B.n160 10.6151
R972 B.n257 B.n160 10.6151
R973 B.n258 B.n257 10.6151
R974 B.n259 B.n258 10.6151
R975 B.n259 B.n158 10.6151
R976 B.n263 B.n158 10.6151
R977 B.n264 B.n263 10.6151
R978 B.n265 B.n264 10.6151
R979 B.n265 B.n156 10.6151
R980 B.n269 B.n156 10.6151
R981 B.n270 B.n269 10.6151
R982 B.n271 B.n270 10.6151
R983 B.n271 B.n154 10.6151
R984 B.n275 B.n154 10.6151
R985 B.n276 B.n275 10.6151
R986 B.n277 B.n276 10.6151
R987 B.n277 B.n152 10.6151
R988 B.n281 B.n152 10.6151
R989 B.n282 B.n281 10.6151
R990 B.n283 B.n282 10.6151
R991 B.n283 B.n150 10.6151
R992 B.n287 B.n150 10.6151
R993 B.n288 B.n287 10.6151
R994 B.n289 B.n288 10.6151
R995 B.n289 B.n148 10.6151
R996 B.n293 B.n148 10.6151
R997 B.n294 B.n293 10.6151
R998 B.n295 B.n294 10.6151
R999 B.n295 B.n146 10.6151
R1000 B.n299 B.n146 10.6151
R1001 B.n300 B.n299 10.6151
R1002 B.n301 B.n300 10.6151
R1003 B.n301 B.n144 10.6151
R1004 B.n305 B.n144 10.6151
R1005 B.n306 B.n305 10.6151
R1006 B.n308 B.n140 10.6151
R1007 B.n312 B.n140 10.6151
R1008 B.n313 B.n312 10.6151
R1009 B.n314 B.n313 10.6151
R1010 B.n314 B.n138 10.6151
R1011 B.n318 B.n138 10.6151
R1012 B.n319 B.n318 10.6151
R1013 B.n323 B.n319 10.6151
R1014 B.n327 B.n136 10.6151
R1015 B.n328 B.n327 10.6151
R1016 B.n329 B.n328 10.6151
R1017 B.n329 B.n134 10.6151
R1018 B.n333 B.n134 10.6151
R1019 B.n334 B.n333 10.6151
R1020 B.n335 B.n334 10.6151
R1021 B.n335 B.n132 10.6151
R1022 B.n339 B.n132 10.6151
R1023 B.n340 B.n339 10.6151
R1024 B.n341 B.n340 10.6151
R1025 B.n341 B.n130 10.6151
R1026 B.n345 B.n130 10.6151
R1027 B.n346 B.n345 10.6151
R1028 B.n347 B.n346 10.6151
R1029 B.n347 B.n128 10.6151
R1030 B.n351 B.n128 10.6151
R1031 B.n352 B.n351 10.6151
R1032 B.n353 B.n352 10.6151
R1033 B.n353 B.n126 10.6151
R1034 B.n357 B.n126 10.6151
R1035 B.n358 B.n357 10.6151
R1036 B.n359 B.n358 10.6151
R1037 B.n359 B.n124 10.6151
R1038 B.n363 B.n124 10.6151
R1039 B.n364 B.n363 10.6151
R1040 B.n365 B.n364 10.6151
R1041 B.n365 B.n122 10.6151
R1042 B.n369 B.n122 10.6151
R1043 B.n370 B.n369 10.6151
R1044 B.n371 B.n370 10.6151
R1045 B.n371 B.n120 10.6151
R1046 B.n375 B.n120 10.6151
R1047 B.n376 B.n375 10.6151
R1048 B.n377 B.n376 10.6151
R1049 B.n377 B.n118 10.6151
R1050 B.n381 B.n118 10.6151
R1051 B.n382 B.n381 10.6151
R1052 B.n383 B.n382 10.6151
R1053 B.n383 B.n116 10.6151
R1054 B.n387 B.n116 10.6151
R1055 B.n388 B.n387 10.6151
R1056 B.n389 B.n388 10.6151
R1057 B.n389 B.n114 10.6151
R1058 B.n393 B.n114 10.6151
R1059 B.n394 B.n393 10.6151
R1060 B.n395 B.n394 10.6151
R1061 B.n395 B.n112 10.6151
R1062 B.n399 B.n112 10.6151
R1063 B.n400 B.n399 10.6151
R1064 B.n401 B.n400 10.6151
R1065 B.n401 B.n110 10.6151
R1066 B.n405 B.n110 10.6151
R1067 B.n406 B.n405 10.6151
R1068 B.n407 B.n406 10.6151
R1069 B.n407 B.n108 10.6151
R1070 B.n411 B.n108 10.6151
R1071 B.n412 B.n411 10.6151
R1072 B.n413 B.n412 10.6151
R1073 B.n413 B.n106 10.6151
R1074 B.n717 B.n0 8.11757
R1075 B.n717 B.n1 8.11757
R1076 B.n591 B.n590 6.5566
R1077 B.n578 B.n52 6.5566
R1078 B.n308 B.n307 6.5566
R1079 B.n323 B.n322 6.5566
R1080 B.n592 B.n591 4.05904
R1081 B.n575 B.n52 4.05904
R1082 B.n307 B.n306 4.05904
R1083 B.n322 B.n136 4.05904
R1084 VP.n3 VP.t6 781.83
R1085 VP.n1 VP.t2 755.009
R1086 VP.n10 VP.t3 755.009
R1087 VP.n11 VP.t5 755.009
R1088 VP.n12 VP.t0 755.009
R1089 VP.n6 VP.t7 755.009
R1090 VP.n5 VP.t4 755.009
R1091 VP.n4 VP.t1 755.009
R1092 VP.n13 VP.n12 161.3
R1093 VP.n7 VP.n6 161.3
R1094 VP.n8 VP.n1 161.3
R1095 VP.n5 VP.n2 80.6037
R1096 VP.n11 VP.n0 80.6037
R1097 VP.n10 VP.n9 80.6037
R1098 VP.n10 VP.n1 48.2005
R1099 VP.n11 VP.n10 48.2005
R1100 VP.n12 VP.n11 48.2005
R1101 VP.n6 VP.n5 48.2005
R1102 VP.n5 VP.n4 48.2005
R1103 VP.n8 VP.n7 46.6747
R1104 VP.n3 VP.n2 45.2318
R1105 VP.n4 VP.n3 13.3799
R1106 VP.n9 VP.n0 0.380177
R1107 VP.n7 VP.n2 0.285035
R1108 VP.n9 VP.n8 0.285035
R1109 VP.n13 VP.n0 0.285035
R1110 VP VP.n13 0.0516364
R1111 VTAIL.n11 VTAIL.t14 56.5936
R1112 VTAIL.n10 VTAIL.t4 56.5936
R1113 VTAIL.n7 VTAIL.t0 56.5936
R1114 VTAIL.n15 VTAIL.t1 56.5925
R1115 VTAIL.n2 VTAIL.t3 56.5925
R1116 VTAIL.n3 VTAIL.t11 56.5925
R1117 VTAIL.n6 VTAIL.t12 56.5925
R1118 VTAIL.n14 VTAIL.t10 56.5924
R1119 VTAIL.n13 VTAIL.n12 54.8279
R1120 VTAIL.n9 VTAIL.n8 54.8279
R1121 VTAIL.n1 VTAIL.n0 54.8277
R1122 VTAIL.n5 VTAIL.n4 54.8277
R1123 VTAIL.n15 VTAIL.n14 29.0738
R1124 VTAIL.n7 VTAIL.n6 29.0738
R1125 VTAIL.n0 VTAIL.t5 1.76612
R1126 VTAIL.n0 VTAIL.t6 1.76612
R1127 VTAIL.n4 VTAIL.t13 1.76612
R1128 VTAIL.n4 VTAIL.t15 1.76612
R1129 VTAIL.n12 VTAIL.t8 1.76612
R1130 VTAIL.n12 VTAIL.t9 1.76612
R1131 VTAIL.n8 VTAIL.t2 1.76612
R1132 VTAIL.n8 VTAIL.t7 1.76612
R1133 VTAIL.n9 VTAIL.n7 0.836707
R1134 VTAIL.n10 VTAIL.n9 0.836707
R1135 VTAIL.n13 VTAIL.n11 0.836707
R1136 VTAIL.n14 VTAIL.n13 0.836707
R1137 VTAIL.n6 VTAIL.n5 0.836707
R1138 VTAIL.n5 VTAIL.n3 0.836707
R1139 VTAIL.n2 VTAIL.n1 0.836707
R1140 VTAIL VTAIL.n15 0.778517
R1141 VTAIL.n11 VTAIL.n10 0.470328
R1142 VTAIL.n3 VTAIL.n2 0.470328
R1143 VTAIL VTAIL.n1 0.0586897
R1144 VDD1 VDD1.n0 71.983
R1145 VDD1.n3 VDD1.n2 71.8693
R1146 VDD1.n3 VDD1.n1 71.8693
R1147 VDD1.n5 VDD1.n4 71.5056
R1148 VDD1.n5 VDD1.n3 43.9319
R1149 VDD1.n4 VDD1.t3 1.76612
R1150 VDD1.n4 VDD1.t0 1.76612
R1151 VDD1.n0 VDD1.t1 1.76612
R1152 VDD1.n0 VDD1.t6 1.76612
R1153 VDD1.n2 VDD1.t2 1.76612
R1154 VDD1.n2 VDD1.t7 1.76612
R1155 VDD1.n1 VDD1.t5 1.76612
R1156 VDD1.n1 VDD1.t4 1.76612
R1157 VDD1 VDD1.n5 0.360414
R1158 VN.n1 VN.t1 781.83
R1159 VN.n7 VN.t2 781.83
R1160 VN.n2 VN.t7 755.009
R1161 VN.n3 VN.t6 755.009
R1162 VN.n4 VN.t3 755.009
R1163 VN.n8 VN.t5 755.009
R1164 VN.n9 VN.t0 755.009
R1165 VN.n10 VN.t4 755.009
R1166 VN.n5 VN.n4 161.3
R1167 VN.n11 VN.n10 161.3
R1168 VN.n9 VN.n6 80.6037
R1169 VN.n3 VN.n0 80.6037
R1170 VN.n3 VN.n2 48.2005
R1171 VN.n4 VN.n3 48.2005
R1172 VN.n9 VN.n8 48.2005
R1173 VN.n10 VN.n9 48.2005
R1174 VN VN.n11 47.0554
R1175 VN.n7 VN.n6 45.2318
R1176 VN.n1 VN.n0 45.2318
R1177 VN.n8 VN.n7 13.3799
R1178 VN.n2 VN.n1 13.3799
R1179 VN.n11 VN.n6 0.285035
R1180 VN.n5 VN.n0 0.285035
R1181 VN VN.n5 0.0516364
R1182 VDD2.n2 VDD2.n1 71.8693
R1183 VDD2.n2 VDD2.n0 71.8693
R1184 VDD2 VDD2.n5 71.8655
R1185 VDD2.n4 VDD2.n3 71.5067
R1186 VDD2.n4 VDD2.n2 43.3489
R1187 VDD2.n5 VDD2.t2 1.76612
R1188 VDD2.n5 VDD2.t5 1.76612
R1189 VDD2.n3 VDD2.t3 1.76612
R1190 VDD2.n3 VDD2.t7 1.76612
R1191 VDD2.n1 VDD2.t1 1.76612
R1192 VDD2.n1 VDD2.t4 1.76612
R1193 VDD2.n0 VDD2.t6 1.76612
R1194 VDD2.n0 VDD2.t0 1.76612
R1195 VDD2 VDD2.n4 0.476793
C0 VDD2 B 1.25919f
C1 VN VP 6.44934f
C2 w_n1940_n4650# B 8.91404f
C3 VTAIL VP 7.35309f
C4 VTAIL VN 7.33898f
C5 VDD1 B 1.22438f
C6 VDD2 VP 0.311147f
C7 VDD2 VN 7.858171f
C8 w_n1940_n4650# VP 3.75427f
C9 w_n1940_n4650# VN 3.5082f
C10 VDD2 VTAIL 16.6335f
C11 VTAIL w_n1940_n4650# 5.84167f
C12 VDD1 VP 8.02069f
C13 VDD1 VN 0.148226f
C14 VTAIL VDD1 16.5922f
C15 VDD2 w_n1940_n4650# 1.48234f
C16 VDD2 VDD1 0.796903f
C17 VDD1 w_n1940_n4650# 1.44998f
C18 B VP 1.24443f
C19 B VN 0.842369f
C20 VTAIL B 5.50248f
C21 VDD2 VSUBS 1.492766f
C22 VDD1 VSUBS 1.78749f
C23 VTAIL VSUBS 1.123947f
C24 VN VSUBS 5.16188f
C25 VP VSUBS 1.829904f
C26 B VSUBS 3.353748f
C27 w_n1940_n4650# VSUBS 0.110277p
C28 VDD2.t6 VSUBS 0.407561f
C29 VDD2.t0 VSUBS 0.407561f
C30 VDD2.n0 VSUBS 3.42322f
C31 VDD2.t1 VSUBS 0.407561f
C32 VDD2.t4 VSUBS 0.407561f
C33 VDD2.n1 VSUBS 3.42322f
C34 VDD2.n2 VSUBS 3.43629f
C35 VDD2.t3 VSUBS 0.407561f
C36 VDD2.t7 VSUBS 0.407561f
C37 VDD2.n3 VSUBS 3.41994f
C38 VDD2.n4 VSUBS 3.39281f
C39 VDD2.t2 VSUBS 0.407561f
C40 VDD2.t5 VSUBS 0.407561f
C41 VDD2.n5 VSUBS 3.42318f
C42 VN.n0 VSUBS 0.260245f
C43 VN.t1 VSUBS 1.77037f
C44 VN.n1 VSUBS 0.638709f
C45 VN.t7 VSUBS 1.74773f
C46 VN.n2 VSUBS 0.6716f
C47 VN.t6 VSUBS 1.74773f
C48 VN.n3 VSUBS 0.6716f
C49 VN.t3 VSUBS 1.74773f
C50 VN.n4 VSUBS 0.659727f
C51 VN.n5 VSUBS 0.058044f
C52 VN.n6 VSUBS 0.260245f
C53 VN.t5 VSUBS 1.74773f
C54 VN.t2 VSUBS 1.77037f
C55 VN.n7 VSUBS 0.638709f
C56 VN.n8 VSUBS 0.6716f
C57 VN.t0 VSUBS 1.74773f
C58 VN.n9 VSUBS 0.6716f
C59 VN.t4 VSUBS 1.74773f
C60 VN.n10 VSUBS 0.659727f
C61 VN.n11 VSUBS 2.61176f
C62 VDD1.t1 VSUBS 0.407503f
C63 VDD1.t6 VSUBS 0.407503f
C64 VDD1.n0 VSUBS 3.42382f
C65 VDD1.t5 VSUBS 0.407503f
C66 VDD1.t4 VSUBS 0.407503f
C67 VDD1.n1 VSUBS 3.42274f
C68 VDD1.t2 VSUBS 0.407503f
C69 VDD1.t7 VSUBS 0.407503f
C70 VDD1.n2 VSUBS 3.42274f
C71 VDD1.n3 VSUBS 3.4952f
C72 VDD1.t3 VSUBS 0.407503f
C73 VDD1.t0 VSUBS 0.407503f
C74 VDD1.n4 VSUBS 3.41945f
C75 VDD1.n5 VSUBS 3.42591f
C76 VTAIL.t5 VSUBS 0.354717f
C77 VTAIL.t6 VSUBS 0.354717f
C78 VTAIL.n0 VSUBS 2.83777f
C79 VTAIL.n1 VSUBS 0.636587f
C80 VTAIL.t3 VSUBS 3.69754f
C81 VTAIL.n2 VSUBS 0.776568f
C82 VTAIL.t11 VSUBS 3.69754f
C83 VTAIL.n3 VSUBS 0.776568f
C84 VTAIL.t13 VSUBS 0.354717f
C85 VTAIL.t15 VSUBS 0.354717f
C86 VTAIL.n4 VSUBS 2.83777f
C87 VTAIL.n5 VSUBS 0.697712f
C88 VTAIL.t12 VSUBS 3.69754f
C89 VTAIL.n6 VSUBS 2.38344f
C90 VTAIL.t0 VSUBS 3.69754f
C91 VTAIL.n7 VSUBS 2.38344f
C92 VTAIL.t2 VSUBS 0.354717f
C93 VTAIL.t7 VSUBS 0.354717f
C94 VTAIL.n8 VSUBS 2.83778f
C95 VTAIL.n9 VSUBS 0.697706f
C96 VTAIL.t4 VSUBS 3.69754f
C97 VTAIL.n10 VSUBS 0.77657f
C98 VTAIL.t14 VSUBS 3.69754f
C99 VTAIL.n11 VSUBS 0.77657f
C100 VTAIL.t8 VSUBS 0.354717f
C101 VTAIL.t9 VSUBS 0.354717f
C102 VTAIL.n12 VSUBS 2.83778f
C103 VTAIL.n13 VSUBS 0.697706f
C104 VTAIL.t10 VSUBS 3.69752f
C105 VTAIL.n14 VSUBS 2.38346f
C106 VTAIL.t1 VSUBS 3.69754f
C107 VTAIL.n15 VSUBS 2.37887f
C108 VP.n0 VSUBS 0.089149f
C109 VP.t2 VSUBS 1.78779f
C110 VP.n1 VSUBS 0.674846f
C111 VP.n2 VSUBS 0.26621f
C112 VP.t7 VSUBS 1.78779f
C113 VP.t4 VSUBS 1.78779f
C114 VP.t1 VSUBS 1.78779f
C115 VP.t6 VSUBS 1.81094f
C116 VP.n3 VSUBS 0.653346f
C117 VP.n4 VSUBS 0.686992f
C118 VP.n5 VSUBS 0.686992f
C119 VP.n6 VSUBS 0.674846f
C120 VP.n7 VSUBS 2.63669f
C121 VP.n8 VSUBS 2.67792f
C122 VP.n9 VSUBS 0.089149f
C123 VP.t3 VSUBS 1.78779f
C124 VP.n10 VSUBS 0.686992f
C125 VP.t5 VSUBS 1.78779f
C126 VP.n11 VSUBS 0.686992f
C127 VP.t0 VSUBS 1.78779f
C128 VP.n12 VSUBS 0.674846f
C129 VP.n13 VSUBS 0.059375f
C130 B.n0 VSUBS 0.006831f
C131 B.n1 VSUBS 0.006831f
C132 B.n2 VSUBS 0.010102f
C133 B.n3 VSUBS 0.007742f
C134 B.n4 VSUBS 0.007742f
C135 B.n5 VSUBS 0.007742f
C136 B.n6 VSUBS 0.007742f
C137 B.n7 VSUBS 0.007742f
C138 B.n8 VSUBS 0.007742f
C139 B.n9 VSUBS 0.007742f
C140 B.n10 VSUBS 0.007742f
C141 B.n11 VSUBS 0.007742f
C142 B.n12 VSUBS 0.007742f
C143 B.n13 VSUBS 0.017221f
C144 B.n14 VSUBS 0.007742f
C145 B.n15 VSUBS 0.007742f
C146 B.n16 VSUBS 0.007742f
C147 B.n17 VSUBS 0.007742f
C148 B.n18 VSUBS 0.007742f
C149 B.n19 VSUBS 0.007742f
C150 B.n20 VSUBS 0.007742f
C151 B.n21 VSUBS 0.007742f
C152 B.n22 VSUBS 0.007742f
C153 B.n23 VSUBS 0.007742f
C154 B.n24 VSUBS 0.007742f
C155 B.n25 VSUBS 0.007742f
C156 B.n26 VSUBS 0.007742f
C157 B.n27 VSUBS 0.007742f
C158 B.n28 VSUBS 0.007742f
C159 B.n29 VSUBS 0.007742f
C160 B.n30 VSUBS 0.007742f
C161 B.n31 VSUBS 0.007742f
C162 B.n32 VSUBS 0.007742f
C163 B.n33 VSUBS 0.007742f
C164 B.n34 VSUBS 0.007742f
C165 B.n35 VSUBS 0.007742f
C166 B.n36 VSUBS 0.007742f
C167 B.n37 VSUBS 0.007742f
C168 B.n38 VSUBS 0.007742f
C169 B.n39 VSUBS 0.007742f
C170 B.n40 VSUBS 0.007742f
C171 B.n41 VSUBS 0.007742f
C172 B.n42 VSUBS 0.007742f
C173 B.n43 VSUBS 0.007742f
C174 B.t4 VSUBS 0.688399f
C175 B.t5 VSUBS 0.697331f
C176 B.t3 VSUBS 0.522019f
C177 B.n44 VSUBS 0.198104f
C178 B.n45 VSUBS 0.070824f
C179 B.n46 VSUBS 0.007742f
C180 B.n47 VSUBS 0.007742f
C181 B.n48 VSUBS 0.007742f
C182 B.n49 VSUBS 0.007742f
C183 B.t10 VSUBS 0.688372f
C184 B.t11 VSUBS 0.697306f
C185 B.t9 VSUBS 0.522019f
C186 B.n50 VSUBS 0.198128f
C187 B.n51 VSUBS 0.07085f
C188 B.n52 VSUBS 0.017936f
C189 B.n53 VSUBS 0.007742f
C190 B.n54 VSUBS 0.007742f
C191 B.n55 VSUBS 0.007742f
C192 B.n56 VSUBS 0.007742f
C193 B.n57 VSUBS 0.007742f
C194 B.n58 VSUBS 0.007742f
C195 B.n59 VSUBS 0.007742f
C196 B.n60 VSUBS 0.007742f
C197 B.n61 VSUBS 0.007742f
C198 B.n62 VSUBS 0.007742f
C199 B.n63 VSUBS 0.007742f
C200 B.n64 VSUBS 0.007742f
C201 B.n65 VSUBS 0.007742f
C202 B.n66 VSUBS 0.007742f
C203 B.n67 VSUBS 0.007742f
C204 B.n68 VSUBS 0.007742f
C205 B.n69 VSUBS 0.007742f
C206 B.n70 VSUBS 0.007742f
C207 B.n71 VSUBS 0.007742f
C208 B.n72 VSUBS 0.007742f
C209 B.n73 VSUBS 0.007742f
C210 B.n74 VSUBS 0.007742f
C211 B.n75 VSUBS 0.007742f
C212 B.n76 VSUBS 0.007742f
C213 B.n77 VSUBS 0.007742f
C214 B.n78 VSUBS 0.007742f
C215 B.n79 VSUBS 0.007742f
C216 B.n80 VSUBS 0.007742f
C217 B.n81 VSUBS 0.007742f
C218 B.n82 VSUBS 0.007742f
C219 B.n83 VSUBS 0.016022f
C220 B.n84 VSUBS 0.007742f
C221 B.n85 VSUBS 0.007742f
C222 B.n86 VSUBS 0.007742f
C223 B.n87 VSUBS 0.007742f
C224 B.n88 VSUBS 0.007742f
C225 B.n89 VSUBS 0.007742f
C226 B.n90 VSUBS 0.007742f
C227 B.n91 VSUBS 0.007742f
C228 B.n92 VSUBS 0.007742f
C229 B.n93 VSUBS 0.007742f
C230 B.n94 VSUBS 0.007742f
C231 B.n95 VSUBS 0.007742f
C232 B.n96 VSUBS 0.007742f
C233 B.n97 VSUBS 0.007742f
C234 B.n98 VSUBS 0.007742f
C235 B.n99 VSUBS 0.007742f
C236 B.n100 VSUBS 0.007742f
C237 B.n101 VSUBS 0.007742f
C238 B.n102 VSUBS 0.007742f
C239 B.n103 VSUBS 0.007742f
C240 B.n104 VSUBS 0.007742f
C241 B.n105 VSUBS 0.007742f
C242 B.n106 VSUBS 0.016175f
C243 B.n107 VSUBS 0.007742f
C244 B.n108 VSUBS 0.007742f
C245 B.n109 VSUBS 0.007742f
C246 B.n110 VSUBS 0.007742f
C247 B.n111 VSUBS 0.007742f
C248 B.n112 VSUBS 0.007742f
C249 B.n113 VSUBS 0.007742f
C250 B.n114 VSUBS 0.007742f
C251 B.n115 VSUBS 0.007742f
C252 B.n116 VSUBS 0.007742f
C253 B.n117 VSUBS 0.007742f
C254 B.n118 VSUBS 0.007742f
C255 B.n119 VSUBS 0.007742f
C256 B.n120 VSUBS 0.007742f
C257 B.n121 VSUBS 0.007742f
C258 B.n122 VSUBS 0.007742f
C259 B.n123 VSUBS 0.007742f
C260 B.n124 VSUBS 0.007742f
C261 B.n125 VSUBS 0.007742f
C262 B.n126 VSUBS 0.007742f
C263 B.n127 VSUBS 0.007742f
C264 B.n128 VSUBS 0.007742f
C265 B.n129 VSUBS 0.007742f
C266 B.n130 VSUBS 0.007742f
C267 B.n131 VSUBS 0.007742f
C268 B.n132 VSUBS 0.007742f
C269 B.n133 VSUBS 0.007742f
C270 B.n134 VSUBS 0.007742f
C271 B.n135 VSUBS 0.007742f
C272 B.n136 VSUBS 0.005351f
C273 B.n137 VSUBS 0.007742f
C274 B.n138 VSUBS 0.007742f
C275 B.n139 VSUBS 0.007742f
C276 B.n140 VSUBS 0.007742f
C277 B.n141 VSUBS 0.007742f
C278 B.t2 VSUBS 0.688399f
C279 B.t1 VSUBS 0.697331f
C280 B.t0 VSUBS 0.522019f
C281 B.n142 VSUBS 0.198104f
C282 B.n143 VSUBS 0.070824f
C283 B.n144 VSUBS 0.007742f
C284 B.n145 VSUBS 0.007742f
C285 B.n146 VSUBS 0.007742f
C286 B.n147 VSUBS 0.007742f
C287 B.n148 VSUBS 0.007742f
C288 B.n149 VSUBS 0.007742f
C289 B.n150 VSUBS 0.007742f
C290 B.n151 VSUBS 0.007742f
C291 B.n152 VSUBS 0.007742f
C292 B.n153 VSUBS 0.007742f
C293 B.n154 VSUBS 0.007742f
C294 B.n155 VSUBS 0.007742f
C295 B.n156 VSUBS 0.007742f
C296 B.n157 VSUBS 0.007742f
C297 B.n158 VSUBS 0.007742f
C298 B.n159 VSUBS 0.007742f
C299 B.n160 VSUBS 0.007742f
C300 B.n161 VSUBS 0.007742f
C301 B.n162 VSUBS 0.007742f
C302 B.n163 VSUBS 0.007742f
C303 B.n164 VSUBS 0.007742f
C304 B.n165 VSUBS 0.007742f
C305 B.n166 VSUBS 0.007742f
C306 B.n167 VSUBS 0.007742f
C307 B.n168 VSUBS 0.007742f
C308 B.n169 VSUBS 0.007742f
C309 B.n170 VSUBS 0.007742f
C310 B.n171 VSUBS 0.007742f
C311 B.n172 VSUBS 0.007742f
C312 B.n173 VSUBS 0.017221f
C313 B.n174 VSUBS 0.007742f
C314 B.n175 VSUBS 0.007742f
C315 B.n176 VSUBS 0.007742f
C316 B.n177 VSUBS 0.007742f
C317 B.n178 VSUBS 0.007742f
C318 B.n179 VSUBS 0.007742f
C319 B.n180 VSUBS 0.007742f
C320 B.n181 VSUBS 0.007742f
C321 B.n182 VSUBS 0.007742f
C322 B.n183 VSUBS 0.007742f
C323 B.n184 VSUBS 0.007742f
C324 B.n185 VSUBS 0.007742f
C325 B.n186 VSUBS 0.007742f
C326 B.n187 VSUBS 0.007742f
C327 B.n188 VSUBS 0.007742f
C328 B.n189 VSUBS 0.007742f
C329 B.n190 VSUBS 0.007742f
C330 B.n191 VSUBS 0.007742f
C331 B.n192 VSUBS 0.007742f
C332 B.n193 VSUBS 0.007742f
C333 B.n194 VSUBS 0.007742f
C334 B.n195 VSUBS 0.007742f
C335 B.n196 VSUBS 0.007742f
C336 B.n197 VSUBS 0.007742f
C337 B.n198 VSUBS 0.007742f
C338 B.n199 VSUBS 0.007742f
C339 B.n200 VSUBS 0.007742f
C340 B.n201 VSUBS 0.007742f
C341 B.n202 VSUBS 0.007742f
C342 B.n203 VSUBS 0.007742f
C343 B.n204 VSUBS 0.007742f
C344 B.n205 VSUBS 0.007742f
C345 B.n206 VSUBS 0.007742f
C346 B.n207 VSUBS 0.007742f
C347 B.n208 VSUBS 0.007742f
C348 B.n209 VSUBS 0.007742f
C349 B.n210 VSUBS 0.007742f
C350 B.n211 VSUBS 0.007742f
C351 B.n212 VSUBS 0.007742f
C352 B.n213 VSUBS 0.007742f
C353 B.n214 VSUBS 0.016022f
C354 B.n215 VSUBS 0.016022f
C355 B.n216 VSUBS 0.017221f
C356 B.n217 VSUBS 0.007742f
C357 B.n218 VSUBS 0.007742f
C358 B.n219 VSUBS 0.007742f
C359 B.n220 VSUBS 0.007742f
C360 B.n221 VSUBS 0.007742f
C361 B.n222 VSUBS 0.007742f
C362 B.n223 VSUBS 0.007742f
C363 B.n224 VSUBS 0.007742f
C364 B.n225 VSUBS 0.007742f
C365 B.n226 VSUBS 0.007742f
C366 B.n227 VSUBS 0.007742f
C367 B.n228 VSUBS 0.007742f
C368 B.n229 VSUBS 0.007742f
C369 B.n230 VSUBS 0.007742f
C370 B.n231 VSUBS 0.007742f
C371 B.n232 VSUBS 0.007742f
C372 B.n233 VSUBS 0.007742f
C373 B.n234 VSUBS 0.007742f
C374 B.n235 VSUBS 0.007742f
C375 B.n236 VSUBS 0.007742f
C376 B.n237 VSUBS 0.007742f
C377 B.n238 VSUBS 0.007742f
C378 B.n239 VSUBS 0.007742f
C379 B.n240 VSUBS 0.007742f
C380 B.n241 VSUBS 0.007742f
C381 B.n242 VSUBS 0.007742f
C382 B.n243 VSUBS 0.007742f
C383 B.n244 VSUBS 0.007742f
C384 B.n245 VSUBS 0.007742f
C385 B.n246 VSUBS 0.007742f
C386 B.n247 VSUBS 0.007742f
C387 B.n248 VSUBS 0.007742f
C388 B.n249 VSUBS 0.007742f
C389 B.n250 VSUBS 0.007742f
C390 B.n251 VSUBS 0.007742f
C391 B.n252 VSUBS 0.007742f
C392 B.n253 VSUBS 0.007742f
C393 B.n254 VSUBS 0.007742f
C394 B.n255 VSUBS 0.007742f
C395 B.n256 VSUBS 0.007742f
C396 B.n257 VSUBS 0.007742f
C397 B.n258 VSUBS 0.007742f
C398 B.n259 VSUBS 0.007742f
C399 B.n260 VSUBS 0.007742f
C400 B.n261 VSUBS 0.007742f
C401 B.n262 VSUBS 0.007742f
C402 B.n263 VSUBS 0.007742f
C403 B.n264 VSUBS 0.007742f
C404 B.n265 VSUBS 0.007742f
C405 B.n266 VSUBS 0.007742f
C406 B.n267 VSUBS 0.007742f
C407 B.n268 VSUBS 0.007742f
C408 B.n269 VSUBS 0.007742f
C409 B.n270 VSUBS 0.007742f
C410 B.n271 VSUBS 0.007742f
C411 B.n272 VSUBS 0.007742f
C412 B.n273 VSUBS 0.007742f
C413 B.n274 VSUBS 0.007742f
C414 B.n275 VSUBS 0.007742f
C415 B.n276 VSUBS 0.007742f
C416 B.n277 VSUBS 0.007742f
C417 B.n278 VSUBS 0.007742f
C418 B.n279 VSUBS 0.007742f
C419 B.n280 VSUBS 0.007742f
C420 B.n281 VSUBS 0.007742f
C421 B.n282 VSUBS 0.007742f
C422 B.n283 VSUBS 0.007742f
C423 B.n284 VSUBS 0.007742f
C424 B.n285 VSUBS 0.007742f
C425 B.n286 VSUBS 0.007742f
C426 B.n287 VSUBS 0.007742f
C427 B.n288 VSUBS 0.007742f
C428 B.n289 VSUBS 0.007742f
C429 B.n290 VSUBS 0.007742f
C430 B.n291 VSUBS 0.007742f
C431 B.n292 VSUBS 0.007742f
C432 B.n293 VSUBS 0.007742f
C433 B.n294 VSUBS 0.007742f
C434 B.n295 VSUBS 0.007742f
C435 B.n296 VSUBS 0.007742f
C436 B.n297 VSUBS 0.007742f
C437 B.n298 VSUBS 0.007742f
C438 B.n299 VSUBS 0.007742f
C439 B.n300 VSUBS 0.007742f
C440 B.n301 VSUBS 0.007742f
C441 B.n302 VSUBS 0.007742f
C442 B.n303 VSUBS 0.007742f
C443 B.n304 VSUBS 0.007742f
C444 B.n305 VSUBS 0.007742f
C445 B.n306 VSUBS 0.005351f
C446 B.n307 VSUBS 0.017936f
C447 B.n308 VSUBS 0.006262f
C448 B.n309 VSUBS 0.007742f
C449 B.n310 VSUBS 0.007742f
C450 B.n311 VSUBS 0.007742f
C451 B.n312 VSUBS 0.007742f
C452 B.n313 VSUBS 0.007742f
C453 B.n314 VSUBS 0.007742f
C454 B.n315 VSUBS 0.007742f
C455 B.n316 VSUBS 0.007742f
C456 B.n317 VSUBS 0.007742f
C457 B.n318 VSUBS 0.007742f
C458 B.n319 VSUBS 0.007742f
C459 B.t8 VSUBS 0.688372f
C460 B.t7 VSUBS 0.697306f
C461 B.t6 VSUBS 0.522019f
C462 B.n320 VSUBS 0.198128f
C463 B.n321 VSUBS 0.07085f
C464 B.n322 VSUBS 0.017936f
C465 B.n323 VSUBS 0.006262f
C466 B.n324 VSUBS 0.007742f
C467 B.n325 VSUBS 0.007742f
C468 B.n326 VSUBS 0.007742f
C469 B.n327 VSUBS 0.007742f
C470 B.n328 VSUBS 0.007742f
C471 B.n329 VSUBS 0.007742f
C472 B.n330 VSUBS 0.007742f
C473 B.n331 VSUBS 0.007742f
C474 B.n332 VSUBS 0.007742f
C475 B.n333 VSUBS 0.007742f
C476 B.n334 VSUBS 0.007742f
C477 B.n335 VSUBS 0.007742f
C478 B.n336 VSUBS 0.007742f
C479 B.n337 VSUBS 0.007742f
C480 B.n338 VSUBS 0.007742f
C481 B.n339 VSUBS 0.007742f
C482 B.n340 VSUBS 0.007742f
C483 B.n341 VSUBS 0.007742f
C484 B.n342 VSUBS 0.007742f
C485 B.n343 VSUBS 0.007742f
C486 B.n344 VSUBS 0.007742f
C487 B.n345 VSUBS 0.007742f
C488 B.n346 VSUBS 0.007742f
C489 B.n347 VSUBS 0.007742f
C490 B.n348 VSUBS 0.007742f
C491 B.n349 VSUBS 0.007742f
C492 B.n350 VSUBS 0.007742f
C493 B.n351 VSUBS 0.007742f
C494 B.n352 VSUBS 0.007742f
C495 B.n353 VSUBS 0.007742f
C496 B.n354 VSUBS 0.007742f
C497 B.n355 VSUBS 0.007742f
C498 B.n356 VSUBS 0.007742f
C499 B.n357 VSUBS 0.007742f
C500 B.n358 VSUBS 0.007742f
C501 B.n359 VSUBS 0.007742f
C502 B.n360 VSUBS 0.007742f
C503 B.n361 VSUBS 0.007742f
C504 B.n362 VSUBS 0.007742f
C505 B.n363 VSUBS 0.007742f
C506 B.n364 VSUBS 0.007742f
C507 B.n365 VSUBS 0.007742f
C508 B.n366 VSUBS 0.007742f
C509 B.n367 VSUBS 0.007742f
C510 B.n368 VSUBS 0.007742f
C511 B.n369 VSUBS 0.007742f
C512 B.n370 VSUBS 0.007742f
C513 B.n371 VSUBS 0.007742f
C514 B.n372 VSUBS 0.007742f
C515 B.n373 VSUBS 0.007742f
C516 B.n374 VSUBS 0.007742f
C517 B.n375 VSUBS 0.007742f
C518 B.n376 VSUBS 0.007742f
C519 B.n377 VSUBS 0.007742f
C520 B.n378 VSUBS 0.007742f
C521 B.n379 VSUBS 0.007742f
C522 B.n380 VSUBS 0.007742f
C523 B.n381 VSUBS 0.007742f
C524 B.n382 VSUBS 0.007742f
C525 B.n383 VSUBS 0.007742f
C526 B.n384 VSUBS 0.007742f
C527 B.n385 VSUBS 0.007742f
C528 B.n386 VSUBS 0.007742f
C529 B.n387 VSUBS 0.007742f
C530 B.n388 VSUBS 0.007742f
C531 B.n389 VSUBS 0.007742f
C532 B.n390 VSUBS 0.007742f
C533 B.n391 VSUBS 0.007742f
C534 B.n392 VSUBS 0.007742f
C535 B.n393 VSUBS 0.007742f
C536 B.n394 VSUBS 0.007742f
C537 B.n395 VSUBS 0.007742f
C538 B.n396 VSUBS 0.007742f
C539 B.n397 VSUBS 0.007742f
C540 B.n398 VSUBS 0.007742f
C541 B.n399 VSUBS 0.007742f
C542 B.n400 VSUBS 0.007742f
C543 B.n401 VSUBS 0.007742f
C544 B.n402 VSUBS 0.007742f
C545 B.n403 VSUBS 0.007742f
C546 B.n404 VSUBS 0.007742f
C547 B.n405 VSUBS 0.007742f
C548 B.n406 VSUBS 0.007742f
C549 B.n407 VSUBS 0.007742f
C550 B.n408 VSUBS 0.007742f
C551 B.n409 VSUBS 0.007742f
C552 B.n410 VSUBS 0.007742f
C553 B.n411 VSUBS 0.007742f
C554 B.n412 VSUBS 0.007742f
C555 B.n413 VSUBS 0.007742f
C556 B.n414 VSUBS 0.007742f
C557 B.n415 VSUBS 0.017221f
C558 B.n416 VSUBS 0.016022f
C559 B.n417 VSUBS 0.017068f
C560 B.n418 VSUBS 0.007742f
C561 B.n419 VSUBS 0.007742f
C562 B.n420 VSUBS 0.007742f
C563 B.n421 VSUBS 0.007742f
C564 B.n422 VSUBS 0.007742f
C565 B.n423 VSUBS 0.007742f
C566 B.n424 VSUBS 0.007742f
C567 B.n425 VSUBS 0.007742f
C568 B.n426 VSUBS 0.007742f
C569 B.n427 VSUBS 0.007742f
C570 B.n428 VSUBS 0.007742f
C571 B.n429 VSUBS 0.007742f
C572 B.n430 VSUBS 0.007742f
C573 B.n431 VSUBS 0.007742f
C574 B.n432 VSUBS 0.007742f
C575 B.n433 VSUBS 0.007742f
C576 B.n434 VSUBS 0.007742f
C577 B.n435 VSUBS 0.007742f
C578 B.n436 VSUBS 0.007742f
C579 B.n437 VSUBS 0.007742f
C580 B.n438 VSUBS 0.007742f
C581 B.n439 VSUBS 0.007742f
C582 B.n440 VSUBS 0.007742f
C583 B.n441 VSUBS 0.007742f
C584 B.n442 VSUBS 0.007742f
C585 B.n443 VSUBS 0.007742f
C586 B.n444 VSUBS 0.007742f
C587 B.n445 VSUBS 0.007742f
C588 B.n446 VSUBS 0.007742f
C589 B.n447 VSUBS 0.007742f
C590 B.n448 VSUBS 0.007742f
C591 B.n449 VSUBS 0.007742f
C592 B.n450 VSUBS 0.007742f
C593 B.n451 VSUBS 0.007742f
C594 B.n452 VSUBS 0.007742f
C595 B.n453 VSUBS 0.007742f
C596 B.n454 VSUBS 0.007742f
C597 B.n455 VSUBS 0.007742f
C598 B.n456 VSUBS 0.007742f
C599 B.n457 VSUBS 0.007742f
C600 B.n458 VSUBS 0.007742f
C601 B.n459 VSUBS 0.007742f
C602 B.n460 VSUBS 0.007742f
C603 B.n461 VSUBS 0.007742f
C604 B.n462 VSUBS 0.007742f
C605 B.n463 VSUBS 0.007742f
C606 B.n464 VSUBS 0.007742f
C607 B.n465 VSUBS 0.007742f
C608 B.n466 VSUBS 0.007742f
C609 B.n467 VSUBS 0.007742f
C610 B.n468 VSUBS 0.007742f
C611 B.n469 VSUBS 0.007742f
C612 B.n470 VSUBS 0.007742f
C613 B.n471 VSUBS 0.007742f
C614 B.n472 VSUBS 0.007742f
C615 B.n473 VSUBS 0.007742f
C616 B.n474 VSUBS 0.007742f
C617 B.n475 VSUBS 0.007742f
C618 B.n476 VSUBS 0.007742f
C619 B.n477 VSUBS 0.007742f
C620 B.n478 VSUBS 0.007742f
C621 B.n479 VSUBS 0.007742f
C622 B.n480 VSUBS 0.007742f
C623 B.n481 VSUBS 0.007742f
C624 B.n482 VSUBS 0.007742f
C625 B.n483 VSUBS 0.007742f
C626 B.n484 VSUBS 0.016022f
C627 B.n485 VSUBS 0.017221f
C628 B.n486 VSUBS 0.017221f
C629 B.n487 VSUBS 0.007742f
C630 B.n488 VSUBS 0.007742f
C631 B.n489 VSUBS 0.007742f
C632 B.n490 VSUBS 0.007742f
C633 B.n491 VSUBS 0.007742f
C634 B.n492 VSUBS 0.007742f
C635 B.n493 VSUBS 0.007742f
C636 B.n494 VSUBS 0.007742f
C637 B.n495 VSUBS 0.007742f
C638 B.n496 VSUBS 0.007742f
C639 B.n497 VSUBS 0.007742f
C640 B.n498 VSUBS 0.007742f
C641 B.n499 VSUBS 0.007742f
C642 B.n500 VSUBS 0.007742f
C643 B.n501 VSUBS 0.007742f
C644 B.n502 VSUBS 0.007742f
C645 B.n503 VSUBS 0.007742f
C646 B.n504 VSUBS 0.007742f
C647 B.n505 VSUBS 0.007742f
C648 B.n506 VSUBS 0.007742f
C649 B.n507 VSUBS 0.007742f
C650 B.n508 VSUBS 0.007742f
C651 B.n509 VSUBS 0.007742f
C652 B.n510 VSUBS 0.007742f
C653 B.n511 VSUBS 0.007742f
C654 B.n512 VSUBS 0.007742f
C655 B.n513 VSUBS 0.007742f
C656 B.n514 VSUBS 0.007742f
C657 B.n515 VSUBS 0.007742f
C658 B.n516 VSUBS 0.007742f
C659 B.n517 VSUBS 0.007742f
C660 B.n518 VSUBS 0.007742f
C661 B.n519 VSUBS 0.007742f
C662 B.n520 VSUBS 0.007742f
C663 B.n521 VSUBS 0.007742f
C664 B.n522 VSUBS 0.007742f
C665 B.n523 VSUBS 0.007742f
C666 B.n524 VSUBS 0.007742f
C667 B.n525 VSUBS 0.007742f
C668 B.n526 VSUBS 0.007742f
C669 B.n527 VSUBS 0.007742f
C670 B.n528 VSUBS 0.007742f
C671 B.n529 VSUBS 0.007742f
C672 B.n530 VSUBS 0.007742f
C673 B.n531 VSUBS 0.007742f
C674 B.n532 VSUBS 0.007742f
C675 B.n533 VSUBS 0.007742f
C676 B.n534 VSUBS 0.007742f
C677 B.n535 VSUBS 0.007742f
C678 B.n536 VSUBS 0.007742f
C679 B.n537 VSUBS 0.007742f
C680 B.n538 VSUBS 0.007742f
C681 B.n539 VSUBS 0.007742f
C682 B.n540 VSUBS 0.007742f
C683 B.n541 VSUBS 0.007742f
C684 B.n542 VSUBS 0.007742f
C685 B.n543 VSUBS 0.007742f
C686 B.n544 VSUBS 0.007742f
C687 B.n545 VSUBS 0.007742f
C688 B.n546 VSUBS 0.007742f
C689 B.n547 VSUBS 0.007742f
C690 B.n548 VSUBS 0.007742f
C691 B.n549 VSUBS 0.007742f
C692 B.n550 VSUBS 0.007742f
C693 B.n551 VSUBS 0.007742f
C694 B.n552 VSUBS 0.007742f
C695 B.n553 VSUBS 0.007742f
C696 B.n554 VSUBS 0.007742f
C697 B.n555 VSUBS 0.007742f
C698 B.n556 VSUBS 0.007742f
C699 B.n557 VSUBS 0.007742f
C700 B.n558 VSUBS 0.007742f
C701 B.n559 VSUBS 0.007742f
C702 B.n560 VSUBS 0.007742f
C703 B.n561 VSUBS 0.007742f
C704 B.n562 VSUBS 0.007742f
C705 B.n563 VSUBS 0.007742f
C706 B.n564 VSUBS 0.007742f
C707 B.n565 VSUBS 0.007742f
C708 B.n566 VSUBS 0.007742f
C709 B.n567 VSUBS 0.007742f
C710 B.n568 VSUBS 0.007742f
C711 B.n569 VSUBS 0.007742f
C712 B.n570 VSUBS 0.007742f
C713 B.n571 VSUBS 0.007742f
C714 B.n572 VSUBS 0.007742f
C715 B.n573 VSUBS 0.007742f
C716 B.n574 VSUBS 0.007742f
C717 B.n575 VSUBS 0.005351f
C718 B.n576 VSUBS 0.007742f
C719 B.n577 VSUBS 0.007742f
C720 B.n578 VSUBS 0.006262f
C721 B.n579 VSUBS 0.007742f
C722 B.n580 VSUBS 0.007742f
C723 B.n581 VSUBS 0.007742f
C724 B.n582 VSUBS 0.007742f
C725 B.n583 VSUBS 0.007742f
C726 B.n584 VSUBS 0.007742f
C727 B.n585 VSUBS 0.007742f
C728 B.n586 VSUBS 0.007742f
C729 B.n587 VSUBS 0.007742f
C730 B.n588 VSUBS 0.007742f
C731 B.n589 VSUBS 0.007742f
C732 B.n590 VSUBS 0.006262f
C733 B.n591 VSUBS 0.017936f
C734 B.n592 VSUBS 0.005351f
C735 B.n593 VSUBS 0.007742f
C736 B.n594 VSUBS 0.007742f
C737 B.n595 VSUBS 0.007742f
C738 B.n596 VSUBS 0.007742f
C739 B.n597 VSUBS 0.007742f
C740 B.n598 VSUBS 0.007742f
C741 B.n599 VSUBS 0.007742f
C742 B.n600 VSUBS 0.007742f
C743 B.n601 VSUBS 0.007742f
C744 B.n602 VSUBS 0.007742f
C745 B.n603 VSUBS 0.007742f
C746 B.n604 VSUBS 0.007742f
C747 B.n605 VSUBS 0.007742f
C748 B.n606 VSUBS 0.007742f
C749 B.n607 VSUBS 0.007742f
C750 B.n608 VSUBS 0.007742f
C751 B.n609 VSUBS 0.007742f
C752 B.n610 VSUBS 0.007742f
C753 B.n611 VSUBS 0.007742f
C754 B.n612 VSUBS 0.007742f
C755 B.n613 VSUBS 0.007742f
C756 B.n614 VSUBS 0.007742f
C757 B.n615 VSUBS 0.007742f
C758 B.n616 VSUBS 0.007742f
C759 B.n617 VSUBS 0.007742f
C760 B.n618 VSUBS 0.007742f
C761 B.n619 VSUBS 0.007742f
C762 B.n620 VSUBS 0.007742f
C763 B.n621 VSUBS 0.007742f
C764 B.n622 VSUBS 0.007742f
C765 B.n623 VSUBS 0.007742f
C766 B.n624 VSUBS 0.007742f
C767 B.n625 VSUBS 0.007742f
C768 B.n626 VSUBS 0.007742f
C769 B.n627 VSUBS 0.007742f
C770 B.n628 VSUBS 0.007742f
C771 B.n629 VSUBS 0.007742f
C772 B.n630 VSUBS 0.007742f
C773 B.n631 VSUBS 0.007742f
C774 B.n632 VSUBS 0.007742f
C775 B.n633 VSUBS 0.007742f
C776 B.n634 VSUBS 0.007742f
C777 B.n635 VSUBS 0.007742f
C778 B.n636 VSUBS 0.007742f
C779 B.n637 VSUBS 0.007742f
C780 B.n638 VSUBS 0.007742f
C781 B.n639 VSUBS 0.007742f
C782 B.n640 VSUBS 0.007742f
C783 B.n641 VSUBS 0.007742f
C784 B.n642 VSUBS 0.007742f
C785 B.n643 VSUBS 0.007742f
C786 B.n644 VSUBS 0.007742f
C787 B.n645 VSUBS 0.007742f
C788 B.n646 VSUBS 0.007742f
C789 B.n647 VSUBS 0.007742f
C790 B.n648 VSUBS 0.007742f
C791 B.n649 VSUBS 0.007742f
C792 B.n650 VSUBS 0.007742f
C793 B.n651 VSUBS 0.007742f
C794 B.n652 VSUBS 0.007742f
C795 B.n653 VSUBS 0.007742f
C796 B.n654 VSUBS 0.007742f
C797 B.n655 VSUBS 0.007742f
C798 B.n656 VSUBS 0.007742f
C799 B.n657 VSUBS 0.007742f
C800 B.n658 VSUBS 0.007742f
C801 B.n659 VSUBS 0.007742f
C802 B.n660 VSUBS 0.007742f
C803 B.n661 VSUBS 0.007742f
C804 B.n662 VSUBS 0.007742f
C805 B.n663 VSUBS 0.007742f
C806 B.n664 VSUBS 0.007742f
C807 B.n665 VSUBS 0.007742f
C808 B.n666 VSUBS 0.007742f
C809 B.n667 VSUBS 0.007742f
C810 B.n668 VSUBS 0.007742f
C811 B.n669 VSUBS 0.007742f
C812 B.n670 VSUBS 0.007742f
C813 B.n671 VSUBS 0.007742f
C814 B.n672 VSUBS 0.007742f
C815 B.n673 VSUBS 0.007742f
C816 B.n674 VSUBS 0.007742f
C817 B.n675 VSUBS 0.007742f
C818 B.n676 VSUBS 0.007742f
C819 B.n677 VSUBS 0.007742f
C820 B.n678 VSUBS 0.007742f
C821 B.n679 VSUBS 0.007742f
C822 B.n680 VSUBS 0.007742f
C823 B.n681 VSUBS 0.007742f
C824 B.n682 VSUBS 0.017221f
C825 B.n683 VSUBS 0.016022f
C826 B.n684 VSUBS 0.016022f
C827 B.n685 VSUBS 0.007742f
C828 B.n686 VSUBS 0.007742f
C829 B.n687 VSUBS 0.007742f
C830 B.n688 VSUBS 0.007742f
C831 B.n689 VSUBS 0.007742f
C832 B.n690 VSUBS 0.007742f
C833 B.n691 VSUBS 0.007742f
C834 B.n692 VSUBS 0.007742f
C835 B.n693 VSUBS 0.007742f
C836 B.n694 VSUBS 0.007742f
C837 B.n695 VSUBS 0.007742f
C838 B.n696 VSUBS 0.007742f
C839 B.n697 VSUBS 0.007742f
C840 B.n698 VSUBS 0.007742f
C841 B.n699 VSUBS 0.007742f
C842 B.n700 VSUBS 0.007742f
C843 B.n701 VSUBS 0.007742f
C844 B.n702 VSUBS 0.007742f
C845 B.n703 VSUBS 0.007742f
C846 B.n704 VSUBS 0.007742f
C847 B.n705 VSUBS 0.007742f
C848 B.n706 VSUBS 0.007742f
C849 B.n707 VSUBS 0.007742f
C850 B.n708 VSUBS 0.007742f
C851 B.n709 VSUBS 0.007742f
C852 B.n710 VSUBS 0.007742f
C853 B.n711 VSUBS 0.007742f
C854 B.n712 VSUBS 0.007742f
C855 B.n713 VSUBS 0.007742f
C856 B.n714 VSUBS 0.007742f
C857 B.n715 VSUBS 0.010102f
C858 B.n716 VSUBS 0.010762f
C859 B.n717 VSUBS 0.021401f
.ends

