* NGSPICE file created from diff_pair_sample_1685.ext - technology: sky130A

.subckt diff_pair_sample_1685 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X1 VTAIL.t16 VN.t1 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X2 VDD2.t2 VN.t2 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X3 VDD1.t9 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X4 VDD2.t8 VN.t3 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=2.27
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=2.27
X6 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=2.27
X7 VDD1.t8 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=2.27
X8 VTAIL.t5 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=2.27
X10 VDD1.t6 VP.t3 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=2.27
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=0 ps=0 w=7.85 l=2.27
X12 VTAIL.t18 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X13 VTAIL.t13 VN.t4 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X14 VDD2.t6 VN.t5 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=2.27
X15 VDD1.t4 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=3.0615 ps=16.48 w=7.85 l=2.27
X16 VTAIL.t1 VP.t6 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X17 VDD2.t1 VN.t6 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X18 VDD2.t9 VN.t7 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=2.27
X19 VDD2.t3 VN.t8 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=2.27
X20 VDD1.t2 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0615 pd=16.48 as=1.29525 ps=8.18 w=7.85 l=2.27
X21 VDD1.t1 VP.t8 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X22 VTAIL.t4 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
X23 VTAIL.t8 VN.t9 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.29525 pd=8.18 as=1.29525 ps=8.18 w=7.85 l=2.27
R0 VN.n71 VN.n37 161.3
R1 VN.n70 VN.n69 161.3
R2 VN.n68 VN.n38 161.3
R3 VN.n67 VN.n66 161.3
R4 VN.n65 VN.n39 161.3
R5 VN.n63 VN.n62 161.3
R6 VN.n61 VN.n40 161.3
R7 VN.n60 VN.n59 161.3
R8 VN.n58 VN.n41 161.3
R9 VN.n57 VN.n56 161.3
R10 VN.n55 VN.n42 161.3
R11 VN.n54 VN.n53 161.3
R12 VN.n52 VN.n43 161.3
R13 VN.n51 VN.n50 161.3
R14 VN.n49 VN.n44 161.3
R15 VN.n48 VN.n47 161.3
R16 VN.n34 VN.n0 161.3
R17 VN.n33 VN.n32 161.3
R18 VN.n31 VN.n1 161.3
R19 VN.n30 VN.n29 161.3
R20 VN.n28 VN.n2 161.3
R21 VN.n26 VN.n25 161.3
R22 VN.n24 VN.n3 161.3
R23 VN.n23 VN.n22 161.3
R24 VN.n21 VN.n4 161.3
R25 VN.n20 VN.n19 161.3
R26 VN.n18 VN.n5 161.3
R27 VN.n17 VN.n16 161.3
R28 VN.n15 VN.n6 161.3
R29 VN.n14 VN.n13 161.3
R30 VN.n12 VN.n7 161.3
R31 VN.n11 VN.n10 161.3
R32 VN.n8 VN.t8 114.216
R33 VN.n45 VN.t5 114.216
R34 VN.n36 VN.n35 100.969
R35 VN.n73 VN.n72 100.969
R36 VN.n5 VN.t2 83.3419
R37 VN.n9 VN.t1 83.3419
R38 VN.n27 VN.t0 83.3419
R39 VN.n35 VN.t3 83.3419
R40 VN.n42 VN.t6 83.3419
R41 VN.n46 VN.t4 83.3419
R42 VN.n64 VN.t9 83.3419
R43 VN.n72 VN.t7 83.3419
R44 VN.n9 VN.n8 67.1934
R45 VN.n46 VN.n45 67.1934
R46 VN.n15 VN.n14 56.5193
R47 VN.n22 VN.n21 56.5193
R48 VN.n52 VN.n51 56.5193
R49 VN.n59 VN.n58 56.5193
R50 VN.n29 VN.n1 50.2061
R51 VN.n66 VN.n38 50.2061
R52 VN VN.n73 48.3921
R53 VN.n33 VN.n1 30.7807
R54 VN.n70 VN.n38 30.7807
R55 VN.n10 VN.n7 24.4675
R56 VN.n14 VN.n7 24.4675
R57 VN.n16 VN.n15 24.4675
R58 VN.n16 VN.n5 24.4675
R59 VN.n20 VN.n5 24.4675
R60 VN.n21 VN.n20 24.4675
R61 VN.n22 VN.n3 24.4675
R62 VN.n26 VN.n3 24.4675
R63 VN.n29 VN.n28 24.4675
R64 VN.n34 VN.n33 24.4675
R65 VN.n51 VN.n44 24.4675
R66 VN.n47 VN.n44 24.4675
R67 VN.n58 VN.n57 24.4675
R68 VN.n57 VN.n42 24.4675
R69 VN.n53 VN.n42 24.4675
R70 VN.n53 VN.n52 24.4675
R71 VN.n66 VN.n65 24.4675
R72 VN.n63 VN.n40 24.4675
R73 VN.n59 VN.n40 24.4675
R74 VN.n71 VN.n70 24.4675
R75 VN.n28 VN.n27 19.5741
R76 VN.n65 VN.n64 19.5741
R77 VN.n48 VN.n45 10.026
R78 VN.n11 VN.n8 10.026
R79 VN.n35 VN.n34 9.7873
R80 VN.n72 VN.n71 9.7873
R81 VN.n10 VN.n9 4.8939
R82 VN.n27 VN.n26 4.8939
R83 VN.n47 VN.n46 4.8939
R84 VN.n64 VN.n63 4.8939
R85 VN.n73 VN.n37 0.278367
R86 VN.n36 VN.n0 0.278367
R87 VN.n69 VN.n37 0.189894
R88 VN.n69 VN.n68 0.189894
R89 VN.n68 VN.n67 0.189894
R90 VN.n67 VN.n39 0.189894
R91 VN.n62 VN.n39 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n60 0.189894
R94 VN.n60 VN.n41 0.189894
R95 VN.n56 VN.n41 0.189894
R96 VN.n56 VN.n55 0.189894
R97 VN.n55 VN.n54 0.189894
R98 VN.n54 VN.n43 0.189894
R99 VN.n50 VN.n43 0.189894
R100 VN.n50 VN.n49 0.189894
R101 VN.n49 VN.n48 0.189894
R102 VN.n12 VN.n11 0.189894
R103 VN.n13 VN.n12 0.189894
R104 VN.n13 VN.n6 0.189894
R105 VN.n17 VN.n6 0.189894
R106 VN.n18 VN.n17 0.189894
R107 VN.n19 VN.n18 0.189894
R108 VN.n19 VN.n4 0.189894
R109 VN.n23 VN.n4 0.189894
R110 VN.n24 VN.n23 0.189894
R111 VN.n25 VN.n24 0.189894
R112 VN.n25 VN.n2 0.189894
R113 VN.n30 VN.n2 0.189894
R114 VN.n31 VN.n30 0.189894
R115 VN.n32 VN.n31 0.189894
R116 VN.n32 VN.n0 0.189894
R117 VN VN.n36 0.153454
R118 VDD2.n81 VDD2.n45 289.615
R119 VDD2.n36 VDD2.n0 289.615
R120 VDD2.n82 VDD2.n81 185
R121 VDD2.n80 VDD2.n47 185
R122 VDD2.n79 VDD2.n78 185
R123 VDD2.n50 VDD2.n48 185
R124 VDD2.n73 VDD2.n72 185
R125 VDD2.n71 VDD2.n70 185
R126 VDD2.n54 VDD2.n53 185
R127 VDD2.n65 VDD2.n64 185
R128 VDD2.n63 VDD2.n62 185
R129 VDD2.n58 VDD2.n57 185
R130 VDD2.n12 VDD2.n11 185
R131 VDD2.n17 VDD2.n16 185
R132 VDD2.n19 VDD2.n18 185
R133 VDD2.n8 VDD2.n7 185
R134 VDD2.n25 VDD2.n24 185
R135 VDD2.n27 VDD2.n26 185
R136 VDD2.n4 VDD2.n3 185
R137 VDD2.n34 VDD2.n33 185
R138 VDD2.n35 VDD2.n2 185
R139 VDD2.n37 VDD2.n36 185
R140 VDD2.n59 VDD2.t9 149.524
R141 VDD2.n13 VDD2.t3 149.524
R142 VDD2.n81 VDD2.n80 104.615
R143 VDD2.n80 VDD2.n79 104.615
R144 VDD2.n79 VDD2.n48 104.615
R145 VDD2.n72 VDD2.n48 104.615
R146 VDD2.n72 VDD2.n71 104.615
R147 VDD2.n71 VDD2.n53 104.615
R148 VDD2.n64 VDD2.n53 104.615
R149 VDD2.n64 VDD2.n63 104.615
R150 VDD2.n63 VDD2.n57 104.615
R151 VDD2.n17 VDD2.n11 104.615
R152 VDD2.n18 VDD2.n17 104.615
R153 VDD2.n18 VDD2.n7 104.615
R154 VDD2.n25 VDD2.n7 104.615
R155 VDD2.n26 VDD2.n25 104.615
R156 VDD2.n26 VDD2.n3 104.615
R157 VDD2.n34 VDD2.n3 104.615
R158 VDD2.n35 VDD2.n34 104.615
R159 VDD2.n36 VDD2.n35 104.615
R160 VDD2.n44 VDD2.n43 66.5732
R161 VDD2 VDD2.n89 66.5703
R162 VDD2.n88 VDD2.n87 64.9477
R163 VDD2.n42 VDD2.n41 64.9475
R164 VDD2.t9 VDD2.n57 52.3082
R165 VDD2.t3 VDD2.n11 52.3082
R166 VDD2.n42 VDD2.n40 52.0752
R167 VDD2.n86 VDD2.n85 49.8338
R168 VDD2.n86 VDD2.n44 41.1291
R169 VDD2.n82 VDD2.n47 13.1884
R170 VDD2.n37 VDD2.n2 13.1884
R171 VDD2.n83 VDD2.n45 12.8005
R172 VDD2.n78 VDD2.n49 12.8005
R173 VDD2.n33 VDD2.n32 12.8005
R174 VDD2.n38 VDD2.n0 12.8005
R175 VDD2.n77 VDD2.n50 12.0247
R176 VDD2.n31 VDD2.n4 12.0247
R177 VDD2.n74 VDD2.n73 11.249
R178 VDD2.n28 VDD2.n27 11.249
R179 VDD2.n70 VDD2.n52 10.4732
R180 VDD2.n24 VDD2.n6 10.4732
R181 VDD2.n59 VDD2.n58 10.2747
R182 VDD2.n13 VDD2.n12 10.2747
R183 VDD2.n69 VDD2.n54 9.69747
R184 VDD2.n23 VDD2.n8 9.69747
R185 VDD2.n85 VDD2.n84 9.45567
R186 VDD2.n40 VDD2.n39 9.45567
R187 VDD2.n61 VDD2.n60 9.3005
R188 VDD2.n56 VDD2.n55 9.3005
R189 VDD2.n67 VDD2.n66 9.3005
R190 VDD2.n69 VDD2.n68 9.3005
R191 VDD2.n52 VDD2.n51 9.3005
R192 VDD2.n75 VDD2.n74 9.3005
R193 VDD2.n77 VDD2.n76 9.3005
R194 VDD2.n49 VDD2.n46 9.3005
R195 VDD2.n84 VDD2.n83 9.3005
R196 VDD2.n39 VDD2.n38 9.3005
R197 VDD2.n15 VDD2.n14 9.3005
R198 VDD2.n10 VDD2.n9 9.3005
R199 VDD2.n21 VDD2.n20 9.3005
R200 VDD2.n23 VDD2.n22 9.3005
R201 VDD2.n6 VDD2.n5 9.3005
R202 VDD2.n29 VDD2.n28 9.3005
R203 VDD2.n31 VDD2.n30 9.3005
R204 VDD2.n32 VDD2.n1 9.3005
R205 VDD2.n66 VDD2.n65 8.92171
R206 VDD2.n20 VDD2.n19 8.92171
R207 VDD2.n62 VDD2.n56 8.14595
R208 VDD2.n16 VDD2.n10 8.14595
R209 VDD2.n61 VDD2.n58 7.3702
R210 VDD2.n15 VDD2.n12 7.3702
R211 VDD2.n62 VDD2.n61 5.81868
R212 VDD2.n16 VDD2.n15 5.81868
R213 VDD2.n65 VDD2.n56 5.04292
R214 VDD2.n19 VDD2.n10 5.04292
R215 VDD2.n66 VDD2.n54 4.26717
R216 VDD2.n20 VDD2.n8 4.26717
R217 VDD2.n70 VDD2.n69 3.49141
R218 VDD2.n24 VDD2.n23 3.49141
R219 VDD2.n60 VDD2.n59 2.84304
R220 VDD2.n14 VDD2.n13 2.84304
R221 VDD2.n73 VDD2.n52 2.71565
R222 VDD2.n27 VDD2.n6 2.71565
R223 VDD2.n89 VDD2.t7 2.52279
R224 VDD2.n89 VDD2.t6 2.52279
R225 VDD2.n87 VDD2.t4 2.52279
R226 VDD2.n87 VDD2.t1 2.52279
R227 VDD2.n43 VDD2.t0 2.52279
R228 VDD2.n43 VDD2.t8 2.52279
R229 VDD2.n41 VDD2.t5 2.52279
R230 VDD2.n41 VDD2.t2 2.52279
R231 VDD2.n88 VDD2.n86 2.24188
R232 VDD2.n74 VDD2.n50 1.93989
R233 VDD2.n28 VDD2.n4 1.93989
R234 VDD2.n85 VDD2.n45 1.16414
R235 VDD2.n78 VDD2.n77 1.16414
R236 VDD2.n33 VDD2.n31 1.16414
R237 VDD2.n40 VDD2.n0 1.16414
R238 VDD2 VDD2.n88 0.619035
R239 VDD2.n44 VDD2.n42 0.505499
R240 VDD2.n83 VDD2.n82 0.388379
R241 VDD2.n49 VDD2.n47 0.388379
R242 VDD2.n32 VDD2.n2 0.388379
R243 VDD2.n38 VDD2.n37 0.388379
R244 VDD2.n84 VDD2.n46 0.155672
R245 VDD2.n76 VDD2.n46 0.155672
R246 VDD2.n76 VDD2.n75 0.155672
R247 VDD2.n75 VDD2.n51 0.155672
R248 VDD2.n68 VDD2.n51 0.155672
R249 VDD2.n68 VDD2.n67 0.155672
R250 VDD2.n67 VDD2.n55 0.155672
R251 VDD2.n60 VDD2.n55 0.155672
R252 VDD2.n14 VDD2.n9 0.155672
R253 VDD2.n21 VDD2.n9 0.155672
R254 VDD2.n22 VDD2.n21 0.155672
R255 VDD2.n22 VDD2.n5 0.155672
R256 VDD2.n29 VDD2.n5 0.155672
R257 VDD2.n30 VDD2.n29 0.155672
R258 VDD2.n30 VDD2.n1 0.155672
R259 VDD2.n39 VDD2.n1 0.155672
R260 VTAIL.n176 VTAIL.n140 289.615
R261 VTAIL.n38 VTAIL.n2 289.615
R262 VTAIL.n134 VTAIL.n98 289.615
R263 VTAIL.n88 VTAIL.n52 289.615
R264 VTAIL.n152 VTAIL.n151 185
R265 VTAIL.n157 VTAIL.n156 185
R266 VTAIL.n159 VTAIL.n158 185
R267 VTAIL.n148 VTAIL.n147 185
R268 VTAIL.n165 VTAIL.n164 185
R269 VTAIL.n167 VTAIL.n166 185
R270 VTAIL.n144 VTAIL.n143 185
R271 VTAIL.n174 VTAIL.n173 185
R272 VTAIL.n175 VTAIL.n142 185
R273 VTAIL.n177 VTAIL.n176 185
R274 VTAIL.n14 VTAIL.n13 185
R275 VTAIL.n19 VTAIL.n18 185
R276 VTAIL.n21 VTAIL.n20 185
R277 VTAIL.n10 VTAIL.n9 185
R278 VTAIL.n27 VTAIL.n26 185
R279 VTAIL.n29 VTAIL.n28 185
R280 VTAIL.n6 VTAIL.n5 185
R281 VTAIL.n36 VTAIL.n35 185
R282 VTAIL.n37 VTAIL.n4 185
R283 VTAIL.n39 VTAIL.n38 185
R284 VTAIL.n135 VTAIL.n134 185
R285 VTAIL.n133 VTAIL.n100 185
R286 VTAIL.n132 VTAIL.n131 185
R287 VTAIL.n103 VTAIL.n101 185
R288 VTAIL.n126 VTAIL.n125 185
R289 VTAIL.n124 VTAIL.n123 185
R290 VTAIL.n107 VTAIL.n106 185
R291 VTAIL.n118 VTAIL.n117 185
R292 VTAIL.n116 VTAIL.n115 185
R293 VTAIL.n111 VTAIL.n110 185
R294 VTAIL.n89 VTAIL.n88 185
R295 VTAIL.n87 VTAIL.n54 185
R296 VTAIL.n86 VTAIL.n85 185
R297 VTAIL.n57 VTAIL.n55 185
R298 VTAIL.n80 VTAIL.n79 185
R299 VTAIL.n78 VTAIL.n77 185
R300 VTAIL.n61 VTAIL.n60 185
R301 VTAIL.n72 VTAIL.n71 185
R302 VTAIL.n70 VTAIL.n69 185
R303 VTAIL.n65 VTAIL.n64 185
R304 VTAIL.n153 VTAIL.t14 149.524
R305 VTAIL.n15 VTAIL.t7 149.524
R306 VTAIL.n112 VTAIL.t3 149.524
R307 VTAIL.n66 VTAIL.t12 149.524
R308 VTAIL.n157 VTAIL.n151 104.615
R309 VTAIL.n158 VTAIL.n157 104.615
R310 VTAIL.n158 VTAIL.n147 104.615
R311 VTAIL.n165 VTAIL.n147 104.615
R312 VTAIL.n166 VTAIL.n165 104.615
R313 VTAIL.n166 VTAIL.n143 104.615
R314 VTAIL.n174 VTAIL.n143 104.615
R315 VTAIL.n175 VTAIL.n174 104.615
R316 VTAIL.n176 VTAIL.n175 104.615
R317 VTAIL.n19 VTAIL.n13 104.615
R318 VTAIL.n20 VTAIL.n19 104.615
R319 VTAIL.n20 VTAIL.n9 104.615
R320 VTAIL.n27 VTAIL.n9 104.615
R321 VTAIL.n28 VTAIL.n27 104.615
R322 VTAIL.n28 VTAIL.n5 104.615
R323 VTAIL.n36 VTAIL.n5 104.615
R324 VTAIL.n37 VTAIL.n36 104.615
R325 VTAIL.n38 VTAIL.n37 104.615
R326 VTAIL.n134 VTAIL.n133 104.615
R327 VTAIL.n133 VTAIL.n132 104.615
R328 VTAIL.n132 VTAIL.n101 104.615
R329 VTAIL.n125 VTAIL.n101 104.615
R330 VTAIL.n125 VTAIL.n124 104.615
R331 VTAIL.n124 VTAIL.n106 104.615
R332 VTAIL.n117 VTAIL.n106 104.615
R333 VTAIL.n117 VTAIL.n116 104.615
R334 VTAIL.n116 VTAIL.n110 104.615
R335 VTAIL.n88 VTAIL.n87 104.615
R336 VTAIL.n87 VTAIL.n86 104.615
R337 VTAIL.n86 VTAIL.n55 104.615
R338 VTAIL.n79 VTAIL.n55 104.615
R339 VTAIL.n79 VTAIL.n78 104.615
R340 VTAIL.n78 VTAIL.n60 104.615
R341 VTAIL.n71 VTAIL.n60 104.615
R342 VTAIL.n71 VTAIL.n70 104.615
R343 VTAIL.n70 VTAIL.n64 104.615
R344 VTAIL.t14 VTAIL.n151 52.3082
R345 VTAIL.t7 VTAIL.n13 52.3082
R346 VTAIL.t3 VTAIL.n110 52.3082
R347 VTAIL.t12 VTAIL.n64 52.3082
R348 VTAIL.n97 VTAIL.n96 48.2689
R349 VTAIL.n95 VTAIL.n94 48.2689
R350 VTAIL.n51 VTAIL.n50 48.2689
R351 VTAIL.n49 VTAIL.n48 48.2689
R352 VTAIL.n183 VTAIL.n182 48.2687
R353 VTAIL.n1 VTAIL.n0 48.2687
R354 VTAIL.n45 VTAIL.n44 48.2687
R355 VTAIL.n47 VTAIL.n46 48.2687
R356 VTAIL.n181 VTAIL.n180 33.155
R357 VTAIL.n43 VTAIL.n42 33.155
R358 VTAIL.n139 VTAIL.n138 33.155
R359 VTAIL.n93 VTAIL.n92 33.155
R360 VTAIL.n49 VTAIL.n47 23.6169
R361 VTAIL.n181 VTAIL.n139 21.3755
R362 VTAIL.n177 VTAIL.n142 13.1884
R363 VTAIL.n39 VTAIL.n4 13.1884
R364 VTAIL.n135 VTAIL.n100 13.1884
R365 VTAIL.n89 VTAIL.n54 13.1884
R366 VTAIL.n173 VTAIL.n172 12.8005
R367 VTAIL.n178 VTAIL.n140 12.8005
R368 VTAIL.n35 VTAIL.n34 12.8005
R369 VTAIL.n40 VTAIL.n2 12.8005
R370 VTAIL.n136 VTAIL.n98 12.8005
R371 VTAIL.n131 VTAIL.n102 12.8005
R372 VTAIL.n90 VTAIL.n52 12.8005
R373 VTAIL.n85 VTAIL.n56 12.8005
R374 VTAIL.n171 VTAIL.n144 12.0247
R375 VTAIL.n33 VTAIL.n6 12.0247
R376 VTAIL.n130 VTAIL.n103 12.0247
R377 VTAIL.n84 VTAIL.n57 12.0247
R378 VTAIL.n168 VTAIL.n167 11.249
R379 VTAIL.n30 VTAIL.n29 11.249
R380 VTAIL.n127 VTAIL.n126 11.249
R381 VTAIL.n81 VTAIL.n80 11.249
R382 VTAIL.n164 VTAIL.n146 10.4732
R383 VTAIL.n26 VTAIL.n8 10.4732
R384 VTAIL.n123 VTAIL.n105 10.4732
R385 VTAIL.n77 VTAIL.n59 10.4732
R386 VTAIL.n153 VTAIL.n152 10.2747
R387 VTAIL.n15 VTAIL.n14 10.2747
R388 VTAIL.n112 VTAIL.n111 10.2747
R389 VTAIL.n66 VTAIL.n65 10.2747
R390 VTAIL.n163 VTAIL.n148 9.69747
R391 VTAIL.n25 VTAIL.n10 9.69747
R392 VTAIL.n122 VTAIL.n107 9.69747
R393 VTAIL.n76 VTAIL.n61 9.69747
R394 VTAIL.n180 VTAIL.n179 9.45567
R395 VTAIL.n42 VTAIL.n41 9.45567
R396 VTAIL.n138 VTAIL.n137 9.45567
R397 VTAIL.n92 VTAIL.n91 9.45567
R398 VTAIL.n179 VTAIL.n178 9.3005
R399 VTAIL.n155 VTAIL.n154 9.3005
R400 VTAIL.n150 VTAIL.n149 9.3005
R401 VTAIL.n161 VTAIL.n160 9.3005
R402 VTAIL.n163 VTAIL.n162 9.3005
R403 VTAIL.n146 VTAIL.n145 9.3005
R404 VTAIL.n169 VTAIL.n168 9.3005
R405 VTAIL.n171 VTAIL.n170 9.3005
R406 VTAIL.n172 VTAIL.n141 9.3005
R407 VTAIL.n41 VTAIL.n40 9.3005
R408 VTAIL.n17 VTAIL.n16 9.3005
R409 VTAIL.n12 VTAIL.n11 9.3005
R410 VTAIL.n23 VTAIL.n22 9.3005
R411 VTAIL.n25 VTAIL.n24 9.3005
R412 VTAIL.n8 VTAIL.n7 9.3005
R413 VTAIL.n31 VTAIL.n30 9.3005
R414 VTAIL.n33 VTAIL.n32 9.3005
R415 VTAIL.n34 VTAIL.n3 9.3005
R416 VTAIL.n114 VTAIL.n113 9.3005
R417 VTAIL.n109 VTAIL.n108 9.3005
R418 VTAIL.n120 VTAIL.n119 9.3005
R419 VTAIL.n122 VTAIL.n121 9.3005
R420 VTAIL.n105 VTAIL.n104 9.3005
R421 VTAIL.n128 VTAIL.n127 9.3005
R422 VTAIL.n130 VTAIL.n129 9.3005
R423 VTAIL.n102 VTAIL.n99 9.3005
R424 VTAIL.n137 VTAIL.n136 9.3005
R425 VTAIL.n68 VTAIL.n67 9.3005
R426 VTAIL.n63 VTAIL.n62 9.3005
R427 VTAIL.n74 VTAIL.n73 9.3005
R428 VTAIL.n76 VTAIL.n75 9.3005
R429 VTAIL.n59 VTAIL.n58 9.3005
R430 VTAIL.n82 VTAIL.n81 9.3005
R431 VTAIL.n84 VTAIL.n83 9.3005
R432 VTAIL.n56 VTAIL.n53 9.3005
R433 VTAIL.n91 VTAIL.n90 9.3005
R434 VTAIL.n160 VTAIL.n159 8.92171
R435 VTAIL.n22 VTAIL.n21 8.92171
R436 VTAIL.n119 VTAIL.n118 8.92171
R437 VTAIL.n73 VTAIL.n72 8.92171
R438 VTAIL.n156 VTAIL.n150 8.14595
R439 VTAIL.n18 VTAIL.n12 8.14595
R440 VTAIL.n115 VTAIL.n109 8.14595
R441 VTAIL.n69 VTAIL.n63 8.14595
R442 VTAIL.n155 VTAIL.n152 7.3702
R443 VTAIL.n17 VTAIL.n14 7.3702
R444 VTAIL.n114 VTAIL.n111 7.3702
R445 VTAIL.n68 VTAIL.n65 7.3702
R446 VTAIL.n156 VTAIL.n155 5.81868
R447 VTAIL.n18 VTAIL.n17 5.81868
R448 VTAIL.n115 VTAIL.n114 5.81868
R449 VTAIL.n69 VTAIL.n68 5.81868
R450 VTAIL.n159 VTAIL.n150 5.04292
R451 VTAIL.n21 VTAIL.n12 5.04292
R452 VTAIL.n118 VTAIL.n109 5.04292
R453 VTAIL.n72 VTAIL.n63 5.04292
R454 VTAIL.n160 VTAIL.n148 4.26717
R455 VTAIL.n22 VTAIL.n10 4.26717
R456 VTAIL.n119 VTAIL.n107 4.26717
R457 VTAIL.n73 VTAIL.n61 4.26717
R458 VTAIL.n164 VTAIL.n163 3.49141
R459 VTAIL.n26 VTAIL.n25 3.49141
R460 VTAIL.n123 VTAIL.n122 3.49141
R461 VTAIL.n77 VTAIL.n76 3.49141
R462 VTAIL.n154 VTAIL.n153 2.84304
R463 VTAIL.n16 VTAIL.n15 2.84304
R464 VTAIL.n113 VTAIL.n112 2.84304
R465 VTAIL.n67 VTAIL.n66 2.84304
R466 VTAIL.n167 VTAIL.n146 2.71565
R467 VTAIL.n29 VTAIL.n8 2.71565
R468 VTAIL.n126 VTAIL.n105 2.71565
R469 VTAIL.n80 VTAIL.n59 2.71565
R470 VTAIL.n182 VTAIL.t15 2.52279
R471 VTAIL.n182 VTAIL.t17 2.52279
R472 VTAIL.n0 VTAIL.t9 2.52279
R473 VTAIL.n0 VTAIL.t16 2.52279
R474 VTAIL.n44 VTAIL.t6 2.52279
R475 VTAIL.n44 VTAIL.t5 2.52279
R476 VTAIL.n46 VTAIL.t19 2.52279
R477 VTAIL.n46 VTAIL.t18 2.52279
R478 VTAIL.n96 VTAIL.t2 2.52279
R479 VTAIL.n96 VTAIL.t1 2.52279
R480 VTAIL.n94 VTAIL.t0 2.52279
R481 VTAIL.n94 VTAIL.t4 2.52279
R482 VTAIL.n50 VTAIL.t11 2.52279
R483 VTAIL.n50 VTAIL.t13 2.52279
R484 VTAIL.n48 VTAIL.t10 2.52279
R485 VTAIL.n48 VTAIL.t8 2.52279
R486 VTAIL.n51 VTAIL.n49 2.24188
R487 VTAIL.n93 VTAIL.n51 2.24188
R488 VTAIL.n97 VTAIL.n95 2.24188
R489 VTAIL.n139 VTAIL.n97 2.24188
R490 VTAIL.n47 VTAIL.n45 2.24188
R491 VTAIL.n45 VTAIL.n43 2.24188
R492 VTAIL.n183 VTAIL.n181 2.24188
R493 VTAIL.n168 VTAIL.n144 1.93989
R494 VTAIL.n30 VTAIL.n6 1.93989
R495 VTAIL.n127 VTAIL.n103 1.93989
R496 VTAIL.n81 VTAIL.n57 1.93989
R497 VTAIL VTAIL.n1 1.73972
R498 VTAIL.n95 VTAIL.n93 1.59102
R499 VTAIL.n43 VTAIL.n1 1.59102
R500 VTAIL.n173 VTAIL.n171 1.16414
R501 VTAIL.n180 VTAIL.n140 1.16414
R502 VTAIL.n35 VTAIL.n33 1.16414
R503 VTAIL.n42 VTAIL.n2 1.16414
R504 VTAIL.n138 VTAIL.n98 1.16414
R505 VTAIL.n131 VTAIL.n130 1.16414
R506 VTAIL.n92 VTAIL.n52 1.16414
R507 VTAIL.n85 VTAIL.n84 1.16414
R508 VTAIL VTAIL.n183 0.502655
R509 VTAIL.n172 VTAIL.n142 0.388379
R510 VTAIL.n178 VTAIL.n177 0.388379
R511 VTAIL.n34 VTAIL.n4 0.388379
R512 VTAIL.n40 VTAIL.n39 0.388379
R513 VTAIL.n136 VTAIL.n135 0.388379
R514 VTAIL.n102 VTAIL.n100 0.388379
R515 VTAIL.n90 VTAIL.n89 0.388379
R516 VTAIL.n56 VTAIL.n54 0.388379
R517 VTAIL.n154 VTAIL.n149 0.155672
R518 VTAIL.n161 VTAIL.n149 0.155672
R519 VTAIL.n162 VTAIL.n161 0.155672
R520 VTAIL.n162 VTAIL.n145 0.155672
R521 VTAIL.n169 VTAIL.n145 0.155672
R522 VTAIL.n170 VTAIL.n169 0.155672
R523 VTAIL.n170 VTAIL.n141 0.155672
R524 VTAIL.n179 VTAIL.n141 0.155672
R525 VTAIL.n16 VTAIL.n11 0.155672
R526 VTAIL.n23 VTAIL.n11 0.155672
R527 VTAIL.n24 VTAIL.n23 0.155672
R528 VTAIL.n24 VTAIL.n7 0.155672
R529 VTAIL.n31 VTAIL.n7 0.155672
R530 VTAIL.n32 VTAIL.n31 0.155672
R531 VTAIL.n32 VTAIL.n3 0.155672
R532 VTAIL.n41 VTAIL.n3 0.155672
R533 VTAIL.n137 VTAIL.n99 0.155672
R534 VTAIL.n129 VTAIL.n99 0.155672
R535 VTAIL.n129 VTAIL.n128 0.155672
R536 VTAIL.n128 VTAIL.n104 0.155672
R537 VTAIL.n121 VTAIL.n104 0.155672
R538 VTAIL.n121 VTAIL.n120 0.155672
R539 VTAIL.n120 VTAIL.n108 0.155672
R540 VTAIL.n113 VTAIL.n108 0.155672
R541 VTAIL.n91 VTAIL.n53 0.155672
R542 VTAIL.n83 VTAIL.n53 0.155672
R543 VTAIL.n83 VTAIL.n82 0.155672
R544 VTAIL.n82 VTAIL.n58 0.155672
R545 VTAIL.n75 VTAIL.n58 0.155672
R546 VTAIL.n75 VTAIL.n74 0.155672
R547 VTAIL.n74 VTAIL.n62 0.155672
R548 VTAIL.n67 VTAIL.n62 0.155672
R549 B.n651 B.n650 585
R550 B.n653 B.n138 585
R551 B.n656 B.n655 585
R552 B.n657 B.n137 585
R553 B.n659 B.n658 585
R554 B.n661 B.n136 585
R555 B.n664 B.n663 585
R556 B.n665 B.n135 585
R557 B.n667 B.n666 585
R558 B.n669 B.n134 585
R559 B.n672 B.n671 585
R560 B.n673 B.n133 585
R561 B.n675 B.n674 585
R562 B.n677 B.n132 585
R563 B.n680 B.n679 585
R564 B.n681 B.n131 585
R565 B.n683 B.n682 585
R566 B.n685 B.n130 585
R567 B.n688 B.n687 585
R568 B.n689 B.n129 585
R569 B.n691 B.n690 585
R570 B.n693 B.n128 585
R571 B.n696 B.n695 585
R572 B.n697 B.n127 585
R573 B.n699 B.n698 585
R574 B.n701 B.n126 585
R575 B.n704 B.n703 585
R576 B.n705 B.n122 585
R577 B.n707 B.n706 585
R578 B.n709 B.n121 585
R579 B.n712 B.n711 585
R580 B.n713 B.n120 585
R581 B.n715 B.n714 585
R582 B.n717 B.n119 585
R583 B.n720 B.n719 585
R584 B.n721 B.n118 585
R585 B.n723 B.n722 585
R586 B.n725 B.n117 585
R587 B.n728 B.n727 585
R588 B.n730 B.n114 585
R589 B.n732 B.n731 585
R590 B.n734 B.n113 585
R591 B.n737 B.n736 585
R592 B.n738 B.n112 585
R593 B.n740 B.n739 585
R594 B.n742 B.n111 585
R595 B.n745 B.n744 585
R596 B.n746 B.n110 585
R597 B.n748 B.n747 585
R598 B.n750 B.n109 585
R599 B.n753 B.n752 585
R600 B.n754 B.n108 585
R601 B.n756 B.n755 585
R602 B.n758 B.n107 585
R603 B.n761 B.n760 585
R604 B.n762 B.n106 585
R605 B.n764 B.n763 585
R606 B.n766 B.n105 585
R607 B.n769 B.n768 585
R608 B.n770 B.n104 585
R609 B.n772 B.n771 585
R610 B.n774 B.n103 585
R611 B.n777 B.n776 585
R612 B.n778 B.n102 585
R613 B.n780 B.n779 585
R614 B.n782 B.n101 585
R615 B.n785 B.n784 585
R616 B.n786 B.n100 585
R617 B.n649 B.n98 585
R618 B.n789 B.n98 585
R619 B.n648 B.n97 585
R620 B.n790 B.n97 585
R621 B.n647 B.n96 585
R622 B.n791 B.n96 585
R623 B.n646 B.n645 585
R624 B.n645 B.n92 585
R625 B.n644 B.n91 585
R626 B.n797 B.n91 585
R627 B.n643 B.n90 585
R628 B.n798 B.n90 585
R629 B.n642 B.n89 585
R630 B.n799 B.n89 585
R631 B.n641 B.n640 585
R632 B.n640 B.n88 585
R633 B.n639 B.n84 585
R634 B.n805 B.n84 585
R635 B.n638 B.n83 585
R636 B.n806 B.n83 585
R637 B.n637 B.n82 585
R638 B.n807 B.n82 585
R639 B.n636 B.n635 585
R640 B.n635 B.n78 585
R641 B.n634 B.n77 585
R642 B.n813 B.n77 585
R643 B.n633 B.n76 585
R644 B.n814 B.n76 585
R645 B.n632 B.n75 585
R646 B.n815 B.n75 585
R647 B.n631 B.n630 585
R648 B.n630 B.n71 585
R649 B.n629 B.n70 585
R650 B.n821 B.n70 585
R651 B.n628 B.n69 585
R652 B.n822 B.n69 585
R653 B.n627 B.n68 585
R654 B.n823 B.n68 585
R655 B.n626 B.n625 585
R656 B.n625 B.n64 585
R657 B.n624 B.n63 585
R658 B.n829 B.n63 585
R659 B.n623 B.n62 585
R660 B.n830 B.n62 585
R661 B.n622 B.n61 585
R662 B.n831 B.n61 585
R663 B.n621 B.n620 585
R664 B.n620 B.n57 585
R665 B.n619 B.n56 585
R666 B.n837 B.n56 585
R667 B.n618 B.n55 585
R668 B.n838 B.n55 585
R669 B.n617 B.n54 585
R670 B.n839 B.n54 585
R671 B.n616 B.n615 585
R672 B.n615 B.n50 585
R673 B.n614 B.n49 585
R674 B.n845 B.n49 585
R675 B.n613 B.n48 585
R676 B.n846 B.n48 585
R677 B.n612 B.n47 585
R678 B.n847 B.n47 585
R679 B.n611 B.n610 585
R680 B.n610 B.n43 585
R681 B.n609 B.n42 585
R682 B.n853 B.n42 585
R683 B.n608 B.n41 585
R684 B.n854 B.n41 585
R685 B.n607 B.n40 585
R686 B.n855 B.n40 585
R687 B.n606 B.n605 585
R688 B.n605 B.n36 585
R689 B.n604 B.n35 585
R690 B.n861 B.n35 585
R691 B.n603 B.n34 585
R692 B.n862 B.n34 585
R693 B.n602 B.n33 585
R694 B.n863 B.n33 585
R695 B.n601 B.n600 585
R696 B.n600 B.n29 585
R697 B.n599 B.n28 585
R698 B.n869 B.n28 585
R699 B.n598 B.n27 585
R700 B.n870 B.n27 585
R701 B.n597 B.n26 585
R702 B.n871 B.n26 585
R703 B.n596 B.n595 585
R704 B.n595 B.n22 585
R705 B.n594 B.n21 585
R706 B.n877 B.n21 585
R707 B.n593 B.n20 585
R708 B.n878 B.n20 585
R709 B.n592 B.n19 585
R710 B.n879 B.n19 585
R711 B.n591 B.n590 585
R712 B.n590 B.n15 585
R713 B.n589 B.n14 585
R714 B.n885 B.n14 585
R715 B.n588 B.n13 585
R716 B.n886 B.n13 585
R717 B.n587 B.n12 585
R718 B.n887 B.n12 585
R719 B.n586 B.n585 585
R720 B.n585 B.n8 585
R721 B.n584 B.n7 585
R722 B.n893 B.n7 585
R723 B.n583 B.n6 585
R724 B.n894 B.n6 585
R725 B.n582 B.n5 585
R726 B.n895 B.n5 585
R727 B.n581 B.n580 585
R728 B.n580 B.n4 585
R729 B.n579 B.n139 585
R730 B.n579 B.n578 585
R731 B.n569 B.n140 585
R732 B.n141 B.n140 585
R733 B.n571 B.n570 585
R734 B.n572 B.n571 585
R735 B.n568 B.n146 585
R736 B.n146 B.n145 585
R737 B.n567 B.n566 585
R738 B.n566 B.n565 585
R739 B.n148 B.n147 585
R740 B.n149 B.n148 585
R741 B.n558 B.n557 585
R742 B.n559 B.n558 585
R743 B.n556 B.n154 585
R744 B.n154 B.n153 585
R745 B.n555 B.n554 585
R746 B.n554 B.n553 585
R747 B.n156 B.n155 585
R748 B.n157 B.n156 585
R749 B.n546 B.n545 585
R750 B.n547 B.n546 585
R751 B.n544 B.n162 585
R752 B.n162 B.n161 585
R753 B.n543 B.n542 585
R754 B.n542 B.n541 585
R755 B.n164 B.n163 585
R756 B.n165 B.n164 585
R757 B.n534 B.n533 585
R758 B.n535 B.n534 585
R759 B.n532 B.n170 585
R760 B.n170 B.n169 585
R761 B.n531 B.n530 585
R762 B.n530 B.n529 585
R763 B.n172 B.n171 585
R764 B.n173 B.n172 585
R765 B.n522 B.n521 585
R766 B.n523 B.n522 585
R767 B.n520 B.n177 585
R768 B.n181 B.n177 585
R769 B.n519 B.n518 585
R770 B.n518 B.n517 585
R771 B.n179 B.n178 585
R772 B.n180 B.n179 585
R773 B.n510 B.n509 585
R774 B.n511 B.n510 585
R775 B.n508 B.n186 585
R776 B.n186 B.n185 585
R777 B.n507 B.n506 585
R778 B.n506 B.n505 585
R779 B.n188 B.n187 585
R780 B.n189 B.n188 585
R781 B.n498 B.n497 585
R782 B.n499 B.n498 585
R783 B.n496 B.n193 585
R784 B.n197 B.n193 585
R785 B.n495 B.n494 585
R786 B.n494 B.n493 585
R787 B.n195 B.n194 585
R788 B.n196 B.n195 585
R789 B.n486 B.n485 585
R790 B.n487 B.n486 585
R791 B.n484 B.n202 585
R792 B.n202 B.n201 585
R793 B.n483 B.n482 585
R794 B.n482 B.n481 585
R795 B.n204 B.n203 585
R796 B.n205 B.n204 585
R797 B.n474 B.n473 585
R798 B.n475 B.n474 585
R799 B.n472 B.n209 585
R800 B.n213 B.n209 585
R801 B.n471 B.n470 585
R802 B.n470 B.n469 585
R803 B.n211 B.n210 585
R804 B.n212 B.n211 585
R805 B.n462 B.n461 585
R806 B.n463 B.n462 585
R807 B.n460 B.n218 585
R808 B.n218 B.n217 585
R809 B.n459 B.n458 585
R810 B.n458 B.n457 585
R811 B.n220 B.n219 585
R812 B.n221 B.n220 585
R813 B.n450 B.n449 585
R814 B.n451 B.n450 585
R815 B.n448 B.n226 585
R816 B.n226 B.n225 585
R817 B.n447 B.n446 585
R818 B.n446 B.n445 585
R819 B.n228 B.n227 585
R820 B.n438 B.n228 585
R821 B.n437 B.n436 585
R822 B.n439 B.n437 585
R823 B.n435 B.n233 585
R824 B.n233 B.n232 585
R825 B.n434 B.n433 585
R826 B.n433 B.n432 585
R827 B.n235 B.n234 585
R828 B.n236 B.n235 585
R829 B.n425 B.n424 585
R830 B.n426 B.n425 585
R831 B.n423 B.n241 585
R832 B.n241 B.n240 585
R833 B.n422 B.n421 585
R834 B.n421 B.n420 585
R835 B.n417 B.n245 585
R836 B.n416 B.n415 585
R837 B.n413 B.n246 585
R838 B.n413 B.n244 585
R839 B.n412 B.n411 585
R840 B.n410 B.n409 585
R841 B.n408 B.n248 585
R842 B.n406 B.n405 585
R843 B.n404 B.n249 585
R844 B.n403 B.n402 585
R845 B.n400 B.n250 585
R846 B.n398 B.n397 585
R847 B.n396 B.n251 585
R848 B.n395 B.n394 585
R849 B.n392 B.n252 585
R850 B.n390 B.n389 585
R851 B.n388 B.n253 585
R852 B.n387 B.n386 585
R853 B.n384 B.n254 585
R854 B.n382 B.n381 585
R855 B.n380 B.n255 585
R856 B.n379 B.n378 585
R857 B.n376 B.n256 585
R858 B.n374 B.n373 585
R859 B.n372 B.n257 585
R860 B.n371 B.n370 585
R861 B.n368 B.n258 585
R862 B.n366 B.n365 585
R863 B.n364 B.n259 585
R864 B.n363 B.n362 585
R865 B.n360 B.n359 585
R866 B.n358 B.n357 585
R867 B.n356 B.n264 585
R868 B.n354 B.n353 585
R869 B.n352 B.n265 585
R870 B.n351 B.n350 585
R871 B.n348 B.n266 585
R872 B.n346 B.n345 585
R873 B.n344 B.n267 585
R874 B.n343 B.n342 585
R875 B.n340 B.n339 585
R876 B.n338 B.n337 585
R877 B.n336 B.n272 585
R878 B.n334 B.n333 585
R879 B.n332 B.n273 585
R880 B.n331 B.n330 585
R881 B.n328 B.n274 585
R882 B.n326 B.n325 585
R883 B.n324 B.n275 585
R884 B.n323 B.n322 585
R885 B.n320 B.n276 585
R886 B.n318 B.n317 585
R887 B.n316 B.n277 585
R888 B.n315 B.n314 585
R889 B.n312 B.n278 585
R890 B.n310 B.n309 585
R891 B.n308 B.n279 585
R892 B.n307 B.n306 585
R893 B.n304 B.n280 585
R894 B.n302 B.n301 585
R895 B.n300 B.n281 585
R896 B.n299 B.n298 585
R897 B.n296 B.n282 585
R898 B.n294 B.n293 585
R899 B.n292 B.n283 585
R900 B.n291 B.n290 585
R901 B.n288 B.n284 585
R902 B.n286 B.n285 585
R903 B.n243 B.n242 585
R904 B.n244 B.n243 585
R905 B.n419 B.n418 585
R906 B.n420 B.n419 585
R907 B.n239 B.n238 585
R908 B.n240 B.n239 585
R909 B.n428 B.n427 585
R910 B.n427 B.n426 585
R911 B.n429 B.n237 585
R912 B.n237 B.n236 585
R913 B.n431 B.n430 585
R914 B.n432 B.n431 585
R915 B.n231 B.n230 585
R916 B.n232 B.n231 585
R917 B.n441 B.n440 585
R918 B.n440 B.n439 585
R919 B.n442 B.n229 585
R920 B.n438 B.n229 585
R921 B.n444 B.n443 585
R922 B.n445 B.n444 585
R923 B.n224 B.n223 585
R924 B.n225 B.n224 585
R925 B.n453 B.n452 585
R926 B.n452 B.n451 585
R927 B.n454 B.n222 585
R928 B.n222 B.n221 585
R929 B.n456 B.n455 585
R930 B.n457 B.n456 585
R931 B.n216 B.n215 585
R932 B.n217 B.n216 585
R933 B.n465 B.n464 585
R934 B.n464 B.n463 585
R935 B.n466 B.n214 585
R936 B.n214 B.n212 585
R937 B.n468 B.n467 585
R938 B.n469 B.n468 585
R939 B.n208 B.n207 585
R940 B.n213 B.n208 585
R941 B.n477 B.n476 585
R942 B.n476 B.n475 585
R943 B.n478 B.n206 585
R944 B.n206 B.n205 585
R945 B.n480 B.n479 585
R946 B.n481 B.n480 585
R947 B.n200 B.n199 585
R948 B.n201 B.n200 585
R949 B.n489 B.n488 585
R950 B.n488 B.n487 585
R951 B.n490 B.n198 585
R952 B.n198 B.n196 585
R953 B.n492 B.n491 585
R954 B.n493 B.n492 585
R955 B.n192 B.n191 585
R956 B.n197 B.n192 585
R957 B.n501 B.n500 585
R958 B.n500 B.n499 585
R959 B.n502 B.n190 585
R960 B.n190 B.n189 585
R961 B.n504 B.n503 585
R962 B.n505 B.n504 585
R963 B.n184 B.n183 585
R964 B.n185 B.n184 585
R965 B.n513 B.n512 585
R966 B.n512 B.n511 585
R967 B.n514 B.n182 585
R968 B.n182 B.n180 585
R969 B.n516 B.n515 585
R970 B.n517 B.n516 585
R971 B.n176 B.n175 585
R972 B.n181 B.n176 585
R973 B.n525 B.n524 585
R974 B.n524 B.n523 585
R975 B.n526 B.n174 585
R976 B.n174 B.n173 585
R977 B.n528 B.n527 585
R978 B.n529 B.n528 585
R979 B.n168 B.n167 585
R980 B.n169 B.n168 585
R981 B.n537 B.n536 585
R982 B.n536 B.n535 585
R983 B.n538 B.n166 585
R984 B.n166 B.n165 585
R985 B.n540 B.n539 585
R986 B.n541 B.n540 585
R987 B.n160 B.n159 585
R988 B.n161 B.n160 585
R989 B.n549 B.n548 585
R990 B.n548 B.n547 585
R991 B.n550 B.n158 585
R992 B.n158 B.n157 585
R993 B.n552 B.n551 585
R994 B.n553 B.n552 585
R995 B.n152 B.n151 585
R996 B.n153 B.n152 585
R997 B.n561 B.n560 585
R998 B.n560 B.n559 585
R999 B.n562 B.n150 585
R1000 B.n150 B.n149 585
R1001 B.n564 B.n563 585
R1002 B.n565 B.n564 585
R1003 B.n144 B.n143 585
R1004 B.n145 B.n144 585
R1005 B.n574 B.n573 585
R1006 B.n573 B.n572 585
R1007 B.n575 B.n142 585
R1008 B.n142 B.n141 585
R1009 B.n577 B.n576 585
R1010 B.n578 B.n577 585
R1011 B.n2 B.n0 585
R1012 B.n4 B.n2 585
R1013 B.n3 B.n1 585
R1014 B.n894 B.n3 585
R1015 B.n892 B.n891 585
R1016 B.n893 B.n892 585
R1017 B.n890 B.n9 585
R1018 B.n9 B.n8 585
R1019 B.n889 B.n888 585
R1020 B.n888 B.n887 585
R1021 B.n11 B.n10 585
R1022 B.n886 B.n11 585
R1023 B.n884 B.n883 585
R1024 B.n885 B.n884 585
R1025 B.n882 B.n16 585
R1026 B.n16 B.n15 585
R1027 B.n881 B.n880 585
R1028 B.n880 B.n879 585
R1029 B.n18 B.n17 585
R1030 B.n878 B.n18 585
R1031 B.n876 B.n875 585
R1032 B.n877 B.n876 585
R1033 B.n874 B.n23 585
R1034 B.n23 B.n22 585
R1035 B.n873 B.n872 585
R1036 B.n872 B.n871 585
R1037 B.n25 B.n24 585
R1038 B.n870 B.n25 585
R1039 B.n868 B.n867 585
R1040 B.n869 B.n868 585
R1041 B.n866 B.n30 585
R1042 B.n30 B.n29 585
R1043 B.n865 B.n864 585
R1044 B.n864 B.n863 585
R1045 B.n32 B.n31 585
R1046 B.n862 B.n32 585
R1047 B.n860 B.n859 585
R1048 B.n861 B.n860 585
R1049 B.n858 B.n37 585
R1050 B.n37 B.n36 585
R1051 B.n857 B.n856 585
R1052 B.n856 B.n855 585
R1053 B.n39 B.n38 585
R1054 B.n854 B.n39 585
R1055 B.n852 B.n851 585
R1056 B.n853 B.n852 585
R1057 B.n850 B.n44 585
R1058 B.n44 B.n43 585
R1059 B.n849 B.n848 585
R1060 B.n848 B.n847 585
R1061 B.n46 B.n45 585
R1062 B.n846 B.n46 585
R1063 B.n844 B.n843 585
R1064 B.n845 B.n844 585
R1065 B.n842 B.n51 585
R1066 B.n51 B.n50 585
R1067 B.n841 B.n840 585
R1068 B.n840 B.n839 585
R1069 B.n53 B.n52 585
R1070 B.n838 B.n53 585
R1071 B.n836 B.n835 585
R1072 B.n837 B.n836 585
R1073 B.n834 B.n58 585
R1074 B.n58 B.n57 585
R1075 B.n833 B.n832 585
R1076 B.n832 B.n831 585
R1077 B.n60 B.n59 585
R1078 B.n830 B.n60 585
R1079 B.n828 B.n827 585
R1080 B.n829 B.n828 585
R1081 B.n826 B.n65 585
R1082 B.n65 B.n64 585
R1083 B.n825 B.n824 585
R1084 B.n824 B.n823 585
R1085 B.n67 B.n66 585
R1086 B.n822 B.n67 585
R1087 B.n820 B.n819 585
R1088 B.n821 B.n820 585
R1089 B.n818 B.n72 585
R1090 B.n72 B.n71 585
R1091 B.n817 B.n816 585
R1092 B.n816 B.n815 585
R1093 B.n74 B.n73 585
R1094 B.n814 B.n74 585
R1095 B.n812 B.n811 585
R1096 B.n813 B.n812 585
R1097 B.n810 B.n79 585
R1098 B.n79 B.n78 585
R1099 B.n809 B.n808 585
R1100 B.n808 B.n807 585
R1101 B.n81 B.n80 585
R1102 B.n806 B.n81 585
R1103 B.n804 B.n803 585
R1104 B.n805 B.n804 585
R1105 B.n802 B.n85 585
R1106 B.n88 B.n85 585
R1107 B.n801 B.n800 585
R1108 B.n800 B.n799 585
R1109 B.n87 B.n86 585
R1110 B.n798 B.n87 585
R1111 B.n796 B.n795 585
R1112 B.n797 B.n796 585
R1113 B.n794 B.n93 585
R1114 B.n93 B.n92 585
R1115 B.n793 B.n792 585
R1116 B.n792 B.n791 585
R1117 B.n95 B.n94 585
R1118 B.n790 B.n95 585
R1119 B.n788 B.n787 585
R1120 B.n789 B.n788 585
R1121 B.n897 B.n896 585
R1122 B.n896 B.n895 585
R1123 B.n419 B.n245 530.939
R1124 B.n788 B.n100 530.939
R1125 B.n421 B.n243 530.939
R1126 B.n651 B.n98 530.939
R1127 B.n268 B.t10 290.829
R1128 B.n260 B.t18 290.829
R1129 B.n115 B.t21 290.829
R1130 B.n123 B.t14 290.829
R1131 B.n268 B.t13 260.807
R1132 B.n123 B.t16 260.807
R1133 B.n260 B.t20 260.807
R1134 B.n115 B.t22 260.807
R1135 B.n652 B.n99 256.663
R1136 B.n654 B.n99 256.663
R1137 B.n660 B.n99 256.663
R1138 B.n662 B.n99 256.663
R1139 B.n668 B.n99 256.663
R1140 B.n670 B.n99 256.663
R1141 B.n676 B.n99 256.663
R1142 B.n678 B.n99 256.663
R1143 B.n684 B.n99 256.663
R1144 B.n686 B.n99 256.663
R1145 B.n692 B.n99 256.663
R1146 B.n694 B.n99 256.663
R1147 B.n700 B.n99 256.663
R1148 B.n702 B.n99 256.663
R1149 B.n708 B.n99 256.663
R1150 B.n710 B.n99 256.663
R1151 B.n716 B.n99 256.663
R1152 B.n718 B.n99 256.663
R1153 B.n724 B.n99 256.663
R1154 B.n726 B.n99 256.663
R1155 B.n733 B.n99 256.663
R1156 B.n735 B.n99 256.663
R1157 B.n741 B.n99 256.663
R1158 B.n743 B.n99 256.663
R1159 B.n749 B.n99 256.663
R1160 B.n751 B.n99 256.663
R1161 B.n757 B.n99 256.663
R1162 B.n759 B.n99 256.663
R1163 B.n765 B.n99 256.663
R1164 B.n767 B.n99 256.663
R1165 B.n773 B.n99 256.663
R1166 B.n775 B.n99 256.663
R1167 B.n781 B.n99 256.663
R1168 B.n783 B.n99 256.663
R1169 B.n414 B.n244 256.663
R1170 B.n247 B.n244 256.663
R1171 B.n407 B.n244 256.663
R1172 B.n401 B.n244 256.663
R1173 B.n399 B.n244 256.663
R1174 B.n393 B.n244 256.663
R1175 B.n391 B.n244 256.663
R1176 B.n385 B.n244 256.663
R1177 B.n383 B.n244 256.663
R1178 B.n377 B.n244 256.663
R1179 B.n375 B.n244 256.663
R1180 B.n369 B.n244 256.663
R1181 B.n367 B.n244 256.663
R1182 B.n361 B.n244 256.663
R1183 B.n263 B.n244 256.663
R1184 B.n355 B.n244 256.663
R1185 B.n349 B.n244 256.663
R1186 B.n347 B.n244 256.663
R1187 B.n341 B.n244 256.663
R1188 B.n271 B.n244 256.663
R1189 B.n335 B.n244 256.663
R1190 B.n329 B.n244 256.663
R1191 B.n327 B.n244 256.663
R1192 B.n321 B.n244 256.663
R1193 B.n319 B.n244 256.663
R1194 B.n313 B.n244 256.663
R1195 B.n311 B.n244 256.663
R1196 B.n305 B.n244 256.663
R1197 B.n303 B.n244 256.663
R1198 B.n297 B.n244 256.663
R1199 B.n295 B.n244 256.663
R1200 B.n289 B.n244 256.663
R1201 B.n287 B.n244 256.663
R1202 B.n269 B.t12 210.382
R1203 B.n124 B.t17 210.382
R1204 B.n261 B.t19 210.382
R1205 B.n116 B.t23 210.382
R1206 B.n419 B.n239 163.367
R1207 B.n427 B.n239 163.367
R1208 B.n427 B.n237 163.367
R1209 B.n431 B.n237 163.367
R1210 B.n431 B.n231 163.367
R1211 B.n440 B.n231 163.367
R1212 B.n440 B.n229 163.367
R1213 B.n444 B.n229 163.367
R1214 B.n444 B.n224 163.367
R1215 B.n452 B.n224 163.367
R1216 B.n452 B.n222 163.367
R1217 B.n456 B.n222 163.367
R1218 B.n456 B.n216 163.367
R1219 B.n464 B.n216 163.367
R1220 B.n464 B.n214 163.367
R1221 B.n468 B.n214 163.367
R1222 B.n468 B.n208 163.367
R1223 B.n476 B.n208 163.367
R1224 B.n476 B.n206 163.367
R1225 B.n480 B.n206 163.367
R1226 B.n480 B.n200 163.367
R1227 B.n488 B.n200 163.367
R1228 B.n488 B.n198 163.367
R1229 B.n492 B.n198 163.367
R1230 B.n492 B.n192 163.367
R1231 B.n500 B.n192 163.367
R1232 B.n500 B.n190 163.367
R1233 B.n504 B.n190 163.367
R1234 B.n504 B.n184 163.367
R1235 B.n512 B.n184 163.367
R1236 B.n512 B.n182 163.367
R1237 B.n516 B.n182 163.367
R1238 B.n516 B.n176 163.367
R1239 B.n524 B.n176 163.367
R1240 B.n524 B.n174 163.367
R1241 B.n528 B.n174 163.367
R1242 B.n528 B.n168 163.367
R1243 B.n536 B.n168 163.367
R1244 B.n536 B.n166 163.367
R1245 B.n540 B.n166 163.367
R1246 B.n540 B.n160 163.367
R1247 B.n548 B.n160 163.367
R1248 B.n548 B.n158 163.367
R1249 B.n552 B.n158 163.367
R1250 B.n552 B.n152 163.367
R1251 B.n560 B.n152 163.367
R1252 B.n560 B.n150 163.367
R1253 B.n564 B.n150 163.367
R1254 B.n564 B.n144 163.367
R1255 B.n573 B.n144 163.367
R1256 B.n573 B.n142 163.367
R1257 B.n577 B.n142 163.367
R1258 B.n577 B.n2 163.367
R1259 B.n896 B.n2 163.367
R1260 B.n896 B.n3 163.367
R1261 B.n892 B.n3 163.367
R1262 B.n892 B.n9 163.367
R1263 B.n888 B.n9 163.367
R1264 B.n888 B.n11 163.367
R1265 B.n884 B.n11 163.367
R1266 B.n884 B.n16 163.367
R1267 B.n880 B.n16 163.367
R1268 B.n880 B.n18 163.367
R1269 B.n876 B.n18 163.367
R1270 B.n876 B.n23 163.367
R1271 B.n872 B.n23 163.367
R1272 B.n872 B.n25 163.367
R1273 B.n868 B.n25 163.367
R1274 B.n868 B.n30 163.367
R1275 B.n864 B.n30 163.367
R1276 B.n864 B.n32 163.367
R1277 B.n860 B.n32 163.367
R1278 B.n860 B.n37 163.367
R1279 B.n856 B.n37 163.367
R1280 B.n856 B.n39 163.367
R1281 B.n852 B.n39 163.367
R1282 B.n852 B.n44 163.367
R1283 B.n848 B.n44 163.367
R1284 B.n848 B.n46 163.367
R1285 B.n844 B.n46 163.367
R1286 B.n844 B.n51 163.367
R1287 B.n840 B.n51 163.367
R1288 B.n840 B.n53 163.367
R1289 B.n836 B.n53 163.367
R1290 B.n836 B.n58 163.367
R1291 B.n832 B.n58 163.367
R1292 B.n832 B.n60 163.367
R1293 B.n828 B.n60 163.367
R1294 B.n828 B.n65 163.367
R1295 B.n824 B.n65 163.367
R1296 B.n824 B.n67 163.367
R1297 B.n820 B.n67 163.367
R1298 B.n820 B.n72 163.367
R1299 B.n816 B.n72 163.367
R1300 B.n816 B.n74 163.367
R1301 B.n812 B.n74 163.367
R1302 B.n812 B.n79 163.367
R1303 B.n808 B.n79 163.367
R1304 B.n808 B.n81 163.367
R1305 B.n804 B.n81 163.367
R1306 B.n804 B.n85 163.367
R1307 B.n800 B.n85 163.367
R1308 B.n800 B.n87 163.367
R1309 B.n796 B.n87 163.367
R1310 B.n796 B.n93 163.367
R1311 B.n792 B.n93 163.367
R1312 B.n792 B.n95 163.367
R1313 B.n788 B.n95 163.367
R1314 B.n415 B.n413 163.367
R1315 B.n413 B.n412 163.367
R1316 B.n409 B.n408 163.367
R1317 B.n406 B.n249 163.367
R1318 B.n402 B.n400 163.367
R1319 B.n398 B.n251 163.367
R1320 B.n394 B.n392 163.367
R1321 B.n390 B.n253 163.367
R1322 B.n386 B.n384 163.367
R1323 B.n382 B.n255 163.367
R1324 B.n378 B.n376 163.367
R1325 B.n374 B.n257 163.367
R1326 B.n370 B.n368 163.367
R1327 B.n366 B.n259 163.367
R1328 B.n362 B.n360 163.367
R1329 B.n357 B.n356 163.367
R1330 B.n354 B.n265 163.367
R1331 B.n350 B.n348 163.367
R1332 B.n346 B.n267 163.367
R1333 B.n342 B.n340 163.367
R1334 B.n337 B.n336 163.367
R1335 B.n334 B.n273 163.367
R1336 B.n330 B.n328 163.367
R1337 B.n326 B.n275 163.367
R1338 B.n322 B.n320 163.367
R1339 B.n318 B.n277 163.367
R1340 B.n314 B.n312 163.367
R1341 B.n310 B.n279 163.367
R1342 B.n306 B.n304 163.367
R1343 B.n302 B.n281 163.367
R1344 B.n298 B.n296 163.367
R1345 B.n294 B.n283 163.367
R1346 B.n290 B.n288 163.367
R1347 B.n286 B.n243 163.367
R1348 B.n421 B.n241 163.367
R1349 B.n425 B.n241 163.367
R1350 B.n425 B.n235 163.367
R1351 B.n433 B.n235 163.367
R1352 B.n433 B.n233 163.367
R1353 B.n437 B.n233 163.367
R1354 B.n437 B.n228 163.367
R1355 B.n446 B.n228 163.367
R1356 B.n446 B.n226 163.367
R1357 B.n450 B.n226 163.367
R1358 B.n450 B.n220 163.367
R1359 B.n458 B.n220 163.367
R1360 B.n458 B.n218 163.367
R1361 B.n462 B.n218 163.367
R1362 B.n462 B.n211 163.367
R1363 B.n470 B.n211 163.367
R1364 B.n470 B.n209 163.367
R1365 B.n474 B.n209 163.367
R1366 B.n474 B.n204 163.367
R1367 B.n482 B.n204 163.367
R1368 B.n482 B.n202 163.367
R1369 B.n486 B.n202 163.367
R1370 B.n486 B.n195 163.367
R1371 B.n494 B.n195 163.367
R1372 B.n494 B.n193 163.367
R1373 B.n498 B.n193 163.367
R1374 B.n498 B.n188 163.367
R1375 B.n506 B.n188 163.367
R1376 B.n506 B.n186 163.367
R1377 B.n510 B.n186 163.367
R1378 B.n510 B.n179 163.367
R1379 B.n518 B.n179 163.367
R1380 B.n518 B.n177 163.367
R1381 B.n522 B.n177 163.367
R1382 B.n522 B.n172 163.367
R1383 B.n530 B.n172 163.367
R1384 B.n530 B.n170 163.367
R1385 B.n534 B.n170 163.367
R1386 B.n534 B.n164 163.367
R1387 B.n542 B.n164 163.367
R1388 B.n542 B.n162 163.367
R1389 B.n546 B.n162 163.367
R1390 B.n546 B.n156 163.367
R1391 B.n554 B.n156 163.367
R1392 B.n554 B.n154 163.367
R1393 B.n558 B.n154 163.367
R1394 B.n558 B.n148 163.367
R1395 B.n566 B.n148 163.367
R1396 B.n566 B.n146 163.367
R1397 B.n571 B.n146 163.367
R1398 B.n571 B.n140 163.367
R1399 B.n579 B.n140 163.367
R1400 B.n580 B.n579 163.367
R1401 B.n580 B.n5 163.367
R1402 B.n6 B.n5 163.367
R1403 B.n7 B.n6 163.367
R1404 B.n585 B.n7 163.367
R1405 B.n585 B.n12 163.367
R1406 B.n13 B.n12 163.367
R1407 B.n14 B.n13 163.367
R1408 B.n590 B.n14 163.367
R1409 B.n590 B.n19 163.367
R1410 B.n20 B.n19 163.367
R1411 B.n21 B.n20 163.367
R1412 B.n595 B.n21 163.367
R1413 B.n595 B.n26 163.367
R1414 B.n27 B.n26 163.367
R1415 B.n28 B.n27 163.367
R1416 B.n600 B.n28 163.367
R1417 B.n600 B.n33 163.367
R1418 B.n34 B.n33 163.367
R1419 B.n35 B.n34 163.367
R1420 B.n605 B.n35 163.367
R1421 B.n605 B.n40 163.367
R1422 B.n41 B.n40 163.367
R1423 B.n42 B.n41 163.367
R1424 B.n610 B.n42 163.367
R1425 B.n610 B.n47 163.367
R1426 B.n48 B.n47 163.367
R1427 B.n49 B.n48 163.367
R1428 B.n615 B.n49 163.367
R1429 B.n615 B.n54 163.367
R1430 B.n55 B.n54 163.367
R1431 B.n56 B.n55 163.367
R1432 B.n620 B.n56 163.367
R1433 B.n620 B.n61 163.367
R1434 B.n62 B.n61 163.367
R1435 B.n63 B.n62 163.367
R1436 B.n625 B.n63 163.367
R1437 B.n625 B.n68 163.367
R1438 B.n69 B.n68 163.367
R1439 B.n70 B.n69 163.367
R1440 B.n630 B.n70 163.367
R1441 B.n630 B.n75 163.367
R1442 B.n76 B.n75 163.367
R1443 B.n77 B.n76 163.367
R1444 B.n635 B.n77 163.367
R1445 B.n635 B.n82 163.367
R1446 B.n83 B.n82 163.367
R1447 B.n84 B.n83 163.367
R1448 B.n640 B.n84 163.367
R1449 B.n640 B.n89 163.367
R1450 B.n90 B.n89 163.367
R1451 B.n91 B.n90 163.367
R1452 B.n645 B.n91 163.367
R1453 B.n645 B.n96 163.367
R1454 B.n97 B.n96 163.367
R1455 B.n98 B.n97 163.367
R1456 B.n784 B.n782 163.367
R1457 B.n780 B.n102 163.367
R1458 B.n776 B.n774 163.367
R1459 B.n772 B.n104 163.367
R1460 B.n768 B.n766 163.367
R1461 B.n764 B.n106 163.367
R1462 B.n760 B.n758 163.367
R1463 B.n756 B.n108 163.367
R1464 B.n752 B.n750 163.367
R1465 B.n748 B.n110 163.367
R1466 B.n744 B.n742 163.367
R1467 B.n740 B.n112 163.367
R1468 B.n736 B.n734 163.367
R1469 B.n732 B.n114 163.367
R1470 B.n727 B.n725 163.367
R1471 B.n723 B.n118 163.367
R1472 B.n719 B.n717 163.367
R1473 B.n715 B.n120 163.367
R1474 B.n711 B.n709 163.367
R1475 B.n707 B.n122 163.367
R1476 B.n703 B.n701 163.367
R1477 B.n699 B.n127 163.367
R1478 B.n695 B.n693 163.367
R1479 B.n691 B.n129 163.367
R1480 B.n687 B.n685 163.367
R1481 B.n683 B.n131 163.367
R1482 B.n679 B.n677 163.367
R1483 B.n675 B.n133 163.367
R1484 B.n671 B.n669 163.367
R1485 B.n667 B.n135 163.367
R1486 B.n663 B.n661 163.367
R1487 B.n659 B.n137 163.367
R1488 B.n655 B.n653 163.367
R1489 B.n420 B.n244 103.087
R1490 B.n789 B.n99 103.087
R1491 B.n414 B.n245 71.676
R1492 B.n412 B.n247 71.676
R1493 B.n408 B.n407 71.676
R1494 B.n401 B.n249 71.676
R1495 B.n400 B.n399 71.676
R1496 B.n393 B.n251 71.676
R1497 B.n392 B.n391 71.676
R1498 B.n385 B.n253 71.676
R1499 B.n384 B.n383 71.676
R1500 B.n377 B.n255 71.676
R1501 B.n376 B.n375 71.676
R1502 B.n369 B.n257 71.676
R1503 B.n368 B.n367 71.676
R1504 B.n361 B.n259 71.676
R1505 B.n360 B.n263 71.676
R1506 B.n356 B.n355 71.676
R1507 B.n349 B.n265 71.676
R1508 B.n348 B.n347 71.676
R1509 B.n341 B.n267 71.676
R1510 B.n340 B.n271 71.676
R1511 B.n336 B.n335 71.676
R1512 B.n329 B.n273 71.676
R1513 B.n328 B.n327 71.676
R1514 B.n321 B.n275 71.676
R1515 B.n320 B.n319 71.676
R1516 B.n313 B.n277 71.676
R1517 B.n312 B.n311 71.676
R1518 B.n305 B.n279 71.676
R1519 B.n304 B.n303 71.676
R1520 B.n297 B.n281 71.676
R1521 B.n296 B.n295 71.676
R1522 B.n289 B.n283 71.676
R1523 B.n288 B.n287 71.676
R1524 B.n783 B.n100 71.676
R1525 B.n782 B.n781 71.676
R1526 B.n775 B.n102 71.676
R1527 B.n774 B.n773 71.676
R1528 B.n767 B.n104 71.676
R1529 B.n766 B.n765 71.676
R1530 B.n759 B.n106 71.676
R1531 B.n758 B.n757 71.676
R1532 B.n751 B.n108 71.676
R1533 B.n750 B.n749 71.676
R1534 B.n743 B.n110 71.676
R1535 B.n742 B.n741 71.676
R1536 B.n735 B.n112 71.676
R1537 B.n734 B.n733 71.676
R1538 B.n726 B.n114 71.676
R1539 B.n725 B.n724 71.676
R1540 B.n718 B.n118 71.676
R1541 B.n717 B.n716 71.676
R1542 B.n710 B.n120 71.676
R1543 B.n709 B.n708 71.676
R1544 B.n702 B.n122 71.676
R1545 B.n701 B.n700 71.676
R1546 B.n694 B.n127 71.676
R1547 B.n693 B.n692 71.676
R1548 B.n686 B.n129 71.676
R1549 B.n685 B.n684 71.676
R1550 B.n678 B.n131 71.676
R1551 B.n677 B.n676 71.676
R1552 B.n670 B.n133 71.676
R1553 B.n669 B.n668 71.676
R1554 B.n662 B.n135 71.676
R1555 B.n661 B.n660 71.676
R1556 B.n654 B.n137 71.676
R1557 B.n653 B.n652 71.676
R1558 B.n652 B.n651 71.676
R1559 B.n655 B.n654 71.676
R1560 B.n660 B.n659 71.676
R1561 B.n663 B.n662 71.676
R1562 B.n668 B.n667 71.676
R1563 B.n671 B.n670 71.676
R1564 B.n676 B.n675 71.676
R1565 B.n679 B.n678 71.676
R1566 B.n684 B.n683 71.676
R1567 B.n687 B.n686 71.676
R1568 B.n692 B.n691 71.676
R1569 B.n695 B.n694 71.676
R1570 B.n700 B.n699 71.676
R1571 B.n703 B.n702 71.676
R1572 B.n708 B.n707 71.676
R1573 B.n711 B.n710 71.676
R1574 B.n716 B.n715 71.676
R1575 B.n719 B.n718 71.676
R1576 B.n724 B.n723 71.676
R1577 B.n727 B.n726 71.676
R1578 B.n733 B.n732 71.676
R1579 B.n736 B.n735 71.676
R1580 B.n741 B.n740 71.676
R1581 B.n744 B.n743 71.676
R1582 B.n749 B.n748 71.676
R1583 B.n752 B.n751 71.676
R1584 B.n757 B.n756 71.676
R1585 B.n760 B.n759 71.676
R1586 B.n765 B.n764 71.676
R1587 B.n768 B.n767 71.676
R1588 B.n773 B.n772 71.676
R1589 B.n776 B.n775 71.676
R1590 B.n781 B.n780 71.676
R1591 B.n784 B.n783 71.676
R1592 B.n415 B.n414 71.676
R1593 B.n409 B.n247 71.676
R1594 B.n407 B.n406 71.676
R1595 B.n402 B.n401 71.676
R1596 B.n399 B.n398 71.676
R1597 B.n394 B.n393 71.676
R1598 B.n391 B.n390 71.676
R1599 B.n386 B.n385 71.676
R1600 B.n383 B.n382 71.676
R1601 B.n378 B.n377 71.676
R1602 B.n375 B.n374 71.676
R1603 B.n370 B.n369 71.676
R1604 B.n367 B.n366 71.676
R1605 B.n362 B.n361 71.676
R1606 B.n357 B.n263 71.676
R1607 B.n355 B.n354 71.676
R1608 B.n350 B.n349 71.676
R1609 B.n347 B.n346 71.676
R1610 B.n342 B.n341 71.676
R1611 B.n337 B.n271 71.676
R1612 B.n335 B.n334 71.676
R1613 B.n330 B.n329 71.676
R1614 B.n327 B.n326 71.676
R1615 B.n322 B.n321 71.676
R1616 B.n319 B.n318 71.676
R1617 B.n314 B.n313 71.676
R1618 B.n311 B.n310 71.676
R1619 B.n306 B.n305 71.676
R1620 B.n303 B.n302 71.676
R1621 B.n298 B.n297 71.676
R1622 B.n295 B.n294 71.676
R1623 B.n290 B.n289 71.676
R1624 B.n287 B.n286 71.676
R1625 B.n270 B.n269 59.5399
R1626 B.n262 B.n261 59.5399
R1627 B.n729 B.n116 59.5399
R1628 B.n125 B.n124 59.5399
R1629 B.n420 B.n240 56.991
R1630 B.n426 B.n240 56.991
R1631 B.n426 B.n236 56.991
R1632 B.n432 B.n236 56.991
R1633 B.n432 B.n232 56.991
R1634 B.n439 B.n232 56.991
R1635 B.n439 B.n438 56.991
R1636 B.n445 B.n225 56.991
R1637 B.n451 B.n225 56.991
R1638 B.n451 B.n221 56.991
R1639 B.n457 B.n221 56.991
R1640 B.n457 B.n217 56.991
R1641 B.n463 B.n217 56.991
R1642 B.n463 B.n212 56.991
R1643 B.n469 B.n212 56.991
R1644 B.n469 B.n213 56.991
R1645 B.n475 B.n205 56.991
R1646 B.n481 B.n205 56.991
R1647 B.n481 B.n201 56.991
R1648 B.n487 B.n201 56.991
R1649 B.n487 B.n196 56.991
R1650 B.n493 B.n196 56.991
R1651 B.n493 B.n197 56.991
R1652 B.n499 B.n189 56.991
R1653 B.n505 B.n189 56.991
R1654 B.n505 B.n185 56.991
R1655 B.n511 B.n185 56.991
R1656 B.n511 B.n180 56.991
R1657 B.n517 B.n180 56.991
R1658 B.n517 B.n181 56.991
R1659 B.n523 B.n173 56.991
R1660 B.n529 B.n173 56.991
R1661 B.n529 B.n169 56.991
R1662 B.n535 B.n169 56.991
R1663 B.n535 B.n165 56.991
R1664 B.n541 B.n165 56.991
R1665 B.n547 B.n161 56.991
R1666 B.n547 B.n157 56.991
R1667 B.n553 B.n157 56.991
R1668 B.n553 B.n153 56.991
R1669 B.n559 B.n153 56.991
R1670 B.n559 B.n149 56.991
R1671 B.n565 B.n149 56.991
R1672 B.n572 B.n145 56.991
R1673 B.n572 B.n141 56.991
R1674 B.n578 B.n141 56.991
R1675 B.n578 B.n4 56.991
R1676 B.n895 B.n4 56.991
R1677 B.n895 B.n894 56.991
R1678 B.n894 B.n893 56.991
R1679 B.n893 B.n8 56.991
R1680 B.n887 B.n8 56.991
R1681 B.n887 B.n886 56.991
R1682 B.n885 B.n15 56.991
R1683 B.n879 B.n15 56.991
R1684 B.n879 B.n878 56.991
R1685 B.n878 B.n877 56.991
R1686 B.n877 B.n22 56.991
R1687 B.n871 B.n22 56.991
R1688 B.n871 B.n870 56.991
R1689 B.n869 B.n29 56.991
R1690 B.n863 B.n29 56.991
R1691 B.n863 B.n862 56.991
R1692 B.n862 B.n861 56.991
R1693 B.n861 B.n36 56.991
R1694 B.n855 B.n36 56.991
R1695 B.n854 B.n853 56.991
R1696 B.n853 B.n43 56.991
R1697 B.n847 B.n43 56.991
R1698 B.n847 B.n846 56.991
R1699 B.n846 B.n845 56.991
R1700 B.n845 B.n50 56.991
R1701 B.n839 B.n50 56.991
R1702 B.n838 B.n837 56.991
R1703 B.n837 B.n57 56.991
R1704 B.n831 B.n57 56.991
R1705 B.n831 B.n830 56.991
R1706 B.n830 B.n829 56.991
R1707 B.n829 B.n64 56.991
R1708 B.n823 B.n64 56.991
R1709 B.n822 B.n821 56.991
R1710 B.n821 B.n71 56.991
R1711 B.n815 B.n71 56.991
R1712 B.n815 B.n814 56.991
R1713 B.n814 B.n813 56.991
R1714 B.n813 B.n78 56.991
R1715 B.n807 B.n78 56.991
R1716 B.n807 B.n806 56.991
R1717 B.n806 B.n805 56.991
R1718 B.n799 B.n88 56.991
R1719 B.n799 B.n798 56.991
R1720 B.n798 B.n797 56.991
R1721 B.n797 B.n92 56.991
R1722 B.n791 B.n92 56.991
R1723 B.n791 B.n790 56.991
R1724 B.n790 B.n789 56.991
R1725 B.n213 B.t9 56.1529
R1726 B.t3 B.n822 56.1529
R1727 B.n541 B.t5 52.8005
R1728 B.t4 B.n869 52.8005
R1729 B.n269 B.n268 50.4247
R1730 B.n261 B.n260 50.4247
R1731 B.n116 B.n115 50.4247
R1732 B.n124 B.n123 50.4247
R1733 B.n445 B.t11 49.4481
R1734 B.n805 B.t15 49.4481
R1735 B.n523 B.t6 41.0672
R1736 B.n855 B.t2 41.0672
R1737 B.n197 B.t8 36.0386
R1738 B.t1 B.n838 36.0386
R1739 B.n787 B.n786 34.4981
R1740 B.n650 B.n649 34.4981
R1741 B.n422 B.n242 34.4981
R1742 B.n418 B.n417 34.4981
R1743 B.n565 B.t7 32.6862
R1744 B.t0 B.n885 32.6862
R1745 B.t7 B.n145 24.3053
R1746 B.n886 B.t0 24.3053
R1747 B.n499 B.t8 20.9529
R1748 B.n839 B.t1 20.9529
R1749 B B.n897 18.0485
R1750 B.n181 B.t6 15.9243
R1751 B.t2 B.n854 15.9243
R1752 B.n786 B.n785 10.6151
R1753 B.n785 B.n101 10.6151
R1754 B.n779 B.n101 10.6151
R1755 B.n779 B.n778 10.6151
R1756 B.n778 B.n777 10.6151
R1757 B.n777 B.n103 10.6151
R1758 B.n771 B.n103 10.6151
R1759 B.n771 B.n770 10.6151
R1760 B.n770 B.n769 10.6151
R1761 B.n769 B.n105 10.6151
R1762 B.n763 B.n105 10.6151
R1763 B.n763 B.n762 10.6151
R1764 B.n762 B.n761 10.6151
R1765 B.n761 B.n107 10.6151
R1766 B.n755 B.n107 10.6151
R1767 B.n755 B.n754 10.6151
R1768 B.n754 B.n753 10.6151
R1769 B.n753 B.n109 10.6151
R1770 B.n747 B.n109 10.6151
R1771 B.n747 B.n746 10.6151
R1772 B.n746 B.n745 10.6151
R1773 B.n745 B.n111 10.6151
R1774 B.n739 B.n111 10.6151
R1775 B.n739 B.n738 10.6151
R1776 B.n738 B.n737 10.6151
R1777 B.n737 B.n113 10.6151
R1778 B.n731 B.n113 10.6151
R1779 B.n731 B.n730 10.6151
R1780 B.n728 B.n117 10.6151
R1781 B.n722 B.n117 10.6151
R1782 B.n722 B.n721 10.6151
R1783 B.n721 B.n720 10.6151
R1784 B.n720 B.n119 10.6151
R1785 B.n714 B.n119 10.6151
R1786 B.n714 B.n713 10.6151
R1787 B.n713 B.n712 10.6151
R1788 B.n712 B.n121 10.6151
R1789 B.n706 B.n705 10.6151
R1790 B.n705 B.n704 10.6151
R1791 B.n704 B.n126 10.6151
R1792 B.n698 B.n126 10.6151
R1793 B.n698 B.n697 10.6151
R1794 B.n697 B.n696 10.6151
R1795 B.n696 B.n128 10.6151
R1796 B.n690 B.n128 10.6151
R1797 B.n690 B.n689 10.6151
R1798 B.n689 B.n688 10.6151
R1799 B.n688 B.n130 10.6151
R1800 B.n682 B.n130 10.6151
R1801 B.n682 B.n681 10.6151
R1802 B.n681 B.n680 10.6151
R1803 B.n680 B.n132 10.6151
R1804 B.n674 B.n132 10.6151
R1805 B.n674 B.n673 10.6151
R1806 B.n673 B.n672 10.6151
R1807 B.n672 B.n134 10.6151
R1808 B.n666 B.n134 10.6151
R1809 B.n666 B.n665 10.6151
R1810 B.n665 B.n664 10.6151
R1811 B.n664 B.n136 10.6151
R1812 B.n658 B.n136 10.6151
R1813 B.n658 B.n657 10.6151
R1814 B.n657 B.n656 10.6151
R1815 B.n656 B.n138 10.6151
R1816 B.n650 B.n138 10.6151
R1817 B.n423 B.n422 10.6151
R1818 B.n424 B.n423 10.6151
R1819 B.n424 B.n234 10.6151
R1820 B.n434 B.n234 10.6151
R1821 B.n435 B.n434 10.6151
R1822 B.n436 B.n435 10.6151
R1823 B.n436 B.n227 10.6151
R1824 B.n447 B.n227 10.6151
R1825 B.n448 B.n447 10.6151
R1826 B.n449 B.n448 10.6151
R1827 B.n449 B.n219 10.6151
R1828 B.n459 B.n219 10.6151
R1829 B.n460 B.n459 10.6151
R1830 B.n461 B.n460 10.6151
R1831 B.n461 B.n210 10.6151
R1832 B.n471 B.n210 10.6151
R1833 B.n472 B.n471 10.6151
R1834 B.n473 B.n472 10.6151
R1835 B.n473 B.n203 10.6151
R1836 B.n483 B.n203 10.6151
R1837 B.n484 B.n483 10.6151
R1838 B.n485 B.n484 10.6151
R1839 B.n485 B.n194 10.6151
R1840 B.n495 B.n194 10.6151
R1841 B.n496 B.n495 10.6151
R1842 B.n497 B.n496 10.6151
R1843 B.n497 B.n187 10.6151
R1844 B.n507 B.n187 10.6151
R1845 B.n508 B.n507 10.6151
R1846 B.n509 B.n508 10.6151
R1847 B.n509 B.n178 10.6151
R1848 B.n519 B.n178 10.6151
R1849 B.n520 B.n519 10.6151
R1850 B.n521 B.n520 10.6151
R1851 B.n521 B.n171 10.6151
R1852 B.n531 B.n171 10.6151
R1853 B.n532 B.n531 10.6151
R1854 B.n533 B.n532 10.6151
R1855 B.n533 B.n163 10.6151
R1856 B.n543 B.n163 10.6151
R1857 B.n544 B.n543 10.6151
R1858 B.n545 B.n544 10.6151
R1859 B.n545 B.n155 10.6151
R1860 B.n555 B.n155 10.6151
R1861 B.n556 B.n555 10.6151
R1862 B.n557 B.n556 10.6151
R1863 B.n557 B.n147 10.6151
R1864 B.n567 B.n147 10.6151
R1865 B.n568 B.n567 10.6151
R1866 B.n570 B.n568 10.6151
R1867 B.n570 B.n569 10.6151
R1868 B.n569 B.n139 10.6151
R1869 B.n581 B.n139 10.6151
R1870 B.n582 B.n581 10.6151
R1871 B.n583 B.n582 10.6151
R1872 B.n584 B.n583 10.6151
R1873 B.n586 B.n584 10.6151
R1874 B.n587 B.n586 10.6151
R1875 B.n588 B.n587 10.6151
R1876 B.n589 B.n588 10.6151
R1877 B.n591 B.n589 10.6151
R1878 B.n592 B.n591 10.6151
R1879 B.n593 B.n592 10.6151
R1880 B.n594 B.n593 10.6151
R1881 B.n596 B.n594 10.6151
R1882 B.n597 B.n596 10.6151
R1883 B.n598 B.n597 10.6151
R1884 B.n599 B.n598 10.6151
R1885 B.n601 B.n599 10.6151
R1886 B.n602 B.n601 10.6151
R1887 B.n603 B.n602 10.6151
R1888 B.n604 B.n603 10.6151
R1889 B.n606 B.n604 10.6151
R1890 B.n607 B.n606 10.6151
R1891 B.n608 B.n607 10.6151
R1892 B.n609 B.n608 10.6151
R1893 B.n611 B.n609 10.6151
R1894 B.n612 B.n611 10.6151
R1895 B.n613 B.n612 10.6151
R1896 B.n614 B.n613 10.6151
R1897 B.n616 B.n614 10.6151
R1898 B.n617 B.n616 10.6151
R1899 B.n618 B.n617 10.6151
R1900 B.n619 B.n618 10.6151
R1901 B.n621 B.n619 10.6151
R1902 B.n622 B.n621 10.6151
R1903 B.n623 B.n622 10.6151
R1904 B.n624 B.n623 10.6151
R1905 B.n626 B.n624 10.6151
R1906 B.n627 B.n626 10.6151
R1907 B.n628 B.n627 10.6151
R1908 B.n629 B.n628 10.6151
R1909 B.n631 B.n629 10.6151
R1910 B.n632 B.n631 10.6151
R1911 B.n633 B.n632 10.6151
R1912 B.n634 B.n633 10.6151
R1913 B.n636 B.n634 10.6151
R1914 B.n637 B.n636 10.6151
R1915 B.n638 B.n637 10.6151
R1916 B.n639 B.n638 10.6151
R1917 B.n641 B.n639 10.6151
R1918 B.n642 B.n641 10.6151
R1919 B.n643 B.n642 10.6151
R1920 B.n644 B.n643 10.6151
R1921 B.n646 B.n644 10.6151
R1922 B.n647 B.n646 10.6151
R1923 B.n648 B.n647 10.6151
R1924 B.n649 B.n648 10.6151
R1925 B.n417 B.n416 10.6151
R1926 B.n416 B.n246 10.6151
R1927 B.n411 B.n246 10.6151
R1928 B.n411 B.n410 10.6151
R1929 B.n410 B.n248 10.6151
R1930 B.n405 B.n248 10.6151
R1931 B.n405 B.n404 10.6151
R1932 B.n404 B.n403 10.6151
R1933 B.n403 B.n250 10.6151
R1934 B.n397 B.n250 10.6151
R1935 B.n397 B.n396 10.6151
R1936 B.n396 B.n395 10.6151
R1937 B.n395 B.n252 10.6151
R1938 B.n389 B.n252 10.6151
R1939 B.n389 B.n388 10.6151
R1940 B.n388 B.n387 10.6151
R1941 B.n387 B.n254 10.6151
R1942 B.n381 B.n254 10.6151
R1943 B.n381 B.n380 10.6151
R1944 B.n380 B.n379 10.6151
R1945 B.n379 B.n256 10.6151
R1946 B.n373 B.n256 10.6151
R1947 B.n373 B.n372 10.6151
R1948 B.n372 B.n371 10.6151
R1949 B.n371 B.n258 10.6151
R1950 B.n365 B.n258 10.6151
R1951 B.n365 B.n364 10.6151
R1952 B.n364 B.n363 10.6151
R1953 B.n359 B.n358 10.6151
R1954 B.n358 B.n264 10.6151
R1955 B.n353 B.n264 10.6151
R1956 B.n353 B.n352 10.6151
R1957 B.n352 B.n351 10.6151
R1958 B.n351 B.n266 10.6151
R1959 B.n345 B.n266 10.6151
R1960 B.n345 B.n344 10.6151
R1961 B.n344 B.n343 10.6151
R1962 B.n339 B.n338 10.6151
R1963 B.n338 B.n272 10.6151
R1964 B.n333 B.n272 10.6151
R1965 B.n333 B.n332 10.6151
R1966 B.n332 B.n331 10.6151
R1967 B.n331 B.n274 10.6151
R1968 B.n325 B.n274 10.6151
R1969 B.n325 B.n324 10.6151
R1970 B.n324 B.n323 10.6151
R1971 B.n323 B.n276 10.6151
R1972 B.n317 B.n276 10.6151
R1973 B.n317 B.n316 10.6151
R1974 B.n316 B.n315 10.6151
R1975 B.n315 B.n278 10.6151
R1976 B.n309 B.n278 10.6151
R1977 B.n309 B.n308 10.6151
R1978 B.n308 B.n307 10.6151
R1979 B.n307 B.n280 10.6151
R1980 B.n301 B.n280 10.6151
R1981 B.n301 B.n300 10.6151
R1982 B.n300 B.n299 10.6151
R1983 B.n299 B.n282 10.6151
R1984 B.n293 B.n282 10.6151
R1985 B.n293 B.n292 10.6151
R1986 B.n292 B.n291 10.6151
R1987 B.n291 B.n284 10.6151
R1988 B.n285 B.n284 10.6151
R1989 B.n285 B.n242 10.6151
R1990 B.n418 B.n238 10.6151
R1991 B.n428 B.n238 10.6151
R1992 B.n429 B.n428 10.6151
R1993 B.n430 B.n429 10.6151
R1994 B.n430 B.n230 10.6151
R1995 B.n441 B.n230 10.6151
R1996 B.n442 B.n441 10.6151
R1997 B.n443 B.n442 10.6151
R1998 B.n443 B.n223 10.6151
R1999 B.n453 B.n223 10.6151
R2000 B.n454 B.n453 10.6151
R2001 B.n455 B.n454 10.6151
R2002 B.n455 B.n215 10.6151
R2003 B.n465 B.n215 10.6151
R2004 B.n466 B.n465 10.6151
R2005 B.n467 B.n466 10.6151
R2006 B.n467 B.n207 10.6151
R2007 B.n477 B.n207 10.6151
R2008 B.n478 B.n477 10.6151
R2009 B.n479 B.n478 10.6151
R2010 B.n479 B.n199 10.6151
R2011 B.n489 B.n199 10.6151
R2012 B.n490 B.n489 10.6151
R2013 B.n491 B.n490 10.6151
R2014 B.n491 B.n191 10.6151
R2015 B.n501 B.n191 10.6151
R2016 B.n502 B.n501 10.6151
R2017 B.n503 B.n502 10.6151
R2018 B.n503 B.n183 10.6151
R2019 B.n513 B.n183 10.6151
R2020 B.n514 B.n513 10.6151
R2021 B.n515 B.n514 10.6151
R2022 B.n515 B.n175 10.6151
R2023 B.n525 B.n175 10.6151
R2024 B.n526 B.n525 10.6151
R2025 B.n527 B.n526 10.6151
R2026 B.n527 B.n167 10.6151
R2027 B.n537 B.n167 10.6151
R2028 B.n538 B.n537 10.6151
R2029 B.n539 B.n538 10.6151
R2030 B.n539 B.n159 10.6151
R2031 B.n549 B.n159 10.6151
R2032 B.n550 B.n549 10.6151
R2033 B.n551 B.n550 10.6151
R2034 B.n551 B.n151 10.6151
R2035 B.n561 B.n151 10.6151
R2036 B.n562 B.n561 10.6151
R2037 B.n563 B.n562 10.6151
R2038 B.n563 B.n143 10.6151
R2039 B.n574 B.n143 10.6151
R2040 B.n575 B.n574 10.6151
R2041 B.n576 B.n575 10.6151
R2042 B.n576 B.n0 10.6151
R2043 B.n891 B.n1 10.6151
R2044 B.n891 B.n890 10.6151
R2045 B.n890 B.n889 10.6151
R2046 B.n889 B.n10 10.6151
R2047 B.n883 B.n10 10.6151
R2048 B.n883 B.n882 10.6151
R2049 B.n882 B.n881 10.6151
R2050 B.n881 B.n17 10.6151
R2051 B.n875 B.n17 10.6151
R2052 B.n875 B.n874 10.6151
R2053 B.n874 B.n873 10.6151
R2054 B.n873 B.n24 10.6151
R2055 B.n867 B.n24 10.6151
R2056 B.n867 B.n866 10.6151
R2057 B.n866 B.n865 10.6151
R2058 B.n865 B.n31 10.6151
R2059 B.n859 B.n31 10.6151
R2060 B.n859 B.n858 10.6151
R2061 B.n858 B.n857 10.6151
R2062 B.n857 B.n38 10.6151
R2063 B.n851 B.n38 10.6151
R2064 B.n851 B.n850 10.6151
R2065 B.n850 B.n849 10.6151
R2066 B.n849 B.n45 10.6151
R2067 B.n843 B.n45 10.6151
R2068 B.n843 B.n842 10.6151
R2069 B.n842 B.n841 10.6151
R2070 B.n841 B.n52 10.6151
R2071 B.n835 B.n52 10.6151
R2072 B.n835 B.n834 10.6151
R2073 B.n834 B.n833 10.6151
R2074 B.n833 B.n59 10.6151
R2075 B.n827 B.n59 10.6151
R2076 B.n827 B.n826 10.6151
R2077 B.n826 B.n825 10.6151
R2078 B.n825 B.n66 10.6151
R2079 B.n819 B.n66 10.6151
R2080 B.n819 B.n818 10.6151
R2081 B.n818 B.n817 10.6151
R2082 B.n817 B.n73 10.6151
R2083 B.n811 B.n73 10.6151
R2084 B.n811 B.n810 10.6151
R2085 B.n810 B.n809 10.6151
R2086 B.n809 B.n80 10.6151
R2087 B.n803 B.n80 10.6151
R2088 B.n803 B.n802 10.6151
R2089 B.n802 B.n801 10.6151
R2090 B.n801 B.n86 10.6151
R2091 B.n795 B.n86 10.6151
R2092 B.n795 B.n794 10.6151
R2093 B.n794 B.n793 10.6151
R2094 B.n793 B.n94 10.6151
R2095 B.n787 B.n94 10.6151
R2096 B.n730 B.n729 9.36635
R2097 B.n706 B.n125 9.36635
R2098 B.n363 B.n262 9.36635
R2099 B.n339 B.n270 9.36635
R2100 B.n438 B.t11 7.54336
R2101 B.n88 B.t15 7.54336
R2102 B.t5 B.n161 4.19098
R2103 B.n870 B.t4 4.19098
R2104 B.n897 B.n0 2.81026
R2105 B.n897 B.n1 2.81026
R2106 B.n729 B.n728 1.24928
R2107 B.n125 B.n121 1.24928
R2108 B.n359 B.n262 1.24928
R2109 B.n343 B.n270 1.24928
R2110 B.n475 B.t9 0.838595
R2111 B.n823 B.t3 0.838595
R2112 VP.n22 VP.n21 161.3
R2113 VP.n23 VP.n18 161.3
R2114 VP.n25 VP.n24 161.3
R2115 VP.n26 VP.n17 161.3
R2116 VP.n28 VP.n27 161.3
R2117 VP.n29 VP.n16 161.3
R2118 VP.n31 VP.n30 161.3
R2119 VP.n32 VP.n15 161.3
R2120 VP.n34 VP.n33 161.3
R2121 VP.n35 VP.n14 161.3
R2122 VP.n37 VP.n36 161.3
R2123 VP.n39 VP.n13 161.3
R2124 VP.n41 VP.n40 161.3
R2125 VP.n42 VP.n12 161.3
R2126 VP.n44 VP.n43 161.3
R2127 VP.n45 VP.n11 161.3
R2128 VP.n82 VP.n0 161.3
R2129 VP.n81 VP.n80 161.3
R2130 VP.n79 VP.n1 161.3
R2131 VP.n78 VP.n77 161.3
R2132 VP.n76 VP.n2 161.3
R2133 VP.n74 VP.n73 161.3
R2134 VP.n72 VP.n3 161.3
R2135 VP.n71 VP.n70 161.3
R2136 VP.n69 VP.n4 161.3
R2137 VP.n68 VP.n67 161.3
R2138 VP.n66 VP.n5 161.3
R2139 VP.n65 VP.n64 161.3
R2140 VP.n63 VP.n6 161.3
R2141 VP.n62 VP.n61 161.3
R2142 VP.n60 VP.n7 161.3
R2143 VP.n59 VP.n58 161.3
R2144 VP.n56 VP.n8 161.3
R2145 VP.n55 VP.n54 161.3
R2146 VP.n53 VP.n9 161.3
R2147 VP.n52 VP.n51 161.3
R2148 VP.n50 VP.n10 161.3
R2149 VP.n19 VP.t7 114.216
R2150 VP.n49 VP.n48 100.969
R2151 VP.n84 VP.n83 100.969
R2152 VP.n47 VP.n46 100.969
R2153 VP.n5 VP.t0 83.3419
R2154 VP.n49 VP.t3 83.3419
R2155 VP.n57 VP.t4 83.3419
R2156 VP.n75 VP.t2 83.3419
R2157 VP.n83 VP.t1 83.3419
R2158 VP.n16 VP.t8 83.3419
R2159 VP.n46 VP.t5 83.3419
R2160 VP.n38 VP.t6 83.3419
R2161 VP.n20 VP.t9 83.3419
R2162 VP.n20 VP.n19 67.1934
R2163 VP.n63 VP.n62 56.5193
R2164 VP.n70 VP.n69 56.5193
R2165 VP.n33 VP.n32 56.5193
R2166 VP.n26 VP.n25 56.5193
R2167 VP.n55 VP.n9 50.2061
R2168 VP.n77 VP.n1 50.2061
R2169 VP.n40 VP.n12 50.2061
R2170 VP.n48 VP.n47 48.1132
R2171 VP.n51 VP.n9 30.7807
R2172 VP.n81 VP.n1 30.7807
R2173 VP.n44 VP.n12 30.7807
R2174 VP.n51 VP.n50 24.4675
R2175 VP.n56 VP.n55 24.4675
R2176 VP.n58 VP.n7 24.4675
R2177 VP.n62 VP.n7 24.4675
R2178 VP.n64 VP.n63 24.4675
R2179 VP.n64 VP.n5 24.4675
R2180 VP.n68 VP.n5 24.4675
R2181 VP.n69 VP.n68 24.4675
R2182 VP.n70 VP.n3 24.4675
R2183 VP.n74 VP.n3 24.4675
R2184 VP.n77 VP.n76 24.4675
R2185 VP.n82 VP.n81 24.4675
R2186 VP.n45 VP.n44 24.4675
R2187 VP.n33 VP.n14 24.4675
R2188 VP.n37 VP.n14 24.4675
R2189 VP.n40 VP.n39 24.4675
R2190 VP.n27 VP.n26 24.4675
R2191 VP.n27 VP.n16 24.4675
R2192 VP.n31 VP.n16 24.4675
R2193 VP.n32 VP.n31 24.4675
R2194 VP.n21 VP.n18 24.4675
R2195 VP.n25 VP.n18 24.4675
R2196 VP.n57 VP.n56 19.5741
R2197 VP.n76 VP.n75 19.5741
R2198 VP.n39 VP.n38 19.5741
R2199 VP.n22 VP.n19 10.026
R2200 VP.n50 VP.n49 9.7873
R2201 VP.n83 VP.n82 9.7873
R2202 VP.n46 VP.n45 9.7873
R2203 VP.n58 VP.n57 4.8939
R2204 VP.n75 VP.n74 4.8939
R2205 VP.n38 VP.n37 4.8939
R2206 VP.n21 VP.n20 4.8939
R2207 VP.n47 VP.n11 0.278367
R2208 VP.n48 VP.n10 0.278367
R2209 VP.n84 VP.n0 0.278367
R2210 VP.n23 VP.n22 0.189894
R2211 VP.n24 VP.n23 0.189894
R2212 VP.n24 VP.n17 0.189894
R2213 VP.n28 VP.n17 0.189894
R2214 VP.n29 VP.n28 0.189894
R2215 VP.n30 VP.n29 0.189894
R2216 VP.n30 VP.n15 0.189894
R2217 VP.n34 VP.n15 0.189894
R2218 VP.n35 VP.n34 0.189894
R2219 VP.n36 VP.n35 0.189894
R2220 VP.n36 VP.n13 0.189894
R2221 VP.n41 VP.n13 0.189894
R2222 VP.n42 VP.n41 0.189894
R2223 VP.n43 VP.n42 0.189894
R2224 VP.n43 VP.n11 0.189894
R2225 VP.n52 VP.n10 0.189894
R2226 VP.n53 VP.n52 0.189894
R2227 VP.n54 VP.n53 0.189894
R2228 VP.n54 VP.n8 0.189894
R2229 VP.n59 VP.n8 0.189894
R2230 VP.n60 VP.n59 0.189894
R2231 VP.n61 VP.n60 0.189894
R2232 VP.n61 VP.n6 0.189894
R2233 VP.n65 VP.n6 0.189894
R2234 VP.n66 VP.n65 0.189894
R2235 VP.n67 VP.n66 0.189894
R2236 VP.n67 VP.n4 0.189894
R2237 VP.n71 VP.n4 0.189894
R2238 VP.n72 VP.n71 0.189894
R2239 VP.n73 VP.n72 0.189894
R2240 VP.n73 VP.n2 0.189894
R2241 VP.n78 VP.n2 0.189894
R2242 VP.n79 VP.n78 0.189894
R2243 VP.n80 VP.n79 0.189894
R2244 VP.n80 VP.n0 0.189894
R2245 VP VP.n84 0.153454
R2246 VDD1.n36 VDD1.n0 289.615
R2247 VDD1.n79 VDD1.n43 289.615
R2248 VDD1.n37 VDD1.n36 185
R2249 VDD1.n35 VDD1.n2 185
R2250 VDD1.n34 VDD1.n33 185
R2251 VDD1.n5 VDD1.n3 185
R2252 VDD1.n28 VDD1.n27 185
R2253 VDD1.n26 VDD1.n25 185
R2254 VDD1.n9 VDD1.n8 185
R2255 VDD1.n20 VDD1.n19 185
R2256 VDD1.n18 VDD1.n17 185
R2257 VDD1.n13 VDD1.n12 185
R2258 VDD1.n55 VDD1.n54 185
R2259 VDD1.n60 VDD1.n59 185
R2260 VDD1.n62 VDD1.n61 185
R2261 VDD1.n51 VDD1.n50 185
R2262 VDD1.n68 VDD1.n67 185
R2263 VDD1.n70 VDD1.n69 185
R2264 VDD1.n47 VDD1.n46 185
R2265 VDD1.n77 VDD1.n76 185
R2266 VDD1.n78 VDD1.n45 185
R2267 VDD1.n80 VDD1.n79 185
R2268 VDD1.n14 VDD1.t2 149.524
R2269 VDD1.n56 VDD1.t6 149.524
R2270 VDD1.n36 VDD1.n35 104.615
R2271 VDD1.n35 VDD1.n34 104.615
R2272 VDD1.n34 VDD1.n3 104.615
R2273 VDD1.n27 VDD1.n3 104.615
R2274 VDD1.n27 VDD1.n26 104.615
R2275 VDD1.n26 VDD1.n8 104.615
R2276 VDD1.n19 VDD1.n8 104.615
R2277 VDD1.n19 VDD1.n18 104.615
R2278 VDD1.n18 VDD1.n12 104.615
R2279 VDD1.n60 VDD1.n54 104.615
R2280 VDD1.n61 VDD1.n60 104.615
R2281 VDD1.n61 VDD1.n50 104.615
R2282 VDD1.n68 VDD1.n50 104.615
R2283 VDD1.n69 VDD1.n68 104.615
R2284 VDD1.n69 VDD1.n46 104.615
R2285 VDD1.n77 VDD1.n46 104.615
R2286 VDD1.n78 VDD1.n77 104.615
R2287 VDD1.n79 VDD1.n78 104.615
R2288 VDD1.n87 VDD1.n86 66.5732
R2289 VDD1.n42 VDD1.n41 64.9477
R2290 VDD1.n89 VDD1.n88 64.9475
R2291 VDD1.n85 VDD1.n84 64.9475
R2292 VDD1.t2 VDD1.n12 52.3082
R2293 VDD1.t6 VDD1.n54 52.3082
R2294 VDD1.n42 VDD1.n40 52.0752
R2295 VDD1.n85 VDD1.n83 52.0752
R2296 VDD1.n89 VDD1.n87 42.8328
R2297 VDD1.n37 VDD1.n2 13.1884
R2298 VDD1.n80 VDD1.n45 13.1884
R2299 VDD1.n38 VDD1.n0 12.8005
R2300 VDD1.n33 VDD1.n4 12.8005
R2301 VDD1.n76 VDD1.n75 12.8005
R2302 VDD1.n81 VDD1.n43 12.8005
R2303 VDD1.n32 VDD1.n5 12.0247
R2304 VDD1.n74 VDD1.n47 12.0247
R2305 VDD1.n29 VDD1.n28 11.249
R2306 VDD1.n71 VDD1.n70 11.249
R2307 VDD1.n25 VDD1.n7 10.4732
R2308 VDD1.n67 VDD1.n49 10.4732
R2309 VDD1.n14 VDD1.n13 10.2747
R2310 VDD1.n56 VDD1.n55 10.2747
R2311 VDD1.n24 VDD1.n9 9.69747
R2312 VDD1.n66 VDD1.n51 9.69747
R2313 VDD1.n40 VDD1.n39 9.45567
R2314 VDD1.n83 VDD1.n82 9.45567
R2315 VDD1.n16 VDD1.n15 9.3005
R2316 VDD1.n11 VDD1.n10 9.3005
R2317 VDD1.n22 VDD1.n21 9.3005
R2318 VDD1.n24 VDD1.n23 9.3005
R2319 VDD1.n7 VDD1.n6 9.3005
R2320 VDD1.n30 VDD1.n29 9.3005
R2321 VDD1.n32 VDD1.n31 9.3005
R2322 VDD1.n4 VDD1.n1 9.3005
R2323 VDD1.n39 VDD1.n38 9.3005
R2324 VDD1.n82 VDD1.n81 9.3005
R2325 VDD1.n58 VDD1.n57 9.3005
R2326 VDD1.n53 VDD1.n52 9.3005
R2327 VDD1.n64 VDD1.n63 9.3005
R2328 VDD1.n66 VDD1.n65 9.3005
R2329 VDD1.n49 VDD1.n48 9.3005
R2330 VDD1.n72 VDD1.n71 9.3005
R2331 VDD1.n74 VDD1.n73 9.3005
R2332 VDD1.n75 VDD1.n44 9.3005
R2333 VDD1.n21 VDD1.n20 8.92171
R2334 VDD1.n63 VDD1.n62 8.92171
R2335 VDD1.n17 VDD1.n11 8.14595
R2336 VDD1.n59 VDD1.n53 8.14595
R2337 VDD1.n16 VDD1.n13 7.3702
R2338 VDD1.n58 VDD1.n55 7.3702
R2339 VDD1.n17 VDD1.n16 5.81868
R2340 VDD1.n59 VDD1.n58 5.81868
R2341 VDD1.n20 VDD1.n11 5.04292
R2342 VDD1.n62 VDD1.n53 5.04292
R2343 VDD1.n21 VDD1.n9 4.26717
R2344 VDD1.n63 VDD1.n51 4.26717
R2345 VDD1.n25 VDD1.n24 3.49141
R2346 VDD1.n67 VDD1.n66 3.49141
R2347 VDD1.n15 VDD1.n14 2.84304
R2348 VDD1.n57 VDD1.n56 2.84304
R2349 VDD1.n28 VDD1.n7 2.71565
R2350 VDD1.n70 VDD1.n49 2.71565
R2351 VDD1.n88 VDD1.t3 2.52279
R2352 VDD1.n88 VDD1.t4 2.52279
R2353 VDD1.n41 VDD1.t0 2.52279
R2354 VDD1.n41 VDD1.t1 2.52279
R2355 VDD1.n86 VDD1.t7 2.52279
R2356 VDD1.n86 VDD1.t8 2.52279
R2357 VDD1.n84 VDD1.t5 2.52279
R2358 VDD1.n84 VDD1.t9 2.52279
R2359 VDD1.n29 VDD1.n5 1.93989
R2360 VDD1.n71 VDD1.n47 1.93989
R2361 VDD1 VDD1.n89 1.62334
R2362 VDD1.n40 VDD1.n0 1.16414
R2363 VDD1.n33 VDD1.n32 1.16414
R2364 VDD1.n76 VDD1.n74 1.16414
R2365 VDD1.n83 VDD1.n43 1.16414
R2366 VDD1 VDD1.n42 0.619035
R2367 VDD1.n87 VDD1.n85 0.505499
R2368 VDD1.n38 VDD1.n37 0.388379
R2369 VDD1.n4 VDD1.n2 0.388379
R2370 VDD1.n75 VDD1.n45 0.388379
R2371 VDD1.n81 VDD1.n80 0.388379
R2372 VDD1.n39 VDD1.n1 0.155672
R2373 VDD1.n31 VDD1.n1 0.155672
R2374 VDD1.n31 VDD1.n30 0.155672
R2375 VDD1.n30 VDD1.n6 0.155672
R2376 VDD1.n23 VDD1.n6 0.155672
R2377 VDD1.n23 VDD1.n22 0.155672
R2378 VDD1.n22 VDD1.n10 0.155672
R2379 VDD1.n15 VDD1.n10 0.155672
R2380 VDD1.n57 VDD1.n52 0.155672
R2381 VDD1.n64 VDD1.n52 0.155672
R2382 VDD1.n65 VDD1.n64 0.155672
R2383 VDD1.n65 VDD1.n48 0.155672
R2384 VDD1.n72 VDD1.n48 0.155672
R2385 VDD1.n73 VDD1.n72 0.155672
R2386 VDD1.n73 VDD1.n44 0.155672
R2387 VDD1.n82 VDD1.n44 0.155672
C0 VN VDD2 6.95152f
C1 VN VP 7.14762f
C2 VTAIL VDD2 8.37354f
C3 VTAIL VP 7.64944f
C4 VDD1 VDD2 1.95934f
C5 VDD1 VP 7.33698f
C6 VN VTAIL 7.6352f
C7 VDD2 VP 0.54116f
C8 VN VDD1 0.152635f
C9 VTAIL VDD1 8.3241f
C10 VDD2 B 6.053424f
C11 VDD1 B 6.050349f
C12 VTAIL B 6.319111f
C13 VN B 16.25001f
C14 VP B 14.805311f
C15 VDD1.n0 B 0.028885f
C16 VDD1.n1 B 0.022612f
C17 VDD1.n2 B 0.012508f
C18 VDD1.n3 B 0.02872f
C19 VDD1.n4 B 0.012151f
C20 VDD1.n5 B 0.012865f
C21 VDD1.n6 B 0.022612f
C22 VDD1.n7 B 0.012151f
C23 VDD1.n8 B 0.02872f
C24 VDD1.n9 B 0.012865f
C25 VDD1.n10 B 0.022612f
C26 VDD1.n11 B 0.012151f
C27 VDD1.n12 B 0.02154f
C28 VDD1.n13 B 0.020303f
C29 VDD1.t2 B 0.048013f
C30 VDD1.n14 B 0.127025f
C31 VDD1.n15 B 0.723315f
C32 VDD1.n16 B 0.012151f
C33 VDD1.n17 B 0.012865f
C34 VDD1.n18 B 0.02872f
C35 VDD1.n19 B 0.02872f
C36 VDD1.n20 B 0.012865f
C37 VDD1.n21 B 0.012151f
C38 VDD1.n22 B 0.022612f
C39 VDD1.n23 B 0.022612f
C40 VDD1.n24 B 0.012151f
C41 VDD1.n25 B 0.012865f
C42 VDD1.n26 B 0.02872f
C43 VDD1.n27 B 0.02872f
C44 VDD1.n28 B 0.012865f
C45 VDD1.n29 B 0.012151f
C46 VDD1.n30 B 0.022612f
C47 VDD1.n31 B 0.022612f
C48 VDD1.n32 B 0.012151f
C49 VDD1.n33 B 0.012865f
C50 VDD1.n34 B 0.02872f
C51 VDD1.n35 B 0.02872f
C52 VDD1.n36 B 0.057048f
C53 VDD1.n37 B 0.012508f
C54 VDD1.n38 B 0.012151f
C55 VDD1.n39 B 0.053811f
C56 VDD1.n40 B 0.055983f
C57 VDD1.t0 B 0.140269f
C58 VDD1.t1 B 0.140269f
C59 VDD1.n41 B 1.2125f
C60 VDD1.n42 B 0.586889f
C61 VDD1.n43 B 0.028885f
C62 VDD1.n44 B 0.022612f
C63 VDD1.n45 B 0.012508f
C64 VDD1.n46 B 0.02872f
C65 VDD1.n47 B 0.012865f
C66 VDD1.n48 B 0.022612f
C67 VDD1.n49 B 0.012151f
C68 VDD1.n50 B 0.02872f
C69 VDD1.n51 B 0.012865f
C70 VDD1.n52 B 0.022612f
C71 VDD1.n53 B 0.012151f
C72 VDD1.n54 B 0.02154f
C73 VDD1.n55 B 0.020303f
C74 VDD1.t6 B 0.048013f
C75 VDD1.n56 B 0.127025f
C76 VDD1.n57 B 0.723315f
C77 VDD1.n58 B 0.012151f
C78 VDD1.n59 B 0.012865f
C79 VDD1.n60 B 0.02872f
C80 VDD1.n61 B 0.02872f
C81 VDD1.n62 B 0.012865f
C82 VDD1.n63 B 0.012151f
C83 VDD1.n64 B 0.022612f
C84 VDD1.n65 B 0.022612f
C85 VDD1.n66 B 0.012151f
C86 VDD1.n67 B 0.012865f
C87 VDD1.n68 B 0.02872f
C88 VDD1.n69 B 0.02872f
C89 VDD1.n70 B 0.012865f
C90 VDD1.n71 B 0.012151f
C91 VDD1.n72 B 0.022612f
C92 VDD1.n73 B 0.022612f
C93 VDD1.n74 B 0.012151f
C94 VDD1.n75 B 0.012151f
C95 VDD1.n76 B 0.012865f
C96 VDD1.n77 B 0.02872f
C97 VDD1.n78 B 0.02872f
C98 VDD1.n79 B 0.057048f
C99 VDD1.n80 B 0.012508f
C100 VDD1.n81 B 0.012151f
C101 VDD1.n82 B 0.053811f
C102 VDD1.n83 B 0.055983f
C103 VDD1.t5 B 0.140269f
C104 VDD1.t9 B 0.140269f
C105 VDD1.n84 B 1.21249f
C106 VDD1.n85 B 0.57966f
C107 VDD1.t7 B 0.140269f
C108 VDD1.t8 B 0.140269f
C109 VDD1.n86 B 1.22399f
C110 VDD1.n87 B 2.33931f
C111 VDD1.t3 B 0.140269f
C112 VDD1.t4 B 0.140269f
C113 VDD1.n88 B 1.21249f
C114 VDD1.n89 B 2.45041f
C115 VP.n0 B 0.03283f
C116 VP.t1 B 1.19075f
C117 VP.n1 B 0.023524f
C118 VP.n2 B 0.024902f
C119 VP.t2 B 1.19075f
C120 VP.n3 B 0.04641f
C121 VP.n4 B 0.024902f
C122 VP.t0 B 1.19075f
C123 VP.n5 B 0.460928f
C124 VP.n6 B 0.024902f
C125 VP.n7 B 0.04641f
C126 VP.n8 B 0.024902f
C127 VP.t4 B 1.19075f
C128 VP.n9 B 0.023524f
C129 VP.n10 B 0.03283f
C130 VP.t3 B 1.19075f
C131 VP.n11 B 0.03283f
C132 VP.t5 B 1.19075f
C133 VP.n12 B 0.023524f
C134 VP.n13 B 0.024902f
C135 VP.t6 B 1.19075f
C136 VP.n14 B 0.04641f
C137 VP.n15 B 0.024902f
C138 VP.t8 B 1.19075f
C139 VP.n16 B 0.460928f
C140 VP.n17 B 0.024902f
C141 VP.n18 B 0.04641f
C142 VP.t7 B 1.34499f
C143 VP.n19 B 0.497012f
C144 VP.t9 B 1.19075f
C145 VP.n20 B 0.497154f
C146 VP.n21 B 0.02808f
C147 VP.n22 B 0.213327f
C148 VP.n23 B 0.024902f
C149 VP.n24 B 0.024902f
C150 VP.n25 B 0.032882f
C151 VP.n26 B 0.039822f
C152 VP.n27 B 0.04641f
C153 VP.n28 B 0.024902f
C154 VP.n29 B 0.024902f
C155 VP.n30 B 0.024902f
C156 VP.n31 B 0.04641f
C157 VP.n32 B 0.039822f
C158 VP.n33 B 0.032882f
C159 VP.n34 B 0.024902f
C160 VP.n35 B 0.024902f
C161 VP.n36 B 0.024902f
C162 VP.n37 B 0.02808f
C163 VP.n38 B 0.437431f
C164 VP.n39 B 0.041828f
C165 VP.n40 B 0.045704f
C166 VP.n41 B 0.024902f
C167 VP.n42 B 0.024902f
C168 VP.n43 B 0.024902f
C169 VP.n44 B 0.049887f
C170 VP.n45 B 0.032663f
C171 VP.n46 B 0.509481f
C172 VP.n47 B 1.30511f
C173 VP.n48 B 1.32372f
C174 VP.n49 B 0.509481f
C175 VP.n50 B 0.032663f
C176 VP.n51 B 0.049887f
C177 VP.n52 B 0.024902f
C178 VP.n53 B 0.024902f
C179 VP.n54 B 0.024902f
C180 VP.n55 B 0.045704f
C181 VP.n56 B 0.041828f
C182 VP.n57 B 0.437431f
C183 VP.n58 B 0.02808f
C184 VP.n59 B 0.024902f
C185 VP.n60 B 0.024902f
C186 VP.n61 B 0.024902f
C187 VP.n62 B 0.032882f
C188 VP.n63 B 0.039822f
C189 VP.n64 B 0.04641f
C190 VP.n65 B 0.024902f
C191 VP.n66 B 0.024902f
C192 VP.n67 B 0.024902f
C193 VP.n68 B 0.04641f
C194 VP.n69 B 0.039822f
C195 VP.n70 B 0.032882f
C196 VP.n71 B 0.024902f
C197 VP.n72 B 0.024902f
C198 VP.n73 B 0.024902f
C199 VP.n74 B 0.02808f
C200 VP.n75 B 0.437431f
C201 VP.n76 B 0.041828f
C202 VP.n77 B 0.045704f
C203 VP.n78 B 0.024902f
C204 VP.n79 B 0.024902f
C205 VP.n80 B 0.024902f
C206 VP.n81 B 0.049887f
C207 VP.n82 B 0.032663f
C208 VP.n83 B 0.509481f
C209 VP.n84 B 0.038069f
C210 VTAIL.t9 B 0.163488f
C211 VTAIL.t16 B 0.163488f
C212 VTAIL.n0 B 1.34255f
C213 VTAIL.n1 B 0.527069f
C214 VTAIL.n2 B 0.033666f
C215 VTAIL.n3 B 0.026355f
C216 VTAIL.n4 B 0.014578f
C217 VTAIL.n5 B 0.033474f
C218 VTAIL.n6 B 0.014995f
C219 VTAIL.n7 B 0.026355f
C220 VTAIL.n8 B 0.014162f
C221 VTAIL.n9 B 0.033474f
C222 VTAIL.n10 B 0.014995f
C223 VTAIL.n11 B 0.026355f
C224 VTAIL.n12 B 0.014162f
C225 VTAIL.n13 B 0.025105f
C226 VTAIL.n14 B 0.023663f
C227 VTAIL.t7 B 0.055961f
C228 VTAIL.n15 B 0.148051f
C229 VTAIL.n16 B 0.843044f
C230 VTAIL.n17 B 0.014162f
C231 VTAIL.n18 B 0.014995f
C232 VTAIL.n19 B 0.033474f
C233 VTAIL.n20 B 0.033474f
C234 VTAIL.n21 B 0.014995f
C235 VTAIL.n22 B 0.014162f
C236 VTAIL.n23 B 0.026355f
C237 VTAIL.n24 B 0.026355f
C238 VTAIL.n25 B 0.014162f
C239 VTAIL.n26 B 0.014995f
C240 VTAIL.n27 B 0.033474f
C241 VTAIL.n28 B 0.033474f
C242 VTAIL.n29 B 0.014995f
C243 VTAIL.n30 B 0.014162f
C244 VTAIL.n31 B 0.026355f
C245 VTAIL.n32 B 0.026355f
C246 VTAIL.n33 B 0.014162f
C247 VTAIL.n34 B 0.014162f
C248 VTAIL.n35 B 0.014995f
C249 VTAIL.n36 B 0.033474f
C250 VTAIL.n37 B 0.033474f
C251 VTAIL.n38 B 0.066491f
C252 VTAIL.n39 B 0.014578f
C253 VTAIL.n40 B 0.014162f
C254 VTAIL.n41 B 0.062718f
C255 VTAIL.n42 B 0.036645f
C256 VTAIL.n43 B 0.348936f
C257 VTAIL.t6 B 0.163488f
C258 VTAIL.t5 B 0.163488f
C259 VTAIL.n44 B 1.34255f
C260 VTAIL.n45 B 0.624985f
C261 VTAIL.t19 B 0.163488f
C262 VTAIL.t18 B 0.163488f
C263 VTAIL.n46 B 1.34255f
C264 VTAIL.n47 B 1.74801f
C265 VTAIL.t10 B 0.163488f
C266 VTAIL.t8 B 0.163488f
C267 VTAIL.n48 B 1.34256f
C268 VTAIL.n49 B 1.748f
C269 VTAIL.t11 B 0.163488f
C270 VTAIL.t13 B 0.163488f
C271 VTAIL.n50 B 1.34256f
C272 VTAIL.n51 B 0.624976f
C273 VTAIL.n52 B 0.033666f
C274 VTAIL.n53 B 0.026355f
C275 VTAIL.n54 B 0.014578f
C276 VTAIL.n55 B 0.033474f
C277 VTAIL.n56 B 0.014162f
C278 VTAIL.n57 B 0.014995f
C279 VTAIL.n58 B 0.026355f
C280 VTAIL.n59 B 0.014162f
C281 VTAIL.n60 B 0.033474f
C282 VTAIL.n61 B 0.014995f
C283 VTAIL.n62 B 0.026355f
C284 VTAIL.n63 B 0.014162f
C285 VTAIL.n64 B 0.025105f
C286 VTAIL.n65 B 0.023663f
C287 VTAIL.t12 B 0.055961f
C288 VTAIL.n66 B 0.148051f
C289 VTAIL.n67 B 0.843044f
C290 VTAIL.n68 B 0.014162f
C291 VTAIL.n69 B 0.014995f
C292 VTAIL.n70 B 0.033474f
C293 VTAIL.n71 B 0.033474f
C294 VTAIL.n72 B 0.014995f
C295 VTAIL.n73 B 0.014162f
C296 VTAIL.n74 B 0.026355f
C297 VTAIL.n75 B 0.026355f
C298 VTAIL.n76 B 0.014162f
C299 VTAIL.n77 B 0.014995f
C300 VTAIL.n78 B 0.033474f
C301 VTAIL.n79 B 0.033474f
C302 VTAIL.n80 B 0.014995f
C303 VTAIL.n81 B 0.014162f
C304 VTAIL.n82 B 0.026355f
C305 VTAIL.n83 B 0.026355f
C306 VTAIL.n84 B 0.014162f
C307 VTAIL.n85 B 0.014995f
C308 VTAIL.n86 B 0.033474f
C309 VTAIL.n87 B 0.033474f
C310 VTAIL.n88 B 0.066491f
C311 VTAIL.n89 B 0.014578f
C312 VTAIL.n90 B 0.014162f
C313 VTAIL.n91 B 0.062718f
C314 VTAIL.n92 B 0.036645f
C315 VTAIL.n93 B 0.348936f
C316 VTAIL.t0 B 0.163488f
C317 VTAIL.t4 B 0.163488f
C318 VTAIL.n94 B 1.34256f
C319 VTAIL.n95 B 0.569704f
C320 VTAIL.t2 B 0.163488f
C321 VTAIL.t1 B 0.163488f
C322 VTAIL.n96 B 1.34256f
C323 VTAIL.n97 B 0.624976f
C324 VTAIL.n98 B 0.033666f
C325 VTAIL.n99 B 0.026355f
C326 VTAIL.n100 B 0.014578f
C327 VTAIL.n101 B 0.033474f
C328 VTAIL.n102 B 0.014162f
C329 VTAIL.n103 B 0.014995f
C330 VTAIL.n104 B 0.026355f
C331 VTAIL.n105 B 0.014162f
C332 VTAIL.n106 B 0.033474f
C333 VTAIL.n107 B 0.014995f
C334 VTAIL.n108 B 0.026355f
C335 VTAIL.n109 B 0.014162f
C336 VTAIL.n110 B 0.025105f
C337 VTAIL.n111 B 0.023663f
C338 VTAIL.t3 B 0.055961f
C339 VTAIL.n112 B 0.148051f
C340 VTAIL.n113 B 0.843044f
C341 VTAIL.n114 B 0.014162f
C342 VTAIL.n115 B 0.014995f
C343 VTAIL.n116 B 0.033474f
C344 VTAIL.n117 B 0.033474f
C345 VTAIL.n118 B 0.014995f
C346 VTAIL.n119 B 0.014162f
C347 VTAIL.n120 B 0.026355f
C348 VTAIL.n121 B 0.026355f
C349 VTAIL.n122 B 0.014162f
C350 VTAIL.n123 B 0.014995f
C351 VTAIL.n124 B 0.033474f
C352 VTAIL.n125 B 0.033474f
C353 VTAIL.n126 B 0.014995f
C354 VTAIL.n127 B 0.014162f
C355 VTAIL.n128 B 0.026355f
C356 VTAIL.n129 B 0.026355f
C357 VTAIL.n130 B 0.014162f
C358 VTAIL.n131 B 0.014995f
C359 VTAIL.n132 B 0.033474f
C360 VTAIL.n133 B 0.033474f
C361 VTAIL.n134 B 0.066491f
C362 VTAIL.n135 B 0.014578f
C363 VTAIL.n136 B 0.014162f
C364 VTAIL.n137 B 0.062718f
C365 VTAIL.n138 B 0.036645f
C366 VTAIL.n139 B 1.33689f
C367 VTAIL.n140 B 0.033666f
C368 VTAIL.n141 B 0.026355f
C369 VTAIL.n142 B 0.014578f
C370 VTAIL.n143 B 0.033474f
C371 VTAIL.n144 B 0.014995f
C372 VTAIL.n145 B 0.026355f
C373 VTAIL.n146 B 0.014162f
C374 VTAIL.n147 B 0.033474f
C375 VTAIL.n148 B 0.014995f
C376 VTAIL.n149 B 0.026355f
C377 VTAIL.n150 B 0.014162f
C378 VTAIL.n151 B 0.025105f
C379 VTAIL.n152 B 0.023663f
C380 VTAIL.t14 B 0.055961f
C381 VTAIL.n153 B 0.148051f
C382 VTAIL.n154 B 0.843044f
C383 VTAIL.n155 B 0.014162f
C384 VTAIL.n156 B 0.014995f
C385 VTAIL.n157 B 0.033474f
C386 VTAIL.n158 B 0.033474f
C387 VTAIL.n159 B 0.014995f
C388 VTAIL.n160 B 0.014162f
C389 VTAIL.n161 B 0.026355f
C390 VTAIL.n162 B 0.026355f
C391 VTAIL.n163 B 0.014162f
C392 VTAIL.n164 B 0.014995f
C393 VTAIL.n165 B 0.033474f
C394 VTAIL.n166 B 0.033474f
C395 VTAIL.n167 B 0.014995f
C396 VTAIL.n168 B 0.014162f
C397 VTAIL.n169 B 0.026355f
C398 VTAIL.n170 B 0.026355f
C399 VTAIL.n171 B 0.014162f
C400 VTAIL.n172 B 0.014162f
C401 VTAIL.n173 B 0.014995f
C402 VTAIL.n174 B 0.033474f
C403 VTAIL.n175 B 0.033474f
C404 VTAIL.n176 B 0.066491f
C405 VTAIL.n177 B 0.014578f
C406 VTAIL.n178 B 0.014162f
C407 VTAIL.n179 B 0.062718f
C408 VTAIL.n180 B 0.036645f
C409 VTAIL.n181 B 1.33689f
C410 VTAIL.t15 B 0.163488f
C411 VTAIL.t17 B 0.163488f
C412 VTAIL.n182 B 1.34255f
C413 VTAIL.n183 B 0.477287f
C414 VDD2.n0 B 0.028668f
C415 VDD2.n1 B 0.022442f
C416 VDD2.n2 B 0.012414f
C417 VDD2.n3 B 0.028504f
C418 VDD2.n4 B 0.012769f
C419 VDD2.n5 B 0.022442f
C420 VDD2.n6 B 0.01206f
C421 VDD2.n7 B 0.028504f
C422 VDD2.n8 B 0.012769f
C423 VDD2.n9 B 0.022442f
C424 VDD2.n10 B 0.01206f
C425 VDD2.n11 B 0.021378f
C426 VDD2.n12 B 0.02015f
C427 VDD2.t3 B 0.047653f
C428 VDD2.n13 B 0.126071f
C429 VDD2.n14 B 0.717885f
C430 VDD2.n15 B 0.01206f
C431 VDD2.n16 B 0.012769f
C432 VDD2.n17 B 0.028504f
C433 VDD2.n18 B 0.028504f
C434 VDD2.n19 B 0.012769f
C435 VDD2.n20 B 0.01206f
C436 VDD2.n21 B 0.022442f
C437 VDD2.n22 B 0.022442f
C438 VDD2.n23 B 0.01206f
C439 VDD2.n24 B 0.012769f
C440 VDD2.n25 B 0.028504f
C441 VDD2.n26 B 0.028504f
C442 VDD2.n27 B 0.012769f
C443 VDD2.n28 B 0.01206f
C444 VDD2.n29 B 0.022442f
C445 VDD2.n30 B 0.022442f
C446 VDD2.n31 B 0.01206f
C447 VDD2.n32 B 0.01206f
C448 VDD2.n33 B 0.012769f
C449 VDD2.n34 B 0.028504f
C450 VDD2.n35 B 0.028504f
C451 VDD2.n36 B 0.056619f
C452 VDD2.n37 B 0.012414f
C453 VDD2.n38 B 0.01206f
C454 VDD2.n39 B 0.053407f
C455 VDD2.n40 B 0.055562f
C456 VDD2.t5 B 0.139216f
C457 VDD2.t2 B 0.139216f
C458 VDD2.n41 B 1.20339f
C459 VDD2.n42 B 0.575308f
C460 VDD2.t0 B 0.139216f
C461 VDD2.t8 B 0.139216f
C462 VDD2.n43 B 1.2148f
C463 VDD2.n44 B 2.22007f
C464 VDD2.n45 B 0.028668f
C465 VDD2.n46 B 0.022442f
C466 VDD2.n47 B 0.012414f
C467 VDD2.n48 B 0.028504f
C468 VDD2.n49 B 0.01206f
C469 VDD2.n50 B 0.012769f
C470 VDD2.n51 B 0.022442f
C471 VDD2.n52 B 0.01206f
C472 VDD2.n53 B 0.028504f
C473 VDD2.n54 B 0.012769f
C474 VDD2.n55 B 0.022442f
C475 VDD2.n56 B 0.01206f
C476 VDD2.n57 B 0.021378f
C477 VDD2.n58 B 0.02015f
C478 VDD2.t9 B 0.047653f
C479 VDD2.n59 B 0.126071f
C480 VDD2.n60 B 0.717885f
C481 VDD2.n61 B 0.01206f
C482 VDD2.n62 B 0.012769f
C483 VDD2.n63 B 0.028504f
C484 VDD2.n64 B 0.028504f
C485 VDD2.n65 B 0.012769f
C486 VDD2.n66 B 0.01206f
C487 VDD2.n67 B 0.022442f
C488 VDD2.n68 B 0.022442f
C489 VDD2.n69 B 0.01206f
C490 VDD2.n70 B 0.012769f
C491 VDD2.n71 B 0.028504f
C492 VDD2.n72 B 0.028504f
C493 VDD2.n73 B 0.012769f
C494 VDD2.n74 B 0.01206f
C495 VDD2.n75 B 0.022442f
C496 VDD2.n76 B 0.022442f
C497 VDD2.n77 B 0.01206f
C498 VDD2.n78 B 0.012769f
C499 VDD2.n79 B 0.028504f
C500 VDD2.n80 B 0.028504f
C501 VDD2.n81 B 0.056619f
C502 VDD2.n82 B 0.012414f
C503 VDD2.n83 B 0.01206f
C504 VDD2.n84 B 0.053407f
C505 VDD2.n85 B 0.046688f
C506 VDD2.n86 B 2.19013f
C507 VDD2.t4 B 0.139216f
C508 VDD2.t1 B 0.139216f
C509 VDD2.n87 B 1.2034f
C510 VDD2.n88 B 0.385182f
C511 VDD2.t7 B 0.139216f
C512 VDD2.t6 B 0.139216f
C513 VDD2.n89 B 1.21477f
C514 VN.n0 B 0.032331f
C515 VN.t3 B 1.17265f
C516 VN.n1 B 0.023166f
C517 VN.n2 B 0.024523f
C518 VN.t0 B 1.17265f
C519 VN.n3 B 0.045705f
C520 VN.n4 B 0.024523f
C521 VN.t2 B 1.17265f
C522 VN.n5 B 0.453921f
C523 VN.n6 B 0.024523f
C524 VN.n7 B 0.045705f
C525 VN.t8 B 1.32454f
C526 VN.n8 B 0.489456f
C527 VN.t1 B 1.17265f
C528 VN.n9 B 0.489595f
C529 VN.n10 B 0.027653f
C530 VN.n11 B 0.210084f
C531 VN.n12 B 0.024523f
C532 VN.n13 B 0.024523f
C533 VN.n14 B 0.032382f
C534 VN.n15 B 0.039216f
C535 VN.n16 B 0.045705f
C536 VN.n17 B 0.024523f
C537 VN.n18 B 0.024523f
C538 VN.n19 B 0.024523f
C539 VN.n20 B 0.045705f
C540 VN.n21 B 0.039216f
C541 VN.n22 B 0.032382f
C542 VN.n23 B 0.024523f
C543 VN.n24 B 0.024523f
C544 VN.n25 B 0.024523f
C545 VN.n26 B 0.027653f
C546 VN.n27 B 0.43078f
C547 VN.n28 B 0.041192f
C548 VN.n29 B 0.045009f
C549 VN.n30 B 0.024523f
C550 VN.n31 B 0.024523f
C551 VN.n32 B 0.024523f
C552 VN.n33 B 0.049128f
C553 VN.n34 B 0.032166f
C554 VN.n35 B 0.501735f
C555 VN.n36 B 0.03749f
C556 VN.n37 B 0.032331f
C557 VN.t7 B 1.17265f
C558 VN.n38 B 0.023166f
C559 VN.n39 B 0.024523f
C560 VN.t9 B 1.17265f
C561 VN.n40 B 0.045705f
C562 VN.n41 B 0.024523f
C563 VN.t6 B 1.17265f
C564 VN.n42 B 0.453921f
C565 VN.n43 B 0.024523f
C566 VN.n44 B 0.045705f
C567 VN.t5 B 1.32454f
C568 VN.n45 B 0.489456f
C569 VN.t4 B 1.17265f
C570 VN.n46 B 0.489595f
C571 VN.n47 B 0.027653f
C572 VN.n48 B 0.210084f
C573 VN.n49 B 0.024523f
C574 VN.n50 B 0.024523f
C575 VN.n51 B 0.032382f
C576 VN.n52 B 0.039216f
C577 VN.n53 B 0.045705f
C578 VN.n54 B 0.024523f
C579 VN.n55 B 0.024523f
C580 VN.n56 B 0.024523f
C581 VN.n57 B 0.045705f
C582 VN.n58 B 0.039216f
C583 VN.n59 B 0.032382f
C584 VN.n60 B 0.024523f
C585 VN.n61 B 0.024523f
C586 VN.n62 B 0.024523f
C587 VN.n63 B 0.027653f
C588 VN.n64 B 0.43078f
C589 VN.n65 B 0.041192f
C590 VN.n66 B 0.045009f
C591 VN.n67 B 0.024523f
C592 VN.n68 B 0.024523f
C593 VN.n69 B 0.024523f
C594 VN.n70 B 0.049128f
C595 VN.n71 B 0.032166f
C596 VN.n72 B 0.501735f
C597 VN.n73 B 1.29853f
.ends

