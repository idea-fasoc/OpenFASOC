* NGSPICE file created from diff_pair_sample_1541.ext - technology: sky130A

.subckt diff_pair_sample_1541 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=5.2065 ps=27.48 w=13.35 l=3.31
X1 VTAIL.t5 VN.t0 VDD2.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=2.20275 ps=13.68 w=13.35 l=3.31
X2 VTAIL.t9 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=2.20275 ps=13.68 w=13.35 l=3.31
X3 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=2.20275 ps=13.68 w=13.35 l=3.31
X4 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=0 ps=0 w=13.35 l=3.31
X5 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=2.20275 ps=13.68 w=13.35 l=3.31
X6 VDD1.t3 VP.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=2.20275 ps=13.68 w=13.35 l=3.31
X7 VTAIL.t6 VP.t3 VDD1.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=2.20275 ps=13.68 w=13.35 l=3.31
X8 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=5.2065 ps=27.48 w=13.35 l=3.31
X9 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=5.2065 ps=27.48 w=13.35 l=3.31
X10 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=0 ps=0 w=13.35 l=3.31
X11 VDD1.t1 VP.t4 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=2.20275 ps=13.68 w=13.35 l=3.31
X12 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=0 ps=0 w=13.35 l=3.31
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=0 ps=0 w=13.35 l=3.31
X14 VDD1.t0 VP.t5 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.20275 pd=13.68 as=5.2065 ps=27.48 w=13.35 l=3.31
X15 VDD2.t0 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.2065 pd=27.48 as=2.20275 ps=13.68 w=13.35 l=3.31
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t4 130.5
R22 VP.n8 VP.t2 97.2014
R23 VP.n4 VP.t1 97.2014
R24 VP.n0 VP.t5 97.2014
R25 VP.n9 VP.t0 97.2014
R26 VP.n13 VP.t3 97.2014
R27 VP.n27 VP.n8 70.9831
R28 VP.n50 VP.n0 70.9831
R29 VP.n26 VP.n9 70.9831
R30 VP.n14 VP.n13 62.0573
R31 VP.n27 VP.n26 52.666
R32 VP.n31 VP.n6 47.2923
R33 VP.n46 VP.n2 47.2923
R34 VP.n22 VP.n11 47.2923
R35 VP.n35 VP.n6 33.6945
R36 VP.n42 VP.n2 33.6945
R37 VP.n18 VP.n11 33.6945
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 19.0848
R51 VP.n48 VP.n0 19.0848
R52 VP.n24 VP.n9 19.0848
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 3.94731
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n290 VTAIL.n224 214.453
R81 VTAIL.n68 VTAIL.n2 214.453
R82 VTAIL.n218 VTAIL.n152 214.453
R83 VTAIL.n144 VTAIL.n78 214.453
R84 VTAIL.n249 VTAIL.n248 185
R85 VTAIL.n251 VTAIL.n250 185
R86 VTAIL.n244 VTAIL.n243 185
R87 VTAIL.n257 VTAIL.n256 185
R88 VTAIL.n259 VTAIL.n258 185
R89 VTAIL.n240 VTAIL.n239 185
R90 VTAIL.n265 VTAIL.n264 185
R91 VTAIL.n267 VTAIL.n266 185
R92 VTAIL.n236 VTAIL.n235 185
R93 VTAIL.n273 VTAIL.n272 185
R94 VTAIL.n275 VTAIL.n274 185
R95 VTAIL.n232 VTAIL.n231 185
R96 VTAIL.n281 VTAIL.n280 185
R97 VTAIL.n283 VTAIL.n282 185
R98 VTAIL.n228 VTAIL.n227 185
R99 VTAIL.n289 VTAIL.n288 185
R100 VTAIL.n291 VTAIL.n290 185
R101 VTAIL.n27 VTAIL.n26 185
R102 VTAIL.n29 VTAIL.n28 185
R103 VTAIL.n22 VTAIL.n21 185
R104 VTAIL.n35 VTAIL.n34 185
R105 VTAIL.n37 VTAIL.n36 185
R106 VTAIL.n18 VTAIL.n17 185
R107 VTAIL.n43 VTAIL.n42 185
R108 VTAIL.n45 VTAIL.n44 185
R109 VTAIL.n14 VTAIL.n13 185
R110 VTAIL.n51 VTAIL.n50 185
R111 VTAIL.n53 VTAIL.n52 185
R112 VTAIL.n10 VTAIL.n9 185
R113 VTAIL.n59 VTAIL.n58 185
R114 VTAIL.n61 VTAIL.n60 185
R115 VTAIL.n6 VTAIL.n5 185
R116 VTAIL.n67 VTAIL.n66 185
R117 VTAIL.n69 VTAIL.n68 185
R118 VTAIL.n219 VTAIL.n218 185
R119 VTAIL.n217 VTAIL.n216 185
R120 VTAIL.n156 VTAIL.n155 185
R121 VTAIL.n211 VTAIL.n210 185
R122 VTAIL.n209 VTAIL.n208 185
R123 VTAIL.n160 VTAIL.n159 185
R124 VTAIL.n203 VTAIL.n202 185
R125 VTAIL.n201 VTAIL.n200 185
R126 VTAIL.n164 VTAIL.n163 185
R127 VTAIL.n195 VTAIL.n194 185
R128 VTAIL.n193 VTAIL.n192 185
R129 VTAIL.n168 VTAIL.n167 185
R130 VTAIL.n187 VTAIL.n186 185
R131 VTAIL.n185 VTAIL.n184 185
R132 VTAIL.n172 VTAIL.n171 185
R133 VTAIL.n179 VTAIL.n178 185
R134 VTAIL.n177 VTAIL.n176 185
R135 VTAIL.n145 VTAIL.n144 185
R136 VTAIL.n143 VTAIL.n142 185
R137 VTAIL.n82 VTAIL.n81 185
R138 VTAIL.n137 VTAIL.n136 185
R139 VTAIL.n135 VTAIL.n134 185
R140 VTAIL.n86 VTAIL.n85 185
R141 VTAIL.n129 VTAIL.n128 185
R142 VTAIL.n127 VTAIL.n126 185
R143 VTAIL.n90 VTAIL.n89 185
R144 VTAIL.n121 VTAIL.n120 185
R145 VTAIL.n119 VTAIL.n118 185
R146 VTAIL.n94 VTAIL.n93 185
R147 VTAIL.n113 VTAIL.n112 185
R148 VTAIL.n111 VTAIL.n110 185
R149 VTAIL.n98 VTAIL.n97 185
R150 VTAIL.n105 VTAIL.n104 185
R151 VTAIL.n103 VTAIL.n102 185
R152 VTAIL.n247 VTAIL.t2 147.659
R153 VTAIL.n25 VTAIL.t7 147.659
R154 VTAIL.n175 VTAIL.t8 147.659
R155 VTAIL.n101 VTAIL.t1 147.659
R156 VTAIL.n250 VTAIL.n249 104.615
R157 VTAIL.n250 VTAIL.n243 104.615
R158 VTAIL.n257 VTAIL.n243 104.615
R159 VTAIL.n258 VTAIL.n257 104.615
R160 VTAIL.n258 VTAIL.n239 104.615
R161 VTAIL.n265 VTAIL.n239 104.615
R162 VTAIL.n266 VTAIL.n265 104.615
R163 VTAIL.n266 VTAIL.n235 104.615
R164 VTAIL.n273 VTAIL.n235 104.615
R165 VTAIL.n274 VTAIL.n273 104.615
R166 VTAIL.n274 VTAIL.n231 104.615
R167 VTAIL.n281 VTAIL.n231 104.615
R168 VTAIL.n282 VTAIL.n281 104.615
R169 VTAIL.n282 VTAIL.n227 104.615
R170 VTAIL.n289 VTAIL.n227 104.615
R171 VTAIL.n290 VTAIL.n289 104.615
R172 VTAIL.n28 VTAIL.n27 104.615
R173 VTAIL.n28 VTAIL.n21 104.615
R174 VTAIL.n35 VTAIL.n21 104.615
R175 VTAIL.n36 VTAIL.n35 104.615
R176 VTAIL.n36 VTAIL.n17 104.615
R177 VTAIL.n43 VTAIL.n17 104.615
R178 VTAIL.n44 VTAIL.n43 104.615
R179 VTAIL.n44 VTAIL.n13 104.615
R180 VTAIL.n51 VTAIL.n13 104.615
R181 VTAIL.n52 VTAIL.n51 104.615
R182 VTAIL.n52 VTAIL.n9 104.615
R183 VTAIL.n59 VTAIL.n9 104.615
R184 VTAIL.n60 VTAIL.n59 104.615
R185 VTAIL.n60 VTAIL.n5 104.615
R186 VTAIL.n67 VTAIL.n5 104.615
R187 VTAIL.n68 VTAIL.n67 104.615
R188 VTAIL.n218 VTAIL.n217 104.615
R189 VTAIL.n217 VTAIL.n155 104.615
R190 VTAIL.n210 VTAIL.n155 104.615
R191 VTAIL.n210 VTAIL.n209 104.615
R192 VTAIL.n209 VTAIL.n159 104.615
R193 VTAIL.n202 VTAIL.n159 104.615
R194 VTAIL.n202 VTAIL.n201 104.615
R195 VTAIL.n201 VTAIL.n163 104.615
R196 VTAIL.n194 VTAIL.n163 104.615
R197 VTAIL.n194 VTAIL.n193 104.615
R198 VTAIL.n193 VTAIL.n167 104.615
R199 VTAIL.n186 VTAIL.n167 104.615
R200 VTAIL.n186 VTAIL.n185 104.615
R201 VTAIL.n185 VTAIL.n171 104.615
R202 VTAIL.n178 VTAIL.n171 104.615
R203 VTAIL.n178 VTAIL.n177 104.615
R204 VTAIL.n144 VTAIL.n143 104.615
R205 VTAIL.n143 VTAIL.n81 104.615
R206 VTAIL.n136 VTAIL.n81 104.615
R207 VTAIL.n136 VTAIL.n135 104.615
R208 VTAIL.n135 VTAIL.n85 104.615
R209 VTAIL.n128 VTAIL.n85 104.615
R210 VTAIL.n128 VTAIL.n127 104.615
R211 VTAIL.n127 VTAIL.n89 104.615
R212 VTAIL.n120 VTAIL.n89 104.615
R213 VTAIL.n120 VTAIL.n119 104.615
R214 VTAIL.n119 VTAIL.n93 104.615
R215 VTAIL.n112 VTAIL.n93 104.615
R216 VTAIL.n112 VTAIL.n111 104.615
R217 VTAIL.n111 VTAIL.n97 104.615
R218 VTAIL.n104 VTAIL.n97 104.615
R219 VTAIL.n104 VTAIL.n103 104.615
R220 VTAIL.n249 VTAIL.t2 52.3082
R221 VTAIL.n27 VTAIL.t7 52.3082
R222 VTAIL.n177 VTAIL.t8 52.3082
R223 VTAIL.n103 VTAIL.t1 52.3082
R224 VTAIL.n151 VTAIL.n150 47.3499
R225 VTAIL.n77 VTAIL.n76 47.3499
R226 VTAIL.n1 VTAIL.n0 47.3498
R227 VTAIL.n75 VTAIL.n74 47.3498
R228 VTAIL.n295 VTAIL.n294 35.0944
R229 VTAIL.n73 VTAIL.n72 35.0944
R230 VTAIL.n223 VTAIL.n222 35.0944
R231 VTAIL.n149 VTAIL.n148 35.0944
R232 VTAIL.n77 VTAIL.n75 30.1514
R233 VTAIL.n295 VTAIL.n223 27.0134
R234 VTAIL.n248 VTAIL.n247 15.6677
R235 VTAIL.n26 VTAIL.n25 15.6677
R236 VTAIL.n176 VTAIL.n175 15.6677
R237 VTAIL.n102 VTAIL.n101 15.6677
R238 VTAIL.n251 VTAIL.n246 12.8005
R239 VTAIL.n292 VTAIL.n291 12.8005
R240 VTAIL.n29 VTAIL.n24 12.8005
R241 VTAIL.n70 VTAIL.n69 12.8005
R242 VTAIL.n220 VTAIL.n219 12.8005
R243 VTAIL.n179 VTAIL.n174 12.8005
R244 VTAIL.n146 VTAIL.n145 12.8005
R245 VTAIL.n105 VTAIL.n100 12.8005
R246 VTAIL.n252 VTAIL.n244 12.0247
R247 VTAIL.n288 VTAIL.n226 12.0247
R248 VTAIL.n30 VTAIL.n22 12.0247
R249 VTAIL.n66 VTAIL.n4 12.0247
R250 VTAIL.n216 VTAIL.n154 12.0247
R251 VTAIL.n180 VTAIL.n172 12.0247
R252 VTAIL.n142 VTAIL.n80 12.0247
R253 VTAIL.n106 VTAIL.n98 12.0247
R254 VTAIL.n256 VTAIL.n255 11.249
R255 VTAIL.n287 VTAIL.n228 11.249
R256 VTAIL.n34 VTAIL.n33 11.249
R257 VTAIL.n65 VTAIL.n6 11.249
R258 VTAIL.n215 VTAIL.n156 11.249
R259 VTAIL.n184 VTAIL.n183 11.249
R260 VTAIL.n141 VTAIL.n82 11.249
R261 VTAIL.n110 VTAIL.n109 11.249
R262 VTAIL.n259 VTAIL.n242 10.4732
R263 VTAIL.n284 VTAIL.n283 10.4732
R264 VTAIL.n37 VTAIL.n20 10.4732
R265 VTAIL.n62 VTAIL.n61 10.4732
R266 VTAIL.n212 VTAIL.n211 10.4732
R267 VTAIL.n187 VTAIL.n170 10.4732
R268 VTAIL.n138 VTAIL.n137 10.4732
R269 VTAIL.n113 VTAIL.n96 10.4732
R270 VTAIL.n260 VTAIL.n240 9.69747
R271 VTAIL.n280 VTAIL.n230 9.69747
R272 VTAIL.n38 VTAIL.n18 9.69747
R273 VTAIL.n58 VTAIL.n8 9.69747
R274 VTAIL.n208 VTAIL.n158 9.69747
R275 VTAIL.n188 VTAIL.n168 9.69747
R276 VTAIL.n134 VTAIL.n84 9.69747
R277 VTAIL.n114 VTAIL.n94 9.69747
R278 VTAIL.n294 VTAIL.n293 9.45567
R279 VTAIL.n72 VTAIL.n71 9.45567
R280 VTAIL.n222 VTAIL.n221 9.45567
R281 VTAIL.n148 VTAIL.n147 9.45567
R282 VTAIL.n269 VTAIL.n268 9.3005
R283 VTAIL.n238 VTAIL.n237 9.3005
R284 VTAIL.n263 VTAIL.n262 9.3005
R285 VTAIL.n261 VTAIL.n260 9.3005
R286 VTAIL.n242 VTAIL.n241 9.3005
R287 VTAIL.n255 VTAIL.n254 9.3005
R288 VTAIL.n253 VTAIL.n252 9.3005
R289 VTAIL.n246 VTAIL.n245 9.3005
R290 VTAIL.n271 VTAIL.n270 9.3005
R291 VTAIL.n234 VTAIL.n233 9.3005
R292 VTAIL.n277 VTAIL.n276 9.3005
R293 VTAIL.n279 VTAIL.n278 9.3005
R294 VTAIL.n230 VTAIL.n229 9.3005
R295 VTAIL.n285 VTAIL.n284 9.3005
R296 VTAIL.n287 VTAIL.n286 9.3005
R297 VTAIL.n226 VTAIL.n225 9.3005
R298 VTAIL.n293 VTAIL.n292 9.3005
R299 VTAIL.n47 VTAIL.n46 9.3005
R300 VTAIL.n16 VTAIL.n15 9.3005
R301 VTAIL.n41 VTAIL.n40 9.3005
R302 VTAIL.n39 VTAIL.n38 9.3005
R303 VTAIL.n20 VTAIL.n19 9.3005
R304 VTAIL.n33 VTAIL.n32 9.3005
R305 VTAIL.n31 VTAIL.n30 9.3005
R306 VTAIL.n24 VTAIL.n23 9.3005
R307 VTAIL.n49 VTAIL.n48 9.3005
R308 VTAIL.n12 VTAIL.n11 9.3005
R309 VTAIL.n55 VTAIL.n54 9.3005
R310 VTAIL.n57 VTAIL.n56 9.3005
R311 VTAIL.n8 VTAIL.n7 9.3005
R312 VTAIL.n63 VTAIL.n62 9.3005
R313 VTAIL.n65 VTAIL.n64 9.3005
R314 VTAIL.n4 VTAIL.n3 9.3005
R315 VTAIL.n71 VTAIL.n70 9.3005
R316 VTAIL.n162 VTAIL.n161 9.3005
R317 VTAIL.n205 VTAIL.n204 9.3005
R318 VTAIL.n207 VTAIL.n206 9.3005
R319 VTAIL.n158 VTAIL.n157 9.3005
R320 VTAIL.n213 VTAIL.n212 9.3005
R321 VTAIL.n215 VTAIL.n214 9.3005
R322 VTAIL.n154 VTAIL.n153 9.3005
R323 VTAIL.n221 VTAIL.n220 9.3005
R324 VTAIL.n199 VTAIL.n198 9.3005
R325 VTAIL.n197 VTAIL.n196 9.3005
R326 VTAIL.n166 VTAIL.n165 9.3005
R327 VTAIL.n191 VTAIL.n190 9.3005
R328 VTAIL.n189 VTAIL.n188 9.3005
R329 VTAIL.n170 VTAIL.n169 9.3005
R330 VTAIL.n183 VTAIL.n182 9.3005
R331 VTAIL.n181 VTAIL.n180 9.3005
R332 VTAIL.n174 VTAIL.n173 9.3005
R333 VTAIL.n88 VTAIL.n87 9.3005
R334 VTAIL.n131 VTAIL.n130 9.3005
R335 VTAIL.n133 VTAIL.n132 9.3005
R336 VTAIL.n84 VTAIL.n83 9.3005
R337 VTAIL.n139 VTAIL.n138 9.3005
R338 VTAIL.n141 VTAIL.n140 9.3005
R339 VTAIL.n80 VTAIL.n79 9.3005
R340 VTAIL.n147 VTAIL.n146 9.3005
R341 VTAIL.n125 VTAIL.n124 9.3005
R342 VTAIL.n123 VTAIL.n122 9.3005
R343 VTAIL.n92 VTAIL.n91 9.3005
R344 VTAIL.n117 VTAIL.n116 9.3005
R345 VTAIL.n115 VTAIL.n114 9.3005
R346 VTAIL.n96 VTAIL.n95 9.3005
R347 VTAIL.n109 VTAIL.n108 9.3005
R348 VTAIL.n107 VTAIL.n106 9.3005
R349 VTAIL.n100 VTAIL.n99 9.3005
R350 VTAIL.n264 VTAIL.n263 8.92171
R351 VTAIL.n279 VTAIL.n232 8.92171
R352 VTAIL.n42 VTAIL.n41 8.92171
R353 VTAIL.n57 VTAIL.n10 8.92171
R354 VTAIL.n207 VTAIL.n160 8.92171
R355 VTAIL.n192 VTAIL.n191 8.92171
R356 VTAIL.n133 VTAIL.n86 8.92171
R357 VTAIL.n118 VTAIL.n117 8.92171
R358 VTAIL.n294 VTAIL.n224 8.2187
R359 VTAIL.n72 VTAIL.n2 8.2187
R360 VTAIL.n222 VTAIL.n152 8.2187
R361 VTAIL.n148 VTAIL.n78 8.2187
R362 VTAIL.n267 VTAIL.n238 8.14595
R363 VTAIL.n276 VTAIL.n275 8.14595
R364 VTAIL.n45 VTAIL.n16 8.14595
R365 VTAIL.n54 VTAIL.n53 8.14595
R366 VTAIL.n204 VTAIL.n203 8.14595
R367 VTAIL.n195 VTAIL.n166 8.14595
R368 VTAIL.n130 VTAIL.n129 8.14595
R369 VTAIL.n121 VTAIL.n92 8.14595
R370 VTAIL.n268 VTAIL.n236 7.3702
R371 VTAIL.n272 VTAIL.n234 7.3702
R372 VTAIL.n46 VTAIL.n14 7.3702
R373 VTAIL.n50 VTAIL.n12 7.3702
R374 VTAIL.n200 VTAIL.n162 7.3702
R375 VTAIL.n196 VTAIL.n164 7.3702
R376 VTAIL.n126 VTAIL.n88 7.3702
R377 VTAIL.n122 VTAIL.n90 7.3702
R378 VTAIL.n271 VTAIL.n236 6.59444
R379 VTAIL.n272 VTAIL.n271 6.59444
R380 VTAIL.n49 VTAIL.n14 6.59444
R381 VTAIL.n50 VTAIL.n49 6.59444
R382 VTAIL.n200 VTAIL.n199 6.59444
R383 VTAIL.n199 VTAIL.n164 6.59444
R384 VTAIL.n126 VTAIL.n125 6.59444
R385 VTAIL.n125 VTAIL.n90 6.59444
R386 VTAIL.n268 VTAIL.n267 5.81868
R387 VTAIL.n275 VTAIL.n234 5.81868
R388 VTAIL.n46 VTAIL.n45 5.81868
R389 VTAIL.n53 VTAIL.n12 5.81868
R390 VTAIL.n203 VTAIL.n162 5.81868
R391 VTAIL.n196 VTAIL.n195 5.81868
R392 VTAIL.n129 VTAIL.n88 5.81868
R393 VTAIL.n122 VTAIL.n121 5.81868
R394 VTAIL.n292 VTAIL.n224 5.3904
R395 VTAIL.n70 VTAIL.n2 5.3904
R396 VTAIL.n220 VTAIL.n152 5.3904
R397 VTAIL.n146 VTAIL.n78 5.3904
R398 VTAIL.n264 VTAIL.n238 5.04292
R399 VTAIL.n276 VTAIL.n232 5.04292
R400 VTAIL.n42 VTAIL.n16 5.04292
R401 VTAIL.n54 VTAIL.n10 5.04292
R402 VTAIL.n204 VTAIL.n160 5.04292
R403 VTAIL.n192 VTAIL.n166 5.04292
R404 VTAIL.n130 VTAIL.n86 5.04292
R405 VTAIL.n118 VTAIL.n92 5.04292
R406 VTAIL.n247 VTAIL.n245 4.38563
R407 VTAIL.n25 VTAIL.n23 4.38563
R408 VTAIL.n175 VTAIL.n173 4.38563
R409 VTAIL.n101 VTAIL.n99 4.38563
R410 VTAIL.n263 VTAIL.n240 4.26717
R411 VTAIL.n280 VTAIL.n279 4.26717
R412 VTAIL.n41 VTAIL.n18 4.26717
R413 VTAIL.n58 VTAIL.n57 4.26717
R414 VTAIL.n208 VTAIL.n207 4.26717
R415 VTAIL.n191 VTAIL.n168 4.26717
R416 VTAIL.n134 VTAIL.n133 4.26717
R417 VTAIL.n117 VTAIL.n94 4.26717
R418 VTAIL.n260 VTAIL.n259 3.49141
R419 VTAIL.n283 VTAIL.n230 3.49141
R420 VTAIL.n38 VTAIL.n37 3.49141
R421 VTAIL.n61 VTAIL.n8 3.49141
R422 VTAIL.n211 VTAIL.n158 3.49141
R423 VTAIL.n188 VTAIL.n187 3.49141
R424 VTAIL.n137 VTAIL.n84 3.49141
R425 VTAIL.n114 VTAIL.n113 3.49141
R426 VTAIL.n149 VTAIL.n77 3.13843
R427 VTAIL.n223 VTAIL.n151 3.13843
R428 VTAIL.n75 VTAIL.n73 3.13843
R429 VTAIL.n256 VTAIL.n242 2.71565
R430 VTAIL.n284 VTAIL.n228 2.71565
R431 VTAIL.n34 VTAIL.n20 2.71565
R432 VTAIL.n62 VTAIL.n6 2.71565
R433 VTAIL.n212 VTAIL.n156 2.71565
R434 VTAIL.n184 VTAIL.n170 2.71565
R435 VTAIL.n138 VTAIL.n82 2.71565
R436 VTAIL.n110 VTAIL.n96 2.71565
R437 VTAIL VTAIL.n295 2.29576
R438 VTAIL.n151 VTAIL.n149 2.03929
R439 VTAIL.n73 VTAIL.n1 2.03929
R440 VTAIL.n255 VTAIL.n244 1.93989
R441 VTAIL.n288 VTAIL.n287 1.93989
R442 VTAIL.n33 VTAIL.n22 1.93989
R443 VTAIL.n66 VTAIL.n65 1.93989
R444 VTAIL.n216 VTAIL.n215 1.93989
R445 VTAIL.n183 VTAIL.n172 1.93989
R446 VTAIL.n142 VTAIL.n141 1.93989
R447 VTAIL.n109 VTAIL.n98 1.93989
R448 VTAIL.n0 VTAIL.t4 1.48365
R449 VTAIL.n0 VTAIL.t5 1.48365
R450 VTAIL.n74 VTAIL.t11 1.48365
R451 VTAIL.n74 VTAIL.t9 1.48365
R452 VTAIL.n150 VTAIL.t10 1.48365
R453 VTAIL.n150 VTAIL.t6 1.48365
R454 VTAIL.n76 VTAIL.t3 1.48365
R455 VTAIL.n76 VTAIL.t0 1.48365
R456 VTAIL.n252 VTAIL.n251 1.16414
R457 VTAIL.n291 VTAIL.n226 1.16414
R458 VTAIL.n30 VTAIL.n29 1.16414
R459 VTAIL.n69 VTAIL.n4 1.16414
R460 VTAIL.n219 VTAIL.n154 1.16414
R461 VTAIL.n180 VTAIL.n179 1.16414
R462 VTAIL.n145 VTAIL.n80 1.16414
R463 VTAIL.n106 VTAIL.n105 1.16414
R464 VTAIL VTAIL.n1 0.843172
R465 VTAIL.n248 VTAIL.n246 0.388379
R466 VTAIL.n26 VTAIL.n24 0.388379
R467 VTAIL.n176 VTAIL.n174 0.388379
R468 VTAIL.n102 VTAIL.n100 0.388379
R469 VTAIL.n253 VTAIL.n245 0.155672
R470 VTAIL.n254 VTAIL.n253 0.155672
R471 VTAIL.n254 VTAIL.n241 0.155672
R472 VTAIL.n261 VTAIL.n241 0.155672
R473 VTAIL.n262 VTAIL.n261 0.155672
R474 VTAIL.n262 VTAIL.n237 0.155672
R475 VTAIL.n269 VTAIL.n237 0.155672
R476 VTAIL.n270 VTAIL.n269 0.155672
R477 VTAIL.n270 VTAIL.n233 0.155672
R478 VTAIL.n277 VTAIL.n233 0.155672
R479 VTAIL.n278 VTAIL.n277 0.155672
R480 VTAIL.n278 VTAIL.n229 0.155672
R481 VTAIL.n285 VTAIL.n229 0.155672
R482 VTAIL.n286 VTAIL.n285 0.155672
R483 VTAIL.n286 VTAIL.n225 0.155672
R484 VTAIL.n293 VTAIL.n225 0.155672
R485 VTAIL.n31 VTAIL.n23 0.155672
R486 VTAIL.n32 VTAIL.n31 0.155672
R487 VTAIL.n32 VTAIL.n19 0.155672
R488 VTAIL.n39 VTAIL.n19 0.155672
R489 VTAIL.n40 VTAIL.n39 0.155672
R490 VTAIL.n40 VTAIL.n15 0.155672
R491 VTAIL.n47 VTAIL.n15 0.155672
R492 VTAIL.n48 VTAIL.n47 0.155672
R493 VTAIL.n48 VTAIL.n11 0.155672
R494 VTAIL.n55 VTAIL.n11 0.155672
R495 VTAIL.n56 VTAIL.n55 0.155672
R496 VTAIL.n56 VTAIL.n7 0.155672
R497 VTAIL.n63 VTAIL.n7 0.155672
R498 VTAIL.n64 VTAIL.n63 0.155672
R499 VTAIL.n64 VTAIL.n3 0.155672
R500 VTAIL.n71 VTAIL.n3 0.155672
R501 VTAIL.n221 VTAIL.n153 0.155672
R502 VTAIL.n214 VTAIL.n153 0.155672
R503 VTAIL.n214 VTAIL.n213 0.155672
R504 VTAIL.n213 VTAIL.n157 0.155672
R505 VTAIL.n206 VTAIL.n157 0.155672
R506 VTAIL.n206 VTAIL.n205 0.155672
R507 VTAIL.n205 VTAIL.n161 0.155672
R508 VTAIL.n198 VTAIL.n161 0.155672
R509 VTAIL.n198 VTAIL.n197 0.155672
R510 VTAIL.n197 VTAIL.n165 0.155672
R511 VTAIL.n190 VTAIL.n165 0.155672
R512 VTAIL.n190 VTAIL.n189 0.155672
R513 VTAIL.n189 VTAIL.n169 0.155672
R514 VTAIL.n182 VTAIL.n169 0.155672
R515 VTAIL.n182 VTAIL.n181 0.155672
R516 VTAIL.n181 VTAIL.n173 0.155672
R517 VTAIL.n147 VTAIL.n79 0.155672
R518 VTAIL.n140 VTAIL.n79 0.155672
R519 VTAIL.n140 VTAIL.n139 0.155672
R520 VTAIL.n139 VTAIL.n83 0.155672
R521 VTAIL.n132 VTAIL.n83 0.155672
R522 VTAIL.n132 VTAIL.n131 0.155672
R523 VTAIL.n131 VTAIL.n87 0.155672
R524 VTAIL.n124 VTAIL.n87 0.155672
R525 VTAIL.n124 VTAIL.n123 0.155672
R526 VTAIL.n123 VTAIL.n91 0.155672
R527 VTAIL.n116 VTAIL.n91 0.155672
R528 VTAIL.n116 VTAIL.n115 0.155672
R529 VTAIL.n115 VTAIL.n95 0.155672
R530 VTAIL.n108 VTAIL.n95 0.155672
R531 VTAIL.n108 VTAIL.n107 0.155672
R532 VTAIL.n107 VTAIL.n99 0.155672
R533 VDD1.n66 VDD1.n0 214.453
R534 VDD1.n137 VDD1.n71 214.453
R535 VDD1.n67 VDD1.n66 185
R536 VDD1.n65 VDD1.n64 185
R537 VDD1.n4 VDD1.n3 185
R538 VDD1.n59 VDD1.n58 185
R539 VDD1.n57 VDD1.n56 185
R540 VDD1.n8 VDD1.n7 185
R541 VDD1.n51 VDD1.n50 185
R542 VDD1.n49 VDD1.n48 185
R543 VDD1.n12 VDD1.n11 185
R544 VDD1.n43 VDD1.n42 185
R545 VDD1.n41 VDD1.n40 185
R546 VDD1.n16 VDD1.n15 185
R547 VDD1.n35 VDD1.n34 185
R548 VDD1.n33 VDD1.n32 185
R549 VDD1.n20 VDD1.n19 185
R550 VDD1.n27 VDD1.n26 185
R551 VDD1.n25 VDD1.n24 185
R552 VDD1.n96 VDD1.n95 185
R553 VDD1.n98 VDD1.n97 185
R554 VDD1.n91 VDD1.n90 185
R555 VDD1.n104 VDD1.n103 185
R556 VDD1.n106 VDD1.n105 185
R557 VDD1.n87 VDD1.n86 185
R558 VDD1.n112 VDD1.n111 185
R559 VDD1.n114 VDD1.n113 185
R560 VDD1.n83 VDD1.n82 185
R561 VDD1.n120 VDD1.n119 185
R562 VDD1.n122 VDD1.n121 185
R563 VDD1.n79 VDD1.n78 185
R564 VDD1.n128 VDD1.n127 185
R565 VDD1.n130 VDD1.n129 185
R566 VDD1.n75 VDD1.n74 185
R567 VDD1.n136 VDD1.n135 185
R568 VDD1.n138 VDD1.n137 185
R569 VDD1.n94 VDD1.t3 147.659
R570 VDD1.n23 VDD1.t1 147.659
R571 VDD1.n66 VDD1.n65 104.615
R572 VDD1.n65 VDD1.n3 104.615
R573 VDD1.n58 VDD1.n3 104.615
R574 VDD1.n58 VDD1.n57 104.615
R575 VDD1.n57 VDD1.n7 104.615
R576 VDD1.n50 VDD1.n7 104.615
R577 VDD1.n50 VDD1.n49 104.615
R578 VDD1.n49 VDD1.n11 104.615
R579 VDD1.n42 VDD1.n11 104.615
R580 VDD1.n42 VDD1.n41 104.615
R581 VDD1.n41 VDD1.n15 104.615
R582 VDD1.n34 VDD1.n15 104.615
R583 VDD1.n34 VDD1.n33 104.615
R584 VDD1.n33 VDD1.n19 104.615
R585 VDD1.n26 VDD1.n19 104.615
R586 VDD1.n26 VDD1.n25 104.615
R587 VDD1.n97 VDD1.n96 104.615
R588 VDD1.n97 VDD1.n90 104.615
R589 VDD1.n104 VDD1.n90 104.615
R590 VDD1.n105 VDD1.n104 104.615
R591 VDD1.n105 VDD1.n86 104.615
R592 VDD1.n112 VDD1.n86 104.615
R593 VDD1.n113 VDD1.n112 104.615
R594 VDD1.n113 VDD1.n82 104.615
R595 VDD1.n120 VDD1.n82 104.615
R596 VDD1.n121 VDD1.n120 104.615
R597 VDD1.n121 VDD1.n78 104.615
R598 VDD1.n128 VDD1.n78 104.615
R599 VDD1.n129 VDD1.n128 104.615
R600 VDD1.n129 VDD1.n74 104.615
R601 VDD1.n136 VDD1.n74 104.615
R602 VDD1.n137 VDD1.n136 104.615
R603 VDD1.n143 VDD1.n142 64.7577
R604 VDD1.n145 VDD1.n144 64.0286
R605 VDD1 VDD1.n70 54.1849
R606 VDD1.n143 VDD1.n141 54.0713
R607 VDD1.n25 VDD1.t1 52.3082
R608 VDD1.n96 VDD1.t3 52.3082
R609 VDD1.n145 VDD1.n143 47.5742
R610 VDD1.n24 VDD1.n23 15.6677
R611 VDD1.n95 VDD1.n94 15.6677
R612 VDD1.n68 VDD1.n67 12.8005
R613 VDD1.n27 VDD1.n22 12.8005
R614 VDD1.n98 VDD1.n93 12.8005
R615 VDD1.n139 VDD1.n138 12.8005
R616 VDD1.n64 VDD1.n2 12.0247
R617 VDD1.n28 VDD1.n20 12.0247
R618 VDD1.n99 VDD1.n91 12.0247
R619 VDD1.n135 VDD1.n73 12.0247
R620 VDD1.n63 VDD1.n4 11.249
R621 VDD1.n32 VDD1.n31 11.249
R622 VDD1.n103 VDD1.n102 11.249
R623 VDD1.n134 VDD1.n75 11.249
R624 VDD1.n60 VDD1.n59 10.4732
R625 VDD1.n35 VDD1.n18 10.4732
R626 VDD1.n106 VDD1.n89 10.4732
R627 VDD1.n131 VDD1.n130 10.4732
R628 VDD1.n56 VDD1.n6 9.69747
R629 VDD1.n36 VDD1.n16 9.69747
R630 VDD1.n107 VDD1.n87 9.69747
R631 VDD1.n127 VDD1.n77 9.69747
R632 VDD1.n70 VDD1.n69 9.45567
R633 VDD1.n141 VDD1.n140 9.45567
R634 VDD1.n10 VDD1.n9 9.3005
R635 VDD1.n53 VDD1.n52 9.3005
R636 VDD1.n55 VDD1.n54 9.3005
R637 VDD1.n6 VDD1.n5 9.3005
R638 VDD1.n61 VDD1.n60 9.3005
R639 VDD1.n63 VDD1.n62 9.3005
R640 VDD1.n2 VDD1.n1 9.3005
R641 VDD1.n69 VDD1.n68 9.3005
R642 VDD1.n47 VDD1.n46 9.3005
R643 VDD1.n45 VDD1.n44 9.3005
R644 VDD1.n14 VDD1.n13 9.3005
R645 VDD1.n39 VDD1.n38 9.3005
R646 VDD1.n37 VDD1.n36 9.3005
R647 VDD1.n18 VDD1.n17 9.3005
R648 VDD1.n31 VDD1.n30 9.3005
R649 VDD1.n29 VDD1.n28 9.3005
R650 VDD1.n22 VDD1.n21 9.3005
R651 VDD1.n116 VDD1.n115 9.3005
R652 VDD1.n85 VDD1.n84 9.3005
R653 VDD1.n110 VDD1.n109 9.3005
R654 VDD1.n108 VDD1.n107 9.3005
R655 VDD1.n89 VDD1.n88 9.3005
R656 VDD1.n102 VDD1.n101 9.3005
R657 VDD1.n100 VDD1.n99 9.3005
R658 VDD1.n93 VDD1.n92 9.3005
R659 VDD1.n118 VDD1.n117 9.3005
R660 VDD1.n81 VDD1.n80 9.3005
R661 VDD1.n124 VDD1.n123 9.3005
R662 VDD1.n126 VDD1.n125 9.3005
R663 VDD1.n77 VDD1.n76 9.3005
R664 VDD1.n132 VDD1.n131 9.3005
R665 VDD1.n134 VDD1.n133 9.3005
R666 VDD1.n73 VDD1.n72 9.3005
R667 VDD1.n140 VDD1.n139 9.3005
R668 VDD1.n55 VDD1.n8 8.92171
R669 VDD1.n40 VDD1.n39 8.92171
R670 VDD1.n111 VDD1.n110 8.92171
R671 VDD1.n126 VDD1.n79 8.92171
R672 VDD1.n70 VDD1.n0 8.2187
R673 VDD1.n141 VDD1.n71 8.2187
R674 VDD1.n52 VDD1.n51 8.14595
R675 VDD1.n43 VDD1.n14 8.14595
R676 VDD1.n114 VDD1.n85 8.14595
R677 VDD1.n123 VDD1.n122 8.14595
R678 VDD1.n48 VDD1.n10 7.3702
R679 VDD1.n44 VDD1.n12 7.3702
R680 VDD1.n115 VDD1.n83 7.3702
R681 VDD1.n119 VDD1.n81 7.3702
R682 VDD1.n48 VDD1.n47 6.59444
R683 VDD1.n47 VDD1.n12 6.59444
R684 VDD1.n118 VDD1.n83 6.59444
R685 VDD1.n119 VDD1.n118 6.59444
R686 VDD1.n51 VDD1.n10 5.81868
R687 VDD1.n44 VDD1.n43 5.81868
R688 VDD1.n115 VDD1.n114 5.81868
R689 VDD1.n122 VDD1.n81 5.81868
R690 VDD1.n68 VDD1.n0 5.3904
R691 VDD1.n139 VDD1.n71 5.3904
R692 VDD1.n52 VDD1.n8 5.04292
R693 VDD1.n40 VDD1.n14 5.04292
R694 VDD1.n111 VDD1.n85 5.04292
R695 VDD1.n123 VDD1.n79 5.04292
R696 VDD1.n94 VDD1.n92 4.38563
R697 VDD1.n23 VDD1.n21 4.38563
R698 VDD1.n56 VDD1.n55 4.26717
R699 VDD1.n39 VDD1.n16 4.26717
R700 VDD1.n110 VDD1.n87 4.26717
R701 VDD1.n127 VDD1.n126 4.26717
R702 VDD1.n59 VDD1.n6 3.49141
R703 VDD1.n36 VDD1.n35 3.49141
R704 VDD1.n107 VDD1.n106 3.49141
R705 VDD1.n130 VDD1.n77 3.49141
R706 VDD1.n60 VDD1.n4 2.71565
R707 VDD1.n32 VDD1.n18 2.71565
R708 VDD1.n103 VDD1.n89 2.71565
R709 VDD1.n131 VDD1.n75 2.71565
R710 VDD1.n64 VDD1.n63 1.93989
R711 VDD1.n31 VDD1.n20 1.93989
R712 VDD1.n102 VDD1.n91 1.93989
R713 VDD1.n135 VDD1.n134 1.93989
R714 VDD1.n144 VDD1.t2 1.48365
R715 VDD1.n144 VDD1.t5 1.48365
R716 VDD1.n142 VDD1.t4 1.48365
R717 VDD1.n142 VDD1.t0 1.48365
R718 VDD1.n67 VDD1.n2 1.16414
R719 VDD1.n28 VDD1.n27 1.16414
R720 VDD1.n99 VDD1.n98 1.16414
R721 VDD1.n138 VDD1.n73 1.16414
R722 VDD1 VDD1.n145 0.726793
R723 VDD1.n24 VDD1.n22 0.388379
R724 VDD1.n95 VDD1.n93 0.388379
R725 VDD1.n69 VDD1.n1 0.155672
R726 VDD1.n62 VDD1.n1 0.155672
R727 VDD1.n62 VDD1.n61 0.155672
R728 VDD1.n61 VDD1.n5 0.155672
R729 VDD1.n54 VDD1.n5 0.155672
R730 VDD1.n54 VDD1.n53 0.155672
R731 VDD1.n53 VDD1.n9 0.155672
R732 VDD1.n46 VDD1.n9 0.155672
R733 VDD1.n46 VDD1.n45 0.155672
R734 VDD1.n45 VDD1.n13 0.155672
R735 VDD1.n38 VDD1.n13 0.155672
R736 VDD1.n38 VDD1.n37 0.155672
R737 VDD1.n37 VDD1.n17 0.155672
R738 VDD1.n30 VDD1.n17 0.155672
R739 VDD1.n30 VDD1.n29 0.155672
R740 VDD1.n29 VDD1.n21 0.155672
R741 VDD1.n100 VDD1.n92 0.155672
R742 VDD1.n101 VDD1.n100 0.155672
R743 VDD1.n101 VDD1.n88 0.155672
R744 VDD1.n108 VDD1.n88 0.155672
R745 VDD1.n109 VDD1.n108 0.155672
R746 VDD1.n109 VDD1.n84 0.155672
R747 VDD1.n116 VDD1.n84 0.155672
R748 VDD1.n117 VDD1.n116 0.155672
R749 VDD1.n117 VDD1.n80 0.155672
R750 VDD1.n124 VDD1.n80 0.155672
R751 VDD1.n125 VDD1.n124 0.155672
R752 VDD1.n125 VDD1.n76 0.155672
R753 VDD1.n132 VDD1.n76 0.155672
R754 VDD1.n133 VDD1.n132 0.155672
R755 VDD1.n133 VDD1.n72 0.155672
R756 VDD1.n140 VDD1.n72 0.155672
R757 B.n924 B.n923 585
R758 B.n925 B.n924 585
R759 B.n347 B.n145 585
R760 B.n346 B.n345 585
R761 B.n344 B.n343 585
R762 B.n342 B.n341 585
R763 B.n340 B.n339 585
R764 B.n338 B.n337 585
R765 B.n336 B.n335 585
R766 B.n334 B.n333 585
R767 B.n332 B.n331 585
R768 B.n330 B.n329 585
R769 B.n328 B.n327 585
R770 B.n326 B.n325 585
R771 B.n324 B.n323 585
R772 B.n322 B.n321 585
R773 B.n320 B.n319 585
R774 B.n318 B.n317 585
R775 B.n316 B.n315 585
R776 B.n314 B.n313 585
R777 B.n312 B.n311 585
R778 B.n310 B.n309 585
R779 B.n308 B.n307 585
R780 B.n306 B.n305 585
R781 B.n304 B.n303 585
R782 B.n302 B.n301 585
R783 B.n300 B.n299 585
R784 B.n298 B.n297 585
R785 B.n296 B.n295 585
R786 B.n294 B.n293 585
R787 B.n292 B.n291 585
R788 B.n290 B.n289 585
R789 B.n288 B.n287 585
R790 B.n286 B.n285 585
R791 B.n284 B.n283 585
R792 B.n282 B.n281 585
R793 B.n280 B.n279 585
R794 B.n278 B.n277 585
R795 B.n276 B.n275 585
R796 B.n274 B.n273 585
R797 B.n272 B.n271 585
R798 B.n270 B.n269 585
R799 B.n268 B.n267 585
R800 B.n266 B.n265 585
R801 B.n264 B.n263 585
R802 B.n262 B.n261 585
R803 B.n260 B.n259 585
R804 B.n257 B.n256 585
R805 B.n255 B.n254 585
R806 B.n253 B.n252 585
R807 B.n251 B.n250 585
R808 B.n249 B.n248 585
R809 B.n247 B.n246 585
R810 B.n245 B.n244 585
R811 B.n243 B.n242 585
R812 B.n241 B.n240 585
R813 B.n239 B.n238 585
R814 B.n237 B.n236 585
R815 B.n235 B.n234 585
R816 B.n233 B.n232 585
R817 B.n231 B.n230 585
R818 B.n229 B.n228 585
R819 B.n227 B.n226 585
R820 B.n225 B.n224 585
R821 B.n223 B.n222 585
R822 B.n221 B.n220 585
R823 B.n219 B.n218 585
R824 B.n217 B.n216 585
R825 B.n215 B.n214 585
R826 B.n213 B.n212 585
R827 B.n211 B.n210 585
R828 B.n209 B.n208 585
R829 B.n207 B.n206 585
R830 B.n205 B.n204 585
R831 B.n203 B.n202 585
R832 B.n201 B.n200 585
R833 B.n199 B.n198 585
R834 B.n197 B.n196 585
R835 B.n195 B.n194 585
R836 B.n193 B.n192 585
R837 B.n191 B.n190 585
R838 B.n189 B.n188 585
R839 B.n187 B.n186 585
R840 B.n185 B.n184 585
R841 B.n183 B.n182 585
R842 B.n181 B.n180 585
R843 B.n179 B.n178 585
R844 B.n177 B.n176 585
R845 B.n175 B.n174 585
R846 B.n173 B.n172 585
R847 B.n171 B.n170 585
R848 B.n169 B.n168 585
R849 B.n167 B.n166 585
R850 B.n165 B.n164 585
R851 B.n163 B.n162 585
R852 B.n161 B.n160 585
R853 B.n159 B.n158 585
R854 B.n157 B.n156 585
R855 B.n155 B.n154 585
R856 B.n153 B.n152 585
R857 B.n95 B.n94 585
R858 B.n928 B.n927 585
R859 B.n922 B.n146 585
R860 B.n146 B.n92 585
R861 B.n921 B.n91 585
R862 B.n932 B.n91 585
R863 B.n920 B.n90 585
R864 B.n933 B.n90 585
R865 B.n919 B.n89 585
R866 B.n934 B.n89 585
R867 B.n918 B.n917 585
R868 B.n917 B.n85 585
R869 B.n916 B.n84 585
R870 B.n940 B.n84 585
R871 B.n915 B.n83 585
R872 B.n941 B.n83 585
R873 B.n914 B.n82 585
R874 B.n942 B.n82 585
R875 B.n913 B.n912 585
R876 B.n912 B.n81 585
R877 B.n911 B.n77 585
R878 B.n948 B.n77 585
R879 B.n910 B.n76 585
R880 B.n949 B.n76 585
R881 B.n909 B.n75 585
R882 B.n950 B.n75 585
R883 B.n908 B.n907 585
R884 B.n907 B.n71 585
R885 B.n906 B.n70 585
R886 B.n956 B.n70 585
R887 B.n905 B.n69 585
R888 B.n957 B.n69 585
R889 B.n904 B.n68 585
R890 B.n958 B.n68 585
R891 B.n903 B.n902 585
R892 B.n902 B.n64 585
R893 B.n901 B.n63 585
R894 B.n964 B.n63 585
R895 B.n900 B.n62 585
R896 B.n965 B.n62 585
R897 B.n899 B.n61 585
R898 B.n966 B.n61 585
R899 B.n898 B.n897 585
R900 B.n897 B.n57 585
R901 B.n896 B.n56 585
R902 B.n972 B.n56 585
R903 B.n895 B.n55 585
R904 B.n973 B.n55 585
R905 B.n894 B.n54 585
R906 B.n974 B.n54 585
R907 B.n893 B.n892 585
R908 B.n892 B.n50 585
R909 B.n891 B.n49 585
R910 B.n980 B.n49 585
R911 B.n890 B.n48 585
R912 B.n981 B.n48 585
R913 B.n889 B.n47 585
R914 B.n982 B.n47 585
R915 B.n888 B.n887 585
R916 B.n887 B.n43 585
R917 B.n886 B.n42 585
R918 B.n988 B.n42 585
R919 B.n885 B.n41 585
R920 B.n989 B.n41 585
R921 B.n884 B.n40 585
R922 B.n990 B.n40 585
R923 B.n883 B.n882 585
R924 B.n882 B.n36 585
R925 B.n881 B.n35 585
R926 B.n996 B.n35 585
R927 B.n880 B.n34 585
R928 B.n997 B.n34 585
R929 B.n879 B.n33 585
R930 B.n998 B.n33 585
R931 B.n878 B.n877 585
R932 B.n877 B.n29 585
R933 B.n876 B.n28 585
R934 B.n1004 B.n28 585
R935 B.n875 B.n27 585
R936 B.n1005 B.n27 585
R937 B.n874 B.n26 585
R938 B.n1006 B.n26 585
R939 B.n873 B.n872 585
R940 B.n872 B.n22 585
R941 B.n871 B.n21 585
R942 B.n1012 B.n21 585
R943 B.n870 B.n20 585
R944 B.n1013 B.n20 585
R945 B.n869 B.n19 585
R946 B.n1014 B.n19 585
R947 B.n868 B.n867 585
R948 B.n867 B.n18 585
R949 B.n866 B.n14 585
R950 B.n1020 B.n14 585
R951 B.n865 B.n13 585
R952 B.n1021 B.n13 585
R953 B.n864 B.n12 585
R954 B.n1022 B.n12 585
R955 B.n863 B.n862 585
R956 B.n862 B.n8 585
R957 B.n861 B.n7 585
R958 B.n1028 B.n7 585
R959 B.n860 B.n6 585
R960 B.n1029 B.n6 585
R961 B.n859 B.n5 585
R962 B.n1030 B.n5 585
R963 B.n858 B.n857 585
R964 B.n857 B.n4 585
R965 B.n856 B.n348 585
R966 B.n856 B.n855 585
R967 B.n846 B.n349 585
R968 B.n350 B.n349 585
R969 B.n848 B.n847 585
R970 B.n849 B.n848 585
R971 B.n845 B.n355 585
R972 B.n355 B.n354 585
R973 B.n844 B.n843 585
R974 B.n843 B.n842 585
R975 B.n357 B.n356 585
R976 B.n835 B.n357 585
R977 B.n834 B.n833 585
R978 B.n836 B.n834 585
R979 B.n832 B.n362 585
R980 B.n362 B.n361 585
R981 B.n831 B.n830 585
R982 B.n830 B.n829 585
R983 B.n364 B.n363 585
R984 B.n365 B.n364 585
R985 B.n822 B.n821 585
R986 B.n823 B.n822 585
R987 B.n820 B.n370 585
R988 B.n370 B.n369 585
R989 B.n819 B.n818 585
R990 B.n818 B.n817 585
R991 B.n372 B.n371 585
R992 B.n373 B.n372 585
R993 B.n810 B.n809 585
R994 B.n811 B.n810 585
R995 B.n808 B.n378 585
R996 B.n378 B.n377 585
R997 B.n807 B.n806 585
R998 B.n806 B.n805 585
R999 B.n380 B.n379 585
R1000 B.n381 B.n380 585
R1001 B.n798 B.n797 585
R1002 B.n799 B.n798 585
R1003 B.n796 B.n386 585
R1004 B.n386 B.n385 585
R1005 B.n795 B.n794 585
R1006 B.n794 B.n793 585
R1007 B.n388 B.n387 585
R1008 B.n389 B.n388 585
R1009 B.n786 B.n785 585
R1010 B.n787 B.n786 585
R1011 B.n784 B.n394 585
R1012 B.n394 B.n393 585
R1013 B.n783 B.n782 585
R1014 B.n782 B.n781 585
R1015 B.n396 B.n395 585
R1016 B.n397 B.n396 585
R1017 B.n774 B.n773 585
R1018 B.n775 B.n774 585
R1019 B.n772 B.n401 585
R1020 B.n405 B.n401 585
R1021 B.n771 B.n770 585
R1022 B.n770 B.n769 585
R1023 B.n403 B.n402 585
R1024 B.n404 B.n403 585
R1025 B.n762 B.n761 585
R1026 B.n763 B.n762 585
R1027 B.n760 B.n410 585
R1028 B.n410 B.n409 585
R1029 B.n759 B.n758 585
R1030 B.n758 B.n757 585
R1031 B.n412 B.n411 585
R1032 B.n413 B.n412 585
R1033 B.n750 B.n749 585
R1034 B.n751 B.n750 585
R1035 B.n748 B.n418 585
R1036 B.n418 B.n417 585
R1037 B.n747 B.n746 585
R1038 B.n746 B.n745 585
R1039 B.n420 B.n419 585
R1040 B.n421 B.n420 585
R1041 B.n738 B.n737 585
R1042 B.n739 B.n738 585
R1043 B.n736 B.n426 585
R1044 B.n426 B.n425 585
R1045 B.n735 B.n734 585
R1046 B.n734 B.n733 585
R1047 B.n428 B.n427 585
R1048 B.n726 B.n428 585
R1049 B.n725 B.n724 585
R1050 B.n727 B.n725 585
R1051 B.n723 B.n433 585
R1052 B.n433 B.n432 585
R1053 B.n722 B.n721 585
R1054 B.n721 B.n720 585
R1055 B.n435 B.n434 585
R1056 B.n436 B.n435 585
R1057 B.n713 B.n712 585
R1058 B.n714 B.n713 585
R1059 B.n711 B.n441 585
R1060 B.n441 B.n440 585
R1061 B.n710 B.n709 585
R1062 B.n709 B.n708 585
R1063 B.n443 B.n442 585
R1064 B.n444 B.n443 585
R1065 B.n704 B.n703 585
R1066 B.n447 B.n446 585
R1067 B.n700 B.n699 585
R1068 B.n701 B.n700 585
R1069 B.n698 B.n497 585
R1070 B.n697 B.n696 585
R1071 B.n695 B.n694 585
R1072 B.n693 B.n692 585
R1073 B.n691 B.n690 585
R1074 B.n689 B.n688 585
R1075 B.n687 B.n686 585
R1076 B.n685 B.n684 585
R1077 B.n683 B.n682 585
R1078 B.n681 B.n680 585
R1079 B.n679 B.n678 585
R1080 B.n677 B.n676 585
R1081 B.n675 B.n674 585
R1082 B.n673 B.n672 585
R1083 B.n671 B.n670 585
R1084 B.n669 B.n668 585
R1085 B.n667 B.n666 585
R1086 B.n665 B.n664 585
R1087 B.n663 B.n662 585
R1088 B.n661 B.n660 585
R1089 B.n659 B.n658 585
R1090 B.n657 B.n656 585
R1091 B.n655 B.n654 585
R1092 B.n653 B.n652 585
R1093 B.n651 B.n650 585
R1094 B.n649 B.n648 585
R1095 B.n647 B.n646 585
R1096 B.n645 B.n644 585
R1097 B.n643 B.n642 585
R1098 B.n641 B.n640 585
R1099 B.n639 B.n638 585
R1100 B.n637 B.n636 585
R1101 B.n635 B.n634 585
R1102 B.n633 B.n632 585
R1103 B.n631 B.n630 585
R1104 B.n629 B.n628 585
R1105 B.n627 B.n626 585
R1106 B.n625 B.n624 585
R1107 B.n623 B.n622 585
R1108 B.n621 B.n620 585
R1109 B.n619 B.n618 585
R1110 B.n617 B.n616 585
R1111 B.n615 B.n614 585
R1112 B.n612 B.n611 585
R1113 B.n610 B.n609 585
R1114 B.n608 B.n607 585
R1115 B.n606 B.n605 585
R1116 B.n604 B.n603 585
R1117 B.n602 B.n601 585
R1118 B.n600 B.n599 585
R1119 B.n598 B.n597 585
R1120 B.n596 B.n595 585
R1121 B.n594 B.n593 585
R1122 B.n592 B.n591 585
R1123 B.n590 B.n589 585
R1124 B.n588 B.n587 585
R1125 B.n586 B.n585 585
R1126 B.n584 B.n583 585
R1127 B.n582 B.n581 585
R1128 B.n580 B.n579 585
R1129 B.n578 B.n577 585
R1130 B.n576 B.n575 585
R1131 B.n574 B.n573 585
R1132 B.n572 B.n571 585
R1133 B.n570 B.n569 585
R1134 B.n568 B.n567 585
R1135 B.n566 B.n565 585
R1136 B.n564 B.n563 585
R1137 B.n562 B.n561 585
R1138 B.n560 B.n559 585
R1139 B.n558 B.n557 585
R1140 B.n556 B.n555 585
R1141 B.n554 B.n553 585
R1142 B.n552 B.n551 585
R1143 B.n550 B.n549 585
R1144 B.n548 B.n547 585
R1145 B.n546 B.n545 585
R1146 B.n544 B.n543 585
R1147 B.n542 B.n541 585
R1148 B.n540 B.n539 585
R1149 B.n538 B.n537 585
R1150 B.n536 B.n535 585
R1151 B.n534 B.n533 585
R1152 B.n532 B.n531 585
R1153 B.n530 B.n529 585
R1154 B.n528 B.n527 585
R1155 B.n526 B.n525 585
R1156 B.n524 B.n523 585
R1157 B.n522 B.n521 585
R1158 B.n520 B.n519 585
R1159 B.n518 B.n517 585
R1160 B.n516 B.n515 585
R1161 B.n514 B.n513 585
R1162 B.n512 B.n511 585
R1163 B.n510 B.n509 585
R1164 B.n508 B.n507 585
R1165 B.n506 B.n505 585
R1166 B.n504 B.n503 585
R1167 B.n705 B.n445 585
R1168 B.n445 B.n444 585
R1169 B.n707 B.n706 585
R1170 B.n708 B.n707 585
R1171 B.n439 B.n438 585
R1172 B.n440 B.n439 585
R1173 B.n716 B.n715 585
R1174 B.n715 B.n714 585
R1175 B.n717 B.n437 585
R1176 B.n437 B.n436 585
R1177 B.n719 B.n718 585
R1178 B.n720 B.n719 585
R1179 B.n431 B.n430 585
R1180 B.n432 B.n431 585
R1181 B.n729 B.n728 585
R1182 B.n728 B.n727 585
R1183 B.n730 B.n429 585
R1184 B.n726 B.n429 585
R1185 B.n732 B.n731 585
R1186 B.n733 B.n732 585
R1187 B.n424 B.n423 585
R1188 B.n425 B.n424 585
R1189 B.n741 B.n740 585
R1190 B.n740 B.n739 585
R1191 B.n742 B.n422 585
R1192 B.n422 B.n421 585
R1193 B.n744 B.n743 585
R1194 B.n745 B.n744 585
R1195 B.n416 B.n415 585
R1196 B.n417 B.n416 585
R1197 B.n753 B.n752 585
R1198 B.n752 B.n751 585
R1199 B.n754 B.n414 585
R1200 B.n414 B.n413 585
R1201 B.n756 B.n755 585
R1202 B.n757 B.n756 585
R1203 B.n408 B.n407 585
R1204 B.n409 B.n408 585
R1205 B.n765 B.n764 585
R1206 B.n764 B.n763 585
R1207 B.n766 B.n406 585
R1208 B.n406 B.n404 585
R1209 B.n768 B.n767 585
R1210 B.n769 B.n768 585
R1211 B.n400 B.n399 585
R1212 B.n405 B.n400 585
R1213 B.n777 B.n776 585
R1214 B.n776 B.n775 585
R1215 B.n778 B.n398 585
R1216 B.n398 B.n397 585
R1217 B.n780 B.n779 585
R1218 B.n781 B.n780 585
R1219 B.n392 B.n391 585
R1220 B.n393 B.n392 585
R1221 B.n789 B.n788 585
R1222 B.n788 B.n787 585
R1223 B.n790 B.n390 585
R1224 B.n390 B.n389 585
R1225 B.n792 B.n791 585
R1226 B.n793 B.n792 585
R1227 B.n384 B.n383 585
R1228 B.n385 B.n384 585
R1229 B.n801 B.n800 585
R1230 B.n800 B.n799 585
R1231 B.n802 B.n382 585
R1232 B.n382 B.n381 585
R1233 B.n804 B.n803 585
R1234 B.n805 B.n804 585
R1235 B.n376 B.n375 585
R1236 B.n377 B.n376 585
R1237 B.n813 B.n812 585
R1238 B.n812 B.n811 585
R1239 B.n814 B.n374 585
R1240 B.n374 B.n373 585
R1241 B.n816 B.n815 585
R1242 B.n817 B.n816 585
R1243 B.n368 B.n367 585
R1244 B.n369 B.n368 585
R1245 B.n825 B.n824 585
R1246 B.n824 B.n823 585
R1247 B.n826 B.n366 585
R1248 B.n366 B.n365 585
R1249 B.n828 B.n827 585
R1250 B.n829 B.n828 585
R1251 B.n360 B.n359 585
R1252 B.n361 B.n360 585
R1253 B.n838 B.n837 585
R1254 B.n837 B.n836 585
R1255 B.n839 B.n358 585
R1256 B.n835 B.n358 585
R1257 B.n841 B.n840 585
R1258 B.n842 B.n841 585
R1259 B.n353 B.n352 585
R1260 B.n354 B.n353 585
R1261 B.n851 B.n850 585
R1262 B.n850 B.n849 585
R1263 B.n852 B.n351 585
R1264 B.n351 B.n350 585
R1265 B.n854 B.n853 585
R1266 B.n855 B.n854 585
R1267 B.n2 B.n0 585
R1268 B.n4 B.n2 585
R1269 B.n3 B.n1 585
R1270 B.n1029 B.n3 585
R1271 B.n1027 B.n1026 585
R1272 B.n1028 B.n1027 585
R1273 B.n1025 B.n9 585
R1274 B.n9 B.n8 585
R1275 B.n1024 B.n1023 585
R1276 B.n1023 B.n1022 585
R1277 B.n11 B.n10 585
R1278 B.n1021 B.n11 585
R1279 B.n1019 B.n1018 585
R1280 B.n1020 B.n1019 585
R1281 B.n1017 B.n15 585
R1282 B.n18 B.n15 585
R1283 B.n1016 B.n1015 585
R1284 B.n1015 B.n1014 585
R1285 B.n17 B.n16 585
R1286 B.n1013 B.n17 585
R1287 B.n1011 B.n1010 585
R1288 B.n1012 B.n1011 585
R1289 B.n1009 B.n23 585
R1290 B.n23 B.n22 585
R1291 B.n1008 B.n1007 585
R1292 B.n1007 B.n1006 585
R1293 B.n25 B.n24 585
R1294 B.n1005 B.n25 585
R1295 B.n1003 B.n1002 585
R1296 B.n1004 B.n1003 585
R1297 B.n1001 B.n30 585
R1298 B.n30 B.n29 585
R1299 B.n1000 B.n999 585
R1300 B.n999 B.n998 585
R1301 B.n32 B.n31 585
R1302 B.n997 B.n32 585
R1303 B.n995 B.n994 585
R1304 B.n996 B.n995 585
R1305 B.n993 B.n37 585
R1306 B.n37 B.n36 585
R1307 B.n992 B.n991 585
R1308 B.n991 B.n990 585
R1309 B.n39 B.n38 585
R1310 B.n989 B.n39 585
R1311 B.n987 B.n986 585
R1312 B.n988 B.n987 585
R1313 B.n985 B.n44 585
R1314 B.n44 B.n43 585
R1315 B.n984 B.n983 585
R1316 B.n983 B.n982 585
R1317 B.n46 B.n45 585
R1318 B.n981 B.n46 585
R1319 B.n979 B.n978 585
R1320 B.n980 B.n979 585
R1321 B.n977 B.n51 585
R1322 B.n51 B.n50 585
R1323 B.n976 B.n975 585
R1324 B.n975 B.n974 585
R1325 B.n53 B.n52 585
R1326 B.n973 B.n53 585
R1327 B.n971 B.n970 585
R1328 B.n972 B.n971 585
R1329 B.n969 B.n58 585
R1330 B.n58 B.n57 585
R1331 B.n968 B.n967 585
R1332 B.n967 B.n966 585
R1333 B.n60 B.n59 585
R1334 B.n965 B.n60 585
R1335 B.n963 B.n962 585
R1336 B.n964 B.n963 585
R1337 B.n961 B.n65 585
R1338 B.n65 B.n64 585
R1339 B.n960 B.n959 585
R1340 B.n959 B.n958 585
R1341 B.n67 B.n66 585
R1342 B.n957 B.n67 585
R1343 B.n955 B.n954 585
R1344 B.n956 B.n955 585
R1345 B.n953 B.n72 585
R1346 B.n72 B.n71 585
R1347 B.n952 B.n951 585
R1348 B.n951 B.n950 585
R1349 B.n74 B.n73 585
R1350 B.n949 B.n74 585
R1351 B.n947 B.n946 585
R1352 B.n948 B.n947 585
R1353 B.n945 B.n78 585
R1354 B.n81 B.n78 585
R1355 B.n944 B.n943 585
R1356 B.n943 B.n942 585
R1357 B.n80 B.n79 585
R1358 B.n941 B.n80 585
R1359 B.n939 B.n938 585
R1360 B.n940 B.n939 585
R1361 B.n937 B.n86 585
R1362 B.n86 B.n85 585
R1363 B.n936 B.n935 585
R1364 B.n935 B.n934 585
R1365 B.n88 B.n87 585
R1366 B.n933 B.n88 585
R1367 B.n931 B.n930 585
R1368 B.n932 B.n931 585
R1369 B.n929 B.n93 585
R1370 B.n93 B.n92 585
R1371 B.n1032 B.n1031 585
R1372 B.n1031 B.n1030 585
R1373 B.n703 B.n445 468.476
R1374 B.n927 B.n93 468.476
R1375 B.n503 B.n443 468.476
R1376 B.n924 B.n146 468.476
R1377 B.n500 B.t12 375.832
R1378 B.n147 B.t7 375.832
R1379 B.n498 B.t15 375.832
R1380 B.n149 B.t17 375.832
R1381 B.n500 B.t9 306.115
R1382 B.n498 B.t13 306.115
R1383 B.n149 B.t16 306.115
R1384 B.n147 B.t5 306.115
R1385 B.n501 B.t11 305.238
R1386 B.n148 B.t8 305.238
R1387 B.n499 B.t14 305.238
R1388 B.n150 B.t18 305.238
R1389 B.n925 B.n144 256.663
R1390 B.n925 B.n143 256.663
R1391 B.n925 B.n142 256.663
R1392 B.n925 B.n141 256.663
R1393 B.n925 B.n140 256.663
R1394 B.n925 B.n139 256.663
R1395 B.n925 B.n138 256.663
R1396 B.n925 B.n137 256.663
R1397 B.n925 B.n136 256.663
R1398 B.n925 B.n135 256.663
R1399 B.n925 B.n134 256.663
R1400 B.n925 B.n133 256.663
R1401 B.n925 B.n132 256.663
R1402 B.n925 B.n131 256.663
R1403 B.n925 B.n130 256.663
R1404 B.n925 B.n129 256.663
R1405 B.n925 B.n128 256.663
R1406 B.n925 B.n127 256.663
R1407 B.n925 B.n126 256.663
R1408 B.n925 B.n125 256.663
R1409 B.n925 B.n124 256.663
R1410 B.n925 B.n123 256.663
R1411 B.n925 B.n122 256.663
R1412 B.n925 B.n121 256.663
R1413 B.n925 B.n120 256.663
R1414 B.n925 B.n119 256.663
R1415 B.n925 B.n118 256.663
R1416 B.n925 B.n117 256.663
R1417 B.n925 B.n116 256.663
R1418 B.n925 B.n115 256.663
R1419 B.n925 B.n114 256.663
R1420 B.n925 B.n113 256.663
R1421 B.n925 B.n112 256.663
R1422 B.n925 B.n111 256.663
R1423 B.n925 B.n110 256.663
R1424 B.n925 B.n109 256.663
R1425 B.n925 B.n108 256.663
R1426 B.n925 B.n107 256.663
R1427 B.n925 B.n106 256.663
R1428 B.n925 B.n105 256.663
R1429 B.n925 B.n104 256.663
R1430 B.n925 B.n103 256.663
R1431 B.n925 B.n102 256.663
R1432 B.n925 B.n101 256.663
R1433 B.n925 B.n100 256.663
R1434 B.n925 B.n99 256.663
R1435 B.n925 B.n98 256.663
R1436 B.n925 B.n97 256.663
R1437 B.n925 B.n96 256.663
R1438 B.n926 B.n925 256.663
R1439 B.n702 B.n701 256.663
R1440 B.n701 B.n448 256.663
R1441 B.n701 B.n449 256.663
R1442 B.n701 B.n450 256.663
R1443 B.n701 B.n451 256.663
R1444 B.n701 B.n452 256.663
R1445 B.n701 B.n453 256.663
R1446 B.n701 B.n454 256.663
R1447 B.n701 B.n455 256.663
R1448 B.n701 B.n456 256.663
R1449 B.n701 B.n457 256.663
R1450 B.n701 B.n458 256.663
R1451 B.n701 B.n459 256.663
R1452 B.n701 B.n460 256.663
R1453 B.n701 B.n461 256.663
R1454 B.n701 B.n462 256.663
R1455 B.n701 B.n463 256.663
R1456 B.n701 B.n464 256.663
R1457 B.n701 B.n465 256.663
R1458 B.n701 B.n466 256.663
R1459 B.n701 B.n467 256.663
R1460 B.n701 B.n468 256.663
R1461 B.n701 B.n469 256.663
R1462 B.n701 B.n470 256.663
R1463 B.n701 B.n471 256.663
R1464 B.n701 B.n472 256.663
R1465 B.n701 B.n473 256.663
R1466 B.n701 B.n474 256.663
R1467 B.n701 B.n475 256.663
R1468 B.n701 B.n476 256.663
R1469 B.n701 B.n477 256.663
R1470 B.n701 B.n478 256.663
R1471 B.n701 B.n479 256.663
R1472 B.n701 B.n480 256.663
R1473 B.n701 B.n481 256.663
R1474 B.n701 B.n482 256.663
R1475 B.n701 B.n483 256.663
R1476 B.n701 B.n484 256.663
R1477 B.n701 B.n485 256.663
R1478 B.n701 B.n486 256.663
R1479 B.n701 B.n487 256.663
R1480 B.n701 B.n488 256.663
R1481 B.n701 B.n489 256.663
R1482 B.n701 B.n490 256.663
R1483 B.n701 B.n491 256.663
R1484 B.n701 B.n492 256.663
R1485 B.n701 B.n493 256.663
R1486 B.n701 B.n494 256.663
R1487 B.n701 B.n495 256.663
R1488 B.n701 B.n496 256.663
R1489 B.n707 B.n445 163.367
R1490 B.n707 B.n439 163.367
R1491 B.n715 B.n439 163.367
R1492 B.n715 B.n437 163.367
R1493 B.n719 B.n437 163.367
R1494 B.n719 B.n431 163.367
R1495 B.n728 B.n431 163.367
R1496 B.n728 B.n429 163.367
R1497 B.n732 B.n429 163.367
R1498 B.n732 B.n424 163.367
R1499 B.n740 B.n424 163.367
R1500 B.n740 B.n422 163.367
R1501 B.n744 B.n422 163.367
R1502 B.n744 B.n416 163.367
R1503 B.n752 B.n416 163.367
R1504 B.n752 B.n414 163.367
R1505 B.n756 B.n414 163.367
R1506 B.n756 B.n408 163.367
R1507 B.n764 B.n408 163.367
R1508 B.n764 B.n406 163.367
R1509 B.n768 B.n406 163.367
R1510 B.n768 B.n400 163.367
R1511 B.n776 B.n400 163.367
R1512 B.n776 B.n398 163.367
R1513 B.n780 B.n398 163.367
R1514 B.n780 B.n392 163.367
R1515 B.n788 B.n392 163.367
R1516 B.n788 B.n390 163.367
R1517 B.n792 B.n390 163.367
R1518 B.n792 B.n384 163.367
R1519 B.n800 B.n384 163.367
R1520 B.n800 B.n382 163.367
R1521 B.n804 B.n382 163.367
R1522 B.n804 B.n376 163.367
R1523 B.n812 B.n376 163.367
R1524 B.n812 B.n374 163.367
R1525 B.n816 B.n374 163.367
R1526 B.n816 B.n368 163.367
R1527 B.n824 B.n368 163.367
R1528 B.n824 B.n366 163.367
R1529 B.n828 B.n366 163.367
R1530 B.n828 B.n360 163.367
R1531 B.n837 B.n360 163.367
R1532 B.n837 B.n358 163.367
R1533 B.n841 B.n358 163.367
R1534 B.n841 B.n353 163.367
R1535 B.n850 B.n353 163.367
R1536 B.n850 B.n351 163.367
R1537 B.n854 B.n351 163.367
R1538 B.n854 B.n2 163.367
R1539 B.n1031 B.n2 163.367
R1540 B.n1031 B.n3 163.367
R1541 B.n1027 B.n3 163.367
R1542 B.n1027 B.n9 163.367
R1543 B.n1023 B.n9 163.367
R1544 B.n1023 B.n11 163.367
R1545 B.n1019 B.n11 163.367
R1546 B.n1019 B.n15 163.367
R1547 B.n1015 B.n15 163.367
R1548 B.n1015 B.n17 163.367
R1549 B.n1011 B.n17 163.367
R1550 B.n1011 B.n23 163.367
R1551 B.n1007 B.n23 163.367
R1552 B.n1007 B.n25 163.367
R1553 B.n1003 B.n25 163.367
R1554 B.n1003 B.n30 163.367
R1555 B.n999 B.n30 163.367
R1556 B.n999 B.n32 163.367
R1557 B.n995 B.n32 163.367
R1558 B.n995 B.n37 163.367
R1559 B.n991 B.n37 163.367
R1560 B.n991 B.n39 163.367
R1561 B.n987 B.n39 163.367
R1562 B.n987 B.n44 163.367
R1563 B.n983 B.n44 163.367
R1564 B.n983 B.n46 163.367
R1565 B.n979 B.n46 163.367
R1566 B.n979 B.n51 163.367
R1567 B.n975 B.n51 163.367
R1568 B.n975 B.n53 163.367
R1569 B.n971 B.n53 163.367
R1570 B.n971 B.n58 163.367
R1571 B.n967 B.n58 163.367
R1572 B.n967 B.n60 163.367
R1573 B.n963 B.n60 163.367
R1574 B.n963 B.n65 163.367
R1575 B.n959 B.n65 163.367
R1576 B.n959 B.n67 163.367
R1577 B.n955 B.n67 163.367
R1578 B.n955 B.n72 163.367
R1579 B.n951 B.n72 163.367
R1580 B.n951 B.n74 163.367
R1581 B.n947 B.n74 163.367
R1582 B.n947 B.n78 163.367
R1583 B.n943 B.n78 163.367
R1584 B.n943 B.n80 163.367
R1585 B.n939 B.n80 163.367
R1586 B.n939 B.n86 163.367
R1587 B.n935 B.n86 163.367
R1588 B.n935 B.n88 163.367
R1589 B.n931 B.n88 163.367
R1590 B.n931 B.n93 163.367
R1591 B.n700 B.n447 163.367
R1592 B.n700 B.n497 163.367
R1593 B.n696 B.n695 163.367
R1594 B.n692 B.n691 163.367
R1595 B.n688 B.n687 163.367
R1596 B.n684 B.n683 163.367
R1597 B.n680 B.n679 163.367
R1598 B.n676 B.n675 163.367
R1599 B.n672 B.n671 163.367
R1600 B.n668 B.n667 163.367
R1601 B.n664 B.n663 163.367
R1602 B.n660 B.n659 163.367
R1603 B.n656 B.n655 163.367
R1604 B.n652 B.n651 163.367
R1605 B.n648 B.n647 163.367
R1606 B.n644 B.n643 163.367
R1607 B.n640 B.n639 163.367
R1608 B.n636 B.n635 163.367
R1609 B.n632 B.n631 163.367
R1610 B.n628 B.n627 163.367
R1611 B.n624 B.n623 163.367
R1612 B.n620 B.n619 163.367
R1613 B.n616 B.n615 163.367
R1614 B.n611 B.n610 163.367
R1615 B.n607 B.n606 163.367
R1616 B.n603 B.n602 163.367
R1617 B.n599 B.n598 163.367
R1618 B.n595 B.n594 163.367
R1619 B.n591 B.n590 163.367
R1620 B.n587 B.n586 163.367
R1621 B.n583 B.n582 163.367
R1622 B.n579 B.n578 163.367
R1623 B.n575 B.n574 163.367
R1624 B.n571 B.n570 163.367
R1625 B.n567 B.n566 163.367
R1626 B.n563 B.n562 163.367
R1627 B.n559 B.n558 163.367
R1628 B.n555 B.n554 163.367
R1629 B.n551 B.n550 163.367
R1630 B.n547 B.n546 163.367
R1631 B.n543 B.n542 163.367
R1632 B.n539 B.n538 163.367
R1633 B.n535 B.n534 163.367
R1634 B.n531 B.n530 163.367
R1635 B.n527 B.n526 163.367
R1636 B.n523 B.n522 163.367
R1637 B.n519 B.n518 163.367
R1638 B.n515 B.n514 163.367
R1639 B.n511 B.n510 163.367
R1640 B.n507 B.n506 163.367
R1641 B.n709 B.n443 163.367
R1642 B.n709 B.n441 163.367
R1643 B.n713 B.n441 163.367
R1644 B.n713 B.n435 163.367
R1645 B.n721 B.n435 163.367
R1646 B.n721 B.n433 163.367
R1647 B.n725 B.n433 163.367
R1648 B.n725 B.n428 163.367
R1649 B.n734 B.n428 163.367
R1650 B.n734 B.n426 163.367
R1651 B.n738 B.n426 163.367
R1652 B.n738 B.n420 163.367
R1653 B.n746 B.n420 163.367
R1654 B.n746 B.n418 163.367
R1655 B.n750 B.n418 163.367
R1656 B.n750 B.n412 163.367
R1657 B.n758 B.n412 163.367
R1658 B.n758 B.n410 163.367
R1659 B.n762 B.n410 163.367
R1660 B.n762 B.n403 163.367
R1661 B.n770 B.n403 163.367
R1662 B.n770 B.n401 163.367
R1663 B.n774 B.n401 163.367
R1664 B.n774 B.n396 163.367
R1665 B.n782 B.n396 163.367
R1666 B.n782 B.n394 163.367
R1667 B.n786 B.n394 163.367
R1668 B.n786 B.n388 163.367
R1669 B.n794 B.n388 163.367
R1670 B.n794 B.n386 163.367
R1671 B.n798 B.n386 163.367
R1672 B.n798 B.n380 163.367
R1673 B.n806 B.n380 163.367
R1674 B.n806 B.n378 163.367
R1675 B.n810 B.n378 163.367
R1676 B.n810 B.n372 163.367
R1677 B.n818 B.n372 163.367
R1678 B.n818 B.n370 163.367
R1679 B.n822 B.n370 163.367
R1680 B.n822 B.n364 163.367
R1681 B.n830 B.n364 163.367
R1682 B.n830 B.n362 163.367
R1683 B.n834 B.n362 163.367
R1684 B.n834 B.n357 163.367
R1685 B.n843 B.n357 163.367
R1686 B.n843 B.n355 163.367
R1687 B.n848 B.n355 163.367
R1688 B.n848 B.n349 163.367
R1689 B.n856 B.n349 163.367
R1690 B.n857 B.n856 163.367
R1691 B.n857 B.n5 163.367
R1692 B.n6 B.n5 163.367
R1693 B.n7 B.n6 163.367
R1694 B.n862 B.n7 163.367
R1695 B.n862 B.n12 163.367
R1696 B.n13 B.n12 163.367
R1697 B.n14 B.n13 163.367
R1698 B.n867 B.n14 163.367
R1699 B.n867 B.n19 163.367
R1700 B.n20 B.n19 163.367
R1701 B.n21 B.n20 163.367
R1702 B.n872 B.n21 163.367
R1703 B.n872 B.n26 163.367
R1704 B.n27 B.n26 163.367
R1705 B.n28 B.n27 163.367
R1706 B.n877 B.n28 163.367
R1707 B.n877 B.n33 163.367
R1708 B.n34 B.n33 163.367
R1709 B.n35 B.n34 163.367
R1710 B.n882 B.n35 163.367
R1711 B.n882 B.n40 163.367
R1712 B.n41 B.n40 163.367
R1713 B.n42 B.n41 163.367
R1714 B.n887 B.n42 163.367
R1715 B.n887 B.n47 163.367
R1716 B.n48 B.n47 163.367
R1717 B.n49 B.n48 163.367
R1718 B.n892 B.n49 163.367
R1719 B.n892 B.n54 163.367
R1720 B.n55 B.n54 163.367
R1721 B.n56 B.n55 163.367
R1722 B.n897 B.n56 163.367
R1723 B.n897 B.n61 163.367
R1724 B.n62 B.n61 163.367
R1725 B.n63 B.n62 163.367
R1726 B.n902 B.n63 163.367
R1727 B.n902 B.n68 163.367
R1728 B.n69 B.n68 163.367
R1729 B.n70 B.n69 163.367
R1730 B.n907 B.n70 163.367
R1731 B.n907 B.n75 163.367
R1732 B.n76 B.n75 163.367
R1733 B.n77 B.n76 163.367
R1734 B.n912 B.n77 163.367
R1735 B.n912 B.n82 163.367
R1736 B.n83 B.n82 163.367
R1737 B.n84 B.n83 163.367
R1738 B.n917 B.n84 163.367
R1739 B.n917 B.n89 163.367
R1740 B.n90 B.n89 163.367
R1741 B.n91 B.n90 163.367
R1742 B.n146 B.n91 163.367
R1743 B.n152 B.n95 163.367
R1744 B.n156 B.n155 163.367
R1745 B.n160 B.n159 163.367
R1746 B.n164 B.n163 163.367
R1747 B.n168 B.n167 163.367
R1748 B.n172 B.n171 163.367
R1749 B.n176 B.n175 163.367
R1750 B.n180 B.n179 163.367
R1751 B.n184 B.n183 163.367
R1752 B.n188 B.n187 163.367
R1753 B.n192 B.n191 163.367
R1754 B.n196 B.n195 163.367
R1755 B.n200 B.n199 163.367
R1756 B.n204 B.n203 163.367
R1757 B.n208 B.n207 163.367
R1758 B.n212 B.n211 163.367
R1759 B.n216 B.n215 163.367
R1760 B.n220 B.n219 163.367
R1761 B.n224 B.n223 163.367
R1762 B.n228 B.n227 163.367
R1763 B.n232 B.n231 163.367
R1764 B.n236 B.n235 163.367
R1765 B.n240 B.n239 163.367
R1766 B.n244 B.n243 163.367
R1767 B.n248 B.n247 163.367
R1768 B.n252 B.n251 163.367
R1769 B.n256 B.n255 163.367
R1770 B.n261 B.n260 163.367
R1771 B.n265 B.n264 163.367
R1772 B.n269 B.n268 163.367
R1773 B.n273 B.n272 163.367
R1774 B.n277 B.n276 163.367
R1775 B.n281 B.n280 163.367
R1776 B.n285 B.n284 163.367
R1777 B.n289 B.n288 163.367
R1778 B.n293 B.n292 163.367
R1779 B.n297 B.n296 163.367
R1780 B.n301 B.n300 163.367
R1781 B.n305 B.n304 163.367
R1782 B.n309 B.n308 163.367
R1783 B.n313 B.n312 163.367
R1784 B.n317 B.n316 163.367
R1785 B.n321 B.n320 163.367
R1786 B.n325 B.n324 163.367
R1787 B.n329 B.n328 163.367
R1788 B.n333 B.n332 163.367
R1789 B.n337 B.n336 163.367
R1790 B.n341 B.n340 163.367
R1791 B.n345 B.n344 163.367
R1792 B.n924 B.n145 163.367
R1793 B.n703 B.n702 71.676
R1794 B.n497 B.n448 71.676
R1795 B.n695 B.n449 71.676
R1796 B.n691 B.n450 71.676
R1797 B.n687 B.n451 71.676
R1798 B.n683 B.n452 71.676
R1799 B.n679 B.n453 71.676
R1800 B.n675 B.n454 71.676
R1801 B.n671 B.n455 71.676
R1802 B.n667 B.n456 71.676
R1803 B.n663 B.n457 71.676
R1804 B.n659 B.n458 71.676
R1805 B.n655 B.n459 71.676
R1806 B.n651 B.n460 71.676
R1807 B.n647 B.n461 71.676
R1808 B.n643 B.n462 71.676
R1809 B.n639 B.n463 71.676
R1810 B.n635 B.n464 71.676
R1811 B.n631 B.n465 71.676
R1812 B.n627 B.n466 71.676
R1813 B.n623 B.n467 71.676
R1814 B.n619 B.n468 71.676
R1815 B.n615 B.n469 71.676
R1816 B.n610 B.n470 71.676
R1817 B.n606 B.n471 71.676
R1818 B.n602 B.n472 71.676
R1819 B.n598 B.n473 71.676
R1820 B.n594 B.n474 71.676
R1821 B.n590 B.n475 71.676
R1822 B.n586 B.n476 71.676
R1823 B.n582 B.n477 71.676
R1824 B.n578 B.n478 71.676
R1825 B.n574 B.n479 71.676
R1826 B.n570 B.n480 71.676
R1827 B.n566 B.n481 71.676
R1828 B.n562 B.n482 71.676
R1829 B.n558 B.n483 71.676
R1830 B.n554 B.n484 71.676
R1831 B.n550 B.n485 71.676
R1832 B.n546 B.n486 71.676
R1833 B.n542 B.n487 71.676
R1834 B.n538 B.n488 71.676
R1835 B.n534 B.n489 71.676
R1836 B.n530 B.n490 71.676
R1837 B.n526 B.n491 71.676
R1838 B.n522 B.n492 71.676
R1839 B.n518 B.n493 71.676
R1840 B.n514 B.n494 71.676
R1841 B.n510 B.n495 71.676
R1842 B.n506 B.n496 71.676
R1843 B.n927 B.n926 71.676
R1844 B.n152 B.n96 71.676
R1845 B.n156 B.n97 71.676
R1846 B.n160 B.n98 71.676
R1847 B.n164 B.n99 71.676
R1848 B.n168 B.n100 71.676
R1849 B.n172 B.n101 71.676
R1850 B.n176 B.n102 71.676
R1851 B.n180 B.n103 71.676
R1852 B.n184 B.n104 71.676
R1853 B.n188 B.n105 71.676
R1854 B.n192 B.n106 71.676
R1855 B.n196 B.n107 71.676
R1856 B.n200 B.n108 71.676
R1857 B.n204 B.n109 71.676
R1858 B.n208 B.n110 71.676
R1859 B.n212 B.n111 71.676
R1860 B.n216 B.n112 71.676
R1861 B.n220 B.n113 71.676
R1862 B.n224 B.n114 71.676
R1863 B.n228 B.n115 71.676
R1864 B.n232 B.n116 71.676
R1865 B.n236 B.n117 71.676
R1866 B.n240 B.n118 71.676
R1867 B.n244 B.n119 71.676
R1868 B.n248 B.n120 71.676
R1869 B.n252 B.n121 71.676
R1870 B.n256 B.n122 71.676
R1871 B.n261 B.n123 71.676
R1872 B.n265 B.n124 71.676
R1873 B.n269 B.n125 71.676
R1874 B.n273 B.n126 71.676
R1875 B.n277 B.n127 71.676
R1876 B.n281 B.n128 71.676
R1877 B.n285 B.n129 71.676
R1878 B.n289 B.n130 71.676
R1879 B.n293 B.n131 71.676
R1880 B.n297 B.n132 71.676
R1881 B.n301 B.n133 71.676
R1882 B.n305 B.n134 71.676
R1883 B.n309 B.n135 71.676
R1884 B.n313 B.n136 71.676
R1885 B.n317 B.n137 71.676
R1886 B.n321 B.n138 71.676
R1887 B.n325 B.n139 71.676
R1888 B.n329 B.n140 71.676
R1889 B.n333 B.n141 71.676
R1890 B.n337 B.n142 71.676
R1891 B.n341 B.n143 71.676
R1892 B.n345 B.n144 71.676
R1893 B.n145 B.n144 71.676
R1894 B.n344 B.n143 71.676
R1895 B.n340 B.n142 71.676
R1896 B.n336 B.n141 71.676
R1897 B.n332 B.n140 71.676
R1898 B.n328 B.n139 71.676
R1899 B.n324 B.n138 71.676
R1900 B.n320 B.n137 71.676
R1901 B.n316 B.n136 71.676
R1902 B.n312 B.n135 71.676
R1903 B.n308 B.n134 71.676
R1904 B.n304 B.n133 71.676
R1905 B.n300 B.n132 71.676
R1906 B.n296 B.n131 71.676
R1907 B.n292 B.n130 71.676
R1908 B.n288 B.n129 71.676
R1909 B.n284 B.n128 71.676
R1910 B.n280 B.n127 71.676
R1911 B.n276 B.n126 71.676
R1912 B.n272 B.n125 71.676
R1913 B.n268 B.n124 71.676
R1914 B.n264 B.n123 71.676
R1915 B.n260 B.n122 71.676
R1916 B.n255 B.n121 71.676
R1917 B.n251 B.n120 71.676
R1918 B.n247 B.n119 71.676
R1919 B.n243 B.n118 71.676
R1920 B.n239 B.n117 71.676
R1921 B.n235 B.n116 71.676
R1922 B.n231 B.n115 71.676
R1923 B.n227 B.n114 71.676
R1924 B.n223 B.n113 71.676
R1925 B.n219 B.n112 71.676
R1926 B.n215 B.n111 71.676
R1927 B.n211 B.n110 71.676
R1928 B.n207 B.n109 71.676
R1929 B.n203 B.n108 71.676
R1930 B.n199 B.n107 71.676
R1931 B.n195 B.n106 71.676
R1932 B.n191 B.n105 71.676
R1933 B.n187 B.n104 71.676
R1934 B.n183 B.n103 71.676
R1935 B.n179 B.n102 71.676
R1936 B.n175 B.n101 71.676
R1937 B.n171 B.n100 71.676
R1938 B.n167 B.n99 71.676
R1939 B.n163 B.n98 71.676
R1940 B.n159 B.n97 71.676
R1941 B.n155 B.n96 71.676
R1942 B.n926 B.n95 71.676
R1943 B.n702 B.n447 71.676
R1944 B.n696 B.n448 71.676
R1945 B.n692 B.n449 71.676
R1946 B.n688 B.n450 71.676
R1947 B.n684 B.n451 71.676
R1948 B.n680 B.n452 71.676
R1949 B.n676 B.n453 71.676
R1950 B.n672 B.n454 71.676
R1951 B.n668 B.n455 71.676
R1952 B.n664 B.n456 71.676
R1953 B.n660 B.n457 71.676
R1954 B.n656 B.n458 71.676
R1955 B.n652 B.n459 71.676
R1956 B.n648 B.n460 71.676
R1957 B.n644 B.n461 71.676
R1958 B.n640 B.n462 71.676
R1959 B.n636 B.n463 71.676
R1960 B.n632 B.n464 71.676
R1961 B.n628 B.n465 71.676
R1962 B.n624 B.n466 71.676
R1963 B.n620 B.n467 71.676
R1964 B.n616 B.n468 71.676
R1965 B.n611 B.n469 71.676
R1966 B.n607 B.n470 71.676
R1967 B.n603 B.n471 71.676
R1968 B.n599 B.n472 71.676
R1969 B.n595 B.n473 71.676
R1970 B.n591 B.n474 71.676
R1971 B.n587 B.n475 71.676
R1972 B.n583 B.n476 71.676
R1973 B.n579 B.n477 71.676
R1974 B.n575 B.n478 71.676
R1975 B.n571 B.n479 71.676
R1976 B.n567 B.n480 71.676
R1977 B.n563 B.n481 71.676
R1978 B.n559 B.n482 71.676
R1979 B.n555 B.n483 71.676
R1980 B.n551 B.n484 71.676
R1981 B.n547 B.n485 71.676
R1982 B.n543 B.n486 71.676
R1983 B.n539 B.n487 71.676
R1984 B.n535 B.n488 71.676
R1985 B.n531 B.n489 71.676
R1986 B.n527 B.n490 71.676
R1987 B.n523 B.n491 71.676
R1988 B.n519 B.n492 71.676
R1989 B.n515 B.n493 71.676
R1990 B.n511 B.n494 71.676
R1991 B.n507 B.n495 71.676
R1992 B.n503 B.n496 71.676
R1993 B.n501 B.n500 70.5944
R1994 B.n499 B.n498 70.5944
R1995 B.n150 B.n149 70.5944
R1996 B.n148 B.n147 70.5944
R1997 B.n701 B.n444 70.2824
R1998 B.n925 B.n92 70.2824
R1999 B.n502 B.n501 59.5399
R2000 B.n613 B.n499 59.5399
R2001 B.n151 B.n150 59.5399
R2002 B.n258 B.n148 59.5399
R2003 B.n708 B.n444 40.1616
R2004 B.n708 B.n440 40.1616
R2005 B.n714 B.n440 40.1616
R2006 B.n714 B.n436 40.1616
R2007 B.n720 B.n436 40.1616
R2008 B.n720 B.n432 40.1616
R2009 B.n727 B.n432 40.1616
R2010 B.n727 B.n726 40.1616
R2011 B.n733 B.n425 40.1616
R2012 B.n739 B.n425 40.1616
R2013 B.n739 B.n421 40.1616
R2014 B.n745 B.n421 40.1616
R2015 B.n745 B.n417 40.1616
R2016 B.n751 B.n417 40.1616
R2017 B.n751 B.n413 40.1616
R2018 B.n757 B.n413 40.1616
R2019 B.n757 B.n409 40.1616
R2020 B.n763 B.n409 40.1616
R2021 B.n763 B.n404 40.1616
R2022 B.n769 B.n404 40.1616
R2023 B.n769 B.n405 40.1616
R2024 B.n775 B.n397 40.1616
R2025 B.n781 B.n397 40.1616
R2026 B.n781 B.n393 40.1616
R2027 B.n787 B.n393 40.1616
R2028 B.n787 B.n389 40.1616
R2029 B.n793 B.n389 40.1616
R2030 B.n793 B.n385 40.1616
R2031 B.n799 B.n385 40.1616
R2032 B.n799 B.n381 40.1616
R2033 B.n805 B.n381 40.1616
R2034 B.n811 B.n377 40.1616
R2035 B.n811 B.n373 40.1616
R2036 B.n817 B.n373 40.1616
R2037 B.n817 B.n369 40.1616
R2038 B.n823 B.n369 40.1616
R2039 B.n823 B.n365 40.1616
R2040 B.n829 B.n365 40.1616
R2041 B.n829 B.n361 40.1616
R2042 B.n836 B.n361 40.1616
R2043 B.n836 B.n835 40.1616
R2044 B.n842 B.n354 40.1616
R2045 B.n849 B.n354 40.1616
R2046 B.n849 B.n350 40.1616
R2047 B.n855 B.n350 40.1616
R2048 B.n855 B.n4 40.1616
R2049 B.n1030 B.n4 40.1616
R2050 B.n1030 B.n1029 40.1616
R2051 B.n1029 B.n1028 40.1616
R2052 B.n1028 B.n8 40.1616
R2053 B.n1022 B.n8 40.1616
R2054 B.n1022 B.n1021 40.1616
R2055 B.n1021 B.n1020 40.1616
R2056 B.n1014 B.n18 40.1616
R2057 B.n1014 B.n1013 40.1616
R2058 B.n1013 B.n1012 40.1616
R2059 B.n1012 B.n22 40.1616
R2060 B.n1006 B.n22 40.1616
R2061 B.n1006 B.n1005 40.1616
R2062 B.n1005 B.n1004 40.1616
R2063 B.n1004 B.n29 40.1616
R2064 B.n998 B.n29 40.1616
R2065 B.n998 B.n997 40.1616
R2066 B.n996 B.n36 40.1616
R2067 B.n990 B.n36 40.1616
R2068 B.n990 B.n989 40.1616
R2069 B.n989 B.n988 40.1616
R2070 B.n988 B.n43 40.1616
R2071 B.n982 B.n43 40.1616
R2072 B.n982 B.n981 40.1616
R2073 B.n981 B.n980 40.1616
R2074 B.n980 B.n50 40.1616
R2075 B.n974 B.n50 40.1616
R2076 B.n973 B.n972 40.1616
R2077 B.n972 B.n57 40.1616
R2078 B.n966 B.n57 40.1616
R2079 B.n966 B.n965 40.1616
R2080 B.n965 B.n964 40.1616
R2081 B.n964 B.n64 40.1616
R2082 B.n958 B.n64 40.1616
R2083 B.n958 B.n957 40.1616
R2084 B.n957 B.n956 40.1616
R2085 B.n956 B.n71 40.1616
R2086 B.n950 B.n71 40.1616
R2087 B.n950 B.n949 40.1616
R2088 B.n949 B.n948 40.1616
R2089 B.n942 B.n81 40.1616
R2090 B.n942 B.n941 40.1616
R2091 B.n941 B.n940 40.1616
R2092 B.n940 B.n85 40.1616
R2093 B.n934 B.n85 40.1616
R2094 B.n934 B.n933 40.1616
R2095 B.n933 B.n932 40.1616
R2096 B.n932 B.n92 40.1616
R2097 B.n842 B.t1 38.3898
R2098 B.n1020 B.t4 38.3898
R2099 B.n929 B.n928 30.4395
R2100 B.n923 B.n922 30.4395
R2101 B.n504 B.n442 30.4395
R2102 B.n705 B.n704 30.4395
R2103 B.n726 B.t10 28.9401
R2104 B.n81 B.t6 28.9401
R2105 B.t0 B.n377 26.5777
R2106 B.n997 B.t19 26.5777
R2107 B.n405 B.t3 25.3965
R2108 B.t2 B.n973 25.3965
R2109 B B.n1032 18.0485
R2110 B.n775 B.t3 14.7656
R2111 B.n974 B.t2 14.7656
R2112 B.n805 B.t0 13.5844
R2113 B.t19 B.n996 13.5844
R2114 B.n733 B.t10 11.222
R2115 B.n948 B.t6 11.222
R2116 B.n928 B.n94 10.6151
R2117 B.n153 B.n94 10.6151
R2118 B.n154 B.n153 10.6151
R2119 B.n157 B.n154 10.6151
R2120 B.n158 B.n157 10.6151
R2121 B.n161 B.n158 10.6151
R2122 B.n162 B.n161 10.6151
R2123 B.n165 B.n162 10.6151
R2124 B.n166 B.n165 10.6151
R2125 B.n169 B.n166 10.6151
R2126 B.n170 B.n169 10.6151
R2127 B.n173 B.n170 10.6151
R2128 B.n174 B.n173 10.6151
R2129 B.n177 B.n174 10.6151
R2130 B.n178 B.n177 10.6151
R2131 B.n181 B.n178 10.6151
R2132 B.n182 B.n181 10.6151
R2133 B.n185 B.n182 10.6151
R2134 B.n186 B.n185 10.6151
R2135 B.n189 B.n186 10.6151
R2136 B.n190 B.n189 10.6151
R2137 B.n193 B.n190 10.6151
R2138 B.n194 B.n193 10.6151
R2139 B.n197 B.n194 10.6151
R2140 B.n198 B.n197 10.6151
R2141 B.n201 B.n198 10.6151
R2142 B.n202 B.n201 10.6151
R2143 B.n205 B.n202 10.6151
R2144 B.n206 B.n205 10.6151
R2145 B.n209 B.n206 10.6151
R2146 B.n210 B.n209 10.6151
R2147 B.n213 B.n210 10.6151
R2148 B.n214 B.n213 10.6151
R2149 B.n217 B.n214 10.6151
R2150 B.n218 B.n217 10.6151
R2151 B.n221 B.n218 10.6151
R2152 B.n222 B.n221 10.6151
R2153 B.n225 B.n222 10.6151
R2154 B.n226 B.n225 10.6151
R2155 B.n229 B.n226 10.6151
R2156 B.n230 B.n229 10.6151
R2157 B.n233 B.n230 10.6151
R2158 B.n234 B.n233 10.6151
R2159 B.n237 B.n234 10.6151
R2160 B.n238 B.n237 10.6151
R2161 B.n242 B.n241 10.6151
R2162 B.n245 B.n242 10.6151
R2163 B.n246 B.n245 10.6151
R2164 B.n249 B.n246 10.6151
R2165 B.n250 B.n249 10.6151
R2166 B.n253 B.n250 10.6151
R2167 B.n254 B.n253 10.6151
R2168 B.n257 B.n254 10.6151
R2169 B.n262 B.n259 10.6151
R2170 B.n263 B.n262 10.6151
R2171 B.n266 B.n263 10.6151
R2172 B.n267 B.n266 10.6151
R2173 B.n270 B.n267 10.6151
R2174 B.n271 B.n270 10.6151
R2175 B.n274 B.n271 10.6151
R2176 B.n275 B.n274 10.6151
R2177 B.n278 B.n275 10.6151
R2178 B.n279 B.n278 10.6151
R2179 B.n282 B.n279 10.6151
R2180 B.n283 B.n282 10.6151
R2181 B.n286 B.n283 10.6151
R2182 B.n287 B.n286 10.6151
R2183 B.n290 B.n287 10.6151
R2184 B.n291 B.n290 10.6151
R2185 B.n294 B.n291 10.6151
R2186 B.n295 B.n294 10.6151
R2187 B.n298 B.n295 10.6151
R2188 B.n299 B.n298 10.6151
R2189 B.n302 B.n299 10.6151
R2190 B.n303 B.n302 10.6151
R2191 B.n306 B.n303 10.6151
R2192 B.n307 B.n306 10.6151
R2193 B.n310 B.n307 10.6151
R2194 B.n311 B.n310 10.6151
R2195 B.n314 B.n311 10.6151
R2196 B.n315 B.n314 10.6151
R2197 B.n318 B.n315 10.6151
R2198 B.n319 B.n318 10.6151
R2199 B.n322 B.n319 10.6151
R2200 B.n323 B.n322 10.6151
R2201 B.n326 B.n323 10.6151
R2202 B.n327 B.n326 10.6151
R2203 B.n330 B.n327 10.6151
R2204 B.n331 B.n330 10.6151
R2205 B.n334 B.n331 10.6151
R2206 B.n335 B.n334 10.6151
R2207 B.n338 B.n335 10.6151
R2208 B.n339 B.n338 10.6151
R2209 B.n342 B.n339 10.6151
R2210 B.n343 B.n342 10.6151
R2211 B.n346 B.n343 10.6151
R2212 B.n347 B.n346 10.6151
R2213 B.n923 B.n347 10.6151
R2214 B.n710 B.n442 10.6151
R2215 B.n711 B.n710 10.6151
R2216 B.n712 B.n711 10.6151
R2217 B.n712 B.n434 10.6151
R2218 B.n722 B.n434 10.6151
R2219 B.n723 B.n722 10.6151
R2220 B.n724 B.n723 10.6151
R2221 B.n724 B.n427 10.6151
R2222 B.n735 B.n427 10.6151
R2223 B.n736 B.n735 10.6151
R2224 B.n737 B.n736 10.6151
R2225 B.n737 B.n419 10.6151
R2226 B.n747 B.n419 10.6151
R2227 B.n748 B.n747 10.6151
R2228 B.n749 B.n748 10.6151
R2229 B.n749 B.n411 10.6151
R2230 B.n759 B.n411 10.6151
R2231 B.n760 B.n759 10.6151
R2232 B.n761 B.n760 10.6151
R2233 B.n761 B.n402 10.6151
R2234 B.n771 B.n402 10.6151
R2235 B.n772 B.n771 10.6151
R2236 B.n773 B.n772 10.6151
R2237 B.n773 B.n395 10.6151
R2238 B.n783 B.n395 10.6151
R2239 B.n784 B.n783 10.6151
R2240 B.n785 B.n784 10.6151
R2241 B.n785 B.n387 10.6151
R2242 B.n795 B.n387 10.6151
R2243 B.n796 B.n795 10.6151
R2244 B.n797 B.n796 10.6151
R2245 B.n797 B.n379 10.6151
R2246 B.n807 B.n379 10.6151
R2247 B.n808 B.n807 10.6151
R2248 B.n809 B.n808 10.6151
R2249 B.n809 B.n371 10.6151
R2250 B.n819 B.n371 10.6151
R2251 B.n820 B.n819 10.6151
R2252 B.n821 B.n820 10.6151
R2253 B.n821 B.n363 10.6151
R2254 B.n831 B.n363 10.6151
R2255 B.n832 B.n831 10.6151
R2256 B.n833 B.n832 10.6151
R2257 B.n833 B.n356 10.6151
R2258 B.n844 B.n356 10.6151
R2259 B.n845 B.n844 10.6151
R2260 B.n847 B.n845 10.6151
R2261 B.n847 B.n846 10.6151
R2262 B.n846 B.n348 10.6151
R2263 B.n858 B.n348 10.6151
R2264 B.n859 B.n858 10.6151
R2265 B.n860 B.n859 10.6151
R2266 B.n861 B.n860 10.6151
R2267 B.n863 B.n861 10.6151
R2268 B.n864 B.n863 10.6151
R2269 B.n865 B.n864 10.6151
R2270 B.n866 B.n865 10.6151
R2271 B.n868 B.n866 10.6151
R2272 B.n869 B.n868 10.6151
R2273 B.n870 B.n869 10.6151
R2274 B.n871 B.n870 10.6151
R2275 B.n873 B.n871 10.6151
R2276 B.n874 B.n873 10.6151
R2277 B.n875 B.n874 10.6151
R2278 B.n876 B.n875 10.6151
R2279 B.n878 B.n876 10.6151
R2280 B.n879 B.n878 10.6151
R2281 B.n880 B.n879 10.6151
R2282 B.n881 B.n880 10.6151
R2283 B.n883 B.n881 10.6151
R2284 B.n884 B.n883 10.6151
R2285 B.n885 B.n884 10.6151
R2286 B.n886 B.n885 10.6151
R2287 B.n888 B.n886 10.6151
R2288 B.n889 B.n888 10.6151
R2289 B.n890 B.n889 10.6151
R2290 B.n891 B.n890 10.6151
R2291 B.n893 B.n891 10.6151
R2292 B.n894 B.n893 10.6151
R2293 B.n895 B.n894 10.6151
R2294 B.n896 B.n895 10.6151
R2295 B.n898 B.n896 10.6151
R2296 B.n899 B.n898 10.6151
R2297 B.n900 B.n899 10.6151
R2298 B.n901 B.n900 10.6151
R2299 B.n903 B.n901 10.6151
R2300 B.n904 B.n903 10.6151
R2301 B.n905 B.n904 10.6151
R2302 B.n906 B.n905 10.6151
R2303 B.n908 B.n906 10.6151
R2304 B.n909 B.n908 10.6151
R2305 B.n910 B.n909 10.6151
R2306 B.n911 B.n910 10.6151
R2307 B.n913 B.n911 10.6151
R2308 B.n914 B.n913 10.6151
R2309 B.n915 B.n914 10.6151
R2310 B.n916 B.n915 10.6151
R2311 B.n918 B.n916 10.6151
R2312 B.n919 B.n918 10.6151
R2313 B.n920 B.n919 10.6151
R2314 B.n921 B.n920 10.6151
R2315 B.n922 B.n921 10.6151
R2316 B.n704 B.n446 10.6151
R2317 B.n699 B.n446 10.6151
R2318 B.n699 B.n698 10.6151
R2319 B.n698 B.n697 10.6151
R2320 B.n697 B.n694 10.6151
R2321 B.n694 B.n693 10.6151
R2322 B.n693 B.n690 10.6151
R2323 B.n690 B.n689 10.6151
R2324 B.n689 B.n686 10.6151
R2325 B.n686 B.n685 10.6151
R2326 B.n685 B.n682 10.6151
R2327 B.n682 B.n681 10.6151
R2328 B.n681 B.n678 10.6151
R2329 B.n678 B.n677 10.6151
R2330 B.n677 B.n674 10.6151
R2331 B.n674 B.n673 10.6151
R2332 B.n673 B.n670 10.6151
R2333 B.n670 B.n669 10.6151
R2334 B.n669 B.n666 10.6151
R2335 B.n666 B.n665 10.6151
R2336 B.n665 B.n662 10.6151
R2337 B.n662 B.n661 10.6151
R2338 B.n661 B.n658 10.6151
R2339 B.n658 B.n657 10.6151
R2340 B.n657 B.n654 10.6151
R2341 B.n654 B.n653 10.6151
R2342 B.n653 B.n650 10.6151
R2343 B.n650 B.n649 10.6151
R2344 B.n649 B.n646 10.6151
R2345 B.n646 B.n645 10.6151
R2346 B.n645 B.n642 10.6151
R2347 B.n642 B.n641 10.6151
R2348 B.n641 B.n638 10.6151
R2349 B.n638 B.n637 10.6151
R2350 B.n637 B.n634 10.6151
R2351 B.n634 B.n633 10.6151
R2352 B.n633 B.n630 10.6151
R2353 B.n630 B.n629 10.6151
R2354 B.n629 B.n626 10.6151
R2355 B.n626 B.n625 10.6151
R2356 B.n625 B.n622 10.6151
R2357 B.n622 B.n621 10.6151
R2358 B.n621 B.n618 10.6151
R2359 B.n618 B.n617 10.6151
R2360 B.n617 B.n614 10.6151
R2361 B.n612 B.n609 10.6151
R2362 B.n609 B.n608 10.6151
R2363 B.n608 B.n605 10.6151
R2364 B.n605 B.n604 10.6151
R2365 B.n604 B.n601 10.6151
R2366 B.n601 B.n600 10.6151
R2367 B.n600 B.n597 10.6151
R2368 B.n597 B.n596 10.6151
R2369 B.n593 B.n592 10.6151
R2370 B.n592 B.n589 10.6151
R2371 B.n589 B.n588 10.6151
R2372 B.n588 B.n585 10.6151
R2373 B.n585 B.n584 10.6151
R2374 B.n584 B.n581 10.6151
R2375 B.n581 B.n580 10.6151
R2376 B.n580 B.n577 10.6151
R2377 B.n577 B.n576 10.6151
R2378 B.n576 B.n573 10.6151
R2379 B.n573 B.n572 10.6151
R2380 B.n572 B.n569 10.6151
R2381 B.n569 B.n568 10.6151
R2382 B.n568 B.n565 10.6151
R2383 B.n565 B.n564 10.6151
R2384 B.n564 B.n561 10.6151
R2385 B.n561 B.n560 10.6151
R2386 B.n560 B.n557 10.6151
R2387 B.n557 B.n556 10.6151
R2388 B.n556 B.n553 10.6151
R2389 B.n553 B.n552 10.6151
R2390 B.n552 B.n549 10.6151
R2391 B.n549 B.n548 10.6151
R2392 B.n548 B.n545 10.6151
R2393 B.n545 B.n544 10.6151
R2394 B.n544 B.n541 10.6151
R2395 B.n541 B.n540 10.6151
R2396 B.n540 B.n537 10.6151
R2397 B.n537 B.n536 10.6151
R2398 B.n536 B.n533 10.6151
R2399 B.n533 B.n532 10.6151
R2400 B.n532 B.n529 10.6151
R2401 B.n529 B.n528 10.6151
R2402 B.n528 B.n525 10.6151
R2403 B.n525 B.n524 10.6151
R2404 B.n524 B.n521 10.6151
R2405 B.n521 B.n520 10.6151
R2406 B.n520 B.n517 10.6151
R2407 B.n517 B.n516 10.6151
R2408 B.n516 B.n513 10.6151
R2409 B.n513 B.n512 10.6151
R2410 B.n512 B.n509 10.6151
R2411 B.n509 B.n508 10.6151
R2412 B.n508 B.n505 10.6151
R2413 B.n505 B.n504 10.6151
R2414 B.n706 B.n705 10.6151
R2415 B.n706 B.n438 10.6151
R2416 B.n716 B.n438 10.6151
R2417 B.n717 B.n716 10.6151
R2418 B.n718 B.n717 10.6151
R2419 B.n718 B.n430 10.6151
R2420 B.n729 B.n430 10.6151
R2421 B.n730 B.n729 10.6151
R2422 B.n731 B.n730 10.6151
R2423 B.n731 B.n423 10.6151
R2424 B.n741 B.n423 10.6151
R2425 B.n742 B.n741 10.6151
R2426 B.n743 B.n742 10.6151
R2427 B.n743 B.n415 10.6151
R2428 B.n753 B.n415 10.6151
R2429 B.n754 B.n753 10.6151
R2430 B.n755 B.n754 10.6151
R2431 B.n755 B.n407 10.6151
R2432 B.n765 B.n407 10.6151
R2433 B.n766 B.n765 10.6151
R2434 B.n767 B.n766 10.6151
R2435 B.n767 B.n399 10.6151
R2436 B.n777 B.n399 10.6151
R2437 B.n778 B.n777 10.6151
R2438 B.n779 B.n778 10.6151
R2439 B.n779 B.n391 10.6151
R2440 B.n789 B.n391 10.6151
R2441 B.n790 B.n789 10.6151
R2442 B.n791 B.n790 10.6151
R2443 B.n791 B.n383 10.6151
R2444 B.n801 B.n383 10.6151
R2445 B.n802 B.n801 10.6151
R2446 B.n803 B.n802 10.6151
R2447 B.n803 B.n375 10.6151
R2448 B.n813 B.n375 10.6151
R2449 B.n814 B.n813 10.6151
R2450 B.n815 B.n814 10.6151
R2451 B.n815 B.n367 10.6151
R2452 B.n825 B.n367 10.6151
R2453 B.n826 B.n825 10.6151
R2454 B.n827 B.n826 10.6151
R2455 B.n827 B.n359 10.6151
R2456 B.n838 B.n359 10.6151
R2457 B.n839 B.n838 10.6151
R2458 B.n840 B.n839 10.6151
R2459 B.n840 B.n352 10.6151
R2460 B.n851 B.n352 10.6151
R2461 B.n852 B.n851 10.6151
R2462 B.n853 B.n852 10.6151
R2463 B.n853 B.n0 10.6151
R2464 B.n1026 B.n1 10.6151
R2465 B.n1026 B.n1025 10.6151
R2466 B.n1025 B.n1024 10.6151
R2467 B.n1024 B.n10 10.6151
R2468 B.n1018 B.n10 10.6151
R2469 B.n1018 B.n1017 10.6151
R2470 B.n1017 B.n1016 10.6151
R2471 B.n1016 B.n16 10.6151
R2472 B.n1010 B.n16 10.6151
R2473 B.n1010 B.n1009 10.6151
R2474 B.n1009 B.n1008 10.6151
R2475 B.n1008 B.n24 10.6151
R2476 B.n1002 B.n24 10.6151
R2477 B.n1002 B.n1001 10.6151
R2478 B.n1001 B.n1000 10.6151
R2479 B.n1000 B.n31 10.6151
R2480 B.n994 B.n31 10.6151
R2481 B.n994 B.n993 10.6151
R2482 B.n993 B.n992 10.6151
R2483 B.n992 B.n38 10.6151
R2484 B.n986 B.n38 10.6151
R2485 B.n986 B.n985 10.6151
R2486 B.n985 B.n984 10.6151
R2487 B.n984 B.n45 10.6151
R2488 B.n978 B.n45 10.6151
R2489 B.n978 B.n977 10.6151
R2490 B.n977 B.n976 10.6151
R2491 B.n976 B.n52 10.6151
R2492 B.n970 B.n52 10.6151
R2493 B.n970 B.n969 10.6151
R2494 B.n969 B.n968 10.6151
R2495 B.n968 B.n59 10.6151
R2496 B.n962 B.n59 10.6151
R2497 B.n962 B.n961 10.6151
R2498 B.n961 B.n960 10.6151
R2499 B.n960 B.n66 10.6151
R2500 B.n954 B.n66 10.6151
R2501 B.n954 B.n953 10.6151
R2502 B.n953 B.n952 10.6151
R2503 B.n952 B.n73 10.6151
R2504 B.n946 B.n73 10.6151
R2505 B.n946 B.n945 10.6151
R2506 B.n945 B.n944 10.6151
R2507 B.n944 B.n79 10.6151
R2508 B.n938 B.n79 10.6151
R2509 B.n938 B.n937 10.6151
R2510 B.n937 B.n936 10.6151
R2511 B.n936 B.n87 10.6151
R2512 B.n930 B.n87 10.6151
R2513 B.n930 B.n929 10.6151
R2514 B.n241 B.n151 6.5566
R2515 B.n258 B.n257 6.5566
R2516 B.n613 B.n612 6.5566
R2517 B.n596 B.n502 6.5566
R2518 B.n238 B.n151 4.05904
R2519 B.n259 B.n258 4.05904
R2520 B.n614 B.n613 4.05904
R2521 B.n593 B.n502 4.05904
R2522 B.n1032 B.n0 2.81026
R2523 B.n1032 B.n1 2.81026
R2524 B.n835 B.t1 1.77231
R2525 B.n18 B.t4 1.77231
R2526 VN.n34 VN.n33 161.3
R2527 VN.n32 VN.n19 161.3
R2528 VN.n31 VN.n30 161.3
R2529 VN.n29 VN.n20 161.3
R2530 VN.n28 VN.n27 161.3
R2531 VN.n26 VN.n21 161.3
R2532 VN.n25 VN.n24 161.3
R2533 VN.n16 VN.n15 161.3
R2534 VN.n14 VN.n1 161.3
R2535 VN.n13 VN.n12 161.3
R2536 VN.n11 VN.n2 161.3
R2537 VN.n10 VN.n9 161.3
R2538 VN.n8 VN.n3 161.3
R2539 VN.n7 VN.n6 161.3
R2540 VN.n23 VN.t4 130.5
R2541 VN.n5 VN.t5 130.5
R2542 VN.n4 VN.t0 97.2014
R2543 VN.n0 VN.t3 97.2014
R2544 VN.n22 VN.t2 97.2014
R2545 VN.n18 VN.t1 97.2014
R2546 VN.n17 VN.n0 70.9831
R2547 VN.n35 VN.n18 70.9831
R2548 VN.n5 VN.n4 62.0573
R2549 VN.n23 VN.n22 62.0573
R2550 VN VN.n35 52.8314
R2551 VN.n13 VN.n2 47.2923
R2552 VN.n31 VN.n20 47.2923
R2553 VN.n9 VN.n2 33.6945
R2554 VN.n27 VN.n20 33.6945
R2555 VN.n8 VN.n7 24.4675
R2556 VN.n9 VN.n8 24.4675
R2557 VN.n14 VN.n13 24.4675
R2558 VN.n15 VN.n14 24.4675
R2559 VN.n27 VN.n26 24.4675
R2560 VN.n26 VN.n25 24.4675
R2561 VN.n33 VN.n32 24.4675
R2562 VN.n32 VN.n31 24.4675
R2563 VN.n15 VN.n0 19.0848
R2564 VN.n33 VN.n18 19.0848
R2565 VN.n7 VN.n4 12.234
R2566 VN.n25 VN.n22 12.234
R2567 VN.n24 VN.n23 3.94734
R2568 VN.n6 VN.n5 3.94734
R2569 VN.n35 VN.n34 0.354971
R2570 VN.n17 VN.n16 0.354971
R2571 VN VN.n17 0.26696
R2572 VN.n34 VN.n19 0.189894
R2573 VN.n30 VN.n19 0.189894
R2574 VN.n30 VN.n29 0.189894
R2575 VN.n29 VN.n28 0.189894
R2576 VN.n28 VN.n21 0.189894
R2577 VN.n24 VN.n21 0.189894
R2578 VN.n6 VN.n3 0.189894
R2579 VN.n10 VN.n3 0.189894
R2580 VN.n11 VN.n10 0.189894
R2581 VN.n12 VN.n11 0.189894
R2582 VN.n12 VN.n1 0.189894
R2583 VN.n16 VN.n1 0.189894
R2584 VDD2.n139 VDD2.n73 214.453
R2585 VDD2.n66 VDD2.n0 214.453
R2586 VDD2.n140 VDD2.n139 185
R2587 VDD2.n138 VDD2.n137 185
R2588 VDD2.n77 VDD2.n76 185
R2589 VDD2.n132 VDD2.n131 185
R2590 VDD2.n130 VDD2.n129 185
R2591 VDD2.n81 VDD2.n80 185
R2592 VDD2.n124 VDD2.n123 185
R2593 VDD2.n122 VDD2.n121 185
R2594 VDD2.n85 VDD2.n84 185
R2595 VDD2.n116 VDD2.n115 185
R2596 VDD2.n114 VDD2.n113 185
R2597 VDD2.n89 VDD2.n88 185
R2598 VDD2.n108 VDD2.n107 185
R2599 VDD2.n106 VDD2.n105 185
R2600 VDD2.n93 VDD2.n92 185
R2601 VDD2.n100 VDD2.n99 185
R2602 VDD2.n98 VDD2.n97 185
R2603 VDD2.n25 VDD2.n24 185
R2604 VDD2.n27 VDD2.n26 185
R2605 VDD2.n20 VDD2.n19 185
R2606 VDD2.n33 VDD2.n32 185
R2607 VDD2.n35 VDD2.n34 185
R2608 VDD2.n16 VDD2.n15 185
R2609 VDD2.n41 VDD2.n40 185
R2610 VDD2.n43 VDD2.n42 185
R2611 VDD2.n12 VDD2.n11 185
R2612 VDD2.n49 VDD2.n48 185
R2613 VDD2.n51 VDD2.n50 185
R2614 VDD2.n8 VDD2.n7 185
R2615 VDD2.n57 VDD2.n56 185
R2616 VDD2.n59 VDD2.n58 185
R2617 VDD2.n4 VDD2.n3 185
R2618 VDD2.n65 VDD2.n64 185
R2619 VDD2.n67 VDD2.n66 185
R2620 VDD2.n23 VDD2.t0 147.659
R2621 VDD2.n96 VDD2.t4 147.659
R2622 VDD2.n139 VDD2.n138 104.615
R2623 VDD2.n138 VDD2.n76 104.615
R2624 VDD2.n131 VDD2.n76 104.615
R2625 VDD2.n131 VDD2.n130 104.615
R2626 VDD2.n130 VDD2.n80 104.615
R2627 VDD2.n123 VDD2.n80 104.615
R2628 VDD2.n123 VDD2.n122 104.615
R2629 VDD2.n122 VDD2.n84 104.615
R2630 VDD2.n115 VDD2.n84 104.615
R2631 VDD2.n115 VDD2.n114 104.615
R2632 VDD2.n114 VDD2.n88 104.615
R2633 VDD2.n107 VDD2.n88 104.615
R2634 VDD2.n107 VDD2.n106 104.615
R2635 VDD2.n106 VDD2.n92 104.615
R2636 VDD2.n99 VDD2.n92 104.615
R2637 VDD2.n99 VDD2.n98 104.615
R2638 VDD2.n26 VDD2.n25 104.615
R2639 VDD2.n26 VDD2.n19 104.615
R2640 VDD2.n33 VDD2.n19 104.615
R2641 VDD2.n34 VDD2.n33 104.615
R2642 VDD2.n34 VDD2.n15 104.615
R2643 VDD2.n41 VDD2.n15 104.615
R2644 VDD2.n42 VDD2.n41 104.615
R2645 VDD2.n42 VDD2.n11 104.615
R2646 VDD2.n49 VDD2.n11 104.615
R2647 VDD2.n50 VDD2.n49 104.615
R2648 VDD2.n50 VDD2.n7 104.615
R2649 VDD2.n57 VDD2.n7 104.615
R2650 VDD2.n58 VDD2.n57 104.615
R2651 VDD2.n58 VDD2.n3 104.615
R2652 VDD2.n65 VDD2.n3 104.615
R2653 VDD2.n66 VDD2.n65 104.615
R2654 VDD2.n72 VDD2.n71 64.7577
R2655 VDD2 VDD2.n145 64.7548
R2656 VDD2.n72 VDD2.n70 54.0713
R2657 VDD2.n98 VDD2.t4 52.3082
R2658 VDD2.n25 VDD2.t0 52.3082
R2659 VDD2.n144 VDD2.n143 51.7732
R2660 VDD2.n144 VDD2.n72 45.4222
R2661 VDD2.n97 VDD2.n96 15.6677
R2662 VDD2.n24 VDD2.n23 15.6677
R2663 VDD2.n141 VDD2.n140 12.8005
R2664 VDD2.n100 VDD2.n95 12.8005
R2665 VDD2.n27 VDD2.n22 12.8005
R2666 VDD2.n68 VDD2.n67 12.8005
R2667 VDD2.n137 VDD2.n75 12.0247
R2668 VDD2.n101 VDD2.n93 12.0247
R2669 VDD2.n28 VDD2.n20 12.0247
R2670 VDD2.n64 VDD2.n2 12.0247
R2671 VDD2.n136 VDD2.n77 11.249
R2672 VDD2.n105 VDD2.n104 11.249
R2673 VDD2.n32 VDD2.n31 11.249
R2674 VDD2.n63 VDD2.n4 11.249
R2675 VDD2.n133 VDD2.n132 10.4732
R2676 VDD2.n108 VDD2.n91 10.4732
R2677 VDD2.n35 VDD2.n18 10.4732
R2678 VDD2.n60 VDD2.n59 10.4732
R2679 VDD2.n129 VDD2.n79 9.69747
R2680 VDD2.n109 VDD2.n89 9.69747
R2681 VDD2.n36 VDD2.n16 9.69747
R2682 VDD2.n56 VDD2.n6 9.69747
R2683 VDD2.n143 VDD2.n142 9.45567
R2684 VDD2.n70 VDD2.n69 9.45567
R2685 VDD2.n83 VDD2.n82 9.3005
R2686 VDD2.n126 VDD2.n125 9.3005
R2687 VDD2.n128 VDD2.n127 9.3005
R2688 VDD2.n79 VDD2.n78 9.3005
R2689 VDD2.n134 VDD2.n133 9.3005
R2690 VDD2.n136 VDD2.n135 9.3005
R2691 VDD2.n75 VDD2.n74 9.3005
R2692 VDD2.n142 VDD2.n141 9.3005
R2693 VDD2.n120 VDD2.n119 9.3005
R2694 VDD2.n118 VDD2.n117 9.3005
R2695 VDD2.n87 VDD2.n86 9.3005
R2696 VDD2.n112 VDD2.n111 9.3005
R2697 VDD2.n110 VDD2.n109 9.3005
R2698 VDD2.n91 VDD2.n90 9.3005
R2699 VDD2.n104 VDD2.n103 9.3005
R2700 VDD2.n102 VDD2.n101 9.3005
R2701 VDD2.n95 VDD2.n94 9.3005
R2702 VDD2.n45 VDD2.n44 9.3005
R2703 VDD2.n14 VDD2.n13 9.3005
R2704 VDD2.n39 VDD2.n38 9.3005
R2705 VDD2.n37 VDD2.n36 9.3005
R2706 VDD2.n18 VDD2.n17 9.3005
R2707 VDD2.n31 VDD2.n30 9.3005
R2708 VDD2.n29 VDD2.n28 9.3005
R2709 VDD2.n22 VDD2.n21 9.3005
R2710 VDD2.n47 VDD2.n46 9.3005
R2711 VDD2.n10 VDD2.n9 9.3005
R2712 VDD2.n53 VDD2.n52 9.3005
R2713 VDD2.n55 VDD2.n54 9.3005
R2714 VDD2.n6 VDD2.n5 9.3005
R2715 VDD2.n61 VDD2.n60 9.3005
R2716 VDD2.n63 VDD2.n62 9.3005
R2717 VDD2.n2 VDD2.n1 9.3005
R2718 VDD2.n69 VDD2.n68 9.3005
R2719 VDD2.n128 VDD2.n81 8.92171
R2720 VDD2.n113 VDD2.n112 8.92171
R2721 VDD2.n40 VDD2.n39 8.92171
R2722 VDD2.n55 VDD2.n8 8.92171
R2723 VDD2.n143 VDD2.n73 8.2187
R2724 VDD2.n70 VDD2.n0 8.2187
R2725 VDD2.n125 VDD2.n124 8.14595
R2726 VDD2.n116 VDD2.n87 8.14595
R2727 VDD2.n43 VDD2.n14 8.14595
R2728 VDD2.n52 VDD2.n51 8.14595
R2729 VDD2.n121 VDD2.n83 7.3702
R2730 VDD2.n117 VDD2.n85 7.3702
R2731 VDD2.n44 VDD2.n12 7.3702
R2732 VDD2.n48 VDD2.n10 7.3702
R2733 VDD2.n121 VDD2.n120 6.59444
R2734 VDD2.n120 VDD2.n85 6.59444
R2735 VDD2.n47 VDD2.n12 6.59444
R2736 VDD2.n48 VDD2.n47 6.59444
R2737 VDD2.n124 VDD2.n83 5.81868
R2738 VDD2.n117 VDD2.n116 5.81868
R2739 VDD2.n44 VDD2.n43 5.81868
R2740 VDD2.n51 VDD2.n10 5.81868
R2741 VDD2.n141 VDD2.n73 5.3904
R2742 VDD2.n68 VDD2.n0 5.3904
R2743 VDD2.n125 VDD2.n81 5.04292
R2744 VDD2.n113 VDD2.n87 5.04292
R2745 VDD2.n40 VDD2.n14 5.04292
R2746 VDD2.n52 VDD2.n8 5.04292
R2747 VDD2.n23 VDD2.n21 4.38563
R2748 VDD2.n96 VDD2.n94 4.38563
R2749 VDD2.n129 VDD2.n128 4.26717
R2750 VDD2.n112 VDD2.n89 4.26717
R2751 VDD2.n39 VDD2.n16 4.26717
R2752 VDD2.n56 VDD2.n55 4.26717
R2753 VDD2.n132 VDD2.n79 3.49141
R2754 VDD2.n109 VDD2.n108 3.49141
R2755 VDD2.n36 VDD2.n35 3.49141
R2756 VDD2.n59 VDD2.n6 3.49141
R2757 VDD2.n133 VDD2.n77 2.71565
R2758 VDD2.n105 VDD2.n91 2.71565
R2759 VDD2.n32 VDD2.n18 2.71565
R2760 VDD2.n60 VDD2.n4 2.71565
R2761 VDD2 VDD2.n144 2.41214
R2762 VDD2.n137 VDD2.n136 1.93989
R2763 VDD2.n104 VDD2.n93 1.93989
R2764 VDD2.n31 VDD2.n20 1.93989
R2765 VDD2.n64 VDD2.n63 1.93989
R2766 VDD2.n145 VDD2.t3 1.48365
R2767 VDD2.n145 VDD2.t1 1.48365
R2768 VDD2.n71 VDD2.t5 1.48365
R2769 VDD2.n71 VDD2.t2 1.48365
R2770 VDD2.n140 VDD2.n75 1.16414
R2771 VDD2.n101 VDD2.n100 1.16414
R2772 VDD2.n28 VDD2.n27 1.16414
R2773 VDD2.n67 VDD2.n2 1.16414
R2774 VDD2.n97 VDD2.n95 0.388379
R2775 VDD2.n24 VDD2.n22 0.388379
R2776 VDD2.n142 VDD2.n74 0.155672
R2777 VDD2.n135 VDD2.n74 0.155672
R2778 VDD2.n135 VDD2.n134 0.155672
R2779 VDD2.n134 VDD2.n78 0.155672
R2780 VDD2.n127 VDD2.n78 0.155672
R2781 VDD2.n127 VDD2.n126 0.155672
R2782 VDD2.n126 VDD2.n82 0.155672
R2783 VDD2.n119 VDD2.n82 0.155672
R2784 VDD2.n119 VDD2.n118 0.155672
R2785 VDD2.n118 VDD2.n86 0.155672
R2786 VDD2.n111 VDD2.n86 0.155672
R2787 VDD2.n111 VDD2.n110 0.155672
R2788 VDD2.n110 VDD2.n90 0.155672
R2789 VDD2.n103 VDD2.n90 0.155672
R2790 VDD2.n103 VDD2.n102 0.155672
R2791 VDD2.n102 VDD2.n94 0.155672
R2792 VDD2.n29 VDD2.n21 0.155672
R2793 VDD2.n30 VDD2.n29 0.155672
R2794 VDD2.n30 VDD2.n17 0.155672
R2795 VDD2.n37 VDD2.n17 0.155672
R2796 VDD2.n38 VDD2.n37 0.155672
R2797 VDD2.n38 VDD2.n13 0.155672
R2798 VDD2.n45 VDD2.n13 0.155672
R2799 VDD2.n46 VDD2.n45 0.155672
R2800 VDD2.n46 VDD2.n9 0.155672
R2801 VDD2.n53 VDD2.n9 0.155672
R2802 VDD2.n54 VDD2.n53 0.155672
R2803 VDD2.n54 VDD2.n5 0.155672
R2804 VDD2.n61 VDD2.n5 0.155672
R2805 VDD2.n62 VDD2.n61 0.155672
R2806 VDD2.n62 VDD2.n1 0.155672
R2807 VDD2.n69 VDD2.n1 0.155672
C0 VDD1 VN 0.151625f
C1 VP VDD2 0.518527f
C2 VDD1 VTAIL 8.39009f
C3 VDD2 VN 7.75287f
C4 VDD2 VTAIL 8.44608f
C5 VP VN 7.86456f
C6 VDD1 VDD2 1.68346f
C7 VP VTAIL 8.034241f
C8 VN VTAIL 8.019979f
C9 VP VDD1 8.1165f
C10 VDD2 B 6.759055f
C11 VDD1 B 6.928947f
C12 VTAIL B 8.819215f
C13 VN B 15.07806f
C14 VP B 13.754593f
C15 VDD2.n0 B 0.029103f
C16 VDD2.n1 B 0.021291f
C17 VDD2.n2 B 0.011441f
C18 VDD2.n3 B 0.027042f
C19 VDD2.n4 B 0.012114f
C20 VDD2.n5 B 0.021291f
C21 VDD2.n6 B 0.011441f
C22 VDD2.n7 B 0.027042f
C23 VDD2.n8 B 0.012114f
C24 VDD2.n9 B 0.021291f
C25 VDD2.n10 B 0.011441f
C26 VDD2.n11 B 0.027042f
C27 VDD2.n12 B 0.012114f
C28 VDD2.n13 B 0.021291f
C29 VDD2.n14 B 0.011441f
C30 VDD2.n15 B 0.027042f
C31 VDD2.n16 B 0.012114f
C32 VDD2.n17 B 0.021291f
C33 VDD2.n18 B 0.011441f
C34 VDD2.n19 B 0.027042f
C35 VDD2.n20 B 0.012114f
C36 VDD2.n21 B 1.22423f
C37 VDD2.n22 B 0.011441f
C38 VDD2.t0 B 0.044469f
C39 VDD2.n23 B 0.130058f
C40 VDD2.n24 B 0.015975f
C41 VDD2.n25 B 0.020282f
C42 VDD2.n26 B 0.027042f
C43 VDD2.n27 B 0.012114f
C44 VDD2.n28 B 0.011441f
C45 VDD2.n29 B 0.021291f
C46 VDD2.n30 B 0.021291f
C47 VDD2.n31 B 0.011441f
C48 VDD2.n32 B 0.012114f
C49 VDD2.n33 B 0.027042f
C50 VDD2.n34 B 0.027042f
C51 VDD2.n35 B 0.012114f
C52 VDD2.n36 B 0.011441f
C53 VDD2.n37 B 0.021291f
C54 VDD2.n38 B 0.021291f
C55 VDD2.n39 B 0.011441f
C56 VDD2.n40 B 0.012114f
C57 VDD2.n41 B 0.027042f
C58 VDD2.n42 B 0.027042f
C59 VDD2.n43 B 0.012114f
C60 VDD2.n44 B 0.011441f
C61 VDD2.n45 B 0.021291f
C62 VDD2.n46 B 0.021291f
C63 VDD2.n47 B 0.011441f
C64 VDD2.n48 B 0.012114f
C65 VDD2.n49 B 0.027042f
C66 VDD2.n50 B 0.027042f
C67 VDD2.n51 B 0.012114f
C68 VDD2.n52 B 0.011441f
C69 VDD2.n53 B 0.021291f
C70 VDD2.n54 B 0.021291f
C71 VDD2.n55 B 0.011441f
C72 VDD2.n56 B 0.012114f
C73 VDD2.n57 B 0.027042f
C74 VDD2.n58 B 0.027042f
C75 VDD2.n59 B 0.012114f
C76 VDD2.n60 B 0.011441f
C77 VDD2.n61 B 0.021291f
C78 VDD2.n62 B 0.021291f
C79 VDD2.n63 B 0.011441f
C80 VDD2.n64 B 0.012114f
C81 VDD2.n65 B 0.027042f
C82 VDD2.n66 B 0.055335f
C83 VDD2.n67 B 0.012114f
C84 VDD2.n68 B 0.022371f
C85 VDD2.n69 B 0.053577f
C86 VDD2.n70 B 0.080341f
C87 VDD2.t5 B 0.224613f
C88 VDD2.t2 B 0.224613f
C89 VDD2.n71 B 2.02635f
C90 VDD2.n72 B 2.61079f
C91 VDD2.n73 B 0.029103f
C92 VDD2.n74 B 0.021291f
C93 VDD2.n75 B 0.011441f
C94 VDD2.n76 B 0.027042f
C95 VDD2.n77 B 0.012114f
C96 VDD2.n78 B 0.021291f
C97 VDD2.n79 B 0.011441f
C98 VDD2.n80 B 0.027042f
C99 VDD2.n81 B 0.012114f
C100 VDD2.n82 B 0.021291f
C101 VDD2.n83 B 0.011441f
C102 VDD2.n84 B 0.027042f
C103 VDD2.n85 B 0.012114f
C104 VDD2.n86 B 0.021291f
C105 VDD2.n87 B 0.011441f
C106 VDD2.n88 B 0.027042f
C107 VDD2.n89 B 0.012114f
C108 VDD2.n90 B 0.021291f
C109 VDD2.n91 B 0.011441f
C110 VDD2.n92 B 0.027042f
C111 VDD2.n93 B 0.012114f
C112 VDD2.n94 B 1.22423f
C113 VDD2.n95 B 0.011441f
C114 VDD2.t4 B 0.044469f
C115 VDD2.n96 B 0.130058f
C116 VDD2.n97 B 0.015975f
C117 VDD2.n98 B 0.020282f
C118 VDD2.n99 B 0.027042f
C119 VDD2.n100 B 0.012114f
C120 VDD2.n101 B 0.011441f
C121 VDD2.n102 B 0.021291f
C122 VDD2.n103 B 0.021291f
C123 VDD2.n104 B 0.011441f
C124 VDD2.n105 B 0.012114f
C125 VDD2.n106 B 0.027042f
C126 VDD2.n107 B 0.027042f
C127 VDD2.n108 B 0.012114f
C128 VDD2.n109 B 0.011441f
C129 VDD2.n110 B 0.021291f
C130 VDD2.n111 B 0.021291f
C131 VDD2.n112 B 0.011441f
C132 VDD2.n113 B 0.012114f
C133 VDD2.n114 B 0.027042f
C134 VDD2.n115 B 0.027042f
C135 VDD2.n116 B 0.012114f
C136 VDD2.n117 B 0.011441f
C137 VDD2.n118 B 0.021291f
C138 VDD2.n119 B 0.021291f
C139 VDD2.n120 B 0.011441f
C140 VDD2.n121 B 0.012114f
C141 VDD2.n122 B 0.027042f
C142 VDD2.n123 B 0.027042f
C143 VDD2.n124 B 0.012114f
C144 VDD2.n125 B 0.011441f
C145 VDD2.n126 B 0.021291f
C146 VDD2.n127 B 0.021291f
C147 VDD2.n128 B 0.011441f
C148 VDD2.n129 B 0.012114f
C149 VDD2.n130 B 0.027042f
C150 VDD2.n131 B 0.027042f
C151 VDD2.n132 B 0.012114f
C152 VDD2.n133 B 0.011441f
C153 VDD2.n134 B 0.021291f
C154 VDD2.n135 B 0.021291f
C155 VDD2.n136 B 0.011441f
C156 VDD2.n137 B 0.012114f
C157 VDD2.n138 B 0.027042f
C158 VDD2.n139 B 0.055335f
C159 VDD2.n140 B 0.012114f
C160 VDD2.n141 B 0.022371f
C161 VDD2.n142 B 0.053577f
C162 VDD2.n143 B 0.071782f
C163 VDD2.n144 B 2.43736f
C164 VDD2.t3 B 0.224613f
C165 VDD2.t1 B 0.224613f
C166 VDD2.n145 B 2.02632f
C167 VN.t3 B 2.37547f
C168 VN.n0 B 0.913718f
C169 VN.n1 B 0.019674f
C170 VN.n2 B 0.017178f
C171 VN.n3 B 0.019674f
C172 VN.t0 B 2.37547f
C173 VN.n4 B 0.895904f
C174 VN.t5 B 2.62427f
C175 VN.n5 B 0.854726f
C176 VN.n6 B 0.229527f
C177 VN.n7 B 0.027615f
C178 VN.n8 B 0.036667f
C179 VN.n9 B 0.039739f
C180 VN.n10 B 0.019674f
C181 VN.n11 B 0.019674f
C182 VN.n12 B 0.019674f
C183 VN.n13 B 0.037189f
C184 VN.n14 B 0.036667f
C185 VN.n15 B 0.032684f
C186 VN.n16 B 0.031753f
C187 VN.n17 B 0.04384f
C188 VN.t1 B 2.37547f
C189 VN.n18 B 0.913718f
C190 VN.n19 B 0.019674f
C191 VN.n20 B 0.017178f
C192 VN.n21 B 0.019674f
C193 VN.t2 B 2.37547f
C194 VN.n22 B 0.895904f
C195 VN.t4 B 2.62427f
C196 VN.n23 B 0.854726f
C197 VN.n24 B 0.229527f
C198 VN.n25 B 0.027615f
C199 VN.n26 B 0.036667f
C200 VN.n27 B 0.039739f
C201 VN.n28 B 0.019674f
C202 VN.n29 B 0.019674f
C203 VN.n30 B 0.019674f
C204 VN.n31 B 0.037189f
C205 VN.n32 B 0.036667f
C206 VN.n33 B 0.032684f
C207 VN.n34 B 0.031753f
C208 VN.n35 B 1.21042f
C209 VDD1.n0 B 0.029499f
C210 VDD1.n1 B 0.021581f
C211 VDD1.n2 B 0.011597f
C212 VDD1.n3 B 0.02741f
C213 VDD1.n4 B 0.012279f
C214 VDD1.n5 B 0.021581f
C215 VDD1.n6 B 0.011597f
C216 VDD1.n7 B 0.02741f
C217 VDD1.n8 B 0.012279f
C218 VDD1.n9 B 0.021581f
C219 VDD1.n10 B 0.011597f
C220 VDD1.n11 B 0.02741f
C221 VDD1.n12 B 0.012279f
C222 VDD1.n13 B 0.021581f
C223 VDD1.n14 B 0.011597f
C224 VDD1.n15 B 0.02741f
C225 VDD1.n16 B 0.012279f
C226 VDD1.n17 B 0.021581f
C227 VDD1.n18 B 0.011597f
C228 VDD1.n19 B 0.02741f
C229 VDD1.n20 B 0.012279f
C230 VDD1.n21 B 1.24088f
C231 VDD1.n22 B 0.011597f
C232 VDD1.t1 B 0.045074f
C233 VDD1.n23 B 0.131826f
C234 VDD1.n24 B 0.016192f
C235 VDD1.n25 B 0.020558f
C236 VDD1.n26 B 0.02741f
C237 VDD1.n27 B 0.012279f
C238 VDD1.n28 B 0.011597f
C239 VDD1.n29 B 0.021581f
C240 VDD1.n30 B 0.021581f
C241 VDD1.n31 B 0.011597f
C242 VDD1.n32 B 0.012279f
C243 VDD1.n33 B 0.02741f
C244 VDD1.n34 B 0.02741f
C245 VDD1.n35 B 0.012279f
C246 VDD1.n36 B 0.011597f
C247 VDD1.n37 B 0.021581f
C248 VDD1.n38 B 0.021581f
C249 VDD1.n39 B 0.011597f
C250 VDD1.n40 B 0.012279f
C251 VDD1.n41 B 0.02741f
C252 VDD1.n42 B 0.02741f
C253 VDD1.n43 B 0.012279f
C254 VDD1.n44 B 0.011597f
C255 VDD1.n45 B 0.021581f
C256 VDD1.n46 B 0.021581f
C257 VDD1.n47 B 0.011597f
C258 VDD1.n48 B 0.012279f
C259 VDD1.n49 B 0.02741f
C260 VDD1.n50 B 0.02741f
C261 VDD1.n51 B 0.012279f
C262 VDD1.n52 B 0.011597f
C263 VDD1.n53 B 0.021581f
C264 VDD1.n54 B 0.021581f
C265 VDD1.n55 B 0.011597f
C266 VDD1.n56 B 0.012279f
C267 VDD1.n57 B 0.02741f
C268 VDD1.n58 B 0.02741f
C269 VDD1.n59 B 0.012279f
C270 VDD1.n60 B 0.011597f
C271 VDD1.n61 B 0.021581f
C272 VDD1.n62 B 0.021581f
C273 VDD1.n63 B 0.011597f
C274 VDD1.n64 B 0.012279f
C275 VDD1.n65 B 0.02741f
C276 VDD1.n66 B 0.056087f
C277 VDD1.n67 B 0.012279f
C278 VDD1.n68 B 0.022675f
C279 VDD1.n69 B 0.054305f
C280 VDD1.n70 B 0.082185f
C281 VDD1.n71 B 0.029499f
C282 VDD1.n72 B 0.021581f
C283 VDD1.n73 B 0.011597f
C284 VDD1.n74 B 0.02741f
C285 VDD1.n75 B 0.012279f
C286 VDD1.n76 B 0.021581f
C287 VDD1.n77 B 0.011597f
C288 VDD1.n78 B 0.02741f
C289 VDD1.n79 B 0.012279f
C290 VDD1.n80 B 0.021581f
C291 VDD1.n81 B 0.011597f
C292 VDD1.n82 B 0.02741f
C293 VDD1.n83 B 0.012279f
C294 VDD1.n84 B 0.021581f
C295 VDD1.n85 B 0.011597f
C296 VDD1.n86 B 0.02741f
C297 VDD1.n87 B 0.012279f
C298 VDD1.n88 B 0.021581f
C299 VDD1.n89 B 0.011597f
C300 VDD1.n90 B 0.02741f
C301 VDD1.n91 B 0.012279f
C302 VDD1.n92 B 1.24088f
C303 VDD1.n93 B 0.011597f
C304 VDD1.t3 B 0.045074f
C305 VDD1.n94 B 0.131826f
C306 VDD1.n95 B 0.016192f
C307 VDD1.n96 B 0.020558f
C308 VDD1.n97 B 0.02741f
C309 VDD1.n98 B 0.012279f
C310 VDD1.n99 B 0.011597f
C311 VDD1.n100 B 0.021581f
C312 VDD1.n101 B 0.021581f
C313 VDD1.n102 B 0.011597f
C314 VDD1.n103 B 0.012279f
C315 VDD1.n104 B 0.02741f
C316 VDD1.n105 B 0.02741f
C317 VDD1.n106 B 0.012279f
C318 VDD1.n107 B 0.011597f
C319 VDD1.n108 B 0.021581f
C320 VDD1.n109 B 0.021581f
C321 VDD1.n110 B 0.011597f
C322 VDD1.n111 B 0.012279f
C323 VDD1.n112 B 0.02741f
C324 VDD1.n113 B 0.02741f
C325 VDD1.n114 B 0.012279f
C326 VDD1.n115 B 0.011597f
C327 VDD1.n116 B 0.021581f
C328 VDD1.n117 B 0.021581f
C329 VDD1.n118 B 0.011597f
C330 VDD1.n119 B 0.012279f
C331 VDD1.n120 B 0.02741f
C332 VDD1.n121 B 0.02741f
C333 VDD1.n122 B 0.012279f
C334 VDD1.n123 B 0.011597f
C335 VDD1.n124 B 0.021581f
C336 VDD1.n125 B 0.021581f
C337 VDD1.n126 B 0.011597f
C338 VDD1.n127 B 0.012279f
C339 VDD1.n128 B 0.02741f
C340 VDD1.n129 B 0.02741f
C341 VDD1.n130 B 0.012279f
C342 VDD1.n131 B 0.011597f
C343 VDD1.n132 B 0.021581f
C344 VDD1.n133 B 0.021581f
C345 VDD1.n134 B 0.011597f
C346 VDD1.n135 B 0.012279f
C347 VDD1.n136 B 0.02741f
C348 VDD1.n137 B 0.056087f
C349 VDD1.n138 B 0.012279f
C350 VDD1.n139 B 0.022675f
C351 VDD1.n140 B 0.054305f
C352 VDD1.n141 B 0.081434f
C353 VDD1.t4 B 0.227667f
C354 VDD1.t0 B 0.227667f
C355 VDD1.n142 B 2.0539f
C356 VDD1.n143 B 2.77065f
C357 VDD1.t2 B 0.227667f
C358 VDD1.t5 B 0.227667f
C359 VDD1.n144 B 2.04883f
C360 VDD1.n145 B 2.66385f
C361 VTAIL.t4 B 0.250288f
C362 VTAIL.t5 B 0.250288f
C363 VTAIL.n0 B 2.18723f
C364 VTAIL.n1 B 0.442697f
C365 VTAIL.n2 B 0.03243f
C366 VTAIL.n3 B 0.023725f
C367 VTAIL.n4 B 0.012749f
C368 VTAIL.n5 B 0.030133f
C369 VTAIL.n6 B 0.013499f
C370 VTAIL.n7 B 0.023725f
C371 VTAIL.n8 B 0.012749f
C372 VTAIL.n9 B 0.030133f
C373 VTAIL.n10 B 0.013499f
C374 VTAIL.n11 B 0.023725f
C375 VTAIL.n12 B 0.012749f
C376 VTAIL.n13 B 0.030133f
C377 VTAIL.n14 B 0.013499f
C378 VTAIL.n15 B 0.023725f
C379 VTAIL.n16 B 0.012749f
C380 VTAIL.n17 B 0.030133f
C381 VTAIL.n18 B 0.013499f
C382 VTAIL.n19 B 0.023725f
C383 VTAIL.n20 B 0.012749f
C384 VTAIL.n21 B 0.030133f
C385 VTAIL.n22 B 0.013499f
C386 VTAIL.n23 B 1.36417f
C387 VTAIL.n24 B 0.012749f
C388 VTAIL.t7 B 0.049552f
C389 VTAIL.n25 B 0.144924f
C390 VTAIL.n26 B 0.017801f
C391 VTAIL.n27 B 0.0226f
C392 VTAIL.n28 B 0.030133f
C393 VTAIL.n29 B 0.013499f
C394 VTAIL.n30 B 0.012749f
C395 VTAIL.n31 B 0.023725f
C396 VTAIL.n32 B 0.023725f
C397 VTAIL.n33 B 0.012749f
C398 VTAIL.n34 B 0.013499f
C399 VTAIL.n35 B 0.030133f
C400 VTAIL.n36 B 0.030133f
C401 VTAIL.n37 B 0.013499f
C402 VTAIL.n38 B 0.012749f
C403 VTAIL.n39 B 0.023725f
C404 VTAIL.n40 B 0.023725f
C405 VTAIL.n41 B 0.012749f
C406 VTAIL.n42 B 0.013499f
C407 VTAIL.n43 B 0.030133f
C408 VTAIL.n44 B 0.030133f
C409 VTAIL.n45 B 0.013499f
C410 VTAIL.n46 B 0.012749f
C411 VTAIL.n47 B 0.023725f
C412 VTAIL.n48 B 0.023725f
C413 VTAIL.n49 B 0.012749f
C414 VTAIL.n50 B 0.013499f
C415 VTAIL.n51 B 0.030133f
C416 VTAIL.n52 B 0.030133f
C417 VTAIL.n53 B 0.013499f
C418 VTAIL.n54 B 0.012749f
C419 VTAIL.n55 B 0.023725f
C420 VTAIL.n56 B 0.023725f
C421 VTAIL.n57 B 0.012749f
C422 VTAIL.n58 B 0.013499f
C423 VTAIL.n59 B 0.030133f
C424 VTAIL.n60 B 0.030133f
C425 VTAIL.n61 B 0.013499f
C426 VTAIL.n62 B 0.012749f
C427 VTAIL.n63 B 0.023725f
C428 VTAIL.n64 B 0.023725f
C429 VTAIL.n65 B 0.012749f
C430 VTAIL.n66 B 0.013499f
C431 VTAIL.n67 B 0.030133f
C432 VTAIL.n68 B 0.06166f
C433 VTAIL.n69 B 0.013499f
C434 VTAIL.n70 B 0.024928f
C435 VTAIL.n71 B 0.059701f
C436 VTAIL.n72 B 0.063641f
C437 VTAIL.n73 B 0.418757f
C438 VTAIL.t11 B 0.250288f
C439 VTAIL.t9 B 0.250288f
C440 VTAIL.n74 B 2.18723f
C441 VTAIL.n75 B 2.14415f
C442 VTAIL.t3 B 0.250288f
C443 VTAIL.t0 B 0.250288f
C444 VTAIL.n76 B 2.18724f
C445 VTAIL.n77 B 2.14413f
C446 VTAIL.n78 B 0.03243f
C447 VTAIL.n79 B 0.023725f
C448 VTAIL.n80 B 0.012749f
C449 VTAIL.n81 B 0.030133f
C450 VTAIL.n82 B 0.013499f
C451 VTAIL.n83 B 0.023725f
C452 VTAIL.n84 B 0.012749f
C453 VTAIL.n85 B 0.030133f
C454 VTAIL.n86 B 0.013499f
C455 VTAIL.n87 B 0.023725f
C456 VTAIL.n88 B 0.012749f
C457 VTAIL.n89 B 0.030133f
C458 VTAIL.n90 B 0.013499f
C459 VTAIL.n91 B 0.023725f
C460 VTAIL.n92 B 0.012749f
C461 VTAIL.n93 B 0.030133f
C462 VTAIL.n94 B 0.013499f
C463 VTAIL.n95 B 0.023725f
C464 VTAIL.n96 B 0.012749f
C465 VTAIL.n97 B 0.030133f
C466 VTAIL.n98 B 0.013499f
C467 VTAIL.n99 B 1.36417f
C468 VTAIL.n100 B 0.012749f
C469 VTAIL.t1 B 0.049552f
C470 VTAIL.n101 B 0.144924f
C471 VTAIL.n102 B 0.017801f
C472 VTAIL.n103 B 0.0226f
C473 VTAIL.n104 B 0.030133f
C474 VTAIL.n105 B 0.013499f
C475 VTAIL.n106 B 0.012749f
C476 VTAIL.n107 B 0.023725f
C477 VTAIL.n108 B 0.023725f
C478 VTAIL.n109 B 0.012749f
C479 VTAIL.n110 B 0.013499f
C480 VTAIL.n111 B 0.030133f
C481 VTAIL.n112 B 0.030133f
C482 VTAIL.n113 B 0.013499f
C483 VTAIL.n114 B 0.012749f
C484 VTAIL.n115 B 0.023725f
C485 VTAIL.n116 B 0.023725f
C486 VTAIL.n117 B 0.012749f
C487 VTAIL.n118 B 0.013499f
C488 VTAIL.n119 B 0.030133f
C489 VTAIL.n120 B 0.030133f
C490 VTAIL.n121 B 0.013499f
C491 VTAIL.n122 B 0.012749f
C492 VTAIL.n123 B 0.023725f
C493 VTAIL.n124 B 0.023725f
C494 VTAIL.n125 B 0.012749f
C495 VTAIL.n126 B 0.013499f
C496 VTAIL.n127 B 0.030133f
C497 VTAIL.n128 B 0.030133f
C498 VTAIL.n129 B 0.013499f
C499 VTAIL.n130 B 0.012749f
C500 VTAIL.n131 B 0.023725f
C501 VTAIL.n132 B 0.023725f
C502 VTAIL.n133 B 0.012749f
C503 VTAIL.n134 B 0.013499f
C504 VTAIL.n135 B 0.030133f
C505 VTAIL.n136 B 0.030133f
C506 VTAIL.n137 B 0.013499f
C507 VTAIL.n138 B 0.012749f
C508 VTAIL.n139 B 0.023725f
C509 VTAIL.n140 B 0.023725f
C510 VTAIL.n141 B 0.012749f
C511 VTAIL.n142 B 0.013499f
C512 VTAIL.n143 B 0.030133f
C513 VTAIL.n144 B 0.06166f
C514 VTAIL.n145 B 0.013499f
C515 VTAIL.n146 B 0.024928f
C516 VTAIL.n147 B 0.059701f
C517 VTAIL.n148 B 0.063641f
C518 VTAIL.n149 B 0.418757f
C519 VTAIL.t10 B 0.250288f
C520 VTAIL.t6 B 0.250288f
C521 VTAIL.n150 B 2.18724f
C522 VTAIL.n151 B 0.61815f
C523 VTAIL.n152 B 0.03243f
C524 VTAIL.n153 B 0.023725f
C525 VTAIL.n154 B 0.012749f
C526 VTAIL.n155 B 0.030133f
C527 VTAIL.n156 B 0.013499f
C528 VTAIL.n157 B 0.023725f
C529 VTAIL.n158 B 0.012749f
C530 VTAIL.n159 B 0.030133f
C531 VTAIL.n160 B 0.013499f
C532 VTAIL.n161 B 0.023725f
C533 VTAIL.n162 B 0.012749f
C534 VTAIL.n163 B 0.030133f
C535 VTAIL.n164 B 0.013499f
C536 VTAIL.n165 B 0.023725f
C537 VTAIL.n166 B 0.012749f
C538 VTAIL.n167 B 0.030133f
C539 VTAIL.n168 B 0.013499f
C540 VTAIL.n169 B 0.023725f
C541 VTAIL.n170 B 0.012749f
C542 VTAIL.n171 B 0.030133f
C543 VTAIL.n172 B 0.013499f
C544 VTAIL.n173 B 1.36417f
C545 VTAIL.n174 B 0.012749f
C546 VTAIL.t8 B 0.049552f
C547 VTAIL.n175 B 0.144924f
C548 VTAIL.n176 B 0.017801f
C549 VTAIL.n177 B 0.0226f
C550 VTAIL.n178 B 0.030133f
C551 VTAIL.n179 B 0.013499f
C552 VTAIL.n180 B 0.012749f
C553 VTAIL.n181 B 0.023725f
C554 VTAIL.n182 B 0.023725f
C555 VTAIL.n183 B 0.012749f
C556 VTAIL.n184 B 0.013499f
C557 VTAIL.n185 B 0.030133f
C558 VTAIL.n186 B 0.030133f
C559 VTAIL.n187 B 0.013499f
C560 VTAIL.n188 B 0.012749f
C561 VTAIL.n189 B 0.023725f
C562 VTAIL.n190 B 0.023725f
C563 VTAIL.n191 B 0.012749f
C564 VTAIL.n192 B 0.013499f
C565 VTAIL.n193 B 0.030133f
C566 VTAIL.n194 B 0.030133f
C567 VTAIL.n195 B 0.013499f
C568 VTAIL.n196 B 0.012749f
C569 VTAIL.n197 B 0.023725f
C570 VTAIL.n198 B 0.023725f
C571 VTAIL.n199 B 0.012749f
C572 VTAIL.n200 B 0.013499f
C573 VTAIL.n201 B 0.030133f
C574 VTAIL.n202 B 0.030133f
C575 VTAIL.n203 B 0.013499f
C576 VTAIL.n204 B 0.012749f
C577 VTAIL.n205 B 0.023725f
C578 VTAIL.n206 B 0.023725f
C579 VTAIL.n207 B 0.012749f
C580 VTAIL.n208 B 0.013499f
C581 VTAIL.n209 B 0.030133f
C582 VTAIL.n210 B 0.030133f
C583 VTAIL.n211 B 0.013499f
C584 VTAIL.n212 B 0.012749f
C585 VTAIL.n213 B 0.023725f
C586 VTAIL.n214 B 0.023725f
C587 VTAIL.n215 B 0.012749f
C588 VTAIL.n216 B 0.013499f
C589 VTAIL.n217 B 0.030133f
C590 VTAIL.n218 B 0.06166f
C591 VTAIL.n219 B 0.013499f
C592 VTAIL.n220 B 0.024928f
C593 VTAIL.n221 B 0.059701f
C594 VTAIL.n222 B 0.063641f
C595 VTAIL.n223 B 1.70486f
C596 VTAIL.n224 B 0.03243f
C597 VTAIL.n225 B 0.023725f
C598 VTAIL.n226 B 0.012749f
C599 VTAIL.n227 B 0.030133f
C600 VTAIL.n228 B 0.013499f
C601 VTAIL.n229 B 0.023725f
C602 VTAIL.n230 B 0.012749f
C603 VTAIL.n231 B 0.030133f
C604 VTAIL.n232 B 0.013499f
C605 VTAIL.n233 B 0.023725f
C606 VTAIL.n234 B 0.012749f
C607 VTAIL.n235 B 0.030133f
C608 VTAIL.n236 B 0.013499f
C609 VTAIL.n237 B 0.023725f
C610 VTAIL.n238 B 0.012749f
C611 VTAIL.n239 B 0.030133f
C612 VTAIL.n240 B 0.013499f
C613 VTAIL.n241 B 0.023725f
C614 VTAIL.n242 B 0.012749f
C615 VTAIL.n243 B 0.030133f
C616 VTAIL.n244 B 0.013499f
C617 VTAIL.n245 B 1.36417f
C618 VTAIL.n246 B 0.012749f
C619 VTAIL.t2 B 0.049552f
C620 VTAIL.n247 B 0.144924f
C621 VTAIL.n248 B 0.017801f
C622 VTAIL.n249 B 0.0226f
C623 VTAIL.n250 B 0.030133f
C624 VTAIL.n251 B 0.013499f
C625 VTAIL.n252 B 0.012749f
C626 VTAIL.n253 B 0.023725f
C627 VTAIL.n254 B 0.023725f
C628 VTAIL.n255 B 0.012749f
C629 VTAIL.n256 B 0.013499f
C630 VTAIL.n257 B 0.030133f
C631 VTAIL.n258 B 0.030133f
C632 VTAIL.n259 B 0.013499f
C633 VTAIL.n260 B 0.012749f
C634 VTAIL.n261 B 0.023725f
C635 VTAIL.n262 B 0.023725f
C636 VTAIL.n263 B 0.012749f
C637 VTAIL.n264 B 0.013499f
C638 VTAIL.n265 B 0.030133f
C639 VTAIL.n266 B 0.030133f
C640 VTAIL.n267 B 0.013499f
C641 VTAIL.n268 B 0.012749f
C642 VTAIL.n269 B 0.023725f
C643 VTAIL.n270 B 0.023725f
C644 VTAIL.n271 B 0.012749f
C645 VTAIL.n272 B 0.013499f
C646 VTAIL.n273 B 0.030133f
C647 VTAIL.n274 B 0.030133f
C648 VTAIL.n275 B 0.013499f
C649 VTAIL.n276 B 0.012749f
C650 VTAIL.n277 B 0.023725f
C651 VTAIL.n278 B 0.023725f
C652 VTAIL.n279 B 0.012749f
C653 VTAIL.n280 B 0.013499f
C654 VTAIL.n281 B 0.030133f
C655 VTAIL.n282 B 0.030133f
C656 VTAIL.n283 B 0.013499f
C657 VTAIL.n284 B 0.012749f
C658 VTAIL.n285 B 0.023725f
C659 VTAIL.n286 B 0.023725f
C660 VTAIL.n287 B 0.012749f
C661 VTAIL.n288 B 0.013499f
C662 VTAIL.n289 B 0.030133f
C663 VTAIL.n290 B 0.06166f
C664 VTAIL.n291 B 0.013499f
C665 VTAIL.n292 B 0.024928f
C666 VTAIL.n293 B 0.059701f
C667 VTAIL.n294 B 0.063641f
C668 VTAIL.n295 B 1.64044f
C669 VP.t5 B 2.40835f
C670 VP.n0 B 0.926365f
C671 VP.n1 B 0.019946f
C672 VP.n2 B 0.017416f
C673 VP.n3 B 0.019946f
C674 VP.t1 B 2.40835f
C675 VP.n4 B 0.841695f
C676 VP.n5 B 0.019946f
C677 VP.n6 B 0.017416f
C678 VP.n7 B 0.019946f
C679 VP.t2 B 2.40835f
C680 VP.n8 B 0.926365f
C681 VP.t0 B 2.40835f
C682 VP.n9 B 0.926365f
C683 VP.n10 B 0.019946f
C684 VP.n11 B 0.017416f
C685 VP.n12 B 0.019946f
C686 VP.t3 B 2.40835f
C687 VP.n13 B 0.908305f
C688 VP.t4 B 2.66059f
C689 VP.n14 B 0.866557f
C690 VP.n15 B 0.232704f
C691 VP.n16 B 0.027997f
C692 VP.n17 B 0.037174f
C693 VP.n18 B 0.040289f
C694 VP.n19 B 0.019946f
C695 VP.n20 B 0.019946f
C696 VP.n21 B 0.019946f
C697 VP.n22 B 0.037704f
C698 VP.n23 B 0.037174f
C699 VP.n24 B 0.033136f
C700 VP.n25 B 0.032192f
C701 VP.n26 B 1.21916f
C702 VP.n27 B 1.23277f
C703 VP.n28 B 0.032192f
C704 VP.n29 B 0.033136f
C705 VP.n30 B 0.037174f
C706 VP.n31 B 0.037704f
C707 VP.n32 B 0.019946f
C708 VP.n33 B 0.019946f
C709 VP.n34 B 0.019946f
C710 VP.n35 B 0.040289f
C711 VP.n36 B 0.037174f
C712 VP.n37 B 0.027997f
C713 VP.n38 B 0.019946f
C714 VP.n39 B 0.019946f
C715 VP.n40 B 0.027997f
C716 VP.n41 B 0.037174f
C717 VP.n42 B 0.040289f
C718 VP.n43 B 0.019946f
C719 VP.n44 B 0.019946f
C720 VP.n45 B 0.019946f
C721 VP.n46 B 0.037704f
C722 VP.n47 B 0.037174f
C723 VP.n48 B 0.033136f
C724 VP.n49 B 0.032192f
C725 VP.n50 B 0.044446f
.ends

