* NGSPICE file created from diff_pair_sample_0887.ext - technology: sky130A

.subckt diff_pair_sample_0887 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=2.43
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=6.0528 ps=31.82 w=15.52 l=2.43
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=2.43
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=2.43
X4 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=6.0528 ps=31.82 w=15.52 l=2.43
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=0 ps=0 w=15.52 l=2.43
X6 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=6.0528 ps=31.82 w=15.52 l=2.43
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.0528 pd=31.82 as=6.0528 ps=31.82 w=15.52 l=2.43
R0 B.n777 B.n776 585
R1 B.n334 B.n105 585
R2 B.n333 B.n332 585
R3 B.n331 B.n330 585
R4 B.n329 B.n328 585
R5 B.n327 B.n326 585
R6 B.n325 B.n324 585
R7 B.n323 B.n322 585
R8 B.n321 B.n320 585
R9 B.n319 B.n318 585
R10 B.n317 B.n316 585
R11 B.n315 B.n314 585
R12 B.n313 B.n312 585
R13 B.n311 B.n310 585
R14 B.n309 B.n308 585
R15 B.n307 B.n306 585
R16 B.n305 B.n304 585
R17 B.n303 B.n302 585
R18 B.n301 B.n300 585
R19 B.n299 B.n298 585
R20 B.n297 B.n296 585
R21 B.n295 B.n294 585
R22 B.n293 B.n292 585
R23 B.n291 B.n290 585
R24 B.n289 B.n288 585
R25 B.n287 B.n286 585
R26 B.n285 B.n284 585
R27 B.n283 B.n282 585
R28 B.n281 B.n280 585
R29 B.n279 B.n278 585
R30 B.n277 B.n276 585
R31 B.n275 B.n274 585
R32 B.n273 B.n272 585
R33 B.n271 B.n270 585
R34 B.n269 B.n268 585
R35 B.n267 B.n266 585
R36 B.n265 B.n264 585
R37 B.n263 B.n262 585
R38 B.n261 B.n260 585
R39 B.n259 B.n258 585
R40 B.n257 B.n256 585
R41 B.n255 B.n254 585
R42 B.n253 B.n252 585
R43 B.n251 B.n250 585
R44 B.n249 B.n248 585
R45 B.n247 B.n246 585
R46 B.n245 B.n244 585
R47 B.n243 B.n242 585
R48 B.n241 B.n240 585
R49 B.n239 B.n238 585
R50 B.n237 B.n236 585
R51 B.n235 B.n234 585
R52 B.n233 B.n232 585
R53 B.n231 B.n230 585
R54 B.n229 B.n228 585
R55 B.n227 B.n226 585
R56 B.n225 B.n224 585
R57 B.n223 B.n222 585
R58 B.n221 B.n220 585
R59 B.n219 B.n218 585
R60 B.n217 B.n216 585
R61 B.n215 B.n214 585
R62 B.n213 B.n212 585
R63 B.n211 B.n210 585
R64 B.n209 B.n208 585
R65 B.n207 B.n206 585
R66 B.n205 B.n204 585
R67 B.n203 B.n202 585
R68 B.n201 B.n200 585
R69 B.n199 B.n198 585
R70 B.n197 B.n196 585
R71 B.n195 B.n194 585
R72 B.n193 B.n192 585
R73 B.n191 B.n190 585
R74 B.n189 B.n188 585
R75 B.n187 B.n186 585
R76 B.n185 B.n184 585
R77 B.n183 B.n182 585
R78 B.n181 B.n180 585
R79 B.n179 B.n178 585
R80 B.n177 B.n176 585
R81 B.n175 B.n174 585
R82 B.n173 B.n172 585
R83 B.n171 B.n170 585
R84 B.n169 B.n168 585
R85 B.n167 B.n166 585
R86 B.n165 B.n164 585
R87 B.n163 B.n162 585
R88 B.n161 B.n160 585
R89 B.n159 B.n158 585
R90 B.n157 B.n156 585
R91 B.n155 B.n154 585
R92 B.n153 B.n152 585
R93 B.n151 B.n150 585
R94 B.n149 B.n148 585
R95 B.n147 B.n146 585
R96 B.n145 B.n144 585
R97 B.n143 B.n142 585
R98 B.n141 B.n140 585
R99 B.n139 B.n138 585
R100 B.n137 B.n136 585
R101 B.n135 B.n134 585
R102 B.n133 B.n132 585
R103 B.n131 B.n130 585
R104 B.n129 B.n128 585
R105 B.n127 B.n126 585
R106 B.n125 B.n124 585
R107 B.n123 B.n122 585
R108 B.n121 B.n120 585
R109 B.n119 B.n118 585
R110 B.n117 B.n116 585
R111 B.n115 B.n114 585
R112 B.n113 B.n112 585
R113 B.n47 B.n46 585
R114 B.n775 B.n48 585
R115 B.n780 B.n48 585
R116 B.n774 B.n773 585
R117 B.n773 B.n44 585
R118 B.n772 B.n43 585
R119 B.n786 B.n43 585
R120 B.n771 B.n42 585
R121 B.n787 B.n42 585
R122 B.n770 B.n41 585
R123 B.n788 B.n41 585
R124 B.n769 B.n768 585
R125 B.n768 B.n37 585
R126 B.n767 B.n36 585
R127 B.n794 B.n36 585
R128 B.n766 B.n35 585
R129 B.n795 B.n35 585
R130 B.n765 B.n34 585
R131 B.n796 B.n34 585
R132 B.n764 B.n763 585
R133 B.n763 B.n30 585
R134 B.n762 B.n29 585
R135 B.n802 B.n29 585
R136 B.n761 B.n28 585
R137 B.n803 B.n28 585
R138 B.n760 B.n27 585
R139 B.n804 B.n27 585
R140 B.n759 B.n758 585
R141 B.n758 B.n23 585
R142 B.n757 B.n22 585
R143 B.n810 B.n22 585
R144 B.n756 B.n21 585
R145 B.n811 B.n21 585
R146 B.n755 B.n20 585
R147 B.n812 B.n20 585
R148 B.n754 B.n753 585
R149 B.n753 B.n16 585
R150 B.n752 B.n15 585
R151 B.n818 B.n15 585
R152 B.n751 B.n14 585
R153 B.n819 B.n14 585
R154 B.n750 B.n13 585
R155 B.n820 B.n13 585
R156 B.n749 B.n748 585
R157 B.n748 B.n12 585
R158 B.n747 B.n746 585
R159 B.n747 B.n8 585
R160 B.n745 B.n7 585
R161 B.n827 B.n7 585
R162 B.n744 B.n6 585
R163 B.n828 B.n6 585
R164 B.n743 B.n5 585
R165 B.n829 B.n5 585
R166 B.n742 B.n741 585
R167 B.n741 B.n4 585
R168 B.n740 B.n335 585
R169 B.n740 B.n739 585
R170 B.n730 B.n336 585
R171 B.n337 B.n336 585
R172 B.n732 B.n731 585
R173 B.n733 B.n732 585
R174 B.n729 B.n342 585
R175 B.n342 B.n341 585
R176 B.n728 B.n727 585
R177 B.n727 B.n726 585
R178 B.n344 B.n343 585
R179 B.n345 B.n344 585
R180 B.n719 B.n718 585
R181 B.n720 B.n719 585
R182 B.n717 B.n350 585
R183 B.n350 B.n349 585
R184 B.n716 B.n715 585
R185 B.n715 B.n714 585
R186 B.n352 B.n351 585
R187 B.n353 B.n352 585
R188 B.n707 B.n706 585
R189 B.n708 B.n707 585
R190 B.n705 B.n358 585
R191 B.n358 B.n357 585
R192 B.n704 B.n703 585
R193 B.n703 B.n702 585
R194 B.n360 B.n359 585
R195 B.n361 B.n360 585
R196 B.n695 B.n694 585
R197 B.n696 B.n695 585
R198 B.n693 B.n365 585
R199 B.n369 B.n365 585
R200 B.n692 B.n691 585
R201 B.n691 B.n690 585
R202 B.n367 B.n366 585
R203 B.n368 B.n367 585
R204 B.n683 B.n682 585
R205 B.n684 B.n683 585
R206 B.n681 B.n374 585
R207 B.n374 B.n373 585
R208 B.n680 B.n679 585
R209 B.n679 B.n678 585
R210 B.n376 B.n375 585
R211 B.n377 B.n376 585
R212 B.n671 B.n670 585
R213 B.n672 B.n671 585
R214 B.n380 B.n379 585
R215 B.n443 B.n441 585
R216 B.n444 B.n440 585
R217 B.n444 B.n381 585
R218 B.n447 B.n446 585
R219 B.n448 B.n439 585
R220 B.n450 B.n449 585
R221 B.n452 B.n438 585
R222 B.n455 B.n454 585
R223 B.n456 B.n437 585
R224 B.n458 B.n457 585
R225 B.n460 B.n436 585
R226 B.n463 B.n462 585
R227 B.n464 B.n435 585
R228 B.n466 B.n465 585
R229 B.n468 B.n434 585
R230 B.n471 B.n470 585
R231 B.n472 B.n433 585
R232 B.n474 B.n473 585
R233 B.n476 B.n432 585
R234 B.n479 B.n478 585
R235 B.n480 B.n431 585
R236 B.n482 B.n481 585
R237 B.n484 B.n430 585
R238 B.n487 B.n486 585
R239 B.n488 B.n429 585
R240 B.n490 B.n489 585
R241 B.n492 B.n428 585
R242 B.n495 B.n494 585
R243 B.n496 B.n427 585
R244 B.n498 B.n497 585
R245 B.n500 B.n426 585
R246 B.n503 B.n502 585
R247 B.n504 B.n425 585
R248 B.n506 B.n505 585
R249 B.n508 B.n424 585
R250 B.n511 B.n510 585
R251 B.n512 B.n423 585
R252 B.n514 B.n513 585
R253 B.n516 B.n422 585
R254 B.n519 B.n518 585
R255 B.n520 B.n421 585
R256 B.n522 B.n521 585
R257 B.n524 B.n420 585
R258 B.n527 B.n526 585
R259 B.n528 B.n419 585
R260 B.n530 B.n529 585
R261 B.n532 B.n418 585
R262 B.n535 B.n534 585
R263 B.n536 B.n417 585
R264 B.n538 B.n537 585
R265 B.n540 B.n416 585
R266 B.n543 B.n542 585
R267 B.n545 B.n413 585
R268 B.n547 B.n546 585
R269 B.n549 B.n412 585
R270 B.n552 B.n551 585
R271 B.n553 B.n411 585
R272 B.n555 B.n554 585
R273 B.n557 B.n410 585
R274 B.n560 B.n559 585
R275 B.n561 B.n409 585
R276 B.n566 B.n565 585
R277 B.n568 B.n408 585
R278 B.n571 B.n570 585
R279 B.n572 B.n407 585
R280 B.n574 B.n573 585
R281 B.n576 B.n406 585
R282 B.n579 B.n578 585
R283 B.n580 B.n405 585
R284 B.n582 B.n581 585
R285 B.n584 B.n404 585
R286 B.n587 B.n586 585
R287 B.n588 B.n403 585
R288 B.n590 B.n589 585
R289 B.n592 B.n402 585
R290 B.n595 B.n594 585
R291 B.n596 B.n401 585
R292 B.n598 B.n597 585
R293 B.n600 B.n400 585
R294 B.n603 B.n602 585
R295 B.n604 B.n399 585
R296 B.n606 B.n605 585
R297 B.n608 B.n398 585
R298 B.n611 B.n610 585
R299 B.n612 B.n397 585
R300 B.n614 B.n613 585
R301 B.n616 B.n396 585
R302 B.n619 B.n618 585
R303 B.n620 B.n395 585
R304 B.n622 B.n621 585
R305 B.n624 B.n394 585
R306 B.n627 B.n626 585
R307 B.n628 B.n393 585
R308 B.n630 B.n629 585
R309 B.n632 B.n392 585
R310 B.n635 B.n634 585
R311 B.n636 B.n391 585
R312 B.n638 B.n637 585
R313 B.n640 B.n390 585
R314 B.n643 B.n642 585
R315 B.n644 B.n389 585
R316 B.n646 B.n645 585
R317 B.n648 B.n388 585
R318 B.n651 B.n650 585
R319 B.n652 B.n387 585
R320 B.n654 B.n653 585
R321 B.n656 B.n386 585
R322 B.n659 B.n658 585
R323 B.n660 B.n385 585
R324 B.n662 B.n661 585
R325 B.n664 B.n384 585
R326 B.n665 B.n383 585
R327 B.n668 B.n667 585
R328 B.n669 B.n382 585
R329 B.n382 B.n381 585
R330 B.n674 B.n673 585
R331 B.n673 B.n672 585
R332 B.n675 B.n378 585
R333 B.n378 B.n377 585
R334 B.n677 B.n676 585
R335 B.n678 B.n677 585
R336 B.n372 B.n371 585
R337 B.n373 B.n372 585
R338 B.n686 B.n685 585
R339 B.n685 B.n684 585
R340 B.n687 B.n370 585
R341 B.n370 B.n368 585
R342 B.n689 B.n688 585
R343 B.n690 B.n689 585
R344 B.n364 B.n363 585
R345 B.n369 B.n364 585
R346 B.n698 B.n697 585
R347 B.n697 B.n696 585
R348 B.n699 B.n362 585
R349 B.n362 B.n361 585
R350 B.n701 B.n700 585
R351 B.n702 B.n701 585
R352 B.n356 B.n355 585
R353 B.n357 B.n356 585
R354 B.n710 B.n709 585
R355 B.n709 B.n708 585
R356 B.n711 B.n354 585
R357 B.n354 B.n353 585
R358 B.n713 B.n712 585
R359 B.n714 B.n713 585
R360 B.n348 B.n347 585
R361 B.n349 B.n348 585
R362 B.n722 B.n721 585
R363 B.n721 B.n720 585
R364 B.n723 B.n346 585
R365 B.n346 B.n345 585
R366 B.n725 B.n724 585
R367 B.n726 B.n725 585
R368 B.n340 B.n339 585
R369 B.n341 B.n340 585
R370 B.n735 B.n734 585
R371 B.n734 B.n733 585
R372 B.n736 B.n338 585
R373 B.n338 B.n337 585
R374 B.n738 B.n737 585
R375 B.n739 B.n738 585
R376 B.n3 B.n0 585
R377 B.n4 B.n3 585
R378 B.n826 B.n1 585
R379 B.n827 B.n826 585
R380 B.n825 B.n824 585
R381 B.n825 B.n8 585
R382 B.n823 B.n9 585
R383 B.n12 B.n9 585
R384 B.n822 B.n821 585
R385 B.n821 B.n820 585
R386 B.n11 B.n10 585
R387 B.n819 B.n11 585
R388 B.n817 B.n816 585
R389 B.n818 B.n817 585
R390 B.n815 B.n17 585
R391 B.n17 B.n16 585
R392 B.n814 B.n813 585
R393 B.n813 B.n812 585
R394 B.n19 B.n18 585
R395 B.n811 B.n19 585
R396 B.n809 B.n808 585
R397 B.n810 B.n809 585
R398 B.n807 B.n24 585
R399 B.n24 B.n23 585
R400 B.n806 B.n805 585
R401 B.n805 B.n804 585
R402 B.n26 B.n25 585
R403 B.n803 B.n26 585
R404 B.n801 B.n800 585
R405 B.n802 B.n801 585
R406 B.n799 B.n31 585
R407 B.n31 B.n30 585
R408 B.n798 B.n797 585
R409 B.n797 B.n796 585
R410 B.n33 B.n32 585
R411 B.n795 B.n33 585
R412 B.n793 B.n792 585
R413 B.n794 B.n793 585
R414 B.n791 B.n38 585
R415 B.n38 B.n37 585
R416 B.n790 B.n789 585
R417 B.n789 B.n788 585
R418 B.n40 B.n39 585
R419 B.n787 B.n40 585
R420 B.n785 B.n784 585
R421 B.n786 B.n785 585
R422 B.n783 B.n45 585
R423 B.n45 B.n44 585
R424 B.n782 B.n781 585
R425 B.n781 B.n780 585
R426 B.n830 B.n829 585
R427 B.n828 B.n2 585
R428 B.n781 B.n47 434.841
R429 B.n777 B.n48 434.841
R430 B.n671 B.n382 434.841
R431 B.n673 B.n380 434.841
R432 B.n106 B.t7 396.425
R433 B.n562 B.t12 396.425
R434 B.n109 B.t4 396.425
R435 B.n414 B.t15 396.425
R436 B.n109 B.t2 361.699
R437 B.n106 B.t6 361.699
R438 B.n562 B.t9 361.699
R439 B.n414 B.t13 361.699
R440 B.n107 B.t8 342.897
R441 B.n563 B.t11 342.897
R442 B.n110 B.t5 342.897
R443 B.n415 B.t14 342.897
R444 B.n779 B.n778 256.663
R445 B.n779 B.n104 256.663
R446 B.n779 B.n103 256.663
R447 B.n779 B.n102 256.663
R448 B.n779 B.n101 256.663
R449 B.n779 B.n100 256.663
R450 B.n779 B.n99 256.663
R451 B.n779 B.n98 256.663
R452 B.n779 B.n97 256.663
R453 B.n779 B.n96 256.663
R454 B.n779 B.n95 256.663
R455 B.n779 B.n94 256.663
R456 B.n779 B.n93 256.663
R457 B.n779 B.n92 256.663
R458 B.n779 B.n91 256.663
R459 B.n779 B.n90 256.663
R460 B.n779 B.n89 256.663
R461 B.n779 B.n88 256.663
R462 B.n779 B.n87 256.663
R463 B.n779 B.n86 256.663
R464 B.n779 B.n85 256.663
R465 B.n779 B.n84 256.663
R466 B.n779 B.n83 256.663
R467 B.n779 B.n82 256.663
R468 B.n779 B.n81 256.663
R469 B.n779 B.n80 256.663
R470 B.n779 B.n79 256.663
R471 B.n779 B.n78 256.663
R472 B.n779 B.n77 256.663
R473 B.n779 B.n76 256.663
R474 B.n779 B.n75 256.663
R475 B.n779 B.n74 256.663
R476 B.n779 B.n73 256.663
R477 B.n779 B.n72 256.663
R478 B.n779 B.n71 256.663
R479 B.n779 B.n70 256.663
R480 B.n779 B.n69 256.663
R481 B.n779 B.n68 256.663
R482 B.n779 B.n67 256.663
R483 B.n779 B.n66 256.663
R484 B.n779 B.n65 256.663
R485 B.n779 B.n64 256.663
R486 B.n779 B.n63 256.663
R487 B.n779 B.n62 256.663
R488 B.n779 B.n61 256.663
R489 B.n779 B.n60 256.663
R490 B.n779 B.n59 256.663
R491 B.n779 B.n58 256.663
R492 B.n779 B.n57 256.663
R493 B.n779 B.n56 256.663
R494 B.n779 B.n55 256.663
R495 B.n779 B.n54 256.663
R496 B.n779 B.n53 256.663
R497 B.n779 B.n52 256.663
R498 B.n779 B.n51 256.663
R499 B.n779 B.n50 256.663
R500 B.n779 B.n49 256.663
R501 B.n442 B.n381 256.663
R502 B.n445 B.n381 256.663
R503 B.n451 B.n381 256.663
R504 B.n453 B.n381 256.663
R505 B.n459 B.n381 256.663
R506 B.n461 B.n381 256.663
R507 B.n467 B.n381 256.663
R508 B.n469 B.n381 256.663
R509 B.n475 B.n381 256.663
R510 B.n477 B.n381 256.663
R511 B.n483 B.n381 256.663
R512 B.n485 B.n381 256.663
R513 B.n491 B.n381 256.663
R514 B.n493 B.n381 256.663
R515 B.n499 B.n381 256.663
R516 B.n501 B.n381 256.663
R517 B.n507 B.n381 256.663
R518 B.n509 B.n381 256.663
R519 B.n515 B.n381 256.663
R520 B.n517 B.n381 256.663
R521 B.n523 B.n381 256.663
R522 B.n525 B.n381 256.663
R523 B.n531 B.n381 256.663
R524 B.n533 B.n381 256.663
R525 B.n539 B.n381 256.663
R526 B.n541 B.n381 256.663
R527 B.n548 B.n381 256.663
R528 B.n550 B.n381 256.663
R529 B.n556 B.n381 256.663
R530 B.n558 B.n381 256.663
R531 B.n567 B.n381 256.663
R532 B.n569 B.n381 256.663
R533 B.n575 B.n381 256.663
R534 B.n577 B.n381 256.663
R535 B.n583 B.n381 256.663
R536 B.n585 B.n381 256.663
R537 B.n591 B.n381 256.663
R538 B.n593 B.n381 256.663
R539 B.n599 B.n381 256.663
R540 B.n601 B.n381 256.663
R541 B.n607 B.n381 256.663
R542 B.n609 B.n381 256.663
R543 B.n615 B.n381 256.663
R544 B.n617 B.n381 256.663
R545 B.n623 B.n381 256.663
R546 B.n625 B.n381 256.663
R547 B.n631 B.n381 256.663
R548 B.n633 B.n381 256.663
R549 B.n639 B.n381 256.663
R550 B.n641 B.n381 256.663
R551 B.n647 B.n381 256.663
R552 B.n649 B.n381 256.663
R553 B.n655 B.n381 256.663
R554 B.n657 B.n381 256.663
R555 B.n663 B.n381 256.663
R556 B.n666 B.n381 256.663
R557 B.n832 B.n831 256.663
R558 B.n114 B.n113 163.367
R559 B.n118 B.n117 163.367
R560 B.n122 B.n121 163.367
R561 B.n126 B.n125 163.367
R562 B.n130 B.n129 163.367
R563 B.n134 B.n133 163.367
R564 B.n138 B.n137 163.367
R565 B.n142 B.n141 163.367
R566 B.n146 B.n145 163.367
R567 B.n150 B.n149 163.367
R568 B.n154 B.n153 163.367
R569 B.n158 B.n157 163.367
R570 B.n162 B.n161 163.367
R571 B.n166 B.n165 163.367
R572 B.n170 B.n169 163.367
R573 B.n174 B.n173 163.367
R574 B.n178 B.n177 163.367
R575 B.n182 B.n181 163.367
R576 B.n186 B.n185 163.367
R577 B.n190 B.n189 163.367
R578 B.n194 B.n193 163.367
R579 B.n198 B.n197 163.367
R580 B.n202 B.n201 163.367
R581 B.n206 B.n205 163.367
R582 B.n210 B.n209 163.367
R583 B.n214 B.n213 163.367
R584 B.n218 B.n217 163.367
R585 B.n222 B.n221 163.367
R586 B.n226 B.n225 163.367
R587 B.n230 B.n229 163.367
R588 B.n234 B.n233 163.367
R589 B.n238 B.n237 163.367
R590 B.n242 B.n241 163.367
R591 B.n246 B.n245 163.367
R592 B.n250 B.n249 163.367
R593 B.n254 B.n253 163.367
R594 B.n258 B.n257 163.367
R595 B.n262 B.n261 163.367
R596 B.n266 B.n265 163.367
R597 B.n270 B.n269 163.367
R598 B.n274 B.n273 163.367
R599 B.n278 B.n277 163.367
R600 B.n282 B.n281 163.367
R601 B.n286 B.n285 163.367
R602 B.n290 B.n289 163.367
R603 B.n294 B.n293 163.367
R604 B.n298 B.n297 163.367
R605 B.n302 B.n301 163.367
R606 B.n306 B.n305 163.367
R607 B.n310 B.n309 163.367
R608 B.n314 B.n313 163.367
R609 B.n318 B.n317 163.367
R610 B.n322 B.n321 163.367
R611 B.n326 B.n325 163.367
R612 B.n330 B.n329 163.367
R613 B.n332 B.n105 163.367
R614 B.n671 B.n376 163.367
R615 B.n679 B.n376 163.367
R616 B.n679 B.n374 163.367
R617 B.n683 B.n374 163.367
R618 B.n683 B.n367 163.367
R619 B.n691 B.n367 163.367
R620 B.n691 B.n365 163.367
R621 B.n695 B.n365 163.367
R622 B.n695 B.n360 163.367
R623 B.n703 B.n360 163.367
R624 B.n703 B.n358 163.367
R625 B.n707 B.n358 163.367
R626 B.n707 B.n352 163.367
R627 B.n715 B.n352 163.367
R628 B.n715 B.n350 163.367
R629 B.n719 B.n350 163.367
R630 B.n719 B.n344 163.367
R631 B.n727 B.n344 163.367
R632 B.n727 B.n342 163.367
R633 B.n732 B.n342 163.367
R634 B.n732 B.n336 163.367
R635 B.n740 B.n336 163.367
R636 B.n741 B.n740 163.367
R637 B.n741 B.n5 163.367
R638 B.n6 B.n5 163.367
R639 B.n7 B.n6 163.367
R640 B.n747 B.n7 163.367
R641 B.n748 B.n747 163.367
R642 B.n748 B.n13 163.367
R643 B.n14 B.n13 163.367
R644 B.n15 B.n14 163.367
R645 B.n753 B.n15 163.367
R646 B.n753 B.n20 163.367
R647 B.n21 B.n20 163.367
R648 B.n22 B.n21 163.367
R649 B.n758 B.n22 163.367
R650 B.n758 B.n27 163.367
R651 B.n28 B.n27 163.367
R652 B.n29 B.n28 163.367
R653 B.n763 B.n29 163.367
R654 B.n763 B.n34 163.367
R655 B.n35 B.n34 163.367
R656 B.n36 B.n35 163.367
R657 B.n768 B.n36 163.367
R658 B.n768 B.n41 163.367
R659 B.n42 B.n41 163.367
R660 B.n43 B.n42 163.367
R661 B.n773 B.n43 163.367
R662 B.n773 B.n48 163.367
R663 B.n444 B.n443 163.367
R664 B.n446 B.n444 163.367
R665 B.n450 B.n439 163.367
R666 B.n454 B.n452 163.367
R667 B.n458 B.n437 163.367
R668 B.n462 B.n460 163.367
R669 B.n466 B.n435 163.367
R670 B.n470 B.n468 163.367
R671 B.n474 B.n433 163.367
R672 B.n478 B.n476 163.367
R673 B.n482 B.n431 163.367
R674 B.n486 B.n484 163.367
R675 B.n490 B.n429 163.367
R676 B.n494 B.n492 163.367
R677 B.n498 B.n427 163.367
R678 B.n502 B.n500 163.367
R679 B.n506 B.n425 163.367
R680 B.n510 B.n508 163.367
R681 B.n514 B.n423 163.367
R682 B.n518 B.n516 163.367
R683 B.n522 B.n421 163.367
R684 B.n526 B.n524 163.367
R685 B.n530 B.n419 163.367
R686 B.n534 B.n532 163.367
R687 B.n538 B.n417 163.367
R688 B.n542 B.n540 163.367
R689 B.n547 B.n413 163.367
R690 B.n551 B.n549 163.367
R691 B.n555 B.n411 163.367
R692 B.n559 B.n557 163.367
R693 B.n566 B.n409 163.367
R694 B.n570 B.n568 163.367
R695 B.n574 B.n407 163.367
R696 B.n578 B.n576 163.367
R697 B.n582 B.n405 163.367
R698 B.n586 B.n584 163.367
R699 B.n590 B.n403 163.367
R700 B.n594 B.n592 163.367
R701 B.n598 B.n401 163.367
R702 B.n602 B.n600 163.367
R703 B.n606 B.n399 163.367
R704 B.n610 B.n608 163.367
R705 B.n614 B.n397 163.367
R706 B.n618 B.n616 163.367
R707 B.n622 B.n395 163.367
R708 B.n626 B.n624 163.367
R709 B.n630 B.n393 163.367
R710 B.n634 B.n632 163.367
R711 B.n638 B.n391 163.367
R712 B.n642 B.n640 163.367
R713 B.n646 B.n389 163.367
R714 B.n650 B.n648 163.367
R715 B.n654 B.n387 163.367
R716 B.n658 B.n656 163.367
R717 B.n662 B.n385 163.367
R718 B.n665 B.n664 163.367
R719 B.n667 B.n382 163.367
R720 B.n673 B.n378 163.367
R721 B.n677 B.n378 163.367
R722 B.n677 B.n372 163.367
R723 B.n685 B.n372 163.367
R724 B.n685 B.n370 163.367
R725 B.n689 B.n370 163.367
R726 B.n689 B.n364 163.367
R727 B.n697 B.n364 163.367
R728 B.n697 B.n362 163.367
R729 B.n701 B.n362 163.367
R730 B.n701 B.n356 163.367
R731 B.n709 B.n356 163.367
R732 B.n709 B.n354 163.367
R733 B.n713 B.n354 163.367
R734 B.n713 B.n348 163.367
R735 B.n721 B.n348 163.367
R736 B.n721 B.n346 163.367
R737 B.n725 B.n346 163.367
R738 B.n725 B.n340 163.367
R739 B.n734 B.n340 163.367
R740 B.n734 B.n338 163.367
R741 B.n738 B.n338 163.367
R742 B.n738 B.n3 163.367
R743 B.n830 B.n3 163.367
R744 B.n826 B.n2 163.367
R745 B.n826 B.n825 163.367
R746 B.n825 B.n9 163.367
R747 B.n821 B.n9 163.367
R748 B.n821 B.n11 163.367
R749 B.n817 B.n11 163.367
R750 B.n817 B.n17 163.367
R751 B.n813 B.n17 163.367
R752 B.n813 B.n19 163.367
R753 B.n809 B.n19 163.367
R754 B.n809 B.n24 163.367
R755 B.n805 B.n24 163.367
R756 B.n805 B.n26 163.367
R757 B.n801 B.n26 163.367
R758 B.n801 B.n31 163.367
R759 B.n797 B.n31 163.367
R760 B.n797 B.n33 163.367
R761 B.n793 B.n33 163.367
R762 B.n793 B.n38 163.367
R763 B.n789 B.n38 163.367
R764 B.n789 B.n40 163.367
R765 B.n785 B.n40 163.367
R766 B.n785 B.n45 163.367
R767 B.n781 B.n45 163.367
R768 B.n49 B.n47 71.676
R769 B.n114 B.n50 71.676
R770 B.n118 B.n51 71.676
R771 B.n122 B.n52 71.676
R772 B.n126 B.n53 71.676
R773 B.n130 B.n54 71.676
R774 B.n134 B.n55 71.676
R775 B.n138 B.n56 71.676
R776 B.n142 B.n57 71.676
R777 B.n146 B.n58 71.676
R778 B.n150 B.n59 71.676
R779 B.n154 B.n60 71.676
R780 B.n158 B.n61 71.676
R781 B.n162 B.n62 71.676
R782 B.n166 B.n63 71.676
R783 B.n170 B.n64 71.676
R784 B.n174 B.n65 71.676
R785 B.n178 B.n66 71.676
R786 B.n182 B.n67 71.676
R787 B.n186 B.n68 71.676
R788 B.n190 B.n69 71.676
R789 B.n194 B.n70 71.676
R790 B.n198 B.n71 71.676
R791 B.n202 B.n72 71.676
R792 B.n206 B.n73 71.676
R793 B.n210 B.n74 71.676
R794 B.n214 B.n75 71.676
R795 B.n218 B.n76 71.676
R796 B.n222 B.n77 71.676
R797 B.n226 B.n78 71.676
R798 B.n230 B.n79 71.676
R799 B.n234 B.n80 71.676
R800 B.n238 B.n81 71.676
R801 B.n242 B.n82 71.676
R802 B.n246 B.n83 71.676
R803 B.n250 B.n84 71.676
R804 B.n254 B.n85 71.676
R805 B.n258 B.n86 71.676
R806 B.n262 B.n87 71.676
R807 B.n266 B.n88 71.676
R808 B.n270 B.n89 71.676
R809 B.n274 B.n90 71.676
R810 B.n278 B.n91 71.676
R811 B.n282 B.n92 71.676
R812 B.n286 B.n93 71.676
R813 B.n290 B.n94 71.676
R814 B.n294 B.n95 71.676
R815 B.n298 B.n96 71.676
R816 B.n302 B.n97 71.676
R817 B.n306 B.n98 71.676
R818 B.n310 B.n99 71.676
R819 B.n314 B.n100 71.676
R820 B.n318 B.n101 71.676
R821 B.n322 B.n102 71.676
R822 B.n326 B.n103 71.676
R823 B.n330 B.n104 71.676
R824 B.n778 B.n105 71.676
R825 B.n778 B.n777 71.676
R826 B.n332 B.n104 71.676
R827 B.n329 B.n103 71.676
R828 B.n325 B.n102 71.676
R829 B.n321 B.n101 71.676
R830 B.n317 B.n100 71.676
R831 B.n313 B.n99 71.676
R832 B.n309 B.n98 71.676
R833 B.n305 B.n97 71.676
R834 B.n301 B.n96 71.676
R835 B.n297 B.n95 71.676
R836 B.n293 B.n94 71.676
R837 B.n289 B.n93 71.676
R838 B.n285 B.n92 71.676
R839 B.n281 B.n91 71.676
R840 B.n277 B.n90 71.676
R841 B.n273 B.n89 71.676
R842 B.n269 B.n88 71.676
R843 B.n265 B.n87 71.676
R844 B.n261 B.n86 71.676
R845 B.n257 B.n85 71.676
R846 B.n253 B.n84 71.676
R847 B.n249 B.n83 71.676
R848 B.n245 B.n82 71.676
R849 B.n241 B.n81 71.676
R850 B.n237 B.n80 71.676
R851 B.n233 B.n79 71.676
R852 B.n229 B.n78 71.676
R853 B.n225 B.n77 71.676
R854 B.n221 B.n76 71.676
R855 B.n217 B.n75 71.676
R856 B.n213 B.n74 71.676
R857 B.n209 B.n73 71.676
R858 B.n205 B.n72 71.676
R859 B.n201 B.n71 71.676
R860 B.n197 B.n70 71.676
R861 B.n193 B.n69 71.676
R862 B.n189 B.n68 71.676
R863 B.n185 B.n67 71.676
R864 B.n181 B.n66 71.676
R865 B.n177 B.n65 71.676
R866 B.n173 B.n64 71.676
R867 B.n169 B.n63 71.676
R868 B.n165 B.n62 71.676
R869 B.n161 B.n61 71.676
R870 B.n157 B.n60 71.676
R871 B.n153 B.n59 71.676
R872 B.n149 B.n58 71.676
R873 B.n145 B.n57 71.676
R874 B.n141 B.n56 71.676
R875 B.n137 B.n55 71.676
R876 B.n133 B.n54 71.676
R877 B.n129 B.n53 71.676
R878 B.n125 B.n52 71.676
R879 B.n121 B.n51 71.676
R880 B.n117 B.n50 71.676
R881 B.n113 B.n49 71.676
R882 B.n442 B.n380 71.676
R883 B.n446 B.n445 71.676
R884 B.n451 B.n450 71.676
R885 B.n454 B.n453 71.676
R886 B.n459 B.n458 71.676
R887 B.n462 B.n461 71.676
R888 B.n467 B.n466 71.676
R889 B.n470 B.n469 71.676
R890 B.n475 B.n474 71.676
R891 B.n478 B.n477 71.676
R892 B.n483 B.n482 71.676
R893 B.n486 B.n485 71.676
R894 B.n491 B.n490 71.676
R895 B.n494 B.n493 71.676
R896 B.n499 B.n498 71.676
R897 B.n502 B.n501 71.676
R898 B.n507 B.n506 71.676
R899 B.n510 B.n509 71.676
R900 B.n515 B.n514 71.676
R901 B.n518 B.n517 71.676
R902 B.n523 B.n522 71.676
R903 B.n526 B.n525 71.676
R904 B.n531 B.n530 71.676
R905 B.n534 B.n533 71.676
R906 B.n539 B.n538 71.676
R907 B.n542 B.n541 71.676
R908 B.n548 B.n547 71.676
R909 B.n551 B.n550 71.676
R910 B.n556 B.n555 71.676
R911 B.n559 B.n558 71.676
R912 B.n567 B.n566 71.676
R913 B.n570 B.n569 71.676
R914 B.n575 B.n574 71.676
R915 B.n578 B.n577 71.676
R916 B.n583 B.n582 71.676
R917 B.n586 B.n585 71.676
R918 B.n591 B.n590 71.676
R919 B.n594 B.n593 71.676
R920 B.n599 B.n598 71.676
R921 B.n602 B.n601 71.676
R922 B.n607 B.n606 71.676
R923 B.n610 B.n609 71.676
R924 B.n615 B.n614 71.676
R925 B.n618 B.n617 71.676
R926 B.n623 B.n622 71.676
R927 B.n626 B.n625 71.676
R928 B.n631 B.n630 71.676
R929 B.n634 B.n633 71.676
R930 B.n639 B.n638 71.676
R931 B.n642 B.n641 71.676
R932 B.n647 B.n646 71.676
R933 B.n650 B.n649 71.676
R934 B.n655 B.n654 71.676
R935 B.n658 B.n657 71.676
R936 B.n663 B.n662 71.676
R937 B.n666 B.n665 71.676
R938 B.n443 B.n442 71.676
R939 B.n445 B.n439 71.676
R940 B.n452 B.n451 71.676
R941 B.n453 B.n437 71.676
R942 B.n460 B.n459 71.676
R943 B.n461 B.n435 71.676
R944 B.n468 B.n467 71.676
R945 B.n469 B.n433 71.676
R946 B.n476 B.n475 71.676
R947 B.n477 B.n431 71.676
R948 B.n484 B.n483 71.676
R949 B.n485 B.n429 71.676
R950 B.n492 B.n491 71.676
R951 B.n493 B.n427 71.676
R952 B.n500 B.n499 71.676
R953 B.n501 B.n425 71.676
R954 B.n508 B.n507 71.676
R955 B.n509 B.n423 71.676
R956 B.n516 B.n515 71.676
R957 B.n517 B.n421 71.676
R958 B.n524 B.n523 71.676
R959 B.n525 B.n419 71.676
R960 B.n532 B.n531 71.676
R961 B.n533 B.n417 71.676
R962 B.n540 B.n539 71.676
R963 B.n541 B.n413 71.676
R964 B.n549 B.n548 71.676
R965 B.n550 B.n411 71.676
R966 B.n557 B.n556 71.676
R967 B.n558 B.n409 71.676
R968 B.n568 B.n567 71.676
R969 B.n569 B.n407 71.676
R970 B.n576 B.n575 71.676
R971 B.n577 B.n405 71.676
R972 B.n584 B.n583 71.676
R973 B.n585 B.n403 71.676
R974 B.n592 B.n591 71.676
R975 B.n593 B.n401 71.676
R976 B.n600 B.n599 71.676
R977 B.n601 B.n399 71.676
R978 B.n608 B.n607 71.676
R979 B.n609 B.n397 71.676
R980 B.n616 B.n615 71.676
R981 B.n617 B.n395 71.676
R982 B.n624 B.n623 71.676
R983 B.n625 B.n393 71.676
R984 B.n632 B.n631 71.676
R985 B.n633 B.n391 71.676
R986 B.n640 B.n639 71.676
R987 B.n641 B.n389 71.676
R988 B.n648 B.n647 71.676
R989 B.n649 B.n387 71.676
R990 B.n656 B.n655 71.676
R991 B.n657 B.n385 71.676
R992 B.n664 B.n663 71.676
R993 B.n667 B.n666 71.676
R994 B.n831 B.n830 71.676
R995 B.n831 B.n2 71.676
R996 B.n672 B.n381 59.7745
R997 B.n780 B.n779 59.7745
R998 B.n111 B.n110 59.5399
R999 B.n108 B.n107 59.5399
R1000 B.n564 B.n563 59.5399
R1001 B.n544 B.n415 59.5399
R1002 B.n110 B.n109 53.5278
R1003 B.n107 B.n106 53.5278
R1004 B.n563 B.n562 53.5278
R1005 B.n415 B.n414 53.5278
R1006 B.n672 B.n377 35.9707
R1007 B.n678 B.n377 35.9707
R1008 B.n678 B.n373 35.9707
R1009 B.n684 B.n373 35.9707
R1010 B.n684 B.n368 35.9707
R1011 B.n690 B.n368 35.9707
R1012 B.n690 B.n369 35.9707
R1013 B.n696 B.n361 35.9707
R1014 B.n702 B.n361 35.9707
R1015 B.n702 B.n357 35.9707
R1016 B.n708 B.n357 35.9707
R1017 B.n708 B.n353 35.9707
R1018 B.n714 B.n353 35.9707
R1019 B.n714 B.n349 35.9707
R1020 B.n720 B.n349 35.9707
R1021 B.n720 B.n345 35.9707
R1022 B.n726 B.n345 35.9707
R1023 B.n733 B.n341 35.9707
R1024 B.n733 B.n337 35.9707
R1025 B.n739 B.n337 35.9707
R1026 B.n739 B.n4 35.9707
R1027 B.n829 B.n4 35.9707
R1028 B.n829 B.n828 35.9707
R1029 B.n828 B.n827 35.9707
R1030 B.n827 B.n8 35.9707
R1031 B.n12 B.n8 35.9707
R1032 B.n820 B.n12 35.9707
R1033 B.n820 B.n819 35.9707
R1034 B.n818 B.n16 35.9707
R1035 B.n812 B.n16 35.9707
R1036 B.n812 B.n811 35.9707
R1037 B.n811 B.n810 35.9707
R1038 B.n810 B.n23 35.9707
R1039 B.n804 B.n23 35.9707
R1040 B.n804 B.n803 35.9707
R1041 B.n803 B.n802 35.9707
R1042 B.n802 B.n30 35.9707
R1043 B.n796 B.n30 35.9707
R1044 B.n795 B.n794 35.9707
R1045 B.n794 B.n37 35.9707
R1046 B.n788 B.n37 35.9707
R1047 B.n788 B.n787 35.9707
R1048 B.n787 B.n786 35.9707
R1049 B.n786 B.n44 35.9707
R1050 B.n780 B.n44 35.9707
R1051 B.n726 B.t1 30.152
R1052 B.t0 B.n818 30.152
R1053 B.n776 B.n775 28.2542
R1054 B.n674 B.n379 28.2542
R1055 B.n670 B.n669 28.2542
R1056 B.n782 B.n46 28.2542
R1057 B.n369 B.t10 18.5146
R1058 B.t3 B.n795 18.5146
R1059 B B.n832 18.0485
R1060 B.n696 B.t10 17.4566
R1061 B.n796 B.t3 17.4566
R1062 B.n675 B.n674 10.6151
R1063 B.n676 B.n675 10.6151
R1064 B.n676 B.n371 10.6151
R1065 B.n686 B.n371 10.6151
R1066 B.n687 B.n686 10.6151
R1067 B.n688 B.n687 10.6151
R1068 B.n688 B.n363 10.6151
R1069 B.n698 B.n363 10.6151
R1070 B.n699 B.n698 10.6151
R1071 B.n700 B.n699 10.6151
R1072 B.n700 B.n355 10.6151
R1073 B.n710 B.n355 10.6151
R1074 B.n711 B.n710 10.6151
R1075 B.n712 B.n711 10.6151
R1076 B.n712 B.n347 10.6151
R1077 B.n722 B.n347 10.6151
R1078 B.n723 B.n722 10.6151
R1079 B.n724 B.n723 10.6151
R1080 B.n724 B.n339 10.6151
R1081 B.n735 B.n339 10.6151
R1082 B.n736 B.n735 10.6151
R1083 B.n737 B.n736 10.6151
R1084 B.n737 B.n0 10.6151
R1085 B.n441 B.n379 10.6151
R1086 B.n441 B.n440 10.6151
R1087 B.n447 B.n440 10.6151
R1088 B.n448 B.n447 10.6151
R1089 B.n449 B.n448 10.6151
R1090 B.n449 B.n438 10.6151
R1091 B.n455 B.n438 10.6151
R1092 B.n456 B.n455 10.6151
R1093 B.n457 B.n456 10.6151
R1094 B.n457 B.n436 10.6151
R1095 B.n463 B.n436 10.6151
R1096 B.n464 B.n463 10.6151
R1097 B.n465 B.n464 10.6151
R1098 B.n465 B.n434 10.6151
R1099 B.n471 B.n434 10.6151
R1100 B.n472 B.n471 10.6151
R1101 B.n473 B.n472 10.6151
R1102 B.n473 B.n432 10.6151
R1103 B.n479 B.n432 10.6151
R1104 B.n480 B.n479 10.6151
R1105 B.n481 B.n480 10.6151
R1106 B.n481 B.n430 10.6151
R1107 B.n487 B.n430 10.6151
R1108 B.n488 B.n487 10.6151
R1109 B.n489 B.n488 10.6151
R1110 B.n489 B.n428 10.6151
R1111 B.n495 B.n428 10.6151
R1112 B.n496 B.n495 10.6151
R1113 B.n497 B.n496 10.6151
R1114 B.n497 B.n426 10.6151
R1115 B.n503 B.n426 10.6151
R1116 B.n504 B.n503 10.6151
R1117 B.n505 B.n504 10.6151
R1118 B.n505 B.n424 10.6151
R1119 B.n511 B.n424 10.6151
R1120 B.n512 B.n511 10.6151
R1121 B.n513 B.n512 10.6151
R1122 B.n513 B.n422 10.6151
R1123 B.n519 B.n422 10.6151
R1124 B.n520 B.n519 10.6151
R1125 B.n521 B.n520 10.6151
R1126 B.n521 B.n420 10.6151
R1127 B.n527 B.n420 10.6151
R1128 B.n528 B.n527 10.6151
R1129 B.n529 B.n528 10.6151
R1130 B.n529 B.n418 10.6151
R1131 B.n535 B.n418 10.6151
R1132 B.n536 B.n535 10.6151
R1133 B.n537 B.n536 10.6151
R1134 B.n537 B.n416 10.6151
R1135 B.n543 B.n416 10.6151
R1136 B.n546 B.n545 10.6151
R1137 B.n546 B.n412 10.6151
R1138 B.n552 B.n412 10.6151
R1139 B.n553 B.n552 10.6151
R1140 B.n554 B.n553 10.6151
R1141 B.n554 B.n410 10.6151
R1142 B.n560 B.n410 10.6151
R1143 B.n561 B.n560 10.6151
R1144 B.n565 B.n561 10.6151
R1145 B.n571 B.n408 10.6151
R1146 B.n572 B.n571 10.6151
R1147 B.n573 B.n572 10.6151
R1148 B.n573 B.n406 10.6151
R1149 B.n579 B.n406 10.6151
R1150 B.n580 B.n579 10.6151
R1151 B.n581 B.n580 10.6151
R1152 B.n581 B.n404 10.6151
R1153 B.n587 B.n404 10.6151
R1154 B.n588 B.n587 10.6151
R1155 B.n589 B.n588 10.6151
R1156 B.n589 B.n402 10.6151
R1157 B.n595 B.n402 10.6151
R1158 B.n596 B.n595 10.6151
R1159 B.n597 B.n596 10.6151
R1160 B.n597 B.n400 10.6151
R1161 B.n603 B.n400 10.6151
R1162 B.n604 B.n603 10.6151
R1163 B.n605 B.n604 10.6151
R1164 B.n605 B.n398 10.6151
R1165 B.n611 B.n398 10.6151
R1166 B.n612 B.n611 10.6151
R1167 B.n613 B.n612 10.6151
R1168 B.n613 B.n396 10.6151
R1169 B.n619 B.n396 10.6151
R1170 B.n620 B.n619 10.6151
R1171 B.n621 B.n620 10.6151
R1172 B.n621 B.n394 10.6151
R1173 B.n627 B.n394 10.6151
R1174 B.n628 B.n627 10.6151
R1175 B.n629 B.n628 10.6151
R1176 B.n629 B.n392 10.6151
R1177 B.n635 B.n392 10.6151
R1178 B.n636 B.n635 10.6151
R1179 B.n637 B.n636 10.6151
R1180 B.n637 B.n390 10.6151
R1181 B.n643 B.n390 10.6151
R1182 B.n644 B.n643 10.6151
R1183 B.n645 B.n644 10.6151
R1184 B.n645 B.n388 10.6151
R1185 B.n651 B.n388 10.6151
R1186 B.n652 B.n651 10.6151
R1187 B.n653 B.n652 10.6151
R1188 B.n653 B.n386 10.6151
R1189 B.n659 B.n386 10.6151
R1190 B.n660 B.n659 10.6151
R1191 B.n661 B.n660 10.6151
R1192 B.n661 B.n384 10.6151
R1193 B.n384 B.n383 10.6151
R1194 B.n668 B.n383 10.6151
R1195 B.n669 B.n668 10.6151
R1196 B.n670 B.n375 10.6151
R1197 B.n680 B.n375 10.6151
R1198 B.n681 B.n680 10.6151
R1199 B.n682 B.n681 10.6151
R1200 B.n682 B.n366 10.6151
R1201 B.n692 B.n366 10.6151
R1202 B.n693 B.n692 10.6151
R1203 B.n694 B.n693 10.6151
R1204 B.n694 B.n359 10.6151
R1205 B.n704 B.n359 10.6151
R1206 B.n705 B.n704 10.6151
R1207 B.n706 B.n705 10.6151
R1208 B.n706 B.n351 10.6151
R1209 B.n716 B.n351 10.6151
R1210 B.n717 B.n716 10.6151
R1211 B.n718 B.n717 10.6151
R1212 B.n718 B.n343 10.6151
R1213 B.n728 B.n343 10.6151
R1214 B.n729 B.n728 10.6151
R1215 B.n731 B.n729 10.6151
R1216 B.n731 B.n730 10.6151
R1217 B.n730 B.n335 10.6151
R1218 B.n742 B.n335 10.6151
R1219 B.n743 B.n742 10.6151
R1220 B.n744 B.n743 10.6151
R1221 B.n745 B.n744 10.6151
R1222 B.n746 B.n745 10.6151
R1223 B.n749 B.n746 10.6151
R1224 B.n750 B.n749 10.6151
R1225 B.n751 B.n750 10.6151
R1226 B.n752 B.n751 10.6151
R1227 B.n754 B.n752 10.6151
R1228 B.n755 B.n754 10.6151
R1229 B.n756 B.n755 10.6151
R1230 B.n757 B.n756 10.6151
R1231 B.n759 B.n757 10.6151
R1232 B.n760 B.n759 10.6151
R1233 B.n761 B.n760 10.6151
R1234 B.n762 B.n761 10.6151
R1235 B.n764 B.n762 10.6151
R1236 B.n765 B.n764 10.6151
R1237 B.n766 B.n765 10.6151
R1238 B.n767 B.n766 10.6151
R1239 B.n769 B.n767 10.6151
R1240 B.n770 B.n769 10.6151
R1241 B.n771 B.n770 10.6151
R1242 B.n772 B.n771 10.6151
R1243 B.n774 B.n772 10.6151
R1244 B.n775 B.n774 10.6151
R1245 B.n824 B.n1 10.6151
R1246 B.n824 B.n823 10.6151
R1247 B.n823 B.n822 10.6151
R1248 B.n822 B.n10 10.6151
R1249 B.n816 B.n10 10.6151
R1250 B.n816 B.n815 10.6151
R1251 B.n815 B.n814 10.6151
R1252 B.n814 B.n18 10.6151
R1253 B.n808 B.n18 10.6151
R1254 B.n808 B.n807 10.6151
R1255 B.n807 B.n806 10.6151
R1256 B.n806 B.n25 10.6151
R1257 B.n800 B.n25 10.6151
R1258 B.n800 B.n799 10.6151
R1259 B.n799 B.n798 10.6151
R1260 B.n798 B.n32 10.6151
R1261 B.n792 B.n32 10.6151
R1262 B.n792 B.n791 10.6151
R1263 B.n791 B.n790 10.6151
R1264 B.n790 B.n39 10.6151
R1265 B.n784 B.n39 10.6151
R1266 B.n784 B.n783 10.6151
R1267 B.n783 B.n782 10.6151
R1268 B.n112 B.n46 10.6151
R1269 B.n115 B.n112 10.6151
R1270 B.n116 B.n115 10.6151
R1271 B.n119 B.n116 10.6151
R1272 B.n120 B.n119 10.6151
R1273 B.n123 B.n120 10.6151
R1274 B.n124 B.n123 10.6151
R1275 B.n127 B.n124 10.6151
R1276 B.n128 B.n127 10.6151
R1277 B.n131 B.n128 10.6151
R1278 B.n132 B.n131 10.6151
R1279 B.n135 B.n132 10.6151
R1280 B.n136 B.n135 10.6151
R1281 B.n139 B.n136 10.6151
R1282 B.n140 B.n139 10.6151
R1283 B.n143 B.n140 10.6151
R1284 B.n144 B.n143 10.6151
R1285 B.n147 B.n144 10.6151
R1286 B.n148 B.n147 10.6151
R1287 B.n151 B.n148 10.6151
R1288 B.n152 B.n151 10.6151
R1289 B.n155 B.n152 10.6151
R1290 B.n156 B.n155 10.6151
R1291 B.n159 B.n156 10.6151
R1292 B.n160 B.n159 10.6151
R1293 B.n163 B.n160 10.6151
R1294 B.n164 B.n163 10.6151
R1295 B.n167 B.n164 10.6151
R1296 B.n168 B.n167 10.6151
R1297 B.n171 B.n168 10.6151
R1298 B.n172 B.n171 10.6151
R1299 B.n175 B.n172 10.6151
R1300 B.n176 B.n175 10.6151
R1301 B.n179 B.n176 10.6151
R1302 B.n180 B.n179 10.6151
R1303 B.n183 B.n180 10.6151
R1304 B.n184 B.n183 10.6151
R1305 B.n187 B.n184 10.6151
R1306 B.n188 B.n187 10.6151
R1307 B.n191 B.n188 10.6151
R1308 B.n192 B.n191 10.6151
R1309 B.n195 B.n192 10.6151
R1310 B.n196 B.n195 10.6151
R1311 B.n199 B.n196 10.6151
R1312 B.n200 B.n199 10.6151
R1313 B.n203 B.n200 10.6151
R1314 B.n204 B.n203 10.6151
R1315 B.n207 B.n204 10.6151
R1316 B.n208 B.n207 10.6151
R1317 B.n211 B.n208 10.6151
R1318 B.n212 B.n211 10.6151
R1319 B.n216 B.n215 10.6151
R1320 B.n219 B.n216 10.6151
R1321 B.n220 B.n219 10.6151
R1322 B.n223 B.n220 10.6151
R1323 B.n224 B.n223 10.6151
R1324 B.n227 B.n224 10.6151
R1325 B.n228 B.n227 10.6151
R1326 B.n231 B.n228 10.6151
R1327 B.n232 B.n231 10.6151
R1328 B.n236 B.n235 10.6151
R1329 B.n239 B.n236 10.6151
R1330 B.n240 B.n239 10.6151
R1331 B.n243 B.n240 10.6151
R1332 B.n244 B.n243 10.6151
R1333 B.n247 B.n244 10.6151
R1334 B.n248 B.n247 10.6151
R1335 B.n251 B.n248 10.6151
R1336 B.n252 B.n251 10.6151
R1337 B.n255 B.n252 10.6151
R1338 B.n256 B.n255 10.6151
R1339 B.n259 B.n256 10.6151
R1340 B.n260 B.n259 10.6151
R1341 B.n263 B.n260 10.6151
R1342 B.n264 B.n263 10.6151
R1343 B.n267 B.n264 10.6151
R1344 B.n268 B.n267 10.6151
R1345 B.n271 B.n268 10.6151
R1346 B.n272 B.n271 10.6151
R1347 B.n275 B.n272 10.6151
R1348 B.n276 B.n275 10.6151
R1349 B.n279 B.n276 10.6151
R1350 B.n280 B.n279 10.6151
R1351 B.n283 B.n280 10.6151
R1352 B.n284 B.n283 10.6151
R1353 B.n287 B.n284 10.6151
R1354 B.n288 B.n287 10.6151
R1355 B.n291 B.n288 10.6151
R1356 B.n292 B.n291 10.6151
R1357 B.n295 B.n292 10.6151
R1358 B.n296 B.n295 10.6151
R1359 B.n299 B.n296 10.6151
R1360 B.n300 B.n299 10.6151
R1361 B.n303 B.n300 10.6151
R1362 B.n304 B.n303 10.6151
R1363 B.n307 B.n304 10.6151
R1364 B.n308 B.n307 10.6151
R1365 B.n311 B.n308 10.6151
R1366 B.n312 B.n311 10.6151
R1367 B.n315 B.n312 10.6151
R1368 B.n316 B.n315 10.6151
R1369 B.n319 B.n316 10.6151
R1370 B.n320 B.n319 10.6151
R1371 B.n323 B.n320 10.6151
R1372 B.n324 B.n323 10.6151
R1373 B.n327 B.n324 10.6151
R1374 B.n328 B.n327 10.6151
R1375 B.n331 B.n328 10.6151
R1376 B.n333 B.n331 10.6151
R1377 B.n334 B.n333 10.6151
R1378 B.n776 B.n334 10.6151
R1379 B.n544 B.n543 9.36635
R1380 B.n564 B.n408 9.36635
R1381 B.n212 B.n111 9.36635
R1382 B.n235 B.n108 9.36635
R1383 B.n832 B.n0 8.11757
R1384 B.n832 B.n1 8.11757
R1385 B.t1 B.n341 5.81921
R1386 B.n819 B.t0 5.81921
R1387 B.n545 B.n544 1.24928
R1388 B.n565 B.n564 1.24928
R1389 B.n215 B.n111 1.24928
R1390 B.n232 B.n108 1.24928
R1391 VP.n0 VP.t1 250.011
R1392 VP.n0 VP.t0 203.138
R1393 VP VP.n0 0.336784
R1394 VTAIL.n338 VTAIL.n258 289.615
R1395 VTAIL.n80 VTAIL.n0 289.615
R1396 VTAIL.n252 VTAIL.n172 289.615
R1397 VTAIL.n166 VTAIL.n86 289.615
R1398 VTAIL.n287 VTAIL.n286 185
R1399 VTAIL.n289 VTAIL.n288 185
R1400 VTAIL.n282 VTAIL.n281 185
R1401 VTAIL.n295 VTAIL.n294 185
R1402 VTAIL.n297 VTAIL.n296 185
R1403 VTAIL.n278 VTAIL.n277 185
R1404 VTAIL.n303 VTAIL.n302 185
R1405 VTAIL.n305 VTAIL.n304 185
R1406 VTAIL.n274 VTAIL.n273 185
R1407 VTAIL.n311 VTAIL.n310 185
R1408 VTAIL.n313 VTAIL.n312 185
R1409 VTAIL.n270 VTAIL.n269 185
R1410 VTAIL.n319 VTAIL.n318 185
R1411 VTAIL.n321 VTAIL.n320 185
R1412 VTAIL.n266 VTAIL.n265 185
R1413 VTAIL.n328 VTAIL.n327 185
R1414 VTAIL.n329 VTAIL.n264 185
R1415 VTAIL.n331 VTAIL.n330 185
R1416 VTAIL.n262 VTAIL.n261 185
R1417 VTAIL.n337 VTAIL.n336 185
R1418 VTAIL.n339 VTAIL.n338 185
R1419 VTAIL.n29 VTAIL.n28 185
R1420 VTAIL.n31 VTAIL.n30 185
R1421 VTAIL.n24 VTAIL.n23 185
R1422 VTAIL.n37 VTAIL.n36 185
R1423 VTAIL.n39 VTAIL.n38 185
R1424 VTAIL.n20 VTAIL.n19 185
R1425 VTAIL.n45 VTAIL.n44 185
R1426 VTAIL.n47 VTAIL.n46 185
R1427 VTAIL.n16 VTAIL.n15 185
R1428 VTAIL.n53 VTAIL.n52 185
R1429 VTAIL.n55 VTAIL.n54 185
R1430 VTAIL.n12 VTAIL.n11 185
R1431 VTAIL.n61 VTAIL.n60 185
R1432 VTAIL.n63 VTAIL.n62 185
R1433 VTAIL.n8 VTAIL.n7 185
R1434 VTAIL.n70 VTAIL.n69 185
R1435 VTAIL.n71 VTAIL.n6 185
R1436 VTAIL.n73 VTAIL.n72 185
R1437 VTAIL.n4 VTAIL.n3 185
R1438 VTAIL.n79 VTAIL.n78 185
R1439 VTAIL.n81 VTAIL.n80 185
R1440 VTAIL.n253 VTAIL.n252 185
R1441 VTAIL.n251 VTAIL.n250 185
R1442 VTAIL.n176 VTAIL.n175 185
R1443 VTAIL.n180 VTAIL.n178 185
R1444 VTAIL.n245 VTAIL.n244 185
R1445 VTAIL.n243 VTAIL.n242 185
R1446 VTAIL.n182 VTAIL.n181 185
R1447 VTAIL.n237 VTAIL.n236 185
R1448 VTAIL.n235 VTAIL.n234 185
R1449 VTAIL.n186 VTAIL.n185 185
R1450 VTAIL.n229 VTAIL.n228 185
R1451 VTAIL.n227 VTAIL.n226 185
R1452 VTAIL.n190 VTAIL.n189 185
R1453 VTAIL.n221 VTAIL.n220 185
R1454 VTAIL.n219 VTAIL.n218 185
R1455 VTAIL.n194 VTAIL.n193 185
R1456 VTAIL.n213 VTAIL.n212 185
R1457 VTAIL.n211 VTAIL.n210 185
R1458 VTAIL.n198 VTAIL.n197 185
R1459 VTAIL.n205 VTAIL.n204 185
R1460 VTAIL.n203 VTAIL.n202 185
R1461 VTAIL.n167 VTAIL.n166 185
R1462 VTAIL.n165 VTAIL.n164 185
R1463 VTAIL.n90 VTAIL.n89 185
R1464 VTAIL.n94 VTAIL.n92 185
R1465 VTAIL.n159 VTAIL.n158 185
R1466 VTAIL.n157 VTAIL.n156 185
R1467 VTAIL.n96 VTAIL.n95 185
R1468 VTAIL.n151 VTAIL.n150 185
R1469 VTAIL.n149 VTAIL.n148 185
R1470 VTAIL.n100 VTAIL.n99 185
R1471 VTAIL.n143 VTAIL.n142 185
R1472 VTAIL.n141 VTAIL.n140 185
R1473 VTAIL.n104 VTAIL.n103 185
R1474 VTAIL.n135 VTAIL.n134 185
R1475 VTAIL.n133 VTAIL.n132 185
R1476 VTAIL.n108 VTAIL.n107 185
R1477 VTAIL.n127 VTAIL.n126 185
R1478 VTAIL.n125 VTAIL.n124 185
R1479 VTAIL.n112 VTAIL.n111 185
R1480 VTAIL.n119 VTAIL.n118 185
R1481 VTAIL.n117 VTAIL.n116 185
R1482 VTAIL.n285 VTAIL.t0 147.659
R1483 VTAIL.n27 VTAIL.t2 147.659
R1484 VTAIL.n201 VTAIL.t3 147.659
R1485 VTAIL.n115 VTAIL.t1 147.659
R1486 VTAIL.n288 VTAIL.n287 104.615
R1487 VTAIL.n288 VTAIL.n281 104.615
R1488 VTAIL.n295 VTAIL.n281 104.615
R1489 VTAIL.n296 VTAIL.n295 104.615
R1490 VTAIL.n296 VTAIL.n277 104.615
R1491 VTAIL.n303 VTAIL.n277 104.615
R1492 VTAIL.n304 VTAIL.n303 104.615
R1493 VTAIL.n304 VTAIL.n273 104.615
R1494 VTAIL.n311 VTAIL.n273 104.615
R1495 VTAIL.n312 VTAIL.n311 104.615
R1496 VTAIL.n312 VTAIL.n269 104.615
R1497 VTAIL.n319 VTAIL.n269 104.615
R1498 VTAIL.n320 VTAIL.n319 104.615
R1499 VTAIL.n320 VTAIL.n265 104.615
R1500 VTAIL.n328 VTAIL.n265 104.615
R1501 VTAIL.n329 VTAIL.n328 104.615
R1502 VTAIL.n330 VTAIL.n329 104.615
R1503 VTAIL.n330 VTAIL.n261 104.615
R1504 VTAIL.n337 VTAIL.n261 104.615
R1505 VTAIL.n338 VTAIL.n337 104.615
R1506 VTAIL.n30 VTAIL.n29 104.615
R1507 VTAIL.n30 VTAIL.n23 104.615
R1508 VTAIL.n37 VTAIL.n23 104.615
R1509 VTAIL.n38 VTAIL.n37 104.615
R1510 VTAIL.n38 VTAIL.n19 104.615
R1511 VTAIL.n45 VTAIL.n19 104.615
R1512 VTAIL.n46 VTAIL.n45 104.615
R1513 VTAIL.n46 VTAIL.n15 104.615
R1514 VTAIL.n53 VTAIL.n15 104.615
R1515 VTAIL.n54 VTAIL.n53 104.615
R1516 VTAIL.n54 VTAIL.n11 104.615
R1517 VTAIL.n61 VTAIL.n11 104.615
R1518 VTAIL.n62 VTAIL.n61 104.615
R1519 VTAIL.n62 VTAIL.n7 104.615
R1520 VTAIL.n70 VTAIL.n7 104.615
R1521 VTAIL.n71 VTAIL.n70 104.615
R1522 VTAIL.n72 VTAIL.n71 104.615
R1523 VTAIL.n72 VTAIL.n3 104.615
R1524 VTAIL.n79 VTAIL.n3 104.615
R1525 VTAIL.n80 VTAIL.n79 104.615
R1526 VTAIL.n252 VTAIL.n251 104.615
R1527 VTAIL.n251 VTAIL.n175 104.615
R1528 VTAIL.n180 VTAIL.n175 104.615
R1529 VTAIL.n244 VTAIL.n180 104.615
R1530 VTAIL.n244 VTAIL.n243 104.615
R1531 VTAIL.n243 VTAIL.n181 104.615
R1532 VTAIL.n236 VTAIL.n181 104.615
R1533 VTAIL.n236 VTAIL.n235 104.615
R1534 VTAIL.n235 VTAIL.n185 104.615
R1535 VTAIL.n228 VTAIL.n185 104.615
R1536 VTAIL.n228 VTAIL.n227 104.615
R1537 VTAIL.n227 VTAIL.n189 104.615
R1538 VTAIL.n220 VTAIL.n189 104.615
R1539 VTAIL.n220 VTAIL.n219 104.615
R1540 VTAIL.n219 VTAIL.n193 104.615
R1541 VTAIL.n212 VTAIL.n193 104.615
R1542 VTAIL.n212 VTAIL.n211 104.615
R1543 VTAIL.n211 VTAIL.n197 104.615
R1544 VTAIL.n204 VTAIL.n197 104.615
R1545 VTAIL.n204 VTAIL.n203 104.615
R1546 VTAIL.n166 VTAIL.n165 104.615
R1547 VTAIL.n165 VTAIL.n89 104.615
R1548 VTAIL.n94 VTAIL.n89 104.615
R1549 VTAIL.n158 VTAIL.n94 104.615
R1550 VTAIL.n158 VTAIL.n157 104.615
R1551 VTAIL.n157 VTAIL.n95 104.615
R1552 VTAIL.n150 VTAIL.n95 104.615
R1553 VTAIL.n150 VTAIL.n149 104.615
R1554 VTAIL.n149 VTAIL.n99 104.615
R1555 VTAIL.n142 VTAIL.n99 104.615
R1556 VTAIL.n142 VTAIL.n141 104.615
R1557 VTAIL.n141 VTAIL.n103 104.615
R1558 VTAIL.n134 VTAIL.n103 104.615
R1559 VTAIL.n134 VTAIL.n133 104.615
R1560 VTAIL.n133 VTAIL.n107 104.615
R1561 VTAIL.n126 VTAIL.n107 104.615
R1562 VTAIL.n126 VTAIL.n125 104.615
R1563 VTAIL.n125 VTAIL.n111 104.615
R1564 VTAIL.n118 VTAIL.n111 104.615
R1565 VTAIL.n118 VTAIL.n117 104.615
R1566 VTAIL.n287 VTAIL.t0 52.3082
R1567 VTAIL.n29 VTAIL.t2 52.3082
R1568 VTAIL.n203 VTAIL.t3 52.3082
R1569 VTAIL.n117 VTAIL.t1 52.3082
R1570 VTAIL.n343 VTAIL.n342 35.2884
R1571 VTAIL.n85 VTAIL.n84 35.2884
R1572 VTAIL.n257 VTAIL.n256 35.2884
R1573 VTAIL.n171 VTAIL.n170 35.2884
R1574 VTAIL.n171 VTAIL.n85 30.5048
R1575 VTAIL.n343 VTAIL.n257 28.1255
R1576 VTAIL.n286 VTAIL.n285 15.6677
R1577 VTAIL.n28 VTAIL.n27 15.6677
R1578 VTAIL.n202 VTAIL.n201 15.6677
R1579 VTAIL.n116 VTAIL.n115 15.6677
R1580 VTAIL.n331 VTAIL.n262 13.1884
R1581 VTAIL.n73 VTAIL.n4 13.1884
R1582 VTAIL.n178 VTAIL.n176 13.1884
R1583 VTAIL.n92 VTAIL.n90 13.1884
R1584 VTAIL.n289 VTAIL.n284 12.8005
R1585 VTAIL.n332 VTAIL.n264 12.8005
R1586 VTAIL.n336 VTAIL.n335 12.8005
R1587 VTAIL.n31 VTAIL.n26 12.8005
R1588 VTAIL.n74 VTAIL.n6 12.8005
R1589 VTAIL.n78 VTAIL.n77 12.8005
R1590 VTAIL.n250 VTAIL.n249 12.8005
R1591 VTAIL.n246 VTAIL.n245 12.8005
R1592 VTAIL.n205 VTAIL.n200 12.8005
R1593 VTAIL.n164 VTAIL.n163 12.8005
R1594 VTAIL.n160 VTAIL.n159 12.8005
R1595 VTAIL.n119 VTAIL.n114 12.8005
R1596 VTAIL.n290 VTAIL.n282 12.0247
R1597 VTAIL.n327 VTAIL.n326 12.0247
R1598 VTAIL.n339 VTAIL.n260 12.0247
R1599 VTAIL.n32 VTAIL.n24 12.0247
R1600 VTAIL.n69 VTAIL.n68 12.0247
R1601 VTAIL.n81 VTAIL.n2 12.0247
R1602 VTAIL.n253 VTAIL.n174 12.0247
R1603 VTAIL.n242 VTAIL.n179 12.0247
R1604 VTAIL.n206 VTAIL.n198 12.0247
R1605 VTAIL.n167 VTAIL.n88 12.0247
R1606 VTAIL.n156 VTAIL.n93 12.0247
R1607 VTAIL.n120 VTAIL.n112 12.0247
R1608 VTAIL.n294 VTAIL.n293 11.249
R1609 VTAIL.n325 VTAIL.n266 11.249
R1610 VTAIL.n340 VTAIL.n258 11.249
R1611 VTAIL.n36 VTAIL.n35 11.249
R1612 VTAIL.n67 VTAIL.n8 11.249
R1613 VTAIL.n82 VTAIL.n0 11.249
R1614 VTAIL.n254 VTAIL.n172 11.249
R1615 VTAIL.n241 VTAIL.n182 11.249
R1616 VTAIL.n210 VTAIL.n209 11.249
R1617 VTAIL.n168 VTAIL.n86 11.249
R1618 VTAIL.n155 VTAIL.n96 11.249
R1619 VTAIL.n124 VTAIL.n123 11.249
R1620 VTAIL.n297 VTAIL.n280 10.4732
R1621 VTAIL.n322 VTAIL.n321 10.4732
R1622 VTAIL.n39 VTAIL.n22 10.4732
R1623 VTAIL.n64 VTAIL.n63 10.4732
R1624 VTAIL.n238 VTAIL.n237 10.4732
R1625 VTAIL.n213 VTAIL.n196 10.4732
R1626 VTAIL.n152 VTAIL.n151 10.4732
R1627 VTAIL.n127 VTAIL.n110 10.4732
R1628 VTAIL.n298 VTAIL.n278 9.69747
R1629 VTAIL.n318 VTAIL.n268 9.69747
R1630 VTAIL.n40 VTAIL.n20 9.69747
R1631 VTAIL.n60 VTAIL.n10 9.69747
R1632 VTAIL.n234 VTAIL.n184 9.69747
R1633 VTAIL.n214 VTAIL.n194 9.69747
R1634 VTAIL.n148 VTAIL.n98 9.69747
R1635 VTAIL.n128 VTAIL.n108 9.69747
R1636 VTAIL.n342 VTAIL.n341 9.45567
R1637 VTAIL.n84 VTAIL.n83 9.45567
R1638 VTAIL.n256 VTAIL.n255 9.45567
R1639 VTAIL.n170 VTAIL.n169 9.45567
R1640 VTAIL.n341 VTAIL.n340 9.3005
R1641 VTAIL.n260 VTAIL.n259 9.3005
R1642 VTAIL.n335 VTAIL.n334 9.3005
R1643 VTAIL.n307 VTAIL.n306 9.3005
R1644 VTAIL.n276 VTAIL.n275 9.3005
R1645 VTAIL.n301 VTAIL.n300 9.3005
R1646 VTAIL.n299 VTAIL.n298 9.3005
R1647 VTAIL.n280 VTAIL.n279 9.3005
R1648 VTAIL.n293 VTAIL.n292 9.3005
R1649 VTAIL.n291 VTAIL.n290 9.3005
R1650 VTAIL.n284 VTAIL.n283 9.3005
R1651 VTAIL.n309 VTAIL.n308 9.3005
R1652 VTAIL.n272 VTAIL.n271 9.3005
R1653 VTAIL.n315 VTAIL.n314 9.3005
R1654 VTAIL.n317 VTAIL.n316 9.3005
R1655 VTAIL.n268 VTAIL.n267 9.3005
R1656 VTAIL.n323 VTAIL.n322 9.3005
R1657 VTAIL.n325 VTAIL.n324 9.3005
R1658 VTAIL.n326 VTAIL.n263 9.3005
R1659 VTAIL.n333 VTAIL.n332 9.3005
R1660 VTAIL.n83 VTAIL.n82 9.3005
R1661 VTAIL.n2 VTAIL.n1 9.3005
R1662 VTAIL.n77 VTAIL.n76 9.3005
R1663 VTAIL.n49 VTAIL.n48 9.3005
R1664 VTAIL.n18 VTAIL.n17 9.3005
R1665 VTAIL.n43 VTAIL.n42 9.3005
R1666 VTAIL.n41 VTAIL.n40 9.3005
R1667 VTAIL.n22 VTAIL.n21 9.3005
R1668 VTAIL.n35 VTAIL.n34 9.3005
R1669 VTAIL.n33 VTAIL.n32 9.3005
R1670 VTAIL.n26 VTAIL.n25 9.3005
R1671 VTAIL.n51 VTAIL.n50 9.3005
R1672 VTAIL.n14 VTAIL.n13 9.3005
R1673 VTAIL.n57 VTAIL.n56 9.3005
R1674 VTAIL.n59 VTAIL.n58 9.3005
R1675 VTAIL.n10 VTAIL.n9 9.3005
R1676 VTAIL.n65 VTAIL.n64 9.3005
R1677 VTAIL.n67 VTAIL.n66 9.3005
R1678 VTAIL.n68 VTAIL.n5 9.3005
R1679 VTAIL.n75 VTAIL.n74 9.3005
R1680 VTAIL.n188 VTAIL.n187 9.3005
R1681 VTAIL.n231 VTAIL.n230 9.3005
R1682 VTAIL.n233 VTAIL.n232 9.3005
R1683 VTAIL.n184 VTAIL.n183 9.3005
R1684 VTAIL.n239 VTAIL.n238 9.3005
R1685 VTAIL.n241 VTAIL.n240 9.3005
R1686 VTAIL.n179 VTAIL.n177 9.3005
R1687 VTAIL.n247 VTAIL.n246 9.3005
R1688 VTAIL.n255 VTAIL.n254 9.3005
R1689 VTAIL.n174 VTAIL.n173 9.3005
R1690 VTAIL.n249 VTAIL.n248 9.3005
R1691 VTAIL.n225 VTAIL.n224 9.3005
R1692 VTAIL.n223 VTAIL.n222 9.3005
R1693 VTAIL.n192 VTAIL.n191 9.3005
R1694 VTAIL.n217 VTAIL.n216 9.3005
R1695 VTAIL.n215 VTAIL.n214 9.3005
R1696 VTAIL.n196 VTAIL.n195 9.3005
R1697 VTAIL.n209 VTAIL.n208 9.3005
R1698 VTAIL.n207 VTAIL.n206 9.3005
R1699 VTAIL.n200 VTAIL.n199 9.3005
R1700 VTAIL.n102 VTAIL.n101 9.3005
R1701 VTAIL.n145 VTAIL.n144 9.3005
R1702 VTAIL.n147 VTAIL.n146 9.3005
R1703 VTAIL.n98 VTAIL.n97 9.3005
R1704 VTAIL.n153 VTAIL.n152 9.3005
R1705 VTAIL.n155 VTAIL.n154 9.3005
R1706 VTAIL.n93 VTAIL.n91 9.3005
R1707 VTAIL.n161 VTAIL.n160 9.3005
R1708 VTAIL.n169 VTAIL.n168 9.3005
R1709 VTAIL.n88 VTAIL.n87 9.3005
R1710 VTAIL.n163 VTAIL.n162 9.3005
R1711 VTAIL.n139 VTAIL.n138 9.3005
R1712 VTAIL.n137 VTAIL.n136 9.3005
R1713 VTAIL.n106 VTAIL.n105 9.3005
R1714 VTAIL.n131 VTAIL.n130 9.3005
R1715 VTAIL.n129 VTAIL.n128 9.3005
R1716 VTAIL.n110 VTAIL.n109 9.3005
R1717 VTAIL.n123 VTAIL.n122 9.3005
R1718 VTAIL.n121 VTAIL.n120 9.3005
R1719 VTAIL.n114 VTAIL.n113 9.3005
R1720 VTAIL.n302 VTAIL.n301 8.92171
R1721 VTAIL.n317 VTAIL.n270 8.92171
R1722 VTAIL.n44 VTAIL.n43 8.92171
R1723 VTAIL.n59 VTAIL.n12 8.92171
R1724 VTAIL.n233 VTAIL.n186 8.92171
R1725 VTAIL.n218 VTAIL.n217 8.92171
R1726 VTAIL.n147 VTAIL.n100 8.92171
R1727 VTAIL.n132 VTAIL.n131 8.92171
R1728 VTAIL.n305 VTAIL.n276 8.14595
R1729 VTAIL.n314 VTAIL.n313 8.14595
R1730 VTAIL.n47 VTAIL.n18 8.14595
R1731 VTAIL.n56 VTAIL.n55 8.14595
R1732 VTAIL.n230 VTAIL.n229 8.14595
R1733 VTAIL.n221 VTAIL.n192 8.14595
R1734 VTAIL.n144 VTAIL.n143 8.14595
R1735 VTAIL.n135 VTAIL.n106 8.14595
R1736 VTAIL.n306 VTAIL.n274 7.3702
R1737 VTAIL.n310 VTAIL.n272 7.3702
R1738 VTAIL.n48 VTAIL.n16 7.3702
R1739 VTAIL.n52 VTAIL.n14 7.3702
R1740 VTAIL.n226 VTAIL.n188 7.3702
R1741 VTAIL.n222 VTAIL.n190 7.3702
R1742 VTAIL.n140 VTAIL.n102 7.3702
R1743 VTAIL.n136 VTAIL.n104 7.3702
R1744 VTAIL.n309 VTAIL.n274 6.59444
R1745 VTAIL.n310 VTAIL.n309 6.59444
R1746 VTAIL.n51 VTAIL.n16 6.59444
R1747 VTAIL.n52 VTAIL.n51 6.59444
R1748 VTAIL.n226 VTAIL.n225 6.59444
R1749 VTAIL.n225 VTAIL.n190 6.59444
R1750 VTAIL.n140 VTAIL.n139 6.59444
R1751 VTAIL.n139 VTAIL.n104 6.59444
R1752 VTAIL.n306 VTAIL.n305 5.81868
R1753 VTAIL.n313 VTAIL.n272 5.81868
R1754 VTAIL.n48 VTAIL.n47 5.81868
R1755 VTAIL.n55 VTAIL.n14 5.81868
R1756 VTAIL.n229 VTAIL.n188 5.81868
R1757 VTAIL.n222 VTAIL.n221 5.81868
R1758 VTAIL.n143 VTAIL.n102 5.81868
R1759 VTAIL.n136 VTAIL.n135 5.81868
R1760 VTAIL.n302 VTAIL.n276 5.04292
R1761 VTAIL.n314 VTAIL.n270 5.04292
R1762 VTAIL.n44 VTAIL.n18 5.04292
R1763 VTAIL.n56 VTAIL.n12 5.04292
R1764 VTAIL.n230 VTAIL.n186 5.04292
R1765 VTAIL.n218 VTAIL.n192 5.04292
R1766 VTAIL.n144 VTAIL.n100 5.04292
R1767 VTAIL.n132 VTAIL.n106 5.04292
R1768 VTAIL.n285 VTAIL.n283 4.38563
R1769 VTAIL.n27 VTAIL.n25 4.38563
R1770 VTAIL.n201 VTAIL.n199 4.38563
R1771 VTAIL.n115 VTAIL.n113 4.38563
R1772 VTAIL.n301 VTAIL.n278 4.26717
R1773 VTAIL.n318 VTAIL.n317 4.26717
R1774 VTAIL.n43 VTAIL.n20 4.26717
R1775 VTAIL.n60 VTAIL.n59 4.26717
R1776 VTAIL.n234 VTAIL.n233 4.26717
R1777 VTAIL.n217 VTAIL.n194 4.26717
R1778 VTAIL.n148 VTAIL.n147 4.26717
R1779 VTAIL.n131 VTAIL.n108 4.26717
R1780 VTAIL.n298 VTAIL.n297 3.49141
R1781 VTAIL.n321 VTAIL.n268 3.49141
R1782 VTAIL.n40 VTAIL.n39 3.49141
R1783 VTAIL.n63 VTAIL.n10 3.49141
R1784 VTAIL.n237 VTAIL.n184 3.49141
R1785 VTAIL.n214 VTAIL.n213 3.49141
R1786 VTAIL.n151 VTAIL.n98 3.49141
R1787 VTAIL.n128 VTAIL.n127 3.49141
R1788 VTAIL.n294 VTAIL.n280 2.71565
R1789 VTAIL.n322 VTAIL.n266 2.71565
R1790 VTAIL.n342 VTAIL.n258 2.71565
R1791 VTAIL.n36 VTAIL.n22 2.71565
R1792 VTAIL.n64 VTAIL.n8 2.71565
R1793 VTAIL.n84 VTAIL.n0 2.71565
R1794 VTAIL.n256 VTAIL.n172 2.71565
R1795 VTAIL.n238 VTAIL.n182 2.71565
R1796 VTAIL.n210 VTAIL.n196 2.71565
R1797 VTAIL.n170 VTAIL.n86 2.71565
R1798 VTAIL.n152 VTAIL.n96 2.71565
R1799 VTAIL.n124 VTAIL.n110 2.71565
R1800 VTAIL.n293 VTAIL.n282 1.93989
R1801 VTAIL.n327 VTAIL.n325 1.93989
R1802 VTAIL.n340 VTAIL.n339 1.93989
R1803 VTAIL.n35 VTAIL.n24 1.93989
R1804 VTAIL.n69 VTAIL.n67 1.93989
R1805 VTAIL.n82 VTAIL.n81 1.93989
R1806 VTAIL.n254 VTAIL.n253 1.93989
R1807 VTAIL.n242 VTAIL.n241 1.93989
R1808 VTAIL.n209 VTAIL.n198 1.93989
R1809 VTAIL.n168 VTAIL.n167 1.93989
R1810 VTAIL.n156 VTAIL.n155 1.93989
R1811 VTAIL.n123 VTAIL.n112 1.93989
R1812 VTAIL.n257 VTAIL.n171 1.65998
R1813 VTAIL.n290 VTAIL.n289 1.16414
R1814 VTAIL.n326 VTAIL.n264 1.16414
R1815 VTAIL.n336 VTAIL.n260 1.16414
R1816 VTAIL.n32 VTAIL.n31 1.16414
R1817 VTAIL.n68 VTAIL.n6 1.16414
R1818 VTAIL.n78 VTAIL.n2 1.16414
R1819 VTAIL.n250 VTAIL.n174 1.16414
R1820 VTAIL.n245 VTAIL.n179 1.16414
R1821 VTAIL.n206 VTAIL.n205 1.16414
R1822 VTAIL.n164 VTAIL.n88 1.16414
R1823 VTAIL.n159 VTAIL.n93 1.16414
R1824 VTAIL.n120 VTAIL.n119 1.16414
R1825 VTAIL VTAIL.n85 1.12334
R1826 VTAIL VTAIL.n343 0.537138
R1827 VTAIL.n286 VTAIL.n284 0.388379
R1828 VTAIL.n332 VTAIL.n331 0.388379
R1829 VTAIL.n335 VTAIL.n262 0.388379
R1830 VTAIL.n28 VTAIL.n26 0.388379
R1831 VTAIL.n74 VTAIL.n73 0.388379
R1832 VTAIL.n77 VTAIL.n4 0.388379
R1833 VTAIL.n249 VTAIL.n176 0.388379
R1834 VTAIL.n246 VTAIL.n178 0.388379
R1835 VTAIL.n202 VTAIL.n200 0.388379
R1836 VTAIL.n163 VTAIL.n90 0.388379
R1837 VTAIL.n160 VTAIL.n92 0.388379
R1838 VTAIL.n116 VTAIL.n114 0.388379
R1839 VTAIL.n291 VTAIL.n283 0.155672
R1840 VTAIL.n292 VTAIL.n291 0.155672
R1841 VTAIL.n292 VTAIL.n279 0.155672
R1842 VTAIL.n299 VTAIL.n279 0.155672
R1843 VTAIL.n300 VTAIL.n299 0.155672
R1844 VTAIL.n300 VTAIL.n275 0.155672
R1845 VTAIL.n307 VTAIL.n275 0.155672
R1846 VTAIL.n308 VTAIL.n307 0.155672
R1847 VTAIL.n308 VTAIL.n271 0.155672
R1848 VTAIL.n315 VTAIL.n271 0.155672
R1849 VTAIL.n316 VTAIL.n315 0.155672
R1850 VTAIL.n316 VTAIL.n267 0.155672
R1851 VTAIL.n323 VTAIL.n267 0.155672
R1852 VTAIL.n324 VTAIL.n323 0.155672
R1853 VTAIL.n324 VTAIL.n263 0.155672
R1854 VTAIL.n333 VTAIL.n263 0.155672
R1855 VTAIL.n334 VTAIL.n333 0.155672
R1856 VTAIL.n334 VTAIL.n259 0.155672
R1857 VTAIL.n341 VTAIL.n259 0.155672
R1858 VTAIL.n33 VTAIL.n25 0.155672
R1859 VTAIL.n34 VTAIL.n33 0.155672
R1860 VTAIL.n34 VTAIL.n21 0.155672
R1861 VTAIL.n41 VTAIL.n21 0.155672
R1862 VTAIL.n42 VTAIL.n41 0.155672
R1863 VTAIL.n42 VTAIL.n17 0.155672
R1864 VTAIL.n49 VTAIL.n17 0.155672
R1865 VTAIL.n50 VTAIL.n49 0.155672
R1866 VTAIL.n50 VTAIL.n13 0.155672
R1867 VTAIL.n57 VTAIL.n13 0.155672
R1868 VTAIL.n58 VTAIL.n57 0.155672
R1869 VTAIL.n58 VTAIL.n9 0.155672
R1870 VTAIL.n65 VTAIL.n9 0.155672
R1871 VTAIL.n66 VTAIL.n65 0.155672
R1872 VTAIL.n66 VTAIL.n5 0.155672
R1873 VTAIL.n75 VTAIL.n5 0.155672
R1874 VTAIL.n76 VTAIL.n75 0.155672
R1875 VTAIL.n76 VTAIL.n1 0.155672
R1876 VTAIL.n83 VTAIL.n1 0.155672
R1877 VTAIL.n255 VTAIL.n173 0.155672
R1878 VTAIL.n248 VTAIL.n173 0.155672
R1879 VTAIL.n248 VTAIL.n247 0.155672
R1880 VTAIL.n247 VTAIL.n177 0.155672
R1881 VTAIL.n240 VTAIL.n177 0.155672
R1882 VTAIL.n240 VTAIL.n239 0.155672
R1883 VTAIL.n239 VTAIL.n183 0.155672
R1884 VTAIL.n232 VTAIL.n183 0.155672
R1885 VTAIL.n232 VTAIL.n231 0.155672
R1886 VTAIL.n231 VTAIL.n187 0.155672
R1887 VTAIL.n224 VTAIL.n187 0.155672
R1888 VTAIL.n224 VTAIL.n223 0.155672
R1889 VTAIL.n223 VTAIL.n191 0.155672
R1890 VTAIL.n216 VTAIL.n191 0.155672
R1891 VTAIL.n216 VTAIL.n215 0.155672
R1892 VTAIL.n215 VTAIL.n195 0.155672
R1893 VTAIL.n208 VTAIL.n195 0.155672
R1894 VTAIL.n208 VTAIL.n207 0.155672
R1895 VTAIL.n207 VTAIL.n199 0.155672
R1896 VTAIL.n169 VTAIL.n87 0.155672
R1897 VTAIL.n162 VTAIL.n87 0.155672
R1898 VTAIL.n162 VTAIL.n161 0.155672
R1899 VTAIL.n161 VTAIL.n91 0.155672
R1900 VTAIL.n154 VTAIL.n91 0.155672
R1901 VTAIL.n154 VTAIL.n153 0.155672
R1902 VTAIL.n153 VTAIL.n97 0.155672
R1903 VTAIL.n146 VTAIL.n97 0.155672
R1904 VTAIL.n146 VTAIL.n145 0.155672
R1905 VTAIL.n145 VTAIL.n101 0.155672
R1906 VTAIL.n138 VTAIL.n101 0.155672
R1907 VTAIL.n138 VTAIL.n137 0.155672
R1908 VTAIL.n137 VTAIL.n105 0.155672
R1909 VTAIL.n130 VTAIL.n105 0.155672
R1910 VTAIL.n130 VTAIL.n129 0.155672
R1911 VTAIL.n129 VTAIL.n109 0.155672
R1912 VTAIL.n122 VTAIL.n109 0.155672
R1913 VTAIL.n122 VTAIL.n121 0.155672
R1914 VTAIL.n121 VTAIL.n113 0.155672
R1915 VDD1.n80 VDD1.n0 289.615
R1916 VDD1.n165 VDD1.n85 289.615
R1917 VDD1.n81 VDD1.n80 185
R1918 VDD1.n79 VDD1.n78 185
R1919 VDD1.n4 VDD1.n3 185
R1920 VDD1.n8 VDD1.n6 185
R1921 VDD1.n73 VDD1.n72 185
R1922 VDD1.n71 VDD1.n70 185
R1923 VDD1.n10 VDD1.n9 185
R1924 VDD1.n65 VDD1.n64 185
R1925 VDD1.n63 VDD1.n62 185
R1926 VDD1.n14 VDD1.n13 185
R1927 VDD1.n57 VDD1.n56 185
R1928 VDD1.n55 VDD1.n54 185
R1929 VDD1.n18 VDD1.n17 185
R1930 VDD1.n49 VDD1.n48 185
R1931 VDD1.n47 VDD1.n46 185
R1932 VDD1.n22 VDD1.n21 185
R1933 VDD1.n41 VDD1.n40 185
R1934 VDD1.n39 VDD1.n38 185
R1935 VDD1.n26 VDD1.n25 185
R1936 VDD1.n33 VDD1.n32 185
R1937 VDD1.n31 VDD1.n30 185
R1938 VDD1.n114 VDD1.n113 185
R1939 VDD1.n116 VDD1.n115 185
R1940 VDD1.n109 VDD1.n108 185
R1941 VDD1.n122 VDD1.n121 185
R1942 VDD1.n124 VDD1.n123 185
R1943 VDD1.n105 VDD1.n104 185
R1944 VDD1.n130 VDD1.n129 185
R1945 VDD1.n132 VDD1.n131 185
R1946 VDD1.n101 VDD1.n100 185
R1947 VDD1.n138 VDD1.n137 185
R1948 VDD1.n140 VDD1.n139 185
R1949 VDD1.n97 VDD1.n96 185
R1950 VDD1.n146 VDD1.n145 185
R1951 VDD1.n148 VDD1.n147 185
R1952 VDD1.n93 VDD1.n92 185
R1953 VDD1.n155 VDD1.n154 185
R1954 VDD1.n156 VDD1.n91 185
R1955 VDD1.n158 VDD1.n157 185
R1956 VDD1.n89 VDD1.n88 185
R1957 VDD1.n164 VDD1.n163 185
R1958 VDD1.n166 VDD1.n165 185
R1959 VDD1.n29 VDD1.t0 147.659
R1960 VDD1.n112 VDD1.t1 147.659
R1961 VDD1.n80 VDD1.n79 104.615
R1962 VDD1.n79 VDD1.n3 104.615
R1963 VDD1.n8 VDD1.n3 104.615
R1964 VDD1.n72 VDD1.n8 104.615
R1965 VDD1.n72 VDD1.n71 104.615
R1966 VDD1.n71 VDD1.n9 104.615
R1967 VDD1.n64 VDD1.n9 104.615
R1968 VDD1.n64 VDD1.n63 104.615
R1969 VDD1.n63 VDD1.n13 104.615
R1970 VDD1.n56 VDD1.n13 104.615
R1971 VDD1.n56 VDD1.n55 104.615
R1972 VDD1.n55 VDD1.n17 104.615
R1973 VDD1.n48 VDD1.n17 104.615
R1974 VDD1.n48 VDD1.n47 104.615
R1975 VDD1.n47 VDD1.n21 104.615
R1976 VDD1.n40 VDD1.n21 104.615
R1977 VDD1.n40 VDD1.n39 104.615
R1978 VDD1.n39 VDD1.n25 104.615
R1979 VDD1.n32 VDD1.n25 104.615
R1980 VDD1.n32 VDD1.n31 104.615
R1981 VDD1.n115 VDD1.n114 104.615
R1982 VDD1.n115 VDD1.n108 104.615
R1983 VDD1.n122 VDD1.n108 104.615
R1984 VDD1.n123 VDD1.n122 104.615
R1985 VDD1.n123 VDD1.n104 104.615
R1986 VDD1.n130 VDD1.n104 104.615
R1987 VDD1.n131 VDD1.n130 104.615
R1988 VDD1.n131 VDD1.n100 104.615
R1989 VDD1.n138 VDD1.n100 104.615
R1990 VDD1.n139 VDD1.n138 104.615
R1991 VDD1.n139 VDD1.n96 104.615
R1992 VDD1.n146 VDD1.n96 104.615
R1993 VDD1.n147 VDD1.n146 104.615
R1994 VDD1.n147 VDD1.n92 104.615
R1995 VDD1.n155 VDD1.n92 104.615
R1996 VDD1.n156 VDD1.n155 104.615
R1997 VDD1.n157 VDD1.n156 104.615
R1998 VDD1.n157 VDD1.n88 104.615
R1999 VDD1.n164 VDD1.n88 104.615
R2000 VDD1.n165 VDD1.n164 104.615
R2001 VDD1 VDD1.n169 94.8842
R2002 VDD1 VDD1.n84 52.6202
R2003 VDD1.n31 VDD1.t0 52.3082
R2004 VDD1.n114 VDD1.t1 52.3082
R2005 VDD1.n30 VDD1.n29 15.6677
R2006 VDD1.n113 VDD1.n112 15.6677
R2007 VDD1.n6 VDD1.n4 13.1884
R2008 VDD1.n158 VDD1.n89 13.1884
R2009 VDD1.n78 VDD1.n77 12.8005
R2010 VDD1.n74 VDD1.n73 12.8005
R2011 VDD1.n33 VDD1.n28 12.8005
R2012 VDD1.n116 VDD1.n111 12.8005
R2013 VDD1.n159 VDD1.n91 12.8005
R2014 VDD1.n163 VDD1.n162 12.8005
R2015 VDD1.n81 VDD1.n2 12.0247
R2016 VDD1.n70 VDD1.n7 12.0247
R2017 VDD1.n34 VDD1.n26 12.0247
R2018 VDD1.n117 VDD1.n109 12.0247
R2019 VDD1.n154 VDD1.n153 12.0247
R2020 VDD1.n166 VDD1.n87 12.0247
R2021 VDD1.n82 VDD1.n0 11.249
R2022 VDD1.n69 VDD1.n10 11.249
R2023 VDD1.n38 VDD1.n37 11.249
R2024 VDD1.n121 VDD1.n120 11.249
R2025 VDD1.n152 VDD1.n93 11.249
R2026 VDD1.n167 VDD1.n85 11.249
R2027 VDD1.n66 VDD1.n65 10.4732
R2028 VDD1.n41 VDD1.n24 10.4732
R2029 VDD1.n124 VDD1.n107 10.4732
R2030 VDD1.n149 VDD1.n148 10.4732
R2031 VDD1.n62 VDD1.n12 9.69747
R2032 VDD1.n42 VDD1.n22 9.69747
R2033 VDD1.n125 VDD1.n105 9.69747
R2034 VDD1.n145 VDD1.n95 9.69747
R2035 VDD1.n84 VDD1.n83 9.45567
R2036 VDD1.n169 VDD1.n168 9.45567
R2037 VDD1.n16 VDD1.n15 9.3005
R2038 VDD1.n59 VDD1.n58 9.3005
R2039 VDD1.n61 VDD1.n60 9.3005
R2040 VDD1.n12 VDD1.n11 9.3005
R2041 VDD1.n67 VDD1.n66 9.3005
R2042 VDD1.n69 VDD1.n68 9.3005
R2043 VDD1.n7 VDD1.n5 9.3005
R2044 VDD1.n75 VDD1.n74 9.3005
R2045 VDD1.n83 VDD1.n82 9.3005
R2046 VDD1.n2 VDD1.n1 9.3005
R2047 VDD1.n77 VDD1.n76 9.3005
R2048 VDD1.n53 VDD1.n52 9.3005
R2049 VDD1.n51 VDD1.n50 9.3005
R2050 VDD1.n20 VDD1.n19 9.3005
R2051 VDD1.n45 VDD1.n44 9.3005
R2052 VDD1.n43 VDD1.n42 9.3005
R2053 VDD1.n24 VDD1.n23 9.3005
R2054 VDD1.n37 VDD1.n36 9.3005
R2055 VDD1.n35 VDD1.n34 9.3005
R2056 VDD1.n28 VDD1.n27 9.3005
R2057 VDD1.n168 VDD1.n167 9.3005
R2058 VDD1.n87 VDD1.n86 9.3005
R2059 VDD1.n162 VDD1.n161 9.3005
R2060 VDD1.n134 VDD1.n133 9.3005
R2061 VDD1.n103 VDD1.n102 9.3005
R2062 VDD1.n128 VDD1.n127 9.3005
R2063 VDD1.n126 VDD1.n125 9.3005
R2064 VDD1.n107 VDD1.n106 9.3005
R2065 VDD1.n120 VDD1.n119 9.3005
R2066 VDD1.n118 VDD1.n117 9.3005
R2067 VDD1.n111 VDD1.n110 9.3005
R2068 VDD1.n136 VDD1.n135 9.3005
R2069 VDD1.n99 VDD1.n98 9.3005
R2070 VDD1.n142 VDD1.n141 9.3005
R2071 VDD1.n144 VDD1.n143 9.3005
R2072 VDD1.n95 VDD1.n94 9.3005
R2073 VDD1.n150 VDD1.n149 9.3005
R2074 VDD1.n152 VDD1.n151 9.3005
R2075 VDD1.n153 VDD1.n90 9.3005
R2076 VDD1.n160 VDD1.n159 9.3005
R2077 VDD1.n61 VDD1.n14 8.92171
R2078 VDD1.n46 VDD1.n45 8.92171
R2079 VDD1.n129 VDD1.n128 8.92171
R2080 VDD1.n144 VDD1.n97 8.92171
R2081 VDD1.n58 VDD1.n57 8.14595
R2082 VDD1.n49 VDD1.n20 8.14595
R2083 VDD1.n132 VDD1.n103 8.14595
R2084 VDD1.n141 VDD1.n140 8.14595
R2085 VDD1.n54 VDD1.n16 7.3702
R2086 VDD1.n50 VDD1.n18 7.3702
R2087 VDD1.n133 VDD1.n101 7.3702
R2088 VDD1.n137 VDD1.n99 7.3702
R2089 VDD1.n54 VDD1.n53 6.59444
R2090 VDD1.n53 VDD1.n18 6.59444
R2091 VDD1.n136 VDD1.n101 6.59444
R2092 VDD1.n137 VDD1.n136 6.59444
R2093 VDD1.n57 VDD1.n16 5.81868
R2094 VDD1.n50 VDD1.n49 5.81868
R2095 VDD1.n133 VDD1.n132 5.81868
R2096 VDD1.n140 VDD1.n99 5.81868
R2097 VDD1.n58 VDD1.n14 5.04292
R2098 VDD1.n46 VDD1.n20 5.04292
R2099 VDD1.n129 VDD1.n103 5.04292
R2100 VDD1.n141 VDD1.n97 5.04292
R2101 VDD1.n29 VDD1.n27 4.38563
R2102 VDD1.n112 VDD1.n110 4.38563
R2103 VDD1.n62 VDD1.n61 4.26717
R2104 VDD1.n45 VDD1.n22 4.26717
R2105 VDD1.n128 VDD1.n105 4.26717
R2106 VDD1.n145 VDD1.n144 4.26717
R2107 VDD1.n65 VDD1.n12 3.49141
R2108 VDD1.n42 VDD1.n41 3.49141
R2109 VDD1.n125 VDD1.n124 3.49141
R2110 VDD1.n148 VDD1.n95 3.49141
R2111 VDD1.n84 VDD1.n0 2.71565
R2112 VDD1.n66 VDD1.n10 2.71565
R2113 VDD1.n38 VDD1.n24 2.71565
R2114 VDD1.n121 VDD1.n107 2.71565
R2115 VDD1.n149 VDD1.n93 2.71565
R2116 VDD1.n169 VDD1.n85 2.71565
R2117 VDD1.n82 VDD1.n81 1.93989
R2118 VDD1.n70 VDD1.n69 1.93989
R2119 VDD1.n37 VDD1.n26 1.93989
R2120 VDD1.n120 VDD1.n109 1.93989
R2121 VDD1.n154 VDD1.n152 1.93989
R2122 VDD1.n167 VDD1.n166 1.93989
R2123 VDD1.n78 VDD1.n2 1.16414
R2124 VDD1.n73 VDD1.n7 1.16414
R2125 VDD1.n34 VDD1.n33 1.16414
R2126 VDD1.n117 VDD1.n116 1.16414
R2127 VDD1.n153 VDD1.n91 1.16414
R2128 VDD1.n163 VDD1.n87 1.16414
R2129 VDD1.n77 VDD1.n4 0.388379
R2130 VDD1.n74 VDD1.n6 0.388379
R2131 VDD1.n30 VDD1.n28 0.388379
R2132 VDD1.n113 VDD1.n111 0.388379
R2133 VDD1.n159 VDD1.n158 0.388379
R2134 VDD1.n162 VDD1.n89 0.388379
R2135 VDD1.n83 VDD1.n1 0.155672
R2136 VDD1.n76 VDD1.n1 0.155672
R2137 VDD1.n76 VDD1.n75 0.155672
R2138 VDD1.n75 VDD1.n5 0.155672
R2139 VDD1.n68 VDD1.n5 0.155672
R2140 VDD1.n68 VDD1.n67 0.155672
R2141 VDD1.n67 VDD1.n11 0.155672
R2142 VDD1.n60 VDD1.n11 0.155672
R2143 VDD1.n60 VDD1.n59 0.155672
R2144 VDD1.n59 VDD1.n15 0.155672
R2145 VDD1.n52 VDD1.n15 0.155672
R2146 VDD1.n52 VDD1.n51 0.155672
R2147 VDD1.n51 VDD1.n19 0.155672
R2148 VDD1.n44 VDD1.n19 0.155672
R2149 VDD1.n44 VDD1.n43 0.155672
R2150 VDD1.n43 VDD1.n23 0.155672
R2151 VDD1.n36 VDD1.n23 0.155672
R2152 VDD1.n36 VDD1.n35 0.155672
R2153 VDD1.n35 VDD1.n27 0.155672
R2154 VDD1.n118 VDD1.n110 0.155672
R2155 VDD1.n119 VDD1.n118 0.155672
R2156 VDD1.n119 VDD1.n106 0.155672
R2157 VDD1.n126 VDD1.n106 0.155672
R2158 VDD1.n127 VDD1.n126 0.155672
R2159 VDD1.n127 VDD1.n102 0.155672
R2160 VDD1.n134 VDD1.n102 0.155672
R2161 VDD1.n135 VDD1.n134 0.155672
R2162 VDD1.n135 VDD1.n98 0.155672
R2163 VDD1.n142 VDD1.n98 0.155672
R2164 VDD1.n143 VDD1.n142 0.155672
R2165 VDD1.n143 VDD1.n94 0.155672
R2166 VDD1.n150 VDD1.n94 0.155672
R2167 VDD1.n151 VDD1.n150 0.155672
R2168 VDD1.n151 VDD1.n90 0.155672
R2169 VDD1.n160 VDD1.n90 0.155672
R2170 VDD1.n161 VDD1.n160 0.155672
R2171 VDD1.n161 VDD1.n86 0.155672
R2172 VDD1.n168 VDD1.n86 0.155672
R2173 VN VN.t0 250.107
R2174 VN VN.t1 203.475
R2175 VDD2.n165 VDD2.n85 289.615
R2176 VDD2.n80 VDD2.n0 289.615
R2177 VDD2.n166 VDD2.n165 185
R2178 VDD2.n164 VDD2.n163 185
R2179 VDD2.n89 VDD2.n88 185
R2180 VDD2.n93 VDD2.n91 185
R2181 VDD2.n158 VDD2.n157 185
R2182 VDD2.n156 VDD2.n155 185
R2183 VDD2.n95 VDD2.n94 185
R2184 VDD2.n150 VDD2.n149 185
R2185 VDD2.n148 VDD2.n147 185
R2186 VDD2.n99 VDD2.n98 185
R2187 VDD2.n142 VDD2.n141 185
R2188 VDD2.n140 VDD2.n139 185
R2189 VDD2.n103 VDD2.n102 185
R2190 VDD2.n134 VDD2.n133 185
R2191 VDD2.n132 VDD2.n131 185
R2192 VDD2.n107 VDD2.n106 185
R2193 VDD2.n126 VDD2.n125 185
R2194 VDD2.n124 VDD2.n123 185
R2195 VDD2.n111 VDD2.n110 185
R2196 VDD2.n118 VDD2.n117 185
R2197 VDD2.n116 VDD2.n115 185
R2198 VDD2.n29 VDD2.n28 185
R2199 VDD2.n31 VDD2.n30 185
R2200 VDD2.n24 VDD2.n23 185
R2201 VDD2.n37 VDD2.n36 185
R2202 VDD2.n39 VDD2.n38 185
R2203 VDD2.n20 VDD2.n19 185
R2204 VDD2.n45 VDD2.n44 185
R2205 VDD2.n47 VDD2.n46 185
R2206 VDD2.n16 VDD2.n15 185
R2207 VDD2.n53 VDD2.n52 185
R2208 VDD2.n55 VDD2.n54 185
R2209 VDD2.n12 VDD2.n11 185
R2210 VDD2.n61 VDD2.n60 185
R2211 VDD2.n63 VDD2.n62 185
R2212 VDD2.n8 VDD2.n7 185
R2213 VDD2.n70 VDD2.n69 185
R2214 VDD2.n71 VDD2.n6 185
R2215 VDD2.n73 VDD2.n72 185
R2216 VDD2.n4 VDD2.n3 185
R2217 VDD2.n79 VDD2.n78 185
R2218 VDD2.n81 VDD2.n80 185
R2219 VDD2.n114 VDD2.t1 147.659
R2220 VDD2.n27 VDD2.t0 147.659
R2221 VDD2.n165 VDD2.n164 104.615
R2222 VDD2.n164 VDD2.n88 104.615
R2223 VDD2.n93 VDD2.n88 104.615
R2224 VDD2.n157 VDD2.n93 104.615
R2225 VDD2.n157 VDD2.n156 104.615
R2226 VDD2.n156 VDD2.n94 104.615
R2227 VDD2.n149 VDD2.n94 104.615
R2228 VDD2.n149 VDD2.n148 104.615
R2229 VDD2.n148 VDD2.n98 104.615
R2230 VDD2.n141 VDD2.n98 104.615
R2231 VDD2.n141 VDD2.n140 104.615
R2232 VDD2.n140 VDD2.n102 104.615
R2233 VDD2.n133 VDD2.n102 104.615
R2234 VDD2.n133 VDD2.n132 104.615
R2235 VDD2.n132 VDD2.n106 104.615
R2236 VDD2.n125 VDD2.n106 104.615
R2237 VDD2.n125 VDD2.n124 104.615
R2238 VDD2.n124 VDD2.n110 104.615
R2239 VDD2.n117 VDD2.n110 104.615
R2240 VDD2.n117 VDD2.n116 104.615
R2241 VDD2.n30 VDD2.n29 104.615
R2242 VDD2.n30 VDD2.n23 104.615
R2243 VDD2.n37 VDD2.n23 104.615
R2244 VDD2.n38 VDD2.n37 104.615
R2245 VDD2.n38 VDD2.n19 104.615
R2246 VDD2.n45 VDD2.n19 104.615
R2247 VDD2.n46 VDD2.n45 104.615
R2248 VDD2.n46 VDD2.n15 104.615
R2249 VDD2.n53 VDD2.n15 104.615
R2250 VDD2.n54 VDD2.n53 104.615
R2251 VDD2.n54 VDD2.n11 104.615
R2252 VDD2.n61 VDD2.n11 104.615
R2253 VDD2.n62 VDD2.n61 104.615
R2254 VDD2.n62 VDD2.n7 104.615
R2255 VDD2.n70 VDD2.n7 104.615
R2256 VDD2.n71 VDD2.n70 104.615
R2257 VDD2.n72 VDD2.n71 104.615
R2258 VDD2.n72 VDD2.n3 104.615
R2259 VDD2.n79 VDD2.n3 104.615
R2260 VDD2.n80 VDD2.n79 104.615
R2261 VDD2.n170 VDD2.n84 93.7645
R2262 VDD2.n116 VDD2.t1 52.3082
R2263 VDD2.n29 VDD2.t0 52.3082
R2264 VDD2.n170 VDD2.n169 51.9672
R2265 VDD2.n115 VDD2.n114 15.6677
R2266 VDD2.n28 VDD2.n27 15.6677
R2267 VDD2.n91 VDD2.n89 13.1884
R2268 VDD2.n73 VDD2.n4 13.1884
R2269 VDD2.n163 VDD2.n162 12.8005
R2270 VDD2.n159 VDD2.n158 12.8005
R2271 VDD2.n118 VDD2.n113 12.8005
R2272 VDD2.n31 VDD2.n26 12.8005
R2273 VDD2.n74 VDD2.n6 12.8005
R2274 VDD2.n78 VDD2.n77 12.8005
R2275 VDD2.n166 VDD2.n87 12.0247
R2276 VDD2.n155 VDD2.n92 12.0247
R2277 VDD2.n119 VDD2.n111 12.0247
R2278 VDD2.n32 VDD2.n24 12.0247
R2279 VDD2.n69 VDD2.n68 12.0247
R2280 VDD2.n81 VDD2.n2 12.0247
R2281 VDD2.n167 VDD2.n85 11.249
R2282 VDD2.n154 VDD2.n95 11.249
R2283 VDD2.n123 VDD2.n122 11.249
R2284 VDD2.n36 VDD2.n35 11.249
R2285 VDD2.n67 VDD2.n8 11.249
R2286 VDD2.n82 VDD2.n0 11.249
R2287 VDD2.n151 VDD2.n150 10.4732
R2288 VDD2.n126 VDD2.n109 10.4732
R2289 VDD2.n39 VDD2.n22 10.4732
R2290 VDD2.n64 VDD2.n63 10.4732
R2291 VDD2.n147 VDD2.n97 9.69747
R2292 VDD2.n127 VDD2.n107 9.69747
R2293 VDD2.n40 VDD2.n20 9.69747
R2294 VDD2.n60 VDD2.n10 9.69747
R2295 VDD2.n169 VDD2.n168 9.45567
R2296 VDD2.n84 VDD2.n83 9.45567
R2297 VDD2.n101 VDD2.n100 9.3005
R2298 VDD2.n144 VDD2.n143 9.3005
R2299 VDD2.n146 VDD2.n145 9.3005
R2300 VDD2.n97 VDD2.n96 9.3005
R2301 VDD2.n152 VDD2.n151 9.3005
R2302 VDD2.n154 VDD2.n153 9.3005
R2303 VDD2.n92 VDD2.n90 9.3005
R2304 VDD2.n160 VDD2.n159 9.3005
R2305 VDD2.n168 VDD2.n167 9.3005
R2306 VDD2.n87 VDD2.n86 9.3005
R2307 VDD2.n162 VDD2.n161 9.3005
R2308 VDD2.n138 VDD2.n137 9.3005
R2309 VDD2.n136 VDD2.n135 9.3005
R2310 VDD2.n105 VDD2.n104 9.3005
R2311 VDD2.n130 VDD2.n129 9.3005
R2312 VDD2.n128 VDD2.n127 9.3005
R2313 VDD2.n109 VDD2.n108 9.3005
R2314 VDD2.n122 VDD2.n121 9.3005
R2315 VDD2.n120 VDD2.n119 9.3005
R2316 VDD2.n113 VDD2.n112 9.3005
R2317 VDD2.n83 VDD2.n82 9.3005
R2318 VDD2.n2 VDD2.n1 9.3005
R2319 VDD2.n77 VDD2.n76 9.3005
R2320 VDD2.n49 VDD2.n48 9.3005
R2321 VDD2.n18 VDD2.n17 9.3005
R2322 VDD2.n43 VDD2.n42 9.3005
R2323 VDD2.n41 VDD2.n40 9.3005
R2324 VDD2.n22 VDD2.n21 9.3005
R2325 VDD2.n35 VDD2.n34 9.3005
R2326 VDD2.n33 VDD2.n32 9.3005
R2327 VDD2.n26 VDD2.n25 9.3005
R2328 VDD2.n51 VDD2.n50 9.3005
R2329 VDD2.n14 VDD2.n13 9.3005
R2330 VDD2.n57 VDD2.n56 9.3005
R2331 VDD2.n59 VDD2.n58 9.3005
R2332 VDD2.n10 VDD2.n9 9.3005
R2333 VDD2.n65 VDD2.n64 9.3005
R2334 VDD2.n67 VDD2.n66 9.3005
R2335 VDD2.n68 VDD2.n5 9.3005
R2336 VDD2.n75 VDD2.n74 9.3005
R2337 VDD2.n146 VDD2.n99 8.92171
R2338 VDD2.n131 VDD2.n130 8.92171
R2339 VDD2.n44 VDD2.n43 8.92171
R2340 VDD2.n59 VDD2.n12 8.92171
R2341 VDD2.n143 VDD2.n142 8.14595
R2342 VDD2.n134 VDD2.n105 8.14595
R2343 VDD2.n47 VDD2.n18 8.14595
R2344 VDD2.n56 VDD2.n55 8.14595
R2345 VDD2.n139 VDD2.n101 7.3702
R2346 VDD2.n135 VDD2.n103 7.3702
R2347 VDD2.n48 VDD2.n16 7.3702
R2348 VDD2.n52 VDD2.n14 7.3702
R2349 VDD2.n139 VDD2.n138 6.59444
R2350 VDD2.n138 VDD2.n103 6.59444
R2351 VDD2.n51 VDD2.n16 6.59444
R2352 VDD2.n52 VDD2.n51 6.59444
R2353 VDD2.n142 VDD2.n101 5.81868
R2354 VDD2.n135 VDD2.n134 5.81868
R2355 VDD2.n48 VDD2.n47 5.81868
R2356 VDD2.n55 VDD2.n14 5.81868
R2357 VDD2.n143 VDD2.n99 5.04292
R2358 VDD2.n131 VDD2.n105 5.04292
R2359 VDD2.n44 VDD2.n18 5.04292
R2360 VDD2.n56 VDD2.n12 5.04292
R2361 VDD2.n114 VDD2.n112 4.38563
R2362 VDD2.n27 VDD2.n25 4.38563
R2363 VDD2.n147 VDD2.n146 4.26717
R2364 VDD2.n130 VDD2.n107 4.26717
R2365 VDD2.n43 VDD2.n20 4.26717
R2366 VDD2.n60 VDD2.n59 4.26717
R2367 VDD2.n150 VDD2.n97 3.49141
R2368 VDD2.n127 VDD2.n126 3.49141
R2369 VDD2.n40 VDD2.n39 3.49141
R2370 VDD2.n63 VDD2.n10 3.49141
R2371 VDD2.n169 VDD2.n85 2.71565
R2372 VDD2.n151 VDD2.n95 2.71565
R2373 VDD2.n123 VDD2.n109 2.71565
R2374 VDD2.n36 VDD2.n22 2.71565
R2375 VDD2.n64 VDD2.n8 2.71565
R2376 VDD2.n84 VDD2.n0 2.71565
R2377 VDD2.n167 VDD2.n166 1.93989
R2378 VDD2.n155 VDD2.n154 1.93989
R2379 VDD2.n122 VDD2.n111 1.93989
R2380 VDD2.n35 VDD2.n24 1.93989
R2381 VDD2.n69 VDD2.n67 1.93989
R2382 VDD2.n82 VDD2.n81 1.93989
R2383 VDD2.n163 VDD2.n87 1.16414
R2384 VDD2.n158 VDD2.n92 1.16414
R2385 VDD2.n119 VDD2.n118 1.16414
R2386 VDD2.n32 VDD2.n31 1.16414
R2387 VDD2.n68 VDD2.n6 1.16414
R2388 VDD2.n78 VDD2.n2 1.16414
R2389 VDD2 VDD2.n170 0.653517
R2390 VDD2.n162 VDD2.n89 0.388379
R2391 VDD2.n159 VDD2.n91 0.388379
R2392 VDD2.n115 VDD2.n113 0.388379
R2393 VDD2.n28 VDD2.n26 0.388379
R2394 VDD2.n74 VDD2.n73 0.388379
R2395 VDD2.n77 VDD2.n4 0.388379
R2396 VDD2.n168 VDD2.n86 0.155672
R2397 VDD2.n161 VDD2.n86 0.155672
R2398 VDD2.n161 VDD2.n160 0.155672
R2399 VDD2.n160 VDD2.n90 0.155672
R2400 VDD2.n153 VDD2.n90 0.155672
R2401 VDD2.n153 VDD2.n152 0.155672
R2402 VDD2.n152 VDD2.n96 0.155672
R2403 VDD2.n145 VDD2.n96 0.155672
R2404 VDD2.n145 VDD2.n144 0.155672
R2405 VDD2.n144 VDD2.n100 0.155672
R2406 VDD2.n137 VDD2.n100 0.155672
R2407 VDD2.n137 VDD2.n136 0.155672
R2408 VDD2.n136 VDD2.n104 0.155672
R2409 VDD2.n129 VDD2.n104 0.155672
R2410 VDD2.n129 VDD2.n128 0.155672
R2411 VDD2.n128 VDD2.n108 0.155672
R2412 VDD2.n121 VDD2.n108 0.155672
R2413 VDD2.n121 VDD2.n120 0.155672
R2414 VDD2.n120 VDD2.n112 0.155672
R2415 VDD2.n33 VDD2.n25 0.155672
R2416 VDD2.n34 VDD2.n33 0.155672
R2417 VDD2.n34 VDD2.n21 0.155672
R2418 VDD2.n41 VDD2.n21 0.155672
R2419 VDD2.n42 VDD2.n41 0.155672
R2420 VDD2.n42 VDD2.n17 0.155672
R2421 VDD2.n49 VDD2.n17 0.155672
R2422 VDD2.n50 VDD2.n49 0.155672
R2423 VDD2.n50 VDD2.n13 0.155672
R2424 VDD2.n57 VDD2.n13 0.155672
R2425 VDD2.n58 VDD2.n57 0.155672
R2426 VDD2.n58 VDD2.n9 0.155672
R2427 VDD2.n65 VDD2.n9 0.155672
R2428 VDD2.n66 VDD2.n65 0.155672
R2429 VDD2.n66 VDD2.n5 0.155672
R2430 VDD2.n75 VDD2.n5 0.155672
R2431 VDD2.n76 VDD2.n75 0.155672
R2432 VDD2.n76 VDD2.n1 0.155672
R2433 VDD2.n83 VDD2.n1 0.155672
C0 VTAIL VDD2 6.03493f
C1 VN VDD1 0.148378f
C2 VTAIL VP 2.99105f
C3 VTAIL VDD1 5.98652f
C4 VN VTAIL 2.9767f
C5 VDD2 VP 0.326562f
C6 VDD1 VDD2 0.654694f
C7 VDD1 VP 3.65954f
C8 VN VDD2 3.48463f
C9 VN VP 6.02403f
C10 VDD2 B 5.002263f
C11 VDD1 B 7.99917f
C12 VTAIL B 8.715515f
C13 VN B 11.36827f
C14 VP B 6.423227f
C15 VDD2.n0 B 0.02809f
C16 VDD2.n1 B 0.019984f
C17 VDD2.n2 B 0.010739f
C18 VDD2.n3 B 0.025383f
C19 VDD2.n4 B 0.011055f
C20 VDD2.n5 B 0.019984f
C21 VDD2.n6 B 0.01137f
C22 VDD2.n7 B 0.025383f
C23 VDD2.n8 B 0.01137f
C24 VDD2.n9 B 0.019984f
C25 VDD2.n10 B 0.010739f
C26 VDD2.n11 B 0.025383f
C27 VDD2.n12 B 0.01137f
C28 VDD2.n13 B 0.019984f
C29 VDD2.n14 B 0.010739f
C30 VDD2.n15 B 0.025383f
C31 VDD2.n16 B 0.01137f
C32 VDD2.n17 B 0.019984f
C33 VDD2.n18 B 0.010739f
C34 VDD2.n19 B 0.025383f
C35 VDD2.n20 B 0.01137f
C36 VDD2.n21 B 0.019984f
C37 VDD2.n22 B 0.010739f
C38 VDD2.n23 B 0.025383f
C39 VDD2.n24 B 0.01137f
C40 VDD2.n25 B 1.34784f
C41 VDD2.n26 B 0.010739f
C42 VDD2.t0 B 0.041888f
C43 VDD2.n27 B 0.132948f
C44 VDD2.n28 B 0.014994f
C45 VDD2.n29 B 0.019037f
C46 VDD2.n30 B 0.025383f
C47 VDD2.n31 B 0.01137f
C48 VDD2.n32 B 0.010739f
C49 VDD2.n33 B 0.019984f
C50 VDD2.n34 B 0.019984f
C51 VDD2.n35 B 0.010739f
C52 VDD2.n36 B 0.01137f
C53 VDD2.n37 B 0.025383f
C54 VDD2.n38 B 0.025383f
C55 VDD2.n39 B 0.01137f
C56 VDD2.n40 B 0.010739f
C57 VDD2.n41 B 0.019984f
C58 VDD2.n42 B 0.019984f
C59 VDD2.n43 B 0.010739f
C60 VDD2.n44 B 0.01137f
C61 VDD2.n45 B 0.025383f
C62 VDD2.n46 B 0.025383f
C63 VDD2.n47 B 0.01137f
C64 VDD2.n48 B 0.010739f
C65 VDD2.n49 B 0.019984f
C66 VDD2.n50 B 0.019984f
C67 VDD2.n51 B 0.010739f
C68 VDD2.n52 B 0.01137f
C69 VDD2.n53 B 0.025383f
C70 VDD2.n54 B 0.025383f
C71 VDD2.n55 B 0.01137f
C72 VDD2.n56 B 0.010739f
C73 VDD2.n57 B 0.019984f
C74 VDD2.n58 B 0.019984f
C75 VDD2.n59 B 0.010739f
C76 VDD2.n60 B 0.01137f
C77 VDD2.n61 B 0.025383f
C78 VDD2.n62 B 0.025383f
C79 VDD2.n63 B 0.01137f
C80 VDD2.n64 B 0.010739f
C81 VDD2.n65 B 0.019984f
C82 VDD2.n66 B 0.019984f
C83 VDD2.n67 B 0.010739f
C84 VDD2.n68 B 0.010739f
C85 VDD2.n69 B 0.01137f
C86 VDD2.n70 B 0.025383f
C87 VDD2.n71 B 0.025383f
C88 VDD2.n72 B 0.025383f
C89 VDD2.n73 B 0.011055f
C90 VDD2.n74 B 0.010739f
C91 VDD2.n75 B 0.019984f
C92 VDD2.n76 B 0.019984f
C93 VDD2.n77 B 0.010739f
C94 VDD2.n78 B 0.01137f
C95 VDD2.n79 B 0.025383f
C96 VDD2.n80 B 0.054949f
C97 VDD2.n81 B 0.01137f
C98 VDD2.n82 B 0.010739f
C99 VDD2.n83 B 0.050561f
C100 VDD2.n84 B 0.661309f
C101 VDD2.n85 B 0.02809f
C102 VDD2.n86 B 0.019984f
C103 VDD2.n87 B 0.010739f
C104 VDD2.n88 B 0.025383f
C105 VDD2.n89 B 0.011055f
C106 VDD2.n90 B 0.019984f
C107 VDD2.n91 B 0.011055f
C108 VDD2.n92 B 0.010739f
C109 VDD2.n93 B 0.025383f
C110 VDD2.n94 B 0.025383f
C111 VDD2.n95 B 0.01137f
C112 VDD2.n96 B 0.019984f
C113 VDD2.n97 B 0.010739f
C114 VDD2.n98 B 0.025383f
C115 VDD2.n99 B 0.01137f
C116 VDD2.n100 B 0.019984f
C117 VDD2.n101 B 0.010739f
C118 VDD2.n102 B 0.025383f
C119 VDD2.n103 B 0.01137f
C120 VDD2.n104 B 0.019984f
C121 VDD2.n105 B 0.010739f
C122 VDD2.n106 B 0.025383f
C123 VDD2.n107 B 0.01137f
C124 VDD2.n108 B 0.019984f
C125 VDD2.n109 B 0.010739f
C126 VDD2.n110 B 0.025383f
C127 VDD2.n111 B 0.01137f
C128 VDD2.n112 B 1.34784f
C129 VDD2.n113 B 0.010739f
C130 VDD2.t1 B 0.041888f
C131 VDD2.n114 B 0.132948f
C132 VDD2.n115 B 0.014994f
C133 VDD2.n116 B 0.019037f
C134 VDD2.n117 B 0.025383f
C135 VDD2.n118 B 0.01137f
C136 VDD2.n119 B 0.010739f
C137 VDD2.n120 B 0.019984f
C138 VDD2.n121 B 0.019984f
C139 VDD2.n122 B 0.010739f
C140 VDD2.n123 B 0.01137f
C141 VDD2.n124 B 0.025383f
C142 VDD2.n125 B 0.025383f
C143 VDD2.n126 B 0.01137f
C144 VDD2.n127 B 0.010739f
C145 VDD2.n128 B 0.019984f
C146 VDD2.n129 B 0.019984f
C147 VDD2.n130 B 0.010739f
C148 VDD2.n131 B 0.01137f
C149 VDD2.n132 B 0.025383f
C150 VDD2.n133 B 0.025383f
C151 VDD2.n134 B 0.01137f
C152 VDD2.n135 B 0.010739f
C153 VDD2.n136 B 0.019984f
C154 VDD2.n137 B 0.019984f
C155 VDD2.n138 B 0.010739f
C156 VDD2.n139 B 0.01137f
C157 VDD2.n140 B 0.025383f
C158 VDD2.n141 B 0.025383f
C159 VDD2.n142 B 0.01137f
C160 VDD2.n143 B 0.010739f
C161 VDD2.n144 B 0.019984f
C162 VDD2.n145 B 0.019984f
C163 VDD2.n146 B 0.010739f
C164 VDD2.n147 B 0.01137f
C165 VDD2.n148 B 0.025383f
C166 VDD2.n149 B 0.025383f
C167 VDD2.n150 B 0.01137f
C168 VDD2.n151 B 0.010739f
C169 VDD2.n152 B 0.019984f
C170 VDD2.n153 B 0.019984f
C171 VDD2.n154 B 0.010739f
C172 VDD2.n155 B 0.01137f
C173 VDD2.n156 B 0.025383f
C174 VDD2.n157 B 0.025383f
C175 VDD2.n158 B 0.01137f
C176 VDD2.n159 B 0.010739f
C177 VDD2.n160 B 0.019984f
C178 VDD2.n161 B 0.019984f
C179 VDD2.n162 B 0.010739f
C180 VDD2.n163 B 0.01137f
C181 VDD2.n164 B 0.025383f
C182 VDD2.n165 B 0.054949f
C183 VDD2.n166 B 0.01137f
C184 VDD2.n167 B 0.010739f
C185 VDD2.n168 B 0.050561f
C186 VDD2.n169 B 0.044643f
C187 VDD2.n170 B 2.72715f
C188 VN.t1 B 3.55063f
C189 VN.t0 B 4.05168f
C190 VDD1.n0 B 0.02846f
C191 VDD1.n1 B 0.020248f
C192 VDD1.n2 B 0.01088f
C193 VDD1.n3 B 0.025717f
C194 VDD1.n4 B 0.0112f
C195 VDD1.n5 B 0.020248f
C196 VDD1.n6 B 0.0112f
C197 VDD1.n7 B 0.01088f
C198 VDD1.n8 B 0.025717f
C199 VDD1.n9 B 0.025717f
C200 VDD1.n10 B 0.01152f
C201 VDD1.n11 B 0.020248f
C202 VDD1.n12 B 0.01088f
C203 VDD1.n13 B 0.025717f
C204 VDD1.n14 B 0.01152f
C205 VDD1.n15 B 0.020248f
C206 VDD1.n16 B 0.01088f
C207 VDD1.n17 B 0.025717f
C208 VDD1.n18 B 0.01152f
C209 VDD1.n19 B 0.020248f
C210 VDD1.n20 B 0.01088f
C211 VDD1.n21 B 0.025717f
C212 VDD1.n22 B 0.01152f
C213 VDD1.n23 B 0.020248f
C214 VDD1.n24 B 0.01088f
C215 VDD1.n25 B 0.025717f
C216 VDD1.n26 B 0.01152f
C217 VDD1.n27 B 1.3656f
C218 VDD1.n28 B 0.01088f
C219 VDD1.t0 B 0.04244f
C220 VDD1.n29 B 0.1347f
C221 VDD1.n30 B 0.015192f
C222 VDD1.n31 B 0.019288f
C223 VDD1.n32 B 0.025717f
C224 VDD1.n33 B 0.01152f
C225 VDD1.n34 B 0.01088f
C226 VDD1.n35 B 0.020248f
C227 VDD1.n36 B 0.020248f
C228 VDD1.n37 B 0.01088f
C229 VDD1.n38 B 0.01152f
C230 VDD1.n39 B 0.025717f
C231 VDD1.n40 B 0.025717f
C232 VDD1.n41 B 0.01152f
C233 VDD1.n42 B 0.01088f
C234 VDD1.n43 B 0.020248f
C235 VDD1.n44 B 0.020248f
C236 VDD1.n45 B 0.01088f
C237 VDD1.n46 B 0.01152f
C238 VDD1.n47 B 0.025717f
C239 VDD1.n48 B 0.025717f
C240 VDD1.n49 B 0.01152f
C241 VDD1.n50 B 0.01088f
C242 VDD1.n51 B 0.020248f
C243 VDD1.n52 B 0.020248f
C244 VDD1.n53 B 0.01088f
C245 VDD1.n54 B 0.01152f
C246 VDD1.n55 B 0.025717f
C247 VDD1.n56 B 0.025717f
C248 VDD1.n57 B 0.01152f
C249 VDD1.n58 B 0.01088f
C250 VDD1.n59 B 0.020248f
C251 VDD1.n60 B 0.020248f
C252 VDD1.n61 B 0.01088f
C253 VDD1.n62 B 0.01152f
C254 VDD1.n63 B 0.025717f
C255 VDD1.n64 B 0.025717f
C256 VDD1.n65 B 0.01152f
C257 VDD1.n66 B 0.01088f
C258 VDD1.n67 B 0.020248f
C259 VDD1.n68 B 0.020248f
C260 VDD1.n69 B 0.01088f
C261 VDD1.n70 B 0.01152f
C262 VDD1.n71 B 0.025717f
C263 VDD1.n72 B 0.025717f
C264 VDD1.n73 B 0.01152f
C265 VDD1.n74 B 0.01088f
C266 VDD1.n75 B 0.020248f
C267 VDD1.n76 B 0.020248f
C268 VDD1.n77 B 0.01088f
C269 VDD1.n78 B 0.01152f
C270 VDD1.n79 B 0.025717f
C271 VDD1.n80 B 0.055673f
C272 VDD1.n81 B 0.01152f
C273 VDD1.n82 B 0.01088f
C274 VDD1.n83 B 0.051227f
C275 VDD1.n84 B 0.046275f
C276 VDD1.n85 B 0.02846f
C277 VDD1.n86 B 0.020248f
C278 VDD1.n87 B 0.01088f
C279 VDD1.n88 B 0.025717f
C280 VDD1.n89 B 0.0112f
C281 VDD1.n90 B 0.020248f
C282 VDD1.n91 B 0.01152f
C283 VDD1.n92 B 0.025717f
C284 VDD1.n93 B 0.01152f
C285 VDD1.n94 B 0.020248f
C286 VDD1.n95 B 0.01088f
C287 VDD1.n96 B 0.025717f
C288 VDD1.n97 B 0.01152f
C289 VDD1.n98 B 0.020248f
C290 VDD1.n99 B 0.01088f
C291 VDD1.n100 B 0.025717f
C292 VDD1.n101 B 0.01152f
C293 VDD1.n102 B 0.020248f
C294 VDD1.n103 B 0.01088f
C295 VDD1.n104 B 0.025717f
C296 VDD1.n105 B 0.01152f
C297 VDD1.n106 B 0.020248f
C298 VDD1.n107 B 0.01088f
C299 VDD1.n108 B 0.025717f
C300 VDD1.n109 B 0.01152f
C301 VDD1.n110 B 1.3656f
C302 VDD1.n111 B 0.01088f
C303 VDD1.t1 B 0.04244f
C304 VDD1.n112 B 0.1347f
C305 VDD1.n113 B 0.015192f
C306 VDD1.n114 B 0.019288f
C307 VDD1.n115 B 0.025717f
C308 VDD1.n116 B 0.01152f
C309 VDD1.n117 B 0.01088f
C310 VDD1.n118 B 0.020248f
C311 VDD1.n119 B 0.020248f
C312 VDD1.n120 B 0.01088f
C313 VDD1.n121 B 0.01152f
C314 VDD1.n122 B 0.025717f
C315 VDD1.n123 B 0.025717f
C316 VDD1.n124 B 0.01152f
C317 VDD1.n125 B 0.01088f
C318 VDD1.n126 B 0.020248f
C319 VDD1.n127 B 0.020248f
C320 VDD1.n128 B 0.01088f
C321 VDD1.n129 B 0.01152f
C322 VDD1.n130 B 0.025717f
C323 VDD1.n131 B 0.025717f
C324 VDD1.n132 B 0.01152f
C325 VDD1.n133 B 0.01088f
C326 VDD1.n134 B 0.020248f
C327 VDD1.n135 B 0.020248f
C328 VDD1.n136 B 0.01088f
C329 VDD1.n137 B 0.01152f
C330 VDD1.n138 B 0.025717f
C331 VDD1.n139 B 0.025717f
C332 VDD1.n140 B 0.01152f
C333 VDD1.n141 B 0.01088f
C334 VDD1.n142 B 0.020248f
C335 VDD1.n143 B 0.020248f
C336 VDD1.n144 B 0.01088f
C337 VDD1.n145 B 0.01152f
C338 VDD1.n146 B 0.025717f
C339 VDD1.n147 B 0.025717f
C340 VDD1.n148 B 0.01152f
C341 VDD1.n149 B 0.01088f
C342 VDD1.n150 B 0.020248f
C343 VDD1.n151 B 0.020248f
C344 VDD1.n152 B 0.01088f
C345 VDD1.n153 B 0.01088f
C346 VDD1.n154 B 0.01152f
C347 VDD1.n155 B 0.025717f
C348 VDD1.n156 B 0.025717f
C349 VDD1.n157 B 0.025717f
C350 VDD1.n158 B 0.0112f
C351 VDD1.n159 B 0.01088f
C352 VDD1.n160 B 0.020248f
C353 VDD1.n161 B 0.020248f
C354 VDD1.n162 B 0.01088f
C355 VDD1.n163 B 0.01152f
C356 VDD1.n164 B 0.025717f
C357 VDD1.n165 B 0.055673f
C358 VDD1.n166 B 0.01152f
C359 VDD1.n167 B 0.01088f
C360 VDD1.n168 B 0.051227f
C361 VDD1.n169 B 0.709735f
C362 VTAIL.n0 B 0.028128f
C363 VTAIL.n1 B 0.020011f
C364 VTAIL.n2 B 0.010753f
C365 VTAIL.n3 B 0.025417f
C366 VTAIL.n4 B 0.011069f
C367 VTAIL.n5 B 0.020011f
C368 VTAIL.n6 B 0.011386f
C369 VTAIL.n7 B 0.025417f
C370 VTAIL.n8 B 0.011386f
C371 VTAIL.n9 B 0.020011f
C372 VTAIL.n10 B 0.010753f
C373 VTAIL.n11 B 0.025417f
C374 VTAIL.n12 B 0.011386f
C375 VTAIL.n13 B 0.020011f
C376 VTAIL.n14 B 0.010753f
C377 VTAIL.n15 B 0.025417f
C378 VTAIL.n16 B 0.011386f
C379 VTAIL.n17 B 0.020011f
C380 VTAIL.n18 B 0.010753f
C381 VTAIL.n19 B 0.025417f
C382 VTAIL.n20 B 0.011386f
C383 VTAIL.n21 B 0.020011f
C384 VTAIL.n22 B 0.010753f
C385 VTAIL.n23 B 0.025417f
C386 VTAIL.n24 B 0.011386f
C387 VTAIL.n25 B 1.34965f
C388 VTAIL.n26 B 0.010753f
C389 VTAIL.t2 B 0.041945f
C390 VTAIL.n27 B 0.133127f
C391 VTAIL.n28 B 0.015014f
C392 VTAIL.n29 B 0.019063f
C393 VTAIL.n30 B 0.025417f
C394 VTAIL.n31 B 0.011386f
C395 VTAIL.n32 B 0.010753f
C396 VTAIL.n33 B 0.020011f
C397 VTAIL.n34 B 0.020011f
C398 VTAIL.n35 B 0.010753f
C399 VTAIL.n36 B 0.011386f
C400 VTAIL.n37 B 0.025417f
C401 VTAIL.n38 B 0.025417f
C402 VTAIL.n39 B 0.011386f
C403 VTAIL.n40 B 0.010753f
C404 VTAIL.n41 B 0.020011f
C405 VTAIL.n42 B 0.020011f
C406 VTAIL.n43 B 0.010753f
C407 VTAIL.n44 B 0.011386f
C408 VTAIL.n45 B 0.025417f
C409 VTAIL.n46 B 0.025417f
C410 VTAIL.n47 B 0.011386f
C411 VTAIL.n48 B 0.010753f
C412 VTAIL.n49 B 0.020011f
C413 VTAIL.n50 B 0.020011f
C414 VTAIL.n51 B 0.010753f
C415 VTAIL.n52 B 0.011386f
C416 VTAIL.n53 B 0.025417f
C417 VTAIL.n54 B 0.025417f
C418 VTAIL.n55 B 0.011386f
C419 VTAIL.n56 B 0.010753f
C420 VTAIL.n57 B 0.020011f
C421 VTAIL.n58 B 0.020011f
C422 VTAIL.n59 B 0.010753f
C423 VTAIL.n60 B 0.011386f
C424 VTAIL.n61 B 0.025417f
C425 VTAIL.n62 B 0.025417f
C426 VTAIL.n63 B 0.011386f
C427 VTAIL.n64 B 0.010753f
C428 VTAIL.n65 B 0.020011f
C429 VTAIL.n66 B 0.020011f
C430 VTAIL.n67 B 0.010753f
C431 VTAIL.n68 B 0.010753f
C432 VTAIL.n69 B 0.011386f
C433 VTAIL.n70 B 0.025417f
C434 VTAIL.n71 B 0.025417f
C435 VTAIL.n72 B 0.025417f
C436 VTAIL.n73 B 0.011069f
C437 VTAIL.n74 B 0.010753f
C438 VTAIL.n75 B 0.020011f
C439 VTAIL.n76 B 0.020011f
C440 VTAIL.n77 B 0.010753f
C441 VTAIL.n78 B 0.011386f
C442 VTAIL.n79 B 0.025417f
C443 VTAIL.n80 B 0.055023f
C444 VTAIL.n81 B 0.011386f
C445 VTAIL.n82 B 0.010753f
C446 VTAIL.n83 B 0.050629f
C447 VTAIL.n84 B 0.030916f
C448 VTAIL.n85 B 1.53334f
C449 VTAIL.n86 B 0.028128f
C450 VTAIL.n87 B 0.020011f
C451 VTAIL.n88 B 0.010753f
C452 VTAIL.n89 B 0.025417f
C453 VTAIL.n90 B 0.011069f
C454 VTAIL.n91 B 0.020011f
C455 VTAIL.n92 B 0.011069f
C456 VTAIL.n93 B 0.010753f
C457 VTAIL.n94 B 0.025417f
C458 VTAIL.n95 B 0.025417f
C459 VTAIL.n96 B 0.011386f
C460 VTAIL.n97 B 0.020011f
C461 VTAIL.n98 B 0.010753f
C462 VTAIL.n99 B 0.025417f
C463 VTAIL.n100 B 0.011386f
C464 VTAIL.n101 B 0.020011f
C465 VTAIL.n102 B 0.010753f
C466 VTAIL.n103 B 0.025417f
C467 VTAIL.n104 B 0.011386f
C468 VTAIL.n105 B 0.020011f
C469 VTAIL.n106 B 0.010753f
C470 VTAIL.n107 B 0.025417f
C471 VTAIL.n108 B 0.011386f
C472 VTAIL.n109 B 0.020011f
C473 VTAIL.n110 B 0.010753f
C474 VTAIL.n111 B 0.025417f
C475 VTAIL.n112 B 0.011386f
C476 VTAIL.n113 B 1.34965f
C477 VTAIL.n114 B 0.010753f
C478 VTAIL.t1 B 0.041945f
C479 VTAIL.n115 B 0.133127f
C480 VTAIL.n116 B 0.015014f
C481 VTAIL.n117 B 0.019063f
C482 VTAIL.n118 B 0.025417f
C483 VTAIL.n119 B 0.011386f
C484 VTAIL.n120 B 0.010753f
C485 VTAIL.n121 B 0.020011f
C486 VTAIL.n122 B 0.020011f
C487 VTAIL.n123 B 0.010753f
C488 VTAIL.n124 B 0.011386f
C489 VTAIL.n125 B 0.025417f
C490 VTAIL.n126 B 0.025417f
C491 VTAIL.n127 B 0.011386f
C492 VTAIL.n128 B 0.010753f
C493 VTAIL.n129 B 0.020011f
C494 VTAIL.n130 B 0.020011f
C495 VTAIL.n131 B 0.010753f
C496 VTAIL.n132 B 0.011386f
C497 VTAIL.n133 B 0.025417f
C498 VTAIL.n134 B 0.025417f
C499 VTAIL.n135 B 0.011386f
C500 VTAIL.n136 B 0.010753f
C501 VTAIL.n137 B 0.020011f
C502 VTAIL.n138 B 0.020011f
C503 VTAIL.n139 B 0.010753f
C504 VTAIL.n140 B 0.011386f
C505 VTAIL.n141 B 0.025417f
C506 VTAIL.n142 B 0.025417f
C507 VTAIL.n143 B 0.011386f
C508 VTAIL.n144 B 0.010753f
C509 VTAIL.n145 B 0.020011f
C510 VTAIL.n146 B 0.020011f
C511 VTAIL.n147 B 0.010753f
C512 VTAIL.n148 B 0.011386f
C513 VTAIL.n149 B 0.025417f
C514 VTAIL.n150 B 0.025417f
C515 VTAIL.n151 B 0.011386f
C516 VTAIL.n152 B 0.010753f
C517 VTAIL.n153 B 0.020011f
C518 VTAIL.n154 B 0.020011f
C519 VTAIL.n155 B 0.010753f
C520 VTAIL.n156 B 0.011386f
C521 VTAIL.n157 B 0.025417f
C522 VTAIL.n158 B 0.025417f
C523 VTAIL.n159 B 0.011386f
C524 VTAIL.n160 B 0.010753f
C525 VTAIL.n161 B 0.020011f
C526 VTAIL.n162 B 0.020011f
C527 VTAIL.n163 B 0.010753f
C528 VTAIL.n164 B 0.011386f
C529 VTAIL.n165 B 0.025417f
C530 VTAIL.n166 B 0.055023f
C531 VTAIL.n167 B 0.011386f
C532 VTAIL.n168 B 0.010753f
C533 VTAIL.n169 B 0.050629f
C534 VTAIL.n170 B 0.030916f
C535 VTAIL.n171 B 1.56795f
C536 VTAIL.n172 B 0.028128f
C537 VTAIL.n173 B 0.020011f
C538 VTAIL.n174 B 0.010753f
C539 VTAIL.n175 B 0.025417f
C540 VTAIL.n176 B 0.011069f
C541 VTAIL.n177 B 0.020011f
C542 VTAIL.n178 B 0.011069f
C543 VTAIL.n179 B 0.010753f
C544 VTAIL.n180 B 0.025417f
C545 VTAIL.n181 B 0.025417f
C546 VTAIL.n182 B 0.011386f
C547 VTAIL.n183 B 0.020011f
C548 VTAIL.n184 B 0.010753f
C549 VTAIL.n185 B 0.025417f
C550 VTAIL.n186 B 0.011386f
C551 VTAIL.n187 B 0.020011f
C552 VTAIL.n188 B 0.010753f
C553 VTAIL.n189 B 0.025417f
C554 VTAIL.n190 B 0.011386f
C555 VTAIL.n191 B 0.020011f
C556 VTAIL.n192 B 0.010753f
C557 VTAIL.n193 B 0.025417f
C558 VTAIL.n194 B 0.011386f
C559 VTAIL.n195 B 0.020011f
C560 VTAIL.n196 B 0.010753f
C561 VTAIL.n197 B 0.025417f
C562 VTAIL.n198 B 0.011386f
C563 VTAIL.n199 B 1.34965f
C564 VTAIL.n200 B 0.010753f
C565 VTAIL.t3 B 0.041945f
C566 VTAIL.n201 B 0.133127f
C567 VTAIL.n202 B 0.015014f
C568 VTAIL.n203 B 0.019063f
C569 VTAIL.n204 B 0.025417f
C570 VTAIL.n205 B 0.011386f
C571 VTAIL.n206 B 0.010753f
C572 VTAIL.n207 B 0.020011f
C573 VTAIL.n208 B 0.020011f
C574 VTAIL.n209 B 0.010753f
C575 VTAIL.n210 B 0.011386f
C576 VTAIL.n211 B 0.025417f
C577 VTAIL.n212 B 0.025417f
C578 VTAIL.n213 B 0.011386f
C579 VTAIL.n214 B 0.010753f
C580 VTAIL.n215 B 0.020011f
C581 VTAIL.n216 B 0.020011f
C582 VTAIL.n217 B 0.010753f
C583 VTAIL.n218 B 0.011386f
C584 VTAIL.n219 B 0.025417f
C585 VTAIL.n220 B 0.025417f
C586 VTAIL.n221 B 0.011386f
C587 VTAIL.n222 B 0.010753f
C588 VTAIL.n223 B 0.020011f
C589 VTAIL.n224 B 0.020011f
C590 VTAIL.n225 B 0.010753f
C591 VTAIL.n226 B 0.011386f
C592 VTAIL.n227 B 0.025417f
C593 VTAIL.n228 B 0.025417f
C594 VTAIL.n229 B 0.011386f
C595 VTAIL.n230 B 0.010753f
C596 VTAIL.n231 B 0.020011f
C597 VTAIL.n232 B 0.020011f
C598 VTAIL.n233 B 0.010753f
C599 VTAIL.n234 B 0.011386f
C600 VTAIL.n235 B 0.025417f
C601 VTAIL.n236 B 0.025417f
C602 VTAIL.n237 B 0.011386f
C603 VTAIL.n238 B 0.010753f
C604 VTAIL.n239 B 0.020011f
C605 VTAIL.n240 B 0.020011f
C606 VTAIL.n241 B 0.010753f
C607 VTAIL.n242 B 0.011386f
C608 VTAIL.n243 B 0.025417f
C609 VTAIL.n244 B 0.025417f
C610 VTAIL.n245 B 0.011386f
C611 VTAIL.n246 B 0.010753f
C612 VTAIL.n247 B 0.020011f
C613 VTAIL.n248 B 0.020011f
C614 VTAIL.n249 B 0.010753f
C615 VTAIL.n250 B 0.011386f
C616 VTAIL.n251 B 0.025417f
C617 VTAIL.n252 B 0.055023f
C618 VTAIL.n253 B 0.011386f
C619 VTAIL.n254 B 0.010753f
C620 VTAIL.n255 B 0.050629f
C621 VTAIL.n256 B 0.030916f
C622 VTAIL.n257 B 1.41453f
C623 VTAIL.n258 B 0.028128f
C624 VTAIL.n259 B 0.020011f
C625 VTAIL.n260 B 0.010753f
C626 VTAIL.n261 B 0.025417f
C627 VTAIL.n262 B 0.011069f
C628 VTAIL.n263 B 0.020011f
C629 VTAIL.n264 B 0.011386f
C630 VTAIL.n265 B 0.025417f
C631 VTAIL.n266 B 0.011386f
C632 VTAIL.n267 B 0.020011f
C633 VTAIL.n268 B 0.010753f
C634 VTAIL.n269 B 0.025417f
C635 VTAIL.n270 B 0.011386f
C636 VTAIL.n271 B 0.020011f
C637 VTAIL.n272 B 0.010753f
C638 VTAIL.n273 B 0.025417f
C639 VTAIL.n274 B 0.011386f
C640 VTAIL.n275 B 0.020011f
C641 VTAIL.n276 B 0.010753f
C642 VTAIL.n277 B 0.025417f
C643 VTAIL.n278 B 0.011386f
C644 VTAIL.n279 B 0.020011f
C645 VTAIL.n280 B 0.010753f
C646 VTAIL.n281 B 0.025417f
C647 VTAIL.n282 B 0.011386f
C648 VTAIL.n283 B 1.34965f
C649 VTAIL.n284 B 0.010753f
C650 VTAIL.t0 B 0.041945f
C651 VTAIL.n285 B 0.133127f
C652 VTAIL.n286 B 0.015014f
C653 VTAIL.n287 B 0.019063f
C654 VTAIL.n288 B 0.025417f
C655 VTAIL.n289 B 0.011386f
C656 VTAIL.n290 B 0.010753f
C657 VTAIL.n291 B 0.020011f
C658 VTAIL.n292 B 0.020011f
C659 VTAIL.n293 B 0.010753f
C660 VTAIL.n294 B 0.011386f
C661 VTAIL.n295 B 0.025417f
C662 VTAIL.n296 B 0.025417f
C663 VTAIL.n297 B 0.011386f
C664 VTAIL.n298 B 0.010753f
C665 VTAIL.n299 B 0.020011f
C666 VTAIL.n300 B 0.020011f
C667 VTAIL.n301 B 0.010753f
C668 VTAIL.n302 B 0.011386f
C669 VTAIL.n303 B 0.025417f
C670 VTAIL.n304 B 0.025417f
C671 VTAIL.n305 B 0.011386f
C672 VTAIL.n306 B 0.010753f
C673 VTAIL.n307 B 0.020011f
C674 VTAIL.n308 B 0.020011f
C675 VTAIL.n309 B 0.010753f
C676 VTAIL.n310 B 0.011386f
C677 VTAIL.n311 B 0.025417f
C678 VTAIL.n312 B 0.025417f
C679 VTAIL.n313 B 0.011386f
C680 VTAIL.n314 B 0.010753f
C681 VTAIL.n315 B 0.020011f
C682 VTAIL.n316 B 0.020011f
C683 VTAIL.n317 B 0.010753f
C684 VTAIL.n318 B 0.011386f
C685 VTAIL.n319 B 0.025417f
C686 VTAIL.n320 B 0.025417f
C687 VTAIL.n321 B 0.011386f
C688 VTAIL.n322 B 0.010753f
C689 VTAIL.n323 B 0.020011f
C690 VTAIL.n324 B 0.020011f
C691 VTAIL.n325 B 0.010753f
C692 VTAIL.n326 B 0.010753f
C693 VTAIL.n327 B 0.011386f
C694 VTAIL.n328 B 0.025417f
C695 VTAIL.n329 B 0.025417f
C696 VTAIL.n330 B 0.025417f
C697 VTAIL.n331 B 0.011069f
C698 VTAIL.n332 B 0.010753f
C699 VTAIL.n333 B 0.020011f
C700 VTAIL.n334 B 0.020011f
C701 VTAIL.n335 B 0.010753f
C702 VTAIL.n336 B 0.011386f
C703 VTAIL.n337 B 0.025417f
C704 VTAIL.n338 B 0.055023f
C705 VTAIL.n339 B 0.011386f
C706 VTAIL.n340 B 0.010753f
C707 VTAIL.n341 B 0.050629f
C708 VTAIL.n342 B 0.030916f
C709 VTAIL.n343 B 1.34213f
C710 VP.t1 B 4.12811f
C711 VP.t0 B 3.61824f
C712 VP.n0 B 4.88241f
.ends

