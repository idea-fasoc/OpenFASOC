* NGSPICE file created from diff_pair_sample_0018.ext - technology: sky130A

.subckt diff_pair_sample_0018 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X1 VTAIL.t16 VP.t1 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X2 VDD2.t9 VN.t0 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=2.83635 ps=17.52 w=17.19 l=2.69
X3 VDD1.t7 VP.t2 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=2.83635 ps=17.52 w=17.19 l=2.69
X4 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=0 ps=0 w=17.19 l=2.69
X5 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=0 ps=0 w=17.19 l=2.69
X6 VDD1.t6 VP.t3 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X7 VTAIL.t5 VN.t1 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X8 VDD2.t7 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=2.83635 ps=17.52 w=17.19 l=2.69
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=0 ps=0 w=17.19 l=2.69
X10 VTAIL.t1 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X11 VTAIL.t13 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X12 VDD2.t5 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X13 VTAIL.t0 VN.t5 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X14 VTAIL.t6 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X15 VDD2.t2 VN.t7 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=6.7041 ps=35.16 w=17.19 l=2.69
X16 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X17 VDD1.t0 VP.t5 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=2.83635 ps=17.52 w=17.19 l=2.69
X18 VDD2.t0 VN.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=6.7041 ps=35.16 w=17.19 l=2.69
X19 VDD1.t5 VP.t6 VTAIL.t11 B.t8 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=6.7041 ps=35.16 w=17.19 l=2.69
X20 VDD1.t4 VP.t7 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=6.7041 ps=35.16 w=17.19 l=2.69
X21 VDD1.t9 VP.t8 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X22 VTAIL.t8 VP.t9 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83635 pd=17.52 as=2.83635 ps=17.52 w=17.19 l=2.69
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7041 pd=35.16 as=0 ps=0 w=17.19 l=2.69
R0 VP.n24 VP.t5 184.72
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n23 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n22 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n34 VP.n21 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n20 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n19 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n18 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n48 VP.n16 161.3
R16 VP.n50 VP.n49 161.3
R17 VP.n51 VP.n15 161.3
R18 VP.n53 VP.n52 161.3
R19 VP.n54 VP.n14 161.3
R20 VP.n96 VP.n0 161.3
R21 VP.n95 VP.n94 161.3
R22 VP.n93 VP.n1 161.3
R23 VP.n92 VP.n91 161.3
R24 VP.n90 VP.n2 161.3
R25 VP.n89 VP.n88 161.3
R26 VP.n87 VP.n86 161.3
R27 VP.n85 VP.n4 161.3
R28 VP.n84 VP.n83 161.3
R29 VP.n82 VP.n5 161.3
R30 VP.n81 VP.n80 161.3
R31 VP.n79 VP.n6 161.3
R32 VP.n78 VP.n77 161.3
R33 VP.n76 VP.n7 161.3
R34 VP.n75 VP.n74 161.3
R35 VP.n73 VP.n8 161.3
R36 VP.n72 VP.n71 161.3
R37 VP.n70 VP.n9 161.3
R38 VP.n69 VP.n68 161.3
R39 VP.n66 VP.n10 161.3
R40 VP.n65 VP.n64 161.3
R41 VP.n63 VP.n11 161.3
R42 VP.n62 VP.n61 161.3
R43 VP.n60 VP.n12 161.3
R44 VP.n59 VP.n58 161.3
R45 VP.n78 VP.t8 154.007
R46 VP.n13 VP.t2 154.007
R47 VP.n67 VP.t0 154.007
R48 VP.n3 VP.t9 154.007
R49 VP.n97 VP.t6 154.007
R50 VP.n36 VP.t3 154.007
R51 VP.n55 VP.t7 154.007
R52 VP.n17 VP.t1 154.007
R53 VP.n25 VP.t4 154.007
R54 VP.n57 VP.n13 108.799
R55 VP.n98 VP.n97 108.799
R56 VP.n56 VP.n55 108.799
R57 VP.n25 VP.n24 72.37
R58 VP.n57 VP.n56 57.4541
R59 VP.n61 VP.n11 43.4072
R60 VP.n91 VP.n1 43.4072
R61 VP.n49 VP.n15 43.4072
R62 VP.n73 VP.n72 41.4647
R63 VP.n84 VP.n5 41.4647
R64 VP.n42 VP.n19 41.4647
R65 VP.n31 VP.n30 41.4647
R66 VP.n74 VP.n73 39.5221
R67 VP.n80 VP.n5 39.5221
R68 VP.n38 VP.n19 39.5221
R69 VP.n32 VP.n31 39.5221
R70 VP.n65 VP.n11 37.5796
R71 VP.n91 VP.n90 37.5796
R72 VP.n49 VP.n48 37.5796
R73 VP.n60 VP.n59 24.4675
R74 VP.n61 VP.n60 24.4675
R75 VP.n66 VP.n65 24.4675
R76 VP.n68 VP.n9 24.4675
R77 VP.n72 VP.n9 24.4675
R78 VP.n74 VP.n7 24.4675
R79 VP.n78 VP.n7 24.4675
R80 VP.n79 VP.n78 24.4675
R81 VP.n80 VP.n79 24.4675
R82 VP.n85 VP.n84 24.4675
R83 VP.n86 VP.n85 24.4675
R84 VP.n90 VP.n89 24.4675
R85 VP.n95 VP.n1 24.4675
R86 VP.n96 VP.n95 24.4675
R87 VP.n53 VP.n15 24.4675
R88 VP.n54 VP.n53 24.4675
R89 VP.n43 VP.n42 24.4675
R90 VP.n44 VP.n43 24.4675
R91 VP.n48 VP.n47 24.4675
R92 VP.n32 VP.n21 24.4675
R93 VP.n36 VP.n21 24.4675
R94 VP.n37 VP.n36 24.4675
R95 VP.n38 VP.n37 24.4675
R96 VP.n26 VP.n23 24.4675
R97 VP.n30 VP.n23 24.4675
R98 VP.n67 VP.n66 23.4888
R99 VP.n89 VP.n3 23.4888
R100 VP.n47 VP.n17 23.4888
R101 VP.n27 VP.n24 7.37486
R102 VP.n59 VP.n13 1.95786
R103 VP.n97 VP.n96 1.95786
R104 VP.n55 VP.n54 1.95786
R105 VP.n68 VP.n67 0.97918
R106 VP.n86 VP.n3 0.97918
R107 VP.n44 VP.n17 0.97918
R108 VP.n26 VP.n25 0.97918
R109 VP.n56 VP.n14 0.278367
R110 VP.n58 VP.n57 0.278367
R111 VP.n98 VP.n0 0.278367
R112 VP.n28 VP.n27 0.189894
R113 VP.n29 VP.n28 0.189894
R114 VP.n29 VP.n22 0.189894
R115 VP.n33 VP.n22 0.189894
R116 VP.n34 VP.n33 0.189894
R117 VP.n35 VP.n34 0.189894
R118 VP.n35 VP.n20 0.189894
R119 VP.n39 VP.n20 0.189894
R120 VP.n40 VP.n39 0.189894
R121 VP.n41 VP.n40 0.189894
R122 VP.n41 VP.n18 0.189894
R123 VP.n45 VP.n18 0.189894
R124 VP.n46 VP.n45 0.189894
R125 VP.n46 VP.n16 0.189894
R126 VP.n50 VP.n16 0.189894
R127 VP.n51 VP.n50 0.189894
R128 VP.n52 VP.n51 0.189894
R129 VP.n52 VP.n14 0.189894
R130 VP.n58 VP.n12 0.189894
R131 VP.n62 VP.n12 0.189894
R132 VP.n63 VP.n62 0.189894
R133 VP.n64 VP.n63 0.189894
R134 VP.n64 VP.n10 0.189894
R135 VP.n69 VP.n10 0.189894
R136 VP.n70 VP.n69 0.189894
R137 VP.n71 VP.n70 0.189894
R138 VP.n71 VP.n8 0.189894
R139 VP.n75 VP.n8 0.189894
R140 VP.n76 VP.n75 0.189894
R141 VP.n77 VP.n76 0.189894
R142 VP.n77 VP.n6 0.189894
R143 VP.n81 VP.n6 0.189894
R144 VP.n82 VP.n81 0.189894
R145 VP.n83 VP.n82 0.189894
R146 VP.n83 VP.n4 0.189894
R147 VP.n87 VP.n4 0.189894
R148 VP.n88 VP.n87 0.189894
R149 VP.n88 VP.n2 0.189894
R150 VP.n92 VP.n2 0.189894
R151 VP.n93 VP.n92 0.189894
R152 VP.n94 VP.n93 0.189894
R153 VP.n94 VP.n0 0.189894
R154 VP VP.n98 0.153454
R155 VDD1.n1 VDD1.t0 65.0391
R156 VDD1.n3 VDD1.t7 65.039
R157 VDD1.n5 VDD1.n4 63.1809
R158 VDD1.n1 VDD1.n0 61.2839
R159 VDD1.n7 VDD1.n6 61.2837
R160 VDD1.n3 VDD1.n2 61.2836
R161 VDD1.n7 VDD1.n5 52.7854
R162 VDD1 VDD1.n7 1.8949
R163 VDD1.n6 VDD1.t2 1.15233
R164 VDD1.n6 VDD1.t4 1.15233
R165 VDD1.n0 VDD1.t1 1.15233
R166 VDD1.n0 VDD1.t6 1.15233
R167 VDD1.n4 VDD1.t8 1.15233
R168 VDD1.n4 VDD1.t5 1.15233
R169 VDD1.n2 VDD1.t3 1.15233
R170 VDD1.n2 VDD1.t9 1.15233
R171 VDD1 VDD1.n1 0.709552
R172 VDD1.n5 VDD1.n3 0.596016
R173 VTAIL.n11 VTAIL.t18 45.7569
R174 VTAIL.n17 VTAIL.t7 45.7567
R175 VTAIL.n2 VTAIL.t11 45.7567
R176 VTAIL.n16 VTAIL.t10 45.7567
R177 VTAIL.n15 VTAIL.n14 44.6051
R178 VTAIL.n13 VTAIL.n12 44.6051
R179 VTAIL.n10 VTAIL.n9 44.6051
R180 VTAIL.n8 VTAIL.n7 44.6051
R181 VTAIL.n19 VTAIL.n18 44.6049
R182 VTAIL.n1 VTAIL.n0 44.6049
R183 VTAIL.n4 VTAIL.n3 44.6049
R184 VTAIL.n6 VTAIL.n5 44.6049
R185 VTAIL.n8 VTAIL.n6 32.3927
R186 VTAIL.n17 VTAIL.n16 29.7893
R187 VTAIL.n10 VTAIL.n8 2.60395
R188 VTAIL.n11 VTAIL.n10 2.60395
R189 VTAIL.n15 VTAIL.n13 2.60395
R190 VTAIL.n16 VTAIL.n15 2.60395
R191 VTAIL.n6 VTAIL.n4 2.60395
R192 VTAIL.n4 VTAIL.n2 2.60395
R193 VTAIL.n19 VTAIL.n17 2.60395
R194 VTAIL VTAIL.n1 2.01128
R195 VTAIL.n13 VTAIL.n11 1.77205
R196 VTAIL.n2 VTAIL.n1 1.77205
R197 VTAIL.n18 VTAIL.t3 1.15233
R198 VTAIL.n18 VTAIL.t6 1.15233
R199 VTAIL.n0 VTAIL.t2 1.15233
R200 VTAIL.n0 VTAIL.t5 1.15233
R201 VTAIL.n3 VTAIL.t9 1.15233
R202 VTAIL.n3 VTAIL.t8 1.15233
R203 VTAIL.n5 VTAIL.t15 1.15233
R204 VTAIL.n5 VTAIL.t17 1.15233
R205 VTAIL.n14 VTAIL.t14 1.15233
R206 VTAIL.n14 VTAIL.t16 1.15233
R207 VTAIL.n12 VTAIL.t12 1.15233
R208 VTAIL.n12 VTAIL.t13 1.15233
R209 VTAIL.n9 VTAIL.t4 1.15233
R210 VTAIL.n9 VTAIL.t0 1.15233
R211 VTAIL.n7 VTAIL.t19 1.15233
R212 VTAIL.n7 VTAIL.t1 1.15233
R213 VTAIL VTAIL.n19 0.593172
R214 B.n1120 B.n1119 585
R215 B.n1121 B.n1120 585
R216 B.n423 B.n174 585
R217 B.n422 B.n421 585
R218 B.n420 B.n419 585
R219 B.n418 B.n417 585
R220 B.n416 B.n415 585
R221 B.n414 B.n413 585
R222 B.n412 B.n411 585
R223 B.n410 B.n409 585
R224 B.n408 B.n407 585
R225 B.n406 B.n405 585
R226 B.n404 B.n403 585
R227 B.n402 B.n401 585
R228 B.n400 B.n399 585
R229 B.n398 B.n397 585
R230 B.n396 B.n395 585
R231 B.n394 B.n393 585
R232 B.n392 B.n391 585
R233 B.n390 B.n389 585
R234 B.n388 B.n387 585
R235 B.n386 B.n385 585
R236 B.n384 B.n383 585
R237 B.n382 B.n381 585
R238 B.n380 B.n379 585
R239 B.n378 B.n377 585
R240 B.n376 B.n375 585
R241 B.n374 B.n373 585
R242 B.n372 B.n371 585
R243 B.n370 B.n369 585
R244 B.n368 B.n367 585
R245 B.n366 B.n365 585
R246 B.n364 B.n363 585
R247 B.n362 B.n361 585
R248 B.n360 B.n359 585
R249 B.n358 B.n357 585
R250 B.n356 B.n355 585
R251 B.n354 B.n353 585
R252 B.n352 B.n351 585
R253 B.n350 B.n349 585
R254 B.n348 B.n347 585
R255 B.n346 B.n345 585
R256 B.n344 B.n343 585
R257 B.n342 B.n341 585
R258 B.n340 B.n339 585
R259 B.n338 B.n337 585
R260 B.n336 B.n335 585
R261 B.n334 B.n333 585
R262 B.n332 B.n331 585
R263 B.n330 B.n329 585
R264 B.n328 B.n327 585
R265 B.n326 B.n325 585
R266 B.n324 B.n323 585
R267 B.n322 B.n321 585
R268 B.n320 B.n319 585
R269 B.n318 B.n317 585
R270 B.n316 B.n315 585
R271 B.n314 B.n313 585
R272 B.n312 B.n311 585
R273 B.n310 B.n309 585
R274 B.n308 B.n307 585
R275 B.n306 B.n305 585
R276 B.n304 B.n303 585
R277 B.n302 B.n301 585
R278 B.n300 B.n299 585
R279 B.n298 B.n297 585
R280 B.n296 B.n295 585
R281 B.n293 B.n292 585
R282 B.n291 B.n290 585
R283 B.n289 B.n288 585
R284 B.n287 B.n286 585
R285 B.n285 B.n284 585
R286 B.n283 B.n282 585
R287 B.n281 B.n280 585
R288 B.n279 B.n278 585
R289 B.n277 B.n276 585
R290 B.n275 B.n274 585
R291 B.n273 B.n272 585
R292 B.n271 B.n270 585
R293 B.n269 B.n268 585
R294 B.n267 B.n266 585
R295 B.n265 B.n264 585
R296 B.n263 B.n262 585
R297 B.n261 B.n260 585
R298 B.n259 B.n258 585
R299 B.n257 B.n256 585
R300 B.n255 B.n254 585
R301 B.n253 B.n252 585
R302 B.n251 B.n250 585
R303 B.n249 B.n248 585
R304 B.n247 B.n246 585
R305 B.n245 B.n244 585
R306 B.n243 B.n242 585
R307 B.n241 B.n240 585
R308 B.n239 B.n238 585
R309 B.n237 B.n236 585
R310 B.n235 B.n234 585
R311 B.n233 B.n232 585
R312 B.n231 B.n230 585
R313 B.n229 B.n228 585
R314 B.n227 B.n226 585
R315 B.n225 B.n224 585
R316 B.n223 B.n222 585
R317 B.n221 B.n220 585
R318 B.n219 B.n218 585
R319 B.n217 B.n216 585
R320 B.n215 B.n214 585
R321 B.n213 B.n212 585
R322 B.n211 B.n210 585
R323 B.n209 B.n208 585
R324 B.n207 B.n206 585
R325 B.n205 B.n204 585
R326 B.n203 B.n202 585
R327 B.n201 B.n200 585
R328 B.n199 B.n198 585
R329 B.n197 B.n196 585
R330 B.n195 B.n194 585
R331 B.n193 B.n192 585
R332 B.n191 B.n190 585
R333 B.n189 B.n188 585
R334 B.n187 B.n186 585
R335 B.n185 B.n184 585
R336 B.n183 B.n182 585
R337 B.n181 B.n180 585
R338 B.n1118 B.n112 585
R339 B.n1122 B.n112 585
R340 B.n1117 B.n111 585
R341 B.n1123 B.n111 585
R342 B.n1116 B.n1115 585
R343 B.n1115 B.n107 585
R344 B.n1114 B.n106 585
R345 B.n1129 B.n106 585
R346 B.n1113 B.n105 585
R347 B.n1130 B.n105 585
R348 B.n1112 B.n104 585
R349 B.n1131 B.n104 585
R350 B.n1111 B.n1110 585
R351 B.n1110 B.n100 585
R352 B.n1109 B.n99 585
R353 B.n1137 B.n99 585
R354 B.n1108 B.n98 585
R355 B.n1138 B.n98 585
R356 B.n1107 B.n97 585
R357 B.n1139 B.n97 585
R358 B.n1106 B.n1105 585
R359 B.n1105 B.n93 585
R360 B.n1104 B.n92 585
R361 B.n1145 B.n92 585
R362 B.n1103 B.n91 585
R363 B.n1146 B.n91 585
R364 B.n1102 B.n90 585
R365 B.n1147 B.n90 585
R366 B.n1101 B.n1100 585
R367 B.n1100 B.n86 585
R368 B.n1099 B.n85 585
R369 B.n1153 B.n85 585
R370 B.n1098 B.n84 585
R371 B.n1154 B.n84 585
R372 B.n1097 B.n83 585
R373 B.n1155 B.n83 585
R374 B.n1096 B.n1095 585
R375 B.n1095 B.n79 585
R376 B.n1094 B.n78 585
R377 B.n1161 B.n78 585
R378 B.n1093 B.n77 585
R379 B.n1162 B.n77 585
R380 B.n1092 B.n76 585
R381 B.n1163 B.n76 585
R382 B.n1091 B.n1090 585
R383 B.n1090 B.n72 585
R384 B.n1089 B.n71 585
R385 B.n1169 B.n71 585
R386 B.n1088 B.n70 585
R387 B.n1170 B.n70 585
R388 B.n1087 B.n69 585
R389 B.n1171 B.n69 585
R390 B.n1086 B.n1085 585
R391 B.n1085 B.n65 585
R392 B.n1084 B.n64 585
R393 B.n1177 B.n64 585
R394 B.n1083 B.n63 585
R395 B.n1178 B.n63 585
R396 B.n1082 B.n62 585
R397 B.n1179 B.n62 585
R398 B.n1081 B.n1080 585
R399 B.n1080 B.n58 585
R400 B.n1079 B.n57 585
R401 B.n1185 B.n57 585
R402 B.n1078 B.n56 585
R403 B.n1186 B.n56 585
R404 B.n1077 B.n55 585
R405 B.n1187 B.n55 585
R406 B.n1076 B.n1075 585
R407 B.n1075 B.n51 585
R408 B.n1074 B.n50 585
R409 B.n1193 B.n50 585
R410 B.n1073 B.n49 585
R411 B.n1194 B.n49 585
R412 B.n1072 B.n48 585
R413 B.n1195 B.n48 585
R414 B.n1071 B.n1070 585
R415 B.n1070 B.n44 585
R416 B.n1069 B.n43 585
R417 B.n1201 B.n43 585
R418 B.n1068 B.n42 585
R419 B.n1202 B.n42 585
R420 B.n1067 B.n41 585
R421 B.n1203 B.n41 585
R422 B.n1066 B.n1065 585
R423 B.n1065 B.n37 585
R424 B.n1064 B.n36 585
R425 B.n1209 B.n36 585
R426 B.n1063 B.n35 585
R427 B.n1210 B.n35 585
R428 B.n1062 B.n34 585
R429 B.n1211 B.n34 585
R430 B.n1061 B.n1060 585
R431 B.n1060 B.n33 585
R432 B.n1059 B.n29 585
R433 B.n1217 B.n29 585
R434 B.n1058 B.n28 585
R435 B.n1218 B.n28 585
R436 B.n1057 B.n27 585
R437 B.n1219 B.n27 585
R438 B.n1056 B.n1055 585
R439 B.n1055 B.n23 585
R440 B.n1054 B.n22 585
R441 B.n1225 B.n22 585
R442 B.n1053 B.n21 585
R443 B.n1226 B.n21 585
R444 B.n1052 B.n20 585
R445 B.n1227 B.n20 585
R446 B.n1051 B.n1050 585
R447 B.n1050 B.n16 585
R448 B.n1049 B.n15 585
R449 B.n1233 B.n15 585
R450 B.n1048 B.n14 585
R451 B.n1234 B.n14 585
R452 B.n1047 B.n13 585
R453 B.n1235 B.n13 585
R454 B.n1046 B.n1045 585
R455 B.n1045 B.n12 585
R456 B.n1044 B.n1043 585
R457 B.n1044 B.n8 585
R458 B.n1042 B.n7 585
R459 B.n1242 B.n7 585
R460 B.n1041 B.n6 585
R461 B.n1243 B.n6 585
R462 B.n1040 B.n5 585
R463 B.n1244 B.n5 585
R464 B.n1039 B.n1038 585
R465 B.n1038 B.n4 585
R466 B.n1037 B.n424 585
R467 B.n1037 B.n1036 585
R468 B.n1027 B.n425 585
R469 B.n426 B.n425 585
R470 B.n1029 B.n1028 585
R471 B.n1030 B.n1029 585
R472 B.n1026 B.n431 585
R473 B.n431 B.n430 585
R474 B.n1025 B.n1024 585
R475 B.n1024 B.n1023 585
R476 B.n433 B.n432 585
R477 B.n434 B.n433 585
R478 B.n1016 B.n1015 585
R479 B.n1017 B.n1016 585
R480 B.n1014 B.n439 585
R481 B.n439 B.n438 585
R482 B.n1013 B.n1012 585
R483 B.n1012 B.n1011 585
R484 B.n441 B.n440 585
R485 B.n442 B.n441 585
R486 B.n1004 B.n1003 585
R487 B.n1005 B.n1004 585
R488 B.n1002 B.n447 585
R489 B.n447 B.n446 585
R490 B.n1001 B.n1000 585
R491 B.n1000 B.n999 585
R492 B.n449 B.n448 585
R493 B.n992 B.n449 585
R494 B.n991 B.n990 585
R495 B.n993 B.n991 585
R496 B.n989 B.n454 585
R497 B.n454 B.n453 585
R498 B.n988 B.n987 585
R499 B.n987 B.n986 585
R500 B.n456 B.n455 585
R501 B.n457 B.n456 585
R502 B.n979 B.n978 585
R503 B.n980 B.n979 585
R504 B.n977 B.n462 585
R505 B.n462 B.n461 585
R506 B.n976 B.n975 585
R507 B.n975 B.n974 585
R508 B.n464 B.n463 585
R509 B.n465 B.n464 585
R510 B.n967 B.n966 585
R511 B.n968 B.n967 585
R512 B.n965 B.n470 585
R513 B.n470 B.n469 585
R514 B.n964 B.n963 585
R515 B.n963 B.n962 585
R516 B.n472 B.n471 585
R517 B.n473 B.n472 585
R518 B.n955 B.n954 585
R519 B.n956 B.n955 585
R520 B.n953 B.n478 585
R521 B.n478 B.n477 585
R522 B.n952 B.n951 585
R523 B.n951 B.n950 585
R524 B.n480 B.n479 585
R525 B.n481 B.n480 585
R526 B.n943 B.n942 585
R527 B.n944 B.n943 585
R528 B.n941 B.n485 585
R529 B.n489 B.n485 585
R530 B.n940 B.n939 585
R531 B.n939 B.n938 585
R532 B.n487 B.n486 585
R533 B.n488 B.n487 585
R534 B.n931 B.n930 585
R535 B.n932 B.n931 585
R536 B.n929 B.n494 585
R537 B.n494 B.n493 585
R538 B.n928 B.n927 585
R539 B.n927 B.n926 585
R540 B.n496 B.n495 585
R541 B.n497 B.n496 585
R542 B.n919 B.n918 585
R543 B.n920 B.n919 585
R544 B.n917 B.n502 585
R545 B.n502 B.n501 585
R546 B.n916 B.n915 585
R547 B.n915 B.n914 585
R548 B.n504 B.n503 585
R549 B.n505 B.n504 585
R550 B.n907 B.n906 585
R551 B.n908 B.n907 585
R552 B.n905 B.n510 585
R553 B.n510 B.n509 585
R554 B.n904 B.n903 585
R555 B.n903 B.n902 585
R556 B.n512 B.n511 585
R557 B.n513 B.n512 585
R558 B.n895 B.n894 585
R559 B.n896 B.n895 585
R560 B.n893 B.n518 585
R561 B.n518 B.n517 585
R562 B.n892 B.n891 585
R563 B.n891 B.n890 585
R564 B.n520 B.n519 585
R565 B.n521 B.n520 585
R566 B.n883 B.n882 585
R567 B.n884 B.n883 585
R568 B.n881 B.n526 585
R569 B.n526 B.n525 585
R570 B.n880 B.n879 585
R571 B.n879 B.n878 585
R572 B.n528 B.n527 585
R573 B.n529 B.n528 585
R574 B.n871 B.n870 585
R575 B.n872 B.n871 585
R576 B.n869 B.n534 585
R577 B.n534 B.n533 585
R578 B.n868 B.n867 585
R579 B.n867 B.n866 585
R580 B.n536 B.n535 585
R581 B.n537 B.n536 585
R582 B.n859 B.n858 585
R583 B.n860 B.n859 585
R584 B.n857 B.n542 585
R585 B.n542 B.n541 585
R586 B.n851 B.n850 585
R587 B.n849 B.n605 585
R588 B.n848 B.n604 585
R589 B.n853 B.n604 585
R590 B.n847 B.n846 585
R591 B.n845 B.n844 585
R592 B.n843 B.n842 585
R593 B.n841 B.n840 585
R594 B.n839 B.n838 585
R595 B.n837 B.n836 585
R596 B.n835 B.n834 585
R597 B.n833 B.n832 585
R598 B.n831 B.n830 585
R599 B.n829 B.n828 585
R600 B.n827 B.n826 585
R601 B.n825 B.n824 585
R602 B.n823 B.n822 585
R603 B.n821 B.n820 585
R604 B.n819 B.n818 585
R605 B.n817 B.n816 585
R606 B.n815 B.n814 585
R607 B.n813 B.n812 585
R608 B.n811 B.n810 585
R609 B.n809 B.n808 585
R610 B.n807 B.n806 585
R611 B.n805 B.n804 585
R612 B.n803 B.n802 585
R613 B.n801 B.n800 585
R614 B.n799 B.n798 585
R615 B.n797 B.n796 585
R616 B.n795 B.n794 585
R617 B.n793 B.n792 585
R618 B.n791 B.n790 585
R619 B.n789 B.n788 585
R620 B.n787 B.n786 585
R621 B.n785 B.n784 585
R622 B.n783 B.n782 585
R623 B.n781 B.n780 585
R624 B.n779 B.n778 585
R625 B.n777 B.n776 585
R626 B.n775 B.n774 585
R627 B.n773 B.n772 585
R628 B.n771 B.n770 585
R629 B.n769 B.n768 585
R630 B.n767 B.n766 585
R631 B.n765 B.n764 585
R632 B.n763 B.n762 585
R633 B.n761 B.n760 585
R634 B.n759 B.n758 585
R635 B.n757 B.n756 585
R636 B.n755 B.n754 585
R637 B.n753 B.n752 585
R638 B.n751 B.n750 585
R639 B.n749 B.n748 585
R640 B.n747 B.n746 585
R641 B.n745 B.n744 585
R642 B.n743 B.n742 585
R643 B.n741 B.n740 585
R644 B.n739 B.n738 585
R645 B.n737 B.n736 585
R646 B.n735 B.n734 585
R647 B.n733 B.n732 585
R648 B.n731 B.n730 585
R649 B.n729 B.n728 585
R650 B.n727 B.n726 585
R651 B.n725 B.n724 585
R652 B.n723 B.n722 585
R653 B.n720 B.n719 585
R654 B.n718 B.n717 585
R655 B.n716 B.n715 585
R656 B.n714 B.n713 585
R657 B.n712 B.n711 585
R658 B.n710 B.n709 585
R659 B.n708 B.n707 585
R660 B.n706 B.n705 585
R661 B.n704 B.n703 585
R662 B.n702 B.n701 585
R663 B.n700 B.n699 585
R664 B.n698 B.n697 585
R665 B.n696 B.n695 585
R666 B.n694 B.n693 585
R667 B.n692 B.n691 585
R668 B.n690 B.n689 585
R669 B.n688 B.n687 585
R670 B.n686 B.n685 585
R671 B.n684 B.n683 585
R672 B.n682 B.n681 585
R673 B.n680 B.n679 585
R674 B.n678 B.n677 585
R675 B.n676 B.n675 585
R676 B.n674 B.n673 585
R677 B.n672 B.n671 585
R678 B.n670 B.n669 585
R679 B.n668 B.n667 585
R680 B.n666 B.n665 585
R681 B.n664 B.n663 585
R682 B.n662 B.n661 585
R683 B.n660 B.n659 585
R684 B.n658 B.n657 585
R685 B.n656 B.n655 585
R686 B.n654 B.n653 585
R687 B.n652 B.n651 585
R688 B.n650 B.n649 585
R689 B.n648 B.n647 585
R690 B.n646 B.n645 585
R691 B.n644 B.n643 585
R692 B.n642 B.n641 585
R693 B.n640 B.n639 585
R694 B.n638 B.n637 585
R695 B.n636 B.n635 585
R696 B.n634 B.n633 585
R697 B.n632 B.n631 585
R698 B.n630 B.n629 585
R699 B.n628 B.n627 585
R700 B.n626 B.n625 585
R701 B.n624 B.n623 585
R702 B.n622 B.n621 585
R703 B.n620 B.n619 585
R704 B.n618 B.n617 585
R705 B.n616 B.n615 585
R706 B.n614 B.n613 585
R707 B.n612 B.n611 585
R708 B.n544 B.n543 585
R709 B.n856 B.n855 585
R710 B.n540 B.n539 585
R711 B.n541 B.n540 585
R712 B.n862 B.n861 585
R713 B.n861 B.n860 585
R714 B.n863 B.n538 585
R715 B.n538 B.n537 585
R716 B.n865 B.n864 585
R717 B.n866 B.n865 585
R718 B.n532 B.n531 585
R719 B.n533 B.n532 585
R720 B.n874 B.n873 585
R721 B.n873 B.n872 585
R722 B.n875 B.n530 585
R723 B.n530 B.n529 585
R724 B.n877 B.n876 585
R725 B.n878 B.n877 585
R726 B.n524 B.n523 585
R727 B.n525 B.n524 585
R728 B.n886 B.n885 585
R729 B.n885 B.n884 585
R730 B.n887 B.n522 585
R731 B.n522 B.n521 585
R732 B.n889 B.n888 585
R733 B.n890 B.n889 585
R734 B.n516 B.n515 585
R735 B.n517 B.n516 585
R736 B.n898 B.n897 585
R737 B.n897 B.n896 585
R738 B.n899 B.n514 585
R739 B.n514 B.n513 585
R740 B.n901 B.n900 585
R741 B.n902 B.n901 585
R742 B.n508 B.n507 585
R743 B.n509 B.n508 585
R744 B.n910 B.n909 585
R745 B.n909 B.n908 585
R746 B.n911 B.n506 585
R747 B.n506 B.n505 585
R748 B.n913 B.n912 585
R749 B.n914 B.n913 585
R750 B.n500 B.n499 585
R751 B.n501 B.n500 585
R752 B.n922 B.n921 585
R753 B.n921 B.n920 585
R754 B.n923 B.n498 585
R755 B.n498 B.n497 585
R756 B.n925 B.n924 585
R757 B.n926 B.n925 585
R758 B.n492 B.n491 585
R759 B.n493 B.n492 585
R760 B.n934 B.n933 585
R761 B.n933 B.n932 585
R762 B.n935 B.n490 585
R763 B.n490 B.n488 585
R764 B.n937 B.n936 585
R765 B.n938 B.n937 585
R766 B.n484 B.n483 585
R767 B.n489 B.n484 585
R768 B.n946 B.n945 585
R769 B.n945 B.n944 585
R770 B.n947 B.n482 585
R771 B.n482 B.n481 585
R772 B.n949 B.n948 585
R773 B.n950 B.n949 585
R774 B.n476 B.n475 585
R775 B.n477 B.n476 585
R776 B.n958 B.n957 585
R777 B.n957 B.n956 585
R778 B.n959 B.n474 585
R779 B.n474 B.n473 585
R780 B.n961 B.n960 585
R781 B.n962 B.n961 585
R782 B.n468 B.n467 585
R783 B.n469 B.n468 585
R784 B.n970 B.n969 585
R785 B.n969 B.n968 585
R786 B.n971 B.n466 585
R787 B.n466 B.n465 585
R788 B.n973 B.n972 585
R789 B.n974 B.n973 585
R790 B.n460 B.n459 585
R791 B.n461 B.n460 585
R792 B.n982 B.n981 585
R793 B.n981 B.n980 585
R794 B.n983 B.n458 585
R795 B.n458 B.n457 585
R796 B.n985 B.n984 585
R797 B.n986 B.n985 585
R798 B.n452 B.n451 585
R799 B.n453 B.n452 585
R800 B.n995 B.n994 585
R801 B.n994 B.n993 585
R802 B.n996 B.n450 585
R803 B.n992 B.n450 585
R804 B.n998 B.n997 585
R805 B.n999 B.n998 585
R806 B.n445 B.n444 585
R807 B.n446 B.n445 585
R808 B.n1007 B.n1006 585
R809 B.n1006 B.n1005 585
R810 B.n1008 B.n443 585
R811 B.n443 B.n442 585
R812 B.n1010 B.n1009 585
R813 B.n1011 B.n1010 585
R814 B.n437 B.n436 585
R815 B.n438 B.n437 585
R816 B.n1019 B.n1018 585
R817 B.n1018 B.n1017 585
R818 B.n1020 B.n435 585
R819 B.n435 B.n434 585
R820 B.n1022 B.n1021 585
R821 B.n1023 B.n1022 585
R822 B.n429 B.n428 585
R823 B.n430 B.n429 585
R824 B.n1032 B.n1031 585
R825 B.n1031 B.n1030 585
R826 B.n1033 B.n427 585
R827 B.n427 B.n426 585
R828 B.n1035 B.n1034 585
R829 B.n1036 B.n1035 585
R830 B.n3 B.n0 585
R831 B.n4 B.n3 585
R832 B.n1241 B.n1 585
R833 B.n1242 B.n1241 585
R834 B.n1240 B.n1239 585
R835 B.n1240 B.n8 585
R836 B.n1238 B.n9 585
R837 B.n12 B.n9 585
R838 B.n1237 B.n1236 585
R839 B.n1236 B.n1235 585
R840 B.n11 B.n10 585
R841 B.n1234 B.n11 585
R842 B.n1232 B.n1231 585
R843 B.n1233 B.n1232 585
R844 B.n1230 B.n17 585
R845 B.n17 B.n16 585
R846 B.n1229 B.n1228 585
R847 B.n1228 B.n1227 585
R848 B.n19 B.n18 585
R849 B.n1226 B.n19 585
R850 B.n1224 B.n1223 585
R851 B.n1225 B.n1224 585
R852 B.n1222 B.n24 585
R853 B.n24 B.n23 585
R854 B.n1221 B.n1220 585
R855 B.n1220 B.n1219 585
R856 B.n26 B.n25 585
R857 B.n1218 B.n26 585
R858 B.n1216 B.n1215 585
R859 B.n1217 B.n1216 585
R860 B.n1214 B.n30 585
R861 B.n33 B.n30 585
R862 B.n1213 B.n1212 585
R863 B.n1212 B.n1211 585
R864 B.n32 B.n31 585
R865 B.n1210 B.n32 585
R866 B.n1208 B.n1207 585
R867 B.n1209 B.n1208 585
R868 B.n1206 B.n38 585
R869 B.n38 B.n37 585
R870 B.n1205 B.n1204 585
R871 B.n1204 B.n1203 585
R872 B.n40 B.n39 585
R873 B.n1202 B.n40 585
R874 B.n1200 B.n1199 585
R875 B.n1201 B.n1200 585
R876 B.n1198 B.n45 585
R877 B.n45 B.n44 585
R878 B.n1197 B.n1196 585
R879 B.n1196 B.n1195 585
R880 B.n47 B.n46 585
R881 B.n1194 B.n47 585
R882 B.n1192 B.n1191 585
R883 B.n1193 B.n1192 585
R884 B.n1190 B.n52 585
R885 B.n52 B.n51 585
R886 B.n1189 B.n1188 585
R887 B.n1188 B.n1187 585
R888 B.n54 B.n53 585
R889 B.n1186 B.n54 585
R890 B.n1184 B.n1183 585
R891 B.n1185 B.n1184 585
R892 B.n1182 B.n59 585
R893 B.n59 B.n58 585
R894 B.n1181 B.n1180 585
R895 B.n1180 B.n1179 585
R896 B.n61 B.n60 585
R897 B.n1178 B.n61 585
R898 B.n1176 B.n1175 585
R899 B.n1177 B.n1176 585
R900 B.n1174 B.n66 585
R901 B.n66 B.n65 585
R902 B.n1173 B.n1172 585
R903 B.n1172 B.n1171 585
R904 B.n68 B.n67 585
R905 B.n1170 B.n68 585
R906 B.n1168 B.n1167 585
R907 B.n1169 B.n1168 585
R908 B.n1166 B.n73 585
R909 B.n73 B.n72 585
R910 B.n1165 B.n1164 585
R911 B.n1164 B.n1163 585
R912 B.n75 B.n74 585
R913 B.n1162 B.n75 585
R914 B.n1160 B.n1159 585
R915 B.n1161 B.n1160 585
R916 B.n1158 B.n80 585
R917 B.n80 B.n79 585
R918 B.n1157 B.n1156 585
R919 B.n1156 B.n1155 585
R920 B.n82 B.n81 585
R921 B.n1154 B.n82 585
R922 B.n1152 B.n1151 585
R923 B.n1153 B.n1152 585
R924 B.n1150 B.n87 585
R925 B.n87 B.n86 585
R926 B.n1149 B.n1148 585
R927 B.n1148 B.n1147 585
R928 B.n89 B.n88 585
R929 B.n1146 B.n89 585
R930 B.n1144 B.n1143 585
R931 B.n1145 B.n1144 585
R932 B.n1142 B.n94 585
R933 B.n94 B.n93 585
R934 B.n1141 B.n1140 585
R935 B.n1140 B.n1139 585
R936 B.n96 B.n95 585
R937 B.n1138 B.n96 585
R938 B.n1136 B.n1135 585
R939 B.n1137 B.n1136 585
R940 B.n1134 B.n101 585
R941 B.n101 B.n100 585
R942 B.n1133 B.n1132 585
R943 B.n1132 B.n1131 585
R944 B.n103 B.n102 585
R945 B.n1130 B.n103 585
R946 B.n1128 B.n1127 585
R947 B.n1129 B.n1128 585
R948 B.n1126 B.n108 585
R949 B.n108 B.n107 585
R950 B.n1125 B.n1124 585
R951 B.n1124 B.n1123 585
R952 B.n110 B.n109 585
R953 B.n1122 B.n110 585
R954 B.n1245 B.n1244 585
R955 B.n1243 B.n2 585
R956 B.n180 B.n110 511.721
R957 B.n1120 B.n112 511.721
R958 B.n855 B.n542 511.721
R959 B.n851 B.n540 511.721
R960 B.n178 B.t14 362.187
R961 B.n175 B.t21 362.187
R962 B.n609 B.t10 362.187
R963 B.n606 B.t18 362.187
R964 B.n1121 B.n173 256.663
R965 B.n1121 B.n172 256.663
R966 B.n1121 B.n171 256.663
R967 B.n1121 B.n170 256.663
R968 B.n1121 B.n169 256.663
R969 B.n1121 B.n168 256.663
R970 B.n1121 B.n167 256.663
R971 B.n1121 B.n166 256.663
R972 B.n1121 B.n165 256.663
R973 B.n1121 B.n164 256.663
R974 B.n1121 B.n163 256.663
R975 B.n1121 B.n162 256.663
R976 B.n1121 B.n161 256.663
R977 B.n1121 B.n160 256.663
R978 B.n1121 B.n159 256.663
R979 B.n1121 B.n158 256.663
R980 B.n1121 B.n157 256.663
R981 B.n1121 B.n156 256.663
R982 B.n1121 B.n155 256.663
R983 B.n1121 B.n154 256.663
R984 B.n1121 B.n153 256.663
R985 B.n1121 B.n152 256.663
R986 B.n1121 B.n151 256.663
R987 B.n1121 B.n150 256.663
R988 B.n1121 B.n149 256.663
R989 B.n1121 B.n148 256.663
R990 B.n1121 B.n147 256.663
R991 B.n1121 B.n146 256.663
R992 B.n1121 B.n145 256.663
R993 B.n1121 B.n144 256.663
R994 B.n1121 B.n143 256.663
R995 B.n1121 B.n142 256.663
R996 B.n1121 B.n141 256.663
R997 B.n1121 B.n140 256.663
R998 B.n1121 B.n139 256.663
R999 B.n1121 B.n138 256.663
R1000 B.n1121 B.n137 256.663
R1001 B.n1121 B.n136 256.663
R1002 B.n1121 B.n135 256.663
R1003 B.n1121 B.n134 256.663
R1004 B.n1121 B.n133 256.663
R1005 B.n1121 B.n132 256.663
R1006 B.n1121 B.n131 256.663
R1007 B.n1121 B.n130 256.663
R1008 B.n1121 B.n129 256.663
R1009 B.n1121 B.n128 256.663
R1010 B.n1121 B.n127 256.663
R1011 B.n1121 B.n126 256.663
R1012 B.n1121 B.n125 256.663
R1013 B.n1121 B.n124 256.663
R1014 B.n1121 B.n123 256.663
R1015 B.n1121 B.n122 256.663
R1016 B.n1121 B.n121 256.663
R1017 B.n1121 B.n120 256.663
R1018 B.n1121 B.n119 256.663
R1019 B.n1121 B.n118 256.663
R1020 B.n1121 B.n117 256.663
R1021 B.n1121 B.n116 256.663
R1022 B.n1121 B.n115 256.663
R1023 B.n1121 B.n114 256.663
R1024 B.n1121 B.n113 256.663
R1025 B.n853 B.n852 256.663
R1026 B.n853 B.n545 256.663
R1027 B.n853 B.n546 256.663
R1028 B.n853 B.n547 256.663
R1029 B.n853 B.n548 256.663
R1030 B.n853 B.n549 256.663
R1031 B.n853 B.n550 256.663
R1032 B.n853 B.n551 256.663
R1033 B.n853 B.n552 256.663
R1034 B.n853 B.n553 256.663
R1035 B.n853 B.n554 256.663
R1036 B.n853 B.n555 256.663
R1037 B.n853 B.n556 256.663
R1038 B.n853 B.n557 256.663
R1039 B.n853 B.n558 256.663
R1040 B.n853 B.n559 256.663
R1041 B.n853 B.n560 256.663
R1042 B.n853 B.n561 256.663
R1043 B.n853 B.n562 256.663
R1044 B.n853 B.n563 256.663
R1045 B.n853 B.n564 256.663
R1046 B.n853 B.n565 256.663
R1047 B.n853 B.n566 256.663
R1048 B.n853 B.n567 256.663
R1049 B.n853 B.n568 256.663
R1050 B.n853 B.n569 256.663
R1051 B.n853 B.n570 256.663
R1052 B.n853 B.n571 256.663
R1053 B.n853 B.n572 256.663
R1054 B.n853 B.n573 256.663
R1055 B.n853 B.n574 256.663
R1056 B.n853 B.n575 256.663
R1057 B.n853 B.n576 256.663
R1058 B.n853 B.n577 256.663
R1059 B.n853 B.n578 256.663
R1060 B.n853 B.n579 256.663
R1061 B.n853 B.n580 256.663
R1062 B.n853 B.n581 256.663
R1063 B.n853 B.n582 256.663
R1064 B.n853 B.n583 256.663
R1065 B.n853 B.n584 256.663
R1066 B.n853 B.n585 256.663
R1067 B.n853 B.n586 256.663
R1068 B.n853 B.n587 256.663
R1069 B.n853 B.n588 256.663
R1070 B.n853 B.n589 256.663
R1071 B.n853 B.n590 256.663
R1072 B.n853 B.n591 256.663
R1073 B.n853 B.n592 256.663
R1074 B.n853 B.n593 256.663
R1075 B.n853 B.n594 256.663
R1076 B.n853 B.n595 256.663
R1077 B.n853 B.n596 256.663
R1078 B.n853 B.n597 256.663
R1079 B.n853 B.n598 256.663
R1080 B.n853 B.n599 256.663
R1081 B.n853 B.n600 256.663
R1082 B.n853 B.n601 256.663
R1083 B.n853 B.n602 256.663
R1084 B.n853 B.n603 256.663
R1085 B.n854 B.n853 256.663
R1086 B.n1247 B.n1246 256.663
R1087 B.n184 B.n183 163.367
R1088 B.n188 B.n187 163.367
R1089 B.n192 B.n191 163.367
R1090 B.n196 B.n195 163.367
R1091 B.n200 B.n199 163.367
R1092 B.n204 B.n203 163.367
R1093 B.n208 B.n207 163.367
R1094 B.n212 B.n211 163.367
R1095 B.n216 B.n215 163.367
R1096 B.n220 B.n219 163.367
R1097 B.n224 B.n223 163.367
R1098 B.n228 B.n227 163.367
R1099 B.n232 B.n231 163.367
R1100 B.n236 B.n235 163.367
R1101 B.n240 B.n239 163.367
R1102 B.n244 B.n243 163.367
R1103 B.n248 B.n247 163.367
R1104 B.n252 B.n251 163.367
R1105 B.n256 B.n255 163.367
R1106 B.n260 B.n259 163.367
R1107 B.n264 B.n263 163.367
R1108 B.n268 B.n267 163.367
R1109 B.n272 B.n271 163.367
R1110 B.n276 B.n275 163.367
R1111 B.n280 B.n279 163.367
R1112 B.n284 B.n283 163.367
R1113 B.n288 B.n287 163.367
R1114 B.n292 B.n291 163.367
R1115 B.n297 B.n296 163.367
R1116 B.n301 B.n300 163.367
R1117 B.n305 B.n304 163.367
R1118 B.n309 B.n308 163.367
R1119 B.n313 B.n312 163.367
R1120 B.n317 B.n316 163.367
R1121 B.n321 B.n320 163.367
R1122 B.n325 B.n324 163.367
R1123 B.n329 B.n328 163.367
R1124 B.n333 B.n332 163.367
R1125 B.n337 B.n336 163.367
R1126 B.n341 B.n340 163.367
R1127 B.n345 B.n344 163.367
R1128 B.n349 B.n348 163.367
R1129 B.n353 B.n352 163.367
R1130 B.n357 B.n356 163.367
R1131 B.n361 B.n360 163.367
R1132 B.n365 B.n364 163.367
R1133 B.n369 B.n368 163.367
R1134 B.n373 B.n372 163.367
R1135 B.n377 B.n376 163.367
R1136 B.n381 B.n380 163.367
R1137 B.n385 B.n384 163.367
R1138 B.n389 B.n388 163.367
R1139 B.n393 B.n392 163.367
R1140 B.n397 B.n396 163.367
R1141 B.n401 B.n400 163.367
R1142 B.n405 B.n404 163.367
R1143 B.n409 B.n408 163.367
R1144 B.n413 B.n412 163.367
R1145 B.n417 B.n416 163.367
R1146 B.n421 B.n420 163.367
R1147 B.n1120 B.n174 163.367
R1148 B.n859 B.n542 163.367
R1149 B.n859 B.n536 163.367
R1150 B.n867 B.n536 163.367
R1151 B.n867 B.n534 163.367
R1152 B.n871 B.n534 163.367
R1153 B.n871 B.n528 163.367
R1154 B.n879 B.n528 163.367
R1155 B.n879 B.n526 163.367
R1156 B.n883 B.n526 163.367
R1157 B.n883 B.n520 163.367
R1158 B.n891 B.n520 163.367
R1159 B.n891 B.n518 163.367
R1160 B.n895 B.n518 163.367
R1161 B.n895 B.n512 163.367
R1162 B.n903 B.n512 163.367
R1163 B.n903 B.n510 163.367
R1164 B.n907 B.n510 163.367
R1165 B.n907 B.n504 163.367
R1166 B.n915 B.n504 163.367
R1167 B.n915 B.n502 163.367
R1168 B.n919 B.n502 163.367
R1169 B.n919 B.n496 163.367
R1170 B.n927 B.n496 163.367
R1171 B.n927 B.n494 163.367
R1172 B.n931 B.n494 163.367
R1173 B.n931 B.n487 163.367
R1174 B.n939 B.n487 163.367
R1175 B.n939 B.n485 163.367
R1176 B.n943 B.n485 163.367
R1177 B.n943 B.n480 163.367
R1178 B.n951 B.n480 163.367
R1179 B.n951 B.n478 163.367
R1180 B.n955 B.n478 163.367
R1181 B.n955 B.n472 163.367
R1182 B.n963 B.n472 163.367
R1183 B.n963 B.n470 163.367
R1184 B.n967 B.n470 163.367
R1185 B.n967 B.n464 163.367
R1186 B.n975 B.n464 163.367
R1187 B.n975 B.n462 163.367
R1188 B.n979 B.n462 163.367
R1189 B.n979 B.n456 163.367
R1190 B.n987 B.n456 163.367
R1191 B.n987 B.n454 163.367
R1192 B.n991 B.n454 163.367
R1193 B.n991 B.n449 163.367
R1194 B.n1000 B.n449 163.367
R1195 B.n1000 B.n447 163.367
R1196 B.n1004 B.n447 163.367
R1197 B.n1004 B.n441 163.367
R1198 B.n1012 B.n441 163.367
R1199 B.n1012 B.n439 163.367
R1200 B.n1016 B.n439 163.367
R1201 B.n1016 B.n433 163.367
R1202 B.n1024 B.n433 163.367
R1203 B.n1024 B.n431 163.367
R1204 B.n1029 B.n431 163.367
R1205 B.n1029 B.n425 163.367
R1206 B.n1037 B.n425 163.367
R1207 B.n1038 B.n1037 163.367
R1208 B.n1038 B.n5 163.367
R1209 B.n6 B.n5 163.367
R1210 B.n7 B.n6 163.367
R1211 B.n1044 B.n7 163.367
R1212 B.n1045 B.n1044 163.367
R1213 B.n1045 B.n13 163.367
R1214 B.n14 B.n13 163.367
R1215 B.n15 B.n14 163.367
R1216 B.n1050 B.n15 163.367
R1217 B.n1050 B.n20 163.367
R1218 B.n21 B.n20 163.367
R1219 B.n22 B.n21 163.367
R1220 B.n1055 B.n22 163.367
R1221 B.n1055 B.n27 163.367
R1222 B.n28 B.n27 163.367
R1223 B.n29 B.n28 163.367
R1224 B.n1060 B.n29 163.367
R1225 B.n1060 B.n34 163.367
R1226 B.n35 B.n34 163.367
R1227 B.n36 B.n35 163.367
R1228 B.n1065 B.n36 163.367
R1229 B.n1065 B.n41 163.367
R1230 B.n42 B.n41 163.367
R1231 B.n43 B.n42 163.367
R1232 B.n1070 B.n43 163.367
R1233 B.n1070 B.n48 163.367
R1234 B.n49 B.n48 163.367
R1235 B.n50 B.n49 163.367
R1236 B.n1075 B.n50 163.367
R1237 B.n1075 B.n55 163.367
R1238 B.n56 B.n55 163.367
R1239 B.n57 B.n56 163.367
R1240 B.n1080 B.n57 163.367
R1241 B.n1080 B.n62 163.367
R1242 B.n63 B.n62 163.367
R1243 B.n64 B.n63 163.367
R1244 B.n1085 B.n64 163.367
R1245 B.n1085 B.n69 163.367
R1246 B.n70 B.n69 163.367
R1247 B.n71 B.n70 163.367
R1248 B.n1090 B.n71 163.367
R1249 B.n1090 B.n76 163.367
R1250 B.n77 B.n76 163.367
R1251 B.n78 B.n77 163.367
R1252 B.n1095 B.n78 163.367
R1253 B.n1095 B.n83 163.367
R1254 B.n84 B.n83 163.367
R1255 B.n85 B.n84 163.367
R1256 B.n1100 B.n85 163.367
R1257 B.n1100 B.n90 163.367
R1258 B.n91 B.n90 163.367
R1259 B.n92 B.n91 163.367
R1260 B.n1105 B.n92 163.367
R1261 B.n1105 B.n97 163.367
R1262 B.n98 B.n97 163.367
R1263 B.n99 B.n98 163.367
R1264 B.n1110 B.n99 163.367
R1265 B.n1110 B.n104 163.367
R1266 B.n105 B.n104 163.367
R1267 B.n106 B.n105 163.367
R1268 B.n1115 B.n106 163.367
R1269 B.n1115 B.n111 163.367
R1270 B.n112 B.n111 163.367
R1271 B.n605 B.n604 163.367
R1272 B.n846 B.n604 163.367
R1273 B.n844 B.n843 163.367
R1274 B.n840 B.n839 163.367
R1275 B.n836 B.n835 163.367
R1276 B.n832 B.n831 163.367
R1277 B.n828 B.n827 163.367
R1278 B.n824 B.n823 163.367
R1279 B.n820 B.n819 163.367
R1280 B.n816 B.n815 163.367
R1281 B.n812 B.n811 163.367
R1282 B.n808 B.n807 163.367
R1283 B.n804 B.n803 163.367
R1284 B.n800 B.n799 163.367
R1285 B.n796 B.n795 163.367
R1286 B.n792 B.n791 163.367
R1287 B.n788 B.n787 163.367
R1288 B.n784 B.n783 163.367
R1289 B.n780 B.n779 163.367
R1290 B.n776 B.n775 163.367
R1291 B.n772 B.n771 163.367
R1292 B.n768 B.n767 163.367
R1293 B.n764 B.n763 163.367
R1294 B.n760 B.n759 163.367
R1295 B.n756 B.n755 163.367
R1296 B.n752 B.n751 163.367
R1297 B.n748 B.n747 163.367
R1298 B.n744 B.n743 163.367
R1299 B.n740 B.n739 163.367
R1300 B.n736 B.n735 163.367
R1301 B.n732 B.n731 163.367
R1302 B.n728 B.n727 163.367
R1303 B.n724 B.n723 163.367
R1304 B.n719 B.n718 163.367
R1305 B.n715 B.n714 163.367
R1306 B.n711 B.n710 163.367
R1307 B.n707 B.n706 163.367
R1308 B.n703 B.n702 163.367
R1309 B.n699 B.n698 163.367
R1310 B.n695 B.n694 163.367
R1311 B.n691 B.n690 163.367
R1312 B.n687 B.n686 163.367
R1313 B.n683 B.n682 163.367
R1314 B.n679 B.n678 163.367
R1315 B.n675 B.n674 163.367
R1316 B.n671 B.n670 163.367
R1317 B.n667 B.n666 163.367
R1318 B.n663 B.n662 163.367
R1319 B.n659 B.n658 163.367
R1320 B.n655 B.n654 163.367
R1321 B.n651 B.n650 163.367
R1322 B.n647 B.n646 163.367
R1323 B.n643 B.n642 163.367
R1324 B.n639 B.n638 163.367
R1325 B.n635 B.n634 163.367
R1326 B.n631 B.n630 163.367
R1327 B.n627 B.n626 163.367
R1328 B.n623 B.n622 163.367
R1329 B.n619 B.n618 163.367
R1330 B.n615 B.n614 163.367
R1331 B.n611 B.n544 163.367
R1332 B.n861 B.n540 163.367
R1333 B.n861 B.n538 163.367
R1334 B.n865 B.n538 163.367
R1335 B.n865 B.n532 163.367
R1336 B.n873 B.n532 163.367
R1337 B.n873 B.n530 163.367
R1338 B.n877 B.n530 163.367
R1339 B.n877 B.n524 163.367
R1340 B.n885 B.n524 163.367
R1341 B.n885 B.n522 163.367
R1342 B.n889 B.n522 163.367
R1343 B.n889 B.n516 163.367
R1344 B.n897 B.n516 163.367
R1345 B.n897 B.n514 163.367
R1346 B.n901 B.n514 163.367
R1347 B.n901 B.n508 163.367
R1348 B.n909 B.n508 163.367
R1349 B.n909 B.n506 163.367
R1350 B.n913 B.n506 163.367
R1351 B.n913 B.n500 163.367
R1352 B.n921 B.n500 163.367
R1353 B.n921 B.n498 163.367
R1354 B.n925 B.n498 163.367
R1355 B.n925 B.n492 163.367
R1356 B.n933 B.n492 163.367
R1357 B.n933 B.n490 163.367
R1358 B.n937 B.n490 163.367
R1359 B.n937 B.n484 163.367
R1360 B.n945 B.n484 163.367
R1361 B.n945 B.n482 163.367
R1362 B.n949 B.n482 163.367
R1363 B.n949 B.n476 163.367
R1364 B.n957 B.n476 163.367
R1365 B.n957 B.n474 163.367
R1366 B.n961 B.n474 163.367
R1367 B.n961 B.n468 163.367
R1368 B.n969 B.n468 163.367
R1369 B.n969 B.n466 163.367
R1370 B.n973 B.n466 163.367
R1371 B.n973 B.n460 163.367
R1372 B.n981 B.n460 163.367
R1373 B.n981 B.n458 163.367
R1374 B.n985 B.n458 163.367
R1375 B.n985 B.n452 163.367
R1376 B.n994 B.n452 163.367
R1377 B.n994 B.n450 163.367
R1378 B.n998 B.n450 163.367
R1379 B.n998 B.n445 163.367
R1380 B.n1006 B.n445 163.367
R1381 B.n1006 B.n443 163.367
R1382 B.n1010 B.n443 163.367
R1383 B.n1010 B.n437 163.367
R1384 B.n1018 B.n437 163.367
R1385 B.n1018 B.n435 163.367
R1386 B.n1022 B.n435 163.367
R1387 B.n1022 B.n429 163.367
R1388 B.n1031 B.n429 163.367
R1389 B.n1031 B.n427 163.367
R1390 B.n1035 B.n427 163.367
R1391 B.n1035 B.n3 163.367
R1392 B.n1245 B.n3 163.367
R1393 B.n1241 B.n2 163.367
R1394 B.n1241 B.n1240 163.367
R1395 B.n1240 B.n9 163.367
R1396 B.n1236 B.n9 163.367
R1397 B.n1236 B.n11 163.367
R1398 B.n1232 B.n11 163.367
R1399 B.n1232 B.n17 163.367
R1400 B.n1228 B.n17 163.367
R1401 B.n1228 B.n19 163.367
R1402 B.n1224 B.n19 163.367
R1403 B.n1224 B.n24 163.367
R1404 B.n1220 B.n24 163.367
R1405 B.n1220 B.n26 163.367
R1406 B.n1216 B.n26 163.367
R1407 B.n1216 B.n30 163.367
R1408 B.n1212 B.n30 163.367
R1409 B.n1212 B.n32 163.367
R1410 B.n1208 B.n32 163.367
R1411 B.n1208 B.n38 163.367
R1412 B.n1204 B.n38 163.367
R1413 B.n1204 B.n40 163.367
R1414 B.n1200 B.n40 163.367
R1415 B.n1200 B.n45 163.367
R1416 B.n1196 B.n45 163.367
R1417 B.n1196 B.n47 163.367
R1418 B.n1192 B.n47 163.367
R1419 B.n1192 B.n52 163.367
R1420 B.n1188 B.n52 163.367
R1421 B.n1188 B.n54 163.367
R1422 B.n1184 B.n54 163.367
R1423 B.n1184 B.n59 163.367
R1424 B.n1180 B.n59 163.367
R1425 B.n1180 B.n61 163.367
R1426 B.n1176 B.n61 163.367
R1427 B.n1176 B.n66 163.367
R1428 B.n1172 B.n66 163.367
R1429 B.n1172 B.n68 163.367
R1430 B.n1168 B.n68 163.367
R1431 B.n1168 B.n73 163.367
R1432 B.n1164 B.n73 163.367
R1433 B.n1164 B.n75 163.367
R1434 B.n1160 B.n75 163.367
R1435 B.n1160 B.n80 163.367
R1436 B.n1156 B.n80 163.367
R1437 B.n1156 B.n82 163.367
R1438 B.n1152 B.n82 163.367
R1439 B.n1152 B.n87 163.367
R1440 B.n1148 B.n87 163.367
R1441 B.n1148 B.n89 163.367
R1442 B.n1144 B.n89 163.367
R1443 B.n1144 B.n94 163.367
R1444 B.n1140 B.n94 163.367
R1445 B.n1140 B.n96 163.367
R1446 B.n1136 B.n96 163.367
R1447 B.n1136 B.n101 163.367
R1448 B.n1132 B.n101 163.367
R1449 B.n1132 B.n103 163.367
R1450 B.n1128 B.n103 163.367
R1451 B.n1128 B.n108 163.367
R1452 B.n1124 B.n108 163.367
R1453 B.n1124 B.n110 163.367
R1454 B.n175 B.t22 129.554
R1455 B.n609 B.t13 129.554
R1456 B.n178 B.t16 129.531
R1457 B.n606 B.t20 129.531
R1458 B.n180 B.n113 71.676
R1459 B.n184 B.n114 71.676
R1460 B.n188 B.n115 71.676
R1461 B.n192 B.n116 71.676
R1462 B.n196 B.n117 71.676
R1463 B.n200 B.n118 71.676
R1464 B.n204 B.n119 71.676
R1465 B.n208 B.n120 71.676
R1466 B.n212 B.n121 71.676
R1467 B.n216 B.n122 71.676
R1468 B.n220 B.n123 71.676
R1469 B.n224 B.n124 71.676
R1470 B.n228 B.n125 71.676
R1471 B.n232 B.n126 71.676
R1472 B.n236 B.n127 71.676
R1473 B.n240 B.n128 71.676
R1474 B.n244 B.n129 71.676
R1475 B.n248 B.n130 71.676
R1476 B.n252 B.n131 71.676
R1477 B.n256 B.n132 71.676
R1478 B.n260 B.n133 71.676
R1479 B.n264 B.n134 71.676
R1480 B.n268 B.n135 71.676
R1481 B.n272 B.n136 71.676
R1482 B.n276 B.n137 71.676
R1483 B.n280 B.n138 71.676
R1484 B.n284 B.n139 71.676
R1485 B.n288 B.n140 71.676
R1486 B.n292 B.n141 71.676
R1487 B.n297 B.n142 71.676
R1488 B.n301 B.n143 71.676
R1489 B.n305 B.n144 71.676
R1490 B.n309 B.n145 71.676
R1491 B.n313 B.n146 71.676
R1492 B.n317 B.n147 71.676
R1493 B.n321 B.n148 71.676
R1494 B.n325 B.n149 71.676
R1495 B.n329 B.n150 71.676
R1496 B.n333 B.n151 71.676
R1497 B.n337 B.n152 71.676
R1498 B.n341 B.n153 71.676
R1499 B.n345 B.n154 71.676
R1500 B.n349 B.n155 71.676
R1501 B.n353 B.n156 71.676
R1502 B.n357 B.n157 71.676
R1503 B.n361 B.n158 71.676
R1504 B.n365 B.n159 71.676
R1505 B.n369 B.n160 71.676
R1506 B.n373 B.n161 71.676
R1507 B.n377 B.n162 71.676
R1508 B.n381 B.n163 71.676
R1509 B.n385 B.n164 71.676
R1510 B.n389 B.n165 71.676
R1511 B.n393 B.n166 71.676
R1512 B.n397 B.n167 71.676
R1513 B.n401 B.n168 71.676
R1514 B.n405 B.n169 71.676
R1515 B.n409 B.n170 71.676
R1516 B.n413 B.n171 71.676
R1517 B.n417 B.n172 71.676
R1518 B.n421 B.n173 71.676
R1519 B.n174 B.n173 71.676
R1520 B.n420 B.n172 71.676
R1521 B.n416 B.n171 71.676
R1522 B.n412 B.n170 71.676
R1523 B.n408 B.n169 71.676
R1524 B.n404 B.n168 71.676
R1525 B.n400 B.n167 71.676
R1526 B.n396 B.n166 71.676
R1527 B.n392 B.n165 71.676
R1528 B.n388 B.n164 71.676
R1529 B.n384 B.n163 71.676
R1530 B.n380 B.n162 71.676
R1531 B.n376 B.n161 71.676
R1532 B.n372 B.n160 71.676
R1533 B.n368 B.n159 71.676
R1534 B.n364 B.n158 71.676
R1535 B.n360 B.n157 71.676
R1536 B.n356 B.n156 71.676
R1537 B.n352 B.n155 71.676
R1538 B.n348 B.n154 71.676
R1539 B.n344 B.n153 71.676
R1540 B.n340 B.n152 71.676
R1541 B.n336 B.n151 71.676
R1542 B.n332 B.n150 71.676
R1543 B.n328 B.n149 71.676
R1544 B.n324 B.n148 71.676
R1545 B.n320 B.n147 71.676
R1546 B.n316 B.n146 71.676
R1547 B.n312 B.n145 71.676
R1548 B.n308 B.n144 71.676
R1549 B.n304 B.n143 71.676
R1550 B.n300 B.n142 71.676
R1551 B.n296 B.n141 71.676
R1552 B.n291 B.n140 71.676
R1553 B.n287 B.n139 71.676
R1554 B.n283 B.n138 71.676
R1555 B.n279 B.n137 71.676
R1556 B.n275 B.n136 71.676
R1557 B.n271 B.n135 71.676
R1558 B.n267 B.n134 71.676
R1559 B.n263 B.n133 71.676
R1560 B.n259 B.n132 71.676
R1561 B.n255 B.n131 71.676
R1562 B.n251 B.n130 71.676
R1563 B.n247 B.n129 71.676
R1564 B.n243 B.n128 71.676
R1565 B.n239 B.n127 71.676
R1566 B.n235 B.n126 71.676
R1567 B.n231 B.n125 71.676
R1568 B.n227 B.n124 71.676
R1569 B.n223 B.n123 71.676
R1570 B.n219 B.n122 71.676
R1571 B.n215 B.n121 71.676
R1572 B.n211 B.n120 71.676
R1573 B.n207 B.n119 71.676
R1574 B.n203 B.n118 71.676
R1575 B.n199 B.n117 71.676
R1576 B.n195 B.n116 71.676
R1577 B.n191 B.n115 71.676
R1578 B.n187 B.n114 71.676
R1579 B.n183 B.n113 71.676
R1580 B.n852 B.n851 71.676
R1581 B.n846 B.n545 71.676
R1582 B.n843 B.n546 71.676
R1583 B.n839 B.n547 71.676
R1584 B.n835 B.n548 71.676
R1585 B.n831 B.n549 71.676
R1586 B.n827 B.n550 71.676
R1587 B.n823 B.n551 71.676
R1588 B.n819 B.n552 71.676
R1589 B.n815 B.n553 71.676
R1590 B.n811 B.n554 71.676
R1591 B.n807 B.n555 71.676
R1592 B.n803 B.n556 71.676
R1593 B.n799 B.n557 71.676
R1594 B.n795 B.n558 71.676
R1595 B.n791 B.n559 71.676
R1596 B.n787 B.n560 71.676
R1597 B.n783 B.n561 71.676
R1598 B.n779 B.n562 71.676
R1599 B.n775 B.n563 71.676
R1600 B.n771 B.n564 71.676
R1601 B.n767 B.n565 71.676
R1602 B.n763 B.n566 71.676
R1603 B.n759 B.n567 71.676
R1604 B.n755 B.n568 71.676
R1605 B.n751 B.n569 71.676
R1606 B.n747 B.n570 71.676
R1607 B.n743 B.n571 71.676
R1608 B.n739 B.n572 71.676
R1609 B.n735 B.n573 71.676
R1610 B.n731 B.n574 71.676
R1611 B.n727 B.n575 71.676
R1612 B.n723 B.n576 71.676
R1613 B.n718 B.n577 71.676
R1614 B.n714 B.n578 71.676
R1615 B.n710 B.n579 71.676
R1616 B.n706 B.n580 71.676
R1617 B.n702 B.n581 71.676
R1618 B.n698 B.n582 71.676
R1619 B.n694 B.n583 71.676
R1620 B.n690 B.n584 71.676
R1621 B.n686 B.n585 71.676
R1622 B.n682 B.n586 71.676
R1623 B.n678 B.n587 71.676
R1624 B.n674 B.n588 71.676
R1625 B.n670 B.n589 71.676
R1626 B.n666 B.n590 71.676
R1627 B.n662 B.n591 71.676
R1628 B.n658 B.n592 71.676
R1629 B.n654 B.n593 71.676
R1630 B.n650 B.n594 71.676
R1631 B.n646 B.n595 71.676
R1632 B.n642 B.n596 71.676
R1633 B.n638 B.n597 71.676
R1634 B.n634 B.n598 71.676
R1635 B.n630 B.n599 71.676
R1636 B.n626 B.n600 71.676
R1637 B.n622 B.n601 71.676
R1638 B.n618 B.n602 71.676
R1639 B.n614 B.n603 71.676
R1640 B.n854 B.n544 71.676
R1641 B.n852 B.n605 71.676
R1642 B.n844 B.n545 71.676
R1643 B.n840 B.n546 71.676
R1644 B.n836 B.n547 71.676
R1645 B.n832 B.n548 71.676
R1646 B.n828 B.n549 71.676
R1647 B.n824 B.n550 71.676
R1648 B.n820 B.n551 71.676
R1649 B.n816 B.n552 71.676
R1650 B.n812 B.n553 71.676
R1651 B.n808 B.n554 71.676
R1652 B.n804 B.n555 71.676
R1653 B.n800 B.n556 71.676
R1654 B.n796 B.n557 71.676
R1655 B.n792 B.n558 71.676
R1656 B.n788 B.n559 71.676
R1657 B.n784 B.n560 71.676
R1658 B.n780 B.n561 71.676
R1659 B.n776 B.n562 71.676
R1660 B.n772 B.n563 71.676
R1661 B.n768 B.n564 71.676
R1662 B.n764 B.n565 71.676
R1663 B.n760 B.n566 71.676
R1664 B.n756 B.n567 71.676
R1665 B.n752 B.n568 71.676
R1666 B.n748 B.n569 71.676
R1667 B.n744 B.n570 71.676
R1668 B.n740 B.n571 71.676
R1669 B.n736 B.n572 71.676
R1670 B.n732 B.n573 71.676
R1671 B.n728 B.n574 71.676
R1672 B.n724 B.n575 71.676
R1673 B.n719 B.n576 71.676
R1674 B.n715 B.n577 71.676
R1675 B.n711 B.n578 71.676
R1676 B.n707 B.n579 71.676
R1677 B.n703 B.n580 71.676
R1678 B.n699 B.n581 71.676
R1679 B.n695 B.n582 71.676
R1680 B.n691 B.n583 71.676
R1681 B.n687 B.n584 71.676
R1682 B.n683 B.n585 71.676
R1683 B.n679 B.n586 71.676
R1684 B.n675 B.n587 71.676
R1685 B.n671 B.n588 71.676
R1686 B.n667 B.n589 71.676
R1687 B.n663 B.n590 71.676
R1688 B.n659 B.n591 71.676
R1689 B.n655 B.n592 71.676
R1690 B.n651 B.n593 71.676
R1691 B.n647 B.n594 71.676
R1692 B.n643 B.n595 71.676
R1693 B.n639 B.n596 71.676
R1694 B.n635 B.n597 71.676
R1695 B.n631 B.n598 71.676
R1696 B.n627 B.n599 71.676
R1697 B.n623 B.n600 71.676
R1698 B.n619 B.n601 71.676
R1699 B.n615 B.n602 71.676
R1700 B.n611 B.n603 71.676
R1701 B.n855 B.n854 71.676
R1702 B.n1246 B.n1245 71.676
R1703 B.n1246 B.n2 71.676
R1704 B.n176 B.t23 70.9841
R1705 B.n610 B.t12 70.9841
R1706 B.n179 B.t17 70.9613
R1707 B.n607 B.t19 70.9613
R1708 B.n294 B.n179 59.5399
R1709 B.n177 B.n176 59.5399
R1710 B.n721 B.n610 59.5399
R1711 B.n608 B.n607 59.5399
R1712 B.n179 B.n178 58.5702
R1713 B.n176 B.n175 58.5702
R1714 B.n610 B.n609 58.5702
R1715 B.n607 B.n606 58.5702
R1716 B.n853 B.n541 57.2896
R1717 B.n1122 B.n1121 57.2896
R1718 B.n860 B.n541 33.2967
R1719 B.n860 B.n537 33.2967
R1720 B.n866 B.n537 33.2967
R1721 B.n866 B.n533 33.2967
R1722 B.n872 B.n533 33.2967
R1723 B.n872 B.n529 33.2967
R1724 B.n878 B.n529 33.2967
R1725 B.n884 B.n525 33.2967
R1726 B.n884 B.n521 33.2967
R1727 B.n890 B.n521 33.2967
R1728 B.n890 B.n517 33.2967
R1729 B.n896 B.n517 33.2967
R1730 B.n896 B.n513 33.2967
R1731 B.n902 B.n513 33.2967
R1732 B.n902 B.n509 33.2967
R1733 B.n908 B.n509 33.2967
R1734 B.n908 B.n505 33.2967
R1735 B.n914 B.n505 33.2967
R1736 B.n920 B.n501 33.2967
R1737 B.n920 B.n497 33.2967
R1738 B.n926 B.n497 33.2967
R1739 B.n926 B.n493 33.2967
R1740 B.n932 B.n493 33.2967
R1741 B.n932 B.n488 33.2967
R1742 B.n938 B.n488 33.2967
R1743 B.n938 B.n489 33.2967
R1744 B.n944 B.n481 33.2967
R1745 B.n950 B.n481 33.2967
R1746 B.n950 B.n477 33.2967
R1747 B.n956 B.n477 33.2967
R1748 B.n956 B.n473 33.2967
R1749 B.n962 B.n473 33.2967
R1750 B.n962 B.n469 33.2967
R1751 B.n968 B.n469 33.2967
R1752 B.n974 B.n465 33.2967
R1753 B.n974 B.n461 33.2967
R1754 B.n980 B.n461 33.2967
R1755 B.n980 B.n457 33.2967
R1756 B.n986 B.n457 33.2967
R1757 B.n986 B.n453 33.2967
R1758 B.n993 B.n453 33.2967
R1759 B.n993 B.n992 33.2967
R1760 B.n999 B.n446 33.2967
R1761 B.n1005 B.n446 33.2967
R1762 B.n1005 B.n442 33.2967
R1763 B.n1011 B.n442 33.2967
R1764 B.n1011 B.n438 33.2967
R1765 B.n1017 B.n438 33.2967
R1766 B.n1017 B.n434 33.2967
R1767 B.n1023 B.n434 33.2967
R1768 B.n1030 B.n430 33.2967
R1769 B.n1030 B.n426 33.2967
R1770 B.n1036 B.n426 33.2967
R1771 B.n1036 B.n4 33.2967
R1772 B.n1244 B.n4 33.2967
R1773 B.n1244 B.n1243 33.2967
R1774 B.n1243 B.n1242 33.2967
R1775 B.n1242 B.n8 33.2967
R1776 B.n12 B.n8 33.2967
R1777 B.n1235 B.n12 33.2967
R1778 B.n1235 B.n1234 33.2967
R1779 B.n1233 B.n16 33.2967
R1780 B.n1227 B.n16 33.2967
R1781 B.n1227 B.n1226 33.2967
R1782 B.n1226 B.n1225 33.2967
R1783 B.n1225 B.n23 33.2967
R1784 B.n1219 B.n23 33.2967
R1785 B.n1219 B.n1218 33.2967
R1786 B.n1218 B.n1217 33.2967
R1787 B.n1211 B.n33 33.2967
R1788 B.n1211 B.n1210 33.2967
R1789 B.n1210 B.n1209 33.2967
R1790 B.n1209 B.n37 33.2967
R1791 B.n1203 B.n37 33.2967
R1792 B.n1203 B.n1202 33.2967
R1793 B.n1202 B.n1201 33.2967
R1794 B.n1201 B.n44 33.2967
R1795 B.n1195 B.n1194 33.2967
R1796 B.n1194 B.n1193 33.2967
R1797 B.n1193 B.n51 33.2967
R1798 B.n1187 B.n51 33.2967
R1799 B.n1187 B.n1186 33.2967
R1800 B.n1186 B.n1185 33.2967
R1801 B.n1185 B.n58 33.2967
R1802 B.n1179 B.n58 33.2967
R1803 B.n1178 B.n1177 33.2967
R1804 B.n1177 B.n65 33.2967
R1805 B.n1171 B.n65 33.2967
R1806 B.n1171 B.n1170 33.2967
R1807 B.n1170 B.n1169 33.2967
R1808 B.n1169 B.n72 33.2967
R1809 B.n1163 B.n72 33.2967
R1810 B.n1163 B.n1162 33.2967
R1811 B.n1161 B.n79 33.2967
R1812 B.n1155 B.n79 33.2967
R1813 B.n1155 B.n1154 33.2967
R1814 B.n1154 B.n1153 33.2967
R1815 B.n1153 B.n86 33.2967
R1816 B.n1147 B.n86 33.2967
R1817 B.n1147 B.n1146 33.2967
R1818 B.n1146 B.n1145 33.2967
R1819 B.n1145 B.n93 33.2967
R1820 B.n1139 B.n93 33.2967
R1821 B.n1139 B.n1138 33.2967
R1822 B.n1137 B.n100 33.2967
R1823 B.n1131 B.n100 33.2967
R1824 B.n1131 B.n1130 33.2967
R1825 B.n1130 B.n1129 33.2967
R1826 B.n1129 B.n107 33.2967
R1827 B.n1123 B.n107 33.2967
R1828 B.n1123 B.n1122 33.2967
R1829 B.n850 B.n539 33.2493
R1830 B.n857 B.n856 33.2493
R1831 B.n1119 B.n1118 33.2493
R1832 B.n181 B.n109 33.2493
R1833 B.n914 B.t9 30.8485
R1834 B.t7 B.n1161 30.8485
R1835 B.n878 B.t11 27.9106
R1836 B.t15 B.n1137 27.9106
R1837 B.n489 B.t1 26.9313
R1838 B.t6 B.n1178 26.9313
R1839 B.n968 B.t4 23.0141
R1840 B.n1195 B.t3 23.0141
R1841 B.n992 B.t0 19.0969
R1842 B.n33 B.t5 19.0969
R1843 B.t8 B.n430 18.1176
R1844 B.n1234 B.t2 18.1176
R1845 B B.n1247 18.0485
R1846 B.n1023 B.t8 15.1797
R1847 B.t2 B.n1233 15.1797
R1848 B.n999 B.t0 14.2004
R1849 B.n1217 B.t5 14.2004
R1850 B.n862 B.n539 10.6151
R1851 B.n863 B.n862 10.6151
R1852 B.n864 B.n863 10.6151
R1853 B.n864 B.n531 10.6151
R1854 B.n874 B.n531 10.6151
R1855 B.n875 B.n874 10.6151
R1856 B.n876 B.n875 10.6151
R1857 B.n876 B.n523 10.6151
R1858 B.n886 B.n523 10.6151
R1859 B.n887 B.n886 10.6151
R1860 B.n888 B.n887 10.6151
R1861 B.n888 B.n515 10.6151
R1862 B.n898 B.n515 10.6151
R1863 B.n899 B.n898 10.6151
R1864 B.n900 B.n899 10.6151
R1865 B.n900 B.n507 10.6151
R1866 B.n910 B.n507 10.6151
R1867 B.n911 B.n910 10.6151
R1868 B.n912 B.n911 10.6151
R1869 B.n912 B.n499 10.6151
R1870 B.n922 B.n499 10.6151
R1871 B.n923 B.n922 10.6151
R1872 B.n924 B.n923 10.6151
R1873 B.n924 B.n491 10.6151
R1874 B.n934 B.n491 10.6151
R1875 B.n935 B.n934 10.6151
R1876 B.n936 B.n935 10.6151
R1877 B.n936 B.n483 10.6151
R1878 B.n946 B.n483 10.6151
R1879 B.n947 B.n946 10.6151
R1880 B.n948 B.n947 10.6151
R1881 B.n948 B.n475 10.6151
R1882 B.n958 B.n475 10.6151
R1883 B.n959 B.n958 10.6151
R1884 B.n960 B.n959 10.6151
R1885 B.n960 B.n467 10.6151
R1886 B.n970 B.n467 10.6151
R1887 B.n971 B.n970 10.6151
R1888 B.n972 B.n971 10.6151
R1889 B.n972 B.n459 10.6151
R1890 B.n982 B.n459 10.6151
R1891 B.n983 B.n982 10.6151
R1892 B.n984 B.n983 10.6151
R1893 B.n984 B.n451 10.6151
R1894 B.n995 B.n451 10.6151
R1895 B.n996 B.n995 10.6151
R1896 B.n997 B.n996 10.6151
R1897 B.n997 B.n444 10.6151
R1898 B.n1007 B.n444 10.6151
R1899 B.n1008 B.n1007 10.6151
R1900 B.n1009 B.n1008 10.6151
R1901 B.n1009 B.n436 10.6151
R1902 B.n1019 B.n436 10.6151
R1903 B.n1020 B.n1019 10.6151
R1904 B.n1021 B.n1020 10.6151
R1905 B.n1021 B.n428 10.6151
R1906 B.n1032 B.n428 10.6151
R1907 B.n1033 B.n1032 10.6151
R1908 B.n1034 B.n1033 10.6151
R1909 B.n1034 B.n0 10.6151
R1910 B.n850 B.n849 10.6151
R1911 B.n849 B.n848 10.6151
R1912 B.n848 B.n847 10.6151
R1913 B.n847 B.n845 10.6151
R1914 B.n845 B.n842 10.6151
R1915 B.n842 B.n841 10.6151
R1916 B.n841 B.n838 10.6151
R1917 B.n838 B.n837 10.6151
R1918 B.n837 B.n834 10.6151
R1919 B.n834 B.n833 10.6151
R1920 B.n833 B.n830 10.6151
R1921 B.n830 B.n829 10.6151
R1922 B.n829 B.n826 10.6151
R1923 B.n826 B.n825 10.6151
R1924 B.n825 B.n822 10.6151
R1925 B.n822 B.n821 10.6151
R1926 B.n821 B.n818 10.6151
R1927 B.n818 B.n817 10.6151
R1928 B.n817 B.n814 10.6151
R1929 B.n814 B.n813 10.6151
R1930 B.n813 B.n810 10.6151
R1931 B.n810 B.n809 10.6151
R1932 B.n809 B.n806 10.6151
R1933 B.n806 B.n805 10.6151
R1934 B.n805 B.n802 10.6151
R1935 B.n802 B.n801 10.6151
R1936 B.n801 B.n798 10.6151
R1937 B.n798 B.n797 10.6151
R1938 B.n797 B.n794 10.6151
R1939 B.n794 B.n793 10.6151
R1940 B.n793 B.n790 10.6151
R1941 B.n790 B.n789 10.6151
R1942 B.n789 B.n786 10.6151
R1943 B.n786 B.n785 10.6151
R1944 B.n785 B.n782 10.6151
R1945 B.n782 B.n781 10.6151
R1946 B.n781 B.n778 10.6151
R1947 B.n778 B.n777 10.6151
R1948 B.n777 B.n774 10.6151
R1949 B.n774 B.n773 10.6151
R1950 B.n773 B.n770 10.6151
R1951 B.n770 B.n769 10.6151
R1952 B.n769 B.n766 10.6151
R1953 B.n766 B.n765 10.6151
R1954 B.n765 B.n762 10.6151
R1955 B.n762 B.n761 10.6151
R1956 B.n761 B.n758 10.6151
R1957 B.n758 B.n757 10.6151
R1958 B.n757 B.n754 10.6151
R1959 B.n754 B.n753 10.6151
R1960 B.n753 B.n750 10.6151
R1961 B.n750 B.n749 10.6151
R1962 B.n749 B.n746 10.6151
R1963 B.n746 B.n745 10.6151
R1964 B.n745 B.n742 10.6151
R1965 B.n742 B.n741 10.6151
R1966 B.n738 B.n737 10.6151
R1967 B.n737 B.n734 10.6151
R1968 B.n734 B.n733 10.6151
R1969 B.n733 B.n730 10.6151
R1970 B.n730 B.n729 10.6151
R1971 B.n729 B.n726 10.6151
R1972 B.n726 B.n725 10.6151
R1973 B.n725 B.n722 10.6151
R1974 B.n720 B.n717 10.6151
R1975 B.n717 B.n716 10.6151
R1976 B.n716 B.n713 10.6151
R1977 B.n713 B.n712 10.6151
R1978 B.n712 B.n709 10.6151
R1979 B.n709 B.n708 10.6151
R1980 B.n708 B.n705 10.6151
R1981 B.n705 B.n704 10.6151
R1982 B.n704 B.n701 10.6151
R1983 B.n701 B.n700 10.6151
R1984 B.n700 B.n697 10.6151
R1985 B.n697 B.n696 10.6151
R1986 B.n696 B.n693 10.6151
R1987 B.n693 B.n692 10.6151
R1988 B.n692 B.n689 10.6151
R1989 B.n689 B.n688 10.6151
R1990 B.n688 B.n685 10.6151
R1991 B.n685 B.n684 10.6151
R1992 B.n684 B.n681 10.6151
R1993 B.n681 B.n680 10.6151
R1994 B.n680 B.n677 10.6151
R1995 B.n677 B.n676 10.6151
R1996 B.n676 B.n673 10.6151
R1997 B.n673 B.n672 10.6151
R1998 B.n672 B.n669 10.6151
R1999 B.n669 B.n668 10.6151
R2000 B.n668 B.n665 10.6151
R2001 B.n665 B.n664 10.6151
R2002 B.n664 B.n661 10.6151
R2003 B.n661 B.n660 10.6151
R2004 B.n660 B.n657 10.6151
R2005 B.n657 B.n656 10.6151
R2006 B.n656 B.n653 10.6151
R2007 B.n653 B.n652 10.6151
R2008 B.n652 B.n649 10.6151
R2009 B.n649 B.n648 10.6151
R2010 B.n648 B.n645 10.6151
R2011 B.n645 B.n644 10.6151
R2012 B.n644 B.n641 10.6151
R2013 B.n641 B.n640 10.6151
R2014 B.n640 B.n637 10.6151
R2015 B.n637 B.n636 10.6151
R2016 B.n636 B.n633 10.6151
R2017 B.n633 B.n632 10.6151
R2018 B.n632 B.n629 10.6151
R2019 B.n629 B.n628 10.6151
R2020 B.n628 B.n625 10.6151
R2021 B.n625 B.n624 10.6151
R2022 B.n624 B.n621 10.6151
R2023 B.n621 B.n620 10.6151
R2024 B.n620 B.n617 10.6151
R2025 B.n617 B.n616 10.6151
R2026 B.n616 B.n613 10.6151
R2027 B.n613 B.n612 10.6151
R2028 B.n612 B.n543 10.6151
R2029 B.n856 B.n543 10.6151
R2030 B.n858 B.n857 10.6151
R2031 B.n858 B.n535 10.6151
R2032 B.n868 B.n535 10.6151
R2033 B.n869 B.n868 10.6151
R2034 B.n870 B.n869 10.6151
R2035 B.n870 B.n527 10.6151
R2036 B.n880 B.n527 10.6151
R2037 B.n881 B.n880 10.6151
R2038 B.n882 B.n881 10.6151
R2039 B.n882 B.n519 10.6151
R2040 B.n892 B.n519 10.6151
R2041 B.n893 B.n892 10.6151
R2042 B.n894 B.n893 10.6151
R2043 B.n894 B.n511 10.6151
R2044 B.n904 B.n511 10.6151
R2045 B.n905 B.n904 10.6151
R2046 B.n906 B.n905 10.6151
R2047 B.n906 B.n503 10.6151
R2048 B.n916 B.n503 10.6151
R2049 B.n917 B.n916 10.6151
R2050 B.n918 B.n917 10.6151
R2051 B.n918 B.n495 10.6151
R2052 B.n928 B.n495 10.6151
R2053 B.n929 B.n928 10.6151
R2054 B.n930 B.n929 10.6151
R2055 B.n930 B.n486 10.6151
R2056 B.n940 B.n486 10.6151
R2057 B.n941 B.n940 10.6151
R2058 B.n942 B.n941 10.6151
R2059 B.n942 B.n479 10.6151
R2060 B.n952 B.n479 10.6151
R2061 B.n953 B.n952 10.6151
R2062 B.n954 B.n953 10.6151
R2063 B.n954 B.n471 10.6151
R2064 B.n964 B.n471 10.6151
R2065 B.n965 B.n964 10.6151
R2066 B.n966 B.n965 10.6151
R2067 B.n966 B.n463 10.6151
R2068 B.n976 B.n463 10.6151
R2069 B.n977 B.n976 10.6151
R2070 B.n978 B.n977 10.6151
R2071 B.n978 B.n455 10.6151
R2072 B.n988 B.n455 10.6151
R2073 B.n989 B.n988 10.6151
R2074 B.n990 B.n989 10.6151
R2075 B.n990 B.n448 10.6151
R2076 B.n1001 B.n448 10.6151
R2077 B.n1002 B.n1001 10.6151
R2078 B.n1003 B.n1002 10.6151
R2079 B.n1003 B.n440 10.6151
R2080 B.n1013 B.n440 10.6151
R2081 B.n1014 B.n1013 10.6151
R2082 B.n1015 B.n1014 10.6151
R2083 B.n1015 B.n432 10.6151
R2084 B.n1025 B.n432 10.6151
R2085 B.n1026 B.n1025 10.6151
R2086 B.n1028 B.n1026 10.6151
R2087 B.n1028 B.n1027 10.6151
R2088 B.n1027 B.n424 10.6151
R2089 B.n1039 B.n424 10.6151
R2090 B.n1040 B.n1039 10.6151
R2091 B.n1041 B.n1040 10.6151
R2092 B.n1042 B.n1041 10.6151
R2093 B.n1043 B.n1042 10.6151
R2094 B.n1046 B.n1043 10.6151
R2095 B.n1047 B.n1046 10.6151
R2096 B.n1048 B.n1047 10.6151
R2097 B.n1049 B.n1048 10.6151
R2098 B.n1051 B.n1049 10.6151
R2099 B.n1052 B.n1051 10.6151
R2100 B.n1053 B.n1052 10.6151
R2101 B.n1054 B.n1053 10.6151
R2102 B.n1056 B.n1054 10.6151
R2103 B.n1057 B.n1056 10.6151
R2104 B.n1058 B.n1057 10.6151
R2105 B.n1059 B.n1058 10.6151
R2106 B.n1061 B.n1059 10.6151
R2107 B.n1062 B.n1061 10.6151
R2108 B.n1063 B.n1062 10.6151
R2109 B.n1064 B.n1063 10.6151
R2110 B.n1066 B.n1064 10.6151
R2111 B.n1067 B.n1066 10.6151
R2112 B.n1068 B.n1067 10.6151
R2113 B.n1069 B.n1068 10.6151
R2114 B.n1071 B.n1069 10.6151
R2115 B.n1072 B.n1071 10.6151
R2116 B.n1073 B.n1072 10.6151
R2117 B.n1074 B.n1073 10.6151
R2118 B.n1076 B.n1074 10.6151
R2119 B.n1077 B.n1076 10.6151
R2120 B.n1078 B.n1077 10.6151
R2121 B.n1079 B.n1078 10.6151
R2122 B.n1081 B.n1079 10.6151
R2123 B.n1082 B.n1081 10.6151
R2124 B.n1083 B.n1082 10.6151
R2125 B.n1084 B.n1083 10.6151
R2126 B.n1086 B.n1084 10.6151
R2127 B.n1087 B.n1086 10.6151
R2128 B.n1088 B.n1087 10.6151
R2129 B.n1089 B.n1088 10.6151
R2130 B.n1091 B.n1089 10.6151
R2131 B.n1092 B.n1091 10.6151
R2132 B.n1093 B.n1092 10.6151
R2133 B.n1094 B.n1093 10.6151
R2134 B.n1096 B.n1094 10.6151
R2135 B.n1097 B.n1096 10.6151
R2136 B.n1098 B.n1097 10.6151
R2137 B.n1099 B.n1098 10.6151
R2138 B.n1101 B.n1099 10.6151
R2139 B.n1102 B.n1101 10.6151
R2140 B.n1103 B.n1102 10.6151
R2141 B.n1104 B.n1103 10.6151
R2142 B.n1106 B.n1104 10.6151
R2143 B.n1107 B.n1106 10.6151
R2144 B.n1108 B.n1107 10.6151
R2145 B.n1109 B.n1108 10.6151
R2146 B.n1111 B.n1109 10.6151
R2147 B.n1112 B.n1111 10.6151
R2148 B.n1113 B.n1112 10.6151
R2149 B.n1114 B.n1113 10.6151
R2150 B.n1116 B.n1114 10.6151
R2151 B.n1117 B.n1116 10.6151
R2152 B.n1118 B.n1117 10.6151
R2153 B.n1239 B.n1 10.6151
R2154 B.n1239 B.n1238 10.6151
R2155 B.n1238 B.n1237 10.6151
R2156 B.n1237 B.n10 10.6151
R2157 B.n1231 B.n10 10.6151
R2158 B.n1231 B.n1230 10.6151
R2159 B.n1230 B.n1229 10.6151
R2160 B.n1229 B.n18 10.6151
R2161 B.n1223 B.n18 10.6151
R2162 B.n1223 B.n1222 10.6151
R2163 B.n1222 B.n1221 10.6151
R2164 B.n1221 B.n25 10.6151
R2165 B.n1215 B.n25 10.6151
R2166 B.n1215 B.n1214 10.6151
R2167 B.n1214 B.n1213 10.6151
R2168 B.n1213 B.n31 10.6151
R2169 B.n1207 B.n31 10.6151
R2170 B.n1207 B.n1206 10.6151
R2171 B.n1206 B.n1205 10.6151
R2172 B.n1205 B.n39 10.6151
R2173 B.n1199 B.n39 10.6151
R2174 B.n1199 B.n1198 10.6151
R2175 B.n1198 B.n1197 10.6151
R2176 B.n1197 B.n46 10.6151
R2177 B.n1191 B.n46 10.6151
R2178 B.n1191 B.n1190 10.6151
R2179 B.n1190 B.n1189 10.6151
R2180 B.n1189 B.n53 10.6151
R2181 B.n1183 B.n53 10.6151
R2182 B.n1183 B.n1182 10.6151
R2183 B.n1182 B.n1181 10.6151
R2184 B.n1181 B.n60 10.6151
R2185 B.n1175 B.n60 10.6151
R2186 B.n1175 B.n1174 10.6151
R2187 B.n1174 B.n1173 10.6151
R2188 B.n1173 B.n67 10.6151
R2189 B.n1167 B.n67 10.6151
R2190 B.n1167 B.n1166 10.6151
R2191 B.n1166 B.n1165 10.6151
R2192 B.n1165 B.n74 10.6151
R2193 B.n1159 B.n74 10.6151
R2194 B.n1159 B.n1158 10.6151
R2195 B.n1158 B.n1157 10.6151
R2196 B.n1157 B.n81 10.6151
R2197 B.n1151 B.n81 10.6151
R2198 B.n1151 B.n1150 10.6151
R2199 B.n1150 B.n1149 10.6151
R2200 B.n1149 B.n88 10.6151
R2201 B.n1143 B.n88 10.6151
R2202 B.n1143 B.n1142 10.6151
R2203 B.n1142 B.n1141 10.6151
R2204 B.n1141 B.n95 10.6151
R2205 B.n1135 B.n95 10.6151
R2206 B.n1135 B.n1134 10.6151
R2207 B.n1134 B.n1133 10.6151
R2208 B.n1133 B.n102 10.6151
R2209 B.n1127 B.n102 10.6151
R2210 B.n1127 B.n1126 10.6151
R2211 B.n1126 B.n1125 10.6151
R2212 B.n1125 B.n109 10.6151
R2213 B.n182 B.n181 10.6151
R2214 B.n185 B.n182 10.6151
R2215 B.n186 B.n185 10.6151
R2216 B.n189 B.n186 10.6151
R2217 B.n190 B.n189 10.6151
R2218 B.n193 B.n190 10.6151
R2219 B.n194 B.n193 10.6151
R2220 B.n197 B.n194 10.6151
R2221 B.n198 B.n197 10.6151
R2222 B.n201 B.n198 10.6151
R2223 B.n202 B.n201 10.6151
R2224 B.n205 B.n202 10.6151
R2225 B.n206 B.n205 10.6151
R2226 B.n209 B.n206 10.6151
R2227 B.n210 B.n209 10.6151
R2228 B.n213 B.n210 10.6151
R2229 B.n214 B.n213 10.6151
R2230 B.n217 B.n214 10.6151
R2231 B.n218 B.n217 10.6151
R2232 B.n221 B.n218 10.6151
R2233 B.n222 B.n221 10.6151
R2234 B.n225 B.n222 10.6151
R2235 B.n226 B.n225 10.6151
R2236 B.n229 B.n226 10.6151
R2237 B.n230 B.n229 10.6151
R2238 B.n233 B.n230 10.6151
R2239 B.n234 B.n233 10.6151
R2240 B.n237 B.n234 10.6151
R2241 B.n238 B.n237 10.6151
R2242 B.n241 B.n238 10.6151
R2243 B.n242 B.n241 10.6151
R2244 B.n245 B.n242 10.6151
R2245 B.n246 B.n245 10.6151
R2246 B.n249 B.n246 10.6151
R2247 B.n250 B.n249 10.6151
R2248 B.n253 B.n250 10.6151
R2249 B.n254 B.n253 10.6151
R2250 B.n257 B.n254 10.6151
R2251 B.n258 B.n257 10.6151
R2252 B.n261 B.n258 10.6151
R2253 B.n262 B.n261 10.6151
R2254 B.n265 B.n262 10.6151
R2255 B.n266 B.n265 10.6151
R2256 B.n269 B.n266 10.6151
R2257 B.n270 B.n269 10.6151
R2258 B.n273 B.n270 10.6151
R2259 B.n274 B.n273 10.6151
R2260 B.n277 B.n274 10.6151
R2261 B.n278 B.n277 10.6151
R2262 B.n281 B.n278 10.6151
R2263 B.n282 B.n281 10.6151
R2264 B.n285 B.n282 10.6151
R2265 B.n286 B.n285 10.6151
R2266 B.n289 B.n286 10.6151
R2267 B.n290 B.n289 10.6151
R2268 B.n293 B.n290 10.6151
R2269 B.n298 B.n295 10.6151
R2270 B.n299 B.n298 10.6151
R2271 B.n302 B.n299 10.6151
R2272 B.n303 B.n302 10.6151
R2273 B.n306 B.n303 10.6151
R2274 B.n307 B.n306 10.6151
R2275 B.n310 B.n307 10.6151
R2276 B.n311 B.n310 10.6151
R2277 B.n315 B.n314 10.6151
R2278 B.n318 B.n315 10.6151
R2279 B.n319 B.n318 10.6151
R2280 B.n322 B.n319 10.6151
R2281 B.n323 B.n322 10.6151
R2282 B.n326 B.n323 10.6151
R2283 B.n327 B.n326 10.6151
R2284 B.n330 B.n327 10.6151
R2285 B.n331 B.n330 10.6151
R2286 B.n334 B.n331 10.6151
R2287 B.n335 B.n334 10.6151
R2288 B.n338 B.n335 10.6151
R2289 B.n339 B.n338 10.6151
R2290 B.n342 B.n339 10.6151
R2291 B.n343 B.n342 10.6151
R2292 B.n346 B.n343 10.6151
R2293 B.n347 B.n346 10.6151
R2294 B.n350 B.n347 10.6151
R2295 B.n351 B.n350 10.6151
R2296 B.n354 B.n351 10.6151
R2297 B.n355 B.n354 10.6151
R2298 B.n358 B.n355 10.6151
R2299 B.n359 B.n358 10.6151
R2300 B.n362 B.n359 10.6151
R2301 B.n363 B.n362 10.6151
R2302 B.n366 B.n363 10.6151
R2303 B.n367 B.n366 10.6151
R2304 B.n370 B.n367 10.6151
R2305 B.n371 B.n370 10.6151
R2306 B.n374 B.n371 10.6151
R2307 B.n375 B.n374 10.6151
R2308 B.n378 B.n375 10.6151
R2309 B.n379 B.n378 10.6151
R2310 B.n382 B.n379 10.6151
R2311 B.n383 B.n382 10.6151
R2312 B.n386 B.n383 10.6151
R2313 B.n387 B.n386 10.6151
R2314 B.n390 B.n387 10.6151
R2315 B.n391 B.n390 10.6151
R2316 B.n394 B.n391 10.6151
R2317 B.n395 B.n394 10.6151
R2318 B.n398 B.n395 10.6151
R2319 B.n399 B.n398 10.6151
R2320 B.n402 B.n399 10.6151
R2321 B.n403 B.n402 10.6151
R2322 B.n406 B.n403 10.6151
R2323 B.n407 B.n406 10.6151
R2324 B.n410 B.n407 10.6151
R2325 B.n411 B.n410 10.6151
R2326 B.n414 B.n411 10.6151
R2327 B.n415 B.n414 10.6151
R2328 B.n418 B.n415 10.6151
R2329 B.n419 B.n418 10.6151
R2330 B.n422 B.n419 10.6151
R2331 B.n423 B.n422 10.6151
R2332 B.n1119 B.n423 10.6151
R2333 B.t4 B.n465 10.2832
R2334 B.t3 B.n44 10.2832
R2335 B.n1247 B.n0 8.11757
R2336 B.n1247 B.n1 8.11757
R2337 B.n738 B.n608 6.5566
R2338 B.n722 B.n721 6.5566
R2339 B.n295 B.n294 6.5566
R2340 B.n311 B.n177 6.5566
R2341 B.n944 B.t1 6.36596
R2342 B.n1179 B.t6 6.36596
R2343 B.t11 B.n525 5.38666
R2344 B.n1138 B.t15 5.38666
R2345 B.n741 B.n608 4.05904
R2346 B.n721 B.n720 4.05904
R2347 B.n294 B.n293 4.05904
R2348 B.n314 B.n177 4.05904
R2349 B.t9 B.n501 2.44875
R2350 B.n1162 B.t7 2.44875
R2351 VN.n10 VN.t2 184.72
R2352 VN.n53 VN.t7 184.72
R2353 VN.n83 VN.n43 161.3
R2354 VN.n82 VN.n81 161.3
R2355 VN.n80 VN.n44 161.3
R2356 VN.n79 VN.n78 161.3
R2357 VN.n77 VN.n45 161.3
R2358 VN.n76 VN.n75 161.3
R2359 VN.n74 VN.n73 161.3
R2360 VN.n72 VN.n47 161.3
R2361 VN.n71 VN.n70 161.3
R2362 VN.n69 VN.n48 161.3
R2363 VN.n68 VN.n67 161.3
R2364 VN.n66 VN.n49 161.3
R2365 VN.n65 VN.n64 161.3
R2366 VN.n63 VN.n50 161.3
R2367 VN.n62 VN.n61 161.3
R2368 VN.n60 VN.n51 161.3
R2369 VN.n59 VN.n58 161.3
R2370 VN.n57 VN.n52 161.3
R2371 VN.n56 VN.n55 161.3
R2372 VN.n40 VN.n0 161.3
R2373 VN.n39 VN.n38 161.3
R2374 VN.n37 VN.n1 161.3
R2375 VN.n36 VN.n35 161.3
R2376 VN.n34 VN.n2 161.3
R2377 VN.n33 VN.n32 161.3
R2378 VN.n31 VN.n30 161.3
R2379 VN.n29 VN.n4 161.3
R2380 VN.n28 VN.n27 161.3
R2381 VN.n26 VN.n5 161.3
R2382 VN.n25 VN.n24 161.3
R2383 VN.n23 VN.n6 161.3
R2384 VN.n22 VN.n21 161.3
R2385 VN.n20 VN.n7 161.3
R2386 VN.n19 VN.n18 161.3
R2387 VN.n17 VN.n8 161.3
R2388 VN.n16 VN.n15 161.3
R2389 VN.n14 VN.n9 161.3
R2390 VN.n13 VN.n12 161.3
R2391 VN.n22 VN.t8 154.007
R2392 VN.n11 VN.t1 154.007
R2393 VN.n3 VN.t6 154.007
R2394 VN.n41 VN.t9 154.007
R2395 VN.n65 VN.t4 154.007
R2396 VN.n54 VN.t5 154.007
R2397 VN.n46 VN.t3 154.007
R2398 VN.n84 VN.t0 154.007
R2399 VN.n42 VN.n41 108.799
R2400 VN.n85 VN.n84 108.799
R2401 VN.n11 VN.n10 72.37
R2402 VN.n54 VN.n53 72.37
R2403 VN VN.n85 57.733
R2404 VN.n35 VN.n1 43.4072
R2405 VN.n78 VN.n44 43.4072
R2406 VN.n17 VN.n16 41.4647
R2407 VN.n28 VN.n5 41.4647
R2408 VN.n60 VN.n59 41.4647
R2409 VN.n71 VN.n48 41.4647
R2410 VN.n18 VN.n17 39.5221
R2411 VN.n24 VN.n5 39.5221
R2412 VN.n61 VN.n60 39.5221
R2413 VN.n67 VN.n48 39.5221
R2414 VN.n35 VN.n34 37.5796
R2415 VN.n78 VN.n77 37.5796
R2416 VN.n12 VN.n9 24.4675
R2417 VN.n16 VN.n9 24.4675
R2418 VN.n18 VN.n7 24.4675
R2419 VN.n22 VN.n7 24.4675
R2420 VN.n23 VN.n22 24.4675
R2421 VN.n24 VN.n23 24.4675
R2422 VN.n29 VN.n28 24.4675
R2423 VN.n30 VN.n29 24.4675
R2424 VN.n34 VN.n33 24.4675
R2425 VN.n39 VN.n1 24.4675
R2426 VN.n40 VN.n39 24.4675
R2427 VN.n59 VN.n52 24.4675
R2428 VN.n55 VN.n52 24.4675
R2429 VN.n67 VN.n66 24.4675
R2430 VN.n66 VN.n65 24.4675
R2431 VN.n65 VN.n50 24.4675
R2432 VN.n61 VN.n50 24.4675
R2433 VN.n77 VN.n76 24.4675
R2434 VN.n73 VN.n72 24.4675
R2435 VN.n72 VN.n71 24.4675
R2436 VN.n83 VN.n82 24.4675
R2437 VN.n82 VN.n44 24.4675
R2438 VN.n33 VN.n3 23.4888
R2439 VN.n76 VN.n46 23.4888
R2440 VN.n56 VN.n53 7.37486
R2441 VN.n13 VN.n10 7.37486
R2442 VN.n41 VN.n40 1.95786
R2443 VN.n84 VN.n83 1.95786
R2444 VN.n12 VN.n11 0.97918
R2445 VN.n30 VN.n3 0.97918
R2446 VN.n55 VN.n54 0.97918
R2447 VN.n73 VN.n46 0.97918
R2448 VN.n85 VN.n43 0.278367
R2449 VN.n42 VN.n0 0.278367
R2450 VN.n81 VN.n43 0.189894
R2451 VN.n81 VN.n80 0.189894
R2452 VN.n80 VN.n79 0.189894
R2453 VN.n79 VN.n45 0.189894
R2454 VN.n75 VN.n45 0.189894
R2455 VN.n75 VN.n74 0.189894
R2456 VN.n74 VN.n47 0.189894
R2457 VN.n70 VN.n47 0.189894
R2458 VN.n70 VN.n69 0.189894
R2459 VN.n69 VN.n68 0.189894
R2460 VN.n68 VN.n49 0.189894
R2461 VN.n64 VN.n49 0.189894
R2462 VN.n64 VN.n63 0.189894
R2463 VN.n63 VN.n62 0.189894
R2464 VN.n62 VN.n51 0.189894
R2465 VN.n58 VN.n51 0.189894
R2466 VN.n58 VN.n57 0.189894
R2467 VN.n57 VN.n56 0.189894
R2468 VN.n14 VN.n13 0.189894
R2469 VN.n15 VN.n14 0.189894
R2470 VN.n15 VN.n8 0.189894
R2471 VN.n19 VN.n8 0.189894
R2472 VN.n20 VN.n19 0.189894
R2473 VN.n21 VN.n20 0.189894
R2474 VN.n21 VN.n6 0.189894
R2475 VN.n25 VN.n6 0.189894
R2476 VN.n26 VN.n25 0.189894
R2477 VN.n27 VN.n26 0.189894
R2478 VN.n27 VN.n4 0.189894
R2479 VN.n31 VN.n4 0.189894
R2480 VN.n32 VN.n31 0.189894
R2481 VN.n32 VN.n2 0.189894
R2482 VN.n36 VN.n2 0.189894
R2483 VN.n37 VN.n36 0.189894
R2484 VN.n38 VN.n37 0.189894
R2485 VN.n38 VN.n0 0.189894
R2486 VN VN.n42 0.153454
R2487 VDD2.n1 VDD2.t7 65.039
R2488 VDD2.n3 VDD2.n2 63.1809
R2489 VDD2 VDD2.n7 63.1781
R2490 VDD2.n4 VDD2.t9 62.4357
R2491 VDD2.n6 VDD2.n5 61.2839
R2492 VDD2.n1 VDD2.n0 61.2836
R2493 VDD2.n4 VDD2.n3 50.9006
R2494 VDD2.n6 VDD2.n4 2.60395
R2495 VDD2.n7 VDD2.t4 1.15233
R2496 VDD2.n7 VDD2.t2 1.15233
R2497 VDD2.n5 VDD2.t6 1.15233
R2498 VDD2.n5 VDD2.t5 1.15233
R2499 VDD2.n2 VDD2.t3 1.15233
R2500 VDD2.n2 VDD2.t0 1.15233
R2501 VDD2.n0 VDD2.t8 1.15233
R2502 VDD2.n0 VDD2.t1 1.15233
R2503 VDD2 VDD2.n6 0.709552
R2504 VDD2.n3 VDD2.n1 0.596016
C0 VTAIL VDD2 12.818f
C1 VP VDD2 0.595093f
C2 VN VDD2 15.1698f
C3 VTAIL VP 15.629f
C4 VDD1 VDD2 2.23098f
C5 VTAIL VN 15.6146f
C6 VP VN 9.49509f
C7 VTAIL VDD1 12.767501f
C8 VDD1 VP 15.6069f
C9 VDD1 VN 0.153196f
C10 VDD2 B 8.220441f
C11 VDD1 B 8.198223f
C12 VTAIL B 10.332709f
C13 VN B 19.00395f
C14 VP B 17.462124f
C15 VDD2.t7 B 3.7391f
C16 VDD2.t8 B 0.320118f
C17 VDD2.t1 B 0.320118f
C18 VDD2.n0 B 2.91133f
C19 VDD2.n1 B 0.885492f
C20 VDD2.t3 B 0.320118f
C21 VDD2.t0 B 0.320118f
C22 VDD2.n2 B 2.92773f
C23 VDD2.n3 B 3.08939f
C24 VDD2.t9 B 3.72048f
C25 VDD2.n4 B 3.35342f
C26 VDD2.t6 B 0.320118f
C27 VDD2.t5 B 0.320118f
C28 VDD2.n5 B 2.91133f
C29 VDD2.n6 B 0.446133f
C30 VDD2.t4 B 0.320118f
C31 VDD2.t2 B 0.320118f
C32 VDD2.n7 B 2.92768f
C33 VN.n0 B 0.026604f
C34 VN.t9 B 2.56425f
C35 VN.n1 B 0.039389f
C36 VN.n2 B 0.020179f
C37 VN.t6 B 2.56425f
C38 VN.n3 B 0.89022f
C39 VN.n4 B 0.020179f
C40 VN.n5 B 0.016339f
C41 VN.n6 B 0.020179f
C42 VN.t8 B 2.56425f
C43 VN.n7 B 0.037608f
C44 VN.n8 B 0.020179f
C45 VN.n9 B 0.037608f
C46 VN.t2 B 2.73307f
C47 VN.n10 B 0.932587f
C48 VN.t1 B 2.56425f
C49 VN.n11 B 0.942788f
C50 VN.n12 B 0.019784f
C51 VN.n13 B 0.196497f
C52 VN.n14 B 0.020179f
C53 VN.n15 B 0.020179f
C54 VN.n16 B 0.03989f
C55 VN.n17 B 0.016339f
C56 VN.n18 B 0.040294f
C57 VN.n19 B 0.020179f
C58 VN.n20 B 0.020179f
C59 VN.n21 B 0.020179f
C60 VN.n22 B 0.909261f
C61 VN.n23 B 0.037608f
C62 VN.n24 B 0.040294f
C63 VN.n25 B 0.020179f
C64 VN.n26 B 0.020179f
C65 VN.n27 B 0.020179f
C66 VN.n28 B 0.03989f
C67 VN.n29 B 0.037608f
C68 VN.n30 B 0.019784f
C69 VN.n31 B 0.020179f
C70 VN.n32 B 0.020179f
C71 VN.n33 B 0.036866f
C72 VN.n34 B 0.040587f
C73 VN.n35 B 0.016547f
C74 VN.n36 B 0.020179f
C75 VN.n37 B 0.020179f
C76 VN.n38 B 0.020179f
C77 VN.n39 B 0.037608f
C78 VN.n40 B 0.020526f
C79 VN.n41 B 0.951673f
C80 VN.n42 B 0.03711f
C81 VN.n43 B 0.026604f
C82 VN.t0 B 2.56425f
C83 VN.n44 B 0.039389f
C84 VN.n45 B 0.020179f
C85 VN.t3 B 2.56425f
C86 VN.n46 B 0.89022f
C87 VN.n47 B 0.020179f
C88 VN.n48 B 0.016339f
C89 VN.n49 B 0.020179f
C90 VN.t4 B 2.56425f
C91 VN.n50 B 0.037608f
C92 VN.n51 B 0.020179f
C93 VN.n52 B 0.037608f
C94 VN.t7 B 2.73307f
C95 VN.n53 B 0.932587f
C96 VN.t5 B 2.56425f
C97 VN.n54 B 0.942788f
C98 VN.n55 B 0.019784f
C99 VN.n56 B 0.196497f
C100 VN.n57 B 0.020179f
C101 VN.n58 B 0.020179f
C102 VN.n59 B 0.03989f
C103 VN.n60 B 0.016339f
C104 VN.n61 B 0.040294f
C105 VN.n62 B 0.020179f
C106 VN.n63 B 0.020179f
C107 VN.n64 B 0.020179f
C108 VN.n65 B 0.909261f
C109 VN.n66 B 0.037608f
C110 VN.n67 B 0.040294f
C111 VN.n68 B 0.020179f
C112 VN.n69 B 0.020179f
C113 VN.n70 B 0.020179f
C114 VN.n71 B 0.03989f
C115 VN.n72 B 0.037608f
C116 VN.n73 B 0.019784f
C117 VN.n74 B 0.020179f
C118 VN.n75 B 0.020179f
C119 VN.n76 B 0.036866f
C120 VN.n77 B 0.040587f
C121 VN.n78 B 0.016547f
C122 VN.n79 B 0.020179f
C123 VN.n80 B 0.020179f
C124 VN.n81 B 0.020179f
C125 VN.n82 B 0.037608f
C126 VN.n83 B 0.020526f
C127 VN.n84 B 0.951673f
C128 VN.n85 B 1.38282f
C129 VTAIL.t2 B 0.32371f
C130 VTAIL.t5 B 0.32371f
C131 VTAIL.n0 B 2.87211f
C132 VTAIL.n1 B 0.526716f
C133 VTAIL.t11 B 3.66857f
C134 VTAIL.n2 B 0.658609f
C135 VTAIL.t9 B 0.32371f
C136 VTAIL.t8 B 0.32371f
C137 VTAIL.n3 B 2.87211f
C138 VTAIL.n4 B 0.636103f
C139 VTAIL.t15 B 0.32371f
C140 VTAIL.t17 B 0.32371f
C141 VTAIL.n5 B 2.87211f
C142 VTAIL.n6 B 2.29761f
C143 VTAIL.t19 B 0.32371f
C144 VTAIL.t1 B 0.32371f
C145 VTAIL.n7 B 2.87212f
C146 VTAIL.n8 B 2.2976f
C147 VTAIL.t4 B 0.32371f
C148 VTAIL.t0 B 0.32371f
C149 VTAIL.n9 B 2.87212f
C150 VTAIL.n10 B 0.636099f
C151 VTAIL.t18 B 3.66859f
C152 VTAIL.n11 B 0.658587f
C153 VTAIL.t12 B 0.32371f
C154 VTAIL.t13 B 0.32371f
C155 VTAIL.n12 B 2.87212f
C156 VTAIL.n13 B 0.572221f
C157 VTAIL.t14 B 0.32371f
C158 VTAIL.t16 B 0.32371f
C159 VTAIL.n14 B 2.87212f
C160 VTAIL.n15 B 0.636099f
C161 VTAIL.t10 B 3.66857f
C162 VTAIL.n16 B 2.18408f
C163 VTAIL.t7 B 3.66857f
C164 VTAIL.n17 B 2.18408f
C165 VTAIL.t3 B 0.32371f
C166 VTAIL.t6 B 0.32371f
C167 VTAIL.n18 B 2.87211f
C168 VTAIL.n19 B 0.481703f
C169 VDD1.t0 B 3.77776f
C170 VDD1.t1 B 0.323426f
C171 VDD1.t6 B 0.323426f
C172 VDD1.n0 B 2.94142f
C173 VDD1.n1 B 0.902408f
C174 VDD1.t7 B 3.77774f
C175 VDD1.t3 B 0.323426f
C176 VDD1.t9 B 0.323426f
C177 VDD1.n2 B 2.94141f
C178 VDD1.n3 B 0.894642f
C179 VDD1.t8 B 0.323426f
C180 VDD1.t5 B 0.323426f
C181 VDD1.n4 B 2.95798f
C182 VDD1.n5 B 3.24578f
C183 VDD1.t2 B 0.323426f
C184 VDD1.t4 B 0.323426f
C185 VDD1.n6 B 2.94141f
C186 VDD1.n7 B 3.43232f
C187 VP.n0 B 0.026887f
C188 VP.t6 B 2.59153f
C189 VP.n1 B 0.039808f
C190 VP.n2 B 0.020394f
C191 VP.t9 B 2.59153f
C192 VP.n3 B 0.899689f
C193 VP.n4 B 0.020394f
C194 VP.n5 B 0.016512f
C195 VP.n6 B 0.020394f
C196 VP.t8 B 2.59153f
C197 VP.n7 B 0.038008f
C198 VP.n8 B 0.020394f
C199 VP.n9 B 0.038008f
C200 VP.n10 B 0.020394f
C201 VP.t0 B 2.59153f
C202 VP.n11 B 0.016723f
C203 VP.n12 B 0.020394f
C204 VP.t2 B 2.59153f
C205 VP.n13 B 0.961796f
C206 VP.n14 B 0.026887f
C207 VP.t7 B 2.59153f
C208 VP.n15 B 0.039808f
C209 VP.n16 B 0.020394f
C210 VP.t1 B 2.59153f
C211 VP.n17 B 0.899689f
C212 VP.n18 B 0.020394f
C213 VP.n19 B 0.016512f
C214 VP.n20 B 0.020394f
C215 VP.t3 B 2.59153f
C216 VP.n21 B 0.038008f
C217 VP.n22 B 0.020394f
C218 VP.n23 B 0.038008f
C219 VP.t5 B 2.76214f
C220 VP.n24 B 0.942506f
C221 VP.t4 B 2.59153f
C222 VP.n25 B 0.952816f
C223 VP.n26 B 0.019994f
C224 VP.n27 B 0.198587f
C225 VP.n28 B 0.020394f
C226 VP.n29 B 0.020394f
C227 VP.n30 B 0.040314f
C228 VP.n31 B 0.016512f
C229 VP.n32 B 0.040723f
C230 VP.n33 B 0.020394f
C231 VP.n34 B 0.020394f
C232 VP.n35 B 0.020394f
C233 VP.n36 B 0.918932f
C234 VP.n37 B 0.038008f
C235 VP.n38 B 0.040723f
C236 VP.n39 B 0.020394f
C237 VP.n40 B 0.020394f
C238 VP.n41 B 0.020394f
C239 VP.n42 B 0.040314f
C240 VP.n43 B 0.038008f
C241 VP.n44 B 0.019994f
C242 VP.n45 B 0.020394f
C243 VP.n46 B 0.020394f
C244 VP.n47 B 0.037258f
C245 VP.n48 B 0.041019f
C246 VP.n49 B 0.016723f
C247 VP.n50 B 0.020394f
C248 VP.n51 B 0.020394f
C249 VP.n52 B 0.020394f
C250 VP.n53 B 0.038008f
C251 VP.n54 B 0.020745f
C252 VP.n55 B 0.961796f
C253 VP.n56 B 1.38679f
C254 VP.n57 B 1.39955f
C255 VP.n58 B 0.026887f
C256 VP.n59 B 0.020745f
C257 VP.n60 B 0.038008f
C258 VP.n61 B 0.039808f
C259 VP.n62 B 0.020394f
C260 VP.n63 B 0.020394f
C261 VP.n64 B 0.020394f
C262 VP.n65 B 0.041019f
C263 VP.n66 B 0.037258f
C264 VP.n67 B 0.899689f
C265 VP.n68 B 0.019994f
C266 VP.n69 B 0.020394f
C267 VP.n70 B 0.020394f
C268 VP.n71 B 0.020394f
C269 VP.n72 B 0.040314f
C270 VP.n73 B 0.016512f
C271 VP.n74 B 0.040723f
C272 VP.n75 B 0.020394f
C273 VP.n76 B 0.020394f
C274 VP.n77 B 0.020394f
C275 VP.n78 B 0.918932f
C276 VP.n79 B 0.038008f
C277 VP.n80 B 0.040723f
C278 VP.n81 B 0.020394f
C279 VP.n82 B 0.020394f
C280 VP.n83 B 0.020394f
C281 VP.n84 B 0.040314f
C282 VP.n85 B 0.038008f
C283 VP.n86 B 0.019994f
C284 VP.n87 B 0.020394f
C285 VP.n88 B 0.020394f
C286 VP.n89 B 0.037258f
C287 VP.n90 B 0.041019f
C288 VP.n91 B 0.016723f
C289 VP.n92 B 0.020394f
C290 VP.n93 B 0.020394f
C291 VP.n94 B 0.020394f
C292 VP.n95 B 0.038008f
C293 VP.n96 B 0.020745f
C294 VP.n97 B 0.961796f
C295 VP.n98 B 0.037505f
.ends

