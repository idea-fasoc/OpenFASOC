* NGSPICE file created from tg_sample_0004.ext - technology: sky130A

.subckt tg_sample_0004 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t1 VGP.t0 VIN.t1 VCC.t8 sky130_fd_pr__pfet_01v8 ad=1.17 pd=6.78 as=1.17 ps=6.78 w=3 l=0.5
X1 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X2 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=0.5
X3 VOUT.t0 VGN.t0 VIN.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.585 ps=3.78 w=1.5 l=0.5
X4 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.5
X5 VSS.t3 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=0.5
R0 VGP VGP.t0 384.51
R1 VIN VIN.t1 142.843
R2 VIN VIN.t0 114.448
R3 VOUT VOUT.t1 148.275
R4 VOUT VOUT.t0 141.881
R5 VCC.n148 VCC.n9 365.854
R6 VCC.n146 VCC.n13 365.854
R7 VCC.n73 VCC.n72 365.854
R8 VCC.n68 VCC.n28 365.854
R9 VCC.n112 VCC.t4 351.009
R10 VCC.n41 VCC.t0 351.009
R11 VCC.n146 VCC.n145 185
R12 VCC.n147 VCC.n146 185
R13 VCC.n14 VCC.n12 185
R14 VCC.n12 VCC.n10 185
R15 VCC.n103 VCC.n102 185
R16 VCC.n102 VCC.n101 185
R17 VCC.n17 VCC.n16 185
R18 VCC.n99 VCC.n17 185
R19 VCC.n97 VCC.n96 185
R20 VCC.n98 VCC.n97 185
R21 VCC.n19 VCC.n18 185
R22 VCC.n18 VCC.t8 185
R23 VCC.n92 VCC.n91 185
R24 VCC.n91 VCC.n90 185
R25 VCC.n22 VCC.n21 185
R26 VCC.n23 VCC.n22 185
R27 VCC.n79 VCC.n78 185
R28 VCC.n80 VCC.n79 185
R29 VCC.n31 VCC.n30 185
R30 VCC.n81 VCC.n30 185
R31 VCC.n74 VCC.n73 185
R32 VCC.n73 VCC.n29 185
R33 VCC.n28 VCC.n27 185
R34 VCC.n29 VCC.n28 185
R35 VCC.n83 VCC.n82 185
R36 VCC.n82 VCC.n81 185
R37 VCC.n25 VCC.n24 185
R38 VCC.n80 VCC.n24 185
R39 VCC.n88 VCC.n87 185
R40 VCC.n88 VCC.n23 185
R41 VCC.n89 VCC.n2 185
R42 VCC.n90 VCC.n89 185
R43 VCC.n156 VCC.n3 185
R44 VCC.t8 VCC.n3 185
R45 VCC.n155 VCC.n4 185
R46 VCC.n98 VCC.n4 185
R47 VCC.n154 VCC.n5 185
R48 VCC.n99 VCC.n5 185
R49 VCC.n100 VCC.n6 185
R50 VCC.n101 VCC.n100 185
R51 VCC.n150 VCC.n8 185
R52 VCC.n10 VCC.n8 185
R53 VCC.n149 VCC.n148 185
R54 VCC.n148 VCC.n147 185
R55 VCC.n143 VCC.n13 185
R56 VCC.n142 VCC.n141 185
R57 VCC.n139 VCC.n106 185
R58 VCC.n137 VCC.n136 185
R59 VCC.n135 VCC.n107 185
R60 VCC.n134 VCC.n133 185
R61 VCC.n131 VCC.n108 185
R62 VCC.n129 VCC.n128 185
R63 VCC.n127 VCC.n109 185
R64 VCC.n126 VCC.n125 185
R65 VCC.n123 VCC.n110 185
R66 VCC.n121 VCC.n120 185
R67 VCC.n119 VCC.n111 185
R68 VCC.n117 VCC.n116 185
R69 VCC.n114 VCC.n9 185
R70 VCC.n11 VCC.n9 185
R71 VCC.n68 VCC.n67 185
R72 VCC.n66 VCC.n40 185
R73 VCC.n64 VCC.n39 185
R74 VCC.n70 VCC.n39 185
R75 VCC.n63 VCC.n62 185
R76 VCC.n61 VCC.n60 185
R77 VCC.n59 VCC.n58 185
R78 VCC.n57 VCC.n56 185
R79 VCC.n55 VCC.n54 185
R80 VCC.n53 VCC.n52 185
R81 VCC.n51 VCC.n50 185
R82 VCC.n49 VCC.n48 185
R83 VCC.n47 VCC.n46 185
R84 VCC.n45 VCC.n44 185
R85 VCC.n43 VCC.n33 185
R86 VCC.n72 VCC.n32 185
R87 VCC.n112 VCC.t6 161.32
R88 VCC.n41 VCC.t3 161.32
R89 VCC.n73 VCC.n30 146.341
R90 VCC.n79 VCC.n30 146.341
R91 VCC.n79 VCC.n22 146.341
R92 VCC.n91 VCC.n22 146.341
R93 VCC.n91 VCC.n18 146.341
R94 VCC.n97 VCC.n18 146.341
R95 VCC.n97 VCC.n17 146.341
R96 VCC.n102 VCC.n17 146.341
R97 VCC.n102 VCC.n12 146.341
R98 VCC.n146 VCC.n12 146.341
R99 VCC.n82 VCC.n28 146.341
R100 VCC.n82 VCC.n24 146.341
R101 VCC.n88 VCC.n24 146.341
R102 VCC.n89 VCC.n88 146.341
R103 VCC.n89 VCC.n3 146.341
R104 VCC.n4 VCC.n3 146.341
R105 VCC.n5 VCC.n4 146.341
R106 VCC.n100 VCC.n5 146.341
R107 VCC.n100 VCC.n8 146.341
R108 VCC.n148 VCC.n8 146.341
R109 VCC.n113 VCC.t7 145.222
R110 VCC.n42 VCC.t2 145.222
R111 VCC.n70 VCC.n29 106.225
R112 VCC.n147 VCC.n11 106.225
R113 VCC.n116 VCC.n9 99.5127
R114 VCC.n121 VCC.n111 99.5127
R115 VCC.n125 VCC.n123 99.5127
R116 VCC.n129 VCC.n109 99.5127
R117 VCC.n133 VCC.n131 99.5127
R118 VCC.n137 VCC.n107 99.5127
R119 VCC.n141 VCC.n139 99.5127
R120 VCC.n40 VCC.n39 99.5127
R121 VCC.n62 VCC.n39 99.5127
R122 VCC.n60 VCC.n59 99.5127
R123 VCC.n56 VCC.n55 99.5127
R124 VCC.n52 VCC.n51 99.5127
R125 VCC.n48 VCC.n47 99.5127
R126 VCC.n44 VCC.n33 99.5127
R127 VCC.n140 VCC.n11 72.8958
R128 VCC.n138 VCC.n11 72.8958
R129 VCC.n132 VCC.n11 72.8958
R130 VCC.n130 VCC.n11 72.8958
R131 VCC.n124 VCC.n11 72.8958
R132 VCC.n122 VCC.n11 72.8958
R133 VCC.n115 VCC.n11 72.8958
R134 VCC.n70 VCC.n69 72.8958
R135 VCC.n70 VCC.n34 72.8958
R136 VCC.n70 VCC.n35 72.8958
R137 VCC.n70 VCC.n36 72.8958
R138 VCC.n70 VCC.n37 72.8958
R139 VCC.n70 VCC.n38 72.8958
R140 VCC.n71 VCC.n70 72.8958
R141 VCC.n81 VCC.n29 66.8078
R142 VCC.n80 VCC.n23 66.8078
R143 VCC.n90 VCC.n23 66.8078
R144 VCC.n90 VCC.t8 66.8078
R145 VCC.n98 VCC.t8 66.8078
R146 VCC.n99 VCC.n98 66.8078
R147 VCC.n101 VCC.n99 66.8078
R148 VCC.n147 VCC.n10 66.8078
R149 VCC.t1 VCC.n80 56.1186
R150 VCC.n101 VCC.t5 56.1186
R151 VCC.n115 VCC.n111 39.2114
R152 VCC.n123 VCC.n122 39.2114
R153 VCC.n124 VCC.n109 39.2114
R154 VCC.n131 VCC.n130 39.2114
R155 VCC.n132 VCC.n107 39.2114
R156 VCC.n139 VCC.n138 39.2114
R157 VCC.n140 VCC.n13 39.2114
R158 VCC.n69 VCC.n68 39.2114
R159 VCC.n62 VCC.n34 39.2114
R160 VCC.n59 VCC.n35 39.2114
R161 VCC.n55 VCC.n36 39.2114
R162 VCC.n51 VCC.n37 39.2114
R163 VCC.n47 VCC.n38 39.2114
R164 VCC.n71 VCC.n33 39.2114
R165 VCC.n141 VCC.n140 39.2114
R166 VCC.n138 VCC.n137 39.2114
R167 VCC.n133 VCC.n132 39.2114
R168 VCC.n130 VCC.n129 39.2114
R169 VCC.n125 VCC.n124 39.2114
R170 VCC.n122 VCC.n121 39.2114
R171 VCC.n116 VCC.n115 39.2114
R172 VCC.n69 VCC.n40 39.2114
R173 VCC.n60 VCC.n34 39.2114
R174 VCC.n56 VCC.n35 39.2114
R175 VCC.n52 VCC.n36 39.2114
R176 VCC.n48 VCC.n37 39.2114
R177 VCC.n44 VCC.n38 39.2114
R178 VCC.n72 VCC.n71 39.2114
R179 VCC.n114 VCC.n7 30.1478
R180 VCC.n144 VCC.n143 30.1478
R181 VCC.n67 VCC.n26 30.1478
R182 VCC.n75 VCC.n32 30.1478
R183 VCC.n118 VCC.n113 29.2853
R184 VCC.n65 VCC.n42 29.2853
R185 VCC.n74 VCC.n31 19.3944
R186 VCC.n78 VCC.n31 19.3944
R187 VCC.n78 VCC.n21 19.3944
R188 VCC.n92 VCC.n21 19.3944
R189 VCC.n92 VCC.n19 19.3944
R190 VCC.n96 VCC.n19 19.3944
R191 VCC.n96 VCC.n16 19.3944
R192 VCC.n103 VCC.n16 19.3944
R193 VCC.n103 VCC.n14 19.3944
R194 VCC.n145 VCC.n14 19.3944
R195 VCC.n83 VCC.n27 19.3944
R196 VCC.n83 VCC.n25 19.3944
R197 VCC.n87 VCC.n25 19.3944
R198 VCC.n87 VCC.n2 19.3944
R199 VCC.n156 VCC.n2 19.3944
R200 VCC.n156 VCC.n155 19.3944
R201 VCC.n155 VCC.n154 19.3944
R202 VCC.n154 VCC.n6 19.3944
R203 VCC.n150 VCC.n6 19.3944
R204 VCC.n150 VCC.n149 19.3944
R205 VCC.n113 VCC.n112 16.0975
R206 VCC.n42 VCC.n41 16.0975
R207 VCC.n81 VCC.t1 10.6897
R208 VCC.t5 VCC.n10 10.6897
R209 VCC.n117 VCC.n114 10.6151
R210 VCC.n120 VCC.n119 10.6151
R211 VCC.n120 VCC.n110 10.6151
R212 VCC.n126 VCC.n110 10.6151
R213 VCC.n127 VCC.n126 10.6151
R214 VCC.n128 VCC.n127 10.6151
R215 VCC.n128 VCC.n108 10.6151
R216 VCC.n134 VCC.n108 10.6151
R217 VCC.n135 VCC.n134 10.6151
R218 VCC.n136 VCC.n135 10.6151
R219 VCC.n136 VCC.n106 10.6151
R220 VCC.n142 VCC.n106 10.6151
R221 VCC.n143 VCC.n142 10.6151
R222 VCC.n67 VCC.n66 10.6151
R223 VCC.n64 VCC.n63 10.6151
R224 VCC.n63 VCC.n61 10.6151
R225 VCC.n61 VCC.n58 10.6151
R226 VCC.n58 VCC.n57 10.6151
R227 VCC.n57 VCC.n54 10.6151
R228 VCC.n54 VCC.n53 10.6151
R229 VCC.n53 VCC.n50 10.6151
R230 VCC.n50 VCC.n49 10.6151
R231 VCC.n49 VCC.n46 10.6151
R232 VCC.n46 VCC.n45 10.6151
R233 VCC.n45 VCC.n43 10.6151
R234 VCC.n43 VCC.n32 10.6151
R235 VCC.n155 VCC.n0 9.3005
R236 VCC.n154 VCC.n153 9.3005
R237 VCC.n152 VCC.n6 9.3005
R238 VCC.n151 VCC.n150 9.3005
R239 VCC.n149 VCC.n7 9.3005
R240 VCC.n76 VCC.n31 9.3005
R241 VCC.n78 VCC.n77 9.3005
R242 VCC.n21 VCC.n20 9.3005
R243 VCC.n93 VCC.n92 9.3005
R244 VCC.n94 VCC.n19 9.3005
R245 VCC.n96 VCC.n95 9.3005
R246 VCC.n16 VCC.n15 9.3005
R247 VCC.n104 VCC.n103 9.3005
R248 VCC.n105 VCC.n14 9.3005
R249 VCC.n145 VCC.n144 9.3005
R250 VCC.n75 VCC.n74 9.3005
R251 VCC.n27 VCC.n26 9.3005
R252 VCC.n84 VCC.n83 9.3005
R253 VCC.n85 VCC.n25 9.3005
R254 VCC.n87 VCC.n86 9.3005
R255 VCC.n2 VCC.n1 9.3005
R256 VCC.n157 VCC.n156 9.3005
R257 VCC.n118 VCC.n117 6.0883
R258 VCC.n66 VCC.n65 6.0883
R259 VCC.n119 VCC.n118 4.52733
R260 VCC.n65 VCC.n64 4.52733
R261 VCC.n153 VCC.n0 0.152939
R262 VCC.n153 VCC.n152 0.152939
R263 VCC.n152 VCC.n151 0.152939
R264 VCC.n151 VCC.n7 0.152939
R265 VCC.n76 VCC.n75 0.152939
R266 VCC.n77 VCC.n76 0.152939
R267 VCC.n77 VCC.n20 0.152939
R268 VCC.n93 VCC.n20 0.152939
R269 VCC.n94 VCC.n93 0.152939
R270 VCC.n95 VCC.n94 0.152939
R271 VCC.n95 VCC.n15 0.152939
R272 VCC.n104 VCC.n15 0.152939
R273 VCC.n105 VCC.n104 0.152939
R274 VCC.n144 VCC.n105 0.152939
R275 VCC.n84 VCC.n26 0.152939
R276 VCC.n85 VCC.n84 0.152939
R277 VCC.n86 VCC.n85 0.152939
R278 VCC.n86 VCC.n1 0.152939
R279 VCC.n157 VCC.n1 0.13922
R280 VCC VCC.n0 0.0767195
R281 VCC VCC.n157 0.063
R282 VGN VGN.t0 312.211
R283 VSS.n305 VSS.n74 4865.35
R284 VSS.n345 VSS.n344 4865.35
R285 VSS.n312 VSS.n74 2953.02
R286 VSS.n313 VSS.n312 2953.02
R287 VSS.n314 VSS.n313 2953.02
R288 VSS.n314 VSS.n68 2953.02
R289 VSS.n322 VSS.n68 2953.02
R290 VSS.n323 VSS.n322 2953.02
R291 VSS.n324 VSS.n323 2953.02
R292 VSS.n324 VSS.n62 2953.02
R293 VSS.n332 VSS.n62 2953.02
R294 VSS.n333 VSS.n332 2953.02
R295 VSS.n334 VSS.n333 2953.02
R296 VSS.n334 VSS.n56 2953.02
R297 VSS.n343 VSS.n56 2953.02
R298 VSS.n344 VSS.n343 2953.02
R299 VSS.n305 VSS.n304 1719.54
R300 VSS.n304 VSS.n303 1719.54
R301 VSS.n303 VSS.n79 1719.54
R302 VSS.n297 VSS.n79 1719.54
R303 VSS.n297 VSS.n296 1719.54
R304 VSS.n296 VSS.n295 1719.54
R305 VSS.n295 VSS.n83 1719.54
R306 VSS.n289 VSS.n83 1719.54
R307 VSS.n289 VSS.n288 1719.54
R308 VSS.n288 VSS.n287 1719.54
R309 VSS.n287 VSS.n87 1719.54
R310 VSS.n281 VSS.n87 1719.54
R311 VSS.n281 VSS.n280 1719.54
R312 VSS.n280 VSS.n279 1719.54
R313 VSS.n279 VSS.n91 1719.54
R314 VSS.n273 VSS.n91 1719.54
R315 VSS.n273 VSS.n272 1719.54
R316 VSS.n272 VSS.n271 1719.54
R317 VSS.n271 VSS.n95 1719.54
R318 VSS.n265 VSS.n95 1719.54
R319 VSS.n345 VSS.n52 1719.54
R320 VSS.n351 VSS.n52 1719.54
R321 VSS.n352 VSS.n351 1719.54
R322 VSS.n353 VSS.n352 1719.54
R323 VSS.n353 VSS.n48 1719.54
R324 VSS.n359 VSS.n48 1719.54
R325 VSS.n360 VSS.n359 1719.54
R326 VSS.n361 VSS.n360 1719.54
R327 VSS.n361 VSS.n44 1719.54
R328 VSS.n367 VSS.n44 1719.54
R329 VSS.n368 VSS.n367 1719.54
R330 VSS.n369 VSS.n368 1719.54
R331 VSS.n369 VSS.n40 1719.54
R332 VSS.n375 VSS.n40 1719.54
R333 VSS.n376 VSS.n375 1719.54
R334 VSS.n377 VSS.n376 1719.54
R335 VSS.n377 VSS.n36 1719.54
R336 VSS.n384 VSS.n36 1719.54
R337 VSS.n385 VSS.n384 1719.54
R338 VSS.n386 VSS.n385 1719.54
R339 VSS.n306 VSS.n75 615.024
R340 VSS.n346 VSS.n55 615.024
R341 VSS.n425 VSS.n21 615.024
R342 VSS.n262 VSS.n101 615.024
R343 VSS.n187 VSS.n153 610.22
R344 VSS.n210 VSS.n209 610.22
R345 VSS.n459 VSS.n14 610.22
R346 VSS.n461 VSS.n9 610.22
R347 VSS.n307 VSS.n306 585
R348 VSS.n306 VSS.n305 585
R349 VSS.n78 VSS.n77 585
R350 VSS.n304 VSS.n78 585
R351 VSS.n302 VSS.n301 585
R352 VSS.n303 VSS.n302 585
R353 VSS.n300 VSS.n80 585
R354 VSS.n80 VSS.n79 585
R355 VSS.n299 VSS.n298 585
R356 VSS.n298 VSS.n297 585
R357 VSS.n82 VSS.n81 585
R358 VSS.n296 VSS.n82 585
R359 VSS.n294 VSS.n293 585
R360 VSS.n295 VSS.n294 585
R361 VSS.n292 VSS.n84 585
R362 VSS.n84 VSS.n83 585
R363 VSS.n291 VSS.n290 585
R364 VSS.n290 VSS.n289 585
R365 VSS.n86 VSS.n85 585
R366 VSS.n288 VSS.n86 585
R367 VSS.n286 VSS.n285 585
R368 VSS.n287 VSS.n286 585
R369 VSS.n284 VSS.n88 585
R370 VSS.n88 VSS.n87 585
R371 VSS.n283 VSS.n282 585
R372 VSS.n282 VSS.n281 585
R373 VSS.n90 VSS.n89 585
R374 VSS.n280 VSS.n90 585
R375 VSS.n278 VSS.n277 585
R376 VSS.n279 VSS.n278 585
R377 VSS.n276 VSS.n92 585
R378 VSS.n92 VSS.n91 585
R379 VSS.n275 VSS.n274 585
R380 VSS.n274 VSS.n273 585
R381 VSS.n94 VSS.n93 585
R382 VSS.n272 VSS.n94 585
R383 VSS.n270 VSS.n269 585
R384 VSS.n271 VSS.n270 585
R385 VSS.n268 VSS.n96 585
R386 VSS.n96 VSS.n95 585
R387 VSS.n267 VSS.n266 585
R388 VSS.n266 VSS.n265 585
R389 VSS.n76 VSS.n75 585
R390 VSS.n75 VSS.n74 585
R391 VSS.n311 VSS.n310 585
R392 VSS.n312 VSS.n311 585
R393 VSS.n73 VSS.n72 585
R394 VSS.n313 VSS.n73 585
R395 VSS.n316 VSS.n315 585
R396 VSS.n315 VSS.n314 585
R397 VSS.n70 VSS.n69 585
R398 VSS.n69 VSS.n68 585
R399 VSS.n321 VSS.n320 585
R400 VSS.n322 VSS.n321 585
R401 VSS.n67 VSS.n66 585
R402 VSS.n323 VSS.n67 585
R403 VSS.n326 VSS.n325 585
R404 VSS.n325 VSS.n324 585
R405 VSS.n64 VSS.n63 585
R406 VSS.n63 VSS.n62 585
R407 VSS.n331 VSS.n330 585
R408 VSS.n332 VSS.n331 585
R409 VSS.n61 VSS.n60 585
R410 VSS.n333 VSS.n61 585
R411 VSS.n336 VSS.n335 585
R412 VSS.n335 VSS.n334 585
R413 VSS.n58 VSS.n57 585
R414 VSS.n57 VSS.n56 585
R415 VSS.n342 VSS.n341 585
R416 VSS.n343 VSS.n342 585
R417 VSS.n340 VSS.n55 585
R418 VSS.n344 VSS.n55 585
R419 VSS.n387 VSS.n34 585
R420 VSS.n387 VSS.n386 585
R421 VSS.n381 VSS.n35 585
R422 VSS.n385 VSS.n35 585
R423 VSS.n383 VSS.n382 585
R424 VSS.n384 VSS.n383 585
R425 VSS.n380 VSS.n37 585
R426 VSS.n37 VSS.n36 585
R427 VSS.n379 VSS.n378 585
R428 VSS.n378 VSS.n377 585
R429 VSS.n39 VSS.n38 585
R430 VSS.n376 VSS.n39 585
R431 VSS.n374 VSS.n373 585
R432 VSS.n375 VSS.n374 585
R433 VSS.n372 VSS.n41 585
R434 VSS.n41 VSS.n40 585
R435 VSS.n371 VSS.n370 585
R436 VSS.n370 VSS.n369 585
R437 VSS.n43 VSS.n42 585
R438 VSS.n368 VSS.n43 585
R439 VSS.n366 VSS.n365 585
R440 VSS.n367 VSS.n366 585
R441 VSS.n364 VSS.n45 585
R442 VSS.n45 VSS.n44 585
R443 VSS.n363 VSS.n362 585
R444 VSS.n362 VSS.n361 585
R445 VSS.n47 VSS.n46 585
R446 VSS.n360 VSS.n47 585
R447 VSS.n358 VSS.n357 585
R448 VSS.n359 VSS.n358 585
R449 VSS.n356 VSS.n49 585
R450 VSS.n49 VSS.n48 585
R451 VSS.n355 VSS.n354 585
R452 VSS.n354 VSS.n353 585
R453 VSS.n51 VSS.n50 585
R454 VSS.n352 VSS.n51 585
R455 VSS.n350 VSS.n349 585
R456 VSS.n351 VSS.n350 585
R457 VSS.n348 VSS.n53 585
R458 VSS.n53 VSS.n52 585
R459 VSS.n347 VSS.n346 585
R460 VSS.n346 VSS.n345 585
R461 VSS.n98 VSS.n97 585
R462 VSS.n113 VSS.n111 585
R463 VSS.n114 VSS.n110 585
R464 VSS.n114 VSS.n99 585
R465 VSS.n117 VSS.n116 585
R466 VSS.n118 VSS.n109 585
R467 VSS.n120 VSS.n119 585
R468 VSS.n122 VSS.n108 585
R469 VSS.n125 VSS.n124 585
R470 VSS.n126 VSS.n107 585
R471 VSS.n128 VSS.n127 585
R472 VSS.n130 VSS.n106 585
R473 VSS.n133 VSS.n132 585
R474 VSS.n134 VSS.n105 585
R475 VSS.n136 VSS.n135 585
R476 VSS.n138 VSS.n104 585
R477 VSS.n139 VSS.n103 585
R478 VSS.n142 VSS.n141 585
R479 VSS.n143 VSS.n101 585
R480 VSS.n101 VSS.n99 585
R481 VSS.n422 VSS.n21 585
R482 VSS.n421 VSS.n420 585
R483 VSS.n25 VSS.n24 585
R484 VSS.n416 VSS.n415 585
R485 VSS.n414 VSS.n33 585
R486 VSS.n413 VSS.n412 585
R487 VSS.n411 VSS.n410 585
R488 VSS.n409 VSS.n408 585
R489 VSS.n407 VSS.n406 585
R490 VSS.n405 VSS.n404 585
R491 VSS.n403 VSS.n402 585
R492 VSS.n401 VSS.n400 585
R493 VSS.n399 VSS.n398 585
R494 VSS.n397 VSS.n396 585
R495 VSS.n395 VSS.n394 585
R496 VSS.n393 VSS.n392 585
R497 VSS.n391 VSS.n390 585
R498 VSS.n389 VSS.n388 585
R499 VSS.n425 VSS.n424 585
R500 VSS.n426 VSS.n425 585
R501 VSS.n22 VSS.n20 585
R502 VSS.n20 VSS.n11 585
R503 VSS.n235 VSS.n12 585
R504 VSS.n460 VSS.n12 585
R505 VSS.n236 VSS.n168 585
R506 VSS.n168 VSS.n10 585
R507 VSS.n238 VSS.n237 585
R508 VSS.n239 VSS.n238 585
R509 VSS.n169 VSS.n167 585
R510 VSS.n167 VSS.n165 585
R511 VSS.n229 VSS.n228 585
R512 VSS.n228 VSS.n227 585
R513 VSS.n172 VSS.n171 585
R514 VSS.t8 VSS.n172 585
R515 VSS.n224 VSS.n223 585
R516 VSS.n225 VSS.n224 585
R517 VSS.n220 VSS.n219 585
R518 VSS.n219 VSS.n173 585
R519 VSS.n149 VSS.n147 585
R520 VSS.n174 VSS.n149 585
R521 VSS.n256 VSS.n255 585
R522 VSS.n255 VSS.n254 585
R523 VSS.n148 VSS.n145 585
R524 VSS.n151 VSS.n148 585
R525 VSS.n260 VSS.n102 585
R526 VSS.n150 VSS.n102 585
R527 VSS.n262 VSS.n261 585
R528 VSS.n263 VSS.n262 585
R529 VSS.n459 VSS.n458 585
R530 VSS.n460 VSS.n459 585
R531 VSS.n15 VSS.n13 585
R532 VSS.n13 VSS.n10 585
R533 VSS.n241 VSS.n240 585
R534 VSS.n240 VSS.n239 585
R535 VSS.n242 VSS.n164 585
R536 VSS.n165 VSS.n164 585
R537 VSS.n226 VSS.n162 585
R538 VSS.n227 VSS.n226 585
R539 VSS.n246 VSS.n161 585
R540 VSS.t8 VSS.n161 585
R541 VSS.n247 VSS.n160 585
R542 VSS.n225 VSS.n160 585
R543 VSS.n248 VSS.n159 585
R544 VSS.n173 VSS.n159 585
R545 VSS.n156 VSS.n154 585
R546 VSS.n174 VSS.n154 585
R547 VSS.n253 VSS.n252 585
R548 VSS.n254 VSS.n253 585
R549 VSS.n155 VSS.n153 585
R550 VSS.n153 VSS.n151 585
R551 VSS.n462 VSS.n461 585
R552 VSS.n461 VSS.n460 585
R553 VSS.n463 VSS.n8 585
R554 VSS.n10 VSS.n8 585
R555 VSS.n166 VSS.n6 585
R556 VSS.n239 VSS.n166 585
R557 VSS.n467 VSS.n5 585
R558 VSS.n165 VSS.n5 585
R559 VSS.n468 VSS.n4 585
R560 VSS.n227 VSS.n4 585
R561 VSS.n469 VSS.n3 585
R562 VSS.t8 VSS.n3 585
R563 VSS.n218 VSS.n2 585
R564 VSS.n225 VSS.n218 585
R565 VSS.n217 VSS.n216 585
R566 VSS.n217 VSS.n173 585
R567 VSS.n176 VSS.n175 585
R568 VSS.n175 VSS.n174 585
R569 VSS.n212 VSS.n152 585
R570 VSS.n254 VSS.n152 585
R571 VSS.n211 VSS.n210 585
R572 VSS.n210 VSS.n151 585
R573 VSS.n434 VSS.n9 585
R574 VSS.n438 VSS.n435 585
R575 VSS.n440 VSS.n439 585
R576 VSS.n442 VSS.n431 585
R577 VSS.n444 VSS.n443 585
R578 VSS.n446 VSS.n429 585
R579 VSS.n448 VSS.n447 585
R580 VSS.n449 VSS.n428 585
R581 VSS.n451 VSS.n450 585
R582 VSS.n453 VSS.n17 585
R583 VSS.n455 VSS.n454 585
R584 VSS.n456 VSS.n14 585
R585 VSS.n187 VSS.n186 585
R586 VSS.n190 VSS.n189 585
R587 VSS.n191 VSS.n185 585
R588 VSS.n185 VSS.n100 585
R589 VSS.n193 VSS.n192 585
R590 VSS.n195 VSS.n184 585
R591 VSS.n198 VSS.n197 585
R592 VSS.n199 VSS.n183 585
R593 VSS.n201 VSS.n200 585
R594 VSS.n203 VSS.n182 585
R595 VSS.n206 VSS.n205 585
R596 VSS.n207 VSS.n178 585
R597 VSS.n209 VSS.n208 585
R598 VSS.n209 VSS.n100 585
R599 VSS.n264 VSS.n263 467.284
R600 VSS.n426 VSS.n19 467.284
R601 VSS.n265 VSS.n264 404.599
R602 VSS.n386 VSS.n19 404.599
R603 VSS.n151 VSS.n150 313.615
R604 VSS.n254 VSS.n151 313.615
R605 VSS.n174 VSS.n173 313.615
R606 VSS.n225 VSS.n173 313.615
R607 VSS.t8 VSS.n225 313.615
R608 VSS.n227 VSS.t8 313.615
R609 VSS.n227 VSS.n165 313.615
R610 VSS.n239 VSS.n165 313.615
R611 VSS.n460 VSS.n10 313.615
R612 VSS.n460 VSS.n11 313.615
R613 VSS.n432 VSS.t4 278.709
R614 VSS.n179 VSS.t0 278.709
R615 VSS.n150 VSS.n100 266.572
R616 VSS.n427 VSS.n11 266.572
R617 VSS.n174 VSS.t1 263.435
R618 VSS.n239 VSS.t5 263.435
R619 VSS.n112 VSS.n99 256.663
R620 VSS.n115 VSS.n99 256.663
R621 VSS.n121 VSS.n99 256.663
R622 VSS.n123 VSS.n99 256.663
R623 VSS.n129 VSS.n99 256.663
R624 VSS.n131 VSS.n99 256.663
R625 VSS.n137 VSS.n99 256.663
R626 VSS.n140 VSS.n99 256.663
R627 VSS.n419 VSS.n418 256.663
R628 VSS.n418 VSS.n417 256.663
R629 VSS.n418 VSS.n32 256.663
R630 VSS.n418 VSS.n31 256.663
R631 VSS.n418 VSS.n30 256.663
R632 VSS.n418 VSS.n29 256.663
R633 VSS.n418 VSS.n28 256.663
R634 VSS.n418 VSS.n27 256.663
R635 VSS.n418 VSS.n26 256.663
R636 VSS.n437 VSS.n427 256.663
R637 VSS.n436 VSS.n427 256.663
R638 VSS.n445 VSS.n427 256.663
R639 VSS.n430 VSS.n427 256.663
R640 VSS.n452 VSS.n427 256.663
R641 VSS.n427 VSS.n18 256.663
R642 VSS.n188 VSS.n100 256.663
R643 VSS.n194 VSS.n100 256.663
R644 VSS.n196 VSS.n100 256.663
R645 VSS.n202 VSS.n100 256.663
R646 VSS.n204 VSS.n100 256.663
R647 VSS.n311 VSS.n75 240.244
R648 VSS.n311 VSS.n73 240.244
R649 VSS.n315 VSS.n73 240.244
R650 VSS.n315 VSS.n69 240.244
R651 VSS.n321 VSS.n69 240.244
R652 VSS.n321 VSS.n67 240.244
R653 VSS.n325 VSS.n67 240.244
R654 VSS.n325 VSS.n63 240.244
R655 VSS.n331 VSS.n63 240.244
R656 VSS.n331 VSS.n61 240.244
R657 VSS.n335 VSS.n61 240.244
R658 VSS.n335 VSS.n57 240.244
R659 VSS.n342 VSS.n57 240.244
R660 VSS.n342 VSS.n55 240.244
R661 VSS.n262 VSS.n102 240.244
R662 VSS.n148 VSS.n102 240.244
R663 VSS.n255 VSS.n148 240.244
R664 VSS.n255 VSS.n149 240.244
R665 VSS.n219 VSS.n149 240.244
R666 VSS.n224 VSS.n219 240.244
R667 VSS.n224 VSS.n172 240.244
R668 VSS.n228 VSS.n172 240.244
R669 VSS.n228 VSS.n167 240.244
R670 VSS.n238 VSS.n167 240.244
R671 VSS.n238 VSS.n168 240.244
R672 VSS.n168 VSS.n12 240.244
R673 VSS.n20 VSS.n12 240.244
R674 VSS.n425 VSS.n20 240.244
R675 VSS.n253 VSS.n153 240.244
R676 VSS.n253 VSS.n154 240.244
R677 VSS.n159 VSS.n154 240.244
R678 VSS.n160 VSS.n159 240.244
R679 VSS.n161 VSS.n160 240.244
R680 VSS.n226 VSS.n161 240.244
R681 VSS.n226 VSS.n164 240.244
R682 VSS.n240 VSS.n164 240.244
R683 VSS.n240 VSS.n13 240.244
R684 VSS.n459 VSS.n13 240.244
R685 VSS.n210 VSS.n152 240.244
R686 VSS.n175 VSS.n152 240.244
R687 VSS.n217 VSS.n175 240.244
R688 VSS.n218 VSS.n217 240.244
R689 VSS.n218 VSS.n3 240.244
R690 VSS.n4 VSS.n3 240.244
R691 VSS.n5 VSS.n4 240.244
R692 VSS.n166 VSS.n5 240.244
R693 VSS.n166 VSS.n8 240.244
R694 VSS.n461 VSS.n8 240.244
R695 VSS.n346 VSS.n53 163.367
R696 VSS.n350 VSS.n53 163.367
R697 VSS.n350 VSS.n51 163.367
R698 VSS.n354 VSS.n51 163.367
R699 VSS.n354 VSS.n49 163.367
R700 VSS.n358 VSS.n49 163.367
R701 VSS.n358 VSS.n47 163.367
R702 VSS.n362 VSS.n47 163.367
R703 VSS.n362 VSS.n45 163.367
R704 VSS.n366 VSS.n45 163.367
R705 VSS.n366 VSS.n43 163.367
R706 VSS.n370 VSS.n43 163.367
R707 VSS.n370 VSS.n41 163.367
R708 VSS.n374 VSS.n41 163.367
R709 VSS.n374 VSS.n39 163.367
R710 VSS.n378 VSS.n39 163.367
R711 VSS.n378 VSS.n37 163.367
R712 VSS.n383 VSS.n37 163.367
R713 VSS.n383 VSS.n35 163.367
R714 VSS.n387 VSS.n35 163.367
R715 VSS.n388 VSS.n387 163.367
R716 VSS.n392 VSS.n391 163.367
R717 VSS.n396 VSS.n395 163.367
R718 VSS.n400 VSS.n399 163.367
R719 VSS.n404 VSS.n403 163.367
R720 VSS.n408 VSS.n407 163.367
R721 VSS.n412 VSS.n411 163.367
R722 VSS.n416 VSS.n33 163.367
R723 VSS.n420 VSS.n25 163.367
R724 VSS.n306 VSS.n78 163.367
R725 VSS.n302 VSS.n78 163.367
R726 VSS.n302 VSS.n80 163.367
R727 VSS.n298 VSS.n80 163.367
R728 VSS.n298 VSS.n82 163.367
R729 VSS.n294 VSS.n82 163.367
R730 VSS.n294 VSS.n84 163.367
R731 VSS.n290 VSS.n84 163.367
R732 VSS.n290 VSS.n86 163.367
R733 VSS.n286 VSS.n86 163.367
R734 VSS.n286 VSS.n88 163.367
R735 VSS.n282 VSS.n88 163.367
R736 VSS.n282 VSS.n90 163.367
R737 VSS.n278 VSS.n90 163.367
R738 VSS.n278 VSS.n92 163.367
R739 VSS.n274 VSS.n92 163.367
R740 VSS.n274 VSS.n94 163.367
R741 VSS.n270 VSS.n94 163.367
R742 VSS.n270 VSS.n96 163.367
R743 VSS.n266 VSS.n96 163.367
R744 VSS.n266 VSS.n98 163.367
R745 VSS.n114 VSS.n113 163.367
R746 VSS.n116 VSS.n114 163.367
R747 VSS.n120 VSS.n109 163.367
R748 VSS.n124 VSS.n122 163.367
R749 VSS.n128 VSS.n107 163.367
R750 VSS.n132 VSS.n130 163.367
R751 VSS.n136 VSS.n105 163.367
R752 VSS.n139 VSS.n138 163.367
R753 VSS.n141 VSS.n101 163.367
R754 VSS.n189 VSS.n185 163.367
R755 VSS.n193 VSS.n185 163.367
R756 VSS.n197 VSS.n195 163.367
R757 VSS.n201 VSS.n183 163.367
R758 VSS.n205 VSS.n203 163.367
R759 VSS.n209 VSS.n178 163.367
R760 VSS.n454 VSS.n453 163.367
R761 VSS.n451 VSS.n428 163.367
R762 VSS.n447 VSS.n446 163.367
R763 VSS.n444 VSS.n431 163.367
R764 VSS.n439 VSS.n438 163.367
R765 VSS.n432 VSS.t6 123.436
R766 VSS.n179 VSS.t3 123.436
R767 VSS.n433 VSS.t7 107.338
R768 VSS.n180 VSS.t2 107.338
R769 VSS.n391 VSS.n26 71.676
R770 VSS.n395 VSS.n27 71.676
R771 VSS.n399 VSS.n28 71.676
R772 VSS.n403 VSS.n29 71.676
R773 VSS.n407 VSS.n30 71.676
R774 VSS.n411 VSS.n31 71.676
R775 VSS.n33 VSS.n32 71.676
R776 VSS.n417 VSS.n25 71.676
R777 VSS.n419 VSS.n21 71.676
R778 VSS.n112 VSS.n98 71.676
R779 VSS.n116 VSS.n115 71.676
R780 VSS.n121 VSS.n120 71.676
R781 VSS.n124 VSS.n123 71.676
R782 VSS.n129 VSS.n128 71.676
R783 VSS.n132 VSS.n131 71.676
R784 VSS.n137 VSS.n136 71.676
R785 VSS.n140 VSS.n139 71.676
R786 VSS.n113 VSS.n112 71.676
R787 VSS.n115 VSS.n109 71.676
R788 VSS.n122 VSS.n121 71.676
R789 VSS.n123 VSS.n107 71.676
R790 VSS.n130 VSS.n129 71.676
R791 VSS.n131 VSS.n105 71.676
R792 VSS.n138 VSS.n137 71.676
R793 VSS.n141 VSS.n140 71.676
R794 VSS.n420 VSS.n419 71.676
R795 VSS.n417 VSS.n416 71.676
R796 VSS.n412 VSS.n32 71.676
R797 VSS.n408 VSS.n31 71.676
R798 VSS.n404 VSS.n30 71.676
R799 VSS.n400 VSS.n29 71.676
R800 VSS.n396 VSS.n28 71.676
R801 VSS.n392 VSS.n27 71.676
R802 VSS.n388 VSS.n26 71.676
R803 VSS.n188 VSS.n187 71.676
R804 VSS.n194 VSS.n193 71.676
R805 VSS.n197 VSS.n196 71.676
R806 VSS.n202 VSS.n201 71.676
R807 VSS.n205 VSS.n204 71.676
R808 VSS.n454 VSS.n18 71.676
R809 VSS.n452 VSS.n451 71.676
R810 VSS.n447 VSS.n430 71.676
R811 VSS.n445 VSS.n444 71.676
R812 VSS.n439 VSS.n436 71.676
R813 VSS.n437 VSS.n9 71.676
R814 VSS.n438 VSS.n437 71.676
R815 VSS.n436 VSS.n431 71.676
R816 VSS.n446 VSS.n445 71.676
R817 VSS.n430 VSS.n428 71.676
R818 VSS.n453 VSS.n452 71.676
R819 VSS.n18 VSS.n14 71.676
R820 VSS.n189 VSS.n188 71.676
R821 VSS.n195 VSS.n194 71.676
R822 VSS.n196 VSS.n183 71.676
R823 VSS.n203 VSS.n202 71.676
R824 VSS.n204 VSS.n178 71.676
R825 VSS.n264 VSS.n99 62.7232
R826 VSS.n418 VSS.n19 62.7232
R827 VSS.n254 VSS.t1 50.1787
R828 VSS.t5 VSS.n10 50.1787
R829 VSS.n263 VSS.n100 47.0426
R830 VSS.n427 VSS.n426 47.0426
R831 VSS.n441 VSS.n433 34.3278
R832 VSS.n181 VSS.n180 34.3278
R833 VSS.n347 VSS.n54 29.5386
R834 VSS.n423 VSS.n422 29.5386
R835 VSS.n308 VSS.n307 29.5386
R836 VSS.n144 VSS.n143 29.5386
R837 VSS.n457 VSS.n456 26.7532
R838 VSS.n434 VSS.n7 26.7532
R839 VSS.n186 VSS.n157 26.7532
R840 VSS.n208 VSS.n177 26.7532
R841 VSS.n310 VSS.n76 19.3944
R842 VSS.n310 VSS.n72 19.3944
R843 VSS.n316 VSS.n72 19.3944
R844 VSS.n316 VSS.n70 19.3944
R845 VSS.n320 VSS.n70 19.3944
R846 VSS.n320 VSS.n66 19.3944
R847 VSS.n326 VSS.n66 19.3944
R848 VSS.n326 VSS.n64 19.3944
R849 VSS.n330 VSS.n64 19.3944
R850 VSS.n330 VSS.n60 19.3944
R851 VSS.n336 VSS.n60 19.3944
R852 VSS.n336 VSS.n58 19.3944
R853 VSS.n341 VSS.n58 19.3944
R854 VSS.n341 VSS.n340 19.3944
R855 VSS.n261 VSS.n260 19.3944
R856 VSS.n260 VSS.n145 19.3944
R857 VSS.n256 VSS.n145 19.3944
R858 VSS.n256 VSS.n147 19.3944
R859 VSS.n220 VSS.n147 19.3944
R860 VSS.n223 VSS.n220 19.3944
R861 VSS.n223 VSS.n171 19.3944
R862 VSS.n229 VSS.n171 19.3944
R863 VSS.n229 VSS.n169 19.3944
R864 VSS.n237 VSS.n169 19.3944
R865 VSS.n237 VSS.n236 19.3944
R866 VSS.n236 VSS.n235 19.3944
R867 VSS.n235 VSS.n22 19.3944
R868 VSS.n424 VSS.n22 19.3944
R869 VSS.n252 VSS.n155 19.3944
R870 VSS.n252 VSS.n156 19.3944
R871 VSS.n248 VSS.n156 19.3944
R872 VSS.n248 VSS.n247 19.3944
R873 VSS.n247 VSS.n246 19.3944
R874 VSS.n246 VSS.n162 19.3944
R875 VSS.n242 VSS.n162 19.3944
R876 VSS.n242 VSS.n241 19.3944
R877 VSS.n241 VSS.n15 19.3944
R878 VSS.n458 VSS.n15 19.3944
R879 VSS.n212 VSS.n211 19.3944
R880 VSS.n212 VSS.n176 19.3944
R881 VSS.n216 VSS.n176 19.3944
R882 VSS.n216 VSS.n2 19.3944
R883 VSS.n469 VSS.n2 19.3944
R884 VSS.n469 VSS.n468 19.3944
R885 VSS.n468 VSS.n467 19.3944
R886 VSS.n467 VSS.n6 19.3944
R887 VSS.n463 VSS.n6 19.3944
R888 VSS.n463 VSS.n462 19.3944
R889 VSS.n433 VSS.n432 16.0975
R890 VSS.n180 VSS.n179 16.0975
R891 VSS.n348 VSS.n347 10.6151
R892 VSS.n349 VSS.n348 10.6151
R893 VSS.n349 VSS.n50 10.6151
R894 VSS.n355 VSS.n50 10.6151
R895 VSS.n356 VSS.n355 10.6151
R896 VSS.n357 VSS.n356 10.6151
R897 VSS.n357 VSS.n46 10.6151
R898 VSS.n363 VSS.n46 10.6151
R899 VSS.n364 VSS.n363 10.6151
R900 VSS.n365 VSS.n364 10.6151
R901 VSS.n365 VSS.n42 10.6151
R902 VSS.n371 VSS.n42 10.6151
R903 VSS.n372 VSS.n371 10.6151
R904 VSS.n373 VSS.n372 10.6151
R905 VSS.n373 VSS.n38 10.6151
R906 VSS.n379 VSS.n38 10.6151
R907 VSS.n380 VSS.n379 10.6151
R908 VSS.n382 VSS.n380 10.6151
R909 VSS.n382 VSS.n381 10.6151
R910 VSS.n381 VSS.n34 10.6151
R911 VSS.n389 VSS.n34 10.6151
R912 VSS.n390 VSS.n389 10.6151
R913 VSS.n393 VSS.n390 10.6151
R914 VSS.n394 VSS.n393 10.6151
R915 VSS.n397 VSS.n394 10.6151
R916 VSS.n398 VSS.n397 10.6151
R917 VSS.n401 VSS.n398 10.6151
R918 VSS.n402 VSS.n401 10.6151
R919 VSS.n405 VSS.n402 10.6151
R920 VSS.n406 VSS.n405 10.6151
R921 VSS.n409 VSS.n406 10.6151
R922 VSS.n410 VSS.n409 10.6151
R923 VSS.n413 VSS.n410 10.6151
R924 VSS.n414 VSS.n413 10.6151
R925 VSS.n415 VSS.n414 10.6151
R926 VSS.n415 VSS.n24 10.6151
R927 VSS.n421 VSS.n24 10.6151
R928 VSS.n422 VSS.n421 10.6151
R929 VSS.n307 VSS.n77 10.6151
R930 VSS.n301 VSS.n77 10.6151
R931 VSS.n301 VSS.n300 10.6151
R932 VSS.n300 VSS.n299 10.6151
R933 VSS.n299 VSS.n81 10.6151
R934 VSS.n293 VSS.n81 10.6151
R935 VSS.n293 VSS.n292 10.6151
R936 VSS.n292 VSS.n291 10.6151
R937 VSS.n291 VSS.n85 10.6151
R938 VSS.n285 VSS.n85 10.6151
R939 VSS.n285 VSS.n284 10.6151
R940 VSS.n284 VSS.n283 10.6151
R941 VSS.n283 VSS.n89 10.6151
R942 VSS.n277 VSS.n89 10.6151
R943 VSS.n277 VSS.n276 10.6151
R944 VSS.n276 VSS.n275 10.6151
R945 VSS.n275 VSS.n93 10.6151
R946 VSS.n269 VSS.n93 10.6151
R947 VSS.n269 VSS.n268 10.6151
R948 VSS.n268 VSS.n267 10.6151
R949 VSS.n267 VSS.n97 10.6151
R950 VSS.n111 VSS.n97 10.6151
R951 VSS.n111 VSS.n110 10.6151
R952 VSS.n117 VSS.n110 10.6151
R953 VSS.n118 VSS.n117 10.6151
R954 VSS.n119 VSS.n118 10.6151
R955 VSS.n119 VSS.n108 10.6151
R956 VSS.n125 VSS.n108 10.6151
R957 VSS.n126 VSS.n125 10.6151
R958 VSS.n127 VSS.n126 10.6151
R959 VSS.n127 VSS.n106 10.6151
R960 VSS.n133 VSS.n106 10.6151
R961 VSS.n134 VSS.n133 10.6151
R962 VSS.n135 VSS.n134 10.6151
R963 VSS.n135 VSS.n104 10.6151
R964 VSS.n104 VSS.n103 10.6151
R965 VSS.n142 VSS.n103 10.6151
R966 VSS.n143 VSS.n142 10.6151
R967 VSS.n456 VSS.n455 10.6151
R968 VSS.n455 VSS.n17 10.6151
R969 VSS.n450 VSS.n17 10.6151
R970 VSS.n450 VSS.n449 10.6151
R971 VSS.n449 VSS.n448 10.6151
R972 VSS.n448 VSS.n429 10.6151
R973 VSS.n443 VSS.n429 10.6151
R974 VSS.n443 VSS.n442 10.6151
R975 VSS.n440 VSS.n435 10.6151
R976 VSS.n435 VSS.n434 10.6151
R977 VSS.n190 VSS.n186 10.6151
R978 VSS.n191 VSS.n190 10.6151
R979 VSS.n192 VSS.n191 10.6151
R980 VSS.n192 VSS.n184 10.6151
R981 VSS.n198 VSS.n184 10.6151
R982 VSS.n199 VSS.n198 10.6151
R983 VSS.n200 VSS.n199 10.6151
R984 VSS.n200 VSS.n182 10.6151
R985 VSS.n207 VSS.n206 10.6151
R986 VSS.n208 VSS.n207 10.6151
R987 VSS.n260 VSS.n259 9.3005
R988 VSS.n258 VSS.n145 9.3005
R989 VSS.n257 VSS.n256 9.3005
R990 VSS.n147 VSS.n146 9.3005
R991 VSS.n221 VSS.n220 9.3005
R992 VSS.n223 VSS.n222 9.3005
R993 VSS.n171 VSS.n170 9.3005
R994 VSS.n230 VSS.n229 9.3005
R995 VSS.n231 VSS.n169 9.3005
R996 VSS.n237 VSS.n232 9.3005
R997 VSS.n236 VSS.n233 9.3005
R998 VSS.n235 VSS.n234 9.3005
R999 VSS.n23 VSS.n22 9.3005
R1000 VSS.n424 VSS.n423 9.3005
R1001 VSS.n261 VSS.n144 9.3005
R1002 VSS.n308 VSS.n76 9.3005
R1003 VSS.n310 VSS.n309 9.3005
R1004 VSS.n72 VSS.n71 9.3005
R1005 VSS.n317 VSS.n316 9.3005
R1006 VSS.n318 VSS.n70 9.3005
R1007 VSS.n320 VSS.n319 9.3005
R1008 VSS.n66 VSS.n65 9.3005
R1009 VSS.n327 VSS.n326 9.3005
R1010 VSS.n328 VSS.n64 9.3005
R1011 VSS.n330 VSS.n329 9.3005
R1012 VSS.n60 VSS.n59 9.3005
R1013 VSS.n337 VSS.n336 9.3005
R1014 VSS.n338 VSS.n58 9.3005
R1015 VSS.n341 VSS.n339 9.3005
R1016 VSS.n340 VSS.n54 9.3005
R1017 VSS.n468 VSS.n0 9.3005
R1018 VSS.n467 VSS.n466 9.3005
R1019 VSS.n465 VSS.n6 9.3005
R1020 VSS.n464 VSS.n463 9.3005
R1021 VSS.n462 VSS.n7 9.3005
R1022 VSS.n252 VSS.n251 9.3005
R1023 VSS.n250 VSS.n156 9.3005
R1024 VSS.n249 VSS.n248 9.3005
R1025 VSS.n247 VSS.n158 9.3005
R1026 VSS.n246 VSS.n245 9.3005
R1027 VSS.n244 VSS.n162 9.3005
R1028 VSS.n243 VSS.n242 9.3005
R1029 VSS.n241 VSS.n163 9.3005
R1030 VSS.n16 VSS.n15 9.3005
R1031 VSS.n458 VSS.n457 9.3005
R1032 VSS.n157 VSS.n155 9.3005
R1033 VSS.n213 VSS.n212 9.3005
R1034 VSS.n214 VSS.n176 9.3005
R1035 VSS.n216 VSS.n215 9.3005
R1036 VSS.n2 VSS.n1 9.3005
R1037 VSS.n211 VSS.n177 9.3005
R1038 VSS.n470 VSS.n469 9.3005
R1039 VSS.n442 VSS.n441 7.64928
R1040 VSS.n182 VSS.n181 7.64928
R1041 VSS.n441 VSS.n440 2.96635
R1042 VSS.n206 VSS.n181 2.96635
R1043 VSS.n259 VSS.n144 0.152939
R1044 VSS.n259 VSS.n258 0.152939
R1045 VSS.n258 VSS.n257 0.152939
R1046 VSS.n257 VSS.n146 0.152939
R1047 VSS.n221 VSS.n146 0.152939
R1048 VSS.n222 VSS.n221 0.152939
R1049 VSS.n222 VSS.n170 0.152939
R1050 VSS.n230 VSS.n170 0.152939
R1051 VSS.n231 VSS.n230 0.152939
R1052 VSS.n232 VSS.n231 0.152939
R1053 VSS.n233 VSS.n232 0.152939
R1054 VSS.n234 VSS.n233 0.152939
R1055 VSS.n234 VSS.n23 0.152939
R1056 VSS.n423 VSS.n23 0.152939
R1057 VSS.n309 VSS.n308 0.152939
R1058 VSS.n309 VSS.n71 0.152939
R1059 VSS.n317 VSS.n71 0.152939
R1060 VSS.n318 VSS.n317 0.152939
R1061 VSS.n319 VSS.n318 0.152939
R1062 VSS.n319 VSS.n65 0.152939
R1063 VSS.n327 VSS.n65 0.152939
R1064 VSS.n328 VSS.n327 0.152939
R1065 VSS.n329 VSS.n328 0.152939
R1066 VSS.n329 VSS.n59 0.152939
R1067 VSS.n337 VSS.n59 0.152939
R1068 VSS.n338 VSS.n337 0.152939
R1069 VSS.n339 VSS.n338 0.152939
R1070 VSS.n339 VSS.n54 0.152939
R1071 VSS.n466 VSS.n0 0.152939
R1072 VSS.n466 VSS.n465 0.152939
R1073 VSS.n465 VSS.n464 0.152939
R1074 VSS.n464 VSS.n7 0.152939
R1075 VSS.n251 VSS.n157 0.152939
R1076 VSS.n251 VSS.n250 0.152939
R1077 VSS.n250 VSS.n249 0.152939
R1078 VSS.n249 VSS.n158 0.152939
R1079 VSS.n245 VSS.n158 0.152939
R1080 VSS.n245 VSS.n244 0.152939
R1081 VSS.n244 VSS.n243 0.152939
R1082 VSS.n243 VSS.n163 0.152939
R1083 VSS.n163 VSS.n16 0.152939
R1084 VSS.n457 VSS.n16 0.152939
R1085 VSS.n213 VSS.n177 0.152939
R1086 VSS.n214 VSS.n213 0.152939
R1087 VSS.n215 VSS.n214 0.152939
R1088 VSS.n215 VSS.n1 0.152939
R1089 VSS.n470 VSS.n1 0.13922
R1090 VSS VSS.n0 0.0767195
R1091 VSS VSS.n470 0.063
C0 VIN VGP 0.151302f
C1 VOUT VIN 0.949141f
C2 VGN VCC 0.001774f
C3 VOUT VGP 0.128336f
C4 VIN VGN 0.096189f
C5 VGP VGN 0.002f
C6 VIN VCC 0.555421f
C7 VOUT VGN 0.071863f
C8 VGP VCC 0.376799f
C9 VOUT VCC 0.678351f
C10 VGN VSS 0.438504f
C11 VOUT VSS 0.734895f
C12 VIN VSS 0.673971f
C13 VGP VSS 0.077729f
C14 VCC VSS 8.186231f
.ends

