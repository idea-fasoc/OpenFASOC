* NGSPICE file created from opamp_sample_0006.ext - technology: sky130A

.subckt opamp_sample_0006 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 a_n10683_10810.t5 a_n10683_10810.t4 a_n10827_11007.t10 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X1 a_n10827_11007.t9 a_n10683_10810.t18 a_n10683_10810.t19 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X2 GND.t23 CS_BIAS.t8 VOUT.t7 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X3 a_n17822_7210.t3 VN.t7 a_n2596_242.t4 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=2.94 as=1.6416 ps=6 w=2.28 l=5.28
X4 VDD.t120 VDD.t118 VDD.t119 VDD.t69 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X5 VDD.t117 VDD.t115 VDD.t116 VDD.t82 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X6 VOUT.t34 a_n17822_7210.t12 VDD.t24 VDD.t11 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X7 a_n10827_11007.t8 a_n10683_10810.t6 a_n10683_10810.t7 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X8 GND.t160 GND.t158 GND.t159 GND.t56 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X9 VOUT.t46 a_n6906_9317.t0 sky130_fd_pr__cap_mim_m3_1 l=15.59 w=6.85
X10 VOUT.t6 CS_BIAS.t9 GND.t22 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X11 VDD.t114 VDD.t112 VDD.t113 VDD.t50 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X12 GND.t157 GND.t155 GND.t156 GND.t56 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X13 VDD.t111 VDD.t109 VDD.t110 VDD.t46 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X14 a_n10827_11007.t15 a_n10683_10810.t20 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X15 VN.t6 GND.t152 GND.t154 GND.t153 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X16 GND.t151 GND.t149 GND.t150 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X17 VDD.t108 VDD.t106 VDD.t107 VDD.t38 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X18 GND.t148 GND.t146 GND.t147 GND.t42 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0 ps=0 w=2.28 l=5.28
X19 GND.t139 GND.t137 GND.t138 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0 ps=0 w=2.28 l=5.28
X20 VOUT.t1 a_n17822_7210.t13 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X21 VDD.t105 VDD.t103 VDD.t104 VDD.t38 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X22 VOUT.t24 a_n17822_7210.t14 VDD.t14 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X23 VDD.t164 a_n17822_7210.t15 VOUT.t40 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X24 VOUT.t45 a_n17822_7210.t16 VDD.t169 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X25 VOUT.t32 a_n17822_7210.t17 VDD.t22 VDD.t4 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X26 VOUT.t28 a_n17822_7210.t18 VDD.t18 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X27 a_n2596_242.t3 VP.t7 a_n10683_10810.t2 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0.7524 ps=2.94 w=2.28 l=5.28
X28 VDD.t1 a_n17822_7210.t19 VOUT.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X29 GND.t145 GND.t143 VP.t6 GND.t144 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X30 a_n17822_7210.t5 a_n10683_10810.t21 a_n6906_9317.t8 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X31 GND.t21 CS_BIAS.t10 VOUT.t5 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X32 VOUT.t3 CS_BIAS.t11 GND.t20 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X33 VOUT.t8 CS_BIAS.t12 GND.t19 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X34 GND.t142 GND.t140 GND.t141 GND.t38 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X35 a_n10683_10810.t0 VP.t8 a_n2596_242.t0 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=2.94 as=1.6416 ps=6 w=2.28 l=5.28
X36 VOUT.t35 a_n17822_7210.t20 VDD.t25 VDD.t11 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X37 a_n6906_9317.t16 a_n10683_10810.t22 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X38 GND.t136 GND.t134 VP.t5 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X39 VDD.t102 VDD.t100 VDD.t101 VDD.t50 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X40 VDD.t99 VDD.t97 VDD.t98 VDD.t34 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X41 VOUT.t13 CS_BIAS.t13 GND.t18 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X42 GND.t17 CS_BIAS.t14 VOUT.t14 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X43 GND.t16 CS_BIAS.t15 VOUT.t15 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X44 VOUT.t31 a_n17822_7210.t21 VDD.t21 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X45 VOUT.t21 a_n17822_7210.t22 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X46 VDD.t96 VDD.t94 VDD.t95 VDD.t38 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X47 VN.t5 GND.t131 GND.t133 GND.t132 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X48 VOUT.t2 CS_BIAS.t16 GND.t15 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X49 VDD.t7 a_n17822_7210.t23 VOUT.t19 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X50 GND.t130 GND.t128 GND.t129 GND.t56 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X51 GND.t127 GND.t125 VP.t4 GND.t126 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X52 a_n10683_10810.t17 a_n10683_10810.t16 a_n10827_11007.t7 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X53 VDD.t93 VDD.t91 VDD.t92 VDD.t38 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X54 GND.t124 GND.t122 GND.t123 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X55 VOUT.t42 a_n17822_7210.t24 VDD.t166 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X56 a_n10827_11007.t14 a_n10683_10810.t23 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X57 a_n10827_11007.t13 a_n10683_10810.t24 VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X58 a_10955_11007# a_10955_11007# a_10955_11007# VDD.t28 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=4.1904 ps=14.52 w=2.91 l=5.29
X59 GND.t121 GND.t119 GND.t120 GND.t38 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X60 GND.t118 GND.t116 VP.t3 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X61 a_n17822_7210.t9 a_n10683_10810.t25 a_n6906_9317.t7 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X62 VDD.t152 a_n10683_10810.t26 a_n10827_11007.t12 VDD.t151 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X63 a_n10827_11007.t1 a_n10683_10810.t27 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X64 VDD.t148 a_n10683_10810.t28 a_n10827_11007.t0 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X65 GND.t11 CS_BIAS.t4 CS_BIAS.t5 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X66 VDD.t90 VDD.t88 VDD.t89 VDD.t34 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X67 a_n6906_9317.t6 a_n10683_10810.t29 a_n17822_7210.t6 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X68 VOUT.t10 CS_BIAS.t17 GND.t14 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X69 VDD.t145 a_n10683_10810.t30 a_n10827_11007.t2 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X70 VOUT.t16 CS_BIAS.t18 GND.t13 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X71 CS_BIAS.t1 CS_BIAS.t0 GND.t12 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X72 VDD.t143 a_n10683_10810.t31 a_n6906_9317.t15 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X73 VOUT.t25 a_n17822_7210.t25 VDD.t15 VDD.t11 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X74 a_n17822_7210.t7 a_n10683_10810.t32 a_n6906_9317.t5 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X75 a_n6906_9317.t4 a_n10683_10810.t33 a_n17822_7210.t4 VDD.t122 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X76 GND.t10 CS_BIAS.t19 VOUT.t4 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X77 a_n6906_9317.t14 a_n10683_10810.t34 VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X78 CS_BIAS.t7 CS_BIAS.t6 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X79 a_n12301_11007# a_n12301_11007# a_n12301_11007# VDD.t27 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=4.1904 ps=14.52 w=2.91 l=5.29
X80 VN.t4 GND.t110 GND.t112 GND.t111 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X81 VDD.t87 VDD.t85 VDD.t86 VDD.t50 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X82 a_n6906_9317.t3 a_n10683_10810.t35 a_n17822_7210.t8 VDD.t124 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X83 VOUT.t27 a_n17822_7210.t26 VDD.t17 VDD.t11 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X84 VDD.t84 VDD.t81 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X85 GND.t7 CS_BIAS.t2 CS_BIAS.t3 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X86 GND.t115 GND.t113 GND.t114 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X87 VDD.t138 a_n10683_10810.t36 a_n6906_9317.t13 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X88 VOUT.t30 a_n17822_7210.t27 VDD.t20 VDD.t4 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X89 VDD.t162 a_n17822_7210.t28 VOUT.t38 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X90 VDD.t136 a_n10683_10810.t37 a_n6906_9317.t12 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X91 VDD.t80 VDD.t78 VDD.t79 VDD.t30 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X92 VDD.t77 VDD.t75 VDD.t76 VDD.t42 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X93 VDD.t134 a_n10683_10810.t38 a_n10827_11007.t11 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X94 VP.t2 GND.t107 GND.t109 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X95 a_n6906_9317.t11 a_n10683_10810.t39 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X96 VOUT.t20 a_n17822_7210.t29 VDD.t8 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X97 VDD.t13 a_n17822_7210.t30 VOUT.t23 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X98 VDD.t74 VDD.t72 VDD.t73 VDD.t34 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X99 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=1.6056 ps=5.9 w=2.23 l=4.26
X100 GND.t106 GND.t104 GND.t105 GND.t38 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X101 a_n17822_7210.t2 VN.t8 a_n2596_242.t7 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=2.94 as=1.6416 ps=6 w=2.28 l=5.28
X102 GND.t6 CS_BIAS.t20 VOUT.t11 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X103 a_n10827_11007.t6 a_n10683_10810.t10 a_n10683_10810.t11 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X104 VDD.t71 VDD.t68 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X105 a_n6906_9317.t10 a_n10683_10810.t40 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X106 GND.t103 GND.t100 GND.t102 GND.t101 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0 ps=0 w=2.28 l=5.28
X107 GND.t99 GND.t96 GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=0 ps=0 w=2.23 l=4.26
X108 a_n17822_7210.t10 a_n10683_10810.t41 a_n6906_9317.t2 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X109 GND.t95 GND.t93 GND.t94 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X110 GND.t92 GND.t90 GND.t91 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X111 VDD.t126 a_n10683_10810.t42 a_n6906_9317.t9 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=2.0952 ps=7.26 w=2.91 l=5.29
X112 VOUT.t12 CS_BIAS.t21 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.9801 pd=3.63 as=2.1384 ps=7.38 w=2.97 l=5.77
X113 VDD.t67 VDD.t65 VDD.t66 VDD.t50 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X114 VOUT.t22 a_n17822_7210.t31 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X115 GND.t89 GND.t87 VN.t3 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X116 VP.t1 GND.t84 GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X117 VDD.t26 a_n17822_7210.t32 VOUT.t36 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X118 VOUT.t33 a_n17822_7210.t33 VDD.t23 VDD.t4 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X119 VDD.t64 VDD.t62 VDD.t63 VDD.t42 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X120 VDD.t61 VDD.t59 VDD.t60 VDD.t42 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X121 GND.t83 GND.t81 GND.t82 GND.t56 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X122 a_n2596_242.t6 VN.t9 a_n17822_7210.t1 GND.t31 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0.7524 ps=2.94 w=2.28 l=5.28
X123 VDD.t168 a_n17822_7210.t34 VOUT.t44 VDD.t6 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X124 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=1.6056 ps=5.9 w=2.23 l=4.26
X125 GND.t80 GND.t78 VN.t2 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X126 VP.t0 GND.t75 GND.t77 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X127 VDD.t58 VDD.t56 VDD.t57 VDD.t34 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X128 GND.t74 GND.t72 GND.t73 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X129 a_n10683_10810.t15 a_n10683_10810.t14 a_n10827_11007.t5 VDD.t124 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X130 VOUT.t39 a_n17822_7210.t35 VDD.t163 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X131 a_n2596_242.t8 DIFFPAIR_BIAS.t4 GND.t162 GND.t161 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=1.6056 ps=5.9 w=2.23 l=4.26
X132 VDD.t165 a_n17822_7210.t36 VOUT.t41 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X133 GND.t71 GND.t69 GND.t70 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X134 a_n10683_10810.t3 VP.t9 a_n2596_242.t9 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.7524 pd=2.94 as=1.6416 ps=6 w=2.28 l=5.28
X135 GND.t68 GND.t66 VN.t1 GND.t67 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X136 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=0 ps=0 w=2.23 l=4.26
X137 a_n2596_242.t1 DIFFPAIR_BIAS.t5 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.6056 pd=5.9 as=1.6056 ps=5.9 w=2.23 l=4.26
X138 a_n2596_242.t5 VN.t10 a_n17822_7210.t0 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0.7524 ps=2.94 w=2.28 l=5.28
X139 GND.t61 GND.t59 VN.t0 GND.t60 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X140 GND.t3 CS_BIAS.t22 VOUT.t17 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X141 GND.t58 GND.t55 GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X142 VDD.t167 a_n17822_7210.t37 VOUT.t43 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X143 GND.t54 GND.t51 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X144 GND.t50 GND.t48 GND.t49 GND.t38 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X145 VDD.t55 VDD.t53 VDD.t54 VDD.t42 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X146 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X147 a_n6906_9317.t1 a_n10683_10810.t43 a_n17822_7210.t11 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X148 GND.t1 CS_BIAS.t23 VOUT.t9 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0.9801 ps=3.63 w=2.97 l=5.77
X149 a_n2596_242.t2 VP.t10 a_n10683_10810.t1 GND.t31 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0.7524 ps=2.94 w=2.28 l=5.28
X150 VDD.t48 VDD.t45 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X151 VOUT.t26 a_n17822_7210.t38 VDD.t16 VDD.t4 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X152 VDD.t44 VDD.t41 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X153 VOUT.t47 a_n6906_9317.t0 sky130_fd_pr__cap_mim_m3_1 l=15.59 w=6.85
X154 VOUT.t29 a_n17822_7210.t39 VDD.t19 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=3.6432 ps=11.56 w=5.06 l=4.69
X155 VDD.t40 VDD.t37 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X156 VDD.t161 a_n17822_7210.t40 VOUT.t37 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.6698 pd=5.72 as=1.6698 ps=5.72 w=5.06 l=4.69
X157 a_n10683_10810.t13 a_n10683_10810.t12 a_n10827_11007.t4 VDD.t122 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0.9603 ps=3.57 w=2.91 l=5.29
X158 VDD.t36 VDD.t33 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=0 ps=0 w=5.06 l=4.69
X159 GND.t47 GND.t45 GND.t46 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X160 GND.t44 GND.t41 GND.t43 GND.t42 sky130_fd_pr__nfet_01v8 ad=1.6416 pd=6 as=0 ps=0 w=2.28 l=5.28
X161 a_n10827_11007.t3 a_n10683_10810.t8 a_n10683_10810.t9 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.9603 pd=3.57 as=0.9603 ps=3.57 w=2.91 l=5.29
X162 VOUT.t18 a_n17822_7210.t41 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=3.6432 pd=11.56 as=1.6698 ps=5.72 w=5.06 l=4.69
X163 GND.t40 GND.t37 GND.t39 GND.t38 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
X164 VDD.t32 VDD.t29 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=2.0952 pd=7.26 as=0 ps=0 w=2.91 l=5.29
X165 GND.t36 GND.t33 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.1384 pd=7.38 as=0 ps=0 w=2.97 l=5.77
R0 a_n10683_10810.n9 a_n10683_10810.n6 1.65239
R1 a_n10683_10810.n10 a_n10683_10810.n0 1.65239
R2 a_n10683_10810.n12 a_n10683_10810.t13 139.797
R3 a_n10683_10810.n11 a_n10683_10810.t11 139.797
R4 a_n10683_10810.n11 a_n10683_10810.t15 138.088
R5 a_n10683_10810.n12 a_n10683_10810.t7 138.087
R6 a_n10683_10810.n14 a_n10683_10810.t2 118.799
R7 a_n10683_10810.n11 a_n10683_10810.n15 115.746
R8 a_n10683_10810.n18 a_n10683_10810.n12 115.746
R9 a_n10683_10810.n14 a_n10683_10810.t1 88.9385
R10 a_n10683_10810.n4 a_n10683_10810.n3 5.3041
R11 a_n10683_10810.n7 a_n10683_10810.n0 2.34331
R12 a_n10683_10810.n17 a_n10683_10810.n7 64.6446
R13 a_n10683_10810.n10 a_n10683_10810.n17 64.6624
R14 a_n10683_10810.t6 a_n10683_10810.n10 33.5923
R15 a_n10683_10810.n8 a_n10683_10810.n6 2.34331
R16 a_n10683_10810.n16 a_n10683_10810.n8 64.6446
R17 a_n10683_10810.n9 a_n10683_10810.n16 64.6624
R18 a_n10683_10810.t25 a_n10683_10810.n9 33.5923
R19 a_n10683_10810.n3 a_n10683_10810.n14 24.432
R20 a_n10683_10810.n15 a_n10683_10810.t19 22.3407
R21 a_n10683_10810.n15 a_n10683_10810.t17 22.3407
R22 a_n10683_10810.n18 a_n10683_10810.t9 22.3407
R23 a_n10683_10810.t5 a_n10683_10810.n18 22.3407
R24 a_n10683_10810.n6 a_n10683_10810.n13 19.2399
R25 a_n10683_10810.n3 a_n10683_10810.n2 6.00387
R26 a_n10683_10810.t1 a_n10683_10810.t3 17.3689
R27 a_n10683_10810.t2 a_n10683_10810.t0 17.3689
R28 a_n10683_10810.n13 a_n10683_10810.n2 5.69867
R29 a_n10683_10810.n1 a_n10683_10810.n0 15.6527
R30 a_n10683_10810.n4 a_n10683_10810.t21 49.6596
R31 a_n10683_10810.n4 a_n10683_10810.t43 42.9336
R32 a_n10683_10810.n3 a_n10683_10810.t41 46.8496
R33 a_n10683_10810.n5 a_n10683_10810.t18 43.7124
R34 a_n10683_10810.n3 a_n10683_10810.t16 44.8617
R35 a_n10683_10810.n3 a_n10683_10810.t10 46.5211
R36 a_n10683_10810.n0 a_n10683_10810.t12 45.0818
R37 a_n10683_10810.n7 a_n10683_10810.t8 44.3575
R38 a_n10683_10810.n17 a_n10683_10810.t4 13.2578
R39 a_n10683_10810.n6 a_n10683_10810.t35 45.0818
R40 a_n10683_10810.n8 a_n10683_10810.t32 44.3575
R41 a_n10683_10810.n16 a_n10683_10810.t29 13.2578
R42 a_n10683_10810.n1 a_n10683_10810.t26 45.5055
R43 a_n10683_10810.n1 a_n10683_10810.t20 45.0124
R44 a_n10683_10810.n1 a_n10683_10810.t38 46.8496
R45 a_n10683_10810.n1 a_n10683_10810.t30 44.2702
R46 a_n10683_10810.n1 a_n10683_10810.t24 44.6185
R47 a_n10683_10810.n1 a_n10683_10810.t28 47.6796
R48 a_n10683_10810.n1 a_n10683_10810.t37 45.5055
R49 a_n10683_10810.n1 a_n10683_10810.t40 45.0124
R50 a_n10683_10810.n1 a_n10683_10810.t42 46.8496
R51 a_n10683_10810.n1 a_n10683_10810.t36 44.3336
R52 a_n10683_10810.n1 a_n10683_10810.t34 44.6185
R53 a_n10683_10810.n1 a_n10683_10810.t31 47.6796
R54 a_n10683_10810.n3 a_n10683_10810.n5 3.66108
R55 a_n10683_10810.n13 a_n10683_10810.n11 10.1708
R56 a_n10683_10810.n0 a_n10683_10810.n6 9.29361
R57 a_n10683_10810.n3 a_n10683_10810.t33 31.8245
R58 a_n10683_10810.n5 a_n10683_10810.t14 35.7049
R59 a_n10683_10810.n1 a_n10683_10810.t23 31.8245
R60 a_n10683_10810.n1 a_n10683_10810.t27 34.3477
R61 a_n10683_10810.n1 a_n10683_10810.t22 31.8245
R62 a_n10683_10810.n1 a_n10683_10810.t39 34.2167
R63 a_n10683_10810.n12 a_n10683_10810.n1 23.526
R64 a_n10683_10810.n2 a_n10683_10810.n1 19.9385
R65 a_n10827_11007.n0 a_n10827_11007.t1 139.797
R66 a_n10827_11007.n1 a_n10827_11007.t11 138.088
R67 a_n10827_11007.n0 a_n10827_11007.t14 138.088
R68 a_n10827_11007.n0 a_n10827_11007.t0 138.088
R69 a_n10827_11007.n9 a_n10827_11007.n2 137.044
R70 a_n10827_11007.n5 a_n10827_11007.n3 136.078
R71 a_n10827_11007.n5 a_n10827_11007.n4 135.334
R72 a_n10827_11007.n10 a_n10827_11007.n9 135.334
R73 a_n10827_11007.n1 a_n10827_11007.n7 115.746
R74 a_n10827_11007.n0 a_n10827_11007.n6 115.746
R75 a_n10827_11007.n2 a_n10827_11007.t4 22.3407
R76 a_n10827_11007.n2 a_n10827_11007.t3 22.3407
R77 a_n10827_11007.n7 a_n10827_11007.t12 22.3407
R78 a_n10827_11007.n7 a_n10827_11007.t15 22.3407
R79 a_n10827_11007.n6 a_n10827_11007.t2 22.3407
R80 a_n10827_11007.n6 a_n10827_11007.t13 22.3407
R81 a_n10827_11007.n4 a_n10827_11007.t7 22.3407
R82 a_n10827_11007.n4 a_n10827_11007.t6 22.3407
R83 a_n10827_11007.n3 a_n10827_11007.t5 22.3407
R84 a_n10827_11007.n3 a_n10827_11007.t9 22.3407
R85 a_n10827_11007.t10 a_n10827_11007.n10 22.3407
R86 a_n10827_11007.n10 a_n10827_11007.t8 22.3407
R87 a_n10827_11007.n8 a_n10827_11007.n5 17.7024
R88 a_n10827_11007.n9 a_n10827_11007.n8 13.2382
R89 a_n10827_11007.n8 a_n10827_11007.n1 5.76343
R90 a_n10827_11007.n1 a_n10827_11007.n0 5.54145
R91 VDD.n3968 VDD.n127 475.611
R92 VDD.n4539 VDD.n4169 475.611
R93 VDD.n4318 VDD.n4167 475.611
R94 VDD.n3970 VDD.n125 475.611
R95 VDD.n2169 VDD.n1211 475.611
R96 VDD.n2172 VDD.n2171 475.611
R97 VDD.n1697 VDD.n1388 475.611
R98 VDD.n1695 VDD.n1390 475.611
R99 VDD.n3742 VDD.n242 355.611
R100 VDD.n3709 VDD.n239 355.611
R101 VDD.n3111 VDD.n2897 355.611
R102 VDD.n3336 VDD.n601 355.611
R103 VDD.n2852 VDD.n632 355.611
R104 VDD.n2818 VDD.n2817 355.611
R105 VDD.n2431 VDD.n987 355.611
R106 VDD.n2465 VDD.n977 355.611
R107 VDD.n3688 VDD.n240 355.611
R108 VDD.n3745 VDD.n3744 355.611
R109 VDD.n3298 VDD.n3112 355.611
R110 VDD.n3334 VDD.n3113 355.611
R111 VDD.n2894 VDD.n621 355.611
R112 VDD.n2859 VDD.n620 355.611
R113 VDD.n2243 VDD.n996 355.611
R114 VDD.n997 VDD.n973 355.611
R115 VDD.n1154 VDD.t48 236.714
R116 VDD.n624 VDD.t116 236.714
R117 VDD.n253 VDD.t31 236.714
R118 VDD.n2900 VDD.t71 236.714
R119 VDD.n634 VDD.t83 236.714
R120 VDD.n1000 VDD.t111 236.714
R121 VDD.n230 VDD.t79 236.714
R122 VDD.n3120 VDD.t120 236.714
R123 VDD.n1490 VDD.t33 235.915
R124 VDD.n1556 VDD.t88 235.915
R125 VDD.n1586 VDD.t97 235.915
R126 VDD.n1641 VDD.t56 235.915
R127 VDD.n1419 VDD.t72 235.915
R128 VDD.n1975 VDD.t75 235.915
R129 VDD.n2035 VDD.t41 235.915
R130 VDD.n1189 VDD.t53 235.915
R131 VDD.n1164 VDD.t59 235.915
R132 VDD.n2004 VDD.t62 235.915
R133 VDD.n206 VDD.t49 235.915
R134 VDD.n3795 VDD.t100 235.915
R135 VDD.n4256 VDD.t91 235.915
R136 VDD.n4320 VDD.t94 235.915
R137 VDD.n4288 VDD.t103 235.915
R138 VDD.n4225 VDD.t106 235.915
R139 VDD.n4508 VDD.t37 235.915
R140 VDD.n150 VDD.t85 235.915
R141 VDD.n177 VDD.t65 235.915
R142 VDD.n3832 VDD.t112 235.915
R143 VDD.n1154 VDD.t45 223.453
R144 VDD.n624 VDD.t115 223.453
R145 VDD.n253 VDD.t29 223.453
R146 VDD.n2900 VDD.t68 223.453
R147 VDD.n634 VDD.t81 223.453
R148 VDD.n1000 VDD.t109 223.453
R149 VDD.n230 VDD.t78 223.453
R150 VDD.n3120 VDD.t118 223.453
R151 VDD.n4320 VDD.t95 198.272
R152 VDD.n177 VDD.t67 198.272
R153 VDD.n3832 VDD.t114 198.272
R154 VDD.n1490 VDD.t36 188.672
R155 VDD.n1556 VDD.t90 188.672
R156 VDD.n1586 VDD.t99 188.672
R157 VDD.n1641 VDD.t58 188.672
R158 VDD.n1419 VDD.t74 188.672
R159 VDD.n1975 VDD.t76 188.672
R160 VDD.n2035 VDD.t43 188.672
R161 VDD.n1189 VDD.t54 188.672
R162 VDD.n1164 VDD.t60 188.672
R163 VDD.n2004 VDD.t63 188.672
R164 VDD.n206 VDD.t52 188.672
R165 VDD.n3795 VDD.t102 188.672
R166 VDD.n4256 VDD.t92 188.672
R167 VDD.n4288 VDD.t104 188.672
R168 VDD.n4225 VDD.t107 188.672
R169 VDD.n4508 VDD.t39 188.672
R170 VDD.n150 VDD.t87 188.672
R171 VDD.n3690 VDD.n240 185
R172 VDD.n3743 VDD.n240 185
R173 VDD.n3692 VDD.n3691 185
R174 VDD.n3691 VDD.n238 185
R175 VDD.n3693 VDD.n261 185
R176 VDD.n3703 VDD.n261 185
R177 VDD.n3694 VDD.n269 185
R178 VDD.n269 VDD.n259 185
R179 VDD.n3696 VDD.n3695 185
R180 VDD.n3697 VDD.n3696 185
R181 VDD.n3668 VDD.n268 185
R182 VDD.n268 VDD.n265 185
R183 VDD.n3667 VDD.n3666 185
R184 VDD.n3666 VDD.n3665 185
R185 VDD.n271 VDD.n270 185
R186 VDD.n272 VDD.n271 185
R187 VDD.n3658 VDD.n3657 185
R188 VDD.n3659 VDD.n3658 185
R189 VDD.n3656 VDD.n281 185
R190 VDD.n281 VDD.n278 185
R191 VDD.n3655 VDD.n3654 185
R192 VDD.n3654 VDD.n3653 185
R193 VDD.n283 VDD.n282 185
R194 VDD.n292 VDD.n283 185
R195 VDD.n3646 VDD.n3645 185
R196 VDD.n3647 VDD.n3646 185
R197 VDD.n3644 VDD.n293 185
R198 VDD.n293 VDD.n289 185
R199 VDD.n3643 VDD.n3642 185
R200 VDD.n3642 VDD.n3641 185
R201 VDD.n295 VDD.n294 185
R202 VDD.n296 VDD.n295 185
R203 VDD.n3634 VDD.n3633 185
R204 VDD.n3635 VDD.n3634 185
R205 VDD.n3632 VDD.n305 185
R206 VDD.n305 VDD.n302 185
R207 VDD.n3631 VDD.n3630 185
R208 VDD.n3630 VDD.n3629 185
R209 VDD.n307 VDD.n306 185
R210 VDD.n308 VDD.n307 185
R211 VDD.n3622 VDD.n3621 185
R212 VDD.n3623 VDD.n3622 185
R213 VDD.n3620 VDD.n317 185
R214 VDD.n317 VDD.n314 185
R215 VDD.n3619 VDD.n3618 185
R216 VDD.n3618 VDD.n3617 185
R217 VDD.n319 VDD.n318 185
R218 VDD.n320 VDD.n319 185
R219 VDD.n3610 VDD.n3609 185
R220 VDD.n3611 VDD.n3610 185
R221 VDD.n3608 VDD.n329 185
R222 VDD.n329 VDD.n326 185
R223 VDD.n3607 VDD.n3606 185
R224 VDD.n3606 VDD.n3605 185
R225 VDD.n331 VDD.n330 185
R226 VDD.n340 VDD.n331 185
R227 VDD.n3598 VDD.n3597 185
R228 VDD.n3599 VDD.n3598 185
R229 VDD.n3596 VDD.n341 185
R230 VDD.n341 VDD.n337 185
R231 VDD.n3595 VDD.n3594 185
R232 VDD.n3594 VDD.n3593 185
R233 VDD.n343 VDD.n342 185
R234 VDD.n344 VDD.n343 185
R235 VDD.n3586 VDD.n3585 185
R236 VDD.n3587 VDD.n3586 185
R237 VDD.n3584 VDD.n353 185
R238 VDD.n353 VDD.n350 185
R239 VDD.n3583 VDD.n3582 185
R240 VDD.n3582 VDD.n3581 185
R241 VDD.n355 VDD.n354 185
R242 VDD.n356 VDD.n355 185
R243 VDD.n3574 VDD.n3573 185
R244 VDD.n3575 VDD.n3574 185
R245 VDD.n3572 VDD.n365 185
R246 VDD.n365 VDD.n362 185
R247 VDD.n3571 VDD.n3570 185
R248 VDD.n3570 VDD.n3569 185
R249 VDD.n367 VDD.n366 185
R250 VDD.n368 VDD.n367 185
R251 VDD.n3562 VDD.n3561 185
R252 VDD.n3563 VDD.n3562 185
R253 VDD.n3560 VDD.n377 185
R254 VDD.n377 VDD.n374 185
R255 VDD.n3559 VDD.n3558 185
R256 VDD.n3558 VDD.n3557 185
R257 VDD.n379 VDD.n378 185
R258 VDD.n380 VDD.n379 185
R259 VDD.n3550 VDD.n3549 185
R260 VDD.n3551 VDD.n3550 185
R261 VDD.n3548 VDD.n389 185
R262 VDD.n389 VDD.n386 185
R263 VDD.n3547 VDD.n3546 185
R264 VDD.n3546 VDD.n3545 185
R265 VDD.n391 VDD.n390 185
R266 VDD.n392 VDD.n391 185
R267 VDD.n3538 VDD.n3537 185
R268 VDD.n3539 VDD.n3538 185
R269 VDD.n3536 VDD.n401 185
R270 VDD.n401 VDD.n398 185
R271 VDD.n3535 VDD.n3534 185
R272 VDD.n3534 VDD.n3533 185
R273 VDD.n403 VDD.n402 185
R274 VDD.n404 VDD.n403 185
R275 VDD.n3526 VDD.n3525 185
R276 VDD.n3527 VDD.n3526 185
R277 VDD.n3524 VDD.n412 185
R278 VDD.n418 VDD.n412 185
R279 VDD.n3523 VDD.n3522 185
R280 VDD.n3522 VDD.n3521 185
R281 VDD.n414 VDD.n413 185
R282 VDD.n415 VDD.n414 185
R283 VDD.n3514 VDD.n3513 185
R284 VDD.n3515 VDD.n3514 185
R285 VDD.n3512 VDD.n425 185
R286 VDD.n425 VDD.n422 185
R287 VDD.n3511 VDD.n3510 185
R288 VDD.n3510 VDD.n3509 185
R289 VDD.n427 VDD.n426 185
R290 VDD.n428 VDD.n427 185
R291 VDD.n3502 VDD.n3501 185
R292 VDD.n3503 VDD.n3502 185
R293 VDD.n3500 VDD.n437 185
R294 VDD.n437 VDD.n434 185
R295 VDD.n3499 VDD.n3498 185
R296 VDD.n3498 VDD.n3497 185
R297 VDD.n439 VDD.n438 185
R298 VDD.n440 VDD.n439 185
R299 VDD.n3490 VDD.n3489 185
R300 VDD.n3491 VDD.n3490 185
R301 VDD.n3488 VDD.n449 185
R302 VDD.n449 VDD.n446 185
R303 VDD.n3487 VDD.n3486 185
R304 VDD.n3486 VDD.n3485 185
R305 VDD.n451 VDD.n450 185
R306 VDD.n460 VDD.n451 185
R307 VDD.n3478 VDD.n3477 185
R308 VDD.n3479 VDD.n3478 185
R309 VDD.n3476 VDD.n461 185
R310 VDD.n461 VDD.n457 185
R311 VDD.n3475 VDD.n3474 185
R312 VDD.n3474 VDD.n3473 185
R313 VDD.n463 VDD.n462 185
R314 VDD.n472 VDD.n463 185
R315 VDD.n3466 VDD.n3465 185
R316 VDD.n3467 VDD.n3466 185
R317 VDD.n3464 VDD.n473 185
R318 VDD.n473 VDD.n469 185
R319 VDD.n3463 VDD.n3462 185
R320 VDD.n3462 VDD.n3461 185
R321 VDD.n475 VDD.n474 185
R322 VDD.n476 VDD.n475 185
R323 VDD.n3454 VDD.n3453 185
R324 VDD.n3455 VDD.n3454 185
R325 VDD.n3452 VDD.n485 185
R326 VDD.n485 VDD.n482 185
R327 VDD.n3451 VDD.n3450 185
R328 VDD.n3450 VDD.n3449 185
R329 VDD.n487 VDD.n486 185
R330 VDD.n488 VDD.n487 185
R331 VDD.n3442 VDD.n3441 185
R332 VDD.n3443 VDD.n3442 185
R333 VDD.n3440 VDD.n497 185
R334 VDD.n497 VDD.n494 185
R335 VDD.n3439 VDD.n3438 185
R336 VDD.n3438 VDD.n3437 185
R337 VDD.n499 VDD.n498 185
R338 VDD.n500 VDD.n499 185
R339 VDD.n3430 VDD.n3429 185
R340 VDD.n3431 VDD.n3430 185
R341 VDD.n3428 VDD.n508 185
R342 VDD.n514 VDD.n508 185
R343 VDD.n3427 VDD.n3426 185
R344 VDD.n3426 VDD.n3425 185
R345 VDD.n510 VDD.n509 185
R346 VDD.n511 VDD.n510 185
R347 VDD.n3418 VDD.n3417 185
R348 VDD.n3419 VDD.n3418 185
R349 VDD.n3416 VDD.n521 185
R350 VDD.n521 VDD.n518 185
R351 VDD.n3415 VDD.n3414 185
R352 VDD.n3414 VDD.n3413 185
R353 VDD.n523 VDD.n522 185
R354 VDD.n524 VDD.n523 185
R355 VDD.n3406 VDD.n3405 185
R356 VDD.n3407 VDD.n3406 185
R357 VDD.n3404 VDD.n533 185
R358 VDD.n533 VDD.n530 185
R359 VDD.n3403 VDD.n3402 185
R360 VDD.n3402 VDD.n3401 185
R361 VDD.n535 VDD.n534 185
R362 VDD.n536 VDD.n535 185
R363 VDD.n3394 VDD.n3393 185
R364 VDD.n3395 VDD.n3394 185
R365 VDD.n3392 VDD.n545 185
R366 VDD.n545 VDD.n542 185
R367 VDD.n3391 VDD.n3390 185
R368 VDD.n3390 VDD.n3389 185
R369 VDD.n547 VDD.n546 185
R370 VDD.n548 VDD.n547 185
R371 VDD.n3382 VDD.n3381 185
R372 VDD.n3383 VDD.n3382 185
R373 VDD.n3380 VDD.n557 185
R374 VDD.n557 VDD.n554 185
R375 VDD.n3379 VDD.n3378 185
R376 VDD.n3378 VDD.n3377 185
R377 VDD.n559 VDD.n558 185
R378 VDD.n560 VDD.n559 185
R379 VDD.n3370 VDD.n3369 185
R380 VDD.n3371 VDD.n3370 185
R381 VDD.n3368 VDD.n569 185
R382 VDD.n569 VDD.n566 185
R383 VDD.n3367 VDD.n3366 185
R384 VDD.n3366 VDD.n3365 185
R385 VDD.n571 VDD.n570 185
R386 VDD.n572 VDD.n571 185
R387 VDD.n3358 VDD.n3357 185
R388 VDD.n3359 VDD.n3358 185
R389 VDD.n3356 VDD.n581 185
R390 VDD.n581 VDD.n578 185
R391 VDD.n3355 VDD.n3354 185
R392 VDD.n3354 VDD.n3353 185
R393 VDD.n583 VDD.n582 185
R394 VDD.n584 VDD.n583 185
R395 VDD.n3346 VDD.n3345 185
R396 VDD.n3347 VDD.n3346 185
R397 VDD.n3344 VDD.n593 185
R398 VDD.n593 VDD.n590 185
R399 VDD.n3343 VDD.n3342 185
R400 VDD.n3342 VDD.n3341 185
R401 VDD.n595 VDD.n594 185
R402 VDD.n596 VDD.n595 185
R403 VDD.n3334 VDD.n3333 185
R404 VDD.n3335 VDD.n3334 185
R405 VDD.n3332 VDD.n3113 185
R406 VDD.n3331 VDD.n3330 185
R407 VDD.n3328 VDD.n3114 185
R408 VDD.n3326 VDD.n3325 185
R409 VDD.n3324 VDD.n3115 185
R410 VDD.n3323 VDD.n3322 185
R411 VDD.n3320 VDD.n3116 185
R412 VDD.n3318 VDD.n3317 185
R413 VDD.n3316 VDD.n3117 185
R414 VDD.n3315 VDD.n3314 185
R415 VDD.n3312 VDD.n3118 185
R416 VDD.n3310 VDD.n3309 185
R417 VDD.n3308 VDD.n3119 185
R418 VDD.n3307 VDD.n3306 185
R419 VDD.n3304 VDD.n3122 185
R420 VDD.n3302 VDD.n3301 185
R421 VDD.n3300 VDD.n3123 185
R422 VDD.n3299 VDD.n3298 185
R423 VDD.n3746 VDD.n3745 185
R424 VDD.n3747 VDD.n234 185
R425 VDD.n3749 VDD.n3748 185
R426 VDD.n3751 VDD.n232 185
R427 VDD.n3753 VDD.n3752 185
R428 VDD.n3754 VDD.n229 185
R429 VDD.n3756 VDD.n3755 185
R430 VDD.n3758 VDD.n226 185
R431 VDD.n3760 VDD.n3759 185
R432 VDD.n3674 VDD.n225 185
R433 VDD.n3676 VDD.n3675 185
R434 VDD.n3678 VDD.n3672 185
R435 VDD.n3680 VDD.n3679 185
R436 VDD.n3681 VDD.n3671 185
R437 VDD.n3683 VDD.n3682 185
R438 VDD.n3685 VDD.n3670 185
R439 VDD.n3686 VDD.n3669 185
R440 VDD.n3689 VDD.n3688 185
R441 VDD.n3744 VDD.n235 185
R442 VDD.n3744 VDD.n3743 185
R443 VDD.n3124 VDD.n237 185
R444 VDD.n238 VDD.n237 185
R445 VDD.n3125 VDD.n260 185
R446 VDD.n3703 VDD.n260 185
R447 VDD.n3127 VDD.n3126 185
R448 VDD.n3126 VDD.n259 185
R449 VDD.n3128 VDD.n267 185
R450 VDD.n3697 VDD.n267 185
R451 VDD.n3130 VDD.n3129 185
R452 VDD.n3129 VDD.n265 185
R453 VDD.n3131 VDD.n274 185
R454 VDD.n3665 VDD.n274 185
R455 VDD.n3133 VDD.n3132 185
R456 VDD.n3132 VDD.n272 185
R457 VDD.n3134 VDD.n280 185
R458 VDD.n3659 VDD.n280 185
R459 VDD.n3136 VDD.n3135 185
R460 VDD.n3135 VDD.n278 185
R461 VDD.n3137 VDD.n285 185
R462 VDD.n3653 VDD.n285 185
R463 VDD.n3139 VDD.n3138 185
R464 VDD.n3138 VDD.n292 185
R465 VDD.n3140 VDD.n291 185
R466 VDD.n3647 VDD.n291 185
R467 VDD.n3142 VDD.n3141 185
R468 VDD.n3141 VDD.n289 185
R469 VDD.n3143 VDD.n298 185
R470 VDD.n3641 VDD.n298 185
R471 VDD.n3145 VDD.n3144 185
R472 VDD.n3144 VDD.n296 185
R473 VDD.n3146 VDD.n304 185
R474 VDD.n3635 VDD.n304 185
R475 VDD.n3148 VDD.n3147 185
R476 VDD.n3147 VDD.n302 185
R477 VDD.n3149 VDD.n310 185
R478 VDD.n3629 VDD.n310 185
R479 VDD.n3151 VDD.n3150 185
R480 VDD.n3150 VDD.n308 185
R481 VDD.n3152 VDD.n316 185
R482 VDD.n3623 VDD.n316 185
R483 VDD.n3154 VDD.n3153 185
R484 VDD.n3153 VDD.n314 185
R485 VDD.n3155 VDD.n322 185
R486 VDD.n3617 VDD.n322 185
R487 VDD.n3157 VDD.n3156 185
R488 VDD.n3156 VDD.n320 185
R489 VDD.n3158 VDD.n328 185
R490 VDD.n3611 VDD.n328 185
R491 VDD.n3160 VDD.n3159 185
R492 VDD.n3159 VDD.n326 185
R493 VDD.n3161 VDD.n333 185
R494 VDD.n3605 VDD.n333 185
R495 VDD.n3163 VDD.n3162 185
R496 VDD.n3162 VDD.n340 185
R497 VDD.n3164 VDD.n339 185
R498 VDD.n3599 VDD.n339 185
R499 VDD.n3166 VDD.n3165 185
R500 VDD.n3165 VDD.n337 185
R501 VDD.n3167 VDD.n346 185
R502 VDD.n3593 VDD.n346 185
R503 VDD.n3169 VDD.n3168 185
R504 VDD.n3168 VDD.n344 185
R505 VDD.n3170 VDD.n352 185
R506 VDD.n3587 VDD.n352 185
R507 VDD.n3172 VDD.n3171 185
R508 VDD.n3171 VDD.n350 185
R509 VDD.n3173 VDD.n358 185
R510 VDD.n3581 VDD.n358 185
R511 VDD.n3175 VDD.n3174 185
R512 VDD.n3174 VDD.n356 185
R513 VDD.n3176 VDD.n364 185
R514 VDD.n3575 VDD.n364 185
R515 VDD.n3178 VDD.n3177 185
R516 VDD.n3177 VDD.n362 185
R517 VDD.n3179 VDD.n370 185
R518 VDD.n3569 VDD.n370 185
R519 VDD.n3181 VDD.n3180 185
R520 VDD.n3180 VDD.n368 185
R521 VDD.n3182 VDD.n376 185
R522 VDD.n3563 VDD.n376 185
R523 VDD.n3184 VDD.n3183 185
R524 VDD.n3183 VDD.n374 185
R525 VDD.n3185 VDD.n382 185
R526 VDD.n3557 VDD.n382 185
R527 VDD.n3187 VDD.n3186 185
R528 VDD.n3186 VDD.n380 185
R529 VDD.n3188 VDD.n388 185
R530 VDD.n3551 VDD.n388 185
R531 VDD.n3190 VDD.n3189 185
R532 VDD.n3189 VDD.n386 185
R533 VDD.n3191 VDD.n394 185
R534 VDD.n3545 VDD.n394 185
R535 VDD.n3193 VDD.n3192 185
R536 VDD.n3192 VDD.n392 185
R537 VDD.n3194 VDD.n400 185
R538 VDD.n3539 VDD.n400 185
R539 VDD.n3196 VDD.n3195 185
R540 VDD.n3195 VDD.n398 185
R541 VDD.n3197 VDD.n406 185
R542 VDD.n3533 VDD.n406 185
R543 VDD.n3199 VDD.n3198 185
R544 VDD.n3198 VDD.n404 185
R545 VDD.n3200 VDD.n411 185
R546 VDD.n3527 VDD.n411 185
R547 VDD.n3202 VDD.n3201 185
R548 VDD.n3201 VDD.n418 185
R549 VDD.n3203 VDD.n417 185
R550 VDD.n3521 VDD.n417 185
R551 VDD.n3205 VDD.n3204 185
R552 VDD.n3204 VDD.n415 185
R553 VDD.n3206 VDD.n424 185
R554 VDD.n3515 VDD.n424 185
R555 VDD.n3208 VDD.n3207 185
R556 VDD.n3207 VDD.n422 185
R557 VDD.n3209 VDD.n430 185
R558 VDD.n3509 VDD.n430 185
R559 VDD.n3211 VDD.n3210 185
R560 VDD.n3210 VDD.n428 185
R561 VDD.n3212 VDD.n436 185
R562 VDD.n3503 VDD.n436 185
R563 VDD.n3214 VDD.n3213 185
R564 VDD.n3213 VDD.n434 185
R565 VDD.n3215 VDD.n442 185
R566 VDD.n3497 VDD.n442 185
R567 VDD.n3217 VDD.n3216 185
R568 VDD.n3216 VDD.n440 185
R569 VDD.n3218 VDD.n448 185
R570 VDD.n3491 VDD.n448 185
R571 VDD.n3220 VDD.n3219 185
R572 VDD.n3219 VDD.n446 185
R573 VDD.n3221 VDD.n453 185
R574 VDD.n3485 VDD.n453 185
R575 VDD.n3223 VDD.n3222 185
R576 VDD.n3222 VDD.n460 185
R577 VDD.n3224 VDD.n459 185
R578 VDD.n3479 VDD.n459 185
R579 VDD.n3226 VDD.n3225 185
R580 VDD.n3225 VDD.n457 185
R581 VDD.n3227 VDD.n465 185
R582 VDD.n3473 VDD.n465 185
R583 VDD.n3229 VDD.n3228 185
R584 VDD.n3228 VDD.n472 185
R585 VDD.n3230 VDD.n471 185
R586 VDD.n3467 VDD.n471 185
R587 VDD.n3232 VDD.n3231 185
R588 VDD.n3231 VDD.n469 185
R589 VDD.n3233 VDD.n478 185
R590 VDD.n3461 VDD.n478 185
R591 VDD.n3235 VDD.n3234 185
R592 VDD.n3234 VDD.n476 185
R593 VDD.n3236 VDD.n484 185
R594 VDD.n3455 VDD.n484 185
R595 VDD.n3238 VDD.n3237 185
R596 VDD.n3237 VDD.n482 185
R597 VDD.n3239 VDD.n490 185
R598 VDD.n3449 VDD.n490 185
R599 VDD.n3241 VDD.n3240 185
R600 VDD.n3240 VDD.n488 185
R601 VDD.n3242 VDD.n496 185
R602 VDD.n3443 VDD.n496 185
R603 VDD.n3244 VDD.n3243 185
R604 VDD.n3243 VDD.n494 185
R605 VDD.n3245 VDD.n502 185
R606 VDD.n3437 VDD.n502 185
R607 VDD.n3247 VDD.n3246 185
R608 VDD.n3246 VDD.n500 185
R609 VDD.n3248 VDD.n507 185
R610 VDD.n3431 VDD.n507 185
R611 VDD.n3250 VDD.n3249 185
R612 VDD.n3249 VDD.n514 185
R613 VDD.n3251 VDD.n513 185
R614 VDD.n3425 VDD.n513 185
R615 VDD.n3253 VDD.n3252 185
R616 VDD.n3252 VDD.n511 185
R617 VDD.n3254 VDD.n520 185
R618 VDD.n3419 VDD.n520 185
R619 VDD.n3256 VDD.n3255 185
R620 VDD.n3255 VDD.n518 185
R621 VDD.n3257 VDD.n526 185
R622 VDD.n3413 VDD.n526 185
R623 VDD.n3259 VDD.n3258 185
R624 VDD.n3258 VDD.n524 185
R625 VDD.n3260 VDD.n532 185
R626 VDD.n3407 VDD.n532 185
R627 VDD.n3262 VDD.n3261 185
R628 VDD.n3261 VDD.n530 185
R629 VDD.n3263 VDD.n538 185
R630 VDD.n3401 VDD.n538 185
R631 VDD.n3265 VDD.n3264 185
R632 VDD.n3264 VDD.n536 185
R633 VDD.n3266 VDD.n544 185
R634 VDD.n3395 VDD.n544 185
R635 VDD.n3268 VDD.n3267 185
R636 VDD.n3267 VDD.n542 185
R637 VDD.n3269 VDD.n550 185
R638 VDD.n3389 VDD.n550 185
R639 VDD.n3271 VDD.n3270 185
R640 VDD.n3270 VDD.n548 185
R641 VDD.n3272 VDD.n556 185
R642 VDD.n3383 VDD.n556 185
R643 VDD.n3274 VDD.n3273 185
R644 VDD.n3273 VDD.n554 185
R645 VDD.n3275 VDD.n562 185
R646 VDD.n3377 VDD.n562 185
R647 VDD.n3277 VDD.n3276 185
R648 VDD.n3276 VDD.n560 185
R649 VDD.n3278 VDD.n568 185
R650 VDD.n3371 VDD.n568 185
R651 VDD.n3280 VDD.n3279 185
R652 VDD.n3279 VDD.n566 185
R653 VDD.n3281 VDD.n574 185
R654 VDD.n3365 VDD.n574 185
R655 VDD.n3283 VDD.n3282 185
R656 VDD.n3282 VDD.n572 185
R657 VDD.n3284 VDD.n580 185
R658 VDD.n3359 VDD.n580 185
R659 VDD.n3286 VDD.n3285 185
R660 VDD.n3285 VDD.n578 185
R661 VDD.n3287 VDD.n586 185
R662 VDD.n3353 VDD.n586 185
R663 VDD.n3289 VDD.n3288 185
R664 VDD.n3288 VDD.n584 185
R665 VDD.n3290 VDD.n592 185
R666 VDD.n3347 VDD.n592 185
R667 VDD.n3292 VDD.n3291 185
R668 VDD.n3291 VDD.n590 185
R669 VDD.n3293 VDD.n598 185
R670 VDD.n3341 VDD.n598 185
R671 VDD.n3295 VDD.n3294 185
R672 VDD.n3294 VDD.n596 185
R673 VDD.n3296 VDD.n3112 185
R674 VDD.n3335 VDD.n3112 185
R675 VDD.n2854 VDD.n632 185
R676 VDD.n632 VDD.n602 185
R677 VDD.n2856 VDD.n2855 185
R678 VDD.n2857 VDD.n2856 185
R679 VDD.n633 VDD.n631 185
R680 VDD.n631 VDD.n628 185
R681 VDD.n2810 VDD.n2809 185
R682 VDD.n2811 VDD.n2810 185
R683 VDD.n2808 VDD.n641 185
R684 VDD.n641 VDD.n638 185
R685 VDD.n2807 VDD.n2806 185
R686 VDD.n2806 VDD.n2805 185
R687 VDD.n643 VDD.n642 185
R688 VDD.n644 VDD.n643 185
R689 VDD.n2793 VDD.n2792 185
R690 VDD.n2794 VDD.n2793 185
R691 VDD.n2791 VDD.n654 185
R692 VDD.n654 VDD.n651 185
R693 VDD.n2790 VDD.n2789 185
R694 VDD.n2789 VDD.n2788 185
R695 VDD.n656 VDD.n655 185
R696 VDD.n657 VDD.n656 185
R697 VDD.n2781 VDD.n2780 185
R698 VDD.n2782 VDD.n2781 185
R699 VDD.n2779 VDD.n666 185
R700 VDD.n666 VDD.n663 185
R701 VDD.n2778 VDD.n2777 185
R702 VDD.n2777 VDD.n2776 185
R703 VDD.n668 VDD.n667 185
R704 VDD.n669 VDD.n668 185
R705 VDD.n2769 VDD.n2768 185
R706 VDD.n2770 VDD.n2769 185
R707 VDD.n2767 VDD.n678 185
R708 VDD.n678 VDD.n675 185
R709 VDD.n2766 VDD.n2765 185
R710 VDD.n2765 VDD.n2764 185
R711 VDD.n680 VDD.n679 185
R712 VDD.n681 VDD.n680 185
R713 VDD.n2757 VDD.n2756 185
R714 VDD.n2758 VDD.n2757 185
R715 VDD.n2755 VDD.n690 185
R716 VDD.n690 VDD.n687 185
R717 VDD.n2754 VDD.n2753 185
R718 VDD.n2753 VDD.n2752 185
R719 VDD.n692 VDD.n691 185
R720 VDD.n693 VDD.n692 185
R721 VDD.n2745 VDD.n2744 185
R722 VDD.n2746 VDD.n2745 185
R723 VDD.n2743 VDD.n702 185
R724 VDD.n702 VDD.n699 185
R725 VDD.n2742 VDD.n2741 185
R726 VDD.n2741 VDD.n2740 185
R727 VDD.n704 VDD.n703 185
R728 VDD.n705 VDD.n704 185
R729 VDD.n2733 VDD.n2732 185
R730 VDD.n2734 VDD.n2733 185
R731 VDD.n2731 VDD.n714 185
R732 VDD.n714 VDD.n711 185
R733 VDD.n2730 VDD.n2729 185
R734 VDD.n2729 VDD.n2728 185
R735 VDD.n716 VDD.n715 185
R736 VDD.n717 VDD.n716 185
R737 VDD.n2721 VDD.n2720 185
R738 VDD.n2722 VDD.n2721 185
R739 VDD.n2719 VDD.n725 185
R740 VDD.n731 VDD.n725 185
R741 VDD.n2718 VDD.n2717 185
R742 VDD.n2717 VDD.n2716 185
R743 VDD.n727 VDD.n726 185
R744 VDD.n728 VDD.n727 185
R745 VDD.n2709 VDD.n2708 185
R746 VDD.n2710 VDD.n2709 185
R747 VDD.n2707 VDD.n738 185
R748 VDD.n738 VDD.n735 185
R749 VDD.n2706 VDD.n2705 185
R750 VDD.n2705 VDD.n2704 185
R751 VDD.n740 VDD.n739 185
R752 VDD.n741 VDD.n740 185
R753 VDD.n2697 VDD.n2696 185
R754 VDD.n2698 VDD.n2697 185
R755 VDD.n2695 VDD.n750 185
R756 VDD.n750 VDD.n747 185
R757 VDD.n2694 VDD.n2693 185
R758 VDD.n2693 VDD.n2692 185
R759 VDD.n752 VDD.n751 185
R760 VDD.n753 VDD.n752 185
R761 VDD.n2685 VDD.n2684 185
R762 VDD.n2686 VDD.n2685 185
R763 VDD.n2683 VDD.n762 185
R764 VDD.n762 VDD.n759 185
R765 VDD.n2682 VDD.n2681 185
R766 VDD.n2681 VDD.n2680 185
R767 VDD.n764 VDD.n763 185
R768 VDD.n773 VDD.n764 185
R769 VDD.n2673 VDD.n2672 185
R770 VDD.n2674 VDD.n2673 185
R771 VDD.n2671 VDD.n774 185
R772 VDD.n774 VDD.n770 185
R773 VDD.n2670 VDD.n2669 185
R774 VDD.n2669 VDD.n2668 185
R775 VDD.n776 VDD.n775 185
R776 VDD.n785 VDD.n776 185
R777 VDD.n2661 VDD.n2660 185
R778 VDD.n2662 VDD.n2661 185
R779 VDD.n2659 VDD.n786 185
R780 VDD.n786 VDD.n782 185
R781 VDD.n2658 VDD.n2657 185
R782 VDD.n2657 VDD.n2656 185
R783 VDD.n788 VDD.n787 185
R784 VDD.n789 VDD.n788 185
R785 VDD.n2649 VDD.n2648 185
R786 VDD.n2650 VDD.n2649 185
R787 VDD.n2647 VDD.n798 185
R788 VDD.n798 VDD.n795 185
R789 VDD.n2646 VDD.n2645 185
R790 VDD.n2645 VDD.n2644 185
R791 VDD.n800 VDD.n799 185
R792 VDD.n801 VDD.n800 185
R793 VDD.n2637 VDD.n2636 185
R794 VDD.n2638 VDD.n2637 185
R795 VDD.n2635 VDD.n810 185
R796 VDD.n810 VDD.n807 185
R797 VDD.n2634 VDD.n2633 185
R798 VDD.n2633 VDD.n2632 185
R799 VDD.n812 VDD.n811 185
R800 VDD.n813 VDD.n812 185
R801 VDD.n2625 VDD.n2624 185
R802 VDD.n2626 VDD.n2625 185
R803 VDD.n2623 VDD.n821 185
R804 VDD.n827 VDD.n821 185
R805 VDD.n2622 VDD.n2621 185
R806 VDD.n2621 VDD.n2620 185
R807 VDD.n823 VDD.n822 185
R808 VDD.n824 VDD.n823 185
R809 VDD.n2613 VDD.n2612 185
R810 VDD.n2614 VDD.n2613 185
R811 VDD.n2611 VDD.n834 185
R812 VDD.n834 VDD.n831 185
R813 VDD.n2610 VDD.n2609 185
R814 VDD.n2609 VDD.n2608 185
R815 VDD.n836 VDD.n835 185
R816 VDD.n837 VDD.n836 185
R817 VDD.n2601 VDD.n2600 185
R818 VDD.n2602 VDD.n2601 185
R819 VDD.n2599 VDD.n846 185
R820 VDD.n846 VDD.n843 185
R821 VDD.n2598 VDD.n2597 185
R822 VDD.n2597 VDD.n2596 185
R823 VDD.n848 VDD.n847 185
R824 VDD.n849 VDD.n848 185
R825 VDD.n2589 VDD.n2588 185
R826 VDD.n2590 VDD.n2589 185
R827 VDD.n2587 VDD.n858 185
R828 VDD.n858 VDD.n855 185
R829 VDD.n2586 VDD.n2585 185
R830 VDD.n2585 VDD.n2584 185
R831 VDD.n860 VDD.n859 185
R832 VDD.n861 VDD.n860 185
R833 VDD.n2577 VDD.n2576 185
R834 VDD.n2578 VDD.n2577 185
R835 VDD.n2575 VDD.n870 185
R836 VDD.n870 VDD.n867 185
R837 VDD.n2574 VDD.n2573 185
R838 VDD.n2573 VDD.n2572 185
R839 VDD.n872 VDD.n871 185
R840 VDD.n873 VDD.n872 185
R841 VDD.n2565 VDD.n2564 185
R842 VDD.n2566 VDD.n2565 185
R843 VDD.n2563 VDD.n882 185
R844 VDD.n882 VDD.n879 185
R845 VDD.n2562 VDD.n2561 185
R846 VDD.n2561 VDD.n2560 185
R847 VDD.n884 VDD.n883 185
R848 VDD.n885 VDD.n884 185
R849 VDD.n2553 VDD.n2552 185
R850 VDD.n2554 VDD.n2553 185
R851 VDD.n2551 VDD.n894 185
R852 VDD.n894 VDD.n891 185
R853 VDD.n2550 VDD.n2549 185
R854 VDD.n2549 VDD.n2548 185
R855 VDD.n896 VDD.n895 185
R856 VDD.n905 VDD.n896 185
R857 VDD.n2541 VDD.n2540 185
R858 VDD.n2542 VDD.n2541 185
R859 VDD.n2539 VDD.n906 185
R860 VDD.n906 VDD.n902 185
R861 VDD.n2538 VDD.n2537 185
R862 VDD.n2537 VDD.n2536 185
R863 VDD.n908 VDD.n907 185
R864 VDD.n909 VDD.n908 185
R865 VDD.n2529 VDD.n2528 185
R866 VDD.n2530 VDD.n2529 185
R867 VDD.n2527 VDD.n918 185
R868 VDD.n918 VDD.n915 185
R869 VDD.n2526 VDD.n2525 185
R870 VDD.n2525 VDD.n2524 185
R871 VDD.n920 VDD.n919 185
R872 VDD.n921 VDD.n920 185
R873 VDD.n2517 VDD.n2516 185
R874 VDD.n2518 VDD.n2517 185
R875 VDD.n2515 VDD.n930 185
R876 VDD.n930 VDD.n927 185
R877 VDD.n2514 VDD.n2513 185
R878 VDD.n2513 VDD.n2512 185
R879 VDD.n932 VDD.n931 185
R880 VDD.n933 VDD.n932 185
R881 VDD.n2505 VDD.n2504 185
R882 VDD.n2506 VDD.n2505 185
R883 VDD.n2503 VDD.n942 185
R884 VDD.n942 VDD.n939 185
R885 VDD.n2502 VDD.n2501 185
R886 VDD.n2501 VDD.n2500 185
R887 VDD.n944 VDD.n943 185
R888 VDD.n2415 VDD.n944 185
R889 VDD.n2493 VDD.n2492 185
R890 VDD.n2494 VDD.n2493 185
R891 VDD.n2491 VDD.n953 185
R892 VDD.n953 VDD.n950 185
R893 VDD.n2490 VDD.n2489 185
R894 VDD.n2489 VDD.n2488 185
R895 VDD.n955 VDD.n954 185
R896 VDD.n956 VDD.n955 185
R897 VDD.n2481 VDD.n2480 185
R898 VDD.n2482 VDD.n2481 185
R899 VDD.n2479 VDD.n965 185
R900 VDD.n965 VDD.n962 185
R901 VDD.n2478 VDD.n2477 185
R902 VDD.n2477 VDD.n2476 185
R903 VDD.n967 VDD.n966 185
R904 VDD.n968 VDD.n967 185
R905 VDD.n2469 VDD.n2468 185
R906 VDD.n2470 VDD.n2469 185
R907 VDD.n2467 VDD.n977 185
R908 VDD.n977 VDD.n974 185
R909 VDD.n2466 VDD.n2465 185
R910 VDD.n979 VDD.n978 185
R911 VDD.n2462 VDD.n2461 185
R912 VDD.n2463 VDD.n2462 185
R913 VDD.n2460 VDD.n998 185
R914 VDD.n2459 VDD.n2458 185
R915 VDD.n2457 VDD.n2456 185
R916 VDD.n2455 VDD.n2454 185
R917 VDD.n2453 VDD.n2452 185
R918 VDD.n2451 VDD.n2450 185
R919 VDD.n2449 VDD.n2448 185
R920 VDD.n2447 VDD.n2446 185
R921 VDD.n2445 VDD.n2444 185
R922 VDD.n2443 VDD.n2442 185
R923 VDD.n2441 VDD.n2440 185
R924 VDD.n2439 VDD.n2438 185
R925 VDD.n2437 VDD.n2436 185
R926 VDD.n2435 VDD.n2434 185
R927 VDD.n2433 VDD.n987 185
R928 VDD.n2463 VDD.n987 185
R929 VDD.n2819 VDD.n2818 185
R930 VDD.n2821 VDD.n2820 185
R931 VDD.n2823 VDD.n2822 185
R932 VDD.n2825 VDD.n2824 185
R933 VDD.n2827 VDD.n2826 185
R934 VDD.n2829 VDD.n2828 185
R935 VDD.n2831 VDD.n2830 185
R936 VDD.n2833 VDD.n2832 185
R937 VDD.n2835 VDD.n2834 185
R938 VDD.n2837 VDD.n2836 185
R939 VDD.n2839 VDD.n2838 185
R940 VDD.n2841 VDD.n2840 185
R941 VDD.n2843 VDD.n2842 185
R942 VDD.n2845 VDD.n2844 185
R943 VDD.n2847 VDD.n2846 185
R944 VDD.n2849 VDD.n2848 185
R945 VDD.n2851 VDD.n2850 185
R946 VDD.n2853 VDD.n2852 185
R947 VDD.n2817 VDD.n2816 185
R948 VDD.n2817 VDD.n602 185
R949 VDD.n2815 VDD.n629 185
R950 VDD.n2857 VDD.n629 185
R951 VDD.n2814 VDD.n2813 185
R952 VDD.n2813 VDD.n628 185
R953 VDD.n2812 VDD.n636 185
R954 VDD.n2812 VDD.n2811 185
R955 VDD.n1002 VDD.n637 185
R956 VDD.n638 VDD.n637 185
R957 VDD.n1003 VDD.n645 185
R958 VDD.n2805 VDD.n645 185
R959 VDD.n1005 VDD.n1004 185
R960 VDD.n1004 VDD.n644 185
R961 VDD.n1006 VDD.n652 185
R962 VDD.n2794 VDD.n652 185
R963 VDD.n1008 VDD.n1007 185
R964 VDD.n1007 VDD.n651 185
R965 VDD.n1009 VDD.n658 185
R966 VDD.n2788 VDD.n658 185
R967 VDD.n1011 VDD.n1010 185
R968 VDD.n1010 VDD.n657 185
R969 VDD.n1012 VDD.n664 185
R970 VDD.n2782 VDD.n664 185
R971 VDD.n1014 VDD.n1013 185
R972 VDD.n1013 VDD.n663 185
R973 VDD.n1015 VDD.n670 185
R974 VDD.n2776 VDD.n670 185
R975 VDD.n1017 VDD.n1016 185
R976 VDD.n1016 VDD.n669 185
R977 VDD.n1018 VDD.n676 185
R978 VDD.n2770 VDD.n676 185
R979 VDD.n1020 VDD.n1019 185
R980 VDD.n1019 VDD.n675 185
R981 VDD.n1021 VDD.n682 185
R982 VDD.n2764 VDD.n682 185
R983 VDD.n1023 VDD.n1022 185
R984 VDD.n1022 VDD.n681 185
R985 VDD.n1024 VDD.n688 185
R986 VDD.n2758 VDD.n688 185
R987 VDD.n1026 VDD.n1025 185
R988 VDD.n1025 VDD.n687 185
R989 VDD.n1027 VDD.n694 185
R990 VDD.n2752 VDD.n694 185
R991 VDD.n1029 VDD.n1028 185
R992 VDD.n1028 VDD.n693 185
R993 VDD.n1030 VDD.n700 185
R994 VDD.n2746 VDD.n700 185
R995 VDD.n1032 VDD.n1031 185
R996 VDD.n1031 VDD.n699 185
R997 VDD.n1033 VDD.n706 185
R998 VDD.n2740 VDD.n706 185
R999 VDD.n1035 VDD.n1034 185
R1000 VDD.n1034 VDD.n705 185
R1001 VDD.n1036 VDD.n712 185
R1002 VDD.n2734 VDD.n712 185
R1003 VDD.n1038 VDD.n1037 185
R1004 VDD.n1037 VDD.n711 185
R1005 VDD.n1039 VDD.n718 185
R1006 VDD.n2728 VDD.n718 185
R1007 VDD.n1041 VDD.n1040 185
R1008 VDD.n1040 VDD.n717 185
R1009 VDD.n1042 VDD.n723 185
R1010 VDD.n2722 VDD.n723 185
R1011 VDD.n1044 VDD.n1043 185
R1012 VDD.n1043 VDD.n731 185
R1013 VDD.n1045 VDD.n729 185
R1014 VDD.n2716 VDD.n729 185
R1015 VDD.n1047 VDD.n1046 185
R1016 VDD.n1046 VDD.n728 185
R1017 VDD.n1048 VDD.n736 185
R1018 VDD.n2710 VDD.n736 185
R1019 VDD.n1050 VDD.n1049 185
R1020 VDD.n1049 VDD.n735 185
R1021 VDD.n1051 VDD.n742 185
R1022 VDD.n2704 VDD.n742 185
R1023 VDD.n1053 VDD.n1052 185
R1024 VDD.n1052 VDD.n741 185
R1025 VDD.n1054 VDD.n748 185
R1026 VDD.n2698 VDD.n748 185
R1027 VDD.n1056 VDD.n1055 185
R1028 VDD.n1055 VDD.n747 185
R1029 VDD.n1057 VDD.n754 185
R1030 VDD.n2692 VDD.n754 185
R1031 VDD.n1059 VDD.n1058 185
R1032 VDD.n1058 VDD.n753 185
R1033 VDD.n1060 VDD.n760 185
R1034 VDD.n2686 VDD.n760 185
R1035 VDD.n1062 VDD.n1061 185
R1036 VDD.n1061 VDD.n759 185
R1037 VDD.n1063 VDD.n765 185
R1038 VDD.n2680 VDD.n765 185
R1039 VDD.n1065 VDD.n1064 185
R1040 VDD.n1064 VDD.n773 185
R1041 VDD.n1066 VDD.n771 185
R1042 VDD.n2674 VDD.n771 185
R1043 VDD.n1068 VDD.n1067 185
R1044 VDD.n1067 VDD.n770 185
R1045 VDD.n1069 VDD.n777 185
R1046 VDD.n2668 VDD.n777 185
R1047 VDD.n1071 VDD.n1070 185
R1048 VDD.n1070 VDD.n785 185
R1049 VDD.n1072 VDD.n783 185
R1050 VDD.n2662 VDD.n783 185
R1051 VDD.n1074 VDD.n1073 185
R1052 VDD.n1073 VDD.n782 185
R1053 VDD.n1075 VDD.n790 185
R1054 VDD.n2656 VDD.n790 185
R1055 VDD.n1077 VDD.n1076 185
R1056 VDD.n1076 VDD.n789 185
R1057 VDD.n1078 VDD.n796 185
R1058 VDD.n2650 VDD.n796 185
R1059 VDD.n1080 VDD.n1079 185
R1060 VDD.n1079 VDD.n795 185
R1061 VDD.n1081 VDD.n802 185
R1062 VDD.n2644 VDD.n802 185
R1063 VDD.n1083 VDD.n1082 185
R1064 VDD.n1082 VDD.n801 185
R1065 VDD.n1084 VDD.n808 185
R1066 VDD.n2638 VDD.n808 185
R1067 VDD.n1086 VDD.n1085 185
R1068 VDD.n1085 VDD.n807 185
R1069 VDD.n1087 VDD.n814 185
R1070 VDD.n2632 VDD.n814 185
R1071 VDD.n1089 VDD.n1088 185
R1072 VDD.n1088 VDD.n813 185
R1073 VDD.n1090 VDD.n819 185
R1074 VDD.n2626 VDD.n819 185
R1075 VDD.n1092 VDD.n1091 185
R1076 VDD.n1091 VDD.n827 185
R1077 VDD.n1093 VDD.n825 185
R1078 VDD.n2620 VDD.n825 185
R1079 VDD.n1095 VDD.n1094 185
R1080 VDD.n1094 VDD.n824 185
R1081 VDD.n1096 VDD.n832 185
R1082 VDD.n2614 VDD.n832 185
R1083 VDD.n1098 VDD.n1097 185
R1084 VDD.n1097 VDD.n831 185
R1085 VDD.n1099 VDD.n838 185
R1086 VDD.n2608 VDD.n838 185
R1087 VDD.n1101 VDD.n1100 185
R1088 VDD.n1100 VDD.n837 185
R1089 VDD.n1102 VDD.n844 185
R1090 VDD.n2602 VDD.n844 185
R1091 VDD.n1104 VDD.n1103 185
R1092 VDD.n1103 VDD.n843 185
R1093 VDD.n1105 VDD.n850 185
R1094 VDD.n2596 VDD.n850 185
R1095 VDD.n1107 VDD.n1106 185
R1096 VDD.n1106 VDD.n849 185
R1097 VDD.n1108 VDD.n856 185
R1098 VDD.n2590 VDD.n856 185
R1099 VDD.n1110 VDD.n1109 185
R1100 VDD.n1109 VDD.n855 185
R1101 VDD.n1111 VDD.n862 185
R1102 VDD.n2584 VDD.n862 185
R1103 VDD.n1113 VDD.n1112 185
R1104 VDD.n1112 VDD.n861 185
R1105 VDD.n1114 VDD.n868 185
R1106 VDD.n2578 VDD.n868 185
R1107 VDD.n1116 VDD.n1115 185
R1108 VDD.n1115 VDD.n867 185
R1109 VDD.n1117 VDD.n874 185
R1110 VDD.n2572 VDD.n874 185
R1111 VDD.n1119 VDD.n1118 185
R1112 VDD.n1118 VDD.n873 185
R1113 VDD.n1120 VDD.n880 185
R1114 VDD.n2566 VDD.n880 185
R1115 VDD.n1122 VDD.n1121 185
R1116 VDD.n1121 VDD.n879 185
R1117 VDD.n1123 VDD.n886 185
R1118 VDD.n2560 VDD.n886 185
R1119 VDD.n1125 VDD.n1124 185
R1120 VDD.n1124 VDD.n885 185
R1121 VDD.n1126 VDD.n892 185
R1122 VDD.n2554 VDD.n892 185
R1123 VDD.n1128 VDD.n1127 185
R1124 VDD.n1127 VDD.n891 185
R1125 VDD.n1129 VDD.n897 185
R1126 VDD.n2548 VDD.n897 185
R1127 VDD.n1131 VDD.n1130 185
R1128 VDD.n1130 VDD.n905 185
R1129 VDD.n1132 VDD.n903 185
R1130 VDD.n2542 VDD.n903 185
R1131 VDD.n1134 VDD.n1133 185
R1132 VDD.n1133 VDD.n902 185
R1133 VDD.n1135 VDD.n910 185
R1134 VDD.n2536 VDD.n910 185
R1135 VDD.n1137 VDD.n1136 185
R1136 VDD.n1136 VDD.n909 185
R1137 VDD.n1138 VDD.n916 185
R1138 VDD.n2530 VDD.n916 185
R1139 VDD.n1140 VDD.n1139 185
R1140 VDD.n1139 VDD.n915 185
R1141 VDD.n1141 VDD.n922 185
R1142 VDD.n2524 VDD.n922 185
R1143 VDD.n1143 VDD.n1142 185
R1144 VDD.n1142 VDD.n921 185
R1145 VDD.n1144 VDD.n928 185
R1146 VDD.n2518 VDD.n928 185
R1147 VDD.n1146 VDD.n1145 185
R1148 VDD.n1145 VDD.n927 185
R1149 VDD.n1147 VDD.n934 185
R1150 VDD.n2512 VDD.n934 185
R1151 VDD.n1149 VDD.n1148 185
R1152 VDD.n1148 VDD.n933 185
R1153 VDD.n1150 VDD.n940 185
R1154 VDD.n2506 VDD.n940 185
R1155 VDD.n1152 VDD.n1151 185
R1156 VDD.n1151 VDD.n939 185
R1157 VDD.n1153 VDD.n945 185
R1158 VDD.n2500 VDD.n945 185
R1159 VDD.n2417 VDD.n2416 185
R1160 VDD.n2416 VDD.n2415 185
R1161 VDD.n2418 VDD.n951 185
R1162 VDD.n2494 VDD.n951 185
R1163 VDD.n2420 VDD.n2419 185
R1164 VDD.n2419 VDD.n950 185
R1165 VDD.n2421 VDD.n957 185
R1166 VDD.n2488 VDD.n957 185
R1167 VDD.n2423 VDD.n2422 185
R1168 VDD.n2422 VDD.n956 185
R1169 VDD.n2424 VDD.n963 185
R1170 VDD.n2482 VDD.n963 185
R1171 VDD.n2426 VDD.n2425 185
R1172 VDD.n2425 VDD.n962 185
R1173 VDD.n2427 VDD.n969 185
R1174 VDD.n2476 VDD.n969 185
R1175 VDD.n2429 VDD.n2428 185
R1176 VDD.n2428 VDD.n968 185
R1177 VDD.n2430 VDD.n975 185
R1178 VDD.n2470 VDD.n975 185
R1179 VDD.n2432 VDD.n2431 185
R1180 VDD.n2431 VDD.n974 185
R1181 VDD.n3742 VDD.n3741 185
R1182 VDD.n3743 VDD.n3742 185
R1183 VDD.n243 VDD.n241 185
R1184 VDD.n241 VDD.n238 185
R1185 VDD.n3702 VDD.n3701 185
R1186 VDD.n3703 VDD.n3702 185
R1187 VDD.n3700 VDD.n262 185
R1188 VDD.n262 VDD.n259 185
R1189 VDD.n3699 VDD.n3698 185
R1190 VDD.n3698 VDD.n3697 185
R1191 VDD.n264 VDD.n263 185
R1192 VDD.n265 VDD.n264 185
R1193 VDD.n3664 VDD.n3663 185
R1194 VDD.n3665 VDD.n3664 185
R1195 VDD.n3662 VDD.n275 185
R1196 VDD.n275 VDD.n272 185
R1197 VDD.n3661 VDD.n3660 185
R1198 VDD.n3660 VDD.n3659 185
R1199 VDD.n277 VDD.n276 185
R1200 VDD.n278 VDD.n277 185
R1201 VDD.n3652 VDD.n3651 185
R1202 VDD.n3653 VDD.n3652 185
R1203 VDD.n3650 VDD.n286 185
R1204 VDD.n292 VDD.n286 185
R1205 VDD.n3649 VDD.n3648 185
R1206 VDD.n3648 VDD.n3647 185
R1207 VDD.n288 VDD.n287 185
R1208 VDD.n289 VDD.n288 185
R1209 VDD.n3640 VDD.n3639 185
R1210 VDD.n3641 VDD.n3640 185
R1211 VDD.n3638 VDD.n299 185
R1212 VDD.n299 VDD.n296 185
R1213 VDD.n3637 VDD.n3636 185
R1214 VDD.n3636 VDD.n3635 185
R1215 VDD.n301 VDD.n300 185
R1216 VDD.n302 VDD.n301 185
R1217 VDD.n3628 VDD.n3627 185
R1218 VDD.n3629 VDD.n3628 185
R1219 VDD.n3626 VDD.n311 185
R1220 VDD.n311 VDD.n308 185
R1221 VDD.n3625 VDD.n3624 185
R1222 VDD.n3624 VDD.n3623 185
R1223 VDD.n313 VDD.n312 185
R1224 VDD.n314 VDD.n313 185
R1225 VDD.n3616 VDD.n3615 185
R1226 VDD.n3617 VDD.n3616 185
R1227 VDD.n3614 VDD.n323 185
R1228 VDD.n323 VDD.n320 185
R1229 VDD.n3613 VDD.n3612 185
R1230 VDD.n3612 VDD.n3611 185
R1231 VDD.n325 VDD.n324 185
R1232 VDD.n326 VDD.n325 185
R1233 VDD.n3604 VDD.n3603 185
R1234 VDD.n3605 VDD.n3604 185
R1235 VDD.n3602 VDD.n334 185
R1236 VDD.n340 VDD.n334 185
R1237 VDD.n3601 VDD.n3600 185
R1238 VDD.n3600 VDD.n3599 185
R1239 VDD.n336 VDD.n335 185
R1240 VDD.n337 VDD.n336 185
R1241 VDD.n3592 VDD.n3591 185
R1242 VDD.n3593 VDD.n3592 185
R1243 VDD.n3590 VDD.n347 185
R1244 VDD.n347 VDD.n344 185
R1245 VDD.n3589 VDD.n3588 185
R1246 VDD.n3588 VDD.n3587 185
R1247 VDD.n349 VDD.n348 185
R1248 VDD.n350 VDD.n349 185
R1249 VDD.n3580 VDD.n3579 185
R1250 VDD.n3581 VDD.n3580 185
R1251 VDD.n3578 VDD.n359 185
R1252 VDD.n359 VDD.n356 185
R1253 VDD.n3577 VDD.n3576 185
R1254 VDD.n3576 VDD.n3575 185
R1255 VDD.n361 VDD.n360 185
R1256 VDD.n362 VDD.n361 185
R1257 VDD.n3568 VDD.n3567 185
R1258 VDD.n3569 VDD.n3568 185
R1259 VDD.n3566 VDD.n371 185
R1260 VDD.n371 VDD.n368 185
R1261 VDD.n3565 VDD.n3564 185
R1262 VDD.n3564 VDD.n3563 185
R1263 VDD.n373 VDD.n372 185
R1264 VDD.n374 VDD.n373 185
R1265 VDD.n3556 VDD.n3555 185
R1266 VDD.n3557 VDD.n3556 185
R1267 VDD.n3554 VDD.n383 185
R1268 VDD.n383 VDD.n380 185
R1269 VDD.n3553 VDD.n3552 185
R1270 VDD.n3552 VDD.n3551 185
R1271 VDD.n385 VDD.n384 185
R1272 VDD.n386 VDD.n385 185
R1273 VDD.n3544 VDD.n3543 185
R1274 VDD.n3545 VDD.n3544 185
R1275 VDD.n3542 VDD.n395 185
R1276 VDD.n395 VDD.n392 185
R1277 VDD.n3541 VDD.n3540 185
R1278 VDD.n3540 VDD.n3539 185
R1279 VDD.n397 VDD.n396 185
R1280 VDD.n398 VDD.n397 185
R1281 VDD.n3532 VDD.n3531 185
R1282 VDD.n3533 VDD.n3532 185
R1283 VDD.n3530 VDD.n407 185
R1284 VDD.n407 VDD.n404 185
R1285 VDD.n3529 VDD.n3528 185
R1286 VDD.n3528 VDD.n3527 185
R1287 VDD.n409 VDD.n408 185
R1288 VDD.n418 VDD.n409 185
R1289 VDD.n3520 VDD.n3519 185
R1290 VDD.n3521 VDD.n3520 185
R1291 VDD.n3518 VDD.n419 185
R1292 VDD.n419 VDD.n415 185
R1293 VDD.n3517 VDD.n3516 185
R1294 VDD.n3516 VDD.n3515 185
R1295 VDD.n421 VDD.n420 185
R1296 VDD.n422 VDD.n421 185
R1297 VDD.n3508 VDD.n3507 185
R1298 VDD.n3509 VDD.n3508 185
R1299 VDD.n3506 VDD.n431 185
R1300 VDD.n431 VDD.n428 185
R1301 VDD.n3505 VDD.n3504 185
R1302 VDD.n3504 VDD.n3503 185
R1303 VDD.n433 VDD.n432 185
R1304 VDD.n434 VDD.n433 185
R1305 VDD.n3496 VDD.n3495 185
R1306 VDD.n3497 VDD.n3496 185
R1307 VDD.n3494 VDD.n443 185
R1308 VDD.n443 VDD.n440 185
R1309 VDD.n3493 VDD.n3492 185
R1310 VDD.n3492 VDD.n3491 185
R1311 VDD.n445 VDD.n444 185
R1312 VDD.n446 VDD.n445 185
R1313 VDD.n3484 VDD.n3483 185
R1314 VDD.n3485 VDD.n3484 185
R1315 VDD.n3482 VDD.n454 185
R1316 VDD.n460 VDD.n454 185
R1317 VDD.n3481 VDD.n3480 185
R1318 VDD.n3480 VDD.n3479 185
R1319 VDD.n456 VDD.n455 185
R1320 VDD.n457 VDD.n456 185
R1321 VDD.n3472 VDD.n3471 185
R1322 VDD.n3473 VDD.n3472 185
R1323 VDD.n3470 VDD.n466 185
R1324 VDD.n472 VDD.n466 185
R1325 VDD.n3469 VDD.n3468 185
R1326 VDD.n3468 VDD.n3467 185
R1327 VDD.n468 VDD.n467 185
R1328 VDD.n469 VDD.n468 185
R1329 VDD.n3460 VDD.n3459 185
R1330 VDD.n3461 VDD.n3460 185
R1331 VDD.n3458 VDD.n479 185
R1332 VDD.n479 VDD.n476 185
R1333 VDD.n3457 VDD.n3456 185
R1334 VDD.n3456 VDD.n3455 185
R1335 VDD.n481 VDD.n480 185
R1336 VDD.n482 VDD.n481 185
R1337 VDD.n3448 VDD.n3447 185
R1338 VDD.n3449 VDD.n3448 185
R1339 VDD.n3446 VDD.n491 185
R1340 VDD.n491 VDD.n488 185
R1341 VDD.n3445 VDD.n3444 185
R1342 VDD.n3444 VDD.n3443 185
R1343 VDD.n493 VDD.n492 185
R1344 VDD.n494 VDD.n493 185
R1345 VDD.n3436 VDD.n3435 185
R1346 VDD.n3437 VDD.n3436 185
R1347 VDD.n3434 VDD.n503 185
R1348 VDD.n503 VDD.n500 185
R1349 VDD.n3433 VDD.n3432 185
R1350 VDD.n3432 VDD.n3431 185
R1351 VDD.n505 VDD.n504 185
R1352 VDD.n514 VDD.n505 185
R1353 VDD.n3424 VDD.n3423 185
R1354 VDD.n3425 VDD.n3424 185
R1355 VDD.n3422 VDD.n515 185
R1356 VDD.n515 VDD.n511 185
R1357 VDD.n3421 VDD.n3420 185
R1358 VDD.n3420 VDD.n3419 185
R1359 VDD.n517 VDD.n516 185
R1360 VDD.n518 VDD.n517 185
R1361 VDD.n3412 VDD.n3411 185
R1362 VDD.n3413 VDD.n3412 185
R1363 VDD.n3410 VDD.n527 185
R1364 VDD.n527 VDD.n524 185
R1365 VDD.n3409 VDD.n3408 185
R1366 VDD.n3408 VDD.n3407 185
R1367 VDD.n529 VDD.n528 185
R1368 VDD.n530 VDD.n529 185
R1369 VDD.n3400 VDD.n3399 185
R1370 VDD.n3401 VDD.n3400 185
R1371 VDD.n3398 VDD.n539 185
R1372 VDD.n539 VDD.n536 185
R1373 VDD.n3397 VDD.n3396 185
R1374 VDD.n3396 VDD.n3395 185
R1375 VDD.n541 VDD.n540 185
R1376 VDD.n542 VDD.n541 185
R1377 VDD.n3388 VDD.n3387 185
R1378 VDD.n3389 VDD.n3388 185
R1379 VDD.n3386 VDD.n551 185
R1380 VDD.n551 VDD.n548 185
R1381 VDD.n3385 VDD.n3384 185
R1382 VDD.n3384 VDD.n3383 185
R1383 VDD.n553 VDD.n552 185
R1384 VDD.n554 VDD.n553 185
R1385 VDD.n3376 VDD.n3375 185
R1386 VDD.n3377 VDD.n3376 185
R1387 VDD.n3374 VDD.n563 185
R1388 VDD.n563 VDD.n560 185
R1389 VDD.n3373 VDD.n3372 185
R1390 VDD.n3372 VDD.n3371 185
R1391 VDD.n565 VDD.n564 185
R1392 VDD.n566 VDD.n565 185
R1393 VDD.n3364 VDD.n3363 185
R1394 VDD.n3365 VDD.n3364 185
R1395 VDD.n3362 VDD.n575 185
R1396 VDD.n575 VDD.n572 185
R1397 VDD.n3361 VDD.n3360 185
R1398 VDD.n3360 VDD.n3359 185
R1399 VDD.n577 VDD.n576 185
R1400 VDD.n578 VDD.n577 185
R1401 VDD.n3352 VDD.n3351 185
R1402 VDD.n3353 VDD.n3352 185
R1403 VDD.n3350 VDD.n587 185
R1404 VDD.n587 VDD.n584 185
R1405 VDD.n3349 VDD.n3348 185
R1406 VDD.n3348 VDD.n3347 185
R1407 VDD.n589 VDD.n588 185
R1408 VDD.n590 VDD.n589 185
R1409 VDD.n3340 VDD.n3339 185
R1410 VDD.n3341 VDD.n3340 185
R1411 VDD.n3338 VDD.n599 185
R1412 VDD.n599 VDD.n596 185
R1413 VDD.n3337 VDD.n3336 185
R1414 VDD.n3336 VDD.n3335 185
R1415 VDD.n601 VDD.n600 185
R1416 VDD.n2911 VDD.n2909 185
R1417 VDD.n2912 VDD.n2908 185
R1418 VDD.n2912 VDD.n2896 185
R1419 VDD.n2915 VDD.n2914 185
R1420 VDD.n2916 VDD.n2907 185
R1421 VDD.n2918 VDD.n2917 185
R1422 VDD.n2920 VDD.n2906 185
R1423 VDD.n2923 VDD.n2922 185
R1424 VDD.n2924 VDD.n2905 185
R1425 VDD.n2926 VDD.n2925 185
R1426 VDD.n2928 VDD.n2904 185
R1427 VDD.n2931 VDD.n2930 185
R1428 VDD.n2932 VDD.n2903 185
R1429 VDD.n2934 VDD.n2933 185
R1430 VDD.n2936 VDD.n2902 185
R1431 VDD.n2937 VDD.n2899 185
R1432 VDD.n2940 VDD.n2939 185
R1433 VDD.n2941 VDD.n2897 185
R1434 VDD.n2897 VDD.n2896 185
R1435 VDD.n3709 VDD.n3708 185
R1436 VDD.n3711 VDD.n255 185
R1437 VDD.n3713 VDD.n3712 185
R1438 VDD.n3714 VDD.n252 185
R1439 VDD.n3716 VDD.n3715 185
R1440 VDD.n3718 VDD.n250 185
R1441 VDD.n3720 VDD.n3719 185
R1442 VDD.n3721 VDD.n249 185
R1443 VDD.n3723 VDD.n3722 185
R1444 VDD.n3726 VDD.n3725 185
R1445 VDD.n3728 VDD.n3727 185
R1446 VDD.n3730 VDD.n247 185
R1447 VDD.n3732 VDD.n3731 185
R1448 VDD.n3733 VDD.n246 185
R1449 VDD.n3735 VDD.n3734 185
R1450 VDD.n3737 VDD.n244 185
R1451 VDD.n3739 VDD.n3738 185
R1452 VDD.n3740 VDD.n242 185
R1453 VDD.n3707 VDD.n239 185
R1454 VDD.n3743 VDD.n239 185
R1455 VDD.n3706 VDD.n3705 185
R1456 VDD.n3705 VDD.n238 185
R1457 VDD.n3704 VDD.n257 185
R1458 VDD.n3704 VDD.n3703 185
R1459 VDD.n2942 VDD.n258 185
R1460 VDD.n259 VDD.n258 185
R1461 VDD.n2943 VDD.n266 185
R1462 VDD.n3697 VDD.n266 185
R1463 VDD.n2945 VDD.n2944 185
R1464 VDD.n2944 VDD.n265 185
R1465 VDD.n2946 VDD.n273 185
R1466 VDD.n3665 VDD.n273 185
R1467 VDD.n2948 VDD.n2947 185
R1468 VDD.n2947 VDD.n272 185
R1469 VDD.n2949 VDD.n279 185
R1470 VDD.n3659 VDD.n279 185
R1471 VDD.n2951 VDD.n2950 185
R1472 VDD.n2950 VDD.n278 185
R1473 VDD.n2952 VDD.n284 185
R1474 VDD.n3653 VDD.n284 185
R1475 VDD.n2954 VDD.n2953 185
R1476 VDD.n2953 VDD.n292 185
R1477 VDD.n2955 VDD.n290 185
R1478 VDD.n3647 VDD.n290 185
R1479 VDD.n2957 VDD.n2956 185
R1480 VDD.n2956 VDD.n289 185
R1481 VDD.n2958 VDD.n297 185
R1482 VDD.n3641 VDD.n297 185
R1483 VDD.n2960 VDD.n2959 185
R1484 VDD.n2959 VDD.n296 185
R1485 VDD.n2961 VDD.n303 185
R1486 VDD.n3635 VDD.n303 185
R1487 VDD.n2963 VDD.n2962 185
R1488 VDD.n2962 VDD.n302 185
R1489 VDD.n2964 VDD.n309 185
R1490 VDD.n3629 VDD.n309 185
R1491 VDD.n2966 VDD.n2965 185
R1492 VDD.n2965 VDD.n308 185
R1493 VDD.n2967 VDD.n315 185
R1494 VDD.n3623 VDD.n315 185
R1495 VDD.n2969 VDD.n2968 185
R1496 VDD.n2968 VDD.n314 185
R1497 VDD.n2970 VDD.n321 185
R1498 VDD.n3617 VDD.n321 185
R1499 VDD.n2972 VDD.n2971 185
R1500 VDD.n2971 VDD.n320 185
R1501 VDD.n2973 VDD.n327 185
R1502 VDD.n3611 VDD.n327 185
R1503 VDD.n2975 VDD.n2974 185
R1504 VDD.n2974 VDD.n326 185
R1505 VDD.n2976 VDD.n332 185
R1506 VDD.n3605 VDD.n332 185
R1507 VDD.n2978 VDD.n2977 185
R1508 VDD.n2977 VDD.n340 185
R1509 VDD.n2979 VDD.n338 185
R1510 VDD.n3599 VDD.n338 185
R1511 VDD.n2981 VDD.n2980 185
R1512 VDD.n2980 VDD.n337 185
R1513 VDD.n2982 VDD.n345 185
R1514 VDD.n3593 VDD.n345 185
R1515 VDD.n2984 VDD.n2983 185
R1516 VDD.n2983 VDD.n344 185
R1517 VDD.n2985 VDD.n351 185
R1518 VDD.n3587 VDD.n351 185
R1519 VDD.n2987 VDD.n2986 185
R1520 VDD.n2986 VDD.n350 185
R1521 VDD.n2988 VDD.n357 185
R1522 VDD.n3581 VDD.n357 185
R1523 VDD.n2990 VDD.n2989 185
R1524 VDD.n2989 VDD.n356 185
R1525 VDD.n2991 VDD.n363 185
R1526 VDD.n3575 VDD.n363 185
R1527 VDD.n2993 VDD.n2992 185
R1528 VDD.n2992 VDD.n362 185
R1529 VDD.n2994 VDD.n369 185
R1530 VDD.n3569 VDD.n369 185
R1531 VDD.n2996 VDD.n2995 185
R1532 VDD.n2995 VDD.n368 185
R1533 VDD.n2997 VDD.n375 185
R1534 VDD.n3563 VDD.n375 185
R1535 VDD.n2999 VDD.n2998 185
R1536 VDD.n2998 VDD.n374 185
R1537 VDD.n3000 VDD.n381 185
R1538 VDD.n3557 VDD.n381 185
R1539 VDD.n3002 VDD.n3001 185
R1540 VDD.n3001 VDD.n380 185
R1541 VDD.n3003 VDD.n387 185
R1542 VDD.n3551 VDD.n387 185
R1543 VDD.n3005 VDD.n3004 185
R1544 VDD.n3004 VDD.n386 185
R1545 VDD.n3006 VDD.n393 185
R1546 VDD.n3545 VDD.n393 185
R1547 VDD.n3008 VDD.n3007 185
R1548 VDD.n3007 VDD.n392 185
R1549 VDD.n3009 VDD.n399 185
R1550 VDD.n3539 VDD.n399 185
R1551 VDD.n3011 VDD.n3010 185
R1552 VDD.n3010 VDD.n398 185
R1553 VDD.n3012 VDD.n405 185
R1554 VDD.n3533 VDD.n405 185
R1555 VDD.n3014 VDD.n3013 185
R1556 VDD.n3013 VDD.n404 185
R1557 VDD.n3015 VDD.n410 185
R1558 VDD.n3527 VDD.n410 185
R1559 VDD.n3017 VDD.n3016 185
R1560 VDD.n3016 VDD.n418 185
R1561 VDD.n3018 VDD.n416 185
R1562 VDD.n3521 VDD.n416 185
R1563 VDD.n3020 VDD.n3019 185
R1564 VDD.n3019 VDD.n415 185
R1565 VDD.n3021 VDD.n423 185
R1566 VDD.n3515 VDD.n423 185
R1567 VDD.n3023 VDD.n3022 185
R1568 VDD.n3022 VDD.n422 185
R1569 VDD.n3024 VDD.n429 185
R1570 VDD.n3509 VDD.n429 185
R1571 VDD.n3026 VDD.n3025 185
R1572 VDD.n3025 VDD.n428 185
R1573 VDD.n3027 VDD.n435 185
R1574 VDD.n3503 VDD.n435 185
R1575 VDD.n3029 VDD.n3028 185
R1576 VDD.n3028 VDD.n434 185
R1577 VDD.n3030 VDD.n441 185
R1578 VDD.n3497 VDD.n441 185
R1579 VDD.n3032 VDD.n3031 185
R1580 VDD.n3031 VDD.n440 185
R1581 VDD.n3033 VDD.n447 185
R1582 VDD.n3491 VDD.n447 185
R1583 VDD.n3035 VDD.n3034 185
R1584 VDD.n3034 VDD.n446 185
R1585 VDD.n3036 VDD.n452 185
R1586 VDD.n3485 VDD.n452 185
R1587 VDD.n3038 VDD.n3037 185
R1588 VDD.n3037 VDD.n460 185
R1589 VDD.n3039 VDD.n458 185
R1590 VDD.n3479 VDD.n458 185
R1591 VDD.n3041 VDD.n3040 185
R1592 VDD.n3040 VDD.n457 185
R1593 VDD.n3042 VDD.n464 185
R1594 VDD.n3473 VDD.n464 185
R1595 VDD.n3044 VDD.n3043 185
R1596 VDD.n3043 VDD.n472 185
R1597 VDD.n3045 VDD.n470 185
R1598 VDD.n3467 VDD.n470 185
R1599 VDD.n3047 VDD.n3046 185
R1600 VDD.n3046 VDD.n469 185
R1601 VDD.n3048 VDD.n477 185
R1602 VDD.n3461 VDD.n477 185
R1603 VDD.n3050 VDD.n3049 185
R1604 VDD.n3049 VDD.n476 185
R1605 VDD.n3051 VDD.n483 185
R1606 VDD.n3455 VDD.n483 185
R1607 VDD.n3053 VDD.n3052 185
R1608 VDD.n3052 VDD.n482 185
R1609 VDD.n3054 VDD.n489 185
R1610 VDD.n3449 VDD.n489 185
R1611 VDD.n3056 VDD.n3055 185
R1612 VDD.n3055 VDD.n488 185
R1613 VDD.n3057 VDD.n495 185
R1614 VDD.n3443 VDD.n495 185
R1615 VDD.n3059 VDD.n3058 185
R1616 VDD.n3058 VDD.n494 185
R1617 VDD.n3060 VDD.n501 185
R1618 VDD.n3437 VDD.n501 185
R1619 VDD.n3062 VDD.n3061 185
R1620 VDD.n3061 VDD.n500 185
R1621 VDD.n3063 VDD.n506 185
R1622 VDD.n3431 VDD.n506 185
R1623 VDD.n3065 VDD.n3064 185
R1624 VDD.n3064 VDD.n514 185
R1625 VDD.n3066 VDD.n512 185
R1626 VDD.n3425 VDD.n512 185
R1627 VDD.n3068 VDD.n3067 185
R1628 VDD.n3067 VDD.n511 185
R1629 VDD.n3069 VDD.n519 185
R1630 VDD.n3419 VDD.n519 185
R1631 VDD.n3071 VDD.n3070 185
R1632 VDD.n3070 VDD.n518 185
R1633 VDD.n3072 VDD.n525 185
R1634 VDD.n3413 VDD.n525 185
R1635 VDD.n3074 VDD.n3073 185
R1636 VDD.n3073 VDD.n524 185
R1637 VDD.n3075 VDD.n531 185
R1638 VDD.n3407 VDD.n531 185
R1639 VDD.n3077 VDD.n3076 185
R1640 VDD.n3076 VDD.n530 185
R1641 VDD.n3078 VDD.n537 185
R1642 VDD.n3401 VDD.n537 185
R1643 VDD.n3080 VDD.n3079 185
R1644 VDD.n3079 VDD.n536 185
R1645 VDD.n3081 VDD.n543 185
R1646 VDD.n3395 VDD.n543 185
R1647 VDD.n3083 VDD.n3082 185
R1648 VDD.n3082 VDD.n542 185
R1649 VDD.n3084 VDD.n549 185
R1650 VDD.n3389 VDD.n549 185
R1651 VDD.n3086 VDD.n3085 185
R1652 VDD.n3085 VDD.n548 185
R1653 VDD.n3087 VDD.n555 185
R1654 VDD.n3383 VDD.n555 185
R1655 VDD.n3089 VDD.n3088 185
R1656 VDD.n3088 VDD.n554 185
R1657 VDD.n3090 VDD.n561 185
R1658 VDD.n3377 VDD.n561 185
R1659 VDD.n3092 VDD.n3091 185
R1660 VDD.n3091 VDD.n560 185
R1661 VDD.n3093 VDD.n567 185
R1662 VDD.n3371 VDD.n567 185
R1663 VDD.n3095 VDD.n3094 185
R1664 VDD.n3094 VDD.n566 185
R1665 VDD.n3096 VDD.n573 185
R1666 VDD.n3365 VDD.n573 185
R1667 VDD.n3098 VDD.n3097 185
R1668 VDD.n3097 VDD.n572 185
R1669 VDD.n3099 VDD.n579 185
R1670 VDD.n3359 VDD.n579 185
R1671 VDD.n3101 VDD.n3100 185
R1672 VDD.n3100 VDD.n578 185
R1673 VDD.n3102 VDD.n585 185
R1674 VDD.n3353 VDD.n585 185
R1675 VDD.n3104 VDD.n3103 185
R1676 VDD.n3103 VDD.n584 185
R1677 VDD.n3105 VDD.n591 185
R1678 VDD.n3347 VDD.n591 185
R1679 VDD.n3107 VDD.n3106 185
R1680 VDD.n3106 VDD.n590 185
R1681 VDD.n3108 VDD.n597 185
R1682 VDD.n3341 VDD.n597 185
R1683 VDD.n3109 VDD.n2898 185
R1684 VDD.n2898 VDD.n596 185
R1685 VDD.n3111 VDD.n3110 185
R1686 VDD.n3335 VDD.n3111 185
R1687 VDD.n2169 VDD.n2168 185
R1688 VDD.n2170 VDD.n2169 185
R1689 VDD.n1212 VDD.n1210 185
R1690 VDD.n1210 VDD.n1209 185
R1691 VDD.n1947 VDD.n1946 185
R1692 VDD.n1946 VDD.n1945 185
R1693 VDD.n1215 VDD.n1214 185
R1694 VDD.n1216 VDD.n1215 185
R1695 VDD.n1934 VDD.n1933 185
R1696 VDD.n1935 VDD.n1934 185
R1697 VDD.n1225 VDD.n1224 185
R1698 VDD.n1224 VDD.n1223 185
R1699 VDD.n1929 VDD.n1928 185
R1700 VDD.n1928 VDD.n1927 185
R1701 VDD.n1228 VDD.n1227 185
R1702 VDD.n1229 VDD.n1228 185
R1703 VDD.n1918 VDD.n1917 185
R1704 VDD.n1919 VDD.n1918 185
R1705 VDD.n1237 VDD.n1236 185
R1706 VDD.n1236 VDD.n1235 185
R1707 VDD.n1913 VDD.n1912 185
R1708 VDD.n1912 VDD.n1911 185
R1709 VDD.n1240 VDD.n1239 185
R1710 VDD.n1241 VDD.n1240 185
R1711 VDD.n1902 VDD.n1901 185
R1712 VDD.n1903 VDD.n1902 185
R1713 VDD.n1249 VDD.n1248 185
R1714 VDD.n1248 VDD.n1247 185
R1715 VDD.n1897 VDD.n1896 185
R1716 VDD.n1896 VDD.n1895 185
R1717 VDD.n1252 VDD.n1251 185
R1718 VDD.n1253 VDD.n1252 185
R1719 VDD.n1886 VDD.n1885 185
R1720 VDD.n1887 VDD.n1886 185
R1721 VDD.n1261 VDD.n1260 185
R1722 VDD.n1260 VDD.n1259 185
R1723 VDD.n1881 VDD.n1880 185
R1724 VDD.n1880 VDD.n1879 185
R1725 VDD.n1264 VDD.n1263 185
R1726 VDD.n1265 VDD.n1264 185
R1727 VDD.n1870 VDD.n1869 185
R1728 VDD.n1871 VDD.n1870 185
R1729 VDD.n1273 VDD.n1272 185
R1730 VDD.n1272 VDD.n1271 185
R1731 VDD.n1865 VDD.n1864 185
R1732 VDD.n1864 VDD.n1863 185
R1733 VDD.n1276 VDD.n1275 185
R1734 VDD.n1277 VDD.n1276 185
R1735 VDD.n1854 VDD.n1853 185
R1736 VDD.n1855 VDD.n1854 185
R1737 VDD.n1285 VDD.n1284 185
R1738 VDD.n1284 VDD.n1283 185
R1739 VDD.n1849 VDD.n1848 185
R1740 VDD.n1848 VDD.n1847 185
R1741 VDD.n1288 VDD.n1287 185
R1742 VDD.n1289 VDD.n1288 185
R1743 VDD.n1838 VDD.n1837 185
R1744 VDD.n1839 VDD.n1838 185
R1745 VDD.n1297 VDD.n1296 185
R1746 VDD.n1296 VDD.n1295 185
R1747 VDD.n1818 VDD.n1817 185
R1748 VDD.n1817 VDD.t0 185
R1749 VDD.n1300 VDD.n1299 185
R1750 VDD.n1301 VDD.n1300 185
R1751 VDD.n1808 VDD.n1807 185
R1752 VDD.n1809 VDD.n1808 185
R1753 VDD.n1309 VDD.n1308 185
R1754 VDD.n1308 VDD.n1307 185
R1755 VDD.n1803 VDD.n1802 185
R1756 VDD.n1802 VDD.n1801 185
R1757 VDD.n1312 VDD.n1311 185
R1758 VDD.n1313 VDD.n1312 185
R1759 VDD.n1792 VDD.n1791 185
R1760 VDD.n1793 VDD.n1792 185
R1761 VDD.n1321 VDD.n1320 185
R1762 VDD.n1320 VDD.n1319 185
R1763 VDD.n1787 VDD.n1786 185
R1764 VDD.n1786 VDD.n1785 185
R1765 VDD.n1324 VDD.n1323 185
R1766 VDD.n1325 VDD.n1324 185
R1767 VDD.n1776 VDD.n1775 185
R1768 VDD.n1777 VDD.n1776 185
R1769 VDD.n1332 VDD.n1331 185
R1770 VDD.n1768 VDD.n1331 185
R1771 VDD.n1771 VDD.n1770 185
R1772 VDD.n1770 VDD.n1769 185
R1773 VDD.n1335 VDD.n1334 185
R1774 VDD.n1336 VDD.n1335 185
R1775 VDD.n1759 VDD.n1758 185
R1776 VDD.n1760 VDD.n1759 185
R1777 VDD.n1344 VDD.n1343 185
R1778 VDD.n1343 VDD.n1342 185
R1779 VDD.n1754 VDD.n1753 185
R1780 VDD.n1753 VDD.n1752 185
R1781 VDD.n1347 VDD.n1346 185
R1782 VDD.n1348 VDD.n1347 185
R1783 VDD.n1743 VDD.n1742 185
R1784 VDD.n1744 VDD.n1743 185
R1785 VDD.n1356 VDD.n1355 185
R1786 VDD.n1355 VDD.n1354 185
R1787 VDD.n1738 VDD.n1737 185
R1788 VDD.n1737 VDD.n1736 185
R1789 VDD.n1359 VDD.n1358 185
R1790 VDD.n1360 VDD.n1359 185
R1791 VDD.n1727 VDD.n1726 185
R1792 VDD.n1728 VDD.n1727 185
R1793 VDD.n1368 VDD.n1367 185
R1794 VDD.n1367 VDD.n1366 185
R1795 VDD.n1722 VDD.n1721 185
R1796 VDD.n1721 VDD.n1720 185
R1797 VDD.n1371 VDD.n1370 185
R1798 VDD.n1378 VDD.n1371 185
R1799 VDD.n1711 VDD.n1710 185
R1800 VDD.n1712 VDD.n1711 185
R1801 VDD.n1380 VDD.n1379 185
R1802 VDD.n1379 VDD.n1377 185
R1803 VDD.n1706 VDD.n1705 185
R1804 VDD.n1705 VDD.n1704 185
R1805 VDD.n1383 VDD.n1382 185
R1806 VDD.n1384 VDD.n1383 185
R1807 VDD.n1695 VDD.n1694 185
R1808 VDD.n1696 VDD.n1695 185
R1809 VDD.n1691 VDD.n1390 185
R1810 VDD.n1690 VDD.n1393 185
R1811 VDD.n1689 VDD.n1394 185
R1812 VDD.n1394 VDD.n1389 185
R1813 VDD.n1397 VDD.n1395 185
R1814 VDD.n1685 VDD.n1399 185
R1815 VDD.n1684 VDD.n1400 185
R1816 VDD.n1683 VDD.n1402 185
R1817 VDD.n1405 VDD.n1403 185
R1818 VDD.n1679 VDD.n1407 185
R1819 VDD.n1678 VDD.n1408 185
R1820 VDD.n1677 VDD.n1410 185
R1821 VDD.n1413 VDD.n1411 185
R1822 VDD.n1673 VDD.n1415 185
R1823 VDD.n1672 VDD.n1416 185
R1824 VDD.n1671 VDD.n1418 185
R1825 VDD.n1668 VDD.n1423 185
R1826 VDD.n1667 VDD.n1425 185
R1827 VDD.n1666 VDD.n1426 185
R1828 VDD.n1430 VDD.n1427 185
R1829 VDD.n1662 VDD.n1431 185
R1830 VDD.n1661 VDD.n1433 185
R1831 VDD.n1660 VDD.n1434 185
R1832 VDD.n1438 VDD.n1435 185
R1833 VDD.n1656 VDD.n1439 185
R1834 VDD.n1655 VDD.n1441 185
R1835 VDD.n1654 VDD.n1442 185
R1836 VDD.n1446 VDD.n1443 185
R1837 VDD.n1650 VDD.n1447 185
R1838 VDD.n1649 VDD.n1449 185
R1839 VDD.n1648 VDD.n1450 185
R1840 VDD.n1454 VDD.n1451 185
R1841 VDD.n1644 VDD.n1455 185
R1842 VDD.n1640 VDD.n1457 185
R1843 VDD.n1639 VDD.n1458 185
R1844 VDD.n1462 VDD.n1459 185
R1845 VDD.n1635 VDD.n1463 185
R1846 VDD.n1634 VDD.n1465 185
R1847 VDD.n1633 VDD.n1466 185
R1848 VDD.n1470 VDD.n1467 185
R1849 VDD.n1629 VDD.n1471 185
R1850 VDD.n1628 VDD.n1473 185
R1851 VDD.n1627 VDD.n1474 185
R1852 VDD.n1478 VDD.n1475 185
R1853 VDD.n1623 VDD.n1479 185
R1854 VDD.n1622 VDD.n1481 185
R1855 VDD.n1621 VDD.n1482 185
R1856 VDD.n1486 VDD.n1483 185
R1857 VDD.n1617 VDD.n1487 185
R1858 VDD.n1616 VDD.n1489 185
R1859 VDD.n1615 VDD.n1614 185
R1860 VDD.n1612 VDD.n1493 185
R1861 VDD.n1611 VDD.n1610 185
R1862 VDD.n1498 VDD.n1495 185
R1863 VDD.n1606 VDD.n1499 185
R1864 VDD.n1605 VDD.n1501 185
R1865 VDD.n1604 VDD.n1502 185
R1866 VDD.n1506 VDD.n1503 185
R1867 VDD.n1600 VDD.n1507 185
R1868 VDD.n1599 VDD.n1509 185
R1869 VDD.n1598 VDD.n1510 185
R1870 VDD.n1514 VDD.n1511 185
R1871 VDD.n1594 VDD.n1515 185
R1872 VDD.n1593 VDD.n1517 185
R1873 VDD.n1592 VDD.n1518 185
R1874 VDD.n1523 VDD.n1519 185
R1875 VDD.n1588 VDD.n1585 185
R1876 VDD.n1583 VDD.n1521 185
R1877 VDD.n1582 VDD.n1581 185
R1878 VDD.n1527 VDD.n1525 185
R1879 VDD.n1577 VDD.n1528 185
R1880 VDD.n1576 VDD.n1530 185
R1881 VDD.n1575 VDD.n1531 185
R1882 VDD.n1535 VDD.n1532 185
R1883 VDD.n1571 VDD.n1536 185
R1884 VDD.n1570 VDD.n1538 185
R1885 VDD.n1569 VDD.n1539 185
R1886 VDD.n1543 VDD.n1540 185
R1887 VDD.n1565 VDD.n1544 185
R1888 VDD.n1564 VDD.n1546 185
R1889 VDD.n1563 VDD.n1547 185
R1890 VDD.n1551 VDD.n1548 185
R1891 VDD.n1559 VDD.n1552 185
R1892 VDD.n1558 VDD.n1555 185
R1893 VDD.n1553 VDD.n1388 185
R1894 VDD.n1389 VDD.n1388 185
R1895 VDD.n2172 VDD.n1188 185
R1896 VDD.n2175 VDD.n2174 185
R1897 VDD.n1191 VDD.n1186 185
R1898 VDD.n2179 VDD.n1185 185
R1899 VDD.n2180 VDD.n1184 185
R1900 VDD.n2181 VDD.n1183 185
R1901 VDD.n1202 VDD.n1181 185
R1902 VDD.n2185 VDD.n1180 185
R1903 VDD.n2186 VDD.n1179 185
R1904 VDD.n2187 VDD.n1178 185
R1905 VDD.n1199 VDD.n1176 185
R1906 VDD.n2191 VDD.n1175 185
R1907 VDD.n2192 VDD.n1174 185
R1908 VDD.n2193 VDD.n1173 185
R1909 VDD.n1196 VDD.n1171 185
R1910 VDD.n2197 VDD.n1170 185
R1911 VDD.n2198 VDD.n1169 185
R1912 VDD.n2199 VDD.n1168 185
R1913 VDD.n1193 VDD.n1166 185
R1914 VDD.n2203 VDD.n1163 185
R1915 VDD.n2204 VDD.n1162 185
R1916 VDD.n2205 VDD.n1161 185
R1917 VDD.n2052 VDD.n1160 185
R1918 VDD.n2055 VDD.n2054 185
R1919 VDD.n2057 VDD.n2056 185
R1920 VDD.n2060 VDD.n2059 185
R1921 VDD.n2062 VDD.n2061 185
R1922 VDD.n2064 VDD.n2050 185
R1923 VDD.n2066 VDD.n2065 185
R1924 VDD.n2067 VDD.n2045 185
R1925 VDD.n2069 VDD.n2068 185
R1926 VDD.n2071 VDD.n2043 185
R1927 VDD.n2073 VDD.n2072 185
R1928 VDD.n2040 VDD.n2039 185
R1929 VDD.n2078 VDD.n2077 185
R1930 VDD.n2080 VDD.n2037 185
R1931 VDD.n2082 VDD.n2081 185
R1932 VDD.n2083 VDD.n2030 185
R1933 VDD.n2085 VDD.n2084 185
R1934 VDD.n2087 VDD.n2028 185
R1935 VDD.n2089 VDD.n2088 185
R1936 VDD.n2090 VDD.n2023 185
R1937 VDD.n2092 VDD.n2091 185
R1938 VDD.n2094 VDD.n2021 185
R1939 VDD.n2096 VDD.n2095 185
R1940 VDD.n2097 VDD.n2016 185
R1941 VDD.n2099 VDD.n2098 185
R1942 VDD.n2101 VDD.n2014 185
R1943 VDD.n2103 VDD.n2102 185
R1944 VDD.n2104 VDD.n2009 185
R1945 VDD.n2106 VDD.n2105 185
R1946 VDD.n2108 VDD.n2008 185
R1947 VDD.n2110 VDD.n2109 185
R1948 VDD.n2111 VDD.n1999 185
R1949 VDD.n2113 VDD.n2112 185
R1950 VDD.n2115 VDD.n1998 185
R1951 VDD.n2116 VDD.n1995 185
R1952 VDD.n2119 VDD.n2118 185
R1953 VDD.n1997 VDD.n1993 185
R1954 VDD.n2123 VDD.n1991 185
R1955 VDD.n2125 VDD.n2124 185
R1956 VDD.n2127 VDD.n1989 185
R1957 VDD.n2129 VDD.n2128 185
R1958 VDD.n2130 VDD.n1984 185
R1959 VDD.n2132 VDD.n2131 185
R1960 VDD.n2134 VDD.n1982 185
R1961 VDD.n2136 VDD.n2135 185
R1962 VDD.n2137 VDD.n1974 185
R1963 VDD.n2139 VDD.n2138 185
R1964 VDD.n2141 VDD.n1972 185
R1965 VDD.n2143 VDD.n2142 185
R1966 VDD.n2144 VDD.n1967 185
R1967 VDD.n2146 VDD.n2145 185
R1968 VDD.n2148 VDD.n1965 185
R1969 VDD.n2150 VDD.n2149 185
R1970 VDD.n2151 VDD.n1960 185
R1971 VDD.n2153 VDD.n2152 185
R1972 VDD.n2155 VDD.n1958 185
R1973 VDD.n2157 VDD.n2156 185
R1974 VDD.n2158 VDD.n1953 185
R1975 VDD.n2160 VDD.n2159 185
R1976 VDD.n2162 VDD.n1951 185
R1977 VDD.n2164 VDD.n2163 185
R1978 VDD.n2165 VDD.n1211 185
R1979 VDD.n2171 VDD.n1208 185
R1980 VDD.n2171 VDD.n2170 185
R1981 VDD.n1219 VDD.n1207 185
R1982 VDD.n1209 VDD.n1207 185
R1983 VDD.n1944 VDD.n1943 185
R1984 VDD.n1945 VDD.n1944 185
R1985 VDD.n1218 VDD.n1217 185
R1986 VDD.n1217 VDD.n1216 185
R1987 VDD.n1937 VDD.n1936 185
R1988 VDD.n1936 VDD.n1935 185
R1989 VDD.n1222 VDD.n1221 185
R1990 VDD.n1223 VDD.n1222 185
R1991 VDD.n1926 VDD.n1925 185
R1992 VDD.n1927 VDD.n1926 185
R1993 VDD.n1231 VDD.n1230 185
R1994 VDD.n1230 VDD.n1229 185
R1995 VDD.n1921 VDD.n1920 185
R1996 VDD.n1920 VDD.n1919 185
R1997 VDD.n1234 VDD.n1233 185
R1998 VDD.n1235 VDD.n1234 185
R1999 VDD.n1910 VDD.n1909 185
R2000 VDD.n1911 VDD.n1910 185
R2001 VDD.n1243 VDD.n1242 185
R2002 VDD.n1242 VDD.n1241 185
R2003 VDD.n1905 VDD.n1904 185
R2004 VDD.n1904 VDD.n1903 185
R2005 VDD.n1246 VDD.n1245 185
R2006 VDD.n1247 VDD.n1246 185
R2007 VDD.n1894 VDD.n1893 185
R2008 VDD.n1895 VDD.n1894 185
R2009 VDD.n1255 VDD.n1254 185
R2010 VDD.n1254 VDD.n1253 185
R2011 VDD.n1889 VDD.n1888 185
R2012 VDD.n1888 VDD.n1887 185
R2013 VDD.n1258 VDD.n1257 185
R2014 VDD.n1259 VDD.n1258 185
R2015 VDD.n1878 VDD.n1877 185
R2016 VDD.n1879 VDD.n1878 185
R2017 VDD.n1267 VDD.n1266 185
R2018 VDD.n1266 VDD.n1265 185
R2019 VDD.n1873 VDD.n1872 185
R2020 VDD.n1872 VDD.n1871 185
R2021 VDD.n1270 VDD.n1269 185
R2022 VDD.n1271 VDD.n1270 185
R2023 VDD.n1862 VDD.n1861 185
R2024 VDD.n1863 VDD.n1862 185
R2025 VDD.n1279 VDD.n1278 185
R2026 VDD.n1278 VDD.n1277 185
R2027 VDD.n1857 VDD.n1856 185
R2028 VDD.n1856 VDD.n1855 185
R2029 VDD.n1282 VDD.n1281 185
R2030 VDD.n1283 VDD.n1282 185
R2031 VDD.n1846 VDD.n1845 185
R2032 VDD.n1847 VDD.n1846 185
R2033 VDD.n1291 VDD.n1290 185
R2034 VDD.n1290 VDD.n1289 185
R2035 VDD.n1841 VDD.n1840 185
R2036 VDD.n1840 VDD.n1839 185
R2037 VDD.n1294 VDD.n1293 185
R2038 VDD.n1295 VDD.n1294 185
R2039 VDD.n1816 VDD.n1815 185
R2040 VDD.t0 VDD.n1816 185
R2041 VDD.n1303 VDD.n1302 185
R2042 VDD.n1302 VDD.n1301 185
R2043 VDD.n1811 VDD.n1810 185
R2044 VDD.n1810 VDD.n1809 185
R2045 VDD.n1306 VDD.n1305 185
R2046 VDD.n1307 VDD.n1306 185
R2047 VDD.n1800 VDD.n1799 185
R2048 VDD.n1801 VDD.n1800 185
R2049 VDD.n1315 VDD.n1314 185
R2050 VDD.n1314 VDD.n1313 185
R2051 VDD.n1795 VDD.n1794 185
R2052 VDD.n1794 VDD.n1793 185
R2053 VDD.n1318 VDD.n1317 185
R2054 VDD.n1319 VDD.n1318 185
R2055 VDD.n1784 VDD.n1783 185
R2056 VDD.n1785 VDD.n1784 185
R2057 VDD.n1327 VDD.n1326 185
R2058 VDD.n1326 VDD.n1325 185
R2059 VDD.n1779 VDD.n1778 185
R2060 VDD.n1778 VDD.n1777 185
R2061 VDD.n1330 VDD.n1329 185
R2062 VDD.n1768 VDD.n1330 185
R2063 VDD.n1767 VDD.n1766 185
R2064 VDD.n1769 VDD.n1767 185
R2065 VDD.n1338 VDD.n1337 185
R2066 VDD.n1337 VDD.n1336 185
R2067 VDD.n1762 VDD.n1761 185
R2068 VDD.n1761 VDD.n1760 185
R2069 VDD.n1341 VDD.n1340 185
R2070 VDD.n1342 VDD.n1341 185
R2071 VDD.n1751 VDD.n1750 185
R2072 VDD.n1752 VDD.n1751 185
R2073 VDD.n1350 VDD.n1349 185
R2074 VDD.n1349 VDD.n1348 185
R2075 VDD.n1746 VDD.n1745 185
R2076 VDD.n1745 VDD.n1744 185
R2077 VDD.n1353 VDD.n1352 185
R2078 VDD.n1354 VDD.n1353 185
R2079 VDD.n1735 VDD.n1734 185
R2080 VDD.n1736 VDD.n1735 185
R2081 VDD.n1362 VDD.n1361 185
R2082 VDD.n1361 VDD.n1360 185
R2083 VDD.n1730 VDD.n1729 185
R2084 VDD.n1729 VDD.n1728 185
R2085 VDD.n1365 VDD.n1364 185
R2086 VDD.n1366 VDD.n1365 185
R2087 VDD.n1719 VDD.n1718 185
R2088 VDD.n1720 VDD.n1719 185
R2089 VDD.n1373 VDD.n1372 185
R2090 VDD.n1378 VDD.n1372 185
R2091 VDD.n1714 VDD.n1713 185
R2092 VDD.n1713 VDD.n1712 185
R2093 VDD.n1376 VDD.n1375 185
R2094 VDD.n1377 VDD.n1376 185
R2095 VDD.n1703 VDD.n1702 185
R2096 VDD.n1704 VDD.n1703 185
R2097 VDD.n1386 VDD.n1385 185
R2098 VDD.n1385 VDD.n1384 185
R2099 VDD.n1698 VDD.n1697 185
R2100 VDD.n1697 VDD.n1696 185
R2101 VDD.n3964 VDD.n127 185
R2102 VDD.n3963 VDD.n3962 185
R2103 VDD.n3960 VDD.n129 185
R2104 VDD.n3960 VDD.n126 185
R2105 VDD.n3959 VDD.n3958 185
R2106 VDD.n3957 VDD.n3956 185
R2107 VDD.n3955 VDD.n134 185
R2108 VDD.n3953 VDD.n3952 185
R2109 VDD.n3951 VDD.n135 185
R2110 VDD.n3950 VDD.n3949 185
R2111 VDD.n3947 VDD.n140 185
R2112 VDD.n3945 VDD.n3944 185
R2113 VDD.n3943 VDD.n141 185
R2114 VDD.n3942 VDD.n3941 185
R2115 VDD.n3939 VDD.n146 185
R2116 VDD.n3937 VDD.n3936 185
R2117 VDD.n3934 VDD.n147 185
R2118 VDD.n3933 VDD.n3932 185
R2119 VDD.n3930 VDD.n154 185
R2120 VDD.n3928 VDD.n3927 185
R2121 VDD.n3926 VDD.n155 185
R2122 VDD.n3925 VDD.n3924 185
R2123 VDD.n3922 VDD.n160 185
R2124 VDD.n3920 VDD.n3919 185
R2125 VDD.n162 VDD.n161 185
R2126 VDD.n167 VDD.n165 185
R2127 VDD.n3914 VDD.n168 185
R2128 VDD.n3913 VDD.n3912 185
R2129 VDD.n3910 VDD.n169 185
R2130 VDD.n3908 VDD.n3907 185
R2131 VDD.n3906 VDD.n170 185
R2132 VDD.n3905 VDD.n3904 185
R2133 VDD.n3902 VDD.n175 185
R2134 VDD.n3900 VDD.n3899 185
R2135 VDD.n3898 VDD.n176 185
R2136 VDD.n3897 VDD.n3896 185
R2137 VDD.n3894 VDD.n184 185
R2138 VDD.n3892 VDD.n3891 185
R2139 VDD.n3890 VDD.n185 185
R2140 VDD.n3889 VDD.n3888 185
R2141 VDD.n3886 VDD.n190 185
R2142 VDD.n3884 VDD.n3883 185
R2143 VDD.n3882 VDD.n191 185
R2144 VDD.n3881 VDD.n3880 185
R2145 VDD.n3878 VDD.n196 185
R2146 VDD.n3876 VDD.n3875 185
R2147 VDD.n3874 VDD.n197 185
R2148 VDD.n3873 VDD.n3872 185
R2149 VDD.n3870 VDD.n202 185
R2150 VDD.n3868 VDD.n3867 185
R2151 VDD.n3866 VDD.n203 185
R2152 VDD.n3865 VDD.n3864 185
R2153 VDD.n3862 VDD.n210 185
R2154 VDD.n3860 VDD.n3859 185
R2155 VDD.n3858 VDD.n211 185
R2156 VDD.n3857 VDD.n3856 185
R2157 VDD.n3854 VDD.n216 185
R2158 VDD.n3852 VDD.n3851 185
R2159 VDD.n3850 VDD.n217 185
R2160 VDD.n3849 VDD.n3848 185
R2161 VDD.n3846 VDD.n3845 185
R2162 VDD.n3844 VDD.n3843 185
R2163 VDD.n3842 VDD.n3841 185
R2164 VDD.n3840 VDD.n3839 185
R2165 VDD.n3838 VDD.n3764 185
R2166 VDD.n3836 VDD.n3835 185
R2167 VDD.n3834 VDD.n3765 185
R2168 VDD.n3772 VDD.n3768 185
R2169 VDD.n3828 VDD.n3827 185
R2170 VDD.n3825 VDD.n3770 185
R2171 VDD.n3824 VDD.n3823 185
R2172 VDD.n3822 VDD.n3821 185
R2173 VDD.n3820 VDD.n3776 185
R2174 VDD.n3818 VDD.n3817 185
R2175 VDD.n3816 VDD.n3777 185
R2176 VDD.n3815 VDD.n3814 185
R2177 VDD.n3812 VDD.n3782 185
R2178 VDD.n3810 VDD.n3809 185
R2179 VDD.n3808 VDD.n3783 185
R2180 VDD.n3807 VDD.n3806 185
R2181 VDD.n3804 VDD.n3788 185
R2182 VDD.n3802 VDD.n3801 185
R2183 VDD.n3800 VDD.n3789 185
R2184 VDD.n3797 VDD.n3794 185
R2185 VDD.n3792 VDD.n125 185
R2186 VDD.n126 VDD.n125 185
R2187 VDD.n4319 VDD.n4318 185
R2188 VDD.n4385 VDD.n4314 185
R2189 VDD.n4387 VDD.n4386 185
R2190 VDD.n4389 VDD.n4312 185
R2191 VDD.n4391 VDD.n4390 185
R2192 VDD.n4392 VDD.n4307 185
R2193 VDD.n4394 VDD.n4393 185
R2194 VDD.n4396 VDD.n4305 185
R2195 VDD.n4398 VDD.n4397 185
R2196 VDD.n4399 VDD.n4300 185
R2197 VDD.n4401 VDD.n4400 185
R2198 VDD.n4403 VDD.n4298 185
R2199 VDD.n4405 VDD.n4404 185
R2200 VDD.n4406 VDD.n4294 185
R2201 VDD.n4408 VDD.n4407 185
R2202 VDD.n4410 VDD.n4292 185
R2203 VDD.n4412 VDD.n4411 185
R2204 VDD.n4287 VDD.n4286 185
R2205 VDD.n4417 VDD.n4416 185
R2206 VDD.n4419 VDD.n4284 185
R2207 VDD.n4421 VDD.n4420 185
R2208 VDD.n4422 VDD.n4279 185
R2209 VDD.n4424 VDD.n4423 185
R2210 VDD.n4426 VDD.n4277 185
R2211 VDD.n4428 VDD.n4427 185
R2212 VDD.n4429 VDD.n4272 185
R2213 VDD.n4431 VDD.n4430 185
R2214 VDD.n4433 VDD.n4270 185
R2215 VDD.n4435 VDD.n4434 185
R2216 VDD.n4436 VDD.n4266 185
R2217 VDD.n4438 VDD.n4437 185
R2218 VDD.n4440 VDD.n4264 185
R2219 VDD.n4442 VDD.n4441 185
R2220 VDD.n4261 VDD.n4260 185
R2221 VDD.n4447 VDD.n4446 185
R2222 VDD.n4449 VDD.n4258 185
R2223 VDD.n4451 VDD.n4450 185
R2224 VDD.n4452 VDD.n4251 185
R2225 VDD.n4454 VDD.n4453 185
R2226 VDD.n4456 VDD.n4249 185
R2227 VDD.n4458 VDD.n4457 185
R2228 VDD.n4459 VDD.n4244 185
R2229 VDD.n4461 VDD.n4460 185
R2230 VDD.n4463 VDD.n4242 185
R2231 VDD.n4465 VDD.n4464 185
R2232 VDD.n4466 VDD.n4237 185
R2233 VDD.n4468 VDD.n4467 185
R2234 VDD.n4470 VDD.n4235 185
R2235 VDD.n4472 VDD.n4471 185
R2236 VDD.n4473 VDD.n4230 185
R2237 VDD.n4475 VDD.n4474 185
R2238 VDD.n4477 VDD.n4229 185
R2239 VDD.n4479 VDD.n4478 185
R2240 VDD.n4480 VDD.n4220 185
R2241 VDD.n4482 VDD.n4481 185
R2242 VDD.n4484 VDD.n4218 185
R2243 VDD.n4486 VDD.n4485 185
R2244 VDD.n4487 VDD.n4213 185
R2245 VDD.n4489 VDD.n4488 185
R2246 VDD.n4491 VDD.n4211 185
R2247 VDD.n4493 VDD.n4492 185
R2248 VDD.n4494 VDD.n4206 185
R2249 VDD.n4496 VDD.n4495 185
R2250 VDD.n4498 VDD.n4204 185
R2251 VDD.n4500 VDD.n4499 185
R2252 VDD.n4501 VDD.n4199 185
R2253 VDD.n4503 VDD.n4502 185
R2254 VDD.n4505 VDD.n4197 185
R2255 VDD.n4507 VDD.n4506 185
R2256 VDD.n4511 VDD.n4192 185
R2257 VDD.n4513 VDD.n4512 185
R2258 VDD.n4515 VDD.n4190 185
R2259 VDD.n4517 VDD.n4516 185
R2260 VDD.n4518 VDD.n4185 185
R2261 VDD.n4520 VDD.n4519 185
R2262 VDD.n4522 VDD.n4183 185
R2263 VDD.n4524 VDD.n4523 185
R2264 VDD.n4525 VDD.n4177 185
R2265 VDD.n4527 VDD.n4526 185
R2266 VDD.n4529 VDD.n4176 185
R2267 VDD.n4530 VDD.n4175 185
R2268 VDD.n4533 VDD.n4532 185
R2269 VDD.n4534 VDD.n4173 185
R2270 VDD.n4535 VDD.n4169 185
R2271 VDD.n4381 VDD.n4167 185
R2272 VDD.n4540 VDD.n4167 185
R2273 VDD.n4380 VDD.n4166 185
R2274 VDD.n4541 VDD.n4166 185
R2275 VDD.n4379 VDD.n4165 185
R2276 VDD.n4542 VDD.n4165 185
R2277 VDD.n4324 VDD.n4323 185
R2278 VDD.n4323 VDD.n4157 185
R2279 VDD.n4375 VDD.n4156 185
R2280 VDD.n4548 VDD.n4156 185
R2281 VDD.n4374 VDD.n4155 185
R2282 VDD.n4549 VDD.n4155 185
R2283 VDD.n4373 VDD.n4154 185
R2284 VDD.n4550 VDD.n4154 185
R2285 VDD.n4327 VDD.n4326 185
R2286 VDD.n4326 VDD.n4146 185
R2287 VDD.n4369 VDD.n4145 185
R2288 VDD.n4556 VDD.n4145 185
R2289 VDD.n4368 VDD.n4144 185
R2290 VDD.n4557 VDD.n4144 185
R2291 VDD.n4367 VDD.n4143 185
R2292 VDD.n4558 VDD.n4143 185
R2293 VDD.n4330 VDD.n4329 185
R2294 VDD.n4329 VDD.n4135 185
R2295 VDD.n4363 VDD.n4134 185
R2296 VDD.n4564 VDD.n4134 185
R2297 VDD.n4362 VDD.n4133 185
R2298 VDD.n4565 VDD.n4133 185
R2299 VDD.n4361 VDD.n4132 185
R2300 VDD.n4566 VDD.n4132 185
R2301 VDD.n4333 VDD.n4332 185
R2302 VDD.n4332 VDD.n4124 185
R2303 VDD.n4357 VDD.n4123 185
R2304 VDD.n4572 VDD.n4123 185
R2305 VDD.n4356 VDD.n4122 185
R2306 VDD.n4573 VDD.n4122 185
R2307 VDD.n4355 VDD.n4121 185
R2308 VDD.n4574 VDD.n4121 185
R2309 VDD.n4336 VDD.n4335 185
R2310 VDD.n4335 VDD.n4120 185
R2311 VDD.n4351 VDD.n4112 185
R2312 VDD.n4580 VDD.n4112 185
R2313 VDD.n4350 VDD.n4111 185
R2314 VDD.n4581 VDD.n4111 185
R2315 VDD.n4349 VDD.n4110 185
R2316 VDD.n4582 VDD.n4110 185
R2317 VDD.n4339 VDD.n4338 185
R2318 VDD.n4338 VDD.n4102 185
R2319 VDD.n4345 VDD.n4101 185
R2320 VDD.n4588 VDD.n4101 185
R2321 VDD.n4344 VDD.n4100 185
R2322 VDD.n4589 VDD.n4100 185
R2323 VDD.n4343 VDD.n4099 185
R2324 VDD.n4590 VDD.n4099 185
R2325 VDD.n4091 VDD.n4090 185
R2326 VDD.n4092 VDD.n4091 185
R2327 VDD.n4598 VDD.n4597 185
R2328 VDD.n4597 VDD.n4596 185
R2329 VDD.n4599 VDD.n39 185
R2330 VDD.n39 VDD.n37 185
R2331 VDD.n4601 VDD.n4600 185
R2332 VDD.t6 VDD.n4601 185
R2333 VDD.n40 VDD.n38 185
R2334 VDD.n38 VDD.n36 185
R2335 VDD.n4084 VDD.n4083 185
R2336 VDD.n4083 VDD.n4082 185
R2337 VDD.n43 VDD.n42 185
R2338 VDD.n44 VDD.n43 185
R2339 VDD.n4073 VDD.n4072 185
R2340 VDD.n4074 VDD.n4073 185
R2341 VDD.n52 VDD.n51 185
R2342 VDD.n51 VDD.n50 185
R2343 VDD.n4068 VDD.n4067 185
R2344 VDD.n4067 VDD.n4066 185
R2345 VDD.n55 VDD.n54 185
R2346 VDD.n56 VDD.n55 185
R2347 VDD.n4057 VDD.n4056 185
R2348 VDD.n4058 VDD.n4057 185
R2349 VDD.n64 VDD.n63 185
R2350 VDD.n63 VDD.n62 185
R2351 VDD.n4052 VDD.n4051 185
R2352 VDD.n4051 VDD.n4050 185
R2353 VDD.n67 VDD.n66 185
R2354 VDD.n4041 VDD.n67 185
R2355 VDD.n4040 VDD.n4039 185
R2356 VDD.n4042 VDD.n4040 185
R2357 VDD.n75 VDD.n74 185
R2358 VDD.n74 VDD.n73 185
R2359 VDD.n4035 VDD.n4034 185
R2360 VDD.n4034 VDD.n4033 185
R2361 VDD.n78 VDD.n77 185
R2362 VDD.n79 VDD.n78 185
R2363 VDD.n4024 VDD.n4023 185
R2364 VDD.n4025 VDD.n4024 185
R2365 VDD.n87 VDD.n86 185
R2366 VDD.n86 VDD.n85 185
R2367 VDD.n4019 VDD.n4018 185
R2368 VDD.n4018 VDD.n4017 185
R2369 VDD.n90 VDD.n89 185
R2370 VDD.n91 VDD.n90 185
R2371 VDD.n4008 VDD.n4007 185
R2372 VDD.n4009 VDD.n4008 185
R2373 VDD.n99 VDD.n98 185
R2374 VDD.n98 VDD.n97 185
R2375 VDD.n4003 VDD.n4002 185
R2376 VDD.n4002 VDD.n4001 185
R2377 VDD.n102 VDD.n101 185
R2378 VDD.n103 VDD.n102 185
R2379 VDD.n3992 VDD.n3991 185
R2380 VDD.n3993 VDD.n3992 185
R2381 VDD.n110 VDD.n109 185
R2382 VDD.n115 VDD.n109 185
R2383 VDD.n3987 VDD.n3986 185
R2384 VDD.n3986 VDD.n3985 185
R2385 VDD.n113 VDD.n112 185
R2386 VDD.n114 VDD.n113 185
R2387 VDD.n3976 VDD.n3975 185
R2388 VDD.n3977 VDD.n3976 185
R2389 VDD.n123 VDD.n122 185
R2390 VDD.n122 VDD.n121 185
R2391 VDD.n3971 VDD.n3970 185
R2392 VDD.n3970 VDD.n3969 185
R2393 VDD.n3968 VDD.n3967 185
R2394 VDD.n3969 VDD.n3968 185
R2395 VDD.n120 VDD.n119 185
R2396 VDD.n121 VDD.n120 185
R2397 VDD.n3979 VDD.n3978 185
R2398 VDD.n3978 VDD.n3977 185
R2399 VDD.n117 VDD.n116 185
R2400 VDD.n116 VDD.n114 185
R2401 VDD.n3984 VDD.n3983 185
R2402 VDD.n3985 VDD.n3984 185
R2403 VDD.n108 VDD.n107 185
R2404 VDD.n115 VDD.n108 185
R2405 VDD.n3995 VDD.n3994 185
R2406 VDD.n3994 VDD.n3993 185
R2407 VDD.n105 VDD.n104 185
R2408 VDD.n104 VDD.n103 185
R2409 VDD.n4000 VDD.n3999 185
R2410 VDD.n4001 VDD.n4000 185
R2411 VDD.n96 VDD.n95 185
R2412 VDD.n97 VDD.n96 185
R2413 VDD.n4011 VDD.n4010 185
R2414 VDD.n4010 VDD.n4009 185
R2415 VDD.n93 VDD.n92 185
R2416 VDD.n92 VDD.n91 185
R2417 VDD.n4016 VDD.n4015 185
R2418 VDD.n4017 VDD.n4016 185
R2419 VDD.n84 VDD.n83 185
R2420 VDD.n85 VDD.n84 185
R2421 VDD.n4027 VDD.n4026 185
R2422 VDD.n4026 VDD.n4025 185
R2423 VDD.n81 VDD.n80 185
R2424 VDD.n80 VDD.n79 185
R2425 VDD.n4032 VDD.n4031 185
R2426 VDD.n4033 VDD.n4032 185
R2427 VDD.n72 VDD.n71 185
R2428 VDD.n73 VDD.n72 185
R2429 VDD.n4044 VDD.n4043 185
R2430 VDD.n4043 VDD.n4042 185
R2431 VDD.n69 VDD.n68 185
R2432 VDD.n4041 VDD.n68 185
R2433 VDD.n4049 VDD.n4048 185
R2434 VDD.n4050 VDD.n4049 185
R2435 VDD.n61 VDD.n60 185
R2436 VDD.n62 VDD.n61 185
R2437 VDD.n4060 VDD.n4059 185
R2438 VDD.n4059 VDD.n4058 185
R2439 VDD.n58 VDD.n57 185
R2440 VDD.n57 VDD.n56 185
R2441 VDD.n4065 VDD.n4064 185
R2442 VDD.n4066 VDD.n4065 185
R2443 VDD.n49 VDD.n48 185
R2444 VDD.n50 VDD.n49 185
R2445 VDD.n4076 VDD.n4075 185
R2446 VDD.n4075 VDD.n4074 185
R2447 VDD.n46 VDD.n45 185
R2448 VDD.n45 VDD.n44 185
R2449 VDD.n4081 VDD.n4080 185
R2450 VDD.n4082 VDD.n4081 185
R2451 VDD.n34 VDD.n32 185
R2452 VDD.n36 VDD.n34 185
R2453 VDD.n4603 VDD.n4602 185
R2454 VDD.n4602 VDD.t6 185
R2455 VDD.n35 VDD.n33 185
R2456 VDD.n37 VDD.n35 185
R2457 VDD.n4595 VDD.n4594 185
R2458 VDD.n4596 VDD.n4595 185
R2459 VDD.n4593 VDD.n4093 185
R2460 VDD.n4093 VDD.n4092 185
R2461 VDD.n4592 VDD.n4591 185
R2462 VDD.n4591 VDD.n4590 185
R2463 VDD.n4098 VDD.n4097 185
R2464 VDD.n4589 VDD.n4098 185
R2465 VDD.n4587 VDD.n4586 185
R2466 VDD.n4588 VDD.n4587 185
R2467 VDD.n4585 VDD.n4103 185
R2468 VDD.n4103 VDD.n4102 185
R2469 VDD.n4584 VDD.n4583 185
R2470 VDD.n4583 VDD.n4582 185
R2471 VDD.n4109 VDD.n4108 185
R2472 VDD.n4581 VDD.n4109 185
R2473 VDD.n4579 VDD.n4578 185
R2474 VDD.n4580 VDD.n4579 185
R2475 VDD.n4577 VDD.n4113 185
R2476 VDD.n4120 VDD.n4113 185
R2477 VDD.n4576 VDD.n4575 185
R2478 VDD.n4575 VDD.n4574 185
R2479 VDD.n4119 VDD.n4118 185
R2480 VDD.n4573 VDD.n4119 185
R2481 VDD.n4571 VDD.n4570 185
R2482 VDD.n4572 VDD.n4571 185
R2483 VDD.n4569 VDD.n4125 185
R2484 VDD.n4125 VDD.n4124 185
R2485 VDD.n4568 VDD.n4567 185
R2486 VDD.n4567 VDD.n4566 185
R2487 VDD.n4131 VDD.n4130 185
R2488 VDD.n4565 VDD.n4131 185
R2489 VDD.n4563 VDD.n4562 185
R2490 VDD.n4564 VDD.n4563 185
R2491 VDD.n4561 VDD.n4136 185
R2492 VDD.n4136 VDD.n4135 185
R2493 VDD.n4560 VDD.n4559 185
R2494 VDD.n4559 VDD.n4558 185
R2495 VDD.n4142 VDD.n4141 185
R2496 VDD.n4557 VDD.n4142 185
R2497 VDD.n4555 VDD.n4554 185
R2498 VDD.n4556 VDD.n4555 185
R2499 VDD.n4553 VDD.n4147 185
R2500 VDD.n4147 VDD.n4146 185
R2501 VDD.n4552 VDD.n4551 185
R2502 VDD.n4551 VDD.n4550 185
R2503 VDD.n4153 VDD.n4152 185
R2504 VDD.n4549 VDD.n4153 185
R2505 VDD.n4547 VDD.n4546 185
R2506 VDD.n4548 VDD.n4547 185
R2507 VDD.n4545 VDD.n4158 185
R2508 VDD.n4158 VDD.n4157 185
R2509 VDD.n4544 VDD.n4543 185
R2510 VDD.n4543 VDD.n4542 185
R2511 VDD.n4164 VDD.n4163 185
R2512 VDD.n4541 VDD.n4164 185
R2513 VDD.n4539 VDD.n4538 185
R2514 VDD.n4540 VDD.n4539 185
R2515 VDD.n623 VDD.n621 185
R2516 VDD.n621 VDD.n602 185
R2517 VDD.n2798 VDD.n630 185
R2518 VDD.n2857 VDD.n630 185
R2519 VDD.n2800 VDD.n2799 185
R2520 VDD.n2799 VDD.n628 185
R2521 VDD.n2801 VDD.n640 185
R2522 VDD.n2811 VDD.n640 185
R2523 VDD.n2802 VDD.n648 185
R2524 VDD.n648 VDD.n638 185
R2525 VDD.n2804 VDD.n2803 185
R2526 VDD.n2805 VDD.n2804 185
R2527 VDD.n2797 VDD.n647 185
R2528 VDD.n647 VDD.n644 185
R2529 VDD.n2796 VDD.n2795 185
R2530 VDD.n2795 VDD.n2794 185
R2531 VDD.n650 VDD.n649 185
R2532 VDD.n651 VDD.n650 185
R2533 VDD.n2787 VDD.n2786 185
R2534 VDD.n2788 VDD.n2787 185
R2535 VDD.n2785 VDD.n660 185
R2536 VDD.n660 VDD.n657 185
R2537 VDD.n2784 VDD.n2783 185
R2538 VDD.n2783 VDD.n2782 185
R2539 VDD.n662 VDD.n661 185
R2540 VDD.n663 VDD.n662 185
R2541 VDD.n2775 VDD.n2774 185
R2542 VDD.n2776 VDD.n2775 185
R2543 VDD.n2773 VDD.n672 185
R2544 VDD.n672 VDD.n669 185
R2545 VDD.n2772 VDD.n2771 185
R2546 VDD.n2771 VDD.n2770 185
R2547 VDD.n674 VDD.n673 185
R2548 VDD.n675 VDD.n674 185
R2549 VDD.n2763 VDD.n2762 185
R2550 VDD.n2764 VDD.n2763 185
R2551 VDD.n2761 VDD.n684 185
R2552 VDD.n684 VDD.n681 185
R2553 VDD.n2760 VDD.n2759 185
R2554 VDD.n2759 VDD.n2758 185
R2555 VDD.n686 VDD.n685 185
R2556 VDD.n687 VDD.n686 185
R2557 VDD.n2751 VDD.n2750 185
R2558 VDD.n2752 VDD.n2751 185
R2559 VDD.n2749 VDD.n696 185
R2560 VDD.n696 VDD.n693 185
R2561 VDD.n2748 VDD.n2747 185
R2562 VDD.n2747 VDD.n2746 185
R2563 VDD.n698 VDD.n697 185
R2564 VDD.n699 VDD.n698 185
R2565 VDD.n2739 VDD.n2738 185
R2566 VDD.n2740 VDD.n2739 185
R2567 VDD.n2737 VDD.n708 185
R2568 VDD.n708 VDD.n705 185
R2569 VDD.n2736 VDD.n2735 185
R2570 VDD.n2735 VDD.n2734 185
R2571 VDD.n710 VDD.n709 185
R2572 VDD.n711 VDD.n710 185
R2573 VDD.n2727 VDD.n2726 185
R2574 VDD.n2728 VDD.n2727 185
R2575 VDD.n2725 VDD.n720 185
R2576 VDD.n720 VDD.n717 185
R2577 VDD.n2724 VDD.n2723 185
R2578 VDD.n2723 VDD.n2722 185
R2579 VDD.n722 VDD.n721 185
R2580 VDD.n731 VDD.n722 185
R2581 VDD.n2715 VDD.n2714 185
R2582 VDD.n2716 VDD.n2715 185
R2583 VDD.n2713 VDD.n732 185
R2584 VDD.n732 VDD.n728 185
R2585 VDD.n2712 VDD.n2711 185
R2586 VDD.n2711 VDD.n2710 185
R2587 VDD.n734 VDD.n733 185
R2588 VDD.n735 VDD.n734 185
R2589 VDD.n2703 VDD.n2702 185
R2590 VDD.n2704 VDD.n2703 185
R2591 VDD.n2701 VDD.n744 185
R2592 VDD.n744 VDD.n741 185
R2593 VDD.n2700 VDD.n2699 185
R2594 VDD.n2699 VDD.n2698 185
R2595 VDD.n746 VDD.n745 185
R2596 VDD.n747 VDD.n746 185
R2597 VDD.n2691 VDD.n2690 185
R2598 VDD.n2692 VDD.n2691 185
R2599 VDD.n2689 VDD.n756 185
R2600 VDD.n756 VDD.n753 185
R2601 VDD.n2688 VDD.n2687 185
R2602 VDD.n2687 VDD.n2686 185
R2603 VDD.n758 VDD.n757 185
R2604 VDD.n759 VDD.n758 185
R2605 VDD.n2679 VDD.n2678 185
R2606 VDD.n2680 VDD.n2679 185
R2607 VDD.n2677 VDD.n767 185
R2608 VDD.n773 VDD.n767 185
R2609 VDD.n2676 VDD.n2675 185
R2610 VDD.n2675 VDD.n2674 185
R2611 VDD.n769 VDD.n768 185
R2612 VDD.n770 VDD.n769 185
R2613 VDD.n2667 VDD.n2666 185
R2614 VDD.n2668 VDD.n2667 185
R2615 VDD.n2665 VDD.n779 185
R2616 VDD.n785 VDD.n779 185
R2617 VDD.n2664 VDD.n2663 185
R2618 VDD.n2663 VDD.n2662 185
R2619 VDD.n781 VDD.n780 185
R2620 VDD.n782 VDD.n781 185
R2621 VDD.n2655 VDD.n2654 185
R2622 VDD.n2656 VDD.n2655 185
R2623 VDD.n2653 VDD.n792 185
R2624 VDD.n792 VDD.n789 185
R2625 VDD.n2652 VDD.n2651 185
R2626 VDD.n2651 VDD.n2650 185
R2627 VDD.n794 VDD.n793 185
R2628 VDD.n795 VDD.n794 185
R2629 VDD.n2643 VDD.n2642 185
R2630 VDD.n2644 VDD.n2643 185
R2631 VDD.n2641 VDD.n804 185
R2632 VDD.n804 VDD.n801 185
R2633 VDD.n2640 VDD.n2639 185
R2634 VDD.n2639 VDD.n2638 185
R2635 VDD.n806 VDD.n805 185
R2636 VDD.n807 VDD.n806 185
R2637 VDD.n2631 VDD.n2630 185
R2638 VDD.n2632 VDD.n2631 185
R2639 VDD.n2629 VDD.n816 185
R2640 VDD.n816 VDD.n813 185
R2641 VDD.n2628 VDD.n2627 185
R2642 VDD.n2627 VDD.n2626 185
R2643 VDD.n818 VDD.n817 185
R2644 VDD.n827 VDD.n818 185
R2645 VDD.n2619 VDD.n2618 185
R2646 VDD.n2620 VDD.n2619 185
R2647 VDD.n2617 VDD.n828 185
R2648 VDD.n828 VDD.n824 185
R2649 VDD.n2616 VDD.n2615 185
R2650 VDD.n2615 VDD.n2614 185
R2651 VDD.n830 VDD.n829 185
R2652 VDD.n831 VDD.n830 185
R2653 VDD.n2607 VDD.n2606 185
R2654 VDD.n2608 VDD.n2607 185
R2655 VDD.n2605 VDD.n840 185
R2656 VDD.n840 VDD.n837 185
R2657 VDD.n2604 VDD.n2603 185
R2658 VDD.n2603 VDD.n2602 185
R2659 VDD.n842 VDD.n841 185
R2660 VDD.n843 VDD.n842 185
R2661 VDD.n2595 VDD.n2594 185
R2662 VDD.n2596 VDD.n2595 185
R2663 VDD.n2593 VDD.n852 185
R2664 VDD.n852 VDD.n849 185
R2665 VDD.n2592 VDD.n2591 185
R2666 VDD.n2591 VDD.n2590 185
R2667 VDD.n854 VDD.n853 185
R2668 VDD.n855 VDD.n854 185
R2669 VDD.n2583 VDD.n2582 185
R2670 VDD.n2584 VDD.n2583 185
R2671 VDD.n2581 VDD.n864 185
R2672 VDD.n864 VDD.n861 185
R2673 VDD.n2580 VDD.n2579 185
R2674 VDD.n2579 VDD.n2578 185
R2675 VDD.n866 VDD.n865 185
R2676 VDD.n867 VDD.n866 185
R2677 VDD.n2571 VDD.n2570 185
R2678 VDD.n2572 VDD.n2571 185
R2679 VDD.n2569 VDD.n876 185
R2680 VDD.n876 VDD.n873 185
R2681 VDD.n2568 VDD.n2567 185
R2682 VDD.n2567 VDD.n2566 185
R2683 VDD.n878 VDD.n877 185
R2684 VDD.n879 VDD.n878 185
R2685 VDD.n2559 VDD.n2558 185
R2686 VDD.n2560 VDD.n2559 185
R2687 VDD.n2557 VDD.n888 185
R2688 VDD.n888 VDD.n885 185
R2689 VDD.n2556 VDD.n2555 185
R2690 VDD.n2555 VDD.n2554 185
R2691 VDD.n890 VDD.n889 185
R2692 VDD.n891 VDD.n890 185
R2693 VDD.n2547 VDD.n2546 185
R2694 VDD.n2548 VDD.n2547 185
R2695 VDD.n2545 VDD.n899 185
R2696 VDD.n905 VDD.n899 185
R2697 VDD.n2544 VDD.n2543 185
R2698 VDD.n2543 VDD.n2542 185
R2699 VDD.n901 VDD.n900 185
R2700 VDD.n902 VDD.n901 185
R2701 VDD.n2535 VDD.n2534 185
R2702 VDD.n2536 VDD.n2535 185
R2703 VDD.n2533 VDD.n912 185
R2704 VDD.n912 VDD.n909 185
R2705 VDD.n2532 VDD.n2531 185
R2706 VDD.n2531 VDD.n2530 185
R2707 VDD.n914 VDD.n913 185
R2708 VDD.n915 VDD.n914 185
R2709 VDD.n2523 VDD.n2522 185
R2710 VDD.n2524 VDD.n2523 185
R2711 VDD.n2521 VDD.n924 185
R2712 VDD.n924 VDD.n921 185
R2713 VDD.n2520 VDD.n2519 185
R2714 VDD.n2519 VDD.n2518 185
R2715 VDD.n926 VDD.n925 185
R2716 VDD.n927 VDD.n926 185
R2717 VDD.n2511 VDD.n2510 185
R2718 VDD.n2512 VDD.n2511 185
R2719 VDD.n2509 VDD.n936 185
R2720 VDD.n936 VDD.n933 185
R2721 VDD.n2508 VDD.n2507 185
R2722 VDD.n2507 VDD.n2506 185
R2723 VDD.n938 VDD.n937 185
R2724 VDD.n939 VDD.n938 185
R2725 VDD.n2499 VDD.n2498 185
R2726 VDD.n2500 VDD.n2499 185
R2727 VDD.n2497 VDD.n947 185
R2728 VDD.n2415 VDD.n947 185
R2729 VDD.n2496 VDD.n2495 185
R2730 VDD.n2495 VDD.n2494 185
R2731 VDD.n949 VDD.n948 185
R2732 VDD.n950 VDD.n949 185
R2733 VDD.n2487 VDD.n2486 185
R2734 VDD.n2488 VDD.n2487 185
R2735 VDD.n2485 VDD.n959 185
R2736 VDD.n959 VDD.n956 185
R2737 VDD.n2484 VDD.n2483 185
R2738 VDD.n2483 VDD.n2482 185
R2739 VDD.n961 VDD.n960 185
R2740 VDD.n962 VDD.n961 185
R2741 VDD.n2475 VDD.n2474 185
R2742 VDD.n2476 VDD.n2475 185
R2743 VDD.n2473 VDD.n971 185
R2744 VDD.n971 VDD.n968 185
R2745 VDD.n2472 VDD.n2471 185
R2746 VDD.n2471 VDD.n2470 185
R2747 VDD.n973 VDD.n972 185
R2748 VDD.n974 VDD.n973 185
R2749 VDD.n2861 VDD.n620 185
R2750 VDD.n2895 VDD.n620 185
R2751 VDD.n2863 VDD.n2862 185
R2752 VDD.n2865 VDD.n2864 185
R2753 VDD.n2867 VDD.n2866 185
R2754 VDD.n2869 VDD.n2868 185
R2755 VDD.n2871 VDD.n2870 185
R2756 VDD.n2873 VDD.n2872 185
R2757 VDD.n2875 VDD.n2874 185
R2758 VDD.n2877 VDD.n2876 185
R2759 VDD.n2879 VDD.n2878 185
R2760 VDD.n2881 VDD.n2880 185
R2761 VDD.n2883 VDD.n2882 185
R2762 VDD.n2885 VDD.n2884 185
R2763 VDD.n2887 VDD.n2886 185
R2764 VDD.n2889 VDD.n2888 185
R2765 VDD.n2891 VDD.n2890 185
R2766 VDD.n2892 VDD.n622 185
R2767 VDD.n2894 VDD.n2893 185
R2768 VDD.n2895 VDD.n2894 185
R2769 VDD.n2860 VDD.n2859 185
R2770 VDD.n2859 VDD.n602 185
R2771 VDD.n2858 VDD.n626 185
R2772 VDD.n2858 VDD.n2857 185
R2773 VDD.n2258 VDD.n627 185
R2774 VDD.n628 VDD.n627 185
R2775 VDD.n2259 VDD.n639 185
R2776 VDD.n2811 VDD.n639 185
R2777 VDD.n2261 VDD.n2260 185
R2778 VDD.n2260 VDD.n638 185
R2779 VDD.n2262 VDD.n646 185
R2780 VDD.n2805 VDD.n646 185
R2781 VDD.n2264 VDD.n2263 185
R2782 VDD.n2263 VDD.n644 185
R2783 VDD.n2265 VDD.n653 185
R2784 VDD.n2794 VDD.n653 185
R2785 VDD.n2267 VDD.n2266 185
R2786 VDD.n2266 VDD.n651 185
R2787 VDD.n2268 VDD.n659 185
R2788 VDD.n2788 VDD.n659 185
R2789 VDD.n2270 VDD.n2269 185
R2790 VDD.n2269 VDD.n657 185
R2791 VDD.n2271 VDD.n665 185
R2792 VDD.n2782 VDD.n665 185
R2793 VDD.n2273 VDD.n2272 185
R2794 VDD.n2272 VDD.n663 185
R2795 VDD.n2274 VDD.n671 185
R2796 VDD.n2776 VDD.n671 185
R2797 VDD.n2276 VDD.n2275 185
R2798 VDD.n2275 VDD.n669 185
R2799 VDD.n2277 VDD.n677 185
R2800 VDD.n2770 VDD.n677 185
R2801 VDD.n2279 VDD.n2278 185
R2802 VDD.n2278 VDD.n675 185
R2803 VDD.n2280 VDD.n683 185
R2804 VDD.n2764 VDD.n683 185
R2805 VDD.n2282 VDD.n2281 185
R2806 VDD.n2281 VDD.n681 185
R2807 VDD.n2283 VDD.n689 185
R2808 VDD.n2758 VDD.n689 185
R2809 VDD.n2285 VDD.n2284 185
R2810 VDD.n2284 VDD.n687 185
R2811 VDD.n2286 VDD.n695 185
R2812 VDD.n2752 VDD.n695 185
R2813 VDD.n2288 VDD.n2287 185
R2814 VDD.n2287 VDD.n693 185
R2815 VDD.n2289 VDD.n701 185
R2816 VDD.n2746 VDD.n701 185
R2817 VDD.n2291 VDD.n2290 185
R2818 VDD.n2290 VDD.n699 185
R2819 VDD.n2292 VDD.n707 185
R2820 VDD.n2740 VDD.n707 185
R2821 VDD.n2294 VDD.n2293 185
R2822 VDD.n2293 VDD.n705 185
R2823 VDD.n2295 VDD.n713 185
R2824 VDD.n2734 VDD.n713 185
R2825 VDD.n2297 VDD.n2296 185
R2826 VDD.n2296 VDD.n711 185
R2827 VDD.n2298 VDD.n719 185
R2828 VDD.n2728 VDD.n719 185
R2829 VDD.n2300 VDD.n2299 185
R2830 VDD.n2299 VDD.n717 185
R2831 VDD.n2301 VDD.n724 185
R2832 VDD.n2722 VDD.n724 185
R2833 VDD.n2303 VDD.n2302 185
R2834 VDD.n2302 VDD.n731 185
R2835 VDD.n2304 VDD.n730 185
R2836 VDD.n2716 VDD.n730 185
R2837 VDD.n2306 VDD.n2305 185
R2838 VDD.n2305 VDD.n728 185
R2839 VDD.n2307 VDD.n737 185
R2840 VDD.n2710 VDD.n737 185
R2841 VDD.n2309 VDD.n2308 185
R2842 VDD.n2308 VDD.n735 185
R2843 VDD.n2310 VDD.n743 185
R2844 VDD.n2704 VDD.n743 185
R2845 VDD.n2312 VDD.n2311 185
R2846 VDD.n2311 VDD.n741 185
R2847 VDD.n2313 VDD.n749 185
R2848 VDD.n2698 VDD.n749 185
R2849 VDD.n2315 VDD.n2314 185
R2850 VDD.n2314 VDD.n747 185
R2851 VDD.n2316 VDD.n755 185
R2852 VDD.n2692 VDD.n755 185
R2853 VDD.n2318 VDD.n2317 185
R2854 VDD.n2317 VDD.n753 185
R2855 VDD.n2319 VDD.n761 185
R2856 VDD.n2686 VDD.n761 185
R2857 VDD.n2321 VDD.n2320 185
R2858 VDD.n2320 VDD.n759 185
R2859 VDD.n2322 VDD.n766 185
R2860 VDD.n2680 VDD.n766 185
R2861 VDD.n2324 VDD.n2323 185
R2862 VDD.n2323 VDD.n773 185
R2863 VDD.n2325 VDD.n772 185
R2864 VDD.n2674 VDD.n772 185
R2865 VDD.n2327 VDD.n2326 185
R2866 VDD.n2326 VDD.n770 185
R2867 VDD.n2328 VDD.n778 185
R2868 VDD.n2668 VDD.n778 185
R2869 VDD.n2330 VDD.n2329 185
R2870 VDD.n2329 VDD.n785 185
R2871 VDD.n2331 VDD.n784 185
R2872 VDD.n2662 VDD.n784 185
R2873 VDD.n2333 VDD.n2332 185
R2874 VDD.n2332 VDD.n782 185
R2875 VDD.n2334 VDD.n791 185
R2876 VDD.n2656 VDD.n791 185
R2877 VDD.n2336 VDD.n2335 185
R2878 VDD.n2335 VDD.n789 185
R2879 VDD.n2337 VDD.n797 185
R2880 VDD.n2650 VDD.n797 185
R2881 VDD.n2339 VDD.n2338 185
R2882 VDD.n2338 VDD.n795 185
R2883 VDD.n2340 VDD.n803 185
R2884 VDD.n2644 VDD.n803 185
R2885 VDD.n2342 VDD.n2341 185
R2886 VDD.n2341 VDD.n801 185
R2887 VDD.n2343 VDD.n809 185
R2888 VDD.n2638 VDD.n809 185
R2889 VDD.n2345 VDD.n2344 185
R2890 VDD.n2344 VDD.n807 185
R2891 VDD.n2346 VDD.n815 185
R2892 VDD.n2632 VDD.n815 185
R2893 VDD.n2348 VDD.n2347 185
R2894 VDD.n2347 VDD.n813 185
R2895 VDD.n2349 VDD.n820 185
R2896 VDD.n2626 VDD.n820 185
R2897 VDD.n2351 VDD.n2350 185
R2898 VDD.n2350 VDD.n827 185
R2899 VDD.n2352 VDD.n826 185
R2900 VDD.n2620 VDD.n826 185
R2901 VDD.n2354 VDD.n2353 185
R2902 VDD.n2353 VDD.n824 185
R2903 VDD.n2355 VDD.n833 185
R2904 VDD.n2614 VDD.n833 185
R2905 VDD.n2357 VDD.n2356 185
R2906 VDD.n2356 VDD.n831 185
R2907 VDD.n2358 VDD.n839 185
R2908 VDD.n2608 VDD.n839 185
R2909 VDD.n2360 VDD.n2359 185
R2910 VDD.n2359 VDD.n837 185
R2911 VDD.n2361 VDD.n845 185
R2912 VDD.n2602 VDD.n845 185
R2913 VDD.n2363 VDD.n2362 185
R2914 VDD.n2362 VDD.n843 185
R2915 VDD.n2364 VDD.n851 185
R2916 VDD.n2596 VDD.n851 185
R2917 VDD.n2366 VDD.n2365 185
R2918 VDD.n2365 VDD.n849 185
R2919 VDD.n2367 VDD.n857 185
R2920 VDD.n2590 VDD.n857 185
R2921 VDD.n2369 VDD.n2368 185
R2922 VDD.n2368 VDD.n855 185
R2923 VDD.n2370 VDD.n863 185
R2924 VDD.n2584 VDD.n863 185
R2925 VDD.n2372 VDD.n2371 185
R2926 VDD.n2371 VDD.n861 185
R2927 VDD.n2373 VDD.n869 185
R2928 VDD.n2578 VDD.n869 185
R2929 VDD.n2375 VDD.n2374 185
R2930 VDD.n2374 VDD.n867 185
R2931 VDD.n2376 VDD.n875 185
R2932 VDD.n2572 VDD.n875 185
R2933 VDD.n2378 VDD.n2377 185
R2934 VDD.n2377 VDD.n873 185
R2935 VDD.n2379 VDD.n881 185
R2936 VDD.n2566 VDD.n881 185
R2937 VDD.n2381 VDD.n2380 185
R2938 VDD.n2380 VDD.n879 185
R2939 VDD.n2382 VDD.n887 185
R2940 VDD.n2560 VDD.n887 185
R2941 VDD.n2384 VDD.n2383 185
R2942 VDD.n2383 VDD.n885 185
R2943 VDD.n2385 VDD.n893 185
R2944 VDD.n2554 VDD.n893 185
R2945 VDD.n2387 VDD.n2386 185
R2946 VDD.n2386 VDD.n891 185
R2947 VDD.n2388 VDD.n898 185
R2948 VDD.n2548 VDD.n898 185
R2949 VDD.n2390 VDD.n2389 185
R2950 VDD.n2389 VDD.n905 185
R2951 VDD.n2391 VDD.n904 185
R2952 VDD.n2542 VDD.n904 185
R2953 VDD.n2393 VDD.n2392 185
R2954 VDD.n2392 VDD.n902 185
R2955 VDD.n2394 VDD.n911 185
R2956 VDD.n2536 VDD.n911 185
R2957 VDD.n2396 VDD.n2395 185
R2958 VDD.n2395 VDD.n909 185
R2959 VDD.n2397 VDD.n917 185
R2960 VDD.n2530 VDD.n917 185
R2961 VDD.n2399 VDD.n2398 185
R2962 VDD.n2398 VDD.n915 185
R2963 VDD.n2400 VDD.n923 185
R2964 VDD.n2524 VDD.n923 185
R2965 VDD.n2402 VDD.n2401 185
R2966 VDD.n2401 VDD.n921 185
R2967 VDD.n2403 VDD.n929 185
R2968 VDD.n2518 VDD.n929 185
R2969 VDD.n2405 VDD.n2404 185
R2970 VDD.n2404 VDD.n927 185
R2971 VDD.n2406 VDD.n935 185
R2972 VDD.n2512 VDD.n935 185
R2973 VDD.n2408 VDD.n2407 185
R2974 VDD.n2407 VDD.n933 185
R2975 VDD.n2409 VDD.n941 185
R2976 VDD.n2506 VDD.n941 185
R2977 VDD.n2411 VDD.n2410 185
R2978 VDD.n2410 VDD.n939 185
R2979 VDD.n2412 VDD.n946 185
R2980 VDD.n2500 VDD.n946 185
R2981 VDD.n2414 VDD.n2413 185
R2982 VDD.n2415 VDD.n2414 185
R2983 VDD.n2257 VDD.n952 185
R2984 VDD.n2494 VDD.n952 185
R2985 VDD.n2256 VDD.n2255 185
R2986 VDD.n2255 VDD.n950 185
R2987 VDD.n2254 VDD.n958 185
R2988 VDD.n2488 VDD.n958 185
R2989 VDD.n2253 VDD.n2252 185
R2990 VDD.n2252 VDD.n956 185
R2991 VDD.n2251 VDD.n964 185
R2992 VDD.n2482 VDD.n964 185
R2993 VDD.n2250 VDD.n2249 185
R2994 VDD.n2249 VDD.n962 185
R2995 VDD.n2248 VDD.n970 185
R2996 VDD.n2476 VDD.n970 185
R2997 VDD.n2247 VDD.n2246 185
R2998 VDD.n2246 VDD.n968 185
R2999 VDD.n2245 VDD.n976 185
R3000 VDD.n2470 VDD.n976 185
R3001 VDD.n2244 VDD.n2243 185
R3002 VDD.n2243 VDD.n974 185
R3003 VDD.n2209 VDD.n997 185
R3004 VDD.n2463 VDD.n997 185
R3005 VDD.n2211 VDD.n2210 185
R3006 VDD.n2213 VDD.n2212 185
R3007 VDD.n2215 VDD.n2214 185
R3008 VDD.n2217 VDD.n2216 185
R3009 VDD.n2219 VDD.n2218 185
R3010 VDD.n2221 VDD.n2220 185
R3011 VDD.n2223 VDD.n2222 185
R3012 VDD.n2225 VDD.n2224 185
R3013 VDD.n2227 VDD.n2226 185
R3014 VDD.n2229 VDD.n2228 185
R3015 VDD.n2231 VDD.n2230 185
R3016 VDD.n2233 VDD.n2232 185
R3017 VDD.n2235 VDD.n2234 185
R3018 VDD.n2237 VDD.n2236 185
R3019 VDD.n2239 VDD.n2238 185
R3020 VDD.n2241 VDD.n2240 185
R3021 VDD.n2242 VDD.n996 185
R3022 VDD.n2463 VDD.n996 185
R3023 VDD.t28 VDD.t131 156.564
R3024 VDD.t133 VDD.t27 156.564
R3025 VDD.n1206 VDD.t28 156.244
R3026 VDD.t27 VDD.n126 156.244
R3027 VDD.n3968 VDD.n120 146.341
R3028 VDD.n3978 VDD.n120 146.341
R3029 VDD.n3978 VDD.n116 146.341
R3030 VDD.n3984 VDD.n116 146.341
R3031 VDD.n3984 VDD.n108 146.341
R3032 VDD.n3994 VDD.n108 146.341
R3033 VDD.n3994 VDD.n104 146.341
R3034 VDD.n4000 VDD.n104 146.341
R3035 VDD.n4000 VDD.n96 146.341
R3036 VDD.n4010 VDD.n96 146.341
R3037 VDD.n4010 VDD.n92 146.341
R3038 VDD.n4016 VDD.n92 146.341
R3039 VDD.n4016 VDD.n84 146.341
R3040 VDD.n4026 VDD.n84 146.341
R3041 VDD.n4026 VDD.n80 146.341
R3042 VDD.n4032 VDD.n80 146.341
R3043 VDD.n4032 VDD.n72 146.341
R3044 VDD.n4043 VDD.n72 146.341
R3045 VDD.n4043 VDD.n68 146.341
R3046 VDD.n4049 VDD.n68 146.341
R3047 VDD.n4049 VDD.n61 146.341
R3048 VDD.n4059 VDD.n61 146.341
R3049 VDD.n4059 VDD.n57 146.341
R3050 VDD.n4065 VDD.n57 146.341
R3051 VDD.n4065 VDD.n49 146.341
R3052 VDD.n4075 VDD.n49 146.341
R3053 VDD.n4075 VDD.n45 146.341
R3054 VDD.n4081 VDD.n45 146.341
R3055 VDD.n4081 VDD.n34 146.341
R3056 VDD.n4602 VDD.n34 146.341
R3057 VDD.n4602 VDD.n35 146.341
R3058 VDD.n4595 VDD.n35 146.341
R3059 VDD.n4595 VDD.n4093 146.341
R3060 VDD.n4591 VDD.n4093 146.341
R3061 VDD.n4591 VDD.n4098 146.341
R3062 VDD.n4587 VDD.n4098 146.341
R3063 VDD.n4587 VDD.n4103 146.341
R3064 VDD.n4583 VDD.n4103 146.341
R3065 VDD.n4583 VDD.n4109 146.341
R3066 VDD.n4579 VDD.n4109 146.341
R3067 VDD.n4579 VDD.n4113 146.341
R3068 VDD.n4575 VDD.n4113 146.341
R3069 VDD.n4575 VDD.n4119 146.341
R3070 VDD.n4571 VDD.n4119 146.341
R3071 VDD.n4571 VDD.n4125 146.341
R3072 VDD.n4567 VDD.n4125 146.341
R3073 VDD.n4567 VDD.n4131 146.341
R3074 VDD.n4563 VDD.n4131 146.341
R3075 VDD.n4563 VDD.n4136 146.341
R3076 VDD.n4559 VDD.n4136 146.341
R3077 VDD.n4559 VDD.n4142 146.341
R3078 VDD.n4555 VDD.n4142 146.341
R3079 VDD.n4555 VDD.n4147 146.341
R3080 VDD.n4551 VDD.n4147 146.341
R3081 VDD.n4551 VDD.n4153 146.341
R3082 VDD.n4547 VDD.n4153 146.341
R3083 VDD.n4547 VDD.n4158 146.341
R3084 VDD.n4543 VDD.n4158 146.341
R3085 VDD.n4543 VDD.n4164 146.341
R3086 VDD.n4539 VDD.n4164 146.341
R3087 VDD.n4532 VDD.n4173 146.341
R3088 VDD.n4530 VDD.n4529 146.341
R3089 VDD.n4527 VDD.n4177 146.341
R3090 VDD.n4523 VDD.n4522 146.341
R3091 VDD.n4520 VDD.n4185 146.341
R3092 VDD.n4516 VDD.n4515 146.341
R3093 VDD.n4513 VDD.n4192 146.341
R3094 VDD.n4506 VDD.n4505 146.341
R3095 VDD.n4503 VDD.n4199 146.341
R3096 VDD.n4499 VDD.n4498 146.341
R3097 VDD.n4496 VDD.n4206 146.341
R3098 VDD.n4492 VDD.n4491 146.341
R3099 VDD.n4489 VDD.n4213 146.341
R3100 VDD.n4485 VDD.n4484 146.341
R3101 VDD.n4482 VDD.n4220 146.341
R3102 VDD.n4478 VDD.n4477 146.341
R3103 VDD.n4475 VDD.n4230 146.341
R3104 VDD.n4471 VDD.n4470 146.341
R3105 VDD.n4468 VDD.n4237 146.341
R3106 VDD.n4464 VDD.n4463 146.341
R3107 VDD.n4461 VDD.n4244 146.341
R3108 VDD.n4457 VDD.n4456 146.341
R3109 VDD.n4454 VDD.n4251 146.341
R3110 VDD.n4450 VDD.n4449 146.341
R3111 VDD.n4447 VDD.n4260 146.341
R3112 VDD.n4441 VDD.n4440 146.341
R3113 VDD.n4438 VDD.n4266 146.341
R3114 VDD.n4434 VDD.n4433 146.341
R3115 VDD.n4431 VDD.n4272 146.341
R3116 VDD.n4427 VDD.n4426 146.341
R3117 VDD.n4424 VDD.n4279 146.341
R3118 VDD.n4420 VDD.n4419 146.341
R3119 VDD.n4417 VDD.n4286 146.341
R3120 VDD.n4411 VDD.n4410 146.341
R3121 VDD.n4408 VDD.n4294 146.341
R3122 VDD.n4404 VDD.n4403 146.341
R3123 VDD.n4401 VDD.n4300 146.341
R3124 VDD.n4397 VDD.n4396 146.341
R3125 VDD.n4394 VDD.n4307 146.341
R3126 VDD.n4390 VDD.n4389 146.341
R3127 VDD.n4387 VDD.n4314 146.341
R3128 VDD.n3970 VDD.n122 146.341
R3129 VDD.n3976 VDD.n122 146.341
R3130 VDD.n3976 VDD.n113 146.341
R3131 VDD.n3986 VDD.n113 146.341
R3132 VDD.n3986 VDD.n109 146.341
R3133 VDD.n3992 VDD.n109 146.341
R3134 VDD.n3992 VDD.n102 146.341
R3135 VDD.n4002 VDD.n102 146.341
R3136 VDD.n4002 VDD.n98 146.341
R3137 VDD.n4008 VDD.n98 146.341
R3138 VDD.n4008 VDD.n90 146.341
R3139 VDD.n4018 VDD.n90 146.341
R3140 VDD.n4018 VDD.n86 146.341
R3141 VDD.n4024 VDD.n86 146.341
R3142 VDD.n4024 VDD.n78 146.341
R3143 VDD.n4034 VDD.n78 146.341
R3144 VDD.n4034 VDD.n74 146.341
R3145 VDD.n4040 VDD.n74 146.341
R3146 VDD.n4040 VDD.n67 146.341
R3147 VDD.n4051 VDD.n67 146.341
R3148 VDD.n4051 VDD.n63 146.341
R3149 VDD.n4057 VDD.n63 146.341
R3150 VDD.n4057 VDD.n55 146.341
R3151 VDD.n4067 VDD.n55 146.341
R3152 VDD.n4067 VDD.n51 146.341
R3153 VDD.n4073 VDD.n51 146.341
R3154 VDD.n4073 VDD.n43 146.341
R3155 VDD.n4083 VDD.n43 146.341
R3156 VDD.n4083 VDD.n38 146.341
R3157 VDD.n4601 VDD.n38 146.341
R3158 VDD.n4601 VDD.n39 146.341
R3159 VDD.n4597 VDD.n39 146.341
R3160 VDD.n4597 VDD.n4091 146.341
R3161 VDD.n4099 VDD.n4091 146.341
R3162 VDD.n4100 VDD.n4099 146.341
R3163 VDD.n4101 VDD.n4100 146.341
R3164 VDD.n4338 VDD.n4101 146.341
R3165 VDD.n4338 VDD.n4110 146.341
R3166 VDD.n4111 VDD.n4110 146.341
R3167 VDD.n4112 VDD.n4111 146.341
R3168 VDD.n4335 VDD.n4112 146.341
R3169 VDD.n4335 VDD.n4121 146.341
R3170 VDD.n4122 VDD.n4121 146.341
R3171 VDD.n4123 VDD.n4122 146.341
R3172 VDD.n4332 VDD.n4123 146.341
R3173 VDD.n4332 VDD.n4132 146.341
R3174 VDD.n4133 VDD.n4132 146.341
R3175 VDD.n4134 VDD.n4133 146.341
R3176 VDD.n4329 VDD.n4134 146.341
R3177 VDD.n4329 VDD.n4143 146.341
R3178 VDD.n4144 VDD.n4143 146.341
R3179 VDD.n4145 VDD.n4144 146.341
R3180 VDD.n4326 VDD.n4145 146.341
R3181 VDD.n4326 VDD.n4154 146.341
R3182 VDD.n4155 VDD.n4154 146.341
R3183 VDD.n4156 VDD.n4155 146.341
R3184 VDD.n4323 VDD.n4156 146.341
R3185 VDD.n4323 VDD.n4165 146.341
R3186 VDD.n4166 VDD.n4165 146.341
R3187 VDD.n4167 VDD.n4166 146.341
R3188 VDD.n3962 VDD.n3960 146.341
R3189 VDD.n3960 VDD.n3959 146.341
R3190 VDD.n3956 VDD.n3955 146.341
R3191 VDD.n3953 VDD.n135 146.341
R3192 VDD.n3949 VDD.n3947 146.341
R3193 VDD.n3945 VDD.n141 146.341
R3194 VDD.n3941 VDD.n3939 146.341
R3195 VDD.n3937 VDD.n147 146.341
R3196 VDD.n3932 VDD.n3930 146.341
R3197 VDD.n3928 VDD.n155 146.341
R3198 VDD.n3924 VDD.n3922 146.341
R3199 VDD.n3920 VDD.n161 146.341
R3200 VDD.n168 VDD.n167 146.341
R3201 VDD.n3912 VDD.n3910 146.341
R3202 VDD.n3908 VDD.n170 146.341
R3203 VDD.n3904 VDD.n3902 146.341
R3204 VDD.n3900 VDD.n176 146.341
R3205 VDD.n3896 VDD.n3894 146.341
R3206 VDD.n3892 VDD.n185 146.341
R3207 VDD.n3888 VDD.n3886 146.341
R3208 VDD.n3884 VDD.n191 146.341
R3209 VDD.n3880 VDD.n3878 146.341
R3210 VDD.n3876 VDD.n197 146.341
R3211 VDD.n3872 VDD.n3870 146.341
R3212 VDD.n3868 VDD.n203 146.341
R3213 VDD.n3864 VDD.n3862 146.341
R3214 VDD.n3860 VDD.n211 146.341
R3215 VDD.n3856 VDD.n3854 146.341
R3216 VDD.n3852 VDD.n217 146.341
R3217 VDD.n3848 VDD.n3846 146.341
R3218 VDD.n3843 VDD.n3842 146.341
R3219 VDD.n3839 VDD.n3838 146.341
R3220 VDD.n3836 VDD.n3765 146.341
R3221 VDD.n3827 VDD.n3772 146.341
R3222 VDD.n3825 VDD.n3824 146.341
R3223 VDD.n3821 VDD.n3820 146.341
R3224 VDD.n3818 VDD.n3777 146.341
R3225 VDD.n3814 VDD.n3812 146.341
R3226 VDD.n3810 VDD.n3783 146.341
R3227 VDD.n3806 VDD.n3804 146.341
R3228 VDD.n3802 VDD.n3789 146.341
R3229 VDD.n3794 VDD.n125 146.341
R3230 VDD.n2163 VDD.n2162 146.341
R3231 VDD.n2160 VDD.n1953 146.341
R3232 VDD.n2156 VDD.n2155 146.341
R3233 VDD.n2153 VDD.n1960 146.341
R3234 VDD.n2149 VDD.n2148 146.341
R3235 VDD.n2146 VDD.n1967 146.341
R3236 VDD.n2142 VDD.n2141 146.341
R3237 VDD.n2139 VDD.n1974 146.341
R3238 VDD.n2135 VDD.n2134 146.341
R3239 VDD.n2132 VDD.n1984 146.341
R3240 VDD.n2128 VDD.n2127 146.341
R3241 VDD.n2125 VDD.n1991 146.341
R3242 VDD.n2118 VDD.n1997 146.341
R3243 VDD.n2116 VDD.n2115 146.341
R3244 VDD.n2113 VDD.n1999 146.341
R3245 VDD.n2109 VDD.n2108 146.341
R3246 VDD.n2106 VDD.n2009 146.341
R3247 VDD.n2102 VDD.n2101 146.341
R3248 VDD.n2099 VDD.n2016 146.341
R3249 VDD.n2095 VDD.n2094 146.341
R3250 VDD.n2092 VDD.n2023 146.341
R3251 VDD.n2088 VDD.n2087 146.341
R3252 VDD.n2085 VDD.n2030 146.341
R3253 VDD.n2081 VDD.n2080 146.341
R3254 VDD.n2078 VDD.n2039 146.341
R3255 VDD.n2072 VDD.n2071 146.341
R3256 VDD.n2069 VDD.n2045 146.341
R3257 VDD.n2065 VDD.n2064 146.341
R3258 VDD.n2062 VDD.n2059 146.341
R3259 VDD.n2057 VDD.n2054 146.341
R3260 VDD.n2052 VDD.n1161 146.341
R3261 VDD.n1163 VDD.n1162 146.341
R3262 VDD.n1193 VDD.n1168 146.341
R3263 VDD.n1170 VDD.n1169 146.341
R3264 VDD.n1196 VDD.n1173 146.341
R3265 VDD.n1175 VDD.n1174 146.341
R3266 VDD.n1199 VDD.n1178 146.341
R3267 VDD.n1180 VDD.n1179 146.341
R3268 VDD.n1202 VDD.n1183 146.341
R3269 VDD.n1185 VDD.n1184 146.341
R3270 VDD.n2174 VDD.n1191 146.341
R3271 VDD.n1697 VDD.n1385 146.341
R3272 VDD.n1703 VDD.n1385 146.341
R3273 VDD.n1703 VDD.n1376 146.341
R3274 VDD.n1713 VDD.n1376 146.341
R3275 VDD.n1713 VDD.n1372 146.341
R3276 VDD.n1719 VDD.n1372 146.341
R3277 VDD.n1719 VDD.n1365 146.341
R3278 VDD.n1729 VDD.n1365 146.341
R3279 VDD.n1729 VDD.n1361 146.341
R3280 VDD.n1735 VDD.n1361 146.341
R3281 VDD.n1735 VDD.n1353 146.341
R3282 VDD.n1745 VDD.n1353 146.341
R3283 VDD.n1745 VDD.n1349 146.341
R3284 VDD.n1751 VDD.n1349 146.341
R3285 VDD.n1751 VDD.n1341 146.341
R3286 VDD.n1761 VDD.n1341 146.341
R3287 VDD.n1761 VDD.n1337 146.341
R3288 VDD.n1767 VDD.n1337 146.341
R3289 VDD.n1767 VDD.n1330 146.341
R3290 VDD.n1778 VDD.n1330 146.341
R3291 VDD.n1778 VDD.n1326 146.341
R3292 VDD.n1784 VDD.n1326 146.341
R3293 VDD.n1784 VDD.n1318 146.341
R3294 VDD.n1794 VDD.n1318 146.341
R3295 VDD.n1794 VDD.n1314 146.341
R3296 VDD.n1800 VDD.n1314 146.341
R3297 VDD.n1800 VDD.n1306 146.341
R3298 VDD.n1810 VDD.n1306 146.341
R3299 VDD.n1810 VDD.n1302 146.341
R3300 VDD.n1816 VDD.n1302 146.341
R3301 VDD.n1816 VDD.n1294 146.341
R3302 VDD.n1840 VDD.n1294 146.341
R3303 VDD.n1840 VDD.n1290 146.341
R3304 VDD.n1846 VDD.n1290 146.341
R3305 VDD.n1846 VDD.n1282 146.341
R3306 VDD.n1856 VDD.n1282 146.341
R3307 VDD.n1856 VDD.n1278 146.341
R3308 VDD.n1862 VDD.n1278 146.341
R3309 VDD.n1862 VDD.n1270 146.341
R3310 VDD.n1872 VDD.n1270 146.341
R3311 VDD.n1872 VDD.n1266 146.341
R3312 VDD.n1878 VDD.n1266 146.341
R3313 VDD.n1878 VDD.n1258 146.341
R3314 VDD.n1888 VDD.n1258 146.341
R3315 VDD.n1888 VDD.n1254 146.341
R3316 VDD.n1894 VDD.n1254 146.341
R3317 VDD.n1894 VDD.n1246 146.341
R3318 VDD.n1904 VDD.n1246 146.341
R3319 VDD.n1904 VDD.n1242 146.341
R3320 VDD.n1910 VDD.n1242 146.341
R3321 VDD.n1910 VDD.n1234 146.341
R3322 VDD.n1920 VDD.n1234 146.341
R3323 VDD.n1920 VDD.n1230 146.341
R3324 VDD.n1926 VDD.n1230 146.341
R3325 VDD.n1926 VDD.n1222 146.341
R3326 VDD.n1936 VDD.n1222 146.341
R3327 VDD.n1936 VDD.n1217 146.341
R3328 VDD.n1944 VDD.n1217 146.341
R3329 VDD.n1944 VDD.n1207 146.341
R3330 VDD.n2171 VDD.n1207 146.341
R3331 VDD.n1394 VDD.n1393 146.341
R3332 VDD.n1397 VDD.n1394 146.341
R3333 VDD.n1400 VDD.n1399 146.341
R3334 VDD.n1405 VDD.n1402 146.341
R3335 VDD.n1408 VDD.n1407 146.341
R3336 VDD.n1413 VDD.n1410 146.341
R3337 VDD.n1416 VDD.n1415 146.341
R3338 VDD.n1423 VDD.n1418 146.341
R3339 VDD.n1426 VDD.n1425 146.341
R3340 VDD.n1431 VDD.n1430 146.341
R3341 VDD.n1434 VDD.n1433 146.341
R3342 VDD.n1439 VDD.n1438 146.341
R3343 VDD.n1442 VDD.n1441 146.341
R3344 VDD.n1447 VDD.n1446 146.341
R3345 VDD.n1450 VDD.n1449 146.341
R3346 VDD.n1455 VDD.n1454 146.341
R3347 VDD.n1458 VDD.n1457 146.341
R3348 VDD.n1463 VDD.n1462 146.341
R3349 VDD.n1466 VDD.n1465 146.341
R3350 VDD.n1471 VDD.n1470 146.341
R3351 VDD.n1474 VDD.n1473 146.341
R3352 VDD.n1479 VDD.n1478 146.341
R3353 VDD.n1482 VDD.n1481 146.341
R3354 VDD.n1487 VDD.n1486 146.341
R3355 VDD.n1614 VDD.n1489 146.341
R3356 VDD.n1612 VDD.n1611 146.341
R3357 VDD.n1499 VDD.n1498 146.341
R3358 VDD.n1502 VDD.n1501 146.341
R3359 VDD.n1507 VDD.n1506 146.341
R3360 VDD.n1510 VDD.n1509 146.341
R3361 VDD.n1515 VDD.n1514 146.341
R3362 VDD.n1518 VDD.n1517 146.341
R3363 VDD.n1585 VDD.n1523 146.341
R3364 VDD.n1583 VDD.n1582 146.341
R3365 VDD.n1528 VDD.n1527 146.341
R3366 VDD.n1531 VDD.n1530 146.341
R3367 VDD.n1536 VDD.n1535 146.341
R3368 VDD.n1539 VDD.n1538 146.341
R3369 VDD.n1544 VDD.n1543 146.341
R3370 VDD.n1547 VDD.n1546 146.341
R3371 VDD.n1552 VDD.n1551 146.341
R3372 VDD.n1555 VDD.n1388 146.341
R3373 VDD.n1695 VDD.n1383 146.341
R3374 VDD.n1705 VDD.n1383 146.341
R3375 VDD.n1705 VDD.n1379 146.341
R3376 VDD.n1711 VDD.n1379 146.341
R3377 VDD.n1711 VDD.n1371 146.341
R3378 VDD.n1721 VDD.n1371 146.341
R3379 VDD.n1721 VDD.n1367 146.341
R3380 VDD.n1727 VDD.n1367 146.341
R3381 VDD.n1727 VDD.n1359 146.341
R3382 VDD.n1737 VDD.n1359 146.341
R3383 VDD.n1737 VDD.n1355 146.341
R3384 VDD.n1743 VDD.n1355 146.341
R3385 VDD.n1743 VDD.n1347 146.341
R3386 VDD.n1753 VDD.n1347 146.341
R3387 VDD.n1753 VDD.n1343 146.341
R3388 VDD.n1759 VDD.n1343 146.341
R3389 VDD.n1759 VDD.n1335 146.341
R3390 VDD.n1770 VDD.n1335 146.341
R3391 VDD.n1770 VDD.n1331 146.341
R3392 VDD.n1776 VDD.n1331 146.341
R3393 VDD.n1776 VDD.n1324 146.341
R3394 VDD.n1786 VDD.n1324 146.341
R3395 VDD.n1786 VDD.n1320 146.341
R3396 VDD.n1792 VDD.n1320 146.341
R3397 VDD.n1792 VDD.n1312 146.341
R3398 VDD.n1802 VDD.n1312 146.341
R3399 VDD.n1802 VDD.n1308 146.341
R3400 VDD.n1808 VDD.n1308 146.341
R3401 VDD.n1808 VDD.n1300 146.341
R3402 VDD.n1817 VDD.n1300 146.341
R3403 VDD.n1817 VDD.n1296 146.341
R3404 VDD.n1838 VDD.n1296 146.341
R3405 VDD.n1838 VDD.n1288 146.341
R3406 VDD.n1848 VDD.n1288 146.341
R3407 VDD.n1848 VDD.n1284 146.341
R3408 VDD.n1854 VDD.n1284 146.341
R3409 VDD.n1854 VDD.n1276 146.341
R3410 VDD.n1864 VDD.n1276 146.341
R3411 VDD.n1864 VDD.n1272 146.341
R3412 VDD.n1870 VDD.n1272 146.341
R3413 VDD.n1870 VDD.n1264 146.341
R3414 VDD.n1880 VDD.n1264 146.341
R3415 VDD.n1880 VDD.n1260 146.341
R3416 VDD.n1886 VDD.n1260 146.341
R3417 VDD.n1886 VDD.n1252 146.341
R3418 VDD.n1896 VDD.n1252 146.341
R3419 VDD.n1896 VDD.n1248 146.341
R3420 VDD.n1902 VDD.n1248 146.341
R3421 VDD.n1902 VDD.n1240 146.341
R3422 VDD.n1912 VDD.n1240 146.341
R3423 VDD.n1912 VDD.n1236 146.341
R3424 VDD.n1918 VDD.n1236 146.341
R3425 VDD.n1918 VDD.n1228 146.341
R3426 VDD.n1928 VDD.n1228 146.341
R3427 VDD.n1928 VDD.n1224 146.341
R3428 VDD.n1934 VDD.n1224 146.341
R3429 VDD.n1934 VDD.n1215 146.341
R3430 VDD.n1946 VDD.n1215 146.341
R3431 VDD.n1946 VDD.n1210 146.341
R3432 VDD.n2169 VDD.n1210 146.341
R3433 VDD.n9 VDD.n7 137.044
R3434 VDD.n2 VDD.n0 137.044
R3435 VDD.n9 VDD.n8 135.334
R3436 VDD.n11 VDD.n10 135.334
R3437 VDD.n13 VDD.n12 135.334
R3438 VDD.n6 VDD.n5 135.334
R3439 VDD.n4 VDD.n3 135.334
R3440 VDD.n2 VDD.n1 135.334
R3441 VDD.n1155 VDD.t47 134.12
R3442 VDD.n625 VDD.t117 134.12
R3443 VDD.n254 VDD.t32 134.12
R3444 VDD.n2901 VDD.t70 134.12
R3445 VDD.n635 VDD.t84 134.12
R3446 VDD.n1001 VDD.t110 134.12
R3447 VDD.n231 VDD.t80 134.12
R3448 VDD.n3121 VDD.t119 134.12
R3449 VDD.t131 VDD.t137 126.398
R3450 VDD.t159 VDD.t133 126.398
R3451 VDD.n4321 VDD.n4320 103.758
R3452 VDD.n178 VDD.n177 103.758
R3453 VDD.n3833 VDD.n3832 103.758
R3454 VDD.n1155 VDD.n1154 102.594
R3455 VDD.n625 VDD.n624 102.594
R3456 VDD.n254 VDD.n253 102.594
R3457 VDD.n2901 VDD.n2900 102.594
R3458 VDD.n635 VDD.n634 102.594
R3459 VDD.n1001 VDD.n1000 102.594
R3460 VDD.n231 VDD.n230 102.594
R3461 VDD.n3121 VDD.n3120 102.594
R3462 VDD.n3738 VDD.n3737 99.5127
R3463 VDD.n3735 VDD.n246 99.5127
R3464 VDD.n3731 VDD.n3730 99.5127
R3465 VDD.n3728 VDD.n3725 99.5127
R3466 VDD.n3723 VDD.n249 99.5127
R3467 VDD.n3719 VDD.n3718 99.5127
R3468 VDD.n3716 VDD.n252 99.5127
R3469 VDD.n3712 VDD.n3711 99.5127
R3470 VDD.n3111 VDD.n2898 99.5127
R3471 VDD.n2898 VDD.n597 99.5127
R3472 VDD.n3106 VDD.n597 99.5127
R3473 VDD.n3106 VDD.n591 99.5127
R3474 VDD.n3103 VDD.n591 99.5127
R3475 VDD.n3103 VDD.n585 99.5127
R3476 VDD.n3100 VDD.n585 99.5127
R3477 VDD.n3100 VDD.n579 99.5127
R3478 VDD.n3097 VDD.n579 99.5127
R3479 VDD.n3097 VDD.n573 99.5127
R3480 VDD.n3094 VDD.n573 99.5127
R3481 VDD.n3094 VDD.n567 99.5127
R3482 VDD.n3091 VDD.n567 99.5127
R3483 VDD.n3091 VDD.n561 99.5127
R3484 VDD.n3088 VDD.n561 99.5127
R3485 VDD.n3088 VDD.n555 99.5127
R3486 VDD.n3085 VDD.n555 99.5127
R3487 VDD.n3085 VDD.n549 99.5127
R3488 VDD.n3082 VDD.n549 99.5127
R3489 VDD.n3082 VDD.n543 99.5127
R3490 VDD.n3079 VDD.n543 99.5127
R3491 VDD.n3079 VDD.n537 99.5127
R3492 VDD.n3076 VDD.n537 99.5127
R3493 VDD.n3076 VDD.n531 99.5127
R3494 VDD.n3073 VDD.n531 99.5127
R3495 VDD.n3073 VDD.n525 99.5127
R3496 VDD.n3070 VDD.n525 99.5127
R3497 VDD.n3070 VDD.n519 99.5127
R3498 VDD.n3067 VDD.n519 99.5127
R3499 VDD.n3067 VDD.n512 99.5127
R3500 VDD.n3064 VDD.n512 99.5127
R3501 VDD.n3064 VDD.n506 99.5127
R3502 VDD.n3061 VDD.n506 99.5127
R3503 VDD.n3061 VDD.n501 99.5127
R3504 VDD.n3058 VDD.n501 99.5127
R3505 VDD.n3058 VDD.n495 99.5127
R3506 VDD.n3055 VDD.n495 99.5127
R3507 VDD.n3055 VDD.n489 99.5127
R3508 VDD.n3052 VDD.n489 99.5127
R3509 VDD.n3052 VDD.n483 99.5127
R3510 VDD.n3049 VDD.n483 99.5127
R3511 VDD.n3049 VDD.n477 99.5127
R3512 VDD.n3046 VDD.n477 99.5127
R3513 VDD.n3046 VDD.n470 99.5127
R3514 VDD.n3043 VDD.n470 99.5127
R3515 VDD.n3043 VDD.n464 99.5127
R3516 VDD.n3040 VDD.n464 99.5127
R3517 VDD.n3040 VDD.n458 99.5127
R3518 VDD.n3037 VDD.n458 99.5127
R3519 VDD.n3037 VDD.n452 99.5127
R3520 VDD.n3034 VDD.n452 99.5127
R3521 VDD.n3034 VDD.n447 99.5127
R3522 VDD.n3031 VDD.n447 99.5127
R3523 VDD.n3031 VDD.n441 99.5127
R3524 VDD.n3028 VDD.n441 99.5127
R3525 VDD.n3028 VDD.n435 99.5127
R3526 VDD.n3025 VDD.n435 99.5127
R3527 VDD.n3025 VDD.n429 99.5127
R3528 VDD.n3022 VDD.n429 99.5127
R3529 VDD.n3022 VDD.n423 99.5127
R3530 VDD.n3019 VDD.n423 99.5127
R3531 VDD.n3019 VDD.n416 99.5127
R3532 VDD.n3016 VDD.n416 99.5127
R3533 VDD.n3016 VDD.n410 99.5127
R3534 VDD.n3013 VDD.n410 99.5127
R3535 VDD.n3013 VDD.n405 99.5127
R3536 VDD.n3010 VDD.n405 99.5127
R3537 VDD.n3010 VDD.n399 99.5127
R3538 VDD.n3007 VDD.n399 99.5127
R3539 VDD.n3007 VDD.n393 99.5127
R3540 VDD.n3004 VDD.n393 99.5127
R3541 VDD.n3004 VDD.n387 99.5127
R3542 VDD.n3001 VDD.n387 99.5127
R3543 VDD.n3001 VDD.n381 99.5127
R3544 VDD.n2998 VDD.n381 99.5127
R3545 VDD.n2998 VDD.n375 99.5127
R3546 VDD.n2995 VDD.n375 99.5127
R3547 VDD.n2995 VDD.n369 99.5127
R3548 VDD.n2992 VDD.n369 99.5127
R3549 VDD.n2992 VDD.n363 99.5127
R3550 VDD.n2989 VDD.n363 99.5127
R3551 VDD.n2989 VDD.n357 99.5127
R3552 VDD.n2986 VDD.n357 99.5127
R3553 VDD.n2986 VDD.n351 99.5127
R3554 VDD.n2983 VDD.n351 99.5127
R3555 VDD.n2983 VDD.n345 99.5127
R3556 VDD.n2980 VDD.n345 99.5127
R3557 VDD.n2980 VDD.n338 99.5127
R3558 VDD.n2977 VDD.n338 99.5127
R3559 VDD.n2977 VDD.n332 99.5127
R3560 VDD.n2974 VDD.n332 99.5127
R3561 VDD.n2974 VDD.n327 99.5127
R3562 VDD.n2971 VDD.n327 99.5127
R3563 VDD.n2971 VDD.n321 99.5127
R3564 VDD.n2968 VDD.n321 99.5127
R3565 VDD.n2968 VDD.n315 99.5127
R3566 VDD.n2965 VDD.n315 99.5127
R3567 VDD.n2965 VDD.n309 99.5127
R3568 VDD.n2962 VDD.n309 99.5127
R3569 VDD.n2962 VDD.n303 99.5127
R3570 VDD.n2959 VDD.n303 99.5127
R3571 VDD.n2959 VDD.n297 99.5127
R3572 VDD.n2956 VDD.n297 99.5127
R3573 VDD.n2956 VDD.n290 99.5127
R3574 VDD.n2953 VDD.n290 99.5127
R3575 VDD.n2953 VDD.n284 99.5127
R3576 VDD.n2950 VDD.n284 99.5127
R3577 VDD.n2950 VDD.n279 99.5127
R3578 VDD.n2947 VDD.n279 99.5127
R3579 VDD.n2947 VDD.n273 99.5127
R3580 VDD.n2944 VDD.n273 99.5127
R3581 VDD.n2944 VDD.n266 99.5127
R3582 VDD.n266 VDD.n258 99.5127
R3583 VDD.n3704 VDD.n258 99.5127
R3584 VDD.n3705 VDD.n3704 99.5127
R3585 VDD.n3705 VDD.n239 99.5127
R3586 VDD.n2912 VDD.n2911 99.5127
R3587 VDD.n2914 VDD.n2912 99.5127
R3588 VDD.n2918 VDD.n2907 99.5127
R3589 VDD.n2922 VDD.n2920 99.5127
R3590 VDD.n2926 VDD.n2905 99.5127
R3591 VDD.n2930 VDD.n2928 99.5127
R3592 VDD.n2934 VDD.n2903 99.5127
R3593 VDD.n2937 VDD.n2936 99.5127
R3594 VDD.n2939 VDD.n2897 99.5127
R3595 VDD.n3336 VDD.n599 99.5127
R3596 VDD.n3340 VDD.n599 99.5127
R3597 VDD.n3340 VDD.n589 99.5127
R3598 VDD.n3348 VDD.n589 99.5127
R3599 VDD.n3348 VDD.n587 99.5127
R3600 VDD.n3352 VDD.n587 99.5127
R3601 VDD.n3352 VDD.n577 99.5127
R3602 VDD.n3360 VDD.n577 99.5127
R3603 VDD.n3360 VDD.n575 99.5127
R3604 VDD.n3364 VDD.n575 99.5127
R3605 VDD.n3364 VDD.n565 99.5127
R3606 VDD.n3372 VDD.n565 99.5127
R3607 VDD.n3372 VDD.n563 99.5127
R3608 VDD.n3376 VDD.n563 99.5127
R3609 VDD.n3376 VDD.n553 99.5127
R3610 VDD.n3384 VDD.n553 99.5127
R3611 VDD.n3384 VDD.n551 99.5127
R3612 VDD.n3388 VDD.n551 99.5127
R3613 VDD.n3388 VDD.n541 99.5127
R3614 VDD.n3396 VDD.n541 99.5127
R3615 VDD.n3396 VDD.n539 99.5127
R3616 VDD.n3400 VDD.n539 99.5127
R3617 VDD.n3400 VDD.n529 99.5127
R3618 VDD.n3408 VDD.n529 99.5127
R3619 VDD.n3408 VDD.n527 99.5127
R3620 VDD.n3412 VDD.n527 99.5127
R3621 VDD.n3412 VDD.n517 99.5127
R3622 VDD.n3420 VDD.n517 99.5127
R3623 VDD.n3420 VDD.n515 99.5127
R3624 VDD.n3424 VDD.n515 99.5127
R3625 VDD.n3424 VDD.n505 99.5127
R3626 VDD.n3432 VDD.n505 99.5127
R3627 VDD.n3432 VDD.n503 99.5127
R3628 VDD.n3436 VDD.n503 99.5127
R3629 VDD.n3436 VDD.n493 99.5127
R3630 VDD.n3444 VDD.n493 99.5127
R3631 VDD.n3444 VDD.n491 99.5127
R3632 VDD.n3448 VDD.n491 99.5127
R3633 VDD.n3448 VDD.n481 99.5127
R3634 VDD.n3456 VDD.n481 99.5127
R3635 VDD.n3456 VDD.n479 99.5127
R3636 VDD.n3460 VDD.n479 99.5127
R3637 VDD.n3460 VDD.n468 99.5127
R3638 VDD.n3468 VDD.n468 99.5127
R3639 VDD.n3468 VDD.n466 99.5127
R3640 VDD.n3472 VDD.n466 99.5127
R3641 VDD.n3472 VDD.n456 99.5127
R3642 VDD.n3480 VDD.n456 99.5127
R3643 VDD.n3480 VDD.n454 99.5127
R3644 VDD.n3484 VDD.n454 99.5127
R3645 VDD.n3484 VDD.n445 99.5127
R3646 VDD.n3492 VDD.n445 99.5127
R3647 VDD.n3492 VDD.n443 99.5127
R3648 VDD.n3496 VDD.n443 99.5127
R3649 VDD.n3496 VDD.n433 99.5127
R3650 VDD.n3504 VDD.n433 99.5127
R3651 VDD.n3504 VDD.n431 99.5127
R3652 VDD.n3508 VDD.n431 99.5127
R3653 VDD.n3508 VDD.n421 99.5127
R3654 VDD.n3516 VDD.n421 99.5127
R3655 VDD.n3516 VDD.n419 99.5127
R3656 VDD.n3520 VDD.n419 99.5127
R3657 VDD.n3520 VDD.n409 99.5127
R3658 VDD.n3528 VDD.n409 99.5127
R3659 VDD.n3528 VDD.n407 99.5127
R3660 VDD.n3532 VDD.n407 99.5127
R3661 VDD.n3532 VDD.n397 99.5127
R3662 VDD.n3540 VDD.n397 99.5127
R3663 VDD.n3540 VDD.n395 99.5127
R3664 VDD.n3544 VDD.n395 99.5127
R3665 VDD.n3544 VDD.n385 99.5127
R3666 VDD.n3552 VDD.n385 99.5127
R3667 VDD.n3552 VDD.n383 99.5127
R3668 VDD.n3556 VDD.n383 99.5127
R3669 VDD.n3556 VDD.n373 99.5127
R3670 VDD.n3564 VDD.n373 99.5127
R3671 VDD.n3564 VDD.n371 99.5127
R3672 VDD.n3568 VDD.n371 99.5127
R3673 VDD.n3568 VDD.n361 99.5127
R3674 VDD.n3576 VDD.n361 99.5127
R3675 VDD.n3576 VDD.n359 99.5127
R3676 VDD.n3580 VDD.n359 99.5127
R3677 VDD.n3580 VDD.n349 99.5127
R3678 VDD.n3588 VDD.n349 99.5127
R3679 VDD.n3588 VDD.n347 99.5127
R3680 VDD.n3592 VDD.n347 99.5127
R3681 VDD.n3592 VDD.n336 99.5127
R3682 VDD.n3600 VDD.n336 99.5127
R3683 VDD.n3600 VDD.n334 99.5127
R3684 VDD.n3604 VDD.n334 99.5127
R3685 VDD.n3604 VDD.n325 99.5127
R3686 VDD.n3612 VDD.n325 99.5127
R3687 VDD.n3612 VDD.n323 99.5127
R3688 VDD.n3616 VDD.n323 99.5127
R3689 VDD.n3616 VDD.n313 99.5127
R3690 VDD.n3624 VDD.n313 99.5127
R3691 VDD.n3624 VDD.n311 99.5127
R3692 VDD.n3628 VDD.n311 99.5127
R3693 VDD.n3628 VDD.n301 99.5127
R3694 VDD.n3636 VDD.n301 99.5127
R3695 VDD.n3636 VDD.n299 99.5127
R3696 VDD.n3640 VDD.n299 99.5127
R3697 VDD.n3640 VDD.n288 99.5127
R3698 VDD.n3648 VDD.n288 99.5127
R3699 VDD.n3648 VDD.n286 99.5127
R3700 VDD.n3652 VDD.n286 99.5127
R3701 VDD.n3652 VDD.n277 99.5127
R3702 VDD.n3660 VDD.n277 99.5127
R3703 VDD.n3660 VDD.n275 99.5127
R3704 VDD.n3664 VDD.n275 99.5127
R3705 VDD.n3664 VDD.n264 99.5127
R3706 VDD.n3698 VDD.n264 99.5127
R3707 VDD.n3698 VDD.n262 99.5127
R3708 VDD.n3702 VDD.n262 99.5127
R3709 VDD.n3702 VDD.n241 99.5127
R3710 VDD.n3742 VDD.n241 99.5127
R3711 VDD.n2850 VDD.n2849 99.5127
R3712 VDD.n2846 VDD.n2845 99.5127
R3713 VDD.n2842 VDD.n2841 99.5127
R3714 VDD.n2838 VDD.n2837 99.5127
R3715 VDD.n2834 VDD.n2833 99.5127
R3716 VDD.n2830 VDD.n2829 99.5127
R3717 VDD.n2826 VDD.n2825 99.5127
R3718 VDD.n2822 VDD.n2821 99.5127
R3719 VDD.n2431 VDD.n975 99.5127
R3720 VDD.n2428 VDD.n975 99.5127
R3721 VDD.n2428 VDD.n969 99.5127
R3722 VDD.n2425 VDD.n969 99.5127
R3723 VDD.n2425 VDD.n963 99.5127
R3724 VDD.n2422 VDD.n963 99.5127
R3725 VDD.n2422 VDD.n957 99.5127
R3726 VDD.n2419 VDD.n957 99.5127
R3727 VDD.n2419 VDD.n951 99.5127
R3728 VDD.n2416 VDD.n951 99.5127
R3729 VDD.n2416 VDD.n945 99.5127
R3730 VDD.n1151 VDD.n945 99.5127
R3731 VDD.n1151 VDD.n940 99.5127
R3732 VDD.n1148 VDD.n940 99.5127
R3733 VDD.n1148 VDD.n934 99.5127
R3734 VDD.n1145 VDD.n934 99.5127
R3735 VDD.n1145 VDD.n928 99.5127
R3736 VDD.n1142 VDD.n928 99.5127
R3737 VDD.n1142 VDD.n922 99.5127
R3738 VDD.n1139 VDD.n922 99.5127
R3739 VDD.n1139 VDD.n916 99.5127
R3740 VDD.n1136 VDD.n916 99.5127
R3741 VDD.n1136 VDD.n910 99.5127
R3742 VDD.n1133 VDD.n910 99.5127
R3743 VDD.n1133 VDD.n903 99.5127
R3744 VDD.n1130 VDD.n903 99.5127
R3745 VDD.n1130 VDD.n897 99.5127
R3746 VDD.n1127 VDD.n897 99.5127
R3747 VDD.n1127 VDD.n892 99.5127
R3748 VDD.n1124 VDD.n892 99.5127
R3749 VDD.n1124 VDD.n886 99.5127
R3750 VDD.n1121 VDD.n886 99.5127
R3751 VDD.n1121 VDD.n880 99.5127
R3752 VDD.n1118 VDD.n880 99.5127
R3753 VDD.n1118 VDD.n874 99.5127
R3754 VDD.n1115 VDD.n874 99.5127
R3755 VDD.n1115 VDD.n868 99.5127
R3756 VDD.n1112 VDD.n868 99.5127
R3757 VDD.n1112 VDD.n862 99.5127
R3758 VDD.n1109 VDD.n862 99.5127
R3759 VDD.n1109 VDD.n856 99.5127
R3760 VDD.n1106 VDD.n856 99.5127
R3761 VDD.n1106 VDD.n850 99.5127
R3762 VDD.n1103 VDD.n850 99.5127
R3763 VDD.n1103 VDD.n844 99.5127
R3764 VDD.n1100 VDD.n844 99.5127
R3765 VDD.n1100 VDD.n838 99.5127
R3766 VDD.n1097 VDD.n838 99.5127
R3767 VDD.n1097 VDD.n832 99.5127
R3768 VDD.n1094 VDD.n832 99.5127
R3769 VDD.n1094 VDD.n825 99.5127
R3770 VDD.n1091 VDD.n825 99.5127
R3771 VDD.n1091 VDD.n819 99.5127
R3772 VDD.n1088 VDD.n819 99.5127
R3773 VDD.n1088 VDD.n814 99.5127
R3774 VDD.n1085 VDD.n814 99.5127
R3775 VDD.n1085 VDD.n808 99.5127
R3776 VDD.n1082 VDD.n808 99.5127
R3777 VDD.n1082 VDD.n802 99.5127
R3778 VDD.n1079 VDD.n802 99.5127
R3779 VDD.n1079 VDD.n796 99.5127
R3780 VDD.n1076 VDD.n796 99.5127
R3781 VDD.n1076 VDD.n790 99.5127
R3782 VDD.n1073 VDD.n790 99.5127
R3783 VDD.n1073 VDD.n783 99.5127
R3784 VDD.n1070 VDD.n783 99.5127
R3785 VDD.n1070 VDD.n777 99.5127
R3786 VDD.n1067 VDD.n777 99.5127
R3787 VDD.n1067 VDD.n771 99.5127
R3788 VDD.n1064 VDD.n771 99.5127
R3789 VDD.n1064 VDD.n765 99.5127
R3790 VDD.n1061 VDD.n765 99.5127
R3791 VDD.n1061 VDD.n760 99.5127
R3792 VDD.n1058 VDD.n760 99.5127
R3793 VDD.n1058 VDD.n754 99.5127
R3794 VDD.n1055 VDD.n754 99.5127
R3795 VDD.n1055 VDD.n748 99.5127
R3796 VDD.n1052 VDD.n748 99.5127
R3797 VDD.n1052 VDD.n742 99.5127
R3798 VDD.n1049 VDD.n742 99.5127
R3799 VDD.n1049 VDD.n736 99.5127
R3800 VDD.n1046 VDD.n736 99.5127
R3801 VDD.n1046 VDD.n729 99.5127
R3802 VDD.n1043 VDD.n729 99.5127
R3803 VDD.n1043 VDD.n723 99.5127
R3804 VDD.n1040 VDD.n723 99.5127
R3805 VDD.n1040 VDD.n718 99.5127
R3806 VDD.n1037 VDD.n718 99.5127
R3807 VDD.n1037 VDD.n712 99.5127
R3808 VDD.n1034 VDD.n712 99.5127
R3809 VDD.n1034 VDD.n706 99.5127
R3810 VDD.n1031 VDD.n706 99.5127
R3811 VDD.n1031 VDD.n700 99.5127
R3812 VDD.n1028 VDD.n700 99.5127
R3813 VDD.n1028 VDD.n694 99.5127
R3814 VDD.n1025 VDD.n694 99.5127
R3815 VDD.n1025 VDD.n688 99.5127
R3816 VDD.n1022 VDD.n688 99.5127
R3817 VDD.n1022 VDD.n682 99.5127
R3818 VDD.n1019 VDD.n682 99.5127
R3819 VDD.n1019 VDD.n676 99.5127
R3820 VDD.n1016 VDD.n676 99.5127
R3821 VDD.n1016 VDD.n670 99.5127
R3822 VDD.n1013 VDD.n670 99.5127
R3823 VDD.n1013 VDD.n664 99.5127
R3824 VDD.n1010 VDD.n664 99.5127
R3825 VDD.n1010 VDD.n658 99.5127
R3826 VDD.n1007 VDD.n658 99.5127
R3827 VDD.n1007 VDD.n652 99.5127
R3828 VDD.n1004 VDD.n652 99.5127
R3829 VDD.n1004 VDD.n645 99.5127
R3830 VDD.n645 VDD.n637 99.5127
R3831 VDD.n2812 VDD.n637 99.5127
R3832 VDD.n2813 VDD.n2812 99.5127
R3833 VDD.n2813 VDD.n629 99.5127
R3834 VDD.n2817 VDD.n629 99.5127
R3835 VDD.n2462 VDD.n979 99.5127
R3836 VDD.n2462 VDD.n998 99.5127
R3837 VDD.n2458 VDD.n2457 99.5127
R3838 VDD.n2454 VDD.n2453 99.5127
R3839 VDD.n2450 VDD.n2449 99.5127
R3840 VDD.n2446 VDD.n2445 99.5127
R3841 VDD.n2442 VDD.n2441 99.5127
R3842 VDD.n2438 VDD.n2437 99.5127
R3843 VDD.n2434 VDD.n987 99.5127
R3844 VDD.n2469 VDD.n977 99.5127
R3845 VDD.n2469 VDD.n967 99.5127
R3846 VDD.n2477 VDD.n967 99.5127
R3847 VDD.n2477 VDD.n965 99.5127
R3848 VDD.n2481 VDD.n965 99.5127
R3849 VDD.n2481 VDD.n955 99.5127
R3850 VDD.n2489 VDD.n955 99.5127
R3851 VDD.n2489 VDD.n953 99.5127
R3852 VDD.n2493 VDD.n953 99.5127
R3853 VDD.n2493 VDD.n944 99.5127
R3854 VDD.n2501 VDD.n944 99.5127
R3855 VDD.n2501 VDD.n942 99.5127
R3856 VDD.n2505 VDD.n942 99.5127
R3857 VDD.n2505 VDD.n932 99.5127
R3858 VDD.n2513 VDD.n932 99.5127
R3859 VDD.n2513 VDD.n930 99.5127
R3860 VDD.n2517 VDD.n930 99.5127
R3861 VDD.n2517 VDD.n920 99.5127
R3862 VDD.n2525 VDD.n920 99.5127
R3863 VDD.n2525 VDD.n918 99.5127
R3864 VDD.n2529 VDD.n918 99.5127
R3865 VDD.n2529 VDD.n908 99.5127
R3866 VDD.n2537 VDD.n908 99.5127
R3867 VDD.n2537 VDD.n906 99.5127
R3868 VDD.n2541 VDD.n906 99.5127
R3869 VDD.n2541 VDD.n896 99.5127
R3870 VDD.n2549 VDD.n896 99.5127
R3871 VDD.n2549 VDD.n894 99.5127
R3872 VDD.n2553 VDD.n894 99.5127
R3873 VDD.n2553 VDD.n884 99.5127
R3874 VDD.n2561 VDD.n884 99.5127
R3875 VDD.n2561 VDD.n882 99.5127
R3876 VDD.n2565 VDD.n882 99.5127
R3877 VDD.n2565 VDD.n872 99.5127
R3878 VDD.n2573 VDD.n872 99.5127
R3879 VDD.n2573 VDD.n870 99.5127
R3880 VDD.n2577 VDD.n870 99.5127
R3881 VDD.n2577 VDD.n860 99.5127
R3882 VDD.n2585 VDD.n860 99.5127
R3883 VDD.n2585 VDD.n858 99.5127
R3884 VDD.n2589 VDD.n858 99.5127
R3885 VDD.n2589 VDD.n848 99.5127
R3886 VDD.n2597 VDD.n848 99.5127
R3887 VDD.n2597 VDD.n846 99.5127
R3888 VDD.n2601 VDD.n846 99.5127
R3889 VDD.n2601 VDD.n836 99.5127
R3890 VDD.n2609 VDD.n836 99.5127
R3891 VDD.n2609 VDD.n834 99.5127
R3892 VDD.n2613 VDD.n834 99.5127
R3893 VDD.n2613 VDD.n823 99.5127
R3894 VDD.n2621 VDD.n823 99.5127
R3895 VDD.n2621 VDD.n821 99.5127
R3896 VDD.n2625 VDD.n821 99.5127
R3897 VDD.n2625 VDD.n812 99.5127
R3898 VDD.n2633 VDD.n812 99.5127
R3899 VDD.n2633 VDD.n810 99.5127
R3900 VDD.n2637 VDD.n810 99.5127
R3901 VDD.n2637 VDD.n800 99.5127
R3902 VDD.n2645 VDD.n800 99.5127
R3903 VDD.n2645 VDD.n798 99.5127
R3904 VDD.n2649 VDD.n798 99.5127
R3905 VDD.n2649 VDD.n788 99.5127
R3906 VDD.n2657 VDD.n788 99.5127
R3907 VDD.n2657 VDD.n786 99.5127
R3908 VDD.n2661 VDD.n786 99.5127
R3909 VDD.n2661 VDD.n776 99.5127
R3910 VDD.n2669 VDD.n776 99.5127
R3911 VDD.n2669 VDD.n774 99.5127
R3912 VDD.n2673 VDD.n774 99.5127
R3913 VDD.n2673 VDD.n764 99.5127
R3914 VDD.n2681 VDD.n764 99.5127
R3915 VDD.n2681 VDD.n762 99.5127
R3916 VDD.n2685 VDD.n762 99.5127
R3917 VDD.n2685 VDD.n752 99.5127
R3918 VDD.n2693 VDD.n752 99.5127
R3919 VDD.n2693 VDD.n750 99.5127
R3920 VDD.n2697 VDD.n750 99.5127
R3921 VDD.n2697 VDD.n740 99.5127
R3922 VDD.n2705 VDD.n740 99.5127
R3923 VDD.n2705 VDD.n738 99.5127
R3924 VDD.n2709 VDD.n738 99.5127
R3925 VDD.n2709 VDD.n727 99.5127
R3926 VDD.n2717 VDD.n727 99.5127
R3927 VDD.n2717 VDD.n725 99.5127
R3928 VDD.n2721 VDD.n725 99.5127
R3929 VDD.n2721 VDD.n716 99.5127
R3930 VDD.n2729 VDD.n716 99.5127
R3931 VDD.n2729 VDD.n714 99.5127
R3932 VDD.n2733 VDD.n714 99.5127
R3933 VDD.n2733 VDD.n704 99.5127
R3934 VDD.n2741 VDD.n704 99.5127
R3935 VDD.n2741 VDD.n702 99.5127
R3936 VDD.n2745 VDD.n702 99.5127
R3937 VDD.n2745 VDD.n692 99.5127
R3938 VDD.n2753 VDD.n692 99.5127
R3939 VDD.n2753 VDD.n690 99.5127
R3940 VDD.n2757 VDD.n690 99.5127
R3941 VDD.n2757 VDD.n680 99.5127
R3942 VDD.n2765 VDD.n680 99.5127
R3943 VDD.n2765 VDD.n678 99.5127
R3944 VDD.n2769 VDD.n678 99.5127
R3945 VDD.n2769 VDD.n668 99.5127
R3946 VDD.n2777 VDD.n668 99.5127
R3947 VDD.n2777 VDD.n666 99.5127
R3948 VDD.n2781 VDD.n666 99.5127
R3949 VDD.n2781 VDD.n656 99.5127
R3950 VDD.n2789 VDD.n656 99.5127
R3951 VDD.n2789 VDD.n654 99.5127
R3952 VDD.n2793 VDD.n654 99.5127
R3953 VDD.n2793 VDD.n643 99.5127
R3954 VDD.n2806 VDD.n643 99.5127
R3955 VDD.n2806 VDD.n641 99.5127
R3956 VDD.n2810 VDD.n641 99.5127
R3957 VDD.n2810 VDD.n631 99.5127
R3958 VDD.n2856 VDD.n631 99.5127
R3959 VDD.n2856 VDD.n632 99.5127
R3960 VDD.n3686 VDD.n3685 99.5127
R3961 VDD.n3683 VDD.n3671 99.5127
R3962 VDD.n3679 VDD.n3678 99.5127
R3963 VDD.n3676 VDD.n3674 99.5127
R3964 VDD.n3759 VDD.n3758 99.5127
R3965 VDD.n3756 VDD.n229 99.5127
R3966 VDD.n3752 VDD.n3751 99.5127
R3967 VDD.n3749 VDD.n234 99.5127
R3968 VDD.n3294 VDD.n3112 99.5127
R3969 VDD.n3294 VDD.n598 99.5127
R3970 VDD.n3291 VDD.n598 99.5127
R3971 VDD.n3291 VDD.n592 99.5127
R3972 VDD.n3288 VDD.n592 99.5127
R3973 VDD.n3288 VDD.n586 99.5127
R3974 VDD.n3285 VDD.n586 99.5127
R3975 VDD.n3285 VDD.n580 99.5127
R3976 VDD.n3282 VDD.n580 99.5127
R3977 VDD.n3282 VDD.n574 99.5127
R3978 VDD.n3279 VDD.n574 99.5127
R3979 VDD.n3279 VDD.n568 99.5127
R3980 VDD.n3276 VDD.n568 99.5127
R3981 VDD.n3276 VDD.n562 99.5127
R3982 VDD.n3273 VDD.n562 99.5127
R3983 VDD.n3273 VDD.n556 99.5127
R3984 VDD.n3270 VDD.n556 99.5127
R3985 VDD.n3270 VDD.n550 99.5127
R3986 VDD.n3267 VDD.n550 99.5127
R3987 VDD.n3267 VDD.n544 99.5127
R3988 VDD.n3264 VDD.n544 99.5127
R3989 VDD.n3264 VDD.n538 99.5127
R3990 VDD.n3261 VDD.n538 99.5127
R3991 VDD.n3261 VDD.n532 99.5127
R3992 VDD.n3258 VDD.n532 99.5127
R3993 VDD.n3258 VDD.n526 99.5127
R3994 VDD.n3255 VDD.n526 99.5127
R3995 VDD.n3255 VDD.n520 99.5127
R3996 VDD.n3252 VDD.n520 99.5127
R3997 VDD.n3252 VDD.n513 99.5127
R3998 VDD.n3249 VDD.n513 99.5127
R3999 VDD.n3249 VDD.n507 99.5127
R4000 VDD.n3246 VDD.n507 99.5127
R4001 VDD.n3246 VDD.n502 99.5127
R4002 VDD.n3243 VDD.n502 99.5127
R4003 VDD.n3243 VDD.n496 99.5127
R4004 VDD.n3240 VDD.n496 99.5127
R4005 VDD.n3240 VDD.n490 99.5127
R4006 VDD.n3237 VDD.n490 99.5127
R4007 VDD.n3237 VDD.n484 99.5127
R4008 VDD.n3234 VDD.n484 99.5127
R4009 VDD.n3234 VDD.n478 99.5127
R4010 VDD.n3231 VDD.n478 99.5127
R4011 VDD.n3231 VDD.n471 99.5127
R4012 VDD.n3228 VDD.n471 99.5127
R4013 VDD.n3228 VDD.n465 99.5127
R4014 VDD.n3225 VDD.n465 99.5127
R4015 VDD.n3225 VDD.n459 99.5127
R4016 VDD.n3222 VDD.n459 99.5127
R4017 VDD.n3222 VDD.n453 99.5127
R4018 VDD.n3219 VDD.n453 99.5127
R4019 VDD.n3219 VDD.n448 99.5127
R4020 VDD.n3216 VDD.n448 99.5127
R4021 VDD.n3216 VDD.n442 99.5127
R4022 VDD.n3213 VDD.n442 99.5127
R4023 VDD.n3213 VDD.n436 99.5127
R4024 VDD.n3210 VDD.n436 99.5127
R4025 VDD.n3210 VDD.n430 99.5127
R4026 VDD.n3207 VDD.n430 99.5127
R4027 VDD.n3207 VDD.n424 99.5127
R4028 VDD.n3204 VDD.n424 99.5127
R4029 VDD.n3204 VDD.n417 99.5127
R4030 VDD.n3201 VDD.n417 99.5127
R4031 VDD.n3201 VDD.n411 99.5127
R4032 VDD.n3198 VDD.n411 99.5127
R4033 VDD.n3198 VDD.n406 99.5127
R4034 VDD.n3195 VDD.n406 99.5127
R4035 VDD.n3195 VDD.n400 99.5127
R4036 VDD.n3192 VDD.n400 99.5127
R4037 VDD.n3192 VDD.n394 99.5127
R4038 VDD.n3189 VDD.n394 99.5127
R4039 VDD.n3189 VDD.n388 99.5127
R4040 VDD.n3186 VDD.n388 99.5127
R4041 VDD.n3186 VDD.n382 99.5127
R4042 VDD.n3183 VDD.n382 99.5127
R4043 VDD.n3183 VDD.n376 99.5127
R4044 VDD.n3180 VDD.n376 99.5127
R4045 VDD.n3180 VDD.n370 99.5127
R4046 VDD.n3177 VDD.n370 99.5127
R4047 VDD.n3177 VDD.n364 99.5127
R4048 VDD.n3174 VDD.n364 99.5127
R4049 VDD.n3174 VDD.n358 99.5127
R4050 VDD.n3171 VDD.n358 99.5127
R4051 VDD.n3171 VDD.n352 99.5127
R4052 VDD.n3168 VDD.n352 99.5127
R4053 VDD.n3168 VDD.n346 99.5127
R4054 VDD.n3165 VDD.n346 99.5127
R4055 VDD.n3165 VDD.n339 99.5127
R4056 VDD.n3162 VDD.n339 99.5127
R4057 VDD.n3162 VDD.n333 99.5127
R4058 VDD.n3159 VDD.n333 99.5127
R4059 VDD.n3159 VDD.n328 99.5127
R4060 VDD.n3156 VDD.n328 99.5127
R4061 VDD.n3156 VDD.n322 99.5127
R4062 VDD.n3153 VDD.n322 99.5127
R4063 VDD.n3153 VDD.n316 99.5127
R4064 VDD.n3150 VDD.n316 99.5127
R4065 VDD.n3150 VDD.n310 99.5127
R4066 VDD.n3147 VDD.n310 99.5127
R4067 VDD.n3147 VDD.n304 99.5127
R4068 VDD.n3144 VDD.n304 99.5127
R4069 VDD.n3144 VDD.n298 99.5127
R4070 VDD.n3141 VDD.n298 99.5127
R4071 VDD.n3141 VDD.n291 99.5127
R4072 VDD.n3138 VDD.n291 99.5127
R4073 VDD.n3138 VDD.n285 99.5127
R4074 VDD.n3135 VDD.n285 99.5127
R4075 VDD.n3135 VDD.n280 99.5127
R4076 VDD.n3132 VDD.n280 99.5127
R4077 VDD.n3132 VDD.n274 99.5127
R4078 VDD.n3129 VDD.n274 99.5127
R4079 VDD.n3129 VDD.n267 99.5127
R4080 VDD.n3126 VDD.n267 99.5127
R4081 VDD.n3126 VDD.n260 99.5127
R4082 VDD.n260 VDD.n237 99.5127
R4083 VDD.n3744 VDD.n237 99.5127
R4084 VDD.n3330 VDD.n3328 99.5127
R4085 VDD.n3326 VDD.n3115 99.5127
R4086 VDD.n3322 VDD.n3320 99.5127
R4087 VDD.n3318 VDD.n3117 99.5127
R4088 VDD.n3314 VDD.n3312 99.5127
R4089 VDD.n3310 VDD.n3119 99.5127
R4090 VDD.n3306 VDD.n3304 99.5127
R4091 VDD.n3302 VDD.n3123 99.5127
R4092 VDD.n3334 VDD.n595 99.5127
R4093 VDD.n3342 VDD.n595 99.5127
R4094 VDD.n3342 VDD.n593 99.5127
R4095 VDD.n3346 VDD.n593 99.5127
R4096 VDD.n3346 VDD.n583 99.5127
R4097 VDD.n3354 VDD.n583 99.5127
R4098 VDD.n3354 VDD.n581 99.5127
R4099 VDD.n3358 VDD.n581 99.5127
R4100 VDD.n3358 VDD.n571 99.5127
R4101 VDD.n3366 VDD.n571 99.5127
R4102 VDD.n3366 VDD.n569 99.5127
R4103 VDD.n3370 VDD.n569 99.5127
R4104 VDD.n3370 VDD.n559 99.5127
R4105 VDD.n3378 VDD.n559 99.5127
R4106 VDD.n3378 VDD.n557 99.5127
R4107 VDD.n3382 VDD.n557 99.5127
R4108 VDD.n3382 VDD.n547 99.5127
R4109 VDD.n3390 VDD.n547 99.5127
R4110 VDD.n3390 VDD.n545 99.5127
R4111 VDD.n3394 VDD.n545 99.5127
R4112 VDD.n3394 VDD.n535 99.5127
R4113 VDD.n3402 VDD.n535 99.5127
R4114 VDD.n3402 VDD.n533 99.5127
R4115 VDD.n3406 VDD.n533 99.5127
R4116 VDD.n3406 VDD.n523 99.5127
R4117 VDD.n3414 VDD.n523 99.5127
R4118 VDD.n3414 VDD.n521 99.5127
R4119 VDD.n3418 VDD.n521 99.5127
R4120 VDD.n3418 VDD.n510 99.5127
R4121 VDD.n3426 VDD.n510 99.5127
R4122 VDD.n3426 VDD.n508 99.5127
R4123 VDD.n3430 VDD.n508 99.5127
R4124 VDD.n3430 VDD.n499 99.5127
R4125 VDD.n3438 VDD.n499 99.5127
R4126 VDD.n3438 VDD.n497 99.5127
R4127 VDD.n3442 VDD.n497 99.5127
R4128 VDD.n3442 VDD.n487 99.5127
R4129 VDD.n3450 VDD.n487 99.5127
R4130 VDD.n3450 VDD.n485 99.5127
R4131 VDD.n3454 VDD.n485 99.5127
R4132 VDD.n3454 VDD.n475 99.5127
R4133 VDD.n3462 VDD.n475 99.5127
R4134 VDD.n3462 VDD.n473 99.5127
R4135 VDD.n3466 VDD.n473 99.5127
R4136 VDD.n3466 VDD.n463 99.5127
R4137 VDD.n3474 VDD.n463 99.5127
R4138 VDD.n3474 VDD.n461 99.5127
R4139 VDD.n3478 VDD.n461 99.5127
R4140 VDD.n3478 VDD.n451 99.5127
R4141 VDD.n3486 VDD.n451 99.5127
R4142 VDD.n3486 VDD.n449 99.5127
R4143 VDD.n3490 VDD.n449 99.5127
R4144 VDD.n3490 VDD.n439 99.5127
R4145 VDD.n3498 VDD.n439 99.5127
R4146 VDD.n3498 VDD.n437 99.5127
R4147 VDD.n3502 VDD.n437 99.5127
R4148 VDD.n3502 VDD.n427 99.5127
R4149 VDD.n3510 VDD.n427 99.5127
R4150 VDD.n3510 VDD.n425 99.5127
R4151 VDD.n3514 VDD.n425 99.5127
R4152 VDD.n3514 VDD.n414 99.5127
R4153 VDD.n3522 VDD.n414 99.5127
R4154 VDD.n3522 VDD.n412 99.5127
R4155 VDD.n3526 VDD.n412 99.5127
R4156 VDD.n3526 VDD.n403 99.5127
R4157 VDD.n3534 VDD.n403 99.5127
R4158 VDD.n3534 VDD.n401 99.5127
R4159 VDD.n3538 VDD.n401 99.5127
R4160 VDD.n3538 VDD.n391 99.5127
R4161 VDD.n3546 VDD.n391 99.5127
R4162 VDD.n3546 VDD.n389 99.5127
R4163 VDD.n3550 VDD.n389 99.5127
R4164 VDD.n3550 VDD.n379 99.5127
R4165 VDD.n3558 VDD.n379 99.5127
R4166 VDD.n3558 VDD.n377 99.5127
R4167 VDD.n3562 VDD.n377 99.5127
R4168 VDD.n3562 VDD.n367 99.5127
R4169 VDD.n3570 VDD.n367 99.5127
R4170 VDD.n3570 VDD.n365 99.5127
R4171 VDD.n3574 VDD.n365 99.5127
R4172 VDD.n3574 VDD.n355 99.5127
R4173 VDD.n3582 VDD.n355 99.5127
R4174 VDD.n3582 VDD.n353 99.5127
R4175 VDD.n3586 VDD.n353 99.5127
R4176 VDD.n3586 VDD.n343 99.5127
R4177 VDD.n3594 VDD.n343 99.5127
R4178 VDD.n3594 VDD.n341 99.5127
R4179 VDD.n3598 VDD.n341 99.5127
R4180 VDD.n3598 VDD.n331 99.5127
R4181 VDD.n3606 VDD.n331 99.5127
R4182 VDD.n3606 VDD.n329 99.5127
R4183 VDD.n3610 VDD.n329 99.5127
R4184 VDD.n3610 VDD.n319 99.5127
R4185 VDD.n3618 VDD.n319 99.5127
R4186 VDD.n3618 VDD.n317 99.5127
R4187 VDD.n3622 VDD.n317 99.5127
R4188 VDD.n3622 VDD.n307 99.5127
R4189 VDD.n3630 VDD.n307 99.5127
R4190 VDD.n3630 VDD.n305 99.5127
R4191 VDD.n3634 VDD.n305 99.5127
R4192 VDD.n3634 VDD.n295 99.5127
R4193 VDD.n3642 VDD.n295 99.5127
R4194 VDD.n3642 VDD.n293 99.5127
R4195 VDD.n3646 VDD.n293 99.5127
R4196 VDD.n3646 VDD.n283 99.5127
R4197 VDD.n3654 VDD.n283 99.5127
R4198 VDD.n3654 VDD.n281 99.5127
R4199 VDD.n3658 VDD.n281 99.5127
R4200 VDD.n3658 VDD.n271 99.5127
R4201 VDD.n3666 VDD.n271 99.5127
R4202 VDD.n3666 VDD.n268 99.5127
R4203 VDD.n3696 VDD.n268 99.5127
R4204 VDD.n3696 VDD.n269 99.5127
R4205 VDD.n269 VDD.n261 99.5127
R4206 VDD.n3691 VDD.n261 99.5127
R4207 VDD.n3691 VDD.n240 99.5127
R4208 VDD.n2894 VDD.n622 99.5127
R4209 VDD.n2890 VDD.n2889 99.5127
R4210 VDD.n2886 VDD.n2885 99.5127
R4211 VDD.n2882 VDD.n2881 99.5127
R4212 VDD.n2878 VDD.n2877 99.5127
R4213 VDD.n2874 VDD.n2873 99.5127
R4214 VDD.n2870 VDD.n2869 99.5127
R4215 VDD.n2866 VDD.n2865 99.5127
R4216 VDD.n2862 VDD.n620 99.5127
R4217 VDD.n2243 VDD.n976 99.5127
R4218 VDD.n2246 VDD.n976 99.5127
R4219 VDD.n2246 VDD.n970 99.5127
R4220 VDD.n2249 VDD.n970 99.5127
R4221 VDD.n2249 VDD.n964 99.5127
R4222 VDD.n2252 VDD.n964 99.5127
R4223 VDD.n2252 VDD.n958 99.5127
R4224 VDD.n2255 VDD.n958 99.5127
R4225 VDD.n2255 VDD.n952 99.5127
R4226 VDD.n2414 VDD.n952 99.5127
R4227 VDD.n2414 VDD.n946 99.5127
R4228 VDD.n2410 VDD.n946 99.5127
R4229 VDD.n2410 VDD.n941 99.5127
R4230 VDD.n2407 VDD.n941 99.5127
R4231 VDD.n2407 VDD.n935 99.5127
R4232 VDD.n2404 VDD.n935 99.5127
R4233 VDD.n2404 VDD.n929 99.5127
R4234 VDD.n2401 VDD.n929 99.5127
R4235 VDD.n2401 VDD.n923 99.5127
R4236 VDD.n2398 VDD.n923 99.5127
R4237 VDD.n2398 VDD.n917 99.5127
R4238 VDD.n2395 VDD.n917 99.5127
R4239 VDD.n2395 VDD.n911 99.5127
R4240 VDD.n2392 VDD.n911 99.5127
R4241 VDD.n2392 VDD.n904 99.5127
R4242 VDD.n2389 VDD.n904 99.5127
R4243 VDD.n2389 VDD.n898 99.5127
R4244 VDD.n2386 VDD.n898 99.5127
R4245 VDD.n2386 VDD.n893 99.5127
R4246 VDD.n2383 VDD.n893 99.5127
R4247 VDD.n2383 VDD.n887 99.5127
R4248 VDD.n2380 VDD.n887 99.5127
R4249 VDD.n2380 VDD.n881 99.5127
R4250 VDD.n2377 VDD.n881 99.5127
R4251 VDD.n2377 VDD.n875 99.5127
R4252 VDD.n2374 VDD.n875 99.5127
R4253 VDD.n2374 VDD.n869 99.5127
R4254 VDD.n2371 VDD.n869 99.5127
R4255 VDD.n2371 VDD.n863 99.5127
R4256 VDD.n2368 VDD.n863 99.5127
R4257 VDD.n2368 VDD.n857 99.5127
R4258 VDD.n2365 VDD.n857 99.5127
R4259 VDD.n2365 VDD.n851 99.5127
R4260 VDD.n2362 VDD.n851 99.5127
R4261 VDD.n2362 VDD.n845 99.5127
R4262 VDD.n2359 VDD.n845 99.5127
R4263 VDD.n2359 VDD.n839 99.5127
R4264 VDD.n2356 VDD.n839 99.5127
R4265 VDD.n2356 VDD.n833 99.5127
R4266 VDD.n2353 VDD.n833 99.5127
R4267 VDD.n2353 VDD.n826 99.5127
R4268 VDD.n2350 VDD.n826 99.5127
R4269 VDD.n2350 VDD.n820 99.5127
R4270 VDD.n2347 VDD.n820 99.5127
R4271 VDD.n2347 VDD.n815 99.5127
R4272 VDD.n2344 VDD.n815 99.5127
R4273 VDD.n2344 VDD.n809 99.5127
R4274 VDD.n2341 VDD.n809 99.5127
R4275 VDD.n2341 VDD.n803 99.5127
R4276 VDD.n2338 VDD.n803 99.5127
R4277 VDD.n2338 VDD.n797 99.5127
R4278 VDD.n2335 VDD.n797 99.5127
R4279 VDD.n2335 VDD.n791 99.5127
R4280 VDD.n2332 VDD.n791 99.5127
R4281 VDD.n2332 VDD.n784 99.5127
R4282 VDD.n2329 VDD.n784 99.5127
R4283 VDD.n2329 VDD.n778 99.5127
R4284 VDD.n2326 VDD.n778 99.5127
R4285 VDD.n2326 VDD.n772 99.5127
R4286 VDD.n2323 VDD.n772 99.5127
R4287 VDD.n2323 VDD.n766 99.5127
R4288 VDD.n2320 VDD.n766 99.5127
R4289 VDD.n2320 VDD.n761 99.5127
R4290 VDD.n2317 VDD.n761 99.5127
R4291 VDD.n2317 VDD.n755 99.5127
R4292 VDD.n2314 VDD.n755 99.5127
R4293 VDD.n2314 VDD.n749 99.5127
R4294 VDD.n2311 VDD.n749 99.5127
R4295 VDD.n2311 VDD.n743 99.5127
R4296 VDD.n2308 VDD.n743 99.5127
R4297 VDD.n2308 VDD.n737 99.5127
R4298 VDD.n2305 VDD.n737 99.5127
R4299 VDD.n2305 VDD.n730 99.5127
R4300 VDD.n2302 VDD.n730 99.5127
R4301 VDD.n2302 VDD.n724 99.5127
R4302 VDD.n2299 VDD.n724 99.5127
R4303 VDD.n2299 VDD.n719 99.5127
R4304 VDD.n2296 VDD.n719 99.5127
R4305 VDD.n2296 VDD.n713 99.5127
R4306 VDD.n2293 VDD.n713 99.5127
R4307 VDD.n2293 VDD.n707 99.5127
R4308 VDD.n2290 VDD.n707 99.5127
R4309 VDD.n2290 VDD.n701 99.5127
R4310 VDD.n2287 VDD.n701 99.5127
R4311 VDD.n2287 VDD.n695 99.5127
R4312 VDD.n2284 VDD.n695 99.5127
R4313 VDD.n2284 VDD.n689 99.5127
R4314 VDD.n2281 VDD.n689 99.5127
R4315 VDD.n2281 VDD.n683 99.5127
R4316 VDD.n2278 VDD.n683 99.5127
R4317 VDD.n2278 VDD.n677 99.5127
R4318 VDD.n2275 VDD.n677 99.5127
R4319 VDD.n2275 VDD.n671 99.5127
R4320 VDD.n2272 VDD.n671 99.5127
R4321 VDD.n2272 VDD.n665 99.5127
R4322 VDD.n2269 VDD.n665 99.5127
R4323 VDD.n2269 VDD.n659 99.5127
R4324 VDD.n2266 VDD.n659 99.5127
R4325 VDD.n2266 VDD.n653 99.5127
R4326 VDD.n2263 VDD.n653 99.5127
R4327 VDD.n2263 VDD.n646 99.5127
R4328 VDD.n2260 VDD.n646 99.5127
R4329 VDD.n2260 VDD.n639 99.5127
R4330 VDD.n639 VDD.n627 99.5127
R4331 VDD.n2858 VDD.n627 99.5127
R4332 VDD.n2859 VDD.n2858 99.5127
R4333 VDD.n2210 VDD.n997 99.5127
R4334 VDD.n2214 VDD.n2213 99.5127
R4335 VDD.n2218 VDD.n2217 99.5127
R4336 VDD.n2222 VDD.n2221 99.5127
R4337 VDD.n2226 VDD.n2225 99.5127
R4338 VDD.n2230 VDD.n2229 99.5127
R4339 VDD.n2234 VDD.n2233 99.5127
R4340 VDD.n2238 VDD.n2237 99.5127
R4341 VDD.n2240 VDD.n996 99.5127
R4342 VDD.n2471 VDD.n973 99.5127
R4343 VDD.n2471 VDD.n971 99.5127
R4344 VDD.n2475 VDD.n971 99.5127
R4345 VDD.n2475 VDD.n961 99.5127
R4346 VDD.n2483 VDD.n961 99.5127
R4347 VDD.n2483 VDD.n959 99.5127
R4348 VDD.n2487 VDD.n959 99.5127
R4349 VDD.n2487 VDD.n949 99.5127
R4350 VDD.n2495 VDD.n949 99.5127
R4351 VDD.n2495 VDD.n947 99.5127
R4352 VDD.n2499 VDD.n947 99.5127
R4353 VDD.n2499 VDD.n938 99.5127
R4354 VDD.n2507 VDD.n938 99.5127
R4355 VDD.n2507 VDD.n936 99.5127
R4356 VDD.n2511 VDD.n936 99.5127
R4357 VDD.n2511 VDD.n926 99.5127
R4358 VDD.n2519 VDD.n926 99.5127
R4359 VDD.n2519 VDD.n924 99.5127
R4360 VDD.n2523 VDD.n924 99.5127
R4361 VDD.n2523 VDD.n914 99.5127
R4362 VDD.n2531 VDD.n914 99.5127
R4363 VDD.n2531 VDD.n912 99.5127
R4364 VDD.n2535 VDD.n912 99.5127
R4365 VDD.n2535 VDD.n901 99.5127
R4366 VDD.n2543 VDD.n901 99.5127
R4367 VDD.n2543 VDD.n899 99.5127
R4368 VDD.n2547 VDD.n899 99.5127
R4369 VDD.n2547 VDD.n890 99.5127
R4370 VDD.n2555 VDD.n890 99.5127
R4371 VDD.n2555 VDD.n888 99.5127
R4372 VDD.n2559 VDD.n888 99.5127
R4373 VDD.n2559 VDD.n878 99.5127
R4374 VDD.n2567 VDD.n878 99.5127
R4375 VDD.n2567 VDD.n876 99.5127
R4376 VDD.n2571 VDD.n876 99.5127
R4377 VDD.n2571 VDD.n866 99.5127
R4378 VDD.n2579 VDD.n866 99.5127
R4379 VDD.n2579 VDD.n864 99.5127
R4380 VDD.n2583 VDD.n864 99.5127
R4381 VDD.n2583 VDD.n854 99.5127
R4382 VDD.n2591 VDD.n854 99.5127
R4383 VDD.n2591 VDD.n852 99.5127
R4384 VDD.n2595 VDD.n852 99.5127
R4385 VDD.n2595 VDD.n842 99.5127
R4386 VDD.n2603 VDD.n842 99.5127
R4387 VDD.n2603 VDD.n840 99.5127
R4388 VDD.n2607 VDD.n840 99.5127
R4389 VDD.n2607 VDD.n830 99.5127
R4390 VDD.n2615 VDD.n830 99.5127
R4391 VDD.n2615 VDD.n828 99.5127
R4392 VDD.n2619 VDD.n828 99.5127
R4393 VDD.n2619 VDD.n818 99.5127
R4394 VDD.n2627 VDD.n818 99.5127
R4395 VDD.n2627 VDD.n816 99.5127
R4396 VDD.n2631 VDD.n816 99.5127
R4397 VDD.n2631 VDD.n806 99.5127
R4398 VDD.n2639 VDD.n806 99.5127
R4399 VDD.n2639 VDD.n804 99.5127
R4400 VDD.n2643 VDD.n804 99.5127
R4401 VDD.n2643 VDD.n794 99.5127
R4402 VDD.n2651 VDD.n794 99.5127
R4403 VDD.n2651 VDD.n792 99.5127
R4404 VDD.n2655 VDD.n792 99.5127
R4405 VDD.n2655 VDD.n781 99.5127
R4406 VDD.n2663 VDD.n781 99.5127
R4407 VDD.n2663 VDD.n779 99.5127
R4408 VDD.n2667 VDD.n779 99.5127
R4409 VDD.n2667 VDD.n769 99.5127
R4410 VDD.n2675 VDD.n769 99.5127
R4411 VDD.n2675 VDD.n767 99.5127
R4412 VDD.n2679 VDD.n767 99.5127
R4413 VDD.n2679 VDD.n758 99.5127
R4414 VDD.n2687 VDD.n758 99.5127
R4415 VDD.n2687 VDD.n756 99.5127
R4416 VDD.n2691 VDD.n756 99.5127
R4417 VDD.n2691 VDD.n746 99.5127
R4418 VDD.n2699 VDD.n746 99.5127
R4419 VDD.n2699 VDD.n744 99.5127
R4420 VDD.n2703 VDD.n744 99.5127
R4421 VDD.n2703 VDD.n734 99.5127
R4422 VDD.n2711 VDD.n734 99.5127
R4423 VDD.n2711 VDD.n732 99.5127
R4424 VDD.n2715 VDD.n732 99.5127
R4425 VDD.n2715 VDD.n722 99.5127
R4426 VDD.n2723 VDD.n722 99.5127
R4427 VDD.n2723 VDD.n720 99.5127
R4428 VDD.n2727 VDD.n720 99.5127
R4429 VDD.n2727 VDD.n710 99.5127
R4430 VDD.n2735 VDD.n710 99.5127
R4431 VDD.n2735 VDD.n708 99.5127
R4432 VDD.n2739 VDD.n708 99.5127
R4433 VDD.n2739 VDD.n698 99.5127
R4434 VDD.n2747 VDD.n698 99.5127
R4435 VDD.n2747 VDD.n696 99.5127
R4436 VDD.n2751 VDD.n696 99.5127
R4437 VDD.n2751 VDD.n686 99.5127
R4438 VDD.n2759 VDD.n686 99.5127
R4439 VDD.n2759 VDD.n684 99.5127
R4440 VDD.n2763 VDD.n684 99.5127
R4441 VDD.n2763 VDD.n674 99.5127
R4442 VDD.n2771 VDD.n674 99.5127
R4443 VDD.n2771 VDD.n672 99.5127
R4444 VDD.n2775 VDD.n672 99.5127
R4445 VDD.n2775 VDD.n662 99.5127
R4446 VDD.n2783 VDD.n662 99.5127
R4447 VDD.n2783 VDD.n660 99.5127
R4448 VDD.n2787 VDD.n660 99.5127
R4449 VDD.n2787 VDD.n650 99.5127
R4450 VDD.n2795 VDD.n650 99.5127
R4451 VDD.n2795 VDD.n647 99.5127
R4452 VDD.n2804 VDD.n647 99.5127
R4453 VDD.n2804 VDD.n648 99.5127
R4454 VDD.n648 VDD.n640 99.5127
R4455 VDD.n2799 VDD.n640 99.5127
R4456 VDD.n2799 VDD.n630 99.5127
R4457 VDD.n630 VDD.n621 99.5127
R4458 VDD.n1491 VDD.t35 97.7139
R4459 VDD.n1557 VDD.t89 97.7139
R4460 VDD.n1587 VDD.t98 97.7139
R4461 VDD.n1642 VDD.t57 97.7139
R4462 VDD.n1420 VDD.t73 97.7139
R4463 VDD.n1976 VDD.t77 97.7139
R4464 VDD.n2036 VDD.t44 97.7139
R4465 VDD.n1190 VDD.t55 97.7139
R4466 VDD.n1165 VDD.t61 97.7139
R4467 VDD.n2005 VDD.t64 97.7139
R4468 VDD.n207 VDD.t51 97.7139
R4469 VDD.n3796 VDD.t101 97.7139
R4470 VDD.n4257 VDD.t93 97.7139
R4471 VDD.n4289 VDD.t105 97.7139
R4472 VDD.n4226 VDD.t108 97.7139
R4473 VDD.n4509 VDD.t40 97.7139
R4474 VDD.n151 VDD.t86 97.7139
R4475 VDD.n4321 VDD.t96 94.5139
R4476 VDD.n178 VDD.t66 94.5139
R4477 VDD.n3833 VDD.t113 94.5139
R4478 VDD.n1831 VDD.t18 92.3973
R4479 VDD.n1828 VDD.t166 92.3973
R4480 VDD.n1825 VDD.t8 92.3973
R4481 VDD.n1822 VDD.t3 92.3973
R4482 VDD.n1820 VDD.t21 92.3973
R4483 VDD.n1491 VDD.n1490 90.9581
R4484 VDD.n1557 VDD.n1556 90.9581
R4485 VDD.n1587 VDD.n1586 90.9581
R4486 VDD.n1642 VDD.n1641 90.9581
R4487 VDD.n1420 VDD.n1419 90.9581
R4488 VDD.n1976 VDD.n1975 90.9581
R4489 VDD.n2036 VDD.n2035 90.9581
R4490 VDD.n1190 VDD.n1189 90.9581
R4491 VDD.n1165 VDD.n1164 90.9581
R4492 VDD.n2005 VDD.n2004 90.9581
R4493 VDD.n207 VDD.n206 90.9581
R4494 VDD.n3796 VDD.n3795 90.9581
R4495 VDD.n4257 VDD.n4256 90.9581
R4496 VDD.n4289 VDD.n4288 90.9581
R4497 VDD.n4226 VDD.n4225 90.9581
R4498 VDD.n4509 VDD.n4508 90.9581
R4499 VDD.n151 VDD.n150 90.9581
R4500 VDD.n28 VDD.t163 90.86
R4501 VDD.n25 VDD.t19 90.86
R4502 VDD.n22 VDD.t169 90.86
R4503 VDD.n19 VDD.t14 90.86
R4504 VDD.n17 VDD.t10 90.86
R4505 VDD.n28 VDD.n27 79.5496
R4506 VDD.n25 VDD.n24 79.5496
R4507 VDD.n22 VDD.n21 79.5496
R4508 VDD.n19 VDD.n18 79.5496
R4509 VDD.n17 VDD.n16 79.5496
R4510 VDD.n1831 VDD.n1830 78.0122
R4511 VDD.n1828 VDD.n1827 78.0122
R4512 VDD.n1825 VDD.n1824 78.0122
R4513 VDD.n1822 VDD.n1821 78.0122
R4514 VDD.n1820 VDD.n1819 78.0122
R4515 VDD.n2896 VDD.n2895 77.1137
R4516 VDD.n3329 VDD.n2896 72.8958
R4517 VDD.n3327 VDD.n2896 72.8958
R4518 VDD.n3321 VDD.n2896 72.8958
R4519 VDD.n3319 VDD.n2896 72.8958
R4520 VDD.n3313 VDD.n2896 72.8958
R4521 VDD.n3311 VDD.n2896 72.8958
R4522 VDD.n3305 VDD.n2896 72.8958
R4523 VDD.n3303 VDD.n2896 72.8958
R4524 VDD.n3297 VDD.n2896 72.8958
R4525 VDD.n236 VDD.n228 72.8958
R4526 VDD.n3750 VDD.n228 72.8958
R4527 VDD.n233 VDD.n228 72.8958
R4528 VDD.n3757 VDD.n228 72.8958
R4529 VDD.n228 VDD.n227 72.8958
R4530 VDD.n3677 VDD.n228 72.8958
R4531 VDD.n3673 VDD.n228 72.8958
R4532 VDD.n3684 VDD.n228 72.8958
R4533 VDD.n3687 VDD.n228 72.8958
R4534 VDD.n2464 VDD.n2463 72.8958
R4535 VDD.n2463 VDD.n980 72.8958
R4536 VDD.n2463 VDD.n981 72.8958
R4537 VDD.n2463 VDD.n982 72.8958
R4538 VDD.n2463 VDD.n983 72.8958
R4539 VDD.n2463 VDD.n984 72.8958
R4540 VDD.n2463 VDD.n985 72.8958
R4541 VDD.n2463 VDD.n986 72.8958
R4542 VDD.n2895 VDD.n611 72.8958
R4543 VDD.n2895 VDD.n610 72.8958
R4544 VDD.n2895 VDD.n609 72.8958
R4545 VDD.n2895 VDD.n608 72.8958
R4546 VDD.n2895 VDD.n607 72.8958
R4547 VDD.n2895 VDD.n606 72.8958
R4548 VDD.n2895 VDD.n605 72.8958
R4549 VDD.n2895 VDD.n604 72.8958
R4550 VDD.n2895 VDD.n603 72.8958
R4551 VDD.n2910 VDD.n2896 72.8958
R4552 VDD.n2913 VDD.n2896 72.8958
R4553 VDD.n2919 VDD.n2896 72.8958
R4554 VDD.n2921 VDD.n2896 72.8958
R4555 VDD.n2927 VDD.n2896 72.8958
R4556 VDD.n2929 VDD.n2896 72.8958
R4557 VDD.n2935 VDD.n2896 72.8958
R4558 VDD.n2938 VDD.n2896 72.8958
R4559 VDD.n3710 VDD.n228 72.8958
R4560 VDD.n256 VDD.n228 72.8958
R4561 VDD.n3717 VDD.n228 72.8958
R4562 VDD.n251 VDD.n228 72.8958
R4563 VDD.n3724 VDD.n228 72.8958
R4564 VDD.n3729 VDD.n228 72.8958
R4565 VDD.n248 VDD.n228 72.8958
R4566 VDD.n3736 VDD.n228 72.8958
R4567 VDD.n245 VDD.n228 72.8958
R4568 VDD.n2895 VDD.n619 72.8958
R4569 VDD.n2895 VDD.n618 72.8958
R4570 VDD.n2895 VDD.n617 72.8958
R4571 VDD.n2895 VDD.n616 72.8958
R4572 VDD.n2895 VDD.n615 72.8958
R4573 VDD.n2895 VDD.n614 72.8958
R4574 VDD.n2895 VDD.n613 72.8958
R4575 VDD.n2895 VDD.n612 72.8958
R4576 VDD.n2463 VDD.n988 72.8958
R4577 VDD.n2463 VDD.n989 72.8958
R4578 VDD.n2463 VDD.n990 72.8958
R4579 VDD.n2463 VDD.n991 72.8958
R4580 VDD.n2463 VDD.n992 72.8958
R4581 VDD.n2463 VDD.n993 72.8958
R4582 VDD.n2463 VDD.n994 72.8958
R4583 VDD.n2463 VDD.n995 72.8958
R4584 VDD.n1392 VDD.n1389 66.2847
R4585 VDD.n1398 VDD.n1389 66.2847
R4586 VDD.n1401 VDD.n1389 66.2847
R4587 VDD.n1406 VDD.n1389 66.2847
R4588 VDD.n1409 VDD.n1389 66.2847
R4589 VDD.n1414 VDD.n1389 66.2847
R4590 VDD.n1417 VDD.n1389 66.2847
R4591 VDD.n1424 VDD.n1389 66.2847
R4592 VDD.n1429 VDD.n1389 66.2847
R4593 VDD.n1432 VDD.n1389 66.2847
R4594 VDD.n1437 VDD.n1389 66.2847
R4595 VDD.n1440 VDD.n1389 66.2847
R4596 VDD.n1445 VDD.n1389 66.2847
R4597 VDD.n1448 VDD.n1389 66.2847
R4598 VDD.n1453 VDD.n1389 66.2847
R4599 VDD.n1456 VDD.n1389 66.2847
R4600 VDD.n1461 VDD.n1389 66.2847
R4601 VDD.n1464 VDD.n1389 66.2847
R4602 VDD.n1469 VDD.n1389 66.2847
R4603 VDD.n1472 VDD.n1389 66.2847
R4604 VDD.n1477 VDD.n1389 66.2847
R4605 VDD.n1480 VDD.n1389 66.2847
R4606 VDD.n1485 VDD.n1389 66.2847
R4607 VDD.n1488 VDD.n1389 66.2847
R4608 VDD.n1613 VDD.n1389 66.2847
R4609 VDD.n1494 VDD.n1389 66.2847
R4610 VDD.n1500 VDD.n1389 66.2847
R4611 VDD.n1505 VDD.n1389 66.2847
R4612 VDD.n1508 VDD.n1389 66.2847
R4613 VDD.n1513 VDD.n1389 66.2847
R4614 VDD.n1516 VDD.n1389 66.2847
R4615 VDD.n1522 VDD.n1389 66.2847
R4616 VDD.n1584 VDD.n1389 66.2847
R4617 VDD.n1524 VDD.n1389 66.2847
R4618 VDD.n1529 VDD.n1389 66.2847
R4619 VDD.n1534 VDD.n1389 66.2847
R4620 VDD.n1537 VDD.n1389 66.2847
R4621 VDD.n1542 VDD.n1389 66.2847
R4622 VDD.n1545 VDD.n1389 66.2847
R4623 VDD.n1550 VDD.n1389 66.2847
R4624 VDD.n1554 VDD.n1389 66.2847
R4625 VDD.n2173 VDD.n1206 66.2847
R4626 VDD.n1206 VDD.n1205 66.2847
R4627 VDD.n1206 VDD.n1204 66.2847
R4628 VDD.n1206 VDD.n1203 66.2847
R4629 VDD.n1206 VDD.n1201 66.2847
R4630 VDD.n1206 VDD.n1200 66.2847
R4631 VDD.n1206 VDD.n1198 66.2847
R4632 VDD.n1206 VDD.n1197 66.2847
R4633 VDD.n1206 VDD.n1195 66.2847
R4634 VDD.n1206 VDD.n1194 66.2847
R4635 VDD.n1206 VDD.n1192 66.2847
R4636 VDD.n2053 VDD.n1206 66.2847
R4637 VDD.n2058 VDD.n1206 66.2847
R4638 VDD.n2063 VDD.n1206 66.2847
R4639 VDD.n2051 VDD.n1206 66.2847
R4640 VDD.n2070 VDD.n1206 66.2847
R4641 VDD.n2044 VDD.n1206 66.2847
R4642 VDD.n2079 VDD.n1206 66.2847
R4643 VDD.n2038 VDD.n1206 66.2847
R4644 VDD.n2086 VDD.n1206 66.2847
R4645 VDD.n2029 VDD.n1206 66.2847
R4646 VDD.n2093 VDD.n1206 66.2847
R4647 VDD.n2022 VDD.n1206 66.2847
R4648 VDD.n2100 VDD.n1206 66.2847
R4649 VDD.n2015 VDD.n1206 66.2847
R4650 VDD.n2107 VDD.n1206 66.2847
R4651 VDD.n2007 VDD.n1206 66.2847
R4652 VDD.n2114 VDD.n1206 66.2847
R4653 VDD.n2117 VDD.n1206 66.2847
R4654 VDD.n1996 VDD.n1206 66.2847
R4655 VDD.n2126 VDD.n1206 66.2847
R4656 VDD.n1990 VDD.n1206 66.2847
R4657 VDD.n2133 VDD.n1206 66.2847
R4658 VDD.n1983 VDD.n1206 66.2847
R4659 VDD.n2140 VDD.n1206 66.2847
R4660 VDD.n1973 VDD.n1206 66.2847
R4661 VDD.n2147 VDD.n1206 66.2847
R4662 VDD.n1966 VDD.n1206 66.2847
R4663 VDD.n2154 VDD.n1206 66.2847
R4664 VDD.n1959 VDD.n1206 66.2847
R4665 VDD.n2161 VDD.n1206 66.2847
R4666 VDD.n1952 VDD.n1206 66.2847
R4667 VDD.n3961 VDD.n126 66.2847
R4668 VDD.n130 VDD.n126 66.2847
R4669 VDD.n3954 VDD.n126 66.2847
R4670 VDD.n3948 VDD.n126 66.2847
R4671 VDD.n3946 VDD.n126 66.2847
R4672 VDD.n3940 VDD.n126 66.2847
R4673 VDD.n3938 VDD.n126 66.2847
R4674 VDD.n3931 VDD.n126 66.2847
R4675 VDD.n3929 VDD.n126 66.2847
R4676 VDD.n3923 VDD.n126 66.2847
R4677 VDD.n3921 VDD.n126 66.2847
R4678 VDD.n166 VDD.n126 66.2847
R4679 VDD.n3911 VDD.n126 66.2847
R4680 VDD.n3909 VDD.n126 66.2847
R4681 VDD.n3903 VDD.n126 66.2847
R4682 VDD.n3901 VDD.n126 66.2847
R4683 VDD.n3895 VDD.n126 66.2847
R4684 VDD.n3893 VDD.n126 66.2847
R4685 VDD.n3887 VDD.n126 66.2847
R4686 VDD.n3885 VDD.n126 66.2847
R4687 VDD.n3879 VDD.n126 66.2847
R4688 VDD.n3877 VDD.n126 66.2847
R4689 VDD.n3871 VDD.n126 66.2847
R4690 VDD.n3869 VDD.n126 66.2847
R4691 VDD.n3863 VDD.n126 66.2847
R4692 VDD.n3861 VDD.n126 66.2847
R4693 VDD.n3855 VDD.n126 66.2847
R4694 VDD.n3853 VDD.n126 66.2847
R4695 VDD.n3847 VDD.n126 66.2847
R4696 VDD.n222 VDD.n126 66.2847
R4697 VDD.n224 VDD.n126 66.2847
R4698 VDD.n3837 VDD.n126 66.2847
R4699 VDD.n3771 VDD.n126 66.2847
R4700 VDD.n3826 VDD.n126 66.2847
R4701 VDD.n3773 VDD.n126 66.2847
R4702 VDD.n3819 VDD.n126 66.2847
R4703 VDD.n3813 VDD.n126 66.2847
R4704 VDD.n3811 VDD.n126 66.2847
R4705 VDD.n3805 VDD.n126 66.2847
R4706 VDD.n3803 VDD.n126 66.2847
R4707 VDD.n3793 VDD.n126 66.2847
R4708 VDD.n4317 VDD.n4168 66.2847
R4709 VDD.n4388 VDD.n4168 66.2847
R4710 VDD.n4313 VDD.n4168 66.2847
R4711 VDD.n4395 VDD.n4168 66.2847
R4712 VDD.n4306 VDD.n4168 66.2847
R4713 VDD.n4402 VDD.n4168 66.2847
R4714 VDD.n4299 VDD.n4168 66.2847
R4715 VDD.n4409 VDD.n4168 66.2847
R4716 VDD.n4293 VDD.n4168 66.2847
R4717 VDD.n4418 VDD.n4168 66.2847
R4718 VDD.n4285 VDD.n4168 66.2847
R4719 VDD.n4425 VDD.n4168 66.2847
R4720 VDD.n4278 VDD.n4168 66.2847
R4721 VDD.n4432 VDD.n4168 66.2847
R4722 VDD.n4271 VDD.n4168 66.2847
R4723 VDD.n4439 VDD.n4168 66.2847
R4724 VDD.n4265 VDD.n4168 66.2847
R4725 VDD.n4448 VDD.n4168 66.2847
R4726 VDD.n4259 VDD.n4168 66.2847
R4727 VDD.n4455 VDD.n4168 66.2847
R4728 VDD.n4250 VDD.n4168 66.2847
R4729 VDD.n4462 VDD.n4168 66.2847
R4730 VDD.n4243 VDD.n4168 66.2847
R4731 VDD.n4469 VDD.n4168 66.2847
R4732 VDD.n4236 VDD.n4168 66.2847
R4733 VDD.n4476 VDD.n4168 66.2847
R4734 VDD.n4228 VDD.n4168 66.2847
R4735 VDD.n4483 VDD.n4168 66.2847
R4736 VDD.n4219 VDD.n4168 66.2847
R4737 VDD.n4490 VDD.n4168 66.2847
R4738 VDD.n4212 VDD.n4168 66.2847
R4739 VDD.n4497 VDD.n4168 66.2847
R4740 VDD.n4205 VDD.n4168 66.2847
R4741 VDD.n4504 VDD.n4168 66.2847
R4742 VDD.n4198 VDD.n4168 66.2847
R4743 VDD.n4514 VDD.n4168 66.2847
R4744 VDD.n4191 VDD.n4168 66.2847
R4745 VDD.n4521 VDD.n4168 66.2847
R4746 VDD.n4184 VDD.n4168 66.2847
R4747 VDD.n4528 VDD.n4168 66.2847
R4748 VDD.n4531 VDD.n4168 66.2847
R4749 VDD.n4172 VDD.n4168 66.2847
R4750 VDD.n4173 VDD.n4172 52.4337
R4751 VDD.n4531 VDD.n4530 52.4337
R4752 VDD.n4528 VDD.n4527 52.4337
R4753 VDD.n4523 VDD.n4184 52.4337
R4754 VDD.n4521 VDD.n4520 52.4337
R4755 VDD.n4516 VDD.n4191 52.4337
R4756 VDD.n4514 VDD.n4513 52.4337
R4757 VDD.n4506 VDD.n4198 52.4337
R4758 VDD.n4504 VDD.n4503 52.4337
R4759 VDD.n4499 VDD.n4205 52.4337
R4760 VDD.n4497 VDD.n4496 52.4337
R4761 VDD.n4492 VDD.n4212 52.4337
R4762 VDD.n4490 VDD.n4489 52.4337
R4763 VDD.n4485 VDD.n4219 52.4337
R4764 VDD.n4483 VDD.n4482 52.4337
R4765 VDD.n4478 VDD.n4228 52.4337
R4766 VDD.n4476 VDD.n4475 52.4337
R4767 VDD.n4471 VDD.n4236 52.4337
R4768 VDD.n4469 VDD.n4468 52.4337
R4769 VDD.n4464 VDD.n4243 52.4337
R4770 VDD.n4462 VDD.n4461 52.4337
R4771 VDD.n4457 VDD.n4250 52.4337
R4772 VDD.n4455 VDD.n4454 52.4337
R4773 VDD.n4450 VDD.n4259 52.4337
R4774 VDD.n4448 VDD.n4447 52.4337
R4775 VDD.n4441 VDD.n4265 52.4337
R4776 VDD.n4439 VDD.n4438 52.4337
R4777 VDD.n4434 VDD.n4271 52.4337
R4778 VDD.n4432 VDD.n4431 52.4337
R4779 VDD.n4427 VDD.n4278 52.4337
R4780 VDD.n4425 VDD.n4424 52.4337
R4781 VDD.n4420 VDD.n4285 52.4337
R4782 VDD.n4418 VDD.n4417 52.4337
R4783 VDD.n4411 VDD.n4293 52.4337
R4784 VDD.n4409 VDD.n4408 52.4337
R4785 VDD.n4404 VDD.n4299 52.4337
R4786 VDD.n4402 VDD.n4401 52.4337
R4787 VDD.n4397 VDD.n4306 52.4337
R4788 VDD.n4395 VDD.n4394 52.4337
R4789 VDD.n4390 VDD.n4313 52.4337
R4790 VDD.n4388 VDD.n4387 52.4337
R4791 VDD.n4318 VDD.n4317 52.4337
R4792 VDD.n3961 VDD.n127 52.4337
R4793 VDD.n3959 VDD.n130 52.4337
R4794 VDD.n3955 VDD.n3954 52.4337
R4795 VDD.n3948 VDD.n135 52.4337
R4796 VDD.n3947 VDD.n3946 52.4337
R4797 VDD.n3940 VDD.n141 52.4337
R4798 VDD.n3939 VDD.n3938 52.4337
R4799 VDD.n3931 VDD.n147 52.4337
R4800 VDD.n3930 VDD.n3929 52.4337
R4801 VDD.n3923 VDD.n155 52.4337
R4802 VDD.n3922 VDD.n3921 52.4337
R4803 VDD.n166 VDD.n161 52.4337
R4804 VDD.n3911 VDD.n168 52.4337
R4805 VDD.n3910 VDD.n3909 52.4337
R4806 VDD.n3903 VDD.n170 52.4337
R4807 VDD.n3902 VDD.n3901 52.4337
R4808 VDD.n3895 VDD.n176 52.4337
R4809 VDD.n3894 VDD.n3893 52.4337
R4810 VDD.n3887 VDD.n185 52.4337
R4811 VDD.n3886 VDD.n3885 52.4337
R4812 VDD.n3879 VDD.n191 52.4337
R4813 VDD.n3878 VDD.n3877 52.4337
R4814 VDD.n3871 VDD.n197 52.4337
R4815 VDD.n3870 VDD.n3869 52.4337
R4816 VDD.n3863 VDD.n203 52.4337
R4817 VDD.n3862 VDD.n3861 52.4337
R4818 VDD.n3855 VDD.n211 52.4337
R4819 VDD.n3854 VDD.n3853 52.4337
R4820 VDD.n3847 VDD.n217 52.4337
R4821 VDD.n3846 VDD.n222 52.4337
R4822 VDD.n3842 VDD.n224 52.4337
R4823 VDD.n3838 VDD.n3837 52.4337
R4824 VDD.n3771 VDD.n3765 52.4337
R4825 VDD.n3827 VDD.n3826 52.4337
R4826 VDD.n3824 VDD.n3773 52.4337
R4827 VDD.n3820 VDD.n3819 52.4337
R4828 VDD.n3813 VDD.n3777 52.4337
R4829 VDD.n3812 VDD.n3811 52.4337
R4830 VDD.n3805 VDD.n3783 52.4337
R4831 VDD.n3804 VDD.n3803 52.4337
R4832 VDD.n3793 VDD.n3789 52.4337
R4833 VDD.n2163 VDD.n1952 52.4337
R4834 VDD.n2161 VDD.n2160 52.4337
R4835 VDD.n2156 VDD.n1959 52.4337
R4836 VDD.n2154 VDD.n2153 52.4337
R4837 VDD.n2149 VDD.n1966 52.4337
R4838 VDD.n2147 VDD.n2146 52.4337
R4839 VDD.n2142 VDD.n1973 52.4337
R4840 VDD.n2140 VDD.n2139 52.4337
R4841 VDD.n2135 VDD.n1983 52.4337
R4842 VDD.n2133 VDD.n2132 52.4337
R4843 VDD.n2128 VDD.n1990 52.4337
R4844 VDD.n2126 VDD.n2125 52.4337
R4845 VDD.n1997 VDD.n1996 52.4337
R4846 VDD.n2117 VDD.n2116 52.4337
R4847 VDD.n2114 VDD.n2113 52.4337
R4848 VDD.n2109 VDD.n2007 52.4337
R4849 VDD.n2107 VDD.n2106 52.4337
R4850 VDD.n2102 VDD.n2015 52.4337
R4851 VDD.n2100 VDD.n2099 52.4337
R4852 VDD.n2095 VDD.n2022 52.4337
R4853 VDD.n2093 VDD.n2092 52.4337
R4854 VDD.n2088 VDD.n2029 52.4337
R4855 VDD.n2086 VDD.n2085 52.4337
R4856 VDD.n2081 VDD.n2038 52.4337
R4857 VDD.n2079 VDD.n2078 52.4337
R4858 VDD.n2072 VDD.n2044 52.4337
R4859 VDD.n2070 VDD.n2069 52.4337
R4860 VDD.n2065 VDD.n2051 52.4337
R4861 VDD.n2063 VDD.n2062 52.4337
R4862 VDD.n2058 VDD.n2057 52.4337
R4863 VDD.n2053 VDD.n2052 52.4337
R4864 VDD.n1192 VDD.n1162 52.4337
R4865 VDD.n1194 VDD.n1193 52.4337
R4866 VDD.n1195 VDD.n1169 52.4337
R4867 VDD.n1197 VDD.n1196 52.4337
R4868 VDD.n1198 VDD.n1174 52.4337
R4869 VDD.n1200 VDD.n1199 52.4337
R4870 VDD.n1201 VDD.n1179 52.4337
R4871 VDD.n1203 VDD.n1202 52.4337
R4872 VDD.n1204 VDD.n1184 52.4337
R4873 VDD.n1205 VDD.n1191 52.4337
R4874 VDD.n2173 VDD.n2172 52.4337
R4875 VDD.n1392 VDD.n1390 52.4337
R4876 VDD.n1398 VDD.n1397 52.4337
R4877 VDD.n1401 VDD.n1400 52.4337
R4878 VDD.n1406 VDD.n1405 52.4337
R4879 VDD.n1409 VDD.n1408 52.4337
R4880 VDD.n1414 VDD.n1413 52.4337
R4881 VDD.n1417 VDD.n1416 52.4337
R4882 VDD.n1424 VDD.n1423 52.4337
R4883 VDD.n1429 VDD.n1426 52.4337
R4884 VDD.n1432 VDD.n1431 52.4337
R4885 VDD.n1437 VDD.n1434 52.4337
R4886 VDD.n1440 VDD.n1439 52.4337
R4887 VDD.n1445 VDD.n1442 52.4337
R4888 VDD.n1448 VDD.n1447 52.4337
R4889 VDD.n1453 VDD.n1450 52.4337
R4890 VDD.n1456 VDD.n1455 52.4337
R4891 VDD.n1461 VDD.n1458 52.4337
R4892 VDD.n1464 VDD.n1463 52.4337
R4893 VDD.n1469 VDD.n1466 52.4337
R4894 VDD.n1472 VDD.n1471 52.4337
R4895 VDD.n1477 VDD.n1474 52.4337
R4896 VDD.n1480 VDD.n1479 52.4337
R4897 VDD.n1485 VDD.n1482 52.4337
R4898 VDD.n1488 VDD.n1487 52.4337
R4899 VDD.n1614 VDD.n1613 52.4337
R4900 VDD.n1611 VDD.n1494 52.4337
R4901 VDD.n1500 VDD.n1499 52.4337
R4902 VDD.n1505 VDD.n1502 52.4337
R4903 VDD.n1508 VDD.n1507 52.4337
R4904 VDD.n1513 VDD.n1510 52.4337
R4905 VDD.n1516 VDD.n1515 52.4337
R4906 VDD.n1522 VDD.n1518 52.4337
R4907 VDD.n1585 VDD.n1584 52.4337
R4908 VDD.n1582 VDD.n1524 52.4337
R4909 VDD.n1529 VDD.n1528 52.4337
R4910 VDD.n1534 VDD.n1531 52.4337
R4911 VDD.n1537 VDD.n1536 52.4337
R4912 VDD.n1542 VDD.n1539 52.4337
R4913 VDD.n1545 VDD.n1544 52.4337
R4914 VDD.n1550 VDD.n1547 52.4337
R4915 VDD.n1554 VDD.n1552 52.4337
R4916 VDD.n1393 VDD.n1392 52.4337
R4917 VDD.n1399 VDD.n1398 52.4337
R4918 VDD.n1402 VDD.n1401 52.4337
R4919 VDD.n1407 VDD.n1406 52.4337
R4920 VDD.n1410 VDD.n1409 52.4337
R4921 VDD.n1415 VDD.n1414 52.4337
R4922 VDD.n1418 VDD.n1417 52.4337
R4923 VDD.n1425 VDD.n1424 52.4337
R4924 VDD.n1430 VDD.n1429 52.4337
R4925 VDD.n1433 VDD.n1432 52.4337
R4926 VDD.n1438 VDD.n1437 52.4337
R4927 VDD.n1441 VDD.n1440 52.4337
R4928 VDD.n1446 VDD.n1445 52.4337
R4929 VDD.n1449 VDD.n1448 52.4337
R4930 VDD.n1454 VDD.n1453 52.4337
R4931 VDD.n1457 VDD.n1456 52.4337
R4932 VDD.n1462 VDD.n1461 52.4337
R4933 VDD.n1465 VDD.n1464 52.4337
R4934 VDD.n1470 VDD.n1469 52.4337
R4935 VDD.n1473 VDD.n1472 52.4337
R4936 VDD.n1478 VDD.n1477 52.4337
R4937 VDD.n1481 VDD.n1480 52.4337
R4938 VDD.n1486 VDD.n1485 52.4337
R4939 VDD.n1489 VDD.n1488 52.4337
R4940 VDD.n1613 VDD.n1612 52.4337
R4941 VDD.n1498 VDD.n1494 52.4337
R4942 VDD.n1501 VDD.n1500 52.4337
R4943 VDD.n1506 VDD.n1505 52.4337
R4944 VDD.n1509 VDD.n1508 52.4337
R4945 VDD.n1514 VDD.n1513 52.4337
R4946 VDD.n1517 VDD.n1516 52.4337
R4947 VDD.n1523 VDD.n1522 52.4337
R4948 VDD.n1584 VDD.n1583 52.4337
R4949 VDD.n1527 VDD.n1524 52.4337
R4950 VDD.n1530 VDD.n1529 52.4337
R4951 VDD.n1535 VDD.n1534 52.4337
R4952 VDD.n1538 VDD.n1537 52.4337
R4953 VDD.n1543 VDD.n1542 52.4337
R4954 VDD.n1546 VDD.n1545 52.4337
R4955 VDD.n1551 VDD.n1550 52.4337
R4956 VDD.n1555 VDD.n1554 52.4337
R4957 VDD.n2174 VDD.n2173 52.4337
R4958 VDD.n1205 VDD.n1185 52.4337
R4959 VDD.n1204 VDD.n1183 52.4337
R4960 VDD.n1203 VDD.n1180 52.4337
R4961 VDD.n1201 VDD.n1178 52.4337
R4962 VDD.n1200 VDD.n1175 52.4337
R4963 VDD.n1198 VDD.n1173 52.4337
R4964 VDD.n1197 VDD.n1170 52.4337
R4965 VDD.n1195 VDD.n1168 52.4337
R4966 VDD.n1194 VDD.n1163 52.4337
R4967 VDD.n1192 VDD.n1161 52.4337
R4968 VDD.n2054 VDD.n2053 52.4337
R4969 VDD.n2059 VDD.n2058 52.4337
R4970 VDD.n2064 VDD.n2063 52.4337
R4971 VDD.n2051 VDD.n2045 52.4337
R4972 VDD.n2071 VDD.n2070 52.4337
R4973 VDD.n2044 VDD.n2039 52.4337
R4974 VDD.n2080 VDD.n2079 52.4337
R4975 VDD.n2038 VDD.n2030 52.4337
R4976 VDD.n2087 VDD.n2086 52.4337
R4977 VDD.n2029 VDD.n2023 52.4337
R4978 VDD.n2094 VDD.n2093 52.4337
R4979 VDD.n2022 VDD.n2016 52.4337
R4980 VDD.n2101 VDD.n2100 52.4337
R4981 VDD.n2015 VDD.n2009 52.4337
R4982 VDD.n2108 VDD.n2107 52.4337
R4983 VDD.n2007 VDD.n1999 52.4337
R4984 VDD.n2115 VDD.n2114 52.4337
R4985 VDD.n2118 VDD.n2117 52.4337
R4986 VDD.n1996 VDD.n1991 52.4337
R4987 VDD.n2127 VDD.n2126 52.4337
R4988 VDD.n1990 VDD.n1984 52.4337
R4989 VDD.n2134 VDD.n2133 52.4337
R4990 VDD.n1983 VDD.n1974 52.4337
R4991 VDD.n2141 VDD.n2140 52.4337
R4992 VDD.n1973 VDD.n1967 52.4337
R4993 VDD.n2148 VDD.n2147 52.4337
R4994 VDD.n1966 VDD.n1960 52.4337
R4995 VDD.n2155 VDD.n2154 52.4337
R4996 VDD.n1959 VDD.n1953 52.4337
R4997 VDD.n2162 VDD.n2161 52.4337
R4998 VDD.n1952 VDD.n1211 52.4337
R4999 VDD.n3962 VDD.n3961 52.4337
R5000 VDD.n3956 VDD.n130 52.4337
R5001 VDD.n3954 VDD.n3953 52.4337
R5002 VDD.n3949 VDD.n3948 52.4337
R5003 VDD.n3946 VDD.n3945 52.4337
R5004 VDD.n3941 VDD.n3940 52.4337
R5005 VDD.n3938 VDD.n3937 52.4337
R5006 VDD.n3932 VDD.n3931 52.4337
R5007 VDD.n3929 VDD.n3928 52.4337
R5008 VDD.n3924 VDD.n3923 52.4337
R5009 VDD.n3921 VDD.n3920 52.4337
R5010 VDD.n167 VDD.n166 52.4337
R5011 VDD.n3912 VDD.n3911 52.4337
R5012 VDD.n3909 VDD.n3908 52.4337
R5013 VDD.n3904 VDD.n3903 52.4337
R5014 VDD.n3901 VDD.n3900 52.4337
R5015 VDD.n3896 VDD.n3895 52.4337
R5016 VDD.n3893 VDD.n3892 52.4337
R5017 VDD.n3888 VDD.n3887 52.4337
R5018 VDD.n3885 VDD.n3884 52.4337
R5019 VDD.n3880 VDD.n3879 52.4337
R5020 VDD.n3877 VDD.n3876 52.4337
R5021 VDD.n3872 VDD.n3871 52.4337
R5022 VDD.n3869 VDD.n3868 52.4337
R5023 VDD.n3864 VDD.n3863 52.4337
R5024 VDD.n3861 VDD.n3860 52.4337
R5025 VDD.n3856 VDD.n3855 52.4337
R5026 VDD.n3853 VDD.n3852 52.4337
R5027 VDD.n3848 VDD.n3847 52.4337
R5028 VDD.n3843 VDD.n222 52.4337
R5029 VDD.n3839 VDD.n224 52.4337
R5030 VDD.n3837 VDD.n3836 52.4337
R5031 VDD.n3772 VDD.n3771 52.4337
R5032 VDD.n3826 VDD.n3825 52.4337
R5033 VDD.n3821 VDD.n3773 52.4337
R5034 VDD.n3819 VDD.n3818 52.4337
R5035 VDD.n3814 VDD.n3813 52.4337
R5036 VDD.n3811 VDD.n3810 52.4337
R5037 VDD.n3806 VDD.n3805 52.4337
R5038 VDD.n3803 VDD.n3802 52.4337
R5039 VDD.n3794 VDD.n3793 52.4337
R5040 VDD.n4317 VDD.n4314 52.4337
R5041 VDD.n4389 VDD.n4388 52.4337
R5042 VDD.n4313 VDD.n4307 52.4337
R5043 VDD.n4396 VDD.n4395 52.4337
R5044 VDD.n4306 VDD.n4300 52.4337
R5045 VDD.n4403 VDD.n4402 52.4337
R5046 VDD.n4299 VDD.n4294 52.4337
R5047 VDD.n4410 VDD.n4409 52.4337
R5048 VDD.n4293 VDD.n4286 52.4337
R5049 VDD.n4419 VDD.n4418 52.4337
R5050 VDD.n4285 VDD.n4279 52.4337
R5051 VDD.n4426 VDD.n4425 52.4337
R5052 VDD.n4278 VDD.n4272 52.4337
R5053 VDD.n4433 VDD.n4432 52.4337
R5054 VDD.n4271 VDD.n4266 52.4337
R5055 VDD.n4440 VDD.n4439 52.4337
R5056 VDD.n4265 VDD.n4260 52.4337
R5057 VDD.n4449 VDD.n4448 52.4337
R5058 VDD.n4259 VDD.n4251 52.4337
R5059 VDD.n4456 VDD.n4455 52.4337
R5060 VDD.n4250 VDD.n4244 52.4337
R5061 VDD.n4463 VDD.n4462 52.4337
R5062 VDD.n4243 VDD.n4237 52.4337
R5063 VDD.n4470 VDD.n4469 52.4337
R5064 VDD.n4236 VDD.n4230 52.4337
R5065 VDD.n4477 VDD.n4476 52.4337
R5066 VDD.n4228 VDD.n4220 52.4337
R5067 VDD.n4484 VDD.n4483 52.4337
R5068 VDD.n4219 VDD.n4213 52.4337
R5069 VDD.n4491 VDD.n4490 52.4337
R5070 VDD.n4212 VDD.n4206 52.4337
R5071 VDD.n4498 VDD.n4497 52.4337
R5072 VDD.n4205 VDD.n4199 52.4337
R5073 VDD.n4505 VDD.n4504 52.4337
R5074 VDD.n4198 VDD.n4192 52.4337
R5075 VDD.n4515 VDD.n4514 52.4337
R5076 VDD.n4191 VDD.n4185 52.4337
R5077 VDD.n4522 VDD.n4521 52.4337
R5078 VDD.n4184 VDD.n4177 52.4337
R5079 VDD.n4529 VDD.n4528 52.4337
R5080 VDD.n4532 VDD.n4531 52.4337
R5081 VDD.n4172 VDD.n4169 52.4337
R5082 VDD.n2463 VDD.t137 45.7798
R5083 VDD.n228 VDD.t159 45.7798
R5084 VDD.n4385 VDD.n4321 43.6369
R5085 VDD.n179 VDD.n178 43.6369
R5086 VDD.n3834 VDD.n3833 43.6369
R5087 VDD.n3738 VDD.n245 39.2114
R5088 VDD.n3736 VDD.n3735 39.2114
R5089 VDD.n3731 VDD.n248 39.2114
R5090 VDD.n3729 VDD.n3728 39.2114
R5091 VDD.n3724 VDD.n3723 39.2114
R5092 VDD.n3719 VDD.n251 39.2114
R5093 VDD.n3717 VDD.n3716 39.2114
R5094 VDD.n3712 VDD.n256 39.2114
R5095 VDD.n3710 VDD.n3709 39.2114
R5096 VDD.n2910 VDD.n601 39.2114
R5097 VDD.n2914 VDD.n2913 39.2114
R5098 VDD.n2919 VDD.n2918 39.2114
R5099 VDD.n2922 VDD.n2921 39.2114
R5100 VDD.n2927 VDD.n2926 39.2114
R5101 VDD.n2930 VDD.n2929 39.2114
R5102 VDD.n2935 VDD.n2934 39.2114
R5103 VDD.n2938 VDD.n2937 39.2114
R5104 VDD.n2850 VDD.n603 39.2114
R5105 VDD.n2846 VDD.n604 39.2114
R5106 VDD.n2842 VDD.n605 39.2114
R5107 VDD.n2838 VDD.n606 39.2114
R5108 VDD.n2834 VDD.n607 39.2114
R5109 VDD.n2830 VDD.n608 39.2114
R5110 VDD.n2826 VDD.n609 39.2114
R5111 VDD.n2822 VDD.n610 39.2114
R5112 VDD.n2818 VDD.n611 39.2114
R5113 VDD.n2465 VDD.n2464 39.2114
R5114 VDD.n998 VDD.n980 39.2114
R5115 VDD.n2457 VDD.n981 39.2114
R5116 VDD.n2453 VDD.n982 39.2114
R5117 VDD.n2449 VDD.n983 39.2114
R5118 VDD.n2445 VDD.n984 39.2114
R5119 VDD.n2441 VDD.n985 39.2114
R5120 VDD.n2437 VDD.n986 39.2114
R5121 VDD.n3687 VDD.n3686 39.2114
R5122 VDD.n3684 VDD.n3683 39.2114
R5123 VDD.n3679 VDD.n3673 39.2114
R5124 VDD.n3677 VDD.n3676 39.2114
R5125 VDD.n3759 VDD.n227 39.2114
R5126 VDD.n3757 VDD.n3756 39.2114
R5127 VDD.n3752 VDD.n233 39.2114
R5128 VDD.n3750 VDD.n3749 39.2114
R5129 VDD.n3745 VDD.n236 39.2114
R5130 VDD.n3329 VDD.n3113 39.2114
R5131 VDD.n3328 VDD.n3327 39.2114
R5132 VDD.n3321 VDD.n3115 39.2114
R5133 VDD.n3320 VDD.n3319 39.2114
R5134 VDD.n3313 VDD.n3117 39.2114
R5135 VDD.n3312 VDD.n3311 39.2114
R5136 VDD.n3305 VDD.n3119 39.2114
R5137 VDD.n3304 VDD.n3303 39.2114
R5138 VDD.n3297 VDD.n3123 39.2114
R5139 VDD.n3330 VDD.n3329 39.2114
R5140 VDD.n3327 VDD.n3326 39.2114
R5141 VDD.n3322 VDD.n3321 39.2114
R5142 VDD.n3319 VDD.n3318 39.2114
R5143 VDD.n3314 VDD.n3313 39.2114
R5144 VDD.n3311 VDD.n3310 39.2114
R5145 VDD.n3306 VDD.n3305 39.2114
R5146 VDD.n3303 VDD.n3302 39.2114
R5147 VDD.n3298 VDD.n3297 39.2114
R5148 VDD.n236 VDD.n234 39.2114
R5149 VDD.n3751 VDD.n3750 39.2114
R5150 VDD.n233 VDD.n229 39.2114
R5151 VDD.n3758 VDD.n3757 39.2114
R5152 VDD.n3674 VDD.n227 39.2114
R5153 VDD.n3678 VDD.n3677 39.2114
R5154 VDD.n3673 VDD.n3671 39.2114
R5155 VDD.n3685 VDD.n3684 39.2114
R5156 VDD.n3688 VDD.n3687 39.2114
R5157 VDD.n2464 VDD.n979 39.2114
R5158 VDD.n2458 VDD.n980 39.2114
R5159 VDD.n2454 VDD.n981 39.2114
R5160 VDD.n2450 VDD.n982 39.2114
R5161 VDD.n2446 VDD.n983 39.2114
R5162 VDD.n2442 VDD.n984 39.2114
R5163 VDD.n2438 VDD.n985 39.2114
R5164 VDD.n2434 VDD.n986 39.2114
R5165 VDD.n2821 VDD.n611 39.2114
R5166 VDD.n2825 VDD.n610 39.2114
R5167 VDD.n2829 VDD.n609 39.2114
R5168 VDD.n2833 VDD.n608 39.2114
R5169 VDD.n2837 VDD.n607 39.2114
R5170 VDD.n2841 VDD.n606 39.2114
R5171 VDD.n2845 VDD.n605 39.2114
R5172 VDD.n2849 VDD.n604 39.2114
R5173 VDD.n2852 VDD.n603 39.2114
R5174 VDD.n2911 VDD.n2910 39.2114
R5175 VDD.n2913 VDD.n2907 39.2114
R5176 VDD.n2920 VDD.n2919 39.2114
R5177 VDD.n2921 VDD.n2905 39.2114
R5178 VDD.n2928 VDD.n2927 39.2114
R5179 VDD.n2929 VDD.n2903 39.2114
R5180 VDD.n2936 VDD.n2935 39.2114
R5181 VDD.n2939 VDD.n2938 39.2114
R5182 VDD.n3711 VDD.n3710 39.2114
R5183 VDD.n256 VDD.n252 39.2114
R5184 VDD.n3718 VDD.n3717 39.2114
R5185 VDD.n251 VDD.n249 39.2114
R5186 VDD.n3725 VDD.n3724 39.2114
R5187 VDD.n3730 VDD.n3729 39.2114
R5188 VDD.n248 VDD.n246 39.2114
R5189 VDD.n3737 VDD.n3736 39.2114
R5190 VDD.n245 VDD.n242 39.2114
R5191 VDD.n622 VDD.n612 39.2114
R5192 VDD.n2889 VDD.n613 39.2114
R5193 VDD.n2885 VDD.n614 39.2114
R5194 VDD.n2881 VDD.n615 39.2114
R5195 VDD.n2877 VDD.n616 39.2114
R5196 VDD.n2873 VDD.n617 39.2114
R5197 VDD.n2869 VDD.n618 39.2114
R5198 VDD.n2865 VDD.n619 39.2114
R5199 VDD.n2210 VDD.n988 39.2114
R5200 VDD.n2214 VDD.n989 39.2114
R5201 VDD.n2218 VDD.n990 39.2114
R5202 VDD.n2222 VDD.n991 39.2114
R5203 VDD.n2226 VDD.n992 39.2114
R5204 VDD.n2230 VDD.n993 39.2114
R5205 VDD.n2234 VDD.n994 39.2114
R5206 VDD.n2238 VDD.n995 39.2114
R5207 VDD.n2862 VDD.n619 39.2114
R5208 VDD.n2866 VDD.n618 39.2114
R5209 VDD.n2870 VDD.n617 39.2114
R5210 VDD.n2874 VDD.n616 39.2114
R5211 VDD.n2878 VDD.n615 39.2114
R5212 VDD.n2882 VDD.n614 39.2114
R5213 VDD.n2886 VDD.n613 39.2114
R5214 VDD.n2890 VDD.n612 39.2114
R5215 VDD.n2213 VDD.n988 39.2114
R5216 VDD.n2217 VDD.n989 39.2114
R5217 VDD.n2221 VDD.n990 39.2114
R5218 VDD.n2225 VDD.n991 39.2114
R5219 VDD.n2229 VDD.n992 39.2114
R5220 VDD.n2233 VDD.n993 39.2114
R5221 VDD.n2237 VDD.n994 39.2114
R5222 VDD.n2240 VDD.n995 39.2114
R5223 VDD.n2854 VDD.n2853 37.9322
R5224 VDD.n2819 VDD.n2816 37.9322
R5225 VDD.n2433 VDD.n2432 37.9322
R5226 VDD.n2467 VDD.n2466 37.9322
R5227 VDD.n3110 VDD.n2941 37.9322
R5228 VDD.n3708 VDD.n3707 37.9322
R5229 VDD.n3337 VDD.n600 37.9322
R5230 VDD.n3741 VDD.n3740 37.9322
R5231 VDD.n3690 VDD.n3689 37.9322
R5232 VDD.n3746 VDD.n235 37.9322
R5233 VDD.n3299 VDD.n3296 37.9322
R5234 VDD.n3333 VDD.n3332 37.9322
R5235 VDD.n2209 VDD.n972 37.9322
R5236 VDD.n2893 VDD.n623 37.9322
R5237 VDD.n2861 VDD.n2860 37.9322
R5238 VDD.n2244 VDD.n2242 37.9322
R5239 VDD.n1616 VDD.n1491 30.8369
R5240 VDD.n1558 VDD.n1557 30.8369
R5241 VDD.n1588 VDD.n1587 30.8369
R5242 VDD.n1643 VDD.n1642 30.8369
R5243 VDD.n1421 VDD.n1420 30.8369
R5244 VDD.n1977 VDD.n1976 30.8369
R5245 VDD.n2037 VDD.n2036 30.8369
R5246 VDD.n2175 VDD.n1190 30.8369
R5247 VDD.n1166 VDD.n1165 30.8369
R5248 VDD.n2006 VDD.n2005 30.8369
R5249 VDD.n3867 VDD.n207 30.8369
R5250 VDD.n3797 VDD.n3796 30.8369
R5251 VDD.n4258 VDD.n4257 30.8369
R5252 VDD.n4416 VDD.n4289 30.8369
R5253 VDD.n4227 VDD.n4226 30.8369
R5254 VDD.n4510 VDD.n4509 30.8369
R5255 VDD.n3935 VDD.n151 30.8369
R5256 VDD.n2236 VDD.n1155 24.049
R5257 VDD.n2867 VDD.n625 24.049
R5258 VDD.n3714 VDD.n254 24.049
R5259 VDD.n2902 VDD.n2901 24.049
R5260 VDD.n2824 VDD.n635 24.049
R5261 VDD.n2439 VDD.n1001 24.049
R5262 VDD.n232 VDD.n231 24.049
R5263 VDD.n3122 VDD.n3121 24.049
R5264 VDD.n7 VDD.t160 22.3407
R5265 VDD.n7 VDD.t134 22.3407
R5266 VDD.n8 VDD.t156 22.3407
R5267 VDD.n8 VDD.t152 22.3407
R5268 VDD.n10 VDD.t154 22.3407
R5269 VDD.n10 VDD.t148 22.3407
R5270 VDD.n12 VDD.t150 22.3407
R5271 VDD.n12 VDD.t145 22.3407
R5272 VDD.n5 VDD.t129 22.3407
R5273 VDD.n5 VDD.t126 22.3407
R5274 VDD.n3 VDD.t158 22.3407
R5275 VDD.n3 VDD.t136 22.3407
R5276 VDD.n1 VDD.t140 22.3407
R5277 VDD.n1 VDD.t143 22.3407
R5278 VDD.n0 VDD.t132 22.3407
R5279 VDD.n0 VDD.t138 22.3407
R5280 VDD.n1696 VDD.n1389 19.5443
R5281 VDD.n2170 VDD.n1206 19.5443
R5282 VDD.n3969 VDD.n126 19.5443
R5283 VDD.n4540 VDD.n4168 19.5443
R5284 VDD.n1698 VDD.n1386 19.3944
R5285 VDD.n1702 VDD.n1386 19.3944
R5286 VDD.n1702 VDD.n1375 19.3944
R5287 VDD.n1714 VDD.n1375 19.3944
R5288 VDD.n1714 VDD.n1373 19.3944
R5289 VDD.n1718 VDD.n1373 19.3944
R5290 VDD.n1718 VDD.n1364 19.3944
R5291 VDD.n1730 VDD.n1364 19.3944
R5292 VDD.n1730 VDD.n1362 19.3944
R5293 VDD.n1734 VDD.n1362 19.3944
R5294 VDD.n1734 VDD.n1352 19.3944
R5295 VDD.n1746 VDD.n1352 19.3944
R5296 VDD.n1746 VDD.n1350 19.3944
R5297 VDD.n1750 VDD.n1350 19.3944
R5298 VDD.n1750 VDD.n1340 19.3944
R5299 VDD.n1762 VDD.n1340 19.3944
R5300 VDD.n1762 VDD.n1338 19.3944
R5301 VDD.n1766 VDD.n1338 19.3944
R5302 VDD.n1766 VDD.n1329 19.3944
R5303 VDD.n1779 VDD.n1329 19.3944
R5304 VDD.n1779 VDD.n1327 19.3944
R5305 VDD.n1783 VDD.n1327 19.3944
R5306 VDD.n1783 VDD.n1317 19.3944
R5307 VDD.n1795 VDD.n1317 19.3944
R5308 VDD.n1795 VDD.n1315 19.3944
R5309 VDD.n1799 VDD.n1315 19.3944
R5310 VDD.n1799 VDD.n1305 19.3944
R5311 VDD.n1811 VDD.n1305 19.3944
R5312 VDD.n1811 VDD.n1303 19.3944
R5313 VDD.n1815 VDD.n1303 19.3944
R5314 VDD.n1815 VDD.n1293 19.3944
R5315 VDD.n1841 VDD.n1293 19.3944
R5316 VDD.n1841 VDD.n1291 19.3944
R5317 VDD.n1845 VDD.n1291 19.3944
R5318 VDD.n1845 VDD.n1281 19.3944
R5319 VDD.n1857 VDD.n1281 19.3944
R5320 VDD.n1857 VDD.n1279 19.3944
R5321 VDD.n1861 VDD.n1279 19.3944
R5322 VDD.n1861 VDD.n1269 19.3944
R5323 VDD.n1873 VDD.n1269 19.3944
R5324 VDD.n1873 VDD.n1267 19.3944
R5325 VDD.n1877 VDD.n1267 19.3944
R5326 VDD.n1877 VDD.n1257 19.3944
R5327 VDD.n1889 VDD.n1257 19.3944
R5328 VDD.n1889 VDD.n1255 19.3944
R5329 VDD.n1893 VDD.n1255 19.3944
R5330 VDD.n1893 VDD.n1245 19.3944
R5331 VDD.n1905 VDD.n1245 19.3944
R5332 VDD.n1905 VDD.n1243 19.3944
R5333 VDD.n1909 VDD.n1243 19.3944
R5334 VDD.n1909 VDD.n1233 19.3944
R5335 VDD.n1921 VDD.n1233 19.3944
R5336 VDD.n1921 VDD.n1231 19.3944
R5337 VDD.n1925 VDD.n1231 19.3944
R5338 VDD.n1925 VDD.n1221 19.3944
R5339 VDD.n1937 VDD.n1221 19.3944
R5340 VDD.n1937 VDD.n1218 19.3944
R5341 VDD.n1943 VDD.n1218 19.3944
R5342 VDD.n1943 VDD.n1219 19.3944
R5343 VDD.n1219 VDD.n1208 19.3944
R5344 VDD.n1581 VDD.n1521 19.3944
R5345 VDD.n1581 VDD.n1525 19.3944
R5346 VDD.n1577 VDD.n1525 19.3944
R5347 VDD.n1577 VDD.n1576 19.3944
R5348 VDD.n1576 VDD.n1575 19.3944
R5349 VDD.n1575 VDD.n1532 19.3944
R5350 VDD.n1571 VDD.n1532 19.3944
R5351 VDD.n1571 VDD.n1570 19.3944
R5352 VDD.n1570 VDD.n1569 19.3944
R5353 VDD.n1569 VDD.n1540 19.3944
R5354 VDD.n1565 VDD.n1540 19.3944
R5355 VDD.n1565 VDD.n1564 19.3944
R5356 VDD.n1564 VDD.n1563 19.3944
R5357 VDD.n1563 VDD.n1548 19.3944
R5358 VDD.n1559 VDD.n1548 19.3944
R5359 VDD.n1615 VDD.n1493 19.3944
R5360 VDD.n1610 VDD.n1493 19.3944
R5361 VDD.n1610 VDD.n1495 19.3944
R5362 VDD.n1606 VDD.n1495 19.3944
R5363 VDD.n1606 VDD.n1605 19.3944
R5364 VDD.n1605 VDD.n1604 19.3944
R5365 VDD.n1604 VDD.n1503 19.3944
R5366 VDD.n1600 VDD.n1503 19.3944
R5367 VDD.n1600 VDD.n1599 19.3944
R5368 VDD.n1599 VDD.n1598 19.3944
R5369 VDD.n1598 VDD.n1511 19.3944
R5370 VDD.n1594 VDD.n1511 19.3944
R5371 VDD.n1594 VDD.n1593 19.3944
R5372 VDD.n1593 VDD.n1592 19.3944
R5373 VDD.n1592 VDD.n1519 19.3944
R5374 VDD.n1640 VDD.n1639 19.3944
R5375 VDD.n1639 VDD.n1459 19.3944
R5376 VDD.n1635 VDD.n1459 19.3944
R5377 VDD.n1635 VDD.n1634 19.3944
R5378 VDD.n1634 VDD.n1633 19.3944
R5379 VDD.n1633 VDD.n1467 19.3944
R5380 VDD.n1629 VDD.n1467 19.3944
R5381 VDD.n1629 VDD.n1628 19.3944
R5382 VDD.n1628 VDD.n1627 19.3944
R5383 VDD.n1627 VDD.n1475 19.3944
R5384 VDD.n1623 VDD.n1475 19.3944
R5385 VDD.n1623 VDD.n1622 19.3944
R5386 VDD.n1622 VDD.n1621 19.3944
R5387 VDD.n1621 VDD.n1483 19.3944
R5388 VDD.n1617 VDD.n1483 19.3944
R5389 VDD.n1617 VDD.n1616 19.3944
R5390 VDD.n1668 VDD.n1667 19.3944
R5391 VDD.n1667 VDD.n1666 19.3944
R5392 VDD.n1666 VDD.n1427 19.3944
R5393 VDD.n1662 VDD.n1427 19.3944
R5394 VDD.n1662 VDD.n1661 19.3944
R5395 VDD.n1661 VDD.n1660 19.3944
R5396 VDD.n1660 VDD.n1435 19.3944
R5397 VDD.n1656 VDD.n1435 19.3944
R5398 VDD.n1656 VDD.n1655 19.3944
R5399 VDD.n1655 VDD.n1654 19.3944
R5400 VDD.n1654 VDD.n1443 19.3944
R5401 VDD.n1650 VDD.n1443 19.3944
R5402 VDD.n1650 VDD.n1649 19.3944
R5403 VDD.n1649 VDD.n1648 19.3944
R5404 VDD.n1648 VDD.n1451 19.3944
R5405 VDD.n1644 VDD.n1451 19.3944
R5406 VDD.n1691 VDD.n1690 19.3944
R5407 VDD.n1690 VDD.n1689 19.3944
R5408 VDD.n1689 VDD.n1395 19.3944
R5409 VDD.n1685 VDD.n1395 19.3944
R5410 VDD.n1685 VDD.n1684 19.3944
R5411 VDD.n1684 VDD.n1683 19.3944
R5412 VDD.n1683 VDD.n1403 19.3944
R5413 VDD.n1679 VDD.n1403 19.3944
R5414 VDD.n1679 VDD.n1678 19.3944
R5415 VDD.n1678 VDD.n1677 19.3944
R5416 VDD.n1677 VDD.n1411 19.3944
R5417 VDD.n1673 VDD.n1411 19.3944
R5418 VDD.n1673 VDD.n1672 19.3944
R5419 VDD.n1672 VDD.n1671 19.3944
R5420 VDD.n1694 VDD.n1382 19.3944
R5421 VDD.n1706 VDD.n1382 19.3944
R5422 VDD.n1706 VDD.n1380 19.3944
R5423 VDD.n1710 VDD.n1380 19.3944
R5424 VDD.n1710 VDD.n1370 19.3944
R5425 VDD.n1722 VDD.n1370 19.3944
R5426 VDD.n1722 VDD.n1368 19.3944
R5427 VDD.n1726 VDD.n1368 19.3944
R5428 VDD.n1726 VDD.n1358 19.3944
R5429 VDD.n1738 VDD.n1358 19.3944
R5430 VDD.n1738 VDD.n1356 19.3944
R5431 VDD.n1742 VDD.n1356 19.3944
R5432 VDD.n1742 VDD.n1346 19.3944
R5433 VDD.n1754 VDD.n1346 19.3944
R5434 VDD.n1754 VDD.n1344 19.3944
R5435 VDD.n1758 VDD.n1344 19.3944
R5436 VDD.n1758 VDD.n1334 19.3944
R5437 VDD.n1771 VDD.n1334 19.3944
R5438 VDD.n1771 VDD.n1332 19.3944
R5439 VDD.n1775 VDD.n1332 19.3944
R5440 VDD.n1775 VDD.n1323 19.3944
R5441 VDD.n1787 VDD.n1323 19.3944
R5442 VDD.n1787 VDD.n1321 19.3944
R5443 VDD.n1791 VDD.n1321 19.3944
R5444 VDD.n1791 VDD.n1311 19.3944
R5445 VDD.n1803 VDD.n1311 19.3944
R5446 VDD.n1803 VDD.n1309 19.3944
R5447 VDD.n1807 VDD.n1309 19.3944
R5448 VDD.n1807 VDD.n1299 19.3944
R5449 VDD.n1818 VDD.n1299 19.3944
R5450 VDD.n1818 VDD.n1297 19.3944
R5451 VDD.n1837 VDD.n1297 19.3944
R5452 VDD.n1837 VDD.n1287 19.3944
R5453 VDD.n1849 VDD.n1287 19.3944
R5454 VDD.n1849 VDD.n1285 19.3944
R5455 VDD.n1853 VDD.n1285 19.3944
R5456 VDD.n1853 VDD.n1275 19.3944
R5457 VDD.n1865 VDD.n1275 19.3944
R5458 VDD.n1865 VDD.n1273 19.3944
R5459 VDD.n1869 VDD.n1273 19.3944
R5460 VDD.n1869 VDD.n1263 19.3944
R5461 VDD.n1881 VDD.n1263 19.3944
R5462 VDD.n1881 VDD.n1261 19.3944
R5463 VDD.n1885 VDD.n1261 19.3944
R5464 VDD.n1885 VDD.n1251 19.3944
R5465 VDD.n1897 VDD.n1251 19.3944
R5466 VDD.n1897 VDD.n1249 19.3944
R5467 VDD.n1901 VDD.n1249 19.3944
R5468 VDD.n1901 VDD.n1239 19.3944
R5469 VDD.n1913 VDD.n1239 19.3944
R5470 VDD.n1913 VDD.n1237 19.3944
R5471 VDD.n1917 VDD.n1237 19.3944
R5472 VDD.n1917 VDD.n1227 19.3944
R5473 VDD.n1929 VDD.n1227 19.3944
R5474 VDD.n1929 VDD.n1225 19.3944
R5475 VDD.n1933 VDD.n1225 19.3944
R5476 VDD.n1933 VDD.n1214 19.3944
R5477 VDD.n1947 VDD.n1214 19.3944
R5478 VDD.n1947 VDD.n1212 19.3944
R5479 VDD.n2168 VDD.n1212 19.3944
R5480 VDD.n2165 VDD.n2164 19.3944
R5481 VDD.n2164 VDD.n1951 19.3944
R5482 VDD.n2159 VDD.n1951 19.3944
R5483 VDD.n2159 VDD.n2158 19.3944
R5484 VDD.n2158 VDD.n2157 19.3944
R5485 VDD.n2157 VDD.n1958 19.3944
R5486 VDD.n2152 VDD.n1958 19.3944
R5487 VDD.n2152 VDD.n2151 19.3944
R5488 VDD.n2151 VDD.n2150 19.3944
R5489 VDD.n2150 VDD.n1965 19.3944
R5490 VDD.n2145 VDD.n1965 19.3944
R5491 VDD.n2145 VDD.n2144 19.3944
R5492 VDD.n2144 VDD.n2143 19.3944
R5493 VDD.n2143 VDD.n1972 19.3944
R5494 VDD.n2199 VDD.n2198 19.3944
R5495 VDD.n2198 VDD.n2197 19.3944
R5496 VDD.n2197 VDD.n1171 19.3944
R5497 VDD.n2193 VDD.n1171 19.3944
R5498 VDD.n2193 VDD.n2192 19.3944
R5499 VDD.n2192 VDD.n2191 19.3944
R5500 VDD.n2191 VDD.n1176 19.3944
R5501 VDD.n2187 VDD.n1176 19.3944
R5502 VDD.n2187 VDD.n2186 19.3944
R5503 VDD.n2186 VDD.n2185 19.3944
R5504 VDD.n2185 VDD.n1181 19.3944
R5505 VDD.n2181 VDD.n1181 19.3944
R5506 VDD.n2181 VDD.n2180 19.3944
R5507 VDD.n2180 VDD.n2179 19.3944
R5508 VDD.n2179 VDD.n1186 19.3944
R5509 VDD.n2077 VDD.n2040 19.3944
R5510 VDD.n2073 VDD.n2040 19.3944
R5511 VDD.n2073 VDD.n2043 19.3944
R5512 VDD.n2068 VDD.n2043 19.3944
R5513 VDD.n2068 VDD.n2067 19.3944
R5514 VDD.n2067 VDD.n2066 19.3944
R5515 VDD.n2066 VDD.n2050 19.3944
R5516 VDD.n2061 VDD.n2050 19.3944
R5517 VDD.n2061 VDD.n2060 19.3944
R5518 VDD.n2056 VDD.n2055 19.3944
R5519 VDD.n2205 VDD.n1160 19.3944
R5520 VDD.n2205 VDD.n2204 19.3944
R5521 VDD.n2204 VDD.n2203 19.3944
R5522 VDD.n2105 VDD.n2008 19.3944
R5523 VDD.n2105 VDD.n2104 19.3944
R5524 VDD.n2104 VDD.n2103 19.3944
R5525 VDD.n2103 VDD.n2014 19.3944
R5526 VDD.n2098 VDD.n2014 19.3944
R5527 VDD.n2098 VDD.n2097 19.3944
R5528 VDD.n2097 VDD.n2096 19.3944
R5529 VDD.n2096 VDD.n2021 19.3944
R5530 VDD.n2091 VDD.n2021 19.3944
R5531 VDD.n2091 VDD.n2090 19.3944
R5532 VDD.n2090 VDD.n2089 19.3944
R5533 VDD.n2089 VDD.n2028 19.3944
R5534 VDD.n2084 VDD.n2028 19.3944
R5535 VDD.n2084 VDD.n2083 19.3944
R5536 VDD.n2083 VDD.n2082 19.3944
R5537 VDD.n2082 VDD.n2037 19.3944
R5538 VDD.n2138 VDD.n2137 19.3944
R5539 VDD.n2137 VDD.n2136 19.3944
R5540 VDD.n2136 VDD.n1982 19.3944
R5541 VDD.n2131 VDD.n1982 19.3944
R5542 VDD.n2131 VDD.n2130 19.3944
R5543 VDD.n2130 VDD.n2129 19.3944
R5544 VDD.n2129 VDD.n1989 19.3944
R5545 VDD.n2124 VDD.n2123 19.3944
R5546 VDD.n2119 VDD.n1993 19.3944
R5547 VDD.n2119 VDD.n1995 19.3944
R5548 VDD.n1998 VDD.n1995 19.3944
R5549 VDD.n2112 VDD.n1998 19.3944
R5550 VDD.n2112 VDD.n2111 19.3944
R5551 VDD.n2111 VDD.n2110 19.3944
R5552 VDD.n3828 VDD.n3768 19.3944
R5553 VDD.n3828 VDD.n3770 19.3944
R5554 VDD.n3823 VDD.n3770 19.3944
R5555 VDD.n3823 VDD.n3822 19.3944
R5556 VDD.n3822 VDD.n3776 19.3944
R5557 VDD.n3817 VDD.n3776 19.3944
R5558 VDD.n3817 VDD.n3816 19.3944
R5559 VDD.n3816 VDD.n3815 19.3944
R5560 VDD.n3815 VDD.n3782 19.3944
R5561 VDD.n3809 VDD.n3782 19.3944
R5562 VDD.n3809 VDD.n3808 19.3944
R5563 VDD.n3808 VDD.n3807 19.3944
R5564 VDD.n3807 VDD.n3788 19.3944
R5565 VDD.n3801 VDD.n3788 19.3944
R5566 VDD.n3801 VDD.n3800 19.3944
R5567 VDD.n3971 VDD.n123 19.3944
R5568 VDD.n3975 VDD.n123 19.3944
R5569 VDD.n3975 VDD.n112 19.3944
R5570 VDD.n3987 VDD.n112 19.3944
R5571 VDD.n3987 VDD.n110 19.3944
R5572 VDD.n3991 VDD.n110 19.3944
R5573 VDD.n3991 VDD.n101 19.3944
R5574 VDD.n4003 VDD.n101 19.3944
R5575 VDD.n4003 VDD.n99 19.3944
R5576 VDD.n4007 VDD.n99 19.3944
R5577 VDD.n4007 VDD.n89 19.3944
R5578 VDD.n4019 VDD.n89 19.3944
R5579 VDD.n4019 VDD.n87 19.3944
R5580 VDD.n4023 VDD.n87 19.3944
R5581 VDD.n4023 VDD.n77 19.3944
R5582 VDD.n4035 VDD.n77 19.3944
R5583 VDD.n4035 VDD.n75 19.3944
R5584 VDD.n4039 VDD.n75 19.3944
R5585 VDD.n4039 VDD.n66 19.3944
R5586 VDD.n4052 VDD.n66 19.3944
R5587 VDD.n4052 VDD.n64 19.3944
R5588 VDD.n4056 VDD.n64 19.3944
R5589 VDD.n4056 VDD.n54 19.3944
R5590 VDD.n4068 VDD.n54 19.3944
R5591 VDD.n4068 VDD.n52 19.3944
R5592 VDD.n4072 VDD.n52 19.3944
R5593 VDD.n4072 VDD.n42 19.3944
R5594 VDD.n4084 VDD.n42 19.3944
R5595 VDD.n4084 VDD.n40 19.3944
R5596 VDD.n4600 VDD.n40 19.3944
R5597 VDD.n4600 VDD.n4599 19.3944
R5598 VDD.n4599 VDD.n4598 19.3944
R5599 VDD.n4598 VDD.n4090 19.3944
R5600 VDD.n4343 VDD.n4090 19.3944
R5601 VDD.n4344 VDD.n4343 19.3944
R5602 VDD.n4345 VDD.n4344 19.3944
R5603 VDD.n4345 VDD.n4339 19.3944
R5604 VDD.n4349 VDD.n4339 19.3944
R5605 VDD.n4350 VDD.n4349 19.3944
R5606 VDD.n4351 VDD.n4350 19.3944
R5607 VDD.n4351 VDD.n4336 19.3944
R5608 VDD.n4355 VDD.n4336 19.3944
R5609 VDD.n4356 VDD.n4355 19.3944
R5610 VDD.n4357 VDD.n4356 19.3944
R5611 VDD.n4357 VDD.n4333 19.3944
R5612 VDD.n4361 VDD.n4333 19.3944
R5613 VDD.n4362 VDD.n4361 19.3944
R5614 VDD.n4363 VDD.n4362 19.3944
R5615 VDD.n4363 VDD.n4330 19.3944
R5616 VDD.n4367 VDD.n4330 19.3944
R5617 VDD.n4368 VDD.n4367 19.3944
R5618 VDD.n4369 VDD.n4368 19.3944
R5619 VDD.n4369 VDD.n4327 19.3944
R5620 VDD.n4373 VDD.n4327 19.3944
R5621 VDD.n4374 VDD.n4373 19.3944
R5622 VDD.n4375 VDD.n4374 19.3944
R5623 VDD.n4375 VDD.n4324 19.3944
R5624 VDD.n4379 VDD.n4324 19.3944
R5625 VDD.n4380 VDD.n4379 19.3944
R5626 VDD.n4381 VDD.n4380 19.3944
R5627 VDD.n4412 VDD.n4287 19.3944
R5628 VDD.n4412 VDD.n4292 19.3944
R5629 VDD.n4407 VDD.n4292 19.3944
R5630 VDD.n4407 VDD.n4406 19.3944
R5631 VDD.n4406 VDD.n4405 19.3944
R5632 VDD.n4405 VDD.n4298 19.3944
R5633 VDD.n4400 VDD.n4298 19.3944
R5634 VDD.n4400 VDD.n4399 19.3944
R5635 VDD.n4399 VDD.n4398 19.3944
R5636 VDD.n4398 VDD.n4305 19.3944
R5637 VDD.n4393 VDD.n4305 19.3944
R5638 VDD.n4393 VDD.n4392 19.3944
R5639 VDD.n4392 VDD.n4391 19.3944
R5640 VDD.n4391 VDD.n4312 19.3944
R5641 VDD.n4386 VDD.n4312 19.3944
R5642 VDD.n4446 VDD.n4261 19.3944
R5643 VDD.n4442 VDD.n4261 19.3944
R5644 VDD.n4442 VDD.n4264 19.3944
R5645 VDD.n4437 VDD.n4264 19.3944
R5646 VDD.n4437 VDD.n4436 19.3944
R5647 VDD.n4436 VDD.n4435 19.3944
R5648 VDD.n4435 VDD.n4270 19.3944
R5649 VDD.n4430 VDD.n4270 19.3944
R5650 VDD.n4430 VDD.n4429 19.3944
R5651 VDD.n4429 VDD.n4428 19.3944
R5652 VDD.n4428 VDD.n4277 19.3944
R5653 VDD.n4423 VDD.n4277 19.3944
R5654 VDD.n4423 VDD.n4422 19.3944
R5655 VDD.n4422 VDD.n4421 19.3944
R5656 VDD.n4421 VDD.n4284 19.3944
R5657 VDD.n4474 VDD.n4229 19.3944
R5658 VDD.n4474 VDD.n4473 19.3944
R5659 VDD.n4473 VDD.n4472 19.3944
R5660 VDD.n4472 VDD.n4235 19.3944
R5661 VDD.n4467 VDD.n4235 19.3944
R5662 VDD.n4467 VDD.n4466 19.3944
R5663 VDD.n4466 VDD.n4465 19.3944
R5664 VDD.n4465 VDD.n4242 19.3944
R5665 VDD.n4460 VDD.n4242 19.3944
R5666 VDD.n4460 VDD.n4459 19.3944
R5667 VDD.n4459 VDD.n4458 19.3944
R5668 VDD.n4458 VDD.n4249 19.3944
R5669 VDD.n4453 VDD.n4249 19.3944
R5670 VDD.n4453 VDD.n4452 19.3944
R5671 VDD.n4452 VDD.n4451 19.3944
R5672 VDD.n4451 VDD.n4258 19.3944
R5673 VDD.n4507 VDD.n4197 19.3944
R5674 VDD.n4502 VDD.n4197 19.3944
R5675 VDD.n4502 VDD.n4501 19.3944
R5676 VDD.n4501 VDD.n4500 19.3944
R5677 VDD.n4500 VDD.n4204 19.3944
R5678 VDD.n4495 VDD.n4204 19.3944
R5679 VDD.n4495 VDD.n4494 19.3944
R5680 VDD.n4494 VDD.n4493 19.3944
R5681 VDD.n4493 VDD.n4211 19.3944
R5682 VDD.n4488 VDD.n4211 19.3944
R5683 VDD.n4488 VDD.n4487 19.3944
R5684 VDD.n4487 VDD.n4486 19.3944
R5685 VDD.n4486 VDD.n4218 19.3944
R5686 VDD.n4481 VDD.n4218 19.3944
R5687 VDD.n4481 VDD.n4480 19.3944
R5688 VDD.n4480 VDD.n4479 19.3944
R5689 VDD.n4535 VDD.n4534 19.3944
R5690 VDD.n4534 VDD.n4533 19.3944
R5691 VDD.n4533 VDD.n4175 19.3944
R5692 VDD.n4176 VDD.n4175 19.3944
R5693 VDD.n4526 VDD.n4176 19.3944
R5694 VDD.n4526 VDD.n4525 19.3944
R5695 VDD.n4525 VDD.n4524 19.3944
R5696 VDD.n4524 VDD.n4183 19.3944
R5697 VDD.n4519 VDD.n4183 19.3944
R5698 VDD.n4519 VDD.n4518 19.3944
R5699 VDD.n4518 VDD.n4517 19.3944
R5700 VDD.n4517 VDD.n4190 19.3944
R5701 VDD.n4512 VDD.n4190 19.3944
R5702 VDD.n4512 VDD.n4511 19.3944
R5703 VDD.n3967 VDD.n119 19.3944
R5704 VDD.n3979 VDD.n119 19.3944
R5705 VDD.n3979 VDD.n117 19.3944
R5706 VDD.n3983 VDD.n117 19.3944
R5707 VDD.n3983 VDD.n107 19.3944
R5708 VDD.n3995 VDD.n107 19.3944
R5709 VDD.n3995 VDD.n105 19.3944
R5710 VDD.n3999 VDD.n105 19.3944
R5711 VDD.n3999 VDD.n95 19.3944
R5712 VDD.n4011 VDD.n95 19.3944
R5713 VDD.n4011 VDD.n93 19.3944
R5714 VDD.n4015 VDD.n93 19.3944
R5715 VDD.n4015 VDD.n83 19.3944
R5716 VDD.n4027 VDD.n83 19.3944
R5717 VDD.n4027 VDD.n81 19.3944
R5718 VDD.n4031 VDD.n81 19.3944
R5719 VDD.n4031 VDD.n71 19.3944
R5720 VDD.n4044 VDD.n71 19.3944
R5721 VDD.n4044 VDD.n69 19.3944
R5722 VDD.n4048 VDD.n69 19.3944
R5723 VDD.n4048 VDD.n60 19.3944
R5724 VDD.n4060 VDD.n60 19.3944
R5725 VDD.n4060 VDD.n58 19.3944
R5726 VDD.n4064 VDD.n58 19.3944
R5727 VDD.n4064 VDD.n48 19.3944
R5728 VDD.n4076 VDD.n48 19.3944
R5729 VDD.n4076 VDD.n46 19.3944
R5730 VDD.n4080 VDD.n46 19.3944
R5731 VDD.n4080 VDD.n32 19.3944
R5732 VDD.n4603 VDD.n32 19.3944
R5733 VDD.n4603 VDD.n33 19.3944
R5734 VDD.n4594 VDD.n33 19.3944
R5735 VDD.n4594 VDD.n4593 19.3944
R5736 VDD.n4593 VDD.n4592 19.3944
R5737 VDD.n4592 VDD.n4097 19.3944
R5738 VDD.n4586 VDD.n4097 19.3944
R5739 VDD.n4586 VDD.n4585 19.3944
R5740 VDD.n4585 VDD.n4584 19.3944
R5741 VDD.n4584 VDD.n4108 19.3944
R5742 VDD.n4578 VDD.n4108 19.3944
R5743 VDD.n4578 VDD.n4577 19.3944
R5744 VDD.n4577 VDD.n4576 19.3944
R5745 VDD.n4576 VDD.n4118 19.3944
R5746 VDD.n4570 VDD.n4118 19.3944
R5747 VDD.n4570 VDD.n4569 19.3944
R5748 VDD.n4569 VDD.n4568 19.3944
R5749 VDD.n4568 VDD.n4130 19.3944
R5750 VDD.n4562 VDD.n4130 19.3944
R5751 VDD.n4562 VDD.n4561 19.3944
R5752 VDD.n4561 VDD.n4560 19.3944
R5753 VDD.n4560 VDD.n4141 19.3944
R5754 VDD.n4554 VDD.n4141 19.3944
R5755 VDD.n4554 VDD.n4553 19.3944
R5756 VDD.n4553 VDD.n4552 19.3944
R5757 VDD.n4552 VDD.n4152 19.3944
R5758 VDD.n4546 VDD.n4152 19.3944
R5759 VDD.n4546 VDD.n4545 19.3944
R5760 VDD.n4545 VDD.n4544 19.3944
R5761 VDD.n4544 VDD.n4163 19.3944
R5762 VDD.n4538 VDD.n4163 19.3944
R5763 VDD.n3964 VDD.n3963 19.3944
R5764 VDD.n3963 VDD.n129 19.3944
R5765 VDD.n3958 VDD.n129 19.3944
R5766 VDD.n3958 VDD.n3957 19.3944
R5767 VDD.n3957 VDD.n134 19.3944
R5768 VDD.n3952 VDD.n134 19.3944
R5769 VDD.n3952 VDD.n3951 19.3944
R5770 VDD.n3951 VDD.n3950 19.3944
R5771 VDD.n3950 VDD.n140 19.3944
R5772 VDD.n3944 VDD.n140 19.3944
R5773 VDD.n3944 VDD.n3943 19.3944
R5774 VDD.n3943 VDD.n3942 19.3944
R5775 VDD.n3942 VDD.n146 19.3944
R5776 VDD.n3936 VDD.n146 19.3944
R5777 VDD.n3899 VDD.n3898 19.3944
R5778 VDD.n3898 VDD.n3897 19.3944
R5779 VDD.n3897 VDD.n184 19.3944
R5780 VDD.n3891 VDD.n184 19.3944
R5781 VDD.n3891 VDD.n3890 19.3944
R5782 VDD.n3890 VDD.n3889 19.3944
R5783 VDD.n3889 VDD.n190 19.3944
R5784 VDD.n3883 VDD.n190 19.3944
R5785 VDD.n3883 VDD.n3882 19.3944
R5786 VDD.n3882 VDD.n3881 19.3944
R5787 VDD.n3881 VDD.n196 19.3944
R5788 VDD.n3875 VDD.n196 19.3944
R5789 VDD.n3875 VDD.n3874 19.3944
R5790 VDD.n3874 VDD.n3873 19.3944
R5791 VDD.n3873 VDD.n202 19.3944
R5792 VDD.n3867 VDD.n202 19.3944
R5793 VDD.n3934 VDD.n3933 19.3944
R5794 VDD.n3933 VDD.n154 19.3944
R5795 VDD.n3927 VDD.n154 19.3944
R5796 VDD.n3927 VDD.n3926 19.3944
R5797 VDD.n3926 VDD.n3925 19.3944
R5798 VDD.n3925 VDD.n160 19.3944
R5799 VDD.n3919 VDD.n160 19.3944
R5800 VDD.n165 VDD.n162 19.3944
R5801 VDD.n3914 VDD.n3913 19.3944
R5802 VDD.n3913 VDD.n169 19.3944
R5803 VDD.n3907 VDD.n169 19.3944
R5804 VDD.n3907 VDD.n3906 19.3944
R5805 VDD.n3906 VDD.n3905 19.3944
R5806 VDD.n3905 VDD.n175 19.3944
R5807 VDD.n3866 VDD.n3865 19.3944
R5808 VDD.n3865 VDD.n210 19.3944
R5809 VDD.n3859 VDD.n210 19.3944
R5810 VDD.n3859 VDD.n3858 19.3944
R5811 VDD.n3858 VDD.n3857 19.3944
R5812 VDD.n3857 VDD.n216 19.3944
R5813 VDD.n3851 VDD.n216 19.3944
R5814 VDD.n3851 VDD.n3850 19.3944
R5815 VDD.n3850 VDD.n3849 19.3944
R5816 VDD.n3845 VDD.n3844 19.3944
R5817 VDD.n3841 VDD.n3840 19.3944
R5818 VDD.n3840 VDD.n3764 19.3944
R5819 VDD.n3835 VDD.n3764 19.3944
R5820 VDD.n1588 VDD.n1519 18.8126
R5821 VDD.n2203 VDD.n1166 18.8126
R5822 VDD.n4416 VDD.n4284 18.8126
R5823 VDD.n3835 VDD.n3834 18.8126
R5824 VDD.n1559 VDD.n1558 18.2308
R5825 VDD.n2175 VDD.n1186 18.2308
R5826 VDD.n3800 VDD.n3797 18.2308
R5827 VDD.n4386 VDD.n4385 18.2308
R5828 VDD.n2463 VDD.n974 14.977
R5829 VDD.n2895 VDD.n602 14.977
R5830 VDD.n3335 VDD.n2896 14.977
R5831 VDD.n3743 VDD.n228 14.977
R5832 VDD.n27 VDD.t20 12.8483
R5833 VDD.n27 VDD.t164 12.8483
R5834 VDD.n24 VDD.t23 12.8483
R5835 VDD.n24 VDD.t7 12.8483
R5836 VDD.n21 VDD.t16 12.8483
R5837 VDD.n21 VDD.t162 12.8483
R5838 VDD.n18 VDD.t5 12.8483
R5839 VDD.n18 VDD.t13 12.8483
R5840 VDD.n16 VDD.t22 12.8483
R5841 VDD.n16 VDD.t168 12.8483
R5842 VDD.n1830 VDD.t24 12.8483
R5843 VDD.n1830 VDD.t165 12.8483
R5844 VDD.n1827 VDD.t25 12.8483
R5845 VDD.n1827 VDD.t161 12.8483
R5846 VDD.n1824 VDD.t15 12.8483
R5847 VDD.n1824 VDD.t1 12.8483
R5848 VDD.n1821 VDD.t17 12.8483
R5849 VDD.n1821 VDD.t26 12.8483
R5850 VDD.n1819 VDD.t12 12.8483
R5851 VDD.n1819 VDD.t167 12.8483
R5852 VDD.n2121 VDD.n999 10.7146
R5853 VDD.n3917 VDD.n164 10.7146
R5854 VDD.n3762 VDD.n3761 10.7146
R5855 VDD.n2208 VDD.n2207 10.7146
R5856 VDD.n1696 VDD.n1384 10.6221
R5857 VDD.n1704 VDD.n1384 10.6221
R5858 VDD.n1704 VDD.n1377 10.6221
R5859 VDD.n1712 VDD.n1377 10.6221
R5860 VDD.n1712 VDD.n1378 10.6221
R5861 VDD.n1720 VDD.n1366 10.6221
R5862 VDD.n1728 VDD.n1366 10.6221
R5863 VDD.n1728 VDD.n1360 10.6221
R5864 VDD.n1736 VDD.n1360 10.6221
R5865 VDD.n1736 VDD.n1354 10.6221
R5866 VDD.n1744 VDD.n1354 10.6221
R5867 VDD.n1744 VDD.n1348 10.6221
R5868 VDD.n1752 VDD.n1348 10.6221
R5869 VDD.n1752 VDD.n1342 10.6221
R5870 VDD.n1760 VDD.n1342 10.6221
R5871 VDD.n1760 VDD.n1336 10.6221
R5872 VDD.n1769 VDD.n1336 10.6221
R5873 VDD.n1769 VDD.n1768 10.6221
R5874 VDD.n1777 VDD.n1325 10.6221
R5875 VDD.n1785 VDD.n1325 10.6221
R5876 VDD.n1785 VDD.n1319 10.6221
R5877 VDD.n1793 VDD.n1319 10.6221
R5878 VDD.n1793 VDD.n1313 10.6221
R5879 VDD.n1801 VDD.n1313 10.6221
R5880 VDD.n1801 VDD.n1307 10.6221
R5881 VDD.n1809 VDD.n1307 10.6221
R5882 VDD.n1809 VDD.n1301 10.6221
R5883 VDD.t0 VDD.n1301 10.6221
R5884 VDD.t0 VDD.n1295 10.6221
R5885 VDD.n1839 VDD.n1295 10.6221
R5886 VDD.n1839 VDD.n1289 10.6221
R5887 VDD.n1847 VDD.n1289 10.6221
R5888 VDD.n1847 VDD.n1283 10.6221
R5889 VDD.n1855 VDD.n1283 10.6221
R5890 VDD.n1855 VDD.n1277 10.6221
R5891 VDD.n1863 VDD.n1277 10.6221
R5892 VDD.n1863 VDD.n1271 10.6221
R5893 VDD.n1871 VDD.n1271 10.6221
R5894 VDD.n1879 VDD.n1265 10.6221
R5895 VDD.n1879 VDD.n1259 10.6221
R5896 VDD.n1887 VDD.n1259 10.6221
R5897 VDD.n1887 VDD.n1253 10.6221
R5898 VDD.n1895 VDD.n1253 10.6221
R5899 VDD.n1895 VDD.n1247 10.6221
R5900 VDD.n1903 VDD.n1247 10.6221
R5901 VDD.n1903 VDD.n1241 10.6221
R5902 VDD.n1911 VDD.n1241 10.6221
R5903 VDD.n1911 VDD.n1235 10.6221
R5904 VDD.n1919 VDD.n1235 10.6221
R5905 VDD.n1919 VDD.n1229 10.6221
R5906 VDD.n1927 VDD.n1229 10.6221
R5907 VDD.n1935 VDD.n1223 10.6221
R5908 VDD.n1935 VDD.n1216 10.6221
R5909 VDD.n1945 VDD.n1216 10.6221
R5910 VDD.n1945 VDD.n1209 10.6221
R5911 VDD.n2170 VDD.n1209 10.6221
R5912 VDD.n3969 VDD.n121 10.6221
R5913 VDD.n3977 VDD.n121 10.6221
R5914 VDD.n3977 VDD.n114 10.6221
R5915 VDD.n3985 VDD.n114 10.6221
R5916 VDD.n3985 VDD.n115 10.6221
R5917 VDD.n3993 VDD.n103 10.6221
R5918 VDD.n4001 VDD.n103 10.6221
R5919 VDD.n4001 VDD.n97 10.6221
R5920 VDD.n4009 VDD.n97 10.6221
R5921 VDD.n4009 VDD.n91 10.6221
R5922 VDD.n4017 VDD.n91 10.6221
R5923 VDD.n4017 VDD.n85 10.6221
R5924 VDD.n4025 VDD.n85 10.6221
R5925 VDD.n4025 VDD.n79 10.6221
R5926 VDD.n4033 VDD.n79 10.6221
R5927 VDD.n4033 VDD.n73 10.6221
R5928 VDD.n4042 VDD.n73 10.6221
R5929 VDD.n4042 VDD.n4041 10.6221
R5930 VDD.n4050 VDD.n62 10.6221
R5931 VDD.n4058 VDD.n62 10.6221
R5932 VDD.n4058 VDD.n56 10.6221
R5933 VDD.n4066 VDD.n56 10.6221
R5934 VDD.n4066 VDD.n50 10.6221
R5935 VDD.n4074 VDD.n50 10.6221
R5936 VDD.n4074 VDD.n44 10.6221
R5937 VDD.n4082 VDD.n44 10.6221
R5938 VDD.n4082 VDD.n36 10.6221
R5939 VDD.t6 VDD.n36 10.6221
R5940 VDD.t6 VDD.n37 10.6221
R5941 VDD.n4596 VDD.n37 10.6221
R5942 VDD.n4596 VDD.n4092 10.6221
R5943 VDD.n4590 VDD.n4092 10.6221
R5944 VDD.n4590 VDD.n4589 10.6221
R5945 VDD.n4589 VDD.n4588 10.6221
R5946 VDD.n4588 VDD.n4102 10.6221
R5947 VDD.n4582 VDD.n4102 10.6221
R5948 VDD.n4582 VDD.n4581 10.6221
R5949 VDD.n4581 VDD.n4580 10.6221
R5950 VDD.n4574 VDD.n4120 10.6221
R5951 VDD.n4574 VDD.n4573 10.6221
R5952 VDD.n4573 VDD.n4572 10.6221
R5953 VDD.n4572 VDD.n4124 10.6221
R5954 VDD.n4566 VDD.n4124 10.6221
R5955 VDD.n4566 VDD.n4565 10.6221
R5956 VDD.n4565 VDD.n4564 10.6221
R5957 VDD.n4564 VDD.n4135 10.6221
R5958 VDD.n4558 VDD.n4135 10.6221
R5959 VDD.n4558 VDD.n4557 10.6221
R5960 VDD.n4557 VDD.n4556 10.6221
R5961 VDD.n4556 VDD.n4146 10.6221
R5962 VDD.n4550 VDD.n4146 10.6221
R5963 VDD.n4549 VDD.n4548 10.6221
R5964 VDD.n4548 VDD.n4157 10.6221
R5965 VDD.n4542 VDD.n4157 10.6221
R5966 VDD.n4542 VDD.n4541 10.6221
R5967 VDD.n4541 VDD.n4540 10.6221
R5968 VDD.n2853 VDD.n2851 10.6151
R5969 VDD.n2851 VDD.n2848 10.6151
R5970 VDD.n2848 VDD.n2847 10.6151
R5971 VDD.n2847 VDD.n2844 10.6151
R5972 VDD.n2844 VDD.n2843 10.6151
R5973 VDD.n2843 VDD.n2840 10.6151
R5974 VDD.n2840 VDD.n2839 10.6151
R5975 VDD.n2839 VDD.n2836 10.6151
R5976 VDD.n2836 VDD.n2835 10.6151
R5977 VDD.n2835 VDD.n2832 10.6151
R5978 VDD.n2832 VDD.n2831 10.6151
R5979 VDD.n2831 VDD.n2828 10.6151
R5980 VDD.n2828 VDD.n2827 10.6151
R5981 VDD.n2827 VDD.n2824 10.6151
R5982 VDD.n2824 VDD.n2823 10.6151
R5983 VDD.n2823 VDD.n2820 10.6151
R5984 VDD.n2820 VDD.n2819 10.6151
R5985 VDD.n2432 VDD.n2430 10.6151
R5986 VDD.n2430 VDD.n2429 10.6151
R5987 VDD.n2429 VDD.n2427 10.6151
R5988 VDD.n2427 VDD.n2426 10.6151
R5989 VDD.n2426 VDD.n2424 10.6151
R5990 VDD.n2424 VDD.n2423 10.6151
R5991 VDD.n2423 VDD.n2421 10.6151
R5992 VDD.n2421 VDD.n2420 10.6151
R5993 VDD.n2420 VDD.n2418 10.6151
R5994 VDD.n2418 VDD.n2417 10.6151
R5995 VDD.n2417 VDD.n1153 10.6151
R5996 VDD.n1153 VDD.n1152 10.6151
R5997 VDD.n1152 VDD.n1150 10.6151
R5998 VDD.n1150 VDD.n1149 10.6151
R5999 VDD.n1149 VDD.n1147 10.6151
R6000 VDD.n1147 VDD.n1146 10.6151
R6001 VDD.n1146 VDD.n1144 10.6151
R6002 VDD.n1144 VDD.n1143 10.6151
R6003 VDD.n1143 VDD.n1141 10.6151
R6004 VDD.n1141 VDD.n1140 10.6151
R6005 VDD.n1140 VDD.n1138 10.6151
R6006 VDD.n1138 VDD.n1137 10.6151
R6007 VDD.n1137 VDD.n1135 10.6151
R6008 VDD.n1135 VDD.n1134 10.6151
R6009 VDD.n1134 VDD.n1132 10.6151
R6010 VDD.n1132 VDD.n1131 10.6151
R6011 VDD.n1131 VDD.n1129 10.6151
R6012 VDD.n1129 VDD.n1128 10.6151
R6013 VDD.n1128 VDD.n1126 10.6151
R6014 VDD.n1126 VDD.n1125 10.6151
R6015 VDD.n1125 VDD.n1123 10.6151
R6016 VDD.n1123 VDD.n1122 10.6151
R6017 VDD.n1122 VDD.n1120 10.6151
R6018 VDD.n1120 VDD.n1119 10.6151
R6019 VDD.n1119 VDD.n1117 10.6151
R6020 VDD.n1117 VDD.n1116 10.6151
R6021 VDD.n1116 VDD.n1114 10.6151
R6022 VDD.n1114 VDD.n1113 10.6151
R6023 VDD.n1113 VDD.n1111 10.6151
R6024 VDD.n1111 VDD.n1110 10.6151
R6025 VDD.n1110 VDD.n1108 10.6151
R6026 VDD.n1108 VDD.n1107 10.6151
R6027 VDD.n1107 VDD.n1105 10.6151
R6028 VDD.n1105 VDD.n1104 10.6151
R6029 VDD.n1104 VDD.n1102 10.6151
R6030 VDD.n1102 VDD.n1101 10.6151
R6031 VDD.n1101 VDD.n1099 10.6151
R6032 VDD.n1099 VDD.n1098 10.6151
R6033 VDD.n1098 VDD.n1096 10.6151
R6034 VDD.n1096 VDD.n1095 10.6151
R6035 VDD.n1095 VDD.n1093 10.6151
R6036 VDD.n1093 VDD.n1092 10.6151
R6037 VDD.n1092 VDD.n1090 10.6151
R6038 VDD.n1090 VDD.n1089 10.6151
R6039 VDD.n1089 VDD.n1087 10.6151
R6040 VDD.n1087 VDD.n1086 10.6151
R6041 VDD.n1086 VDD.n1084 10.6151
R6042 VDD.n1084 VDD.n1083 10.6151
R6043 VDD.n1083 VDD.n1081 10.6151
R6044 VDD.n1081 VDD.n1080 10.6151
R6045 VDD.n1080 VDD.n1078 10.6151
R6046 VDD.n1078 VDD.n1077 10.6151
R6047 VDD.n1077 VDD.n1075 10.6151
R6048 VDD.n1075 VDD.n1074 10.6151
R6049 VDD.n1074 VDD.n1072 10.6151
R6050 VDD.n1072 VDD.n1071 10.6151
R6051 VDD.n1071 VDD.n1069 10.6151
R6052 VDD.n1069 VDD.n1068 10.6151
R6053 VDD.n1068 VDD.n1066 10.6151
R6054 VDD.n1066 VDD.n1065 10.6151
R6055 VDD.n1065 VDD.n1063 10.6151
R6056 VDD.n1063 VDD.n1062 10.6151
R6057 VDD.n1062 VDD.n1060 10.6151
R6058 VDD.n1060 VDD.n1059 10.6151
R6059 VDD.n1059 VDD.n1057 10.6151
R6060 VDD.n1057 VDD.n1056 10.6151
R6061 VDD.n1056 VDD.n1054 10.6151
R6062 VDD.n1054 VDD.n1053 10.6151
R6063 VDD.n1053 VDD.n1051 10.6151
R6064 VDD.n1051 VDD.n1050 10.6151
R6065 VDD.n1050 VDD.n1048 10.6151
R6066 VDD.n1048 VDD.n1047 10.6151
R6067 VDD.n1047 VDD.n1045 10.6151
R6068 VDD.n1045 VDD.n1044 10.6151
R6069 VDD.n1044 VDD.n1042 10.6151
R6070 VDD.n1042 VDD.n1041 10.6151
R6071 VDD.n1041 VDD.n1039 10.6151
R6072 VDD.n1039 VDD.n1038 10.6151
R6073 VDD.n1038 VDD.n1036 10.6151
R6074 VDD.n1036 VDD.n1035 10.6151
R6075 VDD.n1035 VDD.n1033 10.6151
R6076 VDD.n1033 VDD.n1032 10.6151
R6077 VDD.n1032 VDD.n1030 10.6151
R6078 VDD.n1030 VDD.n1029 10.6151
R6079 VDD.n1029 VDD.n1027 10.6151
R6080 VDD.n1027 VDD.n1026 10.6151
R6081 VDD.n1026 VDD.n1024 10.6151
R6082 VDD.n1024 VDD.n1023 10.6151
R6083 VDD.n1023 VDD.n1021 10.6151
R6084 VDD.n1021 VDD.n1020 10.6151
R6085 VDD.n1020 VDD.n1018 10.6151
R6086 VDD.n1018 VDD.n1017 10.6151
R6087 VDD.n1017 VDD.n1015 10.6151
R6088 VDD.n1015 VDD.n1014 10.6151
R6089 VDD.n1014 VDD.n1012 10.6151
R6090 VDD.n1012 VDD.n1011 10.6151
R6091 VDD.n1011 VDD.n1009 10.6151
R6092 VDD.n1009 VDD.n1008 10.6151
R6093 VDD.n1008 VDD.n1006 10.6151
R6094 VDD.n1006 VDD.n1005 10.6151
R6095 VDD.n1005 VDD.n1003 10.6151
R6096 VDD.n1003 VDD.n1002 10.6151
R6097 VDD.n1002 VDD.n636 10.6151
R6098 VDD.n2814 VDD.n636 10.6151
R6099 VDD.n2815 VDD.n2814 10.6151
R6100 VDD.n2816 VDD.n2815 10.6151
R6101 VDD.n2466 VDD.n978 10.6151
R6102 VDD.n2461 VDD.n978 10.6151
R6103 VDD.n2461 VDD.n2460 10.6151
R6104 VDD.n2460 VDD.n2459 10.6151
R6105 VDD.n2459 VDD.n2456 10.6151
R6106 VDD.n2456 VDD.n2455 10.6151
R6107 VDD.n2455 VDD.n2452 10.6151
R6108 VDD.n2452 VDD.n2451 10.6151
R6109 VDD.n2448 VDD.n2447 10.6151
R6110 VDD.n2447 VDD.n2444 10.6151
R6111 VDD.n2444 VDD.n2443 10.6151
R6112 VDD.n2443 VDD.n2440 10.6151
R6113 VDD.n2440 VDD.n2439 10.6151
R6114 VDD.n2439 VDD.n2436 10.6151
R6115 VDD.n2436 VDD.n2435 10.6151
R6116 VDD.n2435 VDD.n2433 10.6151
R6117 VDD.n2468 VDD.n2467 10.6151
R6118 VDD.n2468 VDD.n966 10.6151
R6119 VDD.n2478 VDD.n966 10.6151
R6120 VDD.n2479 VDD.n2478 10.6151
R6121 VDD.n2480 VDD.n2479 10.6151
R6122 VDD.n2480 VDD.n954 10.6151
R6123 VDD.n2490 VDD.n954 10.6151
R6124 VDD.n2491 VDD.n2490 10.6151
R6125 VDD.n2492 VDD.n2491 10.6151
R6126 VDD.n2492 VDD.n943 10.6151
R6127 VDD.n2502 VDD.n943 10.6151
R6128 VDD.n2503 VDD.n2502 10.6151
R6129 VDD.n2504 VDD.n2503 10.6151
R6130 VDD.n2504 VDD.n931 10.6151
R6131 VDD.n2514 VDD.n931 10.6151
R6132 VDD.n2515 VDD.n2514 10.6151
R6133 VDD.n2516 VDD.n2515 10.6151
R6134 VDD.n2516 VDD.n919 10.6151
R6135 VDD.n2526 VDD.n919 10.6151
R6136 VDD.n2527 VDD.n2526 10.6151
R6137 VDD.n2528 VDD.n2527 10.6151
R6138 VDD.n2528 VDD.n907 10.6151
R6139 VDD.n2538 VDD.n907 10.6151
R6140 VDD.n2539 VDD.n2538 10.6151
R6141 VDD.n2540 VDD.n2539 10.6151
R6142 VDD.n2540 VDD.n895 10.6151
R6143 VDD.n2550 VDD.n895 10.6151
R6144 VDD.n2551 VDD.n2550 10.6151
R6145 VDD.n2552 VDD.n2551 10.6151
R6146 VDD.n2552 VDD.n883 10.6151
R6147 VDD.n2562 VDD.n883 10.6151
R6148 VDD.n2563 VDD.n2562 10.6151
R6149 VDD.n2564 VDD.n2563 10.6151
R6150 VDD.n2564 VDD.n871 10.6151
R6151 VDD.n2574 VDD.n871 10.6151
R6152 VDD.n2575 VDD.n2574 10.6151
R6153 VDD.n2576 VDD.n2575 10.6151
R6154 VDD.n2576 VDD.n859 10.6151
R6155 VDD.n2586 VDD.n859 10.6151
R6156 VDD.n2587 VDD.n2586 10.6151
R6157 VDD.n2588 VDD.n2587 10.6151
R6158 VDD.n2588 VDD.n847 10.6151
R6159 VDD.n2598 VDD.n847 10.6151
R6160 VDD.n2599 VDD.n2598 10.6151
R6161 VDD.n2600 VDD.n2599 10.6151
R6162 VDD.n2600 VDD.n835 10.6151
R6163 VDD.n2610 VDD.n835 10.6151
R6164 VDD.n2611 VDD.n2610 10.6151
R6165 VDD.n2612 VDD.n2611 10.6151
R6166 VDD.n2612 VDD.n822 10.6151
R6167 VDD.n2622 VDD.n822 10.6151
R6168 VDD.n2623 VDD.n2622 10.6151
R6169 VDD.n2624 VDD.n2623 10.6151
R6170 VDD.n2624 VDD.n811 10.6151
R6171 VDD.n2634 VDD.n811 10.6151
R6172 VDD.n2635 VDD.n2634 10.6151
R6173 VDD.n2636 VDD.n2635 10.6151
R6174 VDD.n2636 VDD.n799 10.6151
R6175 VDD.n2646 VDD.n799 10.6151
R6176 VDD.n2647 VDD.n2646 10.6151
R6177 VDD.n2648 VDD.n2647 10.6151
R6178 VDD.n2648 VDD.n787 10.6151
R6179 VDD.n2658 VDD.n787 10.6151
R6180 VDD.n2659 VDD.n2658 10.6151
R6181 VDD.n2660 VDD.n2659 10.6151
R6182 VDD.n2660 VDD.n775 10.6151
R6183 VDD.n2670 VDD.n775 10.6151
R6184 VDD.n2671 VDD.n2670 10.6151
R6185 VDD.n2672 VDD.n2671 10.6151
R6186 VDD.n2672 VDD.n763 10.6151
R6187 VDD.n2682 VDD.n763 10.6151
R6188 VDD.n2683 VDD.n2682 10.6151
R6189 VDD.n2684 VDD.n2683 10.6151
R6190 VDD.n2684 VDD.n751 10.6151
R6191 VDD.n2694 VDD.n751 10.6151
R6192 VDD.n2695 VDD.n2694 10.6151
R6193 VDD.n2696 VDD.n2695 10.6151
R6194 VDD.n2696 VDD.n739 10.6151
R6195 VDD.n2706 VDD.n739 10.6151
R6196 VDD.n2707 VDD.n2706 10.6151
R6197 VDD.n2708 VDD.n2707 10.6151
R6198 VDD.n2708 VDD.n726 10.6151
R6199 VDD.n2718 VDD.n726 10.6151
R6200 VDD.n2719 VDD.n2718 10.6151
R6201 VDD.n2720 VDD.n2719 10.6151
R6202 VDD.n2720 VDD.n715 10.6151
R6203 VDD.n2730 VDD.n715 10.6151
R6204 VDD.n2731 VDD.n2730 10.6151
R6205 VDD.n2732 VDD.n2731 10.6151
R6206 VDD.n2732 VDD.n703 10.6151
R6207 VDD.n2742 VDD.n703 10.6151
R6208 VDD.n2743 VDD.n2742 10.6151
R6209 VDD.n2744 VDD.n2743 10.6151
R6210 VDD.n2744 VDD.n691 10.6151
R6211 VDD.n2754 VDD.n691 10.6151
R6212 VDD.n2755 VDD.n2754 10.6151
R6213 VDD.n2756 VDD.n2755 10.6151
R6214 VDD.n2756 VDD.n679 10.6151
R6215 VDD.n2766 VDD.n679 10.6151
R6216 VDD.n2767 VDD.n2766 10.6151
R6217 VDD.n2768 VDD.n2767 10.6151
R6218 VDD.n2768 VDD.n667 10.6151
R6219 VDD.n2778 VDD.n667 10.6151
R6220 VDD.n2779 VDD.n2778 10.6151
R6221 VDD.n2780 VDD.n2779 10.6151
R6222 VDD.n2780 VDD.n655 10.6151
R6223 VDD.n2790 VDD.n655 10.6151
R6224 VDD.n2791 VDD.n2790 10.6151
R6225 VDD.n2792 VDD.n2791 10.6151
R6226 VDD.n2792 VDD.n642 10.6151
R6227 VDD.n2807 VDD.n642 10.6151
R6228 VDD.n2808 VDD.n2807 10.6151
R6229 VDD.n2809 VDD.n2808 10.6151
R6230 VDD.n2809 VDD.n633 10.6151
R6231 VDD.n2855 VDD.n633 10.6151
R6232 VDD.n2855 VDD.n2854 10.6151
R6233 VDD.n3110 VDD.n3109 10.6151
R6234 VDD.n3109 VDD.n3108 10.6151
R6235 VDD.n3108 VDD.n3107 10.6151
R6236 VDD.n3107 VDD.n3105 10.6151
R6237 VDD.n3105 VDD.n3104 10.6151
R6238 VDD.n3104 VDD.n3102 10.6151
R6239 VDD.n3102 VDD.n3101 10.6151
R6240 VDD.n3101 VDD.n3099 10.6151
R6241 VDD.n3099 VDD.n3098 10.6151
R6242 VDD.n3098 VDD.n3096 10.6151
R6243 VDD.n3096 VDD.n3095 10.6151
R6244 VDD.n3095 VDD.n3093 10.6151
R6245 VDD.n3093 VDD.n3092 10.6151
R6246 VDD.n3092 VDD.n3090 10.6151
R6247 VDD.n3090 VDD.n3089 10.6151
R6248 VDD.n3089 VDD.n3087 10.6151
R6249 VDD.n3087 VDD.n3086 10.6151
R6250 VDD.n3086 VDD.n3084 10.6151
R6251 VDD.n3084 VDD.n3083 10.6151
R6252 VDD.n3083 VDD.n3081 10.6151
R6253 VDD.n3081 VDD.n3080 10.6151
R6254 VDD.n3080 VDD.n3078 10.6151
R6255 VDD.n3078 VDD.n3077 10.6151
R6256 VDD.n3077 VDD.n3075 10.6151
R6257 VDD.n3075 VDD.n3074 10.6151
R6258 VDD.n3074 VDD.n3072 10.6151
R6259 VDD.n3072 VDD.n3071 10.6151
R6260 VDD.n3071 VDD.n3069 10.6151
R6261 VDD.n3069 VDD.n3068 10.6151
R6262 VDD.n3068 VDD.n3066 10.6151
R6263 VDD.n3066 VDD.n3065 10.6151
R6264 VDD.n3065 VDD.n3063 10.6151
R6265 VDD.n3063 VDD.n3062 10.6151
R6266 VDD.n3062 VDD.n3060 10.6151
R6267 VDD.n3060 VDD.n3059 10.6151
R6268 VDD.n3059 VDD.n3057 10.6151
R6269 VDD.n3057 VDD.n3056 10.6151
R6270 VDD.n3056 VDD.n3054 10.6151
R6271 VDD.n3054 VDD.n3053 10.6151
R6272 VDD.n3053 VDD.n3051 10.6151
R6273 VDD.n3051 VDD.n3050 10.6151
R6274 VDD.n3050 VDD.n3048 10.6151
R6275 VDD.n3048 VDD.n3047 10.6151
R6276 VDD.n3047 VDD.n3045 10.6151
R6277 VDD.n3045 VDD.n3044 10.6151
R6278 VDD.n3044 VDD.n3042 10.6151
R6279 VDD.n3042 VDD.n3041 10.6151
R6280 VDD.n3041 VDD.n3039 10.6151
R6281 VDD.n3039 VDD.n3038 10.6151
R6282 VDD.n3038 VDD.n3036 10.6151
R6283 VDD.n3036 VDD.n3035 10.6151
R6284 VDD.n3035 VDD.n3033 10.6151
R6285 VDD.n3033 VDD.n3032 10.6151
R6286 VDD.n3032 VDD.n3030 10.6151
R6287 VDD.n3030 VDD.n3029 10.6151
R6288 VDD.n3029 VDD.n3027 10.6151
R6289 VDD.n3027 VDD.n3026 10.6151
R6290 VDD.n3026 VDD.n3024 10.6151
R6291 VDD.n3024 VDD.n3023 10.6151
R6292 VDD.n3023 VDD.n3021 10.6151
R6293 VDD.n3021 VDD.n3020 10.6151
R6294 VDD.n3020 VDD.n3018 10.6151
R6295 VDD.n3018 VDD.n3017 10.6151
R6296 VDD.n3017 VDD.n3015 10.6151
R6297 VDD.n3015 VDD.n3014 10.6151
R6298 VDD.n3014 VDD.n3012 10.6151
R6299 VDD.n3012 VDD.n3011 10.6151
R6300 VDD.n3011 VDD.n3009 10.6151
R6301 VDD.n3009 VDD.n3008 10.6151
R6302 VDD.n3008 VDD.n3006 10.6151
R6303 VDD.n3006 VDD.n3005 10.6151
R6304 VDD.n3005 VDD.n3003 10.6151
R6305 VDD.n3003 VDD.n3002 10.6151
R6306 VDD.n3002 VDD.n3000 10.6151
R6307 VDD.n3000 VDD.n2999 10.6151
R6308 VDD.n2999 VDD.n2997 10.6151
R6309 VDD.n2997 VDD.n2996 10.6151
R6310 VDD.n2996 VDD.n2994 10.6151
R6311 VDD.n2994 VDD.n2993 10.6151
R6312 VDD.n2993 VDD.n2991 10.6151
R6313 VDD.n2991 VDD.n2990 10.6151
R6314 VDD.n2990 VDD.n2988 10.6151
R6315 VDD.n2988 VDD.n2987 10.6151
R6316 VDD.n2987 VDD.n2985 10.6151
R6317 VDD.n2985 VDD.n2984 10.6151
R6318 VDD.n2984 VDD.n2982 10.6151
R6319 VDD.n2982 VDD.n2981 10.6151
R6320 VDD.n2981 VDD.n2979 10.6151
R6321 VDD.n2979 VDD.n2978 10.6151
R6322 VDD.n2978 VDD.n2976 10.6151
R6323 VDD.n2976 VDD.n2975 10.6151
R6324 VDD.n2975 VDD.n2973 10.6151
R6325 VDD.n2973 VDD.n2972 10.6151
R6326 VDD.n2972 VDD.n2970 10.6151
R6327 VDD.n2970 VDD.n2969 10.6151
R6328 VDD.n2969 VDD.n2967 10.6151
R6329 VDD.n2967 VDD.n2966 10.6151
R6330 VDD.n2966 VDD.n2964 10.6151
R6331 VDD.n2964 VDD.n2963 10.6151
R6332 VDD.n2963 VDD.n2961 10.6151
R6333 VDD.n2961 VDD.n2960 10.6151
R6334 VDD.n2960 VDD.n2958 10.6151
R6335 VDD.n2958 VDD.n2957 10.6151
R6336 VDD.n2957 VDD.n2955 10.6151
R6337 VDD.n2955 VDD.n2954 10.6151
R6338 VDD.n2954 VDD.n2952 10.6151
R6339 VDD.n2952 VDD.n2951 10.6151
R6340 VDD.n2951 VDD.n2949 10.6151
R6341 VDD.n2949 VDD.n2948 10.6151
R6342 VDD.n2948 VDD.n2946 10.6151
R6343 VDD.n2946 VDD.n2945 10.6151
R6344 VDD.n2945 VDD.n2943 10.6151
R6345 VDD.n2943 VDD.n2942 10.6151
R6346 VDD.n2942 VDD.n257 10.6151
R6347 VDD.n3706 VDD.n257 10.6151
R6348 VDD.n3707 VDD.n3706 10.6151
R6349 VDD.n2909 VDD.n600 10.6151
R6350 VDD.n2909 VDD.n2908 10.6151
R6351 VDD.n2915 VDD.n2908 10.6151
R6352 VDD.n2916 VDD.n2915 10.6151
R6353 VDD.n2917 VDD.n2916 10.6151
R6354 VDD.n2917 VDD.n2906 10.6151
R6355 VDD.n2923 VDD.n2906 10.6151
R6356 VDD.n2924 VDD.n2923 10.6151
R6357 VDD.n2925 VDD.n2924 10.6151
R6358 VDD.n2925 VDD.n2904 10.6151
R6359 VDD.n2931 VDD.n2904 10.6151
R6360 VDD.n2932 VDD.n2931 10.6151
R6361 VDD.n2933 VDD.n2932 10.6151
R6362 VDD.n2933 VDD.n2902 10.6151
R6363 VDD.n2902 VDD.n2899 10.6151
R6364 VDD.n2940 VDD.n2899 10.6151
R6365 VDD.n2941 VDD.n2940 10.6151
R6366 VDD.n3338 VDD.n3337 10.6151
R6367 VDD.n3339 VDD.n3338 10.6151
R6368 VDD.n3339 VDD.n588 10.6151
R6369 VDD.n3349 VDD.n588 10.6151
R6370 VDD.n3350 VDD.n3349 10.6151
R6371 VDD.n3351 VDD.n3350 10.6151
R6372 VDD.n3351 VDD.n576 10.6151
R6373 VDD.n3361 VDD.n576 10.6151
R6374 VDD.n3362 VDD.n3361 10.6151
R6375 VDD.n3363 VDD.n3362 10.6151
R6376 VDD.n3363 VDD.n564 10.6151
R6377 VDD.n3373 VDD.n564 10.6151
R6378 VDD.n3374 VDD.n3373 10.6151
R6379 VDD.n3375 VDD.n3374 10.6151
R6380 VDD.n3375 VDD.n552 10.6151
R6381 VDD.n3385 VDD.n552 10.6151
R6382 VDD.n3386 VDD.n3385 10.6151
R6383 VDD.n3387 VDD.n3386 10.6151
R6384 VDD.n3387 VDD.n540 10.6151
R6385 VDD.n3397 VDD.n540 10.6151
R6386 VDD.n3398 VDD.n3397 10.6151
R6387 VDD.n3399 VDD.n3398 10.6151
R6388 VDD.n3399 VDD.n528 10.6151
R6389 VDD.n3409 VDD.n528 10.6151
R6390 VDD.n3410 VDD.n3409 10.6151
R6391 VDD.n3411 VDD.n3410 10.6151
R6392 VDD.n3411 VDD.n516 10.6151
R6393 VDD.n3421 VDD.n516 10.6151
R6394 VDD.n3422 VDD.n3421 10.6151
R6395 VDD.n3423 VDD.n3422 10.6151
R6396 VDD.n3423 VDD.n504 10.6151
R6397 VDD.n3433 VDD.n504 10.6151
R6398 VDD.n3434 VDD.n3433 10.6151
R6399 VDD.n3435 VDD.n3434 10.6151
R6400 VDD.n3435 VDD.n492 10.6151
R6401 VDD.n3445 VDD.n492 10.6151
R6402 VDD.n3446 VDD.n3445 10.6151
R6403 VDD.n3447 VDD.n3446 10.6151
R6404 VDD.n3447 VDD.n480 10.6151
R6405 VDD.n3457 VDD.n480 10.6151
R6406 VDD.n3458 VDD.n3457 10.6151
R6407 VDD.n3459 VDD.n3458 10.6151
R6408 VDD.n3459 VDD.n467 10.6151
R6409 VDD.n3469 VDD.n467 10.6151
R6410 VDD.n3470 VDD.n3469 10.6151
R6411 VDD.n3471 VDD.n3470 10.6151
R6412 VDD.n3471 VDD.n455 10.6151
R6413 VDD.n3481 VDD.n455 10.6151
R6414 VDD.n3482 VDD.n3481 10.6151
R6415 VDD.n3483 VDD.n3482 10.6151
R6416 VDD.n3483 VDD.n444 10.6151
R6417 VDD.n3493 VDD.n444 10.6151
R6418 VDD.n3494 VDD.n3493 10.6151
R6419 VDD.n3495 VDD.n3494 10.6151
R6420 VDD.n3495 VDD.n432 10.6151
R6421 VDD.n3505 VDD.n432 10.6151
R6422 VDD.n3506 VDD.n3505 10.6151
R6423 VDD.n3507 VDD.n3506 10.6151
R6424 VDD.n3507 VDD.n420 10.6151
R6425 VDD.n3517 VDD.n420 10.6151
R6426 VDD.n3518 VDD.n3517 10.6151
R6427 VDD.n3519 VDD.n3518 10.6151
R6428 VDD.n3519 VDD.n408 10.6151
R6429 VDD.n3529 VDD.n408 10.6151
R6430 VDD.n3530 VDD.n3529 10.6151
R6431 VDD.n3531 VDD.n3530 10.6151
R6432 VDD.n3531 VDD.n396 10.6151
R6433 VDD.n3541 VDD.n396 10.6151
R6434 VDD.n3542 VDD.n3541 10.6151
R6435 VDD.n3543 VDD.n3542 10.6151
R6436 VDD.n3543 VDD.n384 10.6151
R6437 VDD.n3553 VDD.n384 10.6151
R6438 VDD.n3554 VDD.n3553 10.6151
R6439 VDD.n3555 VDD.n3554 10.6151
R6440 VDD.n3555 VDD.n372 10.6151
R6441 VDD.n3565 VDD.n372 10.6151
R6442 VDD.n3566 VDD.n3565 10.6151
R6443 VDD.n3567 VDD.n3566 10.6151
R6444 VDD.n3567 VDD.n360 10.6151
R6445 VDD.n3577 VDD.n360 10.6151
R6446 VDD.n3578 VDD.n3577 10.6151
R6447 VDD.n3579 VDD.n3578 10.6151
R6448 VDD.n3579 VDD.n348 10.6151
R6449 VDD.n3589 VDD.n348 10.6151
R6450 VDD.n3590 VDD.n3589 10.6151
R6451 VDD.n3591 VDD.n3590 10.6151
R6452 VDD.n3591 VDD.n335 10.6151
R6453 VDD.n3601 VDD.n335 10.6151
R6454 VDD.n3602 VDD.n3601 10.6151
R6455 VDD.n3603 VDD.n3602 10.6151
R6456 VDD.n3603 VDD.n324 10.6151
R6457 VDD.n3613 VDD.n324 10.6151
R6458 VDD.n3614 VDD.n3613 10.6151
R6459 VDD.n3615 VDD.n3614 10.6151
R6460 VDD.n3615 VDD.n312 10.6151
R6461 VDD.n3625 VDD.n312 10.6151
R6462 VDD.n3626 VDD.n3625 10.6151
R6463 VDD.n3627 VDD.n3626 10.6151
R6464 VDD.n3627 VDD.n300 10.6151
R6465 VDD.n3637 VDD.n300 10.6151
R6466 VDD.n3638 VDD.n3637 10.6151
R6467 VDD.n3639 VDD.n3638 10.6151
R6468 VDD.n3639 VDD.n287 10.6151
R6469 VDD.n3649 VDD.n287 10.6151
R6470 VDD.n3650 VDD.n3649 10.6151
R6471 VDD.n3651 VDD.n3650 10.6151
R6472 VDD.n3651 VDD.n276 10.6151
R6473 VDD.n3661 VDD.n276 10.6151
R6474 VDD.n3662 VDD.n3661 10.6151
R6475 VDD.n3663 VDD.n3662 10.6151
R6476 VDD.n3663 VDD.n263 10.6151
R6477 VDD.n3699 VDD.n263 10.6151
R6478 VDD.n3700 VDD.n3699 10.6151
R6479 VDD.n3701 VDD.n3700 10.6151
R6480 VDD.n3701 VDD.n243 10.6151
R6481 VDD.n3741 VDD.n243 10.6151
R6482 VDD.n3740 VDD.n3739 10.6151
R6483 VDD.n3739 VDD.n244 10.6151
R6484 VDD.n3734 VDD.n244 10.6151
R6485 VDD.n3734 VDD.n3733 10.6151
R6486 VDD.n3733 VDD.n3732 10.6151
R6487 VDD.n3732 VDD.n247 10.6151
R6488 VDD.n3727 VDD.n247 10.6151
R6489 VDD.n3727 VDD.n3726 10.6151
R6490 VDD.n3722 VDD.n3721 10.6151
R6491 VDD.n3721 VDD.n3720 10.6151
R6492 VDD.n3720 VDD.n250 10.6151
R6493 VDD.n3715 VDD.n250 10.6151
R6494 VDD.n3715 VDD.n3714 10.6151
R6495 VDD.n3714 VDD.n3713 10.6151
R6496 VDD.n3713 VDD.n255 10.6151
R6497 VDD.n3708 VDD.n255 10.6151
R6498 VDD.n3689 VDD.n3669 10.6151
R6499 VDD.n3670 VDD.n3669 10.6151
R6500 VDD.n3682 VDD.n3670 10.6151
R6501 VDD.n3682 VDD.n3681 10.6151
R6502 VDD.n3681 VDD.n3680 10.6151
R6503 VDD.n3680 VDD.n3672 10.6151
R6504 VDD.n3675 VDD.n3672 10.6151
R6505 VDD.n3675 VDD.n225 10.6151
R6506 VDD.n3760 VDD.n226 10.6151
R6507 VDD.n3755 VDD.n226 10.6151
R6508 VDD.n3755 VDD.n3754 10.6151
R6509 VDD.n3754 VDD.n3753 10.6151
R6510 VDD.n3753 VDD.n232 10.6151
R6511 VDD.n3748 VDD.n232 10.6151
R6512 VDD.n3748 VDD.n3747 10.6151
R6513 VDD.n3747 VDD.n3746 10.6151
R6514 VDD.n3296 VDD.n3295 10.6151
R6515 VDD.n3295 VDD.n3293 10.6151
R6516 VDD.n3293 VDD.n3292 10.6151
R6517 VDD.n3292 VDD.n3290 10.6151
R6518 VDD.n3290 VDD.n3289 10.6151
R6519 VDD.n3289 VDD.n3287 10.6151
R6520 VDD.n3287 VDD.n3286 10.6151
R6521 VDD.n3286 VDD.n3284 10.6151
R6522 VDD.n3284 VDD.n3283 10.6151
R6523 VDD.n3283 VDD.n3281 10.6151
R6524 VDD.n3281 VDD.n3280 10.6151
R6525 VDD.n3280 VDD.n3278 10.6151
R6526 VDD.n3278 VDD.n3277 10.6151
R6527 VDD.n3277 VDD.n3275 10.6151
R6528 VDD.n3275 VDD.n3274 10.6151
R6529 VDD.n3274 VDD.n3272 10.6151
R6530 VDD.n3272 VDD.n3271 10.6151
R6531 VDD.n3271 VDD.n3269 10.6151
R6532 VDD.n3269 VDD.n3268 10.6151
R6533 VDD.n3268 VDD.n3266 10.6151
R6534 VDD.n3266 VDD.n3265 10.6151
R6535 VDD.n3265 VDD.n3263 10.6151
R6536 VDD.n3263 VDD.n3262 10.6151
R6537 VDD.n3262 VDD.n3260 10.6151
R6538 VDD.n3260 VDD.n3259 10.6151
R6539 VDD.n3259 VDD.n3257 10.6151
R6540 VDD.n3257 VDD.n3256 10.6151
R6541 VDD.n3256 VDD.n3254 10.6151
R6542 VDD.n3254 VDD.n3253 10.6151
R6543 VDD.n3253 VDD.n3251 10.6151
R6544 VDD.n3251 VDD.n3250 10.6151
R6545 VDD.n3250 VDD.n3248 10.6151
R6546 VDD.n3248 VDD.n3247 10.6151
R6547 VDD.n3247 VDD.n3245 10.6151
R6548 VDD.n3245 VDD.n3244 10.6151
R6549 VDD.n3244 VDD.n3242 10.6151
R6550 VDD.n3242 VDD.n3241 10.6151
R6551 VDD.n3241 VDD.n3239 10.6151
R6552 VDD.n3239 VDD.n3238 10.6151
R6553 VDD.n3238 VDD.n3236 10.6151
R6554 VDD.n3236 VDD.n3235 10.6151
R6555 VDD.n3235 VDD.n3233 10.6151
R6556 VDD.n3233 VDD.n3232 10.6151
R6557 VDD.n3232 VDD.n3230 10.6151
R6558 VDD.n3230 VDD.n3229 10.6151
R6559 VDD.n3229 VDD.n3227 10.6151
R6560 VDD.n3227 VDD.n3226 10.6151
R6561 VDD.n3226 VDD.n3224 10.6151
R6562 VDD.n3224 VDD.n3223 10.6151
R6563 VDD.n3223 VDD.n3221 10.6151
R6564 VDD.n3221 VDD.n3220 10.6151
R6565 VDD.n3220 VDD.n3218 10.6151
R6566 VDD.n3218 VDD.n3217 10.6151
R6567 VDD.n3217 VDD.n3215 10.6151
R6568 VDD.n3215 VDD.n3214 10.6151
R6569 VDD.n3214 VDD.n3212 10.6151
R6570 VDD.n3212 VDD.n3211 10.6151
R6571 VDD.n3211 VDD.n3209 10.6151
R6572 VDD.n3209 VDD.n3208 10.6151
R6573 VDD.n3208 VDD.n3206 10.6151
R6574 VDD.n3206 VDD.n3205 10.6151
R6575 VDD.n3205 VDD.n3203 10.6151
R6576 VDD.n3203 VDD.n3202 10.6151
R6577 VDD.n3202 VDD.n3200 10.6151
R6578 VDD.n3200 VDD.n3199 10.6151
R6579 VDD.n3199 VDD.n3197 10.6151
R6580 VDD.n3197 VDD.n3196 10.6151
R6581 VDD.n3196 VDD.n3194 10.6151
R6582 VDD.n3194 VDD.n3193 10.6151
R6583 VDD.n3193 VDD.n3191 10.6151
R6584 VDD.n3191 VDD.n3190 10.6151
R6585 VDD.n3190 VDD.n3188 10.6151
R6586 VDD.n3188 VDD.n3187 10.6151
R6587 VDD.n3187 VDD.n3185 10.6151
R6588 VDD.n3185 VDD.n3184 10.6151
R6589 VDD.n3184 VDD.n3182 10.6151
R6590 VDD.n3182 VDD.n3181 10.6151
R6591 VDD.n3181 VDD.n3179 10.6151
R6592 VDD.n3179 VDD.n3178 10.6151
R6593 VDD.n3178 VDD.n3176 10.6151
R6594 VDD.n3176 VDD.n3175 10.6151
R6595 VDD.n3175 VDD.n3173 10.6151
R6596 VDD.n3173 VDD.n3172 10.6151
R6597 VDD.n3172 VDD.n3170 10.6151
R6598 VDD.n3170 VDD.n3169 10.6151
R6599 VDD.n3169 VDD.n3167 10.6151
R6600 VDD.n3167 VDD.n3166 10.6151
R6601 VDD.n3166 VDD.n3164 10.6151
R6602 VDD.n3164 VDD.n3163 10.6151
R6603 VDD.n3163 VDD.n3161 10.6151
R6604 VDD.n3161 VDD.n3160 10.6151
R6605 VDD.n3160 VDD.n3158 10.6151
R6606 VDD.n3158 VDD.n3157 10.6151
R6607 VDD.n3157 VDD.n3155 10.6151
R6608 VDD.n3155 VDD.n3154 10.6151
R6609 VDD.n3154 VDD.n3152 10.6151
R6610 VDD.n3152 VDD.n3151 10.6151
R6611 VDD.n3151 VDD.n3149 10.6151
R6612 VDD.n3149 VDD.n3148 10.6151
R6613 VDD.n3148 VDD.n3146 10.6151
R6614 VDD.n3146 VDD.n3145 10.6151
R6615 VDD.n3145 VDD.n3143 10.6151
R6616 VDD.n3143 VDD.n3142 10.6151
R6617 VDD.n3142 VDD.n3140 10.6151
R6618 VDD.n3140 VDD.n3139 10.6151
R6619 VDD.n3139 VDD.n3137 10.6151
R6620 VDD.n3137 VDD.n3136 10.6151
R6621 VDD.n3136 VDD.n3134 10.6151
R6622 VDD.n3134 VDD.n3133 10.6151
R6623 VDD.n3133 VDD.n3131 10.6151
R6624 VDD.n3131 VDD.n3130 10.6151
R6625 VDD.n3130 VDD.n3128 10.6151
R6626 VDD.n3128 VDD.n3127 10.6151
R6627 VDD.n3127 VDD.n3125 10.6151
R6628 VDD.n3125 VDD.n3124 10.6151
R6629 VDD.n3124 VDD.n235 10.6151
R6630 VDD.n3332 VDD.n3331 10.6151
R6631 VDD.n3331 VDD.n3114 10.6151
R6632 VDD.n3325 VDD.n3114 10.6151
R6633 VDD.n3325 VDD.n3324 10.6151
R6634 VDD.n3324 VDD.n3323 10.6151
R6635 VDD.n3323 VDD.n3116 10.6151
R6636 VDD.n3317 VDD.n3116 10.6151
R6637 VDD.n3317 VDD.n3316 10.6151
R6638 VDD.n3316 VDD.n3315 10.6151
R6639 VDD.n3315 VDD.n3118 10.6151
R6640 VDD.n3309 VDD.n3118 10.6151
R6641 VDD.n3309 VDD.n3308 10.6151
R6642 VDD.n3308 VDD.n3307 10.6151
R6643 VDD.n3307 VDD.n3122 10.6151
R6644 VDD.n3301 VDD.n3122 10.6151
R6645 VDD.n3301 VDD.n3300 10.6151
R6646 VDD.n3300 VDD.n3299 10.6151
R6647 VDD.n3333 VDD.n594 10.6151
R6648 VDD.n3343 VDD.n594 10.6151
R6649 VDD.n3344 VDD.n3343 10.6151
R6650 VDD.n3345 VDD.n3344 10.6151
R6651 VDD.n3345 VDD.n582 10.6151
R6652 VDD.n3355 VDD.n582 10.6151
R6653 VDD.n3356 VDD.n3355 10.6151
R6654 VDD.n3357 VDD.n3356 10.6151
R6655 VDD.n3357 VDD.n570 10.6151
R6656 VDD.n3367 VDD.n570 10.6151
R6657 VDD.n3368 VDD.n3367 10.6151
R6658 VDD.n3369 VDD.n3368 10.6151
R6659 VDD.n3369 VDD.n558 10.6151
R6660 VDD.n3379 VDD.n558 10.6151
R6661 VDD.n3380 VDD.n3379 10.6151
R6662 VDD.n3381 VDD.n3380 10.6151
R6663 VDD.n3381 VDD.n546 10.6151
R6664 VDD.n3391 VDD.n546 10.6151
R6665 VDD.n3392 VDD.n3391 10.6151
R6666 VDD.n3393 VDD.n3392 10.6151
R6667 VDD.n3393 VDD.n534 10.6151
R6668 VDD.n3403 VDD.n534 10.6151
R6669 VDD.n3404 VDD.n3403 10.6151
R6670 VDD.n3405 VDD.n3404 10.6151
R6671 VDD.n3405 VDD.n522 10.6151
R6672 VDD.n3415 VDD.n522 10.6151
R6673 VDD.n3416 VDD.n3415 10.6151
R6674 VDD.n3417 VDD.n3416 10.6151
R6675 VDD.n3417 VDD.n509 10.6151
R6676 VDD.n3427 VDD.n509 10.6151
R6677 VDD.n3428 VDD.n3427 10.6151
R6678 VDD.n3429 VDD.n3428 10.6151
R6679 VDD.n3429 VDD.n498 10.6151
R6680 VDD.n3439 VDD.n498 10.6151
R6681 VDD.n3440 VDD.n3439 10.6151
R6682 VDD.n3441 VDD.n3440 10.6151
R6683 VDD.n3441 VDD.n486 10.6151
R6684 VDD.n3451 VDD.n486 10.6151
R6685 VDD.n3452 VDD.n3451 10.6151
R6686 VDD.n3453 VDD.n3452 10.6151
R6687 VDD.n3453 VDD.n474 10.6151
R6688 VDD.n3463 VDD.n474 10.6151
R6689 VDD.n3464 VDD.n3463 10.6151
R6690 VDD.n3465 VDD.n3464 10.6151
R6691 VDD.n3465 VDD.n462 10.6151
R6692 VDD.n3475 VDD.n462 10.6151
R6693 VDD.n3476 VDD.n3475 10.6151
R6694 VDD.n3477 VDD.n3476 10.6151
R6695 VDD.n3477 VDD.n450 10.6151
R6696 VDD.n3487 VDD.n450 10.6151
R6697 VDD.n3488 VDD.n3487 10.6151
R6698 VDD.n3489 VDD.n3488 10.6151
R6699 VDD.n3489 VDD.n438 10.6151
R6700 VDD.n3499 VDD.n438 10.6151
R6701 VDD.n3500 VDD.n3499 10.6151
R6702 VDD.n3501 VDD.n3500 10.6151
R6703 VDD.n3501 VDD.n426 10.6151
R6704 VDD.n3511 VDD.n426 10.6151
R6705 VDD.n3512 VDD.n3511 10.6151
R6706 VDD.n3513 VDD.n3512 10.6151
R6707 VDD.n3513 VDD.n413 10.6151
R6708 VDD.n3523 VDD.n413 10.6151
R6709 VDD.n3524 VDD.n3523 10.6151
R6710 VDD.n3525 VDD.n3524 10.6151
R6711 VDD.n3525 VDD.n402 10.6151
R6712 VDD.n3535 VDD.n402 10.6151
R6713 VDD.n3536 VDD.n3535 10.6151
R6714 VDD.n3537 VDD.n3536 10.6151
R6715 VDD.n3537 VDD.n390 10.6151
R6716 VDD.n3547 VDD.n390 10.6151
R6717 VDD.n3548 VDD.n3547 10.6151
R6718 VDD.n3549 VDD.n3548 10.6151
R6719 VDD.n3549 VDD.n378 10.6151
R6720 VDD.n3559 VDD.n378 10.6151
R6721 VDD.n3560 VDD.n3559 10.6151
R6722 VDD.n3561 VDD.n3560 10.6151
R6723 VDD.n3561 VDD.n366 10.6151
R6724 VDD.n3571 VDD.n366 10.6151
R6725 VDD.n3572 VDD.n3571 10.6151
R6726 VDD.n3573 VDD.n3572 10.6151
R6727 VDD.n3573 VDD.n354 10.6151
R6728 VDD.n3583 VDD.n354 10.6151
R6729 VDD.n3584 VDD.n3583 10.6151
R6730 VDD.n3585 VDD.n3584 10.6151
R6731 VDD.n3585 VDD.n342 10.6151
R6732 VDD.n3595 VDD.n342 10.6151
R6733 VDD.n3596 VDD.n3595 10.6151
R6734 VDD.n3597 VDD.n3596 10.6151
R6735 VDD.n3597 VDD.n330 10.6151
R6736 VDD.n3607 VDD.n330 10.6151
R6737 VDD.n3608 VDD.n3607 10.6151
R6738 VDD.n3609 VDD.n3608 10.6151
R6739 VDD.n3609 VDD.n318 10.6151
R6740 VDD.n3619 VDD.n318 10.6151
R6741 VDD.n3620 VDD.n3619 10.6151
R6742 VDD.n3621 VDD.n3620 10.6151
R6743 VDD.n3621 VDD.n306 10.6151
R6744 VDD.n3631 VDD.n306 10.6151
R6745 VDD.n3632 VDD.n3631 10.6151
R6746 VDD.n3633 VDD.n3632 10.6151
R6747 VDD.n3633 VDD.n294 10.6151
R6748 VDD.n3643 VDD.n294 10.6151
R6749 VDD.n3644 VDD.n3643 10.6151
R6750 VDD.n3645 VDD.n3644 10.6151
R6751 VDD.n3645 VDD.n282 10.6151
R6752 VDD.n3655 VDD.n282 10.6151
R6753 VDD.n3656 VDD.n3655 10.6151
R6754 VDD.n3657 VDD.n3656 10.6151
R6755 VDD.n3657 VDD.n270 10.6151
R6756 VDD.n3667 VDD.n270 10.6151
R6757 VDD.n3668 VDD.n3667 10.6151
R6758 VDD.n3695 VDD.n3668 10.6151
R6759 VDD.n3695 VDD.n3694 10.6151
R6760 VDD.n3694 VDD.n3693 10.6151
R6761 VDD.n3693 VDD.n3692 10.6151
R6762 VDD.n3692 VDD.n3690 10.6151
R6763 VDD.n2472 VDD.n972 10.6151
R6764 VDD.n2473 VDD.n2472 10.6151
R6765 VDD.n2474 VDD.n2473 10.6151
R6766 VDD.n2474 VDD.n960 10.6151
R6767 VDD.n2484 VDD.n960 10.6151
R6768 VDD.n2485 VDD.n2484 10.6151
R6769 VDD.n2486 VDD.n2485 10.6151
R6770 VDD.n2486 VDD.n948 10.6151
R6771 VDD.n2496 VDD.n948 10.6151
R6772 VDD.n2497 VDD.n2496 10.6151
R6773 VDD.n2498 VDD.n2497 10.6151
R6774 VDD.n2498 VDD.n937 10.6151
R6775 VDD.n2508 VDD.n937 10.6151
R6776 VDD.n2509 VDD.n2508 10.6151
R6777 VDD.n2510 VDD.n2509 10.6151
R6778 VDD.n2510 VDD.n925 10.6151
R6779 VDD.n2520 VDD.n925 10.6151
R6780 VDD.n2521 VDD.n2520 10.6151
R6781 VDD.n2522 VDD.n2521 10.6151
R6782 VDD.n2522 VDD.n913 10.6151
R6783 VDD.n2532 VDD.n913 10.6151
R6784 VDD.n2533 VDD.n2532 10.6151
R6785 VDD.n2534 VDD.n2533 10.6151
R6786 VDD.n2534 VDD.n900 10.6151
R6787 VDD.n2544 VDD.n900 10.6151
R6788 VDD.n2545 VDD.n2544 10.6151
R6789 VDD.n2546 VDD.n2545 10.6151
R6790 VDD.n2546 VDD.n889 10.6151
R6791 VDD.n2556 VDD.n889 10.6151
R6792 VDD.n2557 VDD.n2556 10.6151
R6793 VDD.n2558 VDD.n2557 10.6151
R6794 VDD.n2558 VDD.n877 10.6151
R6795 VDD.n2568 VDD.n877 10.6151
R6796 VDD.n2569 VDD.n2568 10.6151
R6797 VDD.n2570 VDD.n2569 10.6151
R6798 VDD.n2570 VDD.n865 10.6151
R6799 VDD.n2580 VDD.n865 10.6151
R6800 VDD.n2581 VDD.n2580 10.6151
R6801 VDD.n2582 VDD.n2581 10.6151
R6802 VDD.n2582 VDD.n853 10.6151
R6803 VDD.n2592 VDD.n853 10.6151
R6804 VDD.n2593 VDD.n2592 10.6151
R6805 VDD.n2594 VDD.n2593 10.6151
R6806 VDD.n2594 VDD.n841 10.6151
R6807 VDD.n2604 VDD.n841 10.6151
R6808 VDD.n2605 VDD.n2604 10.6151
R6809 VDD.n2606 VDD.n2605 10.6151
R6810 VDD.n2606 VDD.n829 10.6151
R6811 VDD.n2616 VDD.n829 10.6151
R6812 VDD.n2617 VDD.n2616 10.6151
R6813 VDD.n2618 VDD.n2617 10.6151
R6814 VDD.n2618 VDD.n817 10.6151
R6815 VDD.n2628 VDD.n817 10.6151
R6816 VDD.n2629 VDD.n2628 10.6151
R6817 VDD.n2630 VDD.n2629 10.6151
R6818 VDD.n2630 VDD.n805 10.6151
R6819 VDD.n2640 VDD.n805 10.6151
R6820 VDD.n2641 VDD.n2640 10.6151
R6821 VDD.n2642 VDD.n2641 10.6151
R6822 VDD.n2642 VDD.n793 10.6151
R6823 VDD.n2652 VDD.n793 10.6151
R6824 VDD.n2653 VDD.n2652 10.6151
R6825 VDD.n2654 VDD.n2653 10.6151
R6826 VDD.n2654 VDD.n780 10.6151
R6827 VDD.n2664 VDD.n780 10.6151
R6828 VDD.n2665 VDD.n2664 10.6151
R6829 VDD.n2666 VDD.n2665 10.6151
R6830 VDD.n2666 VDD.n768 10.6151
R6831 VDD.n2676 VDD.n768 10.6151
R6832 VDD.n2677 VDD.n2676 10.6151
R6833 VDD.n2678 VDD.n2677 10.6151
R6834 VDD.n2678 VDD.n757 10.6151
R6835 VDD.n2688 VDD.n757 10.6151
R6836 VDD.n2689 VDD.n2688 10.6151
R6837 VDD.n2690 VDD.n2689 10.6151
R6838 VDD.n2690 VDD.n745 10.6151
R6839 VDD.n2700 VDD.n745 10.6151
R6840 VDD.n2701 VDD.n2700 10.6151
R6841 VDD.n2702 VDD.n2701 10.6151
R6842 VDD.n2702 VDD.n733 10.6151
R6843 VDD.n2712 VDD.n733 10.6151
R6844 VDD.n2713 VDD.n2712 10.6151
R6845 VDD.n2714 VDD.n2713 10.6151
R6846 VDD.n2714 VDD.n721 10.6151
R6847 VDD.n2724 VDD.n721 10.6151
R6848 VDD.n2725 VDD.n2724 10.6151
R6849 VDD.n2726 VDD.n2725 10.6151
R6850 VDD.n2726 VDD.n709 10.6151
R6851 VDD.n2736 VDD.n709 10.6151
R6852 VDD.n2737 VDD.n2736 10.6151
R6853 VDD.n2738 VDD.n2737 10.6151
R6854 VDD.n2738 VDD.n697 10.6151
R6855 VDD.n2748 VDD.n697 10.6151
R6856 VDD.n2749 VDD.n2748 10.6151
R6857 VDD.n2750 VDD.n2749 10.6151
R6858 VDD.n2750 VDD.n685 10.6151
R6859 VDD.n2760 VDD.n685 10.6151
R6860 VDD.n2761 VDD.n2760 10.6151
R6861 VDD.n2762 VDD.n2761 10.6151
R6862 VDD.n2762 VDD.n673 10.6151
R6863 VDD.n2772 VDD.n673 10.6151
R6864 VDD.n2773 VDD.n2772 10.6151
R6865 VDD.n2774 VDD.n2773 10.6151
R6866 VDD.n2774 VDD.n661 10.6151
R6867 VDD.n2784 VDD.n661 10.6151
R6868 VDD.n2785 VDD.n2784 10.6151
R6869 VDD.n2786 VDD.n2785 10.6151
R6870 VDD.n2786 VDD.n649 10.6151
R6871 VDD.n2796 VDD.n649 10.6151
R6872 VDD.n2797 VDD.n2796 10.6151
R6873 VDD.n2803 VDD.n2797 10.6151
R6874 VDD.n2803 VDD.n2802 10.6151
R6875 VDD.n2802 VDD.n2801 10.6151
R6876 VDD.n2801 VDD.n2800 10.6151
R6877 VDD.n2800 VDD.n2798 10.6151
R6878 VDD.n2798 VDD.n623 10.6151
R6879 VDD.n2893 VDD.n2892 10.6151
R6880 VDD.n2892 VDD.n2891 10.6151
R6881 VDD.n2891 VDD.n2888 10.6151
R6882 VDD.n2888 VDD.n2887 10.6151
R6883 VDD.n2887 VDD.n2884 10.6151
R6884 VDD.n2884 VDD.n2883 10.6151
R6885 VDD.n2883 VDD.n2880 10.6151
R6886 VDD.n2880 VDD.n2879 10.6151
R6887 VDD.n2879 VDD.n2876 10.6151
R6888 VDD.n2876 VDD.n2875 10.6151
R6889 VDD.n2875 VDD.n2872 10.6151
R6890 VDD.n2872 VDD.n2871 10.6151
R6891 VDD.n2871 VDD.n2868 10.6151
R6892 VDD.n2868 VDD.n2867 10.6151
R6893 VDD.n2867 VDD.n2864 10.6151
R6894 VDD.n2864 VDD.n2863 10.6151
R6895 VDD.n2863 VDD.n2861 10.6151
R6896 VDD.n2245 VDD.n2244 10.6151
R6897 VDD.n2247 VDD.n2245 10.6151
R6898 VDD.n2248 VDD.n2247 10.6151
R6899 VDD.n2250 VDD.n2248 10.6151
R6900 VDD.n2251 VDD.n2250 10.6151
R6901 VDD.n2253 VDD.n2251 10.6151
R6902 VDD.n2254 VDD.n2253 10.6151
R6903 VDD.n2256 VDD.n2254 10.6151
R6904 VDD.n2257 VDD.n2256 10.6151
R6905 VDD.n2413 VDD.n2257 10.6151
R6906 VDD.n2413 VDD.n2412 10.6151
R6907 VDD.n2412 VDD.n2411 10.6151
R6908 VDD.n2411 VDD.n2409 10.6151
R6909 VDD.n2409 VDD.n2408 10.6151
R6910 VDD.n2408 VDD.n2406 10.6151
R6911 VDD.n2406 VDD.n2405 10.6151
R6912 VDD.n2405 VDD.n2403 10.6151
R6913 VDD.n2403 VDD.n2402 10.6151
R6914 VDD.n2402 VDD.n2400 10.6151
R6915 VDD.n2400 VDD.n2399 10.6151
R6916 VDD.n2399 VDD.n2397 10.6151
R6917 VDD.n2397 VDD.n2396 10.6151
R6918 VDD.n2396 VDD.n2394 10.6151
R6919 VDD.n2394 VDD.n2393 10.6151
R6920 VDD.n2393 VDD.n2391 10.6151
R6921 VDD.n2391 VDD.n2390 10.6151
R6922 VDD.n2390 VDD.n2388 10.6151
R6923 VDD.n2388 VDD.n2387 10.6151
R6924 VDD.n2387 VDD.n2385 10.6151
R6925 VDD.n2385 VDD.n2384 10.6151
R6926 VDD.n2384 VDD.n2382 10.6151
R6927 VDD.n2382 VDD.n2381 10.6151
R6928 VDD.n2381 VDD.n2379 10.6151
R6929 VDD.n2379 VDD.n2378 10.6151
R6930 VDD.n2378 VDD.n2376 10.6151
R6931 VDD.n2376 VDD.n2375 10.6151
R6932 VDD.n2375 VDD.n2373 10.6151
R6933 VDD.n2373 VDD.n2372 10.6151
R6934 VDD.n2372 VDD.n2370 10.6151
R6935 VDD.n2370 VDD.n2369 10.6151
R6936 VDD.n2369 VDD.n2367 10.6151
R6937 VDD.n2367 VDD.n2366 10.6151
R6938 VDD.n2366 VDD.n2364 10.6151
R6939 VDD.n2364 VDD.n2363 10.6151
R6940 VDD.n2363 VDD.n2361 10.6151
R6941 VDD.n2361 VDD.n2360 10.6151
R6942 VDD.n2360 VDD.n2358 10.6151
R6943 VDD.n2358 VDD.n2357 10.6151
R6944 VDD.n2357 VDD.n2355 10.6151
R6945 VDD.n2355 VDD.n2354 10.6151
R6946 VDD.n2354 VDD.n2352 10.6151
R6947 VDD.n2352 VDD.n2351 10.6151
R6948 VDD.n2351 VDD.n2349 10.6151
R6949 VDD.n2349 VDD.n2348 10.6151
R6950 VDD.n2348 VDD.n2346 10.6151
R6951 VDD.n2346 VDD.n2345 10.6151
R6952 VDD.n2345 VDD.n2343 10.6151
R6953 VDD.n2343 VDD.n2342 10.6151
R6954 VDD.n2342 VDD.n2340 10.6151
R6955 VDD.n2340 VDD.n2339 10.6151
R6956 VDD.n2339 VDD.n2337 10.6151
R6957 VDD.n2337 VDD.n2336 10.6151
R6958 VDD.n2336 VDD.n2334 10.6151
R6959 VDD.n2334 VDD.n2333 10.6151
R6960 VDD.n2333 VDD.n2331 10.6151
R6961 VDD.n2331 VDD.n2330 10.6151
R6962 VDD.n2330 VDD.n2328 10.6151
R6963 VDD.n2328 VDD.n2327 10.6151
R6964 VDD.n2327 VDD.n2325 10.6151
R6965 VDD.n2325 VDD.n2324 10.6151
R6966 VDD.n2324 VDD.n2322 10.6151
R6967 VDD.n2322 VDD.n2321 10.6151
R6968 VDD.n2321 VDD.n2319 10.6151
R6969 VDD.n2319 VDD.n2318 10.6151
R6970 VDD.n2318 VDD.n2316 10.6151
R6971 VDD.n2316 VDD.n2315 10.6151
R6972 VDD.n2315 VDD.n2313 10.6151
R6973 VDD.n2313 VDD.n2312 10.6151
R6974 VDD.n2312 VDD.n2310 10.6151
R6975 VDD.n2310 VDD.n2309 10.6151
R6976 VDD.n2309 VDD.n2307 10.6151
R6977 VDD.n2307 VDD.n2306 10.6151
R6978 VDD.n2306 VDD.n2304 10.6151
R6979 VDD.n2304 VDD.n2303 10.6151
R6980 VDD.n2303 VDD.n2301 10.6151
R6981 VDD.n2301 VDD.n2300 10.6151
R6982 VDD.n2300 VDD.n2298 10.6151
R6983 VDD.n2298 VDD.n2297 10.6151
R6984 VDD.n2297 VDD.n2295 10.6151
R6985 VDD.n2295 VDD.n2294 10.6151
R6986 VDD.n2294 VDD.n2292 10.6151
R6987 VDD.n2292 VDD.n2291 10.6151
R6988 VDD.n2291 VDD.n2289 10.6151
R6989 VDD.n2289 VDD.n2288 10.6151
R6990 VDD.n2288 VDD.n2286 10.6151
R6991 VDD.n2286 VDD.n2285 10.6151
R6992 VDD.n2285 VDD.n2283 10.6151
R6993 VDD.n2283 VDD.n2282 10.6151
R6994 VDD.n2282 VDD.n2280 10.6151
R6995 VDD.n2280 VDD.n2279 10.6151
R6996 VDD.n2279 VDD.n2277 10.6151
R6997 VDD.n2277 VDD.n2276 10.6151
R6998 VDD.n2276 VDD.n2274 10.6151
R6999 VDD.n2274 VDD.n2273 10.6151
R7000 VDD.n2273 VDD.n2271 10.6151
R7001 VDD.n2271 VDD.n2270 10.6151
R7002 VDD.n2270 VDD.n2268 10.6151
R7003 VDD.n2268 VDD.n2267 10.6151
R7004 VDD.n2267 VDD.n2265 10.6151
R7005 VDD.n2265 VDD.n2264 10.6151
R7006 VDD.n2264 VDD.n2262 10.6151
R7007 VDD.n2262 VDD.n2261 10.6151
R7008 VDD.n2261 VDD.n2259 10.6151
R7009 VDD.n2259 VDD.n2258 10.6151
R7010 VDD.n2258 VDD.n626 10.6151
R7011 VDD.n2860 VDD.n626 10.6151
R7012 VDD.n2211 VDD.n2209 10.6151
R7013 VDD.n2212 VDD.n2211 10.6151
R7014 VDD.n2215 VDD.n2212 10.6151
R7015 VDD.n2216 VDD.n2215 10.6151
R7016 VDD.n2219 VDD.n2216 10.6151
R7017 VDD.n2220 VDD.n2219 10.6151
R7018 VDD.n2223 VDD.n2220 10.6151
R7019 VDD.n2224 VDD.n2223 10.6151
R7020 VDD.n2228 VDD.n2227 10.6151
R7021 VDD.n2231 VDD.n2228 10.6151
R7022 VDD.n2232 VDD.n2231 10.6151
R7023 VDD.n2235 VDD.n2232 10.6151
R7024 VDD.n2236 VDD.n2235 10.6151
R7025 VDD.n2239 VDD.n2236 10.6151
R7026 VDD.n2241 VDD.n2239 10.6151
R7027 VDD.n2242 VDD.n2241 10.6151
R7028 VDD.n1835 VDD.n1297 9.3005
R7029 VDD.n1837 VDD.n1836 9.3005
R7030 VDD.n1287 VDD.n1286 9.3005
R7031 VDD.n1850 VDD.n1849 9.3005
R7032 VDD.n1851 VDD.n1285 9.3005
R7033 VDD.n1853 VDD.n1852 9.3005
R7034 VDD.n1275 VDD.n1274 9.3005
R7035 VDD.n1866 VDD.n1865 9.3005
R7036 VDD.n1867 VDD.n1273 9.3005
R7037 VDD.n1869 VDD.n1868 9.3005
R7038 VDD.n1263 VDD.n1262 9.3005
R7039 VDD.n1882 VDD.n1881 9.3005
R7040 VDD.n1883 VDD.n1261 9.3005
R7041 VDD.n1885 VDD.n1884 9.3005
R7042 VDD.n1251 VDD.n1250 9.3005
R7043 VDD.n1898 VDD.n1897 9.3005
R7044 VDD.n1899 VDD.n1249 9.3005
R7045 VDD.n1901 VDD.n1900 9.3005
R7046 VDD.n1239 VDD.n1238 9.3005
R7047 VDD.n1914 VDD.n1913 9.3005
R7048 VDD.n1915 VDD.n1237 9.3005
R7049 VDD.n1917 VDD.n1916 9.3005
R7050 VDD.n1227 VDD.n1226 9.3005
R7051 VDD.n1930 VDD.n1929 9.3005
R7052 VDD.n1931 VDD.n1225 9.3005
R7053 VDD.n1933 VDD.n1932 9.3005
R7054 VDD.n1214 VDD.n1213 9.3005
R7055 VDD.n1948 VDD.n1947 9.3005
R7056 VDD.n1949 VDD.n1212 9.3005
R7057 VDD.n2168 VDD.n2167 9.3005
R7058 VDD.n2164 VDD.n1950 9.3005
R7059 VDD.n1954 VDD.n1951 9.3005
R7060 VDD.n2159 VDD.n1955 9.3005
R7061 VDD.n2158 VDD.n1956 9.3005
R7062 VDD.n2157 VDD.n1957 9.3005
R7063 VDD.n1961 VDD.n1958 9.3005
R7064 VDD.n2152 VDD.n1962 9.3005
R7065 VDD.n2151 VDD.n1963 9.3005
R7066 VDD.n2150 VDD.n1964 9.3005
R7067 VDD.n1968 VDD.n1965 9.3005
R7068 VDD.n2145 VDD.n1969 9.3005
R7069 VDD.n2144 VDD.n1970 9.3005
R7070 VDD.n2143 VDD.n1971 9.3005
R7071 VDD.n1978 VDD.n1972 9.3005
R7072 VDD.n2166 VDD.n2165 9.3005
R7073 VDD.n2077 VDD.n2076 9.3005
R7074 VDD.n2075 VDD.n2040 9.3005
R7075 VDD.n2074 VDD.n2073 9.3005
R7076 VDD.n2043 VDD.n2042 9.3005
R7077 VDD.n2068 VDD.n2046 9.3005
R7078 VDD.n2067 VDD.n2047 9.3005
R7079 VDD.n2066 VDD.n2048 9.3005
R7080 VDD.n2050 VDD.n2049 9.3005
R7081 VDD.n2061 VDD.n1156 9.3005
R7082 VDD.n2010 VDD.n2008 9.3005
R7083 VDD.n2105 VDD.n2011 9.3005
R7084 VDD.n2104 VDD.n2012 9.3005
R7085 VDD.n2103 VDD.n2013 9.3005
R7086 VDD.n2017 VDD.n2014 9.3005
R7087 VDD.n2098 VDD.n2018 9.3005
R7088 VDD.n2097 VDD.n2019 9.3005
R7089 VDD.n2096 VDD.n2020 9.3005
R7090 VDD.n2024 VDD.n2021 9.3005
R7091 VDD.n2091 VDD.n2025 9.3005
R7092 VDD.n2090 VDD.n2026 9.3005
R7093 VDD.n2089 VDD.n2027 9.3005
R7094 VDD.n2031 VDD.n2028 9.3005
R7095 VDD.n2084 VDD.n2032 9.3005
R7096 VDD.n2083 VDD.n2033 9.3005
R7097 VDD.n2082 VDD.n2034 9.3005
R7098 VDD.n2041 VDD.n2037 9.3005
R7099 VDD.n2138 VDD.n1979 9.3005
R7100 VDD.n2137 VDD.n1980 9.3005
R7101 VDD.n2136 VDD.n1981 9.3005
R7102 VDD.n1985 VDD.n1982 9.3005
R7103 VDD.n2131 VDD.n1986 9.3005
R7104 VDD.n2130 VDD.n1987 9.3005
R7105 VDD.n2129 VDD.n1988 9.3005
R7106 VDD.n2120 VDD.n2119 9.3005
R7107 VDD.n1995 VDD.n1994 9.3005
R7108 VDD.n2000 VDD.n1998 9.3005
R7109 VDD.n2112 VDD.n2001 9.3005
R7110 VDD.n2111 VDD.n2002 9.3005
R7111 VDD.n2110 VDD.n2003 9.3005
R7112 VDD.n204 VDD.n202 9.3005
R7113 VDD.n3873 VDD.n201 9.3005
R7114 VDD.n3874 VDD.n200 9.3005
R7115 VDD.n3875 VDD.n199 9.3005
R7116 VDD.n198 VDD.n196 9.3005
R7117 VDD.n3881 VDD.n195 9.3005
R7118 VDD.n3882 VDD.n194 9.3005
R7119 VDD.n3883 VDD.n193 9.3005
R7120 VDD.n192 VDD.n190 9.3005
R7121 VDD.n3889 VDD.n189 9.3005
R7122 VDD.n3890 VDD.n188 9.3005
R7123 VDD.n3891 VDD.n187 9.3005
R7124 VDD.n186 VDD.n184 9.3005
R7125 VDD.n3897 VDD.n183 9.3005
R7126 VDD.n3898 VDD.n182 9.3005
R7127 VDD.n3899 VDD.n181 9.3005
R7128 VDD.n3867 VDD.n205 9.3005
R7129 VDD.n180 VDD.n175 9.3005
R7130 VDD.n3905 VDD.n174 9.3005
R7131 VDD.n3906 VDD.n173 9.3005
R7132 VDD.n3907 VDD.n172 9.3005
R7133 VDD.n171 VDD.n169 9.3005
R7134 VDD.n3913 VDD.n163 9.3005
R7135 VDD.n3916 VDD.n160 9.3005
R7136 VDD.n3925 VDD.n159 9.3005
R7137 VDD.n3926 VDD.n158 9.3005
R7138 VDD.n3927 VDD.n157 9.3005
R7139 VDD.n156 VDD.n154 9.3005
R7140 VDD.n3933 VDD.n153 9.3005
R7141 VDD.n3934 VDD.n152 9.3005
R7142 VDD.n3936 VDD.n149 9.3005
R7143 VDD.n148 VDD.n146 9.3005
R7144 VDD.n3942 VDD.n145 9.3005
R7145 VDD.n3943 VDD.n144 9.3005
R7146 VDD.n3944 VDD.n143 9.3005
R7147 VDD.n142 VDD.n140 9.3005
R7148 VDD.n3950 VDD.n139 9.3005
R7149 VDD.n3951 VDD.n138 9.3005
R7150 VDD.n3952 VDD.n137 9.3005
R7151 VDD.n136 VDD.n134 9.3005
R7152 VDD.n3957 VDD.n133 9.3005
R7153 VDD.n3958 VDD.n132 9.3005
R7154 VDD.n131 VDD.n129 9.3005
R7155 VDD.n3963 VDD.n128 9.3005
R7156 VDD.n3965 VDD.n3964 9.3005
R7157 VDD.n3967 VDD.n3966 9.3005
R7158 VDD.n119 VDD.n118 9.3005
R7159 VDD.n3980 VDD.n3979 9.3005
R7160 VDD.n3981 VDD.n117 9.3005
R7161 VDD.n3983 VDD.n3982 9.3005
R7162 VDD.n107 VDD.n106 9.3005
R7163 VDD.n3996 VDD.n3995 9.3005
R7164 VDD.n3997 VDD.n105 9.3005
R7165 VDD.n3999 VDD.n3998 9.3005
R7166 VDD.n95 VDD.n94 9.3005
R7167 VDD.n4012 VDD.n4011 9.3005
R7168 VDD.n4013 VDD.n93 9.3005
R7169 VDD.n4015 VDD.n4014 9.3005
R7170 VDD.n83 VDD.n82 9.3005
R7171 VDD.n4028 VDD.n4027 9.3005
R7172 VDD.n4029 VDD.n81 9.3005
R7173 VDD.n4031 VDD.n4030 9.3005
R7174 VDD.n71 VDD.n70 9.3005
R7175 VDD.n4045 VDD.n4044 9.3005
R7176 VDD.n4046 VDD.n69 9.3005
R7177 VDD.n4048 VDD.n4047 9.3005
R7178 VDD.n60 VDD.n59 9.3005
R7179 VDD.n4061 VDD.n4060 9.3005
R7180 VDD.n4062 VDD.n58 9.3005
R7181 VDD.n4064 VDD.n4063 9.3005
R7182 VDD.n48 VDD.n47 9.3005
R7183 VDD.n4077 VDD.n4076 9.3005
R7184 VDD.n4078 VDD.n46 9.3005
R7185 VDD.n4080 VDD.n4079 9.3005
R7186 VDD.n32 VDD.n30 9.3005
R7187 VDD.n4604 VDD.n4603 9.3005
R7188 VDD.n33 VDD.n31 9.3005
R7189 VDD.n4594 VDD.n4094 9.3005
R7190 VDD.n4593 VDD.n4095 9.3005
R7191 VDD.n4592 VDD.n4096 9.3005
R7192 VDD.n4104 VDD.n4097 9.3005
R7193 VDD.n4586 VDD.n4105 9.3005
R7194 VDD.n4585 VDD.n4106 9.3005
R7195 VDD.n4584 VDD.n4107 9.3005
R7196 VDD.n4114 VDD.n4108 9.3005
R7197 VDD.n4578 VDD.n4115 9.3005
R7198 VDD.n4577 VDD.n4116 9.3005
R7199 VDD.n4576 VDD.n4117 9.3005
R7200 VDD.n4126 VDD.n4118 9.3005
R7201 VDD.n4570 VDD.n4127 9.3005
R7202 VDD.n4569 VDD.n4128 9.3005
R7203 VDD.n4568 VDD.n4129 9.3005
R7204 VDD.n4137 VDD.n4130 9.3005
R7205 VDD.n4562 VDD.n4138 9.3005
R7206 VDD.n4561 VDD.n4139 9.3005
R7207 VDD.n4560 VDD.n4140 9.3005
R7208 VDD.n4148 VDD.n4141 9.3005
R7209 VDD.n4554 VDD.n4149 9.3005
R7210 VDD.n4553 VDD.n4150 9.3005
R7211 VDD.n4552 VDD.n4151 9.3005
R7212 VDD.n4159 VDD.n4152 9.3005
R7213 VDD.n4546 VDD.n4160 9.3005
R7214 VDD.n4545 VDD.n4161 9.3005
R7215 VDD.n4544 VDD.n4162 9.3005
R7216 VDD.n4170 VDD.n4163 9.3005
R7217 VDD.n4538 VDD.n4537 9.3005
R7218 VDD.n4534 VDD.n4171 9.3005
R7219 VDD.n4533 VDD.n4174 9.3005
R7220 VDD.n4178 VDD.n4175 9.3005
R7221 VDD.n4179 VDD.n4176 9.3005
R7222 VDD.n4526 VDD.n4180 9.3005
R7223 VDD.n4525 VDD.n4181 9.3005
R7224 VDD.n4524 VDD.n4182 9.3005
R7225 VDD.n4186 VDD.n4183 9.3005
R7226 VDD.n4519 VDD.n4187 9.3005
R7227 VDD.n4518 VDD.n4188 9.3005
R7228 VDD.n4517 VDD.n4189 9.3005
R7229 VDD.n4193 VDD.n4190 9.3005
R7230 VDD.n4512 VDD.n4194 9.3005
R7231 VDD.n4511 VDD.n4195 9.3005
R7232 VDD.n4507 VDD.n4196 9.3005
R7233 VDD.n4200 VDD.n4197 9.3005
R7234 VDD.n4502 VDD.n4201 9.3005
R7235 VDD.n4501 VDD.n4202 9.3005
R7236 VDD.n4500 VDD.n4203 9.3005
R7237 VDD.n4207 VDD.n4204 9.3005
R7238 VDD.n4495 VDD.n4208 9.3005
R7239 VDD.n4494 VDD.n4209 9.3005
R7240 VDD.n4493 VDD.n4210 9.3005
R7241 VDD.n4214 VDD.n4211 9.3005
R7242 VDD.n4488 VDD.n4215 9.3005
R7243 VDD.n4487 VDD.n4216 9.3005
R7244 VDD.n4486 VDD.n4217 9.3005
R7245 VDD.n4221 VDD.n4218 9.3005
R7246 VDD.n4481 VDD.n4222 9.3005
R7247 VDD.n4480 VDD.n4223 9.3005
R7248 VDD.n4479 VDD.n4224 9.3005
R7249 VDD.n4231 VDD.n4229 9.3005
R7250 VDD.n4474 VDD.n4232 9.3005
R7251 VDD.n4473 VDD.n4233 9.3005
R7252 VDD.n4472 VDD.n4234 9.3005
R7253 VDD.n4238 VDD.n4235 9.3005
R7254 VDD.n4467 VDD.n4239 9.3005
R7255 VDD.n4466 VDD.n4240 9.3005
R7256 VDD.n4465 VDD.n4241 9.3005
R7257 VDD.n4245 VDD.n4242 9.3005
R7258 VDD.n4460 VDD.n4246 9.3005
R7259 VDD.n4459 VDD.n4247 9.3005
R7260 VDD.n4458 VDD.n4248 9.3005
R7261 VDD.n4252 VDD.n4249 9.3005
R7262 VDD.n4453 VDD.n4253 9.3005
R7263 VDD.n4452 VDD.n4254 9.3005
R7264 VDD.n4451 VDD.n4255 9.3005
R7265 VDD.n4262 VDD.n4258 9.3005
R7266 VDD.n4446 VDD.n4445 9.3005
R7267 VDD.n4444 VDD.n4261 9.3005
R7268 VDD.n4443 VDD.n4442 9.3005
R7269 VDD.n4264 VDD.n4263 9.3005
R7270 VDD.n4437 VDD.n4267 9.3005
R7271 VDD.n4436 VDD.n4268 9.3005
R7272 VDD.n4435 VDD.n4269 9.3005
R7273 VDD.n4273 VDD.n4270 9.3005
R7274 VDD.n4430 VDD.n4274 9.3005
R7275 VDD.n4429 VDD.n4275 9.3005
R7276 VDD.n4428 VDD.n4276 9.3005
R7277 VDD.n4280 VDD.n4277 9.3005
R7278 VDD.n4423 VDD.n4281 9.3005
R7279 VDD.n4422 VDD.n4282 9.3005
R7280 VDD.n4421 VDD.n4283 9.3005
R7281 VDD.n4290 VDD.n4284 9.3005
R7282 VDD.n4416 VDD.n4415 9.3005
R7283 VDD.n4414 VDD.n4287 9.3005
R7284 VDD.n4413 VDD.n4412 9.3005
R7285 VDD.n4292 VDD.n4291 9.3005
R7286 VDD.n4407 VDD.n4295 9.3005
R7287 VDD.n4406 VDD.n4296 9.3005
R7288 VDD.n4405 VDD.n4297 9.3005
R7289 VDD.n4301 VDD.n4298 9.3005
R7290 VDD.n4400 VDD.n4302 9.3005
R7291 VDD.n4399 VDD.n4303 9.3005
R7292 VDD.n4398 VDD.n4304 9.3005
R7293 VDD.n4308 VDD.n4305 9.3005
R7294 VDD.n4393 VDD.n4309 9.3005
R7295 VDD.n4392 VDD.n4310 9.3005
R7296 VDD.n4391 VDD.n4311 9.3005
R7297 VDD.n4315 VDD.n4312 9.3005
R7298 VDD.n4386 VDD.n4316 9.3005
R7299 VDD.n4385 VDD.n4384 9.3005
R7300 VDD.n4383 VDD.n4319 9.3005
R7301 VDD.n4536 VDD.n4535 9.3005
R7302 VDD.n3973 VDD.n123 9.3005
R7303 VDD.n3975 VDD.n3974 9.3005
R7304 VDD.n112 VDD.n111 9.3005
R7305 VDD.n3988 VDD.n3987 9.3005
R7306 VDD.n3989 VDD.n110 9.3005
R7307 VDD.n3991 VDD.n3990 9.3005
R7308 VDD.n101 VDD.n100 9.3005
R7309 VDD.n4004 VDD.n4003 9.3005
R7310 VDD.n4005 VDD.n99 9.3005
R7311 VDD.n4007 VDD.n4006 9.3005
R7312 VDD.n89 VDD.n88 9.3005
R7313 VDD.n4020 VDD.n4019 9.3005
R7314 VDD.n4021 VDD.n87 9.3005
R7315 VDD.n4023 VDD.n4022 9.3005
R7316 VDD.n77 VDD.n76 9.3005
R7317 VDD.n4036 VDD.n4035 9.3005
R7318 VDD.n4037 VDD.n75 9.3005
R7319 VDD.n4039 VDD.n4038 9.3005
R7320 VDD.n66 VDD.n65 9.3005
R7321 VDD.n4053 VDD.n4052 9.3005
R7322 VDD.n4054 VDD.n64 9.3005
R7323 VDD.n4056 VDD.n4055 9.3005
R7324 VDD.n54 VDD.n53 9.3005
R7325 VDD.n4069 VDD.n4068 9.3005
R7326 VDD.n4070 VDD.n52 9.3005
R7327 VDD.n4072 VDD.n4071 9.3005
R7328 VDD.n42 VDD.n41 9.3005
R7329 VDD.n4085 VDD.n4084 9.3005
R7330 VDD.n4086 VDD.n40 9.3005
R7331 VDD.n4600 VDD.n4087 9.3005
R7332 VDD.n4599 VDD.n4088 9.3005
R7333 VDD.n4598 VDD.n4089 9.3005
R7334 VDD.n4341 VDD.n4090 9.3005
R7335 VDD.n4343 VDD.n4342 9.3005
R7336 VDD.n4344 VDD.n4340 9.3005
R7337 VDD.n4346 VDD.n4345 9.3005
R7338 VDD.n4347 VDD.n4339 9.3005
R7339 VDD.n4349 VDD.n4348 9.3005
R7340 VDD.n4350 VDD.n4337 9.3005
R7341 VDD.n4352 VDD.n4351 9.3005
R7342 VDD.n4353 VDD.n4336 9.3005
R7343 VDD.n4355 VDD.n4354 9.3005
R7344 VDD.n4356 VDD.n4334 9.3005
R7345 VDD.n4358 VDD.n4357 9.3005
R7346 VDD.n4359 VDD.n4333 9.3005
R7347 VDD.n4361 VDD.n4360 9.3005
R7348 VDD.n4362 VDD.n4331 9.3005
R7349 VDD.n4364 VDD.n4363 9.3005
R7350 VDD.n4365 VDD.n4330 9.3005
R7351 VDD.n4367 VDD.n4366 9.3005
R7352 VDD.n4368 VDD.n4328 9.3005
R7353 VDD.n4370 VDD.n4369 9.3005
R7354 VDD.n4371 VDD.n4327 9.3005
R7355 VDD.n4373 VDD.n4372 9.3005
R7356 VDD.n4374 VDD.n4325 9.3005
R7357 VDD.n4376 VDD.n4375 9.3005
R7358 VDD.n4377 VDD.n4324 9.3005
R7359 VDD.n4379 VDD.n4378 9.3005
R7360 VDD.n4380 VDD.n4322 9.3005
R7361 VDD.n4382 VDD.n4381 9.3005
R7362 VDD.n3972 VDD.n3971 9.3005
R7363 VDD.n3800 VDD.n3799 9.3005
R7364 VDD.n3801 VDD.n3791 9.3005
R7365 VDD.n3790 VDD.n3788 9.3005
R7366 VDD.n3807 VDD.n3787 9.3005
R7367 VDD.n3808 VDD.n3786 9.3005
R7368 VDD.n3809 VDD.n3785 9.3005
R7369 VDD.n3784 VDD.n3782 9.3005
R7370 VDD.n3815 VDD.n3781 9.3005
R7371 VDD.n3816 VDD.n3780 9.3005
R7372 VDD.n3817 VDD.n3779 9.3005
R7373 VDD.n3778 VDD.n3776 9.3005
R7374 VDD.n3822 VDD.n3775 9.3005
R7375 VDD.n3823 VDD.n3774 9.3005
R7376 VDD.n3770 VDD.n3769 9.3005
R7377 VDD.n3829 VDD.n3828 9.3005
R7378 VDD.n3830 VDD.n3768 9.3005
R7379 VDD.n3798 VDD.n3797 9.3005
R7380 VDD.n3792 VDD.n124 9.3005
R7381 VDD.n3834 VDD.n3831 9.3005
R7382 VDD.n3835 VDD.n3767 9.3005
R7383 VDD.n3766 VDD.n3764 9.3005
R7384 VDD.n3840 VDD.n3763 9.3005
R7385 VDD.n3850 VDD.n220 9.3005
R7386 VDD.n3851 VDD.n219 9.3005
R7387 VDD.n218 VDD.n216 9.3005
R7388 VDD.n3857 VDD.n215 9.3005
R7389 VDD.n3858 VDD.n214 9.3005
R7390 VDD.n3859 VDD.n213 9.3005
R7391 VDD.n212 VDD.n210 9.3005
R7392 VDD.n3865 VDD.n209 9.3005
R7393 VDD.n3866 VDD.n208 9.3005
R7394 VDD.n2206 VDD.n2205 9.3005
R7395 VDD.n2204 VDD.n1159 9.3005
R7396 VDD.n2203 VDD.n2202 9.3005
R7397 VDD.n2201 VDD.n1166 9.3005
R7398 VDD.n2200 VDD.n2199 9.3005
R7399 VDD.n2198 VDD.n1167 9.3005
R7400 VDD.n2197 VDD.n2196 9.3005
R7401 VDD.n2195 VDD.n1171 9.3005
R7402 VDD.n2194 VDD.n2193 9.3005
R7403 VDD.n2192 VDD.n1172 9.3005
R7404 VDD.n2191 VDD.n2190 9.3005
R7405 VDD.n2189 VDD.n1176 9.3005
R7406 VDD.n2188 VDD.n2187 9.3005
R7407 VDD.n2186 VDD.n1177 9.3005
R7408 VDD.n2185 VDD.n2184 9.3005
R7409 VDD.n2183 VDD.n1181 9.3005
R7410 VDD.n2182 VDD.n2181 9.3005
R7411 VDD.n2180 VDD.n1182 9.3005
R7412 VDD.n2179 VDD.n2178 9.3005
R7413 VDD.n2177 VDD.n1186 9.3005
R7414 VDD.n2176 VDD.n2175 9.3005
R7415 VDD.n1188 VDD.n1187 9.3005
R7416 VDD.n1700 VDD.n1386 9.3005
R7417 VDD.n1702 VDD.n1701 9.3005
R7418 VDD.n1375 VDD.n1374 9.3005
R7419 VDD.n1715 VDD.n1714 9.3005
R7420 VDD.n1716 VDD.n1373 9.3005
R7421 VDD.n1718 VDD.n1717 9.3005
R7422 VDD.n1364 VDD.n1363 9.3005
R7423 VDD.n1731 VDD.n1730 9.3005
R7424 VDD.n1732 VDD.n1362 9.3005
R7425 VDD.n1734 VDD.n1733 9.3005
R7426 VDD.n1352 VDD.n1351 9.3005
R7427 VDD.n1747 VDD.n1746 9.3005
R7428 VDD.n1748 VDD.n1350 9.3005
R7429 VDD.n1750 VDD.n1749 9.3005
R7430 VDD.n1340 VDD.n1339 9.3005
R7431 VDD.n1763 VDD.n1762 9.3005
R7432 VDD.n1764 VDD.n1338 9.3005
R7433 VDD.n1766 VDD.n1765 9.3005
R7434 VDD.n1329 VDD.n1328 9.3005
R7435 VDD.n1780 VDD.n1779 9.3005
R7436 VDD.n1781 VDD.n1327 9.3005
R7437 VDD.n1783 VDD.n1782 9.3005
R7438 VDD.n1317 VDD.n1316 9.3005
R7439 VDD.n1796 VDD.n1795 9.3005
R7440 VDD.n1797 VDD.n1315 9.3005
R7441 VDD.n1799 VDD.n1798 9.3005
R7442 VDD.n1305 VDD.n1304 9.3005
R7443 VDD.n1812 VDD.n1811 9.3005
R7444 VDD.n1813 VDD.n1303 9.3005
R7445 VDD.n1815 VDD.n1814 9.3005
R7446 VDD.n1293 VDD.n1292 9.3005
R7447 VDD.n1842 VDD.n1841 9.3005
R7448 VDD.n1843 VDD.n1291 9.3005
R7449 VDD.n1845 VDD.n1844 9.3005
R7450 VDD.n1281 VDD.n1280 9.3005
R7451 VDD.n1858 VDD.n1857 9.3005
R7452 VDD.n1859 VDD.n1279 9.3005
R7453 VDD.n1861 VDD.n1860 9.3005
R7454 VDD.n1269 VDD.n1268 9.3005
R7455 VDD.n1874 VDD.n1873 9.3005
R7456 VDD.n1875 VDD.n1267 9.3005
R7457 VDD.n1877 VDD.n1876 9.3005
R7458 VDD.n1257 VDD.n1256 9.3005
R7459 VDD.n1890 VDD.n1889 9.3005
R7460 VDD.n1891 VDD.n1255 9.3005
R7461 VDD.n1893 VDD.n1892 9.3005
R7462 VDD.n1245 VDD.n1244 9.3005
R7463 VDD.n1906 VDD.n1905 9.3005
R7464 VDD.n1907 VDD.n1243 9.3005
R7465 VDD.n1909 VDD.n1908 9.3005
R7466 VDD.n1233 VDD.n1232 9.3005
R7467 VDD.n1922 VDD.n1921 9.3005
R7468 VDD.n1923 VDD.n1231 9.3005
R7469 VDD.n1925 VDD.n1924 9.3005
R7470 VDD.n1221 VDD.n1220 9.3005
R7471 VDD.n1938 VDD.n1937 9.3005
R7472 VDD.n1939 VDD.n1218 9.3005
R7473 VDD.n1943 VDD.n1942 9.3005
R7474 VDD.n1941 VDD.n1219 9.3005
R7475 VDD.n1940 VDD.n1208 9.3005
R7476 VDD.n1699 VDD.n1698 9.3005
R7477 VDD.n1560 VDD.n1559 9.3005
R7478 VDD.n1561 VDD.n1548 9.3005
R7479 VDD.n1563 VDD.n1562 9.3005
R7480 VDD.n1564 VDD.n1541 9.3005
R7481 VDD.n1566 VDD.n1565 9.3005
R7482 VDD.n1567 VDD.n1540 9.3005
R7483 VDD.n1569 VDD.n1568 9.3005
R7484 VDD.n1570 VDD.n1533 9.3005
R7485 VDD.n1572 VDD.n1571 9.3005
R7486 VDD.n1573 VDD.n1532 9.3005
R7487 VDD.n1575 VDD.n1574 9.3005
R7488 VDD.n1576 VDD.n1526 9.3005
R7489 VDD.n1578 VDD.n1577 9.3005
R7490 VDD.n1579 VDD.n1525 9.3005
R7491 VDD.n1581 VDD.n1580 9.3005
R7492 VDD.n1521 VDD.n1520 9.3005
R7493 VDD.n1590 VDD.n1519 9.3005
R7494 VDD.n1592 VDD.n1591 9.3005
R7495 VDD.n1593 VDD.n1512 9.3005
R7496 VDD.n1595 VDD.n1594 9.3005
R7497 VDD.n1596 VDD.n1511 9.3005
R7498 VDD.n1598 VDD.n1597 9.3005
R7499 VDD.n1599 VDD.n1504 9.3005
R7500 VDD.n1601 VDD.n1600 9.3005
R7501 VDD.n1602 VDD.n1503 9.3005
R7502 VDD.n1604 VDD.n1603 9.3005
R7503 VDD.n1605 VDD.n1497 9.3005
R7504 VDD.n1607 VDD.n1606 9.3005
R7505 VDD.n1608 VDD.n1495 9.3005
R7506 VDD.n1610 VDD.n1609 9.3005
R7507 VDD.n1496 VDD.n1493 9.3005
R7508 VDD.n1615 VDD.n1492 9.3005
R7509 VDD.n1618 VDD.n1617 9.3005
R7510 VDD.n1619 VDD.n1483 9.3005
R7511 VDD.n1621 VDD.n1620 9.3005
R7512 VDD.n1622 VDD.n1476 9.3005
R7513 VDD.n1624 VDD.n1623 9.3005
R7514 VDD.n1625 VDD.n1475 9.3005
R7515 VDD.n1627 VDD.n1626 9.3005
R7516 VDD.n1628 VDD.n1468 9.3005
R7517 VDD.n1630 VDD.n1629 9.3005
R7518 VDD.n1631 VDD.n1467 9.3005
R7519 VDD.n1633 VDD.n1632 9.3005
R7520 VDD.n1634 VDD.n1460 9.3005
R7521 VDD.n1636 VDD.n1635 9.3005
R7522 VDD.n1637 VDD.n1459 9.3005
R7523 VDD.n1639 VDD.n1638 9.3005
R7524 VDD.n1640 VDD.n1452 9.3005
R7525 VDD.n1645 VDD.n1644 9.3005
R7526 VDD.n1646 VDD.n1451 9.3005
R7527 VDD.n1648 VDD.n1647 9.3005
R7528 VDD.n1649 VDD.n1444 9.3005
R7529 VDD.n1651 VDD.n1650 9.3005
R7530 VDD.n1652 VDD.n1443 9.3005
R7531 VDD.n1654 VDD.n1653 9.3005
R7532 VDD.n1655 VDD.n1436 9.3005
R7533 VDD.n1657 VDD.n1656 9.3005
R7534 VDD.n1658 VDD.n1435 9.3005
R7535 VDD.n1660 VDD.n1659 9.3005
R7536 VDD.n1661 VDD.n1428 9.3005
R7537 VDD.n1663 VDD.n1662 9.3005
R7538 VDD.n1664 VDD.n1427 9.3005
R7539 VDD.n1666 VDD.n1665 9.3005
R7540 VDD.n1667 VDD.n1422 9.3005
R7541 VDD.n1669 VDD.n1668 9.3005
R7542 VDD.n1671 VDD.n1670 9.3005
R7543 VDD.n1672 VDD.n1412 9.3005
R7544 VDD.n1674 VDD.n1673 9.3005
R7545 VDD.n1675 VDD.n1411 9.3005
R7546 VDD.n1677 VDD.n1676 9.3005
R7547 VDD.n1678 VDD.n1404 9.3005
R7548 VDD.n1680 VDD.n1679 9.3005
R7549 VDD.n1681 VDD.n1403 9.3005
R7550 VDD.n1683 VDD.n1682 9.3005
R7551 VDD.n1684 VDD.n1396 9.3005
R7552 VDD.n1686 VDD.n1685 9.3005
R7553 VDD.n1687 VDD.n1395 9.3005
R7554 VDD.n1689 VDD.n1688 9.3005
R7555 VDD.n1690 VDD.n1391 9.3005
R7556 VDD.n1692 VDD.n1691 9.3005
R7557 VDD.n1616 VDD.n1484 9.3005
R7558 VDD.n1589 VDD.n1588 9.3005
R7559 VDD.n1558 VDD.n1549 9.3005
R7560 VDD.n1553 VDD.n1387 9.3005
R7561 VDD.n1382 VDD.n1381 9.3005
R7562 VDD.n1707 VDD.n1706 9.3005
R7563 VDD.n1708 VDD.n1380 9.3005
R7564 VDD.n1710 VDD.n1709 9.3005
R7565 VDD.n1370 VDD.n1369 9.3005
R7566 VDD.n1723 VDD.n1722 9.3005
R7567 VDD.n1724 VDD.n1368 9.3005
R7568 VDD.n1726 VDD.n1725 9.3005
R7569 VDD.n1358 VDD.n1357 9.3005
R7570 VDD.n1739 VDD.n1738 9.3005
R7571 VDD.n1740 VDD.n1356 9.3005
R7572 VDD.n1742 VDD.n1741 9.3005
R7573 VDD.n1346 VDD.n1345 9.3005
R7574 VDD.n1755 VDD.n1754 9.3005
R7575 VDD.n1756 VDD.n1344 9.3005
R7576 VDD.n1758 VDD.n1757 9.3005
R7577 VDD.n1334 VDD.n1333 9.3005
R7578 VDD.n1772 VDD.n1771 9.3005
R7579 VDD.n1773 VDD.n1332 9.3005
R7580 VDD.n1775 VDD.n1774 9.3005
R7581 VDD.n1323 VDD.n1322 9.3005
R7582 VDD.n1788 VDD.n1787 9.3005
R7583 VDD.n1789 VDD.n1321 9.3005
R7584 VDD.n1791 VDD.n1790 9.3005
R7585 VDD.n1311 VDD.n1310 9.3005
R7586 VDD.n1804 VDD.n1803 9.3005
R7587 VDD.n1805 VDD.n1309 9.3005
R7588 VDD.n1807 VDD.n1806 9.3005
R7589 VDD.n1299 VDD.n1298 9.3005
R7590 VDD.n1694 VDD.n1693 9.3005
R7591 VDD.n1834 VDD.n1818 9.3005
R7592 VDD.n15 VDD.n14 8.55753
R7593 VDD.n4605 VDD.n4604 8.07387
R7594 VDD.n1834 VDD.n1833 8.07387
R7595 VDD.n1378 VDD.t34 8.07295
R7596 VDD.t42 VDD.n1223 8.07295
R7597 VDD.n115 VDD.t50 8.07295
R7598 VDD.t38 VDD.n4549 8.07295
R7599 VDD.n1558 VDD.n1553 7.75808
R7600 VDD.n2175 VDD.n1188 7.75808
R7601 VDD.n3797 VDD.n3792 7.75808
R7602 VDD.n4385 VDD.n4319 7.75808
R7603 VDD.n1777 VDD.t11 7.43565
R7604 VDD.n1871 VDD.t2 7.43565
R7605 VDD.n4050 VDD.t4 7.43565
R7606 VDD.n4580 VDD.t9 7.43565
R7607 VDD.n2470 VDD.n974 7.22322
R7608 VDD.n2470 VDD.n968 7.22322
R7609 VDD.n2476 VDD.n968 7.22322
R7610 VDD.n2476 VDD.n962 7.22322
R7611 VDD.n2482 VDD.n962 7.22322
R7612 VDD.n2482 VDD.n956 7.22322
R7613 VDD.n2488 VDD.n956 7.22322
R7614 VDD.n2488 VDD.n950 7.22322
R7615 VDD.n2494 VDD.n950 7.22322
R7616 VDD.n2500 VDD.n939 7.22322
R7617 VDD.n2506 VDD.n939 7.22322
R7618 VDD.n2506 VDD.n933 7.22322
R7619 VDD.n2512 VDD.n933 7.22322
R7620 VDD.n2512 VDD.n927 7.22322
R7621 VDD.n2518 VDD.n927 7.22322
R7622 VDD.n2518 VDD.n921 7.22322
R7623 VDD.n2524 VDD.n921 7.22322
R7624 VDD.n2524 VDD.n915 7.22322
R7625 VDD.n2530 VDD.n915 7.22322
R7626 VDD.n2530 VDD.n909 7.22322
R7627 VDD.n2536 VDD.n909 7.22322
R7628 VDD.n2536 VDD.n902 7.22322
R7629 VDD.n2542 VDD.n902 7.22322
R7630 VDD.n2542 VDD.n905 7.22322
R7631 VDD.n2548 VDD.n891 7.22322
R7632 VDD.n2554 VDD.n891 7.22322
R7633 VDD.n2554 VDD.n885 7.22322
R7634 VDD.n2560 VDD.n885 7.22322
R7635 VDD.n2566 VDD.n879 7.22322
R7636 VDD.n2566 VDD.n873 7.22322
R7637 VDD.n2572 VDD.n873 7.22322
R7638 VDD.n2572 VDD.n867 7.22322
R7639 VDD.n2578 VDD.n867 7.22322
R7640 VDD.n2578 VDD.n861 7.22322
R7641 VDD.n2584 VDD.n861 7.22322
R7642 VDD.n2584 VDD.n855 7.22322
R7643 VDD.n2590 VDD.n855 7.22322
R7644 VDD.n2590 VDD.n849 7.22322
R7645 VDD.n2596 VDD.n849 7.22322
R7646 VDD.n2596 VDD.n843 7.22322
R7647 VDD.n2602 VDD.n843 7.22322
R7648 VDD.n2602 VDD.n837 7.22322
R7649 VDD.n2608 VDD.n837 7.22322
R7650 VDD.n2608 VDD.n831 7.22322
R7651 VDD.n2614 VDD.n831 7.22322
R7652 VDD.n2620 VDD.n824 7.22322
R7653 VDD.n2620 VDD.n827 7.22322
R7654 VDD.n2626 VDD.n813 7.22322
R7655 VDD.n2632 VDD.n813 7.22322
R7656 VDD.n2632 VDD.n807 7.22322
R7657 VDD.n2638 VDD.n807 7.22322
R7658 VDD.n2638 VDD.n801 7.22322
R7659 VDD.n2644 VDD.n801 7.22322
R7660 VDD.n2644 VDD.n795 7.22322
R7661 VDD.n2650 VDD.n795 7.22322
R7662 VDD.n2650 VDD.n789 7.22322
R7663 VDD.n2656 VDD.n789 7.22322
R7664 VDD.n2656 VDD.n782 7.22322
R7665 VDD.n2662 VDD.n782 7.22322
R7666 VDD.n2662 VDD.n785 7.22322
R7667 VDD.n2668 VDD.n770 7.22322
R7668 VDD.n2674 VDD.n770 7.22322
R7669 VDD.n2674 VDD.n773 7.22322
R7670 VDD.n2680 VDD.n759 7.22322
R7671 VDD.n2686 VDD.n759 7.22322
R7672 VDD.n2686 VDD.n753 7.22322
R7673 VDD.n2692 VDD.n753 7.22322
R7674 VDD.n2692 VDD.n747 7.22322
R7675 VDD.n2698 VDD.n747 7.22322
R7676 VDD.n2698 VDD.n741 7.22322
R7677 VDD.n2704 VDD.n741 7.22322
R7678 VDD.n2704 VDD.n735 7.22322
R7679 VDD.n2710 VDD.n735 7.22322
R7680 VDD.n2710 VDD.n728 7.22322
R7681 VDD.n2716 VDD.n728 7.22322
R7682 VDD.n2716 VDD.n731 7.22322
R7683 VDD.n2722 VDD.n717 7.22322
R7684 VDD.n2728 VDD.n717 7.22322
R7685 VDD.n2734 VDD.n711 7.22322
R7686 VDD.n2734 VDD.n705 7.22322
R7687 VDD.n2740 VDD.n705 7.22322
R7688 VDD.n2740 VDD.n699 7.22322
R7689 VDD.n2746 VDD.n699 7.22322
R7690 VDD.n2746 VDD.n693 7.22322
R7691 VDD.n2752 VDD.n693 7.22322
R7692 VDD.n2752 VDD.n687 7.22322
R7693 VDD.n2758 VDD.n687 7.22322
R7694 VDD.n2758 VDD.n681 7.22322
R7695 VDD.n2764 VDD.n681 7.22322
R7696 VDD.n2764 VDD.n675 7.22322
R7697 VDD.n2770 VDD.n675 7.22322
R7698 VDD.n2770 VDD.n669 7.22322
R7699 VDD.n2776 VDD.n669 7.22322
R7700 VDD.n2776 VDD.n663 7.22322
R7701 VDD.n2782 VDD.n663 7.22322
R7702 VDD.n2788 VDD.n657 7.22322
R7703 VDD.n2788 VDD.n651 7.22322
R7704 VDD.n2794 VDD.n651 7.22322
R7705 VDD.n2794 VDD.n644 7.22322
R7706 VDD.n2805 VDD.n644 7.22322
R7707 VDD.n2805 VDD.n638 7.22322
R7708 VDD.n2811 VDD.n638 7.22322
R7709 VDD.n2811 VDD.n628 7.22322
R7710 VDD.n2857 VDD.n628 7.22322
R7711 VDD.n2857 VDD.n602 7.22322
R7712 VDD.n3335 VDD.n596 7.22322
R7713 VDD.n3341 VDD.n596 7.22322
R7714 VDD.n3341 VDD.n590 7.22322
R7715 VDD.n3347 VDD.n590 7.22322
R7716 VDD.n3347 VDD.n584 7.22322
R7717 VDD.n3353 VDD.n584 7.22322
R7718 VDD.n3353 VDD.n578 7.22322
R7719 VDD.n3359 VDD.n578 7.22322
R7720 VDD.n3359 VDD.n572 7.22322
R7721 VDD.n3365 VDD.n572 7.22322
R7722 VDD.n3371 VDD.n566 7.22322
R7723 VDD.n3371 VDD.n560 7.22322
R7724 VDD.n3377 VDD.n560 7.22322
R7725 VDD.n3377 VDD.n554 7.22322
R7726 VDD.n3383 VDD.n554 7.22322
R7727 VDD.n3383 VDD.n548 7.22322
R7728 VDD.n3389 VDD.n548 7.22322
R7729 VDD.n3389 VDD.n542 7.22322
R7730 VDD.n3395 VDD.n542 7.22322
R7731 VDD.n3395 VDD.n536 7.22322
R7732 VDD.n3401 VDD.n536 7.22322
R7733 VDD.n3401 VDD.n530 7.22322
R7734 VDD.n3407 VDD.n530 7.22322
R7735 VDD.n3407 VDD.n524 7.22322
R7736 VDD.n3413 VDD.n524 7.22322
R7737 VDD.n3413 VDD.n518 7.22322
R7738 VDD.n3419 VDD.n518 7.22322
R7739 VDD.n3425 VDD.n511 7.22322
R7740 VDD.n3425 VDD.n514 7.22322
R7741 VDD.n3431 VDD.n500 7.22322
R7742 VDD.n3437 VDD.n500 7.22322
R7743 VDD.n3437 VDD.n494 7.22322
R7744 VDD.n3443 VDD.n494 7.22322
R7745 VDD.n3443 VDD.n488 7.22322
R7746 VDD.n3449 VDD.n488 7.22322
R7747 VDD.n3449 VDD.n482 7.22322
R7748 VDD.n3455 VDD.n482 7.22322
R7749 VDD.n3455 VDD.n476 7.22322
R7750 VDD.n3461 VDD.n476 7.22322
R7751 VDD.n3461 VDD.n469 7.22322
R7752 VDD.n3467 VDD.n469 7.22322
R7753 VDD.n3467 VDD.n472 7.22322
R7754 VDD.n3473 VDD.n457 7.22322
R7755 VDD.n3479 VDD.n457 7.22322
R7756 VDD.n3479 VDD.n460 7.22322
R7757 VDD.n3485 VDD.n446 7.22322
R7758 VDD.n3491 VDD.n446 7.22322
R7759 VDD.n3491 VDD.n440 7.22322
R7760 VDD.n3497 VDD.n440 7.22322
R7761 VDD.n3497 VDD.n434 7.22322
R7762 VDD.n3503 VDD.n434 7.22322
R7763 VDD.n3503 VDD.n428 7.22322
R7764 VDD.n3509 VDD.n428 7.22322
R7765 VDD.n3509 VDD.n422 7.22322
R7766 VDD.n3515 VDD.n422 7.22322
R7767 VDD.n3515 VDD.n415 7.22322
R7768 VDD.n3521 VDD.n415 7.22322
R7769 VDD.n3521 VDD.n418 7.22322
R7770 VDD.n3527 VDD.n404 7.22322
R7771 VDD.n3533 VDD.n404 7.22322
R7772 VDD.n3539 VDD.n398 7.22322
R7773 VDD.n3539 VDD.n392 7.22322
R7774 VDD.n3545 VDD.n392 7.22322
R7775 VDD.n3545 VDD.n386 7.22322
R7776 VDD.n3551 VDD.n386 7.22322
R7777 VDD.n3551 VDD.n380 7.22322
R7778 VDD.n3557 VDD.n380 7.22322
R7779 VDD.n3557 VDD.n374 7.22322
R7780 VDD.n3563 VDD.n374 7.22322
R7781 VDD.n3563 VDD.n368 7.22322
R7782 VDD.n3569 VDD.n368 7.22322
R7783 VDD.n3569 VDD.n362 7.22322
R7784 VDD.n3575 VDD.n362 7.22322
R7785 VDD.n3575 VDD.n356 7.22322
R7786 VDD.n3581 VDD.n356 7.22322
R7787 VDD.n3581 VDD.n350 7.22322
R7788 VDD.n3587 VDD.n350 7.22322
R7789 VDD.n3593 VDD.n344 7.22322
R7790 VDD.n3593 VDD.n337 7.22322
R7791 VDD.n3599 VDD.n337 7.22322
R7792 VDD.n3599 VDD.n340 7.22322
R7793 VDD.n3605 VDD.n326 7.22322
R7794 VDD.n3611 VDD.n326 7.22322
R7795 VDD.n3611 VDD.n320 7.22322
R7796 VDD.n3617 VDD.n320 7.22322
R7797 VDD.n3617 VDD.n314 7.22322
R7798 VDD.n3623 VDD.n314 7.22322
R7799 VDD.n3623 VDD.n308 7.22322
R7800 VDD.n3629 VDD.n308 7.22322
R7801 VDD.n3629 VDD.n302 7.22322
R7802 VDD.n3635 VDD.n302 7.22322
R7803 VDD.n3635 VDD.n296 7.22322
R7804 VDD.n3641 VDD.n296 7.22322
R7805 VDD.n3641 VDD.n289 7.22322
R7806 VDD.n3647 VDD.n289 7.22322
R7807 VDD.n3647 VDD.n292 7.22322
R7808 VDD.n3659 VDD.n278 7.22322
R7809 VDD.n3659 VDD.n272 7.22322
R7810 VDD.n3665 VDD.n272 7.22322
R7811 VDD.n3665 VDD.n265 7.22322
R7812 VDD.n3697 VDD.n265 7.22322
R7813 VDD.n3697 VDD.n259 7.22322
R7814 VDD.n3703 VDD.n259 7.22322
R7815 VDD.n3703 VDD.n238 7.22322
R7816 VDD.n3743 VDD.n238 7.22322
R7817 VDD.n1588 VDD.n1521 7.17626
R7818 VDD.n2199 VDD.n1166 7.17626
R7819 VDD.n3834 VDD.n3768 7.17626
R7820 VDD.n4416 VDD.n4287 7.17626
R7821 VDD.n2680 VDD.t135 7.117
R7822 VDD.n472 VDD.t153 7.117
R7823 VDD.n2500 VDD.t46 6.69214
R7824 VDD.n292 VDD.t30 6.69214
R7825 VDD.n1823 VDD.n1820 6.62622
R7826 VDD.n1616 VDD.n1615 6.59444
R7827 VDD.n2077 VDD.n2037 6.59444
R7828 VDD.n4446 VDD.n4258 6.59444
R7829 VDD.n3867 VDD.n3866 6.59444
R7830 VDD.n2415 VDD.t139 6.58592
R7831 VDD.t125 VDD.t82 6.58592
R7832 VDD.t69 VDD.t149 6.58592
R7833 VDD.n3653 VDD.t151 6.58592
R7834 VDD.n1643 VDD.n1640 6.01262
R7835 VDD.n2008 VDD.n2006 6.01262
R7836 VDD.n4229 VDD.n4227 6.01262
R7837 VDD.n3899 VDD.n179 6.01262
R7838 VDD.n20 VDD.n17 5.85754
R7839 VDD.n1668 VDD.n1421 5.4308
R7840 VDD.n2138 VDD.n1977 5.4308
R7841 VDD.n4510 VDD.n4507 5.4308
R7842 VDD.n3935 VDD.n3934 5.4308
R7843 VDD.n2560 VDD.t124 5.41754
R7844 VDD.t141 VDD.n824 5.41754
R7845 VDD.n785 VDD.t146 5.41754
R7846 VDD.n2722 VDD.t130 5.41754
R7847 VDD.n514 VDD.t122 5.41754
R7848 VDD.n3485 VDD.t121 5.41754
R7849 VDD.n3533 VDD.t123 5.41754
R7850 VDD.t127 VDD.n344 5.41754
R7851 VDD.n1832 VDD.n1831 5.40711
R7852 VDD.n1829 VDD.n1828 5.40711
R7853 VDD.n1826 VDD.n1825 5.40711
R7854 VDD.n1823 VDD.n1822 5.40711
R7855 VDD.n2451 VDD.n999 5.30782
R7856 VDD.n2448 VDD.n999 5.30782
R7857 VDD.n3726 VDD.n164 5.30782
R7858 VDD.n3722 VDD.n164 5.30782
R7859 VDD.n3761 VDD.n225 5.30782
R7860 VDD.n3761 VDD.n3760 5.30782
R7861 VDD.n2224 VDD.n2208 5.30782
R7862 VDD.n2227 VDD.n2208 5.30782
R7863 VDD.n2060 VDD.n1157 4.74817
R7864 VDD.n2055 VDD.n1158 4.74817
R7865 VDD.n1992 VDD.n1989 4.74817
R7866 VDD.n2123 VDD.n2122 4.74817
R7867 VDD.n2124 VDD.n1992 4.74817
R7868 VDD.n2122 VDD.n1993 4.74817
R7869 VDD.n3919 VDD.n3918 4.74817
R7870 VDD.n3915 VDD.n3914 4.74817
R7871 VDD.n3915 VDD.n165 4.74817
R7872 VDD.n3918 VDD.n162 4.74817
R7873 VDD.n3845 VDD.n221 4.74817
R7874 VDD.n3841 VDD.n223 4.74817
R7875 VDD.n3844 VDD.n223 4.74817
R7876 VDD.n3849 VDD.n221 4.74817
R7877 VDD.n2056 VDD.n1157 4.74817
R7878 VDD.n1160 VDD.n1158 4.74817
R7879 VDD.n29 VDD.n28 4.63843
R7880 VDD.n26 VDD.n25 4.63843
R7881 VDD.n23 VDD.n22 4.63843
R7882 VDD.n20 VDD.n19 4.63843
R7883 VDD.n4605 VDD.n29 4.32081
R7884 VDD.n1833 VDD.n1832 4.32081
R7885 VDD.n905 VDD.t142 4.24916
R7886 VDD.n3605 VDD.t155 4.24916
R7887 VDD.n827 VDD.t157 3.71808
R7888 VDD.n2728 VDD.t128 3.71808
R7889 VDD.t144 VDD.n511 3.71808
R7890 VDD.n3527 VDD.t147 3.71808
R7891 VDD.n2626 VDD.t157 3.50564
R7892 VDD.t128 VDD.n711 3.50564
R7893 VDD.n3419 VDD.t144 3.50564
R7894 VDD.n418 VDD.t147 3.50564
R7895 VDD.n1768 VDD.t11 3.18699
R7896 VDD.t2 VDD.n1265 3.18699
R7897 VDD.n4041 VDD.t4 3.18699
R7898 VDD.n4120 VDD.t9 3.18699
R7899 VDD.n2548 VDD.t142 2.97456
R7900 VDD.n340 VDD.t155 2.97456
R7901 VDD.n1720 VDD.t34 2.5497
R7902 VDD.n1927 VDD.t42 2.5497
R7903 VDD.n3993 VDD.t50 2.5497
R7904 VDD.n4550 VDD.t38 2.5497
R7905 VDD.n1833 VDD.n15 2.51234
R7906 VDD VDD.n4605 2.5045
R7907 VDD.n2121 VDD.n1992 2.27742
R7908 VDD.n2122 VDD.n2121 2.27742
R7909 VDD.n3917 VDD.n3915 2.27742
R7910 VDD.n3918 VDD.n3917 2.27742
R7911 VDD.n3762 VDD.n223 2.27742
R7912 VDD.n3762 VDD.n221 2.27742
R7913 VDD.n2207 VDD.n1157 2.27742
R7914 VDD.n2207 VDD.n1158 2.27742
R7915 VDD.n4 VDD.n2 2.12191
R7916 VDD.n11 VDD.n9 2.12191
R7917 VDD.t124 VDD.n879 1.80618
R7918 VDD.n2614 VDD.t141 1.80618
R7919 VDD.n2668 VDD.t146 1.80618
R7920 VDD.n731 VDD.t130 1.80618
R7921 VDD.n3431 VDD.t122 1.80618
R7922 VDD.n460 VDD.t121 1.80618
R7923 VDD.t123 VDD.n398 1.80618
R7924 VDD.n3587 VDD.t127 1.80618
R7925 VDD.n6 VDD.n4 1.71027
R7926 VDD.n13 VDD.n11 1.71027
R7927 VDD.n14 VDD.n6 1.32665
R7928 VDD.n14 VDD.n13 1.32665
R7929 VDD.n29 VDD.n26 1.21961
R7930 VDD.n26 VDD.n23 1.21961
R7931 VDD.n23 VDD.n20 1.21961
R7932 VDD.n1832 VDD.n1829 1.21961
R7933 VDD.n1829 VDD.n1826 1.21961
R7934 VDD.n1826 VDD.n1823 1.21961
R7935 VDD.n1671 VDD.n1421 1.16414
R7936 VDD.n1977 VDD.n1972 1.16414
R7937 VDD.n4511 VDD.n4510 1.16414
R7938 VDD.n3936 VDD.n3935 1.16414
R7939 VDD.n2494 VDD.t139 0.637799
R7940 VDD.t151 VDD.n278 0.637799
R7941 VDD.n1644 VDD.n1643 0.582318
R7942 VDD.n2110 VDD.n2006 0.582318
R7943 VDD.n4479 VDD.n4227 0.582318
R7944 VDD.n179 VDD.n175 0.582318
R7945 VDD.n2415 VDD.t46 0.531582
R7946 VDD.t82 VDD.n657 0.531582
R7947 VDD.n3365 VDD.t69 0.531582
R7948 VDD.n3653 VDD.t30 0.531582
R7949 VDD.n2167 VDD.n2166 0.495927
R7950 VDD.n3966 VDD.n3965 0.495927
R7951 VDD.n4537 VDD.n4536 0.495927
R7952 VDD.n4383 VDD.n4382 0.495927
R7953 VDD.n3972 VDD.n124 0.495927
R7954 VDD.n1940 VDD.n1187 0.495927
R7955 VDD.n1699 VDD.n1387 0.495927
R7956 VDD.n1693 VDD.n1692 0.495927
R7957 VDD.n1836 VDD.n1835 0.152939
R7958 VDD.n1836 VDD.n1286 0.152939
R7959 VDD.n1850 VDD.n1286 0.152939
R7960 VDD.n1851 VDD.n1850 0.152939
R7961 VDD.n1852 VDD.n1851 0.152939
R7962 VDD.n1852 VDD.n1274 0.152939
R7963 VDD.n1866 VDD.n1274 0.152939
R7964 VDD.n1867 VDD.n1866 0.152939
R7965 VDD.n1868 VDD.n1867 0.152939
R7966 VDD.n1868 VDD.n1262 0.152939
R7967 VDD.n1882 VDD.n1262 0.152939
R7968 VDD.n1883 VDD.n1882 0.152939
R7969 VDD.n1884 VDD.n1883 0.152939
R7970 VDD.n1884 VDD.n1250 0.152939
R7971 VDD.n1898 VDD.n1250 0.152939
R7972 VDD.n1899 VDD.n1898 0.152939
R7973 VDD.n1900 VDD.n1899 0.152939
R7974 VDD.n1900 VDD.n1238 0.152939
R7975 VDD.n1914 VDD.n1238 0.152939
R7976 VDD.n1915 VDD.n1914 0.152939
R7977 VDD.n1916 VDD.n1915 0.152939
R7978 VDD.n1916 VDD.n1226 0.152939
R7979 VDD.n1930 VDD.n1226 0.152939
R7980 VDD.n1931 VDD.n1930 0.152939
R7981 VDD.n1932 VDD.n1931 0.152939
R7982 VDD.n1932 VDD.n1213 0.152939
R7983 VDD.n1948 VDD.n1213 0.152939
R7984 VDD.n1949 VDD.n1948 0.152939
R7985 VDD.n2167 VDD.n1949 0.152939
R7986 VDD.n2166 VDD.n1950 0.152939
R7987 VDD.n1954 VDD.n1950 0.152939
R7988 VDD.n1955 VDD.n1954 0.152939
R7989 VDD.n1956 VDD.n1955 0.152939
R7990 VDD.n1957 VDD.n1956 0.152939
R7991 VDD.n1961 VDD.n1957 0.152939
R7992 VDD.n1962 VDD.n1961 0.152939
R7993 VDD.n1963 VDD.n1962 0.152939
R7994 VDD.n1964 VDD.n1963 0.152939
R7995 VDD.n1968 VDD.n1964 0.152939
R7996 VDD.n1969 VDD.n1968 0.152939
R7997 VDD.n1970 VDD.n1969 0.152939
R7998 VDD.n1971 VDD.n1970 0.152939
R7999 VDD.n1978 VDD.n1971 0.152939
R8000 VDD.n1979 VDD.n1978 0.152939
R8001 VDD.n1980 VDD.n1979 0.152939
R8002 VDD.n1981 VDD.n1980 0.152939
R8003 VDD.n1985 VDD.n1981 0.152939
R8004 VDD.n1986 VDD.n1985 0.152939
R8005 VDD.n1987 VDD.n1986 0.152939
R8006 VDD.n1988 VDD.n1987 0.152939
R8007 VDD.n2120 VDD.n1994 0.152939
R8008 VDD.n2000 VDD.n1994 0.152939
R8009 VDD.n2001 VDD.n2000 0.152939
R8010 VDD.n2002 VDD.n2001 0.152939
R8011 VDD.n2003 VDD.n2002 0.152939
R8012 VDD.n2010 VDD.n2003 0.152939
R8013 VDD.n2011 VDD.n2010 0.152939
R8014 VDD.n2012 VDD.n2011 0.152939
R8015 VDD.n2013 VDD.n2012 0.152939
R8016 VDD.n2017 VDD.n2013 0.152939
R8017 VDD.n2018 VDD.n2017 0.152939
R8018 VDD.n2019 VDD.n2018 0.152939
R8019 VDD.n2020 VDD.n2019 0.152939
R8020 VDD.n2024 VDD.n2020 0.152939
R8021 VDD.n2025 VDD.n2024 0.152939
R8022 VDD.n2026 VDD.n2025 0.152939
R8023 VDD.n2027 VDD.n2026 0.152939
R8024 VDD.n2031 VDD.n2027 0.152939
R8025 VDD.n2032 VDD.n2031 0.152939
R8026 VDD.n2033 VDD.n2032 0.152939
R8027 VDD.n2034 VDD.n2033 0.152939
R8028 VDD.n2041 VDD.n2034 0.152939
R8029 VDD.n2076 VDD.n2041 0.152939
R8030 VDD.n2076 VDD.n2075 0.152939
R8031 VDD.n2075 VDD.n2074 0.152939
R8032 VDD.n2074 VDD.n2042 0.152939
R8033 VDD.n2046 VDD.n2042 0.152939
R8034 VDD.n2047 VDD.n2046 0.152939
R8035 VDD.n2048 VDD.n2047 0.152939
R8036 VDD.n2049 VDD.n2048 0.152939
R8037 VDD.n2049 VDD.n1156 0.152939
R8038 VDD.n171 VDD.n163 0.152939
R8039 VDD.n172 VDD.n171 0.152939
R8040 VDD.n173 VDD.n172 0.152939
R8041 VDD.n174 VDD.n173 0.152939
R8042 VDD.n180 VDD.n174 0.152939
R8043 VDD.n181 VDD.n180 0.152939
R8044 VDD.n182 VDD.n181 0.152939
R8045 VDD.n183 VDD.n182 0.152939
R8046 VDD.n186 VDD.n183 0.152939
R8047 VDD.n187 VDD.n186 0.152939
R8048 VDD.n188 VDD.n187 0.152939
R8049 VDD.n189 VDD.n188 0.152939
R8050 VDD.n192 VDD.n189 0.152939
R8051 VDD.n193 VDD.n192 0.152939
R8052 VDD.n194 VDD.n193 0.152939
R8053 VDD.n195 VDD.n194 0.152939
R8054 VDD.n198 VDD.n195 0.152939
R8055 VDD.n199 VDD.n198 0.152939
R8056 VDD.n200 VDD.n199 0.152939
R8057 VDD.n201 VDD.n200 0.152939
R8058 VDD.n204 VDD.n201 0.152939
R8059 VDD.n205 VDD.n204 0.152939
R8060 VDD.n208 VDD.n205 0.152939
R8061 VDD.n209 VDD.n208 0.152939
R8062 VDD.n212 VDD.n209 0.152939
R8063 VDD.n213 VDD.n212 0.152939
R8064 VDD.n214 VDD.n213 0.152939
R8065 VDD.n215 VDD.n214 0.152939
R8066 VDD.n218 VDD.n215 0.152939
R8067 VDD.n219 VDD.n218 0.152939
R8068 VDD.n220 VDD.n219 0.152939
R8069 VDD.n3965 VDD.n128 0.152939
R8070 VDD.n131 VDD.n128 0.152939
R8071 VDD.n132 VDD.n131 0.152939
R8072 VDD.n133 VDD.n132 0.152939
R8073 VDD.n136 VDD.n133 0.152939
R8074 VDD.n137 VDD.n136 0.152939
R8075 VDD.n138 VDD.n137 0.152939
R8076 VDD.n139 VDD.n138 0.152939
R8077 VDD.n142 VDD.n139 0.152939
R8078 VDD.n143 VDD.n142 0.152939
R8079 VDD.n144 VDD.n143 0.152939
R8080 VDD.n145 VDD.n144 0.152939
R8081 VDD.n148 VDD.n145 0.152939
R8082 VDD.n149 VDD.n148 0.152939
R8083 VDD.n152 VDD.n149 0.152939
R8084 VDD.n153 VDD.n152 0.152939
R8085 VDD.n156 VDD.n153 0.152939
R8086 VDD.n157 VDD.n156 0.152939
R8087 VDD.n158 VDD.n157 0.152939
R8088 VDD.n159 VDD.n158 0.152939
R8089 VDD.n3916 VDD.n159 0.152939
R8090 VDD.n3966 VDD.n118 0.152939
R8091 VDD.n3980 VDD.n118 0.152939
R8092 VDD.n3981 VDD.n3980 0.152939
R8093 VDD.n3982 VDD.n3981 0.152939
R8094 VDD.n3982 VDD.n106 0.152939
R8095 VDD.n3996 VDD.n106 0.152939
R8096 VDD.n3997 VDD.n3996 0.152939
R8097 VDD.n3998 VDD.n3997 0.152939
R8098 VDD.n3998 VDD.n94 0.152939
R8099 VDD.n4012 VDD.n94 0.152939
R8100 VDD.n4013 VDD.n4012 0.152939
R8101 VDD.n4014 VDD.n4013 0.152939
R8102 VDD.n4014 VDD.n82 0.152939
R8103 VDD.n4028 VDD.n82 0.152939
R8104 VDD.n4029 VDD.n4028 0.152939
R8105 VDD.n4030 VDD.n4029 0.152939
R8106 VDD.n4030 VDD.n70 0.152939
R8107 VDD.n4045 VDD.n70 0.152939
R8108 VDD.n4046 VDD.n4045 0.152939
R8109 VDD.n4047 VDD.n4046 0.152939
R8110 VDD.n4047 VDD.n59 0.152939
R8111 VDD.n4061 VDD.n59 0.152939
R8112 VDD.n4062 VDD.n4061 0.152939
R8113 VDD.n4063 VDD.n4062 0.152939
R8114 VDD.n4063 VDD.n47 0.152939
R8115 VDD.n4077 VDD.n47 0.152939
R8116 VDD.n4078 VDD.n4077 0.152939
R8117 VDD.n4079 VDD.n4078 0.152939
R8118 VDD.n4079 VDD.n30 0.152939
R8119 VDD.n4094 VDD.n31 0.152939
R8120 VDD.n4095 VDD.n4094 0.152939
R8121 VDD.n4096 VDD.n4095 0.152939
R8122 VDD.n4104 VDD.n4096 0.152939
R8123 VDD.n4105 VDD.n4104 0.152939
R8124 VDD.n4106 VDD.n4105 0.152939
R8125 VDD.n4107 VDD.n4106 0.152939
R8126 VDD.n4114 VDD.n4107 0.152939
R8127 VDD.n4115 VDD.n4114 0.152939
R8128 VDD.n4116 VDD.n4115 0.152939
R8129 VDD.n4117 VDD.n4116 0.152939
R8130 VDD.n4126 VDD.n4117 0.152939
R8131 VDD.n4127 VDD.n4126 0.152939
R8132 VDD.n4128 VDD.n4127 0.152939
R8133 VDD.n4129 VDD.n4128 0.152939
R8134 VDD.n4137 VDD.n4129 0.152939
R8135 VDD.n4138 VDD.n4137 0.152939
R8136 VDD.n4139 VDD.n4138 0.152939
R8137 VDD.n4140 VDD.n4139 0.152939
R8138 VDD.n4148 VDD.n4140 0.152939
R8139 VDD.n4149 VDD.n4148 0.152939
R8140 VDD.n4150 VDD.n4149 0.152939
R8141 VDD.n4151 VDD.n4150 0.152939
R8142 VDD.n4159 VDD.n4151 0.152939
R8143 VDD.n4160 VDD.n4159 0.152939
R8144 VDD.n4161 VDD.n4160 0.152939
R8145 VDD.n4162 VDD.n4161 0.152939
R8146 VDD.n4170 VDD.n4162 0.152939
R8147 VDD.n4537 VDD.n4170 0.152939
R8148 VDD.n4536 VDD.n4171 0.152939
R8149 VDD.n4174 VDD.n4171 0.152939
R8150 VDD.n4178 VDD.n4174 0.152939
R8151 VDD.n4179 VDD.n4178 0.152939
R8152 VDD.n4180 VDD.n4179 0.152939
R8153 VDD.n4181 VDD.n4180 0.152939
R8154 VDD.n4182 VDD.n4181 0.152939
R8155 VDD.n4186 VDD.n4182 0.152939
R8156 VDD.n4187 VDD.n4186 0.152939
R8157 VDD.n4188 VDD.n4187 0.152939
R8158 VDD.n4189 VDD.n4188 0.152939
R8159 VDD.n4193 VDD.n4189 0.152939
R8160 VDD.n4194 VDD.n4193 0.152939
R8161 VDD.n4195 VDD.n4194 0.152939
R8162 VDD.n4196 VDD.n4195 0.152939
R8163 VDD.n4200 VDD.n4196 0.152939
R8164 VDD.n4201 VDD.n4200 0.152939
R8165 VDD.n4202 VDD.n4201 0.152939
R8166 VDD.n4203 VDD.n4202 0.152939
R8167 VDD.n4207 VDD.n4203 0.152939
R8168 VDD.n4208 VDD.n4207 0.152939
R8169 VDD.n4209 VDD.n4208 0.152939
R8170 VDD.n4210 VDD.n4209 0.152939
R8171 VDD.n4214 VDD.n4210 0.152939
R8172 VDD.n4215 VDD.n4214 0.152939
R8173 VDD.n4216 VDD.n4215 0.152939
R8174 VDD.n4217 VDD.n4216 0.152939
R8175 VDD.n4221 VDD.n4217 0.152939
R8176 VDD.n4222 VDD.n4221 0.152939
R8177 VDD.n4223 VDD.n4222 0.152939
R8178 VDD.n4224 VDD.n4223 0.152939
R8179 VDD.n4231 VDD.n4224 0.152939
R8180 VDD.n4232 VDD.n4231 0.152939
R8181 VDD.n4233 VDD.n4232 0.152939
R8182 VDD.n4234 VDD.n4233 0.152939
R8183 VDD.n4238 VDD.n4234 0.152939
R8184 VDD.n4239 VDD.n4238 0.152939
R8185 VDD.n4240 VDD.n4239 0.152939
R8186 VDD.n4241 VDD.n4240 0.152939
R8187 VDD.n4245 VDD.n4241 0.152939
R8188 VDD.n4246 VDD.n4245 0.152939
R8189 VDD.n4247 VDD.n4246 0.152939
R8190 VDD.n4248 VDD.n4247 0.152939
R8191 VDD.n4252 VDD.n4248 0.152939
R8192 VDD.n4253 VDD.n4252 0.152939
R8193 VDD.n4254 VDD.n4253 0.152939
R8194 VDD.n4255 VDD.n4254 0.152939
R8195 VDD.n4262 VDD.n4255 0.152939
R8196 VDD.n4445 VDD.n4262 0.152939
R8197 VDD.n4445 VDD.n4444 0.152939
R8198 VDD.n4444 VDD.n4443 0.152939
R8199 VDD.n4443 VDD.n4263 0.152939
R8200 VDD.n4267 VDD.n4263 0.152939
R8201 VDD.n4268 VDD.n4267 0.152939
R8202 VDD.n4269 VDD.n4268 0.152939
R8203 VDD.n4273 VDD.n4269 0.152939
R8204 VDD.n4274 VDD.n4273 0.152939
R8205 VDD.n4275 VDD.n4274 0.152939
R8206 VDD.n4276 VDD.n4275 0.152939
R8207 VDD.n4280 VDD.n4276 0.152939
R8208 VDD.n4281 VDD.n4280 0.152939
R8209 VDD.n4282 VDD.n4281 0.152939
R8210 VDD.n4283 VDD.n4282 0.152939
R8211 VDD.n4290 VDD.n4283 0.152939
R8212 VDD.n4415 VDD.n4290 0.152939
R8213 VDD.n4415 VDD.n4414 0.152939
R8214 VDD.n4414 VDD.n4413 0.152939
R8215 VDD.n4413 VDD.n4291 0.152939
R8216 VDD.n4295 VDD.n4291 0.152939
R8217 VDD.n4296 VDD.n4295 0.152939
R8218 VDD.n4297 VDD.n4296 0.152939
R8219 VDD.n4301 VDD.n4297 0.152939
R8220 VDD.n4302 VDD.n4301 0.152939
R8221 VDD.n4303 VDD.n4302 0.152939
R8222 VDD.n4304 VDD.n4303 0.152939
R8223 VDD.n4308 VDD.n4304 0.152939
R8224 VDD.n4309 VDD.n4308 0.152939
R8225 VDD.n4310 VDD.n4309 0.152939
R8226 VDD.n4311 VDD.n4310 0.152939
R8227 VDD.n4315 VDD.n4311 0.152939
R8228 VDD.n4316 VDD.n4315 0.152939
R8229 VDD.n4384 VDD.n4316 0.152939
R8230 VDD.n4384 VDD.n4383 0.152939
R8231 VDD.n3973 VDD.n3972 0.152939
R8232 VDD.n3974 VDD.n3973 0.152939
R8233 VDD.n3974 VDD.n111 0.152939
R8234 VDD.n3988 VDD.n111 0.152939
R8235 VDD.n3989 VDD.n3988 0.152939
R8236 VDD.n3990 VDD.n3989 0.152939
R8237 VDD.n3990 VDD.n100 0.152939
R8238 VDD.n4004 VDD.n100 0.152939
R8239 VDD.n4005 VDD.n4004 0.152939
R8240 VDD.n4006 VDD.n4005 0.152939
R8241 VDD.n4006 VDD.n88 0.152939
R8242 VDD.n4020 VDD.n88 0.152939
R8243 VDD.n4021 VDD.n4020 0.152939
R8244 VDD.n4022 VDD.n4021 0.152939
R8245 VDD.n4022 VDD.n76 0.152939
R8246 VDD.n4036 VDD.n76 0.152939
R8247 VDD.n4037 VDD.n4036 0.152939
R8248 VDD.n4038 VDD.n4037 0.152939
R8249 VDD.n4038 VDD.n65 0.152939
R8250 VDD.n4053 VDD.n65 0.152939
R8251 VDD.n4054 VDD.n4053 0.152939
R8252 VDD.n4055 VDD.n4054 0.152939
R8253 VDD.n4055 VDD.n53 0.152939
R8254 VDD.n4069 VDD.n53 0.152939
R8255 VDD.n4070 VDD.n4069 0.152939
R8256 VDD.n4071 VDD.n4070 0.152939
R8257 VDD.n4071 VDD.n41 0.152939
R8258 VDD.n4085 VDD.n41 0.152939
R8259 VDD.n4086 VDD.n4085 0.152939
R8260 VDD.n4087 VDD.n4086 0.152939
R8261 VDD.n4088 VDD.n4087 0.152939
R8262 VDD.n4089 VDD.n4088 0.152939
R8263 VDD.n4341 VDD.n4089 0.152939
R8264 VDD.n4342 VDD.n4341 0.152939
R8265 VDD.n4342 VDD.n4340 0.152939
R8266 VDD.n4346 VDD.n4340 0.152939
R8267 VDD.n4347 VDD.n4346 0.152939
R8268 VDD.n4348 VDD.n4347 0.152939
R8269 VDD.n4348 VDD.n4337 0.152939
R8270 VDD.n4352 VDD.n4337 0.152939
R8271 VDD.n4353 VDD.n4352 0.152939
R8272 VDD.n4354 VDD.n4353 0.152939
R8273 VDD.n4354 VDD.n4334 0.152939
R8274 VDD.n4358 VDD.n4334 0.152939
R8275 VDD.n4359 VDD.n4358 0.152939
R8276 VDD.n4360 VDD.n4359 0.152939
R8277 VDD.n4360 VDD.n4331 0.152939
R8278 VDD.n4364 VDD.n4331 0.152939
R8279 VDD.n4365 VDD.n4364 0.152939
R8280 VDD.n4366 VDD.n4365 0.152939
R8281 VDD.n4366 VDD.n4328 0.152939
R8282 VDD.n4370 VDD.n4328 0.152939
R8283 VDD.n4371 VDD.n4370 0.152939
R8284 VDD.n4372 VDD.n4371 0.152939
R8285 VDD.n4372 VDD.n4325 0.152939
R8286 VDD.n4376 VDD.n4325 0.152939
R8287 VDD.n4377 VDD.n4376 0.152939
R8288 VDD.n4378 VDD.n4377 0.152939
R8289 VDD.n4378 VDD.n4322 0.152939
R8290 VDD.n4382 VDD.n4322 0.152939
R8291 VDD.n3766 VDD.n3763 0.152939
R8292 VDD.n3767 VDD.n3766 0.152939
R8293 VDD.n3831 VDD.n3767 0.152939
R8294 VDD.n3831 VDD.n3830 0.152939
R8295 VDD.n3830 VDD.n3829 0.152939
R8296 VDD.n3829 VDD.n3769 0.152939
R8297 VDD.n3774 VDD.n3769 0.152939
R8298 VDD.n3775 VDD.n3774 0.152939
R8299 VDD.n3778 VDD.n3775 0.152939
R8300 VDD.n3779 VDD.n3778 0.152939
R8301 VDD.n3780 VDD.n3779 0.152939
R8302 VDD.n3781 VDD.n3780 0.152939
R8303 VDD.n3784 VDD.n3781 0.152939
R8304 VDD.n3785 VDD.n3784 0.152939
R8305 VDD.n3786 VDD.n3785 0.152939
R8306 VDD.n3787 VDD.n3786 0.152939
R8307 VDD.n3790 VDD.n3787 0.152939
R8308 VDD.n3791 VDD.n3790 0.152939
R8309 VDD.n3799 VDD.n3791 0.152939
R8310 VDD.n3799 VDD.n3798 0.152939
R8311 VDD.n3798 VDD.n124 0.152939
R8312 VDD.n2206 VDD.n1159 0.152939
R8313 VDD.n2202 VDD.n1159 0.152939
R8314 VDD.n2202 VDD.n2201 0.152939
R8315 VDD.n2201 VDD.n2200 0.152939
R8316 VDD.n2200 VDD.n1167 0.152939
R8317 VDD.n2196 VDD.n1167 0.152939
R8318 VDD.n2196 VDD.n2195 0.152939
R8319 VDD.n2195 VDD.n2194 0.152939
R8320 VDD.n2194 VDD.n1172 0.152939
R8321 VDD.n2190 VDD.n1172 0.152939
R8322 VDD.n2190 VDD.n2189 0.152939
R8323 VDD.n2189 VDD.n2188 0.152939
R8324 VDD.n2188 VDD.n1177 0.152939
R8325 VDD.n2184 VDD.n1177 0.152939
R8326 VDD.n2184 VDD.n2183 0.152939
R8327 VDD.n2183 VDD.n2182 0.152939
R8328 VDD.n2182 VDD.n1182 0.152939
R8329 VDD.n2178 VDD.n1182 0.152939
R8330 VDD.n2178 VDD.n2177 0.152939
R8331 VDD.n2177 VDD.n2176 0.152939
R8332 VDD.n2176 VDD.n1187 0.152939
R8333 VDD.n1700 VDD.n1699 0.152939
R8334 VDD.n1701 VDD.n1700 0.152939
R8335 VDD.n1701 VDD.n1374 0.152939
R8336 VDD.n1715 VDD.n1374 0.152939
R8337 VDD.n1716 VDD.n1715 0.152939
R8338 VDD.n1717 VDD.n1716 0.152939
R8339 VDD.n1717 VDD.n1363 0.152939
R8340 VDD.n1731 VDD.n1363 0.152939
R8341 VDD.n1732 VDD.n1731 0.152939
R8342 VDD.n1733 VDD.n1732 0.152939
R8343 VDD.n1733 VDD.n1351 0.152939
R8344 VDD.n1747 VDD.n1351 0.152939
R8345 VDD.n1748 VDD.n1747 0.152939
R8346 VDD.n1749 VDD.n1748 0.152939
R8347 VDD.n1749 VDD.n1339 0.152939
R8348 VDD.n1763 VDD.n1339 0.152939
R8349 VDD.n1764 VDD.n1763 0.152939
R8350 VDD.n1765 VDD.n1764 0.152939
R8351 VDD.n1765 VDD.n1328 0.152939
R8352 VDD.n1780 VDD.n1328 0.152939
R8353 VDD.n1781 VDD.n1780 0.152939
R8354 VDD.n1782 VDD.n1781 0.152939
R8355 VDD.n1782 VDD.n1316 0.152939
R8356 VDD.n1796 VDD.n1316 0.152939
R8357 VDD.n1797 VDD.n1796 0.152939
R8358 VDD.n1798 VDD.n1797 0.152939
R8359 VDD.n1798 VDD.n1304 0.152939
R8360 VDD.n1812 VDD.n1304 0.152939
R8361 VDD.n1813 VDD.n1812 0.152939
R8362 VDD.n1814 VDD.n1813 0.152939
R8363 VDD.n1814 VDD.n1292 0.152939
R8364 VDD.n1842 VDD.n1292 0.152939
R8365 VDD.n1843 VDD.n1842 0.152939
R8366 VDD.n1844 VDD.n1843 0.152939
R8367 VDD.n1844 VDD.n1280 0.152939
R8368 VDD.n1858 VDD.n1280 0.152939
R8369 VDD.n1859 VDD.n1858 0.152939
R8370 VDD.n1860 VDD.n1859 0.152939
R8371 VDD.n1860 VDD.n1268 0.152939
R8372 VDD.n1874 VDD.n1268 0.152939
R8373 VDD.n1875 VDD.n1874 0.152939
R8374 VDD.n1876 VDD.n1875 0.152939
R8375 VDD.n1876 VDD.n1256 0.152939
R8376 VDD.n1890 VDD.n1256 0.152939
R8377 VDD.n1891 VDD.n1890 0.152939
R8378 VDD.n1892 VDD.n1891 0.152939
R8379 VDD.n1892 VDD.n1244 0.152939
R8380 VDD.n1906 VDD.n1244 0.152939
R8381 VDD.n1907 VDD.n1906 0.152939
R8382 VDD.n1908 VDD.n1907 0.152939
R8383 VDD.n1908 VDD.n1232 0.152939
R8384 VDD.n1922 VDD.n1232 0.152939
R8385 VDD.n1923 VDD.n1922 0.152939
R8386 VDD.n1924 VDD.n1923 0.152939
R8387 VDD.n1924 VDD.n1220 0.152939
R8388 VDD.n1938 VDD.n1220 0.152939
R8389 VDD.n1939 VDD.n1938 0.152939
R8390 VDD.n1942 VDD.n1939 0.152939
R8391 VDD.n1942 VDD.n1941 0.152939
R8392 VDD.n1941 VDD.n1940 0.152939
R8393 VDD.n1692 VDD.n1391 0.152939
R8394 VDD.n1688 VDD.n1391 0.152939
R8395 VDD.n1688 VDD.n1687 0.152939
R8396 VDD.n1687 VDD.n1686 0.152939
R8397 VDD.n1686 VDD.n1396 0.152939
R8398 VDD.n1682 VDD.n1396 0.152939
R8399 VDD.n1682 VDD.n1681 0.152939
R8400 VDD.n1681 VDD.n1680 0.152939
R8401 VDD.n1680 VDD.n1404 0.152939
R8402 VDD.n1676 VDD.n1404 0.152939
R8403 VDD.n1676 VDD.n1675 0.152939
R8404 VDD.n1675 VDD.n1674 0.152939
R8405 VDD.n1674 VDD.n1412 0.152939
R8406 VDD.n1670 VDD.n1412 0.152939
R8407 VDD.n1670 VDD.n1669 0.152939
R8408 VDD.n1669 VDD.n1422 0.152939
R8409 VDD.n1665 VDD.n1422 0.152939
R8410 VDD.n1665 VDD.n1664 0.152939
R8411 VDD.n1664 VDD.n1663 0.152939
R8412 VDD.n1663 VDD.n1428 0.152939
R8413 VDD.n1659 VDD.n1428 0.152939
R8414 VDD.n1659 VDD.n1658 0.152939
R8415 VDD.n1658 VDD.n1657 0.152939
R8416 VDD.n1657 VDD.n1436 0.152939
R8417 VDD.n1653 VDD.n1436 0.152939
R8418 VDD.n1653 VDD.n1652 0.152939
R8419 VDD.n1652 VDD.n1651 0.152939
R8420 VDD.n1651 VDD.n1444 0.152939
R8421 VDD.n1647 VDD.n1444 0.152939
R8422 VDD.n1647 VDD.n1646 0.152939
R8423 VDD.n1646 VDD.n1645 0.152939
R8424 VDD.n1645 VDD.n1452 0.152939
R8425 VDD.n1638 VDD.n1452 0.152939
R8426 VDD.n1638 VDD.n1637 0.152939
R8427 VDD.n1637 VDD.n1636 0.152939
R8428 VDD.n1636 VDD.n1460 0.152939
R8429 VDD.n1632 VDD.n1460 0.152939
R8430 VDD.n1632 VDD.n1631 0.152939
R8431 VDD.n1631 VDD.n1630 0.152939
R8432 VDD.n1630 VDD.n1468 0.152939
R8433 VDD.n1626 VDD.n1468 0.152939
R8434 VDD.n1626 VDD.n1625 0.152939
R8435 VDD.n1625 VDD.n1624 0.152939
R8436 VDD.n1624 VDD.n1476 0.152939
R8437 VDD.n1620 VDD.n1476 0.152939
R8438 VDD.n1620 VDD.n1619 0.152939
R8439 VDD.n1619 VDD.n1618 0.152939
R8440 VDD.n1618 VDD.n1484 0.152939
R8441 VDD.n1492 VDD.n1484 0.152939
R8442 VDD.n1496 VDD.n1492 0.152939
R8443 VDD.n1609 VDD.n1496 0.152939
R8444 VDD.n1609 VDD.n1608 0.152939
R8445 VDD.n1608 VDD.n1607 0.152939
R8446 VDD.n1607 VDD.n1497 0.152939
R8447 VDD.n1603 VDD.n1497 0.152939
R8448 VDD.n1603 VDD.n1602 0.152939
R8449 VDD.n1602 VDD.n1601 0.152939
R8450 VDD.n1601 VDD.n1504 0.152939
R8451 VDD.n1597 VDD.n1504 0.152939
R8452 VDD.n1597 VDD.n1596 0.152939
R8453 VDD.n1596 VDD.n1595 0.152939
R8454 VDD.n1595 VDD.n1512 0.152939
R8455 VDD.n1591 VDD.n1512 0.152939
R8456 VDD.n1591 VDD.n1590 0.152939
R8457 VDD.n1590 VDD.n1589 0.152939
R8458 VDD.n1589 VDD.n1520 0.152939
R8459 VDD.n1580 VDD.n1520 0.152939
R8460 VDD.n1580 VDD.n1579 0.152939
R8461 VDD.n1579 VDD.n1578 0.152939
R8462 VDD.n1578 VDD.n1526 0.152939
R8463 VDD.n1574 VDD.n1526 0.152939
R8464 VDD.n1574 VDD.n1573 0.152939
R8465 VDD.n1573 VDD.n1572 0.152939
R8466 VDD.n1572 VDD.n1533 0.152939
R8467 VDD.n1568 VDD.n1533 0.152939
R8468 VDD.n1568 VDD.n1567 0.152939
R8469 VDD.n1567 VDD.n1566 0.152939
R8470 VDD.n1566 VDD.n1541 0.152939
R8471 VDD.n1562 VDD.n1541 0.152939
R8472 VDD.n1562 VDD.n1561 0.152939
R8473 VDD.n1561 VDD.n1560 0.152939
R8474 VDD.n1560 VDD.n1549 0.152939
R8475 VDD.n1549 VDD.n1387 0.152939
R8476 VDD.n1693 VDD.n1381 0.152939
R8477 VDD.n1707 VDD.n1381 0.152939
R8478 VDD.n1708 VDD.n1707 0.152939
R8479 VDD.n1709 VDD.n1708 0.152939
R8480 VDD.n1709 VDD.n1369 0.152939
R8481 VDD.n1723 VDD.n1369 0.152939
R8482 VDD.n1724 VDD.n1723 0.152939
R8483 VDD.n1725 VDD.n1724 0.152939
R8484 VDD.n1725 VDD.n1357 0.152939
R8485 VDD.n1739 VDD.n1357 0.152939
R8486 VDD.n1740 VDD.n1739 0.152939
R8487 VDD.n1741 VDD.n1740 0.152939
R8488 VDD.n1741 VDD.n1345 0.152939
R8489 VDD.n1755 VDD.n1345 0.152939
R8490 VDD.n1756 VDD.n1755 0.152939
R8491 VDD.n1757 VDD.n1756 0.152939
R8492 VDD.n1757 VDD.n1333 0.152939
R8493 VDD.n1772 VDD.n1333 0.152939
R8494 VDD.n1773 VDD.n1772 0.152939
R8495 VDD.n1774 VDD.n1773 0.152939
R8496 VDD.n1774 VDD.n1322 0.152939
R8497 VDD.n1788 VDD.n1322 0.152939
R8498 VDD.n1789 VDD.n1788 0.152939
R8499 VDD.n1790 VDD.n1789 0.152939
R8500 VDD.n1790 VDD.n1310 0.152939
R8501 VDD.n1804 VDD.n1310 0.152939
R8502 VDD.n1805 VDD.n1804 0.152939
R8503 VDD.n1806 VDD.n1805 0.152939
R8504 VDD.n1806 VDD.n1298 0.152939
R8505 VDD.n1835 VDD.n1834 0.145814
R8506 VDD.n4604 VDD.n30 0.145814
R8507 VDD.n4604 VDD.n31 0.145814
R8508 VDD.n1834 VDD.n1298 0.145814
R8509 VDD.n773 VDD.t135 0.106716
R8510 VDD.n2782 VDD.t125 0.106716
R8511 VDD.t149 VDD.n566 0.106716
R8512 VDD.n3473 VDD.t153 0.106716
R8513 VDD.n2121 VDD.n1988 0.0889146
R8514 VDD.n3917 VDD.n3916 0.0889146
R8515 VDD.n3763 VDD.n3762 0.0889146
R8516 VDD.n2207 VDD.n2206 0.0889146
R8517 VDD.n2121 VDD.n2120 0.0645244
R8518 VDD.n2207 VDD.n1156 0.0645244
R8519 VDD.n3917 VDD.n163 0.0645244
R8520 VDD.n3762 VDD.n220 0.0645244
R8521 VDD VDD.n15 0.00833333
R8522 CS_BIAS.n9 CS_BIAS.n8 161.3
R8523 CS_BIAS.n10 CS_BIAS.n2 161.3
R8524 CS_BIAS.n12 CS_BIAS.n11 161.3
R8525 CS_BIAS.n13 CS_BIAS.n1 161.3
R8526 CS_BIAS.n15 CS_BIAS.n14 161.3
R8527 CS_BIAS.n16 CS_BIAS.n0 161.3
R8528 CS_BIAS.n41 CS_BIAS.n25 161.3
R8529 CS_BIAS.n40 CS_BIAS.n39 161.3
R8530 CS_BIAS.n38 CS_BIAS.n26 161.3
R8531 CS_BIAS.n37 CS_BIAS.n36 161.3
R8532 CS_BIAS.n35 CS_BIAS.n27 161.3
R8533 CS_BIAS.n34 CS_BIAS.n33 161.3
R8534 CS_BIAS.n9 CS_BIAS.n3 122.968
R8535 CS_BIAS.n34 CS_BIAS.n28 122.968
R8536 CS_BIAS.n6 CS_BIAS.n5 78.7033
R8537 CS_BIAS.n31 CS_BIAS.n29 78.7033
R8538 CS_BIAS.n18 CS_BIAS.n17 54.5572
R8539 CS_BIAS.n43 CS_BIAS.n42 54.5572
R8540 CS_BIAS.n23 CS_BIAS.t16 45.9483
R8541 CS_BIAS.n48 CS_BIAS.t23 45.9483
R8542 CS_BIAS.n46 CS_BIAS.t14 45.9483
R8543 CS_BIAS.n44 CS_BIAS.t8 45.9483
R8544 CS_BIAS.n30 CS_BIAS.t2 45.9483
R8545 CS_BIAS.n21 CS_BIAS.t21 45.9479
R8546 CS_BIAS.n19 CS_BIAS.t18 45.9479
R8547 CS_BIAS.n4 CS_BIAS.t0 45.9479
R8548 CS_BIAS.n23 CS_BIAS.t19 43.5984
R8549 CS_BIAS.n21 CS_BIAS.t22 43.5984
R8550 CS_BIAS.n19 CS_BIAS.t20 43.5984
R8551 CS_BIAS.n4 CS_BIAS.t4 43.5984
R8552 CS_BIAS.n48 CS_BIAS.t9 43.5984
R8553 CS_BIAS.n46 CS_BIAS.t17 43.5984
R8554 CS_BIAS.n44 CS_BIAS.t11 43.5984
R8555 CS_BIAS.n30 CS_BIAS.t6 43.5984
R8556 CS_BIAS.n28 CS_BIAS.t15 39.5493
R8557 CS_BIAS.n3 CS_BIAS.t12 39.549
R8558 CS_BIAS.n10 CS_BIAS.n9 32.2376
R8559 CS_BIAS.n35 CS_BIAS.n34 32.2376
R8560 CS_BIAS.n16 CS_BIAS.n15 24.4675
R8561 CS_BIAS.n15 CS_BIAS.n1 24.4675
R8562 CS_BIAS.n11 CS_BIAS.n1 24.4675
R8563 CS_BIAS.n11 CS_BIAS.n10 24.4675
R8564 CS_BIAS.n36 CS_BIAS.n35 24.4675
R8565 CS_BIAS.n36 CS_BIAS.n26 24.4675
R8566 CS_BIAS.n40 CS_BIAS.n26 24.4675
R8567 CS_BIAS.n41 CS_BIAS.n40 24.4675
R8568 CS_BIAS.n17 CS_BIAS.n16 22.7548
R8569 CS_BIAS.n42 CS_BIAS.n41 22.7548
R8570 CS_BIAS.n31 CS_BIAS.n30 13.3368
R8571 CS_BIAS.n6 CS_BIAS.n4 13.3368
R8572 CS_BIAS.n5 CS_BIAS.t5 13.3338
R8573 CS_BIAS.n5 CS_BIAS.t1 13.3338
R8574 CS_BIAS.n29 CS_BIAS.t3 13.3338
R8575 CS_BIAS.n29 CS_BIAS.t7 13.3338
R8576 CS_BIAS.n17 CS_BIAS.t10 12.4055
R8577 CS_BIAS.n42 CS_BIAS.t13 12.4055
R8578 CS_BIAS.n7 CS_BIAS.n6 9.50363
R8579 CS_BIAS.n32 CS_BIAS.n31 9.50363
R8580 CS_BIAS.n50 CS_BIAS.n24 8.62412
R8581 CS_BIAS.n20 CS_BIAS.n18 7.94595
R8582 CS_BIAS.n45 CS_BIAS.n43 7.94595
R8583 CS_BIAS.n50 CS_BIAS.n49 6.52792
R8584 CS_BIAS.n24 CS_BIAS.n23 6.06568
R8585 CS_BIAS.n49 CS_BIAS.n48 6.06568
R8586 CS_BIAS.n47 CS_BIAS.n46 6.06568
R8587 CS_BIAS.n45 CS_BIAS.n44 6.06568
R8588 CS_BIAS.n22 CS_BIAS.n21 6.06567
R8589 CS_BIAS.n20 CS_BIAS.n19 6.06567
R8590 CS_BIAS.n32 CS_BIAS.n28 5.54113
R8591 CS_BIAS.n7 CS_BIAS.n3 5.54106
R8592 CS_BIAS CS_BIAS.n50 5.07654
R8593 CS_BIAS.n22 CS_BIAS.n20 2.38686
R8594 CS_BIAS.n24 CS_BIAS.n22 2.38686
R8595 CS_BIAS.n47 CS_BIAS.n45 2.38686
R8596 CS_BIAS.n49 CS_BIAS.n47 2.38686
R8597 CS_BIAS.n18 CS_BIAS.n0 0.502622
R8598 CS_BIAS.n43 CS_BIAS.n25 0.502622
R8599 CS_BIAS.n14 CS_BIAS.n0 0.189894
R8600 CS_BIAS.n14 CS_BIAS.n13 0.189894
R8601 CS_BIAS.n13 CS_BIAS.n12 0.189894
R8602 CS_BIAS.n12 CS_BIAS.n2 0.189894
R8603 CS_BIAS.n8 CS_BIAS.n2 0.189894
R8604 CS_BIAS.n33 CS_BIAS.n27 0.189894
R8605 CS_BIAS.n37 CS_BIAS.n27 0.189894
R8606 CS_BIAS.n38 CS_BIAS.n37 0.189894
R8607 CS_BIAS.n39 CS_BIAS.n38 0.189894
R8608 CS_BIAS.n39 CS_BIAS.n25 0.189894
R8609 CS_BIAS.n8 CS_BIAS.n7 0.0762576
R8610 CS_BIAS.n33 CS_BIAS.n32 0.0762576
R8611 VOUT.n29 VOUT.t30 111.986
R8612 VOUT.n26 VOUT.t33 111.986
R8613 VOUT.n23 VOUT.t26 111.986
R8614 VOUT.n20 VOUT.t18 111.986
R8615 VOUT.n18 VOUT.t32 111.986
R8616 VOUT.n12 VOUT.t34 110.448
R8617 VOUT.n9 VOUT.t35 110.448
R8618 VOUT.n6 VOUT.t25 110.448
R8619 VOUT.n3 VOUT.t27 110.448
R8620 VOUT.n1 VOUT.t22 110.448
R8621 VOUT.n12 VOUT.n11 99.1374
R8622 VOUT.n9 VOUT.n8 99.1374
R8623 VOUT.n6 VOUT.n5 99.1374
R8624 VOUT.n3 VOUT.n2 99.1374
R8625 VOUT.n1 VOUT.n0 99.1374
R8626 VOUT.n26 VOUT.n25 97.6001
R8627 VOUT.n23 VOUT.n22 97.6001
R8628 VOUT.n20 VOUT.n19 97.6001
R8629 VOUT.n18 VOUT.n17 97.6001
R8630 VOUT.n29 VOUT.n28 97.5999
R8631 VOUT.n34 VOUT.n32 85.3571
R8632 VOUT.n42 VOUT.n40 85.3571
R8633 VOUT.n38 VOUT.n37 84.4375
R8634 VOUT.n36 VOUT.n35 84.4375
R8635 VOUT.n34 VOUT.n33 84.4375
R8636 VOUT.n46 VOUT.n45 84.4375
R8637 VOUT.n44 VOUT.n43 84.4375
R8638 VOUT.n42 VOUT.n41 84.4375
R8639 VOUT.n37 VOUT.t4 13.3338
R8640 VOUT.n37 VOUT.t2 13.3338
R8641 VOUT.n35 VOUT.t17 13.3338
R8642 VOUT.n35 VOUT.t12 13.3338
R8643 VOUT.n33 VOUT.t11 13.3338
R8644 VOUT.n33 VOUT.t16 13.3338
R8645 VOUT.n32 VOUT.t5 13.3338
R8646 VOUT.n32 VOUT.t8 13.3338
R8647 VOUT.n45 VOUT.t9 13.3338
R8648 VOUT.n45 VOUT.t6 13.3338
R8649 VOUT.n43 VOUT.t14 13.3338
R8650 VOUT.n43 VOUT.t10 13.3338
R8651 VOUT.n41 VOUT.t7 13.3338
R8652 VOUT.n41 VOUT.t3 13.3338
R8653 VOUT.n40 VOUT.t15 13.3338
R8654 VOUT.n40 VOUT.t13 13.3338
R8655 VOUT.n28 VOUT.t40 12.8483
R8656 VOUT.n28 VOUT.t39 12.8483
R8657 VOUT.n25 VOUT.t19 12.8483
R8658 VOUT.n25 VOUT.t29 12.8483
R8659 VOUT.n22 VOUT.t38 12.8483
R8660 VOUT.n22 VOUT.t45 12.8483
R8661 VOUT.n19 VOUT.t23 12.8483
R8662 VOUT.n19 VOUT.t24 12.8483
R8663 VOUT.n17 VOUT.t44 12.8483
R8664 VOUT.n17 VOUT.t21 12.8483
R8665 VOUT.n11 VOUT.t41 12.8483
R8666 VOUT.n11 VOUT.t28 12.8483
R8667 VOUT.n8 VOUT.t37 12.8483
R8668 VOUT.n8 VOUT.t42 12.8483
R8669 VOUT.n5 VOUT.t0 12.8483
R8670 VOUT.n5 VOUT.t20 12.8483
R8671 VOUT.n2 VOUT.t36 12.8483
R8672 VOUT.n2 VOUT.t1 12.8483
R8673 VOUT.n0 VOUT.t43 12.8483
R8674 VOUT.n0 VOUT.t31 12.8483
R8675 VOUT.n39 VOUT.n31 10.2716
R8676 VOUT.n21 VOUT.n18 6.79863
R8677 VOUT.n4 VOUT.n1 6.02995
R8678 VOUT.n31 VOUT.n14 5.76051
R8679 VOUT.n30 VOUT.n29 5.57952
R8680 VOUT.n27 VOUT.n26 5.57952
R8681 VOUT.n24 VOUT.n23 5.57952
R8682 VOUT.n21 VOUT.n20 5.57952
R8683 VOUT.n48 VOUT.n14 5.15741
R8684 VOUT.n48 VOUT.n47 5.09514
R8685 VOUT.n13 VOUT.n12 4.81084
R8686 VOUT.n10 VOUT.n9 4.81084
R8687 VOUT.n7 VOUT.n6 4.81084
R8688 VOUT.n4 VOUT.n3 4.81084
R8689 VOUT.n31 VOUT.n30 4.39254
R8690 VOUT.n14 VOUT.n13 4.39254
R8691 VOUT.n39 VOUT.n38 4.24958
R8692 VOUT.n47 VOUT.n46 4.24958
R8693 VOUT.n16 VOUT 3.10955
R8694 VOUT.n47 VOUT.n39 3.01195
R8695 VOUT.n30 VOUT.n27 1.21961
R8696 VOUT.n27 VOUT.n24 1.21961
R8697 VOUT.n24 VOUT.n21 1.21961
R8698 VOUT.n13 VOUT.n10 1.21961
R8699 VOUT.n10 VOUT.n7 1.21961
R8700 VOUT.n7 VOUT.n4 1.21961
R8701 VOUT.n38 VOUT.n36 0.92004
R8702 VOUT.n36 VOUT.n34 0.92004
R8703 VOUT.n46 VOUT.n44 0.92004
R8704 VOUT.n44 VOUT.n42 0.92004
R8705 VOUT.n16 VOUT.n15 0.376486
R8706 VOUT.n48 VOUT.n16 0.302005
R8707 VOUT.n15 VOUT.t46 0.106373
R8708 VOUT.n15 VOUT.t47 0.0345405
R8709 VOUT VOUT.n48 0.0099
R8710 GND.n7339 GND.n679 2269.2
R8711 GND.n6174 GND.n6173 1148.21
R8712 GND.n6357 GND.n1267 766.379
R8713 GND.n7338 GND.n680 766.379
R8714 GND.n7564 GND.n546 766.379
R8715 GND.n6175 GND.n1445 766.379
R8716 GND.n5124 GND.n176 754.366
R8717 GND.n5152 GND.n181 754.366
R8718 GND.n4910 GND.n4801 754.366
R8719 GND.n2902 GND.n2598 754.366
R8720 GND.n6003 GND.n1648 754.366
R8721 GND.n1668 GND.n1646 754.366
R8722 GND.n4222 GND.n4221 754.366
R8723 GND.n5891 GND.n1748 754.366
R8724 GND.n6358 GND.n1266 744.005
R8725 GND.n5522 GND.n2372 703.915
R8726 GND.n5479 GND.n5478 703.915
R8727 GND.n4257 GND.n3079 703.915
R8728 GND.n4255 GND.n3081 703.915
R8729 GND.n378 GND.n171 699.111
R8730 GND.n7739 GND.n180 699.111
R8731 GND.n4908 GND.n4907 699.111
R8732 GND.n5402 GND.n2590 699.111
R8733 GND.n5888 GND.n1782 699.111
R8734 GND.n4224 GND.n3185 699.111
R8735 GND.n3667 GND.n1640 699.111
R8736 GND.n3670 GND.n3483 699.111
R8737 GND.n6353 GND.n1267 585
R8738 GND.n1267 GND.n1266 585
R8739 GND.n6352 GND.n6351 585
R8740 GND.n6351 GND.n6350 585
R8741 GND.n1270 GND.n1269 585
R8742 GND.n6349 GND.n1270 585
R8743 GND.n6347 GND.n6346 585
R8744 GND.n6348 GND.n6347 585
R8745 GND.n6345 GND.n1272 585
R8746 GND.n1272 GND.n1271 585
R8747 GND.n6344 GND.n6343 585
R8748 GND.n6343 GND.n6342 585
R8749 GND.n1278 GND.n1277 585
R8750 GND.n6341 GND.n1278 585
R8751 GND.n6339 GND.n6338 585
R8752 GND.n6340 GND.n6339 585
R8753 GND.n6337 GND.n1280 585
R8754 GND.n1280 GND.n1279 585
R8755 GND.n6336 GND.n6335 585
R8756 GND.n6335 GND.n6334 585
R8757 GND.n1286 GND.n1285 585
R8758 GND.n6333 GND.n1286 585
R8759 GND.n6331 GND.n6330 585
R8760 GND.n6332 GND.n6331 585
R8761 GND.n6329 GND.n1288 585
R8762 GND.n1288 GND.n1287 585
R8763 GND.n6328 GND.n6327 585
R8764 GND.n6327 GND.n6326 585
R8765 GND.n1294 GND.n1293 585
R8766 GND.n6325 GND.n1294 585
R8767 GND.n6323 GND.n6322 585
R8768 GND.n6324 GND.n6323 585
R8769 GND.n6321 GND.n1296 585
R8770 GND.n1296 GND.n1295 585
R8771 GND.n6320 GND.n6319 585
R8772 GND.n6319 GND.n6318 585
R8773 GND.n1302 GND.n1301 585
R8774 GND.n6317 GND.n1302 585
R8775 GND.n6315 GND.n6314 585
R8776 GND.n6316 GND.n6315 585
R8777 GND.n6313 GND.n1304 585
R8778 GND.n1304 GND.n1303 585
R8779 GND.n6312 GND.n6311 585
R8780 GND.n6311 GND.n6310 585
R8781 GND.n1310 GND.n1309 585
R8782 GND.n6309 GND.n1310 585
R8783 GND.n6307 GND.n6306 585
R8784 GND.n6308 GND.n6307 585
R8785 GND.n6305 GND.n1312 585
R8786 GND.n1312 GND.n1311 585
R8787 GND.n6304 GND.n6303 585
R8788 GND.n6303 GND.n6302 585
R8789 GND.n1318 GND.n1317 585
R8790 GND.n6301 GND.n1318 585
R8791 GND.n6299 GND.n6298 585
R8792 GND.n6300 GND.n6299 585
R8793 GND.n6297 GND.n1320 585
R8794 GND.n1320 GND.n1319 585
R8795 GND.n6296 GND.n6295 585
R8796 GND.n6295 GND.n6294 585
R8797 GND.n1326 GND.n1325 585
R8798 GND.n6293 GND.n1326 585
R8799 GND.n6291 GND.n6290 585
R8800 GND.n6292 GND.n6291 585
R8801 GND.n6289 GND.n1328 585
R8802 GND.n1328 GND.n1327 585
R8803 GND.n6288 GND.n6287 585
R8804 GND.n6287 GND.n6286 585
R8805 GND.n1334 GND.n1333 585
R8806 GND.n6285 GND.n1334 585
R8807 GND.n6283 GND.n6282 585
R8808 GND.n6284 GND.n6283 585
R8809 GND.n6281 GND.n1336 585
R8810 GND.n1336 GND.n1335 585
R8811 GND.n6280 GND.n6279 585
R8812 GND.n6279 GND.n6278 585
R8813 GND.n1342 GND.n1341 585
R8814 GND.n6277 GND.n1342 585
R8815 GND.n6275 GND.n6274 585
R8816 GND.n6276 GND.n6275 585
R8817 GND.n6273 GND.n1344 585
R8818 GND.n1344 GND.n1343 585
R8819 GND.n6272 GND.n6271 585
R8820 GND.n6271 GND.n6270 585
R8821 GND.n1350 GND.n1349 585
R8822 GND.n6269 GND.n1350 585
R8823 GND.n6267 GND.n6266 585
R8824 GND.n6268 GND.n6267 585
R8825 GND.n6265 GND.n1352 585
R8826 GND.n1352 GND.n1351 585
R8827 GND.n6264 GND.n6263 585
R8828 GND.n6263 GND.n6262 585
R8829 GND.n1358 GND.n1357 585
R8830 GND.n6261 GND.n1358 585
R8831 GND.n6259 GND.n6258 585
R8832 GND.n6260 GND.n6259 585
R8833 GND.n6257 GND.n1360 585
R8834 GND.n1360 GND.n1359 585
R8835 GND.n6256 GND.n6255 585
R8836 GND.n6255 GND.n6254 585
R8837 GND.n1366 GND.n1365 585
R8838 GND.n6253 GND.n1366 585
R8839 GND.n6251 GND.n6250 585
R8840 GND.n6252 GND.n6251 585
R8841 GND.n6249 GND.n1368 585
R8842 GND.n1368 GND.n1367 585
R8843 GND.n6248 GND.n6247 585
R8844 GND.n6247 GND.n6246 585
R8845 GND.n1374 GND.n1373 585
R8846 GND.n6245 GND.n1374 585
R8847 GND.n6243 GND.n6242 585
R8848 GND.n6244 GND.n6243 585
R8849 GND.n6241 GND.n1376 585
R8850 GND.n1376 GND.n1375 585
R8851 GND.n6240 GND.n6239 585
R8852 GND.n6239 GND.n6238 585
R8853 GND.n1382 GND.n1381 585
R8854 GND.n6237 GND.n1382 585
R8855 GND.n6235 GND.n6234 585
R8856 GND.n6236 GND.n6235 585
R8857 GND.n6233 GND.n1384 585
R8858 GND.n1384 GND.n1383 585
R8859 GND.n6232 GND.n6231 585
R8860 GND.n6231 GND.n6230 585
R8861 GND.n1390 GND.n1389 585
R8862 GND.n6229 GND.n1390 585
R8863 GND.n6227 GND.n6226 585
R8864 GND.n6228 GND.n6227 585
R8865 GND.n6225 GND.n1392 585
R8866 GND.n1392 GND.n1391 585
R8867 GND.n6224 GND.n6223 585
R8868 GND.n6223 GND.n6222 585
R8869 GND.n1398 GND.n1397 585
R8870 GND.n6221 GND.n1398 585
R8871 GND.n6219 GND.n6218 585
R8872 GND.n6220 GND.n6219 585
R8873 GND.n6217 GND.n1400 585
R8874 GND.n1400 GND.n1399 585
R8875 GND.n6216 GND.n6215 585
R8876 GND.n6215 GND.n6214 585
R8877 GND.n1406 GND.n1405 585
R8878 GND.n6213 GND.n1406 585
R8879 GND.n6211 GND.n6210 585
R8880 GND.n6212 GND.n6211 585
R8881 GND.n6209 GND.n1408 585
R8882 GND.n1408 GND.n1407 585
R8883 GND.n6208 GND.n6207 585
R8884 GND.n6207 GND.n6206 585
R8885 GND.n1414 GND.n1413 585
R8886 GND.n6205 GND.n1414 585
R8887 GND.n6203 GND.n6202 585
R8888 GND.n6204 GND.n6203 585
R8889 GND.n6201 GND.n1416 585
R8890 GND.n1416 GND.n1415 585
R8891 GND.n6200 GND.n6199 585
R8892 GND.n6199 GND.n6198 585
R8893 GND.n1422 GND.n1421 585
R8894 GND.n6197 GND.n1422 585
R8895 GND.n6195 GND.n6194 585
R8896 GND.n6196 GND.n6195 585
R8897 GND.n6193 GND.n1424 585
R8898 GND.n1424 GND.n1423 585
R8899 GND.n6192 GND.n6191 585
R8900 GND.n6191 GND.n6190 585
R8901 GND.n1430 GND.n1429 585
R8902 GND.n6189 GND.n1430 585
R8903 GND.n6187 GND.n6186 585
R8904 GND.n6188 GND.n6187 585
R8905 GND.n6185 GND.n1432 585
R8906 GND.n1432 GND.n1431 585
R8907 GND.n6184 GND.n6183 585
R8908 GND.n6183 GND.n6182 585
R8909 GND.n1438 GND.n1437 585
R8910 GND.n6181 GND.n1438 585
R8911 GND.n6179 GND.n6178 585
R8912 GND.n6180 GND.n6179 585
R8913 GND.n6177 GND.n1440 585
R8914 GND.n1440 GND.n1439 585
R8915 GND.n6176 GND.n6175 585
R8916 GND.n6175 GND.n6174 585
R8917 GND.n6357 GND.n6356 585
R8918 GND.n6358 GND.n6357 585
R8919 GND.n1265 GND.n1264 585
R8920 GND.n6359 GND.n1265 585
R8921 GND.n6362 GND.n6361 585
R8922 GND.n6361 GND.n6360 585
R8923 GND.n1262 GND.n1261 585
R8924 GND.n1261 GND.n1260 585
R8925 GND.n6367 GND.n6366 585
R8926 GND.n6368 GND.n6367 585
R8927 GND.n1259 GND.n1258 585
R8928 GND.n6369 GND.n1259 585
R8929 GND.n6372 GND.n6371 585
R8930 GND.n6371 GND.n6370 585
R8931 GND.n1256 GND.n1255 585
R8932 GND.n1255 GND.n1254 585
R8933 GND.n6377 GND.n6376 585
R8934 GND.n6378 GND.n6377 585
R8935 GND.n1253 GND.n1252 585
R8936 GND.n6379 GND.n1253 585
R8937 GND.n6382 GND.n6381 585
R8938 GND.n6381 GND.n6380 585
R8939 GND.n1250 GND.n1249 585
R8940 GND.n1249 GND.n1248 585
R8941 GND.n6387 GND.n6386 585
R8942 GND.n6388 GND.n6387 585
R8943 GND.n1247 GND.n1246 585
R8944 GND.n6389 GND.n1247 585
R8945 GND.n6392 GND.n6391 585
R8946 GND.n6391 GND.n6390 585
R8947 GND.n1244 GND.n1243 585
R8948 GND.n1243 GND.n1242 585
R8949 GND.n6397 GND.n6396 585
R8950 GND.n6398 GND.n6397 585
R8951 GND.n1241 GND.n1240 585
R8952 GND.n6399 GND.n1241 585
R8953 GND.n6402 GND.n6401 585
R8954 GND.n6401 GND.n6400 585
R8955 GND.n1238 GND.n1237 585
R8956 GND.n1237 GND.n1236 585
R8957 GND.n6407 GND.n6406 585
R8958 GND.n6408 GND.n6407 585
R8959 GND.n1235 GND.n1234 585
R8960 GND.n6409 GND.n1235 585
R8961 GND.n6412 GND.n6411 585
R8962 GND.n6411 GND.n6410 585
R8963 GND.n1232 GND.n1231 585
R8964 GND.n1231 GND.n1230 585
R8965 GND.n6417 GND.n6416 585
R8966 GND.n6418 GND.n6417 585
R8967 GND.n1229 GND.n1228 585
R8968 GND.n6419 GND.n1229 585
R8969 GND.n6422 GND.n6421 585
R8970 GND.n6421 GND.n6420 585
R8971 GND.n1226 GND.n1225 585
R8972 GND.n1225 GND.n1224 585
R8973 GND.n6427 GND.n6426 585
R8974 GND.n6428 GND.n6427 585
R8975 GND.n1223 GND.n1222 585
R8976 GND.n6429 GND.n1223 585
R8977 GND.n6432 GND.n6431 585
R8978 GND.n6431 GND.n6430 585
R8979 GND.n1220 GND.n1219 585
R8980 GND.n1219 GND.n1218 585
R8981 GND.n6437 GND.n6436 585
R8982 GND.n6438 GND.n6437 585
R8983 GND.n1217 GND.n1216 585
R8984 GND.n6439 GND.n1217 585
R8985 GND.n6442 GND.n6441 585
R8986 GND.n6441 GND.n6440 585
R8987 GND.n1214 GND.n1213 585
R8988 GND.n1213 GND.n1212 585
R8989 GND.n6447 GND.n6446 585
R8990 GND.n6448 GND.n6447 585
R8991 GND.n1211 GND.n1210 585
R8992 GND.n6449 GND.n1211 585
R8993 GND.n6452 GND.n6451 585
R8994 GND.n6451 GND.n6450 585
R8995 GND.n1208 GND.n1207 585
R8996 GND.n1207 GND.n1206 585
R8997 GND.n6457 GND.n6456 585
R8998 GND.n6458 GND.n6457 585
R8999 GND.n1205 GND.n1204 585
R9000 GND.n6459 GND.n1205 585
R9001 GND.n6462 GND.n6461 585
R9002 GND.n6461 GND.n6460 585
R9003 GND.n1202 GND.n1201 585
R9004 GND.n1201 GND.n1200 585
R9005 GND.n6467 GND.n6466 585
R9006 GND.n6468 GND.n6467 585
R9007 GND.n1199 GND.n1198 585
R9008 GND.n6469 GND.n1199 585
R9009 GND.n6472 GND.n6471 585
R9010 GND.n6471 GND.n6470 585
R9011 GND.n1196 GND.n1195 585
R9012 GND.n1195 GND.n1194 585
R9013 GND.n6477 GND.n6476 585
R9014 GND.n6478 GND.n6477 585
R9015 GND.n1193 GND.n1192 585
R9016 GND.n6479 GND.n1193 585
R9017 GND.n6482 GND.n6481 585
R9018 GND.n6481 GND.n6480 585
R9019 GND.n1190 GND.n1189 585
R9020 GND.n1189 GND.n1188 585
R9021 GND.n6487 GND.n6486 585
R9022 GND.n6488 GND.n6487 585
R9023 GND.n1187 GND.n1186 585
R9024 GND.n6489 GND.n1187 585
R9025 GND.n6492 GND.n6491 585
R9026 GND.n6491 GND.n6490 585
R9027 GND.n1184 GND.n1183 585
R9028 GND.n1183 GND.n1182 585
R9029 GND.n6497 GND.n6496 585
R9030 GND.n6498 GND.n6497 585
R9031 GND.n1181 GND.n1180 585
R9032 GND.n6499 GND.n1181 585
R9033 GND.n6502 GND.n6501 585
R9034 GND.n6501 GND.n6500 585
R9035 GND.n1178 GND.n1177 585
R9036 GND.n1177 GND.n1176 585
R9037 GND.n6507 GND.n6506 585
R9038 GND.n6508 GND.n6507 585
R9039 GND.n1175 GND.n1174 585
R9040 GND.n6509 GND.n1175 585
R9041 GND.n6512 GND.n6511 585
R9042 GND.n6511 GND.n6510 585
R9043 GND.n1172 GND.n1171 585
R9044 GND.n1171 GND.n1170 585
R9045 GND.n6517 GND.n6516 585
R9046 GND.n6518 GND.n6517 585
R9047 GND.n1169 GND.n1168 585
R9048 GND.n6519 GND.n1169 585
R9049 GND.n6522 GND.n6521 585
R9050 GND.n6521 GND.n6520 585
R9051 GND.n1166 GND.n1165 585
R9052 GND.n1165 GND.n1164 585
R9053 GND.n6527 GND.n6526 585
R9054 GND.n6528 GND.n6527 585
R9055 GND.n1163 GND.n1162 585
R9056 GND.n6529 GND.n1163 585
R9057 GND.n6532 GND.n6531 585
R9058 GND.n6531 GND.n6530 585
R9059 GND.n1160 GND.n1159 585
R9060 GND.n1159 GND.n1158 585
R9061 GND.n6537 GND.n6536 585
R9062 GND.n6538 GND.n6537 585
R9063 GND.n1157 GND.n1156 585
R9064 GND.n6539 GND.n1157 585
R9065 GND.n6542 GND.n6541 585
R9066 GND.n6541 GND.n6540 585
R9067 GND.n1154 GND.n1153 585
R9068 GND.n1153 GND.n1152 585
R9069 GND.n6547 GND.n6546 585
R9070 GND.n6548 GND.n6547 585
R9071 GND.n1151 GND.n1150 585
R9072 GND.n6549 GND.n1151 585
R9073 GND.n6552 GND.n6551 585
R9074 GND.n6551 GND.n6550 585
R9075 GND.n1148 GND.n1147 585
R9076 GND.n1147 GND.n1146 585
R9077 GND.n6557 GND.n6556 585
R9078 GND.n6558 GND.n6557 585
R9079 GND.n1145 GND.n1144 585
R9080 GND.n6559 GND.n1145 585
R9081 GND.n6562 GND.n6561 585
R9082 GND.n6561 GND.n6560 585
R9083 GND.n1142 GND.n1141 585
R9084 GND.n1141 GND.n1140 585
R9085 GND.n6567 GND.n6566 585
R9086 GND.n6568 GND.n6567 585
R9087 GND.n1139 GND.n1138 585
R9088 GND.n6569 GND.n1139 585
R9089 GND.n6572 GND.n6571 585
R9090 GND.n6571 GND.n6570 585
R9091 GND.n1136 GND.n1135 585
R9092 GND.n1135 GND.n1134 585
R9093 GND.n6577 GND.n6576 585
R9094 GND.n6578 GND.n6577 585
R9095 GND.n1133 GND.n1132 585
R9096 GND.n6579 GND.n1133 585
R9097 GND.n6582 GND.n6581 585
R9098 GND.n6581 GND.n6580 585
R9099 GND.n1130 GND.n1129 585
R9100 GND.n1129 GND.n1128 585
R9101 GND.n6587 GND.n6586 585
R9102 GND.n6588 GND.n6587 585
R9103 GND.n1127 GND.n1126 585
R9104 GND.n6589 GND.n1127 585
R9105 GND.n6592 GND.n6591 585
R9106 GND.n6591 GND.n6590 585
R9107 GND.n1124 GND.n1123 585
R9108 GND.n1123 GND.n1122 585
R9109 GND.n6597 GND.n6596 585
R9110 GND.n6598 GND.n6597 585
R9111 GND.n1121 GND.n1120 585
R9112 GND.n6599 GND.n1121 585
R9113 GND.n6602 GND.n6601 585
R9114 GND.n6601 GND.n6600 585
R9115 GND.n1118 GND.n1117 585
R9116 GND.n1117 GND.n1116 585
R9117 GND.n6607 GND.n6606 585
R9118 GND.n6608 GND.n6607 585
R9119 GND.n1115 GND.n1114 585
R9120 GND.n6609 GND.n1115 585
R9121 GND.n6612 GND.n6611 585
R9122 GND.n6611 GND.n6610 585
R9123 GND.n1112 GND.n1111 585
R9124 GND.n1111 GND.n1110 585
R9125 GND.n6617 GND.n6616 585
R9126 GND.n6618 GND.n6617 585
R9127 GND.n1109 GND.n1108 585
R9128 GND.n6619 GND.n1109 585
R9129 GND.n6622 GND.n6621 585
R9130 GND.n6621 GND.n6620 585
R9131 GND.n1106 GND.n1105 585
R9132 GND.n1105 GND.n1104 585
R9133 GND.n6627 GND.n6626 585
R9134 GND.n6628 GND.n6627 585
R9135 GND.n1103 GND.n1102 585
R9136 GND.n6629 GND.n1103 585
R9137 GND.n6632 GND.n6631 585
R9138 GND.n6631 GND.n6630 585
R9139 GND.n1100 GND.n1099 585
R9140 GND.n1099 GND.n1098 585
R9141 GND.n6637 GND.n6636 585
R9142 GND.n6638 GND.n6637 585
R9143 GND.n1097 GND.n1096 585
R9144 GND.n6639 GND.n1097 585
R9145 GND.n6642 GND.n6641 585
R9146 GND.n6641 GND.n6640 585
R9147 GND.n1094 GND.n1093 585
R9148 GND.n1093 GND.n1092 585
R9149 GND.n6647 GND.n6646 585
R9150 GND.n6648 GND.n6647 585
R9151 GND.n1091 GND.n1090 585
R9152 GND.n6649 GND.n1091 585
R9153 GND.n6652 GND.n6651 585
R9154 GND.n6651 GND.n6650 585
R9155 GND.n1088 GND.n1087 585
R9156 GND.n1087 GND.n1086 585
R9157 GND.n6657 GND.n6656 585
R9158 GND.n6658 GND.n6657 585
R9159 GND.n1085 GND.n1084 585
R9160 GND.n6659 GND.n1085 585
R9161 GND.n6662 GND.n6661 585
R9162 GND.n6661 GND.n6660 585
R9163 GND.n1082 GND.n1081 585
R9164 GND.n1081 GND.n1080 585
R9165 GND.n6667 GND.n6666 585
R9166 GND.n6668 GND.n6667 585
R9167 GND.n1079 GND.n1078 585
R9168 GND.n6669 GND.n1079 585
R9169 GND.n6672 GND.n6671 585
R9170 GND.n6671 GND.n6670 585
R9171 GND.n1076 GND.n1075 585
R9172 GND.n1075 GND.n1074 585
R9173 GND.n6677 GND.n6676 585
R9174 GND.n6678 GND.n6677 585
R9175 GND.n1073 GND.n1072 585
R9176 GND.n6679 GND.n1073 585
R9177 GND.n6682 GND.n6681 585
R9178 GND.n6681 GND.n6680 585
R9179 GND.n1070 GND.n1069 585
R9180 GND.n1069 GND.n1068 585
R9181 GND.n6687 GND.n6686 585
R9182 GND.n6688 GND.n6687 585
R9183 GND.n1067 GND.n1066 585
R9184 GND.n6689 GND.n1067 585
R9185 GND.n6692 GND.n6691 585
R9186 GND.n6691 GND.n6690 585
R9187 GND.n1064 GND.n1063 585
R9188 GND.n1063 GND.n1062 585
R9189 GND.n6697 GND.n6696 585
R9190 GND.n6698 GND.n6697 585
R9191 GND.n1061 GND.n1060 585
R9192 GND.n6699 GND.n1061 585
R9193 GND.n6702 GND.n6701 585
R9194 GND.n6701 GND.n6700 585
R9195 GND.n1058 GND.n1057 585
R9196 GND.n1057 GND.n1056 585
R9197 GND.n6707 GND.n6706 585
R9198 GND.n6708 GND.n6707 585
R9199 GND.n1055 GND.n1054 585
R9200 GND.n6709 GND.n1055 585
R9201 GND.n6712 GND.n6711 585
R9202 GND.n6711 GND.n6710 585
R9203 GND.n1052 GND.n1051 585
R9204 GND.n1051 GND.n1050 585
R9205 GND.n6717 GND.n6716 585
R9206 GND.n6718 GND.n6717 585
R9207 GND.n1049 GND.n1048 585
R9208 GND.n6719 GND.n1049 585
R9209 GND.n6722 GND.n6721 585
R9210 GND.n6721 GND.n6720 585
R9211 GND.n1046 GND.n1045 585
R9212 GND.n1045 GND.n1044 585
R9213 GND.n6727 GND.n6726 585
R9214 GND.n6728 GND.n6727 585
R9215 GND.n1043 GND.n1042 585
R9216 GND.n6729 GND.n1043 585
R9217 GND.n6732 GND.n6731 585
R9218 GND.n6731 GND.n6730 585
R9219 GND.n1040 GND.n1039 585
R9220 GND.n1039 GND.n1038 585
R9221 GND.n6737 GND.n6736 585
R9222 GND.n6738 GND.n6737 585
R9223 GND.n1037 GND.n1036 585
R9224 GND.n6739 GND.n1037 585
R9225 GND.n6742 GND.n6741 585
R9226 GND.n6741 GND.n6740 585
R9227 GND.n1034 GND.n1033 585
R9228 GND.n1033 GND.n1032 585
R9229 GND.n6747 GND.n6746 585
R9230 GND.n6748 GND.n6747 585
R9231 GND.n1031 GND.n1030 585
R9232 GND.n6749 GND.n1031 585
R9233 GND.n6752 GND.n6751 585
R9234 GND.n6751 GND.n6750 585
R9235 GND.n1028 GND.n1027 585
R9236 GND.n1027 GND.n1026 585
R9237 GND.n6757 GND.n6756 585
R9238 GND.n6758 GND.n6757 585
R9239 GND.n1025 GND.n1024 585
R9240 GND.n6759 GND.n1025 585
R9241 GND.n6762 GND.n6761 585
R9242 GND.n6761 GND.n6760 585
R9243 GND.n1022 GND.n1021 585
R9244 GND.n1021 GND.n1020 585
R9245 GND.n6767 GND.n6766 585
R9246 GND.n6768 GND.n6767 585
R9247 GND.n1019 GND.n1018 585
R9248 GND.n6769 GND.n1019 585
R9249 GND.n6772 GND.n6771 585
R9250 GND.n6771 GND.n6770 585
R9251 GND.n1016 GND.n1015 585
R9252 GND.n1015 GND.n1014 585
R9253 GND.n6777 GND.n6776 585
R9254 GND.n6778 GND.n6777 585
R9255 GND.n1013 GND.n1012 585
R9256 GND.n6779 GND.n1013 585
R9257 GND.n6782 GND.n6781 585
R9258 GND.n6781 GND.n6780 585
R9259 GND.n1010 GND.n1009 585
R9260 GND.n1009 GND.n1008 585
R9261 GND.n6787 GND.n6786 585
R9262 GND.n6788 GND.n6787 585
R9263 GND.n1007 GND.n1006 585
R9264 GND.n6789 GND.n1007 585
R9265 GND.n6792 GND.n6791 585
R9266 GND.n6791 GND.n6790 585
R9267 GND.n1004 GND.n1003 585
R9268 GND.n1003 GND.n1002 585
R9269 GND.n6797 GND.n6796 585
R9270 GND.n6798 GND.n6797 585
R9271 GND.n1001 GND.n1000 585
R9272 GND.n6799 GND.n1001 585
R9273 GND.n6802 GND.n6801 585
R9274 GND.n6801 GND.n6800 585
R9275 GND.n998 GND.n997 585
R9276 GND.n997 GND.n996 585
R9277 GND.n6807 GND.n6806 585
R9278 GND.n6808 GND.n6807 585
R9279 GND.n995 GND.n994 585
R9280 GND.n6809 GND.n995 585
R9281 GND.n6812 GND.n6811 585
R9282 GND.n6811 GND.n6810 585
R9283 GND.n992 GND.n991 585
R9284 GND.n991 GND.n990 585
R9285 GND.n6817 GND.n6816 585
R9286 GND.n6818 GND.n6817 585
R9287 GND.n989 GND.n988 585
R9288 GND.n6819 GND.n989 585
R9289 GND.n6822 GND.n6821 585
R9290 GND.n6821 GND.n6820 585
R9291 GND.n986 GND.n985 585
R9292 GND.n985 GND.n984 585
R9293 GND.n6827 GND.n6826 585
R9294 GND.n6828 GND.n6827 585
R9295 GND.n983 GND.n982 585
R9296 GND.n6829 GND.n983 585
R9297 GND.n6832 GND.n6831 585
R9298 GND.n6831 GND.n6830 585
R9299 GND.n980 GND.n979 585
R9300 GND.n979 GND.n978 585
R9301 GND.n6837 GND.n6836 585
R9302 GND.n6838 GND.n6837 585
R9303 GND.n977 GND.n976 585
R9304 GND.n6839 GND.n977 585
R9305 GND.n6842 GND.n6841 585
R9306 GND.n6841 GND.n6840 585
R9307 GND.n974 GND.n973 585
R9308 GND.n973 GND.n972 585
R9309 GND.n6847 GND.n6846 585
R9310 GND.n6848 GND.n6847 585
R9311 GND.n971 GND.n970 585
R9312 GND.n6849 GND.n971 585
R9313 GND.n6852 GND.n6851 585
R9314 GND.n6851 GND.n6850 585
R9315 GND.n968 GND.n967 585
R9316 GND.n967 GND.n966 585
R9317 GND.n6857 GND.n6856 585
R9318 GND.n6858 GND.n6857 585
R9319 GND.n965 GND.n964 585
R9320 GND.n6859 GND.n965 585
R9321 GND.n6862 GND.n6861 585
R9322 GND.n6861 GND.n6860 585
R9323 GND.n962 GND.n961 585
R9324 GND.n961 GND.n960 585
R9325 GND.n6867 GND.n6866 585
R9326 GND.n6868 GND.n6867 585
R9327 GND.n959 GND.n958 585
R9328 GND.n6869 GND.n959 585
R9329 GND.n6872 GND.n6871 585
R9330 GND.n6871 GND.n6870 585
R9331 GND.n956 GND.n955 585
R9332 GND.n955 GND.n954 585
R9333 GND.n6877 GND.n6876 585
R9334 GND.n6878 GND.n6877 585
R9335 GND.n953 GND.n952 585
R9336 GND.n6879 GND.n953 585
R9337 GND.n6882 GND.n6881 585
R9338 GND.n6881 GND.n6880 585
R9339 GND.n950 GND.n949 585
R9340 GND.n949 GND.n948 585
R9341 GND.n6887 GND.n6886 585
R9342 GND.n6888 GND.n6887 585
R9343 GND.n947 GND.n946 585
R9344 GND.n6889 GND.n947 585
R9345 GND.n6892 GND.n6891 585
R9346 GND.n6891 GND.n6890 585
R9347 GND.n944 GND.n943 585
R9348 GND.n943 GND.n942 585
R9349 GND.n6897 GND.n6896 585
R9350 GND.n6898 GND.n6897 585
R9351 GND.n941 GND.n940 585
R9352 GND.n6899 GND.n941 585
R9353 GND.n6902 GND.n6901 585
R9354 GND.n6901 GND.n6900 585
R9355 GND.n938 GND.n937 585
R9356 GND.n937 GND.n936 585
R9357 GND.n6907 GND.n6906 585
R9358 GND.n6908 GND.n6907 585
R9359 GND.n935 GND.n934 585
R9360 GND.n6909 GND.n935 585
R9361 GND.n6912 GND.n6911 585
R9362 GND.n6911 GND.n6910 585
R9363 GND.n932 GND.n931 585
R9364 GND.n931 GND.n930 585
R9365 GND.n6917 GND.n6916 585
R9366 GND.n6918 GND.n6917 585
R9367 GND.n929 GND.n928 585
R9368 GND.n6919 GND.n929 585
R9369 GND.n6922 GND.n6921 585
R9370 GND.n6921 GND.n6920 585
R9371 GND.n926 GND.n925 585
R9372 GND.n925 GND.n924 585
R9373 GND.n6927 GND.n6926 585
R9374 GND.n6928 GND.n6927 585
R9375 GND.n923 GND.n922 585
R9376 GND.n6929 GND.n923 585
R9377 GND.n6932 GND.n6931 585
R9378 GND.n6931 GND.n6930 585
R9379 GND.n920 GND.n919 585
R9380 GND.n919 GND.n918 585
R9381 GND.n6937 GND.n6936 585
R9382 GND.n6938 GND.n6937 585
R9383 GND.n917 GND.n916 585
R9384 GND.n6939 GND.n917 585
R9385 GND.n6942 GND.n6941 585
R9386 GND.n6941 GND.n6940 585
R9387 GND.n914 GND.n913 585
R9388 GND.n913 GND.n912 585
R9389 GND.n6947 GND.n6946 585
R9390 GND.n6948 GND.n6947 585
R9391 GND.n911 GND.n910 585
R9392 GND.n6949 GND.n911 585
R9393 GND.n6952 GND.n6951 585
R9394 GND.n6951 GND.n6950 585
R9395 GND.n908 GND.n907 585
R9396 GND.n907 GND.n906 585
R9397 GND.n6957 GND.n6956 585
R9398 GND.n6958 GND.n6957 585
R9399 GND.n905 GND.n904 585
R9400 GND.n6959 GND.n905 585
R9401 GND.n6962 GND.n6961 585
R9402 GND.n6961 GND.n6960 585
R9403 GND.n902 GND.n901 585
R9404 GND.n901 GND.n900 585
R9405 GND.n6967 GND.n6966 585
R9406 GND.n6968 GND.n6967 585
R9407 GND.n899 GND.n898 585
R9408 GND.n6969 GND.n899 585
R9409 GND.n6972 GND.n6971 585
R9410 GND.n6971 GND.n6970 585
R9411 GND.n896 GND.n895 585
R9412 GND.n895 GND.n894 585
R9413 GND.n6977 GND.n6976 585
R9414 GND.n6978 GND.n6977 585
R9415 GND.n893 GND.n892 585
R9416 GND.n6979 GND.n893 585
R9417 GND.n6982 GND.n6981 585
R9418 GND.n6981 GND.n6980 585
R9419 GND.n890 GND.n889 585
R9420 GND.n889 GND.n888 585
R9421 GND.n6987 GND.n6986 585
R9422 GND.n6988 GND.n6987 585
R9423 GND.n887 GND.n886 585
R9424 GND.n6989 GND.n887 585
R9425 GND.n6992 GND.n6991 585
R9426 GND.n6991 GND.n6990 585
R9427 GND.n884 GND.n883 585
R9428 GND.n883 GND.n882 585
R9429 GND.n6997 GND.n6996 585
R9430 GND.n6998 GND.n6997 585
R9431 GND.n881 GND.n880 585
R9432 GND.n6999 GND.n881 585
R9433 GND.n7002 GND.n7001 585
R9434 GND.n7001 GND.n7000 585
R9435 GND.n878 GND.n877 585
R9436 GND.n877 GND.n876 585
R9437 GND.n7007 GND.n7006 585
R9438 GND.n7008 GND.n7007 585
R9439 GND.n875 GND.n874 585
R9440 GND.n7009 GND.n875 585
R9441 GND.n7012 GND.n7011 585
R9442 GND.n7011 GND.n7010 585
R9443 GND.n872 GND.n871 585
R9444 GND.n871 GND.n870 585
R9445 GND.n7017 GND.n7016 585
R9446 GND.n7018 GND.n7017 585
R9447 GND.n869 GND.n868 585
R9448 GND.n7019 GND.n869 585
R9449 GND.n7022 GND.n7021 585
R9450 GND.n7021 GND.n7020 585
R9451 GND.n866 GND.n865 585
R9452 GND.n865 GND.n864 585
R9453 GND.n7027 GND.n7026 585
R9454 GND.n7028 GND.n7027 585
R9455 GND.n863 GND.n862 585
R9456 GND.n7029 GND.n863 585
R9457 GND.n7032 GND.n7031 585
R9458 GND.n7031 GND.n7030 585
R9459 GND.n860 GND.n859 585
R9460 GND.n859 GND.n858 585
R9461 GND.n7037 GND.n7036 585
R9462 GND.n7038 GND.n7037 585
R9463 GND.n857 GND.n856 585
R9464 GND.n7039 GND.n857 585
R9465 GND.n7042 GND.n7041 585
R9466 GND.n7041 GND.n7040 585
R9467 GND.n854 GND.n853 585
R9468 GND.n853 GND.n852 585
R9469 GND.n7047 GND.n7046 585
R9470 GND.n7048 GND.n7047 585
R9471 GND.n851 GND.n850 585
R9472 GND.n7049 GND.n851 585
R9473 GND.n7052 GND.n7051 585
R9474 GND.n7051 GND.n7050 585
R9475 GND.n848 GND.n847 585
R9476 GND.n847 GND.n846 585
R9477 GND.n7057 GND.n7056 585
R9478 GND.n7058 GND.n7057 585
R9479 GND.n845 GND.n844 585
R9480 GND.n7059 GND.n845 585
R9481 GND.n7062 GND.n7061 585
R9482 GND.n7061 GND.n7060 585
R9483 GND.n842 GND.n841 585
R9484 GND.n841 GND.n840 585
R9485 GND.n7067 GND.n7066 585
R9486 GND.n7068 GND.n7067 585
R9487 GND.n839 GND.n838 585
R9488 GND.n7069 GND.n839 585
R9489 GND.n7072 GND.n7071 585
R9490 GND.n7071 GND.n7070 585
R9491 GND.n836 GND.n835 585
R9492 GND.n835 GND.n834 585
R9493 GND.n7077 GND.n7076 585
R9494 GND.n7078 GND.n7077 585
R9495 GND.n833 GND.n832 585
R9496 GND.n7079 GND.n833 585
R9497 GND.n7082 GND.n7081 585
R9498 GND.n7081 GND.n7080 585
R9499 GND.n830 GND.n829 585
R9500 GND.n829 GND.n828 585
R9501 GND.n7087 GND.n7086 585
R9502 GND.n7088 GND.n7087 585
R9503 GND.n827 GND.n826 585
R9504 GND.n7089 GND.n827 585
R9505 GND.n7092 GND.n7091 585
R9506 GND.n7091 GND.n7090 585
R9507 GND.n824 GND.n823 585
R9508 GND.n823 GND.n822 585
R9509 GND.n7097 GND.n7096 585
R9510 GND.n7098 GND.n7097 585
R9511 GND.n821 GND.n820 585
R9512 GND.n7099 GND.n821 585
R9513 GND.n7102 GND.n7101 585
R9514 GND.n7101 GND.n7100 585
R9515 GND.n818 GND.n817 585
R9516 GND.n817 GND.n816 585
R9517 GND.n7107 GND.n7106 585
R9518 GND.n7108 GND.n7107 585
R9519 GND.n815 GND.n814 585
R9520 GND.n7109 GND.n815 585
R9521 GND.n7112 GND.n7111 585
R9522 GND.n7111 GND.n7110 585
R9523 GND.n812 GND.n811 585
R9524 GND.n811 GND.n810 585
R9525 GND.n7117 GND.n7116 585
R9526 GND.n7118 GND.n7117 585
R9527 GND.n809 GND.n808 585
R9528 GND.n7119 GND.n809 585
R9529 GND.n7122 GND.n7121 585
R9530 GND.n7121 GND.n7120 585
R9531 GND.n806 GND.n805 585
R9532 GND.n805 GND.n804 585
R9533 GND.n7127 GND.n7126 585
R9534 GND.n7128 GND.n7127 585
R9535 GND.n803 GND.n802 585
R9536 GND.n7129 GND.n803 585
R9537 GND.n7132 GND.n7131 585
R9538 GND.n7131 GND.n7130 585
R9539 GND.n800 GND.n799 585
R9540 GND.n799 GND.n798 585
R9541 GND.n7137 GND.n7136 585
R9542 GND.n7138 GND.n7137 585
R9543 GND.n797 GND.n796 585
R9544 GND.n7139 GND.n797 585
R9545 GND.n7142 GND.n7141 585
R9546 GND.n7141 GND.n7140 585
R9547 GND.n794 GND.n793 585
R9548 GND.n793 GND.n792 585
R9549 GND.n7147 GND.n7146 585
R9550 GND.n7148 GND.n7147 585
R9551 GND.n791 GND.n790 585
R9552 GND.n7149 GND.n791 585
R9553 GND.n7152 GND.n7151 585
R9554 GND.n7151 GND.n7150 585
R9555 GND.n788 GND.n787 585
R9556 GND.n787 GND.n786 585
R9557 GND.n7157 GND.n7156 585
R9558 GND.n7158 GND.n7157 585
R9559 GND.n785 GND.n784 585
R9560 GND.n7159 GND.n785 585
R9561 GND.n7162 GND.n7161 585
R9562 GND.n7161 GND.n7160 585
R9563 GND.n782 GND.n781 585
R9564 GND.n781 GND.n780 585
R9565 GND.n7167 GND.n7166 585
R9566 GND.n7168 GND.n7167 585
R9567 GND.n779 GND.n778 585
R9568 GND.n7169 GND.n779 585
R9569 GND.n7172 GND.n7171 585
R9570 GND.n7171 GND.n7170 585
R9571 GND.n776 GND.n775 585
R9572 GND.n775 GND.n774 585
R9573 GND.n7177 GND.n7176 585
R9574 GND.n7178 GND.n7177 585
R9575 GND.n773 GND.n772 585
R9576 GND.n7179 GND.n773 585
R9577 GND.n7182 GND.n7181 585
R9578 GND.n7181 GND.n7180 585
R9579 GND.n770 GND.n769 585
R9580 GND.n769 GND.n768 585
R9581 GND.n7187 GND.n7186 585
R9582 GND.n7188 GND.n7187 585
R9583 GND.n767 GND.n766 585
R9584 GND.n7189 GND.n767 585
R9585 GND.n7192 GND.n7191 585
R9586 GND.n7191 GND.n7190 585
R9587 GND.n764 GND.n763 585
R9588 GND.n763 GND.n762 585
R9589 GND.n7197 GND.n7196 585
R9590 GND.n7198 GND.n7197 585
R9591 GND.n761 GND.n760 585
R9592 GND.n7199 GND.n761 585
R9593 GND.n7202 GND.n7201 585
R9594 GND.n7201 GND.n7200 585
R9595 GND.n758 GND.n757 585
R9596 GND.n757 GND.n756 585
R9597 GND.n7207 GND.n7206 585
R9598 GND.n7208 GND.n7207 585
R9599 GND.n755 GND.n754 585
R9600 GND.n7209 GND.n755 585
R9601 GND.n7212 GND.n7211 585
R9602 GND.n7211 GND.n7210 585
R9603 GND.n752 GND.n751 585
R9604 GND.n751 GND.n750 585
R9605 GND.n7217 GND.n7216 585
R9606 GND.n7218 GND.n7217 585
R9607 GND.n749 GND.n748 585
R9608 GND.n7219 GND.n749 585
R9609 GND.n7222 GND.n7221 585
R9610 GND.n7221 GND.n7220 585
R9611 GND.n746 GND.n745 585
R9612 GND.n745 GND.n744 585
R9613 GND.n7227 GND.n7226 585
R9614 GND.n7228 GND.n7227 585
R9615 GND.n743 GND.n742 585
R9616 GND.n7229 GND.n743 585
R9617 GND.n7232 GND.n7231 585
R9618 GND.n7231 GND.n7230 585
R9619 GND.n740 GND.n739 585
R9620 GND.n739 GND.n738 585
R9621 GND.n7237 GND.n7236 585
R9622 GND.n7238 GND.n7237 585
R9623 GND.n737 GND.n736 585
R9624 GND.n7239 GND.n737 585
R9625 GND.n7242 GND.n7241 585
R9626 GND.n7241 GND.n7240 585
R9627 GND.n734 GND.n733 585
R9628 GND.n733 GND.n732 585
R9629 GND.n7247 GND.n7246 585
R9630 GND.n7248 GND.n7247 585
R9631 GND.n731 GND.n730 585
R9632 GND.n7249 GND.n731 585
R9633 GND.n7252 GND.n7251 585
R9634 GND.n7251 GND.n7250 585
R9635 GND.n728 GND.n727 585
R9636 GND.n727 GND.n726 585
R9637 GND.n7257 GND.n7256 585
R9638 GND.n7258 GND.n7257 585
R9639 GND.n725 GND.n724 585
R9640 GND.n7259 GND.n725 585
R9641 GND.n7262 GND.n7261 585
R9642 GND.n7261 GND.n7260 585
R9643 GND.n722 GND.n721 585
R9644 GND.n721 GND.n720 585
R9645 GND.n7267 GND.n7266 585
R9646 GND.n7268 GND.n7267 585
R9647 GND.n719 GND.n718 585
R9648 GND.n7269 GND.n719 585
R9649 GND.n7272 GND.n7271 585
R9650 GND.n7271 GND.n7270 585
R9651 GND.n716 GND.n715 585
R9652 GND.n715 GND.n714 585
R9653 GND.n7277 GND.n7276 585
R9654 GND.n7278 GND.n7277 585
R9655 GND.n713 GND.n712 585
R9656 GND.n7279 GND.n713 585
R9657 GND.n7282 GND.n7281 585
R9658 GND.n7281 GND.n7280 585
R9659 GND.n710 GND.n709 585
R9660 GND.n709 GND.n708 585
R9661 GND.n7287 GND.n7286 585
R9662 GND.n7288 GND.n7287 585
R9663 GND.n707 GND.n706 585
R9664 GND.n7289 GND.n707 585
R9665 GND.n7292 GND.n7291 585
R9666 GND.n7291 GND.n7290 585
R9667 GND.n704 GND.n703 585
R9668 GND.n703 GND.n702 585
R9669 GND.n7297 GND.n7296 585
R9670 GND.n7298 GND.n7297 585
R9671 GND.n701 GND.n700 585
R9672 GND.n7299 GND.n701 585
R9673 GND.n7302 GND.n7301 585
R9674 GND.n7301 GND.n7300 585
R9675 GND.n698 GND.n697 585
R9676 GND.n697 GND.n696 585
R9677 GND.n7307 GND.n7306 585
R9678 GND.n7308 GND.n7307 585
R9679 GND.n695 GND.n694 585
R9680 GND.n7309 GND.n695 585
R9681 GND.n7312 GND.n7311 585
R9682 GND.n7311 GND.n7310 585
R9683 GND.n692 GND.n691 585
R9684 GND.n691 GND.n690 585
R9685 GND.n7317 GND.n7316 585
R9686 GND.n7318 GND.n7317 585
R9687 GND.n689 GND.n688 585
R9688 GND.n7319 GND.n689 585
R9689 GND.n7322 GND.n7321 585
R9690 GND.n7321 GND.n7320 585
R9691 GND.n686 GND.n685 585
R9692 GND.n685 GND.n684 585
R9693 GND.n7328 GND.n7327 585
R9694 GND.n7329 GND.n7328 585
R9695 GND.n683 GND.n682 585
R9696 GND.n7330 GND.n683 585
R9697 GND.n7333 GND.n7332 585
R9698 GND.n7332 GND.n7331 585
R9699 GND.n7334 GND.n680 585
R9700 GND.n680 GND.n679 585
R9701 GND.n7558 GND.n546 585
R9702 GND.n7562 GND.n546 585
R9703 GND.n7560 GND.n7559 585
R9704 GND.n7561 GND.n7560 585
R9705 GND.n549 GND.n548 585
R9706 GND.n548 GND.n547 585
R9707 GND.n7553 GND.n7552 585
R9708 GND.n7552 GND.n7551 585
R9709 GND.n552 GND.n551 585
R9710 GND.n7550 GND.n552 585
R9711 GND.n7548 GND.n7547 585
R9712 GND.n7549 GND.n7548 585
R9713 GND.n555 GND.n554 585
R9714 GND.n554 GND.n553 585
R9715 GND.n7543 GND.n7542 585
R9716 GND.n7542 GND.n7541 585
R9717 GND.n558 GND.n557 585
R9718 GND.n7540 GND.n558 585
R9719 GND.n7538 GND.n7537 585
R9720 GND.n7539 GND.n7538 585
R9721 GND.n561 GND.n560 585
R9722 GND.n560 GND.n559 585
R9723 GND.n7533 GND.n7532 585
R9724 GND.n7532 GND.n7531 585
R9725 GND.n564 GND.n563 585
R9726 GND.n7530 GND.n564 585
R9727 GND.n7528 GND.n7527 585
R9728 GND.n7529 GND.n7528 585
R9729 GND.n567 GND.n566 585
R9730 GND.n566 GND.n565 585
R9731 GND.n7523 GND.n7522 585
R9732 GND.n7522 GND.n7521 585
R9733 GND.n570 GND.n569 585
R9734 GND.n7520 GND.n570 585
R9735 GND.n7518 GND.n7517 585
R9736 GND.n7519 GND.n7518 585
R9737 GND.n573 GND.n572 585
R9738 GND.n572 GND.n571 585
R9739 GND.n7513 GND.n7512 585
R9740 GND.n7512 GND.n7511 585
R9741 GND.n576 GND.n575 585
R9742 GND.n7510 GND.n576 585
R9743 GND.n7508 GND.n7507 585
R9744 GND.n7509 GND.n7508 585
R9745 GND.n579 GND.n578 585
R9746 GND.n578 GND.n577 585
R9747 GND.n7503 GND.n7502 585
R9748 GND.n7502 GND.n7501 585
R9749 GND.n582 GND.n581 585
R9750 GND.n7500 GND.n582 585
R9751 GND.n7498 GND.n7497 585
R9752 GND.n7499 GND.n7498 585
R9753 GND.n585 GND.n584 585
R9754 GND.n584 GND.n583 585
R9755 GND.n7493 GND.n7492 585
R9756 GND.n7492 GND.n7491 585
R9757 GND.n588 GND.n587 585
R9758 GND.n7490 GND.n588 585
R9759 GND.n7488 GND.n7487 585
R9760 GND.n7489 GND.n7488 585
R9761 GND.n591 GND.n590 585
R9762 GND.n590 GND.n589 585
R9763 GND.n7483 GND.n7482 585
R9764 GND.n7482 GND.n7481 585
R9765 GND.n594 GND.n593 585
R9766 GND.n7480 GND.n594 585
R9767 GND.n7478 GND.n7477 585
R9768 GND.n7479 GND.n7478 585
R9769 GND.n597 GND.n596 585
R9770 GND.n596 GND.n595 585
R9771 GND.n7473 GND.n7472 585
R9772 GND.n7472 GND.n7471 585
R9773 GND.n600 GND.n599 585
R9774 GND.n7470 GND.n600 585
R9775 GND.n7468 GND.n7467 585
R9776 GND.n7469 GND.n7468 585
R9777 GND.n603 GND.n602 585
R9778 GND.n602 GND.n601 585
R9779 GND.n7463 GND.n7462 585
R9780 GND.n7462 GND.n7461 585
R9781 GND.n606 GND.n605 585
R9782 GND.n7460 GND.n606 585
R9783 GND.n7458 GND.n7457 585
R9784 GND.n7459 GND.n7458 585
R9785 GND.n609 GND.n608 585
R9786 GND.n608 GND.n607 585
R9787 GND.n7453 GND.n7452 585
R9788 GND.n7452 GND.n7451 585
R9789 GND.n612 GND.n611 585
R9790 GND.n7450 GND.n612 585
R9791 GND.n7448 GND.n7447 585
R9792 GND.n7449 GND.n7448 585
R9793 GND.n615 GND.n614 585
R9794 GND.n614 GND.n613 585
R9795 GND.n7443 GND.n7442 585
R9796 GND.n7442 GND.n7441 585
R9797 GND.n618 GND.n617 585
R9798 GND.n7440 GND.n618 585
R9799 GND.n7438 GND.n7437 585
R9800 GND.n7439 GND.n7438 585
R9801 GND.n621 GND.n620 585
R9802 GND.n620 GND.n619 585
R9803 GND.n7433 GND.n7432 585
R9804 GND.n7432 GND.n7431 585
R9805 GND.n624 GND.n623 585
R9806 GND.n7430 GND.n624 585
R9807 GND.n7428 GND.n7427 585
R9808 GND.n7429 GND.n7428 585
R9809 GND.n627 GND.n626 585
R9810 GND.n626 GND.n625 585
R9811 GND.n7423 GND.n7422 585
R9812 GND.n7422 GND.n7421 585
R9813 GND.n630 GND.n629 585
R9814 GND.n7420 GND.n630 585
R9815 GND.n7418 GND.n7417 585
R9816 GND.n7419 GND.n7418 585
R9817 GND.n633 GND.n632 585
R9818 GND.n632 GND.n631 585
R9819 GND.n7413 GND.n7412 585
R9820 GND.n7412 GND.n7411 585
R9821 GND.n636 GND.n635 585
R9822 GND.n7410 GND.n636 585
R9823 GND.n7408 GND.n7407 585
R9824 GND.n7409 GND.n7408 585
R9825 GND.n639 GND.n638 585
R9826 GND.n638 GND.n637 585
R9827 GND.n7403 GND.n7402 585
R9828 GND.n7402 GND.n7401 585
R9829 GND.n642 GND.n641 585
R9830 GND.n7400 GND.n642 585
R9831 GND.n7398 GND.n7397 585
R9832 GND.n7399 GND.n7398 585
R9833 GND.n645 GND.n644 585
R9834 GND.n644 GND.n643 585
R9835 GND.n7393 GND.n7392 585
R9836 GND.n7392 GND.n7391 585
R9837 GND.n648 GND.n647 585
R9838 GND.n7390 GND.n648 585
R9839 GND.n7388 GND.n7387 585
R9840 GND.n7389 GND.n7388 585
R9841 GND.n651 GND.n650 585
R9842 GND.n650 GND.n649 585
R9843 GND.n7383 GND.n7382 585
R9844 GND.n7382 GND.n7381 585
R9845 GND.n654 GND.n653 585
R9846 GND.n7380 GND.n654 585
R9847 GND.n7378 GND.n7377 585
R9848 GND.n7379 GND.n7378 585
R9849 GND.n657 GND.n656 585
R9850 GND.n656 GND.n655 585
R9851 GND.n7373 GND.n7372 585
R9852 GND.n7372 GND.n7371 585
R9853 GND.n660 GND.n659 585
R9854 GND.n7370 GND.n660 585
R9855 GND.n7368 GND.n7367 585
R9856 GND.n7369 GND.n7368 585
R9857 GND.n663 GND.n662 585
R9858 GND.n662 GND.n661 585
R9859 GND.n7363 GND.n7362 585
R9860 GND.n7362 GND.n7361 585
R9861 GND.n666 GND.n665 585
R9862 GND.n7360 GND.n666 585
R9863 GND.n7358 GND.n7357 585
R9864 GND.n7359 GND.n7358 585
R9865 GND.n669 GND.n668 585
R9866 GND.n668 GND.n667 585
R9867 GND.n7353 GND.n7352 585
R9868 GND.n7352 GND.n7351 585
R9869 GND.n672 GND.n671 585
R9870 GND.n7350 GND.n672 585
R9871 GND.n7348 GND.n7347 585
R9872 GND.n7349 GND.n7348 585
R9873 GND.n675 GND.n674 585
R9874 GND.n674 GND.n673 585
R9875 GND.n7343 GND.n7342 585
R9876 GND.n7342 GND.n7341 585
R9877 GND.n678 GND.n677 585
R9878 GND.n7340 GND.n678 585
R9879 GND.n7338 GND.n7337 585
R9880 GND.n7339 GND.n7338 585
R9881 GND.n7742 GND.n176 585
R9882 GND.n7738 GND.n176 585
R9883 GND.n7744 GND.n7743 585
R9884 GND.n7745 GND.n7744 585
R9885 GND.n160 GND.n159 585
R9886 GND.n5161 GND.n160 585
R9887 GND.n7753 GND.n7752 585
R9888 GND.n7752 GND.n7751 585
R9889 GND.n7754 GND.n155 585
R9890 GND.n5167 GND.n155 585
R9891 GND.n7756 GND.n7755 585
R9892 GND.n7757 GND.n7756 585
R9893 GND.n140 GND.n139 585
R9894 GND.n5173 GND.n140 585
R9895 GND.n7765 GND.n7764 585
R9896 GND.n7764 GND.n7763 585
R9897 GND.n7766 GND.n135 585
R9898 GND.n5179 GND.n135 585
R9899 GND.n7768 GND.n7767 585
R9900 GND.n7769 GND.n7768 585
R9901 GND.n119 GND.n118 585
R9902 GND.n5098 GND.n119 585
R9903 GND.n7777 GND.n7776 585
R9904 GND.n7776 GND.n7775 585
R9905 GND.n7778 GND.n114 585
R9906 GND.n5089 GND.n114 585
R9907 GND.n7780 GND.n7779 585
R9908 GND.n7781 GND.n7780 585
R9909 GND.n98 GND.n97 585
R9910 GND.n5083 GND.n98 585
R9911 GND.n7789 GND.n7788 585
R9912 GND.n7788 GND.n7787 585
R9913 GND.n7790 GND.n93 585
R9914 GND.n5075 GND.n93 585
R9915 GND.n7792 GND.n7791 585
R9916 GND.n7793 GND.n7792 585
R9917 GND.n77 GND.n76 585
R9918 GND.n5069 GND.n77 585
R9919 GND.n7801 GND.n7800 585
R9920 GND.n7800 GND.n7799 585
R9921 GND.n7802 GND.n72 585
R9922 GND.n5061 GND.n72 585
R9923 GND.n7804 GND.n7803 585
R9924 GND.n7805 GND.n7804 585
R9925 GND.n58 GND.n57 585
R9926 GND.n5055 GND.n58 585
R9927 GND.n7813 GND.n7812 585
R9928 GND.n7812 GND.n7811 585
R9929 GND.n7814 GND.n52 585
R9930 GND.n5047 GND.n52 585
R9931 GND.n7816 GND.n7815 585
R9932 GND.n7817 GND.n7816 585
R9933 GND.n53 GND.n51 585
R9934 GND.n5040 GND.n51 585
R9935 GND.n2755 GND.n2754 585
R9936 GND.n2759 GND.n2755 585
R9937 GND.n5240 GND.n5239 585
R9938 GND.n5239 GND.n5238 585
R9939 GND.n5241 GND.n31 585
R9940 GND.n7824 GND.n31 585
R9941 GND.n5243 GND.n5242 585
R9942 GND.n5244 GND.n5243 585
R9943 GND.n2750 GND.n2749 585
R9944 GND.n2749 GND.n2747 585
R9945 GND.n5020 GND.n5019 585
R9946 GND.n5019 GND.n2738 585
R9947 GND.n2729 GND.n2728 585
R9948 GND.n5253 GND.n2729 585
R9949 GND.n5259 GND.n5258 585
R9950 GND.n5258 GND.n5257 585
R9951 GND.n5260 GND.n2724 585
R9952 GND.n5013 GND.n2724 585
R9953 GND.n5262 GND.n5261 585
R9954 GND.n5263 GND.n5262 585
R9955 GND.n2709 GND.n2708 585
R9956 GND.n4995 GND.n2709 585
R9957 GND.n5271 GND.n5270 585
R9958 GND.n5270 GND.n5269 585
R9959 GND.n5272 GND.n2704 585
R9960 GND.n4988 GND.n2704 585
R9961 GND.n5274 GND.n5273 585
R9962 GND.n5275 GND.n5274 585
R9963 GND.n2688 GND.n2687 585
R9964 GND.n4980 GND.n2688 585
R9965 GND.n5283 GND.n5282 585
R9966 GND.n5282 GND.n5281 585
R9967 GND.n5284 GND.n2683 585
R9968 GND.n4973 GND.n2683 585
R9969 GND.n5286 GND.n5285 585
R9970 GND.n5287 GND.n5286 585
R9971 GND.n2667 GND.n2666 585
R9972 GND.n4965 GND.n2667 585
R9973 GND.n5295 GND.n5294 585
R9974 GND.n5294 GND.n5293 585
R9975 GND.n5296 GND.n2662 585
R9976 GND.n4958 GND.n2662 585
R9977 GND.n5298 GND.n5297 585
R9978 GND.n5299 GND.n5298 585
R9979 GND.n2646 GND.n2645 585
R9980 GND.n4950 GND.n2646 585
R9981 GND.n5307 GND.n5306 585
R9982 GND.n5306 GND.n5305 585
R9983 GND.n5308 GND.n2640 585
R9984 GND.n4943 GND.n2640 585
R9985 GND.n5310 GND.n5309 585
R9986 GND.n5311 GND.n5310 585
R9987 GND.n2641 GND.n2639 585
R9988 GND.n4935 GND.n2639 585
R9989 GND.n4930 GND.n2622 585
R9990 GND.n5317 GND.n2622 585
R9991 GND.n4929 GND.n4928 585
R9992 GND.n4928 GND.n2618 585
R9993 GND.n4927 GND.n4926 585
R9994 GND.n4927 GND.n2608 585
R9995 GND.n2601 GND.n2599 585
R9996 GND.n5325 GND.n2599 585
R9997 GND.n5331 GND.n5330 585
R9998 GND.n5332 GND.n5331 585
R9999 GND.n2600 GND.n2598 585
R10000 GND.n4909 GND.n2598 585
R10001 GND.n2903 GND.n2902 585
R10002 GND.n2907 GND.n2905 585
R10003 GND.n2909 GND.n2908 585
R10004 GND.n2913 GND.n2911 585
R10005 GND.n2915 GND.n2914 585
R10006 GND.n2919 GND.n2917 585
R10007 GND.n2921 GND.n2920 585
R10008 GND.n2925 GND.n2923 585
R10009 GND.n2927 GND.n2926 585
R10010 GND.n2930 GND.n2928 585
R10011 GND.n2931 GND.n2897 585
R10012 GND.n4801 GND.n4800 585
R10013 GND.n5153 GND.n5152 585
R10014 GND.n5150 GND.n5114 585
R10015 GND.n5149 GND.n5148 585
R10016 GND.n5142 GND.n5116 585
R10017 GND.n5144 GND.n5143 585
R10018 GND.n5140 GND.n5118 585
R10019 GND.n5139 GND.n5138 585
R10020 GND.n5132 GND.n5120 585
R10021 GND.n5134 GND.n5133 585
R10022 GND.n5130 GND.n5122 585
R10023 GND.n5129 GND.n5128 585
R10024 GND.n5125 GND.n5124 585
R10025 GND.n5156 GND.n181 585
R10026 GND.n7738 GND.n181 585
R10027 GND.n5157 GND.n174 585
R10028 GND.n7745 GND.n174 585
R10029 GND.n5163 GND.n5162 585
R10030 GND.n5162 GND.n5161 585
R10031 GND.n5164 GND.n163 585
R10032 GND.n7751 GND.n163 585
R10033 GND.n5166 GND.n5165 585
R10034 GND.n5167 GND.n5166 585
R10035 GND.n2792 GND.n153 585
R10036 GND.n7757 GND.n153 585
R10037 GND.n5175 GND.n5174 585
R10038 GND.n5174 GND.n5173 585
R10039 GND.n5176 GND.n142 585
R10040 GND.n7763 GND.n142 585
R10041 GND.n5178 GND.n5177 585
R10042 GND.n5179 GND.n5178 585
R10043 GND.n2788 GND.n133 585
R10044 GND.n7769 GND.n133 585
R10045 GND.n5097 GND.n5096 585
R10046 GND.n5098 GND.n5097 585
R10047 GND.n2795 GND.n122 585
R10048 GND.n7775 GND.n122 585
R10049 GND.n5091 GND.n5090 585
R10050 GND.n5090 GND.n5089 585
R10051 GND.n2797 GND.n112 585
R10052 GND.n7781 GND.n112 585
R10053 GND.n5082 GND.n5081 585
R10054 GND.n5083 GND.n5082 585
R10055 GND.n2800 GND.n101 585
R10056 GND.n7787 GND.n101 585
R10057 GND.n5077 GND.n5076 585
R10058 GND.n5076 GND.n5075 585
R10059 GND.n2802 GND.n91 585
R10060 GND.n7793 GND.n91 585
R10061 GND.n5068 GND.n5067 585
R10062 GND.n5069 GND.n5068 585
R10063 GND.n2805 GND.n80 585
R10064 GND.n7799 GND.n80 585
R10065 GND.n5063 GND.n5062 585
R10066 GND.n5062 GND.n5061 585
R10067 GND.n2807 GND.n70 585
R10068 GND.n7805 GND.n70 585
R10069 GND.n5054 GND.n5053 585
R10070 GND.n5055 GND.n5054 585
R10071 GND.n2810 GND.n60 585
R10072 GND.n7811 GND.n60 585
R10073 GND.n5049 GND.n5048 585
R10074 GND.n5048 GND.n5047 585
R10075 GND.n2812 GND.n49 585
R10076 GND.n7817 GND.n49 585
R10077 GND.n5039 GND.n5038 585
R10078 GND.n5040 GND.n5039 585
R10079 GND.n5035 GND.n5034 585
R10080 GND.n5034 GND.n2759 585
R10081 GND.n27 GND.n25 585
R10082 GND.n5238 GND.n27 585
R10083 GND.n7826 GND.n7825 585
R10084 GND.n7825 GND.n7824 585
R10085 GND.n26 GND.n24 585
R10086 GND.n5244 GND.n26 585
R10087 GND.n5006 GND.n5005 585
R10088 GND.n5006 GND.n2747 585
R10089 GND.n5008 GND.n5007 585
R10090 GND.n5007 GND.n2738 585
R10091 GND.n5009 GND.n2737 585
R10092 GND.n5253 GND.n2737 585
R10093 GND.n5010 GND.n2732 585
R10094 GND.n5257 GND.n2732 585
R10095 GND.n5012 GND.n5011 585
R10096 GND.n5013 GND.n5012 585
R10097 GND.n2816 GND.n2723 585
R10098 GND.n5263 GND.n2723 585
R10099 GND.n4997 GND.n4996 585
R10100 GND.n4996 GND.n4995 585
R10101 GND.n2818 GND.n2712 585
R10102 GND.n5269 GND.n2712 585
R10103 GND.n4987 GND.n4986 585
R10104 GND.n4988 GND.n4987 585
R10105 GND.n2820 GND.n2702 585
R10106 GND.n5275 GND.n2702 585
R10107 GND.n4982 GND.n4981 585
R10108 GND.n4981 GND.n4980 585
R10109 GND.n2822 GND.n2691 585
R10110 GND.n5281 GND.n2691 585
R10111 GND.n4972 GND.n4971 585
R10112 GND.n4973 GND.n4972 585
R10113 GND.n2824 GND.n2681 585
R10114 GND.n5287 GND.n2681 585
R10115 GND.n4967 GND.n4966 585
R10116 GND.n4966 GND.n4965 585
R10117 GND.n2826 GND.n2670 585
R10118 GND.n5293 GND.n2670 585
R10119 GND.n4957 GND.n4956 585
R10120 GND.n4958 GND.n4957 585
R10121 GND.n2828 GND.n2660 585
R10122 GND.n5299 GND.n2660 585
R10123 GND.n4952 GND.n4951 585
R10124 GND.n4951 GND.n4950 585
R10125 GND.n2830 GND.n2649 585
R10126 GND.n5305 GND.n2649 585
R10127 GND.n4942 GND.n4941 585
R10128 GND.n4943 GND.n4942 585
R10129 GND.n2892 GND.n2638 585
R10130 GND.n5311 GND.n2638 585
R10131 GND.n4937 GND.n4936 585
R10132 GND.n4936 GND.n4935 585
R10133 GND.n4920 GND.n2620 585
R10134 GND.n5317 GND.n2620 585
R10135 GND.n4919 GND.n4918 585
R10136 GND.n4918 GND.n2618 585
R10137 GND.n4917 GND.n2894 585
R10138 GND.n4917 GND.n2608 585
R10139 GND.n4913 GND.n2607 585
R10140 GND.n5325 GND.n2607 585
R10141 GND.n4912 GND.n2596 585
R10142 GND.n5332 GND.n2596 585
R10143 GND.n4911 GND.n4910 585
R10144 GND.n4910 GND.n4909 585
R10145 GND.n5526 GND.n2372 585
R10146 GND.n5477 GND.n2372 585
R10147 GND.n5528 GND.n5527 585
R10148 GND.n5529 GND.n5528 585
R10149 GND.n2360 GND.n2359 585
R10150 GND.n4792 GND.n2360 585
R10151 GND.n5539 GND.n5538 585
R10152 GND.n5538 GND.n5537 585
R10153 GND.n5540 GND.n2354 585
R10154 GND.n2941 GND.n2354 585
R10155 GND.n5542 GND.n5541 585
R10156 GND.n5543 GND.n5542 585
R10157 GND.n2340 GND.n2339 585
R10158 GND.n4752 GND.n2340 585
R10159 GND.n5553 GND.n5552 585
R10160 GND.n5552 GND.n5551 585
R10161 GND.n5554 GND.n2334 585
R10162 GND.n4738 GND.n2334 585
R10163 GND.n5556 GND.n5555 585
R10164 GND.n5557 GND.n5556 585
R10165 GND.n2320 GND.n2319 585
R10166 GND.n4702 GND.n2320 585
R10167 GND.n5567 GND.n5566 585
R10168 GND.n5566 GND.n5565 585
R10169 GND.n5568 GND.n2309 585
R10170 GND.n4694 GND.n2309 585
R10171 GND.n5570 GND.n5569 585
R10172 GND.n5571 GND.n5570 585
R10173 GND.n2310 GND.n2308 585
R10174 GND.n4685 GND.n2308 585
R10175 GND.n2313 GND.n2312 585
R10176 GND.n2312 GND.n2291 585
R10177 GND.n2279 GND.n2278 585
R10178 GND.n2289 GND.n2279 585
R10179 GND.n5588 GND.n5587 585
R10180 GND.n5587 GND.n5586 585
R10181 GND.n5589 GND.n2273 585
R10182 GND.n4674 GND.n2273 585
R10183 GND.n5591 GND.n5590 585
R10184 GND.n5592 GND.n5591 585
R10185 GND.n2274 GND.n2272 585
R10186 GND.n4640 GND.n2272 585
R10187 GND.n4623 GND.n4621 585
R10188 GND.n4623 GND.n4622 585
R10189 GND.n4625 GND.n4624 585
R10190 GND.n4624 GND.n2259 585
R10191 GND.n4626 GND.n4597 585
R10192 GND.n4597 GND.n2253 585
R10193 GND.n4628 GND.n4627 585
R10194 GND.n4629 GND.n4628 585
R10195 GND.n4598 GND.n4596 585
R10196 GND.n4596 GND.n4595 585
R10197 GND.n4613 GND.n4612 585
R10198 GND.n4612 GND.n2236 585
R10199 GND.n4611 GND.n4600 585
R10200 GND.n4611 GND.n2229 585
R10201 GND.n4610 GND.n4609 585
R10202 GND.n4610 GND.n2222 585
R10203 GND.n4602 GND.n4601 585
R10204 GND.n4601 GND.n2220 585
R10205 GND.n4605 GND.n4604 585
R10206 GND.n4604 GND.n2206 585
R10207 GND.n2195 GND.n2194 585
R10208 GND.n4561 GND.n2195 585
R10209 GND.n5642 GND.n5641 585
R10210 GND.n5641 GND.n5640 585
R10211 GND.n5643 GND.n2189 585
R10212 GND.n4544 GND.n2189 585
R10213 GND.n5645 GND.n5644 585
R10214 GND.n5646 GND.n5645 585
R10215 GND.n2190 GND.n2188 585
R10216 GND.n4534 GND.n2188 585
R10217 GND.n4500 GND.n4499 585
R10218 GND.n4500 GND.n2177 585
R10219 GND.n4502 GND.n4501 585
R10220 GND.n4501 GND.n2175 585
R10221 GND.n4503 GND.n3004 585
R10222 GND.n3004 GND.n2169 585
R10223 GND.n4505 GND.n4504 585
R10224 GND.n4506 GND.n4505 585
R10225 GND.n3005 GND.n3003 585
R10226 GND.n4480 GND.n3003 585
R10227 GND.n4491 GND.n4490 585
R10228 GND.n4490 GND.n2157 585
R10229 GND.n4489 GND.n3007 585
R10230 GND.n4489 GND.n2151 585
R10231 GND.n4488 GND.n3009 585
R10232 GND.n4488 GND.n4487 585
R10233 GND.n4454 GND.n3008 585
R10234 GND.n4366 GND.n3008 585
R10235 GND.n4456 GND.n4455 585
R10236 GND.n4455 GND.n2140 585
R10237 GND.n4457 GND.n3019 585
R10238 GND.n3019 GND.n2134 585
R10239 GND.n4459 GND.n4458 585
R10240 GND.n4460 GND.n4459 585
R10241 GND.n3020 GND.n3018 585
R10242 GND.n4377 GND.n3018 585
R10243 GND.n4446 GND.n4445 585
R10244 GND.n4445 GND.n2122 585
R10245 GND.n4444 GND.n3022 585
R10246 GND.n4444 GND.n2116 585
R10247 GND.n4443 GND.n3037 585
R10248 GND.n4443 GND.n4442 585
R10249 GND.n3024 GND.n3023 585
R10250 GND.n4392 GND.n3023 585
R10251 GND.n3033 GND.n3032 585
R10252 GND.n3032 GND.n2104 585
R10253 GND.n3031 GND.n3026 585
R10254 GND.n3031 GND.n2098 585
R10255 GND.n3030 GND.n3029 585
R10256 GND.n3030 GND.n2096 585
R10257 GND.n2079 GND.n2078 585
R10258 GND.n3053 GND.n2079 585
R10259 GND.n5726 GND.n5725 585
R10260 GND.n5725 GND.n5724 585
R10261 GND.n5727 GND.n2065 585
R10262 GND.n4417 GND.n2065 585
R10263 GND.n5729 GND.n5728 585
R10264 GND.n5730 GND.n5729 585
R10265 GND.n2066 GND.n2064 585
R10266 GND.n2064 GND.n2054 585
R10267 GND.n2072 GND.n2071 585
R10268 GND.n2071 GND.n2052 585
R10269 GND.n2070 GND.n2069 585
R10270 GND.n2070 GND.n2037 585
R10271 GND.n2026 GND.n2025 585
R10272 GND.n2036 GND.n2026 585
R10273 GND.n5753 GND.n5752 585
R10274 GND.n5752 GND.n5751 585
R10275 GND.n5754 GND.n2020 585
R10276 GND.n4320 GND.n2020 585
R10277 GND.n5756 GND.n5755 585
R10278 GND.n5757 GND.n5756 585
R10279 GND.n2021 GND.n2019 585
R10280 GND.n4297 GND.n2019 585
R10281 GND.n3068 GND.n3067 585
R10282 GND.n3069 GND.n3068 585
R10283 GND.n1980 GND.n1979 585
R10284 GND.n1989 GND.n1980 585
R10285 GND.n5774 GND.n5773 585
R10286 GND.n5773 GND.n5772 585
R10287 GND.n5775 GND.n1974 585
R10288 GND.n4272 GND.n1974 585
R10289 GND.n5777 GND.n5776 585
R10290 GND.n5778 GND.n5777 585
R10291 GND.n1975 GND.n1973 585
R10292 GND.n4259 GND.n1973 585
R10293 GND.n4255 GND.n4254 585
R10294 GND.n4256 GND.n4255 585
R10295 GND.n4250 GND.n3081 585
R10296 GND.n4249 GND.n4248 585
R10297 GND.n4246 GND.n3083 585
R10298 GND.n4246 GND.n1896 585
R10299 GND.n4245 GND.n4244 585
R10300 GND.n4243 GND.n4242 585
R10301 GND.n4241 GND.n3088 585
R10302 GND.n4239 GND.n4238 585
R10303 GND.n4237 GND.n3089 585
R10304 GND.n4236 GND.n4235 585
R10305 GND.n4233 GND.n3094 585
R10306 GND.n4231 GND.n4230 585
R10307 GND.n3096 GND.n3095 585
R10308 GND.n4217 GND.n4154 585
R10309 GND.n4216 GND.n4155 585
R10310 GND.n4165 GND.n4156 585
R10311 GND.n4209 GND.n4166 585
R10312 GND.n4208 GND.n4168 585
R10313 GND.n4175 GND.n4169 585
R10314 GND.n4201 GND.n4177 585
R10315 GND.n4197 GND.n4178 585
R10316 GND.n4186 GND.n4179 585
R10317 GND.n4190 GND.n4188 585
R10318 GND.n4189 GND.n3079 585
R10319 GND.n5480 GND.n5479 585
R10320 GND.n5482 GND.n5481 585
R10321 GND.n5484 GND.n5483 585
R10322 GND.n5486 GND.n5485 585
R10323 GND.n5488 GND.n5487 585
R10324 GND.n5490 GND.n5489 585
R10325 GND.n5492 GND.n5491 585
R10326 GND.n5494 GND.n5493 585
R10327 GND.n5496 GND.n5495 585
R10328 GND.n5498 GND.n5497 585
R10329 GND.n5500 GND.n5499 585
R10330 GND.n5502 GND.n5501 585
R10331 GND.n5504 GND.n5503 585
R10332 GND.n5506 GND.n5505 585
R10333 GND.n5508 GND.n5507 585
R10334 GND.n5510 GND.n5509 585
R10335 GND.n5512 GND.n5511 585
R10336 GND.n5514 GND.n5513 585
R10337 GND.n5516 GND.n5515 585
R10338 GND.n5517 GND.n2389 585
R10339 GND.n5519 GND.n5518 585
R10340 GND.n2377 GND.n2376 585
R10341 GND.n5523 GND.n5522 585
R10342 GND.n5522 GND.n5521 585
R10343 GND.n5478 GND.n2414 585
R10344 GND.n5478 GND.n5477 585
R10345 GND.n4795 GND.n2370 585
R10346 GND.n5529 GND.n2370 585
R10347 GND.n4794 GND.n4793 585
R10348 GND.n4793 GND.n4792 585
R10349 GND.n2933 GND.n2361 585
R10350 GND.n5537 GND.n2361 585
R10351 GND.n4748 GND.n4747 585
R10352 GND.n4747 GND.n2941 585
R10353 GND.n4749 GND.n2352 585
R10354 GND.n5543 GND.n2352 585
R10355 GND.n4751 GND.n4750 585
R10356 GND.n4752 GND.n4751 585
R10357 GND.n2948 GND.n2342 585
R10358 GND.n5551 GND.n2342 585
R10359 GND.n4740 GND.n4739 585
R10360 GND.n4739 GND.n4738 585
R10361 GND.n2950 GND.n2332 585
R10362 GND.n5557 GND.n2332 585
R10363 GND.n4701 GND.n4700 585
R10364 GND.n4702 GND.n4701 585
R10365 GND.n2954 GND.n2322 585
R10366 GND.n5565 GND.n2322 585
R10367 GND.n4696 GND.n4695 585
R10368 GND.n4695 GND.n4694 585
R10369 GND.n2956 GND.n2306 585
R10370 GND.n5571 GND.n2306 585
R10371 GND.n4684 GND.n4683 585
R10372 GND.n4685 GND.n4684 585
R10373 GND.n2964 GND.n2963 585
R10374 GND.n2963 GND.n2291 585
R10375 GND.n4679 GND.n4678 585
R10376 GND.n4678 GND.n2289 585
R10377 GND.n4677 GND.n2281 585
R10378 GND.n5586 GND.n2281 585
R10379 GND.n4676 GND.n4675 585
R10380 GND.n4675 GND.n4674 585
R10381 GND.n2966 GND.n2270 585
R10382 GND.n5592 GND.n2270 585
R10383 GND.n4639 GND.n4638 585
R10384 GND.n4640 GND.n4639 585
R10385 GND.n2976 GND.n2975 585
R10386 GND.n4622 GND.n2975 585
R10387 GND.n4633 GND.n4632 585
R10388 GND.n4632 GND.n2259 585
R10389 GND.n4631 GND.n2978 585
R10390 GND.n4631 GND.n2253 585
R10391 GND.n4630 GND.n4576 585
R10392 GND.n4630 GND.n4629 585
R10393 GND.n2980 GND.n2979 585
R10394 GND.n4595 GND.n2979 585
R10395 GND.n4572 GND.n4571 585
R10396 GND.n4571 GND.n2236 585
R10397 GND.n4570 GND.n2982 585
R10398 GND.n4570 GND.n2229 585
R10399 GND.n4569 GND.n4568 585
R10400 GND.n4569 GND.n2222 585
R10401 GND.n2984 GND.n2983 585
R10402 GND.n2983 GND.n2220 585
R10403 GND.n4564 GND.n4563 585
R10404 GND.n4563 GND.n2206 585
R10405 GND.n4562 GND.n2986 585
R10406 GND.n4562 GND.n4561 585
R10407 GND.n4541 GND.n2197 585
R10408 GND.n5640 GND.n2197 585
R10409 GND.n4543 GND.n4542 585
R10410 GND.n4544 GND.n4543 585
R10411 GND.n2991 GND.n2186 585
R10412 GND.n5646 GND.n2186 585
R10413 GND.n4536 GND.n4535 585
R10414 GND.n4535 GND.n4534 585
R10415 GND.n2994 GND.n2993 585
R10416 GND.n2994 GND.n2177 585
R10417 GND.n4475 GND.n4474 585
R10418 GND.n4475 GND.n2175 585
R10419 GND.n4477 GND.n4476 585
R10420 GND.n4476 GND.n2169 585
R10421 GND.n4478 GND.n3002 585
R10422 GND.n4506 GND.n3002 585
R10423 GND.n4481 GND.n4479 585
R10424 GND.n4481 GND.n4480 585
R10425 GND.n4483 GND.n4482 585
R10426 GND.n4482 GND.n2157 585
R10427 GND.n4484 GND.n3011 585
R10428 GND.n3011 GND.n2151 585
R10429 GND.n4486 GND.n4485 585
R10430 GND.n4487 GND.n4486 585
R10431 GND.n3012 GND.n3010 585
R10432 GND.n4366 GND.n3010 585
R10433 GND.n4464 GND.n4463 585
R10434 GND.n4463 GND.n2140 585
R10435 GND.n4462 GND.n3014 585
R10436 GND.n4462 GND.n2134 585
R10437 GND.n4461 GND.n3016 585
R10438 GND.n4461 GND.n4460 585
R10439 GND.n4436 GND.n3015 585
R10440 GND.n4377 GND.n3015 585
R10441 GND.n4438 GND.n4437 585
R10442 GND.n4437 GND.n2122 585
R10443 GND.n4439 GND.n3040 585
R10444 GND.n3040 GND.n2116 585
R10445 GND.n4441 GND.n4440 585
R10446 GND.n4442 GND.n4441 585
R10447 GND.n3041 GND.n3039 585
R10448 GND.n4392 GND.n3039 585
R10449 GND.n4428 GND.n4427 585
R10450 GND.n4427 GND.n2104 585
R10451 GND.n4426 GND.n3043 585
R10452 GND.n4426 GND.n2098 585
R10453 GND.n4425 GND.n4424 585
R10454 GND.n4425 GND.n2096 585
R10455 GND.n3045 GND.n3044 585
R10456 GND.n3053 GND.n3044 585
R10457 GND.n4420 GND.n2081 585
R10458 GND.n5724 GND.n2081 585
R10459 GND.n4419 GND.n4418 585
R10460 GND.n4418 GND.n4417 585
R10461 GND.n3047 GND.n2062 585
R10462 GND.n5730 GND.n2062 585
R10463 GND.n4311 GND.n4306 585
R10464 GND.n4306 GND.n2054 585
R10465 GND.n4313 GND.n4312 585
R10466 GND.n4313 GND.n2052 585
R10467 GND.n4314 GND.n4305 585
R10468 GND.n4314 GND.n2037 585
R10469 GND.n4316 GND.n4315 585
R10470 GND.n4315 GND.n2036 585
R10471 GND.n4317 GND.n2028 585
R10472 GND.n5751 GND.n2028 585
R10473 GND.n4319 GND.n4318 585
R10474 GND.n4320 GND.n4319 585
R10475 GND.n3059 GND.n2017 585
R10476 GND.n5757 GND.n2017 585
R10477 GND.n4299 GND.n4298 585
R10478 GND.n4298 GND.n4297 585
R10479 GND.n3062 GND.n3061 585
R10480 GND.n3069 GND.n3062 585
R10481 GND.n4268 GND.n4267 585
R10482 GND.n4267 GND.n1989 585
R10483 GND.n4269 GND.n1982 585
R10484 GND.n5772 GND.n1982 585
R10485 GND.n4271 GND.n4270 585
R10486 GND.n4272 GND.n4271 585
R10487 GND.n3077 GND.n1971 585
R10488 GND.n5778 GND.n1971 585
R10489 GND.n4261 GND.n4260 585
R10490 GND.n4260 GND.n4259 585
R10491 GND.n4257 GND.n3078 585
R10492 GND.n4257 GND.n4256 585
R10493 GND.n2496 GND.n2465 585
R10494 GND.n2465 GND.n2443 585
R10495 GND.n2431 GND.n2430 585
R10496 GND.n2433 GND.n2431 585
R10497 GND.n5460 GND.n5459 585
R10498 GND.n5459 GND.n5458 585
R10499 GND.n5461 GND.n2429 585
R10500 GND.n2429 GND.n2428 585
R10501 GND.n5463 GND.n5462 585
R10502 GND.n5464 GND.n5463 585
R10503 GND.n2419 GND.n2418 585
R10504 GND.n2426 GND.n2419 585
R10505 GND.n5472 GND.n5471 585
R10506 GND.n5471 GND.n5470 585
R10507 GND.n5473 GND.n2417 585
R10508 GND.n2420 GND.n2417 585
R10509 GND.n5475 GND.n5474 585
R10510 GND.n5476 GND.n5475 585
R10511 GND.n2368 GND.n2367 585
R10512 GND.n2371 GND.n2368 585
R10513 GND.n5532 GND.n5531 585
R10514 GND.n5531 GND.n5530 585
R10515 GND.n5533 GND.n2365 585
R10516 GND.n4791 GND.n2365 585
R10517 GND.n5535 GND.n5534 585
R10518 GND.n5536 GND.n5535 585
R10519 GND.n2366 GND.n2364 585
R10520 GND.n4768 GND.n2364 585
R10521 GND.n2944 GND.n2943 585
R10522 GND.n2945 GND.n2944 585
R10523 GND.n2349 GND.n2348 585
R10524 GND.n2353 GND.n2349 585
R10525 GND.n5546 GND.n5545 585
R10526 GND.n5545 GND.n5544 585
R10527 GND.n5547 GND.n2346 585
R10528 GND.n4753 GND.n2346 585
R10529 GND.n5549 GND.n5548 585
R10530 GND.n5550 GND.n5549 585
R10531 GND.n2347 GND.n2345 585
R10532 GND.n2345 GND.n2341 585
R10533 GND.n4712 GND.n4711 585
R10534 GND.n4713 GND.n4712 585
R10535 GND.n2329 GND.n2328 585
R10536 GND.n2333 GND.n2329 585
R10537 GND.n5560 GND.n5559 585
R10538 GND.n5559 GND.n5558 585
R10539 GND.n5561 GND.n2326 585
R10540 GND.n4703 GND.n2326 585
R10541 GND.n5563 GND.n5562 585
R10542 GND.n5564 GND.n5563 585
R10543 GND.n2327 GND.n2325 585
R10544 GND.n2325 GND.n2321 585
R10545 GND.n4692 GND.n4691 585
R10546 GND.n4693 GND.n4692 585
R10547 GND.n4690 GND.n2959 585
R10548 GND.n2959 GND.n2307 585
R10549 GND.n4689 GND.n4688 585
R10550 GND.n4688 GND.n2305 585
R10551 GND.n4687 GND.n2960 585
R10552 GND.n4687 GND.n4686 585
R10553 GND.n2288 GND.n2287 585
R10554 GND.n4663 GND.n2288 585
R10555 GND.n5581 GND.n5580 585
R10556 GND.n5580 GND.n5579 585
R10557 GND.n5582 GND.n2285 585
R10558 GND.n4667 GND.n2285 585
R10559 GND.n5584 GND.n5583 585
R10560 GND.n5585 GND.n5584 585
R10561 GND.n2286 GND.n2284 585
R10562 GND.n4673 GND.n2284 585
R10563 GND.n4643 GND.n4642 585
R10564 GND.n4643 GND.n2969 585
R10565 GND.n4645 GND.n4644 585
R10566 GND.n4644 GND.n2271 585
R10567 GND.n4646 GND.n4641 585
R10568 GND.n4641 GND.n2269 585
R10569 GND.n4648 GND.n4647 585
R10570 GND.n4649 GND.n4648 585
R10571 GND.n2258 GND.n2257 585
R10572 GND.n2261 GND.n2258 585
R10573 GND.n5602 GND.n5601 585
R10574 GND.n5601 GND.n5600 585
R10575 GND.n5603 GND.n2255 585
R10576 GND.n4584 GND.n2255 585
R10577 GND.n5605 GND.n5604 585
R10578 GND.n5606 GND.n5605 585
R10579 GND.n2256 GND.n2254 585
R10580 GND.n2254 GND.n2251 585
R10581 GND.n4592 GND.n4591 585
R10582 GND.n4593 GND.n4592 585
R10583 GND.n2235 GND.n2234 585
R10584 GND.n2238 GND.n2235 585
R10585 GND.n5616 GND.n5615 585
R10586 GND.n5615 GND.n5614 585
R10587 GND.n5617 GND.n2232 585
R10588 GND.n2239 GND.n2232 585
R10589 GND.n5619 GND.n5618 585
R10590 GND.n5620 GND.n5619 585
R10591 GND.n2233 GND.n2231 585
R10592 GND.n2231 GND.n2230 585
R10593 GND.n4549 GND.n2221 585
R10594 GND.n5626 GND.n2221 585
R10595 GND.n4551 GND.n4550 585
R10596 GND.n4552 GND.n4551 585
R10597 GND.n2204 GND.n2203 585
R10598 GND.n4554 GND.n2204 585
R10599 GND.n5635 GND.n5634 585
R10600 GND.n5634 GND.n5633 585
R10601 GND.n5636 GND.n2201 585
R10602 GND.n4560 GND.n2201 585
R10603 GND.n5638 GND.n5637 585
R10604 GND.n5639 GND.n5638 585
R10605 GND.n2202 GND.n2200 585
R10606 GND.n4545 GND.n2200 585
R10607 GND.n4527 GND.n4526 585
R10608 GND.n4527 GND.n2990 585
R10609 GND.n4529 GND.n4528 585
R10610 GND.n4528 GND.n2187 585
R10611 GND.n4530 GND.n4525 585
R10612 GND.n4525 GND.n2185 585
R10613 GND.n4532 GND.n4531 585
R10614 GND.n4533 GND.n4532 585
R10615 GND.n2174 GND.n2173 585
R10616 GND.n2996 GND.n2174 585
R10617 GND.n5656 GND.n5655 585
R10618 GND.n5655 GND.n5654 585
R10619 GND.n5657 GND.n2171 585
R10620 GND.n4515 GND.n2171 585
R10621 GND.n5659 GND.n5658 585
R10622 GND.n5660 GND.n5659 585
R10623 GND.n2172 GND.n2170 585
R10624 GND.n2170 GND.n2167 585
R10625 GND.n4508 GND.n4507 585
R10626 GND.n4509 GND.n4508 585
R10627 GND.n2156 GND.n2155 585
R10628 GND.n2159 GND.n2156 585
R10629 GND.n5670 GND.n5669 585
R10630 GND.n5669 GND.n5668 585
R10631 GND.n5671 GND.n2153 585
R10632 GND.n4355 GND.n2153 585
R10633 GND.n5673 GND.n5672 585
R10634 GND.n5674 GND.n5673 585
R10635 GND.n2154 GND.n2152 585
R10636 GND.n2152 GND.n2149 585
R10637 GND.n4363 GND.n4362 585
R10638 GND.n4364 GND.n4363 585
R10639 GND.n2139 GND.n2138 585
R10640 GND.n4367 GND.n2139 585
R10641 GND.n5684 GND.n5683 585
R10642 GND.n5683 GND.n5682 585
R10643 GND.n5685 GND.n2136 585
R10644 GND.n4371 GND.n2136 585
R10645 GND.n5687 GND.n5686 585
R10646 GND.n5688 GND.n5687 585
R10647 GND.n2137 GND.n2135 585
R10648 GND.n2135 GND.n2132 585
R10649 GND.n4379 GND.n4378 585
R10650 GND.n4380 GND.n4379 585
R10651 GND.n2121 GND.n2120 585
R10652 GND.n2124 GND.n2121 585
R10653 GND.n5698 GND.n5697 585
R10654 GND.n5697 GND.n5696 585
R10655 GND.n5699 GND.n2118 585
R10656 GND.n4386 GND.n2118 585
R10657 GND.n5701 GND.n5700 585
R10658 GND.n5702 GND.n5701 585
R10659 GND.n2119 GND.n2117 585
R10660 GND.n2117 GND.n2114 585
R10661 GND.n4394 GND.n4393 585
R10662 GND.n4395 GND.n4394 585
R10663 GND.n2103 GND.n2102 585
R10664 GND.n2106 GND.n2103 585
R10665 GND.n5712 GND.n5711 585
R10666 GND.n5711 GND.n5710 585
R10667 GND.n5713 GND.n2100 585
R10668 GND.n4401 GND.n2100 585
R10669 GND.n5715 GND.n5714 585
R10670 GND.n5716 GND.n5715 585
R10671 GND.n2101 GND.n2099 585
R10672 GND.n4407 GND.n2099 585
R10673 GND.n4410 GND.n3052 585
R10674 GND.n4410 GND.n4409 585
R10675 GND.n4412 GND.n4411 585
R10676 GND.n4411 GND.n2082 585
R10677 GND.n4413 GND.n3051 585
R10678 GND.n3051 GND.n2080 585
R10679 GND.n4415 GND.n4414 585
R10680 GND.n4416 GND.n4415 585
R10681 GND.n2059 GND.n2058 585
R10682 GND.n3048 GND.n2059 585
R10683 GND.n5733 GND.n5732 585
R10684 GND.n5732 GND.n5731 585
R10685 GND.n5734 GND.n2056 585
R10686 GND.n4337 GND.n2056 585
R10687 GND.n5736 GND.n5735 585
R10688 GND.n5737 GND.n5736 585
R10689 GND.n2057 GND.n2055 585
R10690 GND.n4333 GND.n2055 585
R10691 GND.n2035 GND.n2034 585
R10692 GND.n4331 GND.n2035 585
R10693 GND.n5746 GND.n5745 585
R10694 GND.n5745 GND.n5744 585
R10695 GND.n5747 GND.n2032 585
R10696 GND.n4325 GND.n2032 585
R10697 GND.n5749 GND.n5748 585
R10698 GND.n5750 GND.n5749 585
R10699 GND.n2033 GND.n2031 585
R10700 GND.n4321 GND.n2031 585
R10701 GND.n4290 GND.n4289 585
R10702 GND.n4290 GND.n3058 585
R10703 GND.n4292 GND.n4291 585
R10704 GND.n4291 GND.n2018 585
R10705 GND.n4293 GND.n4288 585
R10706 GND.n4288 GND.n2016 585
R10707 GND.n4295 GND.n4294 585
R10708 GND.n4296 GND.n4295 585
R10709 GND.n1988 GND.n1987 585
R10710 GND.n3070 GND.n1988 585
R10711 GND.n5767 GND.n5766 585
R10712 GND.n5766 GND.n5765 585
R10713 GND.n5768 GND.n1985 585
R10714 GND.n4278 GND.n1985 585
R10715 GND.n5770 GND.n5769 585
R10716 GND.n5771 GND.n5770 585
R10717 GND.n1986 GND.n1984 585
R10718 GND.n4273 GND.n1984 585
R10719 GND.n1968 GND.n1967 585
R10720 GND.n3076 GND.n1968 585
R10721 GND.n5781 GND.n5780 585
R10722 GND.n5780 GND.n5779 585
R10723 GND.n5782 GND.n1966 585
R10724 GND.n4258 GND.n1966 585
R10725 GND.n5784 GND.n5783 585
R10726 GND.n5785 GND.n5784 585
R10727 GND.n1901 GND.n1900 585
R10728 GND.n3080 GND.n1901 585
R10729 GND.n5792 GND.n5791 585
R10730 GND.n5791 GND.t153 585
R10731 GND.n5793 GND.n1898 585
R10732 GND.n1903 GND.n1898 585
R10733 GND.n5795 GND.n5794 585
R10734 GND.n5796 GND.n5795 585
R10735 GND.n1899 GND.n1897 585
R10736 GND.n1897 GND.n1894 585
R10737 GND.n1956 GND.n1955 585
R10738 GND.n1957 GND.n1956 585
R10739 GND.n1882 GND.n1881 585
R10740 GND.n1885 GND.n1882 585
R10741 GND.n5806 GND.n5805 585
R10742 GND.n5805 GND.n5804 585
R10743 GND.n5807 GND.n1850 585
R10744 GND.n1883 GND.n1850 585
R10745 GND.n5845 GND.n5844 585
R10746 GND.n5843 GND.n1849 585
R10747 GND.n5842 GND.n1848 585
R10748 GND.n5847 GND.n1848 585
R10749 GND.n5841 GND.n5840 585
R10750 GND.n5839 GND.n5838 585
R10751 GND.n5837 GND.n5836 585
R10752 GND.n5835 GND.n5834 585
R10753 GND.n5833 GND.n5832 585
R10754 GND.n5831 GND.n5830 585
R10755 GND.n5829 GND.n5828 585
R10756 GND.n5827 GND.n5826 585
R10757 GND.n5825 GND.n5824 585
R10758 GND.n5823 GND.n5822 585
R10759 GND.n5821 GND.n5820 585
R10760 GND.n5819 GND.n5818 585
R10761 GND.n5817 GND.n5816 585
R10762 GND.n5814 GND.n5813 585
R10763 GND.n5812 GND.n5811 585
R10764 GND.n1826 GND.n1825 585
R10765 GND.n5850 GND.n5849 585
R10766 GND.n1910 GND.n1823 585
R10767 GND.n1912 GND.n1911 585
R10768 GND.n1914 GND.n1913 585
R10769 GND.n1916 GND.n1915 585
R10770 GND.n1919 GND.n1918 585
R10771 GND.n1921 GND.n1920 585
R10772 GND.n1923 GND.n1922 585
R10773 GND.n1925 GND.n1924 585
R10774 GND.n1927 GND.n1926 585
R10775 GND.n1929 GND.n1928 585
R10776 GND.n1931 GND.n1930 585
R10777 GND.n1933 GND.n1932 585
R10778 GND.n1935 GND.n1934 585
R10779 GND.n1937 GND.n1936 585
R10780 GND.n1939 GND.n1938 585
R10781 GND.n1941 GND.n1940 585
R10782 GND.n1943 GND.n1942 585
R10783 GND.n1945 GND.n1944 585
R10784 GND.n1947 GND.n1946 585
R10785 GND.n1948 GND.n1846 585
R10786 GND.n5847 GND.n1846 585
R10787 GND.n2509 GND.n2508 585
R10788 GND.n2511 GND.n2510 585
R10789 GND.n2513 GND.n2512 585
R10790 GND.n2515 GND.n2514 585
R10791 GND.n2517 GND.n2516 585
R10792 GND.n2519 GND.n2518 585
R10793 GND.n2521 GND.n2520 585
R10794 GND.n2523 GND.n2522 585
R10795 GND.n2525 GND.n2524 585
R10796 GND.n2527 GND.n2526 585
R10797 GND.n2529 GND.n2528 585
R10798 GND.n2531 GND.n2530 585
R10799 GND.n2533 GND.n2532 585
R10800 GND.n2535 GND.n2534 585
R10801 GND.n2537 GND.n2536 585
R10802 GND.n2539 GND.n2538 585
R10803 GND.n2541 GND.n2540 585
R10804 GND.n2543 GND.n2542 585
R10805 GND.n2545 GND.n2544 585
R10806 GND.n2547 GND.n2546 585
R10807 GND.n5450 GND.n2444 585
R10808 GND.n5411 GND.n5410 585
R10809 GND.n5413 GND.n5412 585
R10810 GND.n5415 GND.n5414 585
R10811 GND.n5417 GND.n5416 585
R10812 GND.n5420 GND.n5419 585
R10813 GND.n5422 GND.n5421 585
R10814 GND.n5424 GND.n5423 585
R10815 GND.n5426 GND.n5425 585
R10816 GND.n5428 GND.n5427 585
R10817 GND.n5430 GND.n5429 585
R10818 GND.n5432 GND.n5431 585
R10819 GND.n5434 GND.n5433 585
R10820 GND.n5436 GND.n5435 585
R10821 GND.n5438 GND.n5437 585
R10822 GND.n5440 GND.n5439 585
R10823 GND.n5442 GND.n5441 585
R10824 GND.n5444 GND.n5443 585
R10825 GND.n5446 GND.n5445 585
R10826 GND.n5447 GND.n2466 585
R10827 GND.n5449 GND.n5448 585
R10828 GND.n5450 GND.n5449 585
R10829 GND.n2507 GND.n2503 585
R10830 GND.n2507 GND.n2443 585
R10831 GND.n2506 GND.n2505 585
R10832 GND.n2506 GND.n2433 585
R10833 GND.n2504 GND.n2432 585
R10834 GND.n5458 GND.n2432 585
R10835 GND.n2425 GND.n2424 585
R10836 GND.n2428 GND.n2425 585
R10837 GND.n5466 GND.n5465 585
R10838 GND.n5465 GND.n5464 585
R10839 GND.n5467 GND.n2422 585
R10840 GND.n2426 GND.n2422 585
R10841 GND.n5469 GND.n5468 585
R10842 GND.n5470 GND.n5469 585
R10843 GND.n2423 GND.n2421 585
R10844 GND.n2421 GND.n2420 585
R10845 GND.n4760 GND.n2416 585
R10846 GND.n5476 GND.n2416 585
R10847 GND.n4762 GND.n4761 585
R10848 GND.n4761 GND.n2371 585
R10849 GND.n4763 GND.n2369 585
R10850 GND.n5530 GND.n2369 585
R10851 GND.n4764 GND.n2934 585
R10852 GND.n4791 GND.n2934 585
R10853 GND.n4765 GND.n2362 585
R10854 GND.n5536 GND.n2362 585
R10855 GND.n4767 GND.n4766 585
R10856 GND.n4768 GND.n4767 585
R10857 GND.n4759 GND.n2946 585
R10858 GND.n2946 GND.n2945 585
R10859 GND.n4758 GND.n4757 585
R10860 GND.n4757 GND.n2353 585
R10861 GND.n4756 GND.n2351 585
R10862 GND.n5544 GND.n2351 585
R10863 GND.n4755 GND.n4754 585
R10864 GND.n4754 GND.n4753 585
R10865 GND.n2947 GND.n2343 585
R10866 GND.n5550 GND.n2343 585
R10867 GND.n4708 GND.n2952 585
R10868 GND.n2952 GND.n2341 585
R10869 GND.n4710 GND.n4709 585
R10870 GND.n4713 GND.n4710 585
R10871 GND.n4707 GND.n2951 585
R10872 GND.n2951 GND.n2333 585
R10873 GND.n4706 GND.n2331 585
R10874 GND.n5558 GND.n2331 585
R10875 GND.n4705 GND.n4704 585
R10876 GND.n4704 GND.n4703 585
R10877 GND.n2953 GND.n2323 585
R10878 GND.n5564 GND.n2323 585
R10879 GND.n4656 GND.n4655 585
R10880 GND.n4655 GND.n2321 585
R10881 GND.n4657 GND.n2958 585
R10882 GND.n4693 GND.n2958 585
R10883 GND.n4659 GND.n4658 585
R10884 GND.n4659 GND.n2307 585
R10885 GND.n4661 GND.n4660 585
R10886 GND.n4660 GND.n2305 585
R10887 GND.n4662 GND.n2962 585
R10888 GND.n4686 GND.n2962 585
R10889 GND.n4665 GND.n4664 585
R10890 GND.n4664 GND.n4663 585
R10891 GND.n4666 GND.n2290 585
R10892 GND.n5579 GND.n2290 585
R10893 GND.n4669 GND.n4668 585
R10894 GND.n4668 GND.n4667 585
R10895 GND.n4670 GND.n2282 585
R10896 GND.n5585 GND.n2282 585
R10897 GND.n4672 GND.n4671 585
R10898 GND.n4673 GND.n4672 585
R10899 GND.n4654 GND.n2970 585
R10900 GND.n2970 GND.n2969 585
R10901 GND.n4653 GND.n4652 585
R10902 GND.n4652 GND.n2271 585
R10903 GND.n4651 GND.n2971 585
R10904 GND.n4651 GND.n2269 585
R10905 GND.n4650 GND.n2973 585
R10906 GND.n4650 GND.n4649 585
R10907 GND.n4581 GND.n2972 585
R10908 GND.n2972 GND.n2261 585
R10909 GND.n4582 GND.n2260 585
R10910 GND.n5600 GND.n2260 585
R10911 GND.n4586 GND.n4585 585
R10912 GND.n4585 GND.n4584 585
R10913 GND.n4587 GND.n2252 585
R10914 GND.n5606 GND.n2252 585
R10915 GND.n4588 GND.n4578 585
R10916 GND.n4578 GND.n2251 585
R10917 GND.n4590 GND.n4589 585
R10918 GND.n4593 GND.n4590 585
R10919 GND.n4580 GND.n4577 585
R10920 GND.n4577 GND.n2238 585
R10921 GND.n4579 GND.n2237 585
R10922 GND.n5614 GND.n2237 585
R10923 GND.n2227 GND.n2226 585
R10924 GND.n2239 GND.n2227 585
R10925 GND.n5622 GND.n5621 585
R10926 GND.n5621 GND.n5620 585
R10927 GND.n5623 GND.n2224 585
R10928 GND.n2230 GND.n2224 585
R10929 GND.n5625 GND.n5624 585
R10930 GND.n5626 GND.n5625 585
R10931 GND.n2225 GND.n2223 585
R10932 GND.n4552 GND.n2223 585
R10933 GND.n4556 GND.n4555 585
R10934 GND.n4555 GND.n4554 585
R10935 GND.n4557 GND.n2205 585
R10936 GND.n5633 GND.n2205 585
R10937 GND.n4559 GND.n4558 585
R10938 GND.n4560 GND.n4559 585
R10939 GND.n4548 GND.n2198 585
R10940 GND.n5639 GND.n2198 585
R10941 GND.n4547 GND.n4546 585
R10942 GND.n4546 GND.n4545 585
R10943 GND.n2988 GND.n2987 585
R10944 GND.n2990 GND.n2988 585
R10945 GND.n4521 GND.n4520 585
R10946 GND.n4520 GND.n2187 585
R10947 GND.n4522 GND.n2998 585
R10948 GND.n2998 GND.n2185 585
R10949 GND.n4524 GND.n4523 585
R10950 GND.n4533 GND.n4524 585
R10951 GND.n4519 GND.n2997 585
R10952 GND.n2997 GND.n2996 585
R10953 GND.n4518 GND.n2176 585
R10954 GND.n5654 GND.n2176 585
R10955 GND.n4517 GND.n4516 585
R10956 GND.n4516 GND.n4515 585
R10957 GND.n4513 GND.n2168 585
R10958 GND.n5660 GND.n2168 585
R10959 GND.n4512 GND.n4511 585
R10960 GND.n4511 GND.n2167 585
R10961 GND.n4510 GND.n2999 585
R10962 GND.n4510 GND.n4509 585
R10963 GND.n4352 GND.n3000 585
R10964 GND.n3000 GND.n2159 585
R10965 GND.n4353 GND.n2158 585
R10966 GND.n5668 GND.n2158 585
R10967 GND.n4357 GND.n4356 585
R10968 GND.n4356 GND.n4355 585
R10969 GND.n4358 GND.n2150 585
R10970 GND.n5674 GND.n2150 585
R10971 GND.n4360 GND.n4359 585
R10972 GND.n4360 GND.n2149 585
R10973 GND.n4361 GND.n4351 585
R10974 GND.n4364 GND.n4361 585
R10975 GND.n4369 GND.n4368 585
R10976 GND.n4368 GND.n4367 585
R10977 GND.n4370 GND.n2141 585
R10978 GND.n5682 GND.n2141 585
R10979 GND.n4373 GND.n4372 585
R10980 GND.n4372 GND.n4371 585
R10981 GND.n4374 GND.n2133 585
R10982 GND.n5688 GND.n2133 585
R10983 GND.n4376 GND.n4375 585
R10984 GND.n4376 GND.n2132 585
R10985 GND.n4381 GND.n4350 585
R10986 GND.n4381 GND.n4380 585
R10987 GND.n4383 GND.n4382 585
R10988 GND.n4382 GND.n2124 585
R10989 GND.n4384 GND.n2123 585
R10990 GND.n5696 GND.n2123 585
R10991 GND.n4388 GND.n4387 585
R10992 GND.n4387 GND.n4386 585
R10993 GND.n4389 GND.n2115 585
R10994 GND.n5702 GND.n2115 585
R10995 GND.n4391 GND.n4390 585
R10996 GND.n4391 GND.n2114 585
R10997 GND.n4396 GND.n4349 585
R10998 GND.n4396 GND.n4395 585
R10999 GND.n4398 GND.n4397 585
R11000 GND.n4397 GND.n2106 585
R11001 GND.n4399 GND.n2105 585
R11002 GND.n5710 GND.n2105 585
R11003 GND.n4403 GND.n4402 585
R11004 GND.n4402 GND.n4401 585
R11005 GND.n4404 GND.n2097 585
R11006 GND.n5716 GND.n2097 585
R11007 GND.n4406 GND.n4405 585
R11008 GND.n4407 GND.n4406 585
R11009 GND.n4348 GND.n3054 585
R11010 GND.n4409 GND.n3054 585
R11011 GND.n4347 GND.n4346 585
R11012 GND.n4346 GND.n2082 585
R11013 GND.n4345 GND.n4344 585
R11014 GND.n4345 GND.n2080 585
R11015 GND.n4343 GND.n3049 585
R11016 GND.n4416 GND.n3049 585
R11017 GND.n4342 GND.n4341 585
R11018 GND.n4341 GND.n3048 585
R11019 GND.n4340 GND.n2061 585
R11020 GND.n5731 GND.n2061 585
R11021 GND.n4339 GND.n4338 585
R11022 GND.n4338 GND.n4337 585
R11023 GND.n4336 GND.n2053 585
R11024 GND.n5737 GND.n2053 585
R11025 GND.n4335 GND.n4334 585
R11026 GND.n4334 GND.n4333 585
R11027 GND.n4330 GND.n4329 585
R11028 GND.n4331 GND.n4330 585
R11029 GND.n4328 GND.n2038 585
R11030 GND.n5744 GND.n2038 585
R11031 GND.n4327 GND.n4326 585
R11032 GND.n4326 GND.n4325 585
R11033 GND.n4324 GND.n2029 585
R11034 GND.n5750 GND.n2029 585
R11035 GND.n4323 GND.n4322 585
R11036 GND.n4322 GND.n4321 585
R11037 GND.n3056 GND.n3055 585
R11038 GND.n3058 GND.n3056 585
R11039 GND.n4284 GND.n4283 585
R11040 GND.n4283 GND.n2018 585
R11041 GND.n4285 GND.n3072 585
R11042 GND.n3072 GND.n2016 585
R11043 GND.n4287 GND.n4286 585
R11044 GND.n4296 GND.n4287 585
R11045 GND.n4282 GND.n3071 585
R11046 GND.n3071 GND.n3070 585
R11047 GND.n4281 GND.n1990 585
R11048 GND.n5765 GND.n1990 585
R11049 GND.n4280 GND.n4279 585
R11050 GND.n4279 GND.n4278 585
R11051 GND.n4276 GND.n1983 585
R11052 GND.n5771 GND.n1983 585
R11053 GND.n4275 GND.n4274 585
R11054 GND.n4274 GND.n4273 585
R11055 GND.n3075 GND.n3074 585
R11056 GND.n3076 GND.n3075 585
R11057 GND.n3073 GND.n1970 585
R11058 GND.n5779 GND.n1970 585
R11059 GND.n1964 GND.n1963 585
R11060 GND.n4258 GND.n1964 585
R11061 GND.n5787 GND.n5786 585
R11062 GND.n5786 GND.n5785 585
R11063 GND.n5788 GND.n1906 585
R11064 GND.n3080 GND.n1906 585
R11065 GND.n5790 GND.n5789 585
R11066 GND.t153 GND.n5790 585
R11067 GND.n1962 GND.n1905 585
R11068 GND.n1905 GND.n1903 585
R11069 GND.n1961 GND.n1895 585
R11070 GND.n5796 GND.n1895 585
R11071 GND.n1960 GND.n1959 585
R11072 GND.n1959 GND.n1894 585
R11073 GND.n1958 GND.n1907 585
R11074 GND.n1958 GND.n1957 585
R11075 GND.n1953 GND.n1952 585
R11076 GND.n1953 GND.n1885 585
R11077 GND.n1951 GND.n1884 585
R11078 GND.n5804 GND.n1884 585
R11079 GND.n1950 GND.n1949 585
R11080 GND.n1949 GND.n1883 585
R11081 GND.n4146 GND.n1782 585
R11082 GND.n4223 GND.n1782 585
R11083 GND.n4148 GND.n4147 585
R11084 GND.n4149 GND.n4148 585
R11085 GND.n3192 GND.n3191 585
R11086 GND.n4133 GND.n3191 585
R11087 GND.n4142 GND.n4141 585
R11088 GND.n4141 GND.n4140 585
R11089 GND.n3195 GND.n3194 585
R11090 GND.n4130 GND.n3195 585
R11091 GND.n4081 GND.n3218 585
R11092 GND.n3218 GND.n3206 585
R11093 GND.n4083 GND.n4082 585
R11094 GND.n4084 GND.n4083 585
R11095 GND.n3219 GND.n3217 585
R11096 GND.n3217 GND.n3213 585
R11097 GND.n4076 GND.n4075 585
R11098 GND.n4075 GND.n4074 585
R11099 GND.n3222 GND.n3221 585
R11100 GND.n4059 GND.n3222 585
R11101 GND.n4044 GND.n3248 585
R11102 GND.n3248 GND.n3235 585
R11103 GND.n4046 GND.n4045 585
R11104 GND.n4047 GND.n4046 585
R11105 GND.n3249 GND.n3247 585
R11106 GND.n3247 GND.n3243 585
R11107 GND.n4039 GND.n4038 585
R11108 GND.n4038 GND.n4037 585
R11109 GND.n3252 GND.n3251 585
R11110 GND.n4022 GND.n3252 585
R11111 GND.n4007 GND.n3277 585
R11112 GND.n3277 GND.n3264 585
R11113 GND.n4009 GND.n4008 585
R11114 GND.n4010 GND.n4009 585
R11115 GND.n3278 GND.n3276 585
R11116 GND.n3276 GND.n3271 585
R11117 GND.n4002 GND.n4001 585
R11118 GND.n4001 GND.n4000 585
R11119 GND.n3281 GND.n3280 585
R11120 GND.n3985 GND.n3281 585
R11121 GND.n3970 GND.n3306 585
R11122 GND.n3306 GND.n3294 585
R11123 GND.n3972 GND.n3971 585
R11124 GND.n3973 GND.n3972 585
R11125 GND.n3307 GND.n3305 585
R11126 GND.n3305 GND.n3301 585
R11127 GND.n3965 GND.n3964 585
R11128 GND.n3964 GND.n3963 585
R11129 GND.n3310 GND.n3309 585
R11130 GND.n3948 GND.n3310 585
R11131 GND.n3911 GND.n3910 585
R11132 GND.n3912 GND.n3911 585
R11133 GND.n3909 GND.n3854 585
R11134 GND.n3859 GND.n3854 585
R11135 GND.n3907 GND.n3906 585
R11136 GND.n3906 GND.n3905 585
R11137 GND.n3856 GND.n3855 585
R11138 GND.n3902 GND.n3856 585
R11139 GND.n3885 GND.n3881 585
R11140 GND.n3881 GND.n3863 585
R11141 GND.n3887 GND.n3886 585
R11142 GND.n3888 GND.n3887 585
R11143 GND.n3882 GND.n3880 585
R11144 GND.n3880 GND.n3879 585
R11145 GND.n3344 GND.n3343 585
R11146 GND.n3869 GND.n3344 585
R11147 GND.n3932 GND.n3931 585
R11148 GND.n3931 GND.n3930 585
R11149 GND.n3934 GND.n3340 585
R11150 GND.n3836 GND.n3340 585
R11151 GND.n3936 GND.n3935 585
R11152 GND.n3937 GND.n3936 585
R11153 GND.n3341 GND.n3339 585
R11154 GND.n3830 GND.n3339 585
R11155 GND.n3825 GND.n3824 585
R11156 GND.n3826 GND.n3825 585
R11157 GND.n3363 GND.n3362 585
R11158 GND.n3371 GND.n3362 585
R11159 GND.n3819 GND.n3818 585
R11160 GND.n3818 GND.n3817 585
R11161 GND.n3366 GND.n3365 585
R11162 GND.n3809 GND.n3366 585
R11163 GND.n3787 GND.n3392 585
R11164 GND.n3392 GND.n3380 585
R11165 GND.n3789 GND.n3788 585
R11166 GND.n3790 GND.n3789 585
R11167 GND.n3393 GND.n3391 585
R11168 GND.n3391 GND.n3387 585
R11169 GND.n3782 GND.n3781 585
R11170 GND.n3781 GND.n3780 585
R11171 GND.n3396 GND.n3395 585
R11172 GND.n3765 GND.n3396 585
R11173 GND.n3750 GND.n3422 585
R11174 GND.n3422 GND.n3409 585
R11175 GND.n3752 GND.n3751 585
R11176 GND.n3753 GND.n3752 585
R11177 GND.n3423 GND.n3421 585
R11178 GND.n3421 GND.n3417 585
R11179 GND.n3745 GND.n3744 585
R11180 GND.n3744 GND.n3743 585
R11181 GND.n3426 GND.n3425 585
R11182 GND.n3728 GND.n3426 585
R11183 GND.n3713 GND.n3451 585
R11184 GND.n3451 GND.n3438 585
R11185 GND.n3715 GND.n3714 585
R11186 GND.n3716 GND.n3715 585
R11187 GND.n3452 GND.n3450 585
R11188 GND.n3450 GND.n3445 585
R11189 GND.n3708 GND.n3707 585
R11190 GND.n3707 GND.n3706 585
R11191 GND.n3455 GND.n3454 585
R11192 GND.n3691 GND.n3455 585
R11193 GND.n3676 GND.n3480 585
R11194 GND.n3480 GND.n3468 585
R11195 GND.n3678 GND.n3677 585
R11196 GND.n3679 GND.n3678 585
R11197 GND.n3481 GND.n3479 585
R11198 GND.n3479 GND.n3475 585
R11199 GND.n3671 GND.n3670 585
R11200 GND.n3670 GND.n3669 585
R11201 GND.n3527 GND.n3483 585
R11202 GND.n3529 GND.n3528 585
R11203 GND.n3531 GND.n3530 585
R11204 GND.n3535 GND.n3525 585
R11205 GND.n3537 GND.n3536 585
R11206 GND.n3539 GND.n3538 585
R11207 GND.n3541 GND.n3540 585
R11208 GND.n3545 GND.n3523 585
R11209 GND.n3547 GND.n3546 585
R11210 GND.n3549 GND.n3548 585
R11211 GND.n3551 GND.n3550 585
R11212 GND.n3555 GND.n3554 585
R11213 GND.n3557 GND.n3556 585
R11214 GND.n3560 GND.n3559 585
R11215 GND.n3558 GND.n3517 585
R11216 GND.n3565 GND.n3564 585
R11217 GND.n3567 GND.n3566 585
R11218 GND.n3570 GND.n3569 585
R11219 GND.n3568 GND.n3515 585
R11220 GND.n3575 GND.n3574 585
R11221 GND.n3577 GND.n3576 585
R11222 GND.n3580 GND.n3579 585
R11223 GND.n3578 GND.n3513 585
R11224 GND.n3585 GND.n3584 585
R11225 GND.n3587 GND.n3586 585
R11226 GND.n3589 GND.n3588 585
R11227 GND.n3591 GND.n3590 585
R11228 GND.n3595 GND.n3507 585
R11229 GND.n3597 GND.n3596 585
R11230 GND.n3599 GND.n3598 585
R11231 GND.n3601 GND.n3600 585
R11232 GND.n3605 GND.n3505 585
R11233 GND.n3607 GND.n3606 585
R11234 GND.n3609 GND.n3608 585
R11235 GND.n3611 GND.n3610 585
R11236 GND.n3502 GND.n3501 585
R11237 GND.n3617 GND.n3503 585
R11238 GND.n3619 GND.n3618 585
R11239 GND.n3621 GND.n3620 585
R11240 GND.n3625 GND.n3499 585
R11241 GND.n3627 GND.n3626 585
R11242 GND.n3629 GND.n3628 585
R11243 GND.n3631 GND.n3630 585
R11244 GND.n3635 GND.n3497 585
R11245 GND.n3637 GND.n3636 585
R11246 GND.n3639 GND.n3638 585
R11247 GND.n3641 GND.n3640 585
R11248 GND.n3645 GND.n3495 585
R11249 GND.n3647 GND.n3646 585
R11250 GND.n3651 GND.n3648 585
R11251 GND.n3652 GND.n1640 585
R11252 GND.n6004 GND.n1640 585
R11253 GND.n3185 GND.n3184 585
R11254 GND.n3183 GND.n3182 585
R11255 GND.n3181 GND.n3104 585
R11256 GND.n3177 GND.n3176 585
R11257 GND.n3175 GND.n3174 585
R11258 GND.n3173 GND.n3110 585
R11259 GND.n3109 GND.n3108 585
R11260 GND.n3169 GND.n3168 585
R11261 GND.n3167 GND.n3166 585
R11262 GND.n3165 GND.n3114 585
R11263 GND.n3113 GND.n3112 585
R11264 GND.n3161 GND.n3160 585
R11265 GND.n3159 GND.n3158 585
R11266 GND.n3157 GND.n3120 585
R11267 GND.n3119 GND.n3118 585
R11268 GND.n3153 GND.n3152 585
R11269 GND.n3151 GND.n3150 585
R11270 GND.n3149 GND.n3124 585
R11271 GND.n3123 GND.n3122 585
R11272 GND.n3145 GND.n3144 585
R11273 GND.n3143 GND.n3142 585
R11274 GND.n3141 GND.n3128 585
R11275 GND.n3127 GND.n3126 585
R11276 GND.n3137 GND.n3136 585
R11277 GND.n3135 GND.n3134 585
R11278 GND.n3133 GND.n3131 585
R11279 GND.n3130 GND.n1819 585
R11280 GND.n1817 GND.n1816 585
R11281 GND.n5856 GND.n1815 585
R11282 GND.n5857 GND.n1814 585
R11283 GND.n5858 GND.n1813 585
R11284 GND.n1811 GND.n1810 585
R11285 GND.n5862 GND.n1809 585
R11286 GND.n5863 GND.n1808 585
R11287 GND.n5864 GND.n1807 585
R11288 GND.n1805 GND.n1804 585
R11289 GND.n5868 GND.n1803 585
R11290 GND.n5869 GND.n1802 585
R11291 GND.n5871 GND.n1799 585
R11292 GND.n1797 GND.n1796 585
R11293 GND.n5875 GND.n1795 585
R11294 GND.n5876 GND.n1794 585
R11295 GND.n5877 GND.n1793 585
R11296 GND.n1791 GND.n1790 585
R11297 GND.n5881 GND.n1789 585
R11298 GND.n5882 GND.n1788 585
R11299 GND.n5883 GND.n1787 585
R11300 GND.n1784 GND.n1783 585
R11301 GND.n5888 GND.n5887 585
R11302 GND.n5889 GND.n5888 585
R11303 GND.n4225 GND.n4224 585
R11304 GND.n4224 GND.n4223 585
R11305 GND.n3103 GND.n3102 585
R11306 GND.n4149 GND.n3103 585
R11307 GND.n4135 GND.n4134 585
R11308 GND.n4134 GND.n4133 585
R11309 GND.n4136 GND.n3197 585
R11310 GND.n4140 GND.n3197 585
R11311 GND.n4132 GND.n4131 585
R11312 GND.n4131 GND.n4130 585
R11313 GND.n3205 GND.n3204 585
R11314 GND.n3206 GND.n3205 585
R11315 GND.n4068 GND.n3214 585
R11316 GND.n4084 GND.n3214 585
R11317 GND.n4069 GND.n4062 585
R11318 GND.n4062 GND.n3213 585
R11319 GND.n4070 GND.n3224 585
R11320 GND.n4074 GND.n3224 585
R11321 GND.n4061 GND.n4060 585
R11322 GND.n4060 GND.n4059 585
R11323 GND.n3234 GND.n3233 585
R11324 GND.n3235 GND.n3234 585
R11325 GND.n4031 GND.n3244 585
R11326 GND.n4047 GND.n3244 585
R11327 GND.n4032 GND.n4025 585
R11328 GND.n4025 GND.n3243 585
R11329 GND.n4033 GND.n3254 585
R11330 GND.n4037 GND.n3254 585
R11331 GND.n4024 GND.n4023 585
R11332 GND.n4023 GND.n4022 585
R11333 GND.n3263 GND.n3262 585
R11334 GND.n3264 GND.n3263 585
R11335 GND.n3994 GND.n3272 585
R11336 GND.n4010 GND.n3272 585
R11337 GND.n3995 GND.n3988 585
R11338 GND.n3988 GND.n3271 585
R11339 GND.n3996 GND.n3283 585
R11340 GND.n4000 GND.n3283 585
R11341 GND.n3987 GND.n3986 585
R11342 GND.n3986 GND.n3985 585
R11343 GND.n3292 GND.n3291 585
R11344 GND.n3294 GND.n3292 585
R11345 GND.n3957 GND.n3302 585
R11346 GND.n3973 GND.n3302 585
R11347 GND.n3958 GND.n3951 585
R11348 GND.n3951 GND.n3301 585
R11349 GND.n3959 GND.n3311 585
R11350 GND.n3963 GND.n3311 585
R11351 GND.n3950 GND.n3949 585
R11352 GND.n3949 GND.n3948 585
R11353 GND.n3320 GND.n3319 585
R11354 GND.n3912 GND.n3320 585
R11355 GND.n3858 GND.n3849 585
R11356 GND.n3859 GND.n3858 585
R11357 GND.n3918 GND.n3848 585
R11358 GND.n3905 GND.n3848 585
R11359 GND.n3919 GND.n3847 585
R11360 GND.n3902 GND.n3847 585
R11361 GND.n3920 GND.n3846 585
R11362 GND.n3863 GND.n3846 585
R11363 GND.n3866 GND.n3841 585
R11364 GND.n3888 GND.n3866 585
R11365 GND.n3924 GND.n3840 585
R11366 GND.n3879 GND.n3840 585
R11367 GND.n3925 GND.n3839 585
R11368 GND.n3869 GND.n3839 585
R11369 GND.n3926 GND.n3346 585
R11370 GND.n3930 GND.n3346 585
R11371 GND.n3838 GND.n3837 585
R11372 GND.n3837 GND.n3836 585
R11373 GND.n3835 GND.n3336 585
R11374 GND.n3937 GND.n3336 585
R11375 GND.n3828 GND.n3354 585
R11376 GND.n3830 GND.n3828 585
R11377 GND.n3827 GND.n3360 585
R11378 GND.n3827 GND.n3826 585
R11379 GND.n3812 GND.n3359 585
R11380 GND.n3371 GND.n3359 585
R11381 GND.n3813 GND.n3368 585
R11382 GND.n3817 GND.n3368 585
R11383 GND.n3811 GND.n3810 585
R11384 GND.n3810 GND.n3809 585
R11385 GND.n3379 GND.n3378 585
R11386 GND.n3380 GND.n3379 585
R11387 GND.n3774 GND.n3388 585
R11388 GND.n3790 GND.n3388 585
R11389 GND.n3775 GND.n3768 585
R11390 GND.n3768 GND.n3387 585
R11391 GND.n3776 GND.n3398 585
R11392 GND.n3780 GND.n3398 585
R11393 GND.n3767 GND.n3766 585
R11394 GND.n3766 GND.n3765 585
R11395 GND.n3408 GND.n3407 585
R11396 GND.n3409 GND.n3408 585
R11397 GND.n3737 GND.n3418 585
R11398 GND.n3753 GND.n3418 585
R11399 GND.n3738 GND.n3731 585
R11400 GND.n3731 GND.n3417 585
R11401 GND.n3739 GND.n3428 585
R11402 GND.n3743 GND.n3428 585
R11403 GND.n3730 GND.n3729 585
R11404 GND.n3729 GND.n3728 585
R11405 GND.n3437 GND.n3436 585
R11406 GND.n3438 GND.n3437 585
R11407 GND.n3700 GND.n3446 585
R11408 GND.n3716 GND.n3446 585
R11409 GND.n3701 GND.n3694 585
R11410 GND.n3694 GND.n3445 585
R11411 GND.n3702 GND.n3457 585
R11412 GND.n3706 GND.n3457 585
R11413 GND.n3693 GND.n3692 585
R11414 GND.n3692 GND.n3691 585
R11415 GND.n3466 GND.n3465 585
R11416 GND.n3468 GND.n3466 585
R11417 GND.n3662 GND.n3476 585
R11418 GND.n3679 GND.n3476 585
R11419 GND.n3493 GND.n3492 585
R11420 GND.n3492 GND.n3475 585
R11421 GND.n3667 GND.n3666 585
R11422 GND.n3669 GND.n3667 585
R11423 GND.n171 GND.n170 585
R11424 GND.n7738 GND.n171 585
R11425 GND.n7747 GND.n7746 585
R11426 GND.n7746 GND.n7745 585
R11427 GND.n7748 GND.n165 585
R11428 GND.n5161 GND.n165 585
R11429 GND.n7750 GND.n7749 585
R11430 GND.n7751 GND.n7750 585
R11431 GND.n150 GND.n149 585
R11432 GND.n5167 GND.n150 585
R11433 GND.n7759 GND.n7758 585
R11434 GND.n7758 GND.n7757 585
R11435 GND.n7760 GND.n144 585
R11436 GND.n5173 GND.n144 585
R11437 GND.n7762 GND.n7761 585
R11438 GND.n7763 GND.n7762 585
R11439 GND.n130 GND.n129 585
R11440 GND.n5179 GND.n130 585
R11441 GND.n7771 GND.n7770 585
R11442 GND.n7770 GND.n7769 585
R11443 GND.n7772 GND.n124 585
R11444 GND.n5098 GND.n124 585
R11445 GND.n7774 GND.n7773 585
R11446 GND.n7775 GND.n7774 585
R11447 GND.n109 GND.n108 585
R11448 GND.n5089 GND.n109 585
R11449 GND.n7783 GND.n7782 585
R11450 GND.n7782 GND.n7781 585
R11451 GND.n7784 GND.n103 585
R11452 GND.n5083 GND.n103 585
R11453 GND.n7786 GND.n7785 585
R11454 GND.n7787 GND.n7786 585
R11455 GND.n88 GND.n87 585
R11456 GND.n5075 GND.n88 585
R11457 GND.n7795 GND.n7794 585
R11458 GND.n7794 GND.n7793 585
R11459 GND.n7796 GND.n82 585
R11460 GND.n5069 GND.n82 585
R11461 GND.n7798 GND.n7797 585
R11462 GND.n7799 GND.n7798 585
R11463 GND.n67 GND.n66 585
R11464 GND.n5061 GND.n67 585
R11465 GND.n7807 GND.n7806 585
R11466 GND.n7806 GND.n7805 585
R11467 GND.n7808 GND.n62 585
R11468 GND.n5055 GND.n62 585
R11469 GND.n7810 GND.n7809 585
R11470 GND.n7811 GND.n7810 585
R11471 GND.n46 GND.n44 585
R11472 GND.n5047 GND.n46 585
R11473 GND.n7819 GND.n7818 585
R11474 GND.n7818 GND.n7817 585
R11475 GND.n45 GND.n43 585
R11476 GND.n5040 GND.n45 585
R11477 GND.n2758 GND.n2757 585
R11478 GND.n2759 GND.n2758 585
R11479 GND.n35 GND.n33 585
R11480 GND.n5238 GND.n33 585
R11481 GND.n7823 GND.n7822 585
R11482 GND.n7824 GND.n7823 585
R11483 GND.n34 GND.n32 585
R11484 GND.n5244 GND.n32 585
R11485 GND.n2746 GND.n2745 585
R11486 GND.n2747 GND.n2746 585
R11487 GND.n2734 GND.n41 585
R11488 GND.n2738 GND.n2734 585
R11489 GND.n5254 GND.n2735 585
R11490 GND.n5254 GND.n5253 585
R11491 GND.n5256 GND.n5255 585
R11492 GND.n5257 GND.n5256 585
R11493 GND.n2720 GND.n2719 585
R11494 GND.n5013 GND.n2720 585
R11495 GND.n5265 GND.n5264 585
R11496 GND.n5264 GND.n5263 585
R11497 GND.n5266 GND.n2714 585
R11498 GND.n4995 GND.n2714 585
R11499 GND.n5268 GND.n5267 585
R11500 GND.n5269 GND.n5268 585
R11501 GND.n2699 GND.n2698 585
R11502 GND.n4988 GND.n2699 585
R11503 GND.n5277 GND.n5276 585
R11504 GND.n5276 GND.n5275 585
R11505 GND.n5278 GND.n2693 585
R11506 GND.n4980 GND.n2693 585
R11507 GND.n5280 GND.n5279 585
R11508 GND.n5281 GND.n5280 585
R11509 GND.n2678 GND.n2677 585
R11510 GND.n4973 GND.n2678 585
R11511 GND.n5289 GND.n5288 585
R11512 GND.n5288 GND.n5287 585
R11513 GND.n5290 GND.n2672 585
R11514 GND.n4965 GND.n2672 585
R11515 GND.n5292 GND.n5291 585
R11516 GND.n5293 GND.n5292 585
R11517 GND.n2657 GND.n2656 585
R11518 GND.n4958 GND.n2657 585
R11519 GND.n5301 GND.n5300 585
R11520 GND.n5300 GND.n5299 585
R11521 GND.n5302 GND.n2651 585
R11522 GND.n4950 GND.n2651 585
R11523 GND.n5304 GND.n5303 585
R11524 GND.n5305 GND.n5304 585
R11525 GND.n2635 GND.n2634 585
R11526 GND.n4943 GND.n2635 585
R11527 GND.n5313 GND.n5312 585
R11528 GND.n5312 GND.n5311 585
R11529 GND.n5314 GND.n2624 585
R11530 GND.n4935 GND.n2624 585
R11531 GND.n5316 GND.n5315 585
R11532 GND.n5317 GND.n5316 585
R11533 GND.n2625 GND.n2623 585
R11534 GND.n2623 GND.n2618 585
R11535 GND.n2628 GND.n2627 585
R11536 GND.n2627 GND.n2608 585
R11537 GND.n2593 GND.n2592 585
R11538 GND.n5325 GND.n2593 585
R11539 GND.n5334 GND.n5333 585
R11540 GND.n5333 GND.n5332 585
R11541 GND.n5335 GND.n2590 585
R11542 GND.n4909 GND.n2590 585
R11543 GND.n5402 GND.n5401 585
R11544 GND.n5400 GND.n2589 585
R11545 GND.n5399 GND.n2588 585
R11546 GND.n5404 GND.n2588 585
R11547 GND.n5398 GND.n5397 585
R11548 GND.n5396 GND.n5395 585
R11549 GND.n5394 GND.n5393 585
R11550 GND.n5392 GND.n5391 585
R11551 GND.n5390 GND.n5389 585
R11552 GND.n5388 GND.n5387 585
R11553 GND.n5386 GND.n5385 585
R11554 GND.n5384 GND.n5383 585
R11555 GND.n5382 GND.n5381 585
R11556 GND.n5380 GND.n5379 585
R11557 GND.n5378 GND.n5377 585
R11558 GND.n5376 GND.n5375 585
R11559 GND.n5374 GND.n5373 585
R11560 GND.n5372 GND.n5371 585
R11561 GND.n5370 GND.n5369 585
R11562 GND.n5368 GND.n5367 585
R11563 GND.n5366 GND.n5365 585
R11564 GND.n5364 GND.n5363 585
R11565 GND.n5362 GND.n2549 585
R11566 GND.n5407 GND.n5406 585
R11567 GND.n2556 GND.n2555 585
R11568 GND.n4843 GND.n4842 585
R11569 GND.n4845 GND.n4844 585
R11570 GND.n4848 GND.n4847 585
R11571 GND.n4846 GND.n4838 585
R11572 GND.n4853 GND.n4852 585
R11573 GND.n4855 GND.n4854 585
R11574 GND.n4858 GND.n4857 585
R11575 GND.n4856 GND.n4836 585
R11576 GND.n4863 GND.n4862 585
R11577 GND.n4865 GND.n4864 585
R11578 GND.n4870 GND.n4867 585
R11579 GND.n4866 GND.n4834 585
R11580 GND.n4875 GND.n4874 585
R11581 GND.n4877 GND.n4876 585
R11582 GND.n4880 GND.n4879 585
R11583 GND.n4878 GND.n4832 585
R11584 GND.n4885 GND.n4884 585
R11585 GND.n4887 GND.n4886 585
R11586 GND.n4890 GND.n4889 585
R11587 GND.n4888 GND.n4830 585
R11588 GND.n4895 GND.n4894 585
R11589 GND.n4897 GND.n4896 585
R11590 GND.n4900 GND.n4899 585
R11591 GND.n4898 GND.n4828 585
R11592 GND.n4907 GND.n4906 585
R11593 GND.n270 GND.n180 585
R11594 GND.n276 GND.n275 585
R11595 GND.n278 GND.n277 585
R11596 GND.n280 GND.n279 585
R11597 GND.n282 GND.n281 585
R11598 GND.n284 GND.n283 585
R11599 GND.n286 GND.n285 585
R11600 GND.n288 GND.n287 585
R11601 GND.n290 GND.n289 585
R11602 GND.n292 GND.n291 585
R11603 GND.n294 GND.n293 585
R11604 GND.n296 GND.n295 585
R11605 GND.n298 GND.n297 585
R11606 GND.n258 GND.n255 585
R11607 GND.n302 GND.n259 585
R11608 GND.n304 GND.n303 585
R11609 GND.n306 GND.n305 585
R11610 GND.n308 GND.n307 585
R11611 GND.n310 GND.n309 585
R11612 GND.n312 GND.n311 585
R11613 GND.n314 GND.n313 585
R11614 GND.n316 GND.n315 585
R11615 GND.n318 GND.n317 585
R11616 GND.n320 GND.n319 585
R11617 GND.n322 GND.n321 585
R11618 GND.n324 GND.n323 585
R11619 GND.n326 GND.n325 585
R11620 GND.n331 GND.n330 585
R11621 GND.n333 GND.n332 585
R11622 GND.n335 GND.n334 585
R11623 GND.n337 GND.n336 585
R11624 GND.n339 GND.n338 585
R11625 GND.n341 GND.n340 585
R11626 GND.n343 GND.n342 585
R11627 GND.n345 GND.n344 585
R11628 GND.n347 GND.n346 585
R11629 GND.n349 GND.n348 585
R11630 GND.n351 GND.n350 585
R11631 GND.n353 GND.n352 585
R11632 GND.n355 GND.n354 585
R11633 GND.n357 GND.n356 585
R11634 GND.n359 GND.n358 585
R11635 GND.n361 GND.n360 585
R11636 GND.n363 GND.n362 585
R11637 GND.n365 GND.n364 585
R11638 GND.n367 GND.n366 585
R11639 GND.n369 GND.n368 585
R11640 GND.n372 GND.n371 585
R11641 GND.n370 GND.n219 585
R11642 GND.n376 GND.n216 585
R11643 GND.n378 GND.n377 585
R11644 GND.n379 GND.n378 585
R11645 GND.n7740 GND.n7739 585
R11646 GND.n7739 GND.n7738 585
R11647 GND.n179 GND.n173 585
R11648 GND.n7745 GND.n173 585
R11649 GND.n5160 GND.n5159 585
R11650 GND.n5161 GND.n5160 585
R11651 GND.n5105 GND.n162 585
R11652 GND.n7751 GND.n162 585
R11653 GND.n5169 GND.n5168 585
R11654 GND.n5168 GND.n5167 585
R11655 GND.n5170 GND.n152 585
R11656 GND.n7757 GND.n152 585
R11657 GND.n5172 GND.n5171 585
R11658 GND.n5173 GND.n5172 585
R11659 GND.n5103 GND.n141 585
R11660 GND.n7763 GND.n141 585
R11661 GND.n5102 GND.n2787 585
R11662 GND.n5179 GND.n2787 585
R11663 GND.n5101 GND.n132 585
R11664 GND.n7769 GND.n132 585
R11665 GND.n5100 GND.n5099 585
R11666 GND.n5099 GND.n5098 585
R11667 GND.n2793 GND.n121 585
R11668 GND.n7775 GND.n121 585
R11669 GND.n5088 GND.n5087 585
R11670 GND.n5089 GND.n5088 585
R11671 GND.n5086 GND.n111 585
R11672 GND.n7781 GND.n111 585
R11673 GND.n5085 GND.n5084 585
R11674 GND.n5084 GND.n5083 585
R11675 GND.n2798 GND.n100 585
R11676 GND.n7787 GND.n100 585
R11677 GND.n5074 GND.n5073 585
R11678 GND.n5075 GND.n5074 585
R11679 GND.n5072 GND.n90 585
R11680 GND.n7793 GND.n90 585
R11681 GND.n5071 GND.n5070 585
R11682 GND.n5070 GND.n5069 585
R11683 GND.n2803 GND.n79 585
R11684 GND.n7799 GND.n79 585
R11685 GND.n5060 GND.n5059 585
R11686 GND.n5061 GND.n5060 585
R11687 GND.n5058 GND.n69 585
R11688 GND.n7805 GND.n69 585
R11689 GND.n5057 GND.n5056 585
R11690 GND.n5056 GND.n5055 585
R11691 GND.n2808 GND.n59 585
R11692 GND.n7811 GND.n59 585
R11693 GND.n5045 GND.n5044 585
R11694 GND.n5047 GND.n5045 585
R11695 GND.n5043 GND.n48 585
R11696 GND.n7817 GND.n48 585
R11697 GND.n5042 GND.n5041 585
R11698 GND.n5041 GND.n5040 585
R11699 GND.n5032 GND.n5029 585
R11700 GND.n5032 GND.n2759 585
R11701 GND.n5028 GND.n2756 585
R11702 GND.n5238 GND.n2756 585
R11703 GND.n5027 GND.n29 585
R11704 GND.n7824 GND.n29 585
R11705 GND.n5026 GND.n2748 585
R11706 GND.n5244 GND.n2748 585
R11707 GND.n5025 GND.n5024 585
R11708 GND.n5024 GND.n2747 585
R11709 GND.n5023 GND.n2813 585
R11710 GND.n5023 GND.n2738 585
R11711 GND.n5017 GND.n2736 585
R11712 GND.n5253 GND.n2736 585
R11713 GND.n5016 GND.n2731 585
R11714 GND.n5257 GND.n2731 585
R11715 GND.n5015 GND.n5014 585
R11716 GND.n5014 GND.n5013 585
R11717 GND.n2814 GND.n2722 585
R11718 GND.n5263 GND.n2722 585
R11719 GND.n4994 GND.n4993 585
R11720 GND.n4995 GND.n4994 585
R11721 GND.n4991 GND.n2711 585
R11722 GND.n5269 GND.n2711 585
R11723 GND.n4990 GND.n4989 585
R11724 GND.n4989 GND.n4988 585
R11725 GND.n2819 GND.n2701 585
R11726 GND.n5275 GND.n2701 585
R11727 GND.n4979 GND.n4978 585
R11728 GND.n4980 GND.n4979 585
R11729 GND.n4976 GND.n2690 585
R11730 GND.n5281 GND.n2690 585
R11731 GND.n4975 GND.n4974 585
R11732 GND.n4974 GND.n4973 585
R11733 GND.n2823 GND.n2680 585
R11734 GND.n5287 GND.n2680 585
R11735 GND.n4964 GND.n4963 585
R11736 GND.n4965 GND.n4964 585
R11737 GND.n4961 GND.n2669 585
R11738 GND.n5293 GND.n2669 585
R11739 GND.n4960 GND.n4959 585
R11740 GND.n4959 GND.n4958 585
R11741 GND.n2827 GND.n2659 585
R11742 GND.n5299 GND.n2659 585
R11743 GND.n4949 GND.n4948 585
R11744 GND.n4950 GND.n4949 585
R11745 GND.n4946 GND.n2648 585
R11746 GND.n5305 GND.n2648 585
R11747 GND.n4945 GND.n4944 585
R11748 GND.n4944 GND.n4943 585
R11749 GND.n2831 GND.n2637 585
R11750 GND.n5311 GND.n2637 585
R11751 GND.n4934 GND.n4933 585
R11752 GND.n4935 GND.n4934 585
R11753 GND.n4921 GND.n2619 585
R11754 GND.n5317 GND.n2619 585
R11755 GND.n4923 GND.n4922 585
R11756 GND.n4922 GND.n2618 585
R11757 GND.n2606 GND.n2605 585
R11758 GND.n2608 GND.n2606 585
R11759 GND.n5327 GND.n5326 585
R11760 GND.n5326 GND.n5325 585
R11761 GND.n5328 GND.n2595 585
R11762 GND.n5332 GND.n2595 585
R11763 GND.n4908 GND.n2604 585
R11764 GND.n4909 GND.n4908 585
R11765 GND.n7565 GND.n7564 585
R11766 GND.n7564 GND.n7563 585
R11767 GND.n7566 GND.n541 585
R11768 GND.n541 GND.n540 585
R11769 GND.n7568 GND.n7567 585
R11770 GND.n7569 GND.n7568 585
R11771 GND.n539 GND.n538 585
R11772 GND.n7570 GND.n539 585
R11773 GND.n7573 GND.n7572 585
R11774 GND.n7572 GND.n7571 585
R11775 GND.n7574 GND.n533 585
R11776 GND.n533 GND.n532 585
R11777 GND.n7576 GND.n7575 585
R11778 GND.n7577 GND.n7576 585
R11779 GND.n531 GND.n530 585
R11780 GND.n7578 GND.n531 585
R11781 GND.n7581 GND.n7580 585
R11782 GND.n7580 GND.n7579 585
R11783 GND.n7582 GND.n525 585
R11784 GND.n525 GND.n524 585
R11785 GND.n7584 GND.n7583 585
R11786 GND.n7585 GND.n7584 585
R11787 GND.n523 GND.n522 585
R11788 GND.n7586 GND.n523 585
R11789 GND.n7589 GND.n7588 585
R11790 GND.n7588 GND.n7587 585
R11791 GND.n7590 GND.n517 585
R11792 GND.n517 GND.n516 585
R11793 GND.n7592 GND.n7591 585
R11794 GND.n7593 GND.n7592 585
R11795 GND.n515 GND.n514 585
R11796 GND.n7594 GND.n515 585
R11797 GND.n7597 GND.n7596 585
R11798 GND.n7596 GND.n7595 585
R11799 GND.n7598 GND.n509 585
R11800 GND.n509 GND.n508 585
R11801 GND.n7600 GND.n7599 585
R11802 GND.n7601 GND.n7600 585
R11803 GND.n507 GND.n506 585
R11804 GND.n7602 GND.n507 585
R11805 GND.n7605 GND.n7604 585
R11806 GND.n7604 GND.n7603 585
R11807 GND.n7606 GND.n501 585
R11808 GND.n501 GND.n500 585
R11809 GND.n7608 GND.n7607 585
R11810 GND.n7609 GND.n7608 585
R11811 GND.n499 GND.n498 585
R11812 GND.n7610 GND.n499 585
R11813 GND.n7613 GND.n7612 585
R11814 GND.n7612 GND.n7611 585
R11815 GND.n7614 GND.n493 585
R11816 GND.n493 GND.n492 585
R11817 GND.n7616 GND.n7615 585
R11818 GND.n7617 GND.n7616 585
R11819 GND.n491 GND.n490 585
R11820 GND.n7618 GND.n491 585
R11821 GND.n7621 GND.n7620 585
R11822 GND.n7620 GND.n7619 585
R11823 GND.n7622 GND.n485 585
R11824 GND.n485 GND.n484 585
R11825 GND.n7624 GND.n7623 585
R11826 GND.n7625 GND.n7624 585
R11827 GND.n483 GND.n482 585
R11828 GND.n7626 GND.n483 585
R11829 GND.n7629 GND.n7628 585
R11830 GND.n7628 GND.n7627 585
R11831 GND.n7630 GND.n477 585
R11832 GND.n477 GND.n476 585
R11833 GND.n7632 GND.n7631 585
R11834 GND.n7633 GND.n7632 585
R11835 GND.n475 GND.n474 585
R11836 GND.n7634 GND.n475 585
R11837 GND.n7637 GND.n7636 585
R11838 GND.n7636 GND.n7635 585
R11839 GND.n7638 GND.n469 585
R11840 GND.n469 GND.n468 585
R11841 GND.n7640 GND.n7639 585
R11842 GND.n7641 GND.n7640 585
R11843 GND.n467 GND.n466 585
R11844 GND.n7642 GND.n467 585
R11845 GND.n7645 GND.n7644 585
R11846 GND.n7644 GND.n7643 585
R11847 GND.n7646 GND.n461 585
R11848 GND.n461 GND.n460 585
R11849 GND.n7648 GND.n7647 585
R11850 GND.n7649 GND.n7648 585
R11851 GND.n459 GND.n458 585
R11852 GND.n7650 GND.n459 585
R11853 GND.n7653 GND.n7652 585
R11854 GND.n7652 GND.n7651 585
R11855 GND.n7654 GND.n453 585
R11856 GND.n453 GND.n452 585
R11857 GND.n7656 GND.n7655 585
R11858 GND.n7657 GND.n7656 585
R11859 GND.n451 GND.n450 585
R11860 GND.n7658 GND.n451 585
R11861 GND.n7661 GND.n7660 585
R11862 GND.n7660 GND.n7659 585
R11863 GND.n7662 GND.n445 585
R11864 GND.n445 GND.n444 585
R11865 GND.n7664 GND.n7663 585
R11866 GND.n7665 GND.n7664 585
R11867 GND.n443 GND.n442 585
R11868 GND.n7666 GND.n443 585
R11869 GND.n7669 GND.n7668 585
R11870 GND.n7668 GND.n7667 585
R11871 GND.n7670 GND.n437 585
R11872 GND.n437 GND.n436 585
R11873 GND.n7672 GND.n7671 585
R11874 GND.n7673 GND.n7672 585
R11875 GND.n435 GND.n434 585
R11876 GND.n7674 GND.n435 585
R11877 GND.n7677 GND.n7676 585
R11878 GND.n7676 GND.n7675 585
R11879 GND.n7678 GND.n429 585
R11880 GND.n429 GND.n428 585
R11881 GND.n7680 GND.n7679 585
R11882 GND.n7681 GND.n7680 585
R11883 GND.n427 GND.n426 585
R11884 GND.n7682 GND.n427 585
R11885 GND.n7685 GND.n7684 585
R11886 GND.n7684 GND.n7683 585
R11887 GND.n7686 GND.n421 585
R11888 GND.n421 GND.n420 585
R11889 GND.n7688 GND.n7687 585
R11890 GND.n7689 GND.n7688 585
R11891 GND.n419 GND.n418 585
R11892 GND.n7690 GND.n419 585
R11893 GND.n7693 GND.n7692 585
R11894 GND.n7692 GND.n7691 585
R11895 GND.n7694 GND.n413 585
R11896 GND.n413 GND.n412 585
R11897 GND.n7696 GND.n7695 585
R11898 GND.n7697 GND.n7696 585
R11899 GND.n411 GND.n410 585
R11900 GND.n7698 GND.n411 585
R11901 GND.n7701 GND.n7700 585
R11902 GND.n7700 GND.n7699 585
R11903 GND.n7702 GND.n405 585
R11904 GND.n405 GND.n404 585
R11905 GND.n7704 GND.n7703 585
R11906 GND.n7705 GND.n7704 585
R11907 GND.n403 GND.n402 585
R11908 GND.n7706 GND.n403 585
R11909 GND.n7709 GND.n7708 585
R11910 GND.n7708 GND.n7707 585
R11911 GND.n7710 GND.n397 585
R11912 GND.n397 GND.n396 585
R11913 GND.n7712 GND.n7711 585
R11914 GND.n7713 GND.n7712 585
R11915 GND.n395 GND.n394 585
R11916 GND.n7714 GND.n395 585
R11917 GND.n7717 GND.n7716 585
R11918 GND.n7716 GND.n7715 585
R11919 GND.n7718 GND.n389 585
R11920 GND.n389 GND.n388 585
R11921 GND.n7720 GND.n7719 585
R11922 GND.n7721 GND.n7720 585
R11923 GND.n387 GND.n386 585
R11924 GND.n7722 GND.n387 585
R11925 GND.n7725 GND.n7724 585
R11926 GND.n7724 GND.n7723 585
R11927 GND.n7726 GND.n381 585
R11928 GND.n381 GND.n380 585
R11929 GND.n7728 GND.n7727 585
R11930 GND.n7729 GND.n7728 585
R11931 GND.n190 GND.n189 585
R11932 GND.n7730 GND.n190 585
R11933 GND.n7733 GND.n7732 585
R11934 GND.n7732 GND.n7731 585
R11935 GND.n7734 GND.n184 585
R11936 GND.n184 GND.n182 585
R11937 GND.n7736 GND.n7735 585
R11938 GND.n7737 GND.n7736 585
R11939 GND.n185 GND.n183 585
R11940 GND.n183 GND.n175 585
R11941 GND.n5195 GND.n5194 585
R11942 GND.n5195 GND.n172 585
R11943 GND.n5197 GND.n5196 585
R11944 GND.n5196 GND.n164 585
R11945 GND.n5198 GND.n5187 585
R11946 GND.n5187 GND.n161 585
R11947 GND.n5200 GND.n5199 585
R11948 GND.n5200 GND.n154 585
R11949 GND.n5201 GND.n5186 585
R11950 GND.n5201 GND.n151 585
R11951 GND.n5203 GND.n5202 585
R11952 GND.n5202 GND.n143 585
R11953 GND.n5204 GND.n5181 585
R11954 GND.n5181 GND.n5180 585
R11955 GND.n5206 GND.n5205 585
R11956 GND.n5206 GND.n134 585
R11957 GND.n5207 GND.n2786 585
R11958 GND.n5207 GND.n131 585
R11959 GND.n5209 GND.n5208 585
R11960 GND.n5208 GND.n123 585
R11961 GND.n5210 GND.n2781 585
R11962 GND.n2781 GND.n120 585
R11963 GND.n5212 GND.n5211 585
R11964 GND.n5212 GND.n113 585
R11965 GND.n5213 GND.n2780 585
R11966 GND.n5213 GND.n110 585
R11967 GND.n5215 GND.n5214 585
R11968 GND.n5214 GND.n102 585
R11969 GND.n5216 GND.n2775 585
R11970 GND.n2775 GND.n99 585
R11971 GND.n5218 GND.n5217 585
R11972 GND.n5218 GND.n92 585
R11973 GND.n5219 GND.n2774 585
R11974 GND.n5219 GND.n89 585
R11975 GND.n5221 GND.n5220 585
R11976 GND.n5220 GND.n81 585
R11977 GND.n5222 GND.n2769 585
R11978 GND.n2769 GND.n78 585
R11979 GND.n5224 GND.n5223 585
R11980 GND.n5224 GND.n71 585
R11981 GND.n5225 GND.n2768 585
R11982 GND.n5225 GND.n68 585
R11983 GND.n5227 GND.n5226 585
R11984 GND.n5226 GND.n61 585
R11985 GND.n5228 GND.n2765 585
R11986 GND.n5046 GND.n2765 585
R11987 GND.n5230 GND.n5229 585
R11988 GND.n5230 GND.n50 585
R11989 GND.n5232 GND.n5231 585
R11990 GND.n5231 GND.n47 585
R11991 GND.n5233 GND.n2761 585
R11992 GND.n5033 GND.n2761 585
R11993 GND.n5236 GND.n5235 585
R11994 GND.n5237 GND.n5236 585
R11995 GND.n2763 GND.n2760 585
R11996 GND.n2760 GND.n30 585
R11997 GND.n2743 GND.n2742 585
R11998 GND.n2743 GND.n28 585
R11999 GND.n5247 GND.n5246 585
R12000 GND.n5246 GND.n5245 585
R12001 GND.n5249 GND.n2740 585
R12002 GND.n2744 GND.n2740 585
R12003 GND.n5251 GND.n5250 585
R12004 GND.n5252 GND.n5251 585
R12005 GND.n2863 GND.n2739 585
R12006 GND.n2739 GND.n2733 585
R12007 GND.n2864 GND.n2859 585
R12008 GND.n2859 GND.n2730 585
R12009 GND.n2866 GND.n2865 585
R12010 GND.n2866 GND.n2815 585
R12011 GND.n2867 GND.n2858 585
R12012 GND.n2867 GND.n2721 585
R12013 GND.n2869 GND.n2868 585
R12014 GND.n2868 GND.n2713 585
R12015 GND.n2870 GND.n2853 585
R12016 GND.n2853 GND.n2710 585
R12017 GND.n2872 GND.n2871 585
R12018 GND.n2872 GND.n2703 585
R12019 GND.n2873 GND.n2852 585
R12020 GND.n2873 GND.n2700 585
R12021 GND.n2875 GND.n2874 585
R12022 GND.n2874 GND.n2692 585
R12023 GND.n2876 GND.n2847 585
R12024 GND.n2847 GND.n2689 585
R12025 GND.n2878 GND.n2877 585
R12026 GND.n2878 GND.n2682 585
R12027 GND.n2879 GND.n2846 585
R12028 GND.n2879 GND.n2679 585
R12029 GND.n2881 GND.n2880 585
R12030 GND.n2880 GND.n2671 585
R12031 GND.n2882 GND.n2841 585
R12032 GND.n2841 GND.n2668 585
R12033 GND.n2884 GND.n2883 585
R12034 GND.n2884 GND.n2661 585
R12035 GND.n2885 GND.n2840 585
R12036 GND.n2885 GND.n2658 585
R12037 GND.n2887 GND.n2886 585
R12038 GND.n2886 GND.n2650 585
R12039 GND.n2888 GND.n2833 585
R12040 GND.n2833 GND.n2647 585
R12041 GND.n2890 GND.n2889 585
R12042 GND.n2891 GND.n2890 585
R12043 GND.n2834 GND.n2832 585
R12044 GND.n2832 GND.n2636 585
R12045 GND.n2616 GND.n2615 585
R12046 GND.n2621 GND.n2616 585
R12047 GND.n5320 GND.n5319 585
R12048 GND.n5319 GND.n5318 585
R12049 GND.n5321 GND.n2610 585
R12050 GND.n2617 GND.n2610 585
R12051 GND.n5323 GND.n5322 585
R12052 GND.n5324 GND.n5323 585
R12053 GND.n2611 GND.n2609 585
R12054 GND.n2609 GND.n2597 585
R12055 GND.n4822 GND.n4803 585
R12056 GND.n4803 GND.n2594 585
R12057 GND.n4824 GND.n4823 585
R12058 GND.n4825 GND.n4824 585
R12059 GND.n4804 GND.n4802 585
R12060 GND.n4802 GND.n2587 585
R12061 GND.n4816 GND.n4815 585
R12062 GND.n4815 GND.n2557 585
R12063 GND.n4814 GND.n4806 585
R12064 GND.n4814 GND.n4813 585
R12065 GND.n4810 GND.n4809 585
R12066 GND.n4812 GND.n4810 585
R12067 GND.n2442 GND.n2441 585
R12068 GND.n4811 GND.n2442 585
R12069 GND.n5453 GND.n5452 585
R12070 GND.n5452 GND.n5451 585
R12071 GND.n5454 GND.n2436 585
R12072 GND.n2443 GND.n2436 585
R12073 GND.n5456 GND.n5455 585
R12074 GND.n5457 GND.n5456 585
R12075 GND.n2437 GND.n2435 585
R12076 GND.n2435 GND.n2434 585
R12077 GND.n4782 GND.n4781 585
R12078 GND.n4782 GND.n2427 585
R12079 GND.n4783 GND.n4777 585
R12080 GND.n4783 GND.n2378 585
R12081 GND.n4786 GND.n4785 585
R12082 GND.n4785 GND.n4784 585
R12083 GND.n4787 GND.n2936 585
R12084 GND.n2936 GND.n2415 585
R12085 GND.n4789 GND.n4788 585
R12086 GND.n4790 GND.n4789 585
R12087 GND.n2937 GND.n2935 585
R12088 GND.n2935 GND.n2363 585
R12089 GND.n4771 GND.n4770 585
R12090 GND.n4770 GND.n4769 585
R12091 GND.n2940 GND.n2939 585
R12092 GND.n2942 GND.n2940 585
R12093 GND.n4733 GND.n4732 585
R12094 GND.n4732 GND.n2350 585
R12095 GND.n4734 GND.n4716 585
R12096 GND.n4716 GND.n2344 585
R12097 GND.n4736 GND.n4735 585
R12098 GND.n4737 GND.n4736 585
R12099 GND.n4717 GND.n4715 585
R12100 GND.n4715 GND.n4714 585
R12101 GND.n4726 GND.n4725 585
R12102 GND.n4725 GND.n2330 585
R12103 GND.n4724 GND.n4719 585
R12104 GND.n4724 GND.n2324 585
R12105 GND.n4723 GND.n4722 585
R12106 GND.n4723 GND.n2321 585
R12107 GND.n2304 GND.n2303 585
R12108 GND.n2957 GND.n2304 585
R12109 GND.n5574 GND.n5573 585
R12110 GND.n5573 GND.n5572 585
R12111 GND.n5575 GND.n2293 585
R12112 GND.n2961 GND.n2293 585
R12113 GND.n5577 GND.n5576 585
R12114 GND.n5578 GND.n5577 585
R12115 GND.n2294 GND.n2292 585
R12116 GND.n2292 GND.n2283 585
R12117 GND.n2297 GND.n2296 585
R12118 GND.n2296 GND.n2280 585
R12119 GND.n2268 GND.n2267 585
R12120 GND.n2968 GND.n2268 585
R12121 GND.n5595 GND.n5594 585
R12122 GND.n5594 GND.n5593 585
R12123 GND.n5596 GND.n2262 585
R12124 GND.n2974 GND.n2262 585
R12125 GND.n5598 GND.n5597 585
R12126 GND.n5599 GND.n5598 585
R12127 GND.n2250 GND.n2249 585
R12128 GND.n4583 GND.n2250 585
R12129 GND.n5609 GND.n5608 585
R12130 GND.n5608 GND.n5607 585
R12131 GND.n5610 GND.n2242 585
R12132 GND.n4594 GND.n2242 585
R12133 GND.n5612 GND.n5611 585
R12134 GND.n5613 GND.n5612 585
R12135 GND.n2243 GND.n2241 585
R12136 GND.n2241 GND.n2240 585
R12137 GND.n2219 GND.n2218 585
R12138 GND.n2228 GND.n2219 585
R12139 GND.n5628 GND.n5627 585
R12140 GND.n5627 GND.n5626 585
R12141 GND.n5629 GND.n2208 585
R12142 GND.n4553 GND.n2208 585
R12143 GND.n5631 GND.n5630 585
R12144 GND.n5632 GND.n5631 585
R12145 GND.n2209 GND.n2207 585
R12146 GND.n2207 GND.n2199 585
R12147 GND.n2212 GND.n2211 585
R12148 GND.n2211 GND.n2196 585
R12149 GND.n2184 GND.n2183 585
R12150 GND.n2989 GND.n2184 585
R12151 GND.n5649 GND.n5648 585
R12152 GND.n5648 GND.n5647 585
R12153 GND.n5650 GND.n2178 585
R12154 GND.n2995 GND.n2178 585
R12155 GND.n5652 GND.n5651 585
R12156 GND.n5653 GND.n5652 585
R12157 GND.n2166 GND.n2165 585
R12158 GND.n4514 GND.n2166 585
R12159 GND.n5663 GND.n5662 585
R12160 GND.n5662 GND.n5661 585
R12161 GND.n5664 GND.n2160 585
R12162 GND.n3001 GND.n2160 585
R12163 GND.n5666 GND.n5665 585
R12164 GND.n5667 GND.n5666 585
R12165 GND.n2148 GND.n2147 585
R12166 GND.n4354 GND.n2148 585
R12167 GND.n5677 GND.n5676 585
R12168 GND.n5676 GND.n5675 585
R12169 GND.n5678 GND.n2142 585
R12170 GND.n4365 GND.n2142 585
R12171 GND.n5680 GND.n5679 585
R12172 GND.n5681 GND.n5680 585
R12173 GND.n2131 GND.n2130 585
R12174 GND.n4371 GND.n2131 585
R12175 GND.n5691 GND.n5690 585
R12176 GND.n5690 GND.n5689 585
R12177 GND.n5692 GND.n2125 585
R12178 GND.n3017 GND.n2125 585
R12179 GND.n5694 GND.n5693 585
R12180 GND.n5695 GND.n5694 585
R12181 GND.n2113 GND.n2112 585
R12182 GND.n4385 GND.n2113 585
R12183 GND.n5705 GND.n5704 585
R12184 GND.n5704 GND.n5703 585
R12185 GND.n5706 GND.n2107 585
R12186 GND.n3038 GND.n2107 585
R12187 GND.n5708 GND.n5707 585
R12188 GND.n5709 GND.n5708 585
R12189 GND.n2095 GND.n2094 585
R12190 GND.n4400 GND.n2095 585
R12191 GND.n5719 GND.n5718 585
R12192 GND.n5718 GND.n5717 585
R12193 GND.n5720 GND.n2084 585
R12194 GND.n4408 GND.n2084 585
R12195 GND.n5722 GND.n5721 585
R12196 GND.n5723 GND.n5722 585
R12197 GND.n2085 GND.n2083 585
R12198 GND.n3050 GND.n2083 585
R12199 GND.n2088 GND.n2087 585
R12200 GND.n2087 GND.n2063 585
R12201 GND.n2051 GND.n2050 585
R12202 GND.n2060 GND.n2051 585
R12203 GND.n5740 GND.n5739 585
R12204 GND.n5739 GND.n5738 585
R12205 GND.n5741 GND.n2040 585
R12206 GND.n4332 GND.n2040 585
R12207 GND.n5743 GND.n5742 585
R12208 GND.n5744 GND.n5743 585
R12209 GND.n2041 GND.n2039 585
R12210 GND.n2039 GND.n2030 585
R12211 GND.n2044 GND.n2043 585
R12212 GND.n2043 GND.n2027 585
R12213 GND.n2015 GND.n2014 585
R12214 GND.n3057 GND.n2015 585
R12215 GND.n5760 GND.n5759 585
R12216 GND.n5759 GND.n5758 585
R12217 GND.n5761 GND.n1992 585
R12218 GND.n3063 GND.n1992 585
R12219 GND.n5763 GND.n5762 585
R12220 GND.n5764 GND.n5763 585
R12221 GND.n1993 GND.n1991 585
R12222 GND.n4277 GND.n1991 585
R12223 GND.n2008 GND.n2007 585
R12224 GND.n2007 GND.n1981 585
R12225 GND.n2006 GND.n1995 585
R12226 GND.n2006 GND.n1972 585
R12227 GND.n2005 GND.n2004 585
R12228 GND.n2005 GND.n1969 585
R12229 GND.n1997 GND.n1996 585
R12230 GND.n1996 GND.n1965 585
R12231 GND.n2000 GND.n1999 585
R12232 GND.n1999 GND.n1904 585
R12233 GND.n1893 GND.n1892 585
R12234 GND.n1902 GND.n1893 585
R12235 GND.n5799 GND.n5798 585
R12236 GND.n5798 GND.n5797 585
R12237 GND.n5800 GND.n1887 585
R12238 GND.n1954 GND.n1887 585
R12239 GND.n5802 GND.n5801 585
R12240 GND.n5803 GND.n5802 585
R12241 GND.n1888 GND.n1886 585
R12242 GND.n1886 GND.n1883 585
R12243 GND.n4108 GND.n4107 585
R12244 GND.n4108 GND.n1847 585
R12245 GND.n4110 GND.n4109 585
R12246 GND.n4109 GND.n1827 585
R12247 GND.n4111 GND.n4100 585
R12248 GND.n4113 GND.n4100 585
R12249 GND.n4115 GND.n4112 585
R12250 GND.n4115 GND.n4114 585
R12251 GND.n4116 GND.n4099 585
R12252 GND.n4116 GND.n1756 585
R12253 GND.n4118 GND.n4117 585
R12254 GND.n4117 GND.n1750 585
R12255 GND.n4119 GND.n4094 585
R12256 GND.n4094 GND.n3187 585
R12257 GND.n4121 GND.n4120 585
R12258 GND.n4121 GND.n3186 585
R12259 GND.n4122 GND.n4093 585
R12260 GND.n4122 GND.n3190 585
R12261 GND.n4124 GND.n4123 585
R12262 GND.n4123 GND.n3198 585
R12263 GND.n4125 GND.n3208 585
R12264 GND.n3208 GND.n3196 585
R12265 GND.n4127 GND.n4126 585
R12266 GND.n4128 GND.n4127 585
R12267 GND.n3209 GND.n3207 585
R12268 GND.n3215 GND.n3207 585
R12269 GND.n4087 GND.n4086 585
R12270 GND.n4086 GND.n4085 585
R12271 GND.n3212 GND.n3211 585
R12272 GND.n3226 GND.n3212 585
R12273 GND.n4055 GND.n3237 585
R12274 GND.n3237 GND.n3223 585
R12275 GND.n4057 GND.n4056 585
R12276 GND.n4058 GND.n4057 585
R12277 GND.n3238 GND.n3236 585
R12278 GND.n3245 GND.n3236 585
R12279 GND.n4050 GND.n4049 585
R12280 GND.n4049 GND.n4048 585
R12281 GND.n3241 GND.n3240 585
R12282 GND.n3255 GND.n3241 585
R12283 GND.n4018 GND.n3266 585
R12284 GND.n3266 GND.n3253 585
R12285 GND.n4020 GND.n4019 585
R12286 GND.n4021 GND.n4020 585
R12287 GND.n3267 GND.n3265 585
R12288 GND.n3274 GND.n3265 585
R12289 GND.n4013 GND.n4012 585
R12290 GND.n4012 GND.n4011 585
R12291 GND.n3270 GND.n3269 585
R12292 GND.n3284 GND.n3270 585
R12293 GND.n3981 GND.n3296 585
R12294 GND.n3296 GND.n3282 585
R12295 GND.n3983 GND.n3982 585
R12296 GND.n3984 GND.n3983 585
R12297 GND.n3297 GND.n3295 585
R12298 GND.n3303 GND.n3295 585
R12299 GND.n3976 GND.n3975 585
R12300 GND.n3975 GND.n3974 585
R12301 GND.n3300 GND.n3299 585
R12302 GND.n3312 GND.n3300 585
R12303 GND.n3946 GND.n3945 585
R12304 GND.n3947 GND.n3946 585
R12305 GND.n3324 GND.n3323 585
R12306 GND.n3323 GND.n3321 585
R12307 GND.n3892 GND.n3891 585
R12308 GND.n3892 GND.n3853 585
R12309 GND.n3894 GND.n3893 585
R12310 GND.n3893 GND.n3860 585
R12311 GND.n3896 GND.n3895 585
R12312 GND.n3896 GND.n3857 585
R12313 GND.n3899 GND.n3898 585
R12314 GND.n3900 GND.n3899 585
R12315 GND.n3897 GND.n3890 585
R12316 GND.n3890 GND.n3889 585
R12317 GND.n3874 GND.n3864 585
R12318 GND.n3865 GND.n3864 585
R12319 GND.n3876 GND.n3875 585
R12320 GND.n3877 GND.n3876 585
R12321 GND.n3873 GND.n3872 585
R12322 GND.n3873 GND.n3347 585
R12323 GND.n3871 GND.n3870 585
R12324 GND.n3870 GND.n3345 585
R12325 GND.n3335 GND.n3333 585
R12326 GND.n3337 GND.n3335 585
R12327 GND.n3940 GND.n3939 585
R12328 GND.n3939 GND.n3938 585
R12329 GND.n3334 GND.n3332 585
R12330 GND.n3358 GND.n3334 585
R12331 GND.n3801 GND.n3800 585
R12332 GND.n3801 GND.n3361 585
R12333 GND.n3803 GND.n3802 585
R12334 GND.n3802 GND.n3369 585
R12335 GND.n3804 GND.n3382 585
R12336 GND.n3382 GND.n3367 585
R12337 GND.n3806 GND.n3805 585
R12338 GND.n3807 GND.n3806 585
R12339 GND.n3383 GND.n3381 585
R12340 GND.n3389 GND.n3381 585
R12341 GND.n3793 GND.n3792 585
R12342 GND.n3792 GND.n3791 585
R12343 GND.n3386 GND.n3385 585
R12344 GND.n3400 GND.n3386 585
R12345 GND.n3761 GND.n3411 585
R12346 GND.n3411 GND.n3397 585
R12347 GND.n3763 GND.n3762 585
R12348 GND.n3764 GND.n3763 585
R12349 GND.n3412 GND.n3410 585
R12350 GND.n3419 GND.n3410 585
R12351 GND.n3756 GND.n3755 585
R12352 GND.n3755 GND.n3754 585
R12353 GND.n3415 GND.n3414 585
R12354 GND.n3429 GND.n3415 585
R12355 GND.n3724 GND.n3440 585
R12356 GND.n3440 GND.n3427 585
R12357 GND.n3726 GND.n3725 585
R12358 GND.n3727 GND.n3726 585
R12359 GND.n3441 GND.n3439 585
R12360 GND.n3448 GND.n3439 585
R12361 GND.n3719 GND.n3718 585
R12362 GND.n3718 GND.n3717 585
R12363 GND.n3444 GND.n3443 585
R12364 GND.n3458 GND.n3444 585
R12365 GND.n3687 GND.n3470 585
R12366 GND.n3470 GND.n3456 585
R12367 GND.n3689 GND.n3688 585
R12368 GND.n3690 GND.n3689 585
R12369 GND.n3471 GND.n3469 585
R12370 GND.n3477 GND.n3469 585
R12371 GND.n3682 GND.n3681 585
R12372 GND.n3681 GND.n3680 585
R12373 GND.n3474 GND.n3473 585
R12374 GND.n3668 GND.n3474 585
R12375 GND.n3490 GND.n3489 585
R12376 GND.n3491 GND.n3490 585
R12377 GND.n3485 GND.n3484 585
R12378 GND.n3484 GND.n1647 585
R12379 GND.n1614 GND.n1613 585
R12380 GND.n6005 GND.n1614 585
R12381 GND.n6008 GND.n6007 585
R12382 GND.n6007 GND.n6006 585
R12383 GND.n6009 GND.n1608 585
R12384 GND.n1608 GND.n1607 585
R12385 GND.n6011 GND.n6010 585
R12386 GND.n6012 GND.n6011 585
R12387 GND.n1606 GND.n1605 585
R12388 GND.n6013 GND.n1606 585
R12389 GND.n6016 GND.n6015 585
R12390 GND.n6015 GND.n6014 585
R12391 GND.n6017 GND.n1600 585
R12392 GND.n1600 GND.n1599 585
R12393 GND.n6019 GND.n6018 585
R12394 GND.n6020 GND.n6019 585
R12395 GND.n1598 GND.n1597 585
R12396 GND.n6021 GND.n1598 585
R12397 GND.n6024 GND.n6023 585
R12398 GND.n6023 GND.n6022 585
R12399 GND.n6025 GND.n1592 585
R12400 GND.n1592 GND.n1591 585
R12401 GND.n6027 GND.n6026 585
R12402 GND.n6028 GND.n6027 585
R12403 GND.n1590 GND.n1589 585
R12404 GND.n6029 GND.n1590 585
R12405 GND.n6032 GND.n6031 585
R12406 GND.n6031 GND.n6030 585
R12407 GND.n6033 GND.n1584 585
R12408 GND.n1584 GND.n1583 585
R12409 GND.n6035 GND.n6034 585
R12410 GND.n6036 GND.n6035 585
R12411 GND.n1582 GND.n1581 585
R12412 GND.n6037 GND.n1582 585
R12413 GND.n6040 GND.n6039 585
R12414 GND.n6039 GND.n6038 585
R12415 GND.n6041 GND.n1576 585
R12416 GND.n1576 GND.n1575 585
R12417 GND.n6043 GND.n6042 585
R12418 GND.n6044 GND.n6043 585
R12419 GND.n1574 GND.n1573 585
R12420 GND.n6045 GND.n1574 585
R12421 GND.n6048 GND.n6047 585
R12422 GND.n6047 GND.n6046 585
R12423 GND.n6049 GND.n1568 585
R12424 GND.n1568 GND.n1567 585
R12425 GND.n6051 GND.n6050 585
R12426 GND.n6052 GND.n6051 585
R12427 GND.n1566 GND.n1565 585
R12428 GND.n6053 GND.n1566 585
R12429 GND.n6056 GND.n6055 585
R12430 GND.n6055 GND.n6054 585
R12431 GND.n6057 GND.n1560 585
R12432 GND.n1560 GND.n1559 585
R12433 GND.n6059 GND.n6058 585
R12434 GND.n6060 GND.n6059 585
R12435 GND.n1558 GND.n1557 585
R12436 GND.n6061 GND.n1558 585
R12437 GND.n6064 GND.n6063 585
R12438 GND.n6063 GND.n6062 585
R12439 GND.n6065 GND.n1552 585
R12440 GND.n1552 GND.n1551 585
R12441 GND.n6067 GND.n6066 585
R12442 GND.n6068 GND.n6067 585
R12443 GND.n1550 GND.n1549 585
R12444 GND.n6069 GND.n1550 585
R12445 GND.n6072 GND.n6071 585
R12446 GND.n6071 GND.n6070 585
R12447 GND.n6073 GND.n1544 585
R12448 GND.n1544 GND.n1543 585
R12449 GND.n6075 GND.n6074 585
R12450 GND.n6076 GND.n6075 585
R12451 GND.n1542 GND.n1541 585
R12452 GND.n6077 GND.n1542 585
R12453 GND.n6080 GND.n6079 585
R12454 GND.n6079 GND.n6078 585
R12455 GND.n6081 GND.n1536 585
R12456 GND.n1536 GND.n1535 585
R12457 GND.n6083 GND.n6082 585
R12458 GND.n6084 GND.n6083 585
R12459 GND.n1534 GND.n1533 585
R12460 GND.n6085 GND.n1534 585
R12461 GND.n6088 GND.n6087 585
R12462 GND.n6087 GND.n6086 585
R12463 GND.n6089 GND.n1528 585
R12464 GND.n1528 GND.n1527 585
R12465 GND.n6091 GND.n6090 585
R12466 GND.n6092 GND.n6091 585
R12467 GND.n1526 GND.n1525 585
R12468 GND.n6093 GND.n1526 585
R12469 GND.n6096 GND.n6095 585
R12470 GND.n6095 GND.n6094 585
R12471 GND.n6097 GND.n1520 585
R12472 GND.n1520 GND.n1519 585
R12473 GND.n6099 GND.n6098 585
R12474 GND.n6100 GND.n6099 585
R12475 GND.n1518 GND.n1517 585
R12476 GND.n6101 GND.n1518 585
R12477 GND.n6104 GND.n6103 585
R12478 GND.n6103 GND.n6102 585
R12479 GND.n6105 GND.n1512 585
R12480 GND.n1512 GND.n1511 585
R12481 GND.n6107 GND.n6106 585
R12482 GND.n6108 GND.n6107 585
R12483 GND.n1510 GND.n1509 585
R12484 GND.n6109 GND.n1510 585
R12485 GND.n6112 GND.n6111 585
R12486 GND.n6111 GND.n6110 585
R12487 GND.n6113 GND.n1504 585
R12488 GND.n1504 GND.n1503 585
R12489 GND.n6115 GND.n6114 585
R12490 GND.n6116 GND.n6115 585
R12491 GND.n1502 GND.n1501 585
R12492 GND.n6117 GND.n1502 585
R12493 GND.n6120 GND.n6119 585
R12494 GND.n6119 GND.n6118 585
R12495 GND.n6121 GND.n1496 585
R12496 GND.n1496 GND.n1495 585
R12497 GND.n6123 GND.n6122 585
R12498 GND.n6124 GND.n6123 585
R12499 GND.n1494 GND.n1493 585
R12500 GND.n6125 GND.n1494 585
R12501 GND.n6128 GND.n6127 585
R12502 GND.n6127 GND.n6126 585
R12503 GND.n6129 GND.n1488 585
R12504 GND.n1488 GND.n1487 585
R12505 GND.n6131 GND.n6130 585
R12506 GND.n6132 GND.n6131 585
R12507 GND.n1486 GND.n1485 585
R12508 GND.n6133 GND.n1486 585
R12509 GND.n6136 GND.n6135 585
R12510 GND.n6135 GND.n6134 585
R12511 GND.n6137 GND.n1480 585
R12512 GND.n1480 GND.n1479 585
R12513 GND.n6139 GND.n6138 585
R12514 GND.n6140 GND.n6139 585
R12515 GND.n1478 GND.n1477 585
R12516 GND.n6141 GND.n1478 585
R12517 GND.n6144 GND.n6143 585
R12518 GND.n6143 GND.n6142 585
R12519 GND.n6145 GND.n1472 585
R12520 GND.n1472 GND.n1471 585
R12521 GND.n6147 GND.n6146 585
R12522 GND.n6148 GND.n6147 585
R12523 GND.n1470 GND.n1469 585
R12524 GND.n6149 GND.n1470 585
R12525 GND.n6152 GND.n6151 585
R12526 GND.n6151 GND.n6150 585
R12527 GND.n6153 GND.n1464 585
R12528 GND.n1464 GND.n1463 585
R12529 GND.n6155 GND.n6154 585
R12530 GND.n6156 GND.n6155 585
R12531 GND.n1462 GND.n1461 585
R12532 GND.n6157 GND.n1462 585
R12533 GND.n6160 GND.n6159 585
R12534 GND.n6159 GND.n6158 585
R12535 GND.n6161 GND.n1456 585
R12536 GND.n1456 GND.n1455 585
R12537 GND.n6163 GND.n6162 585
R12538 GND.n6164 GND.n6163 585
R12539 GND.n1454 GND.n1453 585
R12540 GND.n6165 GND.n1454 585
R12541 GND.n6168 GND.n6167 585
R12542 GND.n6167 GND.n6166 585
R12543 GND.n6169 GND.n1447 585
R12544 GND.n1447 GND.n1446 585
R12545 GND.n6171 GND.n6170 585
R12546 GND.n6172 GND.n6171 585
R12547 GND.n1448 GND.n1445 585
R12548 GND.n6173 GND.n1445 585
R12549 GND.n6003 GND.n6002 585
R12550 GND.n6004 GND.n6003 585
R12551 GND.n6001 GND.n1649 585
R12552 GND.n1653 GND.n1651 585
R12553 GND.n5997 GND.n1654 585
R12554 GND.n5996 GND.n1655 585
R12555 GND.n5995 GND.n1656 585
R12556 GND.n1659 GND.n1657 585
R12557 GND.n5991 GND.n1660 585
R12558 GND.n5990 GND.n1661 585
R12559 GND.n5989 GND.n1662 585
R12560 GND.n1666 GND.n1663 585
R12561 GND.n5985 GND.n1646 585
R12562 GND.n6004 GND.n1646 585
R12563 GND.n4222 GND.n3101 585
R12564 GND.n4223 GND.n4222 585
R12565 GND.n4150 GND.n3189 585
R12566 GND.n4150 GND.n4149 585
R12567 GND.n3201 GND.n3188 585
R12568 GND.n4133 GND.n3188 585
R12569 GND.n4139 GND.n4138 585
R12570 GND.n4140 GND.n4139 585
R12571 GND.n3200 GND.n3199 585
R12572 GND.n4130 GND.n3199 585
R12573 GND.n4065 GND.n4064 585
R12574 GND.n4064 GND.n3206 585
R12575 GND.n4063 GND.n3216 585
R12576 GND.n4084 GND.n3216 585
R12577 GND.n3230 GND.n3228 585
R12578 GND.n3228 GND.n3213 585
R12579 GND.n4073 GND.n4072 585
R12580 GND.n4074 GND.n4073 585
R12581 GND.n3229 GND.n3227 585
R12582 GND.n4059 GND.n3227 585
R12583 GND.n4028 GND.n4027 585
R12584 GND.n4027 GND.n3235 585
R12585 GND.n4026 GND.n3246 585
R12586 GND.n4047 GND.n3246 585
R12587 GND.n3259 GND.n3257 585
R12588 GND.n3257 GND.n3243 585
R12589 GND.n4036 GND.n4035 585
R12590 GND.n4037 GND.n4036 585
R12591 GND.n3258 GND.n3256 585
R12592 GND.n4022 GND.n3256 585
R12593 GND.n3991 GND.n3990 585
R12594 GND.n3990 GND.n3264 585
R12595 GND.n3989 GND.n3275 585
R12596 GND.n4010 GND.n3275 585
R12597 GND.n3288 GND.n3286 585
R12598 GND.n3286 GND.n3271 585
R12599 GND.n3999 GND.n3998 585
R12600 GND.n4000 GND.n3999 585
R12601 GND.n3287 GND.n3285 585
R12602 GND.n3985 GND.n3285 585
R12603 GND.n3954 GND.n3953 585
R12604 GND.n3953 GND.n3294 585
R12605 GND.n3952 GND.n3304 585
R12606 GND.n3973 GND.n3304 585
R12607 GND.n3316 GND.n3314 585
R12608 GND.n3314 GND.n3301 585
R12609 GND.n3962 GND.n3961 585
R12610 GND.n3963 GND.n3962 585
R12611 GND.n3315 GND.n3313 585
R12612 GND.n3948 GND.n3313 585
R12613 GND.n3914 GND.n3913 585
R12614 GND.n3913 GND.n3912 585
R12615 GND.n3852 GND.n3851 585
R12616 GND.n3859 GND.n3852 585
R12617 GND.n3904 GND.n3850 585
R12618 GND.n3905 GND.n3904 585
R12619 GND.n3903 GND.n3862 585
R12620 GND.n3903 GND.n3902 585
R12621 GND.n3861 GND.n3844 585
R12622 GND.n3863 GND.n3861 585
R12623 GND.n3867 GND.n3843 585
R12624 GND.n3888 GND.n3867 585
R12625 GND.n3878 GND.n3842 585
R12626 GND.n3879 GND.n3878 585
R12627 GND.n3351 GND.n3349 585
R12628 GND.n3869 GND.n3349 585
R12629 GND.n3929 GND.n3928 585
R12630 GND.n3930 GND.n3929 585
R12631 GND.n3350 GND.n3348 585
R12632 GND.n3836 GND.n3348 585
R12633 GND.n3833 GND.n3338 585
R12634 GND.n3937 GND.n3338 585
R12635 GND.n3832 GND.n3831 585
R12636 GND.n3831 GND.n3830 585
R12637 GND.n3357 GND.n3356 585
R12638 GND.n3826 GND.n3357 585
R12639 GND.n3374 GND.n3372 585
R12640 GND.n3372 GND.n3371 585
R12641 GND.n3816 GND.n3815 585
R12642 GND.n3817 GND.n3816 585
R12643 GND.n3373 GND.n3370 585
R12644 GND.n3809 GND.n3370 585
R12645 GND.n3771 GND.n3770 585
R12646 GND.n3770 GND.n3380 585
R12647 GND.n3769 GND.n3390 585
R12648 GND.n3790 GND.n3390 585
R12649 GND.n3404 GND.n3402 585
R12650 GND.n3402 GND.n3387 585
R12651 GND.n3779 GND.n3778 585
R12652 GND.n3780 GND.n3779 585
R12653 GND.n3403 GND.n3401 585
R12654 GND.n3765 GND.n3401 585
R12655 GND.n3734 GND.n3733 585
R12656 GND.n3733 GND.n3409 585
R12657 GND.n3732 GND.n3420 585
R12658 GND.n3753 GND.n3420 585
R12659 GND.n3433 GND.n3431 585
R12660 GND.n3431 GND.n3417 585
R12661 GND.n3742 GND.n3741 585
R12662 GND.n3743 GND.n3742 585
R12663 GND.n3432 GND.n3430 585
R12664 GND.n3728 GND.n3430 585
R12665 GND.n3697 GND.n3696 585
R12666 GND.n3696 GND.n3438 585
R12667 GND.n3695 GND.n3449 585
R12668 GND.n3716 GND.n3449 585
R12669 GND.n3462 GND.n3460 585
R12670 GND.n3460 GND.n3445 585
R12671 GND.n3705 GND.n3704 585
R12672 GND.n3706 GND.n3705 585
R12673 GND.n3461 GND.n3459 585
R12674 GND.n3691 GND.n3459 585
R12675 GND.n3660 GND.n3659 585
R12676 GND.n3659 GND.n3468 585
R12677 GND.n3658 GND.n3478 585
R12678 GND.n3679 GND.n3478 585
R12679 GND.n3657 GND.n3656 585
R12680 GND.n3656 GND.n3475 585
R12681 GND.n3655 GND.n1648 585
R12682 GND.n3669 GND.n1648 585
R12683 GND.n5892 GND.n5891 585
R12684 GND.n1749 GND.n1747 585
R12685 GND.n4193 GND.n4183 585
R12686 GND.n4194 GND.n4182 585
R12687 GND.n4181 GND.n4173 585
R12688 GND.n4204 GND.n4172 585
R12689 GND.n4205 GND.n4171 585
R12690 GND.n4162 GND.n4161 585
R12691 GND.n4212 GND.n4160 585
R12692 GND.n4213 GND.n4159 585
R12693 GND.n4158 GND.n4151 585
R12694 GND.n4221 GND.n4220 585
R12695 GND.n1748 GND.n1742 585
R12696 GND.n4223 GND.n1748 585
R12697 GND.n5897 GND.n1741 585
R12698 GND.n4149 GND.n1741 585
R12699 GND.n5898 GND.n1740 585
R12700 GND.n4133 GND.n1740 585
R12701 GND.n5899 GND.n1739 585
R12702 GND.n4140 GND.n1739 585
R12703 GND.n4129 GND.n1737 585
R12704 GND.n4130 GND.n4129 585
R12705 GND.n5903 GND.n1736 585
R12706 GND.n3206 GND.n1736 585
R12707 GND.n5904 GND.n1735 585
R12708 GND.n4084 GND.n1735 585
R12709 GND.n5905 GND.n1734 585
R12710 GND.n3213 GND.n1734 585
R12711 GND.n3225 GND.n1732 585
R12712 GND.n4074 GND.n3225 585
R12713 GND.n5909 GND.n1731 585
R12714 GND.n4059 GND.n1731 585
R12715 GND.n5910 GND.n1730 585
R12716 GND.n3235 GND.n1730 585
R12717 GND.n5911 GND.n1729 585
R12718 GND.n4047 GND.n1729 585
R12719 GND.n3242 GND.n1727 585
R12720 GND.n3243 GND.n3242 585
R12721 GND.n5915 GND.n1726 585
R12722 GND.n4037 GND.n1726 585
R12723 GND.n5916 GND.n1725 585
R12724 GND.n4022 GND.n1725 585
R12725 GND.n5917 GND.n1724 585
R12726 GND.n3264 GND.n1724 585
R12727 GND.n3273 GND.n1722 585
R12728 GND.n4010 GND.n3273 585
R12729 GND.n5921 GND.n1721 585
R12730 GND.n3271 GND.n1721 585
R12731 GND.n5922 GND.n1720 585
R12732 GND.n4000 GND.n1720 585
R12733 GND.n5923 GND.n1719 585
R12734 GND.n3985 GND.n1719 585
R12735 GND.n3293 GND.n1717 585
R12736 GND.n3294 GND.n3293 585
R12737 GND.n5927 GND.n1716 585
R12738 GND.n3973 GND.n1716 585
R12739 GND.n5928 GND.n1715 585
R12740 GND.n3301 GND.n1715 585
R12741 GND.n5929 GND.n1714 585
R12742 GND.n3963 GND.n1714 585
R12743 GND.n3322 GND.n1712 585
R12744 GND.n3948 GND.n3322 585
R12745 GND.n5933 GND.n1711 585
R12746 GND.n3912 GND.n1711 585
R12747 GND.n5934 GND.n1710 585
R12748 GND.n3859 GND.n1710 585
R12749 GND.n5935 GND.n1709 585
R12750 GND.n3905 GND.n1709 585
R12751 GND.n3901 GND.n1706 585
R12752 GND.n3902 GND.n3901 585
R12753 GND.n5939 GND.n1705 585
R12754 GND.n3863 GND.n1705 585
R12755 GND.n5940 GND.n1704 585
R12756 GND.n3888 GND.n1704 585
R12757 GND.n5941 GND.n1703 585
R12758 GND.n3879 GND.n1703 585
R12759 GND.n3868 GND.n1701 585
R12760 GND.n3869 GND.n3868 585
R12761 GND.n5945 GND.n1700 585
R12762 GND.n3930 GND.n1700 585
R12763 GND.n5946 GND.n1699 585
R12764 GND.n3836 GND.n1699 585
R12765 GND.n5947 GND.n1698 585
R12766 GND.n3937 GND.n1698 585
R12767 GND.n3829 GND.n1696 585
R12768 GND.n3830 GND.n3829 585
R12769 GND.n5951 GND.n1695 585
R12770 GND.n3826 GND.n1695 585
R12771 GND.n5952 GND.n1694 585
R12772 GND.n3371 GND.n1694 585
R12773 GND.n5953 GND.n1693 585
R12774 GND.n3817 GND.n1693 585
R12775 GND.n3808 GND.n1691 585
R12776 GND.n3809 GND.n3808 585
R12777 GND.n5957 GND.n1690 585
R12778 GND.n3380 GND.n1690 585
R12779 GND.n5958 GND.n1689 585
R12780 GND.n3790 GND.n1689 585
R12781 GND.n5959 GND.n1688 585
R12782 GND.n3387 GND.n1688 585
R12783 GND.n3399 GND.n1686 585
R12784 GND.n3780 GND.n3399 585
R12785 GND.n5963 GND.n1685 585
R12786 GND.n3765 GND.n1685 585
R12787 GND.n5964 GND.n1684 585
R12788 GND.n3409 GND.n1684 585
R12789 GND.n5965 GND.n1683 585
R12790 GND.n3753 GND.n1683 585
R12791 GND.n3416 GND.n1681 585
R12792 GND.n3417 GND.n3416 585
R12793 GND.n5969 GND.n1680 585
R12794 GND.n3743 GND.n1680 585
R12795 GND.n5970 GND.n1679 585
R12796 GND.n3728 GND.n1679 585
R12797 GND.n5971 GND.n1678 585
R12798 GND.n3438 GND.n1678 585
R12799 GND.n3447 GND.n1676 585
R12800 GND.n3716 GND.n3447 585
R12801 GND.n5975 GND.n1675 585
R12802 GND.n3445 GND.n1675 585
R12803 GND.n5976 GND.n1674 585
R12804 GND.n3706 GND.n1674 585
R12805 GND.n5977 GND.n1673 585
R12806 GND.n3691 GND.n1673 585
R12807 GND.n3467 GND.n1671 585
R12808 GND.n3468 GND.n3467 585
R12809 GND.n5981 GND.n1670 585
R12810 GND.n3679 GND.n1670 585
R12811 GND.n5982 GND.n1669 585
R12812 GND.n3475 GND.n1669 585
R12813 GND.n5983 GND.n1668 585
R12814 GND.n3669 GND.n1668 585
R12815 GND.n5449 GND.n2465 530.939
R12816 GND.n2508 GND.n2507 530.939
R12817 GND.n1949 GND.n1846 530.939
R12818 GND.n5845 GND.n1850 530.939
R12819 GND.n7563 GND.n7562 355.238
R12820 GND.n7340 GND.n7339 301.784
R12821 GND.n7341 GND.n7340 301.784
R12822 GND.n7341 GND.n673 301.784
R12823 GND.n7349 GND.n673 301.784
R12824 GND.n7350 GND.n7349 301.784
R12825 GND.n7351 GND.n7350 301.784
R12826 GND.n7351 GND.n667 301.784
R12827 GND.n7359 GND.n667 301.784
R12828 GND.n7360 GND.n7359 301.784
R12829 GND.n7361 GND.n7360 301.784
R12830 GND.n7361 GND.n661 301.784
R12831 GND.n7369 GND.n661 301.784
R12832 GND.n7370 GND.n7369 301.784
R12833 GND.n7371 GND.n7370 301.784
R12834 GND.n7371 GND.n655 301.784
R12835 GND.n7379 GND.n655 301.784
R12836 GND.n7380 GND.n7379 301.784
R12837 GND.n7381 GND.n7380 301.784
R12838 GND.n7381 GND.n649 301.784
R12839 GND.n7389 GND.n649 301.784
R12840 GND.n7390 GND.n7389 301.784
R12841 GND.n7391 GND.n7390 301.784
R12842 GND.n7391 GND.n643 301.784
R12843 GND.n7399 GND.n643 301.784
R12844 GND.n7400 GND.n7399 301.784
R12845 GND.n7401 GND.n7400 301.784
R12846 GND.n7401 GND.n637 301.784
R12847 GND.n7409 GND.n637 301.784
R12848 GND.n7410 GND.n7409 301.784
R12849 GND.n7411 GND.n7410 301.784
R12850 GND.n7411 GND.n631 301.784
R12851 GND.n7419 GND.n631 301.784
R12852 GND.n7420 GND.n7419 301.784
R12853 GND.n7421 GND.n7420 301.784
R12854 GND.n7421 GND.n625 301.784
R12855 GND.n7429 GND.n625 301.784
R12856 GND.n7430 GND.n7429 301.784
R12857 GND.n7431 GND.n7430 301.784
R12858 GND.n7431 GND.n619 301.784
R12859 GND.n7439 GND.n619 301.784
R12860 GND.n7440 GND.n7439 301.784
R12861 GND.n7441 GND.n7440 301.784
R12862 GND.n7441 GND.n613 301.784
R12863 GND.n7449 GND.n613 301.784
R12864 GND.n7450 GND.n7449 301.784
R12865 GND.n7451 GND.n7450 301.784
R12866 GND.n7451 GND.n607 301.784
R12867 GND.n7459 GND.n607 301.784
R12868 GND.n7460 GND.n7459 301.784
R12869 GND.n7461 GND.n7460 301.784
R12870 GND.n7461 GND.n601 301.784
R12871 GND.n7469 GND.n601 301.784
R12872 GND.n7470 GND.n7469 301.784
R12873 GND.n7471 GND.n7470 301.784
R12874 GND.n7471 GND.n595 301.784
R12875 GND.n7479 GND.n595 301.784
R12876 GND.n7480 GND.n7479 301.784
R12877 GND.n7481 GND.n7480 301.784
R12878 GND.n7481 GND.n589 301.784
R12879 GND.n7489 GND.n589 301.784
R12880 GND.n7490 GND.n7489 301.784
R12881 GND.n7491 GND.n7490 301.784
R12882 GND.n7491 GND.n583 301.784
R12883 GND.n7499 GND.n583 301.784
R12884 GND.n7500 GND.n7499 301.784
R12885 GND.n7501 GND.n7500 301.784
R12886 GND.n7501 GND.n577 301.784
R12887 GND.n7509 GND.n577 301.784
R12888 GND.n7510 GND.n7509 301.784
R12889 GND.n7511 GND.n7510 301.784
R12890 GND.n7511 GND.n571 301.784
R12891 GND.n7519 GND.n571 301.784
R12892 GND.n7520 GND.n7519 301.784
R12893 GND.n7521 GND.n7520 301.784
R12894 GND.n7521 GND.n565 301.784
R12895 GND.n7529 GND.n565 301.784
R12896 GND.n7530 GND.n7529 301.784
R12897 GND.n7531 GND.n7530 301.784
R12898 GND.n7531 GND.n559 301.784
R12899 GND.n7539 GND.n559 301.784
R12900 GND.n7540 GND.n7539 301.784
R12901 GND.n7541 GND.n7540 301.784
R12902 GND.n7541 GND.n553 301.784
R12903 GND.n7549 GND.n553 301.784
R12904 GND.n7550 GND.n7549 301.784
R12905 GND.n7551 GND.n7550 301.784
R12906 GND.n7551 GND.n547 301.784
R12907 GND.n7561 GND.n547 301.784
R12908 GND.n7562 GND.n7561 301.784
R12909 GND.n6359 GND.n6358 280.613
R12910 GND.n6360 GND.n6359 280.613
R12911 GND.n6360 GND.n1260 280.613
R12912 GND.n6368 GND.n1260 280.613
R12913 GND.n6369 GND.n6368 280.613
R12914 GND.n6370 GND.n6369 280.613
R12915 GND.n6370 GND.n1254 280.613
R12916 GND.n6378 GND.n1254 280.613
R12917 GND.n6379 GND.n6378 280.613
R12918 GND.n6380 GND.n6379 280.613
R12919 GND.n6380 GND.n1248 280.613
R12920 GND.n6388 GND.n1248 280.613
R12921 GND.n6389 GND.n6388 280.613
R12922 GND.n6390 GND.n6389 280.613
R12923 GND.n6390 GND.n1242 280.613
R12924 GND.n6398 GND.n1242 280.613
R12925 GND.n6399 GND.n6398 280.613
R12926 GND.n6400 GND.n6399 280.613
R12927 GND.n6400 GND.n1236 280.613
R12928 GND.n6408 GND.n1236 280.613
R12929 GND.n6409 GND.n6408 280.613
R12930 GND.n6410 GND.n6409 280.613
R12931 GND.n6410 GND.n1230 280.613
R12932 GND.n6418 GND.n1230 280.613
R12933 GND.n6419 GND.n6418 280.613
R12934 GND.n6420 GND.n6419 280.613
R12935 GND.n6420 GND.n1224 280.613
R12936 GND.n6428 GND.n1224 280.613
R12937 GND.n6429 GND.n6428 280.613
R12938 GND.n6430 GND.n6429 280.613
R12939 GND.n6430 GND.n1218 280.613
R12940 GND.n6438 GND.n1218 280.613
R12941 GND.n6439 GND.n6438 280.613
R12942 GND.n6440 GND.n6439 280.613
R12943 GND.n6440 GND.n1212 280.613
R12944 GND.n6448 GND.n1212 280.613
R12945 GND.n6449 GND.n6448 280.613
R12946 GND.n6450 GND.n6449 280.613
R12947 GND.n6450 GND.n1206 280.613
R12948 GND.n6458 GND.n1206 280.613
R12949 GND.n6459 GND.n6458 280.613
R12950 GND.n6460 GND.n6459 280.613
R12951 GND.n6460 GND.n1200 280.613
R12952 GND.n6468 GND.n1200 280.613
R12953 GND.n6469 GND.n6468 280.613
R12954 GND.n6470 GND.n6469 280.613
R12955 GND.n6470 GND.n1194 280.613
R12956 GND.n6478 GND.n1194 280.613
R12957 GND.n6479 GND.n6478 280.613
R12958 GND.n6480 GND.n6479 280.613
R12959 GND.n6480 GND.n1188 280.613
R12960 GND.n6488 GND.n1188 280.613
R12961 GND.n6489 GND.n6488 280.613
R12962 GND.n6490 GND.n6489 280.613
R12963 GND.n6490 GND.n1182 280.613
R12964 GND.n6498 GND.n1182 280.613
R12965 GND.n6499 GND.n6498 280.613
R12966 GND.n6500 GND.n6499 280.613
R12967 GND.n6500 GND.n1176 280.613
R12968 GND.n6508 GND.n1176 280.613
R12969 GND.n6509 GND.n6508 280.613
R12970 GND.n6510 GND.n6509 280.613
R12971 GND.n6510 GND.n1170 280.613
R12972 GND.n6518 GND.n1170 280.613
R12973 GND.n6519 GND.n6518 280.613
R12974 GND.n6520 GND.n6519 280.613
R12975 GND.n6520 GND.n1164 280.613
R12976 GND.n6528 GND.n1164 280.613
R12977 GND.n6529 GND.n6528 280.613
R12978 GND.n6530 GND.n6529 280.613
R12979 GND.n6530 GND.n1158 280.613
R12980 GND.n6538 GND.n1158 280.613
R12981 GND.n6539 GND.n6538 280.613
R12982 GND.n6540 GND.n6539 280.613
R12983 GND.n6540 GND.n1152 280.613
R12984 GND.n6548 GND.n1152 280.613
R12985 GND.n6549 GND.n6548 280.613
R12986 GND.n6550 GND.n6549 280.613
R12987 GND.n6550 GND.n1146 280.613
R12988 GND.n6558 GND.n1146 280.613
R12989 GND.n6559 GND.n6558 280.613
R12990 GND.n6560 GND.n6559 280.613
R12991 GND.n6560 GND.n1140 280.613
R12992 GND.n6568 GND.n1140 280.613
R12993 GND.n6569 GND.n6568 280.613
R12994 GND.n6570 GND.n6569 280.613
R12995 GND.n6570 GND.n1134 280.613
R12996 GND.n6578 GND.n1134 280.613
R12997 GND.n6579 GND.n6578 280.613
R12998 GND.n6580 GND.n6579 280.613
R12999 GND.n6580 GND.n1128 280.613
R13000 GND.n6588 GND.n1128 280.613
R13001 GND.n6589 GND.n6588 280.613
R13002 GND.n6590 GND.n6589 280.613
R13003 GND.n6590 GND.n1122 280.613
R13004 GND.n6598 GND.n1122 280.613
R13005 GND.n6599 GND.n6598 280.613
R13006 GND.n6600 GND.n6599 280.613
R13007 GND.n6600 GND.n1116 280.613
R13008 GND.n6608 GND.n1116 280.613
R13009 GND.n6609 GND.n6608 280.613
R13010 GND.n6610 GND.n6609 280.613
R13011 GND.n6610 GND.n1110 280.613
R13012 GND.n6618 GND.n1110 280.613
R13013 GND.n6619 GND.n6618 280.613
R13014 GND.n6620 GND.n6619 280.613
R13015 GND.n6620 GND.n1104 280.613
R13016 GND.n6628 GND.n1104 280.613
R13017 GND.n6629 GND.n6628 280.613
R13018 GND.n6630 GND.n6629 280.613
R13019 GND.n6630 GND.n1098 280.613
R13020 GND.n6638 GND.n1098 280.613
R13021 GND.n6639 GND.n6638 280.613
R13022 GND.n6640 GND.n6639 280.613
R13023 GND.n6640 GND.n1092 280.613
R13024 GND.n6648 GND.n1092 280.613
R13025 GND.n6649 GND.n6648 280.613
R13026 GND.n6650 GND.n6649 280.613
R13027 GND.n6650 GND.n1086 280.613
R13028 GND.n6658 GND.n1086 280.613
R13029 GND.n6659 GND.n6658 280.613
R13030 GND.n6660 GND.n6659 280.613
R13031 GND.n6660 GND.n1080 280.613
R13032 GND.n6668 GND.n1080 280.613
R13033 GND.n6669 GND.n6668 280.613
R13034 GND.n6670 GND.n6669 280.613
R13035 GND.n6670 GND.n1074 280.613
R13036 GND.n6678 GND.n1074 280.613
R13037 GND.n6679 GND.n6678 280.613
R13038 GND.n6680 GND.n6679 280.613
R13039 GND.n6680 GND.n1068 280.613
R13040 GND.n6688 GND.n1068 280.613
R13041 GND.n6689 GND.n6688 280.613
R13042 GND.n6690 GND.n6689 280.613
R13043 GND.n6690 GND.n1062 280.613
R13044 GND.n6698 GND.n1062 280.613
R13045 GND.n6699 GND.n6698 280.613
R13046 GND.n6700 GND.n6699 280.613
R13047 GND.n6700 GND.n1056 280.613
R13048 GND.n6708 GND.n1056 280.613
R13049 GND.n6709 GND.n6708 280.613
R13050 GND.n6710 GND.n6709 280.613
R13051 GND.n6710 GND.n1050 280.613
R13052 GND.n6718 GND.n1050 280.613
R13053 GND.n6719 GND.n6718 280.613
R13054 GND.n6720 GND.n6719 280.613
R13055 GND.n6720 GND.n1044 280.613
R13056 GND.n6728 GND.n1044 280.613
R13057 GND.n6729 GND.n6728 280.613
R13058 GND.n6730 GND.n6729 280.613
R13059 GND.n6730 GND.n1038 280.613
R13060 GND.n6738 GND.n1038 280.613
R13061 GND.n6739 GND.n6738 280.613
R13062 GND.n6740 GND.n6739 280.613
R13063 GND.n6740 GND.n1032 280.613
R13064 GND.n6748 GND.n1032 280.613
R13065 GND.n6749 GND.n6748 280.613
R13066 GND.n6750 GND.n6749 280.613
R13067 GND.n6750 GND.n1026 280.613
R13068 GND.n6758 GND.n1026 280.613
R13069 GND.n6759 GND.n6758 280.613
R13070 GND.n6760 GND.n6759 280.613
R13071 GND.n6760 GND.n1020 280.613
R13072 GND.n6768 GND.n1020 280.613
R13073 GND.n6769 GND.n6768 280.613
R13074 GND.n6770 GND.n6769 280.613
R13075 GND.n6770 GND.n1014 280.613
R13076 GND.n6778 GND.n1014 280.613
R13077 GND.n6779 GND.n6778 280.613
R13078 GND.n6780 GND.n6779 280.613
R13079 GND.n6780 GND.n1008 280.613
R13080 GND.n6788 GND.n1008 280.613
R13081 GND.n6789 GND.n6788 280.613
R13082 GND.n6790 GND.n6789 280.613
R13083 GND.n6790 GND.n1002 280.613
R13084 GND.n6798 GND.n1002 280.613
R13085 GND.n6799 GND.n6798 280.613
R13086 GND.n6800 GND.n6799 280.613
R13087 GND.n6800 GND.n996 280.613
R13088 GND.n6808 GND.n996 280.613
R13089 GND.n6809 GND.n6808 280.613
R13090 GND.n6810 GND.n6809 280.613
R13091 GND.n6810 GND.n990 280.613
R13092 GND.n6818 GND.n990 280.613
R13093 GND.n6819 GND.n6818 280.613
R13094 GND.n6820 GND.n6819 280.613
R13095 GND.n6820 GND.n984 280.613
R13096 GND.n6828 GND.n984 280.613
R13097 GND.n6829 GND.n6828 280.613
R13098 GND.n6830 GND.n6829 280.613
R13099 GND.n6830 GND.n978 280.613
R13100 GND.n6838 GND.n978 280.613
R13101 GND.n6839 GND.n6838 280.613
R13102 GND.n6840 GND.n6839 280.613
R13103 GND.n6840 GND.n972 280.613
R13104 GND.n6848 GND.n972 280.613
R13105 GND.n6849 GND.n6848 280.613
R13106 GND.n6850 GND.n6849 280.613
R13107 GND.n6850 GND.n966 280.613
R13108 GND.n6858 GND.n966 280.613
R13109 GND.n6859 GND.n6858 280.613
R13110 GND.n6860 GND.n6859 280.613
R13111 GND.n6860 GND.n960 280.613
R13112 GND.n6868 GND.n960 280.613
R13113 GND.n6869 GND.n6868 280.613
R13114 GND.n6870 GND.n6869 280.613
R13115 GND.n6870 GND.n954 280.613
R13116 GND.n6878 GND.n954 280.613
R13117 GND.n6879 GND.n6878 280.613
R13118 GND.n6880 GND.n6879 280.613
R13119 GND.n6880 GND.n948 280.613
R13120 GND.n6888 GND.n948 280.613
R13121 GND.n6889 GND.n6888 280.613
R13122 GND.n6890 GND.n6889 280.613
R13123 GND.n6890 GND.n942 280.613
R13124 GND.n6898 GND.n942 280.613
R13125 GND.n6899 GND.n6898 280.613
R13126 GND.n6900 GND.n6899 280.613
R13127 GND.n6900 GND.n936 280.613
R13128 GND.n6908 GND.n936 280.613
R13129 GND.n6909 GND.n6908 280.613
R13130 GND.n6910 GND.n6909 280.613
R13131 GND.n6910 GND.n930 280.613
R13132 GND.n6918 GND.n930 280.613
R13133 GND.n6919 GND.n6918 280.613
R13134 GND.n6920 GND.n6919 280.613
R13135 GND.n6920 GND.n924 280.613
R13136 GND.n6928 GND.n924 280.613
R13137 GND.n6929 GND.n6928 280.613
R13138 GND.n6930 GND.n6929 280.613
R13139 GND.n6930 GND.n918 280.613
R13140 GND.n6938 GND.n918 280.613
R13141 GND.n6939 GND.n6938 280.613
R13142 GND.n6940 GND.n6939 280.613
R13143 GND.n6940 GND.n912 280.613
R13144 GND.n6948 GND.n912 280.613
R13145 GND.n6949 GND.n6948 280.613
R13146 GND.n6950 GND.n6949 280.613
R13147 GND.n6950 GND.n906 280.613
R13148 GND.n6958 GND.n906 280.613
R13149 GND.n6959 GND.n6958 280.613
R13150 GND.n6960 GND.n6959 280.613
R13151 GND.n6960 GND.n900 280.613
R13152 GND.n6968 GND.n900 280.613
R13153 GND.n6969 GND.n6968 280.613
R13154 GND.n6970 GND.n6969 280.613
R13155 GND.n6970 GND.n894 280.613
R13156 GND.n6978 GND.n894 280.613
R13157 GND.n6979 GND.n6978 280.613
R13158 GND.n6980 GND.n6979 280.613
R13159 GND.n6980 GND.n888 280.613
R13160 GND.n6988 GND.n888 280.613
R13161 GND.n6989 GND.n6988 280.613
R13162 GND.n6990 GND.n6989 280.613
R13163 GND.n6990 GND.n882 280.613
R13164 GND.n6998 GND.n882 280.613
R13165 GND.n6999 GND.n6998 280.613
R13166 GND.n7000 GND.n6999 280.613
R13167 GND.n7000 GND.n876 280.613
R13168 GND.n7008 GND.n876 280.613
R13169 GND.n7009 GND.n7008 280.613
R13170 GND.n7010 GND.n7009 280.613
R13171 GND.n7010 GND.n870 280.613
R13172 GND.n7018 GND.n870 280.613
R13173 GND.n7019 GND.n7018 280.613
R13174 GND.n7020 GND.n7019 280.613
R13175 GND.n7020 GND.n864 280.613
R13176 GND.n7028 GND.n864 280.613
R13177 GND.n7029 GND.n7028 280.613
R13178 GND.n7030 GND.n7029 280.613
R13179 GND.n7030 GND.n858 280.613
R13180 GND.n7038 GND.n858 280.613
R13181 GND.n7039 GND.n7038 280.613
R13182 GND.n7040 GND.n7039 280.613
R13183 GND.n7040 GND.n852 280.613
R13184 GND.n7048 GND.n852 280.613
R13185 GND.n7049 GND.n7048 280.613
R13186 GND.n7050 GND.n7049 280.613
R13187 GND.n7050 GND.n846 280.613
R13188 GND.n7058 GND.n846 280.613
R13189 GND.n7059 GND.n7058 280.613
R13190 GND.n7060 GND.n7059 280.613
R13191 GND.n7060 GND.n840 280.613
R13192 GND.n7068 GND.n840 280.613
R13193 GND.n7069 GND.n7068 280.613
R13194 GND.n7070 GND.n7069 280.613
R13195 GND.n7070 GND.n834 280.613
R13196 GND.n7078 GND.n834 280.613
R13197 GND.n7079 GND.n7078 280.613
R13198 GND.n7080 GND.n7079 280.613
R13199 GND.n7080 GND.n828 280.613
R13200 GND.n7088 GND.n828 280.613
R13201 GND.n7089 GND.n7088 280.613
R13202 GND.n7090 GND.n7089 280.613
R13203 GND.n7090 GND.n822 280.613
R13204 GND.n7098 GND.n822 280.613
R13205 GND.n7099 GND.n7098 280.613
R13206 GND.n7100 GND.n7099 280.613
R13207 GND.n7100 GND.n816 280.613
R13208 GND.n7108 GND.n816 280.613
R13209 GND.n7109 GND.n7108 280.613
R13210 GND.n7110 GND.n7109 280.613
R13211 GND.n7110 GND.n810 280.613
R13212 GND.n7118 GND.n810 280.613
R13213 GND.n7119 GND.n7118 280.613
R13214 GND.n7120 GND.n7119 280.613
R13215 GND.n7120 GND.n804 280.613
R13216 GND.n7128 GND.n804 280.613
R13217 GND.n7129 GND.n7128 280.613
R13218 GND.n7130 GND.n7129 280.613
R13219 GND.n7130 GND.n798 280.613
R13220 GND.n7138 GND.n798 280.613
R13221 GND.n7139 GND.n7138 280.613
R13222 GND.n7140 GND.n7139 280.613
R13223 GND.n7140 GND.n792 280.613
R13224 GND.n7148 GND.n792 280.613
R13225 GND.n7149 GND.n7148 280.613
R13226 GND.n7150 GND.n7149 280.613
R13227 GND.n7150 GND.n786 280.613
R13228 GND.n7158 GND.n786 280.613
R13229 GND.n7159 GND.n7158 280.613
R13230 GND.n7160 GND.n7159 280.613
R13231 GND.n7160 GND.n780 280.613
R13232 GND.n7168 GND.n780 280.613
R13233 GND.n7169 GND.n7168 280.613
R13234 GND.n7170 GND.n7169 280.613
R13235 GND.n7170 GND.n774 280.613
R13236 GND.n7178 GND.n774 280.613
R13237 GND.n7179 GND.n7178 280.613
R13238 GND.n7180 GND.n7179 280.613
R13239 GND.n7180 GND.n768 280.613
R13240 GND.n7188 GND.n768 280.613
R13241 GND.n7189 GND.n7188 280.613
R13242 GND.n7190 GND.n7189 280.613
R13243 GND.n7190 GND.n762 280.613
R13244 GND.n7198 GND.n762 280.613
R13245 GND.n7199 GND.n7198 280.613
R13246 GND.n7200 GND.n7199 280.613
R13247 GND.n7200 GND.n756 280.613
R13248 GND.n7208 GND.n756 280.613
R13249 GND.n7209 GND.n7208 280.613
R13250 GND.n7210 GND.n7209 280.613
R13251 GND.n7210 GND.n750 280.613
R13252 GND.n7218 GND.n750 280.613
R13253 GND.n7219 GND.n7218 280.613
R13254 GND.n7220 GND.n7219 280.613
R13255 GND.n7220 GND.n744 280.613
R13256 GND.n7228 GND.n744 280.613
R13257 GND.n7229 GND.n7228 280.613
R13258 GND.n7230 GND.n7229 280.613
R13259 GND.n7230 GND.n738 280.613
R13260 GND.n7238 GND.n738 280.613
R13261 GND.n7239 GND.n7238 280.613
R13262 GND.n7240 GND.n7239 280.613
R13263 GND.n7240 GND.n732 280.613
R13264 GND.n7248 GND.n732 280.613
R13265 GND.n7249 GND.n7248 280.613
R13266 GND.n7250 GND.n7249 280.613
R13267 GND.n7250 GND.n726 280.613
R13268 GND.n7258 GND.n726 280.613
R13269 GND.n7259 GND.n7258 280.613
R13270 GND.n7260 GND.n7259 280.613
R13271 GND.n7260 GND.n720 280.613
R13272 GND.n7268 GND.n720 280.613
R13273 GND.n7269 GND.n7268 280.613
R13274 GND.n7270 GND.n7269 280.613
R13275 GND.n7270 GND.n714 280.613
R13276 GND.n7278 GND.n714 280.613
R13277 GND.n7279 GND.n7278 280.613
R13278 GND.n7280 GND.n7279 280.613
R13279 GND.n7280 GND.n708 280.613
R13280 GND.n7288 GND.n708 280.613
R13281 GND.n7289 GND.n7288 280.613
R13282 GND.n7290 GND.n7289 280.613
R13283 GND.n7290 GND.n702 280.613
R13284 GND.n7298 GND.n702 280.613
R13285 GND.n7299 GND.n7298 280.613
R13286 GND.n7300 GND.n7299 280.613
R13287 GND.n7300 GND.n696 280.613
R13288 GND.n7308 GND.n696 280.613
R13289 GND.n7309 GND.n7308 280.613
R13290 GND.n7310 GND.n7309 280.613
R13291 GND.n7310 GND.n690 280.613
R13292 GND.n7318 GND.n690 280.613
R13293 GND.n7319 GND.n7318 280.613
R13294 GND.n7320 GND.n7319 280.613
R13295 GND.n7320 GND.n684 280.613
R13296 GND.n7329 GND.n684 280.613
R13297 GND.n7330 GND.n7329 280.613
R13298 GND.n7331 GND.n7330 280.613
R13299 GND.n7331 GND.n679 280.613
R13300 GND.n1859 GND.t80 260.649
R13301 GND.n2486 GND.t136 260.649
R13302 GND.n5847 GND.n5846 256.663
R13303 GND.n5847 GND.n1828 256.663
R13304 GND.n5847 GND.n1829 256.663
R13305 GND.n5847 GND.n1830 256.663
R13306 GND.n5847 GND.n1831 256.663
R13307 GND.n5847 GND.n1832 256.663
R13308 GND.n5847 GND.n1833 256.663
R13309 GND.n5847 GND.n1834 256.663
R13310 GND.n5847 GND.n1835 256.663
R13311 GND.n5848 GND.n5847 256.663
R13312 GND.n5851 GND.n1824 256.663
R13313 GND.n5847 GND.n1836 256.663
R13314 GND.n5847 GND.n1837 256.663
R13315 GND.n5847 GND.n1838 256.663
R13316 GND.n5847 GND.n1839 256.663
R13317 GND.n5847 GND.n1840 256.663
R13318 GND.n5847 GND.n1841 256.663
R13319 GND.n5847 GND.n1842 256.663
R13320 GND.n5847 GND.n1843 256.663
R13321 GND.n5847 GND.n1844 256.663
R13322 GND.n5847 GND.n1845 256.663
R13323 GND.n5450 GND.n2454 256.663
R13324 GND.n5450 GND.n2453 256.663
R13325 GND.n5450 GND.n2452 256.663
R13326 GND.n5450 GND.n2451 256.663
R13327 GND.n5450 GND.n2450 256.663
R13328 GND.n5450 GND.n2449 256.663
R13329 GND.n5450 GND.n2448 256.663
R13330 GND.n5450 GND.n2447 256.663
R13331 GND.n5450 GND.n2446 256.663
R13332 GND.n5450 GND.n2445 256.663
R13333 GND.n5409 GND.n2548 256.663
R13334 GND.n5450 GND.n2455 256.663
R13335 GND.n5450 GND.n2456 256.663
R13336 GND.n5450 GND.n2457 256.663
R13337 GND.n5450 GND.n2458 256.663
R13338 GND.n5450 GND.n2459 256.663
R13339 GND.n5450 GND.n2460 256.663
R13340 GND.n5450 GND.n2461 256.663
R13341 GND.n5450 GND.n2462 256.663
R13342 GND.n5450 GND.n2463 256.663
R13343 GND.n5450 GND.n2464 256.663
R13344 GND.n5404 GND.n2581 242.672
R13345 GND.n5404 GND.n2582 242.672
R13346 GND.n5404 GND.n2583 242.672
R13347 GND.n5404 GND.n2584 242.672
R13348 GND.n5404 GND.n2585 242.672
R13349 GND.n5404 GND.n2586 242.672
R13350 GND.n5151 GND.n379 242.672
R13351 GND.n5115 GND.n379 242.672
R13352 GND.n5141 GND.n379 242.672
R13353 GND.n5119 GND.n379 242.672
R13354 GND.n5131 GND.n379 242.672
R13355 GND.n5123 GND.n379 242.672
R13356 GND.n4247 GND.n1896 242.672
R13357 GND.n3084 GND.n1896 242.672
R13358 GND.n4240 GND.n1896 242.672
R13359 GND.n4234 GND.n1896 242.672
R13360 GND.n4232 GND.n1896 242.672
R13361 GND.n4153 GND.n1896 242.672
R13362 GND.n4164 GND.n1896 242.672
R13363 GND.n4167 GND.n1896 242.672
R13364 GND.n4176 GND.n1896 242.672
R13365 GND.n4185 GND.n1896 242.672
R13366 GND.n4187 GND.n1896 242.672
R13367 GND.n5521 GND.n2379 242.672
R13368 GND.n5521 GND.n2380 242.672
R13369 GND.n5521 GND.n2381 242.672
R13370 GND.n5521 GND.n2382 242.672
R13371 GND.n5521 GND.n2383 242.672
R13372 GND.n5521 GND.n2384 242.672
R13373 GND.n5521 GND.n2385 242.672
R13374 GND.n5521 GND.n2386 242.672
R13375 GND.n5521 GND.n2387 242.672
R13376 GND.n5521 GND.n2388 242.672
R13377 GND.n5521 GND.n5520 242.672
R13378 GND.n6004 GND.n1615 242.672
R13379 GND.n6004 GND.n1616 242.672
R13380 GND.n6004 GND.n1617 242.672
R13381 GND.n6004 GND.n1618 242.672
R13382 GND.n6004 GND.n1619 242.672
R13383 GND.n6004 GND.n1620 242.672
R13384 GND.n6004 GND.n1621 242.672
R13385 GND.n6004 GND.n1622 242.672
R13386 GND.n6004 GND.n1623 242.672
R13387 GND.n6004 GND.n1624 242.672
R13388 GND.n6004 GND.n1625 242.672
R13389 GND.n6004 GND.n1626 242.672
R13390 GND.n6004 GND.n1627 242.672
R13391 GND.n6004 GND.n1628 242.672
R13392 GND.n6004 GND.n1629 242.672
R13393 GND.n6004 GND.n1630 242.672
R13394 GND.n6004 GND.n1631 242.672
R13395 GND.n6004 GND.n1632 242.672
R13396 GND.n6004 GND.n1633 242.672
R13397 GND.n6004 GND.n1634 242.672
R13398 GND.n6004 GND.n1635 242.672
R13399 GND.n6004 GND.n1636 242.672
R13400 GND.n6004 GND.n1637 242.672
R13401 GND.n6004 GND.n1638 242.672
R13402 GND.n6004 GND.n1639 242.672
R13403 GND.n5889 GND.n1757 242.672
R13404 GND.n5889 GND.n1758 242.672
R13405 GND.n5889 GND.n1759 242.672
R13406 GND.n5889 GND.n1760 242.672
R13407 GND.n5889 GND.n1761 242.672
R13408 GND.n5889 GND.n1762 242.672
R13409 GND.n5889 GND.n1763 242.672
R13410 GND.n5889 GND.n1764 242.672
R13411 GND.n5889 GND.n1765 242.672
R13412 GND.n5889 GND.n1766 242.672
R13413 GND.n5889 GND.n1767 242.672
R13414 GND.n5889 GND.n1768 242.672
R13415 GND.n5889 GND.n1769 242.672
R13416 GND.n5889 GND.n1770 242.672
R13417 GND.n5852 GND.n1822 242.672
R13418 GND.n5889 GND.n1771 242.672
R13419 GND.n5889 GND.n1772 242.672
R13420 GND.n5889 GND.n1773 242.672
R13421 GND.n5889 GND.n1774 242.672
R13422 GND.n5889 GND.n1775 242.672
R13423 GND.n5889 GND.n1776 242.672
R13424 GND.n5889 GND.n1777 242.672
R13425 GND.n5889 GND.n1778 242.672
R13426 GND.n5889 GND.n1779 242.672
R13427 GND.n5889 GND.n1780 242.672
R13428 GND.n5889 GND.n1781 242.672
R13429 GND.n5404 GND.n5403 242.672
R13430 GND.n5404 GND.n2558 242.672
R13431 GND.n5404 GND.n2559 242.672
R13432 GND.n5404 GND.n2560 242.672
R13433 GND.n5404 GND.n2561 242.672
R13434 GND.n5404 GND.n2562 242.672
R13435 GND.n5404 GND.n2563 242.672
R13436 GND.n5404 GND.n2564 242.672
R13437 GND.n5404 GND.n2565 242.672
R13438 GND.n5404 GND.n2566 242.672
R13439 GND.n5404 GND.n2567 242.672
R13440 GND.n5408 GND.n2550 242.672
R13441 GND.n5405 GND.n5404 242.672
R13442 GND.n5404 GND.n2568 242.672
R13443 GND.n5404 GND.n2569 242.672
R13444 GND.n5404 GND.n2570 242.672
R13445 GND.n5404 GND.n2571 242.672
R13446 GND.n5404 GND.n2572 242.672
R13447 GND.n5404 GND.n2573 242.672
R13448 GND.n5404 GND.n2574 242.672
R13449 GND.n5404 GND.n2575 242.672
R13450 GND.n5404 GND.n2576 242.672
R13451 GND.n5404 GND.n2577 242.672
R13452 GND.n5404 GND.n2578 242.672
R13453 GND.n5404 GND.n2579 242.672
R13454 GND.n5404 GND.n2580 242.672
R13455 GND.n379 GND.n191 242.672
R13456 GND.n379 GND.n192 242.672
R13457 GND.n379 GND.n193 242.672
R13458 GND.n379 GND.n194 242.672
R13459 GND.n379 GND.n195 242.672
R13460 GND.n379 GND.n196 242.672
R13461 GND.n379 GND.n197 242.672
R13462 GND.n379 GND.n198 242.672
R13463 GND.n379 GND.n199 242.672
R13464 GND.n379 GND.n200 242.672
R13465 GND.n379 GND.n201 242.672
R13466 GND.n379 GND.n202 242.672
R13467 GND.n379 GND.n203 242.672
R13468 GND.n379 GND.n204 242.672
R13469 GND.n379 GND.n205 242.672
R13470 GND.n379 GND.n206 242.672
R13471 GND.n379 GND.n207 242.672
R13472 GND.n379 GND.n208 242.672
R13473 GND.n379 GND.n209 242.672
R13474 GND.n379 GND.n210 242.672
R13475 GND.n379 GND.n211 242.672
R13476 GND.n379 GND.n212 242.672
R13477 GND.n379 GND.n213 242.672
R13478 GND.n379 GND.n214 242.672
R13479 GND.n379 GND.n215 242.672
R13480 GND.n6004 GND.n1641 242.672
R13481 GND.n6004 GND.n1642 242.672
R13482 GND.n6004 GND.n1643 242.672
R13483 GND.n6004 GND.n1644 242.672
R13484 GND.n6004 GND.n1645 242.672
R13485 GND.n5890 GND.n5889 242.672
R13486 GND.n5889 GND.n1755 242.672
R13487 GND.n5889 GND.n1754 242.672
R13488 GND.n5889 GND.n1753 242.672
R13489 GND.n5889 GND.n1752 242.672
R13490 GND.n5889 GND.n1751 242.672
R13491 GND.n378 GND.n216 240.244
R13492 GND.n371 GND.n370 240.244
R13493 GND.n368 GND.n367 240.244
R13494 GND.n364 GND.n363 240.244
R13495 GND.n360 GND.n359 240.244
R13496 GND.n356 GND.n355 240.244
R13497 GND.n352 GND.n351 240.244
R13498 GND.n348 GND.n347 240.244
R13499 GND.n344 GND.n343 240.244
R13500 GND.n340 GND.n339 240.244
R13501 GND.n336 GND.n335 240.244
R13502 GND.n332 GND.n331 240.244
R13503 GND.n325 GND.n324 240.244
R13504 GND.n321 GND.n320 240.244
R13505 GND.n317 GND.n316 240.244
R13506 GND.n313 GND.n312 240.244
R13507 GND.n309 GND.n308 240.244
R13508 GND.n305 GND.n304 240.244
R13509 GND.n259 GND.n258 240.244
R13510 GND.n297 GND.n296 240.244
R13511 GND.n293 GND.n292 240.244
R13512 GND.n289 GND.n288 240.244
R13513 GND.n285 GND.n284 240.244
R13514 GND.n281 GND.n280 240.244
R13515 GND.n277 GND.n276 240.244
R13516 GND.n4908 GND.n2595 240.244
R13517 GND.n5326 GND.n2595 240.244
R13518 GND.n5326 GND.n2606 240.244
R13519 GND.n4922 GND.n2606 240.244
R13520 GND.n4922 GND.n2619 240.244
R13521 GND.n4934 GND.n2619 240.244
R13522 GND.n4934 GND.n2637 240.244
R13523 GND.n4944 GND.n2637 240.244
R13524 GND.n4944 GND.n2648 240.244
R13525 GND.n4949 GND.n2648 240.244
R13526 GND.n4949 GND.n2659 240.244
R13527 GND.n4959 GND.n2659 240.244
R13528 GND.n4959 GND.n2669 240.244
R13529 GND.n4964 GND.n2669 240.244
R13530 GND.n4964 GND.n2680 240.244
R13531 GND.n4974 GND.n2680 240.244
R13532 GND.n4974 GND.n2690 240.244
R13533 GND.n4979 GND.n2690 240.244
R13534 GND.n4979 GND.n2701 240.244
R13535 GND.n4989 GND.n2701 240.244
R13536 GND.n4989 GND.n2711 240.244
R13537 GND.n4994 GND.n2711 240.244
R13538 GND.n4994 GND.n2722 240.244
R13539 GND.n5014 GND.n2722 240.244
R13540 GND.n5014 GND.n2731 240.244
R13541 GND.n2736 GND.n2731 240.244
R13542 GND.n5023 GND.n2736 240.244
R13543 GND.n5024 GND.n5023 240.244
R13544 GND.n5024 GND.n2748 240.244
R13545 GND.n2748 GND.n29 240.244
R13546 GND.n2756 GND.n29 240.244
R13547 GND.n5032 GND.n2756 240.244
R13548 GND.n5041 GND.n5032 240.244
R13549 GND.n5041 GND.n48 240.244
R13550 GND.n5045 GND.n48 240.244
R13551 GND.n5045 GND.n59 240.244
R13552 GND.n5056 GND.n59 240.244
R13553 GND.n5056 GND.n69 240.244
R13554 GND.n5060 GND.n69 240.244
R13555 GND.n5060 GND.n79 240.244
R13556 GND.n5070 GND.n79 240.244
R13557 GND.n5070 GND.n90 240.244
R13558 GND.n5074 GND.n90 240.244
R13559 GND.n5074 GND.n100 240.244
R13560 GND.n5084 GND.n100 240.244
R13561 GND.n5084 GND.n111 240.244
R13562 GND.n5088 GND.n111 240.244
R13563 GND.n5088 GND.n121 240.244
R13564 GND.n5099 GND.n121 240.244
R13565 GND.n5099 GND.n132 240.244
R13566 GND.n2787 GND.n132 240.244
R13567 GND.n2787 GND.n141 240.244
R13568 GND.n5172 GND.n141 240.244
R13569 GND.n5172 GND.n152 240.244
R13570 GND.n5168 GND.n152 240.244
R13571 GND.n5168 GND.n162 240.244
R13572 GND.n5160 GND.n162 240.244
R13573 GND.n5160 GND.n173 240.244
R13574 GND.n7739 GND.n173 240.244
R13575 GND.n2589 GND.n2588 240.244
R13576 GND.n5397 GND.n2588 240.244
R13577 GND.n5395 GND.n5394 240.244
R13578 GND.n5391 GND.n5390 240.244
R13579 GND.n5387 GND.n5386 240.244
R13580 GND.n5383 GND.n5382 240.244
R13581 GND.n5379 GND.n5378 240.244
R13582 GND.n5375 GND.n5374 240.244
R13583 GND.n5371 GND.n5370 240.244
R13584 GND.n5367 GND.n5366 240.244
R13585 GND.n5363 GND.n5362 240.244
R13586 GND.n5406 GND.n2556 240.244
R13587 GND.n4844 GND.n4843 240.244
R13588 GND.n4847 GND.n4846 240.244
R13589 GND.n4854 GND.n4853 240.244
R13590 GND.n4857 GND.n4856 240.244
R13591 GND.n4864 GND.n4863 240.244
R13592 GND.n4867 GND.n4866 240.244
R13593 GND.n4876 GND.n4875 240.244
R13594 GND.n4879 GND.n4878 240.244
R13595 GND.n4886 GND.n4885 240.244
R13596 GND.n4889 GND.n4888 240.244
R13597 GND.n4896 GND.n4895 240.244
R13598 GND.n4899 GND.n4898 240.244
R13599 GND.n5333 GND.n2590 240.244
R13600 GND.n5333 GND.n2593 240.244
R13601 GND.n2627 GND.n2593 240.244
R13602 GND.n2627 GND.n2623 240.244
R13603 GND.n5316 GND.n2623 240.244
R13604 GND.n5316 GND.n2624 240.244
R13605 GND.n5312 GND.n2624 240.244
R13606 GND.n5312 GND.n2635 240.244
R13607 GND.n5304 GND.n2635 240.244
R13608 GND.n5304 GND.n2651 240.244
R13609 GND.n5300 GND.n2651 240.244
R13610 GND.n5300 GND.n2657 240.244
R13611 GND.n5292 GND.n2657 240.244
R13612 GND.n5292 GND.n2672 240.244
R13613 GND.n5288 GND.n2672 240.244
R13614 GND.n5288 GND.n2678 240.244
R13615 GND.n5280 GND.n2678 240.244
R13616 GND.n5280 GND.n2693 240.244
R13617 GND.n5276 GND.n2693 240.244
R13618 GND.n5276 GND.n2699 240.244
R13619 GND.n5268 GND.n2699 240.244
R13620 GND.n5268 GND.n2714 240.244
R13621 GND.n5264 GND.n2714 240.244
R13622 GND.n5264 GND.n2720 240.244
R13623 GND.n5256 GND.n2720 240.244
R13624 GND.n5256 GND.n5254 240.244
R13625 GND.n5254 GND.n2734 240.244
R13626 GND.n2746 GND.n2734 240.244
R13627 GND.n2746 GND.n32 240.244
R13628 GND.n7823 GND.n32 240.244
R13629 GND.n7823 GND.n33 240.244
R13630 GND.n2758 GND.n33 240.244
R13631 GND.n2758 GND.n45 240.244
R13632 GND.n7818 GND.n45 240.244
R13633 GND.n7818 GND.n46 240.244
R13634 GND.n7810 GND.n46 240.244
R13635 GND.n7810 GND.n62 240.244
R13636 GND.n7806 GND.n62 240.244
R13637 GND.n7806 GND.n67 240.244
R13638 GND.n7798 GND.n67 240.244
R13639 GND.n7798 GND.n82 240.244
R13640 GND.n7794 GND.n82 240.244
R13641 GND.n7794 GND.n88 240.244
R13642 GND.n7786 GND.n88 240.244
R13643 GND.n7786 GND.n103 240.244
R13644 GND.n7782 GND.n103 240.244
R13645 GND.n7782 GND.n109 240.244
R13646 GND.n7774 GND.n109 240.244
R13647 GND.n7774 GND.n124 240.244
R13648 GND.n7770 GND.n124 240.244
R13649 GND.n7770 GND.n130 240.244
R13650 GND.n7762 GND.n130 240.244
R13651 GND.n7762 GND.n144 240.244
R13652 GND.n7758 GND.n144 240.244
R13653 GND.n7758 GND.n150 240.244
R13654 GND.n7750 GND.n150 240.244
R13655 GND.n7750 GND.n165 240.244
R13656 GND.n7746 GND.n165 240.244
R13657 GND.n7746 GND.n171 240.244
R13658 GND.n5888 GND.n1783 240.244
R13659 GND.n1788 GND.n1787 240.244
R13660 GND.n1790 GND.n1789 240.244
R13661 GND.n1794 GND.n1793 240.244
R13662 GND.n1796 GND.n1795 240.244
R13663 GND.n1802 GND.n1799 240.244
R13664 GND.n1804 GND.n1803 240.244
R13665 GND.n1808 GND.n1807 240.244
R13666 GND.n1810 GND.n1809 240.244
R13667 GND.n1814 GND.n1813 240.244
R13668 GND.n1816 GND.n1815 240.244
R13669 GND.n3131 GND.n3130 240.244
R13670 GND.n3136 GND.n3135 240.244
R13671 GND.n3128 GND.n3127 240.244
R13672 GND.n3144 GND.n3143 240.244
R13673 GND.n3124 GND.n3123 240.244
R13674 GND.n3152 GND.n3151 240.244
R13675 GND.n3120 GND.n3119 240.244
R13676 GND.n3160 GND.n3159 240.244
R13677 GND.n3114 GND.n3113 240.244
R13678 GND.n3168 GND.n3167 240.244
R13679 GND.n3110 GND.n3109 240.244
R13680 GND.n3176 GND.n3175 240.244
R13681 GND.n3182 GND.n3181 240.244
R13682 GND.n3667 GND.n3492 240.244
R13683 GND.n3492 GND.n3476 240.244
R13684 GND.n3476 GND.n3466 240.244
R13685 GND.n3692 GND.n3466 240.244
R13686 GND.n3692 GND.n3457 240.244
R13687 GND.n3694 GND.n3457 240.244
R13688 GND.n3694 GND.n3446 240.244
R13689 GND.n3446 GND.n3437 240.244
R13690 GND.n3729 GND.n3437 240.244
R13691 GND.n3729 GND.n3428 240.244
R13692 GND.n3731 GND.n3428 240.244
R13693 GND.n3731 GND.n3418 240.244
R13694 GND.n3418 GND.n3408 240.244
R13695 GND.n3766 GND.n3408 240.244
R13696 GND.n3766 GND.n3398 240.244
R13697 GND.n3768 GND.n3398 240.244
R13698 GND.n3768 GND.n3388 240.244
R13699 GND.n3388 GND.n3379 240.244
R13700 GND.n3810 GND.n3379 240.244
R13701 GND.n3810 GND.n3368 240.244
R13702 GND.n3368 GND.n3359 240.244
R13703 GND.n3827 GND.n3359 240.244
R13704 GND.n3828 GND.n3827 240.244
R13705 GND.n3828 GND.n3336 240.244
R13706 GND.n3837 GND.n3336 240.244
R13707 GND.n3837 GND.n3346 240.244
R13708 GND.n3839 GND.n3346 240.244
R13709 GND.n3840 GND.n3839 240.244
R13710 GND.n3866 GND.n3840 240.244
R13711 GND.n3866 GND.n3846 240.244
R13712 GND.n3847 GND.n3846 240.244
R13713 GND.n3848 GND.n3847 240.244
R13714 GND.n3858 GND.n3848 240.244
R13715 GND.n3858 GND.n3320 240.244
R13716 GND.n3949 GND.n3320 240.244
R13717 GND.n3949 GND.n3311 240.244
R13718 GND.n3951 GND.n3311 240.244
R13719 GND.n3951 GND.n3302 240.244
R13720 GND.n3302 GND.n3292 240.244
R13721 GND.n3986 GND.n3292 240.244
R13722 GND.n3986 GND.n3283 240.244
R13723 GND.n3988 GND.n3283 240.244
R13724 GND.n3988 GND.n3272 240.244
R13725 GND.n3272 GND.n3263 240.244
R13726 GND.n4023 GND.n3263 240.244
R13727 GND.n4023 GND.n3254 240.244
R13728 GND.n4025 GND.n3254 240.244
R13729 GND.n4025 GND.n3244 240.244
R13730 GND.n3244 GND.n3234 240.244
R13731 GND.n4060 GND.n3234 240.244
R13732 GND.n4060 GND.n3224 240.244
R13733 GND.n4062 GND.n3224 240.244
R13734 GND.n4062 GND.n3214 240.244
R13735 GND.n3214 GND.n3205 240.244
R13736 GND.n4131 GND.n3205 240.244
R13737 GND.n4131 GND.n3197 240.244
R13738 GND.n4134 GND.n3197 240.244
R13739 GND.n4134 GND.n3103 240.244
R13740 GND.n4224 GND.n3103 240.244
R13741 GND.n3530 GND.n3529 240.244
R13742 GND.n3536 GND.n3535 240.244
R13743 GND.n3540 GND.n3539 240.244
R13744 GND.n3546 GND.n3545 240.244
R13745 GND.n3550 GND.n3549 240.244
R13746 GND.n3556 GND.n3555 240.244
R13747 GND.n3559 GND.n3558 240.244
R13748 GND.n3566 GND.n3565 240.244
R13749 GND.n3569 GND.n3568 240.244
R13750 GND.n3576 GND.n3575 240.244
R13751 GND.n3579 GND.n3578 240.244
R13752 GND.n3586 GND.n3585 240.244
R13753 GND.n3590 GND.n3589 240.244
R13754 GND.n3596 GND.n3595 240.244
R13755 GND.n3600 GND.n3599 240.244
R13756 GND.n3606 GND.n3605 240.244
R13757 GND.n3610 GND.n3609 240.244
R13758 GND.n3503 GND.n3502 240.244
R13759 GND.n3620 GND.n3619 240.244
R13760 GND.n3626 GND.n3625 240.244
R13761 GND.n3630 GND.n3629 240.244
R13762 GND.n3636 GND.n3635 240.244
R13763 GND.n3640 GND.n3639 240.244
R13764 GND.n3646 GND.n3645 240.244
R13765 GND.n3648 GND.n1640 240.244
R13766 GND.n3670 GND.n3479 240.244
R13767 GND.n3678 GND.n3479 240.244
R13768 GND.n3678 GND.n3480 240.244
R13769 GND.n3480 GND.n3455 240.244
R13770 GND.n3707 GND.n3455 240.244
R13771 GND.n3707 GND.n3450 240.244
R13772 GND.n3715 GND.n3450 240.244
R13773 GND.n3715 GND.n3451 240.244
R13774 GND.n3451 GND.n3426 240.244
R13775 GND.n3744 GND.n3426 240.244
R13776 GND.n3744 GND.n3421 240.244
R13777 GND.n3752 GND.n3421 240.244
R13778 GND.n3752 GND.n3422 240.244
R13779 GND.n3422 GND.n3396 240.244
R13780 GND.n3781 GND.n3396 240.244
R13781 GND.n3781 GND.n3391 240.244
R13782 GND.n3789 GND.n3391 240.244
R13783 GND.n3789 GND.n3392 240.244
R13784 GND.n3392 GND.n3366 240.244
R13785 GND.n3818 GND.n3366 240.244
R13786 GND.n3818 GND.n3362 240.244
R13787 GND.n3825 GND.n3362 240.244
R13788 GND.n3825 GND.n3339 240.244
R13789 GND.n3936 GND.n3339 240.244
R13790 GND.n3936 GND.n3340 240.244
R13791 GND.n3931 GND.n3340 240.244
R13792 GND.n3931 GND.n3344 240.244
R13793 GND.n3880 GND.n3344 240.244
R13794 GND.n3887 GND.n3880 240.244
R13795 GND.n3887 GND.n3881 240.244
R13796 GND.n3881 GND.n3856 240.244
R13797 GND.n3906 GND.n3856 240.244
R13798 GND.n3906 GND.n3854 240.244
R13799 GND.n3911 GND.n3854 240.244
R13800 GND.n3911 GND.n3310 240.244
R13801 GND.n3964 GND.n3310 240.244
R13802 GND.n3964 GND.n3305 240.244
R13803 GND.n3972 GND.n3305 240.244
R13804 GND.n3972 GND.n3306 240.244
R13805 GND.n3306 GND.n3281 240.244
R13806 GND.n4001 GND.n3281 240.244
R13807 GND.n4001 GND.n3276 240.244
R13808 GND.n4009 GND.n3276 240.244
R13809 GND.n4009 GND.n3277 240.244
R13810 GND.n3277 GND.n3252 240.244
R13811 GND.n4038 GND.n3252 240.244
R13812 GND.n4038 GND.n3247 240.244
R13813 GND.n4046 GND.n3247 240.244
R13814 GND.n4046 GND.n3248 240.244
R13815 GND.n3248 GND.n3222 240.244
R13816 GND.n4075 GND.n3222 240.244
R13817 GND.n4075 GND.n3217 240.244
R13818 GND.n4083 GND.n3217 240.244
R13819 GND.n4083 GND.n3218 240.244
R13820 GND.n3218 GND.n3195 240.244
R13821 GND.n4141 GND.n3195 240.244
R13822 GND.n4141 GND.n3191 240.244
R13823 GND.n4148 GND.n3191 240.244
R13824 GND.n4148 GND.n1782 240.244
R13825 GND.n5522 GND.n2377 240.244
R13826 GND.n5519 GND.n2389 240.244
R13827 GND.n5515 GND.n5514 240.244
R13828 GND.n5511 GND.n5510 240.244
R13829 GND.n5507 GND.n5506 240.244
R13830 GND.n5503 GND.n5502 240.244
R13831 GND.n5499 GND.n5498 240.244
R13832 GND.n5495 GND.n5494 240.244
R13833 GND.n5491 GND.n5490 240.244
R13834 GND.n5487 GND.n5486 240.244
R13835 GND.n5483 GND.n5482 240.244
R13836 GND.n4260 GND.n4257 240.244
R13837 GND.n4260 GND.n1971 240.244
R13838 GND.n4271 GND.n1971 240.244
R13839 GND.n4271 GND.n1982 240.244
R13840 GND.n4267 GND.n1982 240.244
R13841 GND.n4267 GND.n3062 240.244
R13842 GND.n4298 GND.n3062 240.244
R13843 GND.n4298 GND.n2017 240.244
R13844 GND.n4319 GND.n2017 240.244
R13845 GND.n4319 GND.n2028 240.244
R13846 GND.n4315 GND.n2028 240.244
R13847 GND.n4315 GND.n4314 240.244
R13848 GND.n4314 GND.n4313 240.244
R13849 GND.n4313 GND.n4306 240.244
R13850 GND.n4306 GND.n2062 240.244
R13851 GND.n4418 GND.n2062 240.244
R13852 GND.n4418 GND.n2081 240.244
R13853 GND.n3044 GND.n2081 240.244
R13854 GND.n4425 GND.n3044 240.244
R13855 GND.n4426 GND.n4425 240.244
R13856 GND.n4427 GND.n4426 240.244
R13857 GND.n4427 GND.n3039 240.244
R13858 GND.n4441 GND.n3039 240.244
R13859 GND.n4441 GND.n3040 240.244
R13860 GND.n4437 GND.n3040 240.244
R13861 GND.n4437 GND.n3015 240.244
R13862 GND.n4461 GND.n3015 240.244
R13863 GND.n4462 GND.n4461 240.244
R13864 GND.n4463 GND.n4462 240.244
R13865 GND.n4463 GND.n3010 240.244
R13866 GND.n4486 GND.n3010 240.244
R13867 GND.n4486 GND.n3011 240.244
R13868 GND.n4482 GND.n3011 240.244
R13869 GND.n4482 GND.n4481 240.244
R13870 GND.n4481 GND.n3002 240.244
R13871 GND.n4476 GND.n3002 240.244
R13872 GND.n4476 GND.n4475 240.244
R13873 GND.n4475 GND.n2994 240.244
R13874 GND.n4535 GND.n2994 240.244
R13875 GND.n4535 GND.n2186 240.244
R13876 GND.n4543 GND.n2186 240.244
R13877 GND.n4543 GND.n2197 240.244
R13878 GND.n4562 GND.n2197 240.244
R13879 GND.n4563 GND.n4562 240.244
R13880 GND.n4563 GND.n2983 240.244
R13881 GND.n4569 GND.n2983 240.244
R13882 GND.n4570 GND.n4569 240.244
R13883 GND.n4571 GND.n4570 240.244
R13884 GND.n4571 GND.n2979 240.244
R13885 GND.n4630 GND.n2979 240.244
R13886 GND.n4631 GND.n4630 240.244
R13887 GND.n4632 GND.n4631 240.244
R13888 GND.n4632 GND.n2975 240.244
R13889 GND.n4639 GND.n2975 240.244
R13890 GND.n4639 GND.n2270 240.244
R13891 GND.n4675 GND.n2270 240.244
R13892 GND.n4675 GND.n2281 240.244
R13893 GND.n4678 GND.n2281 240.244
R13894 GND.n4678 GND.n2963 240.244
R13895 GND.n4684 GND.n2963 240.244
R13896 GND.n4684 GND.n2306 240.244
R13897 GND.n4695 GND.n2306 240.244
R13898 GND.n4695 GND.n2322 240.244
R13899 GND.n4701 GND.n2322 240.244
R13900 GND.n4701 GND.n2332 240.244
R13901 GND.n4739 GND.n2332 240.244
R13902 GND.n4739 GND.n2342 240.244
R13903 GND.n4751 GND.n2342 240.244
R13904 GND.n4751 GND.n2352 240.244
R13905 GND.n4747 GND.n2352 240.244
R13906 GND.n4747 GND.n2361 240.244
R13907 GND.n4793 GND.n2361 240.244
R13908 GND.n4793 GND.n2370 240.244
R13909 GND.n5478 GND.n2370 240.244
R13910 GND.n4248 GND.n4246 240.244
R13911 GND.n4246 GND.n4245 240.244
R13912 GND.n4242 GND.n4241 240.244
R13913 GND.n4239 GND.n3089 240.244
R13914 GND.n4235 GND.n4233 240.244
R13915 GND.n4231 GND.n3095 240.244
R13916 GND.n4155 GND.n4154 240.244
R13917 GND.n4166 GND.n4165 240.244
R13918 GND.n4175 GND.n4168 240.244
R13919 GND.n4178 GND.n4177 240.244
R13920 GND.n4188 GND.n4186 240.244
R13921 GND.n4255 GND.n1973 240.244
R13922 GND.n5777 GND.n1973 240.244
R13923 GND.n5777 GND.n1974 240.244
R13924 GND.n5773 GND.n1974 240.244
R13925 GND.n5773 GND.n1980 240.244
R13926 GND.n3068 GND.n1980 240.244
R13927 GND.n3068 GND.n2019 240.244
R13928 GND.n5756 GND.n2019 240.244
R13929 GND.n5756 GND.n2020 240.244
R13930 GND.n5752 GND.n2020 240.244
R13931 GND.n5752 GND.n2026 240.244
R13932 GND.n2070 GND.n2026 240.244
R13933 GND.n2071 GND.n2070 240.244
R13934 GND.n2071 GND.n2064 240.244
R13935 GND.n5729 GND.n2064 240.244
R13936 GND.n5729 GND.n2065 240.244
R13937 GND.n5725 GND.n2065 240.244
R13938 GND.n5725 GND.n2079 240.244
R13939 GND.n3030 GND.n2079 240.244
R13940 GND.n3031 GND.n3030 240.244
R13941 GND.n3032 GND.n3031 240.244
R13942 GND.n3032 GND.n3023 240.244
R13943 GND.n4443 GND.n3023 240.244
R13944 GND.n4444 GND.n4443 240.244
R13945 GND.n4445 GND.n4444 240.244
R13946 GND.n4445 GND.n3018 240.244
R13947 GND.n4459 GND.n3018 240.244
R13948 GND.n4459 GND.n3019 240.244
R13949 GND.n4455 GND.n3019 240.244
R13950 GND.n4455 GND.n3008 240.244
R13951 GND.n4488 GND.n3008 240.244
R13952 GND.n4489 GND.n4488 240.244
R13953 GND.n4490 GND.n4489 240.244
R13954 GND.n4490 GND.n3003 240.244
R13955 GND.n4505 GND.n3003 240.244
R13956 GND.n4505 GND.n3004 240.244
R13957 GND.n4501 GND.n3004 240.244
R13958 GND.n4501 GND.n4500 240.244
R13959 GND.n4500 GND.n2188 240.244
R13960 GND.n5645 GND.n2188 240.244
R13961 GND.n5645 GND.n2189 240.244
R13962 GND.n5641 GND.n2189 240.244
R13963 GND.n5641 GND.n2195 240.244
R13964 GND.n4604 GND.n2195 240.244
R13965 GND.n4604 GND.n4601 240.244
R13966 GND.n4610 GND.n4601 240.244
R13967 GND.n4611 GND.n4610 240.244
R13968 GND.n4612 GND.n4611 240.244
R13969 GND.n4612 GND.n4596 240.244
R13970 GND.n4628 GND.n4596 240.244
R13971 GND.n4628 GND.n4597 240.244
R13972 GND.n4624 GND.n4597 240.244
R13973 GND.n4624 GND.n4623 240.244
R13974 GND.n4623 GND.n2272 240.244
R13975 GND.n5591 GND.n2272 240.244
R13976 GND.n5591 GND.n2273 240.244
R13977 GND.n5587 GND.n2273 240.244
R13978 GND.n5587 GND.n2279 240.244
R13979 GND.n2312 GND.n2279 240.244
R13980 GND.n2312 GND.n2308 240.244
R13981 GND.n5570 GND.n2308 240.244
R13982 GND.n5570 GND.n2309 240.244
R13983 GND.n5566 GND.n2309 240.244
R13984 GND.n5566 GND.n2320 240.244
R13985 GND.n5556 GND.n2320 240.244
R13986 GND.n5556 GND.n2334 240.244
R13987 GND.n5552 GND.n2334 240.244
R13988 GND.n5552 GND.n2340 240.244
R13989 GND.n5542 GND.n2340 240.244
R13990 GND.n5542 GND.n2354 240.244
R13991 GND.n5538 GND.n2354 240.244
R13992 GND.n5538 GND.n2360 240.244
R13993 GND.n5528 GND.n2360 240.244
R13994 GND.n5528 GND.n2372 240.244
R13995 GND.n5130 GND.n5129 240.244
R13996 GND.n5133 GND.n5132 240.244
R13997 GND.n5140 GND.n5139 240.244
R13998 GND.n5143 GND.n5142 240.244
R13999 GND.n5150 GND.n5149 240.244
R14000 GND.n4910 GND.n2596 240.244
R14001 GND.n2607 GND.n2596 240.244
R14002 GND.n4917 GND.n2607 240.244
R14003 GND.n4918 GND.n4917 240.244
R14004 GND.n4918 GND.n2620 240.244
R14005 GND.n4936 GND.n2620 240.244
R14006 GND.n4936 GND.n2638 240.244
R14007 GND.n4942 GND.n2638 240.244
R14008 GND.n4942 GND.n2649 240.244
R14009 GND.n4951 GND.n2649 240.244
R14010 GND.n4951 GND.n2660 240.244
R14011 GND.n4957 GND.n2660 240.244
R14012 GND.n4957 GND.n2670 240.244
R14013 GND.n4966 GND.n2670 240.244
R14014 GND.n4966 GND.n2681 240.244
R14015 GND.n4972 GND.n2681 240.244
R14016 GND.n4972 GND.n2691 240.244
R14017 GND.n4981 GND.n2691 240.244
R14018 GND.n4981 GND.n2702 240.244
R14019 GND.n4987 GND.n2702 240.244
R14020 GND.n4987 GND.n2712 240.244
R14021 GND.n4996 GND.n2712 240.244
R14022 GND.n4996 GND.n2723 240.244
R14023 GND.n5012 GND.n2723 240.244
R14024 GND.n5012 GND.n2732 240.244
R14025 GND.n2737 GND.n2732 240.244
R14026 GND.n5007 GND.n2737 240.244
R14027 GND.n5007 GND.n5006 240.244
R14028 GND.n5006 GND.n26 240.244
R14029 GND.n7825 GND.n26 240.244
R14030 GND.n7825 GND.n27 240.244
R14031 GND.n5034 GND.n27 240.244
R14032 GND.n5039 GND.n5034 240.244
R14033 GND.n5039 GND.n49 240.244
R14034 GND.n5048 GND.n49 240.244
R14035 GND.n5048 GND.n60 240.244
R14036 GND.n5054 GND.n60 240.244
R14037 GND.n5054 GND.n70 240.244
R14038 GND.n5062 GND.n70 240.244
R14039 GND.n5062 GND.n80 240.244
R14040 GND.n5068 GND.n80 240.244
R14041 GND.n5068 GND.n91 240.244
R14042 GND.n5076 GND.n91 240.244
R14043 GND.n5076 GND.n101 240.244
R14044 GND.n5082 GND.n101 240.244
R14045 GND.n5082 GND.n112 240.244
R14046 GND.n5090 GND.n112 240.244
R14047 GND.n5090 GND.n122 240.244
R14048 GND.n5097 GND.n122 240.244
R14049 GND.n5097 GND.n133 240.244
R14050 GND.n5178 GND.n133 240.244
R14051 GND.n5178 GND.n142 240.244
R14052 GND.n5174 GND.n142 240.244
R14053 GND.n5174 GND.n153 240.244
R14054 GND.n5166 GND.n153 240.244
R14055 GND.n5166 GND.n163 240.244
R14056 GND.n5162 GND.n163 240.244
R14057 GND.n5162 GND.n174 240.244
R14058 GND.n181 GND.n174 240.244
R14059 GND.n2908 GND.n2907 240.244
R14060 GND.n2914 GND.n2913 240.244
R14061 GND.n2920 GND.n2919 240.244
R14062 GND.n2926 GND.n2925 240.244
R14063 GND.n2928 GND.n2897 240.244
R14064 GND.n5331 GND.n2598 240.244
R14065 GND.n5331 GND.n2599 240.244
R14066 GND.n4927 GND.n2599 240.244
R14067 GND.n4928 GND.n4927 240.244
R14068 GND.n4928 GND.n2622 240.244
R14069 GND.n2639 GND.n2622 240.244
R14070 GND.n5310 GND.n2639 240.244
R14071 GND.n5310 GND.n2640 240.244
R14072 GND.n5306 GND.n2640 240.244
R14073 GND.n5306 GND.n2646 240.244
R14074 GND.n5298 GND.n2646 240.244
R14075 GND.n5298 GND.n2662 240.244
R14076 GND.n5294 GND.n2662 240.244
R14077 GND.n5294 GND.n2667 240.244
R14078 GND.n5286 GND.n2667 240.244
R14079 GND.n5286 GND.n2683 240.244
R14080 GND.n5282 GND.n2683 240.244
R14081 GND.n5282 GND.n2688 240.244
R14082 GND.n5274 GND.n2688 240.244
R14083 GND.n5274 GND.n2704 240.244
R14084 GND.n5270 GND.n2704 240.244
R14085 GND.n5270 GND.n2709 240.244
R14086 GND.n5262 GND.n2709 240.244
R14087 GND.n5262 GND.n2724 240.244
R14088 GND.n5258 GND.n2724 240.244
R14089 GND.n5258 GND.n2729 240.244
R14090 GND.n5019 GND.n2729 240.244
R14091 GND.n5019 GND.n2749 240.244
R14092 GND.n5243 GND.n2749 240.244
R14093 GND.n5243 GND.n31 240.244
R14094 GND.n5239 GND.n31 240.244
R14095 GND.n5239 GND.n2755 240.244
R14096 GND.n2755 GND.n51 240.244
R14097 GND.n7816 GND.n51 240.244
R14098 GND.n7816 GND.n52 240.244
R14099 GND.n7812 GND.n52 240.244
R14100 GND.n7812 GND.n58 240.244
R14101 GND.n7804 GND.n58 240.244
R14102 GND.n7804 GND.n72 240.244
R14103 GND.n7800 GND.n72 240.244
R14104 GND.n7800 GND.n77 240.244
R14105 GND.n7792 GND.n77 240.244
R14106 GND.n7792 GND.n93 240.244
R14107 GND.n7788 GND.n93 240.244
R14108 GND.n7788 GND.n98 240.244
R14109 GND.n7780 GND.n98 240.244
R14110 GND.n7780 GND.n114 240.244
R14111 GND.n7776 GND.n114 240.244
R14112 GND.n7776 GND.n119 240.244
R14113 GND.n7768 GND.n119 240.244
R14114 GND.n7768 GND.n135 240.244
R14115 GND.n7764 GND.n135 240.244
R14116 GND.n7764 GND.n140 240.244
R14117 GND.n7756 GND.n140 240.244
R14118 GND.n7756 GND.n155 240.244
R14119 GND.n7752 GND.n155 240.244
R14120 GND.n7752 GND.n160 240.244
R14121 GND.n7744 GND.n160 240.244
R14122 GND.n7744 GND.n176 240.244
R14123 GND.n6357 GND.n1265 240.244
R14124 GND.n6361 GND.n1265 240.244
R14125 GND.n6361 GND.n1261 240.244
R14126 GND.n6367 GND.n1261 240.244
R14127 GND.n6367 GND.n1259 240.244
R14128 GND.n6371 GND.n1259 240.244
R14129 GND.n6371 GND.n1255 240.244
R14130 GND.n6377 GND.n1255 240.244
R14131 GND.n6377 GND.n1253 240.244
R14132 GND.n6381 GND.n1253 240.244
R14133 GND.n6381 GND.n1249 240.244
R14134 GND.n6387 GND.n1249 240.244
R14135 GND.n6387 GND.n1247 240.244
R14136 GND.n6391 GND.n1247 240.244
R14137 GND.n6391 GND.n1243 240.244
R14138 GND.n6397 GND.n1243 240.244
R14139 GND.n6397 GND.n1241 240.244
R14140 GND.n6401 GND.n1241 240.244
R14141 GND.n6401 GND.n1237 240.244
R14142 GND.n6407 GND.n1237 240.244
R14143 GND.n6407 GND.n1235 240.244
R14144 GND.n6411 GND.n1235 240.244
R14145 GND.n6411 GND.n1231 240.244
R14146 GND.n6417 GND.n1231 240.244
R14147 GND.n6417 GND.n1229 240.244
R14148 GND.n6421 GND.n1229 240.244
R14149 GND.n6421 GND.n1225 240.244
R14150 GND.n6427 GND.n1225 240.244
R14151 GND.n6427 GND.n1223 240.244
R14152 GND.n6431 GND.n1223 240.244
R14153 GND.n6431 GND.n1219 240.244
R14154 GND.n6437 GND.n1219 240.244
R14155 GND.n6437 GND.n1217 240.244
R14156 GND.n6441 GND.n1217 240.244
R14157 GND.n6441 GND.n1213 240.244
R14158 GND.n6447 GND.n1213 240.244
R14159 GND.n6447 GND.n1211 240.244
R14160 GND.n6451 GND.n1211 240.244
R14161 GND.n6451 GND.n1207 240.244
R14162 GND.n6457 GND.n1207 240.244
R14163 GND.n6457 GND.n1205 240.244
R14164 GND.n6461 GND.n1205 240.244
R14165 GND.n6461 GND.n1201 240.244
R14166 GND.n6467 GND.n1201 240.244
R14167 GND.n6467 GND.n1199 240.244
R14168 GND.n6471 GND.n1199 240.244
R14169 GND.n6471 GND.n1195 240.244
R14170 GND.n6477 GND.n1195 240.244
R14171 GND.n6477 GND.n1193 240.244
R14172 GND.n6481 GND.n1193 240.244
R14173 GND.n6481 GND.n1189 240.244
R14174 GND.n6487 GND.n1189 240.244
R14175 GND.n6487 GND.n1187 240.244
R14176 GND.n6491 GND.n1187 240.244
R14177 GND.n6491 GND.n1183 240.244
R14178 GND.n6497 GND.n1183 240.244
R14179 GND.n6497 GND.n1181 240.244
R14180 GND.n6501 GND.n1181 240.244
R14181 GND.n6501 GND.n1177 240.244
R14182 GND.n6507 GND.n1177 240.244
R14183 GND.n6507 GND.n1175 240.244
R14184 GND.n6511 GND.n1175 240.244
R14185 GND.n6511 GND.n1171 240.244
R14186 GND.n6517 GND.n1171 240.244
R14187 GND.n6517 GND.n1169 240.244
R14188 GND.n6521 GND.n1169 240.244
R14189 GND.n6521 GND.n1165 240.244
R14190 GND.n6527 GND.n1165 240.244
R14191 GND.n6527 GND.n1163 240.244
R14192 GND.n6531 GND.n1163 240.244
R14193 GND.n6531 GND.n1159 240.244
R14194 GND.n6537 GND.n1159 240.244
R14195 GND.n6537 GND.n1157 240.244
R14196 GND.n6541 GND.n1157 240.244
R14197 GND.n6541 GND.n1153 240.244
R14198 GND.n6547 GND.n1153 240.244
R14199 GND.n6547 GND.n1151 240.244
R14200 GND.n6551 GND.n1151 240.244
R14201 GND.n6551 GND.n1147 240.244
R14202 GND.n6557 GND.n1147 240.244
R14203 GND.n6557 GND.n1145 240.244
R14204 GND.n6561 GND.n1145 240.244
R14205 GND.n6561 GND.n1141 240.244
R14206 GND.n6567 GND.n1141 240.244
R14207 GND.n6567 GND.n1139 240.244
R14208 GND.n6571 GND.n1139 240.244
R14209 GND.n6571 GND.n1135 240.244
R14210 GND.n6577 GND.n1135 240.244
R14211 GND.n6577 GND.n1133 240.244
R14212 GND.n6581 GND.n1133 240.244
R14213 GND.n6581 GND.n1129 240.244
R14214 GND.n6587 GND.n1129 240.244
R14215 GND.n6587 GND.n1127 240.244
R14216 GND.n6591 GND.n1127 240.244
R14217 GND.n6591 GND.n1123 240.244
R14218 GND.n6597 GND.n1123 240.244
R14219 GND.n6597 GND.n1121 240.244
R14220 GND.n6601 GND.n1121 240.244
R14221 GND.n6601 GND.n1117 240.244
R14222 GND.n6607 GND.n1117 240.244
R14223 GND.n6607 GND.n1115 240.244
R14224 GND.n6611 GND.n1115 240.244
R14225 GND.n6611 GND.n1111 240.244
R14226 GND.n6617 GND.n1111 240.244
R14227 GND.n6617 GND.n1109 240.244
R14228 GND.n6621 GND.n1109 240.244
R14229 GND.n6621 GND.n1105 240.244
R14230 GND.n6627 GND.n1105 240.244
R14231 GND.n6627 GND.n1103 240.244
R14232 GND.n6631 GND.n1103 240.244
R14233 GND.n6631 GND.n1099 240.244
R14234 GND.n6637 GND.n1099 240.244
R14235 GND.n6637 GND.n1097 240.244
R14236 GND.n6641 GND.n1097 240.244
R14237 GND.n6641 GND.n1093 240.244
R14238 GND.n6647 GND.n1093 240.244
R14239 GND.n6647 GND.n1091 240.244
R14240 GND.n6651 GND.n1091 240.244
R14241 GND.n6651 GND.n1087 240.244
R14242 GND.n6657 GND.n1087 240.244
R14243 GND.n6657 GND.n1085 240.244
R14244 GND.n6661 GND.n1085 240.244
R14245 GND.n6661 GND.n1081 240.244
R14246 GND.n6667 GND.n1081 240.244
R14247 GND.n6667 GND.n1079 240.244
R14248 GND.n6671 GND.n1079 240.244
R14249 GND.n6671 GND.n1075 240.244
R14250 GND.n6677 GND.n1075 240.244
R14251 GND.n6677 GND.n1073 240.244
R14252 GND.n6681 GND.n1073 240.244
R14253 GND.n6681 GND.n1069 240.244
R14254 GND.n6687 GND.n1069 240.244
R14255 GND.n6687 GND.n1067 240.244
R14256 GND.n6691 GND.n1067 240.244
R14257 GND.n6691 GND.n1063 240.244
R14258 GND.n6697 GND.n1063 240.244
R14259 GND.n6697 GND.n1061 240.244
R14260 GND.n6701 GND.n1061 240.244
R14261 GND.n6701 GND.n1057 240.244
R14262 GND.n6707 GND.n1057 240.244
R14263 GND.n6707 GND.n1055 240.244
R14264 GND.n6711 GND.n1055 240.244
R14265 GND.n6711 GND.n1051 240.244
R14266 GND.n6717 GND.n1051 240.244
R14267 GND.n6717 GND.n1049 240.244
R14268 GND.n6721 GND.n1049 240.244
R14269 GND.n6721 GND.n1045 240.244
R14270 GND.n6727 GND.n1045 240.244
R14271 GND.n6727 GND.n1043 240.244
R14272 GND.n6731 GND.n1043 240.244
R14273 GND.n6731 GND.n1039 240.244
R14274 GND.n6737 GND.n1039 240.244
R14275 GND.n6737 GND.n1037 240.244
R14276 GND.n6741 GND.n1037 240.244
R14277 GND.n6741 GND.n1033 240.244
R14278 GND.n6747 GND.n1033 240.244
R14279 GND.n6747 GND.n1031 240.244
R14280 GND.n6751 GND.n1031 240.244
R14281 GND.n6751 GND.n1027 240.244
R14282 GND.n6757 GND.n1027 240.244
R14283 GND.n6757 GND.n1025 240.244
R14284 GND.n6761 GND.n1025 240.244
R14285 GND.n6761 GND.n1021 240.244
R14286 GND.n6767 GND.n1021 240.244
R14287 GND.n6767 GND.n1019 240.244
R14288 GND.n6771 GND.n1019 240.244
R14289 GND.n6771 GND.n1015 240.244
R14290 GND.n6777 GND.n1015 240.244
R14291 GND.n6777 GND.n1013 240.244
R14292 GND.n6781 GND.n1013 240.244
R14293 GND.n6781 GND.n1009 240.244
R14294 GND.n6787 GND.n1009 240.244
R14295 GND.n6787 GND.n1007 240.244
R14296 GND.n6791 GND.n1007 240.244
R14297 GND.n6791 GND.n1003 240.244
R14298 GND.n6797 GND.n1003 240.244
R14299 GND.n6797 GND.n1001 240.244
R14300 GND.n6801 GND.n1001 240.244
R14301 GND.n6801 GND.n997 240.244
R14302 GND.n6807 GND.n997 240.244
R14303 GND.n6807 GND.n995 240.244
R14304 GND.n6811 GND.n995 240.244
R14305 GND.n6811 GND.n991 240.244
R14306 GND.n6817 GND.n991 240.244
R14307 GND.n6817 GND.n989 240.244
R14308 GND.n6821 GND.n989 240.244
R14309 GND.n6821 GND.n985 240.244
R14310 GND.n6827 GND.n985 240.244
R14311 GND.n6827 GND.n983 240.244
R14312 GND.n6831 GND.n983 240.244
R14313 GND.n6831 GND.n979 240.244
R14314 GND.n6837 GND.n979 240.244
R14315 GND.n6837 GND.n977 240.244
R14316 GND.n6841 GND.n977 240.244
R14317 GND.n6841 GND.n973 240.244
R14318 GND.n6847 GND.n973 240.244
R14319 GND.n6847 GND.n971 240.244
R14320 GND.n6851 GND.n971 240.244
R14321 GND.n6851 GND.n967 240.244
R14322 GND.n6857 GND.n967 240.244
R14323 GND.n6857 GND.n965 240.244
R14324 GND.n6861 GND.n965 240.244
R14325 GND.n6861 GND.n961 240.244
R14326 GND.n6867 GND.n961 240.244
R14327 GND.n6867 GND.n959 240.244
R14328 GND.n6871 GND.n959 240.244
R14329 GND.n6871 GND.n955 240.244
R14330 GND.n6877 GND.n955 240.244
R14331 GND.n6877 GND.n953 240.244
R14332 GND.n6881 GND.n953 240.244
R14333 GND.n6881 GND.n949 240.244
R14334 GND.n6887 GND.n949 240.244
R14335 GND.n6887 GND.n947 240.244
R14336 GND.n6891 GND.n947 240.244
R14337 GND.n6891 GND.n943 240.244
R14338 GND.n6897 GND.n943 240.244
R14339 GND.n6897 GND.n941 240.244
R14340 GND.n6901 GND.n941 240.244
R14341 GND.n6901 GND.n937 240.244
R14342 GND.n6907 GND.n937 240.244
R14343 GND.n6907 GND.n935 240.244
R14344 GND.n6911 GND.n935 240.244
R14345 GND.n6911 GND.n931 240.244
R14346 GND.n6917 GND.n931 240.244
R14347 GND.n6917 GND.n929 240.244
R14348 GND.n6921 GND.n929 240.244
R14349 GND.n6921 GND.n925 240.244
R14350 GND.n6927 GND.n925 240.244
R14351 GND.n6927 GND.n923 240.244
R14352 GND.n6931 GND.n923 240.244
R14353 GND.n6931 GND.n919 240.244
R14354 GND.n6937 GND.n919 240.244
R14355 GND.n6937 GND.n917 240.244
R14356 GND.n6941 GND.n917 240.244
R14357 GND.n6941 GND.n913 240.244
R14358 GND.n6947 GND.n913 240.244
R14359 GND.n6947 GND.n911 240.244
R14360 GND.n6951 GND.n911 240.244
R14361 GND.n6951 GND.n907 240.244
R14362 GND.n6957 GND.n907 240.244
R14363 GND.n6957 GND.n905 240.244
R14364 GND.n6961 GND.n905 240.244
R14365 GND.n6961 GND.n901 240.244
R14366 GND.n6967 GND.n901 240.244
R14367 GND.n6967 GND.n899 240.244
R14368 GND.n6971 GND.n899 240.244
R14369 GND.n6971 GND.n895 240.244
R14370 GND.n6977 GND.n895 240.244
R14371 GND.n6977 GND.n893 240.244
R14372 GND.n6981 GND.n893 240.244
R14373 GND.n6981 GND.n889 240.244
R14374 GND.n6987 GND.n889 240.244
R14375 GND.n6987 GND.n887 240.244
R14376 GND.n6991 GND.n887 240.244
R14377 GND.n6991 GND.n883 240.244
R14378 GND.n6997 GND.n883 240.244
R14379 GND.n6997 GND.n881 240.244
R14380 GND.n7001 GND.n881 240.244
R14381 GND.n7001 GND.n877 240.244
R14382 GND.n7007 GND.n877 240.244
R14383 GND.n7007 GND.n875 240.244
R14384 GND.n7011 GND.n875 240.244
R14385 GND.n7011 GND.n871 240.244
R14386 GND.n7017 GND.n871 240.244
R14387 GND.n7017 GND.n869 240.244
R14388 GND.n7021 GND.n869 240.244
R14389 GND.n7021 GND.n865 240.244
R14390 GND.n7027 GND.n865 240.244
R14391 GND.n7027 GND.n863 240.244
R14392 GND.n7031 GND.n863 240.244
R14393 GND.n7031 GND.n859 240.244
R14394 GND.n7037 GND.n859 240.244
R14395 GND.n7037 GND.n857 240.244
R14396 GND.n7041 GND.n857 240.244
R14397 GND.n7041 GND.n853 240.244
R14398 GND.n7047 GND.n853 240.244
R14399 GND.n7047 GND.n851 240.244
R14400 GND.n7051 GND.n851 240.244
R14401 GND.n7051 GND.n847 240.244
R14402 GND.n7057 GND.n847 240.244
R14403 GND.n7057 GND.n845 240.244
R14404 GND.n7061 GND.n845 240.244
R14405 GND.n7061 GND.n841 240.244
R14406 GND.n7067 GND.n841 240.244
R14407 GND.n7067 GND.n839 240.244
R14408 GND.n7071 GND.n839 240.244
R14409 GND.n7071 GND.n835 240.244
R14410 GND.n7077 GND.n835 240.244
R14411 GND.n7077 GND.n833 240.244
R14412 GND.n7081 GND.n833 240.244
R14413 GND.n7081 GND.n829 240.244
R14414 GND.n7087 GND.n829 240.244
R14415 GND.n7087 GND.n827 240.244
R14416 GND.n7091 GND.n827 240.244
R14417 GND.n7091 GND.n823 240.244
R14418 GND.n7097 GND.n823 240.244
R14419 GND.n7097 GND.n821 240.244
R14420 GND.n7101 GND.n821 240.244
R14421 GND.n7101 GND.n817 240.244
R14422 GND.n7107 GND.n817 240.244
R14423 GND.n7107 GND.n815 240.244
R14424 GND.n7111 GND.n815 240.244
R14425 GND.n7111 GND.n811 240.244
R14426 GND.n7117 GND.n811 240.244
R14427 GND.n7117 GND.n809 240.244
R14428 GND.n7121 GND.n809 240.244
R14429 GND.n7121 GND.n805 240.244
R14430 GND.n7127 GND.n805 240.244
R14431 GND.n7127 GND.n803 240.244
R14432 GND.n7131 GND.n803 240.244
R14433 GND.n7131 GND.n799 240.244
R14434 GND.n7137 GND.n799 240.244
R14435 GND.n7137 GND.n797 240.244
R14436 GND.n7141 GND.n797 240.244
R14437 GND.n7141 GND.n793 240.244
R14438 GND.n7147 GND.n793 240.244
R14439 GND.n7147 GND.n791 240.244
R14440 GND.n7151 GND.n791 240.244
R14441 GND.n7151 GND.n787 240.244
R14442 GND.n7157 GND.n787 240.244
R14443 GND.n7157 GND.n785 240.244
R14444 GND.n7161 GND.n785 240.244
R14445 GND.n7161 GND.n781 240.244
R14446 GND.n7167 GND.n781 240.244
R14447 GND.n7167 GND.n779 240.244
R14448 GND.n7171 GND.n779 240.244
R14449 GND.n7171 GND.n775 240.244
R14450 GND.n7177 GND.n775 240.244
R14451 GND.n7177 GND.n773 240.244
R14452 GND.n7181 GND.n773 240.244
R14453 GND.n7181 GND.n769 240.244
R14454 GND.n7187 GND.n769 240.244
R14455 GND.n7187 GND.n767 240.244
R14456 GND.n7191 GND.n767 240.244
R14457 GND.n7191 GND.n763 240.244
R14458 GND.n7197 GND.n763 240.244
R14459 GND.n7197 GND.n761 240.244
R14460 GND.n7201 GND.n761 240.244
R14461 GND.n7201 GND.n757 240.244
R14462 GND.n7207 GND.n757 240.244
R14463 GND.n7207 GND.n755 240.244
R14464 GND.n7211 GND.n755 240.244
R14465 GND.n7211 GND.n751 240.244
R14466 GND.n7217 GND.n751 240.244
R14467 GND.n7217 GND.n749 240.244
R14468 GND.n7221 GND.n749 240.244
R14469 GND.n7221 GND.n745 240.244
R14470 GND.n7227 GND.n745 240.244
R14471 GND.n7227 GND.n743 240.244
R14472 GND.n7231 GND.n743 240.244
R14473 GND.n7231 GND.n739 240.244
R14474 GND.n7237 GND.n739 240.244
R14475 GND.n7237 GND.n737 240.244
R14476 GND.n7241 GND.n737 240.244
R14477 GND.n7241 GND.n733 240.244
R14478 GND.n7247 GND.n733 240.244
R14479 GND.n7247 GND.n731 240.244
R14480 GND.n7251 GND.n731 240.244
R14481 GND.n7251 GND.n727 240.244
R14482 GND.n7257 GND.n727 240.244
R14483 GND.n7257 GND.n725 240.244
R14484 GND.n7261 GND.n725 240.244
R14485 GND.n7261 GND.n721 240.244
R14486 GND.n7267 GND.n721 240.244
R14487 GND.n7267 GND.n719 240.244
R14488 GND.n7271 GND.n719 240.244
R14489 GND.n7271 GND.n715 240.244
R14490 GND.n7277 GND.n715 240.244
R14491 GND.n7277 GND.n713 240.244
R14492 GND.n7281 GND.n713 240.244
R14493 GND.n7281 GND.n709 240.244
R14494 GND.n7287 GND.n709 240.244
R14495 GND.n7287 GND.n707 240.244
R14496 GND.n7291 GND.n707 240.244
R14497 GND.n7291 GND.n703 240.244
R14498 GND.n7297 GND.n703 240.244
R14499 GND.n7297 GND.n701 240.244
R14500 GND.n7301 GND.n701 240.244
R14501 GND.n7301 GND.n697 240.244
R14502 GND.n7307 GND.n697 240.244
R14503 GND.n7307 GND.n695 240.244
R14504 GND.n7311 GND.n695 240.244
R14505 GND.n7311 GND.n691 240.244
R14506 GND.n7317 GND.n691 240.244
R14507 GND.n7317 GND.n689 240.244
R14508 GND.n7321 GND.n689 240.244
R14509 GND.n7321 GND.n685 240.244
R14510 GND.n7328 GND.n685 240.244
R14511 GND.n7328 GND.n683 240.244
R14512 GND.n7332 GND.n683 240.244
R14513 GND.n7332 GND.n680 240.244
R14514 GND.n7338 GND.n678 240.244
R14515 GND.n7342 GND.n678 240.244
R14516 GND.n7342 GND.n674 240.244
R14517 GND.n7348 GND.n674 240.244
R14518 GND.n7348 GND.n672 240.244
R14519 GND.n7352 GND.n672 240.244
R14520 GND.n7352 GND.n668 240.244
R14521 GND.n7358 GND.n668 240.244
R14522 GND.n7358 GND.n666 240.244
R14523 GND.n7362 GND.n666 240.244
R14524 GND.n7362 GND.n662 240.244
R14525 GND.n7368 GND.n662 240.244
R14526 GND.n7368 GND.n660 240.244
R14527 GND.n7372 GND.n660 240.244
R14528 GND.n7372 GND.n656 240.244
R14529 GND.n7378 GND.n656 240.244
R14530 GND.n7378 GND.n654 240.244
R14531 GND.n7382 GND.n654 240.244
R14532 GND.n7382 GND.n650 240.244
R14533 GND.n7388 GND.n650 240.244
R14534 GND.n7388 GND.n648 240.244
R14535 GND.n7392 GND.n648 240.244
R14536 GND.n7392 GND.n644 240.244
R14537 GND.n7398 GND.n644 240.244
R14538 GND.n7398 GND.n642 240.244
R14539 GND.n7402 GND.n642 240.244
R14540 GND.n7402 GND.n638 240.244
R14541 GND.n7408 GND.n638 240.244
R14542 GND.n7408 GND.n636 240.244
R14543 GND.n7412 GND.n636 240.244
R14544 GND.n7412 GND.n632 240.244
R14545 GND.n7418 GND.n632 240.244
R14546 GND.n7418 GND.n630 240.244
R14547 GND.n7422 GND.n630 240.244
R14548 GND.n7422 GND.n626 240.244
R14549 GND.n7428 GND.n626 240.244
R14550 GND.n7428 GND.n624 240.244
R14551 GND.n7432 GND.n624 240.244
R14552 GND.n7432 GND.n620 240.244
R14553 GND.n7438 GND.n620 240.244
R14554 GND.n7438 GND.n618 240.244
R14555 GND.n7442 GND.n618 240.244
R14556 GND.n7442 GND.n614 240.244
R14557 GND.n7448 GND.n614 240.244
R14558 GND.n7448 GND.n612 240.244
R14559 GND.n7452 GND.n612 240.244
R14560 GND.n7452 GND.n608 240.244
R14561 GND.n7458 GND.n608 240.244
R14562 GND.n7458 GND.n606 240.244
R14563 GND.n7462 GND.n606 240.244
R14564 GND.n7462 GND.n602 240.244
R14565 GND.n7468 GND.n602 240.244
R14566 GND.n7468 GND.n600 240.244
R14567 GND.n7472 GND.n600 240.244
R14568 GND.n7472 GND.n596 240.244
R14569 GND.n7478 GND.n596 240.244
R14570 GND.n7478 GND.n594 240.244
R14571 GND.n7482 GND.n594 240.244
R14572 GND.n7482 GND.n590 240.244
R14573 GND.n7488 GND.n590 240.244
R14574 GND.n7488 GND.n588 240.244
R14575 GND.n7492 GND.n588 240.244
R14576 GND.n7492 GND.n584 240.244
R14577 GND.n7498 GND.n584 240.244
R14578 GND.n7498 GND.n582 240.244
R14579 GND.n7502 GND.n582 240.244
R14580 GND.n7502 GND.n578 240.244
R14581 GND.n7508 GND.n578 240.244
R14582 GND.n7508 GND.n576 240.244
R14583 GND.n7512 GND.n576 240.244
R14584 GND.n7512 GND.n572 240.244
R14585 GND.n7518 GND.n572 240.244
R14586 GND.n7518 GND.n570 240.244
R14587 GND.n7522 GND.n570 240.244
R14588 GND.n7522 GND.n566 240.244
R14589 GND.n7528 GND.n566 240.244
R14590 GND.n7528 GND.n564 240.244
R14591 GND.n7532 GND.n564 240.244
R14592 GND.n7532 GND.n560 240.244
R14593 GND.n7538 GND.n560 240.244
R14594 GND.n7538 GND.n558 240.244
R14595 GND.n7542 GND.n558 240.244
R14596 GND.n7542 GND.n554 240.244
R14597 GND.n7548 GND.n554 240.244
R14598 GND.n7548 GND.n552 240.244
R14599 GND.n7552 GND.n552 240.244
R14600 GND.n7552 GND.n548 240.244
R14601 GND.n7560 GND.n548 240.244
R14602 GND.n7560 GND.n546 240.244
R14603 GND.n6171 GND.n1445 240.244
R14604 GND.n6171 GND.n1447 240.244
R14605 GND.n6167 GND.n1447 240.244
R14606 GND.n6167 GND.n1454 240.244
R14607 GND.n6163 GND.n1454 240.244
R14608 GND.n6163 GND.n1456 240.244
R14609 GND.n6159 GND.n1456 240.244
R14610 GND.n6159 GND.n1462 240.244
R14611 GND.n6155 GND.n1462 240.244
R14612 GND.n6155 GND.n1464 240.244
R14613 GND.n6151 GND.n1464 240.244
R14614 GND.n6151 GND.n1470 240.244
R14615 GND.n6147 GND.n1470 240.244
R14616 GND.n6147 GND.n1472 240.244
R14617 GND.n6143 GND.n1472 240.244
R14618 GND.n6143 GND.n1478 240.244
R14619 GND.n6139 GND.n1478 240.244
R14620 GND.n6139 GND.n1480 240.244
R14621 GND.n6135 GND.n1480 240.244
R14622 GND.n6135 GND.n1486 240.244
R14623 GND.n6131 GND.n1486 240.244
R14624 GND.n6131 GND.n1488 240.244
R14625 GND.n6127 GND.n1488 240.244
R14626 GND.n6127 GND.n1494 240.244
R14627 GND.n6123 GND.n1494 240.244
R14628 GND.n6123 GND.n1496 240.244
R14629 GND.n6119 GND.n1496 240.244
R14630 GND.n6119 GND.n1502 240.244
R14631 GND.n6115 GND.n1502 240.244
R14632 GND.n6115 GND.n1504 240.244
R14633 GND.n6111 GND.n1504 240.244
R14634 GND.n6111 GND.n1510 240.244
R14635 GND.n6107 GND.n1510 240.244
R14636 GND.n6107 GND.n1512 240.244
R14637 GND.n6103 GND.n1512 240.244
R14638 GND.n6103 GND.n1518 240.244
R14639 GND.n6099 GND.n1518 240.244
R14640 GND.n6099 GND.n1520 240.244
R14641 GND.n6095 GND.n1520 240.244
R14642 GND.n6095 GND.n1526 240.244
R14643 GND.n6091 GND.n1526 240.244
R14644 GND.n6091 GND.n1528 240.244
R14645 GND.n6087 GND.n1528 240.244
R14646 GND.n6087 GND.n1534 240.244
R14647 GND.n6083 GND.n1534 240.244
R14648 GND.n6083 GND.n1536 240.244
R14649 GND.n6079 GND.n1536 240.244
R14650 GND.n6079 GND.n1542 240.244
R14651 GND.n6075 GND.n1542 240.244
R14652 GND.n6075 GND.n1544 240.244
R14653 GND.n6071 GND.n1544 240.244
R14654 GND.n6071 GND.n1550 240.244
R14655 GND.n6067 GND.n1550 240.244
R14656 GND.n6067 GND.n1552 240.244
R14657 GND.n6063 GND.n1552 240.244
R14658 GND.n6063 GND.n1558 240.244
R14659 GND.n6059 GND.n1558 240.244
R14660 GND.n6059 GND.n1560 240.244
R14661 GND.n6055 GND.n1560 240.244
R14662 GND.n6055 GND.n1566 240.244
R14663 GND.n6051 GND.n1566 240.244
R14664 GND.n6051 GND.n1568 240.244
R14665 GND.n6047 GND.n1568 240.244
R14666 GND.n6047 GND.n1574 240.244
R14667 GND.n6043 GND.n1574 240.244
R14668 GND.n6043 GND.n1576 240.244
R14669 GND.n6039 GND.n1576 240.244
R14670 GND.n6039 GND.n1582 240.244
R14671 GND.n6035 GND.n1582 240.244
R14672 GND.n6035 GND.n1584 240.244
R14673 GND.n6031 GND.n1584 240.244
R14674 GND.n6031 GND.n1590 240.244
R14675 GND.n6027 GND.n1590 240.244
R14676 GND.n6027 GND.n1592 240.244
R14677 GND.n6023 GND.n1592 240.244
R14678 GND.n6023 GND.n1598 240.244
R14679 GND.n6019 GND.n1598 240.244
R14680 GND.n6019 GND.n1600 240.244
R14681 GND.n6015 GND.n1600 240.244
R14682 GND.n6015 GND.n1606 240.244
R14683 GND.n6011 GND.n1606 240.244
R14684 GND.n6011 GND.n1608 240.244
R14685 GND.n6007 GND.n1608 240.244
R14686 GND.n6007 GND.n1614 240.244
R14687 GND.n3484 GND.n1614 240.244
R14688 GND.n3490 GND.n3484 240.244
R14689 GND.n3490 GND.n3474 240.244
R14690 GND.n3681 GND.n3474 240.244
R14691 GND.n3681 GND.n3469 240.244
R14692 GND.n3689 GND.n3469 240.244
R14693 GND.n3689 GND.n3470 240.244
R14694 GND.n3470 GND.n3444 240.244
R14695 GND.n3718 GND.n3444 240.244
R14696 GND.n3718 GND.n3439 240.244
R14697 GND.n3726 GND.n3439 240.244
R14698 GND.n3726 GND.n3440 240.244
R14699 GND.n3440 GND.n3415 240.244
R14700 GND.n3755 GND.n3415 240.244
R14701 GND.n3755 GND.n3410 240.244
R14702 GND.n3763 GND.n3410 240.244
R14703 GND.n3763 GND.n3411 240.244
R14704 GND.n3411 GND.n3386 240.244
R14705 GND.n3792 GND.n3386 240.244
R14706 GND.n3792 GND.n3381 240.244
R14707 GND.n3806 GND.n3381 240.244
R14708 GND.n3806 GND.n3382 240.244
R14709 GND.n3802 GND.n3382 240.244
R14710 GND.n3802 GND.n3801 240.244
R14711 GND.n3801 GND.n3334 240.244
R14712 GND.n3939 GND.n3334 240.244
R14713 GND.n3939 GND.n3335 240.244
R14714 GND.n3870 GND.n3335 240.244
R14715 GND.n3873 GND.n3870 240.244
R14716 GND.n3876 GND.n3873 240.244
R14717 GND.n3876 GND.n3864 240.244
R14718 GND.n3890 GND.n3864 240.244
R14719 GND.n3899 GND.n3890 240.244
R14720 GND.n3899 GND.n3896 240.244
R14721 GND.n3896 GND.n3893 240.244
R14722 GND.n3893 GND.n3892 240.244
R14723 GND.n3892 GND.n3323 240.244
R14724 GND.n3946 GND.n3323 240.244
R14725 GND.n3946 GND.n3300 240.244
R14726 GND.n3975 GND.n3300 240.244
R14727 GND.n3975 GND.n3295 240.244
R14728 GND.n3983 GND.n3295 240.244
R14729 GND.n3983 GND.n3296 240.244
R14730 GND.n3296 GND.n3270 240.244
R14731 GND.n4012 GND.n3270 240.244
R14732 GND.n4012 GND.n3265 240.244
R14733 GND.n4020 GND.n3265 240.244
R14734 GND.n4020 GND.n3266 240.244
R14735 GND.n3266 GND.n3241 240.244
R14736 GND.n4049 GND.n3241 240.244
R14737 GND.n4049 GND.n3236 240.244
R14738 GND.n4057 GND.n3236 240.244
R14739 GND.n4057 GND.n3237 240.244
R14740 GND.n3237 GND.n3212 240.244
R14741 GND.n4086 GND.n3212 240.244
R14742 GND.n4086 GND.n3207 240.244
R14743 GND.n4127 GND.n3207 240.244
R14744 GND.n4127 GND.n3208 240.244
R14745 GND.n4123 GND.n3208 240.244
R14746 GND.n4123 GND.n4122 240.244
R14747 GND.n4122 GND.n4121 240.244
R14748 GND.n4121 GND.n4094 240.244
R14749 GND.n4117 GND.n4094 240.244
R14750 GND.n4117 GND.n4116 240.244
R14751 GND.n4116 GND.n4115 240.244
R14752 GND.n4115 GND.n4100 240.244
R14753 GND.n4109 GND.n4100 240.244
R14754 GND.n4109 GND.n4108 240.244
R14755 GND.n4108 GND.n1886 240.244
R14756 GND.n5802 GND.n1886 240.244
R14757 GND.n5802 GND.n1887 240.244
R14758 GND.n5798 GND.n1887 240.244
R14759 GND.n5798 GND.n1893 240.244
R14760 GND.n1999 GND.n1893 240.244
R14761 GND.n1999 GND.n1996 240.244
R14762 GND.n2005 GND.n1996 240.244
R14763 GND.n2006 GND.n2005 240.244
R14764 GND.n2007 GND.n2006 240.244
R14765 GND.n2007 GND.n1991 240.244
R14766 GND.n5763 GND.n1991 240.244
R14767 GND.n5763 GND.n1992 240.244
R14768 GND.n5759 GND.n1992 240.244
R14769 GND.n5759 GND.n2015 240.244
R14770 GND.n2043 GND.n2015 240.244
R14771 GND.n2043 GND.n2039 240.244
R14772 GND.n5743 GND.n2039 240.244
R14773 GND.n5743 GND.n2040 240.244
R14774 GND.n5739 GND.n2040 240.244
R14775 GND.n5739 GND.n2051 240.244
R14776 GND.n2087 GND.n2051 240.244
R14777 GND.n2087 GND.n2083 240.244
R14778 GND.n5722 GND.n2083 240.244
R14779 GND.n5722 GND.n2084 240.244
R14780 GND.n5718 GND.n2084 240.244
R14781 GND.n5718 GND.n2095 240.244
R14782 GND.n5708 GND.n2095 240.244
R14783 GND.n5708 GND.n2107 240.244
R14784 GND.n5704 GND.n2107 240.244
R14785 GND.n5704 GND.n2113 240.244
R14786 GND.n5694 GND.n2113 240.244
R14787 GND.n5694 GND.n2125 240.244
R14788 GND.n5690 GND.n2125 240.244
R14789 GND.n5690 GND.n2131 240.244
R14790 GND.n5680 GND.n2131 240.244
R14791 GND.n5680 GND.n2142 240.244
R14792 GND.n5676 GND.n2142 240.244
R14793 GND.n5676 GND.n2148 240.244
R14794 GND.n5666 GND.n2148 240.244
R14795 GND.n5666 GND.n2160 240.244
R14796 GND.n5662 GND.n2160 240.244
R14797 GND.n5662 GND.n2166 240.244
R14798 GND.n5652 GND.n2166 240.244
R14799 GND.n5652 GND.n2178 240.244
R14800 GND.n5648 GND.n2178 240.244
R14801 GND.n5648 GND.n2184 240.244
R14802 GND.n2211 GND.n2184 240.244
R14803 GND.n2211 GND.n2207 240.244
R14804 GND.n5631 GND.n2207 240.244
R14805 GND.n5631 GND.n2208 240.244
R14806 GND.n5627 GND.n2208 240.244
R14807 GND.n5627 GND.n2219 240.244
R14808 GND.n2241 GND.n2219 240.244
R14809 GND.n5612 GND.n2241 240.244
R14810 GND.n5612 GND.n2242 240.244
R14811 GND.n5608 GND.n2242 240.244
R14812 GND.n5608 GND.n2250 240.244
R14813 GND.n5598 GND.n2250 240.244
R14814 GND.n5598 GND.n2262 240.244
R14815 GND.n5594 GND.n2262 240.244
R14816 GND.n5594 GND.n2268 240.244
R14817 GND.n2296 GND.n2268 240.244
R14818 GND.n2296 GND.n2292 240.244
R14819 GND.n5577 GND.n2292 240.244
R14820 GND.n5577 GND.n2293 240.244
R14821 GND.n5573 GND.n2293 240.244
R14822 GND.n5573 GND.n2304 240.244
R14823 GND.n4723 GND.n2304 240.244
R14824 GND.n4724 GND.n4723 240.244
R14825 GND.n4725 GND.n4724 240.244
R14826 GND.n4725 GND.n4715 240.244
R14827 GND.n4736 GND.n4715 240.244
R14828 GND.n4736 GND.n4716 240.244
R14829 GND.n4732 GND.n4716 240.244
R14830 GND.n4732 GND.n2940 240.244
R14831 GND.n4770 GND.n2940 240.244
R14832 GND.n4770 GND.n2935 240.244
R14833 GND.n4789 GND.n2935 240.244
R14834 GND.n4789 GND.n2936 240.244
R14835 GND.n4785 GND.n2936 240.244
R14836 GND.n4785 GND.n4783 240.244
R14837 GND.n4783 GND.n4782 240.244
R14838 GND.n4782 GND.n2435 240.244
R14839 GND.n5456 GND.n2435 240.244
R14840 GND.n5456 GND.n2436 240.244
R14841 GND.n5452 GND.n2436 240.244
R14842 GND.n5452 GND.n2442 240.244
R14843 GND.n4810 GND.n2442 240.244
R14844 GND.n4814 GND.n4810 240.244
R14845 GND.n4815 GND.n4814 240.244
R14846 GND.n4815 GND.n4802 240.244
R14847 GND.n4824 GND.n4802 240.244
R14848 GND.n4824 GND.n4803 240.244
R14849 GND.n4803 GND.n2609 240.244
R14850 GND.n5323 GND.n2609 240.244
R14851 GND.n5323 GND.n2610 240.244
R14852 GND.n5319 GND.n2610 240.244
R14853 GND.n5319 GND.n2616 240.244
R14854 GND.n2832 GND.n2616 240.244
R14855 GND.n2890 GND.n2832 240.244
R14856 GND.n2890 GND.n2833 240.244
R14857 GND.n2886 GND.n2833 240.244
R14858 GND.n2886 GND.n2885 240.244
R14859 GND.n2885 GND.n2884 240.244
R14860 GND.n2884 GND.n2841 240.244
R14861 GND.n2880 GND.n2841 240.244
R14862 GND.n2880 GND.n2879 240.244
R14863 GND.n2879 GND.n2878 240.244
R14864 GND.n2878 GND.n2847 240.244
R14865 GND.n2874 GND.n2847 240.244
R14866 GND.n2874 GND.n2873 240.244
R14867 GND.n2873 GND.n2872 240.244
R14868 GND.n2872 GND.n2853 240.244
R14869 GND.n2868 GND.n2853 240.244
R14870 GND.n2868 GND.n2867 240.244
R14871 GND.n2867 GND.n2866 240.244
R14872 GND.n2866 GND.n2859 240.244
R14873 GND.n2859 GND.n2739 240.244
R14874 GND.n5251 GND.n2739 240.244
R14875 GND.n5251 GND.n2740 240.244
R14876 GND.n5246 GND.n2740 240.244
R14877 GND.n5246 GND.n2743 240.244
R14878 GND.n2760 GND.n2743 240.244
R14879 GND.n5236 GND.n2760 240.244
R14880 GND.n5236 GND.n2761 240.244
R14881 GND.n5231 GND.n2761 240.244
R14882 GND.n5231 GND.n5230 240.244
R14883 GND.n5230 GND.n2765 240.244
R14884 GND.n5226 GND.n2765 240.244
R14885 GND.n5226 GND.n5225 240.244
R14886 GND.n5225 GND.n5224 240.244
R14887 GND.n5224 GND.n2769 240.244
R14888 GND.n5220 GND.n2769 240.244
R14889 GND.n5220 GND.n5219 240.244
R14890 GND.n5219 GND.n5218 240.244
R14891 GND.n5218 GND.n2775 240.244
R14892 GND.n5214 GND.n2775 240.244
R14893 GND.n5214 GND.n5213 240.244
R14894 GND.n5213 GND.n5212 240.244
R14895 GND.n5212 GND.n2781 240.244
R14896 GND.n5208 GND.n2781 240.244
R14897 GND.n5208 GND.n5207 240.244
R14898 GND.n5207 GND.n5206 240.244
R14899 GND.n5206 GND.n5181 240.244
R14900 GND.n5202 GND.n5181 240.244
R14901 GND.n5202 GND.n5201 240.244
R14902 GND.n5201 GND.n5200 240.244
R14903 GND.n5200 GND.n5187 240.244
R14904 GND.n5196 GND.n5187 240.244
R14905 GND.n5196 GND.n5195 240.244
R14906 GND.n5195 GND.n183 240.244
R14907 GND.n7736 GND.n183 240.244
R14908 GND.n7736 GND.n184 240.244
R14909 GND.n7732 GND.n184 240.244
R14910 GND.n7732 GND.n190 240.244
R14911 GND.n7728 GND.n190 240.244
R14912 GND.n7728 GND.n381 240.244
R14913 GND.n7724 GND.n381 240.244
R14914 GND.n7724 GND.n387 240.244
R14915 GND.n7720 GND.n387 240.244
R14916 GND.n7720 GND.n389 240.244
R14917 GND.n7716 GND.n389 240.244
R14918 GND.n7716 GND.n395 240.244
R14919 GND.n7712 GND.n395 240.244
R14920 GND.n7712 GND.n397 240.244
R14921 GND.n7708 GND.n397 240.244
R14922 GND.n7708 GND.n403 240.244
R14923 GND.n7704 GND.n403 240.244
R14924 GND.n7704 GND.n405 240.244
R14925 GND.n7700 GND.n405 240.244
R14926 GND.n7700 GND.n411 240.244
R14927 GND.n7696 GND.n411 240.244
R14928 GND.n7696 GND.n413 240.244
R14929 GND.n7692 GND.n413 240.244
R14930 GND.n7692 GND.n419 240.244
R14931 GND.n7688 GND.n419 240.244
R14932 GND.n7688 GND.n421 240.244
R14933 GND.n7684 GND.n421 240.244
R14934 GND.n7684 GND.n427 240.244
R14935 GND.n7680 GND.n427 240.244
R14936 GND.n7680 GND.n429 240.244
R14937 GND.n7676 GND.n429 240.244
R14938 GND.n7676 GND.n435 240.244
R14939 GND.n7672 GND.n435 240.244
R14940 GND.n7672 GND.n437 240.244
R14941 GND.n7668 GND.n437 240.244
R14942 GND.n7668 GND.n443 240.244
R14943 GND.n7664 GND.n443 240.244
R14944 GND.n7664 GND.n445 240.244
R14945 GND.n7660 GND.n445 240.244
R14946 GND.n7660 GND.n451 240.244
R14947 GND.n7656 GND.n451 240.244
R14948 GND.n7656 GND.n453 240.244
R14949 GND.n7652 GND.n453 240.244
R14950 GND.n7652 GND.n459 240.244
R14951 GND.n7648 GND.n459 240.244
R14952 GND.n7648 GND.n461 240.244
R14953 GND.n7644 GND.n461 240.244
R14954 GND.n7644 GND.n467 240.244
R14955 GND.n7640 GND.n467 240.244
R14956 GND.n7640 GND.n469 240.244
R14957 GND.n7636 GND.n469 240.244
R14958 GND.n7636 GND.n475 240.244
R14959 GND.n7632 GND.n475 240.244
R14960 GND.n7632 GND.n477 240.244
R14961 GND.n7628 GND.n477 240.244
R14962 GND.n7628 GND.n483 240.244
R14963 GND.n7624 GND.n483 240.244
R14964 GND.n7624 GND.n485 240.244
R14965 GND.n7620 GND.n485 240.244
R14966 GND.n7620 GND.n491 240.244
R14967 GND.n7616 GND.n491 240.244
R14968 GND.n7616 GND.n493 240.244
R14969 GND.n7612 GND.n493 240.244
R14970 GND.n7612 GND.n499 240.244
R14971 GND.n7608 GND.n499 240.244
R14972 GND.n7608 GND.n501 240.244
R14973 GND.n7604 GND.n501 240.244
R14974 GND.n7604 GND.n507 240.244
R14975 GND.n7600 GND.n507 240.244
R14976 GND.n7600 GND.n509 240.244
R14977 GND.n7596 GND.n509 240.244
R14978 GND.n7596 GND.n515 240.244
R14979 GND.n7592 GND.n515 240.244
R14980 GND.n7592 GND.n517 240.244
R14981 GND.n7588 GND.n517 240.244
R14982 GND.n7588 GND.n523 240.244
R14983 GND.n7584 GND.n523 240.244
R14984 GND.n7584 GND.n525 240.244
R14985 GND.n7580 GND.n525 240.244
R14986 GND.n7580 GND.n531 240.244
R14987 GND.n7576 GND.n531 240.244
R14988 GND.n7576 GND.n533 240.244
R14989 GND.n7572 GND.n533 240.244
R14990 GND.n7572 GND.n539 240.244
R14991 GND.n7568 GND.n539 240.244
R14992 GND.n7568 GND.n541 240.244
R14993 GND.n7564 GND.n541 240.244
R14994 GND.n6351 GND.n1267 240.244
R14995 GND.n6351 GND.n1270 240.244
R14996 GND.n6347 GND.n1270 240.244
R14997 GND.n6347 GND.n1272 240.244
R14998 GND.n6343 GND.n1272 240.244
R14999 GND.n6343 GND.n1278 240.244
R15000 GND.n6339 GND.n1278 240.244
R15001 GND.n6339 GND.n1280 240.244
R15002 GND.n6335 GND.n1280 240.244
R15003 GND.n6335 GND.n1286 240.244
R15004 GND.n6331 GND.n1286 240.244
R15005 GND.n6331 GND.n1288 240.244
R15006 GND.n6327 GND.n1288 240.244
R15007 GND.n6327 GND.n1294 240.244
R15008 GND.n6323 GND.n1294 240.244
R15009 GND.n6323 GND.n1296 240.244
R15010 GND.n6319 GND.n1296 240.244
R15011 GND.n6319 GND.n1302 240.244
R15012 GND.n6315 GND.n1302 240.244
R15013 GND.n6315 GND.n1304 240.244
R15014 GND.n6311 GND.n1304 240.244
R15015 GND.n6311 GND.n1310 240.244
R15016 GND.n6307 GND.n1310 240.244
R15017 GND.n6307 GND.n1312 240.244
R15018 GND.n6303 GND.n1312 240.244
R15019 GND.n6303 GND.n1318 240.244
R15020 GND.n6299 GND.n1318 240.244
R15021 GND.n6299 GND.n1320 240.244
R15022 GND.n6295 GND.n1320 240.244
R15023 GND.n6295 GND.n1326 240.244
R15024 GND.n6291 GND.n1326 240.244
R15025 GND.n6291 GND.n1328 240.244
R15026 GND.n6287 GND.n1328 240.244
R15027 GND.n6287 GND.n1334 240.244
R15028 GND.n6283 GND.n1334 240.244
R15029 GND.n6283 GND.n1336 240.244
R15030 GND.n6279 GND.n1336 240.244
R15031 GND.n6279 GND.n1342 240.244
R15032 GND.n6275 GND.n1342 240.244
R15033 GND.n6275 GND.n1344 240.244
R15034 GND.n6271 GND.n1344 240.244
R15035 GND.n6271 GND.n1350 240.244
R15036 GND.n6267 GND.n1350 240.244
R15037 GND.n6267 GND.n1352 240.244
R15038 GND.n6263 GND.n1352 240.244
R15039 GND.n6263 GND.n1358 240.244
R15040 GND.n6259 GND.n1358 240.244
R15041 GND.n6259 GND.n1360 240.244
R15042 GND.n6255 GND.n1360 240.244
R15043 GND.n6255 GND.n1366 240.244
R15044 GND.n6251 GND.n1366 240.244
R15045 GND.n6251 GND.n1368 240.244
R15046 GND.n6247 GND.n1368 240.244
R15047 GND.n6247 GND.n1374 240.244
R15048 GND.n6243 GND.n1374 240.244
R15049 GND.n6243 GND.n1376 240.244
R15050 GND.n6239 GND.n1376 240.244
R15051 GND.n6239 GND.n1382 240.244
R15052 GND.n6235 GND.n1382 240.244
R15053 GND.n6235 GND.n1384 240.244
R15054 GND.n6231 GND.n1384 240.244
R15055 GND.n6231 GND.n1390 240.244
R15056 GND.n6227 GND.n1390 240.244
R15057 GND.n6227 GND.n1392 240.244
R15058 GND.n6223 GND.n1392 240.244
R15059 GND.n6223 GND.n1398 240.244
R15060 GND.n6219 GND.n1398 240.244
R15061 GND.n6219 GND.n1400 240.244
R15062 GND.n6215 GND.n1400 240.244
R15063 GND.n6215 GND.n1406 240.244
R15064 GND.n6211 GND.n1406 240.244
R15065 GND.n6211 GND.n1408 240.244
R15066 GND.n6207 GND.n1408 240.244
R15067 GND.n6207 GND.n1414 240.244
R15068 GND.n6203 GND.n1414 240.244
R15069 GND.n6203 GND.n1416 240.244
R15070 GND.n6199 GND.n1416 240.244
R15071 GND.n6199 GND.n1422 240.244
R15072 GND.n6195 GND.n1422 240.244
R15073 GND.n6195 GND.n1424 240.244
R15074 GND.n6191 GND.n1424 240.244
R15075 GND.n6191 GND.n1430 240.244
R15076 GND.n6187 GND.n1430 240.244
R15077 GND.n6187 GND.n1432 240.244
R15078 GND.n6183 GND.n1432 240.244
R15079 GND.n6183 GND.n1438 240.244
R15080 GND.n6179 GND.n1438 240.244
R15081 GND.n6179 GND.n1440 240.244
R15082 GND.n6175 GND.n1440 240.244
R15083 GND.n6003 GND.n1649 240.244
R15084 GND.n1654 GND.n1653 240.244
R15085 GND.n1656 GND.n1655 240.244
R15086 GND.n1660 GND.n1659 240.244
R15087 GND.n1662 GND.n1661 240.244
R15088 GND.n1663 GND.n1646 240.244
R15089 GND.n3656 GND.n1648 240.244
R15090 GND.n3656 GND.n3478 240.244
R15091 GND.n3659 GND.n3478 240.244
R15092 GND.n3659 GND.n3459 240.244
R15093 GND.n3705 GND.n3459 240.244
R15094 GND.n3705 GND.n3460 240.244
R15095 GND.n3460 GND.n3449 240.244
R15096 GND.n3696 GND.n3449 240.244
R15097 GND.n3696 GND.n3430 240.244
R15098 GND.n3742 GND.n3430 240.244
R15099 GND.n3742 GND.n3431 240.244
R15100 GND.n3431 GND.n3420 240.244
R15101 GND.n3733 GND.n3420 240.244
R15102 GND.n3733 GND.n3401 240.244
R15103 GND.n3779 GND.n3401 240.244
R15104 GND.n3779 GND.n3402 240.244
R15105 GND.n3402 GND.n3390 240.244
R15106 GND.n3770 GND.n3390 240.244
R15107 GND.n3770 GND.n3370 240.244
R15108 GND.n3816 GND.n3370 240.244
R15109 GND.n3816 GND.n3372 240.244
R15110 GND.n3372 GND.n3357 240.244
R15111 GND.n3831 GND.n3357 240.244
R15112 GND.n3831 GND.n3338 240.244
R15113 GND.n3348 GND.n3338 240.244
R15114 GND.n3929 GND.n3348 240.244
R15115 GND.n3929 GND.n3349 240.244
R15116 GND.n3878 GND.n3349 240.244
R15117 GND.n3878 GND.n3867 240.244
R15118 GND.n3867 GND.n3861 240.244
R15119 GND.n3903 GND.n3861 240.244
R15120 GND.n3904 GND.n3903 240.244
R15121 GND.n3904 GND.n3852 240.244
R15122 GND.n3913 GND.n3852 240.244
R15123 GND.n3913 GND.n3313 240.244
R15124 GND.n3962 GND.n3313 240.244
R15125 GND.n3962 GND.n3314 240.244
R15126 GND.n3314 GND.n3304 240.244
R15127 GND.n3953 GND.n3304 240.244
R15128 GND.n3953 GND.n3285 240.244
R15129 GND.n3999 GND.n3285 240.244
R15130 GND.n3999 GND.n3286 240.244
R15131 GND.n3286 GND.n3275 240.244
R15132 GND.n3990 GND.n3275 240.244
R15133 GND.n3990 GND.n3256 240.244
R15134 GND.n4036 GND.n3256 240.244
R15135 GND.n4036 GND.n3257 240.244
R15136 GND.n3257 GND.n3246 240.244
R15137 GND.n4027 GND.n3246 240.244
R15138 GND.n4027 GND.n3227 240.244
R15139 GND.n4073 GND.n3227 240.244
R15140 GND.n4073 GND.n3228 240.244
R15141 GND.n3228 GND.n3216 240.244
R15142 GND.n4064 GND.n3216 240.244
R15143 GND.n4064 GND.n3199 240.244
R15144 GND.n4139 GND.n3199 240.244
R15145 GND.n4139 GND.n3188 240.244
R15146 GND.n4150 GND.n3188 240.244
R15147 GND.n4222 GND.n4150 240.244
R15148 GND.n4159 GND.n4158 240.244
R15149 GND.n4161 GND.n4160 240.244
R15150 GND.n4172 GND.n4171 240.244
R15151 GND.n4182 GND.n4181 240.244
R15152 GND.n4183 GND.n1749 240.244
R15153 GND.n1669 GND.n1668 240.244
R15154 GND.n1670 GND.n1669 240.244
R15155 GND.n3467 GND.n1670 240.244
R15156 GND.n3467 GND.n1673 240.244
R15157 GND.n1674 GND.n1673 240.244
R15158 GND.n1675 GND.n1674 240.244
R15159 GND.n3447 GND.n1675 240.244
R15160 GND.n3447 GND.n1678 240.244
R15161 GND.n1679 GND.n1678 240.244
R15162 GND.n1680 GND.n1679 240.244
R15163 GND.n3416 GND.n1680 240.244
R15164 GND.n3416 GND.n1683 240.244
R15165 GND.n1684 GND.n1683 240.244
R15166 GND.n1685 GND.n1684 240.244
R15167 GND.n3399 GND.n1685 240.244
R15168 GND.n3399 GND.n1688 240.244
R15169 GND.n1689 GND.n1688 240.244
R15170 GND.n1690 GND.n1689 240.244
R15171 GND.n3808 GND.n1690 240.244
R15172 GND.n3808 GND.n1693 240.244
R15173 GND.n1694 GND.n1693 240.244
R15174 GND.n1695 GND.n1694 240.244
R15175 GND.n3829 GND.n1695 240.244
R15176 GND.n3829 GND.n1698 240.244
R15177 GND.n1699 GND.n1698 240.244
R15178 GND.n1700 GND.n1699 240.244
R15179 GND.n3868 GND.n1700 240.244
R15180 GND.n3868 GND.n1703 240.244
R15181 GND.n1704 GND.n1703 240.244
R15182 GND.n1705 GND.n1704 240.244
R15183 GND.n3901 GND.n1705 240.244
R15184 GND.n3901 GND.n1709 240.244
R15185 GND.n1710 GND.n1709 240.244
R15186 GND.n1711 GND.n1710 240.244
R15187 GND.n3322 GND.n1711 240.244
R15188 GND.n3322 GND.n1714 240.244
R15189 GND.n1715 GND.n1714 240.244
R15190 GND.n1716 GND.n1715 240.244
R15191 GND.n3293 GND.n1716 240.244
R15192 GND.n3293 GND.n1719 240.244
R15193 GND.n1720 GND.n1719 240.244
R15194 GND.n1721 GND.n1720 240.244
R15195 GND.n3273 GND.n1721 240.244
R15196 GND.n3273 GND.n1724 240.244
R15197 GND.n1725 GND.n1724 240.244
R15198 GND.n1726 GND.n1725 240.244
R15199 GND.n3242 GND.n1726 240.244
R15200 GND.n3242 GND.n1729 240.244
R15201 GND.n1730 GND.n1729 240.244
R15202 GND.n1731 GND.n1730 240.244
R15203 GND.n3225 GND.n1731 240.244
R15204 GND.n3225 GND.n1734 240.244
R15205 GND.n1735 GND.n1734 240.244
R15206 GND.n1736 GND.n1735 240.244
R15207 GND.n4129 GND.n1736 240.244
R15208 GND.n4129 GND.n1739 240.244
R15209 GND.n1740 GND.n1739 240.244
R15210 GND.n1741 GND.n1740 240.244
R15211 GND.n1748 GND.n1741 240.244
R15212 GND.n1861 GND.n1860 240.132
R15213 GND.n1859 GND.n1858 240.132
R15214 GND.n2488 GND.n2487 240.132
R15215 GND.n2486 GND.n2485 240.132
R15216 GND.n1745 GND.t128 210.554
R15217 GND.n1800 GND.t81 210.554
R15218 GND.n3116 GND.t55 210.554
R15219 GND.n3105 GND.t155 210.554
R15220 GND.n1820 GND.t158 210.554
R15221 GND.n5348 GND.t48 210.554
R15222 GND.n2552 GND.t140 210.554
R15223 GND.n4868 GND.t37 210.554
R15224 GND.n4826 GND.t119 210.554
R15225 GND.n271 GND.t69 210.554
R15226 GND.n256 GND.t72 210.554
R15227 GND.n327 GND.t45 210.554
R15228 GND.n227 GND.t90 210.554
R15229 GND.n5112 GND.t33 210.554
R15230 GND.n2899 GND.t104 210.554
R15231 GND.n3519 GND.t113 210.554
R15232 GND.n3509 GND.t51 210.554
R15233 GND.n3615 GND.t93 210.554
R15234 GND.n3649 GND.t149 210.554
R15235 GND.n1664 GND.t122 210.554
R15236 GND.n5809 GND.t41 210.429
R15237 GND.n1908 GND.t146 210.429
R15238 GND.n2500 GND.t100 210.429
R15239 GND.n2498 GND.t137 210.429
R15240 GND.n2407 GND.t96 209.957
R15241 GND.n4198 GND.t62 209.957
R15242 GND.n2567 GND.n2550 199.319
R15243 GND.n5405 GND.n2550 199.319
R15244 GND.n1822 GND.n1771 199.319
R15245 GND.n1822 GND.n1770 199.319
R15246 GND.n4868 GND.t40 189.087
R15247 GND.n271 GND.t70 189.087
R15248 GND.n1862 GND.n1857 186.49
R15249 GND.n2489 GND.n2484 186.49
R15250 GND.n1908 GND.t148 181.083
R15251 GND.n2500 GND.t102 181.083
R15252 GND.n5809 GND.t44 181.083
R15253 GND.n2498 GND.t138 181.083
R15254 GND.n1745 GND.t129 179.487
R15255 GND.n1800 GND.t82 179.487
R15256 GND.n3116 GND.t57 179.487
R15257 GND.n3105 GND.t156 179.487
R15258 GND.n1820 GND.t159 179.487
R15259 GND.n5348 GND.t50 179.487
R15260 GND.n2552 GND.t142 179.487
R15261 GND.n4826 GND.t121 179.487
R15262 GND.n256 GND.t73 179.487
R15263 GND.n327 GND.t46 179.487
R15264 GND.n227 GND.t91 179.487
R15265 GND.n5112 GND.t35 179.487
R15266 GND.n2899 GND.t106 179.487
R15267 GND.n3519 GND.t115 179.487
R15268 GND.n3509 GND.t54 179.487
R15269 GND.n3615 GND.t95 179.487
R15270 GND.n3649 GND.t151 179.487
R15271 GND.n1664 GND.t124 179.487
R15272 GND.n10 GND.t162 165.251
R15273 GND.n10 GND.t26 164.044
R15274 GND.n5449 GND.n2466 163.367
R15275 GND.n5445 GND.n5444 163.367
R15276 GND.n5441 GND.n5440 163.367
R15277 GND.n5437 GND.n5436 163.367
R15278 GND.n5433 GND.n5432 163.367
R15279 GND.n5429 GND.n5428 163.367
R15280 GND.n5425 GND.n5424 163.367
R15281 GND.n5421 GND.n5420 163.367
R15282 GND.n5416 GND.n5415 163.367
R15283 GND.n5412 GND.n5411 163.367
R15284 GND.n2546 GND.n2444 163.367
R15285 GND.n2544 GND.n2543 163.367
R15286 GND.n2540 GND.n2539 163.367
R15287 GND.n2536 GND.n2535 163.367
R15288 GND.n2532 GND.n2531 163.367
R15289 GND.n2528 GND.n2527 163.367
R15290 GND.n2524 GND.n2523 163.367
R15291 GND.n2520 GND.n2519 163.367
R15292 GND.n2516 GND.n2515 163.367
R15293 GND.n2512 GND.n2511 163.367
R15294 GND.n1949 GND.n1884 163.367
R15295 GND.n1953 GND.n1884 163.367
R15296 GND.n1958 GND.n1953 163.367
R15297 GND.n1959 GND.n1958 163.367
R15298 GND.n1959 GND.n1895 163.367
R15299 GND.n1905 GND.n1895 163.367
R15300 GND.n5790 GND.n1905 163.367
R15301 GND.n5790 GND.n1906 163.367
R15302 GND.n5786 GND.n1906 163.367
R15303 GND.n5786 GND.n1964 163.367
R15304 GND.n1970 GND.n1964 163.367
R15305 GND.n3075 GND.n1970 163.367
R15306 GND.n4274 GND.n3075 163.367
R15307 GND.n4274 GND.n1983 163.367
R15308 GND.n4279 GND.n1983 163.367
R15309 GND.n4279 GND.n1990 163.367
R15310 GND.n3071 GND.n1990 163.367
R15311 GND.n4287 GND.n3071 163.367
R15312 GND.n4287 GND.n3072 163.367
R15313 GND.n4283 GND.n3072 163.367
R15314 GND.n4283 GND.n3056 163.367
R15315 GND.n4322 GND.n3056 163.367
R15316 GND.n4322 GND.n2029 163.367
R15317 GND.n4326 GND.n2029 163.367
R15318 GND.n4326 GND.n2038 163.367
R15319 GND.n4330 GND.n2038 163.367
R15320 GND.n4334 GND.n4330 163.367
R15321 GND.n4334 GND.n2053 163.367
R15322 GND.n4338 GND.n2053 163.367
R15323 GND.n4338 GND.n2061 163.367
R15324 GND.n4341 GND.n2061 163.367
R15325 GND.n4341 GND.n3049 163.367
R15326 GND.n4345 GND.n3049 163.367
R15327 GND.n4346 GND.n4345 163.367
R15328 GND.n4346 GND.n3054 163.367
R15329 GND.n4406 GND.n3054 163.367
R15330 GND.n4406 GND.n2097 163.367
R15331 GND.n4402 GND.n2097 163.367
R15332 GND.n4402 GND.n2105 163.367
R15333 GND.n4397 GND.n2105 163.367
R15334 GND.n4397 GND.n4396 163.367
R15335 GND.n4396 GND.n4391 163.367
R15336 GND.n4391 GND.n2115 163.367
R15337 GND.n4387 GND.n2115 163.367
R15338 GND.n4387 GND.n2123 163.367
R15339 GND.n4382 GND.n2123 163.367
R15340 GND.n4382 GND.n4381 163.367
R15341 GND.n4381 GND.n4376 163.367
R15342 GND.n4376 GND.n2133 163.367
R15343 GND.n4372 GND.n2133 163.367
R15344 GND.n4372 GND.n2141 163.367
R15345 GND.n4368 GND.n2141 163.367
R15346 GND.n4368 GND.n4361 163.367
R15347 GND.n4361 GND.n4360 163.367
R15348 GND.n4360 GND.n2150 163.367
R15349 GND.n4356 GND.n2150 163.367
R15350 GND.n4356 GND.n2158 163.367
R15351 GND.n3000 GND.n2158 163.367
R15352 GND.n4510 GND.n3000 163.367
R15353 GND.n4511 GND.n4510 163.367
R15354 GND.n4511 GND.n2168 163.367
R15355 GND.n4516 GND.n2168 163.367
R15356 GND.n4516 GND.n2176 163.367
R15357 GND.n2997 GND.n2176 163.367
R15358 GND.n4524 GND.n2997 163.367
R15359 GND.n4524 GND.n2998 163.367
R15360 GND.n4520 GND.n2998 163.367
R15361 GND.n4520 GND.n2988 163.367
R15362 GND.n4546 GND.n2988 163.367
R15363 GND.n4546 GND.n2198 163.367
R15364 GND.n4559 GND.n2198 163.367
R15365 GND.n4559 GND.n2205 163.367
R15366 GND.n4555 GND.n2205 163.367
R15367 GND.n4555 GND.n2223 163.367
R15368 GND.n5625 GND.n2223 163.367
R15369 GND.n5625 GND.n2224 163.367
R15370 GND.n5621 GND.n2224 163.367
R15371 GND.n5621 GND.n2227 163.367
R15372 GND.n2237 GND.n2227 163.367
R15373 GND.n4577 GND.n2237 163.367
R15374 GND.n4590 GND.n4577 163.367
R15375 GND.n4590 GND.n4578 163.367
R15376 GND.n4578 GND.n2252 163.367
R15377 GND.n4585 GND.n2252 163.367
R15378 GND.n4585 GND.n2260 163.367
R15379 GND.n2972 GND.n2260 163.367
R15380 GND.n4650 GND.n2972 163.367
R15381 GND.n4651 GND.n4650 163.367
R15382 GND.n4652 GND.n4651 163.367
R15383 GND.n4652 GND.n2970 163.367
R15384 GND.n4672 GND.n2970 163.367
R15385 GND.n4672 GND.n2282 163.367
R15386 GND.n4668 GND.n2282 163.367
R15387 GND.n4668 GND.n2290 163.367
R15388 GND.n4664 GND.n2290 163.367
R15389 GND.n4664 GND.n2962 163.367
R15390 GND.n4660 GND.n2962 163.367
R15391 GND.n4660 GND.n4659 163.367
R15392 GND.n4659 GND.n2958 163.367
R15393 GND.n4655 GND.n2958 163.367
R15394 GND.n4655 GND.n2323 163.367
R15395 GND.n4704 GND.n2323 163.367
R15396 GND.n4704 GND.n2331 163.367
R15397 GND.n2951 GND.n2331 163.367
R15398 GND.n4710 GND.n2951 163.367
R15399 GND.n4710 GND.n2952 163.367
R15400 GND.n2952 GND.n2343 163.367
R15401 GND.n4754 GND.n2343 163.367
R15402 GND.n4754 GND.n2351 163.367
R15403 GND.n4757 GND.n2351 163.367
R15404 GND.n4757 GND.n2946 163.367
R15405 GND.n4767 GND.n2946 163.367
R15406 GND.n4767 GND.n2362 163.367
R15407 GND.n2934 GND.n2362 163.367
R15408 GND.n2934 GND.n2369 163.367
R15409 GND.n4761 GND.n2369 163.367
R15410 GND.n4761 GND.n2416 163.367
R15411 GND.n2421 GND.n2416 163.367
R15412 GND.n5469 GND.n2421 163.367
R15413 GND.n5469 GND.n2422 163.367
R15414 GND.n5465 GND.n2422 163.367
R15415 GND.n5465 GND.n2425 163.367
R15416 GND.n2432 GND.n2425 163.367
R15417 GND.n2506 GND.n2432 163.367
R15418 GND.n2507 GND.n2506 163.367
R15419 GND.n1849 GND.n1848 163.367
R15420 GND.n5840 GND.n1848 163.367
R15421 GND.n5838 GND.n5837 163.367
R15422 GND.n5834 GND.n5833 163.367
R15423 GND.n5830 GND.n5829 163.367
R15424 GND.n5826 GND.n5825 163.367
R15425 GND.n5822 GND.n5821 163.367
R15426 GND.n5818 GND.n5817 163.367
R15427 GND.n5813 GND.n5812 163.367
R15428 GND.n5849 GND.n1826 163.367
R15429 GND.n1911 GND.n1910 163.367
R15430 GND.n1915 GND.n1914 163.367
R15431 GND.n1920 GND.n1919 163.367
R15432 GND.n1924 GND.n1923 163.367
R15433 GND.n1928 GND.n1927 163.367
R15434 GND.n1932 GND.n1931 163.367
R15435 GND.n1936 GND.n1935 163.367
R15436 GND.n1940 GND.n1939 163.367
R15437 GND.n1944 GND.n1943 163.367
R15438 GND.n1946 GND.n1846 163.367
R15439 GND.n5805 GND.n1850 163.367
R15440 GND.n5805 GND.n1882 163.367
R15441 GND.n1956 GND.n1882 163.367
R15442 GND.n1956 GND.n1897 163.367
R15443 GND.n5795 GND.n1897 163.367
R15444 GND.n5795 GND.n1898 163.367
R15445 GND.n5791 GND.n1898 163.367
R15446 GND.n5791 GND.n1901 163.367
R15447 GND.n5784 GND.n1901 163.367
R15448 GND.n5784 GND.n1966 163.367
R15449 GND.n5780 GND.n1966 163.367
R15450 GND.n5780 GND.n1968 163.367
R15451 GND.n1984 GND.n1968 163.367
R15452 GND.n5770 GND.n1984 163.367
R15453 GND.n5770 GND.n1985 163.367
R15454 GND.n5766 GND.n1985 163.367
R15455 GND.n5766 GND.n1988 163.367
R15456 GND.n4295 GND.n1988 163.367
R15457 GND.n4295 GND.n4288 163.367
R15458 GND.n4291 GND.n4288 163.367
R15459 GND.n4291 GND.n4290 163.367
R15460 GND.n4290 GND.n2031 163.367
R15461 GND.n5749 GND.n2031 163.367
R15462 GND.n5749 GND.n2032 163.367
R15463 GND.n5745 GND.n2032 163.367
R15464 GND.n5745 GND.n2035 163.367
R15465 GND.n2055 GND.n2035 163.367
R15466 GND.n5736 GND.n2055 163.367
R15467 GND.n5736 GND.n2056 163.367
R15468 GND.n5732 GND.n2056 163.367
R15469 GND.n5732 GND.n2059 163.367
R15470 GND.n4415 GND.n2059 163.367
R15471 GND.n4415 GND.n3051 163.367
R15472 GND.n4411 GND.n3051 163.367
R15473 GND.n4411 GND.n4410 163.367
R15474 GND.n4410 GND.n2099 163.367
R15475 GND.n5715 GND.n2099 163.367
R15476 GND.n5715 GND.n2100 163.367
R15477 GND.n5711 GND.n2100 163.367
R15478 GND.n5711 GND.n2103 163.367
R15479 GND.n4394 GND.n2103 163.367
R15480 GND.n4394 GND.n2117 163.367
R15481 GND.n5701 GND.n2117 163.367
R15482 GND.n5701 GND.n2118 163.367
R15483 GND.n5697 GND.n2118 163.367
R15484 GND.n5697 GND.n2121 163.367
R15485 GND.n4379 GND.n2121 163.367
R15486 GND.n4379 GND.n2135 163.367
R15487 GND.n5687 GND.n2135 163.367
R15488 GND.n5687 GND.n2136 163.367
R15489 GND.n5683 GND.n2136 163.367
R15490 GND.n5683 GND.n2139 163.367
R15491 GND.n4363 GND.n2139 163.367
R15492 GND.n4363 GND.n2152 163.367
R15493 GND.n5673 GND.n2152 163.367
R15494 GND.n5673 GND.n2153 163.367
R15495 GND.n5669 GND.n2153 163.367
R15496 GND.n5669 GND.n2156 163.367
R15497 GND.n4508 GND.n2156 163.367
R15498 GND.n4508 GND.n2170 163.367
R15499 GND.n5659 GND.n2170 163.367
R15500 GND.n5659 GND.n2171 163.367
R15501 GND.n5655 GND.n2171 163.367
R15502 GND.n5655 GND.n2174 163.367
R15503 GND.n4532 GND.n2174 163.367
R15504 GND.n4532 GND.n4525 163.367
R15505 GND.n4528 GND.n4525 163.367
R15506 GND.n4528 GND.n4527 163.367
R15507 GND.n4527 GND.n2200 163.367
R15508 GND.n5638 GND.n2200 163.367
R15509 GND.n5638 GND.n2201 163.367
R15510 GND.n5634 GND.n2201 163.367
R15511 GND.n5634 GND.n2204 163.367
R15512 GND.n4551 GND.n2204 163.367
R15513 GND.n4551 GND.n2221 163.367
R15514 GND.n2231 GND.n2221 163.367
R15515 GND.n5619 GND.n2231 163.367
R15516 GND.n5619 GND.n2232 163.367
R15517 GND.n5615 GND.n2232 163.367
R15518 GND.n5615 GND.n2235 163.367
R15519 GND.n4592 GND.n2235 163.367
R15520 GND.n4592 GND.n2254 163.367
R15521 GND.n5605 GND.n2254 163.367
R15522 GND.n5605 GND.n2255 163.367
R15523 GND.n5601 GND.n2255 163.367
R15524 GND.n5601 GND.n2258 163.367
R15525 GND.n4648 GND.n2258 163.367
R15526 GND.n4648 GND.n4641 163.367
R15527 GND.n4644 GND.n4641 163.367
R15528 GND.n4644 GND.n4643 163.367
R15529 GND.n4643 GND.n2284 163.367
R15530 GND.n5584 GND.n2284 163.367
R15531 GND.n5584 GND.n2285 163.367
R15532 GND.n5580 GND.n2285 163.367
R15533 GND.n5580 GND.n2288 163.367
R15534 GND.n4687 GND.n2288 163.367
R15535 GND.n4688 GND.n4687 163.367
R15536 GND.n4688 GND.n2959 163.367
R15537 GND.n4692 GND.n2959 163.367
R15538 GND.n4692 GND.n2325 163.367
R15539 GND.n5563 GND.n2325 163.367
R15540 GND.n5563 GND.n2326 163.367
R15541 GND.n5559 GND.n2326 163.367
R15542 GND.n5559 GND.n2329 163.367
R15543 GND.n4712 GND.n2329 163.367
R15544 GND.n4712 GND.n2345 163.367
R15545 GND.n5549 GND.n2345 163.367
R15546 GND.n5549 GND.n2346 163.367
R15547 GND.n5545 GND.n2346 163.367
R15548 GND.n5545 GND.n2349 163.367
R15549 GND.n2944 GND.n2349 163.367
R15550 GND.n2944 GND.n2364 163.367
R15551 GND.n5535 GND.n2364 163.367
R15552 GND.n5535 GND.n2365 163.367
R15553 GND.n5531 GND.n2365 163.367
R15554 GND.n5531 GND.n2368 163.367
R15555 GND.n5475 GND.n2368 163.367
R15556 GND.n5475 GND.n2417 163.367
R15557 GND.n5471 GND.n2417 163.367
R15558 GND.n5471 GND.n2419 163.367
R15559 GND.n5463 GND.n2419 163.367
R15560 GND.n5463 GND.n2429 163.367
R15561 GND.n5459 GND.n2429 163.367
R15562 GND.n5459 GND.n2431 163.367
R15563 GND.n2465 GND.n2431 163.367
R15564 GND.n2407 GND.t98 161.207
R15565 GND.n4198 GND.t65 161.207
R15566 GND.n2495 GND.n2494 157.237
R15567 GND.n1867 GND.n1866 152
R15568 GND.n1868 GND.n1855 152
R15569 GND.n1870 GND.n1869 152
R15570 GND.n1873 GND.n1872 152
R15571 GND.n1874 GND.n1853 152
R15572 GND.n1876 GND.n1875 152
R15573 GND.n1878 GND.n1851 152
R15574 GND.n1880 GND.n1879 152
R15575 GND.n2493 GND.n2467 152
R15576 GND.n2483 GND.n2468 152
R15577 GND.n2482 GND.n2481 152
R15578 GND.n2480 GND.n2469 152
R15579 GND.n2477 GND.n2470 152
R15580 GND.n2476 GND.n2475 152
R15581 GND.n2474 GND.n2471 152
R15582 GND.n2472 GND.t134 149.72
R15583 GND.n2548 GND.n2455 143.351
R15584 GND.n5848 GND.n1824 143.351
R15585 GND.n1836 GND.n1824 143.351
R15586 GND.n1864 GND.t59 129.018
R15587 GND.n1879 GND.t78 126.766
R15588 GND.n1877 GND.t131 126.766
R15589 GND.n1853 GND.t66 126.766
R15590 GND.n1871 GND.t152 126.766
R15591 GND.n1855 GND.t87 126.766
R15592 GND.n1865 GND.t110 126.766
R15593 GND.n2473 GND.t84 126.766
R15594 GND.n2475 GND.t116 126.766
R15595 GND.n2479 GND.t107 126.766
R15596 GND.n2481 GND.t125 126.766
R15597 GND.n2492 GND.t75 126.766
R15598 GND.n2494 GND.t143 126.766
R15599 GND.n4869 GND.n4868 124.704
R15600 GND.n272 GND.n271 124.704
R15601 GND.n1746 GND.n1745 111.903
R15602 GND.n1801 GND.n1800 111.903
R15603 GND.n3117 GND.n3116 111.903
R15604 GND.n3106 GND.n3105 111.903
R15605 GND.n1821 GND.n1820 111.903
R15606 GND.n5349 GND.n5348 111.903
R15607 GND.n2553 GND.n2552 111.903
R15608 GND.n4827 GND.n4826 111.903
R15609 GND.n257 GND.n256 111.903
R15610 GND.n328 GND.n327 111.903
R15611 GND.n228 GND.n227 111.903
R15612 GND.n5113 GND.n5112 111.903
R15613 GND.n2900 GND.n2899 111.903
R15614 GND.n3520 GND.n3519 111.903
R15615 GND.n3510 GND.n3509 111.903
R15616 GND.n3616 GND.n3615 111.903
R15617 GND.n3650 GND.n3649 111.903
R15618 GND.n1665 GND.n1664 111.903
R15619 GND.n5810 GND.n5809 102.4
R15620 GND.n1909 GND.n1908 102.4
R15621 GND.n2501 GND.n2500 102.4
R15622 GND.n2499 GND.n2498 102.4
R15623 GND.n370 GND.n215 99.6594
R15624 GND.n368 GND.n214 99.6594
R15625 GND.n364 GND.n213 99.6594
R15626 GND.n360 GND.n212 99.6594
R15627 GND.n356 GND.n211 99.6594
R15628 GND.n352 GND.n210 99.6594
R15629 GND.n348 GND.n209 99.6594
R15630 GND.n344 GND.n208 99.6594
R15631 GND.n340 GND.n207 99.6594
R15632 GND.n336 GND.n206 99.6594
R15633 GND.n332 GND.n205 99.6594
R15634 GND.n325 GND.n204 99.6594
R15635 GND.n321 GND.n203 99.6594
R15636 GND.n317 GND.n202 99.6594
R15637 GND.n313 GND.n201 99.6594
R15638 GND.n309 GND.n200 99.6594
R15639 GND.n305 GND.n199 99.6594
R15640 GND.n259 GND.n198 99.6594
R15641 GND.n297 GND.n197 99.6594
R15642 GND.n293 GND.n196 99.6594
R15643 GND.n289 GND.n195 99.6594
R15644 GND.n285 GND.n194 99.6594
R15645 GND.n281 GND.n193 99.6594
R15646 GND.n277 GND.n192 99.6594
R15647 GND.n191 GND.n180 99.6594
R15648 GND.n5403 GND.n5402 99.6594
R15649 GND.n5397 GND.n2558 99.6594
R15650 GND.n5394 GND.n2559 99.6594
R15651 GND.n5390 GND.n2560 99.6594
R15652 GND.n5386 GND.n2561 99.6594
R15653 GND.n5382 GND.n2562 99.6594
R15654 GND.n5378 GND.n2563 99.6594
R15655 GND.n5374 GND.n2564 99.6594
R15656 GND.n5370 GND.n2565 99.6594
R15657 GND.n5366 GND.n2566 99.6594
R15658 GND.n5362 GND.n2567 99.6594
R15659 GND.n2568 GND.n2556 99.6594
R15660 GND.n4844 GND.n2569 99.6594
R15661 GND.n4846 GND.n2570 99.6594
R15662 GND.n4854 GND.n2571 99.6594
R15663 GND.n4856 GND.n2572 99.6594
R15664 GND.n4864 GND.n2573 99.6594
R15665 GND.n4866 GND.n2574 99.6594
R15666 GND.n4876 GND.n2575 99.6594
R15667 GND.n4878 GND.n2576 99.6594
R15668 GND.n4886 GND.n2577 99.6594
R15669 GND.n4888 GND.n2578 99.6594
R15670 GND.n4896 GND.n2579 99.6594
R15671 GND.n4898 GND.n2580 99.6594
R15672 GND.n1787 GND.n1781 99.6594
R15673 GND.n1789 GND.n1780 99.6594
R15674 GND.n1793 GND.n1779 99.6594
R15675 GND.n1795 GND.n1778 99.6594
R15676 GND.n1799 GND.n1777 99.6594
R15677 GND.n1803 GND.n1776 99.6594
R15678 GND.n1807 GND.n1775 99.6594
R15679 GND.n1809 GND.n1774 99.6594
R15680 GND.n1813 GND.n1773 99.6594
R15681 GND.n1815 GND.n1772 99.6594
R15682 GND.n3130 GND.n1770 99.6594
R15683 GND.n3135 GND.n1769 99.6594
R15684 GND.n3127 GND.n1768 99.6594
R15685 GND.n3143 GND.n1767 99.6594
R15686 GND.n3123 GND.n1766 99.6594
R15687 GND.n3151 GND.n1765 99.6594
R15688 GND.n3119 GND.n1764 99.6594
R15689 GND.n3159 GND.n1763 99.6594
R15690 GND.n3113 GND.n1762 99.6594
R15691 GND.n3167 GND.n1761 99.6594
R15692 GND.n3109 GND.n1760 99.6594
R15693 GND.n3175 GND.n1759 99.6594
R15694 GND.n3181 GND.n1758 99.6594
R15695 GND.n3185 GND.n1757 99.6594
R15696 GND.n3483 GND.n1615 99.6594
R15697 GND.n3530 GND.n1616 99.6594
R15698 GND.n3536 GND.n1617 99.6594
R15699 GND.n3540 GND.n1618 99.6594
R15700 GND.n3546 GND.n1619 99.6594
R15701 GND.n3550 GND.n1620 99.6594
R15702 GND.n3556 GND.n1621 99.6594
R15703 GND.n3558 GND.n1622 99.6594
R15704 GND.n3566 GND.n1623 99.6594
R15705 GND.n3568 GND.n1624 99.6594
R15706 GND.n3576 GND.n1625 99.6594
R15707 GND.n3578 GND.n1626 99.6594
R15708 GND.n3586 GND.n1627 99.6594
R15709 GND.n3590 GND.n1628 99.6594
R15710 GND.n3596 GND.n1629 99.6594
R15711 GND.n3600 GND.n1630 99.6594
R15712 GND.n3606 GND.n1631 99.6594
R15713 GND.n3610 GND.n1632 99.6594
R15714 GND.n3503 GND.n1633 99.6594
R15715 GND.n3620 GND.n1634 99.6594
R15716 GND.n3626 GND.n1635 99.6594
R15717 GND.n3630 GND.n1636 99.6594
R15718 GND.n3636 GND.n1637 99.6594
R15719 GND.n3640 GND.n1638 99.6594
R15720 GND.n3646 GND.n1639 99.6594
R15721 GND.n5520 GND.n5519 99.6594
R15722 GND.n5515 GND.n2388 99.6594
R15723 GND.n5511 GND.n2387 99.6594
R15724 GND.n5507 GND.n2386 99.6594
R15725 GND.n5503 GND.n2385 99.6594
R15726 GND.n5499 GND.n2384 99.6594
R15727 GND.n5495 GND.n2383 99.6594
R15728 GND.n5491 GND.n2382 99.6594
R15729 GND.n5487 GND.n2381 99.6594
R15730 GND.n5483 GND.n2380 99.6594
R15731 GND.n5479 GND.n2379 99.6594
R15732 GND.n4247 GND.n3081 99.6594
R15733 GND.n4245 GND.n3084 99.6594
R15734 GND.n4241 GND.n4240 99.6594
R15735 GND.n4234 GND.n3089 99.6594
R15736 GND.n4233 GND.n4232 99.6594
R15737 GND.n4153 GND.n3095 99.6594
R15738 GND.n4164 GND.n4155 99.6594
R15739 GND.n4167 GND.n4166 99.6594
R15740 GND.n4176 GND.n4175 99.6594
R15741 GND.n4185 GND.n4178 99.6594
R15742 GND.n4188 GND.n4187 99.6594
R15743 GND.n5129 GND.n5123 99.6594
R15744 GND.n5133 GND.n5131 99.6594
R15745 GND.n5139 GND.n5119 99.6594
R15746 GND.n5143 GND.n5141 99.6594
R15747 GND.n5149 GND.n5115 99.6594
R15748 GND.n5152 GND.n5151 99.6594
R15749 GND.n2902 GND.n2581 99.6594
R15750 GND.n2908 GND.n2582 99.6594
R15751 GND.n2914 GND.n2583 99.6594
R15752 GND.n2920 GND.n2584 99.6594
R15753 GND.n2926 GND.n2585 99.6594
R15754 GND.n2897 GND.n2586 99.6594
R15755 GND.n2907 GND.n2581 99.6594
R15756 GND.n2913 GND.n2582 99.6594
R15757 GND.n2919 GND.n2583 99.6594
R15758 GND.n2925 GND.n2584 99.6594
R15759 GND.n2928 GND.n2585 99.6594
R15760 GND.n4801 GND.n2586 99.6594
R15761 GND.n5151 GND.n5150 99.6594
R15762 GND.n5142 GND.n5115 99.6594
R15763 GND.n5141 GND.n5140 99.6594
R15764 GND.n5132 GND.n5119 99.6594
R15765 GND.n5131 GND.n5130 99.6594
R15766 GND.n5124 GND.n5123 99.6594
R15767 GND.n4248 GND.n4247 99.6594
R15768 GND.n4242 GND.n3084 99.6594
R15769 GND.n4240 GND.n4239 99.6594
R15770 GND.n4235 GND.n4234 99.6594
R15771 GND.n4232 GND.n4231 99.6594
R15772 GND.n4154 GND.n4153 99.6594
R15773 GND.n4165 GND.n4164 99.6594
R15774 GND.n4168 GND.n4167 99.6594
R15775 GND.n4177 GND.n4176 99.6594
R15776 GND.n4186 GND.n4185 99.6594
R15777 GND.n4187 GND.n3079 99.6594
R15778 GND.n5482 GND.n2379 99.6594
R15779 GND.n5486 GND.n2380 99.6594
R15780 GND.n5490 GND.n2381 99.6594
R15781 GND.n5494 GND.n2382 99.6594
R15782 GND.n5498 GND.n2383 99.6594
R15783 GND.n5502 GND.n2384 99.6594
R15784 GND.n5506 GND.n2385 99.6594
R15785 GND.n5510 GND.n2386 99.6594
R15786 GND.n5514 GND.n2387 99.6594
R15787 GND.n2389 GND.n2388 99.6594
R15788 GND.n5520 GND.n2377 99.6594
R15789 GND.n3529 GND.n1615 99.6594
R15790 GND.n3535 GND.n1616 99.6594
R15791 GND.n3539 GND.n1617 99.6594
R15792 GND.n3545 GND.n1618 99.6594
R15793 GND.n3549 GND.n1619 99.6594
R15794 GND.n3555 GND.n1620 99.6594
R15795 GND.n3559 GND.n1621 99.6594
R15796 GND.n3565 GND.n1622 99.6594
R15797 GND.n3569 GND.n1623 99.6594
R15798 GND.n3575 GND.n1624 99.6594
R15799 GND.n3579 GND.n1625 99.6594
R15800 GND.n3585 GND.n1626 99.6594
R15801 GND.n3589 GND.n1627 99.6594
R15802 GND.n3595 GND.n1628 99.6594
R15803 GND.n3599 GND.n1629 99.6594
R15804 GND.n3605 GND.n1630 99.6594
R15805 GND.n3609 GND.n1631 99.6594
R15806 GND.n3502 GND.n1632 99.6594
R15807 GND.n3619 GND.n1633 99.6594
R15808 GND.n3625 GND.n1634 99.6594
R15809 GND.n3629 GND.n1635 99.6594
R15810 GND.n3635 GND.n1636 99.6594
R15811 GND.n3639 GND.n1637 99.6594
R15812 GND.n3645 GND.n1638 99.6594
R15813 GND.n3648 GND.n1639 99.6594
R15814 GND.n3182 GND.n1757 99.6594
R15815 GND.n3176 GND.n1758 99.6594
R15816 GND.n3110 GND.n1759 99.6594
R15817 GND.n3168 GND.n1760 99.6594
R15818 GND.n3114 GND.n1761 99.6594
R15819 GND.n3160 GND.n1762 99.6594
R15820 GND.n3120 GND.n1763 99.6594
R15821 GND.n3152 GND.n1764 99.6594
R15822 GND.n3124 GND.n1765 99.6594
R15823 GND.n3144 GND.n1766 99.6594
R15824 GND.n3128 GND.n1767 99.6594
R15825 GND.n3136 GND.n1768 99.6594
R15826 GND.n3131 GND.n1769 99.6594
R15827 GND.n1816 GND.n1771 99.6594
R15828 GND.n1814 GND.n1772 99.6594
R15829 GND.n1810 GND.n1773 99.6594
R15830 GND.n1808 GND.n1774 99.6594
R15831 GND.n1804 GND.n1775 99.6594
R15832 GND.n1802 GND.n1776 99.6594
R15833 GND.n1796 GND.n1777 99.6594
R15834 GND.n1794 GND.n1778 99.6594
R15835 GND.n1790 GND.n1779 99.6594
R15836 GND.n1788 GND.n1780 99.6594
R15837 GND.n1783 GND.n1781 99.6594
R15838 GND.n5403 GND.n2589 99.6594
R15839 GND.n5395 GND.n2558 99.6594
R15840 GND.n5391 GND.n2559 99.6594
R15841 GND.n5387 GND.n2560 99.6594
R15842 GND.n5383 GND.n2561 99.6594
R15843 GND.n5379 GND.n2562 99.6594
R15844 GND.n5375 GND.n2563 99.6594
R15845 GND.n5371 GND.n2564 99.6594
R15846 GND.n5367 GND.n2565 99.6594
R15847 GND.n5363 GND.n2566 99.6594
R15848 GND.n5406 GND.n5405 99.6594
R15849 GND.n4843 GND.n2568 99.6594
R15850 GND.n4847 GND.n2569 99.6594
R15851 GND.n4853 GND.n2570 99.6594
R15852 GND.n4857 GND.n2571 99.6594
R15853 GND.n4863 GND.n2572 99.6594
R15854 GND.n4867 GND.n2573 99.6594
R15855 GND.n4875 GND.n2574 99.6594
R15856 GND.n4879 GND.n2575 99.6594
R15857 GND.n4885 GND.n2576 99.6594
R15858 GND.n4889 GND.n2577 99.6594
R15859 GND.n4895 GND.n2578 99.6594
R15860 GND.n4899 GND.n2579 99.6594
R15861 GND.n4907 GND.n2580 99.6594
R15862 GND.n276 GND.n191 99.6594
R15863 GND.n280 GND.n192 99.6594
R15864 GND.n284 GND.n193 99.6594
R15865 GND.n288 GND.n194 99.6594
R15866 GND.n292 GND.n195 99.6594
R15867 GND.n296 GND.n196 99.6594
R15868 GND.n258 GND.n197 99.6594
R15869 GND.n304 GND.n198 99.6594
R15870 GND.n308 GND.n199 99.6594
R15871 GND.n312 GND.n200 99.6594
R15872 GND.n316 GND.n201 99.6594
R15873 GND.n320 GND.n202 99.6594
R15874 GND.n324 GND.n203 99.6594
R15875 GND.n331 GND.n204 99.6594
R15876 GND.n335 GND.n205 99.6594
R15877 GND.n339 GND.n206 99.6594
R15878 GND.n343 GND.n207 99.6594
R15879 GND.n347 GND.n208 99.6594
R15880 GND.n351 GND.n209 99.6594
R15881 GND.n355 GND.n210 99.6594
R15882 GND.n359 GND.n211 99.6594
R15883 GND.n363 GND.n212 99.6594
R15884 GND.n367 GND.n213 99.6594
R15885 GND.n371 GND.n214 99.6594
R15886 GND.n216 GND.n215 99.6594
R15887 GND.n1649 GND.n1641 99.6594
R15888 GND.n1654 GND.n1642 99.6594
R15889 GND.n1656 GND.n1643 99.6594
R15890 GND.n1660 GND.n1644 99.6594
R15891 GND.n1662 GND.n1645 99.6594
R15892 GND.n1653 GND.n1641 99.6594
R15893 GND.n1655 GND.n1642 99.6594
R15894 GND.n1659 GND.n1643 99.6594
R15895 GND.n1661 GND.n1644 99.6594
R15896 GND.n1663 GND.n1645 99.6594
R15897 GND.n4221 GND.n1751 99.6594
R15898 GND.n4159 GND.n1752 99.6594
R15899 GND.n4161 GND.n1753 99.6594
R15900 GND.n4172 GND.n1754 99.6594
R15901 GND.n4182 GND.n1755 99.6594
R15902 GND.n5890 GND.n1749 99.6594
R15903 GND.n5891 GND.n5890 99.6594
R15904 GND.n4183 GND.n1755 99.6594
R15905 GND.n4181 GND.n1754 99.6594
R15906 GND.n4171 GND.n1753 99.6594
R15907 GND.n4160 GND.n1752 99.6594
R15908 GND.n4158 GND.n1751 99.6594
R15909 GND.n11 GND.t30 97.7611
R15910 GND.n11 GND.t28 96.5537
R15911 GND.n1864 GND.n1863 83.3186
R15912 GND.n2408 GND.n2407 82.6187
R15913 GND.n4199 GND.n4198 82.6187
R15914 GND.n1909 GND.t147 78.6838
R15915 GND.n2501 GND.t103 78.6838
R15916 GND.n5810 GND.t43 78.6836
R15917 GND.n2499 GND.t139 78.6836
R15918 GND.n2408 GND.t99 78.5881
R15919 GND.n4199 GND.t64 78.5881
R15920 GND.n1 GND.t22 74.2965
R15921 GND.n2 GND.t14 74.2965
R15922 GND.n4 GND.t20 74.2965
R15923 GND.n6 GND.t18 74.2965
R15924 GND.n0 GND.t9 74.2965
R15925 GND.n13 GND.t10 74.2965
R15926 GND.n14 GND.t3 74.2965
R15927 GND.n16 GND.t6 74.2965
R15928 GND.n18 GND.t21 74.2965
R15929 GND.n20 GND.t11 74.2965
R15930 GND.n1865 GND.n1856 72.8411
R15931 GND.n1871 GND.n1854 72.8411
R15932 GND.n1877 GND.n1852 72.8411
R15933 GND.n2492 GND.n2491 72.8411
R15934 GND.n2479 GND.n2478 72.8411
R15935 GND.n6350 GND.n1266 72.812
R15936 GND.n6350 GND.n6349 72.812
R15937 GND.n6349 GND.n6348 72.812
R15938 GND.n6348 GND.n1271 72.812
R15939 GND.n6342 GND.n1271 72.812
R15940 GND.n6342 GND.n6341 72.812
R15941 GND.n6341 GND.n6340 72.812
R15942 GND.n6340 GND.n1279 72.812
R15943 GND.n6334 GND.n1279 72.812
R15944 GND.n6334 GND.n6333 72.812
R15945 GND.n6333 GND.n6332 72.812
R15946 GND.n6332 GND.n1287 72.812
R15947 GND.n6326 GND.n1287 72.812
R15948 GND.n6326 GND.n6325 72.812
R15949 GND.n6325 GND.n6324 72.812
R15950 GND.n6324 GND.n1295 72.812
R15951 GND.n6318 GND.n1295 72.812
R15952 GND.n6318 GND.n6317 72.812
R15953 GND.n6317 GND.n6316 72.812
R15954 GND.n6316 GND.n1303 72.812
R15955 GND.n6310 GND.n1303 72.812
R15956 GND.n6310 GND.n6309 72.812
R15957 GND.n6309 GND.n6308 72.812
R15958 GND.n6308 GND.n1311 72.812
R15959 GND.n6302 GND.n1311 72.812
R15960 GND.n6302 GND.n6301 72.812
R15961 GND.n6301 GND.n6300 72.812
R15962 GND.n6300 GND.n1319 72.812
R15963 GND.n6294 GND.n1319 72.812
R15964 GND.n6294 GND.n6293 72.812
R15965 GND.n6293 GND.n6292 72.812
R15966 GND.n6292 GND.n1327 72.812
R15967 GND.n6286 GND.n1327 72.812
R15968 GND.n6286 GND.n6285 72.812
R15969 GND.n6285 GND.n6284 72.812
R15970 GND.n6284 GND.n1335 72.812
R15971 GND.n6278 GND.n1335 72.812
R15972 GND.n6278 GND.n6277 72.812
R15973 GND.n6277 GND.n6276 72.812
R15974 GND.n6276 GND.n1343 72.812
R15975 GND.n6270 GND.n1343 72.812
R15976 GND.n6270 GND.n6269 72.812
R15977 GND.n6269 GND.n6268 72.812
R15978 GND.n6268 GND.n1351 72.812
R15979 GND.n6262 GND.n1351 72.812
R15980 GND.n6262 GND.n6261 72.812
R15981 GND.n6261 GND.n6260 72.812
R15982 GND.n6260 GND.n1359 72.812
R15983 GND.n6254 GND.n1359 72.812
R15984 GND.n6254 GND.n6253 72.812
R15985 GND.n6253 GND.n6252 72.812
R15986 GND.n6252 GND.n1367 72.812
R15987 GND.n6246 GND.n1367 72.812
R15988 GND.n6246 GND.n6245 72.812
R15989 GND.n6245 GND.n6244 72.812
R15990 GND.n6244 GND.n1375 72.812
R15991 GND.n6238 GND.n1375 72.812
R15992 GND.n6238 GND.n6237 72.812
R15993 GND.n6237 GND.n6236 72.812
R15994 GND.n6236 GND.n1383 72.812
R15995 GND.n6230 GND.n1383 72.812
R15996 GND.n6230 GND.n6229 72.812
R15997 GND.n6229 GND.n6228 72.812
R15998 GND.n6228 GND.n1391 72.812
R15999 GND.n6222 GND.n1391 72.812
R16000 GND.n6222 GND.n6221 72.812
R16001 GND.n6221 GND.n6220 72.812
R16002 GND.n6220 GND.n1399 72.812
R16003 GND.n6214 GND.n1399 72.812
R16004 GND.n6214 GND.n6213 72.812
R16005 GND.n6213 GND.n6212 72.812
R16006 GND.n6212 GND.n1407 72.812
R16007 GND.n6206 GND.n1407 72.812
R16008 GND.n6206 GND.n6205 72.812
R16009 GND.n6205 GND.n6204 72.812
R16010 GND.n6204 GND.n1415 72.812
R16011 GND.n6198 GND.n1415 72.812
R16012 GND.n6198 GND.n6197 72.812
R16013 GND.n6197 GND.n6196 72.812
R16014 GND.n6196 GND.n1423 72.812
R16015 GND.n6190 GND.n1423 72.812
R16016 GND.n6190 GND.n6189 72.812
R16017 GND.n6189 GND.n6188 72.812
R16018 GND.n6188 GND.n1431 72.812
R16019 GND.n6182 GND.n1431 72.812
R16020 GND.n6182 GND.n6181 72.812
R16021 GND.n6181 GND.n6180 72.812
R16022 GND.n6180 GND.n1439 72.812
R16023 GND.n6174 GND.n1439 72.812
R16024 GND.n1 GND.t1 72.4488
R16025 GND.n2 GND.t17 72.4488
R16026 GND.n4 GND.t23 72.4488
R16027 GND.n6 GND.t16 72.4488
R16028 GND.n0 GND.t7 72.4488
R16029 GND.n13 GND.t15 72.4488
R16030 GND.n14 GND.t5 72.4488
R16031 GND.n16 GND.t13 72.4488
R16032 GND.n18 GND.t19 72.4488
R16033 GND.n20 GND.t12 72.4488
R16034 GND.n5445 GND.n2464 71.676
R16035 GND.n5441 GND.n2463 71.676
R16036 GND.n5437 GND.n2462 71.676
R16037 GND.n5433 GND.n2461 71.676
R16038 GND.n5429 GND.n2460 71.676
R16039 GND.n5425 GND.n2459 71.676
R16040 GND.n5421 GND.n2458 71.676
R16041 GND.n5416 GND.n2457 71.676
R16042 GND.n5412 GND.n2456 71.676
R16043 GND.n2548 GND.n2444 71.676
R16044 GND.n2544 GND.n2445 71.676
R16045 GND.n2540 GND.n2446 71.676
R16046 GND.n2536 GND.n2447 71.676
R16047 GND.n2532 GND.n2448 71.676
R16048 GND.n2528 GND.n2449 71.676
R16049 GND.n2524 GND.n2450 71.676
R16050 GND.n2520 GND.n2451 71.676
R16051 GND.n2516 GND.n2452 71.676
R16052 GND.n2512 GND.n2453 71.676
R16053 GND.n2508 GND.n2454 71.676
R16054 GND.n5846 GND.n5845 71.676
R16055 GND.n5840 GND.n1828 71.676
R16056 GND.n5837 GND.n1829 71.676
R16057 GND.n5833 GND.n1830 71.676
R16058 GND.n5829 GND.n1831 71.676
R16059 GND.n5825 GND.n1832 71.676
R16060 GND.n5821 GND.n1833 71.676
R16061 GND.n5817 GND.n1834 71.676
R16062 GND.n5812 GND.n1835 71.676
R16063 GND.n5849 GND.n5848 71.676
R16064 GND.n1911 GND.n1837 71.676
R16065 GND.n1915 GND.n1838 71.676
R16066 GND.n1920 GND.n1839 71.676
R16067 GND.n1924 GND.n1840 71.676
R16068 GND.n1928 GND.n1841 71.676
R16069 GND.n1932 GND.n1842 71.676
R16070 GND.n1936 GND.n1843 71.676
R16071 GND.n1940 GND.n1844 71.676
R16072 GND.n1944 GND.n1845 71.676
R16073 GND.n5846 GND.n1849 71.676
R16074 GND.n5838 GND.n1828 71.676
R16075 GND.n5834 GND.n1829 71.676
R16076 GND.n5830 GND.n1830 71.676
R16077 GND.n5826 GND.n1831 71.676
R16078 GND.n5822 GND.n1832 71.676
R16079 GND.n5818 GND.n1833 71.676
R16080 GND.n5813 GND.n1834 71.676
R16081 GND.n1835 GND.n1826 71.676
R16082 GND.n1910 GND.n1836 71.676
R16083 GND.n1914 GND.n1837 71.676
R16084 GND.n1919 GND.n1838 71.676
R16085 GND.n1923 GND.n1839 71.676
R16086 GND.n1927 GND.n1840 71.676
R16087 GND.n1931 GND.n1841 71.676
R16088 GND.n1935 GND.n1842 71.676
R16089 GND.n1939 GND.n1843 71.676
R16090 GND.n1943 GND.n1844 71.676
R16091 GND.n1946 GND.n1845 71.676
R16092 GND.n2511 GND.n2454 71.676
R16093 GND.n2515 GND.n2453 71.676
R16094 GND.n2519 GND.n2452 71.676
R16095 GND.n2523 GND.n2451 71.676
R16096 GND.n2527 GND.n2450 71.676
R16097 GND.n2531 GND.n2449 71.676
R16098 GND.n2535 GND.n2448 71.676
R16099 GND.n2539 GND.n2447 71.676
R16100 GND.n2543 GND.n2446 71.676
R16101 GND.n2546 GND.n2445 71.676
R16102 GND.n5411 GND.n2455 71.676
R16103 GND.n5415 GND.n2456 71.676
R16104 GND.n5420 GND.n2457 71.676
R16105 GND.n5424 GND.n2458 71.676
R16106 GND.n5428 GND.n2459 71.676
R16107 GND.n5432 GND.n2460 71.676
R16108 GND.n5436 GND.n2461 71.676
R16109 GND.n5440 GND.n2462 71.676
R16110 GND.n5444 GND.n2463 71.676
R16111 GND.n2466 GND.n2464 71.676
R16112 GND.n1746 GND.t130 67.5836
R16113 GND.n1801 GND.t83 67.5836
R16114 GND.n3117 GND.t58 67.5836
R16115 GND.n3106 GND.t157 67.5836
R16116 GND.n1821 GND.t160 67.5836
R16117 GND.n5349 GND.t49 67.5836
R16118 GND.n2553 GND.t141 67.5836
R16119 GND.n4827 GND.t120 67.5836
R16120 GND.n257 GND.t74 67.5836
R16121 GND.n328 GND.t47 67.5836
R16122 GND.n228 GND.t92 67.5836
R16123 GND.n5113 GND.t36 67.5836
R16124 GND.n2900 GND.t105 67.5836
R16125 GND.n3520 GND.t114 67.5836
R16126 GND.n3510 GND.t53 67.5836
R16127 GND.n3616 GND.t94 67.5836
R16128 GND.n3650 GND.t150 67.5836
R16129 GND.n1665 GND.t123 67.5836
R16130 GND.n4869 GND.t39 64.3836
R16131 GND.n272 GND.t71 64.3836
R16132 GND.n5808 GND.n1880 58.4046
R16133 GND.n1862 GND.n1861 54.358
R16134 GND.n2489 GND.n2488 54.358
R16135 GND.n5815 GND.n5810 53.1399
R16136 GND.n1917 GND.n1909 53.1399
R16137 GND.n2502 GND.n2501 53.1399
R16138 GND.n5418 GND.n2499 53.1399
R16139 GND.n2472 GND.n2471 52.3702
R16140 GND.n4870 GND.n4869 48.6793
R16141 GND.n275 GND.n272 48.6793
R16142 GND.n1865 GND.n1864 45.8904
R16143 GND.n2497 GND.n2495 44.3322
R16144 GND.n1878 GND.n1877 43.8187
R16145 GND.n2493 GND.n2492 43.8187
R16146 GND.n1863 GND.n1862 41.6274
R16147 GND.n2490 GND.n2489 41.6274
R16148 GND.n1872 GND.n1871 37.9763
R16149 GND.n1871 GND.n1870 37.9763
R16150 GND.n2479 GND.n2470 37.9763
R16151 GND.n2480 GND.n2479 37.9763
R16152 GND.n6173 GND.n6172 36.7959
R16153 GND.n6172 GND.n1446 36.7959
R16154 GND.n6166 GND.n1446 36.7959
R16155 GND.n6166 GND.n6165 36.7959
R16156 GND.n6165 GND.n6164 36.7959
R16157 GND.n6164 GND.n1455 36.7959
R16158 GND.n6158 GND.n1455 36.7959
R16159 GND.n6158 GND.n6157 36.7959
R16160 GND.n6157 GND.n6156 36.7959
R16161 GND.n6156 GND.n1463 36.7959
R16162 GND.n6150 GND.n1463 36.7959
R16163 GND.n6150 GND.n6149 36.7959
R16164 GND.n6149 GND.n6148 36.7959
R16165 GND.n6148 GND.n1471 36.7959
R16166 GND.n6142 GND.n1471 36.7959
R16167 GND.n6142 GND.n6141 36.7959
R16168 GND.n6141 GND.n6140 36.7959
R16169 GND.n6140 GND.n1479 36.7959
R16170 GND.n6134 GND.n1479 36.7959
R16171 GND.n6134 GND.n6133 36.7959
R16172 GND.n6133 GND.n6132 36.7959
R16173 GND.n6132 GND.n1487 36.7959
R16174 GND.n6126 GND.n1487 36.7959
R16175 GND.n6126 GND.n6125 36.7959
R16176 GND.n6125 GND.n6124 36.7959
R16177 GND.n6124 GND.n1495 36.7959
R16178 GND.n6118 GND.n1495 36.7959
R16179 GND.n6118 GND.n6117 36.7959
R16180 GND.n6117 GND.n6116 36.7959
R16181 GND.n6116 GND.n1503 36.7959
R16182 GND.n6110 GND.n1503 36.7959
R16183 GND.n6110 GND.n6109 36.7959
R16184 GND.n6109 GND.n6108 36.7959
R16185 GND.n6108 GND.n1511 36.7959
R16186 GND.n6102 GND.n1511 36.7959
R16187 GND.n6102 GND.n6101 36.7959
R16188 GND.n6101 GND.n6100 36.7959
R16189 GND.n6100 GND.n1519 36.7959
R16190 GND.n6094 GND.n1519 36.7959
R16191 GND.n6094 GND.n6093 36.7959
R16192 GND.n6093 GND.n6092 36.7959
R16193 GND.n6092 GND.n1527 36.7959
R16194 GND.n6086 GND.n1527 36.7959
R16195 GND.n6086 GND.n6085 36.7959
R16196 GND.n6085 GND.n6084 36.7959
R16197 GND.n6084 GND.n1535 36.7959
R16198 GND.n6078 GND.n1535 36.7959
R16199 GND.n6078 GND.n6077 36.7959
R16200 GND.n6077 GND.n6076 36.7959
R16201 GND.n6076 GND.n1543 36.7959
R16202 GND.n6070 GND.n1543 36.7959
R16203 GND.n6070 GND.n6069 36.7959
R16204 GND.n6069 GND.n6068 36.7959
R16205 GND.n6068 GND.n1551 36.7959
R16206 GND.n6062 GND.n1551 36.7959
R16207 GND.n6062 GND.n6061 36.7959
R16208 GND.n6061 GND.n6060 36.7959
R16209 GND.n6060 GND.n1559 36.7959
R16210 GND.n6054 GND.n1559 36.7959
R16211 GND.n6054 GND.n6053 36.7959
R16212 GND.n6053 GND.n6052 36.7959
R16213 GND.n6052 GND.n1567 36.7959
R16214 GND.n6046 GND.n1567 36.7959
R16215 GND.n6046 GND.n6045 36.7959
R16216 GND.n6045 GND.n6044 36.7959
R16217 GND.n6044 GND.n1575 36.7959
R16218 GND.n6038 GND.n1575 36.7959
R16219 GND.n6038 GND.n6037 36.7959
R16220 GND.n6037 GND.n6036 36.7959
R16221 GND.n6036 GND.n1583 36.7959
R16222 GND.n6030 GND.n1583 36.7959
R16223 GND.n6030 GND.n6029 36.7959
R16224 GND.n6029 GND.n6028 36.7959
R16225 GND.n6028 GND.n1591 36.7959
R16226 GND.n6022 GND.n1591 36.7959
R16227 GND.n6022 GND.n6021 36.7959
R16228 GND.n6021 GND.n6020 36.7959
R16229 GND.n6020 GND.n1599 36.7959
R16230 GND.n6014 GND.n1599 36.7959
R16231 GND.n6014 GND.n6013 36.7959
R16232 GND.n6013 GND.n6012 36.7959
R16233 GND.n6012 GND.n1607 36.7959
R16234 GND.n6006 GND.n1607 36.7959
R16235 GND.n6006 GND.n6005 36.7959
R16236 GND.n3491 GND.n1647 36.7959
R16237 GND.n3187 GND.n1750 36.7959
R16238 GND.n4114 GND.n1756 36.7959
R16239 GND.n4114 GND.n4113 36.7959
R16240 GND.n4113 GND.n1827 36.7959
R16241 GND.n5451 GND.n2443 36.7959
R16242 GND.n4812 GND.n4811 36.7959
R16243 GND.n4813 GND.n4812 36.7959
R16244 GND.n4813 GND.n2557 36.7959
R16245 GND.n4825 GND.n2587 36.7959
R16246 GND.n7737 GND.n182 36.7959
R16247 GND.n7731 GND.n7730 36.7959
R16248 GND.n7730 GND.n7729 36.7959
R16249 GND.n7729 GND.n380 36.7959
R16250 GND.n7723 GND.n380 36.7959
R16251 GND.n7723 GND.n7722 36.7959
R16252 GND.n7722 GND.n7721 36.7959
R16253 GND.n7721 GND.n388 36.7959
R16254 GND.n7715 GND.n388 36.7959
R16255 GND.n7715 GND.n7714 36.7959
R16256 GND.n7714 GND.n7713 36.7959
R16257 GND.n7713 GND.n396 36.7959
R16258 GND.n7707 GND.n396 36.7959
R16259 GND.n7707 GND.n7706 36.7959
R16260 GND.n7706 GND.n7705 36.7959
R16261 GND.n7705 GND.n404 36.7959
R16262 GND.n7699 GND.n404 36.7959
R16263 GND.n7699 GND.n7698 36.7959
R16264 GND.n7698 GND.n7697 36.7959
R16265 GND.n7697 GND.n412 36.7959
R16266 GND.n7691 GND.n412 36.7959
R16267 GND.n7691 GND.n7690 36.7959
R16268 GND.n7690 GND.n7689 36.7959
R16269 GND.n7689 GND.n420 36.7959
R16270 GND.n7683 GND.n420 36.7959
R16271 GND.n7683 GND.n7682 36.7959
R16272 GND.n7682 GND.n7681 36.7959
R16273 GND.n7681 GND.n428 36.7959
R16274 GND.n7675 GND.n428 36.7959
R16275 GND.n7675 GND.n7674 36.7959
R16276 GND.n7674 GND.n7673 36.7959
R16277 GND.n7673 GND.n436 36.7959
R16278 GND.n7667 GND.n436 36.7959
R16279 GND.n7667 GND.n7666 36.7959
R16280 GND.n7666 GND.n7665 36.7959
R16281 GND.n7665 GND.n444 36.7959
R16282 GND.n7659 GND.n444 36.7959
R16283 GND.n7659 GND.n7658 36.7959
R16284 GND.n7658 GND.n7657 36.7959
R16285 GND.n7657 GND.n452 36.7959
R16286 GND.n7651 GND.n452 36.7959
R16287 GND.n7651 GND.n7650 36.7959
R16288 GND.n7650 GND.n7649 36.7959
R16289 GND.n7649 GND.n460 36.7959
R16290 GND.n7643 GND.n460 36.7959
R16291 GND.n7643 GND.n7642 36.7959
R16292 GND.n7642 GND.n7641 36.7959
R16293 GND.n7641 GND.n468 36.7959
R16294 GND.n7635 GND.n468 36.7959
R16295 GND.n7635 GND.n7634 36.7959
R16296 GND.n7634 GND.n7633 36.7959
R16297 GND.n7633 GND.n476 36.7959
R16298 GND.n7627 GND.n476 36.7959
R16299 GND.n7627 GND.n7626 36.7959
R16300 GND.n7626 GND.n7625 36.7959
R16301 GND.n7625 GND.n484 36.7959
R16302 GND.n7619 GND.n484 36.7959
R16303 GND.n7619 GND.n7618 36.7959
R16304 GND.n7618 GND.n7617 36.7959
R16305 GND.n7617 GND.n492 36.7959
R16306 GND.n7611 GND.n492 36.7959
R16307 GND.n7611 GND.n7610 36.7959
R16308 GND.n7610 GND.n7609 36.7959
R16309 GND.n7609 GND.n500 36.7959
R16310 GND.n7603 GND.n500 36.7959
R16311 GND.n7603 GND.n7602 36.7959
R16312 GND.n7602 GND.n7601 36.7959
R16313 GND.n7601 GND.n508 36.7959
R16314 GND.n7595 GND.n508 36.7959
R16315 GND.n7595 GND.n7594 36.7959
R16316 GND.n7594 GND.n7593 36.7959
R16317 GND.n7593 GND.n516 36.7959
R16318 GND.n7587 GND.n516 36.7959
R16319 GND.n7587 GND.n7586 36.7959
R16320 GND.n7586 GND.n7585 36.7959
R16321 GND.n7585 GND.n524 36.7959
R16322 GND.n7579 GND.n524 36.7959
R16323 GND.n7579 GND.n7578 36.7959
R16324 GND.n7578 GND.n7577 36.7959
R16325 GND.n7577 GND.n532 36.7959
R16326 GND.n7571 GND.n532 36.7959
R16327 GND.n7571 GND.n7570 36.7959
R16328 GND.n7570 GND.n7569 36.7959
R16329 GND.n7569 GND.n540 36.7959
R16330 GND.n7563 GND.n540 36.7959
R16331 GND.n5889 GND.n1756 36.428
R16332 GND.n5404 GND.n2557 36.428
R16333 GND.n1747 GND.n1746 35.8793
R16334 GND.n5870 GND.n1801 35.8793
R16335 GND.n3118 GND.n3117 35.8793
R16336 GND.n3183 GND.n3106 35.8793
R16337 GND.n5350 GND.n5349 35.8793
R16338 GND.n4828 GND.n4827 35.8793
R16339 GND.n302 GND.n257 35.8793
R16340 GND.n329 GND.n328 35.8793
R16341 GND.n229 GND.n228 35.8793
R16342 GND.n5114 GND.n5113 35.8793
R16343 GND.n2931 GND.n2900 35.8793
R16344 GND.n2409 GND.n2408 35.8793
R16345 GND.n4200 GND.n4199 35.8793
R16346 GND.n3521 GND.n3520 35.8793
R16347 GND.n3511 GND.n3510 35.8793
R16348 GND.n3617 GND.n3616 35.8793
R16349 GND.n3651 GND.n3650 35.8793
R16350 GND.n1666 GND.n1665 35.8793
R16351 GND.n2509 GND.n2503 34.4981
R16352 GND.n1950 GND.n1948 34.4981
R16353 GND.n1877 GND.n1876 32.1338
R16354 GND.n1866 GND.n1865 32.1338
R16355 GND.n2474 GND.n2473 32.1338
R16356 GND.n2492 GND.n2468 32.1338
R16357 GND.n6005 GND.n6004 32.0125
R16358 GND.n7731 GND.n379 32.0125
R16359 GND.n5852 GND.n5851 30.5925
R16360 GND.n5409 GND.n5408 30.5925
R16361 GND.n5852 GND.n1821 30.5518
R16362 GND.n5408 GND.n2553 30.5518
R16363 GND.n5847 GND.n1827 29.0689
R16364 GND.t79 GND.n1847 28.701
R16365 GND.n5804 GND.n1883 25.0214
R16366 GND.n1957 GND.n1894 25.0214
R16367 GND.t153 GND.n1903 25.0214
R16368 GND.n5470 GND.n2420 25.0214
R16369 GND.n5464 GND.n2428 25.0214
R16370 GND.n4811 GND.t144 23.5496
R16371 GND.n5458 GND.t126 22.0778
R16372 GND.n3669 GND.n3668 20.606
R16373 GND.n3680 GND.n3475 20.606
R16374 GND.n3679 GND.n3477 20.606
R16375 GND.n3690 GND.n3468 20.606
R16376 GND.n3691 GND.n3456 20.606
R16377 GND.n3706 GND.n3458 20.606
R16378 GND.n3717 GND.n3445 20.606
R16379 GND.n3727 GND.n3438 20.606
R16380 GND.n3728 GND.n3427 20.606
R16381 GND.n3743 GND.n3429 20.606
R16382 GND.n3754 GND.n3417 20.606
R16383 GND.n3753 GND.n3419 20.606
R16384 GND.n3764 GND.n3409 20.606
R16385 GND.n3765 GND.n3397 20.606
R16386 GND.n3780 GND.n3400 20.606
R16387 GND.n3791 GND.n3387 20.606
R16388 GND.n3790 GND.n3389 20.606
R16389 GND.n3807 GND.n3380 20.606
R16390 GND.n3809 GND.n3367 20.606
R16391 GND.n3817 GND.n3369 20.606
R16392 GND.n3371 GND.n3361 20.606
R16393 GND.n3826 GND.n3358 20.606
R16394 GND.n3937 GND.n3337 20.606
R16395 GND.n3836 GND.n3345 20.606
R16396 GND.n3930 GND.n3347 20.606
R16397 GND.n3877 GND.n3869 20.606
R16398 GND.n3879 GND.n3865 20.606
R16399 GND.n3889 GND.n3888 20.606
R16400 GND.n3900 GND.n3863 20.606
R16401 GND.n3902 GND.n3857 20.606
R16402 GND.n3905 GND.n3860 20.606
R16403 GND.n3859 GND.n3853 20.606
R16404 GND.n3912 GND.n3321 20.606
R16405 GND.n3948 GND.n3947 20.606
R16406 GND.n3963 GND.n3312 20.606
R16407 GND.n3974 GND.n3301 20.606
R16408 GND.n3973 GND.n3303 20.606
R16409 GND.n3984 GND.n3294 20.606
R16410 GND.n3985 GND.n3282 20.606
R16411 GND.n4000 GND.n3284 20.606
R16412 GND.n4011 GND.n3271 20.606
R16413 GND.n4010 GND.n3274 20.606
R16414 GND.n4021 GND.n3264 20.606
R16415 GND.n4022 GND.n3253 20.606
R16416 GND.n4037 GND.n3255 20.606
R16417 GND.n4048 GND.n3243 20.606
R16418 GND.n4047 GND.n3245 20.606
R16419 GND.n4058 GND.n3235 20.606
R16420 GND.n4059 GND.n3223 20.606
R16421 GND.n4074 GND.n3226 20.606
R16422 GND.n4085 GND.n3213 20.606
R16423 GND.n4084 GND.n3215 20.606
R16424 GND.n4128 GND.n3206 20.606
R16425 GND.n4130 GND.n3196 20.606
R16426 GND.n4140 GND.n3198 20.606
R16427 GND.n4133 GND.n3190 20.606
R16428 GND.n4149 GND.n3186 20.606
R16429 GND.n4223 GND.n3187 20.606
R16430 GND.n1954 GND.t132 20.606
R16431 GND.n4909 GND.n4825 20.606
R16432 GND.n5332 GND.n2594 20.606
R16433 GND.n5325 GND.n2597 20.606
R16434 GND.n5324 GND.n2608 20.606
R16435 GND.n2618 GND.n2617 20.606
R16436 GND.n5318 GND.n5317 20.606
R16437 GND.n4935 GND.n2621 20.606
R16438 GND.n5311 GND.n2636 20.606
R16439 GND.n4943 GND.n2891 20.606
R16440 GND.n5305 GND.n2647 20.606
R16441 GND.n4950 GND.n2650 20.606
R16442 GND.n5299 GND.n2658 20.606
R16443 GND.n4958 GND.n2661 20.606
R16444 GND.n5293 GND.n2668 20.606
R16445 GND.n4965 GND.n2671 20.606
R16446 GND.n5287 GND.n2679 20.606
R16447 GND.n4973 GND.n2682 20.606
R16448 GND.n5281 GND.n2689 20.606
R16449 GND.n4980 GND.n2692 20.606
R16450 GND.n5275 GND.n2700 20.606
R16451 GND.n4988 GND.n2703 20.606
R16452 GND.n5269 GND.n2710 20.606
R16453 GND.n4995 GND.n2713 20.606
R16454 GND.n5263 GND.n2721 20.606
R16455 GND.n5013 GND.n2815 20.606
R16456 GND.n5257 GND.n2730 20.606
R16457 GND.n5253 GND.n2733 20.606
R16458 GND.n5252 GND.n2738 20.606
R16459 GND.n2747 GND.n2744 20.606
R16460 GND.n5245 GND.n5244 20.606
R16461 GND.n7824 GND.n28 20.606
R16462 GND.n5238 GND.n30 20.606
R16463 GND.n5237 GND.n2759 20.606
R16464 GND.n5040 GND.n5033 20.606
R16465 GND.n7817 GND.n47 20.606
R16466 GND.n5047 GND.n50 20.606
R16467 GND.n5055 GND.n61 20.606
R16468 GND.n7805 GND.n68 20.606
R16469 GND.n5061 GND.n71 20.606
R16470 GND.n7799 GND.n78 20.606
R16471 GND.n5069 GND.n81 20.606
R16472 GND.n7793 GND.n89 20.606
R16473 GND.n5075 GND.n92 20.606
R16474 GND.n7787 GND.n99 20.606
R16475 GND.n5083 GND.n102 20.606
R16476 GND.n7781 GND.n110 20.606
R16477 GND.n5089 GND.n113 20.606
R16478 GND.n7775 GND.n120 20.606
R16479 GND.n5098 GND.n123 20.606
R16480 GND.n7769 GND.n131 20.606
R16481 GND.n5179 GND.n134 20.606
R16482 GND.n5173 GND.n143 20.606
R16483 GND.n7757 GND.n151 20.606
R16484 GND.n5167 GND.n154 20.606
R16485 GND.n7751 GND.n161 20.606
R16486 GND.n5161 GND.n164 20.606
R16487 GND.n7745 GND.n172 20.606
R16488 GND.n7738 GND.n175 20.606
R16489 GND.n1860 GND.t154 19.8005
R16490 GND.n1860 GND.t89 19.8005
R16491 GND.n1858 GND.t133 19.8005
R16492 GND.n1858 GND.t68 19.8005
R16493 GND.n1857 GND.t112 19.8005
R16494 GND.n1857 GND.t61 19.8005
R16495 GND.n2487 GND.t109 19.8005
R16496 GND.n2487 GND.t127 19.8005
R16497 GND.n2485 GND.t86 19.8005
R16498 GND.n2485 GND.t118 19.8005
R16499 GND.n2484 GND.t77 19.8005
R16500 GND.n2484 GND.t145 19.8005
R16501 GND.n1852 GND.n1851 19.5087
R16502 GND.n1875 GND.n1852 19.5087
R16503 GND.n1873 GND.n1854 19.5087
R16504 GND.n1869 GND.n1854 19.5087
R16505 GND.n1867 GND.n1856 19.5087
R16506 GND.n2478 GND.n2477 19.5087
R16507 GND.n2478 GND.n2469 19.5087
R16508 GND.n2491 GND.n2483 19.5087
R16509 GND.n4220 GND.n4151 19.3944
R16510 GND.n4213 GND.n4151 19.3944
R16511 GND.n4213 GND.n4212 19.3944
R16512 GND.n4212 GND.n4162 19.3944
R16513 GND.n4205 GND.n4162 19.3944
R16514 GND.n4205 GND.n4204 19.3944
R16515 GND.n4204 GND.n4173 19.3944
R16516 GND.n4194 GND.n4173 19.3944
R16517 GND.n4194 GND.n4193 19.3944
R16518 GND.n3657 GND.n3655 19.3944
R16519 GND.n3658 GND.n3657 19.3944
R16520 GND.n3660 GND.n3658 19.3944
R16521 GND.n3660 GND.n3461 19.3944
R16522 GND.n3704 GND.n3461 19.3944
R16523 GND.n3704 GND.n3462 19.3944
R16524 GND.n3695 GND.n3462 19.3944
R16525 GND.n3697 GND.n3695 19.3944
R16526 GND.n3697 GND.n3432 19.3944
R16527 GND.n3741 GND.n3432 19.3944
R16528 GND.n3741 GND.n3433 19.3944
R16529 GND.n3732 GND.n3433 19.3944
R16530 GND.n3734 GND.n3732 19.3944
R16531 GND.n3734 GND.n3403 19.3944
R16532 GND.n3778 GND.n3403 19.3944
R16533 GND.n3778 GND.n3404 19.3944
R16534 GND.n3769 GND.n3404 19.3944
R16535 GND.n3771 GND.n3769 19.3944
R16536 GND.n3771 GND.n3373 19.3944
R16537 GND.n3815 GND.n3373 19.3944
R16538 GND.n3815 GND.n3374 19.3944
R16539 GND.n3374 GND.n3356 19.3944
R16540 GND.n3832 GND.n3356 19.3944
R16541 GND.n3833 GND.n3832 19.3944
R16542 GND.n3833 GND.n3350 19.3944
R16543 GND.n3928 GND.n3350 19.3944
R16544 GND.n3928 GND.n3351 19.3944
R16545 GND.n3842 GND.n3351 19.3944
R16546 GND.n3843 GND.n3842 19.3944
R16547 GND.n3844 GND.n3843 19.3944
R16548 GND.n3862 GND.n3844 19.3944
R16549 GND.n3862 GND.n3850 19.3944
R16550 GND.n3851 GND.n3850 19.3944
R16551 GND.n3914 GND.n3851 19.3944
R16552 GND.n3914 GND.n3315 19.3944
R16553 GND.n3961 GND.n3315 19.3944
R16554 GND.n3961 GND.n3316 19.3944
R16555 GND.n3952 GND.n3316 19.3944
R16556 GND.n3954 GND.n3952 19.3944
R16557 GND.n3954 GND.n3287 19.3944
R16558 GND.n3998 GND.n3287 19.3944
R16559 GND.n3998 GND.n3288 19.3944
R16560 GND.n3989 GND.n3288 19.3944
R16561 GND.n3991 GND.n3989 19.3944
R16562 GND.n3991 GND.n3258 19.3944
R16563 GND.n4035 GND.n3258 19.3944
R16564 GND.n4035 GND.n3259 19.3944
R16565 GND.n4026 GND.n3259 19.3944
R16566 GND.n4028 GND.n4026 19.3944
R16567 GND.n4028 GND.n3229 19.3944
R16568 GND.n4072 GND.n3229 19.3944
R16569 GND.n4072 GND.n3230 19.3944
R16570 GND.n4063 GND.n3230 19.3944
R16571 GND.n4065 GND.n4063 19.3944
R16572 GND.n4065 GND.n3200 19.3944
R16573 GND.n4138 GND.n3200 19.3944
R16574 GND.n4138 GND.n3201 19.3944
R16575 GND.n3201 GND.n3189 19.3944
R16576 GND.n3189 GND.n3101 19.3944
R16577 GND.n3666 GND.n3493 19.3944
R16578 GND.n3662 GND.n3493 19.3944
R16579 GND.n3662 GND.n3465 19.3944
R16580 GND.n3693 GND.n3465 19.3944
R16581 GND.n3702 GND.n3693 19.3944
R16582 GND.n3702 GND.n3701 19.3944
R16583 GND.n3701 GND.n3700 19.3944
R16584 GND.n3700 GND.n3436 19.3944
R16585 GND.n3730 GND.n3436 19.3944
R16586 GND.n3739 GND.n3730 19.3944
R16587 GND.n3739 GND.n3738 19.3944
R16588 GND.n3738 GND.n3737 19.3944
R16589 GND.n3737 GND.n3407 19.3944
R16590 GND.n3767 GND.n3407 19.3944
R16591 GND.n3776 GND.n3767 19.3944
R16592 GND.n3776 GND.n3775 19.3944
R16593 GND.n3775 GND.n3774 19.3944
R16594 GND.n3774 GND.n3378 19.3944
R16595 GND.n3811 GND.n3378 19.3944
R16596 GND.n3813 GND.n3811 19.3944
R16597 GND.n3813 GND.n3812 19.3944
R16598 GND.n3812 GND.n3360 19.3944
R16599 GND.n3360 GND.n3354 19.3944
R16600 GND.n3835 GND.n3354 19.3944
R16601 GND.n3838 GND.n3835 19.3944
R16602 GND.n3926 GND.n3838 19.3944
R16603 GND.n3926 GND.n3925 19.3944
R16604 GND.n3925 GND.n3924 19.3944
R16605 GND.n3924 GND.n3841 19.3944
R16606 GND.n3920 GND.n3841 19.3944
R16607 GND.n3920 GND.n3919 19.3944
R16608 GND.n3919 GND.n3918 19.3944
R16609 GND.n3918 GND.n3849 19.3944
R16610 GND.n3849 GND.n3319 19.3944
R16611 GND.n3950 GND.n3319 19.3944
R16612 GND.n3959 GND.n3950 19.3944
R16613 GND.n3959 GND.n3958 19.3944
R16614 GND.n3958 GND.n3957 19.3944
R16615 GND.n3957 GND.n3291 19.3944
R16616 GND.n3987 GND.n3291 19.3944
R16617 GND.n3996 GND.n3987 19.3944
R16618 GND.n3996 GND.n3995 19.3944
R16619 GND.n3995 GND.n3994 19.3944
R16620 GND.n3994 GND.n3262 19.3944
R16621 GND.n4024 GND.n3262 19.3944
R16622 GND.n4033 GND.n4024 19.3944
R16623 GND.n4033 GND.n4032 19.3944
R16624 GND.n4032 GND.n4031 19.3944
R16625 GND.n4031 GND.n3233 19.3944
R16626 GND.n4061 GND.n3233 19.3944
R16627 GND.n4070 GND.n4061 19.3944
R16628 GND.n4070 GND.n4069 19.3944
R16629 GND.n4069 GND.n4068 19.3944
R16630 GND.n4068 GND.n3204 19.3944
R16631 GND.n4132 GND.n3204 19.3944
R16632 GND.n4136 GND.n4132 19.3944
R16633 GND.n4136 GND.n4135 19.3944
R16634 GND.n4135 GND.n3102 19.3944
R16635 GND.n4225 GND.n3102 19.3944
R16636 GND.n5887 GND.n1784 19.3944
R16637 GND.n5883 GND.n1784 19.3944
R16638 GND.n5883 GND.n5882 19.3944
R16639 GND.n5882 GND.n5881 19.3944
R16640 GND.n5881 GND.n1791 19.3944
R16641 GND.n5877 GND.n1791 19.3944
R16642 GND.n5877 GND.n5876 19.3944
R16643 GND.n5876 GND.n5875 19.3944
R16644 GND.n5875 GND.n1797 19.3944
R16645 GND.n5871 GND.n1797 19.3944
R16646 GND.n5869 GND.n5868 19.3944
R16647 GND.n5868 GND.n1805 19.3944
R16648 GND.n5864 GND.n1805 19.3944
R16649 GND.n5864 GND.n5863 19.3944
R16650 GND.n5863 GND.n5862 19.3944
R16651 GND.n5862 GND.n1811 19.3944
R16652 GND.n5858 GND.n1811 19.3944
R16653 GND.n5858 GND.n5857 19.3944
R16654 GND.n5857 GND.n5856 19.3944
R16655 GND.n5856 GND.n1817 19.3944
R16656 GND.n3133 GND.n1819 19.3944
R16657 GND.n3134 GND.n3133 19.3944
R16658 GND.n3137 GND.n3134 19.3944
R16659 GND.n3137 GND.n3126 19.3944
R16660 GND.n3141 GND.n3126 19.3944
R16661 GND.n3142 GND.n3141 19.3944
R16662 GND.n3145 GND.n3142 19.3944
R16663 GND.n3145 GND.n3122 19.3944
R16664 GND.n3149 GND.n3122 19.3944
R16665 GND.n3150 GND.n3149 19.3944
R16666 GND.n3153 GND.n3150 19.3944
R16667 GND.n3158 GND.n3157 19.3944
R16668 GND.n3161 GND.n3158 19.3944
R16669 GND.n3161 GND.n3112 19.3944
R16670 GND.n3165 GND.n3112 19.3944
R16671 GND.n3166 GND.n3165 19.3944
R16672 GND.n3169 GND.n3166 19.3944
R16673 GND.n3169 GND.n3108 19.3944
R16674 GND.n3173 GND.n3108 19.3944
R16675 GND.n3174 GND.n3173 19.3944
R16676 GND.n3177 GND.n3174 19.3944
R16677 GND.n3177 GND.n3104 19.3944
R16678 GND.n7337 GND.n677 19.3944
R16679 GND.n7343 GND.n677 19.3944
R16680 GND.n7343 GND.n675 19.3944
R16681 GND.n7347 GND.n675 19.3944
R16682 GND.n7347 GND.n671 19.3944
R16683 GND.n7353 GND.n671 19.3944
R16684 GND.n7353 GND.n669 19.3944
R16685 GND.n7357 GND.n669 19.3944
R16686 GND.n7357 GND.n665 19.3944
R16687 GND.n7363 GND.n665 19.3944
R16688 GND.n7363 GND.n663 19.3944
R16689 GND.n7367 GND.n663 19.3944
R16690 GND.n7367 GND.n659 19.3944
R16691 GND.n7373 GND.n659 19.3944
R16692 GND.n7373 GND.n657 19.3944
R16693 GND.n7377 GND.n657 19.3944
R16694 GND.n7377 GND.n653 19.3944
R16695 GND.n7383 GND.n653 19.3944
R16696 GND.n7383 GND.n651 19.3944
R16697 GND.n7387 GND.n651 19.3944
R16698 GND.n7387 GND.n647 19.3944
R16699 GND.n7393 GND.n647 19.3944
R16700 GND.n7393 GND.n645 19.3944
R16701 GND.n7397 GND.n645 19.3944
R16702 GND.n7397 GND.n641 19.3944
R16703 GND.n7403 GND.n641 19.3944
R16704 GND.n7403 GND.n639 19.3944
R16705 GND.n7407 GND.n639 19.3944
R16706 GND.n7407 GND.n635 19.3944
R16707 GND.n7413 GND.n635 19.3944
R16708 GND.n7413 GND.n633 19.3944
R16709 GND.n7417 GND.n633 19.3944
R16710 GND.n7417 GND.n629 19.3944
R16711 GND.n7423 GND.n629 19.3944
R16712 GND.n7423 GND.n627 19.3944
R16713 GND.n7427 GND.n627 19.3944
R16714 GND.n7427 GND.n623 19.3944
R16715 GND.n7433 GND.n623 19.3944
R16716 GND.n7433 GND.n621 19.3944
R16717 GND.n7437 GND.n621 19.3944
R16718 GND.n7437 GND.n617 19.3944
R16719 GND.n7443 GND.n617 19.3944
R16720 GND.n7443 GND.n615 19.3944
R16721 GND.n7447 GND.n615 19.3944
R16722 GND.n7447 GND.n611 19.3944
R16723 GND.n7453 GND.n611 19.3944
R16724 GND.n7453 GND.n609 19.3944
R16725 GND.n7457 GND.n609 19.3944
R16726 GND.n7457 GND.n605 19.3944
R16727 GND.n7463 GND.n605 19.3944
R16728 GND.n7463 GND.n603 19.3944
R16729 GND.n7467 GND.n603 19.3944
R16730 GND.n7467 GND.n599 19.3944
R16731 GND.n7473 GND.n599 19.3944
R16732 GND.n7473 GND.n597 19.3944
R16733 GND.n7477 GND.n597 19.3944
R16734 GND.n7477 GND.n593 19.3944
R16735 GND.n7483 GND.n593 19.3944
R16736 GND.n7483 GND.n591 19.3944
R16737 GND.n7487 GND.n591 19.3944
R16738 GND.n7487 GND.n587 19.3944
R16739 GND.n7493 GND.n587 19.3944
R16740 GND.n7493 GND.n585 19.3944
R16741 GND.n7497 GND.n585 19.3944
R16742 GND.n7497 GND.n581 19.3944
R16743 GND.n7503 GND.n581 19.3944
R16744 GND.n7503 GND.n579 19.3944
R16745 GND.n7507 GND.n579 19.3944
R16746 GND.n7507 GND.n575 19.3944
R16747 GND.n7513 GND.n575 19.3944
R16748 GND.n7513 GND.n573 19.3944
R16749 GND.n7517 GND.n573 19.3944
R16750 GND.n7517 GND.n569 19.3944
R16751 GND.n7523 GND.n569 19.3944
R16752 GND.n7523 GND.n567 19.3944
R16753 GND.n7527 GND.n567 19.3944
R16754 GND.n7527 GND.n563 19.3944
R16755 GND.n7533 GND.n563 19.3944
R16756 GND.n7533 GND.n561 19.3944
R16757 GND.n7537 GND.n561 19.3944
R16758 GND.n7537 GND.n557 19.3944
R16759 GND.n7543 GND.n557 19.3944
R16760 GND.n7543 GND.n555 19.3944
R16761 GND.n7547 GND.n555 19.3944
R16762 GND.n7547 GND.n551 19.3944
R16763 GND.n7553 GND.n551 19.3944
R16764 GND.n7553 GND.n549 19.3944
R16765 GND.n7559 GND.n549 19.3944
R16766 GND.n7559 GND.n7558 19.3944
R16767 GND.n6356 GND.n1264 19.3944
R16768 GND.n6362 GND.n1264 19.3944
R16769 GND.n6362 GND.n1262 19.3944
R16770 GND.n6366 GND.n1262 19.3944
R16771 GND.n6366 GND.n1258 19.3944
R16772 GND.n6372 GND.n1258 19.3944
R16773 GND.n6372 GND.n1256 19.3944
R16774 GND.n6376 GND.n1256 19.3944
R16775 GND.n6376 GND.n1252 19.3944
R16776 GND.n6382 GND.n1252 19.3944
R16777 GND.n6382 GND.n1250 19.3944
R16778 GND.n6386 GND.n1250 19.3944
R16779 GND.n6386 GND.n1246 19.3944
R16780 GND.n6392 GND.n1246 19.3944
R16781 GND.n6392 GND.n1244 19.3944
R16782 GND.n6396 GND.n1244 19.3944
R16783 GND.n6396 GND.n1240 19.3944
R16784 GND.n6402 GND.n1240 19.3944
R16785 GND.n6402 GND.n1238 19.3944
R16786 GND.n6406 GND.n1238 19.3944
R16787 GND.n6406 GND.n1234 19.3944
R16788 GND.n6412 GND.n1234 19.3944
R16789 GND.n6412 GND.n1232 19.3944
R16790 GND.n6416 GND.n1232 19.3944
R16791 GND.n6416 GND.n1228 19.3944
R16792 GND.n6422 GND.n1228 19.3944
R16793 GND.n6422 GND.n1226 19.3944
R16794 GND.n6426 GND.n1226 19.3944
R16795 GND.n6426 GND.n1222 19.3944
R16796 GND.n6432 GND.n1222 19.3944
R16797 GND.n6432 GND.n1220 19.3944
R16798 GND.n6436 GND.n1220 19.3944
R16799 GND.n6436 GND.n1216 19.3944
R16800 GND.n6442 GND.n1216 19.3944
R16801 GND.n6442 GND.n1214 19.3944
R16802 GND.n6446 GND.n1214 19.3944
R16803 GND.n6446 GND.n1210 19.3944
R16804 GND.n6452 GND.n1210 19.3944
R16805 GND.n6452 GND.n1208 19.3944
R16806 GND.n6456 GND.n1208 19.3944
R16807 GND.n6456 GND.n1204 19.3944
R16808 GND.n6462 GND.n1204 19.3944
R16809 GND.n6462 GND.n1202 19.3944
R16810 GND.n6466 GND.n1202 19.3944
R16811 GND.n6466 GND.n1198 19.3944
R16812 GND.n6472 GND.n1198 19.3944
R16813 GND.n6472 GND.n1196 19.3944
R16814 GND.n6476 GND.n1196 19.3944
R16815 GND.n6476 GND.n1192 19.3944
R16816 GND.n6482 GND.n1192 19.3944
R16817 GND.n6482 GND.n1190 19.3944
R16818 GND.n6486 GND.n1190 19.3944
R16819 GND.n6486 GND.n1186 19.3944
R16820 GND.n6492 GND.n1186 19.3944
R16821 GND.n6492 GND.n1184 19.3944
R16822 GND.n6496 GND.n1184 19.3944
R16823 GND.n6496 GND.n1180 19.3944
R16824 GND.n6502 GND.n1180 19.3944
R16825 GND.n6502 GND.n1178 19.3944
R16826 GND.n6506 GND.n1178 19.3944
R16827 GND.n6506 GND.n1174 19.3944
R16828 GND.n6512 GND.n1174 19.3944
R16829 GND.n6512 GND.n1172 19.3944
R16830 GND.n6516 GND.n1172 19.3944
R16831 GND.n6516 GND.n1168 19.3944
R16832 GND.n6522 GND.n1168 19.3944
R16833 GND.n6522 GND.n1166 19.3944
R16834 GND.n6526 GND.n1166 19.3944
R16835 GND.n6526 GND.n1162 19.3944
R16836 GND.n6532 GND.n1162 19.3944
R16837 GND.n6532 GND.n1160 19.3944
R16838 GND.n6536 GND.n1160 19.3944
R16839 GND.n6536 GND.n1156 19.3944
R16840 GND.n6542 GND.n1156 19.3944
R16841 GND.n6542 GND.n1154 19.3944
R16842 GND.n6546 GND.n1154 19.3944
R16843 GND.n6546 GND.n1150 19.3944
R16844 GND.n6552 GND.n1150 19.3944
R16845 GND.n6552 GND.n1148 19.3944
R16846 GND.n6556 GND.n1148 19.3944
R16847 GND.n6556 GND.n1144 19.3944
R16848 GND.n6562 GND.n1144 19.3944
R16849 GND.n6562 GND.n1142 19.3944
R16850 GND.n6566 GND.n1142 19.3944
R16851 GND.n6566 GND.n1138 19.3944
R16852 GND.n6572 GND.n1138 19.3944
R16853 GND.n6572 GND.n1136 19.3944
R16854 GND.n6576 GND.n1136 19.3944
R16855 GND.n6576 GND.n1132 19.3944
R16856 GND.n6582 GND.n1132 19.3944
R16857 GND.n6582 GND.n1130 19.3944
R16858 GND.n6586 GND.n1130 19.3944
R16859 GND.n6586 GND.n1126 19.3944
R16860 GND.n6592 GND.n1126 19.3944
R16861 GND.n6592 GND.n1124 19.3944
R16862 GND.n6596 GND.n1124 19.3944
R16863 GND.n6596 GND.n1120 19.3944
R16864 GND.n6602 GND.n1120 19.3944
R16865 GND.n6602 GND.n1118 19.3944
R16866 GND.n6606 GND.n1118 19.3944
R16867 GND.n6606 GND.n1114 19.3944
R16868 GND.n6612 GND.n1114 19.3944
R16869 GND.n6612 GND.n1112 19.3944
R16870 GND.n6616 GND.n1112 19.3944
R16871 GND.n6616 GND.n1108 19.3944
R16872 GND.n6622 GND.n1108 19.3944
R16873 GND.n6622 GND.n1106 19.3944
R16874 GND.n6626 GND.n1106 19.3944
R16875 GND.n6626 GND.n1102 19.3944
R16876 GND.n6632 GND.n1102 19.3944
R16877 GND.n6632 GND.n1100 19.3944
R16878 GND.n6636 GND.n1100 19.3944
R16879 GND.n6636 GND.n1096 19.3944
R16880 GND.n6642 GND.n1096 19.3944
R16881 GND.n6642 GND.n1094 19.3944
R16882 GND.n6646 GND.n1094 19.3944
R16883 GND.n6646 GND.n1090 19.3944
R16884 GND.n6652 GND.n1090 19.3944
R16885 GND.n6652 GND.n1088 19.3944
R16886 GND.n6656 GND.n1088 19.3944
R16887 GND.n6656 GND.n1084 19.3944
R16888 GND.n6662 GND.n1084 19.3944
R16889 GND.n6662 GND.n1082 19.3944
R16890 GND.n6666 GND.n1082 19.3944
R16891 GND.n6666 GND.n1078 19.3944
R16892 GND.n6672 GND.n1078 19.3944
R16893 GND.n6672 GND.n1076 19.3944
R16894 GND.n6676 GND.n1076 19.3944
R16895 GND.n6676 GND.n1072 19.3944
R16896 GND.n6682 GND.n1072 19.3944
R16897 GND.n6682 GND.n1070 19.3944
R16898 GND.n6686 GND.n1070 19.3944
R16899 GND.n6686 GND.n1066 19.3944
R16900 GND.n6692 GND.n1066 19.3944
R16901 GND.n6692 GND.n1064 19.3944
R16902 GND.n6696 GND.n1064 19.3944
R16903 GND.n6696 GND.n1060 19.3944
R16904 GND.n6702 GND.n1060 19.3944
R16905 GND.n6702 GND.n1058 19.3944
R16906 GND.n6706 GND.n1058 19.3944
R16907 GND.n6706 GND.n1054 19.3944
R16908 GND.n6712 GND.n1054 19.3944
R16909 GND.n6712 GND.n1052 19.3944
R16910 GND.n6716 GND.n1052 19.3944
R16911 GND.n6716 GND.n1048 19.3944
R16912 GND.n6722 GND.n1048 19.3944
R16913 GND.n6722 GND.n1046 19.3944
R16914 GND.n6726 GND.n1046 19.3944
R16915 GND.n6726 GND.n1042 19.3944
R16916 GND.n6732 GND.n1042 19.3944
R16917 GND.n6732 GND.n1040 19.3944
R16918 GND.n6736 GND.n1040 19.3944
R16919 GND.n6736 GND.n1036 19.3944
R16920 GND.n6742 GND.n1036 19.3944
R16921 GND.n6742 GND.n1034 19.3944
R16922 GND.n6746 GND.n1034 19.3944
R16923 GND.n6746 GND.n1030 19.3944
R16924 GND.n6752 GND.n1030 19.3944
R16925 GND.n6752 GND.n1028 19.3944
R16926 GND.n6756 GND.n1028 19.3944
R16927 GND.n6756 GND.n1024 19.3944
R16928 GND.n6762 GND.n1024 19.3944
R16929 GND.n6762 GND.n1022 19.3944
R16930 GND.n6766 GND.n1022 19.3944
R16931 GND.n6766 GND.n1018 19.3944
R16932 GND.n6772 GND.n1018 19.3944
R16933 GND.n6772 GND.n1016 19.3944
R16934 GND.n6776 GND.n1016 19.3944
R16935 GND.n6776 GND.n1012 19.3944
R16936 GND.n6782 GND.n1012 19.3944
R16937 GND.n6782 GND.n1010 19.3944
R16938 GND.n6786 GND.n1010 19.3944
R16939 GND.n6786 GND.n1006 19.3944
R16940 GND.n6792 GND.n1006 19.3944
R16941 GND.n6792 GND.n1004 19.3944
R16942 GND.n6796 GND.n1004 19.3944
R16943 GND.n6796 GND.n1000 19.3944
R16944 GND.n6802 GND.n1000 19.3944
R16945 GND.n6802 GND.n998 19.3944
R16946 GND.n6806 GND.n998 19.3944
R16947 GND.n6806 GND.n994 19.3944
R16948 GND.n6812 GND.n994 19.3944
R16949 GND.n6812 GND.n992 19.3944
R16950 GND.n6816 GND.n992 19.3944
R16951 GND.n6816 GND.n988 19.3944
R16952 GND.n6822 GND.n988 19.3944
R16953 GND.n6822 GND.n986 19.3944
R16954 GND.n6826 GND.n986 19.3944
R16955 GND.n6826 GND.n982 19.3944
R16956 GND.n6832 GND.n982 19.3944
R16957 GND.n6832 GND.n980 19.3944
R16958 GND.n6836 GND.n980 19.3944
R16959 GND.n6836 GND.n976 19.3944
R16960 GND.n6842 GND.n976 19.3944
R16961 GND.n6842 GND.n974 19.3944
R16962 GND.n6846 GND.n974 19.3944
R16963 GND.n6846 GND.n970 19.3944
R16964 GND.n6852 GND.n970 19.3944
R16965 GND.n6852 GND.n968 19.3944
R16966 GND.n6856 GND.n968 19.3944
R16967 GND.n6856 GND.n964 19.3944
R16968 GND.n6862 GND.n964 19.3944
R16969 GND.n6862 GND.n962 19.3944
R16970 GND.n6866 GND.n962 19.3944
R16971 GND.n6866 GND.n958 19.3944
R16972 GND.n6872 GND.n958 19.3944
R16973 GND.n6872 GND.n956 19.3944
R16974 GND.n6876 GND.n956 19.3944
R16975 GND.n6876 GND.n952 19.3944
R16976 GND.n6882 GND.n952 19.3944
R16977 GND.n6882 GND.n950 19.3944
R16978 GND.n6886 GND.n950 19.3944
R16979 GND.n6886 GND.n946 19.3944
R16980 GND.n6892 GND.n946 19.3944
R16981 GND.n6892 GND.n944 19.3944
R16982 GND.n6896 GND.n944 19.3944
R16983 GND.n6896 GND.n940 19.3944
R16984 GND.n6902 GND.n940 19.3944
R16985 GND.n6902 GND.n938 19.3944
R16986 GND.n6906 GND.n938 19.3944
R16987 GND.n6906 GND.n934 19.3944
R16988 GND.n6912 GND.n934 19.3944
R16989 GND.n6912 GND.n932 19.3944
R16990 GND.n6916 GND.n932 19.3944
R16991 GND.n6916 GND.n928 19.3944
R16992 GND.n6922 GND.n928 19.3944
R16993 GND.n6922 GND.n926 19.3944
R16994 GND.n6926 GND.n926 19.3944
R16995 GND.n6926 GND.n922 19.3944
R16996 GND.n6932 GND.n922 19.3944
R16997 GND.n6932 GND.n920 19.3944
R16998 GND.n6936 GND.n920 19.3944
R16999 GND.n6936 GND.n916 19.3944
R17000 GND.n6942 GND.n916 19.3944
R17001 GND.n6942 GND.n914 19.3944
R17002 GND.n6946 GND.n914 19.3944
R17003 GND.n6946 GND.n910 19.3944
R17004 GND.n6952 GND.n910 19.3944
R17005 GND.n6952 GND.n908 19.3944
R17006 GND.n6956 GND.n908 19.3944
R17007 GND.n6956 GND.n904 19.3944
R17008 GND.n6962 GND.n904 19.3944
R17009 GND.n6962 GND.n902 19.3944
R17010 GND.n6966 GND.n902 19.3944
R17011 GND.n6966 GND.n898 19.3944
R17012 GND.n6972 GND.n898 19.3944
R17013 GND.n6972 GND.n896 19.3944
R17014 GND.n6976 GND.n896 19.3944
R17015 GND.n6976 GND.n892 19.3944
R17016 GND.n6982 GND.n892 19.3944
R17017 GND.n6982 GND.n890 19.3944
R17018 GND.n6986 GND.n890 19.3944
R17019 GND.n6986 GND.n886 19.3944
R17020 GND.n6992 GND.n886 19.3944
R17021 GND.n6992 GND.n884 19.3944
R17022 GND.n6996 GND.n884 19.3944
R17023 GND.n6996 GND.n880 19.3944
R17024 GND.n7002 GND.n880 19.3944
R17025 GND.n7002 GND.n878 19.3944
R17026 GND.n7006 GND.n878 19.3944
R17027 GND.n7006 GND.n874 19.3944
R17028 GND.n7012 GND.n874 19.3944
R17029 GND.n7012 GND.n872 19.3944
R17030 GND.n7016 GND.n872 19.3944
R17031 GND.n7016 GND.n868 19.3944
R17032 GND.n7022 GND.n868 19.3944
R17033 GND.n7022 GND.n866 19.3944
R17034 GND.n7026 GND.n866 19.3944
R17035 GND.n7026 GND.n862 19.3944
R17036 GND.n7032 GND.n862 19.3944
R17037 GND.n7032 GND.n860 19.3944
R17038 GND.n7036 GND.n860 19.3944
R17039 GND.n7036 GND.n856 19.3944
R17040 GND.n7042 GND.n856 19.3944
R17041 GND.n7042 GND.n854 19.3944
R17042 GND.n7046 GND.n854 19.3944
R17043 GND.n7046 GND.n850 19.3944
R17044 GND.n7052 GND.n850 19.3944
R17045 GND.n7052 GND.n848 19.3944
R17046 GND.n7056 GND.n848 19.3944
R17047 GND.n7056 GND.n844 19.3944
R17048 GND.n7062 GND.n844 19.3944
R17049 GND.n7062 GND.n842 19.3944
R17050 GND.n7066 GND.n842 19.3944
R17051 GND.n7066 GND.n838 19.3944
R17052 GND.n7072 GND.n838 19.3944
R17053 GND.n7072 GND.n836 19.3944
R17054 GND.n7076 GND.n836 19.3944
R17055 GND.n7076 GND.n832 19.3944
R17056 GND.n7082 GND.n832 19.3944
R17057 GND.n7082 GND.n830 19.3944
R17058 GND.n7086 GND.n830 19.3944
R17059 GND.n7086 GND.n826 19.3944
R17060 GND.n7092 GND.n826 19.3944
R17061 GND.n7092 GND.n824 19.3944
R17062 GND.n7096 GND.n824 19.3944
R17063 GND.n7096 GND.n820 19.3944
R17064 GND.n7102 GND.n820 19.3944
R17065 GND.n7102 GND.n818 19.3944
R17066 GND.n7106 GND.n818 19.3944
R17067 GND.n7106 GND.n814 19.3944
R17068 GND.n7112 GND.n814 19.3944
R17069 GND.n7112 GND.n812 19.3944
R17070 GND.n7116 GND.n812 19.3944
R17071 GND.n7116 GND.n808 19.3944
R17072 GND.n7122 GND.n808 19.3944
R17073 GND.n7122 GND.n806 19.3944
R17074 GND.n7126 GND.n806 19.3944
R17075 GND.n7126 GND.n802 19.3944
R17076 GND.n7132 GND.n802 19.3944
R17077 GND.n7132 GND.n800 19.3944
R17078 GND.n7136 GND.n800 19.3944
R17079 GND.n7136 GND.n796 19.3944
R17080 GND.n7142 GND.n796 19.3944
R17081 GND.n7142 GND.n794 19.3944
R17082 GND.n7146 GND.n794 19.3944
R17083 GND.n7146 GND.n790 19.3944
R17084 GND.n7152 GND.n790 19.3944
R17085 GND.n7152 GND.n788 19.3944
R17086 GND.n7156 GND.n788 19.3944
R17087 GND.n7156 GND.n784 19.3944
R17088 GND.n7162 GND.n784 19.3944
R17089 GND.n7162 GND.n782 19.3944
R17090 GND.n7166 GND.n782 19.3944
R17091 GND.n7166 GND.n778 19.3944
R17092 GND.n7172 GND.n778 19.3944
R17093 GND.n7172 GND.n776 19.3944
R17094 GND.n7176 GND.n776 19.3944
R17095 GND.n7176 GND.n772 19.3944
R17096 GND.n7182 GND.n772 19.3944
R17097 GND.n7182 GND.n770 19.3944
R17098 GND.n7186 GND.n770 19.3944
R17099 GND.n7186 GND.n766 19.3944
R17100 GND.n7192 GND.n766 19.3944
R17101 GND.n7192 GND.n764 19.3944
R17102 GND.n7196 GND.n764 19.3944
R17103 GND.n7196 GND.n760 19.3944
R17104 GND.n7202 GND.n760 19.3944
R17105 GND.n7202 GND.n758 19.3944
R17106 GND.n7206 GND.n758 19.3944
R17107 GND.n7206 GND.n754 19.3944
R17108 GND.n7212 GND.n754 19.3944
R17109 GND.n7212 GND.n752 19.3944
R17110 GND.n7216 GND.n752 19.3944
R17111 GND.n7216 GND.n748 19.3944
R17112 GND.n7222 GND.n748 19.3944
R17113 GND.n7222 GND.n746 19.3944
R17114 GND.n7226 GND.n746 19.3944
R17115 GND.n7226 GND.n742 19.3944
R17116 GND.n7232 GND.n742 19.3944
R17117 GND.n7232 GND.n740 19.3944
R17118 GND.n7236 GND.n740 19.3944
R17119 GND.n7236 GND.n736 19.3944
R17120 GND.n7242 GND.n736 19.3944
R17121 GND.n7242 GND.n734 19.3944
R17122 GND.n7246 GND.n734 19.3944
R17123 GND.n7246 GND.n730 19.3944
R17124 GND.n7252 GND.n730 19.3944
R17125 GND.n7252 GND.n728 19.3944
R17126 GND.n7256 GND.n728 19.3944
R17127 GND.n7256 GND.n724 19.3944
R17128 GND.n7262 GND.n724 19.3944
R17129 GND.n7262 GND.n722 19.3944
R17130 GND.n7266 GND.n722 19.3944
R17131 GND.n7266 GND.n718 19.3944
R17132 GND.n7272 GND.n718 19.3944
R17133 GND.n7272 GND.n716 19.3944
R17134 GND.n7276 GND.n716 19.3944
R17135 GND.n7276 GND.n712 19.3944
R17136 GND.n7282 GND.n712 19.3944
R17137 GND.n7282 GND.n710 19.3944
R17138 GND.n7286 GND.n710 19.3944
R17139 GND.n7286 GND.n706 19.3944
R17140 GND.n7292 GND.n706 19.3944
R17141 GND.n7292 GND.n704 19.3944
R17142 GND.n7296 GND.n704 19.3944
R17143 GND.n7296 GND.n700 19.3944
R17144 GND.n7302 GND.n700 19.3944
R17145 GND.n7302 GND.n698 19.3944
R17146 GND.n7306 GND.n698 19.3944
R17147 GND.n7306 GND.n694 19.3944
R17148 GND.n7312 GND.n694 19.3944
R17149 GND.n7312 GND.n692 19.3944
R17150 GND.n7316 GND.n692 19.3944
R17151 GND.n7316 GND.n688 19.3944
R17152 GND.n7322 GND.n688 19.3944
R17153 GND.n7322 GND.n686 19.3944
R17154 GND.n7327 GND.n686 19.3944
R17155 GND.n7327 GND.n682 19.3944
R17156 GND.n7333 GND.n682 19.3944
R17157 GND.n7334 GND.n7333 19.3944
R17158 GND.n5401 GND.n5400 19.3944
R17159 GND.n5400 GND.n5399 19.3944
R17160 GND.n5399 GND.n5398 19.3944
R17161 GND.n5398 GND.n5396 19.3944
R17162 GND.n5396 GND.n5393 19.3944
R17163 GND.n5393 GND.n5392 19.3944
R17164 GND.n5392 GND.n5389 19.3944
R17165 GND.n5389 GND.n5388 19.3944
R17166 GND.n5388 GND.n5385 19.3944
R17167 GND.n5385 GND.n5384 19.3944
R17168 GND.n5381 GND.n5380 19.3944
R17169 GND.n5380 GND.n5377 19.3944
R17170 GND.n5377 GND.n5376 19.3944
R17171 GND.n5376 GND.n5373 19.3944
R17172 GND.n5373 GND.n5372 19.3944
R17173 GND.n5372 GND.n5369 19.3944
R17174 GND.n5369 GND.n5368 19.3944
R17175 GND.n5368 GND.n5365 19.3944
R17176 GND.n5365 GND.n5364 19.3944
R17177 GND.n5364 GND.n2549 19.3944
R17178 GND.n5407 GND.n2555 19.3944
R17179 GND.n4842 GND.n2555 19.3944
R17180 GND.n4845 GND.n4842 19.3944
R17181 GND.n4848 GND.n4845 19.3944
R17182 GND.n4848 GND.n4838 19.3944
R17183 GND.n4852 GND.n4838 19.3944
R17184 GND.n4855 GND.n4852 19.3944
R17185 GND.n4858 GND.n4855 19.3944
R17186 GND.n4858 GND.n4836 19.3944
R17187 GND.n4862 GND.n4836 19.3944
R17188 GND.n4865 GND.n4862 19.3944
R17189 GND.n4874 GND.n4834 19.3944
R17190 GND.n4877 GND.n4874 19.3944
R17191 GND.n4880 GND.n4877 19.3944
R17192 GND.n4880 GND.n4832 19.3944
R17193 GND.n4884 GND.n4832 19.3944
R17194 GND.n4887 GND.n4884 19.3944
R17195 GND.n4890 GND.n4887 19.3944
R17196 GND.n4890 GND.n4830 19.3944
R17197 GND.n4894 GND.n4830 19.3944
R17198 GND.n4897 GND.n4894 19.3944
R17199 GND.n4900 GND.n4897 19.3944
R17200 GND.n5328 GND.n2604 19.3944
R17201 GND.n5328 GND.n5327 19.3944
R17202 GND.n5327 GND.n2605 19.3944
R17203 GND.n4923 GND.n2605 19.3944
R17204 GND.n4923 GND.n4921 19.3944
R17205 GND.n4933 GND.n4921 19.3944
R17206 GND.n4933 GND.n2831 19.3944
R17207 GND.n4945 GND.n2831 19.3944
R17208 GND.n4946 GND.n4945 19.3944
R17209 GND.n4948 GND.n4946 19.3944
R17210 GND.n4948 GND.n2827 19.3944
R17211 GND.n4960 GND.n2827 19.3944
R17212 GND.n4961 GND.n4960 19.3944
R17213 GND.n4963 GND.n4961 19.3944
R17214 GND.n4963 GND.n2823 19.3944
R17215 GND.n4975 GND.n2823 19.3944
R17216 GND.n4976 GND.n4975 19.3944
R17217 GND.n4978 GND.n4976 19.3944
R17218 GND.n4978 GND.n2819 19.3944
R17219 GND.n4990 GND.n2819 19.3944
R17220 GND.n4991 GND.n4990 19.3944
R17221 GND.n4993 GND.n4991 19.3944
R17222 GND.n4993 GND.n2814 19.3944
R17223 GND.n5015 GND.n2814 19.3944
R17224 GND.n5016 GND.n5015 19.3944
R17225 GND.n5017 GND.n5016 19.3944
R17226 GND.n5017 GND.n2813 19.3944
R17227 GND.n5025 GND.n2813 19.3944
R17228 GND.n5026 GND.n5025 19.3944
R17229 GND.n5027 GND.n5026 19.3944
R17230 GND.n5028 GND.n5027 19.3944
R17231 GND.n5029 GND.n5028 19.3944
R17232 GND.n5042 GND.n5029 19.3944
R17233 GND.n5043 GND.n5042 19.3944
R17234 GND.n5044 GND.n5043 19.3944
R17235 GND.n5044 GND.n2808 19.3944
R17236 GND.n5057 GND.n2808 19.3944
R17237 GND.n5058 GND.n5057 19.3944
R17238 GND.n5059 GND.n5058 19.3944
R17239 GND.n5059 GND.n2803 19.3944
R17240 GND.n5071 GND.n2803 19.3944
R17241 GND.n5072 GND.n5071 19.3944
R17242 GND.n5073 GND.n5072 19.3944
R17243 GND.n5073 GND.n2798 19.3944
R17244 GND.n5085 GND.n2798 19.3944
R17245 GND.n5086 GND.n5085 19.3944
R17246 GND.n5087 GND.n5086 19.3944
R17247 GND.n5087 GND.n2793 19.3944
R17248 GND.n5100 GND.n2793 19.3944
R17249 GND.n5101 GND.n5100 19.3944
R17250 GND.n5102 GND.n5101 19.3944
R17251 GND.n5103 GND.n5102 19.3944
R17252 GND.n5171 GND.n5103 19.3944
R17253 GND.n5171 GND.n5170 19.3944
R17254 GND.n5170 GND.n5169 19.3944
R17255 GND.n5169 GND.n5105 19.3944
R17256 GND.n5159 GND.n5105 19.3944
R17257 GND.n5159 GND.n179 19.3944
R17258 GND.n7740 GND.n179 19.3944
R17259 GND.n5330 GND.n2600 19.3944
R17260 GND.n5330 GND.n2601 19.3944
R17261 GND.n4926 GND.n2601 19.3944
R17262 GND.n4929 GND.n4926 19.3944
R17263 GND.n4930 GND.n4929 19.3944
R17264 GND.n4930 GND.n2641 19.3944
R17265 GND.n5309 GND.n2641 19.3944
R17266 GND.n5309 GND.n5308 19.3944
R17267 GND.n5308 GND.n5307 19.3944
R17268 GND.n5307 GND.n2645 19.3944
R17269 GND.n5297 GND.n2645 19.3944
R17270 GND.n5297 GND.n5296 19.3944
R17271 GND.n5296 GND.n5295 19.3944
R17272 GND.n5295 GND.n2666 19.3944
R17273 GND.n5285 GND.n2666 19.3944
R17274 GND.n5285 GND.n5284 19.3944
R17275 GND.n5284 GND.n5283 19.3944
R17276 GND.n5283 GND.n2687 19.3944
R17277 GND.n5273 GND.n2687 19.3944
R17278 GND.n5273 GND.n5272 19.3944
R17279 GND.n5272 GND.n5271 19.3944
R17280 GND.n5271 GND.n2708 19.3944
R17281 GND.n5261 GND.n2708 19.3944
R17282 GND.n5261 GND.n5260 19.3944
R17283 GND.n5260 GND.n5259 19.3944
R17284 GND.n5259 GND.n2728 19.3944
R17285 GND.n5020 GND.n2728 19.3944
R17286 GND.n5020 GND.n2750 19.3944
R17287 GND.n5242 GND.n2750 19.3944
R17288 GND.n5242 GND.n5241 19.3944
R17289 GND.n5241 GND.n5240 19.3944
R17290 GND.n5240 GND.n2754 19.3944
R17291 GND.n2754 GND.n53 19.3944
R17292 GND.n7815 GND.n53 19.3944
R17293 GND.n7815 GND.n7814 19.3944
R17294 GND.n7814 GND.n7813 19.3944
R17295 GND.n7813 GND.n57 19.3944
R17296 GND.n7803 GND.n57 19.3944
R17297 GND.n7803 GND.n7802 19.3944
R17298 GND.n7802 GND.n7801 19.3944
R17299 GND.n7801 GND.n76 19.3944
R17300 GND.n7791 GND.n76 19.3944
R17301 GND.n7791 GND.n7790 19.3944
R17302 GND.n7790 GND.n7789 19.3944
R17303 GND.n7789 GND.n97 19.3944
R17304 GND.n7779 GND.n97 19.3944
R17305 GND.n7779 GND.n7778 19.3944
R17306 GND.n7778 GND.n7777 19.3944
R17307 GND.n7777 GND.n118 19.3944
R17308 GND.n7767 GND.n118 19.3944
R17309 GND.n7767 GND.n7766 19.3944
R17310 GND.n7766 GND.n7765 19.3944
R17311 GND.n7765 GND.n139 19.3944
R17312 GND.n7755 GND.n139 19.3944
R17313 GND.n7755 GND.n7754 19.3944
R17314 GND.n7754 GND.n7753 19.3944
R17315 GND.n7753 GND.n159 19.3944
R17316 GND.n7743 GND.n159 19.3944
R17317 GND.n7743 GND.n7742 19.3944
R17318 GND.n298 GND.n255 19.3944
R17319 GND.n298 GND.n295 19.3944
R17320 GND.n295 GND.n294 19.3944
R17321 GND.n294 GND.n291 19.3944
R17322 GND.n291 GND.n290 19.3944
R17323 GND.n290 GND.n287 19.3944
R17324 GND.n287 GND.n286 19.3944
R17325 GND.n286 GND.n283 19.3944
R17326 GND.n283 GND.n282 19.3944
R17327 GND.n282 GND.n279 19.3944
R17328 GND.n279 GND.n278 19.3944
R17329 GND.n326 GND.n323 19.3944
R17330 GND.n323 GND.n322 19.3944
R17331 GND.n322 GND.n319 19.3944
R17332 GND.n319 GND.n318 19.3944
R17333 GND.n318 GND.n315 19.3944
R17334 GND.n315 GND.n314 19.3944
R17335 GND.n314 GND.n311 19.3944
R17336 GND.n311 GND.n310 19.3944
R17337 GND.n310 GND.n307 19.3944
R17338 GND.n307 GND.n306 19.3944
R17339 GND.n306 GND.n303 19.3944
R17340 GND.n354 GND.n353 19.3944
R17341 GND.n353 GND.n350 19.3944
R17342 GND.n350 GND.n349 19.3944
R17343 GND.n349 GND.n346 19.3944
R17344 GND.n346 GND.n345 19.3944
R17345 GND.n345 GND.n342 19.3944
R17346 GND.n342 GND.n341 19.3944
R17347 GND.n341 GND.n338 19.3944
R17348 GND.n338 GND.n337 19.3944
R17349 GND.n337 GND.n334 19.3944
R17350 GND.n334 GND.n333 19.3944
R17351 GND.n333 GND.n330 19.3944
R17352 GND.n377 GND.n376 19.3944
R17353 GND.n376 GND.n219 19.3944
R17354 GND.n372 GND.n219 19.3944
R17355 GND.n372 GND.n369 19.3944
R17356 GND.n369 GND.n366 19.3944
R17357 GND.n366 GND.n365 19.3944
R17358 GND.n365 GND.n362 19.3944
R17359 GND.n362 GND.n361 19.3944
R17360 GND.n361 GND.n358 19.3944
R17361 GND.n358 GND.n357 19.3944
R17362 GND.n5128 GND.n5125 19.3944
R17363 GND.n5128 GND.n5122 19.3944
R17364 GND.n5134 GND.n5122 19.3944
R17365 GND.n5134 GND.n5120 19.3944
R17366 GND.n5138 GND.n5120 19.3944
R17367 GND.n5138 GND.n5118 19.3944
R17368 GND.n5144 GND.n5118 19.3944
R17369 GND.n5144 GND.n5116 19.3944
R17370 GND.n5148 GND.n5116 19.3944
R17371 GND.n4912 GND.n4911 19.3944
R17372 GND.n4913 GND.n4912 19.3944
R17373 GND.n4913 GND.n2894 19.3944
R17374 GND.n4919 GND.n2894 19.3944
R17375 GND.n4920 GND.n4919 19.3944
R17376 GND.n4937 GND.n4920 19.3944
R17377 GND.n4937 GND.n2892 19.3944
R17378 GND.n4941 GND.n2892 19.3944
R17379 GND.n4941 GND.n2830 19.3944
R17380 GND.n4952 GND.n2830 19.3944
R17381 GND.n4952 GND.n2828 19.3944
R17382 GND.n4956 GND.n2828 19.3944
R17383 GND.n4956 GND.n2826 19.3944
R17384 GND.n4967 GND.n2826 19.3944
R17385 GND.n4967 GND.n2824 19.3944
R17386 GND.n4971 GND.n2824 19.3944
R17387 GND.n4971 GND.n2822 19.3944
R17388 GND.n4982 GND.n2822 19.3944
R17389 GND.n4982 GND.n2820 19.3944
R17390 GND.n4986 GND.n2820 19.3944
R17391 GND.n4986 GND.n2818 19.3944
R17392 GND.n4997 GND.n2818 19.3944
R17393 GND.n4997 GND.n2816 19.3944
R17394 GND.n5011 GND.n2816 19.3944
R17395 GND.n5011 GND.n5010 19.3944
R17396 GND.n5010 GND.n5009 19.3944
R17397 GND.n5009 GND.n5008 19.3944
R17398 GND.n5008 GND.n5005 19.3944
R17399 GND.n5005 GND.n24 19.3944
R17400 GND.n7826 GND.n24 19.3944
R17401 GND.n7826 GND.n25 19.3944
R17402 GND.n5035 GND.n25 19.3944
R17403 GND.n5038 GND.n5035 19.3944
R17404 GND.n5038 GND.n2812 19.3944
R17405 GND.n5049 GND.n2812 19.3944
R17406 GND.n5049 GND.n2810 19.3944
R17407 GND.n5053 GND.n2810 19.3944
R17408 GND.n5053 GND.n2807 19.3944
R17409 GND.n5063 GND.n2807 19.3944
R17410 GND.n5063 GND.n2805 19.3944
R17411 GND.n5067 GND.n2805 19.3944
R17412 GND.n5067 GND.n2802 19.3944
R17413 GND.n5077 GND.n2802 19.3944
R17414 GND.n5077 GND.n2800 19.3944
R17415 GND.n5081 GND.n2800 19.3944
R17416 GND.n5081 GND.n2797 19.3944
R17417 GND.n5091 GND.n2797 19.3944
R17418 GND.n5091 GND.n2795 19.3944
R17419 GND.n5096 GND.n2795 19.3944
R17420 GND.n5096 GND.n2788 19.3944
R17421 GND.n5177 GND.n2788 19.3944
R17422 GND.n5177 GND.n5176 19.3944
R17423 GND.n5176 GND.n5175 19.3944
R17424 GND.n5175 GND.n2792 19.3944
R17425 GND.n5165 GND.n2792 19.3944
R17426 GND.n5165 GND.n5164 19.3944
R17427 GND.n5164 GND.n5163 19.3944
R17428 GND.n5163 GND.n5157 19.3944
R17429 GND.n5157 GND.n5156 19.3944
R17430 GND.n2905 GND.n2903 19.3944
R17431 GND.n2909 GND.n2905 19.3944
R17432 GND.n2911 GND.n2909 19.3944
R17433 GND.n2915 GND.n2911 19.3944
R17434 GND.n2917 GND.n2915 19.3944
R17435 GND.n2921 GND.n2917 19.3944
R17436 GND.n2923 GND.n2921 19.3944
R17437 GND.n2927 GND.n2923 19.3944
R17438 GND.n2930 GND.n2927 19.3944
R17439 GND.n4261 GND.n3078 19.3944
R17440 GND.n4261 GND.n3077 19.3944
R17441 GND.n4270 GND.n3077 19.3944
R17442 GND.n4270 GND.n4269 19.3944
R17443 GND.n4269 GND.n4268 19.3944
R17444 GND.n4268 GND.n3061 19.3944
R17445 GND.n4299 GND.n3061 19.3944
R17446 GND.n4299 GND.n3059 19.3944
R17447 GND.n4318 GND.n3059 19.3944
R17448 GND.n4318 GND.n4317 19.3944
R17449 GND.n4317 GND.n4316 19.3944
R17450 GND.n4316 GND.n4305 19.3944
R17451 GND.n4312 GND.n4305 19.3944
R17452 GND.n4312 GND.n4311 19.3944
R17453 GND.n4311 GND.n3047 19.3944
R17454 GND.n4419 GND.n3047 19.3944
R17455 GND.n4420 GND.n4419 19.3944
R17456 GND.n4420 GND.n3045 19.3944
R17457 GND.n4424 GND.n3045 19.3944
R17458 GND.n4424 GND.n3043 19.3944
R17459 GND.n4428 GND.n3043 19.3944
R17460 GND.n4428 GND.n3041 19.3944
R17461 GND.n4440 GND.n3041 19.3944
R17462 GND.n4440 GND.n4439 19.3944
R17463 GND.n4439 GND.n4438 19.3944
R17464 GND.n4438 GND.n4436 19.3944
R17465 GND.n4436 GND.n3016 19.3944
R17466 GND.n3016 GND.n3014 19.3944
R17467 GND.n4464 GND.n3014 19.3944
R17468 GND.n4464 GND.n3012 19.3944
R17469 GND.n4485 GND.n3012 19.3944
R17470 GND.n4485 GND.n4484 19.3944
R17471 GND.n4484 GND.n4483 19.3944
R17472 GND.n4483 GND.n4479 19.3944
R17473 GND.n4479 GND.n4478 19.3944
R17474 GND.n4478 GND.n4477 19.3944
R17475 GND.n4477 GND.n4474 19.3944
R17476 GND.n4474 GND.n2993 19.3944
R17477 GND.n4536 GND.n2993 19.3944
R17478 GND.n4536 GND.n2991 19.3944
R17479 GND.n4542 GND.n2991 19.3944
R17480 GND.n4542 GND.n4541 19.3944
R17481 GND.n4541 GND.n2986 19.3944
R17482 GND.n4564 GND.n2986 19.3944
R17483 GND.n4564 GND.n2984 19.3944
R17484 GND.n4568 GND.n2984 19.3944
R17485 GND.n4568 GND.n2982 19.3944
R17486 GND.n4572 GND.n2982 19.3944
R17487 GND.n4572 GND.n2980 19.3944
R17488 GND.n4576 GND.n2980 19.3944
R17489 GND.n4576 GND.n2978 19.3944
R17490 GND.n4633 GND.n2978 19.3944
R17491 GND.n4633 GND.n2976 19.3944
R17492 GND.n4638 GND.n2976 19.3944
R17493 GND.n4638 GND.n2966 19.3944
R17494 GND.n4676 GND.n2966 19.3944
R17495 GND.n4677 GND.n4676 19.3944
R17496 GND.n4679 GND.n4677 19.3944
R17497 GND.n4679 GND.n2964 19.3944
R17498 GND.n4683 GND.n2964 19.3944
R17499 GND.n4683 GND.n2956 19.3944
R17500 GND.n4696 GND.n2956 19.3944
R17501 GND.n4696 GND.n2954 19.3944
R17502 GND.n4700 GND.n2954 19.3944
R17503 GND.n4700 GND.n2950 19.3944
R17504 GND.n4740 GND.n2950 19.3944
R17505 GND.n4740 GND.n2948 19.3944
R17506 GND.n4750 GND.n2948 19.3944
R17507 GND.n4750 GND.n4749 19.3944
R17508 GND.n4749 GND.n4748 19.3944
R17509 GND.n4748 GND.n2933 19.3944
R17510 GND.n4794 GND.n2933 19.3944
R17511 GND.n4795 GND.n4794 19.3944
R17512 GND.n4795 GND.n2414 19.3944
R17513 GND.n5485 GND.n5484 19.3944
R17514 GND.n5484 GND.n5481 19.3944
R17515 GND.n5481 GND.n5480 19.3944
R17516 GND.n5523 GND.n2376 19.3944
R17517 GND.n5518 GND.n2376 19.3944
R17518 GND.n5518 GND.n5517 19.3944
R17519 GND.n5517 GND.n5516 19.3944
R17520 GND.n5516 GND.n5513 19.3944
R17521 GND.n5513 GND.n5512 19.3944
R17522 GND.n5512 GND.n5509 19.3944
R17523 GND.n5509 GND.n5508 19.3944
R17524 GND.n5508 GND.n5505 19.3944
R17525 GND.n5505 GND.n5504 19.3944
R17526 GND.n5504 GND.n5501 19.3944
R17527 GND.n5501 GND.n5500 19.3944
R17528 GND.n5500 GND.n5497 19.3944
R17529 GND.n5497 GND.n5496 19.3944
R17530 GND.n5496 GND.n5493 19.3944
R17531 GND.n5493 GND.n5492 19.3944
R17532 GND.n5492 GND.n5489 19.3944
R17533 GND.n5489 GND.n5488 19.3944
R17534 GND.n4254 GND.n1975 19.3944
R17535 GND.n5776 GND.n1975 19.3944
R17536 GND.n5776 GND.n5775 19.3944
R17537 GND.n5775 GND.n5774 19.3944
R17538 GND.n5774 GND.n1979 19.3944
R17539 GND.n3067 GND.n1979 19.3944
R17540 GND.n3067 GND.n2021 19.3944
R17541 GND.n5755 GND.n2021 19.3944
R17542 GND.n5755 GND.n5754 19.3944
R17543 GND.n5754 GND.n5753 19.3944
R17544 GND.n5753 GND.n2025 19.3944
R17545 GND.n2069 GND.n2025 19.3944
R17546 GND.n2072 GND.n2069 19.3944
R17547 GND.n2072 GND.n2066 19.3944
R17548 GND.n5728 GND.n2066 19.3944
R17549 GND.n5728 GND.n5727 19.3944
R17550 GND.n5727 GND.n5726 19.3944
R17551 GND.n5726 GND.n2078 19.3944
R17552 GND.n3029 GND.n2078 19.3944
R17553 GND.n3029 GND.n3026 19.3944
R17554 GND.n3033 GND.n3026 19.3944
R17555 GND.n3033 GND.n3024 19.3944
R17556 GND.n3037 GND.n3024 19.3944
R17557 GND.n3037 GND.n3022 19.3944
R17558 GND.n4446 GND.n3022 19.3944
R17559 GND.n4446 GND.n3020 19.3944
R17560 GND.n4458 GND.n3020 19.3944
R17561 GND.n4458 GND.n4457 19.3944
R17562 GND.n4457 GND.n4456 19.3944
R17563 GND.n4456 GND.n4454 19.3944
R17564 GND.n4454 GND.n3009 19.3944
R17565 GND.n3009 GND.n3007 19.3944
R17566 GND.n4491 GND.n3007 19.3944
R17567 GND.n4491 GND.n3005 19.3944
R17568 GND.n4504 GND.n3005 19.3944
R17569 GND.n4504 GND.n4503 19.3944
R17570 GND.n4503 GND.n4502 19.3944
R17571 GND.n4502 GND.n4499 19.3944
R17572 GND.n4499 GND.n2190 19.3944
R17573 GND.n5644 GND.n2190 19.3944
R17574 GND.n5644 GND.n5643 19.3944
R17575 GND.n5643 GND.n5642 19.3944
R17576 GND.n5642 GND.n2194 19.3944
R17577 GND.n4605 GND.n2194 19.3944
R17578 GND.n4605 GND.n4602 19.3944
R17579 GND.n4609 GND.n4602 19.3944
R17580 GND.n4609 GND.n4600 19.3944
R17581 GND.n4613 GND.n4600 19.3944
R17582 GND.n4613 GND.n4598 19.3944
R17583 GND.n4627 GND.n4598 19.3944
R17584 GND.n4627 GND.n4626 19.3944
R17585 GND.n4626 GND.n4625 19.3944
R17586 GND.n4625 GND.n4621 19.3944
R17587 GND.n4621 GND.n2274 19.3944
R17588 GND.n5590 GND.n2274 19.3944
R17589 GND.n5590 GND.n5589 19.3944
R17590 GND.n5589 GND.n5588 19.3944
R17591 GND.n5588 GND.n2278 19.3944
R17592 GND.n2313 GND.n2278 19.3944
R17593 GND.n2313 GND.n2310 19.3944
R17594 GND.n5569 GND.n2310 19.3944
R17595 GND.n5569 GND.n5568 19.3944
R17596 GND.n5568 GND.n5567 19.3944
R17597 GND.n5567 GND.n2319 19.3944
R17598 GND.n5555 GND.n2319 19.3944
R17599 GND.n5555 GND.n5554 19.3944
R17600 GND.n5554 GND.n5553 19.3944
R17601 GND.n5553 GND.n2339 19.3944
R17602 GND.n5541 GND.n2339 19.3944
R17603 GND.n5541 GND.n5540 19.3944
R17604 GND.n5540 GND.n5539 19.3944
R17605 GND.n5539 GND.n2359 19.3944
R17606 GND.n5527 GND.n2359 19.3944
R17607 GND.n5527 GND.n5526 19.3944
R17608 GND.n4197 GND.n4179 19.3944
R17609 GND.n4190 GND.n4179 19.3944
R17610 GND.n4190 GND.n4189 19.3944
R17611 GND.n4250 GND.n4249 19.3944
R17612 GND.n4249 GND.n3083 19.3944
R17613 GND.n4244 GND.n3083 19.3944
R17614 GND.n4244 GND.n4243 19.3944
R17615 GND.n4243 GND.n3088 19.3944
R17616 GND.n4238 GND.n3088 19.3944
R17617 GND.n4238 GND.n4237 19.3944
R17618 GND.n4237 GND.n4236 19.3944
R17619 GND.n4236 GND.n3094 19.3944
R17620 GND.n4230 GND.n3094 19.3944
R17621 GND.n4230 GND.n3096 19.3944
R17622 GND.n4217 GND.n3096 19.3944
R17623 GND.n4217 GND.n4216 19.3944
R17624 GND.n4216 GND.n4156 19.3944
R17625 GND.n4209 GND.n4156 19.3944
R17626 GND.n4209 GND.n4208 19.3944
R17627 GND.n4208 GND.n4169 19.3944
R17628 GND.n4201 GND.n4169 19.3944
R17629 GND.n5335 GND.n5334 19.3944
R17630 GND.n5334 GND.n2592 19.3944
R17631 GND.n2628 GND.n2592 19.3944
R17632 GND.n2628 GND.n2625 19.3944
R17633 GND.n5315 GND.n2625 19.3944
R17634 GND.n5315 GND.n5314 19.3944
R17635 GND.n5314 GND.n5313 19.3944
R17636 GND.n5313 GND.n2634 19.3944
R17637 GND.n5303 GND.n2634 19.3944
R17638 GND.n5303 GND.n5302 19.3944
R17639 GND.n5302 GND.n5301 19.3944
R17640 GND.n5301 GND.n2656 19.3944
R17641 GND.n5291 GND.n2656 19.3944
R17642 GND.n5291 GND.n5290 19.3944
R17643 GND.n5290 GND.n5289 19.3944
R17644 GND.n5289 GND.n2677 19.3944
R17645 GND.n5279 GND.n2677 19.3944
R17646 GND.n5279 GND.n5278 19.3944
R17647 GND.n5278 GND.n5277 19.3944
R17648 GND.n5277 GND.n2698 19.3944
R17649 GND.n5267 GND.n2698 19.3944
R17650 GND.n5267 GND.n5266 19.3944
R17651 GND.n5266 GND.n5265 19.3944
R17652 GND.n5265 GND.n2719 19.3944
R17653 GND.n5255 GND.n2719 19.3944
R17654 GND.n2735 GND.n41 19.3944
R17655 GND.n2745 GND.n41 19.3944
R17656 GND.n7822 GND.n34 19.3944
R17657 GND.n2757 GND.n35 19.3944
R17658 GND.n7819 GND.n43 19.3944
R17659 GND.n7819 GND.n44 19.3944
R17660 GND.n7809 GND.n44 19.3944
R17661 GND.n7809 GND.n7808 19.3944
R17662 GND.n7808 GND.n7807 19.3944
R17663 GND.n7807 GND.n66 19.3944
R17664 GND.n7797 GND.n66 19.3944
R17665 GND.n7797 GND.n7796 19.3944
R17666 GND.n7796 GND.n7795 19.3944
R17667 GND.n7795 GND.n87 19.3944
R17668 GND.n7785 GND.n87 19.3944
R17669 GND.n7785 GND.n7784 19.3944
R17670 GND.n7784 GND.n7783 19.3944
R17671 GND.n7783 GND.n108 19.3944
R17672 GND.n7773 GND.n108 19.3944
R17673 GND.n7773 GND.n7772 19.3944
R17674 GND.n7772 GND.n7771 19.3944
R17675 GND.n7771 GND.n129 19.3944
R17676 GND.n7761 GND.n129 19.3944
R17677 GND.n7761 GND.n7760 19.3944
R17678 GND.n7760 GND.n7759 19.3944
R17679 GND.n7759 GND.n149 19.3944
R17680 GND.n7749 GND.n149 19.3944
R17681 GND.n7749 GND.n7748 19.3944
R17682 GND.n7748 GND.n7747 19.3944
R17683 GND.n7747 GND.n170 19.3944
R17684 GND.n6170 GND.n1448 19.3944
R17685 GND.n6170 GND.n6169 19.3944
R17686 GND.n6169 GND.n6168 19.3944
R17687 GND.n6168 GND.n1453 19.3944
R17688 GND.n6162 GND.n1453 19.3944
R17689 GND.n6162 GND.n6161 19.3944
R17690 GND.n6161 GND.n6160 19.3944
R17691 GND.n6160 GND.n1461 19.3944
R17692 GND.n6154 GND.n1461 19.3944
R17693 GND.n6154 GND.n6153 19.3944
R17694 GND.n6153 GND.n6152 19.3944
R17695 GND.n6152 GND.n1469 19.3944
R17696 GND.n6146 GND.n1469 19.3944
R17697 GND.n6146 GND.n6145 19.3944
R17698 GND.n6145 GND.n6144 19.3944
R17699 GND.n6144 GND.n1477 19.3944
R17700 GND.n6138 GND.n1477 19.3944
R17701 GND.n6138 GND.n6137 19.3944
R17702 GND.n6137 GND.n6136 19.3944
R17703 GND.n6136 GND.n1485 19.3944
R17704 GND.n6130 GND.n1485 19.3944
R17705 GND.n6130 GND.n6129 19.3944
R17706 GND.n6129 GND.n6128 19.3944
R17707 GND.n6128 GND.n1493 19.3944
R17708 GND.n6122 GND.n1493 19.3944
R17709 GND.n6122 GND.n6121 19.3944
R17710 GND.n6121 GND.n6120 19.3944
R17711 GND.n6120 GND.n1501 19.3944
R17712 GND.n6114 GND.n1501 19.3944
R17713 GND.n6114 GND.n6113 19.3944
R17714 GND.n6113 GND.n6112 19.3944
R17715 GND.n6112 GND.n1509 19.3944
R17716 GND.n6106 GND.n1509 19.3944
R17717 GND.n6106 GND.n6105 19.3944
R17718 GND.n6105 GND.n6104 19.3944
R17719 GND.n6104 GND.n1517 19.3944
R17720 GND.n6098 GND.n1517 19.3944
R17721 GND.n6098 GND.n6097 19.3944
R17722 GND.n6097 GND.n6096 19.3944
R17723 GND.n6096 GND.n1525 19.3944
R17724 GND.n6090 GND.n1525 19.3944
R17725 GND.n6090 GND.n6089 19.3944
R17726 GND.n6089 GND.n6088 19.3944
R17727 GND.n6088 GND.n1533 19.3944
R17728 GND.n6082 GND.n1533 19.3944
R17729 GND.n6082 GND.n6081 19.3944
R17730 GND.n6081 GND.n6080 19.3944
R17731 GND.n6080 GND.n1541 19.3944
R17732 GND.n6074 GND.n1541 19.3944
R17733 GND.n6074 GND.n6073 19.3944
R17734 GND.n6073 GND.n6072 19.3944
R17735 GND.n6072 GND.n1549 19.3944
R17736 GND.n6066 GND.n1549 19.3944
R17737 GND.n6066 GND.n6065 19.3944
R17738 GND.n6065 GND.n6064 19.3944
R17739 GND.n6064 GND.n1557 19.3944
R17740 GND.n6058 GND.n1557 19.3944
R17741 GND.n6058 GND.n6057 19.3944
R17742 GND.n6057 GND.n6056 19.3944
R17743 GND.n6056 GND.n1565 19.3944
R17744 GND.n6050 GND.n1565 19.3944
R17745 GND.n6050 GND.n6049 19.3944
R17746 GND.n6049 GND.n6048 19.3944
R17747 GND.n6048 GND.n1573 19.3944
R17748 GND.n6042 GND.n1573 19.3944
R17749 GND.n6042 GND.n6041 19.3944
R17750 GND.n6041 GND.n6040 19.3944
R17751 GND.n6040 GND.n1581 19.3944
R17752 GND.n6034 GND.n1581 19.3944
R17753 GND.n6034 GND.n6033 19.3944
R17754 GND.n6033 GND.n6032 19.3944
R17755 GND.n6032 GND.n1589 19.3944
R17756 GND.n6026 GND.n1589 19.3944
R17757 GND.n6026 GND.n6025 19.3944
R17758 GND.n6025 GND.n6024 19.3944
R17759 GND.n6024 GND.n1597 19.3944
R17760 GND.n6018 GND.n1597 19.3944
R17761 GND.n6018 GND.n6017 19.3944
R17762 GND.n6017 GND.n6016 19.3944
R17763 GND.n6016 GND.n1605 19.3944
R17764 GND.n6010 GND.n1605 19.3944
R17765 GND.n6010 GND.n6009 19.3944
R17766 GND.n6009 GND.n6008 19.3944
R17767 GND.n6008 GND.n1613 19.3944
R17768 GND.n3485 GND.n1613 19.3944
R17769 GND.n3489 GND.n3485 19.3944
R17770 GND.n3489 GND.n3473 19.3944
R17771 GND.n3682 GND.n3473 19.3944
R17772 GND.n3682 GND.n3471 19.3944
R17773 GND.n3688 GND.n3471 19.3944
R17774 GND.n3688 GND.n3687 19.3944
R17775 GND.n3687 GND.n3443 19.3944
R17776 GND.n3719 GND.n3443 19.3944
R17777 GND.n3719 GND.n3441 19.3944
R17778 GND.n3725 GND.n3441 19.3944
R17779 GND.n3725 GND.n3724 19.3944
R17780 GND.n3724 GND.n3414 19.3944
R17781 GND.n3756 GND.n3414 19.3944
R17782 GND.n3756 GND.n3412 19.3944
R17783 GND.n3762 GND.n3412 19.3944
R17784 GND.n3762 GND.n3761 19.3944
R17785 GND.n3761 GND.n3385 19.3944
R17786 GND.n3793 GND.n3385 19.3944
R17787 GND.n3793 GND.n3383 19.3944
R17788 GND.n3805 GND.n3383 19.3944
R17789 GND.n3805 GND.n3804 19.3944
R17790 GND.n3804 GND.n3803 19.3944
R17791 GND.n3803 GND.n3800 19.3944
R17792 GND.n3800 GND.n3332 19.3944
R17793 GND.n3940 GND.n3332 19.3944
R17794 GND.n3940 GND.n3333 19.3944
R17795 GND.n3872 GND.n3871 19.3944
R17796 GND.n3875 GND.n3874 19.3944
R17797 GND.n3898 GND.n3897 19.3944
R17798 GND.n3895 GND.n3894 19.3944
R17799 GND.n3891 GND.n3324 19.3944
R17800 GND.n3945 GND.n3324 19.3944
R17801 GND.n3945 GND.n3299 19.3944
R17802 GND.n3976 GND.n3299 19.3944
R17803 GND.n3976 GND.n3297 19.3944
R17804 GND.n3982 GND.n3297 19.3944
R17805 GND.n3982 GND.n3981 19.3944
R17806 GND.n3981 GND.n3269 19.3944
R17807 GND.n4013 GND.n3269 19.3944
R17808 GND.n4013 GND.n3267 19.3944
R17809 GND.n4019 GND.n3267 19.3944
R17810 GND.n4019 GND.n4018 19.3944
R17811 GND.n4018 GND.n3240 19.3944
R17812 GND.n4050 GND.n3240 19.3944
R17813 GND.n4050 GND.n3238 19.3944
R17814 GND.n4056 GND.n3238 19.3944
R17815 GND.n4056 GND.n4055 19.3944
R17816 GND.n4055 GND.n3211 19.3944
R17817 GND.n4087 GND.n3211 19.3944
R17818 GND.n4087 GND.n3209 19.3944
R17819 GND.n4126 GND.n3209 19.3944
R17820 GND.n4126 GND.n4125 19.3944
R17821 GND.n4125 GND.n4124 19.3944
R17822 GND.n4124 GND.n4093 19.3944
R17823 GND.n4120 GND.n4093 19.3944
R17824 GND.n4120 GND.n4119 19.3944
R17825 GND.n4119 GND.n4118 19.3944
R17826 GND.n4118 GND.n4099 19.3944
R17827 GND.n4112 GND.n4099 19.3944
R17828 GND.n4112 GND.n4111 19.3944
R17829 GND.n4111 GND.n4110 19.3944
R17830 GND.n4110 GND.n4107 19.3944
R17831 GND.n4107 GND.n1888 19.3944
R17832 GND.n5801 GND.n1888 19.3944
R17833 GND.n5801 GND.n5800 19.3944
R17834 GND.n5800 GND.n5799 19.3944
R17835 GND.n5799 GND.n1892 19.3944
R17836 GND.n2000 GND.n1892 19.3944
R17837 GND.n2000 GND.n1997 19.3944
R17838 GND.n2004 GND.n1997 19.3944
R17839 GND.n2004 GND.n1995 19.3944
R17840 GND.n2008 GND.n1995 19.3944
R17841 GND.n2008 GND.n1993 19.3944
R17842 GND.n5762 GND.n1993 19.3944
R17843 GND.n5762 GND.n5761 19.3944
R17844 GND.n5761 GND.n5760 19.3944
R17845 GND.n5760 GND.n2014 19.3944
R17846 GND.n2044 GND.n2014 19.3944
R17847 GND.n2044 GND.n2041 19.3944
R17848 GND.n5742 GND.n2041 19.3944
R17849 GND.n5742 GND.n5741 19.3944
R17850 GND.n5741 GND.n5740 19.3944
R17851 GND.n5740 GND.n2050 19.3944
R17852 GND.n2088 GND.n2050 19.3944
R17853 GND.n2088 GND.n2085 19.3944
R17854 GND.n5721 GND.n2085 19.3944
R17855 GND.n5721 GND.n5720 19.3944
R17856 GND.n5720 GND.n5719 19.3944
R17857 GND.n5719 GND.n2094 19.3944
R17858 GND.n5707 GND.n2094 19.3944
R17859 GND.n5707 GND.n5706 19.3944
R17860 GND.n5706 GND.n5705 19.3944
R17861 GND.n5705 GND.n2112 19.3944
R17862 GND.n5693 GND.n2112 19.3944
R17863 GND.n5693 GND.n5692 19.3944
R17864 GND.n5692 GND.n5691 19.3944
R17865 GND.n5691 GND.n2130 19.3944
R17866 GND.n5679 GND.n2130 19.3944
R17867 GND.n5679 GND.n5678 19.3944
R17868 GND.n5678 GND.n5677 19.3944
R17869 GND.n5677 GND.n2147 19.3944
R17870 GND.n5665 GND.n2147 19.3944
R17871 GND.n5665 GND.n5664 19.3944
R17872 GND.n5664 GND.n5663 19.3944
R17873 GND.n5663 GND.n2165 19.3944
R17874 GND.n5651 GND.n2165 19.3944
R17875 GND.n5651 GND.n5650 19.3944
R17876 GND.n5650 GND.n5649 19.3944
R17877 GND.n5649 GND.n2183 19.3944
R17878 GND.n2212 GND.n2183 19.3944
R17879 GND.n2212 GND.n2209 19.3944
R17880 GND.n5630 GND.n2209 19.3944
R17881 GND.n5630 GND.n5629 19.3944
R17882 GND.n5629 GND.n5628 19.3944
R17883 GND.n5628 GND.n2218 19.3944
R17884 GND.n2243 GND.n2218 19.3944
R17885 GND.n5611 GND.n2243 19.3944
R17886 GND.n5611 GND.n5610 19.3944
R17887 GND.n5610 GND.n5609 19.3944
R17888 GND.n5609 GND.n2249 19.3944
R17889 GND.n5597 GND.n2249 19.3944
R17890 GND.n5597 GND.n5596 19.3944
R17891 GND.n5596 GND.n5595 19.3944
R17892 GND.n5595 GND.n2267 19.3944
R17893 GND.n2297 GND.n2267 19.3944
R17894 GND.n2297 GND.n2294 19.3944
R17895 GND.n5576 GND.n2294 19.3944
R17896 GND.n5576 GND.n5575 19.3944
R17897 GND.n5575 GND.n5574 19.3944
R17898 GND.n5574 GND.n2303 19.3944
R17899 GND.n4722 GND.n2303 19.3944
R17900 GND.n4722 GND.n4719 19.3944
R17901 GND.n4726 GND.n4719 19.3944
R17902 GND.n4726 GND.n4717 19.3944
R17903 GND.n4735 GND.n4717 19.3944
R17904 GND.n4735 GND.n4734 19.3944
R17905 GND.n4734 GND.n4733 19.3944
R17906 GND.n4733 GND.n2939 19.3944
R17907 GND.n4771 GND.n2939 19.3944
R17908 GND.n4771 GND.n2937 19.3944
R17909 GND.n4788 GND.n2937 19.3944
R17910 GND.n4788 GND.n4787 19.3944
R17911 GND.n4787 GND.n4786 19.3944
R17912 GND.n4786 GND.n4777 19.3944
R17913 GND.n4781 GND.n4777 19.3944
R17914 GND.n4781 GND.n2437 19.3944
R17915 GND.n5455 GND.n2437 19.3944
R17916 GND.n5455 GND.n5454 19.3944
R17917 GND.n5454 GND.n5453 19.3944
R17918 GND.n5453 GND.n2441 19.3944
R17919 GND.n4809 GND.n2441 19.3944
R17920 GND.n4809 GND.n4806 19.3944
R17921 GND.n4816 GND.n4806 19.3944
R17922 GND.n4816 GND.n4804 19.3944
R17923 GND.n4823 GND.n4804 19.3944
R17924 GND.n4823 GND.n4822 19.3944
R17925 GND.n4822 GND.n2611 19.3944
R17926 GND.n5322 GND.n2611 19.3944
R17927 GND.n5322 GND.n5321 19.3944
R17928 GND.n5321 GND.n5320 19.3944
R17929 GND.n5320 GND.n2615 19.3944
R17930 GND.n2834 GND.n2615 19.3944
R17931 GND.n2889 GND.n2834 19.3944
R17932 GND.n2889 GND.n2888 19.3944
R17933 GND.n2888 GND.n2887 19.3944
R17934 GND.n2887 GND.n2840 19.3944
R17935 GND.n2883 GND.n2840 19.3944
R17936 GND.n2883 GND.n2882 19.3944
R17937 GND.n2882 GND.n2881 19.3944
R17938 GND.n2881 GND.n2846 19.3944
R17939 GND.n2877 GND.n2846 19.3944
R17940 GND.n2877 GND.n2876 19.3944
R17941 GND.n2876 GND.n2875 19.3944
R17942 GND.n2875 GND.n2852 19.3944
R17943 GND.n2871 GND.n2852 19.3944
R17944 GND.n2871 GND.n2870 19.3944
R17945 GND.n2870 GND.n2869 19.3944
R17946 GND.n2869 GND.n2858 19.3944
R17947 GND.n2865 GND.n2858 19.3944
R17948 GND.n2865 GND.n2864 19.3944
R17949 GND.n2864 GND.n2863 19.3944
R17950 GND.n5250 GND.n5249 19.3944
R17951 GND.n5247 GND.n2742 19.3944
R17952 GND.n5235 GND.n2763 19.3944
R17953 GND.n5233 GND.n5232 19.3944
R17954 GND.n5229 GND.n5228 19.3944
R17955 GND.n5228 GND.n5227 19.3944
R17956 GND.n5227 GND.n2768 19.3944
R17957 GND.n5223 GND.n2768 19.3944
R17958 GND.n5223 GND.n5222 19.3944
R17959 GND.n5222 GND.n5221 19.3944
R17960 GND.n5221 GND.n2774 19.3944
R17961 GND.n5217 GND.n2774 19.3944
R17962 GND.n5217 GND.n5216 19.3944
R17963 GND.n5216 GND.n5215 19.3944
R17964 GND.n5215 GND.n2780 19.3944
R17965 GND.n5211 GND.n2780 19.3944
R17966 GND.n5211 GND.n5210 19.3944
R17967 GND.n5210 GND.n5209 19.3944
R17968 GND.n5209 GND.n2786 19.3944
R17969 GND.n5205 GND.n2786 19.3944
R17970 GND.n5205 GND.n5204 19.3944
R17971 GND.n5204 GND.n5203 19.3944
R17972 GND.n5203 GND.n5186 19.3944
R17973 GND.n5199 GND.n5186 19.3944
R17974 GND.n5199 GND.n5198 19.3944
R17975 GND.n5198 GND.n5197 19.3944
R17976 GND.n5197 GND.n5194 19.3944
R17977 GND.n5194 GND.n185 19.3944
R17978 GND.n7735 GND.n185 19.3944
R17979 GND.n7735 GND.n7734 19.3944
R17980 GND.n7734 GND.n7733 19.3944
R17981 GND.n7733 GND.n189 19.3944
R17982 GND.n7727 GND.n189 19.3944
R17983 GND.n7727 GND.n7726 19.3944
R17984 GND.n7726 GND.n7725 19.3944
R17985 GND.n7725 GND.n386 19.3944
R17986 GND.n7719 GND.n386 19.3944
R17987 GND.n7719 GND.n7718 19.3944
R17988 GND.n7718 GND.n7717 19.3944
R17989 GND.n7717 GND.n394 19.3944
R17990 GND.n7711 GND.n394 19.3944
R17991 GND.n7711 GND.n7710 19.3944
R17992 GND.n7710 GND.n7709 19.3944
R17993 GND.n7709 GND.n402 19.3944
R17994 GND.n7703 GND.n402 19.3944
R17995 GND.n7703 GND.n7702 19.3944
R17996 GND.n7702 GND.n7701 19.3944
R17997 GND.n7701 GND.n410 19.3944
R17998 GND.n7695 GND.n410 19.3944
R17999 GND.n7695 GND.n7694 19.3944
R18000 GND.n7694 GND.n7693 19.3944
R18001 GND.n7693 GND.n418 19.3944
R18002 GND.n7687 GND.n418 19.3944
R18003 GND.n7687 GND.n7686 19.3944
R18004 GND.n7686 GND.n7685 19.3944
R18005 GND.n7685 GND.n426 19.3944
R18006 GND.n7679 GND.n426 19.3944
R18007 GND.n7679 GND.n7678 19.3944
R18008 GND.n7678 GND.n7677 19.3944
R18009 GND.n7677 GND.n434 19.3944
R18010 GND.n7671 GND.n434 19.3944
R18011 GND.n7671 GND.n7670 19.3944
R18012 GND.n7670 GND.n7669 19.3944
R18013 GND.n7669 GND.n442 19.3944
R18014 GND.n7663 GND.n442 19.3944
R18015 GND.n7663 GND.n7662 19.3944
R18016 GND.n7662 GND.n7661 19.3944
R18017 GND.n7661 GND.n450 19.3944
R18018 GND.n7655 GND.n450 19.3944
R18019 GND.n7655 GND.n7654 19.3944
R18020 GND.n7654 GND.n7653 19.3944
R18021 GND.n7653 GND.n458 19.3944
R18022 GND.n7647 GND.n458 19.3944
R18023 GND.n7647 GND.n7646 19.3944
R18024 GND.n7646 GND.n7645 19.3944
R18025 GND.n7645 GND.n466 19.3944
R18026 GND.n7639 GND.n466 19.3944
R18027 GND.n7639 GND.n7638 19.3944
R18028 GND.n7638 GND.n7637 19.3944
R18029 GND.n7637 GND.n474 19.3944
R18030 GND.n7631 GND.n474 19.3944
R18031 GND.n7631 GND.n7630 19.3944
R18032 GND.n7630 GND.n7629 19.3944
R18033 GND.n7629 GND.n482 19.3944
R18034 GND.n7623 GND.n482 19.3944
R18035 GND.n7623 GND.n7622 19.3944
R18036 GND.n7622 GND.n7621 19.3944
R18037 GND.n7621 GND.n490 19.3944
R18038 GND.n7615 GND.n490 19.3944
R18039 GND.n7615 GND.n7614 19.3944
R18040 GND.n7614 GND.n7613 19.3944
R18041 GND.n7613 GND.n498 19.3944
R18042 GND.n7607 GND.n498 19.3944
R18043 GND.n7607 GND.n7606 19.3944
R18044 GND.n7606 GND.n7605 19.3944
R18045 GND.n7605 GND.n506 19.3944
R18046 GND.n7599 GND.n506 19.3944
R18047 GND.n7599 GND.n7598 19.3944
R18048 GND.n7598 GND.n7597 19.3944
R18049 GND.n7597 GND.n514 19.3944
R18050 GND.n7591 GND.n514 19.3944
R18051 GND.n7591 GND.n7590 19.3944
R18052 GND.n7590 GND.n7589 19.3944
R18053 GND.n7589 GND.n522 19.3944
R18054 GND.n7583 GND.n522 19.3944
R18055 GND.n7583 GND.n7582 19.3944
R18056 GND.n7582 GND.n7581 19.3944
R18057 GND.n7581 GND.n530 19.3944
R18058 GND.n7575 GND.n530 19.3944
R18059 GND.n7575 GND.n7574 19.3944
R18060 GND.n7574 GND.n7573 19.3944
R18061 GND.n7573 GND.n538 19.3944
R18062 GND.n7567 GND.n538 19.3944
R18063 GND.n7567 GND.n7566 19.3944
R18064 GND.n7566 GND.n7565 19.3944
R18065 GND.n3528 GND.n3527 19.3944
R18066 GND.n3531 GND.n3528 19.3944
R18067 GND.n3531 GND.n3525 19.3944
R18068 GND.n3537 GND.n3525 19.3944
R18069 GND.n3538 GND.n3537 19.3944
R18070 GND.n3541 GND.n3538 19.3944
R18071 GND.n3541 GND.n3523 19.3944
R18072 GND.n3547 GND.n3523 19.3944
R18073 GND.n3548 GND.n3547 19.3944
R18074 GND.n3551 GND.n3548 19.3944
R18075 GND.n3557 GND.n3554 19.3944
R18076 GND.n3560 GND.n3557 19.3944
R18077 GND.n3560 GND.n3517 19.3944
R18078 GND.n3564 GND.n3517 19.3944
R18079 GND.n3567 GND.n3564 19.3944
R18080 GND.n3570 GND.n3567 19.3944
R18081 GND.n3570 GND.n3515 19.3944
R18082 GND.n3574 GND.n3515 19.3944
R18083 GND.n3577 GND.n3574 19.3944
R18084 GND.n3580 GND.n3577 19.3944
R18085 GND.n3580 GND.n3513 19.3944
R18086 GND.n3584 GND.n3513 19.3944
R18087 GND.n3588 GND.n3587 19.3944
R18088 GND.n3591 GND.n3588 19.3944
R18089 GND.n3591 GND.n3507 19.3944
R18090 GND.n3597 GND.n3507 19.3944
R18091 GND.n3598 GND.n3597 19.3944
R18092 GND.n3601 GND.n3598 19.3944
R18093 GND.n3601 GND.n3505 19.3944
R18094 GND.n3607 GND.n3505 19.3944
R18095 GND.n3608 GND.n3607 19.3944
R18096 GND.n3611 GND.n3608 19.3944
R18097 GND.n3611 GND.n3501 19.3944
R18098 GND.n3621 GND.n3618 19.3944
R18099 GND.n3621 GND.n3499 19.3944
R18100 GND.n3627 GND.n3499 19.3944
R18101 GND.n3628 GND.n3627 19.3944
R18102 GND.n3631 GND.n3628 19.3944
R18103 GND.n3631 GND.n3497 19.3944
R18104 GND.n3637 GND.n3497 19.3944
R18105 GND.n3638 GND.n3637 19.3944
R18106 GND.n3641 GND.n3638 19.3944
R18107 GND.n3641 GND.n3495 19.3944
R18108 GND.n3647 GND.n3495 19.3944
R18109 GND.n3671 GND.n3481 19.3944
R18110 GND.n3677 GND.n3481 19.3944
R18111 GND.n3677 GND.n3676 19.3944
R18112 GND.n3676 GND.n3454 19.3944
R18113 GND.n3708 GND.n3454 19.3944
R18114 GND.n3708 GND.n3452 19.3944
R18115 GND.n3714 GND.n3452 19.3944
R18116 GND.n3714 GND.n3713 19.3944
R18117 GND.n3713 GND.n3425 19.3944
R18118 GND.n3745 GND.n3425 19.3944
R18119 GND.n3745 GND.n3423 19.3944
R18120 GND.n3751 GND.n3423 19.3944
R18121 GND.n3751 GND.n3750 19.3944
R18122 GND.n3750 GND.n3395 19.3944
R18123 GND.n3782 GND.n3395 19.3944
R18124 GND.n3782 GND.n3393 19.3944
R18125 GND.n3788 GND.n3393 19.3944
R18126 GND.n3788 GND.n3787 19.3944
R18127 GND.n3787 GND.n3365 19.3944
R18128 GND.n3819 GND.n3365 19.3944
R18129 GND.n3819 GND.n3363 19.3944
R18130 GND.n3824 GND.n3363 19.3944
R18131 GND.n3824 GND.n3341 19.3944
R18132 GND.n3935 GND.n3341 19.3944
R18133 GND.n3935 GND.n3934 19.3944
R18134 GND.n3932 GND.n3343 19.3944
R18135 GND.n3882 GND.n3343 19.3944
R18136 GND.n3886 GND.n3885 19.3944
R18137 GND.n3907 GND.n3855 19.3944
R18138 GND.n3910 GND.n3909 19.3944
R18139 GND.n3910 GND.n3309 19.3944
R18140 GND.n3965 GND.n3309 19.3944
R18141 GND.n3965 GND.n3307 19.3944
R18142 GND.n3971 GND.n3307 19.3944
R18143 GND.n3971 GND.n3970 19.3944
R18144 GND.n3970 GND.n3280 19.3944
R18145 GND.n4002 GND.n3280 19.3944
R18146 GND.n4002 GND.n3278 19.3944
R18147 GND.n4008 GND.n3278 19.3944
R18148 GND.n4008 GND.n4007 19.3944
R18149 GND.n4007 GND.n3251 19.3944
R18150 GND.n4039 GND.n3251 19.3944
R18151 GND.n4039 GND.n3249 19.3944
R18152 GND.n4045 GND.n3249 19.3944
R18153 GND.n4045 GND.n4044 19.3944
R18154 GND.n4044 GND.n3221 19.3944
R18155 GND.n4076 GND.n3221 19.3944
R18156 GND.n4076 GND.n3219 19.3944
R18157 GND.n4082 GND.n3219 19.3944
R18158 GND.n4082 GND.n4081 19.3944
R18159 GND.n4081 GND.n3194 19.3944
R18160 GND.n4142 GND.n3194 19.3944
R18161 GND.n4142 GND.n3192 19.3944
R18162 GND.n4147 GND.n3192 19.3944
R18163 GND.n4147 GND.n4146 19.3944
R18164 GND.n6353 GND.n6352 19.3944
R18165 GND.n6352 GND.n1269 19.3944
R18166 GND.n6346 GND.n1269 19.3944
R18167 GND.n6346 GND.n6345 19.3944
R18168 GND.n6345 GND.n6344 19.3944
R18169 GND.n6344 GND.n1277 19.3944
R18170 GND.n6338 GND.n1277 19.3944
R18171 GND.n6338 GND.n6337 19.3944
R18172 GND.n6337 GND.n6336 19.3944
R18173 GND.n6336 GND.n1285 19.3944
R18174 GND.n6330 GND.n1285 19.3944
R18175 GND.n6330 GND.n6329 19.3944
R18176 GND.n6329 GND.n6328 19.3944
R18177 GND.n6328 GND.n1293 19.3944
R18178 GND.n6322 GND.n1293 19.3944
R18179 GND.n6322 GND.n6321 19.3944
R18180 GND.n6321 GND.n6320 19.3944
R18181 GND.n6320 GND.n1301 19.3944
R18182 GND.n6314 GND.n1301 19.3944
R18183 GND.n6314 GND.n6313 19.3944
R18184 GND.n6313 GND.n6312 19.3944
R18185 GND.n6312 GND.n1309 19.3944
R18186 GND.n6306 GND.n1309 19.3944
R18187 GND.n6306 GND.n6305 19.3944
R18188 GND.n6305 GND.n6304 19.3944
R18189 GND.n6304 GND.n1317 19.3944
R18190 GND.n6298 GND.n1317 19.3944
R18191 GND.n6298 GND.n6297 19.3944
R18192 GND.n6297 GND.n6296 19.3944
R18193 GND.n6296 GND.n1325 19.3944
R18194 GND.n6290 GND.n1325 19.3944
R18195 GND.n6290 GND.n6289 19.3944
R18196 GND.n6289 GND.n6288 19.3944
R18197 GND.n6288 GND.n1333 19.3944
R18198 GND.n6282 GND.n1333 19.3944
R18199 GND.n6282 GND.n6281 19.3944
R18200 GND.n6281 GND.n6280 19.3944
R18201 GND.n6280 GND.n1341 19.3944
R18202 GND.n6274 GND.n1341 19.3944
R18203 GND.n6274 GND.n6273 19.3944
R18204 GND.n6273 GND.n6272 19.3944
R18205 GND.n6272 GND.n1349 19.3944
R18206 GND.n6266 GND.n1349 19.3944
R18207 GND.n6266 GND.n6265 19.3944
R18208 GND.n6265 GND.n6264 19.3944
R18209 GND.n6264 GND.n1357 19.3944
R18210 GND.n6258 GND.n1357 19.3944
R18211 GND.n6258 GND.n6257 19.3944
R18212 GND.n6257 GND.n6256 19.3944
R18213 GND.n6256 GND.n1365 19.3944
R18214 GND.n6250 GND.n1365 19.3944
R18215 GND.n6250 GND.n6249 19.3944
R18216 GND.n6249 GND.n6248 19.3944
R18217 GND.n6248 GND.n1373 19.3944
R18218 GND.n6242 GND.n1373 19.3944
R18219 GND.n6242 GND.n6241 19.3944
R18220 GND.n6241 GND.n6240 19.3944
R18221 GND.n6240 GND.n1381 19.3944
R18222 GND.n6234 GND.n1381 19.3944
R18223 GND.n6234 GND.n6233 19.3944
R18224 GND.n6233 GND.n6232 19.3944
R18225 GND.n6232 GND.n1389 19.3944
R18226 GND.n6226 GND.n1389 19.3944
R18227 GND.n6226 GND.n6225 19.3944
R18228 GND.n6225 GND.n6224 19.3944
R18229 GND.n6224 GND.n1397 19.3944
R18230 GND.n6218 GND.n1397 19.3944
R18231 GND.n6218 GND.n6217 19.3944
R18232 GND.n6217 GND.n6216 19.3944
R18233 GND.n6216 GND.n1405 19.3944
R18234 GND.n6210 GND.n1405 19.3944
R18235 GND.n6210 GND.n6209 19.3944
R18236 GND.n6209 GND.n6208 19.3944
R18237 GND.n6208 GND.n1413 19.3944
R18238 GND.n6202 GND.n1413 19.3944
R18239 GND.n6202 GND.n6201 19.3944
R18240 GND.n6201 GND.n6200 19.3944
R18241 GND.n6200 GND.n1421 19.3944
R18242 GND.n6194 GND.n1421 19.3944
R18243 GND.n6194 GND.n6193 19.3944
R18244 GND.n6193 GND.n6192 19.3944
R18245 GND.n6192 GND.n1429 19.3944
R18246 GND.n6186 GND.n1429 19.3944
R18247 GND.n6186 GND.n6185 19.3944
R18248 GND.n6185 GND.n6184 19.3944
R18249 GND.n6184 GND.n1437 19.3944
R18250 GND.n6178 GND.n1437 19.3944
R18251 GND.n6178 GND.n6177 19.3944
R18252 GND.n6177 GND.n6176 19.3944
R18253 GND.n6002 GND.n6001 19.3944
R18254 GND.n6001 GND.n1651 19.3944
R18255 GND.n5997 GND.n1651 19.3944
R18256 GND.n5997 GND.n5996 19.3944
R18257 GND.n5996 GND.n5995 19.3944
R18258 GND.n5995 GND.n1657 19.3944
R18259 GND.n5991 GND.n1657 19.3944
R18260 GND.n5991 GND.n5990 19.3944
R18261 GND.n5990 GND.n5989 19.3944
R18262 GND.n5983 GND.n5982 19.3944
R18263 GND.n5982 GND.n5981 19.3944
R18264 GND.n5981 GND.n1671 19.3944
R18265 GND.n5977 GND.n1671 19.3944
R18266 GND.n5977 GND.n5976 19.3944
R18267 GND.n5976 GND.n5975 19.3944
R18268 GND.n5975 GND.n1676 19.3944
R18269 GND.n5971 GND.n1676 19.3944
R18270 GND.n5971 GND.n5970 19.3944
R18271 GND.n5970 GND.n5969 19.3944
R18272 GND.n5969 GND.n1681 19.3944
R18273 GND.n5965 GND.n1681 19.3944
R18274 GND.n5965 GND.n5964 19.3944
R18275 GND.n5964 GND.n5963 19.3944
R18276 GND.n5963 GND.n1686 19.3944
R18277 GND.n5959 GND.n1686 19.3944
R18278 GND.n5959 GND.n5958 19.3944
R18279 GND.n5958 GND.n5957 19.3944
R18280 GND.n5957 GND.n1691 19.3944
R18281 GND.n5953 GND.n1691 19.3944
R18282 GND.n5953 GND.n5952 19.3944
R18283 GND.n5952 GND.n5951 19.3944
R18284 GND.n5951 GND.n1696 19.3944
R18285 GND.n5947 GND.n1696 19.3944
R18286 GND.n5947 GND.n5946 19.3944
R18287 GND.n5946 GND.n5945 19.3944
R18288 GND.n5945 GND.n1701 19.3944
R18289 GND.n5941 GND.n1701 19.3944
R18290 GND.n5941 GND.n5940 19.3944
R18291 GND.n5940 GND.n5939 19.3944
R18292 GND.n5939 GND.n1706 19.3944
R18293 GND.n5935 GND.n1706 19.3944
R18294 GND.n5935 GND.n5934 19.3944
R18295 GND.n5934 GND.n5933 19.3944
R18296 GND.n5933 GND.n1712 19.3944
R18297 GND.n5929 GND.n1712 19.3944
R18298 GND.n5929 GND.n5928 19.3944
R18299 GND.n5928 GND.n5927 19.3944
R18300 GND.n5927 GND.n1717 19.3944
R18301 GND.n5923 GND.n1717 19.3944
R18302 GND.n5923 GND.n5922 19.3944
R18303 GND.n5922 GND.n5921 19.3944
R18304 GND.n5921 GND.n1722 19.3944
R18305 GND.n5917 GND.n1722 19.3944
R18306 GND.n5917 GND.n5916 19.3944
R18307 GND.n5916 GND.n5915 19.3944
R18308 GND.n5915 GND.n1727 19.3944
R18309 GND.n5911 GND.n1727 19.3944
R18310 GND.n5911 GND.n5910 19.3944
R18311 GND.n5910 GND.n5909 19.3944
R18312 GND.n5909 GND.n1732 19.3944
R18313 GND.n5905 GND.n1732 19.3944
R18314 GND.n5905 GND.n5904 19.3944
R18315 GND.n5904 GND.n5903 19.3944
R18316 GND.n5903 GND.n1737 19.3944
R18317 GND.n5899 GND.n1737 19.3944
R18318 GND.n5899 GND.n5898 19.3944
R18319 GND.n5898 GND.n5897 19.3944
R18320 GND.n5897 GND.n1742 19.3944
R18321 GND.n4193 GND.n1747 19.2005
R18322 GND.n5148 GND.n5114 19.2005
R18323 GND.n2931 GND.n2930 19.2005
R18324 GND.n5989 GND.n1666 19.2005
R18325 GND.n5808 GND.n5807 18.8883
R18326 GND.n2497 GND.n2496 18.8883
R18327 GND.n5852 GND.n1817 18.4247
R18328 GND.n5408 GND.n2549 18.4247
R18329 GND.n4256 GND.n1965 18.3982
R18330 GND.n5778 GND.n1972 18.3982
R18331 GND.n5772 GND.n1981 18.3982
R18332 GND.n5758 GND.n5757 18.3982
R18333 GND.n5751 GND.n2027 18.3982
R18334 GND.n5744 GND.n2036 18.3982
R18335 GND.n5744 GND.n2037 18.3982
R18336 GND.n5738 GND.n2052 18.3982
R18337 GND.n5730 GND.n2063 18.3982
R18338 GND.n5724 GND.n5723 18.3982
R18339 GND.n5717 GND.n2096 18.3982
R18340 GND.n4400 GND.n2104 18.3982
R18341 GND.n4442 GND.n3038 18.3982
R18342 GND.n4385 GND.n2122 18.3982
R18343 GND.n4460 GND.n3017 18.3982
R18344 GND.n4371 GND.n2134 18.3982
R18345 GND.n4371 GND.n2140 18.3982
R18346 GND.n4366 GND.n4365 18.3982
R18347 GND.n4354 GND.n2151 18.3982
R18348 GND.n4480 GND.n3001 18.3982
R18349 GND.n4514 GND.n2169 18.3982
R18350 GND.n5653 GND.n2177 18.3982
R18351 GND.n5647 GND.n5646 18.3982
R18352 GND.n5640 GND.n2196 18.3982
R18353 GND.n5632 GND.n2206 18.3982
R18354 GND.n5626 GND.n2220 18.3982
R18355 GND.n5626 GND.n2222 18.3982
R18356 GND.n2240 GND.n2229 18.3982
R18357 GND.n4595 GND.n4594 18.3982
R18358 GND.n4583 GND.n2253 18.3982
R18359 GND.n4622 GND.n2974 18.3982
R18360 GND.n5593 GND.n5592 18.3982
R18361 GND.n5586 GND.n2280 18.3982
R18362 GND.n5578 GND.n2291 18.3982
R18363 GND.n5572 GND.n5571 18.3982
R18364 GND.n4694 GND.n2321 18.3982
R18365 GND.n5565 GND.n2321 18.3982
R18366 GND.n4702 GND.n2330 18.3982
R18367 GND.n4738 GND.n4737 18.3982
R18368 GND.n4769 GND.n2941 18.3982
R18369 GND.n4792 GND.n2363 18.3982
R18370 GND.n5477 GND.n2415 18.3982
R18371 GND.n3938 GND.t0 18.0303
R18372 GND.n5046 GND.t4 18.0303
R18373 GND.n5779 GND.n1969 17.6623
R18374 GND.n4408 GND.n4407 17.6623
R18375 GND.n5710 GND.n5709 17.6623
R18376 GND.n5661 GND.n5660 17.6623
R18377 GND.n2996 GND.n2995 17.6623
R18378 GND.n5599 GND.n2261 17.6623
R18379 GND.n2968 GND.n2271 17.6623
R18380 GND.n2945 GND.n2942 17.6623
R18381 GND.n4791 GND.n4790 17.6623
R18382 GND.n4321 GND.n4320 16.9264
R18383 GND.n5737 GND.n2054 16.9264
R18384 GND.n4380 GND.n4377 16.9264
R18385 GND.n2239 GND.n2236 16.9264
R18386 GND.n4685 GND.n2305 16.9264
R18387 GND.n5558 GND.n5557 16.9264
R18388 GND.n3669 GND.n3491 16.1905
R18389 GND.n3668 GND.n3475 16.1905
R18390 GND.n3680 GND.n3679 16.1905
R18391 GND.n3477 GND.n3468 16.1905
R18392 GND.n3691 GND.n3690 16.1905
R18393 GND.n3706 GND.n3456 16.1905
R18394 GND.n3458 GND.n3445 16.1905
R18395 GND.n3717 GND.n3716 16.1905
R18396 GND.n3448 GND.n3438 16.1905
R18397 GND.n3728 GND.n3727 16.1905
R18398 GND.n3743 GND.n3427 16.1905
R18399 GND.n3429 GND.n3417 16.1905
R18400 GND.n3754 GND.n3753 16.1905
R18401 GND.n3419 GND.n3409 16.1905
R18402 GND.n3765 GND.n3764 16.1905
R18403 GND.n3780 GND.n3397 16.1905
R18404 GND.n3400 GND.n3387 16.1905
R18405 GND.n3791 GND.n3790 16.1905
R18406 GND.n3389 GND.n3380 16.1905
R18407 GND.n3809 GND.n3807 16.1905
R18408 GND.n3817 GND.n3367 16.1905
R18409 GND.n3371 GND.n3369 16.1905
R18410 GND.n3826 GND.n3361 16.1905
R18411 GND.n3830 GND.n3358 16.1905
R18412 GND.n3938 GND.n3937 16.1905
R18413 GND.n3836 GND.n3337 16.1905
R18414 GND.n3930 GND.n3345 16.1905
R18415 GND.n3869 GND.n3347 16.1905
R18416 GND.n3879 GND.n3877 16.1905
R18417 GND.n3888 GND.n3865 16.1905
R18418 GND.n3889 GND.n3863 16.1905
R18419 GND.n3902 GND.n3900 16.1905
R18420 GND.n3905 GND.n3857 16.1905
R18421 GND.n3860 GND.n3859 16.1905
R18422 GND.n3912 GND.n3853 16.1905
R18423 GND.n3948 GND.n3321 16.1905
R18424 GND.n3312 GND.n3301 16.1905
R18425 GND.n3974 GND.n3973 16.1905
R18426 GND.n3303 GND.n3294 16.1905
R18427 GND.n3985 GND.n3984 16.1905
R18428 GND.n4000 GND.n3282 16.1905
R18429 GND.n3284 GND.n3271 16.1905
R18430 GND.n4011 GND.n4010 16.1905
R18431 GND.n3274 GND.n3264 16.1905
R18432 GND.n4022 GND.n4021 16.1905
R18433 GND.n4037 GND.n3253 16.1905
R18434 GND.n3255 GND.n3243 16.1905
R18435 GND.n4048 GND.n4047 16.1905
R18436 GND.n3245 GND.n3235 16.1905
R18437 GND.n4059 GND.n4058 16.1905
R18438 GND.n4074 GND.n3223 16.1905
R18439 GND.n4085 GND.n4084 16.1905
R18440 GND.n3215 GND.n3206 16.1905
R18441 GND.n4130 GND.n4128 16.1905
R18442 GND.n4140 GND.n3196 16.1905
R18443 GND.n4133 GND.n3198 16.1905
R18444 GND.n4149 GND.n3190 16.1905
R18445 GND.n4223 GND.n3186 16.1905
R18446 GND.n3080 GND.n1904 16.1905
R18447 GND.n3070 GND.n3063 16.1905
R18448 GND.n3050 GND.n2080 16.1905
R18449 GND.n5703 GND.n2114 16.1905
R18450 GND.n5667 GND.n2159 16.1905
R18451 GND.n2989 GND.n2187 16.1905
R18452 GND.n5607 GND.n5606 16.1905
R18453 GND.n5585 GND.n2283 16.1905
R18454 GND.n4753 GND.n2344 16.1905
R18455 GND.n4909 GND.n2594 16.1905
R18456 GND.n5332 GND.n2597 16.1905
R18457 GND.n5325 GND.n5324 16.1905
R18458 GND.n2617 GND.n2608 16.1905
R18459 GND.n5318 GND.n2618 16.1905
R18460 GND.n5317 GND.n2621 16.1905
R18461 GND.n4935 GND.n2636 16.1905
R18462 GND.n4943 GND.n2647 16.1905
R18463 GND.n5305 GND.n2650 16.1905
R18464 GND.n4950 GND.n2658 16.1905
R18465 GND.n5299 GND.n2661 16.1905
R18466 GND.n4958 GND.n2668 16.1905
R18467 GND.n5293 GND.n2671 16.1905
R18468 GND.n4965 GND.n2679 16.1905
R18469 GND.n5287 GND.n2682 16.1905
R18470 GND.n4973 GND.n2689 16.1905
R18471 GND.n5281 GND.n2692 16.1905
R18472 GND.n4980 GND.n2700 16.1905
R18473 GND.n5275 GND.n2703 16.1905
R18474 GND.n4988 GND.n2710 16.1905
R18475 GND.n5269 GND.n2713 16.1905
R18476 GND.n4995 GND.n2721 16.1905
R18477 GND.n5013 GND.n2730 16.1905
R18478 GND.n5257 GND.n2733 16.1905
R18479 GND.n5253 GND.n5252 16.1905
R18480 GND.n2744 GND.n2738 16.1905
R18481 GND.n5245 GND.n2747 16.1905
R18482 GND.n5244 GND.n28 16.1905
R18483 GND.n7824 GND.n30 16.1905
R18484 GND.n5238 GND.n5237 16.1905
R18485 GND.n5033 GND.n2759 16.1905
R18486 GND.n5040 GND.n47 16.1905
R18487 GND.n7817 GND.n50 16.1905
R18488 GND.n5047 GND.n5046 16.1905
R18489 GND.n7811 GND.n61 16.1905
R18490 GND.n5055 GND.n68 16.1905
R18491 GND.n7805 GND.n71 16.1905
R18492 GND.n5061 GND.n78 16.1905
R18493 GND.n7799 GND.n81 16.1905
R18494 GND.n5069 GND.n89 16.1905
R18495 GND.n7793 GND.n92 16.1905
R18496 GND.n5075 GND.n99 16.1905
R18497 GND.n7787 GND.n102 16.1905
R18498 GND.n5083 GND.n110 16.1905
R18499 GND.n7781 GND.n113 16.1905
R18500 GND.n5089 GND.n120 16.1905
R18501 GND.n7775 GND.n123 16.1905
R18502 GND.n5098 GND.n131 16.1905
R18503 GND.n7769 GND.n134 16.1905
R18504 GND.n5180 GND.n5179 16.1905
R18505 GND.n7763 GND.n143 16.1905
R18506 GND.n5173 GND.n151 16.1905
R18507 GND.n7757 GND.n154 16.1905
R18508 GND.n5167 GND.n161 16.1905
R18509 GND.n7751 GND.n164 16.1905
R18510 GND.n5161 GND.n172 16.1905
R18511 GND.n7745 GND.n175 16.1905
R18512 GND.n7738 GND.n7737 16.1905
R18513 GND.n1876 GND.n1853 16.0672
R18514 GND.n1866 GND.n1855 16.0672
R18515 GND.n2475 GND.n2474 16.0672
R18516 GND.n2481 GND.n2468 16.0672
R18517 GND.n3153 GND.n3118 15.7096
R18518 GND.n4870 GND.n4865 15.7096
R18519 GND.n303 GND.n302 15.7096
R18520 GND.n3617 GND.n3501 15.7096
R18521 GND.n5844 GND.n5808 15.6103
R18522 GND.n5448 GND.n2497 15.6103
R18523 GND.n4297 GND.n2016 15.4546
R18524 GND.n4417 GND.n3048 15.4546
R18525 GND.n4386 GND.n2116 15.4546
R18526 GND.n4355 GND.n2157 15.4546
R18527 GND.n4545 GND.n4544 15.4546
R18528 GND.n4629 GND.n4593 15.4546
R18529 GND.n5579 GND.n2289 15.4546
R18530 GND.n5551 GND.n2341 15.4546
R18531 GND.n2473 GND.n2472 15.4533
R18532 GND.n3057 GND.n2018 14.7187
R18533 GND.n5731 GND.n2060 14.7187
R18534 GND.n5696 GND.n5695 14.7187
R18535 GND.n5675 GND.n5674 14.7187
R18536 GND.n5639 GND.n2199 14.7187
R18537 GND.n5613 GND.n2238 14.7187
R18538 GND.n4663 GND.n2961 14.7187
R18539 GND.n4714 GND.n4713 14.7187
R18540 GND.n2427 GND.n2426 14.7187
R18541 GND.n1863 GND.n1856 14.2723
R18542 GND.n2491 GND.n2490 14.2723
R18543 GND.n3184 GND.n3183 14.1581
R18544 GND.n4906 GND.n4828 14.1581
R18545 GND.n275 GND.n270 14.1581
R18546 GND.n3652 GND.n3651 14.1581
R18547 GND.n5765 GND.n1989 13.9828
R18548 GND.n4395 GND.n4392 13.9828
R18549 GND.n4509 GND.n4506 13.9828
R18550 GND.n4534 GND.n2185 13.9828
R18551 GND.n4584 GND.n2259 13.9828
R18552 GND.n5544 GND.n5543 13.9828
R18553 GND.n5529 GND.n2371 13.9828
R18554 GND.t76 GND.n2433 13.9828
R18555 GND.n3716 GND.t52 13.6148
R18556 GND.n3947 GND.t8 13.6148
R18557 GND.t56 GND.n3213 13.6148
R18558 GND.n3069 GND.t63 13.6148
R18559 GND.n4752 GND.t97 13.6148
R18560 GND.n5311 GND.t38 13.6148
R18561 GND.n2815 GND.t2 13.6148
R18562 GND.n7763 GND.t34 13.6148
R18563 GND.n5803 GND.n1885 13.2469
R18564 GND.n5750 GND.n2030 13.2469
R18565 GND.n4333 GND.n4332 13.2469
R18566 GND.n5689 GND.n2132 13.2469
R18567 GND.n5620 GND.n2228 13.2469
R18568 GND.n2957 GND.n2307 13.2469
R18569 GND.n4703 GND.n2324 13.2469
R18570 GND.n5458 GND.n5457 13.2469
R18571 GND.n1880 GND.n1851 13.1884
R18572 GND.n1875 GND.n1874 13.1884
R18573 GND.n1874 GND.n1873 13.1884
R18574 GND.n1869 GND.n1868 13.1884
R18575 GND.n1868 GND.n1867 13.1884
R18576 GND.n2476 GND.n2471 13.1884
R18577 GND.n2477 GND.n2476 13.1884
R18578 GND.n2482 GND.n2469 13.1884
R18579 GND.n2483 GND.n2482 13.1884
R18580 GND.n4272 GND.n3076 12.511
R18581 GND.n5716 GND.n2098 12.511
R18582 GND.n4401 GND.n2098 12.511
R18583 GND.n4515 GND.n2175 12.511
R18584 GND.n5654 GND.n2175 12.511
R18585 GND.n4649 GND.n4640 12.511
R18586 GND.n4640 GND.n2269 12.511
R18587 GND.n5537 GND.n5536 12.511
R18588 GND.n3183 GND.n3104 11.8308
R18589 GND.n4900 GND.n4828 11.8308
R18590 GND.n278 GND.n275 11.8308
R18591 GND.n3651 GND.n3647 11.8308
R18592 GND.n5804 GND.n5803 11.775
R18593 GND.n4325 GND.n2030 11.775
R18594 GND.n4332 GND.n4331 11.775
R18595 GND.n5689 GND.n5688 11.775
R18596 GND.n5682 GND.n5681 11.775
R18597 GND.n4553 GND.n4552 11.775
R18598 GND.n2230 GND.n2228 11.775
R18599 GND.n4693 GND.n2957 11.775
R18600 GND.n5564 GND.n2324 11.775
R18601 GND.n5457 GND.n2433 11.775
R18602 GND.t67 GND.n5796 11.0391
R18603 GND.n5796 GND.n1896 11.0391
R18604 GND.n1902 GND.n1896 11.0391
R18605 GND.n5785 GND.t88 11.0391
R18606 GND.n4259 GND.n4258 11.0391
R18607 GND.n4273 GND.t42 11.0391
R18608 GND.n4278 GND.n1989 11.0391
R18609 GND.n4409 GND.n3053 11.0391
R18610 GND.n4392 GND.n2106 11.0391
R18611 GND.n4506 GND.n2167 11.0391
R18612 GND.n4534 GND.n4533 11.0391
R18613 GND.n5600 GND.n2259 11.0391
R18614 GND.n4674 GND.n2969 11.0391
R18615 GND.n5543 GND.n2353 11.0391
R18616 GND.n5530 GND.n5529 11.0391
R18617 GND.n5521 GND.n2378 11.0391
R18618 GND.n2443 GND.t76 11.0391
R18619 GND.n2547 GND.n2545 10.6151
R18620 GND.n2545 GND.n2542 10.6151
R18621 GND.n2542 GND.n2541 10.6151
R18622 GND.n2538 GND.n2537 10.6151
R18623 GND.n2537 GND.n2534 10.6151
R18624 GND.n2534 GND.n2533 10.6151
R18625 GND.n2533 GND.n2530 10.6151
R18626 GND.n2530 GND.n2529 10.6151
R18627 GND.n2529 GND.n2526 10.6151
R18628 GND.n2526 GND.n2525 10.6151
R18629 GND.n2525 GND.n2522 10.6151
R18630 GND.n2522 GND.n2521 10.6151
R18631 GND.n2521 GND.n2518 10.6151
R18632 GND.n2518 GND.n2517 10.6151
R18633 GND.n2517 GND.n2514 10.6151
R18634 GND.n2514 GND.n2513 10.6151
R18635 GND.n2513 GND.n2510 10.6151
R18636 GND.n2510 GND.n2509 10.6151
R18637 GND.n1951 GND.n1950 10.6151
R18638 GND.n1952 GND.n1951 10.6151
R18639 GND.n1952 GND.n1907 10.6151
R18640 GND.n1960 GND.n1907 10.6151
R18641 GND.n1961 GND.n1960 10.6151
R18642 GND.n1962 GND.n1961 10.6151
R18643 GND.n5789 GND.n1962 10.6151
R18644 GND.n5789 GND.n5788 10.6151
R18645 GND.n5788 GND.n5787 10.6151
R18646 GND.n5787 GND.n1963 10.6151
R18647 GND.n3073 GND.n1963 10.6151
R18648 GND.n3074 GND.n3073 10.6151
R18649 GND.n4275 GND.n3074 10.6151
R18650 GND.n4276 GND.n4275 10.6151
R18651 GND.n4280 GND.n4276 10.6151
R18652 GND.n4281 GND.n4280 10.6151
R18653 GND.n4282 GND.n4281 10.6151
R18654 GND.n4286 GND.n4282 10.6151
R18655 GND.n4286 GND.n4285 10.6151
R18656 GND.n4285 GND.n4284 10.6151
R18657 GND.n4284 GND.n3055 10.6151
R18658 GND.n4323 GND.n3055 10.6151
R18659 GND.n4324 GND.n4323 10.6151
R18660 GND.n4327 GND.n4324 10.6151
R18661 GND.n4328 GND.n4327 10.6151
R18662 GND.n4329 GND.n4328 10.6151
R18663 GND.n4335 GND.n4329 10.6151
R18664 GND.n4336 GND.n4335 10.6151
R18665 GND.n4339 GND.n4336 10.6151
R18666 GND.n4340 GND.n4339 10.6151
R18667 GND.n4342 GND.n4340 10.6151
R18668 GND.n4343 GND.n4342 10.6151
R18669 GND.n4344 GND.n4343 10.6151
R18670 GND.n4347 GND.n4344 10.6151
R18671 GND.n4348 GND.n4347 10.6151
R18672 GND.n4405 GND.n4348 10.6151
R18673 GND.n4405 GND.n4404 10.6151
R18674 GND.n4404 GND.n4403 10.6151
R18675 GND.n4403 GND.n4399 10.6151
R18676 GND.n4399 GND.n4398 10.6151
R18677 GND.n4398 GND.n4349 10.6151
R18678 GND.n4390 GND.n4349 10.6151
R18679 GND.n4390 GND.n4389 10.6151
R18680 GND.n4389 GND.n4388 10.6151
R18681 GND.n4388 GND.n4384 10.6151
R18682 GND.n4384 GND.n4383 10.6151
R18683 GND.n4383 GND.n4350 10.6151
R18684 GND.n4375 GND.n4350 10.6151
R18685 GND.n4375 GND.n4374 10.6151
R18686 GND.n4374 GND.n4373 10.6151
R18687 GND.n4373 GND.n4370 10.6151
R18688 GND.n4370 GND.n4369 10.6151
R18689 GND.n4369 GND.n4351 10.6151
R18690 GND.n4359 GND.n4351 10.6151
R18691 GND.n4359 GND.n4358 10.6151
R18692 GND.n4358 GND.n4357 10.6151
R18693 GND.n4357 GND.n4353 10.6151
R18694 GND.n4353 GND.n4352 10.6151
R18695 GND.n4352 GND.n2999 10.6151
R18696 GND.n4512 GND.n2999 10.6151
R18697 GND.n4513 GND.n4512 10.6151
R18698 GND.n4517 GND.n4513 10.6151
R18699 GND.n4518 GND.n4517 10.6151
R18700 GND.n4519 GND.n4518 10.6151
R18701 GND.n4523 GND.n4519 10.6151
R18702 GND.n4523 GND.n4522 10.6151
R18703 GND.n4522 GND.n4521 10.6151
R18704 GND.n4521 GND.n2987 10.6151
R18705 GND.n4547 GND.n2987 10.6151
R18706 GND.n4548 GND.n4547 10.6151
R18707 GND.n4558 GND.n4548 10.6151
R18708 GND.n4558 GND.n4557 10.6151
R18709 GND.n4557 GND.n4556 10.6151
R18710 GND.n4556 GND.n2225 10.6151
R18711 GND.n5624 GND.n2225 10.6151
R18712 GND.n5624 GND.n5623 10.6151
R18713 GND.n5623 GND.n5622 10.6151
R18714 GND.n5622 GND.n2226 10.6151
R18715 GND.n4579 GND.n2226 10.6151
R18716 GND.n4580 GND.n4579 10.6151
R18717 GND.n4589 GND.n4580 10.6151
R18718 GND.n4589 GND.n4588 10.6151
R18719 GND.n4588 GND.n4587 10.6151
R18720 GND.n4587 GND.n4586 10.6151
R18721 GND.n4586 GND.n4582 10.6151
R18722 GND.n4582 GND.n4581 10.6151
R18723 GND.n4581 GND.n2973 10.6151
R18724 GND.n2973 GND.n2971 10.6151
R18725 GND.n4653 GND.n2971 10.6151
R18726 GND.n4654 GND.n4653 10.6151
R18727 GND.n4671 GND.n4654 10.6151
R18728 GND.n4671 GND.n4670 10.6151
R18729 GND.n4670 GND.n4669 10.6151
R18730 GND.n4669 GND.n4666 10.6151
R18731 GND.n4666 GND.n4665 10.6151
R18732 GND.n4665 GND.n4662 10.6151
R18733 GND.n4662 GND.n4661 10.6151
R18734 GND.n4661 GND.n4658 10.6151
R18735 GND.n4658 GND.n4657 10.6151
R18736 GND.n4657 GND.n4656 10.6151
R18737 GND.n4656 GND.n2953 10.6151
R18738 GND.n4705 GND.n2953 10.6151
R18739 GND.n4706 GND.n4705 10.6151
R18740 GND.n4707 GND.n4706 10.6151
R18741 GND.n4709 GND.n4707 10.6151
R18742 GND.n4709 GND.n4708 10.6151
R18743 GND.n4708 GND.n2947 10.6151
R18744 GND.n4755 GND.n2947 10.6151
R18745 GND.n4756 GND.n4755 10.6151
R18746 GND.n4758 GND.n4756 10.6151
R18747 GND.n4759 GND.n4758 10.6151
R18748 GND.n4766 GND.n4759 10.6151
R18749 GND.n4766 GND.n4765 10.6151
R18750 GND.n4765 GND.n4764 10.6151
R18751 GND.n4764 GND.n4763 10.6151
R18752 GND.n4763 GND.n4762 10.6151
R18753 GND.n4762 GND.n4760 10.6151
R18754 GND.n4760 GND.n2423 10.6151
R18755 GND.n5468 GND.n2423 10.6151
R18756 GND.n5468 GND.n5467 10.6151
R18757 GND.n5467 GND.n5466 10.6151
R18758 GND.n5466 GND.n2424 10.6151
R18759 GND.n2504 GND.n2424 10.6151
R18760 GND.n2505 GND.n2504 10.6151
R18761 GND.n2505 GND.n2503 10.6151
R18762 GND.n1912 GND.n1823 10.6151
R18763 GND.n1913 GND.n1912 10.6151
R18764 GND.n1916 GND.n1913 10.6151
R18765 GND.n1921 GND.n1918 10.6151
R18766 GND.n1922 GND.n1921 10.6151
R18767 GND.n1925 GND.n1922 10.6151
R18768 GND.n1926 GND.n1925 10.6151
R18769 GND.n1929 GND.n1926 10.6151
R18770 GND.n1930 GND.n1929 10.6151
R18771 GND.n1933 GND.n1930 10.6151
R18772 GND.n1934 GND.n1933 10.6151
R18773 GND.n1937 GND.n1934 10.6151
R18774 GND.n1938 GND.n1937 10.6151
R18775 GND.n1941 GND.n1938 10.6151
R18776 GND.n1942 GND.n1941 10.6151
R18777 GND.n1945 GND.n1942 10.6151
R18778 GND.n1947 GND.n1945 10.6151
R18779 GND.n1948 GND.n1947 10.6151
R18780 GND.n5844 GND.n5843 10.6151
R18781 GND.n5843 GND.n5842 10.6151
R18782 GND.n5842 GND.n5841 10.6151
R18783 GND.n5841 GND.n5839 10.6151
R18784 GND.n5839 GND.n5836 10.6151
R18785 GND.n5836 GND.n5835 10.6151
R18786 GND.n5835 GND.n5832 10.6151
R18787 GND.n5832 GND.n5831 10.6151
R18788 GND.n5831 GND.n5828 10.6151
R18789 GND.n5828 GND.n5827 10.6151
R18790 GND.n5827 GND.n5824 10.6151
R18791 GND.n5824 GND.n5823 10.6151
R18792 GND.n5823 GND.n5820 10.6151
R18793 GND.n5820 GND.n5819 10.6151
R18794 GND.n5819 GND.n5816 10.6151
R18795 GND.n5814 GND.n5811 10.6151
R18796 GND.n5811 GND.n1825 10.6151
R18797 GND.n5850 GND.n1825 10.6151
R18798 GND.n5448 GND.n5447 10.6151
R18799 GND.n5447 GND.n5446 10.6151
R18800 GND.n5446 GND.n5443 10.6151
R18801 GND.n5443 GND.n5442 10.6151
R18802 GND.n5442 GND.n5439 10.6151
R18803 GND.n5439 GND.n5438 10.6151
R18804 GND.n5438 GND.n5435 10.6151
R18805 GND.n5435 GND.n5434 10.6151
R18806 GND.n5434 GND.n5431 10.6151
R18807 GND.n5431 GND.n5430 10.6151
R18808 GND.n5430 GND.n5427 10.6151
R18809 GND.n5427 GND.n5426 10.6151
R18810 GND.n5426 GND.n5423 10.6151
R18811 GND.n5423 GND.n5422 10.6151
R18812 GND.n5422 GND.n5419 10.6151
R18813 GND.n5417 GND.n5414 10.6151
R18814 GND.n5414 GND.n5413 10.6151
R18815 GND.n5413 GND.n5410 10.6151
R18816 GND.n5807 GND.n5806 10.6151
R18817 GND.n5806 GND.n1881 10.6151
R18818 GND.n1955 GND.n1881 10.6151
R18819 GND.n1955 GND.n1899 10.6151
R18820 GND.n5794 GND.n1899 10.6151
R18821 GND.n5794 GND.n5793 10.6151
R18822 GND.n5793 GND.n5792 10.6151
R18823 GND.n5792 GND.n1900 10.6151
R18824 GND.n5783 GND.n1900 10.6151
R18825 GND.n5783 GND.n5782 10.6151
R18826 GND.n5782 GND.n5781 10.6151
R18827 GND.n5781 GND.n1967 10.6151
R18828 GND.n1986 GND.n1967 10.6151
R18829 GND.n5769 GND.n1986 10.6151
R18830 GND.n5769 GND.n5768 10.6151
R18831 GND.n5768 GND.n5767 10.6151
R18832 GND.n5767 GND.n1987 10.6151
R18833 GND.n4294 GND.n1987 10.6151
R18834 GND.n4294 GND.n4293 10.6151
R18835 GND.n4293 GND.n4292 10.6151
R18836 GND.n4292 GND.n4289 10.6151
R18837 GND.n4289 GND.n2033 10.6151
R18838 GND.n5748 GND.n2033 10.6151
R18839 GND.n5748 GND.n5747 10.6151
R18840 GND.n5747 GND.n5746 10.6151
R18841 GND.n5746 GND.n2034 10.6151
R18842 GND.n2057 GND.n2034 10.6151
R18843 GND.n5735 GND.n2057 10.6151
R18844 GND.n5735 GND.n5734 10.6151
R18845 GND.n5734 GND.n5733 10.6151
R18846 GND.n5733 GND.n2058 10.6151
R18847 GND.n4414 GND.n2058 10.6151
R18848 GND.n4414 GND.n4413 10.6151
R18849 GND.n4413 GND.n4412 10.6151
R18850 GND.n4412 GND.n3052 10.6151
R18851 GND.n3052 GND.n2101 10.6151
R18852 GND.n5714 GND.n2101 10.6151
R18853 GND.n5714 GND.n5713 10.6151
R18854 GND.n5713 GND.n5712 10.6151
R18855 GND.n5712 GND.n2102 10.6151
R18856 GND.n4393 GND.n2102 10.6151
R18857 GND.n4393 GND.n2119 10.6151
R18858 GND.n5700 GND.n2119 10.6151
R18859 GND.n5700 GND.n5699 10.6151
R18860 GND.n5699 GND.n5698 10.6151
R18861 GND.n5698 GND.n2120 10.6151
R18862 GND.n4378 GND.n2120 10.6151
R18863 GND.n4378 GND.n2137 10.6151
R18864 GND.n5686 GND.n2137 10.6151
R18865 GND.n5686 GND.n5685 10.6151
R18866 GND.n5685 GND.n5684 10.6151
R18867 GND.n5684 GND.n2138 10.6151
R18868 GND.n4362 GND.n2138 10.6151
R18869 GND.n4362 GND.n2154 10.6151
R18870 GND.n5672 GND.n2154 10.6151
R18871 GND.n5672 GND.n5671 10.6151
R18872 GND.n5671 GND.n5670 10.6151
R18873 GND.n5670 GND.n2155 10.6151
R18874 GND.n4507 GND.n2155 10.6151
R18875 GND.n4507 GND.n2172 10.6151
R18876 GND.n5658 GND.n2172 10.6151
R18877 GND.n5658 GND.n5657 10.6151
R18878 GND.n5657 GND.n5656 10.6151
R18879 GND.n5656 GND.n2173 10.6151
R18880 GND.n4531 GND.n2173 10.6151
R18881 GND.n4531 GND.n4530 10.6151
R18882 GND.n4530 GND.n4529 10.6151
R18883 GND.n4529 GND.n4526 10.6151
R18884 GND.n4526 GND.n2202 10.6151
R18885 GND.n5637 GND.n2202 10.6151
R18886 GND.n5637 GND.n5636 10.6151
R18887 GND.n5636 GND.n5635 10.6151
R18888 GND.n5635 GND.n2203 10.6151
R18889 GND.n4550 GND.n2203 10.6151
R18890 GND.n4550 GND.n4549 10.6151
R18891 GND.n4549 GND.n2233 10.6151
R18892 GND.n5618 GND.n2233 10.6151
R18893 GND.n5618 GND.n5617 10.6151
R18894 GND.n5617 GND.n5616 10.6151
R18895 GND.n5616 GND.n2234 10.6151
R18896 GND.n4591 GND.n2234 10.6151
R18897 GND.n4591 GND.n2256 10.6151
R18898 GND.n5604 GND.n2256 10.6151
R18899 GND.n5604 GND.n5603 10.6151
R18900 GND.n5603 GND.n5602 10.6151
R18901 GND.n5602 GND.n2257 10.6151
R18902 GND.n4647 GND.n2257 10.6151
R18903 GND.n4647 GND.n4646 10.6151
R18904 GND.n4646 GND.n4645 10.6151
R18905 GND.n4645 GND.n4642 10.6151
R18906 GND.n4642 GND.n2286 10.6151
R18907 GND.n5583 GND.n2286 10.6151
R18908 GND.n5583 GND.n5582 10.6151
R18909 GND.n5582 GND.n5581 10.6151
R18910 GND.n5581 GND.n2287 10.6151
R18911 GND.n2960 GND.n2287 10.6151
R18912 GND.n4689 GND.n2960 10.6151
R18913 GND.n4690 GND.n4689 10.6151
R18914 GND.n4691 GND.n4690 10.6151
R18915 GND.n4691 GND.n2327 10.6151
R18916 GND.n5562 GND.n2327 10.6151
R18917 GND.n5562 GND.n5561 10.6151
R18918 GND.n5561 GND.n5560 10.6151
R18919 GND.n5560 GND.n2328 10.6151
R18920 GND.n4711 GND.n2328 10.6151
R18921 GND.n4711 GND.n2347 10.6151
R18922 GND.n5548 GND.n2347 10.6151
R18923 GND.n5548 GND.n5547 10.6151
R18924 GND.n5547 GND.n5546 10.6151
R18925 GND.n5546 GND.n2348 10.6151
R18926 GND.n2943 GND.n2348 10.6151
R18927 GND.n2943 GND.n2366 10.6151
R18928 GND.n5534 GND.n2366 10.6151
R18929 GND.n5534 GND.n5533 10.6151
R18930 GND.n5533 GND.n5532 10.6151
R18931 GND.n5532 GND.n2367 10.6151
R18932 GND.n5474 GND.n2367 10.6151
R18933 GND.n5474 GND.n5473 10.6151
R18934 GND.n5473 GND.n5472 10.6151
R18935 GND.n5472 GND.n2418 10.6151
R18936 GND.n5462 GND.n2418 10.6151
R18937 GND.n5462 GND.n5461 10.6151
R18938 GND.n5461 GND.n5460 10.6151
R18939 GND.n5460 GND.n2430 10.6151
R18940 GND.n2496 GND.n2430 10.6151
R18941 GND.n5797 GND.n1894 10.3032
R18942 GND.n3058 GND.n3057 10.3032
R18943 GND.n4337 GND.n2060 10.3032
R18944 GND.n5695 GND.n2124 10.3032
R18945 GND.n5675 GND.n2149 10.3032
R18946 GND.n4560 GND.n2199 10.3032
R18947 GND.n5614 GND.n5613 10.3032
R18948 GND.n4686 GND.n2961 10.3032
R18949 GND.n4714 GND.n2333 10.3032
R18950 GND.n4784 GND.t117 10.3032
R18951 GND.n5464 GND.n2427 10.3032
R18952 GND.n3157 GND.n3118 10.2793
R18953 GND.n4870 GND.n4834 10.2793
R18954 GND.n302 GND.n255 10.2793
R18955 GND.n3618 GND.n3617 10.2793
R18956 GND.n1872 GND.n1853 10.2247
R18957 GND.n1870 GND.n1855 10.2247
R18958 GND.n2475 GND.n2470 10.2247
R18959 GND.n2481 GND.n2480 10.2247
R18960 GND.n4277 GND.t60 9.56732
R18961 GND.n4297 GND.n4296 9.56732
R18962 GND.n4417 GND.n4416 9.56732
R18963 GND.n5702 GND.n2116 9.56732
R18964 GND.n5668 GND.n2157 9.56732
R18965 GND.n4544 GND.n2990 9.56732
R18966 GND.n4629 GND.n2251 9.56732
R18967 GND.n4667 GND.n2289 9.56732
R18968 GND.n5551 GND.n5550 9.56732
R18969 GND.n2538 GND.n2502 9.36635
R18970 GND.n1918 GND.n1917 9.36635
R18971 GND.n5816 GND.n5815 9.36635
R18972 GND.n5419 GND.n5418 9.36635
R18973 GND.n6356 GND.n6355 9.3005
R18974 GND.n1264 GND.n1263 9.3005
R18975 GND.n6363 GND.n6362 9.3005
R18976 GND.n6364 GND.n1262 9.3005
R18977 GND.n6366 GND.n6365 9.3005
R18978 GND.n1258 GND.n1257 9.3005
R18979 GND.n6373 GND.n6372 9.3005
R18980 GND.n6374 GND.n1256 9.3005
R18981 GND.n6376 GND.n6375 9.3005
R18982 GND.n1252 GND.n1251 9.3005
R18983 GND.n6383 GND.n6382 9.3005
R18984 GND.n6384 GND.n1250 9.3005
R18985 GND.n6386 GND.n6385 9.3005
R18986 GND.n1246 GND.n1245 9.3005
R18987 GND.n6393 GND.n6392 9.3005
R18988 GND.n6394 GND.n1244 9.3005
R18989 GND.n6396 GND.n6395 9.3005
R18990 GND.n1240 GND.n1239 9.3005
R18991 GND.n6403 GND.n6402 9.3005
R18992 GND.n6404 GND.n1238 9.3005
R18993 GND.n6406 GND.n6405 9.3005
R18994 GND.n1234 GND.n1233 9.3005
R18995 GND.n6413 GND.n6412 9.3005
R18996 GND.n6414 GND.n1232 9.3005
R18997 GND.n6416 GND.n6415 9.3005
R18998 GND.n1228 GND.n1227 9.3005
R18999 GND.n6423 GND.n6422 9.3005
R19000 GND.n6424 GND.n1226 9.3005
R19001 GND.n6426 GND.n6425 9.3005
R19002 GND.n1222 GND.n1221 9.3005
R19003 GND.n6433 GND.n6432 9.3005
R19004 GND.n6434 GND.n1220 9.3005
R19005 GND.n6436 GND.n6435 9.3005
R19006 GND.n1216 GND.n1215 9.3005
R19007 GND.n6443 GND.n6442 9.3005
R19008 GND.n6444 GND.n1214 9.3005
R19009 GND.n6446 GND.n6445 9.3005
R19010 GND.n1210 GND.n1209 9.3005
R19011 GND.n6453 GND.n6452 9.3005
R19012 GND.n6454 GND.n1208 9.3005
R19013 GND.n6456 GND.n6455 9.3005
R19014 GND.n1204 GND.n1203 9.3005
R19015 GND.n6463 GND.n6462 9.3005
R19016 GND.n6464 GND.n1202 9.3005
R19017 GND.n6466 GND.n6465 9.3005
R19018 GND.n1198 GND.n1197 9.3005
R19019 GND.n6473 GND.n6472 9.3005
R19020 GND.n6474 GND.n1196 9.3005
R19021 GND.n6476 GND.n6475 9.3005
R19022 GND.n1192 GND.n1191 9.3005
R19023 GND.n6483 GND.n6482 9.3005
R19024 GND.n6484 GND.n1190 9.3005
R19025 GND.n6486 GND.n6485 9.3005
R19026 GND.n1186 GND.n1185 9.3005
R19027 GND.n6493 GND.n6492 9.3005
R19028 GND.n6494 GND.n1184 9.3005
R19029 GND.n6496 GND.n6495 9.3005
R19030 GND.n1180 GND.n1179 9.3005
R19031 GND.n6503 GND.n6502 9.3005
R19032 GND.n6504 GND.n1178 9.3005
R19033 GND.n6506 GND.n6505 9.3005
R19034 GND.n1174 GND.n1173 9.3005
R19035 GND.n6513 GND.n6512 9.3005
R19036 GND.n6514 GND.n1172 9.3005
R19037 GND.n6516 GND.n6515 9.3005
R19038 GND.n1168 GND.n1167 9.3005
R19039 GND.n6523 GND.n6522 9.3005
R19040 GND.n6524 GND.n1166 9.3005
R19041 GND.n6526 GND.n6525 9.3005
R19042 GND.n1162 GND.n1161 9.3005
R19043 GND.n6533 GND.n6532 9.3005
R19044 GND.n6534 GND.n1160 9.3005
R19045 GND.n6536 GND.n6535 9.3005
R19046 GND.n1156 GND.n1155 9.3005
R19047 GND.n6543 GND.n6542 9.3005
R19048 GND.n6544 GND.n1154 9.3005
R19049 GND.n6546 GND.n6545 9.3005
R19050 GND.n1150 GND.n1149 9.3005
R19051 GND.n6553 GND.n6552 9.3005
R19052 GND.n6554 GND.n1148 9.3005
R19053 GND.n6556 GND.n6555 9.3005
R19054 GND.n1144 GND.n1143 9.3005
R19055 GND.n6563 GND.n6562 9.3005
R19056 GND.n6564 GND.n1142 9.3005
R19057 GND.n6566 GND.n6565 9.3005
R19058 GND.n1138 GND.n1137 9.3005
R19059 GND.n6573 GND.n6572 9.3005
R19060 GND.n6574 GND.n1136 9.3005
R19061 GND.n6576 GND.n6575 9.3005
R19062 GND.n1132 GND.n1131 9.3005
R19063 GND.n6583 GND.n6582 9.3005
R19064 GND.n6584 GND.n1130 9.3005
R19065 GND.n6586 GND.n6585 9.3005
R19066 GND.n1126 GND.n1125 9.3005
R19067 GND.n6593 GND.n6592 9.3005
R19068 GND.n6594 GND.n1124 9.3005
R19069 GND.n6596 GND.n6595 9.3005
R19070 GND.n1120 GND.n1119 9.3005
R19071 GND.n6603 GND.n6602 9.3005
R19072 GND.n6604 GND.n1118 9.3005
R19073 GND.n6606 GND.n6605 9.3005
R19074 GND.n1114 GND.n1113 9.3005
R19075 GND.n6613 GND.n6612 9.3005
R19076 GND.n6614 GND.n1112 9.3005
R19077 GND.n6616 GND.n6615 9.3005
R19078 GND.n1108 GND.n1107 9.3005
R19079 GND.n6623 GND.n6622 9.3005
R19080 GND.n6624 GND.n1106 9.3005
R19081 GND.n6626 GND.n6625 9.3005
R19082 GND.n1102 GND.n1101 9.3005
R19083 GND.n6633 GND.n6632 9.3005
R19084 GND.n6634 GND.n1100 9.3005
R19085 GND.n6636 GND.n6635 9.3005
R19086 GND.n1096 GND.n1095 9.3005
R19087 GND.n6643 GND.n6642 9.3005
R19088 GND.n6644 GND.n1094 9.3005
R19089 GND.n6646 GND.n6645 9.3005
R19090 GND.n1090 GND.n1089 9.3005
R19091 GND.n6653 GND.n6652 9.3005
R19092 GND.n6654 GND.n1088 9.3005
R19093 GND.n6656 GND.n6655 9.3005
R19094 GND.n1084 GND.n1083 9.3005
R19095 GND.n6663 GND.n6662 9.3005
R19096 GND.n6664 GND.n1082 9.3005
R19097 GND.n6666 GND.n6665 9.3005
R19098 GND.n1078 GND.n1077 9.3005
R19099 GND.n6673 GND.n6672 9.3005
R19100 GND.n6674 GND.n1076 9.3005
R19101 GND.n6676 GND.n6675 9.3005
R19102 GND.n1072 GND.n1071 9.3005
R19103 GND.n6683 GND.n6682 9.3005
R19104 GND.n6684 GND.n1070 9.3005
R19105 GND.n6686 GND.n6685 9.3005
R19106 GND.n1066 GND.n1065 9.3005
R19107 GND.n6693 GND.n6692 9.3005
R19108 GND.n6694 GND.n1064 9.3005
R19109 GND.n6696 GND.n6695 9.3005
R19110 GND.n1060 GND.n1059 9.3005
R19111 GND.n6703 GND.n6702 9.3005
R19112 GND.n6704 GND.n1058 9.3005
R19113 GND.n6706 GND.n6705 9.3005
R19114 GND.n1054 GND.n1053 9.3005
R19115 GND.n6713 GND.n6712 9.3005
R19116 GND.n6714 GND.n1052 9.3005
R19117 GND.n6716 GND.n6715 9.3005
R19118 GND.n1048 GND.n1047 9.3005
R19119 GND.n6723 GND.n6722 9.3005
R19120 GND.n6724 GND.n1046 9.3005
R19121 GND.n6726 GND.n6725 9.3005
R19122 GND.n1042 GND.n1041 9.3005
R19123 GND.n6733 GND.n6732 9.3005
R19124 GND.n6734 GND.n1040 9.3005
R19125 GND.n6736 GND.n6735 9.3005
R19126 GND.n1036 GND.n1035 9.3005
R19127 GND.n6743 GND.n6742 9.3005
R19128 GND.n6744 GND.n1034 9.3005
R19129 GND.n6746 GND.n6745 9.3005
R19130 GND.n1030 GND.n1029 9.3005
R19131 GND.n6753 GND.n6752 9.3005
R19132 GND.n6754 GND.n1028 9.3005
R19133 GND.n6756 GND.n6755 9.3005
R19134 GND.n1024 GND.n1023 9.3005
R19135 GND.n6763 GND.n6762 9.3005
R19136 GND.n6764 GND.n1022 9.3005
R19137 GND.n6766 GND.n6765 9.3005
R19138 GND.n1018 GND.n1017 9.3005
R19139 GND.n6773 GND.n6772 9.3005
R19140 GND.n6774 GND.n1016 9.3005
R19141 GND.n6776 GND.n6775 9.3005
R19142 GND.n1012 GND.n1011 9.3005
R19143 GND.n6783 GND.n6782 9.3005
R19144 GND.n6784 GND.n1010 9.3005
R19145 GND.n6786 GND.n6785 9.3005
R19146 GND.n1006 GND.n1005 9.3005
R19147 GND.n6793 GND.n6792 9.3005
R19148 GND.n6794 GND.n1004 9.3005
R19149 GND.n6796 GND.n6795 9.3005
R19150 GND.n1000 GND.n999 9.3005
R19151 GND.n6803 GND.n6802 9.3005
R19152 GND.n6804 GND.n998 9.3005
R19153 GND.n6806 GND.n6805 9.3005
R19154 GND.n994 GND.n993 9.3005
R19155 GND.n6813 GND.n6812 9.3005
R19156 GND.n6814 GND.n992 9.3005
R19157 GND.n6816 GND.n6815 9.3005
R19158 GND.n988 GND.n987 9.3005
R19159 GND.n6823 GND.n6822 9.3005
R19160 GND.n6824 GND.n986 9.3005
R19161 GND.n6826 GND.n6825 9.3005
R19162 GND.n982 GND.n981 9.3005
R19163 GND.n6833 GND.n6832 9.3005
R19164 GND.n6834 GND.n980 9.3005
R19165 GND.n6836 GND.n6835 9.3005
R19166 GND.n976 GND.n975 9.3005
R19167 GND.n6843 GND.n6842 9.3005
R19168 GND.n6844 GND.n974 9.3005
R19169 GND.n6846 GND.n6845 9.3005
R19170 GND.n970 GND.n969 9.3005
R19171 GND.n6853 GND.n6852 9.3005
R19172 GND.n6854 GND.n968 9.3005
R19173 GND.n6856 GND.n6855 9.3005
R19174 GND.n964 GND.n963 9.3005
R19175 GND.n6863 GND.n6862 9.3005
R19176 GND.n6864 GND.n962 9.3005
R19177 GND.n6866 GND.n6865 9.3005
R19178 GND.n958 GND.n957 9.3005
R19179 GND.n6873 GND.n6872 9.3005
R19180 GND.n6874 GND.n956 9.3005
R19181 GND.n6876 GND.n6875 9.3005
R19182 GND.n952 GND.n951 9.3005
R19183 GND.n6883 GND.n6882 9.3005
R19184 GND.n6884 GND.n950 9.3005
R19185 GND.n6886 GND.n6885 9.3005
R19186 GND.n946 GND.n945 9.3005
R19187 GND.n6893 GND.n6892 9.3005
R19188 GND.n6894 GND.n944 9.3005
R19189 GND.n6896 GND.n6895 9.3005
R19190 GND.n940 GND.n939 9.3005
R19191 GND.n6903 GND.n6902 9.3005
R19192 GND.n6904 GND.n938 9.3005
R19193 GND.n6906 GND.n6905 9.3005
R19194 GND.n934 GND.n933 9.3005
R19195 GND.n6913 GND.n6912 9.3005
R19196 GND.n6914 GND.n932 9.3005
R19197 GND.n6916 GND.n6915 9.3005
R19198 GND.n928 GND.n927 9.3005
R19199 GND.n6923 GND.n6922 9.3005
R19200 GND.n6924 GND.n926 9.3005
R19201 GND.n6926 GND.n6925 9.3005
R19202 GND.n922 GND.n921 9.3005
R19203 GND.n6933 GND.n6932 9.3005
R19204 GND.n6934 GND.n920 9.3005
R19205 GND.n6936 GND.n6935 9.3005
R19206 GND.n916 GND.n915 9.3005
R19207 GND.n6943 GND.n6942 9.3005
R19208 GND.n6944 GND.n914 9.3005
R19209 GND.n6946 GND.n6945 9.3005
R19210 GND.n910 GND.n909 9.3005
R19211 GND.n6953 GND.n6952 9.3005
R19212 GND.n6954 GND.n908 9.3005
R19213 GND.n6956 GND.n6955 9.3005
R19214 GND.n904 GND.n903 9.3005
R19215 GND.n6963 GND.n6962 9.3005
R19216 GND.n6964 GND.n902 9.3005
R19217 GND.n6966 GND.n6965 9.3005
R19218 GND.n898 GND.n897 9.3005
R19219 GND.n6973 GND.n6972 9.3005
R19220 GND.n6974 GND.n896 9.3005
R19221 GND.n6976 GND.n6975 9.3005
R19222 GND.n892 GND.n891 9.3005
R19223 GND.n6983 GND.n6982 9.3005
R19224 GND.n6984 GND.n890 9.3005
R19225 GND.n6986 GND.n6985 9.3005
R19226 GND.n886 GND.n885 9.3005
R19227 GND.n6993 GND.n6992 9.3005
R19228 GND.n6994 GND.n884 9.3005
R19229 GND.n6996 GND.n6995 9.3005
R19230 GND.n880 GND.n879 9.3005
R19231 GND.n7003 GND.n7002 9.3005
R19232 GND.n7004 GND.n878 9.3005
R19233 GND.n7006 GND.n7005 9.3005
R19234 GND.n874 GND.n873 9.3005
R19235 GND.n7013 GND.n7012 9.3005
R19236 GND.n7014 GND.n872 9.3005
R19237 GND.n7016 GND.n7015 9.3005
R19238 GND.n868 GND.n867 9.3005
R19239 GND.n7023 GND.n7022 9.3005
R19240 GND.n7024 GND.n866 9.3005
R19241 GND.n7026 GND.n7025 9.3005
R19242 GND.n862 GND.n861 9.3005
R19243 GND.n7033 GND.n7032 9.3005
R19244 GND.n7034 GND.n860 9.3005
R19245 GND.n7036 GND.n7035 9.3005
R19246 GND.n856 GND.n855 9.3005
R19247 GND.n7043 GND.n7042 9.3005
R19248 GND.n7044 GND.n854 9.3005
R19249 GND.n7046 GND.n7045 9.3005
R19250 GND.n850 GND.n849 9.3005
R19251 GND.n7053 GND.n7052 9.3005
R19252 GND.n7054 GND.n848 9.3005
R19253 GND.n7056 GND.n7055 9.3005
R19254 GND.n844 GND.n843 9.3005
R19255 GND.n7063 GND.n7062 9.3005
R19256 GND.n7064 GND.n842 9.3005
R19257 GND.n7066 GND.n7065 9.3005
R19258 GND.n838 GND.n837 9.3005
R19259 GND.n7073 GND.n7072 9.3005
R19260 GND.n7074 GND.n836 9.3005
R19261 GND.n7076 GND.n7075 9.3005
R19262 GND.n832 GND.n831 9.3005
R19263 GND.n7083 GND.n7082 9.3005
R19264 GND.n7084 GND.n830 9.3005
R19265 GND.n7086 GND.n7085 9.3005
R19266 GND.n826 GND.n825 9.3005
R19267 GND.n7093 GND.n7092 9.3005
R19268 GND.n7094 GND.n824 9.3005
R19269 GND.n7096 GND.n7095 9.3005
R19270 GND.n820 GND.n819 9.3005
R19271 GND.n7103 GND.n7102 9.3005
R19272 GND.n7104 GND.n818 9.3005
R19273 GND.n7106 GND.n7105 9.3005
R19274 GND.n814 GND.n813 9.3005
R19275 GND.n7113 GND.n7112 9.3005
R19276 GND.n7114 GND.n812 9.3005
R19277 GND.n7116 GND.n7115 9.3005
R19278 GND.n808 GND.n807 9.3005
R19279 GND.n7123 GND.n7122 9.3005
R19280 GND.n7124 GND.n806 9.3005
R19281 GND.n7126 GND.n7125 9.3005
R19282 GND.n802 GND.n801 9.3005
R19283 GND.n7133 GND.n7132 9.3005
R19284 GND.n7134 GND.n800 9.3005
R19285 GND.n7136 GND.n7135 9.3005
R19286 GND.n796 GND.n795 9.3005
R19287 GND.n7143 GND.n7142 9.3005
R19288 GND.n7144 GND.n794 9.3005
R19289 GND.n7146 GND.n7145 9.3005
R19290 GND.n790 GND.n789 9.3005
R19291 GND.n7153 GND.n7152 9.3005
R19292 GND.n7154 GND.n788 9.3005
R19293 GND.n7156 GND.n7155 9.3005
R19294 GND.n784 GND.n783 9.3005
R19295 GND.n7163 GND.n7162 9.3005
R19296 GND.n7164 GND.n782 9.3005
R19297 GND.n7166 GND.n7165 9.3005
R19298 GND.n778 GND.n777 9.3005
R19299 GND.n7173 GND.n7172 9.3005
R19300 GND.n7174 GND.n776 9.3005
R19301 GND.n7176 GND.n7175 9.3005
R19302 GND.n772 GND.n771 9.3005
R19303 GND.n7183 GND.n7182 9.3005
R19304 GND.n7184 GND.n770 9.3005
R19305 GND.n7186 GND.n7185 9.3005
R19306 GND.n766 GND.n765 9.3005
R19307 GND.n7193 GND.n7192 9.3005
R19308 GND.n7194 GND.n764 9.3005
R19309 GND.n7196 GND.n7195 9.3005
R19310 GND.n760 GND.n759 9.3005
R19311 GND.n7203 GND.n7202 9.3005
R19312 GND.n7204 GND.n758 9.3005
R19313 GND.n7206 GND.n7205 9.3005
R19314 GND.n754 GND.n753 9.3005
R19315 GND.n7213 GND.n7212 9.3005
R19316 GND.n7214 GND.n752 9.3005
R19317 GND.n7216 GND.n7215 9.3005
R19318 GND.n748 GND.n747 9.3005
R19319 GND.n7223 GND.n7222 9.3005
R19320 GND.n7224 GND.n746 9.3005
R19321 GND.n7226 GND.n7225 9.3005
R19322 GND.n742 GND.n741 9.3005
R19323 GND.n7233 GND.n7232 9.3005
R19324 GND.n7234 GND.n740 9.3005
R19325 GND.n7236 GND.n7235 9.3005
R19326 GND.n736 GND.n735 9.3005
R19327 GND.n7243 GND.n7242 9.3005
R19328 GND.n7244 GND.n734 9.3005
R19329 GND.n7246 GND.n7245 9.3005
R19330 GND.n730 GND.n729 9.3005
R19331 GND.n7253 GND.n7252 9.3005
R19332 GND.n7254 GND.n728 9.3005
R19333 GND.n7256 GND.n7255 9.3005
R19334 GND.n724 GND.n723 9.3005
R19335 GND.n7263 GND.n7262 9.3005
R19336 GND.n7264 GND.n722 9.3005
R19337 GND.n7266 GND.n7265 9.3005
R19338 GND.n718 GND.n717 9.3005
R19339 GND.n7273 GND.n7272 9.3005
R19340 GND.n7274 GND.n716 9.3005
R19341 GND.n7276 GND.n7275 9.3005
R19342 GND.n712 GND.n711 9.3005
R19343 GND.n7283 GND.n7282 9.3005
R19344 GND.n7284 GND.n710 9.3005
R19345 GND.n7286 GND.n7285 9.3005
R19346 GND.n706 GND.n705 9.3005
R19347 GND.n7293 GND.n7292 9.3005
R19348 GND.n7294 GND.n704 9.3005
R19349 GND.n7296 GND.n7295 9.3005
R19350 GND.n700 GND.n699 9.3005
R19351 GND.n7303 GND.n7302 9.3005
R19352 GND.n7304 GND.n698 9.3005
R19353 GND.n7306 GND.n7305 9.3005
R19354 GND.n694 GND.n693 9.3005
R19355 GND.n7313 GND.n7312 9.3005
R19356 GND.n7314 GND.n692 9.3005
R19357 GND.n7316 GND.n7315 9.3005
R19358 GND.n688 GND.n687 9.3005
R19359 GND.n7323 GND.n7322 9.3005
R19360 GND.n7324 GND.n686 9.3005
R19361 GND.n7327 GND.n7326 9.3005
R19362 GND.n7325 GND.n682 9.3005
R19363 GND.n7333 GND.n681 9.3005
R19364 GND.n7335 GND.n7334 9.3005
R19365 GND.n677 GND.n676 9.3005
R19366 GND.n7344 GND.n7343 9.3005
R19367 GND.n7345 GND.n675 9.3005
R19368 GND.n7347 GND.n7346 9.3005
R19369 GND.n671 GND.n670 9.3005
R19370 GND.n7354 GND.n7353 9.3005
R19371 GND.n7355 GND.n669 9.3005
R19372 GND.n7357 GND.n7356 9.3005
R19373 GND.n665 GND.n664 9.3005
R19374 GND.n7364 GND.n7363 9.3005
R19375 GND.n7365 GND.n663 9.3005
R19376 GND.n7367 GND.n7366 9.3005
R19377 GND.n659 GND.n658 9.3005
R19378 GND.n7374 GND.n7373 9.3005
R19379 GND.n7375 GND.n657 9.3005
R19380 GND.n7377 GND.n7376 9.3005
R19381 GND.n653 GND.n652 9.3005
R19382 GND.n7384 GND.n7383 9.3005
R19383 GND.n7385 GND.n651 9.3005
R19384 GND.n7387 GND.n7386 9.3005
R19385 GND.n647 GND.n646 9.3005
R19386 GND.n7394 GND.n7393 9.3005
R19387 GND.n7395 GND.n645 9.3005
R19388 GND.n7397 GND.n7396 9.3005
R19389 GND.n641 GND.n640 9.3005
R19390 GND.n7404 GND.n7403 9.3005
R19391 GND.n7405 GND.n639 9.3005
R19392 GND.n7407 GND.n7406 9.3005
R19393 GND.n635 GND.n634 9.3005
R19394 GND.n7414 GND.n7413 9.3005
R19395 GND.n7415 GND.n633 9.3005
R19396 GND.n7417 GND.n7416 9.3005
R19397 GND.n629 GND.n628 9.3005
R19398 GND.n7424 GND.n7423 9.3005
R19399 GND.n7425 GND.n627 9.3005
R19400 GND.n7427 GND.n7426 9.3005
R19401 GND.n623 GND.n622 9.3005
R19402 GND.n7434 GND.n7433 9.3005
R19403 GND.n7435 GND.n621 9.3005
R19404 GND.n7437 GND.n7436 9.3005
R19405 GND.n617 GND.n616 9.3005
R19406 GND.n7444 GND.n7443 9.3005
R19407 GND.n7445 GND.n615 9.3005
R19408 GND.n7447 GND.n7446 9.3005
R19409 GND.n611 GND.n610 9.3005
R19410 GND.n7454 GND.n7453 9.3005
R19411 GND.n7455 GND.n609 9.3005
R19412 GND.n7457 GND.n7456 9.3005
R19413 GND.n605 GND.n604 9.3005
R19414 GND.n7464 GND.n7463 9.3005
R19415 GND.n7465 GND.n603 9.3005
R19416 GND.n7467 GND.n7466 9.3005
R19417 GND.n599 GND.n598 9.3005
R19418 GND.n7474 GND.n7473 9.3005
R19419 GND.n7475 GND.n597 9.3005
R19420 GND.n7477 GND.n7476 9.3005
R19421 GND.n593 GND.n592 9.3005
R19422 GND.n7484 GND.n7483 9.3005
R19423 GND.n7485 GND.n591 9.3005
R19424 GND.n7487 GND.n7486 9.3005
R19425 GND.n587 GND.n586 9.3005
R19426 GND.n7494 GND.n7493 9.3005
R19427 GND.n7495 GND.n585 9.3005
R19428 GND.n7497 GND.n7496 9.3005
R19429 GND.n581 GND.n580 9.3005
R19430 GND.n7504 GND.n7503 9.3005
R19431 GND.n7505 GND.n579 9.3005
R19432 GND.n7507 GND.n7506 9.3005
R19433 GND.n575 GND.n574 9.3005
R19434 GND.n7514 GND.n7513 9.3005
R19435 GND.n7515 GND.n573 9.3005
R19436 GND.n7517 GND.n7516 9.3005
R19437 GND.n569 GND.n568 9.3005
R19438 GND.n7524 GND.n7523 9.3005
R19439 GND.n7525 GND.n567 9.3005
R19440 GND.n7527 GND.n7526 9.3005
R19441 GND.n563 GND.n562 9.3005
R19442 GND.n7534 GND.n7533 9.3005
R19443 GND.n7535 GND.n561 9.3005
R19444 GND.n7537 GND.n7536 9.3005
R19445 GND.n557 GND.n556 9.3005
R19446 GND.n7544 GND.n7543 9.3005
R19447 GND.n7545 GND.n555 9.3005
R19448 GND.n7547 GND.n7546 9.3005
R19449 GND.n551 GND.n550 9.3005
R19450 GND.n7554 GND.n7553 9.3005
R19451 GND.n7555 GND.n549 9.3005
R19452 GND.n7559 GND.n7556 9.3005
R19453 GND.n7558 GND.n7557 9.3005
R19454 GND.n7337 GND.n7336 9.3005
R19455 GND.n4262 GND.n4261 9.3005
R19456 GND.n4263 GND.n3077 9.3005
R19457 GND.n4270 GND.n4264 9.3005
R19458 GND.n4269 GND.n4265 9.3005
R19459 GND.n4268 GND.n4266 9.3005
R19460 GND.n3061 GND.n3060 9.3005
R19461 GND.n4300 GND.n4299 9.3005
R19462 GND.n4301 GND.n3059 9.3005
R19463 GND.n4318 GND.n4302 9.3005
R19464 GND.n4317 GND.n4303 9.3005
R19465 GND.n4316 GND.n4304 9.3005
R19466 GND.n4307 GND.n4305 9.3005
R19467 GND.n4312 GND.n4308 9.3005
R19468 GND.n4311 GND.n4310 9.3005
R19469 GND.n4309 GND.n3047 9.3005
R19470 GND.n4419 GND.n3046 9.3005
R19471 GND.n4421 GND.n4420 9.3005
R19472 GND.n4422 GND.n3045 9.3005
R19473 GND.n4424 GND.n4423 9.3005
R19474 GND.n3043 GND.n3042 9.3005
R19475 GND.n4429 GND.n4428 9.3005
R19476 GND.n4430 GND.n3041 9.3005
R19477 GND.n4440 GND.n4431 9.3005
R19478 GND.n4439 GND.n4432 9.3005
R19479 GND.n4438 GND.n4433 9.3005
R19480 GND.n4436 GND.n4435 9.3005
R19481 GND.n4434 GND.n3016 9.3005
R19482 GND.n3014 GND.n3013 9.3005
R19483 GND.n4465 GND.n4464 9.3005
R19484 GND.n4466 GND.n3012 9.3005
R19485 GND.n4485 GND.n4467 9.3005
R19486 GND.n4484 GND.n4468 9.3005
R19487 GND.n4483 GND.n4469 9.3005
R19488 GND.n4479 GND.n4470 9.3005
R19489 GND.n4478 GND.n4471 9.3005
R19490 GND.n4477 GND.n4472 9.3005
R19491 GND.n4474 GND.n4473 9.3005
R19492 GND.n2993 GND.n2992 9.3005
R19493 GND.n4537 GND.n4536 9.3005
R19494 GND.n4538 GND.n2991 9.3005
R19495 GND.n4542 GND.n4539 9.3005
R19496 GND.n4541 GND.n4540 9.3005
R19497 GND.n2986 GND.n2985 9.3005
R19498 GND.n4565 GND.n4564 9.3005
R19499 GND.n4566 GND.n2984 9.3005
R19500 GND.n4568 GND.n4567 9.3005
R19501 GND.n2982 GND.n2981 9.3005
R19502 GND.n4573 GND.n4572 9.3005
R19503 GND.n4574 GND.n2980 9.3005
R19504 GND.n4576 GND.n4575 9.3005
R19505 GND.n2978 GND.n2977 9.3005
R19506 GND.n4634 GND.n4633 9.3005
R19507 GND.n4635 GND.n2976 9.3005
R19508 GND.n4638 GND.n4637 9.3005
R19509 GND.n4636 GND.n2966 9.3005
R19510 GND.n4676 GND.n2967 9.3005
R19511 GND.n4677 GND.n2965 9.3005
R19512 GND.n4680 GND.n4679 9.3005
R19513 GND.n4681 GND.n2964 9.3005
R19514 GND.n4683 GND.n4682 9.3005
R19515 GND.n2956 GND.n2955 9.3005
R19516 GND.n4697 GND.n4696 9.3005
R19517 GND.n4698 GND.n2954 9.3005
R19518 GND.n4700 GND.n4699 9.3005
R19519 GND.n2950 GND.n2949 9.3005
R19520 GND.n4741 GND.n4740 9.3005
R19521 GND.n4742 GND.n2948 9.3005
R19522 GND.n4750 GND.n4743 9.3005
R19523 GND.n4749 GND.n4744 9.3005
R19524 GND.n4748 GND.n4746 9.3005
R19525 GND.n4745 GND.n2933 9.3005
R19526 GND.n4794 GND.n2932 9.3005
R19527 GND.n4796 GND.n4795 9.3005
R19528 GND.n4797 GND.n2414 9.3005
R19529 GND.n3078 GND.n1743 9.3005
R19530 GND.n4230 GND.n4229 9.3005
R19531 GND.n3097 GND.n3094 9.3005
R19532 GND.n4236 GND.n3093 9.3005
R19533 GND.n4237 GND.n3092 9.3005
R19534 GND.n4238 GND.n3091 9.3005
R19535 GND.n3090 GND.n3088 9.3005
R19536 GND.n4243 GND.n3087 9.3005
R19537 GND.n4244 GND.n3086 9.3005
R19538 GND.n3085 GND.n3083 9.3005
R19539 GND.n4249 GND.n3082 9.3005
R19540 GND.n4251 GND.n4250 9.3005
R19541 GND.n4252 GND.n1975 9.3005
R19542 GND.n5776 GND.n1976 9.3005
R19543 GND.n5775 GND.n1977 9.3005
R19544 GND.n5774 GND.n1978 9.3005
R19545 GND.n3064 GND.n1979 9.3005
R19546 GND.n3067 GND.n3066 9.3005
R19547 GND.n3065 GND.n2021 9.3005
R19548 GND.n5755 GND.n2022 9.3005
R19549 GND.n5754 GND.n2023 9.3005
R19550 GND.n5753 GND.n2024 9.3005
R19551 GND.n2067 GND.n2025 9.3005
R19552 GND.n2069 GND.n2068 9.3005
R19553 GND.n2073 GND.n2072 9.3005
R19554 GND.n2074 GND.n2066 9.3005
R19555 GND.n5728 GND.n2075 9.3005
R19556 GND.n5727 GND.n2076 9.3005
R19557 GND.n5726 GND.n2077 9.3005
R19558 GND.n3027 GND.n2078 9.3005
R19559 GND.n3029 GND.n3028 9.3005
R19560 GND.n3026 GND.n3025 9.3005
R19561 GND.n3034 GND.n3033 9.3005
R19562 GND.n3035 GND.n3024 9.3005
R19563 GND.n3037 GND.n3036 9.3005
R19564 GND.n3022 GND.n3021 9.3005
R19565 GND.n4447 GND.n4446 9.3005
R19566 GND.n4448 GND.n3020 9.3005
R19567 GND.n4458 GND.n4449 9.3005
R19568 GND.n4457 GND.n4450 9.3005
R19569 GND.n4456 GND.n4451 9.3005
R19570 GND.n4454 GND.n4453 9.3005
R19571 GND.n4452 GND.n3009 9.3005
R19572 GND.n3007 GND.n3006 9.3005
R19573 GND.n4492 GND.n4491 9.3005
R19574 GND.n4493 GND.n3005 9.3005
R19575 GND.n4504 GND.n4494 9.3005
R19576 GND.n4503 GND.n4495 9.3005
R19577 GND.n4502 GND.n4496 9.3005
R19578 GND.n4499 GND.n4498 9.3005
R19579 GND.n4497 GND.n2190 9.3005
R19580 GND.n5644 GND.n2191 9.3005
R19581 GND.n5643 GND.n2192 9.3005
R19582 GND.n5642 GND.n2193 9.3005
R19583 GND.n4603 GND.n2194 9.3005
R19584 GND.n4606 GND.n4605 9.3005
R19585 GND.n4607 GND.n4602 9.3005
R19586 GND.n4609 GND.n4608 9.3005
R19587 GND.n4600 GND.n4599 9.3005
R19588 GND.n4614 GND.n4613 9.3005
R19589 GND.n4615 GND.n4598 9.3005
R19590 GND.n4627 GND.n4616 9.3005
R19591 GND.n4626 GND.n4617 9.3005
R19592 GND.n4625 GND.n4618 9.3005
R19593 GND.n4621 GND.n4620 9.3005
R19594 GND.n4619 GND.n2274 9.3005
R19595 GND.n5590 GND.n2275 9.3005
R19596 GND.n5589 GND.n2276 9.3005
R19597 GND.n5588 GND.n2277 9.3005
R19598 GND.n2311 GND.n2278 9.3005
R19599 GND.n2314 GND.n2313 9.3005
R19600 GND.n2315 GND.n2310 9.3005
R19601 GND.n5569 GND.n2316 9.3005
R19602 GND.n5568 GND.n2317 9.3005
R19603 GND.n5567 GND.n2318 9.3005
R19604 GND.n2335 GND.n2319 9.3005
R19605 GND.n5555 GND.n2336 9.3005
R19606 GND.n5554 GND.n2337 9.3005
R19607 GND.n5553 GND.n2338 9.3005
R19608 GND.n2355 GND.n2339 9.3005
R19609 GND.n5541 GND.n2356 9.3005
R19610 GND.n5540 GND.n2357 9.3005
R19611 GND.n5539 GND.n2358 9.3005
R19612 GND.n2373 GND.n2359 9.3005
R19613 GND.n5527 GND.n2374 9.3005
R19614 GND.n5526 GND.n5525 9.3005
R19615 GND.n4254 GND.n4253 9.3005
R19616 GND.n2376 GND.n2375 9.3005
R19617 GND.n5518 GND.n2390 9.3005
R19618 GND.n5517 GND.n2391 9.3005
R19619 GND.n5516 GND.n2392 9.3005
R19620 GND.n5513 GND.n2393 9.3005
R19621 GND.n5512 GND.n2394 9.3005
R19622 GND.n5509 GND.n2395 9.3005
R19623 GND.n5508 GND.n2396 9.3005
R19624 GND.n5505 GND.n2397 9.3005
R19625 GND.n5504 GND.n2398 9.3005
R19626 GND.n5524 GND.n5523 9.3005
R19627 GND.n2930 GND.n2929 9.3005
R19628 GND.n2927 GND.n2924 9.3005
R19629 GND.n2923 GND.n2922 9.3005
R19630 GND.n2921 GND.n2918 9.3005
R19631 GND.n2917 GND.n2916 9.3005
R19632 GND.n2915 GND.n2912 9.3005
R19633 GND.n2911 GND.n2910 9.3005
R19634 GND.n2909 GND.n2906 9.3005
R19635 GND.n2905 GND.n2904 9.3005
R19636 GND.n2903 GND.n2901 9.3005
R19637 GND.n2931 GND.n2898 9.3005
R19638 GND.n4800 GND.n4799 9.3005
R19639 GND.n5501 GND.n2399 9.3005
R19640 GND.n5500 GND.n2400 9.3005
R19641 GND.n5497 GND.n2401 9.3005
R19642 GND.n5496 GND.n2402 9.3005
R19643 GND.n5493 GND.n2403 9.3005
R19644 GND.n5492 GND.n2404 9.3005
R19645 GND.n5489 GND.n2405 9.3005
R19646 GND.n5488 GND.n2406 9.3005
R19647 GND.n5485 GND.n2410 9.3005
R19648 GND.n5484 GND.n2411 9.3005
R19649 GND.n5481 GND.n2412 9.3005
R19650 GND.n5480 GND.n2413 9.3005
R19651 GND.n4912 GND.n2895 9.3005
R19652 GND.n4914 GND.n4913 9.3005
R19653 GND.n4915 GND.n2894 9.3005
R19654 GND.n4919 GND.n4916 9.3005
R19655 GND.n4920 GND.n2893 9.3005
R19656 GND.n4938 GND.n4937 9.3005
R19657 GND.n4939 GND.n2892 9.3005
R19658 GND.n4941 GND.n4940 9.3005
R19659 GND.n2830 GND.n2829 9.3005
R19660 GND.n4953 GND.n4952 9.3005
R19661 GND.n4954 GND.n2828 9.3005
R19662 GND.n4956 GND.n4955 9.3005
R19663 GND.n2826 GND.n2825 9.3005
R19664 GND.n4968 GND.n4967 9.3005
R19665 GND.n4969 GND.n2824 9.3005
R19666 GND.n4971 GND.n4970 9.3005
R19667 GND.n2822 GND.n2821 9.3005
R19668 GND.n4983 GND.n4982 9.3005
R19669 GND.n4984 GND.n2820 9.3005
R19670 GND.n4986 GND.n4985 9.3005
R19671 GND.n2818 GND.n2817 9.3005
R19672 GND.n4998 GND.n4997 9.3005
R19673 GND.n4999 GND.n2816 9.3005
R19674 GND.n5011 GND.n5000 9.3005
R19675 GND.n5010 GND.n5001 9.3005
R19676 GND.n5009 GND.n5002 9.3005
R19677 GND.n5008 GND.n5003 9.3005
R19678 GND.n5005 GND.n5004 9.3005
R19679 GND.n24 GND.n22 9.3005
R19680 GND.n4911 GND.n2896 9.3005
R19681 GND.n7827 GND.n7826 9.3005
R19682 GND.n25 GND.n23 9.3005
R19683 GND.n5036 GND.n5035 9.3005
R19684 GND.n5038 GND.n5037 9.3005
R19685 GND.n2812 GND.n2811 9.3005
R19686 GND.n5050 GND.n5049 9.3005
R19687 GND.n5051 GND.n2810 9.3005
R19688 GND.n5053 GND.n5052 9.3005
R19689 GND.n2807 GND.n2806 9.3005
R19690 GND.n5064 GND.n5063 9.3005
R19691 GND.n5065 GND.n2805 9.3005
R19692 GND.n5067 GND.n5066 9.3005
R19693 GND.n2802 GND.n2801 9.3005
R19694 GND.n5078 GND.n5077 9.3005
R19695 GND.n5079 GND.n2800 9.3005
R19696 GND.n5081 GND.n5080 9.3005
R19697 GND.n2797 GND.n2796 9.3005
R19698 GND.n5092 GND.n5091 9.3005
R19699 GND.n5093 GND.n2795 9.3005
R19700 GND.n5096 GND.n5095 9.3005
R19701 GND.n5094 GND.n2788 9.3005
R19702 GND.n5177 GND.n2789 9.3005
R19703 GND.n5176 GND.n2790 9.3005
R19704 GND.n5175 GND.n2791 9.3005
R19705 GND.n5106 GND.n2792 9.3005
R19706 GND.n5165 GND.n5107 9.3005
R19707 GND.n5164 GND.n5108 9.3005
R19708 GND.n5163 GND.n5109 9.3005
R19709 GND.n5157 GND.n5110 9.3005
R19710 GND.n5156 GND.n5155 9.3005
R19711 GND.n5128 GND.n5127 9.3005
R19712 GND.n5122 GND.n5121 9.3005
R19713 GND.n5135 GND.n5134 9.3005
R19714 GND.n5136 GND.n5120 9.3005
R19715 GND.n5138 GND.n5137 9.3005
R19716 GND.n5118 GND.n5117 9.3005
R19717 GND.n5145 GND.n5144 9.3005
R19718 GND.n5146 GND.n5116 9.3005
R19719 GND.n5148 GND.n5147 9.3005
R19720 GND.n5114 GND.n5111 9.3005
R19721 GND.n5154 GND.n5153 9.3005
R19722 GND.n5126 GND.n5125 9.3005
R19723 GND.n376 GND.n375 9.3005
R19724 GND.n374 GND.n219 9.3005
R19725 GND.n373 GND.n372 9.3005
R19726 GND.n369 GND.n220 9.3005
R19727 GND.n366 GND.n221 9.3005
R19728 GND.n365 GND.n222 9.3005
R19729 GND.n362 GND.n223 9.3005
R19730 GND.n361 GND.n224 9.3005
R19731 GND.n358 GND.n225 9.3005
R19732 GND.n357 GND.n226 9.3005
R19733 GND.n354 GND.n230 9.3005
R19734 GND.n353 GND.n231 9.3005
R19735 GND.n350 GND.n232 9.3005
R19736 GND.n349 GND.n233 9.3005
R19737 GND.n346 GND.n234 9.3005
R19738 GND.n345 GND.n235 9.3005
R19739 GND.n342 GND.n236 9.3005
R19740 GND.n341 GND.n237 9.3005
R19741 GND.n338 GND.n238 9.3005
R19742 GND.n337 GND.n239 9.3005
R19743 GND.n334 GND.n240 9.3005
R19744 GND.n333 GND.n241 9.3005
R19745 GND.n330 GND.n242 9.3005
R19746 GND.n326 GND.n243 9.3005
R19747 GND.n323 GND.n244 9.3005
R19748 GND.n322 GND.n245 9.3005
R19749 GND.n319 GND.n246 9.3005
R19750 GND.n318 GND.n247 9.3005
R19751 GND.n315 GND.n248 9.3005
R19752 GND.n314 GND.n249 9.3005
R19753 GND.n311 GND.n250 9.3005
R19754 GND.n310 GND.n251 9.3005
R19755 GND.n307 GND.n252 9.3005
R19756 GND.n306 GND.n253 9.3005
R19757 GND.n303 GND.n254 9.3005
R19758 GND.n302 GND.n301 9.3005
R19759 GND.n300 GND.n255 9.3005
R19760 GND.n299 GND.n298 9.3005
R19761 GND.n295 GND.n260 9.3005
R19762 GND.n294 GND.n261 9.3005
R19763 GND.n291 GND.n262 9.3005
R19764 GND.n290 GND.n263 9.3005
R19765 GND.n287 GND.n264 9.3005
R19766 GND.n286 GND.n265 9.3005
R19767 GND.n283 GND.n266 9.3005
R19768 GND.n282 GND.n267 9.3005
R19769 GND.n279 GND.n268 9.3005
R19770 GND.n278 GND.n269 9.3005
R19771 GND.n275 GND.n274 9.3005
R19772 GND.n273 GND.n270 9.3005
R19773 GND.n377 GND.n218 9.3005
R19774 GND.n5330 GND.n5329 9.3005
R19775 GND.n2603 GND.n2601 9.3005
R19776 GND.n4926 GND.n4925 9.3005
R19777 GND.n4929 GND.n4924 9.3005
R19778 GND.n4931 GND.n4930 9.3005
R19779 GND.n4932 GND.n2641 9.3005
R19780 GND.n5309 GND.n2642 9.3005
R19781 GND.n5308 GND.n2643 9.3005
R19782 GND.n5307 GND.n2644 9.3005
R19783 GND.n4947 GND.n2645 9.3005
R19784 GND.n5297 GND.n2663 9.3005
R19785 GND.n5296 GND.n2664 9.3005
R19786 GND.n5295 GND.n2665 9.3005
R19787 GND.n4962 GND.n2666 9.3005
R19788 GND.n5285 GND.n2684 9.3005
R19789 GND.n5284 GND.n2685 9.3005
R19790 GND.n5283 GND.n2686 9.3005
R19791 GND.n4977 GND.n2687 9.3005
R19792 GND.n5273 GND.n2705 9.3005
R19793 GND.n5272 GND.n2706 9.3005
R19794 GND.n5271 GND.n2707 9.3005
R19795 GND.n4992 GND.n2708 9.3005
R19796 GND.n5261 GND.n2725 9.3005
R19797 GND.n5260 GND.n2726 9.3005
R19798 GND.n5259 GND.n2727 9.3005
R19799 GND.n5018 GND.n2728 9.3005
R19800 GND.n5021 GND.n5020 9.3005
R19801 GND.n5022 GND.n2750 9.3005
R19802 GND.n5242 GND.n2751 9.3005
R19803 GND.n5241 GND.n2752 9.3005
R19804 GND.n5240 GND.n2753 9.3005
R19805 GND.n5030 GND.n2754 9.3005
R19806 GND.n5031 GND.n53 9.3005
R19807 GND.n7815 GND.n54 9.3005
R19808 GND.n7814 GND.n55 9.3005
R19809 GND.n7813 GND.n56 9.3005
R19810 GND.n2809 GND.n57 9.3005
R19811 GND.n7803 GND.n73 9.3005
R19812 GND.n7802 GND.n74 9.3005
R19813 GND.n7801 GND.n75 9.3005
R19814 GND.n2804 GND.n76 9.3005
R19815 GND.n7791 GND.n94 9.3005
R19816 GND.n7790 GND.n95 9.3005
R19817 GND.n7789 GND.n96 9.3005
R19818 GND.n2799 GND.n97 9.3005
R19819 GND.n7779 GND.n115 9.3005
R19820 GND.n7778 GND.n116 9.3005
R19821 GND.n7777 GND.n117 9.3005
R19822 GND.n2794 GND.n118 9.3005
R19823 GND.n7767 GND.n136 9.3005
R19824 GND.n7766 GND.n137 9.3005
R19825 GND.n7765 GND.n138 9.3005
R19826 GND.n5104 GND.n139 9.3005
R19827 GND.n7755 GND.n156 9.3005
R19828 GND.n7754 GND.n157 9.3005
R19829 GND.n7753 GND.n158 9.3005
R19830 GND.n5158 GND.n159 9.3005
R19831 GND.n7743 GND.n177 9.3005
R19832 GND.n7742 GND.n7741 9.3005
R19833 GND.n2602 GND.n2600 9.3005
R19834 GND.n5329 GND.n5328 9.3005
R19835 GND.n5327 GND.n2603 9.3005
R19836 GND.n4925 GND.n2605 9.3005
R19837 GND.n4924 GND.n4923 9.3005
R19838 GND.n4931 GND.n4921 9.3005
R19839 GND.n4933 GND.n4932 9.3005
R19840 GND.n2831 GND.n2642 9.3005
R19841 GND.n4945 GND.n2643 9.3005
R19842 GND.n4946 GND.n2644 9.3005
R19843 GND.n4948 GND.n4947 9.3005
R19844 GND.n2827 GND.n2663 9.3005
R19845 GND.n4960 GND.n2664 9.3005
R19846 GND.n4961 GND.n2665 9.3005
R19847 GND.n4963 GND.n4962 9.3005
R19848 GND.n2823 GND.n2684 9.3005
R19849 GND.n4975 GND.n2685 9.3005
R19850 GND.n4976 GND.n2686 9.3005
R19851 GND.n4978 GND.n4977 9.3005
R19852 GND.n2819 GND.n2705 9.3005
R19853 GND.n4990 GND.n2706 9.3005
R19854 GND.n4991 GND.n2707 9.3005
R19855 GND.n4993 GND.n4992 9.3005
R19856 GND.n2814 GND.n2725 9.3005
R19857 GND.n5015 GND.n2726 9.3005
R19858 GND.n5016 GND.n2727 9.3005
R19859 GND.n5018 GND.n5017 9.3005
R19860 GND.n5021 GND.n2813 9.3005
R19861 GND.n5025 GND.n5022 9.3005
R19862 GND.n5026 GND.n2751 9.3005
R19863 GND.n5027 GND.n2752 9.3005
R19864 GND.n5028 GND.n2753 9.3005
R19865 GND.n5030 GND.n5029 9.3005
R19866 GND.n5042 GND.n5031 9.3005
R19867 GND.n5043 GND.n54 9.3005
R19868 GND.n5044 GND.n55 9.3005
R19869 GND.n2808 GND.n56 9.3005
R19870 GND.n5057 GND.n2809 9.3005
R19871 GND.n5058 GND.n73 9.3005
R19872 GND.n5059 GND.n74 9.3005
R19873 GND.n2803 GND.n75 9.3005
R19874 GND.n5071 GND.n2804 9.3005
R19875 GND.n5072 GND.n94 9.3005
R19876 GND.n5073 GND.n95 9.3005
R19877 GND.n2798 GND.n96 9.3005
R19878 GND.n5085 GND.n2799 9.3005
R19879 GND.n5086 GND.n115 9.3005
R19880 GND.n5087 GND.n116 9.3005
R19881 GND.n2793 GND.n117 9.3005
R19882 GND.n5100 GND.n2794 9.3005
R19883 GND.n5101 GND.n136 9.3005
R19884 GND.n5102 GND.n137 9.3005
R19885 GND.n5103 GND.n138 9.3005
R19886 GND.n5171 GND.n5104 9.3005
R19887 GND.n5170 GND.n156 9.3005
R19888 GND.n5169 GND.n157 9.3005
R19889 GND.n5105 GND.n158 9.3005
R19890 GND.n5159 GND.n5158 9.3005
R19891 GND.n179 GND.n177 9.3005
R19892 GND.n7741 GND.n7740 9.3005
R19893 GND.n2604 GND.n2602 9.3005
R19894 GND.n4902 GND.n4828 9.3005
R19895 GND.n4901 GND.n4900 9.3005
R19896 GND.n4897 GND.n4829 9.3005
R19897 GND.n4894 GND.n4893 9.3005
R19898 GND.n4892 GND.n4830 9.3005
R19899 GND.n4891 GND.n4890 9.3005
R19900 GND.n4887 GND.n4831 9.3005
R19901 GND.n4884 GND.n4883 9.3005
R19902 GND.n4882 GND.n4832 9.3005
R19903 GND.n4881 GND.n4880 9.3005
R19904 GND.n4877 GND.n4833 9.3005
R19905 GND.n4874 GND.n4873 9.3005
R19906 GND.n4872 GND.n4834 9.3005
R19907 GND.n4865 GND.n4835 9.3005
R19908 GND.n4862 GND.n4861 9.3005
R19909 GND.n4860 GND.n4836 9.3005
R19910 GND.n4859 GND.n4858 9.3005
R19911 GND.n4855 GND.n4837 9.3005
R19912 GND.n4852 GND.n4851 9.3005
R19913 GND.n4850 GND.n4838 9.3005
R19914 GND.n4849 GND.n4848 9.3005
R19915 GND.n4845 GND.n4839 9.3005
R19916 GND.n4842 GND.n4841 9.3005
R19917 GND.n4840 GND.n2555 9.3005
R19918 GND.n5407 GND.n2554 9.3005
R19919 GND.n5360 GND.n2549 9.3005
R19920 GND.n5364 GND.n5361 9.3005
R19921 GND.n5365 GND.n5359 9.3005
R19922 GND.n5368 GND.n5358 9.3005
R19923 GND.n5369 GND.n5357 9.3005
R19924 GND.n5372 GND.n5356 9.3005
R19925 GND.n5373 GND.n5355 9.3005
R19926 GND.n5376 GND.n5354 9.3005
R19927 GND.n5377 GND.n5353 9.3005
R19928 GND.n5380 GND.n5352 9.3005
R19929 GND.n5381 GND.n5351 9.3005
R19930 GND.n5384 GND.n5347 9.3005
R19931 GND.n5385 GND.n5346 9.3005
R19932 GND.n5388 GND.n5345 9.3005
R19933 GND.n5389 GND.n5344 9.3005
R19934 GND.n5392 GND.n5343 9.3005
R19935 GND.n5393 GND.n5342 9.3005
R19936 GND.n5396 GND.n5341 9.3005
R19937 GND.n5398 GND.n5340 9.3005
R19938 GND.n5399 GND.n5339 9.3005
R19939 GND.n5400 GND.n5338 9.3005
R19940 GND.n5401 GND.n5337 9.3005
R19941 GND.n4871 GND.n4870 9.3005
R19942 GND.n4906 GND.n4905 9.3005
R19943 GND.n5334 GND.n2591 9.3005
R19944 GND.n2626 GND.n2592 9.3005
R19945 GND.n2629 GND.n2628 9.3005
R19946 GND.n2630 GND.n2625 9.3005
R19947 GND.n5315 GND.n2631 9.3005
R19948 GND.n5314 GND.n2632 9.3005
R19949 GND.n5313 GND.n2633 9.3005
R19950 GND.n2652 GND.n2634 9.3005
R19951 GND.n5303 GND.n2653 9.3005
R19952 GND.n5302 GND.n2654 9.3005
R19953 GND.n5301 GND.n2655 9.3005
R19954 GND.n2673 GND.n2656 9.3005
R19955 GND.n5291 GND.n2674 9.3005
R19956 GND.n5290 GND.n2675 9.3005
R19957 GND.n5289 GND.n2676 9.3005
R19958 GND.n2694 GND.n2677 9.3005
R19959 GND.n5279 GND.n2695 9.3005
R19960 GND.n5278 GND.n2696 9.3005
R19961 GND.n5277 GND.n2697 9.3005
R19962 GND.n2715 GND.n2698 9.3005
R19963 GND.n5267 GND.n2716 9.3005
R19964 GND.n5266 GND.n2717 9.3005
R19965 GND.n5265 GND.n2718 9.3005
R19966 GND.n2719 GND.n37 9.3005
R19967 GND.n44 GND.n36 9.3005
R19968 GND.n7809 GND.n63 9.3005
R19969 GND.n7808 GND.n64 9.3005
R19970 GND.n7807 GND.n65 9.3005
R19971 GND.n83 GND.n66 9.3005
R19972 GND.n7797 GND.n84 9.3005
R19973 GND.n7796 GND.n85 9.3005
R19974 GND.n7795 GND.n86 9.3005
R19975 GND.n104 GND.n87 9.3005
R19976 GND.n7785 GND.n105 9.3005
R19977 GND.n7784 GND.n106 9.3005
R19978 GND.n7783 GND.n107 9.3005
R19979 GND.n125 GND.n108 9.3005
R19980 GND.n7773 GND.n126 9.3005
R19981 GND.n7772 GND.n127 9.3005
R19982 GND.n7771 GND.n128 9.3005
R19983 GND.n145 GND.n129 9.3005
R19984 GND.n7761 GND.n146 9.3005
R19985 GND.n7760 GND.n147 9.3005
R19986 GND.n7759 GND.n148 9.3005
R19987 GND.n166 GND.n149 9.3005
R19988 GND.n7749 GND.n167 9.3005
R19989 GND.n7748 GND.n168 9.3005
R19990 GND.n7747 GND.n169 9.3005
R19991 GND.n217 GND.n170 9.3005
R19992 GND.n5336 GND.n5335 9.3005
R19993 GND.n7820 GND.n41 9.3005
R19994 GND.n7820 GND.n7819 9.3005
R19995 GND.n3943 GND.n3324 9.3005
R19996 GND.n3945 GND.n3944 9.3005
R19997 GND.n3299 GND.n3298 9.3005
R19998 GND.n3977 GND.n3976 9.3005
R19999 GND.n3978 GND.n3297 9.3005
R20000 GND.n3982 GND.n3979 9.3005
R20001 GND.n3981 GND.n3980 9.3005
R20002 GND.n3269 GND.n3268 9.3005
R20003 GND.n4014 GND.n4013 9.3005
R20004 GND.n4015 GND.n3267 9.3005
R20005 GND.n4019 GND.n4016 9.3005
R20006 GND.n4018 GND.n4017 9.3005
R20007 GND.n3240 GND.n3239 9.3005
R20008 GND.n4051 GND.n4050 9.3005
R20009 GND.n4052 GND.n3238 9.3005
R20010 GND.n4056 GND.n4053 9.3005
R20011 GND.n4055 GND.n4054 9.3005
R20012 GND.n3211 GND.n3210 9.3005
R20013 GND.n4088 GND.n4087 9.3005
R20014 GND.n4089 GND.n3209 9.3005
R20015 GND.n4126 GND.n4090 9.3005
R20016 GND.n4125 GND.n4091 9.3005
R20017 GND.n4124 GND.n4092 9.3005
R20018 GND.n4095 GND.n4093 9.3005
R20019 GND.n4120 GND.n4096 9.3005
R20020 GND.n4119 GND.n4097 9.3005
R20021 GND.n4118 GND.n4098 9.3005
R20022 GND.n4101 GND.n4099 9.3005
R20023 GND.n4112 GND.n4102 9.3005
R20024 GND.n4111 GND.n4103 9.3005
R20025 GND.n4110 GND.n4104 9.3005
R20026 GND.n4107 GND.n4106 9.3005
R20027 GND.n4105 GND.n1888 9.3005
R20028 GND.n5801 GND.n1889 9.3005
R20029 GND.n5800 GND.n1890 9.3005
R20030 GND.n5799 GND.n1891 9.3005
R20031 GND.n1998 GND.n1892 9.3005
R20032 GND.n2001 GND.n2000 9.3005
R20033 GND.n2002 GND.n1997 9.3005
R20034 GND.n2004 GND.n2003 9.3005
R20035 GND.n1995 GND.n1994 9.3005
R20036 GND.n2009 GND.n2008 9.3005
R20037 GND.n2010 GND.n1993 9.3005
R20038 GND.n5762 GND.n2011 9.3005
R20039 GND.n5761 GND.n2012 9.3005
R20040 GND.n5760 GND.n2013 9.3005
R20041 GND.n2042 GND.n2014 9.3005
R20042 GND.n2045 GND.n2044 9.3005
R20043 GND.n2046 GND.n2041 9.3005
R20044 GND.n5742 GND.n2047 9.3005
R20045 GND.n5741 GND.n2048 9.3005
R20046 GND.n5740 GND.n2049 9.3005
R20047 GND.n2086 GND.n2050 9.3005
R20048 GND.n2089 GND.n2088 9.3005
R20049 GND.n2090 GND.n2085 9.3005
R20050 GND.n5721 GND.n2091 9.3005
R20051 GND.n5720 GND.n2092 9.3005
R20052 GND.n5719 GND.n2093 9.3005
R20053 GND.n2108 GND.n2094 9.3005
R20054 GND.n5707 GND.n2109 9.3005
R20055 GND.n5706 GND.n2110 9.3005
R20056 GND.n5705 GND.n2111 9.3005
R20057 GND.n2126 GND.n2112 9.3005
R20058 GND.n5693 GND.n2127 9.3005
R20059 GND.n5692 GND.n2128 9.3005
R20060 GND.n5691 GND.n2129 9.3005
R20061 GND.n2143 GND.n2130 9.3005
R20062 GND.n5679 GND.n2144 9.3005
R20063 GND.n5678 GND.n2145 9.3005
R20064 GND.n5677 GND.n2146 9.3005
R20065 GND.n2161 GND.n2147 9.3005
R20066 GND.n5665 GND.n2162 9.3005
R20067 GND.n5664 GND.n2163 9.3005
R20068 GND.n5663 GND.n2164 9.3005
R20069 GND.n2179 GND.n2165 9.3005
R20070 GND.n5651 GND.n2180 9.3005
R20071 GND.n5650 GND.n2181 9.3005
R20072 GND.n5649 GND.n2182 9.3005
R20073 GND.n2210 GND.n2183 9.3005
R20074 GND.n2213 GND.n2212 9.3005
R20075 GND.n2214 GND.n2209 9.3005
R20076 GND.n5630 GND.n2215 9.3005
R20077 GND.n5629 GND.n2216 9.3005
R20078 GND.n5628 GND.n2217 9.3005
R20079 GND.n2244 GND.n2218 9.3005
R20080 GND.n2245 GND.n2243 9.3005
R20081 GND.n5611 GND.n2246 9.3005
R20082 GND.n5610 GND.n2247 9.3005
R20083 GND.n5609 GND.n2248 9.3005
R20084 GND.n2263 GND.n2249 9.3005
R20085 GND.n5597 GND.n2264 9.3005
R20086 GND.n5596 GND.n2265 9.3005
R20087 GND.n5595 GND.n2266 9.3005
R20088 GND.n2295 GND.n2267 9.3005
R20089 GND.n2298 GND.n2297 9.3005
R20090 GND.n2299 GND.n2294 9.3005
R20091 GND.n5576 GND.n2300 9.3005
R20092 GND.n5575 GND.n2301 9.3005
R20093 GND.n5574 GND.n2302 9.3005
R20094 GND.n4720 GND.n2303 9.3005
R20095 GND.n4722 GND.n4721 9.3005
R20096 GND.n4719 GND.n4718 9.3005
R20097 GND.n4727 GND.n4726 9.3005
R20098 GND.n4728 GND.n4717 9.3005
R20099 GND.n4735 GND.n4729 9.3005
R20100 GND.n4734 GND.n4730 9.3005
R20101 GND.n4733 GND.n4731 9.3005
R20102 GND.n2939 GND.n2938 9.3005
R20103 GND.n4772 GND.n4771 9.3005
R20104 GND.n4773 GND.n2937 9.3005
R20105 GND.n4788 GND.n4774 9.3005
R20106 GND.n4787 GND.n4775 9.3005
R20107 GND.n4786 GND.n4776 9.3005
R20108 GND.n4778 GND.n4777 9.3005
R20109 GND.n4781 GND.n4780 9.3005
R20110 GND.n4779 GND.n2437 9.3005
R20111 GND.n5455 GND.n2438 9.3005
R20112 GND.n5454 GND.n2439 9.3005
R20113 GND.n5453 GND.n2440 9.3005
R20114 GND.n4807 GND.n2441 9.3005
R20115 GND.n4809 GND.n4808 9.3005
R20116 GND.n4806 GND.n4805 9.3005
R20117 GND.n4817 GND.n4816 9.3005
R20118 GND.n4818 GND.n4804 9.3005
R20119 GND.n4823 GND.n4819 9.3005
R20120 GND.n4822 GND.n4821 9.3005
R20121 GND.n4820 GND.n2611 9.3005
R20122 GND.n5322 GND.n2612 9.3005
R20123 GND.n5321 GND.n2613 9.3005
R20124 GND.n5320 GND.n2614 9.3005
R20125 GND.n2835 GND.n2615 9.3005
R20126 GND.n2836 GND.n2834 9.3005
R20127 GND.n2889 GND.n2837 9.3005
R20128 GND.n2888 GND.n2838 9.3005
R20129 GND.n2887 GND.n2839 9.3005
R20130 GND.n2842 GND.n2840 9.3005
R20131 GND.n2883 GND.n2843 9.3005
R20132 GND.n2882 GND.n2844 9.3005
R20133 GND.n2881 GND.n2845 9.3005
R20134 GND.n2848 GND.n2846 9.3005
R20135 GND.n2877 GND.n2849 9.3005
R20136 GND.n2876 GND.n2850 9.3005
R20137 GND.n2875 GND.n2851 9.3005
R20138 GND.n2854 GND.n2852 9.3005
R20139 GND.n2871 GND.n2855 9.3005
R20140 GND.n2870 GND.n2856 9.3005
R20141 GND.n2869 GND.n2857 9.3005
R20142 GND.n2860 GND.n2858 9.3005
R20143 GND.n2865 GND.n2861 9.3005
R20144 GND.n2864 GND.n2862 9.3005
R20145 GND.n5228 GND.n2766 9.3005
R20146 GND.n5227 GND.n2767 9.3005
R20147 GND.n2770 GND.n2768 9.3005
R20148 GND.n5223 GND.n2771 9.3005
R20149 GND.n5222 GND.n2772 9.3005
R20150 GND.n5221 GND.n2773 9.3005
R20151 GND.n2776 GND.n2774 9.3005
R20152 GND.n5217 GND.n2777 9.3005
R20153 GND.n5216 GND.n2778 9.3005
R20154 GND.n5215 GND.n2779 9.3005
R20155 GND.n2782 GND.n2780 9.3005
R20156 GND.n5211 GND.n2783 9.3005
R20157 GND.n5210 GND.n2784 9.3005
R20158 GND.n5209 GND.n2785 9.3005
R20159 GND.n5182 GND.n2786 9.3005
R20160 GND.n5205 GND.n5183 9.3005
R20161 GND.n5204 GND.n5184 9.3005
R20162 GND.n5203 GND.n5185 9.3005
R20163 GND.n5188 GND.n5186 9.3005
R20164 GND.n5199 GND.n5189 9.3005
R20165 GND.n5198 GND.n5190 9.3005
R20166 GND.n5197 GND.n5191 9.3005
R20167 GND.n5194 GND.n5193 9.3005
R20168 GND.n5192 GND.n185 9.3005
R20169 GND.n7735 GND.n186 9.3005
R20170 GND.n7734 GND.n187 9.3005
R20171 GND.n7733 GND.n188 9.3005
R20172 GND.n382 GND.n189 9.3005
R20173 GND.n7727 GND.n383 9.3005
R20174 GND.n7726 GND.n384 9.3005
R20175 GND.n7725 GND.n385 9.3005
R20176 GND.n390 GND.n386 9.3005
R20177 GND.n7719 GND.n391 9.3005
R20178 GND.n7718 GND.n392 9.3005
R20179 GND.n7717 GND.n393 9.3005
R20180 GND.n398 GND.n394 9.3005
R20181 GND.n7711 GND.n399 9.3005
R20182 GND.n7710 GND.n400 9.3005
R20183 GND.n7709 GND.n401 9.3005
R20184 GND.n406 GND.n402 9.3005
R20185 GND.n7703 GND.n407 9.3005
R20186 GND.n7702 GND.n408 9.3005
R20187 GND.n7701 GND.n409 9.3005
R20188 GND.n414 GND.n410 9.3005
R20189 GND.n7695 GND.n415 9.3005
R20190 GND.n7694 GND.n416 9.3005
R20191 GND.n7693 GND.n417 9.3005
R20192 GND.n422 GND.n418 9.3005
R20193 GND.n7687 GND.n423 9.3005
R20194 GND.n7686 GND.n424 9.3005
R20195 GND.n7685 GND.n425 9.3005
R20196 GND.n430 GND.n426 9.3005
R20197 GND.n7679 GND.n431 9.3005
R20198 GND.n7678 GND.n432 9.3005
R20199 GND.n7677 GND.n433 9.3005
R20200 GND.n438 GND.n434 9.3005
R20201 GND.n7671 GND.n439 9.3005
R20202 GND.n7670 GND.n440 9.3005
R20203 GND.n7669 GND.n441 9.3005
R20204 GND.n446 GND.n442 9.3005
R20205 GND.n7663 GND.n447 9.3005
R20206 GND.n7662 GND.n448 9.3005
R20207 GND.n7661 GND.n449 9.3005
R20208 GND.n454 GND.n450 9.3005
R20209 GND.n7655 GND.n455 9.3005
R20210 GND.n7654 GND.n456 9.3005
R20211 GND.n7653 GND.n457 9.3005
R20212 GND.n462 GND.n458 9.3005
R20213 GND.n7647 GND.n463 9.3005
R20214 GND.n7646 GND.n464 9.3005
R20215 GND.n7645 GND.n465 9.3005
R20216 GND.n470 GND.n466 9.3005
R20217 GND.n7639 GND.n471 9.3005
R20218 GND.n7638 GND.n472 9.3005
R20219 GND.n7637 GND.n473 9.3005
R20220 GND.n478 GND.n474 9.3005
R20221 GND.n7631 GND.n479 9.3005
R20222 GND.n7630 GND.n480 9.3005
R20223 GND.n7629 GND.n481 9.3005
R20224 GND.n486 GND.n482 9.3005
R20225 GND.n7623 GND.n487 9.3005
R20226 GND.n7622 GND.n488 9.3005
R20227 GND.n7621 GND.n489 9.3005
R20228 GND.n494 GND.n490 9.3005
R20229 GND.n7615 GND.n495 9.3005
R20230 GND.n7614 GND.n496 9.3005
R20231 GND.n7613 GND.n497 9.3005
R20232 GND.n502 GND.n498 9.3005
R20233 GND.n7607 GND.n503 9.3005
R20234 GND.n7606 GND.n504 9.3005
R20235 GND.n7605 GND.n505 9.3005
R20236 GND.n510 GND.n506 9.3005
R20237 GND.n7599 GND.n511 9.3005
R20238 GND.n7598 GND.n512 9.3005
R20239 GND.n7597 GND.n513 9.3005
R20240 GND.n518 GND.n514 9.3005
R20241 GND.n7591 GND.n519 9.3005
R20242 GND.n7590 GND.n520 9.3005
R20243 GND.n7589 GND.n521 9.3005
R20244 GND.n526 GND.n522 9.3005
R20245 GND.n7583 GND.n527 9.3005
R20246 GND.n7582 GND.n528 9.3005
R20247 GND.n7581 GND.n529 9.3005
R20248 GND.n534 GND.n530 9.3005
R20249 GND.n7575 GND.n535 9.3005
R20250 GND.n7574 GND.n536 9.3005
R20251 GND.n7573 GND.n537 9.3005
R20252 GND.n542 GND.n538 9.3005
R20253 GND.n7567 GND.n543 9.3005
R20254 GND.n7566 GND.n544 9.3005
R20255 GND.n7565 GND.n545 9.3005
R20256 GND.n3651 GND.n3494 9.3005
R20257 GND.n3647 GND.n3644 9.3005
R20258 GND.n3643 GND.n3495 9.3005
R20259 GND.n3642 GND.n3641 9.3005
R20260 GND.n3638 GND.n3496 9.3005
R20261 GND.n3637 GND.n3634 9.3005
R20262 GND.n3633 GND.n3497 9.3005
R20263 GND.n3632 GND.n3631 9.3005
R20264 GND.n3628 GND.n3498 9.3005
R20265 GND.n3627 GND.n3624 9.3005
R20266 GND.n3623 GND.n3499 9.3005
R20267 GND.n3622 GND.n3621 9.3005
R20268 GND.n3618 GND.n3500 9.3005
R20269 GND.n3613 GND.n3501 9.3005
R20270 GND.n3612 GND.n3611 9.3005
R20271 GND.n3608 GND.n3504 9.3005
R20272 GND.n3607 GND.n3604 9.3005
R20273 GND.n3603 GND.n3505 9.3005
R20274 GND.n3602 GND.n3601 9.3005
R20275 GND.n3598 GND.n3506 9.3005
R20276 GND.n3597 GND.n3594 9.3005
R20277 GND.n3593 GND.n3507 9.3005
R20278 GND.n3592 GND.n3591 9.3005
R20279 GND.n3588 GND.n3508 9.3005
R20280 GND.n3587 GND.n3512 9.3005
R20281 GND.n3582 GND.n3513 9.3005
R20282 GND.n3581 GND.n3580 9.3005
R20283 GND.n3577 GND.n3514 9.3005
R20284 GND.n3574 GND.n3573 9.3005
R20285 GND.n3572 GND.n3515 9.3005
R20286 GND.n3571 GND.n3570 9.3005
R20287 GND.n3567 GND.n3516 9.3005
R20288 GND.n3564 GND.n3563 9.3005
R20289 GND.n3562 GND.n3517 9.3005
R20290 GND.n3561 GND.n3560 9.3005
R20291 GND.n3557 GND.n3518 9.3005
R20292 GND.n3554 GND.n3553 9.3005
R20293 GND.n3552 GND.n3551 9.3005
R20294 GND.n3548 GND.n3522 9.3005
R20295 GND.n3547 GND.n3544 9.3005
R20296 GND.n3543 GND.n3523 9.3005
R20297 GND.n3542 GND.n3541 9.3005
R20298 GND.n3538 GND.n3524 9.3005
R20299 GND.n3537 GND.n3534 9.3005
R20300 GND.n3533 GND.n3525 9.3005
R20301 GND.n3532 GND.n3531 9.3005
R20302 GND.n3528 GND.n3526 9.3005
R20303 GND.n3527 GND.n3482 9.3005
R20304 GND.n3584 GND.n3583 9.3005
R20305 GND.n3617 GND.n3614 9.3005
R20306 GND.n3653 GND.n3652 9.3005
R20307 GND.n3673 GND.n3481 9.3005
R20308 GND.n3677 GND.n3674 9.3005
R20309 GND.n3676 GND.n3675 9.3005
R20310 GND.n3454 GND.n3453 9.3005
R20311 GND.n3709 GND.n3708 9.3005
R20312 GND.n3710 GND.n3452 9.3005
R20313 GND.n3714 GND.n3711 9.3005
R20314 GND.n3713 GND.n3712 9.3005
R20315 GND.n3425 GND.n3424 9.3005
R20316 GND.n3746 GND.n3745 9.3005
R20317 GND.n3747 GND.n3423 9.3005
R20318 GND.n3751 GND.n3748 9.3005
R20319 GND.n3750 GND.n3749 9.3005
R20320 GND.n3395 GND.n3394 9.3005
R20321 GND.n3783 GND.n3782 9.3005
R20322 GND.n3784 GND.n3393 9.3005
R20323 GND.n3788 GND.n3785 9.3005
R20324 GND.n3787 GND.n3786 9.3005
R20325 GND.n3365 GND.n3364 9.3005
R20326 GND.n3820 GND.n3819 9.3005
R20327 GND.n3821 GND.n3363 9.3005
R20328 GND.n3824 GND.n3823 9.3005
R20329 GND.n3822 GND.n3341 9.3005
R20330 GND.n3935 GND.n3342 9.3005
R20331 GND.n3309 GND.n3308 9.3005
R20332 GND.n3966 GND.n3965 9.3005
R20333 GND.n3967 GND.n3307 9.3005
R20334 GND.n3971 GND.n3968 9.3005
R20335 GND.n3970 GND.n3969 9.3005
R20336 GND.n3280 GND.n3279 9.3005
R20337 GND.n4003 GND.n4002 9.3005
R20338 GND.n4004 GND.n3278 9.3005
R20339 GND.n4008 GND.n4005 9.3005
R20340 GND.n4007 GND.n4006 9.3005
R20341 GND.n3251 GND.n3250 9.3005
R20342 GND.n4040 GND.n4039 9.3005
R20343 GND.n4041 GND.n3249 9.3005
R20344 GND.n4045 GND.n4042 9.3005
R20345 GND.n4044 GND.n4043 9.3005
R20346 GND.n3221 GND.n3220 9.3005
R20347 GND.n4077 GND.n4076 9.3005
R20348 GND.n4078 GND.n3219 9.3005
R20349 GND.n4082 GND.n4079 9.3005
R20350 GND.n4081 GND.n4080 9.3005
R20351 GND.n3194 GND.n3193 9.3005
R20352 GND.n4143 GND.n4142 9.3005
R20353 GND.n4144 GND.n3192 9.3005
R20354 GND.n4147 GND.n4145 9.3005
R20355 GND.n4146 GND.n1785 9.3005
R20356 GND.n3672 GND.n3671 9.3005
R20357 GND.n3343 GND.n3329 9.3005
R20358 GND.n3910 GND.n3329 9.3005
R20359 GND.n6170 GND.n1450 9.3005
R20360 GND.n6169 GND.n1451 9.3005
R20361 GND.n6168 GND.n1452 9.3005
R20362 GND.n1457 GND.n1453 9.3005
R20363 GND.n6162 GND.n1458 9.3005
R20364 GND.n6161 GND.n1459 9.3005
R20365 GND.n6160 GND.n1460 9.3005
R20366 GND.n1465 GND.n1461 9.3005
R20367 GND.n6154 GND.n1466 9.3005
R20368 GND.n6153 GND.n1467 9.3005
R20369 GND.n6152 GND.n1468 9.3005
R20370 GND.n1473 GND.n1469 9.3005
R20371 GND.n6146 GND.n1474 9.3005
R20372 GND.n6145 GND.n1475 9.3005
R20373 GND.n6144 GND.n1476 9.3005
R20374 GND.n1481 GND.n1477 9.3005
R20375 GND.n6138 GND.n1482 9.3005
R20376 GND.n6137 GND.n1483 9.3005
R20377 GND.n6136 GND.n1484 9.3005
R20378 GND.n1489 GND.n1485 9.3005
R20379 GND.n6130 GND.n1490 9.3005
R20380 GND.n6129 GND.n1491 9.3005
R20381 GND.n6128 GND.n1492 9.3005
R20382 GND.n1497 GND.n1493 9.3005
R20383 GND.n6122 GND.n1498 9.3005
R20384 GND.n6121 GND.n1499 9.3005
R20385 GND.n6120 GND.n1500 9.3005
R20386 GND.n1505 GND.n1501 9.3005
R20387 GND.n6114 GND.n1506 9.3005
R20388 GND.n6113 GND.n1507 9.3005
R20389 GND.n6112 GND.n1508 9.3005
R20390 GND.n1513 GND.n1509 9.3005
R20391 GND.n6106 GND.n1514 9.3005
R20392 GND.n6105 GND.n1515 9.3005
R20393 GND.n6104 GND.n1516 9.3005
R20394 GND.n1521 GND.n1517 9.3005
R20395 GND.n6098 GND.n1522 9.3005
R20396 GND.n6097 GND.n1523 9.3005
R20397 GND.n6096 GND.n1524 9.3005
R20398 GND.n1529 GND.n1525 9.3005
R20399 GND.n6090 GND.n1530 9.3005
R20400 GND.n6089 GND.n1531 9.3005
R20401 GND.n6088 GND.n1532 9.3005
R20402 GND.n1537 GND.n1533 9.3005
R20403 GND.n6082 GND.n1538 9.3005
R20404 GND.n6081 GND.n1539 9.3005
R20405 GND.n6080 GND.n1540 9.3005
R20406 GND.n1545 GND.n1541 9.3005
R20407 GND.n6074 GND.n1546 9.3005
R20408 GND.n6073 GND.n1547 9.3005
R20409 GND.n6072 GND.n1548 9.3005
R20410 GND.n1553 GND.n1549 9.3005
R20411 GND.n6066 GND.n1554 9.3005
R20412 GND.n6065 GND.n1555 9.3005
R20413 GND.n6064 GND.n1556 9.3005
R20414 GND.n1561 GND.n1557 9.3005
R20415 GND.n6058 GND.n1562 9.3005
R20416 GND.n6057 GND.n1563 9.3005
R20417 GND.n6056 GND.n1564 9.3005
R20418 GND.n1569 GND.n1565 9.3005
R20419 GND.n6050 GND.n1570 9.3005
R20420 GND.n6049 GND.n1571 9.3005
R20421 GND.n6048 GND.n1572 9.3005
R20422 GND.n1577 GND.n1573 9.3005
R20423 GND.n6042 GND.n1578 9.3005
R20424 GND.n6041 GND.n1579 9.3005
R20425 GND.n6040 GND.n1580 9.3005
R20426 GND.n1585 GND.n1581 9.3005
R20427 GND.n6034 GND.n1586 9.3005
R20428 GND.n6033 GND.n1587 9.3005
R20429 GND.n6032 GND.n1588 9.3005
R20430 GND.n1593 GND.n1589 9.3005
R20431 GND.n6026 GND.n1594 9.3005
R20432 GND.n6025 GND.n1595 9.3005
R20433 GND.n6024 GND.n1596 9.3005
R20434 GND.n1601 GND.n1597 9.3005
R20435 GND.n6018 GND.n1602 9.3005
R20436 GND.n6017 GND.n1603 9.3005
R20437 GND.n6016 GND.n1604 9.3005
R20438 GND.n1609 GND.n1605 9.3005
R20439 GND.n6010 GND.n1610 9.3005
R20440 GND.n6009 GND.n1611 9.3005
R20441 GND.n6008 GND.n1612 9.3005
R20442 GND.n3486 GND.n1613 9.3005
R20443 GND.n3487 GND.n3485 9.3005
R20444 GND.n3489 GND.n3488 9.3005
R20445 GND.n3473 GND.n3472 9.3005
R20446 GND.n3683 GND.n3682 9.3005
R20447 GND.n3684 GND.n3471 9.3005
R20448 GND.n3688 GND.n3685 9.3005
R20449 GND.n3687 GND.n3686 9.3005
R20450 GND.n3443 GND.n3442 9.3005
R20451 GND.n3720 GND.n3719 9.3005
R20452 GND.n3721 GND.n3441 9.3005
R20453 GND.n3725 GND.n3722 9.3005
R20454 GND.n3724 GND.n3723 9.3005
R20455 GND.n3414 GND.n3413 9.3005
R20456 GND.n3757 GND.n3756 9.3005
R20457 GND.n3758 GND.n3412 9.3005
R20458 GND.n3762 GND.n3759 9.3005
R20459 GND.n3761 GND.n3760 9.3005
R20460 GND.n3385 GND.n3384 9.3005
R20461 GND.n3794 GND.n3793 9.3005
R20462 GND.n3795 GND.n3383 9.3005
R20463 GND.n3805 GND.n3796 9.3005
R20464 GND.n3804 GND.n3797 9.3005
R20465 GND.n3803 GND.n3798 9.3005
R20466 GND.n3800 GND.n3799 9.3005
R20467 GND.n3332 GND.n3331 9.3005
R20468 GND.n3941 GND.n3940 9.3005
R20469 GND.n1449 GND.n1448 9.3005
R20470 GND.n6177 GND.n1443 9.3005
R20471 GND.n6178 GND.n1442 9.3005
R20472 GND.n1441 GND.n1437 9.3005
R20473 GND.n6184 GND.n1436 9.3005
R20474 GND.n6185 GND.n1435 9.3005
R20475 GND.n6186 GND.n1434 9.3005
R20476 GND.n1433 GND.n1429 9.3005
R20477 GND.n6192 GND.n1428 9.3005
R20478 GND.n6193 GND.n1427 9.3005
R20479 GND.n6194 GND.n1426 9.3005
R20480 GND.n1425 GND.n1421 9.3005
R20481 GND.n6200 GND.n1420 9.3005
R20482 GND.n6201 GND.n1419 9.3005
R20483 GND.n6202 GND.n1418 9.3005
R20484 GND.n1417 GND.n1413 9.3005
R20485 GND.n6208 GND.n1412 9.3005
R20486 GND.n6209 GND.n1411 9.3005
R20487 GND.n6210 GND.n1410 9.3005
R20488 GND.n1409 GND.n1405 9.3005
R20489 GND.n6216 GND.n1404 9.3005
R20490 GND.n6217 GND.n1403 9.3005
R20491 GND.n6218 GND.n1402 9.3005
R20492 GND.n1401 GND.n1397 9.3005
R20493 GND.n6224 GND.n1396 9.3005
R20494 GND.n6225 GND.n1395 9.3005
R20495 GND.n6226 GND.n1394 9.3005
R20496 GND.n1393 GND.n1389 9.3005
R20497 GND.n6232 GND.n1388 9.3005
R20498 GND.n6233 GND.n1387 9.3005
R20499 GND.n6234 GND.n1386 9.3005
R20500 GND.n1385 GND.n1381 9.3005
R20501 GND.n6240 GND.n1380 9.3005
R20502 GND.n6241 GND.n1379 9.3005
R20503 GND.n6242 GND.n1378 9.3005
R20504 GND.n1377 GND.n1373 9.3005
R20505 GND.n6248 GND.n1372 9.3005
R20506 GND.n6249 GND.n1371 9.3005
R20507 GND.n6250 GND.n1370 9.3005
R20508 GND.n1369 GND.n1365 9.3005
R20509 GND.n6256 GND.n1364 9.3005
R20510 GND.n6257 GND.n1363 9.3005
R20511 GND.n6258 GND.n1362 9.3005
R20512 GND.n1361 GND.n1357 9.3005
R20513 GND.n6264 GND.n1356 9.3005
R20514 GND.n6265 GND.n1355 9.3005
R20515 GND.n6266 GND.n1354 9.3005
R20516 GND.n1353 GND.n1349 9.3005
R20517 GND.n6272 GND.n1348 9.3005
R20518 GND.n6273 GND.n1347 9.3005
R20519 GND.n6274 GND.n1346 9.3005
R20520 GND.n1345 GND.n1341 9.3005
R20521 GND.n6280 GND.n1340 9.3005
R20522 GND.n6281 GND.n1339 9.3005
R20523 GND.n6282 GND.n1338 9.3005
R20524 GND.n1337 GND.n1333 9.3005
R20525 GND.n6288 GND.n1332 9.3005
R20526 GND.n6289 GND.n1331 9.3005
R20527 GND.n6290 GND.n1330 9.3005
R20528 GND.n1329 GND.n1325 9.3005
R20529 GND.n6296 GND.n1324 9.3005
R20530 GND.n6297 GND.n1323 9.3005
R20531 GND.n6298 GND.n1322 9.3005
R20532 GND.n1321 GND.n1317 9.3005
R20533 GND.n6304 GND.n1316 9.3005
R20534 GND.n6305 GND.n1315 9.3005
R20535 GND.n6306 GND.n1314 9.3005
R20536 GND.n1313 GND.n1309 9.3005
R20537 GND.n6312 GND.n1308 9.3005
R20538 GND.n6313 GND.n1307 9.3005
R20539 GND.n6314 GND.n1306 9.3005
R20540 GND.n1305 GND.n1301 9.3005
R20541 GND.n6320 GND.n1300 9.3005
R20542 GND.n6321 GND.n1299 9.3005
R20543 GND.n6322 GND.n1298 9.3005
R20544 GND.n1297 GND.n1293 9.3005
R20545 GND.n6328 GND.n1292 9.3005
R20546 GND.n6329 GND.n1291 9.3005
R20547 GND.n6330 GND.n1290 9.3005
R20548 GND.n1289 GND.n1285 9.3005
R20549 GND.n6336 GND.n1284 9.3005
R20550 GND.n6337 GND.n1283 9.3005
R20551 GND.n6338 GND.n1282 9.3005
R20552 GND.n1281 GND.n1277 9.3005
R20553 GND.n6344 GND.n1276 9.3005
R20554 GND.n6345 GND.n1275 9.3005
R20555 GND.n6346 GND.n1274 9.3005
R20556 GND.n1273 GND.n1269 9.3005
R20557 GND.n6352 GND.n1268 9.3005
R20558 GND.n6354 GND.n6353 9.3005
R20559 GND.n6176 GND.n1444 9.3005
R20560 GND.n5939 GND.n5938 9.3005
R20561 GND.n5937 GND.n1706 9.3005
R20562 GND.n5936 GND.n5935 9.3005
R20563 GND.n5934 GND.n1708 9.3005
R20564 GND.n5933 GND.n5932 9.3005
R20565 GND.n5931 GND.n1712 9.3005
R20566 GND.n5930 GND.n5929 9.3005
R20567 GND.n5928 GND.n1713 9.3005
R20568 GND.n5927 GND.n5926 9.3005
R20569 GND.n5925 GND.n1717 9.3005
R20570 GND.n5924 GND.n5923 9.3005
R20571 GND.n5922 GND.n1718 9.3005
R20572 GND.n5921 GND.n5920 9.3005
R20573 GND.n5919 GND.n1722 9.3005
R20574 GND.n5918 GND.n5917 9.3005
R20575 GND.n5916 GND.n1723 9.3005
R20576 GND.n5915 GND.n5914 9.3005
R20577 GND.n5913 GND.n1727 9.3005
R20578 GND.n5912 GND.n5911 9.3005
R20579 GND.n5910 GND.n1728 9.3005
R20580 GND.n5909 GND.n5908 9.3005
R20581 GND.n5907 GND.n1732 9.3005
R20582 GND.n5906 GND.n5905 9.3005
R20583 GND.n5904 GND.n1733 9.3005
R20584 GND.n5903 GND.n5902 9.3005
R20585 GND.n5901 GND.n1737 9.3005
R20586 GND.n5900 GND.n5899 9.3005
R20587 GND.n5898 GND.n1738 9.3005
R20588 GND.n5897 GND.n5896 9.3005
R20589 GND.n5895 GND.n1742 9.3005
R20590 GND.n4152 GND.n4151 9.3005
R20591 GND.n4214 GND.n4213 9.3005
R20592 GND.n4212 GND.n4211 9.3005
R20593 GND.n4163 GND.n4162 9.3005
R20594 GND.n4206 GND.n4205 9.3005
R20595 GND.n4204 GND.n4203 9.3005
R20596 GND.n4174 GND.n4173 9.3005
R20597 GND.n4195 GND.n4194 9.3005
R20598 GND.n4193 GND.n4192 9.3005
R20599 GND.n4184 GND.n1747 9.3005
R20600 GND.n5893 GND.n5892 9.3005
R20601 GND.n4220 GND.n4219 9.3005
R20602 GND.n4191 GND.n4190 9.3005
R20603 GND.n4180 GND.n4179 9.3005
R20604 GND.n4197 GND.n4196 9.3005
R20605 GND.n4170 GND.n4169 9.3005
R20606 GND.n4208 GND.n4207 9.3005
R20607 GND.n4210 GND.n4209 9.3005
R20608 GND.n4157 GND.n4156 9.3005
R20609 GND.n4216 GND.n4215 9.3005
R20610 GND.n4218 GND.n4217 9.3005
R20611 GND.n3098 GND.n3096 9.3005
R20612 GND.n4202 GND.n4201 9.3005
R20613 GND.n4189 GND.n1744 9.3005
R20614 GND.n5854 GND.n1817 9.3005
R20615 GND.n5856 GND.n5855 9.3005
R20616 GND.n5857 GND.n1812 9.3005
R20617 GND.n5859 GND.n5858 9.3005
R20618 GND.n5860 GND.n1811 9.3005
R20619 GND.n5862 GND.n5861 9.3005
R20620 GND.n5863 GND.n1806 9.3005
R20621 GND.n5865 GND.n5864 9.3005
R20622 GND.n5866 GND.n1805 9.3005
R20623 GND.n5868 GND.n5867 9.3005
R20624 GND.n5869 GND.n1798 9.3005
R20625 GND.n5872 GND.n5871 9.3005
R20626 GND.n5873 GND.n1797 9.3005
R20627 GND.n5875 GND.n5874 9.3005
R20628 GND.n5876 GND.n1792 9.3005
R20629 GND.n5878 GND.n5877 9.3005
R20630 GND.n5879 GND.n1791 9.3005
R20631 GND.n5881 GND.n5880 9.3005
R20632 GND.n5882 GND.n1786 9.3005
R20633 GND.n5884 GND.n5883 9.3005
R20634 GND.n5885 GND.n1784 9.3005
R20635 GND.n5887 GND.n5886 9.3005
R20636 GND.n1819 GND.n1818 9.3005
R20637 GND.n3133 GND.n3132 9.3005
R20638 GND.n3134 GND.n3129 9.3005
R20639 GND.n3138 GND.n3137 9.3005
R20640 GND.n3139 GND.n3126 9.3005
R20641 GND.n3141 GND.n3140 9.3005
R20642 GND.n3142 GND.n3125 9.3005
R20643 GND.n3146 GND.n3145 9.3005
R20644 GND.n3147 GND.n3122 9.3005
R20645 GND.n3149 GND.n3148 9.3005
R20646 GND.n3150 GND.n3121 9.3005
R20647 GND.n3154 GND.n3153 9.3005
R20648 GND.n3155 GND.n3118 9.3005
R20649 GND.n3157 GND.n3156 9.3005
R20650 GND.n3158 GND.n3115 9.3005
R20651 GND.n3162 GND.n3161 9.3005
R20652 GND.n3163 GND.n3112 9.3005
R20653 GND.n3165 GND.n3164 9.3005
R20654 GND.n3166 GND.n3111 9.3005
R20655 GND.n3170 GND.n3169 9.3005
R20656 GND.n3171 GND.n3108 9.3005
R20657 GND.n3173 GND.n3172 9.3005
R20658 GND.n3174 GND.n3107 9.3005
R20659 GND.n3178 GND.n3177 9.3005
R20660 GND.n3179 GND.n3104 9.3005
R20661 GND.n3183 GND.n3180 9.3005
R20662 GND.n3184 GND.n3099 9.3005
R20663 GND.n3664 GND.n3657 9.3005
R20664 GND.n3663 GND.n3658 9.3005
R20665 GND.n3661 GND.n3660 9.3005
R20666 GND.n3463 GND.n3461 9.3005
R20667 GND.n3704 GND.n3703 9.3005
R20668 GND.n3464 GND.n3462 9.3005
R20669 GND.n3699 GND.n3695 9.3005
R20670 GND.n3698 GND.n3697 9.3005
R20671 GND.n3434 GND.n3432 9.3005
R20672 GND.n3741 GND.n3740 9.3005
R20673 GND.n3435 GND.n3433 9.3005
R20674 GND.n3736 GND.n3732 9.3005
R20675 GND.n3735 GND.n3734 9.3005
R20676 GND.n3405 GND.n3403 9.3005
R20677 GND.n3778 GND.n3777 9.3005
R20678 GND.n3406 GND.n3404 9.3005
R20679 GND.n3773 GND.n3769 9.3005
R20680 GND.n3772 GND.n3771 9.3005
R20681 GND.n3375 GND.n3373 9.3005
R20682 GND.n3815 GND.n3814 9.3005
R20683 GND.n3377 GND.n3374 9.3005
R20684 GND.n3376 GND.n3356 9.3005
R20685 GND.n3832 GND.n3355 9.3005
R20686 GND.n3834 GND.n3833 9.3005
R20687 GND.n3352 GND.n3350 9.3005
R20688 GND.n3928 GND.n3927 9.3005
R20689 GND.n3353 GND.n3351 9.3005
R20690 GND.n3923 GND.n3842 9.3005
R20691 GND.n3922 GND.n3843 9.3005
R20692 GND.n3921 GND.n3844 9.3005
R20693 GND.n3862 GND.n3845 9.3005
R20694 GND.n3917 GND.n3850 9.3005
R20695 GND.n3916 GND.n3851 9.3005
R20696 GND.n3915 GND.n3914 9.3005
R20697 GND.n3317 GND.n3315 9.3005
R20698 GND.n3961 GND.n3960 9.3005
R20699 GND.n3318 GND.n3316 9.3005
R20700 GND.n3956 GND.n3952 9.3005
R20701 GND.n3955 GND.n3954 9.3005
R20702 GND.n3289 GND.n3287 9.3005
R20703 GND.n3998 GND.n3997 9.3005
R20704 GND.n3290 GND.n3288 9.3005
R20705 GND.n3993 GND.n3989 9.3005
R20706 GND.n3992 GND.n3991 9.3005
R20707 GND.n3260 GND.n3258 9.3005
R20708 GND.n4035 GND.n4034 9.3005
R20709 GND.n3261 GND.n3259 9.3005
R20710 GND.n4030 GND.n4026 9.3005
R20711 GND.n4029 GND.n4028 9.3005
R20712 GND.n3231 GND.n3229 9.3005
R20713 GND.n4072 GND.n4071 9.3005
R20714 GND.n3232 GND.n3230 9.3005
R20715 GND.n4067 GND.n4063 9.3005
R20716 GND.n4066 GND.n4065 9.3005
R20717 GND.n3202 GND.n3200 9.3005
R20718 GND.n4138 GND.n4137 9.3005
R20719 GND.n3203 GND.n3201 9.3005
R20720 GND.n3189 GND.n3100 9.3005
R20721 GND.n4226 GND.n3101 9.3005
R20722 GND.n3665 GND.n3655 9.3005
R20723 GND.n3664 GND.n3493 9.3005
R20724 GND.n3663 GND.n3662 9.3005
R20725 GND.n3661 GND.n3465 9.3005
R20726 GND.n3693 GND.n3463 9.3005
R20727 GND.n3703 GND.n3702 9.3005
R20728 GND.n3701 GND.n3464 9.3005
R20729 GND.n3700 GND.n3699 9.3005
R20730 GND.n3698 GND.n3436 9.3005
R20731 GND.n3730 GND.n3434 9.3005
R20732 GND.n3740 GND.n3739 9.3005
R20733 GND.n3738 GND.n3435 9.3005
R20734 GND.n3737 GND.n3736 9.3005
R20735 GND.n3735 GND.n3407 9.3005
R20736 GND.n3767 GND.n3405 9.3005
R20737 GND.n3777 GND.n3776 9.3005
R20738 GND.n3775 GND.n3406 9.3005
R20739 GND.n3774 GND.n3773 9.3005
R20740 GND.n3772 GND.n3378 9.3005
R20741 GND.n3811 GND.n3375 9.3005
R20742 GND.n3814 GND.n3813 9.3005
R20743 GND.n3812 GND.n3377 9.3005
R20744 GND.n3376 GND.n3360 9.3005
R20745 GND.n3355 GND.n3354 9.3005
R20746 GND.n3835 GND.n3834 9.3005
R20747 GND.n3838 GND.n3352 9.3005
R20748 GND.n3927 GND.n3926 9.3005
R20749 GND.n3925 GND.n3353 9.3005
R20750 GND.n3924 GND.n3923 9.3005
R20751 GND.n3922 GND.n3841 9.3005
R20752 GND.n3921 GND.n3920 9.3005
R20753 GND.n3919 GND.n3845 9.3005
R20754 GND.n3918 GND.n3917 9.3005
R20755 GND.n3916 GND.n3849 9.3005
R20756 GND.n3915 GND.n3319 9.3005
R20757 GND.n3950 GND.n3317 9.3005
R20758 GND.n3960 GND.n3959 9.3005
R20759 GND.n3958 GND.n3318 9.3005
R20760 GND.n3957 GND.n3956 9.3005
R20761 GND.n3955 GND.n3291 9.3005
R20762 GND.n3987 GND.n3289 9.3005
R20763 GND.n3997 GND.n3996 9.3005
R20764 GND.n3995 GND.n3290 9.3005
R20765 GND.n3994 GND.n3993 9.3005
R20766 GND.n3992 GND.n3262 9.3005
R20767 GND.n4024 GND.n3260 9.3005
R20768 GND.n4034 GND.n4033 9.3005
R20769 GND.n4032 GND.n3261 9.3005
R20770 GND.n4031 GND.n4030 9.3005
R20771 GND.n4029 GND.n3233 9.3005
R20772 GND.n4061 GND.n3231 9.3005
R20773 GND.n4071 GND.n4070 9.3005
R20774 GND.n4069 GND.n3232 9.3005
R20775 GND.n4068 GND.n4067 9.3005
R20776 GND.n4066 GND.n3204 9.3005
R20777 GND.n4132 GND.n3202 9.3005
R20778 GND.n4137 GND.n4136 9.3005
R20779 GND.n4135 GND.n3203 9.3005
R20780 GND.n3102 GND.n3100 9.3005
R20781 GND.n4226 GND.n4225 9.3005
R20782 GND.n3666 GND.n3665 9.3005
R20783 GND.n5989 GND.n5988 9.3005
R20784 GND.n5990 GND.n1658 9.3005
R20785 GND.n5992 GND.n5991 9.3005
R20786 GND.n5993 GND.n1657 9.3005
R20787 GND.n5995 GND.n5994 9.3005
R20788 GND.n5996 GND.n1652 9.3005
R20789 GND.n5998 GND.n5997 9.3005
R20790 GND.n5999 GND.n1651 9.3005
R20791 GND.n6001 GND.n6000 9.3005
R20792 GND.n6002 GND.n1650 9.3005
R20793 GND.n5987 GND.n1666 9.3005
R20794 GND.n5986 GND.n5985 9.3005
R20795 GND.n5982 GND.n1667 9.3005
R20796 GND.n5981 GND.n5980 9.3005
R20797 GND.n5979 GND.n1671 9.3005
R20798 GND.n5978 GND.n5977 9.3005
R20799 GND.n5976 GND.n1672 9.3005
R20800 GND.n5975 GND.n5974 9.3005
R20801 GND.n5973 GND.n1676 9.3005
R20802 GND.n5972 GND.n5971 9.3005
R20803 GND.n5970 GND.n1677 9.3005
R20804 GND.n5969 GND.n5968 9.3005
R20805 GND.n5967 GND.n1681 9.3005
R20806 GND.n5966 GND.n5965 9.3005
R20807 GND.n5964 GND.n1682 9.3005
R20808 GND.n5963 GND.n5962 9.3005
R20809 GND.n5961 GND.n1686 9.3005
R20810 GND.n5960 GND.n5959 9.3005
R20811 GND.n5958 GND.n1687 9.3005
R20812 GND.n5957 GND.n5956 9.3005
R20813 GND.n5955 GND.n1691 9.3005
R20814 GND.n5954 GND.n5953 9.3005
R20815 GND.n5952 GND.n1692 9.3005
R20816 GND.n5951 GND.n5950 9.3005
R20817 GND.n5949 GND.n1696 9.3005
R20818 GND.n5948 GND.n5947 9.3005
R20819 GND.n5946 GND.n1697 9.3005
R20820 GND.n5945 GND.n5944 9.3005
R20821 GND.n5943 GND.n1701 9.3005
R20822 GND.n5942 GND.n5941 9.3005
R20823 GND.n5940 GND.n1702 9.3005
R20824 GND.n5984 GND.n5983 9.3005
R20825 GND.t153 GND.n1904 8.83141
R20826 GND.n4296 GND.n3063 8.83141
R20827 GND.n4416 GND.n3050 8.83141
R20828 GND.n3053 GND.t31 8.83141
R20829 GND.n5703 GND.n5702 8.83141
R20830 GND.n5668 GND.n5667 8.83141
R20831 GND.n2990 GND.n2989 8.83141
R20832 GND.n5607 GND.n2251 8.83141
R20833 GND.n4674 GND.t24 8.83141
R20834 GND.n4667 GND.n2283 8.83141
R20835 GND.n5550 GND.n2344 8.83141
R20836 GND.n4768 GND.t135 8.83141
R20837 GND.n4784 GND.n2420 8.83141
R20838 GND.n4364 GND.t29 8.46345
R20839 GND.n4487 GND.t29 8.46345
R20840 GND.n4561 GND.t25 8.46345
R20841 GND.n5633 GND.t25 8.46345
R20842 GND.n1883 GND.t79 8.0955
R20843 GND.n5771 GND.t60 8.0955
R20844 GND.n4320 GND.n3058 8.0955
R20845 GND.n4337 GND.n2054 8.0955
R20846 GND.n4377 GND.n2124 8.0955
R20847 GND.n4367 GND.t163 8.0955
R20848 GND.n4487 GND.n2149 8.0955
R20849 GND.n4561 GND.n4560 8.0955
R20850 GND.n4554 GND.t32 8.0955
R20851 GND.n5614 GND.n2236 8.0955
R20852 GND.n4686 GND.n4685 8.0955
R20853 GND.n5557 GND.n2333 8.0955
R20854 GND.n2426 GND.t108 8.0955
R20855 GND.n7829 GND.n7828 8.09467
R20856 GND.n1707 GND.n9 8.09467
R20857 GND.n2495 GND.n2467 7.95202
R20858 GND.n5847 GND.n1847 7.72754
R20859 GND.n5451 GND.n5450 7.72754
R20860 GND.n4258 GND.n1969 7.35959
R20861 GND.n4278 GND.n4277 7.35959
R20862 GND.n5709 GND.n2106 7.35959
R20863 GND.n5661 GND.n2167 7.35959
R20864 GND.n4533 GND.n2995 7.35959
R20865 GND.n5600 GND.n5599 7.35959
R20866 GND.n2942 GND.n2353 7.35959
R20867 GND.t52 GND.n3448 6.99164
R20868 GND.t161 GND.n4408 6.99164
R20869 GND.t27 GND.n2968 6.99164
R20870 GND.n5180 GND.t34 6.99164
R20871 GND.n5892 GND.n1747 6.78838
R20872 GND.n5153 GND.n5114 6.78838
R20873 GND.n4800 GND.n2931 6.78838
R20874 GND.n5985 GND.n1666 6.78838
R20875 GND.n4325 GND.n2036 6.62368
R20876 GND.n4331 GND.n2037 6.62368
R20877 GND.n5688 GND.n2134 6.62368
R20878 GND.n5682 GND.n2140 6.62368
R20879 GND.n4552 GND.n2220 6.62368
R20880 GND.n2230 GND.n2222 6.62368
R20881 GND.n4694 GND.n4693 6.62368
R20882 GND.n5565 GND.n5564 6.62368
R20883 GND.n329 GND.n326 6.4005
R20884 GND.n5485 GND.n2409 6.4005
R20885 GND.n4200 GND.n4197 6.4005
R20886 GND.n3587 GND.n3511 6.4005
R20887 GND.n4273 GND.n1981 5.88777
R20888 GND.n5717 GND.n5716 5.88777
R20889 GND.n4401 GND.n4400 5.88777
R20890 GND.n4515 GND.n4514 5.88777
R20891 GND.n5654 GND.n5653 5.88777
R20892 GND.n4649 GND.n2974 5.88777
R20893 GND.n5593 GND.n2269 5.88777
R20894 GND.n4769 GND.n4768 5.88777
R20895 GND.n5536 GND.n2363 5.88777
R20896 GND.n5476 GND.t117 5.88777
R20897 GND.n3 GND.n1 5.55797
R20898 GND.n15 GND.n13 5.55797
R20899 GND.n5450 GND.t144 5.51982
R20900 GND.n2490 GND.n2467 5.23686
R20901 GND.n5751 GND.n5750 5.15186
R20902 GND.n4333 GND.n2052 5.15186
R20903 GND.t31 GND.n2082 5.15186
R20904 GND.n4460 GND.n2132 5.15186
R20905 GND.n5681 GND.t163 5.15186
R20906 GND.n4367 GND.n4366 5.15186
R20907 GND.n4554 GND.n2206 5.15186
R20908 GND.t32 GND.n4553 5.15186
R20909 GND.n5620 GND.n2229 5.15186
R20910 GND.t24 GND.n4673 5.15186
R20911 GND.n5571 GND.n2307 5.15186
R20912 GND.n4703 GND.n4702 5.15186
R20913 GND.n5530 GND.t85 5.15186
R20914 GND.n6004 GND.n1647 4.78391
R20915 GND.n5764 GND.t63 4.78391
R20916 GND.t97 GND.n2350 4.78391
R20917 GND.n379 GND.n182 4.78391
R20918 GND.n5255 GND.n42 4.74817
R20919 GND.n40 GND.n34 4.74817
R20920 GND.n7821 GND.n35 4.74817
R20921 GND.n43 GND.n39 4.74817
R20922 GND.n2735 GND.n42 4.74817
R20923 GND.n2745 GND.n40 4.74817
R20924 GND.n7822 GND.n7821 4.74817
R20925 GND.n2757 GND.n39 4.74817
R20926 GND.n3333 GND.n3330 4.74817
R20927 GND.n3875 GND.n3328 4.74817
R20928 GND.n3897 GND.n3327 4.74817
R20929 GND.n3895 GND.n3326 4.74817
R20930 GND.n3891 GND.n3325 4.74817
R20931 GND.n5250 GND.n2741 4.74817
R20932 GND.n5248 GND.n5247 4.74817
R20933 GND.n2763 GND.n2762 4.74817
R20934 GND.n5234 GND.n5233 4.74817
R20935 GND.n5229 GND.n2764 4.74817
R20936 GND.n2863 GND.n2741 4.74817
R20937 GND.n5249 GND.n5248 4.74817
R20938 GND.n2762 GND.n2742 4.74817
R20939 GND.n5235 GND.n5234 4.74817
R20940 GND.n5232 GND.n2764 4.74817
R20941 GND.n3934 GND.n3933 4.74817
R20942 GND.n3886 GND.n3883 4.74817
R20943 GND.n3884 GND.n3855 4.74817
R20944 GND.n3909 GND.n3908 4.74817
R20945 GND.n3933 GND.n3932 4.74817
R20946 GND.n3883 GND.n3882 4.74817
R20947 GND.n3885 GND.n3884 4.74817
R20948 GND.n3908 GND.n3907 4.74817
R20949 GND.n3871 GND.n3330 4.74817
R20950 GND.n3872 GND.n3328 4.74817
R20951 GND.n3874 GND.n3327 4.74817
R20952 GND.n3898 GND.n3326 4.74817
R20953 GND.n3894 GND.n3325 4.74817
R20954 GND.n8 GND.n0 4.70093
R20955 GND.n21 GND.n20 4.70093
R20956 GND.n3 GND.n2 4.63843
R20957 GND.n5 GND.n4 4.63843
R20958 GND.n7 GND.n6 4.63843
R20959 GND.n15 GND.n14 4.63843
R20960 GND.n17 GND.n16 4.63843
R20961 GND.n19 GND.n18 4.63843
R20962 GND.n5408 GND.n2551 4.6132
R20963 GND.n5853 GND.n5852 4.6132
R20964 GND.n9 GND.n8 4.57909
R20965 GND.n7829 GND.n21 4.57909
R20966 GND.n5785 GND.n1965 4.41595
R20967 GND.n5765 GND.n5764 4.41595
R20968 GND.n5723 GND.n2082 4.41595
R20969 GND.n4395 GND.n3038 4.41595
R20970 GND.n4509 GND.n3001 4.41595
R20971 GND.n5647 GND.n2185 4.41595
R20972 GND.n4584 GND.n4583 4.41595
R20973 GND.n4673 GND.n2280 4.41595
R20974 GND.n5544 GND.n2350 4.41595
R20975 GND.n2415 GND.n2371 4.41595
R20976 GND.n1879 GND.n1878 4.38232
R20977 GND.n2494 GND.n2493 4.38232
R20978 GND.n12 GND.n10 4.24406
R20979 GND.n5871 GND.n5870 4.07323
R20980 GND.n5384 GND.n5350 4.07323
R20981 GND.n357 GND.n229 4.07323
R20982 GND.n3551 GND.n3521 4.07323
R20983 GND.n5797 GND.t67 3.68005
R20984 GND.n5757 GND.n2018 3.68005
R20985 GND.n5731 GND.n5730 3.68005
R20986 GND.n5696 GND.n2122 3.68005
R20987 GND.n5674 GND.n2151 3.68005
R20988 GND.n5640 GND.n5639 3.68005
R20989 GND.n4595 GND.n2238 3.68005
R20990 GND.n4663 GND.n2291 3.68005
R20991 GND.n4738 GND.n4713 3.68005
R20992 GND.n12 GND.n11 3.53792
R20993 GND.t132 GND.n1885 2.94414
R20994 GND.n1903 GND.n1902 2.94414
R20995 GND.n4259 GND.t88 2.94414
R20996 GND.t111 GND.n1972 2.94414
R20997 GND.n3076 GND.t111 2.94414
R20998 GND.n5758 GND.n2016 2.94414
R20999 GND.n3048 GND.n2063 2.94414
R21000 GND.n4386 GND.n4385 2.94414
R21001 GND.n4355 GND.n4354 2.94414
R21002 GND.n4545 GND.n2196 2.94414
R21003 GND.n4594 GND.n4593 2.94414
R21004 GND.n5579 GND.n5578 2.94414
R21005 GND.n4737 GND.n2341 2.94414
R21006 GND.n5470 GND.n2378 2.94414
R21007 GND.n5521 GND.t108 2.94414
R21008 GND.n3830 GND.t0 2.57618
R21009 GND.n3963 GND.t8 2.57618
R21010 GND.n3226 GND.t56 2.57618
R21011 GND.n2891 GND.t38 2.57618
R21012 GND.n5263 GND.t2 2.57618
R21013 GND.n7811 GND.t4 2.57618
R21014 GND.n5870 GND.n5869 2.52171
R21015 GND.n5381 GND.n5350 2.52171
R21016 GND.n354 GND.n229 2.52171
R21017 GND.n3554 GND.n3521 2.52171
R21018 GND.n7820 GND.n42 2.27742
R21019 GND.n7820 GND.n40 2.27742
R21020 GND.n7821 GND.n7820 2.27742
R21021 GND.n7820 GND.n39 2.27742
R21022 GND.n2741 GND.n38 2.27742
R21023 GND.n5248 GND.n38 2.27742
R21024 GND.n2762 GND.n38 2.27742
R21025 GND.n5234 GND.n38 2.27742
R21026 GND.n2764 GND.n38 2.27742
R21027 GND.n3933 GND.n3329 2.27742
R21028 GND.n3883 GND.n3329 2.27742
R21029 GND.n3884 GND.n3329 2.27742
R21030 GND.n3908 GND.n3329 2.27742
R21031 GND.n3942 GND.n3330 2.27742
R21032 GND.n3942 GND.n3328 2.27742
R21033 GND.n3942 GND.n3327 2.27742
R21034 GND.n3942 GND.n3326 2.27742
R21035 GND.n3942 GND.n3325 2.27742
R21036 GND.n4256 GND.n3080 2.20823
R21037 GND.n3070 GND.n3069 2.20823
R21038 GND.n5724 GND.n2080 2.20823
R21039 GND.n4442 GND.n2114 2.20823
R21040 GND.n4480 GND.n2159 2.20823
R21041 GND.n5646 GND.n2187 2.20823
R21042 GND.n5606 GND.n2253 2.20823
R21043 GND.n5586 GND.n5585 2.20823
R21044 GND.n4753 GND.n4752 2.20823
R21045 GND.t135 GND.t101 2.20823
R21046 GND.n4790 GND.t85 2.20823
R21047 GND.n5477 GND.n5476 2.20823
R21048 GND.n5895 GND.n5894 2.1585
R21049 GND.n4798 GND.n2896 2.15419
R21050 GND.n1957 GND.n1954 1.47232
R21051 GND.t42 GND.n4272 1.47232
R21052 GND.n4321 GND.n2027 1.47232
R21053 GND.n5738 GND.n5737 1.47232
R21054 GND.n4380 GND.n3017 1.47232
R21055 GND.n4365 GND.n4364 1.47232
R21056 GND.n5633 GND.n5632 1.47232
R21057 GND.n2240 GND.n2239 1.47232
R21058 GND.n5572 GND.n2305 1.47232
R21059 GND.n5558 GND.n2330 1.47232
R21060 GND.n5537 GND.t101 1.47232
R21061 GND.n2434 GND.n2428 1.47232
R21062 GND.n2434 GND.t126 1.47232
R21063 GND.n8 GND.n7 1.25984
R21064 GND.n21 GND.n19 1.25984
R21065 GND.n2541 GND.n2502 1.24928
R21066 GND.n1917 GND.n1916 1.24928
R21067 GND.n5815 GND.n5814 1.24928
R21068 GND.n5418 GND.n5417 1.24928
R21069 GND GND.n9 1.22344
R21070 GND.n5852 GND.n1819 0.970197
R21071 GND.n5408 GND.n5407 0.970197
R21072 GND.n5 GND.n3 0.92004
R21073 GND.n7 GND.n5 0.92004
R21074 GND.n17 GND.n15 0.92004
R21075 GND.n19 GND.n17 0.92004
R21076 GND.n7830 GND.n7829 0.83193
R21077 GND.n5779 GND.n5778 0.736409
R21078 GND.n5772 GND.n5771 0.736409
R21079 GND.n4407 GND.n2096 0.736409
R21080 GND.n5710 GND.n2104 0.736409
R21081 GND.n5660 GND.n2169 0.736409
R21082 GND.n2996 GND.n2177 0.736409
R21083 GND.n4622 GND.n2261 0.736409
R21084 GND.n5592 GND.n2271 0.736409
R21085 GND.n2945 GND.n2941 0.736409
R21086 GND.n4792 GND.n4791 0.736409
R21087 GND.n1861 GND.n1859 0.716017
R21088 GND.n2488 GND.n2486 0.716017
R21089 GND.n6355 GND.n6354 0.486781
R21090 GND.n7336 GND.n7335 0.486781
R21091 GND.n7557 GND.n545 0.486781
R21092 GND.n1449 GND.n1444 0.486781
R21093 GND.n5986 GND.n5984 0.479159
R21094 GND.n5155 GND.n5154 0.479158
R21095 GND.n4253 GND.n4251 0.447146
R21096 GND.n5525 GND.n5524 0.447146
R21097 GND.n5337 GND.n5336 0.444098
R21098 GND.n3672 GND.n3482 0.444098
R21099 GND.n218 GND.n217 0.444098
R21100 GND.n5886 GND.n1785 0.444098
R21101 GND.n7820 GND.n38 0.40325
R21102 GND.n3942 GND.n3329 0.40325
R21103 GND.n5889 GND.n1750 0.368454
R21104 GND.n4409 GND.t161 0.368454
R21105 GND.n2969 GND.t27 0.368454
R21106 GND.n5404 GND.n2587 0.368454
R21107 GND.n5409 GND.n2547 0.312695
R21108 GND.n5851 GND.n1823 0.312695
R21109 GND.n5851 GND.n5850 0.312695
R21110 GND.n5410 GND.n5409 0.312695
R21111 GND.n5126 GND.n178 0.302329
R21112 GND.n3654 GND.n1650 0.302329
R21113 GND.n273 GND.n178 0.267268
R21114 GND.n4905 GND.n4904 0.267268
R21115 GND.n3654 GND.n3653 0.267268
R21116 GND.n4227 GND.n3099 0.267268
R21117 GND.n7830 GND.n12 0.24114
R21118 GND.n5360 GND.n2551 0.229039
R21119 GND.n2554 GND.n2551 0.229039
R21120 GND.n5854 GND.n5853 0.229039
R21121 GND.n5853 GND.n1818 0.229039
R21122 GND.n5894 GND.n1743 0.21239
R21123 GND.n4798 GND.n4797 0.21239
R21124 GND GND.n7830 0.198213
R21125 GND.n330 GND.n329 0.194439
R21126 GND.n5488 GND.n2409 0.194439
R21127 GND.n4201 GND.n4200 0.194439
R21128 GND.n3584 GND.n3511 0.194439
R21129 GND.n6355 GND.n1263 0.152939
R21130 GND.n6363 GND.n1263 0.152939
R21131 GND.n6364 GND.n6363 0.152939
R21132 GND.n6365 GND.n6364 0.152939
R21133 GND.n6365 GND.n1257 0.152939
R21134 GND.n6373 GND.n1257 0.152939
R21135 GND.n6374 GND.n6373 0.152939
R21136 GND.n6375 GND.n6374 0.152939
R21137 GND.n6375 GND.n1251 0.152939
R21138 GND.n6383 GND.n1251 0.152939
R21139 GND.n6384 GND.n6383 0.152939
R21140 GND.n6385 GND.n6384 0.152939
R21141 GND.n6385 GND.n1245 0.152939
R21142 GND.n6393 GND.n1245 0.152939
R21143 GND.n6394 GND.n6393 0.152939
R21144 GND.n6395 GND.n6394 0.152939
R21145 GND.n6395 GND.n1239 0.152939
R21146 GND.n6403 GND.n1239 0.152939
R21147 GND.n6404 GND.n6403 0.152939
R21148 GND.n6405 GND.n6404 0.152939
R21149 GND.n6405 GND.n1233 0.152939
R21150 GND.n6413 GND.n1233 0.152939
R21151 GND.n6414 GND.n6413 0.152939
R21152 GND.n6415 GND.n6414 0.152939
R21153 GND.n6415 GND.n1227 0.152939
R21154 GND.n6423 GND.n1227 0.152939
R21155 GND.n6424 GND.n6423 0.152939
R21156 GND.n6425 GND.n6424 0.152939
R21157 GND.n6425 GND.n1221 0.152939
R21158 GND.n6433 GND.n1221 0.152939
R21159 GND.n6434 GND.n6433 0.152939
R21160 GND.n6435 GND.n6434 0.152939
R21161 GND.n6435 GND.n1215 0.152939
R21162 GND.n6443 GND.n1215 0.152939
R21163 GND.n6444 GND.n6443 0.152939
R21164 GND.n6445 GND.n6444 0.152939
R21165 GND.n6445 GND.n1209 0.152939
R21166 GND.n6453 GND.n1209 0.152939
R21167 GND.n6454 GND.n6453 0.152939
R21168 GND.n6455 GND.n6454 0.152939
R21169 GND.n6455 GND.n1203 0.152939
R21170 GND.n6463 GND.n1203 0.152939
R21171 GND.n6464 GND.n6463 0.152939
R21172 GND.n6465 GND.n6464 0.152939
R21173 GND.n6465 GND.n1197 0.152939
R21174 GND.n6473 GND.n1197 0.152939
R21175 GND.n6474 GND.n6473 0.152939
R21176 GND.n6475 GND.n6474 0.152939
R21177 GND.n6475 GND.n1191 0.152939
R21178 GND.n6483 GND.n1191 0.152939
R21179 GND.n6484 GND.n6483 0.152939
R21180 GND.n6485 GND.n6484 0.152939
R21181 GND.n6485 GND.n1185 0.152939
R21182 GND.n6493 GND.n1185 0.152939
R21183 GND.n6494 GND.n6493 0.152939
R21184 GND.n6495 GND.n6494 0.152939
R21185 GND.n6495 GND.n1179 0.152939
R21186 GND.n6503 GND.n1179 0.152939
R21187 GND.n6504 GND.n6503 0.152939
R21188 GND.n6505 GND.n6504 0.152939
R21189 GND.n6505 GND.n1173 0.152939
R21190 GND.n6513 GND.n1173 0.152939
R21191 GND.n6514 GND.n6513 0.152939
R21192 GND.n6515 GND.n6514 0.152939
R21193 GND.n6515 GND.n1167 0.152939
R21194 GND.n6523 GND.n1167 0.152939
R21195 GND.n6524 GND.n6523 0.152939
R21196 GND.n6525 GND.n6524 0.152939
R21197 GND.n6525 GND.n1161 0.152939
R21198 GND.n6533 GND.n1161 0.152939
R21199 GND.n6534 GND.n6533 0.152939
R21200 GND.n6535 GND.n6534 0.152939
R21201 GND.n6535 GND.n1155 0.152939
R21202 GND.n6543 GND.n1155 0.152939
R21203 GND.n6544 GND.n6543 0.152939
R21204 GND.n6545 GND.n6544 0.152939
R21205 GND.n6545 GND.n1149 0.152939
R21206 GND.n6553 GND.n1149 0.152939
R21207 GND.n6554 GND.n6553 0.152939
R21208 GND.n6555 GND.n6554 0.152939
R21209 GND.n6555 GND.n1143 0.152939
R21210 GND.n6563 GND.n1143 0.152939
R21211 GND.n6564 GND.n6563 0.152939
R21212 GND.n6565 GND.n6564 0.152939
R21213 GND.n6565 GND.n1137 0.152939
R21214 GND.n6573 GND.n1137 0.152939
R21215 GND.n6574 GND.n6573 0.152939
R21216 GND.n6575 GND.n6574 0.152939
R21217 GND.n6575 GND.n1131 0.152939
R21218 GND.n6583 GND.n1131 0.152939
R21219 GND.n6584 GND.n6583 0.152939
R21220 GND.n6585 GND.n6584 0.152939
R21221 GND.n6585 GND.n1125 0.152939
R21222 GND.n6593 GND.n1125 0.152939
R21223 GND.n6594 GND.n6593 0.152939
R21224 GND.n6595 GND.n6594 0.152939
R21225 GND.n6595 GND.n1119 0.152939
R21226 GND.n6603 GND.n1119 0.152939
R21227 GND.n6604 GND.n6603 0.152939
R21228 GND.n6605 GND.n6604 0.152939
R21229 GND.n6605 GND.n1113 0.152939
R21230 GND.n6613 GND.n1113 0.152939
R21231 GND.n6614 GND.n6613 0.152939
R21232 GND.n6615 GND.n6614 0.152939
R21233 GND.n6615 GND.n1107 0.152939
R21234 GND.n6623 GND.n1107 0.152939
R21235 GND.n6624 GND.n6623 0.152939
R21236 GND.n6625 GND.n6624 0.152939
R21237 GND.n6625 GND.n1101 0.152939
R21238 GND.n6633 GND.n1101 0.152939
R21239 GND.n6634 GND.n6633 0.152939
R21240 GND.n6635 GND.n6634 0.152939
R21241 GND.n6635 GND.n1095 0.152939
R21242 GND.n6643 GND.n1095 0.152939
R21243 GND.n6644 GND.n6643 0.152939
R21244 GND.n6645 GND.n6644 0.152939
R21245 GND.n6645 GND.n1089 0.152939
R21246 GND.n6653 GND.n1089 0.152939
R21247 GND.n6654 GND.n6653 0.152939
R21248 GND.n6655 GND.n6654 0.152939
R21249 GND.n6655 GND.n1083 0.152939
R21250 GND.n6663 GND.n1083 0.152939
R21251 GND.n6664 GND.n6663 0.152939
R21252 GND.n6665 GND.n6664 0.152939
R21253 GND.n6665 GND.n1077 0.152939
R21254 GND.n6673 GND.n1077 0.152939
R21255 GND.n6674 GND.n6673 0.152939
R21256 GND.n6675 GND.n6674 0.152939
R21257 GND.n6675 GND.n1071 0.152939
R21258 GND.n6683 GND.n1071 0.152939
R21259 GND.n6684 GND.n6683 0.152939
R21260 GND.n6685 GND.n6684 0.152939
R21261 GND.n6685 GND.n1065 0.152939
R21262 GND.n6693 GND.n1065 0.152939
R21263 GND.n6694 GND.n6693 0.152939
R21264 GND.n6695 GND.n6694 0.152939
R21265 GND.n6695 GND.n1059 0.152939
R21266 GND.n6703 GND.n1059 0.152939
R21267 GND.n6704 GND.n6703 0.152939
R21268 GND.n6705 GND.n6704 0.152939
R21269 GND.n6705 GND.n1053 0.152939
R21270 GND.n6713 GND.n1053 0.152939
R21271 GND.n6714 GND.n6713 0.152939
R21272 GND.n6715 GND.n6714 0.152939
R21273 GND.n6715 GND.n1047 0.152939
R21274 GND.n6723 GND.n1047 0.152939
R21275 GND.n6724 GND.n6723 0.152939
R21276 GND.n6725 GND.n6724 0.152939
R21277 GND.n6725 GND.n1041 0.152939
R21278 GND.n6733 GND.n1041 0.152939
R21279 GND.n6734 GND.n6733 0.152939
R21280 GND.n6735 GND.n6734 0.152939
R21281 GND.n6735 GND.n1035 0.152939
R21282 GND.n6743 GND.n1035 0.152939
R21283 GND.n6744 GND.n6743 0.152939
R21284 GND.n6745 GND.n6744 0.152939
R21285 GND.n6745 GND.n1029 0.152939
R21286 GND.n6753 GND.n1029 0.152939
R21287 GND.n6754 GND.n6753 0.152939
R21288 GND.n6755 GND.n6754 0.152939
R21289 GND.n6755 GND.n1023 0.152939
R21290 GND.n6763 GND.n1023 0.152939
R21291 GND.n6764 GND.n6763 0.152939
R21292 GND.n6765 GND.n6764 0.152939
R21293 GND.n6765 GND.n1017 0.152939
R21294 GND.n6773 GND.n1017 0.152939
R21295 GND.n6774 GND.n6773 0.152939
R21296 GND.n6775 GND.n6774 0.152939
R21297 GND.n6775 GND.n1011 0.152939
R21298 GND.n6783 GND.n1011 0.152939
R21299 GND.n6784 GND.n6783 0.152939
R21300 GND.n6785 GND.n6784 0.152939
R21301 GND.n6785 GND.n1005 0.152939
R21302 GND.n6793 GND.n1005 0.152939
R21303 GND.n6794 GND.n6793 0.152939
R21304 GND.n6795 GND.n6794 0.152939
R21305 GND.n6795 GND.n999 0.152939
R21306 GND.n6803 GND.n999 0.152939
R21307 GND.n6804 GND.n6803 0.152939
R21308 GND.n6805 GND.n6804 0.152939
R21309 GND.n6805 GND.n993 0.152939
R21310 GND.n6813 GND.n993 0.152939
R21311 GND.n6814 GND.n6813 0.152939
R21312 GND.n6815 GND.n6814 0.152939
R21313 GND.n6815 GND.n987 0.152939
R21314 GND.n6823 GND.n987 0.152939
R21315 GND.n6824 GND.n6823 0.152939
R21316 GND.n6825 GND.n6824 0.152939
R21317 GND.n6825 GND.n981 0.152939
R21318 GND.n6833 GND.n981 0.152939
R21319 GND.n6834 GND.n6833 0.152939
R21320 GND.n6835 GND.n6834 0.152939
R21321 GND.n6835 GND.n975 0.152939
R21322 GND.n6843 GND.n975 0.152939
R21323 GND.n6844 GND.n6843 0.152939
R21324 GND.n6845 GND.n6844 0.152939
R21325 GND.n6845 GND.n969 0.152939
R21326 GND.n6853 GND.n969 0.152939
R21327 GND.n6854 GND.n6853 0.152939
R21328 GND.n6855 GND.n6854 0.152939
R21329 GND.n6855 GND.n963 0.152939
R21330 GND.n6863 GND.n963 0.152939
R21331 GND.n6864 GND.n6863 0.152939
R21332 GND.n6865 GND.n6864 0.152939
R21333 GND.n6865 GND.n957 0.152939
R21334 GND.n6873 GND.n957 0.152939
R21335 GND.n6874 GND.n6873 0.152939
R21336 GND.n6875 GND.n6874 0.152939
R21337 GND.n6875 GND.n951 0.152939
R21338 GND.n6883 GND.n951 0.152939
R21339 GND.n6884 GND.n6883 0.152939
R21340 GND.n6885 GND.n6884 0.152939
R21341 GND.n6885 GND.n945 0.152939
R21342 GND.n6893 GND.n945 0.152939
R21343 GND.n6894 GND.n6893 0.152939
R21344 GND.n6895 GND.n6894 0.152939
R21345 GND.n6895 GND.n939 0.152939
R21346 GND.n6903 GND.n939 0.152939
R21347 GND.n6904 GND.n6903 0.152939
R21348 GND.n6905 GND.n6904 0.152939
R21349 GND.n6905 GND.n933 0.152939
R21350 GND.n6913 GND.n933 0.152939
R21351 GND.n6914 GND.n6913 0.152939
R21352 GND.n6915 GND.n6914 0.152939
R21353 GND.n6915 GND.n927 0.152939
R21354 GND.n6923 GND.n927 0.152939
R21355 GND.n6924 GND.n6923 0.152939
R21356 GND.n6925 GND.n6924 0.152939
R21357 GND.n6925 GND.n921 0.152939
R21358 GND.n6933 GND.n921 0.152939
R21359 GND.n6934 GND.n6933 0.152939
R21360 GND.n6935 GND.n6934 0.152939
R21361 GND.n6935 GND.n915 0.152939
R21362 GND.n6943 GND.n915 0.152939
R21363 GND.n6944 GND.n6943 0.152939
R21364 GND.n6945 GND.n6944 0.152939
R21365 GND.n6945 GND.n909 0.152939
R21366 GND.n6953 GND.n909 0.152939
R21367 GND.n6954 GND.n6953 0.152939
R21368 GND.n6955 GND.n6954 0.152939
R21369 GND.n6955 GND.n903 0.152939
R21370 GND.n6963 GND.n903 0.152939
R21371 GND.n6964 GND.n6963 0.152939
R21372 GND.n6965 GND.n6964 0.152939
R21373 GND.n6965 GND.n897 0.152939
R21374 GND.n6973 GND.n897 0.152939
R21375 GND.n6974 GND.n6973 0.152939
R21376 GND.n6975 GND.n6974 0.152939
R21377 GND.n6975 GND.n891 0.152939
R21378 GND.n6983 GND.n891 0.152939
R21379 GND.n6984 GND.n6983 0.152939
R21380 GND.n6985 GND.n6984 0.152939
R21381 GND.n6985 GND.n885 0.152939
R21382 GND.n6993 GND.n885 0.152939
R21383 GND.n6994 GND.n6993 0.152939
R21384 GND.n6995 GND.n6994 0.152939
R21385 GND.n6995 GND.n879 0.152939
R21386 GND.n7003 GND.n879 0.152939
R21387 GND.n7004 GND.n7003 0.152939
R21388 GND.n7005 GND.n7004 0.152939
R21389 GND.n7005 GND.n873 0.152939
R21390 GND.n7013 GND.n873 0.152939
R21391 GND.n7014 GND.n7013 0.152939
R21392 GND.n7015 GND.n7014 0.152939
R21393 GND.n7015 GND.n867 0.152939
R21394 GND.n7023 GND.n867 0.152939
R21395 GND.n7024 GND.n7023 0.152939
R21396 GND.n7025 GND.n7024 0.152939
R21397 GND.n7025 GND.n861 0.152939
R21398 GND.n7033 GND.n861 0.152939
R21399 GND.n7034 GND.n7033 0.152939
R21400 GND.n7035 GND.n7034 0.152939
R21401 GND.n7035 GND.n855 0.152939
R21402 GND.n7043 GND.n855 0.152939
R21403 GND.n7044 GND.n7043 0.152939
R21404 GND.n7045 GND.n7044 0.152939
R21405 GND.n7045 GND.n849 0.152939
R21406 GND.n7053 GND.n849 0.152939
R21407 GND.n7054 GND.n7053 0.152939
R21408 GND.n7055 GND.n7054 0.152939
R21409 GND.n7055 GND.n843 0.152939
R21410 GND.n7063 GND.n843 0.152939
R21411 GND.n7064 GND.n7063 0.152939
R21412 GND.n7065 GND.n7064 0.152939
R21413 GND.n7065 GND.n837 0.152939
R21414 GND.n7073 GND.n837 0.152939
R21415 GND.n7074 GND.n7073 0.152939
R21416 GND.n7075 GND.n7074 0.152939
R21417 GND.n7075 GND.n831 0.152939
R21418 GND.n7083 GND.n831 0.152939
R21419 GND.n7084 GND.n7083 0.152939
R21420 GND.n7085 GND.n7084 0.152939
R21421 GND.n7085 GND.n825 0.152939
R21422 GND.n7093 GND.n825 0.152939
R21423 GND.n7094 GND.n7093 0.152939
R21424 GND.n7095 GND.n7094 0.152939
R21425 GND.n7095 GND.n819 0.152939
R21426 GND.n7103 GND.n819 0.152939
R21427 GND.n7104 GND.n7103 0.152939
R21428 GND.n7105 GND.n7104 0.152939
R21429 GND.n7105 GND.n813 0.152939
R21430 GND.n7113 GND.n813 0.152939
R21431 GND.n7114 GND.n7113 0.152939
R21432 GND.n7115 GND.n7114 0.152939
R21433 GND.n7115 GND.n807 0.152939
R21434 GND.n7123 GND.n807 0.152939
R21435 GND.n7124 GND.n7123 0.152939
R21436 GND.n7125 GND.n7124 0.152939
R21437 GND.n7125 GND.n801 0.152939
R21438 GND.n7133 GND.n801 0.152939
R21439 GND.n7134 GND.n7133 0.152939
R21440 GND.n7135 GND.n7134 0.152939
R21441 GND.n7135 GND.n795 0.152939
R21442 GND.n7143 GND.n795 0.152939
R21443 GND.n7144 GND.n7143 0.152939
R21444 GND.n7145 GND.n7144 0.152939
R21445 GND.n7145 GND.n789 0.152939
R21446 GND.n7153 GND.n789 0.152939
R21447 GND.n7154 GND.n7153 0.152939
R21448 GND.n7155 GND.n7154 0.152939
R21449 GND.n7155 GND.n783 0.152939
R21450 GND.n7163 GND.n783 0.152939
R21451 GND.n7164 GND.n7163 0.152939
R21452 GND.n7165 GND.n7164 0.152939
R21453 GND.n7165 GND.n777 0.152939
R21454 GND.n7173 GND.n777 0.152939
R21455 GND.n7174 GND.n7173 0.152939
R21456 GND.n7175 GND.n7174 0.152939
R21457 GND.n7175 GND.n771 0.152939
R21458 GND.n7183 GND.n771 0.152939
R21459 GND.n7184 GND.n7183 0.152939
R21460 GND.n7185 GND.n7184 0.152939
R21461 GND.n7185 GND.n765 0.152939
R21462 GND.n7193 GND.n765 0.152939
R21463 GND.n7194 GND.n7193 0.152939
R21464 GND.n7195 GND.n7194 0.152939
R21465 GND.n7195 GND.n759 0.152939
R21466 GND.n7203 GND.n759 0.152939
R21467 GND.n7204 GND.n7203 0.152939
R21468 GND.n7205 GND.n7204 0.152939
R21469 GND.n7205 GND.n753 0.152939
R21470 GND.n7213 GND.n753 0.152939
R21471 GND.n7214 GND.n7213 0.152939
R21472 GND.n7215 GND.n7214 0.152939
R21473 GND.n7215 GND.n747 0.152939
R21474 GND.n7223 GND.n747 0.152939
R21475 GND.n7224 GND.n7223 0.152939
R21476 GND.n7225 GND.n7224 0.152939
R21477 GND.n7225 GND.n741 0.152939
R21478 GND.n7233 GND.n741 0.152939
R21479 GND.n7234 GND.n7233 0.152939
R21480 GND.n7235 GND.n7234 0.152939
R21481 GND.n7235 GND.n735 0.152939
R21482 GND.n7243 GND.n735 0.152939
R21483 GND.n7244 GND.n7243 0.152939
R21484 GND.n7245 GND.n7244 0.152939
R21485 GND.n7245 GND.n729 0.152939
R21486 GND.n7253 GND.n729 0.152939
R21487 GND.n7254 GND.n7253 0.152939
R21488 GND.n7255 GND.n7254 0.152939
R21489 GND.n7255 GND.n723 0.152939
R21490 GND.n7263 GND.n723 0.152939
R21491 GND.n7264 GND.n7263 0.152939
R21492 GND.n7265 GND.n7264 0.152939
R21493 GND.n7265 GND.n717 0.152939
R21494 GND.n7273 GND.n717 0.152939
R21495 GND.n7274 GND.n7273 0.152939
R21496 GND.n7275 GND.n7274 0.152939
R21497 GND.n7275 GND.n711 0.152939
R21498 GND.n7283 GND.n711 0.152939
R21499 GND.n7284 GND.n7283 0.152939
R21500 GND.n7285 GND.n7284 0.152939
R21501 GND.n7285 GND.n705 0.152939
R21502 GND.n7293 GND.n705 0.152939
R21503 GND.n7294 GND.n7293 0.152939
R21504 GND.n7295 GND.n7294 0.152939
R21505 GND.n7295 GND.n699 0.152939
R21506 GND.n7303 GND.n699 0.152939
R21507 GND.n7304 GND.n7303 0.152939
R21508 GND.n7305 GND.n7304 0.152939
R21509 GND.n7305 GND.n693 0.152939
R21510 GND.n7313 GND.n693 0.152939
R21511 GND.n7314 GND.n7313 0.152939
R21512 GND.n7315 GND.n7314 0.152939
R21513 GND.n7315 GND.n687 0.152939
R21514 GND.n7323 GND.n687 0.152939
R21515 GND.n7324 GND.n7323 0.152939
R21516 GND.n7326 GND.n7324 0.152939
R21517 GND.n7326 GND.n7325 0.152939
R21518 GND.n7325 GND.n681 0.152939
R21519 GND.n7335 GND.n681 0.152939
R21520 GND.n7336 GND.n676 0.152939
R21521 GND.n7344 GND.n676 0.152939
R21522 GND.n7345 GND.n7344 0.152939
R21523 GND.n7346 GND.n7345 0.152939
R21524 GND.n7346 GND.n670 0.152939
R21525 GND.n7354 GND.n670 0.152939
R21526 GND.n7355 GND.n7354 0.152939
R21527 GND.n7356 GND.n7355 0.152939
R21528 GND.n7356 GND.n664 0.152939
R21529 GND.n7364 GND.n664 0.152939
R21530 GND.n7365 GND.n7364 0.152939
R21531 GND.n7366 GND.n7365 0.152939
R21532 GND.n7366 GND.n658 0.152939
R21533 GND.n7374 GND.n658 0.152939
R21534 GND.n7375 GND.n7374 0.152939
R21535 GND.n7376 GND.n7375 0.152939
R21536 GND.n7376 GND.n652 0.152939
R21537 GND.n7384 GND.n652 0.152939
R21538 GND.n7385 GND.n7384 0.152939
R21539 GND.n7386 GND.n7385 0.152939
R21540 GND.n7386 GND.n646 0.152939
R21541 GND.n7394 GND.n646 0.152939
R21542 GND.n7395 GND.n7394 0.152939
R21543 GND.n7396 GND.n7395 0.152939
R21544 GND.n7396 GND.n640 0.152939
R21545 GND.n7404 GND.n640 0.152939
R21546 GND.n7405 GND.n7404 0.152939
R21547 GND.n7406 GND.n7405 0.152939
R21548 GND.n7406 GND.n634 0.152939
R21549 GND.n7414 GND.n634 0.152939
R21550 GND.n7415 GND.n7414 0.152939
R21551 GND.n7416 GND.n7415 0.152939
R21552 GND.n7416 GND.n628 0.152939
R21553 GND.n7424 GND.n628 0.152939
R21554 GND.n7425 GND.n7424 0.152939
R21555 GND.n7426 GND.n7425 0.152939
R21556 GND.n7426 GND.n622 0.152939
R21557 GND.n7434 GND.n622 0.152939
R21558 GND.n7435 GND.n7434 0.152939
R21559 GND.n7436 GND.n7435 0.152939
R21560 GND.n7436 GND.n616 0.152939
R21561 GND.n7444 GND.n616 0.152939
R21562 GND.n7445 GND.n7444 0.152939
R21563 GND.n7446 GND.n7445 0.152939
R21564 GND.n7446 GND.n610 0.152939
R21565 GND.n7454 GND.n610 0.152939
R21566 GND.n7455 GND.n7454 0.152939
R21567 GND.n7456 GND.n7455 0.152939
R21568 GND.n7456 GND.n604 0.152939
R21569 GND.n7464 GND.n604 0.152939
R21570 GND.n7465 GND.n7464 0.152939
R21571 GND.n7466 GND.n7465 0.152939
R21572 GND.n7466 GND.n598 0.152939
R21573 GND.n7474 GND.n598 0.152939
R21574 GND.n7475 GND.n7474 0.152939
R21575 GND.n7476 GND.n7475 0.152939
R21576 GND.n7476 GND.n592 0.152939
R21577 GND.n7484 GND.n592 0.152939
R21578 GND.n7485 GND.n7484 0.152939
R21579 GND.n7486 GND.n7485 0.152939
R21580 GND.n7486 GND.n586 0.152939
R21581 GND.n7494 GND.n586 0.152939
R21582 GND.n7495 GND.n7494 0.152939
R21583 GND.n7496 GND.n7495 0.152939
R21584 GND.n7496 GND.n580 0.152939
R21585 GND.n7504 GND.n580 0.152939
R21586 GND.n7505 GND.n7504 0.152939
R21587 GND.n7506 GND.n7505 0.152939
R21588 GND.n7506 GND.n574 0.152939
R21589 GND.n7514 GND.n574 0.152939
R21590 GND.n7515 GND.n7514 0.152939
R21591 GND.n7516 GND.n7515 0.152939
R21592 GND.n7516 GND.n568 0.152939
R21593 GND.n7524 GND.n568 0.152939
R21594 GND.n7525 GND.n7524 0.152939
R21595 GND.n7526 GND.n7525 0.152939
R21596 GND.n7526 GND.n562 0.152939
R21597 GND.n7534 GND.n562 0.152939
R21598 GND.n7535 GND.n7534 0.152939
R21599 GND.n7536 GND.n7535 0.152939
R21600 GND.n7536 GND.n556 0.152939
R21601 GND.n7544 GND.n556 0.152939
R21602 GND.n7545 GND.n7544 0.152939
R21603 GND.n7546 GND.n7545 0.152939
R21604 GND.n7546 GND.n550 0.152939
R21605 GND.n7554 GND.n550 0.152939
R21606 GND.n7555 GND.n7554 0.152939
R21607 GND.n7556 GND.n7555 0.152939
R21608 GND.n7557 GND.n7556 0.152939
R21609 GND.n2767 GND.n2766 0.152939
R21610 GND.n2770 GND.n2767 0.152939
R21611 GND.n2771 GND.n2770 0.152939
R21612 GND.n2772 GND.n2771 0.152939
R21613 GND.n2773 GND.n2772 0.152939
R21614 GND.n2776 GND.n2773 0.152939
R21615 GND.n2777 GND.n2776 0.152939
R21616 GND.n2778 GND.n2777 0.152939
R21617 GND.n2779 GND.n2778 0.152939
R21618 GND.n2782 GND.n2779 0.152939
R21619 GND.n2783 GND.n2782 0.152939
R21620 GND.n2784 GND.n2783 0.152939
R21621 GND.n2785 GND.n2784 0.152939
R21622 GND.n5182 GND.n2785 0.152939
R21623 GND.n5183 GND.n5182 0.152939
R21624 GND.n5184 GND.n5183 0.152939
R21625 GND.n5185 GND.n5184 0.152939
R21626 GND.n5188 GND.n5185 0.152939
R21627 GND.n5189 GND.n5188 0.152939
R21628 GND.n5190 GND.n5189 0.152939
R21629 GND.n5191 GND.n5190 0.152939
R21630 GND.n5193 GND.n5191 0.152939
R21631 GND.n5193 GND.n5192 0.152939
R21632 GND.n5192 GND.n186 0.152939
R21633 GND.n187 GND.n186 0.152939
R21634 GND.n188 GND.n187 0.152939
R21635 GND.n382 GND.n188 0.152939
R21636 GND.n383 GND.n382 0.152939
R21637 GND.n384 GND.n383 0.152939
R21638 GND.n385 GND.n384 0.152939
R21639 GND.n390 GND.n385 0.152939
R21640 GND.n391 GND.n390 0.152939
R21641 GND.n392 GND.n391 0.152939
R21642 GND.n393 GND.n392 0.152939
R21643 GND.n398 GND.n393 0.152939
R21644 GND.n399 GND.n398 0.152939
R21645 GND.n400 GND.n399 0.152939
R21646 GND.n401 GND.n400 0.152939
R21647 GND.n406 GND.n401 0.152939
R21648 GND.n407 GND.n406 0.152939
R21649 GND.n408 GND.n407 0.152939
R21650 GND.n409 GND.n408 0.152939
R21651 GND.n414 GND.n409 0.152939
R21652 GND.n415 GND.n414 0.152939
R21653 GND.n416 GND.n415 0.152939
R21654 GND.n417 GND.n416 0.152939
R21655 GND.n422 GND.n417 0.152939
R21656 GND.n423 GND.n422 0.152939
R21657 GND.n424 GND.n423 0.152939
R21658 GND.n425 GND.n424 0.152939
R21659 GND.n430 GND.n425 0.152939
R21660 GND.n431 GND.n430 0.152939
R21661 GND.n432 GND.n431 0.152939
R21662 GND.n433 GND.n432 0.152939
R21663 GND.n438 GND.n433 0.152939
R21664 GND.n439 GND.n438 0.152939
R21665 GND.n440 GND.n439 0.152939
R21666 GND.n441 GND.n440 0.152939
R21667 GND.n446 GND.n441 0.152939
R21668 GND.n447 GND.n446 0.152939
R21669 GND.n448 GND.n447 0.152939
R21670 GND.n449 GND.n448 0.152939
R21671 GND.n454 GND.n449 0.152939
R21672 GND.n455 GND.n454 0.152939
R21673 GND.n456 GND.n455 0.152939
R21674 GND.n457 GND.n456 0.152939
R21675 GND.n462 GND.n457 0.152939
R21676 GND.n463 GND.n462 0.152939
R21677 GND.n464 GND.n463 0.152939
R21678 GND.n465 GND.n464 0.152939
R21679 GND.n470 GND.n465 0.152939
R21680 GND.n471 GND.n470 0.152939
R21681 GND.n472 GND.n471 0.152939
R21682 GND.n473 GND.n472 0.152939
R21683 GND.n478 GND.n473 0.152939
R21684 GND.n479 GND.n478 0.152939
R21685 GND.n480 GND.n479 0.152939
R21686 GND.n481 GND.n480 0.152939
R21687 GND.n486 GND.n481 0.152939
R21688 GND.n487 GND.n486 0.152939
R21689 GND.n488 GND.n487 0.152939
R21690 GND.n489 GND.n488 0.152939
R21691 GND.n494 GND.n489 0.152939
R21692 GND.n495 GND.n494 0.152939
R21693 GND.n496 GND.n495 0.152939
R21694 GND.n497 GND.n496 0.152939
R21695 GND.n502 GND.n497 0.152939
R21696 GND.n503 GND.n502 0.152939
R21697 GND.n504 GND.n503 0.152939
R21698 GND.n505 GND.n504 0.152939
R21699 GND.n510 GND.n505 0.152939
R21700 GND.n511 GND.n510 0.152939
R21701 GND.n512 GND.n511 0.152939
R21702 GND.n513 GND.n512 0.152939
R21703 GND.n518 GND.n513 0.152939
R21704 GND.n519 GND.n518 0.152939
R21705 GND.n520 GND.n519 0.152939
R21706 GND.n521 GND.n520 0.152939
R21707 GND.n526 GND.n521 0.152939
R21708 GND.n527 GND.n526 0.152939
R21709 GND.n528 GND.n527 0.152939
R21710 GND.n529 GND.n528 0.152939
R21711 GND.n534 GND.n529 0.152939
R21712 GND.n535 GND.n534 0.152939
R21713 GND.n536 GND.n535 0.152939
R21714 GND.n537 GND.n536 0.152939
R21715 GND.n542 GND.n537 0.152939
R21716 GND.n543 GND.n542 0.152939
R21717 GND.n544 GND.n543 0.152939
R21718 GND.n545 GND.n544 0.152939
R21719 GND.n63 GND.n36 0.152939
R21720 GND.n64 GND.n63 0.152939
R21721 GND.n65 GND.n64 0.152939
R21722 GND.n83 GND.n65 0.152939
R21723 GND.n84 GND.n83 0.152939
R21724 GND.n85 GND.n84 0.152939
R21725 GND.n86 GND.n85 0.152939
R21726 GND.n104 GND.n86 0.152939
R21727 GND.n105 GND.n104 0.152939
R21728 GND.n106 GND.n105 0.152939
R21729 GND.n107 GND.n106 0.152939
R21730 GND.n125 GND.n107 0.152939
R21731 GND.n126 GND.n125 0.152939
R21732 GND.n127 GND.n126 0.152939
R21733 GND.n128 GND.n127 0.152939
R21734 GND.n145 GND.n128 0.152939
R21735 GND.n146 GND.n145 0.152939
R21736 GND.n147 GND.n146 0.152939
R21737 GND.n148 GND.n147 0.152939
R21738 GND.n166 GND.n148 0.152939
R21739 GND.n167 GND.n166 0.152939
R21740 GND.n168 GND.n167 0.152939
R21741 GND.n169 GND.n168 0.152939
R21742 GND.n217 GND.n169 0.152939
R21743 GND.n4262 GND.n1743 0.152939
R21744 GND.n4263 GND.n4262 0.152939
R21745 GND.n4264 GND.n4263 0.152939
R21746 GND.n4265 GND.n4264 0.152939
R21747 GND.n4266 GND.n4265 0.152939
R21748 GND.n4266 GND.n3060 0.152939
R21749 GND.n4300 GND.n3060 0.152939
R21750 GND.n4301 GND.n4300 0.152939
R21751 GND.n4302 GND.n4301 0.152939
R21752 GND.n4303 GND.n4302 0.152939
R21753 GND.n4304 GND.n4303 0.152939
R21754 GND.n4307 GND.n4304 0.152939
R21755 GND.n4308 GND.n4307 0.152939
R21756 GND.n4310 GND.n4308 0.152939
R21757 GND.n4310 GND.n4309 0.152939
R21758 GND.n4309 GND.n3046 0.152939
R21759 GND.n4421 GND.n3046 0.152939
R21760 GND.n4422 GND.n4421 0.152939
R21761 GND.n4423 GND.n4422 0.152939
R21762 GND.n4423 GND.n3042 0.152939
R21763 GND.n4429 GND.n3042 0.152939
R21764 GND.n4430 GND.n4429 0.152939
R21765 GND.n4431 GND.n4430 0.152939
R21766 GND.n4432 GND.n4431 0.152939
R21767 GND.n4433 GND.n4432 0.152939
R21768 GND.n4435 GND.n4433 0.152939
R21769 GND.n4435 GND.n4434 0.152939
R21770 GND.n4434 GND.n3013 0.152939
R21771 GND.n4465 GND.n3013 0.152939
R21772 GND.n4466 GND.n4465 0.152939
R21773 GND.n4467 GND.n4466 0.152939
R21774 GND.n4468 GND.n4467 0.152939
R21775 GND.n4469 GND.n4468 0.152939
R21776 GND.n4470 GND.n4469 0.152939
R21777 GND.n4471 GND.n4470 0.152939
R21778 GND.n4472 GND.n4471 0.152939
R21779 GND.n4473 GND.n4472 0.152939
R21780 GND.n4473 GND.n2992 0.152939
R21781 GND.n4537 GND.n2992 0.152939
R21782 GND.n4538 GND.n4537 0.152939
R21783 GND.n4539 GND.n4538 0.152939
R21784 GND.n4540 GND.n4539 0.152939
R21785 GND.n4540 GND.n2985 0.152939
R21786 GND.n4565 GND.n2985 0.152939
R21787 GND.n4566 GND.n4565 0.152939
R21788 GND.n4567 GND.n4566 0.152939
R21789 GND.n4567 GND.n2981 0.152939
R21790 GND.n4573 GND.n2981 0.152939
R21791 GND.n4574 GND.n4573 0.152939
R21792 GND.n4575 GND.n4574 0.152939
R21793 GND.n4575 GND.n2977 0.152939
R21794 GND.n4634 GND.n2977 0.152939
R21795 GND.n4635 GND.n4634 0.152939
R21796 GND.n4637 GND.n4635 0.152939
R21797 GND.n4637 GND.n4636 0.152939
R21798 GND.n4636 GND.n2967 0.152939
R21799 GND.n2967 GND.n2965 0.152939
R21800 GND.n4680 GND.n2965 0.152939
R21801 GND.n4681 GND.n4680 0.152939
R21802 GND.n4682 GND.n4681 0.152939
R21803 GND.n4682 GND.n2955 0.152939
R21804 GND.n4697 GND.n2955 0.152939
R21805 GND.n4698 GND.n4697 0.152939
R21806 GND.n4699 GND.n4698 0.152939
R21807 GND.n4699 GND.n2949 0.152939
R21808 GND.n4741 GND.n2949 0.152939
R21809 GND.n4742 GND.n4741 0.152939
R21810 GND.n4743 GND.n4742 0.152939
R21811 GND.n4744 GND.n4743 0.152939
R21812 GND.n4746 GND.n4744 0.152939
R21813 GND.n4746 GND.n4745 0.152939
R21814 GND.n4745 GND.n2932 0.152939
R21815 GND.n4796 GND.n2932 0.152939
R21816 GND.n4797 GND.n4796 0.152939
R21817 GND.n4251 GND.n3082 0.152939
R21818 GND.n3085 GND.n3082 0.152939
R21819 GND.n3086 GND.n3085 0.152939
R21820 GND.n3087 GND.n3086 0.152939
R21821 GND.n3090 GND.n3087 0.152939
R21822 GND.n3091 GND.n3090 0.152939
R21823 GND.n3092 GND.n3091 0.152939
R21824 GND.n3093 GND.n3092 0.152939
R21825 GND.n3097 GND.n3093 0.152939
R21826 GND.n4229 GND.n3097 0.152939
R21827 GND.n4253 GND.n4252 0.152939
R21828 GND.n4252 GND.n1976 0.152939
R21829 GND.n1977 GND.n1976 0.152939
R21830 GND.n1978 GND.n1977 0.152939
R21831 GND.n3064 GND.n1978 0.152939
R21832 GND.n3066 GND.n3064 0.152939
R21833 GND.n3066 GND.n3065 0.152939
R21834 GND.n3065 GND.n2022 0.152939
R21835 GND.n2023 GND.n2022 0.152939
R21836 GND.n2024 GND.n2023 0.152939
R21837 GND.n2067 GND.n2024 0.152939
R21838 GND.n2068 GND.n2067 0.152939
R21839 GND.n2073 GND.n2068 0.152939
R21840 GND.n2074 GND.n2073 0.152939
R21841 GND.n2075 GND.n2074 0.152939
R21842 GND.n2076 GND.n2075 0.152939
R21843 GND.n2077 GND.n2076 0.152939
R21844 GND.n3027 GND.n2077 0.152939
R21845 GND.n3028 GND.n3027 0.152939
R21846 GND.n3028 GND.n3025 0.152939
R21847 GND.n3034 GND.n3025 0.152939
R21848 GND.n3035 GND.n3034 0.152939
R21849 GND.n3036 GND.n3035 0.152939
R21850 GND.n3036 GND.n3021 0.152939
R21851 GND.n4447 GND.n3021 0.152939
R21852 GND.n4448 GND.n4447 0.152939
R21853 GND.n4449 GND.n4448 0.152939
R21854 GND.n4450 GND.n4449 0.152939
R21855 GND.n4451 GND.n4450 0.152939
R21856 GND.n4453 GND.n4451 0.152939
R21857 GND.n4453 GND.n4452 0.152939
R21858 GND.n4452 GND.n3006 0.152939
R21859 GND.n4492 GND.n3006 0.152939
R21860 GND.n4493 GND.n4492 0.152939
R21861 GND.n4494 GND.n4493 0.152939
R21862 GND.n4495 GND.n4494 0.152939
R21863 GND.n4496 GND.n4495 0.152939
R21864 GND.n4498 GND.n4496 0.152939
R21865 GND.n4498 GND.n4497 0.152939
R21866 GND.n4497 GND.n2191 0.152939
R21867 GND.n2192 GND.n2191 0.152939
R21868 GND.n2193 GND.n2192 0.152939
R21869 GND.n4603 GND.n2193 0.152939
R21870 GND.n4606 GND.n4603 0.152939
R21871 GND.n4607 GND.n4606 0.152939
R21872 GND.n4608 GND.n4607 0.152939
R21873 GND.n4608 GND.n4599 0.152939
R21874 GND.n4614 GND.n4599 0.152939
R21875 GND.n4615 GND.n4614 0.152939
R21876 GND.n4616 GND.n4615 0.152939
R21877 GND.n4617 GND.n4616 0.152939
R21878 GND.n4618 GND.n4617 0.152939
R21879 GND.n4620 GND.n4618 0.152939
R21880 GND.n4620 GND.n4619 0.152939
R21881 GND.n4619 GND.n2275 0.152939
R21882 GND.n2276 GND.n2275 0.152939
R21883 GND.n2277 GND.n2276 0.152939
R21884 GND.n2311 GND.n2277 0.152939
R21885 GND.n2314 GND.n2311 0.152939
R21886 GND.n2315 GND.n2314 0.152939
R21887 GND.n2316 GND.n2315 0.152939
R21888 GND.n2317 GND.n2316 0.152939
R21889 GND.n2318 GND.n2317 0.152939
R21890 GND.n2335 GND.n2318 0.152939
R21891 GND.n2336 GND.n2335 0.152939
R21892 GND.n2337 GND.n2336 0.152939
R21893 GND.n2338 GND.n2337 0.152939
R21894 GND.n2355 GND.n2338 0.152939
R21895 GND.n2356 GND.n2355 0.152939
R21896 GND.n2357 GND.n2356 0.152939
R21897 GND.n2358 GND.n2357 0.152939
R21898 GND.n2373 GND.n2358 0.152939
R21899 GND.n2374 GND.n2373 0.152939
R21900 GND.n5525 GND.n2374 0.152939
R21901 GND.n5524 GND.n2375 0.152939
R21902 GND.n2390 GND.n2375 0.152939
R21903 GND.n2391 GND.n2390 0.152939
R21904 GND.n2392 GND.n2391 0.152939
R21905 GND.n2393 GND.n2392 0.152939
R21906 GND.n2394 GND.n2393 0.152939
R21907 GND.n2395 GND.n2394 0.152939
R21908 GND.n2396 GND.n2395 0.152939
R21909 GND.n2397 GND.n2396 0.152939
R21910 GND.n2398 GND.n2397 0.152939
R21911 GND.n2896 GND.n2895 0.152939
R21912 GND.n4914 GND.n2895 0.152939
R21913 GND.n4915 GND.n4914 0.152939
R21914 GND.n4916 GND.n4915 0.152939
R21915 GND.n4916 GND.n2893 0.152939
R21916 GND.n4938 GND.n2893 0.152939
R21917 GND.n4939 GND.n4938 0.152939
R21918 GND.n4940 GND.n4939 0.152939
R21919 GND.n4940 GND.n2829 0.152939
R21920 GND.n4953 GND.n2829 0.152939
R21921 GND.n4954 GND.n4953 0.152939
R21922 GND.n4955 GND.n4954 0.152939
R21923 GND.n4955 GND.n2825 0.152939
R21924 GND.n4968 GND.n2825 0.152939
R21925 GND.n4969 GND.n4968 0.152939
R21926 GND.n4970 GND.n4969 0.152939
R21927 GND.n4970 GND.n2821 0.152939
R21928 GND.n4983 GND.n2821 0.152939
R21929 GND.n4984 GND.n4983 0.152939
R21930 GND.n4985 GND.n4984 0.152939
R21931 GND.n4985 GND.n2817 0.152939
R21932 GND.n4998 GND.n2817 0.152939
R21933 GND.n4999 GND.n4998 0.152939
R21934 GND.n5000 GND.n4999 0.152939
R21935 GND.n5001 GND.n5000 0.152939
R21936 GND.n5002 GND.n5001 0.152939
R21937 GND.n5003 GND.n5002 0.152939
R21938 GND.n5004 GND.n5003 0.152939
R21939 GND.n5004 GND.n22 0.152939
R21940 GND.n7827 GND.n23 0.152939
R21941 GND.n5036 GND.n23 0.152939
R21942 GND.n5037 GND.n5036 0.152939
R21943 GND.n5037 GND.n2811 0.152939
R21944 GND.n5050 GND.n2811 0.152939
R21945 GND.n5051 GND.n5050 0.152939
R21946 GND.n5052 GND.n5051 0.152939
R21947 GND.n5052 GND.n2806 0.152939
R21948 GND.n5064 GND.n2806 0.152939
R21949 GND.n5065 GND.n5064 0.152939
R21950 GND.n5066 GND.n5065 0.152939
R21951 GND.n5066 GND.n2801 0.152939
R21952 GND.n5078 GND.n2801 0.152939
R21953 GND.n5079 GND.n5078 0.152939
R21954 GND.n5080 GND.n5079 0.152939
R21955 GND.n5080 GND.n2796 0.152939
R21956 GND.n5092 GND.n2796 0.152939
R21957 GND.n5093 GND.n5092 0.152939
R21958 GND.n5095 GND.n5093 0.152939
R21959 GND.n5095 GND.n5094 0.152939
R21960 GND.n5094 GND.n2789 0.152939
R21961 GND.n2790 GND.n2789 0.152939
R21962 GND.n2791 GND.n2790 0.152939
R21963 GND.n5106 GND.n2791 0.152939
R21964 GND.n5107 GND.n5106 0.152939
R21965 GND.n5108 GND.n5107 0.152939
R21966 GND.n5109 GND.n5108 0.152939
R21967 GND.n5110 GND.n5109 0.152939
R21968 GND.n5155 GND.n5110 0.152939
R21969 GND.n5127 GND.n5126 0.152939
R21970 GND.n5127 GND.n5121 0.152939
R21971 GND.n5135 GND.n5121 0.152939
R21972 GND.n5136 GND.n5135 0.152939
R21973 GND.n5137 GND.n5136 0.152939
R21974 GND.n5137 GND.n5117 0.152939
R21975 GND.n5145 GND.n5117 0.152939
R21976 GND.n5146 GND.n5145 0.152939
R21977 GND.n5147 GND.n5146 0.152939
R21978 GND.n5147 GND.n5111 0.152939
R21979 GND.n5154 GND.n5111 0.152939
R21980 GND.n375 GND.n218 0.152939
R21981 GND.n375 GND.n374 0.152939
R21982 GND.n374 GND.n373 0.152939
R21983 GND.n373 GND.n220 0.152939
R21984 GND.n221 GND.n220 0.152939
R21985 GND.n222 GND.n221 0.152939
R21986 GND.n223 GND.n222 0.152939
R21987 GND.n224 GND.n223 0.152939
R21988 GND.n225 GND.n224 0.152939
R21989 GND.n226 GND.n225 0.152939
R21990 GND.n230 GND.n226 0.152939
R21991 GND.n231 GND.n230 0.152939
R21992 GND.n232 GND.n231 0.152939
R21993 GND.n233 GND.n232 0.152939
R21994 GND.n234 GND.n233 0.152939
R21995 GND.n235 GND.n234 0.152939
R21996 GND.n236 GND.n235 0.152939
R21997 GND.n237 GND.n236 0.152939
R21998 GND.n238 GND.n237 0.152939
R21999 GND.n239 GND.n238 0.152939
R22000 GND.n240 GND.n239 0.152939
R22001 GND.n241 GND.n240 0.152939
R22002 GND.n242 GND.n241 0.152939
R22003 GND.n243 GND.n242 0.152939
R22004 GND.n244 GND.n243 0.152939
R22005 GND.n245 GND.n244 0.152939
R22006 GND.n246 GND.n245 0.152939
R22007 GND.n247 GND.n246 0.152939
R22008 GND.n248 GND.n247 0.152939
R22009 GND.n249 GND.n248 0.152939
R22010 GND.n250 GND.n249 0.152939
R22011 GND.n251 GND.n250 0.152939
R22012 GND.n252 GND.n251 0.152939
R22013 GND.n253 GND.n252 0.152939
R22014 GND.n254 GND.n253 0.152939
R22015 GND.n301 GND.n254 0.152939
R22016 GND.n301 GND.n300 0.152939
R22017 GND.n300 GND.n299 0.152939
R22018 GND.n299 GND.n260 0.152939
R22019 GND.n261 GND.n260 0.152939
R22020 GND.n262 GND.n261 0.152939
R22021 GND.n263 GND.n262 0.152939
R22022 GND.n264 GND.n263 0.152939
R22023 GND.n265 GND.n264 0.152939
R22024 GND.n266 GND.n265 0.152939
R22025 GND.n267 GND.n266 0.152939
R22026 GND.n268 GND.n267 0.152939
R22027 GND.n269 GND.n268 0.152939
R22028 GND.n274 GND.n269 0.152939
R22029 GND.n274 GND.n273 0.152939
R22030 GND.n5338 GND.n5337 0.152939
R22031 GND.n5339 GND.n5338 0.152939
R22032 GND.n5340 GND.n5339 0.152939
R22033 GND.n5341 GND.n5340 0.152939
R22034 GND.n5342 GND.n5341 0.152939
R22035 GND.n5343 GND.n5342 0.152939
R22036 GND.n5344 GND.n5343 0.152939
R22037 GND.n5345 GND.n5344 0.152939
R22038 GND.n5346 GND.n5345 0.152939
R22039 GND.n5347 GND.n5346 0.152939
R22040 GND.n5351 GND.n5347 0.152939
R22041 GND.n5352 GND.n5351 0.152939
R22042 GND.n5353 GND.n5352 0.152939
R22043 GND.n5354 GND.n5353 0.152939
R22044 GND.n5355 GND.n5354 0.152939
R22045 GND.n5356 GND.n5355 0.152939
R22046 GND.n5357 GND.n5356 0.152939
R22047 GND.n5358 GND.n5357 0.152939
R22048 GND.n5359 GND.n5358 0.152939
R22049 GND.n5361 GND.n5359 0.152939
R22050 GND.n5361 GND.n5360 0.152939
R22051 GND.n4840 GND.n2554 0.152939
R22052 GND.n4841 GND.n4840 0.152939
R22053 GND.n4841 GND.n4839 0.152939
R22054 GND.n4849 GND.n4839 0.152939
R22055 GND.n4850 GND.n4849 0.152939
R22056 GND.n4851 GND.n4850 0.152939
R22057 GND.n4851 GND.n4837 0.152939
R22058 GND.n4859 GND.n4837 0.152939
R22059 GND.n4860 GND.n4859 0.152939
R22060 GND.n4861 GND.n4860 0.152939
R22061 GND.n4861 GND.n4835 0.152939
R22062 GND.n4871 GND.n4835 0.152939
R22063 GND.n4872 GND.n4871 0.152939
R22064 GND.n4873 GND.n4872 0.152939
R22065 GND.n4873 GND.n4833 0.152939
R22066 GND.n4881 GND.n4833 0.152939
R22067 GND.n4882 GND.n4881 0.152939
R22068 GND.n4883 GND.n4882 0.152939
R22069 GND.n4883 GND.n4831 0.152939
R22070 GND.n4891 GND.n4831 0.152939
R22071 GND.n4892 GND.n4891 0.152939
R22072 GND.n4893 GND.n4892 0.152939
R22073 GND.n4893 GND.n4829 0.152939
R22074 GND.n4901 GND.n4829 0.152939
R22075 GND.n4902 GND.n4901 0.152939
R22076 GND.n4905 GND.n4902 0.152939
R22077 GND.n5336 GND.n2591 0.152939
R22078 GND.n2626 GND.n2591 0.152939
R22079 GND.n2629 GND.n2626 0.152939
R22080 GND.n2630 GND.n2629 0.152939
R22081 GND.n2631 GND.n2630 0.152939
R22082 GND.n2632 GND.n2631 0.152939
R22083 GND.n2633 GND.n2632 0.152939
R22084 GND.n2652 GND.n2633 0.152939
R22085 GND.n2653 GND.n2652 0.152939
R22086 GND.n2654 GND.n2653 0.152939
R22087 GND.n2655 GND.n2654 0.152939
R22088 GND.n2673 GND.n2655 0.152939
R22089 GND.n2674 GND.n2673 0.152939
R22090 GND.n2675 GND.n2674 0.152939
R22091 GND.n2676 GND.n2675 0.152939
R22092 GND.n2694 GND.n2676 0.152939
R22093 GND.n2695 GND.n2694 0.152939
R22094 GND.n2696 GND.n2695 0.152939
R22095 GND.n2697 GND.n2696 0.152939
R22096 GND.n2715 GND.n2697 0.152939
R22097 GND.n2716 GND.n2715 0.152939
R22098 GND.n2717 GND.n2716 0.152939
R22099 GND.n2718 GND.n2717 0.152939
R22100 GND.n2718 GND.n37 0.152939
R22101 GND.n3944 GND.n3943 0.152939
R22102 GND.n3944 GND.n3298 0.152939
R22103 GND.n3977 GND.n3298 0.152939
R22104 GND.n3978 GND.n3977 0.152939
R22105 GND.n3979 GND.n3978 0.152939
R22106 GND.n3980 GND.n3979 0.152939
R22107 GND.n3980 GND.n3268 0.152939
R22108 GND.n4014 GND.n3268 0.152939
R22109 GND.n4015 GND.n4014 0.152939
R22110 GND.n4016 GND.n4015 0.152939
R22111 GND.n4017 GND.n4016 0.152939
R22112 GND.n4017 GND.n3239 0.152939
R22113 GND.n4051 GND.n3239 0.152939
R22114 GND.n4052 GND.n4051 0.152939
R22115 GND.n4053 GND.n4052 0.152939
R22116 GND.n4054 GND.n4053 0.152939
R22117 GND.n4054 GND.n3210 0.152939
R22118 GND.n4088 GND.n3210 0.152939
R22119 GND.n4089 GND.n4088 0.152939
R22120 GND.n4090 GND.n4089 0.152939
R22121 GND.n4091 GND.n4090 0.152939
R22122 GND.n4092 GND.n4091 0.152939
R22123 GND.n4095 GND.n4092 0.152939
R22124 GND.n4096 GND.n4095 0.152939
R22125 GND.n4097 GND.n4096 0.152939
R22126 GND.n4098 GND.n4097 0.152939
R22127 GND.n4101 GND.n4098 0.152939
R22128 GND.n4102 GND.n4101 0.152939
R22129 GND.n4103 GND.n4102 0.152939
R22130 GND.n4104 GND.n4103 0.152939
R22131 GND.n4106 GND.n4104 0.152939
R22132 GND.n4106 GND.n4105 0.152939
R22133 GND.n4105 GND.n1889 0.152939
R22134 GND.n1890 GND.n1889 0.152939
R22135 GND.n1891 GND.n1890 0.152939
R22136 GND.n1998 GND.n1891 0.152939
R22137 GND.n2001 GND.n1998 0.152939
R22138 GND.n2002 GND.n2001 0.152939
R22139 GND.n2003 GND.n2002 0.152939
R22140 GND.n2003 GND.n1994 0.152939
R22141 GND.n2009 GND.n1994 0.152939
R22142 GND.n2010 GND.n2009 0.152939
R22143 GND.n2011 GND.n2010 0.152939
R22144 GND.n2012 GND.n2011 0.152939
R22145 GND.n2013 GND.n2012 0.152939
R22146 GND.n2042 GND.n2013 0.152939
R22147 GND.n2045 GND.n2042 0.152939
R22148 GND.n2046 GND.n2045 0.152939
R22149 GND.n2047 GND.n2046 0.152939
R22150 GND.n2048 GND.n2047 0.152939
R22151 GND.n2049 GND.n2048 0.152939
R22152 GND.n2086 GND.n2049 0.152939
R22153 GND.n2089 GND.n2086 0.152939
R22154 GND.n2090 GND.n2089 0.152939
R22155 GND.n2091 GND.n2090 0.152939
R22156 GND.n2092 GND.n2091 0.152939
R22157 GND.n2093 GND.n2092 0.152939
R22158 GND.n2108 GND.n2093 0.152939
R22159 GND.n2109 GND.n2108 0.152939
R22160 GND.n2110 GND.n2109 0.152939
R22161 GND.n2111 GND.n2110 0.152939
R22162 GND.n2126 GND.n2111 0.152939
R22163 GND.n2127 GND.n2126 0.152939
R22164 GND.n2128 GND.n2127 0.152939
R22165 GND.n2129 GND.n2128 0.152939
R22166 GND.n2143 GND.n2129 0.152939
R22167 GND.n2144 GND.n2143 0.152939
R22168 GND.n2145 GND.n2144 0.152939
R22169 GND.n2146 GND.n2145 0.152939
R22170 GND.n2161 GND.n2146 0.152939
R22171 GND.n2162 GND.n2161 0.152939
R22172 GND.n2163 GND.n2162 0.152939
R22173 GND.n2164 GND.n2163 0.152939
R22174 GND.n2179 GND.n2164 0.152939
R22175 GND.n2180 GND.n2179 0.152939
R22176 GND.n2181 GND.n2180 0.152939
R22177 GND.n2182 GND.n2181 0.152939
R22178 GND.n2210 GND.n2182 0.152939
R22179 GND.n2213 GND.n2210 0.152939
R22180 GND.n2214 GND.n2213 0.152939
R22181 GND.n2215 GND.n2214 0.152939
R22182 GND.n2216 GND.n2215 0.152939
R22183 GND.n2217 GND.n2216 0.152939
R22184 GND.n2244 GND.n2217 0.152939
R22185 GND.n2245 GND.n2244 0.152939
R22186 GND.n2246 GND.n2245 0.152939
R22187 GND.n2247 GND.n2246 0.152939
R22188 GND.n2248 GND.n2247 0.152939
R22189 GND.n2263 GND.n2248 0.152939
R22190 GND.n2264 GND.n2263 0.152939
R22191 GND.n2265 GND.n2264 0.152939
R22192 GND.n2266 GND.n2265 0.152939
R22193 GND.n2295 GND.n2266 0.152939
R22194 GND.n2298 GND.n2295 0.152939
R22195 GND.n2299 GND.n2298 0.152939
R22196 GND.n2300 GND.n2299 0.152939
R22197 GND.n2301 GND.n2300 0.152939
R22198 GND.n2302 GND.n2301 0.152939
R22199 GND.n4720 GND.n2302 0.152939
R22200 GND.n4721 GND.n4720 0.152939
R22201 GND.n4721 GND.n4718 0.152939
R22202 GND.n4727 GND.n4718 0.152939
R22203 GND.n4728 GND.n4727 0.152939
R22204 GND.n4729 GND.n4728 0.152939
R22205 GND.n4730 GND.n4729 0.152939
R22206 GND.n4731 GND.n4730 0.152939
R22207 GND.n4731 GND.n2938 0.152939
R22208 GND.n4772 GND.n2938 0.152939
R22209 GND.n4773 GND.n4772 0.152939
R22210 GND.n4774 GND.n4773 0.152939
R22211 GND.n4775 GND.n4774 0.152939
R22212 GND.n4776 GND.n4775 0.152939
R22213 GND.n4778 GND.n4776 0.152939
R22214 GND.n4780 GND.n4778 0.152939
R22215 GND.n4780 GND.n4779 0.152939
R22216 GND.n4779 GND.n2438 0.152939
R22217 GND.n2439 GND.n2438 0.152939
R22218 GND.n2440 GND.n2439 0.152939
R22219 GND.n4807 GND.n2440 0.152939
R22220 GND.n4808 GND.n4807 0.152939
R22221 GND.n4808 GND.n4805 0.152939
R22222 GND.n4817 GND.n4805 0.152939
R22223 GND.n4818 GND.n4817 0.152939
R22224 GND.n4819 GND.n4818 0.152939
R22225 GND.n4821 GND.n4819 0.152939
R22226 GND.n4821 GND.n4820 0.152939
R22227 GND.n4820 GND.n2612 0.152939
R22228 GND.n2613 GND.n2612 0.152939
R22229 GND.n2614 GND.n2613 0.152939
R22230 GND.n2835 GND.n2614 0.152939
R22231 GND.n2836 GND.n2835 0.152939
R22232 GND.n2837 GND.n2836 0.152939
R22233 GND.n2838 GND.n2837 0.152939
R22234 GND.n2839 GND.n2838 0.152939
R22235 GND.n2842 GND.n2839 0.152939
R22236 GND.n2843 GND.n2842 0.152939
R22237 GND.n2844 GND.n2843 0.152939
R22238 GND.n2845 GND.n2844 0.152939
R22239 GND.n2848 GND.n2845 0.152939
R22240 GND.n2849 GND.n2848 0.152939
R22241 GND.n2850 GND.n2849 0.152939
R22242 GND.n2851 GND.n2850 0.152939
R22243 GND.n2854 GND.n2851 0.152939
R22244 GND.n2855 GND.n2854 0.152939
R22245 GND.n2856 GND.n2855 0.152939
R22246 GND.n2857 GND.n2856 0.152939
R22247 GND.n2860 GND.n2857 0.152939
R22248 GND.n2861 GND.n2860 0.152939
R22249 GND.n2862 GND.n2861 0.152939
R22250 GND.n3966 GND.n3308 0.152939
R22251 GND.n3967 GND.n3966 0.152939
R22252 GND.n3968 GND.n3967 0.152939
R22253 GND.n3969 GND.n3968 0.152939
R22254 GND.n3969 GND.n3279 0.152939
R22255 GND.n4003 GND.n3279 0.152939
R22256 GND.n4004 GND.n4003 0.152939
R22257 GND.n4005 GND.n4004 0.152939
R22258 GND.n4006 GND.n4005 0.152939
R22259 GND.n4006 GND.n3250 0.152939
R22260 GND.n4040 GND.n3250 0.152939
R22261 GND.n4041 GND.n4040 0.152939
R22262 GND.n4042 GND.n4041 0.152939
R22263 GND.n4043 GND.n4042 0.152939
R22264 GND.n4043 GND.n3220 0.152939
R22265 GND.n4077 GND.n3220 0.152939
R22266 GND.n4078 GND.n4077 0.152939
R22267 GND.n4079 GND.n4078 0.152939
R22268 GND.n4080 GND.n4079 0.152939
R22269 GND.n4080 GND.n3193 0.152939
R22270 GND.n4143 GND.n3193 0.152939
R22271 GND.n4144 GND.n4143 0.152939
R22272 GND.n4145 GND.n4144 0.152939
R22273 GND.n4145 GND.n1785 0.152939
R22274 GND.n3526 GND.n3482 0.152939
R22275 GND.n3532 GND.n3526 0.152939
R22276 GND.n3533 GND.n3532 0.152939
R22277 GND.n3534 GND.n3533 0.152939
R22278 GND.n3534 GND.n3524 0.152939
R22279 GND.n3542 GND.n3524 0.152939
R22280 GND.n3543 GND.n3542 0.152939
R22281 GND.n3544 GND.n3543 0.152939
R22282 GND.n3544 GND.n3522 0.152939
R22283 GND.n3552 GND.n3522 0.152939
R22284 GND.n3553 GND.n3552 0.152939
R22285 GND.n3553 GND.n3518 0.152939
R22286 GND.n3561 GND.n3518 0.152939
R22287 GND.n3562 GND.n3561 0.152939
R22288 GND.n3563 GND.n3562 0.152939
R22289 GND.n3563 GND.n3516 0.152939
R22290 GND.n3571 GND.n3516 0.152939
R22291 GND.n3572 GND.n3571 0.152939
R22292 GND.n3573 GND.n3572 0.152939
R22293 GND.n3573 GND.n3514 0.152939
R22294 GND.n3581 GND.n3514 0.152939
R22295 GND.n3582 GND.n3581 0.152939
R22296 GND.n3583 GND.n3582 0.152939
R22297 GND.n3583 GND.n3512 0.152939
R22298 GND.n3512 GND.n3508 0.152939
R22299 GND.n3592 GND.n3508 0.152939
R22300 GND.n3593 GND.n3592 0.152939
R22301 GND.n3594 GND.n3593 0.152939
R22302 GND.n3594 GND.n3506 0.152939
R22303 GND.n3602 GND.n3506 0.152939
R22304 GND.n3603 GND.n3602 0.152939
R22305 GND.n3604 GND.n3603 0.152939
R22306 GND.n3604 GND.n3504 0.152939
R22307 GND.n3612 GND.n3504 0.152939
R22308 GND.n3613 GND.n3612 0.152939
R22309 GND.n3614 GND.n3613 0.152939
R22310 GND.n3614 GND.n3500 0.152939
R22311 GND.n3622 GND.n3500 0.152939
R22312 GND.n3623 GND.n3622 0.152939
R22313 GND.n3624 GND.n3623 0.152939
R22314 GND.n3624 GND.n3498 0.152939
R22315 GND.n3632 GND.n3498 0.152939
R22316 GND.n3633 GND.n3632 0.152939
R22317 GND.n3634 GND.n3633 0.152939
R22318 GND.n3634 GND.n3496 0.152939
R22319 GND.n3642 GND.n3496 0.152939
R22320 GND.n3643 GND.n3642 0.152939
R22321 GND.n3644 GND.n3643 0.152939
R22322 GND.n3644 GND.n3494 0.152939
R22323 GND.n3653 GND.n3494 0.152939
R22324 GND.n3673 GND.n3672 0.152939
R22325 GND.n3674 GND.n3673 0.152939
R22326 GND.n3675 GND.n3674 0.152939
R22327 GND.n3675 GND.n3453 0.152939
R22328 GND.n3709 GND.n3453 0.152939
R22329 GND.n3710 GND.n3709 0.152939
R22330 GND.n3711 GND.n3710 0.152939
R22331 GND.n3712 GND.n3711 0.152939
R22332 GND.n3712 GND.n3424 0.152939
R22333 GND.n3746 GND.n3424 0.152939
R22334 GND.n3747 GND.n3746 0.152939
R22335 GND.n3748 GND.n3747 0.152939
R22336 GND.n3749 GND.n3748 0.152939
R22337 GND.n3749 GND.n3394 0.152939
R22338 GND.n3783 GND.n3394 0.152939
R22339 GND.n3784 GND.n3783 0.152939
R22340 GND.n3785 GND.n3784 0.152939
R22341 GND.n3786 GND.n3785 0.152939
R22342 GND.n3786 GND.n3364 0.152939
R22343 GND.n3820 GND.n3364 0.152939
R22344 GND.n3821 GND.n3820 0.152939
R22345 GND.n3823 GND.n3821 0.152939
R22346 GND.n3823 GND.n3822 0.152939
R22347 GND.n3822 GND.n3342 0.152939
R22348 GND.n1450 GND.n1449 0.152939
R22349 GND.n1451 GND.n1450 0.152939
R22350 GND.n1452 GND.n1451 0.152939
R22351 GND.n1457 GND.n1452 0.152939
R22352 GND.n1458 GND.n1457 0.152939
R22353 GND.n1459 GND.n1458 0.152939
R22354 GND.n1460 GND.n1459 0.152939
R22355 GND.n1465 GND.n1460 0.152939
R22356 GND.n1466 GND.n1465 0.152939
R22357 GND.n1467 GND.n1466 0.152939
R22358 GND.n1468 GND.n1467 0.152939
R22359 GND.n1473 GND.n1468 0.152939
R22360 GND.n1474 GND.n1473 0.152939
R22361 GND.n1475 GND.n1474 0.152939
R22362 GND.n1476 GND.n1475 0.152939
R22363 GND.n1481 GND.n1476 0.152939
R22364 GND.n1482 GND.n1481 0.152939
R22365 GND.n1483 GND.n1482 0.152939
R22366 GND.n1484 GND.n1483 0.152939
R22367 GND.n1489 GND.n1484 0.152939
R22368 GND.n1490 GND.n1489 0.152939
R22369 GND.n1491 GND.n1490 0.152939
R22370 GND.n1492 GND.n1491 0.152939
R22371 GND.n1497 GND.n1492 0.152939
R22372 GND.n1498 GND.n1497 0.152939
R22373 GND.n1499 GND.n1498 0.152939
R22374 GND.n1500 GND.n1499 0.152939
R22375 GND.n1505 GND.n1500 0.152939
R22376 GND.n1506 GND.n1505 0.152939
R22377 GND.n1507 GND.n1506 0.152939
R22378 GND.n1508 GND.n1507 0.152939
R22379 GND.n1513 GND.n1508 0.152939
R22380 GND.n1514 GND.n1513 0.152939
R22381 GND.n1515 GND.n1514 0.152939
R22382 GND.n1516 GND.n1515 0.152939
R22383 GND.n1521 GND.n1516 0.152939
R22384 GND.n1522 GND.n1521 0.152939
R22385 GND.n1523 GND.n1522 0.152939
R22386 GND.n1524 GND.n1523 0.152939
R22387 GND.n1529 GND.n1524 0.152939
R22388 GND.n1530 GND.n1529 0.152939
R22389 GND.n1531 GND.n1530 0.152939
R22390 GND.n1532 GND.n1531 0.152939
R22391 GND.n1537 GND.n1532 0.152939
R22392 GND.n1538 GND.n1537 0.152939
R22393 GND.n1539 GND.n1538 0.152939
R22394 GND.n1540 GND.n1539 0.152939
R22395 GND.n1545 GND.n1540 0.152939
R22396 GND.n1546 GND.n1545 0.152939
R22397 GND.n1547 GND.n1546 0.152939
R22398 GND.n1548 GND.n1547 0.152939
R22399 GND.n1553 GND.n1548 0.152939
R22400 GND.n1554 GND.n1553 0.152939
R22401 GND.n1555 GND.n1554 0.152939
R22402 GND.n1556 GND.n1555 0.152939
R22403 GND.n1561 GND.n1556 0.152939
R22404 GND.n1562 GND.n1561 0.152939
R22405 GND.n1563 GND.n1562 0.152939
R22406 GND.n1564 GND.n1563 0.152939
R22407 GND.n1569 GND.n1564 0.152939
R22408 GND.n1570 GND.n1569 0.152939
R22409 GND.n1571 GND.n1570 0.152939
R22410 GND.n1572 GND.n1571 0.152939
R22411 GND.n1577 GND.n1572 0.152939
R22412 GND.n1578 GND.n1577 0.152939
R22413 GND.n1579 GND.n1578 0.152939
R22414 GND.n1580 GND.n1579 0.152939
R22415 GND.n1585 GND.n1580 0.152939
R22416 GND.n1586 GND.n1585 0.152939
R22417 GND.n1587 GND.n1586 0.152939
R22418 GND.n1588 GND.n1587 0.152939
R22419 GND.n1593 GND.n1588 0.152939
R22420 GND.n1594 GND.n1593 0.152939
R22421 GND.n1595 GND.n1594 0.152939
R22422 GND.n1596 GND.n1595 0.152939
R22423 GND.n1601 GND.n1596 0.152939
R22424 GND.n1602 GND.n1601 0.152939
R22425 GND.n1603 GND.n1602 0.152939
R22426 GND.n1604 GND.n1603 0.152939
R22427 GND.n1609 GND.n1604 0.152939
R22428 GND.n1610 GND.n1609 0.152939
R22429 GND.n1611 GND.n1610 0.152939
R22430 GND.n1612 GND.n1611 0.152939
R22431 GND.n3486 GND.n1612 0.152939
R22432 GND.n3487 GND.n3486 0.152939
R22433 GND.n3488 GND.n3487 0.152939
R22434 GND.n3488 GND.n3472 0.152939
R22435 GND.n3683 GND.n3472 0.152939
R22436 GND.n3684 GND.n3683 0.152939
R22437 GND.n3685 GND.n3684 0.152939
R22438 GND.n3686 GND.n3685 0.152939
R22439 GND.n3686 GND.n3442 0.152939
R22440 GND.n3720 GND.n3442 0.152939
R22441 GND.n3721 GND.n3720 0.152939
R22442 GND.n3722 GND.n3721 0.152939
R22443 GND.n3723 GND.n3722 0.152939
R22444 GND.n3723 GND.n3413 0.152939
R22445 GND.n3757 GND.n3413 0.152939
R22446 GND.n3758 GND.n3757 0.152939
R22447 GND.n3759 GND.n3758 0.152939
R22448 GND.n3760 GND.n3759 0.152939
R22449 GND.n3760 GND.n3384 0.152939
R22450 GND.n3794 GND.n3384 0.152939
R22451 GND.n3795 GND.n3794 0.152939
R22452 GND.n3796 GND.n3795 0.152939
R22453 GND.n3797 GND.n3796 0.152939
R22454 GND.n3798 GND.n3797 0.152939
R22455 GND.n3799 GND.n3798 0.152939
R22456 GND.n3799 GND.n3331 0.152939
R22457 GND.n3941 GND.n3331 0.152939
R22458 GND.n6354 GND.n1268 0.152939
R22459 GND.n1273 GND.n1268 0.152939
R22460 GND.n1274 GND.n1273 0.152939
R22461 GND.n1275 GND.n1274 0.152939
R22462 GND.n1276 GND.n1275 0.152939
R22463 GND.n1281 GND.n1276 0.152939
R22464 GND.n1282 GND.n1281 0.152939
R22465 GND.n1283 GND.n1282 0.152939
R22466 GND.n1284 GND.n1283 0.152939
R22467 GND.n1289 GND.n1284 0.152939
R22468 GND.n1290 GND.n1289 0.152939
R22469 GND.n1291 GND.n1290 0.152939
R22470 GND.n1292 GND.n1291 0.152939
R22471 GND.n1297 GND.n1292 0.152939
R22472 GND.n1298 GND.n1297 0.152939
R22473 GND.n1299 GND.n1298 0.152939
R22474 GND.n1300 GND.n1299 0.152939
R22475 GND.n1305 GND.n1300 0.152939
R22476 GND.n1306 GND.n1305 0.152939
R22477 GND.n1307 GND.n1306 0.152939
R22478 GND.n1308 GND.n1307 0.152939
R22479 GND.n1313 GND.n1308 0.152939
R22480 GND.n1314 GND.n1313 0.152939
R22481 GND.n1315 GND.n1314 0.152939
R22482 GND.n1316 GND.n1315 0.152939
R22483 GND.n1321 GND.n1316 0.152939
R22484 GND.n1322 GND.n1321 0.152939
R22485 GND.n1323 GND.n1322 0.152939
R22486 GND.n1324 GND.n1323 0.152939
R22487 GND.n1329 GND.n1324 0.152939
R22488 GND.n1330 GND.n1329 0.152939
R22489 GND.n1331 GND.n1330 0.152939
R22490 GND.n1332 GND.n1331 0.152939
R22491 GND.n1337 GND.n1332 0.152939
R22492 GND.n1338 GND.n1337 0.152939
R22493 GND.n1339 GND.n1338 0.152939
R22494 GND.n1340 GND.n1339 0.152939
R22495 GND.n1345 GND.n1340 0.152939
R22496 GND.n1346 GND.n1345 0.152939
R22497 GND.n1347 GND.n1346 0.152939
R22498 GND.n1348 GND.n1347 0.152939
R22499 GND.n1353 GND.n1348 0.152939
R22500 GND.n1354 GND.n1353 0.152939
R22501 GND.n1355 GND.n1354 0.152939
R22502 GND.n1356 GND.n1355 0.152939
R22503 GND.n1361 GND.n1356 0.152939
R22504 GND.n1362 GND.n1361 0.152939
R22505 GND.n1363 GND.n1362 0.152939
R22506 GND.n1364 GND.n1363 0.152939
R22507 GND.n1369 GND.n1364 0.152939
R22508 GND.n1370 GND.n1369 0.152939
R22509 GND.n1371 GND.n1370 0.152939
R22510 GND.n1372 GND.n1371 0.152939
R22511 GND.n1377 GND.n1372 0.152939
R22512 GND.n1378 GND.n1377 0.152939
R22513 GND.n1379 GND.n1378 0.152939
R22514 GND.n1380 GND.n1379 0.152939
R22515 GND.n1385 GND.n1380 0.152939
R22516 GND.n1386 GND.n1385 0.152939
R22517 GND.n1387 GND.n1386 0.152939
R22518 GND.n1388 GND.n1387 0.152939
R22519 GND.n1393 GND.n1388 0.152939
R22520 GND.n1394 GND.n1393 0.152939
R22521 GND.n1395 GND.n1394 0.152939
R22522 GND.n1396 GND.n1395 0.152939
R22523 GND.n1401 GND.n1396 0.152939
R22524 GND.n1402 GND.n1401 0.152939
R22525 GND.n1403 GND.n1402 0.152939
R22526 GND.n1404 GND.n1403 0.152939
R22527 GND.n1409 GND.n1404 0.152939
R22528 GND.n1410 GND.n1409 0.152939
R22529 GND.n1411 GND.n1410 0.152939
R22530 GND.n1412 GND.n1411 0.152939
R22531 GND.n1417 GND.n1412 0.152939
R22532 GND.n1418 GND.n1417 0.152939
R22533 GND.n1419 GND.n1418 0.152939
R22534 GND.n1420 GND.n1419 0.152939
R22535 GND.n1425 GND.n1420 0.152939
R22536 GND.n1426 GND.n1425 0.152939
R22537 GND.n1427 GND.n1426 0.152939
R22538 GND.n1428 GND.n1427 0.152939
R22539 GND.n1433 GND.n1428 0.152939
R22540 GND.n1434 GND.n1433 0.152939
R22541 GND.n1435 GND.n1434 0.152939
R22542 GND.n1436 GND.n1435 0.152939
R22543 GND.n1441 GND.n1436 0.152939
R22544 GND.n1442 GND.n1441 0.152939
R22545 GND.n1443 GND.n1442 0.152939
R22546 GND.n1444 GND.n1443 0.152939
R22547 GND.n5938 GND.n5937 0.152939
R22548 GND.n5937 GND.n5936 0.152939
R22549 GND.n5936 GND.n1708 0.152939
R22550 GND.n5932 GND.n1708 0.152939
R22551 GND.n5932 GND.n5931 0.152939
R22552 GND.n5931 GND.n5930 0.152939
R22553 GND.n5930 GND.n1713 0.152939
R22554 GND.n5926 GND.n1713 0.152939
R22555 GND.n5926 GND.n5925 0.152939
R22556 GND.n5925 GND.n5924 0.152939
R22557 GND.n5924 GND.n1718 0.152939
R22558 GND.n5920 GND.n1718 0.152939
R22559 GND.n5920 GND.n5919 0.152939
R22560 GND.n5919 GND.n5918 0.152939
R22561 GND.n5918 GND.n1723 0.152939
R22562 GND.n5914 GND.n1723 0.152939
R22563 GND.n5914 GND.n5913 0.152939
R22564 GND.n5913 GND.n5912 0.152939
R22565 GND.n5912 GND.n1728 0.152939
R22566 GND.n5908 GND.n1728 0.152939
R22567 GND.n5908 GND.n5907 0.152939
R22568 GND.n5907 GND.n5906 0.152939
R22569 GND.n5906 GND.n1733 0.152939
R22570 GND.n5902 GND.n1733 0.152939
R22571 GND.n5902 GND.n5901 0.152939
R22572 GND.n5901 GND.n5900 0.152939
R22573 GND.n5900 GND.n1738 0.152939
R22574 GND.n5896 GND.n1738 0.152939
R22575 GND.n5896 GND.n5895 0.152939
R22576 GND.n5886 GND.n5885 0.152939
R22577 GND.n5885 GND.n5884 0.152939
R22578 GND.n5884 GND.n1786 0.152939
R22579 GND.n5880 GND.n1786 0.152939
R22580 GND.n5880 GND.n5879 0.152939
R22581 GND.n5879 GND.n5878 0.152939
R22582 GND.n5878 GND.n1792 0.152939
R22583 GND.n5874 GND.n1792 0.152939
R22584 GND.n5874 GND.n5873 0.152939
R22585 GND.n5873 GND.n5872 0.152939
R22586 GND.n5872 GND.n1798 0.152939
R22587 GND.n5867 GND.n1798 0.152939
R22588 GND.n5867 GND.n5866 0.152939
R22589 GND.n5866 GND.n5865 0.152939
R22590 GND.n5865 GND.n1806 0.152939
R22591 GND.n5861 GND.n1806 0.152939
R22592 GND.n5861 GND.n5860 0.152939
R22593 GND.n5860 GND.n5859 0.152939
R22594 GND.n5859 GND.n1812 0.152939
R22595 GND.n5855 GND.n1812 0.152939
R22596 GND.n5855 GND.n5854 0.152939
R22597 GND.n3132 GND.n1818 0.152939
R22598 GND.n3132 GND.n3129 0.152939
R22599 GND.n3138 GND.n3129 0.152939
R22600 GND.n3139 GND.n3138 0.152939
R22601 GND.n3140 GND.n3139 0.152939
R22602 GND.n3140 GND.n3125 0.152939
R22603 GND.n3146 GND.n3125 0.152939
R22604 GND.n3147 GND.n3146 0.152939
R22605 GND.n3148 GND.n3147 0.152939
R22606 GND.n3148 GND.n3121 0.152939
R22607 GND.n3154 GND.n3121 0.152939
R22608 GND.n3155 GND.n3154 0.152939
R22609 GND.n3156 GND.n3155 0.152939
R22610 GND.n3156 GND.n3115 0.152939
R22611 GND.n3162 GND.n3115 0.152939
R22612 GND.n3163 GND.n3162 0.152939
R22613 GND.n3164 GND.n3163 0.152939
R22614 GND.n3164 GND.n3111 0.152939
R22615 GND.n3170 GND.n3111 0.152939
R22616 GND.n3171 GND.n3170 0.152939
R22617 GND.n3172 GND.n3171 0.152939
R22618 GND.n3172 GND.n3107 0.152939
R22619 GND.n3178 GND.n3107 0.152939
R22620 GND.n3179 GND.n3178 0.152939
R22621 GND.n3180 GND.n3179 0.152939
R22622 GND.n3180 GND.n3099 0.152939
R22623 GND.n6000 GND.n1650 0.152939
R22624 GND.n6000 GND.n5999 0.152939
R22625 GND.n5999 GND.n5998 0.152939
R22626 GND.n5998 GND.n1652 0.152939
R22627 GND.n5994 GND.n1652 0.152939
R22628 GND.n5994 GND.n5993 0.152939
R22629 GND.n5993 GND.n5992 0.152939
R22630 GND.n5992 GND.n1658 0.152939
R22631 GND.n5988 GND.n1658 0.152939
R22632 GND.n5988 GND.n5987 0.152939
R22633 GND.n5987 GND.n5986 0.152939
R22634 GND.n5984 GND.n1667 0.152939
R22635 GND.n5980 GND.n1667 0.152939
R22636 GND.n5980 GND.n5979 0.152939
R22637 GND.n5979 GND.n5978 0.152939
R22638 GND.n5978 GND.n1672 0.152939
R22639 GND.n5974 GND.n1672 0.152939
R22640 GND.n5974 GND.n5973 0.152939
R22641 GND.n5973 GND.n5972 0.152939
R22642 GND.n5972 GND.n1677 0.152939
R22643 GND.n5968 GND.n1677 0.152939
R22644 GND.n5968 GND.n5967 0.152939
R22645 GND.n5967 GND.n5966 0.152939
R22646 GND.n5966 GND.n1682 0.152939
R22647 GND.n5962 GND.n1682 0.152939
R22648 GND.n5962 GND.n5961 0.152939
R22649 GND.n5961 GND.n5960 0.152939
R22650 GND.n5960 GND.n1687 0.152939
R22651 GND.n5956 GND.n1687 0.152939
R22652 GND.n5956 GND.n5955 0.152939
R22653 GND.n5955 GND.n5954 0.152939
R22654 GND.n5954 GND.n1692 0.152939
R22655 GND.n5950 GND.n1692 0.152939
R22656 GND.n5950 GND.n5949 0.152939
R22657 GND.n5949 GND.n5948 0.152939
R22658 GND.n5948 GND.n1697 0.152939
R22659 GND.n5944 GND.n1697 0.152939
R22660 GND.n5944 GND.n5943 0.152939
R22661 GND.n5943 GND.n5942 0.152939
R22662 GND.n5942 GND.n1702 0.152939
R22663 GND.n2766 GND.n38 0.143793
R22664 GND.n3942 GND.n3941 0.143793
R22665 GND.n7820 GND.n36 0.0767195
R22666 GND.n7820 GND.n37 0.0767195
R22667 GND.n3329 GND.n3308 0.0767195
R22668 GND.n3342 GND.n3329 0.0767195
R22669 GND.n7828 GND.n22 0.0695946
R22670 GND.n7828 GND.n7827 0.0695946
R22671 GND.n5938 GND.n1707 0.0695946
R22672 GND.n1707 GND.n1702 0.0695946
R22673 GND.n4904 GND.n4903 0.063
R22674 GND.n4228 GND.n4227 0.063
R22675 GND.n4904 GND.n2602 0.0399022
R22676 GND.n7741 GND.n178 0.0399022
R22677 GND.n3665 GND.n3654 0.0399022
R22678 GND.n4227 GND.n4226 0.0399022
R22679 GND.n5329 GND.n2602 0.0344674
R22680 GND.n5329 GND.n2603 0.0344674
R22681 GND.n4925 GND.n2603 0.0344674
R22682 GND.n4925 GND.n4924 0.0344674
R22683 GND.n4931 GND.n4924 0.0344674
R22684 GND.n4932 GND.n4931 0.0344674
R22685 GND.n4932 GND.n2642 0.0344674
R22686 GND.n2643 GND.n2642 0.0344674
R22687 GND.n2644 GND.n2643 0.0344674
R22688 GND.n4947 GND.n2644 0.0344674
R22689 GND.n4947 GND.n2663 0.0344674
R22690 GND.n2664 GND.n2663 0.0344674
R22691 GND.n2665 GND.n2664 0.0344674
R22692 GND.n4962 GND.n2665 0.0344674
R22693 GND.n4962 GND.n2684 0.0344674
R22694 GND.n2685 GND.n2684 0.0344674
R22695 GND.n2686 GND.n2685 0.0344674
R22696 GND.n4977 GND.n2686 0.0344674
R22697 GND.n4977 GND.n2705 0.0344674
R22698 GND.n2706 GND.n2705 0.0344674
R22699 GND.n2707 GND.n2706 0.0344674
R22700 GND.n4992 GND.n2707 0.0344674
R22701 GND.n4992 GND.n2725 0.0344674
R22702 GND.n2726 GND.n2725 0.0344674
R22703 GND.n2727 GND.n2726 0.0344674
R22704 GND.n5018 GND.n2727 0.0344674
R22705 GND.n5021 GND.n5018 0.0344674
R22706 GND.n5022 GND.n5021 0.0344674
R22707 GND.n5022 GND.n2751 0.0344674
R22708 GND.n2752 GND.n2751 0.0344674
R22709 GND.n2753 GND.n2752 0.0344674
R22710 GND.n5030 GND.n2753 0.0344674
R22711 GND.n5031 GND.n5030 0.0344674
R22712 GND.n5031 GND.n54 0.0344674
R22713 GND.n55 GND.n54 0.0344674
R22714 GND.n56 GND.n55 0.0344674
R22715 GND.n2809 GND.n56 0.0344674
R22716 GND.n2809 GND.n73 0.0344674
R22717 GND.n74 GND.n73 0.0344674
R22718 GND.n75 GND.n74 0.0344674
R22719 GND.n2804 GND.n75 0.0344674
R22720 GND.n2804 GND.n94 0.0344674
R22721 GND.n95 GND.n94 0.0344674
R22722 GND.n96 GND.n95 0.0344674
R22723 GND.n2799 GND.n96 0.0344674
R22724 GND.n2799 GND.n115 0.0344674
R22725 GND.n116 GND.n115 0.0344674
R22726 GND.n117 GND.n116 0.0344674
R22727 GND.n2794 GND.n117 0.0344674
R22728 GND.n2794 GND.n136 0.0344674
R22729 GND.n137 GND.n136 0.0344674
R22730 GND.n138 GND.n137 0.0344674
R22731 GND.n5104 GND.n138 0.0344674
R22732 GND.n5104 GND.n156 0.0344674
R22733 GND.n157 GND.n156 0.0344674
R22734 GND.n158 GND.n157 0.0344674
R22735 GND.n5158 GND.n158 0.0344674
R22736 GND.n5158 GND.n177 0.0344674
R22737 GND.n7741 GND.n177 0.0344674
R22738 GND.n3665 GND.n3664 0.0344674
R22739 GND.n3664 GND.n3663 0.0344674
R22740 GND.n3663 GND.n3661 0.0344674
R22741 GND.n3661 GND.n3463 0.0344674
R22742 GND.n3703 GND.n3463 0.0344674
R22743 GND.n3703 GND.n3464 0.0344674
R22744 GND.n3699 GND.n3464 0.0344674
R22745 GND.n3699 GND.n3698 0.0344674
R22746 GND.n3698 GND.n3434 0.0344674
R22747 GND.n3740 GND.n3434 0.0344674
R22748 GND.n3740 GND.n3435 0.0344674
R22749 GND.n3736 GND.n3435 0.0344674
R22750 GND.n3736 GND.n3735 0.0344674
R22751 GND.n3735 GND.n3405 0.0344674
R22752 GND.n3777 GND.n3405 0.0344674
R22753 GND.n3777 GND.n3406 0.0344674
R22754 GND.n3773 GND.n3406 0.0344674
R22755 GND.n3773 GND.n3772 0.0344674
R22756 GND.n3772 GND.n3375 0.0344674
R22757 GND.n3814 GND.n3375 0.0344674
R22758 GND.n3814 GND.n3377 0.0344674
R22759 GND.n3377 GND.n3376 0.0344674
R22760 GND.n3376 GND.n3355 0.0344674
R22761 GND.n3834 GND.n3355 0.0344674
R22762 GND.n3834 GND.n3352 0.0344674
R22763 GND.n3927 GND.n3352 0.0344674
R22764 GND.n3927 GND.n3353 0.0344674
R22765 GND.n3923 GND.n3353 0.0344674
R22766 GND.n3923 GND.n3922 0.0344674
R22767 GND.n3922 GND.n3921 0.0344674
R22768 GND.n3921 GND.n3845 0.0344674
R22769 GND.n3917 GND.n3845 0.0344674
R22770 GND.n3917 GND.n3916 0.0344674
R22771 GND.n3916 GND.n3915 0.0344674
R22772 GND.n3915 GND.n3317 0.0344674
R22773 GND.n3960 GND.n3317 0.0344674
R22774 GND.n3960 GND.n3318 0.0344674
R22775 GND.n3956 GND.n3318 0.0344674
R22776 GND.n3956 GND.n3955 0.0344674
R22777 GND.n3955 GND.n3289 0.0344674
R22778 GND.n3997 GND.n3289 0.0344674
R22779 GND.n3997 GND.n3290 0.0344674
R22780 GND.n3993 GND.n3290 0.0344674
R22781 GND.n3993 GND.n3992 0.0344674
R22782 GND.n3992 GND.n3260 0.0344674
R22783 GND.n4034 GND.n3260 0.0344674
R22784 GND.n4034 GND.n3261 0.0344674
R22785 GND.n4030 GND.n3261 0.0344674
R22786 GND.n4030 GND.n4029 0.0344674
R22787 GND.n4029 GND.n3231 0.0344674
R22788 GND.n4071 GND.n3231 0.0344674
R22789 GND.n4071 GND.n3232 0.0344674
R22790 GND.n4067 GND.n3232 0.0344674
R22791 GND.n4067 GND.n4066 0.0344674
R22792 GND.n4066 GND.n3202 0.0344674
R22793 GND.n4137 GND.n3202 0.0344674
R22794 GND.n4137 GND.n3203 0.0344674
R22795 GND.n3203 GND.n3100 0.0344674
R22796 GND.n4226 GND.n3100 0.0344674
R22797 GND.n4229 GND.n4228 0.0157439
R22798 GND.n4903 GND.n2398 0.0157439
R22799 GND.n4903 GND.n2399 0.0112041
R22800 GND.n4228 GND.n3098 0.0112041
R22801 GND.n4799 GND.n4798 0.0108473
R22802 GND.n5894 GND.n5893 0.0108473
R22803 GND.n3943 GND.n3942 0.00964634
R22804 GND.n2862 GND.n38 0.00964634
R22805 GND.n2901 GND.n2399 0.0084686
R22806 GND.n2904 GND.n2400 0.0084686
R22807 GND.n2906 GND.n2401 0.0084686
R22808 GND.n2910 GND.n2402 0.0084686
R22809 GND.n2912 GND.n2403 0.0084686
R22810 GND.n2916 GND.n2404 0.0084686
R22811 GND.n2918 GND.n2405 0.0084686
R22812 GND.n2922 GND.n2406 0.0084686
R22813 GND.n2924 GND.n2410 0.0084686
R22814 GND.n2929 GND.n2411 0.0084686
R22815 GND.n2898 GND.n2412 0.0084686
R22816 GND.n4799 GND.n2413 0.0084686
R22817 GND.n4219 GND.n3098 0.0084686
R22818 GND.n4218 GND.n4152 0.0084686
R22819 GND.n4215 GND.n4214 0.0084686
R22820 GND.n4211 GND.n4157 0.0084686
R22821 GND.n4210 GND.n4163 0.0084686
R22822 GND.n4207 GND.n4206 0.0084686
R22823 GND.n4203 GND.n4170 0.0084686
R22824 GND.n4202 GND.n4174 0.0084686
R22825 GND.n4196 GND.n4195 0.0084686
R22826 GND.n4192 GND.n4180 0.0084686
R22827 GND.n4191 GND.n4184 0.0084686
R22828 GND.n5893 GND.n1744 0.0084686
R22829 GND.n2901 GND.n2400 0.00442483
R22830 GND.n2904 GND.n2401 0.00442483
R22831 GND.n2906 GND.n2402 0.00442483
R22832 GND.n2910 GND.n2403 0.00442483
R22833 GND.n2912 GND.n2404 0.00442483
R22834 GND.n2916 GND.n2405 0.00442483
R22835 GND.n2918 GND.n2406 0.00442483
R22836 GND.n2922 GND.n2410 0.00442483
R22837 GND.n2924 GND.n2411 0.00442483
R22838 GND.n2929 GND.n2412 0.00442483
R22839 GND.n2898 GND.n2413 0.00442483
R22840 GND.n4219 GND.n4218 0.00442483
R22841 GND.n4215 GND.n4152 0.00442483
R22842 GND.n4214 GND.n4157 0.00442483
R22843 GND.n4211 GND.n4210 0.00442483
R22844 GND.n4207 GND.n4163 0.00442483
R22845 GND.n4206 GND.n4170 0.00442483
R22846 GND.n4203 GND.n4202 0.00442483
R22847 GND.n4196 GND.n4174 0.00442483
R22848 GND.n4195 GND.n4180 0.00442483
R22849 GND.n4192 GND.n4191 0.00442483
R22850 GND.n4184 GND.n1744 0.00442483
R22851 VN.n4 VN.t0 243.97
R22852 VN.n4 VN.n3 223.454
R22853 VN.n6 VN.n5 223.454
R22854 VN.n8 VN.n7 223.454
R22855 VN.n1 VN.t10 44.8721
R22856 VN.n0 VN.t8 44.8719
R22857 VN.n1 VN.t7 42.7258
R22858 VN.n0 VN.t9 42.7258
R22859 VN.n2 VN.n1 38.6431
R22860 VN.n3 VN.t3 19.8005
R22861 VN.n3 VN.t4 19.8005
R22862 VN.n5 VN.t1 19.8005
R22863 VN.n5 VN.t6 19.8005
R22864 VN.n7 VN.t2 19.8005
R22865 VN.n7 VN.t5 19.8005
R22866 VN VN.n9 18.0539
R22867 VN.n2 VN.n0 13.4878
R22868 VN.n9 VN.n8 5.40567
R22869 VN.n9 VN.n2 1.188
R22870 VN.n8 VN.n6 0.716017
R22871 VN.n6 VN.n4 0.716017
R22872 a_n2596_242.n0 a_n2596_242.t8 194.494
R22873 a_n2596_242.t1 a_n2596_242.n0 194.494
R22874 a_n2596_242.n0 a_n2596_242.t2 96.9377
R22875 a_n2596_242.n0 a_n2596_242.t0 86.719
R22876 a_n2596_242.n0 a_n2596_242.t3 86.719
R22877 a_n2596_242.n0 a_n2596_242.t7 86.719
R22878 a_n2596_242.n0 a_n2596_242.t6 86.719
R22879 a_n2596_242.n0 a_n2596_242.t4 86.719
R22880 a_n2596_242.n0 a_n2596_242.t5 86.7188
R22881 a_n2596_242.n0 a_n2596_242.t9 86.7188
R22882 a_n17822_7210.n30 a_n17822_7210.n28 137.044
R22883 a_n17822_7210.n27 a_n17822_7210.n25 137.044
R22884 a_n17822_7210.n30 a_n17822_7210.n29 135.334
R22885 a_n17822_7210.n27 a_n17822_7210.n26 135.334
R22886 a_n17822_7210.n33 a_n17822_7210.n32 119.757
R22887 a_n17822_7210.n34 a_n17822_7210.n33 88.9373
R22888 a_n17822_7210.n18 a_n17822_7210.n19 0.920017
R22889 a_n17822_7210.n16 a_n17822_7210.n17 0.920017
R22890 a_n17822_7210.n14 a_n17822_7210.n15 0.920017
R22891 a_n17822_7210.n12 a_n17822_7210.n13 0.920017
R22892 a_n17822_7210.n10 a_n17822_7210.n11 0.920018
R22893 a_n17822_7210.n8 a_n17822_7210.n9 0.836337
R22894 a_n17822_7210.n6 a_n17822_7210.n7 0.836337
R22895 a_n17822_7210.n4 a_n17822_7210.n5 0.836337
R22896 a_n17822_7210.n2 a_n17822_7210.n3 0.836337
R22897 a_n17822_7210.n0 a_n17822_7210.n1 0.836337
R22898 a_n17822_7210.n10 a_n17822_7210.t35 59.5667
R22899 a_n17822_7210.n8 a_n17822_7210.t31 59.5667
R22900 a_n17822_7210.n6 a_n17822_7210.t26 59.5667
R22901 a_n17822_7210.n4 a_n17822_7210.t25 59.5667
R22902 a_n17822_7210.n2 a_n17822_7210.t20 59.5667
R22903 a_n17822_7210.n0 a_n17822_7210.t12 59.5667
R22904 a_n17822_7210.n18 a_n17822_7210.t22 59.5665
R22905 a_n17822_7210.n16 a_n17822_7210.t14 59.5665
R22906 a_n17822_7210.n14 a_n17822_7210.t16 59.5665
R22907 a_n17822_7210.n12 a_n17822_7210.t39 59.5665
R22908 a_n17822_7210.n31 a_n17822_7210.n27 33.3106
R22909 a_n17822_7210.n19 a_n17822_7210.t17 58.1638
R22910 a_n17822_7210.n19 a_n17822_7210.t34 60.6625
R22911 a_n17822_7210.n17 a_n17822_7210.t41 58.1638
R22912 a_n17822_7210.n17 a_n17822_7210.t30 60.6625
R22913 a_n17822_7210.n15 a_n17822_7210.t38 58.1638
R22914 a_n17822_7210.n15 a_n17822_7210.t28 60.6625
R22915 a_n17822_7210.n13 a_n17822_7210.t33 58.1638
R22916 a_n17822_7210.n13 a_n17822_7210.t23 60.6625
R22917 a_n17822_7210.n11 a_n17822_7210.t15 60.6625
R22918 a_n17822_7210.n11 a_n17822_7210.t27 58.1638
R22919 a_n17822_7210.n9 a_n17822_7210.t37 57.4776
R22920 a_n17822_7210.n9 a_n17822_7210.t21 61.4742
R22921 a_n17822_7210.n7 a_n17822_7210.t32 57.4776
R22922 a_n17822_7210.n7 a_n17822_7210.t13 61.4742
R22923 a_n17822_7210.n5 a_n17822_7210.t19 57.4776
R22924 a_n17822_7210.n5 a_n17822_7210.t29 61.4742
R22925 a_n17822_7210.n3 a_n17822_7210.t40 57.4776
R22926 a_n17822_7210.n3 a_n17822_7210.t24 61.4742
R22927 a_n17822_7210.n1 a_n17822_7210.t36 57.4776
R22928 a_n17822_7210.n1 a_n17822_7210.t18 61.4742
R22929 a_n17822_7210.n31 a_n17822_7210.n30 24.6118
R22930 a_n17822_7210.n29 a_n17822_7210.t11 22.3407
R22931 a_n17822_7210.n29 a_n17822_7210.t10 22.3407
R22932 a_n17822_7210.n28 a_n17822_7210.t4 22.3407
R22933 a_n17822_7210.n28 a_n17822_7210.t5 22.3407
R22934 a_n17822_7210.n25 a_n17822_7210.t6 22.3407
R22935 a_n17822_7210.n25 a_n17822_7210.t9 22.3407
R22936 a_n17822_7210.n26 a_n17822_7210.t8 22.3407
R22937 a_n17822_7210.n26 a_n17822_7210.t7 22.3407
R22938 a_n17822_7210.n32 a_n17822_7210.t1 17.3689
R22939 a_n17822_7210.n32 a_n17822_7210.t2 17.3689
R22940 a_n17822_7210.n34 a_n17822_7210.t0 17.3689
R22941 a_n17822_7210.t3 a_n17822_7210.n34 17.3689
R22942 a_n17822_7210.n33 a_n17822_7210.n20 12.4007
R22943 a_n17822_7210.n20 a_n17822_7210.n31 11.9628
R22944 a_n17822_7210.n20 a_n17822_7210.n22 10.0448
R22945 a_n17822_7210.n21 a_n17822_7210.n10 8.47786
R22946 a_n17822_7210.n23 a_n17822_7210.n0 8.47786
R22947 a_n17822_7210.n23 a_n17822_7210.n4 8.47786
R22948 a_n17822_7210.n21 a_n17822_7210.n14 8.47786
R22949 a_n17822_7210.n20 a_n17822_7210.n24 7.05156
R22950 a_n17822_7210.n24 a_n17822_7210.n23 6.35277
R22951 a_n17822_7210.n22 a_n17822_7210.n21 6.35277
R22952 a_n17822_7210.n22 a_n17822_7210.n18 5.30172
R22953 a_n17822_7210.n22 a_n17822_7210.n16 5.30172
R22954 a_n17822_7210.n21 a_n17822_7210.n12 5.30172
R22955 a_n17822_7210.n24 a_n17822_7210.n8 5.30172
R22956 a_n17822_7210.n24 a_n17822_7210.n6 5.30172
R22957 a_n17822_7210.n23 a_n17822_7210.n2 5.30172
R22958 a_n6906_9317.n3 a_n6906_9317.t2 139.797
R22959 a_n6906_9317.n1 a_n6906_9317.t9 139.797
R22960 a_n6906_9317.n0 a_n6906_9317.t7 139.797
R22961 a_n6906_9317.n3 a_n6906_9317.t4 138.088
R22962 a_n6906_9317.n0 a_n6906_9317.t3 138.088
R22963 a_n6906_9317.n1 a_n6906_9317.t16 138.088
R22964 a_n6906_9317.n1 a_n6906_9317.t15 138.088
R22965 a_n6906_9317.n2 a_n6906_9317.t11 138.088
R22966 a_n6906_9317.n0 a_n6906_9317.n4 115.746
R22967 a_n6906_9317.n1 a_n6906_9317.n6 115.746
R22968 a_n6906_9317.n2 a_n6906_9317.n7 115.746
R22969 a_n6906_9317.n9 a_n6906_9317.n3 115.746
R22970 a_n6906_9317.n3 a_n6906_9317.n8 28.1107
R22971 a_n6906_9317.n4 a_n6906_9317.t5 22.3407
R22972 a_n6906_9317.n4 a_n6906_9317.t6 22.3407
R22973 a_n6906_9317.n6 a_n6906_9317.t12 22.3407
R22974 a_n6906_9317.n6 a_n6906_9317.t10 22.3407
R22975 a_n6906_9317.n7 a_n6906_9317.t13 22.3407
R22976 a_n6906_9317.n7 a_n6906_9317.t14 22.3407
R22977 a_n6906_9317.t8 a_n6906_9317.n9 22.3407
R22978 a_n6906_9317.n9 a_n6906_9317.t1 22.3407
R22979 a_n6906_9317.n5 a_n6906_9317.t0 17.1466
R22980 a_n6906_9317.n5 a_n6906_9317.n0 10.29
R22981 a_n6906_9317.n8 a_n6906_9317.n2 5.76343
R22982 a_n6906_9317.n2 a_n6906_9317.n1 5.54145
R22983 a_n6906_9317.n8 a_n6906_9317.n5 3.58762
R22984 VP.n8 VP.t6 243.255
R22985 VP.n5 VP.n3 224.169
R22986 VP.n7 VP.n6 223.454
R22987 VP.n5 VP.n4 223.454
R22988 VP.n0 VP.t7 44.8721
R22989 VP.n1 VP.t9 44.8719
R22990 VP.n1 VP.t10 42.7258
R22991 VP.n0 VP.t8 42.7258
R22992 VP.n2 VP.n1 38.859
R22993 VP.n6 VP.t4 19.8005
R22994 VP.n6 VP.t0 19.8005
R22995 VP.n4 VP.t3 19.8005
R22996 VP.n4 VP.t2 19.8005
R22997 VP.n3 VP.t5 19.8005
R22998 VP.n3 VP.t1 19.8005
R22999 VP VP.n9 14.2554
R23000 VP.n2 VP.n0 13.7037
R23001 VP.n9 VP.n8 4.80222
R23002 VP.n9 VP.n2 0.972091
R23003 VP.n7 VP.n5 0.716017
R23004 VP.n8 VP.n7 0.716017
R23005 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t3 128.209
R23006 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t1 127.002
R23007 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t2 46.923
R23008 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t5 43.4256
R23009 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t0 43.2987
R23010 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t4 42.6649
R23011 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 6.38688
R23012 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 4.61307
R23013 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n0 4.34443
R23014 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 2.57317
R23015 DIFFPAIR_BIAS DIFFPAIR_BIAS.n4 0.753625
C0 VDD VOUT 64.9369f
C1 VOUT VP 4.82961f
C2 VDD VN 0.188398f
C3 a_n12301_11007# VDD 1.80787f
C4 VOUT VN 1.09056f
C5 VP VN 12.9376f
C6 VOUT CS_BIAS 19.625801f
C7 VP CS_BIAS 0.333631f
C8 VP DIFFPAIR_BIAS 3.21e-20
C9 VN CS_BIAS 0.288971f
C10 VN DIFFPAIR_BIAS 9.01e-20
C11 a_10955_11007# VDD 1.80788f
C12 DIFFPAIR_BIAS GND 25.161499f
C13 CS_BIAS GND 98.310875f
C14 VN GND 40.931038f
C15 VP GND 35.679066f
C16 VOUT GND 78.551f
C17 VDD GND 1.073463p
C18 a_10955_11007# GND 0.679905f
C19 a_n12301_11007# GND 0.679905f
C20 VP.t8 GND 0.860307f
C21 VP.t7 GND 0.88538f
C22 VP.n0 GND 1.24445f
C23 VP.t9 GND 0.885379f
C24 VP.t10 GND 0.860307f
C25 VP.n1 GND 1.76849f
C26 VP.n2 GND 1.15029f
C27 VP.t5 GND 0.006002f
C28 VP.t1 GND 0.006002f
C29 VP.n3 GND 0.019735f
C30 VP.t3 GND 0.006002f
C31 VP.t2 GND 0.006002f
C32 VP.n4 GND 0.019465f
C33 VP.n5 GND 0.166122f
C34 VP.t4 GND 0.006002f
C35 VP.t0 GND 0.006002f
C36 VP.n6 GND 0.019465f
C37 VP.n7 GND 0.081667f
C38 VP.t6 GND 0.033405f
C39 VP.n8 GND 0.090651f
C40 VP.n9 GND 2.58022f
C41 a_n6906_9317.n0 GND 6.28071f
C42 a_n6906_9317.n1 GND 5.1637f
C43 a_n6906_9317.n2 GND 3.64828f
C44 a_n6906_9317.n3 GND 8.00118f
C45 a_n6906_9317.t0 GND 38.9884f
C46 a_n6906_9317.t1 GND 0.063311f
C47 a_n6906_9317.t7 GND 0.344107f
C48 a_n6906_9317.t5 GND 0.063311f
C49 a_n6906_9317.t6 GND 0.063311f
C50 a_n6906_9317.n4 GND 0.233095f
C51 a_n6906_9317.t3 GND 0.33106f
C52 a_n6906_9317.n5 GND 5.9593f
C53 a_n6906_9317.t9 GND 0.344108f
C54 a_n6906_9317.t12 GND 0.063311f
C55 a_n6906_9317.t10 GND 0.063311f
C56 a_n6906_9317.n6 GND 0.233095f
C57 a_n6906_9317.t16 GND 0.33106f
C58 a_n6906_9317.t15 GND 0.33106f
C59 a_n6906_9317.t13 GND 0.063311f
C60 a_n6906_9317.t14 GND 0.063311f
C61 a_n6906_9317.n7 GND 0.233095f
C62 a_n6906_9317.t11 GND 0.33106f
C63 a_n6906_9317.n8 GND 5.23198f
C64 a_n6906_9317.t4 GND 0.33106f
C65 a_n6906_9317.t2 GND 0.344108f
C66 a_n6906_9317.n9 GND 0.233096f
C67 a_n6906_9317.t8 GND 0.063311f
C68 a_n17822_7210.n0 GND 1.88958f
C69 a_n17822_7210.n1 GND 1.06501f
C70 a_n17822_7210.n2 GND 1.82295f
C71 a_n17822_7210.n3 GND 1.06501f
C72 a_n17822_7210.n4 GND 1.82295f
C73 a_n17822_7210.n5 GND 1.06501f
C74 a_n17822_7210.n6 GND 1.82295f
C75 a_n17822_7210.n7 GND 1.06501f
C76 a_n17822_7210.n8 GND 1.82295f
C77 a_n17822_7210.n9 GND 1.06501f
C78 a_n17822_7210.n10 GND 1.88958f
C79 a_n17822_7210.n11 GND 1.06527f
C80 a_n17822_7210.n12 GND 1.82295f
C81 a_n17822_7210.n13 GND 1.06527f
C82 a_n17822_7210.n14 GND 1.82295f
C83 a_n17822_7210.n15 GND 1.06527f
C84 a_n17822_7210.n16 GND 1.82295f
C85 a_n17822_7210.n17 GND 1.06527f
C86 a_n17822_7210.n18 GND 1.82295f
C87 a_n17822_7210.n19 GND 1.06527f
C88 a_n17822_7210.n20 GND 23.474699f
C89 a_n17822_7210.n21 GND 0.757534f
C90 a_n17822_7210.n22 GND 2.50277f
C91 a_n17822_7210.n23 GND 0.757534f
C92 a_n17822_7210.n24 GND 3.113f
C93 a_n17822_7210.t0 GND 0.041125f
C94 a_n17822_7210.t6 GND 0.052488f
C95 a_n17822_7210.t9 GND 0.052488f
C96 a_n17822_7210.n25 GND 0.258428f
C97 a_n17822_7210.t8 GND 0.052488f
C98 a_n17822_7210.t7 GND 0.052488f
C99 a_n17822_7210.n26 GND 0.24055f
C100 a_n17822_7210.n27 GND 6.9299f
C101 a_n17822_7210.t4 GND 0.052488f
C102 a_n17822_7210.t5 GND 0.052488f
C103 a_n17822_7210.n28 GND 0.258428f
C104 a_n17822_7210.t11 GND 0.052488f
C105 a_n17822_7210.t10 GND 0.052488f
C106 a_n17822_7210.n29 GND 0.24055f
C107 a_n17822_7210.n30 GND 6.35108f
C108 a_n17822_7210.n31 GND 11.5894f
C109 a_n17822_7210.t18 GND 2.3544f
C110 a_n17822_7210.t12 GND 2.34255f
C111 a_n17822_7210.t36 GND 2.30996f
C112 a_n17822_7210.t24 GND 2.3544f
C113 a_n17822_7210.t20 GND 2.34255f
C114 a_n17822_7210.t40 GND 2.30996f
C115 a_n17822_7210.t29 GND 2.3544f
C116 a_n17822_7210.t25 GND 2.34255f
C117 a_n17822_7210.t19 GND 2.30996f
C118 a_n17822_7210.t13 GND 2.3544f
C119 a_n17822_7210.t26 GND 2.34255f
C120 a_n17822_7210.t32 GND 2.30996f
C121 a_n17822_7210.t21 GND 2.3544f
C122 a_n17822_7210.t31 GND 2.34255f
C123 a_n17822_7210.t37 GND 2.30996f
C124 a_n17822_7210.t27 GND 2.32216f
C125 a_n17822_7210.t35 GND 2.34255f
C126 a_n17822_7210.t15 GND 2.34195f
C127 a_n17822_7210.t33 GND 2.32216f
C128 a_n17822_7210.t39 GND 2.34254f
C129 a_n17822_7210.t23 GND 2.34195f
C130 a_n17822_7210.t38 GND 2.32216f
C131 a_n17822_7210.t16 GND 2.34254f
C132 a_n17822_7210.t28 GND 2.34195f
C133 a_n17822_7210.t41 GND 2.32216f
C134 a_n17822_7210.t14 GND 2.34254f
C135 a_n17822_7210.t30 GND 2.34195f
C136 a_n17822_7210.t17 GND 2.32216f
C137 a_n17822_7210.t22 GND 2.34254f
C138 a_n17822_7210.t34 GND 2.34195f
C139 a_n17822_7210.t1 GND 0.041125f
C140 a_n17822_7210.t2 GND 0.041125f
C141 a_n17822_7210.n32 GND 1.10971f
C142 a_n17822_7210.n33 GND 6.299181f
C143 a_n17822_7210.n34 GND 0.250903f
C144 a_n17822_7210.t3 GND 0.041125f
C145 a_n2596_242.n0 GND 14.1385f
C146 a_n2596_242.t8 GND 0.390363f
C147 a_n2596_242.t4 GND 0.197598f
C148 a_n2596_242.t5 GND 0.197599f
C149 a_n2596_242.t9 GND 0.197599f
C150 a_n2596_242.t2 GND 0.197599f
C151 a_n2596_242.t6 GND 0.197598f
C152 a_n2596_242.t7 GND 0.197598f
C153 a_n2596_242.t3 GND 0.197598f
C154 a_n2596_242.t0 GND 0.197598f
C155 a_n2596_242.t1 GND 0.390363f
C156 VN.t8 GND 0.591728f
C157 VN.t9 GND 0.574972f
C158 VN.n0 GND 0.828589f
C159 VN.t7 GND 0.574972f
C160 VN.t10 GND 0.591729f
C161 VN.n1 GND 1.17686f
C162 VN.n2 GND 0.763262f
C163 VN.t0 GND 0.022462f
C164 VN.t3 GND 0.004011f
C165 VN.t4 GND 0.004011f
C166 VN.n3 GND 0.013009f
C167 VN.n4 GND 0.100989f
C168 VN.t1 GND 0.004011f
C169 VN.t6 GND 0.004011f
C170 VN.n5 GND 0.013009f
C171 VN.n6 GND 0.054581f
C172 VN.t2 GND 0.004011f
C173 VN.t5 GND 0.004011f
C174 VN.n7 GND 0.013009f
C175 VN.n8 GND 0.075805f
C176 VN.n9 GND 3.03902f
C177 VOUT.t43 GND 0.058408f
C178 VOUT.t31 GND 0.058408f
C179 VOUT.n0 GND 0.328939f
C180 VOUT.t22 GND 0.407473f
C181 VOUT.n1 GND 1.64356f
C182 VOUT.t36 GND 0.058408f
C183 VOUT.t1 GND 0.058408f
C184 VOUT.n2 GND 0.328939f
C185 VOUT.t27 GND 0.407473f
C186 VOUT.n3 GND 1.58768f
C187 VOUT.n4 GND 0.742013f
C188 VOUT.t0 GND 0.058408f
C189 VOUT.t20 GND 0.058408f
C190 VOUT.n5 GND 0.328939f
C191 VOUT.t25 GND 0.407473f
C192 VOUT.n6 GND 1.58768f
C193 VOUT.n7 GND 0.521512f
C194 VOUT.t37 GND 0.058408f
C195 VOUT.t42 GND 0.058408f
C196 VOUT.n8 GND 0.328939f
C197 VOUT.t35 GND 0.407473f
C198 VOUT.n9 GND 1.58768f
C199 VOUT.n10 GND 0.521512f
C200 VOUT.t41 GND 0.058408f
C201 VOUT.t28 GND 0.058408f
C202 VOUT.n11 GND 0.328939f
C203 VOUT.t34 GND 0.407473f
C204 VOUT.n12 GND 1.58768f
C205 VOUT.n13 GND 0.734819f
C206 VOUT.n14 GND 12.0007f
C207 VOUT.t46 GND 12.8818f
C208 VOUT.t47 GND 8.16504f
C209 VOUT.n15 GND 10.7432f
C210 VOUT.n16 GND 2.41432f
C211 VOUT.t32 GND 0.415648f
C212 VOUT.t44 GND 0.058408f
C213 VOUT.t21 GND 0.058408f
C214 VOUT.n17 GND 0.315368f
C215 VOUT.n18 GND 1.60846f
C216 VOUT.t18 GND 0.415648f
C217 VOUT.t23 GND 0.058408f
C218 VOUT.t24 GND 0.058408f
C219 VOUT.n19 GND 0.315368f
C220 VOUT.n20 GND 1.55143f
C221 VOUT.n21 GND 0.824159f
C222 VOUT.t26 GND 0.415648f
C223 VOUT.t38 GND 0.058408f
C224 VOUT.t45 GND 0.058408f
C225 VOUT.n22 GND 0.315368f
C226 VOUT.n23 GND 1.55143f
C227 VOUT.n24 GND 0.563159f
C228 VOUT.t33 GND 0.415648f
C229 VOUT.t19 GND 0.058408f
C230 VOUT.t29 GND 0.058408f
C231 VOUT.n25 GND 0.315368f
C232 VOUT.n26 GND 1.55143f
C233 VOUT.n27 GND 0.563159f
C234 VOUT.t30 GND 0.415648f
C235 VOUT.t40 GND 0.058408f
C236 VOUT.t39 GND 0.058408f
C237 VOUT.n28 GND 0.315367f
C238 VOUT.n29 GND 1.55143f
C239 VOUT.n30 GND 0.776466f
C240 VOUT.n31 GND 16.237902f
C241 VOUT.t5 GND 0.034283f
C242 VOUT.t8 GND 0.034283f
C243 VOUT.n32 GND 0.302212f
C244 VOUT.t11 GND 0.034283f
C245 VOUT.t16 GND 0.034283f
C246 VOUT.n33 GND 0.289307f
C247 VOUT.n34 GND 2.5646f
C248 VOUT.t17 GND 0.034283f
C249 VOUT.t12 GND 0.034283f
C250 VOUT.n35 GND 0.289307f
C251 VOUT.n36 GND 1.37959f
C252 VOUT.t4 GND 0.034283f
C253 VOUT.t2 GND 0.034283f
C254 VOUT.n37 GND 0.289307f
C255 VOUT.n38 GND 1.61063f
C256 VOUT.n39 GND 14.141701f
C257 VOUT.t15 GND 0.034283f
C258 VOUT.t13 GND 0.034283f
C259 VOUT.n40 GND 0.302212f
C260 VOUT.t7 GND 0.034283f
C261 VOUT.t3 GND 0.034283f
C262 VOUT.n41 GND 0.289307f
C263 VOUT.n42 GND 2.5646f
C264 VOUT.t14 GND 0.034283f
C265 VOUT.t10 GND 0.034283f
C266 VOUT.n43 GND 0.289307f
C267 VOUT.n44 GND 1.37959f
C268 VOUT.t9 GND 0.034283f
C269 VOUT.t6 GND 0.034283f
C270 VOUT.n45 GND 0.289307f
C271 VOUT.n46 GND 1.61063f
C272 VOUT.n47 GND 9.86513f
C273 VOUT.n48 GND 8.60515f
C274 CS_BIAS.n0 GND 0.013689f
C275 CS_BIAS.t10 GND 0.251791f
C276 CS_BIAS.n1 GND 0.011007f
C277 CS_BIAS.n2 GND 0.005906f
C278 CS_BIAS.t12 GND 0.351512f
C279 CS_BIAS.n3 GND 0.088545f
C280 CS_BIAS.t4 GND 0.359096f
C281 CS_BIAS.t0 GND 0.368704f
C282 CS_BIAS.n4 GND 0.407887f
C283 CS_BIAS.t5 GND 0.010814f
C284 CS_BIAS.t1 GND 0.010814f
C285 CS_BIAS.n5 GND 0.069862f
C286 CS_BIAS.n6 GND 0.364691f
C287 CS_BIAS.n7 GND 0.136658f
C288 CS_BIAS.n8 GND 0.005159f
C289 CS_BIAS.n9 GND 0.013517f
C290 CS_BIAS.n10 GND 0.011897f
C291 CS_BIAS.n11 GND 0.011007f
C292 CS_BIAS.n12 GND 0.005906f
C293 CS_BIAS.n13 GND 0.005906f
C294 CS_BIAS.n14 GND 0.005906f
C295 CS_BIAS.n15 GND 0.011007f
C296 CS_BIAS.n16 GND 0.010626f
C297 CS_BIAS.n17 GND 0.127991f
C298 CS_BIAS.n18 GND 0.07598f
C299 CS_BIAS.t20 GND 0.359096f
C300 CS_BIAS.t18 GND 0.368704f
C301 CS_BIAS.n19 GND 0.360452f
C302 CS_BIAS.n20 GND 0.084384f
C303 CS_BIAS.t22 GND 0.359096f
C304 CS_BIAS.t21 GND 0.368704f
C305 CS_BIAS.n21 GND 0.360452f
C306 CS_BIAS.n22 GND 0.062575f
C307 CS_BIAS.t16 GND 0.368705f
C308 CS_BIAS.t19 GND 0.359096f
C309 CS_BIAS.n23 GND 0.360451f
C310 CS_BIAS.n24 GND 0.394928f
C311 CS_BIAS.n25 GND 0.013689f
C312 CS_BIAS.t13 GND 0.251791f
C313 CS_BIAS.n26 GND 0.011007f
C314 CS_BIAS.n27 GND 0.005906f
C315 CS_BIAS.t15 GND 0.351513f
C316 CS_BIAS.n28 GND 0.088545f
C317 CS_BIAS.t3 GND 0.010814f
C318 CS_BIAS.t7 GND 0.010814f
C319 CS_BIAS.n29 GND 0.069862f
C320 CS_BIAS.t2 GND 0.368705f
C321 CS_BIAS.t6 GND 0.359096f
C322 CS_BIAS.n30 GND 0.407887f
C323 CS_BIAS.n31 GND 0.364691f
C324 CS_BIAS.n32 GND 0.136657f
C325 CS_BIAS.n33 GND 0.005159f
C326 CS_BIAS.n34 GND 0.013517f
C327 CS_BIAS.n35 GND 0.011897f
C328 CS_BIAS.n36 GND 0.011007f
C329 CS_BIAS.n37 GND 0.005906f
C330 CS_BIAS.n38 GND 0.005906f
C331 CS_BIAS.n39 GND 0.005906f
C332 CS_BIAS.n40 GND 0.011007f
C333 CS_BIAS.n41 GND 0.010626f
C334 CS_BIAS.n42 GND 0.127991f
C335 CS_BIAS.n43 GND 0.07598f
C336 CS_BIAS.t8 GND 0.368705f
C337 CS_BIAS.t11 GND 0.359096f
C338 CS_BIAS.n44 GND 0.360451f
C339 CS_BIAS.n45 GND 0.084384f
C340 CS_BIAS.t14 GND 0.368705f
C341 CS_BIAS.t17 GND 0.359096f
C342 CS_BIAS.n46 GND 0.360451f
C343 CS_BIAS.n47 GND 0.062575f
C344 CS_BIAS.t23 GND 0.368705f
C345 CS_BIAS.t9 GND 0.359096f
C346 CS_BIAS.n48 GND 0.360451f
C347 CS_BIAS.n49 GND 0.110677f
C348 CS_BIAS.n50 GND 4.161241f
C349 VDD.t132 GND 0.012474f
C350 VDD.t138 GND 0.012474f
C351 VDD.n0 GND 0.061416f
C352 VDD.t140 GND 0.012474f
C353 VDD.t143 GND 0.012474f
C354 VDD.n1 GND 0.057167f
C355 VDD.n2 GND 0.705965f
C356 VDD.t158 GND 0.012474f
C357 VDD.t136 GND 0.012474f
C358 VDD.n3 GND 0.057167f
C359 VDD.n4 GND 0.369657f
C360 VDD.t129 GND 0.012474f
C361 VDD.t126 GND 0.012474f
C362 VDD.n5 GND 0.057167f
C363 VDD.n6 GND 0.307107f
C364 VDD.t160 GND 0.012474f
C365 VDD.t134 GND 0.012474f
C366 VDD.n7 GND 0.061416f
C367 VDD.t156 GND 0.012474f
C368 VDD.t152 GND 0.012474f
C369 VDD.n8 GND 0.057167f
C370 VDD.n9 GND 0.705965f
C371 VDD.t154 GND 0.012474f
C372 VDD.t148 GND 0.012474f
C373 VDD.n10 GND 0.057167f
C374 VDD.n11 GND 0.369657f
C375 VDD.t150 GND 0.012474f
C376 VDD.t145 GND 0.012474f
C377 VDD.n12 GND 0.057167f
C378 VDD.n13 GND 0.307107f
C379 VDD.n14 GND 0.245391f
C380 VDD.n15 GND 2.53232f
C381 VDD.t22 GND 0.02169f
C382 VDD.t168 GND 0.02169f
C383 VDD.n16 GND 0.103858f
C384 VDD.t10 GND 0.130827f
C385 VDD.n17 GND 0.5891f
C386 VDD.t5 GND 0.02169f
C387 VDD.t13 GND 0.02169f
C388 VDD.n18 GND 0.103858f
C389 VDD.t14 GND 0.130827f
C390 VDD.n19 GND 0.568033f
C391 VDD.n20 GND 0.27239f
C392 VDD.t16 GND 0.02169f
C393 VDD.t162 GND 0.02169f
C394 VDD.n21 GND 0.103858f
C395 VDD.t169 GND 0.130827f
C396 VDD.n22 GND 0.568033f
C397 VDD.n23 GND 0.192243f
C398 VDD.t23 GND 0.02169f
C399 VDD.t7 GND 0.02169f
C400 VDD.n24 GND 0.103858f
C401 VDD.t19 GND 0.130827f
C402 VDD.n25 GND 0.568033f
C403 VDD.n26 GND 0.192243f
C404 VDD.t20 GND 0.02169f
C405 VDD.t164 GND 0.02169f
C406 VDD.n27 GND 0.103858f
C407 VDD.t163 GND 0.130827f
C408 VDD.n28 GND 0.568033f
C409 VDD.n29 GND 0.243428f
C410 VDD.n30 GND 0.005307f
C411 VDD.n31 GND 0.005307f
C412 VDD.n32 GND 0.004287f
C413 VDD.n33 GND 0.004287f
C414 VDD.n34 GND 0.005326f
C415 VDD.n35 GND 0.005326f
C416 VDD.n36 GND 0.58089f
C417 VDD.n37 GND 0.58089f
C418 VDD.n38 GND 0.005326f
C419 VDD.n39 GND 0.005326f
C420 VDD.n40 GND 0.004287f
C421 VDD.n41 GND 0.005326f
C422 VDD.n42 GND 0.004287f
C423 VDD.n43 GND 0.005326f
C424 VDD.n44 GND 0.58089f
C425 VDD.n45 GND 0.005326f
C426 VDD.n46 GND 0.004287f
C427 VDD.n47 GND 0.005326f
C428 VDD.n48 GND 0.004287f
C429 VDD.n49 GND 0.005326f
C430 VDD.n50 GND 0.58089f
C431 VDD.n51 GND 0.005326f
C432 VDD.n52 GND 0.004287f
C433 VDD.n53 GND 0.005326f
C434 VDD.n54 GND 0.004287f
C435 VDD.n55 GND 0.005326f
C436 VDD.n56 GND 0.58089f
C437 VDD.n57 GND 0.005326f
C438 VDD.n58 GND 0.004287f
C439 VDD.n59 GND 0.005326f
C440 VDD.n60 GND 0.004287f
C441 VDD.n61 GND 0.005326f
C442 VDD.n62 GND 0.58089f
C443 VDD.n63 GND 0.005326f
C444 VDD.n64 GND 0.004287f
C445 VDD.n65 GND 0.005326f
C446 VDD.n66 GND 0.004287f
C447 VDD.n67 GND 0.005326f
C448 VDD.t4 GND 0.290445f
C449 VDD.n68 GND 0.005326f
C450 VDD.n69 GND 0.004287f
C451 VDD.n70 GND 0.005326f
C452 VDD.n71 GND 0.004287f
C453 VDD.n72 GND 0.005326f
C454 VDD.n73 GND 0.58089f
C455 VDD.n74 GND 0.005326f
C456 VDD.n75 GND 0.004287f
C457 VDD.n76 GND 0.005326f
C458 VDD.n77 GND 0.004287f
C459 VDD.n78 GND 0.005326f
C460 VDD.n79 GND 0.58089f
C461 VDD.n80 GND 0.005326f
C462 VDD.n81 GND 0.004287f
C463 VDD.n82 GND 0.005326f
C464 VDD.n83 GND 0.004287f
C465 VDD.n84 GND 0.005326f
C466 VDD.n85 GND 0.58089f
C467 VDD.n86 GND 0.005326f
C468 VDD.n87 GND 0.004287f
C469 VDD.n88 GND 0.005326f
C470 VDD.n89 GND 0.004287f
C471 VDD.n90 GND 0.005326f
C472 VDD.n91 GND 0.58089f
C473 VDD.n92 GND 0.005326f
C474 VDD.n93 GND 0.004287f
C475 VDD.n94 GND 0.005326f
C476 VDD.n95 GND 0.004287f
C477 VDD.n96 GND 0.005326f
C478 VDD.n97 GND 0.58089f
C479 VDD.n98 GND 0.005326f
C480 VDD.n99 GND 0.004287f
C481 VDD.n100 GND 0.005326f
C482 VDD.n101 GND 0.004287f
C483 VDD.n102 GND 0.005326f
C484 VDD.n103 GND 0.58089f
C485 VDD.n104 GND 0.005326f
C486 VDD.n105 GND 0.004287f
C487 VDD.n106 GND 0.005326f
C488 VDD.n107 GND 0.004287f
C489 VDD.n108 GND 0.005326f
C490 VDD.t50 GND 0.290445f
C491 VDD.n109 GND 0.005326f
C492 VDD.n110 GND 0.004287f
C493 VDD.n111 GND 0.005326f
C494 VDD.n112 GND 0.004287f
C495 VDD.n113 GND 0.005326f
C496 VDD.n114 GND 0.58089f
C497 VDD.n115 GND 0.511183f
C498 VDD.n116 GND 0.005326f
C499 VDD.n117 GND 0.004287f
C500 VDD.n118 GND 0.005326f
C501 VDD.n119 GND 0.004287f
C502 VDD.n120 GND 0.005326f
C503 VDD.n121 GND 0.58089f
C504 VDD.n122 GND 0.005326f
C505 VDD.n123 GND 0.004287f
C506 VDD.n124 GND 0.012553f
C507 VDD.n125 GND 0.012553f
C508 VDD.n126 GND 4.80687f
C509 VDD.n127 GND 0.012553f
C510 VDD.n128 GND 0.005326f
C511 VDD.n129 GND 0.004287f
C512 VDD.n131 GND 0.005326f
C513 VDD.n132 GND 0.005326f
C514 VDD.n133 GND 0.005326f
C515 VDD.n134 GND 0.004287f
C516 VDD.n135 GND 0.005326f
C517 VDD.n136 GND 0.005326f
C518 VDD.n137 GND 0.005326f
C519 VDD.n138 GND 0.005326f
C520 VDD.n139 GND 0.005326f
C521 VDD.n140 GND 0.004287f
C522 VDD.n141 GND 0.005326f
C523 VDD.n142 GND 0.005326f
C524 VDD.n143 GND 0.005326f
C525 VDD.n144 GND 0.005326f
C526 VDD.n145 GND 0.005326f
C527 VDD.n146 GND 0.004287f
C528 VDD.n147 GND 0.005326f
C529 VDD.n148 GND 0.005326f
C530 VDD.n149 GND 0.005326f
C531 VDD.t87 GND 0.159105f
C532 VDD.t85 GND 0.597454f
C533 VDD.n150 GND 0.084294f
C534 VDD.t86 GND 0.119732f
C535 VDD.n151 GND 0.085079f
C536 VDD.n152 GND 0.005326f
C537 VDD.n153 GND 0.005326f
C538 VDD.n154 GND 0.004287f
C539 VDD.n155 GND 0.005326f
C540 VDD.n156 GND 0.005326f
C541 VDD.n157 GND 0.005326f
C542 VDD.n158 GND 0.005326f
C543 VDD.n159 GND 0.005326f
C544 VDD.n160 GND 0.004287f
C545 VDD.n161 GND 0.005326f
C546 VDD.n162 GND 0.004287f
C547 VDD.n163 GND 0.003781f
C548 VDD.n164 GND 0.078438f
C549 VDD.n165 GND 0.004287f
C550 VDD.n167 GND 0.005326f
C551 VDD.n168 GND 0.005326f
C552 VDD.n169 GND 0.004287f
C553 VDD.n170 GND 0.005326f
C554 VDD.n171 GND 0.005326f
C555 VDD.n172 GND 0.005326f
C556 VDD.n173 GND 0.005326f
C557 VDD.n174 GND 0.005326f
C558 VDD.n175 GND 0.002208f
C559 VDD.n176 GND 0.005326f
C560 VDD.t66 GND 0.117451f
C561 VDD.t67 GND 0.160644f
C562 VDD.t65 GND 0.597454f
C563 VDD.n177 GND 0.084171f
C564 VDD.n178 GND 0.084531f
C565 VDD.n179 GND 0.007309f
C566 VDD.n180 GND 0.005326f
C567 VDD.n181 GND 0.005326f
C568 VDD.n182 GND 0.005326f
C569 VDD.n183 GND 0.005326f
C570 VDD.n184 GND 0.004287f
C571 VDD.n185 GND 0.005326f
C572 VDD.n186 GND 0.005326f
C573 VDD.n187 GND 0.005326f
C574 VDD.n188 GND 0.005326f
C575 VDD.n189 GND 0.005326f
C576 VDD.n190 GND 0.004287f
C577 VDD.n191 GND 0.005326f
C578 VDD.n192 GND 0.005326f
C579 VDD.n193 GND 0.005326f
C580 VDD.n194 GND 0.005326f
C581 VDD.n195 GND 0.005326f
C582 VDD.n196 GND 0.004287f
C583 VDD.n197 GND 0.005326f
C584 VDD.n198 GND 0.005326f
C585 VDD.n199 GND 0.005326f
C586 VDD.n200 GND 0.005326f
C587 VDD.n201 GND 0.005326f
C588 VDD.n202 GND 0.004287f
C589 VDD.n203 GND 0.005326f
C590 VDD.n204 GND 0.005326f
C591 VDD.n205 GND 0.005326f
C592 VDD.t52 GND 0.159105f
C593 VDD.t49 GND 0.597454f
C594 VDD.n206 GND 0.084294f
C595 VDD.t51 GND 0.119732f
C596 VDD.n207 GND 0.085079f
C597 VDD.n208 GND 0.005326f
C598 VDD.n209 GND 0.005326f
C599 VDD.n210 GND 0.004287f
C600 VDD.n211 GND 0.005326f
C601 VDD.n212 GND 0.005326f
C602 VDD.n213 GND 0.005326f
C603 VDD.n214 GND 0.005326f
C604 VDD.n215 GND 0.005326f
C605 VDD.n216 GND 0.004287f
C606 VDD.n217 GND 0.005326f
C607 VDD.n218 GND 0.005326f
C608 VDD.n219 GND 0.005326f
C609 VDD.n220 GND 0.003781f
C610 VDD.n225 GND 0.002716f
C611 VDD.n226 GND 0.003621f
C612 VDD.t27 GND 8.553611f
C613 VDD.t133 GND 7.73746f
C614 VDD.t159 GND 4.70812f
C615 VDD.n228 GND 1.66135f
C616 VDD.n229 GND 0.003621f
C617 VDD.t79 GND 0.087165f
C618 VDD.t78 GND 0.39322f
C619 VDD.n230 GND 0.070647f
C620 VDD.t80 GND 0.057758f
C621 VDD.n231 GND 0.070509f
C622 VDD.n232 GND 0.006279f
C623 VDD.n234 GND 0.003621f
C624 VDD.n235 GND 0.009566f
C625 VDD.n237 GND 0.003621f
C626 VDD.n238 GND 0.395005f
C627 VDD.n239 GND 0.009198f
C628 VDD.n240 GND 0.009198f
C629 VDD.n241 GND 0.003621f
C630 VDD.n242 GND 0.009548f
C631 VDD.n243 GND 0.003621f
C632 VDD.n244 GND 0.003621f
C633 VDD.n246 GND 0.003621f
C634 VDD.n247 GND 0.003621f
C635 VDD.n249 GND 0.003621f
C636 VDD.n250 GND 0.003621f
C637 VDD.n252 GND 0.003621f
C638 VDD.t31 GND 0.087165f
C639 VDD.t29 GND 0.39322f
C640 VDD.n253 GND 0.070647f
C641 VDD.t32 GND 0.057758f
C642 VDD.n254 GND 0.070509f
C643 VDD.n255 GND 0.003621f
C644 VDD.n257 GND 0.003621f
C645 VDD.n258 GND 0.003621f
C646 VDD.n259 GND 0.395005f
C647 VDD.n260 GND 0.003621f
C648 VDD.n261 GND 0.003621f
C649 VDD.n262 GND 0.003621f
C650 VDD.n263 GND 0.003621f
C651 VDD.n264 GND 0.003621f
C652 VDD.n265 GND 0.395005f
C653 VDD.n266 GND 0.003621f
C654 VDD.n267 GND 0.003621f
C655 VDD.n268 GND 0.003621f
C656 VDD.n269 GND 0.003621f
C657 VDD.n270 GND 0.003621f
C658 VDD.n271 GND 0.003621f
C659 VDD.n272 GND 0.395005f
C660 VDD.n273 GND 0.003621f
C661 VDD.n274 GND 0.003621f
C662 VDD.n275 GND 0.003621f
C663 VDD.n276 GND 0.003621f
C664 VDD.n277 GND 0.003621f
C665 VDD.n278 GND 0.214929f
C666 VDD.n279 GND 0.003621f
C667 VDD.n280 GND 0.003621f
C668 VDD.n281 GND 0.003621f
C669 VDD.n282 GND 0.003621f
C670 VDD.n283 GND 0.003621f
C671 VDD.t30 GND 0.197503f
C672 VDD.n284 GND 0.003621f
C673 VDD.n285 GND 0.003621f
C674 VDD.t151 GND 0.197503f
C675 VDD.n286 GND 0.003621f
C676 VDD.n287 GND 0.003621f
C677 VDD.n288 GND 0.003621f
C678 VDD.n289 GND 0.395005f
C679 VDD.n290 GND 0.003621f
C680 VDD.n291 GND 0.003621f
C681 VDD.n292 GND 0.380483f
C682 VDD.n293 GND 0.003621f
C683 VDD.n294 GND 0.003621f
C684 VDD.n295 GND 0.003621f
C685 VDD.n296 GND 0.395005f
C686 VDD.n297 GND 0.003621f
C687 VDD.n298 GND 0.003621f
C688 VDD.n299 GND 0.003621f
C689 VDD.n300 GND 0.003621f
C690 VDD.n301 GND 0.003621f
C691 VDD.n302 GND 0.395005f
C692 VDD.n303 GND 0.003621f
C693 VDD.n304 GND 0.003621f
C694 VDD.n305 GND 0.003621f
C695 VDD.n306 GND 0.003621f
C696 VDD.n307 GND 0.003621f
C697 VDD.n308 GND 0.395005f
C698 VDD.n309 GND 0.003621f
C699 VDD.n310 GND 0.003621f
C700 VDD.n311 GND 0.003621f
C701 VDD.n312 GND 0.003621f
C702 VDD.n313 GND 0.003621f
C703 VDD.n314 GND 0.395005f
C704 VDD.n315 GND 0.003621f
C705 VDD.n316 GND 0.003621f
C706 VDD.n317 GND 0.003621f
C707 VDD.n318 GND 0.003621f
C708 VDD.n319 GND 0.003621f
C709 VDD.n320 GND 0.395005f
C710 VDD.n321 GND 0.003621f
C711 VDD.n322 GND 0.003621f
C712 VDD.n323 GND 0.003621f
C713 VDD.n324 GND 0.003621f
C714 VDD.n325 GND 0.003621f
C715 VDD.n326 GND 0.395005f
C716 VDD.n327 GND 0.003621f
C717 VDD.n328 GND 0.003621f
C718 VDD.n329 GND 0.003621f
C719 VDD.n330 GND 0.003621f
C720 VDD.n331 GND 0.003621f
C721 VDD.t155 GND 0.197503f
C722 VDD.n332 GND 0.003621f
C723 VDD.n333 GND 0.003621f
C724 VDD.n334 GND 0.003621f
C725 VDD.n335 GND 0.003621f
C726 VDD.n336 GND 0.003621f
C727 VDD.n337 GND 0.395005f
C728 VDD.n338 GND 0.003621f
C729 VDD.n339 GND 0.003621f
C730 VDD.n340 GND 0.278827f
C731 VDD.n341 GND 0.003621f
C732 VDD.n342 GND 0.003621f
C733 VDD.n343 GND 0.003621f
C734 VDD.n344 GND 0.34563f
C735 VDD.n345 GND 0.003621f
C736 VDD.n346 GND 0.003621f
C737 VDD.n347 GND 0.003621f
C738 VDD.n348 GND 0.003621f
C739 VDD.n349 GND 0.003621f
C740 VDD.n350 GND 0.395005f
C741 VDD.n351 GND 0.003621f
C742 VDD.n352 GND 0.003621f
C743 VDD.t127 GND 0.197503f
C744 VDD.n353 GND 0.003621f
C745 VDD.n354 GND 0.003621f
C746 VDD.n355 GND 0.003621f
C747 VDD.n356 GND 0.395005f
C748 VDD.n357 GND 0.003621f
C749 VDD.n358 GND 0.003621f
C750 VDD.n359 GND 0.003621f
C751 VDD.n360 GND 0.003621f
C752 VDD.n361 GND 0.003621f
C753 VDD.n362 GND 0.395005f
C754 VDD.n363 GND 0.003621f
C755 VDD.n364 GND 0.003621f
C756 VDD.n365 GND 0.003621f
C757 VDD.n366 GND 0.003621f
C758 VDD.n367 GND 0.003621f
C759 VDD.n368 GND 0.395005f
C760 VDD.n369 GND 0.003621f
C761 VDD.n370 GND 0.003621f
C762 VDD.n371 GND 0.003621f
C763 VDD.n372 GND 0.003621f
C764 VDD.n373 GND 0.003621f
C765 VDD.n374 GND 0.395005f
C766 VDD.n375 GND 0.003621f
C767 VDD.n376 GND 0.003621f
C768 VDD.n377 GND 0.003621f
C769 VDD.n378 GND 0.003621f
C770 VDD.n379 GND 0.003621f
C771 VDD.n380 GND 0.395005f
C772 VDD.n381 GND 0.003621f
C773 VDD.n382 GND 0.003621f
C774 VDD.n383 GND 0.003621f
C775 VDD.n384 GND 0.003621f
C776 VDD.n385 GND 0.003621f
C777 VDD.n386 GND 0.395005f
C778 VDD.n387 GND 0.003621f
C779 VDD.n388 GND 0.003621f
C780 VDD.n389 GND 0.003621f
C781 VDD.n390 GND 0.003621f
C782 VDD.n391 GND 0.003621f
C783 VDD.n392 GND 0.395005f
C784 VDD.n393 GND 0.003621f
C785 VDD.n394 GND 0.003621f
C786 VDD.n395 GND 0.003621f
C787 VDD.n396 GND 0.003621f
C788 VDD.n397 GND 0.003621f
C789 VDD.n398 GND 0.246878f
C790 VDD.n399 GND 0.003621f
C791 VDD.n400 GND 0.003621f
C792 VDD.n401 GND 0.003621f
C793 VDD.n402 GND 0.003621f
C794 VDD.n403 GND 0.003621f
C795 VDD.n404 GND 0.395005f
C796 VDD.n405 GND 0.003621f
C797 VDD.n406 GND 0.003621f
C798 VDD.t123 GND 0.197503f
C799 VDD.n407 GND 0.003621f
C800 VDD.n408 GND 0.003621f
C801 VDD.n409 GND 0.003621f
C802 VDD.t147 GND 0.197503f
C803 VDD.n410 GND 0.003621f
C804 VDD.n411 GND 0.003621f
C805 VDD.n412 GND 0.003621f
C806 VDD.n413 GND 0.003621f
C807 VDD.n414 GND 0.003621f
C808 VDD.n415 GND 0.395005f
C809 VDD.n416 GND 0.003621f
C810 VDD.n417 GND 0.003621f
C811 VDD.n418 GND 0.29335f
C812 VDD.n419 GND 0.003621f
C813 VDD.n420 GND 0.003621f
C814 VDD.n421 GND 0.003621f
C815 VDD.n422 GND 0.395005f
C816 VDD.n423 GND 0.003621f
C817 VDD.n424 GND 0.003621f
C818 VDD.n425 GND 0.003621f
C819 VDD.n426 GND 0.003621f
C820 VDD.n427 GND 0.003621f
C821 VDD.n428 GND 0.395005f
C822 VDD.n429 GND 0.003621f
C823 VDD.n430 GND 0.003621f
C824 VDD.n431 GND 0.003621f
C825 VDD.n432 GND 0.003621f
C826 VDD.n433 GND 0.003621f
C827 VDD.n434 GND 0.395005f
C828 VDD.n435 GND 0.003621f
C829 VDD.n436 GND 0.003621f
C830 VDD.n437 GND 0.003621f
C831 VDD.n438 GND 0.003621f
C832 VDD.n439 GND 0.003621f
C833 VDD.n440 GND 0.395005f
C834 VDD.n441 GND 0.003621f
C835 VDD.n442 GND 0.003621f
C836 VDD.n443 GND 0.003621f
C837 VDD.n444 GND 0.003621f
C838 VDD.n445 GND 0.003621f
C839 VDD.n446 GND 0.395005f
C840 VDD.n447 GND 0.003621f
C841 VDD.n448 GND 0.003621f
C842 VDD.n449 GND 0.003621f
C843 VDD.n450 GND 0.003621f
C844 VDD.n451 GND 0.003621f
C845 VDD.t121 GND 0.197503f
C846 VDD.n452 GND 0.003621f
C847 VDD.n453 GND 0.003621f
C848 VDD.n454 GND 0.003621f
C849 VDD.n455 GND 0.003621f
C850 VDD.n456 GND 0.003621f
C851 VDD.n457 GND 0.395005f
C852 VDD.n458 GND 0.003621f
C853 VDD.n459 GND 0.003621f
C854 VDD.n460 GND 0.246878f
C855 VDD.n461 GND 0.003621f
C856 VDD.n462 GND 0.003621f
C857 VDD.n463 GND 0.003621f
C858 VDD.t153 GND 0.197503f
C859 VDD.n464 GND 0.003621f
C860 VDD.n465 GND 0.003621f
C861 VDD.n466 GND 0.003621f
C862 VDD.n467 GND 0.003621f
C863 VDD.n468 GND 0.003621f
C864 VDD.n469 GND 0.395005f
C865 VDD.n470 GND 0.003621f
C866 VDD.n471 GND 0.003621f
C867 VDD.n472 GND 0.392101f
C868 VDD.n473 GND 0.003621f
C869 VDD.n474 GND 0.003621f
C870 VDD.n475 GND 0.003621f
C871 VDD.n476 GND 0.395005f
C872 VDD.n477 GND 0.003621f
C873 VDD.n478 GND 0.003621f
C874 VDD.n479 GND 0.003621f
C875 VDD.n480 GND 0.003621f
C876 VDD.n481 GND 0.003621f
C877 VDD.n482 GND 0.395005f
C878 VDD.n483 GND 0.003621f
C879 VDD.n484 GND 0.003621f
C880 VDD.n485 GND 0.003621f
C881 VDD.n486 GND 0.003621f
C882 VDD.n487 GND 0.003621f
C883 VDD.n488 GND 0.395005f
C884 VDD.n489 GND 0.003621f
C885 VDD.n490 GND 0.003621f
C886 VDD.n491 GND 0.003621f
C887 VDD.n492 GND 0.003621f
C888 VDD.n493 GND 0.003621f
C889 VDD.n494 GND 0.395005f
C890 VDD.n495 GND 0.003621f
C891 VDD.n496 GND 0.003621f
C892 VDD.n497 GND 0.003621f
C893 VDD.n498 GND 0.003621f
C894 VDD.n499 GND 0.003621f
C895 VDD.n500 GND 0.395005f
C896 VDD.n501 GND 0.003621f
C897 VDD.n502 GND 0.003621f
C898 VDD.n503 GND 0.003621f
C899 VDD.n504 GND 0.003621f
C900 VDD.n505 GND 0.003621f
C901 VDD.t122 GND 0.197503f
C902 VDD.n506 GND 0.003621f
C903 VDD.n507 GND 0.003621f
C904 VDD.n508 GND 0.003621f
C905 VDD.n509 GND 0.003621f
C906 VDD.n510 GND 0.003621f
C907 VDD.n511 GND 0.299158f
C908 VDD.n512 GND 0.003621f
C909 VDD.n513 GND 0.003621f
C910 VDD.n514 GND 0.34563f
C911 VDD.n515 GND 0.003621f
C912 VDD.n516 GND 0.003621f
C913 VDD.n517 GND 0.003621f
C914 VDD.n518 GND 0.395005f
C915 VDD.n519 GND 0.003621f
C916 VDD.n520 GND 0.003621f
C917 VDD.t144 GND 0.197503f
C918 VDD.n521 GND 0.003621f
C919 VDD.n522 GND 0.003621f
C920 VDD.n523 GND 0.003621f
C921 VDD.n524 GND 0.395005f
C922 VDD.n525 GND 0.003621f
C923 VDD.n526 GND 0.003621f
C924 VDD.n527 GND 0.003621f
C925 VDD.n528 GND 0.003621f
C926 VDD.n529 GND 0.003621f
C927 VDD.n530 GND 0.395005f
C928 VDD.n531 GND 0.003621f
C929 VDD.n532 GND 0.003621f
C930 VDD.n533 GND 0.003621f
C931 VDD.n534 GND 0.003621f
C932 VDD.n535 GND 0.003621f
C933 VDD.n536 GND 0.395005f
C934 VDD.n537 GND 0.003621f
C935 VDD.n538 GND 0.003621f
C936 VDD.n539 GND 0.003621f
C937 VDD.n540 GND 0.003621f
C938 VDD.n541 GND 0.003621f
C939 VDD.n542 GND 0.395005f
C940 VDD.n543 GND 0.003621f
C941 VDD.n544 GND 0.003621f
C942 VDD.n545 GND 0.003621f
C943 VDD.n546 GND 0.003621f
C944 VDD.n547 GND 0.003621f
C945 VDD.n548 GND 0.395005f
C946 VDD.n549 GND 0.003621f
C947 VDD.n550 GND 0.003621f
C948 VDD.n551 GND 0.003621f
C949 VDD.n552 GND 0.003621f
C950 VDD.n553 GND 0.003621f
C951 VDD.n554 GND 0.395005f
C952 VDD.n555 GND 0.003621f
C953 VDD.n556 GND 0.003621f
C954 VDD.n557 GND 0.003621f
C955 VDD.n558 GND 0.003621f
C956 VDD.n559 GND 0.003621f
C957 VDD.n560 GND 0.395005f
C958 VDD.n561 GND 0.003621f
C959 VDD.n562 GND 0.003621f
C960 VDD.n563 GND 0.003621f
C961 VDD.n564 GND 0.003621f
C962 VDD.n565 GND 0.003621f
C963 VDD.n566 GND 0.200407f
C964 VDD.n567 GND 0.003621f
C965 VDD.n568 GND 0.003621f
C966 VDD.n569 GND 0.003621f
C967 VDD.n570 GND 0.003621f
C968 VDD.n571 GND 0.003621f
C969 VDD.n572 GND 0.395005f
C970 VDD.n573 GND 0.003621f
C971 VDD.n574 GND 0.003621f
C972 VDD.t149 GND 0.18298f
C973 VDD.t69 GND 0.194598f
C974 VDD.n575 GND 0.003621f
C975 VDD.n576 GND 0.003621f
C976 VDD.n577 GND 0.003621f
C977 VDD.n578 GND 0.395005f
C978 VDD.n579 GND 0.003621f
C979 VDD.n580 GND 0.003621f
C980 VDD.n581 GND 0.003621f
C981 VDD.n582 GND 0.003621f
C982 VDD.n583 GND 0.003621f
C983 VDD.n584 GND 0.395005f
C984 VDD.n585 GND 0.003621f
C985 VDD.n586 GND 0.003621f
C986 VDD.n587 GND 0.003621f
C987 VDD.n588 GND 0.003621f
C988 VDD.n589 GND 0.003621f
C989 VDD.n590 GND 0.395005f
C990 VDD.n591 GND 0.003621f
C991 VDD.n592 GND 0.003621f
C992 VDD.n593 GND 0.003621f
C993 VDD.n594 GND 0.003621f
C994 VDD.n595 GND 0.003621f
C995 VDD.n596 GND 0.395005f
C996 VDD.n597 GND 0.003621f
C997 VDD.n598 GND 0.003621f
C998 VDD.n599 GND 0.003621f
C999 VDD.n600 GND 0.009548f
C1000 VDD.n601 GND 0.009548f
C1001 VDD.n602 GND 0.60703f
C1002 VDD.n620 GND 0.009548f
C1003 VDD.n621 GND 0.009198f
C1004 VDD.n622 GND 0.003621f
C1005 VDD.n623 GND 0.009198f
C1006 VDD.t116 GND 0.087165f
C1007 VDD.t115 GND 0.39322f
C1008 VDD.n624 GND 0.070647f
C1009 VDD.t117 GND 0.057758f
C1010 VDD.n625 GND 0.070509f
C1011 VDD.n626 GND 0.003621f
C1012 VDD.n627 GND 0.003621f
C1013 VDD.n628 GND 0.395005f
C1014 VDD.n629 GND 0.003621f
C1015 VDD.n630 GND 0.003621f
C1016 VDD.n631 GND 0.003621f
C1017 VDD.n632 GND 0.009198f
C1018 VDD.n633 GND 0.003621f
C1019 VDD.t83 GND 0.087165f
C1020 VDD.t81 GND 0.39322f
C1021 VDD.n634 GND 0.070647f
C1022 VDD.t84 GND 0.057758f
C1023 VDD.n635 GND 0.070509f
C1024 VDD.n636 GND 0.003621f
C1025 VDD.n637 GND 0.003621f
C1026 VDD.n638 GND 0.395005f
C1027 VDD.n639 GND 0.003621f
C1028 VDD.n640 GND 0.003621f
C1029 VDD.n641 GND 0.003621f
C1030 VDD.n642 GND 0.003621f
C1031 VDD.n643 GND 0.003621f
C1032 VDD.n644 GND 0.395005f
C1033 VDD.n645 GND 0.003621f
C1034 VDD.n646 GND 0.003621f
C1035 VDD.n647 GND 0.003621f
C1036 VDD.n648 GND 0.003621f
C1037 VDD.n649 GND 0.003621f
C1038 VDD.n650 GND 0.003621f
C1039 VDD.n651 GND 0.395005f
C1040 VDD.n652 GND 0.003621f
C1041 VDD.n653 GND 0.003621f
C1042 VDD.n654 GND 0.003621f
C1043 VDD.n655 GND 0.003621f
C1044 VDD.n656 GND 0.003621f
C1045 VDD.n657 GND 0.212025f
C1046 VDD.n658 GND 0.003621f
C1047 VDD.n659 GND 0.003621f
C1048 VDD.n660 GND 0.003621f
C1049 VDD.n661 GND 0.003621f
C1050 VDD.n662 GND 0.003621f
C1051 VDD.n663 GND 0.395005f
C1052 VDD.n664 GND 0.003621f
C1053 VDD.n665 GND 0.003621f
C1054 VDD.t82 GND 0.194598f
C1055 VDD.t125 GND 0.18298f
C1056 VDD.n666 GND 0.003621f
C1057 VDD.n667 GND 0.003621f
C1058 VDD.n668 GND 0.003621f
C1059 VDD.n669 GND 0.395005f
C1060 VDD.n670 GND 0.003621f
C1061 VDD.n671 GND 0.003621f
C1062 VDD.n672 GND 0.003621f
C1063 VDD.n673 GND 0.003621f
C1064 VDD.n674 GND 0.003621f
C1065 VDD.n675 GND 0.395005f
C1066 VDD.n676 GND 0.003621f
C1067 VDD.n677 GND 0.003621f
C1068 VDD.n678 GND 0.003621f
C1069 VDD.n679 GND 0.003621f
C1070 VDD.n680 GND 0.003621f
C1071 VDD.n681 GND 0.395005f
C1072 VDD.n682 GND 0.003621f
C1073 VDD.n683 GND 0.003621f
C1074 VDD.n684 GND 0.003621f
C1075 VDD.n685 GND 0.003621f
C1076 VDD.n686 GND 0.003621f
C1077 VDD.n687 GND 0.395005f
C1078 VDD.n688 GND 0.003621f
C1079 VDD.n689 GND 0.003621f
C1080 VDD.n690 GND 0.003621f
C1081 VDD.n691 GND 0.003621f
C1082 VDD.n692 GND 0.003621f
C1083 VDD.n693 GND 0.395005f
C1084 VDD.n694 GND 0.003621f
C1085 VDD.n695 GND 0.003621f
C1086 VDD.n696 GND 0.003621f
C1087 VDD.n697 GND 0.003621f
C1088 VDD.n698 GND 0.003621f
C1089 VDD.n699 GND 0.395005f
C1090 VDD.n700 GND 0.003621f
C1091 VDD.n701 GND 0.003621f
C1092 VDD.n702 GND 0.003621f
C1093 VDD.n703 GND 0.003621f
C1094 VDD.n704 GND 0.003621f
C1095 VDD.n705 GND 0.395005f
C1096 VDD.n706 GND 0.003621f
C1097 VDD.n707 GND 0.003621f
C1098 VDD.n708 GND 0.003621f
C1099 VDD.n709 GND 0.003621f
C1100 VDD.n710 GND 0.003621f
C1101 VDD.n711 GND 0.29335f
C1102 VDD.n712 GND 0.003621f
C1103 VDD.n713 GND 0.003621f
C1104 VDD.n714 GND 0.003621f
C1105 VDD.n715 GND 0.003621f
C1106 VDD.n716 GND 0.003621f
C1107 VDD.n717 GND 0.395005f
C1108 VDD.n718 GND 0.003621f
C1109 VDD.n719 GND 0.003621f
C1110 VDD.t128 GND 0.197503f
C1111 VDD.n720 GND 0.003621f
C1112 VDD.n721 GND 0.003621f
C1113 VDD.n722 GND 0.003621f
C1114 VDD.t130 GND 0.197503f
C1115 VDD.n723 GND 0.003621f
C1116 VDD.n724 GND 0.003621f
C1117 VDD.n725 GND 0.003621f
C1118 VDD.n726 GND 0.003621f
C1119 VDD.n727 GND 0.003621f
C1120 VDD.n728 GND 0.395005f
C1121 VDD.n729 GND 0.003621f
C1122 VDD.n730 GND 0.003621f
C1123 VDD.n731 GND 0.246878f
C1124 VDD.n732 GND 0.003621f
C1125 VDD.n733 GND 0.003621f
C1126 VDD.n734 GND 0.003621f
C1127 VDD.n735 GND 0.395005f
C1128 VDD.n736 GND 0.003621f
C1129 VDD.n737 GND 0.003621f
C1130 VDD.n738 GND 0.003621f
C1131 VDD.n739 GND 0.003621f
C1132 VDD.n740 GND 0.003621f
C1133 VDD.n741 GND 0.395005f
C1134 VDD.n742 GND 0.003621f
C1135 VDD.n743 GND 0.003621f
C1136 VDD.n744 GND 0.003621f
C1137 VDD.n745 GND 0.003621f
C1138 VDD.n746 GND 0.003621f
C1139 VDD.n747 GND 0.395005f
C1140 VDD.n748 GND 0.003621f
C1141 VDD.n749 GND 0.003621f
C1142 VDD.n750 GND 0.003621f
C1143 VDD.n751 GND 0.003621f
C1144 VDD.n752 GND 0.003621f
C1145 VDD.n753 GND 0.395005f
C1146 VDD.n754 GND 0.003621f
C1147 VDD.n755 GND 0.003621f
C1148 VDD.n756 GND 0.003621f
C1149 VDD.n757 GND 0.003621f
C1150 VDD.n758 GND 0.003621f
C1151 VDD.n759 GND 0.395005f
C1152 VDD.n760 GND 0.003621f
C1153 VDD.n761 GND 0.003621f
C1154 VDD.n762 GND 0.003621f
C1155 VDD.n763 GND 0.003621f
C1156 VDD.n764 GND 0.003621f
C1157 VDD.t135 GND 0.197503f
C1158 VDD.n765 GND 0.003621f
C1159 VDD.n766 GND 0.003621f
C1160 VDD.n767 GND 0.003621f
C1161 VDD.n768 GND 0.003621f
C1162 VDD.n769 GND 0.003621f
C1163 VDD.n770 GND 0.395005f
C1164 VDD.n771 GND 0.003621f
C1165 VDD.n772 GND 0.003621f
C1166 VDD.n773 GND 0.200407f
C1167 VDD.n774 GND 0.003621f
C1168 VDD.n775 GND 0.003621f
C1169 VDD.n776 GND 0.003621f
C1170 VDD.t146 GND 0.197503f
C1171 VDD.n777 GND 0.003621f
C1172 VDD.n778 GND 0.003621f
C1173 VDD.n779 GND 0.003621f
C1174 VDD.n780 GND 0.003621f
C1175 VDD.n781 GND 0.003621f
C1176 VDD.n782 GND 0.395005f
C1177 VDD.n783 GND 0.003621f
C1178 VDD.n784 GND 0.003621f
C1179 VDD.n785 GND 0.34563f
C1180 VDD.n786 GND 0.003621f
C1181 VDD.n787 GND 0.003621f
C1182 VDD.n788 GND 0.003621f
C1183 VDD.n789 GND 0.395005f
C1184 VDD.n790 GND 0.003621f
C1185 VDD.n791 GND 0.003621f
C1186 VDD.n792 GND 0.003621f
C1187 VDD.n793 GND 0.003621f
C1188 VDD.n794 GND 0.003621f
C1189 VDD.n795 GND 0.395005f
C1190 VDD.n796 GND 0.003621f
C1191 VDD.n797 GND 0.003621f
C1192 VDD.n798 GND 0.003621f
C1193 VDD.n799 GND 0.003621f
C1194 VDD.n800 GND 0.003621f
C1195 VDD.n801 GND 0.395005f
C1196 VDD.n802 GND 0.003621f
C1197 VDD.n803 GND 0.003621f
C1198 VDD.n804 GND 0.003621f
C1199 VDD.n805 GND 0.003621f
C1200 VDD.n806 GND 0.003621f
C1201 VDD.n807 GND 0.395005f
C1202 VDD.n808 GND 0.003621f
C1203 VDD.n809 GND 0.003621f
C1204 VDD.n810 GND 0.003621f
C1205 VDD.n811 GND 0.003621f
C1206 VDD.n812 GND 0.003621f
C1207 VDD.n813 GND 0.395005f
C1208 VDD.n814 GND 0.003621f
C1209 VDD.n815 GND 0.003621f
C1210 VDD.n816 GND 0.003621f
C1211 VDD.n817 GND 0.003621f
C1212 VDD.n818 GND 0.003621f
C1213 VDD.t157 GND 0.197503f
C1214 VDD.n819 GND 0.003621f
C1215 VDD.n820 GND 0.003621f
C1216 VDD.n821 GND 0.003621f
C1217 VDD.n822 GND 0.003621f
C1218 VDD.n823 GND 0.003621f
C1219 VDD.n824 GND 0.34563f
C1220 VDD.n825 GND 0.003621f
C1221 VDD.n826 GND 0.003621f
C1222 VDD.n827 GND 0.299158f
C1223 VDD.n828 GND 0.003621f
C1224 VDD.n829 GND 0.003621f
C1225 VDD.n830 GND 0.003621f
C1226 VDD.n831 GND 0.395005f
C1227 VDD.n832 GND 0.003621f
C1228 VDD.n833 GND 0.003621f
C1229 VDD.t141 GND 0.197503f
C1230 VDD.n834 GND 0.003621f
C1231 VDD.n835 GND 0.003621f
C1232 VDD.n836 GND 0.003621f
C1233 VDD.n837 GND 0.395005f
C1234 VDD.n838 GND 0.003621f
C1235 VDD.n839 GND 0.003621f
C1236 VDD.n840 GND 0.003621f
C1237 VDD.n841 GND 0.003621f
C1238 VDD.n842 GND 0.003621f
C1239 VDD.n843 GND 0.395005f
C1240 VDD.n844 GND 0.003621f
C1241 VDD.n845 GND 0.003621f
C1242 VDD.n846 GND 0.003621f
C1243 VDD.n847 GND 0.003621f
C1244 VDD.n848 GND 0.003621f
C1245 VDD.n849 GND 0.395005f
C1246 VDD.n850 GND 0.003621f
C1247 VDD.n851 GND 0.003621f
C1248 VDD.n852 GND 0.003621f
C1249 VDD.n853 GND 0.003621f
C1250 VDD.n854 GND 0.003621f
C1251 VDD.n855 GND 0.395005f
C1252 VDD.n856 GND 0.003621f
C1253 VDD.n857 GND 0.003621f
C1254 VDD.n858 GND 0.003621f
C1255 VDD.n859 GND 0.003621f
C1256 VDD.n860 GND 0.003621f
C1257 VDD.n861 GND 0.395005f
C1258 VDD.n862 GND 0.003621f
C1259 VDD.n863 GND 0.003621f
C1260 VDD.n864 GND 0.003621f
C1261 VDD.n865 GND 0.003621f
C1262 VDD.n866 GND 0.003621f
C1263 VDD.n867 GND 0.395005f
C1264 VDD.n868 GND 0.003621f
C1265 VDD.n869 GND 0.003621f
C1266 VDD.n870 GND 0.003621f
C1267 VDD.n871 GND 0.003621f
C1268 VDD.n872 GND 0.003621f
C1269 VDD.n873 GND 0.395005f
C1270 VDD.n874 GND 0.003621f
C1271 VDD.n875 GND 0.003621f
C1272 VDD.n876 GND 0.003621f
C1273 VDD.n877 GND 0.003621f
C1274 VDD.n878 GND 0.003621f
C1275 VDD.n879 GND 0.246878f
C1276 VDD.n880 GND 0.003621f
C1277 VDD.n881 GND 0.003621f
C1278 VDD.n882 GND 0.003621f
C1279 VDD.n883 GND 0.003621f
C1280 VDD.n884 GND 0.003621f
C1281 VDD.n885 GND 0.395005f
C1282 VDD.n886 GND 0.003621f
C1283 VDD.n887 GND 0.003621f
C1284 VDD.t124 GND 0.197503f
C1285 VDD.n888 GND 0.003621f
C1286 VDD.n889 GND 0.003621f
C1287 VDD.n890 GND 0.003621f
C1288 VDD.n891 GND 0.395005f
C1289 VDD.n892 GND 0.003621f
C1290 VDD.n893 GND 0.003621f
C1291 VDD.n894 GND 0.003621f
C1292 VDD.n895 GND 0.003621f
C1293 VDD.n896 GND 0.003621f
C1294 VDD.t142 GND 0.197503f
C1295 VDD.n897 GND 0.003621f
C1296 VDD.n898 GND 0.003621f
C1297 VDD.n899 GND 0.003621f
C1298 VDD.n900 GND 0.003621f
C1299 VDD.n901 GND 0.003621f
C1300 VDD.n902 GND 0.395005f
C1301 VDD.n903 GND 0.003621f
C1302 VDD.n904 GND 0.003621f
C1303 VDD.n905 GND 0.313681f
C1304 VDD.n906 GND 0.003621f
C1305 VDD.n907 GND 0.003621f
C1306 VDD.n908 GND 0.003621f
C1307 VDD.n909 GND 0.395005f
C1308 VDD.n910 GND 0.003621f
C1309 VDD.n911 GND 0.003621f
C1310 VDD.n912 GND 0.003621f
C1311 VDD.n913 GND 0.003621f
C1312 VDD.n914 GND 0.003621f
C1313 VDD.n915 GND 0.395005f
C1314 VDD.n916 GND 0.003621f
C1315 VDD.n917 GND 0.003621f
C1316 VDD.n918 GND 0.003621f
C1317 VDD.n919 GND 0.003621f
C1318 VDD.n920 GND 0.003621f
C1319 VDD.n921 GND 0.395005f
C1320 VDD.n922 GND 0.003621f
C1321 VDD.n923 GND 0.003621f
C1322 VDD.n924 GND 0.003621f
C1323 VDD.n925 GND 0.003621f
C1324 VDD.n926 GND 0.003621f
C1325 VDD.n927 GND 0.395005f
C1326 VDD.n928 GND 0.003621f
C1327 VDD.n929 GND 0.003621f
C1328 VDD.n930 GND 0.003621f
C1329 VDD.n931 GND 0.003621f
C1330 VDD.n932 GND 0.003621f
C1331 VDD.n933 GND 0.395005f
C1332 VDD.n934 GND 0.003621f
C1333 VDD.n935 GND 0.003621f
C1334 VDD.n936 GND 0.003621f
C1335 VDD.n937 GND 0.003621f
C1336 VDD.n938 GND 0.003621f
C1337 VDD.n939 GND 0.395005f
C1338 VDD.n940 GND 0.003621f
C1339 VDD.n941 GND 0.003621f
C1340 VDD.n942 GND 0.003621f
C1341 VDD.n943 GND 0.003621f
C1342 VDD.n944 GND 0.003621f
C1343 VDD.t46 GND 0.197503f
C1344 VDD.n945 GND 0.003621f
C1345 VDD.n946 GND 0.003621f
C1346 VDD.n947 GND 0.003621f
C1347 VDD.n948 GND 0.003621f
C1348 VDD.n949 GND 0.003621f
C1349 VDD.n950 GND 0.395005f
C1350 VDD.n951 GND 0.003621f
C1351 VDD.n952 GND 0.003621f
C1352 VDD.t139 GND 0.197503f
C1353 VDD.n953 GND 0.003621f
C1354 VDD.n954 GND 0.003621f
C1355 VDD.n955 GND 0.003621f
C1356 VDD.n956 GND 0.395005f
C1357 VDD.n957 GND 0.003621f
C1358 VDD.n958 GND 0.003621f
C1359 VDD.n959 GND 0.003621f
C1360 VDD.n960 GND 0.003621f
C1361 VDD.n961 GND 0.003621f
C1362 VDD.n962 GND 0.395005f
C1363 VDD.n963 GND 0.003621f
C1364 VDD.n964 GND 0.003621f
C1365 VDD.n965 GND 0.003621f
C1366 VDD.n966 GND 0.003621f
C1367 VDD.n967 GND 0.003621f
C1368 VDD.n968 GND 0.395005f
C1369 VDD.n969 GND 0.003621f
C1370 VDD.n970 GND 0.003621f
C1371 VDD.n971 GND 0.003621f
C1372 VDD.n972 GND 0.009198f
C1373 VDD.n973 GND 0.009198f
C1374 VDD.n974 GND 0.60703f
C1375 VDD.n975 GND 0.003621f
C1376 VDD.n976 GND 0.003621f
C1377 VDD.n977 GND 0.009198f
C1378 VDD.n978 GND 0.003621f
C1379 VDD.n979 GND 0.003621f
C1380 VDD.t137 GND 4.70812f
C1381 VDD.n987 GND 0.009548f
C1382 VDD.n996 GND 0.009548f
C1383 VDD.n997 GND 0.009548f
C1384 VDD.n998 GND 0.003621f
C1385 VDD.n999 GND 0.080335f
C1386 VDD.t111 GND 0.087165f
C1387 VDD.t109 GND 0.39322f
C1388 VDD.n1000 GND 0.070647f
C1389 VDD.t110 GND 0.057758f
C1390 VDD.n1001 GND 0.070509f
C1391 VDD.n1002 GND 0.003621f
C1392 VDD.n1003 GND 0.003621f
C1393 VDD.n1004 GND 0.003621f
C1394 VDD.n1005 GND 0.003621f
C1395 VDD.n1006 GND 0.003621f
C1396 VDD.n1007 GND 0.003621f
C1397 VDD.n1008 GND 0.003621f
C1398 VDD.n1009 GND 0.003621f
C1399 VDD.n1010 GND 0.003621f
C1400 VDD.n1011 GND 0.003621f
C1401 VDD.n1012 GND 0.003621f
C1402 VDD.n1013 GND 0.003621f
C1403 VDD.n1014 GND 0.003621f
C1404 VDD.n1015 GND 0.003621f
C1405 VDD.n1016 GND 0.003621f
C1406 VDD.n1017 GND 0.003621f
C1407 VDD.n1018 GND 0.003621f
C1408 VDD.n1019 GND 0.003621f
C1409 VDD.n1020 GND 0.003621f
C1410 VDD.n1021 GND 0.003621f
C1411 VDD.n1022 GND 0.003621f
C1412 VDD.n1023 GND 0.003621f
C1413 VDD.n1024 GND 0.003621f
C1414 VDD.n1025 GND 0.003621f
C1415 VDD.n1026 GND 0.003621f
C1416 VDD.n1027 GND 0.003621f
C1417 VDD.n1028 GND 0.003621f
C1418 VDD.n1029 GND 0.003621f
C1419 VDD.n1030 GND 0.003621f
C1420 VDD.n1031 GND 0.003621f
C1421 VDD.n1032 GND 0.003621f
C1422 VDD.n1033 GND 0.003621f
C1423 VDD.n1034 GND 0.003621f
C1424 VDD.n1035 GND 0.003621f
C1425 VDD.n1036 GND 0.003621f
C1426 VDD.n1037 GND 0.003621f
C1427 VDD.n1038 GND 0.003621f
C1428 VDD.n1039 GND 0.003621f
C1429 VDD.n1040 GND 0.003621f
C1430 VDD.n1041 GND 0.003621f
C1431 VDD.n1042 GND 0.003621f
C1432 VDD.n1043 GND 0.003621f
C1433 VDD.n1044 GND 0.003621f
C1434 VDD.n1045 GND 0.003621f
C1435 VDD.n1046 GND 0.003621f
C1436 VDD.n1047 GND 0.003621f
C1437 VDD.n1048 GND 0.003621f
C1438 VDD.n1049 GND 0.003621f
C1439 VDD.n1050 GND 0.003621f
C1440 VDD.n1051 GND 0.003621f
C1441 VDD.n1052 GND 0.003621f
C1442 VDD.n1053 GND 0.003621f
C1443 VDD.n1054 GND 0.003621f
C1444 VDD.n1055 GND 0.003621f
C1445 VDD.n1056 GND 0.003621f
C1446 VDD.n1057 GND 0.003621f
C1447 VDD.n1058 GND 0.003621f
C1448 VDD.n1059 GND 0.003621f
C1449 VDD.n1060 GND 0.003621f
C1450 VDD.n1061 GND 0.003621f
C1451 VDD.n1062 GND 0.003621f
C1452 VDD.n1063 GND 0.003621f
C1453 VDD.n1064 GND 0.003621f
C1454 VDD.n1065 GND 0.003621f
C1455 VDD.n1066 GND 0.003621f
C1456 VDD.n1067 GND 0.003621f
C1457 VDD.n1068 GND 0.003621f
C1458 VDD.n1069 GND 0.003621f
C1459 VDD.n1070 GND 0.003621f
C1460 VDD.n1071 GND 0.003621f
C1461 VDD.n1072 GND 0.003621f
C1462 VDD.n1073 GND 0.003621f
C1463 VDD.n1074 GND 0.003621f
C1464 VDD.n1075 GND 0.003621f
C1465 VDD.n1076 GND 0.003621f
C1466 VDD.n1077 GND 0.003621f
C1467 VDD.n1078 GND 0.003621f
C1468 VDD.n1079 GND 0.003621f
C1469 VDD.n1080 GND 0.003621f
C1470 VDD.n1081 GND 0.003621f
C1471 VDD.n1082 GND 0.003621f
C1472 VDD.n1083 GND 0.003621f
C1473 VDD.n1084 GND 0.003621f
C1474 VDD.n1085 GND 0.003621f
C1475 VDD.n1086 GND 0.003621f
C1476 VDD.n1087 GND 0.003621f
C1477 VDD.n1088 GND 0.003621f
C1478 VDD.n1089 GND 0.003621f
C1479 VDD.n1090 GND 0.003621f
C1480 VDD.n1091 GND 0.003621f
C1481 VDD.n1092 GND 0.003621f
C1482 VDD.n1093 GND 0.003621f
C1483 VDD.n1094 GND 0.003621f
C1484 VDD.n1095 GND 0.003621f
C1485 VDD.n1096 GND 0.003621f
C1486 VDD.n1097 GND 0.003621f
C1487 VDD.n1098 GND 0.003621f
C1488 VDD.n1099 GND 0.003621f
C1489 VDD.n1100 GND 0.003621f
C1490 VDD.n1101 GND 0.003621f
C1491 VDD.n1102 GND 0.003621f
C1492 VDD.n1103 GND 0.003621f
C1493 VDD.n1104 GND 0.003621f
C1494 VDD.n1105 GND 0.003621f
C1495 VDD.n1106 GND 0.003621f
C1496 VDD.n1107 GND 0.003621f
C1497 VDD.n1108 GND 0.003621f
C1498 VDD.n1109 GND 0.003621f
C1499 VDD.n1110 GND 0.003621f
C1500 VDD.n1111 GND 0.003621f
C1501 VDD.n1112 GND 0.003621f
C1502 VDD.n1113 GND 0.003621f
C1503 VDD.n1114 GND 0.003621f
C1504 VDD.n1115 GND 0.003621f
C1505 VDD.n1116 GND 0.003621f
C1506 VDD.n1117 GND 0.003621f
C1507 VDD.n1118 GND 0.003621f
C1508 VDD.n1119 GND 0.003621f
C1509 VDD.n1120 GND 0.003621f
C1510 VDD.n1121 GND 0.003621f
C1511 VDD.n1122 GND 0.003621f
C1512 VDD.n1123 GND 0.003621f
C1513 VDD.n1124 GND 0.003621f
C1514 VDD.n1125 GND 0.003621f
C1515 VDD.n1126 GND 0.003621f
C1516 VDD.n1127 GND 0.003621f
C1517 VDD.n1128 GND 0.003621f
C1518 VDD.n1129 GND 0.003621f
C1519 VDD.n1130 GND 0.003621f
C1520 VDD.n1131 GND 0.003621f
C1521 VDD.n1132 GND 0.003621f
C1522 VDD.n1133 GND 0.003621f
C1523 VDD.n1134 GND 0.003621f
C1524 VDD.n1135 GND 0.003621f
C1525 VDD.n1136 GND 0.003621f
C1526 VDD.n1137 GND 0.003621f
C1527 VDD.n1138 GND 0.003621f
C1528 VDD.n1139 GND 0.003621f
C1529 VDD.n1140 GND 0.003621f
C1530 VDD.n1141 GND 0.003621f
C1531 VDD.n1142 GND 0.003621f
C1532 VDD.n1143 GND 0.003621f
C1533 VDD.n1144 GND 0.003621f
C1534 VDD.n1145 GND 0.003621f
C1535 VDD.n1146 GND 0.003621f
C1536 VDD.n1147 GND 0.003621f
C1537 VDD.n1148 GND 0.003621f
C1538 VDD.n1149 GND 0.003621f
C1539 VDD.n1150 GND 0.003621f
C1540 VDD.n1151 GND 0.003621f
C1541 VDD.n1152 GND 0.003621f
C1542 VDD.n1153 GND 0.003621f
C1543 VDD.t48 GND 0.087165f
C1544 VDD.t45 GND 0.39322f
C1545 VDD.n1154 GND 0.070647f
C1546 VDD.t47 GND 0.057758f
C1547 VDD.n1155 GND 0.070509f
C1548 VDD.n1156 GND 0.003781f
C1549 VDD.n1159 GND 0.005326f
C1550 VDD.n1160 GND 0.004287f
C1551 VDD.n1161 GND 0.005326f
C1552 VDD.n1162 GND 0.005326f
C1553 VDD.n1163 GND 0.005326f
C1554 VDD.t60 GND 0.159105f
C1555 VDD.t59 GND 0.597454f
C1556 VDD.n1164 GND 0.084294f
C1557 VDD.t61 GND 0.119732f
C1558 VDD.n1165 GND 0.085079f
C1559 VDD.n1166 GND 0.008037f
C1560 VDD.n1167 GND 0.005326f
C1561 VDD.n1168 GND 0.005326f
C1562 VDD.n1169 GND 0.005326f
C1563 VDD.n1170 GND 0.005326f
C1564 VDD.n1171 GND 0.004287f
C1565 VDD.n1172 GND 0.005326f
C1566 VDD.n1173 GND 0.005326f
C1567 VDD.n1174 GND 0.005326f
C1568 VDD.n1175 GND 0.005326f
C1569 VDD.n1176 GND 0.004287f
C1570 VDD.n1177 GND 0.005326f
C1571 VDD.n1178 GND 0.005326f
C1572 VDD.n1179 GND 0.005326f
C1573 VDD.n1180 GND 0.005326f
C1574 VDD.n1181 GND 0.004287f
C1575 VDD.n1182 GND 0.005326f
C1576 VDD.n1183 GND 0.005326f
C1577 VDD.n1184 GND 0.005326f
C1578 VDD.n1185 GND 0.005326f
C1579 VDD.n1186 GND 0.004158f
C1580 VDD.n1187 GND 0.012553f
C1581 VDD.n1188 GND 0.002272f
C1582 VDD.t54 GND 0.159105f
C1583 VDD.t53 GND 0.597454f
C1584 VDD.n1189 GND 0.084294f
C1585 VDD.t55 GND 0.119732f
C1586 VDD.n1190 GND 0.085079f
C1587 VDD.n1191 GND 0.005326f
C1588 VDD.n1193 GND 0.005326f
C1589 VDD.n1196 GND 0.005326f
C1590 VDD.n1199 GND 0.005326f
C1591 VDD.n1202 GND 0.005326f
C1592 VDD.t131 GND 7.73746f
C1593 VDD.t28 GND 8.553611f
C1594 VDD.n1206 GND 4.80687f
C1595 VDD.n1207 GND 0.005326f
C1596 VDD.n1208 GND 0.003558f
C1597 VDD.n1209 GND 0.58089f
C1598 VDD.n1210 GND 0.005326f
C1599 VDD.n1211 GND 0.012553f
C1600 VDD.n1212 GND 0.004287f
C1601 VDD.n1213 GND 0.005326f
C1602 VDD.n1214 GND 0.004287f
C1603 VDD.n1215 GND 0.005326f
C1604 VDD.n1216 GND 0.58089f
C1605 VDD.n1217 GND 0.005326f
C1606 VDD.n1218 GND 0.004287f
C1607 VDD.n1219 GND 0.004287f
C1608 VDD.n1220 GND 0.005326f
C1609 VDD.n1221 GND 0.004287f
C1610 VDD.n1222 GND 0.005326f
C1611 VDD.n1223 GND 0.511183f
C1612 VDD.n1224 GND 0.005326f
C1613 VDD.n1225 GND 0.004287f
C1614 VDD.n1226 GND 0.005326f
C1615 VDD.n1227 GND 0.004287f
C1616 VDD.n1228 GND 0.005326f
C1617 VDD.n1229 GND 0.58089f
C1618 VDD.n1230 GND 0.005326f
C1619 VDD.n1231 GND 0.004287f
C1620 VDD.n1232 GND 0.005326f
C1621 VDD.n1233 GND 0.004287f
C1622 VDD.n1234 GND 0.005326f
C1623 VDD.n1235 GND 0.58089f
C1624 VDD.n1236 GND 0.005326f
C1625 VDD.n1237 GND 0.004287f
C1626 VDD.n1238 GND 0.005326f
C1627 VDD.n1239 GND 0.004287f
C1628 VDD.n1240 GND 0.005326f
C1629 VDD.n1241 GND 0.58089f
C1630 VDD.n1242 GND 0.005326f
C1631 VDD.n1243 GND 0.004287f
C1632 VDD.n1244 GND 0.005326f
C1633 VDD.n1245 GND 0.004287f
C1634 VDD.n1246 GND 0.005326f
C1635 VDD.n1247 GND 0.58089f
C1636 VDD.n1248 GND 0.005326f
C1637 VDD.n1249 GND 0.004287f
C1638 VDD.n1250 GND 0.005326f
C1639 VDD.n1251 GND 0.004287f
C1640 VDD.n1252 GND 0.005326f
C1641 VDD.n1253 GND 0.58089f
C1642 VDD.n1254 GND 0.005326f
C1643 VDD.n1255 GND 0.004287f
C1644 VDD.n1256 GND 0.005326f
C1645 VDD.n1257 GND 0.004287f
C1646 VDD.n1258 GND 0.005326f
C1647 VDD.n1259 GND 0.58089f
C1648 VDD.n1260 GND 0.005326f
C1649 VDD.n1261 GND 0.004287f
C1650 VDD.n1262 GND 0.005326f
C1651 VDD.n1263 GND 0.004287f
C1652 VDD.n1264 GND 0.005326f
C1653 VDD.n1265 GND 0.377579f
C1654 VDD.n1266 GND 0.005326f
C1655 VDD.n1267 GND 0.004287f
C1656 VDD.n1268 GND 0.005326f
C1657 VDD.n1269 GND 0.004287f
C1658 VDD.n1270 GND 0.005326f
C1659 VDD.n1271 GND 0.58089f
C1660 VDD.t2 GND 0.290445f
C1661 VDD.n1272 GND 0.005326f
C1662 VDD.n1273 GND 0.004287f
C1663 VDD.n1274 GND 0.005326f
C1664 VDD.n1275 GND 0.004287f
C1665 VDD.n1276 GND 0.005326f
C1666 VDD.n1277 GND 0.58089f
C1667 VDD.n1278 GND 0.005326f
C1668 VDD.n1279 GND 0.004287f
C1669 VDD.n1280 GND 0.005326f
C1670 VDD.n1281 GND 0.004287f
C1671 VDD.n1282 GND 0.005326f
C1672 VDD.n1283 GND 0.58089f
C1673 VDD.n1284 GND 0.005326f
C1674 VDD.n1285 GND 0.004287f
C1675 VDD.n1286 GND 0.005326f
C1676 VDD.n1287 GND 0.004287f
C1677 VDD.n1288 GND 0.005326f
C1678 VDD.n1289 GND 0.58089f
C1679 VDD.n1290 GND 0.005326f
C1680 VDD.n1291 GND 0.004287f
C1681 VDD.n1292 GND 0.005326f
C1682 VDD.n1293 GND 0.004287f
C1683 VDD.n1294 GND 0.005326f
C1684 VDD.n1295 GND 0.58089f
C1685 VDD.n1296 GND 0.005326f
C1686 VDD.n1297 GND 0.004287f
C1687 VDD.n1298 GND 0.005307f
C1688 VDD.n1299 GND 0.004287f
C1689 VDD.n1300 GND 0.005326f
C1690 VDD.n1301 GND 0.58089f
C1691 VDD.n1302 GND 0.005326f
C1692 VDD.n1303 GND 0.004287f
C1693 VDD.n1304 GND 0.005326f
C1694 VDD.n1305 GND 0.004287f
C1695 VDD.n1306 GND 0.005326f
C1696 VDD.n1307 GND 0.58089f
C1697 VDD.n1308 GND 0.005326f
C1698 VDD.n1309 GND 0.004287f
C1699 VDD.n1310 GND 0.005326f
C1700 VDD.n1311 GND 0.004287f
C1701 VDD.n1312 GND 0.005326f
C1702 VDD.n1313 GND 0.58089f
C1703 VDD.n1314 GND 0.005326f
C1704 VDD.n1315 GND 0.004287f
C1705 VDD.n1316 GND 0.005326f
C1706 VDD.n1317 GND 0.004287f
C1707 VDD.n1318 GND 0.005326f
C1708 VDD.n1319 GND 0.58089f
C1709 VDD.n1320 GND 0.005326f
C1710 VDD.n1321 GND 0.004287f
C1711 VDD.n1322 GND 0.005326f
C1712 VDD.n1323 GND 0.004287f
C1713 VDD.n1324 GND 0.005326f
C1714 VDD.n1325 GND 0.58089f
C1715 VDD.n1326 GND 0.005326f
C1716 VDD.n1327 GND 0.004287f
C1717 VDD.n1328 GND 0.005326f
C1718 VDD.n1329 GND 0.004287f
C1719 VDD.n1330 GND 0.005326f
C1720 VDD.t11 GND 0.290445f
C1721 VDD.n1331 GND 0.005326f
C1722 VDD.n1332 GND 0.004287f
C1723 VDD.n1333 GND 0.005326f
C1724 VDD.n1334 GND 0.004287f
C1725 VDD.n1335 GND 0.005326f
C1726 VDD.n1336 GND 0.58089f
C1727 VDD.n1337 GND 0.005326f
C1728 VDD.n1338 GND 0.004287f
C1729 VDD.n1339 GND 0.005326f
C1730 VDD.n1340 GND 0.004287f
C1731 VDD.n1341 GND 0.005326f
C1732 VDD.n1342 GND 0.58089f
C1733 VDD.n1343 GND 0.005326f
C1734 VDD.n1344 GND 0.004287f
C1735 VDD.n1345 GND 0.005326f
C1736 VDD.n1346 GND 0.004287f
C1737 VDD.n1347 GND 0.005326f
C1738 VDD.n1348 GND 0.58089f
C1739 VDD.n1349 GND 0.005326f
C1740 VDD.n1350 GND 0.004287f
C1741 VDD.n1351 GND 0.005326f
C1742 VDD.n1352 GND 0.004287f
C1743 VDD.n1353 GND 0.005326f
C1744 VDD.n1354 GND 0.58089f
C1745 VDD.n1355 GND 0.005326f
C1746 VDD.n1356 GND 0.004287f
C1747 VDD.n1357 GND 0.005326f
C1748 VDD.n1358 GND 0.004287f
C1749 VDD.n1359 GND 0.005326f
C1750 VDD.n1360 GND 0.58089f
C1751 VDD.n1361 GND 0.005326f
C1752 VDD.n1362 GND 0.004287f
C1753 VDD.n1363 GND 0.005326f
C1754 VDD.n1364 GND 0.004287f
C1755 VDD.n1365 GND 0.005326f
C1756 VDD.n1366 GND 0.58089f
C1757 VDD.n1367 GND 0.005326f
C1758 VDD.n1368 GND 0.004287f
C1759 VDD.n1369 GND 0.005326f
C1760 VDD.n1370 GND 0.004287f
C1761 VDD.n1371 GND 0.005326f
C1762 VDD.t34 GND 0.290445f
C1763 VDD.n1372 GND 0.005326f
C1764 VDD.n1373 GND 0.004287f
C1765 VDD.n1374 GND 0.005326f
C1766 VDD.n1375 GND 0.004287f
C1767 VDD.n1376 GND 0.005326f
C1768 VDD.n1377 GND 0.58089f
C1769 VDD.n1378 GND 0.511183f
C1770 VDD.n1379 GND 0.005326f
C1771 VDD.n1380 GND 0.004287f
C1772 VDD.n1381 GND 0.005326f
C1773 VDD.n1382 GND 0.004287f
C1774 VDD.n1383 GND 0.005326f
C1775 VDD.n1384 GND 0.58089f
C1776 VDD.n1385 GND 0.005326f
C1777 VDD.n1386 GND 0.004287f
C1778 VDD.n1387 GND 0.012553f
C1779 VDD.n1388 GND 0.012553f
C1780 VDD.n1389 GND 1.34186f
C1781 VDD.n1390 GND 0.012553f
C1782 VDD.n1391 GND 0.005326f
C1783 VDD.n1393 GND 0.005326f
C1784 VDD.n1394 GND 0.005326f
C1785 VDD.n1395 GND 0.004287f
C1786 VDD.n1396 GND 0.005326f
C1787 VDD.n1397 GND 0.005326f
C1788 VDD.n1399 GND 0.005326f
C1789 VDD.n1400 GND 0.005326f
C1790 VDD.n1402 GND 0.005326f
C1791 VDD.n1403 GND 0.004287f
C1792 VDD.n1404 GND 0.005326f
C1793 VDD.n1405 GND 0.005326f
C1794 VDD.n1407 GND 0.005326f
C1795 VDD.n1408 GND 0.005326f
C1796 VDD.n1410 GND 0.005326f
C1797 VDD.n1411 GND 0.004287f
C1798 VDD.n1412 GND 0.005326f
C1799 VDD.n1413 GND 0.005326f
C1800 VDD.n1415 GND 0.005326f
C1801 VDD.n1416 GND 0.005326f
C1802 VDD.n1418 GND 0.005326f
C1803 VDD.t74 GND 0.159105f
C1804 VDD.t72 GND 0.597454f
C1805 VDD.n1419 GND 0.084294f
C1806 VDD.t73 GND 0.119732f
C1807 VDD.n1420 GND 0.085079f
C1808 VDD.n1421 GND 0.005894f
C1809 VDD.n1422 GND 0.005326f
C1810 VDD.n1423 GND 0.005326f
C1811 VDD.n1425 GND 0.005326f
C1812 VDD.n1426 GND 0.005326f
C1813 VDD.n1427 GND 0.004287f
C1814 VDD.n1428 GND 0.005326f
C1815 VDD.n1430 GND 0.005326f
C1816 VDD.n1431 GND 0.005326f
C1817 VDD.n1433 GND 0.005326f
C1818 VDD.n1434 GND 0.005326f
C1819 VDD.n1435 GND 0.004287f
C1820 VDD.n1436 GND 0.005326f
C1821 VDD.n1438 GND 0.005326f
C1822 VDD.n1439 GND 0.005326f
C1823 VDD.n1441 GND 0.005326f
C1824 VDD.n1442 GND 0.005326f
C1825 VDD.n1443 GND 0.004287f
C1826 VDD.n1444 GND 0.005326f
C1827 VDD.n1446 GND 0.005326f
C1828 VDD.n1447 GND 0.005326f
C1829 VDD.n1449 GND 0.005326f
C1830 VDD.n1450 GND 0.005326f
C1831 VDD.n1451 GND 0.004287f
C1832 VDD.n1452 GND 0.005326f
C1833 VDD.n1454 GND 0.005326f
C1834 VDD.n1455 GND 0.005326f
C1835 VDD.n1457 GND 0.005326f
C1836 VDD.n1458 GND 0.005326f
C1837 VDD.n1459 GND 0.004287f
C1838 VDD.n1460 GND 0.005326f
C1839 VDD.n1462 GND 0.005326f
C1840 VDD.n1463 GND 0.005326f
C1841 VDD.n1465 GND 0.005326f
C1842 VDD.n1466 GND 0.005326f
C1843 VDD.n1467 GND 0.004287f
C1844 VDD.n1468 GND 0.005326f
C1845 VDD.n1470 GND 0.005326f
C1846 VDD.n1471 GND 0.005326f
C1847 VDD.n1473 GND 0.005326f
C1848 VDD.n1474 GND 0.005326f
C1849 VDD.n1475 GND 0.004287f
C1850 VDD.n1476 GND 0.005326f
C1851 VDD.n1478 GND 0.005326f
C1852 VDD.n1479 GND 0.005326f
C1853 VDD.n1481 GND 0.005326f
C1854 VDD.n1482 GND 0.005326f
C1855 VDD.n1483 GND 0.004287f
C1856 VDD.n1484 GND 0.005326f
C1857 VDD.n1486 GND 0.005326f
C1858 VDD.n1487 GND 0.005326f
C1859 VDD.n1489 GND 0.005326f
C1860 VDD.t36 GND 0.159105f
C1861 VDD.t33 GND 0.597454f
C1862 VDD.n1490 GND 0.084294f
C1863 VDD.t35 GND 0.119732f
C1864 VDD.n1491 GND 0.085079f
C1865 VDD.n1492 GND 0.005326f
C1866 VDD.n1493 GND 0.004287f
C1867 VDD.n1495 GND 0.004287f
C1868 VDD.n1496 GND 0.005326f
C1869 VDD.n1497 GND 0.005326f
C1870 VDD.n1498 GND 0.005326f
C1871 VDD.n1499 GND 0.005326f
C1872 VDD.n1501 GND 0.005326f
C1873 VDD.n1502 GND 0.005326f
C1874 VDD.n1503 GND 0.004287f
C1875 VDD.n1504 GND 0.005326f
C1876 VDD.n1506 GND 0.005326f
C1877 VDD.n1507 GND 0.005326f
C1878 VDD.n1509 GND 0.005326f
C1879 VDD.n1510 GND 0.005326f
C1880 VDD.n1511 GND 0.004287f
C1881 VDD.n1512 GND 0.005326f
C1882 VDD.n1514 GND 0.005326f
C1883 VDD.n1515 GND 0.005326f
C1884 VDD.n1517 GND 0.005326f
C1885 VDD.n1518 GND 0.005326f
C1886 VDD.n1519 GND 0.004222f
C1887 VDD.n1520 GND 0.005326f
C1888 VDD.n1521 GND 0.002936f
C1889 VDD.n1523 GND 0.005326f
C1890 VDD.n1525 GND 0.004287f
C1891 VDD.n1526 GND 0.005326f
C1892 VDD.n1527 GND 0.005326f
C1893 VDD.n1528 GND 0.005326f
C1894 VDD.n1530 GND 0.005326f
C1895 VDD.n1531 GND 0.005326f
C1896 VDD.n1532 GND 0.004287f
C1897 VDD.n1533 GND 0.005326f
C1898 VDD.n1535 GND 0.005326f
C1899 VDD.n1536 GND 0.005326f
C1900 VDD.n1538 GND 0.005326f
C1901 VDD.n1539 GND 0.005326f
C1902 VDD.n1540 GND 0.004287f
C1903 VDD.n1541 GND 0.005326f
C1904 VDD.n1543 GND 0.005326f
C1905 VDD.n1544 GND 0.005326f
C1906 VDD.n1546 GND 0.005326f
C1907 VDD.n1547 GND 0.005326f
C1908 VDD.n1548 GND 0.004287f
C1909 VDD.n1549 GND 0.005326f
C1910 VDD.n1551 GND 0.005326f
C1911 VDD.n1552 GND 0.005326f
C1912 VDD.n1553 GND 0.002272f
C1913 VDD.n1555 GND 0.005326f
C1914 VDD.t90 GND 0.159105f
C1915 VDD.t88 GND 0.597454f
C1916 VDD.n1556 GND 0.084294f
C1917 VDD.t89 GND 0.119732f
C1918 VDD.n1557 GND 0.085079f
C1919 VDD.n1558 GND 0.008037f
C1920 VDD.n1559 GND 0.004158f
C1921 VDD.n1560 GND 0.005326f
C1922 VDD.n1561 GND 0.005326f
C1923 VDD.n1562 GND 0.005326f
C1924 VDD.n1563 GND 0.004287f
C1925 VDD.n1564 GND 0.004287f
C1926 VDD.n1565 GND 0.004287f
C1927 VDD.n1566 GND 0.005326f
C1928 VDD.n1567 GND 0.005326f
C1929 VDD.n1568 GND 0.005326f
C1930 VDD.n1569 GND 0.004287f
C1931 VDD.n1570 GND 0.004287f
C1932 VDD.n1571 GND 0.004287f
C1933 VDD.n1572 GND 0.005326f
C1934 VDD.n1573 GND 0.005326f
C1935 VDD.n1574 GND 0.005326f
C1936 VDD.n1575 GND 0.004287f
C1937 VDD.n1576 GND 0.004287f
C1938 VDD.n1577 GND 0.004287f
C1939 VDD.n1578 GND 0.005326f
C1940 VDD.n1579 GND 0.005326f
C1941 VDD.n1580 GND 0.005326f
C1942 VDD.n1581 GND 0.004287f
C1943 VDD.n1582 GND 0.005326f
C1944 VDD.n1583 GND 0.005326f
C1945 VDD.n1585 GND 0.005326f
C1946 VDD.t99 GND 0.159105f
C1947 VDD.t97 GND 0.597454f
C1948 VDD.n1586 GND 0.084294f
C1949 VDD.t98 GND 0.119732f
C1950 VDD.n1587 GND 0.085079f
C1951 VDD.n1588 GND 0.008037f
C1952 VDD.n1589 GND 0.005326f
C1953 VDD.n1590 GND 0.005326f
C1954 VDD.n1591 GND 0.005326f
C1955 VDD.n1592 GND 0.004287f
C1956 VDD.n1593 GND 0.004287f
C1957 VDD.n1594 GND 0.004287f
C1958 VDD.n1595 GND 0.005326f
C1959 VDD.n1596 GND 0.005326f
C1960 VDD.n1597 GND 0.005326f
C1961 VDD.n1598 GND 0.004287f
C1962 VDD.n1599 GND 0.004287f
C1963 VDD.n1600 GND 0.004287f
C1964 VDD.n1601 GND 0.005326f
C1965 VDD.n1602 GND 0.005326f
C1966 VDD.n1603 GND 0.005326f
C1967 VDD.n1604 GND 0.004287f
C1968 VDD.n1605 GND 0.004287f
C1969 VDD.n1606 GND 0.004287f
C1970 VDD.n1607 GND 0.005326f
C1971 VDD.n1608 GND 0.005326f
C1972 VDD.n1609 GND 0.005326f
C1973 VDD.n1610 GND 0.004287f
C1974 VDD.n1611 GND 0.005326f
C1975 VDD.n1612 GND 0.005326f
C1976 VDD.n1614 GND 0.005326f
C1977 VDD.n1615 GND 0.002872f
C1978 VDD.n1616 GND 0.008037f
C1979 VDD.n1617 GND 0.004287f
C1980 VDD.n1618 GND 0.005326f
C1981 VDD.n1619 GND 0.005326f
C1982 VDD.n1620 GND 0.005326f
C1983 VDD.n1621 GND 0.004287f
C1984 VDD.n1622 GND 0.004287f
C1985 VDD.n1623 GND 0.004287f
C1986 VDD.n1624 GND 0.005326f
C1987 VDD.n1625 GND 0.005326f
C1988 VDD.n1626 GND 0.005326f
C1989 VDD.n1627 GND 0.004287f
C1990 VDD.n1628 GND 0.004287f
C1991 VDD.n1629 GND 0.004287f
C1992 VDD.n1630 GND 0.005326f
C1993 VDD.n1631 GND 0.005326f
C1994 VDD.n1632 GND 0.005326f
C1995 VDD.n1633 GND 0.004287f
C1996 VDD.n1634 GND 0.004287f
C1997 VDD.n1635 GND 0.004287f
C1998 VDD.n1636 GND 0.005326f
C1999 VDD.n1637 GND 0.005326f
C2000 VDD.n1638 GND 0.005326f
C2001 VDD.n1639 GND 0.004287f
C2002 VDD.n1640 GND 0.002808f
C2003 VDD.t58 GND 0.159105f
C2004 VDD.t56 GND 0.597454f
C2005 VDD.n1641 GND 0.084294f
C2006 VDD.t57 GND 0.119732f
C2007 VDD.n1642 GND 0.085079f
C2008 VDD.n1643 GND 0.005894f
C2009 VDD.n1644 GND 0.002208f
C2010 VDD.n1645 GND 0.005326f
C2011 VDD.n1646 GND 0.005326f
C2012 VDD.n1647 GND 0.005326f
C2013 VDD.n1648 GND 0.004287f
C2014 VDD.n1649 GND 0.004287f
C2015 VDD.n1650 GND 0.004287f
C2016 VDD.n1651 GND 0.005326f
C2017 VDD.n1652 GND 0.005326f
C2018 VDD.n1653 GND 0.005326f
C2019 VDD.n1654 GND 0.004287f
C2020 VDD.n1655 GND 0.004287f
C2021 VDD.n1656 GND 0.004287f
C2022 VDD.n1657 GND 0.005326f
C2023 VDD.n1658 GND 0.005326f
C2024 VDD.n1659 GND 0.005326f
C2025 VDD.n1660 GND 0.004287f
C2026 VDD.n1661 GND 0.004287f
C2027 VDD.n1662 GND 0.004287f
C2028 VDD.n1663 GND 0.005326f
C2029 VDD.n1664 GND 0.005326f
C2030 VDD.n1665 GND 0.005326f
C2031 VDD.n1666 GND 0.004287f
C2032 VDD.n1667 GND 0.004287f
C2033 VDD.n1668 GND 0.002743f
C2034 VDD.n1669 GND 0.005326f
C2035 VDD.n1670 GND 0.005326f
C2036 VDD.n1671 GND 0.002272f
C2037 VDD.n1672 GND 0.004287f
C2038 VDD.n1673 GND 0.004287f
C2039 VDD.n1674 GND 0.005326f
C2040 VDD.n1675 GND 0.005326f
C2041 VDD.n1676 GND 0.005326f
C2042 VDD.n1677 GND 0.004287f
C2043 VDD.n1678 GND 0.004287f
C2044 VDD.n1679 GND 0.004287f
C2045 VDD.n1680 GND 0.005326f
C2046 VDD.n1681 GND 0.005326f
C2047 VDD.n1682 GND 0.005326f
C2048 VDD.n1683 GND 0.004287f
C2049 VDD.n1684 GND 0.004287f
C2050 VDD.n1685 GND 0.004287f
C2051 VDD.n1686 GND 0.005326f
C2052 VDD.n1687 GND 0.005326f
C2053 VDD.n1688 GND 0.005326f
C2054 VDD.n1689 GND 0.004287f
C2055 VDD.n1690 GND 0.004287f
C2056 VDD.n1691 GND 0.003558f
C2057 VDD.n1692 GND 0.012553f
C2058 VDD.n1693 GND 0.012264f
C2059 VDD.n1694 GND 0.003558f
C2060 VDD.n1695 GND 0.012264f
C2061 VDD.n1696 GND 0.824864f
C2062 VDD.n1697 GND 0.012264f
C2063 VDD.n1698 GND 0.003558f
C2064 VDD.n1699 GND 0.012264f
C2065 VDD.n1700 GND 0.005326f
C2066 VDD.n1701 GND 0.005326f
C2067 VDD.n1702 GND 0.004287f
C2068 VDD.n1703 GND 0.005326f
C2069 VDD.n1704 GND 0.58089f
C2070 VDD.n1705 GND 0.005326f
C2071 VDD.n1706 GND 0.004287f
C2072 VDD.n1707 GND 0.005326f
C2073 VDD.n1708 GND 0.005326f
C2074 VDD.n1709 GND 0.005326f
C2075 VDD.n1710 GND 0.004287f
C2076 VDD.n1711 GND 0.005326f
C2077 VDD.n1712 GND 0.58089f
C2078 VDD.n1713 GND 0.005326f
C2079 VDD.n1714 GND 0.004287f
C2080 VDD.n1715 GND 0.005326f
C2081 VDD.n1716 GND 0.005326f
C2082 VDD.n1717 GND 0.005326f
C2083 VDD.n1718 GND 0.004287f
C2084 VDD.n1719 GND 0.005326f
C2085 VDD.n1720 GND 0.360152f
C2086 VDD.n1721 GND 0.005326f
C2087 VDD.n1722 GND 0.004287f
C2088 VDD.n1723 GND 0.005326f
C2089 VDD.n1724 GND 0.005326f
C2090 VDD.n1725 GND 0.005326f
C2091 VDD.n1726 GND 0.004287f
C2092 VDD.n1727 GND 0.005326f
C2093 VDD.n1728 GND 0.58089f
C2094 VDD.n1729 GND 0.005326f
C2095 VDD.n1730 GND 0.004287f
C2096 VDD.n1731 GND 0.005326f
C2097 VDD.n1732 GND 0.005326f
C2098 VDD.n1733 GND 0.005326f
C2099 VDD.n1734 GND 0.004287f
C2100 VDD.n1735 GND 0.005326f
C2101 VDD.n1736 GND 0.58089f
C2102 VDD.n1737 GND 0.005326f
C2103 VDD.n1738 GND 0.004287f
C2104 VDD.n1739 GND 0.005326f
C2105 VDD.n1740 GND 0.005326f
C2106 VDD.n1741 GND 0.005326f
C2107 VDD.n1742 GND 0.004287f
C2108 VDD.n1743 GND 0.005326f
C2109 VDD.n1744 GND 0.58089f
C2110 VDD.n1745 GND 0.005326f
C2111 VDD.n1746 GND 0.004287f
C2112 VDD.n1747 GND 0.005326f
C2113 VDD.n1748 GND 0.005326f
C2114 VDD.n1749 GND 0.005326f
C2115 VDD.n1750 GND 0.004287f
C2116 VDD.n1751 GND 0.005326f
C2117 VDD.n1752 GND 0.58089f
C2118 VDD.n1753 GND 0.005326f
C2119 VDD.n1754 GND 0.004287f
C2120 VDD.n1755 GND 0.005326f
C2121 VDD.n1756 GND 0.005326f
C2122 VDD.n1757 GND 0.005326f
C2123 VDD.n1758 GND 0.004287f
C2124 VDD.n1759 GND 0.005326f
C2125 VDD.n1760 GND 0.58089f
C2126 VDD.n1761 GND 0.005326f
C2127 VDD.n1762 GND 0.004287f
C2128 VDD.n1763 GND 0.005326f
C2129 VDD.n1764 GND 0.005326f
C2130 VDD.n1765 GND 0.005326f
C2131 VDD.n1766 GND 0.004287f
C2132 VDD.n1767 GND 0.005326f
C2133 VDD.n1768 GND 0.377579f
C2134 VDD.n1769 GND 0.58089f
C2135 VDD.n1770 GND 0.005326f
C2136 VDD.n1771 GND 0.004287f
C2137 VDD.n1772 GND 0.005326f
C2138 VDD.n1773 GND 0.005326f
C2139 VDD.n1774 GND 0.005326f
C2140 VDD.n1775 GND 0.004287f
C2141 VDD.n1776 GND 0.005326f
C2142 VDD.n1777 GND 0.493757f
C2143 VDD.n1778 GND 0.005326f
C2144 VDD.n1779 GND 0.004287f
C2145 VDD.n1780 GND 0.005326f
C2146 VDD.n1781 GND 0.005326f
C2147 VDD.n1782 GND 0.005326f
C2148 VDD.n1783 GND 0.004287f
C2149 VDD.n1784 GND 0.005326f
C2150 VDD.n1785 GND 0.58089f
C2151 VDD.n1786 GND 0.005326f
C2152 VDD.n1787 GND 0.004287f
C2153 VDD.n1788 GND 0.005326f
C2154 VDD.n1789 GND 0.005326f
C2155 VDD.n1790 GND 0.005326f
C2156 VDD.n1791 GND 0.004287f
C2157 VDD.n1792 GND 0.005326f
C2158 VDD.n1793 GND 0.58089f
C2159 VDD.n1794 GND 0.005326f
C2160 VDD.n1795 GND 0.004287f
C2161 VDD.n1796 GND 0.005326f
C2162 VDD.n1797 GND 0.005326f
C2163 VDD.n1798 GND 0.005326f
C2164 VDD.n1799 GND 0.004287f
C2165 VDD.n1800 GND 0.005326f
C2166 VDD.n1801 GND 0.58089f
C2167 VDD.n1802 GND 0.005326f
C2168 VDD.n1803 GND 0.004287f
C2169 VDD.n1804 GND 0.005326f
C2170 VDD.n1805 GND 0.005326f
C2171 VDD.n1806 GND 0.005326f
C2172 VDD.n1807 GND 0.004287f
C2173 VDD.n1808 GND 0.005326f
C2174 VDD.n1809 GND 0.58089f
C2175 VDD.n1810 GND 0.005326f
C2176 VDD.n1811 GND 0.004287f
C2177 VDD.n1812 GND 0.005326f
C2178 VDD.n1813 GND 0.005326f
C2179 VDD.n1814 GND 0.005326f
C2180 VDD.n1815 GND 0.004287f
C2181 VDD.n1816 GND 0.005326f
C2182 VDD.t0 GND 0.58089f
C2183 VDD.n1817 GND 0.005326f
C2184 VDD.n1818 GND 0.004287f
C2185 VDD.t21 GND 0.134559f
C2186 VDD.t12 GND 0.02169f
C2187 VDD.t167 GND 0.02169f
C2188 VDD.n1819 GND 0.097534f
C2189 VDD.n1820 GND 0.579207f
C2190 VDD.t3 GND 0.134559f
C2191 VDD.t17 GND 0.02169f
C2192 VDD.t26 GND 0.02169f
C2193 VDD.n1821 GND 0.097534f
C2194 VDD.n1822 GND 0.55832f
C2195 VDD.n1823 GND 0.29718f
C2196 VDD.t8 GND 0.134559f
C2197 VDD.t15 GND 0.02169f
C2198 VDD.t1 GND 0.02169f
C2199 VDD.n1824 GND 0.097534f
C2200 VDD.n1825 GND 0.55832f
C2201 VDD.n1826 GND 0.204548f
C2202 VDD.t166 GND 0.134559f
C2203 VDD.t25 GND 0.02169f
C2204 VDD.t161 GND 0.02169f
C2205 VDD.n1827 GND 0.097534f
C2206 VDD.n1828 GND 0.55832f
C2207 VDD.n1829 GND 0.204548f
C2208 VDD.t18 GND 0.134559f
C2209 VDD.t24 GND 0.02169f
C2210 VDD.t165 GND 0.02169f
C2211 VDD.n1830 GND 0.097534f
C2212 VDD.n1831 GND 0.55832f
C2213 VDD.n1832 GND 0.255733f
C2214 VDD.n1833 GND 2.08058f
C2215 VDD.n1834 GND 0.118204f
C2216 VDD.n1835 GND 0.005307f
C2217 VDD.n1836 GND 0.005326f
C2218 VDD.n1837 GND 0.004287f
C2219 VDD.n1838 GND 0.005326f
C2220 VDD.n1839 GND 0.58089f
C2221 VDD.n1840 GND 0.005326f
C2222 VDD.n1841 GND 0.004287f
C2223 VDD.n1842 GND 0.005326f
C2224 VDD.n1843 GND 0.005326f
C2225 VDD.n1844 GND 0.005326f
C2226 VDD.n1845 GND 0.004287f
C2227 VDD.n1846 GND 0.005326f
C2228 VDD.n1847 GND 0.58089f
C2229 VDD.n1848 GND 0.005326f
C2230 VDD.n1849 GND 0.004287f
C2231 VDD.n1850 GND 0.005326f
C2232 VDD.n1851 GND 0.005326f
C2233 VDD.n1852 GND 0.005326f
C2234 VDD.n1853 GND 0.004287f
C2235 VDD.n1854 GND 0.005326f
C2236 VDD.n1855 GND 0.58089f
C2237 VDD.n1856 GND 0.005326f
C2238 VDD.n1857 GND 0.004287f
C2239 VDD.n1858 GND 0.005326f
C2240 VDD.n1859 GND 0.005326f
C2241 VDD.n1860 GND 0.005326f
C2242 VDD.n1861 GND 0.004287f
C2243 VDD.n1862 GND 0.005326f
C2244 VDD.n1863 GND 0.58089f
C2245 VDD.n1864 GND 0.005326f
C2246 VDD.n1865 GND 0.004287f
C2247 VDD.n1866 GND 0.005326f
C2248 VDD.n1867 GND 0.005326f
C2249 VDD.n1868 GND 0.005326f
C2250 VDD.n1869 GND 0.004287f
C2251 VDD.n1870 GND 0.005326f
C2252 VDD.n1871 GND 0.493757f
C2253 VDD.n1872 GND 0.005326f
C2254 VDD.n1873 GND 0.004287f
C2255 VDD.n1874 GND 0.005326f
C2256 VDD.n1875 GND 0.005326f
C2257 VDD.n1876 GND 0.005326f
C2258 VDD.n1877 GND 0.004287f
C2259 VDD.n1878 GND 0.005326f
C2260 VDD.n1879 GND 0.58089f
C2261 VDD.n1880 GND 0.005326f
C2262 VDD.n1881 GND 0.004287f
C2263 VDD.n1882 GND 0.005326f
C2264 VDD.n1883 GND 0.005326f
C2265 VDD.n1884 GND 0.005326f
C2266 VDD.n1885 GND 0.004287f
C2267 VDD.n1886 GND 0.005326f
C2268 VDD.n1887 GND 0.58089f
C2269 VDD.n1888 GND 0.005326f
C2270 VDD.n1889 GND 0.004287f
C2271 VDD.n1890 GND 0.005326f
C2272 VDD.n1891 GND 0.005326f
C2273 VDD.n1892 GND 0.005326f
C2274 VDD.n1893 GND 0.004287f
C2275 VDD.n1894 GND 0.005326f
C2276 VDD.n1895 GND 0.58089f
C2277 VDD.n1896 GND 0.005326f
C2278 VDD.n1897 GND 0.004287f
C2279 VDD.n1898 GND 0.005326f
C2280 VDD.n1899 GND 0.005326f
C2281 VDD.n1900 GND 0.005326f
C2282 VDD.n1901 GND 0.004287f
C2283 VDD.n1902 GND 0.005326f
C2284 VDD.n1903 GND 0.58089f
C2285 VDD.n1904 GND 0.005326f
C2286 VDD.n1905 GND 0.004287f
C2287 VDD.n1906 GND 0.005326f
C2288 VDD.n1907 GND 0.005326f
C2289 VDD.n1908 GND 0.005326f
C2290 VDD.n1909 GND 0.004287f
C2291 VDD.n1910 GND 0.005326f
C2292 VDD.n1911 GND 0.58089f
C2293 VDD.n1912 GND 0.005326f
C2294 VDD.n1913 GND 0.004287f
C2295 VDD.n1914 GND 0.005326f
C2296 VDD.n1915 GND 0.005326f
C2297 VDD.n1916 GND 0.005326f
C2298 VDD.n1917 GND 0.004287f
C2299 VDD.n1918 GND 0.005326f
C2300 VDD.n1919 GND 0.58089f
C2301 VDD.n1920 GND 0.005326f
C2302 VDD.n1921 GND 0.004287f
C2303 VDD.n1922 GND 0.005326f
C2304 VDD.n1923 GND 0.005326f
C2305 VDD.n1924 GND 0.005326f
C2306 VDD.n1925 GND 0.004287f
C2307 VDD.n1926 GND 0.005326f
C2308 VDD.t42 GND 0.290445f
C2309 VDD.n1927 GND 0.360152f
C2310 VDD.n1928 GND 0.005326f
C2311 VDD.n1929 GND 0.004287f
C2312 VDD.n1930 GND 0.005326f
C2313 VDD.n1931 GND 0.005326f
C2314 VDD.n1932 GND 0.005326f
C2315 VDD.n1933 GND 0.004287f
C2316 VDD.n1934 GND 0.005326f
C2317 VDD.n1935 GND 0.58089f
C2318 VDD.n1936 GND 0.005326f
C2319 VDD.n1937 GND 0.004287f
C2320 VDD.n1938 GND 0.005326f
C2321 VDD.n1939 GND 0.005326f
C2322 VDD.n1940 GND 0.012264f
C2323 VDD.n1941 GND 0.005326f
C2324 VDD.n1942 GND 0.005326f
C2325 VDD.n1943 GND 0.004287f
C2326 VDD.n1944 GND 0.005326f
C2327 VDD.n1945 GND 0.58089f
C2328 VDD.n1946 GND 0.005326f
C2329 VDD.n1947 GND 0.004287f
C2330 VDD.n1948 GND 0.005326f
C2331 VDD.n1949 GND 0.005326f
C2332 VDD.n1950 GND 0.005326f
C2333 VDD.n1951 GND 0.004287f
C2334 VDD.n1953 GND 0.005326f
C2335 VDD.n1954 GND 0.005326f
C2336 VDD.n1955 GND 0.005326f
C2337 VDD.n1956 GND 0.005326f
C2338 VDD.n1957 GND 0.005326f
C2339 VDD.n1958 GND 0.004287f
C2340 VDD.n1960 GND 0.005326f
C2341 VDD.n1961 GND 0.005326f
C2342 VDD.n1962 GND 0.005326f
C2343 VDD.n1963 GND 0.005326f
C2344 VDD.n1964 GND 0.005326f
C2345 VDD.n1965 GND 0.004287f
C2346 VDD.n1967 GND 0.005326f
C2347 VDD.n1968 GND 0.005326f
C2348 VDD.n1969 GND 0.005326f
C2349 VDD.n1970 GND 0.005326f
C2350 VDD.n1971 GND 0.005326f
C2351 VDD.n1972 GND 0.002272f
C2352 VDD.n1974 GND 0.005326f
C2353 VDD.t76 GND 0.159105f
C2354 VDD.t75 GND 0.597454f
C2355 VDD.n1975 GND 0.084294f
C2356 VDD.t77 GND 0.119732f
C2357 VDD.n1976 GND 0.085079f
C2358 VDD.n1977 GND 0.005894f
C2359 VDD.n1978 GND 0.005326f
C2360 VDD.n1979 GND 0.005326f
C2361 VDD.n1980 GND 0.005326f
C2362 VDD.n1981 GND 0.005326f
C2363 VDD.n1982 GND 0.004287f
C2364 VDD.n1984 GND 0.005326f
C2365 VDD.n1985 GND 0.005326f
C2366 VDD.n1986 GND 0.005326f
C2367 VDD.n1987 GND 0.005326f
C2368 VDD.n1988 GND 0.004207f
C2369 VDD.n1989 GND 0.004287f
C2370 VDD.n1991 GND 0.005326f
C2371 VDD.n1993 GND 0.004287f
C2372 VDD.n1994 GND 0.005326f
C2373 VDD.n1995 GND 0.004287f
C2374 VDD.n1997 GND 0.005326f
C2375 VDD.n1998 GND 0.004287f
C2376 VDD.n1999 GND 0.005326f
C2377 VDD.n2000 GND 0.005326f
C2378 VDD.n2001 GND 0.005326f
C2379 VDD.n2002 GND 0.005326f
C2380 VDD.n2003 GND 0.005326f
C2381 VDD.t63 GND 0.159105f
C2382 VDD.t62 GND 0.597454f
C2383 VDD.n2004 GND 0.084294f
C2384 VDD.t64 GND 0.119732f
C2385 VDD.n2005 GND 0.085079f
C2386 VDD.n2006 GND 0.005894f
C2387 VDD.n2008 GND 0.002808f
C2388 VDD.n2009 GND 0.005326f
C2389 VDD.n2010 GND 0.005326f
C2390 VDD.n2011 GND 0.005326f
C2391 VDD.n2012 GND 0.005326f
C2392 VDD.n2013 GND 0.005326f
C2393 VDD.n2014 GND 0.004287f
C2394 VDD.n2016 GND 0.005326f
C2395 VDD.n2017 GND 0.005326f
C2396 VDD.n2018 GND 0.005326f
C2397 VDD.n2019 GND 0.005326f
C2398 VDD.n2020 GND 0.005326f
C2399 VDD.n2021 GND 0.004287f
C2400 VDD.n2023 GND 0.005326f
C2401 VDD.n2024 GND 0.005326f
C2402 VDD.n2025 GND 0.005326f
C2403 VDD.n2026 GND 0.005326f
C2404 VDD.n2027 GND 0.005326f
C2405 VDD.n2028 GND 0.004287f
C2406 VDD.n2030 GND 0.005326f
C2407 VDD.n2031 GND 0.005326f
C2408 VDD.n2032 GND 0.005326f
C2409 VDD.n2033 GND 0.005326f
C2410 VDD.n2034 GND 0.005326f
C2411 VDD.t43 GND 0.159105f
C2412 VDD.t41 GND 0.597454f
C2413 VDD.n2035 GND 0.084294f
C2414 VDD.t44 GND 0.119732f
C2415 VDD.n2036 GND 0.085079f
C2416 VDD.n2037 GND 0.008037f
C2417 VDD.n2039 GND 0.005326f
C2418 VDD.n2040 GND 0.004287f
C2419 VDD.n2041 GND 0.005326f
C2420 VDD.n2042 GND 0.005326f
C2421 VDD.n2043 GND 0.004287f
C2422 VDD.n2045 GND 0.005326f
C2423 VDD.n2046 GND 0.005326f
C2424 VDD.n2047 GND 0.005326f
C2425 VDD.n2048 GND 0.005326f
C2426 VDD.n2049 GND 0.005326f
C2427 VDD.n2050 GND 0.004287f
C2428 VDD.n2052 GND 0.005326f
C2429 VDD.n2054 GND 0.005326f
C2430 VDD.n2055 GND 0.004287f
C2431 VDD.n2056 GND 0.004287f
C2432 VDD.n2057 GND 0.005326f
C2433 VDD.n2059 GND 0.005326f
C2434 VDD.n2060 GND 0.004287f
C2435 VDD.n2061 GND 0.004287f
C2436 VDD.n2062 GND 0.005326f
C2437 VDD.n2064 GND 0.005326f
C2438 VDD.n2065 GND 0.005326f
C2439 VDD.n2066 GND 0.004287f
C2440 VDD.n2067 GND 0.004287f
C2441 VDD.n2068 GND 0.004287f
C2442 VDD.n2069 GND 0.005326f
C2443 VDD.n2071 GND 0.005326f
C2444 VDD.n2072 GND 0.005326f
C2445 VDD.n2073 GND 0.004287f
C2446 VDD.n2074 GND 0.005326f
C2447 VDD.n2075 GND 0.005326f
C2448 VDD.n2076 GND 0.005326f
C2449 VDD.n2077 GND 0.002872f
C2450 VDD.n2078 GND 0.005326f
C2451 VDD.n2080 GND 0.005326f
C2452 VDD.n2081 GND 0.005326f
C2453 VDD.n2082 GND 0.004287f
C2454 VDD.n2083 GND 0.004287f
C2455 VDD.n2084 GND 0.004287f
C2456 VDD.n2085 GND 0.005326f
C2457 VDD.n2087 GND 0.005326f
C2458 VDD.n2088 GND 0.005326f
C2459 VDD.n2089 GND 0.004287f
C2460 VDD.n2090 GND 0.004287f
C2461 VDD.n2091 GND 0.004287f
C2462 VDD.n2092 GND 0.005326f
C2463 VDD.n2094 GND 0.005326f
C2464 VDD.n2095 GND 0.005326f
C2465 VDD.n2096 GND 0.004287f
C2466 VDD.n2097 GND 0.004287f
C2467 VDD.n2098 GND 0.004287f
C2468 VDD.n2099 GND 0.005326f
C2469 VDD.n2101 GND 0.005326f
C2470 VDD.n2102 GND 0.005326f
C2471 VDD.n2103 GND 0.004287f
C2472 VDD.n2104 GND 0.004287f
C2473 VDD.n2105 GND 0.004287f
C2474 VDD.n2106 GND 0.005326f
C2475 VDD.n2108 GND 0.005326f
C2476 VDD.n2109 GND 0.005326f
C2477 VDD.n2110 GND 0.002208f
C2478 VDD.n2111 GND 0.004287f
C2479 VDD.n2112 GND 0.004287f
C2480 VDD.n2113 GND 0.005326f
C2481 VDD.n2115 GND 0.005326f
C2482 VDD.n2116 GND 0.005326f
C2483 VDD.n2118 GND 0.005326f
C2484 VDD.n2119 GND 0.004287f
C2485 VDD.n2120 GND 0.003781f
C2486 VDD.n2121 GND 1.11034f
C2487 VDD.n2123 GND 0.004287f
C2488 VDD.n2124 GND 0.004287f
C2489 VDD.n2125 GND 0.005326f
C2490 VDD.n2127 GND 0.005326f
C2491 VDD.n2128 GND 0.005326f
C2492 VDD.n2129 GND 0.004287f
C2493 VDD.n2130 GND 0.004287f
C2494 VDD.n2131 GND 0.004287f
C2495 VDD.n2132 GND 0.005326f
C2496 VDD.n2134 GND 0.005326f
C2497 VDD.n2135 GND 0.005326f
C2498 VDD.n2136 GND 0.004287f
C2499 VDD.n2137 GND 0.004287f
C2500 VDD.n2138 GND 0.002743f
C2501 VDD.n2139 GND 0.005326f
C2502 VDD.n2141 GND 0.005326f
C2503 VDD.n2142 GND 0.005326f
C2504 VDD.n2143 GND 0.004287f
C2505 VDD.n2144 GND 0.004287f
C2506 VDD.n2145 GND 0.004287f
C2507 VDD.n2146 GND 0.005326f
C2508 VDD.n2148 GND 0.005326f
C2509 VDD.n2149 GND 0.005326f
C2510 VDD.n2150 GND 0.004287f
C2511 VDD.n2151 GND 0.004287f
C2512 VDD.n2152 GND 0.004287f
C2513 VDD.n2153 GND 0.005326f
C2514 VDD.n2155 GND 0.005326f
C2515 VDD.n2156 GND 0.005326f
C2516 VDD.n2157 GND 0.004287f
C2517 VDD.n2158 GND 0.004287f
C2518 VDD.n2159 GND 0.004287f
C2519 VDD.n2160 GND 0.005326f
C2520 VDD.n2162 GND 0.005326f
C2521 VDD.n2163 GND 0.005326f
C2522 VDD.n2164 GND 0.004287f
C2523 VDD.n2165 GND 0.003558f
C2524 VDD.n2166 GND 0.012553f
C2525 VDD.n2167 GND 0.012264f
C2526 VDD.n2168 GND 0.003558f
C2527 VDD.n2169 GND 0.012264f
C2528 VDD.n2170 GND 0.824864f
C2529 VDD.n2171 GND 0.012264f
C2530 VDD.n2172 GND 0.012553f
C2531 VDD.n2174 GND 0.005326f
C2532 VDD.n2175 GND 0.008037f
C2533 VDD.n2176 GND 0.005326f
C2534 VDD.n2177 GND 0.005326f
C2535 VDD.n2178 GND 0.005326f
C2536 VDD.n2179 GND 0.004287f
C2537 VDD.n2180 GND 0.004287f
C2538 VDD.n2181 GND 0.004287f
C2539 VDD.n2182 GND 0.005326f
C2540 VDD.n2183 GND 0.005326f
C2541 VDD.n2184 GND 0.005326f
C2542 VDD.n2185 GND 0.004287f
C2543 VDD.n2186 GND 0.004287f
C2544 VDD.n2187 GND 0.004287f
C2545 VDD.n2188 GND 0.005326f
C2546 VDD.n2189 GND 0.005326f
C2547 VDD.n2190 GND 0.005326f
C2548 VDD.n2191 GND 0.004287f
C2549 VDD.n2192 GND 0.004287f
C2550 VDD.n2193 GND 0.004287f
C2551 VDD.n2194 GND 0.005326f
C2552 VDD.n2195 GND 0.005326f
C2553 VDD.n2196 GND 0.005326f
C2554 VDD.n2197 GND 0.004287f
C2555 VDD.n2198 GND 0.004287f
C2556 VDD.n2199 GND 0.002936f
C2557 VDD.n2200 GND 0.005326f
C2558 VDD.n2201 GND 0.005326f
C2559 VDD.n2202 GND 0.005326f
C2560 VDD.n2203 GND 0.004222f
C2561 VDD.n2204 GND 0.004287f
C2562 VDD.n2205 GND 0.004287f
C2563 VDD.n2206 GND 0.004207f
C2564 VDD.n2207 GND 1.11034f
C2565 VDD.n2208 GND 0.080335f
C2566 VDD.n2209 GND 0.009548f
C2567 VDD.n2210 GND 0.003621f
C2568 VDD.n2211 GND 0.003621f
C2569 VDD.n2212 GND 0.003621f
C2570 VDD.n2213 GND 0.003621f
C2571 VDD.n2214 GND 0.003621f
C2572 VDD.n2215 GND 0.003621f
C2573 VDD.n2216 GND 0.003621f
C2574 VDD.n2217 GND 0.003621f
C2575 VDD.n2218 GND 0.003621f
C2576 VDD.n2219 GND 0.003621f
C2577 VDD.n2220 GND 0.003621f
C2578 VDD.n2221 GND 0.003621f
C2579 VDD.n2222 GND 0.003621f
C2580 VDD.n2223 GND 0.003621f
C2581 VDD.n2224 GND 0.002716f
C2582 VDD.n2225 GND 0.003621f
C2583 VDD.n2226 GND 0.003621f
C2584 VDD.n2227 GND 0.002716f
C2585 VDD.n2228 GND 0.003621f
C2586 VDD.n2229 GND 0.003621f
C2587 VDD.n2230 GND 0.003621f
C2588 VDD.n2231 GND 0.003621f
C2589 VDD.n2232 GND 0.003621f
C2590 VDD.n2233 GND 0.003621f
C2591 VDD.n2234 GND 0.003621f
C2592 VDD.n2235 GND 0.003621f
C2593 VDD.n2236 GND 0.006279f
C2594 VDD.n2237 GND 0.003621f
C2595 VDD.n2238 GND 0.003621f
C2596 VDD.n2239 GND 0.003621f
C2597 VDD.n2240 GND 0.003621f
C2598 VDD.n2241 GND 0.003621f
C2599 VDD.n2242 GND 0.009548f
C2600 VDD.n2243 GND 0.009198f
C2601 VDD.n2244 GND 0.009198f
C2602 VDD.n2245 GND 0.003621f
C2603 VDD.n2246 GND 0.003621f
C2604 VDD.n2247 GND 0.003621f
C2605 VDD.n2248 GND 0.003621f
C2606 VDD.n2249 GND 0.003621f
C2607 VDD.n2250 GND 0.003621f
C2608 VDD.n2251 GND 0.003621f
C2609 VDD.n2252 GND 0.003621f
C2610 VDD.n2253 GND 0.003621f
C2611 VDD.n2254 GND 0.003621f
C2612 VDD.n2255 GND 0.003621f
C2613 VDD.n2256 GND 0.003621f
C2614 VDD.n2257 GND 0.003621f
C2615 VDD.n2258 GND 0.003621f
C2616 VDD.n2259 GND 0.003621f
C2617 VDD.n2260 GND 0.003621f
C2618 VDD.n2261 GND 0.003621f
C2619 VDD.n2262 GND 0.003621f
C2620 VDD.n2263 GND 0.003621f
C2621 VDD.n2264 GND 0.003621f
C2622 VDD.n2265 GND 0.003621f
C2623 VDD.n2266 GND 0.003621f
C2624 VDD.n2267 GND 0.003621f
C2625 VDD.n2268 GND 0.003621f
C2626 VDD.n2269 GND 0.003621f
C2627 VDD.n2270 GND 0.003621f
C2628 VDD.n2271 GND 0.003621f
C2629 VDD.n2272 GND 0.003621f
C2630 VDD.n2273 GND 0.003621f
C2631 VDD.n2274 GND 0.003621f
C2632 VDD.n2275 GND 0.003621f
C2633 VDD.n2276 GND 0.003621f
C2634 VDD.n2277 GND 0.003621f
C2635 VDD.n2278 GND 0.003621f
C2636 VDD.n2279 GND 0.003621f
C2637 VDD.n2280 GND 0.003621f
C2638 VDD.n2281 GND 0.003621f
C2639 VDD.n2282 GND 0.003621f
C2640 VDD.n2283 GND 0.003621f
C2641 VDD.n2284 GND 0.003621f
C2642 VDD.n2285 GND 0.003621f
C2643 VDD.n2286 GND 0.003621f
C2644 VDD.n2287 GND 0.003621f
C2645 VDD.n2288 GND 0.003621f
C2646 VDD.n2289 GND 0.003621f
C2647 VDD.n2290 GND 0.003621f
C2648 VDD.n2291 GND 0.003621f
C2649 VDD.n2292 GND 0.003621f
C2650 VDD.n2293 GND 0.003621f
C2651 VDD.n2294 GND 0.003621f
C2652 VDD.n2295 GND 0.003621f
C2653 VDD.n2296 GND 0.003621f
C2654 VDD.n2297 GND 0.003621f
C2655 VDD.n2298 GND 0.003621f
C2656 VDD.n2299 GND 0.003621f
C2657 VDD.n2300 GND 0.003621f
C2658 VDD.n2301 GND 0.003621f
C2659 VDD.n2302 GND 0.003621f
C2660 VDD.n2303 GND 0.003621f
C2661 VDD.n2304 GND 0.003621f
C2662 VDD.n2305 GND 0.003621f
C2663 VDD.n2306 GND 0.003621f
C2664 VDD.n2307 GND 0.003621f
C2665 VDD.n2308 GND 0.003621f
C2666 VDD.n2309 GND 0.003621f
C2667 VDD.n2310 GND 0.003621f
C2668 VDD.n2311 GND 0.003621f
C2669 VDD.n2312 GND 0.003621f
C2670 VDD.n2313 GND 0.003621f
C2671 VDD.n2314 GND 0.003621f
C2672 VDD.n2315 GND 0.003621f
C2673 VDD.n2316 GND 0.003621f
C2674 VDD.n2317 GND 0.003621f
C2675 VDD.n2318 GND 0.003621f
C2676 VDD.n2319 GND 0.003621f
C2677 VDD.n2320 GND 0.003621f
C2678 VDD.n2321 GND 0.003621f
C2679 VDD.n2322 GND 0.003621f
C2680 VDD.n2323 GND 0.003621f
C2681 VDD.n2324 GND 0.003621f
C2682 VDD.n2325 GND 0.003621f
C2683 VDD.n2326 GND 0.003621f
C2684 VDD.n2327 GND 0.003621f
C2685 VDD.n2328 GND 0.003621f
C2686 VDD.n2329 GND 0.003621f
C2687 VDD.n2330 GND 0.003621f
C2688 VDD.n2331 GND 0.003621f
C2689 VDD.n2332 GND 0.003621f
C2690 VDD.n2333 GND 0.003621f
C2691 VDD.n2334 GND 0.003621f
C2692 VDD.n2335 GND 0.003621f
C2693 VDD.n2336 GND 0.003621f
C2694 VDD.n2337 GND 0.003621f
C2695 VDD.n2338 GND 0.003621f
C2696 VDD.n2339 GND 0.003621f
C2697 VDD.n2340 GND 0.003621f
C2698 VDD.n2341 GND 0.003621f
C2699 VDD.n2342 GND 0.003621f
C2700 VDD.n2343 GND 0.003621f
C2701 VDD.n2344 GND 0.003621f
C2702 VDD.n2345 GND 0.003621f
C2703 VDD.n2346 GND 0.003621f
C2704 VDD.n2347 GND 0.003621f
C2705 VDD.n2348 GND 0.003621f
C2706 VDD.n2349 GND 0.003621f
C2707 VDD.n2350 GND 0.003621f
C2708 VDD.n2351 GND 0.003621f
C2709 VDD.n2352 GND 0.003621f
C2710 VDD.n2353 GND 0.003621f
C2711 VDD.n2354 GND 0.003621f
C2712 VDD.n2355 GND 0.003621f
C2713 VDD.n2356 GND 0.003621f
C2714 VDD.n2357 GND 0.003621f
C2715 VDD.n2358 GND 0.003621f
C2716 VDD.n2359 GND 0.003621f
C2717 VDD.n2360 GND 0.003621f
C2718 VDD.n2361 GND 0.003621f
C2719 VDD.n2362 GND 0.003621f
C2720 VDD.n2363 GND 0.003621f
C2721 VDD.n2364 GND 0.003621f
C2722 VDD.n2365 GND 0.003621f
C2723 VDD.n2366 GND 0.003621f
C2724 VDD.n2367 GND 0.003621f
C2725 VDD.n2368 GND 0.003621f
C2726 VDD.n2369 GND 0.003621f
C2727 VDD.n2370 GND 0.003621f
C2728 VDD.n2371 GND 0.003621f
C2729 VDD.n2372 GND 0.003621f
C2730 VDD.n2373 GND 0.003621f
C2731 VDD.n2374 GND 0.003621f
C2732 VDD.n2375 GND 0.003621f
C2733 VDD.n2376 GND 0.003621f
C2734 VDD.n2377 GND 0.003621f
C2735 VDD.n2378 GND 0.003621f
C2736 VDD.n2379 GND 0.003621f
C2737 VDD.n2380 GND 0.003621f
C2738 VDD.n2381 GND 0.003621f
C2739 VDD.n2382 GND 0.003621f
C2740 VDD.n2383 GND 0.003621f
C2741 VDD.n2384 GND 0.003621f
C2742 VDD.n2385 GND 0.003621f
C2743 VDD.n2386 GND 0.003621f
C2744 VDD.n2387 GND 0.003621f
C2745 VDD.n2388 GND 0.003621f
C2746 VDD.n2389 GND 0.003621f
C2747 VDD.n2390 GND 0.003621f
C2748 VDD.n2391 GND 0.003621f
C2749 VDD.n2392 GND 0.003621f
C2750 VDD.n2393 GND 0.003621f
C2751 VDD.n2394 GND 0.003621f
C2752 VDD.n2395 GND 0.003621f
C2753 VDD.n2396 GND 0.003621f
C2754 VDD.n2397 GND 0.003621f
C2755 VDD.n2398 GND 0.003621f
C2756 VDD.n2399 GND 0.003621f
C2757 VDD.n2400 GND 0.003621f
C2758 VDD.n2401 GND 0.003621f
C2759 VDD.n2402 GND 0.003621f
C2760 VDD.n2403 GND 0.003621f
C2761 VDD.n2404 GND 0.003621f
C2762 VDD.n2405 GND 0.003621f
C2763 VDD.n2406 GND 0.003621f
C2764 VDD.n2407 GND 0.003621f
C2765 VDD.n2408 GND 0.003621f
C2766 VDD.n2409 GND 0.003621f
C2767 VDD.n2410 GND 0.003621f
C2768 VDD.n2411 GND 0.003621f
C2769 VDD.n2412 GND 0.003621f
C2770 VDD.n2413 GND 0.003621f
C2771 VDD.n2414 GND 0.003621f
C2772 VDD.n2415 GND 0.194598f
C2773 VDD.n2416 GND 0.003621f
C2774 VDD.n2417 GND 0.003621f
C2775 VDD.n2418 GND 0.003621f
C2776 VDD.n2419 GND 0.003621f
C2777 VDD.n2420 GND 0.003621f
C2778 VDD.n2421 GND 0.003621f
C2779 VDD.n2422 GND 0.003621f
C2780 VDD.n2423 GND 0.003621f
C2781 VDD.n2424 GND 0.003621f
C2782 VDD.n2425 GND 0.003621f
C2783 VDD.n2426 GND 0.003621f
C2784 VDD.n2427 GND 0.003621f
C2785 VDD.n2428 GND 0.003621f
C2786 VDD.n2429 GND 0.003621f
C2787 VDD.n2430 GND 0.003621f
C2788 VDD.n2431 GND 0.009198f
C2789 VDD.n2432 GND 0.009198f
C2790 VDD.n2433 GND 0.009548f
C2791 VDD.n2434 GND 0.003621f
C2792 VDD.n2435 GND 0.003621f
C2793 VDD.n2436 GND 0.003621f
C2794 VDD.n2437 GND 0.003621f
C2795 VDD.n2438 GND 0.003621f
C2796 VDD.n2439 GND 0.006279f
C2797 VDD.n2440 GND 0.003621f
C2798 VDD.n2441 GND 0.003621f
C2799 VDD.n2442 GND 0.003621f
C2800 VDD.n2443 GND 0.003621f
C2801 VDD.n2444 GND 0.003621f
C2802 VDD.n2445 GND 0.003621f
C2803 VDD.n2446 GND 0.003621f
C2804 VDD.n2447 GND 0.003621f
C2805 VDD.n2448 GND 0.002716f
C2806 VDD.n2449 GND 0.003621f
C2807 VDD.n2450 GND 0.003621f
C2808 VDD.n2451 GND 0.002716f
C2809 VDD.n2452 GND 0.003621f
C2810 VDD.n2453 GND 0.003621f
C2811 VDD.n2454 GND 0.003621f
C2812 VDD.n2455 GND 0.003621f
C2813 VDD.n2456 GND 0.003621f
C2814 VDD.n2457 GND 0.003621f
C2815 VDD.n2458 GND 0.003621f
C2816 VDD.n2459 GND 0.003621f
C2817 VDD.n2460 GND 0.003621f
C2818 VDD.n2461 GND 0.003621f
C2819 VDD.n2462 GND 0.003621f
C2820 VDD.n2463 GND 1.66135f
C2821 VDD.n2465 GND 0.009548f
C2822 VDD.n2466 GND 0.009548f
C2823 VDD.n2467 GND 0.009198f
C2824 VDD.n2468 GND 0.003621f
C2825 VDD.n2469 GND 0.003621f
C2826 VDD.n2470 GND 0.395005f
C2827 VDD.n2471 GND 0.003621f
C2828 VDD.n2472 GND 0.003621f
C2829 VDD.n2473 GND 0.003621f
C2830 VDD.n2474 GND 0.003621f
C2831 VDD.n2475 GND 0.003621f
C2832 VDD.n2476 GND 0.395005f
C2833 VDD.n2477 GND 0.003621f
C2834 VDD.n2478 GND 0.003621f
C2835 VDD.n2479 GND 0.003621f
C2836 VDD.n2480 GND 0.003621f
C2837 VDD.n2481 GND 0.003621f
C2838 VDD.n2482 GND 0.395005f
C2839 VDD.n2483 GND 0.003621f
C2840 VDD.n2484 GND 0.003621f
C2841 VDD.n2485 GND 0.003621f
C2842 VDD.n2486 GND 0.003621f
C2843 VDD.n2487 GND 0.003621f
C2844 VDD.n2488 GND 0.395005f
C2845 VDD.n2489 GND 0.003621f
C2846 VDD.n2490 GND 0.003621f
C2847 VDD.n2491 GND 0.003621f
C2848 VDD.n2492 GND 0.003621f
C2849 VDD.n2493 GND 0.003621f
C2850 VDD.n2494 GND 0.214929f
C2851 VDD.n2495 GND 0.003621f
C2852 VDD.n2496 GND 0.003621f
C2853 VDD.n2497 GND 0.003621f
C2854 VDD.n2498 GND 0.003621f
C2855 VDD.n2499 GND 0.003621f
C2856 VDD.n2500 GND 0.380483f
C2857 VDD.n2501 GND 0.003621f
C2858 VDD.n2502 GND 0.003621f
C2859 VDD.n2503 GND 0.003621f
C2860 VDD.n2504 GND 0.003621f
C2861 VDD.n2505 GND 0.003621f
C2862 VDD.n2506 GND 0.395005f
C2863 VDD.n2507 GND 0.003621f
C2864 VDD.n2508 GND 0.003621f
C2865 VDD.n2509 GND 0.003621f
C2866 VDD.n2510 GND 0.003621f
C2867 VDD.n2511 GND 0.003621f
C2868 VDD.n2512 GND 0.395005f
C2869 VDD.n2513 GND 0.003621f
C2870 VDD.n2514 GND 0.003621f
C2871 VDD.n2515 GND 0.003621f
C2872 VDD.n2516 GND 0.003621f
C2873 VDD.n2517 GND 0.003621f
C2874 VDD.n2518 GND 0.395005f
C2875 VDD.n2519 GND 0.003621f
C2876 VDD.n2520 GND 0.003621f
C2877 VDD.n2521 GND 0.003621f
C2878 VDD.n2522 GND 0.003621f
C2879 VDD.n2523 GND 0.003621f
C2880 VDD.n2524 GND 0.395005f
C2881 VDD.n2525 GND 0.003621f
C2882 VDD.n2526 GND 0.003621f
C2883 VDD.n2527 GND 0.003621f
C2884 VDD.n2528 GND 0.003621f
C2885 VDD.n2529 GND 0.003621f
C2886 VDD.n2530 GND 0.395005f
C2887 VDD.n2531 GND 0.003621f
C2888 VDD.n2532 GND 0.003621f
C2889 VDD.n2533 GND 0.003621f
C2890 VDD.n2534 GND 0.003621f
C2891 VDD.n2535 GND 0.003621f
C2892 VDD.n2536 GND 0.395005f
C2893 VDD.n2537 GND 0.003621f
C2894 VDD.n2538 GND 0.003621f
C2895 VDD.n2539 GND 0.003621f
C2896 VDD.n2540 GND 0.003621f
C2897 VDD.n2541 GND 0.003621f
C2898 VDD.n2542 GND 0.395005f
C2899 VDD.n2543 GND 0.003621f
C2900 VDD.n2544 GND 0.003621f
C2901 VDD.n2545 GND 0.003621f
C2902 VDD.n2546 GND 0.003621f
C2903 VDD.n2547 GND 0.003621f
C2904 VDD.n2548 GND 0.278827f
C2905 VDD.n2549 GND 0.003621f
C2906 VDD.n2550 GND 0.003621f
C2907 VDD.n2551 GND 0.003621f
C2908 VDD.n2552 GND 0.003621f
C2909 VDD.n2553 GND 0.003621f
C2910 VDD.n2554 GND 0.395005f
C2911 VDD.n2555 GND 0.003621f
C2912 VDD.n2556 GND 0.003621f
C2913 VDD.n2557 GND 0.003621f
C2914 VDD.n2558 GND 0.003621f
C2915 VDD.n2559 GND 0.003621f
C2916 VDD.n2560 GND 0.34563f
C2917 VDD.n2561 GND 0.003621f
C2918 VDD.n2562 GND 0.003621f
C2919 VDD.n2563 GND 0.003621f
C2920 VDD.n2564 GND 0.003621f
C2921 VDD.n2565 GND 0.003621f
C2922 VDD.n2566 GND 0.395005f
C2923 VDD.n2567 GND 0.003621f
C2924 VDD.n2568 GND 0.003621f
C2925 VDD.n2569 GND 0.003621f
C2926 VDD.n2570 GND 0.003621f
C2927 VDD.n2571 GND 0.003621f
C2928 VDD.n2572 GND 0.395005f
C2929 VDD.n2573 GND 0.003621f
C2930 VDD.n2574 GND 0.003621f
C2931 VDD.n2575 GND 0.003621f
C2932 VDD.n2576 GND 0.003621f
C2933 VDD.n2577 GND 0.003621f
C2934 VDD.n2578 GND 0.395005f
C2935 VDD.n2579 GND 0.003621f
C2936 VDD.n2580 GND 0.003621f
C2937 VDD.n2581 GND 0.003621f
C2938 VDD.n2582 GND 0.003621f
C2939 VDD.n2583 GND 0.003621f
C2940 VDD.n2584 GND 0.395005f
C2941 VDD.n2585 GND 0.003621f
C2942 VDD.n2586 GND 0.003621f
C2943 VDD.n2587 GND 0.003621f
C2944 VDD.n2588 GND 0.003621f
C2945 VDD.n2589 GND 0.003621f
C2946 VDD.n2590 GND 0.395005f
C2947 VDD.n2591 GND 0.003621f
C2948 VDD.n2592 GND 0.003621f
C2949 VDD.n2593 GND 0.003621f
C2950 VDD.n2594 GND 0.003621f
C2951 VDD.n2595 GND 0.003621f
C2952 VDD.n2596 GND 0.395005f
C2953 VDD.n2597 GND 0.003621f
C2954 VDD.n2598 GND 0.003621f
C2955 VDD.n2599 GND 0.003621f
C2956 VDD.n2600 GND 0.003621f
C2957 VDD.n2601 GND 0.003621f
C2958 VDD.n2602 GND 0.395005f
C2959 VDD.n2603 GND 0.003621f
C2960 VDD.n2604 GND 0.003621f
C2961 VDD.n2605 GND 0.003621f
C2962 VDD.n2606 GND 0.003621f
C2963 VDD.n2607 GND 0.003621f
C2964 VDD.n2608 GND 0.395005f
C2965 VDD.n2609 GND 0.003621f
C2966 VDD.n2610 GND 0.003621f
C2967 VDD.n2611 GND 0.003621f
C2968 VDD.n2612 GND 0.003621f
C2969 VDD.n2613 GND 0.003621f
C2970 VDD.n2614 GND 0.246878f
C2971 VDD.n2615 GND 0.003621f
C2972 VDD.n2616 GND 0.003621f
C2973 VDD.n2617 GND 0.003621f
C2974 VDD.n2618 GND 0.003621f
C2975 VDD.n2619 GND 0.003621f
C2976 VDD.n2620 GND 0.395005f
C2977 VDD.n2621 GND 0.003621f
C2978 VDD.n2622 GND 0.003621f
C2979 VDD.n2623 GND 0.003621f
C2980 VDD.n2624 GND 0.003621f
C2981 VDD.n2625 GND 0.003621f
C2982 VDD.n2626 GND 0.29335f
C2983 VDD.n2627 GND 0.003621f
C2984 VDD.n2628 GND 0.003621f
C2985 VDD.n2629 GND 0.003621f
C2986 VDD.n2630 GND 0.003621f
C2987 VDD.n2631 GND 0.003621f
C2988 VDD.n2632 GND 0.395005f
C2989 VDD.n2633 GND 0.003621f
C2990 VDD.n2634 GND 0.003621f
C2991 VDD.n2635 GND 0.003621f
C2992 VDD.n2636 GND 0.003621f
C2993 VDD.n2637 GND 0.003621f
C2994 VDD.n2638 GND 0.395005f
C2995 VDD.n2639 GND 0.003621f
C2996 VDD.n2640 GND 0.003621f
C2997 VDD.n2641 GND 0.003621f
C2998 VDD.n2642 GND 0.003621f
C2999 VDD.n2643 GND 0.003621f
C3000 VDD.n2644 GND 0.395005f
C3001 VDD.n2645 GND 0.003621f
C3002 VDD.n2646 GND 0.003621f
C3003 VDD.n2647 GND 0.003621f
C3004 VDD.n2648 GND 0.003621f
C3005 VDD.n2649 GND 0.003621f
C3006 VDD.n2650 GND 0.395005f
C3007 VDD.n2651 GND 0.003621f
C3008 VDD.n2652 GND 0.003621f
C3009 VDD.n2653 GND 0.003621f
C3010 VDD.n2654 GND 0.003621f
C3011 VDD.n2655 GND 0.003621f
C3012 VDD.n2656 GND 0.395005f
C3013 VDD.n2657 GND 0.003621f
C3014 VDD.n2658 GND 0.003621f
C3015 VDD.n2659 GND 0.003621f
C3016 VDD.n2660 GND 0.003621f
C3017 VDD.n2661 GND 0.003621f
C3018 VDD.n2662 GND 0.395005f
C3019 VDD.n2663 GND 0.003621f
C3020 VDD.n2664 GND 0.003621f
C3021 VDD.n2665 GND 0.003621f
C3022 VDD.n2666 GND 0.003621f
C3023 VDD.n2667 GND 0.003621f
C3024 VDD.n2668 GND 0.246878f
C3025 VDD.n2669 GND 0.003621f
C3026 VDD.n2670 GND 0.003621f
C3027 VDD.n2671 GND 0.003621f
C3028 VDD.n2672 GND 0.003621f
C3029 VDD.n2673 GND 0.003621f
C3030 VDD.n2674 GND 0.395005f
C3031 VDD.n2675 GND 0.003621f
C3032 VDD.n2676 GND 0.003621f
C3033 VDD.n2677 GND 0.003621f
C3034 VDD.n2678 GND 0.003621f
C3035 VDD.n2679 GND 0.003621f
C3036 VDD.n2680 GND 0.392101f
C3037 VDD.n2681 GND 0.003621f
C3038 VDD.n2682 GND 0.003621f
C3039 VDD.n2683 GND 0.003621f
C3040 VDD.n2684 GND 0.003621f
C3041 VDD.n2685 GND 0.003621f
C3042 VDD.n2686 GND 0.395005f
C3043 VDD.n2687 GND 0.003621f
C3044 VDD.n2688 GND 0.003621f
C3045 VDD.n2689 GND 0.003621f
C3046 VDD.n2690 GND 0.003621f
C3047 VDD.n2691 GND 0.003621f
C3048 VDD.n2692 GND 0.395005f
C3049 VDD.n2693 GND 0.003621f
C3050 VDD.n2694 GND 0.003621f
C3051 VDD.n2695 GND 0.003621f
C3052 VDD.n2696 GND 0.003621f
C3053 VDD.n2697 GND 0.003621f
C3054 VDD.n2698 GND 0.395005f
C3055 VDD.n2699 GND 0.003621f
C3056 VDD.n2700 GND 0.003621f
C3057 VDD.n2701 GND 0.003621f
C3058 VDD.n2702 GND 0.003621f
C3059 VDD.n2703 GND 0.003621f
C3060 VDD.n2704 GND 0.395005f
C3061 VDD.n2705 GND 0.003621f
C3062 VDD.n2706 GND 0.003621f
C3063 VDD.n2707 GND 0.003621f
C3064 VDD.n2708 GND 0.003621f
C3065 VDD.n2709 GND 0.003621f
C3066 VDD.n2710 GND 0.395005f
C3067 VDD.n2711 GND 0.003621f
C3068 VDD.n2712 GND 0.003621f
C3069 VDD.n2713 GND 0.003621f
C3070 VDD.n2714 GND 0.003621f
C3071 VDD.n2715 GND 0.003621f
C3072 VDD.n2716 GND 0.395005f
C3073 VDD.n2717 GND 0.003621f
C3074 VDD.n2718 GND 0.003621f
C3075 VDD.n2719 GND 0.003621f
C3076 VDD.n2720 GND 0.003621f
C3077 VDD.n2721 GND 0.003621f
C3078 VDD.n2722 GND 0.34563f
C3079 VDD.n2723 GND 0.003621f
C3080 VDD.n2724 GND 0.003621f
C3081 VDD.n2725 GND 0.003621f
C3082 VDD.n2726 GND 0.003621f
C3083 VDD.n2727 GND 0.003621f
C3084 VDD.n2728 GND 0.299158f
C3085 VDD.n2729 GND 0.003621f
C3086 VDD.n2730 GND 0.003621f
C3087 VDD.n2731 GND 0.003621f
C3088 VDD.n2732 GND 0.003621f
C3089 VDD.n2733 GND 0.003621f
C3090 VDD.n2734 GND 0.395005f
C3091 VDD.n2735 GND 0.003621f
C3092 VDD.n2736 GND 0.003621f
C3093 VDD.n2737 GND 0.003621f
C3094 VDD.n2738 GND 0.003621f
C3095 VDD.n2739 GND 0.003621f
C3096 VDD.n2740 GND 0.395005f
C3097 VDD.n2741 GND 0.003621f
C3098 VDD.n2742 GND 0.003621f
C3099 VDD.n2743 GND 0.003621f
C3100 VDD.n2744 GND 0.003621f
C3101 VDD.n2745 GND 0.003621f
C3102 VDD.n2746 GND 0.395005f
C3103 VDD.n2747 GND 0.003621f
C3104 VDD.n2748 GND 0.003621f
C3105 VDD.n2749 GND 0.003621f
C3106 VDD.n2750 GND 0.003621f
C3107 VDD.n2751 GND 0.003621f
C3108 VDD.n2752 GND 0.395005f
C3109 VDD.n2753 GND 0.003621f
C3110 VDD.n2754 GND 0.003621f
C3111 VDD.n2755 GND 0.003621f
C3112 VDD.n2756 GND 0.003621f
C3113 VDD.n2757 GND 0.003621f
C3114 VDD.n2758 GND 0.395005f
C3115 VDD.n2759 GND 0.003621f
C3116 VDD.n2760 GND 0.003621f
C3117 VDD.n2761 GND 0.003621f
C3118 VDD.n2762 GND 0.003621f
C3119 VDD.n2763 GND 0.003621f
C3120 VDD.n2764 GND 0.395005f
C3121 VDD.n2765 GND 0.003621f
C3122 VDD.n2766 GND 0.003621f
C3123 VDD.n2767 GND 0.003621f
C3124 VDD.n2768 GND 0.003621f
C3125 VDD.n2769 GND 0.003621f
C3126 VDD.n2770 GND 0.395005f
C3127 VDD.n2771 GND 0.003621f
C3128 VDD.n2772 GND 0.003621f
C3129 VDD.n2773 GND 0.003621f
C3130 VDD.n2774 GND 0.003621f
C3131 VDD.n2775 GND 0.003621f
C3132 VDD.n2776 GND 0.395005f
C3133 VDD.n2777 GND 0.003621f
C3134 VDD.n2778 GND 0.003621f
C3135 VDD.n2779 GND 0.003621f
C3136 VDD.n2780 GND 0.003621f
C3137 VDD.n2781 GND 0.003621f
C3138 VDD.n2782 GND 0.200407f
C3139 VDD.n2783 GND 0.003621f
C3140 VDD.n2784 GND 0.003621f
C3141 VDD.n2785 GND 0.003621f
C3142 VDD.n2786 GND 0.003621f
C3143 VDD.n2787 GND 0.003621f
C3144 VDD.n2788 GND 0.395005f
C3145 VDD.n2789 GND 0.003621f
C3146 VDD.n2790 GND 0.003621f
C3147 VDD.n2791 GND 0.003621f
C3148 VDD.n2792 GND 0.003621f
C3149 VDD.n2793 GND 0.003621f
C3150 VDD.n2794 GND 0.395005f
C3151 VDD.n2795 GND 0.003621f
C3152 VDD.n2796 GND 0.003621f
C3153 VDD.n2797 GND 0.003621f
C3154 VDD.n2798 GND 0.003621f
C3155 VDD.n2799 GND 0.003621f
C3156 VDD.n2800 GND 0.003621f
C3157 VDD.n2801 GND 0.003621f
C3158 VDD.n2802 GND 0.003621f
C3159 VDD.n2803 GND 0.003621f
C3160 VDD.n2804 GND 0.003621f
C3161 VDD.n2805 GND 0.395005f
C3162 VDD.n2806 GND 0.003621f
C3163 VDD.n2807 GND 0.003621f
C3164 VDD.n2808 GND 0.003621f
C3165 VDD.n2809 GND 0.003621f
C3166 VDD.n2810 GND 0.003621f
C3167 VDD.n2811 GND 0.395005f
C3168 VDD.n2812 GND 0.003621f
C3169 VDD.n2813 GND 0.003621f
C3170 VDD.n2814 GND 0.003621f
C3171 VDD.n2815 GND 0.003621f
C3172 VDD.n2816 GND 0.009566f
C3173 VDD.n2817 GND 0.009198f
C3174 VDD.n2818 GND 0.009548f
C3175 VDD.n2819 GND 0.00918f
C3176 VDD.n2820 GND 0.003621f
C3177 VDD.n2821 GND 0.003621f
C3178 VDD.n2822 GND 0.003621f
C3179 VDD.n2823 GND 0.003621f
C3180 VDD.n2824 GND 0.006279f
C3181 VDD.n2825 GND 0.003621f
C3182 VDD.n2826 GND 0.003621f
C3183 VDD.n2827 GND 0.003621f
C3184 VDD.n2828 GND 0.003621f
C3185 VDD.n2829 GND 0.003621f
C3186 VDD.n2830 GND 0.003621f
C3187 VDD.n2831 GND 0.003621f
C3188 VDD.n2832 GND 0.003621f
C3189 VDD.n2833 GND 0.003621f
C3190 VDD.n2834 GND 0.003621f
C3191 VDD.n2835 GND 0.003621f
C3192 VDD.n2836 GND 0.003621f
C3193 VDD.n2837 GND 0.003621f
C3194 VDD.n2838 GND 0.003621f
C3195 VDD.n2839 GND 0.003621f
C3196 VDD.n2840 GND 0.003621f
C3197 VDD.n2841 GND 0.003621f
C3198 VDD.n2842 GND 0.003621f
C3199 VDD.n2843 GND 0.003621f
C3200 VDD.n2844 GND 0.003621f
C3201 VDD.n2845 GND 0.003621f
C3202 VDD.n2846 GND 0.003621f
C3203 VDD.n2847 GND 0.003621f
C3204 VDD.n2848 GND 0.003621f
C3205 VDD.n2849 GND 0.003621f
C3206 VDD.n2850 GND 0.003621f
C3207 VDD.n2851 GND 0.003621f
C3208 VDD.n2852 GND 0.009548f
C3209 VDD.n2853 GND 0.009548f
C3210 VDD.n2854 GND 0.009198f
C3211 VDD.n2855 GND 0.003621f
C3212 VDD.n2856 GND 0.003621f
C3213 VDD.n2857 GND 0.395005f
C3214 VDD.n2858 GND 0.003621f
C3215 VDD.n2859 GND 0.009198f
C3216 VDD.n2860 GND 0.009566f
C3217 VDD.n2861 GND 0.00918f
C3218 VDD.n2862 GND 0.003621f
C3219 VDD.n2863 GND 0.003621f
C3220 VDD.n2864 GND 0.003621f
C3221 VDD.n2865 GND 0.003621f
C3222 VDD.n2866 GND 0.003621f
C3223 VDD.n2867 GND 0.006279f
C3224 VDD.n2868 GND 0.003621f
C3225 VDD.n2869 GND 0.003621f
C3226 VDD.n2870 GND 0.003621f
C3227 VDD.n2871 GND 0.003621f
C3228 VDD.n2872 GND 0.003621f
C3229 VDD.n2873 GND 0.003621f
C3230 VDD.n2874 GND 0.003621f
C3231 VDD.n2875 GND 0.003621f
C3232 VDD.n2876 GND 0.003621f
C3233 VDD.n2877 GND 0.003621f
C3234 VDD.n2878 GND 0.003621f
C3235 VDD.n2879 GND 0.003621f
C3236 VDD.n2880 GND 0.003621f
C3237 VDD.n2881 GND 0.003621f
C3238 VDD.n2882 GND 0.003621f
C3239 VDD.n2883 GND 0.003621f
C3240 VDD.n2884 GND 0.003621f
C3241 VDD.n2885 GND 0.003621f
C3242 VDD.n2886 GND 0.003621f
C3243 VDD.n2887 GND 0.003621f
C3244 VDD.n2888 GND 0.003621f
C3245 VDD.n2889 GND 0.003621f
C3246 VDD.n2890 GND 0.003621f
C3247 VDD.n2891 GND 0.003621f
C3248 VDD.n2892 GND 0.003621f
C3249 VDD.n2893 GND 0.009548f
C3250 VDD.n2894 GND 0.009548f
C3251 VDD.n2895 GND 2.51816f
C3252 VDD.n2896 GND 2.51816f
C3253 VDD.n2897 GND 0.009548f
C3254 VDD.n2898 GND 0.003621f
C3255 VDD.n2899 GND 0.003621f
C3256 VDD.t71 GND 0.087165f
C3257 VDD.t68 GND 0.39322f
C3258 VDD.n2900 GND 0.070647f
C3259 VDD.t70 GND 0.057758f
C3260 VDD.n2901 GND 0.070509f
C3261 VDD.n2902 GND 0.006279f
C3262 VDD.n2903 GND 0.003621f
C3263 VDD.n2904 GND 0.003621f
C3264 VDD.n2905 GND 0.003621f
C3265 VDD.n2906 GND 0.003621f
C3266 VDD.n2907 GND 0.003621f
C3267 VDD.n2908 GND 0.003621f
C3268 VDD.n2909 GND 0.003621f
C3269 VDD.n2911 GND 0.003621f
C3270 VDD.n2912 GND 0.003621f
C3271 VDD.n2914 GND 0.003621f
C3272 VDD.n2915 GND 0.003621f
C3273 VDD.n2916 GND 0.003621f
C3274 VDD.n2917 GND 0.003621f
C3275 VDD.n2918 GND 0.003621f
C3276 VDD.n2920 GND 0.003621f
C3277 VDD.n2922 GND 0.003621f
C3278 VDD.n2923 GND 0.003621f
C3279 VDD.n2924 GND 0.003621f
C3280 VDD.n2925 GND 0.003621f
C3281 VDD.n2926 GND 0.003621f
C3282 VDD.n2928 GND 0.003621f
C3283 VDD.n2930 GND 0.003621f
C3284 VDD.n2931 GND 0.003621f
C3285 VDD.n2932 GND 0.003621f
C3286 VDD.n2933 GND 0.003621f
C3287 VDD.n2934 GND 0.003621f
C3288 VDD.n2936 GND 0.003621f
C3289 VDD.n2937 GND 0.003621f
C3290 VDD.n2939 GND 0.003621f
C3291 VDD.n2940 GND 0.003621f
C3292 VDD.n2941 GND 0.009548f
C3293 VDD.n2942 GND 0.003621f
C3294 VDD.n2943 GND 0.003621f
C3295 VDD.n2944 GND 0.003621f
C3296 VDD.n2945 GND 0.003621f
C3297 VDD.n2946 GND 0.003621f
C3298 VDD.n2947 GND 0.003621f
C3299 VDD.n2948 GND 0.003621f
C3300 VDD.n2949 GND 0.003621f
C3301 VDD.n2950 GND 0.003621f
C3302 VDD.n2951 GND 0.003621f
C3303 VDD.n2952 GND 0.003621f
C3304 VDD.n2953 GND 0.003621f
C3305 VDD.n2954 GND 0.003621f
C3306 VDD.n2955 GND 0.003621f
C3307 VDD.n2956 GND 0.003621f
C3308 VDD.n2957 GND 0.003621f
C3309 VDD.n2958 GND 0.003621f
C3310 VDD.n2959 GND 0.003621f
C3311 VDD.n2960 GND 0.003621f
C3312 VDD.n2961 GND 0.003621f
C3313 VDD.n2962 GND 0.003621f
C3314 VDD.n2963 GND 0.003621f
C3315 VDD.n2964 GND 0.003621f
C3316 VDD.n2965 GND 0.003621f
C3317 VDD.n2966 GND 0.003621f
C3318 VDD.n2967 GND 0.003621f
C3319 VDD.n2968 GND 0.003621f
C3320 VDD.n2969 GND 0.003621f
C3321 VDD.n2970 GND 0.003621f
C3322 VDD.n2971 GND 0.003621f
C3323 VDD.n2972 GND 0.003621f
C3324 VDD.n2973 GND 0.003621f
C3325 VDD.n2974 GND 0.003621f
C3326 VDD.n2975 GND 0.003621f
C3327 VDD.n2976 GND 0.003621f
C3328 VDD.n2977 GND 0.003621f
C3329 VDD.n2978 GND 0.003621f
C3330 VDD.n2979 GND 0.003621f
C3331 VDD.n2980 GND 0.003621f
C3332 VDD.n2981 GND 0.003621f
C3333 VDD.n2982 GND 0.003621f
C3334 VDD.n2983 GND 0.003621f
C3335 VDD.n2984 GND 0.003621f
C3336 VDD.n2985 GND 0.003621f
C3337 VDD.n2986 GND 0.003621f
C3338 VDD.n2987 GND 0.003621f
C3339 VDD.n2988 GND 0.003621f
C3340 VDD.n2989 GND 0.003621f
C3341 VDD.n2990 GND 0.003621f
C3342 VDD.n2991 GND 0.003621f
C3343 VDD.n2992 GND 0.003621f
C3344 VDD.n2993 GND 0.003621f
C3345 VDD.n2994 GND 0.003621f
C3346 VDD.n2995 GND 0.003621f
C3347 VDD.n2996 GND 0.003621f
C3348 VDD.n2997 GND 0.003621f
C3349 VDD.n2998 GND 0.003621f
C3350 VDD.n2999 GND 0.003621f
C3351 VDD.n3000 GND 0.003621f
C3352 VDD.n3001 GND 0.003621f
C3353 VDD.n3002 GND 0.003621f
C3354 VDD.n3003 GND 0.003621f
C3355 VDD.n3004 GND 0.003621f
C3356 VDD.n3005 GND 0.003621f
C3357 VDD.n3006 GND 0.003621f
C3358 VDD.n3007 GND 0.003621f
C3359 VDD.n3008 GND 0.003621f
C3360 VDD.n3009 GND 0.003621f
C3361 VDD.n3010 GND 0.003621f
C3362 VDD.n3011 GND 0.003621f
C3363 VDD.n3012 GND 0.003621f
C3364 VDD.n3013 GND 0.003621f
C3365 VDD.n3014 GND 0.003621f
C3366 VDD.n3015 GND 0.003621f
C3367 VDD.n3016 GND 0.003621f
C3368 VDD.n3017 GND 0.003621f
C3369 VDD.n3018 GND 0.003621f
C3370 VDD.n3019 GND 0.003621f
C3371 VDD.n3020 GND 0.003621f
C3372 VDD.n3021 GND 0.003621f
C3373 VDD.n3022 GND 0.003621f
C3374 VDD.n3023 GND 0.003621f
C3375 VDD.n3024 GND 0.003621f
C3376 VDD.n3025 GND 0.003621f
C3377 VDD.n3026 GND 0.003621f
C3378 VDD.n3027 GND 0.003621f
C3379 VDD.n3028 GND 0.003621f
C3380 VDD.n3029 GND 0.003621f
C3381 VDD.n3030 GND 0.003621f
C3382 VDD.n3031 GND 0.003621f
C3383 VDD.n3032 GND 0.003621f
C3384 VDD.n3033 GND 0.003621f
C3385 VDD.n3034 GND 0.003621f
C3386 VDD.n3035 GND 0.003621f
C3387 VDD.n3036 GND 0.003621f
C3388 VDD.n3037 GND 0.003621f
C3389 VDD.n3038 GND 0.003621f
C3390 VDD.n3039 GND 0.003621f
C3391 VDD.n3040 GND 0.003621f
C3392 VDD.n3041 GND 0.003621f
C3393 VDD.n3042 GND 0.003621f
C3394 VDD.n3043 GND 0.003621f
C3395 VDD.n3044 GND 0.003621f
C3396 VDD.n3045 GND 0.003621f
C3397 VDD.n3046 GND 0.003621f
C3398 VDD.n3047 GND 0.003621f
C3399 VDD.n3048 GND 0.003621f
C3400 VDD.n3049 GND 0.003621f
C3401 VDD.n3050 GND 0.003621f
C3402 VDD.n3051 GND 0.003621f
C3403 VDD.n3052 GND 0.003621f
C3404 VDD.n3053 GND 0.003621f
C3405 VDD.n3054 GND 0.003621f
C3406 VDD.n3055 GND 0.003621f
C3407 VDD.n3056 GND 0.003621f
C3408 VDD.n3057 GND 0.003621f
C3409 VDD.n3058 GND 0.003621f
C3410 VDD.n3059 GND 0.003621f
C3411 VDD.n3060 GND 0.003621f
C3412 VDD.n3061 GND 0.003621f
C3413 VDD.n3062 GND 0.003621f
C3414 VDD.n3063 GND 0.003621f
C3415 VDD.n3064 GND 0.003621f
C3416 VDD.n3065 GND 0.003621f
C3417 VDD.n3066 GND 0.003621f
C3418 VDD.n3067 GND 0.003621f
C3419 VDD.n3068 GND 0.003621f
C3420 VDD.n3069 GND 0.003621f
C3421 VDD.n3070 GND 0.003621f
C3422 VDD.n3071 GND 0.003621f
C3423 VDD.n3072 GND 0.003621f
C3424 VDD.n3073 GND 0.003621f
C3425 VDD.n3074 GND 0.003621f
C3426 VDD.n3075 GND 0.003621f
C3427 VDD.n3076 GND 0.003621f
C3428 VDD.n3077 GND 0.003621f
C3429 VDD.n3078 GND 0.003621f
C3430 VDD.n3079 GND 0.003621f
C3431 VDD.n3080 GND 0.003621f
C3432 VDD.n3081 GND 0.003621f
C3433 VDD.n3082 GND 0.003621f
C3434 VDD.n3083 GND 0.003621f
C3435 VDD.n3084 GND 0.003621f
C3436 VDD.n3085 GND 0.003621f
C3437 VDD.n3086 GND 0.003621f
C3438 VDD.n3087 GND 0.003621f
C3439 VDD.n3088 GND 0.003621f
C3440 VDD.n3089 GND 0.003621f
C3441 VDD.n3090 GND 0.003621f
C3442 VDD.n3091 GND 0.003621f
C3443 VDD.n3092 GND 0.003621f
C3444 VDD.n3093 GND 0.003621f
C3445 VDD.n3094 GND 0.003621f
C3446 VDD.n3095 GND 0.003621f
C3447 VDD.n3096 GND 0.003621f
C3448 VDD.n3097 GND 0.003621f
C3449 VDD.n3098 GND 0.003621f
C3450 VDD.n3099 GND 0.003621f
C3451 VDD.n3100 GND 0.003621f
C3452 VDD.n3101 GND 0.003621f
C3453 VDD.n3102 GND 0.003621f
C3454 VDD.n3103 GND 0.003621f
C3455 VDD.n3104 GND 0.003621f
C3456 VDD.n3105 GND 0.003621f
C3457 VDD.n3106 GND 0.003621f
C3458 VDD.n3107 GND 0.003621f
C3459 VDD.n3108 GND 0.003621f
C3460 VDD.n3109 GND 0.003621f
C3461 VDD.n3110 GND 0.009198f
C3462 VDD.n3111 GND 0.009198f
C3463 VDD.n3112 GND 0.009198f
C3464 VDD.n3113 GND 0.009548f
C3465 VDD.n3114 GND 0.003621f
C3466 VDD.n3115 GND 0.003621f
C3467 VDD.n3116 GND 0.003621f
C3468 VDD.n3117 GND 0.003621f
C3469 VDD.n3118 GND 0.003621f
C3470 VDD.n3119 GND 0.003621f
C3471 VDD.t120 GND 0.087165f
C3472 VDD.t118 GND 0.39322f
C3473 VDD.n3120 GND 0.070647f
C3474 VDD.t119 GND 0.057758f
C3475 VDD.n3121 GND 0.070509f
C3476 VDD.n3122 GND 0.006279f
C3477 VDD.n3123 GND 0.003621f
C3478 VDD.n3124 GND 0.003621f
C3479 VDD.n3125 GND 0.003621f
C3480 VDD.n3126 GND 0.003621f
C3481 VDD.n3127 GND 0.003621f
C3482 VDD.n3128 GND 0.003621f
C3483 VDD.n3129 GND 0.003621f
C3484 VDD.n3130 GND 0.003621f
C3485 VDD.n3131 GND 0.003621f
C3486 VDD.n3132 GND 0.003621f
C3487 VDD.n3133 GND 0.003621f
C3488 VDD.n3134 GND 0.003621f
C3489 VDD.n3135 GND 0.003621f
C3490 VDD.n3136 GND 0.003621f
C3491 VDD.n3137 GND 0.003621f
C3492 VDD.n3138 GND 0.003621f
C3493 VDD.n3139 GND 0.003621f
C3494 VDD.n3140 GND 0.003621f
C3495 VDD.n3141 GND 0.003621f
C3496 VDD.n3142 GND 0.003621f
C3497 VDD.n3143 GND 0.003621f
C3498 VDD.n3144 GND 0.003621f
C3499 VDD.n3145 GND 0.003621f
C3500 VDD.n3146 GND 0.003621f
C3501 VDD.n3147 GND 0.003621f
C3502 VDD.n3148 GND 0.003621f
C3503 VDD.n3149 GND 0.003621f
C3504 VDD.n3150 GND 0.003621f
C3505 VDD.n3151 GND 0.003621f
C3506 VDD.n3152 GND 0.003621f
C3507 VDD.n3153 GND 0.003621f
C3508 VDD.n3154 GND 0.003621f
C3509 VDD.n3155 GND 0.003621f
C3510 VDD.n3156 GND 0.003621f
C3511 VDD.n3157 GND 0.003621f
C3512 VDD.n3158 GND 0.003621f
C3513 VDD.n3159 GND 0.003621f
C3514 VDD.n3160 GND 0.003621f
C3515 VDD.n3161 GND 0.003621f
C3516 VDD.n3162 GND 0.003621f
C3517 VDD.n3163 GND 0.003621f
C3518 VDD.n3164 GND 0.003621f
C3519 VDD.n3165 GND 0.003621f
C3520 VDD.n3166 GND 0.003621f
C3521 VDD.n3167 GND 0.003621f
C3522 VDD.n3168 GND 0.003621f
C3523 VDD.n3169 GND 0.003621f
C3524 VDD.n3170 GND 0.003621f
C3525 VDD.n3171 GND 0.003621f
C3526 VDD.n3172 GND 0.003621f
C3527 VDD.n3173 GND 0.003621f
C3528 VDD.n3174 GND 0.003621f
C3529 VDD.n3175 GND 0.003621f
C3530 VDD.n3176 GND 0.003621f
C3531 VDD.n3177 GND 0.003621f
C3532 VDD.n3178 GND 0.003621f
C3533 VDD.n3179 GND 0.003621f
C3534 VDD.n3180 GND 0.003621f
C3535 VDD.n3181 GND 0.003621f
C3536 VDD.n3182 GND 0.003621f
C3537 VDD.n3183 GND 0.003621f
C3538 VDD.n3184 GND 0.003621f
C3539 VDD.n3185 GND 0.003621f
C3540 VDD.n3186 GND 0.003621f
C3541 VDD.n3187 GND 0.003621f
C3542 VDD.n3188 GND 0.003621f
C3543 VDD.n3189 GND 0.003621f
C3544 VDD.n3190 GND 0.003621f
C3545 VDD.n3191 GND 0.003621f
C3546 VDD.n3192 GND 0.003621f
C3547 VDD.n3193 GND 0.003621f
C3548 VDD.n3194 GND 0.003621f
C3549 VDD.n3195 GND 0.003621f
C3550 VDD.n3196 GND 0.003621f
C3551 VDD.n3197 GND 0.003621f
C3552 VDD.n3198 GND 0.003621f
C3553 VDD.n3199 GND 0.003621f
C3554 VDD.n3200 GND 0.003621f
C3555 VDD.n3201 GND 0.003621f
C3556 VDD.n3202 GND 0.003621f
C3557 VDD.n3203 GND 0.003621f
C3558 VDD.n3204 GND 0.003621f
C3559 VDD.n3205 GND 0.003621f
C3560 VDD.n3206 GND 0.003621f
C3561 VDD.n3207 GND 0.003621f
C3562 VDD.n3208 GND 0.003621f
C3563 VDD.n3209 GND 0.003621f
C3564 VDD.n3210 GND 0.003621f
C3565 VDD.n3211 GND 0.003621f
C3566 VDD.n3212 GND 0.003621f
C3567 VDD.n3213 GND 0.003621f
C3568 VDD.n3214 GND 0.003621f
C3569 VDD.n3215 GND 0.003621f
C3570 VDD.n3216 GND 0.003621f
C3571 VDD.n3217 GND 0.003621f
C3572 VDD.n3218 GND 0.003621f
C3573 VDD.n3219 GND 0.003621f
C3574 VDD.n3220 GND 0.003621f
C3575 VDD.n3221 GND 0.003621f
C3576 VDD.n3222 GND 0.003621f
C3577 VDD.n3223 GND 0.003621f
C3578 VDD.n3224 GND 0.003621f
C3579 VDD.n3225 GND 0.003621f
C3580 VDD.n3226 GND 0.003621f
C3581 VDD.n3227 GND 0.003621f
C3582 VDD.n3228 GND 0.003621f
C3583 VDD.n3229 GND 0.003621f
C3584 VDD.n3230 GND 0.003621f
C3585 VDD.n3231 GND 0.003621f
C3586 VDD.n3232 GND 0.003621f
C3587 VDD.n3233 GND 0.003621f
C3588 VDD.n3234 GND 0.003621f
C3589 VDD.n3235 GND 0.003621f
C3590 VDD.n3236 GND 0.003621f
C3591 VDD.n3237 GND 0.003621f
C3592 VDD.n3238 GND 0.003621f
C3593 VDD.n3239 GND 0.003621f
C3594 VDD.n3240 GND 0.003621f
C3595 VDD.n3241 GND 0.003621f
C3596 VDD.n3242 GND 0.003621f
C3597 VDD.n3243 GND 0.003621f
C3598 VDD.n3244 GND 0.003621f
C3599 VDD.n3245 GND 0.003621f
C3600 VDD.n3246 GND 0.003621f
C3601 VDD.n3247 GND 0.003621f
C3602 VDD.n3248 GND 0.003621f
C3603 VDD.n3249 GND 0.003621f
C3604 VDD.n3250 GND 0.003621f
C3605 VDD.n3251 GND 0.003621f
C3606 VDD.n3252 GND 0.003621f
C3607 VDD.n3253 GND 0.003621f
C3608 VDD.n3254 GND 0.003621f
C3609 VDD.n3255 GND 0.003621f
C3610 VDD.n3256 GND 0.003621f
C3611 VDD.n3257 GND 0.003621f
C3612 VDD.n3258 GND 0.003621f
C3613 VDD.n3259 GND 0.003621f
C3614 VDD.n3260 GND 0.003621f
C3615 VDD.n3261 GND 0.003621f
C3616 VDD.n3262 GND 0.003621f
C3617 VDD.n3263 GND 0.003621f
C3618 VDD.n3264 GND 0.003621f
C3619 VDD.n3265 GND 0.003621f
C3620 VDD.n3266 GND 0.003621f
C3621 VDD.n3267 GND 0.003621f
C3622 VDD.n3268 GND 0.003621f
C3623 VDD.n3269 GND 0.003621f
C3624 VDD.n3270 GND 0.003621f
C3625 VDD.n3271 GND 0.003621f
C3626 VDD.n3272 GND 0.003621f
C3627 VDD.n3273 GND 0.003621f
C3628 VDD.n3274 GND 0.003621f
C3629 VDD.n3275 GND 0.003621f
C3630 VDD.n3276 GND 0.003621f
C3631 VDD.n3277 GND 0.003621f
C3632 VDD.n3278 GND 0.003621f
C3633 VDD.n3279 GND 0.003621f
C3634 VDD.n3280 GND 0.003621f
C3635 VDD.n3281 GND 0.003621f
C3636 VDD.n3282 GND 0.003621f
C3637 VDD.n3283 GND 0.003621f
C3638 VDD.n3284 GND 0.003621f
C3639 VDD.n3285 GND 0.003621f
C3640 VDD.n3286 GND 0.003621f
C3641 VDD.n3287 GND 0.003621f
C3642 VDD.n3288 GND 0.003621f
C3643 VDD.n3289 GND 0.003621f
C3644 VDD.n3290 GND 0.003621f
C3645 VDD.n3291 GND 0.003621f
C3646 VDD.n3292 GND 0.003621f
C3647 VDD.n3293 GND 0.003621f
C3648 VDD.n3294 GND 0.003621f
C3649 VDD.n3295 GND 0.003621f
C3650 VDD.n3296 GND 0.009198f
C3651 VDD.n3298 GND 0.009548f
C3652 VDD.n3299 GND 0.009548f
C3653 VDD.n3300 GND 0.003621f
C3654 VDD.n3301 GND 0.003621f
C3655 VDD.n3302 GND 0.003621f
C3656 VDD.n3304 GND 0.003621f
C3657 VDD.n3306 GND 0.003621f
C3658 VDD.n3307 GND 0.003621f
C3659 VDD.n3308 GND 0.003621f
C3660 VDD.n3309 GND 0.003621f
C3661 VDD.n3310 GND 0.003621f
C3662 VDD.n3312 GND 0.003621f
C3663 VDD.n3314 GND 0.003621f
C3664 VDD.n3315 GND 0.003621f
C3665 VDD.n3316 GND 0.003621f
C3666 VDD.n3317 GND 0.003621f
C3667 VDD.n3318 GND 0.003621f
C3668 VDD.n3320 GND 0.003621f
C3669 VDD.n3322 GND 0.003621f
C3670 VDD.n3323 GND 0.003621f
C3671 VDD.n3324 GND 0.003621f
C3672 VDD.n3325 GND 0.003621f
C3673 VDD.n3326 GND 0.003621f
C3674 VDD.n3328 GND 0.003621f
C3675 VDD.n3330 GND 0.003621f
C3676 VDD.n3331 GND 0.003621f
C3677 VDD.n3332 GND 0.009548f
C3678 VDD.n3333 GND 0.009198f
C3679 VDD.n3334 GND 0.009198f
C3680 VDD.n3335 GND 0.60703f
C3681 VDD.n3336 GND 0.009198f
C3682 VDD.n3337 GND 0.009198f
C3683 VDD.n3338 GND 0.003621f
C3684 VDD.n3339 GND 0.003621f
C3685 VDD.n3340 GND 0.003621f
C3686 VDD.n3341 GND 0.395005f
C3687 VDD.n3342 GND 0.003621f
C3688 VDD.n3343 GND 0.003621f
C3689 VDD.n3344 GND 0.003621f
C3690 VDD.n3345 GND 0.003621f
C3691 VDD.n3346 GND 0.003621f
C3692 VDD.n3347 GND 0.395005f
C3693 VDD.n3348 GND 0.003621f
C3694 VDD.n3349 GND 0.003621f
C3695 VDD.n3350 GND 0.003621f
C3696 VDD.n3351 GND 0.003621f
C3697 VDD.n3352 GND 0.003621f
C3698 VDD.n3353 GND 0.395005f
C3699 VDD.n3354 GND 0.003621f
C3700 VDD.n3355 GND 0.003621f
C3701 VDD.n3356 GND 0.003621f
C3702 VDD.n3357 GND 0.003621f
C3703 VDD.n3358 GND 0.003621f
C3704 VDD.n3359 GND 0.395005f
C3705 VDD.n3360 GND 0.003621f
C3706 VDD.n3361 GND 0.003621f
C3707 VDD.n3362 GND 0.003621f
C3708 VDD.n3363 GND 0.003621f
C3709 VDD.n3364 GND 0.003621f
C3710 VDD.n3365 GND 0.212025f
C3711 VDD.n3366 GND 0.003621f
C3712 VDD.n3367 GND 0.003621f
C3713 VDD.n3368 GND 0.003621f
C3714 VDD.n3369 GND 0.003621f
C3715 VDD.n3370 GND 0.003621f
C3716 VDD.n3371 GND 0.395005f
C3717 VDD.n3372 GND 0.003621f
C3718 VDD.n3373 GND 0.003621f
C3719 VDD.n3374 GND 0.003621f
C3720 VDD.n3375 GND 0.003621f
C3721 VDD.n3376 GND 0.003621f
C3722 VDD.n3377 GND 0.395005f
C3723 VDD.n3378 GND 0.003621f
C3724 VDD.n3379 GND 0.003621f
C3725 VDD.n3380 GND 0.003621f
C3726 VDD.n3381 GND 0.003621f
C3727 VDD.n3382 GND 0.003621f
C3728 VDD.n3383 GND 0.395005f
C3729 VDD.n3384 GND 0.003621f
C3730 VDD.n3385 GND 0.003621f
C3731 VDD.n3386 GND 0.003621f
C3732 VDD.n3387 GND 0.003621f
C3733 VDD.n3388 GND 0.003621f
C3734 VDD.n3389 GND 0.395005f
C3735 VDD.n3390 GND 0.003621f
C3736 VDD.n3391 GND 0.003621f
C3737 VDD.n3392 GND 0.003621f
C3738 VDD.n3393 GND 0.003621f
C3739 VDD.n3394 GND 0.003621f
C3740 VDD.n3395 GND 0.395005f
C3741 VDD.n3396 GND 0.003621f
C3742 VDD.n3397 GND 0.003621f
C3743 VDD.n3398 GND 0.003621f
C3744 VDD.n3399 GND 0.003621f
C3745 VDD.n3400 GND 0.003621f
C3746 VDD.n3401 GND 0.395005f
C3747 VDD.n3402 GND 0.003621f
C3748 VDD.n3403 GND 0.003621f
C3749 VDD.n3404 GND 0.003621f
C3750 VDD.n3405 GND 0.003621f
C3751 VDD.n3406 GND 0.003621f
C3752 VDD.n3407 GND 0.395005f
C3753 VDD.n3408 GND 0.003621f
C3754 VDD.n3409 GND 0.003621f
C3755 VDD.n3410 GND 0.003621f
C3756 VDD.n3411 GND 0.003621f
C3757 VDD.n3412 GND 0.003621f
C3758 VDD.n3413 GND 0.395005f
C3759 VDD.n3414 GND 0.003621f
C3760 VDD.n3415 GND 0.003621f
C3761 VDD.n3416 GND 0.003621f
C3762 VDD.n3417 GND 0.003621f
C3763 VDD.n3418 GND 0.003621f
C3764 VDD.n3419 GND 0.29335f
C3765 VDD.n3420 GND 0.003621f
C3766 VDD.n3421 GND 0.003621f
C3767 VDD.n3422 GND 0.003621f
C3768 VDD.n3423 GND 0.003621f
C3769 VDD.n3424 GND 0.003621f
C3770 VDD.n3425 GND 0.395005f
C3771 VDD.n3426 GND 0.003621f
C3772 VDD.n3427 GND 0.003621f
C3773 VDD.n3428 GND 0.003621f
C3774 VDD.n3429 GND 0.003621f
C3775 VDD.n3430 GND 0.003621f
C3776 VDD.n3431 GND 0.246878f
C3777 VDD.n3432 GND 0.003621f
C3778 VDD.n3433 GND 0.003621f
C3779 VDD.n3434 GND 0.003621f
C3780 VDD.n3435 GND 0.003621f
C3781 VDD.n3436 GND 0.003621f
C3782 VDD.n3437 GND 0.395005f
C3783 VDD.n3438 GND 0.003621f
C3784 VDD.n3439 GND 0.003621f
C3785 VDD.n3440 GND 0.003621f
C3786 VDD.n3441 GND 0.003621f
C3787 VDD.n3442 GND 0.003621f
C3788 VDD.n3443 GND 0.395005f
C3789 VDD.n3444 GND 0.003621f
C3790 VDD.n3445 GND 0.003621f
C3791 VDD.n3446 GND 0.003621f
C3792 VDD.n3447 GND 0.003621f
C3793 VDD.n3448 GND 0.003621f
C3794 VDD.n3449 GND 0.395005f
C3795 VDD.n3450 GND 0.003621f
C3796 VDD.n3451 GND 0.003621f
C3797 VDD.n3452 GND 0.003621f
C3798 VDD.n3453 GND 0.003621f
C3799 VDD.n3454 GND 0.003621f
C3800 VDD.n3455 GND 0.395005f
C3801 VDD.n3456 GND 0.003621f
C3802 VDD.n3457 GND 0.003621f
C3803 VDD.n3458 GND 0.003621f
C3804 VDD.n3459 GND 0.003621f
C3805 VDD.n3460 GND 0.003621f
C3806 VDD.n3461 GND 0.395005f
C3807 VDD.n3462 GND 0.003621f
C3808 VDD.n3463 GND 0.003621f
C3809 VDD.n3464 GND 0.003621f
C3810 VDD.n3465 GND 0.003621f
C3811 VDD.n3466 GND 0.003621f
C3812 VDD.n3467 GND 0.395005f
C3813 VDD.n3468 GND 0.003621f
C3814 VDD.n3469 GND 0.003621f
C3815 VDD.n3470 GND 0.003621f
C3816 VDD.n3471 GND 0.003621f
C3817 VDD.n3472 GND 0.003621f
C3818 VDD.n3473 GND 0.200407f
C3819 VDD.n3474 GND 0.003621f
C3820 VDD.n3475 GND 0.003621f
C3821 VDD.n3476 GND 0.003621f
C3822 VDD.n3477 GND 0.003621f
C3823 VDD.n3478 GND 0.003621f
C3824 VDD.n3479 GND 0.395005f
C3825 VDD.n3480 GND 0.003621f
C3826 VDD.n3481 GND 0.003621f
C3827 VDD.n3482 GND 0.003621f
C3828 VDD.n3483 GND 0.003621f
C3829 VDD.n3484 GND 0.003621f
C3830 VDD.n3485 GND 0.34563f
C3831 VDD.n3486 GND 0.003621f
C3832 VDD.n3487 GND 0.003621f
C3833 VDD.n3488 GND 0.003621f
C3834 VDD.n3489 GND 0.003621f
C3835 VDD.n3490 GND 0.003621f
C3836 VDD.n3491 GND 0.395005f
C3837 VDD.n3492 GND 0.003621f
C3838 VDD.n3493 GND 0.003621f
C3839 VDD.n3494 GND 0.003621f
C3840 VDD.n3495 GND 0.003621f
C3841 VDD.n3496 GND 0.003621f
C3842 VDD.n3497 GND 0.395005f
C3843 VDD.n3498 GND 0.003621f
C3844 VDD.n3499 GND 0.003621f
C3845 VDD.n3500 GND 0.003621f
C3846 VDD.n3501 GND 0.003621f
C3847 VDD.n3502 GND 0.003621f
C3848 VDD.n3503 GND 0.395005f
C3849 VDD.n3504 GND 0.003621f
C3850 VDD.n3505 GND 0.003621f
C3851 VDD.n3506 GND 0.003621f
C3852 VDD.n3507 GND 0.003621f
C3853 VDD.n3508 GND 0.003621f
C3854 VDD.n3509 GND 0.395005f
C3855 VDD.n3510 GND 0.003621f
C3856 VDD.n3511 GND 0.003621f
C3857 VDD.n3512 GND 0.003621f
C3858 VDD.n3513 GND 0.003621f
C3859 VDD.n3514 GND 0.003621f
C3860 VDD.n3515 GND 0.395005f
C3861 VDD.n3516 GND 0.003621f
C3862 VDD.n3517 GND 0.003621f
C3863 VDD.n3518 GND 0.003621f
C3864 VDD.n3519 GND 0.003621f
C3865 VDD.n3520 GND 0.003621f
C3866 VDD.n3521 GND 0.395005f
C3867 VDD.n3522 GND 0.003621f
C3868 VDD.n3523 GND 0.003621f
C3869 VDD.n3524 GND 0.003621f
C3870 VDD.n3525 GND 0.003621f
C3871 VDD.n3526 GND 0.003621f
C3872 VDD.n3527 GND 0.299158f
C3873 VDD.n3528 GND 0.003621f
C3874 VDD.n3529 GND 0.003621f
C3875 VDD.n3530 GND 0.003621f
C3876 VDD.n3531 GND 0.003621f
C3877 VDD.n3532 GND 0.003621f
C3878 VDD.n3533 GND 0.34563f
C3879 VDD.n3534 GND 0.003621f
C3880 VDD.n3535 GND 0.003621f
C3881 VDD.n3536 GND 0.003621f
C3882 VDD.n3537 GND 0.003621f
C3883 VDD.n3538 GND 0.003621f
C3884 VDD.n3539 GND 0.395005f
C3885 VDD.n3540 GND 0.003621f
C3886 VDD.n3541 GND 0.003621f
C3887 VDD.n3542 GND 0.003621f
C3888 VDD.n3543 GND 0.003621f
C3889 VDD.n3544 GND 0.003621f
C3890 VDD.n3545 GND 0.395005f
C3891 VDD.n3546 GND 0.003621f
C3892 VDD.n3547 GND 0.003621f
C3893 VDD.n3548 GND 0.003621f
C3894 VDD.n3549 GND 0.003621f
C3895 VDD.n3550 GND 0.003621f
C3896 VDD.n3551 GND 0.395005f
C3897 VDD.n3552 GND 0.003621f
C3898 VDD.n3553 GND 0.003621f
C3899 VDD.n3554 GND 0.003621f
C3900 VDD.n3555 GND 0.003621f
C3901 VDD.n3556 GND 0.003621f
C3902 VDD.n3557 GND 0.395005f
C3903 VDD.n3558 GND 0.003621f
C3904 VDD.n3559 GND 0.003621f
C3905 VDD.n3560 GND 0.003621f
C3906 VDD.n3561 GND 0.003621f
C3907 VDD.n3562 GND 0.003621f
C3908 VDD.n3563 GND 0.395005f
C3909 VDD.n3564 GND 0.003621f
C3910 VDD.n3565 GND 0.003621f
C3911 VDD.n3566 GND 0.003621f
C3912 VDD.n3567 GND 0.003621f
C3913 VDD.n3568 GND 0.003621f
C3914 VDD.n3569 GND 0.395005f
C3915 VDD.n3570 GND 0.003621f
C3916 VDD.n3571 GND 0.003621f
C3917 VDD.n3572 GND 0.003621f
C3918 VDD.n3573 GND 0.003621f
C3919 VDD.n3574 GND 0.003621f
C3920 VDD.n3575 GND 0.395005f
C3921 VDD.n3576 GND 0.003621f
C3922 VDD.n3577 GND 0.003621f
C3923 VDD.n3578 GND 0.003621f
C3924 VDD.n3579 GND 0.003621f
C3925 VDD.n3580 GND 0.003621f
C3926 VDD.n3581 GND 0.395005f
C3927 VDD.n3582 GND 0.003621f
C3928 VDD.n3583 GND 0.003621f
C3929 VDD.n3584 GND 0.003621f
C3930 VDD.n3585 GND 0.003621f
C3931 VDD.n3586 GND 0.003621f
C3932 VDD.n3587 GND 0.246878f
C3933 VDD.n3588 GND 0.003621f
C3934 VDD.n3589 GND 0.003621f
C3935 VDD.n3590 GND 0.003621f
C3936 VDD.n3591 GND 0.003621f
C3937 VDD.n3592 GND 0.003621f
C3938 VDD.n3593 GND 0.395005f
C3939 VDD.n3594 GND 0.003621f
C3940 VDD.n3595 GND 0.003621f
C3941 VDD.n3596 GND 0.003621f
C3942 VDD.n3597 GND 0.003621f
C3943 VDD.n3598 GND 0.003621f
C3944 VDD.n3599 GND 0.395005f
C3945 VDD.n3600 GND 0.003621f
C3946 VDD.n3601 GND 0.003621f
C3947 VDD.n3602 GND 0.003621f
C3948 VDD.n3603 GND 0.003621f
C3949 VDD.n3604 GND 0.003621f
C3950 VDD.n3605 GND 0.313681f
C3951 VDD.n3606 GND 0.003621f
C3952 VDD.n3607 GND 0.003621f
C3953 VDD.n3608 GND 0.003621f
C3954 VDD.n3609 GND 0.003621f
C3955 VDD.n3610 GND 0.003621f
C3956 VDD.n3611 GND 0.395005f
C3957 VDD.n3612 GND 0.003621f
C3958 VDD.n3613 GND 0.003621f
C3959 VDD.n3614 GND 0.003621f
C3960 VDD.n3615 GND 0.003621f
C3961 VDD.n3616 GND 0.003621f
C3962 VDD.n3617 GND 0.395005f
C3963 VDD.n3618 GND 0.003621f
C3964 VDD.n3619 GND 0.003621f
C3965 VDD.n3620 GND 0.003621f
C3966 VDD.n3621 GND 0.003621f
C3967 VDD.n3622 GND 0.003621f
C3968 VDD.n3623 GND 0.395005f
C3969 VDD.n3624 GND 0.003621f
C3970 VDD.n3625 GND 0.003621f
C3971 VDD.n3626 GND 0.003621f
C3972 VDD.n3627 GND 0.003621f
C3973 VDD.n3628 GND 0.003621f
C3974 VDD.n3629 GND 0.395005f
C3975 VDD.n3630 GND 0.003621f
C3976 VDD.n3631 GND 0.003621f
C3977 VDD.n3632 GND 0.003621f
C3978 VDD.n3633 GND 0.003621f
C3979 VDD.n3634 GND 0.003621f
C3980 VDD.n3635 GND 0.395005f
C3981 VDD.n3636 GND 0.003621f
C3982 VDD.n3637 GND 0.003621f
C3983 VDD.n3638 GND 0.003621f
C3984 VDD.n3639 GND 0.003621f
C3985 VDD.n3640 GND 0.003621f
C3986 VDD.n3641 GND 0.395005f
C3987 VDD.n3642 GND 0.003621f
C3988 VDD.n3643 GND 0.003621f
C3989 VDD.n3644 GND 0.003621f
C3990 VDD.n3645 GND 0.003621f
C3991 VDD.n3646 GND 0.003621f
C3992 VDD.n3647 GND 0.395005f
C3993 VDD.n3648 GND 0.003621f
C3994 VDD.n3649 GND 0.003621f
C3995 VDD.n3650 GND 0.003621f
C3996 VDD.n3651 GND 0.003621f
C3997 VDD.n3652 GND 0.003621f
C3998 VDD.n3653 GND 0.194598f
C3999 VDD.n3654 GND 0.003621f
C4000 VDD.n3655 GND 0.003621f
C4001 VDD.n3656 GND 0.003621f
C4002 VDD.n3657 GND 0.003621f
C4003 VDD.n3658 GND 0.003621f
C4004 VDD.n3659 GND 0.395005f
C4005 VDD.n3660 GND 0.003621f
C4006 VDD.n3661 GND 0.003621f
C4007 VDD.n3662 GND 0.003621f
C4008 VDD.n3663 GND 0.003621f
C4009 VDD.n3664 GND 0.003621f
C4010 VDD.n3665 GND 0.395005f
C4011 VDD.n3666 GND 0.003621f
C4012 VDD.n3667 GND 0.003621f
C4013 VDD.n3668 GND 0.003621f
C4014 VDD.n3669 GND 0.003621f
C4015 VDD.n3670 GND 0.003621f
C4016 VDD.n3671 GND 0.003621f
C4017 VDD.n3672 GND 0.003621f
C4018 VDD.n3674 GND 0.003621f
C4019 VDD.n3675 GND 0.003621f
C4020 VDD.n3676 GND 0.003621f
C4021 VDD.n3678 GND 0.003621f
C4022 VDD.n3679 GND 0.003621f
C4023 VDD.n3680 GND 0.003621f
C4024 VDD.n3681 GND 0.003621f
C4025 VDD.n3682 GND 0.003621f
C4026 VDD.n3683 GND 0.003621f
C4027 VDD.n3685 GND 0.003621f
C4028 VDD.n3686 GND 0.003621f
C4029 VDD.n3688 GND 0.009548f
C4030 VDD.n3689 GND 0.009548f
C4031 VDD.n3690 GND 0.009198f
C4032 VDD.n3691 GND 0.003621f
C4033 VDD.n3692 GND 0.003621f
C4034 VDD.n3693 GND 0.003621f
C4035 VDD.n3694 GND 0.003621f
C4036 VDD.n3695 GND 0.003621f
C4037 VDD.n3696 GND 0.003621f
C4038 VDD.n3697 GND 0.395005f
C4039 VDD.n3698 GND 0.003621f
C4040 VDD.n3699 GND 0.003621f
C4041 VDD.n3700 GND 0.003621f
C4042 VDD.n3701 GND 0.003621f
C4043 VDD.n3702 GND 0.003621f
C4044 VDD.n3703 GND 0.395005f
C4045 VDD.n3704 GND 0.003621f
C4046 VDD.n3705 GND 0.003621f
C4047 VDD.n3706 GND 0.003621f
C4048 VDD.n3707 GND 0.009566f
C4049 VDD.n3708 GND 0.00918f
C4050 VDD.n3709 GND 0.009548f
C4051 VDD.n3711 GND 0.003621f
C4052 VDD.n3712 GND 0.003621f
C4053 VDD.n3713 GND 0.003621f
C4054 VDD.n3714 GND 0.006279f
C4055 VDD.n3715 GND 0.003621f
C4056 VDD.n3716 GND 0.003621f
C4057 VDD.n3718 GND 0.003621f
C4058 VDD.n3719 GND 0.003621f
C4059 VDD.n3720 GND 0.003621f
C4060 VDD.n3721 GND 0.003621f
C4061 VDD.n3722 GND 0.002716f
C4062 VDD.n3723 GND 0.003621f
C4063 VDD.n3725 GND 0.003621f
C4064 VDD.n3726 GND 0.002716f
C4065 VDD.n3727 GND 0.003621f
C4066 VDD.n3728 GND 0.003621f
C4067 VDD.n3730 GND 0.003621f
C4068 VDD.n3731 GND 0.003621f
C4069 VDD.n3732 GND 0.003621f
C4070 VDD.n3733 GND 0.003621f
C4071 VDD.n3734 GND 0.003621f
C4072 VDD.n3735 GND 0.003621f
C4073 VDD.n3737 GND 0.003621f
C4074 VDD.n3738 GND 0.003621f
C4075 VDD.n3739 GND 0.003621f
C4076 VDD.n3740 GND 0.009548f
C4077 VDD.n3741 GND 0.009198f
C4078 VDD.n3742 GND 0.009198f
C4079 VDD.n3743 GND 0.60703f
C4080 VDD.n3744 GND 0.009198f
C4081 VDD.n3745 GND 0.009548f
C4082 VDD.n3746 GND 0.00918f
C4083 VDD.n3747 GND 0.003621f
C4084 VDD.n3748 GND 0.003621f
C4085 VDD.n3749 GND 0.003621f
C4086 VDD.n3751 GND 0.003621f
C4087 VDD.n3752 GND 0.003621f
C4088 VDD.n3753 GND 0.003621f
C4089 VDD.n3754 GND 0.003621f
C4090 VDD.n3755 GND 0.003621f
C4091 VDD.n3756 GND 0.003621f
C4092 VDD.n3758 GND 0.003621f
C4093 VDD.n3759 GND 0.003621f
C4094 VDD.n3760 GND 0.002716f
C4095 VDD.n3761 GND 0.078438f
C4096 VDD.n3762 GND 1.11224f
C4097 VDD.n3763 GND 0.004207f
C4098 VDD.n3764 GND 0.004287f
C4099 VDD.n3765 GND 0.005326f
C4100 VDD.n3766 GND 0.005326f
C4101 VDD.n3767 GND 0.005326f
C4102 VDD.n3768 GND 0.002936f
C4103 VDD.n3769 GND 0.005326f
C4104 VDD.n3770 GND 0.004287f
C4105 VDD.n3772 GND 0.005326f
C4106 VDD.n3774 GND 0.005326f
C4107 VDD.n3775 GND 0.005326f
C4108 VDD.n3776 GND 0.004287f
C4109 VDD.n3777 GND 0.005326f
C4110 VDD.n3778 GND 0.005326f
C4111 VDD.n3779 GND 0.005326f
C4112 VDD.n3780 GND 0.005326f
C4113 VDD.n3781 GND 0.005326f
C4114 VDD.n3782 GND 0.004287f
C4115 VDD.n3783 GND 0.005326f
C4116 VDD.n3784 GND 0.005326f
C4117 VDD.n3785 GND 0.005326f
C4118 VDD.n3786 GND 0.005326f
C4119 VDD.n3787 GND 0.005326f
C4120 VDD.n3788 GND 0.004287f
C4121 VDD.n3789 GND 0.005326f
C4122 VDD.n3790 GND 0.005326f
C4123 VDD.n3791 GND 0.005326f
C4124 VDD.n3792 GND 0.002272f
C4125 VDD.n3794 GND 0.005326f
C4126 VDD.t102 GND 0.159105f
C4127 VDD.t100 GND 0.597454f
C4128 VDD.n3795 GND 0.084294f
C4129 VDD.t101 GND 0.119732f
C4130 VDD.n3796 GND 0.085079f
C4131 VDD.n3797 GND 0.008037f
C4132 VDD.n3798 GND 0.005326f
C4133 VDD.n3799 GND 0.005326f
C4134 VDD.n3800 GND 0.004158f
C4135 VDD.n3801 GND 0.004287f
C4136 VDD.n3802 GND 0.005326f
C4137 VDD.n3804 GND 0.005326f
C4138 VDD.n3806 GND 0.005326f
C4139 VDD.n3807 GND 0.004287f
C4140 VDD.n3808 GND 0.004287f
C4141 VDD.n3809 GND 0.004287f
C4142 VDD.n3810 GND 0.005326f
C4143 VDD.n3812 GND 0.005326f
C4144 VDD.n3814 GND 0.005326f
C4145 VDD.n3815 GND 0.004287f
C4146 VDD.n3816 GND 0.004287f
C4147 VDD.n3817 GND 0.004287f
C4148 VDD.n3818 GND 0.005326f
C4149 VDD.n3820 GND 0.005326f
C4150 VDD.n3821 GND 0.005326f
C4151 VDD.n3822 GND 0.004287f
C4152 VDD.n3823 GND 0.004287f
C4153 VDD.n3824 GND 0.005326f
C4154 VDD.n3825 GND 0.005326f
C4155 VDD.n3827 GND 0.005326f
C4156 VDD.n3828 GND 0.004287f
C4157 VDD.n3829 GND 0.005326f
C4158 VDD.n3830 GND 0.005326f
C4159 VDD.n3831 GND 0.005326f
C4160 VDD.t113 GND 0.117451f
C4161 VDD.t114 GND 0.160644f
C4162 VDD.t112 GND 0.597454f
C4163 VDD.n3832 GND 0.084171f
C4164 VDD.n3833 GND 0.084531f
C4165 VDD.n3834 GND 0.009452f
C4166 VDD.n3835 GND 0.004222f
C4167 VDD.n3836 GND 0.005326f
C4168 VDD.n3838 GND 0.005326f
C4169 VDD.n3839 GND 0.005326f
C4170 VDD.n3840 GND 0.004287f
C4171 VDD.n3841 GND 0.004287f
C4172 VDD.n3842 GND 0.005326f
C4173 VDD.n3843 GND 0.005326f
C4174 VDD.n3844 GND 0.004287f
C4175 VDD.n3845 GND 0.004287f
C4176 VDD.n3846 GND 0.005326f
C4177 VDD.n3848 GND 0.005326f
C4178 VDD.n3849 GND 0.004287f
C4179 VDD.n3850 GND 0.004287f
C4180 VDD.n3851 GND 0.004287f
C4181 VDD.n3852 GND 0.005326f
C4182 VDD.n3854 GND 0.005326f
C4183 VDD.n3856 GND 0.005326f
C4184 VDD.n3857 GND 0.004287f
C4185 VDD.n3858 GND 0.004287f
C4186 VDD.n3859 GND 0.004287f
C4187 VDD.n3860 GND 0.005326f
C4188 VDD.n3862 GND 0.005326f
C4189 VDD.n3864 GND 0.005326f
C4190 VDD.n3865 GND 0.004287f
C4191 VDD.n3866 GND 0.002872f
C4192 VDD.n3867 GND 0.008037f
C4193 VDD.n3868 GND 0.005326f
C4194 VDD.n3870 GND 0.005326f
C4195 VDD.n3872 GND 0.005326f
C4196 VDD.n3873 GND 0.004287f
C4197 VDD.n3874 GND 0.004287f
C4198 VDD.n3875 GND 0.004287f
C4199 VDD.n3876 GND 0.005326f
C4200 VDD.n3878 GND 0.005326f
C4201 VDD.n3880 GND 0.005326f
C4202 VDD.n3881 GND 0.004287f
C4203 VDD.n3882 GND 0.004287f
C4204 VDD.n3883 GND 0.004287f
C4205 VDD.n3884 GND 0.005326f
C4206 VDD.n3886 GND 0.005326f
C4207 VDD.n3888 GND 0.005326f
C4208 VDD.n3889 GND 0.004287f
C4209 VDD.n3890 GND 0.004287f
C4210 VDD.n3891 GND 0.004287f
C4211 VDD.n3892 GND 0.005326f
C4212 VDD.n3894 GND 0.005326f
C4213 VDD.n3896 GND 0.005326f
C4214 VDD.n3897 GND 0.004287f
C4215 VDD.n3898 GND 0.004287f
C4216 VDD.n3899 GND 0.002808f
C4217 VDD.n3900 GND 0.005326f
C4218 VDD.n3902 GND 0.005326f
C4219 VDD.n3904 GND 0.005326f
C4220 VDD.n3905 GND 0.004287f
C4221 VDD.n3906 GND 0.004287f
C4222 VDD.n3907 GND 0.004287f
C4223 VDD.n3908 GND 0.005326f
C4224 VDD.n3910 GND 0.005326f
C4225 VDD.n3912 GND 0.005326f
C4226 VDD.n3913 GND 0.004287f
C4227 VDD.n3914 GND 0.004287f
C4228 VDD.n3916 GND 0.004207f
C4229 VDD.n3917 GND 1.11224f
C4230 VDD.n3919 GND 0.004287f
C4231 VDD.n3920 GND 0.005326f
C4232 VDD.n3922 GND 0.005326f
C4233 VDD.n3924 GND 0.005326f
C4234 VDD.n3925 GND 0.004287f
C4235 VDD.n3926 GND 0.004287f
C4236 VDD.n3927 GND 0.004287f
C4237 VDD.n3928 GND 0.005326f
C4238 VDD.n3930 GND 0.005326f
C4239 VDD.n3932 GND 0.005326f
C4240 VDD.n3933 GND 0.004287f
C4241 VDD.n3934 GND 0.002743f
C4242 VDD.n3935 GND 0.005894f
C4243 VDD.n3936 GND 0.002272f
C4244 VDD.n3937 GND 0.005326f
C4245 VDD.n3939 GND 0.005326f
C4246 VDD.n3941 GND 0.005326f
C4247 VDD.n3942 GND 0.004287f
C4248 VDD.n3943 GND 0.004287f
C4249 VDD.n3944 GND 0.004287f
C4250 VDD.n3945 GND 0.005326f
C4251 VDD.n3947 GND 0.005326f
C4252 VDD.n3949 GND 0.005326f
C4253 VDD.n3950 GND 0.004287f
C4254 VDD.n3951 GND 0.004287f
C4255 VDD.n3952 GND 0.004287f
C4256 VDD.n3953 GND 0.005326f
C4257 VDD.n3955 GND 0.005326f
C4258 VDD.n3956 GND 0.005326f
C4259 VDD.n3957 GND 0.004287f
C4260 VDD.n3958 GND 0.004287f
C4261 VDD.n3959 GND 0.005326f
C4262 VDD.n3960 GND 0.005326f
C4263 VDD.n3962 GND 0.005326f
C4264 VDD.n3963 GND 0.004287f
C4265 VDD.n3964 GND 0.003558f
C4266 VDD.n3965 GND 0.012553f
C4267 VDD.n3966 GND 0.012264f
C4268 VDD.n3967 GND 0.003558f
C4269 VDD.n3968 GND 0.012264f
C4270 VDD.n3969 GND 0.824864f
C4271 VDD.n3970 GND 0.012264f
C4272 VDD.n3971 GND 0.003558f
C4273 VDD.n3972 GND 0.012264f
C4274 VDD.n3973 GND 0.005326f
C4275 VDD.n3974 GND 0.005326f
C4276 VDD.n3975 GND 0.004287f
C4277 VDD.n3976 GND 0.005326f
C4278 VDD.n3977 GND 0.58089f
C4279 VDD.n3978 GND 0.005326f
C4280 VDD.n3979 GND 0.004287f
C4281 VDD.n3980 GND 0.005326f
C4282 VDD.n3981 GND 0.005326f
C4283 VDD.n3982 GND 0.005326f
C4284 VDD.n3983 GND 0.004287f
C4285 VDD.n3984 GND 0.005326f
C4286 VDD.n3985 GND 0.58089f
C4287 VDD.n3986 GND 0.005326f
C4288 VDD.n3987 GND 0.004287f
C4289 VDD.n3988 GND 0.005326f
C4290 VDD.n3989 GND 0.005326f
C4291 VDD.n3990 GND 0.005326f
C4292 VDD.n3991 GND 0.004287f
C4293 VDD.n3992 GND 0.005326f
C4294 VDD.n3993 GND 0.360152f
C4295 VDD.n3994 GND 0.005326f
C4296 VDD.n3995 GND 0.004287f
C4297 VDD.n3996 GND 0.005326f
C4298 VDD.n3997 GND 0.005326f
C4299 VDD.n3998 GND 0.005326f
C4300 VDD.n3999 GND 0.004287f
C4301 VDD.n4000 GND 0.005326f
C4302 VDD.n4001 GND 0.58089f
C4303 VDD.n4002 GND 0.005326f
C4304 VDD.n4003 GND 0.004287f
C4305 VDD.n4004 GND 0.005326f
C4306 VDD.n4005 GND 0.005326f
C4307 VDD.n4006 GND 0.005326f
C4308 VDD.n4007 GND 0.004287f
C4309 VDD.n4008 GND 0.005326f
C4310 VDD.n4009 GND 0.58089f
C4311 VDD.n4010 GND 0.005326f
C4312 VDD.n4011 GND 0.004287f
C4313 VDD.n4012 GND 0.005326f
C4314 VDD.n4013 GND 0.005326f
C4315 VDD.n4014 GND 0.005326f
C4316 VDD.n4015 GND 0.004287f
C4317 VDD.n4016 GND 0.005326f
C4318 VDD.n4017 GND 0.58089f
C4319 VDD.n4018 GND 0.005326f
C4320 VDD.n4019 GND 0.004287f
C4321 VDD.n4020 GND 0.005326f
C4322 VDD.n4021 GND 0.005326f
C4323 VDD.n4022 GND 0.005326f
C4324 VDD.n4023 GND 0.004287f
C4325 VDD.n4024 GND 0.005326f
C4326 VDD.n4025 GND 0.58089f
C4327 VDD.n4026 GND 0.005326f
C4328 VDD.n4027 GND 0.004287f
C4329 VDD.n4028 GND 0.005326f
C4330 VDD.n4029 GND 0.005326f
C4331 VDD.n4030 GND 0.005326f
C4332 VDD.n4031 GND 0.004287f
C4333 VDD.n4032 GND 0.005326f
C4334 VDD.n4033 GND 0.58089f
C4335 VDD.n4034 GND 0.005326f
C4336 VDD.n4035 GND 0.004287f
C4337 VDD.n4036 GND 0.005326f
C4338 VDD.n4037 GND 0.005326f
C4339 VDD.n4038 GND 0.005326f
C4340 VDD.n4039 GND 0.004287f
C4341 VDD.n4040 GND 0.005326f
C4342 VDD.n4041 GND 0.377579f
C4343 VDD.n4042 GND 0.58089f
C4344 VDD.n4043 GND 0.005326f
C4345 VDD.n4044 GND 0.004287f
C4346 VDD.n4045 GND 0.005326f
C4347 VDD.n4046 GND 0.005326f
C4348 VDD.n4047 GND 0.005326f
C4349 VDD.n4048 GND 0.004287f
C4350 VDD.n4049 GND 0.005326f
C4351 VDD.n4050 GND 0.493757f
C4352 VDD.n4051 GND 0.005326f
C4353 VDD.n4052 GND 0.004287f
C4354 VDD.n4053 GND 0.005326f
C4355 VDD.n4054 GND 0.005326f
C4356 VDD.n4055 GND 0.005326f
C4357 VDD.n4056 GND 0.004287f
C4358 VDD.n4057 GND 0.005326f
C4359 VDD.n4058 GND 0.58089f
C4360 VDD.n4059 GND 0.005326f
C4361 VDD.n4060 GND 0.004287f
C4362 VDD.n4061 GND 0.005326f
C4363 VDD.n4062 GND 0.005326f
C4364 VDD.n4063 GND 0.005326f
C4365 VDD.n4064 GND 0.004287f
C4366 VDD.n4065 GND 0.005326f
C4367 VDD.n4066 GND 0.58089f
C4368 VDD.n4067 GND 0.005326f
C4369 VDD.n4068 GND 0.004287f
C4370 VDD.n4069 GND 0.005326f
C4371 VDD.n4070 GND 0.005326f
C4372 VDD.n4071 GND 0.005326f
C4373 VDD.n4072 GND 0.004287f
C4374 VDD.n4073 GND 0.005326f
C4375 VDD.n4074 GND 0.58089f
C4376 VDD.n4075 GND 0.005326f
C4377 VDD.n4076 GND 0.004287f
C4378 VDD.n4077 GND 0.005326f
C4379 VDD.n4078 GND 0.005326f
C4380 VDD.n4079 GND 0.005326f
C4381 VDD.n4080 GND 0.004287f
C4382 VDD.n4081 GND 0.005326f
C4383 VDD.n4082 GND 0.58089f
C4384 VDD.n4083 GND 0.005326f
C4385 VDD.n4084 GND 0.004287f
C4386 VDD.n4085 GND 0.005326f
C4387 VDD.n4086 GND 0.005326f
C4388 VDD.n4087 GND 0.005326f
C4389 VDD.n4088 GND 0.005326f
C4390 VDD.n4089 GND 0.005326f
C4391 VDD.n4090 GND 0.004287f
C4392 VDD.n4091 GND 0.005326f
C4393 VDD.n4092 GND 0.58089f
C4394 VDD.n4093 GND 0.005326f
C4395 VDD.n4094 GND 0.005326f
C4396 VDD.n4095 GND 0.005326f
C4397 VDD.n4096 GND 0.005326f
C4398 VDD.n4097 GND 0.004287f
C4399 VDD.n4098 GND 0.005326f
C4400 VDD.n4099 GND 0.005326f
C4401 VDD.n4100 GND 0.005326f
C4402 VDD.n4101 GND 0.005326f
C4403 VDD.n4102 GND 0.58089f
C4404 VDD.n4103 GND 0.005326f
C4405 VDD.n4104 GND 0.005326f
C4406 VDD.n4105 GND 0.005326f
C4407 VDD.n4106 GND 0.005326f
C4408 VDD.n4107 GND 0.005326f
C4409 VDD.n4108 GND 0.004287f
C4410 VDD.n4109 GND 0.005326f
C4411 VDD.n4110 GND 0.005326f
C4412 VDD.n4111 GND 0.005326f
C4413 VDD.n4112 GND 0.005326f
C4414 VDD.t9 GND 0.290445f
C4415 VDD.n4113 GND 0.005326f
C4416 VDD.n4114 GND 0.005326f
C4417 VDD.n4115 GND 0.005326f
C4418 VDD.n4116 GND 0.005326f
C4419 VDD.n4117 GND 0.005326f
C4420 VDD.n4118 GND 0.004287f
C4421 VDD.n4119 GND 0.005326f
C4422 VDD.n4120 GND 0.377579f
C4423 VDD.n4121 GND 0.005326f
C4424 VDD.n4122 GND 0.005326f
C4425 VDD.n4123 GND 0.005326f
C4426 VDD.n4124 GND 0.58089f
C4427 VDD.n4125 GND 0.005326f
C4428 VDD.n4126 GND 0.005326f
C4429 VDD.n4127 GND 0.005326f
C4430 VDD.n4128 GND 0.005326f
C4431 VDD.n4129 GND 0.005326f
C4432 VDD.n4130 GND 0.004287f
C4433 VDD.n4131 GND 0.005326f
C4434 VDD.n4132 GND 0.005326f
C4435 VDD.n4133 GND 0.005326f
C4436 VDD.n4134 GND 0.005326f
C4437 VDD.n4135 GND 0.58089f
C4438 VDD.n4136 GND 0.005326f
C4439 VDD.n4137 GND 0.005326f
C4440 VDD.n4138 GND 0.005326f
C4441 VDD.n4139 GND 0.005326f
C4442 VDD.n4140 GND 0.005326f
C4443 VDD.n4141 GND 0.004287f
C4444 VDD.n4142 GND 0.005326f
C4445 VDD.n4143 GND 0.005326f
C4446 VDD.n4144 GND 0.005326f
C4447 VDD.n4145 GND 0.005326f
C4448 VDD.n4146 GND 0.58089f
C4449 VDD.n4147 GND 0.005326f
C4450 VDD.n4148 GND 0.005326f
C4451 VDD.n4149 GND 0.005326f
C4452 VDD.n4150 GND 0.005326f
C4453 VDD.n4151 GND 0.005326f
C4454 VDD.n4152 GND 0.004287f
C4455 VDD.n4153 GND 0.005326f
C4456 VDD.n4154 GND 0.005326f
C4457 VDD.n4155 GND 0.005326f
C4458 VDD.n4156 GND 0.005326f
C4459 VDD.n4157 GND 0.58089f
C4460 VDD.n4158 GND 0.005326f
C4461 VDD.n4159 GND 0.005326f
C4462 VDD.n4160 GND 0.005326f
C4463 VDD.n4161 GND 0.005326f
C4464 VDD.n4162 GND 0.005326f
C4465 VDD.n4163 GND 0.004287f
C4466 VDD.n4164 GND 0.005326f
C4467 VDD.n4165 GND 0.005326f
C4468 VDD.n4166 GND 0.005326f
C4469 VDD.n4167 GND 0.012264f
C4470 VDD.n4168 GND 1.34186f
C4471 VDD.n4169 GND 0.012553f
C4472 VDD.n4170 GND 0.005326f
C4473 VDD.n4171 GND 0.005326f
C4474 VDD.n4173 GND 0.005326f
C4475 VDD.n4174 GND 0.005326f
C4476 VDD.n4175 GND 0.004287f
C4477 VDD.n4176 GND 0.004287f
C4478 VDD.n4177 GND 0.005326f
C4479 VDD.n4178 GND 0.005326f
C4480 VDD.n4179 GND 0.005326f
C4481 VDD.n4180 GND 0.005326f
C4482 VDD.n4181 GND 0.005326f
C4483 VDD.n4182 GND 0.005326f
C4484 VDD.n4183 GND 0.004287f
C4485 VDD.n4185 GND 0.005326f
C4486 VDD.n4186 GND 0.005326f
C4487 VDD.n4187 GND 0.005326f
C4488 VDD.n4188 GND 0.005326f
C4489 VDD.n4189 GND 0.005326f
C4490 VDD.n4190 GND 0.004287f
C4491 VDD.n4192 GND 0.005326f
C4492 VDD.n4193 GND 0.005326f
C4493 VDD.n4194 GND 0.005326f
C4494 VDD.n4195 GND 0.005326f
C4495 VDD.n4196 GND 0.005326f
C4496 VDD.n4197 GND 0.004287f
C4497 VDD.n4199 GND 0.005326f
C4498 VDD.n4200 GND 0.005326f
C4499 VDD.n4201 GND 0.005326f
C4500 VDD.n4202 GND 0.005326f
C4501 VDD.n4203 GND 0.005326f
C4502 VDD.n4204 GND 0.004287f
C4503 VDD.n4206 GND 0.005326f
C4504 VDD.n4207 GND 0.005326f
C4505 VDD.n4208 GND 0.005326f
C4506 VDD.n4209 GND 0.005326f
C4507 VDD.n4210 GND 0.005326f
C4508 VDD.n4211 GND 0.004287f
C4509 VDD.n4213 GND 0.005326f
C4510 VDD.n4214 GND 0.005326f
C4511 VDD.n4215 GND 0.005326f
C4512 VDD.n4216 GND 0.005326f
C4513 VDD.n4217 GND 0.005326f
C4514 VDD.n4218 GND 0.004287f
C4515 VDD.n4220 GND 0.005326f
C4516 VDD.n4221 GND 0.005326f
C4517 VDD.n4222 GND 0.005326f
C4518 VDD.n4223 GND 0.005326f
C4519 VDD.n4224 GND 0.005326f
C4520 VDD.t107 GND 0.159105f
C4521 VDD.t106 GND 0.597454f
C4522 VDD.n4225 GND 0.084294f
C4523 VDD.t108 GND 0.119732f
C4524 VDD.n4226 GND 0.085079f
C4525 VDD.n4227 GND 0.005894f
C4526 VDD.n4229 GND 0.002808f
C4527 VDD.n4230 GND 0.005326f
C4528 VDD.n4231 GND 0.005326f
C4529 VDD.n4232 GND 0.005326f
C4530 VDD.n4233 GND 0.005326f
C4531 VDD.n4234 GND 0.005326f
C4532 VDD.n4235 GND 0.004287f
C4533 VDD.n4237 GND 0.005326f
C4534 VDD.n4238 GND 0.005326f
C4535 VDD.n4239 GND 0.005326f
C4536 VDD.n4240 GND 0.005326f
C4537 VDD.n4241 GND 0.005326f
C4538 VDD.n4242 GND 0.004287f
C4539 VDD.n4244 GND 0.005326f
C4540 VDD.n4245 GND 0.005326f
C4541 VDD.n4246 GND 0.005326f
C4542 VDD.n4247 GND 0.005326f
C4543 VDD.n4248 GND 0.005326f
C4544 VDD.n4249 GND 0.004287f
C4545 VDD.n4251 GND 0.005326f
C4546 VDD.n4252 GND 0.005326f
C4547 VDD.n4253 GND 0.005326f
C4548 VDD.n4254 GND 0.005326f
C4549 VDD.n4255 GND 0.005326f
C4550 VDD.t92 GND 0.159105f
C4551 VDD.t91 GND 0.597454f
C4552 VDD.n4256 GND 0.084294f
C4553 VDD.t93 GND 0.119732f
C4554 VDD.n4257 GND 0.085079f
C4555 VDD.n4258 GND 0.008037f
C4556 VDD.n4260 GND 0.005326f
C4557 VDD.n4261 GND 0.004287f
C4558 VDD.n4262 GND 0.005326f
C4559 VDD.n4263 GND 0.005326f
C4560 VDD.n4264 GND 0.004287f
C4561 VDD.n4266 GND 0.005326f
C4562 VDD.n4267 GND 0.005326f
C4563 VDD.n4268 GND 0.005326f
C4564 VDD.n4269 GND 0.005326f
C4565 VDD.n4270 GND 0.004287f
C4566 VDD.n4272 GND 0.005326f
C4567 VDD.n4273 GND 0.005326f
C4568 VDD.n4274 GND 0.005326f
C4569 VDD.n4275 GND 0.005326f
C4570 VDD.n4276 GND 0.005326f
C4571 VDD.n4277 GND 0.004287f
C4572 VDD.n4279 GND 0.005326f
C4573 VDD.n4280 GND 0.005326f
C4574 VDD.n4281 GND 0.005326f
C4575 VDD.n4282 GND 0.005326f
C4576 VDD.n4283 GND 0.005326f
C4577 VDD.n4284 GND 0.004222f
C4578 VDD.n4286 GND 0.005326f
C4579 VDD.n4287 GND 0.002936f
C4580 VDD.t104 GND 0.159105f
C4581 VDD.t103 GND 0.597454f
C4582 VDD.n4288 GND 0.084294f
C4583 VDD.t105 GND 0.119732f
C4584 VDD.n4289 GND 0.085079f
C4585 VDD.n4290 GND 0.005326f
C4586 VDD.n4291 GND 0.005326f
C4587 VDD.n4292 GND 0.004287f
C4588 VDD.n4294 GND 0.005326f
C4589 VDD.n4295 GND 0.005326f
C4590 VDD.n4296 GND 0.005326f
C4591 VDD.n4297 GND 0.005326f
C4592 VDD.n4298 GND 0.004287f
C4593 VDD.n4300 GND 0.005326f
C4594 VDD.n4301 GND 0.005326f
C4595 VDD.n4302 GND 0.005326f
C4596 VDD.n4303 GND 0.005326f
C4597 VDD.n4304 GND 0.005326f
C4598 VDD.n4305 GND 0.004287f
C4599 VDD.n4307 GND 0.005326f
C4600 VDD.n4308 GND 0.005326f
C4601 VDD.n4309 GND 0.005326f
C4602 VDD.n4310 GND 0.005326f
C4603 VDD.n4311 GND 0.005326f
C4604 VDD.n4312 GND 0.004287f
C4605 VDD.n4314 GND 0.005326f
C4606 VDD.n4315 GND 0.005326f
C4607 VDD.n4316 GND 0.005326f
C4608 VDD.n4318 GND 0.012553f
C4609 VDD.n4319 GND 0.002272f
C4610 VDD.t96 GND 0.117451f
C4611 VDD.t95 GND 0.160644f
C4612 VDD.t94 GND 0.597454f
C4613 VDD.n4320 GND 0.084171f
C4614 VDD.n4321 GND 0.084531f
C4615 VDD.n4322 GND 0.005326f
C4616 VDD.n4323 GND 0.005326f
C4617 VDD.n4324 GND 0.004287f
C4618 VDD.n4325 GND 0.005326f
C4619 VDD.n4326 GND 0.005326f
C4620 VDD.n4327 GND 0.004287f
C4621 VDD.n4328 GND 0.005326f
C4622 VDD.n4329 GND 0.005326f
C4623 VDD.n4330 GND 0.004287f
C4624 VDD.n4331 GND 0.005326f
C4625 VDD.n4332 GND 0.005326f
C4626 VDD.n4333 GND 0.004287f
C4627 VDD.n4334 GND 0.005326f
C4628 VDD.n4335 GND 0.005326f
C4629 VDD.n4336 GND 0.004287f
C4630 VDD.n4337 GND 0.005326f
C4631 VDD.n4338 GND 0.005326f
C4632 VDD.n4339 GND 0.004287f
C4633 VDD.n4340 GND 0.005326f
C4634 VDD.n4341 GND 0.005326f
C4635 VDD.n4342 GND 0.005326f
C4636 VDD.n4343 GND 0.004287f
C4637 VDD.n4344 GND 0.004287f
C4638 VDD.n4345 GND 0.004287f
C4639 VDD.n4346 GND 0.005326f
C4640 VDD.n4347 GND 0.005326f
C4641 VDD.n4348 GND 0.005326f
C4642 VDD.n4349 GND 0.004287f
C4643 VDD.n4350 GND 0.004287f
C4644 VDD.n4351 GND 0.004287f
C4645 VDD.n4352 GND 0.005326f
C4646 VDD.n4353 GND 0.005326f
C4647 VDD.n4354 GND 0.005326f
C4648 VDD.n4355 GND 0.004287f
C4649 VDD.n4356 GND 0.004287f
C4650 VDD.n4357 GND 0.004287f
C4651 VDD.n4358 GND 0.005326f
C4652 VDD.n4359 GND 0.005326f
C4653 VDD.n4360 GND 0.005326f
C4654 VDD.n4361 GND 0.004287f
C4655 VDD.n4362 GND 0.004287f
C4656 VDD.n4363 GND 0.004287f
C4657 VDD.n4364 GND 0.005326f
C4658 VDD.n4365 GND 0.005326f
C4659 VDD.n4366 GND 0.005326f
C4660 VDD.n4367 GND 0.004287f
C4661 VDD.n4368 GND 0.004287f
C4662 VDD.n4369 GND 0.004287f
C4663 VDD.n4370 GND 0.005326f
C4664 VDD.n4371 GND 0.005326f
C4665 VDD.n4372 GND 0.005326f
C4666 VDD.n4373 GND 0.004287f
C4667 VDD.n4374 GND 0.004287f
C4668 VDD.n4375 GND 0.004287f
C4669 VDD.n4376 GND 0.005326f
C4670 VDD.n4377 GND 0.005326f
C4671 VDD.n4378 GND 0.005326f
C4672 VDD.n4379 GND 0.004287f
C4673 VDD.n4380 GND 0.004287f
C4674 VDD.n4381 GND 0.003558f
C4675 VDD.n4382 GND 0.012264f
C4676 VDD.n4383 GND 0.012553f
C4677 VDD.n4384 GND 0.005326f
C4678 VDD.n4385 GND 0.009452f
C4679 VDD.n4386 GND 0.004158f
C4680 VDD.n4387 GND 0.005326f
C4681 VDD.n4389 GND 0.005326f
C4682 VDD.n4390 GND 0.005326f
C4683 VDD.n4391 GND 0.004287f
C4684 VDD.n4392 GND 0.004287f
C4685 VDD.n4393 GND 0.004287f
C4686 VDD.n4394 GND 0.005326f
C4687 VDD.n4396 GND 0.005326f
C4688 VDD.n4397 GND 0.005326f
C4689 VDD.n4398 GND 0.004287f
C4690 VDD.n4399 GND 0.004287f
C4691 VDD.n4400 GND 0.004287f
C4692 VDD.n4401 GND 0.005326f
C4693 VDD.n4403 GND 0.005326f
C4694 VDD.n4404 GND 0.005326f
C4695 VDD.n4405 GND 0.004287f
C4696 VDD.n4406 GND 0.004287f
C4697 VDD.n4407 GND 0.004287f
C4698 VDD.n4408 GND 0.005326f
C4699 VDD.n4410 GND 0.005326f
C4700 VDD.n4411 GND 0.005326f
C4701 VDD.n4412 GND 0.004287f
C4702 VDD.n4413 GND 0.005326f
C4703 VDD.n4414 GND 0.005326f
C4704 VDD.n4415 GND 0.005326f
C4705 VDD.n4416 GND 0.008037f
C4706 VDD.n4417 GND 0.005326f
C4707 VDD.n4419 GND 0.005326f
C4708 VDD.n4420 GND 0.005326f
C4709 VDD.n4421 GND 0.004287f
C4710 VDD.n4422 GND 0.004287f
C4711 VDD.n4423 GND 0.004287f
C4712 VDD.n4424 GND 0.005326f
C4713 VDD.n4426 GND 0.005326f
C4714 VDD.n4427 GND 0.005326f
C4715 VDD.n4428 GND 0.004287f
C4716 VDD.n4429 GND 0.004287f
C4717 VDD.n4430 GND 0.004287f
C4718 VDD.n4431 GND 0.005326f
C4719 VDD.n4433 GND 0.005326f
C4720 VDD.n4434 GND 0.005326f
C4721 VDD.n4435 GND 0.004287f
C4722 VDD.n4436 GND 0.004287f
C4723 VDD.n4437 GND 0.004287f
C4724 VDD.n4438 GND 0.005326f
C4725 VDD.n4440 GND 0.005326f
C4726 VDD.n4441 GND 0.005326f
C4727 VDD.n4442 GND 0.004287f
C4728 VDD.n4443 GND 0.005326f
C4729 VDD.n4444 GND 0.005326f
C4730 VDD.n4445 GND 0.005326f
C4731 VDD.n4446 GND 0.002872f
C4732 VDD.n4447 GND 0.005326f
C4733 VDD.n4449 GND 0.005326f
C4734 VDD.n4450 GND 0.005326f
C4735 VDD.n4451 GND 0.004287f
C4736 VDD.n4452 GND 0.004287f
C4737 VDD.n4453 GND 0.004287f
C4738 VDD.n4454 GND 0.005326f
C4739 VDD.n4456 GND 0.005326f
C4740 VDD.n4457 GND 0.005326f
C4741 VDD.n4458 GND 0.004287f
C4742 VDD.n4459 GND 0.004287f
C4743 VDD.n4460 GND 0.004287f
C4744 VDD.n4461 GND 0.005326f
C4745 VDD.n4463 GND 0.005326f
C4746 VDD.n4464 GND 0.005326f
C4747 VDD.n4465 GND 0.004287f
C4748 VDD.n4466 GND 0.004287f
C4749 VDD.n4467 GND 0.004287f
C4750 VDD.n4468 GND 0.005326f
C4751 VDD.n4470 GND 0.005326f
C4752 VDD.n4471 GND 0.005326f
C4753 VDD.n4472 GND 0.004287f
C4754 VDD.n4473 GND 0.004287f
C4755 VDD.n4474 GND 0.004287f
C4756 VDD.n4475 GND 0.005326f
C4757 VDD.n4477 GND 0.005326f
C4758 VDD.n4478 GND 0.005326f
C4759 VDD.n4479 GND 0.002208f
C4760 VDD.n4480 GND 0.004287f
C4761 VDD.n4481 GND 0.004287f
C4762 VDD.n4482 GND 0.005326f
C4763 VDD.n4484 GND 0.005326f
C4764 VDD.n4485 GND 0.005326f
C4765 VDD.n4486 GND 0.004287f
C4766 VDD.n4487 GND 0.004287f
C4767 VDD.n4488 GND 0.004287f
C4768 VDD.n4489 GND 0.005326f
C4769 VDD.n4491 GND 0.005326f
C4770 VDD.n4492 GND 0.005326f
C4771 VDD.n4493 GND 0.004287f
C4772 VDD.n4494 GND 0.004287f
C4773 VDD.n4495 GND 0.004287f
C4774 VDD.n4496 GND 0.005326f
C4775 VDD.n4498 GND 0.005326f
C4776 VDD.n4499 GND 0.005326f
C4777 VDD.n4500 GND 0.004287f
C4778 VDD.n4501 GND 0.004287f
C4779 VDD.n4502 GND 0.004287f
C4780 VDD.n4503 GND 0.005326f
C4781 VDD.n4505 GND 0.005326f
C4782 VDD.n4506 GND 0.005326f
C4783 VDD.n4507 GND 0.002743f
C4784 VDD.t39 GND 0.159105f
C4785 VDD.t37 GND 0.597454f
C4786 VDD.n4508 GND 0.084294f
C4787 VDD.t40 GND 0.119732f
C4788 VDD.n4509 GND 0.085079f
C4789 VDD.n4510 GND 0.005894f
C4790 VDD.n4511 GND 0.002272f
C4791 VDD.n4512 GND 0.004287f
C4792 VDD.n4513 GND 0.005326f
C4793 VDD.n4515 GND 0.005326f
C4794 VDD.n4516 GND 0.005326f
C4795 VDD.n4517 GND 0.004287f
C4796 VDD.n4518 GND 0.004287f
C4797 VDD.n4519 GND 0.004287f
C4798 VDD.n4520 GND 0.005326f
C4799 VDD.n4522 GND 0.005326f
C4800 VDD.n4523 GND 0.005326f
C4801 VDD.n4524 GND 0.004287f
C4802 VDD.n4525 GND 0.004287f
C4803 VDD.n4526 GND 0.004287f
C4804 VDD.n4527 GND 0.005326f
C4805 VDD.n4529 GND 0.005326f
C4806 VDD.n4530 GND 0.005326f
C4807 VDD.n4532 GND 0.005326f
C4808 VDD.n4533 GND 0.004287f
C4809 VDD.n4534 GND 0.004287f
C4810 VDD.n4535 GND 0.003558f
C4811 VDD.n4536 GND 0.012553f
C4812 VDD.n4537 GND 0.012264f
C4813 VDD.n4538 GND 0.003558f
C4814 VDD.n4539 GND 0.012264f
C4815 VDD.n4540 GND 0.824864f
C4816 VDD.n4541 GND 0.58089f
C4817 VDD.n4542 GND 0.58089f
C4818 VDD.n4543 GND 0.005326f
C4819 VDD.n4544 GND 0.004287f
C4820 VDD.n4545 GND 0.004287f
C4821 VDD.n4546 GND 0.004287f
C4822 VDD.n4547 GND 0.005326f
C4823 VDD.n4548 GND 0.58089f
C4824 VDD.n4549 GND 0.511183f
C4825 VDD.t38 GND 0.290445f
C4826 VDD.n4550 GND 0.360152f
C4827 VDD.n4551 GND 0.005326f
C4828 VDD.n4552 GND 0.004287f
C4829 VDD.n4553 GND 0.004287f
C4830 VDD.n4554 GND 0.004287f
C4831 VDD.n4555 GND 0.005326f
C4832 VDD.n4556 GND 0.58089f
C4833 VDD.n4557 GND 0.58089f
C4834 VDD.n4558 GND 0.58089f
C4835 VDD.n4559 GND 0.005326f
C4836 VDD.n4560 GND 0.004287f
C4837 VDD.n4561 GND 0.004287f
C4838 VDD.n4562 GND 0.004287f
C4839 VDD.n4563 GND 0.005326f
C4840 VDD.n4564 GND 0.58089f
C4841 VDD.n4565 GND 0.58089f
C4842 VDD.n4566 GND 0.58089f
C4843 VDD.n4567 GND 0.005326f
C4844 VDD.n4568 GND 0.004287f
C4845 VDD.n4569 GND 0.004287f
C4846 VDD.n4570 GND 0.004287f
C4847 VDD.n4571 GND 0.005326f
C4848 VDD.n4572 GND 0.58089f
C4849 VDD.n4573 GND 0.58089f
C4850 VDD.n4574 GND 0.58089f
C4851 VDD.n4575 GND 0.005326f
C4852 VDD.n4576 GND 0.004287f
C4853 VDD.n4577 GND 0.004287f
C4854 VDD.n4578 GND 0.004287f
C4855 VDD.n4579 GND 0.005326f
C4856 VDD.n4580 GND 0.493757f
C4857 VDD.n4581 GND 0.58089f
C4858 VDD.n4582 GND 0.58089f
C4859 VDD.n4583 GND 0.005326f
C4860 VDD.n4584 GND 0.004287f
C4861 VDD.n4585 GND 0.004287f
C4862 VDD.n4586 GND 0.004287f
C4863 VDD.n4587 GND 0.005326f
C4864 VDD.n4588 GND 0.58089f
C4865 VDD.n4589 GND 0.58089f
C4866 VDD.n4590 GND 0.58089f
C4867 VDD.n4591 GND 0.005326f
C4868 VDD.n4592 GND 0.004287f
C4869 VDD.n4593 GND 0.004287f
C4870 VDD.n4594 GND 0.004287f
C4871 VDD.n4595 GND 0.005326f
C4872 VDD.n4596 GND 0.58089f
C4873 VDD.n4597 GND 0.005326f
C4874 VDD.n4598 GND 0.004287f
C4875 VDD.n4599 GND 0.004287f
C4876 VDD.n4600 GND 0.004287f
C4877 VDD.n4601 GND 0.005326f
C4878 VDD.t6 GND 0.58089f
C4879 VDD.n4602 GND 0.005326f
C4880 VDD.n4603 GND 0.004287f
C4881 VDD.n4604 GND 0.118204f
C4882 VDD.n4605 GND 2.0753f
C4883 a_n10827_11007.n0 GND 7.81229f
C4884 a_n10827_11007.n1 GND 5.51957f
C4885 a_n10827_11007.t8 GND 0.095784f
C4886 a_n10827_11007.t4 GND 0.095784f
C4887 a_n10827_11007.t3 GND 0.095784f
C4888 a_n10827_11007.n2 GND 0.471602f
C4889 a_n10827_11007.t5 GND 0.095784f
C4890 a_n10827_11007.t9 GND 0.095784f
C4891 a_n10827_11007.n3 GND 0.468109f
C4892 a_n10827_11007.t7 GND 0.095784f
C4893 a_n10827_11007.t6 GND 0.095784f
C4894 a_n10827_11007.n4 GND 0.438976f
C4895 a_n10827_11007.n5 GND 19.267302f
C4896 a_n10827_11007.t1 GND 0.520609f
C4897 a_n10827_11007.t2 GND 0.095784f
C4898 a_n10827_11007.t13 GND 0.095784f
C4899 a_n10827_11007.n6 GND 0.352656f
C4900 a_n10827_11007.t0 GND 0.50087f
C4901 a_n10827_11007.t14 GND 0.50087f
C4902 a_n10827_11007.t12 GND 0.095784f
C4903 a_n10827_11007.t15 GND 0.095784f
C4904 a_n10827_11007.n7 GND 0.352656f
C4905 a_n10827_11007.t11 GND 0.50087f
C4906 a_n10827_11007.n8 GND 6.29434f
C4907 a_n10827_11007.n9 GND 9.110929f
C4908 a_n10827_11007.n10 GND 0.438976f
C4909 a_n10827_11007.t10 GND 0.095784f
C4910 a_n10683_10810.t39 GND 2.34869f
C4911 a_n10683_10810.t36 GND 2.05497f
C4912 a_n10683_10810.n0 GND 4.11996f
C4913 a_n10683_10810.n1 GND 20.598f
C4914 a_n10683_10810.t41 GND 2.08053f
C4915 a_n10683_10810.n3 GND 12.0365f
C4916 a_n10683_10810.n4 GND 0.892299f
C4917 a_n10683_10810.t27 GND 2.35023f
C4918 a_n10683_10810.t30 GND 2.05459f
C4919 a_n10683_10810.n5 GND 0.654624f
C4920 a_n10683_10810.t26 GND 2.07072f
C4921 a_n10683_10810.t20 GND 2.06176f
C4922 a_n10683_10810.t37 GND 2.07072f
C4923 a_n10683_10810.t40 GND 2.06176f
C4924 a_n10683_10810.t31 GND 2.09237f
C4925 a_n10683_10810.t34 GND 2.0507f
C4926 a_n10683_10810.t28 GND 2.09237f
C4927 a_n10683_10810.t24 GND 2.0507f
C4928 a_n10683_10810.t38 GND 2.08053f
C4929 a_n10683_10810.t42 GND 2.08053f
C4930 a_n10683_10810.t33 GND 2.31839f
C4931 a_n10683_10810.t12 GND 2.05916f
C4932 a_n10683_10810.n6 GND 4.25616f
C4933 a_n10683_10810.n7 GND 0.691856f
C4934 a_n10683_10810.t35 GND 2.05916f
C4935 a_n10683_10810.n8 GND 0.691856f
C4936 a_n10683_10810.t23 GND 2.31839f
C4937 a_n10683_10810.t22 GND 2.31839f
C4938 a_n10683_10810.t16 GND 2.05224f
C4939 a_n10683_10810.t10 GND 2.07628f
C4940 a_n10683_10810.n9 GND 0.425763f
C4941 a_n10683_10810.n10 GND 0.425763f
C4942 a_n10683_10810.n11 GND 6.62334f
C4943 a_n10683_10810.n12 GND 6.76462f
C4944 a_n10683_10810.n13 GND 2.57188f
C4945 a_n10683_10810.t9 GND 0.067488f
C4946 a_n10683_10810.t13 GND 0.366812f
C4947 a_n10683_10810.t6 GND 2.33455f
C4948 a_n10683_10810.t25 GND 2.33455f
C4949 a_n10683_10810.t14 GND 2.36549f
C4950 a_n10683_10810.t18 GND 2.05316f
C4951 a_n10683_10810.t21 GND 2.12898f
C4952 a_n10683_10810.t43 GND 2.05093f
C4953 a_n10683_10810.t2 GND 1.44433f
C4954 a_n10683_10810.t0 GND 0.052877f
C4955 a_n10683_10810.t1 GND 0.375484f
C4956 a_n10683_10810.t3 GND 0.052877f
C4957 a_n10683_10810.n14 GND 10.284201f
C4958 a_n10683_10810.t11 GND 0.366812f
C4959 a_n10683_10810.t19 GND 0.067488f
C4960 a_n10683_10810.t17 GND 0.067488f
C4961 a_n10683_10810.n15 GND 0.248475f
C4962 a_n10683_10810.t15 GND 0.352904f
C4963 a_n10683_10810.t32 GND 2.05511f
C4964 a_n10683_10810.t29 GND 1.4369f
C4965 a_n10683_10810.n16 GND 0.88835f
C4966 a_n10683_10810.t8 GND 2.05511f
C4967 a_n10683_10810.t4 GND 1.4369f
C4968 a_n10683_10810.n17 GND 0.88835f
C4969 a_n10683_10810.t7 GND 0.352904f
C4970 a_n10683_10810.n18 GND 0.248476f
C4971 a_n10683_10810.t5 GND 0.067488f
.ends

