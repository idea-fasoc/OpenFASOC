* NGSPICE file created from diff_pair_sample_0388.ext - technology: sky130A

.subckt diff_pair_sample_0388 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t15 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X1 B.t11 B.t9 B.t10 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=0 ps=0 w=13.37 l=2.63
X2 VDD1.t7 VP.t0 VTAIL.t1 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X3 VDD2.t6 VN.t1 VTAIL.t14 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X4 VTAIL.t13 VN.t2 VDD2.t5 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X5 VDD1.t6 VP.t1 VTAIL.t4 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=5.2143 ps=27.52 w=13.37 l=2.63
X6 VTAIL.t3 VP.t2 VDD1.t5 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=2.20605 ps=13.7 w=13.37 l=2.63
X7 VDD1.t4 VP.t3 VTAIL.t2 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X8 B.t8 B.t6 B.t7 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=0 ps=0 w=13.37 l=2.63
X9 VDD2.t4 VN.t3 VTAIL.t8 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=5.2143 ps=27.52 w=13.37 l=2.63
X10 VDD1.t3 VP.t4 VTAIL.t6 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=5.2143 ps=27.52 w=13.37 l=2.63
X11 VTAIL.t7 VP.t5 VDD1.t2 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X12 VTAIL.t5 VP.t6 VDD1.t1 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=2.20605 ps=13.7 w=13.37 l=2.63
X13 B.t5 B.t3 B.t4 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=0 ps=0 w=13.37 l=2.63
X14 B.t2 B.t0 B.t1 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=0 ps=0 w=13.37 l=2.63
X15 VDD2.t3 VN.t4 VTAIL.t9 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=5.2143 ps=27.52 w=13.37 l=2.63
X16 VTAIL.t10 VN.t5 VDD2.t2 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X17 VTAIL.t0 VP.t7 VDD1.t0 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=2.20605 pd=13.7 as=2.20605 ps=13.7 w=13.37 l=2.63
X18 VTAIL.t11 VN.t6 VDD2.t1 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=2.20605 ps=13.7 w=13.37 l=2.63
X19 VTAIL.t12 VN.t7 VDD2.t0 w_n3930_n3642# sky130_fd_pr__pfet_01v8 ad=5.2143 pd=27.52 as=2.20605 ps=13.7 w=13.37 l=2.63
R0 VN.n55 VN.n29 161.3
R1 VN.n54 VN.n53 161.3
R2 VN.n52 VN.n30 161.3
R3 VN.n51 VN.n50 161.3
R4 VN.n49 VN.n31 161.3
R5 VN.n48 VN.n47 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n26 VN.n0 161.3
R13 VN.n25 VN.n24 161.3
R14 VN.n23 VN.n1 161.3
R15 VN.n22 VN.n21 161.3
R16 VN.n20 VN.n2 161.3
R17 VN.n19 VN.n18 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n7 VN.t6 155.923
R25 VN.n36 VN.t3 155.923
R26 VN.n8 VN.t0 122.516
R27 VN.n3 VN.t5 122.516
R28 VN.n27 VN.t4 122.516
R29 VN.n37 VN.t2 122.516
R30 VN.n32 VN.t1 122.516
R31 VN.n56 VN.t7 122.516
R32 VN.n28 VN.n27 101.459
R33 VN.n57 VN.n56 101.459
R34 VN.n8 VN.n7 61.154
R35 VN.n37 VN.n36 61.154
R36 VN.n14 VN.n5 56.5193
R37 VN.n21 VN.n1 56.5193
R38 VN.n43 VN.n34 56.5193
R39 VN.n50 VN.n30 56.5193
R40 VN VN.n57 52.3694
R41 VN.n10 VN.n9 24.4675
R42 VN.n10 VN.n5 24.4675
R43 VN.n15 VN.n14 24.4675
R44 VN.n16 VN.n15 24.4675
R45 VN.n20 VN.n19 24.4675
R46 VN.n21 VN.n20 24.4675
R47 VN.n25 VN.n1 24.4675
R48 VN.n26 VN.n25 24.4675
R49 VN.n39 VN.n34 24.4675
R50 VN.n39 VN.n38 24.4675
R51 VN.n50 VN.n49 24.4675
R52 VN.n49 VN.n48 24.4675
R53 VN.n45 VN.n44 24.4675
R54 VN.n44 VN.n43 24.4675
R55 VN.n55 VN.n54 24.4675
R56 VN.n54 VN.n30 24.4675
R57 VN.n19 VN.n3 13.2127
R58 VN.n48 VN.n32 13.2127
R59 VN.n9 VN.n8 11.2553
R60 VN.n16 VN.n3 11.2553
R61 VN.n38 VN.n37 11.2553
R62 VN.n45 VN.n32 11.2553
R63 VN.n27 VN.n26 9.29796
R64 VN.n56 VN.n55 9.29796
R65 VN.n36 VN.n35 6.89416
R66 VN.n7 VN.n6 6.89416
R67 VN.n57 VN.n29 0.278367
R68 VN.n28 VN.n0 0.278367
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153454
R92 VTAIL.n537 VTAIL.n536 585
R93 VTAIL.n539 VTAIL.n538 585
R94 VTAIL.n532 VTAIL.n531 585
R95 VTAIL.n545 VTAIL.n544 585
R96 VTAIL.n547 VTAIL.n546 585
R97 VTAIL.n528 VTAIL.n527 585
R98 VTAIL.n553 VTAIL.n552 585
R99 VTAIL.n555 VTAIL.n554 585
R100 VTAIL.n524 VTAIL.n523 585
R101 VTAIL.n561 VTAIL.n560 585
R102 VTAIL.n563 VTAIL.n562 585
R103 VTAIL.n520 VTAIL.n519 585
R104 VTAIL.n569 VTAIL.n568 585
R105 VTAIL.n571 VTAIL.n570 585
R106 VTAIL.n516 VTAIL.n515 585
R107 VTAIL.n577 VTAIL.n576 585
R108 VTAIL.n579 VTAIL.n578 585
R109 VTAIL.n27 VTAIL.n26 585
R110 VTAIL.n29 VTAIL.n28 585
R111 VTAIL.n22 VTAIL.n21 585
R112 VTAIL.n35 VTAIL.n34 585
R113 VTAIL.n37 VTAIL.n36 585
R114 VTAIL.n18 VTAIL.n17 585
R115 VTAIL.n43 VTAIL.n42 585
R116 VTAIL.n45 VTAIL.n44 585
R117 VTAIL.n14 VTAIL.n13 585
R118 VTAIL.n51 VTAIL.n50 585
R119 VTAIL.n53 VTAIL.n52 585
R120 VTAIL.n10 VTAIL.n9 585
R121 VTAIL.n59 VTAIL.n58 585
R122 VTAIL.n61 VTAIL.n60 585
R123 VTAIL.n6 VTAIL.n5 585
R124 VTAIL.n67 VTAIL.n66 585
R125 VTAIL.n69 VTAIL.n68 585
R126 VTAIL.n99 VTAIL.n98 585
R127 VTAIL.n101 VTAIL.n100 585
R128 VTAIL.n94 VTAIL.n93 585
R129 VTAIL.n107 VTAIL.n106 585
R130 VTAIL.n109 VTAIL.n108 585
R131 VTAIL.n90 VTAIL.n89 585
R132 VTAIL.n115 VTAIL.n114 585
R133 VTAIL.n117 VTAIL.n116 585
R134 VTAIL.n86 VTAIL.n85 585
R135 VTAIL.n123 VTAIL.n122 585
R136 VTAIL.n125 VTAIL.n124 585
R137 VTAIL.n82 VTAIL.n81 585
R138 VTAIL.n131 VTAIL.n130 585
R139 VTAIL.n133 VTAIL.n132 585
R140 VTAIL.n78 VTAIL.n77 585
R141 VTAIL.n139 VTAIL.n138 585
R142 VTAIL.n141 VTAIL.n140 585
R143 VTAIL.n173 VTAIL.n172 585
R144 VTAIL.n175 VTAIL.n174 585
R145 VTAIL.n168 VTAIL.n167 585
R146 VTAIL.n181 VTAIL.n180 585
R147 VTAIL.n183 VTAIL.n182 585
R148 VTAIL.n164 VTAIL.n163 585
R149 VTAIL.n189 VTAIL.n188 585
R150 VTAIL.n191 VTAIL.n190 585
R151 VTAIL.n160 VTAIL.n159 585
R152 VTAIL.n197 VTAIL.n196 585
R153 VTAIL.n199 VTAIL.n198 585
R154 VTAIL.n156 VTAIL.n155 585
R155 VTAIL.n205 VTAIL.n204 585
R156 VTAIL.n207 VTAIL.n206 585
R157 VTAIL.n152 VTAIL.n151 585
R158 VTAIL.n213 VTAIL.n212 585
R159 VTAIL.n215 VTAIL.n214 585
R160 VTAIL.n507 VTAIL.n506 585
R161 VTAIL.n505 VTAIL.n504 585
R162 VTAIL.n444 VTAIL.n443 585
R163 VTAIL.n499 VTAIL.n498 585
R164 VTAIL.n497 VTAIL.n496 585
R165 VTAIL.n448 VTAIL.n447 585
R166 VTAIL.n491 VTAIL.n490 585
R167 VTAIL.n489 VTAIL.n488 585
R168 VTAIL.n452 VTAIL.n451 585
R169 VTAIL.n483 VTAIL.n482 585
R170 VTAIL.n481 VTAIL.n480 585
R171 VTAIL.n456 VTAIL.n455 585
R172 VTAIL.n475 VTAIL.n474 585
R173 VTAIL.n473 VTAIL.n472 585
R174 VTAIL.n460 VTAIL.n459 585
R175 VTAIL.n467 VTAIL.n466 585
R176 VTAIL.n465 VTAIL.n464 585
R177 VTAIL.n433 VTAIL.n432 585
R178 VTAIL.n431 VTAIL.n430 585
R179 VTAIL.n370 VTAIL.n369 585
R180 VTAIL.n425 VTAIL.n424 585
R181 VTAIL.n423 VTAIL.n422 585
R182 VTAIL.n374 VTAIL.n373 585
R183 VTAIL.n417 VTAIL.n416 585
R184 VTAIL.n415 VTAIL.n414 585
R185 VTAIL.n378 VTAIL.n377 585
R186 VTAIL.n409 VTAIL.n408 585
R187 VTAIL.n407 VTAIL.n406 585
R188 VTAIL.n382 VTAIL.n381 585
R189 VTAIL.n401 VTAIL.n400 585
R190 VTAIL.n399 VTAIL.n398 585
R191 VTAIL.n386 VTAIL.n385 585
R192 VTAIL.n393 VTAIL.n392 585
R193 VTAIL.n391 VTAIL.n390 585
R194 VTAIL.n361 VTAIL.n360 585
R195 VTAIL.n359 VTAIL.n358 585
R196 VTAIL.n298 VTAIL.n297 585
R197 VTAIL.n353 VTAIL.n352 585
R198 VTAIL.n351 VTAIL.n350 585
R199 VTAIL.n302 VTAIL.n301 585
R200 VTAIL.n345 VTAIL.n344 585
R201 VTAIL.n343 VTAIL.n342 585
R202 VTAIL.n306 VTAIL.n305 585
R203 VTAIL.n337 VTAIL.n336 585
R204 VTAIL.n335 VTAIL.n334 585
R205 VTAIL.n310 VTAIL.n309 585
R206 VTAIL.n329 VTAIL.n328 585
R207 VTAIL.n327 VTAIL.n326 585
R208 VTAIL.n314 VTAIL.n313 585
R209 VTAIL.n321 VTAIL.n320 585
R210 VTAIL.n319 VTAIL.n318 585
R211 VTAIL.n287 VTAIL.n286 585
R212 VTAIL.n285 VTAIL.n284 585
R213 VTAIL.n224 VTAIL.n223 585
R214 VTAIL.n279 VTAIL.n278 585
R215 VTAIL.n277 VTAIL.n276 585
R216 VTAIL.n228 VTAIL.n227 585
R217 VTAIL.n271 VTAIL.n270 585
R218 VTAIL.n269 VTAIL.n268 585
R219 VTAIL.n232 VTAIL.n231 585
R220 VTAIL.n263 VTAIL.n262 585
R221 VTAIL.n261 VTAIL.n260 585
R222 VTAIL.n236 VTAIL.n235 585
R223 VTAIL.n255 VTAIL.n254 585
R224 VTAIL.n253 VTAIL.n252 585
R225 VTAIL.n240 VTAIL.n239 585
R226 VTAIL.n247 VTAIL.n246 585
R227 VTAIL.n245 VTAIL.n244 585
R228 VTAIL.n578 VTAIL.n512 498.474
R229 VTAIL.n68 VTAIL.n2 498.474
R230 VTAIL.n140 VTAIL.n74 498.474
R231 VTAIL.n214 VTAIL.n148 498.474
R232 VTAIL.n506 VTAIL.n440 498.474
R233 VTAIL.n432 VTAIL.n366 498.474
R234 VTAIL.n360 VTAIL.n294 498.474
R235 VTAIL.n286 VTAIL.n220 498.474
R236 VTAIL.n535 VTAIL.t9 327.466
R237 VTAIL.n25 VTAIL.t11 327.466
R238 VTAIL.n97 VTAIL.t4 327.466
R239 VTAIL.n171 VTAIL.t5 327.466
R240 VTAIL.n463 VTAIL.t6 327.466
R241 VTAIL.n389 VTAIL.t3 327.466
R242 VTAIL.n317 VTAIL.t8 327.466
R243 VTAIL.n243 VTAIL.t12 327.466
R244 VTAIL.n538 VTAIL.n537 171.744
R245 VTAIL.n538 VTAIL.n531 171.744
R246 VTAIL.n545 VTAIL.n531 171.744
R247 VTAIL.n546 VTAIL.n545 171.744
R248 VTAIL.n546 VTAIL.n527 171.744
R249 VTAIL.n553 VTAIL.n527 171.744
R250 VTAIL.n554 VTAIL.n553 171.744
R251 VTAIL.n554 VTAIL.n523 171.744
R252 VTAIL.n561 VTAIL.n523 171.744
R253 VTAIL.n562 VTAIL.n561 171.744
R254 VTAIL.n562 VTAIL.n519 171.744
R255 VTAIL.n569 VTAIL.n519 171.744
R256 VTAIL.n570 VTAIL.n569 171.744
R257 VTAIL.n570 VTAIL.n515 171.744
R258 VTAIL.n577 VTAIL.n515 171.744
R259 VTAIL.n578 VTAIL.n577 171.744
R260 VTAIL.n28 VTAIL.n27 171.744
R261 VTAIL.n28 VTAIL.n21 171.744
R262 VTAIL.n35 VTAIL.n21 171.744
R263 VTAIL.n36 VTAIL.n35 171.744
R264 VTAIL.n36 VTAIL.n17 171.744
R265 VTAIL.n43 VTAIL.n17 171.744
R266 VTAIL.n44 VTAIL.n43 171.744
R267 VTAIL.n44 VTAIL.n13 171.744
R268 VTAIL.n51 VTAIL.n13 171.744
R269 VTAIL.n52 VTAIL.n51 171.744
R270 VTAIL.n52 VTAIL.n9 171.744
R271 VTAIL.n59 VTAIL.n9 171.744
R272 VTAIL.n60 VTAIL.n59 171.744
R273 VTAIL.n60 VTAIL.n5 171.744
R274 VTAIL.n67 VTAIL.n5 171.744
R275 VTAIL.n68 VTAIL.n67 171.744
R276 VTAIL.n100 VTAIL.n99 171.744
R277 VTAIL.n100 VTAIL.n93 171.744
R278 VTAIL.n107 VTAIL.n93 171.744
R279 VTAIL.n108 VTAIL.n107 171.744
R280 VTAIL.n108 VTAIL.n89 171.744
R281 VTAIL.n115 VTAIL.n89 171.744
R282 VTAIL.n116 VTAIL.n115 171.744
R283 VTAIL.n116 VTAIL.n85 171.744
R284 VTAIL.n123 VTAIL.n85 171.744
R285 VTAIL.n124 VTAIL.n123 171.744
R286 VTAIL.n124 VTAIL.n81 171.744
R287 VTAIL.n131 VTAIL.n81 171.744
R288 VTAIL.n132 VTAIL.n131 171.744
R289 VTAIL.n132 VTAIL.n77 171.744
R290 VTAIL.n139 VTAIL.n77 171.744
R291 VTAIL.n140 VTAIL.n139 171.744
R292 VTAIL.n174 VTAIL.n173 171.744
R293 VTAIL.n174 VTAIL.n167 171.744
R294 VTAIL.n181 VTAIL.n167 171.744
R295 VTAIL.n182 VTAIL.n181 171.744
R296 VTAIL.n182 VTAIL.n163 171.744
R297 VTAIL.n189 VTAIL.n163 171.744
R298 VTAIL.n190 VTAIL.n189 171.744
R299 VTAIL.n190 VTAIL.n159 171.744
R300 VTAIL.n197 VTAIL.n159 171.744
R301 VTAIL.n198 VTAIL.n197 171.744
R302 VTAIL.n198 VTAIL.n155 171.744
R303 VTAIL.n205 VTAIL.n155 171.744
R304 VTAIL.n206 VTAIL.n205 171.744
R305 VTAIL.n206 VTAIL.n151 171.744
R306 VTAIL.n213 VTAIL.n151 171.744
R307 VTAIL.n214 VTAIL.n213 171.744
R308 VTAIL.n506 VTAIL.n505 171.744
R309 VTAIL.n505 VTAIL.n443 171.744
R310 VTAIL.n498 VTAIL.n443 171.744
R311 VTAIL.n498 VTAIL.n497 171.744
R312 VTAIL.n497 VTAIL.n447 171.744
R313 VTAIL.n490 VTAIL.n447 171.744
R314 VTAIL.n490 VTAIL.n489 171.744
R315 VTAIL.n489 VTAIL.n451 171.744
R316 VTAIL.n482 VTAIL.n451 171.744
R317 VTAIL.n482 VTAIL.n481 171.744
R318 VTAIL.n481 VTAIL.n455 171.744
R319 VTAIL.n474 VTAIL.n455 171.744
R320 VTAIL.n474 VTAIL.n473 171.744
R321 VTAIL.n473 VTAIL.n459 171.744
R322 VTAIL.n466 VTAIL.n459 171.744
R323 VTAIL.n466 VTAIL.n465 171.744
R324 VTAIL.n432 VTAIL.n431 171.744
R325 VTAIL.n431 VTAIL.n369 171.744
R326 VTAIL.n424 VTAIL.n369 171.744
R327 VTAIL.n424 VTAIL.n423 171.744
R328 VTAIL.n423 VTAIL.n373 171.744
R329 VTAIL.n416 VTAIL.n373 171.744
R330 VTAIL.n416 VTAIL.n415 171.744
R331 VTAIL.n415 VTAIL.n377 171.744
R332 VTAIL.n408 VTAIL.n377 171.744
R333 VTAIL.n408 VTAIL.n407 171.744
R334 VTAIL.n407 VTAIL.n381 171.744
R335 VTAIL.n400 VTAIL.n381 171.744
R336 VTAIL.n400 VTAIL.n399 171.744
R337 VTAIL.n399 VTAIL.n385 171.744
R338 VTAIL.n392 VTAIL.n385 171.744
R339 VTAIL.n392 VTAIL.n391 171.744
R340 VTAIL.n360 VTAIL.n359 171.744
R341 VTAIL.n359 VTAIL.n297 171.744
R342 VTAIL.n352 VTAIL.n297 171.744
R343 VTAIL.n352 VTAIL.n351 171.744
R344 VTAIL.n351 VTAIL.n301 171.744
R345 VTAIL.n344 VTAIL.n301 171.744
R346 VTAIL.n344 VTAIL.n343 171.744
R347 VTAIL.n343 VTAIL.n305 171.744
R348 VTAIL.n336 VTAIL.n305 171.744
R349 VTAIL.n336 VTAIL.n335 171.744
R350 VTAIL.n335 VTAIL.n309 171.744
R351 VTAIL.n328 VTAIL.n309 171.744
R352 VTAIL.n328 VTAIL.n327 171.744
R353 VTAIL.n327 VTAIL.n313 171.744
R354 VTAIL.n320 VTAIL.n313 171.744
R355 VTAIL.n320 VTAIL.n319 171.744
R356 VTAIL.n286 VTAIL.n285 171.744
R357 VTAIL.n285 VTAIL.n223 171.744
R358 VTAIL.n278 VTAIL.n223 171.744
R359 VTAIL.n278 VTAIL.n277 171.744
R360 VTAIL.n277 VTAIL.n227 171.744
R361 VTAIL.n270 VTAIL.n227 171.744
R362 VTAIL.n270 VTAIL.n269 171.744
R363 VTAIL.n269 VTAIL.n231 171.744
R364 VTAIL.n262 VTAIL.n231 171.744
R365 VTAIL.n262 VTAIL.n261 171.744
R366 VTAIL.n261 VTAIL.n235 171.744
R367 VTAIL.n254 VTAIL.n235 171.744
R368 VTAIL.n254 VTAIL.n253 171.744
R369 VTAIL.n253 VTAIL.n239 171.744
R370 VTAIL.n246 VTAIL.n239 171.744
R371 VTAIL.n246 VTAIL.n245 171.744
R372 VTAIL.n537 VTAIL.t9 85.8723
R373 VTAIL.n27 VTAIL.t11 85.8723
R374 VTAIL.n99 VTAIL.t4 85.8723
R375 VTAIL.n173 VTAIL.t5 85.8723
R376 VTAIL.n465 VTAIL.t6 85.8723
R377 VTAIL.n391 VTAIL.t3 85.8723
R378 VTAIL.n319 VTAIL.t8 85.8723
R379 VTAIL.n245 VTAIL.t12 85.8723
R380 VTAIL.n439 VTAIL.n438 58.5847
R381 VTAIL.n293 VTAIL.n292 58.5847
R382 VTAIL.n1 VTAIL.n0 58.5846
R383 VTAIL.n147 VTAIL.n146 58.5846
R384 VTAIL.n583 VTAIL.n582 35.4823
R385 VTAIL.n73 VTAIL.n72 35.4823
R386 VTAIL.n145 VTAIL.n144 35.4823
R387 VTAIL.n219 VTAIL.n218 35.4823
R388 VTAIL.n511 VTAIL.n510 35.4823
R389 VTAIL.n437 VTAIL.n436 35.4823
R390 VTAIL.n365 VTAIL.n364 35.4823
R391 VTAIL.n291 VTAIL.n290 35.4823
R392 VTAIL.n583 VTAIL.n511 26.4445
R393 VTAIL.n291 VTAIL.n219 26.4445
R394 VTAIL.n536 VTAIL.n535 16.3895
R395 VTAIL.n26 VTAIL.n25 16.3895
R396 VTAIL.n98 VTAIL.n97 16.3895
R397 VTAIL.n172 VTAIL.n171 16.3895
R398 VTAIL.n464 VTAIL.n463 16.3895
R399 VTAIL.n390 VTAIL.n389 16.3895
R400 VTAIL.n318 VTAIL.n317 16.3895
R401 VTAIL.n244 VTAIL.n243 16.3895
R402 VTAIL.n539 VTAIL.n534 12.8005
R403 VTAIL.n580 VTAIL.n579 12.8005
R404 VTAIL.n29 VTAIL.n24 12.8005
R405 VTAIL.n70 VTAIL.n69 12.8005
R406 VTAIL.n101 VTAIL.n96 12.8005
R407 VTAIL.n142 VTAIL.n141 12.8005
R408 VTAIL.n175 VTAIL.n170 12.8005
R409 VTAIL.n216 VTAIL.n215 12.8005
R410 VTAIL.n508 VTAIL.n507 12.8005
R411 VTAIL.n467 VTAIL.n462 12.8005
R412 VTAIL.n434 VTAIL.n433 12.8005
R413 VTAIL.n393 VTAIL.n388 12.8005
R414 VTAIL.n362 VTAIL.n361 12.8005
R415 VTAIL.n321 VTAIL.n316 12.8005
R416 VTAIL.n288 VTAIL.n287 12.8005
R417 VTAIL.n247 VTAIL.n242 12.8005
R418 VTAIL.n540 VTAIL.n532 12.0247
R419 VTAIL.n576 VTAIL.n514 12.0247
R420 VTAIL.n30 VTAIL.n22 12.0247
R421 VTAIL.n66 VTAIL.n4 12.0247
R422 VTAIL.n102 VTAIL.n94 12.0247
R423 VTAIL.n138 VTAIL.n76 12.0247
R424 VTAIL.n176 VTAIL.n168 12.0247
R425 VTAIL.n212 VTAIL.n150 12.0247
R426 VTAIL.n504 VTAIL.n442 12.0247
R427 VTAIL.n468 VTAIL.n460 12.0247
R428 VTAIL.n430 VTAIL.n368 12.0247
R429 VTAIL.n394 VTAIL.n386 12.0247
R430 VTAIL.n358 VTAIL.n296 12.0247
R431 VTAIL.n322 VTAIL.n314 12.0247
R432 VTAIL.n284 VTAIL.n222 12.0247
R433 VTAIL.n248 VTAIL.n240 12.0247
R434 VTAIL.n544 VTAIL.n543 11.249
R435 VTAIL.n575 VTAIL.n516 11.249
R436 VTAIL.n34 VTAIL.n33 11.249
R437 VTAIL.n65 VTAIL.n6 11.249
R438 VTAIL.n106 VTAIL.n105 11.249
R439 VTAIL.n137 VTAIL.n78 11.249
R440 VTAIL.n180 VTAIL.n179 11.249
R441 VTAIL.n211 VTAIL.n152 11.249
R442 VTAIL.n503 VTAIL.n444 11.249
R443 VTAIL.n472 VTAIL.n471 11.249
R444 VTAIL.n429 VTAIL.n370 11.249
R445 VTAIL.n398 VTAIL.n397 11.249
R446 VTAIL.n357 VTAIL.n298 11.249
R447 VTAIL.n326 VTAIL.n325 11.249
R448 VTAIL.n283 VTAIL.n224 11.249
R449 VTAIL.n252 VTAIL.n251 11.249
R450 VTAIL.n547 VTAIL.n530 10.4732
R451 VTAIL.n572 VTAIL.n571 10.4732
R452 VTAIL.n37 VTAIL.n20 10.4732
R453 VTAIL.n62 VTAIL.n61 10.4732
R454 VTAIL.n109 VTAIL.n92 10.4732
R455 VTAIL.n134 VTAIL.n133 10.4732
R456 VTAIL.n183 VTAIL.n166 10.4732
R457 VTAIL.n208 VTAIL.n207 10.4732
R458 VTAIL.n500 VTAIL.n499 10.4732
R459 VTAIL.n475 VTAIL.n458 10.4732
R460 VTAIL.n426 VTAIL.n425 10.4732
R461 VTAIL.n401 VTAIL.n384 10.4732
R462 VTAIL.n354 VTAIL.n353 10.4732
R463 VTAIL.n329 VTAIL.n312 10.4732
R464 VTAIL.n280 VTAIL.n279 10.4732
R465 VTAIL.n255 VTAIL.n238 10.4732
R466 VTAIL.n548 VTAIL.n528 9.69747
R467 VTAIL.n568 VTAIL.n518 9.69747
R468 VTAIL.n38 VTAIL.n18 9.69747
R469 VTAIL.n58 VTAIL.n8 9.69747
R470 VTAIL.n110 VTAIL.n90 9.69747
R471 VTAIL.n130 VTAIL.n80 9.69747
R472 VTAIL.n184 VTAIL.n164 9.69747
R473 VTAIL.n204 VTAIL.n154 9.69747
R474 VTAIL.n496 VTAIL.n446 9.69747
R475 VTAIL.n476 VTAIL.n456 9.69747
R476 VTAIL.n422 VTAIL.n372 9.69747
R477 VTAIL.n402 VTAIL.n382 9.69747
R478 VTAIL.n350 VTAIL.n300 9.69747
R479 VTAIL.n330 VTAIL.n310 9.69747
R480 VTAIL.n276 VTAIL.n226 9.69747
R481 VTAIL.n256 VTAIL.n236 9.69747
R482 VTAIL.n582 VTAIL.n581 9.45567
R483 VTAIL.n72 VTAIL.n71 9.45567
R484 VTAIL.n144 VTAIL.n143 9.45567
R485 VTAIL.n218 VTAIL.n217 9.45567
R486 VTAIL.n510 VTAIL.n509 9.45567
R487 VTAIL.n436 VTAIL.n435 9.45567
R488 VTAIL.n364 VTAIL.n363 9.45567
R489 VTAIL.n290 VTAIL.n289 9.45567
R490 VTAIL.n557 VTAIL.n556 9.3005
R491 VTAIL.n526 VTAIL.n525 9.3005
R492 VTAIL.n551 VTAIL.n550 9.3005
R493 VTAIL.n549 VTAIL.n548 9.3005
R494 VTAIL.n530 VTAIL.n529 9.3005
R495 VTAIL.n543 VTAIL.n542 9.3005
R496 VTAIL.n541 VTAIL.n540 9.3005
R497 VTAIL.n534 VTAIL.n533 9.3005
R498 VTAIL.n559 VTAIL.n558 9.3005
R499 VTAIL.n522 VTAIL.n521 9.3005
R500 VTAIL.n565 VTAIL.n564 9.3005
R501 VTAIL.n567 VTAIL.n566 9.3005
R502 VTAIL.n518 VTAIL.n517 9.3005
R503 VTAIL.n573 VTAIL.n572 9.3005
R504 VTAIL.n575 VTAIL.n574 9.3005
R505 VTAIL.n514 VTAIL.n513 9.3005
R506 VTAIL.n581 VTAIL.n580 9.3005
R507 VTAIL.n47 VTAIL.n46 9.3005
R508 VTAIL.n16 VTAIL.n15 9.3005
R509 VTAIL.n41 VTAIL.n40 9.3005
R510 VTAIL.n39 VTAIL.n38 9.3005
R511 VTAIL.n20 VTAIL.n19 9.3005
R512 VTAIL.n33 VTAIL.n32 9.3005
R513 VTAIL.n31 VTAIL.n30 9.3005
R514 VTAIL.n24 VTAIL.n23 9.3005
R515 VTAIL.n49 VTAIL.n48 9.3005
R516 VTAIL.n12 VTAIL.n11 9.3005
R517 VTAIL.n55 VTAIL.n54 9.3005
R518 VTAIL.n57 VTAIL.n56 9.3005
R519 VTAIL.n8 VTAIL.n7 9.3005
R520 VTAIL.n63 VTAIL.n62 9.3005
R521 VTAIL.n65 VTAIL.n64 9.3005
R522 VTAIL.n4 VTAIL.n3 9.3005
R523 VTAIL.n71 VTAIL.n70 9.3005
R524 VTAIL.n119 VTAIL.n118 9.3005
R525 VTAIL.n88 VTAIL.n87 9.3005
R526 VTAIL.n113 VTAIL.n112 9.3005
R527 VTAIL.n111 VTAIL.n110 9.3005
R528 VTAIL.n92 VTAIL.n91 9.3005
R529 VTAIL.n105 VTAIL.n104 9.3005
R530 VTAIL.n103 VTAIL.n102 9.3005
R531 VTAIL.n96 VTAIL.n95 9.3005
R532 VTAIL.n121 VTAIL.n120 9.3005
R533 VTAIL.n84 VTAIL.n83 9.3005
R534 VTAIL.n127 VTAIL.n126 9.3005
R535 VTAIL.n129 VTAIL.n128 9.3005
R536 VTAIL.n80 VTAIL.n79 9.3005
R537 VTAIL.n135 VTAIL.n134 9.3005
R538 VTAIL.n137 VTAIL.n136 9.3005
R539 VTAIL.n76 VTAIL.n75 9.3005
R540 VTAIL.n143 VTAIL.n142 9.3005
R541 VTAIL.n193 VTAIL.n192 9.3005
R542 VTAIL.n162 VTAIL.n161 9.3005
R543 VTAIL.n187 VTAIL.n186 9.3005
R544 VTAIL.n185 VTAIL.n184 9.3005
R545 VTAIL.n166 VTAIL.n165 9.3005
R546 VTAIL.n179 VTAIL.n178 9.3005
R547 VTAIL.n177 VTAIL.n176 9.3005
R548 VTAIL.n170 VTAIL.n169 9.3005
R549 VTAIL.n195 VTAIL.n194 9.3005
R550 VTAIL.n158 VTAIL.n157 9.3005
R551 VTAIL.n201 VTAIL.n200 9.3005
R552 VTAIL.n203 VTAIL.n202 9.3005
R553 VTAIL.n154 VTAIL.n153 9.3005
R554 VTAIL.n209 VTAIL.n208 9.3005
R555 VTAIL.n211 VTAIL.n210 9.3005
R556 VTAIL.n150 VTAIL.n149 9.3005
R557 VTAIL.n217 VTAIL.n216 9.3005
R558 VTAIL.n450 VTAIL.n449 9.3005
R559 VTAIL.n493 VTAIL.n492 9.3005
R560 VTAIL.n495 VTAIL.n494 9.3005
R561 VTAIL.n446 VTAIL.n445 9.3005
R562 VTAIL.n501 VTAIL.n500 9.3005
R563 VTAIL.n503 VTAIL.n502 9.3005
R564 VTAIL.n442 VTAIL.n441 9.3005
R565 VTAIL.n509 VTAIL.n508 9.3005
R566 VTAIL.n487 VTAIL.n486 9.3005
R567 VTAIL.n485 VTAIL.n484 9.3005
R568 VTAIL.n454 VTAIL.n453 9.3005
R569 VTAIL.n479 VTAIL.n478 9.3005
R570 VTAIL.n477 VTAIL.n476 9.3005
R571 VTAIL.n458 VTAIL.n457 9.3005
R572 VTAIL.n471 VTAIL.n470 9.3005
R573 VTAIL.n469 VTAIL.n468 9.3005
R574 VTAIL.n462 VTAIL.n461 9.3005
R575 VTAIL.n376 VTAIL.n375 9.3005
R576 VTAIL.n419 VTAIL.n418 9.3005
R577 VTAIL.n421 VTAIL.n420 9.3005
R578 VTAIL.n372 VTAIL.n371 9.3005
R579 VTAIL.n427 VTAIL.n426 9.3005
R580 VTAIL.n429 VTAIL.n428 9.3005
R581 VTAIL.n368 VTAIL.n367 9.3005
R582 VTAIL.n435 VTAIL.n434 9.3005
R583 VTAIL.n413 VTAIL.n412 9.3005
R584 VTAIL.n411 VTAIL.n410 9.3005
R585 VTAIL.n380 VTAIL.n379 9.3005
R586 VTAIL.n405 VTAIL.n404 9.3005
R587 VTAIL.n403 VTAIL.n402 9.3005
R588 VTAIL.n384 VTAIL.n383 9.3005
R589 VTAIL.n397 VTAIL.n396 9.3005
R590 VTAIL.n395 VTAIL.n394 9.3005
R591 VTAIL.n388 VTAIL.n387 9.3005
R592 VTAIL.n304 VTAIL.n303 9.3005
R593 VTAIL.n347 VTAIL.n346 9.3005
R594 VTAIL.n349 VTAIL.n348 9.3005
R595 VTAIL.n300 VTAIL.n299 9.3005
R596 VTAIL.n355 VTAIL.n354 9.3005
R597 VTAIL.n357 VTAIL.n356 9.3005
R598 VTAIL.n296 VTAIL.n295 9.3005
R599 VTAIL.n363 VTAIL.n362 9.3005
R600 VTAIL.n341 VTAIL.n340 9.3005
R601 VTAIL.n339 VTAIL.n338 9.3005
R602 VTAIL.n308 VTAIL.n307 9.3005
R603 VTAIL.n333 VTAIL.n332 9.3005
R604 VTAIL.n331 VTAIL.n330 9.3005
R605 VTAIL.n312 VTAIL.n311 9.3005
R606 VTAIL.n325 VTAIL.n324 9.3005
R607 VTAIL.n323 VTAIL.n322 9.3005
R608 VTAIL.n316 VTAIL.n315 9.3005
R609 VTAIL.n230 VTAIL.n229 9.3005
R610 VTAIL.n273 VTAIL.n272 9.3005
R611 VTAIL.n275 VTAIL.n274 9.3005
R612 VTAIL.n226 VTAIL.n225 9.3005
R613 VTAIL.n281 VTAIL.n280 9.3005
R614 VTAIL.n283 VTAIL.n282 9.3005
R615 VTAIL.n222 VTAIL.n221 9.3005
R616 VTAIL.n289 VTAIL.n288 9.3005
R617 VTAIL.n267 VTAIL.n266 9.3005
R618 VTAIL.n265 VTAIL.n264 9.3005
R619 VTAIL.n234 VTAIL.n233 9.3005
R620 VTAIL.n259 VTAIL.n258 9.3005
R621 VTAIL.n257 VTAIL.n256 9.3005
R622 VTAIL.n238 VTAIL.n237 9.3005
R623 VTAIL.n251 VTAIL.n250 9.3005
R624 VTAIL.n249 VTAIL.n248 9.3005
R625 VTAIL.n242 VTAIL.n241 9.3005
R626 VTAIL.n552 VTAIL.n551 8.92171
R627 VTAIL.n567 VTAIL.n520 8.92171
R628 VTAIL.n42 VTAIL.n41 8.92171
R629 VTAIL.n57 VTAIL.n10 8.92171
R630 VTAIL.n114 VTAIL.n113 8.92171
R631 VTAIL.n129 VTAIL.n82 8.92171
R632 VTAIL.n188 VTAIL.n187 8.92171
R633 VTAIL.n203 VTAIL.n156 8.92171
R634 VTAIL.n495 VTAIL.n448 8.92171
R635 VTAIL.n480 VTAIL.n479 8.92171
R636 VTAIL.n421 VTAIL.n374 8.92171
R637 VTAIL.n406 VTAIL.n405 8.92171
R638 VTAIL.n349 VTAIL.n302 8.92171
R639 VTAIL.n334 VTAIL.n333 8.92171
R640 VTAIL.n275 VTAIL.n228 8.92171
R641 VTAIL.n260 VTAIL.n259 8.92171
R642 VTAIL.n555 VTAIL.n526 8.14595
R643 VTAIL.n564 VTAIL.n563 8.14595
R644 VTAIL.n45 VTAIL.n16 8.14595
R645 VTAIL.n54 VTAIL.n53 8.14595
R646 VTAIL.n117 VTAIL.n88 8.14595
R647 VTAIL.n126 VTAIL.n125 8.14595
R648 VTAIL.n191 VTAIL.n162 8.14595
R649 VTAIL.n200 VTAIL.n199 8.14595
R650 VTAIL.n492 VTAIL.n491 8.14595
R651 VTAIL.n483 VTAIL.n454 8.14595
R652 VTAIL.n418 VTAIL.n417 8.14595
R653 VTAIL.n409 VTAIL.n380 8.14595
R654 VTAIL.n346 VTAIL.n345 8.14595
R655 VTAIL.n337 VTAIL.n308 8.14595
R656 VTAIL.n272 VTAIL.n271 8.14595
R657 VTAIL.n263 VTAIL.n234 8.14595
R658 VTAIL.n582 VTAIL.n512 7.75445
R659 VTAIL.n72 VTAIL.n2 7.75445
R660 VTAIL.n144 VTAIL.n74 7.75445
R661 VTAIL.n218 VTAIL.n148 7.75445
R662 VTAIL.n510 VTAIL.n440 7.75445
R663 VTAIL.n436 VTAIL.n366 7.75445
R664 VTAIL.n364 VTAIL.n294 7.75445
R665 VTAIL.n290 VTAIL.n220 7.75445
R666 VTAIL.n556 VTAIL.n524 7.3702
R667 VTAIL.n560 VTAIL.n522 7.3702
R668 VTAIL.n46 VTAIL.n14 7.3702
R669 VTAIL.n50 VTAIL.n12 7.3702
R670 VTAIL.n118 VTAIL.n86 7.3702
R671 VTAIL.n122 VTAIL.n84 7.3702
R672 VTAIL.n192 VTAIL.n160 7.3702
R673 VTAIL.n196 VTAIL.n158 7.3702
R674 VTAIL.n488 VTAIL.n450 7.3702
R675 VTAIL.n484 VTAIL.n452 7.3702
R676 VTAIL.n414 VTAIL.n376 7.3702
R677 VTAIL.n410 VTAIL.n378 7.3702
R678 VTAIL.n342 VTAIL.n304 7.3702
R679 VTAIL.n338 VTAIL.n306 7.3702
R680 VTAIL.n268 VTAIL.n230 7.3702
R681 VTAIL.n264 VTAIL.n232 7.3702
R682 VTAIL.n559 VTAIL.n524 6.59444
R683 VTAIL.n560 VTAIL.n559 6.59444
R684 VTAIL.n49 VTAIL.n14 6.59444
R685 VTAIL.n50 VTAIL.n49 6.59444
R686 VTAIL.n121 VTAIL.n86 6.59444
R687 VTAIL.n122 VTAIL.n121 6.59444
R688 VTAIL.n195 VTAIL.n160 6.59444
R689 VTAIL.n196 VTAIL.n195 6.59444
R690 VTAIL.n488 VTAIL.n487 6.59444
R691 VTAIL.n487 VTAIL.n452 6.59444
R692 VTAIL.n414 VTAIL.n413 6.59444
R693 VTAIL.n413 VTAIL.n378 6.59444
R694 VTAIL.n342 VTAIL.n341 6.59444
R695 VTAIL.n341 VTAIL.n306 6.59444
R696 VTAIL.n268 VTAIL.n267 6.59444
R697 VTAIL.n267 VTAIL.n232 6.59444
R698 VTAIL.n580 VTAIL.n512 6.08283
R699 VTAIL.n70 VTAIL.n2 6.08283
R700 VTAIL.n142 VTAIL.n74 6.08283
R701 VTAIL.n216 VTAIL.n148 6.08283
R702 VTAIL.n508 VTAIL.n440 6.08283
R703 VTAIL.n434 VTAIL.n366 6.08283
R704 VTAIL.n362 VTAIL.n294 6.08283
R705 VTAIL.n288 VTAIL.n220 6.08283
R706 VTAIL.n556 VTAIL.n555 5.81868
R707 VTAIL.n563 VTAIL.n522 5.81868
R708 VTAIL.n46 VTAIL.n45 5.81868
R709 VTAIL.n53 VTAIL.n12 5.81868
R710 VTAIL.n118 VTAIL.n117 5.81868
R711 VTAIL.n125 VTAIL.n84 5.81868
R712 VTAIL.n192 VTAIL.n191 5.81868
R713 VTAIL.n199 VTAIL.n158 5.81868
R714 VTAIL.n491 VTAIL.n450 5.81868
R715 VTAIL.n484 VTAIL.n483 5.81868
R716 VTAIL.n417 VTAIL.n376 5.81868
R717 VTAIL.n410 VTAIL.n409 5.81868
R718 VTAIL.n345 VTAIL.n304 5.81868
R719 VTAIL.n338 VTAIL.n337 5.81868
R720 VTAIL.n271 VTAIL.n230 5.81868
R721 VTAIL.n264 VTAIL.n263 5.81868
R722 VTAIL.n552 VTAIL.n526 5.04292
R723 VTAIL.n564 VTAIL.n520 5.04292
R724 VTAIL.n42 VTAIL.n16 5.04292
R725 VTAIL.n54 VTAIL.n10 5.04292
R726 VTAIL.n114 VTAIL.n88 5.04292
R727 VTAIL.n126 VTAIL.n82 5.04292
R728 VTAIL.n188 VTAIL.n162 5.04292
R729 VTAIL.n200 VTAIL.n156 5.04292
R730 VTAIL.n492 VTAIL.n448 5.04292
R731 VTAIL.n480 VTAIL.n454 5.04292
R732 VTAIL.n418 VTAIL.n374 5.04292
R733 VTAIL.n406 VTAIL.n380 5.04292
R734 VTAIL.n346 VTAIL.n302 5.04292
R735 VTAIL.n334 VTAIL.n308 5.04292
R736 VTAIL.n272 VTAIL.n228 5.04292
R737 VTAIL.n260 VTAIL.n234 5.04292
R738 VTAIL.n551 VTAIL.n528 4.26717
R739 VTAIL.n568 VTAIL.n567 4.26717
R740 VTAIL.n41 VTAIL.n18 4.26717
R741 VTAIL.n58 VTAIL.n57 4.26717
R742 VTAIL.n113 VTAIL.n90 4.26717
R743 VTAIL.n130 VTAIL.n129 4.26717
R744 VTAIL.n187 VTAIL.n164 4.26717
R745 VTAIL.n204 VTAIL.n203 4.26717
R746 VTAIL.n496 VTAIL.n495 4.26717
R747 VTAIL.n479 VTAIL.n456 4.26717
R748 VTAIL.n422 VTAIL.n421 4.26717
R749 VTAIL.n405 VTAIL.n382 4.26717
R750 VTAIL.n350 VTAIL.n349 4.26717
R751 VTAIL.n333 VTAIL.n310 4.26717
R752 VTAIL.n276 VTAIL.n275 4.26717
R753 VTAIL.n259 VTAIL.n236 4.26717
R754 VTAIL.n535 VTAIL.n533 3.70982
R755 VTAIL.n25 VTAIL.n23 3.70982
R756 VTAIL.n97 VTAIL.n95 3.70982
R757 VTAIL.n171 VTAIL.n169 3.70982
R758 VTAIL.n463 VTAIL.n461 3.70982
R759 VTAIL.n389 VTAIL.n387 3.70982
R760 VTAIL.n317 VTAIL.n315 3.70982
R761 VTAIL.n243 VTAIL.n241 3.70982
R762 VTAIL.n548 VTAIL.n547 3.49141
R763 VTAIL.n571 VTAIL.n518 3.49141
R764 VTAIL.n38 VTAIL.n37 3.49141
R765 VTAIL.n61 VTAIL.n8 3.49141
R766 VTAIL.n110 VTAIL.n109 3.49141
R767 VTAIL.n133 VTAIL.n80 3.49141
R768 VTAIL.n184 VTAIL.n183 3.49141
R769 VTAIL.n207 VTAIL.n154 3.49141
R770 VTAIL.n499 VTAIL.n446 3.49141
R771 VTAIL.n476 VTAIL.n475 3.49141
R772 VTAIL.n425 VTAIL.n372 3.49141
R773 VTAIL.n402 VTAIL.n401 3.49141
R774 VTAIL.n353 VTAIL.n300 3.49141
R775 VTAIL.n330 VTAIL.n329 3.49141
R776 VTAIL.n279 VTAIL.n226 3.49141
R777 VTAIL.n256 VTAIL.n255 3.49141
R778 VTAIL.n544 VTAIL.n530 2.71565
R779 VTAIL.n572 VTAIL.n516 2.71565
R780 VTAIL.n34 VTAIL.n20 2.71565
R781 VTAIL.n62 VTAIL.n6 2.71565
R782 VTAIL.n106 VTAIL.n92 2.71565
R783 VTAIL.n134 VTAIL.n78 2.71565
R784 VTAIL.n180 VTAIL.n166 2.71565
R785 VTAIL.n208 VTAIL.n152 2.71565
R786 VTAIL.n500 VTAIL.n444 2.71565
R787 VTAIL.n472 VTAIL.n458 2.71565
R788 VTAIL.n426 VTAIL.n370 2.71565
R789 VTAIL.n398 VTAIL.n384 2.71565
R790 VTAIL.n354 VTAIL.n298 2.71565
R791 VTAIL.n326 VTAIL.n312 2.71565
R792 VTAIL.n280 VTAIL.n224 2.71565
R793 VTAIL.n252 VTAIL.n238 2.71565
R794 VTAIL.n293 VTAIL.n291 2.55222
R795 VTAIL.n365 VTAIL.n293 2.55222
R796 VTAIL.n439 VTAIL.n437 2.55222
R797 VTAIL.n511 VTAIL.n439 2.55222
R798 VTAIL.n219 VTAIL.n147 2.55222
R799 VTAIL.n147 VTAIL.n145 2.55222
R800 VTAIL.n73 VTAIL.n1 2.55222
R801 VTAIL VTAIL.n583 2.49403
R802 VTAIL.n0 VTAIL.t15 2.43169
R803 VTAIL.n0 VTAIL.t10 2.43169
R804 VTAIL.n146 VTAIL.t2 2.43169
R805 VTAIL.n146 VTAIL.t7 2.43169
R806 VTAIL.n438 VTAIL.t1 2.43169
R807 VTAIL.n438 VTAIL.t0 2.43169
R808 VTAIL.n292 VTAIL.t14 2.43169
R809 VTAIL.n292 VTAIL.t13 2.43169
R810 VTAIL.n543 VTAIL.n532 1.93989
R811 VTAIL.n576 VTAIL.n575 1.93989
R812 VTAIL.n33 VTAIL.n22 1.93989
R813 VTAIL.n66 VTAIL.n65 1.93989
R814 VTAIL.n105 VTAIL.n94 1.93989
R815 VTAIL.n138 VTAIL.n137 1.93989
R816 VTAIL.n179 VTAIL.n168 1.93989
R817 VTAIL.n212 VTAIL.n211 1.93989
R818 VTAIL.n504 VTAIL.n503 1.93989
R819 VTAIL.n471 VTAIL.n460 1.93989
R820 VTAIL.n430 VTAIL.n429 1.93989
R821 VTAIL.n397 VTAIL.n386 1.93989
R822 VTAIL.n358 VTAIL.n357 1.93989
R823 VTAIL.n325 VTAIL.n314 1.93989
R824 VTAIL.n284 VTAIL.n283 1.93989
R825 VTAIL.n251 VTAIL.n240 1.93989
R826 VTAIL.n540 VTAIL.n539 1.16414
R827 VTAIL.n579 VTAIL.n514 1.16414
R828 VTAIL.n30 VTAIL.n29 1.16414
R829 VTAIL.n69 VTAIL.n4 1.16414
R830 VTAIL.n102 VTAIL.n101 1.16414
R831 VTAIL.n141 VTAIL.n76 1.16414
R832 VTAIL.n176 VTAIL.n175 1.16414
R833 VTAIL.n215 VTAIL.n150 1.16414
R834 VTAIL.n507 VTAIL.n442 1.16414
R835 VTAIL.n468 VTAIL.n467 1.16414
R836 VTAIL.n433 VTAIL.n368 1.16414
R837 VTAIL.n394 VTAIL.n393 1.16414
R838 VTAIL.n361 VTAIL.n296 1.16414
R839 VTAIL.n322 VTAIL.n321 1.16414
R840 VTAIL.n287 VTAIL.n222 1.16414
R841 VTAIL.n248 VTAIL.n247 1.16414
R842 VTAIL.n437 VTAIL.n365 0.470328
R843 VTAIL.n145 VTAIL.n73 0.470328
R844 VTAIL.n536 VTAIL.n534 0.388379
R845 VTAIL.n26 VTAIL.n24 0.388379
R846 VTAIL.n98 VTAIL.n96 0.388379
R847 VTAIL.n172 VTAIL.n170 0.388379
R848 VTAIL.n464 VTAIL.n462 0.388379
R849 VTAIL.n390 VTAIL.n388 0.388379
R850 VTAIL.n318 VTAIL.n316 0.388379
R851 VTAIL.n244 VTAIL.n242 0.388379
R852 VTAIL.n541 VTAIL.n533 0.155672
R853 VTAIL.n542 VTAIL.n541 0.155672
R854 VTAIL.n542 VTAIL.n529 0.155672
R855 VTAIL.n549 VTAIL.n529 0.155672
R856 VTAIL.n550 VTAIL.n549 0.155672
R857 VTAIL.n550 VTAIL.n525 0.155672
R858 VTAIL.n557 VTAIL.n525 0.155672
R859 VTAIL.n558 VTAIL.n557 0.155672
R860 VTAIL.n558 VTAIL.n521 0.155672
R861 VTAIL.n565 VTAIL.n521 0.155672
R862 VTAIL.n566 VTAIL.n565 0.155672
R863 VTAIL.n566 VTAIL.n517 0.155672
R864 VTAIL.n573 VTAIL.n517 0.155672
R865 VTAIL.n574 VTAIL.n573 0.155672
R866 VTAIL.n574 VTAIL.n513 0.155672
R867 VTAIL.n581 VTAIL.n513 0.155672
R868 VTAIL.n31 VTAIL.n23 0.155672
R869 VTAIL.n32 VTAIL.n31 0.155672
R870 VTAIL.n32 VTAIL.n19 0.155672
R871 VTAIL.n39 VTAIL.n19 0.155672
R872 VTAIL.n40 VTAIL.n39 0.155672
R873 VTAIL.n40 VTAIL.n15 0.155672
R874 VTAIL.n47 VTAIL.n15 0.155672
R875 VTAIL.n48 VTAIL.n47 0.155672
R876 VTAIL.n48 VTAIL.n11 0.155672
R877 VTAIL.n55 VTAIL.n11 0.155672
R878 VTAIL.n56 VTAIL.n55 0.155672
R879 VTAIL.n56 VTAIL.n7 0.155672
R880 VTAIL.n63 VTAIL.n7 0.155672
R881 VTAIL.n64 VTAIL.n63 0.155672
R882 VTAIL.n64 VTAIL.n3 0.155672
R883 VTAIL.n71 VTAIL.n3 0.155672
R884 VTAIL.n103 VTAIL.n95 0.155672
R885 VTAIL.n104 VTAIL.n103 0.155672
R886 VTAIL.n104 VTAIL.n91 0.155672
R887 VTAIL.n111 VTAIL.n91 0.155672
R888 VTAIL.n112 VTAIL.n111 0.155672
R889 VTAIL.n112 VTAIL.n87 0.155672
R890 VTAIL.n119 VTAIL.n87 0.155672
R891 VTAIL.n120 VTAIL.n119 0.155672
R892 VTAIL.n120 VTAIL.n83 0.155672
R893 VTAIL.n127 VTAIL.n83 0.155672
R894 VTAIL.n128 VTAIL.n127 0.155672
R895 VTAIL.n128 VTAIL.n79 0.155672
R896 VTAIL.n135 VTAIL.n79 0.155672
R897 VTAIL.n136 VTAIL.n135 0.155672
R898 VTAIL.n136 VTAIL.n75 0.155672
R899 VTAIL.n143 VTAIL.n75 0.155672
R900 VTAIL.n177 VTAIL.n169 0.155672
R901 VTAIL.n178 VTAIL.n177 0.155672
R902 VTAIL.n178 VTAIL.n165 0.155672
R903 VTAIL.n185 VTAIL.n165 0.155672
R904 VTAIL.n186 VTAIL.n185 0.155672
R905 VTAIL.n186 VTAIL.n161 0.155672
R906 VTAIL.n193 VTAIL.n161 0.155672
R907 VTAIL.n194 VTAIL.n193 0.155672
R908 VTAIL.n194 VTAIL.n157 0.155672
R909 VTAIL.n201 VTAIL.n157 0.155672
R910 VTAIL.n202 VTAIL.n201 0.155672
R911 VTAIL.n202 VTAIL.n153 0.155672
R912 VTAIL.n209 VTAIL.n153 0.155672
R913 VTAIL.n210 VTAIL.n209 0.155672
R914 VTAIL.n210 VTAIL.n149 0.155672
R915 VTAIL.n217 VTAIL.n149 0.155672
R916 VTAIL.n509 VTAIL.n441 0.155672
R917 VTAIL.n502 VTAIL.n441 0.155672
R918 VTAIL.n502 VTAIL.n501 0.155672
R919 VTAIL.n501 VTAIL.n445 0.155672
R920 VTAIL.n494 VTAIL.n445 0.155672
R921 VTAIL.n494 VTAIL.n493 0.155672
R922 VTAIL.n493 VTAIL.n449 0.155672
R923 VTAIL.n486 VTAIL.n449 0.155672
R924 VTAIL.n486 VTAIL.n485 0.155672
R925 VTAIL.n485 VTAIL.n453 0.155672
R926 VTAIL.n478 VTAIL.n453 0.155672
R927 VTAIL.n478 VTAIL.n477 0.155672
R928 VTAIL.n477 VTAIL.n457 0.155672
R929 VTAIL.n470 VTAIL.n457 0.155672
R930 VTAIL.n470 VTAIL.n469 0.155672
R931 VTAIL.n469 VTAIL.n461 0.155672
R932 VTAIL.n435 VTAIL.n367 0.155672
R933 VTAIL.n428 VTAIL.n367 0.155672
R934 VTAIL.n428 VTAIL.n427 0.155672
R935 VTAIL.n427 VTAIL.n371 0.155672
R936 VTAIL.n420 VTAIL.n371 0.155672
R937 VTAIL.n420 VTAIL.n419 0.155672
R938 VTAIL.n419 VTAIL.n375 0.155672
R939 VTAIL.n412 VTAIL.n375 0.155672
R940 VTAIL.n412 VTAIL.n411 0.155672
R941 VTAIL.n411 VTAIL.n379 0.155672
R942 VTAIL.n404 VTAIL.n379 0.155672
R943 VTAIL.n404 VTAIL.n403 0.155672
R944 VTAIL.n403 VTAIL.n383 0.155672
R945 VTAIL.n396 VTAIL.n383 0.155672
R946 VTAIL.n396 VTAIL.n395 0.155672
R947 VTAIL.n395 VTAIL.n387 0.155672
R948 VTAIL.n363 VTAIL.n295 0.155672
R949 VTAIL.n356 VTAIL.n295 0.155672
R950 VTAIL.n356 VTAIL.n355 0.155672
R951 VTAIL.n355 VTAIL.n299 0.155672
R952 VTAIL.n348 VTAIL.n299 0.155672
R953 VTAIL.n348 VTAIL.n347 0.155672
R954 VTAIL.n347 VTAIL.n303 0.155672
R955 VTAIL.n340 VTAIL.n303 0.155672
R956 VTAIL.n340 VTAIL.n339 0.155672
R957 VTAIL.n339 VTAIL.n307 0.155672
R958 VTAIL.n332 VTAIL.n307 0.155672
R959 VTAIL.n332 VTAIL.n331 0.155672
R960 VTAIL.n331 VTAIL.n311 0.155672
R961 VTAIL.n324 VTAIL.n311 0.155672
R962 VTAIL.n324 VTAIL.n323 0.155672
R963 VTAIL.n323 VTAIL.n315 0.155672
R964 VTAIL.n289 VTAIL.n221 0.155672
R965 VTAIL.n282 VTAIL.n221 0.155672
R966 VTAIL.n282 VTAIL.n281 0.155672
R967 VTAIL.n281 VTAIL.n225 0.155672
R968 VTAIL.n274 VTAIL.n225 0.155672
R969 VTAIL.n274 VTAIL.n273 0.155672
R970 VTAIL.n273 VTAIL.n229 0.155672
R971 VTAIL.n266 VTAIL.n229 0.155672
R972 VTAIL.n266 VTAIL.n265 0.155672
R973 VTAIL.n265 VTAIL.n233 0.155672
R974 VTAIL.n258 VTAIL.n233 0.155672
R975 VTAIL.n258 VTAIL.n257 0.155672
R976 VTAIL.n257 VTAIL.n237 0.155672
R977 VTAIL.n250 VTAIL.n237 0.155672
R978 VTAIL.n250 VTAIL.n249 0.155672
R979 VTAIL.n249 VTAIL.n241 0.155672
R980 VTAIL VTAIL.n1 0.0586897
R981 VDD2.n2 VDD2.n1 76.4839
R982 VDD2.n2 VDD2.n0 76.4839
R983 VDD2 VDD2.n5 76.481
R984 VDD2.n4 VDD2.n3 75.2635
R985 VDD2.n4 VDD2.n2 46.7239
R986 VDD2.n5 VDD2.t5 2.43169
R987 VDD2.n5 VDD2.t4 2.43169
R988 VDD2.n3 VDD2.t0 2.43169
R989 VDD2.n3 VDD2.t6 2.43169
R990 VDD2.n1 VDD2.t2 2.43169
R991 VDD2.n1 VDD2.t3 2.43169
R992 VDD2.n0 VDD2.t1 2.43169
R993 VDD2.n0 VDD2.t7 2.43169
R994 VDD2 VDD2.n4 1.33455
R995 B.n442 B.n135 585
R996 B.n441 B.n440 585
R997 B.n439 B.n136 585
R998 B.n438 B.n437 585
R999 B.n436 B.n137 585
R1000 B.n435 B.n434 585
R1001 B.n433 B.n138 585
R1002 B.n432 B.n431 585
R1003 B.n430 B.n139 585
R1004 B.n429 B.n428 585
R1005 B.n427 B.n140 585
R1006 B.n426 B.n425 585
R1007 B.n424 B.n141 585
R1008 B.n423 B.n422 585
R1009 B.n421 B.n142 585
R1010 B.n420 B.n419 585
R1011 B.n418 B.n143 585
R1012 B.n417 B.n416 585
R1013 B.n415 B.n144 585
R1014 B.n414 B.n413 585
R1015 B.n412 B.n145 585
R1016 B.n411 B.n410 585
R1017 B.n409 B.n146 585
R1018 B.n408 B.n407 585
R1019 B.n406 B.n147 585
R1020 B.n405 B.n404 585
R1021 B.n403 B.n148 585
R1022 B.n402 B.n401 585
R1023 B.n400 B.n149 585
R1024 B.n399 B.n398 585
R1025 B.n397 B.n150 585
R1026 B.n396 B.n395 585
R1027 B.n394 B.n151 585
R1028 B.n393 B.n392 585
R1029 B.n391 B.n152 585
R1030 B.n390 B.n389 585
R1031 B.n388 B.n153 585
R1032 B.n387 B.n386 585
R1033 B.n385 B.n154 585
R1034 B.n384 B.n383 585
R1035 B.n382 B.n155 585
R1036 B.n381 B.n380 585
R1037 B.n379 B.n156 585
R1038 B.n378 B.n377 585
R1039 B.n376 B.n157 585
R1040 B.n375 B.n374 585
R1041 B.n372 B.n158 585
R1042 B.n371 B.n370 585
R1043 B.n369 B.n161 585
R1044 B.n368 B.n367 585
R1045 B.n366 B.n162 585
R1046 B.n365 B.n364 585
R1047 B.n363 B.n163 585
R1048 B.n362 B.n361 585
R1049 B.n360 B.n164 585
R1050 B.n358 B.n357 585
R1051 B.n356 B.n167 585
R1052 B.n355 B.n354 585
R1053 B.n353 B.n168 585
R1054 B.n352 B.n351 585
R1055 B.n350 B.n169 585
R1056 B.n349 B.n348 585
R1057 B.n347 B.n170 585
R1058 B.n346 B.n345 585
R1059 B.n344 B.n171 585
R1060 B.n343 B.n342 585
R1061 B.n341 B.n172 585
R1062 B.n340 B.n339 585
R1063 B.n338 B.n173 585
R1064 B.n337 B.n336 585
R1065 B.n335 B.n174 585
R1066 B.n334 B.n333 585
R1067 B.n332 B.n175 585
R1068 B.n331 B.n330 585
R1069 B.n329 B.n176 585
R1070 B.n328 B.n327 585
R1071 B.n326 B.n177 585
R1072 B.n325 B.n324 585
R1073 B.n323 B.n178 585
R1074 B.n322 B.n321 585
R1075 B.n320 B.n179 585
R1076 B.n319 B.n318 585
R1077 B.n317 B.n180 585
R1078 B.n316 B.n315 585
R1079 B.n314 B.n181 585
R1080 B.n313 B.n312 585
R1081 B.n311 B.n182 585
R1082 B.n310 B.n309 585
R1083 B.n308 B.n183 585
R1084 B.n307 B.n306 585
R1085 B.n305 B.n184 585
R1086 B.n304 B.n303 585
R1087 B.n302 B.n185 585
R1088 B.n301 B.n300 585
R1089 B.n299 B.n186 585
R1090 B.n298 B.n297 585
R1091 B.n296 B.n187 585
R1092 B.n295 B.n294 585
R1093 B.n293 B.n188 585
R1094 B.n292 B.n291 585
R1095 B.n290 B.n189 585
R1096 B.n444 B.n443 585
R1097 B.n445 B.n134 585
R1098 B.n447 B.n446 585
R1099 B.n448 B.n133 585
R1100 B.n450 B.n449 585
R1101 B.n451 B.n132 585
R1102 B.n453 B.n452 585
R1103 B.n454 B.n131 585
R1104 B.n456 B.n455 585
R1105 B.n457 B.n130 585
R1106 B.n459 B.n458 585
R1107 B.n460 B.n129 585
R1108 B.n462 B.n461 585
R1109 B.n463 B.n128 585
R1110 B.n465 B.n464 585
R1111 B.n466 B.n127 585
R1112 B.n468 B.n467 585
R1113 B.n469 B.n126 585
R1114 B.n471 B.n470 585
R1115 B.n472 B.n125 585
R1116 B.n474 B.n473 585
R1117 B.n475 B.n124 585
R1118 B.n477 B.n476 585
R1119 B.n478 B.n123 585
R1120 B.n480 B.n479 585
R1121 B.n481 B.n122 585
R1122 B.n483 B.n482 585
R1123 B.n484 B.n121 585
R1124 B.n486 B.n485 585
R1125 B.n487 B.n120 585
R1126 B.n489 B.n488 585
R1127 B.n490 B.n119 585
R1128 B.n492 B.n491 585
R1129 B.n493 B.n118 585
R1130 B.n495 B.n494 585
R1131 B.n496 B.n117 585
R1132 B.n498 B.n497 585
R1133 B.n499 B.n116 585
R1134 B.n501 B.n500 585
R1135 B.n502 B.n115 585
R1136 B.n504 B.n503 585
R1137 B.n505 B.n114 585
R1138 B.n507 B.n506 585
R1139 B.n508 B.n113 585
R1140 B.n510 B.n509 585
R1141 B.n511 B.n112 585
R1142 B.n513 B.n512 585
R1143 B.n514 B.n111 585
R1144 B.n516 B.n515 585
R1145 B.n517 B.n110 585
R1146 B.n519 B.n518 585
R1147 B.n520 B.n109 585
R1148 B.n522 B.n521 585
R1149 B.n523 B.n108 585
R1150 B.n525 B.n524 585
R1151 B.n526 B.n107 585
R1152 B.n528 B.n527 585
R1153 B.n529 B.n106 585
R1154 B.n531 B.n530 585
R1155 B.n532 B.n105 585
R1156 B.n534 B.n533 585
R1157 B.n535 B.n104 585
R1158 B.n537 B.n536 585
R1159 B.n538 B.n103 585
R1160 B.n540 B.n539 585
R1161 B.n541 B.n102 585
R1162 B.n543 B.n542 585
R1163 B.n544 B.n101 585
R1164 B.n546 B.n545 585
R1165 B.n547 B.n100 585
R1166 B.n549 B.n548 585
R1167 B.n550 B.n99 585
R1168 B.n552 B.n551 585
R1169 B.n553 B.n98 585
R1170 B.n555 B.n554 585
R1171 B.n556 B.n97 585
R1172 B.n558 B.n557 585
R1173 B.n559 B.n96 585
R1174 B.n561 B.n560 585
R1175 B.n562 B.n95 585
R1176 B.n564 B.n563 585
R1177 B.n565 B.n94 585
R1178 B.n567 B.n566 585
R1179 B.n568 B.n93 585
R1180 B.n570 B.n569 585
R1181 B.n571 B.n92 585
R1182 B.n573 B.n572 585
R1183 B.n574 B.n91 585
R1184 B.n576 B.n575 585
R1185 B.n577 B.n90 585
R1186 B.n579 B.n578 585
R1187 B.n580 B.n89 585
R1188 B.n582 B.n581 585
R1189 B.n583 B.n88 585
R1190 B.n585 B.n584 585
R1191 B.n586 B.n87 585
R1192 B.n588 B.n587 585
R1193 B.n589 B.n86 585
R1194 B.n591 B.n590 585
R1195 B.n592 B.n85 585
R1196 B.n594 B.n593 585
R1197 B.n595 B.n84 585
R1198 B.n597 B.n596 585
R1199 B.n598 B.n83 585
R1200 B.n751 B.n750 585
R1201 B.n749 B.n28 585
R1202 B.n748 B.n747 585
R1203 B.n746 B.n29 585
R1204 B.n745 B.n744 585
R1205 B.n743 B.n30 585
R1206 B.n742 B.n741 585
R1207 B.n740 B.n31 585
R1208 B.n739 B.n738 585
R1209 B.n737 B.n32 585
R1210 B.n736 B.n735 585
R1211 B.n734 B.n33 585
R1212 B.n733 B.n732 585
R1213 B.n731 B.n34 585
R1214 B.n730 B.n729 585
R1215 B.n728 B.n35 585
R1216 B.n727 B.n726 585
R1217 B.n725 B.n36 585
R1218 B.n724 B.n723 585
R1219 B.n722 B.n37 585
R1220 B.n721 B.n720 585
R1221 B.n719 B.n38 585
R1222 B.n718 B.n717 585
R1223 B.n716 B.n39 585
R1224 B.n715 B.n714 585
R1225 B.n713 B.n40 585
R1226 B.n712 B.n711 585
R1227 B.n710 B.n41 585
R1228 B.n709 B.n708 585
R1229 B.n707 B.n42 585
R1230 B.n706 B.n705 585
R1231 B.n704 B.n43 585
R1232 B.n703 B.n702 585
R1233 B.n701 B.n44 585
R1234 B.n700 B.n699 585
R1235 B.n698 B.n45 585
R1236 B.n697 B.n696 585
R1237 B.n695 B.n46 585
R1238 B.n694 B.n693 585
R1239 B.n692 B.n47 585
R1240 B.n691 B.n690 585
R1241 B.n689 B.n48 585
R1242 B.n688 B.n687 585
R1243 B.n686 B.n49 585
R1244 B.n685 B.n684 585
R1245 B.n683 B.n50 585
R1246 B.n682 B.n681 585
R1247 B.n680 B.n51 585
R1248 B.n679 B.n678 585
R1249 B.n677 B.n55 585
R1250 B.n676 B.n675 585
R1251 B.n674 B.n56 585
R1252 B.n673 B.n672 585
R1253 B.n671 B.n57 585
R1254 B.n670 B.n669 585
R1255 B.n667 B.n58 585
R1256 B.n666 B.n665 585
R1257 B.n664 B.n61 585
R1258 B.n663 B.n662 585
R1259 B.n661 B.n62 585
R1260 B.n660 B.n659 585
R1261 B.n658 B.n63 585
R1262 B.n657 B.n656 585
R1263 B.n655 B.n64 585
R1264 B.n654 B.n653 585
R1265 B.n652 B.n65 585
R1266 B.n651 B.n650 585
R1267 B.n649 B.n66 585
R1268 B.n648 B.n647 585
R1269 B.n646 B.n67 585
R1270 B.n645 B.n644 585
R1271 B.n643 B.n68 585
R1272 B.n642 B.n641 585
R1273 B.n640 B.n69 585
R1274 B.n639 B.n638 585
R1275 B.n637 B.n70 585
R1276 B.n636 B.n635 585
R1277 B.n634 B.n71 585
R1278 B.n633 B.n632 585
R1279 B.n631 B.n72 585
R1280 B.n630 B.n629 585
R1281 B.n628 B.n73 585
R1282 B.n627 B.n626 585
R1283 B.n625 B.n74 585
R1284 B.n624 B.n623 585
R1285 B.n622 B.n75 585
R1286 B.n621 B.n620 585
R1287 B.n619 B.n76 585
R1288 B.n618 B.n617 585
R1289 B.n616 B.n77 585
R1290 B.n615 B.n614 585
R1291 B.n613 B.n78 585
R1292 B.n612 B.n611 585
R1293 B.n610 B.n79 585
R1294 B.n609 B.n608 585
R1295 B.n607 B.n80 585
R1296 B.n606 B.n605 585
R1297 B.n604 B.n81 585
R1298 B.n603 B.n602 585
R1299 B.n601 B.n82 585
R1300 B.n600 B.n599 585
R1301 B.n752 B.n27 585
R1302 B.n754 B.n753 585
R1303 B.n755 B.n26 585
R1304 B.n757 B.n756 585
R1305 B.n758 B.n25 585
R1306 B.n760 B.n759 585
R1307 B.n761 B.n24 585
R1308 B.n763 B.n762 585
R1309 B.n764 B.n23 585
R1310 B.n766 B.n765 585
R1311 B.n767 B.n22 585
R1312 B.n769 B.n768 585
R1313 B.n770 B.n21 585
R1314 B.n772 B.n771 585
R1315 B.n773 B.n20 585
R1316 B.n775 B.n774 585
R1317 B.n776 B.n19 585
R1318 B.n778 B.n777 585
R1319 B.n779 B.n18 585
R1320 B.n781 B.n780 585
R1321 B.n782 B.n17 585
R1322 B.n784 B.n783 585
R1323 B.n785 B.n16 585
R1324 B.n787 B.n786 585
R1325 B.n788 B.n15 585
R1326 B.n790 B.n789 585
R1327 B.n791 B.n14 585
R1328 B.n793 B.n792 585
R1329 B.n794 B.n13 585
R1330 B.n796 B.n795 585
R1331 B.n797 B.n12 585
R1332 B.n799 B.n798 585
R1333 B.n800 B.n11 585
R1334 B.n802 B.n801 585
R1335 B.n803 B.n10 585
R1336 B.n805 B.n804 585
R1337 B.n806 B.n9 585
R1338 B.n808 B.n807 585
R1339 B.n809 B.n8 585
R1340 B.n811 B.n810 585
R1341 B.n812 B.n7 585
R1342 B.n814 B.n813 585
R1343 B.n815 B.n6 585
R1344 B.n817 B.n816 585
R1345 B.n818 B.n5 585
R1346 B.n820 B.n819 585
R1347 B.n821 B.n4 585
R1348 B.n823 B.n822 585
R1349 B.n824 B.n3 585
R1350 B.n826 B.n825 585
R1351 B.n827 B.n0 585
R1352 B.n2 B.n1 585
R1353 B.n215 B.n214 585
R1354 B.n217 B.n216 585
R1355 B.n218 B.n213 585
R1356 B.n220 B.n219 585
R1357 B.n221 B.n212 585
R1358 B.n223 B.n222 585
R1359 B.n224 B.n211 585
R1360 B.n226 B.n225 585
R1361 B.n227 B.n210 585
R1362 B.n229 B.n228 585
R1363 B.n230 B.n209 585
R1364 B.n232 B.n231 585
R1365 B.n233 B.n208 585
R1366 B.n235 B.n234 585
R1367 B.n236 B.n207 585
R1368 B.n238 B.n237 585
R1369 B.n239 B.n206 585
R1370 B.n241 B.n240 585
R1371 B.n242 B.n205 585
R1372 B.n244 B.n243 585
R1373 B.n245 B.n204 585
R1374 B.n247 B.n246 585
R1375 B.n248 B.n203 585
R1376 B.n250 B.n249 585
R1377 B.n251 B.n202 585
R1378 B.n253 B.n252 585
R1379 B.n254 B.n201 585
R1380 B.n256 B.n255 585
R1381 B.n257 B.n200 585
R1382 B.n259 B.n258 585
R1383 B.n260 B.n199 585
R1384 B.n262 B.n261 585
R1385 B.n263 B.n198 585
R1386 B.n265 B.n264 585
R1387 B.n266 B.n197 585
R1388 B.n268 B.n267 585
R1389 B.n269 B.n196 585
R1390 B.n271 B.n270 585
R1391 B.n272 B.n195 585
R1392 B.n274 B.n273 585
R1393 B.n275 B.n194 585
R1394 B.n277 B.n276 585
R1395 B.n278 B.n193 585
R1396 B.n280 B.n279 585
R1397 B.n281 B.n192 585
R1398 B.n283 B.n282 585
R1399 B.n284 B.n191 585
R1400 B.n286 B.n285 585
R1401 B.n287 B.n190 585
R1402 B.n289 B.n288 585
R1403 B.n290 B.n289 511.721
R1404 B.n443 B.n442 511.721
R1405 B.n599 B.n598 511.721
R1406 B.n750 B.n27 511.721
R1407 B.n159 B.t1 457.625
R1408 B.n59 B.t8 457.625
R1409 B.n165 B.t4 457.625
R1410 B.n52 B.t11 457.625
R1411 B.n160 B.t2 400.219
R1412 B.n60 B.t7 400.219
R1413 B.n166 B.t5 400.219
R1414 B.n53 B.t10 400.219
R1415 B.n165 B.t3 330.608
R1416 B.n159 B.t0 330.608
R1417 B.n59 B.t6 330.608
R1418 B.n52 B.t9 330.608
R1419 B.n829 B.n828 256.663
R1420 B.n828 B.n827 235.042
R1421 B.n828 B.n2 235.042
R1422 B.n291 B.n290 163.367
R1423 B.n291 B.n188 163.367
R1424 B.n295 B.n188 163.367
R1425 B.n296 B.n295 163.367
R1426 B.n297 B.n296 163.367
R1427 B.n297 B.n186 163.367
R1428 B.n301 B.n186 163.367
R1429 B.n302 B.n301 163.367
R1430 B.n303 B.n302 163.367
R1431 B.n303 B.n184 163.367
R1432 B.n307 B.n184 163.367
R1433 B.n308 B.n307 163.367
R1434 B.n309 B.n308 163.367
R1435 B.n309 B.n182 163.367
R1436 B.n313 B.n182 163.367
R1437 B.n314 B.n313 163.367
R1438 B.n315 B.n314 163.367
R1439 B.n315 B.n180 163.367
R1440 B.n319 B.n180 163.367
R1441 B.n320 B.n319 163.367
R1442 B.n321 B.n320 163.367
R1443 B.n321 B.n178 163.367
R1444 B.n325 B.n178 163.367
R1445 B.n326 B.n325 163.367
R1446 B.n327 B.n326 163.367
R1447 B.n327 B.n176 163.367
R1448 B.n331 B.n176 163.367
R1449 B.n332 B.n331 163.367
R1450 B.n333 B.n332 163.367
R1451 B.n333 B.n174 163.367
R1452 B.n337 B.n174 163.367
R1453 B.n338 B.n337 163.367
R1454 B.n339 B.n338 163.367
R1455 B.n339 B.n172 163.367
R1456 B.n343 B.n172 163.367
R1457 B.n344 B.n343 163.367
R1458 B.n345 B.n344 163.367
R1459 B.n345 B.n170 163.367
R1460 B.n349 B.n170 163.367
R1461 B.n350 B.n349 163.367
R1462 B.n351 B.n350 163.367
R1463 B.n351 B.n168 163.367
R1464 B.n355 B.n168 163.367
R1465 B.n356 B.n355 163.367
R1466 B.n357 B.n356 163.367
R1467 B.n357 B.n164 163.367
R1468 B.n362 B.n164 163.367
R1469 B.n363 B.n362 163.367
R1470 B.n364 B.n363 163.367
R1471 B.n364 B.n162 163.367
R1472 B.n368 B.n162 163.367
R1473 B.n369 B.n368 163.367
R1474 B.n370 B.n369 163.367
R1475 B.n370 B.n158 163.367
R1476 B.n375 B.n158 163.367
R1477 B.n376 B.n375 163.367
R1478 B.n377 B.n376 163.367
R1479 B.n377 B.n156 163.367
R1480 B.n381 B.n156 163.367
R1481 B.n382 B.n381 163.367
R1482 B.n383 B.n382 163.367
R1483 B.n383 B.n154 163.367
R1484 B.n387 B.n154 163.367
R1485 B.n388 B.n387 163.367
R1486 B.n389 B.n388 163.367
R1487 B.n389 B.n152 163.367
R1488 B.n393 B.n152 163.367
R1489 B.n394 B.n393 163.367
R1490 B.n395 B.n394 163.367
R1491 B.n395 B.n150 163.367
R1492 B.n399 B.n150 163.367
R1493 B.n400 B.n399 163.367
R1494 B.n401 B.n400 163.367
R1495 B.n401 B.n148 163.367
R1496 B.n405 B.n148 163.367
R1497 B.n406 B.n405 163.367
R1498 B.n407 B.n406 163.367
R1499 B.n407 B.n146 163.367
R1500 B.n411 B.n146 163.367
R1501 B.n412 B.n411 163.367
R1502 B.n413 B.n412 163.367
R1503 B.n413 B.n144 163.367
R1504 B.n417 B.n144 163.367
R1505 B.n418 B.n417 163.367
R1506 B.n419 B.n418 163.367
R1507 B.n419 B.n142 163.367
R1508 B.n423 B.n142 163.367
R1509 B.n424 B.n423 163.367
R1510 B.n425 B.n424 163.367
R1511 B.n425 B.n140 163.367
R1512 B.n429 B.n140 163.367
R1513 B.n430 B.n429 163.367
R1514 B.n431 B.n430 163.367
R1515 B.n431 B.n138 163.367
R1516 B.n435 B.n138 163.367
R1517 B.n436 B.n435 163.367
R1518 B.n437 B.n436 163.367
R1519 B.n437 B.n136 163.367
R1520 B.n441 B.n136 163.367
R1521 B.n442 B.n441 163.367
R1522 B.n598 B.n597 163.367
R1523 B.n597 B.n84 163.367
R1524 B.n593 B.n84 163.367
R1525 B.n593 B.n592 163.367
R1526 B.n592 B.n591 163.367
R1527 B.n591 B.n86 163.367
R1528 B.n587 B.n86 163.367
R1529 B.n587 B.n586 163.367
R1530 B.n586 B.n585 163.367
R1531 B.n585 B.n88 163.367
R1532 B.n581 B.n88 163.367
R1533 B.n581 B.n580 163.367
R1534 B.n580 B.n579 163.367
R1535 B.n579 B.n90 163.367
R1536 B.n575 B.n90 163.367
R1537 B.n575 B.n574 163.367
R1538 B.n574 B.n573 163.367
R1539 B.n573 B.n92 163.367
R1540 B.n569 B.n92 163.367
R1541 B.n569 B.n568 163.367
R1542 B.n568 B.n567 163.367
R1543 B.n567 B.n94 163.367
R1544 B.n563 B.n94 163.367
R1545 B.n563 B.n562 163.367
R1546 B.n562 B.n561 163.367
R1547 B.n561 B.n96 163.367
R1548 B.n557 B.n96 163.367
R1549 B.n557 B.n556 163.367
R1550 B.n556 B.n555 163.367
R1551 B.n555 B.n98 163.367
R1552 B.n551 B.n98 163.367
R1553 B.n551 B.n550 163.367
R1554 B.n550 B.n549 163.367
R1555 B.n549 B.n100 163.367
R1556 B.n545 B.n100 163.367
R1557 B.n545 B.n544 163.367
R1558 B.n544 B.n543 163.367
R1559 B.n543 B.n102 163.367
R1560 B.n539 B.n102 163.367
R1561 B.n539 B.n538 163.367
R1562 B.n538 B.n537 163.367
R1563 B.n537 B.n104 163.367
R1564 B.n533 B.n104 163.367
R1565 B.n533 B.n532 163.367
R1566 B.n532 B.n531 163.367
R1567 B.n531 B.n106 163.367
R1568 B.n527 B.n106 163.367
R1569 B.n527 B.n526 163.367
R1570 B.n526 B.n525 163.367
R1571 B.n525 B.n108 163.367
R1572 B.n521 B.n108 163.367
R1573 B.n521 B.n520 163.367
R1574 B.n520 B.n519 163.367
R1575 B.n519 B.n110 163.367
R1576 B.n515 B.n110 163.367
R1577 B.n515 B.n514 163.367
R1578 B.n514 B.n513 163.367
R1579 B.n513 B.n112 163.367
R1580 B.n509 B.n112 163.367
R1581 B.n509 B.n508 163.367
R1582 B.n508 B.n507 163.367
R1583 B.n507 B.n114 163.367
R1584 B.n503 B.n114 163.367
R1585 B.n503 B.n502 163.367
R1586 B.n502 B.n501 163.367
R1587 B.n501 B.n116 163.367
R1588 B.n497 B.n116 163.367
R1589 B.n497 B.n496 163.367
R1590 B.n496 B.n495 163.367
R1591 B.n495 B.n118 163.367
R1592 B.n491 B.n118 163.367
R1593 B.n491 B.n490 163.367
R1594 B.n490 B.n489 163.367
R1595 B.n489 B.n120 163.367
R1596 B.n485 B.n120 163.367
R1597 B.n485 B.n484 163.367
R1598 B.n484 B.n483 163.367
R1599 B.n483 B.n122 163.367
R1600 B.n479 B.n122 163.367
R1601 B.n479 B.n478 163.367
R1602 B.n478 B.n477 163.367
R1603 B.n477 B.n124 163.367
R1604 B.n473 B.n124 163.367
R1605 B.n473 B.n472 163.367
R1606 B.n472 B.n471 163.367
R1607 B.n471 B.n126 163.367
R1608 B.n467 B.n126 163.367
R1609 B.n467 B.n466 163.367
R1610 B.n466 B.n465 163.367
R1611 B.n465 B.n128 163.367
R1612 B.n461 B.n128 163.367
R1613 B.n461 B.n460 163.367
R1614 B.n460 B.n459 163.367
R1615 B.n459 B.n130 163.367
R1616 B.n455 B.n130 163.367
R1617 B.n455 B.n454 163.367
R1618 B.n454 B.n453 163.367
R1619 B.n453 B.n132 163.367
R1620 B.n449 B.n132 163.367
R1621 B.n449 B.n448 163.367
R1622 B.n448 B.n447 163.367
R1623 B.n447 B.n134 163.367
R1624 B.n443 B.n134 163.367
R1625 B.n750 B.n749 163.367
R1626 B.n749 B.n748 163.367
R1627 B.n748 B.n29 163.367
R1628 B.n744 B.n29 163.367
R1629 B.n744 B.n743 163.367
R1630 B.n743 B.n742 163.367
R1631 B.n742 B.n31 163.367
R1632 B.n738 B.n31 163.367
R1633 B.n738 B.n737 163.367
R1634 B.n737 B.n736 163.367
R1635 B.n736 B.n33 163.367
R1636 B.n732 B.n33 163.367
R1637 B.n732 B.n731 163.367
R1638 B.n731 B.n730 163.367
R1639 B.n730 B.n35 163.367
R1640 B.n726 B.n35 163.367
R1641 B.n726 B.n725 163.367
R1642 B.n725 B.n724 163.367
R1643 B.n724 B.n37 163.367
R1644 B.n720 B.n37 163.367
R1645 B.n720 B.n719 163.367
R1646 B.n719 B.n718 163.367
R1647 B.n718 B.n39 163.367
R1648 B.n714 B.n39 163.367
R1649 B.n714 B.n713 163.367
R1650 B.n713 B.n712 163.367
R1651 B.n712 B.n41 163.367
R1652 B.n708 B.n41 163.367
R1653 B.n708 B.n707 163.367
R1654 B.n707 B.n706 163.367
R1655 B.n706 B.n43 163.367
R1656 B.n702 B.n43 163.367
R1657 B.n702 B.n701 163.367
R1658 B.n701 B.n700 163.367
R1659 B.n700 B.n45 163.367
R1660 B.n696 B.n45 163.367
R1661 B.n696 B.n695 163.367
R1662 B.n695 B.n694 163.367
R1663 B.n694 B.n47 163.367
R1664 B.n690 B.n47 163.367
R1665 B.n690 B.n689 163.367
R1666 B.n689 B.n688 163.367
R1667 B.n688 B.n49 163.367
R1668 B.n684 B.n49 163.367
R1669 B.n684 B.n683 163.367
R1670 B.n683 B.n682 163.367
R1671 B.n682 B.n51 163.367
R1672 B.n678 B.n51 163.367
R1673 B.n678 B.n677 163.367
R1674 B.n677 B.n676 163.367
R1675 B.n676 B.n56 163.367
R1676 B.n672 B.n56 163.367
R1677 B.n672 B.n671 163.367
R1678 B.n671 B.n670 163.367
R1679 B.n670 B.n58 163.367
R1680 B.n665 B.n58 163.367
R1681 B.n665 B.n664 163.367
R1682 B.n664 B.n663 163.367
R1683 B.n663 B.n62 163.367
R1684 B.n659 B.n62 163.367
R1685 B.n659 B.n658 163.367
R1686 B.n658 B.n657 163.367
R1687 B.n657 B.n64 163.367
R1688 B.n653 B.n64 163.367
R1689 B.n653 B.n652 163.367
R1690 B.n652 B.n651 163.367
R1691 B.n651 B.n66 163.367
R1692 B.n647 B.n66 163.367
R1693 B.n647 B.n646 163.367
R1694 B.n646 B.n645 163.367
R1695 B.n645 B.n68 163.367
R1696 B.n641 B.n68 163.367
R1697 B.n641 B.n640 163.367
R1698 B.n640 B.n639 163.367
R1699 B.n639 B.n70 163.367
R1700 B.n635 B.n70 163.367
R1701 B.n635 B.n634 163.367
R1702 B.n634 B.n633 163.367
R1703 B.n633 B.n72 163.367
R1704 B.n629 B.n72 163.367
R1705 B.n629 B.n628 163.367
R1706 B.n628 B.n627 163.367
R1707 B.n627 B.n74 163.367
R1708 B.n623 B.n74 163.367
R1709 B.n623 B.n622 163.367
R1710 B.n622 B.n621 163.367
R1711 B.n621 B.n76 163.367
R1712 B.n617 B.n76 163.367
R1713 B.n617 B.n616 163.367
R1714 B.n616 B.n615 163.367
R1715 B.n615 B.n78 163.367
R1716 B.n611 B.n78 163.367
R1717 B.n611 B.n610 163.367
R1718 B.n610 B.n609 163.367
R1719 B.n609 B.n80 163.367
R1720 B.n605 B.n80 163.367
R1721 B.n605 B.n604 163.367
R1722 B.n604 B.n603 163.367
R1723 B.n603 B.n82 163.367
R1724 B.n599 B.n82 163.367
R1725 B.n754 B.n27 163.367
R1726 B.n755 B.n754 163.367
R1727 B.n756 B.n755 163.367
R1728 B.n756 B.n25 163.367
R1729 B.n760 B.n25 163.367
R1730 B.n761 B.n760 163.367
R1731 B.n762 B.n761 163.367
R1732 B.n762 B.n23 163.367
R1733 B.n766 B.n23 163.367
R1734 B.n767 B.n766 163.367
R1735 B.n768 B.n767 163.367
R1736 B.n768 B.n21 163.367
R1737 B.n772 B.n21 163.367
R1738 B.n773 B.n772 163.367
R1739 B.n774 B.n773 163.367
R1740 B.n774 B.n19 163.367
R1741 B.n778 B.n19 163.367
R1742 B.n779 B.n778 163.367
R1743 B.n780 B.n779 163.367
R1744 B.n780 B.n17 163.367
R1745 B.n784 B.n17 163.367
R1746 B.n785 B.n784 163.367
R1747 B.n786 B.n785 163.367
R1748 B.n786 B.n15 163.367
R1749 B.n790 B.n15 163.367
R1750 B.n791 B.n790 163.367
R1751 B.n792 B.n791 163.367
R1752 B.n792 B.n13 163.367
R1753 B.n796 B.n13 163.367
R1754 B.n797 B.n796 163.367
R1755 B.n798 B.n797 163.367
R1756 B.n798 B.n11 163.367
R1757 B.n802 B.n11 163.367
R1758 B.n803 B.n802 163.367
R1759 B.n804 B.n803 163.367
R1760 B.n804 B.n9 163.367
R1761 B.n808 B.n9 163.367
R1762 B.n809 B.n808 163.367
R1763 B.n810 B.n809 163.367
R1764 B.n810 B.n7 163.367
R1765 B.n814 B.n7 163.367
R1766 B.n815 B.n814 163.367
R1767 B.n816 B.n815 163.367
R1768 B.n816 B.n5 163.367
R1769 B.n820 B.n5 163.367
R1770 B.n821 B.n820 163.367
R1771 B.n822 B.n821 163.367
R1772 B.n822 B.n3 163.367
R1773 B.n826 B.n3 163.367
R1774 B.n827 B.n826 163.367
R1775 B.n214 B.n2 163.367
R1776 B.n217 B.n214 163.367
R1777 B.n218 B.n217 163.367
R1778 B.n219 B.n218 163.367
R1779 B.n219 B.n212 163.367
R1780 B.n223 B.n212 163.367
R1781 B.n224 B.n223 163.367
R1782 B.n225 B.n224 163.367
R1783 B.n225 B.n210 163.367
R1784 B.n229 B.n210 163.367
R1785 B.n230 B.n229 163.367
R1786 B.n231 B.n230 163.367
R1787 B.n231 B.n208 163.367
R1788 B.n235 B.n208 163.367
R1789 B.n236 B.n235 163.367
R1790 B.n237 B.n236 163.367
R1791 B.n237 B.n206 163.367
R1792 B.n241 B.n206 163.367
R1793 B.n242 B.n241 163.367
R1794 B.n243 B.n242 163.367
R1795 B.n243 B.n204 163.367
R1796 B.n247 B.n204 163.367
R1797 B.n248 B.n247 163.367
R1798 B.n249 B.n248 163.367
R1799 B.n249 B.n202 163.367
R1800 B.n253 B.n202 163.367
R1801 B.n254 B.n253 163.367
R1802 B.n255 B.n254 163.367
R1803 B.n255 B.n200 163.367
R1804 B.n259 B.n200 163.367
R1805 B.n260 B.n259 163.367
R1806 B.n261 B.n260 163.367
R1807 B.n261 B.n198 163.367
R1808 B.n265 B.n198 163.367
R1809 B.n266 B.n265 163.367
R1810 B.n267 B.n266 163.367
R1811 B.n267 B.n196 163.367
R1812 B.n271 B.n196 163.367
R1813 B.n272 B.n271 163.367
R1814 B.n273 B.n272 163.367
R1815 B.n273 B.n194 163.367
R1816 B.n277 B.n194 163.367
R1817 B.n278 B.n277 163.367
R1818 B.n279 B.n278 163.367
R1819 B.n279 B.n192 163.367
R1820 B.n283 B.n192 163.367
R1821 B.n284 B.n283 163.367
R1822 B.n285 B.n284 163.367
R1823 B.n285 B.n190 163.367
R1824 B.n289 B.n190 163.367
R1825 B.n359 B.n166 59.5399
R1826 B.n373 B.n160 59.5399
R1827 B.n668 B.n60 59.5399
R1828 B.n54 B.n53 59.5399
R1829 B.n166 B.n165 57.4066
R1830 B.n160 B.n159 57.4066
R1831 B.n60 B.n59 57.4066
R1832 B.n53 B.n52 57.4066
R1833 B.n752 B.n751 33.2493
R1834 B.n600 B.n83 33.2493
R1835 B.n444 B.n135 33.2493
R1836 B.n288 B.n189 33.2493
R1837 B B.n829 18.0485
R1838 B.n753 B.n752 10.6151
R1839 B.n753 B.n26 10.6151
R1840 B.n757 B.n26 10.6151
R1841 B.n758 B.n757 10.6151
R1842 B.n759 B.n758 10.6151
R1843 B.n759 B.n24 10.6151
R1844 B.n763 B.n24 10.6151
R1845 B.n764 B.n763 10.6151
R1846 B.n765 B.n764 10.6151
R1847 B.n765 B.n22 10.6151
R1848 B.n769 B.n22 10.6151
R1849 B.n770 B.n769 10.6151
R1850 B.n771 B.n770 10.6151
R1851 B.n771 B.n20 10.6151
R1852 B.n775 B.n20 10.6151
R1853 B.n776 B.n775 10.6151
R1854 B.n777 B.n776 10.6151
R1855 B.n777 B.n18 10.6151
R1856 B.n781 B.n18 10.6151
R1857 B.n782 B.n781 10.6151
R1858 B.n783 B.n782 10.6151
R1859 B.n783 B.n16 10.6151
R1860 B.n787 B.n16 10.6151
R1861 B.n788 B.n787 10.6151
R1862 B.n789 B.n788 10.6151
R1863 B.n789 B.n14 10.6151
R1864 B.n793 B.n14 10.6151
R1865 B.n794 B.n793 10.6151
R1866 B.n795 B.n794 10.6151
R1867 B.n795 B.n12 10.6151
R1868 B.n799 B.n12 10.6151
R1869 B.n800 B.n799 10.6151
R1870 B.n801 B.n800 10.6151
R1871 B.n801 B.n10 10.6151
R1872 B.n805 B.n10 10.6151
R1873 B.n806 B.n805 10.6151
R1874 B.n807 B.n806 10.6151
R1875 B.n807 B.n8 10.6151
R1876 B.n811 B.n8 10.6151
R1877 B.n812 B.n811 10.6151
R1878 B.n813 B.n812 10.6151
R1879 B.n813 B.n6 10.6151
R1880 B.n817 B.n6 10.6151
R1881 B.n818 B.n817 10.6151
R1882 B.n819 B.n818 10.6151
R1883 B.n819 B.n4 10.6151
R1884 B.n823 B.n4 10.6151
R1885 B.n824 B.n823 10.6151
R1886 B.n825 B.n824 10.6151
R1887 B.n825 B.n0 10.6151
R1888 B.n751 B.n28 10.6151
R1889 B.n747 B.n28 10.6151
R1890 B.n747 B.n746 10.6151
R1891 B.n746 B.n745 10.6151
R1892 B.n745 B.n30 10.6151
R1893 B.n741 B.n30 10.6151
R1894 B.n741 B.n740 10.6151
R1895 B.n740 B.n739 10.6151
R1896 B.n739 B.n32 10.6151
R1897 B.n735 B.n32 10.6151
R1898 B.n735 B.n734 10.6151
R1899 B.n734 B.n733 10.6151
R1900 B.n733 B.n34 10.6151
R1901 B.n729 B.n34 10.6151
R1902 B.n729 B.n728 10.6151
R1903 B.n728 B.n727 10.6151
R1904 B.n727 B.n36 10.6151
R1905 B.n723 B.n36 10.6151
R1906 B.n723 B.n722 10.6151
R1907 B.n722 B.n721 10.6151
R1908 B.n721 B.n38 10.6151
R1909 B.n717 B.n38 10.6151
R1910 B.n717 B.n716 10.6151
R1911 B.n716 B.n715 10.6151
R1912 B.n715 B.n40 10.6151
R1913 B.n711 B.n40 10.6151
R1914 B.n711 B.n710 10.6151
R1915 B.n710 B.n709 10.6151
R1916 B.n709 B.n42 10.6151
R1917 B.n705 B.n42 10.6151
R1918 B.n705 B.n704 10.6151
R1919 B.n704 B.n703 10.6151
R1920 B.n703 B.n44 10.6151
R1921 B.n699 B.n44 10.6151
R1922 B.n699 B.n698 10.6151
R1923 B.n698 B.n697 10.6151
R1924 B.n697 B.n46 10.6151
R1925 B.n693 B.n46 10.6151
R1926 B.n693 B.n692 10.6151
R1927 B.n692 B.n691 10.6151
R1928 B.n691 B.n48 10.6151
R1929 B.n687 B.n48 10.6151
R1930 B.n687 B.n686 10.6151
R1931 B.n686 B.n685 10.6151
R1932 B.n685 B.n50 10.6151
R1933 B.n681 B.n680 10.6151
R1934 B.n680 B.n679 10.6151
R1935 B.n679 B.n55 10.6151
R1936 B.n675 B.n55 10.6151
R1937 B.n675 B.n674 10.6151
R1938 B.n674 B.n673 10.6151
R1939 B.n673 B.n57 10.6151
R1940 B.n669 B.n57 10.6151
R1941 B.n667 B.n666 10.6151
R1942 B.n666 B.n61 10.6151
R1943 B.n662 B.n61 10.6151
R1944 B.n662 B.n661 10.6151
R1945 B.n661 B.n660 10.6151
R1946 B.n660 B.n63 10.6151
R1947 B.n656 B.n63 10.6151
R1948 B.n656 B.n655 10.6151
R1949 B.n655 B.n654 10.6151
R1950 B.n654 B.n65 10.6151
R1951 B.n650 B.n65 10.6151
R1952 B.n650 B.n649 10.6151
R1953 B.n649 B.n648 10.6151
R1954 B.n648 B.n67 10.6151
R1955 B.n644 B.n67 10.6151
R1956 B.n644 B.n643 10.6151
R1957 B.n643 B.n642 10.6151
R1958 B.n642 B.n69 10.6151
R1959 B.n638 B.n69 10.6151
R1960 B.n638 B.n637 10.6151
R1961 B.n637 B.n636 10.6151
R1962 B.n636 B.n71 10.6151
R1963 B.n632 B.n71 10.6151
R1964 B.n632 B.n631 10.6151
R1965 B.n631 B.n630 10.6151
R1966 B.n630 B.n73 10.6151
R1967 B.n626 B.n73 10.6151
R1968 B.n626 B.n625 10.6151
R1969 B.n625 B.n624 10.6151
R1970 B.n624 B.n75 10.6151
R1971 B.n620 B.n75 10.6151
R1972 B.n620 B.n619 10.6151
R1973 B.n619 B.n618 10.6151
R1974 B.n618 B.n77 10.6151
R1975 B.n614 B.n77 10.6151
R1976 B.n614 B.n613 10.6151
R1977 B.n613 B.n612 10.6151
R1978 B.n612 B.n79 10.6151
R1979 B.n608 B.n79 10.6151
R1980 B.n608 B.n607 10.6151
R1981 B.n607 B.n606 10.6151
R1982 B.n606 B.n81 10.6151
R1983 B.n602 B.n81 10.6151
R1984 B.n602 B.n601 10.6151
R1985 B.n601 B.n600 10.6151
R1986 B.n596 B.n83 10.6151
R1987 B.n596 B.n595 10.6151
R1988 B.n595 B.n594 10.6151
R1989 B.n594 B.n85 10.6151
R1990 B.n590 B.n85 10.6151
R1991 B.n590 B.n589 10.6151
R1992 B.n589 B.n588 10.6151
R1993 B.n588 B.n87 10.6151
R1994 B.n584 B.n87 10.6151
R1995 B.n584 B.n583 10.6151
R1996 B.n583 B.n582 10.6151
R1997 B.n582 B.n89 10.6151
R1998 B.n578 B.n89 10.6151
R1999 B.n578 B.n577 10.6151
R2000 B.n577 B.n576 10.6151
R2001 B.n576 B.n91 10.6151
R2002 B.n572 B.n91 10.6151
R2003 B.n572 B.n571 10.6151
R2004 B.n571 B.n570 10.6151
R2005 B.n570 B.n93 10.6151
R2006 B.n566 B.n93 10.6151
R2007 B.n566 B.n565 10.6151
R2008 B.n565 B.n564 10.6151
R2009 B.n564 B.n95 10.6151
R2010 B.n560 B.n95 10.6151
R2011 B.n560 B.n559 10.6151
R2012 B.n559 B.n558 10.6151
R2013 B.n558 B.n97 10.6151
R2014 B.n554 B.n97 10.6151
R2015 B.n554 B.n553 10.6151
R2016 B.n553 B.n552 10.6151
R2017 B.n552 B.n99 10.6151
R2018 B.n548 B.n99 10.6151
R2019 B.n548 B.n547 10.6151
R2020 B.n547 B.n546 10.6151
R2021 B.n546 B.n101 10.6151
R2022 B.n542 B.n101 10.6151
R2023 B.n542 B.n541 10.6151
R2024 B.n541 B.n540 10.6151
R2025 B.n540 B.n103 10.6151
R2026 B.n536 B.n103 10.6151
R2027 B.n536 B.n535 10.6151
R2028 B.n535 B.n534 10.6151
R2029 B.n534 B.n105 10.6151
R2030 B.n530 B.n105 10.6151
R2031 B.n530 B.n529 10.6151
R2032 B.n529 B.n528 10.6151
R2033 B.n528 B.n107 10.6151
R2034 B.n524 B.n107 10.6151
R2035 B.n524 B.n523 10.6151
R2036 B.n523 B.n522 10.6151
R2037 B.n522 B.n109 10.6151
R2038 B.n518 B.n109 10.6151
R2039 B.n518 B.n517 10.6151
R2040 B.n517 B.n516 10.6151
R2041 B.n516 B.n111 10.6151
R2042 B.n512 B.n111 10.6151
R2043 B.n512 B.n511 10.6151
R2044 B.n511 B.n510 10.6151
R2045 B.n510 B.n113 10.6151
R2046 B.n506 B.n113 10.6151
R2047 B.n506 B.n505 10.6151
R2048 B.n505 B.n504 10.6151
R2049 B.n504 B.n115 10.6151
R2050 B.n500 B.n115 10.6151
R2051 B.n500 B.n499 10.6151
R2052 B.n499 B.n498 10.6151
R2053 B.n498 B.n117 10.6151
R2054 B.n494 B.n117 10.6151
R2055 B.n494 B.n493 10.6151
R2056 B.n493 B.n492 10.6151
R2057 B.n492 B.n119 10.6151
R2058 B.n488 B.n119 10.6151
R2059 B.n488 B.n487 10.6151
R2060 B.n487 B.n486 10.6151
R2061 B.n486 B.n121 10.6151
R2062 B.n482 B.n121 10.6151
R2063 B.n482 B.n481 10.6151
R2064 B.n481 B.n480 10.6151
R2065 B.n480 B.n123 10.6151
R2066 B.n476 B.n123 10.6151
R2067 B.n476 B.n475 10.6151
R2068 B.n475 B.n474 10.6151
R2069 B.n474 B.n125 10.6151
R2070 B.n470 B.n125 10.6151
R2071 B.n470 B.n469 10.6151
R2072 B.n469 B.n468 10.6151
R2073 B.n468 B.n127 10.6151
R2074 B.n464 B.n127 10.6151
R2075 B.n464 B.n463 10.6151
R2076 B.n463 B.n462 10.6151
R2077 B.n462 B.n129 10.6151
R2078 B.n458 B.n129 10.6151
R2079 B.n458 B.n457 10.6151
R2080 B.n457 B.n456 10.6151
R2081 B.n456 B.n131 10.6151
R2082 B.n452 B.n131 10.6151
R2083 B.n452 B.n451 10.6151
R2084 B.n451 B.n450 10.6151
R2085 B.n450 B.n133 10.6151
R2086 B.n446 B.n133 10.6151
R2087 B.n446 B.n445 10.6151
R2088 B.n445 B.n444 10.6151
R2089 B.n215 B.n1 10.6151
R2090 B.n216 B.n215 10.6151
R2091 B.n216 B.n213 10.6151
R2092 B.n220 B.n213 10.6151
R2093 B.n221 B.n220 10.6151
R2094 B.n222 B.n221 10.6151
R2095 B.n222 B.n211 10.6151
R2096 B.n226 B.n211 10.6151
R2097 B.n227 B.n226 10.6151
R2098 B.n228 B.n227 10.6151
R2099 B.n228 B.n209 10.6151
R2100 B.n232 B.n209 10.6151
R2101 B.n233 B.n232 10.6151
R2102 B.n234 B.n233 10.6151
R2103 B.n234 B.n207 10.6151
R2104 B.n238 B.n207 10.6151
R2105 B.n239 B.n238 10.6151
R2106 B.n240 B.n239 10.6151
R2107 B.n240 B.n205 10.6151
R2108 B.n244 B.n205 10.6151
R2109 B.n245 B.n244 10.6151
R2110 B.n246 B.n245 10.6151
R2111 B.n246 B.n203 10.6151
R2112 B.n250 B.n203 10.6151
R2113 B.n251 B.n250 10.6151
R2114 B.n252 B.n251 10.6151
R2115 B.n252 B.n201 10.6151
R2116 B.n256 B.n201 10.6151
R2117 B.n257 B.n256 10.6151
R2118 B.n258 B.n257 10.6151
R2119 B.n258 B.n199 10.6151
R2120 B.n262 B.n199 10.6151
R2121 B.n263 B.n262 10.6151
R2122 B.n264 B.n263 10.6151
R2123 B.n264 B.n197 10.6151
R2124 B.n268 B.n197 10.6151
R2125 B.n269 B.n268 10.6151
R2126 B.n270 B.n269 10.6151
R2127 B.n270 B.n195 10.6151
R2128 B.n274 B.n195 10.6151
R2129 B.n275 B.n274 10.6151
R2130 B.n276 B.n275 10.6151
R2131 B.n276 B.n193 10.6151
R2132 B.n280 B.n193 10.6151
R2133 B.n281 B.n280 10.6151
R2134 B.n282 B.n281 10.6151
R2135 B.n282 B.n191 10.6151
R2136 B.n286 B.n191 10.6151
R2137 B.n287 B.n286 10.6151
R2138 B.n288 B.n287 10.6151
R2139 B.n292 B.n189 10.6151
R2140 B.n293 B.n292 10.6151
R2141 B.n294 B.n293 10.6151
R2142 B.n294 B.n187 10.6151
R2143 B.n298 B.n187 10.6151
R2144 B.n299 B.n298 10.6151
R2145 B.n300 B.n299 10.6151
R2146 B.n300 B.n185 10.6151
R2147 B.n304 B.n185 10.6151
R2148 B.n305 B.n304 10.6151
R2149 B.n306 B.n305 10.6151
R2150 B.n306 B.n183 10.6151
R2151 B.n310 B.n183 10.6151
R2152 B.n311 B.n310 10.6151
R2153 B.n312 B.n311 10.6151
R2154 B.n312 B.n181 10.6151
R2155 B.n316 B.n181 10.6151
R2156 B.n317 B.n316 10.6151
R2157 B.n318 B.n317 10.6151
R2158 B.n318 B.n179 10.6151
R2159 B.n322 B.n179 10.6151
R2160 B.n323 B.n322 10.6151
R2161 B.n324 B.n323 10.6151
R2162 B.n324 B.n177 10.6151
R2163 B.n328 B.n177 10.6151
R2164 B.n329 B.n328 10.6151
R2165 B.n330 B.n329 10.6151
R2166 B.n330 B.n175 10.6151
R2167 B.n334 B.n175 10.6151
R2168 B.n335 B.n334 10.6151
R2169 B.n336 B.n335 10.6151
R2170 B.n336 B.n173 10.6151
R2171 B.n340 B.n173 10.6151
R2172 B.n341 B.n340 10.6151
R2173 B.n342 B.n341 10.6151
R2174 B.n342 B.n171 10.6151
R2175 B.n346 B.n171 10.6151
R2176 B.n347 B.n346 10.6151
R2177 B.n348 B.n347 10.6151
R2178 B.n348 B.n169 10.6151
R2179 B.n352 B.n169 10.6151
R2180 B.n353 B.n352 10.6151
R2181 B.n354 B.n353 10.6151
R2182 B.n354 B.n167 10.6151
R2183 B.n358 B.n167 10.6151
R2184 B.n361 B.n360 10.6151
R2185 B.n361 B.n163 10.6151
R2186 B.n365 B.n163 10.6151
R2187 B.n366 B.n365 10.6151
R2188 B.n367 B.n366 10.6151
R2189 B.n367 B.n161 10.6151
R2190 B.n371 B.n161 10.6151
R2191 B.n372 B.n371 10.6151
R2192 B.n374 B.n157 10.6151
R2193 B.n378 B.n157 10.6151
R2194 B.n379 B.n378 10.6151
R2195 B.n380 B.n379 10.6151
R2196 B.n380 B.n155 10.6151
R2197 B.n384 B.n155 10.6151
R2198 B.n385 B.n384 10.6151
R2199 B.n386 B.n385 10.6151
R2200 B.n386 B.n153 10.6151
R2201 B.n390 B.n153 10.6151
R2202 B.n391 B.n390 10.6151
R2203 B.n392 B.n391 10.6151
R2204 B.n392 B.n151 10.6151
R2205 B.n396 B.n151 10.6151
R2206 B.n397 B.n396 10.6151
R2207 B.n398 B.n397 10.6151
R2208 B.n398 B.n149 10.6151
R2209 B.n402 B.n149 10.6151
R2210 B.n403 B.n402 10.6151
R2211 B.n404 B.n403 10.6151
R2212 B.n404 B.n147 10.6151
R2213 B.n408 B.n147 10.6151
R2214 B.n409 B.n408 10.6151
R2215 B.n410 B.n409 10.6151
R2216 B.n410 B.n145 10.6151
R2217 B.n414 B.n145 10.6151
R2218 B.n415 B.n414 10.6151
R2219 B.n416 B.n415 10.6151
R2220 B.n416 B.n143 10.6151
R2221 B.n420 B.n143 10.6151
R2222 B.n421 B.n420 10.6151
R2223 B.n422 B.n421 10.6151
R2224 B.n422 B.n141 10.6151
R2225 B.n426 B.n141 10.6151
R2226 B.n427 B.n426 10.6151
R2227 B.n428 B.n427 10.6151
R2228 B.n428 B.n139 10.6151
R2229 B.n432 B.n139 10.6151
R2230 B.n433 B.n432 10.6151
R2231 B.n434 B.n433 10.6151
R2232 B.n434 B.n137 10.6151
R2233 B.n438 B.n137 10.6151
R2234 B.n439 B.n438 10.6151
R2235 B.n440 B.n439 10.6151
R2236 B.n440 B.n135 10.6151
R2237 B.n829 B.n0 8.11757
R2238 B.n829 B.n1 8.11757
R2239 B.n681 B.n54 6.5566
R2240 B.n669 B.n668 6.5566
R2241 B.n360 B.n359 6.5566
R2242 B.n373 B.n372 6.5566
R2243 B.n54 B.n50 4.05904
R2244 B.n668 B.n667 4.05904
R2245 B.n359 B.n358 4.05904
R2246 B.n374 B.n373 4.05904
R2247 VP.n19 VP.n16 161.3
R2248 VP.n21 VP.n20 161.3
R2249 VP.n22 VP.n15 161.3
R2250 VP.n24 VP.n23 161.3
R2251 VP.n25 VP.n14 161.3
R2252 VP.n27 VP.n26 161.3
R2253 VP.n29 VP.n28 161.3
R2254 VP.n30 VP.n12 161.3
R2255 VP.n32 VP.n31 161.3
R2256 VP.n33 VP.n11 161.3
R2257 VP.n35 VP.n34 161.3
R2258 VP.n36 VP.n10 161.3
R2259 VP.n68 VP.n0 161.3
R2260 VP.n67 VP.n66 161.3
R2261 VP.n65 VP.n1 161.3
R2262 VP.n64 VP.n63 161.3
R2263 VP.n62 VP.n2 161.3
R2264 VP.n61 VP.n60 161.3
R2265 VP.n59 VP.n58 161.3
R2266 VP.n57 VP.n4 161.3
R2267 VP.n56 VP.n55 161.3
R2268 VP.n54 VP.n5 161.3
R2269 VP.n53 VP.n52 161.3
R2270 VP.n51 VP.n6 161.3
R2271 VP.n49 VP.n48 161.3
R2272 VP.n47 VP.n7 161.3
R2273 VP.n46 VP.n45 161.3
R2274 VP.n44 VP.n8 161.3
R2275 VP.n43 VP.n42 161.3
R2276 VP.n41 VP.n9 161.3
R2277 VP.n17 VP.t2 155.923
R2278 VP.n39 VP.t6 122.516
R2279 VP.n50 VP.t3 122.516
R2280 VP.n3 VP.t5 122.516
R2281 VP.n69 VP.t1 122.516
R2282 VP.n37 VP.t4 122.516
R2283 VP.n13 VP.t7 122.516
R2284 VP.n18 VP.t0 122.516
R2285 VP.n40 VP.n39 101.459
R2286 VP.n70 VP.n69 101.459
R2287 VP.n38 VP.n37 101.459
R2288 VP.n18 VP.n17 61.154
R2289 VP.n45 VP.n44 56.5193
R2290 VP.n56 VP.n5 56.5193
R2291 VP.n63 VP.n1 56.5193
R2292 VP.n31 VP.n11 56.5193
R2293 VP.n24 VP.n15 56.5193
R2294 VP.n40 VP.n38 52.0905
R2295 VP.n43 VP.n9 24.4675
R2296 VP.n44 VP.n43 24.4675
R2297 VP.n45 VP.n7 24.4675
R2298 VP.n49 VP.n7 24.4675
R2299 VP.n52 VP.n51 24.4675
R2300 VP.n52 VP.n5 24.4675
R2301 VP.n57 VP.n56 24.4675
R2302 VP.n58 VP.n57 24.4675
R2303 VP.n62 VP.n61 24.4675
R2304 VP.n63 VP.n62 24.4675
R2305 VP.n67 VP.n1 24.4675
R2306 VP.n68 VP.n67 24.4675
R2307 VP.n35 VP.n11 24.4675
R2308 VP.n36 VP.n35 24.4675
R2309 VP.n25 VP.n24 24.4675
R2310 VP.n26 VP.n25 24.4675
R2311 VP.n30 VP.n29 24.4675
R2312 VP.n31 VP.n30 24.4675
R2313 VP.n20 VP.n19 24.4675
R2314 VP.n20 VP.n15 24.4675
R2315 VP.n50 VP.n49 13.2127
R2316 VP.n61 VP.n3 13.2127
R2317 VP.n29 VP.n13 13.2127
R2318 VP.n51 VP.n50 11.2553
R2319 VP.n58 VP.n3 11.2553
R2320 VP.n26 VP.n13 11.2553
R2321 VP.n19 VP.n18 11.2553
R2322 VP.n39 VP.n9 9.29796
R2323 VP.n69 VP.n68 9.29796
R2324 VP.n37 VP.n36 9.29796
R2325 VP.n17 VP.n16 6.89416
R2326 VP.n38 VP.n10 0.278367
R2327 VP.n41 VP.n40 0.278367
R2328 VP.n70 VP.n0 0.278367
R2329 VP.n21 VP.n16 0.189894
R2330 VP.n22 VP.n21 0.189894
R2331 VP.n23 VP.n22 0.189894
R2332 VP.n23 VP.n14 0.189894
R2333 VP.n27 VP.n14 0.189894
R2334 VP.n28 VP.n27 0.189894
R2335 VP.n28 VP.n12 0.189894
R2336 VP.n32 VP.n12 0.189894
R2337 VP.n33 VP.n32 0.189894
R2338 VP.n34 VP.n33 0.189894
R2339 VP.n34 VP.n10 0.189894
R2340 VP.n42 VP.n41 0.189894
R2341 VP.n42 VP.n8 0.189894
R2342 VP.n46 VP.n8 0.189894
R2343 VP.n47 VP.n46 0.189894
R2344 VP.n48 VP.n47 0.189894
R2345 VP.n48 VP.n6 0.189894
R2346 VP.n53 VP.n6 0.189894
R2347 VP.n54 VP.n53 0.189894
R2348 VP.n55 VP.n54 0.189894
R2349 VP.n55 VP.n4 0.189894
R2350 VP.n59 VP.n4 0.189894
R2351 VP.n60 VP.n59 0.189894
R2352 VP.n60 VP.n2 0.189894
R2353 VP.n64 VP.n2 0.189894
R2354 VP.n65 VP.n64 0.189894
R2355 VP.n66 VP.n65 0.189894
R2356 VP.n66 VP.n0 0.189894
R2357 VP VP.n70 0.153454
R2358 VDD1 VDD1.n0 76.5976
R2359 VDD1.n3 VDD1.n2 76.4839
R2360 VDD1.n3 VDD1.n1 76.4839
R2361 VDD1.n5 VDD1.n4 75.2634
R2362 VDD1.n5 VDD1.n3 47.3069
R2363 VDD1.n4 VDD1.t0 2.43169
R2364 VDD1.n4 VDD1.t3 2.43169
R2365 VDD1.n0 VDD1.t5 2.43169
R2366 VDD1.n0 VDD1.t7 2.43169
R2367 VDD1.n2 VDD1.t2 2.43169
R2368 VDD1.n2 VDD1.t6 2.43169
R2369 VDD1.n1 VDD1.t1 2.43169
R2370 VDD1.n1 VDD1.t4 2.43169
R2371 VDD1 VDD1.n5 1.21817
C0 w_n3930_n3642# B 10.5459f
C1 VP VN 7.95178f
C2 VDD1 VDD2 1.79374f
C3 w_n3930_n3642# VN 8.02392f
C4 VDD1 B 1.69434f
C5 VDD1 VN 0.151889f
C6 VDD2 B 1.79131f
C7 VDD2 VN 9.65168f
C8 VP VTAIL 10.0112f
C9 B VN 1.24831f
C10 w_n3930_n3642# VTAIL 4.5243f
C11 VDD1 VTAIL 8.54197f
C12 VDD2 VTAIL 8.59659f
C13 B VTAIL 5.44754f
C14 VN VTAIL 9.99709f
C15 w_n3930_n3642# VP 8.5342f
C16 VDD1 VP 10.0213f
C17 VDD1 w_n3930_n3642# 2.00388f
C18 VDD2 VP 0.52297f
C19 B VP 2.10388f
C20 VDD2 w_n3930_n3642# 2.11985f
C21 VDD2 VSUBS 1.923505f
C22 VDD1 VSUBS 2.56838f
C23 VTAIL VSUBS 1.40244f
C24 VN VSUBS 6.82626f
C25 VP VSUBS 3.666134f
C26 B VSUBS 5.155122f
C27 w_n3930_n3642# VSUBS 0.17586p
C28 VDD1.t5 VSUBS 0.286786f
C29 VDD1.t7 VSUBS 0.286786f
C30 VDD1.n0 VSUBS 2.31582f
C31 VDD1.t1 VSUBS 0.286786f
C32 VDD1.t4 VSUBS 0.286786f
C33 VDD1.n1 VSUBS 2.31443f
C34 VDD1.t2 VSUBS 0.286786f
C35 VDD1.t6 VSUBS 0.286786f
C36 VDD1.n2 VSUBS 2.31443f
C37 VDD1.n3 VSUBS 4.26928f
C38 VDD1.t0 VSUBS 0.286786f
C39 VDD1.t3 VSUBS 0.286786f
C40 VDD1.n4 VSUBS 2.30105f
C41 VDD1.n5 VSUBS 3.63467f
C42 VP.n0 VSUBS 0.040052f
C43 VP.t1 VSUBS 2.91902f
C44 VP.n1 VSUBS 0.047734f
C45 VP.n2 VSUBS 0.030379f
C46 VP.t5 VSUBS 2.91902f
C47 VP.n3 VSUBS 1.02584f
C48 VP.n4 VSUBS 0.030379f
C49 VP.n5 VSUBS 0.044348f
C50 VP.n6 VSUBS 0.030379f
C51 VP.t3 VSUBS 2.91902f
C52 VP.n7 VSUBS 0.056619f
C53 VP.n8 VSUBS 0.030379f
C54 VP.n9 VSUBS 0.039288f
C55 VP.n10 VSUBS 0.040052f
C56 VP.t4 VSUBS 2.91902f
C57 VP.n11 VSUBS 0.047734f
C58 VP.n12 VSUBS 0.030379f
C59 VP.t7 VSUBS 2.91902f
C60 VP.n13 VSUBS 1.02584f
C61 VP.n14 VSUBS 0.030379f
C62 VP.n15 VSUBS 0.044348f
C63 VP.n16 VSUBS 0.29458f
C64 VP.t0 VSUBS 2.91902f
C65 VP.t2 VSUBS 3.17943f
C66 VP.n17 VSUBS 1.08291f
C67 VP.n18 VSUBS 1.11286f
C68 VP.n19 VSUBS 0.041524f
C69 VP.n20 VSUBS 0.056619f
C70 VP.n21 VSUBS 0.030379f
C71 VP.n22 VSUBS 0.030379f
C72 VP.n23 VSUBS 0.030379f
C73 VP.n24 VSUBS 0.044348f
C74 VP.n25 VSUBS 0.056619f
C75 VP.n26 VSUBS 0.041524f
C76 VP.n27 VSUBS 0.030379f
C77 VP.n28 VSUBS 0.030379f
C78 VP.n29 VSUBS 0.043761f
C79 VP.n30 VSUBS 0.056619f
C80 VP.n31 VSUBS 0.040962f
C81 VP.n32 VSUBS 0.030379f
C82 VP.n33 VSUBS 0.030379f
C83 VP.n34 VSUBS 0.030379f
C84 VP.n35 VSUBS 0.056619f
C85 VP.n36 VSUBS 0.039288f
C86 VP.n37 VSUBS 1.12783f
C87 VP.n38 VSUBS 1.7952f
C88 VP.t6 VSUBS 2.91902f
C89 VP.n39 VSUBS 1.12783f
C90 VP.n40 VSUBS 1.81616f
C91 VP.n41 VSUBS 0.040052f
C92 VP.n42 VSUBS 0.030379f
C93 VP.n43 VSUBS 0.056619f
C94 VP.n44 VSUBS 0.047734f
C95 VP.n45 VSUBS 0.040962f
C96 VP.n46 VSUBS 0.030379f
C97 VP.n47 VSUBS 0.030379f
C98 VP.n48 VSUBS 0.030379f
C99 VP.n49 VSUBS 0.043761f
C100 VP.n50 VSUBS 1.02584f
C101 VP.n51 VSUBS 0.041524f
C102 VP.n52 VSUBS 0.056619f
C103 VP.n53 VSUBS 0.030379f
C104 VP.n54 VSUBS 0.030379f
C105 VP.n55 VSUBS 0.030379f
C106 VP.n56 VSUBS 0.044348f
C107 VP.n57 VSUBS 0.056619f
C108 VP.n58 VSUBS 0.041524f
C109 VP.n59 VSUBS 0.030379f
C110 VP.n60 VSUBS 0.030379f
C111 VP.n61 VSUBS 0.043761f
C112 VP.n62 VSUBS 0.056619f
C113 VP.n63 VSUBS 0.040962f
C114 VP.n64 VSUBS 0.030379f
C115 VP.n65 VSUBS 0.030379f
C116 VP.n66 VSUBS 0.030379f
C117 VP.n67 VSUBS 0.056619f
C118 VP.n68 VSUBS 0.039288f
C119 VP.n69 VSUBS 1.12783f
C120 VP.n70 VSUBS 0.050255f
C121 B.n0 VSUBS 0.006464f
C122 B.n1 VSUBS 0.006464f
C123 B.n2 VSUBS 0.00956f
C124 B.n3 VSUBS 0.007326f
C125 B.n4 VSUBS 0.007326f
C126 B.n5 VSUBS 0.007326f
C127 B.n6 VSUBS 0.007326f
C128 B.n7 VSUBS 0.007326f
C129 B.n8 VSUBS 0.007326f
C130 B.n9 VSUBS 0.007326f
C131 B.n10 VSUBS 0.007326f
C132 B.n11 VSUBS 0.007326f
C133 B.n12 VSUBS 0.007326f
C134 B.n13 VSUBS 0.007326f
C135 B.n14 VSUBS 0.007326f
C136 B.n15 VSUBS 0.007326f
C137 B.n16 VSUBS 0.007326f
C138 B.n17 VSUBS 0.007326f
C139 B.n18 VSUBS 0.007326f
C140 B.n19 VSUBS 0.007326f
C141 B.n20 VSUBS 0.007326f
C142 B.n21 VSUBS 0.007326f
C143 B.n22 VSUBS 0.007326f
C144 B.n23 VSUBS 0.007326f
C145 B.n24 VSUBS 0.007326f
C146 B.n25 VSUBS 0.007326f
C147 B.n26 VSUBS 0.007326f
C148 B.n27 VSUBS 0.016795f
C149 B.n28 VSUBS 0.007326f
C150 B.n29 VSUBS 0.007326f
C151 B.n30 VSUBS 0.007326f
C152 B.n31 VSUBS 0.007326f
C153 B.n32 VSUBS 0.007326f
C154 B.n33 VSUBS 0.007326f
C155 B.n34 VSUBS 0.007326f
C156 B.n35 VSUBS 0.007326f
C157 B.n36 VSUBS 0.007326f
C158 B.n37 VSUBS 0.007326f
C159 B.n38 VSUBS 0.007326f
C160 B.n39 VSUBS 0.007326f
C161 B.n40 VSUBS 0.007326f
C162 B.n41 VSUBS 0.007326f
C163 B.n42 VSUBS 0.007326f
C164 B.n43 VSUBS 0.007326f
C165 B.n44 VSUBS 0.007326f
C166 B.n45 VSUBS 0.007326f
C167 B.n46 VSUBS 0.007326f
C168 B.n47 VSUBS 0.007326f
C169 B.n48 VSUBS 0.007326f
C170 B.n49 VSUBS 0.007326f
C171 B.n50 VSUBS 0.005063f
C172 B.n51 VSUBS 0.007326f
C173 B.t10 VSUBS 0.253077f
C174 B.t11 VSUBS 0.287303f
C175 B.t9 VSUBS 1.66611f
C176 B.n52 VSUBS 0.451776f
C177 B.n53 VSUBS 0.283287f
C178 B.n54 VSUBS 0.016973f
C179 B.n55 VSUBS 0.007326f
C180 B.n56 VSUBS 0.007326f
C181 B.n57 VSUBS 0.007326f
C182 B.n58 VSUBS 0.007326f
C183 B.t7 VSUBS 0.25308f
C184 B.t8 VSUBS 0.287306f
C185 B.t6 VSUBS 1.66611f
C186 B.n59 VSUBS 0.451773f
C187 B.n60 VSUBS 0.283284f
C188 B.n61 VSUBS 0.007326f
C189 B.n62 VSUBS 0.007326f
C190 B.n63 VSUBS 0.007326f
C191 B.n64 VSUBS 0.007326f
C192 B.n65 VSUBS 0.007326f
C193 B.n66 VSUBS 0.007326f
C194 B.n67 VSUBS 0.007326f
C195 B.n68 VSUBS 0.007326f
C196 B.n69 VSUBS 0.007326f
C197 B.n70 VSUBS 0.007326f
C198 B.n71 VSUBS 0.007326f
C199 B.n72 VSUBS 0.007326f
C200 B.n73 VSUBS 0.007326f
C201 B.n74 VSUBS 0.007326f
C202 B.n75 VSUBS 0.007326f
C203 B.n76 VSUBS 0.007326f
C204 B.n77 VSUBS 0.007326f
C205 B.n78 VSUBS 0.007326f
C206 B.n79 VSUBS 0.007326f
C207 B.n80 VSUBS 0.007326f
C208 B.n81 VSUBS 0.007326f
C209 B.n82 VSUBS 0.007326f
C210 B.n83 VSUBS 0.016795f
C211 B.n84 VSUBS 0.007326f
C212 B.n85 VSUBS 0.007326f
C213 B.n86 VSUBS 0.007326f
C214 B.n87 VSUBS 0.007326f
C215 B.n88 VSUBS 0.007326f
C216 B.n89 VSUBS 0.007326f
C217 B.n90 VSUBS 0.007326f
C218 B.n91 VSUBS 0.007326f
C219 B.n92 VSUBS 0.007326f
C220 B.n93 VSUBS 0.007326f
C221 B.n94 VSUBS 0.007326f
C222 B.n95 VSUBS 0.007326f
C223 B.n96 VSUBS 0.007326f
C224 B.n97 VSUBS 0.007326f
C225 B.n98 VSUBS 0.007326f
C226 B.n99 VSUBS 0.007326f
C227 B.n100 VSUBS 0.007326f
C228 B.n101 VSUBS 0.007326f
C229 B.n102 VSUBS 0.007326f
C230 B.n103 VSUBS 0.007326f
C231 B.n104 VSUBS 0.007326f
C232 B.n105 VSUBS 0.007326f
C233 B.n106 VSUBS 0.007326f
C234 B.n107 VSUBS 0.007326f
C235 B.n108 VSUBS 0.007326f
C236 B.n109 VSUBS 0.007326f
C237 B.n110 VSUBS 0.007326f
C238 B.n111 VSUBS 0.007326f
C239 B.n112 VSUBS 0.007326f
C240 B.n113 VSUBS 0.007326f
C241 B.n114 VSUBS 0.007326f
C242 B.n115 VSUBS 0.007326f
C243 B.n116 VSUBS 0.007326f
C244 B.n117 VSUBS 0.007326f
C245 B.n118 VSUBS 0.007326f
C246 B.n119 VSUBS 0.007326f
C247 B.n120 VSUBS 0.007326f
C248 B.n121 VSUBS 0.007326f
C249 B.n122 VSUBS 0.007326f
C250 B.n123 VSUBS 0.007326f
C251 B.n124 VSUBS 0.007326f
C252 B.n125 VSUBS 0.007326f
C253 B.n126 VSUBS 0.007326f
C254 B.n127 VSUBS 0.007326f
C255 B.n128 VSUBS 0.007326f
C256 B.n129 VSUBS 0.007326f
C257 B.n130 VSUBS 0.007326f
C258 B.n131 VSUBS 0.007326f
C259 B.n132 VSUBS 0.007326f
C260 B.n133 VSUBS 0.007326f
C261 B.n134 VSUBS 0.007326f
C262 B.n135 VSUBS 0.017044f
C263 B.n136 VSUBS 0.007326f
C264 B.n137 VSUBS 0.007326f
C265 B.n138 VSUBS 0.007326f
C266 B.n139 VSUBS 0.007326f
C267 B.n140 VSUBS 0.007326f
C268 B.n141 VSUBS 0.007326f
C269 B.n142 VSUBS 0.007326f
C270 B.n143 VSUBS 0.007326f
C271 B.n144 VSUBS 0.007326f
C272 B.n145 VSUBS 0.007326f
C273 B.n146 VSUBS 0.007326f
C274 B.n147 VSUBS 0.007326f
C275 B.n148 VSUBS 0.007326f
C276 B.n149 VSUBS 0.007326f
C277 B.n150 VSUBS 0.007326f
C278 B.n151 VSUBS 0.007326f
C279 B.n152 VSUBS 0.007326f
C280 B.n153 VSUBS 0.007326f
C281 B.n154 VSUBS 0.007326f
C282 B.n155 VSUBS 0.007326f
C283 B.n156 VSUBS 0.007326f
C284 B.n157 VSUBS 0.007326f
C285 B.n158 VSUBS 0.007326f
C286 B.t2 VSUBS 0.25308f
C287 B.t1 VSUBS 0.287306f
C288 B.t0 VSUBS 1.66611f
C289 B.n159 VSUBS 0.451773f
C290 B.n160 VSUBS 0.283284f
C291 B.n161 VSUBS 0.007326f
C292 B.n162 VSUBS 0.007326f
C293 B.n163 VSUBS 0.007326f
C294 B.n164 VSUBS 0.007326f
C295 B.t5 VSUBS 0.253077f
C296 B.t4 VSUBS 0.287303f
C297 B.t3 VSUBS 1.66611f
C298 B.n165 VSUBS 0.451776f
C299 B.n166 VSUBS 0.283287f
C300 B.n167 VSUBS 0.007326f
C301 B.n168 VSUBS 0.007326f
C302 B.n169 VSUBS 0.007326f
C303 B.n170 VSUBS 0.007326f
C304 B.n171 VSUBS 0.007326f
C305 B.n172 VSUBS 0.007326f
C306 B.n173 VSUBS 0.007326f
C307 B.n174 VSUBS 0.007326f
C308 B.n175 VSUBS 0.007326f
C309 B.n176 VSUBS 0.007326f
C310 B.n177 VSUBS 0.007326f
C311 B.n178 VSUBS 0.007326f
C312 B.n179 VSUBS 0.007326f
C313 B.n180 VSUBS 0.007326f
C314 B.n181 VSUBS 0.007326f
C315 B.n182 VSUBS 0.007326f
C316 B.n183 VSUBS 0.007326f
C317 B.n184 VSUBS 0.007326f
C318 B.n185 VSUBS 0.007326f
C319 B.n186 VSUBS 0.007326f
C320 B.n187 VSUBS 0.007326f
C321 B.n188 VSUBS 0.007326f
C322 B.n189 VSUBS 0.017894f
C323 B.n190 VSUBS 0.007326f
C324 B.n191 VSUBS 0.007326f
C325 B.n192 VSUBS 0.007326f
C326 B.n193 VSUBS 0.007326f
C327 B.n194 VSUBS 0.007326f
C328 B.n195 VSUBS 0.007326f
C329 B.n196 VSUBS 0.007326f
C330 B.n197 VSUBS 0.007326f
C331 B.n198 VSUBS 0.007326f
C332 B.n199 VSUBS 0.007326f
C333 B.n200 VSUBS 0.007326f
C334 B.n201 VSUBS 0.007326f
C335 B.n202 VSUBS 0.007326f
C336 B.n203 VSUBS 0.007326f
C337 B.n204 VSUBS 0.007326f
C338 B.n205 VSUBS 0.007326f
C339 B.n206 VSUBS 0.007326f
C340 B.n207 VSUBS 0.007326f
C341 B.n208 VSUBS 0.007326f
C342 B.n209 VSUBS 0.007326f
C343 B.n210 VSUBS 0.007326f
C344 B.n211 VSUBS 0.007326f
C345 B.n212 VSUBS 0.007326f
C346 B.n213 VSUBS 0.007326f
C347 B.n214 VSUBS 0.007326f
C348 B.n215 VSUBS 0.007326f
C349 B.n216 VSUBS 0.007326f
C350 B.n217 VSUBS 0.007326f
C351 B.n218 VSUBS 0.007326f
C352 B.n219 VSUBS 0.007326f
C353 B.n220 VSUBS 0.007326f
C354 B.n221 VSUBS 0.007326f
C355 B.n222 VSUBS 0.007326f
C356 B.n223 VSUBS 0.007326f
C357 B.n224 VSUBS 0.007326f
C358 B.n225 VSUBS 0.007326f
C359 B.n226 VSUBS 0.007326f
C360 B.n227 VSUBS 0.007326f
C361 B.n228 VSUBS 0.007326f
C362 B.n229 VSUBS 0.007326f
C363 B.n230 VSUBS 0.007326f
C364 B.n231 VSUBS 0.007326f
C365 B.n232 VSUBS 0.007326f
C366 B.n233 VSUBS 0.007326f
C367 B.n234 VSUBS 0.007326f
C368 B.n235 VSUBS 0.007326f
C369 B.n236 VSUBS 0.007326f
C370 B.n237 VSUBS 0.007326f
C371 B.n238 VSUBS 0.007326f
C372 B.n239 VSUBS 0.007326f
C373 B.n240 VSUBS 0.007326f
C374 B.n241 VSUBS 0.007326f
C375 B.n242 VSUBS 0.007326f
C376 B.n243 VSUBS 0.007326f
C377 B.n244 VSUBS 0.007326f
C378 B.n245 VSUBS 0.007326f
C379 B.n246 VSUBS 0.007326f
C380 B.n247 VSUBS 0.007326f
C381 B.n248 VSUBS 0.007326f
C382 B.n249 VSUBS 0.007326f
C383 B.n250 VSUBS 0.007326f
C384 B.n251 VSUBS 0.007326f
C385 B.n252 VSUBS 0.007326f
C386 B.n253 VSUBS 0.007326f
C387 B.n254 VSUBS 0.007326f
C388 B.n255 VSUBS 0.007326f
C389 B.n256 VSUBS 0.007326f
C390 B.n257 VSUBS 0.007326f
C391 B.n258 VSUBS 0.007326f
C392 B.n259 VSUBS 0.007326f
C393 B.n260 VSUBS 0.007326f
C394 B.n261 VSUBS 0.007326f
C395 B.n262 VSUBS 0.007326f
C396 B.n263 VSUBS 0.007326f
C397 B.n264 VSUBS 0.007326f
C398 B.n265 VSUBS 0.007326f
C399 B.n266 VSUBS 0.007326f
C400 B.n267 VSUBS 0.007326f
C401 B.n268 VSUBS 0.007326f
C402 B.n269 VSUBS 0.007326f
C403 B.n270 VSUBS 0.007326f
C404 B.n271 VSUBS 0.007326f
C405 B.n272 VSUBS 0.007326f
C406 B.n273 VSUBS 0.007326f
C407 B.n274 VSUBS 0.007326f
C408 B.n275 VSUBS 0.007326f
C409 B.n276 VSUBS 0.007326f
C410 B.n277 VSUBS 0.007326f
C411 B.n278 VSUBS 0.007326f
C412 B.n279 VSUBS 0.007326f
C413 B.n280 VSUBS 0.007326f
C414 B.n281 VSUBS 0.007326f
C415 B.n282 VSUBS 0.007326f
C416 B.n283 VSUBS 0.007326f
C417 B.n284 VSUBS 0.007326f
C418 B.n285 VSUBS 0.007326f
C419 B.n286 VSUBS 0.007326f
C420 B.n287 VSUBS 0.007326f
C421 B.n288 VSUBS 0.016795f
C422 B.n289 VSUBS 0.016795f
C423 B.n290 VSUBS 0.017894f
C424 B.n291 VSUBS 0.007326f
C425 B.n292 VSUBS 0.007326f
C426 B.n293 VSUBS 0.007326f
C427 B.n294 VSUBS 0.007326f
C428 B.n295 VSUBS 0.007326f
C429 B.n296 VSUBS 0.007326f
C430 B.n297 VSUBS 0.007326f
C431 B.n298 VSUBS 0.007326f
C432 B.n299 VSUBS 0.007326f
C433 B.n300 VSUBS 0.007326f
C434 B.n301 VSUBS 0.007326f
C435 B.n302 VSUBS 0.007326f
C436 B.n303 VSUBS 0.007326f
C437 B.n304 VSUBS 0.007326f
C438 B.n305 VSUBS 0.007326f
C439 B.n306 VSUBS 0.007326f
C440 B.n307 VSUBS 0.007326f
C441 B.n308 VSUBS 0.007326f
C442 B.n309 VSUBS 0.007326f
C443 B.n310 VSUBS 0.007326f
C444 B.n311 VSUBS 0.007326f
C445 B.n312 VSUBS 0.007326f
C446 B.n313 VSUBS 0.007326f
C447 B.n314 VSUBS 0.007326f
C448 B.n315 VSUBS 0.007326f
C449 B.n316 VSUBS 0.007326f
C450 B.n317 VSUBS 0.007326f
C451 B.n318 VSUBS 0.007326f
C452 B.n319 VSUBS 0.007326f
C453 B.n320 VSUBS 0.007326f
C454 B.n321 VSUBS 0.007326f
C455 B.n322 VSUBS 0.007326f
C456 B.n323 VSUBS 0.007326f
C457 B.n324 VSUBS 0.007326f
C458 B.n325 VSUBS 0.007326f
C459 B.n326 VSUBS 0.007326f
C460 B.n327 VSUBS 0.007326f
C461 B.n328 VSUBS 0.007326f
C462 B.n329 VSUBS 0.007326f
C463 B.n330 VSUBS 0.007326f
C464 B.n331 VSUBS 0.007326f
C465 B.n332 VSUBS 0.007326f
C466 B.n333 VSUBS 0.007326f
C467 B.n334 VSUBS 0.007326f
C468 B.n335 VSUBS 0.007326f
C469 B.n336 VSUBS 0.007326f
C470 B.n337 VSUBS 0.007326f
C471 B.n338 VSUBS 0.007326f
C472 B.n339 VSUBS 0.007326f
C473 B.n340 VSUBS 0.007326f
C474 B.n341 VSUBS 0.007326f
C475 B.n342 VSUBS 0.007326f
C476 B.n343 VSUBS 0.007326f
C477 B.n344 VSUBS 0.007326f
C478 B.n345 VSUBS 0.007326f
C479 B.n346 VSUBS 0.007326f
C480 B.n347 VSUBS 0.007326f
C481 B.n348 VSUBS 0.007326f
C482 B.n349 VSUBS 0.007326f
C483 B.n350 VSUBS 0.007326f
C484 B.n351 VSUBS 0.007326f
C485 B.n352 VSUBS 0.007326f
C486 B.n353 VSUBS 0.007326f
C487 B.n354 VSUBS 0.007326f
C488 B.n355 VSUBS 0.007326f
C489 B.n356 VSUBS 0.007326f
C490 B.n357 VSUBS 0.007326f
C491 B.n358 VSUBS 0.005063f
C492 B.n359 VSUBS 0.016973f
C493 B.n360 VSUBS 0.005925f
C494 B.n361 VSUBS 0.007326f
C495 B.n362 VSUBS 0.007326f
C496 B.n363 VSUBS 0.007326f
C497 B.n364 VSUBS 0.007326f
C498 B.n365 VSUBS 0.007326f
C499 B.n366 VSUBS 0.007326f
C500 B.n367 VSUBS 0.007326f
C501 B.n368 VSUBS 0.007326f
C502 B.n369 VSUBS 0.007326f
C503 B.n370 VSUBS 0.007326f
C504 B.n371 VSUBS 0.007326f
C505 B.n372 VSUBS 0.005925f
C506 B.n373 VSUBS 0.016973f
C507 B.n374 VSUBS 0.005063f
C508 B.n375 VSUBS 0.007326f
C509 B.n376 VSUBS 0.007326f
C510 B.n377 VSUBS 0.007326f
C511 B.n378 VSUBS 0.007326f
C512 B.n379 VSUBS 0.007326f
C513 B.n380 VSUBS 0.007326f
C514 B.n381 VSUBS 0.007326f
C515 B.n382 VSUBS 0.007326f
C516 B.n383 VSUBS 0.007326f
C517 B.n384 VSUBS 0.007326f
C518 B.n385 VSUBS 0.007326f
C519 B.n386 VSUBS 0.007326f
C520 B.n387 VSUBS 0.007326f
C521 B.n388 VSUBS 0.007326f
C522 B.n389 VSUBS 0.007326f
C523 B.n390 VSUBS 0.007326f
C524 B.n391 VSUBS 0.007326f
C525 B.n392 VSUBS 0.007326f
C526 B.n393 VSUBS 0.007326f
C527 B.n394 VSUBS 0.007326f
C528 B.n395 VSUBS 0.007326f
C529 B.n396 VSUBS 0.007326f
C530 B.n397 VSUBS 0.007326f
C531 B.n398 VSUBS 0.007326f
C532 B.n399 VSUBS 0.007326f
C533 B.n400 VSUBS 0.007326f
C534 B.n401 VSUBS 0.007326f
C535 B.n402 VSUBS 0.007326f
C536 B.n403 VSUBS 0.007326f
C537 B.n404 VSUBS 0.007326f
C538 B.n405 VSUBS 0.007326f
C539 B.n406 VSUBS 0.007326f
C540 B.n407 VSUBS 0.007326f
C541 B.n408 VSUBS 0.007326f
C542 B.n409 VSUBS 0.007326f
C543 B.n410 VSUBS 0.007326f
C544 B.n411 VSUBS 0.007326f
C545 B.n412 VSUBS 0.007326f
C546 B.n413 VSUBS 0.007326f
C547 B.n414 VSUBS 0.007326f
C548 B.n415 VSUBS 0.007326f
C549 B.n416 VSUBS 0.007326f
C550 B.n417 VSUBS 0.007326f
C551 B.n418 VSUBS 0.007326f
C552 B.n419 VSUBS 0.007326f
C553 B.n420 VSUBS 0.007326f
C554 B.n421 VSUBS 0.007326f
C555 B.n422 VSUBS 0.007326f
C556 B.n423 VSUBS 0.007326f
C557 B.n424 VSUBS 0.007326f
C558 B.n425 VSUBS 0.007326f
C559 B.n426 VSUBS 0.007326f
C560 B.n427 VSUBS 0.007326f
C561 B.n428 VSUBS 0.007326f
C562 B.n429 VSUBS 0.007326f
C563 B.n430 VSUBS 0.007326f
C564 B.n431 VSUBS 0.007326f
C565 B.n432 VSUBS 0.007326f
C566 B.n433 VSUBS 0.007326f
C567 B.n434 VSUBS 0.007326f
C568 B.n435 VSUBS 0.007326f
C569 B.n436 VSUBS 0.007326f
C570 B.n437 VSUBS 0.007326f
C571 B.n438 VSUBS 0.007326f
C572 B.n439 VSUBS 0.007326f
C573 B.n440 VSUBS 0.007326f
C574 B.n441 VSUBS 0.007326f
C575 B.n442 VSUBS 0.017894f
C576 B.n443 VSUBS 0.016795f
C577 B.n444 VSUBS 0.017645f
C578 B.n445 VSUBS 0.007326f
C579 B.n446 VSUBS 0.007326f
C580 B.n447 VSUBS 0.007326f
C581 B.n448 VSUBS 0.007326f
C582 B.n449 VSUBS 0.007326f
C583 B.n450 VSUBS 0.007326f
C584 B.n451 VSUBS 0.007326f
C585 B.n452 VSUBS 0.007326f
C586 B.n453 VSUBS 0.007326f
C587 B.n454 VSUBS 0.007326f
C588 B.n455 VSUBS 0.007326f
C589 B.n456 VSUBS 0.007326f
C590 B.n457 VSUBS 0.007326f
C591 B.n458 VSUBS 0.007326f
C592 B.n459 VSUBS 0.007326f
C593 B.n460 VSUBS 0.007326f
C594 B.n461 VSUBS 0.007326f
C595 B.n462 VSUBS 0.007326f
C596 B.n463 VSUBS 0.007326f
C597 B.n464 VSUBS 0.007326f
C598 B.n465 VSUBS 0.007326f
C599 B.n466 VSUBS 0.007326f
C600 B.n467 VSUBS 0.007326f
C601 B.n468 VSUBS 0.007326f
C602 B.n469 VSUBS 0.007326f
C603 B.n470 VSUBS 0.007326f
C604 B.n471 VSUBS 0.007326f
C605 B.n472 VSUBS 0.007326f
C606 B.n473 VSUBS 0.007326f
C607 B.n474 VSUBS 0.007326f
C608 B.n475 VSUBS 0.007326f
C609 B.n476 VSUBS 0.007326f
C610 B.n477 VSUBS 0.007326f
C611 B.n478 VSUBS 0.007326f
C612 B.n479 VSUBS 0.007326f
C613 B.n480 VSUBS 0.007326f
C614 B.n481 VSUBS 0.007326f
C615 B.n482 VSUBS 0.007326f
C616 B.n483 VSUBS 0.007326f
C617 B.n484 VSUBS 0.007326f
C618 B.n485 VSUBS 0.007326f
C619 B.n486 VSUBS 0.007326f
C620 B.n487 VSUBS 0.007326f
C621 B.n488 VSUBS 0.007326f
C622 B.n489 VSUBS 0.007326f
C623 B.n490 VSUBS 0.007326f
C624 B.n491 VSUBS 0.007326f
C625 B.n492 VSUBS 0.007326f
C626 B.n493 VSUBS 0.007326f
C627 B.n494 VSUBS 0.007326f
C628 B.n495 VSUBS 0.007326f
C629 B.n496 VSUBS 0.007326f
C630 B.n497 VSUBS 0.007326f
C631 B.n498 VSUBS 0.007326f
C632 B.n499 VSUBS 0.007326f
C633 B.n500 VSUBS 0.007326f
C634 B.n501 VSUBS 0.007326f
C635 B.n502 VSUBS 0.007326f
C636 B.n503 VSUBS 0.007326f
C637 B.n504 VSUBS 0.007326f
C638 B.n505 VSUBS 0.007326f
C639 B.n506 VSUBS 0.007326f
C640 B.n507 VSUBS 0.007326f
C641 B.n508 VSUBS 0.007326f
C642 B.n509 VSUBS 0.007326f
C643 B.n510 VSUBS 0.007326f
C644 B.n511 VSUBS 0.007326f
C645 B.n512 VSUBS 0.007326f
C646 B.n513 VSUBS 0.007326f
C647 B.n514 VSUBS 0.007326f
C648 B.n515 VSUBS 0.007326f
C649 B.n516 VSUBS 0.007326f
C650 B.n517 VSUBS 0.007326f
C651 B.n518 VSUBS 0.007326f
C652 B.n519 VSUBS 0.007326f
C653 B.n520 VSUBS 0.007326f
C654 B.n521 VSUBS 0.007326f
C655 B.n522 VSUBS 0.007326f
C656 B.n523 VSUBS 0.007326f
C657 B.n524 VSUBS 0.007326f
C658 B.n525 VSUBS 0.007326f
C659 B.n526 VSUBS 0.007326f
C660 B.n527 VSUBS 0.007326f
C661 B.n528 VSUBS 0.007326f
C662 B.n529 VSUBS 0.007326f
C663 B.n530 VSUBS 0.007326f
C664 B.n531 VSUBS 0.007326f
C665 B.n532 VSUBS 0.007326f
C666 B.n533 VSUBS 0.007326f
C667 B.n534 VSUBS 0.007326f
C668 B.n535 VSUBS 0.007326f
C669 B.n536 VSUBS 0.007326f
C670 B.n537 VSUBS 0.007326f
C671 B.n538 VSUBS 0.007326f
C672 B.n539 VSUBS 0.007326f
C673 B.n540 VSUBS 0.007326f
C674 B.n541 VSUBS 0.007326f
C675 B.n542 VSUBS 0.007326f
C676 B.n543 VSUBS 0.007326f
C677 B.n544 VSUBS 0.007326f
C678 B.n545 VSUBS 0.007326f
C679 B.n546 VSUBS 0.007326f
C680 B.n547 VSUBS 0.007326f
C681 B.n548 VSUBS 0.007326f
C682 B.n549 VSUBS 0.007326f
C683 B.n550 VSUBS 0.007326f
C684 B.n551 VSUBS 0.007326f
C685 B.n552 VSUBS 0.007326f
C686 B.n553 VSUBS 0.007326f
C687 B.n554 VSUBS 0.007326f
C688 B.n555 VSUBS 0.007326f
C689 B.n556 VSUBS 0.007326f
C690 B.n557 VSUBS 0.007326f
C691 B.n558 VSUBS 0.007326f
C692 B.n559 VSUBS 0.007326f
C693 B.n560 VSUBS 0.007326f
C694 B.n561 VSUBS 0.007326f
C695 B.n562 VSUBS 0.007326f
C696 B.n563 VSUBS 0.007326f
C697 B.n564 VSUBS 0.007326f
C698 B.n565 VSUBS 0.007326f
C699 B.n566 VSUBS 0.007326f
C700 B.n567 VSUBS 0.007326f
C701 B.n568 VSUBS 0.007326f
C702 B.n569 VSUBS 0.007326f
C703 B.n570 VSUBS 0.007326f
C704 B.n571 VSUBS 0.007326f
C705 B.n572 VSUBS 0.007326f
C706 B.n573 VSUBS 0.007326f
C707 B.n574 VSUBS 0.007326f
C708 B.n575 VSUBS 0.007326f
C709 B.n576 VSUBS 0.007326f
C710 B.n577 VSUBS 0.007326f
C711 B.n578 VSUBS 0.007326f
C712 B.n579 VSUBS 0.007326f
C713 B.n580 VSUBS 0.007326f
C714 B.n581 VSUBS 0.007326f
C715 B.n582 VSUBS 0.007326f
C716 B.n583 VSUBS 0.007326f
C717 B.n584 VSUBS 0.007326f
C718 B.n585 VSUBS 0.007326f
C719 B.n586 VSUBS 0.007326f
C720 B.n587 VSUBS 0.007326f
C721 B.n588 VSUBS 0.007326f
C722 B.n589 VSUBS 0.007326f
C723 B.n590 VSUBS 0.007326f
C724 B.n591 VSUBS 0.007326f
C725 B.n592 VSUBS 0.007326f
C726 B.n593 VSUBS 0.007326f
C727 B.n594 VSUBS 0.007326f
C728 B.n595 VSUBS 0.007326f
C729 B.n596 VSUBS 0.007326f
C730 B.n597 VSUBS 0.007326f
C731 B.n598 VSUBS 0.016795f
C732 B.n599 VSUBS 0.017894f
C733 B.n600 VSUBS 0.017894f
C734 B.n601 VSUBS 0.007326f
C735 B.n602 VSUBS 0.007326f
C736 B.n603 VSUBS 0.007326f
C737 B.n604 VSUBS 0.007326f
C738 B.n605 VSUBS 0.007326f
C739 B.n606 VSUBS 0.007326f
C740 B.n607 VSUBS 0.007326f
C741 B.n608 VSUBS 0.007326f
C742 B.n609 VSUBS 0.007326f
C743 B.n610 VSUBS 0.007326f
C744 B.n611 VSUBS 0.007326f
C745 B.n612 VSUBS 0.007326f
C746 B.n613 VSUBS 0.007326f
C747 B.n614 VSUBS 0.007326f
C748 B.n615 VSUBS 0.007326f
C749 B.n616 VSUBS 0.007326f
C750 B.n617 VSUBS 0.007326f
C751 B.n618 VSUBS 0.007326f
C752 B.n619 VSUBS 0.007326f
C753 B.n620 VSUBS 0.007326f
C754 B.n621 VSUBS 0.007326f
C755 B.n622 VSUBS 0.007326f
C756 B.n623 VSUBS 0.007326f
C757 B.n624 VSUBS 0.007326f
C758 B.n625 VSUBS 0.007326f
C759 B.n626 VSUBS 0.007326f
C760 B.n627 VSUBS 0.007326f
C761 B.n628 VSUBS 0.007326f
C762 B.n629 VSUBS 0.007326f
C763 B.n630 VSUBS 0.007326f
C764 B.n631 VSUBS 0.007326f
C765 B.n632 VSUBS 0.007326f
C766 B.n633 VSUBS 0.007326f
C767 B.n634 VSUBS 0.007326f
C768 B.n635 VSUBS 0.007326f
C769 B.n636 VSUBS 0.007326f
C770 B.n637 VSUBS 0.007326f
C771 B.n638 VSUBS 0.007326f
C772 B.n639 VSUBS 0.007326f
C773 B.n640 VSUBS 0.007326f
C774 B.n641 VSUBS 0.007326f
C775 B.n642 VSUBS 0.007326f
C776 B.n643 VSUBS 0.007326f
C777 B.n644 VSUBS 0.007326f
C778 B.n645 VSUBS 0.007326f
C779 B.n646 VSUBS 0.007326f
C780 B.n647 VSUBS 0.007326f
C781 B.n648 VSUBS 0.007326f
C782 B.n649 VSUBS 0.007326f
C783 B.n650 VSUBS 0.007326f
C784 B.n651 VSUBS 0.007326f
C785 B.n652 VSUBS 0.007326f
C786 B.n653 VSUBS 0.007326f
C787 B.n654 VSUBS 0.007326f
C788 B.n655 VSUBS 0.007326f
C789 B.n656 VSUBS 0.007326f
C790 B.n657 VSUBS 0.007326f
C791 B.n658 VSUBS 0.007326f
C792 B.n659 VSUBS 0.007326f
C793 B.n660 VSUBS 0.007326f
C794 B.n661 VSUBS 0.007326f
C795 B.n662 VSUBS 0.007326f
C796 B.n663 VSUBS 0.007326f
C797 B.n664 VSUBS 0.007326f
C798 B.n665 VSUBS 0.007326f
C799 B.n666 VSUBS 0.007326f
C800 B.n667 VSUBS 0.005063f
C801 B.n668 VSUBS 0.016973f
C802 B.n669 VSUBS 0.005925f
C803 B.n670 VSUBS 0.007326f
C804 B.n671 VSUBS 0.007326f
C805 B.n672 VSUBS 0.007326f
C806 B.n673 VSUBS 0.007326f
C807 B.n674 VSUBS 0.007326f
C808 B.n675 VSUBS 0.007326f
C809 B.n676 VSUBS 0.007326f
C810 B.n677 VSUBS 0.007326f
C811 B.n678 VSUBS 0.007326f
C812 B.n679 VSUBS 0.007326f
C813 B.n680 VSUBS 0.007326f
C814 B.n681 VSUBS 0.005925f
C815 B.n682 VSUBS 0.007326f
C816 B.n683 VSUBS 0.007326f
C817 B.n684 VSUBS 0.007326f
C818 B.n685 VSUBS 0.007326f
C819 B.n686 VSUBS 0.007326f
C820 B.n687 VSUBS 0.007326f
C821 B.n688 VSUBS 0.007326f
C822 B.n689 VSUBS 0.007326f
C823 B.n690 VSUBS 0.007326f
C824 B.n691 VSUBS 0.007326f
C825 B.n692 VSUBS 0.007326f
C826 B.n693 VSUBS 0.007326f
C827 B.n694 VSUBS 0.007326f
C828 B.n695 VSUBS 0.007326f
C829 B.n696 VSUBS 0.007326f
C830 B.n697 VSUBS 0.007326f
C831 B.n698 VSUBS 0.007326f
C832 B.n699 VSUBS 0.007326f
C833 B.n700 VSUBS 0.007326f
C834 B.n701 VSUBS 0.007326f
C835 B.n702 VSUBS 0.007326f
C836 B.n703 VSUBS 0.007326f
C837 B.n704 VSUBS 0.007326f
C838 B.n705 VSUBS 0.007326f
C839 B.n706 VSUBS 0.007326f
C840 B.n707 VSUBS 0.007326f
C841 B.n708 VSUBS 0.007326f
C842 B.n709 VSUBS 0.007326f
C843 B.n710 VSUBS 0.007326f
C844 B.n711 VSUBS 0.007326f
C845 B.n712 VSUBS 0.007326f
C846 B.n713 VSUBS 0.007326f
C847 B.n714 VSUBS 0.007326f
C848 B.n715 VSUBS 0.007326f
C849 B.n716 VSUBS 0.007326f
C850 B.n717 VSUBS 0.007326f
C851 B.n718 VSUBS 0.007326f
C852 B.n719 VSUBS 0.007326f
C853 B.n720 VSUBS 0.007326f
C854 B.n721 VSUBS 0.007326f
C855 B.n722 VSUBS 0.007326f
C856 B.n723 VSUBS 0.007326f
C857 B.n724 VSUBS 0.007326f
C858 B.n725 VSUBS 0.007326f
C859 B.n726 VSUBS 0.007326f
C860 B.n727 VSUBS 0.007326f
C861 B.n728 VSUBS 0.007326f
C862 B.n729 VSUBS 0.007326f
C863 B.n730 VSUBS 0.007326f
C864 B.n731 VSUBS 0.007326f
C865 B.n732 VSUBS 0.007326f
C866 B.n733 VSUBS 0.007326f
C867 B.n734 VSUBS 0.007326f
C868 B.n735 VSUBS 0.007326f
C869 B.n736 VSUBS 0.007326f
C870 B.n737 VSUBS 0.007326f
C871 B.n738 VSUBS 0.007326f
C872 B.n739 VSUBS 0.007326f
C873 B.n740 VSUBS 0.007326f
C874 B.n741 VSUBS 0.007326f
C875 B.n742 VSUBS 0.007326f
C876 B.n743 VSUBS 0.007326f
C877 B.n744 VSUBS 0.007326f
C878 B.n745 VSUBS 0.007326f
C879 B.n746 VSUBS 0.007326f
C880 B.n747 VSUBS 0.007326f
C881 B.n748 VSUBS 0.007326f
C882 B.n749 VSUBS 0.007326f
C883 B.n750 VSUBS 0.017894f
C884 B.n751 VSUBS 0.017894f
C885 B.n752 VSUBS 0.016795f
C886 B.n753 VSUBS 0.007326f
C887 B.n754 VSUBS 0.007326f
C888 B.n755 VSUBS 0.007326f
C889 B.n756 VSUBS 0.007326f
C890 B.n757 VSUBS 0.007326f
C891 B.n758 VSUBS 0.007326f
C892 B.n759 VSUBS 0.007326f
C893 B.n760 VSUBS 0.007326f
C894 B.n761 VSUBS 0.007326f
C895 B.n762 VSUBS 0.007326f
C896 B.n763 VSUBS 0.007326f
C897 B.n764 VSUBS 0.007326f
C898 B.n765 VSUBS 0.007326f
C899 B.n766 VSUBS 0.007326f
C900 B.n767 VSUBS 0.007326f
C901 B.n768 VSUBS 0.007326f
C902 B.n769 VSUBS 0.007326f
C903 B.n770 VSUBS 0.007326f
C904 B.n771 VSUBS 0.007326f
C905 B.n772 VSUBS 0.007326f
C906 B.n773 VSUBS 0.007326f
C907 B.n774 VSUBS 0.007326f
C908 B.n775 VSUBS 0.007326f
C909 B.n776 VSUBS 0.007326f
C910 B.n777 VSUBS 0.007326f
C911 B.n778 VSUBS 0.007326f
C912 B.n779 VSUBS 0.007326f
C913 B.n780 VSUBS 0.007326f
C914 B.n781 VSUBS 0.007326f
C915 B.n782 VSUBS 0.007326f
C916 B.n783 VSUBS 0.007326f
C917 B.n784 VSUBS 0.007326f
C918 B.n785 VSUBS 0.007326f
C919 B.n786 VSUBS 0.007326f
C920 B.n787 VSUBS 0.007326f
C921 B.n788 VSUBS 0.007326f
C922 B.n789 VSUBS 0.007326f
C923 B.n790 VSUBS 0.007326f
C924 B.n791 VSUBS 0.007326f
C925 B.n792 VSUBS 0.007326f
C926 B.n793 VSUBS 0.007326f
C927 B.n794 VSUBS 0.007326f
C928 B.n795 VSUBS 0.007326f
C929 B.n796 VSUBS 0.007326f
C930 B.n797 VSUBS 0.007326f
C931 B.n798 VSUBS 0.007326f
C932 B.n799 VSUBS 0.007326f
C933 B.n800 VSUBS 0.007326f
C934 B.n801 VSUBS 0.007326f
C935 B.n802 VSUBS 0.007326f
C936 B.n803 VSUBS 0.007326f
C937 B.n804 VSUBS 0.007326f
C938 B.n805 VSUBS 0.007326f
C939 B.n806 VSUBS 0.007326f
C940 B.n807 VSUBS 0.007326f
C941 B.n808 VSUBS 0.007326f
C942 B.n809 VSUBS 0.007326f
C943 B.n810 VSUBS 0.007326f
C944 B.n811 VSUBS 0.007326f
C945 B.n812 VSUBS 0.007326f
C946 B.n813 VSUBS 0.007326f
C947 B.n814 VSUBS 0.007326f
C948 B.n815 VSUBS 0.007326f
C949 B.n816 VSUBS 0.007326f
C950 B.n817 VSUBS 0.007326f
C951 B.n818 VSUBS 0.007326f
C952 B.n819 VSUBS 0.007326f
C953 B.n820 VSUBS 0.007326f
C954 B.n821 VSUBS 0.007326f
C955 B.n822 VSUBS 0.007326f
C956 B.n823 VSUBS 0.007326f
C957 B.n824 VSUBS 0.007326f
C958 B.n825 VSUBS 0.007326f
C959 B.n826 VSUBS 0.007326f
C960 B.n827 VSUBS 0.00956f
C961 B.n828 VSUBS 0.010184f
C962 B.n829 VSUBS 0.020251f
C963 VDD2.t1 VSUBS 0.28679f
C964 VDD2.t7 VSUBS 0.28679f
C965 VDD2.n0 VSUBS 2.31446f
C966 VDD2.t2 VSUBS 0.28679f
C967 VDD2.t3 VSUBS 0.28679f
C968 VDD2.n1 VSUBS 2.31446f
C969 VDD2.n2 VSUBS 4.21287f
C970 VDD2.t0 VSUBS 0.28679f
C971 VDD2.t6 VSUBS 0.28679f
C972 VDD2.n3 VSUBS 2.30109f
C973 VDD2.n4 VSUBS 3.60108f
C974 VDD2.t5 VSUBS 0.28679f
C975 VDD2.t4 VSUBS 0.28679f
C976 VDD2.n5 VSUBS 2.31441f
C977 VTAIL.t15 VSUBS 0.260118f
C978 VTAIL.t10 VSUBS 0.260118f
C979 VTAIL.n0 VSUBS 1.96011f
C980 VTAIL.n1 VSUBS 0.751177f
C981 VTAIL.n2 VSUBS 0.026754f
C982 VTAIL.n3 VSUBS 0.02462f
C983 VTAIL.n4 VSUBS 0.01323f
C984 VTAIL.n5 VSUBS 0.03127f
C985 VTAIL.n6 VSUBS 0.014008f
C986 VTAIL.n7 VSUBS 0.02462f
C987 VTAIL.n8 VSUBS 0.01323f
C988 VTAIL.n9 VSUBS 0.03127f
C989 VTAIL.n10 VSUBS 0.014008f
C990 VTAIL.n11 VSUBS 0.02462f
C991 VTAIL.n12 VSUBS 0.01323f
C992 VTAIL.n13 VSUBS 0.03127f
C993 VTAIL.n14 VSUBS 0.014008f
C994 VTAIL.n15 VSUBS 0.02462f
C995 VTAIL.n16 VSUBS 0.01323f
C996 VTAIL.n17 VSUBS 0.03127f
C997 VTAIL.n18 VSUBS 0.014008f
C998 VTAIL.n19 VSUBS 0.02462f
C999 VTAIL.n20 VSUBS 0.01323f
C1000 VTAIL.n21 VSUBS 0.03127f
C1001 VTAIL.n22 VSUBS 0.014008f
C1002 VTAIL.n23 VSUBS 1.38984f
C1003 VTAIL.n24 VSUBS 0.01323f
C1004 VTAIL.t11 VSUBS 0.066844f
C1005 VTAIL.n25 VSUBS 0.161713f
C1006 VTAIL.n26 VSUBS 0.019893f
C1007 VTAIL.n27 VSUBS 0.023452f
C1008 VTAIL.n28 VSUBS 0.03127f
C1009 VTAIL.n29 VSUBS 0.014008f
C1010 VTAIL.n30 VSUBS 0.01323f
C1011 VTAIL.n31 VSUBS 0.02462f
C1012 VTAIL.n32 VSUBS 0.02462f
C1013 VTAIL.n33 VSUBS 0.01323f
C1014 VTAIL.n34 VSUBS 0.014008f
C1015 VTAIL.n35 VSUBS 0.03127f
C1016 VTAIL.n36 VSUBS 0.03127f
C1017 VTAIL.n37 VSUBS 0.014008f
C1018 VTAIL.n38 VSUBS 0.01323f
C1019 VTAIL.n39 VSUBS 0.02462f
C1020 VTAIL.n40 VSUBS 0.02462f
C1021 VTAIL.n41 VSUBS 0.01323f
C1022 VTAIL.n42 VSUBS 0.014008f
C1023 VTAIL.n43 VSUBS 0.03127f
C1024 VTAIL.n44 VSUBS 0.03127f
C1025 VTAIL.n45 VSUBS 0.014008f
C1026 VTAIL.n46 VSUBS 0.01323f
C1027 VTAIL.n47 VSUBS 0.02462f
C1028 VTAIL.n48 VSUBS 0.02462f
C1029 VTAIL.n49 VSUBS 0.01323f
C1030 VTAIL.n50 VSUBS 0.014008f
C1031 VTAIL.n51 VSUBS 0.03127f
C1032 VTAIL.n52 VSUBS 0.03127f
C1033 VTAIL.n53 VSUBS 0.014008f
C1034 VTAIL.n54 VSUBS 0.01323f
C1035 VTAIL.n55 VSUBS 0.02462f
C1036 VTAIL.n56 VSUBS 0.02462f
C1037 VTAIL.n57 VSUBS 0.01323f
C1038 VTAIL.n58 VSUBS 0.014008f
C1039 VTAIL.n59 VSUBS 0.03127f
C1040 VTAIL.n60 VSUBS 0.03127f
C1041 VTAIL.n61 VSUBS 0.014008f
C1042 VTAIL.n62 VSUBS 0.01323f
C1043 VTAIL.n63 VSUBS 0.02462f
C1044 VTAIL.n64 VSUBS 0.02462f
C1045 VTAIL.n65 VSUBS 0.01323f
C1046 VTAIL.n66 VSUBS 0.014008f
C1047 VTAIL.n67 VSUBS 0.03127f
C1048 VTAIL.n68 VSUBS 0.078096f
C1049 VTAIL.n69 VSUBS 0.014008f
C1050 VTAIL.n70 VSUBS 0.02598f
C1051 VTAIL.n71 VSUBS 0.062625f
C1052 VTAIL.n72 VSUBS 0.060047f
C1053 VTAIL.n73 VSUBS 0.263963f
C1054 VTAIL.n74 VSUBS 0.026754f
C1055 VTAIL.n75 VSUBS 0.02462f
C1056 VTAIL.n76 VSUBS 0.01323f
C1057 VTAIL.n77 VSUBS 0.03127f
C1058 VTAIL.n78 VSUBS 0.014008f
C1059 VTAIL.n79 VSUBS 0.02462f
C1060 VTAIL.n80 VSUBS 0.01323f
C1061 VTAIL.n81 VSUBS 0.03127f
C1062 VTAIL.n82 VSUBS 0.014008f
C1063 VTAIL.n83 VSUBS 0.02462f
C1064 VTAIL.n84 VSUBS 0.01323f
C1065 VTAIL.n85 VSUBS 0.03127f
C1066 VTAIL.n86 VSUBS 0.014008f
C1067 VTAIL.n87 VSUBS 0.02462f
C1068 VTAIL.n88 VSUBS 0.01323f
C1069 VTAIL.n89 VSUBS 0.03127f
C1070 VTAIL.n90 VSUBS 0.014008f
C1071 VTAIL.n91 VSUBS 0.02462f
C1072 VTAIL.n92 VSUBS 0.01323f
C1073 VTAIL.n93 VSUBS 0.03127f
C1074 VTAIL.n94 VSUBS 0.014008f
C1075 VTAIL.n95 VSUBS 1.38984f
C1076 VTAIL.n96 VSUBS 0.01323f
C1077 VTAIL.t4 VSUBS 0.066844f
C1078 VTAIL.n97 VSUBS 0.161713f
C1079 VTAIL.n98 VSUBS 0.019893f
C1080 VTAIL.n99 VSUBS 0.023452f
C1081 VTAIL.n100 VSUBS 0.03127f
C1082 VTAIL.n101 VSUBS 0.014008f
C1083 VTAIL.n102 VSUBS 0.01323f
C1084 VTAIL.n103 VSUBS 0.02462f
C1085 VTAIL.n104 VSUBS 0.02462f
C1086 VTAIL.n105 VSUBS 0.01323f
C1087 VTAIL.n106 VSUBS 0.014008f
C1088 VTAIL.n107 VSUBS 0.03127f
C1089 VTAIL.n108 VSUBS 0.03127f
C1090 VTAIL.n109 VSUBS 0.014008f
C1091 VTAIL.n110 VSUBS 0.01323f
C1092 VTAIL.n111 VSUBS 0.02462f
C1093 VTAIL.n112 VSUBS 0.02462f
C1094 VTAIL.n113 VSUBS 0.01323f
C1095 VTAIL.n114 VSUBS 0.014008f
C1096 VTAIL.n115 VSUBS 0.03127f
C1097 VTAIL.n116 VSUBS 0.03127f
C1098 VTAIL.n117 VSUBS 0.014008f
C1099 VTAIL.n118 VSUBS 0.01323f
C1100 VTAIL.n119 VSUBS 0.02462f
C1101 VTAIL.n120 VSUBS 0.02462f
C1102 VTAIL.n121 VSUBS 0.01323f
C1103 VTAIL.n122 VSUBS 0.014008f
C1104 VTAIL.n123 VSUBS 0.03127f
C1105 VTAIL.n124 VSUBS 0.03127f
C1106 VTAIL.n125 VSUBS 0.014008f
C1107 VTAIL.n126 VSUBS 0.01323f
C1108 VTAIL.n127 VSUBS 0.02462f
C1109 VTAIL.n128 VSUBS 0.02462f
C1110 VTAIL.n129 VSUBS 0.01323f
C1111 VTAIL.n130 VSUBS 0.014008f
C1112 VTAIL.n131 VSUBS 0.03127f
C1113 VTAIL.n132 VSUBS 0.03127f
C1114 VTAIL.n133 VSUBS 0.014008f
C1115 VTAIL.n134 VSUBS 0.01323f
C1116 VTAIL.n135 VSUBS 0.02462f
C1117 VTAIL.n136 VSUBS 0.02462f
C1118 VTAIL.n137 VSUBS 0.01323f
C1119 VTAIL.n138 VSUBS 0.014008f
C1120 VTAIL.n139 VSUBS 0.03127f
C1121 VTAIL.n140 VSUBS 0.078096f
C1122 VTAIL.n141 VSUBS 0.014008f
C1123 VTAIL.n142 VSUBS 0.02598f
C1124 VTAIL.n143 VSUBS 0.062625f
C1125 VTAIL.n144 VSUBS 0.060047f
C1126 VTAIL.n145 VSUBS 0.263963f
C1127 VTAIL.t2 VSUBS 0.260118f
C1128 VTAIL.t7 VSUBS 0.260118f
C1129 VTAIL.n146 VSUBS 1.96011f
C1130 VTAIL.n147 VSUBS 0.948991f
C1131 VTAIL.n148 VSUBS 0.026754f
C1132 VTAIL.n149 VSUBS 0.02462f
C1133 VTAIL.n150 VSUBS 0.01323f
C1134 VTAIL.n151 VSUBS 0.03127f
C1135 VTAIL.n152 VSUBS 0.014008f
C1136 VTAIL.n153 VSUBS 0.02462f
C1137 VTAIL.n154 VSUBS 0.01323f
C1138 VTAIL.n155 VSUBS 0.03127f
C1139 VTAIL.n156 VSUBS 0.014008f
C1140 VTAIL.n157 VSUBS 0.02462f
C1141 VTAIL.n158 VSUBS 0.01323f
C1142 VTAIL.n159 VSUBS 0.03127f
C1143 VTAIL.n160 VSUBS 0.014008f
C1144 VTAIL.n161 VSUBS 0.02462f
C1145 VTAIL.n162 VSUBS 0.01323f
C1146 VTAIL.n163 VSUBS 0.03127f
C1147 VTAIL.n164 VSUBS 0.014008f
C1148 VTAIL.n165 VSUBS 0.02462f
C1149 VTAIL.n166 VSUBS 0.01323f
C1150 VTAIL.n167 VSUBS 0.03127f
C1151 VTAIL.n168 VSUBS 0.014008f
C1152 VTAIL.n169 VSUBS 1.38984f
C1153 VTAIL.n170 VSUBS 0.01323f
C1154 VTAIL.t5 VSUBS 0.066844f
C1155 VTAIL.n171 VSUBS 0.161713f
C1156 VTAIL.n172 VSUBS 0.019893f
C1157 VTAIL.n173 VSUBS 0.023452f
C1158 VTAIL.n174 VSUBS 0.03127f
C1159 VTAIL.n175 VSUBS 0.014008f
C1160 VTAIL.n176 VSUBS 0.01323f
C1161 VTAIL.n177 VSUBS 0.02462f
C1162 VTAIL.n178 VSUBS 0.02462f
C1163 VTAIL.n179 VSUBS 0.01323f
C1164 VTAIL.n180 VSUBS 0.014008f
C1165 VTAIL.n181 VSUBS 0.03127f
C1166 VTAIL.n182 VSUBS 0.03127f
C1167 VTAIL.n183 VSUBS 0.014008f
C1168 VTAIL.n184 VSUBS 0.01323f
C1169 VTAIL.n185 VSUBS 0.02462f
C1170 VTAIL.n186 VSUBS 0.02462f
C1171 VTAIL.n187 VSUBS 0.01323f
C1172 VTAIL.n188 VSUBS 0.014008f
C1173 VTAIL.n189 VSUBS 0.03127f
C1174 VTAIL.n190 VSUBS 0.03127f
C1175 VTAIL.n191 VSUBS 0.014008f
C1176 VTAIL.n192 VSUBS 0.01323f
C1177 VTAIL.n193 VSUBS 0.02462f
C1178 VTAIL.n194 VSUBS 0.02462f
C1179 VTAIL.n195 VSUBS 0.01323f
C1180 VTAIL.n196 VSUBS 0.014008f
C1181 VTAIL.n197 VSUBS 0.03127f
C1182 VTAIL.n198 VSUBS 0.03127f
C1183 VTAIL.n199 VSUBS 0.014008f
C1184 VTAIL.n200 VSUBS 0.01323f
C1185 VTAIL.n201 VSUBS 0.02462f
C1186 VTAIL.n202 VSUBS 0.02462f
C1187 VTAIL.n203 VSUBS 0.01323f
C1188 VTAIL.n204 VSUBS 0.014008f
C1189 VTAIL.n205 VSUBS 0.03127f
C1190 VTAIL.n206 VSUBS 0.03127f
C1191 VTAIL.n207 VSUBS 0.014008f
C1192 VTAIL.n208 VSUBS 0.01323f
C1193 VTAIL.n209 VSUBS 0.02462f
C1194 VTAIL.n210 VSUBS 0.02462f
C1195 VTAIL.n211 VSUBS 0.01323f
C1196 VTAIL.n212 VSUBS 0.014008f
C1197 VTAIL.n213 VSUBS 0.03127f
C1198 VTAIL.n214 VSUBS 0.078096f
C1199 VTAIL.n215 VSUBS 0.014008f
C1200 VTAIL.n216 VSUBS 0.02598f
C1201 VTAIL.n217 VSUBS 0.062625f
C1202 VTAIL.n218 VSUBS 0.060047f
C1203 VTAIL.n219 VSUBS 1.67791f
C1204 VTAIL.n220 VSUBS 0.026754f
C1205 VTAIL.n221 VSUBS 0.02462f
C1206 VTAIL.n222 VSUBS 0.01323f
C1207 VTAIL.n223 VSUBS 0.03127f
C1208 VTAIL.n224 VSUBS 0.014008f
C1209 VTAIL.n225 VSUBS 0.02462f
C1210 VTAIL.n226 VSUBS 0.01323f
C1211 VTAIL.n227 VSUBS 0.03127f
C1212 VTAIL.n228 VSUBS 0.014008f
C1213 VTAIL.n229 VSUBS 0.02462f
C1214 VTAIL.n230 VSUBS 0.01323f
C1215 VTAIL.n231 VSUBS 0.03127f
C1216 VTAIL.n232 VSUBS 0.014008f
C1217 VTAIL.n233 VSUBS 0.02462f
C1218 VTAIL.n234 VSUBS 0.01323f
C1219 VTAIL.n235 VSUBS 0.03127f
C1220 VTAIL.n236 VSUBS 0.014008f
C1221 VTAIL.n237 VSUBS 0.02462f
C1222 VTAIL.n238 VSUBS 0.01323f
C1223 VTAIL.n239 VSUBS 0.03127f
C1224 VTAIL.n240 VSUBS 0.014008f
C1225 VTAIL.n241 VSUBS 1.38984f
C1226 VTAIL.n242 VSUBS 0.01323f
C1227 VTAIL.t12 VSUBS 0.066844f
C1228 VTAIL.n243 VSUBS 0.161713f
C1229 VTAIL.n244 VSUBS 0.019893f
C1230 VTAIL.n245 VSUBS 0.023452f
C1231 VTAIL.n246 VSUBS 0.03127f
C1232 VTAIL.n247 VSUBS 0.014008f
C1233 VTAIL.n248 VSUBS 0.01323f
C1234 VTAIL.n249 VSUBS 0.02462f
C1235 VTAIL.n250 VSUBS 0.02462f
C1236 VTAIL.n251 VSUBS 0.01323f
C1237 VTAIL.n252 VSUBS 0.014008f
C1238 VTAIL.n253 VSUBS 0.03127f
C1239 VTAIL.n254 VSUBS 0.03127f
C1240 VTAIL.n255 VSUBS 0.014008f
C1241 VTAIL.n256 VSUBS 0.01323f
C1242 VTAIL.n257 VSUBS 0.02462f
C1243 VTAIL.n258 VSUBS 0.02462f
C1244 VTAIL.n259 VSUBS 0.01323f
C1245 VTAIL.n260 VSUBS 0.014008f
C1246 VTAIL.n261 VSUBS 0.03127f
C1247 VTAIL.n262 VSUBS 0.03127f
C1248 VTAIL.n263 VSUBS 0.014008f
C1249 VTAIL.n264 VSUBS 0.01323f
C1250 VTAIL.n265 VSUBS 0.02462f
C1251 VTAIL.n266 VSUBS 0.02462f
C1252 VTAIL.n267 VSUBS 0.01323f
C1253 VTAIL.n268 VSUBS 0.014008f
C1254 VTAIL.n269 VSUBS 0.03127f
C1255 VTAIL.n270 VSUBS 0.03127f
C1256 VTAIL.n271 VSUBS 0.014008f
C1257 VTAIL.n272 VSUBS 0.01323f
C1258 VTAIL.n273 VSUBS 0.02462f
C1259 VTAIL.n274 VSUBS 0.02462f
C1260 VTAIL.n275 VSUBS 0.01323f
C1261 VTAIL.n276 VSUBS 0.014008f
C1262 VTAIL.n277 VSUBS 0.03127f
C1263 VTAIL.n278 VSUBS 0.03127f
C1264 VTAIL.n279 VSUBS 0.014008f
C1265 VTAIL.n280 VSUBS 0.01323f
C1266 VTAIL.n281 VSUBS 0.02462f
C1267 VTAIL.n282 VSUBS 0.02462f
C1268 VTAIL.n283 VSUBS 0.01323f
C1269 VTAIL.n284 VSUBS 0.014008f
C1270 VTAIL.n285 VSUBS 0.03127f
C1271 VTAIL.n286 VSUBS 0.078096f
C1272 VTAIL.n287 VSUBS 0.014008f
C1273 VTAIL.n288 VSUBS 0.02598f
C1274 VTAIL.n289 VSUBS 0.062625f
C1275 VTAIL.n290 VSUBS 0.060047f
C1276 VTAIL.n291 VSUBS 1.67791f
C1277 VTAIL.t14 VSUBS 0.260118f
C1278 VTAIL.t13 VSUBS 0.260118f
C1279 VTAIL.n292 VSUBS 1.96013f
C1280 VTAIL.n293 VSUBS 0.948978f
C1281 VTAIL.n294 VSUBS 0.026754f
C1282 VTAIL.n295 VSUBS 0.02462f
C1283 VTAIL.n296 VSUBS 0.01323f
C1284 VTAIL.n297 VSUBS 0.03127f
C1285 VTAIL.n298 VSUBS 0.014008f
C1286 VTAIL.n299 VSUBS 0.02462f
C1287 VTAIL.n300 VSUBS 0.01323f
C1288 VTAIL.n301 VSUBS 0.03127f
C1289 VTAIL.n302 VSUBS 0.014008f
C1290 VTAIL.n303 VSUBS 0.02462f
C1291 VTAIL.n304 VSUBS 0.01323f
C1292 VTAIL.n305 VSUBS 0.03127f
C1293 VTAIL.n306 VSUBS 0.014008f
C1294 VTAIL.n307 VSUBS 0.02462f
C1295 VTAIL.n308 VSUBS 0.01323f
C1296 VTAIL.n309 VSUBS 0.03127f
C1297 VTAIL.n310 VSUBS 0.014008f
C1298 VTAIL.n311 VSUBS 0.02462f
C1299 VTAIL.n312 VSUBS 0.01323f
C1300 VTAIL.n313 VSUBS 0.03127f
C1301 VTAIL.n314 VSUBS 0.014008f
C1302 VTAIL.n315 VSUBS 1.38984f
C1303 VTAIL.n316 VSUBS 0.01323f
C1304 VTAIL.t8 VSUBS 0.066844f
C1305 VTAIL.n317 VSUBS 0.161713f
C1306 VTAIL.n318 VSUBS 0.019893f
C1307 VTAIL.n319 VSUBS 0.023452f
C1308 VTAIL.n320 VSUBS 0.03127f
C1309 VTAIL.n321 VSUBS 0.014008f
C1310 VTAIL.n322 VSUBS 0.01323f
C1311 VTAIL.n323 VSUBS 0.02462f
C1312 VTAIL.n324 VSUBS 0.02462f
C1313 VTAIL.n325 VSUBS 0.01323f
C1314 VTAIL.n326 VSUBS 0.014008f
C1315 VTAIL.n327 VSUBS 0.03127f
C1316 VTAIL.n328 VSUBS 0.03127f
C1317 VTAIL.n329 VSUBS 0.014008f
C1318 VTAIL.n330 VSUBS 0.01323f
C1319 VTAIL.n331 VSUBS 0.02462f
C1320 VTAIL.n332 VSUBS 0.02462f
C1321 VTAIL.n333 VSUBS 0.01323f
C1322 VTAIL.n334 VSUBS 0.014008f
C1323 VTAIL.n335 VSUBS 0.03127f
C1324 VTAIL.n336 VSUBS 0.03127f
C1325 VTAIL.n337 VSUBS 0.014008f
C1326 VTAIL.n338 VSUBS 0.01323f
C1327 VTAIL.n339 VSUBS 0.02462f
C1328 VTAIL.n340 VSUBS 0.02462f
C1329 VTAIL.n341 VSUBS 0.01323f
C1330 VTAIL.n342 VSUBS 0.014008f
C1331 VTAIL.n343 VSUBS 0.03127f
C1332 VTAIL.n344 VSUBS 0.03127f
C1333 VTAIL.n345 VSUBS 0.014008f
C1334 VTAIL.n346 VSUBS 0.01323f
C1335 VTAIL.n347 VSUBS 0.02462f
C1336 VTAIL.n348 VSUBS 0.02462f
C1337 VTAIL.n349 VSUBS 0.01323f
C1338 VTAIL.n350 VSUBS 0.014008f
C1339 VTAIL.n351 VSUBS 0.03127f
C1340 VTAIL.n352 VSUBS 0.03127f
C1341 VTAIL.n353 VSUBS 0.014008f
C1342 VTAIL.n354 VSUBS 0.01323f
C1343 VTAIL.n355 VSUBS 0.02462f
C1344 VTAIL.n356 VSUBS 0.02462f
C1345 VTAIL.n357 VSUBS 0.01323f
C1346 VTAIL.n358 VSUBS 0.014008f
C1347 VTAIL.n359 VSUBS 0.03127f
C1348 VTAIL.n360 VSUBS 0.078096f
C1349 VTAIL.n361 VSUBS 0.014008f
C1350 VTAIL.n362 VSUBS 0.02598f
C1351 VTAIL.n363 VSUBS 0.062625f
C1352 VTAIL.n364 VSUBS 0.060047f
C1353 VTAIL.n365 VSUBS 0.263963f
C1354 VTAIL.n366 VSUBS 0.026754f
C1355 VTAIL.n367 VSUBS 0.02462f
C1356 VTAIL.n368 VSUBS 0.01323f
C1357 VTAIL.n369 VSUBS 0.03127f
C1358 VTAIL.n370 VSUBS 0.014008f
C1359 VTAIL.n371 VSUBS 0.02462f
C1360 VTAIL.n372 VSUBS 0.01323f
C1361 VTAIL.n373 VSUBS 0.03127f
C1362 VTAIL.n374 VSUBS 0.014008f
C1363 VTAIL.n375 VSUBS 0.02462f
C1364 VTAIL.n376 VSUBS 0.01323f
C1365 VTAIL.n377 VSUBS 0.03127f
C1366 VTAIL.n378 VSUBS 0.014008f
C1367 VTAIL.n379 VSUBS 0.02462f
C1368 VTAIL.n380 VSUBS 0.01323f
C1369 VTAIL.n381 VSUBS 0.03127f
C1370 VTAIL.n382 VSUBS 0.014008f
C1371 VTAIL.n383 VSUBS 0.02462f
C1372 VTAIL.n384 VSUBS 0.01323f
C1373 VTAIL.n385 VSUBS 0.03127f
C1374 VTAIL.n386 VSUBS 0.014008f
C1375 VTAIL.n387 VSUBS 1.38984f
C1376 VTAIL.n388 VSUBS 0.01323f
C1377 VTAIL.t3 VSUBS 0.066844f
C1378 VTAIL.n389 VSUBS 0.161713f
C1379 VTAIL.n390 VSUBS 0.019893f
C1380 VTAIL.n391 VSUBS 0.023452f
C1381 VTAIL.n392 VSUBS 0.03127f
C1382 VTAIL.n393 VSUBS 0.014008f
C1383 VTAIL.n394 VSUBS 0.01323f
C1384 VTAIL.n395 VSUBS 0.02462f
C1385 VTAIL.n396 VSUBS 0.02462f
C1386 VTAIL.n397 VSUBS 0.01323f
C1387 VTAIL.n398 VSUBS 0.014008f
C1388 VTAIL.n399 VSUBS 0.03127f
C1389 VTAIL.n400 VSUBS 0.03127f
C1390 VTAIL.n401 VSUBS 0.014008f
C1391 VTAIL.n402 VSUBS 0.01323f
C1392 VTAIL.n403 VSUBS 0.02462f
C1393 VTAIL.n404 VSUBS 0.02462f
C1394 VTAIL.n405 VSUBS 0.01323f
C1395 VTAIL.n406 VSUBS 0.014008f
C1396 VTAIL.n407 VSUBS 0.03127f
C1397 VTAIL.n408 VSUBS 0.03127f
C1398 VTAIL.n409 VSUBS 0.014008f
C1399 VTAIL.n410 VSUBS 0.01323f
C1400 VTAIL.n411 VSUBS 0.02462f
C1401 VTAIL.n412 VSUBS 0.02462f
C1402 VTAIL.n413 VSUBS 0.01323f
C1403 VTAIL.n414 VSUBS 0.014008f
C1404 VTAIL.n415 VSUBS 0.03127f
C1405 VTAIL.n416 VSUBS 0.03127f
C1406 VTAIL.n417 VSUBS 0.014008f
C1407 VTAIL.n418 VSUBS 0.01323f
C1408 VTAIL.n419 VSUBS 0.02462f
C1409 VTAIL.n420 VSUBS 0.02462f
C1410 VTAIL.n421 VSUBS 0.01323f
C1411 VTAIL.n422 VSUBS 0.014008f
C1412 VTAIL.n423 VSUBS 0.03127f
C1413 VTAIL.n424 VSUBS 0.03127f
C1414 VTAIL.n425 VSUBS 0.014008f
C1415 VTAIL.n426 VSUBS 0.01323f
C1416 VTAIL.n427 VSUBS 0.02462f
C1417 VTAIL.n428 VSUBS 0.02462f
C1418 VTAIL.n429 VSUBS 0.01323f
C1419 VTAIL.n430 VSUBS 0.014008f
C1420 VTAIL.n431 VSUBS 0.03127f
C1421 VTAIL.n432 VSUBS 0.078096f
C1422 VTAIL.n433 VSUBS 0.014008f
C1423 VTAIL.n434 VSUBS 0.02598f
C1424 VTAIL.n435 VSUBS 0.062625f
C1425 VTAIL.n436 VSUBS 0.060047f
C1426 VTAIL.n437 VSUBS 0.263963f
C1427 VTAIL.t1 VSUBS 0.260118f
C1428 VTAIL.t0 VSUBS 0.260118f
C1429 VTAIL.n438 VSUBS 1.96013f
C1430 VTAIL.n439 VSUBS 0.948978f
C1431 VTAIL.n440 VSUBS 0.026754f
C1432 VTAIL.n441 VSUBS 0.02462f
C1433 VTAIL.n442 VSUBS 0.01323f
C1434 VTAIL.n443 VSUBS 0.03127f
C1435 VTAIL.n444 VSUBS 0.014008f
C1436 VTAIL.n445 VSUBS 0.02462f
C1437 VTAIL.n446 VSUBS 0.01323f
C1438 VTAIL.n447 VSUBS 0.03127f
C1439 VTAIL.n448 VSUBS 0.014008f
C1440 VTAIL.n449 VSUBS 0.02462f
C1441 VTAIL.n450 VSUBS 0.01323f
C1442 VTAIL.n451 VSUBS 0.03127f
C1443 VTAIL.n452 VSUBS 0.014008f
C1444 VTAIL.n453 VSUBS 0.02462f
C1445 VTAIL.n454 VSUBS 0.01323f
C1446 VTAIL.n455 VSUBS 0.03127f
C1447 VTAIL.n456 VSUBS 0.014008f
C1448 VTAIL.n457 VSUBS 0.02462f
C1449 VTAIL.n458 VSUBS 0.01323f
C1450 VTAIL.n459 VSUBS 0.03127f
C1451 VTAIL.n460 VSUBS 0.014008f
C1452 VTAIL.n461 VSUBS 1.38984f
C1453 VTAIL.n462 VSUBS 0.01323f
C1454 VTAIL.t6 VSUBS 0.066844f
C1455 VTAIL.n463 VSUBS 0.161713f
C1456 VTAIL.n464 VSUBS 0.019893f
C1457 VTAIL.n465 VSUBS 0.023452f
C1458 VTAIL.n466 VSUBS 0.03127f
C1459 VTAIL.n467 VSUBS 0.014008f
C1460 VTAIL.n468 VSUBS 0.01323f
C1461 VTAIL.n469 VSUBS 0.02462f
C1462 VTAIL.n470 VSUBS 0.02462f
C1463 VTAIL.n471 VSUBS 0.01323f
C1464 VTAIL.n472 VSUBS 0.014008f
C1465 VTAIL.n473 VSUBS 0.03127f
C1466 VTAIL.n474 VSUBS 0.03127f
C1467 VTAIL.n475 VSUBS 0.014008f
C1468 VTAIL.n476 VSUBS 0.01323f
C1469 VTAIL.n477 VSUBS 0.02462f
C1470 VTAIL.n478 VSUBS 0.02462f
C1471 VTAIL.n479 VSUBS 0.01323f
C1472 VTAIL.n480 VSUBS 0.014008f
C1473 VTAIL.n481 VSUBS 0.03127f
C1474 VTAIL.n482 VSUBS 0.03127f
C1475 VTAIL.n483 VSUBS 0.014008f
C1476 VTAIL.n484 VSUBS 0.01323f
C1477 VTAIL.n485 VSUBS 0.02462f
C1478 VTAIL.n486 VSUBS 0.02462f
C1479 VTAIL.n487 VSUBS 0.01323f
C1480 VTAIL.n488 VSUBS 0.014008f
C1481 VTAIL.n489 VSUBS 0.03127f
C1482 VTAIL.n490 VSUBS 0.03127f
C1483 VTAIL.n491 VSUBS 0.014008f
C1484 VTAIL.n492 VSUBS 0.01323f
C1485 VTAIL.n493 VSUBS 0.02462f
C1486 VTAIL.n494 VSUBS 0.02462f
C1487 VTAIL.n495 VSUBS 0.01323f
C1488 VTAIL.n496 VSUBS 0.014008f
C1489 VTAIL.n497 VSUBS 0.03127f
C1490 VTAIL.n498 VSUBS 0.03127f
C1491 VTAIL.n499 VSUBS 0.014008f
C1492 VTAIL.n500 VSUBS 0.01323f
C1493 VTAIL.n501 VSUBS 0.02462f
C1494 VTAIL.n502 VSUBS 0.02462f
C1495 VTAIL.n503 VSUBS 0.01323f
C1496 VTAIL.n504 VSUBS 0.014008f
C1497 VTAIL.n505 VSUBS 0.03127f
C1498 VTAIL.n506 VSUBS 0.078096f
C1499 VTAIL.n507 VSUBS 0.014008f
C1500 VTAIL.n508 VSUBS 0.02598f
C1501 VTAIL.n509 VSUBS 0.062625f
C1502 VTAIL.n510 VSUBS 0.060047f
C1503 VTAIL.n511 VSUBS 1.67791f
C1504 VTAIL.n512 VSUBS 0.026754f
C1505 VTAIL.n513 VSUBS 0.02462f
C1506 VTAIL.n514 VSUBS 0.01323f
C1507 VTAIL.n515 VSUBS 0.03127f
C1508 VTAIL.n516 VSUBS 0.014008f
C1509 VTAIL.n517 VSUBS 0.02462f
C1510 VTAIL.n518 VSUBS 0.01323f
C1511 VTAIL.n519 VSUBS 0.03127f
C1512 VTAIL.n520 VSUBS 0.014008f
C1513 VTAIL.n521 VSUBS 0.02462f
C1514 VTAIL.n522 VSUBS 0.01323f
C1515 VTAIL.n523 VSUBS 0.03127f
C1516 VTAIL.n524 VSUBS 0.014008f
C1517 VTAIL.n525 VSUBS 0.02462f
C1518 VTAIL.n526 VSUBS 0.01323f
C1519 VTAIL.n527 VSUBS 0.03127f
C1520 VTAIL.n528 VSUBS 0.014008f
C1521 VTAIL.n529 VSUBS 0.02462f
C1522 VTAIL.n530 VSUBS 0.01323f
C1523 VTAIL.n531 VSUBS 0.03127f
C1524 VTAIL.n532 VSUBS 0.014008f
C1525 VTAIL.n533 VSUBS 1.38984f
C1526 VTAIL.n534 VSUBS 0.01323f
C1527 VTAIL.t9 VSUBS 0.066844f
C1528 VTAIL.n535 VSUBS 0.161713f
C1529 VTAIL.n536 VSUBS 0.019893f
C1530 VTAIL.n537 VSUBS 0.023452f
C1531 VTAIL.n538 VSUBS 0.03127f
C1532 VTAIL.n539 VSUBS 0.014008f
C1533 VTAIL.n540 VSUBS 0.01323f
C1534 VTAIL.n541 VSUBS 0.02462f
C1535 VTAIL.n542 VSUBS 0.02462f
C1536 VTAIL.n543 VSUBS 0.01323f
C1537 VTAIL.n544 VSUBS 0.014008f
C1538 VTAIL.n545 VSUBS 0.03127f
C1539 VTAIL.n546 VSUBS 0.03127f
C1540 VTAIL.n547 VSUBS 0.014008f
C1541 VTAIL.n548 VSUBS 0.01323f
C1542 VTAIL.n549 VSUBS 0.02462f
C1543 VTAIL.n550 VSUBS 0.02462f
C1544 VTAIL.n551 VSUBS 0.01323f
C1545 VTAIL.n552 VSUBS 0.014008f
C1546 VTAIL.n553 VSUBS 0.03127f
C1547 VTAIL.n554 VSUBS 0.03127f
C1548 VTAIL.n555 VSUBS 0.014008f
C1549 VTAIL.n556 VSUBS 0.01323f
C1550 VTAIL.n557 VSUBS 0.02462f
C1551 VTAIL.n558 VSUBS 0.02462f
C1552 VTAIL.n559 VSUBS 0.01323f
C1553 VTAIL.n560 VSUBS 0.014008f
C1554 VTAIL.n561 VSUBS 0.03127f
C1555 VTAIL.n562 VSUBS 0.03127f
C1556 VTAIL.n563 VSUBS 0.014008f
C1557 VTAIL.n564 VSUBS 0.01323f
C1558 VTAIL.n565 VSUBS 0.02462f
C1559 VTAIL.n566 VSUBS 0.02462f
C1560 VTAIL.n567 VSUBS 0.01323f
C1561 VTAIL.n568 VSUBS 0.014008f
C1562 VTAIL.n569 VSUBS 0.03127f
C1563 VTAIL.n570 VSUBS 0.03127f
C1564 VTAIL.n571 VSUBS 0.014008f
C1565 VTAIL.n572 VSUBS 0.01323f
C1566 VTAIL.n573 VSUBS 0.02462f
C1567 VTAIL.n574 VSUBS 0.02462f
C1568 VTAIL.n575 VSUBS 0.01323f
C1569 VTAIL.n576 VSUBS 0.014008f
C1570 VTAIL.n577 VSUBS 0.03127f
C1571 VTAIL.n578 VSUBS 0.078096f
C1572 VTAIL.n579 VSUBS 0.014008f
C1573 VTAIL.n580 VSUBS 0.02598f
C1574 VTAIL.n581 VSUBS 0.062625f
C1575 VTAIL.n582 VSUBS 0.060047f
C1576 VTAIL.n583 VSUBS 1.67329f
C1577 VN.n0 VSUBS 0.037002f
C1578 VN.t4 VSUBS 2.69673f
C1579 VN.n1 VSUBS 0.044099f
C1580 VN.n2 VSUBS 0.028066f
C1581 VN.t5 VSUBS 2.69673f
C1582 VN.n3 VSUBS 0.94772f
C1583 VN.n4 VSUBS 0.028066f
C1584 VN.n5 VSUBS 0.040971f
C1585 VN.n6 VSUBS 0.272147f
C1586 VN.t0 VSUBS 2.69673f
C1587 VN.t6 VSUBS 2.93731f
C1588 VN.n7 VSUBS 1.00044f
C1589 VN.n8 VSUBS 1.02811f
C1590 VN.n9 VSUBS 0.038362f
C1591 VN.n10 VSUBS 0.052307f
C1592 VN.n11 VSUBS 0.028066f
C1593 VN.n12 VSUBS 0.028066f
C1594 VN.n13 VSUBS 0.028066f
C1595 VN.n14 VSUBS 0.040971f
C1596 VN.n15 VSUBS 0.052307f
C1597 VN.n16 VSUBS 0.038362f
C1598 VN.n17 VSUBS 0.028066f
C1599 VN.n18 VSUBS 0.028066f
C1600 VN.n19 VSUBS 0.040428f
C1601 VN.n20 VSUBS 0.052307f
C1602 VN.n21 VSUBS 0.037842f
C1603 VN.n22 VSUBS 0.028066f
C1604 VN.n23 VSUBS 0.028066f
C1605 VN.n24 VSUBS 0.028066f
C1606 VN.n25 VSUBS 0.052307f
C1607 VN.n26 VSUBS 0.036296f
C1608 VN.n27 VSUBS 1.04194f
C1609 VN.n28 VSUBS 0.046428f
C1610 VN.n29 VSUBS 0.037002f
C1611 VN.t7 VSUBS 2.69673f
C1612 VN.n30 VSUBS 0.044099f
C1613 VN.n31 VSUBS 0.028066f
C1614 VN.t1 VSUBS 2.69673f
C1615 VN.n32 VSUBS 0.94772f
C1616 VN.n33 VSUBS 0.028066f
C1617 VN.n34 VSUBS 0.040971f
C1618 VN.n35 VSUBS 0.272147f
C1619 VN.t2 VSUBS 2.69673f
C1620 VN.t3 VSUBS 2.93731f
C1621 VN.n36 VSUBS 1.00044f
C1622 VN.n37 VSUBS 1.02811f
C1623 VN.n38 VSUBS 0.038362f
C1624 VN.n39 VSUBS 0.052307f
C1625 VN.n40 VSUBS 0.028066f
C1626 VN.n41 VSUBS 0.028066f
C1627 VN.n42 VSUBS 0.028066f
C1628 VN.n43 VSUBS 0.040971f
C1629 VN.n44 VSUBS 0.052307f
C1630 VN.n45 VSUBS 0.038362f
C1631 VN.n46 VSUBS 0.028066f
C1632 VN.n47 VSUBS 0.028066f
C1633 VN.n48 VSUBS 0.040428f
C1634 VN.n49 VSUBS 0.052307f
C1635 VN.n50 VSUBS 0.037842f
C1636 VN.n51 VSUBS 0.028066f
C1637 VN.n52 VSUBS 0.028066f
C1638 VN.n53 VSUBS 0.028066f
C1639 VN.n54 VSUBS 0.052307f
C1640 VN.n55 VSUBS 0.036296f
C1641 VN.n56 VSUBS 1.04194f
C1642 VN.n57 VSUBS 1.67347f
.ends

