* NGSPICE file created from diff_pair_sample_0598.ext - technology: sky130A

.subckt diff_pair_sample_0598 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=2.59
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=2.59
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=2.59
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=1.9188 ps=10.62 w=4.92 l=2.59
X4 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=1.9188 ps=10.62 w=4.92 l=2.59
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=0 ps=0 w=4.92 l=2.59
X6 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=1.9188 ps=10.62 w=4.92 l=2.59
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9188 pd=10.62 as=1.9188 ps=10.62 w=4.92 l=2.59
R0 B.n469 B.n468 585
R1 B.n470 B.n469 585
R2 B.n179 B.n74 585
R3 B.n178 B.n177 585
R4 B.n176 B.n175 585
R5 B.n174 B.n173 585
R6 B.n172 B.n171 585
R7 B.n170 B.n169 585
R8 B.n168 B.n167 585
R9 B.n166 B.n165 585
R10 B.n164 B.n163 585
R11 B.n162 B.n161 585
R12 B.n160 B.n159 585
R13 B.n158 B.n157 585
R14 B.n156 B.n155 585
R15 B.n154 B.n153 585
R16 B.n152 B.n151 585
R17 B.n150 B.n149 585
R18 B.n148 B.n147 585
R19 B.n146 B.n145 585
R20 B.n144 B.n143 585
R21 B.n142 B.n141 585
R22 B.n140 B.n139 585
R23 B.n138 B.n137 585
R24 B.n136 B.n135 585
R25 B.n134 B.n133 585
R26 B.n132 B.n131 585
R27 B.n130 B.n129 585
R28 B.n128 B.n127 585
R29 B.n126 B.n125 585
R30 B.n124 B.n123 585
R31 B.n121 B.n120 585
R32 B.n119 B.n118 585
R33 B.n117 B.n116 585
R34 B.n115 B.n114 585
R35 B.n113 B.n112 585
R36 B.n111 B.n110 585
R37 B.n109 B.n108 585
R38 B.n107 B.n106 585
R39 B.n105 B.n104 585
R40 B.n103 B.n102 585
R41 B.n101 B.n100 585
R42 B.n99 B.n98 585
R43 B.n97 B.n96 585
R44 B.n95 B.n94 585
R45 B.n93 B.n92 585
R46 B.n91 B.n90 585
R47 B.n89 B.n88 585
R48 B.n87 B.n86 585
R49 B.n85 B.n84 585
R50 B.n83 B.n82 585
R51 B.n81 B.n80 585
R52 B.n467 B.n48 585
R53 B.n471 B.n48 585
R54 B.n466 B.n47 585
R55 B.n472 B.n47 585
R56 B.n465 B.n464 585
R57 B.n464 B.n43 585
R58 B.n463 B.n42 585
R59 B.n478 B.n42 585
R60 B.n462 B.n41 585
R61 B.n479 B.n41 585
R62 B.n461 B.n40 585
R63 B.n480 B.n40 585
R64 B.n460 B.n459 585
R65 B.n459 B.n36 585
R66 B.n458 B.n35 585
R67 B.n486 B.n35 585
R68 B.n457 B.n34 585
R69 B.n487 B.n34 585
R70 B.n456 B.n33 585
R71 B.n488 B.n33 585
R72 B.n455 B.n454 585
R73 B.n454 B.n29 585
R74 B.n453 B.n28 585
R75 B.n494 B.n28 585
R76 B.n452 B.n27 585
R77 B.n495 B.n27 585
R78 B.n451 B.n26 585
R79 B.n496 B.n26 585
R80 B.n450 B.n449 585
R81 B.n449 B.n22 585
R82 B.n448 B.n21 585
R83 B.n502 B.n21 585
R84 B.n447 B.n20 585
R85 B.n503 B.n20 585
R86 B.n446 B.n19 585
R87 B.n504 B.n19 585
R88 B.n445 B.n444 585
R89 B.n444 B.n15 585
R90 B.n443 B.n14 585
R91 B.n510 B.n14 585
R92 B.n442 B.n13 585
R93 B.n511 B.n13 585
R94 B.n441 B.n12 585
R95 B.n512 B.n12 585
R96 B.n440 B.n439 585
R97 B.n439 B.n8 585
R98 B.n438 B.n7 585
R99 B.n518 B.n7 585
R100 B.n437 B.n6 585
R101 B.n519 B.n6 585
R102 B.n436 B.n5 585
R103 B.n520 B.n5 585
R104 B.n435 B.n434 585
R105 B.n434 B.n4 585
R106 B.n433 B.n180 585
R107 B.n433 B.n432 585
R108 B.n423 B.n181 585
R109 B.n182 B.n181 585
R110 B.n425 B.n424 585
R111 B.n426 B.n425 585
R112 B.n422 B.n187 585
R113 B.n187 B.n186 585
R114 B.n421 B.n420 585
R115 B.n420 B.n419 585
R116 B.n189 B.n188 585
R117 B.n190 B.n189 585
R118 B.n412 B.n411 585
R119 B.n413 B.n412 585
R120 B.n410 B.n195 585
R121 B.n195 B.n194 585
R122 B.n409 B.n408 585
R123 B.n408 B.n407 585
R124 B.n197 B.n196 585
R125 B.n198 B.n197 585
R126 B.n400 B.n399 585
R127 B.n401 B.n400 585
R128 B.n398 B.n203 585
R129 B.n203 B.n202 585
R130 B.n397 B.n396 585
R131 B.n396 B.n395 585
R132 B.n205 B.n204 585
R133 B.n206 B.n205 585
R134 B.n388 B.n387 585
R135 B.n389 B.n388 585
R136 B.n386 B.n211 585
R137 B.n211 B.n210 585
R138 B.n385 B.n384 585
R139 B.n384 B.n383 585
R140 B.n213 B.n212 585
R141 B.n214 B.n213 585
R142 B.n376 B.n375 585
R143 B.n377 B.n376 585
R144 B.n374 B.n219 585
R145 B.n219 B.n218 585
R146 B.n373 B.n372 585
R147 B.n372 B.n371 585
R148 B.n221 B.n220 585
R149 B.n222 B.n221 585
R150 B.n364 B.n363 585
R151 B.n365 B.n364 585
R152 B.n362 B.n227 585
R153 B.n227 B.n226 585
R154 B.n356 B.n355 585
R155 B.n354 B.n254 585
R156 B.n353 B.n253 585
R157 B.n358 B.n253 585
R158 B.n352 B.n351 585
R159 B.n350 B.n349 585
R160 B.n348 B.n347 585
R161 B.n346 B.n345 585
R162 B.n344 B.n343 585
R163 B.n342 B.n341 585
R164 B.n340 B.n339 585
R165 B.n338 B.n337 585
R166 B.n336 B.n335 585
R167 B.n334 B.n333 585
R168 B.n332 B.n331 585
R169 B.n330 B.n329 585
R170 B.n328 B.n327 585
R171 B.n326 B.n325 585
R172 B.n324 B.n323 585
R173 B.n322 B.n321 585
R174 B.n320 B.n319 585
R175 B.n318 B.n317 585
R176 B.n316 B.n315 585
R177 B.n314 B.n313 585
R178 B.n312 B.n311 585
R179 B.n310 B.n309 585
R180 B.n308 B.n307 585
R181 B.n306 B.n305 585
R182 B.n304 B.n303 585
R183 B.n302 B.n301 585
R184 B.n300 B.n299 585
R185 B.n297 B.n296 585
R186 B.n295 B.n294 585
R187 B.n293 B.n292 585
R188 B.n291 B.n290 585
R189 B.n289 B.n288 585
R190 B.n287 B.n286 585
R191 B.n285 B.n284 585
R192 B.n283 B.n282 585
R193 B.n281 B.n280 585
R194 B.n279 B.n278 585
R195 B.n277 B.n276 585
R196 B.n275 B.n274 585
R197 B.n273 B.n272 585
R198 B.n271 B.n270 585
R199 B.n269 B.n268 585
R200 B.n267 B.n266 585
R201 B.n265 B.n264 585
R202 B.n263 B.n262 585
R203 B.n261 B.n260 585
R204 B.n229 B.n228 585
R205 B.n361 B.n360 585
R206 B.n225 B.n224 585
R207 B.n226 B.n225 585
R208 B.n367 B.n366 585
R209 B.n366 B.n365 585
R210 B.n368 B.n223 585
R211 B.n223 B.n222 585
R212 B.n370 B.n369 585
R213 B.n371 B.n370 585
R214 B.n217 B.n216 585
R215 B.n218 B.n217 585
R216 B.n379 B.n378 585
R217 B.n378 B.n377 585
R218 B.n380 B.n215 585
R219 B.n215 B.n214 585
R220 B.n382 B.n381 585
R221 B.n383 B.n382 585
R222 B.n209 B.n208 585
R223 B.n210 B.n209 585
R224 B.n391 B.n390 585
R225 B.n390 B.n389 585
R226 B.n392 B.n207 585
R227 B.n207 B.n206 585
R228 B.n394 B.n393 585
R229 B.n395 B.n394 585
R230 B.n201 B.n200 585
R231 B.n202 B.n201 585
R232 B.n403 B.n402 585
R233 B.n402 B.n401 585
R234 B.n404 B.n199 585
R235 B.n199 B.n198 585
R236 B.n406 B.n405 585
R237 B.n407 B.n406 585
R238 B.n193 B.n192 585
R239 B.n194 B.n193 585
R240 B.n415 B.n414 585
R241 B.n414 B.n413 585
R242 B.n416 B.n191 585
R243 B.n191 B.n190 585
R244 B.n418 B.n417 585
R245 B.n419 B.n418 585
R246 B.n185 B.n184 585
R247 B.n186 B.n185 585
R248 B.n428 B.n427 585
R249 B.n427 B.n426 585
R250 B.n429 B.n183 585
R251 B.n183 B.n182 585
R252 B.n431 B.n430 585
R253 B.n432 B.n431 585
R254 B.n2 B.n0 585
R255 B.n4 B.n2 585
R256 B.n3 B.n1 585
R257 B.n519 B.n3 585
R258 B.n517 B.n516 585
R259 B.n518 B.n517 585
R260 B.n515 B.n9 585
R261 B.n9 B.n8 585
R262 B.n514 B.n513 585
R263 B.n513 B.n512 585
R264 B.n11 B.n10 585
R265 B.n511 B.n11 585
R266 B.n509 B.n508 585
R267 B.n510 B.n509 585
R268 B.n507 B.n16 585
R269 B.n16 B.n15 585
R270 B.n506 B.n505 585
R271 B.n505 B.n504 585
R272 B.n18 B.n17 585
R273 B.n503 B.n18 585
R274 B.n501 B.n500 585
R275 B.n502 B.n501 585
R276 B.n499 B.n23 585
R277 B.n23 B.n22 585
R278 B.n498 B.n497 585
R279 B.n497 B.n496 585
R280 B.n25 B.n24 585
R281 B.n495 B.n25 585
R282 B.n493 B.n492 585
R283 B.n494 B.n493 585
R284 B.n491 B.n30 585
R285 B.n30 B.n29 585
R286 B.n490 B.n489 585
R287 B.n489 B.n488 585
R288 B.n32 B.n31 585
R289 B.n487 B.n32 585
R290 B.n485 B.n484 585
R291 B.n486 B.n485 585
R292 B.n483 B.n37 585
R293 B.n37 B.n36 585
R294 B.n482 B.n481 585
R295 B.n481 B.n480 585
R296 B.n39 B.n38 585
R297 B.n479 B.n39 585
R298 B.n477 B.n476 585
R299 B.n478 B.n477 585
R300 B.n475 B.n44 585
R301 B.n44 B.n43 585
R302 B.n474 B.n473 585
R303 B.n473 B.n472 585
R304 B.n46 B.n45 585
R305 B.n471 B.n46 585
R306 B.n522 B.n521 585
R307 B.n521 B.n520 585
R308 B.n356 B.n225 559.769
R309 B.n80 B.n46 559.769
R310 B.n360 B.n227 559.769
R311 B.n469 B.n48 559.769
R312 B.n470 B.n73 256.663
R313 B.n470 B.n72 256.663
R314 B.n470 B.n71 256.663
R315 B.n470 B.n70 256.663
R316 B.n470 B.n69 256.663
R317 B.n470 B.n68 256.663
R318 B.n470 B.n67 256.663
R319 B.n470 B.n66 256.663
R320 B.n470 B.n65 256.663
R321 B.n470 B.n64 256.663
R322 B.n470 B.n63 256.663
R323 B.n470 B.n62 256.663
R324 B.n470 B.n61 256.663
R325 B.n470 B.n60 256.663
R326 B.n470 B.n59 256.663
R327 B.n470 B.n58 256.663
R328 B.n470 B.n57 256.663
R329 B.n470 B.n56 256.663
R330 B.n470 B.n55 256.663
R331 B.n470 B.n54 256.663
R332 B.n470 B.n53 256.663
R333 B.n470 B.n52 256.663
R334 B.n470 B.n51 256.663
R335 B.n470 B.n50 256.663
R336 B.n470 B.n49 256.663
R337 B.n358 B.n357 256.663
R338 B.n358 B.n230 256.663
R339 B.n358 B.n231 256.663
R340 B.n358 B.n232 256.663
R341 B.n358 B.n233 256.663
R342 B.n358 B.n234 256.663
R343 B.n358 B.n235 256.663
R344 B.n358 B.n236 256.663
R345 B.n358 B.n237 256.663
R346 B.n358 B.n238 256.663
R347 B.n358 B.n239 256.663
R348 B.n358 B.n240 256.663
R349 B.n358 B.n241 256.663
R350 B.n358 B.n242 256.663
R351 B.n358 B.n243 256.663
R352 B.n358 B.n244 256.663
R353 B.n358 B.n245 256.663
R354 B.n358 B.n246 256.663
R355 B.n358 B.n247 256.663
R356 B.n358 B.n248 256.663
R357 B.n358 B.n249 256.663
R358 B.n358 B.n250 256.663
R359 B.n358 B.n251 256.663
R360 B.n358 B.n252 256.663
R361 B.n359 B.n358 256.663
R362 B.n258 B.t6 253.812
R363 B.n255 B.t2 253.812
R364 B.n78 B.t9 253.812
R365 B.n75 B.t13 253.812
R366 B.n366 B.n225 163.367
R367 B.n366 B.n223 163.367
R368 B.n370 B.n223 163.367
R369 B.n370 B.n217 163.367
R370 B.n378 B.n217 163.367
R371 B.n378 B.n215 163.367
R372 B.n382 B.n215 163.367
R373 B.n382 B.n209 163.367
R374 B.n390 B.n209 163.367
R375 B.n390 B.n207 163.367
R376 B.n394 B.n207 163.367
R377 B.n394 B.n201 163.367
R378 B.n402 B.n201 163.367
R379 B.n402 B.n199 163.367
R380 B.n406 B.n199 163.367
R381 B.n406 B.n193 163.367
R382 B.n414 B.n193 163.367
R383 B.n414 B.n191 163.367
R384 B.n418 B.n191 163.367
R385 B.n418 B.n185 163.367
R386 B.n427 B.n185 163.367
R387 B.n427 B.n183 163.367
R388 B.n431 B.n183 163.367
R389 B.n431 B.n2 163.367
R390 B.n521 B.n2 163.367
R391 B.n521 B.n3 163.367
R392 B.n517 B.n3 163.367
R393 B.n517 B.n9 163.367
R394 B.n513 B.n9 163.367
R395 B.n513 B.n11 163.367
R396 B.n509 B.n11 163.367
R397 B.n509 B.n16 163.367
R398 B.n505 B.n16 163.367
R399 B.n505 B.n18 163.367
R400 B.n501 B.n18 163.367
R401 B.n501 B.n23 163.367
R402 B.n497 B.n23 163.367
R403 B.n497 B.n25 163.367
R404 B.n493 B.n25 163.367
R405 B.n493 B.n30 163.367
R406 B.n489 B.n30 163.367
R407 B.n489 B.n32 163.367
R408 B.n485 B.n32 163.367
R409 B.n485 B.n37 163.367
R410 B.n481 B.n37 163.367
R411 B.n481 B.n39 163.367
R412 B.n477 B.n39 163.367
R413 B.n477 B.n44 163.367
R414 B.n473 B.n44 163.367
R415 B.n473 B.n46 163.367
R416 B.n254 B.n253 163.367
R417 B.n351 B.n253 163.367
R418 B.n349 B.n348 163.367
R419 B.n345 B.n344 163.367
R420 B.n341 B.n340 163.367
R421 B.n337 B.n336 163.367
R422 B.n333 B.n332 163.367
R423 B.n329 B.n328 163.367
R424 B.n325 B.n324 163.367
R425 B.n321 B.n320 163.367
R426 B.n317 B.n316 163.367
R427 B.n313 B.n312 163.367
R428 B.n309 B.n308 163.367
R429 B.n305 B.n304 163.367
R430 B.n301 B.n300 163.367
R431 B.n296 B.n295 163.367
R432 B.n292 B.n291 163.367
R433 B.n288 B.n287 163.367
R434 B.n284 B.n283 163.367
R435 B.n280 B.n279 163.367
R436 B.n276 B.n275 163.367
R437 B.n272 B.n271 163.367
R438 B.n268 B.n267 163.367
R439 B.n264 B.n263 163.367
R440 B.n260 B.n229 163.367
R441 B.n364 B.n227 163.367
R442 B.n364 B.n221 163.367
R443 B.n372 B.n221 163.367
R444 B.n372 B.n219 163.367
R445 B.n376 B.n219 163.367
R446 B.n376 B.n213 163.367
R447 B.n384 B.n213 163.367
R448 B.n384 B.n211 163.367
R449 B.n388 B.n211 163.367
R450 B.n388 B.n205 163.367
R451 B.n396 B.n205 163.367
R452 B.n396 B.n203 163.367
R453 B.n400 B.n203 163.367
R454 B.n400 B.n197 163.367
R455 B.n408 B.n197 163.367
R456 B.n408 B.n195 163.367
R457 B.n412 B.n195 163.367
R458 B.n412 B.n189 163.367
R459 B.n420 B.n189 163.367
R460 B.n420 B.n187 163.367
R461 B.n425 B.n187 163.367
R462 B.n425 B.n181 163.367
R463 B.n433 B.n181 163.367
R464 B.n434 B.n433 163.367
R465 B.n434 B.n5 163.367
R466 B.n6 B.n5 163.367
R467 B.n7 B.n6 163.367
R468 B.n439 B.n7 163.367
R469 B.n439 B.n12 163.367
R470 B.n13 B.n12 163.367
R471 B.n14 B.n13 163.367
R472 B.n444 B.n14 163.367
R473 B.n444 B.n19 163.367
R474 B.n20 B.n19 163.367
R475 B.n21 B.n20 163.367
R476 B.n449 B.n21 163.367
R477 B.n449 B.n26 163.367
R478 B.n27 B.n26 163.367
R479 B.n28 B.n27 163.367
R480 B.n454 B.n28 163.367
R481 B.n454 B.n33 163.367
R482 B.n34 B.n33 163.367
R483 B.n35 B.n34 163.367
R484 B.n459 B.n35 163.367
R485 B.n459 B.n40 163.367
R486 B.n41 B.n40 163.367
R487 B.n42 B.n41 163.367
R488 B.n464 B.n42 163.367
R489 B.n464 B.n47 163.367
R490 B.n48 B.n47 163.367
R491 B.n84 B.n83 163.367
R492 B.n88 B.n87 163.367
R493 B.n92 B.n91 163.367
R494 B.n96 B.n95 163.367
R495 B.n100 B.n99 163.367
R496 B.n104 B.n103 163.367
R497 B.n108 B.n107 163.367
R498 B.n112 B.n111 163.367
R499 B.n116 B.n115 163.367
R500 B.n120 B.n119 163.367
R501 B.n125 B.n124 163.367
R502 B.n129 B.n128 163.367
R503 B.n133 B.n132 163.367
R504 B.n137 B.n136 163.367
R505 B.n141 B.n140 163.367
R506 B.n145 B.n144 163.367
R507 B.n149 B.n148 163.367
R508 B.n153 B.n152 163.367
R509 B.n157 B.n156 163.367
R510 B.n161 B.n160 163.367
R511 B.n165 B.n164 163.367
R512 B.n169 B.n168 163.367
R513 B.n173 B.n172 163.367
R514 B.n177 B.n176 163.367
R515 B.n469 B.n74 163.367
R516 B.n358 B.n226 154.292
R517 B.n471 B.n470 154.292
R518 B.n258 B.t8 129.986
R519 B.n75 B.t14 129.986
R520 B.n255 B.t5 129.981
R521 B.n78 B.t11 129.981
R522 B.n365 B.n226 73.3698
R523 B.n365 B.n222 73.3698
R524 B.n371 B.n222 73.3698
R525 B.n371 B.n218 73.3698
R526 B.n377 B.n218 73.3698
R527 B.n377 B.n214 73.3698
R528 B.n383 B.n214 73.3698
R529 B.n389 B.n210 73.3698
R530 B.n389 B.n206 73.3698
R531 B.n395 B.n206 73.3698
R532 B.n395 B.n202 73.3698
R533 B.n401 B.n202 73.3698
R534 B.n401 B.n198 73.3698
R535 B.n407 B.n198 73.3698
R536 B.n407 B.n194 73.3698
R537 B.n413 B.n194 73.3698
R538 B.n413 B.n190 73.3698
R539 B.n419 B.n190 73.3698
R540 B.n426 B.n186 73.3698
R541 B.n426 B.n182 73.3698
R542 B.n432 B.n182 73.3698
R543 B.n432 B.n4 73.3698
R544 B.n520 B.n4 73.3698
R545 B.n520 B.n519 73.3698
R546 B.n519 B.n518 73.3698
R547 B.n518 B.n8 73.3698
R548 B.n512 B.n8 73.3698
R549 B.n512 B.n511 73.3698
R550 B.n510 B.n15 73.3698
R551 B.n504 B.n15 73.3698
R552 B.n504 B.n503 73.3698
R553 B.n503 B.n502 73.3698
R554 B.n502 B.n22 73.3698
R555 B.n496 B.n22 73.3698
R556 B.n496 B.n495 73.3698
R557 B.n495 B.n494 73.3698
R558 B.n494 B.n29 73.3698
R559 B.n488 B.n29 73.3698
R560 B.n488 B.n487 73.3698
R561 B.n486 B.n36 73.3698
R562 B.n480 B.n36 73.3698
R563 B.n480 B.n479 73.3698
R564 B.n479 B.n478 73.3698
R565 B.n478 B.n43 73.3698
R566 B.n472 B.n43 73.3698
R567 B.n472 B.n471 73.3698
R568 B.n259 B.t7 73.3553
R569 B.n76 B.t15 73.3553
R570 B.n256 B.t4 73.3505
R571 B.n79 B.t12 73.3505
R572 B.n357 B.n356 71.676
R573 B.n351 B.n230 71.676
R574 B.n348 B.n231 71.676
R575 B.n344 B.n232 71.676
R576 B.n340 B.n233 71.676
R577 B.n336 B.n234 71.676
R578 B.n332 B.n235 71.676
R579 B.n328 B.n236 71.676
R580 B.n324 B.n237 71.676
R581 B.n320 B.n238 71.676
R582 B.n316 B.n239 71.676
R583 B.n312 B.n240 71.676
R584 B.n308 B.n241 71.676
R585 B.n304 B.n242 71.676
R586 B.n300 B.n243 71.676
R587 B.n295 B.n244 71.676
R588 B.n291 B.n245 71.676
R589 B.n287 B.n246 71.676
R590 B.n283 B.n247 71.676
R591 B.n279 B.n248 71.676
R592 B.n275 B.n249 71.676
R593 B.n271 B.n250 71.676
R594 B.n267 B.n251 71.676
R595 B.n263 B.n252 71.676
R596 B.n359 B.n229 71.676
R597 B.n80 B.n49 71.676
R598 B.n84 B.n50 71.676
R599 B.n88 B.n51 71.676
R600 B.n92 B.n52 71.676
R601 B.n96 B.n53 71.676
R602 B.n100 B.n54 71.676
R603 B.n104 B.n55 71.676
R604 B.n108 B.n56 71.676
R605 B.n112 B.n57 71.676
R606 B.n116 B.n58 71.676
R607 B.n120 B.n59 71.676
R608 B.n125 B.n60 71.676
R609 B.n129 B.n61 71.676
R610 B.n133 B.n62 71.676
R611 B.n137 B.n63 71.676
R612 B.n141 B.n64 71.676
R613 B.n145 B.n65 71.676
R614 B.n149 B.n66 71.676
R615 B.n153 B.n67 71.676
R616 B.n157 B.n68 71.676
R617 B.n161 B.n69 71.676
R618 B.n165 B.n70 71.676
R619 B.n169 B.n71 71.676
R620 B.n173 B.n72 71.676
R621 B.n177 B.n73 71.676
R622 B.n74 B.n73 71.676
R623 B.n176 B.n72 71.676
R624 B.n172 B.n71 71.676
R625 B.n168 B.n70 71.676
R626 B.n164 B.n69 71.676
R627 B.n160 B.n68 71.676
R628 B.n156 B.n67 71.676
R629 B.n152 B.n66 71.676
R630 B.n148 B.n65 71.676
R631 B.n144 B.n64 71.676
R632 B.n140 B.n63 71.676
R633 B.n136 B.n62 71.676
R634 B.n132 B.n61 71.676
R635 B.n128 B.n60 71.676
R636 B.n124 B.n59 71.676
R637 B.n119 B.n58 71.676
R638 B.n115 B.n57 71.676
R639 B.n111 B.n56 71.676
R640 B.n107 B.n55 71.676
R641 B.n103 B.n54 71.676
R642 B.n99 B.n53 71.676
R643 B.n95 B.n52 71.676
R644 B.n91 B.n51 71.676
R645 B.n87 B.n50 71.676
R646 B.n83 B.n49 71.676
R647 B.n357 B.n254 71.676
R648 B.n349 B.n230 71.676
R649 B.n345 B.n231 71.676
R650 B.n341 B.n232 71.676
R651 B.n337 B.n233 71.676
R652 B.n333 B.n234 71.676
R653 B.n329 B.n235 71.676
R654 B.n325 B.n236 71.676
R655 B.n321 B.n237 71.676
R656 B.n317 B.n238 71.676
R657 B.n313 B.n239 71.676
R658 B.n309 B.n240 71.676
R659 B.n305 B.n241 71.676
R660 B.n301 B.n242 71.676
R661 B.n296 B.n243 71.676
R662 B.n292 B.n244 71.676
R663 B.n288 B.n245 71.676
R664 B.n284 B.n246 71.676
R665 B.n280 B.n247 71.676
R666 B.n276 B.n248 71.676
R667 B.n272 B.n249 71.676
R668 B.n268 B.n250 71.676
R669 B.n264 B.n251 71.676
R670 B.n260 B.n252 71.676
R671 B.n360 B.n359 71.676
R672 B.t1 B.n186 65.8171
R673 B.n511 B.t0 65.8171
R674 B.n298 B.n259 59.5399
R675 B.n257 B.n256 59.5399
R676 B.n122 B.n79 59.5399
R677 B.n77 B.n76 59.5399
R678 B.n259 B.n258 56.6308
R679 B.n256 B.n255 56.6308
R680 B.n79 B.n78 56.6308
R681 B.n76 B.n75 56.6308
R682 B.t3 B.n210 50.7116
R683 B.n487 B.t10 50.7116
R684 B.n468 B.n467 36.3712
R685 B.n81 B.n45 36.3712
R686 B.n362 B.n361 36.3712
R687 B.n355 B.n224 36.3712
R688 B.n383 B.t3 22.6587
R689 B.t10 B.n486 22.6587
R690 B B.n522 18.0485
R691 B.n82 B.n81 10.6151
R692 B.n85 B.n82 10.6151
R693 B.n86 B.n85 10.6151
R694 B.n89 B.n86 10.6151
R695 B.n90 B.n89 10.6151
R696 B.n93 B.n90 10.6151
R697 B.n94 B.n93 10.6151
R698 B.n97 B.n94 10.6151
R699 B.n98 B.n97 10.6151
R700 B.n101 B.n98 10.6151
R701 B.n102 B.n101 10.6151
R702 B.n105 B.n102 10.6151
R703 B.n106 B.n105 10.6151
R704 B.n109 B.n106 10.6151
R705 B.n110 B.n109 10.6151
R706 B.n113 B.n110 10.6151
R707 B.n114 B.n113 10.6151
R708 B.n117 B.n114 10.6151
R709 B.n118 B.n117 10.6151
R710 B.n121 B.n118 10.6151
R711 B.n126 B.n123 10.6151
R712 B.n127 B.n126 10.6151
R713 B.n130 B.n127 10.6151
R714 B.n131 B.n130 10.6151
R715 B.n134 B.n131 10.6151
R716 B.n135 B.n134 10.6151
R717 B.n138 B.n135 10.6151
R718 B.n139 B.n138 10.6151
R719 B.n143 B.n142 10.6151
R720 B.n146 B.n143 10.6151
R721 B.n147 B.n146 10.6151
R722 B.n150 B.n147 10.6151
R723 B.n151 B.n150 10.6151
R724 B.n154 B.n151 10.6151
R725 B.n155 B.n154 10.6151
R726 B.n158 B.n155 10.6151
R727 B.n159 B.n158 10.6151
R728 B.n162 B.n159 10.6151
R729 B.n163 B.n162 10.6151
R730 B.n166 B.n163 10.6151
R731 B.n167 B.n166 10.6151
R732 B.n170 B.n167 10.6151
R733 B.n171 B.n170 10.6151
R734 B.n174 B.n171 10.6151
R735 B.n175 B.n174 10.6151
R736 B.n178 B.n175 10.6151
R737 B.n179 B.n178 10.6151
R738 B.n468 B.n179 10.6151
R739 B.n363 B.n362 10.6151
R740 B.n363 B.n220 10.6151
R741 B.n373 B.n220 10.6151
R742 B.n374 B.n373 10.6151
R743 B.n375 B.n374 10.6151
R744 B.n375 B.n212 10.6151
R745 B.n385 B.n212 10.6151
R746 B.n386 B.n385 10.6151
R747 B.n387 B.n386 10.6151
R748 B.n387 B.n204 10.6151
R749 B.n397 B.n204 10.6151
R750 B.n398 B.n397 10.6151
R751 B.n399 B.n398 10.6151
R752 B.n399 B.n196 10.6151
R753 B.n409 B.n196 10.6151
R754 B.n410 B.n409 10.6151
R755 B.n411 B.n410 10.6151
R756 B.n411 B.n188 10.6151
R757 B.n421 B.n188 10.6151
R758 B.n422 B.n421 10.6151
R759 B.n424 B.n422 10.6151
R760 B.n424 B.n423 10.6151
R761 B.n423 B.n180 10.6151
R762 B.n435 B.n180 10.6151
R763 B.n436 B.n435 10.6151
R764 B.n437 B.n436 10.6151
R765 B.n438 B.n437 10.6151
R766 B.n440 B.n438 10.6151
R767 B.n441 B.n440 10.6151
R768 B.n442 B.n441 10.6151
R769 B.n443 B.n442 10.6151
R770 B.n445 B.n443 10.6151
R771 B.n446 B.n445 10.6151
R772 B.n447 B.n446 10.6151
R773 B.n448 B.n447 10.6151
R774 B.n450 B.n448 10.6151
R775 B.n451 B.n450 10.6151
R776 B.n452 B.n451 10.6151
R777 B.n453 B.n452 10.6151
R778 B.n455 B.n453 10.6151
R779 B.n456 B.n455 10.6151
R780 B.n457 B.n456 10.6151
R781 B.n458 B.n457 10.6151
R782 B.n460 B.n458 10.6151
R783 B.n461 B.n460 10.6151
R784 B.n462 B.n461 10.6151
R785 B.n463 B.n462 10.6151
R786 B.n465 B.n463 10.6151
R787 B.n466 B.n465 10.6151
R788 B.n467 B.n466 10.6151
R789 B.n355 B.n354 10.6151
R790 B.n354 B.n353 10.6151
R791 B.n353 B.n352 10.6151
R792 B.n352 B.n350 10.6151
R793 B.n350 B.n347 10.6151
R794 B.n347 B.n346 10.6151
R795 B.n346 B.n343 10.6151
R796 B.n343 B.n342 10.6151
R797 B.n342 B.n339 10.6151
R798 B.n339 B.n338 10.6151
R799 B.n338 B.n335 10.6151
R800 B.n335 B.n334 10.6151
R801 B.n334 B.n331 10.6151
R802 B.n331 B.n330 10.6151
R803 B.n330 B.n327 10.6151
R804 B.n327 B.n326 10.6151
R805 B.n326 B.n323 10.6151
R806 B.n323 B.n322 10.6151
R807 B.n322 B.n319 10.6151
R808 B.n319 B.n318 10.6151
R809 B.n315 B.n314 10.6151
R810 B.n314 B.n311 10.6151
R811 B.n311 B.n310 10.6151
R812 B.n310 B.n307 10.6151
R813 B.n307 B.n306 10.6151
R814 B.n306 B.n303 10.6151
R815 B.n303 B.n302 10.6151
R816 B.n302 B.n299 10.6151
R817 B.n297 B.n294 10.6151
R818 B.n294 B.n293 10.6151
R819 B.n293 B.n290 10.6151
R820 B.n290 B.n289 10.6151
R821 B.n289 B.n286 10.6151
R822 B.n286 B.n285 10.6151
R823 B.n285 B.n282 10.6151
R824 B.n282 B.n281 10.6151
R825 B.n281 B.n278 10.6151
R826 B.n278 B.n277 10.6151
R827 B.n277 B.n274 10.6151
R828 B.n274 B.n273 10.6151
R829 B.n273 B.n270 10.6151
R830 B.n270 B.n269 10.6151
R831 B.n269 B.n266 10.6151
R832 B.n266 B.n265 10.6151
R833 B.n265 B.n262 10.6151
R834 B.n262 B.n261 10.6151
R835 B.n261 B.n228 10.6151
R836 B.n361 B.n228 10.6151
R837 B.n367 B.n224 10.6151
R838 B.n368 B.n367 10.6151
R839 B.n369 B.n368 10.6151
R840 B.n369 B.n216 10.6151
R841 B.n379 B.n216 10.6151
R842 B.n380 B.n379 10.6151
R843 B.n381 B.n380 10.6151
R844 B.n381 B.n208 10.6151
R845 B.n391 B.n208 10.6151
R846 B.n392 B.n391 10.6151
R847 B.n393 B.n392 10.6151
R848 B.n393 B.n200 10.6151
R849 B.n403 B.n200 10.6151
R850 B.n404 B.n403 10.6151
R851 B.n405 B.n404 10.6151
R852 B.n405 B.n192 10.6151
R853 B.n415 B.n192 10.6151
R854 B.n416 B.n415 10.6151
R855 B.n417 B.n416 10.6151
R856 B.n417 B.n184 10.6151
R857 B.n428 B.n184 10.6151
R858 B.n429 B.n428 10.6151
R859 B.n430 B.n429 10.6151
R860 B.n430 B.n0 10.6151
R861 B.n516 B.n1 10.6151
R862 B.n516 B.n515 10.6151
R863 B.n515 B.n514 10.6151
R864 B.n514 B.n10 10.6151
R865 B.n508 B.n10 10.6151
R866 B.n508 B.n507 10.6151
R867 B.n507 B.n506 10.6151
R868 B.n506 B.n17 10.6151
R869 B.n500 B.n17 10.6151
R870 B.n500 B.n499 10.6151
R871 B.n499 B.n498 10.6151
R872 B.n498 B.n24 10.6151
R873 B.n492 B.n24 10.6151
R874 B.n492 B.n491 10.6151
R875 B.n491 B.n490 10.6151
R876 B.n490 B.n31 10.6151
R877 B.n484 B.n31 10.6151
R878 B.n484 B.n483 10.6151
R879 B.n483 B.n482 10.6151
R880 B.n482 B.n38 10.6151
R881 B.n476 B.n38 10.6151
R882 B.n476 B.n475 10.6151
R883 B.n475 B.n474 10.6151
R884 B.n474 B.n45 10.6151
R885 B.n419 B.t1 7.55322
R886 B.t0 B.n510 7.55322
R887 B.n123 B.n122 6.5566
R888 B.n139 B.n77 6.5566
R889 B.n315 B.n257 6.5566
R890 B.n299 B.n298 6.5566
R891 B.n122 B.n121 4.05904
R892 B.n142 B.n77 4.05904
R893 B.n318 B.n257 4.05904
R894 B.n298 B.n297 4.05904
R895 B.n522 B.n0 2.81026
R896 B.n522 B.n1 2.81026
R897 VP.n0 VP.t0 134.262
R898 VP.n0 VP.t1 94.9962
R899 VP VP.n0 0.336784
R900 VTAIL.n1 VTAIL.t1 56.9126
R901 VTAIL.n3 VTAIL.t0 56.9125
R902 VTAIL.n0 VTAIL.t2 56.9125
R903 VTAIL.n2 VTAIL.t3 56.9125
R904 VTAIL.n1 VTAIL.n0 21.6427
R905 VTAIL.n3 VTAIL.n2 19.1255
R906 VTAIL.n2 VTAIL.n1 1.72895
R907 VTAIL VTAIL.n0 1.15783
R908 VTAIL VTAIL.n3 0.571621
R909 VDD1 VDD1.t0 107.68
R910 VDD1 VDD1.t1 74.2788
R911 VN VN.t1 134.359
R912 VN VN.t0 95.3325
R913 VDD2.n0 VDD2.t1 106.526
R914 VDD2.n0 VDD2.t0 73.5913
R915 VDD2 VDD2.n0 0.688
C0 VTAIL VP 1.38508f
C1 VDD2 VTAIL 3.24552f
C2 VP VN 4.13351f
C3 VDD2 VN 1.28964f
C4 VTAIL VDD1 3.19333f
C5 VDD2 VP 0.336508f
C6 VDD1 VN 0.15224f
C7 VDD1 VP 1.47228f
C8 VDD2 VDD1 0.672578f
C9 VTAIL VN 1.37089f
C10 VDD2 B 3.111776f
C11 VDD1 B 4.97513f
C12 VTAIL B 4.255972f
C13 VN B 7.72838f
C14 VP B 5.755975f
C15 VDD2.t1 B 0.846098f
C16 VDD2.t0 B 0.601286f
C17 VDD2.n0 B 1.65816f
C18 VN.t0 B 0.938246f
C19 VN.t1 B 1.25828f
C20 VDD1.t1 B 0.592783f
C21 VDD1.t0 B 0.852479f
C22 VTAIL.t2 B 0.634869f
C23 VTAIL.n0 B 1.00293f
C24 VTAIL.t1 B 0.634873f
C25 VTAIL.n1 B 1.03433f
C26 VTAIL.t3 B 0.634869f
C27 VTAIL.n2 B 0.895931f
C28 VTAIL.t0 B 0.634869f
C29 VTAIL.n3 B 0.8323f
C30 VP.t0 B 1.26468f
C31 VP.t1 B 0.944185f
C32 VP.n0 B 1.83931f
.ends

