* NGSPICE file created from diff_pair_sample_1554.ext - technology: sky130A

.subckt diff_pair_sample_1554 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=2.0823 ps=12.95 w=12.62 l=0.33
X1 B.t11 B.t9 B.t10 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=0 ps=0 w=12.62 l=0.33
X2 VTAIL.t5 VN.t0 VDD2.t5 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=2.0823 ps=12.95 w=12.62 l=0.33
X3 VDD1.t4 VP.t1 VTAIL.t8 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=4.9218 ps=26.02 w=12.62 l=0.33
X4 B.t8 B.t6 B.t7 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=0 ps=0 w=12.62 l=0.33
X5 VDD2.t4 VN.t1 VTAIL.t0 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=2.0823 ps=12.95 w=12.62 l=0.33
X6 B.t5 B.t3 B.t4 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=0 ps=0 w=12.62 l=0.33
X7 VTAIL.t6 VP.t2 VDD1.t3 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=2.0823 ps=12.95 w=12.62 l=0.33
X8 VDD2.t3 VN.t2 VTAIL.t4 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=4.9218 ps=26.02 w=12.62 l=0.33
X9 VDD2.t2 VN.t3 VTAIL.t3 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=4.9218 ps=26.02 w=12.62 l=0.33
X10 VDD2.t1 VN.t4 VTAIL.t1 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=2.0823 ps=12.95 w=12.62 l=0.33
X11 VDD1.t2 VP.t3 VTAIL.t9 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=4.9218 ps=26.02 w=12.62 l=0.33
X12 VDD1.t1 VP.t4 VTAIL.t10 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=2.0823 ps=12.95 w=12.62 l=0.33
X13 B.t2 B.t0 B.t1 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=4.9218 pd=26.02 as=0 ps=0 w=12.62 l=0.33
X14 VTAIL.t2 VN.t5 VDD2.t0 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=2.0823 ps=12.95 w=12.62 l=0.33
X15 VTAIL.t7 VP.t5 VDD1.t0 w_n1498_n3492# sky130_fd_pr__pfet_01v8 ad=2.0823 pd=12.95 as=2.0823 ps=12.95 w=12.62 l=0.33
R0 VP.n1 VP.t0 1069.75
R1 VP.n8 VP.t1 1039.95
R2 VP.n6 VP.t4 1039.95
R3 VP.n3 VP.t3 1039.95
R4 VP.n7 VP.t5 1016.58
R5 VP.n2 VP.t2 1016.58
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n7 VP.n0 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n7 VP.n6 73.0308
R11 VP.n8 VP.n7 73.0308
R12 VP.n3 VP.n2 73.0308
R13 VP.n4 VP.n1 65.9987
R14 VP.n5 VP.n4 40.2278
R15 VP.n2 VP.n1 29.7615
R16 VP.n5 VP.n0 0.189894
R17 VP.n9 VP.n0 0.189894
R18 VP VP.n9 0.0516364
R19 VTAIL.n286 VTAIL.n285 756.745
R20 VTAIL.n70 VTAIL.n69 756.745
R21 VTAIL.n216 VTAIL.n215 756.745
R22 VTAIL.n144 VTAIL.n143 756.745
R23 VTAIL.n240 VTAIL.n239 585
R24 VTAIL.n245 VTAIL.n244 585
R25 VTAIL.n247 VTAIL.n246 585
R26 VTAIL.n236 VTAIL.n235 585
R27 VTAIL.n253 VTAIL.n252 585
R28 VTAIL.n255 VTAIL.n254 585
R29 VTAIL.n232 VTAIL.n231 585
R30 VTAIL.n261 VTAIL.n260 585
R31 VTAIL.n263 VTAIL.n262 585
R32 VTAIL.n228 VTAIL.n227 585
R33 VTAIL.n269 VTAIL.n268 585
R34 VTAIL.n271 VTAIL.n270 585
R35 VTAIL.n224 VTAIL.n223 585
R36 VTAIL.n277 VTAIL.n276 585
R37 VTAIL.n279 VTAIL.n278 585
R38 VTAIL.n220 VTAIL.n219 585
R39 VTAIL.n285 VTAIL.n284 585
R40 VTAIL.n24 VTAIL.n23 585
R41 VTAIL.n29 VTAIL.n28 585
R42 VTAIL.n31 VTAIL.n30 585
R43 VTAIL.n20 VTAIL.n19 585
R44 VTAIL.n37 VTAIL.n36 585
R45 VTAIL.n39 VTAIL.n38 585
R46 VTAIL.n16 VTAIL.n15 585
R47 VTAIL.n45 VTAIL.n44 585
R48 VTAIL.n47 VTAIL.n46 585
R49 VTAIL.n12 VTAIL.n11 585
R50 VTAIL.n53 VTAIL.n52 585
R51 VTAIL.n55 VTAIL.n54 585
R52 VTAIL.n8 VTAIL.n7 585
R53 VTAIL.n61 VTAIL.n60 585
R54 VTAIL.n63 VTAIL.n62 585
R55 VTAIL.n4 VTAIL.n3 585
R56 VTAIL.n69 VTAIL.n68 585
R57 VTAIL.n215 VTAIL.n214 585
R58 VTAIL.n150 VTAIL.n149 585
R59 VTAIL.n209 VTAIL.n208 585
R60 VTAIL.n207 VTAIL.n206 585
R61 VTAIL.n154 VTAIL.n153 585
R62 VTAIL.n201 VTAIL.n200 585
R63 VTAIL.n199 VTAIL.n198 585
R64 VTAIL.n158 VTAIL.n157 585
R65 VTAIL.n193 VTAIL.n192 585
R66 VTAIL.n191 VTAIL.n190 585
R67 VTAIL.n162 VTAIL.n161 585
R68 VTAIL.n185 VTAIL.n184 585
R69 VTAIL.n183 VTAIL.n182 585
R70 VTAIL.n166 VTAIL.n165 585
R71 VTAIL.n177 VTAIL.n176 585
R72 VTAIL.n175 VTAIL.n174 585
R73 VTAIL.n170 VTAIL.n169 585
R74 VTAIL.n143 VTAIL.n142 585
R75 VTAIL.n78 VTAIL.n77 585
R76 VTAIL.n137 VTAIL.n136 585
R77 VTAIL.n135 VTAIL.n134 585
R78 VTAIL.n82 VTAIL.n81 585
R79 VTAIL.n129 VTAIL.n128 585
R80 VTAIL.n127 VTAIL.n126 585
R81 VTAIL.n86 VTAIL.n85 585
R82 VTAIL.n121 VTAIL.n120 585
R83 VTAIL.n119 VTAIL.n118 585
R84 VTAIL.n90 VTAIL.n89 585
R85 VTAIL.n113 VTAIL.n112 585
R86 VTAIL.n111 VTAIL.n110 585
R87 VTAIL.n94 VTAIL.n93 585
R88 VTAIL.n105 VTAIL.n104 585
R89 VTAIL.n103 VTAIL.n102 585
R90 VTAIL.n98 VTAIL.n97 585
R91 VTAIL.n241 VTAIL.t3 327.466
R92 VTAIL.n25 VTAIL.t8 327.466
R93 VTAIL.n171 VTAIL.t9 327.466
R94 VTAIL.n99 VTAIL.t4 327.466
R95 VTAIL.n245 VTAIL.n239 171.744
R96 VTAIL.n246 VTAIL.n245 171.744
R97 VTAIL.n246 VTAIL.n235 171.744
R98 VTAIL.n253 VTAIL.n235 171.744
R99 VTAIL.n254 VTAIL.n253 171.744
R100 VTAIL.n254 VTAIL.n231 171.744
R101 VTAIL.n261 VTAIL.n231 171.744
R102 VTAIL.n262 VTAIL.n261 171.744
R103 VTAIL.n262 VTAIL.n227 171.744
R104 VTAIL.n269 VTAIL.n227 171.744
R105 VTAIL.n270 VTAIL.n269 171.744
R106 VTAIL.n270 VTAIL.n223 171.744
R107 VTAIL.n277 VTAIL.n223 171.744
R108 VTAIL.n278 VTAIL.n277 171.744
R109 VTAIL.n278 VTAIL.n219 171.744
R110 VTAIL.n285 VTAIL.n219 171.744
R111 VTAIL.n29 VTAIL.n23 171.744
R112 VTAIL.n30 VTAIL.n29 171.744
R113 VTAIL.n30 VTAIL.n19 171.744
R114 VTAIL.n37 VTAIL.n19 171.744
R115 VTAIL.n38 VTAIL.n37 171.744
R116 VTAIL.n38 VTAIL.n15 171.744
R117 VTAIL.n45 VTAIL.n15 171.744
R118 VTAIL.n46 VTAIL.n45 171.744
R119 VTAIL.n46 VTAIL.n11 171.744
R120 VTAIL.n53 VTAIL.n11 171.744
R121 VTAIL.n54 VTAIL.n53 171.744
R122 VTAIL.n54 VTAIL.n7 171.744
R123 VTAIL.n61 VTAIL.n7 171.744
R124 VTAIL.n62 VTAIL.n61 171.744
R125 VTAIL.n62 VTAIL.n3 171.744
R126 VTAIL.n69 VTAIL.n3 171.744
R127 VTAIL.n215 VTAIL.n149 171.744
R128 VTAIL.n208 VTAIL.n149 171.744
R129 VTAIL.n208 VTAIL.n207 171.744
R130 VTAIL.n207 VTAIL.n153 171.744
R131 VTAIL.n200 VTAIL.n153 171.744
R132 VTAIL.n200 VTAIL.n199 171.744
R133 VTAIL.n199 VTAIL.n157 171.744
R134 VTAIL.n192 VTAIL.n157 171.744
R135 VTAIL.n192 VTAIL.n191 171.744
R136 VTAIL.n191 VTAIL.n161 171.744
R137 VTAIL.n184 VTAIL.n161 171.744
R138 VTAIL.n184 VTAIL.n183 171.744
R139 VTAIL.n183 VTAIL.n165 171.744
R140 VTAIL.n176 VTAIL.n165 171.744
R141 VTAIL.n176 VTAIL.n175 171.744
R142 VTAIL.n175 VTAIL.n169 171.744
R143 VTAIL.n143 VTAIL.n77 171.744
R144 VTAIL.n136 VTAIL.n77 171.744
R145 VTAIL.n136 VTAIL.n135 171.744
R146 VTAIL.n135 VTAIL.n81 171.744
R147 VTAIL.n128 VTAIL.n81 171.744
R148 VTAIL.n128 VTAIL.n127 171.744
R149 VTAIL.n127 VTAIL.n85 171.744
R150 VTAIL.n120 VTAIL.n85 171.744
R151 VTAIL.n120 VTAIL.n119 171.744
R152 VTAIL.n119 VTAIL.n89 171.744
R153 VTAIL.n112 VTAIL.n89 171.744
R154 VTAIL.n112 VTAIL.n111 171.744
R155 VTAIL.n111 VTAIL.n93 171.744
R156 VTAIL.n104 VTAIL.n93 171.744
R157 VTAIL.n104 VTAIL.n103 171.744
R158 VTAIL.n103 VTAIL.n97 171.744
R159 VTAIL.t3 VTAIL.n239 85.8723
R160 VTAIL.t8 VTAIL.n23 85.8723
R161 VTAIL.t9 VTAIL.n169 85.8723
R162 VTAIL.t4 VTAIL.n97 85.8723
R163 VTAIL.n147 VTAIL.n146 58.6922
R164 VTAIL.n75 VTAIL.n74 58.6922
R165 VTAIL.n1 VTAIL.n0 58.6912
R166 VTAIL.n73 VTAIL.n72 58.6912
R167 VTAIL.n287 VTAIL.n286 34.5126
R168 VTAIL.n71 VTAIL.n70 34.5126
R169 VTAIL.n217 VTAIL.n216 34.5126
R170 VTAIL.n145 VTAIL.n144 34.5126
R171 VTAIL.n75 VTAIL.n73 24.3841
R172 VTAIL.n287 VTAIL.n217 23.8152
R173 VTAIL.n241 VTAIL.n240 16.3895
R174 VTAIL.n25 VTAIL.n24 16.3895
R175 VTAIL.n171 VTAIL.n170 16.3895
R176 VTAIL.n99 VTAIL.n98 16.3895
R177 VTAIL.n244 VTAIL.n243 12.8005
R178 VTAIL.n284 VTAIL.n218 12.8005
R179 VTAIL.n28 VTAIL.n27 12.8005
R180 VTAIL.n68 VTAIL.n2 12.8005
R181 VTAIL.n214 VTAIL.n148 12.8005
R182 VTAIL.n174 VTAIL.n173 12.8005
R183 VTAIL.n142 VTAIL.n76 12.8005
R184 VTAIL.n102 VTAIL.n101 12.8005
R185 VTAIL.n247 VTAIL.n238 12.0247
R186 VTAIL.n283 VTAIL.n220 12.0247
R187 VTAIL.n31 VTAIL.n22 12.0247
R188 VTAIL.n67 VTAIL.n4 12.0247
R189 VTAIL.n213 VTAIL.n150 12.0247
R190 VTAIL.n177 VTAIL.n168 12.0247
R191 VTAIL.n141 VTAIL.n78 12.0247
R192 VTAIL.n105 VTAIL.n96 12.0247
R193 VTAIL.n248 VTAIL.n236 11.249
R194 VTAIL.n280 VTAIL.n279 11.249
R195 VTAIL.n32 VTAIL.n20 11.249
R196 VTAIL.n64 VTAIL.n63 11.249
R197 VTAIL.n210 VTAIL.n209 11.249
R198 VTAIL.n178 VTAIL.n166 11.249
R199 VTAIL.n138 VTAIL.n137 11.249
R200 VTAIL.n106 VTAIL.n94 11.249
R201 VTAIL.n252 VTAIL.n251 10.4732
R202 VTAIL.n276 VTAIL.n222 10.4732
R203 VTAIL.n36 VTAIL.n35 10.4732
R204 VTAIL.n60 VTAIL.n6 10.4732
R205 VTAIL.n206 VTAIL.n152 10.4732
R206 VTAIL.n182 VTAIL.n181 10.4732
R207 VTAIL.n134 VTAIL.n80 10.4732
R208 VTAIL.n110 VTAIL.n109 10.4732
R209 VTAIL.n255 VTAIL.n234 9.69747
R210 VTAIL.n275 VTAIL.n224 9.69747
R211 VTAIL.n39 VTAIL.n18 9.69747
R212 VTAIL.n59 VTAIL.n8 9.69747
R213 VTAIL.n205 VTAIL.n154 9.69747
R214 VTAIL.n185 VTAIL.n164 9.69747
R215 VTAIL.n133 VTAIL.n82 9.69747
R216 VTAIL.n113 VTAIL.n92 9.69747
R217 VTAIL.n282 VTAIL.n218 9.45567
R218 VTAIL.n66 VTAIL.n2 9.45567
R219 VTAIL.n212 VTAIL.n148 9.45567
R220 VTAIL.n140 VTAIL.n76 9.45567
R221 VTAIL.n265 VTAIL.n264 9.3005
R222 VTAIL.n267 VTAIL.n266 9.3005
R223 VTAIL.n226 VTAIL.n225 9.3005
R224 VTAIL.n273 VTAIL.n272 9.3005
R225 VTAIL.n275 VTAIL.n274 9.3005
R226 VTAIL.n222 VTAIL.n221 9.3005
R227 VTAIL.n281 VTAIL.n280 9.3005
R228 VTAIL.n283 VTAIL.n282 9.3005
R229 VTAIL.n259 VTAIL.n258 9.3005
R230 VTAIL.n257 VTAIL.n256 9.3005
R231 VTAIL.n234 VTAIL.n233 9.3005
R232 VTAIL.n251 VTAIL.n250 9.3005
R233 VTAIL.n249 VTAIL.n248 9.3005
R234 VTAIL.n238 VTAIL.n237 9.3005
R235 VTAIL.n243 VTAIL.n242 9.3005
R236 VTAIL.n230 VTAIL.n229 9.3005
R237 VTAIL.n49 VTAIL.n48 9.3005
R238 VTAIL.n51 VTAIL.n50 9.3005
R239 VTAIL.n10 VTAIL.n9 9.3005
R240 VTAIL.n57 VTAIL.n56 9.3005
R241 VTAIL.n59 VTAIL.n58 9.3005
R242 VTAIL.n6 VTAIL.n5 9.3005
R243 VTAIL.n65 VTAIL.n64 9.3005
R244 VTAIL.n67 VTAIL.n66 9.3005
R245 VTAIL.n43 VTAIL.n42 9.3005
R246 VTAIL.n41 VTAIL.n40 9.3005
R247 VTAIL.n18 VTAIL.n17 9.3005
R248 VTAIL.n35 VTAIL.n34 9.3005
R249 VTAIL.n33 VTAIL.n32 9.3005
R250 VTAIL.n22 VTAIL.n21 9.3005
R251 VTAIL.n27 VTAIL.n26 9.3005
R252 VTAIL.n14 VTAIL.n13 9.3005
R253 VTAIL.n213 VTAIL.n212 9.3005
R254 VTAIL.n211 VTAIL.n210 9.3005
R255 VTAIL.n152 VTAIL.n151 9.3005
R256 VTAIL.n205 VTAIL.n204 9.3005
R257 VTAIL.n203 VTAIL.n202 9.3005
R258 VTAIL.n156 VTAIL.n155 9.3005
R259 VTAIL.n197 VTAIL.n196 9.3005
R260 VTAIL.n195 VTAIL.n194 9.3005
R261 VTAIL.n160 VTAIL.n159 9.3005
R262 VTAIL.n189 VTAIL.n188 9.3005
R263 VTAIL.n187 VTAIL.n186 9.3005
R264 VTAIL.n164 VTAIL.n163 9.3005
R265 VTAIL.n181 VTAIL.n180 9.3005
R266 VTAIL.n179 VTAIL.n178 9.3005
R267 VTAIL.n168 VTAIL.n167 9.3005
R268 VTAIL.n173 VTAIL.n172 9.3005
R269 VTAIL.n125 VTAIL.n124 9.3005
R270 VTAIL.n84 VTAIL.n83 9.3005
R271 VTAIL.n131 VTAIL.n130 9.3005
R272 VTAIL.n133 VTAIL.n132 9.3005
R273 VTAIL.n80 VTAIL.n79 9.3005
R274 VTAIL.n139 VTAIL.n138 9.3005
R275 VTAIL.n141 VTAIL.n140 9.3005
R276 VTAIL.n123 VTAIL.n122 9.3005
R277 VTAIL.n88 VTAIL.n87 9.3005
R278 VTAIL.n117 VTAIL.n116 9.3005
R279 VTAIL.n115 VTAIL.n114 9.3005
R280 VTAIL.n92 VTAIL.n91 9.3005
R281 VTAIL.n109 VTAIL.n108 9.3005
R282 VTAIL.n107 VTAIL.n106 9.3005
R283 VTAIL.n96 VTAIL.n95 9.3005
R284 VTAIL.n101 VTAIL.n100 9.3005
R285 VTAIL.n256 VTAIL.n232 8.92171
R286 VTAIL.n272 VTAIL.n271 8.92171
R287 VTAIL.n40 VTAIL.n16 8.92171
R288 VTAIL.n56 VTAIL.n55 8.92171
R289 VTAIL.n202 VTAIL.n201 8.92171
R290 VTAIL.n186 VTAIL.n162 8.92171
R291 VTAIL.n130 VTAIL.n129 8.92171
R292 VTAIL.n114 VTAIL.n90 8.92171
R293 VTAIL.n260 VTAIL.n259 8.14595
R294 VTAIL.n268 VTAIL.n226 8.14595
R295 VTAIL.n44 VTAIL.n43 8.14595
R296 VTAIL.n52 VTAIL.n10 8.14595
R297 VTAIL.n198 VTAIL.n156 8.14595
R298 VTAIL.n190 VTAIL.n189 8.14595
R299 VTAIL.n126 VTAIL.n84 8.14595
R300 VTAIL.n118 VTAIL.n117 8.14595
R301 VTAIL.n263 VTAIL.n230 7.3702
R302 VTAIL.n267 VTAIL.n228 7.3702
R303 VTAIL.n47 VTAIL.n14 7.3702
R304 VTAIL.n51 VTAIL.n12 7.3702
R305 VTAIL.n197 VTAIL.n158 7.3702
R306 VTAIL.n193 VTAIL.n160 7.3702
R307 VTAIL.n125 VTAIL.n86 7.3702
R308 VTAIL.n121 VTAIL.n88 7.3702
R309 VTAIL.n264 VTAIL.n263 6.59444
R310 VTAIL.n264 VTAIL.n228 6.59444
R311 VTAIL.n48 VTAIL.n47 6.59444
R312 VTAIL.n48 VTAIL.n12 6.59444
R313 VTAIL.n194 VTAIL.n158 6.59444
R314 VTAIL.n194 VTAIL.n193 6.59444
R315 VTAIL.n122 VTAIL.n86 6.59444
R316 VTAIL.n122 VTAIL.n121 6.59444
R317 VTAIL.n260 VTAIL.n230 5.81868
R318 VTAIL.n268 VTAIL.n267 5.81868
R319 VTAIL.n44 VTAIL.n14 5.81868
R320 VTAIL.n52 VTAIL.n51 5.81868
R321 VTAIL.n198 VTAIL.n197 5.81868
R322 VTAIL.n190 VTAIL.n160 5.81868
R323 VTAIL.n126 VTAIL.n125 5.81868
R324 VTAIL.n118 VTAIL.n88 5.81868
R325 VTAIL.n259 VTAIL.n232 5.04292
R326 VTAIL.n271 VTAIL.n226 5.04292
R327 VTAIL.n43 VTAIL.n16 5.04292
R328 VTAIL.n55 VTAIL.n10 5.04292
R329 VTAIL.n201 VTAIL.n156 5.04292
R330 VTAIL.n189 VTAIL.n162 5.04292
R331 VTAIL.n129 VTAIL.n84 5.04292
R332 VTAIL.n117 VTAIL.n90 5.04292
R333 VTAIL.n256 VTAIL.n255 4.26717
R334 VTAIL.n272 VTAIL.n224 4.26717
R335 VTAIL.n40 VTAIL.n39 4.26717
R336 VTAIL.n56 VTAIL.n8 4.26717
R337 VTAIL.n202 VTAIL.n154 4.26717
R338 VTAIL.n186 VTAIL.n185 4.26717
R339 VTAIL.n130 VTAIL.n82 4.26717
R340 VTAIL.n114 VTAIL.n113 4.26717
R341 VTAIL.n242 VTAIL.n241 3.70982
R342 VTAIL.n26 VTAIL.n25 3.70982
R343 VTAIL.n172 VTAIL.n171 3.70982
R344 VTAIL.n100 VTAIL.n99 3.70982
R345 VTAIL.n252 VTAIL.n234 3.49141
R346 VTAIL.n276 VTAIL.n275 3.49141
R347 VTAIL.n36 VTAIL.n18 3.49141
R348 VTAIL.n60 VTAIL.n59 3.49141
R349 VTAIL.n206 VTAIL.n205 3.49141
R350 VTAIL.n182 VTAIL.n164 3.49141
R351 VTAIL.n134 VTAIL.n133 3.49141
R352 VTAIL.n110 VTAIL.n92 3.49141
R353 VTAIL.n251 VTAIL.n236 2.71565
R354 VTAIL.n279 VTAIL.n222 2.71565
R355 VTAIL.n35 VTAIL.n20 2.71565
R356 VTAIL.n63 VTAIL.n6 2.71565
R357 VTAIL.n209 VTAIL.n152 2.71565
R358 VTAIL.n181 VTAIL.n166 2.71565
R359 VTAIL.n137 VTAIL.n80 2.71565
R360 VTAIL.n109 VTAIL.n94 2.71565
R361 VTAIL.n0 VTAIL.t1 2.57617
R362 VTAIL.n0 VTAIL.t5 2.57617
R363 VTAIL.n72 VTAIL.t10 2.57617
R364 VTAIL.n72 VTAIL.t7 2.57617
R365 VTAIL.n146 VTAIL.t11 2.57617
R366 VTAIL.n146 VTAIL.t6 2.57617
R367 VTAIL.n74 VTAIL.t0 2.57617
R368 VTAIL.n74 VTAIL.t2 2.57617
R369 VTAIL.n248 VTAIL.n247 1.93989
R370 VTAIL.n280 VTAIL.n220 1.93989
R371 VTAIL.n32 VTAIL.n31 1.93989
R372 VTAIL.n64 VTAIL.n4 1.93989
R373 VTAIL.n210 VTAIL.n150 1.93989
R374 VTAIL.n178 VTAIL.n177 1.93989
R375 VTAIL.n138 VTAIL.n78 1.93989
R376 VTAIL.n106 VTAIL.n105 1.93989
R377 VTAIL.n244 VTAIL.n238 1.16414
R378 VTAIL.n284 VTAIL.n283 1.16414
R379 VTAIL.n28 VTAIL.n22 1.16414
R380 VTAIL.n68 VTAIL.n67 1.16414
R381 VTAIL.n214 VTAIL.n213 1.16414
R382 VTAIL.n174 VTAIL.n168 1.16414
R383 VTAIL.n142 VTAIL.n141 1.16414
R384 VTAIL.n102 VTAIL.n96 1.16414
R385 VTAIL.n147 VTAIL.n145 0.75481
R386 VTAIL.n71 VTAIL.n1 0.75481
R387 VTAIL.n145 VTAIL.n75 0.569465
R388 VTAIL.n217 VTAIL.n147 0.569465
R389 VTAIL.n73 VTAIL.n71 0.569465
R390 VTAIL.n243 VTAIL.n240 0.388379
R391 VTAIL.n286 VTAIL.n218 0.388379
R392 VTAIL.n27 VTAIL.n24 0.388379
R393 VTAIL.n70 VTAIL.n2 0.388379
R394 VTAIL.n216 VTAIL.n148 0.388379
R395 VTAIL.n173 VTAIL.n170 0.388379
R396 VTAIL.n144 VTAIL.n76 0.388379
R397 VTAIL.n101 VTAIL.n98 0.388379
R398 VTAIL VTAIL.n287 0.369034
R399 VTAIL VTAIL.n1 0.200931
R400 VTAIL.n242 VTAIL.n237 0.155672
R401 VTAIL.n249 VTAIL.n237 0.155672
R402 VTAIL.n250 VTAIL.n249 0.155672
R403 VTAIL.n250 VTAIL.n233 0.155672
R404 VTAIL.n257 VTAIL.n233 0.155672
R405 VTAIL.n258 VTAIL.n257 0.155672
R406 VTAIL.n258 VTAIL.n229 0.155672
R407 VTAIL.n265 VTAIL.n229 0.155672
R408 VTAIL.n266 VTAIL.n265 0.155672
R409 VTAIL.n266 VTAIL.n225 0.155672
R410 VTAIL.n273 VTAIL.n225 0.155672
R411 VTAIL.n274 VTAIL.n273 0.155672
R412 VTAIL.n274 VTAIL.n221 0.155672
R413 VTAIL.n281 VTAIL.n221 0.155672
R414 VTAIL.n282 VTAIL.n281 0.155672
R415 VTAIL.n26 VTAIL.n21 0.155672
R416 VTAIL.n33 VTAIL.n21 0.155672
R417 VTAIL.n34 VTAIL.n33 0.155672
R418 VTAIL.n34 VTAIL.n17 0.155672
R419 VTAIL.n41 VTAIL.n17 0.155672
R420 VTAIL.n42 VTAIL.n41 0.155672
R421 VTAIL.n42 VTAIL.n13 0.155672
R422 VTAIL.n49 VTAIL.n13 0.155672
R423 VTAIL.n50 VTAIL.n49 0.155672
R424 VTAIL.n50 VTAIL.n9 0.155672
R425 VTAIL.n57 VTAIL.n9 0.155672
R426 VTAIL.n58 VTAIL.n57 0.155672
R427 VTAIL.n58 VTAIL.n5 0.155672
R428 VTAIL.n65 VTAIL.n5 0.155672
R429 VTAIL.n66 VTAIL.n65 0.155672
R430 VTAIL.n212 VTAIL.n211 0.155672
R431 VTAIL.n211 VTAIL.n151 0.155672
R432 VTAIL.n204 VTAIL.n151 0.155672
R433 VTAIL.n204 VTAIL.n203 0.155672
R434 VTAIL.n203 VTAIL.n155 0.155672
R435 VTAIL.n196 VTAIL.n155 0.155672
R436 VTAIL.n196 VTAIL.n195 0.155672
R437 VTAIL.n195 VTAIL.n159 0.155672
R438 VTAIL.n188 VTAIL.n159 0.155672
R439 VTAIL.n188 VTAIL.n187 0.155672
R440 VTAIL.n187 VTAIL.n163 0.155672
R441 VTAIL.n180 VTAIL.n163 0.155672
R442 VTAIL.n180 VTAIL.n179 0.155672
R443 VTAIL.n179 VTAIL.n167 0.155672
R444 VTAIL.n172 VTAIL.n167 0.155672
R445 VTAIL.n140 VTAIL.n139 0.155672
R446 VTAIL.n139 VTAIL.n79 0.155672
R447 VTAIL.n132 VTAIL.n79 0.155672
R448 VTAIL.n132 VTAIL.n131 0.155672
R449 VTAIL.n131 VTAIL.n83 0.155672
R450 VTAIL.n124 VTAIL.n83 0.155672
R451 VTAIL.n124 VTAIL.n123 0.155672
R452 VTAIL.n123 VTAIL.n87 0.155672
R453 VTAIL.n116 VTAIL.n87 0.155672
R454 VTAIL.n116 VTAIL.n115 0.155672
R455 VTAIL.n115 VTAIL.n91 0.155672
R456 VTAIL.n108 VTAIL.n91 0.155672
R457 VTAIL.n108 VTAIL.n107 0.155672
R458 VTAIL.n107 VTAIL.n95 0.155672
R459 VTAIL.n100 VTAIL.n95 0.155672
R460 VDD1.n68 VDD1.n67 756.745
R461 VDD1.n137 VDD1.n136 756.745
R462 VDD1.n67 VDD1.n66 585
R463 VDD1.n2 VDD1.n1 585
R464 VDD1.n61 VDD1.n60 585
R465 VDD1.n59 VDD1.n58 585
R466 VDD1.n6 VDD1.n5 585
R467 VDD1.n53 VDD1.n52 585
R468 VDD1.n51 VDD1.n50 585
R469 VDD1.n10 VDD1.n9 585
R470 VDD1.n45 VDD1.n44 585
R471 VDD1.n43 VDD1.n42 585
R472 VDD1.n14 VDD1.n13 585
R473 VDD1.n37 VDD1.n36 585
R474 VDD1.n35 VDD1.n34 585
R475 VDD1.n18 VDD1.n17 585
R476 VDD1.n29 VDD1.n28 585
R477 VDD1.n27 VDD1.n26 585
R478 VDD1.n22 VDD1.n21 585
R479 VDD1.n91 VDD1.n90 585
R480 VDD1.n96 VDD1.n95 585
R481 VDD1.n98 VDD1.n97 585
R482 VDD1.n87 VDD1.n86 585
R483 VDD1.n104 VDD1.n103 585
R484 VDD1.n106 VDD1.n105 585
R485 VDD1.n83 VDD1.n82 585
R486 VDD1.n112 VDD1.n111 585
R487 VDD1.n114 VDD1.n113 585
R488 VDD1.n79 VDD1.n78 585
R489 VDD1.n120 VDD1.n119 585
R490 VDD1.n122 VDD1.n121 585
R491 VDD1.n75 VDD1.n74 585
R492 VDD1.n128 VDD1.n127 585
R493 VDD1.n130 VDD1.n129 585
R494 VDD1.n71 VDD1.n70 585
R495 VDD1.n136 VDD1.n135 585
R496 VDD1.n23 VDD1.t5 327.466
R497 VDD1.n92 VDD1.t1 327.466
R498 VDD1.n67 VDD1.n1 171.744
R499 VDD1.n60 VDD1.n1 171.744
R500 VDD1.n60 VDD1.n59 171.744
R501 VDD1.n59 VDD1.n5 171.744
R502 VDD1.n52 VDD1.n5 171.744
R503 VDD1.n52 VDD1.n51 171.744
R504 VDD1.n51 VDD1.n9 171.744
R505 VDD1.n44 VDD1.n9 171.744
R506 VDD1.n44 VDD1.n43 171.744
R507 VDD1.n43 VDD1.n13 171.744
R508 VDD1.n36 VDD1.n13 171.744
R509 VDD1.n36 VDD1.n35 171.744
R510 VDD1.n35 VDD1.n17 171.744
R511 VDD1.n28 VDD1.n17 171.744
R512 VDD1.n28 VDD1.n27 171.744
R513 VDD1.n27 VDD1.n21 171.744
R514 VDD1.n96 VDD1.n90 171.744
R515 VDD1.n97 VDD1.n96 171.744
R516 VDD1.n97 VDD1.n86 171.744
R517 VDD1.n104 VDD1.n86 171.744
R518 VDD1.n105 VDD1.n104 171.744
R519 VDD1.n105 VDD1.n82 171.744
R520 VDD1.n112 VDD1.n82 171.744
R521 VDD1.n113 VDD1.n112 171.744
R522 VDD1.n113 VDD1.n78 171.744
R523 VDD1.n120 VDD1.n78 171.744
R524 VDD1.n121 VDD1.n120 171.744
R525 VDD1.n121 VDD1.n74 171.744
R526 VDD1.n128 VDD1.n74 171.744
R527 VDD1.n129 VDD1.n128 171.744
R528 VDD1.n129 VDD1.n70 171.744
R529 VDD1.n136 VDD1.n70 171.744
R530 VDD1.t5 VDD1.n21 85.8723
R531 VDD1.t1 VDD1.n90 85.8723
R532 VDD1.n139 VDD1.n138 75.4568
R533 VDD1.n141 VDD1.n140 75.3699
R534 VDD1 VDD1.n68 51.6763
R535 VDD1.n139 VDD1.n137 51.5628
R536 VDD1.n141 VDD1.n139 37.3112
R537 VDD1.n23 VDD1.n22 16.3895
R538 VDD1.n92 VDD1.n91 16.3895
R539 VDD1.n66 VDD1.n0 12.8005
R540 VDD1.n26 VDD1.n25 12.8005
R541 VDD1.n95 VDD1.n94 12.8005
R542 VDD1.n135 VDD1.n69 12.8005
R543 VDD1.n65 VDD1.n2 12.0247
R544 VDD1.n29 VDD1.n20 12.0247
R545 VDD1.n98 VDD1.n89 12.0247
R546 VDD1.n134 VDD1.n71 12.0247
R547 VDD1.n62 VDD1.n61 11.249
R548 VDD1.n30 VDD1.n18 11.249
R549 VDD1.n99 VDD1.n87 11.249
R550 VDD1.n131 VDD1.n130 11.249
R551 VDD1.n58 VDD1.n4 10.4732
R552 VDD1.n34 VDD1.n33 10.4732
R553 VDD1.n103 VDD1.n102 10.4732
R554 VDD1.n127 VDD1.n73 10.4732
R555 VDD1.n57 VDD1.n6 9.69747
R556 VDD1.n37 VDD1.n16 9.69747
R557 VDD1.n106 VDD1.n85 9.69747
R558 VDD1.n126 VDD1.n75 9.69747
R559 VDD1.n64 VDD1.n0 9.45567
R560 VDD1.n133 VDD1.n69 9.45567
R561 VDD1.n49 VDD1.n48 9.3005
R562 VDD1.n8 VDD1.n7 9.3005
R563 VDD1.n55 VDD1.n54 9.3005
R564 VDD1.n57 VDD1.n56 9.3005
R565 VDD1.n4 VDD1.n3 9.3005
R566 VDD1.n63 VDD1.n62 9.3005
R567 VDD1.n65 VDD1.n64 9.3005
R568 VDD1.n47 VDD1.n46 9.3005
R569 VDD1.n12 VDD1.n11 9.3005
R570 VDD1.n41 VDD1.n40 9.3005
R571 VDD1.n39 VDD1.n38 9.3005
R572 VDD1.n16 VDD1.n15 9.3005
R573 VDD1.n33 VDD1.n32 9.3005
R574 VDD1.n31 VDD1.n30 9.3005
R575 VDD1.n20 VDD1.n19 9.3005
R576 VDD1.n25 VDD1.n24 9.3005
R577 VDD1.n116 VDD1.n115 9.3005
R578 VDD1.n118 VDD1.n117 9.3005
R579 VDD1.n77 VDD1.n76 9.3005
R580 VDD1.n124 VDD1.n123 9.3005
R581 VDD1.n126 VDD1.n125 9.3005
R582 VDD1.n73 VDD1.n72 9.3005
R583 VDD1.n132 VDD1.n131 9.3005
R584 VDD1.n134 VDD1.n133 9.3005
R585 VDD1.n110 VDD1.n109 9.3005
R586 VDD1.n108 VDD1.n107 9.3005
R587 VDD1.n85 VDD1.n84 9.3005
R588 VDD1.n102 VDD1.n101 9.3005
R589 VDD1.n100 VDD1.n99 9.3005
R590 VDD1.n89 VDD1.n88 9.3005
R591 VDD1.n94 VDD1.n93 9.3005
R592 VDD1.n81 VDD1.n80 9.3005
R593 VDD1.n54 VDD1.n53 8.92171
R594 VDD1.n38 VDD1.n14 8.92171
R595 VDD1.n107 VDD1.n83 8.92171
R596 VDD1.n123 VDD1.n122 8.92171
R597 VDD1.n50 VDD1.n8 8.14595
R598 VDD1.n42 VDD1.n41 8.14595
R599 VDD1.n111 VDD1.n110 8.14595
R600 VDD1.n119 VDD1.n77 8.14595
R601 VDD1.n49 VDD1.n10 7.3702
R602 VDD1.n45 VDD1.n12 7.3702
R603 VDD1.n114 VDD1.n81 7.3702
R604 VDD1.n118 VDD1.n79 7.3702
R605 VDD1.n46 VDD1.n10 6.59444
R606 VDD1.n46 VDD1.n45 6.59444
R607 VDD1.n115 VDD1.n114 6.59444
R608 VDD1.n115 VDD1.n79 6.59444
R609 VDD1.n50 VDD1.n49 5.81868
R610 VDD1.n42 VDD1.n12 5.81868
R611 VDD1.n111 VDD1.n81 5.81868
R612 VDD1.n119 VDD1.n118 5.81868
R613 VDD1.n53 VDD1.n8 5.04292
R614 VDD1.n41 VDD1.n14 5.04292
R615 VDD1.n110 VDD1.n83 5.04292
R616 VDD1.n122 VDD1.n77 5.04292
R617 VDD1.n54 VDD1.n6 4.26717
R618 VDD1.n38 VDD1.n37 4.26717
R619 VDD1.n107 VDD1.n106 4.26717
R620 VDD1.n123 VDD1.n75 4.26717
R621 VDD1.n24 VDD1.n23 3.70982
R622 VDD1.n93 VDD1.n92 3.70982
R623 VDD1.n58 VDD1.n57 3.49141
R624 VDD1.n34 VDD1.n16 3.49141
R625 VDD1.n103 VDD1.n85 3.49141
R626 VDD1.n127 VDD1.n126 3.49141
R627 VDD1.n61 VDD1.n4 2.71565
R628 VDD1.n33 VDD1.n18 2.71565
R629 VDD1.n102 VDD1.n87 2.71565
R630 VDD1.n130 VDD1.n73 2.71565
R631 VDD1.n140 VDD1.t3 2.57617
R632 VDD1.n140 VDD1.t2 2.57617
R633 VDD1.n138 VDD1.t0 2.57617
R634 VDD1.n138 VDD1.t4 2.57617
R635 VDD1.n62 VDD1.n2 1.93989
R636 VDD1.n30 VDD1.n29 1.93989
R637 VDD1.n99 VDD1.n98 1.93989
R638 VDD1.n131 VDD1.n71 1.93989
R639 VDD1.n66 VDD1.n65 1.16414
R640 VDD1.n26 VDD1.n20 1.16414
R641 VDD1.n95 VDD1.n89 1.16414
R642 VDD1.n135 VDD1.n134 1.16414
R643 VDD1.n68 VDD1.n0 0.388379
R644 VDD1.n25 VDD1.n22 0.388379
R645 VDD1.n94 VDD1.n91 0.388379
R646 VDD1.n137 VDD1.n69 0.388379
R647 VDD1.n64 VDD1.n63 0.155672
R648 VDD1.n63 VDD1.n3 0.155672
R649 VDD1.n56 VDD1.n3 0.155672
R650 VDD1.n56 VDD1.n55 0.155672
R651 VDD1.n55 VDD1.n7 0.155672
R652 VDD1.n48 VDD1.n7 0.155672
R653 VDD1.n48 VDD1.n47 0.155672
R654 VDD1.n47 VDD1.n11 0.155672
R655 VDD1.n40 VDD1.n11 0.155672
R656 VDD1.n40 VDD1.n39 0.155672
R657 VDD1.n39 VDD1.n15 0.155672
R658 VDD1.n32 VDD1.n15 0.155672
R659 VDD1.n32 VDD1.n31 0.155672
R660 VDD1.n31 VDD1.n19 0.155672
R661 VDD1.n24 VDD1.n19 0.155672
R662 VDD1.n93 VDD1.n88 0.155672
R663 VDD1.n100 VDD1.n88 0.155672
R664 VDD1.n101 VDD1.n100 0.155672
R665 VDD1.n101 VDD1.n84 0.155672
R666 VDD1.n108 VDD1.n84 0.155672
R667 VDD1.n109 VDD1.n108 0.155672
R668 VDD1.n109 VDD1.n80 0.155672
R669 VDD1.n116 VDD1.n80 0.155672
R670 VDD1.n117 VDD1.n116 0.155672
R671 VDD1.n117 VDD1.n76 0.155672
R672 VDD1.n124 VDD1.n76 0.155672
R673 VDD1.n125 VDD1.n124 0.155672
R674 VDD1.n125 VDD1.n72 0.155672
R675 VDD1.n132 VDD1.n72 0.155672
R676 VDD1.n133 VDD1.n132 0.155672
R677 VDD1 VDD1.n141 0.0845517
R678 B.n101 B.t6 1134.26
R679 B.n109 B.t9 1134.26
R680 B.n32 B.t0 1134.26
R681 B.n40 B.t3 1134.26
R682 B.n358 B.n357 585
R683 B.n359 B.n62 585
R684 B.n361 B.n360 585
R685 B.n362 B.n61 585
R686 B.n364 B.n363 585
R687 B.n365 B.n60 585
R688 B.n367 B.n366 585
R689 B.n368 B.n59 585
R690 B.n370 B.n369 585
R691 B.n371 B.n58 585
R692 B.n373 B.n372 585
R693 B.n374 B.n57 585
R694 B.n376 B.n375 585
R695 B.n377 B.n56 585
R696 B.n379 B.n378 585
R697 B.n380 B.n55 585
R698 B.n382 B.n381 585
R699 B.n383 B.n54 585
R700 B.n385 B.n384 585
R701 B.n386 B.n53 585
R702 B.n388 B.n387 585
R703 B.n389 B.n52 585
R704 B.n391 B.n390 585
R705 B.n392 B.n51 585
R706 B.n394 B.n393 585
R707 B.n395 B.n50 585
R708 B.n397 B.n396 585
R709 B.n398 B.n49 585
R710 B.n400 B.n399 585
R711 B.n401 B.n48 585
R712 B.n403 B.n402 585
R713 B.n404 B.n47 585
R714 B.n406 B.n405 585
R715 B.n407 B.n46 585
R716 B.n409 B.n408 585
R717 B.n410 B.n45 585
R718 B.n412 B.n411 585
R719 B.n413 B.n44 585
R720 B.n415 B.n414 585
R721 B.n416 B.n43 585
R722 B.n418 B.n417 585
R723 B.n419 B.n39 585
R724 B.n421 B.n420 585
R725 B.n422 B.n38 585
R726 B.n424 B.n423 585
R727 B.n425 B.n37 585
R728 B.n427 B.n426 585
R729 B.n428 B.n36 585
R730 B.n430 B.n429 585
R731 B.n431 B.n35 585
R732 B.n433 B.n432 585
R733 B.n434 B.n34 585
R734 B.n436 B.n435 585
R735 B.n438 B.n31 585
R736 B.n440 B.n439 585
R737 B.n441 B.n30 585
R738 B.n443 B.n442 585
R739 B.n444 B.n29 585
R740 B.n446 B.n445 585
R741 B.n447 B.n28 585
R742 B.n449 B.n448 585
R743 B.n450 B.n27 585
R744 B.n452 B.n451 585
R745 B.n453 B.n26 585
R746 B.n455 B.n454 585
R747 B.n456 B.n25 585
R748 B.n458 B.n457 585
R749 B.n459 B.n24 585
R750 B.n461 B.n460 585
R751 B.n462 B.n23 585
R752 B.n464 B.n463 585
R753 B.n465 B.n22 585
R754 B.n467 B.n466 585
R755 B.n468 B.n21 585
R756 B.n470 B.n469 585
R757 B.n471 B.n20 585
R758 B.n473 B.n472 585
R759 B.n474 B.n19 585
R760 B.n476 B.n475 585
R761 B.n477 B.n18 585
R762 B.n479 B.n478 585
R763 B.n480 B.n17 585
R764 B.n482 B.n481 585
R765 B.n483 B.n16 585
R766 B.n485 B.n484 585
R767 B.n486 B.n15 585
R768 B.n488 B.n487 585
R769 B.n489 B.n14 585
R770 B.n491 B.n490 585
R771 B.n492 B.n13 585
R772 B.n494 B.n493 585
R773 B.n495 B.n12 585
R774 B.n497 B.n496 585
R775 B.n498 B.n11 585
R776 B.n500 B.n499 585
R777 B.n501 B.n10 585
R778 B.n356 B.n63 585
R779 B.n355 B.n354 585
R780 B.n353 B.n64 585
R781 B.n352 B.n351 585
R782 B.n350 B.n65 585
R783 B.n349 B.n348 585
R784 B.n347 B.n66 585
R785 B.n346 B.n345 585
R786 B.n344 B.n67 585
R787 B.n343 B.n342 585
R788 B.n341 B.n68 585
R789 B.n340 B.n339 585
R790 B.n338 B.n69 585
R791 B.n337 B.n336 585
R792 B.n335 B.n70 585
R793 B.n334 B.n333 585
R794 B.n332 B.n71 585
R795 B.n331 B.n330 585
R796 B.n329 B.n72 585
R797 B.n328 B.n327 585
R798 B.n326 B.n73 585
R799 B.n325 B.n324 585
R800 B.n323 B.n74 585
R801 B.n322 B.n321 585
R802 B.n320 B.n75 585
R803 B.n319 B.n318 585
R804 B.n317 B.n76 585
R805 B.n316 B.n315 585
R806 B.n314 B.n77 585
R807 B.n313 B.n312 585
R808 B.n311 B.n78 585
R809 B.n310 B.n309 585
R810 B.n308 B.n79 585
R811 B.n163 B.n162 585
R812 B.n164 B.n131 585
R813 B.n166 B.n165 585
R814 B.n167 B.n130 585
R815 B.n169 B.n168 585
R816 B.n170 B.n129 585
R817 B.n172 B.n171 585
R818 B.n173 B.n128 585
R819 B.n175 B.n174 585
R820 B.n176 B.n127 585
R821 B.n178 B.n177 585
R822 B.n179 B.n126 585
R823 B.n181 B.n180 585
R824 B.n182 B.n125 585
R825 B.n184 B.n183 585
R826 B.n185 B.n124 585
R827 B.n187 B.n186 585
R828 B.n188 B.n123 585
R829 B.n190 B.n189 585
R830 B.n191 B.n122 585
R831 B.n193 B.n192 585
R832 B.n194 B.n121 585
R833 B.n196 B.n195 585
R834 B.n197 B.n120 585
R835 B.n199 B.n198 585
R836 B.n200 B.n119 585
R837 B.n202 B.n201 585
R838 B.n203 B.n118 585
R839 B.n205 B.n204 585
R840 B.n206 B.n117 585
R841 B.n208 B.n207 585
R842 B.n209 B.n116 585
R843 B.n211 B.n210 585
R844 B.n212 B.n115 585
R845 B.n214 B.n213 585
R846 B.n215 B.n114 585
R847 B.n217 B.n216 585
R848 B.n218 B.n113 585
R849 B.n220 B.n219 585
R850 B.n221 B.n112 585
R851 B.n223 B.n222 585
R852 B.n224 B.n111 585
R853 B.n226 B.n225 585
R854 B.n228 B.n108 585
R855 B.n230 B.n229 585
R856 B.n231 B.n107 585
R857 B.n233 B.n232 585
R858 B.n234 B.n106 585
R859 B.n236 B.n235 585
R860 B.n237 B.n105 585
R861 B.n239 B.n238 585
R862 B.n240 B.n104 585
R863 B.n242 B.n241 585
R864 B.n244 B.n243 585
R865 B.n245 B.n100 585
R866 B.n247 B.n246 585
R867 B.n248 B.n99 585
R868 B.n250 B.n249 585
R869 B.n251 B.n98 585
R870 B.n253 B.n252 585
R871 B.n254 B.n97 585
R872 B.n256 B.n255 585
R873 B.n257 B.n96 585
R874 B.n259 B.n258 585
R875 B.n260 B.n95 585
R876 B.n262 B.n261 585
R877 B.n263 B.n94 585
R878 B.n265 B.n264 585
R879 B.n266 B.n93 585
R880 B.n268 B.n267 585
R881 B.n269 B.n92 585
R882 B.n271 B.n270 585
R883 B.n272 B.n91 585
R884 B.n274 B.n273 585
R885 B.n275 B.n90 585
R886 B.n277 B.n276 585
R887 B.n278 B.n89 585
R888 B.n280 B.n279 585
R889 B.n281 B.n88 585
R890 B.n283 B.n282 585
R891 B.n284 B.n87 585
R892 B.n286 B.n285 585
R893 B.n287 B.n86 585
R894 B.n289 B.n288 585
R895 B.n290 B.n85 585
R896 B.n292 B.n291 585
R897 B.n293 B.n84 585
R898 B.n295 B.n294 585
R899 B.n296 B.n83 585
R900 B.n298 B.n297 585
R901 B.n299 B.n82 585
R902 B.n301 B.n300 585
R903 B.n302 B.n81 585
R904 B.n304 B.n303 585
R905 B.n305 B.n80 585
R906 B.n307 B.n306 585
R907 B.n161 B.n132 585
R908 B.n160 B.n159 585
R909 B.n158 B.n133 585
R910 B.n157 B.n156 585
R911 B.n155 B.n134 585
R912 B.n154 B.n153 585
R913 B.n152 B.n135 585
R914 B.n151 B.n150 585
R915 B.n149 B.n136 585
R916 B.n148 B.n147 585
R917 B.n146 B.n137 585
R918 B.n145 B.n144 585
R919 B.n143 B.n138 585
R920 B.n142 B.n141 585
R921 B.n140 B.n139 585
R922 B.n2 B.n0 585
R923 B.n525 B.n1 585
R924 B.n524 B.n523 585
R925 B.n522 B.n3 585
R926 B.n521 B.n520 585
R927 B.n519 B.n4 585
R928 B.n518 B.n517 585
R929 B.n516 B.n5 585
R930 B.n515 B.n514 585
R931 B.n513 B.n6 585
R932 B.n512 B.n511 585
R933 B.n510 B.n7 585
R934 B.n509 B.n508 585
R935 B.n507 B.n8 585
R936 B.n506 B.n505 585
R937 B.n504 B.n9 585
R938 B.n503 B.n502 585
R939 B.n527 B.n526 585
R940 B.n163 B.n132 516.524
R941 B.n502 B.n501 516.524
R942 B.n308 B.n307 516.524
R943 B.n357 B.n356 516.524
R944 B.n101 B.t8 399.413
R945 B.n40 B.t4 399.413
R946 B.n109 B.t11 399.413
R947 B.n32 B.t1 399.413
R948 B.n102 B.t7 386.613
R949 B.n41 B.t5 386.613
R950 B.n110 B.t10 386.613
R951 B.n33 B.t2 386.613
R952 B.n159 B.n132 163.367
R953 B.n159 B.n158 163.367
R954 B.n158 B.n157 163.367
R955 B.n157 B.n134 163.367
R956 B.n153 B.n134 163.367
R957 B.n153 B.n152 163.367
R958 B.n152 B.n151 163.367
R959 B.n151 B.n136 163.367
R960 B.n147 B.n136 163.367
R961 B.n147 B.n146 163.367
R962 B.n146 B.n145 163.367
R963 B.n145 B.n138 163.367
R964 B.n141 B.n138 163.367
R965 B.n141 B.n140 163.367
R966 B.n140 B.n2 163.367
R967 B.n526 B.n2 163.367
R968 B.n526 B.n525 163.367
R969 B.n525 B.n524 163.367
R970 B.n524 B.n3 163.367
R971 B.n520 B.n3 163.367
R972 B.n520 B.n519 163.367
R973 B.n519 B.n518 163.367
R974 B.n518 B.n5 163.367
R975 B.n514 B.n5 163.367
R976 B.n514 B.n513 163.367
R977 B.n513 B.n512 163.367
R978 B.n512 B.n7 163.367
R979 B.n508 B.n7 163.367
R980 B.n508 B.n507 163.367
R981 B.n507 B.n506 163.367
R982 B.n506 B.n9 163.367
R983 B.n502 B.n9 163.367
R984 B.n164 B.n163 163.367
R985 B.n165 B.n164 163.367
R986 B.n165 B.n130 163.367
R987 B.n169 B.n130 163.367
R988 B.n170 B.n169 163.367
R989 B.n171 B.n170 163.367
R990 B.n171 B.n128 163.367
R991 B.n175 B.n128 163.367
R992 B.n176 B.n175 163.367
R993 B.n177 B.n176 163.367
R994 B.n177 B.n126 163.367
R995 B.n181 B.n126 163.367
R996 B.n182 B.n181 163.367
R997 B.n183 B.n182 163.367
R998 B.n183 B.n124 163.367
R999 B.n187 B.n124 163.367
R1000 B.n188 B.n187 163.367
R1001 B.n189 B.n188 163.367
R1002 B.n189 B.n122 163.367
R1003 B.n193 B.n122 163.367
R1004 B.n194 B.n193 163.367
R1005 B.n195 B.n194 163.367
R1006 B.n195 B.n120 163.367
R1007 B.n199 B.n120 163.367
R1008 B.n200 B.n199 163.367
R1009 B.n201 B.n200 163.367
R1010 B.n201 B.n118 163.367
R1011 B.n205 B.n118 163.367
R1012 B.n206 B.n205 163.367
R1013 B.n207 B.n206 163.367
R1014 B.n207 B.n116 163.367
R1015 B.n211 B.n116 163.367
R1016 B.n212 B.n211 163.367
R1017 B.n213 B.n212 163.367
R1018 B.n213 B.n114 163.367
R1019 B.n217 B.n114 163.367
R1020 B.n218 B.n217 163.367
R1021 B.n219 B.n218 163.367
R1022 B.n219 B.n112 163.367
R1023 B.n223 B.n112 163.367
R1024 B.n224 B.n223 163.367
R1025 B.n225 B.n224 163.367
R1026 B.n225 B.n108 163.367
R1027 B.n230 B.n108 163.367
R1028 B.n231 B.n230 163.367
R1029 B.n232 B.n231 163.367
R1030 B.n232 B.n106 163.367
R1031 B.n236 B.n106 163.367
R1032 B.n237 B.n236 163.367
R1033 B.n238 B.n237 163.367
R1034 B.n238 B.n104 163.367
R1035 B.n242 B.n104 163.367
R1036 B.n243 B.n242 163.367
R1037 B.n243 B.n100 163.367
R1038 B.n247 B.n100 163.367
R1039 B.n248 B.n247 163.367
R1040 B.n249 B.n248 163.367
R1041 B.n249 B.n98 163.367
R1042 B.n253 B.n98 163.367
R1043 B.n254 B.n253 163.367
R1044 B.n255 B.n254 163.367
R1045 B.n255 B.n96 163.367
R1046 B.n259 B.n96 163.367
R1047 B.n260 B.n259 163.367
R1048 B.n261 B.n260 163.367
R1049 B.n261 B.n94 163.367
R1050 B.n265 B.n94 163.367
R1051 B.n266 B.n265 163.367
R1052 B.n267 B.n266 163.367
R1053 B.n267 B.n92 163.367
R1054 B.n271 B.n92 163.367
R1055 B.n272 B.n271 163.367
R1056 B.n273 B.n272 163.367
R1057 B.n273 B.n90 163.367
R1058 B.n277 B.n90 163.367
R1059 B.n278 B.n277 163.367
R1060 B.n279 B.n278 163.367
R1061 B.n279 B.n88 163.367
R1062 B.n283 B.n88 163.367
R1063 B.n284 B.n283 163.367
R1064 B.n285 B.n284 163.367
R1065 B.n285 B.n86 163.367
R1066 B.n289 B.n86 163.367
R1067 B.n290 B.n289 163.367
R1068 B.n291 B.n290 163.367
R1069 B.n291 B.n84 163.367
R1070 B.n295 B.n84 163.367
R1071 B.n296 B.n295 163.367
R1072 B.n297 B.n296 163.367
R1073 B.n297 B.n82 163.367
R1074 B.n301 B.n82 163.367
R1075 B.n302 B.n301 163.367
R1076 B.n303 B.n302 163.367
R1077 B.n303 B.n80 163.367
R1078 B.n307 B.n80 163.367
R1079 B.n309 B.n308 163.367
R1080 B.n309 B.n78 163.367
R1081 B.n313 B.n78 163.367
R1082 B.n314 B.n313 163.367
R1083 B.n315 B.n314 163.367
R1084 B.n315 B.n76 163.367
R1085 B.n319 B.n76 163.367
R1086 B.n320 B.n319 163.367
R1087 B.n321 B.n320 163.367
R1088 B.n321 B.n74 163.367
R1089 B.n325 B.n74 163.367
R1090 B.n326 B.n325 163.367
R1091 B.n327 B.n326 163.367
R1092 B.n327 B.n72 163.367
R1093 B.n331 B.n72 163.367
R1094 B.n332 B.n331 163.367
R1095 B.n333 B.n332 163.367
R1096 B.n333 B.n70 163.367
R1097 B.n337 B.n70 163.367
R1098 B.n338 B.n337 163.367
R1099 B.n339 B.n338 163.367
R1100 B.n339 B.n68 163.367
R1101 B.n343 B.n68 163.367
R1102 B.n344 B.n343 163.367
R1103 B.n345 B.n344 163.367
R1104 B.n345 B.n66 163.367
R1105 B.n349 B.n66 163.367
R1106 B.n350 B.n349 163.367
R1107 B.n351 B.n350 163.367
R1108 B.n351 B.n64 163.367
R1109 B.n355 B.n64 163.367
R1110 B.n356 B.n355 163.367
R1111 B.n501 B.n500 163.367
R1112 B.n500 B.n11 163.367
R1113 B.n496 B.n11 163.367
R1114 B.n496 B.n495 163.367
R1115 B.n495 B.n494 163.367
R1116 B.n494 B.n13 163.367
R1117 B.n490 B.n13 163.367
R1118 B.n490 B.n489 163.367
R1119 B.n489 B.n488 163.367
R1120 B.n488 B.n15 163.367
R1121 B.n484 B.n15 163.367
R1122 B.n484 B.n483 163.367
R1123 B.n483 B.n482 163.367
R1124 B.n482 B.n17 163.367
R1125 B.n478 B.n17 163.367
R1126 B.n478 B.n477 163.367
R1127 B.n477 B.n476 163.367
R1128 B.n476 B.n19 163.367
R1129 B.n472 B.n19 163.367
R1130 B.n472 B.n471 163.367
R1131 B.n471 B.n470 163.367
R1132 B.n470 B.n21 163.367
R1133 B.n466 B.n21 163.367
R1134 B.n466 B.n465 163.367
R1135 B.n465 B.n464 163.367
R1136 B.n464 B.n23 163.367
R1137 B.n460 B.n23 163.367
R1138 B.n460 B.n459 163.367
R1139 B.n459 B.n458 163.367
R1140 B.n458 B.n25 163.367
R1141 B.n454 B.n25 163.367
R1142 B.n454 B.n453 163.367
R1143 B.n453 B.n452 163.367
R1144 B.n452 B.n27 163.367
R1145 B.n448 B.n27 163.367
R1146 B.n448 B.n447 163.367
R1147 B.n447 B.n446 163.367
R1148 B.n446 B.n29 163.367
R1149 B.n442 B.n29 163.367
R1150 B.n442 B.n441 163.367
R1151 B.n441 B.n440 163.367
R1152 B.n440 B.n31 163.367
R1153 B.n435 B.n31 163.367
R1154 B.n435 B.n434 163.367
R1155 B.n434 B.n433 163.367
R1156 B.n433 B.n35 163.367
R1157 B.n429 B.n35 163.367
R1158 B.n429 B.n428 163.367
R1159 B.n428 B.n427 163.367
R1160 B.n427 B.n37 163.367
R1161 B.n423 B.n37 163.367
R1162 B.n423 B.n422 163.367
R1163 B.n422 B.n421 163.367
R1164 B.n421 B.n39 163.367
R1165 B.n417 B.n39 163.367
R1166 B.n417 B.n416 163.367
R1167 B.n416 B.n415 163.367
R1168 B.n415 B.n44 163.367
R1169 B.n411 B.n44 163.367
R1170 B.n411 B.n410 163.367
R1171 B.n410 B.n409 163.367
R1172 B.n409 B.n46 163.367
R1173 B.n405 B.n46 163.367
R1174 B.n405 B.n404 163.367
R1175 B.n404 B.n403 163.367
R1176 B.n403 B.n48 163.367
R1177 B.n399 B.n48 163.367
R1178 B.n399 B.n398 163.367
R1179 B.n398 B.n397 163.367
R1180 B.n397 B.n50 163.367
R1181 B.n393 B.n50 163.367
R1182 B.n393 B.n392 163.367
R1183 B.n392 B.n391 163.367
R1184 B.n391 B.n52 163.367
R1185 B.n387 B.n52 163.367
R1186 B.n387 B.n386 163.367
R1187 B.n386 B.n385 163.367
R1188 B.n385 B.n54 163.367
R1189 B.n381 B.n54 163.367
R1190 B.n381 B.n380 163.367
R1191 B.n380 B.n379 163.367
R1192 B.n379 B.n56 163.367
R1193 B.n375 B.n56 163.367
R1194 B.n375 B.n374 163.367
R1195 B.n374 B.n373 163.367
R1196 B.n373 B.n58 163.367
R1197 B.n369 B.n58 163.367
R1198 B.n369 B.n368 163.367
R1199 B.n368 B.n367 163.367
R1200 B.n367 B.n60 163.367
R1201 B.n363 B.n60 163.367
R1202 B.n363 B.n362 163.367
R1203 B.n362 B.n361 163.367
R1204 B.n361 B.n62 163.367
R1205 B.n357 B.n62 163.367
R1206 B.n103 B.n102 59.5399
R1207 B.n227 B.n110 59.5399
R1208 B.n437 B.n33 59.5399
R1209 B.n42 B.n41 59.5399
R1210 B.n503 B.n10 33.5615
R1211 B.n358 B.n63 33.5615
R1212 B.n306 B.n79 33.5615
R1213 B.n162 B.n161 33.5615
R1214 B B.n527 18.0485
R1215 B.n102 B.n101 12.8005
R1216 B.n110 B.n109 12.8005
R1217 B.n33 B.n32 12.8005
R1218 B.n41 B.n40 12.8005
R1219 B.n499 B.n10 10.6151
R1220 B.n499 B.n498 10.6151
R1221 B.n498 B.n497 10.6151
R1222 B.n497 B.n12 10.6151
R1223 B.n493 B.n12 10.6151
R1224 B.n493 B.n492 10.6151
R1225 B.n492 B.n491 10.6151
R1226 B.n491 B.n14 10.6151
R1227 B.n487 B.n14 10.6151
R1228 B.n487 B.n486 10.6151
R1229 B.n486 B.n485 10.6151
R1230 B.n485 B.n16 10.6151
R1231 B.n481 B.n16 10.6151
R1232 B.n481 B.n480 10.6151
R1233 B.n480 B.n479 10.6151
R1234 B.n479 B.n18 10.6151
R1235 B.n475 B.n18 10.6151
R1236 B.n475 B.n474 10.6151
R1237 B.n474 B.n473 10.6151
R1238 B.n473 B.n20 10.6151
R1239 B.n469 B.n20 10.6151
R1240 B.n469 B.n468 10.6151
R1241 B.n468 B.n467 10.6151
R1242 B.n467 B.n22 10.6151
R1243 B.n463 B.n22 10.6151
R1244 B.n463 B.n462 10.6151
R1245 B.n462 B.n461 10.6151
R1246 B.n461 B.n24 10.6151
R1247 B.n457 B.n24 10.6151
R1248 B.n457 B.n456 10.6151
R1249 B.n456 B.n455 10.6151
R1250 B.n455 B.n26 10.6151
R1251 B.n451 B.n26 10.6151
R1252 B.n451 B.n450 10.6151
R1253 B.n450 B.n449 10.6151
R1254 B.n449 B.n28 10.6151
R1255 B.n445 B.n28 10.6151
R1256 B.n445 B.n444 10.6151
R1257 B.n444 B.n443 10.6151
R1258 B.n443 B.n30 10.6151
R1259 B.n439 B.n30 10.6151
R1260 B.n439 B.n438 10.6151
R1261 B.n436 B.n34 10.6151
R1262 B.n432 B.n34 10.6151
R1263 B.n432 B.n431 10.6151
R1264 B.n431 B.n430 10.6151
R1265 B.n430 B.n36 10.6151
R1266 B.n426 B.n36 10.6151
R1267 B.n426 B.n425 10.6151
R1268 B.n425 B.n424 10.6151
R1269 B.n424 B.n38 10.6151
R1270 B.n420 B.n419 10.6151
R1271 B.n419 B.n418 10.6151
R1272 B.n418 B.n43 10.6151
R1273 B.n414 B.n43 10.6151
R1274 B.n414 B.n413 10.6151
R1275 B.n413 B.n412 10.6151
R1276 B.n412 B.n45 10.6151
R1277 B.n408 B.n45 10.6151
R1278 B.n408 B.n407 10.6151
R1279 B.n407 B.n406 10.6151
R1280 B.n406 B.n47 10.6151
R1281 B.n402 B.n47 10.6151
R1282 B.n402 B.n401 10.6151
R1283 B.n401 B.n400 10.6151
R1284 B.n400 B.n49 10.6151
R1285 B.n396 B.n49 10.6151
R1286 B.n396 B.n395 10.6151
R1287 B.n395 B.n394 10.6151
R1288 B.n394 B.n51 10.6151
R1289 B.n390 B.n51 10.6151
R1290 B.n390 B.n389 10.6151
R1291 B.n389 B.n388 10.6151
R1292 B.n388 B.n53 10.6151
R1293 B.n384 B.n53 10.6151
R1294 B.n384 B.n383 10.6151
R1295 B.n383 B.n382 10.6151
R1296 B.n382 B.n55 10.6151
R1297 B.n378 B.n55 10.6151
R1298 B.n378 B.n377 10.6151
R1299 B.n377 B.n376 10.6151
R1300 B.n376 B.n57 10.6151
R1301 B.n372 B.n57 10.6151
R1302 B.n372 B.n371 10.6151
R1303 B.n371 B.n370 10.6151
R1304 B.n370 B.n59 10.6151
R1305 B.n366 B.n59 10.6151
R1306 B.n366 B.n365 10.6151
R1307 B.n365 B.n364 10.6151
R1308 B.n364 B.n61 10.6151
R1309 B.n360 B.n61 10.6151
R1310 B.n360 B.n359 10.6151
R1311 B.n359 B.n358 10.6151
R1312 B.n310 B.n79 10.6151
R1313 B.n311 B.n310 10.6151
R1314 B.n312 B.n311 10.6151
R1315 B.n312 B.n77 10.6151
R1316 B.n316 B.n77 10.6151
R1317 B.n317 B.n316 10.6151
R1318 B.n318 B.n317 10.6151
R1319 B.n318 B.n75 10.6151
R1320 B.n322 B.n75 10.6151
R1321 B.n323 B.n322 10.6151
R1322 B.n324 B.n323 10.6151
R1323 B.n324 B.n73 10.6151
R1324 B.n328 B.n73 10.6151
R1325 B.n329 B.n328 10.6151
R1326 B.n330 B.n329 10.6151
R1327 B.n330 B.n71 10.6151
R1328 B.n334 B.n71 10.6151
R1329 B.n335 B.n334 10.6151
R1330 B.n336 B.n335 10.6151
R1331 B.n336 B.n69 10.6151
R1332 B.n340 B.n69 10.6151
R1333 B.n341 B.n340 10.6151
R1334 B.n342 B.n341 10.6151
R1335 B.n342 B.n67 10.6151
R1336 B.n346 B.n67 10.6151
R1337 B.n347 B.n346 10.6151
R1338 B.n348 B.n347 10.6151
R1339 B.n348 B.n65 10.6151
R1340 B.n352 B.n65 10.6151
R1341 B.n353 B.n352 10.6151
R1342 B.n354 B.n353 10.6151
R1343 B.n354 B.n63 10.6151
R1344 B.n162 B.n131 10.6151
R1345 B.n166 B.n131 10.6151
R1346 B.n167 B.n166 10.6151
R1347 B.n168 B.n167 10.6151
R1348 B.n168 B.n129 10.6151
R1349 B.n172 B.n129 10.6151
R1350 B.n173 B.n172 10.6151
R1351 B.n174 B.n173 10.6151
R1352 B.n174 B.n127 10.6151
R1353 B.n178 B.n127 10.6151
R1354 B.n179 B.n178 10.6151
R1355 B.n180 B.n179 10.6151
R1356 B.n180 B.n125 10.6151
R1357 B.n184 B.n125 10.6151
R1358 B.n185 B.n184 10.6151
R1359 B.n186 B.n185 10.6151
R1360 B.n186 B.n123 10.6151
R1361 B.n190 B.n123 10.6151
R1362 B.n191 B.n190 10.6151
R1363 B.n192 B.n191 10.6151
R1364 B.n192 B.n121 10.6151
R1365 B.n196 B.n121 10.6151
R1366 B.n197 B.n196 10.6151
R1367 B.n198 B.n197 10.6151
R1368 B.n198 B.n119 10.6151
R1369 B.n202 B.n119 10.6151
R1370 B.n203 B.n202 10.6151
R1371 B.n204 B.n203 10.6151
R1372 B.n204 B.n117 10.6151
R1373 B.n208 B.n117 10.6151
R1374 B.n209 B.n208 10.6151
R1375 B.n210 B.n209 10.6151
R1376 B.n210 B.n115 10.6151
R1377 B.n214 B.n115 10.6151
R1378 B.n215 B.n214 10.6151
R1379 B.n216 B.n215 10.6151
R1380 B.n216 B.n113 10.6151
R1381 B.n220 B.n113 10.6151
R1382 B.n221 B.n220 10.6151
R1383 B.n222 B.n221 10.6151
R1384 B.n222 B.n111 10.6151
R1385 B.n226 B.n111 10.6151
R1386 B.n229 B.n228 10.6151
R1387 B.n229 B.n107 10.6151
R1388 B.n233 B.n107 10.6151
R1389 B.n234 B.n233 10.6151
R1390 B.n235 B.n234 10.6151
R1391 B.n235 B.n105 10.6151
R1392 B.n239 B.n105 10.6151
R1393 B.n240 B.n239 10.6151
R1394 B.n241 B.n240 10.6151
R1395 B.n245 B.n244 10.6151
R1396 B.n246 B.n245 10.6151
R1397 B.n246 B.n99 10.6151
R1398 B.n250 B.n99 10.6151
R1399 B.n251 B.n250 10.6151
R1400 B.n252 B.n251 10.6151
R1401 B.n252 B.n97 10.6151
R1402 B.n256 B.n97 10.6151
R1403 B.n257 B.n256 10.6151
R1404 B.n258 B.n257 10.6151
R1405 B.n258 B.n95 10.6151
R1406 B.n262 B.n95 10.6151
R1407 B.n263 B.n262 10.6151
R1408 B.n264 B.n263 10.6151
R1409 B.n264 B.n93 10.6151
R1410 B.n268 B.n93 10.6151
R1411 B.n269 B.n268 10.6151
R1412 B.n270 B.n269 10.6151
R1413 B.n270 B.n91 10.6151
R1414 B.n274 B.n91 10.6151
R1415 B.n275 B.n274 10.6151
R1416 B.n276 B.n275 10.6151
R1417 B.n276 B.n89 10.6151
R1418 B.n280 B.n89 10.6151
R1419 B.n281 B.n280 10.6151
R1420 B.n282 B.n281 10.6151
R1421 B.n282 B.n87 10.6151
R1422 B.n286 B.n87 10.6151
R1423 B.n287 B.n286 10.6151
R1424 B.n288 B.n287 10.6151
R1425 B.n288 B.n85 10.6151
R1426 B.n292 B.n85 10.6151
R1427 B.n293 B.n292 10.6151
R1428 B.n294 B.n293 10.6151
R1429 B.n294 B.n83 10.6151
R1430 B.n298 B.n83 10.6151
R1431 B.n299 B.n298 10.6151
R1432 B.n300 B.n299 10.6151
R1433 B.n300 B.n81 10.6151
R1434 B.n304 B.n81 10.6151
R1435 B.n305 B.n304 10.6151
R1436 B.n306 B.n305 10.6151
R1437 B.n161 B.n160 10.6151
R1438 B.n160 B.n133 10.6151
R1439 B.n156 B.n133 10.6151
R1440 B.n156 B.n155 10.6151
R1441 B.n155 B.n154 10.6151
R1442 B.n154 B.n135 10.6151
R1443 B.n150 B.n135 10.6151
R1444 B.n150 B.n149 10.6151
R1445 B.n149 B.n148 10.6151
R1446 B.n148 B.n137 10.6151
R1447 B.n144 B.n137 10.6151
R1448 B.n144 B.n143 10.6151
R1449 B.n143 B.n142 10.6151
R1450 B.n142 B.n139 10.6151
R1451 B.n139 B.n0 10.6151
R1452 B.n523 B.n1 10.6151
R1453 B.n523 B.n522 10.6151
R1454 B.n522 B.n521 10.6151
R1455 B.n521 B.n4 10.6151
R1456 B.n517 B.n4 10.6151
R1457 B.n517 B.n516 10.6151
R1458 B.n516 B.n515 10.6151
R1459 B.n515 B.n6 10.6151
R1460 B.n511 B.n6 10.6151
R1461 B.n511 B.n510 10.6151
R1462 B.n510 B.n509 10.6151
R1463 B.n509 B.n8 10.6151
R1464 B.n505 B.n8 10.6151
R1465 B.n505 B.n504 10.6151
R1466 B.n504 B.n503 10.6151
R1467 B.n438 B.n437 9.36635
R1468 B.n420 B.n42 9.36635
R1469 B.n227 B.n226 9.36635
R1470 B.n244 B.n103 9.36635
R1471 B.n527 B.n0 2.81026
R1472 B.n527 B.n1 2.81026
R1473 B.n437 B.n436 1.24928
R1474 B.n42 B.n38 1.24928
R1475 B.n228 B.n227 1.24928
R1476 B.n241 B.n103 1.24928
R1477 VN.n0 VN.t4 1069.75
R1478 VN.n4 VN.t2 1069.75
R1479 VN.n2 VN.t3 1039.95
R1480 VN.n6 VN.t1 1039.95
R1481 VN.n1 VN.t0 1016.58
R1482 VN.n5 VN.t5 1016.58
R1483 VN.n3 VN.n2 161.3
R1484 VN.n7 VN.n6 161.3
R1485 VN.n2 VN.n1 73.0308
R1486 VN.n6 VN.n5 73.0308
R1487 VN.n7 VN.n4 65.9987
R1488 VN.n3 VN.n0 65.9987
R1489 VN VN.n7 40.6085
R1490 VN.n5 VN.n4 29.7615
R1491 VN.n1 VN.n0 29.7615
R1492 VN VN.n3 0.0516364
R1493 VDD2.n139 VDD2.n138 756.745
R1494 VDD2.n68 VDD2.n67 756.745
R1495 VDD2.n138 VDD2.n137 585
R1496 VDD2.n73 VDD2.n72 585
R1497 VDD2.n132 VDD2.n131 585
R1498 VDD2.n130 VDD2.n129 585
R1499 VDD2.n77 VDD2.n76 585
R1500 VDD2.n124 VDD2.n123 585
R1501 VDD2.n122 VDD2.n121 585
R1502 VDD2.n81 VDD2.n80 585
R1503 VDD2.n116 VDD2.n115 585
R1504 VDD2.n114 VDD2.n113 585
R1505 VDD2.n85 VDD2.n84 585
R1506 VDD2.n108 VDD2.n107 585
R1507 VDD2.n106 VDD2.n105 585
R1508 VDD2.n89 VDD2.n88 585
R1509 VDD2.n100 VDD2.n99 585
R1510 VDD2.n98 VDD2.n97 585
R1511 VDD2.n93 VDD2.n92 585
R1512 VDD2.n22 VDD2.n21 585
R1513 VDD2.n27 VDD2.n26 585
R1514 VDD2.n29 VDD2.n28 585
R1515 VDD2.n18 VDD2.n17 585
R1516 VDD2.n35 VDD2.n34 585
R1517 VDD2.n37 VDD2.n36 585
R1518 VDD2.n14 VDD2.n13 585
R1519 VDD2.n43 VDD2.n42 585
R1520 VDD2.n45 VDD2.n44 585
R1521 VDD2.n10 VDD2.n9 585
R1522 VDD2.n51 VDD2.n50 585
R1523 VDD2.n53 VDD2.n52 585
R1524 VDD2.n6 VDD2.n5 585
R1525 VDD2.n59 VDD2.n58 585
R1526 VDD2.n61 VDD2.n60 585
R1527 VDD2.n2 VDD2.n1 585
R1528 VDD2.n67 VDD2.n66 585
R1529 VDD2.n94 VDD2.t4 327.466
R1530 VDD2.n23 VDD2.t1 327.466
R1531 VDD2.n138 VDD2.n72 171.744
R1532 VDD2.n131 VDD2.n72 171.744
R1533 VDD2.n131 VDD2.n130 171.744
R1534 VDD2.n130 VDD2.n76 171.744
R1535 VDD2.n123 VDD2.n76 171.744
R1536 VDD2.n123 VDD2.n122 171.744
R1537 VDD2.n122 VDD2.n80 171.744
R1538 VDD2.n115 VDD2.n80 171.744
R1539 VDD2.n115 VDD2.n114 171.744
R1540 VDD2.n114 VDD2.n84 171.744
R1541 VDD2.n107 VDD2.n84 171.744
R1542 VDD2.n107 VDD2.n106 171.744
R1543 VDD2.n106 VDD2.n88 171.744
R1544 VDD2.n99 VDD2.n88 171.744
R1545 VDD2.n99 VDD2.n98 171.744
R1546 VDD2.n98 VDD2.n92 171.744
R1547 VDD2.n27 VDD2.n21 171.744
R1548 VDD2.n28 VDD2.n27 171.744
R1549 VDD2.n28 VDD2.n17 171.744
R1550 VDD2.n35 VDD2.n17 171.744
R1551 VDD2.n36 VDD2.n35 171.744
R1552 VDD2.n36 VDD2.n13 171.744
R1553 VDD2.n43 VDD2.n13 171.744
R1554 VDD2.n44 VDD2.n43 171.744
R1555 VDD2.n44 VDD2.n9 171.744
R1556 VDD2.n51 VDD2.n9 171.744
R1557 VDD2.n52 VDD2.n51 171.744
R1558 VDD2.n52 VDD2.n5 171.744
R1559 VDD2.n59 VDD2.n5 171.744
R1560 VDD2.n60 VDD2.n59 171.744
R1561 VDD2.n60 VDD2.n1 171.744
R1562 VDD2.n67 VDD2.n1 171.744
R1563 VDD2.t4 VDD2.n92 85.8723
R1564 VDD2.t1 VDD2.n21 85.8723
R1565 VDD2.n70 VDD2.n69 75.4568
R1566 VDD2 VDD2.n141 75.4539
R1567 VDD2.n70 VDD2.n68 51.5628
R1568 VDD2.n140 VDD2.n139 51.1914
R1569 VDD2.n140 VDD2.n70 36.4437
R1570 VDD2.n94 VDD2.n93 16.3895
R1571 VDD2.n23 VDD2.n22 16.3895
R1572 VDD2.n137 VDD2.n71 12.8005
R1573 VDD2.n97 VDD2.n96 12.8005
R1574 VDD2.n26 VDD2.n25 12.8005
R1575 VDD2.n66 VDD2.n0 12.8005
R1576 VDD2.n136 VDD2.n73 12.0247
R1577 VDD2.n100 VDD2.n91 12.0247
R1578 VDD2.n29 VDD2.n20 12.0247
R1579 VDD2.n65 VDD2.n2 12.0247
R1580 VDD2.n133 VDD2.n132 11.249
R1581 VDD2.n101 VDD2.n89 11.249
R1582 VDD2.n30 VDD2.n18 11.249
R1583 VDD2.n62 VDD2.n61 11.249
R1584 VDD2.n129 VDD2.n75 10.4732
R1585 VDD2.n105 VDD2.n104 10.4732
R1586 VDD2.n34 VDD2.n33 10.4732
R1587 VDD2.n58 VDD2.n4 10.4732
R1588 VDD2.n128 VDD2.n77 9.69747
R1589 VDD2.n108 VDD2.n87 9.69747
R1590 VDD2.n37 VDD2.n16 9.69747
R1591 VDD2.n57 VDD2.n6 9.69747
R1592 VDD2.n135 VDD2.n71 9.45567
R1593 VDD2.n64 VDD2.n0 9.45567
R1594 VDD2.n120 VDD2.n119 9.3005
R1595 VDD2.n79 VDD2.n78 9.3005
R1596 VDD2.n126 VDD2.n125 9.3005
R1597 VDD2.n128 VDD2.n127 9.3005
R1598 VDD2.n75 VDD2.n74 9.3005
R1599 VDD2.n134 VDD2.n133 9.3005
R1600 VDD2.n136 VDD2.n135 9.3005
R1601 VDD2.n118 VDD2.n117 9.3005
R1602 VDD2.n83 VDD2.n82 9.3005
R1603 VDD2.n112 VDD2.n111 9.3005
R1604 VDD2.n110 VDD2.n109 9.3005
R1605 VDD2.n87 VDD2.n86 9.3005
R1606 VDD2.n104 VDD2.n103 9.3005
R1607 VDD2.n102 VDD2.n101 9.3005
R1608 VDD2.n91 VDD2.n90 9.3005
R1609 VDD2.n96 VDD2.n95 9.3005
R1610 VDD2.n47 VDD2.n46 9.3005
R1611 VDD2.n49 VDD2.n48 9.3005
R1612 VDD2.n8 VDD2.n7 9.3005
R1613 VDD2.n55 VDD2.n54 9.3005
R1614 VDD2.n57 VDD2.n56 9.3005
R1615 VDD2.n4 VDD2.n3 9.3005
R1616 VDD2.n63 VDD2.n62 9.3005
R1617 VDD2.n65 VDD2.n64 9.3005
R1618 VDD2.n41 VDD2.n40 9.3005
R1619 VDD2.n39 VDD2.n38 9.3005
R1620 VDD2.n16 VDD2.n15 9.3005
R1621 VDD2.n33 VDD2.n32 9.3005
R1622 VDD2.n31 VDD2.n30 9.3005
R1623 VDD2.n20 VDD2.n19 9.3005
R1624 VDD2.n25 VDD2.n24 9.3005
R1625 VDD2.n12 VDD2.n11 9.3005
R1626 VDD2.n125 VDD2.n124 8.92171
R1627 VDD2.n109 VDD2.n85 8.92171
R1628 VDD2.n38 VDD2.n14 8.92171
R1629 VDD2.n54 VDD2.n53 8.92171
R1630 VDD2.n121 VDD2.n79 8.14595
R1631 VDD2.n113 VDD2.n112 8.14595
R1632 VDD2.n42 VDD2.n41 8.14595
R1633 VDD2.n50 VDD2.n8 8.14595
R1634 VDD2.n120 VDD2.n81 7.3702
R1635 VDD2.n116 VDD2.n83 7.3702
R1636 VDD2.n45 VDD2.n12 7.3702
R1637 VDD2.n49 VDD2.n10 7.3702
R1638 VDD2.n117 VDD2.n81 6.59444
R1639 VDD2.n117 VDD2.n116 6.59444
R1640 VDD2.n46 VDD2.n45 6.59444
R1641 VDD2.n46 VDD2.n10 6.59444
R1642 VDD2.n121 VDD2.n120 5.81868
R1643 VDD2.n113 VDD2.n83 5.81868
R1644 VDD2.n42 VDD2.n12 5.81868
R1645 VDD2.n50 VDD2.n49 5.81868
R1646 VDD2.n124 VDD2.n79 5.04292
R1647 VDD2.n112 VDD2.n85 5.04292
R1648 VDD2.n41 VDD2.n14 5.04292
R1649 VDD2.n53 VDD2.n8 5.04292
R1650 VDD2.n125 VDD2.n77 4.26717
R1651 VDD2.n109 VDD2.n108 4.26717
R1652 VDD2.n38 VDD2.n37 4.26717
R1653 VDD2.n54 VDD2.n6 4.26717
R1654 VDD2.n95 VDD2.n94 3.70982
R1655 VDD2.n24 VDD2.n23 3.70982
R1656 VDD2.n129 VDD2.n128 3.49141
R1657 VDD2.n105 VDD2.n87 3.49141
R1658 VDD2.n34 VDD2.n16 3.49141
R1659 VDD2.n58 VDD2.n57 3.49141
R1660 VDD2.n132 VDD2.n75 2.71565
R1661 VDD2.n104 VDD2.n89 2.71565
R1662 VDD2.n33 VDD2.n18 2.71565
R1663 VDD2.n61 VDD2.n4 2.71565
R1664 VDD2.n141 VDD2.t0 2.57617
R1665 VDD2.n141 VDD2.t3 2.57617
R1666 VDD2.n69 VDD2.t5 2.57617
R1667 VDD2.n69 VDD2.t2 2.57617
R1668 VDD2.n133 VDD2.n73 1.93989
R1669 VDD2.n101 VDD2.n100 1.93989
R1670 VDD2.n30 VDD2.n29 1.93989
R1671 VDD2.n62 VDD2.n2 1.93989
R1672 VDD2.n137 VDD2.n136 1.16414
R1673 VDD2.n97 VDD2.n91 1.16414
R1674 VDD2.n26 VDD2.n20 1.16414
R1675 VDD2.n66 VDD2.n65 1.16414
R1676 VDD2 VDD2.n140 0.485414
R1677 VDD2.n139 VDD2.n71 0.388379
R1678 VDD2.n96 VDD2.n93 0.388379
R1679 VDD2.n25 VDD2.n22 0.388379
R1680 VDD2.n68 VDD2.n0 0.388379
R1681 VDD2.n135 VDD2.n134 0.155672
R1682 VDD2.n134 VDD2.n74 0.155672
R1683 VDD2.n127 VDD2.n74 0.155672
R1684 VDD2.n127 VDD2.n126 0.155672
R1685 VDD2.n126 VDD2.n78 0.155672
R1686 VDD2.n119 VDD2.n78 0.155672
R1687 VDD2.n119 VDD2.n118 0.155672
R1688 VDD2.n118 VDD2.n82 0.155672
R1689 VDD2.n111 VDD2.n82 0.155672
R1690 VDD2.n111 VDD2.n110 0.155672
R1691 VDD2.n110 VDD2.n86 0.155672
R1692 VDD2.n103 VDD2.n86 0.155672
R1693 VDD2.n103 VDD2.n102 0.155672
R1694 VDD2.n102 VDD2.n90 0.155672
R1695 VDD2.n95 VDD2.n90 0.155672
R1696 VDD2.n24 VDD2.n19 0.155672
R1697 VDD2.n31 VDD2.n19 0.155672
R1698 VDD2.n32 VDD2.n31 0.155672
R1699 VDD2.n32 VDD2.n15 0.155672
R1700 VDD2.n39 VDD2.n15 0.155672
R1701 VDD2.n40 VDD2.n39 0.155672
R1702 VDD2.n40 VDD2.n11 0.155672
R1703 VDD2.n47 VDD2.n11 0.155672
R1704 VDD2.n48 VDD2.n47 0.155672
R1705 VDD2.n48 VDD2.n7 0.155672
R1706 VDD2.n55 VDD2.n7 0.155672
R1707 VDD2.n56 VDD2.n55 0.155672
R1708 VDD2.n56 VDD2.n3 0.155672
R1709 VDD2.n63 VDD2.n3 0.155672
R1710 VDD2.n64 VDD2.n63 0.155672
C0 VP B 0.993795f
C1 VTAIL VP 2.53481f
C2 VN VDD2 2.99764f
C3 B VDD2 1.50637f
C4 VTAIL VDD2 14.048599f
C5 VN B 0.692432f
C6 VN VTAIL 2.52003f
C7 w_n1498_n3492# VP 2.4901f
C8 VTAIL B 2.54734f
C9 w_n1498_n3492# VDD2 1.76534f
C10 VP VDD1 3.11128f
C11 w_n1498_n3492# VN 2.30275f
C12 VDD2 VDD1 0.581314f
C13 w_n1498_n3492# B 6.71925f
C14 w_n1498_n3492# VTAIL 3.09836f
C15 VN VDD1 0.148022f
C16 B VDD1 1.48558f
C17 VTAIL VDD1 14.0191f
C18 VP VDD2 0.266964f
C19 VN VP 4.83648f
C20 w_n1498_n3492# VDD1 1.7524f
C21 VDD2 VSUBS 1.334223f
C22 VDD1 VSUBS 1.057283f
C23 VTAIL VSUBS 0.615846f
C24 VN VSUBS 4.46718f
C25 VP VSUBS 1.209681f
C26 B VSUBS 2.431375f
C27 w_n1498_n3492# VSUBS 64.336105f
C28 VDD2.n0 VSUBS 0.015275f
C29 VDD2.n1 VSUBS 0.034495f
C30 VDD2.n2 VSUBS 0.015453f
C31 VDD2.n3 VSUBS 0.027159f
C32 VDD2.n4 VSUBS 0.014594f
C33 VDD2.n5 VSUBS 0.034495f
C34 VDD2.n6 VSUBS 0.015453f
C35 VDD2.n7 VSUBS 0.027159f
C36 VDD2.n8 VSUBS 0.014594f
C37 VDD2.n9 VSUBS 0.034495f
C38 VDD2.n10 VSUBS 0.015453f
C39 VDD2.n11 VSUBS 0.027159f
C40 VDD2.n12 VSUBS 0.014594f
C41 VDD2.n13 VSUBS 0.034495f
C42 VDD2.n14 VSUBS 0.015453f
C43 VDD2.n15 VSUBS 0.027159f
C44 VDD2.n16 VSUBS 0.014594f
C45 VDD2.n17 VSUBS 0.034495f
C46 VDD2.n18 VSUBS 0.015453f
C47 VDD2.n19 VSUBS 0.027159f
C48 VDD2.n20 VSUBS 0.014594f
C49 VDD2.n21 VSUBS 0.025871f
C50 VDD2.n22 VSUBS 0.021944f
C51 VDD2.t1 VSUBS 0.073689f
C52 VDD2.n23 VSUBS 0.172385f
C53 VDD2.n24 VSUBS 1.44072f
C54 VDD2.n25 VSUBS 0.014594f
C55 VDD2.n26 VSUBS 0.015453f
C56 VDD2.n27 VSUBS 0.034495f
C57 VDD2.n28 VSUBS 0.034495f
C58 VDD2.n29 VSUBS 0.015453f
C59 VDD2.n30 VSUBS 0.014594f
C60 VDD2.n31 VSUBS 0.027159f
C61 VDD2.n32 VSUBS 0.027159f
C62 VDD2.n33 VSUBS 0.014594f
C63 VDD2.n34 VSUBS 0.015453f
C64 VDD2.n35 VSUBS 0.034495f
C65 VDD2.n36 VSUBS 0.034495f
C66 VDD2.n37 VSUBS 0.015453f
C67 VDD2.n38 VSUBS 0.014594f
C68 VDD2.n39 VSUBS 0.027159f
C69 VDD2.n40 VSUBS 0.027159f
C70 VDD2.n41 VSUBS 0.014594f
C71 VDD2.n42 VSUBS 0.015453f
C72 VDD2.n43 VSUBS 0.034495f
C73 VDD2.n44 VSUBS 0.034495f
C74 VDD2.n45 VSUBS 0.015453f
C75 VDD2.n46 VSUBS 0.014594f
C76 VDD2.n47 VSUBS 0.027159f
C77 VDD2.n48 VSUBS 0.027159f
C78 VDD2.n49 VSUBS 0.014594f
C79 VDD2.n50 VSUBS 0.015453f
C80 VDD2.n51 VSUBS 0.034495f
C81 VDD2.n52 VSUBS 0.034495f
C82 VDD2.n53 VSUBS 0.015453f
C83 VDD2.n54 VSUBS 0.014594f
C84 VDD2.n55 VSUBS 0.027159f
C85 VDD2.n56 VSUBS 0.027159f
C86 VDD2.n57 VSUBS 0.014594f
C87 VDD2.n58 VSUBS 0.015453f
C88 VDD2.n59 VSUBS 0.034495f
C89 VDD2.n60 VSUBS 0.034495f
C90 VDD2.n61 VSUBS 0.015453f
C91 VDD2.n62 VSUBS 0.014594f
C92 VDD2.n63 VSUBS 0.027159f
C93 VDD2.n64 VSUBS 0.067971f
C94 VDD2.n65 VSUBS 0.014594f
C95 VDD2.n66 VSUBS 0.015453f
C96 VDD2.n67 VSUBS 0.076064f
C97 VDD2.n68 VSUBS 0.06938f
C98 VDD2.t5 VSUBS 0.27085f
C99 VDD2.t2 VSUBS 0.27085f
C100 VDD2.n69 VSUBS 2.15311f
C101 VDD2.n70 VSUBS 2.14984f
C102 VDD2.n71 VSUBS 0.015275f
C103 VDD2.n72 VSUBS 0.034495f
C104 VDD2.n73 VSUBS 0.015453f
C105 VDD2.n74 VSUBS 0.027159f
C106 VDD2.n75 VSUBS 0.014594f
C107 VDD2.n76 VSUBS 0.034495f
C108 VDD2.n77 VSUBS 0.015453f
C109 VDD2.n78 VSUBS 0.027159f
C110 VDD2.n79 VSUBS 0.014594f
C111 VDD2.n80 VSUBS 0.034495f
C112 VDD2.n81 VSUBS 0.015453f
C113 VDD2.n82 VSUBS 0.027159f
C114 VDD2.n83 VSUBS 0.014594f
C115 VDD2.n84 VSUBS 0.034495f
C116 VDD2.n85 VSUBS 0.015453f
C117 VDD2.n86 VSUBS 0.027159f
C118 VDD2.n87 VSUBS 0.014594f
C119 VDD2.n88 VSUBS 0.034495f
C120 VDD2.n89 VSUBS 0.015453f
C121 VDD2.n90 VSUBS 0.027159f
C122 VDD2.n91 VSUBS 0.014594f
C123 VDD2.n92 VSUBS 0.025871f
C124 VDD2.n93 VSUBS 0.021944f
C125 VDD2.t4 VSUBS 0.073689f
C126 VDD2.n94 VSUBS 0.172385f
C127 VDD2.n95 VSUBS 1.44072f
C128 VDD2.n96 VSUBS 0.014594f
C129 VDD2.n97 VSUBS 0.015453f
C130 VDD2.n98 VSUBS 0.034495f
C131 VDD2.n99 VSUBS 0.034495f
C132 VDD2.n100 VSUBS 0.015453f
C133 VDD2.n101 VSUBS 0.014594f
C134 VDD2.n102 VSUBS 0.027159f
C135 VDD2.n103 VSUBS 0.027159f
C136 VDD2.n104 VSUBS 0.014594f
C137 VDD2.n105 VSUBS 0.015453f
C138 VDD2.n106 VSUBS 0.034495f
C139 VDD2.n107 VSUBS 0.034495f
C140 VDD2.n108 VSUBS 0.015453f
C141 VDD2.n109 VSUBS 0.014594f
C142 VDD2.n110 VSUBS 0.027159f
C143 VDD2.n111 VSUBS 0.027159f
C144 VDD2.n112 VSUBS 0.014594f
C145 VDD2.n113 VSUBS 0.015453f
C146 VDD2.n114 VSUBS 0.034495f
C147 VDD2.n115 VSUBS 0.034495f
C148 VDD2.n116 VSUBS 0.015453f
C149 VDD2.n117 VSUBS 0.014594f
C150 VDD2.n118 VSUBS 0.027159f
C151 VDD2.n119 VSUBS 0.027159f
C152 VDD2.n120 VSUBS 0.014594f
C153 VDD2.n121 VSUBS 0.015453f
C154 VDD2.n122 VSUBS 0.034495f
C155 VDD2.n123 VSUBS 0.034495f
C156 VDD2.n124 VSUBS 0.015453f
C157 VDD2.n125 VSUBS 0.014594f
C158 VDD2.n126 VSUBS 0.027159f
C159 VDD2.n127 VSUBS 0.027159f
C160 VDD2.n128 VSUBS 0.014594f
C161 VDD2.n129 VSUBS 0.015453f
C162 VDD2.n130 VSUBS 0.034495f
C163 VDD2.n131 VSUBS 0.034495f
C164 VDD2.n132 VSUBS 0.015453f
C165 VDD2.n133 VSUBS 0.014594f
C166 VDD2.n134 VSUBS 0.027159f
C167 VDD2.n135 VSUBS 0.067971f
C168 VDD2.n136 VSUBS 0.014594f
C169 VDD2.n137 VSUBS 0.015453f
C170 VDD2.n138 VSUBS 0.076064f
C171 VDD2.n139 VSUBS 0.068738f
C172 VDD2.n140 VSUBS 2.1667f
C173 VDD2.t0 VSUBS 0.27085f
C174 VDD2.t3 VSUBS 0.27085f
C175 VDD2.n141 VSUBS 2.15308f
C176 VN.t4 VSUBS 0.823039f
C177 VN.n0 VSUBS 0.328463f
C178 VN.t0 VSUBS 0.806563f
C179 VN.n1 VSUBS 0.338099f
C180 VN.t3 VSUBS 0.81364f
C181 VN.n2 VSUBS 0.337363f
C182 VN.n3 VSUBS 0.196104f
C183 VN.t2 VSUBS 0.823039f
C184 VN.n4 VSUBS 0.328463f
C185 VN.t1 VSUBS 0.81364f
C186 VN.t5 VSUBS 0.806563f
C187 VN.n5 VSUBS 0.338099f
C188 VN.n6 VSUBS 0.337363f
C189 VN.n7 VSUBS 2.81905f
C190 B.n0 VSUBS 0.004804f
C191 B.n1 VSUBS 0.004804f
C192 B.n2 VSUBS 0.007597f
C193 B.n3 VSUBS 0.007597f
C194 B.n4 VSUBS 0.007597f
C195 B.n5 VSUBS 0.007597f
C196 B.n6 VSUBS 0.007597f
C197 B.n7 VSUBS 0.007597f
C198 B.n8 VSUBS 0.007597f
C199 B.n9 VSUBS 0.007597f
C200 B.n10 VSUBS 0.018257f
C201 B.n11 VSUBS 0.007597f
C202 B.n12 VSUBS 0.007597f
C203 B.n13 VSUBS 0.007597f
C204 B.n14 VSUBS 0.007597f
C205 B.n15 VSUBS 0.007597f
C206 B.n16 VSUBS 0.007597f
C207 B.n17 VSUBS 0.007597f
C208 B.n18 VSUBS 0.007597f
C209 B.n19 VSUBS 0.007597f
C210 B.n20 VSUBS 0.007597f
C211 B.n21 VSUBS 0.007597f
C212 B.n22 VSUBS 0.007597f
C213 B.n23 VSUBS 0.007597f
C214 B.n24 VSUBS 0.007597f
C215 B.n25 VSUBS 0.007597f
C216 B.n26 VSUBS 0.007597f
C217 B.n27 VSUBS 0.007597f
C218 B.n28 VSUBS 0.007597f
C219 B.n29 VSUBS 0.007597f
C220 B.n30 VSUBS 0.007597f
C221 B.n31 VSUBS 0.007597f
C222 B.t2 VSUBS 0.243849f
C223 B.t1 VSUBS 0.252237f
C224 B.t0 VSUBS 0.177948f
C225 B.n32 VSUBS 0.314223f
C226 B.n33 VSUBS 0.272576f
C227 B.n34 VSUBS 0.007597f
C228 B.n35 VSUBS 0.007597f
C229 B.n36 VSUBS 0.007597f
C230 B.n37 VSUBS 0.007597f
C231 B.n38 VSUBS 0.004245f
C232 B.n39 VSUBS 0.007597f
C233 B.t5 VSUBS 0.243852f
C234 B.t4 VSUBS 0.25224f
C235 B.t3 VSUBS 0.177948f
C236 B.n40 VSUBS 0.31422f
C237 B.n41 VSUBS 0.272573f
C238 B.n42 VSUBS 0.0176f
C239 B.n43 VSUBS 0.007597f
C240 B.n44 VSUBS 0.007597f
C241 B.n45 VSUBS 0.007597f
C242 B.n46 VSUBS 0.007597f
C243 B.n47 VSUBS 0.007597f
C244 B.n48 VSUBS 0.007597f
C245 B.n49 VSUBS 0.007597f
C246 B.n50 VSUBS 0.007597f
C247 B.n51 VSUBS 0.007597f
C248 B.n52 VSUBS 0.007597f
C249 B.n53 VSUBS 0.007597f
C250 B.n54 VSUBS 0.007597f
C251 B.n55 VSUBS 0.007597f
C252 B.n56 VSUBS 0.007597f
C253 B.n57 VSUBS 0.007597f
C254 B.n58 VSUBS 0.007597f
C255 B.n59 VSUBS 0.007597f
C256 B.n60 VSUBS 0.007597f
C257 B.n61 VSUBS 0.007597f
C258 B.n62 VSUBS 0.007597f
C259 B.n63 VSUBS 0.018811f
C260 B.n64 VSUBS 0.007597f
C261 B.n65 VSUBS 0.007597f
C262 B.n66 VSUBS 0.007597f
C263 B.n67 VSUBS 0.007597f
C264 B.n68 VSUBS 0.007597f
C265 B.n69 VSUBS 0.007597f
C266 B.n70 VSUBS 0.007597f
C267 B.n71 VSUBS 0.007597f
C268 B.n72 VSUBS 0.007597f
C269 B.n73 VSUBS 0.007597f
C270 B.n74 VSUBS 0.007597f
C271 B.n75 VSUBS 0.007597f
C272 B.n76 VSUBS 0.007597f
C273 B.n77 VSUBS 0.007597f
C274 B.n78 VSUBS 0.007597f
C275 B.n79 VSUBS 0.017938f
C276 B.n80 VSUBS 0.007597f
C277 B.n81 VSUBS 0.007597f
C278 B.n82 VSUBS 0.007597f
C279 B.n83 VSUBS 0.007597f
C280 B.n84 VSUBS 0.007597f
C281 B.n85 VSUBS 0.007597f
C282 B.n86 VSUBS 0.007597f
C283 B.n87 VSUBS 0.007597f
C284 B.n88 VSUBS 0.007597f
C285 B.n89 VSUBS 0.007597f
C286 B.n90 VSUBS 0.007597f
C287 B.n91 VSUBS 0.007597f
C288 B.n92 VSUBS 0.007597f
C289 B.n93 VSUBS 0.007597f
C290 B.n94 VSUBS 0.007597f
C291 B.n95 VSUBS 0.007597f
C292 B.n96 VSUBS 0.007597f
C293 B.n97 VSUBS 0.007597f
C294 B.n98 VSUBS 0.007597f
C295 B.n99 VSUBS 0.007597f
C296 B.n100 VSUBS 0.007597f
C297 B.t7 VSUBS 0.243852f
C298 B.t8 VSUBS 0.25224f
C299 B.t6 VSUBS 0.177948f
C300 B.n101 VSUBS 0.31422f
C301 B.n102 VSUBS 0.272573f
C302 B.n103 VSUBS 0.0176f
C303 B.n104 VSUBS 0.007597f
C304 B.n105 VSUBS 0.007597f
C305 B.n106 VSUBS 0.007597f
C306 B.n107 VSUBS 0.007597f
C307 B.n108 VSUBS 0.007597f
C308 B.t10 VSUBS 0.243849f
C309 B.t11 VSUBS 0.252237f
C310 B.t9 VSUBS 0.177948f
C311 B.n109 VSUBS 0.314223f
C312 B.n110 VSUBS 0.272576f
C313 B.n111 VSUBS 0.007597f
C314 B.n112 VSUBS 0.007597f
C315 B.n113 VSUBS 0.007597f
C316 B.n114 VSUBS 0.007597f
C317 B.n115 VSUBS 0.007597f
C318 B.n116 VSUBS 0.007597f
C319 B.n117 VSUBS 0.007597f
C320 B.n118 VSUBS 0.007597f
C321 B.n119 VSUBS 0.007597f
C322 B.n120 VSUBS 0.007597f
C323 B.n121 VSUBS 0.007597f
C324 B.n122 VSUBS 0.007597f
C325 B.n123 VSUBS 0.007597f
C326 B.n124 VSUBS 0.007597f
C327 B.n125 VSUBS 0.007597f
C328 B.n126 VSUBS 0.007597f
C329 B.n127 VSUBS 0.007597f
C330 B.n128 VSUBS 0.007597f
C331 B.n129 VSUBS 0.007597f
C332 B.n130 VSUBS 0.007597f
C333 B.n131 VSUBS 0.007597f
C334 B.n132 VSUBS 0.017938f
C335 B.n133 VSUBS 0.007597f
C336 B.n134 VSUBS 0.007597f
C337 B.n135 VSUBS 0.007597f
C338 B.n136 VSUBS 0.007597f
C339 B.n137 VSUBS 0.007597f
C340 B.n138 VSUBS 0.007597f
C341 B.n139 VSUBS 0.007597f
C342 B.n140 VSUBS 0.007597f
C343 B.n141 VSUBS 0.007597f
C344 B.n142 VSUBS 0.007597f
C345 B.n143 VSUBS 0.007597f
C346 B.n144 VSUBS 0.007597f
C347 B.n145 VSUBS 0.007597f
C348 B.n146 VSUBS 0.007597f
C349 B.n147 VSUBS 0.007597f
C350 B.n148 VSUBS 0.007597f
C351 B.n149 VSUBS 0.007597f
C352 B.n150 VSUBS 0.007597f
C353 B.n151 VSUBS 0.007597f
C354 B.n152 VSUBS 0.007597f
C355 B.n153 VSUBS 0.007597f
C356 B.n154 VSUBS 0.007597f
C357 B.n155 VSUBS 0.007597f
C358 B.n156 VSUBS 0.007597f
C359 B.n157 VSUBS 0.007597f
C360 B.n158 VSUBS 0.007597f
C361 B.n159 VSUBS 0.007597f
C362 B.n160 VSUBS 0.007597f
C363 B.n161 VSUBS 0.017938f
C364 B.n162 VSUBS 0.018257f
C365 B.n163 VSUBS 0.018257f
C366 B.n164 VSUBS 0.007597f
C367 B.n165 VSUBS 0.007597f
C368 B.n166 VSUBS 0.007597f
C369 B.n167 VSUBS 0.007597f
C370 B.n168 VSUBS 0.007597f
C371 B.n169 VSUBS 0.007597f
C372 B.n170 VSUBS 0.007597f
C373 B.n171 VSUBS 0.007597f
C374 B.n172 VSUBS 0.007597f
C375 B.n173 VSUBS 0.007597f
C376 B.n174 VSUBS 0.007597f
C377 B.n175 VSUBS 0.007597f
C378 B.n176 VSUBS 0.007597f
C379 B.n177 VSUBS 0.007597f
C380 B.n178 VSUBS 0.007597f
C381 B.n179 VSUBS 0.007597f
C382 B.n180 VSUBS 0.007597f
C383 B.n181 VSUBS 0.007597f
C384 B.n182 VSUBS 0.007597f
C385 B.n183 VSUBS 0.007597f
C386 B.n184 VSUBS 0.007597f
C387 B.n185 VSUBS 0.007597f
C388 B.n186 VSUBS 0.007597f
C389 B.n187 VSUBS 0.007597f
C390 B.n188 VSUBS 0.007597f
C391 B.n189 VSUBS 0.007597f
C392 B.n190 VSUBS 0.007597f
C393 B.n191 VSUBS 0.007597f
C394 B.n192 VSUBS 0.007597f
C395 B.n193 VSUBS 0.007597f
C396 B.n194 VSUBS 0.007597f
C397 B.n195 VSUBS 0.007597f
C398 B.n196 VSUBS 0.007597f
C399 B.n197 VSUBS 0.007597f
C400 B.n198 VSUBS 0.007597f
C401 B.n199 VSUBS 0.007597f
C402 B.n200 VSUBS 0.007597f
C403 B.n201 VSUBS 0.007597f
C404 B.n202 VSUBS 0.007597f
C405 B.n203 VSUBS 0.007597f
C406 B.n204 VSUBS 0.007597f
C407 B.n205 VSUBS 0.007597f
C408 B.n206 VSUBS 0.007597f
C409 B.n207 VSUBS 0.007597f
C410 B.n208 VSUBS 0.007597f
C411 B.n209 VSUBS 0.007597f
C412 B.n210 VSUBS 0.007597f
C413 B.n211 VSUBS 0.007597f
C414 B.n212 VSUBS 0.007597f
C415 B.n213 VSUBS 0.007597f
C416 B.n214 VSUBS 0.007597f
C417 B.n215 VSUBS 0.007597f
C418 B.n216 VSUBS 0.007597f
C419 B.n217 VSUBS 0.007597f
C420 B.n218 VSUBS 0.007597f
C421 B.n219 VSUBS 0.007597f
C422 B.n220 VSUBS 0.007597f
C423 B.n221 VSUBS 0.007597f
C424 B.n222 VSUBS 0.007597f
C425 B.n223 VSUBS 0.007597f
C426 B.n224 VSUBS 0.007597f
C427 B.n225 VSUBS 0.007597f
C428 B.n226 VSUBS 0.00715f
C429 B.n227 VSUBS 0.0176f
C430 B.n228 VSUBS 0.004245f
C431 B.n229 VSUBS 0.007597f
C432 B.n230 VSUBS 0.007597f
C433 B.n231 VSUBS 0.007597f
C434 B.n232 VSUBS 0.007597f
C435 B.n233 VSUBS 0.007597f
C436 B.n234 VSUBS 0.007597f
C437 B.n235 VSUBS 0.007597f
C438 B.n236 VSUBS 0.007597f
C439 B.n237 VSUBS 0.007597f
C440 B.n238 VSUBS 0.007597f
C441 B.n239 VSUBS 0.007597f
C442 B.n240 VSUBS 0.007597f
C443 B.n241 VSUBS 0.004245f
C444 B.n242 VSUBS 0.007597f
C445 B.n243 VSUBS 0.007597f
C446 B.n244 VSUBS 0.00715f
C447 B.n245 VSUBS 0.007597f
C448 B.n246 VSUBS 0.007597f
C449 B.n247 VSUBS 0.007597f
C450 B.n248 VSUBS 0.007597f
C451 B.n249 VSUBS 0.007597f
C452 B.n250 VSUBS 0.007597f
C453 B.n251 VSUBS 0.007597f
C454 B.n252 VSUBS 0.007597f
C455 B.n253 VSUBS 0.007597f
C456 B.n254 VSUBS 0.007597f
C457 B.n255 VSUBS 0.007597f
C458 B.n256 VSUBS 0.007597f
C459 B.n257 VSUBS 0.007597f
C460 B.n258 VSUBS 0.007597f
C461 B.n259 VSUBS 0.007597f
C462 B.n260 VSUBS 0.007597f
C463 B.n261 VSUBS 0.007597f
C464 B.n262 VSUBS 0.007597f
C465 B.n263 VSUBS 0.007597f
C466 B.n264 VSUBS 0.007597f
C467 B.n265 VSUBS 0.007597f
C468 B.n266 VSUBS 0.007597f
C469 B.n267 VSUBS 0.007597f
C470 B.n268 VSUBS 0.007597f
C471 B.n269 VSUBS 0.007597f
C472 B.n270 VSUBS 0.007597f
C473 B.n271 VSUBS 0.007597f
C474 B.n272 VSUBS 0.007597f
C475 B.n273 VSUBS 0.007597f
C476 B.n274 VSUBS 0.007597f
C477 B.n275 VSUBS 0.007597f
C478 B.n276 VSUBS 0.007597f
C479 B.n277 VSUBS 0.007597f
C480 B.n278 VSUBS 0.007597f
C481 B.n279 VSUBS 0.007597f
C482 B.n280 VSUBS 0.007597f
C483 B.n281 VSUBS 0.007597f
C484 B.n282 VSUBS 0.007597f
C485 B.n283 VSUBS 0.007597f
C486 B.n284 VSUBS 0.007597f
C487 B.n285 VSUBS 0.007597f
C488 B.n286 VSUBS 0.007597f
C489 B.n287 VSUBS 0.007597f
C490 B.n288 VSUBS 0.007597f
C491 B.n289 VSUBS 0.007597f
C492 B.n290 VSUBS 0.007597f
C493 B.n291 VSUBS 0.007597f
C494 B.n292 VSUBS 0.007597f
C495 B.n293 VSUBS 0.007597f
C496 B.n294 VSUBS 0.007597f
C497 B.n295 VSUBS 0.007597f
C498 B.n296 VSUBS 0.007597f
C499 B.n297 VSUBS 0.007597f
C500 B.n298 VSUBS 0.007597f
C501 B.n299 VSUBS 0.007597f
C502 B.n300 VSUBS 0.007597f
C503 B.n301 VSUBS 0.007597f
C504 B.n302 VSUBS 0.007597f
C505 B.n303 VSUBS 0.007597f
C506 B.n304 VSUBS 0.007597f
C507 B.n305 VSUBS 0.007597f
C508 B.n306 VSUBS 0.018257f
C509 B.n307 VSUBS 0.018257f
C510 B.n308 VSUBS 0.017938f
C511 B.n309 VSUBS 0.007597f
C512 B.n310 VSUBS 0.007597f
C513 B.n311 VSUBS 0.007597f
C514 B.n312 VSUBS 0.007597f
C515 B.n313 VSUBS 0.007597f
C516 B.n314 VSUBS 0.007597f
C517 B.n315 VSUBS 0.007597f
C518 B.n316 VSUBS 0.007597f
C519 B.n317 VSUBS 0.007597f
C520 B.n318 VSUBS 0.007597f
C521 B.n319 VSUBS 0.007597f
C522 B.n320 VSUBS 0.007597f
C523 B.n321 VSUBS 0.007597f
C524 B.n322 VSUBS 0.007597f
C525 B.n323 VSUBS 0.007597f
C526 B.n324 VSUBS 0.007597f
C527 B.n325 VSUBS 0.007597f
C528 B.n326 VSUBS 0.007597f
C529 B.n327 VSUBS 0.007597f
C530 B.n328 VSUBS 0.007597f
C531 B.n329 VSUBS 0.007597f
C532 B.n330 VSUBS 0.007597f
C533 B.n331 VSUBS 0.007597f
C534 B.n332 VSUBS 0.007597f
C535 B.n333 VSUBS 0.007597f
C536 B.n334 VSUBS 0.007597f
C537 B.n335 VSUBS 0.007597f
C538 B.n336 VSUBS 0.007597f
C539 B.n337 VSUBS 0.007597f
C540 B.n338 VSUBS 0.007597f
C541 B.n339 VSUBS 0.007597f
C542 B.n340 VSUBS 0.007597f
C543 B.n341 VSUBS 0.007597f
C544 B.n342 VSUBS 0.007597f
C545 B.n343 VSUBS 0.007597f
C546 B.n344 VSUBS 0.007597f
C547 B.n345 VSUBS 0.007597f
C548 B.n346 VSUBS 0.007597f
C549 B.n347 VSUBS 0.007597f
C550 B.n348 VSUBS 0.007597f
C551 B.n349 VSUBS 0.007597f
C552 B.n350 VSUBS 0.007597f
C553 B.n351 VSUBS 0.007597f
C554 B.n352 VSUBS 0.007597f
C555 B.n353 VSUBS 0.007597f
C556 B.n354 VSUBS 0.007597f
C557 B.n355 VSUBS 0.007597f
C558 B.n356 VSUBS 0.017938f
C559 B.n357 VSUBS 0.018257f
C560 B.n358 VSUBS 0.017384f
C561 B.n359 VSUBS 0.007597f
C562 B.n360 VSUBS 0.007597f
C563 B.n361 VSUBS 0.007597f
C564 B.n362 VSUBS 0.007597f
C565 B.n363 VSUBS 0.007597f
C566 B.n364 VSUBS 0.007597f
C567 B.n365 VSUBS 0.007597f
C568 B.n366 VSUBS 0.007597f
C569 B.n367 VSUBS 0.007597f
C570 B.n368 VSUBS 0.007597f
C571 B.n369 VSUBS 0.007597f
C572 B.n370 VSUBS 0.007597f
C573 B.n371 VSUBS 0.007597f
C574 B.n372 VSUBS 0.007597f
C575 B.n373 VSUBS 0.007597f
C576 B.n374 VSUBS 0.007597f
C577 B.n375 VSUBS 0.007597f
C578 B.n376 VSUBS 0.007597f
C579 B.n377 VSUBS 0.007597f
C580 B.n378 VSUBS 0.007597f
C581 B.n379 VSUBS 0.007597f
C582 B.n380 VSUBS 0.007597f
C583 B.n381 VSUBS 0.007597f
C584 B.n382 VSUBS 0.007597f
C585 B.n383 VSUBS 0.007597f
C586 B.n384 VSUBS 0.007597f
C587 B.n385 VSUBS 0.007597f
C588 B.n386 VSUBS 0.007597f
C589 B.n387 VSUBS 0.007597f
C590 B.n388 VSUBS 0.007597f
C591 B.n389 VSUBS 0.007597f
C592 B.n390 VSUBS 0.007597f
C593 B.n391 VSUBS 0.007597f
C594 B.n392 VSUBS 0.007597f
C595 B.n393 VSUBS 0.007597f
C596 B.n394 VSUBS 0.007597f
C597 B.n395 VSUBS 0.007597f
C598 B.n396 VSUBS 0.007597f
C599 B.n397 VSUBS 0.007597f
C600 B.n398 VSUBS 0.007597f
C601 B.n399 VSUBS 0.007597f
C602 B.n400 VSUBS 0.007597f
C603 B.n401 VSUBS 0.007597f
C604 B.n402 VSUBS 0.007597f
C605 B.n403 VSUBS 0.007597f
C606 B.n404 VSUBS 0.007597f
C607 B.n405 VSUBS 0.007597f
C608 B.n406 VSUBS 0.007597f
C609 B.n407 VSUBS 0.007597f
C610 B.n408 VSUBS 0.007597f
C611 B.n409 VSUBS 0.007597f
C612 B.n410 VSUBS 0.007597f
C613 B.n411 VSUBS 0.007597f
C614 B.n412 VSUBS 0.007597f
C615 B.n413 VSUBS 0.007597f
C616 B.n414 VSUBS 0.007597f
C617 B.n415 VSUBS 0.007597f
C618 B.n416 VSUBS 0.007597f
C619 B.n417 VSUBS 0.007597f
C620 B.n418 VSUBS 0.007597f
C621 B.n419 VSUBS 0.007597f
C622 B.n420 VSUBS 0.00715f
C623 B.n421 VSUBS 0.007597f
C624 B.n422 VSUBS 0.007597f
C625 B.n423 VSUBS 0.007597f
C626 B.n424 VSUBS 0.007597f
C627 B.n425 VSUBS 0.007597f
C628 B.n426 VSUBS 0.007597f
C629 B.n427 VSUBS 0.007597f
C630 B.n428 VSUBS 0.007597f
C631 B.n429 VSUBS 0.007597f
C632 B.n430 VSUBS 0.007597f
C633 B.n431 VSUBS 0.007597f
C634 B.n432 VSUBS 0.007597f
C635 B.n433 VSUBS 0.007597f
C636 B.n434 VSUBS 0.007597f
C637 B.n435 VSUBS 0.007597f
C638 B.n436 VSUBS 0.004245f
C639 B.n437 VSUBS 0.0176f
C640 B.n438 VSUBS 0.00715f
C641 B.n439 VSUBS 0.007597f
C642 B.n440 VSUBS 0.007597f
C643 B.n441 VSUBS 0.007597f
C644 B.n442 VSUBS 0.007597f
C645 B.n443 VSUBS 0.007597f
C646 B.n444 VSUBS 0.007597f
C647 B.n445 VSUBS 0.007597f
C648 B.n446 VSUBS 0.007597f
C649 B.n447 VSUBS 0.007597f
C650 B.n448 VSUBS 0.007597f
C651 B.n449 VSUBS 0.007597f
C652 B.n450 VSUBS 0.007597f
C653 B.n451 VSUBS 0.007597f
C654 B.n452 VSUBS 0.007597f
C655 B.n453 VSUBS 0.007597f
C656 B.n454 VSUBS 0.007597f
C657 B.n455 VSUBS 0.007597f
C658 B.n456 VSUBS 0.007597f
C659 B.n457 VSUBS 0.007597f
C660 B.n458 VSUBS 0.007597f
C661 B.n459 VSUBS 0.007597f
C662 B.n460 VSUBS 0.007597f
C663 B.n461 VSUBS 0.007597f
C664 B.n462 VSUBS 0.007597f
C665 B.n463 VSUBS 0.007597f
C666 B.n464 VSUBS 0.007597f
C667 B.n465 VSUBS 0.007597f
C668 B.n466 VSUBS 0.007597f
C669 B.n467 VSUBS 0.007597f
C670 B.n468 VSUBS 0.007597f
C671 B.n469 VSUBS 0.007597f
C672 B.n470 VSUBS 0.007597f
C673 B.n471 VSUBS 0.007597f
C674 B.n472 VSUBS 0.007597f
C675 B.n473 VSUBS 0.007597f
C676 B.n474 VSUBS 0.007597f
C677 B.n475 VSUBS 0.007597f
C678 B.n476 VSUBS 0.007597f
C679 B.n477 VSUBS 0.007597f
C680 B.n478 VSUBS 0.007597f
C681 B.n479 VSUBS 0.007597f
C682 B.n480 VSUBS 0.007597f
C683 B.n481 VSUBS 0.007597f
C684 B.n482 VSUBS 0.007597f
C685 B.n483 VSUBS 0.007597f
C686 B.n484 VSUBS 0.007597f
C687 B.n485 VSUBS 0.007597f
C688 B.n486 VSUBS 0.007597f
C689 B.n487 VSUBS 0.007597f
C690 B.n488 VSUBS 0.007597f
C691 B.n489 VSUBS 0.007597f
C692 B.n490 VSUBS 0.007597f
C693 B.n491 VSUBS 0.007597f
C694 B.n492 VSUBS 0.007597f
C695 B.n493 VSUBS 0.007597f
C696 B.n494 VSUBS 0.007597f
C697 B.n495 VSUBS 0.007597f
C698 B.n496 VSUBS 0.007597f
C699 B.n497 VSUBS 0.007597f
C700 B.n498 VSUBS 0.007597f
C701 B.n499 VSUBS 0.007597f
C702 B.n500 VSUBS 0.007597f
C703 B.n501 VSUBS 0.018257f
C704 B.n502 VSUBS 0.017938f
C705 B.n503 VSUBS 0.017938f
C706 B.n504 VSUBS 0.007597f
C707 B.n505 VSUBS 0.007597f
C708 B.n506 VSUBS 0.007597f
C709 B.n507 VSUBS 0.007597f
C710 B.n508 VSUBS 0.007597f
C711 B.n509 VSUBS 0.007597f
C712 B.n510 VSUBS 0.007597f
C713 B.n511 VSUBS 0.007597f
C714 B.n512 VSUBS 0.007597f
C715 B.n513 VSUBS 0.007597f
C716 B.n514 VSUBS 0.007597f
C717 B.n515 VSUBS 0.007597f
C718 B.n516 VSUBS 0.007597f
C719 B.n517 VSUBS 0.007597f
C720 B.n518 VSUBS 0.007597f
C721 B.n519 VSUBS 0.007597f
C722 B.n520 VSUBS 0.007597f
C723 B.n521 VSUBS 0.007597f
C724 B.n522 VSUBS 0.007597f
C725 B.n523 VSUBS 0.007597f
C726 B.n524 VSUBS 0.007597f
C727 B.n525 VSUBS 0.007597f
C728 B.n526 VSUBS 0.007597f
C729 B.n527 VSUBS 0.017201f
C730 VDD1.n0 VSUBS 0.015275f
C731 VDD1.n1 VSUBS 0.034495f
C732 VDD1.n2 VSUBS 0.015452f
C733 VDD1.n3 VSUBS 0.027159f
C734 VDD1.n4 VSUBS 0.014594f
C735 VDD1.n5 VSUBS 0.034495f
C736 VDD1.n6 VSUBS 0.015452f
C737 VDD1.n7 VSUBS 0.027159f
C738 VDD1.n8 VSUBS 0.014594f
C739 VDD1.n9 VSUBS 0.034495f
C740 VDD1.n10 VSUBS 0.015452f
C741 VDD1.n11 VSUBS 0.027159f
C742 VDD1.n12 VSUBS 0.014594f
C743 VDD1.n13 VSUBS 0.034495f
C744 VDD1.n14 VSUBS 0.015452f
C745 VDD1.n15 VSUBS 0.027159f
C746 VDD1.n16 VSUBS 0.014594f
C747 VDD1.n17 VSUBS 0.034495f
C748 VDD1.n18 VSUBS 0.015452f
C749 VDD1.n19 VSUBS 0.027159f
C750 VDD1.n20 VSUBS 0.014594f
C751 VDD1.n21 VSUBS 0.025871f
C752 VDD1.n22 VSUBS 0.021944f
C753 VDD1.t5 VSUBS 0.073688f
C754 VDD1.n23 VSUBS 0.172382f
C755 VDD1.n24 VSUBS 1.44069f
C756 VDD1.n25 VSUBS 0.014594f
C757 VDD1.n26 VSUBS 0.015452f
C758 VDD1.n27 VSUBS 0.034495f
C759 VDD1.n28 VSUBS 0.034495f
C760 VDD1.n29 VSUBS 0.015452f
C761 VDD1.n30 VSUBS 0.014594f
C762 VDD1.n31 VSUBS 0.027159f
C763 VDD1.n32 VSUBS 0.027159f
C764 VDD1.n33 VSUBS 0.014594f
C765 VDD1.n34 VSUBS 0.015452f
C766 VDD1.n35 VSUBS 0.034495f
C767 VDD1.n36 VSUBS 0.034495f
C768 VDD1.n37 VSUBS 0.015452f
C769 VDD1.n38 VSUBS 0.014594f
C770 VDD1.n39 VSUBS 0.027159f
C771 VDD1.n40 VSUBS 0.027159f
C772 VDD1.n41 VSUBS 0.014594f
C773 VDD1.n42 VSUBS 0.015452f
C774 VDD1.n43 VSUBS 0.034495f
C775 VDD1.n44 VSUBS 0.034495f
C776 VDD1.n45 VSUBS 0.015452f
C777 VDD1.n46 VSUBS 0.014594f
C778 VDD1.n47 VSUBS 0.027159f
C779 VDD1.n48 VSUBS 0.027159f
C780 VDD1.n49 VSUBS 0.014594f
C781 VDD1.n50 VSUBS 0.015452f
C782 VDD1.n51 VSUBS 0.034495f
C783 VDD1.n52 VSUBS 0.034495f
C784 VDD1.n53 VSUBS 0.015452f
C785 VDD1.n54 VSUBS 0.014594f
C786 VDD1.n55 VSUBS 0.027159f
C787 VDD1.n56 VSUBS 0.027159f
C788 VDD1.n57 VSUBS 0.014594f
C789 VDD1.n58 VSUBS 0.015452f
C790 VDD1.n59 VSUBS 0.034495f
C791 VDD1.n60 VSUBS 0.034495f
C792 VDD1.n61 VSUBS 0.015452f
C793 VDD1.n62 VSUBS 0.014594f
C794 VDD1.n63 VSUBS 0.027159f
C795 VDD1.n64 VSUBS 0.06797f
C796 VDD1.n65 VSUBS 0.014594f
C797 VDD1.n66 VSUBS 0.015452f
C798 VDD1.n67 VSUBS 0.076062f
C799 VDD1.n68 VSUBS 0.06965f
C800 VDD1.n69 VSUBS 0.015275f
C801 VDD1.n70 VSUBS 0.034495f
C802 VDD1.n71 VSUBS 0.015452f
C803 VDD1.n72 VSUBS 0.027159f
C804 VDD1.n73 VSUBS 0.014594f
C805 VDD1.n74 VSUBS 0.034495f
C806 VDD1.n75 VSUBS 0.015452f
C807 VDD1.n76 VSUBS 0.027159f
C808 VDD1.n77 VSUBS 0.014594f
C809 VDD1.n78 VSUBS 0.034495f
C810 VDD1.n79 VSUBS 0.015452f
C811 VDD1.n80 VSUBS 0.027159f
C812 VDD1.n81 VSUBS 0.014594f
C813 VDD1.n82 VSUBS 0.034495f
C814 VDD1.n83 VSUBS 0.015452f
C815 VDD1.n84 VSUBS 0.027159f
C816 VDD1.n85 VSUBS 0.014594f
C817 VDD1.n86 VSUBS 0.034495f
C818 VDD1.n87 VSUBS 0.015452f
C819 VDD1.n88 VSUBS 0.027159f
C820 VDD1.n89 VSUBS 0.014594f
C821 VDD1.n90 VSUBS 0.025871f
C822 VDD1.n91 VSUBS 0.021944f
C823 VDD1.t1 VSUBS 0.073688f
C824 VDD1.n92 VSUBS 0.172382f
C825 VDD1.n93 VSUBS 1.44069f
C826 VDD1.n94 VSUBS 0.014594f
C827 VDD1.n95 VSUBS 0.015452f
C828 VDD1.n96 VSUBS 0.034495f
C829 VDD1.n97 VSUBS 0.034495f
C830 VDD1.n98 VSUBS 0.015452f
C831 VDD1.n99 VSUBS 0.014594f
C832 VDD1.n100 VSUBS 0.027159f
C833 VDD1.n101 VSUBS 0.027159f
C834 VDD1.n102 VSUBS 0.014594f
C835 VDD1.n103 VSUBS 0.015452f
C836 VDD1.n104 VSUBS 0.034495f
C837 VDD1.n105 VSUBS 0.034495f
C838 VDD1.n106 VSUBS 0.015452f
C839 VDD1.n107 VSUBS 0.014594f
C840 VDD1.n108 VSUBS 0.027159f
C841 VDD1.n109 VSUBS 0.027159f
C842 VDD1.n110 VSUBS 0.014594f
C843 VDD1.n111 VSUBS 0.015452f
C844 VDD1.n112 VSUBS 0.034495f
C845 VDD1.n113 VSUBS 0.034495f
C846 VDD1.n114 VSUBS 0.015452f
C847 VDD1.n115 VSUBS 0.014594f
C848 VDD1.n116 VSUBS 0.027159f
C849 VDD1.n117 VSUBS 0.027159f
C850 VDD1.n118 VSUBS 0.014594f
C851 VDD1.n119 VSUBS 0.015452f
C852 VDD1.n120 VSUBS 0.034495f
C853 VDD1.n121 VSUBS 0.034495f
C854 VDD1.n122 VSUBS 0.015452f
C855 VDD1.n123 VSUBS 0.014594f
C856 VDD1.n124 VSUBS 0.027159f
C857 VDD1.n125 VSUBS 0.027159f
C858 VDD1.n126 VSUBS 0.014594f
C859 VDD1.n127 VSUBS 0.015452f
C860 VDD1.n128 VSUBS 0.034495f
C861 VDD1.n129 VSUBS 0.034495f
C862 VDD1.n130 VSUBS 0.015452f
C863 VDD1.n131 VSUBS 0.014594f
C864 VDD1.n132 VSUBS 0.027159f
C865 VDD1.n133 VSUBS 0.06797f
C866 VDD1.n134 VSUBS 0.014594f
C867 VDD1.n135 VSUBS 0.015452f
C868 VDD1.n136 VSUBS 0.076062f
C869 VDD1.n137 VSUBS 0.069378f
C870 VDD1.t0 VSUBS 0.270845f
C871 VDD1.t4 VSUBS 0.270845f
C872 VDD1.n138 VSUBS 2.15308f
C873 VDD1.n139 VSUBS 2.22452f
C874 VDD1.t3 VSUBS 0.270845f
C875 VDD1.t2 VSUBS 0.270845f
C876 VDD1.n140 VSUBS 2.15241f
C877 VDD1.n141 VSUBS 2.65689f
C878 VTAIL.t1 VSUBS 0.324264f
C879 VTAIL.t5 VSUBS 0.324264f
C880 VTAIL.n0 VSUBS 2.41069f
C881 VTAIL.n1 VSUBS 0.813304f
C882 VTAIL.n2 VSUBS 0.018288f
C883 VTAIL.n3 VSUBS 0.041298f
C884 VTAIL.n4 VSUBS 0.0185f
C885 VTAIL.n5 VSUBS 0.032515f
C886 VTAIL.n6 VSUBS 0.017472f
C887 VTAIL.n7 VSUBS 0.041298f
C888 VTAIL.n8 VSUBS 0.0185f
C889 VTAIL.n9 VSUBS 0.032515f
C890 VTAIL.n10 VSUBS 0.017472f
C891 VTAIL.n11 VSUBS 0.041298f
C892 VTAIL.n12 VSUBS 0.0185f
C893 VTAIL.n13 VSUBS 0.032515f
C894 VTAIL.n14 VSUBS 0.017472f
C895 VTAIL.n15 VSUBS 0.041298f
C896 VTAIL.n16 VSUBS 0.0185f
C897 VTAIL.n17 VSUBS 0.032515f
C898 VTAIL.n18 VSUBS 0.017472f
C899 VTAIL.n19 VSUBS 0.041298f
C900 VTAIL.n20 VSUBS 0.0185f
C901 VTAIL.n21 VSUBS 0.032515f
C902 VTAIL.n22 VSUBS 0.017472f
C903 VTAIL.n23 VSUBS 0.030973f
C904 VTAIL.n24 VSUBS 0.026272f
C905 VTAIL.t8 VSUBS 0.088221f
C906 VTAIL.n25 VSUBS 0.206381f
C907 VTAIL.n26 VSUBS 1.72484f
C908 VTAIL.n27 VSUBS 0.017472f
C909 VTAIL.n28 VSUBS 0.0185f
C910 VTAIL.n29 VSUBS 0.041298f
C911 VTAIL.n30 VSUBS 0.041298f
C912 VTAIL.n31 VSUBS 0.0185f
C913 VTAIL.n32 VSUBS 0.017472f
C914 VTAIL.n33 VSUBS 0.032515f
C915 VTAIL.n34 VSUBS 0.032515f
C916 VTAIL.n35 VSUBS 0.017472f
C917 VTAIL.n36 VSUBS 0.0185f
C918 VTAIL.n37 VSUBS 0.041298f
C919 VTAIL.n38 VSUBS 0.041298f
C920 VTAIL.n39 VSUBS 0.0185f
C921 VTAIL.n40 VSUBS 0.017472f
C922 VTAIL.n41 VSUBS 0.032515f
C923 VTAIL.n42 VSUBS 0.032515f
C924 VTAIL.n43 VSUBS 0.017472f
C925 VTAIL.n44 VSUBS 0.0185f
C926 VTAIL.n45 VSUBS 0.041298f
C927 VTAIL.n46 VSUBS 0.041298f
C928 VTAIL.n47 VSUBS 0.0185f
C929 VTAIL.n48 VSUBS 0.017472f
C930 VTAIL.n49 VSUBS 0.032515f
C931 VTAIL.n50 VSUBS 0.032515f
C932 VTAIL.n51 VSUBS 0.017472f
C933 VTAIL.n52 VSUBS 0.0185f
C934 VTAIL.n53 VSUBS 0.041298f
C935 VTAIL.n54 VSUBS 0.041298f
C936 VTAIL.n55 VSUBS 0.0185f
C937 VTAIL.n56 VSUBS 0.017472f
C938 VTAIL.n57 VSUBS 0.032515f
C939 VTAIL.n58 VSUBS 0.032515f
C940 VTAIL.n59 VSUBS 0.017472f
C941 VTAIL.n60 VSUBS 0.0185f
C942 VTAIL.n61 VSUBS 0.041298f
C943 VTAIL.n62 VSUBS 0.041298f
C944 VTAIL.n63 VSUBS 0.0185f
C945 VTAIL.n64 VSUBS 0.017472f
C946 VTAIL.n65 VSUBS 0.032515f
C947 VTAIL.n66 VSUBS 0.081376f
C948 VTAIL.n67 VSUBS 0.017472f
C949 VTAIL.n68 VSUBS 0.0185f
C950 VTAIL.n69 VSUBS 0.091064f
C951 VTAIL.n70 VSUBS 0.059882f
C952 VTAIL.n71 VSUBS 0.169425f
C953 VTAIL.t10 VSUBS 0.324264f
C954 VTAIL.t7 VSUBS 0.324264f
C955 VTAIL.n72 VSUBS 2.41069f
C956 VTAIL.n73 VSUBS 2.47363f
C957 VTAIL.t0 VSUBS 0.324264f
C958 VTAIL.t2 VSUBS 0.324264f
C959 VTAIL.n74 VSUBS 2.41069f
C960 VTAIL.n75 VSUBS 2.47362f
C961 VTAIL.n76 VSUBS 0.018288f
C962 VTAIL.n77 VSUBS 0.041298f
C963 VTAIL.n78 VSUBS 0.0185f
C964 VTAIL.n79 VSUBS 0.032515f
C965 VTAIL.n80 VSUBS 0.017472f
C966 VTAIL.n81 VSUBS 0.041298f
C967 VTAIL.n82 VSUBS 0.0185f
C968 VTAIL.n83 VSUBS 0.032515f
C969 VTAIL.n84 VSUBS 0.017472f
C970 VTAIL.n85 VSUBS 0.041298f
C971 VTAIL.n86 VSUBS 0.0185f
C972 VTAIL.n87 VSUBS 0.032515f
C973 VTAIL.n88 VSUBS 0.017472f
C974 VTAIL.n89 VSUBS 0.041298f
C975 VTAIL.n90 VSUBS 0.0185f
C976 VTAIL.n91 VSUBS 0.032515f
C977 VTAIL.n92 VSUBS 0.017472f
C978 VTAIL.n93 VSUBS 0.041298f
C979 VTAIL.n94 VSUBS 0.0185f
C980 VTAIL.n95 VSUBS 0.032515f
C981 VTAIL.n96 VSUBS 0.017472f
C982 VTAIL.n97 VSUBS 0.030973f
C983 VTAIL.n98 VSUBS 0.026272f
C984 VTAIL.t4 VSUBS 0.088221f
C985 VTAIL.n99 VSUBS 0.206381f
C986 VTAIL.n100 VSUBS 1.72484f
C987 VTAIL.n101 VSUBS 0.017472f
C988 VTAIL.n102 VSUBS 0.0185f
C989 VTAIL.n103 VSUBS 0.041298f
C990 VTAIL.n104 VSUBS 0.041298f
C991 VTAIL.n105 VSUBS 0.0185f
C992 VTAIL.n106 VSUBS 0.017472f
C993 VTAIL.n107 VSUBS 0.032515f
C994 VTAIL.n108 VSUBS 0.032515f
C995 VTAIL.n109 VSUBS 0.017472f
C996 VTAIL.n110 VSUBS 0.0185f
C997 VTAIL.n111 VSUBS 0.041298f
C998 VTAIL.n112 VSUBS 0.041298f
C999 VTAIL.n113 VSUBS 0.0185f
C1000 VTAIL.n114 VSUBS 0.017472f
C1001 VTAIL.n115 VSUBS 0.032515f
C1002 VTAIL.n116 VSUBS 0.032515f
C1003 VTAIL.n117 VSUBS 0.017472f
C1004 VTAIL.n118 VSUBS 0.0185f
C1005 VTAIL.n119 VSUBS 0.041298f
C1006 VTAIL.n120 VSUBS 0.041298f
C1007 VTAIL.n121 VSUBS 0.0185f
C1008 VTAIL.n122 VSUBS 0.017472f
C1009 VTAIL.n123 VSUBS 0.032515f
C1010 VTAIL.n124 VSUBS 0.032515f
C1011 VTAIL.n125 VSUBS 0.017472f
C1012 VTAIL.n126 VSUBS 0.0185f
C1013 VTAIL.n127 VSUBS 0.041298f
C1014 VTAIL.n128 VSUBS 0.041298f
C1015 VTAIL.n129 VSUBS 0.0185f
C1016 VTAIL.n130 VSUBS 0.017472f
C1017 VTAIL.n131 VSUBS 0.032515f
C1018 VTAIL.n132 VSUBS 0.032515f
C1019 VTAIL.n133 VSUBS 0.017472f
C1020 VTAIL.n134 VSUBS 0.0185f
C1021 VTAIL.n135 VSUBS 0.041298f
C1022 VTAIL.n136 VSUBS 0.041298f
C1023 VTAIL.n137 VSUBS 0.0185f
C1024 VTAIL.n138 VSUBS 0.017472f
C1025 VTAIL.n139 VSUBS 0.032515f
C1026 VTAIL.n140 VSUBS 0.081376f
C1027 VTAIL.n141 VSUBS 0.017472f
C1028 VTAIL.n142 VSUBS 0.0185f
C1029 VTAIL.n143 VSUBS 0.091064f
C1030 VTAIL.n144 VSUBS 0.059882f
C1031 VTAIL.n145 VSUBS 0.169425f
C1032 VTAIL.t11 VSUBS 0.324264f
C1033 VTAIL.t6 VSUBS 0.324264f
C1034 VTAIL.n146 VSUBS 2.41069f
C1035 VTAIL.n147 VSUBS 0.851911f
C1036 VTAIL.n148 VSUBS 0.018288f
C1037 VTAIL.n149 VSUBS 0.041298f
C1038 VTAIL.n150 VSUBS 0.0185f
C1039 VTAIL.n151 VSUBS 0.032515f
C1040 VTAIL.n152 VSUBS 0.017472f
C1041 VTAIL.n153 VSUBS 0.041298f
C1042 VTAIL.n154 VSUBS 0.0185f
C1043 VTAIL.n155 VSUBS 0.032515f
C1044 VTAIL.n156 VSUBS 0.017472f
C1045 VTAIL.n157 VSUBS 0.041298f
C1046 VTAIL.n158 VSUBS 0.0185f
C1047 VTAIL.n159 VSUBS 0.032515f
C1048 VTAIL.n160 VSUBS 0.017472f
C1049 VTAIL.n161 VSUBS 0.041298f
C1050 VTAIL.n162 VSUBS 0.0185f
C1051 VTAIL.n163 VSUBS 0.032515f
C1052 VTAIL.n164 VSUBS 0.017472f
C1053 VTAIL.n165 VSUBS 0.041298f
C1054 VTAIL.n166 VSUBS 0.0185f
C1055 VTAIL.n167 VSUBS 0.032515f
C1056 VTAIL.n168 VSUBS 0.017472f
C1057 VTAIL.n169 VSUBS 0.030973f
C1058 VTAIL.n170 VSUBS 0.026272f
C1059 VTAIL.t9 VSUBS 0.088221f
C1060 VTAIL.n171 VSUBS 0.206381f
C1061 VTAIL.n172 VSUBS 1.72484f
C1062 VTAIL.n173 VSUBS 0.017472f
C1063 VTAIL.n174 VSUBS 0.0185f
C1064 VTAIL.n175 VSUBS 0.041298f
C1065 VTAIL.n176 VSUBS 0.041298f
C1066 VTAIL.n177 VSUBS 0.0185f
C1067 VTAIL.n178 VSUBS 0.017472f
C1068 VTAIL.n179 VSUBS 0.032515f
C1069 VTAIL.n180 VSUBS 0.032515f
C1070 VTAIL.n181 VSUBS 0.017472f
C1071 VTAIL.n182 VSUBS 0.0185f
C1072 VTAIL.n183 VSUBS 0.041298f
C1073 VTAIL.n184 VSUBS 0.041298f
C1074 VTAIL.n185 VSUBS 0.0185f
C1075 VTAIL.n186 VSUBS 0.017472f
C1076 VTAIL.n187 VSUBS 0.032515f
C1077 VTAIL.n188 VSUBS 0.032515f
C1078 VTAIL.n189 VSUBS 0.017472f
C1079 VTAIL.n190 VSUBS 0.0185f
C1080 VTAIL.n191 VSUBS 0.041298f
C1081 VTAIL.n192 VSUBS 0.041298f
C1082 VTAIL.n193 VSUBS 0.0185f
C1083 VTAIL.n194 VSUBS 0.017472f
C1084 VTAIL.n195 VSUBS 0.032515f
C1085 VTAIL.n196 VSUBS 0.032515f
C1086 VTAIL.n197 VSUBS 0.017472f
C1087 VTAIL.n198 VSUBS 0.0185f
C1088 VTAIL.n199 VSUBS 0.041298f
C1089 VTAIL.n200 VSUBS 0.041298f
C1090 VTAIL.n201 VSUBS 0.0185f
C1091 VTAIL.n202 VSUBS 0.017472f
C1092 VTAIL.n203 VSUBS 0.032515f
C1093 VTAIL.n204 VSUBS 0.032515f
C1094 VTAIL.n205 VSUBS 0.017472f
C1095 VTAIL.n206 VSUBS 0.0185f
C1096 VTAIL.n207 VSUBS 0.041298f
C1097 VTAIL.n208 VSUBS 0.041298f
C1098 VTAIL.n209 VSUBS 0.0185f
C1099 VTAIL.n210 VSUBS 0.017472f
C1100 VTAIL.n211 VSUBS 0.032515f
C1101 VTAIL.n212 VSUBS 0.081376f
C1102 VTAIL.n213 VSUBS 0.017472f
C1103 VTAIL.n214 VSUBS 0.0185f
C1104 VTAIL.n215 VSUBS 0.091064f
C1105 VTAIL.n216 VSUBS 0.059882f
C1106 VTAIL.n217 VSUBS 1.73152f
C1107 VTAIL.n218 VSUBS 0.018288f
C1108 VTAIL.n219 VSUBS 0.041298f
C1109 VTAIL.n220 VSUBS 0.0185f
C1110 VTAIL.n221 VSUBS 0.032515f
C1111 VTAIL.n222 VSUBS 0.017472f
C1112 VTAIL.n223 VSUBS 0.041298f
C1113 VTAIL.n224 VSUBS 0.0185f
C1114 VTAIL.n225 VSUBS 0.032515f
C1115 VTAIL.n226 VSUBS 0.017472f
C1116 VTAIL.n227 VSUBS 0.041298f
C1117 VTAIL.n228 VSUBS 0.0185f
C1118 VTAIL.n229 VSUBS 0.032515f
C1119 VTAIL.n230 VSUBS 0.017472f
C1120 VTAIL.n231 VSUBS 0.041298f
C1121 VTAIL.n232 VSUBS 0.0185f
C1122 VTAIL.n233 VSUBS 0.032515f
C1123 VTAIL.n234 VSUBS 0.017472f
C1124 VTAIL.n235 VSUBS 0.041298f
C1125 VTAIL.n236 VSUBS 0.0185f
C1126 VTAIL.n237 VSUBS 0.032515f
C1127 VTAIL.n238 VSUBS 0.017472f
C1128 VTAIL.n239 VSUBS 0.030973f
C1129 VTAIL.n240 VSUBS 0.026272f
C1130 VTAIL.t3 VSUBS 0.088221f
C1131 VTAIL.n241 VSUBS 0.206381f
C1132 VTAIL.n242 VSUBS 1.72484f
C1133 VTAIL.n243 VSUBS 0.017472f
C1134 VTAIL.n244 VSUBS 0.0185f
C1135 VTAIL.n245 VSUBS 0.041298f
C1136 VTAIL.n246 VSUBS 0.041298f
C1137 VTAIL.n247 VSUBS 0.0185f
C1138 VTAIL.n248 VSUBS 0.017472f
C1139 VTAIL.n249 VSUBS 0.032515f
C1140 VTAIL.n250 VSUBS 0.032515f
C1141 VTAIL.n251 VSUBS 0.017472f
C1142 VTAIL.n252 VSUBS 0.0185f
C1143 VTAIL.n253 VSUBS 0.041298f
C1144 VTAIL.n254 VSUBS 0.041298f
C1145 VTAIL.n255 VSUBS 0.0185f
C1146 VTAIL.n256 VSUBS 0.017472f
C1147 VTAIL.n257 VSUBS 0.032515f
C1148 VTAIL.n258 VSUBS 0.032515f
C1149 VTAIL.n259 VSUBS 0.017472f
C1150 VTAIL.n260 VSUBS 0.0185f
C1151 VTAIL.n261 VSUBS 0.041298f
C1152 VTAIL.n262 VSUBS 0.041298f
C1153 VTAIL.n263 VSUBS 0.0185f
C1154 VTAIL.n264 VSUBS 0.017472f
C1155 VTAIL.n265 VSUBS 0.032515f
C1156 VTAIL.n266 VSUBS 0.032515f
C1157 VTAIL.n267 VSUBS 0.017472f
C1158 VTAIL.n268 VSUBS 0.0185f
C1159 VTAIL.n269 VSUBS 0.041298f
C1160 VTAIL.n270 VSUBS 0.041298f
C1161 VTAIL.n271 VSUBS 0.0185f
C1162 VTAIL.n272 VSUBS 0.017472f
C1163 VTAIL.n273 VSUBS 0.032515f
C1164 VTAIL.n274 VSUBS 0.032515f
C1165 VTAIL.n275 VSUBS 0.017472f
C1166 VTAIL.n276 VSUBS 0.0185f
C1167 VTAIL.n277 VSUBS 0.041298f
C1168 VTAIL.n278 VSUBS 0.041298f
C1169 VTAIL.n279 VSUBS 0.0185f
C1170 VTAIL.n280 VSUBS 0.017472f
C1171 VTAIL.n281 VSUBS 0.032515f
C1172 VTAIL.n282 VSUBS 0.081376f
C1173 VTAIL.n283 VSUBS 0.017472f
C1174 VTAIL.n284 VSUBS 0.0185f
C1175 VTAIL.n285 VSUBS 0.091064f
C1176 VTAIL.n286 VSUBS 0.059882f
C1177 VTAIL.n287 VSUBS 1.71052f
C1178 VP.n0 VSUBS 0.070738f
C1179 VP.t5 VSUBS 0.832132f
C1180 VP.t4 VSUBS 0.839433f
C1181 VP.t0 VSUBS 0.84913f
C1182 VP.n1 VSUBS 0.338876f
C1183 VP.t2 VSUBS 0.832132f
C1184 VP.n2 VSUBS 0.348817f
C1185 VP.t3 VSUBS 0.839433f
C1186 VP.n3 VSUBS 0.348058f
C1187 VP.n4 VSUBS 2.86186f
C1188 VP.n5 VSUBS 2.77775f
C1189 VP.n6 VSUBS 0.348058f
C1190 VP.n7 VSUBS 0.348817f
C1191 VP.t1 VSUBS 0.839433f
C1192 VP.n8 VSUBS 0.348058f
C1193 VP.n9 VSUBS 0.054819f
.ends

