* NGSPICE file created from diff_pair_sample_0306.ext - technology: sky130A

.subckt diff_pair_sample_0306 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=0 ps=0 w=18.4 l=2.42
X2 VTAIL.t6 VP.t0 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=3.036 ps=18.73 w=18.4 l=2.42
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=0 ps=0 w=18.4 l=2.42
X4 VDD1.t6 VP.t1 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X5 VDD1.t5 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X6 VDD2.t6 VN.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=0 ps=0 w=18.4 l=2.42
X8 VDD1.t4 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=7.176 ps=37.58 w=18.4 l=2.42
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=0 ps=0 w=18.4 l=2.42
X10 VDD2.t5 VN.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=7.176 ps=37.58 w=18.4 l=2.42
X11 VTAIL.t14 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=3.036 ps=18.73 w=18.4 l=2.42
X12 VTAIL.t12 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X13 VTAIL.t7 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=3.036 ps=18.73 w=18.4 l=2.42
X14 VTAIL.t2 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.176 pd=37.58 as=3.036 ps=18.73 w=18.4 l=2.42
X15 VDD1.t2 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=7.176 ps=37.58 w=18.4 l=2.42
X16 VTAIL.t11 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X17 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
X18 VDD2.t0 VN.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=7.176 ps=37.58 w=18.4 l=2.42
X19 VTAIL.t1 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.036 pd=18.73 as=3.036 ps=18.73 w=18.4 l=2.42
R0 VN.n6 VN.t5 215.745
R1 VN.n33 VN.t2 215.745
R2 VN.n7 VN.t0 183.24
R3 VN.n3 VN.t4 183.24
R4 VN.n25 VN.t7 183.24
R5 VN.n34 VN.t6 183.24
R6 VN.n30 VN.t1 183.24
R7 VN.n52 VN.t3 183.24
R8 VN.n51 VN.n27 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n28 161.3
R11 VN.n47 VN.n46 161.3
R12 VN.n45 VN.n29 161.3
R13 VN.n44 VN.n43 161.3
R14 VN.n42 VN.n41 161.3
R15 VN.n40 VN.n31 161.3
R16 VN.n39 VN.n38 161.3
R17 VN.n37 VN.n32 161.3
R18 VN.n36 VN.n35 161.3
R19 VN.n24 VN.n0 161.3
R20 VN.n23 VN.n22 161.3
R21 VN.n21 VN.n1 161.3
R22 VN.n20 VN.n19 161.3
R23 VN.n18 VN.n2 161.3
R24 VN.n17 VN.n16 161.3
R25 VN.n15 VN.n14 161.3
R26 VN.n13 VN.n4 161.3
R27 VN.n12 VN.n11 161.3
R28 VN.n10 VN.n5 161.3
R29 VN.n9 VN.n8 161.3
R30 VN.n26 VN.n25 104.76
R31 VN.n53 VN.n52 104.76
R32 VN.n19 VN.n1 56.5617
R33 VN.n46 VN.n28 56.5617
R34 VN VN.n53 55.0967
R35 VN.n7 VN.n6 53.9941
R36 VN.n34 VN.n33 53.9941
R37 VN.n12 VN.n5 40.577
R38 VN.n13 VN.n12 40.577
R39 VN.n39 VN.n32 40.577
R40 VN.n40 VN.n39 40.577
R41 VN.n8 VN.n5 24.5923
R42 VN.n14 VN.n13 24.5923
R43 VN.n18 VN.n17 24.5923
R44 VN.n19 VN.n18 24.5923
R45 VN.n23 VN.n1 24.5923
R46 VN.n24 VN.n23 24.5923
R47 VN.n35 VN.n32 24.5923
R48 VN.n46 VN.n45 24.5923
R49 VN.n45 VN.n44 24.5923
R50 VN.n41 VN.n40 24.5923
R51 VN.n51 VN.n50 24.5923
R52 VN.n50 VN.n28 24.5923
R53 VN.n8 VN.n7 18.4444
R54 VN.n14 VN.n3 18.4444
R55 VN.n35 VN.n34 18.4444
R56 VN.n41 VN.n30 18.4444
R57 VN.n36 VN.n33 7.07482
R58 VN.n9 VN.n6 7.07482
R59 VN.n17 VN.n3 6.14846
R60 VN.n25 VN.n24 6.14846
R61 VN.n44 VN.n30 6.14846
R62 VN.n52 VN.n51 6.14846
R63 VN.n53 VN.n27 0.278335
R64 VN.n26 VN.n0 0.278335
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n43 VN.n29 0.189894
R70 VN.n43 VN.n42 0.189894
R71 VN.n42 VN.n31 0.189894
R72 VN.n38 VN.n31 0.189894
R73 VN.n38 VN.n37 0.189894
R74 VN.n37 VN.n36 0.189894
R75 VN.n10 VN.n9 0.189894
R76 VN.n11 VN.n10 0.189894
R77 VN.n11 VN.n4 0.189894
R78 VN.n15 VN.n4 0.189894
R79 VN.n16 VN.n15 0.189894
R80 VN.n16 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153485
R86 VTAIL.n11 VTAIL.t6 47.6381
R87 VTAIL.n10 VTAIL.t13 47.6381
R88 VTAIL.n7 VTAIL.t14 47.6381
R89 VTAIL.n15 VTAIL.t8 47.6371
R90 VTAIL.n2 VTAIL.t7 47.6371
R91 VTAIL.n3 VTAIL.t0 47.6371
R92 VTAIL.n6 VTAIL.t2 47.6371
R93 VTAIL.n14 VTAIL.t5 47.6371
R94 VTAIL.n13 VTAIL.n12 46.562
R95 VTAIL.n9 VTAIL.n8 46.562
R96 VTAIL.n1 VTAIL.n0 46.5618
R97 VTAIL.n5 VTAIL.n4 46.5618
R98 VTAIL.n15 VTAIL.n14 30.5996
R99 VTAIL.n7 VTAIL.n6 30.5996
R100 VTAIL.n9 VTAIL.n7 2.37119
R101 VTAIL.n10 VTAIL.n9 2.37119
R102 VTAIL.n13 VTAIL.n11 2.37119
R103 VTAIL.n14 VTAIL.n13 2.37119
R104 VTAIL.n6 VTAIL.n5 2.37119
R105 VTAIL.n5 VTAIL.n3 2.37119
R106 VTAIL.n2 VTAIL.n1 2.37119
R107 VTAIL VTAIL.n15 2.313
R108 VTAIL.n0 VTAIL.t9 1.07659
R109 VTAIL.n0 VTAIL.t12 1.07659
R110 VTAIL.n4 VTAIL.t3 1.07659
R111 VTAIL.n4 VTAIL.t1 1.07659
R112 VTAIL.n12 VTAIL.t15 1.07659
R113 VTAIL.n12 VTAIL.t4 1.07659
R114 VTAIL.n8 VTAIL.t10 1.07659
R115 VTAIL.n8 VTAIL.t11 1.07659
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 VDD2.n2 VDD2.n1 64.3706
R120 VDD2.n2 VDD2.n0 64.3706
R121 VDD2 VDD2.n5 64.3669
R122 VDD2.n4 VDD2.n3 63.2408
R123 VDD2.n4 VDD2.n2 50.2455
R124 VDD2 VDD2.n4 1.24403
R125 VDD2.n5 VDD2.t1 1.07659
R126 VDD2.n5 VDD2.t5 1.07659
R127 VDD2.n3 VDD2.t4 1.07659
R128 VDD2.n3 VDD2.t6 1.07659
R129 VDD2.n1 VDD2.t3 1.07659
R130 VDD2.n1 VDD2.t0 1.07659
R131 VDD2.n0 VDD2.t2 1.07659
R132 VDD2.n0 VDD2.t7 1.07659
R133 B.n1049 B.n1048 585
R134 B.n416 B.n155 585
R135 B.n415 B.n414 585
R136 B.n413 B.n412 585
R137 B.n411 B.n410 585
R138 B.n409 B.n408 585
R139 B.n407 B.n406 585
R140 B.n405 B.n404 585
R141 B.n403 B.n402 585
R142 B.n401 B.n400 585
R143 B.n399 B.n398 585
R144 B.n397 B.n396 585
R145 B.n395 B.n394 585
R146 B.n393 B.n392 585
R147 B.n391 B.n390 585
R148 B.n389 B.n388 585
R149 B.n387 B.n386 585
R150 B.n385 B.n384 585
R151 B.n383 B.n382 585
R152 B.n381 B.n380 585
R153 B.n379 B.n378 585
R154 B.n377 B.n376 585
R155 B.n375 B.n374 585
R156 B.n373 B.n372 585
R157 B.n371 B.n370 585
R158 B.n369 B.n368 585
R159 B.n367 B.n366 585
R160 B.n365 B.n364 585
R161 B.n363 B.n362 585
R162 B.n361 B.n360 585
R163 B.n359 B.n358 585
R164 B.n357 B.n356 585
R165 B.n355 B.n354 585
R166 B.n353 B.n352 585
R167 B.n351 B.n350 585
R168 B.n349 B.n348 585
R169 B.n347 B.n346 585
R170 B.n345 B.n344 585
R171 B.n343 B.n342 585
R172 B.n341 B.n340 585
R173 B.n339 B.n338 585
R174 B.n337 B.n336 585
R175 B.n335 B.n334 585
R176 B.n333 B.n332 585
R177 B.n331 B.n330 585
R178 B.n329 B.n328 585
R179 B.n327 B.n326 585
R180 B.n325 B.n324 585
R181 B.n323 B.n322 585
R182 B.n321 B.n320 585
R183 B.n319 B.n318 585
R184 B.n317 B.n316 585
R185 B.n315 B.n314 585
R186 B.n313 B.n312 585
R187 B.n311 B.n310 585
R188 B.n309 B.n308 585
R189 B.n307 B.n306 585
R190 B.n305 B.n304 585
R191 B.n303 B.n302 585
R192 B.n301 B.n300 585
R193 B.n299 B.n298 585
R194 B.n297 B.n296 585
R195 B.n295 B.n294 585
R196 B.n293 B.n292 585
R197 B.n291 B.n290 585
R198 B.n289 B.n288 585
R199 B.n287 B.n286 585
R200 B.n285 B.n284 585
R201 B.n283 B.n282 585
R202 B.n281 B.n280 585
R203 B.n279 B.n278 585
R204 B.n277 B.n276 585
R205 B.n275 B.n274 585
R206 B.n273 B.n272 585
R207 B.n271 B.n270 585
R208 B.n269 B.n268 585
R209 B.n267 B.n266 585
R210 B.n265 B.n264 585
R211 B.n263 B.n262 585
R212 B.n261 B.n260 585
R213 B.n259 B.n258 585
R214 B.n257 B.n256 585
R215 B.n255 B.n254 585
R216 B.n253 B.n252 585
R217 B.n251 B.n250 585
R218 B.n249 B.n248 585
R219 B.n247 B.n246 585
R220 B.n245 B.n244 585
R221 B.n243 B.n242 585
R222 B.n241 B.n240 585
R223 B.n239 B.n238 585
R224 B.n237 B.n236 585
R225 B.n235 B.n234 585
R226 B.n233 B.n232 585
R227 B.n231 B.n230 585
R228 B.n229 B.n228 585
R229 B.n227 B.n226 585
R230 B.n225 B.n224 585
R231 B.n223 B.n222 585
R232 B.n221 B.n220 585
R233 B.n219 B.n218 585
R234 B.n217 B.n216 585
R235 B.n215 B.n214 585
R236 B.n213 B.n212 585
R237 B.n211 B.n210 585
R238 B.n209 B.n208 585
R239 B.n207 B.n206 585
R240 B.n205 B.n204 585
R241 B.n203 B.n202 585
R242 B.n201 B.n200 585
R243 B.n199 B.n198 585
R244 B.n197 B.n196 585
R245 B.n195 B.n194 585
R246 B.n193 B.n192 585
R247 B.n191 B.n190 585
R248 B.n189 B.n188 585
R249 B.n187 B.n186 585
R250 B.n185 B.n184 585
R251 B.n183 B.n182 585
R252 B.n181 B.n180 585
R253 B.n179 B.n178 585
R254 B.n177 B.n176 585
R255 B.n175 B.n174 585
R256 B.n173 B.n172 585
R257 B.n171 B.n170 585
R258 B.n169 B.n168 585
R259 B.n167 B.n166 585
R260 B.n165 B.n164 585
R261 B.n163 B.n162 585
R262 B.n89 B.n88 585
R263 B.n1047 B.n90 585
R264 B.n1052 B.n90 585
R265 B.n1046 B.n1045 585
R266 B.n1045 B.n86 585
R267 B.n1044 B.n85 585
R268 B.n1058 B.n85 585
R269 B.n1043 B.n84 585
R270 B.n1059 B.n84 585
R271 B.n1042 B.n83 585
R272 B.n1060 B.n83 585
R273 B.n1041 B.n1040 585
R274 B.n1040 B.n79 585
R275 B.n1039 B.n78 585
R276 B.n1066 B.n78 585
R277 B.n1038 B.n77 585
R278 B.n1067 B.n77 585
R279 B.n1037 B.n76 585
R280 B.n1068 B.n76 585
R281 B.n1036 B.n1035 585
R282 B.n1035 B.n72 585
R283 B.n1034 B.n71 585
R284 B.n1074 B.n71 585
R285 B.n1033 B.n70 585
R286 B.n1075 B.n70 585
R287 B.n1032 B.n69 585
R288 B.n1076 B.n69 585
R289 B.n1031 B.n1030 585
R290 B.n1030 B.n65 585
R291 B.n1029 B.n64 585
R292 B.n1082 B.n64 585
R293 B.n1028 B.n63 585
R294 B.n1083 B.n63 585
R295 B.n1027 B.n62 585
R296 B.n1084 B.n62 585
R297 B.n1026 B.n1025 585
R298 B.n1025 B.n58 585
R299 B.n1024 B.n57 585
R300 B.n1090 B.n57 585
R301 B.n1023 B.n56 585
R302 B.n1091 B.n56 585
R303 B.n1022 B.n55 585
R304 B.n1092 B.n55 585
R305 B.n1021 B.n1020 585
R306 B.n1020 B.n51 585
R307 B.n1019 B.n50 585
R308 B.n1098 B.n50 585
R309 B.n1018 B.n49 585
R310 B.n1099 B.n49 585
R311 B.n1017 B.n48 585
R312 B.n1100 B.n48 585
R313 B.n1016 B.n1015 585
R314 B.n1015 B.n44 585
R315 B.n1014 B.n43 585
R316 B.n1106 B.n43 585
R317 B.n1013 B.n42 585
R318 B.n1107 B.n42 585
R319 B.n1012 B.n41 585
R320 B.n1108 B.n41 585
R321 B.n1011 B.n1010 585
R322 B.n1010 B.n37 585
R323 B.n1009 B.n36 585
R324 B.n1114 B.n36 585
R325 B.n1008 B.n35 585
R326 B.n1115 B.n35 585
R327 B.n1007 B.n34 585
R328 B.n1116 B.n34 585
R329 B.n1006 B.n1005 585
R330 B.n1005 B.n30 585
R331 B.n1004 B.n29 585
R332 B.n1122 B.n29 585
R333 B.n1003 B.n28 585
R334 B.n1123 B.n28 585
R335 B.n1002 B.n27 585
R336 B.n1124 B.n27 585
R337 B.n1001 B.n1000 585
R338 B.n1000 B.n23 585
R339 B.n999 B.n22 585
R340 B.n1130 B.n22 585
R341 B.n998 B.n21 585
R342 B.n1131 B.n21 585
R343 B.n997 B.n20 585
R344 B.n1132 B.n20 585
R345 B.n996 B.n995 585
R346 B.n995 B.n16 585
R347 B.n994 B.n15 585
R348 B.n1138 B.n15 585
R349 B.n993 B.n14 585
R350 B.n1139 B.n14 585
R351 B.n992 B.n13 585
R352 B.n1140 B.n13 585
R353 B.n991 B.n990 585
R354 B.n990 B.n12 585
R355 B.n989 B.n988 585
R356 B.n989 B.n8 585
R357 B.n987 B.n7 585
R358 B.n1147 B.n7 585
R359 B.n986 B.n6 585
R360 B.n1148 B.n6 585
R361 B.n985 B.n5 585
R362 B.n1149 B.n5 585
R363 B.n984 B.n983 585
R364 B.n983 B.n4 585
R365 B.n982 B.n417 585
R366 B.n982 B.n981 585
R367 B.n972 B.n418 585
R368 B.n419 B.n418 585
R369 B.n974 B.n973 585
R370 B.n975 B.n974 585
R371 B.n971 B.n424 585
R372 B.n424 B.n423 585
R373 B.n970 B.n969 585
R374 B.n969 B.n968 585
R375 B.n426 B.n425 585
R376 B.n427 B.n426 585
R377 B.n961 B.n960 585
R378 B.n962 B.n961 585
R379 B.n959 B.n432 585
R380 B.n432 B.n431 585
R381 B.n958 B.n957 585
R382 B.n957 B.n956 585
R383 B.n434 B.n433 585
R384 B.n435 B.n434 585
R385 B.n949 B.n948 585
R386 B.n950 B.n949 585
R387 B.n947 B.n440 585
R388 B.n440 B.n439 585
R389 B.n946 B.n945 585
R390 B.n945 B.n944 585
R391 B.n442 B.n441 585
R392 B.n443 B.n442 585
R393 B.n937 B.n936 585
R394 B.n938 B.n937 585
R395 B.n935 B.n448 585
R396 B.n448 B.n447 585
R397 B.n934 B.n933 585
R398 B.n933 B.n932 585
R399 B.n450 B.n449 585
R400 B.n451 B.n450 585
R401 B.n925 B.n924 585
R402 B.n926 B.n925 585
R403 B.n923 B.n456 585
R404 B.n456 B.n455 585
R405 B.n922 B.n921 585
R406 B.n921 B.n920 585
R407 B.n458 B.n457 585
R408 B.n459 B.n458 585
R409 B.n913 B.n912 585
R410 B.n914 B.n913 585
R411 B.n911 B.n464 585
R412 B.n464 B.n463 585
R413 B.n910 B.n909 585
R414 B.n909 B.n908 585
R415 B.n466 B.n465 585
R416 B.n467 B.n466 585
R417 B.n901 B.n900 585
R418 B.n902 B.n901 585
R419 B.n899 B.n472 585
R420 B.n472 B.n471 585
R421 B.n898 B.n897 585
R422 B.n897 B.n896 585
R423 B.n474 B.n473 585
R424 B.n475 B.n474 585
R425 B.n889 B.n888 585
R426 B.n890 B.n889 585
R427 B.n887 B.n480 585
R428 B.n480 B.n479 585
R429 B.n886 B.n885 585
R430 B.n885 B.n884 585
R431 B.n482 B.n481 585
R432 B.n483 B.n482 585
R433 B.n877 B.n876 585
R434 B.n878 B.n877 585
R435 B.n875 B.n488 585
R436 B.n488 B.n487 585
R437 B.n874 B.n873 585
R438 B.n873 B.n872 585
R439 B.n490 B.n489 585
R440 B.n491 B.n490 585
R441 B.n865 B.n864 585
R442 B.n866 B.n865 585
R443 B.n863 B.n495 585
R444 B.n499 B.n495 585
R445 B.n862 B.n861 585
R446 B.n861 B.n860 585
R447 B.n497 B.n496 585
R448 B.n498 B.n497 585
R449 B.n853 B.n852 585
R450 B.n854 B.n853 585
R451 B.n851 B.n504 585
R452 B.n504 B.n503 585
R453 B.n850 B.n849 585
R454 B.n849 B.n848 585
R455 B.n506 B.n505 585
R456 B.n507 B.n506 585
R457 B.n841 B.n840 585
R458 B.n842 B.n841 585
R459 B.n510 B.n509 585
R460 B.n581 B.n579 585
R461 B.n582 B.n578 585
R462 B.n582 B.n511 585
R463 B.n585 B.n584 585
R464 B.n586 B.n577 585
R465 B.n588 B.n587 585
R466 B.n590 B.n576 585
R467 B.n593 B.n592 585
R468 B.n594 B.n575 585
R469 B.n596 B.n595 585
R470 B.n598 B.n574 585
R471 B.n601 B.n600 585
R472 B.n602 B.n573 585
R473 B.n604 B.n603 585
R474 B.n606 B.n572 585
R475 B.n609 B.n608 585
R476 B.n610 B.n571 585
R477 B.n612 B.n611 585
R478 B.n614 B.n570 585
R479 B.n617 B.n616 585
R480 B.n618 B.n569 585
R481 B.n620 B.n619 585
R482 B.n622 B.n568 585
R483 B.n625 B.n624 585
R484 B.n626 B.n567 585
R485 B.n628 B.n627 585
R486 B.n630 B.n566 585
R487 B.n633 B.n632 585
R488 B.n634 B.n565 585
R489 B.n636 B.n635 585
R490 B.n638 B.n564 585
R491 B.n641 B.n640 585
R492 B.n642 B.n563 585
R493 B.n644 B.n643 585
R494 B.n646 B.n562 585
R495 B.n649 B.n648 585
R496 B.n650 B.n561 585
R497 B.n652 B.n651 585
R498 B.n654 B.n560 585
R499 B.n657 B.n656 585
R500 B.n658 B.n559 585
R501 B.n660 B.n659 585
R502 B.n662 B.n558 585
R503 B.n665 B.n664 585
R504 B.n666 B.n557 585
R505 B.n668 B.n667 585
R506 B.n670 B.n556 585
R507 B.n673 B.n672 585
R508 B.n674 B.n555 585
R509 B.n676 B.n675 585
R510 B.n678 B.n554 585
R511 B.n681 B.n680 585
R512 B.n682 B.n553 585
R513 B.n684 B.n683 585
R514 B.n686 B.n552 585
R515 B.n689 B.n688 585
R516 B.n690 B.n551 585
R517 B.n692 B.n691 585
R518 B.n694 B.n550 585
R519 B.n697 B.n696 585
R520 B.n699 B.n547 585
R521 B.n701 B.n700 585
R522 B.n703 B.n546 585
R523 B.n706 B.n705 585
R524 B.n707 B.n545 585
R525 B.n709 B.n708 585
R526 B.n711 B.n544 585
R527 B.n714 B.n713 585
R528 B.n715 B.n543 585
R529 B.n720 B.n719 585
R530 B.n722 B.n542 585
R531 B.n725 B.n724 585
R532 B.n726 B.n541 585
R533 B.n728 B.n727 585
R534 B.n730 B.n540 585
R535 B.n733 B.n732 585
R536 B.n734 B.n539 585
R537 B.n736 B.n735 585
R538 B.n738 B.n538 585
R539 B.n741 B.n740 585
R540 B.n742 B.n537 585
R541 B.n744 B.n743 585
R542 B.n746 B.n536 585
R543 B.n749 B.n748 585
R544 B.n750 B.n535 585
R545 B.n752 B.n751 585
R546 B.n754 B.n534 585
R547 B.n757 B.n756 585
R548 B.n758 B.n533 585
R549 B.n760 B.n759 585
R550 B.n762 B.n532 585
R551 B.n765 B.n764 585
R552 B.n766 B.n531 585
R553 B.n768 B.n767 585
R554 B.n770 B.n530 585
R555 B.n773 B.n772 585
R556 B.n774 B.n529 585
R557 B.n776 B.n775 585
R558 B.n778 B.n528 585
R559 B.n781 B.n780 585
R560 B.n782 B.n527 585
R561 B.n784 B.n783 585
R562 B.n786 B.n526 585
R563 B.n789 B.n788 585
R564 B.n790 B.n525 585
R565 B.n792 B.n791 585
R566 B.n794 B.n524 585
R567 B.n797 B.n796 585
R568 B.n798 B.n523 585
R569 B.n800 B.n799 585
R570 B.n802 B.n522 585
R571 B.n805 B.n804 585
R572 B.n806 B.n521 585
R573 B.n808 B.n807 585
R574 B.n810 B.n520 585
R575 B.n813 B.n812 585
R576 B.n814 B.n519 585
R577 B.n816 B.n815 585
R578 B.n818 B.n518 585
R579 B.n821 B.n820 585
R580 B.n822 B.n517 585
R581 B.n824 B.n823 585
R582 B.n826 B.n516 585
R583 B.n829 B.n828 585
R584 B.n830 B.n515 585
R585 B.n832 B.n831 585
R586 B.n834 B.n514 585
R587 B.n835 B.n513 585
R588 B.n838 B.n837 585
R589 B.n839 B.n512 585
R590 B.n512 B.n511 585
R591 B.n844 B.n843 585
R592 B.n843 B.n842 585
R593 B.n845 B.n508 585
R594 B.n508 B.n507 585
R595 B.n847 B.n846 585
R596 B.n848 B.n847 585
R597 B.n502 B.n501 585
R598 B.n503 B.n502 585
R599 B.n856 B.n855 585
R600 B.n855 B.n854 585
R601 B.n857 B.n500 585
R602 B.n500 B.n498 585
R603 B.n859 B.n858 585
R604 B.n860 B.n859 585
R605 B.n494 B.n493 585
R606 B.n499 B.n494 585
R607 B.n868 B.n867 585
R608 B.n867 B.n866 585
R609 B.n869 B.n492 585
R610 B.n492 B.n491 585
R611 B.n871 B.n870 585
R612 B.n872 B.n871 585
R613 B.n486 B.n485 585
R614 B.n487 B.n486 585
R615 B.n880 B.n879 585
R616 B.n879 B.n878 585
R617 B.n881 B.n484 585
R618 B.n484 B.n483 585
R619 B.n883 B.n882 585
R620 B.n884 B.n883 585
R621 B.n478 B.n477 585
R622 B.n479 B.n478 585
R623 B.n892 B.n891 585
R624 B.n891 B.n890 585
R625 B.n893 B.n476 585
R626 B.n476 B.n475 585
R627 B.n895 B.n894 585
R628 B.n896 B.n895 585
R629 B.n470 B.n469 585
R630 B.n471 B.n470 585
R631 B.n904 B.n903 585
R632 B.n903 B.n902 585
R633 B.n905 B.n468 585
R634 B.n468 B.n467 585
R635 B.n907 B.n906 585
R636 B.n908 B.n907 585
R637 B.n462 B.n461 585
R638 B.n463 B.n462 585
R639 B.n916 B.n915 585
R640 B.n915 B.n914 585
R641 B.n917 B.n460 585
R642 B.n460 B.n459 585
R643 B.n919 B.n918 585
R644 B.n920 B.n919 585
R645 B.n454 B.n453 585
R646 B.n455 B.n454 585
R647 B.n928 B.n927 585
R648 B.n927 B.n926 585
R649 B.n929 B.n452 585
R650 B.n452 B.n451 585
R651 B.n931 B.n930 585
R652 B.n932 B.n931 585
R653 B.n446 B.n445 585
R654 B.n447 B.n446 585
R655 B.n940 B.n939 585
R656 B.n939 B.n938 585
R657 B.n941 B.n444 585
R658 B.n444 B.n443 585
R659 B.n943 B.n942 585
R660 B.n944 B.n943 585
R661 B.n438 B.n437 585
R662 B.n439 B.n438 585
R663 B.n952 B.n951 585
R664 B.n951 B.n950 585
R665 B.n953 B.n436 585
R666 B.n436 B.n435 585
R667 B.n955 B.n954 585
R668 B.n956 B.n955 585
R669 B.n430 B.n429 585
R670 B.n431 B.n430 585
R671 B.n964 B.n963 585
R672 B.n963 B.n962 585
R673 B.n965 B.n428 585
R674 B.n428 B.n427 585
R675 B.n967 B.n966 585
R676 B.n968 B.n967 585
R677 B.n422 B.n421 585
R678 B.n423 B.n422 585
R679 B.n977 B.n976 585
R680 B.n976 B.n975 585
R681 B.n978 B.n420 585
R682 B.n420 B.n419 585
R683 B.n980 B.n979 585
R684 B.n981 B.n980 585
R685 B.n3 B.n0 585
R686 B.n4 B.n3 585
R687 B.n1146 B.n1 585
R688 B.n1147 B.n1146 585
R689 B.n1145 B.n1144 585
R690 B.n1145 B.n8 585
R691 B.n1143 B.n9 585
R692 B.n12 B.n9 585
R693 B.n1142 B.n1141 585
R694 B.n1141 B.n1140 585
R695 B.n11 B.n10 585
R696 B.n1139 B.n11 585
R697 B.n1137 B.n1136 585
R698 B.n1138 B.n1137 585
R699 B.n1135 B.n17 585
R700 B.n17 B.n16 585
R701 B.n1134 B.n1133 585
R702 B.n1133 B.n1132 585
R703 B.n19 B.n18 585
R704 B.n1131 B.n19 585
R705 B.n1129 B.n1128 585
R706 B.n1130 B.n1129 585
R707 B.n1127 B.n24 585
R708 B.n24 B.n23 585
R709 B.n1126 B.n1125 585
R710 B.n1125 B.n1124 585
R711 B.n26 B.n25 585
R712 B.n1123 B.n26 585
R713 B.n1121 B.n1120 585
R714 B.n1122 B.n1121 585
R715 B.n1119 B.n31 585
R716 B.n31 B.n30 585
R717 B.n1118 B.n1117 585
R718 B.n1117 B.n1116 585
R719 B.n33 B.n32 585
R720 B.n1115 B.n33 585
R721 B.n1113 B.n1112 585
R722 B.n1114 B.n1113 585
R723 B.n1111 B.n38 585
R724 B.n38 B.n37 585
R725 B.n1110 B.n1109 585
R726 B.n1109 B.n1108 585
R727 B.n40 B.n39 585
R728 B.n1107 B.n40 585
R729 B.n1105 B.n1104 585
R730 B.n1106 B.n1105 585
R731 B.n1103 B.n45 585
R732 B.n45 B.n44 585
R733 B.n1102 B.n1101 585
R734 B.n1101 B.n1100 585
R735 B.n47 B.n46 585
R736 B.n1099 B.n47 585
R737 B.n1097 B.n1096 585
R738 B.n1098 B.n1097 585
R739 B.n1095 B.n52 585
R740 B.n52 B.n51 585
R741 B.n1094 B.n1093 585
R742 B.n1093 B.n1092 585
R743 B.n54 B.n53 585
R744 B.n1091 B.n54 585
R745 B.n1089 B.n1088 585
R746 B.n1090 B.n1089 585
R747 B.n1087 B.n59 585
R748 B.n59 B.n58 585
R749 B.n1086 B.n1085 585
R750 B.n1085 B.n1084 585
R751 B.n61 B.n60 585
R752 B.n1083 B.n61 585
R753 B.n1081 B.n1080 585
R754 B.n1082 B.n1081 585
R755 B.n1079 B.n66 585
R756 B.n66 B.n65 585
R757 B.n1078 B.n1077 585
R758 B.n1077 B.n1076 585
R759 B.n68 B.n67 585
R760 B.n1075 B.n68 585
R761 B.n1073 B.n1072 585
R762 B.n1074 B.n1073 585
R763 B.n1071 B.n73 585
R764 B.n73 B.n72 585
R765 B.n1070 B.n1069 585
R766 B.n1069 B.n1068 585
R767 B.n75 B.n74 585
R768 B.n1067 B.n75 585
R769 B.n1065 B.n1064 585
R770 B.n1066 B.n1065 585
R771 B.n1063 B.n80 585
R772 B.n80 B.n79 585
R773 B.n1062 B.n1061 585
R774 B.n1061 B.n1060 585
R775 B.n82 B.n81 585
R776 B.n1059 B.n82 585
R777 B.n1057 B.n1056 585
R778 B.n1058 B.n1057 585
R779 B.n1055 B.n87 585
R780 B.n87 B.n86 585
R781 B.n1054 B.n1053 585
R782 B.n1053 B.n1052 585
R783 B.n1150 B.n1149 585
R784 B.n1148 B.n2 585
R785 B.n1053 B.n89 545.355
R786 B.n1049 B.n90 545.355
R787 B.n841 B.n512 545.355
R788 B.n843 B.n510 545.355
R789 B.n159 B.t8 390.998
R790 B.n156 B.t16 390.998
R791 B.n716 B.t19 390.998
R792 B.n548 B.t12 390.998
R793 B.n1051 B.n1050 256.663
R794 B.n1051 B.n154 256.663
R795 B.n1051 B.n153 256.663
R796 B.n1051 B.n152 256.663
R797 B.n1051 B.n151 256.663
R798 B.n1051 B.n150 256.663
R799 B.n1051 B.n149 256.663
R800 B.n1051 B.n148 256.663
R801 B.n1051 B.n147 256.663
R802 B.n1051 B.n146 256.663
R803 B.n1051 B.n145 256.663
R804 B.n1051 B.n144 256.663
R805 B.n1051 B.n143 256.663
R806 B.n1051 B.n142 256.663
R807 B.n1051 B.n141 256.663
R808 B.n1051 B.n140 256.663
R809 B.n1051 B.n139 256.663
R810 B.n1051 B.n138 256.663
R811 B.n1051 B.n137 256.663
R812 B.n1051 B.n136 256.663
R813 B.n1051 B.n135 256.663
R814 B.n1051 B.n134 256.663
R815 B.n1051 B.n133 256.663
R816 B.n1051 B.n132 256.663
R817 B.n1051 B.n131 256.663
R818 B.n1051 B.n130 256.663
R819 B.n1051 B.n129 256.663
R820 B.n1051 B.n128 256.663
R821 B.n1051 B.n127 256.663
R822 B.n1051 B.n126 256.663
R823 B.n1051 B.n125 256.663
R824 B.n1051 B.n124 256.663
R825 B.n1051 B.n123 256.663
R826 B.n1051 B.n122 256.663
R827 B.n1051 B.n121 256.663
R828 B.n1051 B.n120 256.663
R829 B.n1051 B.n119 256.663
R830 B.n1051 B.n118 256.663
R831 B.n1051 B.n117 256.663
R832 B.n1051 B.n116 256.663
R833 B.n1051 B.n115 256.663
R834 B.n1051 B.n114 256.663
R835 B.n1051 B.n113 256.663
R836 B.n1051 B.n112 256.663
R837 B.n1051 B.n111 256.663
R838 B.n1051 B.n110 256.663
R839 B.n1051 B.n109 256.663
R840 B.n1051 B.n108 256.663
R841 B.n1051 B.n107 256.663
R842 B.n1051 B.n106 256.663
R843 B.n1051 B.n105 256.663
R844 B.n1051 B.n104 256.663
R845 B.n1051 B.n103 256.663
R846 B.n1051 B.n102 256.663
R847 B.n1051 B.n101 256.663
R848 B.n1051 B.n100 256.663
R849 B.n1051 B.n99 256.663
R850 B.n1051 B.n98 256.663
R851 B.n1051 B.n97 256.663
R852 B.n1051 B.n96 256.663
R853 B.n1051 B.n95 256.663
R854 B.n1051 B.n94 256.663
R855 B.n1051 B.n93 256.663
R856 B.n1051 B.n92 256.663
R857 B.n1051 B.n91 256.663
R858 B.n580 B.n511 256.663
R859 B.n583 B.n511 256.663
R860 B.n589 B.n511 256.663
R861 B.n591 B.n511 256.663
R862 B.n597 B.n511 256.663
R863 B.n599 B.n511 256.663
R864 B.n605 B.n511 256.663
R865 B.n607 B.n511 256.663
R866 B.n613 B.n511 256.663
R867 B.n615 B.n511 256.663
R868 B.n621 B.n511 256.663
R869 B.n623 B.n511 256.663
R870 B.n629 B.n511 256.663
R871 B.n631 B.n511 256.663
R872 B.n637 B.n511 256.663
R873 B.n639 B.n511 256.663
R874 B.n645 B.n511 256.663
R875 B.n647 B.n511 256.663
R876 B.n653 B.n511 256.663
R877 B.n655 B.n511 256.663
R878 B.n661 B.n511 256.663
R879 B.n663 B.n511 256.663
R880 B.n669 B.n511 256.663
R881 B.n671 B.n511 256.663
R882 B.n677 B.n511 256.663
R883 B.n679 B.n511 256.663
R884 B.n685 B.n511 256.663
R885 B.n687 B.n511 256.663
R886 B.n693 B.n511 256.663
R887 B.n695 B.n511 256.663
R888 B.n702 B.n511 256.663
R889 B.n704 B.n511 256.663
R890 B.n710 B.n511 256.663
R891 B.n712 B.n511 256.663
R892 B.n721 B.n511 256.663
R893 B.n723 B.n511 256.663
R894 B.n729 B.n511 256.663
R895 B.n731 B.n511 256.663
R896 B.n737 B.n511 256.663
R897 B.n739 B.n511 256.663
R898 B.n745 B.n511 256.663
R899 B.n747 B.n511 256.663
R900 B.n753 B.n511 256.663
R901 B.n755 B.n511 256.663
R902 B.n761 B.n511 256.663
R903 B.n763 B.n511 256.663
R904 B.n769 B.n511 256.663
R905 B.n771 B.n511 256.663
R906 B.n777 B.n511 256.663
R907 B.n779 B.n511 256.663
R908 B.n785 B.n511 256.663
R909 B.n787 B.n511 256.663
R910 B.n793 B.n511 256.663
R911 B.n795 B.n511 256.663
R912 B.n801 B.n511 256.663
R913 B.n803 B.n511 256.663
R914 B.n809 B.n511 256.663
R915 B.n811 B.n511 256.663
R916 B.n817 B.n511 256.663
R917 B.n819 B.n511 256.663
R918 B.n825 B.n511 256.663
R919 B.n827 B.n511 256.663
R920 B.n833 B.n511 256.663
R921 B.n836 B.n511 256.663
R922 B.n1152 B.n1151 256.663
R923 B.n164 B.n163 163.367
R924 B.n168 B.n167 163.367
R925 B.n172 B.n171 163.367
R926 B.n176 B.n175 163.367
R927 B.n180 B.n179 163.367
R928 B.n184 B.n183 163.367
R929 B.n188 B.n187 163.367
R930 B.n192 B.n191 163.367
R931 B.n196 B.n195 163.367
R932 B.n200 B.n199 163.367
R933 B.n204 B.n203 163.367
R934 B.n208 B.n207 163.367
R935 B.n212 B.n211 163.367
R936 B.n216 B.n215 163.367
R937 B.n220 B.n219 163.367
R938 B.n224 B.n223 163.367
R939 B.n228 B.n227 163.367
R940 B.n232 B.n231 163.367
R941 B.n236 B.n235 163.367
R942 B.n240 B.n239 163.367
R943 B.n244 B.n243 163.367
R944 B.n248 B.n247 163.367
R945 B.n252 B.n251 163.367
R946 B.n256 B.n255 163.367
R947 B.n260 B.n259 163.367
R948 B.n264 B.n263 163.367
R949 B.n268 B.n267 163.367
R950 B.n272 B.n271 163.367
R951 B.n276 B.n275 163.367
R952 B.n280 B.n279 163.367
R953 B.n284 B.n283 163.367
R954 B.n288 B.n287 163.367
R955 B.n292 B.n291 163.367
R956 B.n296 B.n295 163.367
R957 B.n300 B.n299 163.367
R958 B.n304 B.n303 163.367
R959 B.n308 B.n307 163.367
R960 B.n312 B.n311 163.367
R961 B.n316 B.n315 163.367
R962 B.n320 B.n319 163.367
R963 B.n324 B.n323 163.367
R964 B.n328 B.n327 163.367
R965 B.n332 B.n331 163.367
R966 B.n336 B.n335 163.367
R967 B.n340 B.n339 163.367
R968 B.n344 B.n343 163.367
R969 B.n348 B.n347 163.367
R970 B.n352 B.n351 163.367
R971 B.n356 B.n355 163.367
R972 B.n360 B.n359 163.367
R973 B.n364 B.n363 163.367
R974 B.n368 B.n367 163.367
R975 B.n372 B.n371 163.367
R976 B.n376 B.n375 163.367
R977 B.n380 B.n379 163.367
R978 B.n384 B.n383 163.367
R979 B.n388 B.n387 163.367
R980 B.n392 B.n391 163.367
R981 B.n396 B.n395 163.367
R982 B.n400 B.n399 163.367
R983 B.n404 B.n403 163.367
R984 B.n408 B.n407 163.367
R985 B.n412 B.n411 163.367
R986 B.n414 B.n155 163.367
R987 B.n841 B.n506 163.367
R988 B.n849 B.n506 163.367
R989 B.n849 B.n504 163.367
R990 B.n853 B.n504 163.367
R991 B.n853 B.n497 163.367
R992 B.n861 B.n497 163.367
R993 B.n861 B.n495 163.367
R994 B.n865 B.n495 163.367
R995 B.n865 B.n490 163.367
R996 B.n873 B.n490 163.367
R997 B.n873 B.n488 163.367
R998 B.n877 B.n488 163.367
R999 B.n877 B.n482 163.367
R1000 B.n885 B.n482 163.367
R1001 B.n885 B.n480 163.367
R1002 B.n889 B.n480 163.367
R1003 B.n889 B.n474 163.367
R1004 B.n897 B.n474 163.367
R1005 B.n897 B.n472 163.367
R1006 B.n901 B.n472 163.367
R1007 B.n901 B.n466 163.367
R1008 B.n909 B.n466 163.367
R1009 B.n909 B.n464 163.367
R1010 B.n913 B.n464 163.367
R1011 B.n913 B.n458 163.367
R1012 B.n921 B.n458 163.367
R1013 B.n921 B.n456 163.367
R1014 B.n925 B.n456 163.367
R1015 B.n925 B.n450 163.367
R1016 B.n933 B.n450 163.367
R1017 B.n933 B.n448 163.367
R1018 B.n937 B.n448 163.367
R1019 B.n937 B.n442 163.367
R1020 B.n945 B.n442 163.367
R1021 B.n945 B.n440 163.367
R1022 B.n949 B.n440 163.367
R1023 B.n949 B.n434 163.367
R1024 B.n957 B.n434 163.367
R1025 B.n957 B.n432 163.367
R1026 B.n961 B.n432 163.367
R1027 B.n961 B.n426 163.367
R1028 B.n969 B.n426 163.367
R1029 B.n969 B.n424 163.367
R1030 B.n974 B.n424 163.367
R1031 B.n974 B.n418 163.367
R1032 B.n982 B.n418 163.367
R1033 B.n983 B.n982 163.367
R1034 B.n983 B.n5 163.367
R1035 B.n6 B.n5 163.367
R1036 B.n7 B.n6 163.367
R1037 B.n989 B.n7 163.367
R1038 B.n990 B.n989 163.367
R1039 B.n990 B.n13 163.367
R1040 B.n14 B.n13 163.367
R1041 B.n15 B.n14 163.367
R1042 B.n995 B.n15 163.367
R1043 B.n995 B.n20 163.367
R1044 B.n21 B.n20 163.367
R1045 B.n22 B.n21 163.367
R1046 B.n1000 B.n22 163.367
R1047 B.n1000 B.n27 163.367
R1048 B.n28 B.n27 163.367
R1049 B.n29 B.n28 163.367
R1050 B.n1005 B.n29 163.367
R1051 B.n1005 B.n34 163.367
R1052 B.n35 B.n34 163.367
R1053 B.n36 B.n35 163.367
R1054 B.n1010 B.n36 163.367
R1055 B.n1010 B.n41 163.367
R1056 B.n42 B.n41 163.367
R1057 B.n43 B.n42 163.367
R1058 B.n1015 B.n43 163.367
R1059 B.n1015 B.n48 163.367
R1060 B.n49 B.n48 163.367
R1061 B.n50 B.n49 163.367
R1062 B.n1020 B.n50 163.367
R1063 B.n1020 B.n55 163.367
R1064 B.n56 B.n55 163.367
R1065 B.n57 B.n56 163.367
R1066 B.n1025 B.n57 163.367
R1067 B.n1025 B.n62 163.367
R1068 B.n63 B.n62 163.367
R1069 B.n64 B.n63 163.367
R1070 B.n1030 B.n64 163.367
R1071 B.n1030 B.n69 163.367
R1072 B.n70 B.n69 163.367
R1073 B.n71 B.n70 163.367
R1074 B.n1035 B.n71 163.367
R1075 B.n1035 B.n76 163.367
R1076 B.n77 B.n76 163.367
R1077 B.n78 B.n77 163.367
R1078 B.n1040 B.n78 163.367
R1079 B.n1040 B.n83 163.367
R1080 B.n84 B.n83 163.367
R1081 B.n85 B.n84 163.367
R1082 B.n1045 B.n85 163.367
R1083 B.n1045 B.n90 163.367
R1084 B.n582 B.n581 163.367
R1085 B.n584 B.n582 163.367
R1086 B.n588 B.n577 163.367
R1087 B.n592 B.n590 163.367
R1088 B.n596 B.n575 163.367
R1089 B.n600 B.n598 163.367
R1090 B.n604 B.n573 163.367
R1091 B.n608 B.n606 163.367
R1092 B.n612 B.n571 163.367
R1093 B.n616 B.n614 163.367
R1094 B.n620 B.n569 163.367
R1095 B.n624 B.n622 163.367
R1096 B.n628 B.n567 163.367
R1097 B.n632 B.n630 163.367
R1098 B.n636 B.n565 163.367
R1099 B.n640 B.n638 163.367
R1100 B.n644 B.n563 163.367
R1101 B.n648 B.n646 163.367
R1102 B.n652 B.n561 163.367
R1103 B.n656 B.n654 163.367
R1104 B.n660 B.n559 163.367
R1105 B.n664 B.n662 163.367
R1106 B.n668 B.n557 163.367
R1107 B.n672 B.n670 163.367
R1108 B.n676 B.n555 163.367
R1109 B.n680 B.n678 163.367
R1110 B.n684 B.n553 163.367
R1111 B.n688 B.n686 163.367
R1112 B.n692 B.n551 163.367
R1113 B.n696 B.n694 163.367
R1114 B.n701 B.n547 163.367
R1115 B.n705 B.n703 163.367
R1116 B.n709 B.n545 163.367
R1117 B.n713 B.n711 163.367
R1118 B.n720 B.n543 163.367
R1119 B.n724 B.n722 163.367
R1120 B.n728 B.n541 163.367
R1121 B.n732 B.n730 163.367
R1122 B.n736 B.n539 163.367
R1123 B.n740 B.n738 163.367
R1124 B.n744 B.n537 163.367
R1125 B.n748 B.n746 163.367
R1126 B.n752 B.n535 163.367
R1127 B.n756 B.n754 163.367
R1128 B.n760 B.n533 163.367
R1129 B.n764 B.n762 163.367
R1130 B.n768 B.n531 163.367
R1131 B.n772 B.n770 163.367
R1132 B.n776 B.n529 163.367
R1133 B.n780 B.n778 163.367
R1134 B.n784 B.n527 163.367
R1135 B.n788 B.n786 163.367
R1136 B.n792 B.n525 163.367
R1137 B.n796 B.n794 163.367
R1138 B.n800 B.n523 163.367
R1139 B.n804 B.n802 163.367
R1140 B.n808 B.n521 163.367
R1141 B.n812 B.n810 163.367
R1142 B.n816 B.n519 163.367
R1143 B.n820 B.n818 163.367
R1144 B.n824 B.n517 163.367
R1145 B.n828 B.n826 163.367
R1146 B.n832 B.n515 163.367
R1147 B.n835 B.n834 163.367
R1148 B.n837 B.n512 163.367
R1149 B.n843 B.n508 163.367
R1150 B.n847 B.n508 163.367
R1151 B.n847 B.n502 163.367
R1152 B.n855 B.n502 163.367
R1153 B.n855 B.n500 163.367
R1154 B.n859 B.n500 163.367
R1155 B.n859 B.n494 163.367
R1156 B.n867 B.n494 163.367
R1157 B.n867 B.n492 163.367
R1158 B.n871 B.n492 163.367
R1159 B.n871 B.n486 163.367
R1160 B.n879 B.n486 163.367
R1161 B.n879 B.n484 163.367
R1162 B.n883 B.n484 163.367
R1163 B.n883 B.n478 163.367
R1164 B.n891 B.n478 163.367
R1165 B.n891 B.n476 163.367
R1166 B.n895 B.n476 163.367
R1167 B.n895 B.n470 163.367
R1168 B.n903 B.n470 163.367
R1169 B.n903 B.n468 163.367
R1170 B.n907 B.n468 163.367
R1171 B.n907 B.n462 163.367
R1172 B.n915 B.n462 163.367
R1173 B.n915 B.n460 163.367
R1174 B.n919 B.n460 163.367
R1175 B.n919 B.n454 163.367
R1176 B.n927 B.n454 163.367
R1177 B.n927 B.n452 163.367
R1178 B.n931 B.n452 163.367
R1179 B.n931 B.n446 163.367
R1180 B.n939 B.n446 163.367
R1181 B.n939 B.n444 163.367
R1182 B.n943 B.n444 163.367
R1183 B.n943 B.n438 163.367
R1184 B.n951 B.n438 163.367
R1185 B.n951 B.n436 163.367
R1186 B.n955 B.n436 163.367
R1187 B.n955 B.n430 163.367
R1188 B.n963 B.n430 163.367
R1189 B.n963 B.n428 163.367
R1190 B.n967 B.n428 163.367
R1191 B.n967 B.n422 163.367
R1192 B.n976 B.n422 163.367
R1193 B.n976 B.n420 163.367
R1194 B.n980 B.n420 163.367
R1195 B.n980 B.n3 163.367
R1196 B.n1150 B.n3 163.367
R1197 B.n1146 B.n2 163.367
R1198 B.n1146 B.n1145 163.367
R1199 B.n1145 B.n9 163.367
R1200 B.n1141 B.n9 163.367
R1201 B.n1141 B.n11 163.367
R1202 B.n1137 B.n11 163.367
R1203 B.n1137 B.n17 163.367
R1204 B.n1133 B.n17 163.367
R1205 B.n1133 B.n19 163.367
R1206 B.n1129 B.n19 163.367
R1207 B.n1129 B.n24 163.367
R1208 B.n1125 B.n24 163.367
R1209 B.n1125 B.n26 163.367
R1210 B.n1121 B.n26 163.367
R1211 B.n1121 B.n31 163.367
R1212 B.n1117 B.n31 163.367
R1213 B.n1117 B.n33 163.367
R1214 B.n1113 B.n33 163.367
R1215 B.n1113 B.n38 163.367
R1216 B.n1109 B.n38 163.367
R1217 B.n1109 B.n40 163.367
R1218 B.n1105 B.n40 163.367
R1219 B.n1105 B.n45 163.367
R1220 B.n1101 B.n45 163.367
R1221 B.n1101 B.n47 163.367
R1222 B.n1097 B.n47 163.367
R1223 B.n1097 B.n52 163.367
R1224 B.n1093 B.n52 163.367
R1225 B.n1093 B.n54 163.367
R1226 B.n1089 B.n54 163.367
R1227 B.n1089 B.n59 163.367
R1228 B.n1085 B.n59 163.367
R1229 B.n1085 B.n61 163.367
R1230 B.n1081 B.n61 163.367
R1231 B.n1081 B.n66 163.367
R1232 B.n1077 B.n66 163.367
R1233 B.n1077 B.n68 163.367
R1234 B.n1073 B.n68 163.367
R1235 B.n1073 B.n73 163.367
R1236 B.n1069 B.n73 163.367
R1237 B.n1069 B.n75 163.367
R1238 B.n1065 B.n75 163.367
R1239 B.n1065 B.n80 163.367
R1240 B.n1061 B.n80 163.367
R1241 B.n1061 B.n82 163.367
R1242 B.n1057 B.n82 163.367
R1243 B.n1057 B.n87 163.367
R1244 B.n1053 B.n87 163.367
R1245 B.n156 B.t17 121.335
R1246 B.n716 B.t21 121.335
R1247 B.n159 B.t10 121.309
R1248 B.n548 B.t15 121.309
R1249 B.n91 B.n89 71.676
R1250 B.n164 B.n92 71.676
R1251 B.n168 B.n93 71.676
R1252 B.n172 B.n94 71.676
R1253 B.n176 B.n95 71.676
R1254 B.n180 B.n96 71.676
R1255 B.n184 B.n97 71.676
R1256 B.n188 B.n98 71.676
R1257 B.n192 B.n99 71.676
R1258 B.n196 B.n100 71.676
R1259 B.n200 B.n101 71.676
R1260 B.n204 B.n102 71.676
R1261 B.n208 B.n103 71.676
R1262 B.n212 B.n104 71.676
R1263 B.n216 B.n105 71.676
R1264 B.n220 B.n106 71.676
R1265 B.n224 B.n107 71.676
R1266 B.n228 B.n108 71.676
R1267 B.n232 B.n109 71.676
R1268 B.n236 B.n110 71.676
R1269 B.n240 B.n111 71.676
R1270 B.n244 B.n112 71.676
R1271 B.n248 B.n113 71.676
R1272 B.n252 B.n114 71.676
R1273 B.n256 B.n115 71.676
R1274 B.n260 B.n116 71.676
R1275 B.n264 B.n117 71.676
R1276 B.n268 B.n118 71.676
R1277 B.n272 B.n119 71.676
R1278 B.n276 B.n120 71.676
R1279 B.n280 B.n121 71.676
R1280 B.n284 B.n122 71.676
R1281 B.n288 B.n123 71.676
R1282 B.n292 B.n124 71.676
R1283 B.n296 B.n125 71.676
R1284 B.n300 B.n126 71.676
R1285 B.n304 B.n127 71.676
R1286 B.n308 B.n128 71.676
R1287 B.n312 B.n129 71.676
R1288 B.n316 B.n130 71.676
R1289 B.n320 B.n131 71.676
R1290 B.n324 B.n132 71.676
R1291 B.n328 B.n133 71.676
R1292 B.n332 B.n134 71.676
R1293 B.n336 B.n135 71.676
R1294 B.n340 B.n136 71.676
R1295 B.n344 B.n137 71.676
R1296 B.n348 B.n138 71.676
R1297 B.n352 B.n139 71.676
R1298 B.n356 B.n140 71.676
R1299 B.n360 B.n141 71.676
R1300 B.n364 B.n142 71.676
R1301 B.n368 B.n143 71.676
R1302 B.n372 B.n144 71.676
R1303 B.n376 B.n145 71.676
R1304 B.n380 B.n146 71.676
R1305 B.n384 B.n147 71.676
R1306 B.n388 B.n148 71.676
R1307 B.n392 B.n149 71.676
R1308 B.n396 B.n150 71.676
R1309 B.n400 B.n151 71.676
R1310 B.n404 B.n152 71.676
R1311 B.n408 B.n153 71.676
R1312 B.n412 B.n154 71.676
R1313 B.n1050 B.n155 71.676
R1314 B.n1050 B.n1049 71.676
R1315 B.n414 B.n154 71.676
R1316 B.n411 B.n153 71.676
R1317 B.n407 B.n152 71.676
R1318 B.n403 B.n151 71.676
R1319 B.n399 B.n150 71.676
R1320 B.n395 B.n149 71.676
R1321 B.n391 B.n148 71.676
R1322 B.n387 B.n147 71.676
R1323 B.n383 B.n146 71.676
R1324 B.n379 B.n145 71.676
R1325 B.n375 B.n144 71.676
R1326 B.n371 B.n143 71.676
R1327 B.n367 B.n142 71.676
R1328 B.n363 B.n141 71.676
R1329 B.n359 B.n140 71.676
R1330 B.n355 B.n139 71.676
R1331 B.n351 B.n138 71.676
R1332 B.n347 B.n137 71.676
R1333 B.n343 B.n136 71.676
R1334 B.n339 B.n135 71.676
R1335 B.n335 B.n134 71.676
R1336 B.n331 B.n133 71.676
R1337 B.n327 B.n132 71.676
R1338 B.n323 B.n131 71.676
R1339 B.n319 B.n130 71.676
R1340 B.n315 B.n129 71.676
R1341 B.n311 B.n128 71.676
R1342 B.n307 B.n127 71.676
R1343 B.n303 B.n126 71.676
R1344 B.n299 B.n125 71.676
R1345 B.n295 B.n124 71.676
R1346 B.n291 B.n123 71.676
R1347 B.n287 B.n122 71.676
R1348 B.n283 B.n121 71.676
R1349 B.n279 B.n120 71.676
R1350 B.n275 B.n119 71.676
R1351 B.n271 B.n118 71.676
R1352 B.n267 B.n117 71.676
R1353 B.n263 B.n116 71.676
R1354 B.n259 B.n115 71.676
R1355 B.n255 B.n114 71.676
R1356 B.n251 B.n113 71.676
R1357 B.n247 B.n112 71.676
R1358 B.n243 B.n111 71.676
R1359 B.n239 B.n110 71.676
R1360 B.n235 B.n109 71.676
R1361 B.n231 B.n108 71.676
R1362 B.n227 B.n107 71.676
R1363 B.n223 B.n106 71.676
R1364 B.n219 B.n105 71.676
R1365 B.n215 B.n104 71.676
R1366 B.n211 B.n103 71.676
R1367 B.n207 B.n102 71.676
R1368 B.n203 B.n101 71.676
R1369 B.n199 B.n100 71.676
R1370 B.n195 B.n99 71.676
R1371 B.n191 B.n98 71.676
R1372 B.n187 B.n97 71.676
R1373 B.n183 B.n96 71.676
R1374 B.n179 B.n95 71.676
R1375 B.n175 B.n94 71.676
R1376 B.n171 B.n93 71.676
R1377 B.n167 B.n92 71.676
R1378 B.n163 B.n91 71.676
R1379 B.n580 B.n510 71.676
R1380 B.n584 B.n583 71.676
R1381 B.n589 B.n588 71.676
R1382 B.n592 B.n591 71.676
R1383 B.n597 B.n596 71.676
R1384 B.n600 B.n599 71.676
R1385 B.n605 B.n604 71.676
R1386 B.n608 B.n607 71.676
R1387 B.n613 B.n612 71.676
R1388 B.n616 B.n615 71.676
R1389 B.n621 B.n620 71.676
R1390 B.n624 B.n623 71.676
R1391 B.n629 B.n628 71.676
R1392 B.n632 B.n631 71.676
R1393 B.n637 B.n636 71.676
R1394 B.n640 B.n639 71.676
R1395 B.n645 B.n644 71.676
R1396 B.n648 B.n647 71.676
R1397 B.n653 B.n652 71.676
R1398 B.n656 B.n655 71.676
R1399 B.n661 B.n660 71.676
R1400 B.n664 B.n663 71.676
R1401 B.n669 B.n668 71.676
R1402 B.n672 B.n671 71.676
R1403 B.n677 B.n676 71.676
R1404 B.n680 B.n679 71.676
R1405 B.n685 B.n684 71.676
R1406 B.n688 B.n687 71.676
R1407 B.n693 B.n692 71.676
R1408 B.n696 B.n695 71.676
R1409 B.n702 B.n701 71.676
R1410 B.n705 B.n704 71.676
R1411 B.n710 B.n709 71.676
R1412 B.n713 B.n712 71.676
R1413 B.n721 B.n720 71.676
R1414 B.n724 B.n723 71.676
R1415 B.n729 B.n728 71.676
R1416 B.n732 B.n731 71.676
R1417 B.n737 B.n736 71.676
R1418 B.n740 B.n739 71.676
R1419 B.n745 B.n744 71.676
R1420 B.n748 B.n747 71.676
R1421 B.n753 B.n752 71.676
R1422 B.n756 B.n755 71.676
R1423 B.n761 B.n760 71.676
R1424 B.n764 B.n763 71.676
R1425 B.n769 B.n768 71.676
R1426 B.n772 B.n771 71.676
R1427 B.n777 B.n776 71.676
R1428 B.n780 B.n779 71.676
R1429 B.n785 B.n784 71.676
R1430 B.n788 B.n787 71.676
R1431 B.n793 B.n792 71.676
R1432 B.n796 B.n795 71.676
R1433 B.n801 B.n800 71.676
R1434 B.n804 B.n803 71.676
R1435 B.n809 B.n808 71.676
R1436 B.n812 B.n811 71.676
R1437 B.n817 B.n816 71.676
R1438 B.n820 B.n819 71.676
R1439 B.n825 B.n824 71.676
R1440 B.n828 B.n827 71.676
R1441 B.n833 B.n832 71.676
R1442 B.n836 B.n835 71.676
R1443 B.n581 B.n580 71.676
R1444 B.n583 B.n577 71.676
R1445 B.n590 B.n589 71.676
R1446 B.n591 B.n575 71.676
R1447 B.n598 B.n597 71.676
R1448 B.n599 B.n573 71.676
R1449 B.n606 B.n605 71.676
R1450 B.n607 B.n571 71.676
R1451 B.n614 B.n613 71.676
R1452 B.n615 B.n569 71.676
R1453 B.n622 B.n621 71.676
R1454 B.n623 B.n567 71.676
R1455 B.n630 B.n629 71.676
R1456 B.n631 B.n565 71.676
R1457 B.n638 B.n637 71.676
R1458 B.n639 B.n563 71.676
R1459 B.n646 B.n645 71.676
R1460 B.n647 B.n561 71.676
R1461 B.n654 B.n653 71.676
R1462 B.n655 B.n559 71.676
R1463 B.n662 B.n661 71.676
R1464 B.n663 B.n557 71.676
R1465 B.n670 B.n669 71.676
R1466 B.n671 B.n555 71.676
R1467 B.n678 B.n677 71.676
R1468 B.n679 B.n553 71.676
R1469 B.n686 B.n685 71.676
R1470 B.n687 B.n551 71.676
R1471 B.n694 B.n693 71.676
R1472 B.n695 B.n547 71.676
R1473 B.n703 B.n702 71.676
R1474 B.n704 B.n545 71.676
R1475 B.n711 B.n710 71.676
R1476 B.n712 B.n543 71.676
R1477 B.n722 B.n721 71.676
R1478 B.n723 B.n541 71.676
R1479 B.n730 B.n729 71.676
R1480 B.n731 B.n539 71.676
R1481 B.n738 B.n737 71.676
R1482 B.n739 B.n537 71.676
R1483 B.n746 B.n745 71.676
R1484 B.n747 B.n535 71.676
R1485 B.n754 B.n753 71.676
R1486 B.n755 B.n533 71.676
R1487 B.n762 B.n761 71.676
R1488 B.n763 B.n531 71.676
R1489 B.n770 B.n769 71.676
R1490 B.n771 B.n529 71.676
R1491 B.n778 B.n777 71.676
R1492 B.n779 B.n527 71.676
R1493 B.n786 B.n785 71.676
R1494 B.n787 B.n525 71.676
R1495 B.n794 B.n793 71.676
R1496 B.n795 B.n523 71.676
R1497 B.n802 B.n801 71.676
R1498 B.n803 B.n521 71.676
R1499 B.n810 B.n809 71.676
R1500 B.n811 B.n519 71.676
R1501 B.n818 B.n817 71.676
R1502 B.n819 B.n517 71.676
R1503 B.n826 B.n825 71.676
R1504 B.n827 B.n515 71.676
R1505 B.n834 B.n833 71.676
R1506 B.n837 B.n836 71.676
R1507 B.n1151 B.n1150 71.676
R1508 B.n1151 B.n2 71.676
R1509 B.n157 B.t18 68.0012
R1510 B.n717 B.t20 68.0012
R1511 B.n160 B.t11 67.9765
R1512 B.n549 B.t14 67.9765
R1513 B.n161 B.n160 59.5399
R1514 B.n158 B.n157 59.5399
R1515 B.n718 B.n717 59.5399
R1516 B.n698 B.n549 59.5399
R1517 B.n842 B.n511 59.0079
R1518 B.n1052 B.n1051 59.0079
R1519 B.n160 B.n159 53.3338
R1520 B.n157 B.n156 53.3338
R1521 B.n717 B.n716 53.3338
R1522 B.n549 B.n548 53.3338
R1523 B.n844 B.n509 35.4346
R1524 B.n840 B.n839 35.4346
R1525 B.n1048 B.n1047 35.4346
R1526 B.n1054 B.n88 35.4346
R1527 B.n842 B.n507 31.595
R1528 B.n848 B.n507 31.595
R1529 B.n848 B.n503 31.595
R1530 B.n854 B.n503 31.595
R1531 B.n854 B.n498 31.595
R1532 B.n860 B.n498 31.595
R1533 B.n860 B.n499 31.595
R1534 B.n866 B.n491 31.595
R1535 B.n872 B.n491 31.595
R1536 B.n872 B.n487 31.595
R1537 B.n878 B.n487 31.595
R1538 B.n878 B.n483 31.595
R1539 B.n884 B.n483 31.595
R1540 B.n884 B.n479 31.595
R1541 B.n890 B.n479 31.595
R1542 B.n890 B.n475 31.595
R1543 B.n896 B.n475 31.595
R1544 B.n902 B.n471 31.595
R1545 B.n902 B.n467 31.595
R1546 B.n908 B.n467 31.595
R1547 B.n908 B.n463 31.595
R1548 B.n914 B.n463 31.595
R1549 B.n914 B.n459 31.595
R1550 B.n920 B.n459 31.595
R1551 B.n926 B.n455 31.595
R1552 B.n926 B.n451 31.595
R1553 B.n932 B.n451 31.595
R1554 B.n932 B.n447 31.595
R1555 B.n938 B.n447 31.595
R1556 B.n938 B.n443 31.595
R1557 B.n944 B.n443 31.595
R1558 B.n950 B.n439 31.595
R1559 B.n950 B.n435 31.595
R1560 B.n956 B.n435 31.595
R1561 B.n956 B.n431 31.595
R1562 B.n962 B.n431 31.595
R1563 B.n962 B.n427 31.595
R1564 B.n968 B.n427 31.595
R1565 B.n975 B.n423 31.595
R1566 B.n975 B.n419 31.595
R1567 B.n981 B.n419 31.595
R1568 B.n981 B.n4 31.595
R1569 B.n1149 B.n4 31.595
R1570 B.n1149 B.n1148 31.595
R1571 B.n1148 B.n1147 31.595
R1572 B.n1147 B.n8 31.595
R1573 B.n12 B.n8 31.595
R1574 B.n1140 B.n12 31.595
R1575 B.n1140 B.n1139 31.595
R1576 B.n1138 B.n16 31.595
R1577 B.n1132 B.n16 31.595
R1578 B.n1132 B.n1131 31.595
R1579 B.n1131 B.n1130 31.595
R1580 B.n1130 B.n23 31.595
R1581 B.n1124 B.n23 31.595
R1582 B.n1124 B.n1123 31.595
R1583 B.n1122 B.n30 31.595
R1584 B.n1116 B.n30 31.595
R1585 B.n1116 B.n1115 31.595
R1586 B.n1115 B.n1114 31.595
R1587 B.n1114 B.n37 31.595
R1588 B.n1108 B.n37 31.595
R1589 B.n1108 B.n1107 31.595
R1590 B.n1106 B.n44 31.595
R1591 B.n1100 B.n44 31.595
R1592 B.n1100 B.n1099 31.595
R1593 B.n1099 B.n1098 31.595
R1594 B.n1098 B.n51 31.595
R1595 B.n1092 B.n51 31.595
R1596 B.n1092 B.n1091 31.595
R1597 B.n1090 B.n58 31.595
R1598 B.n1084 B.n58 31.595
R1599 B.n1084 B.n1083 31.595
R1600 B.n1083 B.n1082 31.595
R1601 B.n1082 B.n65 31.595
R1602 B.n1076 B.n65 31.595
R1603 B.n1076 B.n1075 31.595
R1604 B.n1075 B.n1074 31.595
R1605 B.n1074 B.n72 31.595
R1606 B.n1068 B.n72 31.595
R1607 B.n1067 B.n1066 31.595
R1608 B.n1066 B.n79 31.595
R1609 B.n1060 B.n79 31.595
R1610 B.n1060 B.n1059 31.595
R1611 B.n1059 B.n1058 31.595
R1612 B.n1058 B.n86 31.595
R1613 B.n1052 B.n86 31.595
R1614 B.n968 B.t0 26.9488
R1615 B.t6 B.n1138 26.9488
R1616 B.n944 B.t1 24.161
R1617 B.t7 B.n1122 24.161
R1618 B.n866 B.t13 22.3025
R1619 B.n1068 B.t9 22.3025
R1620 B.n920 B.t3 21.3733
R1621 B.t4 B.n1106 21.3733
R1622 B.n896 B.t2 18.5855
R1623 B.t5 B.n1090 18.5855
R1624 B B.n1152 18.0485
R1625 B.t2 B.n471 13.01
R1626 B.n1091 B.t5 13.01
R1627 B.n845 B.n844 10.6151
R1628 B.n846 B.n845 10.6151
R1629 B.n846 B.n501 10.6151
R1630 B.n856 B.n501 10.6151
R1631 B.n857 B.n856 10.6151
R1632 B.n858 B.n857 10.6151
R1633 B.n858 B.n493 10.6151
R1634 B.n868 B.n493 10.6151
R1635 B.n869 B.n868 10.6151
R1636 B.n870 B.n869 10.6151
R1637 B.n870 B.n485 10.6151
R1638 B.n880 B.n485 10.6151
R1639 B.n881 B.n880 10.6151
R1640 B.n882 B.n881 10.6151
R1641 B.n882 B.n477 10.6151
R1642 B.n892 B.n477 10.6151
R1643 B.n893 B.n892 10.6151
R1644 B.n894 B.n893 10.6151
R1645 B.n894 B.n469 10.6151
R1646 B.n904 B.n469 10.6151
R1647 B.n905 B.n904 10.6151
R1648 B.n906 B.n905 10.6151
R1649 B.n906 B.n461 10.6151
R1650 B.n916 B.n461 10.6151
R1651 B.n917 B.n916 10.6151
R1652 B.n918 B.n917 10.6151
R1653 B.n918 B.n453 10.6151
R1654 B.n928 B.n453 10.6151
R1655 B.n929 B.n928 10.6151
R1656 B.n930 B.n929 10.6151
R1657 B.n930 B.n445 10.6151
R1658 B.n940 B.n445 10.6151
R1659 B.n941 B.n940 10.6151
R1660 B.n942 B.n941 10.6151
R1661 B.n942 B.n437 10.6151
R1662 B.n952 B.n437 10.6151
R1663 B.n953 B.n952 10.6151
R1664 B.n954 B.n953 10.6151
R1665 B.n954 B.n429 10.6151
R1666 B.n964 B.n429 10.6151
R1667 B.n965 B.n964 10.6151
R1668 B.n966 B.n965 10.6151
R1669 B.n966 B.n421 10.6151
R1670 B.n977 B.n421 10.6151
R1671 B.n978 B.n977 10.6151
R1672 B.n979 B.n978 10.6151
R1673 B.n979 B.n0 10.6151
R1674 B.n579 B.n509 10.6151
R1675 B.n579 B.n578 10.6151
R1676 B.n585 B.n578 10.6151
R1677 B.n586 B.n585 10.6151
R1678 B.n587 B.n586 10.6151
R1679 B.n587 B.n576 10.6151
R1680 B.n593 B.n576 10.6151
R1681 B.n594 B.n593 10.6151
R1682 B.n595 B.n594 10.6151
R1683 B.n595 B.n574 10.6151
R1684 B.n601 B.n574 10.6151
R1685 B.n602 B.n601 10.6151
R1686 B.n603 B.n602 10.6151
R1687 B.n603 B.n572 10.6151
R1688 B.n609 B.n572 10.6151
R1689 B.n610 B.n609 10.6151
R1690 B.n611 B.n610 10.6151
R1691 B.n611 B.n570 10.6151
R1692 B.n617 B.n570 10.6151
R1693 B.n618 B.n617 10.6151
R1694 B.n619 B.n618 10.6151
R1695 B.n619 B.n568 10.6151
R1696 B.n625 B.n568 10.6151
R1697 B.n626 B.n625 10.6151
R1698 B.n627 B.n626 10.6151
R1699 B.n627 B.n566 10.6151
R1700 B.n633 B.n566 10.6151
R1701 B.n634 B.n633 10.6151
R1702 B.n635 B.n634 10.6151
R1703 B.n635 B.n564 10.6151
R1704 B.n641 B.n564 10.6151
R1705 B.n642 B.n641 10.6151
R1706 B.n643 B.n642 10.6151
R1707 B.n643 B.n562 10.6151
R1708 B.n649 B.n562 10.6151
R1709 B.n650 B.n649 10.6151
R1710 B.n651 B.n650 10.6151
R1711 B.n651 B.n560 10.6151
R1712 B.n657 B.n560 10.6151
R1713 B.n658 B.n657 10.6151
R1714 B.n659 B.n658 10.6151
R1715 B.n659 B.n558 10.6151
R1716 B.n665 B.n558 10.6151
R1717 B.n666 B.n665 10.6151
R1718 B.n667 B.n666 10.6151
R1719 B.n667 B.n556 10.6151
R1720 B.n673 B.n556 10.6151
R1721 B.n674 B.n673 10.6151
R1722 B.n675 B.n674 10.6151
R1723 B.n675 B.n554 10.6151
R1724 B.n681 B.n554 10.6151
R1725 B.n682 B.n681 10.6151
R1726 B.n683 B.n682 10.6151
R1727 B.n683 B.n552 10.6151
R1728 B.n689 B.n552 10.6151
R1729 B.n690 B.n689 10.6151
R1730 B.n691 B.n690 10.6151
R1731 B.n691 B.n550 10.6151
R1732 B.n697 B.n550 10.6151
R1733 B.n700 B.n699 10.6151
R1734 B.n700 B.n546 10.6151
R1735 B.n706 B.n546 10.6151
R1736 B.n707 B.n706 10.6151
R1737 B.n708 B.n707 10.6151
R1738 B.n708 B.n544 10.6151
R1739 B.n714 B.n544 10.6151
R1740 B.n715 B.n714 10.6151
R1741 B.n719 B.n715 10.6151
R1742 B.n725 B.n542 10.6151
R1743 B.n726 B.n725 10.6151
R1744 B.n727 B.n726 10.6151
R1745 B.n727 B.n540 10.6151
R1746 B.n733 B.n540 10.6151
R1747 B.n734 B.n733 10.6151
R1748 B.n735 B.n734 10.6151
R1749 B.n735 B.n538 10.6151
R1750 B.n741 B.n538 10.6151
R1751 B.n742 B.n741 10.6151
R1752 B.n743 B.n742 10.6151
R1753 B.n743 B.n536 10.6151
R1754 B.n749 B.n536 10.6151
R1755 B.n750 B.n749 10.6151
R1756 B.n751 B.n750 10.6151
R1757 B.n751 B.n534 10.6151
R1758 B.n757 B.n534 10.6151
R1759 B.n758 B.n757 10.6151
R1760 B.n759 B.n758 10.6151
R1761 B.n759 B.n532 10.6151
R1762 B.n765 B.n532 10.6151
R1763 B.n766 B.n765 10.6151
R1764 B.n767 B.n766 10.6151
R1765 B.n767 B.n530 10.6151
R1766 B.n773 B.n530 10.6151
R1767 B.n774 B.n773 10.6151
R1768 B.n775 B.n774 10.6151
R1769 B.n775 B.n528 10.6151
R1770 B.n781 B.n528 10.6151
R1771 B.n782 B.n781 10.6151
R1772 B.n783 B.n782 10.6151
R1773 B.n783 B.n526 10.6151
R1774 B.n789 B.n526 10.6151
R1775 B.n790 B.n789 10.6151
R1776 B.n791 B.n790 10.6151
R1777 B.n791 B.n524 10.6151
R1778 B.n797 B.n524 10.6151
R1779 B.n798 B.n797 10.6151
R1780 B.n799 B.n798 10.6151
R1781 B.n799 B.n522 10.6151
R1782 B.n805 B.n522 10.6151
R1783 B.n806 B.n805 10.6151
R1784 B.n807 B.n806 10.6151
R1785 B.n807 B.n520 10.6151
R1786 B.n813 B.n520 10.6151
R1787 B.n814 B.n813 10.6151
R1788 B.n815 B.n814 10.6151
R1789 B.n815 B.n518 10.6151
R1790 B.n821 B.n518 10.6151
R1791 B.n822 B.n821 10.6151
R1792 B.n823 B.n822 10.6151
R1793 B.n823 B.n516 10.6151
R1794 B.n829 B.n516 10.6151
R1795 B.n830 B.n829 10.6151
R1796 B.n831 B.n830 10.6151
R1797 B.n831 B.n514 10.6151
R1798 B.n514 B.n513 10.6151
R1799 B.n838 B.n513 10.6151
R1800 B.n839 B.n838 10.6151
R1801 B.n840 B.n505 10.6151
R1802 B.n850 B.n505 10.6151
R1803 B.n851 B.n850 10.6151
R1804 B.n852 B.n851 10.6151
R1805 B.n852 B.n496 10.6151
R1806 B.n862 B.n496 10.6151
R1807 B.n863 B.n862 10.6151
R1808 B.n864 B.n863 10.6151
R1809 B.n864 B.n489 10.6151
R1810 B.n874 B.n489 10.6151
R1811 B.n875 B.n874 10.6151
R1812 B.n876 B.n875 10.6151
R1813 B.n876 B.n481 10.6151
R1814 B.n886 B.n481 10.6151
R1815 B.n887 B.n886 10.6151
R1816 B.n888 B.n887 10.6151
R1817 B.n888 B.n473 10.6151
R1818 B.n898 B.n473 10.6151
R1819 B.n899 B.n898 10.6151
R1820 B.n900 B.n899 10.6151
R1821 B.n900 B.n465 10.6151
R1822 B.n910 B.n465 10.6151
R1823 B.n911 B.n910 10.6151
R1824 B.n912 B.n911 10.6151
R1825 B.n912 B.n457 10.6151
R1826 B.n922 B.n457 10.6151
R1827 B.n923 B.n922 10.6151
R1828 B.n924 B.n923 10.6151
R1829 B.n924 B.n449 10.6151
R1830 B.n934 B.n449 10.6151
R1831 B.n935 B.n934 10.6151
R1832 B.n936 B.n935 10.6151
R1833 B.n936 B.n441 10.6151
R1834 B.n946 B.n441 10.6151
R1835 B.n947 B.n946 10.6151
R1836 B.n948 B.n947 10.6151
R1837 B.n948 B.n433 10.6151
R1838 B.n958 B.n433 10.6151
R1839 B.n959 B.n958 10.6151
R1840 B.n960 B.n959 10.6151
R1841 B.n960 B.n425 10.6151
R1842 B.n970 B.n425 10.6151
R1843 B.n971 B.n970 10.6151
R1844 B.n973 B.n971 10.6151
R1845 B.n973 B.n972 10.6151
R1846 B.n972 B.n417 10.6151
R1847 B.n984 B.n417 10.6151
R1848 B.n985 B.n984 10.6151
R1849 B.n986 B.n985 10.6151
R1850 B.n987 B.n986 10.6151
R1851 B.n988 B.n987 10.6151
R1852 B.n991 B.n988 10.6151
R1853 B.n992 B.n991 10.6151
R1854 B.n993 B.n992 10.6151
R1855 B.n994 B.n993 10.6151
R1856 B.n996 B.n994 10.6151
R1857 B.n997 B.n996 10.6151
R1858 B.n998 B.n997 10.6151
R1859 B.n999 B.n998 10.6151
R1860 B.n1001 B.n999 10.6151
R1861 B.n1002 B.n1001 10.6151
R1862 B.n1003 B.n1002 10.6151
R1863 B.n1004 B.n1003 10.6151
R1864 B.n1006 B.n1004 10.6151
R1865 B.n1007 B.n1006 10.6151
R1866 B.n1008 B.n1007 10.6151
R1867 B.n1009 B.n1008 10.6151
R1868 B.n1011 B.n1009 10.6151
R1869 B.n1012 B.n1011 10.6151
R1870 B.n1013 B.n1012 10.6151
R1871 B.n1014 B.n1013 10.6151
R1872 B.n1016 B.n1014 10.6151
R1873 B.n1017 B.n1016 10.6151
R1874 B.n1018 B.n1017 10.6151
R1875 B.n1019 B.n1018 10.6151
R1876 B.n1021 B.n1019 10.6151
R1877 B.n1022 B.n1021 10.6151
R1878 B.n1023 B.n1022 10.6151
R1879 B.n1024 B.n1023 10.6151
R1880 B.n1026 B.n1024 10.6151
R1881 B.n1027 B.n1026 10.6151
R1882 B.n1028 B.n1027 10.6151
R1883 B.n1029 B.n1028 10.6151
R1884 B.n1031 B.n1029 10.6151
R1885 B.n1032 B.n1031 10.6151
R1886 B.n1033 B.n1032 10.6151
R1887 B.n1034 B.n1033 10.6151
R1888 B.n1036 B.n1034 10.6151
R1889 B.n1037 B.n1036 10.6151
R1890 B.n1038 B.n1037 10.6151
R1891 B.n1039 B.n1038 10.6151
R1892 B.n1041 B.n1039 10.6151
R1893 B.n1042 B.n1041 10.6151
R1894 B.n1043 B.n1042 10.6151
R1895 B.n1044 B.n1043 10.6151
R1896 B.n1046 B.n1044 10.6151
R1897 B.n1047 B.n1046 10.6151
R1898 B.n1144 B.n1 10.6151
R1899 B.n1144 B.n1143 10.6151
R1900 B.n1143 B.n1142 10.6151
R1901 B.n1142 B.n10 10.6151
R1902 B.n1136 B.n10 10.6151
R1903 B.n1136 B.n1135 10.6151
R1904 B.n1135 B.n1134 10.6151
R1905 B.n1134 B.n18 10.6151
R1906 B.n1128 B.n18 10.6151
R1907 B.n1128 B.n1127 10.6151
R1908 B.n1127 B.n1126 10.6151
R1909 B.n1126 B.n25 10.6151
R1910 B.n1120 B.n25 10.6151
R1911 B.n1120 B.n1119 10.6151
R1912 B.n1119 B.n1118 10.6151
R1913 B.n1118 B.n32 10.6151
R1914 B.n1112 B.n32 10.6151
R1915 B.n1112 B.n1111 10.6151
R1916 B.n1111 B.n1110 10.6151
R1917 B.n1110 B.n39 10.6151
R1918 B.n1104 B.n39 10.6151
R1919 B.n1104 B.n1103 10.6151
R1920 B.n1103 B.n1102 10.6151
R1921 B.n1102 B.n46 10.6151
R1922 B.n1096 B.n46 10.6151
R1923 B.n1096 B.n1095 10.6151
R1924 B.n1095 B.n1094 10.6151
R1925 B.n1094 B.n53 10.6151
R1926 B.n1088 B.n53 10.6151
R1927 B.n1088 B.n1087 10.6151
R1928 B.n1087 B.n1086 10.6151
R1929 B.n1086 B.n60 10.6151
R1930 B.n1080 B.n60 10.6151
R1931 B.n1080 B.n1079 10.6151
R1932 B.n1079 B.n1078 10.6151
R1933 B.n1078 B.n67 10.6151
R1934 B.n1072 B.n67 10.6151
R1935 B.n1072 B.n1071 10.6151
R1936 B.n1071 B.n1070 10.6151
R1937 B.n1070 B.n74 10.6151
R1938 B.n1064 B.n74 10.6151
R1939 B.n1064 B.n1063 10.6151
R1940 B.n1063 B.n1062 10.6151
R1941 B.n1062 B.n81 10.6151
R1942 B.n1056 B.n81 10.6151
R1943 B.n1056 B.n1055 10.6151
R1944 B.n1055 B.n1054 10.6151
R1945 B.n162 B.n88 10.6151
R1946 B.n165 B.n162 10.6151
R1947 B.n166 B.n165 10.6151
R1948 B.n169 B.n166 10.6151
R1949 B.n170 B.n169 10.6151
R1950 B.n173 B.n170 10.6151
R1951 B.n174 B.n173 10.6151
R1952 B.n177 B.n174 10.6151
R1953 B.n178 B.n177 10.6151
R1954 B.n181 B.n178 10.6151
R1955 B.n182 B.n181 10.6151
R1956 B.n185 B.n182 10.6151
R1957 B.n186 B.n185 10.6151
R1958 B.n189 B.n186 10.6151
R1959 B.n190 B.n189 10.6151
R1960 B.n193 B.n190 10.6151
R1961 B.n194 B.n193 10.6151
R1962 B.n197 B.n194 10.6151
R1963 B.n198 B.n197 10.6151
R1964 B.n201 B.n198 10.6151
R1965 B.n202 B.n201 10.6151
R1966 B.n205 B.n202 10.6151
R1967 B.n206 B.n205 10.6151
R1968 B.n209 B.n206 10.6151
R1969 B.n210 B.n209 10.6151
R1970 B.n213 B.n210 10.6151
R1971 B.n214 B.n213 10.6151
R1972 B.n217 B.n214 10.6151
R1973 B.n218 B.n217 10.6151
R1974 B.n221 B.n218 10.6151
R1975 B.n222 B.n221 10.6151
R1976 B.n225 B.n222 10.6151
R1977 B.n226 B.n225 10.6151
R1978 B.n229 B.n226 10.6151
R1979 B.n230 B.n229 10.6151
R1980 B.n233 B.n230 10.6151
R1981 B.n234 B.n233 10.6151
R1982 B.n237 B.n234 10.6151
R1983 B.n238 B.n237 10.6151
R1984 B.n241 B.n238 10.6151
R1985 B.n242 B.n241 10.6151
R1986 B.n245 B.n242 10.6151
R1987 B.n246 B.n245 10.6151
R1988 B.n249 B.n246 10.6151
R1989 B.n250 B.n249 10.6151
R1990 B.n253 B.n250 10.6151
R1991 B.n254 B.n253 10.6151
R1992 B.n257 B.n254 10.6151
R1993 B.n258 B.n257 10.6151
R1994 B.n261 B.n258 10.6151
R1995 B.n262 B.n261 10.6151
R1996 B.n265 B.n262 10.6151
R1997 B.n266 B.n265 10.6151
R1998 B.n269 B.n266 10.6151
R1999 B.n270 B.n269 10.6151
R2000 B.n273 B.n270 10.6151
R2001 B.n274 B.n273 10.6151
R2002 B.n277 B.n274 10.6151
R2003 B.n278 B.n277 10.6151
R2004 B.n282 B.n281 10.6151
R2005 B.n285 B.n282 10.6151
R2006 B.n286 B.n285 10.6151
R2007 B.n289 B.n286 10.6151
R2008 B.n290 B.n289 10.6151
R2009 B.n293 B.n290 10.6151
R2010 B.n294 B.n293 10.6151
R2011 B.n297 B.n294 10.6151
R2012 B.n298 B.n297 10.6151
R2013 B.n302 B.n301 10.6151
R2014 B.n305 B.n302 10.6151
R2015 B.n306 B.n305 10.6151
R2016 B.n309 B.n306 10.6151
R2017 B.n310 B.n309 10.6151
R2018 B.n313 B.n310 10.6151
R2019 B.n314 B.n313 10.6151
R2020 B.n317 B.n314 10.6151
R2021 B.n318 B.n317 10.6151
R2022 B.n321 B.n318 10.6151
R2023 B.n322 B.n321 10.6151
R2024 B.n325 B.n322 10.6151
R2025 B.n326 B.n325 10.6151
R2026 B.n329 B.n326 10.6151
R2027 B.n330 B.n329 10.6151
R2028 B.n333 B.n330 10.6151
R2029 B.n334 B.n333 10.6151
R2030 B.n337 B.n334 10.6151
R2031 B.n338 B.n337 10.6151
R2032 B.n341 B.n338 10.6151
R2033 B.n342 B.n341 10.6151
R2034 B.n345 B.n342 10.6151
R2035 B.n346 B.n345 10.6151
R2036 B.n349 B.n346 10.6151
R2037 B.n350 B.n349 10.6151
R2038 B.n353 B.n350 10.6151
R2039 B.n354 B.n353 10.6151
R2040 B.n357 B.n354 10.6151
R2041 B.n358 B.n357 10.6151
R2042 B.n361 B.n358 10.6151
R2043 B.n362 B.n361 10.6151
R2044 B.n365 B.n362 10.6151
R2045 B.n366 B.n365 10.6151
R2046 B.n369 B.n366 10.6151
R2047 B.n370 B.n369 10.6151
R2048 B.n373 B.n370 10.6151
R2049 B.n374 B.n373 10.6151
R2050 B.n377 B.n374 10.6151
R2051 B.n378 B.n377 10.6151
R2052 B.n381 B.n378 10.6151
R2053 B.n382 B.n381 10.6151
R2054 B.n385 B.n382 10.6151
R2055 B.n386 B.n385 10.6151
R2056 B.n389 B.n386 10.6151
R2057 B.n390 B.n389 10.6151
R2058 B.n393 B.n390 10.6151
R2059 B.n394 B.n393 10.6151
R2060 B.n397 B.n394 10.6151
R2061 B.n398 B.n397 10.6151
R2062 B.n401 B.n398 10.6151
R2063 B.n402 B.n401 10.6151
R2064 B.n405 B.n402 10.6151
R2065 B.n406 B.n405 10.6151
R2066 B.n409 B.n406 10.6151
R2067 B.n410 B.n409 10.6151
R2068 B.n413 B.n410 10.6151
R2069 B.n415 B.n413 10.6151
R2070 B.n416 B.n415 10.6151
R2071 B.n1048 B.n416 10.6151
R2072 B.t3 B.n455 10.2223
R2073 B.n1107 B.t4 10.2223
R2074 B.n698 B.n697 9.36635
R2075 B.n718 B.n542 9.36635
R2076 B.n278 B.n161 9.36635
R2077 B.n301 B.n158 9.36635
R2078 B.n499 B.t13 9.293
R2079 B.t9 B.n1067 9.293
R2080 B.n1152 B.n0 8.11757
R2081 B.n1152 B.n1 8.11757
R2082 B.t1 B.n439 7.4345
R2083 B.n1123 B.t7 7.4345
R2084 B.t0 B.n423 4.64675
R2085 B.n1139 B.t6 4.64675
R2086 B.n699 B.n698 1.24928
R2087 B.n719 B.n718 1.24928
R2088 B.n281 B.n161 1.24928
R2089 B.n298 B.n158 1.24928
R2090 VP.n16 VP.t0 215.745
R2091 VP.n9 VP.t4 183.24
R2092 VP.n47 VP.t2 183.24
R2093 VP.n3 VP.t7 183.24
R2094 VP.n65 VP.t3 183.24
R2095 VP.n35 VP.t5 183.24
R2096 VP.n13 VP.t6 183.24
R2097 VP.n17 VP.t1 183.24
R2098 VP.n19 VP.n18 161.3
R2099 VP.n20 VP.n15 161.3
R2100 VP.n22 VP.n21 161.3
R2101 VP.n23 VP.n14 161.3
R2102 VP.n25 VP.n24 161.3
R2103 VP.n27 VP.n26 161.3
R2104 VP.n28 VP.n12 161.3
R2105 VP.n30 VP.n29 161.3
R2106 VP.n31 VP.n11 161.3
R2107 VP.n33 VP.n32 161.3
R2108 VP.n34 VP.n10 161.3
R2109 VP.n64 VP.n0 161.3
R2110 VP.n63 VP.n62 161.3
R2111 VP.n61 VP.n1 161.3
R2112 VP.n60 VP.n59 161.3
R2113 VP.n58 VP.n2 161.3
R2114 VP.n57 VP.n56 161.3
R2115 VP.n55 VP.n54 161.3
R2116 VP.n53 VP.n4 161.3
R2117 VP.n52 VP.n51 161.3
R2118 VP.n50 VP.n5 161.3
R2119 VP.n49 VP.n48 161.3
R2120 VP.n46 VP.n6 161.3
R2121 VP.n45 VP.n44 161.3
R2122 VP.n43 VP.n7 161.3
R2123 VP.n42 VP.n41 161.3
R2124 VP.n40 VP.n8 161.3
R2125 VP.n39 VP.n38 161.3
R2126 VP.n37 VP.n9 104.76
R2127 VP.n66 VP.n65 104.76
R2128 VP.n36 VP.n35 104.76
R2129 VP.n41 VP.n7 56.5617
R2130 VP.n59 VP.n1 56.5617
R2131 VP.n29 VP.n11 56.5617
R2132 VP.n37 VP.n36 54.8178
R2133 VP.n17 VP.n16 53.9941
R2134 VP.n52 VP.n5 40.577
R2135 VP.n53 VP.n52 40.577
R2136 VP.n23 VP.n22 40.577
R2137 VP.n22 VP.n15 40.577
R2138 VP.n40 VP.n39 24.5923
R2139 VP.n41 VP.n40 24.5923
R2140 VP.n45 VP.n7 24.5923
R2141 VP.n46 VP.n45 24.5923
R2142 VP.n48 VP.n5 24.5923
R2143 VP.n54 VP.n53 24.5923
R2144 VP.n58 VP.n57 24.5923
R2145 VP.n59 VP.n58 24.5923
R2146 VP.n63 VP.n1 24.5923
R2147 VP.n64 VP.n63 24.5923
R2148 VP.n33 VP.n11 24.5923
R2149 VP.n34 VP.n33 24.5923
R2150 VP.n24 VP.n23 24.5923
R2151 VP.n28 VP.n27 24.5923
R2152 VP.n29 VP.n28 24.5923
R2153 VP.n18 VP.n15 24.5923
R2154 VP.n48 VP.n47 18.4444
R2155 VP.n54 VP.n3 18.4444
R2156 VP.n24 VP.n13 18.4444
R2157 VP.n18 VP.n17 18.4444
R2158 VP.n19 VP.n16 7.07482
R2159 VP.n39 VP.n9 6.14846
R2160 VP.n47 VP.n46 6.14846
R2161 VP.n57 VP.n3 6.14846
R2162 VP.n65 VP.n64 6.14846
R2163 VP.n35 VP.n34 6.14846
R2164 VP.n27 VP.n13 6.14846
R2165 VP.n36 VP.n10 0.278335
R2166 VP.n38 VP.n37 0.278335
R2167 VP.n66 VP.n0 0.278335
R2168 VP.n20 VP.n19 0.189894
R2169 VP.n21 VP.n20 0.189894
R2170 VP.n21 VP.n14 0.189894
R2171 VP.n25 VP.n14 0.189894
R2172 VP.n26 VP.n25 0.189894
R2173 VP.n26 VP.n12 0.189894
R2174 VP.n30 VP.n12 0.189894
R2175 VP.n31 VP.n30 0.189894
R2176 VP.n32 VP.n31 0.189894
R2177 VP.n32 VP.n10 0.189894
R2178 VP.n38 VP.n8 0.189894
R2179 VP.n42 VP.n8 0.189894
R2180 VP.n43 VP.n42 0.189894
R2181 VP.n44 VP.n43 0.189894
R2182 VP.n44 VP.n6 0.189894
R2183 VP.n49 VP.n6 0.189894
R2184 VP.n50 VP.n49 0.189894
R2185 VP.n51 VP.n50 0.189894
R2186 VP.n51 VP.n4 0.189894
R2187 VP.n55 VP.n4 0.189894
R2188 VP.n56 VP.n55 0.189894
R2189 VP.n56 VP.n2 0.189894
R2190 VP.n60 VP.n2 0.189894
R2191 VP.n61 VP.n60 0.189894
R2192 VP.n62 VP.n61 0.189894
R2193 VP.n62 VP.n0 0.189894
R2194 VP VP.n66 0.153485
R2195 VDD1 VDD1.n0 64.4844
R2196 VDD1.n3 VDD1.n2 64.3706
R2197 VDD1.n3 VDD1.n1 64.3706
R2198 VDD1.n5 VDD1.n4 63.2398
R2199 VDD1.n5 VDD1.n3 50.8285
R2200 VDD1 VDD1.n5 1.12766
R2201 VDD1.n4 VDD1.t1 1.07659
R2202 VDD1.n4 VDD1.t2 1.07659
R2203 VDD1.n0 VDD1.t7 1.07659
R2204 VDD1.n0 VDD1.t6 1.07659
R2205 VDD1.n2 VDD1.t0 1.07659
R2206 VDD1.n2 VDD1.t4 1.07659
R2207 VDD1.n1 VDD1.t3 1.07659
R2208 VDD1.n1 VDD1.t5 1.07659
C0 VDD2 VDD1 1.68443f
C1 VTAIL VDD2 10.346999f
C2 VP VN 8.62622f
C3 VP VDD1 13.2453f
C4 VTAIL VP 12.9775f
C5 VP VDD2 0.500949f
C6 VDD1 VN 0.151835f
C7 VTAIL VN 12.963401f
C8 VTAIL VDD1 10.2938f
C9 VDD2 VN 12.8975f
C10 VDD2 B 5.661216f
C11 VDD1 B 6.076883f
C12 VTAIL B 14.176244f
C13 VN B 15.374169f
C14 VP B 13.818741f
C15 VDD1.t7 B 0.357076f
C16 VDD1.t6 B 0.357076f
C17 VDD1.n0 B 3.27408f
C18 VDD1.t3 B 0.357076f
C19 VDD1.t5 B 0.357076f
C20 VDD1.n1 B 3.27308f
C21 VDD1.t0 B 0.357076f
C22 VDD1.t4 B 0.357076f
C23 VDD1.n2 B 3.27308f
C24 VDD1.n3 B 3.55276f
C25 VDD1.t1 B 0.357076f
C26 VDD1.t2 B 0.357076f
C27 VDD1.n4 B 3.2646f
C28 VDD1.n5 B 3.33629f
C29 VP.n0 B 0.029561f
C30 VP.t3 B 2.74741f
C31 VP.n1 B 0.032595f
C32 VP.n2 B 0.022423f
C33 VP.t7 B 2.74741f
C34 VP.n3 B 0.953227f
C35 VP.n4 B 0.022423f
C36 VP.n5 B 0.04433f
C37 VP.n6 B 0.022423f
C38 VP.t2 B 2.74741f
C39 VP.n7 B 0.032595f
C40 VP.n8 B 0.022423f
C41 VP.t4 B 2.74741f
C42 VP.n9 B 1.01798f
C43 VP.n10 B 0.029561f
C44 VP.t5 B 2.74741f
C45 VP.n11 B 0.032595f
C46 VP.n12 B 0.022423f
C47 VP.t6 B 2.74741f
C48 VP.n13 B 0.953227f
C49 VP.n14 B 0.022423f
C50 VP.n15 B 0.04433f
C51 VP.t0 B 2.91059f
C52 VP.n16 B 1.00061f
C53 VP.t1 B 2.74741f
C54 VP.n17 B 1.02031f
C55 VP.n18 B 0.036449f
C56 VP.n19 B 0.212249f
C57 VP.n20 B 0.022423f
C58 VP.n21 B 0.022423f
C59 VP.n22 B 0.01811f
C60 VP.n23 B 0.04433f
C61 VP.n24 B 0.036449f
C62 VP.n25 B 0.022423f
C63 VP.n26 B 0.022423f
C64 VP.n27 B 0.026185f
C65 VP.n28 B 0.041581f
C66 VP.n29 B 0.032595f
C67 VP.n30 B 0.022423f
C68 VP.n31 B 0.022423f
C69 VP.n32 B 0.022423f
C70 VP.n33 B 0.041581f
C71 VP.n34 B 0.026185f
C72 VP.n35 B 1.01798f
C73 VP.n36 B 1.42369f
C74 VP.n37 B 1.43843f
C75 VP.n38 B 0.029561f
C76 VP.n39 B 0.026185f
C77 VP.n40 B 0.041581f
C78 VP.n41 B 0.032595f
C79 VP.n42 B 0.022423f
C80 VP.n43 B 0.022423f
C81 VP.n44 B 0.022423f
C82 VP.n45 B 0.041581f
C83 VP.n46 B 0.026185f
C84 VP.n47 B 0.953227f
C85 VP.n48 B 0.036449f
C86 VP.n49 B 0.022423f
C87 VP.n50 B 0.022423f
C88 VP.n51 B 0.022423f
C89 VP.n52 B 0.01811f
C90 VP.n53 B 0.04433f
C91 VP.n54 B 0.036449f
C92 VP.n55 B 0.022423f
C93 VP.n56 B 0.022423f
C94 VP.n57 B 0.026185f
C95 VP.n58 B 0.041581f
C96 VP.n59 B 0.032595f
C97 VP.n60 B 0.022423f
C98 VP.n61 B 0.022423f
C99 VP.n62 B 0.022423f
C100 VP.n63 B 0.041581f
C101 VP.n64 B 0.026185f
C102 VP.n65 B 1.01798f
C103 VP.n66 B 0.037076f
C104 VDD2.t2 B 0.353883f
C105 VDD2.t7 B 0.353883f
C106 VDD2.n0 B 3.24381f
C107 VDD2.t3 B 0.353883f
C108 VDD2.t0 B 0.353883f
C109 VDD2.n1 B 3.24381f
C110 VDD2.n2 B 3.47048f
C111 VDD2.t4 B 0.353883f
C112 VDD2.t6 B 0.353883f
C113 VDD2.n3 B 3.23541f
C114 VDD2.n4 B 3.27621f
C115 VDD2.t1 B 0.353883f
C116 VDD2.t5 B 0.353883f
C117 VDD2.n5 B 3.24378f
C118 VTAIL.t9 B 0.268279f
C119 VTAIL.t12 B 0.268279f
C120 VTAIL.n0 B 2.40141f
C121 VTAIL.n1 B 0.317586f
C122 VTAIL.t7 B 3.06838f
C123 VTAIL.n2 B 0.406762f
C124 VTAIL.t0 B 3.06838f
C125 VTAIL.n3 B 0.406762f
C126 VTAIL.t3 B 0.268279f
C127 VTAIL.t1 B 0.268279f
C128 VTAIL.n4 B 2.40141f
C129 VTAIL.n5 B 0.45507f
C130 VTAIL.t2 B 3.06838f
C131 VTAIL.n6 B 1.71345f
C132 VTAIL.t14 B 3.06837f
C133 VTAIL.n7 B 1.71346f
C134 VTAIL.t10 B 0.268279f
C135 VTAIL.t11 B 0.268279f
C136 VTAIL.n8 B 2.40141f
C137 VTAIL.n9 B 0.455069f
C138 VTAIL.t13 B 3.06837f
C139 VTAIL.n10 B 0.40677f
C140 VTAIL.t6 B 3.06837f
C141 VTAIL.n11 B 0.40677f
C142 VTAIL.t15 B 0.268279f
C143 VTAIL.t4 B 0.268279f
C144 VTAIL.n12 B 2.40141f
C145 VTAIL.n13 B 0.455069f
C146 VTAIL.t5 B 3.06837f
C147 VTAIL.n14 B 1.71346f
C148 VTAIL.t8 B 3.06838f
C149 VTAIL.n15 B 1.70999f
C150 VN.n0 B 0.029279f
C151 VN.t7 B 2.72126f
C152 VN.n1 B 0.032285f
C153 VN.n2 B 0.022209f
C154 VN.t4 B 2.72126f
C155 VN.n3 B 0.944155f
C156 VN.n4 B 0.022209f
C157 VN.n5 B 0.043908f
C158 VN.t5 B 2.88288f
C159 VN.n6 B 0.991087f
C160 VN.t0 B 2.72126f
C161 VN.n7 B 1.0106f
C162 VN.n8 B 0.036102f
C163 VN.n9 B 0.210229f
C164 VN.n10 B 0.022209f
C165 VN.n11 B 0.022209f
C166 VN.n12 B 0.017938f
C167 VN.n13 B 0.043908f
C168 VN.n14 B 0.036102f
C169 VN.n15 B 0.022209f
C170 VN.n16 B 0.022209f
C171 VN.n17 B 0.025936f
C172 VN.n18 B 0.041185f
C173 VN.n19 B 0.032285f
C174 VN.n20 B 0.022209f
C175 VN.n21 B 0.022209f
C176 VN.n22 B 0.022209f
C177 VN.n23 B 0.041185f
C178 VN.n24 B 0.025936f
C179 VN.n25 B 1.00829f
C180 VN.n26 B 0.036723f
C181 VN.n27 B 0.029279f
C182 VN.t3 B 2.72126f
C183 VN.n28 B 0.032285f
C184 VN.n29 B 0.022209f
C185 VN.t1 B 2.72126f
C186 VN.n30 B 0.944155f
C187 VN.n31 B 0.022209f
C188 VN.n32 B 0.043908f
C189 VN.t2 B 2.88288f
C190 VN.n33 B 0.991087f
C191 VN.t6 B 2.72126f
C192 VN.n34 B 1.0106f
C193 VN.n35 B 0.036102f
C194 VN.n36 B 0.210229f
C195 VN.n37 B 0.022209f
C196 VN.n38 B 0.022209f
C197 VN.n39 B 0.017938f
C198 VN.n40 B 0.043908f
C199 VN.n41 B 0.036102f
C200 VN.n42 B 0.022209f
C201 VN.n43 B 0.022209f
C202 VN.n44 B 0.025936f
C203 VN.n45 B 0.041185f
C204 VN.n46 B 0.032285f
C205 VN.n47 B 0.022209f
C206 VN.n48 B 0.022209f
C207 VN.n49 B 0.022209f
C208 VN.n50 B 0.041185f
C209 VN.n51 B 0.025936f
C210 VN.n52 B 1.00829f
C211 VN.n53 B 1.42191f
.ends

