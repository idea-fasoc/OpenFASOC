* NGSPICE file created from diff_pair_sample_0432.ext - technology: sky130A

.subckt diff_pair_sample_0432 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X1 VTAIL.t5 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X2 VTAIL.t13 VP.t1 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X3 VDD2.t6 VN.t1 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X4 VDD1.t5 VP.t2 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=0 ps=0 w=11.52 l=1.02
X6 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X7 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=0 ps=0 w=11.52 l=1.02
X8 VDD1.t2 VP.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X9 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=4.4928 ps=23.82 w=11.52 l=1.02
X10 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=1.9008 ps=11.85 w=11.52 l=1.02
X11 VDD1.t6 VP.t4 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=4.4928 ps=23.82 w=11.52 l=1.02
X12 VTAIL.t9 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=1.9008 ps=11.85 w=11.52 l=1.02
X13 VTAIL.t8 VP.t6 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=1.9008 ps=11.85 w=11.52 l=1.02
X14 VDD2.t2 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=4.4928 ps=23.82 w=11.52 l=1.02
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=0 ps=0 w=11.52 l=1.02
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=0 ps=0 w=11.52 l=1.02
X17 VDD1.t7 VP.t7 VTAIL.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=4.4928 ps=23.82 w=11.52 l=1.02
X18 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9008 pd=11.85 as=1.9008 ps=11.85 w=11.52 l=1.02
X19 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4928 pd=23.82 as=1.9008 ps=11.85 w=11.52 l=1.02
R0 VP.n9 VP.t6 326.95
R1 VP.n21 VP.t5 310.702
R2 VP.n33 VP.t4 310.702
R3 VP.n18 VP.t7 310.702
R4 VP.n3 VP.t2 272.188
R5 VP.n1 VP.t0 272.188
R6 VP.n6 VP.t1 272.188
R7 VP.n8 VP.t3 272.188
R8 VP.n34 VP.n33 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n12 VP.n7 161.3
R11 VP.n14 VP.n13 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n5 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n32 VP.n0 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n29 VP.n28 161.3
R18 VP.n27 VP.n2 161.3
R19 VP.n26 VP.n25 161.3
R20 VP.n24 VP.n23 161.3
R21 VP.n22 VP.n4 161.3
R22 VP.n21 VP.n20 161.3
R23 VP.n23 VP.n22 55.1086
R24 VP.n32 VP.n31 55.1086
R25 VP.n17 VP.n16 55.1086
R26 VP.n9 VP.n8 46.4196
R27 VP.n10 VP.n9 43.7016
R28 VP.n20 VP.n19 43.1899
R29 VP.n27 VP.n26 40.577
R30 VP.n28 VP.n27 40.577
R31 VP.n13 VP.n12 40.577
R32 VP.n12 VP.n11 40.577
R33 VP.n23 VP.n3 15.9852
R34 VP.n31 VP.n1 15.9852
R35 VP.n16 VP.n6 15.9852
R36 VP.n26 VP.n3 8.60764
R37 VP.n28 VP.n1 8.60764
R38 VP.n13 VP.n6 8.60764
R39 VP.n11 VP.n8 8.60764
R40 VP.n22 VP.n21 2.19141
R41 VP.n33 VP.n32 2.19141
R42 VP.n18 VP.n17 2.19141
R43 VP.n10 VP.n7 0.189894
R44 VP.n14 VP.n7 0.189894
R45 VP.n15 VP.n14 0.189894
R46 VP.n15 VP.n5 0.189894
R47 VP.n19 VP.n5 0.189894
R48 VP.n20 VP.n4 0.189894
R49 VP.n24 VP.n4 0.189894
R50 VP.n25 VP.n24 0.189894
R51 VP.n25 VP.n2 0.189894
R52 VP.n29 VP.n2 0.189894
R53 VP.n30 VP.n29 0.189894
R54 VP.n30 VP.n0 0.189894
R55 VP.n34 VP.n0 0.189894
R56 VP VP.n34 0.0516364
R57 VDD1 VDD1.n0 65.0573
R58 VDD1.n3 VDD1.n2 64.9436
R59 VDD1.n3 VDD1.n1 64.9436
R60 VDD1.n5 VDD1.n4 64.417
R61 VDD1.n5 VDD1.n3 39.4664
R62 VDD1.n4 VDD1.t3 1.71925
R63 VDD1.n4 VDD1.t7 1.71925
R64 VDD1.n0 VDD1.t4 1.71925
R65 VDD1.n0 VDD1.t2 1.71925
R66 VDD1.n2 VDD1.t1 1.71925
R67 VDD1.n2 VDD1.t6 1.71925
R68 VDD1.n1 VDD1.t0 1.71925
R69 VDD1.n1 VDD1.t5 1.71925
R70 VDD1 VDD1.n5 0.524207
R71 VTAIL.n498 VTAIL.n442 289.615
R72 VTAIL.n58 VTAIL.n2 289.615
R73 VTAIL.n120 VTAIL.n64 289.615
R74 VTAIL.n184 VTAIL.n128 289.615
R75 VTAIL.n436 VTAIL.n380 289.615
R76 VTAIL.n372 VTAIL.n316 289.615
R77 VTAIL.n310 VTAIL.n254 289.615
R78 VTAIL.n246 VTAIL.n190 289.615
R79 VTAIL.n463 VTAIL.n462 185
R80 VTAIL.n465 VTAIL.n464 185
R81 VTAIL.n458 VTAIL.n457 185
R82 VTAIL.n471 VTAIL.n470 185
R83 VTAIL.n473 VTAIL.n472 185
R84 VTAIL.n454 VTAIL.n453 185
R85 VTAIL.n480 VTAIL.n479 185
R86 VTAIL.n481 VTAIL.n452 185
R87 VTAIL.n483 VTAIL.n482 185
R88 VTAIL.n450 VTAIL.n449 185
R89 VTAIL.n489 VTAIL.n488 185
R90 VTAIL.n491 VTAIL.n490 185
R91 VTAIL.n446 VTAIL.n445 185
R92 VTAIL.n497 VTAIL.n496 185
R93 VTAIL.n499 VTAIL.n498 185
R94 VTAIL.n23 VTAIL.n22 185
R95 VTAIL.n25 VTAIL.n24 185
R96 VTAIL.n18 VTAIL.n17 185
R97 VTAIL.n31 VTAIL.n30 185
R98 VTAIL.n33 VTAIL.n32 185
R99 VTAIL.n14 VTAIL.n13 185
R100 VTAIL.n40 VTAIL.n39 185
R101 VTAIL.n41 VTAIL.n12 185
R102 VTAIL.n43 VTAIL.n42 185
R103 VTAIL.n10 VTAIL.n9 185
R104 VTAIL.n49 VTAIL.n48 185
R105 VTAIL.n51 VTAIL.n50 185
R106 VTAIL.n6 VTAIL.n5 185
R107 VTAIL.n57 VTAIL.n56 185
R108 VTAIL.n59 VTAIL.n58 185
R109 VTAIL.n85 VTAIL.n84 185
R110 VTAIL.n87 VTAIL.n86 185
R111 VTAIL.n80 VTAIL.n79 185
R112 VTAIL.n93 VTAIL.n92 185
R113 VTAIL.n95 VTAIL.n94 185
R114 VTAIL.n76 VTAIL.n75 185
R115 VTAIL.n102 VTAIL.n101 185
R116 VTAIL.n103 VTAIL.n74 185
R117 VTAIL.n105 VTAIL.n104 185
R118 VTAIL.n72 VTAIL.n71 185
R119 VTAIL.n111 VTAIL.n110 185
R120 VTAIL.n113 VTAIL.n112 185
R121 VTAIL.n68 VTAIL.n67 185
R122 VTAIL.n119 VTAIL.n118 185
R123 VTAIL.n121 VTAIL.n120 185
R124 VTAIL.n149 VTAIL.n148 185
R125 VTAIL.n151 VTAIL.n150 185
R126 VTAIL.n144 VTAIL.n143 185
R127 VTAIL.n157 VTAIL.n156 185
R128 VTAIL.n159 VTAIL.n158 185
R129 VTAIL.n140 VTAIL.n139 185
R130 VTAIL.n166 VTAIL.n165 185
R131 VTAIL.n167 VTAIL.n138 185
R132 VTAIL.n169 VTAIL.n168 185
R133 VTAIL.n136 VTAIL.n135 185
R134 VTAIL.n175 VTAIL.n174 185
R135 VTAIL.n177 VTAIL.n176 185
R136 VTAIL.n132 VTAIL.n131 185
R137 VTAIL.n183 VTAIL.n182 185
R138 VTAIL.n185 VTAIL.n184 185
R139 VTAIL.n437 VTAIL.n436 185
R140 VTAIL.n435 VTAIL.n434 185
R141 VTAIL.n384 VTAIL.n383 185
R142 VTAIL.n429 VTAIL.n428 185
R143 VTAIL.n427 VTAIL.n426 185
R144 VTAIL.n388 VTAIL.n387 185
R145 VTAIL.n392 VTAIL.n390 185
R146 VTAIL.n421 VTAIL.n420 185
R147 VTAIL.n419 VTAIL.n418 185
R148 VTAIL.n394 VTAIL.n393 185
R149 VTAIL.n413 VTAIL.n412 185
R150 VTAIL.n411 VTAIL.n410 185
R151 VTAIL.n398 VTAIL.n397 185
R152 VTAIL.n405 VTAIL.n404 185
R153 VTAIL.n403 VTAIL.n402 185
R154 VTAIL.n373 VTAIL.n372 185
R155 VTAIL.n371 VTAIL.n370 185
R156 VTAIL.n320 VTAIL.n319 185
R157 VTAIL.n365 VTAIL.n364 185
R158 VTAIL.n363 VTAIL.n362 185
R159 VTAIL.n324 VTAIL.n323 185
R160 VTAIL.n328 VTAIL.n326 185
R161 VTAIL.n357 VTAIL.n356 185
R162 VTAIL.n355 VTAIL.n354 185
R163 VTAIL.n330 VTAIL.n329 185
R164 VTAIL.n349 VTAIL.n348 185
R165 VTAIL.n347 VTAIL.n346 185
R166 VTAIL.n334 VTAIL.n333 185
R167 VTAIL.n341 VTAIL.n340 185
R168 VTAIL.n339 VTAIL.n338 185
R169 VTAIL.n311 VTAIL.n310 185
R170 VTAIL.n309 VTAIL.n308 185
R171 VTAIL.n258 VTAIL.n257 185
R172 VTAIL.n303 VTAIL.n302 185
R173 VTAIL.n301 VTAIL.n300 185
R174 VTAIL.n262 VTAIL.n261 185
R175 VTAIL.n266 VTAIL.n264 185
R176 VTAIL.n295 VTAIL.n294 185
R177 VTAIL.n293 VTAIL.n292 185
R178 VTAIL.n268 VTAIL.n267 185
R179 VTAIL.n287 VTAIL.n286 185
R180 VTAIL.n285 VTAIL.n284 185
R181 VTAIL.n272 VTAIL.n271 185
R182 VTAIL.n279 VTAIL.n278 185
R183 VTAIL.n277 VTAIL.n276 185
R184 VTAIL.n247 VTAIL.n246 185
R185 VTAIL.n245 VTAIL.n244 185
R186 VTAIL.n194 VTAIL.n193 185
R187 VTAIL.n239 VTAIL.n238 185
R188 VTAIL.n237 VTAIL.n236 185
R189 VTAIL.n198 VTAIL.n197 185
R190 VTAIL.n202 VTAIL.n200 185
R191 VTAIL.n231 VTAIL.n230 185
R192 VTAIL.n229 VTAIL.n228 185
R193 VTAIL.n204 VTAIL.n203 185
R194 VTAIL.n223 VTAIL.n222 185
R195 VTAIL.n221 VTAIL.n220 185
R196 VTAIL.n208 VTAIL.n207 185
R197 VTAIL.n215 VTAIL.n214 185
R198 VTAIL.n213 VTAIL.n212 185
R199 VTAIL.n461 VTAIL.t6 149.524
R200 VTAIL.n21 VTAIL.t3 149.524
R201 VTAIL.n83 VTAIL.t10 149.524
R202 VTAIL.n147 VTAIL.t9 149.524
R203 VTAIL.n401 VTAIL.t7 149.524
R204 VTAIL.n337 VTAIL.t8 149.524
R205 VTAIL.n275 VTAIL.t1 149.524
R206 VTAIL.n211 VTAIL.t0 149.524
R207 VTAIL.n464 VTAIL.n463 104.615
R208 VTAIL.n464 VTAIL.n457 104.615
R209 VTAIL.n471 VTAIL.n457 104.615
R210 VTAIL.n472 VTAIL.n471 104.615
R211 VTAIL.n472 VTAIL.n453 104.615
R212 VTAIL.n480 VTAIL.n453 104.615
R213 VTAIL.n481 VTAIL.n480 104.615
R214 VTAIL.n482 VTAIL.n481 104.615
R215 VTAIL.n482 VTAIL.n449 104.615
R216 VTAIL.n489 VTAIL.n449 104.615
R217 VTAIL.n490 VTAIL.n489 104.615
R218 VTAIL.n490 VTAIL.n445 104.615
R219 VTAIL.n497 VTAIL.n445 104.615
R220 VTAIL.n498 VTAIL.n497 104.615
R221 VTAIL.n24 VTAIL.n23 104.615
R222 VTAIL.n24 VTAIL.n17 104.615
R223 VTAIL.n31 VTAIL.n17 104.615
R224 VTAIL.n32 VTAIL.n31 104.615
R225 VTAIL.n32 VTAIL.n13 104.615
R226 VTAIL.n40 VTAIL.n13 104.615
R227 VTAIL.n41 VTAIL.n40 104.615
R228 VTAIL.n42 VTAIL.n41 104.615
R229 VTAIL.n42 VTAIL.n9 104.615
R230 VTAIL.n49 VTAIL.n9 104.615
R231 VTAIL.n50 VTAIL.n49 104.615
R232 VTAIL.n50 VTAIL.n5 104.615
R233 VTAIL.n57 VTAIL.n5 104.615
R234 VTAIL.n58 VTAIL.n57 104.615
R235 VTAIL.n86 VTAIL.n85 104.615
R236 VTAIL.n86 VTAIL.n79 104.615
R237 VTAIL.n93 VTAIL.n79 104.615
R238 VTAIL.n94 VTAIL.n93 104.615
R239 VTAIL.n94 VTAIL.n75 104.615
R240 VTAIL.n102 VTAIL.n75 104.615
R241 VTAIL.n103 VTAIL.n102 104.615
R242 VTAIL.n104 VTAIL.n103 104.615
R243 VTAIL.n104 VTAIL.n71 104.615
R244 VTAIL.n111 VTAIL.n71 104.615
R245 VTAIL.n112 VTAIL.n111 104.615
R246 VTAIL.n112 VTAIL.n67 104.615
R247 VTAIL.n119 VTAIL.n67 104.615
R248 VTAIL.n120 VTAIL.n119 104.615
R249 VTAIL.n150 VTAIL.n149 104.615
R250 VTAIL.n150 VTAIL.n143 104.615
R251 VTAIL.n157 VTAIL.n143 104.615
R252 VTAIL.n158 VTAIL.n157 104.615
R253 VTAIL.n158 VTAIL.n139 104.615
R254 VTAIL.n166 VTAIL.n139 104.615
R255 VTAIL.n167 VTAIL.n166 104.615
R256 VTAIL.n168 VTAIL.n167 104.615
R257 VTAIL.n168 VTAIL.n135 104.615
R258 VTAIL.n175 VTAIL.n135 104.615
R259 VTAIL.n176 VTAIL.n175 104.615
R260 VTAIL.n176 VTAIL.n131 104.615
R261 VTAIL.n183 VTAIL.n131 104.615
R262 VTAIL.n184 VTAIL.n183 104.615
R263 VTAIL.n436 VTAIL.n435 104.615
R264 VTAIL.n435 VTAIL.n383 104.615
R265 VTAIL.n428 VTAIL.n383 104.615
R266 VTAIL.n428 VTAIL.n427 104.615
R267 VTAIL.n427 VTAIL.n387 104.615
R268 VTAIL.n392 VTAIL.n387 104.615
R269 VTAIL.n420 VTAIL.n392 104.615
R270 VTAIL.n420 VTAIL.n419 104.615
R271 VTAIL.n419 VTAIL.n393 104.615
R272 VTAIL.n412 VTAIL.n393 104.615
R273 VTAIL.n412 VTAIL.n411 104.615
R274 VTAIL.n411 VTAIL.n397 104.615
R275 VTAIL.n404 VTAIL.n397 104.615
R276 VTAIL.n404 VTAIL.n403 104.615
R277 VTAIL.n372 VTAIL.n371 104.615
R278 VTAIL.n371 VTAIL.n319 104.615
R279 VTAIL.n364 VTAIL.n319 104.615
R280 VTAIL.n364 VTAIL.n363 104.615
R281 VTAIL.n363 VTAIL.n323 104.615
R282 VTAIL.n328 VTAIL.n323 104.615
R283 VTAIL.n356 VTAIL.n328 104.615
R284 VTAIL.n356 VTAIL.n355 104.615
R285 VTAIL.n355 VTAIL.n329 104.615
R286 VTAIL.n348 VTAIL.n329 104.615
R287 VTAIL.n348 VTAIL.n347 104.615
R288 VTAIL.n347 VTAIL.n333 104.615
R289 VTAIL.n340 VTAIL.n333 104.615
R290 VTAIL.n340 VTAIL.n339 104.615
R291 VTAIL.n310 VTAIL.n309 104.615
R292 VTAIL.n309 VTAIL.n257 104.615
R293 VTAIL.n302 VTAIL.n257 104.615
R294 VTAIL.n302 VTAIL.n301 104.615
R295 VTAIL.n301 VTAIL.n261 104.615
R296 VTAIL.n266 VTAIL.n261 104.615
R297 VTAIL.n294 VTAIL.n266 104.615
R298 VTAIL.n294 VTAIL.n293 104.615
R299 VTAIL.n293 VTAIL.n267 104.615
R300 VTAIL.n286 VTAIL.n267 104.615
R301 VTAIL.n286 VTAIL.n285 104.615
R302 VTAIL.n285 VTAIL.n271 104.615
R303 VTAIL.n278 VTAIL.n271 104.615
R304 VTAIL.n278 VTAIL.n277 104.615
R305 VTAIL.n246 VTAIL.n245 104.615
R306 VTAIL.n245 VTAIL.n193 104.615
R307 VTAIL.n238 VTAIL.n193 104.615
R308 VTAIL.n238 VTAIL.n237 104.615
R309 VTAIL.n237 VTAIL.n197 104.615
R310 VTAIL.n202 VTAIL.n197 104.615
R311 VTAIL.n230 VTAIL.n202 104.615
R312 VTAIL.n230 VTAIL.n229 104.615
R313 VTAIL.n229 VTAIL.n203 104.615
R314 VTAIL.n222 VTAIL.n203 104.615
R315 VTAIL.n222 VTAIL.n221 104.615
R316 VTAIL.n221 VTAIL.n207 104.615
R317 VTAIL.n214 VTAIL.n207 104.615
R318 VTAIL.n214 VTAIL.n213 104.615
R319 VTAIL.n463 VTAIL.t6 52.3082
R320 VTAIL.n23 VTAIL.t3 52.3082
R321 VTAIL.n85 VTAIL.t10 52.3082
R322 VTAIL.n149 VTAIL.t9 52.3082
R323 VTAIL.n403 VTAIL.t7 52.3082
R324 VTAIL.n339 VTAIL.t8 52.3082
R325 VTAIL.n277 VTAIL.t1 52.3082
R326 VTAIL.n213 VTAIL.t0 52.3082
R327 VTAIL.n379 VTAIL.n378 47.7384
R328 VTAIL.n253 VTAIL.n252 47.7384
R329 VTAIL.n1 VTAIL.n0 47.7382
R330 VTAIL.n127 VTAIL.n126 47.7382
R331 VTAIL.n503 VTAIL.n502 34.5126
R332 VTAIL.n63 VTAIL.n62 34.5126
R333 VTAIL.n125 VTAIL.n124 34.5126
R334 VTAIL.n189 VTAIL.n188 34.5126
R335 VTAIL.n441 VTAIL.n440 34.5126
R336 VTAIL.n377 VTAIL.n376 34.5126
R337 VTAIL.n315 VTAIL.n314 34.5126
R338 VTAIL.n251 VTAIL.n250 34.5126
R339 VTAIL.n503 VTAIL.n441 23.4617
R340 VTAIL.n251 VTAIL.n189 23.4617
R341 VTAIL.n483 VTAIL.n450 13.1884
R342 VTAIL.n43 VTAIL.n10 13.1884
R343 VTAIL.n105 VTAIL.n72 13.1884
R344 VTAIL.n169 VTAIL.n136 13.1884
R345 VTAIL.n390 VTAIL.n388 13.1884
R346 VTAIL.n326 VTAIL.n324 13.1884
R347 VTAIL.n264 VTAIL.n262 13.1884
R348 VTAIL.n200 VTAIL.n198 13.1884
R349 VTAIL.n484 VTAIL.n452 12.8005
R350 VTAIL.n488 VTAIL.n487 12.8005
R351 VTAIL.n44 VTAIL.n12 12.8005
R352 VTAIL.n48 VTAIL.n47 12.8005
R353 VTAIL.n106 VTAIL.n74 12.8005
R354 VTAIL.n110 VTAIL.n109 12.8005
R355 VTAIL.n170 VTAIL.n138 12.8005
R356 VTAIL.n174 VTAIL.n173 12.8005
R357 VTAIL.n426 VTAIL.n425 12.8005
R358 VTAIL.n422 VTAIL.n421 12.8005
R359 VTAIL.n362 VTAIL.n361 12.8005
R360 VTAIL.n358 VTAIL.n357 12.8005
R361 VTAIL.n300 VTAIL.n299 12.8005
R362 VTAIL.n296 VTAIL.n295 12.8005
R363 VTAIL.n236 VTAIL.n235 12.8005
R364 VTAIL.n232 VTAIL.n231 12.8005
R365 VTAIL.n479 VTAIL.n478 12.0247
R366 VTAIL.n491 VTAIL.n448 12.0247
R367 VTAIL.n39 VTAIL.n38 12.0247
R368 VTAIL.n51 VTAIL.n8 12.0247
R369 VTAIL.n101 VTAIL.n100 12.0247
R370 VTAIL.n113 VTAIL.n70 12.0247
R371 VTAIL.n165 VTAIL.n164 12.0247
R372 VTAIL.n177 VTAIL.n134 12.0247
R373 VTAIL.n429 VTAIL.n386 12.0247
R374 VTAIL.n418 VTAIL.n391 12.0247
R375 VTAIL.n365 VTAIL.n322 12.0247
R376 VTAIL.n354 VTAIL.n327 12.0247
R377 VTAIL.n303 VTAIL.n260 12.0247
R378 VTAIL.n292 VTAIL.n265 12.0247
R379 VTAIL.n239 VTAIL.n196 12.0247
R380 VTAIL.n228 VTAIL.n201 12.0247
R381 VTAIL.n477 VTAIL.n454 11.249
R382 VTAIL.n492 VTAIL.n446 11.249
R383 VTAIL.n37 VTAIL.n14 11.249
R384 VTAIL.n52 VTAIL.n6 11.249
R385 VTAIL.n99 VTAIL.n76 11.249
R386 VTAIL.n114 VTAIL.n68 11.249
R387 VTAIL.n163 VTAIL.n140 11.249
R388 VTAIL.n178 VTAIL.n132 11.249
R389 VTAIL.n430 VTAIL.n384 11.249
R390 VTAIL.n417 VTAIL.n394 11.249
R391 VTAIL.n366 VTAIL.n320 11.249
R392 VTAIL.n353 VTAIL.n330 11.249
R393 VTAIL.n304 VTAIL.n258 11.249
R394 VTAIL.n291 VTAIL.n268 11.249
R395 VTAIL.n240 VTAIL.n194 11.249
R396 VTAIL.n227 VTAIL.n204 11.249
R397 VTAIL.n474 VTAIL.n473 10.4732
R398 VTAIL.n496 VTAIL.n495 10.4732
R399 VTAIL.n34 VTAIL.n33 10.4732
R400 VTAIL.n56 VTAIL.n55 10.4732
R401 VTAIL.n96 VTAIL.n95 10.4732
R402 VTAIL.n118 VTAIL.n117 10.4732
R403 VTAIL.n160 VTAIL.n159 10.4732
R404 VTAIL.n182 VTAIL.n181 10.4732
R405 VTAIL.n434 VTAIL.n433 10.4732
R406 VTAIL.n414 VTAIL.n413 10.4732
R407 VTAIL.n370 VTAIL.n369 10.4732
R408 VTAIL.n350 VTAIL.n349 10.4732
R409 VTAIL.n308 VTAIL.n307 10.4732
R410 VTAIL.n288 VTAIL.n287 10.4732
R411 VTAIL.n244 VTAIL.n243 10.4732
R412 VTAIL.n224 VTAIL.n223 10.4732
R413 VTAIL.n462 VTAIL.n461 10.2747
R414 VTAIL.n22 VTAIL.n21 10.2747
R415 VTAIL.n84 VTAIL.n83 10.2747
R416 VTAIL.n148 VTAIL.n147 10.2747
R417 VTAIL.n402 VTAIL.n401 10.2747
R418 VTAIL.n338 VTAIL.n337 10.2747
R419 VTAIL.n276 VTAIL.n275 10.2747
R420 VTAIL.n212 VTAIL.n211 10.2747
R421 VTAIL.n470 VTAIL.n456 9.69747
R422 VTAIL.n499 VTAIL.n444 9.69747
R423 VTAIL.n30 VTAIL.n16 9.69747
R424 VTAIL.n59 VTAIL.n4 9.69747
R425 VTAIL.n92 VTAIL.n78 9.69747
R426 VTAIL.n121 VTAIL.n66 9.69747
R427 VTAIL.n156 VTAIL.n142 9.69747
R428 VTAIL.n185 VTAIL.n130 9.69747
R429 VTAIL.n437 VTAIL.n382 9.69747
R430 VTAIL.n410 VTAIL.n396 9.69747
R431 VTAIL.n373 VTAIL.n318 9.69747
R432 VTAIL.n346 VTAIL.n332 9.69747
R433 VTAIL.n311 VTAIL.n256 9.69747
R434 VTAIL.n284 VTAIL.n270 9.69747
R435 VTAIL.n247 VTAIL.n192 9.69747
R436 VTAIL.n220 VTAIL.n206 9.69747
R437 VTAIL.n502 VTAIL.n501 9.45567
R438 VTAIL.n62 VTAIL.n61 9.45567
R439 VTAIL.n124 VTAIL.n123 9.45567
R440 VTAIL.n188 VTAIL.n187 9.45567
R441 VTAIL.n440 VTAIL.n439 9.45567
R442 VTAIL.n376 VTAIL.n375 9.45567
R443 VTAIL.n314 VTAIL.n313 9.45567
R444 VTAIL.n250 VTAIL.n249 9.45567
R445 VTAIL.n501 VTAIL.n500 9.3005
R446 VTAIL.n444 VTAIL.n443 9.3005
R447 VTAIL.n495 VTAIL.n494 9.3005
R448 VTAIL.n493 VTAIL.n492 9.3005
R449 VTAIL.n448 VTAIL.n447 9.3005
R450 VTAIL.n487 VTAIL.n486 9.3005
R451 VTAIL.n460 VTAIL.n459 9.3005
R452 VTAIL.n467 VTAIL.n466 9.3005
R453 VTAIL.n469 VTAIL.n468 9.3005
R454 VTAIL.n456 VTAIL.n455 9.3005
R455 VTAIL.n475 VTAIL.n474 9.3005
R456 VTAIL.n477 VTAIL.n476 9.3005
R457 VTAIL.n478 VTAIL.n451 9.3005
R458 VTAIL.n485 VTAIL.n484 9.3005
R459 VTAIL.n61 VTAIL.n60 9.3005
R460 VTAIL.n4 VTAIL.n3 9.3005
R461 VTAIL.n55 VTAIL.n54 9.3005
R462 VTAIL.n53 VTAIL.n52 9.3005
R463 VTAIL.n8 VTAIL.n7 9.3005
R464 VTAIL.n47 VTAIL.n46 9.3005
R465 VTAIL.n20 VTAIL.n19 9.3005
R466 VTAIL.n27 VTAIL.n26 9.3005
R467 VTAIL.n29 VTAIL.n28 9.3005
R468 VTAIL.n16 VTAIL.n15 9.3005
R469 VTAIL.n35 VTAIL.n34 9.3005
R470 VTAIL.n37 VTAIL.n36 9.3005
R471 VTAIL.n38 VTAIL.n11 9.3005
R472 VTAIL.n45 VTAIL.n44 9.3005
R473 VTAIL.n123 VTAIL.n122 9.3005
R474 VTAIL.n66 VTAIL.n65 9.3005
R475 VTAIL.n117 VTAIL.n116 9.3005
R476 VTAIL.n115 VTAIL.n114 9.3005
R477 VTAIL.n70 VTAIL.n69 9.3005
R478 VTAIL.n109 VTAIL.n108 9.3005
R479 VTAIL.n82 VTAIL.n81 9.3005
R480 VTAIL.n89 VTAIL.n88 9.3005
R481 VTAIL.n91 VTAIL.n90 9.3005
R482 VTAIL.n78 VTAIL.n77 9.3005
R483 VTAIL.n97 VTAIL.n96 9.3005
R484 VTAIL.n99 VTAIL.n98 9.3005
R485 VTAIL.n100 VTAIL.n73 9.3005
R486 VTAIL.n107 VTAIL.n106 9.3005
R487 VTAIL.n187 VTAIL.n186 9.3005
R488 VTAIL.n130 VTAIL.n129 9.3005
R489 VTAIL.n181 VTAIL.n180 9.3005
R490 VTAIL.n179 VTAIL.n178 9.3005
R491 VTAIL.n134 VTAIL.n133 9.3005
R492 VTAIL.n173 VTAIL.n172 9.3005
R493 VTAIL.n146 VTAIL.n145 9.3005
R494 VTAIL.n153 VTAIL.n152 9.3005
R495 VTAIL.n155 VTAIL.n154 9.3005
R496 VTAIL.n142 VTAIL.n141 9.3005
R497 VTAIL.n161 VTAIL.n160 9.3005
R498 VTAIL.n163 VTAIL.n162 9.3005
R499 VTAIL.n164 VTAIL.n137 9.3005
R500 VTAIL.n171 VTAIL.n170 9.3005
R501 VTAIL.n400 VTAIL.n399 9.3005
R502 VTAIL.n407 VTAIL.n406 9.3005
R503 VTAIL.n409 VTAIL.n408 9.3005
R504 VTAIL.n396 VTAIL.n395 9.3005
R505 VTAIL.n415 VTAIL.n414 9.3005
R506 VTAIL.n417 VTAIL.n416 9.3005
R507 VTAIL.n391 VTAIL.n389 9.3005
R508 VTAIL.n423 VTAIL.n422 9.3005
R509 VTAIL.n439 VTAIL.n438 9.3005
R510 VTAIL.n382 VTAIL.n381 9.3005
R511 VTAIL.n433 VTAIL.n432 9.3005
R512 VTAIL.n431 VTAIL.n430 9.3005
R513 VTAIL.n386 VTAIL.n385 9.3005
R514 VTAIL.n425 VTAIL.n424 9.3005
R515 VTAIL.n336 VTAIL.n335 9.3005
R516 VTAIL.n343 VTAIL.n342 9.3005
R517 VTAIL.n345 VTAIL.n344 9.3005
R518 VTAIL.n332 VTAIL.n331 9.3005
R519 VTAIL.n351 VTAIL.n350 9.3005
R520 VTAIL.n353 VTAIL.n352 9.3005
R521 VTAIL.n327 VTAIL.n325 9.3005
R522 VTAIL.n359 VTAIL.n358 9.3005
R523 VTAIL.n375 VTAIL.n374 9.3005
R524 VTAIL.n318 VTAIL.n317 9.3005
R525 VTAIL.n369 VTAIL.n368 9.3005
R526 VTAIL.n367 VTAIL.n366 9.3005
R527 VTAIL.n322 VTAIL.n321 9.3005
R528 VTAIL.n361 VTAIL.n360 9.3005
R529 VTAIL.n274 VTAIL.n273 9.3005
R530 VTAIL.n281 VTAIL.n280 9.3005
R531 VTAIL.n283 VTAIL.n282 9.3005
R532 VTAIL.n270 VTAIL.n269 9.3005
R533 VTAIL.n289 VTAIL.n288 9.3005
R534 VTAIL.n291 VTAIL.n290 9.3005
R535 VTAIL.n265 VTAIL.n263 9.3005
R536 VTAIL.n297 VTAIL.n296 9.3005
R537 VTAIL.n313 VTAIL.n312 9.3005
R538 VTAIL.n256 VTAIL.n255 9.3005
R539 VTAIL.n307 VTAIL.n306 9.3005
R540 VTAIL.n305 VTAIL.n304 9.3005
R541 VTAIL.n260 VTAIL.n259 9.3005
R542 VTAIL.n299 VTAIL.n298 9.3005
R543 VTAIL.n210 VTAIL.n209 9.3005
R544 VTAIL.n217 VTAIL.n216 9.3005
R545 VTAIL.n219 VTAIL.n218 9.3005
R546 VTAIL.n206 VTAIL.n205 9.3005
R547 VTAIL.n225 VTAIL.n224 9.3005
R548 VTAIL.n227 VTAIL.n226 9.3005
R549 VTAIL.n201 VTAIL.n199 9.3005
R550 VTAIL.n233 VTAIL.n232 9.3005
R551 VTAIL.n249 VTAIL.n248 9.3005
R552 VTAIL.n192 VTAIL.n191 9.3005
R553 VTAIL.n243 VTAIL.n242 9.3005
R554 VTAIL.n241 VTAIL.n240 9.3005
R555 VTAIL.n196 VTAIL.n195 9.3005
R556 VTAIL.n235 VTAIL.n234 9.3005
R557 VTAIL.n469 VTAIL.n458 8.92171
R558 VTAIL.n500 VTAIL.n442 8.92171
R559 VTAIL.n29 VTAIL.n18 8.92171
R560 VTAIL.n60 VTAIL.n2 8.92171
R561 VTAIL.n91 VTAIL.n80 8.92171
R562 VTAIL.n122 VTAIL.n64 8.92171
R563 VTAIL.n155 VTAIL.n144 8.92171
R564 VTAIL.n186 VTAIL.n128 8.92171
R565 VTAIL.n438 VTAIL.n380 8.92171
R566 VTAIL.n409 VTAIL.n398 8.92171
R567 VTAIL.n374 VTAIL.n316 8.92171
R568 VTAIL.n345 VTAIL.n334 8.92171
R569 VTAIL.n312 VTAIL.n254 8.92171
R570 VTAIL.n283 VTAIL.n272 8.92171
R571 VTAIL.n248 VTAIL.n190 8.92171
R572 VTAIL.n219 VTAIL.n208 8.92171
R573 VTAIL.n466 VTAIL.n465 8.14595
R574 VTAIL.n26 VTAIL.n25 8.14595
R575 VTAIL.n88 VTAIL.n87 8.14595
R576 VTAIL.n152 VTAIL.n151 8.14595
R577 VTAIL.n406 VTAIL.n405 8.14595
R578 VTAIL.n342 VTAIL.n341 8.14595
R579 VTAIL.n280 VTAIL.n279 8.14595
R580 VTAIL.n216 VTAIL.n215 8.14595
R581 VTAIL.n462 VTAIL.n460 7.3702
R582 VTAIL.n22 VTAIL.n20 7.3702
R583 VTAIL.n84 VTAIL.n82 7.3702
R584 VTAIL.n148 VTAIL.n146 7.3702
R585 VTAIL.n402 VTAIL.n400 7.3702
R586 VTAIL.n338 VTAIL.n336 7.3702
R587 VTAIL.n276 VTAIL.n274 7.3702
R588 VTAIL.n212 VTAIL.n210 7.3702
R589 VTAIL.n465 VTAIL.n460 5.81868
R590 VTAIL.n25 VTAIL.n20 5.81868
R591 VTAIL.n87 VTAIL.n82 5.81868
R592 VTAIL.n151 VTAIL.n146 5.81868
R593 VTAIL.n405 VTAIL.n400 5.81868
R594 VTAIL.n341 VTAIL.n336 5.81868
R595 VTAIL.n279 VTAIL.n274 5.81868
R596 VTAIL.n215 VTAIL.n210 5.81868
R597 VTAIL.n466 VTAIL.n458 5.04292
R598 VTAIL.n502 VTAIL.n442 5.04292
R599 VTAIL.n26 VTAIL.n18 5.04292
R600 VTAIL.n62 VTAIL.n2 5.04292
R601 VTAIL.n88 VTAIL.n80 5.04292
R602 VTAIL.n124 VTAIL.n64 5.04292
R603 VTAIL.n152 VTAIL.n144 5.04292
R604 VTAIL.n188 VTAIL.n128 5.04292
R605 VTAIL.n440 VTAIL.n380 5.04292
R606 VTAIL.n406 VTAIL.n398 5.04292
R607 VTAIL.n376 VTAIL.n316 5.04292
R608 VTAIL.n342 VTAIL.n334 5.04292
R609 VTAIL.n314 VTAIL.n254 5.04292
R610 VTAIL.n280 VTAIL.n272 5.04292
R611 VTAIL.n250 VTAIL.n190 5.04292
R612 VTAIL.n216 VTAIL.n208 5.04292
R613 VTAIL.n470 VTAIL.n469 4.26717
R614 VTAIL.n500 VTAIL.n499 4.26717
R615 VTAIL.n30 VTAIL.n29 4.26717
R616 VTAIL.n60 VTAIL.n59 4.26717
R617 VTAIL.n92 VTAIL.n91 4.26717
R618 VTAIL.n122 VTAIL.n121 4.26717
R619 VTAIL.n156 VTAIL.n155 4.26717
R620 VTAIL.n186 VTAIL.n185 4.26717
R621 VTAIL.n438 VTAIL.n437 4.26717
R622 VTAIL.n410 VTAIL.n409 4.26717
R623 VTAIL.n374 VTAIL.n373 4.26717
R624 VTAIL.n346 VTAIL.n345 4.26717
R625 VTAIL.n312 VTAIL.n311 4.26717
R626 VTAIL.n284 VTAIL.n283 4.26717
R627 VTAIL.n248 VTAIL.n247 4.26717
R628 VTAIL.n220 VTAIL.n219 4.26717
R629 VTAIL.n473 VTAIL.n456 3.49141
R630 VTAIL.n496 VTAIL.n444 3.49141
R631 VTAIL.n33 VTAIL.n16 3.49141
R632 VTAIL.n56 VTAIL.n4 3.49141
R633 VTAIL.n95 VTAIL.n78 3.49141
R634 VTAIL.n118 VTAIL.n66 3.49141
R635 VTAIL.n159 VTAIL.n142 3.49141
R636 VTAIL.n182 VTAIL.n130 3.49141
R637 VTAIL.n434 VTAIL.n382 3.49141
R638 VTAIL.n413 VTAIL.n396 3.49141
R639 VTAIL.n370 VTAIL.n318 3.49141
R640 VTAIL.n349 VTAIL.n332 3.49141
R641 VTAIL.n308 VTAIL.n256 3.49141
R642 VTAIL.n287 VTAIL.n270 3.49141
R643 VTAIL.n244 VTAIL.n192 3.49141
R644 VTAIL.n223 VTAIL.n206 3.49141
R645 VTAIL.n461 VTAIL.n459 2.84303
R646 VTAIL.n21 VTAIL.n19 2.84303
R647 VTAIL.n83 VTAIL.n81 2.84303
R648 VTAIL.n147 VTAIL.n145 2.84303
R649 VTAIL.n401 VTAIL.n399 2.84303
R650 VTAIL.n337 VTAIL.n335 2.84303
R651 VTAIL.n275 VTAIL.n273 2.84303
R652 VTAIL.n211 VTAIL.n209 2.84303
R653 VTAIL.n474 VTAIL.n454 2.71565
R654 VTAIL.n495 VTAIL.n446 2.71565
R655 VTAIL.n34 VTAIL.n14 2.71565
R656 VTAIL.n55 VTAIL.n6 2.71565
R657 VTAIL.n96 VTAIL.n76 2.71565
R658 VTAIL.n117 VTAIL.n68 2.71565
R659 VTAIL.n160 VTAIL.n140 2.71565
R660 VTAIL.n181 VTAIL.n132 2.71565
R661 VTAIL.n433 VTAIL.n384 2.71565
R662 VTAIL.n414 VTAIL.n394 2.71565
R663 VTAIL.n369 VTAIL.n320 2.71565
R664 VTAIL.n350 VTAIL.n330 2.71565
R665 VTAIL.n307 VTAIL.n258 2.71565
R666 VTAIL.n288 VTAIL.n268 2.71565
R667 VTAIL.n243 VTAIL.n194 2.71565
R668 VTAIL.n224 VTAIL.n204 2.71565
R669 VTAIL.n479 VTAIL.n477 1.93989
R670 VTAIL.n492 VTAIL.n491 1.93989
R671 VTAIL.n39 VTAIL.n37 1.93989
R672 VTAIL.n52 VTAIL.n51 1.93989
R673 VTAIL.n101 VTAIL.n99 1.93989
R674 VTAIL.n114 VTAIL.n113 1.93989
R675 VTAIL.n165 VTAIL.n163 1.93989
R676 VTAIL.n178 VTAIL.n177 1.93989
R677 VTAIL.n430 VTAIL.n429 1.93989
R678 VTAIL.n418 VTAIL.n417 1.93989
R679 VTAIL.n366 VTAIL.n365 1.93989
R680 VTAIL.n354 VTAIL.n353 1.93989
R681 VTAIL.n304 VTAIL.n303 1.93989
R682 VTAIL.n292 VTAIL.n291 1.93989
R683 VTAIL.n240 VTAIL.n239 1.93989
R684 VTAIL.n228 VTAIL.n227 1.93989
R685 VTAIL.n0 VTAIL.t4 1.71925
R686 VTAIL.n0 VTAIL.t5 1.71925
R687 VTAIL.n126 VTAIL.t12 1.71925
R688 VTAIL.n126 VTAIL.t14 1.71925
R689 VTAIL.n378 VTAIL.t11 1.71925
R690 VTAIL.n378 VTAIL.t13 1.71925
R691 VTAIL.n252 VTAIL.t15 1.71925
R692 VTAIL.n252 VTAIL.t2 1.71925
R693 VTAIL.n253 VTAIL.n251 1.16429
R694 VTAIL.n315 VTAIL.n253 1.16429
R695 VTAIL.n379 VTAIL.n377 1.16429
R696 VTAIL.n441 VTAIL.n379 1.16429
R697 VTAIL.n189 VTAIL.n127 1.16429
R698 VTAIL.n127 VTAIL.n125 1.16429
R699 VTAIL.n63 VTAIL.n1 1.16429
R700 VTAIL.n478 VTAIL.n452 1.16414
R701 VTAIL.n488 VTAIL.n448 1.16414
R702 VTAIL.n38 VTAIL.n12 1.16414
R703 VTAIL.n48 VTAIL.n8 1.16414
R704 VTAIL.n100 VTAIL.n74 1.16414
R705 VTAIL.n110 VTAIL.n70 1.16414
R706 VTAIL.n164 VTAIL.n138 1.16414
R707 VTAIL.n174 VTAIL.n134 1.16414
R708 VTAIL.n426 VTAIL.n386 1.16414
R709 VTAIL.n421 VTAIL.n391 1.16414
R710 VTAIL.n362 VTAIL.n322 1.16414
R711 VTAIL.n357 VTAIL.n327 1.16414
R712 VTAIL.n300 VTAIL.n260 1.16414
R713 VTAIL.n295 VTAIL.n265 1.16414
R714 VTAIL.n236 VTAIL.n196 1.16414
R715 VTAIL.n231 VTAIL.n201 1.16414
R716 VTAIL VTAIL.n503 1.1061
R717 VTAIL.n377 VTAIL.n315 0.470328
R718 VTAIL.n125 VTAIL.n63 0.470328
R719 VTAIL.n484 VTAIL.n483 0.388379
R720 VTAIL.n487 VTAIL.n450 0.388379
R721 VTAIL.n44 VTAIL.n43 0.388379
R722 VTAIL.n47 VTAIL.n10 0.388379
R723 VTAIL.n106 VTAIL.n105 0.388379
R724 VTAIL.n109 VTAIL.n72 0.388379
R725 VTAIL.n170 VTAIL.n169 0.388379
R726 VTAIL.n173 VTAIL.n136 0.388379
R727 VTAIL.n425 VTAIL.n388 0.388379
R728 VTAIL.n422 VTAIL.n390 0.388379
R729 VTAIL.n361 VTAIL.n324 0.388379
R730 VTAIL.n358 VTAIL.n326 0.388379
R731 VTAIL.n299 VTAIL.n262 0.388379
R732 VTAIL.n296 VTAIL.n264 0.388379
R733 VTAIL.n235 VTAIL.n198 0.388379
R734 VTAIL.n232 VTAIL.n200 0.388379
R735 VTAIL.n467 VTAIL.n459 0.155672
R736 VTAIL.n468 VTAIL.n467 0.155672
R737 VTAIL.n468 VTAIL.n455 0.155672
R738 VTAIL.n475 VTAIL.n455 0.155672
R739 VTAIL.n476 VTAIL.n475 0.155672
R740 VTAIL.n476 VTAIL.n451 0.155672
R741 VTAIL.n485 VTAIL.n451 0.155672
R742 VTAIL.n486 VTAIL.n485 0.155672
R743 VTAIL.n486 VTAIL.n447 0.155672
R744 VTAIL.n493 VTAIL.n447 0.155672
R745 VTAIL.n494 VTAIL.n493 0.155672
R746 VTAIL.n494 VTAIL.n443 0.155672
R747 VTAIL.n501 VTAIL.n443 0.155672
R748 VTAIL.n27 VTAIL.n19 0.155672
R749 VTAIL.n28 VTAIL.n27 0.155672
R750 VTAIL.n28 VTAIL.n15 0.155672
R751 VTAIL.n35 VTAIL.n15 0.155672
R752 VTAIL.n36 VTAIL.n35 0.155672
R753 VTAIL.n36 VTAIL.n11 0.155672
R754 VTAIL.n45 VTAIL.n11 0.155672
R755 VTAIL.n46 VTAIL.n45 0.155672
R756 VTAIL.n46 VTAIL.n7 0.155672
R757 VTAIL.n53 VTAIL.n7 0.155672
R758 VTAIL.n54 VTAIL.n53 0.155672
R759 VTAIL.n54 VTAIL.n3 0.155672
R760 VTAIL.n61 VTAIL.n3 0.155672
R761 VTAIL.n89 VTAIL.n81 0.155672
R762 VTAIL.n90 VTAIL.n89 0.155672
R763 VTAIL.n90 VTAIL.n77 0.155672
R764 VTAIL.n97 VTAIL.n77 0.155672
R765 VTAIL.n98 VTAIL.n97 0.155672
R766 VTAIL.n98 VTAIL.n73 0.155672
R767 VTAIL.n107 VTAIL.n73 0.155672
R768 VTAIL.n108 VTAIL.n107 0.155672
R769 VTAIL.n108 VTAIL.n69 0.155672
R770 VTAIL.n115 VTAIL.n69 0.155672
R771 VTAIL.n116 VTAIL.n115 0.155672
R772 VTAIL.n116 VTAIL.n65 0.155672
R773 VTAIL.n123 VTAIL.n65 0.155672
R774 VTAIL.n153 VTAIL.n145 0.155672
R775 VTAIL.n154 VTAIL.n153 0.155672
R776 VTAIL.n154 VTAIL.n141 0.155672
R777 VTAIL.n161 VTAIL.n141 0.155672
R778 VTAIL.n162 VTAIL.n161 0.155672
R779 VTAIL.n162 VTAIL.n137 0.155672
R780 VTAIL.n171 VTAIL.n137 0.155672
R781 VTAIL.n172 VTAIL.n171 0.155672
R782 VTAIL.n172 VTAIL.n133 0.155672
R783 VTAIL.n179 VTAIL.n133 0.155672
R784 VTAIL.n180 VTAIL.n179 0.155672
R785 VTAIL.n180 VTAIL.n129 0.155672
R786 VTAIL.n187 VTAIL.n129 0.155672
R787 VTAIL.n439 VTAIL.n381 0.155672
R788 VTAIL.n432 VTAIL.n381 0.155672
R789 VTAIL.n432 VTAIL.n431 0.155672
R790 VTAIL.n431 VTAIL.n385 0.155672
R791 VTAIL.n424 VTAIL.n385 0.155672
R792 VTAIL.n424 VTAIL.n423 0.155672
R793 VTAIL.n423 VTAIL.n389 0.155672
R794 VTAIL.n416 VTAIL.n389 0.155672
R795 VTAIL.n416 VTAIL.n415 0.155672
R796 VTAIL.n415 VTAIL.n395 0.155672
R797 VTAIL.n408 VTAIL.n395 0.155672
R798 VTAIL.n408 VTAIL.n407 0.155672
R799 VTAIL.n407 VTAIL.n399 0.155672
R800 VTAIL.n375 VTAIL.n317 0.155672
R801 VTAIL.n368 VTAIL.n317 0.155672
R802 VTAIL.n368 VTAIL.n367 0.155672
R803 VTAIL.n367 VTAIL.n321 0.155672
R804 VTAIL.n360 VTAIL.n321 0.155672
R805 VTAIL.n360 VTAIL.n359 0.155672
R806 VTAIL.n359 VTAIL.n325 0.155672
R807 VTAIL.n352 VTAIL.n325 0.155672
R808 VTAIL.n352 VTAIL.n351 0.155672
R809 VTAIL.n351 VTAIL.n331 0.155672
R810 VTAIL.n344 VTAIL.n331 0.155672
R811 VTAIL.n344 VTAIL.n343 0.155672
R812 VTAIL.n343 VTAIL.n335 0.155672
R813 VTAIL.n313 VTAIL.n255 0.155672
R814 VTAIL.n306 VTAIL.n255 0.155672
R815 VTAIL.n306 VTAIL.n305 0.155672
R816 VTAIL.n305 VTAIL.n259 0.155672
R817 VTAIL.n298 VTAIL.n259 0.155672
R818 VTAIL.n298 VTAIL.n297 0.155672
R819 VTAIL.n297 VTAIL.n263 0.155672
R820 VTAIL.n290 VTAIL.n263 0.155672
R821 VTAIL.n290 VTAIL.n289 0.155672
R822 VTAIL.n289 VTAIL.n269 0.155672
R823 VTAIL.n282 VTAIL.n269 0.155672
R824 VTAIL.n282 VTAIL.n281 0.155672
R825 VTAIL.n281 VTAIL.n273 0.155672
R826 VTAIL.n249 VTAIL.n191 0.155672
R827 VTAIL.n242 VTAIL.n191 0.155672
R828 VTAIL.n242 VTAIL.n241 0.155672
R829 VTAIL.n241 VTAIL.n195 0.155672
R830 VTAIL.n234 VTAIL.n195 0.155672
R831 VTAIL.n234 VTAIL.n233 0.155672
R832 VTAIL.n233 VTAIL.n199 0.155672
R833 VTAIL.n226 VTAIL.n199 0.155672
R834 VTAIL.n226 VTAIL.n225 0.155672
R835 VTAIL.n225 VTAIL.n205 0.155672
R836 VTAIL.n218 VTAIL.n205 0.155672
R837 VTAIL.n218 VTAIL.n217 0.155672
R838 VTAIL.n217 VTAIL.n209 0.155672
R839 VTAIL VTAIL.n1 0.0586897
R840 B.n686 B.n685 585
R841 B.n280 B.n99 585
R842 B.n279 B.n278 585
R843 B.n277 B.n276 585
R844 B.n275 B.n274 585
R845 B.n273 B.n272 585
R846 B.n271 B.n270 585
R847 B.n269 B.n268 585
R848 B.n267 B.n266 585
R849 B.n265 B.n264 585
R850 B.n263 B.n262 585
R851 B.n261 B.n260 585
R852 B.n259 B.n258 585
R853 B.n257 B.n256 585
R854 B.n255 B.n254 585
R855 B.n253 B.n252 585
R856 B.n251 B.n250 585
R857 B.n249 B.n248 585
R858 B.n247 B.n246 585
R859 B.n245 B.n244 585
R860 B.n243 B.n242 585
R861 B.n241 B.n240 585
R862 B.n239 B.n238 585
R863 B.n237 B.n236 585
R864 B.n235 B.n234 585
R865 B.n233 B.n232 585
R866 B.n231 B.n230 585
R867 B.n229 B.n228 585
R868 B.n227 B.n226 585
R869 B.n225 B.n224 585
R870 B.n223 B.n222 585
R871 B.n221 B.n220 585
R872 B.n219 B.n218 585
R873 B.n217 B.n216 585
R874 B.n215 B.n214 585
R875 B.n213 B.n212 585
R876 B.n211 B.n210 585
R877 B.n209 B.n208 585
R878 B.n207 B.n206 585
R879 B.n205 B.n204 585
R880 B.n203 B.n202 585
R881 B.n201 B.n200 585
R882 B.n199 B.n198 585
R883 B.n197 B.n196 585
R884 B.n195 B.n194 585
R885 B.n193 B.n192 585
R886 B.n191 B.n190 585
R887 B.n189 B.n188 585
R888 B.n187 B.n186 585
R889 B.n185 B.n184 585
R890 B.n183 B.n182 585
R891 B.n181 B.n180 585
R892 B.n179 B.n178 585
R893 B.n177 B.n176 585
R894 B.n175 B.n174 585
R895 B.n173 B.n172 585
R896 B.n171 B.n170 585
R897 B.n169 B.n168 585
R898 B.n167 B.n166 585
R899 B.n165 B.n164 585
R900 B.n163 B.n162 585
R901 B.n161 B.n160 585
R902 B.n159 B.n158 585
R903 B.n157 B.n156 585
R904 B.n155 B.n154 585
R905 B.n153 B.n152 585
R906 B.n151 B.n150 585
R907 B.n149 B.n148 585
R908 B.n147 B.n146 585
R909 B.n145 B.n144 585
R910 B.n143 B.n142 585
R911 B.n141 B.n140 585
R912 B.n139 B.n138 585
R913 B.n137 B.n136 585
R914 B.n135 B.n134 585
R915 B.n133 B.n132 585
R916 B.n131 B.n130 585
R917 B.n129 B.n128 585
R918 B.n127 B.n126 585
R919 B.n125 B.n124 585
R920 B.n123 B.n122 585
R921 B.n121 B.n120 585
R922 B.n119 B.n118 585
R923 B.n117 B.n116 585
R924 B.n115 B.n114 585
R925 B.n113 B.n112 585
R926 B.n111 B.n110 585
R927 B.n109 B.n108 585
R928 B.n107 B.n106 585
R929 B.n53 B.n52 585
R930 B.n684 B.n54 585
R931 B.n689 B.n54 585
R932 B.n683 B.n682 585
R933 B.n682 B.n50 585
R934 B.n681 B.n49 585
R935 B.n695 B.n49 585
R936 B.n680 B.n48 585
R937 B.n696 B.n48 585
R938 B.n679 B.n47 585
R939 B.n697 B.n47 585
R940 B.n678 B.n677 585
R941 B.n677 B.n46 585
R942 B.n676 B.n42 585
R943 B.n703 B.n42 585
R944 B.n675 B.n41 585
R945 B.n704 B.n41 585
R946 B.n674 B.n40 585
R947 B.n705 B.n40 585
R948 B.n673 B.n672 585
R949 B.n672 B.n36 585
R950 B.n671 B.n35 585
R951 B.n711 B.n35 585
R952 B.n670 B.n34 585
R953 B.n712 B.n34 585
R954 B.n669 B.n33 585
R955 B.n713 B.n33 585
R956 B.n668 B.n667 585
R957 B.n667 B.n29 585
R958 B.n666 B.n28 585
R959 B.n719 B.n28 585
R960 B.n665 B.n27 585
R961 B.n720 B.n27 585
R962 B.n664 B.n26 585
R963 B.n721 B.n26 585
R964 B.n663 B.n662 585
R965 B.n662 B.n22 585
R966 B.n661 B.n21 585
R967 B.n727 B.n21 585
R968 B.n660 B.n20 585
R969 B.n728 B.n20 585
R970 B.n659 B.n19 585
R971 B.n729 B.n19 585
R972 B.n658 B.n657 585
R973 B.n657 B.n15 585
R974 B.n656 B.n14 585
R975 B.n735 B.n14 585
R976 B.n655 B.n13 585
R977 B.n736 B.n13 585
R978 B.n654 B.n12 585
R979 B.n737 B.n12 585
R980 B.n653 B.n652 585
R981 B.n652 B.n8 585
R982 B.n651 B.n7 585
R983 B.n743 B.n7 585
R984 B.n650 B.n6 585
R985 B.n744 B.n6 585
R986 B.n649 B.n5 585
R987 B.n745 B.n5 585
R988 B.n648 B.n647 585
R989 B.n647 B.n4 585
R990 B.n646 B.n281 585
R991 B.n646 B.n645 585
R992 B.n636 B.n282 585
R993 B.n283 B.n282 585
R994 B.n638 B.n637 585
R995 B.n639 B.n638 585
R996 B.n635 B.n288 585
R997 B.n288 B.n287 585
R998 B.n634 B.n633 585
R999 B.n633 B.n632 585
R1000 B.n290 B.n289 585
R1001 B.n291 B.n290 585
R1002 B.n625 B.n624 585
R1003 B.n626 B.n625 585
R1004 B.n623 B.n296 585
R1005 B.n296 B.n295 585
R1006 B.n622 B.n621 585
R1007 B.n621 B.n620 585
R1008 B.n298 B.n297 585
R1009 B.n299 B.n298 585
R1010 B.n613 B.n612 585
R1011 B.n614 B.n613 585
R1012 B.n611 B.n304 585
R1013 B.n304 B.n303 585
R1014 B.n610 B.n609 585
R1015 B.n609 B.n608 585
R1016 B.n306 B.n305 585
R1017 B.n307 B.n306 585
R1018 B.n601 B.n600 585
R1019 B.n602 B.n601 585
R1020 B.n599 B.n312 585
R1021 B.n312 B.n311 585
R1022 B.n598 B.n597 585
R1023 B.n597 B.n596 585
R1024 B.n314 B.n313 585
R1025 B.n315 B.n314 585
R1026 B.n589 B.n588 585
R1027 B.n590 B.n589 585
R1028 B.n587 B.n320 585
R1029 B.n320 B.n319 585
R1030 B.n586 B.n585 585
R1031 B.n585 B.n584 585
R1032 B.n322 B.n321 585
R1033 B.n577 B.n322 585
R1034 B.n576 B.n575 585
R1035 B.n578 B.n576 585
R1036 B.n574 B.n327 585
R1037 B.n327 B.n326 585
R1038 B.n573 B.n572 585
R1039 B.n572 B.n571 585
R1040 B.n329 B.n328 585
R1041 B.n330 B.n329 585
R1042 B.n564 B.n563 585
R1043 B.n565 B.n564 585
R1044 B.n333 B.n332 585
R1045 B.n384 B.n382 585
R1046 B.n385 B.n381 585
R1047 B.n385 B.n334 585
R1048 B.n388 B.n387 585
R1049 B.n389 B.n380 585
R1050 B.n391 B.n390 585
R1051 B.n393 B.n379 585
R1052 B.n396 B.n395 585
R1053 B.n397 B.n378 585
R1054 B.n399 B.n398 585
R1055 B.n401 B.n377 585
R1056 B.n404 B.n403 585
R1057 B.n405 B.n376 585
R1058 B.n407 B.n406 585
R1059 B.n409 B.n375 585
R1060 B.n412 B.n411 585
R1061 B.n413 B.n374 585
R1062 B.n415 B.n414 585
R1063 B.n417 B.n373 585
R1064 B.n420 B.n419 585
R1065 B.n421 B.n372 585
R1066 B.n423 B.n422 585
R1067 B.n425 B.n371 585
R1068 B.n428 B.n427 585
R1069 B.n429 B.n370 585
R1070 B.n431 B.n430 585
R1071 B.n433 B.n369 585
R1072 B.n436 B.n435 585
R1073 B.n437 B.n368 585
R1074 B.n439 B.n438 585
R1075 B.n441 B.n367 585
R1076 B.n444 B.n443 585
R1077 B.n445 B.n366 585
R1078 B.n447 B.n446 585
R1079 B.n449 B.n365 585
R1080 B.n452 B.n451 585
R1081 B.n453 B.n364 585
R1082 B.n455 B.n454 585
R1083 B.n457 B.n363 585
R1084 B.n460 B.n459 585
R1085 B.n462 B.n360 585
R1086 B.n464 B.n463 585
R1087 B.n466 B.n359 585
R1088 B.n469 B.n468 585
R1089 B.n470 B.n358 585
R1090 B.n472 B.n471 585
R1091 B.n474 B.n357 585
R1092 B.n477 B.n476 585
R1093 B.n478 B.n356 585
R1094 B.n483 B.n482 585
R1095 B.n485 B.n355 585
R1096 B.n488 B.n487 585
R1097 B.n489 B.n354 585
R1098 B.n491 B.n490 585
R1099 B.n493 B.n353 585
R1100 B.n496 B.n495 585
R1101 B.n497 B.n352 585
R1102 B.n499 B.n498 585
R1103 B.n501 B.n351 585
R1104 B.n504 B.n503 585
R1105 B.n505 B.n350 585
R1106 B.n507 B.n506 585
R1107 B.n509 B.n349 585
R1108 B.n512 B.n511 585
R1109 B.n513 B.n348 585
R1110 B.n515 B.n514 585
R1111 B.n517 B.n347 585
R1112 B.n520 B.n519 585
R1113 B.n521 B.n346 585
R1114 B.n523 B.n522 585
R1115 B.n525 B.n345 585
R1116 B.n528 B.n527 585
R1117 B.n529 B.n344 585
R1118 B.n531 B.n530 585
R1119 B.n533 B.n343 585
R1120 B.n536 B.n535 585
R1121 B.n537 B.n342 585
R1122 B.n539 B.n538 585
R1123 B.n541 B.n341 585
R1124 B.n544 B.n543 585
R1125 B.n545 B.n340 585
R1126 B.n547 B.n546 585
R1127 B.n549 B.n339 585
R1128 B.n552 B.n551 585
R1129 B.n553 B.n338 585
R1130 B.n555 B.n554 585
R1131 B.n557 B.n337 585
R1132 B.n558 B.n336 585
R1133 B.n561 B.n560 585
R1134 B.n562 B.n335 585
R1135 B.n335 B.n334 585
R1136 B.n567 B.n566 585
R1137 B.n566 B.n565 585
R1138 B.n568 B.n331 585
R1139 B.n331 B.n330 585
R1140 B.n570 B.n569 585
R1141 B.n571 B.n570 585
R1142 B.n325 B.n324 585
R1143 B.n326 B.n325 585
R1144 B.n580 B.n579 585
R1145 B.n579 B.n578 585
R1146 B.n581 B.n323 585
R1147 B.n577 B.n323 585
R1148 B.n583 B.n582 585
R1149 B.n584 B.n583 585
R1150 B.n318 B.n317 585
R1151 B.n319 B.n318 585
R1152 B.n592 B.n591 585
R1153 B.n591 B.n590 585
R1154 B.n593 B.n316 585
R1155 B.n316 B.n315 585
R1156 B.n595 B.n594 585
R1157 B.n596 B.n595 585
R1158 B.n310 B.n309 585
R1159 B.n311 B.n310 585
R1160 B.n604 B.n603 585
R1161 B.n603 B.n602 585
R1162 B.n605 B.n308 585
R1163 B.n308 B.n307 585
R1164 B.n607 B.n606 585
R1165 B.n608 B.n607 585
R1166 B.n302 B.n301 585
R1167 B.n303 B.n302 585
R1168 B.n616 B.n615 585
R1169 B.n615 B.n614 585
R1170 B.n617 B.n300 585
R1171 B.n300 B.n299 585
R1172 B.n619 B.n618 585
R1173 B.n620 B.n619 585
R1174 B.n294 B.n293 585
R1175 B.n295 B.n294 585
R1176 B.n628 B.n627 585
R1177 B.n627 B.n626 585
R1178 B.n629 B.n292 585
R1179 B.n292 B.n291 585
R1180 B.n631 B.n630 585
R1181 B.n632 B.n631 585
R1182 B.n286 B.n285 585
R1183 B.n287 B.n286 585
R1184 B.n641 B.n640 585
R1185 B.n640 B.n639 585
R1186 B.n642 B.n284 585
R1187 B.n284 B.n283 585
R1188 B.n644 B.n643 585
R1189 B.n645 B.n644 585
R1190 B.n2 B.n0 585
R1191 B.n4 B.n2 585
R1192 B.n3 B.n1 585
R1193 B.n744 B.n3 585
R1194 B.n742 B.n741 585
R1195 B.n743 B.n742 585
R1196 B.n740 B.n9 585
R1197 B.n9 B.n8 585
R1198 B.n739 B.n738 585
R1199 B.n738 B.n737 585
R1200 B.n11 B.n10 585
R1201 B.n736 B.n11 585
R1202 B.n734 B.n733 585
R1203 B.n735 B.n734 585
R1204 B.n732 B.n16 585
R1205 B.n16 B.n15 585
R1206 B.n731 B.n730 585
R1207 B.n730 B.n729 585
R1208 B.n18 B.n17 585
R1209 B.n728 B.n18 585
R1210 B.n726 B.n725 585
R1211 B.n727 B.n726 585
R1212 B.n724 B.n23 585
R1213 B.n23 B.n22 585
R1214 B.n723 B.n722 585
R1215 B.n722 B.n721 585
R1216 B.n25 B.n24 585
R1217 B.n720 B.n25 585
R1218 B.n718 B.n717 585
R1219 B.n719 B.n718 585
R1220 B.n716 B.n30 585
R1221 B.n30 B.n29 585
R1222 B.n715 B.n714 585
R1223 B.n714 B.n713 585
R1224 B.n32 B.n31 585
R1225 B.n712 B.n32 585
R1226 B.n710 B.n709 585
R1227 B.n711 B.n710 585
R1228 B.n708 B.n37 585
R1229 B.n37 B.n36 585
R1230 B.n707 B.n706 585
R1231 B.n706 B.n705 585
R1232 B.n39 B.n38 585
R1233 B.n704 B.n39 585
R1234 B.n702 B.n701 585
R1235 B.n703 B.n702 585
R1236 B.n700 B.n43 585
R1237 B.n46 B.n43 585
R1238 B.n699 B.n698 585
R1239 B.n698 B.n697 585
R1240 B.n45 B.n44 585
R1241 B.n696 B.n45 585
R1242 B.n694 B.n693 585
R1243 B.n695 B.n694 585
R1244 B.n692 B.n51 585
R1245 B.n51 B.n50 585
R1246 B.n691 B.n690 585
R1247 B.n690 B.n689 585
R1248 B.n747 B.n746 585
R1249 B.n746 B.n745 585
R1250 B.n566 B.n333 492.5
R1251 B.n690 B.n53 492.5
R1252 B.n564 B.n335 492.5
R1253 B.n686 B.n54 492.5
R1254 B.n479 B.t12 475.248
R1255 B.n361 B.t16 475.248
R1256 B.n103 B.t19 475.248
R1257 B.n100 B.t8 475.248
R1258 B.n479 B.t15 300.356
R1259 B.n100 B.t10 300.356
R1260 B.n361 B.t18 300.356
R1261 B.n103 B.t20 300.356
R1262 B.n480 B.t14 274.175
R1263 B.n101 B.t11 274.175
R1264 B.n362 B.t17 274.175
R1265 B.n104 B.t21 274.175
R1266 B.n688 B.n687 256.663
R1267 B.n688 B.n98 256.663
R1268 B.n688 B.n97 256.663
R1269 B.n688 B.n96 256.663
R1270 B.n688 B.n95 256.663
R1271 B.n688 B.n94 256.663
R1272 B.n688 B.n93 256.663
R1273 B.n688 B.n92 256.663
R1274 B.n688 B.n91 256.663
R1275 B.n688 B.n90 256.663
R1276 B.n688 B.n89 256.663
R1277 B.n688 B.n88 256.663
R1278 B.n688 B.n87 256.663
R1279 B.n688 B.n86 256.663
R1280 B.n688 B.n85 256.663
R1281 B.n688 B.n84 256.663
R1282 B.n688 B.n83 256.663
R1283 B.n688 B.n82 256.663
R1284 B.n688 B.n81 256.663
R1285 B.n688 B.n80 256.663
R1286 B.n688 B.n79 256.663
R1287 B.n688 B.n78 256.663
R1288 B.n688 B.n77 256.663
R1289 B.n688 B.n76 256.663
R1290 B.n688 B.n75 256.663
R1291 B.n688 B.n74 256.663
R1292 B.n688 B.n73 256.663
R1293 B.n688 B.n72 256.663
R1294 B.n688 B.n71 256.663
R1295 B.n688 B.n70 256.663
R1296 B.n688 B.n69 256.663
R1297 B.n688 B.n68 256.663
R1298 B.n688 B.n67 256.663
R1299 B.n688 B.n66 256.663
R1300 B.n688 B.n65 256.663
R1301 B.n688 B.n64 256.663
R1302 B.n688 B.n63 256.663
R1303 B.n688 B.n62 256.663
R1304 B.n688 B.n61 256.663
R1305 B.n688 B.n60 256.663
R1306 B.n688 B.n59 256.663
R1307 B.n688 B.n58 256.663
R1308 B.n688 B.n57 256.663
R1309 B.n688 B.n56 256.663
R1310 B.n688 B.n55 256.663
R1311 B.n383 B.n334 256.663
R1312 B.n386 B.n334 256.663
R1313 B.n392 B.n334 256.663
R1314 B.n394 B.n334 256.663
R1315 B.n400 B.n334 256.663
R1316 B.n402 B.n334 256.663
R1317 B.n408 B.n334 256.663
R1318 B.n410 B.n334 256.663
R1319 B.n416 B.n334 256.663
R1320 B.n418 B.n334 256.663
R1321 B.n424 B.n334 256.663
R1322 B.n426 B.n334 256.663
R1323 B.n432 B.n334 256.663
R1324 B.n434 B.n334 256.663
R1325 B.n440 B.n334 256.663
R1326 B.n442 B.n334 256.663
R1327 B.n448 B.n334 256.663
R1328 B.n450 B.n334 256.663
R1329 B.n456 B.n334 256.663
R1330 B.n458 B.n334 256.663
R1331 B.n465 B.n334 256.663
R1332 B.n467 B.n334 256.663
R1333 B.n473 B.n334 256.663
R1334 B.n475 B.n334 256.663
R1335 B.n484 B.n334 256.663
R1336 B.n486 B.n334 256.663
R1337 B.n492 B.n334 256.663
R1338 B.n494 B.n334 256.663
R1339 B.n500 B.n334 256.663
R1340 B.n502 B.n334 256.663
R1341 B.n508 B.n334 256.663
R1342 B.n510 B.n334 256.663
R1343 B.n516 B.n334 256.663
R1344 B.n518 B.n334 256.663
R1345 B.n524 B.n334 256.663
R1346 B.n526 B.n334 256.663
R1347 B.n532 B.n334 256.663
R1348 B.n534 B.n334 256.663
R1349 B.n540 B.n334 256.663
R1350 B.n542 B.n334 256.663
R1351 B.n548 B.n334 256.663
R1352 B.n550 B.n334 256.663
R1353 B.n556 B.n334 256.663
R1354 B.n559 B.n334 256.663
R1355 B.n566 B.n331 163.367
R1356 B.n570 B.n331 163.367
R1357 B.n570 B.n325 163.367
R1358 B.n579 B.n325 163.367
R1359 B.n579 B.n323 163.367
R1360 B.n583 B.n323 163.367
R1361 B.n583 B.n318 163.367
R1362 B.n591 B.n318 163.367
R1363 B.n591 B.n316 163.367
R1364 B.n595 B.n316 163.367
R1365 B.n595 B.n310 163.367
R1366 B.n603 B.n310 163.367
R1367 B.n603 B.n308 163.367
R1368 B.n607 B.n308 163.367
R1369 B.n607 B.n302 163.367
R1370 B.n615 B.n302 163.367
R1371 B.n615 B.n300 163.367
R1372 B.n619 B.n300 163.367
R1373 B.n619 B.n294 163.367
R1374 B.n627 B.n294 163.367
R1375 B.n627 B.n292 163.367
R1376 B.n631 B.n292 163.367
R1377 B.n631 B.n286 163.367
R1378 B.n640 B.n286 163.367
R1379 B.n640 B.n284 163.367
R1380 B.n644 B.n284 163.367
R1381 B.n644 B.n2 163.367
R1382 B.n746 B.n2 163.367
R1383 B.n746 B.n3 163.367
R1384 B.n742 B.n3 163.367
R1385 B.n742 B.n9 163.367
R1386 B.n738 B.n9 163.367
R1387 B.n738 B.n11 163.367
R1388 B.n734 B.n11 163.367
R1389 B.n734 B.n16 163.367
R1390 B.n730 B.n16 163.367
R1391 B.n730 B.n18 163.367
R1392 B.n726 B.n18 163.367
R1393 B.n726 B.n23 163.367
R1394 B.n722 B.n23 163.367
R1395 B.n722 B.n25 163.367
R1396 B.n718 B.n25 163.367
R1397 B.n718 B.n30 163.367
R1398 B.n714 B.n30 163.367
R1399 B.n714 B.n32 163.367
R1400 B.n710 B.n32 163.367
R1401 B.n710 B.n37 163.367
R1402 B.n706 B.n37 163.367
R1403 B.n706 B.n39 163.367
R1404 B.n702 B.n39 163.367
R1405 B.n702 B.n43 163.367
R1406 B.n698 B.n43 163.367
R1407 B.n698 B.n45 163.367
R1408 B.n694 B.n45 163.367
R1409 B.n694 B.n51 163.367
R1410 B.n690 B.n51 163.367
R1411 B.n385 B.n384 163.367
R1412 B.n387 B.n385 163.367
R1413 B.n391 B.n380 163.367
R1414 B.n395 B.n393 163.367
R1415 B.n399 B.n378 163.367
R1416 B.n403 B.n401 163.367
R1417 B.n407 B.n376 163.367
R1418 B.n411 B.n409 163.367
R1419 B.n415 B.n374 163.367
R1420 B.n419 B.n417 163.367
R1421 B.n423 B.n372 163.367
R1422 B.n427 B.n425 163.367
R1423 B.n431 B.n370 163.367
R1424 B.n435 B.n433 163.367
R1425 B.n439 B.n368 163.367
R1426 B.n443 B.n441 163.367
R1427 B.n447 B.n366 163.367
R1428 B.n451 B.n449 163.367
R1429 B.n455 B.n364 163.367
R1430 B.n459 B.n457 163.367
R1431 B.n464 B.n360 163.367
R1432 B.n468 B.n466 163.367
R1433 B.n472 B.n358 163.367
R1434 B.n476 B.n474 163.367
R1435 B.n483 B.n356 163.367
R1436 B.n487 B.n485 163.367
R1437 B.n491 B.n354 163.367
R1438 B.n495 B.n493 163.367
R1439 B.n499 B.n352 163.367
R1440 B.n503 B.n501 163.367
R1441 B.n507 B.n350 163.367
R1442 B.n511 B.n509 163.367
R1443 B.n515 B.n348 163.367
R1444 B.n519 B.n517 163.367
R1445 B.n523 B.n346 163.367
R1446 B.n527 B.n525 163.367
R1447 B.n531 B.n344 163.367
R1448 B.n535 B.n533 163.367
R1449 B.n539 B.n342 163.367
R1450 B.n543 B.n541 163.367
R1451 B.n547 B.n340 163.367
R1452 B.n551 B.n549 163.367
R1453 B.n555 B.n338 163.367
R1454 B.n558 B.n557 163.367
R1455 B.n560 B.n335 163.367
R1456 B.n564 B.n329 163.367
R1457 B.n572 B.n329 163.367
R1458 B.n572 B.n327 163.367
R1459 B.n576 B.n327 163.367
R1460 B.n576 B.n322 163.367
R1461 B.n585 B.n322 163.367
R1462 B.n585 B.n320 163.367
R1463 B.n589 B.n320 163.367
R1464 B.n589 B.n314 163.367
R1465 B.n597 B.n314 163.367
R1466 B.n597 B.n312 163.367
R1467 B.n601 B.n312 163.367
R1468 B.n601 B.n306 163.367
R1469 B.n609 B.n306 163.367
R1470 B.n609 B.n304 163.367
R1471 B.n613 B.n304 163.367
R1472 B.n613 B.n298 163.367
R1473 B.n621 B.n298 163.367
R1474 B.n621 B.n296 163.367
R1475 B.n625 B.n296 163.367
R1476 B.n625 B.n290 163.367
R1477 B.n633 B.n290 163.367
R1478 B.n633 B.n288 163.367
R1479 B.n638 B.n288 163.367
R1480 B.n638 B.n282 163.367
R1481 B.n646 B.n282 163.367
R1482 B.n647 B.n646 163.367
R1483 B.n647 B.n5 163.367
R1484 B.n6 B.n5 163.367
R1485 B.n7 B.n6 163.367
R1486 B.n652 B.n7 163.367
R1487 B.n652 B.n12 163.367
R1488 B.n13 B.n12 163.367
R1489 B.n14 B.n13 163.367
R1490 B.n657 B.n14 163.367
R1491 B.n657 B.n19 163.367
R1492 B.n20 B.n19 163.367
R1493 B.n21 B.n20 163.367
R1494 B.n662 B.n21 163.367
R1495 B.n662 B.n26 163.367
R1496 B.n27 B.n26 163.367
R1497 B.n28 B.n27 163.367
R1498 B.n667 B.n28 163.367
R1499 B.n667 B.n33 163.367
R1500 B.n34 B.n33 163.367
R1501 B.n35 B.n34 163.367
R1502 B.n672 B.n35 163.367
R1503 B.n672 B.n40 163.367
R1504 B.n41 B.n40 163.367
R1505 B.n42 B.n41 163.367
R1506 B.n677 B.n42 163.367
R1507 B.n677 B.n47 163.367
R1508 B.n48 B.n47 163.367
R1509 B.n49 B.n48 163.367
R1510 B.n682 B.n49 163.367
R1511 B.n682 B.n54 163.367
R1512 B.n108 B.n107 163.367
R1513 B.n112 B.n111 163.367
R1514 B.n116 B.n115 163.367
R1515 B.n120 B.n119 163.367
R1516 B.n124 B.n123 163.367
R1517 B.n128 B.n127 163.367
R1518 B.n132 B.n131 163.367
R1519 B.n136 B.n135 163.367
R1520 B.n140 B.n139 163.367
R1521 B.n144 B.n143 163.367
R1522 B.n148 B.n147 163.367
R1523 B.n152 B.n151 163.367
R1524 B.n156 B.n155 163.367
R1525 B.n160 B.n159 163.367
R1526 B.n164 B.n163 163.367
R1527 B.n168 B.n167 163.367
R1528 B.n172 B.n171 163.367
R1529 B.n176 B.n175 163.367
R1530 B.n180 B.n179 163.367
R1531 B.n184 B.n183 163.367
R1532 B.n188 B.n187 163.367
R1533 B.n192 B.n191 163.367
R1534 B.n196 B.n195 163.367
R1535 B.n200 B.n199 163.367
R1536 B.n204 B.n203 163.367
R1537 B.n208 B.n207 163.367
R1538 B.n212 B.n211 163.367
R1539 B.n216 B.n215 163.367
R1540 B.n220 B.n219 163.367
R1541 B.n224 B.n223 163.367
R1542 B.n228 B.n227 163.367
R1543 B.n232 B.n231 163.367
R1544 B.n236 B.n235 163.367
R1545 B.n240 B.n239 163.367
R1546 B.n244 B.n243 163.367
R1547 B.n248 B.n247 163.367
R1548 B.n252 B.n251 163.367
R1549 B.n256 B.n255 163.367
R1550 B.n260 B.n259 163.367
R1551 B.n264 B.n263 163.367
R1552 B.n268 B.n267 163.367
R1553 B.n272 B.n271 163.367
R1554 B.n276 B.n275 163.367
R1555 B.n278 B.n99 163.367
R1556 B.n565 B.n334 79.2503
R1557 B.n689 B.n688 79.2503
R1558 B.n383 B.n333 71.676
R1559 B.n387 B.n386 71.676
R1560 B.n392 B.n391 71.676
R1561 B.n395 B.n394 71.676
R1562 B.n400 B.n399 71.676
R1563 B.n403 B.n402 71.676
R1564 B.n408 B.n407 71.676
R1565 B.n411 B.n410 71.676
R1566 B.n416 B.n415 71.676
R1567 B.n419 B.n418 71.676
R1568 B.n424 B.n423 71.676
R1569 B.n427 B.n426 71.676
R1570 B.n432 B.n431 71.676
R1571 B.n435 B.n434 71.676
R1572 B.n440 B.n439 71.676
R1573 B.n443 B.n442 71.676
R1574 B.n448 B.n447 71.676
R1575 B.n451 B.n450 71.676
R1576 B.n456 B.n455 71.676
R1577 B.n459 B.n458 71.676
R1578 B.n465 B.n464 71.676
R1579 B.n468 B.n467 71.676
R1580 B.n473 B.n472 71.676
R1581 B.n476 B.n475 71.676
R1582 B.n484 B.n483 71.676
R1583 B.n487 B.n486 71.676
R1584 B.n492 B.n491 71.676
R1585 B.n495 B.n494 71.676
R1586 B.n500 B.n499 71.676
R1587 B.n503 B.n502 71.676
R1588 B.n508 B.n507 71.676
R1589 B.n511 B.n510 71.676
R1590 B.n516 B.n515 71.676
R1591 B.n519 B.n518 71.676
R1592 B.n524 B.n523 71.676
R1593 B.n527 B.n526 71.676
R1594 B.n532 B.n531 71.676
R1595 B.n535 B.n534 71.676
R1596 B.n540 B.n539 71.676
R1597 B.n543 B.n542 71.676
R1598 B.n548 B.n547 71.676
R1599 B.n551 B.n550 71.676
R1600 B.n556 B.n555 71.676
R1601 B.n559 B.n558 71.676
R1602 B.n55 B.n53 71.676
R1603 B.n108 B.n56 71.676
R1604 B.n112 B.n57 71.676
R1605 B.n116 B.n58 71.676
R1606 B.n120 B.n59 71.676
R1607 B.n124 B.n60 71.676
R1608 B.n128 B.n61 71.676
R1609 B.n132 B.n62 71.676
R1610 B.n136 B.n63 71.676
R1611 B.n140 B.n64 71.676
R1612 B.n144 B.n65 71.676
R1613 B.n148 B.n66 71.676
R1614 B.n152 B.n67 71.676
R1615 B.n156 B.n68 71.676
R1616 B.n160 B.n69 71.676
R1617 B.n164 B.n70 71.676
R1618 B.n168 B.n71 71.676
R1619 B.n172 B.n72 71.676
R1620 B.n176 B.n73 71.676
R1621 B.n180 B.n74 71.676
R1622 B.n184 B.n75 71.676
R1623 B.n188 B.n76 71.676
R1624 B.n192 B.n77 71.676
R1625 B.n196 B.n78 71.676
R1626 B.n200 B.n79 71.676
R1627 B.n204 B.n80 71.676
R1628 B.n208 B.n81 71.676
R1629 B.n212 B.n82 71.676
R1630 B.n216 B.n83 71.676
R1631 B.n220 B.n84 71.676
R1632 B.n224 B.n85 71.676
R1633 B.n228 B.n86 71.676
R1634 B.n232 B.n87 71.676
R1635 B.n236 B.n88 71.676
R1636 B.n240 B.n89 71.676
R1637 B.n244 B.n90 71.676
R1638 B.n248 B.n91 71.676
R1639 B.n252 B.n92 71.676
R1640 B.n256 B.n93 71.676
R1641 B.n260 B.n94 71.676
R1642 B.n264 B.n95 71.676
R1643 B.n268 B.n96 71.676
R1644 B.n272 B.n97 71.676
R1645 B.n276 B.n98 71.676
R1646 B.n687 B.n99 71.676
R1647 B.n687 B.n686 71.676
R1648 B.n278 B.n98 71.676
R1649 B.n275 B.n97 71.676
R1650 B.n271 B.n96 71.676
R1651 B.n267 B.n95 71.676
R1652 B.n263 B.n94 71.676
R1653 B.n259 B.n93 71.676
R1654 B.n255 B.n92 71.676
R1655 B.n251 B.n91 71.676
R1656 B.n247 B.n90 71.676
R1657 B.n243 B.n89 71.676
R1658 B.n239 B.n88 71.676
R1659 B.n235 B.n87 71.676
R1660 B.n231 B.n86 71.676
R1661 B.n227 B.n85 71.676
R1662 B.n223 B.n84 71.676
R1663 B.n219 B.n83 71.676
R1664 B.n215 B.n82 71.676
R1665 B.n211 B.n81 71.676
R1666 B.n207 B.n80 71.676
R1667 B.n203 B.n79 71.676
R1668 B.n199 B.n78 71.676
R1669 B.n195 B.n77 71.676
R1670 B.n191 B.n76 71.676
R1671 B.n187 B.n75 71.676
R1672 B.n183 B.n74 71.676
R1673 B.n179 B.n73 71.676
R1674 B.n175 B.n72 71.676
R1675 B.n171 B.n71 71.676
R1676 B.n167 B.n70 71.676
R1677 B.n163 B.n69 71.676
R1678 B.n159 B.n68 71.676
R1679 B.n155 B.n67 71.676
R1680 B.n151 B.n66 71.676
R1681 B.n147 B.n65 71.676
R1682 B.n143 B.n64 71.676
R1683 B.n139 B.n63 71.676
R1684 B.n135 B.n62 71.676
R1685 B.n131 B.n61 71.676
R1686 B.n127 B.n60 71.676
R1687 B.n123 B.n59 71.676
R1688 B.n119 B.n58 71.676
R1689 B.n115 B.n57 71.676
R1690 B.n111 B.n56 71.676
R1691 B.n107 B.n55 71.676
R1692 B.n384 B.n383 71.676
R1693 B.n386 B.n380 71.676
R1694 B.n393 B.n392 71.676
R1695 B.n394 B.n378 71.676
R1696 B.n401 B.n400 71.676
R1697 B.n402 B.n376 71.676
R1698 B.n409 B.n408 71.676
R1699 B.n410 B.n374 71.676
R1700 B.n417 B.n416 71.676
R1701 B.n418 B.n372 71.676
R1702 B.n425 B.n424 71.676
R1703 B.n426 B.n370 71.676
R1704 B.n433 B.n432 71.676
R1705 B.n434 B.n368 71.676
R1706 B.n441 B.n440 71.676
R1707 B.n442 B.n366 71.676
R1708 B.n449 B.n448 71.676
R1709 B.n450 B.n364 71.676
R1710 B.n457 B.n456 71.676
R1711 B.n458 B.n360 71.676
R1712 B.n466 B.n465 71.676
R1713 B.n467 B.n358 71.676
R1714 B.n474 B.n473 71.676
R1715 B.n475 B.n356 71.676
R1716 B.n485 B.n484 71.676
R1717 B.n486 B.n354 71.676
R1718 B.n493 B.n492 71.676
R1719 B.n494 B.n352 71.676
R1720 B.n501 B.n500 71.676
R1721 B.n502 B.n350 71.676
R1722 B.n509 B.n508 71.676
R1723 B.n510 B.n348 71.676
R1724 B.n517 B.n516 71.676
R1725 B.n518 B.n346 71.676
R1726 B.n525 B.n524 71.676
R1727 B.n526 B.n344 71.676
R1728 B.n533 B.n532 71.676
R1729 B.n534 B.n342 71.676
R1730 B.n541 B.n540 71.676
R1731 B.n542 B.n340 71.676
R1732 B.n549 B.n548 71.676
R1733 B.n550 B.n338 71.676
R1734 B.n557 B.n556 71.676
R1735 B.n560 B.n559 71.676
R1736 B.n481 B.n480 59.5399
R1737 B.n461 B.n362 59.5399
R1738 B.n105 B.n104 59.5399
R1739 B.n102 B.n101 59.5399
R1740 B.n565 B.n330 44.5376
R1741 B.n571 B.n330 44.5376
R1742 B.n571 B.n326 44.5376
R1743 B.n578 B.n326 44.5376
R1744 B.n578 B.n577 44.5376
R1745 B.n584 B.n319 44.5376
R1746 B.n590 B.n319 44.5376
R1747 B.n590 B.n315 44.5376
R1748 B.n596 B.n315 44.5376
R1749 B.n596 B.n311 44.5376
R1750 B.n602 B.n311 44.5376
R1751 B.n608 B.n307 44.5376
R1752 B.n608 B.n303 44.5376
R1753 B.n614 B.n303 44.5376
R1754 B.n620 B.n299 44.5376
R1755 B.n620 B.n295 44.5376
R1756 B.n626 B.n295 44.5376
R1757 B.n632 B.n291 44.5376
R1758 B.n632 B.n287 44.5376
R1759 B.n639 B.n287 44.5376
R1760 B.n645 B.n283 44.5376
R1761 B.n645 B.n4 44.5376
R1762 B.n745 B.n4 44.5376
R1763 B.n745 B.n744 44.5376
R1764 B.n744 B.n743 44.5376
R1765 B.n743 B.n8 44.5376
R1766 B.n737 B.n736 44.5376
R1767 B.n736 B.n735 44.5376
R1768 B.n735 B.n15 44.5376
R1769 B.n729 B.n728 44.5376
R1770 B.n728 B.n727 44.5376
R1771 B.n727 B.n22 44.5376
R1772 B.n721 B.n720 44.5376
R1773 B.n720 B.n719 44.5376
R1774 B.n719 B.n29 44.5376
R1775 B.n713 B.n712 44.5376
R1776 B.n712 B.n711 44.5376
R1777 B.n711 B.n36 44.5376
R1778 B.n705 B.n36 44.5376
R1779 B.n705 B.n704 44.5376
R1780 B.n704 B.n703 44.5376
R1781 B.n697 B.n46 44.5376
R1782 B.n697 B.n696 44.5376
R1783 B.n696 B.n695 44.5376
R1784 B.n695 B.n50 44.5376
R1785 B.n689 B.n50 44.5376
R1786 B.n691 B.n52 32.0005
R1787 B.n685 B.n684 32.0005
R1788 B.n563 B.n562 32.0005
R1789 B.n567 B.n332 32.0005
R1790 B.n584 B.t13 30.1285
R1791 B.n703 B.t9 30.1285
R1792 B.t1 B.n283 26.1988
R1793 B.t3 B.n8 26.1988
R1794 B.n480 B.n479 26.1823
R1795 B.n362 B.n361 26.1823
R1796 B.n104 B.n103 26.1823
R1797 B.n101 B.n100 26.1823
R1798 B.t2 B.n291 24.8889
R1799 B.t4 B.n15 24.8889
R1800 B.t7 B.n299 23.5789
R1801 B.t5 B.n22 23.5789
R1802 B.n602 B.t0 22.269
R1803 B.t0 B.n307 22.269
R1804 B.t6 B.n29 22.269
R1805 B.n713 B.t6 22.269
R1806 B.n614 B.t7 20.9591
R1807 B.n721 B.t5 20.9591
R1808 B.n626 B.t2 19.6492
R1809 B.n729 B.t4 19.6492
R1810 B.n639 B.t1 18.3393
R1811 B.n737 B.t3 18.3393
R1812 B B.n747 18.0485
R1813 B.n577 B.t13 14.4096
R1814 B.n46 B.t9 14.4096
R1815 B.n106 B.n52 10.6151
R1816 B.n109 B.n106 10.6151
R1817 B.n110 B.n109 10.6151
R1818 B.n113 B.n110 10.6151
R1819 B.n114 B.n113 10.6151
R1820 B.n117 B.n114 10.6151
R1821 B.n118 B.n117 10.6151
R1822 B.n121 B.n118 10.6151
R1823 B.n122 B.n121 10.6151
R1824 B.n125 B.n122 10.6151
R1825 B.n126 B.n125 10.6151
R1826 B.n129 B.n126 10.6151
R1827 B.n130 B.n129 10.6151
R1828 B.n133 B.n130 10.6151
R1829 B.n134 B.n133 10.6151
R1830 B.n137 B.n134 10.6151
R1831 B.n138 B.n137 10.6151
R1832 B.n141 B.n138 10.6151
R1833 B.n142 B.n141 10.6151
R1834 B.n145 B.n142 10.6151
R1835 B.n146 B.n145 10.6151
R1836 B.n149 B.n146 10.6151
R1837 B.n150 B.n149 10.6151
R1838 B.n153 B.n150 10.6151
R1839 B.n154 B.n153 10.6151
R1840 B.n157 B.n154 10.6151
R1841 B.n158 B.n157 10.6151
R1842 B.n161 B.n158 10.6151
R1843 B.n162 B.n161 10.6151
R1844 B.n165 B.n162 10.6151
R1845 B.n166 B.n165 10.6151
R1846 B.n169 B.n166 10.6151
R1847 B.n170 B.n169 10.6151
R1848 B.n173 B.n170 10.6151
R1849 B.n174 B.n173 10.6151
R1850 B.n177 B.n174 10.6151
R1851 B.n178 B.n177 10.6151
R1852 B.n181 B.n178 10.6151
R1853 B.n182 B.n181 10.6151
R1854 B.n186 B.n185 10.6151
R1855 B.n189 B.n186 10.6151
R1856 B.n190 B.n189 10.6151
R1857 B.n193 B.n190 10.6151
R1858 B.n194 B.n193 10.6151
R1859 B.n197 B.n194 10.6151
R1860 B.n198 B.n197 10.6151
R1861 B.n201 B.n198 10.6151
R1862 B.n202 B.n201 10.6151
R1863 B.n206 B.n205 10.6151
R1864 B.n209 B.n206 10.6151
R1865 B.n210 B.n209 10.6151
R1866 B.n213 B.n210 10.6151
R1867 B.n214 B.n213 10.6151
R1868 B.n217 B.n214 10.6151
R1869 B.n218 B.n217 10.6151
R1870 B.n221 B.n218 10.6151
R1871 B.n222 B.n221 10.6151
R1872 B.n225 B.n222 10.6151
R1873 B.n226 B.n225 10.6151
R1874 B.n229 B.n226 10.6151
R1875 B.n230 B.n229 10.6151
R1876 B.n233 B.n230 10.6151
R1877 B.n234 B.n233 10.6151
R1878 B.n237 B.n234 10.6151
R1879 B.n238 B.n237 10.6151
R1880 B.n241 B.n238 10.6151
R1881 B.n242 B.n241 10.6151
R1882 B.n245 B.n242 10.6151
R1883 B.n246 B.n245 10.6151
R1884 B.n249 B.n246 10.6151
R1885 B.n250 B.n249 10.6151
R1886 B.n253 B.n250 10.6151
R1887 B.n254 B.n253 10.6151
R1888 B.n257 B.n254 10.6151
R1889 B.n258 B.n257 10.6151
R1890 B.n261 B.n258 10.6151
R1891 B.n262 B.n261 10.6151
R1892 B.n265 B.n262 10.6151
R1893 B.n266 B.n265 10.6151
R1894 B.n269 B.n266 10.6151
R1895 B.n270 B.n269 10.6151
R1896 B.n273 B.n270 10.6151
R1897 B.n274 B.n273 10.6151
R1898 B.n277 B.n274 10.6151
R1899 B.n279 B.n277 10.6151
R1900 B.n280 B.n279 10.6151
R1901 B.n685 B.n280 10.6151
R1902 B.n563 B.n328 10.6151
R1903 B.n573 B.n328 10.6151
R1904 B.n574 B.n573 10.6151
R1905 B.n575 B.n574 10.6151
R1906 B.n575 B.n321 10.6151
R1907 B.n586 B.n321 10.6151
R1908 B.n587 B.n586 10.6151
R1909 B.n588 B.n587 10.6151
R1910 B.n588 B.n313 10.6151
R1911 B.n598 B.n313 10.6151
R1912 B.n599 B.n598 10.6151
R1913 B.n600 B.n599 10.6151
R1914 B.n600 B.n305 10.6151
R1915 B.n610 B.n305 10.6151
R1916 B.n611 B.n610 10.6151
R1917 B.n612 B.n611 10.6151
R1918 B.n612 B.n297 10.6151
R1919 B.n622 B.n297 10.6151
R1920 B.n623 B.n622 10.6151
R1921 B.n624 B.n623 10.6151
R1922 B.n624 B.n289 10.6151
R1923 B.n634 B.n289 10.6151
R1924 B.n635 B.n634 10.6151
R1925 B.n637 B.n635 10.6151
R1926 B.n637 B.n636 10.6151
R1927 B.n636 B.n281 10.6151
R1928 B.n648 B.n281 10.6151
R1929 B.n649 B.n648 10.6151
R1930 B.n650 B.n649 10.6151
R1931 B.n651 B.n650 10.6151
R1932 B.n653 B.n651 10.6151
R1933 B.n654 B.n653 10.6151
R1934 B.n655 B.n654 10.6151
R1935 B.n656 B.n655 10.6151
R1936 B.n658 B.n656 10.6151
R1937 B.n659 B.n658 10.6151
R1938 B.n660 B.n659 10.6151
R1939 B.n661 B.n660 10.6151
R1940 B.n663 B.n661 10.6151
R1941 B.n664 B.n663 10.6151
R1942 B.n665 B.n664 10.6151
R1943 B.n666 B.n665 10.6151
R1944 B.n668 B.n666 10.6151
R1945 B.n669 B.n668 10.6151
R1946 B.n670 B.n669 10.6151
R1947 B.n671 B.n670 10.6151
R1948 B.n673 B.n671 10.6151
R1949 B.n674 B.n673 10.6151
R1950 B.n675 B.n674 10.6151
R1951 B.n676 B.n675 10.6151
R1952 B.n678 B.n676 10.6151
R1953 B.n679 B.n678 10.6151
R1954 B.n680 B.n679 10.6151
R1955 B.n681 B.n680 10.6151
R1956 B.n683 B.n681 10.6151
R1957 B.n684 B.n683 10.6151
R1958 B.n382 B.n332 10.6151
R1959 B.n382 B.n381 10.6151
R1960 B.n388 B.n381 10.6151
R1961 B.n389 B.n388 10.6151
R1962 B.n390 B.n389 10.6151
R1963 B.n390 B.n379 10.6151
R1964 B.n396 B.n379 10.6151
R1965 B.n397 B.n396 10.6151
R1966 B.n398 B.n397 10.6151
R1967 B.n398 B.n377 10.6151
R1968 B.n404 B.n377 10.6151
R1969 B.n405 B.n404 10.6151
R1970 B.n406 B.n405 10.6151
R1971 B.n406 B.n375 10.6151
R1972 B.n412 B.n375 10.6151
R1973 B.n413 B.n412 10.6151
R1974 B.n414 B.n413 10.6151
R1975 B.n414 B.n373 10.6151
R1976 B.n420 B.n373 10.6151
R1977 B.n421 B.n420 10.6151
R1978 B.n422 B.n421 10.6151
R1979 B.n422 B.n371 10.6151
R1980 B.n428 B.n371 10.6151
R1981 B.n429 B.n428 10.6151
R1982 B.n430 B.n429 10.6151
R1983 B.n430 B.n369 10.6151
R1984 B.n436 B.n369 10.6151
R1985 B.n437 B.n436 10.6151
R1986 B.n438 B.n437 10.6151
R1987 B.n438 B.n367 10.6151
R1988 B.n444 B.n367 10.6151
R1989 B.n445 B.n444 10.6151
R1990 B.n446 B.n445 10.6151
R1991 B.n446 B.n365 10.6151
R1992 B.n452 B.n365 10.6151
R1993 B.n453 B.n452 10.6151
R1994 B.n454 B.n453 10.6151
R1995 B.n454 B.n363 10.6151
R1996 B.n460 B.n363 10.6151
R1997 B.n463 B.n462 10.6151
R1998 B.n463 B.n359 10.6151
R1999 B.n469 B.n359 10.6151
R2000 B.n470 B.n469 10.6151
R2001 B.n471 B.n470 10.6151
R2002 B.n471 B.n357 10.6151
R2003 B.n477 B.n357 10.6151
R2004 B.n478 B.n477 10.6151
R2005 B.n482 B.n478 10.6151
R2006 B.n488 B.n355 10.6151
R2007 B.n489 B.n488 10.6151
R2008 B.n490 B.n489 10.6151
R2009 B.n490 B.n353 10.6151
R2010 B.n496 B.n353 10.6151
R2011 B.n497 B.n496 10.6151
R2012 B.n498 B.n497 10.6151
R2013 B.n498 B.n351 10.6151
R2014 B.n504 B.n351 10.6151
R2015 B.n505 B.n504 10.6151
R2016 B.n506 B.n505 10.6151
R2017 B.n506 B.n349 10.6151
R2018 B.n512 B.n349 10.6151
R2019 B.n513 B.n512 10.6151
R2020 B.n514 B.n513 10.6151
R2021 B.n514 B.n347 10.6151
R2022 B.n520 B.n347 10.6151
R2023 B.n521 B.n520 10.6151
R2024 B.n522 B.n521 10.6151
R2025 B.n522 B.n345 10.6151
R2026 B.n528 B.n345 10.6151
R2027 B.n529 B.n528 10.6151
R2028 B.n530 B.n529 10.6151
R2029 B.n530 B.n343 10.6151
R2030 B.n536 B.n343 10.6151
R2031 B.n537 B.n536 10.6151
R2032 B.n538 B.n537 10.6151
R2033 B.n538 B.n341 10.6151
R2034 B.n544 B.n341 10.6151
R2035 B.n545 B.n544 10.6151
R2036 B.n546 B.n545 10.6151
R2037 B.n546 B.n339 10.6151
R2038 B.n552 B.n339 10.6151
R2039 B.n553 B.n552 10.6151
R2040 B.n554 B.n553 10.6151
R2041 B.n554 B.n337 10.6151
R2042 B.n337 B.n336 10.6151
R2043 B.n561 B.n336 10.6151
R2044 B.n562 B.n561 10.6151
R2045 B.n568 B.n567 10.6151
R2046 B.n569 B.n568 10.6151
R2047 B.n569 B.n324 10.6151
R2048 B.n580 B.n324 10.6151
R2049 B.n581 B.n580 10.6151
R2050 B.n582 B.n581 10.6151
R2051 B.n582 B.n317 10.6151
R2052 B.n592 B.n317 10.6151
R2053 B.n593 B.n592 10.6151
R2054 B.n594 B.n593 10.6151
R2055 B.n594 B.n309 10.6151
R2056 B.n604 B.n309 10.6151
R2057 B.n605 B.n604 10.6151
R2058 B.n606 B.n605 10.6151
R2059 B.n606 B.n301 10.6151
R2060 B.n616 B.n301 10.6151
R2061 B.n617 B.n616 10.6151
R2062 B.n618 B.n617 10.6151
R2063 B.n618 B.n293 10.6151
R2064 B.n628 B.n293 10.6151
R2065 B.n629 B.n628 10.6151
R2066 B.n630 B.n629 10.6151
R2067 B.n630 B.n285 10.6151
R2068 B.n641 B.n285 10.6151
R2069 B.n642 B.n641 10.6151
R2070 B.n643 B.n642 10.6151
R2071 B.n643 B.n0 10.6151
R2072 B.n741 B.n1 10.6151
R2073 B.n741 B.n740 10.6151
R2074 B.n740 B.n739 10.6151
R2075 B.n739 B.n10 10.6151
R2076 B.n733 B.n10 10.6151
R2077 B.n733 B.n732 10.6151
R2078 B.n732 B.n731 10.6151
R2079 B.n731 B.n17 10.6151
R2080 B.n725 B.n17 10.6151
R2081 B.n725 B.n724 10.6151
R2082 B.n724 B.n723 10.6151
R2083 B.n723 B.n24 10.6151
R2084 B.n717 B.n24 10.6151
R2085 B.n717 B.n716 10.6151
R2086 B.n716 B.n715 10.6151
R2087 B.n715 B.n31 10.6151
R2088 B.n709 B.n31 10.6151
R2089 B.n709 B.n708 10.6151
R2090 B.n708 B.n707 10.6151
R2091 B.n707 B.n38 10.6151
R2092 B.n701 B.n38 10.6151
R2093 B.n701 B.n700 10.6151
R2094 B.n700 B.n699 10.6151
R2095 B.n699 B.n44 10.6151
R2096 B.n693 B.n44 10.6151
R2097 B.n693 B.n692 10.6151
R2098 B.n692 B.n691 10.6151
R2099 B.n182 B.n105 9.36635
R2100 B.n205 B.n102 9.36635
R2101 B.n461 B.n460 9.36635
R2102 B.n481 B.n355 9.36635
R2103 B.n747 B.n0 2.81026
R2104 B.n747 B.n1 2.81026
R2105 B.n185 B.n105 1.24928
R2106 B.n202 B.n102 1.24928
R2107 B.n462 B.n461 1.24928
R2108 B.n482 B.n481 1.24928
R2109 VN.n4 VN.t4 326.95
R2110 VN.n19 VN.t5 326.95
R2111 VN.n13 VN.t3 310.702
R2112 VN.n28 VN.t7 310.702
R2113 VN.n3 VN.t6 272.188
R2114 VN.n1 VN.t0 272.188
R2115 VN.n18 VN.t2 272.188
R2116 VN.n16 VN.t1 272.188
R2117 VN.n14 VN.n13 161.3
R2118 VN.n29 VN.n28 161.3
R2119 VN.n27 VN.n15 161.3
R2120 VN.n26 VN.n25 161.3
R2121 VN.n24 VN.n23 161.3
R2122 VN.n22 VN.n17 161.3
R2123 VN.n21 VN.n20 161.3
R2124 VN.n12 VN.n0 161.3
R2125 VN.n11 VN.n10 161.3
R2126 VN.n9 VN.n8 161.3
R2127 VN.n7 VN.n2 161.3
R2128 VN.n6 VN.n5 161.3
R2129 VN.n12 VN.n11 55.1086
R2130 VN.n27 VN.n26 55.1086
R2131 VN.n4 VN.n3 46.4196
R2132 VN.n19 VN.n18 46.4196
R2133 VN.n20 VN.n19 43.7016
R2134 VN.n5 VN.n4 43.7016
R2135 VN VN.n29 43.5706
R2136 VN.n7 VN.n6 40.577
R2137 VN.n8 VN.n7 40.577
R2138 VN.n22 VN.n21 40.577
R2139 VN.n23 VN.n22 40.577
R2140 VN.n11 VN.n1 15.9852
R2141 VN.n26 VN.n16 15.9852
R2142 VN.n6 VN.n3 8.60764
R2143 VN.n8 VN.n1 8.60764
R2144 VN.n21 VN.n18 8.60764
R2145 VN.n23 VN.n16 8.60764
R2146 VN.n13 VN.n12 2.19141
R2147 VN.n28 VN.n27 2.19141
R2148 VN.n29 VN.n15 0.189894
R2149 VN.n25 VN.n15 0.189894
R2150 VN.n25 VN.n24 0.189894
R2151 VN.n24 VN.n17 0.189894
R2152 VN.n20 VN.n17 0.189894
R2153 VN.n5 VN.n2 0.189894
R2154 VN.n9 VN.n2 0.189894
R2155 VN.n10 VN.n9 0.189894
R2156 VN.n10 VN.n0 0.189894
R2157 VN.n14 VN.n0 0.189894
R2158 VN VN.n14 0.0516364
R2159 VDD2.n2 VDD2.n1 64.9436
R2160 VDD2.n2 VDD2.n0 64.9436
R2161 VDD2 VDD2.n5 64.9407
R2162 VDD2.n4 VDD2.n3 64.4172
R2163 VDD2.n4 VDD2.n2 38.8834
R2164 VDD2.n5 VDD2.t5 1.71925
R2165 VDD2.n5 VDD2.t2 1.71925
R2166 VDD2.n3 VDD2.t0 1.71925
R2167 VDD2.n3 VDD2.t6 1.71925
R2168 VDD2.n1 VDD2.t7 1.71925
R2169 VDD2.n1 VDD2.t4 1.71925
R2170 VDD2.n0 VDD2.t3 1.71925
R2171 VDD2.n0 VDD2.t1 1.71925
R2172 VDD2 VDD2.n4 0.640586
C0 VN VDD2 6.31802f
C1 VP VTAIL 6.24387f
C2 VDD1 VP 6.52009f
C3 VN VTAIL 6.22976f
C4 VDD1 VN 0.149186f
C5 VTAIL VDD2 9.26253f
C6 VDD1 VDD2 0.985761f
C7 VN VP 5.6345f
C8 VP VDD2 0.351857f
C9 VDD1 VTAIL 9.21871f
C10 VDD2 B 3.761202f
C11 VDD1 B 4.027636f
C12 VTAIL B 8.962445f
C13 VN B 9.603939f
C14 VP B 7.844721f
C15 VDD2.t3 B 0.235759f
C16 VDD2.t1 B 0.235759f
C17 VDD2.n0 B 2.10062f
C18 VDD2.t7 B 0.235759f
C19 VDD2.t4 B 0.235759f
C20 VDD2.n1 B 2.10062f
C21 VDD2.n2 B 2.41003f
C22 VDD2.t0 B 0.235759f
C23 VDD2.t6 B 0.235759f
C24 VDD2.n3 B 2.09768f
C25 VDD2.n4 B 2.44741f
C26 VDD2.t5 B 0.235759f
C27 VDD2.t2 B 0.235759f
C28 VDD2.n5 B 2.1006f
C29 VN.n0 B 0.03757f
C30 VN.t0 B 1.20138f
C31 VN.n1 B 0.446788f
C32 VN.n2 B 0.03757f
C33 VN.t6 B 1.20138f
C34 VN.n3 B 0.481478f
C35 VN.t4 B 1.28492f
C36 VN.n4 B 0.501053f
C37 VN.n5 B 0.162671f
C38 VN.n6 B 0.05192f
C39 VN.n7 B 0.030344f
C40 VN.n8 B 0.05192f
C41 VN.n9 B 0.03757f
C42 VN.n10 B 0.03757f
C43 VN.n11 B 0.05268f
C44 VN.n12 B 0.011831f
C45 VN.t3 B 1.25973f
C46 VN.n13 B 0.4956f
C47 VN.n14 B 0.029115f
C48 VN.n15 B 0.03757f
C49 VN.t1 B 1.20138f
C50 VN.n16 B 0.446788f
C51 VN.n17 B 0.03757f
C52 VN.t2 B 1.20138f
C53 VN.n18 B 0.481478f
C54 VN.t5 B 1.28492f
C55 VN.n19 B 0.501053f
C56 VN.n20 B 0.162671f
C57 VN.n21 B 0.05192f
C58 VN.n22 B 0.030344f
C59 VN.n23 B 0.05192f
C60 VN.n24 B 0.03757f
C61 VN.n25 B 0.03757f
C62 VN.n26 B 0.05268f
C63 VN.n27 B 0.011831f
C64 VN.t7 B 1.25973f
C65 VN.n28 B 0.4956f
C66 VN.n29 B 1.64855f
C67 VTAIL.t4 B 0.177082f
C68 VTAIL.t5 B 0.177082f
C69 VTAIL.n0 B 1.52138f
C70 VTAIL.n1 B 0.263234f
C71 VTAIL.n2 B 0.028392f
C72 VTAIL.n3 B 0.019452f
C73 VTAIL.n4 B 0.010453f
C74 VTAIL.n5 B 0.024706f
C75 VTAIL.n6 B 0.011068f
C76 VTAIL.n7 B 0.019452f
C77 VTAIL.n8 B 0.010453f
C78 VTAIL.n9 B 0.024706f
C79 VTAIL.n10 B 0.01076f
C80 VTAIL.n11 B 0.019452f
C81 VTAIL.n12 B 0.011068f
C82 VTAIL.n13 B 0.024706f
C83 VTAIL.n14 B 0.011068f
C84 VTAIL.n15 B 0.019452f
C85 VTAIL.n16 B 0.010453f
C86 VTAIL.n17 B 0.024706f
C87 VTAIL.n18 B 0.011068f
C88 VTAIL.n19 B 0.939798f
C89 VTAIL.n20 B 0.010453f
C90 VTAIL.t3 B 0.041678f
C91 VTAIL.n21 B 0.136664f
C92 VTAIL.n22 B 0.017466f
C93 VTAIL.n23 B 0.01853f
C94 VTAIL.n24 B 0.024706f
C95 VTAIL.n25 B 0.011068f
C96 VTAIL.n26 B 0.010453f
C97 VTAIL.n27 B 0.019452f
C98 VTAIL.n28 B 0.019452f
C99 VTAIL.n29 B 0.010453f
C100 VTAIL.n30 B 0.011068f
C101 VTAIL.n31 B 0.024706f
C102 VTAIL.n32 B 0.024706f
C103 VTAIL.n33 B 0.011068f
C104 VTAIL.n34 B 0.010453f
C105 VTAIL.n35 B 0.019452f
C106 VTAIL.n36 B 0.019452f
C107 VTAIL.n37 B 0.010453f
C108 VTAIL.n38 B 0.010453f
C109 VTAIL.n39 B 0.011068f
C110 VTAIL.n40 B 0.024706f
C111 VTAIL.n41 B 0.024706f
C112 VTAIL.n42 B 0.024706f
C113 VTAIL.n43 B 0.01076f
C114 VTAIL.n44 B 0.010453f
C115 VTAIL.n45 B 0.019452f
C116 VTAIL.n46 B 0.019452f
C117 VTAIL.n47 B 0.010453f
C118 VTAIL.n48 B 0.011068f
C119 VTAIL.n49 B 0.024706f
C120 VTAIL.n50 B 0.024706f
C121 VTAIL.n51 B 0.011068f
C122 VTAIL.n52 B 0.010453f
C123 VTAIL.n53 B 0.019452f
C124 VTAIL.n54 B 0.019452f
C125 VTAIL.n55 B 0.010453f
C126 VTAIL.n56 B 0.011068f
C127 VTAIL.n57 B 0.024706f
C128 VTAIL.n58 B 0.055342f
C129 VTAIL.n59 B 0.011068f
C130 VTAIL.n60 B 0.010453f
C131 VTAIL.n61 B 0.048152f
C132 VTAIL.n62 B 0.031252f
C133 VTAIL.n63 B 0.12081f
C134 VTAIL.n64 B 0.028392f
C135 VTAIL.n65 B 0.019452f
C136 VTAIL.n66 B 0.010453f
C137 VTAIL.n67 B 0.024706f
C138 VTAIL.n68 B 0.011068f
C139 VTAIL.n69 B 0.019452f
C140 VTAIL.n70 B 0.010453f
C141 VTAIL.n71 B 0.024706f
C142 VTAIL.n72 B 0.01076f
C143 VTAIL.n73 B 0.019452f
C144 VTAIL.n74 B 0.011068f
C145 VTAIL.n75 B 0.024706f
C146 VTAIL.n76 B 0.011068f
C147 VTAIL.n77 B 0.019452f
C148 VTAIL.n78 B 0.010453f
C149 VTAIL.n79 B 0.024706f
C150 VTAIL.n80 B 0.011068f
C151 VTAIL.n81 B 0.939798f
C152 VTAIL.n82 B 0.010453f
C153 VTAIL.t10 B 0.041678f
C154 VTAIL.n83 B 0.136664f
C155 VTAIL.n84 B 0.017466f
C156 VTAIL.n85 B 0.01853f
C157 VTAIL.n86 B 0.024706f
C158 VTAIL.n87 B 0.011068f
C159 VTAIL.n88 B 0.010453f
C160 VTAIL.n89 B 0.019452f
C161 VTAIL.n90 B 0.019452f
C162 VTAIL.n91 B 0.010453f
C163 VTAIL.n92 B 0.011068f
C164 VTAIL.n93 B 0.024706f
C165 VTAIL.n94 B 0.024706f
C166 VTAIL.n95 B 0.011068f
C167 VTAIL.n96 B 0.010453f
C168 VTAIL.n97 B 0.019452f
C169 VTAIL.n98 B 0.019452f
C170 VTAIL.n99 B 0.010453f
C171 VTAIL.n100 B 0.010453f
C172 VTAIL.n101 B 0.011068f
C173 VTAIL.n102 B 0.024706f
C174 VTAIL.n103 B 0.024706f
C175 VTAIL.n104 B 0.024706f
C176 VTAIL.n105 B 0.01076f
C177 VTAIL.n106 B 0.010453f
C178 VTAIL.n107 B 0.019452f
C179 VTAIL.n108 B 0.019452f
C180 VTAIL.n109 B 0.010453f
C181 VTAIL.n110 B 0.011068f
C182 VTAIL.n111 B 0.024706f
C183 VTAIL.n112 B 0.024706f
C184 VTAIL.n113 B 0.011068f
C185 VTAIL.n114 B 0.010453f
C186 VTAIL.n115 B 0.019452f
C187 VTAIL.n116 B 0.019452f
C188 VTAIL.n117 B 0.010453f
C189 VTAIL.n118 B 0.011068f
C190 VTAIL.n119 B 0.024706f
C191 VTAIL.n120 B 0.055342f
C192 VTAIL.n121 B 0.011068f
C193 VTAIL.n122 B 0.010453f
C194 VTAIL.n123 B 0.048152f
C195 VTAIL.n124 B 0.031252f
C196 VTAIL.n125 B 0.12081f
C197 VTAIL.t12 B 0.177082f
C198 VTAIL.t14 B 0.177082f
C199 VTAIL.n126 B 1.52138f
C200 VTAIL.n127 B 0.332533f
C201 VTAIL.n128 B 0.028392f
C202 VTAIL.n129 B 0.019452f
C203 VTAIL.n130 B 0.010453f
C204 VTAIL.n131 B 0.024706f
C205 VTAIL.n132 B 0.011068f
C206 VTAIL.n133 B 0.019452f
C207 VTAIL.n134 B 0.010453f
C208 VTAIL.n135 B 0.024706f
C209 VTAIL.n136 B 0.01076f
C210 VTAIL.n137 B 0.019452f
C211 VTAIL.n138 B 0.011068f
C212 VTAIL.n139 B 0.024706f
C213 VTAIL.n140 B 0.011068f
C214 VTAIL.n141 B 0.019452f
C215 VTAIL.n142 B 0.010453f
C216 VTAIL.n143 B 0.024706f
C217 VTAIL.n144 B 0.011068f
C218 VTAIL.n145 B 0.939798f
C219 VTAIL.n146 B 0.010453f
C220 VTAIL.t9 B 0.041678f
C221 VTAIL.n147 B 0.136664f
C222 VTAIL.n148 B 0.017466f
C223 VTAIL.n149 B 0.01853f
C224 VTAIL.n150 B 0.024706f
C225 VTAIL.n151 B 0.011068f
C226 VTAIL.n152 B 0.010453f
C227 VTAIL.n153 B 0.019452f
C228 VTAIL.n154 B 0.019452f
C229 VTAIL.n155 B 0.010453f
C230 VTAIL.n156 B 0.011068f
C231 VTAIL.n157 B 0.024706f
C232 VTAIL.n158 B 0.024706f
C233 VTAIL.n159 B 0.011068f
C234 VTAIL.n160 B 0.010453f
C235 VTAIL.n161 B 0.019452f
C236 VTAIL.n162 B 0.019452f
C237 VTAIL.n163 B 0.010453f
C238 VTAIL.n164 B 0.010453f
C239 VTAIL.n165 B 0.011068f
C240 VTAIL.n166 B 0.024706f
C241 VTAIL.n167 B 0.024706f
C242 VTAIL.n168 B 0.024706f
C243 VTAIL.n169 B 0.01076f
C244 VTAIL.n170 B 0.010453f
C245 VTAIL.n171 B 0.019452f
C246 VTAIL.n172 B 0.019452f
C247 VTAIL.n173 B 0.010453f
C248 VTAIL.n174 B 0.011068f
C249 VTAIL.n175 B 0.024706f
C250 VTAIL.n176 B 0.024706f
C251 VTAIL.n177 B 0.011068f
C252 VTAIL.n178 B 0.010453f
C253 VTAIL.n179 B 0.019452f
C254 VTAIL.n180 B 0.019452f
C255 VTAIL.n181 B 0.010453f
C256 VTAIL.n182 B 0.011068f
C257 VTAIL.n183 B 0.024706f
C258 VTAIL.n184 B 0.055342f
C259 VTAIL.n185 B 0.011068f
C260 VTAIL.n186 B 0.010453f
C261 VTAIL.n187 B 0.048152f
C262 VTAIL.n188 B 0.031252f
C263 VTAIL.n189 B 1.05101f
C264 VTAIL.n190 B 0.028392f
C265 VTAIL.n191 B 0.019452f
C266 VTAIL.n192 B 0.010453f
C267 VTAIL.n193 B 0.024706f
C268 VTAIL.n194 B 0.011068f
C269 VTAIL.n195 B 0.019452f
C270 VTAIL.n196 B 0.010453f
C271 VTAIL.n197 B 0.024706f
C272 VTAIL.n198 B 0.01076f
C273 VTAIL.n199 B 0.019452f
C274 VTAIL.n200 B 0.01076f
C275 VTAIL.n201 B 0.010453f
C276 VTAIL.n202 B 0.024706f
C277 VTAIL.n203 B 0.024706f
C278 VTAIL.n204 B 0.011068f
C279 VTAIL.n205 B 0.019452f
C280 VTAIL.n206 B 0.010453f
C281 VTAIL.n207 B 0.024706f
C282 VTAIL.n208 B 0.011068f
C283 VTAIL.n209 B 0.939798f
C284 VTAIL.n210 B 0.010453f
C285 VTAIL.t0 B 0.041678f
C286 VTAIL.n211 B 0.136664f
C287 VTAIL.n212 B 0.017466f
C288 VTAIL.n213 B 0.01853f
C289 VTAIL.n214 B 0.024706f
C290 VTAIL.n215 B 0.011068f
C291 VTAIL.n216 B 0.010453f
C292 VTAIL.n217 B 0.019452f
C293 VTAIL.n218 B 0.019452f
C294 VTAIL.n219 B 0.010453f
C295 VTAIL.n220 B 0.011068f
C296 VTAIL.n221 B 0.024706f
C297 VTAIL.n222 B 0.024706f
C298 VTAIL.n223 B 0.011068f
C299 VTAIL.n224 B 0.010453f
C300 VTAIL.n225 B 0.019452f
C301 VTAIL.n226 B 0.019452f
C302 VTAIL.n227 B 0.010453f
C303 VTAIL.n228 B 0.011068f
C304 VTAIL.n229 B 0.024706f
C305 VTAIL.n230 B 0.024706f
C306 VTAIL.n231 B 0.011068f
C307 VTAIL.n232 B 0.010453f
C308 VTAIL.n233 B 0.019452f
C309 VTAIL.n234 B 0.019452f
C310 VTAIL.n235 B 0.010453f
C311 VTAIL.n236 B 0.011068f
C312 VTAIL.n237 B 0.024706f
C313 VTAIL.n238 B 0.024706f
C314 VTAIL.n239 B 0.011068f
C315 VTAIL.n240 B 0.010453f
C316 VTAIL.n241 B 0.019452f
C317 VTAIL.n242 B 0.019452f
C318 VTAIL.n243 B 0.010453f
C319 VTAIL.n244 B 0.011068f
C320 VTAIL.n245 B 0.024706f
C321 VTAIL.n246 B 0.055342f
C322 VTAIL.n247 B 0.011068f
C323 VTAIL.n248 B 0.010453f
C324 VTAIL.n249 B 0.048152f
C325 VTAIL.n250 B 0.031252f
C326 VTAIL.n251 B 1.05101f
C327 VTAIL.t15 B 0.177082f
C328 VTAIL.t2 B 0.177082f
C329 VTAIL.n252 B 1.52139f
C330 VTAIL.n253 B 0.332524f
C331 VTAIL.n254 B 0.028392f
C332 VTAIL.n255 B 0.019452f
C333 VTAIL.n256 B 0.010453f
C334 VTAIL.n257 B 0.024706f
C335 VTAIL.n258 B 0.011068f
C336 VTAIL.n259 B 0.019452f
C337 VTAIL.n260 B 0.010453f
C338 VTAIL.n261 B 0.024706f
C339 VTAIL.n262 B 0.01076f
C340 VTAIL.n263 B 0.019452f
C341 VTAIL.n264 B 0.01076f
C342 VTAIL.n265 B 0.010453f
C343 VTAIL.n266 B 0.024706f
C344 VTAIL.n267 B 0.024706f
C345 VTAIL.n268 B 0.011068f
C346 VTAIL.n269 B 0.019452f
C347 VTAIL.n270 B 0.010453f
C348 VTAIL.n271 B 0.024706f
C349 VTAIL.n272 B 0.011068f
C350 VTAIL.n273 B 0.939798f
C351 VTAIL.n274 B 0.010453f
C352 VTAIL.t1 B 0.041678f
C353 VTAIL.n275 B 0.136664f
C354 VTAIL.n276 B 0.017466f
C355 VTAIL.n277 B 0.01853f
C356 VTAIL.n278 B 0.024706f
C357 VTAIL.n279 B 0.011068f
C358 VTAIL.n280 B 0.010453f
C359 VTAIL.n281 B 0.019452f
C360 VTAIL.n282 B 0.019452f
C361 VTAIL.n283 B 0.010453f
C362 VTAIL.n284 B 0.011068f
C363 VTAIL.n285 B 0.024706f
C364 VTAIL.n286 B 0.024706f
C365 VTAIL.n287 B 0.011068f
C366 VTAIL.n288 B 0.010453f
C367 VTAIL.n289 B 0.019452f
C368 VTAIL.n290 B 0.019452f
C369 VTAIL.n291 B 0.010453f
C370 VTAIL.n292 B 0.011068f
C371 VTAIL.n293 B 0.024706f
C372 VTAIL.n294 B 0.024706f
C373 VTAIL.n295 B 0.011068f
C374 VTAIL.n296 B 0.010453f
C375 VTAIL.n297 B 0.019452f
C376 VTAIL.n298 B 0.019452f
C377 VTAIL.n299 B 0.010453f
C378 VTAIL.n300 B 0.011068f
C379 VTAIL.n301 B 0.024706f
C380 VTAIL.n302 B 0.024706f
C381 VTAIL.n303 B 0.011068f
C382 VTAIL.n304 B 0.010453f
C383 VTAIL.n305 B 0.019452f
C384 VTAIL.n306 B 0.019452f
C385 VTAIL.n307 B 0.010453f
C386 VTAIL.n308 B 0.011068f
C387 VTAIL.n309 B 0.024706f
C388 VTAIL.n310 B 0.055342f
C389 VTAIL.n311 B 0.011068f
C390 VTAIL.n312 B 0.010453f
C391 VTAIL.n313 B 0.048152f
C392 VTAIL.n314 B 0.031252f
C393 VTAIL.n315 B 0.12081f
C394 VTAIL.n316 B 0.028392f
C395 VTAIL.n317 B 0.019452f
C396 VTAIL.n318 B 0.010453f
C397 VTAIL.n319 B 0.024706f
C398 VTAIL.n320 B 0.011068f
C399 VTAIL.n321 B 0.019452f
C400 VTAIL.n322 B 0.010453f
C401 VTAIL.n323 B 0.024706f
C402 VTAIL.n324 B 0.01076f
C403 VTAIL.n325 B 0.019452f
C404 VTAIL.n326 B 0.01076f
C405 VTAIL.n327 B 0.010453f
C406 VTAIL.n328 B 0.024706f
C407 VTAIL.n329 B 0.024706f
C408 VTAIL.n330 B 0.011068f
C409 VTAIL.n331 B 0.019452f
C410 VTAIL.n332 B 0.010453f
C411 VTAIL.n333 B 0.024706f
C412 VTAIL.n334 B 0.011068f
C413 VTAIL.n335 B 0.939798f
C414 VTAIL.n336 B 0.010453f
C415 VTAIL.t8 B 0.041678f
C416 VTAIL.n337 B 0.136664f
C417 VTAIL.n338 B 0.017466f
C418 VTAIL.n339 B 0.01853f
C419 VTAIL.n340 B 0.024706f
C420 VTAIL.n341 B 0.011068f
C421 VTAIL.n342 B 0.010453f
C422 VTAIL.n343 B 0.019452f
C423 VTAIL.n344 B 0.019452f
C424 VTAIL.n345 B 0.010453f
C425 VTAIL.n346 B 0.011068f
C426 VTAIL.n347 B 0.024706f
C427 VTAIL.n348 B 0.024706f
C428 VTAIL.n349 B 0.011068f
C429 VTAIL.n350 B 0.010453f
C430 VTAIL.n351 B 0.019452f
C431 VTAIL.n352 B 0.019452f
C432 VTAIL.n353 B 0.010453f
C433 VTAIL.n354 B 0.011068f
C434 VTAIL.n355 B 0.024706f
C435 VTAIL.n356 B 0.024706f
C436 VTAIL.n357 B 0.011068f
C437 VTAIL.n358 B 0.010453f
C438 VTAIL.n359 B 0.019452f
C439 VTAIL.n360 B 0.019452f
C440 VTAIL.n361 B 0.010453f
C441 VTAIL.n362 B 0.011068f
C442 VTAIL.n363 B 0.024706f
C443 VTAIL.n364 B 0.024706f
C444 VTAIL.n365 B 0.011068f
C445 VTAIL.n366 B 0.010453f
C446 VTAIL.n367 B 0.019452f
C447 VTAIL.n368 B 0.019452f
C448 VTAIL.n369 B 0.010453f
C449 VTAIL.n370 B 0.011068f
C450 VTAIL.n371 B 0.024706f
C451 VTAIL.n372 B 0.055342f
C452 VTAIL.n373 B 0.011068f
C453 VTAIL.n374 B 0.010453f
C454 VTAIL.n375 B 0.048152f
C455 VTAIL.n376 B 0.031252f
C456 VTAIL.n377 B 0.12081f
C457 VTAIL.t11 B 0.177082f
C458 VTAIL.t13 B 0.177082f
C459 VTAIL.n378 B 1.52139f
C460 VTAIL.n379 B 0.332524f
C461 VTAIL.n380 B 0.028392f
C462 VTAIL.n381 B 0.019452f
C463 VTAIL.n382 B 0.010453f
C464 VTAIL.n383 B 0.024706f
C465 VTAIL.n384 B 0.011068f
C466 VTAIL.n385 B 0.019452f
C467 VTAIL.n386 B 0.010453f
C468 VTAIL.n387 B 0.024706f
C469 VTAIL.n388 B 0.01076f
C470 VTAIL.n389 B 0.019452f
C471 VTAIL.n390 B 0.01076f
C472 VTAIL.n391 B 0.010453f
C473 VTAIL.n392 B 0.024706f
C474 VTAIL.n393 B 0.024706f
C475 VTAIL.n394 B 0.011068f
C476 VTAIL.n395 B 0.019452f
C477 VTAIL.n396 B 0.010453f
C478 VTAIL.n397 B 0.024706f
C479 VTAIL.n398 B 0.011068f
C480 VTAIL.n399 B 0.939798f
C481 VTAIL.n400 B 0.010453f
C482 VTAIL.t7 B 0.041678f
C483 VTAIL.n401 B 0.136664f
C484 VTAIL.n402 B 0.017466f
C485 VTAIL.n403 B 0.01853f
C486 VTAIL.n404 B 0.024706f
C487 VTAIL.n405 B 0.011068f
C488 VTAIL.n406 B 0.010453f
C489 VTAIL.n407 B 0.019452f
C490 VTAIL.n408 B 0.019452f
C491 VTAIL.n409 B 0.010453f
C492 VTAIL.n410 B 0.011068f
C493 VTAIL.n411 B 0.024706f
C494 VTAIL.n412 B 0.024706f
C495 VTAIL.n413 B 0.011068f
C496 VTAIL.n414 B 0.010453f
C497 VTAIL.n415 B 0.019452f
C498 VTAIL.n416 B 0.019452f
C499 VTAIL.n417 B 0.010453f
C500 VTAIL.n418 B 0.011068f
C501 VTAIL.n419 B 0.024706f
C502 VTAIL.n420 B 0.024706f
C503 VTAIL.n421 B 0.011068f
C504 VTAIL.n422 B 0.010453f
C505 VTAIL.n423 B 0.019452f
C506 VTAIL.n424 B 0.019452f
C507 VTAIL.n425 B 0.010453f
C508 VTAIL.n426 B 0.011068f
C509 VTAIL.n427 B 0.024706f
C510 VTAIL.n428 B 0.024706f
C511 VTAIL.n429 B 0.011068f
C512 VTAIL.n430 B 0.010453f
C513 VTAIL.n431 B 0.019452f
C514 VTAIL.n432 B 0.019452f
C515 VTAIL.n433 B 0.010453f
C516 VTAIL.n434 B 0.011068f
C517 VTAIL.n435 B 0.024706f
C518 VTAIL.n436 B 0.055342f
C519 VTAIL.n437 B 0.011068f
C520 VTAIL.n438 B 0.010453f
C521 VTAIL.n439 B 0.048152f
C522 VTAIL.n440 B 0.031252f
C523 VTAIL.n441 B 1.05101f
C524 VTAIL.n442 B 0.028392f
C525 VTAIL.n443 B 0.019452f
C526 VTAIL.n444 B 0.010453f
C527 VTAIL.n445 B 0.024706f
C528 VTAIL.n446 B 0.011068f
C529 VTAIL.n447 B 0.019452f
C530 VTAIL.n448 B 0.010453f
C531 VTAIL.n449 B 0.024706f
C532 VTAIL.n450 B 0.01076f
C533 VTAIL.n451 B 0.019452f
C534 VTAIL.n452 B 0.011068f
C535 VTAIL.n453 B 0.024706f
C536 VTAIL.n454 B 0.011068f
C537 VTAIL.n455 B 0.019452f
C538 VTAIL.n456 B 0.010453f
C539 VTAIL.n457 B 0.024706f
C540 VTAIL.n458 B 0.011068f
C541 VTAIL.n459 B 0.939798f
C542 VTAIL.n460 B 0.010453f
C543 VTAIL.t6 B 0.041678f
C544 VTAIL.n461 B 0.136664f
C545 VTAIL.n462 B 0.017466f
C546 VTAIL.n463 B 0.01853f
C547 VTAIL.n464 B 0.024706f
C548 VTAIL.n465 B 0.011068f
C549 VTAIL.n466 B 0.010453f
C550 VTAIL.n467 B 0.019452f
C551 VTAIL.n468 B 0.019452f
C552 VTAIL.n469 B 0.010453f
C553 VTAIL.n470 B 0.011068f
C554 VTAIL.n471 B 0.024706f
C555 VTAIL.n472 B 0.024706f
C556 VTAIL.n473 B 0.011068f
C557 VTAIL.n474 B 0.010453f
C558 VTAIL.n475 B 0.019452f
C559 VTAIL.n476 B 0.019452f
C560 VTAIL.n477 B 0.010453f
C561 VTAIL.n478 B 0.010453f
C562 VTAIL.n479 B 0.011068f
C563 VTAIL.n480 B 0.024706f
C564 VTAIL.n481 B 0.024706f
C565 VTAIL.n482 B 0.024706f
C566 VTAIL.n483 B 0.01076f
C567 VTAIL.n484 B 0.010453f
C568 VTAIL.n485 B 0.019452f
C569 VTAIL.n486 B 0.019452f
C570 VTAIL.n487 B 0.010453f
C571 VTAIL.n488 B 0.011068f
C572 VTAIL.n489 B 0.024706f
C573 VTAIL.n490 B 0.024706f
C574 VTAIL.n491 B 0.011068f
C575 VTAIL.n492 B 0.010453f
C576 VTAIL.n493 B 0.019452f
C577 VTAIL.n494 B 0.019452f
C578 VTAIL.n495 B 0.010453f
C579 VTAIL.n496 B 0.011068f
C580 VTAIL.n497 B 0.024706f
C581 VTAIL.n498 B 0.055342f
C582 VTAIL.n499 B 0.011068f
C583 VTAIL.n500 B 0.010453f
C584 VTAIL.n501 B 0.048152f
C585 VTAIL.n502 B 0.031252f
C586 VTAIL.n503 B 1.04736f
C587 VDD1.t4 B 0.235825f
C588 VDD1.t2 B 0.235825f
C589 VDD1.n0 B 2.10193f
C590 VDD1.t0 B 0.235825f
C591 VDD1.t5 B 0.235825f
C592 VDD1.n1 B 2.10121f
C593 VDD1.t1 B 0.235825f
C594 VDD1.t6 B 0.235825f
C595 VDD1.n2 B 2.10121f
C596 VDD1.n3 B 2.46575f
C597 VDD1.t3 B 0.235825f
C598 VDD1.t7 B 0.235825f
C599 VDD1.n4 B 2.09825f
C600 VDD1.n5 B 2.47902f
C601 VP.n0 B 0.038096f
C602 VP.t0 B 1.21821f
C603 VP.n1 B 0.453047f
C604 VP.n2 B 0.038096f
C605 VP.t2 B 1.21821f
C606 VP.n3 B 0.453047f
C607 VP.n4 B 0.038096f
C608 VP.n5 B 0.038096f
C609 VP.t7 B 1.27738f
C610 VP.t1 B 1.21821f
C611 VP.n6 B 0.453047f
C612 VP.n7 B 0.038096f
C613 VP.t3 B 1.21821f
C614 VP.n8 B 0.488222f
C615 VP.t6 B 1.30292f
C616 VP.n9 B 0.508072f
C617 VP.n10 B 0.164949f
C618 VP.n11 B 0.052648f
C619 VP.n12 B 0.030769f
C620 VP.n13 B 0.052648f
C621 VP.n14 B 0.038096f
C622 VP.n15 B 0.038096f
C623 VP.n16 B 0.053418f
C624 VP.n17 B 0.011997f
C625 VP.n18 B 0.502543f
C626 VP.n19 B 1.64668f
C627 VP.n20 B 1.67848f
C628 VP.t5 B 1.27738f
C629 VP.n21 B 0.502543f
C630 VP.n22 B 0.011997f
C631 VP.n23 B 0.053418f
C632 VP.n24 B 0.038096f
C633 VP.n25 B 0.038096f
C634 VP.n26 B 0.052648f
C635 VP.n27 B 0.030769f
C636 VP.n28 B 0.052648f
C637 VP.n29 B 0.038096f
C638 VP.n30 B 0.038096f
C639 VP.n31 B 0.053418f
C640 VP.n32 B 0.011997f
C641 VP.t4 B 1.27738f
C642 VP.n33 B 0.502543f
C643 VP.n34 B 0.029523f
.ends

