* NGSPICE file created from diff_pair_sample_1650.ext - technology: sky130A

.subckt diff_pair_sample_1650 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.58
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.58
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0.6357 ps=4.04 w=1.63 l=2.58
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0.6357 ps=4.04 w=1.63 l=2.58
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.58
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0.6357 ps=4.04 w=1.63 l=2.58
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0.6357 ps=4.04 w=1.63 l=2.58
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6357 pd=4.04 as=0 ps=0 w=1.63 l=2.58
R0 B.n373 B.n372 585
R1 B.n131 B.n64 585
R2 B.n130 B.n129 585
R3 B.n128 B.n127 585
R4 B.n126 B.n125 585
R5 B.n124 B.n123 585
R6 B.n122 B.n121 585
R7 B.n120 B.n119 585
R8 B.n118 B.n117 585
R9 B.n116 B.n115 585
R10 B.n114 B.n113 585
R11 B.n111 B.n110 585
R12 B.n109 B.n108 585
R13 B.n107 B.n106 585
R14 B.n105 B.n104 585
R15 B.n103 B.n102 585
R16 B.n101 B.n100 585
R17 B.n99 B.n98 585
R18 B.n97 B.n96 585
R19 B.n95 B.n94 585
R20 B.n93 B.n92 585
R21 B.n90 B.n89 585
R22 B.n88 B.n87 585
R23 B.n86 B.n85 585
R24 B.n84 B.n83 585
R25 B.n82 B.n81 585
R26 B.n80 B.n79 585
R27 B.n78 B.n77 585
R28 B.n76 B.n75 585
R29 B.n74 B.n73 585
R30 B.n72 B.n71 585
R31 B.n70 B.n69 585
R32 B.n371 B.n48 585
R33 B.n376 B.n48 585
R34 B.n370 B.n47 585
R35 B.n377 B.n47 585
R36 B.n369 B.n368 585
R37 B.n368 B.n43 585
R38 B.n367 B.n42 585
R39 B.n383 B.n42 585
R40 B.n366 B.n41 585
R41 B.n384 B.n41 585
R42 B.n365 B.n40 585
R43 B.n385 B.n40 585
R44 B.n364 B.n363 585
R45 B.n363 B.n36 585
R46 B.n362 B.n35 585
R47 B.n391 B.n35 585
R48 B.n361 B.n34 585
R49 B.n392 B.n34 585
R50 B.n360 B.n33 585
R51 B.n393 B.n33 585
R52 B.n359 B.n358 585
R53 B.n358 B.n29 585
R54 B.n357 B.n28 585
R55 B.n399 B.n28 585
R56 B.n356 B.n27 585
R57 B.n400 B.n27 585
R58 B.n355 B.n26 585
R59 B.n401 B.n26 585
R60 B.n354 B.n353 585
R61 B.n353 B.n22 585
R62 B.n352 B.n21 585
R63 B.n407 B.n21 585
R64 B.n351 B.n20 585
R65 B.n408 B.n20 585
R66 B.n350 B.n19 585
R67 B.n409 B.n19 585
R68 B.n349 B.n348 585
R69 B.n348 B.n15 585
R70 B.n347 B.n14 585
R71 B.n415 B.n14 585
R72 B.n346 B.n13 585
R73 B.n416 B.n13 585
R74 B.n345 B.n12 585
R75 B.n417 B.n12 585
R76 B.n344 B.n343 585
R77 B.n343 B.n8 585
R78 B.n342 B.n7 585
R79 B.n423 B.n7 585
R80 B.n341 B.n6 585
R81 B.n424 B.n6 585
R82 B.n340 B.n5 585
R83 B.n425 B.n5 585
R84 B.n339 B.n338 585
R85 B.n338 B.n4 585
R86 B.n337 B.n132 585
R87 B.n337 B.n336 585
R88 B.n327 B.n133 585
R89 B.n134 B.n133 585
R90 B.n329 B.n328 585
R91 B.n330 B.n329 585
R92 B.n326 B.n139 585
R93 B.n139 B.n138 585
R94 B.n325 B.n324 585
R95 B.n324 B.n323 585
R96 B.n141 B.n140 585
R97 B.n142 B.n141 585
R98 B.n316 B.n315 585
R99 B.n317 B.n316 585
R100 B.n314 B.n147 585
R101 B.n147 B.n146 585
R102 B.n313 B.n312 585
R103 B.n312 B.n311 585
R104 B.n149 B.n148 585
R105 B.n150 B.n149 585
R106 B.n304 B.n303 585
R107 B.n305 B.n304 585
R108 B.n302 B.n155 585
R109 B.n155 B.n154 585
R110 B.n301 B.n300 585
R111 B.n300 B.n299 585
R112 B.n157 B.n156 585
R113 B.n158 B.n157 585
R114 B.n292 B.n291 585
R115 B.n293 B.n292 585
R116 B.n290 B.n163 585
R117 B.n163 B.n162 585
R118 B.n289 B.n288 585
R119 B.n288 B.n287 585
R120 B.n165 B.n164 585
R121 B.n166 B.n165 585
R122 B.n280 B.n279 585
R123 B.n281 B.n280 585
R124 B.n278 B.n171 585
R125 B.n171 B.n170 585
R126 B.n277 B.n276 585
R127 B.n276 B.n275 585
R128 B.n173 B.n172 585
R129 B.n174 B.n173 585
R130 B.n268 B.n267 585
R131 B.n269 B.n268 585
R132 B.n266 B.n179 585
R133 B.n179 B.n178 585
R134 B.n261 B.n260 585
R135 B.n259 B.n197 585
R136 B.n258 B.n196 585
R137 B.n263 B.n196 585
R138 B.n257 B.n256 585
R139 B.n255 B.n254 585
R140 B.n253 B.n252 585
R141 B.n251 B.n250 585
R142 B.n249 B.n248 585
R143 B.n247 B.n246 585
R144 B.n245 B.n244 585
R145 B.n243 B.n242 585
R146 B.n241 B.n240 585
R147 B.n239 B.n238 585
R148 B.n237 B.n236 585
R149 B.n235 B.n234 585
R150 B.n233 B.n232 585
R151 B.n231 B.n230 585
R152 B.n229 B.n228 585
R153 B.n227 B.n226 585
R154 B.n225 B.n224 585
R155 B.n223 B.n222 585
R156 B.n221 B.n220 585
R157 B.n219 B.n218 585
R158 B.n217 B.n216 585
R159 B.n215 B.n214 585
R160 B.n213 B.n212 585
R161 B.n211 B.n210 585
R162 B.n209 B.n208 585
R163 B.n207 B.n206 585
R164 B.n205 B.n204 585
R165 B.n181 B.n180 585
R166 B.n265 B.n264 585
R167 B.n264 B.n263 585
R168 B.n177 B.n176 585
R169 B.n178 B.n177 585
R170 B.n271 B.n270 585
R171 B.n270 B.n269 585
R172 B.n272 B.n175 585
R173 B.n175 B.n174 585
R174 B.n274 B.n273 585
R175 B.n275 B.n274 585
R176 B.n169 B.n168 585
R177 B.n170 B.n169 585
R178 B.n283 B.n282 585
R179 B.n282 B.n281 585
R180 B.n284 B.n167 585
R181 B.n167 B.n166 585
R182 B.n286 B.n285 585
R183 B.n287 B.n286 585
R184 B.n161 B.n160 585
R185 B.n162 B.n161 585
R186 B.n295 B.n294 585
R187 B.n294 B.n293 585
R188 B.n296 B.n159 585
R189 B.n159 B.n158 585
R190 B.n298 B.n297 585
R191 B.n299 B.n298 585
R192 B.n153 B.n152 585
R193 B.n154 B.n153 585
R194 B.n307 B.n306 585
R195 B.n306 B.n305 585
R196 B.n308 B.n151 585
R197 B.n151 B.n150 585
R198 B.n310 B.n309 585
R199 B.n311 B.n310 585
R200 B.n145 B.n144 585
R201 B.n146 B.n145 585
R202 B.n319 B.n318 585
R203 B.n318 B.n317 585
R204 B.n320 B.n143 585
R205 B.n143 B.n142 585
R206 B.n322 B.n321 585
R207 B.n323 B.n322 585
R208 B.n137 B.n136 585
R209 B.n138 B.n137 585
R210 B.n332 B.n331 585
R211 B.n331 B.n330 585
R212 B.n333 B.n135 585
R213 B.n135 B.n134 585
R214 B.n335 B.n334 585
R215 B.n336 B.n335 585
R216 B.n2 B.n0 585
R217 B.n4 B.n2 585
R218 B.n3 B.n1 585
R219 B.n424 B.n3 585
R220 B.n422 B.n421 585
R221 B.n423 B.n422 585
R222 B.n420 B.n9 585
R223 B.n9 B.n8 585
R224 B.n419 B.n418 585
R225 B.n418 B.n417 585
R226 B.n11 B.n10 585
R227 B.n416 B.n11 585
R228 B.n414 B.n413 585
R229 B.n415 B.n414 585
R230 B.n412 B.n16 585
R231 B.n16 B.n15 585
R232 B.n411 B.n410 585
R233 B.n410 B.n409 585
R234 B.n18 B.n17 585
R235 B.n408 B.n18 585
R236 B.n406 B.n405 585
R237 B.n407 B.n406 585
R238 B.n404 B.n23 585
R239 B.n23 B.n22 585
R240 B.n403 B.n402 585
R241 B.n402 B.n401 585
R242 B.n25 B.n24 585
R243 B.n400 B.n25 585
R244 B.n398 B.n397 585
R245 B.n399 B.n398 585
R246 B.n396 B.n30 585
R247 B.n30 B.n29 585
R248 B.n395 B.n394 585
R249 B.n394 B.n393 585
R250 B.n32 B.n31 585
R251 B.n392 B.n32 585
R252 B.n390 B.n389 585
R253 B.n391 B.n390 585
R254 B.n388 B.n37 585
R255 B.n37 B.n36 585
R256 B.n387 B.n386 585
R257 B.n386 B.n385 585
R258 B.n39 B.n38 585
R259 B.n384 B.n39 585
R260 B.n382 B.n381 585
R261 B.n383 B.n382 585
R262 B.n380 B.n44 585
R263 B.n44 B.n43 585
R264 B.n379 B.n378 585
R265 B.n378 B.n377 585
R266 B.n46 B.n45 585
R267 B.n376 B.n46 585
R268 B.n427 B.n426 585
R269 B.n426 B.n425 585
R270 B.n261 B.n177 521.33
R271 B.n69 B.n46 521.33
R272 B.n264 B.n179 521.33
R273 B.n373 B.n48 521.33
R274 B.n375 B.n374 256.663
R275 B.n375 B.n63 256.663
R276 B.n375 B.n62 256.663
R277 B.n375 B.n61 256.663
R278 B.n375 B.n60 256.663
R279 B.n375 B.n59 256.663
R280 B.n375 B.n58 256.663
R281 B.n375 B.n57 256.663
R282 B.n375 B.n56 256.663
R283 B.n375 B.n55 256.663
R284 B.n375 B.n54 256.663
R285 B.n375 B.n53 256.663
R286 B.n375 B.n52 256.663
R287 B.n375 B.n51 256.663
R288 B.n375 B.n50 256.663
R289 B.n375 B.n49 256.663
R290 B.n263 B.n262 256.663
R291 B.n263 B.n182 256.663
R292 B.n263 B.n183 256.663
R293 B.n263 B.n184 256.663
R294 B.n263 B.n185 256.663
R295 B.n263 B.n186 256.663
R296 B.n263 B.n187 256.663
R297 B.n263 B.n188 256.663
R298 B.n263 B.n189 256.663
R299 B.n263 B.n190 256.663
R300 B.n263 B.n191 256.663
R301 B.n263 B.n192 256.663
R302 B.n263 B.n193 256.663
R303 B.n263 B.n194 256.663
R304 B.n263 B.n195 256.663
R305 B.n201 B.t6 223.243
R306 B.n198 B.t13 223.243
R307 B.n67 B.t10 223.243
R308 B.n65 B.t2 223.243
R309 B.n263 B.n178 221.435
R310 B.n376 B.n375 221.435
R311 B.n201 B.t9 165.244
R312 B.n65 B.t4 165.244
R313 B.n198 B.t15 165.244
R314 B.n67 B.t11 165.244
R315 B.n270 B.n177 163.367
R316 B.n270 B.n175 163.367
R317 B.n274 B.n175 163.367
R318 B.n274 B.n169 163.367
R319 B.n282 B.n169 163.367
R320 B.n282 B.n167 163.367
R321 B.n286 B.n167 163.367
R322 B.n286 B.n161 163.367
R323 B.n294 B.n161 163.367
R324 B.n294 B.n159 163.367
R325 B.n298 B.n159 163.367
R326 B.n298 B.n153 163.367
R327 B.n306 B.n153 163.367
R328 B.n306 B.n151 163.367
R329 B.n310 B.n151 163.367
R330 B.n310 B.n145 163.367
R331 B.n318 B.n145 163.367
R332 B.n318 B.n143 163.367
R333 B.n322 B.n143 163.367
R334 B.n322 B.n137 163.367
R335 B.n331 B.n137 163.367
R336 B.n331 B.n135 163.367
R337 B.n335 B.n135 163.367
R338 B.n335 B.n2 163.367
R339 B.n426 B.n2 163.367
R340 B.n426 B.n3 163.367
R341 B.n422 B.n3 163.367
R342 B.n422 B.n9 163.367
R343 B.n418 B.n9 163.367
R344 B.n418 B.n11 163.367
R345 B.n414 B.n11 163.367
R346 B.n414 B.n16 163.367
R347 B.n410 B.n16 163.367
R348 B.n410 B.n18 163.367
R349 B.n406 B.n18 163.367
R350 B.n406 B.n23 163.367
R351 B.n402 B.n23 163.367
R352 B.n402 B.n25 163.367
R353 B.n398 B.n25 163.367
R354 B.n398 B.n30 163.367
R355 B.n394 B.n30 163.367
R356 B.n394 B.n32 163.367
R357 B.n390 B.n32 163.367
R358 B.n390 B.n37 163.367
R359 B.n386 B.n37 163.367
R360 B.n386 B.n39 163.367
R361 B.n382 B.n39 163.367
R362 B.n382 B.n44 163.367
R363 B.n378 B.n44 163.367
R364 B.n378 B.n46 163.367
R365 B.n197 B.n196 163.367
R366 B.n256 B.n196 163.367
R367 B.n254 B.n253 163.367
R368 B.n250 B.n249 163.367
R369 B.n246 B.n245 163.367
R370 B.n242 B.n241 163.367
R371 B.n238 B.n237 163.367
R372 B.n234 B.n233 163.367
R373 B.n230 B.n229 163.367
R374 B.n226 B.n225 163.367
R375 B.n222 B.n221 163.367
R376 B.n218 B.n217 163.367
R377 B.n214 B.n213 163.367
R378 B.n210 B.n209 163.367
R379 B.n206 B.n205 163.367
R380 B.n264 B.n181 163.367
R381 B.n268 B.n179 163.367
R382 B.n268 B.n173 163.367
R383 B.n276 B.n173 163.367
R384 B.n276 B.n171 163.367
R385 B.n280 B.n171 163.367
R386 B.n280 B.n165 163.367
R387 B.n288 B.n165 163.367
R388 B.n288 B.n163 163.367
R389 B.n292 B.n163 163.367
R390 B.n292 B.n157 163.367
R391 B.n300 B.n157 163.367
R392 B.n300 B.n155 163.367
R393 B.n304 B.n155 163.367
R394 B.n304 B.n149 163.367
R395 B.n312 B.n149 163.367
R396 B.n312 B.n147 163.367
R397 B.n316 B.n147 163.367
R398 B.n316 B.n141 163.367
R399 B.n324 B.n141 163.367
R400 B.n324 B.n139 163.367
R401 B.n329 B.n139 163.367
R402 B.n329 B.n133 163.367
R403 B.n337 B.n133 163.367
R404 B.n338 B.n337 163.367
R405 B.n338 B.n5 163.367
R406 B.n6 B.n5 163.367
R407 B.n7 B.n6 163.367
R408 B.n343 B.n7 163.367
R409 B.n343 B.n12 163.367
R410 B.n13 B.n12 163.367
R411 B.n14 B.n13 163.367
R412 B.n348 B.n14 163.367
R413 B.n348 B.n19 163.367
R414 B.n20 B.n19 163.367
R415 B.n21 B.n20 163.367
R416 B.n353 B.n21 163.367
R417 B.n353 B.n26 163.367
R418 B.n27 B.n26 163.367
R419 B.n28 B.n27 163.367
R420 B.n358 B.n28 163.367
R421 B.n358 B.n33 163.367
R422 B.n34 B.n33 163.367
R423 B.n35 B.n34 163.367
R424 B.n363 B.n35 163.367
R425 B.n363 B.n40 163.367
R426 B.n41 B.n40 163.367
R427 B.n42 B.n41 163.367
R428 B.n368 B.n42 163.367
R429 B.n368 B.n47 163.367
R430 B.n48 B.n47 163.367
R431 B.n73 B.n72 163.367
R432 B.n77 B.n76 163.367
R433 B.n81 B.n80 163.367
R434 B.n85 B.n84 163.367
R435 B.n89 B.n88 163.367
R436 B.n94 B.n93 163.367
R437 B.n98 B.n97 163.367
R438 B.n102 B.n101 163.367
R439 B.n106 B.n105 163.367
R440 B.n110 B.n109 163.367
R441 B.n115 B.n114 163.367
R442 B.n119 B.n118 163.367
R443 B.n123 B.n122 163.367
R444 B.n127 B.n126 163.367
R445 B.n129 B.n64 163.367
R446 B.n202 B.t8 108.808
R447 B.n66 B.t5 108.808
R448 B.n199 B.t14 108.808
R449 B.n68 B.t12 108.808
R450 B.n269 B.n178 108.328
R451 B.n269 B.n174 108.328
R452 B.n275 B.n174 108.328
R453 B.n275 B.n170 108.328
R454 B.n281 B.n170 108.328
R455 B.n281 B.n166 108.328
R456 B.n287 B.n166 108.328
R457 B.n293 B.n162 108.328
R458 B.n293 B.n158 108.328
R459 B.n299 B.n158 108.328
R460 B.n299 B.n154 108.328
R461 B.n305 B.n154 108.328
R462 B.n305 B.n150 108.328
R463 B.n311 B.n150 108.328
R464 B.n311 B.n146 108.328
R465 B.n317 B.n146 108.328
R466 B.n317 B.n142 108.328
R467 B.n323 B.n142 108.328
R468 B.n330 B.n138 108.328
R469 B.n330 B.n134 108.328
R470 B.n336 B.n134 108.328
R471 B.n336 B.n4 108.328
R472 B.n425 B.n4 108.328
R473 B.n425 B.n424 108.328
R474 B.n424 B.n423 108.328
R475 B.n423 B.n8 108.328
R476 B.n417 B.n8 108.328
R477 B.n417 B.n416 108.328
R478 B.n415 B.n15 108.328
R479 B.n409 B.n15 108.328
R480 B.n409 B.n408 108.328
R481 B.n408 B.n407 108.328
R482 B.n407 B.n22 108.328
R483 B.n401 B.n22 108.328
R484 B.n401 B.n400 108.328
R485 B.n400 B.n399 108.328
R486 B.n399 B.n29 108.328
R487 B.n393 B.n29 108.328
R488 B.n393 B.n392 108.328
R489 B.n391 B.n36 108.328
R490 B.n385 B.n36 108.328
R491 B.n385 B.n384 108.328
R492 B.n384 B.n383 108.328
R493 B.n383 B.n43 108.328
R494 B.n377 B.n43 108.328
R495 B.n377 B.n376 108.328
R496 B.t1 B.n138 95.5834
R497 B.n416 B.t0 95.5834
R498 B.n262 B.n261 71.676
R499 B.n256 B.n182 71.676
R500 B.n253 B.n183 71.676
R501 B.n249 B.n184 71.676
R502 B.n245 B.n185 71.676
R503 B.n241 B.n186 71.676
R504 B.n237 B.n187 71.676
R505 B.n233 B.n188 71.676
R506 B.n229 B.n189 71.676
R507 B.n225 B.n190 71.676
R508 B.n221 B.n191 71.676
R509 B.n217 B.n192 71.676
R510 B.n213 B.n193 71.676
R511 B.n209 B.n194 71.676
R512 B.n205 B.n195 71.676
R513 B.n69 B.n49 71.676
R514 B.n73 B.n50 71.676
R515 B.n77 B.n51 71.676
R516 B.n81 B.n52 71.676
R517 B.n85 B.n53 71.676
R518 B.n89 B.n54 71.676
R519 B.n94 B.n55 71.676
R520 B.n98 B.n56 71.676
R521 B.n102 B.n57 71.676
R522 B.n106 B.n58 71.676
R523 B.n110 B.n59 71.676
R524 B.n115 B.n60 71.676
R525 B.n119 B.n61 71.676
R526 B.n123 B.n62 71.676
R527 B.n127 B.n63 71.676
R528 B.n374 B.n64 71.676
R529 B.n374 B.n373 71.676
R530 B.n129 B.n63 71.676
R531 B.n126 B.n62 71.676
R532 B.n122 B.n61 71.676
R533 B.n118 B.n60 71.676
R534 B.n114 B.n59 71.676
R535 B.n109 B.n58 71.676
R536 B.n105 B.n57 71.676
R537 B.n101 B.n56 71.676
R538 B.n97 B.n55 71.676
R539 B.n93 B.n54 71.676
R540 B.n88 B.n53 71.676
R541 B.n84 B.n52 71.676
R542 B.n80 B.n51 71.676
R543 B.n76 B.n50 71.676
R544 B.n72 B.n49 71.676
R545 B.n262 B.n197 71.676
R546 B.n254 B.n182 71.676
R547 B.n250 B.n183 71.676
R548 B.n246 B.n184 71.676
R549 B.n242 B.n185 71.676
R550 B.n238 B.n186 71.676
R551 B.n234 B.n187 71.676
R552 B.n230 B.n188 71.676
R553 B.n226 B.n189 71.676
R554 B.n222 B.n190 71.676
R555 B.n218 B.n191 71.676
R556 B.n214 B.n192 71.676
R557 B.n210 B.n193 71.676
R558 B.n206 B.n194 71.676
R559 B.n195 B.n181 71.676
R560 B.t7 B.n162 70.0946
R561 B.n392 B.t3 70.0946
R562 B.n203 B.n202 59.5399
R563 B.n200 B.n199 59.5399
R564 B.n91 B.n68 59.5399
R565 B.n112 B.n66 59.5399
R566 B.n202 B.n201 56.4369
R567 B.n199 B.n198 56.4369
R568 B.n68 B.n67 56.4369
R569 B.n66 B.n65 56.4369
R570 B.n287 B.t7 38.2337
R571 B.t3 B.n391 38.2337
R572 B.n70 B.n45 33.8737
R573 B.n372 B.n371 33.8737
R574 B.n266 B.n265 33.8737
R575 B.n260 B.n176 33.8737
R576 B B.n427 18.0485
R577 B.n323 B.t1 12.7449
R578 B.t0 B.n415 12.7449
R579 B.n71 B.n70 10.6151
R580 B.n74 B.n71 10.6151
R581 B.n75 B.n74 10.6151
R582 B.n78 B.n75 10.6151
R583 B.n79 B.n78 10.6151
R584 B.n82 B.n79 10.6151
R585 B.n83 B.n82 10.6151
R586 B.n86 B.n83 10.6151
R587 B.n87 B.n86 10.6151
R588 B.n90 B.n87 10.6151
R589 B.n95 B.n92 10.6151
R590 B.n96 B.n95 10.6151
R591 B.n99 B.n96 10.6151
R592 B.n100 B.n99 10.6151
R593 B.n103 B.n100 10.6151
R594 B.n104 B.n103 10.6151
R595 B.n107 B.n104 10.6151
R596 B.n108 B.n107 10.6151
R597 B.n111 B.n108 10.6151
R598 B.n116 B.n113 10.6151
R599 B.n117 B.n116 10.6151
R600 B.n120 B.n117 10.6151
R601 B.n121 B.n120 10.6151
R602 B.n124 B.n121 10.6151
R603 B.n125 B.n124 10.6151
R604 B.n128 B.n125 10.6151
R605 B.n130 B.n128 10.6151
R606 B.n131 B.n130 10.6151
R607 B.n372 B.n131 10.6151
R608 B.n267 B.n266 10.6151
R609 B.n267 B.n172 10.6151
R610 B.n277 B.n172 10.6151
R611 B.n278 B.n277 10.6151
R612 B.n279 B.n278 10.6151
R613 B.n279 B.n164 10.6151
R614 B.n289 B.n164 10.6151
R615 B.n290 B.n289 10.6151
R616 B.n291 B.n290 10.6151
R617 B.n291 B.n156 10.6151
R618 B.n301 B.n156 10.6151
R619 B.n302 B.n301 10.6151
R620 B.n303 B.n302 10.6151
R621 B.n303 B.n148 10.6151
R622 B.n313 B.n148 10.6151
R623 B.n314 B.n313 10.6151
R624 B.n315 B.n314 10.6151
R625 B.n315 B.n140 10.6151
R626 B.n325 B.n140 10.6151
R627 B.n326 B.n325 10.6151
R628 B.n328 B.n326 10.6151
R629 B.n328 B.n327 10.6151
R630 B.n327 B.n132 10.6151
R631 B.n339 B.n132 10.6151
R632 B.n340 B.n339 10.6151
R633 B.n341 B.n340 10.6151
R634 B.n342 B.n341 10.6151
R635 B.n344 B.n342 10.6151
R636 B.n345 B.n344 10.6151
R637 B.n346 B.n345 10.6151
R638 B.n347 B.n346 10.6151
R639 B.n349 B.n347 10.6151
R640 B.n350 B.n349 10.6151
R641 B.n351 B.n350 10.6151
R642 B.n352 B.n351 10.6151
R643 B.n354 B.n352 10.6151
R644 B.n355 B.n354 10.6151
R645 B.n356 B.n355 10.6151
R646 B.n357 B.n356 10.6151
R647 B.n359 B.n357 10.6151
R648 B.n360 B.n359 10.6151
R649 B.n361 B.n360 10.6151
R650 B.n362 B.n361 10.6151
R651 B.n364 B.n362 10.6151
R652 B.n365 B.n364 10.6151
R653 B.n366 B.n365 10.6151
R654 B.n367 B.n366 10.6151
R655 B.n369 B.n367 10.6151
R656 B.n370 B.n369 10.6151
R657 B.n371 B.n370 10.6151
R658 B.n260 B.n259 10.6151
R659 B.n259 B.n258 10.6151
R660 B.n258 B.n257 10.6151
R661 B.n257 B.n255 10.6151
R662 B.n255 B.n252 10.6151
R663 B.n252 B.n251 10.6151
R664 B.n251 B.n248 10.6151
R665 B.n248 B.n247 10.6151
R666 B.n247 B.n244 10.6151
R667 B.n244 B.n243 10.6151
R668 B.n240 B.n239 10.6151
R669 B.n239 B.n236 10.6151
R670 B.n236 B.n235 10.6151
R671 B.n235 B.n232 10.6151
R672 B.n232 B.n231 10.6151
R673 B.n231 B.n228 10.6151
R674 B.n228 B.n227 10.6151
R675 B.n227 B.n224 10.6151
R676 B.n224 B.n223 10.6151
R677 B.n220 B.n219 10.6151
R678 B.n219 B.n216 10.6151
R679 B.n216 B.n215 10.6151
R680 B.n215 B.n212 10.6151
R681 B.n212 B.n211 10.6151
R682 B.n211 B.n208 10.6151
R683 B.n208 B.n207 10.6151
R684 B.n207 B.n204 10.6151
R685 B.n204 B.n180 10.6151
R686 B.n265 B.n180 10.6151
R687 B.n271 B.n176 10.6151
R688 B.n272 B.n271 10.6151
R689 B.n273 B.n272 10.6151
R690 B.n273 B.n168 10.6151
R691 B.n283 B.n168 10.6151
R692 B.n284 B.n283 10.6151
R693 B.n285 B.n284 10.6151
R694 B.n285 B.n160 10.6151
R695 B.n295 B.n160 10.6151
R696 B.n296 B.n295 10.6151
R697 B.n297 B.n296 10.6151
R698 B.n297 B.n152 10.6151
R699 B.n307 B.n152 10.6151
R700 B.n308 B.n307 10.6151
R701 B.n309 B.n308 10.6151
R702 B.n309 B.n144 10.6151
R703 B.n319 B.n144 10.6151
R704 B.n320 B.n319 10.6151
R705 B.n321 B.n320 10.6151
R706 B.n321 B.n136 10.6151
R707 B.n332 B.n136 10.6151
R708 B.n333 B.n332 10.6151
R709 B.n334 B.n333 10.6151
R710 B.n334 B.n0 10.6151
R711 B.n421 B.n1 10.6151
R712 B.n421 B.n420 10.6151
R713 B.n420 B.n419 10.6151
R714 B.n419 B.n10 10.6151
R715 B.n413 B.n10 10.6151
R716 B.n413 B.n412 10.6151
R717 B.n412 B.n411 10.6151
R718 B.n411 B.n17 10.6151
R719 B.n405 B.n17 10.6151
R720 B.n405 B.n404 10.6151
R721 B.n404 B.n403 10.6151
R722 B.n403 B.n24 10.6151
R723 B.n397 B.n24 10.6151
R724 B.n397 B.n396 10.6151
R725 B.n396 B.n395 10.6151
R726 B.n395 B.n31 10.6151
R727 B.n389 B.n31 10.6151
R728 B.n389 B.n388 10.6151
R729 B.n388 B.n387 10.6151
R730 B.n387 B.n38 10.6151
R731 B.n381 B.n38 10.6151
R732 B.n381 B.n380 10.6151
R733 B.n380 B.n379 10.6151
R734 B.n379 B.n45 10.6151
R735 B.n91 B.n90 9.36635
R736 B.n113 B.n112 9.36635
R737 B.n243 B.n200 9.36635
R738 B.n220 B.n203 9.36635
R739 B.n427 B.n0 2.81026
R740 B.n427 B.n1 2.81026
R741 B.n92 B.n91 1.24928
R742 B.n112 B.n111 1.24928
R743 B.n240 B.n200 1.24928
R744 B.n223 B.n203 1.24928
R745 VN VN.t0 101.24
R746 VN VN.t1 64.7331
R747 VTAIL.n3 VTAIL.t2 111.251
R748 VTAIL.n0 VTAIL.t1 111.251
R749 VTAIL.n2 VTAIL.t0 111.251
R750 VTAIL.n1 VTAIL.t3 111.251
R751 VTAIL.n1 VTAIL.n0 18.7893
R752 VTAIL.n3 VTAIL.n2 16.2807
R753 VTAIL.n2 VTAIL.n1 1.72464
R754 VTAIL VTAIL.n0 1.15567
R755 VTAIL VTAIL.n3 0.569465
R756 VDD2.n0 VDD2.t0 158.012
R757 VDD2.n0 VDD2.t1 127.93
R758 VDD2 VDD2.n0 0.685845
R759 VP.n0 VP.t1 101.144
R760 VP.n0 VP.t0 64.3968
R761 VP VP.n0 0.336784
R762 VDD1 VDD1.t1 159.163
R763 VDD1 VDD1.t0 128.614
C0 VP VDD2 0.339117f
C1 VDD2 VN 0.598362f
C2 VP VDD1 0.780843f
C3 VN VDD1 0.154971f
C4 VDD2 VTAIL 2.37145f
C5 VTAIL VDD1 2.31856f
C6 VP VN 3.53061f
C7 VDD2 VDD1 0.670986f
C8 VP VTAIL 0.935203f
C9 VTAIL VN 0.921072f
C10 VDD2 B 2.529697f
C11 VDD1 B 4.42006f
C12 VTAIL B 2.794317f
C13 VN B 7.48603f
C14 VP B 5.435647f
C15 VDD1.t0 B 0.171391f
C16 VDD1.t1 B 0.326487f
C17 VP.t1 B 0.980283f
C18 VP.t0 B 0.549384f
C19 VP.n0 B 1.89913f
C20 VDD2.t0 B 0.334441f
C21 VDD2.t1 B 0.182809f
C22 VDD2.n0 B 1.76802f
C23 VTAIL.t1 B 0.195714f
C24 VTAIL.n0 B 1.02848f
C25 VTAIL.t3 B 0.195715f
C26 VTAIL.n1 B 1.06932f
C27 VTAIL.t0 B 0.195715f
C28 VTAIL.n2 B 0.889252f
C29 VTAIL.t2 B 0.195714f
C30 VTAIL.n3 B 0.806335f
C31 VN.t1 B 0.543915f
C32 VN.t0 B 0.973584f
.ends

