* NGSPICE file created from diff_pair_sample_0867.ext - technology: sky130A

.subckt diff_pair_sample_0867 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=0 ps=0 w=8.37 l=1.65
X1 VDD1.t5 VP.t0 VTAIL.t8 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=1.38105 ps=8.7 w=8.37 l=1.65
X2 B.t8 B.t6 B.t7 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=0 ps=0 w=8.37 l=1.65
X3 VDD2.t5 VN.t0 VTAIL.t5 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=3.2643 ps=17.52 w=8.37 l=1.65
X4 VDD1.t4 VP.t1 VTAIL.t9 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=3.2643 ps=17.52 w=8.37 l=1.65
X5 B.t5 B.t3 B.t4 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=0 ps=0 w=8.37 l=1.65
X6 VTAIL.t7 VP.t2 VDD1.t3 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=1.38105 ps=8.7 w=8.37 l=1.65
X7 VTAIL.t2 VN.t1 VDD2.t4 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=1.38105 ps=8.7 w=8.37 l=1.65
X8 VDD2.t3 VN.t2 VTAIL.t3 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=3.2643 ps=17.52 w=8.37 l=1.65
X9 B.t2 B.t0 B.t1 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=0 ps=0 w=8.37 l=1.65
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=1.38105 ps=8.7 w=8.37 l=1.65
X11 VDD1.t2 VP.t3 VTAIL.t11 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=1.38105 ps=8.7 w=8.37 l=1.65
X12 VDD2.t1 VN.t4 VTAIL.t1 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=3.2643 pd=17.52 as=1.38105 ps=8.7 w=8.37 l=1.65
X13 VTAIL.t0 VN.t5 VDD2.t0 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=1.38105 ps=8.7 w=8.37 l=1.65
X14 VDD1.t1 VP.t4 VTAIL.t10 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=3.2643 ps=17.52 w=8.37 l=1.65
X15 VTAIL.t6 VP.t5 VDD1.t0 w_n2554_n2642# sky130_fd_pr__pfet_01v8 ad=1.38105 pd=8.7 as=1.38105 ps=8.7 w=8.37 l=1.65
R0 B.n296 B.n89 585
R1 B.n295 B.n294 585
R2 B.n293 B.n90 585
R3 B.n292 B.n291 585
R4 B.n290 B.n91 585
R5 B.n289 B.n288 585
R6 B.n287 B.n92 585
R7 B.n286 B.n285 585
R8 B.n284 B.n93 585
R9 B.n283 B.n282 585
R10 B.n281 B.n94 585
R11 B.n280 B.n279 585
R12 B.n278 B.n95 585
R13 B.n277 B.n276 585
R14 B.n275 B.n96 585
R15 B.n274 B.n273 585
R16 B.n272 B.n97 585
R17 B.n271 B.n270 585
R18 B.n269 B.n98 585
R19 B.n268 B.n267 585
R20 B.n266 B.n99 585
R21 B.n265 B.n264 585
R22 B.n263 B.n100 585
R23 B.n262 B.n261 585
R24 B.n260 B.n101 585
R25 B.n259 B.n258 585
R26 B.n257 B.n102 585
R27 B.n256 B.n255 585
R28 B.n254 B.n103 585
R29 B.n253 B.n252 585
R30 B.n251 B.n104 585
R31 B.n250 B.n249 585
R32 B.n245 B.n105 585
R33 B.n244 B.n243 585
R34 B.n242 B.n106 585
R35 B.n241 B.n240 585
R36 B.n239 B.n107 585
R37 B.n238 B.n237 585
R38 B.n236 B.n108 585
R39 B.n235 B.n234 585
R40 B.n232 B.n109 585
R41 B.n231 B.n230 585
R42 B.n229 B.n112 585
R43 B.n228 B.n227 585
R44 B.n226 B.n113 585
R45 B.n225 B.n224 585
R46 B.n223 B.n114 585
R47 B.n222 B.n221 585
R48 B.n220 B.n115 585
R49 B.n219 B.n218 585
R50 B.n217 B.n116 585
R51 B.n216 B.n215 585
R52 B.n214 B.n117 585
R53 B.n213 B.n212 585
R54 B.n211 B.n118 585
R55 B.n210 B.n209 585
R56 B.n208 B.n119 585
R57 B.n207 B.n206 585
R58 B.n205 B.n120 585
R59 B.n204 B.n203 585
R60 B.n202 B.n121 585
R61 B.n201 B.n200 585
R62 B.n199 B.n122 585
R63 B.n198 B.n197 585
R64 B.n196 B.n123 585
R65 B.n195 B.n194 585
R66 B.n193 B.n124 585
R67 B.n192 B.n191 585
R68 B.n190 B.n125 585
R69 B.n189 B.n188 585
R70 B.n187 B.n126 585
R71 B.n298 B.n297 585
R72 B.n299 B.n88 585
R73 B.n301 B.n300 585
R74 B.n302 B.n87 585
R75 B.n304 B.n303 585
R76 B.n305 B.n86 585
R77 B.n307 B.n306 585
R78 B.n308 B.n85 585
R79 B.n310 B.n309 585
R80 B.n311 B.n84 585
R81 B.n313 B.n312 585
R82 B.n314 B.n83 585
R83 B.n316 B.n315 585
R84 B.n317 B.n82 585
R85 B.n319 B.n318 585
R86 B.n320 B.n81 585
R87 B.n322 B.n321 585
R88 B.n323 B.n80 585
R89 B.n325 B.n324 585
R90 B.n326 B.n79 585
R91 B.n328 B.n327 585
R92 B.n329 B.n78 585
R93 B.n331 B.n330 585
R94 B.n332 B.n77 585
R95 B.n334 B.n333 585
R96 B.n335 B.n76 585
R97 B.n337 B.n336 585
R98 B.n338 B.n75 585
R99 B.n340 B.n339 585
R100 B.n341 B.n74 585
R101 B.n343 B.n342 585
R102 B.n344 B.n73 585
R103 B.n346 B.n345 585
R104 B.n347 B.n72 585
R105 B.n349 B.n348 585
R106 B.n350 B.n71 585
R107 B.n352 B.n351 585
R108 B.n353 B.n70 585
R109 B.n355 B.n354 585
R110 B.n356 B.n69 585
R111 B.n358 B.n357 585
R112 B.n359 B.n68 585
R113 B.n361 B.n360 585
R114 B.n362 B.n67 585
R115 B.n364 B.n363 585
R116 B.n365 B.n66 585
R117 B.n367 B.n366 585
R118 B.n368 B.n65 585
R119 B.n370 B.n369 585
R120 B.n371 B.n64 585
R121 B.n373 B.n372 585
R122 B.n374 B.n63 585
R123 B.n376 B.n375 585
R124 B.n377 B.n62 585
R125 B.n379 B.n378 585
R126 B.n380 B.n61 585
R127 B.n382 B.n381 585
R128 B.n383 B.n60 585
R129 B.n385 B.n384 585
R130 B.n386 B.n59 585
R131 B.n388 B.n387 585
R132 B.n389 B.n58 585
R133 B.n391 B.n390 585
R134 B.n392 B.n57 585
R135 B.n501 B.n500 585
R136 B.n499 B.n18 585
R137 B.n498 B.n497 585
R138 B.n496 B.n19 585
R139 B.n495 B.n494 585
R140 B.n493 B.n20 585
R141 B.n492 B.n491 585
R142 B.n490 B.n21 585
R143 B.n489 B.n488 585
R144 B.n487 B.n22 585
R145 B.n486 B.n485 585
R146 B.n484 B.n23 585
R147 B.n483 B.n482 585
R148 B.n481 B.n24 585
R149 B.n480 B.n479 585
R150 B.n478 B.n25 585
R151 B.n477 B.n476 585
R152 B.n475 B.n26 585
R153 B.n474 B.n473 585
R154 B.n472 B.n27 585
R155 B.n471 B.n470 585
R156 B.n469 B.n28 585
R157 B.n468 B.n467 585
R158 B.n466 B.n29 585
R159 B.n465 B.n464 585
R160 B.n463 B.n30 585
R161 B.n462 B.n461 585
R162 B.n460 B.n31 585
R163 B.n459 B.n458 585
R164 B.n457 B.n32 585
R165 B.n456 B.n455 585
R166 B.n453 B.n33 585
R167 B.n452 B.n451 585
R168 B.n450 B.n36 585
R169 B.n449 B.n448 585
R170 B.n447 B.n37 585
R171 B.n446 B.n445 585
R172 B.n444 B.n38 585
R173 B.n443 B.n442 585
R174 B.n441 B.n39 585
R175 B.n439 B.n438 585
R176 B.n437 B.n42 585
R177 B.n436 B.n435 585
R178 B.n434 B.n43 585
R179 B.n433 B.n432 585
R180 B.n431 B.n44 585
R181 B.n430 B.n429 585
R182 B.n428 B.n45 585
R183 B.n427 B.n426 585
R184 B.n425 B.n46 585
R185 B.n424 B.n423 585
R186 B.n422 B.n47 585
R187 B.n421 B.n420 585
R188 B.n419 B.n48 585
R189 B.n418 B.n417 585
R190 B.n416 B.n49 585
R191 B.n415 B.n414 585
R192 B.n413 B.n50 585
R193 B.n412 B.n411 585
R194 B.n410 B.n51 585
R195 B.n409 B.n408 585
R196 B.n407 B.n52 585
R197 B.n406 B.n405 585
R198 B.n404 B.n53 585
R199 B.n403 B.n402 585
R200 B.n401 B.n54 585
R201 B.n400 B.n399 585
R202 B.n398 B.n55 585
R203 B.n397 B.n396 585
R204 B.n395 B.n56 585
R205 B.n394 B.n393 585
R206 B.n502 B.n17 585
R207 B.n504 B.n503 585
R208 B.n505 B.n16 585
R209 B.n507 B.n506 585
R210 B.n508 B.n15 585
R211 B.n510 B.n509 585
R212 B.n511 B.n14 585
R213 B.n513 B.n512 585
R214 B.n514 B.n13 585
R215 B.n516 B.n515 585
R216 B.n517 B.n12 585
R217 B.n519 B.n518 585
R218 B.n520 B.n11 585
R219 B.n522 B.n521 585
R220 B.n523 B.n10 585
R221 B.n525 B.n524 585
R222 B.n526 B.n9 585
R223 B.n528 B.n527 585
R224 B.n529 B.n8 585
R225 B.n531 B.n530 585
R226 B.n532 B.n7 585
R227 B.n534 B.n533 585
R228 B.n535 B.n6 585
R229 B.n537 B.n536 585
R230 B.n538 B.n5 585
R231 B.n540 B.n539 585
R232 B.n541 B.n4 585
R233 B.n543 B.n542 585
R234 B.n544 B.n3 585
R235 B.n546 B.n545 585
R236 B.n547 B.n0 585
R237 B.n2 B.n1 585
R238 B.n142 B.n141 585
R239 B.n144 B.n143 585
R240 B.n145 B.n140 585
R241 B.n147 B.n146 585
R242 B.n148 B.n139 585
R243 B.n150 B.n149 585
R244 B.n151 B.n138 585
R245 B.n153 B.n152 585
R246 B.n154 B.n137 585
R247 B.n156 B.n155 585
R248 B.n157 B.n136 585
R249 B.n159 B.n158 585
R250 B.n160 B.n135 585
R251 B.n162 B.n161 585
R252 B.n163 B.n134 585
R253 B.n165 B.n164 585
R254 B.n166 B.n133 585
R255 B.n168 B.n167 585
R256 B.n169 B.n132 585
R257 B.n171 B.n170 585
R258 B.n172 B.n131 585
R259 B.n174 B.n173 585
R260 B.n175 B.n130 585
R261 B.n177 B.n176 585
R262 B.n178 B.n129 585
R263 B.n180 B.n179 585
R264 B.n181 B.n128 585
R265 B.n183 B.n182 585
R266 B.n184 B.n127 585
R267 B.n186 B.n185 585
R268 B.n187 B.n186 521.33
R269 B.n298 B.n89 521.33
R270 B.n394 B.n57 521.33
R271 B.n500 B.n17 521.33
R272 B.n110 B.t3 328.211
R273 B.n246 B.t0 328.211
R274 B.n40 B.t9 328.211
R275 B.n34 B.t6 328.211
R276 B.n549 B.n548 256.663
R277 B.n548 B.n547 235.042
R278 B.n548 B.n2 235.042
R279 B.n188 B.n187 163.367
R280 B.n188 B.n125 163.367
R281 B.n192 B.n125 163.367
R282 B.n193 B.n192 163.367
R283 B.n194 B.n193 163.367
R284 B.n194 B.n123 163.367
R285 B.n198 B.n123 163.367
R286 B.n199 B.n198 163.367
R287 B.n200 B.n199 163.367
R288 B.n200 B.n121 163.367
R289 B.n204 B.n121 163.367
R290 B.n205 B.n204 163.367
R291 B.n206 B.n205 163.367
R292 B.n206 B.n119 163.367
R293 B.n210 B.n119 163.367
R294 B.n211 B.n210 163.367
R295 B.n212 B.n211 163.367
R296 B.n212 B.n117 163.367
R297 B.n216 B.n117 163.367
R298 B.n217 B.n216 163.367
R299 B.n218 B.n217 163.367
R300 B.n218 B.n115 163.367
R301 B.n222 B.n115 163.367
R302 B.n223 B.n222 163.367
R303 B.n224 B.n223 163.367
R304 B.n224 B.n113 163.367
R305 B.n228 B.n113 163.367
R306 B.n229 B.n228 163.367
R307 B.n230 B.n229 163.367
R308 B.n230 B.n109 163.367
R309 B.n235 B.n109 163.367
R310 B.n236 B.n235 163.367
R311 B.n237 B.n236 163.367
R312 B.n237 B.n107 163.367
R313 B.n241 B.n107 163.367
R314 B.n242 B.n241 163.367
R315 B.n243 B.n242 163.367
R316 B.n243 B.n105 163.367
R317 B.n250 B.n105 163.367
R318 B.n251 B.n250 163.367
R319 B.n252 B.n251 163.367
R320 B.n252 B.n103 163.367
R321 B.n256 B.n103 163.367
R322 B.n257 B.n256 163.367
R323 B.n258 B.n257 163.367
R324 B.n258 B.n101 163.367
R325 B.n262 B.n101 163.367
R326 B.n263 B.n262 163.367
R327 B.n264 B.n263 163.367
R328 B.n264 B.n99 163.367
R329 B.n268 B.n99 163.367
R330 B.n269 B.n268 163.367
R331 B.n270 B.n269 163.367
R332 B.n270 B.n97 163.367
R333 B.n274 B.n97 163.367
R334 B.n275 B.n274 163.367
R335 B.n276 B.n275 163.367
R336 B.n276 B.n95 163.367
R337 B.n280 B.n95 163.367
R338 B.n281 B.n280 163.367
R339 B.n282 B.n281 163.367
R340 B.n282 B.n93 163.367
R341 B.n286 B.n93 163.367
R342 B.n287 B.n286 163.367
R343 B.n288 B.n287 163.367
R344 B.n288 B.n91 163.367
R345 B.n292 B.n91 163.367
R346 B.n293 B.n292 163.367
R347 B.n294 B.n293 163.367
R348 B.n294 B.n89 163.367
R349 B.n390 B.n57 163.367
R350 B.n390 B.n389 163.367
R351 B.n389 B.n388 163.367
R352 B.n388 B.n59 163.367
R353 B.n384 B.n59 163.367
R354 B.n384 B.n383 163.367
R355 B.n383 B.n382 163.367
R356 B.n382 B.n61 163.367
R357 B.n378 B.n61 163.367
R358 B.n378 B.n377 163.367
R359 B.n377 B.n376 163.367
R360 B.n376 B.n63 163.367
R361 B.n372 B.n63 163.367
R362 B.n372 B.n371 163.367
R363 B.n371 B.n370 163.367
R364 B.n370 B.n65 163.367
R365 B.n366 B.n65 163.367
R366 B.n366 B.n365 163.367
R367 B.n365 B.n364 163.367
R368 B.n364 B.n67 163.367
R369 B.n360 B.n67 163.367
R370 B.n360 B.n359 163.367
R371 B.n359 B.n358 163.367
R372 B.n358 B.n69 163.367
R373 B.n354 B.n69 163.367
R374 B.n354 B.n353 163.367
R375 B.n353 B.n352 163.367
R376 B.n352 B.n71 163.367
R377 B.n348 B.n71 163.367
R378 B.n348 B.n347 163.367
R379 B.n347 B.n346 163.367
R380 B.n346 B.n73 163.367
R381 B.n342 B.n73 163.367
R382 B.n342 B.n341 163.367
R383 B.n341 B.n340 163.367
R384 B.n340 B.n75 163.367
R385 B.n336 B.n75 163.367
R386 B.n336 B.n335 163.367
R387 B.n335 B.n334 163.367
R388 B.n334 B.n77 163.367
R389 B.n330 B.n77 163.367
R390 B.n330 B.n329 163.367
R391 B.n329 B.n328 163.367
R392 B.n328 B.n79 163.367
R393 B.n324 B.n79 163.367
R394 B.n324 B.n323 163.367
R395 B.n323 B.n322 163.367
R396 B.n322 B.n81 163.367
R397 B.n318 B.n81 163.367
R398 B.n318 B.n317 163.367
R399 B.n317 B.n316 163.367
R400 B.n316 B.n83 163.367
R401 B.n312 B.n83 163.367
R402 B.n312 B.n311 163.367
R403 B.n311 B.n310 163.367
R404 B.n310 B.n85 163.367
R405 B.n306 B.n85 163.367
R406 B.n306 B.n305 163.367
R407 B.n305 B.n304 163.367
R408 B.n304 B.n87 163.367
R409 B.n300 B.n87 163.367
R410 B.n300 B.n299 163.367
R411 B.n299 B.n298 163.367
R412 B.n500 B.n499 163.367
R413 B.n499 B.n498 163.367
R414 B.n498 B.n19 163.367
R415 B.n494 B.n19 163.367
R416 B.n494 B.n493 163.367
R417 B.n493 B.n492 163.367
R418 B.n492 B.n21 163.367
R419 B.n488 B.n21 163.367
R420 B.n488 B.n487 163.367
R421 B.n487 B.n486 163.367
R422 B.n486 B.n23 163.367
R423 B.n482 B.n23 163.367
R424 B.n482 B.n481 163.367
R425 B.n481 B.n480 163.367
R426 B.n480 B.n25 163.367
R427 B.n476 B.n25 163.367
R428 B.n476 B.n475 163.367
R429 B.n475 B.n474 163.367
R430 B.n474 B.n27 163.367
R431 B.n470 B.n27 163.367
R432 B.n470 B.n469 163.367
R433 B.n469 B.n468 163.367
R434 B.n468 B.n29 163.367
R435 B.n464 B.n29 163.367
R436 B.n464 B.n463 163.367
R437 B.n463 B.n462 163.367
R438 B.n462 B.n31 163.367
R439 B.n458 B.n31 163.367
R440 B.n458 B.n457 163.367
R441 B.n457 B.n456 163.367
R442 B.n456 B.n33 163.367
R443 B.n451 B.n33 163.367
R444 B.n451 B.n450 163.367
R445 B.n450 B.n449 163.367
R446 B.n449 B.n37 163.367
R447 B.n445 B.n37 163.367
R448 B.n445 B.n444 163.367
R449 B.n444 B.n443 163.367
R450 B.n443 B.n39 163.367
R451 B.n438 B.n39 163.367
R452 B.n438 B.n437 163.367
R453 B.n437 B.n436 163.367
R454 B.n436 B.n43 163.367
R455 B.n432 B.n43 163.367
R456 B.n432 B.n431 163.367
R457 B.n431 B.n430 163.367
R458 B.n430 B.n45 163.367
R459 B.n426 B.n45 163.367
R460 B.n426 B.n425 163.367
R461 B.n425 B.n424 163.367
R462 B.n424 B.n47 163.367
R463 B.n420 B.n47 163.367
R464 B.n420 B.n419 163.367
R465 B.n419 B.n418 163.367
R466 B.n418 B.n49 163.367
R467 B.n414 B.n49 163.367
R468 B.n414 B.n413 163.367
R469 B.n413 B.n412 163.367
R470 B.n412 B.n51 163.367
R471 B.n408 B.n51 163.367
R472 B.n408 B.n407 163.367
R473 B.n407 B.n406 163.367
R474 B.n406 B.n53 163.367
R475 B.n402 B.n53 163.367
R476 B.n402 B.n401 163.367
R477 B.n401 B.n400 163.367
R478 B.n400 B.n55 163.367
R479 B.n396 B.n55 163.367
R480 B.n396 B.n395 163.367
R481 B.n395 B.n394 163.367
R482 B.n504 B.n17 163.367
R483 B.n505 B.n504 163.367
R484 B.n506 B.n505 163.367
R485 B.n506 B.n15 163.367
R486 B.n510 B.n15 163.367
R487 B.n511 B.n510 163.367
R488 B.n512 B.n511 163.367
R489 B.n512 B.n13 163.367
R490 B.n516 B.n13 163.367
R491 B.n517 B.n516 163.367
R492 B.n518 B.n517 163.367
R493 B.n518 B.n11 163.367
R494 B.n522 B.n11 163.367
R495 B.n523 B.n522 163.367
R496 B.n524 B.n523 163.367
R497 B.n524 B.n9 163.367
R498 B.n528 B.n9 163.367
R499 B.n529 B.n528 163.367
R500 B.n530 B.n529 163.367
R501 B.n530 B.n7 163.367
R502 B.n534 B.n7 163.367
R503 B.n535 B.n534 163.367
R504 B.n536 B.n535 163.367
R505 B.n536 B.n5 163.367
R506 B.n540 B.n5 163.367
R507 B.n541 B.n540 163.367
R508 B.n542 B.n541 163.367
R509 B.n542 B.n3 163.367
R510 B.n546 B.n3 163.367
R511 B.n547 B.n546 163.367
R512 B.n141 B.n2 163.367
R513 B.n144 B.n141 163.367
R514 B.n145 B.n144 163.367
R515 B.n146 B.n145 163.367
R516 B.n146 B.n139 163.367
R517 B.n150 B.n139 163.367
R518 B.n151 B.n150 163.367
R519 B.n152 B.n151 163.367
R520 B.n152 B.n137 163.367
R521 B.n156 B.n137 163.367
R522 B.n157 B.n156 163.367
R523 B.n158 B.n157 163.367
R524 B.n158 B.n135 163.367
R525 B.n162 B.n135 163.367
R526 B.n163 B.n162 163.367
R527 B.n164 B.n163 163.367
R528 B.n164 B.n133 163.367
R529 B.n168 B.n133 163.367
R530 B.n169 B.n168 163.367
R531 B.n170 B.n169 163.367
R532 B.n170 B.n131 163.367
R533 B.n174 B.n131 163.367
R534 B.n175 B.n174 163.367
R535 B.n176 B.n175 163.367
R536 B.n176 B.n129 163.367
R537 B.n180 B.n129 163.367
R538 B.n181 B.n180 163.367
R539 B.n182 B.n181 163.367
R540 B.n182 B.n127 163.367
R541 B.n186 B.n127 163.367
R542 B.n246 B.t1 150.917
R543 B.n40 B.t11 150.917
R544 B.n110 B.t4 150.909
R545 B.n34 B.t8 150.909
R546 B.n247 B.t2 112.517
R547 B.n41 B.t10 112.517
R548 B.n111 B.t5 112.508
R549 B.n35 B.t7 112.508
R550 B.n233 B.n111 59.5399
R551 B.n248 B.n247 59.5399
R552 B.n440 B.n41 59.5399
R553 B.n454 B.n35 59.5399
R554 B.n111 B.n110 38.4005
R555 B.n247 B.n246 38.4005
R556 B.n41 B.n40 38.4005
R557 B.n35 B.n34 38.4005
R558 B.n502 B.n501 33.8737
R559 B.n393 B.n392 33.8737
R560 B.n297 B.n296 33.8737
R561 B.n185 B.n126 33.8737
R562 B B.n549 18.0485
R563 B.n503 B.n502 10.6151
R564 B.n503 B.n16 10.6151
R565 B.n507 B.n16 10.6151
R566 B.n508 B.n507 10.6151
R567 B.n509 B.n508 10.6151
R568 B.n509 B.n14 10.6151
R569 B.n513 B.n14 10.6151
R570 B.n514 B.n513 10.6151
R571 B.n515 B.n514 10.6151
R572 B.n515 B.n12 10.6151
R573 B.n519 B.n12 10.6151
R574 B.n520 B.n519 10.6151
R575 B.n521 B.n520 10.6151
R576 B.n521 B.n10 10.6151
R577 B.n525 B.n10 10.6151
R578 B.n526 B.n525 10.6151
R579 B.n527 B.n526 10.6151
R580 B.n527 B.n8 10.6151
R581 B.n531 B.n8 10.6151
R582 B.n532 B.n531 10.6151
R583 B.n533 B.n532 10.6151
R584 B.n533 B.n6 10.6151
R585 B.n537 B.n6 10.6151
R586 B.n538 B.n537 10.6151
R587 B.n539 B.n538 10.6151
R588 B.n539 B.n4 10.6151
R589 B.n543 B.n4 10.6151
R590 B.n544 B.n543 10.6151
R591 B.n545 B.n544 10.6151
R592 B.n545 B.n0 10.6151
R593 B.n501 B.n18 10.6151
R594 B.n497 B.n18 10.6151
R595 B.n497 B.n496 10.6151
R596 B.n496 B.n495 10.6151
R597 B.n495 B.n20 10.6151
R598 B.n491 B.n20 10.6151
R599 B.n491 B.n490 10.6151
R600 B.n490 B.n489 10.6151
R601 B.n489 B.n22 10.6151
R602 B.n485 B.n22 10.6151
R603 B.n485 B.n484 10.6151
R604 B.n484 B.n483 10.6151
R605 B.n483 B.n24 10.6151
R606 B.n479 B.n24 10.6151
R607 B.n479 B.n478 10.6151
R608 B.n478 B.n477 10.6151
R609 B.n477 B.n26 10.6151
R610 B.n473 B.n26 10.6151
R611 B.n473 B.n472 10.6151
R612 B.n472 B.n471 10.6151
R613 B.n471 B.n28 10.6151
R614 B.n467 B.n28 10.6151
R615 B.n467 B.n466 10.6151
R616 B.n466 B.n465 10.6151
R617 B.n465 B.n30 10.6151
R618 B.n461 B.n30 10.6151
R619 B.n461 B.n460 10.6151
R620 B.n460 B.n459 10.6151
R621 B.n459 B.n32 10.6151
R622 B.n455 B.n32 10.6151
R623 B.n453 B.n452 10.6151
R624 B.n452 B.n36 10.6151
R625 B.n448 B.n36 10.6151
R626 B.n448 B.n447 10.6151
R627 B.n447 B.n446 10.6151
R628 B.n446 B.n38 10.6151
R629 B.n442 B.n38 10.6151
R630 B.n442 B.n441 10.6151
R631 B.n439 B.n42 10.6151
R632 B.n435 B.n42 10.6151
R633 B.n435 B.n434 10.6151
R634 B.n434 B.n433 10.6151
R635 B.n433 B.n44 10.6151
R636 B.n429 B.n44 10.6151
R637 B.n429 B.n428 10.6151
R638 B.n428 B.n427 10.6151
R639 B.n427 B.n46 10.6151
R640 B.n423 B.n46 10.6151
R641 B.n423 B.n422 10.6151
R642 B.n422 B.n421 10.6151
R643 B.n421 B.n48 10.6151
R644 B.n417 B.n48 10.6151
R645 B.n417 B.n416 10.6151
R646 B.n416 B.n415 10.6151
R647 B.n415 B.n50 10.6151
R648 B.n411 B.n50 10.6151
R649 B.n411 B.n410 10.6151
R650 B.n410 B.n409 10.6151
R651 B.n409 B.n52 10.6151
R652 B.n405 B.n52 10.6151
R653 B.n405 B.n404 10.6151
R654 B.n404 B.n403 10.6151
R655 B.n403 B.n54 10.6151
R656 B.n399 B.n54 10.6151
R657 B.n399 B.n398 10.6151
R658 B.n398 B.n397 10.6151
R659 B.n397 B.n56 10.6151
R660 B.n393 B.n56 10.6151
R661 B.n392 B.n391 10.6151
R662 B.n391 B.n58 10.6151
R663 B.n387 B.n58 10.6151
R664 B.n387 B.n386 10.6151
R665 B.n386 B.n385 10.6151
R666 B.n385 B.n60 10.6151
R667 B.n381 B.n60 10.6151
R668 B.n381 B.n380 10.6151
R669 B.n380 B.n379 10.6151
R670 B.n379 B.n62 10.6151
R671 B.n375 B.n62 10.6151
R672 B.n375 B.n374 10.6151
R673 B.n374 B.n373 10.6151
R674 B.n373 B.n64 10.6151
R675 B.n369 B.n64 10.6151
R676 B.n369 B.n368 10.6151
R677 B.n368 B.n367 10.6151
R678 B.n367 B.n66 10.6151
R679 B.n363 B.n66 10.6151
R680 B.n363 B.n362 10.6151
R681 B.n362 B.n361 10.6151
R682 B.n361 B.n68 10.6151
R683 B.n357 B.n68 10.6151
R684 B.n357 B.n356 10.6151
R685 B.n356 B.n355 10.6151
R686 B.n355 B.n70 10.6151
R687 B.n351 B.n70 10.6151
R688 B.n351 B.n350 10.6151
R689 B.n350 B.n349 10.6151
R690 B.n349 B.n72 10.6151
R691 B.n345 B.n72 10.6151
R692 B.n345 B.n344 10.6151
R693 B.n344 B.n343 10.6151
R694 B.n343 B.n74 10.6151
R695 B.n339 B.n74 10.6151
R696 B.n339 B.n338 10.6151
R697 B.n338 B.n337 10.6151
R698 B.n337 B.n76 10.6151
R699 B.n333 B.n76 10.6151
R700 B.n333 B.n332 10.6151
R701 B.n332 B.n331 10.6151
R702 B.n331 B.n78 10.6151
R703 B.n327 B.n78 10.6151
R704 B.n327 B.n326 10.6151
R705 B.n326 B.n325 10.6151
R706 B.n325 B.n80 10.6151
R707 B.n321 B.n80 10.6151
R708 B.n321 B.n320 10.6151
R709 B.n320 B.n319 10.6151
R710 B.n319 B.n82 10.6151
R711 B.n315 B.n82 10.6151
R712 B.n315 B.n314 10.6151
R713 B.n314 B.n313 10.6151
R714 B.n313 B.n84 10.6151
R715 B.n309 B.n84 10.6151
R716 B.n309 B.n308 10.6151
R717 B.n308 B.n307 10.6151
R718 B.n307 B.n86 10.6151
R719 B.n303 B.n86 10.6151
R720 B.n303 B.n302 10.6151
R721 B.n302 B.n301 10.6151
R722 B.n301 B.n88 10.6151
R723 B.n297 B.n88 10.6151
R724 B.n142 B.n1 10.6151
R725 B.n143 B.n142 10.6151
R726 B.n143 B.n140 10.6151
R727 B.n147 B.n140 10.6151
R728 B.n148 B.n147 10.6151
R729 B.n149 B.n148 10.6151
R730 B.n149 B.n138 10.6151
R731 B.n153 B.n138 10.6151
R732 B.n154 B.n153 10.6151
R733 B.n155 B.n154 10.6151
R734 B.n155 B.n136 10.6151
R735 B.n159 B.n136 10.6151
R736 B.n160 B.n159 10.6151
R737 B.n161 B.n160 10.6151
R738 B.n161 B.n134 10.6151
R739 B.n165 B.n134 10.6151
R740 B.n166 B.n165 10.6151
R741 B.n167 B.n166 10.6151
R742 B.n167 B.n132 10.6151
R743 B.n171 B.n132 10.6151
R744 B.n172 B.n171 10.6151
R745 B.n173 B.n172 10.6151
R746 B.n173 B.n130 10.6151
R747 B.n177 B.n130 10.6151
R748 B.n178 B.n177 10.6151
R749 B.n179 B.n178 10.6151
R750 B.n179 B.n128 10.6151
R751 B.n183 B.n128 10.6151
R752 B.n184 B.n183 10.6151
R753 B.n185 B.n184 10.6151
R754 B.n189 B.n126 10.6151
R755 B.n190 B.n189 10.6151
R756 B.n191 B.n190 10.6151
R757 B.n191 B.n124 10.6151
R758 B.n195 B.n124 10.6151
R759 B.n196 B.n195 10.6151
R760 B.n197 B.n196 10.6151
R761 B.n197 B.n122 10.6151
R762 B.n201 B.n122 10.6151
R763 B.n202 B.n201 10.6151
R764 B.n203 B.n202 10.6151
R765 B.n203 B.n120 10.6151
R766 B.n207 B.n120 10.6151
R767 B.n208 B.n207 10.6151
R768 B.n209 B.n208 10.6151
R769 B.n209 B.n118 10.6151
R770 B.n213 B.n118 10.6151
R771 B.n214 B.n213 10.6151
R772 B.n215 B.n214 10.6151
R773 B.n215 B.n116 10.6151
R774 B.n219 B.n116 10.6151
R775 B.n220 B.n219 10.6151
R776 B.n221 B.n220 10.6151
R777 B.n221 B.n114 10.6151
R778 B.n225 B.n114 10.6151
R779 B.n226 B.n225 10.6151
R780 B.n227 B.n226 10.6151
R781 B.n227 B.n112 10.6151
R782 B.n231 B.n112 10.6151
R783 B.n232 B.n231 10.6151
R784 B.n234 B.n108 10.6151
R785 B.n238 B.n108 10.6151
R786 B.n239 B.n238 10.6151
R787 B.n240 B.n239 10.6151
R788 B.n240 B.n106 10.6151
R789 B.n244 B.n106 10.6151
R790 B.n245 B.n244 10.6151
R791 B.n249 B.n245 10.6151
R792 B.n253 B.n104 10.6151
R793 B.n254 B.n253 10.6151
R794 B.n255 B.n254 10.6151
R795 B.n255 B.n102 10.6151
R796 B.n259 B.n102 10.6151
R797 B.n260 B.n259 10.6151
R798 B.n261 B.n260 10.6151
R799 B.n261 B.n100 10.6151
R800 B.n265 B.n100 10.6151
R801 B.n266 B.n265 10.6151
R802 B.n267 B.n266 10.6151
R803 B.n267 B.n98 10.6151
R804 B.n271 B.n98 10.6151
R805 B.n272 B.n271 10.6151
R806 B.n273 B.n272 10.6151
R807 B.n273 B.n96 10.6151
R808 B.n277 B.n96 10.6151
R809 B.n278 B.n277 10.6151
R810 B.n279 B.n278 10.6151
R811 B.n279 B.n94 10.6151
R812 B.n283 B.n94 10.6151
R813 B.n284 B.n283 10.6151
R814 B.n285 B.n284 10.6151
R815 B.n285 B.n92 10.6151
R816 B.n289 B.n92 10.6151
R817 B.n290 B.n289 10.6151
R818 B.n291 B.n290 10.6151
R819 B.n291 B.n90 10.6151
R820 B.n295 B.n90 10.6151
R821 B.n296 B.n295 10.6151
R822 B.n549 B.n0 8.11757
R823 B.n549 B.n1 8.11757
R824 B.n454 B.n453 6.5566
R825 B.n441 B.n440 6.5566
R826 B.n234 B.n233 6.5566
R827 B.n249 B.n248 6.5566
R828 B.n455 B.n454 4.05904
R829 B.n440 B.n439 4.05904
R830 B.n233 B.n232 4.05904
R831 B.n248 B.n104 4.05904
R832 VP.n17 VP.n16 174.512
R833 VP.n32 VP.n31 174.512
R834 VP.n15 VP.n14 174.512
R835 VP.n9 VP.n8 161.3
R836 VP.n10 VP.n5 161.3
R837 VP.n12 VP.n11 161.3
R838 VP.n13 VP.n4 161.3
R839 VP.n30 VP.n0 161.3
R840 VP.n29 VP.n28 161.3
R841 VP.n27 VP.n1 161.3
R842 VP.n26 VP.n25 161.3
R843 VP.n23 VP.n2 161.3
R844 VP.n22 VP.n21 161.3
R845 VP.n20 VP.n3 161.3
R846 VP.n19 VP.n18 161.3
R847 VP.n6 VP.t3 156.63
R848 VP.n17 VP.t0 122.254
R849 VP.n24 VP.t2 122.254
R850 VP.n31 VP.t1 122.254
R851 VP.n14 VP.t4 122.254
R852 VP.n7 VP.t5 122.254
R853 VP.n22 VP.n3 56.5193
R854 VP.n29 VP.n1 56.5193
R855 VP.n12 VP.n5 56.5193
R856 VP.n7 VP.n6 54.2622
R857 VP.n16 VP.n15 42.1823
R858 VP.n18 VP.n3 24.4675
R859 VP.n23 VP.n22 24.4675
R860 VP.n25 VP.n1 24.4675
R861 VP.n30 VP.n29 24.4675
R862 VP.n13 VP.n12 24.4675
R863 VP.n8 VP.n5 24.4675
R864 VP.n9 VP.n6 17.6611
R865 VP.n24 VP.n23 12.234
R866 VP.n25 VP.n24 12.234
R867 VP.n8 VP.n7 12.234
R868 VP.n18 VP.n17 11.2553
R869 VP.n31 VP.n30 11.2553
R870 VP.n14 VP.n13 11.2553
R871 VP.n10 VP.n9 0.189894
R872 VP.n11 VP.n10 0.189894
R873 VP.n11 VP.n4 0.189894
R874 VP.n15 VP.n4 0.189894
R875 VP.n19 VP.n16 0.189894
R876 VP.n20 VP.n19 0.189894
R877 VP.n21 VP.n20 0.189894
R878 VP.n21 VP.n2 0.189894
R879 VP.n26 VP.n2 0.189894
R880 VP.n27 VP.n26 0.189894
R881 VP.n28 VP.n27 0.189894
R882 VP.n28 VP.n0 0.189894
R883 VP.n32 VP.n0 0.189894
R884 VP VP.n32 0.0516364
R885 VTAIL.n7 VTAIL.t5 72.5622
R886 VTAIL.n11 VTAIL.t3 72.5621
R887 VTAIL.n2 VTAIL.t9 72.5621
R888 VTAIL.n10 VTAIL.t10 72.5621
R889 VTAIL.n9 VTAIL.n8 68.6788
R890 VTAIL.n6 VTAIL.n5 68.6788
R891 VTAIL.n1 VTAIL.n0 68.6785
R892 VTAIL.n4 VTAIL.n3 68.6785
R893 VTAIL.n6 VTAIL.n4 22.9962
R894 VTAIL.n11 VTAIL.n10 21.2893
R895 VTAIL.n0 VTAIL.t1 3.88401
R896 VTAIL.n0 VTAIL.t0 3.88401
R897 VTAIL.n3 VTAIL.t8 3.88401
R898 VTAIL.n3 VTAIL.t7 3.88401
R899 VTAIL.n8 VTAIL.t11 3.88401
R900 VTAIL.n8 VTAIL.t6 3.88401
R901 VTAIL.n5 VTAIL.t4 3.88401
R902 VTAIL.n5 VTAIL.t2 3.88401
R903 VTAIL.n7 VTAIL.n6 1.7074
R904 VTAIL.n10 VTAIL.n9 1.7074
R905 VTAIL.n4 VTAIL.n2 1.7074
R906 VTAIL.n9 VTAIL.n7 1.32378
R907 VTAIL.n2 VTAIL.n1 1.32378
R908 VTAIL VTAIL.n11 1.22248
R909 VTAIL VTAIL.n1 0.485414
R910 VDD1 VDD1.t2 90.5794
R911 VDD1.n1 VDD1.t5 90.4657
R912 VDD1.n1 VDD1.n0 85.7287
R913 VDD1.n3 VDD1.n2 85.3574
R914 VDD1.n3 VDD1.n1 37.9147
R915 VDD1.n2 VDD1.t0 3.88401
R916 VDD1.n2 VDD1.t1 3.88401
R917 VDD1.n0 VDD1.t3 3.88401
R918 VDD1.n0 VDD1.t4 3.88401
R919 VDD1 VDD1.n3 0.369034
R920 VN.n11 VN.n10 174.512
R921 VN.n23 VN.n22 174.512
R922 VN.n21 VN.n12 161.3
R923 VN.n20 VN.n19 161.3
R924 VN.n18 VN.n13 161.3
R925 VN.n17 VN.n16 161.3
R926 VN.n9 VN.n0 161.3
R927 VN.n8 VN.n7 161.3
R928 VN.n6 VN.n1 161.3
R929 VN.n5 VN.n4 161.3
R930 VN.n2 VN.t4 156.63
R931 VN.n14 VN.t0 156.63
R932 VN.n3 VN.t5 122.254
R933 VN.n10 VN.t2 122.254
R934 VN.n15 VN.t1 122.254
R935 VN.n22 VN.t3 122.254
R936 VN.n8 VN.n1 56.5193
R937 VN.n20 VN.n13 56.5193
R938 VN.n3 VN.n2 54.2622
R939 VN.n15 VN.n14 54.2622
R940 VN VN.n23 42.563
R941 VN.n4 VN.n1 24.4675
R942 VN.n9 VN.n8 24.4675
R943 VN.n16 VN.n13 24.4675
R944 VN.n21 VN.n20 24.4675
R945 VN.n17 VN.n14 17.6611
R946 VN.n5 VN.n2 17.6611
R947 VN.n4 VN.n3 12.234
R948 VN.n16 VN.n15 12.234
R949 VN.n10 VN.n9 11.2553
R950 VN.n22 VN.n21 11.2553
R951 VN.n23 VN.n12 0.189894
R952 VN.n19 VN.n12 0.189894
R953 VN.n19 VN.n18 0.189894
R954 VN.n18 VN.n17 0.189894
R955 VN.n6 VN.n5 0.189894
R956 VN.n7 VN.n6 0.189894
R957 VN.n7 VN.n0 0.189894
R958 VN.n11 VN.n0 0.189894
R959 VN VN.n11 0.0516364
R960 VDD2.n1 VDD2.t1 90.4657
R961 VDD2.n2 VDD2.t2 89.241
R962 VDD2.n1 VDD2.n0 85.7287
R963 VDD2 VDD2.n3 85.7259
R964 VDD2.n2 VDD2.n1 36.4782
R965 VDD2.n3 VDD2.t4 3.88401
R966 VDD2.n3 VDD2.t5 3.88401
R967 VDD2.n0 VDD2.t0 3.88401
R968 VDD2.n0 VDD2.t3 3.88401
R969 VDD2 VDD2.n2 1.33886
C0 w_n2554_n2642# VN 4.52914f
C1 B VDD1 1.55844f
C2 VDD1 VDD2 1.06366f
C3 VTAIL VN 4.40831f
C4 VP VN 5.32777f
C5 w_n2554_n2642# VTAIL 2.38898f
C6 w_n2554_n2642# VP 4.85669f
C7 VP VTAIL 4.42261f
C8 B VN 0.923601f
C9 VDD2 VN 4.32259f
C10 B w_n2554_n2642# 7.34656f
C11 VDD1 VN 0.149509f
C12 w_n2554_n2642# VDD2 1.85615f
C13 B VTAIL 2.51544f
C14 VDD2 VTAIL 6.33064f
C15 w_n2554_n2642# VDD1 1.80155f
C16 B VP 1.4657f
C17 VDD1 VTAIL 6.2863f
C18 VP VDD2 0.37755f
C19 VDD1 VP 4.54789f
C20 B VDD2 1.60982f
C21 VDD2 VSUBS 1.305878f
C22 VDD1 VSUBS 1.692135f
C23 VTAIL VSUBS 0.871897f
C24 VN VSUBS 4.80622f
C25 VP VSUBS 2.057956f
C26 B VSUBS 3.390795f
C27 w_n2554_n2642# VSUBS 83.6384f
C28 VDD2.t1 VSUBS 1.39474f
C29 VDD2.t0 VSUBS 0.143498f
C30 VDD2.t3 VSUBS 0.143498f
C31 VDD2.n0 VSUBS 1.05523f
C32 VDD2.n1 VSUBS 2.35219f
C33 VDD2.t2 VSUBS 1.38772f
C34 VDD2.n2 VSUBS 2.14237f
C35 VDD2.t4 VSUBS 0.143498f
C36 VDD2.t5 VSUBS 0.143498f
C37 VDD2.n3 VSUBS 1.05521f
C38 VN.n0 VSUBS 0.041754f
C39 VN.t2 VSUBS 1.55166f
C40 VN.n1 VSUBS 0.059789f
C41 VN.t4 VSUBS 1.71711f
C42 VN.n2 VSUBS 0.669725f
C43 VN.t5 VSUBS 1.55166f
C44 VN.n3 VSUBS 0.660172f
C45 VN.n4 VSUBS 0.058609f
C46 VN.n5 VSUBS 0.269654f
C47 VN.n6 VSUBS 0.041754f
C48 VN.n7 VSUBS 0.041754f
C49 VN.n8 VSUBS 0.062116f
C50 VN.n9 VSUBS 0.057072f
C51 VN.n10 VSUBS 0.676005f
C52 VN.n11 VSUBS 0.04046f
C53 VN.n12 VSUBS 0.041754f
C54 VN.t3 VSUBS 1.55166f
C55 VN.n13 VSUBS 0.059789f
C56 VN.t0 VSUBS 1.71711f
C57 VN.n14 VSUBS 0.669725f
C58 VN.t1 VSUBS 1.55166f
C59 VN.n15 VSUBS 0.660172f
C60 VN.n16 VSUBS 0.058609f
C61 VN.n17 VSUBS 0.269654f
C62 VN.n18 VSUBS 0.041754f
C63 VN.n19 VSUBS 0.041754f
C64 VN.n20 VSUBS 0.062116f
C65 VN.n21 VSUBS 0.057072f
C66 VN.n22 VSUBS 0.676005f
C67 VN.n23 VSUBS 1.77144f
C68 VDD1.t2 VSUBS 1.41116f
C69 VDD1.t5 VSUBS 1.41039f
C70 VDD1.t3 VSUBS 0.145109f
C71 VDD1.t4 VSUBS 0.145109f
C72 VDD1.n0 VSUBS 1.06707f
C73 VDD1.n1 VSUBS 2.46419f
C74 VDD1.t0 VSUBS 0.145109f
C75 VDD1.t1 VSUBS 0.145109f
C76 VDD1.n2 VSUBS 1.06478f
C77 VDD1.n3 VSUBS 2.1567f
C78 VTAIL.t1 VSUBS 0.197804f
C79 VTAIL.t0 VSUBS 0.197804f
C80 VTAIL.n0 VSUBS 1.32977f
C81 VTAIL.n1 VSUBS 0.762065f
C82 VTAIL.t9 VSUBS 1.77977f
C83 VTAIL.n2 VSUBS 0.969278f
C84 VTAIL.t8 VSUBS 0.197804f
C85 VTAIL.t7 VSUBS 0.197804f
C86 VTAIL.n3 VSUBS 1.32977f
C87 VTAIL.n4 VSUBS 2.18282f
C88 VTAIL.t4 VSUBS 0.197804f
C89 VTAIL.t2 VSUBS 0.197804f
C90 VTAIL.n5 VSUBS 1.32977f
C91 VTAIL.n6 VSUBS 2.18281f
C92 VTAIL.t5 VSUBS 1.77978f
C93 VTAIL.n7 VSUBS 0.969266f
C94 VTAIL.t11 VSUBS 0.197804f
C95 VTAIL.t6 VSUBS 0.197804f
C96 VTAIL.n8 VSUBS 1.32977f
C97 VTAIL.n9 VSUBS 0.879814f
C98 VTAIL.t10 VSUBS 1.77977f
C99 VTAIL.n10 VSUBS 2.10779f
C100 VTAIL.t3 VSUBS 1.77977f
C101 VTAIL.n11 VSUBS 2.06107f
C102 VP.n0 VSUBS 0.043245f
C103 VP.t1 VSUBS 1.60708f
C104 VP.n1 VSUBS 0.061925f
C105 VP.n2 VSUBS 0.043245f
C106 VP.t2 VSUBS 1.60708f
C107 VP.n3 VSUBS 0.064335f
C108 VP.n4 VSUBS 0.043245f
C109 VP.t4 VSUBS 1.60708f
C110 VP.n5 VSUBS 0.061925f
C111 VP.t3 VSUBS 1.77845f
C112 VP.n6 VSUBS 0.693647f
C113 VP.t5 VSUBS 1.60708f
C114 VP.n7 VSUBS 0.683752f
C115 VP.n8 VSUBS 0.060702f
C116 VP.n9 VSUBS 0.279286f
C117 VP.n10 VSUBS 0.043245f
C118 VP.n11 VSUBS 0.043245f
C119 VP.n12 VSUBS 0.064335f
C120 VP.n13 VSUBS 0.05911f
C121 VP.n14 VSUBS 0.700151f
C122 VP.n15 VSUBS 1.80633f
C123 VP.n16 VSUBS 1.84318f
C124 VP.t0 VSUBS 1.60708f
C125 VP.n17 VSUBS 0.700151f
C126 VP.n18 VSUBS 0.05911f
C127 VP.n19 VSUBS 0.043245f
C128 VP.n20 VSUBS 0.043245f
C129 VP.n21 VSUBS 0.043245f
C130 VP.n22 VSUBS 0.061925f
C131 VP.n23 VSUBS 0.060702f
C132 VP.n24 VSUBS 0.597703f
C133 VP.n25 VSUBS 0.060702f
C134 VP.n26 VSUBS 0.043245f
C135 VP.n27 VSUBS 0.043245f
C136 VP.n28 VSUBS 0.043245f
C137 VP.n29 VSUBS 0.064335f
C138 VP.n30 VSUBS 0.05911f
C139 VP.n31 VSUBS 0.700151f
C140 VP.n32 VSUBS 0.041905f
C141 B.n0 VSUBS 0.00641f
C142 B.n1 VSUBS 0.00641f
C143 B.n2 VSUBS 0.00948f
C144 B.n3 VSUBS 0.007265f
C145 B.n4 VSUBS 0.007265f
C146 B.n5 VSUBS 0.007265f
C147 B.n6 VSUBS 0.007265f
C148 B.n7 VSUBS 0.007265f
C149 B.n8 VSUBS 0.007265f
C150 B.n9 VSUBS 0.007265f
C151 B.n10 VSUBS 0.007265f
C152 B.n11 VSUBS 0.007265f
C153 B.n12 VSUBS 0.007265f
C154 B.n13 VSUBS 0.007265f
C155 B.n14 VSUBS 0.007265f
C156 B.n15 VSUBS 0.007265f
C157 B.n16 VSUBS 0.007265f
C158 B.n17 VSUBS 0.017242f
C159 B.n18 VSUBS 0.007265f
C160 B.n19 VSUBS 0.007265f
C161 B.n20 VSUBS 0.007265f
C162 B.n21 VSUBS 0.007265f
C163 B.n22 VSUBS 0.007265f
C164 B.n23 VSUBS 0.007265f
C165 B.n24 VSUBS 0.007265f
C166 B.n25 VSUBS 0.007265f
C167 B.n26 VSUBS 0.007265f
C168 B.n27 VSUBS 0.007265f
C169 B.n28 VSUBS 0.007265f
C170 B.n29 VSUBS 0.007265f
C171 B.n30 VSUBS 0.007265f
C172 B.n31 VSUBS 0.007265f
C173 B.n32 VSUBS 0.007265f
C174 B.n33 VSUBS 0.007265f
C175 B.t7 VSUBS 0.269989f
C176 B.t8 VSUBS 0.285186f
C177 B.t6 VSUBS 0.647102f
C178 B.n34 VSUBS 0.139848f
C179 B.n35 VSUBS 0.070083f
C180 B.n36 VSUBS 0.007265f
C181 B.n37 VSUBS 0.007265f
C182 B.n38 VSUBS 0.007265f
C183 B.n39 VSUBS 0.007265f
C184 B.t10 VSUBS 0.269987f
C185 B.t11 VSUBS 0.285183f
C186 B.t9 VSUBS 0.647102f
C187 B.n40 VSUBS 0.13985f
C188 B.n41 VSUBS 0.070086f
C189 B.n42 VSUBS 0.007265f
C190 B.n43 VSUBS 0.007265f
C191 B.n44 VSUBS 0.007265f
C192 B.n45 VSUBS 0.007265f
C193 B.n46 VSUBS 0.007265f
C194 B.n47 VSUBS 0.007265f
C195 B.n48 VSUBS 0.007265f
C196 B.n49 VSUBS 0.007265f
C197 B.n50 VSUBS 0.007265f
C198 B.n51 VSUBS 0.007265f
C199 B.n52 VSUBS 0.007265f
C200 B.n53 VSUBS 0.007265f
C201 B.n54 VSUBS 0.007265f
C202 B.n55 VSUBS 0.007265f
C203 B.n56 VSUBS 0.007265f
C204 B.n57 VSUBS 0.017242f
C205 B.n58 VSUBS 0.007265f
C206 B.n59 VSUBS 0.007265f
C207 B.n60 VSUBS 0.007265f
C208 B.n61 VSUBS 0.007265f
C209 B.n62 VSUBS 0.007265f
C210 B.n63 VSUBS 0.007265f
C211 B.n64 VSUBS 0.007265f
C212 B.n65 VSUBS 0.007265f
C213 B.n66 VSUBS 0.007265f
C214 B.n67 VSUBS 0.007265f
C215 B.n68 VSUBS 0.007265f
C216 B.n69 VSUBS 0.007265f
C217 B.n70 VSUBS 0.007265f
C218 B.n71 VSUBS 0.007265f
C219 B.n72 VSUBS 0.007265f
C220 B.n73 VSUBS 0.007265f
C221 B.n74 VSUBS 0.007265f
C222 B.n75 VSUBS 0.007265f
C223 B.n76 VSUBS 0.007265f
C224 B.n77 VSUBS 0.007265f
C225 B.n78 VSUBS 0.007265f
C226 B.n79 VSUBS 0.007265f
C227 B.n80 VSUBS 0.007265f
C228 B.n81 VSUBS 0.007265f
C229 B.n82 VSUBS 0.007265f
C230 B.n83 VSUBS 0.007265f
C231 B.n84 VSUBS 0.007265f
C232 B.n85 VSUBS 0.007265f
C233 B.n86 VSUBS 0.007265f
C234 B.n87 VSUBS 0.007265f
C235 B.n88 VSUBS 0.007265f
C236 B.n89 VSUBS 0.017586f
C237 B.n90 VSUBS 0.007265f
C238 B.n91 VSUBS 0.007265f
C239 B.n92 VSUBS 0.007265f
C240 B.n93 VSUBS 0.007265f
C241 B.n94 VSUBS 0.007265f
C242 B.n95 VSUBS 0.007265f
C243 B.n96 VSUBS 0.007265f
C244 B.n97 VSUBS 0.007265f
C245 B.n98 VSUBS 0.007265f
C246 B.n99 VSUBS 0.007265f
C247 B.n100 VSUBS 0.007265f
C248 B.n101 VSUBS 0.007265f
C249 B.n102 VSUBS 0.007265f
C250 B.n103 VSUBS 0.007265f
C251 B.n104 VSUBS 0.005021f
C252 B.n105 VSUBS 0.007265f
C253 B.n106 VSUBS 0.007265f
C254 B.n107 VSUBS 0.007265f
C255 B.n108 VSUBS 0.007265f
C256 B.n109 VSUBS 0.007265f
C257 B.t5 VSUBS 0.269989f
C258 B.t4 VSUBS 0.285186f
C259 B.t3 VSUBS 0.647102f
C260 B.n110 VSUBS 0.139848f
C261 B.n111 VSUBS 0.070083f
C262 B.n112 VSUBS 0.007265f
C263 B.n113 VSUBS 0.007265f
C264 B.n114 VSUBS 0.007265f
C265 B.n115 VSUBS 0.007265f
C266 B.n116 VSUBS 0.007265f
C267 B.n117 VSUBS 0.007265f
C268 B.n118 VSUBS 0.007265f
C269 B.n119 VSUBS 0.007265f
C270 B.n120 VSUBS 0.007265f
C271 B.n121 VSUBS 0.007265f
C272 B.n122 VSUBS 0.007265f
C273 B.n123 VSUBS 0.007265f
C274 B.n124 VSUBS 0.007265f
C275 B.n125 VSUBS 0.007265f
C276 B.n126 VSUBS 0.017586f
C277 B.n127 VSUBS 0.007265f
C278 B.n128 VSUBS 0.007265f
C279 B.n129 VSUBS 0.007265f
C280 B.n130 VSUBS 0.007265f
C281 B.n131 VSUBS 0.007265f
C282 B.n132 VSUBS 0.007265f
C283 B.n133 VSUBS 0.007265f
C284 B.n134 VSUBS 0.007265f
C285 B.n135 VSUBS 0.007265f
C286 B.n136 VSUBS 0.007265f
C287 B.n137 VSUBS 0.007265f
C288 B.n138 VSUBS 0.007265f
C289 B.n139 VSUBS 0.007265f
C290 B.n140 VSUBS 0.007265f
C291 B.n141 VSUBS 0.007265f
C292 B.n142 VSUBS 0.007265f
C293 B.n143 VSUBS 0.007265f
C294 B.n144 VSUBS 0.007265f
C295 B.n145 VSUBS 0.007265f
C296 B.n146 VSUBS 0.007265f
C297 B.n147 VSUBS 0.007265f
C298 B.n148 VSUBS 0.007265f
C299 B.n149 VSUBS 0.007265f
C300 B.n150 VSUBS 0.007265f
C301 B.n151 VSUBS 0.007265f
C302 B.n152 VSUBS 0.007265f
C303 B.n153 VSUBS 0.007265f
C304 B.n154 VSUBS 0.007265f
C305 B.n155 VSUBS 0.007265f
C306 B.n156 VSUBS 0.007265f
C307 B.n157 VSUBS 0.007265f
C308 B.n158 VSUBS 0.007265f
C309 B.n159 VSUBS 0.007265f
C310 B.n160 VSUBS 0.007265f
C311 B.n161 VSUBS 0.007265f
C312 B.n162 VSUBS 0.007265f
C313 B.n163 VSUBS 0.007265f
C314 B.n164 VSUBS 0.007265f
C315 B.n165 VSUBS 0.007265f
C316 B.n166 VSUBS 0.007265f
C317 B.n167 VSUBS 0.007265f
C318 B.n168 VSUBS 0.007265f
C319 B.n169 VSUBS 0.007265f
C320 B.n170 VSUBS 0.007265f
C321 B.n171 VSUBS 0.007265f
C322 B.n172 VSUBS 0.007265f
C323 B.n173 VSUBS 0.007265f
C324 B.n174 VSUBS 0.007265f
C325 B.n175 VSUBS 0.007265f
C326 B.n176 VSUBS 0.007265f
C327 B.n177 VSUBS 0.007265f
C328 B.n178 VSUBS 0.007265f
C329 B.n179 VSUBS 0.007265f
C330 B.n180 VSUBS 0.007265f
C331 B.n181 VSUBS 0.007265f
C332 B.n182 VSUBS 0.007265f
C333 B.n183 VSUBS 0.007265f
C334 B.n184 VSUBS 0.007265f
C335 B.n185 VSUBS 0.017242f
C336 B.n186 VSUBS 0.017242f
C337 B.n187 VSUBS 0.017586f
C338 B.n188 VSUBS 0.007265f
C339 B.n189 VSUBS 0.007265f
C340 B.n190 VSUBS 0.007265f
C341 B.n191 VSUBS 0.007265f
C342 B.n192 VSUBS 0.007265f
C343 B.n193 VSUBS 0.007265f
C344 B.n194 VSUBS 0.007265f
C345 B.n195 VSUBS 0.007265f
C346 B.n196 VSUBS 0.007265f
C347 B.n197 VSUBS 0.007265f
C348 B.n198 VSUBS 0.007265f
C349 B.n199 VSUBS 0.007265f
C350 B.n200 VSUBS 0.007265f
C351 B.n201 VSUBS 0.007265f
C352 B.n202 VSUBS 0.007265f
C353 B.n203 VSUBS 0.007265f
C354 B.n204 VSUBS 0.007265f
C355 B.n205 VSUBS 0.007265f
C356 B.n206 VSUBS 0.007265f
C357 B.n207 VSUBS 0.007265f
C358 B.n208 VSUBS 0.007265f
C359 B.n209 VSUBS 0.007265f
C360 B.n210 VSUBS 0.007265f
C361 B.n211 VSUBS 0.007265f
C362 B.n212 VSUBS 0.007265f
C363 B.n213 VSUBS 0.007265f
C364 B.n214 VSUBS 0.007265f
C365 B.n215 VSUBS 0.007265f
C366 B.n216 VSUBS 0.007265f
C367 B.n217 VSUBS 0.007265f
C368 B.n218 VSUBS 0.007265f
C369 B.n219 VSUBS 0.007265f
C370 B.n220 VSUBS 0.007265f
C371 B.n221 VSUBS 0.007265f
C372 B.n222 VSUBS 0.007265f
C373 B.n223 VSUBS 0.007265f
C374 B.n224 VSUBS 0.007265f
C375 B.n225 VSUBS 0.007265f
C376 B.n226 VSUBS 0.007265f
C377 B.n227 VSUBS 0.007265f
C378 B.n228 VSUBS 0.007265f
C379 B.n229 VSUBS 0.007265f
C380 B.n230 VSUBS 0.007265f
C381 B.n231 VSUBS 0.007265f
C382 B.n232 VSUBS 0.005021f
C383 B.n233 VSUBS 0.016832f
C384 B.n234 VSUBS 0.005876f
C385 B.n235 VSUBS 0.007265f
C386 B.n236 VSUBS 0.007265f
C387 B.n237 VSUBS 0.007265f
C388 B.n238 VSUBS 0.007265f
C389 B.n239 VSUBS 0.007265f
C390 B.n240 VSUBS 0.007265f
C391 B.n241 VSUBS 0.007265f
C392 B.n242 VSUBS 0.007265f
C393 B.n243 VSUBS 0.007265f
C394 B.n244 VSUBS 0.007265f
C395 B.n245 VSUBS 0.007265f
C396 B.t2 VSUBS 0.269987f
C397 B.t1 VSUBS 0.285183f
C398 B.t0 VSUBS 0.647102f
C399 B.n246 VSUBS 0.13985f
C400 B.n247 VSUBS 0.070086f
C401 B.n248 VSUBS 0.016832f
C402 B.n249 VSUBS 0.005876f
C403 B.n250 VSUBS 0.007265f
C404 B.n251 VSUBS 0.007265f
C405 B.n252 VSUBS 0.007265f
C406 B.n253 VSUBS 0.007265f
C407 B.n254 VSUBS 0.007265f
C408 B.n255 VSUBS 0.007265f
C409 B.n256 VSUBS 0.007265f
C410 B.n257 VSUBS 0.007265f
C411 B.n258 VSUBS 0.007265f
C412 B.n259 VSUBS 0.007265f
C413 B.n260 VSUBS 0.007265f
C414 B.n261 VSUBS 0.007265f
C415 B.n262 VSUBS 0.007265f
C416 B.n263 VSUBS 0.007265f
C417 B.n264 VSUBS 0.007265f
C418 B.n265 VSUBS 0.007265f
C419 B.n266 VSUBS 0.007265f
C420 B.n267 VSUBS 0.007265f
C421 B.n268 VSUBS 0.007265f
C422 B.n269 VSUBS 0.007265f
C423 B.n270 VSUBS 0.007265f
C424 B.n271 VSUBS 0.007265f
C425 B.n272 VSUBS 0.007265f
C426 B.n273 VSUBS 0.007265f
C427 B.n274 VSUBS 0.007265f
C428 B.n275 VSUBS 0.007265f
C429 B.n276 VSUBS 0.007265f
C430 B.n277 VSUBS 0.007265f
C431 B.n278 VSUBS 0.007265f
C432 B.n279 VSUBS 0.007265f
C433 B.n280 VSUBS 0.007265f
C434 B.n281 VSUBS 0.007265f
C435 B.n282 VSUBS 0.007265f
C436 B.n283 VSUBS 0.007265f
C437 B.n284 VSUBS 0.007265f
C438 B.n285 VSUBS 0.007265f
C439 B.n286 VSUBS 0.007265f
C440 B.n287 VSUBS 0.007265f
C441 B.n288 VSUBS 0.007265f
C442 B.n289 VSUBS 0.007265f
C443 B.n290 VSUBS 0.007265f
C444 B.n291 VSUBS 0.007265f
C445 B.n292 VSUBS 0.007265f
C446 B.n293 VSUBS 0.007265f
C447 B.n294 VSUBS 0.007265f
C448 B.n295 VSUBS 0.007265f
C449 B.n296 VSUBS 0.016758f
C450 B.n297 VSUBS 0.01807f
C451 B.n298 VSUBS 0.017242f
C452 B.n299 VSUBS 0.007265f
C453 B.n300 VSUBS 0.007265f
C454 B.n301 VSUBS 0.007265f
C455 B.n302 VSUBS 0.007265f
C456 B.n303 VSUBS 0.007265f
C457 B.n304 VSUBS 0.007265f
C458 B.n305 VSUBS 0.007265f
C459 B.n306 VSUBS 0.007265f
C460 B.n307 VSUBS 0.007265f
C461 B.n308 VSUBS 0.007265f
C462 B.n309 VSUBS 0.007265f
C463 B.n310 VSUBS 0.007265f
C464 B.n311 VSUBS 0.007265f
C465 B.n312 VSUBS 0.007265f
C466 B.n313 VSUBS 0.007265f
C467 B.n314 VSUBS 0.007265f
C468 B.n315 VSUBS 0.007265f
C469 B.n316 VSUBS 0.007265f
C470 B.n317 VSUBS 0.007265f
C471 B.n318 VSUBS 0.007265f
C472 B.n319 VSUBS 0.007265f
C473 B.n320 VSUBS 0.007265f
C474 B.n321 VSUBS 0.007265f
C475 B.n322 VSUBS 0.007265f
C476 B.n323 VSUBS 0.007265f
C477 B.n324 VSUBS 0.007265f
C478 B.n325 VSUBS 0.007265f
C479 B.n326 VSUBS 0.007265f
C480 B.n327 VSUBS 0.007265f
C481 B.n328 VSUBS 0.007265f
C482 B.n329 VSUBS 0.007265f
C483 B.n330 VSUBS 0.007265f
C484 B.n331 VSUBS 0.007265f
C485 B.n332 VSUBS 0.007265f
C486 B.n333 VSUBS 0.007265f
C487 B.n334 VSUBS 0.007265f
C488 B.n335 VSUBS 0.007265f
C489 B.n336 VSUBS 0.007265f
C490 B.n337 VSUBS 0.007265f
C491 B.n338 VSUBS 0.007265f
C492 B.n339 VSUBS 0.007265f
C493 B.n340 VSUBS 0.007265f
C494 B.n341 VSUBS 0.007265f
C495 B.n342 VSUBS 0.007265f
C496 B.n343 VSUBS 0.007265f
C497 B.n344 VSUBS 0.007265f
C498 B.n345 VSUBS 0.007265f
C499 B.n346 VSUBS 0.007265f
C500 B.n347 VSUBS 0.007265f
C501 B.n348 VSUBS 0.007265f
C502 B.n349 VSUBS 0.007265f
C503 B.n350 VSUBS 0.007265f
C504 B.n351 VSUBS 0.007265f
C505 B.n352 VSUBS 0.007265f
C506 B.n353 VSUBS 0.007265f
C507 B.n354 VSUBS 0.007265f
C508 B.n355 VSUBS 0.007265f
C509 B.n356 VSUBS 0.007265f
C510 B.n357 VSUBS 0.007265f
C511 B.n358 VSUBS 0.007265f
C512 B.n359 VSUBS 0.007265f
C513 B.n360 VSUBS 0.007265f
C514 B.n361 VSUBS 0.007265f
C515 B.n362 VSUBS 0.007265f
C516 B.n363 VSUBS 0.007265f
C517 B.n364 VSUBS 0.007265f
C518 B.n365 VSUBS 0.007265f
C519 B.n366 VSUBS 0.007265f
C520 B.n367 VSUBS 0.007265f
C521 B.n368 VSUBS 0.007265f
C522 B.n369 VSUBS 0.007265f
C523 B.n370 VSUBS 0.007265f
C524 B.n371 VSUBS 0.007265f
C525 B.n372 VSUBS 0.007265f
C526 B.n373 VSUBS 0.007265f
C527 B.n374 VSUBS 0.007265f
C528 B.n375 VSUBS 0.007265f
C529 B.n376 VSUBS 0.007265f
C530 B.n377 VSUBS 0.007265f
C531 B.n378 VSUBS 0.007265f
C532 B.n379 VSUBS 0.007265f
C533 B.n380 VSUBS 0.007265f
C534 B.n381 VSUBS 0.007265f
C535 B.n382 VSUBS 0.007265f
C536 B.n383 VSUBS 0.007265f
C537 B.n384 VSUBS 0.007265f
C538 B.n385 VSUBS 0.007265f
C539 B.n386 VSUBS 0.007265f
C540 B.n387 VSUBS 0.007265f
C541 B.n388 VSUBS 0.007265f
C542 B.n389 VSUBS 0.007265f
C543 B.n390 VSUBS 0.007265f
C544 B.n391 VSUBS 0.007265f
C545 B.n392 VSUBS 0.017242f
C546 B.n393 VSUBS 0.017586f
C547 B.n394 VSUBS 0.017586f
C548 B.n395 VSUBS 0.007265f
C549 B.n396 VSUBS 0.007265f
C550 B.n397 VSUBS 0.007265f
C551 B.n398 VSUBS 0.007265f
C552 B.n399 VSUBS 0.007265f
C553 B.n400 VSUBS 0.007265f
C554 B.n401 VSUBS 0.007265f
C555 B.n402 VSUBS 0.007265f
C556 B.n403 VSUBS 0.007265f
C557 B.n404 VSUBS 0.007265f
C558 B.n405 VSUBS 0.007265f
C559 B.n406 VSUBS 0.007265f
C560 B.n407 VSUBS 0.007265f
C561 B.n408 VSUBS 0.007265f
C562 B.n409 VSUBS 0.007265f
C563 B.n410 VSUBS 0.007265f
C564 B.n411 VSUBS 0.007265f
C565 B.n412 VSUBS 0.007265f
C566 B.n413 VSUBS 0.007265f
C567 B.n414 VSUBS 0.007265f
C568 B.n415 VSUBS 0.007265f
C569 B.n416 VSUBS 0.007265f
C570 B.n417 VSUBS 0.007265f
C571 B.n418 VSUBS 0.007265f
C572 B.n419 VSUBS 0.007265f
C573 B.n420 VSUBS 0.007265f
C574 B.n421 VSUBS 0.007265f
C575 B.n422 VSUBS 0.007265f
C576 B.n423 VSUBS 0.007265f
C577 B.n424 VSUBS 0.007265f
C578 B.n425 VSUBS 0.007265f
C579 B.n426 VSUBS 0.007265f
C580 B.n427 VSUBS 0.007265f
C581 B.n428 VSUBS 0.007265f
C582 B.n429 VSUBS 0.007265f
C583 B.n430 VSUBS 0.007265f
C584 B.n431 VSUBS 0.007265f
C585 B.n432 VSUBS 0.007265f
C586 B.n433 VSUBS 0.007265f
C587 B.n434 VSUBS 0.007265f
C588 B.n435 VSUBS 0.007265f
C589 B.n436 VSUBS 0.007265f
C590 B.n437 VSUBS 0.007265f
C591 B.n438 VSUBS 0.007265f
C592 B.n439 VSUBS 0.005021f
C593 B.n440 VSUBS 0.016832f
C594 B.n441 VSUBS 0.005876f
C595 B.n442 VSUBS 0.007265f
C596 B.n443 VSUBS 0.007265f
C597 B.n444 VSUBS 0.007265f
C598 B.n445 VSUBS 0.007265f
C599 B.n446 VSUBS 0.007265f
C600 B.n447 VSUBS 0.007265f
C601 B.n448 VSUBS 0.007265f
C602 B.n449 VSUBS 0.007265f
C603 B.n450 VSUBS 0.007265f
C604 B.n451 VSUBS 0.007265f
C605 B.n452 VSUBS 0.007265f
C606 B.n453 VSUBS 0.005876f
C607 B.n454 VSUBS 0.016832f
C608 B.n455 VSUBS 0.005021f
C609 B.n456 VSUBS 0.007265f
C610 B.n457 VSUBS 0.007265f
C611 B.n458 VSUBS 0.007265f
C612 B.n459 VSUBS 0.007265f
C613 B.n460 VSUBS 0.007265f
C614 B.n461 VSUBS 0.007265f
C615 B.n462 VSUBS 0.007265f
C616 B.n463 VSUBS 0.007265f
C617 B.n464 VSUBS 0.007265f
C618 B.n465 VSUBS 0.007265f
C619 B.n466 VSUBS 0.007265f
C620 B.n467 VSUBS 0.007265f
C621 B.n468 VSUBS 0.007265f
C622 B.n469 VSUBS 0.007265f
C623 B.n470 VSUBS 0.007265f
C624 B.n471 VSUBS 0.007265f
C625 B.n472 VSUBS 0.007265f
C626 B.n473 VSUBS 0.007265f
C627 B.n474 VSUBS 0.007265f
C628 B.n475 VSUBS 0.007265f
C629 B.n476 VSUBS 0.007265f
C630 B.n477 VSUBS 0.007265f
C631 B.n478 VSUBS 0.007265f
C632 B.n479 VSUBS 0.007265f
C633 B.n480 VSUBS 0.007265f
C634 B.n481 VSUBS 0.007265f
C635 B.n482 VSUBS 0.007265f
C636 B.n483 VSUBS 0.007265f
C637 B.n484 VSUBS 0.007265f
C638 B.n485 VSUBS 0.007265f
C639 B.n486 VSUBS 0.007265f
C640 B.n487 VSUBS 0.007265f
C641 B.n488 VSUBS 0.007265f
C642 B.n489 VSUBS 0.007265f
C643 B.n490 VSUBS 0.007265f
C644 B.n491 VSUBS 0.007265f
C645 B.n492 VSUBS 0.007265f
C646 B.n493 VSUBS 0.007265f
C647 B.n494 VSUBS 0.007265f
C648 B.n495 VSUBS 0.007265f
C649 B.n496 VSUBS 0.007265f
C650 B.n497 VSUBS 0.007265f
C651 B.n498 VSUBS 0.007265f
C652 B.n499 VSUBS 0.007265f
C653 B.n500 VSUBS 0.017586f
C654 B.n501 VSUBS 0.017586f
C655 B.n502 VSUBS 0.017242f
C656 B.n503 VSUBS 0.007265f
C657 B.n504 VSUBS 0.007265f
C658 B.n505 VSUBS 0.007265f
C659 B.n506 VSUBS 0.007265f
C660 B.n507 VSUBS 0.007265f
C661 B.n508 VSUBS 0.007265f
C662 B.n509 VSUBS 0.007265f
C663 B.n510 VSUBS 0.007265f
C664 B.n511 VSUBS 0.007265f
C665 B.n512 VSUBS 0.007265f
C666 B.n513 VSUBS 0.007265f
C667 B.n514 VSUBS 0.007265f
C668 B.n515 VSUBS 0.007265f
C669 B.n516 VSUBS 0.007265f
C670 B.n517 VSUBS 0.007265f
C671 B.n518 VSUBS 0.007265f
C672 B.n519 VSUBS 0.007265f
C673 B.n520 VSUBS 0.007265f
C674 B.n521 VSUBS 0.007265f
C675 B.n522 VSUBS 0.007265f
C676 B.n523 VSUBS 0.007265f
C677 B.n524 VSUBS 0.007265f
C678 B.n525 VSUBS 0.007265f
C679 B.n526 VSUBS 0.007265f
C680 B.n527 VSUBS 0.007265f
C681 B.n528 VSUBS 0.007265f
C682 B.n529 VSUBS 0.007265f
C683 B.n530 VSUBS 0.007265f
C684 B.n531 VSUBS 0.007265f
C685 B.n532 VSUBS 0.007265f
C686 B.n533 VSUBS 0.007265f
C687 B.n534 VSUBS 0.007265f
C688 B.n535 VSUBS 0.007265f
C689 B.n536 VSUBS 0.007265f
C690 B.n537 VSUBS 0.007265f
C691 B.n538 VSUBS 0.007265f
C692 B.n539 VSUBS 0.007265f
C693 B.n540 VSUBS 0.007265f
C694 B.n541 VSUBS 0.007265f
C695 B.n542 VSUBS 0.007265f
C696 B.n543 VSUBS 0.007265f
C697 B.n544 VSUBS 0.007265f
C698 B.n545 VSUBS 0.007265f
C699 B.n546 VSUBS 0.007265f
C700 B.n547 VSUBS 0.00948f
C701 B.n548 VSUBS 0.010099f
C702 B.n549 VSUBS 0.020082f
.ends

