* NGSPICE file created from diff_pair_sample_0714.ext - technology: sky130A

.subckt diff_pair_sample_0714 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0.4059 ps=2.79 w=2.46 l=0.89
X1 B.t11 B.t9 B.t10 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0 ps=0 w=2.46 l=0.89
X2 VDD1.t4 VP.t1 VTAIL.t10 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.9594 ps=5.7 w=2.46 l=0.89
X3 VDD1.t3 VP.t2 VTAIL.t9 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.9594 ps=5.7 w=2.46 l=0.89
X4 VDD2.t5 VN.t0 VTAIL.t1 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.9594 ps=5.7 w=2.46 l=0.89
X5 VTAIL.t0 VN.t1 VDD2.t4 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.4059 ps=2.79 w=2.46 l=0.89
X6 VTAIL.t3 VN.t2 VDD2.t3 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.4059 ps=2.79 w=2.46 l=0.89
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.9594 ps=5.7 w=2.46 l=0.89
X8 B.t8 B.t6 B.t7 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0 ps=0 w=2.46 l=0.89
X9 VTAIL.t7 VP.t3 VDD1.t2 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.4059 ps=2.79 w=2.46 l=0.89
X10 B.t5 B.t3 B.t4 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0 ps=0 w=2.46 l=0.89
X11 VDD2.t1 VN.t4 VTAIL.t2 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0.4059 ps=2.79 w=2.46 l=0.89
X12 B.t2 B.t0 B.t1 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0 ps=0 w=2.46 l=0.89
X13 VDD1.t1 VP.t4 VTAIL.t11 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0.4059 ps=2.79 w=2.46 l=0.89
X14 VDD2.t0 VN.t5 VTAIL.t5 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.9594 pd=5.7 as=0.4059 ps=2.79 w=2.46 l=0.89
X15 VTAIL.t6 VP.t5 VDD1.t0 w_n1946_n1460# sky130_fd_pr__pfet_01v8 ad=0.4059 pd=2.79 as=0.4059 ps=2.79 w=2.46 l=0.89
R0 VP.n20 VP.n19 161.3
R1 VP.n7 VP.n6 161.3
R2 VP.n8 VP.n3 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n18 VP.n0 161.3
R5 VP.n17 VP.n16 161.3
R6 VP.n15 VP.n14 161.3
R7 VP.n13 VP.n2 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n5 VP.t4 127.615
R10 VP.n12 VP.t0 110.752
R11 VP.n19 VP.t2 110.752
R12 VP.n9 VP.t1 110.752
R13 VP.n1 VP.t3 66.614
R14 VP.n4 VP.t5 66.614
R15 VP.n14 VP.n13 54.1398
R16 VP.n18 VP.n17 54.1398
R17 VP.n8 VP.n7 54.1398
R18 VP.n6 VP.n5 43.5964
R19 VP.n5 VP.n4 42.6566
R20 VP.n11 VP.n10 34.7202
R21 VP.n14 VP.n1 12.2964
R22 VP.n17 VP.n1 12.2964
R23 VP.n7 VP.n4 12.2964
R24 VP.n13 VP.n12 3.65202
R25 VP.n19 VP.n18 3.65202
R26 VP.n9 VP.n8 3.65202
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VTAIL.n50 VTAIL.n44 756.745
R36 VTAIL.n8 VTAIL.n2 756.745
R37 VTAIL.n38 VTAIL.n32 756.745
R38 VTAIL.n24 VTAIL.n18 756.745
R39 VTAIL.n49 VTAIL.n48 585
R40 VTAIL.n51 VTAIL.n50 585
R41 VTAIL.n7 VTAIL.n6 585
R42 VTAIL.n9 VTAIL.n8 585
R43 VTAIL.n39 VTAIL.n38 585
R44 VTAIL.n37 VTAIL.n36 585
R45 VTAIL.n25 VTAIL.n24 585
R46 VTAIL.n23 VTAIL.n22 585
R47 VTAIL.n47 VTAIL.t4 355.474
R48 VTAIL.n5 VTAIL.t9 355.474
R49 VTAIL.n35 VTAIL.t10 355.474
R50 VTAIL.n21 VTAIL.t1 355.474
R51 VTAIL.n50 VTAIL.n49 171.744
R52 VTAIL.n8 VTAIL.n7 171.744
R53 VTAIL.n38 VTAIL.n37 171.744
R54 VTAIL.n24 VTAIL.n23 171.744
R55 VTAIL.n31 VTAIL.n30 136.206
R56 VTAIL.n17 VTAIL.n16 136.206
R57 VTAIL.n1 VTAIL.n0 136.206
R58 VTAIL.n15 VTAIL.n14 136.206
R59 VTAIL.n49 VTAIL.t4 85.8723
R60 VTAIL.n7 VTAIL.t9 85.8723
R61 VTAIL.n37 VTAIL.t10 85.8723
R62 VTAIL.n23 VTAIL.t1 85.8723
R63 VTAIL.n55 VTAIL.n54 33.349
R64 VTAIL.n13 VTAIL.n12 33.349
R65 VTAIL.n43 VTAIL.n42 33.349
R66 VTAIL.n29 VTAIL.n28 33.349
R67 VTAIL.n17 VTAIL.n15 16.591
R68 VTAIL.n48 VTAIL.n47 15.8418
R69 VTAIL.n6 VTAIL.n5 15.8418
R70 VTAIL.n36 VTAIL.n35 15.8418
R71 VTAIL.n22 VTAIL.n21 15.8418
R72 VTAIL.n55 VTAIL.n43 15.5393
R73 VTAIL.n0 VTAIL.t5 13.2139
R74 VTAIL.n0 VTAIL.t0 13.2139
R75 VTAIL.n14 VTAIL.t8 13.2139
R76 VTAIL.n14 VTAIL.t7 13.2139
R77 VTAIL.n30 VTAIL.t11 13.2139
R78 VTAIL.n30 VTAIL.t6 13.2139
R79 VTAIL.n16 VTAIL.t2 13.2139
R80 VTAIL.n16 VTAIL.t3 13.2139
R81 VTAIL.n51 VTAIL.n46 12.8005
R82 VTAIL.n9 VTAIL.n4 12.8005
R83 VTAIL.n39 VTAIL.n34 12.8005
R84 VTAIL.n25 VTAIL.n20 12.8005
R85 VTAIL.n52 VTAIL.n44 12.0247
R86 VTAIL.n10 VTAIL.n2 12.0247
R87 VTAIL.n40 VTAIL.n32 12.0247
R88 VTAIL.n26 VTAIL.n18 12.0247
R89 VTAIL.n54 VTAIL.n53 9.45567
R90 VTAIL.n12 VTAIL.n11 9.45567
R91 VTAIL.n42 VTAIL.n41 9.45567
R92 VTAIL.n28 VTAIL.n27 9.45567
R93 VTAIL.n53 VTAIL.n52 9.3005
R94 VTAIL.n46 VTAIL.n45 9.3005
R95 VTAIL.n11 VTAIL.n10 9.3005
R96 VTAIL.n4 VTAIL.n3 9.3005
R97 VTAIL.n41 VTAIL.n40 9.3005
R98 VTAIL.n34 VTAIL.n33 9.3005
R99 VTAIL.n27 VTAIL.n26 9.3005
R100 VTAIL.n20 VTAIL.n19 9.3005
R101 VTAIL.n35 VTAIL.n33 4.29255
R102 VTAIL.n21 VTAIL.n19 4.29255
R103 VTAIL.n47 VTAIL.n45 4.29255
R104 VTAIL.n5 VTAIL.n3 4.29255
R105 VTAIL.n54 VTAIL.n44 1.93989
R106 VTAIL.n12 VTAIL.n2 1.93989
R107 VTAIL.n42 VTAIL.n32 1.93989
R108 VTAIL.n28 VTAIL.n18 1.93989
R109 VTAIL.n52 VTAIL.n51 1.16414
R110 VTAIL.n10 VTAIL.n9 1.16414
R111 VTAIL.n40 VTAIL.n39 1.16414
R112 VTAIL.n26 VTAIL.n25 1.16414
R113 VTAIL.n29 VTAIL.n17 1.05222
R114 VTAIL.n43 VTAIL.n31 1.05222
R115 VTAIL.n15 VTAIL.n13 1.05222
R116 VTAIL.n31 VTAIL.n29 0.99619
R117 VTAIL.n13 VTAIL.n1 0.99619
R118 VTAIL VTAIL.n55 0.731103
R119 VTAIL.n48 VTAIL.n46 0.388379
R120 VTAIL.n6 VTAIL.n4 0.388379
R121 VTAIL.n36 VTAIL.n34 0.388379
R122 VTAIL.n22 VTAIL.n20 0.388379
R123 VTAIL VTAIL.n1 0.321621
R124 VTAIL.n53 VTAIL.n45 0.155672
R125 VTAIL.n11 VTAIL.n3 0.155672
R126 VTAIL.n41 VTAIL.n33 0.155672
R127 VTAIL.n27 VTAIL.n19 0.155672
R128 VDD1.n6 VDD1.n0 756.745
R129 VDD1.n17 VDD1.n11 756.745
R130 VDD1.n7 VDD1.n6 585
R131 VDD1.n5 VDD1.n4 585
R132 VDD1.n16 VDD1.n15 585
R133 VDD1.n18 VDD1.n17 585
R134 VDD1.n3 VDD1.t1 355.474
R135 VDD1.n14 VDD1.t5 355.474
R136 VDD1.n6 VDD1.n5 171.744
R137 VDD1.n17 VDD1.n16 171.744
R138 VDD1.n23 VDD1.n22 153.091
R139 VDD1.n25 VDD1.n24 152.883
R140 VDD1.n5 VDD1.t1 85.8723
R141 VDD1.n16 VDD1.t5 85.8723
R142 VDD1 VDD1.n10 50.8748
R143 VDD1.n23 VDD1.n21 50.7612
R144 VDD1.n25 VDD1.n23 30.363
R145 VDD1.n4 VDD1.n3 15.8418
R146 VDD1.n15 VDD1.n14 15.8418
R147 VDD1.n24 VDD1.t0 13.2139
R148 VDD1.n24 VDD1.t4 13.2139
R149 VDD1.n22 VDD1.t2 13.2139
R150 VDD1.n22 VDD1.t3 13.2139
R151 VDD1.n7 VDD1.n2 12.8005
R152 VDD1.n18 VDD1.n13 12.8005
R153 VDD1.n8 VDD1.n0 12.0247
R154 VDD1.n19 VDD1.n11 12.0247
R155 VDD1.n10 VDD1.n9 9.45567
R156 VDD1.n21 VDD1.n20 9.45567
R157 VDD1.n9 VDD1.n8 9.3005
R158 VDD1.n2 VDD1.n1 9.3005
R159 VDD1.n20 VDD1.n19 9.3005
R160 VDD1.n13 VDD1.n12 9.3005
R161 VDD1.n3 VDD1.n1 4.29255
R162 VDD1.n14 VDD1.n12 4.29255
R163 VDD1.n10 VDD1.n0 1.93989
R164 VDD1.n21 VDD1.n11 1.93989
R165 VDD1.n8 VDD1.n7 1.16414
R166 VDD1.n19 VDD1.n18 1.16414
R167 VDD1.n4 VDD1.n2 0.388379
R168 VDD1.n15 VDD1.n13 0.388379
R169 VDD1 VDD1.n25 0.205241
R170 VDD1.n9 VDD1.n1 0.155672
R171 VDD1.n20 VDD1.n12 0.155672
R172 B.n180 B.n59 585
R173 B.n179 B.n178 585
R174 B.n177 B.n60 585
R175 B.n176 B.n175 585
R176 B.n174 B.n61 585
R177 B.n173 B.n172 585
R178 B.n171 B.n62 585
R179 B.n170 B.n169 585
R180 B.n168 B.n63 585
R181 B.n167 B.n166 585
R182 B.n165 B.n64 585
R183 B.n164 B.n163 585
R184 B.n162 B.n65 585
R185 B.n161 B.n160 585
R186 B.n159 B.n158 585
R187 B.n157 B.n69 585
R188 B.n156 B.n155 585
R189 B.n154 B.n70 585
R190 B.n153 B.n152 585
R191 B.n151 B.n71 585
R192 B.n150 B.n149 585
R193 B.n148 B.n72 585
R194 B.n147 B.n146 585
R195 B.n144 B.n73 585
R196 B.n143 B.n142 585
R197 B.n141 B.n76 585
R198 B.n140 B.n139 585
R199 B.n138 B.n77 585
R200 B.n137 B.n136 585
R201 B.n135 B.n78 585
R202 B.n134 B.n133 585
R203 B.n132 B.n79 585
R204 B.n131 B.n130 585
R205 B.n129 B.n80 585
R206 B.n128 B.n127 585
R207 B.n126 B.n81 585
R208 B.n125 B.n124 585
R209 B.n182 B.n181 585
R210 B.n183 B.n58 585
R211 B.n185 B.n184 585
R212 B.n186 B.n57 585
R213 B.n188 B.n187 585
R214 B.n189 B.n56 585
R215 B.n191 B.n190 585
R216 B.n192 B.n55 585
R217 B.n194 B.n193 585
R218 B.n195 B.n54 585
R219 B.n197 B.n196 585
R220 B.n198 B.n53 585
R221 B.n200 B.n199 585
R222 B.n201 B.n52 585
R223 B.n203 B.n202 585
R224 B.n204 B.n51 585
R225 B.n206 B.n205 585
R226 B.n207 B.n50 585
R227 B.n209 B.n208 585
R228 B.n210 B.n49 585
R229 B.n212 B.n211 585
R230 B.n213 B.n48 585
R231 B.n215 B.n214 585
R232 B.n216 B.n47 585
R233 B.n218 B.n217 585
R234 B.n219 B.n46 585
R235 B.n221 B.n220 585
R236 B.n222 B.n45 585
R237 B.n224 B.n223 585
R238 B.n225 B.n44 585
R239 B.n227 B.n226 585
R240 B.n228 B.n43 585
R241 B.n230 B.n229 585
R242 B.n231 B.n42 585
R243 B.n233 B.n232 585
R244 B.n234 B.n41 585
R245 B.n236 B.n235 585
R246 B.n237 B.n40 585
R247 B.n239 B.n238 585
R248 B.n240 B.n39 585
R249 B.n242 B.n241 585
R250 B.n243 B.n38 585
R251 B.n245 B.n244 585
R252 B.n246 B.n37 585
R253 B.n248 B.n247 585
R254 B.n249 B.n36 585
R255 B.n306 B.n13 585
R256 B.n305 B.n304 585
R257 B.n303 B.n14 585
R258 B.n302 B.n301 585
R259 B.n300 B.n15 585
R260 B.n299 B.n298 585
R261 B.n297 B.n16 585
R262 B.n296 B.n295 585
R263 B.n294 B.n17 585
R264 B.n293 B.n292 585
R265 B.n291 B.n18 585
R266 B.n290 B.n289 585
R267 B.n288 B.n19 585
R268 B.n287 B.n286 585
R269 B.n285 B.n284 585
R270 B.n283 B.n23 585
R271 B.n282 B.n281 585
R272 B.n280 B.n24 585
R273 B.n279 B.n278 585
R274 B.n277 B.n25 585
R275 B.n276 B.n275 585
R276 B.n274 B.n26 585
R277 B.n273 B.n272 585
R278 B.n270 B.n27 585
R279 B.n269 B.n268 585
R280 B.n267 B.n30 585
R281 B.n266 B.n265 585
R282 B.n264 B.n31 585
R283 B.n263 B.n262 585
R284 B.n261 B.n32 585
R285 B.n260 B.n259 585
R286 B.n258 B.n33 585
R287 B.n257 B.n256 585
R288 B.n255 B.n34 585
R289 B.n254 B.n253 585
R290 B.n252 B.n35 585
R291 B.n251 B.n250 585
R292 B.n308 B.n307 585
R293 B.n309 B.n12 585
R294 B.n311 B.n310 585
R295 B.n312 B.n11 585
R296 B.n314 B.n313 585
R297 B.n315 B.n10 585
R298 B.n317 B.n316 585
R299 B.n318 B.n9 585
R300 B.n320 B.n319 585
R301 B.n321 B.n8 585
R302 B.n323 B.n322 585
R303 B.n324 B.n7 585
R304 B.n326 B.n325 585
R305 B.n327 B.n6 585
R306 B.n329 B.n328 585
R307 B.n330 B.n5 585
R308 B.n332 B.n331 585
R309 B.n333 B.n4 585
R310 B.n335 B.n334 585
R311 B.n336 B.n3 585
R312 B.n338 B.n337 585
R313 B.n339 B.n0 585
R314 B.n2 B.n1 585
R315 B.n93 B.n92 585
R316 B.n95 B.n94 585
R317 B.n96 B.n91 585
R318 B.n98 B.n97 585
R319 B.n99 B.n90 585
R320 B.n101 B.n100 585
R321 B.n102 B.n89 585
R322 B.n104 B.n103 585
R323 B.n105 B.n88 585
R324 B.n107 B.n106 585
R325 B.n108 B.n87 585
R326 B.n110 B.n109 585
R327 B.n111 B.n86 585
R328 B.n113 B.n112 585
R329 B.n114 B.n85 585
R330 B.n116 B.n115 585
R331 B.n117 B.n84 585
R332 B.n119 B.n118 585
R333 B.n120 B.n83 585
R334 B.n122 B.n121 585
R335 B.n123 B.n82 585
R336 B.n124 B.n123 468.476
R337 B.n182 B.n59 468.476
R338 B.n250 B.n249 468.476
R339 B.n308 B.n13 468.476
R340 B.n74 B.t0 268.731
R341 B.n66 B.t9 268.731
R342 B.n28 B.t3 268.731
R343 B.n20 B.t6 268.731
R344 B.n341 B.n340 256.663
R345 B.n66 B.t10 247.137
R346 B.n28 B.t5 247.137
R347 B.n74 B.t1 247.137
R348 B.n20 B.t8 247.137
R349 B.n340 B.n339 235.042
R350 B.n340 B.n2 235.042
R351 B.n67 B.t11 223.476
R352 B.n29 B.t4 223.476
R353 B.n75 B.t2 223.476
R354 B.n21 B.t7 223.476
R355 B.n124 B.n81 163.367
R356 B.n128 B.n81 163.367
R357 B.n129 B.n128 163.367
R358 B.n130 B.n129 163.367
R359 B.n130 B.n79 163.367
R360 B.n134 B.n79 163.367
R361 B.n135 B.n134 163.367
R362 B.n136 B.n135 163.367
R363 B.n136 B.n77 163.367
R364 B.n140 B.n77 163.367
R365 B.n141 B.n140 163.367
R366 B.n142 B.n141 163.367
R367 B.n142 B.n73 163.367
R368 B.n147 B.n73 163.367
R369 B.n148 B.n147 163.367
R370 B.n149 B.n148 163.367
R371 B.n149 B.n71 163.367
R372 B.n153 B.n71 163.367
R373 B.n154 B.n153 163.367
R374 B.n155 B.n154 163.367
R375 B.n155 B.n69 163.367
R376 B.n159 B.n69 163.367
R377 B.n160 B.n159 163.367
R378 B.n160 B.n65 163.367
R379 B.n164 B.n65 163.367
R380 B.n165 B.n164 163.367
R381 B.n166 B.n165 163.367
R382 B.n166 B.n63 163.367
R383 B.n170 B.n63 163.367
R384 B.n171 B.n170 163.367
R385 B.n172 B.n171 163.367
R386 B.n172 B.n61 163.367
R387 B.n176 B.n61 163.367
R388 B.n177 B.n176 163.367
R389 B.n178 B.n177 163.367
R390 B.n178 B.n59 163.367
R391 B.n249 B.n248 163.367
R392 B.n248 B.n37 163.367
R393 B.n244 B.n37 163.367
R394 B.n244 B.n243 163.367
R395 B.n243 B.n242 163.367
R396 B.n242 B.n39 163.367
R397 B.n238 B.n39 163.367
R398 B.n238 B.n237 163.367
R399 B.n237 B.n236 163.367
R400 B.n236 B.n41 163.367
R401 B.n232 B.n41 163.367
R402 B.n232 B.n231 163.367
R403 B.n231 B.n230 163.367
R404 B.n230 B.n43 163.367
R405 B.n226 B.n43 163.367
R406 B.n226 B.n225 163.367
R407 B.n225 B.n224 163.367
R408 B.n224 B.n45 163.367
R409 B.n220 B.n45 163.367
R410 B.n220 B.n219 163.367
R411 B.n219 B.n218 163.367
R412 B.n218 B.n47 163.367
R413 B.n214 B.n47 163.367
R414 B.n214 B.n213 163.367
R415 B.n213 B.n212 163.367
R416 B.n212 B.n49 163.367
R417 B.n208 B.n49 163.367
R418 B.n208 B.n207 163.367
R419 B.n207 B.n206 163.367
R420 B.n206 B.n51 163.367
R421 B.n202 B.n51 163.367
R422 B.n202 B.n201 163.367
R423 B.n201 B.n200 163.367
R424 B.n200 B.n53 163.367
R425 B.n196 B.n53 163.367
R426 B.n196 B.n195 163.367
R427 B.n195 B.n194 163.367
R428 B.n194 B.n55 163.367
R429 B.n190 B.n55 163.367
R430 B.n190 B.n189 163.367
R431 B.n189 B.n188 163.367
R432 B.n188 B.n57 163.367
R433 B.n184 B.n57 163.367
R434 B.n184 B.n183 163.367
R435 B.n183 B.n182 163.367
R436 B.n304 B.n13 163.367
R437 B.n304 B.n303 163.367
R438 B.n303 B.n302 163.367
R439 B.n302 B.n15 163.367
R440 B.n298 B.n15 163.367
R441 B.n298 B.n297 163.367
R442 B.n297 B.n296 163.367
R443 B.n296 B.n17 163.367
R444 B.n292 B.n17 163.367
R445 B.n292 B.n291 163.367
R446 B.n291 B.n290 163.367
R447 B.n290 B.n19 163.367
R448 B.n286 B.n19 163.367
R449 B.n286 B.n285 163.367
R450 B.n285 B.n23 163.367
R451 B.n281 B.n23 163.367
R452 B.n281 B.n280 163.367
R453 B.n280 B.n279 163.367
R454 B.n279 B.n25 163.367
R455 B.n275 B.n25 163.367
R456 B.n275 B.n274 163.367
R457 B.n274 B.n273 163.367
R458 B.n273 B.n27 163.367
R459 B.n268 B.n27 163.367
R460 B.n268 B.n267 163.367
R461 B.n267 B.n266 163.367
R462 B.n266 B.n31 163.367
R463 B.n262 B.n31 163.367
R464 B.n262 B.n261 163.367
R465 B.n261 B.n260 163.367
R466 B.n260 B.n33 163.367
R467 B.n256 B.n33 163.367
R468 B.n256 B.n255 163.367
R469 B.n255 B.n254 163.367
R470 B.n254 B.n35 163.367
R471 B.n250 B.n35 163.367
R472 B.n309 B.n308 163.367
R473 B.n310 B.n309 163.367
R474 B.n310 B.n11 163.367
R475 B.n314 B.n11 163.367
R476 B.n315 B.n314 163.367
R477 B.n316 B.n315 163.367
R478 B.n316 B.n9 163.367
R479 B.n320 B.n9 163.367
R480 B.n321 B.n320 163.367
R481 B.n322 B.n321 163.367
R482 B.n322 B.n7 163.367
R483 B.n326 B.n7 163.367
R484 B.n327 B.n326 163.367
R485 B.n328 B.n327 163.367
R486 B.n328 B.n5 163.367
R487 B.n332 B.n5 163.367
R488 B.n333 B.n332 163.367
R489 B.n334 B.n333 163.367
R490 B.n334 B.n3 163.367
R491 B.n338 B.n3 163.367
R492 B.n339 B.n338 163.367
R493 B.n93 B.n2 163.367
R494 B.n94 B.n93 163.367
R495 B.n94 B.n91 163.367
R496 B.n98 B.n91 163.367
R497 B.n99 B.n98 163.367
R498 B.n100 B.n99 163.367
R499 B.n100 B.n89 163.367
R500 B.n104 B.n89 163.367
R501 B.n105 B.n104 163.367
R502 B.n106 B.n105 163.367
R503 B.n106 B.n87 163.367
R504 B.n110 B.n87 163.367
R505 B.n111 B.n110 163.367
R506 B.n112 B.n111 163.367
R507 B.n112 B.n85 163.367
R508 B.n116 B.n85 163.367
R509 B.n117 B.n116 163.367
R510 B.n118 B.n117 163.367
R511 B.n118 B.n83 163.367
R512 B.n122 B.n83 163.367
R513 B.n123 B.n122 163.367
R514 B.n145 B.n75 59.5399
R515 B.n68 B.n67 59.5399
R516 B.n271 B.n29 59.5399
R517 B.n22 B.n21 59.5399
R518 B.n307 B.n306 30.4395
R519 B.n251 B.n36 30.4395
R520 B.n181 B.n180 30.4395
R521 B.n125 B.n82 30.4395
R522 B.n75 B.n74 23.6611
R523 B.n67 B.n66 23.6611
R524 B.n29 B.n28 23.6611
R525 B.n21 B.n20 23.6611
R526 B B.n341 18.0485
R527 B.n307 B.n12 10.6151
R528 B.n311 B.n12 10.6151
R529 B.n312 B.n311 10.6151
R530 B.n313 B.n312 10.6151
R531 B.n313 B.n10 10.6151
R532 B.n317 B.n10 10.6151
R533 B.n318 B.n317 10.6151
R534 B.n319 B.n318 10.6151
R535 B.n319 B.n8 10.6151
R536 B.n323 B.n8 10.6151
R537 B.n324 B.n323 10.6151
R538 B.n325 B.n324 10.6151
R539 B.n325 B.n6 10.6151
R540 B.n329 B.n6 10.6151
R541 B.n330 B.n329 10.6151
R542 B.n331 B.n330 10.6151
R543 B.n331 B.n4 10.6151
R544 B.n335 B.n4 10.6151
R545 B.n336 B.n335 10.6151
R546 B.n337 B.n336 10.6151
R547 B.n337 B.n0 10.6151
R548 B.n306 B.n305 10.6151
R549 B.n305 B.n14 10.6151
R550 B.n301 B.n14 10.6151
R551 B.n301 B.n300 10.6151
R552 B.n300 B.n299 10.6151
R553 B.n299 B.n16 10.6151
R554 B.n295 B.n16 10.6151
R555 B.n295 B.n294 10.6151
R556 B.n294 B.n293 10.6151
R557 B.n293 B.n18 10.6151
R558 B.n289 B.n18 10.6151
R559 B.n289 B.n288 10.6151
R560 B.n288 B.n287 10.6151
R561 B.n284 B.n283 10.6151
R562 B.n283 B.n282 10.6151
R563 B.n282 B.n24 10.6151
R564 B.n278 B.n24 10.6151
R565 B.n278 B.n277 10.6151
R566 B.n277 B.n276 10.6151
R567 B.n276 B.n26 10.6151
R568 B.n272 B.n26 10.6151
R569 B.n270 B.n269 10.6151
R570 B.n269 B.n30 10.6151
R571 B.n265 B.n30 10.6151
R572 B.n265 B.n264 10.6151
R573 B.n264 B.n263 10.6151
R574 B.n263 B.n32 10.6151
R575 B.n259 B.n32 10.6151
R576 B.n259 B.n258 10.6151
R577 B.n258 B.n257 10.6151
R578 B.n257 B.n34 10.6151
R579 B.n253 B.n34 10.6151
R580 B.n253 B.n252 10.6151
R581 B.n252 B.n251 10.6151
R582 B.n247 B.n36 10.6151
R583 B.n247 B.n246 10.6151
R584 B.n246 B.n245 10.6151
R585 B.n245 B.n38 10.6151
R586 B.n241 B.n38 10.6151
R587 B.n241 B.n240 10.6151
R588 B.n240 B.n239 10.6151
R589 B.n239 B.n40 10.6151
R590 B.n235 B.n40 10.6151
R591 B.n235 B.n234 10.6151
R592 B.n234 B.n233 10.6151
R593 B.n233 B.n42 10.6151
R594 B.n229 B.n42 10.6151
R595 B.n229 B.n228 10.6151
R596 B.n228 B.n227 10.6151
R597 B.n227 B.n44 10.6151
R598 B.n223 B.n44 10.6151
R599 B.n223 B.n222 10.6151
R600 B.n222 B.n221 10.6151
R601 B.n221 B.n46 10.6151
R602 B.n217 B.n46 10.6151
R603 B.n217 B.n216 10.6151
R604 B.n216 B.n215 10.6151
R605 B.n215 B.n48 10.6151
R606 B.n211 B.n48 10.6151
R607 B.n211 B.n210 10.6151
R608 B.n210 B.n209 10.6151
R609 B.n209 B.n50 10.6151
R610 B.n205 B.n50 10.6151
R611 B.n205 B.n204 10.6151
R612 B.n204 B.n203 10.6151
R613 B.n203 B.n52 10.6151
R614 B.n199 B.n52 10.6151
R615 B.n199 B.n198 10.6151
R616 B.n198 B.n197 10.6151
R617 B.n197 B.n54 10.6151
R618 B.n193 B.n54 10.6151
R619 B.n193 B.n192 10.6151
R620 B.n192 B.n191 10.6151
R621 B.n191 B.n56 10.6151
R622 B.n187 B.n56 10.6151
R623 B.n187 B.n186 10.6151
R624 B.n186 B.n185 10.6151
R625 B.n185 B.n58 10.6151
R626 B.n181 B.n58 10.6151
R627 B.n92 B.n1 10.6151
R628 B.n95 B.n92 10.6151
R629 B.n96 B.n95 10.6151
R630 B.n97 B.n96 10.6151
R631 B.n97 B.n90 10.6151
R632 B.n101 B.n90 10.6151
R633 B.n102 B.n101 10.6151
R634 B.n103 B.n102 10.6151
R635 B.n103 B.n88 10.6151
R636 B.n107 B.n88 10.6151
R637 B.n108 B.n107 10.6151
R638 B.n109 B.n108 10.6151
R639 B.n109 B.n86 10.6151
R640 B.n113 B.n86 10.6151
R641 B.n114 B.n113 10.6151
R642 B.n115 B.n114 10.6151
R643 B.n115 B.n84 10.6151
R644 B.n119 B.n84 10.6151
R645 B.n120 B.n119 10.6151
R646 B.n121 B.n120 10.6151
R647 B.n121 B.n82 10.6151
R648 B.n126 B.n125 10.6151
R649 B.n127 B.n126 10.6151
R650 B.n127 B.n80 10.6151
R651 B.n131 B.n80 10.6151
R652 B.n132 B.n131 10.6151
R653 B.n133 B.n132 10.6151
R654 B.n133 B.n78 10.6151
R655 B.n137 B.n78 10.6151
R656 B.n138 B.n137 10.6151
R657 B.n139 B.n138 10.6151
R658 B.n139 B.n76 10.6151
R659 B.n143 B.n76 10.6151
R660 B.n144 B.n143 10.6151
R661 B.n146 B.n72 10.6151
R662 B.n150 B.n72 10.6151
R663 B.n151 B.n150 10.6151
R664 B.n152 B.n151 10.6151
R665 B.n152 B.n70 10.6151
R666 B.n156 B.n70 10.6151
R667 B.n157 B.n156 10.6151
R668 B.n158 B.n157 10.6151
R669 B.n162 B.n161 10.6151
R670 B.n163 B.n162 10.6151
R671 B.n163 B.n64 10.6151
R672 B.n167 B.n64 10.6151
R673 B.n168 B.n167 10.6151
R674 B.n169 B.n168 10.6151
R675 B.n169 B.n62 10.6151
R676 B.n173 B.n62 10.6151
R677 B.n174 B.n173 10.6151
R678 B.n175 B.n174 10.6151
R679 B.n175 B.n60 10.6151
R680 B.n179 B.n60 10.6151
R681 B.n180 B.n179 10.6151
R682 B.n341 B.n0 8.11757
R683 B.n341 B.n1 8.11757
R684 B.n284 B.n22 6.5566
R685 B.n272 B.n271 6.5566
R686 B.n146 B.n145 6.5566
R687 B.n158 B.n68 6.5566
R688 B.n287 B.n22 4.05904
R689 B.n271 B.n270 4.05904
R690 B.n145 B.n144 4.05904
R691 B.n161 B.n68 4.05904
R692 VN.n7 VN.n6 161.3
R693 VN.n15 VN.n14 161.3
R694 VN.n13 VN.n8 161.3
R695 VN.n12 VN.n11 161.3
R696 VN.n5 VN.n0 161.3
R697 VN.n4 VN.n3 161.3
R698 VN.n2 VN.t5 127.615
R699 VN.n10 VN.t0 127.615
R700 VN.n6 VN.t3 110.752
R701 VN.n14 VN.t4 110.752
R702 VN.n1 VN.t1 66.614
R703 VN.n9 VN.t2 66.614
R704 VN.n5 VN.n4 54.1398
R705 VN.n13 VN.n12 54.1398
R706 VN.n11 VN.n10 43.5964
R707 VN.n3 VN.n2 43.5964
R708 VN.n2 VN.n1 42.6566
R709 VN.n10 VN.n9 42.6566
R710 VN VN.n15 35.1009
R711 VN.n4 VN.n1 12.2964
R712 VN.n12 VN.n9 12.2964
R713 VN.n6 VN.n5 3.65202
R714 VN.n14 VN.n13 3.65202
R715 VN.n15 VN.n8 0.189894
R716 VN.n11 VN.n8 0.189894
R717 VN.n3 VN.n0 0.189894
R718 VN.n7 VN.n0 0.189894
R719 VN VN.n7 0.0516364
R720 VDD2.n19 VDD2.n13 756.745
R721 VDD2.n6 VDD2.n0 756.745
R722 VDD2.n20 VDD2.n19 585
R723 VDD2.n18 VDD2.n17 585
R724 VDD2.n5 VDD2.n4 585
R725 VDD2.n7 VDD2.n6 585
R726 VDD2.n16 VDD2.t1 355.474
R727 VDD2.n3 VDD2.t0 355.474
R728 VDD2.n19 VDD2.n18 171.744
R729 VDD2.n6 VDD2.n5 171.744
R730 VDD2.n12 VDD2.n11 153.091
R731 VDD2 VDD2.n25 153.089
R732 VDD2.n18 VDD2.t1 85.8723
R733 VDD2.n5 VDD2.t0 85.8723
R734 VDD2.n12 VDD2.n10 50.7612
R735 VDD2.n24 VDD2.n23 50.0278
R736 VDD2.n24 VDD2.n12 29.2541
R737 VDD2.n17 VDD2.n16 15.8418
R738 VDD2.n4 VDD2.n3 15.8418
R739 VDD2.n25 VDD2.t3 13.2139
R740 VDD2.n25 VDD2.t5 13.2139
R741 VDD2.n11 VDD2.t4 13.2139
R742 VDD2.n11 VDD2.t2 13.2139
R743 VDD2.n20 VDD2.n15 12.8005
R744 VDD2.n7 VDD2.n2 12.8005
R745 VDD2.n21 VDD2.n13 12.0247
R746 VDD2.n8 VDD2.n0 12.0247
R747 VDD2.n23 VDD2.n22 9.45567
R748 VDD2.n10 VDD2.n9 9.45567
R749 VDD2.n22 VDD2.n21 9.3005
R750 VDD2.n15 VDD2.n14 9.3005
R751 VDD2.n9 VDD2.n8 9.3005
R752 VDD2.n2 VDD2.n1 9.3005
R753 VDD2.n16 VDD2.n14 4.29255
R754 VDD2.n3 VDD2.n1 4.29255
R755 VDD2.n23 VDD2.n13 1.93989
R756 VDD2.n10 VDD2.n0 1.93989
R757 VDD2.n21 VDD2.n20 1.16414
R758 VDD2.n8 VDD2.n7 1.16414
R759 VDD2 VDD2.n24 0.847483
R760 VDD2.n17 VDD2.n15 0.388379
R761 VDD2.n4 VDD2.n2 0.388379
R762 VDD2.n22 VDD2.n14 0.155672
R763 VDD2.n9 VDD2.n1 0.155672
C0 VN w_n1946_n1460# 3.06945f
C1 VN VTAIL 1.49749f
C2 VDD1 B 0.912414f
C3 VP B 1.09165f
C4 VDD1 VDD2 0.777578f
C5 VP VDD2 0.319038f
C6 VDD1 w_n1946_n1460# 1.16027f
C7 VDD1 VTAIL 3.47593f
C8 VP w_n1946_n1460# 3.31296f
C9 VP VTAIL 1.51169f
C10 VDD1 VN 0.154498f
C11 VP VN 3.50294f
C12 VDD1 VP 1.42921f
C13 B VDD2 0.94599f
C14 w_n1946_n1460# B 4.63546f
C15 VTAIL B 1.03257f
C16 w_n1946_n1460# VDD2 1.18983f
C17 VTAIL VDD2 3.51675f
C18 VTAIL w_n1946_n1460# 1.40962f
C19 VN B 0.688745f
C20 VN VDD2 1.26661f
C21 VDD2 VSUBS 0.74487f
C22 VDD1 VSUBS 0.828412f
C23 VTAIL VSUBS 0.330222f
C24 VN VSUBS 3.36136f
C25 VP VSUBS 1.144935f
C26 B VSUBS 2.028087f
C27 w_n1946_n1460# VSUBS 36.1255f
C28 VDD2.n0 VSUBS 0.017466f
C29 VDD2.n1 VSUBS 0.117043f
C30 VDD2.n2 VSUBS 0.009066f
C31 VDD2.t0 VSUBS 0.047272f
C32 VDD2.n3 VSUBS 0.05537f
C33 VDD2.n4 VSUBS 0.012635f
C34 VDD2.n5 VSUBS 0.016071f
C35 VDD2.n6 VSUBS 0.048225f
C36 VDD2.n7 VSUBS 0.009599f
C37 VDD2.n8 VSUBS 0.009066f
C38 VDD2.n9 VSUBS 0.04038f
C39 VDD2.n10 VSUBS 0.036835f
C40 VDD2.t4 VSUBS 0.032797f
C41 VDD2.t2 VSUBS 0.032797f
C42 VDD2.n11 VSUBS 0.160021f
C43 VDD2.n12 VSUBS 0.987375f
C44 VDD2.n13 VSUBS 0.017466f
C45 VDD2.n14 VSUBS 0.117043f
C46 VDD2.n15 VSUBS 0.009066f
C47 VDD2.t1 VSUBS 0.047272f
C48 VDD2.n16 VSUBS 0.05537f
C49 VDD2.n17 VSUBS 0.012635f
C50 VDD2.n18 VSUBS 0.016071f
C51 VDD2.n19 VSUBS 0.048225f
C52 VDD2.n20 VSUBS 0.009599f
C53 VDD2.n21 VSUBS 0.009066f
C54 VDD2.n22 VSUBS 0.04038f
C55 VDD2.n23 VSUBS 0.03577f
C56 VDD2.n24 VSUBS 0.897148f
C57 VDD2.t3 VSUBS 0.032797f
C58 VDD2.t5 VSUBS 0.032797f
C59 VDD2.n25 VSUBS 0.160013f
C60 VN.n0 VSUBS 0.048145f
C61 VN.t1 VSUBS 0.255378f
C62 VN.n1 VSUBS 0.186995f
C63 VN.t5 VSUBS 0.34781f
C64 VN.n2 VSUBS 0.198879f
C65 VN.n3 VSUBS 0.201389f
C66 VN.n4 VSUBS 0.061951f
C67 VN.n5 VSUBS 0.015574f
C68 VN.t3 VSUBS 0.320624f
C69 VN.n6 VSUBS 0.192004f
C70 VN.n7 VSUBS 0.037311f
C71 VN.n8 VSUBS 0.048145f
C72 VN.t2 VSUBS 0.255378f
C73 VN.n9 VSUBS 0.186995f
C74 VN.t0 VSUBS 0.34781f
C75 VN.n10 VSUBS 0.198879f
C76 VN.n11 VSUBS 0.201389f
C77 VN.n12 VSUBS 0.061951f
C78 VN.n13 VSUBS 0.015574f
C79 VN.t4 VSUBS 0.320624f
C80 VN.n14 VSUBS 0.192004f
C81 VN.n15 VSUBS 1.44444f
C82 B.n0 VSUBS 0.007333f
C83 B.n1 VSUBS 0.007333f
C84 B.n2 VSUBS 0.010844f
C85 B.n3 VSUBS 0.00831f
C86 B.n4 VSUBS 0.00831f
C87 B.n5 VSUBS 0.00831f
C88 B.n6 VSUBS 0.00831f
C89 B.n7 VSUBS 0.00831f
C90 B.n8 VSUBS 0.00831f
C91 B.n9 VSUBS 0.00831f
C92 B.n10 VSUBS 0.00831f
C93 B.n11 VSUBS 0.00831f
C94 B.n12 VSUBS 0.00831f
C95 B.n13 VSUBS 0.01918f
C96 B.n14 VSUBS 0.00831f
C97 B.n15 VSUBS 0.00831f
C98 B.n16 VSUBS 0.00831f
C99 B.n17 VSUBS 0.00831f
C100 B.n18 VSUBS 0.00831f
C101 B.n19 VSUBS 0.00831f
C102 B.t7 VSUBS 0.045198f
C103 B.t8 VSUBS 0.052336f
C104 B.t6 VSUBS 0.12271f
C105 B.n20 VSUBS 0.093718f
C106 B.n21 VSUBS 0.086407f
C107 B.n22 VSUBS 0.019254f
C108 B.n23 VSUBS 0.00831f
C109 B.n24 VSUBS 0.00831f
C110 B.n25 VSUBS 0.00831f
C111 B.n26 VSUBS 0.00831f
C112 B.n27 VSUBS 0.00831f
C113 B.t4 VSUBS 0.045198f
C114 B.t5 VSUBS 0.052336f
C115 B.t3 VSUBS 0.12271f
C116 B.n28 VSUBS 0.093718f
C117 B.n29 VSUBS 0.086407f
C118 B.n30 VSUBS 0.00831f
C119 B.n31 VSUBS 0.00831f
C120 B.n32 VSUBS 0.00831f
C121 B.n33 VSUBS 0.00831f
C122 B.n34 VSUBS 0.00831f
C123 B.n35 VSUBS 0.00831f
C124 B.n36 VSUBS 0.017972f
C125 B.n37 VSUBS 0.00831f
C126 B.n38 VSUBS 0.00831f
C127 B.n39 VSUBS 0.00831f
C128 B.n40 VSUBS 0.00831f
C129 B.n41 VSUBS 0.00831f
C130 B.n42 VSUBS 0.00831f
C131 B.n43 VSUBS 0.00831f
C132 B.n44 VSUBS 0.00831f
C133 B.n45 VSUBS 0.00831f
C134 B.n46 VSUBS 0.00831f
C135 B.n47 VSUBS 0.00831f
C136 B.n48 VSUBS 0.00831f
C137 B.n49 VSUBS 0.00831f
C138 B.n50 VSUBS 0.00831f
C139 B.n51 VSUBS 0.00831f
C140 B.n52 VSUBS 0.00831f
C141 B.n53 VSUBS 0.00831f
C142 B.n54 VSUBS 0.00831f
C143 B.n55 VSUBS 0.00831f
C144 B.n56 VSUBS 0.00831f
C145 B.n57 VSUBS 0.00831f
C146 B.n58 VSUBS 0.00831f
C147 B.n59 VSUBS 0.01918f
C148 B.n60 VSUBS 0.00831f
C149 B.n61 VSUBS 0.00831f
C150 B.n62 VSUBS 0.00831f
C151 B.n63 VSUBS 0.00831f
C152 B.n64 VSUBS 0.00831f
C153 B.n65 VSUBS 0.00831f
C154 B.t11 VSUBS 0.045198f
C155 B.t10 VSUBS 0.052336f
C156 B.t9 VSUBS 0.12271f
C157 B.n66 VSUBS 0.093718f
C158 B.n67 VSUBS 0.086407f
C159 B.n68 VSUBS 0.019254f
C160 B.n69 VSUBS 0.00831f
C161 B.n70 VSUBS 0.00831f
C162 B.n71 VSUBS 0.00831f
C163 B.n72 VSUBS 0.00831f
C164 B.n73 VSUBS 0.00831f
C165 B.t2 VSUBS 0.045198f
C166 B.t1 VSUBS 0.052336f
C167 B.t0 VSUBS 0.12271f
C168 B.n74 VSUBS 0.093718f
C169 B.n75 VSUBS 0.086407f
C170 B.n76 VSUBS 0.00831f
C171 B.n77 VSUBS 0.00831f
C172 B.n78 VSUBS 0.00831f
C173 B.n79 VSUBS 0.00831f
C174 B.n80 VSUBS 0.00831f
C175 B.n81 VSUBS 0.00831f
C176 B.n82 VSUBS 0.017972f
C177 B.n83 VSUBS 0.00831f
C178 B.n84 VSUBS 0.00831f
C179 B.n85 VSUBS 0.00831f
C180 B.n86 VSUBS 0.00831f
C181 B.n87 VSUBS 0.00831f
C182 B.n88 VSUBS 0.00831f
C183 B.n89 VSUBS 0.00831f
C184 B.n90 VSUBS 0.00831f
C185 B.n91 VSUBS 0.00831f
C186 B.n92 VSUBS 0.00831f
C187 B.n93 VSUBS 0.00831f
C188 B.n94 VSUBS 0.00831f
C189 B.n95 VSUBS 0.00831f
C190 B.n96 VSUBS 0.00831f
C191 B.n97 VSUBS 0.00831f
C192 B.n98 VSUBS 0.00831f
C193 B.n99 VSUBS 0.00831f
C194 B.n100 VSUBS 0.00831f
C195 B.n101 VSUBS 0.00831f
C196 B.n102 VSUBS 0.00831f
C197 B.n103 VSUBS 0.00831f
C198 B.n104 VSUBS 0.00831f
C199 B.n105 VSUBS 0.00831f
C200 B.n106 VSUBS 0.00831f
C201 B.n107 VSUBS 0.00831f
C202 B.n108 VSUBS 0.00831f
C203 B.n109 VSUBS 0.00831f
C204 B.n110 VSUBS 0.00831f
C205 B.n111 VSUBS 0.00831f
C206 B.n112 VSUBS 0.00831f
C207 B.n113 VSUBS 0.00831f
C208 B.n114 VSUBS 0.00831f
C209 B.n115 VSUBS 0.00831f
C210 B.n116 VSUBS 0.00831f
C211 B.n117 VSUBS 0.00831f
C212 B.n118 VSUBS 0.00831f
C213 B.n119 VSUBS 0.00831f
C214 B.n120 VSUBS 0.00831f
C215 B.n121 VSUBS 0.00831f
C216 B.n122 VSUBS 0.00831f
C217 B.n123 VSUBS 0.017972f
C218 B.n124 VSUBS 0.01918f
C219 B.n125 VSUBS 0.01918f
C220 B.n126 VSUBS 0.00831f
C221 B.n127 VSUBS 0.00831f
C222 B.n128 VSUBS 0.00831f
C223 B.n129 VSUBS 0.00831f
C224 B.n130 VSUBS 0.00831f
C225 B.n131 VSUBS 0.00831f
C226 B.n132 VSUBS 0.00831f
C227 B.n133 VSUBS 0.00831f
C228 B.n134 VSUBS 0.00831f
C229 B.n135 VSUBS 0.00831f
C230 B.n136 VSUBS 0.00831f
C231 B.n137 VSUBS 0.00831f
C232 B.n138 VSUBS 0.00831f
C233 B.n139 VSUBS 0.00831f
C234 B.n140 VSUBS 0.00831f
C235 B.n141 VSUBS 0.00831f
C236 B.n142 VSUBS 0.00831f
C237 B.n143 VSUBS 0.00831f
C238 B.n144 VSUBS 0.005744f
C239 B.n145 VSUBS 0.019254f
C240 B.n146 VSUBS 0.006721f
C241 B.n147 VSUBS 0.00831f
C242 B.n148 VSUBS 0.00831f
C243 B.n149 VSUBS 0.00831f
C244 B.n150 VSUBS 0.00831f
C245 B.n151 VSUBS 0.00831f
C246 B.n152 VSUBS 0.00831f
C247 B.n153 VSUBS 0.00831f
C248 B.n154 VSUBS 0.00831f
C249 B.n155 VSUBS 0.00831f
C250 B.n156 VSUBS 0.00831f
C251 B.n157 VSUBS 0.00831f
C252 B.n158 VSUBS 0.006721f
C253 B.n159 VSUBS 0.00831f
C254 B.n160 VSUBS 0.00831f
C255 B.n161 VSUBS 0.005744f
C256 B.n162 VSUBS 0.00831f
C257 B.n163 VSUBS 0.00831f
C258 B.n164 VSUBS 0.00831f
C259 B.n165 VSUBS 0.00831f
C260 B.n166 VSUBS 0.00831f
C261 B.n167 VSUBS 0.00831f
C262 B.n168 VSUBS 0.00831f
C263 B.n169 VSUBS 0.00831f
C264 B.n170 VSUBS 0.00831f
C265 B.n171 VSUBS 0.00831f
C266 B.n172 VSUBS 0.00831f
C267 B.n173 VSUBS 0.00831f
C268 B.n174 VSUBS 0.00831f
C269 B.n175 VSUBS 0.00831f
C270 B.n176 VSUBS 0.00831f
C271 B.n177 VSUBS 0.00831f
C272 B.n178 VSUBS 0.00831f
C273 B.n179 VSUBS 0.00831f
C274 B.n180 VSUBS 0.018126f
C275 B.n181 VSUBS 0.019025f
C276 B.n182 VSUBS 0.017972f
C277 B.n183 VSUBS 0.00831f
C278 B.n184 VSUBS 0.00831f
C279 B.n185 VSUBS 0.00831f
C280 B.n186 VSUBS 0.00831f
C281 B.n187 VSUBS 0.00831f
C282 B.n188 VSUBS 0.00831f
C283 B.n189 VSUBS 0.00831f
C284 B.n190 VSUBS 0.00831f
C285 B.n191 VSUBS 0.00831f
C286 B.n192 VSUBS 0.00831f
C287 B.n193 VSUBS 0.00831f
C288 B.n194 VSUBS 0.00831f
C289 B.n195 VSUBS 0.00831f
C290 B.n196 VSUBS 0.00831f
C291 B.n197 VSUBS 0.00831f
C292 B.n198 VSUBS 0.00831f
C293 B.n199 VSUBS 0.00831f
C294 B.n200 VSUBS 0.00831f
C295 B.n201 VSUBS 0.00831f
C296 B.n202 VSUBS 0.00831f
C297 B.n203 VSUBS 0.00831f
C298 B.n204 VSUBS 0.00831f
C299 B.n205 VSUBS 0.00831f
C300 B.n206 VSUBS 0.00831f
C301 B.n207 VSUBS 0.00831f
C302 B.n208 VSUBS 0.00831f
C303 B.n209 VSUBS 0.00831f
C304 B.n210 VSUBS 0.00831f
C305 B.n211 VSUBS 0.00831f
C306 B.n212 VSUBS 0.00831f
C307 B.n213 VSUBS 0.00831f
C308 B.n214 VSUBS 0.00831f
C309 B.n215 VSUBS 0.00831f
C310 B.n216 VSUBS 0.00831f
C311 B.n217 VSUBS 0.00831f
C312 B.n218 VSUBS 0.00831f
C313 B.n219 VSUBS 0.00831f
C314 B.n220 VSUBS 0.00831f
C315 B.n221 VSUBS 0.00831f
C316 B.n222 VSUBS 0.00831f
C317 B.n223 VSUBS 0.00831f
C318 B.n224 VSUBS 0.00831f
C319 B.n225 VSUBS 0.00831f
C320 B.n226 VSUBS 0.00831f
C321 B.n227 VSUBS 0.00831f
C322 B.n228 VSUBS 0.00831f
C323 B.n229 VSUBS 0.00831f
C324 B.n230 VSUBS 0.00831f
C325 B.n231 VSUBS 0.00831f
C326 B.n232 VSUBS 0.00831f
C327 B.n233 VSUBS 0.00831f
C328 B.n234 VSUBS 0.00831f
C329 B.n235 VSUBS 0.00831f
C330 B.n236 VSUBS 0.00831f
C331 B.n237 VSUBS 0.00831f
C332 B.n238 VSUBS 0.00831f
C333 B.n239 VSUBS 0.00831f
C334 B.n240 VSUBS 0.00831f
C335 B.n241 VSUBS 0.00831f
C336 B.n242 VSUBS 0.00831f
C337 B.n243 VSUBS 0.00831f
C338 B.n244 VSUBS 0.00831f
C339 B.n245 VSUBS 0.00831f
C340 B.n246 VSUBS 0.00831f
C341 B.n247 VSUBS 0.00831f
C342 B.n248 VSUBS 0.00831f
C343 B.n249 VSUBS 0.017972f
C344 B.n250 VSUBS 0.01918f
C345 B.n251 VSUBS 0.01918f
C346 B.n252 VSUBS 0.00831f
C347 B.n253 VSUBS 0.00831f
C348 B.n254 VSUBS 0.00831f
C349 B.n255 VSUBS 0.00831f
C350 B.n256 VSUBS 0.00831f
C351 B.n257 VSUBS 0.00831f
C352 B.n258 VSUBS 0.00831f
C353 B.n259 VSUBS 0.00831f
C354 B.n260 VSUBS 0.00831f
C355 B.n261 VSUBS 0.00831f
C356 B.n262 VSUBS 0.00831f
C357 B.n263 VSUBS 0.00831f
C358 B.n264 VSUBS 0.00831f
C359 B.n265 VSUBS 0.00831f
C360 B.n266 VSUBS 0.00831f
C361 B.n267 VSUBS 0.00831f
C362 B.n268 VSUBS 0.00831f
C363 B.n269 VSUBS 0.00831f
C364 B.n270 VSUBS 0.005744f
C365 B.n271 VSUBS 0.019254f
C366 B.n272 VSUBS 0.006721f
C367 B.n273 VSUBS 0.00831f
C368 B.n274 VSUBS 0.00831f
C369 B.n275 VSUBS 0.00831f
C370 B.n276 VSUBS 0.00831f
C371 B.n277 VSUBS 0.00831f
C372 B.n278 VSUBS 0.00831f
C373 B.n279 VSUBS 0.00831f
C374 B.n280 VSUBS 0.00831f
C375 B.n281 VSUBS 0.00831f
C376 B.n282 VSUBS 0.00831f
C377 B.n283 VSUBS 0.00831f
C378 B.n284 VSUBS 0.006721f
C379 B.n285 VSUBS 0.00831f
C380 B.n286 VSUBS 0.00831f
C381 B.n287 VSUBS 0.005744f
C382 B.n288 VSUBS 0.00831f
C383 B.n289 VSUBS 0.00831f
C384 B.n290 VSUBS 0.00831f
C385 B.n291 VSUBS 0.00831f
C386 B.n292 VSUBS 0.00831f
C387 B.n293 VSUBS 0.00831f
C388 B.n294 VSUBS 0.00831f
C389 B.n295 VSUBS 0.00831f
C390 B.n296 VSUBS 0.00831f
C391 B.n297 VSUBS 0.00831f
C392 B.n298 VSUBS 0.00831f
C393 B.n299 VSUBS 0.00831f
C394 B.n300 VSUBS 0.00831f
C395 B.n301 VSUBS 0.00831f
C396 B.n302 VSUBS 0.00831f
C397 B.n303 VSUBS 0.00831f
C398 B.n304 VSUBS 0.00831f
C399 B.n305 VSUBS 0.00831f
C400 B.n306 VSUBS 0.01918f
C401 B.n307 VSUBS 0.017972f
C402 B.n308 VSUBS 0.017972f
C403 B.n309 VSUBS 0.00831f
C404 B.n310 VSUBS 0.00831f
C405 B.n311 VSUBS 0.00831f
C406 B.n312 VSUBS 0.00831f
C407 B.n313 VSUBS 0.00831f
C408 B.n314 VSUBS 0.00831f
C409 B.n315 VSUBS 0.00831f
C410 B.n316 VSUBS 0.00831f
C411 B.n317 VSUBS 0.00831f
C412 B.n318 VSUBS 0.00831f
C413 B.n319 VSUBS 0.00831f
C414 B.n320 VSUBS 0.00831f
C415 B.n321 VSUBS 0.00831f
C416 B.n322 VSUBS 0.00831f
C417 B.n323 VSUBS 0.00831f
C418 B.n324 VSUBS 0.00831f
C419 B.n325 VSUBS 0.00831f
C420 B.n326 VSUBS 0.00831f
C421 B.n327 VSUBS 0.00831f
C422 B.n328 VSUBS 0.00831f
C423 B.n329 VSUBS 0.00831f
C424 B.n330 VSUBS 0.00831f
C425 B.n331 VSUBS 0.00831f
C426 B.n332 VSUBS 0.00831f
C427 B.n333 VSUBS 0.00831f
C428 B.n334 VSUBS 0.00831f
C429 B.n335 VSUBS 0.00831f
C430 B.n336 VSUBS 0.00831f
C431 B.n337 VSUBS 0.00831f
C432 B.n338 VSUBS 0.00831f
C433 B.n339 VSUBS 0.010844f
C434 B.n340 VSUBS 0.011552f
C435 B.n341 VSUBS 0.022972f
C436 VDD1.n0 VSUBS 0.017161f
C437 VDD1.n1 VSUBS 0.114996f
C438 VDD1.n2 VSUBS 0.008907f
C439 VDD1.t1 VSUBS 0.046445f
C440 VDD1.n3 VSUBS 0.054401f
C441 VDD1.n4 VSUBS 0.012414f
C442 VDD1.n5 VSUBS 0.01579f
C443 VDD1.n6 VSUBS 0.047382f
C444 VDD1.n7 VSUBS 0.009431f
C445 VDD1.n8 VSUBS 0.008907f
C446 VDD1.n9 VSUBS 0.039674f
C447 VDD1.n10 VSUBS 0.036442f
C448 VDD1.n11 VSUBS 0.017161f
C449 VDD1.n12 VSUBS 0.114996f
C450 VDD1.n13 VSUBS 0.008907f
C451 VDD1.t5 VSUBS 0.046445f
C452 VDD1.n14 VSUBS 0.054401f
C453 VDD1.n15 VSUBS 0.012414f
C454 VDD1.n16 VSUBS 0.01579f
C455 VDD1.n17 VSUBS 0.047382f
C456 VDD1.n18 VSUBS 0.009431f
C457 VDD1.n19 VSUBS 0.008907f
C458 VDD1.n20 VSUBS 0.039674f
C459 VDD1.n21 VSUBS 0.036191f
C460 VDD1.t2 VSUBS 0.032224f
C461 VDD1.t3 VSUBS 0.032224f
C462 VDD1.n22 VSUBS 0.157222f
C463 VDD1.n23 VSUBS 1.02054f
C464 VDD1.t0 VSUBS 0.032224f
C465 VDD1.t4 VSUBS 0.032224f
C466 VDD1.n24 VSUBS 0.156859f
C467 VDD1.n25 VSUBS 1.08003f
C468 VTAIL.t5 VSUBS 0.040479f
C469 VTAIL.t0 VSUBS 0.040479f
C470 VTAIL.n0 VSUBS 0.168008f
C471 VTAIL.n1 VSUBS 0.330196f
C472 VTAIL.n2 VSUBS 0.021557f
C473 VTAIL.n3 VSUBS 0.144459f
C474 VTAIL.n4 VSUBS 0.011189f
C475 VTAIL.t9 VSUBS 0.058345f
C476 VTAIL.n5 VSUBS 0.068339f
C477 VTAIL.n6 VSUBS 0.015594f
C478 VTAIL.n7 VSUBS 0.019836f
C479 VTAIL.n8 VSUBS 0.059521f
C480 VTAIL.n9 VSUBS 0.011848f
C481 VTAIL.n10 VSUBS 0.011189f
C482 VTAIL.n11 VSUBS 0.049838f
C483 VTAIL.n12 VSUBS 0.029784f
C484 VTAIL.n13 VSUBS 0.156123f
C485 VTAIL.t8 VSUBS 0.040479f
C486 VTAIL.t7 VSUBS 0.040479f
C487 VTAIL.n14 VSUBS 0.168008f
C488 VTAIL.n15 VSUBS 0.878693f
C489 VTAIL.t2 VSUBS 0.040479f
C490 VTAIL.t3 VSUBS 0.040479f
C491 VTAIL.n16 VSUBS 0.168009f
C492 VTAIL.n17 VSUBS 0.878692f
C493 VTAIL.n18 VSUBS 0.021557f
C494 VTAIL.n19 VSUBS 0.144459f
C495 VTAIL.n20 VSUBS 0.011189f
C496 VTAIL.t1 VSUBS 0.058345f
C497 VTAIL.n21 VSUBS 0.068339f
C498 VTAIL.n22 VSUBS 0.015594f
C499 VTAIL.n23 VSUBS 0.019836f
C500 VTAIL.n24 VSUBS 0.059521f
C501 VTAIL.n25 VSUBS 0.011848f
C502 VTAIL.n26 VSUBS 0.011189f
C503 VTAIL.n27 VSUBS 0.049838f
C504 VTAIL.n28 VSUBS 0.029784f
C505 VTAIL.n29 VSUBS 0.156123f
C506 VTAIL.t11 VSUBS 0.040479f
C507 VTAIL.t6 VSUBS 0.040479f
C508 VTAIL.n30 VSUBS 0.168009f
C509 VTAIL.n31 VSUBS 0.379216f
C510 VTAIL.n32 VSUBS 0.021557f
C511 VTAIL.n33 VSUBS 0.144459f
C512 VTAIL.n34 VSUBS 0.011189f
C513 VTAIL.t10 VSUBS 0.058345f
C514 VTAIL.n35 VSUBS 0.068339f
C515 VTAIL.n36 VSUBS 0.015594f
C516 VTAIL.n37 VSUBS 0.019836f
C517 VTAIL.n38 VSUBS 0.059521f
C518 VTAIL.n39 VSUBS 0.011848f
C519 VTAIL.n40 VSUBS 0.011189f
C520 VTAIL.n41 VSUBS 0.049838f
C521 VTAIL.n42 VSUBS 0.029784f
C522 VTAIL.n43 VSUBS 0.585032f
C523 VTAIL.n44 VSUBS 0.021557f
C524 VTAIL.n45 VSUBS 0.144459f
C525 VTAIL.n46 VSUBS 0.011189f
C526 VTAIL.t4 VSUBS 0.058345f
C527 VTAIL.n47 VSUBS 0.068339f
C528 VTAIL.n48 VSUBS 0.015594f
C529 VTAIL.n49 VSUBS 0.019836f
C530 VTAIL.n50 VSUBS 0.059521f
C531 VTAIL.n51 VSUBS 0.011848f
C532 VTAIL.n52 VSUBS 0.011189f
C533 VTAIL.n53 VSUBS 0.049838f
C534 VTAIL.n54 VSUBS 0.029784f
C535 VTAIL.n55 VSUBS 0.563486f
C536 VP.n0 VSUBS 0.050118f
C537 VP.t3 VSUBS 0.265843f
C538 VP.n1 VSUBS 0.148385f
C539 VP.n2 VSUBS 0.050118f
C540 VP.n3 VSUBS 0.050118f
C541 VP.t1 VSUBS 0.333762f
C542 VP.t5 VSUBS 0.265843f
C543 VP.n4 VSUBS 0.194658f
C544 VP.t4 VSUBS 0.362063f
C545 VP.n5 VSUBS 0.207029f
C546 VP.n6 VSUBS 0.209641f
C547 VP.n7 VSUBS 0.06449f
C548 VP.n8 VSUBS 0.016212f
C549 VP.n9 VSUBS 0.199872f
C550 VP.n10 VSUBS 1.47029f
C551 VP.n11 VSUBS 1.52233f
C552 VP.t0 VSUBS 0.333762f
C553 VP.n12 VSUBS 0.199872f
C554 VP.n13 VSUBS 0.016212f
C555 VP.n14 VSUBS 0.06449f
C556 VP.n15 VSUBS 0.050118f
C557 VP.n16 VSUBS 0.050118f
C558 VP.n17 VSUBS 0.06449f
C559 VP.n18 VSUBS 0.016212f
C560 VP.t2 VSUBS 0.333762f
C561 VP.n19 VSUBS 0.199872f
C562 VP.n20 VSUBS 0.03884f
.ends

