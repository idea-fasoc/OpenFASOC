* NGSPICE file created from diff_pair_sample_1216.ext - technology: sky130A

.subckt diff_pair_sample_1216 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=0 ps=0 w=8.87 l=3.45
X1 VTAIL.t11 VP.t0 VDD1.t0 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=1.46355 ps=9.2 w=8.87 l=3.45
X2 VDD1.t1 VP.t1 VTAIL.t10 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=3.4593 ps=18.52 w=8.87 l=3.45
X3 VTAIL.t5 VN.t0 VDD2.t5 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=1.46355 ps=9.2 w=8.87 l=3.45
X4 VDD2.t4 VN.t1 VTAIL.t0 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=1.46355 ps=9.2 w=8.87 l=3.45
X5 B.t8 B.t6 B.t7 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=0 ps=0 w=8.87 l=3.45
X6 B.t5 B.t3 B.t4 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=0 ps=0 w=8.87 l=3.45
X7 VTAIL.t4 VN.t2 VDD2.t3 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=1.46355 ps=9.2 w=8.87 l=3.45
X8 B.t2 B.t0 B.t1 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=0 ps=0 w=8.87 l=3.45
X9 VDD2.t2 VN.t3 VTAIL.t3 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=3.4593 ps=18.52 w=8.87 l=3.45
X10 VTAIL.t9 VP.t2 VDD1.t2 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=1.46355 ps=9.2 w=8.87 l=3.45
X11 VDD1.t3 VP.t3 VTAIL.t8 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=1.46355 ps=9.2 w=8.87 l=3.45
X12 VDD2.t1 VN.t4 VTAIL.t2 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=3.4593 ps=18.52 w=8.87 l=3.45
X13 VDD1.t4 VP.t4 VTAIL.t7 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=1.46355 ps=9.2 w=8.87 l=3.45
X14 VDD1.t5 VP.t5 VTAIL.t6 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=1.46355 pd=9.2 as=3.4593 ps=18.52 w=8.87 l=3.45
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n3994_n2742# sky130_fd_pr__pfet_01v8 ad=3.4593 pd=18.52 as=1.46355 ps=9.2 w=8.87 l=3.45
R0 B.n378 B.n377 585
R1 B.n376 B.n123 585
R2 B.n375 B.n374 585
R3 B.n373 B.n124 585
R4 B.n372 B.n371 585
R5 B.n370 B.n125 585
R6 B.n369 B.n368 585
R7 B.n367 B.n126 585
R8 B.n366 B.n365 585
R9 B.n364 B.n127 585
R10 B.n363 B.n362 585
R11 B.n361 B.n128 585
R12 B.n360 B.n359 585
R13 B.n358 B.n129 585
R14 B.n357 B.n356 585
R15 B.n355 B.n130 585
R16 B.n354 B.n353 585
R17 B.n352 B.n131 585
R18 B.n351 B.n350 585
R19 B.n349 B.n132 585
R20 B.n348 B.n347 585
R21 B.n346 B.n133 585
R22 B.n345 B.n344 585
R23 B.n343 B.n134 585
R24 B.n342 B.n341 585
R25 B.n340 B.n135 585
R26 B.n339 B.n338 585
R27 B.n337 B.n136 585
R28 B.n336 B.n335 585
R29 B.n334 B.n137 585
R30 B.n333 B.n332 585
R31 B.n331 B.n138 585
R32 B.n330 B.n329 585
R33 B.n325 B.n139 585
R34 B.n324 B.n323 585
R35 B.n322 B.n140 585
R36 B.n321 B.n320 585
R37 B.n319 B.n141 585
R38 B.n318 B.n317 585
R39 B.n316 B.n142 585
R40 B.n315 B.n314 585
R41 B.n313 B.n143 585
R42 B.n311 B.n310 585
R43 B.n309 B.n146 585
R44 B.n308 B.n307 585
R45 B.n306 B.n147 585
R46 B.n305 B.n304 585
R47 B.n303 B.n148 585
R48 B.n302 B.n301 585
R49 B.n300 B.n149 585
R50 B.n299 B.n298 585
R51 B.n297 B.n150 585
R52 B.n296 B.n295 585
R53 B.n294 B.n151 585
R54 B.n293 B.n292 585
R55 B.n291 B.n152 585
R56 B.n290 B.n289 585
R57 B.n288 B.n153 585
R58 B.n287 B.n286 585
R59 B.n285 B.n154 585
R60 B.n284 B.n283 585
R61 B.n282 B.n155 585
R62 B.n281 B.n280 585
R63 B.n279 B.n156 585
R64 B.n278 B.n277 585
R65 B.n276 B.n157 585
R66 B.n275 B.n274 585
R67 B.n273 B.n158 585
R68 B.n272 B.n271 585
R69 B.n270 B.n159 585
R70 B.n269 B.n268 585
R71 B.n267 B.n160 585
R72 B.n266 B.n265 585
R73 B.n264 B.n161 585
R74 B.n379 B.n122 585
R75 B.n381 B.n380 585
R76 B.n382 B.n121 585
R77 B.n384 B.n383 585
R78 B.n385 B.n120 585
R79 B.n387 B.n386 585
R80 B.n388 B.n119 585
R81 B.n390 B.n389 585
R82 B.n391 B.n118 585
R83 B.n393 B.n392 585
R84 B.n394 B.n117 585
R85 B.n396 B.n395 585
R86 B.n397 B.n116 585
R87 B.n399 B.n398 585
R88 B.n400 B.n115 585
R89 B.n402 B.n401 585
R90 B.n403 B.n114 585
R91 B.n405 B.n404 585
R92 B.n406 B.n113 585
R93 B.n408 B.n407 585
R94 B.n409 B.n112 585
R95 B.n411 B.n410 585
R96 B.n412 B.n111 585
R97 B.n414 B.n413 585
R98 B.n415 B.n110 585
R99 B.n417 B.n416 585
R100 B.n418 B.n109 585
R101 B.n420 B.n419 585
R102 B.n421 B.n108 585
R103 B.n423 B.n422 585
R104 B.n424 B.n107 585
R105 B.n426 B.n425 585
R106 B.n427 B.n106 585
R107 B.n429 B.n428 585
R108 B.n430 B.n105 585
R109 B.n432 B.n431 585
R110 B.n433 B.n104 585
R111 B.n435 B.n434 585
R112 B.n436 B.n103 585
R113 B.n438 B.n437 585
R114 B.n439 B.n102 585
R115 B.n441 B.n440 585
R116 B.n442 B.n101 585
R117 B.n444 B.n443 585
R118 B.n445 B.n100 585
R119 B.n447 B.n446 585
R120 B.n448 B.n99 585
R121 B.n450 B.n449 585
R122 B.n451 B.n98 585
R123 B.n453 B.n452 585
R124 B.n454 B.n97 585
R125 B.n456 B.n455 585
R126 B.n457 B.n96 585
R127 B.n459 B.n458 585
R128 B.n460 B.n95 585
R129 B.n462 B.n461 585
R130 B.n463 B.n94 585
R131 B.n465 B.n464 585
R132 B.n466 B.n93 585
R133 B.n468 B.n467 585
R134 B.n469 B.n92 585
R135 B.n471 B.n470 585
R136 B.n472 B.n91 585
R137 B.n474 B.n473 585
R138 B.n475 B.n90 585
R139 B.n477 B.n476 585
R140 B.n478 B.n89 585
R141 B.n480 B.n479 585
R142 B.n481 B.n88 585
R143 B.n483 B.n482 585
R144 B.n484 B.n87 585
R145 B.n486 B.n485 585
R146 B.n487 B.n86 585
R147 B.n489 B.n488 585
R148 B.n490 B.n85 585
R149 B.n492 B.n491 585
R150 B.n493 B.n84 585
R151 B.n495 B.n494 585
R152 B.n496 B.n83 585
R153 B.n498 B.n497 585
R154 B.n499 B.n82 585
R155 B.n501 B.n500 585
R156 B.n502 B.n81 585
R157 B.n504 B.n503 585
R158 B.n505 B.n80 585
R159 B.n507 B.n506 585
R160 B.n508 B.n79 585
R161 B.n510 B.n509 585
R162 B.n511 B.n78 585
R163 B.n513 B.n512 585
R164 B.n514 B.n77 585
R165 B.n516 B.n515 585
R166 B.n517 B.n76 585
R167 B.n519 B.n518 585
R168 B.n520 B.n75 585
R169 B.n522 B.n521 585
R170 B.n523 B.n74 585
R171 B.n525 B.n524 585
R172 B.n526 B.n73 585
R173 B.n528 B.n527 585
R174 B.n529 B.n72 585
R175 B.n531 B.n530 585
R176 B.n532 B.n71 585
R177 B.n534 B.n533 585
R178 B.n535 B.n70 585
R179 B.n537 B.n536 585
R180 B.n649 B.n28 585
R181 B.n648 B.n647 585
R182 B.n646 B.n29 585
R183 B.n645 B.n644 585
R184 B.n643 B.n30 585
R185 B.n642 B.n641 585
R186 B.n640 B.n31 585
R187 B.n639 B.n638 585
R188 B.n637 B.n32 585
R189 B.n636 B.n635 585
R190 B.n634 B.n33 585
R191 B.n633 B.n632 585
R192 B.n631 B.n34 585
R193 B.n630 B.n629 585
R194 B.n628 B.n35 585
R195 B.n627 B.n626 585
R196 B.n625 B.n36 585
R197 B.n624 B.n623 585
R198 B.n622 B.n37 585
R199 B.n621 B.n620 585
R200 B.n619 B.n38 585
R201 B.n618 B.n617 585
R202 B.n616 B.n39 585
R203 B.n615 B.n614 585
R204 B.n613 B.n40 585
R205 B.n612 B.n611 585
R206 B.n610 B.n41 585
R207 B.n609 B.n608 585
R208 B.n607 B.n42 585
R209 B.n606 B.n605 585
R210 B.n604 B.n43 585
R211 B.n603 B.n602 585
R212 B.n601 B.n600 585
R213 B.n599 B.n47 585
R214 B.n598 B.n597 585
R215 B.n596 B.n48 585
R216 B.n595 B.n594 585
R217 B.n593 B.n49 585
R218 B.n592 B.n591 585
R219 B.n590 B.n50 585
R220 B.n589 B.n588 585
R221 B.n587 B.n51 585
R222 B.n585 B.n584 585
R223 B.n583 B.n54 585
R224 B.n582 B.n581 585
R225 B.n580 B.n55 585
R226 B.n579 B.n578 585
R227 B.n577 B.n56 585
R228 B.n576 B.n575 585
R229 B.n574 B.n57 585
R230 B.n573 B.n572 585
R231 B.n571 B.n58 585
R232 B.n570 B.n569 585
R233 B.n568 B.n59 585
R234 B.n567 B.n566 585
R235 B.n565 B.n60 585
R236 B.n564 B.n563 585
R237 B.n562 B.n61 585
R238 B.n561 B.n560 585
R239 B.n559 B.n62 585
R240 B.n558 B.n557 585
R241 B.n556 B.n63 585
R242 B.n555 B.n554 585
R243 B.n553 B.n64 585
R244 B.n552 B.n551 585
R245 B.n550 B.n65 585
R246 B.n549 B.n548 585
R247 B.n547 B.n66 585
R248 B.n546 B.n545 585
R249 B.n544 B.n67 585
R250 B.n543 B.n542 585
R251 B.n541 B.n68 585
R252 B.n540 B.n539 585
R253 B.n538 B.n69 585
R254 B.n651 B.n650 585
R255 B.n652 B.n27 585
R256 B.n654 B.n653 585
R257 B.n655 B.n26 585
R258 B.n657 B.n656 585
R259 B.n658 B.n25 585
R260 B.n660 B.n659 585
R261 B.n661 B.n24 585
R262 B.n663 B.n662 585
R263 B.n664 B.n23 585
R264 B.n666 B.n665 585
R265 B.n667 B.n22 585
R266 B.n669 B.n668 585
R267 B.n670 B.n21 585
R268 B.n672 B.n671 585
R269 B.n673 B.n20 585
R270 B.n675 B.n674 585
R271 B.n676 B.n19 585
R272 B.n678 B.n677 585
R273 B.n679 B.n18 585
R274 B.n681 B.n680 585
R275 B.n682 B.n17 585
R276 B.n684 B.n683 585
R277 B.n685 B.n16 585
R278 B.n687 B.n686 585
R279 B.n688 B.n15 585
R280 B.n690 B.n689 585
R281 B.n691 B.n14 585
R282 B.n693 B.n692 585
R283 B.n694 B.n13 585
R284 B.n696 B.n695 585
R285 B.n697 B.n12 585
R286 B.n699 B.n698 585
R287 B.n700 B.n11 585
R288 B.n702 B.n701 585
R289 B.n703 B.n10 585
R290 B.n705 B.n704 585
R291 B.n706 B.n9 585
R292 B.n708 B.n707 585
R293 B.n709 B.n8 585
R294 B.n711 B.n710 585
R295 B.n712 B.n7 585
R296 B.n714 B.n713 585
R297 B.n715 B.n6 585
R298 B.n717 B.n716 585
R299 B.n718 B.n5 585
R300 B.n720 B.n719 585
R301 B.n721 B.n4 585
R302 B.n723 B.n722 585
R303 B.n724 B.n3 585
R304 B.n726 B.n725 585
R305 B.n727 B.n0 585
R306 B.n2 B.n1 585
R307 B.n188 B.n187 585
R308 B.n189 B.n186 585
R309 B.n191 B.n190 585
R310 B.n192 B.n185 585
R311 B.n194 B.n193 585
R312 B.n195 B.n184 585
R313 B.n197 B.n196 585
R314 B.n198 B.n183 585
R315 B.n200 B.n199 585
R316 B.n201 B.n182 585
R317 B.n203 B.n202 585
R318 B.n204 B.n181 585
R319 B.n206 B.n205 585
R320 B.n207 B.n180 585
R321 B.n209 B.n208 585
R322 B.n210 B.n179 585
R323 B.n212 B.n211 585
R324 B.n213 B.n178 585
R325 B.n215 B.n214 585
R326 B.n216 B.n177 585
R327 B.n218 B.n217 585
R328 B.n219 B.n176 585
R329 B.n221 B.n220 585
R330 B.n222 B.n175 585
R331 B.n224 B.n223 585
R332 B.n225 B.n174 585
R333 B.n227 B.n226 585
R334 B.n228 B.n173 585
R335 B.n230 B.n229 585
R336 B.n231 B.n172 585
R337 B.n233 B.n232 585
R338 B.n234 B.n171 585
R339 B.n236 B.n235 585
R340 B.n237 B.n170 585
R341 B.n239 B.n238 585
R342 B.n240 B.n169 585
R343 B.n242 B.n241 585
R344 B.n243 B.n168 585
R345 B.n245 B.n244 585
R346 B.n246 B.n167 585
R347 B.n248 B.n247 585
R348 B.n249 B.n166 585
R349 B.n251 B.n250 585
R350 B.n252 B.n165 585
R351 B.n254 B.n253 585
R352 B.n255 B.n164 585
R353 B.n257 B.n256 585
R354 B.n258 B.n163 585
R355 B.n260 B.n259 585
R356 B.n261 B.n162 585
R357 B.n263 B.n262 585
R358 B.n262 B.n161 545.355
R359 B.n379 B.n378 545.355
R360 B.n536 B.n69 545.355
R361 B.n650 B.n649 545.355
R362 B.n144 B.t9 271.01
R363 B.n326 B.t6 271.01
R364 B.n52 B.t3 271.01
R365 B.n44 B.t0 271.01
R366 B.n729 B.n728 256.663
R367 B.n728 B.n727 235.042
R368 B.n728 B.n2 235.042
R369 B.n326 B.t7 182.038
R370 B.n52 B.t5 182.038
R371 B.n144 B.t10 182.028
R372 B.n44 B.t2 182.028
R373 B.n266 B.n161 163.367
R374 B.n267 B.n266 163.367
R375 B.n268 B.n267 163.367
R376 B.n268 B.n159 163.367
R377 B.n272 B.n159 163.367
R378 B.n273 B.n272 163.367
R379 B.n274 B.n273 163.367
R380 B.n274 B.n157 163.367
R381 B.n278 B.n157 163.367
R382 B.n279 B.n278 163.367
R383 B.n280 B.n279 163.367
R384 B.n280 B.n155 163.367
R385 B.n284 B.n155 163.367
R386 B.n285 B.n284 163.367
R387 B.n286 B.n285 163.367
R388 B.n286 B.n153 163.367
R389 B.n290 B.n153 163.367
R390 B.n291 B.n290 163.367
R391 B.n292 B.n291 163.367
R392 B.n292 B.n151 163.367
R393 B.n296 B.n151 163.367
R394 B.n297 B.n296 163.367
R395 B.n298 B.n297 163.367
R396 B.n298 B.n149 163.367
R397 B.n302 B.n149 163.367
R398 B.n303 B.n302 163.367
R399 B.n304 B.n303 163.367
R400 B.n304 B.n147 163.367
R401 B.n308 B.n147 163.367
R402 B.n309 B.n308 163.367
R403 B.n310 B.n309 163.367
R404 B.n310 B.n143 163.367
R405 B.n315 B.n143 163.367
R406 B.n316 B.n315 163.367
R407 B.n317 B.n316 163.367
R408 B.n317 B.n141 163.367
R409 B.n321 B.n141 163.367
R410 B.n322 B.n321 163.367
R411 B.n323 B.n322 163.367
R412 B.n323 B.n139 163.367
R413 B.n330 B.n139 163.367
R414 B.n331 B.n330 163.367
R415 B.n332 B.n331 163.367
R416 B.n332 B.n137 163.367
R417 B.n336 B.n137 163.367
R418 B.n337 B.n336 163.367
R419 B.n338 B.n337 163.367
R420 B.n338 B.n135 163.367
R421 B.n342 B.n135 163.367
R422 B.n343 B.n342 163.367
R423 B.n344 B.n343 163.367
R424 B.n344 B.n133 163.367
R425 B.n348 B.n133 163.367
R426 B.n349 B.n348 163.367
R427 B.n350 B.n349 163.367
R428 B.n350 B.n131 163.367
R429 B.n354 B.n131 163.367
R430 B.n355 B.n354 163.367
R431 B.n356 B.n355 163.367
R432 B.n356 B.n129 163.367
R433 B.n360 B.n129 163.367
R434 B.n361 B.n360 163.367
R435 B.n362 B.n361 163.367
R436 B.n362 B.n127 163.367
R437 B.n366 B.n127 163.367
R438 B.n367 B.n366 163.367
R439 B.n368 B.n367 163.367
R440 B.n368 B.n125 163.367
R441 B.n372 B.n125 163.367
R442 B.n373 B.n372 163.367
R443 B.n374 B.n373 163.367
R444 B.n374 B.n123 163.367
R445 B.n378 B.n123 163.367
R446 B.n536 B.n535 163.367
R447 B.n535 B.n534 163.367
R448 B.n534 B.n71 163.367
R449 B.n530 B.n71 163.367
R450 B.n530 B.n529 163.367
R451 B.n529 B.n528 163.367
R452 B.n528 B.n73 163.367
R453 B.n524 B.n73 163.367
R454 B.n524 B.n523 163.367
R455 B.n523 B.n522 163.367
R456 B.n522 B.n75 163.367
R457 B.n518 B.n75 163.367
R458 B.n518 B.n517 163.367
R459 B.n517 B.n516 163.367
R460 B.n516 B.n77 163.367
R461 B.n512 B.n77 163.367
R462 B.n512 B.n511 163.367
R463 B.n511 B.n510 163.367
R464 B.n510 B.n79 163.367
R465 B.n506 B.n79 163.367
R466 B.n506 B.n505 163.367
R467 B.n505 B.n504 163.367
R468 B.n504 B.n81 163.367
R469 B.n500 B.n81 163.367
R470 B.n500 B.n499 163.367
R471 B.n499 B.n498 163.367
R472 B.n498 B.n83 163.367
R473 B.n494 B.n83 163.367
R474 B.n494 B.n493 163.367
R475 B.n493 B.n492 163.367
R476 B.n492 B.n85 163.367
R477 B.n488 B.n85 163.367
R478 B.n488 B.n487 163.367
R479 B.n487 B.n486 163.367
R480 B.n486 B.n87 163.367
R481 B.n482 B.n87 163.367
R482 B.n482 B.n481 163.367
R483 B.n481 B.n480 163.367
R484 B.n480 B.n89 163.367
R485 B.n476 B.n89 163.367
R486 B.n476 B.n475 163.367
R487 B.n475 B.n474 163.367
R488 B.n474 B.n91 163.367
R489 B.n470 B.n91 163.367
R490 B.n470 B.n469 163.367
R491 B.n469 B.n468 163.367
R492 B.n468 B.n93 163.367
R493 B.n464 B.n93 163.367
R494 B.n464 B.n463 163.367
R495 B.n463 B.n462 163.367
R496 B.n462 B.n95 163.367
R497 B.n458 B.n95 163.367
R498 B.n458 B.n457 163.367
R499 B.n457 B.n456 163.367
R500 B.n456 B.n97 163.367
R501 B.n452 B.n97 163.367
R502 B.n452 B.n451 163.367
R503 B.n451 B.n450 163.367
R504 B.n450 B.n99 163.367
R505 B.n446 B.n99 163.367
R506 B.n446 B.n445 163.367
R507 B.n445 B.n444 163.367
R508 B.n444 B.n101 163.367
R509 B.n440 B.n101 163.367
R510 B.n440 B.n439 163.367
R511 B.n439 B.n438 163.367
R512 B.n438 B.n103 163.367
R513 B.n434 B.n103 163.367
R514 B.n434 B.n433 163.367
R515 B.n433 B.n432 163.367
R516 B.n432 B.n105 163.367
R517 B.n428 B.n105 163.367
R518 B.n428 B.n427 163.367
R519 B.n427 B.n426 163.367
R520 B.n426 B.n107 163.367
R521 B.n422 B.n107 163.367
R522 B.n422 B.n421 163.367
R523 B.n421 B.n420 163.367
R524 B.n420 B.n109 163.367
R525 B.n416 B.n109 163.367
R526 B.n416 B.n415 163.367
R527 B.n415 B.n414 163.367
R528 B.n414 B.n111 163.367
R529 B.n410 B.n111 163.367
R530 B.n410 B.n409 163.367
R531 B.n409 B.n408 163.367
R532 B.n408 B.n113 163.367
R533 B.n404 B.n113 163.367
R534 B.n404 B.n403 163.367
R535 B.n403 B.n402 163.367
R536 B.n402 B.n115 163.367
R537 B.n398 B.n115 163.367
R538 B.n398 B.n397 163.367
R539 B.n397 B.n396 163.367
R540 B.n396 B.n117 163.367
R541 B.n392 B.n117 163.367
R542 B.n392 B.n391 163.367
R543 B.n391 B.n390 163.367
R544 B.n390 B.n119 163.367
R545 B.n386 B.n119 163.367
R546 B.n386 B.n385 163.367
R547 B.n385 B.n384 163.367
R548 B.n384 B.n121 163.367
R549 B.n380 B.n121 163.367
R550 B.n380 B.n379 163.367
R551 B.n649 B.n648 163.367
R552 B.n648 B.n29 163.367
R553 B.n644 B.n29 163.367
R554 B.n644 B.n643 163.367
R555 B.n643 B.n642 163.367
R556 B.n642 B.n31 163.367
R557 B.n638 B.n31 163.367
R558 B.n638 B.n637 163.367
R559 B.n637 B.n636 163.367
R560 B.n636 B.n33 163.367
R561 B.n632 B.n33 163.367
R562 B.n632 B.n631 163.367
R563 B.n631 B.n630 163.367
R564 B.n630 B.n35 163.367
R565 B.n626 B.n35 163.367
R566 B.n626 B.n625 163.367
R567 B.n625 B.n624 163.367
R568 B.n624 B.n37 163.367
R569 B.n620 B.n37 163.367
R570 B.n620 B.n619 163.367
R571 B.n619 B.n618 163.367
R572 B.n618 B.n39 163.367
R573 B.n614 B.n39 163.367
R574 B.n614 B.n613 163.367
R575 B.n613 B.n612 163.367
R576 B.n612 B.n41 163.367
R577 B.n608 B.n41 163.367
R578 B.n608 B.n607 163.367
R579 B.n607 B.n606 163.367
R580 B.n606 B.n43 163.367
R581 B.n602 B.n43 163.367
R582 B.n602 B.n601 163.367
R583 B.n601 B.n47 163.367
R584 B.n597 B.n47 163.367
R585 B.n597 B.n596 163.367
R586 B.n596 B.n595 163.367
R587 B.n595 B.n49 163.367
R588 B.n591 B.n49 163.367
R589 B.n591 B.n590 163.367
R590 B.n590 B.n589 163.367
R591 B.n589 B.n51 163.367
R592 B.n584 B.n51 163.367
R593 B.n584 B.n583 163.367
R594 B.n583 B.n582 163.367
R595 B.n582 B.n55 163.367
R596 B.n578 B.n55 163.367
R597 B.n578 B.n577 163.367
R598 B.n577 B.n576 163.367
R599 B.n576 B.n57 163.367
R600 B.n572 B.n57 163.367
R601 B.n572 B.n571 163.367
R602 B.n571 B.n570 163.367
R603 B.n570 B.n59 163.367
R604 B.n566 B.n59 163.367
R605 B.n566 B.n565 163.367
R606 B.n565 B.n564 163.367
R607 B.n564 B.n61 163.367
R608 B.n560 B.n61 163.367
R609 B.n560 B.n559 163.367
R610 B.n559 B.n558 163.367
R611 B.n558 B.n63 163.367
R612 B.n554 B.n63 163.367
R613 B.n554 B.n553 163.367
R614 B.n553 B.n552 163.367
R615 B.n552 B.n65 163.367
R616 B.n548 B.n65 163.367
R617 B.n548 B.n547 163.367
R618 B.n547 B.n546 163.367
R619 B.n546 B.n67 163.367
R620 B.n542 B.n67 163.367
R621 B.n542 B.n541 163.367
R622 B.n541 B.n540 163.367
R623 B.n540 B.n69 163.367
R624 B.n650 B.n27 163.367
R625 B.n654 B.n27 163.367
R626 B.n655 B.n654 163.367
R627 B.n656 B.n655 163.367
R628 B.n656 B.n25 163.367
R629 B.n660 B.n25 163.367
R630 B.n661 B.n660 163.367
R631 B.n662 B.n661 163.367
R632 B.n662 B.n23 163.367
R633 B.n666 B.n23 163.367
R634 B.n667 B.n666 163.367
R635 B.n668 B.n667 163.367
R636 B.n668 B.n21 163.367
R637 B.n672 B.n21 163.367
R638 B.n673 B.n672 163.367
R639 B.n674 B.n673 163.367
R640 B.n674 B.n19 163.367
R641 B.n678 B.n19 163.367
R642 B.n679 B.n678 163.367
R643 B.n680 B.n679 163.367
R644 B.n680 B.n17 163.367
R645 B.n684 B.n17 163.367
R646 B.n685 B.n684 163.367
R647 B.n686 B.n685 163.367
R648 B.n686 B.n15 163.367
R649 B.n690 B.n15 163.367
R650 B.n691 B.n690 163.367
R651 B.n692 B.n691 163.367
R652 B.n692 B.n13 163.367
R653 B.n696 B.n13 163.367
R654 B.n697 B.n696 163.367
R655 B.n698 B.n697 163.367
R656 B.n698 B.n11 163.367
R657 B.n702 B.n11 163.367
R658 B.n703 B.n702 163.367
R659 B.n704 B.n703 163.367
R660 B.n704 B.n9 163.367
R661 B.n708 B.n9 163.367
R662 B.n709 B.n708 163.367
R663 B.n710 B.n709 163.367
R664 B.n710 B.n7 163.367
R665 B.n714 B.n7 163.367
R666 B.n715 B.n714 163.367
R667 B.n716 B.n715 163.367
R668 B.n716 B.n5 163.367
R669 B.n720 B.n5 163.367
R670 B.n721 B.n720 163.367
R671 B.n722 B.n721 163.367
R672 B.n722 B.n3 163.367
R673 B.n726 B.n3 163.367
R674 B.n727 B.n726 163.367
R675 B.n188 B.n2 163.367
R676 B.n189 B.n188 163.367
R677 B.n190 B.n189 163.367
R678 B.n190 B.n185 163.367
R679 B.n194 B.n185 163.367
R680 B.n195 B.n194 163.367
R681 B.n196 B.n195 163.367
R682 B.n196 B.n183 163.367
R683 B.n200 B.n183 163.367
R684 B.n201 B.n200 163.367
R685 B.n202 B.n201 163.367
R686 B.n202 B.n181 163.367
R687 B.n206 B.n181 163.367
R688 B.n207 B.n206 163.367
R689 B.n208 B.n207 163.367
R690 B.n208 B.n179 163.367
R691 B.n212 B.n179 163.367
R692 B.n213 B.n212 163.367
R693 B.n214 B.n213 163.367
R694 B.n214 B.n177 163.367
R695 B.n218 B.n177 163.367
R696 B.n219 B.n218 163.367
R697 B.n220 B.n219 163.367
R698 B.n220 B.n175 163.367
R699 B.n224 B.n175 163.367
R700 B.n225 B.n224 163.367
R701 B.n226 B.n225 163.367
R702 B.n226 B.n173 163.367
R703 B.n230 B.n173 163.367
R704 B.n231 B.n230 163.367
R705 B.n232 B.n231 163.367
R706 B.n232 B.n171 163.367
R707 B.n236 B.n171 163.367
R708 B.n237 B.n236 163.367
R709 B.n238 B.n237 163.367
R710 B.n238 B.n169 163.367
R711 B.n242 B.n169 163.367
R712 B.n243 B.n242 163.367
R713 B.n244 B.n243 163.367
R714 B.n244 B.n167 163.367
R715 B.n248 B.n167 163.367
R716 B.n249 B.n248 163.367
R717 B.n250 B.n249 163.367
R718 B.n250 B.n165 163.367
R719 B.n254 B.n165 163.367
R720 B.n255 B.n254 163.367
R721 B.n256 B.n255 163.367
R722 B.n256 B.n163 163.367
R723 B.n260 B.n163 163.367
R724 B.n261 B.n260 163.367
R725 B.n262 B.n261 163.367
R726 B.n327 B.t8 108.728
R727 B.n53 B.t4 108.728
R728 B.n145 B.t11 108.719
R729 B.n45 B.t1 108.719
R730 B.n145 B.n144 73.3096
R731 B.n327 B.n326 73.3096
R732 B.n53 B.n52 73.3096
R733 B.n45 B.n44 73.3096
R734 B.n312 B.n145 59.5399
R735 B.n328 B.n327 59.5399
R736 B.n586 B.n53 59.5399
R737 B.n46 B.n45 59.5399
R738 B.n651 B.n28 35.4346
R739 B.n538 B.n537 35.4346
R740 B.n264 B.n263 35.4346
R741 B.n377 B.n122 35.4346
R742 B B.n729 18.0485
R743 B.n652 B.n651 10.6151
R744 B.n653 B.n652 10.6151
R745 B.n653 B.n26 10.6151
R746 B.n657 B.n26 10.6151
R747 B.n658 B.n657 10.6151
R748 B.n659 B.n658 10.6151
R749 B.n659 B.n24 10.6151
R750 B.n663 B.n24 10.6151
R751 B.n664 B.n663 10.6151
R752 B.n665 B.n664 10.6151
R753 B.n665 B.n22 10.6151
R754 B.n669 B.n22 10.6151
R755 B.n670 B.n669 10.6151
R756 B.n671 B.n670 10.6151
R757 B.n671 B.n20 10.6151
R758 B.n675 B.n20 10.6151
R759 B.n676 B.n675 10.6151
R760 B.n677 B.n676 10.6151
R761 B.n677 B.n18 10.6151
R762 B.n681 B.n18 10.6151
R763 B.n682 B.n681 10.6151
R764 B.n683 B.n682 10.6151
R765 B.n683 B.n16 10.6151
R766 B.n687 B.n16 10.6151
R767 B.n688 B.n687 10.6151
R768 B.n689 B.n688 10.6151
R769 B.n689 B.n14 10.6151
R770 B.n693 B.n14 10.6151
R771 B.n694 B.n693 10.6151
R772 B.n695 B.n694 10.6151
R773 B.n695 B.n12 10.6151
R774 B.n699 B.n12 10.6151
R775 B.n700 B.n699 10.6151
R776 B.n701 B.n700 10.6151
R777 B.n701 B.n10 10.6151
R778 B.n705 B.n10 10.6151
R779 B.n706 B.n705 10.6151
R780 B.n707 B.n706 10.6151
R781 B.n707 B.n8 10.6151
R782 B.n711 B.n8 10.6151
R783 B.n712 B.n711 10.6151
R784 B.n713 B.n712 10.6151
R785 B.n713 B.n6 10.6151
R786 B.n717 B.n6 10.6151
R787 B.n718 B.n717 10.6151
R788 B.n719 B.n718 10.6151
R789 B.n719 B.n4 10.6151
R790 B.n723 B.n4 10.6151
R791 B.n724 B.n723 10.6151
R792 B.n725 B.n724 10.6151
R793 B.n725 B.n0 10.6151
R794 B.n647 B.n28 10.6151
R795 B.n647 B.n646 10.6151
R796 B.n646 B.n645 10.6151
R797 B.n645 B.n30 10.6151
R798 B.n641 B.n30 10.6151
R799 B.n641 B.n640 10.6151
R800 B.n640 B.n639 10.6151
R801 B.n639 B.n32 10.6151
R802 B.n635 B.n32 10.6151
R803 B.n635 B.n634 10.6151
R804 B.n634 B.n633 10.6151
R805 B.n633 B.n34 10.6151
R806 B.n629 B.n34 10.6151
R807 B.n629 B.n628 10.6151
R808 B.n628 B.n627 10.6151
R809 B.n627 B.n36 10.6151
R810 B.n623 B.n36 10.6151
R811 B.n623 B.n622 10.6151
R812 B.n622 B.n621 10.6151
R813 B.n621 B.n38 10.6151
R814 B.n617 B.n38 10.6151
R815 B.n617 B.n616 10.6151
R816 B.n616 B.n615 10.6151
R817 B.n615 B.n40 10.6151
R818 B.n611 B.n40 10.6151
R819 B.n611 B.n610 10.6151
R820 B.n610 B.n609 10.6151
R821 B.n609 B.n42 10.6151
R822 B.n605 B.n42 10.6151
R823 B.n605 B.n604 10.6151
R824 B.n604 B.n603 10.6151
R825 B.n600 B.n599 10.6151
R826 B.n599 B.n598 10.6151
R827 B.n598 B.n48 10.6151
R828 B.n594 B.n48 10.6151
R829 B.n594 B.n593 10.6151
R830 B.n593 B.n592 10.6151
R831 B.n592 B.n50 10.6151
R832 B.n588 B.n50 10.6151
R833 B.n588 B.n587 10.6151
R834 B.n585 B.n54 10.6151
R835 B.n581 B.n54 10.6151
R836 B.n581 B.n580 10.6151
R837 B.n580 B.n579 10.6151
R838 B.n579 B.n56 10.6151
R839 B.n575 B.n56 10.6151
R840 B.n575 B.n574 10.6151
R841 B.n574 B.n573 10.6151
R842 B.n573 B.n58 10.6151
R843 B.n569 B.n58 10.6151
R844 B.n569 B.n568 10.6151
R845 B.n568 B.n567 10.6151
R846 B.n567 B.n60 10.6151
R847 B.n563 B.n60 10.6151
R848 B.n563 B.n562 10.6151
R849 B.n562 B.n561 10.6151
R850 B.n561 B.n62 10.6151
R851 B.n557 B.n62 10.6151
R852 B.n557 B.n556 10.6151
R853 B.n556 B.n555 10.6151
R854 B.n555 B.n64 10.6151
R855 B.n551 B.n64 10.6151
R856 B.n551 B.n550 10.6151
R857 B.n550 B.n549 10.6151
R858 B.n549 B.n66 10.6151
R859 B.n545 B.n66 10.6151
R860 B.n545 B.n544 10.6151
R861 B.n544 B.n543 10.6151
R862 B.n543 B.n68 10.6151
R863 B.n539 B.n68 10.6151
R864 B.n539 B.n538 10.6151
R865 B.n537 B.n70 10.6151
R866 B.n533 B.n70 10.6151
R867 B.n533 B.n532 10.6151
R868 B.n532 B.n531 10.6151
R869 B.n531 B.n72 10.6151
R870 B.n527 B.n72 10.6151
R871 B.n527 B.n526 10.6151
R872 B.n526 B.n525 10.6151
R873 B.n525 B.n74 10.6151
R874 B.n521 B.n74 10.6151
R875 B.n521 B.n520 10.6151
R876 B.n520 B.n519 10.6151
R877 B.n519 B.n76 10.6151
R878 B.n515 B.n76 10.6151
R879 B.n515 B.n514 10.6151
R880 B.n514 B.n513 10.6151
R881 B.n513 B.n78 10.6151
R882 B.n509 B.n78 10.6151
R883 B.n509 B.n508 10.6151
R884 B.n508 B.n507 10.6151
R885 B.n507 B.n80 10.6151
R886 B.n503 B.n80 10.6151
R887 B.n503 B.n502 10.6151
R888 B.n502 B.n501 10.6151
R889 B.n501 B.n82 10.6151
R890 B.n497 B.n82 10.6151
R891 B.n497 B.n496 10.6151
R892 B.n496 B.n495 10.6151
R893 B.n495 B.n84 10.6151
R894 B.n491 B.n84 10.6151
R895 B.n491 B.n490 10.6151
R896 B.n490 B.n489 10.6151
R897 B.n489 B.n86 10.6151
R898 B.n485 B.n86 10.6151
R899 B.n485 B.n484 10.6151
R900 B.n484 B.n483 10.6151
R901 B.n483 B.n88 10.6151
R902 B.n479 B.n88 10.6151
R903 B.n479 B.n478 10.6151
R904 B.n478 B.n477 10.6151
R905 B.n477 B.n90 10.6151
R906 B.n473 B.n90 10.6151
R907 B.n473 B.n472 10.6151
R908 B.n472 B.n471 10.6151
R909 B.n471 B.n92 10.6151
R910 B.n467 B.n92 10.6151
R911 B.n467 B.n466 10.6151
R912 B.n466 B.n465 10.6151
R913 B.n465 B.n94 10.6151
R914 B.n461 B.n94 10.6151
R915 B.n461 B.n460 10.6151
R916 B.n460 B.n459 10.6151
R917 B.n459 B.n96 10.6151
R918 B.n455 B.n96 10.6151
R919 B.n455 B.n454 10.6151
R920 B.n454 B.n453 10.6151
R921 B.n453 B.n98 10.6151
R922 B.n449 B.n98 10.6151
R923 B.n449 B.n448 10.6151
R924 B.n448 B.n447 10.6151
R925 B.n447 B.n100 10.6151
R926 B.n443 B.n100 10.6151
R927 B.n443 B.n442 10.6151
R928 B.n442 B.n441 10.6151
R929 B.n441 B.n102 10.6151
R930 B.n437 B.n102 10.6151
R931 B.n437 B.n436 10.6151
R932 B.n436 B.n435 10.6151
R933 B.n435 B.n104 10.6151
R934 B.n431 B.n104 10.6151
R935 B.n431 B.n430 10.6151
R936 B.n430 B.n429 10.6151
R937 B.n429 B.n106 10.6151
R938 B.n425 B.n106 10.6151
R939 B.n425 B.n424 10.6151
R940 B.n424 B.n423 10.6151
R941 B.n423 B.n108 10.6151
R942 B.n419 B.n108 10.6151
R943 B.n419 B.n418 10.6151
R944 B.n418 B.n417 10.6151
R945 B.n417 B.n110 10.6151
R946 B.n413 B.n110 10.6151
R947 B.n413 B.n412 10.6151
R948 B.n412 B.n411 10.6151
R949 B.n411 B.n112 10.6151
R950 B.n407 B.n112 10.6151
R951 B.n407 B.n406 10.6151
R952 B.n406 B.n405 10.6151
R953 B.n405 B.n114 10.6151
R954 B.n401 B.n114 10.6151
R955 B.n401 B.n400 10.6151
R956 B.n400 B.n399 10.6151
R957 B.n399 B.n116 10.6151
R958 B.n395 B.n116 10.6151
R959 B.n395 B.n394 10.6151
R960 B.n394 B.n393 10.6151
R961 B.n393 B.n118 10.6151
R962 B.n389 B.n118 10.6151
R963 B.n389 B.n388 10.6151
R964 B.n388 B.n387 10.6151
R965 B.n387 B.n120 10.6151
R966 B.n383 B.n120 10.6151
R967 B.n383 B.n382 10.6151
R968 B.n382 B.n381 10.6151
R969 B.n381 B.n122 10.6151
R970 B.n187 B.n1 10.6151
R971 B.n187 B.n186 10.6151
R972 B.n191 B.n186 10.6151
R973 B.n192 B.n191 10.6151
R974 B.n193 B.n192 10.6151
R975 B.n193 B.n184 10.6151
R976 B.n197 B.n184 10.6151
R977 B.n198 B.n197 10.6151
R978 B.n199 B.n198 10.6151
R979 B.n199 B.n182 10.6151
R980 B.n203 B.n182 10.6151
R981 B.n204 B.n203 10.6151
R982 B.n205 B.n204 10.6151
R983 B.n205 B.n180 10.6151
R984 B.n209 B.n180 10.6151
R985 B.n210 B.n209 10.6151
R986 B.n211 B.n210 10.6151
R987 B.n211 B.n178 10.6151
R988 B.n215 B.n178 10.6151
R989 B.n216 B.n215 10.6151
R990 B.n217 B.n216 10.6151
R991 B.n217 B.n176 10.6151
R992 B.n221 B.n176 10.6151
R993 B.n222 B.n221 10.6151
R994 B.n223 B.n222 10.6151
R995 B.n223 B.n174 10.6151
R996 B.n227 B.n174 10.6151
R997 B.n228 B.n227 10.6151
R998 B.n229 B.n228 10.6151
R999 B.n229 B.n172 10.6151
R1000 B.n233 B.n172 10.6151
R1001 B.n234 B.n233 10.6151
R1002 B.n235 B.n234 10.6151
R1003 B.n235 B.n170 10.6151
R1004 B.n239 B.n170 10.6151
R1005 B.n240 B.n239 10.6151
R1006 B.n241 B.n240 10.6151
R1007 B.n241 B.n168 10.6151
R1008 B.n245 B.n168 10.6151
R1009 B.n246 B.n245 10.6151
R1010 B.n247 B.n246 10.6151
R1011 B.n247 B.n166 10.6151
R1012 B.n251 B.n166 10.6151
R1013 B.n252 B.n251 10.6151
R1014 B.n253 B.n252 10.6151
R1015 B.n253 B.n164 10.6151
R1016 B.n257 B.n164 10.6151
R1017 B.n258 B.n257 10.6151
R1018 B.n259 B.n258 10.6151
R1019 B.n259 B.n162 10.6151
R1020 B.n263 B.n162 10.6151
R1021 B.n265 B.n264 10.6151
R1022 B.n265 B.n160 10.6151
R1023 B.n269 B.n160 10.6151
R1024 B.n270 B.n269 10.6151
R1025 B.n271 B.n270 10.6151
R1026 B.n271 B.n158 10.6151
R1027 B.n275 B.n158 10.6151
R1028 B.n276 B.n275 10.6151
R1029 B.n277 B.n276 10.6151
R1030 B.n277 B.n156 10.6151
R1031 B.n281 B.n156 10.6151
R1032 B.n282 B.n281 10.6151
R1033 B.n283 B.n282 10.6151
R1034 B.n283 B.n154 10.6151
R1035 B.n287 B.n154 10.6151
R1036 B.n288 B.n287 10.6151
R1037 B.n289 B.n288 10.6151
R1038 B.n289 B.n152 10.6151
R1039 B.n293 B.n152 10.6151
R1040 B.n294 B.n293 10.6151
R1041 B.n295 B.n294 10.6151
R1042 B.n295 B.n150 10.6151
R1043 B.n299 B.n150 10.6151
R1044 B.n300 B.n299 10.6151
R1045 B.n301 B.n300 10.6151
R1046 B.n301 B.n148 10.6151
R1047 B.n305 B.n148 10.6151
R1048 B.n306 B.n305 10.6151
R1049 B.n307 B.n306 10.6151
R1050 B.n307 B.n146 10.6151
R1051 B.n311 B.n146 10.6151
R1052 B.n314 B.n313 10.6151
R1053 B.n314 B.n142 10.6151
R1054 B.n318 B.n142 10.6151
R1055 B.n319 B.n318 10.6151
R1056 B.n320 B.n319 10.6151
R1057 B.n320 B.n140 10.6151
R1058 B.n324 B.n140 10.6151
R1059 B.n325 B.n324 10.6151
R1060 B.n329 B.n325 10.6151
R1061 B.n333 B.n138 10.6151
R1062 B.n334 B.n333 10.6151
R1063 B.n335 B.n334 10.6151
R1064 B.n335 B.n136 10.6151
R1065 B.n339 B.n136 10.6151
R1066 B.n340 B.n339 10.6151
R1067 B.n341 B.n340 10.6151
R1068 B.n341 B.n134 10.6151
R1069 B.n345 B.n134 10.6151
R1070 B.n346 B.n345 10.6151
R1071 B.n347 B.n346 10.6151
R1072 B.n347 B.n132 10.6151
R1073 B.n351 B.n132 10.6151
R1074 B.n352 B.n351 10.6151
R1075 B.n353 B.n352 10.6151
R1076 B.n353 B.n130 10.6151
R1077 B.n357 B.n130 10.6151
R1078 B.n358 B.n357 10.6151
R1079 B.n359 B.n358 10.6151
R1080 B.n359 B.n128 10.6151
R1081 B.n363 B.n128 10.6151
R1082 B.n364 B.n363 10.6151
R1083 B.n365 B.n364 10.6151
R1084 B.n365 B.n126 10.6151
R1085 B.n369 B.n126 10.6151
R1086 B.n370 B.n369 10.6151
R1087 B.n371 B.n370 10.6151
R1088 B.n371 B.n124 10.6151
R1089 B.n375 B.n124 10.6151
R1090 B.n376 B.n375 10.6151
R1091 B.n377 B.n376 10.6151
R1092 B.n603 B.n46 9.36635
R1093 B.n586 B.n585 9.36635
R1094 B.n312 B.n311 9.36635
R1095 B.n328 B.n138 9.36635
R1096 B.n729 B.n0 8.11757
R1097 B.n729 B.n1 8.11757
R1098 B.n600 B.n46 1.24928
R1099 B.n587 B.n586 1.24928
R1100 B.n313 B.n312 1.24928
R1101 B.n329 B.n328 1.24928
R1102 VP.n16 VP.n15 161.3
R1103 VP.n17 VP.n12 161.3
R1104 VP.n19 VP.n18 161.3
R1105 VP.n20 VP.n11 161.3
R1106 VP.n22 VP.n21 161.3
R1107 VP.n23 VP.n10 161.3
R1108 VP.n25 VP.n24 161.3
R1109 VP.n50 VP.n49 161.3
R1110 VP.n48 VP.n1 161.3
R1111 VP.n47 VP.n46 161.3
R1112 VP.n45 VP.n2 161.3
R1113 VP.n44 VP.n43 161.3
R1114 VP.n42 VP.n3 161.3
R1115 VP.n41 VP.n40 161.3
R1116 VP.n39 VP.n4 161.3
R1117 VP.n38 VP.n37 161.3
R1118 VP.n36 VP.n5 161.3
R1119 VP.n35 VP.n34 161.3
R1120 VP.n33 VP.n6 161.3
R1121 VP.n32 VP.n31 161.3
R1122 VP.n30 VP.n7 161.3
R1123 VP.n29 VP.n28 161.3
R1124 VP.n14 VP.t3 95.9312
R1125 VP.n27 VP.n8 76.3659
R1126 VP.n51 VP.n0 76.3659
R1127 VP.n26 VP.n9 76.3659
R1128 VP.n4 VP.t2 61.9619
R1129 VP.n8 VP.t4 61.9619
R1130 VP.n0 VP.t1 61.9619
R1131 VP.n13 VP.t0 61.9619
R1132 VP.n9 VP.t5 61.9619
R1133 VP.n35 VP.n6 51.1773
R1134 VP.n43 VP.n2 51.1773
R1135 VP.n18 VP.n11 51.1773
R1136 VP.n14 VP.n13 50.1803
R1137 VP.n27 VP.n26 49.7721
R1138 VP.n31 VP.n6 29.8095
R1139 VP.n47 VP.n2 29.8095
R1140 VP.n22 VP.n11 29.8095
R1141 VP.n30 VP.n29 24.4675
R1142 VP.n31 VP.n30 24.4675
R1143 VP.n36 VP.n35 24.4675
R1144 VP.n37 VP.n36 24.4675
R1145 VP.n37 VP.n4 24.4675
R1146 VP.n41 VP.n4 24.4675
R1147 VP.n42 VP.n41 24.4675
R1148 VP.n43 VP.n42 24.4675
R1149 VP.n48 VP.n47 24.4675
R1150 VP.n49 VP.n48 24.4675
R1151 VP.n23 VP.n22 24.4675
R1152 VP.n24 VP.n23 24.4675
R1153 VP.n16 VP.n13 24.4675
R1154 VP.n17 VP.n16 24.4675
R1155 VP.n18 VP.n17 24.4675
R1156 VP.n29 VP.n8 13.702
R1157 VP.n49 VP.n0 13.702
R1158 VP.n24 VP.n9 13.702
R1159 VP.n15 VP.n14 3.0269
R1160 VP.n26 VP.n25 0.354971
R1161 VP.n28 VP.n27 0.354971
R1162 VP.n51 VP.n50 0.354971
R1163 VP VP.n51 0.26696
R1164 VP.n15 VP.n12 0.189894
R1165 VP.n19 VP.n12 0.189894
R1166 VP.n20 VP.n19 0.189894
R1167 VP.n21 VP.n20 0.189894
R1168 VP.n21 VP.n10 0.189894
R1169 VP.n25 VP.n10 0.189894
R1170 VP.n28 VP.n7 0.189894
R1171 VP.n32 VP.n7 0.189894
R1172 VP.n33 VP.n32 0.189894
R1173 VP.n34 VP.n33 0.189894
R1174 VP.n34 VP.n5 0.189894
R1175 VP.n38 VP.n5 0.189894
R1176 VP.n39 VP.n38 0.189894
R1177 VP.n40 VP.n39 0.189894
R1178 VP.n40 VP.n3 0.189894
R1179 VP.n44 VP.n3 0.189894
R1180 VP.n45 VP.n44 0.189894
R1181 VP.n46 VP.n45 0.189894
R1182 VP.n46 VP.n1 0.189894
R1183 VP.n50 VP.n1 0.189894
R1184 VDD1 VDD1.t3 85.3784
R1185 VDD1.n1 VDD1.t4 85.2645
R1186 VDD1.n1 VDD1.n0 79.9706
R1187 VDD1.n3 VDD1.n2 79.2114
R1188 VDD1.n3 VDD1.n1 44.1647
R1189 VDD1.n2 VDD1.t0 3.6651
R1190 VDD1.n2 VDD1.t5 3.6651
R1191 VDD1.n0 VDD1.t2 3.6651
R1192 VDD1.n0 VDD1.t1 3.6651
R1193 VDD1 VDD1.n3 0.756965
R1194 VTAIL.n7 VTAIL.t3 66.1974
R1195 VTAIL.n10 VTAIL.t6 66.1971
R1196 VTAIL.n11 VTAIL.t2 66.1971
R1197 VTAIL.n2 VTAIL.t10 66.1971
R1198 VTAIL.n9 VTAIL.n8 62.5328
R1199 VTAIL.n6 VTAIL.n5 62.5328
R1200 VTAIL.n1 VTAIL.n0 62.5325
R1201 VTAIL.n4 VTAIL.n3 62.5325
R1202 VTAIL.n6 VTAIL.n4 26.5307
R1203 VTAIL.n11 VTAIL.n10 23.2721
R1204 VTAIL.n0 VTAIL.t1 3.6651
R1205 VTAIL.n0 VTAIL.t4 3.6651
R1206 VTAIL.n3 VTAIL.t7 3.6651
R1207 VTAIL.n3 VTAIL.t9 3.6651
R1208 VTAIL.n8 VTAIL.t8 3.6651
R1209 VTAIL.n8 VTAIL.t11 3.6651
R1210 VTAIL.n5 VTAIL.t0 3.6651
R1211 VTAIL.n5 VTAIL.t5 3.6651
R1212 VTAIL.n7 VTAIL.n6 3.25912
R1213 VTAIL.n10 VTAIL.n9 3.25912
R1214 VTAIL.n4 VTAIL.n2 3.25912
R1215 VTAIL VTAIL.n11 2.38628
R1216 VTAIL.n9 VTAIL.n7 2.09964
R1217 VTAIL.n2 VTAIL.n1 2.09964
R1218 VTAIL VTAIL.n1 0.873345
R1219 VN.n34 VN.n33 161.3
R1220 VN.n32 VN.n19 161.3
R1221 VN.n31 VN.n30 161.3
R1222 VN.n29 VN.n20 161.3
R1223 VN.n28 VN.n27 161.3
R1224 VN.n26 VN.n21 161.3
R1225 VN.n25 VN.n24 161.3
R1226 VN.n16 VN.n15 161.3
R1227 VN.n14 VN.n1 161.3
R1228 VN.n13 VN.n12 161.3
R1229 VN.n11 VN.n2 161.3
R1230 VN.n10 VN.n9 161.3
R1231 VN.n8 VN.n3 161.3
R1232 VN.n7 VN.n6 161.3
R1233 VN.n23 VN.t3 95.9314
R1234 VN.n5 VN.t5 95.9314
R1235 VN.n17 VN.n0 76.3659
R1236 VN.n35 VN.n18 76.3659
R1237 VN.n4 VN.t2 61.9619
R1238 VN.n0 VN.t4 61.9619
R1239 VN.n22 VN.t0 61.9619
R1240 VN.n18 VN.t1 61.9619
R1241 VN.n9 VN.n2 51.1773
R1242 VN.n27 VN.n20 51.1773
R1243 VN.n23 VN.n22 50.1803
R1244 VN.n5 VN.n4 50.1803
R1245 VN VN.n35 49.9374
R1246 VN.n13 VN.n2 29.8095
R1247 VN.n31 VN.n20 29.8095
R1248 VN.n7 VN.n4 24.4675
R1249 VN.n8 VN.n7 24.4675
R1250 VN.n9 VN.n8 24.4675
R1251 VN.n14 VN.n13 24.4675
R1252 VN.n15 VN.n14 24.4675
R1253 VN.n27 VN.n26 24.4675
R1254 VN.n26 VN.n25 24.4675
R1255 VN.n25 VN.n22 24.4675
R1256 VN.n33 VN.n32 24.4675
R1257 VN.n32 VN.n31 24.4675
R1258 VN.n15 VN.n0 13.702
R1259 VN.n33 VN.n18 13.702
R1260 VN.n24 VN.n23 3.02692
R1261 VN.n6 VN.n5 3.02692
R1262 VN.n35 VN.n34 0.354971
R1263 VN.n17 VN.n16 0.354971
R1264 VN VN.n17 0.26696
R1265 VN.n34 VN.n19 0.189894
R1266 VN.n30 VN.n19 0.189894
R1267 VN.n30 VN.n29 0.189894
R1268 VN.n29 VN.n28 0.189894
R1269 VN.n28 VN.n21 0.189894
R1270 VN.n24 VN.n21 0.189894
R1271 VN.n6 VN.n3 0.189894
R1272 VN.n10 VN.n3 0.189894
R1273 VN.n11 VN.n10 0.189894
R1274 VN.n12 VN.n11 0.189894
R1275 VN.n12 VN.n1 0.189894
R1276 VN.n16 VN.n1 0.189894
R1277 VDD2.n1 VDD2.t0 85.2645
R1278 VDD2.n2 VDD2.t4 82.8762
R1279 VDD2.n1 VDD2.n0 79.9706
R1280 VDD2 VDD2.n3 79.9679
R1281 VDD2.n2 VDD2.n1 41.9524
R1282 VDD2.n3 VDD2.t5 3.6651
R1283 VDD2.n3 VDD2.t2 3.6651
R1284 VDD2.n0 VDD2.t3 3.6651
R1285 VDD2.n0 VDD2.t1 3.6651
R1286 VDD2 VDD2.n2 2.50266
C0 VTAIL VN 5.82545f
C1 w_n3994_n2742# VTAIL 2.62377f
C2 VDD2 VN 5.31473f
C3 VN VP 7.17239f
C4 VDD2 w_n3994_n2742# 2.39534f
C5 w_n3994_n2742# VP 8.22908f
C6 VDD2 VTAIL 7.0304f
C7 VTAIL VP 5.83965f
C8 VDD1 VN 0.151889f
C9 VN B 1.30981f
C10 VDD2 VP 0.530189f
C11 VDD1 w_n3994_n2742# 2.2831f
C12 w_n3994_n2742# B 9.9725f
C13 VDD1 VTAIL 6.972589f
C14 VTAIL B 3.27977f
C15 VDD2 VDD1 1.73823f
C16 VDD2 B 2.15753f
C17 VDD1 VP 5.6904f
C18 VP B 2.18018f
C19 VDD1 B 2.06305f
C20 w_n3994_n2742# VN 7.71034f
C21 VDD2 VSUBS 2.056026f
C22 VDD1 VSUBS 2.60612f
C23 VTAIL VSUBS 1.248365f
C24 VN VSUBS 6.61431f
C25 VP VSUBS 3.492917f
C26 B VSUBS 5.214114f
C27 w_n3994_n2742# VSUBS 0.135588p
C28 VDD2.t0 VSUBS 2.02896f
C29 VDD2.t3 VSUBS 0.206864f
C30 VDD2.t1 VSUBS 0.206864f
C31 VDD2.n0 VSUBS 1.53309f
C32 VDD2.n1 VSUBS 4.18876f
C33 VDD2.t4 VSUBS 2.00539f
C34 VDD2.n2 VSUBS 3.5693f
C35 VDD2.t5 VSUBS 0.206864f
C36 VDD2.t2 VSUBS 0.206864f
C37 VDD2.n3 VSUBS 1.53305f
C38 VN.t4 VSUBS 2.39803f
C39 VN.n0 VSUBS 0.974498f
C40 VN.n1 VSUBS 0.029054f
C41 VN.n2 VSUBS 0.02834f
C42 VN.n3 VSUBS 0.029054f
C43 VN.t2 VSUBS 2.39803f
C44 VN.n4 VSUBS 0.972675f
C45 VN.t5 VSUBS 2.77933f
C46 VN.n5 VSUBS 0.909513f
C47 VN.n6 VSUBS 0.354846f
C48 VN.n7 VSUBS 0.054149f
C49 VN.n8 VSUBS 0.054149f
C50 VN.n9 VSUBS 0.052752f
C51 VN.n10 VSUBS 0.029054f
C52 VN.n11 VSUBS 0.029054f
C53 VN.n12 VSUBS 0.029054f
C54 VN.n13 VSUBS 0.057885f
C55 VN.n14 VSUBS 0.054149f
C56 VN.n15 VSUBS 0.042387f
C57 VN.n16 VSUBS 0.046893f
C58 VN.n17 VSUBS 0.073279f
C59 VN.t1 VSUBS 2.39803f
C60 VN.n18 VSUBS 0.974498f
C61 VN.n19 VSUBS 0.029054f
C62 VN.n20 VSUBS 0.02834f
C63 VN.n21 VSUBS 0.029054f
C64 VN.t0 VSUBS 2.39803f
C65 VN.n22 VSUBS 0.972675f
C66 VN.t3 VSUBS 2.77933f
C67 VN.n23 VSUBS 0.909513f
C68 VN.n24 VSUBS 0.354846f
C69 VN.n25 VSUBS 0.054149f
C70 VN.n26 VSUBS 0.054149f
C71 VN.n27 VSUBS 0.052752f
C72 VN.n28 VSUBS 0.029054f
C73 VN.n29 VSUBS 0.029054f
C74 VN.n30 VSUBS 0.029054f
C75 VN.n31 VSUBS 0.057885f
C76 VN.n32 VSUBS 0.054149f
C77 VN.n33 VSUBS 0.042387f
C78 VN.n34 VSUBS 0.046893f
C79 VN.n35 VSUBS 1.65809f
C80 VTAIL.t1 VSUBS 0.220237f
C81 VTAIL.t4 VSUBS 0.220237f
C82 VTAIL.n0 VSUBS 1.47717f
C83 VTAIL.n1 VSUBS 0.956556f
C84 VTAIL.t10 VSUBS 1.97499f
C85 VTAIL.n2 VSUBS 1.30094f
C86 VTAIL.t7 VSUBS 0.220237f
C87 VTAIL.t9 VSUBS 0.220237f
C88 VTAIL.n3 VSUBS 1.47717f
C89 VTAIL.n4 VSUBS 2.84639f
C90 VTAIL.t0 VSUBS 0.220237f
C91 VTAIL.t5 VSUBS 0.220237f
C92 VTAIL.n5 VSUBS 1.47718f
C93 VTAIL.n6 VSUBS 2.84638f
C94 VTAIL.t3 VSUBS 1.97499f
C95 VTAIL.n7 VSUBS 1.30093f
C96 VTAIL.t8 VSUBS 0.220237f
C97 VTAIL.t11 VSUBS 0.220237f
C98 VTAIL.n8 VSUBS 1.47718f
C99 VTAIL.n9 VSUBS 1.1981f
C100 VTAIL.t6 VSUBS 1.97499f
C101 VTAIL.n10 VSUBS 2.6193f
C102 VTAIL.t2 VSUBS 1.97499f
C103 VTAIL.n11 VSUBS 2.53093f
C104 VDD1.t3 VSUBS 2.04122f
C105 VDD1.t4 VSUBS 2.03982f
C106 VDD1.t2 VSUBS 0.207971f
C107 VDD1.t1 VSUBS 0.207971f
C108 VDD1.n0 VSUBS 1.5413f
C109 VDD1.n1 VSUBS 4.38161f
C110 VDD1.t0 VSUBS 0.207971f
C111 VDD1.t5 VSUBS 0.207971f
C112 VDD1.n2 VSUBS 1.53257f
C113 VDD1.n3 VSUBS 3.58855f
C114 VP.t1 VSUBS 2.68817f
C115 VP.n0 VSUBS 1.0924f
C116 VP.n1 VSUBS 0.032569f
C117 VP.n2 VSUBS 0.031769f
C118 VP.n3 VSUBS 0.032569f
C119 VP.t2 VSUBS 2.68817f
C120 VP.n4 VSUBS 0.991747f
C121 VP.n5 VSUBS 0.032569f
C122 VP.n6 VSUBS 0.031769f
C123 VP.n7 VSUBS 0.032569f
C124 VP.t4 VSUBS 2.68817f
C125 VP.n8 VSUBS 1.0924f
C126 VP.t5 VSUBS 2.68817f
C127 VP.n9 VSUBS 1.0924f
C128 VP.n10 VSUBS 0.032569f
C129 VP.n11 VSUBS 0.031769f
C130 VP.n12 VSUBS 0.032569f
C131 VP.t0 VSUBS 2.68817f
C132 VP.n13 VSUBS 1.09036f
C133 VP.t3 VSUBS 3.11561f
C134 VP.n14 VSUBS 1.01956f
C135 VP.n15 VSUBS 0.39778f
C136 VP.n16 VSUBS 0.060701f
C137 VP.n17 VSUBS 0.060701f
C138 VP.n18 VSUBS 0.059134f
C139 VP.n19 VSUBS 0.032569f
C140 VP.n20 VSUBS 0.032569f
C141 VP.n21 VSUBS 0.032569f
C142 VP.n22 VSUBS 0.064888f
C143 VP.n23 VSUBS 0.060701f
C144 VP.n24 VSUBS 0.047515f
C145 VP.n25 VSUBS 0.052566f
C146 VP.n26 VSUBS 1.84536f
C147 VP.n27 VSUBS 1.86889f
C148 VP.n28 VSUBS 0.052566f
C149 VP.n29 VSUBS 0.047515f
C150 VP.n30 VSUBS 0.060701f
C151 VP.n31 VSUBS 0.064888f
C152 VP.n32 VSUBS 0.032569f
C153 VP.n33 VSUBS 0.032569f
C154 VP.n34 VSUBS 0.032569f
C155 VP.n35 VSUBS 0.059134f
C156 VP.n36 VSUBS 0.060701f
C157 VP.n37 VSUBS 0.060701f
C158 VP.n38 VSUBS 0.032569f
C159 VP.n39 VSUBS 0.032569f
C160 VP.n40 VSUBS 0.032569f
C161 VP.n41 VSUBS 0.060701f
C162 VP.n42 VSUBS 0.060701f
C163 VP.n43 VSUBS 0.059134f
C164 VP.n44 VSUBS 0.032569f
C165 VP.n45 VSUBS 0.032569f
C166 VP.n46 VSUBS 0.032569f
C167 VP.n47 VSUBS 0.064888f
C168 VP.n48 VSUBS 0.060701f
C169 VP.n49 VSUBS 0.047515f
C170 VP.n50 VSUBS 0.052566f
C171 VP.n51 VSUBS 0.082145f
C172 B.n0 VSUBS 0.008524f
C173 B.n1 VSUBS 0.008524f
C174 B.n2 VSUBS 0.012606f
C175 B.n3 VSUBS 0.00966f
C176 B.n4 VSUBS 0.00966f
C177 B.n5 VSUBS 0.00966f
C178 B.n6 VSUBS 0.00966f
C179 B.n7 VSUBS 0.00966f
C180 B.n8 VSUBS 0.00966f
C181 B.n9 VSUBS 0.00966f
C182 B.n10 VSUBS 0.00966f
C183 B.n11 VSUBS 0.00966f
C184 B.n12 VSUBS 0.00966f
C185 B.n13 VSUBS 0.00966f
C186 B.n14 VSUBS 0.00966f
C187 B.n15 VSUBS 0.00966f
C188 B.n16 VSUBS 0.00966f
C189 B.n17 VSUBS 0.00966f
C190 B.n18 VSUBS 0.00966f
C191 B.n19 VSUBS 0.00966f
C192 B.n20 VSUBS 0.00966f
C193 B.n21 VSUBS 0.00966f
C194 B.n22 VSUBS 0.00966f
C195 B.n23 VSUBS 0.00966f
C196 B.n24 VSUBS 0.00966f
C197 B.n25 VSUBS 0.00966f
C198 B.n26 VSUBS 0.00966f
C199 B.n27 VSUBS 0.00966f
C200 B.n28 VSUBS 0.024264f
C201 B.n29 VSUBS 0.00966f
C202 B.n30 VSUBS 0.00966f
C203 B.n31 VSUBS 0.00966f
C204 B.n32 VSUBS 0.00966f
C205 B.n33 VSUBS 0.00966f
C206 B.n34 VSUBS 0.00966f
C207 B.n35 VSUBS 0.00966f
C208 B.n36 VSUBS 0.00966f
C209 B.n37 VSUBS 0.00966f
C210 B.n38 VSUBS 0.00966f
C211 B.n39 VSUBS 0.00966f
C212 B.n40 VSUBS 0.00966f
C213 B.n41 VSUBS 0.00966f
C214 B.n42 VSUBS 0.00966f
C215 B.n43 VSUBS 0.00966f
C216 B.t1 VSUBS 0.383921f
C217 B.t2 VSUBS 0.420063f
C218 B.t0 VSUBS 1.98907f
C219 B.n44 VSUBS 0.235903f
C220 B.n45 VSUBS 0.10352f
C221 B.n46 VSUBS 0.022381f
C222 B.n47 VSUBS 0.00966f
C223 B.n48 VSUBS 0.00966f
C224 B.n49 VSUBS 0.00966f
C225 B.n50 VSUBS 0.00966f
C226 B.n51 VSUBS 0.00966f
C227 B.t4 VSUBS 0.383917f
C228 B.t5 VSUBS 0.420059f
C229 B.t3 VSUBS 1.98907f
C230 B.n52 VSUBS 0.235907f
C231 B.n53 VSUBS 0.103524f
C232 B.n54 VSUBS 0.00966f
C233 B.n55 VSUBS 0.00966f
C234 B.n56 VSUBS 0.00966f
C235 B.n57 VSUBS 0.00966f
C236 B.n58 VSUBS 0.00966f
C237 B.n59 VSUBS 0.00966f
C238 B.n60 VSUBS 0.00966f
C239 B.n61 VSUBS 0.00966f
C240 B.n62 VSUBS 0.00966f
C241 B.n63 VSUBS 0.00966f
C242 B.n64 VSUBS 0.00966f
C243 B.n65 VSUBS 0.00966f
C244 B.n66 VSUBS 0.00966f
C245 B.n67 VSUBS 0.00966f
C246 B.n68 VSUBS 0.00966f
C247 B.n69 VSUBS 0.024264f
C248 B.n70 VSUBS 0.00966f
C249 B.n71 VSUBS 0.00966f
C250 B.n72 VSUBS 0.00966f
C251 B.n73 VSUBS 0.00966f
C252 B.n74 VSUBS 0.00966f
C253 B.n75 VSUBS 0.00966f
C254 B.n76 VSUBS 0.00966f
C255 B.n77 VSUBS 0.00966f
C256 B.n78 VSUBS 0.00966f
C257 B.n79 VSUBS 0.00966f
C258 B.n80 VSUBS 0.00966f
C259 B.n81 VSUBS 0.00966f
C260 B.n82 VSUBS 0.00966f
C261 B.n83 VSUBS 0.00966f
C262 B.n84 VSUBS 0.00966f
C263 B.n85 VSUBS 0.00966f
C264 B.n86 VSUBS 0.00966f
C265 B.n87 VSUBS 0.00966f
C266 B.n88 VSUBS 0.00966f
C267 B.n89 VSUBS 0.00966f
C268 B.n90 VSUBS 0.00966f
C269 B.n91 VSUBS 0.00966f
C270 B.n92 VSUBS 0.00966f
C271 B.n93 VSUBS 0.00966f
C272 B.n94 VSUBS 0.00966f
C273 B.n95 VSUBS 0.00966f
C274 B.n96 VSUBS 0.00966f
C275 B.n97 VSUBS 0.00966f
C276 B.n98 VSUBS 0.00966f
C277 B.n99 VSUBS 0.00966f
C278 B.n100 VSUBS 0.00966f
C279 B.n101 VSUBS 0.00966f
C280 B.n102 VSUBS 0.00966f
C281 B.n103 VSUBS 0.00966f
C282 B.n104 VSUBS 0.00966f
C283 B.n105 VSUBS 0.00966f
C284 B.n106 VSUBS 0.00966f
C285 B.n107 VSUBS 0.00966f
C286 B.n108 VSUBS 0.00966f
C287 B.n109 VSUBS 0.00966f
C288 B.n110 VSUBS 0.00966f
C289 B.n111 VSUBS 0.00966f
C290 B.n112 VSUBS 0.00966f
C291 B.n113 VSUBS 0.00966f
C292 B.n114 VSUBS 0.00966f
C293 B.n115 VSUBS 0.00966f
C294 B.n116 VSUBS 0.00966f
C295 B.n117 VSUBS 0.00966f
C296 B.n118 VSUBS 0.00966f
C297 B.n119 VSUBS 0.00966f
C298 B.n120 VSUBS 0.00966f
C299 B.n121 VSUBS 0.00966f
C300 B.n122 VSUBS 0.02452f
C301 B.n123 VSUBS 0.00966f
C302 B.n124 VSUBS 0.00966f
C303 B.n125 VSUBS 0.00966f
C304 B.n126 VSUBS 0.00966f
C305 B.n127 VSUBS 0.00966f
C306 B.n128 VSUBS 0.00966f
C307 B.n129 VSUBS 0.00966f
C308 B.n130 VSUBS 0.00966f
C309 B.n131 VSUBS 0.00966f
C310 B.n132 VSUBS 0.00966f
C311 B.n133 VSUBS 0.00966f
C312 B.n134 VSUBS 0.00966f
C313 B.n135 VSUBS 0.00966f
C314 B.n136 VSUBS 0.00966f
C315 B.n137 VSUBS 0.00966f
C316 B.n138 VSUBS 0.009092f
C317 B.n139 VSUBS 0.00966f
C318 B.n140 VSUBS 0.00966f
C319 B.n141 VSUBS 0.00966f
C320 B.n142 VSUBS 0.00966f
C321 B.n143 VSUBS 0.00966f
C322 B.t11 VSUBS 0.383921f
C323 B.t10 VSUBS 0.420063f
C324 B.t9 VSUBS 1.98907f
C325 B.n144 VSUBS 0.235903f
C326 B.n145 VSUBS 0.10352f
C327 B.n146 VSUBS 0.00966f
C328 B.n147 VSUBS 0.00966f
C329 B.n148 VSUBS 0.00966f
C330 B.n149 VSUBS 0.00966f
C331 B.n150 VSUBS 0.00966f
C332 B.n151 VSUBS 0.00966f
C333 B.n152 VSUBS 0.00966f
C334 B.n153 VSUBS 0.00966f
C335 B.n154 VSUBS 0.00966f
C336 B.n155 VSUBS 0.00966f
C337 B.n156 VSUBS 0.00966f
C338 B.n157 VSUBS 0.00966f
C339 B.n158 VSUBS 0.00966f
C340 B.n159 VSUBS 0.00966f
C341 B.n160 VSUBS 0.00966f
C342 B.n161 VSUBS 0.024264f
C343 B.n162 VSUBS 0.00966f
C344 B.n163 VSUBS 0.00966f
C345 B.n164 VSUBS 0.00966f
C346 B.n165 VSUBS 0.00966f
C347 B.n166 VSUBS 0.00966f
C348 B.n167 VSUBS 0.00966f
C349 B.n168 VSUBS 0.00966f
C350 B.n169 VSUBS 0.00966f
C351 B.n170 VSUBS 0.00966f
C352 B.n171 VSUBS 0.00966f
C353 B.n172 VSUBS 0.00966f
C354 B.n173 VSUBS 0.00966f
C355 B.n174 VSUBS 0.00966f
C356 B.n175 VSUBS 0.00966f
C357 B.n176 VSUBS 0.00966f
C358 B.n177 VSUBS 0.00966f
C359 B.n178 VSUBS 0.00966f
C360 B.n179 VSUBS 0.00966f
C361 B.n180 VSUBS 0.00966f
C362 B.n181 VSUBS 0.00966f
C363 B.n182 VSUBS 0.00966f
C364 B.n183 VSUBS 0.00966f
C365 B.n184 VSUBS 0.00966f
C366 B.n185 VSUBS 0.00966f
C367 B.n186 VSUBS 0.00966f
C368 B.n187 VSUBS 0.00966f
C369 B.n188 VSUBS 0.00966f
C370 B.n189 VSUBS 0.00966f
C371 B.n190 VSUBS 0.00966f
C372 B.n191 VSUBS 0.00966f
C373 B.n192 VSUBS 0.00966f
C374 B.n193 VSUBS 0.00966f
C375 B.n194 VSUBS 0.00966f
C376 B.n195 VSUBS 0.00966f
C377 B.n196 VSUBS 0.00966f
C378 B.n197 VSUBS 0.00966f
C379 B.n198 VSUBS 0.00966f
C380 B.n199 VSUBS 0.00966f
C381 B.n200 VSUBS 0.00966f
C382 B.n201 VSUBS 0.00966f
C383 B.n202 VSUBS 0.00966f
C384 B.n203 VSUBS 0.00966f
C385 B.n204 VSUBS 0.00966f
C386 B.n205 VSUBS 0.00966f
C387 B.n206 VSUBS 0.00966f
C388 B.n207 VSUBS 0.00966f
C389 B.n208 VSUBS 0.00966f
C390 B.n209 VSUBS 0.00966f
C391 B.n210 VSUBS 0.00966f
C392 B.n211 VSUBS 0.00966f
C393 B.n212 VSUBS 0.00966f
C394 B.n213 VSUBS 0.00966f
C395 B.n214 VSUBS 0.00966f
C396 B.n215 VSUBS 0.00966f
C397 B.n216 VSUBS 0.00966f
C398 B.n217 VSUBS 0.00966f
C399 B.n218 VSUBS 0.00966f
C400 B.n219 VSUBS 0.00966f
C401 B.n220 VSUBS 0.00966f
C402 B.n221 VSUBS 0.00966f
C403 B.n222 VSUBS 0.00966f
C404 B.n223 VSUBS 0.00966f
C405 B.n224 VSUBS 0.00966f
C406 B.n225 VSUBS 0.00966f
C407 B.n226 VSUBS 0.00966f
C408 B.n227 VSUBS 0.00966f
C409 B.n228 VSUBS 0.00966f
C410 B.n229 VSUBS 0.00966f
C411 B.n230 VSUBS 0.00966f
C412 B.n231 VSUBS 0.00966f
C413 B.n232 VSUBS 0.00966f
C414 B.n233 VSUBS 0.00966f
C415 B.n234 VSUBS 0.00966f
C416 B.n235 VSUBS 0.00966f
C417 B.n236 VSUBS 0.00966f
C418 B.n237 VSUBS 0.00966f
C419 B.n238 VSUBS 0.00966f
C420 B.n239 VSUBS 0.00966f
C421 B.n240 VSUBS 0.00966f
C422 B.n241 VSUBS 0.00966f
C423 B.n242 VSUBS 0.00966f
C424 B.n243 VSUBS 0.00966f
C425 B.n244 VSUBS 0.00966f
C426 B.n245 VSUBS 0.00966f
C427 B.n246 VSUBS 0.00966f
C428 B.n247 VSUBS 0.00966f
C429 B.n248 VSUBS 0.00966f
C430 B.n249 VSUBS 0.00966f
C431 B.n250 VSUBS 0.00966f
C432 B.n251 VSUBS 0.00966f
C433 B.n252 VSUBS 0.00966f
C434 B.n253 VSUBS 0.00966f
C435 B.n254 VSUBS 0.00966f
C436 B.n255 VSUBS 0.00966f
C437 B.n256 VSUBS 0.00966f
C438 B.n257 VSUBS 0.00966f
C439 B.n258 VSUBS 0.00966f
C440 B.n259 VSUBS 0.00966f
C441 B.n260 VSUBS 0.00966f
C442 B.n261 VSUBS 0.00966f
C443 B.n262 VSUBS 0.023468f
C444 B.n263 VSUBS 0.023468f
C445 B.n264 VSUBS 0.024264f
C446 B.n265 VSUBS 0.00966f
C447 B.n266 VSUBS 0.00966f
C448 B.n267 VSUBS 0.00966f
C449 B.n268 VSUBS 0.00966f
C450 B.n269 VSUBS 0.00966f
C451 B.n270 VSUBS 0.00966f
C452 B.n271 VSUBS 0.00966f
C453 B.n272 VSUBS 0.00966f
C454 B.n273 VSUBS 0.00966f
C455 B.n274 VSUBS 0.00966f
C456 B.n275 VSUBS 0.00966f
C457 B.n276 VSUBS 0.00966f
C458 B.n277 VSUBS 0.00966f
C459 B.n278 VSUBS 0.00966f
C460 B.n279 VSUBS 0.00966f
C461 B.n280 VSUBS 0.00966f
C462 B.n281 VSUBS 0.00966f
C463 B.n282 VSUBS 0.00966f
C464 B.n283 VSUBS 0.00966f
C465 B.n284 VSUBS 0.00966f
C466 B.n285 VSUBS 0.00966f
C467 B.n286 VSUBS 0.00966f
C468 B.n287 VSUBS 0.00966f
C469 B.n288 VSUBS 0.00966f
C470 B.n289 VSUBS 0.00966f
C471 B.n290 VSUBS 0.00966f
C472 B.n291 VSUBS 0.00966f
C473 B.n292 VSUBS 0.00966f
C474 B.n293 VSUBS 0.00966f
C475 B.n294 VSUBS 0.00966f
C476 B.n295 VSUBS 0.00966f
C477 B.n296 VSUBS 0.00966f
C478 B.n297 VSUBS 0.00966f
C479 B.n298 VSUBS 0.00966f
C480 B.n299 VSUBS 0.00966f
C481 B.n300 VSUBS 0.00966f
C482 B.n301 VSUBS 0.00966f
C483 B.n302 VSUBS 0.00966f
C484 B.n303 VSUBS 0.00966f
C485 B.n304 VSUBS 0.00966f
C486 B.n305 VSUBS 0.00966f
C487 B.n306 VSUBS 0.00966f
C488 B.n307 VSUBS 0.00966f
C489 B.n308 VSUBS 0.00966f
C490 B.n309 VSUBS 0.00966f
C491 B.n310 VSUBS 0.00966f
C492 B.n311 VSUBS 0.009092f
C493 B.n312 VSUBS 0.022381f
C494 B.n313 VSUBS 0.005398f
C495 B.n314 VSUBS 0.00966f
C496 B.n315 VSUBS 0.00966f
C497 B.n316 VSUBS 0.00966f
C498 B.n317 VSUBS 0.00966f
C499 B.n318 VSUBS 0.00966f
C500 B.n319 VSUBS 0.00966f
C501 B.n320 VSUBS 0.00966f
C502 B.n321 VSUBS 0.00966f
C503 B.n322 VSUBS 0.00966f
C504 B.n323 VSUBS 0.00966f
C505 B.n324 VSUBS 0.00966f
C506 B.n325 VSUBS 0.00966f
C507 B.t8 VSUBS 0.383917f
C508 B.t7 VSUBS 0.420059f
C509 B.t6 VSUBS 1.98907f
C510 B.n326 VSUBS 0.235907f
C511 B.n327 VSUBS 0.103524f
C512 B.n328 VSUBS 0.022381f
C513 B.n329 VSUBS 0.005398f
C514 B.n330 VSUBS 0.00966f
C515 B.n331 VSUBS 0.00966f
C516 B.n332 VSUBS 0.00966f
C517 B.n333 VSUBS 0.00966f
C518 B.n334 VSUBS 0.00966f
C519 B.n335 VSUBS 0.00966f
C520 B.n336 VSUBS 0.00966f
C521 B.n337 VSUBS 0.00966f
C522 B.n338 VSUBS 0.00966f
C523 B.n339 VSUBS 0.00966f
C524 B.n340 VSUBS 0.00966f
C525 B.n341 VSUBS 0.00966f
C526 B.n342 VSUBS 0.00966f
C527 B.n343 VSUBS 0.00966f
C528 B.n344 VSUBS 0.00966f
C529 B.n345 VSUBS 0.00966f
C530 B.n346 VSUBS 0.00966f
C531 B.n347 VSUBS 0.00966f
C532 B.n348 VSUBS 0.00966f
C533 B.n349 VSUBS 0.00966f
C534 B.n350 VSUBS 0.00966f
C535 B.n351 VSUBS 0.00966f
C536 B.n352 VSUBS 0.00966f
C537 B.n353 VSUBS 0.00966f
C538 B.n354 VSUBS 0.00966f
C539 B.n355 VSUBS 0.00966f
C540 B.n356 VSUBS 0.00966f
C541 B.n357 VSUBS 0.00966f
C542 B.n358 VSUBS 0.00966f
C543 B.n359 VSUBS 0.00966f
C544 B.n360 VSUBS 0.00966f
C545 B.n361 VSUBS 0.00966f
C546 B.n362 VSUBS 0.00966f
C547 B.n363 VSUBS 0.00966f
C548 B.n364 VSUBS 0.00966f
C549 B.n365 VSUBS 0.00966f
C550 B.n366 VSUBS 0.00966f
C551 B.n367 VSUBS 0.00966f
C552 B.n368 VSUBS 0.00966f
C553 B.n369 VSUBS 0.00966f
C554 B.n370 VSUBS 0.00966f
C555 B.n371 VSUBS 0.00966f
C556 B.n372 VSUBS 0.00966f
C557 B.n373 VSUBS 0.00966f
C558 B.n374 VSUBS 0.00966f
C559 B.n375 VSUBS 0.00966f
C560 B.n376 VSUBS 0.00966f
C561 B.n377 VSUBS 0.023212f
C562 B.n378 VSUBS 0.024264f
C563 B.n379 VSUBS 0.023468f
C564 B.n380 VSUBS 0.00966f
C565 B.n381 VSUBS 0.00966f
C566 B.n382 VSUBS 0.00966f
C567 B.n383 VSUBS 0.00966f
C568 B.n384 VSUBS 0.00966f
C569 B.n385 VSUBS 0.00966f
C570 B.n386 VSUBS 0.00966f
C571 B.n387 VSUBS 0.00966f
C572 B.n388 VSUBS 0.00966f
C573 B.n389 VSUBS 0.00966f
C574 B.n390 VSUBS 0.00966f
C575 B.n391 VSUBS 0.00966f
C576 B.n392 VSUBS 0.00966f
C577 B.n393 VSUBS 0.00966f
C578 B.n394 VSUBS 0.00966f
C579 B.n395 VSUBS 0.00966f
C580 B.n396 VSUBS 0.00966f
C581 B.n397 VSUBS 0.00966f
C582 B.n398 VSUBS 0.00966f
C583 B.n399 VSUBS 0.00966f
C584 B.n400 VSUBS 0.00966f
C585 B.n401 VSUBS 0.00966f
C586 B.n402 VSUBS 0.00966f
C587 B.n403 VSUBS 0.00966f
C588 B.n404 VSUBS 0.00966f
C589 B.n405 VSUBS 0.00966f
C590 B.n406 VSUBS 0.00966f
C591 B.n407 VSUBS 0.00966f
C592 B.n408 VSUBS 0.00966f
C593 B.n409 VSUBS 0.00966f
C594 B.n410 VSUBS 0.00966f
C595 B.n411 VSUBS 0.00966f
C596 B.n412 VSUBS 0.00966f
C597 B.n413 VSUBS 0.00966f
C598 B.n414 VSUBS 0.00966f
C599 B.n415 VSUBS 0.00966f
C600 B.n416 VSUBS 0.00966f
C601 B.n417 VSUBS 0.00966f
C602 B.n418 VSUBS 0.00966f
C603 B.n419 VSUBS 0.00966f
C604 B.n420 VSUBS 0.00966f
C605 B.n421 VSUBS 0.00966f
C606 B.n422 VSUBS 0.00966f
C607 B.n423 VSUBS 0.00966f
C608 B.n424 VSUBS 0.00966f
C609 B.n425 VSUBS 0.00966f
C610 B.n426 VSUBS 0.00966f
C611 B.n427 VSUBS 0.00966f
C612 B.n428 VSUBS 0.00966f
C613 B.n429 VSUBS 0.00966f
C614 B.n430 VSUBS 0.00966f
C615 B.n431 VSUBS 0.00966f
C616 B.n432 VSUBS 0.00966f
C617 B.n433 VSUBS 0.00966f
C618 B.n434 VSUBS 0.00966f
C619 B.n435 VSUBS 0.00966f
C620 B.n436 VSUBS 0.00966f
C621 B.n437 VSUBS 0.00966f
C622 B.n438 VSUBS 0.00966f
C623 B.n439 VSUBS 0.00966f
C624 B.n440 VSUBS 0.00966f
C625 B.n441 VSUBS 0.00966f
C626 B.n442 VSUBS 0.00966f
C627 B.n443 VSUBS 0.00966f
C628 B.n444 VSUBS 0.00966f
C629 B.n445 VSUBS 0.00966f
C630 B.n446 VSUBS 0.00966f
C631 B.n447 VSUBS 0.00966f
C632 B.n448 VSUBS 0.00966f
C633 B.n449 VSUBS 0.00966f
C634 B.n450 VSUBS 0.00966f
C635 B.n451 VSUBS 0.00966f
C636 B.n452 VSUBS 0.00966f
C637 B.n453 VSUBS 0.00966f
C638 B.n454 VSUBS 0.00966f
C639 B.n455 VSUBS 0.00966f
C640 B.n456 VSUBS 0.00966f
C641 B.n457 VSUBS 0.00966f
C642 B.n458 VSUBS 0.00966f
C643 B.n459 VSUBS 0.00966f
C644 B.n460 VSUBS 0.00966f
C645 B.n461 VSUBS 0.00966f
C646 B.n462 VSUBS 0.00966f
C647 B.n463 VSUBS 0.00966f
C648 B.n464 VSUBS 0.00966f
C649 B.n465 VSUBS 0.00966f
C650 B.n466 VSUBS 0.00966f
C651 B.n467 VSUBS 0.00966f
C652 B.n468 VSUBS 0.00966f
C653 B.n469 VSUBS 0.00966f
C654 B.n470 VSUBS 0.00966f
C655 B.n471 VSUBS 0.00966f
C656 B.n472 VSUBS 0.00966f
C657 B.n473 VSUBS 0.00966f
C658 B.n474 VSUBS 0.00966f
C659 B.n475 VSUBS 0.00966f
C660 B.n476 VSUBS 0.00966f
C661 B.n477 VSUBS 0.00966f
C662 B.n478 VSUBS 0.00966f
C663 B.n479 VSUBS 0.00966f
C664 B.n480 VSUBS 0.00966f
C665 B.n481 VSUBS 0.00966f
C666 B.n482 VSUBS 0.00966f
C667 B.n483 VSUBS 0.00966f
C668 B.n484 VSUBS 0.00966f
C669 B.n485 VSUBS 0.00966f
C670 B.n486 VSUBS 0.00966f
C671 B.n487 VSUBS 0.00966f
C672 B.n488 VSUBS 0.00966f
C673 B.n489 VSUBS 0.00966f
C674 B.n490 VSUBS 0.00966f
C675 B.n491 VSUBS 0.00966f
C676 B.n492 VSUBS 0.00966f
C677 B.n493 VSUBS 0.00966f
C678 B.n494 VSUBS 0.00966f
C679 B.n495 VSUBS 0.00966f
C680 B.n496 VSUBS 0.00966f
C681 B.n497 VSUBS 0.00966f
C682 B.n498 VSUBS 0.00966f
C683 B.n499 VSUBS 0.00966f
C684 B.n500 VSUBS 0.00966f
C685 B.n501 VSUBS 0.00966f
C686 B.n502 VSUBS 0.00966f
C687 B.n503 VSUBS 0.00966f
C688 B.n504 VSUBS 0.00966f
C689 B.n505 VSUBS 0.00966f
C690 B.n506 VSUBS 0.00966f
C691 B.n507 VSUBS 0.00966f
C692 B.n508 VSUBS 0.00966f
C693 B.n509 VSUBS 0.00966f
C694 B.n510 VSUBS 0.00966f
C695 B.n511 VSUBS 0.00966f
C696 B.n512 VSUBS 0.00966f
C697 B.n513 VSUBS 0.00966f
C698 B.n514 VSUBS 0.00966f
C699 B.n515 VSUBS 0.00966f
C700 B.n516 VSUBS 0.00966f
C701 B.n517 VSUBS 0.00966f
C702 B.n518 VSUBS 0.00966f
C703 B.n519 VSUBS 0.00966f
C704 B.n520 VSUBS 0.00966f
C705 B.n521 VSUBS 0.00966f
C706 B.n522 VSUBS 0.00966f
C707 B.n523 VSUBS 0.00966f
C708 B.n524 VSUBS 0.00966f
C709 B.n525 VSUBS 0.00966f
C710 B.n526 VSUBS 0.00966f
C711 B.n527 VSUBS 0.00966f
C712 B.n528 VSUBS 0.00966f
C713 B.n529 VSUBS 0.00966f
C714 B.n530 VSUBS 0.00966f
C715 B.n531 VSUBS 0.00966f
C716 B.n532 VSUBS 0.00966f
C717 B.n533 VSUBS 0.00966f
C718 B.n534 VSUBS 0.00966f
C719 B.n535 VSUBS 0.00966f
C720 B.n536 VSUBS 0.023468f
C721 B.n537 VSUBS 0.023468f
C722 B.n538 VSUBS 0.024264f
C723 B.n539 VSUBS 0.00966f
C724 B.n540 VSUBS 0.00966f
C725 B.n541 VSUBS 0.00966f
C726 B.n542 VSUBS 0.00966f
C727 B.n543 VSUBS 0.00966f
C728 B.n544 VSUBS 0.00966f
C729 B.n545 VSUBS 0.00966f
C730 B.n546 VSUBS 0.00966f
C731 B.n547 VSUBS 0.00966f
C732 B.n548 VSUBS 0.00966f
C733 B.n549 VSUBS 0.00966f
C734 B.n550 VSUBS 0.00966f
C735 B.n551 VSUBS 0.00966f
C736 B.n552 VSUBS 0.00966f
C737 B.n553 VSUBS 0.00966f
C738 B.n554 VSUBS 0.00966f
C739 B.n555 VSUBS 0.00966f
C740 B.n556 VSUBS 0.00966f
C741 B.n557 VSUBS 0.00966f
C742 B.n558 VSUBS 0.00966f
C743 B.n559 VSUBS 0.00966f
C744 B.n560 VSUBS 0.00966f
C745 B.n561 VSUBS 0.00966f
C746 B.n562 VSUBS 0.00966f
C747 B.n563 VSUBS 0.00966f
C748 B.n564 VSUBS 0.00966f
C749 B.n565 VSUBS 0.00966f
C750 B.n566 VSUBS 0.00966f
C751 B.n567 VSUBS 0.00966f
C752 B.n568 VSUBS 0.00966f
C753 B.n569 VSUBS 0.00966f
C754 B.n570 VSUBS 0.00966f
C755 B.n571 VSUBS 0.00966f
C756 B.n572 VSUBS 0.00966f
C757 B.n573 VSUBS 0.00966f
C758 B.n574 VSUBS 0.00966f
C759 B.n575 VSUBS 0.00966f
C760 B.n576 VSUBS 0.00966f
C761 B.n577 VSUBS 0.00966f
C762 B.n578 VSUBS 0.00966f
C763 B.n579 VSUBS 0.00966f
C764 B.n580 VSUBS 0.00966f
C765 B.n581 VSUBS 0.00966f
C766 B.n582 VSUBS 0.00966f
C767 B.n583 VSUBS 0.00966f
C768 B.n584 VSUBS 0.00966f
C769 B.n585 VSUBS 0.009092f
C770 B.n586 VSUBS 0.022381f
C771 B.n587 VSUBS 0.005398f
C772 B.n588 VSUBS 0.00966f
C773 B.n589 VSUBS 0.00966f
C774 B.n590 VSUBS 0.00966f
C775 B.n591 VSUBS 0.00966f
C776 B.n592 VSUBS 0.00966f
C777 B.n593 VSUBS 0.00966f
C778 B.n594 VSUBS 0.00966f
C779 B.n595 VSUBS 0.00966f
C780 B.n596 VSUBS 0.00966f
C781 B.n597 VSUBS 0.00966f
C782 B.n598 VSUBS 0.00966f
C783 B.n599 VSUBS 0.00966f
C784 B.n600 VSUBS 0.005398f
C785 B.n601 VSUBS 0.00966f
C786 B.n602 VSUBS 0.00966f
C787 B.n603 VSUBS 0.009092f
C788 B.n604 VSUBS 0.00966f
C789 B.n605 VSUBS 0.00966f
C790 B.n606 VSUBS 0.00966f
C791 B.n607 VSUBS 0.00966f
C792 B.n608 VSUBS 0.00966f
C793 B.n609 VSUBS 0.00966f
C794 B.n610 VSUBS 0.00966f
C795 B.n611 VSUBS 0.00966f
C796 B.n612 VSUBS 0.00966f
C797 B.n613 VSUBS 0.00966f
C798 B.n614 VSUBS 0.00966f
C799 B.n615 VSUBS 0.00966f
C800 B.n616 VSUBS 0.00966f
C801 B.n617 VSUBS 0.00966f
C802 B.n618 VSUBS 0.00966f
C803 B.n619 VSUBS 0.00966f
C804 B.n620 VSUBS 0.00966f
C805 B.n621 VSUBS 0.00966f
C806 B.n622 VSUBS 0.00966f
C807 B.n623 VSUBS 0.00966f
C808 B.n624 VSUBS 0.00966f
C809 B.n625 VSUBS 0.00966f
C810 B.n626 VSUBS 0.00966f
C811 B.n627 VSUBS 0.00966f
C812 B.n628 VSUBS 0.00966f
C813 B.n629 VSUBS 0.00966f
C814 B.n630 VSUBS 0.00966f
C815 B.n631 VSUBS 0.00966f
C816 B.n632 VSUBS 0.00966f
C817 B.n633 VSUBS 0.00966f
C818 B.n634 VSUBS 0.00966f
C819 B.n635 VSUBS 0.00966f
C820 B.n636 VSUBS 0.00966f
C821 B.n637 VSUBS 0.00966f
C822 B.n638 VSUBS 0.00966f
C823 B.n639 VSUBS 0.00966f
C824 B.n640 VSUBS 0.00966f
C825 B.n641 VSUBS 0.00966f
C826 B.n642 VSUBS 0.00966f
C827 B.n643 VSUBS 0.00966f
C828 B.n644 VSUBS 0.00966f
C829 B.n645 VSUBS 0.00966f
C830 B.n646 VSUBS 0.00966f
C831 B.n647 VSUBS 0.00966f
C832 B.n648 VSUBS 0.00966f
C833 B.n649 VSUBS 0.024264f
C834 B.n650 VSUBS 0.023468f
C835 B.n651 VSUBS 0.023468f
C836 B.n652 VSUBS 0.00966f
C837 B.n653 VSUBS 0.00966f
C838 B.n654 VSUBS 0.00966f
C839 B.n655 VSUBS 0.00966f
C840 B.n656 VSUBS 0.00966f
C841 B.n657 VSUBS 0.00966f
C842 B.n658 VSUBS 0.00966f
C843 B.n659 VSUBS 0.00966f
C844 B.n660 VSUBS 0.00966f
C845 B.n661 VSUBS 0.00966f
C846 B.n662 VSUBS 0.00966f
C847 B.n663 VSUBS 0.00966f
C848 B.n664 VSUBS 0.00966f
C849 B.n665 VSUBS 0.00966f
C850 B.n666 VSUBS 0.00966f
C851 B.n667 VSUBS 0.00966f
C852 B.n668 VSUBS 0.00966f
C853 B.n669 VSUBS 0.00966f
C854 B.n670 VSUBS 0.00966f
C855 B.n671 VSUBS 0.00966f
C856 B.n672 VSUBS 0.00966f
C857 B.n673 VSUBS 0.00966f
C858 B.n674 VSUBS 0.00966f
C859 B.n675 VSUBS 0.00966f
C860 B.n676 VSUBS 0.00966f
C861 B.n677 VSUBS 0.00966f
C862 B.n678 VSUBS 0.00966f
C863 B.n679 VSUBS 0.00966f
C864 B.n680 VSUBS 0.00966f
C865 B.n681 VSUBS 0.00966f
C866 B.n682 VSUBS 0.00966f
C867 B.n683 VSUBS 0.00966f
C868 B.n684 VSUBS 0.00966f
C869 B.n685 VSUBS 0.00966f
C870 B.n686 VSUBS 0.00966f
C871 B.n687 VSUBS 0.00966f
C872 B.n688 VSUBS 0.00966f
C873 B.n689 VSUBS 0.00966f
C874 B.n690 VSUBS 0.00966f
C875 B.n691 VSUBS 0.00966f
C876 B.n692 VSUBS 0.00966f
C877 B.n693 VSUBS 0.00966f
C878 B.n694 VSUBS 0.00966f
C879 B.n695 VSUBS 0.00966f
C880 B.n696 VSUBS 0.00966f
C881 B.n697 VSUBS 0.00966f
C882 B.n698 VSUBS 0.00966f
C883 B.n699 VSUBS 0.00966f
C884 B.n700 VSUBS 0.00966f
C885 B.n701 VSUBS 0.00966f
C886 B.n702 VSUBS 0.00966f
C887 B.n703 VSUBS 0.00966f
C888 B.n704 VSUBS 0.00966f
C889 B.n705 VSUBS 0.00966f
C890 B.n706 VSUBS 0.00966f
C891 B.n707 VSUBS 0.00966f
C892 B.n708 VSUBS 0.00966f
C893 B.n709 VSUBS 0.00966f
C894 B.n710 VSUBS 0.00966f
C895 B.n711 VSUBS 0.00966f
C896 B.n712 VSUBS 0.00966f
C897 B.n713 VSUBS 0.00966f
C898 B.n714 VSUBS 0.00966f
C899 B.n715 VSUBS 0.00966f
C900 B.n716 VSUBS 0.00966f
C901 B.n717 VSUBS 0.00966f
C902 B.n718 VSUBS 0.00966f
C903 B.n719 VSUBS 0.00966f
C904 B.n720 VSUBS 0.00966f
C905 B.n721 VSUBS 0.00966f
C906 B.n722 VSUBS 0.00966f
C907 B.n723 VSUBS 0.00966f
C908 B.n724 VSUBS 0.00966f
C909 B.n725 VSUBS 0.00966f
C910 B.n726 VSUBS 0.00966f
C911 B.n727 VSUBS 0.012606f
C912 B.n728 VSUBS 0.013429f
C913 B.n729 VSUBS 0.026704f
.ends

