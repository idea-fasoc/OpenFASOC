* NGSPICE file created from diff_pair_sample_1371.ext - technology: sky130A

.subckt diff_pair_sample_1371 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=1.9041 ps=11.87 w=11.54 l=1.24
X1 B.t11 B.t9 B.t10 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=0 ps=0 w=11.54 l=1.24
X2 B.t8 B.t6 B.t7 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=0 ps=0 w=11.54 l=1.24
X3 VTAIL.t6 VP.t1 VDD1.t1 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=1.9041 ps=11.87 w=11.54 l=1.24
X4 B.t5 B.t3 B.t4 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=0 ps=0 w=11.54 l=1.24
X5 VDD2.t3 VN.t0 VTAIL.t3 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=1.9041 pd=11.87 as=4.5006 ps=23.86 w=11.54 l=1.24
X6 VTAIL.t2 VN.t1 VDD2.t2 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=1.9041 ps=11.87 w=11.54 l=1.24
X7 VDD1.t3 VP.t2 VTAIL.t5 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=1.9041 pd=11.87 as=4.5006 ps=23.86 w=11.54 l=1.24
X8 VDD2.t1 VN.t2 VTAIL.t1 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=1.9041 pd=11.87 as=4.5006 ps=23.86 w=11.54 l=1.24
X9 B.t2 B.t0 B.t1 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=0 ps=0 w=11.54 l=1.24
X10 VDD1.t2 VP.t3 VTAIL.t4 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=1.9041 pd=11.87 as=4.5006 ps=23.86 w=11.54 l=1.24
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n1912_n3276# sky130_fd_pr__pfet_01v8 ad=4.5006 pd=23.86 as=1.9041 ps=11.87 w=11.54 l=1.24
R0 VP.n2 VP.t1 260.993
R1 VP.n2 VP.t3 260.772
R2 VP.n3 VP.t0 224.286
R3 VP.n9 VP.t2 224.286
R4 VP.n4 VP.n3 171.875
R5 VP.n10 VP.n9 171.875
R6 VP.n8 VP.n0 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n5 VP.n1 161.3
R9 VP.n4 VP.n2 59.9579
R10 VP.n7 VP.n1 40.577
R11 VP.n8 VP.n7 40.577
R12 VP.n3 VP.n1 14.0178
R13 VP.n9 VP.n8 14.0178
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 115.746
R20 VDD1 VDD1.n0 77.5561
R21 VDD1.n0 VDD1.t1 2.81722
R22 VDD1.n0 VDD1.t2 2.81722
R23 VDD1.n1 VDD1.t0 2.81722
R24 VDD1.n1 VDD1.t3 2.81722
R25 VTAIL.n490 VTAIL.n434 756.745
R26 VTAIL.n56 VTAIL.n0 756.745
R27 VTAIL.n118 VTAIL.n62 756.745
R28 VTAIL.n180 VTAIL.n124 756.745
R29 VTAIL.n428 VTAIL.n372 756.745
R30 VTAIL.n366 VTAIL.n310 756.745
R31 VTAIL.n304 VTAIL.n248 756.745
R32 VTAIL.n242 VTAIL.n186 756.745
R33 VTAIL.n455 VTAIL.n454 585
R34 VTAIL.n457 VTAIL.n456 585
R35 VTAIL.n450 VTAIL.n449 585
R36 VTAIL.n463 VTAIL.n462 585
R37 VTAIL.n465 VTAIL.n464 585
R38 VTAIL.n446 VTAIL.n445 585
R39 VTAIL.n472 VTAIL.n471 585
R40 VTAIL.n473 VTAIL.n444 585
R41 VTAIL.n475 VTAIL.n474 585
R42 VTAIL.n442 VTAIL.n441 585
R43 VTAIL.n481 VTAIL.n480 585
R44 VTAIL.n483 VTAIL.n482 585
R45 VTAIL.n438 VTAIL.n437 585
R46 VTAIL.n489 VTAIL.n488 585
R47 VTAIL.n491 VTAIL.n490 585
R48 VTAIL.n21 VTAIL.n20 585
R49 VTAIL.n23 VTAIL.n22 585
R50 VTAIL.n16 VTAIL.n15 585
R51 VTAIL.n29 VTAIL.n28 585
R52 VTAIL.n31 VTAIL.n30 585
R53 VTAIL.n12 VTAIL.n11 585
R54 VTAIL.n38 VTAIL.n37 585
R55 VTAIL.n39 VTAIL.n10 585
R56 VTAIL.n41 VTAIL.n40 585
R57 VTAIL.n8 VTAIL.n7 585
R58 VTAIL.n47 VTAIL.n46 585
R59 VTAIL.n49 VTAIL.n48 585
R60 VTAIL.n4 VTAIL.n3 585
R61 VTAIL.n55 VTAIL.n54 585
R62 VTAIL.n57 VTAIL.n56 585
R63 VTAIL.n83 VTAIL.n82 585
R64 VTAIL.n85 VTAIL.n84 585
R65 VTAIL.n78 VTAIL.n77 585
R66 VTAIL.n91 VTAIL.n90 585
R67 VTAIL.n93 VTAIL.n92 585
R68 VTAIL.n74 VTAIL.n73 585
R69 VTAIL.n100 VTAIL.n99 585
R70 VTAIL.n101 VTAIL.n72 585
R71 VTAIL.n103 VTAIL.n102 585
R72 VTAIL.n70 VTAIL.n69 585
R73 VTAIL.n109 VTAIL.n108 585
R74 VTAIL.n111 VTAIL.n110 585
R75 VTAIL.n66 VTAIL.n65 585
R76 VTAIL.n117 VTAIL.n116 585
R77 VTAIL.n119 VTAIL.n118 585
R78 VTAIL.n145 VTAIL.n144 585
R79 VTAIL.n147 VTAIL.n146 585
R80 VTAIL.n140 VTAIL.n139 585
R81 VTAIL.n153 VTAIL.n152 585
R82 VTAIL.n155 VTAIL.n154 585
R83 VTAIL.n136 VTAIL.n135 585
R84 VTAIL.n162 VTAIL.n161 585
R85 VTAIL.n163 VTAIL.n134 585
R86 VTAIL.n165 VTAIL.n164 585
R87 VTAIL.n132 VTAIL.n131 585
R88 VTAIL.n171 VTAIL.n170 585
R89 VTAIL.n173 VTAIL.n172 585
R90 VTAIL.n128 VTAIL.n127 585
R91 VTAIL.n179 VTAIL.n178 585
R92 VTAIL.n181 VTAIL.n180 585
R93 VTAIL.n429 VTAIL.n428 585
R94 VTAIL.n427 VTAIL.n426 585
R95 VTAIL.n376 VTAIL.n375 585
R96 VTAIL.n421 VTAIL.n420 585
R97 VTAIL.n419 VTAIL.n418 585
R98 VTAIL.n380 VTAIL.n379 585
R99 VTAIL.n384 VTAIL.n382 585
R100 VTAIL.n413 VTAIL.n412 585
R101 VTAIL.n411 VTAIL.n410 585
R102 VTAIL.n386 VTAIL.n385 585
R103 VTAIL.n405 VTAIL.n404 585
R104 VTAIL.n403 VTAIL.n402 585
R105 VTAIL.n390 VTAIL.n389 585
R106 VTAIL.n397 VTAIL.n396 585
R107 VTAIL.n395 VTAIL.n394 585
R108 VTAIL.n367 VTAIL.n366 585
R109 VTAIL.n365 VTAIL.n364 585
R110 VTAIL.n314 VTAIL.n313 585
R111 VTAIL.n359 VTAIL.n358 585
R112 VTAIL.n357 VTAIL.n356 585
R113 VTAIL.n318 VTAIL.n317 585
R114 VTAIL.n322 VTAIL.n320 585
R115 VTAIL.n351 VTAIL.n350 585
R116 VTAIL.n349 VTAIL.n348 585
R117 VTAIL.n324 VTAIL.n323 585
R118 VTAIL.n343 VTAIL.n342 585
R119 VTAIL.n341 VTAIL.n340 585
R120 VTAIL.n328 VTAIL.n327 585
R121 VTAIL.n335 VTAIL.n334 585
R122 VTAIL.n333 VTAIL.n332 585
R123 VTAIL.n305 VTAIL.n304 585
R124 VTAIL.n303 VTAIL.n302 585
R125 VTAIL.n252 VTAIL.n251 585
R126 VTAIL.n297 VTAIL.n296 585
R127 VTAIL.n295 VTAIL.n294 585
R128 VTAIL.n256 VTAIL.n255 585
R129 VTAIL.n260 VTAIL.n258 585
R130 VTAIL.n289 VTAIL.n288 585
R131 VTAIL.n287 VTAIL.n286 585
R132 VTAIL.n262 VTAIL.n261 585
R133 VTAIL.n281 VTAIL.n280 585
R134 VTAIL.n279 VTAIL.n278 585
R135 VTAIL.n266 VTAIL.n265 585
R136 VTAIL.n273 VTAIL.n272 585
R137 VTAIL.n271 VTAIL.n270 585
R138 VTAIL.n243 VTAIL.n242 585
R139 VTAIL.n241 VTAIL.n240 585
R140 VTAIL.n190 VTAIL.n189 585
R141 VTAIL.n235 VTAIL.n234 585
R142 VTAIL.n233 VTAIL.n232 585
R143 VTAIL.n194 VTAIL.n193 585
R144 VTAIL.n198 VTAIL.n196 585
R145 VTAIL.n227 VTAIL.n226 585
R146 VTAIL.n225 VTAIL.n224 585
R147 VTAIL.n200 VTAIL.n199 585
R148 VTAIL.n219 VTAIL.n218 585
R149 VTAIL.n217 VTAIL.n216 585
R150 VTAIL.n204 VTAIL.n203 585
R151 VTAIL.n211 VTAIL.n210 585
R152 VTAIL.n209 VTAIL.n208 585
R153 VTAIL.n453 VTAIL.t1 329.036
R154 VTAIL.n19 VTAIL.t2 329.036
R155 VTAIL.n81 VTAIL.t5 329.036
R156 VTAIL.n143 VTAIL.t7 329.036
R157 VTAIL.n393 VTAIL.t4 329.036
R158 VTAIL.n331 VTAIL.t6 329.036
R159 VTAIL.n269 VTAIL.t3 329.036
R160 VTAIL.n207 VTAIL.t0 329.036
R161 VTAIL.n456 VTAIL.n455 171.744
R162 VTAIL.n456 VTAIL.n449 171.744
R163 VTAIL.n463 VTAIL.n449 171.744
R164 VTAIL.n464 VTAIL.n463 171.744
R165 VTAIL.n464 VTAIL.n445 171.744
R166 VTAIL.n472 VTAIL.n445 171.744
R167 VTAIL.n473 VTAIL.n472 171.744
R168 VTAIL.n474 VTAIL.n473 171.744
R169 VTAIL.n474 VTAIL.n441 171.744
R170 VTAIL.n481 VTAIL.n441 171.744
R171 VTAIL.n482 VTAIL.n481 171.744
R172 VTAIL.n482 VTAIL.n437 171.744
R173 VTAIL.n489 VTAIL.n437 171.744
R174 VTAIL.n490 VTAIL.n489 171.744
R175 VTAIL.n22 VTAIL.n21 171.744
R176 VTAIL.n22 VTAIL.n15 171.744
R177 VTAIL.n29 VTAIL.n15 171.744
R178 VTAIL.n30 VTAIL.n29 171.744
R179 VTAIL.n30 VTAIL.n11 171.744
R180 VTAIL.n38 VTAIL.n11 171.744
R181 VTAIL.n39 VTAIL.n38 171.744
R182 VTAIL.n40 VTAIL.n39 171.744
R183 VTAIL.n40 VTAIL.n7 171.744
R184 VTAIL.n47 VTAIL.n7 171.744
R185 VTAIL.n48 VTAIL.n47 171.744
R186 VTAIL.n48 VTAIL.n3 171.744
R187 VTAIL.n55 VTAIL.n3 171.744
R188 VTAIL.n56 VTAIL.n55 171.744
R189 VTAIL.n84 VTAIL.n83 171.744
R190 VTAIL.n84 VTAIL.n77 171.744
R191 VTAIL.n91 VTAIL.n77 171.744
R192 VTAIL.n92 VTAIL.n91 171.744
R193 VTAIL.n92 VTAIL.n73 171.744
R194 VTAIL.n100 VTAIL.n73 171.744
R195 VTAIL.n101 VTAIL.n100 171.744
R196 VTAIL.n102 VTAIL.n101 171.744
R197 VTAIL.n102 VTAIL.n69 171.744
R198 VTAIL.n109 VTAIL.n69 171.744
R199 VTAIL.n110 VTAIL.n109 171.744
R200 VTAIL.n110 VTAIL.n65 171.744
R201 VTAIL.n117 VTAIL.n65 171.744
R202 VTAIL.n118 VTAIL.n117 171.744
R203 VTAIL.n146 VTAIL.n145 171.744
R204 VTAIL.n146 VTAIL.n139 171.744
R205 VTAIL.n153 VTAIL.n139 171.744
R206 VTAIL.n154 VTAIL.n153 171.744
R207 VTAIL.n154 VTAIL.n135 171.744
R208 VTAIL.n162 VTAIL.n135 171.744
R209 VTAIL.n163 VTAIL.n162 171.744
R210 VTAIL.n164 VTAIL.n163 171.744
R211 VTAIL.n164 VTAIL.n131 171.744
R212 VTAIL.n171 VTAIL.n131 171.744
R213 VTAIL.n172 VTAIL.n171 171.744
R214 VTAIL.n172 VTAIL.n127 171.744
R215 VTAIL.n179 VTAIL.n127 171.744
R216 VTAIL.n180 VTAIL.n179 171.744
R217 VTAIL.n428 VTAIL.n427 171.744
R218 VTAIL.n427 VTAIL.n375 171.744
R219 VTAIL.n420 VTAIL.n375 171.744
R220 VTAIL.n420 VTAIL.n419 171.744
R221 VTAIL.n419 VTAIL.n379 171.744
R222 VTAIL.n384 VTAIL.n379 171.744
R223 VTAIL.n412 VTAIL.n384 171.744
R224 VTAIL.n412 VTAIL.n411 171.744
R225 VTAIL.n411 VTAIL.n385 171.744
R226 VTAIL.n404 VTAIL.n385 171.744
R227 VTAIL.n404 VTAIL.n403 171.744
R228 VTAIL.n403 VTAIL.n389 171.744
R229 VTAIL.n396 VTAIL.n389 171.744
R230 VTAIL.n396 VTAIL.n395 171.744
R231 VTAIL.n366 VTAIL.n365 171.744
R232 VTAIL.n365 VTAIL.n313 171.744
R233 VTAIL.n358 VTAIL.n313 171.744
R234 VTAIL.n358 VTAIL.n357 171.744
R235 VTAIL.n357 VTAIL.n317 171.744
R236 VTAIL.n322 VTAIL.n317 171.744
R237 VTAIL.n350 VTAIL.n322 171.744
R238 VTAIL.n350 VTAIL.n349 171.744
R239 VTAIL.n349 VTAIL.n323 171.744
R240 VTAIL.n342 VTAIL.n323 171.744
R241 VTAIL.n342 VTAIL.n341 171.744
R242 VTAIL.n341 VTAIL.n327 171.744
R243 VTAIL.n334 VTAIL.n327 171.744
R244 VTAIL.n334 VTAIL.n333 171.744
R245 VTAIL.n304 VTAIL.n303 171.744
R246 VTAIL.n303 VTAIL.n251 171.744
R247 VTAIL.n296 VTAIL.n251 171.744
R248 VTAIL.n296 VTAIL.n295 171.744
R249 VTAIL.n295 VTAIL.n255 171.744
R250 VTAIL.n260 VTAIL.n255 171.744
R251 VTAIL.n288 VTAIL.n260 171.744
R252 VTAIL.n288 VTAIL.n287 171.744
R253 VTAIL.n287 VTAIL.n261 171.744
R254 VTAIL.n280 VTAIL.n261 171.744
R255 VTAIL.n280 VTAIL.n279 171.744
R256 VTAIL.n279 VTAIL.n265 171.744
R257 VTAIL.n272 VTAIL.n265 171.744
R258 VTAIL.n272 VTAIL.n271 171.744
R259 VTAIL.n242 VTAIL.n241 171.744
R260 VTAIL.n241 VTAIL.n189 171.744
R261 VTAIL.n234 VTAIL.n189 171.744
R262 VTAIL.n234 VTAIL.n233 171.744
R263 VTAIL.n233 VTAIL.n193 171.744
R264 VTAIL.n198 VTAIL.n193 171.744
R265 VTAIL.n226 VTAIL.n198 171.744
R266 VTAIL.n226 VTAIL.n225 171.744
R267 VTAIL.n225 VTAIL.n199 171.744
R268 VTAIL.n218 VTAIL.n199 171.744
R269 VTAIL.n218 VTAIL.n217 171.744
R270 VTAIL.n217 VTAIL.n203 171.744
R271 VTAIL.n210 VTAIL.n203 171.744
R272 VTAIL.n210 VTAIL.n209 171.744
R273 VTAIL.n455 VTAIL.t1 85.8723
R274 VTAIL.n21 VTAIL.t2 85.8723
R275 VTAIL.n83 VTAIL.t5 85.8723
R276 VTAIL.n145 VTAIL.t7 85.8723
R277 VTAIL.n395 VTAIL.t4 85.8723
R278 VTAIL.n333 VTAIL.t6 85.8723
R279 VTAIL.n271 VTAIL.t3 85.8723
R280 VTAIL.n209 VTAIL.t0 85.8723
R281 VTAIL.n495 VTAIL.n494 34.9005
R282 VTAIL.n61 VTAIL.n60 34.9005
R283 VTAIL.n123 VTAIL.n122 34.9005
R284 VTAIL.n185 VTAIL.n184 34.9005
R285 VTAIL.n433 VTAIL.n432 34.9005
R286 VTAIL.n371 VTAIL.n370 34.9005
R287 VTAIL.n309 VTAIL.n308 34.9005
R288 VTAIL.n247 VTAIL.n246 34.9005
R289 VTAIL.n495 VTAIL.n433 23.6686
R290 VTAIL.n247 VTAIL.n185 23.6686
R291 VTAIL.n475 VTAIL.n442 13.1884
R292 VTAIL.n41 VTAIL.n8 13.1884
R293 VTAIL.n103 VTAIL.n70 13.1884
R294 VTAIL.n165 VTAIL.n132 13.1884
R295 VTAIL.n382 VTAIL.n380 13.1884
R296 VTAIL.n320 VTAIL.n318 13.1884
R297 VTAIL.n258 VTAIL.n256 13.1884
R298 VTAIL.n196 VTAIL.n194 13.1884
R299 VTAIL.n476 VTAIL.n444 12.8005
R300 VTAIL.n480 VTAIL.n479 12.8005
R301 VTAIL.n42 VTAIL.n10 12.8005
R302 VTAIL.n46 VTAIL.n45 12.8005
R303 VTAIL.n104 VTAIL.n72 12.8005
R304 VTAIL.n108 VTAIL.n107 12.8005
R305 VTAIL.n166 VTAIL.n134 12.8005
R306 VTAIL.n170 VTAIL.n169 12.8005
R307 VTAIL.n418 VTAIL.n417 12.8005
R308 VTAIL.n414 VTAIL.n413 12.8005
R309 VTAIL.n356 VTAIL.n355 12.8005
R310 VTAIL.n352 VTAIL.n351 12.8005
R311 VTAIL.n294 VTAIL.n293 12.8005
R312 VTAIL.n290 VTAIL.n289 12.8005
R313 VTAIL.n232 VTAIL.n231 12.8005
R314 VTAIL.n228 VTAIL.n227 12.8005
R315 VTAIL.n471 VTAIL.n470 12.0247
R316 VTAIL.n483 VTAIL.n440 12.0247
R317 VTAIL.n37 VTAIL.n36 12.0247
R318 VTAIL.n49 VTAIL.n6 12.0247
R319 VTAIL.n99 VTAIL.n98 12.0247
R320 VTAIL.n111 VTAIL.n68 12.0247
R321 VTAIL.n161 VTAIL.n160 12.0247
R322 VTAIL.n173 VTAIL.n130 12.0247
R323 VTAIL.n421 VTAIL.n378 12.0247
R324 VTAIL.n410 VTAIL.n383 12.0247
R325 VTAIL.n359 VTAIL.n316 12.0247
R326 VTAIL.n348 VTAIL.n321 12.0247
R327 VTAIL.n297 VTAIL.n254 12.0247
R328 VTAIL.n286 VTAIL.n259 12.0247
R329 VTAIL.n235 VTAIL.n192 12.0247
R330 VTAIL.n224 VTAIL.n197 12.0247
R331 VTAIL.n469 VTAIL.n446 11.249
R332 VTAIL.n484 VTAIL.n438 11.249
R333 VTAIL.n35 VTAIL.n12 11.249
R334 VTAIL.n50 VTAIL.n4 11.249
R335 VTAIL.n97 VTAIL.n74 11.249
R336 VTAIL.n112 VTAIL.n66 11.249
R337 VTAIL.n159 VTAIL.n136 11.249
R338 VTAIL.n174 VTAIL.n128 11.249
R339 VTAIL.n422 VTAIL.n376 11.249
R340 VTAIL.n409 VTAIL.n386 11.249
R341 VTAIL.n360 VTAIL.n314 11.249
R342 VTAIL.n347 VTAIL.n324 11.249
R343 VTAIL.n298 VTAIL.n252 11.249
R344 VTAIL.n285 VTAIL.n262 11.249
R345 VTAIL.n236 VTAIL.n190 11.249
R346 VTAIL.n223 VTAIL.n200 11.249
R347 VTAIL.n454 VTAIL.n453 10.7239
R348 VTAIL.n20 VTAIL.n19 10.7239
R349 VTAIL.n82 VTAIL.n81 10.7239
R350 VTAIL.n144 VTAIL.n143 10.7239
R351 VTAIL.n394 VTAIL.n393 10.7239
R352 VTAIL.n332 VTAIL.n331 10.7239
R353 VTAIL.n270 VTAIL.n269 10.7239
R354 VTAIL.n208 VTAIL.n207 10.7239
R355 VTAIL.n466 VTAIL.n465 10.4732
R356 VTAIL.n488 VTAIL.n487 10.4732
R357 VTAIL.n32 VTAIL.n31 10.4732
R358 VTAIL.n54 VTAIL.n53 10.4732
R359 VTAIL.n94 VTAIL.n93 10.4732
R360 VTAIL.n116 VTAIL.n115 10.4732
R361 VTAIL.n156 VTAIL.n155 10.4732
R362 VTAIL.n178 VTAIL.n177 10.4732
R363 VTAIL.n426 VTAIL.n425 10.4732
R364 VTAIL.n406 VTAIL.n405 10.4732
R365 VTAIL.n364 VTAIL.n363 10.4732
R366 VTAIL.n344 VTAIL.n343 10.4732
R367 VTAIL.n302 VTAIL.n301 10.4732
R368 VTAIL.n282 VTAIL.n281 10.4732
R369 VTAIL.n240 VTAIL.n239 10.4732
R370 VTAIL.n220 VTAIL.n219 10.4732
R371 VTAIL.n462 VTAIL.n448 9.69747
R372 VTAIL.n491 VTAIL.n436 9.69747
R373 VTAIL.n28 VTAIL.n14 9.69747
R374 VTAIL.n57 VTAIL.n2 9.69747
R375 VTAIL.n90 VTAIL.n76 9.69747
R376 VTAIL.n119 VTAIL.n64 9.69747
R377 VTAIL.n152 VTAIL.n138 9.69747
R378 VTAIL.n181 VTAIL.n126 9.69747
R379 VTAIL.n429 VTAIL.n374 9.69747
R380 VTAIL.n402 VTAIL.n388 9.69747
R381 VTAIL.n367 VTAIL.n312 9.69747
R382 VTAIL.n340 VTAIL.n326 9.69747
R383 VTAIL.n305 VTAIL.n250 9.69747
R384 VTAIL.n278 VTAIL.n264 9.69747
R385 VTAIL.n243 VTAIL.n188 9.69747
R386 VTAIL.n216 VTAIL.n202 9.69747
R387 VTAIL.n494 VTAIL.n493 9.45567
R388 VTAIL.n60 VTAIL.n59 9.45567
R389 VTAIL.n122 VTAIL.n121 9.45567
R390 VTAIL.n184 VTAIL.n183 9.45567
R391 VTAIL.n432 VTAIL.n431 9.45567
R392 VTAIL.n370 VTAIL.n369 9.45567
R393 VTAIL.n308 VTAIL.n307 9.45567
R394 VTAIL.n246 VTAIL.n245 9.45567
R395 VTAIL.n493 VTAIL.n492 9.3005
R396 VTAIL.n436 VTAIL.n435 9.3005
R397 VTAIL.n487 VTAIL.n486 9.3005
R398 VTAIL.n485 VTAIL.n484 9.3005
R399 VTAIL.n440 VTAIL.n439 9.3005
R400 VTAIL.n479 VTAIL.n478 9.3005
R401 VTAIL.n452 VTAIL.n451 9.3005
R402 VTAIL.n459 VTAIL.n458 9.3005
R403 VTAIL.n461 VTAIL.n460 9.3005
R404 VTAIL.n448 VTAIL.n447 9.3005
R405 VTAIL.n467 VTAIL.n466 9.3005
R406 VTAIL.n469 VTAIL.n468 9.3005
R407 VTAIL.n470 VTAIL.n443 9.3005
R408 VTAIL.n477 VTAIL.n476 9.3005
R409 VTAIL.n59 VTAIL.n58 9.3005
R410 VTAIL.n2 VTAIL.n1 9.3005
R411 VTAIL.n53 VTAIL.n52 9.3005
R412 VTAIL.n51 VTAIL.n50 9.3005
R413 VTAIL.n6 VTAIL.n5 9.3005
R414 VTAIL.n45 VTAIL.n44 9.3005
R415 VTAIL.n18 VTAIL.n17 9.3005
R416 VTAIL.n25 VTAIL.n24 9.3005
R417 VTAIL.n27 VTAIL.n26 9.3005
R418 VTAIL.n14 VTAIL.n13 9.3005
R419 VTAIL.n33 VTAIL.n32 9.3005
R420 VTAIL.n35 VTAIL.n34 9.3005
R421 VTAIL.n36 VTAIL.n9 9.3005
R422 VTAIL.n43 VTAIL.n42 9.3005
R423 VTAIL.n121 VTAIL.n120 9.3005
R424 VTAIL.n64 VTAIL.n63 9.3005
R425 VTAIL.n115 VTAIL.n114 9.3005
R426 VTAIL.n113 VTAIL.n112 9.3005
R427 VTAIL.n68 VTAIL.n67 9.3005
R428 VTAIL.n107 VTAIL.n106 9.3005
R429 VTAIL.n80 VTAIL.n79 9.3005
R430 VTAIL.n87 VTAIL.n86 9.3005
R431 VTAIL.n89 VTAIL.n88 9.3005
R432 VTAIL.n76 VTAIL.n75 9.3005
R433 VTAIL.n95 VTAIL.n94 9.3005
R434 VTAIL.n97 VTAIL.n96 9.3005
R435 VTAIL.n98 VTAIL.n71 9.3005
R436 VTAIL.n105 VTAIL.n104 9.3005
R437 VTAIL.n183 VTAIL.n182 9.3005
R438 VTAIL.n126 VTAIL.n125 9.3005
R439 VTAIL.n177 VTAIL.n176 9.3005
R440 VTAIL.n175 VTAIL.n174 9.3005
R441 VTAIL.n130 VTAIL.n129 9.3005
R442 VTAIL.n169 VTAIL.n168 9.3005
R443 VTAIL.n142 VTAIL.n141 9.3005
R444 VTAIL.n149 VTAIL.n148 9.3005
R445 VTAIL.n151 VTAIL.n150 9.3005
R446 VTAIL.n138 VTAIL.n137 9.3005
R447 VTAIL.n157 VTAIL.n156 9.3005
R448 VTAIL.n159 VTAIL.n158 9.3005
R449 VTAIL.n160 VTAIL.n133 9.3005
R450 VTAIL.n167 VTAIL.n166 9.3005
R451 VTAIL.n392 VTAIL.n391 9.3005
R452 VTAIL.n399 VTAIL.n398 9.3005
R453 VTAIL.n401 VTAIL.n400 9.3005
R454 VTAIL.n388 VTAIL.n387 9.3005
R455 VTAIL.n407 VTAIL.n406 9.3005
R456 VTAIL.n409 VTAIL.n408 9.3005
R457 VTAIL.n383 VTAIL.n381 9.3005
R458 VTAIL.n415 VTAIL.n414 9.3005
R459 VTAIL.n431 VTAIL.n430 9.3005
R460 VTAIL.n374 VTAIL.n373 9.3005
R461 VTAIL.n425 VTAIL.n424 9.3005
R462 VTAIL.n423 VTAIL.n422 9.3005
R463 VTAIL.n378 VTAIL.n377 9.3005
R464 VTAIL.n417 VTAIL.n416 9.3005
R465 VTAIL.n330 VTAIL.n329 9.3005
R466 VTAIL.n337 VTAIL.n336 9.3005
R467 VTAIL.n339 VTAIL.n338 9.3005
R468 VTAIL.n326 VTAIL.n325 9.3005
R469 VTAIL.n345 VTAIL.n344 9.3005
R470 VTAIL.n347 VTAIL.n346 9.3005
R471 VTAIL.n321 VTAIL.n319 9.3005
R472 VTAIL.n353 VTAIL.n352 9.3005
R473 VTAIL.n369 VTAIL.n368 9.3005
R474 VTAIL.n312 VTAIL.n311 9.3005
R475 VTAIL.n363 VTAIL.n362 9.3005
R476 VTAIL.n361 VTAIL.n360 9.3005
R477 VTAIL.n316 VTAIL.n315 9.3005
R478 VTAIL.n355 VTAIL.n354 9.3005
R479 VTAIL.n268 VTAIL.n267 9.3005
R480 VTAIL.n275 VTAIL.n274 9.3005
R481 VTAIL.n277 VTAIL.n276 9.3005
R482 VTAIL.n264 VTAIL.n263 9.3005
R483 VTAIL.n283 VTAIL.n282 9.3005
R484 VTAIL.n285 VTAIL.n284 9.3005
R485 VTAIL.n259 VTAIL.n257 9.3005
R486 VTAIL.n291 VTAIL.n290 9.3005
R487 VTAIL.n307 VTAIL.n306 9.3005
R488 VTAIL.n250 VTAIL.n249 9.3005
R489 VTAIL.n301 VTAIL.n300 9.3005
R490 VTAIL.n299 VTAIL.n298 9.3005
R491 VTAIL.n254 VTAIL.n253 9.3005
R492 VTAIL.n293 VTAIL.n292 9.3005
R493 VTAIL.n206 VTAIL.n205 9.3005
R494 VTAIL.n213 VTAIL.n212 9.3005
R495 VTAIL.n215 VTAIL.n214 9.3005
R496 VTAIL.n202 VTAIL.n201 9.3005
R497 VTAIL.n221 VTAIL.n220 9.3005
R498 VTAIL.n223 VTAIL.n222 9.3005
R499 VTAIL.n197 VTAIL.n195 9.3005
R500 VTAIL.n229 VTAIL.n228 9.3005
R501 VTAIL.n245 VTAIL.n244 9.3005
R502 VTAIL.n188 VTAIL.n187 9.3005
R503 VTAIL.n239 VTAIL.n238 9.3005
R504 VTAIL.n237 VTAIL.n236 9.3005
R505 VTAIL.n192 VTAIL.n191 9.3005
R506 VTAIL.n231 VTAIL.n230 9.3005
R507 VTAIL.n461 VTAIL.n450 8.92171
R508 VTAIL.n492 VTAIL.n434 8.92171
R509 VTAIL.n27 VTAIL.n16 8.92171
R510 VTAIL.n58 VTAIL.n0 8.92171
R511 VTAIL.n89 VTAIL.n78 8.92171
R512 VTAIL.n120 VTAIL.n62 8.92171
R513 VTAIL.n151 VTAIL.n140 8.92171
R514 VTAIL.n182 VTAIL.n124 8.92171
R515 VTAIL.n430 VTAIL.n372 8.92171
R516 VTAIL.n401 VTAIL.n390 8.92171
R517 VTAIL.n368 VTAIL.n310 8.92171
R518 VTAIL.n339 VTAIL.n328 8.92171
R519 VTAIL.n306 VTAIL.n248 8.92171
R520 VTAIL.n277 VTAIL.n266 8.92171
R521 VTAIL.n244 VTAIL.n186 8.92171
R522 VTAIL.n215 VTAIL.n204 8.92171
R523 VTAIL.n458 VTAIL.n457 8.14595
R524 VTAIL.n24 VTAIL.n23 8.14595
R525 VTAIL.n86 VTAIL.n85 8.14595
R526 VTAIL.n148 VTAIL.n147 8.14595
R527 VTAIL.n398 VTAIL.n397 8.14595
R528 VTAIL.n336 VTAIL.n335 8.14595
R529 VTAIL.n274 VTAIL.n273 8.14595
R530 VTAIL.n212 VTAIL.n211 8.14595
R531 VTAIL.n454 VTAIL.n452 7.3702
R532 VTAIL.n20 VTAIL.n18 7.3702
R533 VTAIL.n82 VTAIL.n80 7.3702
R534 VTAIL.n144 VTAIL.n142 7.3702
R535 VTAIL.n394 VTAIL.n392 7.3702
R536 VTAIL.n332 VTAIL.n330 7.3702
R537 VTAIL.n270 VTAIL.n268 7.3702
R538 VTAIL.n208 VTAIL.n206 7.3702
R539 VTAIL.n457 VTAIL.n452 5.81868
R540 VTAIL.n23 VTAIL.n18 5.81868
R541 VTAIL.n85 VTAIL.n80 5.81868
R542 VTAIL.n147 VTAIL.n142 5.81868
R543 VTAIL.n397 VTAIL.n392 5.81868
R544 VTAIL.n335 VTAIL.n330 5.81868
R545 VTAIL.n273 VTAIL.n268 5.81868
R546 VTAIL.n211 VTAIL.n206 5.81868
R547 VTAIL.n458 VTAIL.n450 5.04292
R548 VTAIL.n494 VTAIL.n434 5.04292
R549 VTAIL.n24 VTAIL.n16 5.04292
R550 VTAIL.n60 VTAIL.n0 5.04292
R551 VTAIL.n86 VTAIL.n78 5.04292
R552 VTAIL.n122 VTAIL.n62 5.04292
R553 VTAIL.n148 VTAIL.n140 5.04292
R554 VTAIL.n184 VTAIL.n124 5.04292
R555 VTAIL.n432 VTAIL.n372 5.04292
R556 VTAIL.n398 VTAIL.n390 5.04292
R557 VTAIL.n370 VTAIL.n310 5.04292
R558 VTAIL.n336 VTAIL.n328 5.04292
R559 VTAIL.n308 VTAIL.n248 5.04292
R560 VTAIL.n274 VTAIL.n266 5.04292
R561 VTAIL.n246 VTAIL.n186 5.04292
R562 VTAIL.n212 VTAIL.n204 5.04292
R563 VTAIL.n462 VTAIL.n461 4.26717
R564 VTAIL.n492 VTAIL.n491 4.26717
R565 VTAIL.n28 VTAIL.n27 4.26717
R566 VTAIL.n58 VTAIL.n57 4.26717
R567 VTAIL.n90 VTAIL.n89 4.26717
R568 VTAIL.n120 VTAIL.n119 4.26717
R569 VTAIL.n152 VTAIL.n151 4.26717
R570 VTAIL.n182 VTAIL.n181 4.26717
R571 VTAIL.n430 VTAIL.n429 4.26717
R572 VTAIL.n402 VTAIL.n401 4.26717
R573 VTAIL.n368 VTAIL.n367 4.26717
R574 VTAIL.n340 VTAIL.n339 4.26717
R575 VTAIL.n306 VTAIL.n305 4.26717
R576 VTAIL.n278 VTAIL.n277 4.26717
R577 VTAIL.n244 VTAIL.n243 4.26717
R578 VTAIL.n216 VTAIL.n215 4.26717
R579 VTAIL.n465 VTAIL.n448 3.49141
R580 VTAIL.n488 VTAIL.n436 3.49141
R581 VTAIL.n31 VTAIL.n14 3.49141
R582 VTAIL.n54 VTAIL.n2 3.49141
R583 VTAIL.n93 VTAIL.n76 3.49141
R584 VTAIL.n116 VTAIL.n64 3.49141
R585 VTAIL.n155 VTAIL.n138 3.49141
R586 VTAIL.n178 VTAIL.n126 3.49141
R587 VTAIL.n426 VTAIL.n374 3.49141
R588 VTAIL.n405 VTAIL.n388 3.49141
R589 VTAIL.n364 VTAIL.n312 3.49141
R590 VTAIL.n343 VTAIL.n326 3.49141
R591 VTAIL.n302 VTAIL.n250 3.49141
R592 VTAIL.n281 VTAIL.n264 3.49141
R593 VTAIL.n240 VTAIL.n188 3.49141
R594 VTAIL.n219 VTAIL.n202 3.49141
R595 VTAIL.n466 VTAIL.n446 2.71565
R596 VTAIL.n487 VTAIL.n438 2.71565
R597 VTAIL.n32 VTAIL.n12 2.71565
R598 VTAIL.n53 VTAIL.n4 2.71565
R599 VTAIL.n94 VTAIL.n74 2.71565
R600 VTAIL.n115 VTAIL.n66 2.71565
R601 VTAIL.n156 VTAIL.n136 2.71565
R602 VTAIL.n177 VTAIL.n128 2.71565
R603 VTAIL.n425 VTAIL.n376 2.71565
R604 VTAIL.n406 VTAIL.n386 2.71565
R605 VTAIL.n363 VTAIL.n314 2.71565
R606 VTAIL.n344 VTAIL.n324 2.71565
R607 VTAIL.n301 VTAIL.n252 2.71565
R608 VTAIL.n282 VTAIL.n262 2.71565
R609 VTAIL.n239 VTAIL.n190 2.71565
R610 VTAIL.n220 VTAIL.n200 2.71565
R611 VTAIL.n453 VTAIL.n451 2.41282
R612 VTAIL.n19 VTAIL.n17 2.41282
R613 VTAIL.n81 VTAIL.n79 2.41282
R614 VTAIL.n143 VTAIL.n141 2.41282
R615 VTAIL.n393 VTAIL.n391 2.41282
R616 VTAIL.n331 VTAIL.n329 2.41282
R617 VTAIL.n269 VTAIL.n267 2.41282
R618 VTAIL.n207 VTAIL.n205 2.41282
R619 VTAIL.n471 VTAIL.n469 1.93989
R620 VTAIL.n484 VTAIL.n483 1.93989
R621 VTAIL.n37 VTAIL.n35 1.93989
R622 VTAIL.n50 VTAIL.n49 1.93989
R623 VTAIL.n99 VTAIL.n97 1.93989
R624 VTAIL.n112 VTAIL.n111 1.93989
R625 VTAIL.n161 VTAIL.n159 1.93989
R626 VTAIL.n174 VTAIL.n173 1.93989
R627 VTAIL.n422 VTAIL.n421 1.93989
R628 VTAIL.n410 VTAIL.n409 1.93989
R629 VTAIL.n360 VTAIL.n359 1.93989
R630 VTAIL.n348 VTAIL.n347 1.93989
R631 VTAIL.n298 VTAIL.n297 1.93989
R632 VTAIL.n286 VTAIL.n285 1.93989
R633 VTAIL.n236 VTAIL.n235 1.93989
R634 VTAIL.n224 VTAIL.n223 1.93989
R635 VTAIL.n309 VTAIL.n247 1.35395
R636 VTAIL.n433 VTAIL.n371 1.35395
R637 VTAIL.n185 VTAIL.n123 1.35395
R638 VTAIL.n470 VTAIL.n444 1.16414
R639 VTAIL.n480 VTAIL.n440 1.16414
R640 VTAIL.n36 VTAIL.n10 1.16414
R641 VTAIL.n46 VTAIL.n6 1.16414
R642 VTAIL.n98 VTAIL.n72 1.16414
R643 VTAIL.n108 VTAIL.n68 1.16414
R644 VTAIL.n160 VTAIL.n134 1.16414
R645 VTAIL.n170 VTAIL.n130 1.16414
R646 VTAIL.n418 VTAIL.n378 1.16414
R647 VTAIL.n413 VTAIL.n383 1.16414
R648 VTAIL.n356 VTAIL.n316 1.16414
R649 VTAIL.n351 VTAIL.n321 1.16414
R650 VTAIL.n294 VTAIL.n254 1.16414
R651 VTAIL.n289 VTAIL.n259 1.16414
R652 VTAIL.n232 VTAIL.n192 1.16414
R653 VTAIL.n227 VTAIL.n197 1.16414
R654 VTAIL VTAIL.n61 0.735414
R655 VTAIL VTAIL.n495 0.619035
R656 VTAIL.n371 VTAIL.n309 0.470328
R657 VTAIL.n123 VTAIL.n61 0.470328
R658 VTAIL.n476 VTAIL.n475 0.388379
R659 VTAIL.n479 VTAIL.n442 0.388379
R660 VTAIL.n42 VTAIL.n41 0.388379
R661 VTAIL.n45 VTAIL.n8 0.388379
R662 VTAIL.n104 VTAIL.n103 0.388379
R663 VTAIL.n107 VTAIL.n70 0.388379
R664 VTAIL.n166 VTAIL.n165 0.388379
R665 VTAIL.n169 VTAIL.n132 0.388379
R666 VTAIL.n417 VTAIL.n380 0.388379
R667 VTAIL.n414 VTAIL.n382 0.388379
R668 VTAIL.n355 VTAIL.n318 0.388379
R669 VTAIL.n352 VTAIL.n320 0.388379
R670 VTAIL.n293 VTAIL.n256 0.388379
R671 VTAIL.n290 VTAIL.n258 0.388379
R672 VTAIL.n231 VTAIL.n194 0.388379
R673 VTAIL.n228 VTAIL.n196 0.388379
R674 VTAIL.n459 VTAIL.n451 0.155672
R675 VTAIL.n460 VTAIL.n459 0.155672
R676 VTAIL.n460 VTAIL.n447 0.155672
R677 VTAIL.n467 VTAIL.n447 0.155672
R678 VTAIL.n468 VTAIL.n467 0.155672
R679 VTAIL.n468 VTAIL.n443 0.155672
R680 VTAIL.n477 VTAIL.n443 0.155672
R681 VTAIL.n478 VTAIL.n477 0.155672
R682 VTAIL.n478 VTAIL.n439 0.155672
R683 VTAIL.n485 VTAIL.n439 0.155672
R684 VTAIL.n486 VTAIL.n485 0.155672
R685 VTAIL.n486 VTAIL.n435 0.155672
R686 VTAIL.n493 VTAIL.n435 0.155672
R687 VTAIL.n25 VTAIL.n17 0.155672
R688 VTAIL.n26 VTAIL.n25 0.155672
R689 VTAIL.n26 VTAIL.n13 0.155672
R690 VTAIL.n33 VTAIL.n13 0.155672
R691 VTAIL.n34 VTAIL.n33 0.155672
R692 VTAIL.n34 VTAIL.n9 0.155672
R693 VTAIL.n43 VTAIL.n9 0.155672
R694 VTAIL.n44 VTAIL.n43 0.155672
R695 VTAIL.n44 VTAIL.n5 0.155672
R696 VTAIL.n51 VTAIL.n5 0.155672
R697 VTAIL.n52 VTAIL.n51 0.155672
R698 VTAIL.n52 VTAIL.n1 0.155672
R699 VTAIL.n59 VTAIL.n1 0.155672
R700 VTAIL.n87 VTAIL.n79 0.155672
R701 VTAIL.n88 VTAIL.n87 0.155672
R702 VTAIL.n88 VTAIL.n75 0.155672
R703 VTAIL.n95 VTAIL.n75 0.155672
R704 VTAIL.n96 VTAIL.n95 0.155672
R705 VTAIL.n96 VTAIL.n71 0.155672
R706 VTAIL.n105 VTAIL.n71 0.155672
R707 VTAIL.n106 VTAIL.n105 0.155672
R708 VTAIL.n106 VTAIL.n67 0.155672
R709 VTAIL.n113 VTAIL.n67 0.155672
R710 VTAIL.n114 VTAIL.n113 0.155672
R711 VTAIL.n114 VTAIL.n63 0.155672
R712 VTAIL.n121 VTAIL.n63 0.155672
R713 VTAIL.n149 VTAIL.n141 0.155672
R714 VTAIL.n150 VTAIL.n149 0.155672
R715 VTAIL.n150 VTAIL.n137 0.155672
R716 VTAIL.n157 VTAIL.n137 0.155672
R717 VTAIL.n158 VTAIL.n157 0.155672
R718 VTAIL.n158 VTAIL.n133 0.155672
R719 VTAIL.n167 VTAIL.n133 0.155672
R720 VTAIL.n168 VTAIL.n167 0.155672
R721 VTAIL.n168 VTAIL.n129 0.155672
R722 VTAIL.n175 VTAIL.n129 0.155672
R723 VTAIL.n176 VTAIL.n175 0.155672
R724 VTAIL.n176 VTAIL.n125 0.155672
R725 VTAIL.n183 VTAIL.n125 0.155672
R726 VTAIL.n431 VTAIL.n373 0.155672
R727 VTAIL.n424 VTAIL.n373 0.155672
R728 VTAIL.n424 VTAIL.n423 0.155672
R729 VTAIL.n423 VTAIL.n377 0.155672
R730 VTAIL.n416 VTAIL.n377 0.155672
R731 VTAIL.n416 VTAIL.n415 0.155672
R732 VTAIL.n415 VTAIL.n381 0.155672
R733 VTAIL.n408 VTAIL.n381 0.155672
R734 VTAIL.n408 VTAIL.n407 0.155672
R735 VTAIL.n407 VTAIL.n387 0.155672
R736 VTAIL.n400 VTAIL.n387 0.155672
R737 VTAIL.n400 VTAIL.n399 0.155672
R738 VTAIL.n399 VTAIL.n391 0.155672
R739 VTAIL.n369 VTAIL.n311 0.155672
R740 VTAIL.n362 VTAIL.n311 0.155672
R741 VTAIL.n362 VTAIL.n361 0.155672
R742 VTAIL.n361 VTAIL.n315 0.155672
R743 VTAIL.n354 VTAIL.n315 0.155672
R744 VTAIL.n354 VTAIL.n353 0.155672
R745 VTAIL.n353 VTAIL.n319 0.155672
R746 VTAIL.n346 VTAIL.n319 0.155672
R747 VTAIL.n346 VTAIL.n345 0.155672
R748 VTAIL.n345 VTAIL.n325 0.155672
R749 VTAIL.n338 VTAIL.n325 0.155672
R750 VTAIL.n338 VTAIL.n337 0.155672
R751 VTAIL.n337 VTAIL.n329 0.155672
R752 VTAIL.n307 VTAIL.n249 0.155672
R753 VTAIL.n300 VTAIL.n249 0.155672
R754 VTAIL.n300 VTAIL.n299 0.155672
R755 VTAIL.n299 VTAIL.n253 0.155672
R756 VTAIL.n292 VTAIL.n253 0.155672
R757 VTAIL.n292 VTAIL.n291 0.155672
R758 VTAIL.n291 VTAIL.n257 0.155672
R759 VTAIL.n284 VTAIL.n257 0.155672
R760 VTAIL.n284 VTAIL.n283 0.155672
R761 VTAIL.n283 VTAIL.n263 0.155672
R762 VTAIL.n276 VTAIL.n263 0.155672
R763 VTAIL.n276 VTAIL.n275 0.155672
R764 VTAIL.n275 VTAIL.n267 0.155672
R765 VTAIL.n245 VTAIL.n187 0.155672
R766 VTAIL.n238 VTAIL.n187 0.155672
R767 VTAIL.n238 VTAIL.n237 0.155672
R768 VTAIL.n237 VTAIL.n191 0.155672
R769 VTAIL.n230 VTAIL.n191 0.155672
R770 VTAIL.n230 VTAIL.n229 0.155672
R771 VTAIL.n229 VTAIL.n195 0.155672
R772 VTAIL.n222 VTAIL.n195 0.155672
R773 VTAIL.n222 VTAIL.n221 0.155672
R774 VTAIL.n221 VTAIL.n201 0.155672
R775 VTAIL.n214 VTAIL.n201 0.155672
R776 VTAIL.n214 VTAIL.n213 0.155672
R777 VTAIL.n213 VTAIL.n205 0.155672
R778 B.n381 B.n62 585
R779 B.n383 B.n382 585
R780 B.n384 B.n61 585
R781 B.n386 B.n385 585
R782 B.n387 B.n60 585
R783 B.n389 B.n388 585
R784 B.n390 B.n59 585
R785 B.n392 B.n391 585
R786 B.n393 B.n58 585
R787 B.n395 B.n394 585
R788 B.n396 B.n57 585
R789 B.n398 B.n397 585
R790 B.n399 B.n56 585
R791 B.n401 B.n400 585
R792 B.n402 B.n55 585
R793 B.n404 B.n403 585
R794 B.n405 B.n54 585
R795 B.n407 B.n406 585
R796 B.n408 B.n53 585
R797 B.n410 B.n409 585
R798 B.n411 B.n52 585
R799 B.n413 B.n412 585
R800 B.n414 B.n51 585
R801 B.n416 B.n415 585
R802 B.n417 B.n50 585
R803 B.n419 B.n418 585
R804 B.n420 B.n49 585
R805 B.n422 B.n421 585
R806 B.n423 B.n48 585
R807 B.n425 B.n424 585
R808 B.n426 B.n47 585
R809 B.n428 B.n427 585
R810 B.n429 B.n46 585
R811 B.n431 B.n430 585
R812 B.n432 B.n45 585
R813 B.n434 B.n433 585
R814 B.n435 B.n44 585
R815 B.n437 B.n436 585
R816 B.n438 B.n43 585
R817 B.n440 B.n439 585
R818 B.n442 B.n441 585
R819 B.n443 B.n39 585
R820 B.n445 B.n444 585
R821 B.n446 B.n38 585
R822 B.n448 B.n447 585
R823 B.n449 B.n37 585
R824 B.n451 B.n450 585
R825 B.n452 B.n36 585
R826 B.n454 B.n453 585
R827 B.n455 B.n33 585
R828 B.n458 B.n457 585
R829 B.n459 B.n32 585
R830 B.n461 B.n460 585
R831 B.n462 B.n31 585
R832 B.n464 B.n463 585
R833 B.n465 B.n30 585
R834 B.n467 B.n466 585
R835 B.n468 B.n29 585
R836 B.n470 B.n469 585
R837 B.n471 B.n28 585
R838 B.n473 B.n472 585
R839 B.n474 B.n27 585
R840 B.n476 B.n475 585
R841 B.n477 B.n26 585
R842 B.n479 B.n478 585
R843 B.n480 B.n25 585
R844 B.n482 B.n481 585
R845 B.n483 B.n24 585
R846 B.n485 B.n484 585
R847 B.n486 B.n23 585
R848 B.n488 B.n487 585
R849 B.n489 B.n22 585
R850 B.n491 B.n490 585
R851 B.n492 B.n21 585
R852 B.n494 B.n493 585
R853 B.n495 B.n20 585
R854 B.n497 B.n496 585
R855 B.n498 B.n19 585
R856 B.n500 B.n499 585
R857 B.n501 B.n18 585
R858 B.n503 B.n502 585
R859 B.n504 B.n17 585
R860 B.n506 B.n505 585
R861 B.n507 B.n16 585
R862 B.n509 B.n508 585
R863 B.n510 B.n15 585
R864 B.n512 B.n511 585
R865 B.n513 B.n14 585
R866 B.n515 B.n514 585
R867 B.n516 B.n13 585
R868 B.n380 B.n379 585
R869 B.n378 B.n63 585
R870 B.n377 B.n376 585
R871 B.n375 B.n64 585
R872 B.n374 B.n373 585
R873 B.n372 B.n65 585
R874 B.n371 B.n370 585
R875 B.n369 B.n66 585
R876 B.n368 B.n367 585
R877 B.n366 B.n67 585
R878 B.n365 B.n364 585
R879 B.n363 B.n68 585
R880 B.n362 B.n361 585
R881 B.n360 B.n69 585
R882 B.n359 B.n358 585
R883 B.n357 B.n70 585
R884 B.n356 B.n355 585
R885 B.n354 B.n71 585
R886 B.n353 B.n352 585
R887 B.n351 B.n72 585
R888 B.n350 B.n349 585
R889 B.n348 B.n73 585
R890 B.n347 B.n346 585
R891 B.n345 B.n74 585
R892 B.n344 B.n343 585
R893 B.n342 B.n75 585
R894 B.n341 B.n340 585
R895 B.n339 B.n76 585
R896 B.n338 B.n337 585
R897 B.n336 B.n77 585
R898 B.n335 B.n334 585
R899 B.n333 B.n78 585
R900 B.n332 B.n331 585
R901 B.n330 B.n79 585
R902 B.n329 B.n328 585
R903 B.n327 B.n80 585
R904 B.n326 B.n325 585
R905 B.n324 B.n81 585
R906 B.n323 B.n322 585
R907 B.n321 B.n82 585
R908 B.n320 B.n319 585
R909 B.n318 B.n83 585
R910 B.n317 B.n316 585
R911 B.n315 B.n84 585
R912 B.n314 B.n313 585
R913 B.n177 B.n134 585
R914 B.n179 B.n178 585
R915 B.n180 B.n133 585
R916 B.n182 B.n181 585
R917 B.n183 B.n132 585
R918 B.n185 B.n184 585
R919 B.n186 B.n131 585
R920 B.n188 B.n187 585
R921 B.n189 B.n130 585
R922 B.n191 B.n190 585
R923 B.n192 B.n129 585
R924 B.n194 B.n193 585
R925 B.n195 B.n128 585
R926 B.n197 B.n196 585
R927 B.n198 B.n127 585
R928 B.n200 B.n199 585
R929 B.n201 B.n126 585
R930 B.n203 B.n202 585
R931 B.n204 B.n125 585
R932 B.n206 B.n205 585
R933 B.n207 B.n124 585
R934 B.n209 B.n208 585
R935 B.n210 B.n123 585
R936 B.n212 B.n211 585
R937 B.n213 B.n122 585
R938 B.n215 B.n214 585
R939 B.n216 B.n121 585
R940 B.n218 B.n217 585
R941 B.n219 B.n120 585
R942 B.n221 B.n220 585
R943 B.n222 B.n119 585
R944 B.n224 B.n223 585
R945 B.n225 B.n118 585
R946 B.n227 B.n226 585
R947 B.n228 B.n117 585
R948 B.n230 B.n229 585
R949 B.n231 B.n116 585
R950 B.n233 B.n232 585
R951 B.n234 B.n115 585
R952 B.n236 B.n235 585
R953 B.n238 B.n237 585
R954 B.n239 B.n111 585
R955 B.n241 B.n240 585
R956 B.n242 B.n110 585
R957 B.n244 B.n243 585
R958 B.n245 B.n109 585
R959 B.n247 B.n246 585
R960 B.n248 B.n108 585
R961 B.n250 B.n249 585
R962 B.n251 B.n105 585
R963 B.n254 B.n253 585
R964 B.n255 B.n104 585
R965 B.n257 B.n256 585
R966 B.n258 B.n103 585
R967 B.n260 B.n259 585
R968 B.n261 B.n102 585
R969 B.n263 B.n262 585
R970 B.n264 B.n101 585
R971 B.n266 B.n265 585
R972 B.n267 B.n100 585
R973 B.n269 B.n268 585
R974 B.n270 B.n99 585
R975 B.n272 B.n271 585
R976 B.n273 B.n98 585
R977 B.n275 B.n274 585
R978 B.n276 B.n97 585
R979 B.n278 B.n277 585
R980 B.n279 B.n96 585
R981 B.n281 B.n280 585
R982 B.n282 B.n95 585
R983 B.n284 B.n283 585
R984 B.n285 B.n94 585
R985 B.n287 B.n286 585
R986 B.n288 B.n93 585
R987 B.n290 B.n289 585
R988 B.n291 B.n92 585
R989 B.n293 B.n292 585
R990 B.n294 B.n91 585
R991 B.n296 B.n295 585
R992 B.n297 B.n90 585
R993 B.n299 B.n298 585
R994 B.n300 B.n89 585
R995 B.n302 B.n301 585
R996 B.n303 B.n88 585
R997 B.n305 B.n304 585
R998 B.n306 B.n87 585
R999 B.n308 B.n307 585
R1000 B.n309 B.n86 585
R1001 B.n311 B.n310 585
R1002 B.n312 B.n85 585
R1003 B.n176 B.n175 585
R1004 B.n174 B.n135 585
R1005 B.n173 B.n172 585
R1006 B.n171 B.n136 585
R1007 B.n170 B.n169 585
R1008 B.n168 B.n137 585
R1009 B.n167 B.n166 585
R1010 B.n165 B.n138 585
R1011 B.n164 B.n163 585
R1012 B.n162 B.n139 585
R1013 B.n161 B.n160 585
R1014 B.n159 B.n140 585
R1015 B.n158 B.n157 585
R1016 B.n156 B.n141 585
R1017 B.n155 B.n154 585
R1018 B.n153 B.n142 585
R1019 B.n152 B.n151 585
R1020 B.n150 B.n143 585
R1021 B.n149 B.n148 585
R1022 B.n147 B.n144 585
R1023 B.n146 B.n145 585
R1024 B.n2 B.n0 585
R1025 B.n549 B.n1 585
R1026 B.n548 B.n547 585
R1027 B.n546 B.n3 585
R1028 B.n545 B.n544 585
R1029 B.n543 B.n4 585
R1030 B.n542 B.n541 585
R1031 B.n540 B.n5 585
R1032 B.n539 B.n538 585
R1033 B.n537 B.n6 585
R1034 B.n536 B.n535 585
R1035 B.n534 B.n7 585
R1036 B.n533 B.n532 585
R1037 B.n531 B.n8 585
R1038 B.n530 B.n529 585
R1039 B.n528 B.n9 585
R1040 B.n527 B.n526 585
R1041 B.n525 B.n10 585
R1042 B.n524 B.n523 585
R1043 B.n522 B.n11 585
R1044 B.n521 B.n520 585
R1045 B.n519 B.n12 585
R1046 B.n518 B.n517 585
R1047 B.n551 B.n550 585
R1048 B.n177 B.n176 502.111
R1049 B.n518 B.n13 502.111
R1050 B.n314 B.n85 502.111
R1051 B.n381 B.n380 502.111
R1052 B.n106 B.t3 428.606
R1053 B.n112 B.t9 428.606
R1054 B.n34 B.t0 428.606
R1055 B.n40 B.t6 428.606
R1056 B.n106 B.t5 398
R1057 B.n40 B.t7 398
R1058 B.n112 B.t11 398
R1059 B.n34 B.t1 398
R1060 B.n107 B.t4 367.551
R1061 B.n41 B.t8 367.551
R1062 B.n113 B.t10 367.55
R1063 B.n35 B.t2 367.55
R1064 B.n176 B.n135 163.367
R1065 B.n172 B.n135 163.367
R1066 B.n172 B.n171 163.367
R1067 B.n171 B.n170 163.367
R1068 B.n170 B.n137 163.367
R1069 B.n166 B.n137 163.367
R1070 B.n166 B.n165 163.367
R1071 B.n165 B.n164 163.367
R1072 B.n164 B.n139 163.367
R1073 B.n160 B.n139 163.367
R1074 B.n160 B.n159 163.367
R1075 B.n159 B.n158 163.367
R1076 B.n158 B.n141 163.367
R1077 B.n154 B.n141 163.367
R1078 B.n154 B.n153 163.367
R1079 B.n153 B.n152 163.367
R1080 B.n152 B.n143 163.367
R1081 B.n148 B.n143 163.367
R1082 B.n148 B.n147 163.367
R1083 B.n147 B.n146 163.367
R1084 B.n146 B.n2 163.367
R1085 B.n550 B.n2 163.367
R1086 B.n550 B.n549 163.367
R1087 B.n549 B.n548 163.367
R1088 B.n548 B.n3 163.367
R1089 B.n544 B.n3 163.367
R1090 B.n544 B.n543 163.367
R1091 B.n543 B.n542 163.367
R1092 B.n542 B.n5 163.367
R1093 B.n538 B.n5 163.367
R1094 B.n538 B.n537 163.367
R1095 B.n537 B.n536 163.367
R1096 B.n536 B.n7 163.367
R1097 B.n532 B.n7 163.367
R1098 B.n532 B.n531 163.367
R1099 B.n531 B.n530 163.367
R1100 B.n530 B.n9 163.367
R1101 B.n526 B.n9 163.367
R1102 B.n526 B.n525 163.367
R1103 B.n525 B.n524 163.367
R1104 B.n524 B.n11 163.367
R1105 B.n520 B.n11 163.367
R1106 B.n520 B.n519 163.367
R1107 B.n519 B.n518 163.367
R1108 B.n178 B.n177 163.367
R1109 B.n178 B.n133 163.367
R1110 B.n182 B.n133 163.367
R1111 B.n183 B.n182 163.367
R1112 B.n184 B.n183 163.367
R1113 B.n184 B.n131 163.367
R1114 B.n188 B.n131 163.367
R1115 B.n189 B.n188 163.367
R1116 B.n190 B.n189 163.367
R1117 B.n190 B.n129 163.367
R1118 B.n194 B.n129 163.367
R1119 B.n195 B.n194 163.367
R1120 B.n196 B.n195 163.367
R1121 B.n196 B.n127 163.367
R1122 B.n200 B.n127 163.367
R1123 B.n201 B.n200 163.367
R1124 B.n202 B.n201 163.367
R1125 B.n202 B.n125 163.367
R1126 B.n206 B.n125 163.367
R1127 B.n207 B.n206 163.367
R1128 B.n208 B.n207 163.367
R1129 B.n208 B.n123 163.367
R1130 B.n212 B.n123 163.367
R1131 B.n213 B.n212 163.367
R1132 B.n214 B.n213 163.367
R1133 B.n214 B.n121 163.367
R1134 B.n218 B.n121 163.367
R1135 B.n219 B.n218 163.367
R1136 B.n220 B.n219 163.367
R1137 B.n220 B.n119 163.367
R1138 B.n224 B.n119 163.367
R1139 B.n225 B.n224 163.367
R1140 B.n226 B.n225 163.367
R1141 B.n226 B.n117 163.367
R1142 B.n230 B.n117 163.367
R1143 B.n231 B.n230 163.367
R1144 B.n232 B.n231 163.367
R1145 B.n232 B.n115 163.367
R1146 B.n236 B.n115 163.367
R1147 B.n237 B.n236 163.367
R1148 B.n237 B.n111 163.367
R1149 B.n241 B.n111 163.367
R1150 B.n242 B.n241 163.367
R1151 B.n243 B.n242 163.367
R1152 B.n243 B.n109 163.367
R1153 B.n247 B.n109 163.367
R1154 B.n248 B.n247 163.367
R1155 B.n249 B.n248 163.367
R1156 B.n249 B.n105 163.367
R1157 B.n254 B.n105 163.367
R1158 B.n255 B.n254 163.367
R1159 B.n256 B.n255 163.367
R1160 B.n256 B.n103 163.367
R1161 B.n260 B.n103 163.367
R1162 B.n261 B.n260 163.367
R1163 B.n262 B.n261 163.367
R1164 B.n262 B.n101 163.367
R1165 B.n266 B.n101 163.367
R1166 B.n267 B.n266 163.367
R1167 B.n268 B.n267 163.367
R1168 B.n268 B.n99 163.367
R1169 B.n272 B.n99 163.367
R1170 B.n273 B.n272 163.367
R1171 B.n274 B.n273 163.367
R1172 B.n274 B.n97 163.367
R1173 B.n278 B.n97 163.367
R1174 B.n279 B.n278 163.367
R1175 B.n280 B.n279 163.367
R1176 B.n280 B.n95 163.367
R1177 B.n284 B.n95 163.367
R1178 B.n285 B.n284 163.367
R1179 B.n286 B.n285 163.367
R1180 B.n286 B.n93 163.367
R1181 B.n290 B.n93 163.367
R1182 B.n291 B.n290 163.367
R1183 B.n292 B.n291 163.367
R1184 B.n292 B.n91 163.367
R1185 B.n296 B.n91 163.367
R1186 B.n297 B.n296 163.367
R1187 B.n298 B.n297 163.367
R1188 B.n298 B.n89 163.367
R1189 B.n302 B.n89 163.367
R1190 B.n303 B.n302 163.367
R1191 B.n304 B.n303 163.367
R1192 B.n304 B.n87 163.367
R1193 B.n308 B.n87 163.367
R1194 B.n309 B.n308 163.367
R1195 B.n310 B.n309 163.367
R1196 B.n310 B.n85 163.367
R1197 B.n315 B.n314 163.367
R1198 B.n316 B.n315 163.367
R1199 B.n316 B.n83 163.367
R1200 B.n320 B.n83 163.367
R1201 B.n321 B.n320 163.367
R1202 B.n322 B.n321 163.367
R1203 B.n322 B.n81 163.367
R1204 B.n326 B.n81 163.367
R1205 B.n327 B.n326 163.367
R1206 B.n328 B.n327 163.367
R1207 B.n328 B.n79 163.367
R1208 B.n332 B.n79 163.367
R1209 B.n333 B.n332 163.367
R1210 B.n334 B.n333 163.367
R1211 B.n334 B.n77 163.367
R1212 B.n338 B.n77 163.367
R1213 B.n339 B.n338 163.367
R1214 B.n340 B.n339 163.367
R1215 B.n340 B.n75 163.367
R1216 B.n344 B.n75 163.367
R1217 B.n345 B.n344 163.367
R1218 B.n346 B.n345 163.367
R1219 B.n346 B.n73 163.367
R1220 B.n350 B.n73 163.367
R1221 B.n351 B.n350 163.367
R1222 B.n352 B.n351 163.367
R1223 B.n352 B.n71 163.367
R1224 B.n356 B.n71 163.367
R1225 B.n357 B.n356 163.367
R1226 B.n358 B.n357 163.367
R1227 B.n358 B.n69 163.367
R1228 B.n362 B.n69 163.367
R1229 B.n363 B.n362 163.367
R1230 B.n364 B.n363 163.367
R1231 B.n364 B.n67 163.367
R1232 B.n368 B.n67 163.367
R1233 B.n369 B.n368 163.367
R1234 B.n370 B.n369 163.367
R1235 B.n370 B.n65 163.367
R1236 B.n374 B.n65 163.367
R1237 B.n375 B.n374 163.367
R1238 B.n376 B.n375 163.367
R1239 B.n376 B.n63 163.367
R1240 B.n380 B.n63 163.367
R1241 B.n514 B.n13 163.367
R1242 B.n514 B.n513 163.367
R1243 B.n513 B.n512 163.367
R1244 B.n512 B.n15 163.367
R1245 B.n508 B.n15 163.367
R1246 B.n508 B.n507 163.367
R1247 B.n507 B.n506 163.367
R1248 B.n506 B.n17 163.367
R1249 B.n502 B.n17 163.367
R1250 B.n502 B.n501 163.367
R1251 B.n501 B.n500 163.367
R1252 B.n500 B.n19 163.367
R1253 B.n496 B.n19 163.367
R1254 B.n496 B.n495 163.367
R1255 B.n495 B.n494 163.367
R1256 B.n494 B.n21 163.367
R1257 B.n490 B.n21 163.367
R1258 B.n490 B.n489 163.367
R1259 B.n489 B.n488 163.367
R1260 B.n488 B.n23 163.367
R1261 B.n484 B.n23 163.367
R1262 B.n484 B.n483 163.367
R1263 B.n483 B.n482 163.367
R1264 B.n482 B.n25 163.367
R1265 B.n478 B.n25 163.367
R1266 B.n478 B.n477 163.367
R1267 B.n477 B.n476 163.367
R1268 B.n476 B.n27 163.367
R1269 B.n472 B.n27 163.367
R1270 B.n472 B.n471 163.367
R1271 B.n471 B.n470 163.367
R1272 B.n470 B.n29 163.367
R1273 B.n466 B.n29 163.367
R1274 B.n466 B.n465 163.367
R1275 B.n465 B.n464 163.367
R1276 B.n464 B.n31 163.367
R1277 B.n460 B.n31 163.367
R1278 B.n460 B.n459 163.367
R1279 B.n459 B.n458 163.367
R1280 B.n458 B.n33 163.367
R1281 B.n453 B.n33 163.367
R1282 B.n453 B.n452 163.367
R1283 B.n452 B.n451 163.367
R1284 B.n451 B.n37 163.367
R1285 B.n447 B.n37 163.367
R1286 B.n447 B.n446 163.367
R1287 B.n446 B.n445 163.367
R1288 B.n445 B.n39 163.367
R1289 B.n441 B.n39 163.367
R1290 B.n441 B.n440 163.367
R1291 B.n440 B.n43 163.367
R1292 B.n436 B.n43 163.367
R1293 B.n436 B.n435 163.367
R1294 B.n435 B.n434 163.367
R1295 B.n434 B.n45 163.367
R1296 B.n430 B.n45 163.367
R1297 B.n430 B.n429 163.367
R1298 B.n429 B.n428 163.367
R1299 B.n428 B.n47 163.367
R1300 B.n424 B.n47 163.367
R1301 B.n424 B.n423 163.367
R1302 B.n423 B.n422 163.367
R1303 B.n422 B.n49 163.367
R1304 B.n418 B.n49 163.367
R1305 B.n418 B.n417 163.367
R1306 B.n417 B.n416 163.367
R1307 B.n416 B.n51 163.367
R1308 B.n412 B.n51 163.367
R1309 B.n412 B.n411 163.367
R1310 B.n411 B.n410 163.367
R1311 B.n410 B.n53 163.367
R1312 B.n406 B.n53 163.367
R1313 B.n406 B.n405 163.367
R1314 B.n405 B.n404 163.367
R1315 B.n404 B.n55 163.367
R1316 B.n400 B.n55 163.367
R1317 B.n400 B.n399 163.367
R1318 B.n399 B.n398 163.367
R1319 B.n398 B.n57 163.367
R1320 B.n394 B.n57 163.367
R1321 B.n394 B.n393 163.367
R1322 B.n393 B.n392 163.367
R1323 B.n392 B.n59 163.367
R1324 B.n388 B.n59 163.367
R1325 B.n388 B.n387 163.367
R1326 B.n387 B.n386 163.367
R1327 B.n386 B.n61 163.367
R1328 B.n382 B.n61 163.367
R1329 B.n382 B.n381 163.367
R1330 B.n252 B.n107 59.5399
R1331 B.n114 B.n113 59.5399
R1332 B.n456 B.n35 59.5399
R1333 B.n42 B.n41 59.5399
R1334 B.n517 B.n516 32.6249
R1335 B.n379 B.n62 32.6249
R1336 B.n313 B.n312 32.6249
R1337 B.n175 B.n134 32.6249
R1338 B.n107 B.n106 30.449
R1339 B.n113 B.n112 30.449
R1340 B.n35 B.n34 30.449
R1341 B.n41 B.n40 30.449
R1342 B B.n551 18.0485
R1343 B.n516 B.n515 10.6151
R1344 B.n515 B.n14 10.6151
R1345 B.n511 B.n14 10.6151
R1346 B.n511 B.n510 10.6151
R1347 B.n510 B.n509 10.6151
R1348 B.n509 B.n16 10.6151
R1349 B.n505 B.n16 10.6151
R1350 B.n505 B.n504 10.6151
R1351 B.n504 B.n503 10.6151
R1352 B.n503 B.n18 10.6151
R1353 B.n499 B.n18 10.6151
R1354 B.n499 B.n498 10.6151
R1355 B.n498 B.n497 10.6151
R1356 B.n497 B.n20 10.6151
R1357 B.n493 B.n20 10.6151
R1358 B.n493 B.n492 10.6151
R1359 B.n492 B.n491 10.6151
R1360 B.n491 B.n22 10.6151
R1361 B.n487 B.n22 10.6151
R1362 B.n487 B.n486 10.6151
R1363 B.n486 B.n485 10.6151
R1364 B.n485 B.n24 10.6151
R1365 B.n481 B.n24 10.6151
R1366 B.n481 B.n480 10.6151
R1367 B.n480 B.n479 10.6151
R1368 B.n479 B.n26 10.6151
R1369 B.n475 B.n26 10.6151
R1370 B.n475 B.n474 10.6151
R1371 B.n474 B.n473 10.6151
R1372 B.n473 B.n28 10.6151
R1373 B.n469 B.n28 10.6151
R1374 B.n469 B.n468 10.6151
R1375 B.n468 B.n467 10.6151
R1376 B.n467 B.n30 10.6151
R1377 B.n463 B.n30 10.6151
R1378 B.n463 B.n462 10.6151
R1379 B.n462 B.n461 10.6151
R1380 B.n461 B.n32 10.6151
R1381 B.n457 B.n32 10.6151
R1382 B.n455 B.n454 10.6151
R1383 B.n454 B.n36 10.6151
R1384 B.n450 B.n36 10.6151
R1385 B.n450 B.n449 10.6151
R1386 B.n449 B.n448 10.6151
R1387 B.n448 B.n38 10.6151
R1388 B.n444 B.n38 10.6151
R1389 B.n444 B.n443 10.6151
R1390 B.n443 B.n442 10.6151
R1391 B.n439 B.n438 10.6151
R1392 B.n438 B.n437 10.6151
R1393 B.n437 B.n44 10.6151
R1394 B.n433 B.n44 10.6151
R1395 B.n433 B.n432 10.6151
R1396 B.n432 B.n431 10.6151
R1397 B.n431 B.n46 10.6151
R1398 B.n427 B.n46 10.6151
R1399 B.n427 B.n426 10.6151
R1400 B.n426 B.n425 10.6151
R1401 B.n425 B.n48 10.6151
R1402 B.n421 B.n48 10.6151
R1403 B.n421 B.n420 10.6151
R1404 B.n420 B.n419 10.6151
R1405 B.n419 B.n50 10.6151
R1406 B.n415 B.n50 10.6151
R1407 B.n415 B.n414 10.6151
R1408 B.n414 B.n413 10.6151
R1409 B.n413 B.n52 10.6151
R1410 B.n409 B.n52 10.6151
R1411 B.n409 B.n408 10.6151
R1412 B.n408 B.n407 10.6151
R1413 B.n407 B.n54 10.6151
R1414 B.n403 B.n54 10.6151
R1415 B.n403 B.n402 10.6151
R1416 B.n402 B.n401 10.6151
R1417 B.n401 B.n56 10.6151
R1418 B.n397 B.n56 10.6151
R1419 B.n397 B.n396 10.6151
R1420 B.n396 B.n395 10.6151
R1421 B.n395 B.n58 10.6151
R1422 B.n391 B.n58 10.6151
R1423 B.n391 B.n390 10.6151
R1424 B.n390 B.n389 10.6151
R1425 B.n389 B.n60 10.6151
R1426 B.n385 B.n60 10.6151
R1427 B.n385 B.n384 10.6151
R1428 B.n384 B.n383 10.6151
R1429 B.n383 B.n62 10.6151
R1430 B.n313 B.n84 10.6151
R1431 B.n317 B.n84 10.6151
R1432 B.n318 B.n317 10.6151
R1433 B.n319 B.n318 10.6151
R1434 B.n319 B.n82 10.6151
R1435 B.n323 B.n82 10.6151
R1436 B.n324 B.n323 10.6151
R1437 B.n325 B.n324 10.6151
R1438 B.n325 B.n80 10.6151
R1439 B.n329 B.n80 10.6151
R1440 B.n330 B.n329 10.6151
R1441 B.n331 B.n330 10.6151
R1442 B.n331 B.n78 10.6151
R1443 B.n335 B.n78 10.6151
R1444 B.n336 B.n335 10.6151
R1445 B.n337 B.n336 10.6151
R1446 B.n337 B.n76 10.6151
R1447 B.n341 B.n76 10.6151
R1448 B.n342 B.n341 10.6151
R1449 B.n343 B.n342 10.6151
R1450 B.n343 B.n74 10.6151
R1451 B.n347 B.n74 10.6151
R1452 B.n348 B.n347 10.6151
R1453 B.n349 B.n348 10.6151
R1454 B.n349 B.n72 10.6151
R1455 B.n353 B.n72 10.6151
R1456 B.n354 B.n353 10.6151
R1457 B.n355 B.n354 10.6151
R1458 B.n355 B.n70 10.6151
R1459 B.n359 B.n70 10.6151
R1460 B.n360 B.n359 10.6151
R1461 B.n361 B.n360 10.6151
R1462 B.n361 B.n68 10.6151
R1463 B.n365 B.n68 10.6151
R1464 B.n366 B.n365 10.6151
R1465 B.n367 B.n366 10.6151
R1466 B.n367 B.n66 10.6151
R1467 B.n371 B.n66 10.6151
R1468 B.n372 B.n371 10.6151
R1469 B.n373 B.n372 10.6151
R1470 B.n373 B.n64 10.6151
R1471 B.n377 B.n64 10.6151
R1472 B.n378 B.n377 10.6151
R1473 B.n379 B.n378 10.6151
R1474 B.n179 B.n134 10.6151
R1475 B.n180 B.n179 10.6151
R1476 B.n181 B.n180 10.6151
R1477 B.n181 B.n132 10.6151
R1478 B.n185 B.n132 10.6151
R1479 B.n186 B.n185 10.6151
R1480 B.n187 B.n186 10.6151
R1481 B.n187 B.n130 10.6151
R1482 B.n191 B.n130 10.6151
R1483 B.n192 B.n191 10.6151
R1484 B.n193 B.n192 10.6151
R1485 B.n193 B.n128 10.6151
R1486 B.n197 B.n128 10.6151
R1487 B.n198 B.n197 10.6151
R1488 B.n199 B.n198 10.6151
R1489 B.n199 B.n126 10.6151
R1490 B.n203 B.n126 10.6151
R1491 B.n204 B.n203 10.6151
R1492 B.n205 B.n204 10.6151
R1493 B.n205 B.n124 10.6151
R1494 B.n209 B.n124 10.6151
R1495 B.n210 B.n209 10.6151
R1496 B.n211 B.n210 10.6151
R1497 B.n211 B.n122 10.6151
R1498 B.n215 B.n122 10.6151
R1499 B.n216 B.n215 10.6151
R1500 B.n217 B.n216 10.6151
R1501 B.n217 B.n120 10.6151
R1502 B.n221 B.n120 10.6151
R1503 B.n222 B.n221 10.6151
R1504 B.n223 B.n222 10.6151
R1505 B.n223 B.n118 10.6151
R1506 B.n227 B.n118 10.6151
R1507 B.n228 B.n227 10.6151
R1508 B.n229 B.n228 10.6151
R1509 B.n229 B.n116 10.6151
R1510 B.n233 B.n116 10.6151
R1511 B.n234 B.n233 10.6151
R1512 B.n235 B.n234 10.6151
R1513 B.n239 B.n238 10.6151
R1514 B.n240 B.n239 10.6151
R1515 B.n240 B.n110 10.6151
R1516 B.n244 B.n110 10.6151
R1517 B.n245 B.n244 10.6151
R1518 B.n246 B.n245 10.6151
R1519 B.n246 B.n108 10.6151
R1520 B.n250 B.n108 10.6151
R1521 B.n251 B.n250 10.6151
R1522 B.n253 B.n104 10.6151
R1523 B.n257 B.n104 10.6151
R1524 B.n258 B.n257 10.6151
R1525 B.n259 B.n258 10.6151
R1526 B.n259 B.n102 10.6151
R1527 B.n263 B.n102 10.6151
R1528 B.n264 B.n263 10.6151
R1529 B.n265 B.n264 10.6151
R1530 B.n265 B.n100 10.6151
R1531 B.n269 B.n100 10.6151
R1532 B.n270 B.n269 10.6151
R1533 B.n271 B.n270 10.6151
R1534 B.n271 B.n98 10.6151
R1535 B.n275 B.n98 10.6151
R1536 B.n276 B.n275 10.6151
R1537 B.n277 B.n276 10.6151
R1538 B.n277 B.n96 10.6151
R1539 B.n281 B.n96 10.6151
R1540 B.n282 B.n281 10.6151
R1541 B.n283 B.n282 10.6151
R1542 B.n283 B.n94 10.6151
R1543 B.n287 B.n94 10.6151
R1544 B.n288 B.n287 10.6151
R1545 B.n289 B.n288 10.6151
R1546 B.n289 B.n92 10.6151
R1547 B.n293 B.n92 10.6151
R1548 B.n294 B.n293 10.6151
R1549 B.n295 B.n294 10.6151
R1550 B.n295 B.n90 10.6151
R1551 B.n299 B.n90 10.6151
R1552 B.n300 B.n299 10.6151
R1553 B.n301 B.n300 10.6151
R1554 B.n301 B.n88 10.6151
R1555 B.n305 B.n88 10.6151
R1556 B.n306 B.n305 10.6151
R1557 B.n307 B.n306 10.6151
R1558 B.n307 B.n86 10.6151
R1559 B.n311 B.n86 10.6151
R1560 B.n312 B.n311 10.6151
R1561 B.n175 B.n174 10.6151
R1562 B.n174 B.n173 10.6151
R1563 B.n173 B.n136 10.6151
R1564 B.n169 B.n136 10.6151
R1565 B.n169 B.n168 10.6151
R1566 B.n168 B.n167 10.6151
R1567 B.n167 B.n138 10.6151
R1568 B.n163 B.n138 10.6151
R1569 B.n163 B.n162 10.6151
R1570 B.n162 B.n161 10.6151
R1571 B.n161 B.n140 10.6151
R1572 B.n157 B.n140 10.6151
R1573 B.n157 B.n156 10.6151
R1574 B.n156 B.n155 10.6151
R1575 B.n155 B.n142 10.6151
R1576 B.n151 B.n142 10.6151
R1577 B.n151 B.n150 10.6151
R1578 B.n150 B.n149 10.6151
R1579 B.n149 B.n144 10.6151
R1580 B.n145 B.n144 10.6151
R1581 B.n145 B.n0 10.6151
R1582 B.n547 B.n1 10.6151
R1583 B.n547 B.n546 10.6151
R1584 B.n546 B.n545 10.6151
R1585 B.n545 B.n4 10.6151
R1586 B.n541 B.n4 10.6151
R1587 B.n541 B.n540 10.6151
R1588 B.n540 B.n539 10.6151
R1589 B.n539 B.n6 10.6151
R1590 B.n535 B.n6 10.6151
R1591 B.n535 B.n534 10.6151
R1592 B.n534 B.n533 10.6151
R1593 B.n533 B.n8 10.6151
R1594 B.n529 B.n8 10.6151
R1595 B.n529 B.n528 10.6151
R1596 B.n528 B.n527 10.6151
R1597 B.n527 B.n10 10.6151
R1598 B.n523 B.n10 10.6151
R1599 B.n523 B.n522 10.6151
R1600 B.n522 B.n521 10.6151
R1601 B.n521 B.n12 10.6151
R1602 B.n517 B.n12 10.6151
R1603 B.n457 B.n456 9.36635
R1604 B.n439 B.n42 9.36635
R1605 B.n235 B.n114 9.36635
R1606 B.n253 B.n252 9.36635
R1607 B.n551 B.n0 2.81026
R1608 B.n551 B.n1 2.81026
R1609 B.n456 B.n455 1.24928
R1610 B.n442 B.n42 1.24928
R1611 B.n238 B.n114 1.24928
R1612 B.n252 B.n251 1.24928
R1613 VN.n0 VN.t1 260.993
R1614 VN.n1 VN.t0 260.993
R1615 VN.n0 VN.t2 260.772
R1616 VN.n1 VN.t3 260.772
R1617 VN VN.n1 60.3386
R1618 VN VN.n0 18.2817
R1619 VDD2.n2 VDD2.n0 115.222
R1620 VDD2.n2 VDD2.n1 77.498
R1621 VDD2.n1 VDD2.t0 2.81722
R1622 VDD2.n1 VDD2.t3 2.81722
R1623 VDD2.n0 VDD2.t2 2.81722
R1624 VDD2.n0 VDD2.t1 2.81722
R1625 VDD2 VDD2.n2 0.0586897
C0 VN VDD1 0.147918f
C1 VP w_n1912_n3276# 3.22316f
C2 B w_n1912_n3276# 7.44286f
C3 VDD2 w_n1912_n3276# 1.19225f
C4 VP VTAIL 3.54154f
C5 VTAIL B 4.07514f
C6 VDD2 VTAIL 5.62573f
C7 VN VP 5.12403f
C8 VP VDD1 3.97204f
C9 VN B 0.847592f
C10 VDD1 B 1.00953f
C11 VN VDD2 3.81244f
C12 VDD2 VDD1 0.694072f
C13 VTAIL w_n1912_n3276# 3.93405f
C14 VN w_n1912_n3276# 2.98081f
C15 VDD1 w_n1912_n3276# 1.16631f
C16 VP B 1.24344f
C17 VDD2 VP 0.307914f
C18 VDD2 B 1.03952f
C19 VN VTAIL 3.52743f
C20 VDD1 VTAIL 5.58064f
C21 VDD2 VSUBS 0.73354f
C22 VDD1 VSUBS 5.006402f
C23 VTAIL VSUBS 0.958353f
C24 VN VSUBS 5.18972f
C25 VP VSUBS 1.546229f
C26 B VSUBS 3.054572f
C27 w_n1912_n3276# VSUBS 77.160706f
C28 VDD2.t2 VSUBS 0.244441f
C29 VDD2.t1 VSUBS 0.244441f
C30 VDD2.n0 VSUBS 2.49994f
C31 VDD2.t0 VSUBS 0.244441f
C32 VDD2.t3 VSUBS 0.244441f
C33 VDD2.n1 VSUBS 1.90374f
C34 VDD2.n2 VSUBS 3.89589f
C35 VN.t1 VSUBS 1.98821f
C36 VN.t2 VSUBS 1.98746f
C37 VN.n0 VSUBS 1.50033f
C38 VN.t0 VSUBS 1.98821f
C39 VN.t3 VSUBS 1.98746f
C40 VN.n1 VSUBS 3.03616f
C41 B.n0 VSUBS 0.004882f
C42 B.n1 VSUBS 0.004882f
C43 B.n2 VSUBS 0.007721f
C44 B.n3 VSUBS 0.007721f
C45 B.n4 VSUBS 0.007721f
C46 B.n5 VSUBS 0.007721f
C47 B.n6 VSUBS 0.007721f
C48 B.n7 VSUBS 0.007721f
C49 B.n8 VSUBS 0.007721f
C50 B.n9 VSUBS 0.007721f
C51 B.n10 VSUBS 0.007721f
C52 B.n11 VSUBS 0.007721f
C53 B.n12 VSUBS 0.007721f
C54 B.n13 VSUBS 0.018421f
C55 B.n14 VSUBS 0.007721f
C56 B.n15 VSUBS 0.007721f
C57 B.n16 VSUBS 0.007721f
C58 B.n17 VSUBS 0.007721f
C59 B.n18 VSUBS 0.007721f
C60 B.n19 VSUBS 0.007721f
C61 B.n20 VSUBS 0.007721f
C62 B.n21 VSUBS 0.007721f
C63 B.n22 VSUBS 0.007721f
C64 B.n23 VSUBS 0.007721f
C65 B.n24 VSUBS 0.007721f
C66 B.n25 VSUBS 0.007721f
C67 B.n26 VSUBS 0.007721f
C68 B.n27 VSUBS 0.007721f
C69 B.n28 VSUBS 0.007721f
C70 B.n29 VSUBS 0.007721f
C71 B.n30 VSUBS 0.007721f
C72 B.n31 VSUBS 0.007721f
C73 B.n32 VSUBS 0.007721f
C74 B.n33 VSUBS 0.007721f
C75 B.t2 VSUBS 0.221782f
C76 B.t1 VSUBS 0.241151f
C77 B.t0 VSUBS 0.681912f
C78 B.n34 VSUBS 0.364831f
C79 B.n35 VSUBS 0.264185f
C80 B.n36 VSUBS 0.007721f
C81 B.n37 VSUBS 0.007721f
C82 B.n38 VSUBS 0.007721f
C83 B.n39 VSUBS 0.007721f
C84 B.t8 VSUBS 0.221785f
C85 B.t7 VSUBS 0.241154f
C86 B.t6 VSUBS 0.681912f
C87 B.n40 VSUBS 0.364828f
C88 B.n41 VSUBS 0.264182f
C89 B.n42 VSUBS 0.017889f
C90 B.n43 VSUBS 0.007721f
C91 B.n44 VSUBS 0.007721f
C92 B.n45 VSUBS 0.007721f
C93 B.n46 VSUBS 0.007721f
C94 B.n47 VSUBS 0.007721f
C95 B.n48 VSUBS 0.007721f
C96 B.n49 VSUBS 0.007721f
C97 B.n50 VSUBS 0.007721f
C98 B.n51 VSUBS 0.007721f
C99 B.n52 VSUBS 0.007721f
C100 B.n53 VSUBS 0.007721f
C101 B.n54 VSUBS 0.007721f
C102 B.n55 VSUBS 0.007721f
C103 B.n56 VSUBS 0.007721f
C104 B.n57 VSUBS 0.007721f
C105 B.n58 VSUBS 0.007721f
C106 B.n59 VSUBS 0.007721f
C107 B.n60 VSUBS 0.007721f
C108 B.n61 VSUBS 0.007721f
C109 B.n62 VSUBS 0.017507f
C110 B.n63 VSUBS 0.007721f
C111 B.n64 VSUBS 0.007721f
C112 B.n65 VSUBS 0.007721f
C113 B.n66 VSUBS 0.007721f
C114 B.n67 VSUBS 0.007721f
C115 B.n68 VSUBS 0.007721f
C116 B.n69 VSUBS 0.007721f
C117 B.n70 VSUBS 0.007721f
C118 B.n71 VSUBS 0.007721f
C119 B.n72 VSUBS 0.007721f
C120 B.n73 VSUBS 0.007721f
C121 B.n74 VSUBS 0.007721f
C122 B.n75 VSUBS 0.007721f
C123 B.n76 VSUBS 0.007721f
C124 B.n77 VSUBS 0.007721f
C125 B.n78 VSUBS 0.007721f
C126 B.n79 VSUBS 0.007721f
C127 B.n80 VSUBS 0.007721f
C128 B.n81 VSUBS 0.007721f
C129 B.n82 VSUBS 0.007721f
C130 B.n83 VSUBS 0.007721f
C131 B.n84 VSUBS 0.007721f
C132 B.n85 VSUBS 0.018421f
C133 B.n86 VSUBS 0.007721f
C134 B.n87 VSUBS 0.007721f
C135 B.n88 VSUBS 0.007721f
C136 B.n89 VSUBS 0.007721f
C137 B.n90 VSUBS 0.007721f
C138 B.n91 VSUBS 0.007721f
C139 B.n92 VSUBS 0.007721f
C140 B.n93 VSUBS 0.007721f
C141 B.n94 VSUBS 0.007721f
C142 B.n95 VSUBS 0.007721f
C143 B.n96 VSUBS 0.007721f
C144 B.n97 VSUBS 0.007721f
C145 B.n98 VSUBS 0.007721f
C146 B.n99 VSUBS 0.007721f
C147 B.n100 VSUBS 0.007721f
C148 B.n101 VSUBS 0.007721f
C149 B.n102 VSUBS 0.007721f
C150 B.n103 VSUBS 0.007721f
C151 B.n104 VSUBS 0.007721f
C152 B.n105 VSUBS 0.007721f
C153 B.t4 VSUBS 0.221785f
C154 B.t5 VSUBS 0.241154f
C155 B.t3 VSUBS 0.681912f
C156 B.n106 VSUBS 0.364828f
C157 B.n107 VSUBS 0.264182f
C158 B.n108 VSUBS 0.007721f
C159 B.n109 VSUBS 0.007721f
C160 B.n110 VSUBS 0.007721f
C161 B.n111 VSUBS 0.007721f
C162 B.t10 VSUBS 0.221782f
C163 B.t11 VSUBS 0.241151f
C164 B.t9 VSUBS 0.681912f
C165 B.n112 VSUBS 0.364831f
C166 B.n113 VSUBS 0.264185f
C167 B.n114 VSUBS 0.017889f
C168 B.n115 VSUBS 0.007721f
C169 B.n116 VSUBS 0.007721f
C170 B.n117 VSUBS 0.007721f
C171 B.n118 VSUBS 0.007721f
C172 B.n119 VSUBS 0.007721f
C173 B.n120 VSUBS 0.007721f
C174 B.n121 VSUBS 0.007721f
C175 B.n122 VSUBS 0.007721f
C176 B.n123 VSUBS 0.007721f
C177 B.n124 VSUBS 0.007721f
C178 B.n125 VSUBS 0.007721f
C179 B.n126 VSUBS 0.007721f
C180 B.n127 VSUBS 0.007721f
C181 B.n128 VSUBS 0.007721f
C182 B.n129 VSUBS 0.007721f
C183 B.n130 VSUBS 0.007721f
C184 B.n131 VSUBS 0.007721f
C185 B.n132 VSUBS 0.007721f
C186 B.n133 VSUBS 0.007721f
C187 B.n134 VSUBS 0.018421f
C188 B.n135 VSUBS 0.007721f
C189 B.n136 VSUBS 0.007721f
C190 B.n137 VSUBS 0.007721f
C191 B.n138 VSUBS 0.007721f
C192 B.n139 VSUBS 0.007721f
C193 B.n140 VSUBS 0.007721f
C194 B.n141 VSUBS 0.007721f
C195 B.n142 VSUBS 0.007721f
C196 B.n143 VSUBS 0.007721f
C197 B.n144 VSUBS 0.007721f
C198 B.n145 VSUBS 0.007721f
C199 B.n146 VSUBS 0.007721f
C200 B.n147 VSUBS 0.007721f
C201 B.n148 VSUBS 0.007721f
C202 B.n149 VSUBS 0.007721f
C203 B.n150 VSUBS 0.007721f
C204 B.n151 VSUBS 0.007721f
C205 B.n152 VSUBS 0.007721f
C206 B.n153 VSUBS 0.007721f
C207 B.n154 VSUBS 0.007721f
C208 B.n155 VSUBS 0.007721f
C209 B.n156 VSUBS 0.007721f
C210 B.n157 VSUBS 0.007721f
C211 B.n158 VSUBS 0.007721f
C212 B.n159 VSUBS 0.007721f
C213 B.n160 VSUBS 0.007721f
C214 B.n161 VSUBS 0.007721f
C215 B.n162 VSUBS 0.007721f
C216 B.n163 VSUBS 0.007721f
C217 B.n164 VSUBS 0.007721f
C218 B.n165 VSUBS 0.007721f
C219 B.n166 VSUBS 0.007721f
C220 B.n167 VSUBS 0.007721f
C221 B.n168 VSUBS 0.007721f
C222 B.n169 VSUBS 0.007721f
C223 B.n170 VSUBS 0.007721f
C224 B.n171 VSUBS 0.007721f
C225 B.n172 VSUBS 0.007721f
C226 B.n173 VSUBS 0.007721f
C227 B.n174 VSUBS 0.007721f
C228 B.n175 VSUBS 0.017686f
C229 B.n176 VSUBS 0.017686f
C230 B.n177 VSUBS 0.018421f
C231 B.n178 VSUBS 0.007721f
C232 B.n179 VSUBS 0.007721f
C233 B.n180 VSUBS 0.007721f
C234 B.n181 VSUBS 0.007721f
C235 B.n182 VSUBS 0.007721f
C236 B.n183 VSUBS 0.007721f
C237 B.n184 VSUBS 0.007721f
C238 B.n185 VSUBS 0.007721f
C239 B.n186 VSUBS 0.007721f
C240 B.n187 VSUBS 0.007721f
C241 B.n188 VSUBS 0.007721f
C242 B.n189 VSUBS 0.007721f
C243 B.n190 VSUBS 0.007721f
C244 B.n191 VSUBS 0.007721f
C245 B.n192 VSUBS 0.007721f
C246 B.n193 VSUBS 0.007721f
C247 B.n194 VSUBS 0.007721f
C248 B.n195 VSUBS 0.007721f
C249 B.n196 VSUBS 0.007721f
C250 B.n197 VSUBS 0.007721f
C251 B.n198 VSUBS 0.007721f
C252 B.n199 VSUBS 0.007721f
C253 B.n200 VSUBS 0.007721f
C254 B.n201 VSUBS 0.007721f
C255 B.n202 VSUBS 0.007721f
C256 B.n203 VSUBS 0.007721f
C257 B.n204 VSUBS 0.007721f
C258 B.n205 VSUBS 0.007721f
C259 B.n206 VSUBS 0.007721f
C260 B.n207 VSUBS 0.007721f
C261 B.n208 VSUBS 0.007721f
C262 B.n209 VSUBS 0.007721f
C263 B.n210 VSUBS 0.007721f
C264 B.n211 VSUBS 0.007721f
C265 B.n212 VSUBS 0.007721f
C266 B.n213 VSUBS 0.007721f
C267 B.n214 VSUBS 0.007721f
C268 B.n215 VSUBS 0.007721f
C269 B.n216 VSUBS 0.007721f
C270 B.n217 VSUBS 0.007721f
C271 B.n218 VSUBS 0.007721f
C272 B.n219 VSUBS 0.007721f
C273 B.n220 VSUBS 0.007721f
C274 B.n221 VSUBS 0.007721f
C275 B.n222 VSUBS 0.007721f
C276 B.n223 VSUBS 0.007721f
C277 B.n224 VSUBS 0.007721f
C278 B.n225 VSUBS 0.007721f
C279 B.n226 VSUBS 0.007721f
C280 B.n227 VSUBS 0.007721f
C281 B.n228 VSUBS 0.007721f
C282 B.n229 VSUBS 0.007721f
C283 B.n230 VSUBS 0.007721f
C284 B.n231 VSUBS 0.007721f
C285 B.n232 VSUBS 0.007721f
C286 B.n233 VSUBS 0.007721f
C287 B.n234 VSUBS 0.007721f
C288 B.n235 VSUBS 0.007267f
C289 B.n236 VSUBS 0.007721f
C290 B.n237 VSUBS 0.007721f
C291 B.n238 VSUBS 0.004315f
C292 B.n239 VSUBS 0.007721f
C293 B.n240 VSUBS 0.007721f
C294 B.n241 VSUBS 0.007721f
C295 B.n242 VSUBS 0.007721f
C296 B.n243 VSUBS 0.007721f
C297 B.n244 VSUBS 0.007721f
C298 B.n245 VSUBS 0.007721f
C299 B.n246 VSUBS 0.007721f
C300 B.n247 VSUBS 0.007721f
C301 B.n248 VSUBS 0.007721f
C302 B.n249 VSUBS 0.007721f
C303 B.n250 VSUBS 0.007721f
C304 B.n251 VSUBS 0.004315f
C305 B.n252 VSUBS 0.017889f
C306 B.n253 VSUBS 0.007267f
C307 B.n254 VSUBS 0.007721f
C308 B.n255 VSUBS 0.007721f
C309 B.n256 VSUBS 0.007721f
C310 B.n257 VSUBS 0.007721f
C311 B.n258 VSUBS 0.007721f
C312 B.n259 VSUBS 0.007721f
C313 B.n260 VSUBS 0.007721f
C314 B.n261 VSUBS 0.007721f
C315 B.n262 VSUBS 0.007721f
C316 B.n263 VSUBS 0.007721f
C317 B.n264 VSUBS 0.007721f
C318 B.n265 VSUBS 0.007721f
C319 B.n266 VSUBS 0.007721f
C320 B.n267 VSUBS 0.007721f
C321 B.n268 VSUBS 0.007721f
C322 B.n269 VSUBS 0.007721f
C323 B.n270 VSUBS 0.007721f
C324 B.n271 VSUBS 0.007721f
C325 B.n272 VSUBS 0.007721f
C326 B.n273 VSUBS 0.007721f
C327 B.n274 VSUBS 0.007721f
C328 B.n275 VSUBS 0.007721f
C329 B.n276 VSUBS 0.007721f
C330 B.n277 VSUBS 0.007721f
C331 B.n278 VSUBS 0.007721f
C332 B.n279 VSUBS 0.007721f
C333 B.n280 VSUBS 0.007721f
C334 B.n281 VSUBS 0.007721f
C335 B.n282 VSUBS 0.007721f
C336 B.n283 VSUBS 0.007721f
C337 B.n284 VSUBS 0.007721f
C338 B.n285 VSUBS 0.007721f
C339 B.n286 VSUBS 0.007721f
C340 B.n287 VSUBS 0.007721f
C341 B.n288 VSUBS 0.007721f
C342 B.n289 VSUBS 0.007721f
C343 B.n290 VSUBS 0.007721f
C344 B.n291 VSUBS 0.007721f
C345 B.n292 VSUBS 0.007721f
C346 B.n293 VSUBS 0.007721f
C347 B.n294 VSUBS 0.007721f
C348 B.n295 VSUBS 0.007721f
C349 B.n296 VSUBS 0.007721f
C350 B.n297 VSUBS 0.007721f
C351 B.n298 VSUBS 0.007721f
C352 B.n299 VSUBS 0.007721f
C353 B.n300 VSUBS 0.007721f
C354 B.n301 VSUBS 0.007721f
C355 B.n302 VSUBS 0.007721f
C356 B.n303 VSUBS 0.007721f
C357 B.n304 VSUBS 0.007721f
C358 B.n305 VSUBS 0.007721f
C359 B.n306 VSUBS 0.007721f
C360 B.n307 VSUBS 0.007721f
C361 B.n308 VSUBS 0.007721f
C362 B.n309 VSUBS 0.007721f
C363 B.n310 VSUBS 0.007721f
C364 B.n311 VSUBS 0.007721f
C365 B.n312 VSUBS 0.018421f
C366 B.n313 VSUBS 0.017686f
C367 B.n314 VSUBS 0.017686f
C368 B.n315 VSUBS 0.007721f
C369 B.n316 VSUBS 0.007721f
C370 B.n317 VSUBS 0.007721f
C371 B.n318 VSUBS 0.007721f
C372 B.n319 VSUBS 0.007721f
C373 B.n320 VSUBS 0.007721f
C374 B.n321 VSUBS 0.007721f
C375 B.n322 VSUBS 0.007721f
C376 B.n323 VSUBS 0.007721f
C377 B.n324 VSUBS 0.007721f
C378 B.n325 VSUBS 0.007721f
C379 B.n326 VSUBS 0.007721f
C380 B.n327 VSUBS 0.007721f
C381 B.n328 VSUBS 0.007721f
C382 B.n329 VSUBS 0.007721f
C383 B.n330 VSUBS 0.007721f
C384 B.n331 VSUBS 0.007721f
C385 B.n332 VSUBS 0.007721f
C386 B.n333 VSUBS 0.007721f
C387 B.n334 VSUBS 0.007721f
C388 B.n335 VSUBS 0.007721f
C389 B.n336 VSUBS 0.007721f
C390 B.n337 VSUBS 0.007721f
C391 B.n338 VSUBS 0.007721f
C392 B.n339 VSUBS 0.007721f
C393 B.n340 VSUBS 0.007721f
C394 B.n341 VSUBS 0.007721f
C395 B.n342 VSUBS 0.007721f
C396 B.n343 VSUBS 0.007721f
C397 B.n344 VSUBS 0.007721f
C398 B.n345 VSUBS 0.007721f
C399 B.n346 VSUBS 0.007721f
C400 B.n347 VSUBS 0.007721f
C401 B.n348 VSUBS 0.007721f
C402 B.n349 VSUBS 0.007721f
C403 B.n350 VSUBS 0.007721f
C404 B.n351 VSUBS 0.007721f
C405 B.n352 VSUBS 0.007721f
C406 B.n353 VSUBS 0.007721f
C407 B.n354 VSUBS 0.007721f
C408 B.n355 VSUBS 0.007721f
C409 B.n356 VSUBS 0.007721f
C410 B.n357 VSUBS 0.007721f
C411 B.n358 VSUBS 0.007721f
C412 B.n359 VSUBS 0.007721f
C413 B.n360 VSUBS 0.007721f
C414 B.n361 VSUBS 0.007721f
C415 B.n362 VSUBS 0.007721f
C416 B.n363 VSUBS 0.007721f
C417 B.n364 VSUBS 0.007721f
C418 B.n365 VSUBS 0.007721f
C419 B.n366 VSUBS 0.007721f
C420 B.n367 VSUBS 0.007721f
C421 B.n368 VSUBS 0.007721f
C422 B.n369 VSUBS 0.007721f
C423 B.n370 VSUBS 0.007721f
C424 B.n371 VSUBS 0.007721f
C425 B.n372 VSUBS 0.007721f
C426 B.n373 VSUBS 0.007721f
C427 B.n374 VSUBS 0.007721f
C428 B.n375 VSUBS 0.007721f
C429 B.n376 VSUBS 0.007721f
C430 B.n377 VSUBS 0.007721f
C431 B.n378 VSUBS 0.007721f
C432 B.n379 VSUBS 0.018599f
C433 B.n380 VSUBS 0.017686f
C434 B.n381 VSUBS 0.018421f
C435 B.n382 VSUBS 0.007721f
C436 B.n383 VSUBS 0.007721f
C437 B.n384 VSUBS 0.007721f
C438 B.n385 VSUBS 0.007721f
C439 B.n386 VSUBS 0.007721f
C440 B.n387 VSUBS 0.007721f
C441 B.n388 VSUBS 0.007721f
C442 B.n389 VSUBS 0.007721f
C443 B.n390 VSUBS 0.007721f
C444 B.n391 VSUBS 0.007721f
C445 B.n392 VSUBS 0.007721f
C446 B.n393 VSUBS 0.007721f
C447 B.n394 VSUBS 0.007721f
C448 B.n395 VSUBS 0.007721f
C449 B.n396 VSUBS 0.007721f
C450 B.n397 VSUBS 0.007721f
C451 B.n398 VSUBS 0.007721f
C452 B.n399 VSUBS 0.007721f
C453 B.n400 VSUBS 0.007721f
C454 B.n401 VSUBS 0.007721f
C455 B.n402 VSUBS 0.007721f
C456 B.n403 VSUBS 0.007721f
C457 B.n404 VSUBS 0.007721f
C458 B.n405 VSUBS 0.007721f
C459 B.n406 VSUBS 0.007721f
C460 B.n407 VSUBS 0.007721f
C461 B.n408 VSUBS 0.007721f
C462 B.n409 VSUBS 0.007721f
C463 B.n410 VSUBS 0.007721f
C464 B.n411 VSUBS 0.007721f
C465 B.n412 VSUBS 0.007721f
C466 B.n413 VSUBS 0.007721f
C467 B.n414 VSUBS 0.007721f
C468 B.n415 VSUBS 0.007721f
C469 B.n416 VSUBS 0.007721f
C470 B.n417 VSUBS 0.007721f
C471 B.n418 VSUBS 0.007721f
C472 B.n419 VSUBS 0.007721f
C473 B.n420 VSUBS 0.007721f
C474 B.n421 VSUBS 0.007721f
C475 B.n422 VSUBS 0.007721f
C476 B.n423 VSUBS 0.007721f
C477 B.n424 VSUBS 0.007721f
C478 B.n425 VSUBS 0.007721f
C479 B.n426 VSUBS 0.007721f
C480 B.n427 VSUBS 0.007721f
C481 B.n428 VSUBS 0.007721f
C482 B.n429 VSUBS 0.007721f
C483 B.n430 VSUBS 0.007721f
C484 B.n431 VSUBS 0.007721f
C485 B.n432 VSUBS 0.007721f
C486 B.n433 VSUBS 0.007721f
C487 B.n434 VSUBS 0.007721f
C488 B.n435 VSUBS 0.007721f
C489 B.n436 VSUBS 0.007721f
C490 B.n437 VSUBS 0.007721f
C491 B.n438 VSUBS 0.007721f
C492 B.n439 VSUBS 0.007267f
C493 B.n440 VSUBS 0.007721f
C494 B.n441 VSUBS 0.007721f
C495 B.n442 VSUBS 0.004315f
C496 B.n443 VSUBS 0.007721f
C497 B.n444 VSUBS 0.007721f
C498 B.n445 VSUBS 0.007721f
C499 B.n446 VSUBS 0.007721f
C500 B.n447 VSUBS 0.007721f
C501 B.n448 VSUBS 0.007721f
C502 B.n449 VSUBS 0.007721f
C503 B.n450 VSUBS 0.007721f
C504 B.n451 VSUBS 0.007721f
C505 B.n452 VSUBS 0.007721f
C506 B.n453 VSUBS 0.007721f
C507 B.n454 VSUBS 0.007721f
C508 B.n455 VSUBS 0.004315f
C509 B.n456 VSUBS 0.017889f
C510 B.n457 VSUBS 0.007267f
C511 B.n458 VSUBS 0.007721f
C512 B.n459 VSUBS 0.007721f
C513 B.n460 VSUBS 0.007721f
C514 B.n461 VSUBS 0.007721f
C515 B.n462 VSUBS 0.007721f
C516 B.n463 VSUBS 0.007721f
C517 B.n464 VSUBS 0.007721f
C518 B.n465 VSUBS 0.007721f
C519 B.n466 VSUBS 0.007721f
C520 B.n467 VSUBS 0.007721f
C521 B.n468 VSUBS 0.007721f
C522 B.n469 VSUBS 0.007721f
C523 B.n470 VSUBS 0.007721f
C524 B.n471 VSUBS 0.007721f
C525 B.n472 VSUBS 0.007721f
C526 B.n473 VSUBS 0.007721f
C527 B.n474 VSUBS 0.007721f
C528 B.n475 VSUBS 0.007721f
C529 B.n476 VSUBS 0.007721f
C530 B.n477 VSUBS 0.007721f
C531 B.n478 VSUBS 0.007721f
C532 B.n479 VSUBS 0.007721f
C533 B.n480 VSUBS 0.007721f
C534 B.n481 VSUBS 0.007721f
C535 B.n482 VSUBS 0.007721f
C536 B.n483 VSUBS 0.007721f
C537 B.n484 VSUBS 0.007721f
C538 B.n485 VSUBS 0.007721f
C539 B.n486 VSUBS 0.007721f
C540 B.n487 VSUBS 0.007721f
C541 B.n488 VSUBS 0.007721f
C542 B.n489 VSUBS 0.007721f
C543 B.n490 VSUBS 0.007721f
C544 B.n491 VSUBS 0.007721f
C545 B.n492 VSUBS 0.007721f
C546 B.n493 VSUBS 0.007721f
C547 B.n494 VSUBS 0.007721f
C548 B.n495 VSUBS 0.007721f
C549 B.n496 VSUBS 0.007721f
C550 B.n497 VSUBS 0.007721f
C551 B.n498 VSUBS 0.007721f
C552 B.n499 VSUBS 0.007721f
C553 B.n500 VSUBS 0.007721f
C554 B.n501 VSUBS 0.007721f
C555 B.n502 VSUBS 0.007721f
C556 B.n503 VSUBS 0.007721f
C557 B.n504 VSUBS 0.007721f
C558 B.n505 VSUBS 0.007721f
C559 B.n506 VSUBS 0.007721f
C560 B.n507 VSUBS 0.007721f
C561 B.n508 VSUBS 0.007721f
C562 B.n509 VSUBS 0.007721f
C563 B.n510 VSUBS 0.007721f
C564 B.n511 VSUBS 0.007721f
C565 B.n512 VSUBS 0.007721f
C566 B.n513 VSUBS 0.007721f
C567 B.n514 VSUBS 0.007721f
C568 B.n515 VSUBS 0.007721f
C569 B.n516 VSUBS 0.018421f
C570 B.n517 VSUBS 0.017686f
C571 B.n518 VSUBS 0.017686f
C572 B.n519 VSUBS 0.007721f
C573 B.n520 VSUBS 0.007721f
C574 B.n521 VSUBS 0.007721f
C575 B.n522 VSUBS 0.007721f
C576 B.n523 VSUBS 0.007721f
C577 B.n524 VSUBS 0.007721f
C578 B.n525 VSUBS 0.007721f
C579 B.n526 VSUBS 0.007721f
C580 B.n527 VSUBS 0.007721f
C581 B.n528 VSUBS 0.007721f
C582 B.n529 VSUBS 0.007721f
C583 B.n530 VSUBS 0.007721f
C584 B.n531 VSUBS 0.007721f
C585 B.n532 VSUBS 0.007721f
C586 B.n533 VSUBS 0.007721f
C587 B.n534 VSUBS 0.007721f
C588 B.n535 VSUBS 0.007721f
C589 B.n536 VSUBS 0.007721f
C590 B.n537 VSUBS 0.007721f
C591 B.n538 VSUBS 0.007721f
C592 B.n539 VSUBS 0.007721f
C593 B.n540 VSUBS 0.007721f
C594 B.n541 VSUBS 0.007721f
C595 B.n542 VSUBS 0.007721f
C596 B.n543 VSUBS 0.007721f
C597 B.n544 VSUBS 0.007721f
C598 B.n545 VSUBS 0.007721f
C599 B.n546 VSUBS 0.007721f
C600 B.n547 VSUBS 0.007721f
C601 B.n548 VSUBS 0.007721f
C602 B.n549 VSUBS 0.007721f
C603 B.n550 VSUBS 0.007721f
C604 B.n551 VSUBS 0.017483f
C605 VTAIL.n0 VSUBS 0.026049f
C606 VTAIL.n1 VSUBS 0.022911f
C607 VTAIL.n2 VSUBS 0.012311f
C608 VTAIL.n3 VSUBS 0.029099f
C609 VTAIL.n4 VSUBS 0.013035f
C610 VTAIL.n5 VSUBS 0.022911f
C611 VTAIL.n6 VSUBS 0.012311f
C612 VTAIL.n7 VSUBS 0.029099f
C613 VTAIL.n8 VSUBS 0.012673f
C614 VTAIL.n9 VSUBS 0.022911f
C615 VTAIL.n10 VSUBS 0.013035f
C616 VTAIL.n11 VSUBS 0.029099f
C617 VTAIL.n12 VSUBS 0.013035f
C618 VTAIL.n13 VSUBS 0.022911f
C619 VTAIL.n14 VSUBS 0.012311f
C620 VTAIL.n15 VSUBS 0.029099f
C621 VTAIL.n16 VSUBS 0.013035f
C622 VTAIL.n17 VSUBS 1.07949f
C623 VTAIL.n18 VSUBS 0.012311f
C624 VTAIL.t2 VSUBS 0.062676f
C625 VTAIL.n19 VSUBS 0.175676f
C626 VTAIL.n20 VSUBS 0.02189f
C627 VTAIL.n21 VSUBS 0.021825f
C628 VTAIL.n22 VSUBS 0.029099f
C629 VTAIL.n23 VSUBS 0.013035f
C630 VTAIL.n24 VSUBS 0.012311f
C631 VTAIL.n25 VSUBS 0.022911f
C632 VTAIL.n26 VSUBS 0.022911f
C633 VTAIL.n27 VSUBS 0.012311f
C634 VTAIL.n28 VSUBS 0.013035f
C635 VTAIL.n29 VSUBS 0.029099f
C636 VTAIL.n30 VSUBS 0.029099f
C637 VTAIL.n31 VSUBS 0.013035f
C638 VTAIL.n32 VSUBS 0.012311f
C639 VTAIL.n33 VSUBS 0.022911f
C640 VTAIL.n34 VSUBS 0.022911f
C641 VTAIL.n35 VSUBS 0.012311f
C642 VTAIL.n36 VSUBS 0.012311f
C643 VTAIL.n37 VSUBS 0.013035f
C644 VTAIL.n38 VSUBS 0.029099f
C645 VTAIL.n39 VSUBS 0.029099f
C646 VTAIL.n40 VSUBS 0.029099f
C647 VTAIL.n41 VSUBS 0.012673f
C648 VTAIL.n42 VSUBS 0.012311f
C649 VTAIL.n43 VSUBS 0.022911f
C650 VTAIL.n44 VSUBS 0.022911f
C651 VTAIL.n45 VSUBS 0.012311f
C652 VTAIL.n46 VSUBS 0.013035f
C653 VTAIL.n47 VSUBS 0.029099f
C654 VTAIL.n48 VSUBS 0.029099f
C655 VTAIL.n49 VSUBS 0.013035f
C656 VTAIL.n50 VSUBS 0.012311f
C657 VTAIL.n51 VSUBS 0.022911f
C658 VTAIL.n52 VSUBS 0.022911f
C659 VTAIL.n53 VSUBS 0.012311f
C660 VTAIL.n54 VSUBS 0.013035f
C661 VTAIL.n55 VSUBS 0.029099f
C662 VTAIL.n56 VSUBS 0.073428f
C663 VTAIL.n57 VSUBS 0.013035f
C664 VTAIL.n58 VSUBS 0.012311f
C665 VTAIL.n59 VSUBS 0.057339f
C666 VTAIL.n60 VSUBS 0.037189f
C667 VTAIL.n61 VSUBS 0.110984f
C668 VTAIL.n62 VSUBS 0.026049f
C669 VTAIL.n63 VSUBS 0.022911f
C670 VTAIL.n64 VSUBS 0.012311f
C671 VTAIL.n65 VSUBS 0.029099f
C672 VTAIL.n66 VSUBS 0.013035f
C673 VTAIL.n67 VSUBS 0.022911f
C674 VTAIL.n68 VSUBS 0.012311f
C675 VTAIL.n69 VSUBS 0.029099f
C676 VTAIL.n70 VSUBS 0.012673f
C677 VTAIL.n71 VSUBS 0.022911f
C678 VTAIL.n72 VSUBS 0.013035f
C679 VTAIL.n73 VSUBS 0.029099f
C680 VTAIL.n74 VSUBS 0.013035f
C681 VTAIL.n75 VSUBS 0.022911f
C682 VTAIL.n76 VSUBS 0.012311f
C683 VTAIL.n77 VSUBS 0.029099f
C684 VTAIL.n78 VSUBS 0.013035f
C685 VTAIL.n79 VSUBS 1.07949f
C686 VTAIL.n80 VSUBS 0.012311f
C687 VTAIL.t5 VSUBS 0.062676f
C688 VTAIL.n81 VSUBS 0.175676f
C689 VTAIL.n82 VSUBS 0.02189f
C690 VTAIL.n83 VSUBS 0.021825f
C691 VTAIL.n84 VSUBS 0.029099f
C692 VTAIL.n85 VSUBS 0.013035f
C693 VTAIL.n86 VSUBS 0.012311f
C694 VTAIL.n87 VSUBS 0.022911f
C695 VTAIL.n88 VSUBS 0.022911f
C696 VTAIL.n89 VSUBS 0.012311f
C697 VTAIL.n90 VSUBS 0.013035f
C698 VTAIL.n91 VSUBS 0.029099f
C699 VTAIL.n92 VSUBS 0.029099f
C700 VTAIL.n93 VSUBS 0.013035f
C701 VTAIL.n94 VSUBS 0.012311f
C702 VTAIL.n95 VSUBS 0.022911f
C703 VTAIL.n96 VSUBS 0.022911f
C704 VTAIL.n97 VSUBS 0.012311f
C705 VTAIL.n98 VSUBS 0.012311f
C706 VTAIL.n99 VSUBS 0.013035f
C707 VTAIL.n100 VSUBS 0.029099f
C708 VTAIL.n101 VSUBS 0.029099f
C709 VTAIL.n102 VSUBS 0.029099f
C710 VTAIL.n103 VSUBS 0.012673f
C711 VTAIL.n104 VSUBS 0.012311f
C712 VTAIL.n105 VSUBS 0.022911f
C713 VTAIL.n106 VSUBS 0.022911f
C714 VTAIL.n107 VSUBS 0.012311f
C715 VTAIL.n108 VSUBS 0.013035f
C716 VTAIL.n109 VSUBS 0.029099f
C717 VTAIL.n110 VSUBS 0.029099f
C718 VTAIL.n111 VSUBS 0.013035f
C719 VTAIL.n112 VSUBS 0.012311f
C720 VTAIL.n113 VSUBS 0.022911f
C721 VTAIL.n114 VSUBS 0.022911f
C722 VTAIL.n115 VSUBS 0.012311f
C723 VTAIL.n116 VSUBS 0.013035f
C724 VTAIL.n117 VSUBS 0.029099f
C725 VTAIL.n118 VSUBS 0.073428f
C726 VTAIL.n119 VSUBS 0.013035f
C727 VTAIL.n120 VSUBS 0.012311f
C728 VTAIL.n121 VSUBS 0.057339f
C729 VTAIL.n122 VSUBS 0.037189f
C730 VTAIL.n123 VSUBS 0.156647f
C731 VTAIL.n124 VSUBS 0.026049f
C732 VTAIL.n125 VSUBS 0.022911f
C733 VTAIL.n126 VSUBS 0.012311f
C734 VTAIL.n127 VSUBS 0.029099f
C735 VTAIL.n128 VSUBS 0.013035f
C736 VTAIL.n129 VSUBS 0.022911f
C737 VTAIL.n130 VSUBS 0.012311f
C738 VTAIL.n131 VSUBS 0.029099f
C739 VTAIL.n132 VSUBS 0.012673f
C740 VTAIL.n133 VSUBS 0.022911f
C741 VTAIL.n134 VSUBS 0.013035f
C742 VTAIL.n135 VSUBS 0.029099f
C743 VTAIL.n136 VSUBS 0.013035f
C744 VTAIL.n137 VSUBS 0.022911f
C745 VTAIL.n138 VSUBS 0.012311f
C746 VTAIL.n139 VSUBS 0.029099f
C747 VTAIL.n140 VSUBS 0.013035f
C748 VTAIL.n141 VSUBS 1.07949f
C749 VTAIL.n142 VSUBS 0.012311f
C750 VTAIL.t7 VSUBS 0.062676f
C751 VTAIL.n143 VSUBS 0.175676f
C752 VTAIL.n144 VSUBS 0.02189f
C753 VTAIL.n145 VSUBS 0.021825f
C754 VTAIL.n146 VSUBS 0.029099f
C755 VTAIL.n147 VSUBS 0.013035f
C756 VTAIL.n148 VSUBS 0.012311f
C757 VTAIL.n149 VSUBS 0.022911f
C758 VTAIL.n150 VSUBS 0.022911f
C759 VTAIL.n151 VSUBS 0.012311f
C760 VTAIL.n152 VSUBS 0.013035f
C761 VTAIL.n153 VSUBS 0.029099f
C762 VTAIL.n154 VSUBS 0.029099f
C763 VTAIL.n155 VSUBS 0.013035f
C764 VTAIL.n156 VSUBS 0.012311f
C765 VTAIL.n157 VSUBS 0.022911f
C766 VTAIL.n158 VSUBS 0.022911f
C767 VTAIL.n159 VSUBS 0.012311f
C768 VTAIL.n160 VSUBS 0.012311f
C769 VTAIL.n161 VSUBS 0.013035f
C770 VTAIL.n162 VSUBS 0.029099f
C771 VTAIL.n163 VSUBS 0.029099f
C772 VTAIL.n164 VSUBS 0.029099f
C773 VTAIL.n165 VSUBS 0.012673f
C774 VTAIL.n166 VSUBS 0.012311f
C775 VTAIL.n167 VSUBS 0.022911f
C776 VTAIL.n168 VSUBS 0.022911f
C777 VTAIL.n169 VSUBS 0.012311f
C778 VTAIL.n170 VSUBS 0.013035f
C779 VTAIL.n171 VSUBS 0.029099f
C780 VTAIL.n172 VSUBS 0.029099f
C781 VTAIL.n173 VSUBS 0.013035f
C782 VTAIL.n174 VSUBS 0.012311f
C783 VTAIL.n175 VSUBS 0.022911f
C784 VTAIL.n176 VSUBS 0.022911f
C785 VTAIL.n177 VSUBS 0.012311f
C786 VTAIL.n178 VSUBS 0.013035f
C787 VTAIL.n179 VSUBS 0.029099f
C788 VTAIL.n180 VSUBS 0.073428f
C789 VTAIL.n181 VSUBS 0.013035f
C790 VTAIL.n182 VSUBS 0.012311f
C791 VTAIL.n183 VSUBS 0.057339f
C792 VTAIL.n184 VSUBS 0.037189f
C793 VTAIL.n185 VSUBS 1.26752f
C794 VTAIL.n186 VSUBS 0.026049f
C795 VTAIL.n187 VSUBS 0.022911f
C796 VTAIL.n188 VSUBS 0.012311f
C797 VTAIL.n189 VSUBS 0.029099f
C798 VTAIL.n190 VSUBS 0.013035f
C799 VTAIL.n191 VSUBS 0.022911f
C800 VTAIL.n192 VSUBS 0.012311f
C801 VTAIL.n193 VSUBS 0.029099f
C802 VTAIL.n194 VSUBS 0.012673f
C803 VTAIL.n195 VSUBS 0.022911f
C804 VTAIL.n196 VSUBS 0.012673f
C805 VTAIL.n197 VSUBS 0.012311f
C806 VTAIL.n198 VSUBS 0.029099f
C807 VTAIL.n199 VSUBS 0.029099f
C808 VTAIL.n200 VSUBS 0.013035f
C809 VTAIL.n201 VSUBS 0.022911f
C810 VTAIL.n202 VSUBS 0.012311f
C811 VTAIL.n203 VSUBS 0.029099f
C812 VTAIL.n204 VSUBS 0.013035f
C813 VTAIL.n205 VSUBS 1.07949f
C814 VTAIL.n206 VSUBS 0.012311f
C815 VTAIL.t0 VSUBS 0.062676f
C816 VTAIL.n207 VSUBS 0.175676f
C817 VTAIL.n208 VSUBS 0.02189f
C818 VTAIL.n209 VSUBS 0.021825f
C819 VTAIL.n210 VSUBS 0.029099f
C820 VTAIL.n211 VSUBS 0.013035f
C821 VTAIL.n212 VSUBS 0.012311f
C822 VTAIL.n213 VSUBS 0.022911f
C823 VTAIL.n214 VSUBS 0.022911f
C824 VTAIL.n215 VSUBS 0.012311f
C825 VTAIL.n216 VSUBS 0.013035f
C826 VTAIL.n217 VSUBS 0.029099f
C827 VTAIL.n218 VSUBS 0.029099f
C828 VTAIL.n219 VSUBS 0.013035f
C829 VTAIL.n220 VSUBS 0.012311f
C830 VTAIL.n221 VSUBS 0.022911f
C831 VTAIL.n222 VSUBS 0.022911f
C832 VTAIL.n223 VSUBS 0.012311f
C833 VTAIL.n224 VSUBS 0.013035f
C834 VTAIL.n225 VSUBS 0.029099f
C835 VTAIL.n226 VSUBS 0.029099f
C836 VTAIL.n227 VSUBS 0.013035f
C837 VTAIL.n228 VSUBS 0.012311f
C838 VTAIL.n229 VSUBS 0.022911f
C839 VTAIL.n230 VSUBS 0.022911f
C840 VTAIL.n231 VSUBS 0.012311f
C841 VTAIL.n232 VSUBS 0.013035f
C842 VTAIL.n233 VSUBS 0.029099f
C843 VTAIL.n234 VSUBS 0.029099f
C844 VTAIL.n235 VSUBS 0.013035f
C845 VTAIL.n236 VSUBS 0.012311f
C846 VTAIL.n237 VSUBS 0.022911f
C847 VTAIL.n238 VSUBS 0.022911f
C848 VTAIL.n239 VSUBS 0.012311f
C849 VTAIL.n240 VSUBS 0.013035f
C850 VTAIL.n241 VSUBS 0.029099f
C851 VTAIL.n242 VSUBS 0.073428f
C852 VTAIL.n243 VSUBS 0.013035f
C853 VTAIL.n244 VSUBS 0.012311f
C854 VTAIL.n245 VSUBS 0.057339f
C855 VTAIL.n246 VSUBS 0.037189f
C856 VTAIL.n247 VSUBS 1.26752f
C857 VTAIL.n248 VSUBS 0.026049f
C858 VTAIL.n249 VSUBS 0.022911f
C859 VTAIL.n250 VSUBS 0.012311f
C860 VTAIL.n251 VSUBS 0.029099f
C861 VTAIL.n252 VSUBS 0.013035f
C862 VTAIL.n253 VSUBS 0.022911f
C863 VTAIL.n254 VSUBS 0.012311f
C864 VTAIL.n255 VSUBS 0.029099f
C865 VTAIL.n256 VSUBS 0.012673f
C866 VTAIL.n257 VSUBS 0.022911f
C867 VTAIL.n258 VSUBS 0.012673f
C868 VTAIL.n259 VSUBS 0.012311f
C869 VTAIL.n260 VSUBS 0.029099f
C870 VTAIL.n261 VSUBS 0.029099f
C871 VTAIL.n262 VSUBS 0.013035f
C872 VTAIL.n263 VSUBS 0.022911f
C873 VTAIL.n264 VSUBS 0.012311f
C874 VTAIL.n265 VSUBS 0.029099f
C875 VTAIL.n266 VSUBS 0.013035f
C876 VTAIL.n267 VSUBS 1.07949f
C877 VTAIL.n268 VSUBS 0.012311f
C878 VTAIL.t3 VSUBS 0.062676f
C879 VTAIL.n269 VSUBS 0.175676f
C880 VTAIL.n270 VSUBS 0.02189f
C881 VTAIL.n271 VSUBS 0.021825f
C882 VTAIL.n272 VSUBS 0.029099f
C883 VTAIL.n273 VSUBS 0.013035f
C884 VTAIL.n274 VSUBS 0.012311f
C885 VTAIL.n275 VSUBS 0.022911f
C886 VTAIL.n276 VSUBS 0.022911f
C887 VTAIL.n277 VSUBS 0.012311f
C888 VTAIL.n278 VSUBS 0.013035f
C889 VTAIL.n279 VSUBS 0.029099f
C890 VTAIL.n280 VSUBS 0.029099f
C891 VTAIL.n281 VSUBS 0.013035f
C892 VTAIL.n282 VSUBS 0.012311f
C893 VTAIL.n283 VSUBS 0.022911f
C894 VTAIL.n284 VSUBS 0.022911f
C895 VTAIL.n285 VSUBS 0.012311f
C896 VTAIL.n286 VSUBS 0.013035f
C897 VTAIL.n287 VSUBS 0.029099f
C898 VTAIL.n288 VSUBS 0.029099f
C899 VTAIL.n289 VSUBS 0.013035f
C900 VTAIL.n290 VSUBS 0.012311f
C901 VTAIL.n291 VSUBS 0.022911f
C902 VTAIL.n292 VSUBS 0.022911f
C903 VTAIL.n293 VSUBS 0.012311f
C904 VTAIL.n294 VSUBS 0.013035f
C905 VTAIL.n295 VSUBS 0.029099f
C906 VTAIL.n296 VSUBS 0.029099f
C907 VTAIL.n297 VSUBS 0.013035f
C908 VTAIL.n298 VSUBS 0.012311f
C909 VTAIL.n299 VSUBS 0.022911f
C910 VTAIL.n300 VSUBS 0.022911f
C911 VTAIL.n301 VSUBS 0.012311f
C912 VTAIL.n302 VSUBS 0.013035f
C913 VTAIL.n303 VSUBS 0.029099f
C914 VTAIL.n304 VSUBS 0.073428f
C915 VTAIL.n305 VSUBS 0.013035f
C916 VTAIL.n306 VSUBS 0.012311f
C917 VTAIL.n307 VSUBS 0.057339f
C918 VTAIL.n308 VSUBS 0.037189f
C919 VTAIL.n309 VSUBS 0.156647f
C920 VTAIL.n310 VSUBS 0.026049f
C921 VTAIL.n311 VSUBS 0.022911f
C922 VTAIL.n312 VSUBS 0.012311f
C923 VTAIL.n313 VSUBS 0.029099f
C924 VTAIL.n314 VSUBS 0.013035f
C925 VTAIL.n315 VSUBS 0.022911f
C926 VTAIL.n316 VSUBS 0.012311f
C927 VTAIL.n317 VSUBS 0.029099f
C928 VTAIL.n318 VSUBS 0.012673f
C929 VTAIL.n319 VSUBS 0.022911f
C930 VTAIL.n320 VSUBS 0.012673f
C931 VTAIL.n321 VSUBS 0.012311f
C932 VTAIL.n322 VSUBS 0.029099f
C933 VTAIL.n323 VSUBS 0.029099f
C934 VTAIL.n324 VSUBS 0.013035f
C935 VTAIL.n325 VSUBS 0.022911f
C936 VTAIL.n326 VSUBS 0.012311f
C937 VTAIL.n327 VSUBS 0.029099f
C938 VTAIL.n328 VSUBS 0.013035f
C939 VTAIL.n329 VSUBS 1.07949f
C940 VTAIL.n330 VSUBS 0.012311f
C941 VTAIL.t6 VSUBS 0.062676f
C942 VTAIL.n331 VSUBS 0.175676f
C943 VTAIL.n332 VSUBS 0.02189f
C944 VTAIL.n333 VSUBS 0.021825f
C945 VTAIL.n334 VSUBS 0.029099f
C946 VTAIL.n335 VSUBS 0.013035f
C947 VTAIL.n336 VSUBS 0.012311f
C948 VTAIL.n337 VSUBS 0.022911f
C949 VTAIL.n338 VSUBS 0.022911f
C950 VTAIL.n339 VSUBS 0.012311f
C951 VTAIL.n340 VSUBS 0.013035f
C952 VTAIL.n341 VSUBS 0.029099f
C953 VTAIL.n342 VSUBS 0.029099f
C954 VTAIL.n343 VSUBS 0.013035f
C955 VTAIL.n344 VSUBS 0.012311f
C956 VTAIL.n345 VSUBS 0.022911f
C957 VTAIL.n346 VSUBS 0.022911f
C958 VTAIL.n347 VSUBS 0.012311f
C959 VTAIL.n348 VSUBS 0.013035f
C960 VTAIL.n349 VSUBS 0.029099f
C961 VTAIL.n350 VSUBS 0.029099f
C962 VTAIL.n351 VSUBS 0.013035f
C963 VTAIL.n352 VSUBS 0.012311f
C964 VTAIL.n353 VSUBS 0.022911f
C965 VTAIL.n354 VSUBS 0.022911f
C966 VTAIL.n355 VSUBS 0.012311f
C967 VTAIL.n356 VSUBS 0.013035f
C968 VTAIL.n357 VSUBS 0.029099f
C969 VTAIL.n358 VSUBS 0.029099f
C970 VTAIL.n359 VSUBS 0.013035f
C971 VTAIL.n360 VSUBS 0.012311f
C972 VTAIL.n361 VSUBS 0.022911f
C973 VTAIL.n362 VSUBS 0.022911f
C974 VTAIL.n363 VSUBS 0.012311f
C975 VTAIL.n364 VSUBS 0.013035f
C976 VTAIL.n365 VSUBS 0.029099f
C977 VTAIL.n366 VSUBS 0.073428f
C978 VTAIL.n367 VSUBS 0.013035f
C979 VTAIL.n368 VSUBS 0.012311f
C980 VTAIL.n369 VSUBS 0.057339f
C981 VTAIL.n370 VSUBS 0.037189f
C982 VTAIL.n371 VSUBS 0.156647f
C983 VTAIL.n372 VSUBS 0.026049f
C984 VTAIL.n373 VSUBS 0.022911f
C985 VTAIL.n374 VSUBS 0.012311f
C986 VTAIL.n375 VSUBS 0.029099f
C987 VTAIL.n376 VSUBS 0.013035f
C988 VTAIL.n377 VSUBS 0.022911f
C989 VTAIL.n378 VSUBS 0.012311f
C990 VTAIL.n379 VSUBS 0.029099f
C991 VTAIL.n380 VSUBS 0.012673f
C992 VTAIL.n381 VSUBS 0.022911f
C993 VTAIL.n382 VSUBS 0.012673f
C994 VTAIL.n383 VSUBS 0.012311f
C995 VTAIL.n384 VSUBS 0.029099f
C996 VTAIL.n385 VSUBS 0.029099f
C997 VTAIL.n386 VSUBS 0.013035f
C998 VTAIL.n387 VSUBS 0.022911f
C999 VTAIL.n388 VSUBS 0.012311f
C1000 VTAIL.n389 VSUBS 0.029099f
C1001 VTAIL.n390 VSUBS 0.013035f
C1002 VTAIL.n391 VSUBS 1.07949f
C1003 VTAIL.n392 VSUBS 0.012311f
C1004 VTAIL.t4 VSUBS 0.062676f
C1005 VTAIL.n393 VSUBS 0.175676f
C1006 VTAIL.n394 VSUBS 0.02189f
C1007 VTAIL.n395 VSUBS 0.021825f
C1008 VTAIL.n396 VSUBS 0.029099f
C1009 VTAIL.n397 VSUBS 0.013035f
C1010 VTAIL.n398 VSUBS 0.012311f
C1011 VTAIL.n399 VSUBS 0.022911f
C1012 VTAIL.n400 VSUBS 0.022911f
C1013 VTAIL.n401 VSUBS 0.012311f
C1014 VTAIL.n402 VSUBS 0.013035f
C1015 VTAIL.n403 VSUBS 0.029099f
C1016 VTAIL.n404 VSUBS 0.029099f
C1017 VTAIL.n405 VSUBS 0.013035f
C1018 VTAIL.n406 VSUBS 0.012311f
C1019 VTAIL.n407 VSUBS 0.022911f
C1020 VTAIL.n408 VSUBS 0.022911f
C1021 VTAIL.n409 VSUBS 0.012311f
C1022 VTAIL.n410 VSUBS 0.013035f
C1023 VTAIL.n411 VSUBS 0.029099f
C1024 VTAIL.n412 VSUBS 0.029099f
C1025 VTAIL.n413 VSUBS 0.013035f
C1026 VTAIL.n414 VSUBS 0.012311f
C1027 VTAIL.n415 VSUBS 0.022911f
C1028 VTAIL.n416 VSUBS 0.022911f
C1029 VTAIL.n417 VSUBS 0.012311f
C1030 VTAIL.n418 VSUBS 0.013035f
C1031 VTAIL.n419 VSUBS 0.029099f
C1032 VTAIL.n420 VSUBS 0.029099f
C1033 VTAIL.n421 VSUBS 0.013035f
C1034 VTAIL.n422 VSUBS 0.012311f
C1035 VTAIL.n423 VSUBS 0.022911f
C1036 VTAIL.n424 VSUBS 0.022911f
C1037 VTAIL.n425 VSUBS 0.012311f
C1038 VTAIL.n426 VSUBS 0.013035f
C1039 VTAIL.n427 VSUBS 0.029099f
C1040 VTAIL.n428 VSUBS 0.073428f
C1041 VTAIL.n429 VSUBS 0.013035f
C1042 VTAIL.n430 VSUBS 0.012311f
C1043 VTAIL.n431 VSUBS 0.057339f
C1044 VTAIL.n432 VSUBS 0.037189f
C1045 VTAIL.n433 VSUBS 1.26752f
C1046 VTAIL.n434 VSUBS 0.026049f
C1047 VTAIL.n435 VSUBS 0.022911f
C1048 VTAIL.n436 VSUBS 0.012311f
C1049 VTAIL.n437 VSUBS 0.029099f
C1050 VTAIL.n438 VSUBS 0.013035f
C1051 VTAIL.n439 VSUBS 0.022911f
C1052 VTAIL.n440 VSUBS 0.012311f
C1053 VTAIL.n441 VSUBS 0.029099f
C1054 VTAIL.n442 VSUBS 0.012673f
C1055 VTAIL.n443 VSUBS 0.022911f
C1056 VTAIL.n444 VSUBS 0.013035f
C1057 VTAIL.n445 VSUBS 0.029099f
C1058 VTAIL.n446 VSUBS 0.013035f
C1059 VTAIL.n447 VSUBS 0.022911f
C1060 VTAIL.n448 VSUBS 0.012311f
C1061 VTAIL.n449 VSUBS 0.029099f
C1062 VTAIL.n450 VSUBS 0.013035f
C1063 VTAIL.n451 VSUBS 1.07949f
C1064 VTAIL.n452 VSUBS 0.012311f
C1065 VTAIL.t1 VSUBS 0.062676f
C1066 VTAIL.n453 VSUBS 0.175676f
C1067 VTAIL.n454 VSUBS 0.02189f
C1068 VTAIL.n455 VSUBS 0.021825f
C1069 VTAIL.n456 VSUBS 0.029099f
C1070 VTAIL.n457 VSUBS 0.013035f
C1071 VTAIL.n458 VSUBS 0.012311f
C1072 VTAIL.n459 VSUBS 0.022911f
C1073 VTAIL.n460 VSUBS 0.022911f
C1074 VTAIL.n461 VSUBS 0.012311f
C1075 VTAIL.n462 VSUBS 0.013035f
C1076 VTAIL.n463 VSUBS 0.029099f
C1077 VTAIL.n464 VSUBS 0.029099f
C1078 VTAIL.n465 VSUBS 0.013035f
C1079 VTAIL.n466 VSUBS 0.012311f
C1080 VTAIL.n467 VSUBS 0.022911f
C1081 VTAIL.n468 VSUBS 0.022911f
C1082 VTAIL.n469 VSUBS 0.012311f
C1083 VTAIL.n470 VSUBS 0.012311f
C1084 VTAIL.n471 VSUBS 0.013035f
C1085 VTAIL.n472 VSUBS 0.029099f
C1086 VTAIL.n473 VSUBS 0.029099f
C1087 VTAIL.n474 VSUBS 0.029099f
C1088 VTAIL.n475 VSUBS 0.012673f
C1089 VTAIL.n476 VSUBS 0.012311f
C1090 VTAIL.n477 VSUBS 0.022911f
C1091 VTAIL.n478 VSUBS 0.022911f
C1092 VTAIL.n479 VSUBS 0.012311f
C1093 VTAIL.n480 VSUBS 0.013035f
C1094 VTAIL.n481 VSUBS 0.029099f
C1095 VTAIL.n482 VSUBS 0.029099f
C1096 VTAIL.n483 VSUBS 0.013035f
C1097 VTAIL.n484 VSUBS 0.012311f
C1098 VTAIL.n485 VSUBS 0.022911f
C1099 VTAIL.n486 VSUBS 0.022911f
C1100 VTAIL.n487 VSUBS 0.012311f
C1101 VTAIL.n488 VSUBS 0.013035f
C1102 VTAIL.n489 VSUBS 0.029099f
C1103 VTAIL.n490 VSUBS 0.073428f
C1104 VTAIL.n491 VSUBS 0.013035f
C1105 VTAIL.n492 VSUBS 0.012311f
C1106 VTAIL.n493 VSUBS 0.057339f
C1107 VTAIL.n494 VSUBS 0.037189f
C1108 VTAIL.n495 VSUBS 1.21326f
C1109 VDD1.t1 VSUBS 0.24704f
C1110 VDD1.t2 VSUBS 0.24704f
C1111 VDD1.n0 VSUBS 1.92445f
C1112 VDD1.t0 VSUBS 0.24704f
C1113 VDD1.t3 VSUBS 0.24704f
C1114 VDD1.n1 VSUBS 2.55021f
C1115 VP.n0 VSUBS 0.049474f
C1116 VP.t2 VSUBS 1.92669f
C1117 VP.n1 VSUBS 0.078335f
C1118 VP.t1 VSUBS 2.04883f
C1119 VP.t3 VSUBS 2.04806f
C1120 VP.n2 VSUBS 3.10177f
C1121 VP.t0 VSUBS 1.92669f
C1122 VP.n3 VSUBS 0.79485f
C1123 VP.n4 VSUBS 2.7485f
C1124 VP.n5 VSUBS 0.049474f
C1125 VP.n6 VSUBS 0.049474f
C1126 VP.n7 VSUBS 0.039958f
C1127 VP.n8 VSUBS 0.078335f
C1128 VP.n9 VSUBS 0.79485f
C1129 VP.n10 VSUBS 0.044124f
.ends

