* NGSPICE file created from diff_pair_sample_1553.ext - technology: sky130A

.subckt diff_pair_sample_1553 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X1 VTAIL.t15 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=1.87935 ps=11.72 w=11.39 l=2.29
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=0 ps=0 w=11.39 l=2.29
X3 VDD2.t6 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X4 VDD1.t4 VP.t1 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=4.4421 ps=23.56 w=11.39 l=2.29
X5 VTAIL.t3 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=0 ps=0 w=11.39 l=2.29
X7 VDD1.t2 VP.t2 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X8 VTAIL.t14 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X9 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X10 VDD1.t3 VP.t3 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
X11 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=1.87935 ps=11.72 w=11.39 l=2.29
X12 VDD1.t6 VP.t4 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=4.4421 ps=23.56 w=11.39 l=2.29
X13 VTAIL.t8 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=1.87935 ps=11.72 w=11.39 l=2.29
X14 VTAIL.t7 VP.t6 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=1.87935 ps=11.72 w=11.39 l=2.29
X15 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=4.4421 ps=23.56 w=11.39 l=2.29
X16 VDD2.t0 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=4.4421 ps=23.56 w=11.39 l=2.29
X17 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=0 ps=0 w=11.39 l=2.29
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4421 pd=23.56 as=0 ps=0 w=11.39 l=2.29
X19 VTAIL.t6 VP.t7 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=1.87935 pd=11.72 as=1.87935 ps=11.72 w=11.39 l=2.29
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n26 VP.n10 161.3
R7 VP.n28 VP.n27 161.3
R8 VP.n29 VP.n9 161.3
R9 VP.n31 VP.n30 161.3
R10 VP.n32 VP.n8 161.3
R11 VP.n62 VP.n0 161.3
R12 VP.n61 VP.n60 161.3
R13 VP.n59 VP.n1 161.3
R14 VP.n58 VP.n57 161.3
R15 VP.n56 VP.n2 161.3
R16 VP.n54 VP.n53 161.3
R17 VP.n52 VP.n3 161.3
R18 VP.n51 VP.n50 161.3
R19 VP.n49 VP.n4 161.3
R20 VP.n48 VP.n47 161.3
R21 VP.n46 VP.n5 161.3
R22 VP.n45 VP.n44 161.3
R23 VP.n42 VP.n6 161.3
R24 VP.n41 VP.n40 161.3
R25 VP.n39 VP.n7 161.3
R26 VP.n38 VP.n37 161.3
R27 VP.n15 VP.t5 150.291
R28 VP.n36 VP.t6 119.87
R29 VP.n43 VP.t3 119.87
R30 VP.n55 VP.t7 119.87
R31 VP.n63 VP.t1 119.87
R32 VP.n33 VP.t4 119.87
R33 VP.n25 VP.t0 119.87
R34 VP.n14 VP.t2 119.87
R35 VP.n36 VP.n35 101.948
R36 VP.n64 VP.n63 101.948
R37 VP.n34 VP.n33 101.948
R38 VP.n15 VP.n14 69.279
R39 VP.n50 VP.n49 56.5193
R40 VP.n20 VP.n19 56.5193
R41 VP.n42 VP.n41 53.1199
R42 VP.n57 VP.n1 53.1199
R43 VP.n27 VP.n9 53.1199
R44 VP.n35 VP.n34 48.9087
R45 VP.n41 VP.n7 27.8669
R46 VP.n61 VP.n1 27.8669
R47 VP.n31 VP.n9 27.8669
R48 VP.n37 VP.n7 24.4675
R49 VP.n44 VP.n42 24.4675
R50 VP.n48 VP.n5 24.4675
R51 VP.n49 VP.n48 24.4675
R52 VP.n50 VP.n3 24.4675
R53 VP.n54 VP.n3 24.4675
R54 VP.n57 VP.n56 24.4675
R55 VP.n62 VP.n61 24.4675
R56 VP.n32 VP.n31 24.4675
R57 VP.n20 VP.n11 24.4675
R58 VP.n24 VP.n11 24.4675
R59 VP.n27 VP.n26 24.4675
R60 VP.n18 VP.n13 24.4675
R61 VP.n19 VP.n18 24.4675
R62 VP.n44 VP.n43 21.5315
R63 VP.n56 VP.n55 21.5315
R64 VP.n26 VP.n25 21.5315
R65 VP.n16 VP.n15 10.1472
R66 VP.n37 VP.n36 8.80862
R67 VP.n63 VP.n62 8.80862
R68 VP.n33 VP.n32 8.80862
R69 VP.n43 VP.n5 2.93654
R70 VP.n55 VP.n54 2.93654
R71 VP.n25 VP.n24 2.93654
R72 VP.n14 VP.n13 2.93654
R73 VP.n34 VP.n8 0.278367
R74 VP.n38 VP.n35 0.278367
R75 VP.n64 VP.n0 0.278367
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153454
R102 VDD1 VDD1.n0 63.0835
R103 VDD1.n3 VDD1.n2 62.9698
R104 VDD1.n3 VDD1.n1 62.9698
R105 VDD1.n5 VDD1.n4 61.8958
R106 VDD1.n5 VDD1.n3 44.2811
R107 VDD1.n4 VDD1.t7 1.73887
R108 VDD1.n4 VDD1.t6 1.73887
R109 VDD1.n0 VDD1.t0 1.73887
R110 VDD1.n0 VDD1.t2 1.73887
R111 VDD1.n2 VDD1.t1 1.73887
R112 VDD1.n2 VDD1.t4 1.73887
R113 VDD1.n1 VDD1.t5 1.73887
R114 VDD1.n1 VDD1.t3 1.73887
R115 VDD1 VDD1.n5 1.07162
R116 VTAIL.n498 VTAIL.n442 289.615
R117 VTAIL.n58 VTAIL.n2 289.615
R118 VTAIL.n120 VTAIL.n64 289.615
R119 VTAIL.n184 VTAIL.n128 289.615
R120 VTAIL.n436 VTAIL.n380 289.615
R121 VTAIL.n372 VTAIL.n316 289.615
R122 VTAIL.n310 VTAIL.n254 289.615
R123 VTAIL.n246 VTAIL.n190 289.615
R124 VTAIL.n463 VTAIL.n462 185
R125 VTAIL.n465 VTAIL.n464 185
R126 VTAIL.n458 VTAIL.n457 185
R127 VTAIL.n471 VTAIL.n470 185
R128 VTAIL.n473 VTAIL.n472 185
R129 VTAIL.n454 VTAIL.n453 185
R130 VTAIL.n480 VTAIL.n479 185
R131 VTAIL.n481 VTAIL.n452 185
R132 VTAIL.n483 VTAIL.n482 185
R133 VTAIL.n450 VTAIL.n449 185
R134 VTAIL.n489 VTAIL.n488 185
R135 VTAIL.n491 VTAIL.n490 185
R136 VTAIL.n446 VTAIL.n445 185
R137 VTAIL.n497 VTAIL.n496 185
R138 VTAIL.n499 VTAIL.n498 185
R139 VTAIL.n23 VTAIL.n22 185
R140 VTAIL.n25 VTAIL.n24 185
R141 VTAIL.n18 VTAIL.n17 185
R142 VTAIL.n31 VTAIL.n30 185
R143 VTAIL.n33 VTAIL.n32 185
R144 VTAIL.n14 VTAIL.n13 185
R145 VTAIL.n40 VTAIL.n39 185
R146 VTAIL.n41 VTAIL.n12 185
R147 VTAIL.n43 VTAIL.n42 185
R148 VTAIL.n10 VTAIL.n9 185
R149 VTAIL.n49 VTAIL.n48 185
R150 VTAIL.n51 VTAIL.n50 185
R151 VTAIL.n6 VTAIL.n5 185
R152 VTAIL.n57 VTAIL.n56 185
R153 VTAIL.n59 VTAIL.n58 185
R154 VTAIL.n85 VTAIL.n84 185
R155 VTAIL.n87 VTAIL.n86 185
R156 VTAIL.n80 VTAIL.n79 185
R157 VTAIL.n93 VTAIL.n92 185
R158 VTAIL.n95 VTAIL.n94 185
R159 VTAIL.n76 VTAIL.n75 185
R160 VTAIL.n102 VTAIL.n101 185
R161 VTAIL.n103 VTAIL.n74 185
R162 VTAIL.n105 VTAIL.n104 185
R163 VTAIL.n72 VTAIL.n71 185
R164 VTAIL.n111 VTAIL.n110 185
R165 VTAIL.n113 VTAIL.n112 185
R166 VTAIL.n68 VTAIL.n67 185
R167 VTAIL.n119 VTAIL.n118 185
R168 VTAIL.n121 VTAIL.n120 185
R169 VTAIL.n149 VTAIL.n148 185
R170 VTAIL.n151 VTAIL.n150 185
R171 VTAIL.n144 VTAIL.n143 185
R172 VTAIL.n157 VTAIL.n156 185
R173 VTAIL.n159 VTAIL.n158 185
R174 VTAIL.n140 VTAIL.n139 185
R175 VTAIL.n166 VTAIL.n165 185
R176 VTAIL.n167 VTAIL.n138 185
R177 VTAIL.n169 VTAIL.n168 185
R178 VTAIL.n136 VTAIL.n135 185
R179 VTAIL.n175 VTAIL.n174 185
R180 VTAIL.n177 VTAIL.n176 185
R181 VTAIL.n132 VTAIL.n131 185
R182 VTAIL.n183 VTAIL.n182 185
R183 VTAIL.n185 VTAIL.n184 185
R184 VTAIL.n437 VTAIL.n436 185
R185 VTAIL.n435 VTAIL.n434 185
R186 VTAIL.n384 VTAIL.n383 185
R187 VTAIL.n429 VTAIL.n428 185
R188 VTAIL.n427 VTAIL.n426 185
R189 VTAIL.n388 VTAIL.n387 185
R190 VTAIL.n392 VTAIL.n390 185
R191 VTAIL.n421 VTAIL.n420 185
R192 VTAIL.n419 VTAIL.n418 185
R193 VTAIL.n394 VTAIL.n393 185
R194 VTAIL.n413 VTAIL.n412 185
R195 VTAIL.n411 VTAIL.n410 185
R196 VTAIL.n398 VTAIL.n397 185
R197 VTAIL.n405 VTAIL.n404 185
R198 VTAIL.n403 VTAIL.n402 185
R199 VTAIL.n373 VTAIL.n372 185
R200 VTAIL.n371 VTAIL.n370 185
R201 VTAIL.n320 VTAIL.n319 185
R202 VTAIL.n365 VTAIL.n364 185
R203 VTAIL.n363 VTAIL.n362 185
R204 VTAIL.n324 VTAIL.n323 185
R205 VTAIL.n328 VTAIL.n326 185
R206 VTAIL.n357 VTAIL.n356 185
R207 VTAIL.n355 VTAIL.n354 185
R208 VTAIL.n330 VTAIL.n329 185
R209 VTAIL.n349 VTAIL.n348 185
R210 VTAIL.n347 VTAIL.n346 185
R211 VTAIL.n334 VTAIL.n333 185
R212 VTAIL.n341 VTAIL.n340 185
R213 VTAIL.n339 VTAIL.n338 185
R214 VTAIL.n311 VTAIL.n310 185
R215 VTAIL.n309 VTAIL.n308 185
R216 VTAIL.n258 VTAIL.n257 185
R217 VTAIL.n303 VTAIL.n302 185
R218 VTAIL.n301 VTAIL.n300 185
R219 VTAIL.n262 VTAIL.n261 185
R220 VTAIL.n266 VTAIL.n264 185
R221 VTAIL.n295 VTAIL.n294 185
R222 VTAIL.n293 VTAIL.n292 185
R223 VTAIL.n268 VTAIL.n267 185
R224 VTAIL.n287 VTAIL.n286 185
R225 VTAIL.n285 VTAIL.n284 185
R226 VTAIL.n272 VTAIL.n271 185
R227 VTAIL.n279 VTAIL.n278 185
R228 VTAIL.n277 VTAIL.n276 185
R229 VTAIL.n247 VTAIL.n246 185
R230 VTAIL.n245 VTAIL.n244 185
R231 VTAIL.n194 VTAIL.n193 185
R232 VTAIL.n239 VTAIL.n238 185
R233 VTAIL.n237 VTAIL.n236 185
R234 VTAIL.n198 VTAIL.n197 185
R235 VTAIL.n202 VTAIL.n200 185
R236 VTAIL.n231 VTAIL.n230 185
R237 VTAIL.n229 VTAIL.n228 185
R238 VTAIL.n204 VTAIL.n203 185
R239 VTAIL.n223 VTAIL.n222 185
R240 VTAIL.n221 VTAIL.n220 185
R241 VTAIL.n208 VTAIL.n207 185
R242 VTAIL.n215 VTAIL.n214 185
R243 VTAIL.n213 VTAIL.n212 185
R244 VTAIL.n461 VTAIL.t1 149.524
R245 VTAIL.n21 VTAIL.t0 149.524
R246 VTAIL.n83 VTAIL.t12 149.524
R247 VTAIL.n147 VTAIL.t7 149.524
R248 VTAIL.n401 VTAIL.t9 149.524
R249 VTAIL.n337 VTAIL.t8 149.524
R250 VTAIL.n275 VTAIL.t2 149.524
R251 VTAIL.n211 VTAIL.t15 149.524
R252 VTAIL.n464 VTAIL.n463 104.615
R253 VTAIL.n464 VTAIL.n457 104.615
R254 VTAIL.n471 VTAIL.n457 104.615
R255 VTAIL.n472 VTAIL.n471 104.615
R256 VTAIL.n472 VTAIL.n453 104.615
R257 VTAIL.n480 VTAIL.n453 104.615
R258 VTAIL.n481 VTAIL.n480 104.615
R259 VTAIL.n482 VTAIL.n481 104.615
R260 VTAIL.n482 VTAIL.n449 104.615
R261 VTAIL.n489 VTAIL.n449 104.615
R262 VTAIL.n490 VTAIL.n489 104.615
R263 VTAIL.n490 VTAIL.n445 104.615
R264 VTAIL.n497 VTAIL.n445 104.615
R265 VTAIL.n498 VTAIL.n497 104.615
R266 VTAIL.n24 VTAIL.n23 104.615
R267 VTAIL.n24 VTAIL.n17 104.615
R268 VTAIL.n31 VTAIL.n17 104.615
R269 VTAIL.n32 VTAIL.n31 104.615
R270 VTAIL.n32 VTAIL.n13 104.615
R271 VTAIL.n40 VTAIL.n13 104.615
R272 VTAIL.n41 VTAIL.n40 104.615
R273 VTAIL.n42 VTAIL.n41 104.615
R274 VTAIL.n42 VTAIL.n9 104.615
R275 VTAIL.n49 VTAIL.n9 104.615
R276 VTAIL.n50 VTAIL.n49 104.615
R277 VTAIL.n50 VTAIL.n5 104.615
R278 VTAIL.n57 VTAIL.n5 104.615
R279 VTAIL.n58 VTAIL.n57 104.615
R280 VTAIL.n86 VTAIL.n85 104.615
R281 VTAIL.n86 VTAIL.n79 104.615
R282 VTAIL.n93 VTAIL.n79 104.615
R283 VTAIL.n94 VTAIL.n93 104.615
R284 VTAIL.n94 VTAIL.n75 104.615
R285 VTAIL.n102 VTAIL.n75 104.615
R286 VTAIL.n103 VTAIL.n102 104.615
R287 VTAIL.n104 VTAIL.n103 104.615
R288 VTAIL.n104 VTAIL.n71 104.615
R289 VTAIL.n111 VTAIL.n71 104.615
R290 VTAIL.n112 VTAIL.n111 104.615
R291 VTAIL.n112 VTAIL.n67 104.615
R292 VTAIL.n119 VTAIL.n67 104.615
R293 VTAIL.n120 VTAIL.n119 104.615
R294 VTAIL.n150 VTAIL.n149 104.615
R295 VTAIL.n150 VTAIL.n143 104.615
R296 VTAIL.n157 VTAIL.n143 104.615
R297 VTAIL.n158 VTAIL.n157 104.615
R298 VTAIL.n158 VTAIL.n139 104.615
R299 VTAIL.n166 VTAIL.n139 104.615
R300 VTAIL.n167 VTAIL.n166 104.615
R301 VTAIL.n168 VTAIL.n167 104.615
R302 VTAIL.n168 VTAIL.n135 104.615
R303 VTAIL.n175 VTAIL.n135 104.615
R304 VTAIL.n176 VTAIL.n175 104.615
R305 VTAIL.n176 VTAIL.n131 104.615
R306 VTAIL.n183 VTAIL.n131 104.615
R307 VTAIL.n184 VTAIL.n183 104.615
R308 VTAIL.n436 VTAIL.n435 104.615
R309 VTAIL.n435 VTAIL.n383 104.615
R310 VTAIL.n428 VTAIL.n383 104.615
R311 VTAIL.n428 VTAIL.n427 104.615
R312 VTAIL.n427 VTAIL.n387 104.615
R313 VTAIL.n392 VTAIL.n387 104.615
R314 VTAIL.n420 VTAIL.n392 104.615
R315 VTAIL.n420 VTAIL.n419 104.615
R316 VTAIL.n419 VTAIL.n393 104.615
R317 VTAIL.n412 VTAIL.n393 104.615
R318 VTAIL.n412 VTAIL.n411 104.615
R319 VTAIL.n411 VTAIL.n397 104.615
R320 VTAIL.n404 VTAIL.n397 104.615
R321 VTAIL.n404 VTAIL.n403 104.615
R322 VTAIL.n372 VTAIL.n371 104.615
R323 VTAIL.n371 VTAIL.n319 104.615
R324 VTAIL.n364 VTAIL.n319 104.615
R325 VTAIL.n364 VTAIL.n363 104.615
R326 VTAIL.n363 VTAIL.n323 104.615
R327 VTAIL.n328 VTAIL.n323 104.615
R328 VTAIL.n356 VTAIL.n328 104.615
R329 VTAIL.n356 VTAIL.n355 104.615
R330 VTAIL.n355 VTAIL.n329 104.615
R331 VTAIL.n348 VTAIL.n329 104.615
R332 VTAIL.n348 VTAIL.n347 104.615
R333 VTAIL.n347 VTAIL.n333 104.615
R334 VTAIL.n340 VTAIL.n333 104.615
R335 VTAIL.n340 VTAIL.n339 104.615
R336 VTAIL.n310 VTAIL.n309 104.615
R337 VTAIL.n309 VTAIL.n257 104.615
R338 VTAIL.n302 VTAIL.n257 104.615
R339 VTAIL.n302 VTAIL.n301 104.615
R340 VTAIL.n301 VTAIL.n261 104.615
R341 VTAIL.n266 VTAIL.n261 104.615
R342 VTAIL.n294 VTAIL.n266 104.615
R343 VTAIL.n294 VTAIL.n293 104.615
R344 VTAIL.n293 VTAIL.n267 104.615
R345 VTAIL.n286 VTAIL.n267 104.615
R346 VTAIL.n286 VTAIL.n285 104.615
R347 VTAIL.n285 VTAIL.n271 104.615
R348 VTAIL.n278 VTAIL.n271 104.615
R349 VTAIL.n278 VTAIL.n277 104.615
R350 VTAIL.n246 VTAIL.n245 104.615
R351 VTAIL.n245 VTAIL.n193 104.615
R352 VTAIL.n238 VTAIL.n193 104.615
R353 VTAIL.n238 VTAIL.n237 104.615
R354 VTAIL.n237 VTAIL.n197 104.615
R355 VTAIL.n202 VTAIL.n197 104.615
R356 VTAIL.n230 VTAIL.n202 104.615
R357 VTAIL.n230 VTAIL.n229 104.615
R358 VTAIL.n229 VTAIL.n203 104.615
R359 VTAIL.n222 VTAIL.n203 104.615
R360 VTAIL.n222 VTAIL.n221 104.615
R361 VTAIL.n221 VTAIL.n207 104.615
R362 VTAIL.n214 VTAIL.n207 104.615
R363 VTAIL.n214 VTAIL.n213 104.615
R364 VTAIL.n463 VTAIL.t1 52.3082
R365 VTAIL.n23 VTAIL.t0 52.3082
R366 VTAIL.n85 VTAIL.t12 52.3082
R367 VTAIL.n149 VTAIL.t7 52.3082
R368 VTAIL.n403 VTAIL.t9 52.3082
R369 VTAIL.n339 VTAIL.t8 52.3082
R370 VTAIL.n277 VTAIL.t2 52.3082
R371 VTAIL.n213 VTAIL.t15 52.3082
R372 VTAIL.n379 VTAIL.n378 45.2172
R373 VTAIL.n253 VTAIL.n252 45.2172
R374 VTAIL.n1 VTAIL.n0 45.217
R375 VTAIL.n127 VTAIL.n126 45.217
R376 VTAIL.n503 VTAIL.n502 31.9914
R377 VTAIL.n63 VTAIL.n62 31.9914
R378 VTAIL.n125 VTAIL.n124 31.9914
R379 VTAIL.n189 VTAIL.n188 31.9914
R380 VTAIL.n441 VTAIL.n440 31.9914
R381 VTAIL.n377 VTAIL.n376 31.9914
R382 VTAIL.n315 VTAIL.n314 31.9914
R383 VTAIL.n251 VTAIL.n250 31.9914
R384 VTAIL.n503 VTAIL.n441 24.4445
R385 VTAIL.n251 VTAIL.n189 24.4445
R386 VTAIL.n483 VTAIL.n450 13.1884
R387 VTAIL.n43 VTAIL.n10 13.1884
R388 VTAIL.n105 VTAIL.n72 13.1884
R389 VTAIL.n169 VTAIL.n136 13.1884
R390 VTAIL.n390 VTAIL.n388 13.1884
R391 VTAIL.n326 VTAIL.n324 13.1884
R392 VTAIL.n264 VTAIL.n262 13.1884
R393 VTAIL.n200 VTAIL.n198 13.1884
R394 VTAIL.n484 VTAIL.n452 12.8005
R395 VTAIL.n488 VTAIL.n487 12.8005
R396 VTAIL.n44 VTAIL.n12 12.8005
R397 VTAIL.n48 VTAIL.n47 12.8005
R398 VTAIL.n106 VTAIL.n74 12.8005
R399 VTAIL.n110 VTAIL.n109 12.8005
R400 VTAIL.n170 VTAIL.n138 12.8005
R401 VTAIL.n174 VTAIL.n173 12.8005
R402 VTAIL.n426 VTAIL.n425 12.8005
R403 VTAIL.n422 VTAIL.n421 12.8005
R404 VTAIL.n362 VTAIL.n361 12.8005
R405 VTAIL.n358 VTAIL.n357 12.8005
R406 VTAIL.n300 VTAIL.n299 12.8005
R407 VTAIL.n296 VTAIL.n295 12.8005
R408 VTAIL.n236 VTAIL.n235 12.8005
R409 VTAIL.n232 VTAIL.n231 12.8005
R410 VTAIL.n479 VTAIL.n478 12.0247
R411 VTAIL.n491 VTAIL.n448 12.0247
R412 VTAIL.n39 VTAIL.n38 12.0247
R413 VTAIL.n51 VTAIL.n8 12.0247
R414 VTAIL.n101 VTAIL.n100 12.0247
R415 VTAIL.n113 VTAIL.n70 12.0247
R416 VTAIL.n165 VTAIL.n164 12.0247
R417 VTAIL.n177 VTAIL.n134 12.0247
R418 VTAIL.n429 VTAIL.n386 12.0247
R419 VTAIL.n418 VTAIL.n391 12.0247
R420 VTAIL.n365 VTAIL.n322 12.0247
R421 VTAIL.n354 VTAIL.n327 12.0247
R422 VTAIL.n303 VTAIL.n260 12.0247
R423 VTAIL.n292 VTAIL.n265 12.0247
R424 VTAIL.n239 VTAIL.n196 12.0247
R425 VTAIL.n228 VTAIL.n201 12.0247
R426 VTAIL.n477 VTAIL.n454 11.249
R427 VTAIL.n492 VTAIL.n446 11.249
R428 VTAIL.n37 VTAIL.n14 11.249
R429 VTAIL.n52 VTAIL.n6 11.249
R430 VTAIL.n99 VTAIL.n76 11.249
R431 VTAIL.n114 VTAIL.n68 11.249
R432 VTAIL.n163 VTAIL.n140 11.249
R433 VTAIL.n178 VTAIL.n132 11.249
R434 VTAIL.n430 VTAIL.n384 11.249
R435 VTAIL.n417 VTAIL.n394 11.249
R436 VTAIL.n366 VTAIL.n320 11.249
R437 VTAIL.n353 VTAIL.n330 11.249
R438 VTAIL.n304 VTAIL.n258 11.249
R439 VTAIL.n291 VTAIL.n268 11.249
R440 VTAIL.n240 VTAIL.n194 11.249
R441 VTAIL.n227 VTAIL.n204 11.249
R442 VTAIL.n474 VTAIL.n473 10.4732
R443 VTAIL.n496 VTAIL.n495 10.4732
R444 VTAIL.n34 VTAIL.n33 10.4732
R445 VTAIL.n56 VTAIL.n55 10.4732
R446 VTAIL.n96 VTAIL.n95 10.4732
R447 VTAIL.n118 VTAIL.n117 10.4732
R448 VTAIL.n160 VTAIL.n159 10.4732
R449 VTAIL.n182 VTAIL.n181 10.4732
R450 VTAIL.n434 VTAIL.n433 10.4732
R451 VTAIL.n414 VTAIL.n413 10.4732
R452 VTAIL.n370 VTAIL.n369 10.4732
R453 VTAIL.n350 VTAIL.n349 10.4732
R454 VTAIL.n308 VTAIL.n307 10.4732
R455 VTAIL.n288 VTAIL.n287 10.4732
R456 VTAIL.n244 VTAIL.n243 10.4732
R457 VTAIL.n224 VTAIL.n223 10.4732
R458 VTAIL.n462 VTAIL.n461 10.2747
R459 VTAIL.n22 VTAIL.n21 10.2747
R460 VTAIL.n84 VTAIL.n83 10.2747
R461 VTAIL.n148 VTAIL.n147 10.2747
R462 VTAIL.n402 VTAIL.n401 10.2747
R463 VTAIL.n338 VTAIL.n337 10.2747
R464 VTAIL.n276 VTAIL.n275 10.2747
R465 VTAIL.n212 VTAIL.n211 10.2747
R466 VTAIL.n470 VTAIL.n456 9.69747
R467 VTAIL.n499 VTAIL.n444 9.69747
R468 VTAIL.n30 VTAIL.n16 9.69747
R469 VTAIL.n59 VTAIL.n4 9.69747
R470 VTAIL.n92 VTAIL.n78 9.69747
R471 VTAIL.n121 VTAIL.n66 9.69747
R472 VTAIL.n156 VTAIL.n142 9.69747
R473 VTAIL.n185 VTAIL.n130 9.69747
R474 VTAIL.n437 VTAIL.n382 9.69747
R475 VTAIL.n410 VTAIL.n396 9.69747
R476 VTAIL.n373 VTAIL.n318 9.69747
R477 VTAIL.n346 VTAIL.n332 9.69747
R478 VTAIL.n311 VTAIL.n256 9.69747
R479 VTAIL.n284 VTAIL.n270 9.69747
R480 VTAIL.n247 VTAIL.n192 9.69747
R481 VTAIL.n220 VTAIL.n206 9.69747
R482 VTAIL.n502 VTAIL.n501 9.45567
R483 VTAIL.n62 VTAIL.n61 9.45567
R484 VTAIL.n124 VTAIL.n123 9.45567
R485 VTAIL.n188 VTAIL.n187 9.45567
R486 VTAIL.n440 VTAIL.n439 9.45567
R487 VTAIL.n376 VTAIL.n375 9.45567
R488 VTAIL.n314 VTAIL.n313 9.45567
R489 VTAIL.n250 VTAIL.n249 9.45567
R490 VTAIL.n501 VTAIL.n500 9.3005
R491 VTAIL.n444 VTAIL.n443 9.3005
R492 VTAIL.n495 VTAIL.n494 9.3005
R493 VTAIL.n493 VTAIL.n492 9.3005
R494 VTAIL.n448 VTAIL.n447 9.3005
R495 VTAIL.n487 VTAIL.n486 9.3005
R496 VTAIL.n460 VTAIL.n459 9.3005
R497 VTAIL.n467 VTAIL.n466 9.3005
R498 VTAIL.n469 VTAIL.n468 9.3005
R499 VTAIL.n456 VTAIL.n455 9.3005
R500 VTAIL.n475 VTAIL.n474 9.3005
R501 VTAIL.n477 VTAIL.n476 9.3005
R502 VTAIL.n478 VTAIL.n451 9.3005
R503 VTAIL.n485 VTAIL.n484 9.3005
R504 VTAIL.n61 VTAIL.n60 9.3005
R505 VTAIL.n4 VTAIL.n3 9.3005
R506 VTAIL.n55 VTAIL.n54 9.3005
R507 VTAIL.n53 VTAIL.n52 9.3005
R508 VTAIL.n8 VTAIL.n7 9.3005
R509 VTAIL.n47 VTAIL.n46 9.3005
R510 VTAIL.n20 VTAIL.n19 9.3005
R511 VTAIL.n27 VTAIL.n26 9.3005
R512 VTAIL.n29 VTAIL.n28 9.3005
R513 VTAIL.n16 VTAIL.n15 9.3005
R514 VTAIL.n35 VTAIL.n34 9.3005
R515 VTAIL.n37 VTAIL.n36 9.3005
R516 VTAIL.n38 VTAIL.n11 9.3005
R517 VTAIL.n45 VTAIL.n44 9.3005
R518 VTAIL.n123 VTAIL.n122 9.3005
R519 VTAIL.n66 VTAIL.n65 9.3005
R520 VTAIL.n117 VTAIL.n116 9.3005
R521 VTAIL.n115 VTAIL.n114 9.3005
R522 VTAIL.n70 VTAIL.n69 9.3005
R523 VTAIL.n109 VTAIL.n108 9.3005
R524 VTAIL.n82 VTAIL.n81 9.3005
R525 VTAIL.n89 VTAIL.n88 9.3005
R526 VTAIL.n91 VTAIL.n90 9.3005
R527 VTAIL.n78 VTAIL.n77 9.3005
R528 VTAIL.n97 VTAIL.n96 9.3005
R529 VTAIL.n99 VTAIL.n98 9.3005
R530 VTAIL.n100 VTAIL.n73 9.3005
R531 VTAIL.n107 VTAIL.n106 9.3005
R532 VTAIL.n187 VTAIL.n186 9.3005
R533 VTAIL.n130 VTAIL.n129 9.3005
R534 VTAIL.n181 VTAIL.n180 9.3005
R535 VTAIL.n179 VTAIL.n178 9.3005
R536 VTAIL.n134 VTAIL.n133 9.3005
R537 VTAIL.n173 VTAIL.n172 9.3005
R538 VTAIL.n146 VTAIL.n145 9.3005
R539 VTAIL.n153 VTAIL.n152 9.3005
R540 VTAIL.n155 VTAIL.n154 9.3005
R541 VTAIL.n142 VTAIL.n141 9.3005
R542 VTAIL.n161 VTAIL.n160 9.3005
R543 VTAIL.n163 VTAIL.n162 9.3005
R544 VTAIL.n164 VTAIL.n137 9.3005
R545 VTAIL.n171 VTAIL.n170 9.3005
R546 VTAIL.n400 VTAIL.n399 9.3005
R547 VTAIL.n407 VTAIL.n406 9.3005
R548 VTAIL.n409 VTAIL.n408 9.3005
R549 VTAIL.n396 VTAIL.n395 9.3005
R550 VTAIL.n415 VTAIL.n414 9.3005
R551 VTAIL.n417 VTAIL.n416 9.3005
R552 VTAIL.n391 VTAIL.n389 9.3005
R553 VTAIL.n423 VTAIL.n422 9.3005
R554 VTAIL.n439 VTAIL.n438 9.3005
R555 VTAIL.n382 VTAIL.n381 9.3005
R556 VTAIL.n433 VTAIL.n432 9.3005
R557 VTAIL.n431 VTAIL.n430 9.3005
R558 VTAIL.n386 VTAIL.n385 9.3005
R559 VTAIL.n425 VTAIL.n424 9.3005
R560 VTAIL.n336 VTAIL.n335 9.3005
R561 VTAIL.n343 VTAIL.n342 9.3005
R562 VTAIL.n345 VTAIL.n344 9.3005
R563 VTAIL.n332 VTAIL.n331 9.3005
R564 VTAIL.n351 VTAIL.n350 9.3005
R565 VTAIL.n353 VTAIL.n352 9.3005
R566 VTAIL.n327 VTAIL.n325 9.3005
R567 VTAIL.n359 VTAIL.n358 9.3005
R568 VTAIL.n375 VTAIL.n374 9.3005
R569 VTAIL.n318 VTAIL.n317 9.3005
R570 VTAIL.n369 VTAIL.n368 9.3005
R571 VTAIL.n367 VTAIL.n366 9.3005
R572 VTAIL.n322 VTAIL.n321 9.3005
R573 VTAIL.n361 VTAIL.n360 9.3005
R574 VTAIL.n274 VTAIL.n273 9.3005
R575 VTAIL.n281 VTAIL.n280 9.3005
R576 VTAIL.n283 VTAIL.n282 9.3005
R577 VTAIL.n270 VTAIL.n269 9.3005
R578 VTAIL.n289 VTAIL.n288 9.3005
R579 VTAIL.n291 VTAIL.n290 9.3005
R580 VTAIL.n265 VTAIL.n263 9.3005
R581 VTAIL.n297 VTAIL.n296 9.3005
R582 VTAIL.n313 VTAIL.n312 9.3005
R583 VTAIL.n256 VTAIL.n255 9.3005
R584 VTAIL.n307 VTAIL.n306 9.3005
R585 VTAIL.n305 VTAIL.n304 9.3005
R586 VTAIL.n260 VTAIL.n259 9.3005
R587 VTAIL.n299 VTAIL.n298 9.3005
R588 VTAIL.n210 VTAIL.n209 9.3005
R589 VTAIL.n217 VTAIL.n216 9.3005
R590 VTAIL.n219 VTAIL.n218 9.3005
R591 VTAIL.n206 VTAIL.n205 9.3005
R592 VTAIL.n225 VTAIL.n224 9.3005
R593 VTAIL.n227 VTAIL.n226 9.3005
R594 VTAIL.n201 VTAIL.n199 9.3005
R595 VTAIL.n233 VTAIL.n232 9.3005
R596 VTAIL.n249 VTAIL.n248 9.3005
R597 VTAIL.n192 VTAIL.n191 9.3005
R598 VTAIL.n243 VTAIL.n242 9.3005
R599 VTAIL.n241 VTAIL.n240 9.3005
R600 VTAIL.n196 VTAIL.n195 9.3005
R601 VTAIL.n235 VTAIL.n234 9.3005
R602 VTAIL.n469 VTAIL.n458 8.92171
R603 VTAIL.n500 VTAIL.n442 8.92171
R604 VTAIL.n29 VTAIL.n18 8.92171
R605 VTAIL.n60 VTAIL.n2 8.92171
R606 VTAIL.n91 VTAIL.n80 8.92171
R607 VTAIL.n122 VTAIL.n64 8.92171
R608 VTAIL.n155 VTAIL.n144 8.92171
R609 VTAIL.n186 VTAIL.n128 8.92171
R610 VTAIL.n438 VTAIL.n380 8.92171
R611 VTAIL.n409 VTAIL.n398 8.92171
R612 VTAIL.n374 VTAIL.n316 8.92171
R613 VTAIL.n345 VTAIL.n334 8.92171
R614 VTAIL.n312 VTAIL.n254 8.92171
R615 VTAIL.n283 VTAIL.n272 8.92171
R616 VTAIL.n248 VTAIL.n190 8.92171
R617 VTAIL.n219 VTAIL.n208 8.92171
R618 VTAIL.n466 VTAIL.n465 8.14595
R619 VTAIL.n26 VTAIL.n25 8.14595
R620 VTAIL.n88 VTAIL.n87 8.14595
R621 VTAIL.n152 VTAIL.n151 8.14595
R622 VTAIL.n406 VTAIL.n405 8.14595
R623 VTAIL.n342 VTAIL.n341 8.14595
R624 VTAIL.n280 VTAIL.n279 8.14595
R625 VTAIL.n216 VTAIL.n215 8.14595
R626 VTAIL.n462 VTAIL.n460 7.3702
R627 VTAIL.n22 VTAIL.n20 7.3702
R628 VTAIL.n84 VTAIL.n82 7.3702
R629 VTAIL.n148 VTAIL.n146 7.3702
R630 VTAIL.n402 VTAIL.n400 7.3702
R631 VTAIL.n338 VTAIL.n336 7.3702
R632 VTAIL.n276 VTAIL.n274 7.3702
R633 VTAIL.n212 VTAIL.n210 7.3702
R634 VTAIL.n465 VTAIL.n460 5.81868
R635 VTAIL.n25 VTAIL.n20 5.81868
R636 VTAIL.n87 VTAIL.n82 5.81868
R637 VTAIL.n151 VTAIL.n146 5.81868
R638 VTAIL.n405 VTAIL.n400 5.81868
R639 VTAIL.n341 VTAIL.n336 5.81868
R640 VTAIL.n279 VTAIL.n274 5.81868
R641 VTAIL.n215 VTAIL.n210 5.81868
R642 VTAIL.n466 VTAIL.n458 5.04292
R643 VTAIL.n502 VTAIL.n442 5.04292
R644 VTAIL.n26 VTAIL.n18 5.04292
R645 VTAIL.n62 VTAIL.n2 5.04292
R646 VTAIL.n88 VTAIL.n80 5.04292
R647 VTAIL.n124 VTAIL.n64 5.04292
R648 VTAIL.n152 VTAIL.n144 5.04292
R649 VTAIL.n188 VTAIL.n128 5.04292
R650 VTAIL.n440 VTAIL.n380 5.04292
R651 VTAIL.n406 VTAIL.n398 5.04292
R652 VTAIL.n376 VTAIL.n316 5.04292
R653 VTAIL.n342 VTAIL.n334 5.04292
R654 VTAIL.n314 VTAIL.n254 5.04292
R655 VTAIL.n280 VTAIL.n272 5.04292
R656 VTAIL.n250 VTAIL.n190 5.04292
R657 VTAIL.n216 VTAIL.n208 5.04292
R658 VTAIL.n470 VTAIL.n469 4.26717
R659 VTAIL.n500 VTAIL.n499 4.26717
R660 VTAIL.n30 VTAIL.n29 4.26717
R661 VTAIL.n60 VTAIL.n59 4.26717
R662 VTAIL.n92 VTAIL.n91 4.26717
R663 VTAIL.n122 VTAIL.n121 4.26717
R664 VTAIL.n156 VTAIL.n155 4.26717
R665 VTAIL.n186 VTAIL.n185 4.26717
R666 VTAIL.n438 VTAIL.n437 4.26717
R667 VTAIL.n410 VTAIL.n409 4.26717
R668 VTAIL.n374 VTAIL.n373 4.26717
R669 VTAIL.n346 VTAIL.n345 4.26717
R670 VTAIL.n312 VTAIL.n311 4.26717
R671 VTAIL.n284 VTAIL.n283 4.26717
R672 VTAIL.n248 VTAIL.n247 4.26717
R673 VTAIL.n220 VTAIL.n219 4.26717
R674 VTAIL.n473 VTAIL.n456 3.49141
R675 VTAIL.n496 VTAIL.n444 3.49141
R676 VTAIL.n33 VTAIL.n16 3.49141
R677 VTAIL.n56 VTAIL.n4 3.49141
R678 VTAIL.n95 VTAIL.n78 3.49141
R679 VTAIL.n118 VTAIL.n66 3.49141
R680 VTAIL.n159 VTAIL.n142 3.49141
R681 VTAIL.n182 VTAIL.n130 3.49141
R682 VTAIL.n434 VTAIL.n382 3.49141
R683 VTAIL.n413 VTAIL.n396 3.49141
R684 VTAIL.n370 VTAIL.n318 3.49141
R685 VTAIL.n349 VTAIL.n332 3.49141
R686 VTAIL.n308 VTAIL.n256 3.49141
R687 VTAIL.n287 VTAIL.n270 3.49141
R688 VTAIL.n244 VTAIL.n192 3.49141
R689 VTAIL.n223 VTAIL.n206 3.49141
R690 VTAIL.n461 VTAIL.n459 2.84303
R691 VTAIL.n21 VTAIL.n19 2.84303
R692 VTAIL.n83 VTAIL.n81 2.84303
R693 VTAIL.n147 VTAIL.n145 2.84303
R694 VTAIL.n401 VTAIL.n399 2.84303
R695 VTAIL.n337 VTAIL.n335 2.84303
R696 VTAIL.n275 VTAIL.n273 2.84303
R697 VTAIL.n211 VTAIL.n209 2.84303
R698 VTAIL.n474 VTAIL.n454 2.71565
R699 VTAIL.n495 VTAIL.n446 2.71565
R700 VTAIL.n34 VTAIL.n14 2.71565
R701 VTAIL.n55 VTAIL.n6 2.71565
R702 VTAIL.n96 VTAIL.n76 2.71565
R703 VTAIL.n117 VTAIL.n68 2.71565
R704 VTAIL.n160 VTAIL.n140 2.71565
R705 VTAIL.n181 VTAIL.n132 2.71565
R706 VTAIL.n433 VTAIL.n384 2.71565
R707 VTAIL.n414 VTAIL.n394 2.71565
R708 VTAIL.n369 VTAIL.n320 2.71565
R709 VTAIL.n350 VTAIL.n330 2.71565
R710 VTAIL.n307 VTAIL.n258 2.71565
R711 VTAIL.n288 VTAIL.n268 2.71565
R712 VTAIL.n243 VTAIL.n194 2.71565
R713 VTAIL.n224 VTAIL.n204 2.71565
R714 VTAIL.n253 VTAIL.n251 2.25912
R715 VTAIL.n315 VTAIL.n253 2.25912
R716 VTAIL.n379 VTAIL.n377 2.25912
R717 VTAIL.n441 VTAIL.n379 2.25912
R718 VTAIL.n189 VTAIL.n127 2.25912
R719 VTAIL.n127 VTAIL.n125 2.25912
R720 VTAIL.n63 VTAIL.n1 2.25912
R721 VTAIL VTAIL.n503 2.20093
R722 VTAIL.n479 VTAIL.n477 1.93989
R723 VTAIL.n492 VTAIL.n491 1.93989
R724 VTAIL.n39 VTAIL.n37 1.93989
R725 VTAIL.n52 VTAIL.n51 1.93989
R726 VTAIL.n101 VTAIL.n99 1.93989
R727 VTAIL.n114 VTAIL.n113 1.93989
R728 VTAIL.n165 VTAIL.n163 1.93989
R729 VTAIL.n178 VTAIL.n177 1.93989
R730 VTAIL.n430 VTAIL.n429 1.93989
R731 VTAIL.n418 VTAIL.n417 1.93989
R732 VTAIL.n366 VTAIL.n365 1.93989
R733 VTAIL.n354 VTAIL.n353 1.93989
R734 VTAIL.n304 VTAIL.n303 1.93989
R735 VTAIL.n292 VTAIL.n291 1.93989
R736 VTAIL.n240 VTAIL.n239 1.93989
R737 VTAIL.n228 VTAIL.n227 1.93989
R738 VTAIL.n0 VTAIL.t4 1.73887
R739 VTAIL.n0 VTAIL.t3 1.73887
R740 VTAIL.n126 VTAIL.t10 1.73887
R741 VTAIL.n126 VTAIL.t6 1.73887
R742 VTAIL.n378 VTAIL.t11 1.73887
R743 VTAIL.n378 VTAIL.t13 1.73887
R744 VTAIL.n252 VTAIL.t5 1.73887
R745 VTAIL.n252 VTAIL.t14 1.73887
R746 VTAIL.n478 VTAIL.n452 1.16414
R747 VTAIL.n488 VTAIL.n448 1.16414
R748 VTAIL.n38 VTAIL.n12 1.16414
R749 VTAIL.n48 VTAIL.n8 1.16414
R750 VTAIL.n100 VTAIL.n74 1.16414
R751 VTAIL.n110 VTAIL.n70 1.16414
R752 VTAIL.n164 VTAIL.n138 1.16414
R753 VTAIL.n174 VTAIL.n134 1.16414
R754 VTAIL.n426 VTAIL.n386 1.16414
R755 VTAIL.n421 VTAIL.n391 1.16414
R756 VTAIL.n362 VTAIL.n322 1.16414
R757 VTAIL.n357 VTAIL.n327 1.16414
R758 VTAIL.n300 VTAIL.n260 1.16414
R759 VTAIL.n295 VTAIL.n265 1.16414
R760 VTAIL.n236 VTAIL.n196 1.16414
R761 VTAIL.n231 VTAIL.n201 1.16414
R762 VTAIL.n377 VTAIL.n315 0.470328
R763 VTAIL.n125 VTAIL.n63 0.470328
R764 VTAIL.n484 VTAIL.n483 0.388379
R765 VTAIL.n487 VTAIL.n450 0.388379
R766 VTAIL.n44 VTAIL.n43 0.388379
R767 VTAIL.n47 VTAIL.n10 0.388379
R768 VTAIL.n106 VTAIL.n105 0.388379
R769 VTAIL.n109 VTAIL.n72 0.388379
R770 VTAIL.n170 VTAIL.n169 0.388379
R771 VTAIL.n173 VTAIL.n136 0.388379
R772 VTAIL.n425 VTAIL.n388 0.388379
R773 VTAIL.n422 VTAIL.n390 0.388379
R774 VTAIL.n361 VTAIL.n324 0.388379
R775 VTAIL.n358 VTAIL.n326 0.388379
R776 VTAIL.n299 VTAIL.n262 0.388379
R777 VTAIL.n296 VTAIL.n264 0.388379
R778 VTAIL.n235 VTAIL.n198 0.388379
R779 VTAIL.n232 VTAIL.n200 0.388379
R780 VTAIL.n467 VTAIL.n459 0.155672
R781 VTAIL.n468 VTAIL.n467 0.155672
R782 VTAIL.n468 VTAIL.n455 0.155672
R783 VTAIL.n475 VTAIL.n455 0.155672
R784 VTAIL.n476 VTAIL.n475 0.155672
R785 VTAIL.n476 VTAIL.n451 0.155672
R786 VTAIL.n485 VTAIL.n451 0.155672
R787 VTAIL.n486 VTAIL.n485 0.155672
R788 VTAIL.n486 VTAIL.n447 0.155672
R789 VTAIL.n493 VTAIL.n447 0.155672
R790 VTAIL.n494 VTAIL.n493 0.155672
R791 VTAIL.n494 VTAIL.n443 0.155672
R792 VTAIL.n501 VTAIL.n443 0.155672
R793 VTAIL.n27 VTAIL.n19 0.155672
R794 VTAIL.n28 VTAIL.n27 0.155672
R795 VTAIL.n28 VTAIL.n15 0.155672
R796 VTAIL.n35 VTAIL.n15 0.155672
R797 VTAIL.n36 VTAIL.n35 0.155672
R798 VTAIL.n36 VTAIL.n11 0.155672
R799 VTAIL.n45 VTAIL.n11 0.155672
R800 VTAIL.n46 VTAIL.n45 0.155672
R801 VTAIL.n46 VTAIL.n7 0.155672
R802 VTAIL.n53 VTAIL.n7 0.155672
R803 VTAIL.n54 VTAIL.n53 0.155672
R804 VTAIL.n54 VTAIL.n3 0.155672
R805 VTAIL.n61 VTAIL.n3 0.155672
R806 VTAIL.n89 VTAIL.n81 0.155672
R807 VTAIL.n90 VTAIL.n89 0.155672
R808 VTAIL.n90 VTAIL.n77 0.155672
R809 VTAIL.n97 VTAIL.n77 0.155672
R810 VTAIL.n98 VTAIL.n97 0.155672
R811 VTAIL.n98 VTAIL.n73 0.155672
R812 VTAIL.n107 VTAIL.n73 0.155672
R813 VTAIL.n108 VTAIL.n107 0.155672
R814 VTAIL.n108 VTAIL.n69 0.155672
R815 VTAIL.n115 VTAIL.n69 0.155672
R816 VTAIL.n116 VTAIL.n115 0.155672
R817 VTAIL.n116 VTAIL.n65 0.155672
R818 VTAIL.n123 VTAIL.n65 0.155672
R819 VTAIL.n153 VTAIL.n145 0.155672
R820 VTAIL.n154 VTAIL.n153 0.155672
R821 VTAIL.n154 VTAIL.n141 0.155672
R822 VTAIL.n161 VTAIL.n141 0.155672
R823 VTAIL.n162 VTAIL.n161 0.155672
R824 VTAIL.n162 VTAIL.n137 0.155672
R825 VTAIL.n171 VTAIL.n137 0.155672
R826 VTAIL.n172 VTAIL.n171 0.155672
R827 VTAIL.n172 VTAIL.n133 0.155672
R828 VTAIL.n179 VTAIL.n133 0.155672
R829 VTAIL.n180 VTAIL.n179 0.155672
R830 VTAIL.n180 VTAIL.n129 0.155672
R831 VTAIL.n187 VTAIL.n129 0.155672
R832 VTAIL.n439 VTAIL.n381 0.155672
R833 VTAIL.n432 VTAIL.n381 0.155672
R834 VTAIL.n432 VTAIL.n431 0.155672
R835 VTAIL.n431 VTAIL.n385 0.155672
R836 VTAIL.n424 VTAIL.n385 0.155672
R837 VTAIL.n424 VTAIL.n423 0.155672
R838 VTAIL.n423 VTAIL.n389 0.155672
R839 VTAIL.n416 VTAIL.n389 0.155672
R840 VTAIL.n416 VTAIL.n415 0.155672
R841 VTAIL.n415 VTAIL.n395 0.155672
R842 VTAIL.n408 VTAIL.n395 0.155672
R843 VTAIL.n408 VTAIL.n407 0.155672
R844 VTAIL.n407 VTAIL.n399 0.155672
R845 VTAIL.n375 VTAIL.n317 0.155672
R846 VTAIL.n368 VTAIL.n317 0.155672
R847 VTAIL.n368 VTAIL.n367 0.155672
R848 VTAIL.n367 VTAIL.n321 0.155672
R849 VTAIL.n360 VTAIL.n321 0.155672
R850 VTAIL.n360 VTAIL.n359 0.155672
R851 VTAIL.n359 VTAIL.n325 0.155672
R852 VTAIL.n352 VTAIL.n325 0.155672
R853 VTAIL.n352 VTAIL.n351 0.155672
R854 VTAIL.n351 VTAIL.n331 0.155672
R855 VTAIL.n344 VTAIL.n331 0.155672
R856 VTAIL.n344 VTAIL.n343 0.155672
R857 VTAIL.n343 VTAIL.n335 0.155672
R858 VTAIL.n313 VTAIL.n255 0.155672
R859 VTAIL.n306 VTAIL.n255 0.155672
R860 VTAIL.n306 VTAIL.n305 0.155672
R861 VTAIL.n305 VTAIL.n259 0.155672
R862 VTAIL.n298 VTAIL.n259 0.155672
R863 VTAIL.n298 VTAIL.n297 0.155672
R864 VTAIL.n297 VTAIL.n263 0.155672
R865 VTAIL.n290 VTAIL.n263 0.155672
R866 VTAIL.n290 VTAIL.n289 0.155672
R867 VTAIL.n289 VTAIL.n269 0.155672
R868 VTAIL.n282 VTAIL.n269 0.155672
R869 VTAIL.n282 VTAIL.n281 0.155672
R870 VTAIL.n281 VTAIL.n273 0.155672
R871 VTAIL.n249 VTAIL.n191 0.155672
R872 VTAIL.n242 VTAIL.n191 0.155672
R873 VTAIL.n242 VTAIL.n241 0.155672
R874 VTAIL.n241 VTAIL.n195 0.155672
R875 VTAIL.n234 VTAIL.n195 0.155672
R876 VTAIL.n234 VTAIL.n233 0.155672
R877 VTAIL.n233 VTAIL.n199 0.155672
R878 VTAIL.n226 VTAIL.n199 0.155672
R879 VTAIL.n226 VTAIL.n225 0.155672
R880 VTAIL.n225 VTAIL.n205 0.155672
R881 VTAIL.n218 VTAIL.n205 0.155672
R882 VTAIL.n218 VTAIL.n217 0.155672
R883 VTAIL.n217 VTAIL.n209 0.155672
R884 VTAIL VTAIL.n1 0.0586897
R885 B.n652 B.n135 585
R886 B.n135 B.n86 585
R887 B.n654 B.n653 585
R888 B.n656 B.n134 585
R889 B.n659 B.n658 585
R890 B.n660 B.n133 585
R891 B.n662 B.n661 585
R892 B.n664 B.n132 585
R893 B.n667 B.n666 585
R894 B.n668 B.n131 585
R895 B.n670 B.n669 585
R896 B.n672 B.n130 585
R897 B.n675 B.n674 585
R898 B.n676 B.n129 585
R899 B.n678 B.n677 585
R900 B.n680 B.n128 585
R901 B.n683 B.n682 585
R902 B.n684 B.n127 585
R903 B.n686 B.n685 585
R904 B.n688 B.n126 585
R905 B.n691 B.n690 585
R906 B.n692 B.n125 585
R907 B.n694 B.n693 585
R908 B.n696 B.n124 585
R909 B.n699 B.n698 585
R910 B.n700 B.n123 585
R911 B.n702 B.n701 585
R912 B.n704 B.n122 585
R913 B.n707 B.n706 585
R914 B.n708 B.n121 585
R915 B.n710 B.n709 585
R916 B.n712 B.n120 585
R917 B.n715 B.n714 585
R918 B.n716 B.n119 585
R919 B.n718 B.n717 585
R920 B.n720 B.n118 585
R921 B.n723 B.n722 585
R922 B.n724 B.n117 585
R923 B.n726 B.n725 585
R924 B.n728 B.n116 585
R925 B.n731 B.n730 585
R926 B.n733 B.n113 585
R927 B.n735 B.n734 585
R928 B.n737 B.n112 585
R929 B.n740 B.n739 585
R930 B.n741 B.n111 585
R931 B.n743 B.n742 585
R932 B.n745 B.n110 585
R933 B.n748 B.n747 585
R934 B.n749 B.n107 585
R935 B.n752 B.n751 585
R936 B.n754 B.n106 585
R937 B.n757 B.n756 585
R938 B.n758 B.n105 585
R939 B.n760 B.n759 585
R940 B.n762 B.n104 585
R941 B.n765 B.n764 585
R942 B.n766 B.n103 585
R943 B.n768 B.n767 585
R944 B.n770 B.n102 585
R945 B.n773 B.n772 585
R946 B.n774 B.n101 585
R947 B.n776 B.n775 585
R948 B.n778 B.n100 585
R949 B.n781 B.n780 585
R950 B.n782 B.n99 585
R951 B.n784 B.n783 585
R952 B.n786 B.n98 585
R953 B.n789 B.n788 585
R954 B.n790 B.n97 585
R955 B.n792 B.n791 585
R956 B.n794 B.n96 585
R957 B.n797 B.n796 585
R958 B.n798 B.n95 585
R959 B.n800 B.n799 585
R960 B.n802 B.n94 585
R961 B.n805 B.n804 585
R962 B.n806 B.n93 585
R963 B.n808 B.n807 585
R964 B.n810 B.n92 585
R965 B.n813 B.n812 585
R966 B.n814 B.n91 585
R967 B.n816 B.n815 585
R968 B.n818 B.n90 585
R969 B.n821 B.n820 585
R970 B.n822 B.n89 585
R971 B.n824 B.n823 585
R972 B.n826 B.n88 585
R973 B.n829 B.n828 585
R974 B.n830 B.n87 585
R975 B.n651 B.n85 585
R976 B.n833 B.n85 585
R977 B.n650 B.n84 585
R978 B.n834 B.n84 585
R979 B.n649 B.n83 585
R980 B.n835 B.n83 585
R981 B.n648 B.n647 585
R982 B.n647 B.n79 585
R983 B.n646 B.n78 585
R984 B.n841 B.n78 585
R985 B.n645 B.n77 585
R986 B.n842 B.n77 585
R987 B.n644 B.n76 585
R988 B.n843 B.n76 585
R989 B.n643 B.n642 585
R990 B.n642 B.n75 585
R991 B.n641 B.n71 585
R992 B.n849 B.n71 585
R993 B.n640 B.n70 585
R994 B.n850 B.n70 585
R995 B.n639 B.n69 585
R996 B.n851 B.n69 585
R997 B.n638 B.n637 585
R998 B.n637 B.n65 585
R999 B.n636 B.n64 585
R1000 B.n857 B.n64 585
R1001 B.n635 B.n63 585
R1002 B.n858 B.n63 585
R1003 B.n634 B.n62 585
R1004 B.n859 B.n62 585
R1005 B.n633 B.n632 585
R1006 B.n632 B.n58 585
R1007 B.n631 B.n57 585
R1008 B.n865 B.n57 585
R1009 B.n630 B.n56 585
R1010 B.n866 B.n56 585
R1011 B.n629 B.n55 585
R1012 B.n867 B.n55 585
R1013 B.n628 B.n627 585
R1014 B.n627 B.n51 585
R1015 B.n626 B.n50 585
R1016 B.n873 B.n50 585
R1017 B.n625 B.n49 585
R1018 B.n874 B.n49 585
R1019 B.n624 B.n48 585
R1020 B.n875 B.n48 585
R1021 B.n623 B.n622 585
R1022 B.n622 B.n44 585
R1023 B.n621 B.n43 585
R1024 B.n881 B.n43 585
R1025 B.n620 B.n42 585
R1026 B.n882 B.n42 585
R1027 B.n619 B.n41 585
R1028 B.n883 B.n41 585
R1029 B.n618 B.n617 585
R1030 B.n617 B.n37 585
R1031 B.n616 B.n36 585
R1032 B.n889 B.n36 585
R1033 B.n615 B.n35 585
R1034 B.n890 B.n35 585
R1035 B.n614 B.n34 585
R1036 B.n891 B.n34 585
R1037 B.n613 B.n612 585
R1038 B.n612 B.n30 585
R1039 B.n611 B.n29 585
R1040 B.n897 B.n29 585
R1041 B.n610 B.n28 585
R1042 B.n898 B.n28 585
R1043 B.n609 B.n27 585
R1044 B.n899 B.n27 585
R1045 B.n608 B.n607 585
R1046 B.n607 B.n23 585
R1047 B.n606 B.n22 585
R1048 B.n905 B.n22 585
R1049 B.n605 B.n21 585
R1050 B.n906 B.n21 585
R1051 B.n604 B.n20 585
R1052 B.n907 B.n20 585
R1053 B.n603 B.n602 585
R1054 B.n602 B.n16 585
R1055 B.n601 B.n15 585
R1056 B.n913 B.n15 585
R1057 B.n600 B.n14 585
R1058 B.n914 B.n14 585
R1059 B.n599 B.n13 585
R1060 B.n915 B.n13 585
R1061 B.n598 B.n597 585
R1062 B.n597 B.n12 585
R1063 B.n596 B.n595 585
R1064 B.n596 B.n8 585
R1065 B.n594 B.n7 585
R1066 B.n922 B.n7 585
R1067 B.n593 B.n6 585
R1068 B.n923 B.n6 585
R1069 B.n592 B.n5 585
R1070 B.n924 B.n5 585
R1071 B.n591 B.n590 585
R1072 B.n590 B.n4 585
R1073 B.n589 B.n136 585
R1074 B.n589 B.n588 585
R1075 B.n579 B.n137 585
R1076 B.n138 B.n137 585
R1077 B.n581 B.n580 585
R1078 B.n582 B.n581 585
R1079 B.n578 B.n142 585
R1080 B.n146 B.n142 585
R1081 B.n577 B.n576 585
R1082 B.n576 B.n575 585
R1083 B.n144 B.n143 585
R1084 B.n145 B.n144 585
R1085 B.n568 B.n567 585
R1086 B.n569 B.n568 585
R1087 B.n566 B.n151 585
R1088 B.n151 B.n150 585
R1089 B.n565 B.n564 585
R1090 B.n564 B.n563 585
R1091 B.n153 B.n152 585
R1092 B.n154 B.n153 585
R1093 B.n556 B.n555 585
R1094 B.n557 B.n556 585
R1095 B.n554 B.n158 585
R1096 B.n162 B.n158 585
R1097 B.n553 B.n552 585
R1098 B.n552 B.n551 585
R1099 B.n160 B.n159 585
R1100 B.n161 B.n160 585
R1101 B.n544 B.n543 585
R1102 B.n545 B.n544 585
R1103 B.n542 B.n167 585
R1104 B.n167 B.n166 585
R1105 B.n541 B.n540 585
R1106 B.n540 B.n539 585
R1107 B.n169 B.n168 585
R1108 B.n170 B.n169 585
R1109 B.n532 B.n531 585
R1110 B.n533 B.n532 585
R1111 B.n530 B.n174 585
R1112 B.n178 B.n174 585
R1113 B.n529 B.n528 585
R1114 B.n528 B.n527 585
R1115 B.n176 B.n175 585
R1116 B.n177 B.n176 585
R1117 B.n520 B.n519 585
R1118 B.n521 B.n520 585
R1119 B.n518 B.n183 585
R1120 B.n183 B.n182 585
R1121 B.n517 B.n516 585
R1122 B.n516 B.n515 585
R1123 B.n185 B.n184 585
R1124 B.n186 B.n185 585
R1125 B.n508 B.n507 585
R1126 B.n509 B.n508 585
R1127 B.n506 B.n190 585
R1128 B.n194 B.n190 585
R1129 B.n505 B.n504 585
R1130 B.n504 B.n503 585
R1131 B.n192 B.n191 585
R1132 B.n193 B.n192 585
R1133 B.n496 B.n495 585
R1134 B.n497 B.n496 585
R1135 B.n494 B.n199 585
R1136 B.n199 B.n198 585
R1137 B.n493 B.n492 585
R1138 B.n492 B.n491 585
R1139 B.n201 B.n200 585
R1140 B.n202 B.n201 585
R1141 B.n484 B.n483 585
R1142 B.n485 B.n484 585
R1143 B.n482 B.n207 585
R1144 B.n207 B.n206 585
R1145 B.n481 B.n480 585
R1146 B.n480 B.n479 585
R1147 B.n209 B.n208 585
R1148 B.n472 B.n209 585
R1149 B.n471 B.n470 585
R1150 B.n473 B.n471 585
R1151 B.n469 B.n214 585
R1152 B.n214 B.n213 585
R1153 B.n468 B.n467 585
R1154 B.n467 B.n466 585
R1155 B.n216 B.n215 585
R1156 B.n217 B.n216 585
R1157 B.n459 B.n458 585
R1158 B.n460 B.n459 585
R1159 B.n457 B.n222 585
R1160 B.n222 B.n221 585
R1161 B.n456 B.n455 585
R1162 B.n455 B.n454 585
R1163 B.n451 B.n226 585
R1164 B.n450 B.n449 585
R1165 B.n447 B.n227 585
R1166 B.n447 B.n225 585
R1167 B.n446 B.n445 585
R1168 B.n444 B.n443 585
R1169 B.n442 B.n229 585
R1170 B.n440 B.n439 585
R1171 B.n438 B.n230 585
R1172 B.n437 B.n436 585
R1173 B.n434 B.n231 585
R1174 B.n432 B.n431 585
R1175 B.n430 B.n232 585
R1176 B.n429 B.n428 585
R1177 B.n426 B.n233 585
R1178 B.n424 B.n423 585
R1179 B.n422 B.n234 585
R1180 B.n421 B.n420 585
R1181 B.n418 B.n235 585
R1182 B.n416 B.n415 585
R1183 B.n414 B.n236 585
R1184 B.n413 B.n412 585
R1185 B.n410 B.n237 585
R1186 B.n408 B.n407 585
R1187 B.n406 B.n238 585
R1188 B.n405 B.n404 585
R1189 B.n402 B.n239 585
R1190 B.n400 B.n399 585
R1191 B.n398 B.n240 585
R1192 B.n397 B.n396 585
R1193 B.n394 B.n241 585
R1194 B.n392 B.n391 585
R1195 B.n390 B.n242 585
R1196 B.n389 B.n388 585
R1197 B.n386 B.n243 585
R1198 B.n384 B.n383 585
R1199 B.n382 B.n244 585
R1200 B.n381 B.n380 585
R1201 B.n378 B.n245 585
R1202 B.n376 B.n375 585
R1203 B.n374 B.n246 585
R1204 B.n372 B.n371 585
R1205 B.n369 B.n249 585
R1206 B.n367 B.n366 585
R1207 B.n365 B.n250 585
R1208 B.n364 B.n363 585
R1209 B.n361 B.n251 585
R1210 B.n359 B.n358 585
R1211 B.n357 B.n252 585
R1212 B.n356 B.n355 585
R1213 B.n353 B.n352 585
R1214 B.n351 B.n350 585
R1215 B.n349 B.n257 585
R1216 B.n347 B.n346 585
R1217 B.n345 B.n258 585
R1218 B.n344 B.n343 585
R1219 B.n341 B.n259 585
R1220 B.n339 B.n338 585
R1221 B.n337 B.n260 585
R1222 B.n336 B.n335 585
R1223 B.n333 B.n261 585
R1224 B.n331 B.n330 585
R1225 B.n329 B.n262 585
R1226 B.n328 B.n327 585
R1227 B.n325 B.n263 585
R1228 B.n323 B.n322 585
R1229 B.n321 B.n264 585
R1230 B.n320 B.n319 585
R1231 B.n317 B.n265 585
R1232 B.n315 B.n314 585
R1233 B.n313 B.n266 585
R1234 B.n312 B.n311 585
R1235 B.n309 B.n267 585
R1236 B.n307 B.n306 585
R1237 B.n305 B.n268 585
R1238 B.n304 B.n303 585
R1239 B.n301 B.n269 585
R1240 B.n299 B.n298 585
R1241 B.n297 B.n270 585
R1242 B.n296 B.n295 585
R1243 B.n293 B.n271 585
R1244 B.n291 B.n290 585
R1245 B.n289 B.n272 585
R1246 B.n288 B.n287 585
R1247 B.n285 B.n273 585
R1248 B.n283 B.n282 585
R1249 B.n281 B.n274 585
R1250 B.n280 B.n279 585
R1251 B.n277 B.n275 585
R1252 B.n224 B.n223 585
R1253 B.n453 B.n452 585
R1254 B.n454 B.n453 585
R1255 B.n220 B.n219 585
R1256 B.n221 B.n220 585
R1257 B.n462 B.n461 585
R1258 B.n461 B.n460 585
R1259 B.n463 B.n218 585
R1260 B.n218 B.n217 585
R1261 B.n465 B.n464 585
R1262 B.n466 B.n465 585
R1263 B.n212 B.n211 585
R1264 B.n213 B.n212 585
R1265 B.n475 B.n474 585
R1266 B.n474 B.n473 585
R1267 B.n476 B.n210 585
R1268 B.n472 B.n210 585
R1269 B.n478 B.n477 585
R1270 B.n479 B.n478 585
R1271 B.n205 B.n204 585
R1272 B.n206 B.n205 585
R1273 B.n487 B.n486 585
R1274 B.n486 B.n485 585
R1275 B.n488 B.n203 585
R1276 B.n203 B.n202 585
R1277 B.n490 B.n489 585
R1278 B.n491 B.n490 585
R1279 B.n197 B.n196 585
R1280 B.n198 B.n197 585
R1281 B.n499 B.n498 585
R1282 B.n498 B.n497 585
R1283 B.n500 B.n195 585
R1284 B.n195 B.n193 585
R1285 B.n502 B.n501 585
R1286 B.n503 B.n502 585
R1287 B.n189 B.n188 585
R1288 B.n194 B.n189 585
R1289 B.n511 B.n510 585
R1290 B.n510 B.n509 585
R1291 B.n512 B.n187 585
R1292 B.n187 B.n186 585
R1293 B.n514 B.n513 585
R1294 B.n515 B.n514 585
R1295 B.n181 B.n180 585
R1296 B.n182 B.n181 585
R1297 B.n523 B.n522 585
R1298 B.n522 B.n521 585
R1299 B.n524 B.n179 585
R1300 B.n179 B.n177 585
R1301 B.n526 B.n525 585
R1302 B.n527 B.n526 585
R1303 B.n173 B.n172 585
R1304 B.n178 B.n173 585
R1305 B.n535 B.n534 585
R1306 B.n534 B.n533 585
R1307 B.n536 B.n171 585
R1308 B.n171 B.n170 585
R1309 B.n538 B.n537 585
R1310 B.n539 B.n538 585
R1311 B.n165 B.n164 585
R1312 B.n166 B.n165 585
R1313 B.n547 B.n546 585
R1314 B.n546 B.n545 585
R1315 B.n548 B.n163 585
R1316 B.n163 B.n161 585
R1317 B.n550 B.n549 585
R1318 B.n551 B.n550 585
R1319 B.n157 B.n156 585
R1320 B.n162 B.n157 585
R1321 B.n559 B.n558 585
R1322 B.n558 B.n557 585
R1323 B.n560 B.n155 585
R1324 B.n155 B.n154 585
R1325 B.n562 B.n561 585
R1326 B.n563 B.n562 585
R1327 B.n149 B.n148 585
R1328 B.n150 B.n149 585
R1329 B.n571 B.n570 585
R1330 B.n570 B.n569 585
R1331 B.n572 B.n147 585
R1332 B.n147 B.n145 585
R1333 B.n574 B.n573 585
R1334 B.n575 B.n574 585
R1335 B.n141 B.n140 585
R1336 B.n146 B.n141 585
R1337 B.n584 B.n583 585
R1338 B.n583 B.n582 585
R1339 B.n585 B.n139 585
R1340 B.n139 B.n138 585
R1341 B.n587 B.n586 585
R1342 B.n588 B.n587 585
R1343 B.n3 B.n0 585
R1344 B.n4 B.n3 585
R1345 B.n921 B.n1 585
R1346 B.n922 B.n921 585
R1347 B.n920 B.n919 585
R1348 B.n920 B.n8 585
R1349 B.n918 B.n9 585
R1350 B.n12 B.n9 585
R1351 B.n917 B.n916 585
R1352 B.n916 B.n915 585
R1353 B.n11 B.n10 585
R1354 B.n914 B.n11 585
R1355 B.n912 B.n911 585
R1356 B.n913 B.n912 585
R1357 B.n910 B.n17 585
R1358 B.n17 B.n16 585
R1359 B.n909 B.n908 585
R1360 B.n908 B.n907 585
R1361 B.n19 B.n18 585
R1362 B.n906 B.n19 585
R1363 B.n904 B.n903 585
R1364 B.n905 B.n904 585
R1365 B.n902 B.n24 585
R1366 B.n24 B.n23 585
R1367 B.n901 B.n900 585
R1368 B.n900 B.n899 585
R1369 B.n26 B.n25 585
R1370 B.n898 B.n26 585
R1371 B.n896 B.n895 585
R1372 B.n897 B.n896 585
R1373 B.n894 B.n31 585
R1374 B.n31 B.n30 585
R1375 B.n893 B.n892 585
R1376 B.n892 B.n891 585
R1377 B.n33 B.n32 585
R1378 B.n890 B.n33 585
R1379 B.n888 B.n887 585
R1380 B.n889 B.n888 585
R1381 B.n886 B.n38 585
R1382 B.n38 B.n37 585
R1383 B.n885 B.n884 585
R1384 B.n884 B.n883 585
R1385 B.n40 B.n39 585
R1386 B.n882 B.n40 585
R1387 B.n880 B.n879 585
R1388 B.n881 B.n880 585
R1389 B.n878 B.n45 585
R1390 B.n45 B.n44 585
R1391 B.n877 B.n876 585
R1392 B.n876 B.n875 585
R1393 B.n47 B.n46 585
R1394 B.n874 B.n47 585
R1395 B.n872 B.n871 585
R1396 B.n873 B.n872 585
R1397 B.n870 B.n52 585
R1398 B.n52 B.n51 585
R1399 B.n869 B.n868 585
R1400 B.n868 B.n867 585
R1401 B.n54 B.n53 585
R1402 B.n866 B.n54 585
R1403 B.n864 B.n863 585
R1404 B.n865 B.n864 585
R1405 B.n862 B.n59 585
R1406 B.n59 B.n58 585
R1407 B.n861 B.n860 585
R1408 B.n860 B.n859 585
R1409 B.n61 B.n60 585
R1410 B.n858 B.n61 585
R1411 B.n856 B.n855 585
R1412 B.n857 B.n856 585
R1413 B.n854 B.n66 585
R1414 B.n66 B.n65 585
R1415 B.n853 B.n852 585
R1416 B.n852 B.n851 585
R1417 B.n68 B.n67 585
R1418 B.n850 B.n68 585
R1419 B.n848 B.n847 585
R1420 B.n849 B.n848 585
R1421 B.n846 B.n72 585
R1422 B.n75 B.n72 585
R1423 B.n845 B.n844 585
R1424 B.n844 B.n843 585
R1425 B.n74 B.n73 585
R1426 B.n842 B.n74 585
R1427 B.n840 B.n839 585
R1428 B.n841 B.n840 585
R1429 B.n838 B.n80 585
R1430 B.n80 B.n79 585
R1431 B.n837 B.n836 585
R1432 B.n836 B.n835 585
R1433 B.n82 B.n81 585
R1434 B.n834 B.n82 585
R1435 B.n832 B.n831 585
R1436 B.n833 B.n832 585
R1437 B.n925 B.n924 585
R1438 B.n923 B.n2 585
R1439 B.n832 B.n87 540.549
R1440 B.n135 B.n85 540.549
R1441 B.n455 B.n224 540.549
R1442 B.n453 B.n226 540.549
R1443 B.n108 B.t8 327.394
R1444 B.n114 B.t12 327.394
R1445 B.n253 B.t15 327.394
R1446 B.n247 B.t19 327.394
R1447 B.n114 B.t13 322.466
R1448 B.n253 B.t18 322.466
R1449 B.n108 B.t10 322.466
R1450 B.n247 B.t21 322.466
R1451 B.n115 B.t14 271.654
R1452 B.n254 B.t17 271.654
R1453 B.n109 B.t11 271.654
R1454 B.n248 B.t20 271.654
R1455 B.n655 B.n86 256.663
R1456 B.n657 B.n86 256.663
R1457 B.n663 B.n86 256.663
R1458 B.n665 B.n86 256.663
R1459 B.n671 B.n86 256.663
R1460 B.n673 B.n86 256.663
R1461 B.n679 B.n86 256.663
R1462 B.n681 B.n86 256.663
R1463 B.n687 B.n86 256.663
R1464 B.n689 B.n86 256.663
R1465 B.n695 B.n86 256.663
R1466 B.n697 B.n86 256.663
R1467 B.n703 B.n86 256.663
R1468 B.n705 B.n86 256.663
R1469 B.n711 B.n86 256.663
R1470 B.n713 B.n86 256.663
R1471 B.n719 B.n86 256.663
R1472 B.n721 B.n86 256.663
R1473 B.n727 B.n86 256.663
R1474 B.n729 B.n86 256.663
R1475 B.n736 B.n86 256.663
R1476 B.n738 B.n86 256.663
R1477 B.n744 B.n86 256.663
R1478 B.n746 B.n86 256.663
R1479 B.n753 B.n86 256.663
R1480 B.n755 B.n86 256.663
R1481 B.n761 B.n86 256.663
R1482 B.n763 B.n86 256.663
R1483 B.n769 B.n86 256.663
R1484 B.n771 B.n86 256.663
R1485 B.n777 B.n86 256.663
R1486 B.n779 B.n86 256.663
R1487 B.n785 B.n86 256.663
R1488 B.n787 B.n86 256.663
R1489 B.n793 B.n86 256.663
R1490 B.n795 B.n86 256.663
R1491 B.n801 B.n86 256.663
R1492 B.n803 B.n86 256.663
R1493 B.n809 B.n86 256.663
R1494 B.n811 B.n86 256.663
R1495 B.n817 B.n86 256.663
R1496 B.n819 B.n86 256.663
R1497 B.n825 B.n86 256.663
R1498 B.n827 B.n86 256.663
R1499 B.n448 B.n225 256.663
R1500 B.n228 B.n225 256.663
R1501 B.n441 B.n225 256.663
R1502 B.n435 B.n225 256.663
R1503 B.n433 B.n225 256.663
R1504 B.n427 B.n225 256.663
R1505 B.n425 B.n225 256.663
R1506 B.n419 B.n225 256.663
R1507 B.n417 B.n225 256.663
R1508 B.n411 B.n225 256.663
R1509 B.n409 B.n225 256.663
R1510 B.n403 B.n225 256.663
R1511 B.n401 B.n225 256.663
R1512 B.n395 B.n225 256.663
R1513 B.n393 B.n225 256.663
R1514 B.n387 B.n225 256.663
R1515 B.n385 B.n225 256.663
R1516 B.n379 B.n225 256.663
R1517 B.n377 B.n225 256.663
R1518 B.n370 B.n225 256.663
R1519 B.n368 B.n225 256.663
R1520 B.n362 B.n225 256.663
R1521 B.n360 B.n225 256.663
R1522 B.n354 B.n225 256.663
R1523 B.n256 B.n225 256.663
R1524 B.n348 B.n225 256.663
R1525 B.n342 B.n225 256.663
R1526 B.n340 B.n225 256.663
R1527 B.n334 B.n225 256.663
R1528 B.n332 B.n225 256.663
R1529 B.n326 B.n225 256.663
R1530 B.n324 B.n225 256.663
R1531 B.n318 B.n225 256.663
R1532 B.n316 B.n225 256.663
R1533 B.n310 B.n225 256.663
R1534 B.n308 B.n225 256.663
R1535 B.n302 B.n225 256.663
R1536 B.n300 B.n225 256.663
R1537 B.n294 B.n225 256.663
R1538 B.n292 B.n225 256.663
R1539 B.n286 B.n225 256.663
R1540 B.n284 B.n225 256.663
R1541 B.n278 B.n225 256.663
R1542 B.n276 B.n225 256.663
R1543 B.n927 B.n926 256.663
R1544 B.n828 B.n826 163.367
R1545 B.n824 B.n89 163.367
R1546 B.n820 B.n818 163.367
R1547 B.n816 B.n91 163.367
R1548 B.n812 B.n810 163.367
R1549 B.n808 B.n93 163.367
R1550 B.n804 B.n802 163.367
R1551 B.n800 B.n95 163.367
R1552 B.n796 B.n794 163.367
R1553 B.n792 B.n97 163.367
R1554 B.n788 B.n786 163.367
R1555 B.n784 B.n99 163.367
R1556 B.n780 B.n778 163.367
R1557 B.n776 B.n101 163.367
R1558 B.n772 B.n770 163.367
R1559 B.n768 B.n103 163.367
R1560 B.n764 B.n762 163.367
R1561 B.n760 B.n105 163.367
R1562 B.n756 B.n754 163.367
R1563 B.n752 B.n107 163.367
R1564 B.n747 B.n745 163.367
R1565 B.n743 B.n111 163.367
R1566 B.n739 B.n737 163.367
R1567 B.n735 B.n113 163.367
R1568 B.n730 B.n728 163.367
R1569 B.n726 B.n117 163.367
R1570 B.n722 B.n720 163.367
R1571 B.n718 B.n119 163.367
R1572 B.n714 B.n712 163.367
R1573 B.n710 B.n121 163.367
R1574 B.n706 B.n704 163.367
R1575 B.n702 B.n123 163.367
R1576 B.n698 B.n696 163.367
R1577 B.n694 B.n125 163.367
R1578 B.n690 B.n688 163.367
R1579 B.n686 B.n127 163.367
R1580 B.n682 B.n680 163.367
R1581 B.n678 B.n129 163.367
R1582 B.n674 B.n672 163.367
R1583 B.n670 B.n131 163.367
R1584 B.n666 B.n664 163.367
R1585 B.n662 B.n133 163.367
R1586 B.n658 B.n656 163.367
R1587 B.n654 B.n135 163.367
R1588 B.n455 B.n222 163.367
R1589 B.n459 B.n222 163.367
R1590 B.n459 B.n216 163.367
R1591 B.n467 B.n216 163.367
R1592 B.n467 B.n214 163.367
R1593 B.n471 B.n214 163.367
R1594 B.n471 B.n209 163.367
R1595 B.n480 B.n209 163.367
R1596 B.n480 B.n207 163.367
R1597 B.n484 B.n207 163.367
R1598 B.n484 B.n201 163.367
R1599 B.n492 B.n201 163.367
R1600 B.n492 B.n199 163.367
R1601 B.n496 B.n199 163.367
R1602 B.n496 B.n192 163.367
R1603 B.n504 B.n192 163.367
R1604 B.n504 B.n190 163.367
R1605 B.n508 B.n190 163.367
R1606 B.n508 B.n185 163.367
R1607 B.n516 B.n185 163.367
R1608 B.n516 B.n183 163.367
R1609 B.n520 B.n183 163.367
R1610 B.n520 B.n176 163.367
R1611 B.n528 B.n176 163.367
R1612 B.n528 B.n174 163.367
R1613 B.n532 B.n174 163.367
R1614 B.n532 B.n169 163.367
R1615 B.n540 B.n169 163.367
R1616 B.n540 B.n167 163.367
R1617 B.n544 B.n167 163.367
R1618 B.n544 B.n160 163.367
R1619 B.n552 B.n160 163.367
R1620 B.n552 B.n158 163.367
R1621 B.n556 B.n158 163.367
R1622 B.n556 B.n153 163.367
R1623 B.n564 B.n153 163.367
R1624 B.n564 B.n151 163.367
R1625 B.n568 B.n151 163.367
R1626 B.n568 B.n144 163.367
R1627 B.n576 B.n144 163.367
R1628 B.n576 B.n142 163.367
R1629 B.n581 B.n142 163.367
R1630 B.n581 B.n137 163.367
R1631 B.n589 B.n137 163.367
R1632 B.n590 B.n589 163.367
R1633 B.n590 B.n5 163.367
R1634 B.n6 B.n5 163.367
R1635 B.n7 B.n6 163.367
R1636 B.n596 B.n7 163.367
R1637 B.n597 B.n596 163.367
R1638 B.n597 B.n13 163.367
R1639 B.n14 B.n13 163.367
R1640 B.n15 B.n14 163.367
R1641 B.n602 B.n15 163.367
R1642 B.n602 B.n20 163.367
R1643 B.n21 B.n20 163.367
R1644 B.n22 B.n21 163.367
R1645 B.n607 B.n22 163.367
R1646 B.n607 B.n27 163.367
R1647 B.n28 B.n27 163.367
R1648 B.n29 B.n28 163.367
R1649 B.n612 B.n29 163.367
R1650 B.n612 B.n34 163.367
R1651 B.n35 B.n34 163.367
R1652 B.n36 B.n35 163.367
R1653 B.n617 B.n36 163.367
R1654 B.n617 B.n41 163.367
R1655 B.n42 B.n41 163.367
R1656 B.n43 B.n42 163.367
R1657 B.n622 B.n43 163.367
R1658 B.n622 B.n48 163.367
R1659 B.n49 B.n48 163.367
R1660 B.n50 B.n49 163.367
R1661 B.n627 B.n50 163.367
R1662 B.n627 B.n55 163.367
R1663 B.n56 B.n55 163.367
R1664 B.n57 B.n56 163.367
R1665 B.n632 B.n57 163.367
R1666 B.n632 B.n62 163.367
R1667 B.n63 B.n62 163.367
R1668 B.n64 B.n63 163.367
R1669 B.n637 B.n64 163.367
R1670 B.n637 B.n69 163.367
R1671 B.n70 B.n69 163.367
R1672 B.n71 B.n70 163.367
R1673 B.n642 B.n71 163.367
R1674 B.n642 B.n76 163.367
R1675 B.n77 B.n76 163.367
R1676 B.n78 B.n77 163.367
R1677 B.n647 B.n78 163.367
R1678 B.n647 B.n83 163.367
R1679 B.n84 B.n83 163.367
R1680 B.n85 B.n84 163.367
R1681 B.n449 B.n447 163.367
R1682 B.n447 B.n446 163.367
R1683 B.n443 B.n442 163.367
R1684 B.n440 B.n230 163.367
R1685 B.n436 B.n434 163.367
R1686 B.n432 B.n232 163.367
R1687 B.n428 B.n426 163.367
R1688 B.n424 B.n234 163.367
R1689 B.n420 B.n418 163.367
R1690 B.n416 B.n236 163.367
R1691 B.n412 B.n410 163.367
R1692 B.n408 B.n238 163.367
R1693 B.n404 B.n402 163.367
R1694 B.n400 B.n240 163.367
R1695 B.n396 B.n394 163.367
R1696 B.n392 B.n242 163.367
R1697 B.n388 B.n386 163.367
R1698 B.n384 B.n244 163.367
R1699 B.n380 B.n378 163.367
R1700 B.n376 B.n246 163.367
R1701 B.n371 B.n369 163.367
R1702 B.n367 B.n250 163.367
R1703 B.n363 B.n361 163.367
R1704 B.n359 B.n252 163.367
R1705 B.n355 B.n353 163.367
R1706 B.n350 B.n349 163.367
R1707 B.n347 B.n258 163.367
R1708 B.n343 B.n341 163.367
R1709 B.n339 B.n260 163.367
R1710 B.n335 B.n333 163.367
R1711 B.n331 B.n262 163.367
R1712 B.n327 B.n325 163.367
R1713 B.n323 B.n264 163.367
R1714 B.n319 B.n317 163.367
R1715 B.n315 B.n266 163.367
R1716 B.n311 B.n309 163.367
R1717 B.n307 B.n268 163.367
R1718 B.n303 B.n301 163.367
R1719 B.n299 B.n270 163.367
R1720 B.n295 B.n293 163.367
R1721 B.n291 B.n272 163.367
R1722 B.n287 B.n285 163.367
R1723 B.n283 B.n274 163.367
R1724 B.n279 B.n277 163.367
R1725 B.n453 B.n220 163.367
R1726 B.n461 B.n220 163.367
R1727 B.n461 B.n218 163.367
R1728 B.n465 B.n218 163.367
R1729 B.n465 B.n212 163.367
R1730 B.n474 B.n212 163.367
R1731 B.n474 B.n210 163.367
R1732 B.n478 B.n210 163.367
R1733 B.n478 B.n205 163.367
R1734 B.n486 B.n205 163.367
R1735 B.n486 B.n203 163.367
R1736 B.n490 B.n203 163.367
R1737 B.n490 B.n197 163.367
R1738 B.n498 B.n197 163.367
R1739 B.n498 B.n195 163.367
R1740 B.n502 B.n195 163.367
R1741 B.n502 B.n189 163.367
R1742 B.n510 B.n189 163.367
R1743 B.n510 B.n187 163.367
R1744 B.n514 B.n187 163.367
R1745 B.n514 B.n181 163.367
R1746 B.n522 B.n181 163.367
R1747 B.n522 B.n179 163.367
R1748 B.n526 B.n179 163.367
R1749 B.n526 B.n173 163.367
R1750 B.n534 B.n173 163.367
R1751 B.n534 B.n171 163.367
R1752 B.n538 B.n171 163.367
R1753 B.n538 B.n165 163.367
R1754 B.n546 B.n165 163.367
R1755 B.n546 B.n163 163.367
R1756 B.n550 B.n163 163.367
R1757 B.n550 B.n157 163.367
R1758 B.n558 B.n157 163.367
R1759 B.n558 B.n155 163.367
R1760 B.n562 B.n155 163.367
R1761 B.n562 B.n149 163.367
R1762 B.n570 B.n149 163.367
R1763 B.n570 B.n147 163.367
R1764 B.n574 B.n147 163.367
R1765 B.n574 B.n141 163.367
R1766 B.n583 B.n141 163.367
R1767 B.n583 B.n139 163.367
R1768 B.n587 B.n139 163.367
R1769 B.n587 B.n3 163.367
R1770 B.n925 B.n3 163.367
R1771 B.n921 B.n2 163.367
R1772 B.n921 B.n920 163.367
R1773 B.n920 B.n9 163.367
R1774 B.n916 B.n9 163.367
R1775 B.n916 B.n11 163.367
R1776 B.n912 B.n11 163.367
R1777 B.n912 B.n17 163.367
R1778 B.n908 B.n17 163.367
R1779 B.n908 B.n19 163.367
R1780 B.n904 B.n19 163.367
R1781 B.n904 B.n24 163.367
R1782 B.n900 B.n24 163.367
R1783 B.n900 B.n26 163.367
R1784 B.n896 B.n26 163.367
R1785 B.n896 B.n31 163.367
R1786 B.n892 B.n31 163.367
R1787 B.n892 B.n33 163.367
R1788 B.n888 B.n33 163.367
R1789 B.n888 B.n38 163.367
R1790 B.n884 B.n38 163.367
R1791 B.n884 B.n40 163.367
R1792 B.n880 B.n40 163.367
R1793 B.n880 B.n45 163.367
R1794 B.n876 B.n45 163.367
R1795 B.n876 B.n47 163.367
R1796 B.n872 B.n47 163.367
R1797 B.n872 B.n52 163.367
R1798 B.n868 B.n52 163.367
R1799 B.n868 B.n54 163.367
R1800 B.n864 B.n54 163.367
R1801 B.n864 B.n59 163.367
R1802 B.n860 B.n59 163.367
R1803 B.n860 B.n61 163.367
R1804 B.n856 B.n61 163.367
R1805 B.n856 B.n66 163.367
R1806 B.n852 B.n66 163.367
R1807 B.n852 B.n68 163.367
R1808 B.n848 B.n68 163.367
R1809 B.n848 B.n72 163.367
R1810 B.n844 B.n72 163.367
R1811 B.n844 B.n74 163.367
R1812 B.n840 B.n74 163.367
R1813 B.n840 B.n80 163.367
R1814 B.n836 B.n80 163.367
R1815 B.n836 B.n82 163.367
R1816 B.n832 B.n82 163.367
R1817 B.n454 B.n225 87.7893
R1818 B.n833 B.n86 87.7893
R1819 B.n827 B.n87 71.676
R1820 B.n826 B.n825 71.676
R1821 B.n819 B.n89 71.676
R1822 B.n818 B.n817 71.676
R1823 B.n811 B.n91 71.676
R1824 B.n810 B.n809 71.676
R1825 B.n803 B.n93 71.676
R1826 B.n802 B.n801 71.676
R1827 B.n795 B.n95 71.676
R1828 B.n794 B.n793 71.676
R1829 B.n787 B.n97 71.676
R1830 B.n786 B.n785 71.676
R1831 B.n779 B.n99 71.676
R1832 B.n778 B.n777 71.676
R1833 B.n771 B.n101 71.676
R1834 B.n770 B.n769 71.676
R1835 B.n763 B.n103 71.676
R1836 B.n762 B.n761 71.676
R1837 B.n755 B.n105 71.676
R1838 B.n754 B.n753 71.676
R1839 B.n746 B.n107 71.676
R1840 B.n745 B.n744 71.676
R1841 B.n738 B.n111 71.676
R1842 B.n737 B.n736 71.676
R1843 B.n729 B.n113 71.676
R1844 B.n728 B.n727 71.676
R1845 B.n721 B.n117 71.676
R1846 B.n720 B.n719 71.676
R1847 B.n713 B.n119 71.676
R1848 B.n712 B.n711 71.676
R1849 B.n705 B.n121 71.676
R1850 B.n704 B.n703 71.676
R1851 B.n697 B.n123 71.676
R1852 B.n696 B.n695 71.676
R1853 B.n689 B.n125 71.676
R1854 B.n688 B.n687 71.676
R1855 B.n681 B.n127 71.676
R1856 B.n680 B.n679 71.676
R1857 B.n673 B.n129 71.676
R1858 B.n672 B.n671 71.676
R1859 B.n665 B.n131 71.676
R1860 B.n664 B.n663 71.676
R1861 B.n657 B.n133 71.676
R1862 B.n656 B.n655 71.676
R1863 B.n655 B.n654 71.676
R1864 B.n658 B.n657 71.676
R1865 B.n663 B.n662 71.676
R1866 B.n666 B.n665 71.676
R1867 B.n671 B.n670 71.676
R1868 B.n674 B.n673 71.676
R1869 B.n679 B.n678 71.676
R1870 B.n682 B.n681 71.676
R1871 B.n687 B.n686 71.676
R1872 B.n690 B.n689 71.676
R1873 B.n695 B.n694 71.676
R1874 B.n698 B.n697 71.676
R1875 B.n703 B.n702 71.676
R1876 B.n706 B.n705 71.676
R1877 B.n711 B.n710 71.676
R1878 B.n714 B.n713 71.676
R1879 B.n719 B.n718 71.676
R1880 B.n722 B.n721 71.676
R1881 B.n727 B.n726 71.676
R1882 B.n730 B.n729 71.676
R1883 B.n736 B.n735 71.676
R1884 B.n739 B.n738 71.676
R1885 B.n744 B.n743 71.676
R1886 B.n747 B.n746 71.676
R1887 B.n753 B.n752 71.676
R1888 B.n756 B.n755 71.676
R1889 B.n761 B.n760 71.676
R1890 B.n764 B.n763 71.676
R1891 B.n769 B.n768 71.676
R1892 B.n772 B.n771 71.676
R1893 B.n777 B.n776 71.676
R1894 B.n780 B.n779 71.676
R1895 B.n785 B.n784 71.676
R1896 B.n788 B.n787 71.676
R1897 B.n793 B.n792 71.676
R1898 B.n796 B.n795 71.676
R1899 B.n801 B.n800 71.676
R1900 B.n804 B.n803 71.676
R1901 B.n809 B.n808 71.676
R1902 B.n812 B.n811 71.676
R1903 B.n817 B.n816 71.676
R1904 B.n820 B.n819 71.676
R1905 B.n825 B.n824 71.676
R1906 B.n828 B.n827 71.676
R1907 B.n448 B.n226 71.676
R1908 B.n446 B.n228 71.676
R1909 B.n442 B.n441 71.676
R1910 B.n435 B.n230 71.676
R1911 B.n434 B.n433 71.676
R1912 B.n427 B.n232 71.676
R1913 B.n426 B.n425 71.676
R1914 B.n419 B.n234 71.676
R1915 B.n418 B.n417 71.676
R1916 B.n411 B.n236 71.676
R1917 B.n410 B.n409 71.676
R1918 B.n403 B.n238 71.676
R1919 B.n402 B.n401 71.676
R1920 B.n395 B.n240 71.676
R1921 B.n394 B.n393 71.676
R1922 B.n387 B.n242 71.676
R1923 B.n386 B.n385 71.676
R1924 B.n379 B.n244 71.676
R1925 B.n378 B.n377 71.676
R1926 B.n370 B.n246 71.676
R1927 B.n369 B.n368 71.676
R1928 B.n362 B.n250 71.676
R1929 B.n361 B.n360 71.676
R1930 B.n354 B.n252 71.676
R1931 B.n353 B.n256 71.676
R1932 B.n349 B.n348 71.676
R1933 B.n342 B.n258 71.676
R1934 B.n341 B.n340 71.676
R1935 B.n334 B.n260 71.676
R1936 B.n333 B.n332 71.676
R1937 B.n326 B.n262 71.676
R1938 B.n325 B.n324 71.676
R1939 B.n318 B.n264 71.676
R1940 B.n317 B.n316 71.676
R1941 B.n310 B.n266 71.676
R1942 B.n309 B.n308 71.676
R1943 B.n302 B.n268 71.676
R1944 B.n301 B.n300 71.676
R1945 B.n294 B.n270 71.676
R1946 B.n293 B.n292 71.676
R1947 B.n286 B.n272 71.676
R1948 B.n285 B.n284 71.676
R1949 B.n278 B.n274 71.676
R1950 B.n277 B.n276 71.676
R1951 B.n449 B.n448 71.676
R1952 B.n443 B.n228 71.676
R1953 B.n441 B.n440 71.676
R1954 B.n436 B.n435 71.676
R1955 B.n433 B.n432 71.676
R1956 B.n428 B.n427 71.676
R1957 B.n425 B.n424 71.676
R1958 B.n420 B.n419 71.676
R1959 B.n417 B.n416 71.676
R1960 B.n412 B.n411 71.676
R1961 B.n409 B.n408 71.676
R1962 B.n404 B.n403 71.676
R1963 B.n401 B.n400 71.676
R1964 B.n396 B.n395 71.676
R1965 B.n393 B.n392 71.676
R1966 B.n388 B.n387 71.676
R1967 B.n385 B.n384 71.676
R1968 B.n380 B.n379 71.676
R1969 B.n377 B.n376 71.676
R1970 B.n371 B.n370 71.676
R1971 B.n368 B.n367 71.676
R1972 B.n363 B.n362 71.676
R1973 B.n360 B.n359 71.676
R1974 B.n355 B.n354 71.676
R1975 B.n350 B.n256 71.676
R1976 B.n348 B.n347 71.676
R1977 B.n343 B.n342 71.676
R1978 B.n340 B.n339 71.676
R1979 B.n335 B.n334 71.676
R1980 B.n332 B.n331 71.676
R1981 B.n327 B.n326 71.676
R1982 B.n324 B.n323 71.676
R1983 B.n319 B.n318 71.676
R1984 B.n316 B.n315 71.676
R1985 B.n311 B.n310 71.676
R1986 B.n308 B.n307 71.676
R1987 B.n303 B.n302 71.676
R1988 B.n300 B.n299 71.676
R1989 B.n295 B.n294 71.676
R1990 B.n292 B.n291 71.676
R1991 B.n287 B.n286 71.676
R1992 B.n284 B.n283 71.676
R1993 B.n279 B.n278 71.676
R1994 B.n276 B.n224 71.676
R1995 B.n926 B.n925 71.676
R1996 B.n926 B.n2 71.676
R1997 B.n750 B.n109 59.5399
R1998 B.n732 B.n115 59.5399
R1999 B.n255 B.n254 59.5399
R2000 B.n373 B.n248 59.5399
R2001 B.n109 B.n108 50.8126
R2002 B.n115 B.n114 50.8126
R2003 B.n254 B.n253 50.8126
R2004 B.n248 B.n247 50.8126
R2005 B.n454 B.n221 44.885
R2006 B.n460 B.n221 44.885
R2007 B.n460 B.n217 44.885
R2008 B.n466 B.n217 44.885
R2009 B.n466 B.n213 44.885
R2010 B.n473 B.n213 44.885
R2011 B.n473 B.n472 44.885
R2012 B.n479 B.n206 44.885
R2013 B.n485 B.n206 44.885
R2014 B.n485 B.n202 44.885
R2015 B.n491 B.n202 44.885
R2016 B.n491 B.n198 44.885
R2017 B.n497 B.n198 44.885
R2018 B.n497 B.n193 44.885
R2019 B.n503 B.n193 44.885
R2020 B.n503 B.n194 44.885
R2021 B.n509 B.n186 44.885
R2022 B.n515 B.n186 44.885
R2023 B.n515 B.n182 44.885
R2024 B.n521 B.n182 44.885
R2025 B.n521 B.n177 44.885
R2026 B.n527 B.n177 44.885
R2027 B.n527 B.n178 44.885
R2028 B.n533 B.n170 44.885
R2029 B.n539 B.n170 44.885
R2030 B.n539 B.n166 44.885
R2031 B.n545 B.n166 44.885
R2032 B.n545 B.n161 44.885
R2033 B.n551 B.n161 44.885
R2034 B.n551 B.n162 44.885
R2035 B.n557 B.n154 44.885
R2036 B.n563 B.n154 44.885
R2037 B.n563 B.n150 44.885
R2038 B.n569 B.n150 44.885
R2039 B.n569 B.n145 44.885
R2040 B.n575 B.n145 44.885
R2041 B.n575 B.n146 44.885
R2042 B.n582 B.n138 44.885
R2043 B.n588 B.n138 44.885
R2044 B.n588 B.n4 44.885
R2045 B.n924 B.n4 44.885
R2046 B.n924 B.n923 44.885
R2047 B.n923 B.n922 44.885
R2048 B.n922 B.n8 44.885
R2049 B.n12 B.n8 44.885
R2050 B.n915 B.n12 44.885
R2051 B.n914 B.n913 44.885
R2052 B.n913 B.n16 44.885
R2053 B.n907 B.n16 44.885
R2054 B.n907 B.n906 44.885
R2055 B.n906 B.n905 44.885
R2056 B.n905 B.n23 44.885
R2057 B.n899 B.n23 44.885
R2058 B.n898 B.n897 44.885
R2059 B.n897 B.n30 44.885
R2060 B.n891 B.n30 44.885
R2061 B.n891 B.n890 44.885
R2062 B.n890 B.n889 44.885
R2063 B.n889 B.n37 44.885
R2064 B.n883 B.n37 44.885
R2065 B.n882 B.n881 44.885
R2066 B.n881 B.n44 44.885
R2067 B.n875 B.n44 44.885
R2068 B.n875 B.n874 44.885
R2069 B.n874 B.n873 44.885
R2070 B.n873 B.n51 44.885
R2071 B.n867 B.n51 44.885
R2072 B.n866 B.n865 44.885
R2073 B.n865 B.n58 44.885
R2074 B.n859 B.n58 44.885
R2075 B.n859 B.n858 44.885
R2076 B.n858 B.n857 44.885
R2077 B.n857 B.n65 44.885
R2078 B.n851 B.n65 44.885
R2079 B.n851 B.n850 44.885
R2080 B.n850 B.n849 44.885
R2081 B.n843 B.n75 44.885
R2082 B.n843 B.n842 44.885
R2083 B.n842 B.n841 44.885
R2084 B.n841 B.n79 44.885
R2085 B.n835 B.n79 44.885
R2086 B.n835 B.n834 44.885
R2087 B.n834 B.n833 44.885
R2088 B.n479 B.t16 44.2249
R2089 B.n849 B.t9 44.2249
R2090 B.n582 B.t2 42.9048
R2091 B.n915 B.t0 42.9048
R2092 B.n194 B.t7 41.5847
R2093 B.t1 B.n866 41.5847
R2094 B.n452 B.n451 35.1225
R2095 B.n456 B.n223 35.1225
R2096 B.n652 B.n651 35.1225
R2097 B.n831 B.n830 35.1225
R2098 B.n557 B.t6 29.7035
R2099 B.n899 B.t4 29.7035
R2100 B.n178 B.t5 28.3833
R2101 B.t3 B.n882 28.3833
R2102 B B.n927 18.0485
R2103 B.n533 B.t5 16.5021
R2104 B.n883 B.t3 16.5021
R2105 B.n162 B.t6 15.182
R2106 B.t4 B.n898 15.182
R2107 B.n452 B.n219 10.6151
R2108 B.n462 B.n219 10.6151
R2109 B.n463 B.n462 10.6151
R2110 B.n464 B.n463 10.6151
R2111 B.n464 B.n211 10.6151
R2112 B.n475 B.n211 10.6151
R2113 B.n476 B.n475 10.6151
R2114 B.n477 B.n476 10.6151
R2115 B.n477 B.n204 10.6151
R2116 B.n487 B.n204 10.6151
R2117 B.n488 B.n487 10.6151
R2118 B.n489 B.n488 10.6151
R2119 B.n489 B.n196 10.6151
R2120 B.n499 B.n196 10.6151
R2121 B.n500 B.n499 10.6151
R2122 B.n501 B.n500 10.6151
R2123 B.n501 B.n188 10.6151
R2124 B.n511 B.n188 10.6151
R2125 B.n512 B.n511 10.6151
R2126 B.n513 B.n512 10.6151
R2127 B.n513 B.n180 10.6151
R2128 B.n523 B.n180 10.6151
R2129 B.n524 B.n523 10.6151
R2130 B.n525 B.n524 10.6151
R2131 B.n525 B.n172 10.6151
R2132 B.n535 B.n172 10.6151
R2133 B.n536 B.n535 10.6151
R2134 B.n537 B.n536 10.6151
R2135 B.n537 B.n164 10.6151
R2136 B.n547 B.n164 10.6151
R2137 B.n548 B.n547 10.6151
R2138 B.n549 B.n548 10.6151
R2139 B.n549 B.n156 10.6151
R2140 B.n559 B.n156 10.6151
R2141 B.n560 B.n559 10.6151
R2142 B.n561 B.n560 10.6151
R2143 B.n561 B.n148 10.6151
R2144 B.n571 B.n148 10.6151
R2145 B.n572 B.n571 10.6151
R2146 B.n573 B.n572 10.6151
R2147 B.n573 B.n140 10.6151
R2148 B.n584 B.n140 10.6151
R2149 B.n585 B.n584 10.6151
R2150 B.n586 B.n585 10.6151
R2151 B.n586 B.n0 10.6151
R2152 B.n451 B.n450 10.6151
R2153 B.n450 B.n227 10.6151
R2154 B.n445 B.n227 10.6151
R2155 B.n445 B.n444 10.6151
R2156 B.n444 B.n229 10.6151
R2157 B.n439 B.n229 10.6151
R2158 B.n439 B.n438 10.6151
R2159 B.n438 B.n437 10.6151
R2160 B.n437 B.n231 10.6151
R2161 B.n431 B.n231 10.6151
R2162 B.n431 B.n430 10.6151
R2163 B.n430 B.n429 10.6151
R2164 B.n429 B.n233 10.6151
R2165 B.n423 B.n233 10.6151
R2166 B.n423 B.n422 10.6151
R2167 B.n422 B.n421 10.6151
R2168 B.n421 B.n235 10.6151
R2169 B.n415 B.n235 10.6151
R2170 B.n415 B.n414 10.6151
R2171 B.n414 B.n413 10.6151
R2172 B.n413 B.n237 10.6151
R2173 B.n407 B.n237 10.6151
R2174 B.n407 B.n406 10.6151
R2175 B.n406 B.n405 10.6151
R2176 B.n405 B.n239 10.6151
R2177 B.n399 B.n239 10.6151
R2178 B.n399 B.n398 10.6151
R2179 B.n398 B.n397 10.6151
R2180 B.n397 B.n241 10.6151
R2181 B.n391 B.n241 10.6151
R2182 B.n391 B.n390 10.6151
R2183 B.n390 B.n389 10.6151
R2184 B.n389 B.n243 10.6151
R2185 B.n383 B.n243 10.6151
R2186 B.n383 B.n382 10.6151
R2187 B.n382 B.n381 10.6151
R2188 B.n381 B.n245 10.6151
R2189 B.n375 B.n245 10.6151
R2190 B.n375 B.n374 10.6151
R2191 B.n372 B.n249 10.6151
R2192 B.n366 B.n249 10.6151
R2193 B.n366 B.n365 10.6151
R2194 B.n365 B.n364 10.6151
R2195 B.n364 B.n251 10.6151
R2196 B.n358 B.n251 10.6151
R2197 B.n358 B.n357 10.6151
R2198 B.n357 B.n356 10.6151
R2199 B.n352 B.n351 10.6151
R2200 B.n351 B.n257 10.6151
R2201 B.n346 B.n257 10.6151
R2202 B.n346 B.n345 10.6151
R2203 B.n345 B.n344 10.6151
R2204 B.n344 B.n259 10.6151
R2205 B.n338 B.n259 10.6151
R2206 B.n338 B.n337 10.6151
R2207 B.n337 B.n336 10.6151
R2208 B.n336 B.n261 10.6151
R2209 B.n330 B.n261 10.6151
R2210 B.n330 B.n329 10.6151
R2211 B.n329 B.n328 10.6151
R2212 B.n328 B.n263 10.6151
R2213 B.n322 B.n263 10.6151
R2214 B.n322 B.n321 10.6151
R2215 B.n321 B.n320 10.6151
R2216 B.n320 B.n265 10.6151
R2217 B.n314 B.n265 10.6151
R2218 B.n314 B.n313 10.6151
R2219 B.n313 B.n312 10.6151
R2220 B.n312 B.n267 10.6151
R2221 B.n306 B.n267 10.6151
R2222 B.n306 B.n305 10.6151
R2223 B.n305 B.n304 10.6151
R2224 B.n304 B.n269 10.6151
R2225 B.n298 B.n269 10.6151
R2226 B.n298 B.n297 10.6151
R2227 B.n297 B.n296 10.6151
R2228 B.n296 B.n271 10.6151
R2229 B.n290 B.n271 10.6151
R2230 B.n290 B.n289 10.6151
R2231 B.n289 B.n288 10.6151
R2232 B.n288 B.n273 10.6151
R2233 B.n282 B.n273 10.6151
R2234 B.n282 B.n281 10.6151
R2235 B.n281 B.n280 10.6151
R2236 B.n280 B.n275 10.6151
R2237 B.n275 B.n223 10.6151
R2238 B.n457 B.n456 10.6151
R2239 B.n458 B.n457 10.6151
R2240 B.n458 B.n215 10.6151
R2241 B.n468 B.n215 10.6151
R2242 B.n469 B.n468 10.6151
R2243 B.n470 B.n469 10.6151
R2244 B.n470 B.n208 10.6151
R2245 B.n481 B.n208 10.6151
R2246 B.n482 B.n481 10.6151
R2247 B.n483 B.n482 10.6151
R2248 B.n483 B.n200 10.6151
R2249 B.n493 B.n200 10.6151
R2250 B.n494 B.n493 10.6151
R2251 B.n495 B.n494 10.6151
R2252 B.n495 B.n191 10.6151
R2253 B.n505 B.n191 10.6151
R2254 B.n506 B.n505 10.6151
R2255 B.n507 B.n506 10.6151
R2256 B.n507 B.n184 10.6151
R2257 B.n517 B.n184 10.6151
R2258 B.n518 B.n517 10.6151
R2259 B.n519 B.n518 10.6151
R2260 B.n519 B.n175 10.6151
R2261 B.n529 B.n175 10.6151
R2262 B.n530 B.n529 10.6151
R2263 B.n531 B.n530 10.6151
R2264 B.n531 B.n168 10.6151
R2265 B.n541 B.n168 10.6151
R2266 B.n542 B.n541 10.6151
R2267 B.n543 B.n542 10.6151
R2268 B.n543 B.n159 10.6151
R2269 B.n553 B.n159 10.6151
R2270 B.n554 B.n553 10.6151
R2271 B.n555 B.n554 10.6151
R2272 B.n555 B.n152 10.6151
R2273 B.n565 B.n152 10.6151
R2274 B.n566 B.n565 10.6151
R2275 B.n567 B.n566 10.6151
R2276 B.n567 B.n143 10.6151
R2277 B.n577 B.n143 10.6151
R2278 B.n578 B.n577 10.6151
R2279 B.n580 B.n578 10.6151
R2280 B.n580 B.n579 10.6151
R2281 B.n579 B.n136 10.6151
R2282 B.n591 B.n136 10.6151
R2283 B.n592 B.n591 10.6151
R2284 B.n593 B.n592 10.6151
R2285 B.n594 B.n593 10.6151
R2286 B.n595 B.n594 10.6151
R2287 B.n598 B.n595 10.6151
R2288 B.n599 B.n598 10.6151
R2289 B.n600 B.n599 10.6151
R2290 B.n601 B.n600 10.6151
R2291 B.n603 B.n601 10.6151
R2292 B.n604 B.n603 10.6151
R2293 B.n605 B.n604 10.6151
R2294 B.n606 B.n605 10.6151
R2295 B.n608 B.n606 10.6151
R2296 B.n609 B.n608 10.6151
R2297 B.n610 B.n609 10.6151
R2298 B.n611 B.n610 10.6151
R2299 B.n613 B.n611 10.6151
R2300 B.n614 B.n613 10.6151
R2301 B.n615 B.n614 10.6151
R2302 B.n616 B.n615 10.6151
R2303 B.n618 B.n616 10.6151
R2304 B.n619 B.n618 10.6151
R2305 B.n620 B.n619 10.6151
R2306 B.n621 B.n620 10.6151
R2307 B.n623 B.n621 10.6151
R2308 B.n624 B.n623 10.6151
R2309 B.n625 B.n624 10.6151
R2310 B.n626 B.n625 10.6151
R2311 B.n628 B.n626 10.6151
R2312 B.n629 B.n628 10.6151
R2313 B.n630 B.n629 10.6151
R2314 B.n631 B.n630 10.6151
R2315 B.n633 B.n631 10.6151
R2316 B.n634 B.n633 10.6151
R2317 B.n635 B.n634 10.6151
R2318 B.n636 B.n635 10.6151
R2319 B.n638 B.n636 10.6151
R2320 B.n639 B.n638 10.6151
R2321 B.n640 B.n639 10.6151
R2322 B.n641 B.n640 10.6151
R2323 B.n643 B.n641 10.6151
R2324 B.n644 B.n643 10.6151
R2325 B.n645 B.n644 10.6151
R2326 B.n646 B.n645 10.6151
R2327 B.n648 B.n646 10.6151
R2328 B.n649 B.n648 10.6151
R2329 B.n650 B.n649 10.6151
R2330 B.n651 B.n650 10.6151
R2331 B.n919 B.n1 10.6151
R2332 B.n919 B.n918 10.6151
R2333 B.n918 B.n917 10.6151
R2334 B.n917 B.n10 10.6151
R2335 B.n911 B.n10 10.6151
R2336 B.n911 B.n910 10.6151
R2337 B.n910 B.n909 10.6151
R2338 B.n909 B.n18 10.6151
R2339 B.n903 B.n18 10.6151
R2340 B.n903 B.n902 10.6151
R2341 B.n902 B.n901 10.6151
R2342 B.n901 B.n25 10.6151
R2343 B.n895 B.n25 10.6151
R2344 B.n895 B.n894 10.6151
R2345 B.n894 B.n893 10.6151
R2346 B.n893 B.n32 10.6151
R2347 B.n887 B.n32 10.6151
R2348 B.n887 B.n886 10.6151
R2349 B.n886 B.n885 10.6151
R2350 B.n885 B.n39 10.6151
R2351 B.n879 B.n39 10.6151
R2352 B.n879 B.n878 10.6151
R2353 B.n878 B.n877 10.6151
R2354 B.n877 B.n46 10.6151
R2355 B.n871 B.n46 10.6151
R2356 B.n871 B.n870 10.6151
R2357 B.n870 B.n869 10.6151
R2358 B.n869 B.n53 10.6151
R2359 B.n863 B.n53 10.6151
R2360 B.n863 B.n862 10.6151
R2361 B.n862 B.n861 10.6151
R2362 B.n861 B.n60 10.6151
R2363 B.n855 B.n60 10.6151
R2364 B.n855 B.n854 10.6151
R2365 B.n854 B.n853 10.6151
R2366 B.n853 B.n67 10.6151
R2367 B.n847 B.n67 10.6151
R2368 B.n847 B.n846 10.6151
R2369 B.n846 B.n845 10.6151
R2370 B.n845 B.n73 10.6151
R2371 B.n839 B.n73 10.6151
R2372 B.n839 B.n838 10.6151
R2373 B.n838 B.n837 10.6151
R2374 B.n837 B.n81 10.6151
R2375 B.n831 B.n81 10.6151
R2376 B.n830 B.n829 10.6151
R2377 B.n829 B.n88 10.6151
R2378 B.n823 B.n88 10.6151
R2379 B.n823 B.n822 10.6151
R2380 B.n822 B.n821 10.6151
R2381 B.n821 B.n90 10.6151
R2382 B.n815 B.n90 10.6151
R2383 B.n815 B.n814 10.6151
R2384 B.n814 B.n813 10.6151
R2385 B.n813 B.n92 10.6151
R2386 B.n807 B.n92 10.6151
R2387 B.n807 B.n806 10.6151
R2388 B.n806 B.n805 10.6151
R2389 B.n805 B.n94 10.6151
R2390 B.n799 B.n94 10.6151
R2391 B.n799 B.n798 10.6151
R2392 B.n798 B.n797 10.6151
R2393 B.n797 B.n96 10.6151
R2394 B.n791 B.n96 10.6151
R2395 B.n791 B.n790 10.6151
R2396 B.n790 B.n789 10.6151
R2397 B.n789 B.n98 10.6151
R2398 B.n783 B.n98 10.6151
R2399 B.n783 B.n782 10.6151
R2400 B.n782 B.n781 10.6151
R2401 B.n781 B.n100 10.6151
R2402 B.n775 B.n100 10.6151
R2403 B.n775 B.n774 10.6151
R2404 B.n774 B.n773 10.6151
R2405 B.n773 B.n102 10.6151
R2406 B.n767 B.n102 10.6151
R2407 B.n767 B.n766 10.6151
R2408 B.n766 B.n765 10.6151
R2409 B.n765 B.n104 10.6151
R2410 B.n759 B.n104 10.6151
R2411 B.n759 B.n758 10.6151
R2412 B.n758 B.n757 10.6151
R2413 B.n757 B.n106 10.6151
R2414 B.n751 B.n106 10.6151
R2415 B.n749 B.n748 10.6151
R2416 B.n748 B.n110 10.6151
R2417 B.n742 B.n110 10.6151
R2418 B.n742 B.n741 10.6151
R2419 B.n741 B.n740 10.6151
R2420 B.n740 B.n112 10.6151
R2421 B.n734 B.n112 10.6151
R2422 B.n734 B.n733 10.6151
R2423 B.n731 B.n116 10.6151
R2424 B.n725 B.n116 10.6151
R2425 B.n725 B.n724 10.6151
R2426 B.n724 B.n723 10.6151
R2427 B.n723 B.n118 10.6151
R2428 B.n717 B.n118 10.6151
R2429 B.n717 B.n716 10.6151
R2430 B.n716 B.n715 10.6151
R2431 B.n715 B.n120 10.6151
R2432 B.n709 B.n120 10.6151
R2433 B.n709 B.n708 10.6151
R2434 B.n708 B.n707 10.6151
R2435 B.n707 B.n122 10.6151
R2436 B.n701 B.n122 10.6151
R2437 B.n701 B.n700 10.6151
R2438 B.n700 B.n699 10.6151
R2439 B.n699 B.n124 10.6151
R2440 B.n693 B.n124 10.6151
R2441 B.n693 B.n692 10.6151
R2442 B.n692 B.n691 10.6151
R2443 B.n691 B.n126 10.6151
R2444 B.n685 B.n126 10.6151
R2445 B.n685 B.n684 10.6151
R2446 B.n684 B.n683 10.6151
R2447 B.n683 B.n128 10.6151
R2448 B.n677 B.n128 10.6151
R2449 B.n677 B.n676 10.6151
R2450 B.n676 B.n675 10.6151
R2451 B.n675 B.n130 10.6151
R2452 B.n669 B.n130 10.6151
R2453 B.n669 B.n668 10.6151
R2454 B.n668 B.n667 10.6151
R2455 B.n667 B.n132 10.6151
R2456 B.n661 B.n132 10.6151
R2457 B.n661 B.n660 10.6151
R2458 B.n660 B.n659 10.6151
R2459 B.n659 B.n134 10.6151
R2460 B.n653 B.n134 10.6151
R2461 B.n653 B.n652 10.6151
R2462 B.n927 B.n0 8.11757
R2463 B.n927 B.n1 8.11757
R2464 B.n373 B.n372 6.5566
R2465 B.n356 B.n255 6.5566
R2466 B.n750 B.n749 6.5566
R2467 B.n733 B.n732 6.5566
R2468 B.n374 B.n373 4.05904
R2469 B.n352 B.n255 4.05904
R2470 B.n751 B.n750 4.05904
R2471 B.n732 B.n731 4.05904
R2472 B.n509 B.t7 3.30083
R2473 B.n867 B.t1 3.30083
R2474 B.n146 B.t2 1.9807
R2475 B.t0 B.n914 1.9807
R2476 B.n472 B.t16 0.660566
R2477 B.n75 B.t9 0.660566
R2478 VN.n51 VN.n27 161.3
R2479 VN.n50 VN.n49 161.3
R2480 VN.n48 VN.n28 161.3
R2481 VN.n47 VN.n46 161.3
R2482 VN.n45 VN.n29 161.3
R2483 VN.n43 VN.n42 161.3
R2484 VN.n41 VN.n30 161.3
R2485 VN.n40 VN.n39 161.3
R2486 VN.n38 VN.n31 161.3
R2487 VN.n37 VN.n36 161.3
R2488 VN.n35 VN.n32 161.3
R2489 VN.n24 VN.n0 161.3
R2490 VN.n23 VN.n22 161.3
R2491 VN.n21 VN.n1 161.3
R2492 VN.n20 VN.n19 161.3
R2493 VN.n18 VN.n2 161.3
R2494 VN.n16 VN.n15 161.3
R2495 VN.n14 VN.n3 161.3
R2496 VN.n13 VN.n12 161.3
R2497 VN.n11 VN.n4 161.3
R2498 VN.n10 VN.n9 161.3
R2499 VN.n8 VN.n5 161.3
R2500 VN.n7 VN.t5 150.291
R2501 VN.n34 VN.t6 150.291
R2502 VN.n6 VN.t4 119.87
R2503 VN.n17 VN.t2 119.87
R2504 VN.n25 VN.t7 119.87
R2505 VN.n33 VN.t3 119.87
R2506 VN.n44 VN.t1 119.87
R2507 VN.n52 VN.t0 119.87
R2508 VN.n26 VN.n25 101.948
R2509 VN.n53 VN.n52 101.948
R2510 VN.n7 VN.n6 69.279
R2511 VN.n34 VN.n33 69.279
R2512 VN.n12 VN.n11 56.5193
R2513 VN.n39 VN.n38 56.5193
R2514 VN.n19 VN.n1 53.1199
R2515 VN.n46 VN.n28 53.1199
R2516 VN VN.n53 49.1875
R2517 VN.n23 VN.n1 27.8669
R2518 VN.n50 VN.n28 27.8669
R2519 VN.n10 VN.n5 24.4675
R2520 VN.n11 VN.n10 24.4675
R2521 VN.n12 VN.n3 24.4675
R2522 VN.n16 VN.n3 24.4675
R2523 VN.n19 VN.n18 24.4675
R2524 VN.n24 VN.n23 24.4675
R2525 VN.n38 VN.n37 24.4675
R2526 VN.n37 VN.n32 24.4675
R2527 VN.n46 VN.n45 24.4675
R2528 VN.n43 VN.n30 24.4675
R2529 VN.n39 VN.n30 24.4675
R2530 VN.n51 VN.n50 24.4675
R2531 VN.n18 VN.n17 21.5315
R2532 VN.n45 VN.n44 21.5315
R2533 VN.n35 VN.n34 10.1472
R2534 VN.n8 VN.n7 10.1472
R2535 VN.n25 VN.n24 8.80862
R2536 VN.n52 VN.n51 8.80862
R2537 VN.n6 VN.n5 2.93654
R2538 VN.n17 VN.n16 2.93654
R2539 VN.n33 VN.n32 2.93654
R2540 VN.n44 VN.n43 2.93654
R2541 VN.n53 VN.n27 0.278367
R2542 VN.n26 VN.n0 0.278367
R2543 VN.n49 VN.n27 0.189894
R2544 VN.n49 VN.n48 0.189894
R2545 VN.n48 VN.n47 0.189894
R2546 VN.n47 VN.n29 0.189894
R2547 VN.n42 VN.n29 0.189894
R2548 VN.n42 VN.n41 0.189894
R2549 VN.n41 VN.n40 0.189894
R2550 VN.n40 VN.n31 0.189894
R2551 VN.n36 VN.n31 0.189894
R2552 VN.n36 VN.n35 0.189894
R2553 VN.n9 VN.n8 0.189894
R2554 VN.n9 VN.n4 0.189894
R2555 VN.n13 VN.n4 0.189894
R2556 VN.n14 VN.n13 0.189894
R2557 VN.n15 VN.n14 0.189894
R2558 VN.n15 VN.n2 0.189894
R2559 VN.n20 VN.n2 0.189894
R2560 VN.n21 VN.n20 0.189894
R2561 VN.n22 VN.n21 0.189894
R2562 VN.n22 VN.n0 0.189894
R2563 VN VN.n26 0.153454
R2564 VDD2.n2 VDD2.n1 62.9698
R2565 VDD2.n2 VDD2.n0 62.9698
R2566 VDD2 VDD2.n5 62.9669
R2567 VDD2.n4 VDD2.n3 61.896
R2568 VDD2.n4 VDD2.n2 43.6981
R2569 VDD2.n5 VDD2.t4 1.73887
R2570 VDD2.n5 VDD2.t1 1.73887
R2571 VDD2.n3 VDD2.t7 1.73887
R2572 VDD2.n3 VDD2.t6 1.73887
R2573 VDD2.n1 VDD2.t5 1.73887
R2574 VDD2.n1 VDD2.t0 1.73887
R2575 VDD2.n0 VDD2.t2 1.73887
R2576 VDD2.n0 VDD2.t3 1.73887
R2577 VDD2 VDD2.n4 1.188
C0 VP VN 7.17499f
C1 VN VDD1 0.151121f
C2 VP VTAIL 8.3908f
C3 VTAIL VDD1 7.83276f
C4 VP VDD1 8.39125f
C5 VN VDD2 8.05698f
C6 VTAIL VDD2 7.8851f
C7 VP VDD2 0.486637f
C8 VDD1 VDD2 1.61574f
C9 VN VTAIL 8.376691f
C10 VDD2 B 5.004424f
C11 VDD1 B 5.405201f
C12 VTAIL B 9.910336f
C13 VN B 14.28618f
C14 VP B 12.841186f
C15 VDD2.t2 B 0.220417f
C16 VDD2.t3 B 0.220417f
C17 VDD2.n0 B 1.96553f
C18 VDD2.t5 B 0.220417f
C19 VDD2.t0 B 0.220417f
C20 VDD2.n1 B 1.96553f
C21 VDD2.n2 B 2.99863f
C22 VDD2.t7 B 0.220417f
C23 VDD2.t6 B 0.220417f
C24 VDD2.n3 B 1.95743f
C25 VDD2.n4 B 2.73909f
C26 VDD2.t4 B 0.220417f
C27 VDD2.t1 B 0.220417f
C28 VDD2.n5 B 1.9655f
C29 VN.n0 B 0.031942f
C30 VN.t7 B 1.71914f
C31 VN.n1 B 0.025411f
C32 VN.n2 B 0.024228f
C33 VN.t2 B 1.71914f
C34 VN.n3 B 0.045154f
C35 VN.n4 B 0.024228f
C36 VN.n5 B 0.025536f
C37 VN.t5 B 1.86938f
C38 VN.t4 B 1.71914f
C39 VN.n6 B 0.669689f
C40 VN.n7 B 0.671667f
C41 VN.n8 B 0.207917f
C42 VN.n9 B 0.024228f
C43 VN.n10 B 0.045154f
C44 VN.n11 B 0.035368f
C45 VN.n12 B 0.035368f
C46 VN.n13 B 0.024228f
C47 VN.n14 B 0.024228f
C48 VN.n15 B 0.024228f
C49 VN.n16 B 0.025536f
C50 VN.n17 B 0.612615f
C51 VN.n18 B 0.042479f
C52 VN.n19 B 0.042988f
C53 VN.n20 B 0.024228f
C54 VN.n21 B 0.024228f
C55 VN.n22 B 0.024228f
C56 VN.n23 B 0.047492f
C57 VN.n24 B 0.030887f
C58 VN.n25 B 0.682141f
C59 VN.n26 B 0.03769f
C60 VN.n27 B 0.031942f
C61 VN.t0 B 1.71914f
C62 VN.n28 B 0.025411f
C63 VN.n29 B 0.024228f
C64 VN.t1 B 1.71914f
C65 VN.n30 B 0.045154f
C66 VN.n31 B 0.024228f
C67 VN.n32 B 0.025536f
C68 VN.t6 B 1.86938f
C69 VN.t3 B 1.71914f
C70 VN.n33 B 0.669689f
C71 VN.n34 B 0.671667f
C72 VN.n35 B 0.207917f
C73 VN.n36 B 0.024228f
C74 VN.n37 B 0.045154f
C75 VN.n38 B 0.035368f
C76 VN.n39 B 0.035368f
C77 VN.n40 B 0.024228f
C78 VN.n41 B 0.024228f
C79 VN.n42 B 0.024228f
C80 VN.n43 B 0.025536f
C81 VN.n44 B 0.612615f
C82 VN.n45 B 0.042479f
C83 VN.n46 B 0.042988f
C84 VN.n47 B 0.024228f
C85 VN.n48 B 0.024228f
C86 VN.n49 B 0.024228f
C87 VN.n50 B 0.047492f
C88 VN.n51 B 0.030887f
C89 VN.n52 B 0.682141f
C90 VN.n53 B 1.31494f
C91 VTAIL.t4 B 0.178061f
C92 VTAIL.t3 B 0.178061f
C93 VTAIL.n0 B 1.52241f
C94 VTAIL.n1 B 0.343f
C95 VTAIL.n2 B 0.027139f
C96 VTAIL.n3 B 0.019783f
C97 VTAIL.n4 B 0.010631f
C98 VTAIL.n5 B 0.025127f
C99 VTAIL.n6 B 0.011256f
C100 VTAIL.n7 B 0.019783f
C101 VTAIL.n8 B 0.010631f
C102 VTAIL.n9 B 0.025127f
C103 VTAIL.n10 B 0.010943f
C104 VTAIL.n11 B 0.019783f
C105 VTAIL.n12 B 0.011256f
C106 VTAIL.n13 B 0.025127f
C107 VTAIL.n14 B 0.011256f
C108 VTAIL.n15 B 0.019783f
C109 VTAIL.n16 B 0.010631f
C110 VTAIL.n17 B 0.025127f
C111 VTAIL.n18 B 0.011256f
C112 VTAIL.n19 B 0.944339f
C113 VTAIL.n20 B 0.010631f
C114 VTAIL.t0 B 0.042372f
C115 VTAIL.n21 B 0.138f
C116 VTAIL.n22 B 0.017763f
C117 VTAIL.n23 B 0.018845f
C118 VTAIL.n24 B 0.025127f
C119 VTAIL.n25 B 0.011256f
C120 VTAIL.n26 B 0.010631f
C121 VTAIL.n27 B 0.019783f
C122 VTAIL.n28 B 0.019783f
C123 VTAIL.n29 B 0.010631f
C124 VTAIL.n30 B 0.011256f
C125 VTAIL.n31 B 0.025127f
C126 VTAIL.n32 B 0.025127f
C127 VTAIL.n33 B 0.011256f
C128 VTAIL.n34 B 0.010631f
C129 VTAIL.n35 B 0.019783f
C130 VTAIL.n36 B 0.019783f
C131 VTAIL.n37 B 0.010631f
C132 VTAIL.n38 B 0.010631f
C133 VTAIL.n39 B 0.011256f
C134 VTAIL.n40 B 0.025127f
C135 VTAIL.n41 B 0.025127f
C136 VTAIL.n42 B 0.025127f
C137 VTAIL.n43 B 0.010943f
C138 VTAIL.n44 B 0.010631f
C139 VTAIL.n45 B 0.019783f
C140 VTAIL.n46 B 0.019783f
C141 VTAIL.n47 B 0.010631f
C142 VTAIL.n48 B 0.011256f
C143 VTAIL.n49 B 0.025127f
C144 VTAIL.n50 B 0.025127f
C145 VTAIL.n51 B 0.011256f
C146 VTAIL.n52 B 0.010631f
C147 VTAIL.n53 B 0.019783f
C148 VTAIL.n54 B 0.019783f
C149 VTAIL.n55 B 0.010631f
C150 VTAIL.n56 B 0.011256f
C151 VTAIL.n57 B 0.025127f
C152 VTAIL.n58 B 0.053215f
C153 VTAIL.n59 B 0.011256f
C154 VTAIL.n60 B 0.010631f
C155 VTAIL.n61 B 0.045457f
C156 VTAIL.n62 B 0.029646f
C157 VTAIL.n63 B 0.190669f
C158 VTAIL.n64 B 0.027139f
C159 VTAIL.n65 B 0.019783f
C160 VTAIL.n66 B 0.010631f
C161 VTAIL.n67 B 0.025127f
C162 VTAIL.n68 B 0.011256f
C163 VTAIL.n69 B 0.019783f
C164 VTAIL.n70 B 0.010631f
C165 VTAIL.n71 B 0.025127f
C166 VTAIL.n72 B 0.010943f
C167 VTAIL.n73 B 0.019783f
C168 VTAIL.n74 B 0.011256f
C169 VTAIL.n75 B 0.025127f
C170 VTAIL.n76 B 0.011256f
C171 VTAIL.n77 B 0.019783f
C172 VTAIL.n78 B 0.010631f
C173 VTAIL.n79 B 0.025127f
C174 VTAIL.n80 B 0.011256f
C175 VTAIL.n81 B 0.944339f
C176 VTAIL.n82 B 0.010631f
C177 VTAIL.t12 B 0.042372f
C178 VTAIL.n83 B 0.138f
C179 VTAIL.n84 B 0.017763f
C180 VTAIL.n85 B 0.018845f
C181 VTAIL.n86 B 0.025127f
C182 VTAIL.n87 B 0.011256f
C183 VTAIL.n88 B 0.010631f
C184 VTAIL.n89 B 0.019783f
C185 VTAIL.n90 B 0.019783f
C186 VTAIL.n91 B 0.010631f
C187 VTAIL.n92 B 0.011256f
C188 VTAIL.n93 B 0.025127f
C189 VTAIL.n94 B 0.025127f
C190 VTAIL.n95 B 0.011256f
C191 VTAIL.n96 B 0.010631f
C192 VTAIL.n97 B 0.019783f
C193 VTAIL.n98 B 0.019783f
C194 VTAIL.n99 B 0.010631f
C195 VTAIL.n100 B 0.010631f
C196 VTAIL.n101 B 0.011256f
C197 VTAIL.n102 B 0.025127f
C198 VTAIL.n103 B 0.025127f
C199 VTAIL.n104 B 0.025127f
C200 VTAIL.n105 B 0.010943f
C201 VTAIL.n106 B 0.010631f
C202 VTAIL.n107 B 0.019783f
C203 VTAIL.n108 B 0.019783f
C204 VTAIL.n109 B 0.010631f
C205 VTAIL.n110 B 0.011256f
C206 VTAIL.n111 B 0.025127f
C207 VTAIL.n112 B 0.025127f
C208 VTAIL.n113 B 0.011256f
C209 VTAIL.n114 B 0.010631f
C210 VTAIL.n115 B 0.019783f
C211 VTAIL.n116 B 0.019783f
C212 VTAIL.n117 B 0.010631f
C213 VTAIL.n118 B 0.011256f
C214 VTAIL.n119 B 0.025127f
C215 VTAIL.n120 B 0.053215f
C216 VTAIL.n121 B 0.011256f
C217 VTAIL.n122 B 0.010631f
C218 VTAIL.n123 B 0.045457f
C219 VTAIL.n124 B 0.029646f
C220 VTAIL.n125 B 0.190669f
C221 VTAIL.t10 B 0.178061f
C222 VTAIL.t6 B 0.178061f
C223 VTAIL.n126 B 1.52241f
C224 VTAIL.n127 B 0.483266f
C225 VTAIL.n128 B 0.027139f
C226 VTAIL.n129 B 0.019783f
C227 VTAIL.n130 B 0.010631f
C228 VTAIL.n131 B 0.025127f
C229 VTAIL.n132 B 0.011256f
C230 VTAIL.n133 B 0.019783f
C231 VTAIL.n134 B 0.010631f
C232 VTAIL.n135 B 0.025127f
C233 VTAIL.n136 B 0.010943f
C234 VTAIL.n137 B 0.019783f
C235 VTAIL.n138 B 0.011256f
C236 VTAIL.n139 B 0.025127f
C237 VTAIL.n140 B 0.011256f
C238 VTAIL.n141 B 0.019783f
C239 VTAIL.n142 B 0.010631f
C240 VTAIL.n143 B 0.025127f
C241 VTAIL.n144 B 0.011256f
C242 VTAIL.n145 B 0.944339f
C243 VTAIL.n146 B 0.010631f
C244 VTAIL.t7 B 0.042372f
C245 VTAIL.n147 B 0.138f
C246 VTAIL.n148 B 0.017763f
C247 VTAIL.n149 B 0.018845f
C248 VTAIL.n150 B 0.025127f
C249 VTAIL.n151 B 0.011256f
C250 VTAIL.n152 B 0.010631f
C251 VTAIL.n153 B 0.019783f
C252 VTAIL.n154 B 0.019783f
C253 VTAIL.n155 B 0.010631f
C254 VTAIL.n156 B 0.011256f
C255 VTAIL.n157 B 0.025127f
C256 VTAIL.n158 B 0.025127f
C257 VTAIL.n159 B 0.011256f
C258 VTAIL.n160 B 0.010631f
C259 VTAIL.n161 B 0.019783f
C260 VTAIL.n162 B 0.019783f
C261 VTAIL.n163 B 0.010631f
C262 VTAIL.n164 B 0.010631f
C263 VTAIL.n165 B 0.011256f
C264 VTAIL.n166 B 0.025127f
C265 VTAIL.n167 B 0.025127f
C266 VTAIL.n168 B 0.025127f
C267 VTAIL.n169 B 0.010943f
C268 VTAIL.n170 B 0.010631f
C269 VTAIL.n171 B 0.019783f
C270 VTAIL.n172 B 0.019783f
C271 VTAIL.n173 B 0.010631f
C272 VTAIL.n174 B 0.011256f
C273 VTAIL.n175 B 0.025127f
C274 VTAIL.n176 B 0.025127f
C275 VTAIL.n177 B 0.011256f
C276 VTAIL.n178 B 0.010631f
C277 VTAIL.n179 B 0.019783f
C278 VTAIL.n180 B 0.019783f
C279 VTAIL.n181 B 0.010631f
C280 VTAIL.n182 B 0.011256f
C281 VTAIL.n183 B 0.025127f
C282 VTAIL.n184 B 0.053215f
C283 VTAIL.n185 B 0.011256f
C284 VTAIL.n186 B 0.010631f
C285 VTAIL.n187 B 0.045457f
C286 VTAIL.n188 B 0.029646f
C287 VTAIL.n189 B 1.19933f
C288 VTAIL.n190 B 0.027139f
C289 VTAIL.n191 B 0.019783f
C290 VTAIL.n192 B 0.010631f
C291 VTAIL.n193 B 0.025127f
C292 VTAIL.n194 B 0.011256f
C293 VTAIL.n195 B 0.019783f
C294 VTAIL.n196 B 0.010631f
C295 VTAIL.n197 B 0.025127f
C296 VTAIL.n198 B 0.010943f
C297 VTAIL.n199 B 0.019783f
C298 VTAIL.n200 B 0.010943f
C299 VTAIL.n201 B 0.010631f
C300 VTAIL.n202 B 0.025127f
C301 VTAIL.n203 B 0.025127f
C302 VTAIL.n204 B 0.011256f
C303 VTAIL.n205 B 0.019783f
C304 VTAIL.n206 B 0.010631f
C305 VTAIL.n207 B 0.025127f
C306 VTAIL.n208 B 0.011256f
C307 VTAIL.n209 B 0.944339f
C308 VTAIL.n210 B 0.010631f
C309 VTAIL.t15 B 0.042372f
C310 VTAIL.n211 B 0.138f
C311 VTAIL.n212 B 0.017763f
C312 VTAIL.n213 B 0.018845f
C313 VTAIL.n214 B 0.025127f
C314 VTAIL.n215 B 0.011256f
C315 VTAIL.n216 B 0.010631f
C316 VTAIL.n217 B 0.019783f
C317 VTAIL.n218 B 0.019783f
C318 VTAIL.n219 B 0.010631f
C319 VTAIL.n220 B 0.011256f
C320 VTAIL.n221 B 0.025127f
C321 VTAIL.n222 B 0.025127f
C322 VTAIL.n223 B 0.011256f
C323 VTAIL.n224 B 0.010631f
C324 VTAIL.n225 B 0.019783f
C325 VTAIL.n226 B 0.019783f
C326 VTAIL.n227 B 0.010631f
C327 VTAIL.n228 B 0.011256f
C328 VTAIL.n229 B 0.025127f
C329 VTAIL.n230 B 0.025127f
C330 VTAIL.n231 B 0.011256f
C331 VTAIL.n232 B 0.010631f
C332 VTAIL.n233 B 0.019783f
C333 VTAIL.n234 B 0.019783f
C334 VTAIL.n235 B 0.010631f
C335 VTAIL.n236 B 0.011256f
C336 VTAIL.n237 B 0.025127f
C337 VTAIL.n238 B 0.025127f
C338 VTAIL.n239 B 0.011256f
C339 VTAIL.n240 B 0.010631f
C340 VTAIL.n241 B 0.019783f
C341 VTAIL.n242 B 0.019783f
C342 VTAIL.n243 B 0.010631f
C343 VTAIL.n244 B 0.011256f
C344 VTAIL.n245 B 0.025127f
C345 VTAIL.n246 B 0.053215f
C346 VTAIL.n247 B 0.011256f
C347 VTAIL.n248 B 0.010631f
C348 VTAIL.n249 B 0.045457f
C349 VTAIL.n250 B 0.029646f
C350 VTAIL.n251 B 1.19933f
C351 VTAIL.t5 B 0.178061f
C352 VTAIL.t14 B 0.178061f
C353 VTAIL.n252 B 1.52242f
C354 VTAIL.n253 B 0.483257f
C355 VTAIL.n254 B 0.027139f
C356 VTAIL.n255 B 0.019783f
C357 VTAIL.n256 B 0.010631f
C358 VTAIL.n257 B 0.025127f
C359 VTAIL.n258 B 0.011256f
C360 VTAIL.n259 B 0.019783f
C361 VTAIL.n260 B 0.010631f
C362 VTAIL.n261 B 0.025127f
C363 VTAIL.n262 B 0.010943f
C364 VTAIL.n263 B 0.019783f
C365 VTAIL.n264 B 0.010943f
C366 VTAIL.n265 B 0.010631f
C367 VTAIL.n266 B 0.025127f
C368 VTAIL.n267 B 0.025127f
C369 VTAIL.n268 B 0.011256f
C370 VTAIL.n269 B 0.019783f
C371 VTAIL.n270 B 0.010631f
C372 VTAIL.n271 B 0.025127f
C373 VTAIL.n272 B 0.011256f
C374 VTAIL.n273 B 0.944339f
C375 VTAIL.n274 B 0.010631f
C376 VTAIL.t2 B 0.042372f
C377 VTAIL.n275 B 0.138f
C378 VTAIL.n276 B 0.017763f
C379 VTAIL.n277 B 0.018845f
C380 VTAIL.n278 B 0.025127f
C381 VTAIL.n279 B 0.011256f
C382 VTAIL.n280 B 0.010631f
C383 VTAIL.n281 B 0.019783f
C384 VTAIL.n282 B 0.019783f
C385 VTAIL.n283 B 0.010631f
C386 VTAIL.n284 B 0.011256f
C387 VTAIL.n285 B 0.025127f
C388 VTAIL.n286 B 0.025127f
C389 VTAIL.n287 B 0.011256f
C390 VTAIL.n288 B 0.010631f
C391 VTAIL.n289 B 0.019783f
C392 VTAIL.n290 B 0.019783f
C393 VTAIL.n291 B 0.010631f
C394 VTAIL.n292 B 0.011256f
C395 VTAIL.n293 B 0.025127f
C396 VTAIL.n294 B 0.025127f
C397 VTAIL.n295 B 0.011256f
C398 VTAIL.n296 B 0.010631f
C399 VTAIL.n297 B 0.019783f
C400 VTAIL.n298 B 0.019783f
C401 VTAIL.n299 B 0.010631f
C402 VTAIL.n300 B 0.011256f
C403 VTAIL.n301 B 0.025127f
C404 VTAIL.n302 B 0.025127f
C405 VTAIL.n303 B 0.011256f
C406 VTAIL.n304 B 0.010631f
C407 VTAIL.n305 B 0.019783f
C408 VTAIL.n306 B 0.019783f
C409 VTAIL.n307 B 0.010631f
C410 VTAIL.n308 B 0.011256f
C411 VTAIL.n309 B 0.025127f
C412 VTAIL.n310 B 0.053215f
C413 VTAIL.n311 B 0.011256f
C414 VTAIL.n312 B 0.010631f
C415 VTAIL.n313 B 0.045457f
C416 VTAIL.n314 B 0.029646f
C417 VTAIL.n315 B 0.190669f
C418 VTAIL.n316 B 0.027139f
C419 VTAIL.n317 B 0.019783f
C420 VTAIL.n318 B 0.010631f
C421 VTAIL.n319 B 0.025127f
C422 VTAIL.n320 B 0.011256f
C423 VTAIL.n321 B 0.019783f
C424 VTAIL.n322 B 0.010631f
C425 VTAIL.n323 B 0.025127f
C426 VTAIL.n324 B 0.010943f
C427 VTAIL.n325 B 0.019783f
C428 VTAIL.n326 B 0.010943f
C429 VTAIL.n327 B 0.010631f
C430 VTAIL.n328 B 0.025127f
C431 VTAIL.n329 B 0.025127f
C432 VTAIL.n330 B 0.011256f
C433 VTAIL.n331 B 0.019783f
C434 VTAIL.n332 B 0.010631f
C435 VTAIL.n333 B 0.025127f
C436 VTAIL.n334 B 0.011256f
C437 VTAIL.n335 B 0.944339f
C438 VTAIL.n336 B 0.010631f
C439 VTAIL.t8 B 0.042372f
C440 VTAIL.n337 B 0.138f
C441 VTAIL.n338 B 0.017763f
C442 VTAIL.n339 B 0.018845f
C443 VTAIL.n340 B 0.025127f
C444 VTAIL.n341 B 0.011256f
C445 VTAIL.n342 B 0.010631f
C446 VTAIL.n343 B 0.019783f
C447 VTAIL.n344 B 0.019783f
C448 VTAIL.n345 B 0.010631f
C449 VTAIL.n346 B 0.011256f
C450 VTAIL.n347 B 0.025127f
C451 VTAIL.n348 B 0.025127f
C452 VTAIL.n349 B 0.011256f
C453 VTAIL.n350 B 0.010631f
C454 VTAIL.n351 B 0.019783f
C455 VTAIL.n352 B 0.019783f
C456 VTAIL.n353 B 0.010631f
C457 VTAIL.n354 B 0.011256f
C458 VTAIL.n355 B 0.025127f
C459 VTAIL.n356 B 0.025127f
C460 VTAIL.n357 B 0.011256f
C461 VTAIL.n358 B 0.010631f
C462 VTAIL.n359 B 0.019783f
C463 VTAIL.n360 B 0.019783f
C464 VTAIL.n361 B 0.010631f
C465 VTAIL.n362 B 0.011256f
C466 VTAIL.n363 B 0.025127f
C467 VTAIL.n364 B 0.025127f
C468 VTAIL.n365 B 0.011256f
C469 VTAIL.n366 B 0.010631f
C470 VTAIL.n367 B 0.019783f
C471 VTAIL.n368 B 0.019783f
C472 VTAIL.n369 B 0.010631f
C473 VTAIL.n370 B 0.011256f
C474 VTAIL.n371 B 0.025127f
C475 VTAIL.n372 B 0.053215f
C476 VTAIL.n373 B 0.011256f
C477 VTAIL.n374 B 0.010631f
C478 VTAIL.n375 B 0.045457f
C479 VTAIL.n376 B 0.029646f
C480 VTAIL.n377 B 0.190669f
C481 VTAIL.t11 B 0.178061f
C482 VTAIL.t13 B 0.178061f
C483 VTAIL.n378 B 1.52242f
C484 VTAIL.n379 B 0.483257f
C485 VTAIL.n380 B 0.027139f
C486 VTAIL.n381 B 0.019783f
C487 VTAIL.n382 B 0.010631f
C488 VTAIL.n383 B 0.025127f
C489 VTAIL.n384 B 0.011256f
C490 VTAIL.n385 B 0.019783f
C491 VTAIL.n386 B 0.010631f
C492 VTAIL.n387 B 0.025127f
C493 VTAIL.n388 B 0.010943f
C494 VTAIL.n389 B 0.019783f
C495 VTAIL.n390 B 0.010943f
C496 VTAIL.n391 B 0.010631f
C497 VTAIL.n392 B 0.025127f
C498 VTAIL.n393 B 0.025127f
C499 VTAIL.n394 B 0.011256f
C500 VTAIL.n395 B 0.019783f
C501 VTAIL.n396 B 0.010631f
C502 VTAIL.n397 B 0.025127f
C503 VTAIL.n398 B 0.011256f
C504 VTAIL.n399 B 0.944339f
C505 VTAIL.n400 B 0.010631f
C506 VTAIL.t9 B 0.042372f
C507 VTAIL.n401 B 0.138f
C508 VTAIL.n402 B 0.017763f
C509 VTAIL.n403 B 0.018845f
C510 VTAIL.n404 B 0.025127f
C511 VTAIL.n405 B 0.011256f
C512 VTAIL.n406 B 0.010631f
C513 VTAIL.n407 B 0.019783f
C514 VTAIL.n408 B 0.019783f
C515 VTAIL.n409 B 0.010631f
C516 VTAIL.n410 B 0.011256f
C517 VTAIL.n411 B 0.025127f
C518 VTAIL.n412 B 0.025127f
C519 VTAIL.n413 B 0.011256f
C520 VTAIL.n414 B 0.010631f
C521 VTAIL.n415 B 0.019783f
C522 VTAIL.n416 B 0.019783f
C523 VTAIL.n417 B 0.010631f
C524 VTAIL.n418 B 0.011256f
C525 VTAIL.n419 B 0.025127f
C526 VTAIL.n420 B 0.025127f
C527 VTAIL.n421 B 0.011256f
C528 VTAIL.n422 B 0.010631f
C529 VTAIL.n423 B 0.019783f
C530 VTAIL.n424 B 0.019783f
C531 VTAIL.n425 B 0.010631f
C532 VTAIL.n426 B 0.011256f
C533 VTAIL.n427 B 0.025127f
C534 VTAIL.n428 B 0.025127f
C535 VTAIL.n429 B 0.011256f
C536 VTAIL.n430 B 0.010631f
C537 VTAIL.n431 B 0.019783f
C538 VTAIL.n432 B 0.019783f
C539 VTAIL.n433 B 0.010631f
C540 VTAIL.n434 B 0.011256f
C541 VTAIL.n435 B 0.025127f
C542 VTAIL.n436 B 0.053215f
C543 VTAIL.n437 B 0.011256f
C544 VTAIL.n438 B 0.010631f
C545 VTAIL.n439 B 0.045457f
C546 VTAIL.n440 B 0.029646f
C547 VTAIL.n441 B 1.19933f
C548 VTAIL.n442 B 0.027139f
C549 VTAIL.n443 B 0.019783f
C550 VTAIL.n444 B 0.010631f
C551 VTAIL.n445 B 0.025127f
C552 VTAIL.n446 B 0.011256f
C553 VTAIL.n447 B 0.019783f
C554 VTAIL.n448 B 0.010631f
C555 VTAIL.n449 B 0.025127f
C556 VTAIL.n450 B 0.010943f
C557 VTAIL.n451 B 0.019783f
C558 VTAIL.n452 B 0.011256f
C559 VTAIL.n453 B 0.025127f
C560 VTAIL.n454 B 0.011256f
C561 VTAIL.n455 B 0.019783f
C562 VTAIL.n456 B 0.010631f
C563 VTAIL.n457 B 0.025127f
C564 VTAIL.n458 B 0.011256f
C565 VTAIL.n459 B 0.944339f
C566 VTAIL.n460 B 0.010631f
C567 VTAIL.t1 B 0.042372f
C568 VTAIL.n461 B 0.138f
C569 VTAIL.n462 B 0.017763f
C570 VTAIL.n463 B 0.018845f
C571 VTAIL.n464 B 0.025127f
C572 VTAIL.n465 B 0.011256f
C573 VTAIL.n466 B 0.010631f
C574 VTAIL.n467 B 0.019783f
C575 VTAIL.n468 B 0.019783f
C576 VTAIL.n469 B 0.010631f
C577 VTAIL.n470 B 0.011256f
C578 VTAIL.n471 B 0.025127f
C579 VTAIL.n472 B 0.025127f
C580 VTAIL.n473 B 0.011256f
C581 VTAIL.n474 B 0.010631f
C582 VTAIL.n475 B 0.019783f
C583 VTAIL.n476 B 0.019783f
C584 VTAIL.n477 B 0.010631f
C585 VTAIL.n478 B 0.010631f
C586 VTAIL.n479 B 0.011256f
C587 VTAIL.n480 B 0.025127f
C588 VTAIL.n481 B 0.025127f
C589 VTAIL.n482 B 0.025127f
C590 VTAIL.n483 B 0.010943f
C591 VTAIL.n484 B 0.010631f
C592 VTAIL.n485 B 0.019783f
C593 VTAIL.n486 B 0.019783f
C594 VTAIL.n487 B 0.010631f
C595 VTAIL.n488 B 0.011256f
C596 VTAIL.n489 B 0.025127f
C597 VTAIL.n490 B 0.025127f
C598 VTAIL.n491 B 0.011256f
C599 VTAIL.n492 B 0.010631f
C600 VTAIL.n493 B 0.019783f
C601 VTAIL.n494 B 0.019783f
C602 VTAIL.n495 B 0.010631f
C603 VTAIL.n496 B 0.011256f
C604 VTAIL.n497 B 0.025127f
C605 VTAIL.n498 B 0.053215f
C606 VTAIL.n499 B 0.011256f
C607 VTAIL.n500 B 0.010631f
C608 VTAIL.n501 B 0.045457f
C609 VTAIL.n502 B 0.029646f
C610 VTAIL.n503 B 1.19562f
C611 VDD1.t0 B 0.221918f
C612 VDD1.t2 B 0.221918f
C613 VDD1.n0 B 1.97993f
C614 VDD1.t5 B 0.221918f
C615 VDD1.t3 B 0.221918f
C616 VDD1.n1 B 1.97891f
C617 VDD1.t1 B 0.221918f
C618 VDD1.t4 B 0.221918f
C619 VDD1.n2 B 1.97891f
C620 VDD1.n3 B 3.0706f
C621 VDD1.t7 B 0.221918f
C622 VDD1.t6 B 0.221918f
C623 VDD1.n4 B 1.97075f
C624 VDD1.n5 B 2.78801f
C625 VP.n0 B 0.032393f
C626 VP.t1 B 1.74341f
C627 VP.n1 B 0.025769f
C628 VP.n2 B 0.02457f
C629 VP.t7 B 1.74341f
C630 VP.n3 B 0.045792f
C631 VP.n4 B 0.02457f
C632 VP.n5 B 0.025897f
C633 VP.n6 B 0.02457f
C634 VP.n7 B 0.048162f
C635 VP.n8 B 0.032393f
C636 VP.t4 B 1.74341f
C637 VP.n9 B 0.025769f
C638 VP.n10 B 0.02457f
C639 VP.t0 B 1.74341f
C640 VP.n11 B 0.045792f
C641 VP.n12 B 0.02457f
C642 VP.n13 B 0.025897f
C643 VP.t5 B 1.89577f
C644 VP.t2 B 1.74341f
C645 VP.n14 B 0.679142f
C646 VP.n15 B 0.681148f
C647 VP.n16 B 0.210852f
C648 VP.n17 B 0.02457f
C649 VP.n18 B 0.045792f
C650 VP.n19 B 0.035867f
C651 VP.n20 B 0.035867f
C652 VP.n21 B 0.02457f
C653 VP.n22 B 0.02457f
C654 VP.n23 B 0.02457f
C655 VP.n24 B 0.025897f
C656 VP.n25 B 0.621263f
C657 VP.n26 B 0.043079f
C658 VP.n27 B 0.043595f
C659 VP.n28 B 0.02457f
C660 VP.n29 B 0.02457f
C661 VP.n30 B 0.02457f
C662 VP.n31 B 0.048162f
C663 VP.n32 B 0.031323f
C664 VP.n33 B 0.69177f
C665 VP.n34 B 1.32025f
C666 VP.n35 B 1.33831f
C667 VP.t6 B 1.74341f
C668 VP.n36 B 0.69177f
C669 VP.n37 B 0.031323f
C670 VP.n38 B 0.032393f
C671 VP.n39 B 0.02457f
C672 VP.n40 B 0.02457f
C673 VP.n41 B 0.025769f
C674 VP.n42 B 0.043595f
C675 VP.t3 B 1.74341f
C676 VP.n43 B 0.621263f
C677 VP.n44 B 0.043079f
C678 VP.n45 B 0.02457f
C679 VP.n46 B 0.02457f
C680 VP.n47 B 0.02457f
C681 VP.n48 B 0.045792f
C682 VP.n49 B 0.035867f
C683 VP.n50 B 0.035867f
C684 VP.n51 B 0.02457f
C685 VP.n52 B 0.02457f
C686 VP.n53 B 0.02457f
C687 VP.n54 B 0.025897f
C688 VP.n55 B 0.621263f
C689 VP.n56 B 0.043079f
C690 VP.n57 B 0.043595f
C691 VP.n58 B 0.02457f
C692 VP.n59 B 0.02457f
C693 VP.n60 B 0.02457f
C694 VP.n61 B 0.048162f
C695 VP.n62 B 0.031323f
C696 VP.n63 B 0.69177f
C697 VP.n64 B 0.038222f
.ends

