* NGSPICE file created from diff_pair_sample_1349.ext - technology: sky130A

.subckt diff_pair_sample_1349 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X1 VDD2.t6 VN.t1 VTAIL.t14 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X2 B.t11 B.t9 B.t10 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=1.13
X3 VTAIL.t3 VP.t0 VDD1.t7 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=1.96515 ps=12.24 w=11.91 l=1.13
X4 VTAIL.t13 VN.t2 VDD2.t1 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X5 VDD1.t6 VP.t1 VTAIL.t2 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=4.6449 ps=24.6 w=11.91 l=1.13
X6 VTAIL.t6 VP.t2 VDD1.t5 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X7 VDD2.t5 VN.t3 VTAIL.t12 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=4.6449 ps=24.6 w=11.91 l=1.13
X8 B.t8 B.t6 B.t7 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=1.13
X9 VDD2.t7 VN.t4 VTAIL.t11 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=4.6449 ps=24.6 w=11.91 l=1.13
X10 VTAIL.t0 VP.t3 VDD1.t4 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X11 VTAIL.t10 VN.t5 VDD2.t0 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=1.96515 ps=12.24 w=11.91 l=1.13
X12 VDD1.t3 VP.t4 VTAIL.t4 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X13 VTAIL.t9 VN.t6 VDD2.t4 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=1.96515 ps=12.24 w=11.91 l=1.13
X14 VDD2.t2 VN.t7 VTAIL.t8 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
X15 VTAIL.t1 VP.t5 VDD1.t2 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=1.96515 ps=12.24 w=11.91 l=1.13
X16 B.t5 B.t3 B.t4 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=1.13
X17 B.t2 B.t0 B.t1 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=4.6449 pd=24.6 as=0 ps=0 w=11.91 l=1.13
X18 VDD1.t1 VP.t6 VTAIL.t5 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=4.6449 ps=24.6 w=11.91 l=1.13
X19 VDD1.t0 VP.t7 VTAIL.t7 w_n2430_n3350# sky130_fd_pr__pfet_01v8 ad=1.96515 pd=12.24 as=1.96515 ps=12.24 w=11.91 l=1.13
R0 VN.n3 VN.t6 311.981
R1 VN.n16 VN.t3 311.981
R2 VN.n11 VN.t4 288.988
R3 VN.n24 VN.t5 288.988
R4 VN.n4 VN.t1 254.011
R5 VN.n1 VN.t2 254.011
R6 VN.n17 VN.t0 254.011
R7 VN.n14 VN.t7 254.011
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN.n11 VN.n10 50.4025
R21 VN.n24 VN.n23 50.4025
R22 VN VN.n25 44.4384
R23 VN.n4 VN.n3 33.6057
R24 VN.n17 VN.n16 33.6057
R25 VN.n16 VN.n15 28.1515
R26 VN.n3 VN.n2 28.1515
R27 VN.n10 VN.n9 24.4675
R28 VN.n23 VN.n22 24.4675
R29 VN.n5 VN.n4 23.4888
R30 VN.n6 VN.n1 23.4888
R31 VN.n18 VN.n17 23.4888
R32 VN.n19 VN.n14 23.4888
R33 VN.n9 VN.n1 0.97918
R34 VN.n22 VN.n14 0.97918
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VDD2.n2 VDD2.n1 76.8988
R45 VDD2.n2 VDD2.n0 76.8988
R46 VDD2 VDD2.n5 76.895
R47 VDD2.n4 VDD2.n3 76.325
R48 VDD2.n4 VDD2.n2 39.6463
R49 VDD2.n5 VDD2.t3 2.72972
R50 VDD2.n5 VDD2.t5 2.72972
R51 VDD2.n3 VDD2.t0 2.72972
R52 VDD2.n3 VDD2.t2 2.72972
R53 VDD2.n1 VDD2.t1 2.72972
R54 VDD2.n1 VDD2.t7 2.72972
R55 VDD2.n0 VDD2.t4 2.72972
R56 VDD2.n0 VDD2.t6 2.72972
R57 VDD2 VDD2.n4 0.688
R58 VTAIL.n534 VTAIL.n533 756.745
R59 VTAIL.n66 VTAIL.n65 756.745
R60 VTAIL.n132 VTAIL.n131 756.745
R61 VTAIL.n200 VTAIL.n199 756.745
R62 VTAIL.n468 VTAIL.n467 756.745
R63 VTAIL.n400 VTAIL.n399 756.745
R64 VTAIL.n334 VTAIL.n333 756.745
R65 VTAIL.n266 VTAIL.n265 756.745
R66 VTAIL.n493 VTAIL.n492 585
R67 VTAIL.n495 VTAIL.n494 585
R68 VTAIL.n488 VTAIL.n487 585
R69 VTAIL.n501 VTAIL.n500 585
R70 VTAIL.n503 VTAIL.n502 585
R71 VTAIL.n484 VTAIL.n483 585
R72 VTAIL.n509 VTAIL.n508 585
R73 VTAIL.n511 VTAIL.n510 585
R74 VTAIL.n480 VTAIL.n479 585
R75 VTAIL.n517 VTAIL.n516 585
R76 VTAIL.n519 VTAIL.n518 585
R77 VTAIL.n476 VTAIL.n475 585
R78 VTAIL.n525 VTAIL.n524 585
R79 VTAIL.n527 VTAIL.n526 585
R80 VTAIL.n472 VTAIL.n471 585
R81 VTAIL.n533 VTAIL.n532 585
R82 VTAIL.n25 VTAIL.n24 585
R83 VTAIL.n27 VTAIL.n26 585
R84 VTAIL.n20 VTAIL.n19 585
R85 VTAIL.n33 VTAIL.n32 585
R86 VTAIL.n35 VTAIL.n34 585
R87 VTAIL.n16 VTAIL.n15 585
R88 VTAIL.n41 VTAIL.n40 585
R89 VTAIL.n43 VTAIL.n42 585
R90 VTAIL.n12 VTAIL.n11 585
R91 VTAIL.n49 VTAIL.n48 585
R92 VTAIL.n51 VTAIL.n50 585
R93 VTAIL.n8 VTAIL.n7 585
R94 VTAIL.n57 VTAIL.n56 585
R95 VTAIL.n59 VTAIL.n58 585
R96 VTAIL.n4 VTAIL.n3 585
R97 VTAIL.n65 VTAIL.n64 585
R98 VTAIL.n91 VTAIL.n90 585
R99 VTAIL.n93 VTAIL.n92 585
R100 VTAIL.n86 VTAIL.n85 585
R101 VTAIL.n99 VTAIL.n98 585
R102 VTAIL.n101 VTAIL.n100 585
R103 VTAIL.n82 VTAIL.n81 585
R104 VTAIL.n107 VTAIL.n106 585
R105 VTAIL.n109 VTAIL.n108 585
R106 VTAIL.n78 VTAIL.n77 585
R107 VTAIL.n115 VTAIL.n114 585
R108 VTAIL.n117 VTAIL.n116 585
R109 VTAIL.n74 VTAIL.n73 585
R110 VTAIL.n123 VTAIL.n122 585
R111 VTAIL.n125 VTAIL.n124 585
R112 VTAIL.n70 VTAIL.n69 585
R113 VTAIL.n131 VTAIL.n130 585
R114 VTAIL.n159 VTAIL.n158 585
R115 VTAIL.n161 VTAIL.n160 585
R116 VTAIL.n154 VTAIL.n153 585
R117 VTAIL.n167 VTAIL.n166 585
R118 VTAIL.n169 VTAIL.n168 585
R119 VTAIL.n150 VTAIL.n149 585
R120 VTAIL.n175 VTAIL.n174 585
R121 VTAIL.n177 VTAIL.n176 585
R122 VTAIL.n146 VTAIL.n145 585
R123 VTAIL.n183 VTAIL.n182 585
R124 VTAIL.n185 VTAIL.n184 585
R125 VTAIL.n142 VTAIL.n141 585
R126 VTAIL.n191 VTAIL.n190 585
R127 VTAIL.n193 VTAIL.n192 585
R128 VTAIL.n138 VTAIL.n137 585
R129 VTAIL.n199 VTAIL.n198 585
R130 VTAIL.n467 VTAIL.n466 585
R131 VTAIL.n406 VTAIL.n405 585
R132 VTAIL.n461 VTAIL.n460 585
R133 VTAIL.n459 VTAIL.n458 585
R134 VTAIL.n410 VTAIL.n409 585
R135 VTAIL.n453 VTAIL.n452 585
R136 VTAIL.n451 VTAIL.n450 585
R137 VTAIL.n414 VTAIL.n413 585
R138 VTAIL.n445 VTAIL.n444 585
R139 VTAIL.n443 VTAIL.n442 585
R140 VTAIL.n418 VTAIL.n417 585
R141 VTAIL.n437 VTAIL.n436 585
R142 VTAIL.n435 VTAIL.n434 585
R143 VTAIL.n422 VTAIL.n421 585
R144 VTAIL.n429 VTAIL.n428 585
R145 VTAIL.n427 VTAIL.n426 585
R146 VTAIL.n399 VTAIL.n398 585
R147 VTAIL.n338 VTAIL.n337 585
R148 VTAIL.n393 VTAIL.n392 585
R149 VTAIL.n391 VTAIL.n390 585
R150 VTAIL.n342 VTAIL.n341 585
R151 VTAIL.n385 VTAIL.n384 585
R152 VTAIL.n383 VTAIL.n382 585
R153 VTAIL.n346 VTAIL.n345 585
R154 VTAIL.n377 VTAIL.n376 585
R155 VTAIL.n375 VTAIL.n374 585
R156 VTAIL.n350 VTAIL.n349 585
R157 VTAIL.n369 VTAIL.n368 585
R158 VTAIL.n367 VTAIL.n366 585
R159 VTAIL.n354 VTAIL.n353 585
R160 VTAIL.n361 VTAIL.n360 585
R161 VTAIL.n359 VTAIL.n358 585
R162 VTAIL.n333 VTAIL.n332 585
R163 VTAIL.n272 VTAIL.n271 585
R164 VTAIL.n327 VTAIL.n326 585
R165 VTAIL.n325 VTAIL.n324 585
R166 VTAIL.n276 VTAIL.n275 585
R167 VTAIL.n319 VTAIL.n318 585
R168 VTAIL.n317 VTAIL.n316 585
R169 VTAIL.n280 VTAIL.n279 585
R170 VTAIL.n311 VTAIL.n310 585
R171 VTAIL.n309 VTAIL.n308 585
R172 VTAIL.n284 VTAIL.n283 585
R173 VTAIL.n303 VTAIL.n302 585
R174 VTAIL.n301 VTAIL.n300 585
R175 VTAIL.n288 VTAIL.n287 585
R176 VTAIL.n295 VTAIL.n294 585
R177 VTAIL.n293 VTAIL.n292 585
R178 VTAIL.n265 VTAIL.n264 585
R179 VTAIL.n204 VTAIL.n203 585
R180 VTAIL.n259 VTAIL.n258 585
R181 VTAIL.n257 VTAIL.n256 585
R182 VTAIL.n208 VTAIL.n207 585
R183 VTAIL.n251 VTAIL.n250 585
R184 VTAIL.n249 VTAIL.n248 585
R185 VTAIL.n212 VTAIL.n211 585
R186 VTAIL.n243 VTAIL.n242 585
R187 VTAIL.n241 VTAIL.n240 585
R188 VTAIL.n216 VTAIL.n215 585
R189 VTAIL.n235 VTAIL.n234 585
R190 VTAIL.n233 VTAIL.n232 585
R191 VTAIL.n220 VTAIL.n219 585
R192 VTAIL.n227 VTAIL.n226 585
R193 VTAIL.n225 VTAIL.n224 585
R194 VTAIL.n425 VTAIL.t2 327.466
R195 VTAIL.n357 VTAIL.t3 327.466
R196 VTAIL.n291 VTAIL.t12 327.466
R197 VTAIL.n223 VTAIL.t10 327.466
R198 VTAIL.n491 VTAIL.t11 327.466
R199 VTAIL.n23 VTAIL.t9 327.466
R200 VTAIL.n89 VTAIL.t5 327.466
R201 VTAIL.n157 VTAIL.t1 327.466
R202 VTAIL.n494 VTAIL.n493 171.744
R203 VTAIL.n494 VTAIL.n487 171.744
R204 VTAIL.n501 VTAIL.n487 171.744
R205 VTAIL.n502 VTAIL.n501 171.744
R206 VTAIL.n502 VTAIL.n483 171.744
R207 VTAIL.n509 VTAIL.n483 171.744
R208 VTAIL.n510 VTAIL.n509 171.744
R209 VTAIL.n510 VTAIL.n479 171.744
R210 VTAIL.n517 VTAIL.n479 171.744
R211 VTAIL.n518 VTAIL.n517 171.744
R212 VTAIL.n518 VTAIL.n475 171.744
R213 VTAIL.n525 VTAIL.n475 171.744
R214 VTAIL.n526 VTAIL.n525 171.744
R215 VTAIL.n526 VTAIL.n471 171.744
R216 VTAIL.n533 VTAIL.n471 171.744
R217 VTAIL.n26 VTAIL.n25 171.744
R218 VTAIL.n26 VTAIL.n19 171.744
R219 VTAIL.n33 VTAIL.n19 171.744
R220 VTAIL.n34 VTAIL.n33 171.744
R221 VTAIL.n34 VTAIL.n15 171.744
R222 VTAIL.n41 VTAIL.n15 171.744
R223 VTAIL.n42 VTAIL.n41 171.744
R224 VTAIL.n42 VTAIL.n11 171.744
R225 VTAIL.n49 VTAIL.n11 171.744
R226 VTAIL.n50 VTAIL.n49 171.744
R227 VTAIL.n50 VTAIL.n7 171.744
R228 VTAIL.n57 VTAIL.n7 171.744
R229 VTAIL.n58 VTAIL.n57 171.744
R230 VTAIL.n58 VTAIL.n3 171.744
R231 VTAIL.n65 VTAIL.n3 171.744
R232 VTAIL.n92 VTAIL.n91 171.744
R233 VTAIL.n92 VTAIL.n85 171.744
R234 VTAIL.n99 VTAIL.n85 171.744
R235 VTAIL.n100 VTAIL.n99 171.744
R236 VTAIL.n100 VTAIL.n81 171.744
R237 VTAIL.n107 VTAIL.n81 171.744
R238 VTAIL.n108 VTAIL.n107 171.744
R239 VTAIL.n108 VTAIL.n77 171.744
R240 VTAIL.n115 VTAIL.n77 171.744
R241 VTAIL.n116 VTAIL.n115 171.744
R242 VTAIL.n116 VTAIL.n73 171.744
R243 VTAIL.n123 VTAIL.n73 171.744
R244 VTAIL.n124 VTAIL.n123 171.744
R245 VTAIL.n124 VTAIL.n69 171.744
R246 VTAIL.n131 VTAIL.n69 171.744
R247 VTAIL.n160 VTAIL.n159 171.744
R248 VTAIL.n160 VTAIL.n153 171.744
R249 VTAIL.n167 VTAIL.n153 171.744
R250 VTAIL.n168 VTAIL.n167 171.744
R251 VTAIL.n168 VTAIL.n149 171.744
R252 VTAIL.n175 VTAIL.n149 171.744
R253 VTAIL.n176 VTAIL.n175 171.744
R254 VTAIL.n176 VTAIL.n145 171.744
R255 VTAIL.n183 VTAIL.n145 171.744
R256 VTAIL.n184 VTAIL.n183 171.744
R257 VTAIL.n184 VTAIL.n141 171.744
R258 VTAIL.n191 VTAIL.n141 171.744
R259 VTAIL.n192 VTAIL.n191 171.744
R260 VTAIL.n192 VTAIL.n137 171.744
R261 VTAIL.n199 VTAIL.n137 171.744
R262 VTAIL.n467 VTAIL.n405 171.744
R263 VTAIL.n460 VTAIL.n405 171.744
R264 VTAIL.n460 VTAIL.n459 171.744
R265 VTAIL.n459 VTAIL.n409 171.744
R266 VTAIL.n452 VTAIL.n409 171.744
R267 VTAIL.n452 VTAIL.n451 171.744
R268 VTAIL.n451 VTAIL.n413 171.744
R269 VTAIL.n444 VTAIL.n413 171.744
R270 VTAIL.n444 VTAIL.n443 171.744
R271 VTAIL.n443 VTAIL.n417 171.744
R272 VTAIL.n436 VTAIL.n417 171.744
R273 VTAIL.n436 VTAIL.n435 171.744
R274 VTAIL.n435 VTAIL.n421 171.744
R275 VTAIL.n428 VTAIL.n421 171.744
R276 VTAIL.n428 VTAIL.n427 171.744
R277 VTAIL.n399 VTAIL.n337 171.744
R278 VTAIL.n392 VTAIL.n337 171.744
R279 VTAIL.n392 VTAIL.n391 171.744
R280 VTAIL.n391 VTAIL.n341 171.744
R281 VTAIL.n384 VTAIL.n341 171.744
R282 VTAIL.n384 VTAIL.n383 171.744
R283 VTAIL.n383 VTAIL.n345 171.744
R284 VTAIL.n376 VTAIL.n345 171.744
R285 VTAIL.n376 VTAIL.n375 171.744
R286 VTAIL.n375 VTAIL.n349 171.744
R287 VTAIL.n368 VTAIL.n349 171.744
R288 VTAIL.n368 VTAIL.n367 171.744
R289 VTAIL.n367 VTAIL.n353 171.744
R290 VTAIL.n360 VTAIL.n353 171.744
R291 VTAIL.n360 VTAIL.n359 171.744
R292 VTAIL.n333 VTAIL.n271 171.744
R293 VTAIL.n326 VTAIL.n271 171.744
R294 VTAIL.n326 VTAIL.n325 171.744
R295 VTAIL.n325 VTAIL.n275 171.744
R296 VTAIL.n318 VTAIL.n275 171.744
R297 VTAIL.n318 VTAIL.n317 171.744
R298 VTAIL.n317 VTAIL.n279 171.744
R299 VTAIL.n310 VTAIL.n279 171.744
R300 VTAIL.n310 VTAIL.n309 171.744
R301 VTAIL.n309 VTAIL.n283 171.744
R302 VTAIL.n302 VTAIL.n283 171.744
R303 VTAIL.n302 VTAIL.n301 171.744
R304 VTAIL.n301 VTAIL.n287 171.744
R305 VTAIL.n294 VTAIL.n287 171.744
R306 VTAIL.n294 VTAIL.n293 171.744
R307 VTAIL.n265 VTAIL.n203 171.744
R308 VTAIL.n258 VTAIL.n203 171.744
R309 VTAIL.n258 VTAIL.n257 171.744
R310 VTAIL.n257 VTAIL.n207 171.744
R311 VTAIL.n250 VTAIL.n207 171.744
R312 VTAIL.n250 VTAIL.n249 171.744
R313 VTAIL.n249 VTAIL.n211 171.744
R314 VTAIL.n242 VTAIL.n211 171.744
R315 VTAIL.n242 VTAIL.n241 171.744
R316 VTAIL.n241 VTAIL.n215 171.744
R317 VTAIL.n234 VTAIL.n215 171.744
R318 VTAIL.n234 VTAIL.n233 171.744
R319 VTAIL.n233 VTAIL.n219 171.744
R320 VTAIL.n226 VTAIL.n219 171.744
R321 VTAIL.n226 VTAIL.n225 171.744
R322 VTAIL.n493 VTAIL.t11 85.8723
R323 VTAIL.n25 VTAIL.t9 85.8723
R324 VTAIL.n91 VTAIL.t5 85.8723
R325 VTAIL.n159 VTAIL.t1 85.8723
R326 VTAIL.n427 VTAIL.t2 85.8723
R327 VTAIL.n359 VTAIL.t3 85.8723
R328 VTAIL.n293 VTAIL.t12 85.8723
R329 VTAIL.n225 VTAIL.t10 85.8723
R330 VTAIL.n403 VTAIL.n402 59.6462
R331 VTAIL.n269 VTAIL.n268 59.6462
R332 VTAIL.n1 VTAIL.n0 59.646
R333 VTAIL.n135 VTAIL.n134 59.646
R334 VTAIL.n535 VTAIL.n534 33.9308
R335 VTAIL.n67 VTAIL.n66 33.9308
R336 VTAIL.n133 VTAIL.n132 33.9308
R337 VTAIL.n201 VTAIL.n200 33.9308
R338 VTAIL.n469 VTAIL.n468 33.9308
R339 VTAIL.n401 VTAIL.n400 33.9308
R340 VTAIL.n335 VTAIL.n334 33.9308
R341 VTAIL.n267 VTAIL.n266 33.9308
R342 VTAIL.n535 VTAIL.n469 23.8927
R343 VTAIL.n267 VTAIL.n201 23.8927
R344 VTAIL.n492 VTAIL.n491 16.3895
R345 VTAIL.n24 VTAIL.n23 16.3895
R346 VTAIL.n90 VTAIL.n89 16.3895
R347 VTAIL.n158 VTAIL.n157 16.3895
R348 VTAIL.n426 VTAIL.n425 16.3895
R349 VTAIL.n358 VTAIL.n357 16.3895
R350 VTAIL.n292 VTAIL.n291 16.3895
R351 VTAIL.n224 VTAIL.n223 16.3895
R352 VTAIL.n495 VTAIL.n490 12.8005
R353 VTAIL.n27 VTAIL.n22 12.8005
R354 VTAIL.n93 VTAIL.n88 12.8005
R355 VTAIL.n161 VTAIL.n156 12.8005
R356 VTAIL.n429 VTAIL.n424 12.8005
R357 VTAIL.n361 VTAIL.n356 12.8005
R358 VTAIL.n295 VTAIL.n290 12.8005
R359 VTAIL.n227 VTAIL.n222 12.8005
R360 VTAIL.n496 VTAIL.n488 12.0247
R361 VTAIL.n532 VTAIL.n470 12.0247
R362 VTAIL.n28 VTAIL.n20 12.0247
R363 VTAIL.n64 VTAIL.n2 12.0247
R364 VTAIL.n94 VTAIL.n86 12.0247
R365 VTAIL.n130 VTAIL.n68 12.0247
R366 VTAIL.n162 VTAIL.n154 12.0247
R367 VTAIL.n198 VTAIL.n136 12.0247
R368 VTAIL.n466 VTAIL.n404 12.0247
R369 VTAIL.n430 VTAIL.n422 12.0247
R370 VTAIL.n398 VTAIL.n336 12.0247
R371 VTAIL.n362 VTAIL.n354 12.0247
R372 VTAIL.n332 VTAIL.n270 12.0247
R373 VTAIL.n296 VTAIL.n288 12.0247
R374 VTAIL.n264 VTAIL.n202 12.0247
R375 VTAIL.n228 VTAIL.n220 12.0247
R376 VTAIL.n500 VTAIL.n499 11.249
R377 VTAIL.n531 VTAIL.n472 11.249
R378 VTAIL.n32 VTAIL.n31 11.249
R379 VTAIL.n63 VTAIL.n4 11.249
R380 VTAIL.n98 VTAIL.n97 11.249
R381 VTAIL.n129 VTAIL.n70 11.249
R382 VTAIL.n166 VTAIL.n165 11.249
R383 VTAIL.n197 VTAIL.n138 11.249
R384 VTAIL.n465 VTAIL.n406 11.249
R385 VTAIL.n434 VTAIL.n433 11.249
R386 VTAIL.n397 VTAIL.n338 11.249
R387 VTAIL.n366 VTAIL.n365 11.249
R388 VTAIL.n331 VTAIL.n272 11.249
R389 VTAIL.n300 VTAIL.n299 11.249
R390 VTAIL.n263 VTAIL.n204 11.249
R391 VTAIL.n232 VTAIL.n231 11.249
R392 VTAIL.n503 VTAIL.n486 10.4732
R393 VTAIL.n528 VTAIL.n527 10.4732
R394 VTAIL.n35 VTAIL.n18 10.4732
R395 VTAIL.n60 VTAIL.n59 10.4732
R396 VTAIL.n101 VTAIL.n84 10.4732
R397 VTAIL.n126 VTAIL.n125 10.4732
R398 VTAIL.n169 VTAIL.n152 10.4732
R399 VTAIL.n194 VTAIL.n193 10.4732
R400 VTAIL.n462 VTAIL.n461 10.4732
R401 VTAIL.n437 VTAIL.n420 10.4732
R402 VTAIL.n394 VTAIL.n393 10.4732
R403 VTAIL.n369 VTAIL.n352 10.4732
R404 VTAIL.n328 VTAIL.n327 10.4732
R405 VTAIL.n303 VTAIL.n286 10.4732
R406 VTAIL.n260 VTAIL.n259 10.4732
R407 VTAIL.n235 VTAIL.n218 10.4732
R408 VTAIL.n504 VTAIL.n484 9.69747
R409 VTAIL.n524 VTAIL.n474 9.69747
R410 VTAIL.n36 VTAIL.n16 9.69747
R411 VTAIL.n56 VTAIL.n6 9.69747
R412 VTAIL.n102 VTAIL.n82 9.69747
R413 VTAIL.n122 VTAIL.n72 9.69747
R414 VTAIL.n170 VTAIL.n150 9.69747
R415 VTAIL.n190 VTAIL.n140 9.69747
R416 VTAIL.n458 VTAIL.n408 9.69747
R417 VTAIL.n438 VTAIL.n418 9.69747
R418 VTAIL.n390 VTAIL.n340 9.69747
R419 VTAIL.n370 VTAIL.n350 9.69747
R420 VTAIL.n324 VTAIL.n274 9.69747
R421 VTAIL.n304 VTAIL.n284 9.69747
R422 VTAIL.n256 VTAIL.n206 9.69747
R423 VTAIL.n236 VTAIL.n216 9.69747
R424 VTAIL.n530 VTAIL.n470 9.45567
R425 VTAIL.n62 VTAIL.n2 9.45567
R426 VTAIL.n128 VTAIL.n68 9.45567
R427 VTAIL.n196 VTAIL.n136 9.45567
R428 VTAIL.n464 VTAIL.n404 9.45567
R429 VTAIL.n396 VTAIL.n336 9.45567
R430 VTAIL.n330 VTAIL.n270 9.45567
R431 VTAIL.n262 VTAIL.n202 9.45567
R432 VTAIL.n515 VTAIL.n514 9.3005
R433 VTAIL.n478 VTAIL.n477 9.3005
R434 VTAIL.n521 VTAIL.n520 9.3005
R435 VTAIL.n523 VTAIL.n522 9.3005
R436 VTAIL.n474 VTAIL.n473 9.3005
R437 VTAIL.n529 VTAIL.n528 9.3005
R438 VTAIL.n531 VTAIL.n530 9.3005
R439 VTAIL.n482 VTAIL.n481 9.3005
R440 VTAIL.n507 VTAIL.n506 9.3005
R441 VTAIL.n505 VTAIL.n504 9.3005
R442 VTAIL.n486 VTAIL.n485 9.3005
R443 VTAIL.n499 VTAIL.n498 9.3005
R444 VTAIL.n497 VTAIL.n496 9.3005
R445 VTAIL.n490 VTAIL.n489 9.3005
R446 VTAIL.n513 VTAIL.n512 9.3005
R447 VTAIL.n47 VTAIL.n46 9.3005
R448 VTAIL.n10 VTAIL.n9 9.3005
R449 VTAIL.n53 VTAIL.n52 9.3005
R450 VTAIL.n55 VTAIL.n54 9.3005
R451 VTAIL.n6 VTAIL.n5 9.3005
R452 VTAIL.n61 VTAIL.n60 9.3005
R453 VTAIL.n63 VTAIL.n62 9.3005
R454 VTAIL.n14 VTAIL.n13 9.3005
R455 VTAIL.n39 VTAIL.n38 9.3005
R456 VTAIL.n37 VTAIL.n36 9.3005
R457 VTAIL.n18 VTAIL.n17 9.3005
R458 VTAIL.n31 VTAIL.n30 9.3005
R459 VTAIL.n29 VTAIL.n28 9.3005
R460 VTAIL.n22 VTAIL.n21 9.3005
R461 VTAIL.n45 VTAIL.n44 9.3005
R462 VTAIL.n113 VTAIL.n112 9.3005
R463 VTAIL.n76 VTAIL.n75 9.3005
R464 VTAIL.n119 VTAIL.n118 9.3005
R465 VTAIL.n121 VTAIL.n120 9.3005
R466 VTAIL.n72 VTAIL.n71 9.3005
R467 VTAIL.n127 VTAIL.n126 9.3005
R468 VTAIL.n129 VTAIL.n128 9.3005
R469 VTAIL.n80 VTAIL.n79 9.3005
R470 VTAIL.n105 VTAIL.n104 9.3005
R471 VTAIL.n103 VTAIL.n102 9.3005
R472 VTAIL.n84 VTAIL.n83 9.3005
R473 VTAIL.n97 VTAIL.n96 9.3005
R474 VTAIL.n95 VTAIL.n94 9.3005
R475 VTAIL.n88 VTAIL.n87 9.3005
R476 VTAIL.n111 VTAIL.n110 9.3005
R477 VTAIL.n181 VTAIL.n180 9.3005
R478 VTAIL.n144 VTAIL.n143 9.3005
R479 VTAIL.n187 VTAIL.n186 9.3005
R480 VTAIL.n189 VTAIL.n188 9.3005
R481 VTAIL.n140 VTAIL.n139 9.3005
R482 VTAIL.n195 VTAIL.n194 9.3005
R483 VTAIL.n197 VTAIL.n196 9.3005
R484 VTAIL.n148 VTAIL.n147 9.3005
R485 VTAIL.n173 VTAIL.n172 9.3005
R486 VTAIL.n171 VTAIL.n170 9.3005
R487 VTAIL.n152 VTAIL.n151 9.3005
R488 VTAIL.n165 VTAIL.n164 9.3005
R489 VTAIL.n163 VTAIL.n162 9.3005
R490 VTAIL.n156 VTAIL.n155 9.3005
R491 VTAIL.n179 VTAIL.n178 9.3005
R492 VTAIL.n465 VTAIL.n464 9.3005
R493 VTAIL.n463 VTAIL.n462 9.3005
R494 VTAIL.n408 VTAIL.n407 9.3005
R495 VTAIL.n457 VTAIL.n456 9.3005
R496 VTAIL.n455 VTAIL.n454 9.3005
R497 VTAIL.n412 VTAIL.n411 9.3005
R498 VTAIL.n449 VTAIL.n448 9.3005
R499 VTAIL.n447 VTAIL.n446 9.3005
R500 VTAIL.n416 VTAIL.n415 9.3005
R501 VTAIL.n441 VTAIL.n440 9.3005
R502 VTAIL.n439 VTAIL.n438 9.3005
R503 VTAIL.n420 VTAIL.n419 9.3005
R504 VTAIL.n433 VTAIL.n432 9.3005
R505 VTAIL.n431 VTAIL.n430 9.3005
R506 VTAIL.n424 VTAIL.n423 9.3005
R507 VTAIL.n344 VTAIL.n343 9.3005
R508 VTAIL.n387 VTAIL.n386 9.3005
R509 VTAIL.n389 VTAIL.n388 9.3005
R510 VTAIL.n340 VTAIL.n339 9.3005
R511 VTAIL.n395 VTAIL.n394 9.3005
R512 VTAIL.n397 VTAIL.n396 9.3005
R513 VTAIL.n381 VTAIL.n380 9.3005
R514 VTAIL.n379 VTAIL.n378 9.3005
R515 VTAIL.n348 VTAIL.n347 9.3005
R516 VTAIL.n373 VTAIL.n372 9.3005
R517 VTAIL.n371 VTAIL.n370 9.3005
R518 VTAIL.n352 VTAIL.n351 9.3005
R519 VTAIL.n365 VTAIL.n364 9.3005
R520 VTAIL.n363 VTAIL.n362 9.3005
R521 VTAIL.n356 VTAIL.n355 9.3005
R522 VTAIL.n278 VTAIL.n277 9.3005
R523 VTAIL.n321 VTAIL.n320 9.3005
R524 VTAIL.n323 VTAIL.n322 9.3005
R525 VTAIL.n274 VTAIL.n273 9.3005
R526 VTAIL.n329 VTAIL.n328 9.3005
R527 VTAIL.n331 VTAIL.n330 9.3005
R528 VTAIL.n315 VTAIL.n314 9.3005
R529 VTAIL.n313 VTAIL.n312 9.3005
R530 VTAIL.n282 VTAIL.n281 9.3005
R531 VTAIL.n307 VTAIL.n306 9.3005
R532 VTAIL.n305 VTAIL.n304 9.3005
R533 VTAIL.n286 VTAIL.n285 9.3005
R534 VTAIL.n299 VTAIL.n298 9.3005
R535 VTAIL.n297 VTAIL.n296 9.3005
R536 VTAIL.n290 VTAIL.n289 9.3005
R537 VTAIL.n210 VTAIL.n209 9.3005
R538 VTAIL.n253 VTAIL.n252 9.3005
R539 VTAIL.n255 VTAIL.n254 9.3005
R540 VTAIL.n206 VTAIL.n205 9.3005
R541 VTAIL.n261 VTAIL.n260 9.3005
R542 VTAIL.n263 VTAIL.n262 9.3005
R543 VTAIL.n247 VTAIL.n246 9.3005
R544 VTAIL.n245 VTAIL.n244 9.3005
R545 VTAIL.n214 VTAIL.n213 9.3005
R546 VTAIL.n239 VTAIL.n238 9.3005
R547 VTAIL.n237 VTAIL.n236 9.3005
R548 VTAIL.n218 VTAIL.n217 9.3005
R549 VTAIL.n231 VTAIL.n230 9.3005
R550 VTAIL.n229 VTAIL.n228 9.3005
R551 VTAIL.n222 VTAIL.n221 9.3005
R552 VTAIL.n508 VTAIL.n507 8.92171
R553 VTAIL.n523 VTAIL.n476 8.92171
R554 VTAIL.n40 VTAIL.n39 8.92171
R555 VTAIL.n55 VTAIL.n8 8.92171
R556 VTAIL.n106 VTAIL.n105 8.92171
R557 VTAIL.n121 VTAIL.n74 8.92171
R558 VTAIL.n174 VTAIL.n173 8.92171
R559 VTAIL.n189 VTAIL.n142 8.92171
R560 VTAIL.n457 VTAIL.n410 8.92171
R561 VTAIL.n442 VTAIL.n441 8.92171
R562 VTAIL.n389 VTAIL.n342 8.92171
R563 VTAIL.n374 VTAIL.n373 8.92171
R564 VTAIL.n323 VTAIL.n276 8.92171
R565 VTAIL.n308 VTAIL.n307 8.92171
R566 VTAIL.n255 VTAIL.n208 8.92171
R567 VTAIL.n240 VTAIL.n239 8.92171
R568 VTAIL.n511 VTAIL.n482 8.14595
R569 VTAIL.n520 VTAIL.n519 8.14595
R570 VTAIL.n43 VTAIL.n14 8.14595
R571 VTAIL.n52 VTAIL.n51 8.14595
R572 VTAIL.n109 VTAIL.n80 8.14595
R573 VTAIL.n118 VTAIL.n117 8.14595
R574 VTAIL.n177 VTAIL.n148 8.14595
R575 VTAIL.n186 VTAIL.n185 8.14595
R576 VTAIL.n454 VTAIL.n453 8.14595
R577 VTAIL.n445 VTAIL.n416 8.14595
R578 VTAIL.n386 VTAIL.n385 8.14595
R579 VTAIL.n377 VTAIL.n348 8.14595
R580 VTAIL.n320 VTAIL.n319 8.14595
R581 VTAIL.n311 VTAIL.n282 8.14595
R582 VTAIL.n252 VTAIL.n251 8.14595
R583 VTAIL.n243 VTAIL.n214 8.14595
R584 VTAIL.n512 VTAIL.n480 7.3702
R585 VTAIL.n516 VTAIL.n478 7.3702
R586 VTAIL.n44 VTAIL.n12 7.3702
R587 VTAIL.n48 VTAIL.n10 7.3702
R588 VTAIL.n110 VTAIL.n78 7.3702
R589 VTAIL.n114 VTAIL.n76 7.3702
R590 VTAIL.n178 VTAIL.n146 7.3702
R591 VTAIL.n182 VTAIL.n144 7.3702
R592 VTAIL.n450 VTAIL.n412 7.3702
R593 VTAIL.n446 VTAIL.n414 7.3702
R594 VTAIL.n382 VTAIL.n344 7.3702
R595 VTAIL.n378 VTAIL.n346 7.3702
R596 VTAIL.n316 VTAIL.n278 7.3702
R597 VTAIL.n312 VTAIL.n280 7.3702
R598 VTAIL.n248 VTAIL.n210 7.3702
R599 VTAIL.n244 VTAIL.n212 7.3702
R600 VTAIL.n515 VTAIL.n480 6.59444
R601 VTAIL.n516 VTAIL.n515 6.59444
R602 VTAIL.n47 VTAIL.n12 6.59444
R603 VTAIL.n48 VTAIL.n47 6.59444
R604 VTAIL.n113 VTAIL.n78 6.59444
R605 VTAIL.n114 VTAIL.n113 6.59444
R606 VTAIL.n181 VTAIL.n146 6.59444
R607 VTAIL.n182 VTAIL.n181 6.59444
R608 VTAIL.n450 VTAIL.n449 6.59444
R609 VTAIL.n449 VTAIL.n414 6.59444
R610 VTAIL.n382 VTAIL.n381 6.59444
R611 VTAIL.n381 VTAIL.n346 6.59444
R612 VTAIL.n316 VTAIL.n315 6.59444
R613 VTAIL.n315 VTAIL.n280 6.59444
R614 VTAIL.n248 VTAIL.n247 6.59444
R615 VTAIL.n247 VTAIL.n212 6.59444
R616 VTAIL.n512 VTAIL.n511 5.81868
R617 VTAIL.n519 VTAIL.n478 5.81868
R618 VTAIL.n44 VTAIL.n43 5.81868
R619 VTAIL.n51 VTAIL.n10 5.81868
R620 VTAIL.n110 VTAIL.n109 5.81868
R621 VTAIL.n117 VTAIL.n76 5.81868
R622 VTAIL.n178 VTAIL.n177 5.81868
R623 VTAIL.n185 VTAIL.n144 5.81868
R624 VTAIL.n453 VTAIL.n412 5.81868
R625 VTAIL.n446 VTAIL.n445 5.81868
R626 VTAIL.n385 VTAIL.n344 5.81868
R627 VTAIL.n378 VTAIL.n377 5.81868
R628 VTAIL.n319 VTAIL.n278 5.81868
R629 VTAIL.n312 VTAIL.n311 5.81868
R630 VTAIL.n251 VTAIL.n210 5.81868
R631 VTAIL.n244 VTAIL.n243 5.81868
R632 VTAIL.n508 VTAIL.n482 5.04292
R633 VTAIL.n520 VTAIL.n476 5.04292
R634 VTAIL.n40 VTAIL.n14 5.04292
R635 VTAIL.n52 VTAIL.n8 5.04292
R636 VTAIL.n106 VTAIL.n80 5.04292
R637 VTAIL.n118 VTAIL.n74 5.04292
R638 VTAIL.n174 VTAIL.n148 5.04292
R639 VTAIL.n186 VTAIL.n142 5.04292
R640 VTAIL.n454 VTAIL.n410 5.04292
R641 VTAIL.n442 VTAIL.n416 5.04292
R642 VTAIL.n386 VTAIL.n342 5.04292
R643 VTAIL.n374 VTAIL.n348 5.04292
R644 VTAIL.n320 VTAIL.n276 5.04292
R645 VTAIL.n308 VTAIL.n282 5.04292
R646 VTAIL.n252 VTAIL.n208 5.04292
R647 VTAIL.n240 VTAIL.n214 5.04292
R648 VTAIL.n507 VTAIL.n484 4.26717
R649 VTAIL.n524 VTAIL.n523 4.26717
R650 VTAIL.n39 VTAIL.n16 4.26717
R651 VTAIL.n56 VTAIL.n55 4.26717
R652 VTAIL.n105 VTAIL.n82 4.26717
R653 VTAIL.n122 VTAIL.n121 4.26717
R654 VTAIL.n173 VTAIL.n150 4.26717
R655 VTAIL.n190 VTAIL.n189 4.26717
R656 VTAIL.n458 VTAIL.n457 4.26717
R657 VTAIL.n441 VTAIL.n418 4.26717
R658 VTAIL.n390 VTAIL.n389 4.26717
R659 VTAIL.n373 VTAIL.n350 4.26717
R660 VTAIL.n324 VTAIL.n323 4.26717
R661 VTAIL.n307 VTAIL.n284 4.26717
R662 VTAIL.n256 VTAIL.n255 4.26717
R663 VTAIL.n239 VTAIL.n216 4.26717
R664 VTAIL.n425 VTAIL.n423 3.70982
R665 VTAIL.n357 VTAIL.n355 3.70982
R666 VTAIL.n291 VTAIL.n289 3.70982
R667 VTAIL.n223 VTAIL.n221 3.70982
R668 VTAIL.n491 VTAIL.n489 3.70982
R669 VTAIL.n23 VTAIL.n21 3.70982
R670 VTAIL.n89 VTAIL.n87 3.70982
R671 VTAIL.n157 VTAIL.n155 3.70982
R672 VTAIL.n504 VTAIL.n503 3.49141
R673 VTAIL.n527 VTAIL.n474 3.49141
R674 VTAIL.n36 VTAIL.n35 3.49141
R675 VTAIL.n59 VTAIL.n6 3.49141
R676 VTAIL.n102 VTAIL.n101 3.49141
R677 VTAIL.n125 VTAIL.n72 3.49141
R678 VTAIL.n170 VTAIL.n169 3.49141
R679 VTAIL.n193 VTAIL.n140 3.49141
R680 VTAIL.n461 VTAIL.n408 3.49141
R681 VTAIL.n438 VTAIL.n437 3.49141
R682 VTAIL.n393 VTAIL.n340 3.49141
R683 VTAIL.n370 VTAIL.n369 3.49141
R684 VTAIL.n327 VTAIL.n274 3.49141
R685 VTAIL.n304 VTAIL.n303 3.49141
R686 VTAIL.n259 VTAIL.n206 3.49141
R687 VTAIL.n236 VTAIL.n235 3.49141
R688 VTAIL.n0 VTAIL.t14 2.72972
R689 VTAIL.n0 VTAIL.t13 2.72972
R690 VTAIL.n134 VTAIL.t4 2.72972
R691 VTAIL.n134 VTAIL.t6 2.72972
R692 VTAIL.n402 VTAIL.t7 2.72972
R693 VTAIL.n402 VTAIL.t0 2.72972
R694 VTAIL.n268 VTAIL.t8 2.72972
R695 VTAIL.n268 VTAIL.t15 2.72972
R696 VTAIL.n500 VTAIL.n486 2.71565
R697 VTAIL.n528 VTAIL.n472 2.71565
R698 VTAIL.n32 VTAIL.n18 2.71565
R699 VTAIL.n60 VTAIL.n4 2.71565
R700 VTAIL.n98 VTAIL.n84 2.71565
R701 VTAIL.n126 VTAIL.n70 2.71565
R702 VTAIL.n166 VTAIL.n152 2.71565
R703 VTAIL.n194 VTAIL.n138 2.71565
R704 VTAIL.n462 VTAIL.n406 2.71565
R705 VTAIL.n434 VTAIL.n420 2.71565
R706 VTAIL.n394 VTAIL.n338 2.71565
R707 VTAIL.n366 VTAIL.n352 2.71565
R708 VTAIL.n328 VTAIL.n272 2.71565
R709 VTAIL.n300 VTAIL.n286 2.71565
R710 VTAIL.n260 VTAIL.n204 2.71565
R711 VTAIL.n232 VTAIL.n218 2.71565
R712 VTAIL.n499 VTAIL.n488 1.93989
R713 VTAIL.n532 VTAIL.n531 1.93989
R714 VTAIL.n31 VTAIL.n20 1.93989
R715 VTAIL.n64 VTAIL.n63 1.93989
R716 VTAIL.n97 VTAIL.n86 1.93989
R717 VTAIL.n130 VTAIL.n129 1.93989
R718 VTAIL.n165 VTAIL.n154 1.93989
R719 VTAIL.n198 VTAIL.n197 1.93989
R720 VTAIL.n466 VTAIL.n465 1.93989
R721 VTAIL.n433 VTAIL.n422 1.93989
R722 VTAIL.n398 VTAIL.n397 1.93989
R723 VTAIL.n365 VTAIL.n354 1.93989
R724 VTAIL.n332 VTAIL.n331 1.93989
R725 VTAIL.n299 VTAIL.n288 1.93989
R726 VTAIL.n264 VTAIL.n263 1.93989
R727 VTAIL.n231 VTAIL.n220 1.93989
R728 VTAIL.n269 VTAIL.n267 1.25912
R729 VTAIL.n335 VTAIL.n269 1.25912
R730 VTAIL.n403 VTAIL.n401 1.25912
R731 VTAIL.n469 VTAIL.n403 1.25912
R732 VTAIL.n201 VTAIL.n135 1.25912
R733 VTAIL.n135 VTAIL.n133 1.25912
R734 VTAIL.n67 VTAIL.n1 1.25912
R735 VTAIL VTAIL.n535 1.20093
R736 VTAIL.n496 VTAIL.n495 1.16414
R737 VTAIL.n534 VTAIL.n470 1.16414
R738 VTAIL.n28 VTAIL.n27 1.16414
R739 VTAIL.n66 VTAIL.n2 1.16414
R740 VTAIL.n94 VTAIL.n93 1.16414
R741 VTAIL.n132 VTAIL.n68 1.16414
R742 VTAIL.n162 VTAIL.n161 1.16414
R743 VTAIL.n200 VTAIL.n136 1.16414
R744 VTAIL.n468 VTAIL.n404 1.16414
R745 VTAIL.n430 VTAIL.n429 1.16414
R746 VTAIL.n400 VTAIL.n336 1.16414
R747 VTAIL.n362 VTAIL.n361 1.16414
R748 VTAIL.n334 VTAIL.n270 1.16414
R749 VTAIL.n296 VTAIL.n295 1.16414
R750 VTAIL.n266 VTAIL.n202 1.16414
R751 VTAIL.n228 VTAIL.n227 1.16414
R752 VTAIL.n401 VTAIL.n335 0.470328
R753 VTAIL.n133 VTAIL.n67 0.470328
R754 VTAIL.n492 VTAIL.n490 0.388379
R755 VTAIL.n24 VTAIL.n22 0.388379
R756 VTAIL.n90 VTAIL.n88 0.388379
R757 VTAIL.n158 VTAIL.n156 0.388379
R758 VTAIL.n426 VTAIL.n424 0.388379
R759 VTAIL.n358 VTAIL.n356 0.388379
R760 VTAIL.n292 VTAIL.n290 0.388379
R761 VTAIL.n224 VTAIL.n222 0.388379
R762 VTAIL.n497 VTAIL.n489 0.155672
R763 VTAIL.n498 VTAIL.n497 0.155672
R764 VTAIL.n498 VTAIL.n485 0.155672
R765 VTAIL.n505 VTAIL.n485 0.155672
R766 VTAIL.n506 VTAIL.n505 0.155672
R767 VTAIL.n506 VTAIL.n481 0.155672
R768 VTAIL.n513 VTAIL.n481 0.155672
R769 VTAIL.n514 VTAIL.n513 0.155672
R770 VTAIL.n514 VTAIL.n477 0.155672
R771 VTAIL.n521 VTAIL.n477 0.155672
R772 VTAIL.n522 VTAIL.n521 0.155672
R773 VTAIL.n522 VTAIL.n473 0.155672
R774 VTAIL.n529 VTAIL.n473 0.155672
R775 VTAIL.n530 VTAIL.n529 0.155672
R776 VTAIL.n29 VTAIL.n21 0.155672
R777 VTAIL.n30 VTAIL.n29 0.155672
R778 VTAIL.n30 VTAIL.n17 0.155672
R779 VTAIL.n37 VTAIL.n17 0.155672
R780 VTAIL.n38 VTAIL.n37 0.155672
R781 VTAIL.n38 VTAIL.n13 0.155672
R782 VTAIL.n45 VTAIL.n13 0.155672
R783 VTAIL.n46 VTAIL.n45 0.155672
R784 VTAIL.n46 VTAIL.n9 0.155672
R785 VTAIL.n53 VTAIL.n9 0.155672
R786 VTAIL.n54 VTAIL.n53 0.155672
R787 VTAIL.n54 VTAIL.n5 0.155672
R788 VTAIL.n61 VTAIL.n5 0.155672
R789 VTAIL.n62 VTAIL.n61 0.155672
R790 VTAIL.n95 VTAIL.n87 0.155672
R791 VTAIL.n96 VTAIL.n95 0.155672
R792 VTAIL.n96 VTAIL.n83 0.155672
R793 VTAIL.n103 VTAIL.n83 0.155672
R794 VTAIL.n104 VTAIL.n103 0.155672
R795 VTAIL.n104 VTAIL.n79 0.155672
R796 VTAIL.n111 VTAIL.n79 0.155672
R797 VTAIL.n112 VTAIL.n111 0.155672
R798 VTAIL.n112 VTAIL.n75 0.155672
R799 VTAIL.n119 VTAIL.n75 0.155672
R800 VTAIL.n120 VTAIL.n119 0.155672
R801 VTAIL.n120 VTAIL.n71 0.155672
R802 VTAIL.n127 VTAIL.n71 0.155672
R803 VTAIL.n128 VTAIL.n127 0.155672
R804 VTAIL.n163 VTAIL.n155 0.155672
R805 VTAIL.n164 VTAIL.n163 0.155672
R806 VTAIL.n164 VTAIL.n151 0.155672
R807 VTAIL.n171 VTAIL.n151 0.155672
R808 VTAIL.n172 VTAIL.n171 0.155672
R809 VTAIL.n172 VTAIL.n147 0.155672
R810 VTAIL.n179 VTAIL.n147 0.155672
R811 VTAIL.n180 VTAIL.n179 0.155672
R812 VTAIL.n180 VTAIL.n143 0.155672
R813 VTAIL.n187 VTAIL.n143 0.155672
R814 VTAIL.n188 VTAIL.n187 0.155672
R815 VTAIL.n188 VTAIL.n139 0.155672
R816 VTAIL.n195 VTAIL.n139 0.155672
R817 VTAIL.n196 VTAIL.n195 0.155672
R818 VTAIL.n464 VTAIL.n463 0.155672
R819 VTAIL.n463 VTAIL.n407 0.155672
R820 VTAIL.n456 VTAIL.n407 0.155672
R821 VTAIL.n456 VTAIL.n455 0.155672
R822 VTAIL.n455 VTAIL.n411 0.155672
R823 VTAIL.n448 VTAIL.n411 0.155672
R824 VTAIL.n448 VTAIL.n447 0.155672
R825 VTAIL.n447 VTAIL.n415 0.155672
R826 VTAIL.n440 VTAIL.n415 0.155672
R827 VTAIL.n440 VTAIL.n439 0.155672
R828 VTAIL.n439 VTAIL.n419 0.155672
R829 VTAIL.n432 VTAIL.n419 0.155672
R830 VTAIL.n432 VTAIL.n431 0.155672
R831 VTAIL.n431 VTAIL.n423 0.155672
R832 VTAIL.n396 VTAIL.n395 0.155672
R833 VTAIL.n395 VTAIL.n339 0.155672
R834 VTAIL.n388 VTAIL.n339 0.155672
R835 VTAIL.n388 VTAIL.n387 0.155672
R836 VTAIL.n387 VTAIL.n343 0.155672
R837 VTAIL.n380 VTAIL.n343 0.155672
R838 VTAIL.n380 VTAIL.n379 0.155672
R839 VTAIL.n379 VTAIL.n347 0.155672
R840 VTAIL.n372 VTAIL.n347 0.155672
R841 VTAIL.n372 VTAIL.n371 0.155672
R842 VTAIL.n371 VTAIL.n351 0.155672
R843 VTAIL.n364 VTAIL.n351 0.155672
R844 VTAIL.n364 VTAIL.n363 0.155672
R845 VTAIL.n363 VTAIL.n355 0.155672
R846 VTAIL.n330 VTAIL.n329 0.155672
R847 VTAIL.n329 VTAIL.n273 0.155672
R848 VTAIL.n322 VTAIL.n273 0.155672
R849 VTAIL.n322 VTAIL.n321 0.155672
R850 VTAIL.n321 VTAIL.n277 0.155672
R851 VTAIL.n314 VTAIL.n277 0.155672
R852 VTAIL.n314 VTAIL.n313 0.155672
R853 VTAIL.n313 VTAIL.n281 0.155672
R854 VTAIL.n306 VTAIL.n281 0.155672
R855 VTAIL.n306 VTAIL.n305 0.155672
R856 VTAIL.n305 VTAIL.n285 0.155672
R857 VTAIL.n298 VTAIL.n285 0.155672
R858 VTAIL.n298 VTAIL.n297 0.155672
R859 VTAIL.n297 VTAIL.n289 0.155672
R860 VTAIL.n262 VTAIL.n261 0.155672
R861 VTAIL.n261 VTAIL.n205 0.155672
R862 VTAIL.n254 VTAIL.n205 0.155672
R863 VTAIL.n254 VTAIL.n253 0.155672
R864 VTAIL.n253 VTAIL.n209 0.155672
R865 VTAIL.n246 VTAIL.n209 0.155672
R866 VTAIL.n246 VTAIL.n245 0.155672
R867 VTAIL.n245 VTAIL.n213 0.155672
R868 VTAIL.n238 VTAIL.n213 0.155672
R869 VTAIL.n238 VTAIL.n237 0.155672
R870 VTAIL.n237 VTAIL.n217 0.155672
R871 VTAIL.n230 VTAIL.n217 0.155672
R872 VTAIL.n230 VTAIL.n229 0.155672
R873 VTAIL.n229 VTAIL.n221 0.155672
R874 VTAIL VTAIL.n1 0.0586897
R875 B.n342 B.n97 585
R876 B.n341 B.n340 585
R877 B.n339 B.n98 585
R878 B.n338 B.n337 585
R879 B.n336 B.n99 585
R880 B.n335 B.n334 585
R881 B.n333 B.n100 585
R882 B.n332 B.n331 585
R883 B.n330 B.n101 585
R884 B.n329 B.n328 585
R885 B.n327 B.n102 585
R886 B.n326 B.n325 585
R887 B.n324 B.n103 585
R888 B.n323 B.n322 585
R889 B.n321 B.n104 585
R890 B.n320 B.n319 585
R891 B.n318 B.n105 585
R892 B.n317 B.n316 585
R893 B.n315 B.n106 585
R894 B.n314 B.n313 585
R895 B.n312 B.n107 585
R896 B.n311 B.n310 585
R897 B.n309 B.n108 585
R898 B.n308 B.n307 585
R899 B.n306 B.n109 585
R900 B.n305 B.n304 585
R901 B.n303 B.n110 585
R902 B.n302 B.n301 585
R903 B.n300 B.n111 585
R904 B.n299 B.n298 585
R905 B.n297 B.n112 585
R906 B.n296 B.n295 585
R907 B.n294 B.n113 585
R908 B.n293 B.n292 585
R909 B.n291 B.n114 585
R910 B.n290 B.n289 585
R911 B.n288 B.n115 585
R912 B.n287 B.n286 585
R913 B.n285 B.n116 585
R914 B.n284 B.n283 585
R915 B.n282 B.n117 585
R916 B.n280 B.n279 585
R917 B.n278 B.n120 585
R918 B.n277 B.n276 585
R919 B.n275 B.n121 585
R920 B.n274 B.n273 585
R921 B.n272 B.n122 585
R922 B.n271 B.n270 585
R923 B.n269 B.n123 585
R924 B.n268 B.n267 585
R925 B.n266 B.n124 585
R926 B.n265 B.n264 585
R927 B.n260 B.n125 585
R928 B.n259 B.n258 585
R929 B.n257 B.n126 585
R930 B.n256 B.n255 585
R931 B.n254 B.n127 585
R932 B.n253 B.n252 585
R933 B.n251 B.n128 585
R934 B.n250 B.n249 585
R935 B.n248 B.n129 585
R936 B.n247 B.n246 585
R937 B.n245 B.n130 585
R938 B.n244 B.n243 585
R939 B.n242 B.n131 585
R940 B.n241 B.n240 585
R941 B.n239 B.n132 585
R942 B.n238 B.n237 585
R943 B.n236 B.n133 585
R944 B.n235 B.n234 585
R945 B.n233 B.n134 585
R946 B.n232 B.n231 585
R947 B.n230 B.n135 585
R948 B.n229 B.n228 585
R949 B.n227 B.n136 585
R950 B.n226 B.n225 585
R951 B.n224 B.n137 585
R952 B.n223 B.n222 585
R953 B.n221 B.n138 585
R954 B.n220 B.n219 585
R955 B.n218 B.n139 585
R956 B.n217 B.n216 585
R957 B.n215 B.n140 585
R958 B.n214 B.n213 585
R959 B.n212 B.n141 585
R960 B.n211 B.n210 585
R961 B.n209 B.n142 585
R962 B.n208 B.n207 585
R963 B.n206 B.n143 585
R964 B.n205 B.n204 585
R965 B.n203 B.n144 585
R966 B.n202 B.n201 585
R967 B.n344 B.n343 585
R968 B.n345 B.n96 585
R969 B.n347 B.n346 585
R970 B.n348 B.n95 585
R971 B.n350 B.n349 585
R972 B.n351 B.n94 585
R973 B.n353 B.n352 585
R974 B.n354 B.n93 585
R975 B.n356 B.n355 585
R976 B.n357 B.n92 585
R977 B.n359 B.n358 585
R978 B.n360 B.n91 585
R979 B.n362 B.n361 585
R980 B.n363 B.n90 585
R981 B.n365 B.n364 585
R982 B.n366 B.n89 585
R983 B.n368 B.n367 585
R984 B.n369 B.n88 585
R985 B.n371 B.n370 585
R986 B.n372 B.n87 585
R987 B.n374 B.n373 585
R988 B.n375 B.n86 585
R989 B.n377 B.n376 585
R990 B.n378 B.n85 585
R991 B.n380 B.n379 585
R992 B.n381 B.n84 585
R993 B.n383 B.n382 585
R994 B.n384 B.n83 585
R995 B.n386 B.n385 585
R996 B.n387 B.n82 585
R997 B.n389 B.n388 585
R998 B.n390 B.n81 585
R999 B.n392 B.n391 585
R1000 B.n393 B.n80 585
R1001 B.n395 B.n394 585
R1002 B.n396 B.n79 585
R1003 B.n398 B.n397 585
R1004 B.n399 B.n78 585
R1005 B.n401 B.n400 585
R1006 B.n402 B.n77 585
R1007 B.n404 B.n403 585
R1008 B.n405 B.n76 585
R1009 B.n407 B.n406 585
R1010 B.n408 B.n75 585
R1011 B.n410 B.n409 585
R1012 B.n411 B.n74 585
R1013 B.n413 B.n412 585
R1014 B.n414 B.n73 585
R1015 B.n416 B.n415 585
R1016 B.n417 B.n72 585
R1017 B.n419 B.n418 585
R1018 B.n420 B.n71 585
R1019 B.n422 B.n421 585
R1020 B.n423 B.n70 585
R1021 B.n425 B.n424 585
R1022 B.n426 B.n69 585
R1023 B.n428 B.n427 585
R1024 B.n429 B.n68 585
R1025 B.n431 B.n430 585
R1026 B.n432 B.n67 585
R1027 B.n572 B.n571 585
R1028 B.n570 B.n17 585
R1029 B.n569 B.n568 585
R1030 B.n567 B.n18 585
R1031 B.n566 B.n565 585
R1032 B.n564 B.n19 585
R1033 B.n563 B.n562 585
R1034 B.n561 B.n20 585
R1035 B.n560 B.n559 585
R1036 B.n558 B.n21 585
R1037 B.n557 B.n556 585
R1038 B.n555 B.n22 585
R1039 B.n554 B.n553 585
R1040 B.n552 B.n23 585
R1041 B.n551 B.n550 585
R1042 B.n549 B.n24 585
R1043 B.n548 B.n547 585
R1044 B.n546 B.n25 585
R1045 B.n545 B.n544 585
R1046 B.n543 B.n26 585
R1047 B.n542 B.n541 585
R1048 B.n540 B.n27 585
R1049 B.n539 B.n538 585
R1050 B.n537 B.n28 585
R1051 B.n536 B.n535 585
R1052 B.n534 B.n29 585
R1053 B.n533 B.n532 585
R1054 B.n531 B.n30 585
R1055 B.n530 B.n529 585
R1056 B.n528 B.n31 585
R1057 B.n527 B.n526 585
R1058 B.n525 B.n32 585
R1059 B.n524 B.n523 585
R1060 B.n522 B.n33 585
R1061 B.n521 B.n520 585
R1062 B.n519 B.n34 585
R1063 B.n518 B.n517 585
R1064 B.n516 B.n35 585
R1065 B.n515 B.n514 585
R1066 B.n513 B.n36 585
R1067 B.n512 B.n511 585
R1068 B.n509 B.n37 585
R1069 B.n508 B.n507 585
R1070 B.n506 B.n40 585
R1071 B.n505 B.n504 585
R1072 B.n503 B.n41 585
R1073 B.n502 B.n501 585
R1074 B.n500 B.n42 585
R1075 B.n499 B.n498 585
R1076 B.n497 B.n43 585
R1077 B.n496 B.n495 585
R1078 B.n494 B.n493 585
R1079 B.n492 B.n47 585
R1080 B.n491 B.n490 585
R1081 B.n489 B.n48 585
R1082 B.n488 B.n487 585
R1083 B.n486 B.n49 585
R1084 B.n485 B.n484 585
R1085 B.n483 B.n50 585
R1086 B.n482 B.n481 585
R1087 B.n480 B.n51 585
R1088 B.n479 B.n478 585
R1089 B.n477 B.n52 585
R1090 B.n476 B.n475 585
R1091 B.n474 B.n53 585
R1092 B.n473 B.n472 585
R1093 B.n471 B.n54 585
R1094 B.n470 B.n469 585
R1095 B.n468 B.n55 585
R1096 B.n467 B.n466 585
R1097 B.n465 B.n56 585
R1098 B.n464 B.n463 585
R1099 B.n462 B.n57 585
R1100 B.n461 B.n460 585
R1101 B.n459 B.n58 585
R1102 B.n458 B.n457 585
R1103 B.n456 B.n59 585
R1104 B.n455 B.n454 585
R1105 B.n453 B.n60 585
R1106 B.n452 B.n451 585
R1107 B.n450 B.n61 585
R1108 B.n449 B.n448 585
R1109 B.n447 B.n62 585
R1110 B.n446 B.n445 585
R1111 B.n444 B.n63 585
R1112 B.n443 B.n442 585
R1113 B.n441 B.n64 585
R1114 B.n440 B.n439 585
R1115 B.n438 B.n65 585
R1116 B.n437 B.n436 585
R1117 B.n435 B.n66 585
R1118 B.n434 B.n433 585
R1119 B.n573 B.n16 585
R1120 B.n575 B.n574 585
R1121 B.n576 B.n15 585
R1122 B.n578 B.n577 585
R1123 B.n579 B.n14 585
R1124 B.n581 B.n580 585
R1125 B.n582 B.n13 585
R1126 B.n584 B.n583 585
R1127 B.n585 B.n12 585
R1128 B.n587 B.n586 585
R1129 B.n588 B.n11 585
R1130 B.n590 B.n589 585
R1131 B.n591 B.n10 585
R1132 B.n593 B.n592 585
R1133 B.n594 B.n9 585
R1134 B.n596 B.n595 585
R1135 B.n597 B.n8 585
R1136 B.n599 B.n598 585
R1137 B.n600 B.n7 585
R1138 B.n602 B.n601 585
R1139 B.n603 B.n6 585
R1140 B.n605 B.n604 585
R1141 B.n606 B.n5 585
R1142 B.n608 B.n607 585
R1143 B.n609 B.n4 585
R1144 B.n611 B.n610 585
R1145 B.n612 B.n3 585
R1146 B.n614 B.n613 585
R1147 B.n615 B.n0 585
R1148 B.n2 B.n1 585
R1149 B.n160 B.n159 585
R1150 B.n161 B.n158 585
R1151 B.n163 B.n162 585
R1152 B.n164 B.n157 585
R1153 B.n166 B.n165 585
R1154 B.n167 B.n156 585
R1155 B.n169 B.n168 585
R1156 B.n170 B.n155 585
R1157 B.n172 B.n171 585
R1158 B.n173 B.n154 585
R1159 B.n175 B.n174 585
R1160 B.n176 B.n153 585
R1161 B.n178 B.n177 585
R1162 B.n179 B.n152 585
R1163 B.n181 B.n180 585
R1164 B.n182 B.n151 585
R1165 B.n184 B.n183 585
R1166 B.n185 B.n150 585
R1167 B.n187 B.n186 585
R1168 B.n188 B.n149 585
R1169 B.n190 B.n189 585
R1170 B.n191 B.n148 585
R1171 B.n193 B.n192 585
R1172 B.n194 B.n147 585
R1173 B.n196 B.n195 585
R1174 B.n197 B.n146 585
R1175 B.n199 B.n198 585
R1176 B.n200 B.n145 585
R1177 B.n202 B.n145 535.745
R1178 B.n344 B.n97 535.745
R1179 B.n434 B.n67 535.745
R1180 B.n573 B.n572 535.745
R1181 B.n261 B.t6 457.745
R1182 B.n118 B.t0 457.745
R1183 B.n44 B.t9 457.745
R1184 B.n38 B.t3 457.745
R1185 B.n118 B.t1 402.099
R1186 B.n44 B.t11 402.099
R1187 B.n261 B.t7 402.099
R1188 B.n38 B.t5 402.099
R1189 B.n119 B.t2 373.784
R1190 B.n45 B.t10 373.784
R1191 B.n262 B.t8 373.784
R1192 B.n39 B.t4 373.784
R1193 B.n617 B.n616 256.663
R1194 B.n616 B.n615 235.042
R1195 B.n616 B.n2 235.042
R1196 B.n203 B.n202 163.367
R1197 B.n204 B.n203 163.367
R1198 B.n204 B.n143 163.367
R1199 B.n208 B.n143 163.367
R1200 B.n209 B.n208 163.367
R1201 B.n210 B.n209 163.367
R1202 B.n210 B.n141 163.367
R1203 B.n214 B.n141 163.367
R1204 B.n215 B.n214 163.367
R1205 B.n216 B.n215 163.367
R1206 B.n216 B.n139 163.367
R1207 B.n220 B.n139 163.367
R1208 B.n221 B.n220 163.367
R1209 B.n222 B.n221 163.367
R1210 B.n222 B.n137 163.367
R1211 B.n226 B.n137 163.367
R1212 B.n227 B.n226 163.367
R1213 B.n228 B.n227 163.367
R1214 B.n228 B.n135 163.367
R1215 B.n232 B.n135 163.367
R1216 B.n233 B.n232 163.367
R1217 B.n234 B.n233 163.367
R1218 B.n234 B.n133 163.367
R1219 B.n238 B.n133 163.367
R1220 B.n239 B.n238 163.367
R1221 B.n240 B.n239 163.367
R1222 B.n240 B.n131 163.367
R1223 B.n244 B.n131 163.367
R1224 B.n245 B.n244 163.367
R1225 B.n246 B.n245 163.367
R1226 B.n246 B.n129 163.367
R1227 B.n250 B.n129 163.367
R1228 B.n251 B.n250 163.367
R1229 B.n252 B.n251 163.367
R1230 B.n252 B.n127 163.367
R1231 B.n256 B.n127 163.367
R1232 B.n257 B.n256 163.367
R1233 B.n258 B.n257 163.367
R1234 B.n258 B.n125 163.367
R1235 B.n265 B.n125 163.367
R1236 B.n266 B.n265 163.367
R1237 B.n267 B.n266 163.367
R1238 B.n267 B.n123 163.367
R1239 B.n271 B.n123 163.367
R1240 B.n272 B.n271 163.367
R1241 B.n273 B.n272 163.367
R1242 B.n273 B.n121 163.367
R1243 B.n277 B.n121 163.367
R1244 B.n278 B.n277 163.367
R1245 B.n279 B.n278 163.367
R1246 B.n279 B.n117 163.367
R1247 B.n284 B.n117 163.367
R1248 B.n285 B.n284 163.367
R1249 B.n286 B.n285 163.367
R1250 B.n286 B.n115 163.367
R1251 B.n290 B.n115 163.367
R1252 B.n291 B.n290 163.367
R1253 B.n292 B.n291 163.367
R1254 B.n292 B.n113 163.367
R1255 B.n296 B.n113 163.367
R1256 B.n297 B.n296 163.367
R1257 B.n298 B.n297 163.367
R1258 B.n298 B.n111 163.367
R1259 B.n302 B.n111 163.367
R1260 B.n303 B.n302 163.367
R1261 B.n304 B.n303 163.367
R1262 B.n304 B.n109 163.367
R1263 B.n308 B.n109 163.367
R1264 B.n309 B.n308 163.367
R1265 B.n310 B.n309 163.367
R1266 B.n310 B.n107 163.367
R1267 B.n314 B.n107 163.367
R1268 B.n315 B.n314 163.367
R1269 B.n316 B.n315 163.367
R1270 B.n316 B.n105 163.367
R1271 B.n320 B.n105 163.367
R1272 B.n321 B.n320 163.367
R1273 B.n322 B.n321 163.367
R1274 B.n322 B.n103 163.367
R1275 B.n326 B.n103 163.367
R1276 B.n327 B.n326 163.367
R1277 B.n328 B.n327 163.367
R1278 B.n328 B.n101 163.367
R1279 B.n332 B.n101 163.367
R1280 B.n333 B.n332 163.367
R1281 B.n334 B.n333 163.367
R1282 B.n334 B.n99 163.367
R1283 B.n338 B.n99 163.367
R1284 B.n339 B.n338 163.367
R1285 B.n340 B.n339 163.367
R1286 B.n340 B.n97 163.367
R1287 B.n430 B.n67 163.367
R1288 B.n430 B.n429 163.367
R1289 B.n429 B.n428 163.367
R1290 B.n428 B.n69 163.367
R1291 B.n424 B.n69 163.367
R1292 B.n424 B.n423 163.367
R1293 B.n423 B.n422 163.367
R1294 B.n422 B.n71 163.367
R1295 B.n418 B.n71 163.367
R1296 B.n418 B.n417 163.367
R1297 B.n417 B.n416 163.367
R1298 B.n416 B.n73 163.367
R1299 B.n412 B.n73 163.367
R1300 B.n412 B.n411 163.367
R1301 B.n411 B.n410 163.367
R1302 B.n410 B.n75 163.367
R1303 B.n406 B.n75 163.367
R1304 B.n406 B.n405 163.367
R1305 B.n405 B.n404 163.367
R1306 B.n404 B.n77 163.367
R1307 B.n400 B.n77 163.367
R1308 B.n400 B.n399 163.367
R1309 B.n399 B.n398 163.367
R1310 B.n398 B.n79 163.367
R1311 B.n394 B.n79 163.367
R1312 B.n394 B.n393 163.367
R1313 B.n393 B.n392 163.367
R1314 B.n392 B.n81 163.367
R1315 B.n388 B.n81 163.367
R1316 B.n388 B.n387 163.367
R1317 B.n387 B.n386 163.367
R1318 B.n386 B.n83 163.367
R1319 B.n382 B.n83 163.367
R1320 B.n382 B.n381 163.367
R1321 B.n381 B.n380 163.367
R1322 B.n380 B.n85 163.367
R1323 B.n376 B.n85 163.367
R1324 B.n376 B.n375 163.367
R1325 B.n375 B.n374 163.367
R1326 B.n374 B.n87 163.367
R1327 B.n370 B.n87 163.367
R1328 B.n370 B.n369 163.367
R1329 B.n369 B.n368 163.367
R1330 B.n368 B.n89 163.367
R1331 B.n364 B.n89 163.367
R1332 B.n364 B.n363 163.367
R1333 B.n363 B.n362 163.367
R1334 B.n362 B.n91 163.367
R1335 B.n358 B.n91 163.367
R1336 B.n358 B.n357 163.367
R1337 B.n357 B.n356 163.367
R1338 B.n356 B.n93 163.367
R1339 B.n352 B.n93 163.367
R1340 B.n352 B.n351 163.367
R1341 B.n351 B.n350 163.367
R1342 B.n350 B.n95 163.367
R1343 B.n346 B.n95 163.367
R1344 B.n346 B.n345 163.367
R1345 B.n345 B.n344 163.367
R1346 B.n572 B.n17 163.367
R1347 B.n568 B.n17 163.367
R1348 B.n568 B.n567 163.367
R1349 B.n567 B.n566 163.367
R1350 B.n566 B.n19 163.367
R1351 B.n562 B.n19 163.367
R1352 B.n562 B.n561 163.367
R1353 B.n561 B.n560 163.367
R1354 B.n560 B.n21 163.367
R1355 B.n556 B.n21 163.367
R1356 B.n556 B.n555 163.367
R1357 B.n555 B.n554 163.367
R1358 B.n554 B.n23 163.367
R1359 B.n550 B.n23 163.367
R1360 B.n550 B.n549 163.367
R1361 B.n549 B.n548 163.367
R1362 B.n548 B.n25 163.367
R1363 B.n544 B.n25 163.367
R1364 B.n544 B.n543 163.367
R1365 B.n543 B.n542 163.367
R1366 B.n542 B.n27 163.367
R1367 B.n538 B.n27 163.367
R1368 B.n538 B.n537 163.367
R1369 B.n537 B.n536 163.367
R1370 B.n536 B.n29 163.367
R1371 B.n532 B.n29 163.367
R1372 B.n532 B.n531 163.367
R1373 B.n531 B.n530 163.367
R1374 B.n530 B.n31 163.367
R1375 B.n526 B.n31 163.367
R1376 B.n526 B.n525 163.367
R1377 B.n525 B.n524 163.367
R1378 B.n524 B.n33 163.367
R1379 B.n520 B.n33 163.367
R1380 B.n520 B.n519 163.367
R1381 B.n519 B.n518 163.367
R1382 B.n518 B.n35 163.367
R1383 B.n514 B.n35 163.367
R1384 B.n514 B.n513 163.367
R1385 B.n513 B.n512 163.367
R1386 B.n512 B.n37 163.367
R1387 B.n507 B.n37 163.367
R1388 B.n507 B.n506 163.367
R1389 B.n506 B.n505 163.367
R1390 B.n505 B.n41 163.367
R1391 B.n501 B.n41 163.367
R1392 B.n501 B.n500 163.367
R1393 B.n500 B.n499 163.367
R1394 B.n499 B.n43 163.367
R1395 B.n495 B.n43 163.367
R1396 B.n495 B.n494 163.367
R1397 B.n494 B.n47 163.367
R1398 B.n490 B.n47 163.367
R1399 B.n490 B.n489 163.367
R1400 B.n489 B.n488 163.367
R1401 B.n488 B.n49 163.367
R1402 B.n484 B.n49 163.367
R1403 B.n484 B.n483 163.367
R1404 B.n483 B.n482 163.367
R1405 B.n482 B.n51 163.367
R1406 B.n478 B.n51 163.367
R1407 B.n478 B.n477 163.367
R1408 B.n477 B.n476 163.367
R1409 B.n476 B.n53 163.367
R1410 B.n472 B.n53 163.367
R1411 B.n472 B.n471 163.367
R1412 B.n471 B.n470 163.367
R1413 B.n470 B.n55 163.367
R1414 B.n466 B.n55 163.367
R1415 B.n466 B.n465 163.367
R1416 B.n465 B.n464 163.367
R1417 B.n464 B.n57 163.367
R1418 B.n460 B.n57 163.367
R1419 B.n460 B.n459 163.367
R1420 B.n459 B.n458 163.367
R1421 B.n458 B.n59 163.367
R1422 B.n454 B.n59 163.367
R1423 B.n454 B.n453 163.367
R1424 B.n453 B.n452 163.367
R1425 B.n452 B.n61 163.367
R1426 B.n448 B.n61 163.367
R1427 B.n448 B.n447 163.367
R1428 B.n447 B.n446 163.367
R1429 B.n446 B.n63 163.367
R1430 B.n442 B.n63 163.367
R1431 B.n442 B.n441 163.367
R1432 B.n441 B.n440 163.367
R1433 B.n440 B.n65 163.367
R1434 B.n436 B.n65 163.367
R1435 B.n436 B.n435 163.367
R1436 B.n435 B.n434 163.367
R1437 B.n574 B.n573 163.367
R1438 B.n574 B.n15 163.367
R1439 B.n578 B.n15 163.367
R1440 B.n579 B.n578 163.367
R1441 B.n580 B.n579 163.367
R1442 B.n580 B.n13 163.367
R1443 B.n584 B.n13 163.367
R1444 B.n585 B.n584 163.367
R1445 B.n586 B.n585 163.367
R1446 B.n586 B.n11 163.367
R1447 B.n590 B.n11 163.367
R1448 B.n591 B.n590 163.367
R1449 B.n592 B.n591 163.367
R1450 B.n592 B.n9 163.367
R1451 B.n596 B.n9 163.367
R1452 B.n597 B.n596 163.367
R1453 B.n598 B.n597 163.367
R1454 B.n598 B.n7 163.367
R1455 B.n602 B.n7 163.367
R1456 B.n603 B.n602 163.367
R1457 B.n604 B.n603 163.367
R1458 B.n604 B.n5 163.367
R1459 B.n608 B.n5 163.367
R1460 B.n609 B.n608 163.367
R1461 B.n610 B.n609 163.367
R1462 B.n610 B.n3 163.367
R1463 B.n614 B.n3 163.367
R1464 B.n615 B.n614 163.367
R1465 B.n160 B.n2 163.367
R1466 B.n161 B.n160 163.367
R1467 B.n162 B.n161 163.367
R1468 B.n162 B.n157 163.367
R1469 B.n166 B.n157 163.367
R1470 B.n167 B.n166 163.367
R1471 B.n168 B.n167 163.367
R1472 B.n168 B.n155 163.367
R1473 B.n172 B.n155 163.367
R1474 B.n173 B.n172 163.367
R1475 B.n174 B.n173 163.367
R1476 B.n174 B.n153 163.367
R1477 B.n178 B.n153 163.367
R1478 B.n179 B.n178 163.367
R1479 B.n180 B.n179 163.367
R1480 B.n180 B.n151 163.367
R1481 B.n184 B.n151 163.367
R1482 B.n185 B.n184 163.367
R1483 B.n186 B.n185 163.367
R1484 B.n186 B.n149 163.367
R1485 B.n190 B.n149 163.367
R1486 B.n191 B.n190 163.367
R1487 B.n192 B.n191 163.367
R1488 B.n192 B.n147 163.367
R1489 B.n196 B.n147 163.367
R1490 B.n197 B.n196 163.367
R1491 B.n198 B.n197 163.367
R1492 B.n198 B.n145 163.367
R1493 B.n263 B.n262 59.5399
R1494 B.n281 B.n119 59.5399
R1495 B.n46 B.n45 59.5399
R1496 B.n510 B.n39 59.5399
R1497 B.n571 B.n16 34.8103
R1498 B.n433 B.n432 34.8103
R1499 B.n201 B.n200 34.8103
R1500 B.n343 B.n342 34.8103
R1501 B.n262 B.n261 28.3157
R1502 B.n119 B.n118 28.3157
R1503 B.n45 B.n44 28.3157
R1504 B.n39 B.n38 28.3157
R1505 B B.n617 18.0485
R1506 B.n575 B.n16 10.6151
R1507 B.n576 B.n575 10.6151
R1508 B.n577 B.n576 10.6151
R1509 B.n577 B.n14 10.6151
R1510 B.n581 B.n14 10.6151
R1511 B.n582 B.n581 10.6151
R1512 B.n583 B.n582 10.6151
R1513 B.n583 B.n12 10.6151
R1514 B.n587 B.n12 10.6151
R1515 B.n588 B.n587 10.6151
R1516 B.n589 B.n588 10.6151
R1517 B.n589 B.n10 10.6151
R1518 B.n593 B.n10 10.6151
R1519 B.n594 B.n593 10.6151
R1520 B.n595 B.n594 10.6151
R1521 B.n595 B.n8 10.6151
R1522 B.n599 B.n8 10.6151
R1523 B.n600 B.n599 10.6151
R1524 B.n601 B.n600 10.6151
R1525 B.n601 B.n6 10.6151
R1526 B.n605 B.n6 10.6151
R1527 B.n606 B.n605 10.6151
R1528 B.n607 B.n606 10.6151
R1529 B.n607 B.n4 10.6151
R1530 B.n611 B.n4 10.6151
R1531 B.n612 B.n611 10.6151
R1532 B.n613 B.n612 10.6151
R1533 B.n613 B.n0 10.6151
R1534 B.n571 B.n570 10.6151
R1535 B.n570 B.n569 10.6151
R1536 B.n569 B.n18 10.6151
R1537 B.n565 B.n18 10.6151
R1538 B.n565 B.n564 10.6151
R1539 B.n564 B.n563 10.6151
R1540 B.n563 B.n20 10.6151
R1541 B.n559 B.n20 10.6151
R1542 B.n559 B.n558 10.6151
R1543 B.n558 B.n557 10.6151
R1544 B.n557 B.n22 10.6151
R1545 B.n553 B.n22 10.6151
R1546 B.n553 B.n552 10.6151
R1547 B.n552 B.n551 10.6151
R1548 B.n551 B.n24 10.6151
R1549 B.n547 B.n24 10.6151
R1550 B.n547 B.n546 10.6151
R1551 B.n546 B.n545 10.6151
R1552 B.n545 B.n26 10.6151
R1553 B.n541 B.n26 10.6151
R1554 B.n541 B.n540 10.6151
R1555 B.n540 B.n539 10.6151
R1556 B.n539 B.n28 10.6151
R1557 B.n535 B.n28 10.6151
R1558 B.n535 B.n534 10.6151
R1559 B.n534 B.n533 10.6151
R1560 B.n533 B.n30 10.6151
R1561 B.n529 B.n30 10.6151
R1562 B.n529 B.n528 10.6151
R1563 B.n528 B.n527 10.6151
R1564 B.n527 B.n32 10.6151
R1565 B.n523 B.n32 10.6151
R1566 B.n523 B.n522 10.6151
R1567 B.n522 B.n521 10.6151
R1568 B.n521 B.n34 10.6151
R1569 B.n517 B.n34 10.6151
R1570 B.n517 B.n516 10.6151
R1571 B.n516 B.n515 10.6151
R1572 B.n515 B.n36 10.6151
R1573 B.n511 B.n36 10.6151
R1574 B.n509 B.n508 10.6151
R1575 B.n508 B.n40 10.6151
R1576 B.n504 B.n40 10.6151
R1577 B.n504 B.n503 10.6151
R1578 B.n503 B.n502 10.6151
R1579 B.n502 B.n42 10.6151
R1580 B.n498 B.n42 10.6151
R1581 B.n498 B.n497 10.6151
R1582 B.n497 B.n496 10.6151
R1583 B.n493 B.n492 10.6151
R1584 B.n492 B.n491 10.6151
R1585 B.n491 B.n48 10.6151
R1586 B.n487 B.n48 10.6151
R1587 B.n487 B.n486 10.6151
R1588 B.n486 B.n485 10.6151
R1589 B.n485 B.n50 10.6151
R1590 B.n481 B.n50 10.6151
R1591 B.n481 B.n480 10.6151
R1592 B.n480 B.n479 10.6151
R1593 B.n479 B.n52 10.6151
R1594 B.n475 B.n52 10.6151
R1595 B.n475 B.n474 10.6151
R1596 B.n474 B.n473 10.6151
R1597 B.n473 B.n54 10.6151
R1598 B.n469 B.n54 10.6151
R1599 B.n469 B.n468 10.6151
R1600 B.n468 B.n467 10.6151
R1601 B.n467 B.n56 10.6151
R1602 B.n463 B.n56 10.6151
R1603 B.n463 B.n462 10.6151
R1604 B.n462 B.n461 10.6151
R1605 B.n461 B.n58 10.6151
R1606 B.n457 B.n58 10.6151
R1607 B.n457 B.n456 10.6151
R1608 B.n456 B.n455 10.6151
R1609 B.n455 B.n60 10.6151
R1610 B.n451 B.n60 10.6151
R1611 B.n451 B.n450 10.6151
R1612 B.n450 B.n449 10.6151
R1613 B.n449 B.n62 10.6151
R1614 B.n445 B.n62 10.6151
R1615 B.n445 B.n444 10.6151
R1616 B.n444 B.n443 10.6151
R1617 B.n443 B.n64 10.6151
R1618 B.n439 B.n64 10.6151
R1619 B.n439 B.n438 10.6151
R1620 B.n438 B.n437 10.6151
R1621 B.n437 B.n66 10.6151
R1622 B.n433 B.n66 10.6151
R1623 B.n432 B.n431 10.6151
R1624 B.n431 B.n68 10.6151
R1625 B.n427 B.n68 10.6151
R1626 B.n427 B.n426 10.6151
R1627 B.n426 B.n425 10.6151
R1628 B.n425 B.n70 10.6151
R1629 B.n421 B.n70 10.6151
R1630 B.n421 B.n420 10.6151
R1631 B.n420 B.n419 10.6151
R1632 B.n419 B.n72 10.6151
R1633 B.n415 B.n72 10.6151
R1634 B.n415 B.n414 10.6151
R1635 B.n414 B.n413 10.6151
R1636 B.n413 B.n74 10.6151
R1637 B.n409 B.n74 10.6151
R1638 B.n409 B.n408 10.6151
R1639 B.n408 B.n407 10.6151
R1640 B.n407 B.n76 10.6151
R1641 B.n403 B.n76 10.6151
R1642 B.n403 B.n402 10.6151
R1643 B.n402 B.n401 10.6151
R1644 B.n401 B.n78 10.6151
R1645 B.n397 B.n78 10.6151
R1646 B.n397 B.n396 10.6151
R1647 B.n396 B.n395 10.6151
R1648 B.n395 B.n80 10.6151
R1649 B.n391 B.n80 10.6151
R1650 B.n391 B.n390 10.6151
R1651 B.n390 B.n389 10.6151
R1652 B.n389 B.n82 10.6151
R1653 B.n385 B.n82 10.6151
R1654 B.n385 B.n384 10.6151
R1655 B.n384 B.n383 10.6151
R1656 B.n383 B.n84 10.6151
R1657 B.n379 B.n84 10.6151
R1658 B.n379 B.n378 10.6151
R1659 B.n378 B.n377 10.6151
R1660 B.n377 B.n86 10.6151
R1661 B.n373 B.n86 10.6151
R1662 B.n373 B.n372 10.6151
R1663 B.n372 B.n371 10.6151
R1664 B.n371 B.n88 10.6151
R1665 B.n367 B.n88 10.6151
R1666 B.n367 B.n366 10.6151
R1667 B.n366 B.n365 10.6151
R1668 B.n365 B.n90 10.6151
R1669 B.n361 B.n90 10.6151
R1670 B.n361 B.n360 10.6151
R1671 B.n360 B.n359 10.6151
R1672 B.n359 B.n92 10.6151
R1673 B.n355 B.n92 10.6151
R1674 B.n355 B.n354 10.6151
R1675 B.n354 B.n353 10.6151
R1676 B.n353 B.n94 10.6151
R1677 B.n349 B.n94 10.6151
R1678 B.n349 B.n348 10.6151
R1679 B.n348 B.n347 10.6151
R1680 B.n347 B.n96 10.6151
R1681 B.n343 B.n96 10.6151
R1682 B.n159 B.n1 10.6151
R1683 B.n159 B.n158 10.6151
R1684 B.n163 B.n158 10.6151
R1685 B.n164 B.n163 10.6151
R1686 B.n165 B.n164 10.6151
R1687 B.n165 B.n156 10.6151
R1688 B.n169 B.n156 10.6151
R1689 B.n170 B.n169 10.6151
R1690 B.n171 B.n170 10.6151
R1691 B.n171 B.n154 10.6151
R1692 B.n175 B.n154 10.6151
R1693 B.n176 B.n175 10.6151
R1694 B.n177 B.n176 10.6151
R1695 B.n177 B.n152 10.6151
R1696 B.n181 B.n152 10.6151
R1697 B.n182 B.n181 10.6151
R1698 B.n183 B.n182 10.6151
R1699 B.n183 B.n150 10.6151
R1700 B.n187 B.n150 10.6151
R1701 B.n188 B.n187 10.6151
R1702 B.n189 B.n188 10.6151
R1703 B.n189 B.n148 10.6151
R1704 B.n193 B.n148 10.6151
R1705 B.n194 B.n193 10.6151
R1706 B.n195 B.n194 10.6151
R1707 B.n195 B.n146 10.6151
R1708 B.n199 B.n146 10.6151
R1709 B.n200 B.n199 10.6151
R1710 B.n201 B.n144 10.6151
R1711 B.n205 B.n144 10.6151
R1712 B.n206 B.n205 10.6151
R1713 B.n207 B.n206 10.6151
R1714 B.n207 B.n142 10.6151
R1715 B.n211 B.n142 10.6151
R1716 B.n212 B.n211 10.6151
R1717 B.n213 B.n212 10.6151
R1718 B.n213 B.n140 10.6151
R1719 B.n217 B.n140 10.6151
R1720 B.n218 B.n217 10.6151
R1721 B.n219 B.n218 10.6151
R1722 B.n219 B.n138 10.6151
R1723 B.n223 B.n138 10.6151
R1724 B.n224 B.n223 10.6151
R1725 B.n225 B.n224 10.6151
R1726 B.n225 B.n136 10.6151
R1727 B.n229 B.n136 10.6151
R1728 B.n230 B.n229 10.6151
R1729 B.n231 B.n230 10.6151
R1730 B.n231 B.n134 10.6151
R1731 B.n235 B.n134 10.6151
R1732 B.n236 B.n235 10.6151
R1733 B.n237 B.n236 10.6151
R1734 B.n237 B.n132 10.6151
R1735 B.n241 B.n132 10.6151
R1736 B.n242 B.n241 10.6151
R1737 B.n243 B.n242 10.6151
R1738 B.n243 B.n130 10.6151
R1739 B.n247 B.n130 10.6151
R1740 B.n248 B.n247 10.6151
R1741 B.n249 B.n248 10.6151
R1742 B.n249 B.n128 10.6151
R1743 B.n253 B.n128 10.6151
R1744 B.n254 B.n253 10.6151
R1745 B.n255 B.n254 10.6151
R1746 B.n255 B.n126 10.6151
R1747 B.n259 B.n126 10.6151
R1748 B.n260 B.n259 10.6151
R1749 B.n264 B.n260 10.6151
R1750 B.n268 B.n124 10.6151
R1751 B.n269 B.n268 10.6151
R1752 B.n270 B.n269 10.6151
R1753 B.n270 B.n122 10.6151
R1754 B.n274 B.n122 10.6151
R1755 B.n275 B.n274 10.6151
R1756 B.n276 B.n275 10.6151
R1757 B.n276 B.n120 10.6151
R1758 B.n280 B.n120 10.6151
R1759 B.n283 B.n282 10.6151
R1760 B.n283 B.n116 10.6151
R1761 B.n287 B.n116 10.6151
R1762 B.n288 B.n287 10.6151
R1763 B.n289 B.n288 10.6151
R1764 B.n289 B.n114 10.6151
R1765 B.n293 B.n114 10.6151
R1766 B.n294 B.n293 10.6151
R1767 B.n295 B.n294 10.6151
R1768 B.n295 B.n112 10.6151
R1769 B.n299 B.n112 10.6151
R1770 B.n300 B.n299 10.6151
R1771 B.n301 B.n300 10.6151
R1772 B.n301 B.n110 10.6151
R1773 B.n305 B.n110 10.6151
R1774 B.n306 B.n305 10.6151
R1775 B.n307 B.n306 10.6151
R1776 B.n307 B.n108 10.6151
R1777 B.n311 B.n108 10.6151
R1778 B.n312 B.n311 10.6151
R1779 B.n313 B.n312 10.6151
R1780 B.n313 B.n106 10.6151
R1781 B.n317 B.n106 10.6151
R1782 B.n318 B.n317 10.6151
R1783 B.n319 B.n318 10.6151
R1784 B.n319 B.n104 10.6151
R1785 B.n323 B.n104 10.6151
R1786 B.n324 B.n323 10.6151
R1787 B.n325 B.n324 10.6151
R1788 B.n325 B.n102 10.6151
R1789 B.n329 B.n102 10.6151
R1790 B.n330 B.n329 10.6151
R1791 B.n331 B.n330 10.6151
R1792 B.n331 B.n100 10.6151
R1793 B.n335 B.n100 10.6151
R1794 B.n336 B.n335 10.6151
R1795 B.n337 B.n336 10.6151
R1796 B.n337 B.n98 10.6151
R1797 B.n341 B.n98 10.6151
R1798 B.n342 B.n341 10.6151
R1799 B.n511 B.n510 9.36635
R1800 B.n493 B.n46 9.36635
R1801 B.n264 B.n263 9.36635
R1802 B.n282 B.n281 9.36635
R1803 B.n617 B.n0 8.11757
R1804 B.n617 B.n1 8.11757
R1805 B.n510 B.n509 1.24928
R1806 B.n496 B.n46 1.24928
R1807 B.n263 B.n124 1.24928
R1808 B.n281 B.n280 1.24928
R1809 VP.n7 VP.t0 311.981
R1810 VP.n17 VP.t5 288.988
R1811 VP.n29 VP.t6 288.988
R1812 VP.n15 VP.t1 288.988
R1813 VP.n22 VP.t4 254.011
R1814 VP.n1 VP.t2 254.011
R1815 VP.n5 VP.t3 254.011
R1816 VP.n8 VP.t7 254.011
R1817 VP.n9 VP.n6 161.3
R1818 VP.n11 VP.n10 161.3
R1819 VP.n13 VP.n12 161.3
R1820 VP.n14 VP.n4 161.3
R1821 VP.n28 VP.n0 161.3
R1822 VP.n27 VP.n26 161.3
R1823 VP.n25 VP.n24 161.3
R1824 VP.n23 VP.n2 161.3
R1825 VP.n21 VP.n20 161.3
R1826 VP.n19 VP.n3 161.3
R1827 VP.n16 VP.n15 80.6037
R1828 VP.n30 VP.n29 80.6037
R1829 VP.n18 VP.n17 80.6037
R1830 VP.n24 VP.n23 56.5193
R1831 VP.n10 VP.n9 56.5193
R1832 VP.n17 VP.n3 50.4025
R1833 VP.n29 VP.n28 50.4025
R1834 VP.n15 VP.n14 50.4025
R1835 VP.n18 VP.n16 44.1529
R1836 VP.n8 VP.n7 33.6057
R1837 VP.n7 VP.n6 28.1515
R1838 VP.n21 VP.n3 24.4675
R1839 VP.n28 VP.n27 24.4675
R1840 VP.n14 VP.n13 24.4675
R1841 VP.n23 VP.n22 23.4888
R1842 VP.n24 VP.n1 23.4888
R1843 VP.n10 VP.n5 23.4888
R1844 VP.n9 VP.n8 23.4888
R1845 VP.n22 VP.n21 0.97918
R1846 VP.n27 VP.n1 0.97918
R1847 VP.n13 VP.n5 0.97918
R1848 VP.n16 VP.n4 0.285035
R1849 VP.n19 VP.n18 0.285035
R1850 VP.n30 VP.n0 0.285035
R1851 VP.n11 VP.n6 0.189894
R1852 VP.n12 VP.n11 0.189894
R1853 VP.n12 VP.n4 0.189894
R1854 VP.n20 VP.n19 0.189894
R1855 VP.n20 VP.n2 0.189894
R1856 VP.n25 VP.n2 0.189894
R1857 VP.n26 VP.n25 0.189894
R1858 VP.n26 VP.n0 0.189894
R1859 VP VP.n30 0.146778
R1860 VDD1 VDD1.n0 77.0125
R1861 VDD1.n3 VDD1.n2 76.8988
R1862 VDD1.n3 VDD1.n1 76.8988
R1863 VDD1.n5 VDD1.n4 76.3239
R1864 VDD1.n5 VDD1.n3 40.2293
R1865 VDD1.n4 VDD1.t4 2.72972
R1866 VDD1.n4 VDD1.t6 2.72972
R1867 VDD1.n0 VDD1.t7 2.72972
R1868 VDD1.n0 VDD1.t0 2.72972
R1869 VDD1.n2 VDD1.t5 2.72972
R1870 VDD1.n2 VDD1.t1 2.72972
R1871 VDD1.n1 VDD1.t2 2.72972
R1872 VDD1.n1 VDD1.t3 2.72972
R1873 VDD1 VDD1.n5 0.571621
C0 VP VDD2 0.363304f
C1 VTAIL VN 6.71712f
C2 VDD2 w_n2430_n3350# 1.51308f
C3 VP B 1.39508f
C4 B w_n2430_n3350# 7.8401f
C5 VP VDD1 7.00523f
C6 VDD1 w_n2430_n3350# 1.46021f
C7 VDD2 VN 6.79171f
C8 B VN 0.881358f
C9 VDD2 VTAIL 9.16424f
C10 VP w_n2430_n3350# 4.83465f
C11 VDD1 VN 0.149127f
C12 B VTAIL 4.1361f
C13 VDD1 VTAIL 9.119679f
C14 VP VN 5.8459f
C15 w_n2430_n3350# VN 4.52352f
C16 VP VTAIL 6.73123f
C17 VDD2 B 1.24898f
C18 w_n2430_n3350# VTAIL 4.1394f
C19 VDD2 VDD1 1.04164f
C20 B VDD1 1.19901f
C21 VDD2 VSUBS 1.38746f
C22 VDD1 VSUBS 1.767789f
C23 VTAIL VSUBS 1.036568f
C24 VN VSUBS 5.03126f
C25 VP VSUBS 2.100402f
C26 B VSUBS 3.356914f
C27 w_n2430_n3350# VSUBS 0.100223p
C28 VDD1.t7 VSUBS 0.24155f
C29 VDD1.t0 VSUBS 0.24155f
C30 VDD1.n0 VSUBS 1.90869f
C31 VDD1.t2 VSUBS 0.24155f
C32 VDD1.t3 VSUBS 0.24155f
C33 VDD1.n1 VSUBS 1.90769f
C34 VDD1.t5 VSUBS 0.24155f
C35 VDD1.t1 VSUBS 0.24155f
C36 VDD1.n2 VSUBS 1.90769f
C37 VDD1.n3 VSUBS 3.03264f
C38 VDD1.t4 VSUBS 0.24155f
C39 VDD1.t6 VSUBS 0.24155f
C40 VDD1.n4 VSUBS 1.90304f
C41 VDD1.n5 VSUBS 2.77747f
C42 VP.n0 VSUBS 0.060217f
C43 VP.t2 VSUBS 1.65441f
C44 VP.n1 VSUBS 0.608874f
C45 VP.n2 VSUBS 0.045127f
C46 VP.t4 VSUBS 1.65441f
C47 VP.n3 VSUBS 0.05867f
C48 VP.n4 VSUBS 0.060217f
C49 VP.t1 VSUBS 1.73254f
C50 VP.t3 VSUBS 1.65441f
C51 VP.n5 VSUBS 0.608874f
C52 VP.n6 VSUBS 0.237578f
C53 VP.t7 VSUBS 1.65441f
C54 VP.t0 VSUBS 1.78414f
C55 VP.n7 VSUBS 0.669093f
C56 VP.n8 VSUBS 0.682119f
C57 VP.n9 VSUBS 0.064217f
C58 VP.n10 VSUBS 0.064217f
C59 VP.n11 VSUBS 0.045127f
C60 VP.n12 VSUBS 0.045127f
C61 VP.n13 VSUBS 0.044243f
C62 VP.n14 VSUBS 0.05867f
C63 VP.n15 VSUBS 0.688777f
C64 VP.n16 VSUBS 2.03786f
C65 VP.t5 VSUBS 1.73254f
C66 VP.n17 VSUBS 0.688777f
C67 VP.n18 VSUBS 2.0746f
C68 VP.n19 VSUBS 0.060217f
C69 VP.n20 VSUBS 0.045127f
C70 VP.n21 VSUBS 0.044243f
C71 VP.n22 VSUBS 0.608874f
C72 VP.n23 VSUBS 0.064217f
C73 VP.n24 VSUBS 0.064217f
C74 VP.n25 VSUBS 0.045127f
C75 VP.n26 VSUBS 0.045127f
C76 VP.n27 VSUBS 0.044243f
C77 VP.n28 VSUBS 0.05867f
C78 VP.t6 VSUBS 1.73254f
C79 VP.n29 VSUBS 0.688777f
C80 VP.n30 VSUBS 0.042264f
C81 B.n0 VSUBS 0.006779f
C82 B.n1 VSUBS 0.006779f
C83 B.n2 VSUBS 0.010026f
C84 B.n3 VSUBS 0.007683f
C85 B.n4 VSUBS 0.007683f
C86 B.n5 VSUBS 0.007683f
C87 B.n6 VSUBS 0.007683f
C88 B.n7 VSUBS 0.007683f
C89 B.n8 VSUBS 0.007683f
C90 B.n9 VSUBS 0.007683f
C91 B.n10 VSUBS 0.007683f
C92 B.n11 VSUBS 0.007683f
C93 B.n12 VSUBS 0.007683f
C94 B.n13 VSUBS 0.007683f
C95 B.n14 VSUBS 0.007683f
C96 B.n15 VSUBS 0.007683f
C97 B.n16 VSUBS 0.018391f
C98 B.n17 VSUBS 0.007683f
C99 B.n18 VSUBS 0.007683f
C100 B.n19 VSUBS 0.007683f
C101 B.n20 VSUBS 0.007683f
C102 B.n21 VSUBS 0.007683f
C103 B.n22 VSUBS 0.007683f
C104 B.n23 VSUBS 0.007683f
C105 B.n24 VSUBS 0.007683f
C106 B.n25 VSUBS 0.007683f
C107 B.n26 VSUBS 0.007683f
C108 B.n27 VSUBS 0.007683f
C109 B.n28 VSUBS 0.007683f
C110 B.n29 VSUBS 0.007683f
C111 B.n30 VSUBS 0.007683f
C112 B.n31 VSUBS 0.007683f
C113 B.n32 VSUBS 0.007683f
C114 B.n33 VSUBS 0.007683f
C115 B.n34 VSUBS 0.007683f
C116 B.n35 VSUBS 0.007683f
C117 B.n36 VSUBS 0.007683f
C118 B.n37 VSUBS 0.007683f
C119 B.t4 VSUBS 0.229125f
C120 B.t5 VSUBS 0.247269f
C121 B.t3 VSUBS 0.632085f
C122 B.n38 VSUBS 0.368436f
C123 B.n39 VSUBS 0.268621f
C124 B.n40 VSUBS 0.007683f
C125 B.n41 VSUBS 0.007683f
C126 B.n42 VSUBS 0.007683f
C127 B.n43 VSUBS 0.007683f
C128 B.t10 VSUBS 0.229128f
C129 B.t11 VSUBS 0.247272f
C130 B.t9 VSUBS 0.632085f
C131 B.n44 VSUBS 0.368433f
C132 B.n45 VSUBS 0.268618f
C133 B.n46 VSUBS 0.0178f
C134 B.n47 VSUBS 0.007683f
C135 B.n48 VSUBS 0.007683f
C136 B.n49 VSUBS 0.007683f
C137 B.n50 VSUBS 0.007683f
C138 B.n51 VSUBS 0.007683f
C139 B.n52 VSUBS 0.007683f
C140 B.n53 VSUBS 0.007683f
C141 B.n54 VSUBS 0.007683f
C142 B.n55 VSUBS 0.007683f
C143 B.n56 VSUBS 0.007683f
C144 B.n57 VSUBS 0.007683f
C145 B.n58 VSUBS 0.007683f
C146 B.n59 VSUBS 0.007683f
C147 B.n60 VSUBS 0.007683f
C148 B.n61 VSUBS 0.007683f
C149 B.n62 VSUBS 0.007683f
C150 B.n63 VSUBS 0.007683f
C151 B.n64 VSUBS 0.007683f
C152 B.n65 VSUBS 0.007683f
C153 B.n66 VSUBS 0.007683f
C154 B.n67 VSUBS 0.018391f
C155 B.n68 VSUBS 0.007683f
C156 B.n69 VSUBS 0.007683f
C157 B.n70 VSUBS 0.007683f
C158 B.n71 VSUBS 0.007683f
C159 B.n72 VSUBS 0.007683f
C160 B.n73 VSUBS 0.007683f
C161 B.n74 VSUBS 0.007683f
C162 B.n75 VSUBS 0.007683f
C163 B.n76 VSUBS 0.007683f
C164 B.n77 VSUBS 0.007683f
C165 B.n78 VSUBS 0.007683f
C166 B.n79 VSUBS 0.007683f
C167 B.n80 VSUBS 0.007683f
C168 B.n81 VSUBS 0.007683f
C169 B.n82 VSUBS 0.007683f
C170 B.n83 VSUBS 0.007683f
C171 B.n84 VSUBS 0.007683f
C172 B.n85 VSUBS 0.007683f
C173 B.n86 VSUBS 0.007683f
C174 B.n87 VSUBS 0.007683f
C175 B.n88 VSUBS 0.007683f
C176 B.n89 VSUBS 0.007683f
C177 B.n90 VSUBS 0.007683f
C178 B.n91 VSUBS 0.007683f
C179 B.n92 VSUBS 0.007683f
C180 B.n93 VSUBS 0.007683f
C181 B.n94 VSUBS 0.007683f
C182 B.n95 VSUBS 0.007683f
C183 B.n96 VSUBS 0.007683f
C184 B.n97 VSUBS 0.019118f
C185 B.n98 VSUBS 0.007683f
C186 B.n99 VSUBS 0.007683f
C187 B.n100 VSUBS 0.007683f
C188 B.n101 VSUBS 0.007683f
C189 B.n102 VSUBS 0.007683f
C190 B.n103 VSUBS 0.007683f
C191 B.n104 VSUBS 0.007683f
C192 B.n105 VSUBS 0.007683f
C193 B.n106 VSUBS 0.007683f
C194 B.n107 VSUBS 0.007683f
C195 B.n108 VSUBS 0.007683f
C196 B.n109 VSUBS 0.007683f
C197 B.n110 VSUBS 0.007683f
C198 B.n111 VSUBS 0.007683f
C199 B.n112 VSUBS 0.007683f
C200 B.n113 VSUBS 0.007683f
C201 B.n114 VSUBS 0.007683f
C202 B.n115 VSUBS 0.007683f
C203 B.n116 VSUBS 0.007683f
C204 B.n117 VSUBS 0.007683f
C205 B.t2 VSUBS 0.229128f
C206 B.t1 VSUBS 0.247272f
C207 B.t0 VSUBS 0.632085f
C208 B.n118 VSUBS 0.368433f
C209 B.n119 VSUBS 0.268618f
C210 B.n120 VSUBS 0.007683f
C211 B.n121 VSUBS 0.007683f
C212 B.n122 VSUBS 0.007683f
C213 B.n123 VSUBS 0.007683f
C214 B.n124 VSUBS 0.004293f
C215 B.n125 VSUBS 0.007683f
C216 B.n126 VSUBS 0.007683f
C217 B.n127 VSUBS 0.007683f
C218 B.n128 VSUBS 0.007683f
C219 B.n129 VSUBS 0.007683f
C220 B.n130 VSUBS 0.007683f
C221 B.n131 VSUBS 0.007683f
C222 B.n132 VSUBS 0.007683f
C223 B.n133 VSUBS 0.007683f
C224 B.n134 VSUBS 0.007683f
C225 B.n135 VSUBS 0.007683f
C226 B.n136 VSUBS 0.007683f
C227 B.n137 VSUBS 0.007683f
C228 B.n138 VSUBS 0.007683f
C229 B.n139 VSUBS 0.007683f
C230 B.n140 VSUBS 0.007683f
C231 B.n141 VSUBS 0.007683f
C232 B.n142 VSUBS 0.007683f
C233 B.n143 VSUBS 0.007683f
C234 B.n144 VSUBS 0.007683f
C235 B.n145 VSUBS 0.018391f
C236 B.n146 VSUBS 0.007683f
C237 B.n147 VSUBS 0.007683f
C238 B.n148 VSUBS 0.007683f
C239 B.n149 VSUBS 0.007683f
C240 B.n150 VSUBS 0.007683f
C241 B.n151 VSUBS 0.007683f
C242 B.n152 VSUBS 0.007683f
C243 B.n153 VSUBS 0.007683f
C244 B.n154 VSUBS 0.007683f
C245 B.n155 VSUBS 0.007683f
C246 B.n156 VSUBS 0.007683f
C247 B.n157 VSUBS 0.007683f
C248 B.n158 VSUBS 0.007683f
C249 B.n159 VSUBS 0.007683f
C250 B.n160 VSUBS 0.007683f
C251 B.n161 VSUBS 0.007683f
C252 B.n162 VSUBS 0.007683f
C253 B.n163 VSUBS 0.007683f
C254 B.n164 VSUBS 0.007683f
C255 B.n165 VSUBS 0.007683f
C256 B.n166 VSUBS 0.007683f
C257 B.n167 VSUBS 0.007683f
C258 B.n168 VSUBS 0.007683f
C259 B.n169 VSUBS 0.007683f
C260 B.n170 VSUBS 0.007683f
C261 B.n171 VSUBS 0.007683f
C262 B.n172 VSUBS 0.007683f
C263 B.n173 VSUBS 0.007683f
C264 B.n174 VSUBS 0.007683f
C265 B.n175 VSUBS 0.007683f
C266 B.n176 VSUBS 0.007683f
C267 B.n177 VSUBS 0.007683f
C268 B.n178 VSUBS 0.007683f
C269 B.n179 VSUBS 0.007683f
C270 B.n180 VSUBS 0.007683f
C271 B.n181 VSUBS 0.007683f
C272 B.n182 VSUBS 0.007683f
C273 B.n183 VSUBS 0.007683f
C274 B.n184 VSUBS 0.007683f
C275 B.n185 VSUBS 0.007683f
C276 B.n186 VSUBS 0.007683f
C277 B.n187 VSUBS 0.007683f
C278 B.n188 VSUBS 0.007683f
C279 B.n189 VSUBS 0.007683f
C280 B.n190 VSUBS 0.007683f
C281 B.n191 VSUBS 0.007683f
C282 B.n192 VSUBS 0.007683f
C283 B.n193 VSUBS 0.007683f
C284 B.n194 VSUBS 0.007683f
C285 B.n195 VSUBS 0.007683f
C286 B.n196 VSUBS 0.007683f
C287 B.n197 VSUBS 0.007683f
C288 B.n198 VSUBS 0.007683f
C289 B.n199 VSUBS 0.007683f
C290 B.n200 VSUBS 0.018391f
C291 B.n201 VSUBS 0.019118f
C292 B.n202 VSUBS 0.019118f
C293 B.n203 VSUBS 0.007683f
C294 B.n204 VSUBS 0.007683f
C295 B.n205 VSUBS 0.007683f
C296 B.n206 VSUBS 0.007683f
C297 B.n207 VSUBS 0.007683f
C298 B.n208 VSUBS 0.007683f
C299 B.n209 VSUBS 0.007683f
C300 B.n210 VSUBS 0.007683f
C301 B.n211 VSUBS 0.007683f
C302 B.n212 VSUBS 0.007683f
C303 B.n213 VSUBS 0.007683f
C304 B.n214 VSUBS 0.007683f
C305 B.n215 VSUBS 0.007683f
C306 B.n216 VSUBS 0.007683f
C307 B.n217 VSUBS 0.007683f
C308 B.n218 VSUBS 0.007683f
C309 B.n219 VSUBS 0.007683f
C310 B.n220 VSUBS 0.007683f
C311 B.n221 VSUBS 0.007683f
C312 B.n222 VSUBS 0.007683f
C313 B.n223 VSUBS 0.007683f
C314 B.n224 VSUBS 0.007683f
C315 B.n225 VSUBS 0.007683f
C316 B.n226 VSUBS 0.007683f
C317 B.n227 VSUBS 0.007683f
C318 B.n228 VSUBS 0.007683f
C319 B.n229 VSUBS 0.007683f
C320 B.n230 VSUBS 0.007683f
C321 B.n231 VSUBS 0.007683f
C322 B.n232 VSUBS 0.007683f
C323 B.n233 VSUBS 0.007683f
C324 B.n234 VSUBS 0.007683f
C325 B.n235 VSUBS 0.007683f
C326 B.n236 VSUBS 0.007683f
C327 B.n237 VSUBS 0.007683f
C328 B.n238 VSUBS 0.007683f
C329 B.n239 VSUBS 0.007683f
C330 B.n240 VSUBS 0.007683f
C331 B.n241 VSUBS 0.007683f
C332 B.n242 VSUBS 0.007683f
C333 B.n243 VSUBS 0.007683f
C334 B.n244 VSUBS 0.007683f
C335 B.n245 VSUBS 0.007683f
C336 B.n246 VSUBS 0.007683f
C337 B.n247 VSUBS 0.007683f
C338 B.n248 VSUBS 0.007683f
C339 B.n249 VSUBS 0.007683f
C340 B.n250 VSUBS 0.007683f
C341 B.n251 VSUBS 0.007683f
C342 B.n252 VSUBS 0.007683f
C343 B.n253 VSUBS 0.007683f
C344 B.n254 VSUBS 0.007683f
C345 B.n255 VSUBS 0.007683f
C346 B.n256 VSUBS 0.007683f
C347 B.n257 VSUBS 0.007683f
C348 B.n258 VSUBS 0.007683f
C349 B.n259 VSUBS 0.007683f
C350 B.n260 VSUBS 0.007683f
C351 B.t8 VSUBS 0.229125f
C352 B.t7 VSUBS 0.247269f
C353 B.t6 VSUBS 0.632085f
C354 B.n261 VSUBS 0.368436f
C355 B.n262 VSUBS 0.268621f
C356 B.n263 VSUBS 0.0178f
C357 B.n264 VSUBS 0.007231f
C358 B.n265 VSUBS 0.007683f
C359 B.n266 VSUBS 0.007683f
C360 B.n267 VSUBS 0.007683f
C361 B.n268 VSUBS 0.007683f
C362 B.n269 VSUBS 0.007683f
C363 B.n270 VSUBS 0.007683f
C364 B.n271 VSUBS 0.007683f
C365 B.n272 VSUBS 0.007683f
C366 B.n273 VSUBS 0.007683f
C367 B.n274 VSUBS 0.007683f
C368 B.n275 VSUBS 0.007683f
C369 B.n276 VSUBS 0.007683f
C370 B.n277 VSUBS 0.007683f
C371 B.n278 VSUBS 0.007683f
C372 B.n279 VSUBS 0.007683f
C373 B.n280 VSUBS 0.004293f
C374 B.n281 VSUBS 0.0178f
C375 B.n282 VSUBS 0.007231f
C376 B.n283 VSUBS 0.007683f
C377 B.n284 VSUBS 0.007683f
C378 B.n285 VSUBS 0.007683f
C379 B.n286 VSUBS 0.007683f
C380 B.n287 VSUBS 0.007683f
C381 B.n288 VSUBS 0.007683f
C382 B.n289 VSUBS 0.007683f
C383 B.n290 VSUBS 0.007683f
C384 B.n291 VSUBS 0.007683f
C385 B.n292 VSUBS 0.007683f
C386 B.n293 VSUBS 0.007683f
C387 B.n294 VSUBS 0.007683f
C388 B.n295 VSUBS 0.007683f
C389 B.n296 VSUBS 0.007683f
C390 B.n297 VSUBS 0.007683f
C391 B.n298 VSUBS 0.007683f
C392 B.n299 VSUBS 0.007683f
C393 B.n300 VSUBS 0.007683f
C394 B.n301 VSUBS 0.007683f
C395 B.n302 VSUBS 0.007683f
C396 B.n303 VSUBS 0.007683f
C397 B.n304 VSUBS 0.007683f
C398 B.n305 VSUBS 0.007683f
C399 B.n306 VSUBS 0.007683f
C400 B.n307 VSUBS 0.007683f
C401 B.n308 VSUBS 0.007683f
C402 B.n309 VSUBS 0.007683f
C403 B.n310 VSUBS 0.007683f
C404 B.n311 VSUBS 0.007683f
C405 B.n312 VSUBS 0.007683f
C406 B.n313 VSUBS 0.007683f
C407 B.n314 VSUBS 0.007683f
C408 B.n315 VSUBS 0.007683f
C409 B.n316 VSUBS 0.007683f
C410 B.n317 VSUBS 0.007683f
C411 B.n318 VSUBS 0.007683f
C412 B.n319 VSUBS 0.007683f
C413 B.n320 VSUBS 0.007683f
C414 B.n321 VSUBS 0.007683f
C415 B.n322 VSUBS 0.007683f
C416 B.n323 VSUBS 0.007683f
C417 B.n324 VSUBS 0.007683f
C418 B.n325 VSUBS 0.007683f
C419 B.n326 VSUBS 0.007683f
C420 B.n327 VSUBS 0.007683f
C421 B.n328 VSUBS 0.007683f
C422 B.n329 VSUBS 0.007683f
C423 B.n330 VSUBS 0.007683f
C424 B.n331 VSUBS 0.007683f
C425 B.n332 VSUBS 0.007683f
C426 B.n333 VSUBS 0.007683f
C427 B.n334 VSUBS 0.007683f
C428 B.n335 VSUBS 0.007683f
C429 B.n336 VSUBS 0.007683f
C430 B.n337 VSUBS 0.007683f
C431 B.n338 VSUBS 0.007683f
C432 B.n339 VSUBS 0.007683f
C433 B.n340 VSUBS 0.007683f
C434 B.n341 VSUBS 0.007683f
C435 B.n342 VSUBS 0.018267f
C436 B.n343 VSUBS 0.019243f
C437 B.n344 VSUBS 0.018391f
C438 B.n345 VSUBS 0.007683f
C439 B.n346 VSUBS 0.007683f
C440 B.n347 VSUBS 0.007683f
C441 B.n348 VSUBS 0.007683f
C442 B.n349 VSUBS 0.007683f
C443 B.n350 VSUBS 0.007683f
C444 B.n351 VSUBS 0.007683f
C445 B.n352 VSUBS 0.007683f
C446 B.n353 VSUBS 0.007683f
C447 B.n354 VSUBS 0.007683f
C448 B.n355 VSUBS 0.007683f
C449 B.n356 VSUBS 0.007683f
C450 B.n357 VSUBS 0.007683f
C451 B.n358 VSUBS 0.007683f
C452 B.n359 VSUBS 0.007683f
C453 B.n360 VSUBS 0.007683f
C454 B.n361 VSUBS 0.007683f
C455 B.n362 VSUBS 0.007683f
C456 B.n363 VSUBS 0.007683f
C457 B.n364 VSUBS 0.007683f
C458 B.n365 VSUBS 0.007683f
C459 B.n366 VSUBS 0.007683f
C460 B.n367 VSUBS 0.007683f
C461 B.n368 VSUBS 0.007683f
C462 B.n369 VSUBS 0.007683f
C463 B.n370 VSUBS 0.007683f
C464 B.n371 VSUBS 0.007683f
C465 B.n372 VSUBS 0.007683f
C466 B.n373 VSUBS 0.007683f
C467 B.n374 VSUBS 0.007683f
C468 B.n375 VSUBS 0.007683f
C469 B.n376 VSUBS 0.007683f
C470 B.n377 VSUBS 0.007683f
C471 B.n378 VSUBS 0.007683f
C472 B.n379 VSUBS 0.007683f
C473 B.n380 VSUBS 0.007683f
C474 B.n381 VSUBS 0.007683f
C475 B.n382 VSUBS 0.007683f
C476 B.n383 VSUBS 0.007683f
C477 B.n384 VSUBS 0.007683f
C478 B.n385 VSUBS 0.007683f
C479 B.n386 VSUBS 0.007683f
C480 B.n387 VSUBS 0.007683f
C481 B.n388 VSUBS 0.007683f
C482 B.n389 VSUBS 0.007683f
C483 B.n390 VSUBS 0.007683f
C484 B.n391 VSUBS 0.007683f
C485 B.n392 VSUBS 0.007683f
C486 B.n393 VSUBS 0.007683f
C487 B.n394 VSUBS 0.007683f
C488 B.n395 VSUBS 0.007683f
C489 B.n396 VSUBS 0.007683f
C490 B.n397 VSUBS 0.007683f
C491 B.n398 VSUBS 0.007683f
C492 B.n399 VSUBS 0.007683f
C493 B.n400 VSUBS 0.007683f
C494 B.n401 VSUBS 0.007683f
C495 B.n402 VSUBS 0.007683f
C496 B.n403 VSUBS 0.007683f
C497 B.n404 VSUBS 0.007683f
C498 B.n405 VSUBS 0.007683f
C499 B.n406 VSUBS 0.007683f
C500 B.n407 VSUBS 0.007683f
C501 B.n408 VSUBS 0.007683f
C502 B.n409 VSUBS 0.007683f
C503 B.n410 VSUBS 0.007683f
C504 B.n411 VSUBS 0.007683f
C505 B.n412 VSUBS 0.007683f
C506 B.n413 VSUBS 0.007683f
C507 B.n414 VSUBS 0.007683f
C508 B.n415 VSUBS 0.007683f
C509 B.n416 VSUBS 0.007683f
C510 B.n417 VSUBS 0.007683f
C511 B.n418 VSUBS 0.007683f
C512 B.n419 VSUBS 0.007683f
C513 B.n420 VSUBS 0.007683f
C514 B.n421 VSUBS 0.007683f
C515 B.n422 VSUBS 0.007683f
C516 B.n423 VSUBS 0.007683f
C517 B.n424 VSUBS 0.007683f
C518 B.n425 VSUBS 0.007683f
C519 B.n426 VSUBS 0.007683f
C520 B.n427 VSUBS 0.007683f
C521 B.n428 VSUBS 0.007683f
C522 B.n429 VSUBS 0.007683f
C523 B.n430 VSUBS 0.007683f
C524 B.n431 VSUBS 0.007683f
C525 B.n432 VSUBS 0.018391f
C526 B.n433 VSUBS 0.019118f
C527 B.n434 VSUBS 0.019118f
C528 B.n435 VSUBS 0.007683f
C529 B.n436 VSUBS 0.007683f
C530 B.n437 VSUBS 0.007683f
C531 B.n438 VSUBS 0.007683f
C532 B.n439 VSUBS 0.007683f
C533 B.n440 VSUBS 0.007683f
C534 B.n441 VSUBS 0.007683f
C535 B.n442 VSUBS 0.007683f
C536 B.n443 VSUBS 0.007683f
C537 B.n444 VSUBS 0.007683f
C538 B.n445 VSUBS 0.007683f
C539 B.n446 VSUBS 0.007683f
C540 B.n447 VSUBS 0.007683f
C541 B.n448 VSUBS 0.007683f
C542 B.n449 VSUBS 0.007683f
C543 B.n450 VSUBS 0.007683f
C544 B.n451 VSUBS 0.007683f
C545 B.n452 VSUBS 0.007683f
C546 B.n453 VSUBS 0.007683f
C547 B.n454 VSUBS 0.007683f
C548 B.n455 VSUBS 0.007683f
C549 B.n456 VSUBS 0.007683f
C550 B.n457 VSUBS 0.007683f
C551 B.n458 VSUBS 0.007683f
C552 B.n459 VSUBS 0.007683f
C553 B.n460 VSUBS 0.007683f
C554 B.n461 VSUBS 0.007683f
C555 B.n462 VSUBS 0.007683f
C556 B.n463 VSUBS 0.007683f
C557 B.n464 VSUBS 0.007683f
C558 B.n465 VSUBS 0.007683f
C559 B.n466 VSUBS 0.007683f
C560 B.n467 VSUBS 0.007683f
C561 B.n468 VSUBS 0.007683f
C562 B.n469 VSUBS 0.007683f
C563 B.n470 VSUBS 0.007683f
C564 B.n471 VSUBS 0.007683f
C565 B.n472 VSUBS 0.007683f
C566 B.n473 VSUBS 0.007683f
C567 B.n474 VSUBS 0.007683f
C568 B.n475 VSUBS 0.007683f
C569 B.n476 VSUBS 0.007683f
C570 B.n477 VSUBS 0.007683f
C571 B.n478 VSUBS 0.007683f
C572 B.n479 VSUBS 0.007683f
C573 B.n480 VSUBS 0.007683f
C574 B.n481 VSUBS 0.007683f
C575 B.n482 VSUBS 0.007683f
C576 B.n483 VSUBS 0.007683f
C577 B.n484 VSUBS 0.007683f
C578 B.n485 VSUBS 0.007683f
C579 B.n486 VSUBS 0.007683f
C580 B.n487 VSUBS 0.007683f
C581 B.n488 VSUBS 0.007683f
C582 B.n489 VSUBS 0.007683f
C583 B.n490 VSUBS 0.007683f
C584 B.n491 VSUBS 0.007683f
C585 B.n492 VSUBS 0.007683f
C586 B.n493 VSUBS 0.007231f
C587 B.n494 VSUBS 0.007683f
C588 B.n495 VSUBS 0.007683f
C589 B.n496 VSUBS 0.004293f
C590 B.n497 VSUBS 0.007683f
C591 B.n498 VSUBS 0.007683f
C592 B.n499 VSUBS 0.007683f
C593 B.n500 VSUBS 0.007683f
C594 B.n501 VSUBS 0.007683f
C595 B.n502 VSUBS 0.007683f
C596 B.n503 VSUBS 0.007683f
C597 B.n504 VSUBS 0.007683f
C598 B.n505 VSUBS 0.007683f
C599 B.n506 VSUBS 0.007683f
C600 B.n507 VSUBS 0.007683f
C601 B.n508 VSUBS 0.007683f
C602 B.n509 VSUBS 0.004293f
C603 B.n510 VSUBS 0.0178f
C604 B.n511 VSUBS 0.007231f
C605 B.n512 VSUBS 0.007683f
C606 B.n513 VSUBS 0.007683f
C607 B.n514 VSUBS 0.007683f
C608 B.n515 VSUBS 0.007683f
C609 B.n516 VSUBS 0.007683f
C610 B.n517 VSUBS 0.007683f
C611 B.n518 VSUBS 0.007683f
C612 B.n519 VSUBS 0.007683f
C613 B.n520 VSUBS 0.007683f
C614 B.n521 VSUBS 0.007683f
C615 B.n522 VSUBS 0.007683f
C616 B.n523 VSUBS 0.007683f
C617 B.n524 VSUBS 0.007683f
C618 B.n525 VSUBS 0.007683f
C619 B.n526 VSUBS 0.007683f
C620 B.n527 VSUBS 0.007683f
C621 B.n528 VSUBS 0.007683f
C622 B.n529 VSUBS 0.007683f
C623 B.n530 VSUBS 0.007683f
C624 B.n531 VSUBS 0.007683f
C625 B.n532 VSUBS 0.007683f
C626 B.n533 VSUBS 0.007683f
C627 B.n534 VSUBS 0.007683f
C628 B.n535 VSUBS 0.007683f
C629 B.n536 VSUBS 0.007683f
C630 B.n537 VSUBS 0.007683f
C631 B.n538 VSUBS 0.007683f
C632 B.n539 VSUBS 0.007683f
C633 B.n540 VSUBS 0.007683f
C634 B.n541 VSUBS 0.007683f
C635 B.n542 VSUBS 0.007683f
C636 B.n543 VSUBS 0.007683f
C637 B.n544 VSUBS 0.007683f
C638 B.n545 VSUBS 0.007683f
C639 B.n546 VSUBS 0.007683f
C640 B.n547 VSUBS 0.007683f
C641 B.n548 VSUBS 0.007683f
C642 B.n549 VSUBS 0.007683f
C643 B.n550 VSUBS 0.007683f
C644 B.n551 VSUBS 0.007683f
C645 B.n552 VSUBS 0.007683f
C646 B.n553 VSUBS 0.007683f
C647 B.n554 VSUBS 0.007683f
C648 B.n555 VSUBS 0.007683f
C649 B.n556 VSUBS 0.007683f
C650 B.n557 VSUBS 0.007683f
C651 B.n558 VSUBS 0.007683f
C652 B.n559 VSUBS 0.007683f
C653 B.n560 VSUBS 0.007683f
C654 B.n561 VSUBS 0.007683f
C655 B.n562 VSUBS 0.007683f
C656 B.n563 VSUBS 0.007683f
C657 B.n564 VSUBS 0.007683f
C658 B.n565 VSUBS 0.007683f
C659 B.n566 VSUBS 0.007683f
C660 B.n567 VSUBS 0.007683f
C661 B.n568 VSUBS 0.007683f
C662 B.n569 VSUBS 0.007683f
C663 B.n570 VSUBS 0.007683f
C664 B.n571 VSUBS 0.019118f
C665 B.n572 VSUBS 0.019118f
C666 B.n573 VSUBS 0.018391f
C667 B.n574 VSUBS 0.007683f
C668 B.n575 VSUBS 0.007683f
C669 B.n576 VSUBS 0.007683f
C670 B.n577 VSUBS 0.007683f
C671 B.n578 VSUBS 0.007683f
C672 B.n579 VSUBS 0.007683f
C673 B.n580 VSUBS 0.007683f
C674 B.n581 VSUBS 0.007683f
C675 B.n582 VSUBS 0.007683f
C676 B.n583 VSUBS 0.007683f
C677 B.n584 VSUBS 0.007683f
C678 B.n585 VSUBS 0.007683f
C679 B.n586 VSUBS 0.007683f
C680 B.n587 VSUBS 0.007683f
C681 B.n588 VSUBS 0.007683f
C682 B.n589 VSUBS 0.007683f
C683 B.n590 VSUBS 0.007683f
C684 B.n591 VSUBS 0.007683f
C685 B.n592 VSUBS 0.007683f
C686 B.n593 VSUBS 0.007683f
C687 B.n594 VSUBS 0.007683f
C688 B.n595 VSUBS 0.007683f
C689 B.n596 VSUBS 0.007683f
C690 B.n597 VSUBS 0.007683f
C691 B.n598 VSUBS 0.007683f
C692 B.n599 VSUBS 0.007683f
C693 B.n600 VSUBS 0.007683f
C694 B.n601 VSUBS 0.007683f
C695 B.n602 VSUBS 0.007683f
C696 B.n603 VSUBS 0.007683f
C697 B.n604 VSUBS 0.007683f
C698 B.n605 VSUBS 0.007683f
C699 B.n606 VSUBS 0.007683f
C700 B.n607 VSUBS 0.007683f
C701 B.n608 VSUBS 0.007683f
C702 B.n609 VSUBS 0.007683f
C703 B.n610 VSUBS 0.007683f
C704 B.n611 VSUBS 0.007683f
C705 B.n612 VSUBS 0.007683f
C706 B.n613 VSUBS 0.007683f
C707 B.n614 VSUBS 0.007683f
C708 B.n615 VSUBS 0.010026f
C709 B.n616 VSUBS 0.01068f
C710 B.n617 VSUBS 0.021238f
C711 VTAIL.t14 VSUBS 0.228514f
C712 VTAIL.t13 VSUBS 0.228514f
C713 VTAIL.n0 VSUBS 1.67976f
C714 VTAIL.n1 VSUBS 0.626379f
C715 VTAIL.n2 VSUBS 0.013661f
C716 VTAIL.n3 VSUBS 0.030838f
C717 VTAIL.n4 VSUBS 0.013814f
C718 VTAIL.n5 VSUBS 0.02428f
C719 VTAIL.n6 VSUBS 0.013047f
C720 VTAIL.n7 VSUBS 0.030838f
C721 VTAIL.n8 VSUBS 0.013814f
C722 VTAIL.n9 VSUBS 0.02428f
C723 VTAIL.n10 VSUBS 0.013047f
C724 VTAIL.n11 VSUBS 0.030838f
C725 VTAIL.n12 VSUBS 0.013814f
C726 VTAIL.n13 VSUBS 0.02428f
C727 VTAIL.n14 VSUBS 0.013047f
C728 VTAIL.n15 VSUBS 0.030838f
C729 VTAIL.n16 VSUBS 0.013814f
C730 VTAIL.n17 VSUBS 0.02428f
C731 VTAIL.n18 VSUBS 0.013047f
C732 VTAIL.n19 VSUBS 0.030838f
C733 VTAIL.n20 VSUBS 0.013814f
C734 VTAIL.n21 VSUBS 1.20972f
C735 VTAIL.n22 VSUBS 0.013047f
C736 VTAIL.t9 VSUBS 0.065835f
C737 VTAIL.n23 VSUBS 0.149026f
C738 VTAIL.n24 VSUBS 0.019618f
C739 VTAIL.n25 VSUBS 0.023129f
C740 VTAIL.n26 VSUBS 0.030838f
C741 VTAIL.n27 VSUBS 0.013814f
C742 VTAIL.n28 VSUBS 0.013047f
C743 VTAIL.n29 VSUBS 0.02428f
C744 VTAIL.n30 VSUBS 0.02428f
C745 VTAIL.n31 VSUBS 0.013047f
C746 VTAIL.n32 VSUBS 0.013814f
C747 VTAIL.n33 VSUBS 0.030838f
C748 VTAIL.n34 VSUBS 0.030838f
C749 VTAIL.n35 VSUBS 0.013814f
C750 VTAIL.n36 VSUBS 0.013047f
C751 VTAIL.n37 VSUBS 0.02428f
C752 VTAIL.n38 VSUBS 0.02428f
C753 VTAIL.n39 VSUBS 0.013047f
C754 VTAIL.n40 VSUBS 0.013814f
C755 VTAIL.n41 VSUBS 0.030838f
C756 VTAIL.n42 VSUBS 0.030838f
C757 VTAIL.n43 VSUBS 0.013814f
C758 VTAIL.n44 VSUBS 0.013047f
C759 VTAIL.n45 VSUBS 0.02428f
C760 VTAIL.n46 VSUBS 0.02428f
C761 VTAIL.n47 VSUBS 0.013047f
C762 VTAIL.n48 VSUBS 0.013814f
C763 VTAIL.n49 VSUBS 0.030838f
C764 VTAIL.n50 VSUBS 0.030838f
C765 VTAIL.n51 VSUBS 0.013814f
C766 VTAIL.n52 VSUBS 0.013047f
C767 VTAIL.n53 VSUBS 0.02428f
C768 VTAIL.n54 VSUBS 0.02428f
C769 VTAIL.n55 VSUBS 0.013047f
C770 VTAIL.n56 VSUBS 0.013814f
C771 VTAIL.n57 VSUBS 0.030838f
C772 VTAIL.n58 VSUBS 0.030838f
C773 VTAIL.n59 VSUBS 0.013814f
C774 VTAIL.n60 VSUBS 0.013047f
C775 VTAIL.n61 VSUBS 0.02428f
C776 VTAIL.n62 VSUBS 0.061097f
C777 VTAIL.n63 VSUBS 0.013047f
C778 VTAIL.n64 VSUBS 0.013814f
C779 VTAIL.n65 VSUBS 0.066948f
C780 VTAIL.n66 VSUBS 0.044586f
C781 VTAIL.n67 VSUBS 0.157649f
C782 VTAIL.n68 VSUBS 0.013661f
C783 VTAIL.n69 VSUBS 0.030838f
C784 VTAIL.n70 VSUBS 0.013814f
C785 VTAIL.n71 VSUBS 0.02428f
C786 VTAIL.n72 VSUBS 0.013047f
C787 VTAIL.n73 VSUBS 0.030838f
C788 VTAIL.n74 VSUBS 0.013814f
C789 VTAIL.n75 VSUBS 0.02428f
C790 VTAIL.n76 VSUBS 0.013047f
C791 VTAIL.n77 VSUBS 0.030838f
C792 VTAIL.n78 VSUBS 0.013814f
C793 VTAIL.n79 VSUBS 0.02428f
C794 VTAIL.n80 VSUBS 0.013047f
C795 VTAIL.n81 VSUBS 0.030838f
C796 VTAIL.n82 VSUBS 0.013814f
C797 VTAIL.n83 VSUBS 0.02428f
C798 VTAIL.n84 VSUBS 0.013047f
C799 VTAIL.n85 VSUBS 0.030838f
C800 VTAIL.n86 VSUBS 0.013814f
C801 VTAIL.n87 VSUBS 1.20972f
C802 VTAIL.n88 VSUBS 0.013047f
C803 VTAIL.t5 VSUBS 0.065835f
C804 VTAIL.n89 VSUBS 0.149026f
C805 VTAIL.n90 VSUBS 0.019618f
C806 VTAIL.n91 VSUBS 0.023129f
C807 VTAIL.n92 VSUBS 0.030838f
C808 VTAIL.n93 VSUBS 0.013814f
C809 VTAIL.n94 VSUBS 0.013047f
C810 VTAIL.n95 VSUBS 0.02428f
C811 VTAIL.n96 VSUBS 0.02428f
C812 VTAIL.n97 VSUBS 0.013047f
C813 VTAIL.n98 VSUBS 0.013814f
C814 VTAIL.n99 VSUBS 0.030838f
C815 VTAIL.n100 VSUBS 0.030838f
C816 VTAIL.n101 VSUBS 0.013814f
C817 VTAIL.n102 VSUBS 0.013047f
C818 VTAIL.n103 VSUBS 0.02428f
C819 VTAIL.n104 VSUBS 0.02428f
C820 VTAIL.n105 VSUBS 0.013047f
C821 VTAIL.n106 VSUBS 0.013814f
C822 VTAIL.n107 VSUBS 0.030838f
C823 VTAIL.n108 VSUBS 0.030838f
C824 VTAIL.n109 VSUBS 0.013814f
C825 VTAIL.n110 VSUBS 0.013047f
C826 VTAIL.n111 VSUBS 0.02428f
C827 VTAIL.n112 VSUBS 0.02428f
C828 VTAIL.n113 VSUBS 0.013047f
C829 VTAIL.n114 VSUBS 0.013814f
C830 VTAIL.n115 VSUBS 0.030838f
C831 VTAIL.n116 VSUBS 0.030838f
C832 VTAIL.n117 VSUBS 0.013814f
C833 VTAIL.n118 VSUBS 0.013047f
C834 VTAIL.n119 VSUBS 0.02428f
C835 VTAIL.n120 VSUBS 0.02428f
C836 VTAIL.n121 VSUBS 0.013047f
C837 VTAIL.n122 VSUBS 0.013814f
C838 VTAIL.n123 VSUBS 0.030838f
C839 VTAIL.n124 VSUBS 0.030838f
C840 VTAIL.n125 VSUBS 0.013814f
C841 VTAIL.n126 VSUBS 0.013047f
C842 VTAIL.n127 VSUBS 0.02428f
C843 VTAIL.n128 VSUBS 0.061097f
C844 VTAIL.n129 VSUBS 0.013047f
C845 VTAIL.n130 VSUBS 0.013814f
C846 VTAIL.n131 VSUBS 0.066948f
C847 VTAIL.n132 VSUBS 0.044586f
C848 VTAIL.n133 VSUBS 0.157649f
C849 VTAIL.t4 VSUBS 0.228514f
C850 VTAIL.t6 VSUBS 0.228514f
C851 VTAIL.n134 VSUBS 1.67976f
C852 VTAIL.n135 VSUBS 0.720295f
C853 VTAIL.n136 VSUBS 0.013661f
C854 VTAIL.n137 VSUBS 0.030838f
C855 VTAIL.n138 VSUBS 0.013814f
C856 VTAIL.n139 VSUBS 0.02428f
C857 VTAIL.n140 VSUBS 0.013047f
C858 VTAIL.n141 VSUBS 0.030838f
C859 VTAIL.n142 VSUBS 0.013814f
C860 VTAIL.n143 VSUBS 0.02428f
C861 VTAIL.n144 VSUBS 0.013047f
C862 VTAIL.n145 VSUBS 0.030838f
C863 VTAIL.n146 VSUBS 0.013814f
C864 VTAIL.n147 VSUBS 0.02428f
C865 VTAIL.n148 VSUBS 0.013047f
C866 VTAIL.n149 VSUBS 0.030838f
C867 VTAIL.n150 VSUBS 0.013814f
C868 VTAIL.n151 VSUBS 0.02428f
C869 VTAIL.n152 VSUBS 0.013047f
C870 VTAIL.n153 VSUBS 0.030838f
C871 VTAIL.n154 VSUBS 0.013814f
C872 VTAIL.n155 VSUBS 1.20972f
C873 VTAIL.n156 VSUBS 0.013047f
C874 VTAIL.t1 VSUBS 0.065835f
C875 VTAIL.n157 VSUBS 0.149026f
C876 VTAIL.n158 VSUBS 0.019618f
C877 VTAIL.n159 VSUBS 0.023129f
C878 VTAIL.n160 VSUBS 0.030838f
C879 VTAIL.n161 VSUBS 0.013814f
C880 VTAIL.n162 VSUBS 0.013047f
C881 VTAIL.n163 VSUBS 0.02428f
C882 VTAIL.n164 VSUBS 0.02428f
C883 VTAIL.n165 VSUBS 0.013047f
C884 VTAIL.n166 VSUBS 0.013814f
C885 VTAIL.n167 VSUBS 0.030838f
C886 VTAIL.n168 VSUBS 0.030838f
C887 VTAIL.n169 VSUBS 0.013814f
C888 VTAIL.n170 VSUBS 0.013047f
C889 VTAIL.n171 VSUBS 0.02428f
C890 VTAIL.n172 VSUBS 0.02428f
C891 VTAIL.n173 VSUBS 0.013047f
C892 VTAIL.n174 VSUBS 0.013814f
C893 VTAIL.n175 VSUBS 0.030838f
C894 VTAIL.n176 VSUBS 0.030838f
C895 VTAIL.n177 VSUBS 0.013814f
C896 VTAIL.n178 VSUBS 0.013047f
C897 VTAIL.n179 VSUBS 0.02428f
C898 VTAIL.n180 VSUBS 0.02428f
C899 VTAIL.n181 VSUBS 0.013047f
C900 VTAIL.n182 VSUBS 0.013814f
C901 VTAIL.n183 VSUBS 0.030838f
C902 VTAIL.n184 VSUBS 0.030838f
C903 VTAIL.n185 VSUBS 0.013814f
C904 VTAIL.n186 VSUBS 0.013047f
C905 VTAIL.n187 VSUBS 0.02428f
C906 VTAIL.n188 VSUBS 0.02428f
C907 VTAIL.n189 VSUBS 0.013047f
C908 VTAIL.n190 VSUBS 0.013814f
C909 VTAIL.n191 VSUBS 0.030838f
C910 VTAIL.n192 VSUBS 0.030838f
C911 VTAIL.n193 VSUBS 0.013814f
C912 VTAIL.n194 VSUBS 0.013047f
C913 VTAIL.n195 VSUBS 0.02428f
C914 VTAIL.n196 VSUBS 0.061097f
C915 VTAIL.n197 VSUBS 0.013047f
C916 VTAIL.n198 VSUBS 0.013814f
C917 VTAIL.n199 VSUBS 0.066948f
C918 VTAIL.n200 VSUBS 0.044586f
C919 VTAIL.n201 VSUBS 1.35243f
C920 VTAIL.n202 VSUBS 0.013661f
C921 VTAIL.n203 VSUBS 0.030838f
C922 VTAIL.n204 VSUBS 0.013814f
C923 VTAIL.n205 VSUBS 0.02428f
C924 VTAIL.n206 VSUBS 0.013047f
C925 VTAIL.n207 VSUBS 0.030838f
C926 VTAIL.n208 VSUBS 0.013814f
C927 VTAIL.n209 VSUBS 0.02428f
C928 VTAIL.n210 VSUBS 0.013047f
C929 VTAIL.n211 VSUBS 0.030838f
C930 VTAIL.n212 VSUBS 0.013814f
C931 VTAIL.n213 VSUBS 0.02428f
C932 VTAIL.n214 VSUBS 0.013047f
C933 VTAIL.n215 VSUBS 0.030838f
C934 VTAIL.n216 VSUBS 0.013814f
C935 VTAIL.n217 VSUBS 0.02428f
C936 VTAIL.n218 VSUBS 0.013047f
C937 VTAIL.n219 VSUBS 0.030838f
C938 VTAIL.n220 VSUBS 0.013814f
C939 VTAIL.n221 VSUBS 1.20972f
C940 VTAIL.n222 VSUBS 0.013047f
C941 VTAIL.t10 VSUBS 0.065835f
C942 VTAIL.n223 VSUBS 0.149026f
C943 VTAIL.n224 VSUBS 0.019618f
C944 VTAIL.n225 VSUBS 0.023129f
C945 VTAIL.n226 VSUBS 0.030838f
C946 VTAIL.n227 VSUBS 0.013814f
C947 VTAIL.n228 VSUBS 0.013047f
C948 VTAIL.n229 VSUBS 0.02428f
C949 VTAIL.n230 VSUBS 0.02428f
C950 VTAIL.n231 VSUBS 0.013047f
C951 VTAIL.n232 VSUBS 0.013814f
C952 VTAIL.n233 VSUBS 0.030838f
C953 VTAIL.n234 VSUBS 0.030838f
C954 VTAIL.n235 VSUBS 0.013814f
C955 VTAIL.n236 VSUBS 0.013047f
C956 VTAIL.n237 VSUBS 0.02428f
C957 VTAIL.n238 VSUBS 0.02428f
C958 VTAIL.n239 VSUBS 0.013047f
C959 VTAIL.n240 VSUBS 0.013814f
C960 VTAIL.n241 VSUBS 0.030838f
C961 VTAIL.n242 VSUBS 0.030838f
C962 VTAIL.n243 VSUBS 0.013814f
C963 VTAIL.n244 VSUBS 0.013047f
C964 VTAIL.n245 VSUBS 0.02428f
C965 VTAIL.n246 VSUBS 0.02428f
C966 VTAIL.n247 VSUBS 0.013047f
C967 VTAIL.n248 VSUBS 0.013814f
C968 VTAIL.n249 VSUBS 0.030838f
C969 VTAIL.n250 VSUBS 0.030838f
C970 VTAIL.n251 VSUBS 0.013814f
C971 VTAIL.n252 VSUBS 0.013047f
C972 VTAIL.n253 VSUBS 0.02428f
C973 VTAIL.n254 VSUBS 0.02428f
C974 VTAIL.n255 VSUBS 0.013047f
C975 VTAIL.n256 VSUBS 0.013814f
C976 VTAIL.n257 VSUBS 0.030838f
C977 VTAIL.n258 VSUBS 0.030838f
C978 VTAIL.n259 VSUBS 0.013814f
C979 VTAIL.n260 VSUBS 0.013047f
C980 VTAIL.n261 VSUBS 0.02428f
C981 VTAIL.n262 VSUBS 0.061097f
C982 VTAIL.n263 VSUBS 0.013047f
C983 VTAIL.n264 VSUBS 0.013814f
C984 VTAIL.n265 VSUBS 0.066948f
C985 VTAIL.n266 VSUBS 0.044586f
C986 VTAIL.n267 VSUBS 1.35243f
C987 VTAIL.t8 VSUBS 0.228514f
C988 VTAIL.t15 VSUBS 0.228514f
C989 VTAIL.n268 VSUBS 1.67977f
C990 VTAIL.n269 VSUBS 0.720286f
C991 VTAIL.n270 VSUBS 0.013661f
C992 VTAIL.n271 VSUBS 0.030838f
C993 VTAIL.n272 VSUBS 0.013814f
C994 VTAIL.n273 VSUBS 0.02428f
C995 VTAIL.n274 VSUBS 0.013047f
C996 VTAIL.n275 VSUBS 0.030838f
C997 VTAIL.n276 VSUBS 0.013814f
C998 VTAIL.n277 VSUBS 0.02428f
C999 VTAIL.n278 VSUBS 0.013047f
C1000 VTAIL.n279 VSUBS 0.030838f
C1001 VTAIL.n280 VSUBS 0.013814f
C1002 VTAIL.n281 VSUBS 0.02428f
C1003 VTAIL.n282 VSUBS 0.013047f
C1004 VTAIL.n283 VSUBS 0.030838f
C1005 VTAIL.n284 VSUBS 0.013814f
C1006 VTAIL.n285 VSUBS 0.02428f
C1007 VTAIL.n286 VSUBS 0.013047f
C1008 VTAIL.n287 VSUBS 0.030838f
C1009 VTAIL.n288 VSUBS 0.013814f
C1010 VTAIL.n289 VSUBS 1.20972f
C1011 VTAIL.n290 VSUBS 0.013047f
C1012 VTAIL.t12 VSUBS 0.065835f
C1013 VTAIL.n291 VSUBS 0.149026f
C1014 VTAIL.n292 VSUBS 0.019618f
C1015 VTAIL.n293 VSUBS 0.023129f
C1016 VTAIL.n294 VSUBS 0.030838f
C1017 VTAIL.n295 VSUBS 0.013814f
C1018 VTAIL.n296 VSUBS 0.013047f
C1019 VTAIL.n297 VSUBS 0.02428f
C1020 VTAIL.n298 VSUBS 0.02428f
C1021 VTAIL.n299 VSUBS 0.013047f
C1022 VTAIL.n300 VSUBS 0.013814f
C1023 VTAIL.n301 VSUBS 0.030838f
C1024 VTAIL.n302 VSUBS 0.030838f
C1025 VTAIL.n303 VSUBS 0.013814f
C1026 VTAIL.n304 VSUBS 0.013047f
C1027 VTAIL.n305 VSUBS 0.02428f
C1028 VTAIL.n306 VSUBS 0.02428f
C1029 VTAIL.n307 VSUBS 0.013047f
C1030 VTAIL.n308 VSUBS 0.013814f
C1031 VTAIL.n309 VSUBS 0.030838f
C1032 VTAIL.n310 VSUBS 0.030838f
C1033 VTAIL.n311 VSUBS 0.013814f
C1034 VTAIL.n312 VSUBS 0.013047f
C1035 VTAIL.n313 VSUBS 0.02428f
C1036 VTAIL.n314 VSUBS 0.02428f
C1037 VTAIL.n315 VSUBS 0.013047f
C1038 VTAIL.n316 VSUBS 0.013814f
C1039 VTAIL.n317 VSUBS 0.030838f
C1040 VTAIL.n318 VSUBS 0.030838f
C1041 VTAIL.n319 VSUBS 0.013814f
C1042 VTAIL.n320 VSUBS 0.013047f
C1043 VTAIL.n321 VSUBS 0.02428f
C1044 VTAIL.n322 VSUBS 0.02428f
C1045 VTAIL.n323 VSUBS 0.013047f
C1046 VTAIL.n324 VSUBS 0.013814f
C1047 VTAIL.n325 VSUBS 0.030838f
C1048 VTAIL.n326 VSUBS 0.030838f
C1049 VTAIL.n327 VSUBS 0.013814f
C1050 VTAIL.n328 VSUBS 0.013047f
C1051 VTAIL.n329 VSUBS 0.02428f
C1052 VTAIL.n330 VSUBS 0.061097f
C1053 VTAIL.n331 VSUBS 0.013047f
C1054 VTAIL.n332 VSUBS 0.013814f
C1055 VTAIL.n333 VSUBS 0.066948f
C1056 VTAIL.n334 VSUBS 0.044586f
C1057 VTAIL.n335 VSUBS 0.157649f
C1058 VTAIL.n336 VSUBS 0.013661f
C1059 VTAIL.n337 VSUBS 0.030838f
C1060 VTAIL.n338 VSUBS 0.013814f
C1061 VTAIL.n339 VSUBS 0.02428f
C1062 VTAIL.n340 VSUBS 0.013047f
C1063 VTAIL.n341 VSUBS 0.030838f
C1064 VTAIL.n342 VSUBS 0.013814f
C1065 VTAIL.n343 VSUBS 0.02428f
C1066 VTAIL.n344 VSUBS 0.013047f
C1067 VTAIL.n345 VSUBS 0.030838f
C1068 VTAIL.n346 VSUBS 0.013814f
C1069 VTAIL.n347 VSUBS 0.02428f
C1070 VTAIL.n348 VSUBS 0.013047f
C1071 VTAIL.n349 VSUBS 0.030838f
C1072 VTAIL.n350 VSUBS 0.013814f
C1073 VTAIL.n351 VSUBS 0.02428f
C1074 VTAIL.n352 VSUBS 0.013047f
C1075 VTAIL.n353 VSUBS 0.030838f
C1076 VTAIL.n354 VSUBS 0.013814f
C1077 VTAIL.n355 VSUBS 1.20972f
C1078 VTAIL.n356 VSUBS 0.013047f
C1079 VTAIL.t3 VSUBS 0.065835f
C1080 VTAIL.n357 VSUBS 0.149026f
C1081 VTAIL.n358 VSUBS 0.019618f
C1082 VTAIL.n359 VSUBS 0.023129f
C1083 VTAIL.n360 VSUBS 0.030838f
C1084 VTAIL.n361 VSUBS 0.013814f
C1085 VTAIL.n362 VSUBS 0.013047f
C1086 VTAIL.n363 VSUBS 0.02428f
C1087 VTAIL.n364 VSUBS 0.02428f
C1088 VTAIL.n365 VSUBS 0.013047f
C1089 VTAIL.n366 VSUBS 0.013814f
C1090 VTAIL.n367 VSUBS 0.030838f
C1091 VTAIL.n368 VSUBS 0.030838f
C1092 VTAIL.n369 VSUBS 0.013814f
C1093 VTAIL.n370 VSUBS 0.013047f
C1094 VTAIL.n371 VSUBS 0.02428f
C1095 VTAIL.n372 VSUBS 0.02428f
C1096 VTAIL.n373 VSUBS 0.013047f
C1097 VTAIL.n374 VSUBS 0.013814f
C1098 VTAIL.n375 VSUBS 0.030838f
C1099 VTAIL.n376 VSUBS 0.030838f
C1100 VTAIL.n377 VSUBS 0.013814f
C1101 VTAIL.n378 VSUBS 0.013047f
C1102 VTAIL.n379 VSUBS 0.02428f
C1103 VTAIL.n380 VSUBS 0.02428f
C1104 VTAIL.n381 VSUBS 0.013047f
C1105 VTAIL.n382 VSUBS 0.013814f
C1106 VTAIL.n383 VSUBS 0.030838f
C1107 VTAIL.n384 VSUBS 0.030838f
C1108 VTAIL.n385 VSUBS 0.013814f
C1109 VTAIL.n386 VSUBS 0.013047f
C1110 VTAIL.n387 VSUBS 0.02428f
C1111 VTAIL.n388 VSUBS 0.02428f
C1112 VTAIL.n389 VSUBS 0.013047f
C1113 VTAIL.n390 VSUBS 0.013814f
C1114 VTAIL.n391 VSUBS 0.030838f
C1115 VTAIL.n392 VSUBS 0.030838f
C1116 VTAIL.n393 VSUBS 0.013814f
C1117 VTAIL.n394 VSUBS 0.013047f
C1118 VTAIL.n395 VSUBS 0.02428f
C1119 VTAIL.n396 VSUBS 0.061097f
C1120 VTAIL.n397 VSUBS 0.013047f
C1121 VTAIL.n398 VSUBS 0.013814f
C1122 VTAIL.n399 VSUBS 0.066948f
C1123 VTAIL.n400 VSUBS 0.044586f
C1124 VTAIL.n401 VSUBS 0.157649f
C1125 VTAIL.t7 VSUBS 0.228514f
C1126 VTAIL.t0 VSUBS 0.228514f
C1127 VTAIL.n402 VSUBS 1.67977f
C1128 VTAIL.n403 VSUBS 0.720286f
C1129 VTAIL.n404 VSUBS 0.013661f
C1130 VTAIL.n405 VSUBS 0.030838f
C1131 VTAIL.n406 VSUBS 0.013814f
C1132 VTAIL.n407 VSUBS 0.02428f
C1133 VTAIL.n408 VSUBS 0.013047f
C1134 VTAIL.n409 VSUBS 0.030838f
C1135 VTAIL.n410 VSUBS 0.013814f
C1136 VTAIL.n411 VSUBS 0.02428f
C1137 VTAIL.n412 VSUBS 0.013047f
C1138 VTAIL.n413 VSUBS 0.030838f
C1139 VTAIL.n414 VSUBS 0.013814f
C1140 VTAIL.n415 VSUBS 0.02428f
C1141 VTAIL.n416 VSUBS 0.013047f
C1142 VTAIL.n417 VSUBS 0.030838f
C1143 VTAIL.n418 VSUBS 0.013814f
C1144 VTAIL.n419 VSUBS 0.02428f
C1145 VTAIL.n420 VSUBS 0.013047f
C1146 VTAIL.n421 VSUBS 0.030838f
C1147 VTAIL.n422 VSUBS 0.013814f
C1148 VTAIL.n423 VSUBS 1.20972f
C1149 VTAIL.n424 VSUBS 0.013047f
C1150 VTAIL.t2 VSUBS 0.065835f
C1151 VTAIL.n425 VSUBS 0.149026f
C1152 VTAIL.n426 VSUBS 0.019618f
C1153 VTAIL.n427 VSUBS 0.023129f
C1154 VTAIL.n428 VSUBS 0.030838f
C1155 VTAIL.n429 VSUBS 0.013814f
C1156 VTAIL.n430 VSUBS 0.013047f
C1157 VTAIL.n431 VSUBS 0.02428f
C1158 VTAIL.n432 VSUBS 0.02428f
C1159 VTAIL.n433 VSUBS 0.013047f
C1160 VTAIL.n434 VSUBS 0.013814f
C1161 VTAIL.n435 VSUBS 0.030838f
C1162 VTAIL.n436 VSUBS 0.030838f
C1163 VTAIL.n437 VSUBS 0.013814f
C1164 VTAIL.n438 VSUBS 0.013047f
C1165 VTAIL.n439 VSUBS 0.02428f
C1166 VTAIL.n440 VSUBS 0.02428f
C1167 VTAIL.n441 VSUBS 0.013047f
C1168 VTAIL.n442 VSUBS 0.013814f
C1169 VTAIL.n443 VSUBS 0.030838f
C1170 VTAIL.n444 VSUBS 0.030838f
C1171 VTAIL.n445 VSUBS 0.013814f
C1172 VTAIL.n446 VSUBS 0.013047f
C1173 VTAIL.n447 VSUBS 0.02428f
C1174 VTAIL.n448 VSUBS 0.02428f
C1175 VTAIL.n449 VSUBS 0.013047f
C1176 VTAIL.n450 VSUBS 0.013814f
C1177 VTAIL.n451 VSUBS 0.030838f
C1178 VTAIL.n452 VSUBS 0.030838f
C1179 VTAIL.n453 VSUBS 0.013814f
C1180 VTAIL.n454 VSUBS 0.013047f
C1181 VTAIL.n455 VSUBS 0.02428f
C1182 VTAIL.n456 VSUBS 0.02428f
C1183 VTAIL.n457 VSUBS 0.013047f
C1184 VTAIL.n458 VSUBS 0.013814f
C1185 VTAIL.n459 VSUBS 0.030838f
C1186 VTAIL.n460 VSUBS 0.030838f
C1187 VTAIL.n461 VSUBS 0.013814f
C1188 VTAIL.n462 VSUBS 0.013047f
C1189 VTAIL.n463 VSUBS 0.02428f
C1190 VTAIL.n464 VSUBS 0.061097f
C1191 VTAIL.n465 VSUBS 0.013047f
C1192 VTAIL.n466 VSUBS 0.013814f
C1193 VTAIL.n467 VSUBS 0.066948f
C1194 VTAIL.n468 VSUBS 0.044586f
C1195 VTAIL.n469 VSUBS 1.35243f
C1196 VTAIL.n470 VSUBS 0.013661f
C1197 VTAIL.n471 VSUBS 0.030838f
C1198 VTAIL.n472 VSUBS 0.013814f
C1199 VTAIL.n473 VSUBS 0.02428f
C1200 VTAIL.n474 VSUBS 0.013047f
C1201 VTAIL.n475 VSUBS 0.030838f
C1202 VTAIL.n476 VSUBS 0.013814f
C1203 VTAIL.n477 VSUBS 0.02428f
C1204 VTAIL.n478 VSUBS 0.013047f
C1205 VTAIL.n479 VSUBS 0.030838f
C1206 VTAIL.n480 VSUBS 0.013814f
C1207 VTAIL.n481 VSUBS 0.02428f
C1208 VTAIL.n482 VSUBS 0.013047f
C1209 VTAIL.n483 VSUBS 0.030838f
C1210 VTAIL.n484 VSUBS 0.013814f
C1211 VTAIL.n485 VSUBS 0.02428f
C1212 VTAIL.n486 VSUBS 0.013047f
C1213 VTAIL.n487 VSUBS 0.030838f
C1214 VTAIL.n488 VSUBS 0.013814f
C1215 VTAIL.n489 VSUBS 1.20972f
C1216 VTAIL.n490 VSUBS 0.013047f
C1217 VTAIL.t11 VSUBS 0.065835f
C1218 VTAIL.n491 VSUBS 0.149026f
C1219 VTAIL.n492 VSUBS 0.019618f
C1220 VTAIL.n493 VSUBS 0.023129f
C1221 VTAIL.n494 VSUBS 0.030838f
C1222 VTAIL.n495 VSUBS 0.013814f
C1223 VTAIL.n496 VSUBS 0.013047f
C1224 VTAIL.n497 VSUBS 0.02428f
C1225 VTAIL.n498 VSUBS 0.02428f
C1226 VTAIL.n499 VSUBS 0.013047f
C1227 VTAIL.n500 VSUBS 0.013814f
C1228 VTAIL.n501 VSUBS 0.030838f
C1229 VTAIL.n502 VSUBS 0.030838f
C1230 VTAIL.n503 VSUBS 0.013814f
C1231 VTAIL.n504 VSUBS 0.013047f
C1232 VTAIL.n505 VSUBS 0.02428f
C1233 VTAIL.n506 VSUBS 0.02428f
C1234 VTAIL.n507 VSUBS 0.013047f
C1235 VTAIL.n508 VSUBS 0.013814f
C1236 VTAIL.n509 VSUBS 0.030838f
C1237 VTAIL.n510 VSUBS 0.030838f
C1238 VTAIL.n511 VSUBS 0.013814f
C1239 VTAIL.n512 VSUBS 0.013047f
C1240 VTAIL.n513 VSUBS 0.02428f
C1241 VTAIL.n514 VSUBS 0.02428f
C1242 VTAIL.n515 VSUBS 0.013047f
C1243 VTAIL.n516 VSUBS 0.013814f
C1244 VTAIL.n517 VSUBS 0.030838f
C1245 VTAIL.n518 VSUBS 0.030838f
C1246 VTAIL.n519 VSUBS 0.013814f
C1247 VTAIL.n520 VSUBS 0.013047f
C1248 VTAIL.n521 VSUBS 0.02428f
C1249 VTAIL.n522 VSUBS 0.02428f
C1250 VTAIL.n523 VSUBS 0.013047f
C1251 VTAIL.n524 VSUBS 0.013814f
C1252 VTAIL.n525 VSUBS 0.030838f
C1253 VTAIL.n526 VSUBS 0.030838f
C1254 VTAIL.n527 VSUBS 0.013814f
C1255 VTAIL.n528 VSUBS 0.013047f
C1256 VTAIL.n529 VSUBS 0.02428f
C1257 VTAIL.n530 VSUBS 0.061097f
C1258 VTAIL.n531 VSUBS 0.013047f
C1259 VTAIL.n532 VSUBS 0.013814f
C1260 VTAIL.n533 VSUBS 0.066948f
C1261 VTAIL.n534 VSUBS 0.044586f
C1262 VTAIL.n535 VSUBS 1.34788f
C1263 VDD2.t4 VSUBS 0.241472f
C1264 VDD2.t6 VSUBS 0.241472f
C1265 VDD2.n0 VSUBS 1.90707f
C1266 VDD2.t1 VSUBS 0.241472f
C1267 VDD2.t7 VSUBS 0.241472f
C1268 VDD2.n1 VSUBS 1.90707f
C1269 VDD2.n2 VSUBS 2.97724f
C1270 VDD2.t0 VSUBS 0.241472f
C1271 VDD2.t2 VSUBS 0.241472f
C1272 VDD2.n3 VSUBS 1.90243f
C1273 VDD2.n4 VSUBS 2.74584f
C1274 VDD2.t3 VSUBS 0.241472f
C1275 VDD2.t5 VSUBS 0.241472f
C1276 VDD2.n5 VSUBS 1.90704f
C1277 VN.n0 VSUBS 0.058824f
C1278 VN.t2 VSUBS 1.61615f
C1279 VN.n1 VSUBS 0.594793f
C1280 VN.n2 VSUBS 0.232084f
C1281 VN.t1 VSUBS 1.61615f
C1282 VN.t6 VSUBS 1.74288f
C1283 VN.n3 VSUBS 0.653619f
C1284 VN.n4 VSUBS 0.666344f
C1285 VN.n5 VSUBS 0.062732f
C1286 VN.n6 VSUBS 0.062732f
C1287 VN.n7 VSUBS 0.044084f
C1288 VN.n8 VSUBS 0.044084f
C1289 VN.n9 VSUBS 0.04322f
C1290 VN.n10 VSUBS 0.057313f
C1291 VN.t4 VSUBS 1.69247f
C1292 VN.n11 VSUBS 0.672849f
C1293 VN.n12 VSUBS 0.041286f
C1294 VN.n13 VSUBS 0.058824f
C1295 VN.t7 VSUBS 1.61615f
C1296 VN.n14 VSUBS 0.594793f
C1297 VN.n15 VSUBS 0.232084f
C1298 VN.t0 VSUBS 1.61615f
C1299 VN.t3 VSUBS 1.74288f
C1300 VN.n16 VSUBS 0.653619f
C1301 VN.n17 VSUBS 0.666344f
C1302 VN.n18 VSUBS 0.062732f
C1303 VN.n19 VSUBS 0.062732f
C1304 VN.n20 VSUBS 0.044084f
C1305 VN.n21 VSUBS 0.044084f
C1306 VN.n22 VSUBS 0.04322f
C1307 VN.n23 VSUBS 0.057313f
C1308 VN.t5 VSUBS 1.69247f
C1309 VN.n24 VSUBS 0.672849f
C1310 VN.n25 VSUBS 2.01526f
.ends

