* NGSPICE file created from diff_pair_sample_0928.ext - technology: sky130A

.subckt diff_pair_sample_0928 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0.23265 ps=1.74 w=1.41 l=3.33
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0 ps=0 w=1.41 l=3.33
X2 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0.23265 ps=1.74 w=1.41 l=3.33
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0 ps=0 w=1.41 l=3.33
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0 ps=0 w=1.41 l=3.33
X5 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0.23265 ps=1.74 w=1.41 l=3.33
X6 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.23265 pd=1.74 as=0.5499 ps=3.6 w=1.41 l=3.33
X7 VDD2.t3 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.23265 pd=1.74 as=0.5499 ps=3.6 w=1.41 l=3.33
X8 VDD2.t2 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.23265 pd=1.74 as=0.5499 ps=3.6 w=1.41 l=3.33
X9 VTAIL.t4 VN.t3 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0.23265 ps=1.74 w=1.41 l=3.33
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5499 pd=3.6 as=0 ps=0 w=1.41 l=3.33
X11 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.23265 pd=1.74 as=0.5499 ps=3.6 w=1.41 l=3.33
R0 VN.n1 VN.t2 45.208
R1 VN.n0 VN.t3 45.208
R2 VN.n0 VN.t1 44.0817
R3 VN.n1 VN.t0 44.0817
R4 VN VN.n1 43.2305
R5 VN VN.n0 2.44645
R6 VDD2.n2 VDD2.n0 150.214
R7 VDD2.n2 VDD2.n1 115.819
R8 VDD2.n1 VDD2.t0 14.0431
R9 VDD2.n1 VDD2.t2 14.0431
R10 VDD2.n0 VDD2.t1 14.0431
R11 VDD2.n0 VDD2.t3 14.0431
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t2 113.183
R14 VTAIL.n4 VTAIL.t5 113.183
R15 VTAIL.n3 VTAIL.t7 113.183
R16 VTAIL.n7 VTAIL.t6 113.183
R17 VTAIL.n0 VTAIL.t4 113.183
R18 VTAIL.n1 VTAIL.t3 113.183
R19 VTAIL.n2 VTAIL.t1 113.183
R20 VTAIL.n6 VTAIL.t0 113.183
R21 VTAIL.n7 VTAIL.n6 16.7376
R22 VTAIL.n3 VTAIL.n2 16.7376
R23 VTAIL.n4 VTAIL.n3 3.15567
R24 VTAIL.n6 VTAIL.n5 3.15567
R25 VTAIL.n2 VTAIL.n1 3.15567
R26 VTAIL VTAIL.n0 1.63628
R27 VTAIL VTAIL.n7 1.5199
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n491 B.n490 585
R31 B.n492 B.n491 585
R32 B.n155 B.n92 585
R33 B.n154 B.n153 585
R34 B.n152 B.n151 585
R35 B.n150 B.n149 585
R36 B.n148 B.n147 585
R37 B.n146 B.n145 585
R38 B.n144 B.n143 585
R39 B.n142 B.n141 585
R40 B.n140 B.n139 585
R41 B.n138 B.n137 585
R42 B.n136 B.n135 585
R43 B.n134 B.n133 585
R44 B.n132 B.n131 585
R45 B.n130 B.n129 585
R46 B.n128 B.n127 585
R47 B.n126 B.n125 585
R48 B.n124 B.n123 585
R49 B.n122 B.n121 585
R50 B.n120 B.n119 585
R51 B.n117 B.n116 585
R52 B.n115 B.n114 585
R53 B.n113 B.n112 585
R54 B.n111 B.n110 585
R55 B.n109 B.n108 585
R56 B.n107 B.n106 585
R57 B.n105 B.n104 585
R58 B.n103 B.n102 585
R59 B.n101 B.n100 585
R60 B.n99 B.n98 585
R61 B.n75 B.n74 585
R62 B.n489 B.n76 585
R63 B.n493 B.n76 585
R64 B.n488 B.n487 585
R65 B.n487 B.n72 585
R66 B.n486 B.n71 585
R67 B.n499 B.n71 585
R68 B.n485 B.n70 585
R69 B.n500 B.n70 585
R70 B.n484 B.n69 585
R71 B.n501 B.n69 585
R72 B.n483 B.n482 585
R73 B.n482 B.n65 585
R74 B.n481 B.n64 585
R75 B.n507 B.n64 585
R76 B.n480 B.n63 585
R77 B.n508 B.n63 585
R78 B.n479 B.n62 585
R79 B.n509 B.n62 585
R80 B.n478 B.n477 585
R81 B.n477 B.n58 585
R82 B.n476 B.n57 585
R83 B.n515 B.n57 585
R84 B.n475 B.n56 585
R85 B.n516 B.n56 585
R86 B.n474 B.n55 585
R87 B.n517 B.n55 585
R88 B.n473 B.n472 585
R89 B.n472 B.n51 585
R90 B.n471 B.n50 585
R91 B.n523 B.n50 585
R92 B.n470 B.n49 585
R93 B.n524 B.n49 585
R94 B.n469 B.n48 585
R95 B.n525 B.n48 585
R96 B.n468 B.n467 585
R97 B.n467 B.n44 585
R98 B.n466 B.n43 585
R99 B.n531 B.n43 585
R100 B.n465 B.n42 585
R101 B.n532 B.n42 585
R102 B.n464 B.n41 585
R103 B.n533 B.n41 585
R104 B.n463 B.n462 585
R105 B.n462 B.n37 585
R106 B.n461 B.n36 585
R107 B.n539 B.n36 585
R108 B.n460 B.n35 585
R109 B.n540 B.n35 585
R110 B.n459 B.n34 585
R111 B.n541 B.n34 585
R112 B.n458 B.n457 585
R113 B.n457 B.n30 585
R114 B.n456 B.n29 585
R115 B.n547 B.n29 585
R116 B.n455 B.n28 585
R117 B.n548 B.n28 585
R118 B.n454 B.n27 585
R119 B.n549 B.n27 585
R120 B.n453 B.n452 585
R121 B.n452 B.n23 585
R122 B.n451 B.n22 585
R123 B.n555 B.n22 585
R124 B.n450 B.n21 585
R125 B.n556 B.n21 585
R126 B.n449 B.n20 585
R127 B.n557 B.n20 585
R128 B.n448 B.n447 585
R129 B.n447 B.n19 585
R130 B.n446 B.n15 585
R131 B.n563 B.n15 585
R132 B.n445 B.n14 585
R133 B.n564 B.n14 585
R134 B.n444 B.n13 585
R135 B.n565 B.n13 585
R136 B.n443 B.n442 585
R137 B.n442 B.n12 585
R138 B.n441 B.n440 585
R139 B.n441 B.n8 585
R140 B.n439 B.n7 585
R141 B.n572 B.n7 585
R142 B.n438 B.n6 585
R143 B.n573 B.n6 585
R144 B.n437 B.n5 585
R145 B.n574 B.n5 585
R146 B.n436 B.n435 585
R147 B.n435 B.n4 585
R148 B.n434 B.n156 585
R149 B.n434 B.n433 585
R150 B.n424 B.n157 585
R151 B.n158 B.n157 585
R152 B.n426 B.n425 585
R153 B.n427 B.n426 585
R154 B.n423 B.n163 585
R155 B.n163 B.n162 585
R156 B.n422 B.n421 585
R157 B.n421 B.n420 585
R158 B.n165 B.n164 585
R159 B.n413 B.n165 585
R160 B.n412 B.n411 585
R161 B.n414 B.n412 585
R162 B.n410 B.n170 585
R163 B.n170 B.n169 585
R164 B.n409 B.n408 585
R165 B.n408 B.n407 585
R166 B.n172 B.n171 585
R167 B.n173 B.n172 585
R168 B.n400 B.n399 585
R169 B.n401 B.n400 585
R170 B.n398 B.n178 585
R171 B.n178 B.n177 585
R172 B.n397 B.n396 585
R173 B.n396 B.n395 585
R174 B.n180 B.n179 585
R175 B.n181 B.n180 585
R176 B.n388 B.n387 585
R177 B.n389 B.n388 585
R178 B.n386 B.n186 585
R179 B.n186 B.n185 585
R180 B.n385 B.n384 585
R181 B.n384 B.n383 585
R182 B.n188 B.n187 585
R183 B.n189 B.n188 585
R184 B.n376 B.n375 585
R185 B.n377 B.n376 585
R186 B.n374 B.n194 585
R187 B.n194 B.n193 585
R188 B.n373 B.n372 585
R189 B.n372 B.n371 585
R190 B.n196 B.n195 585
R191 B.n197 B.n196 585
R192 B.n364 B.n363 585
R193 B.n365 B.n364 585
R194 B.n362 B.n202 585
R195 B.n202 B.n201 585
R196 B.n361 B.n360 585
R197 B.n360 B.n359 585
R198 B.n204 B.n203 585
R199 B.n205 B.n204 585
R200 B.n352 B.n351 585
R201 B.n353 B.n352 585
R202 B.n350 B.n210 585
R203 B.n210 B.n209 585
R204 B.n349 B.n348 585
R205 B.n348 B.n347 585
R206 B.n212 B.n211 585
R207 B.n213 B.n212 585
R208 B.n340 B.n339 585
R209 B.n341 B.n340 585
R210 B.n338 B.n218 585
R211 B.n218 B.n217 585
R212 B.n337 B.n336 585
R213 B.n336 B.n335 585
R214 B.n220 B.n219 585
R215 B.n221 B.n220 585
R216 B.n328 B.n327 585
R217 B.n329 B.n328 585
R218 B.n326 B.n226 585
R219 B.n226 B.n225 585
R220 B.n325 B.n324 585
R221 B.n324 B.n323 585
R222 B.n228 B.n227 585
R223 B.n229 B.n228 585
R224 B.n316 B.n315 585
R225 B.n317 B.n316 585
R226 B.n232 B.n231 585
R227 B.n253 B.n252 585
R228 B.n254 B.n250 585
R229 B.n250 B.n233 585
R230 B.n256 B.n255 585
R231 B.n258 B.n249 585
R232 B.n261 B.n260 585
R233 B.n262 B.n248 585
R234 B.n264 B.n263 585
R235 B.n266 B.n247 585
R236 B.n269 B.n268 585
R237 B.n270 B.n244 585
R238 B.n273 B.n272 585
R239 B.n275 B.n243 585
R240 B.n278 B.n277 585
R241 B.n279 B.n242 585
R242 B.n281 B.n280 585
R243 B.n283 B.n241 585
R244 B.n286 B.n285 585
R245 B.n287 B.n240 585
R246 B.n292 B.n291 585
R247 B.n294 B.n239 585
R248 B.n297 B.n296 585
R249 B.n298 B.n238 585
R250 B.n300 B.n299 585
R251 B.n302 B.n237 585
R252 B.n305 B.n304 585
R253 B.n306 B.n236 585
R254 B.n308 B.n307 585
R255 B.n310 B.n235 585
R256 B.n313 B.n312 585
R257 B.n314 B.n234 585
R258 B.n319 B.n318 585
R259 B.n318 B.n317 585
R260 B.n320 B.n230 585
R261 B.n230 B.n229 585
R262 B.n322 B.n321 585
R263 B.n323 B.n322 585
R264 B.n224 B.n223 585
R265 B.n225 B.n224 585
R266 B.n331 B.n330 585
R267 B.n330 B.n329 585
R268 B.n332 B.n222 585
R269 B.n222 B.n221 585
R270 B.n334 B.n333 585
R271 B.n335 B.n334 585
R272 B.n216 B.n215 585
R273 B.n217 B.n216 585
R274 B.n343 B.n342 585
R275 B.n342 B.n341 585
R276 B.n344 B.n214 585
R277 B.n214 B.n213 585
R278 B.n346 B.n345 585
R279 B.n347 B.n346 585
R280 B.n208 B.n207 585
R281 B.n209 B.n208 585
R282 B.n355 B.n354 585
R283 B.n354 B.n353 585
R284 B.n356 B.n206 585
R285 B.n206 B.n205 585
R286 B.n358 B.n357 585
R287 B.n359 B.n358 585
R288 B.n200 B.n199 585
R289 B.n201 B.n200 585
R290 B.n367 B.n366 585
R291 B.n366 B.n365 585
R292 B.n368 B.n198 585
R293 B.n198 B.n197 585
R294 B.n370 B.n369 585
R295 B.n371 B.n370 585
R296 B.n192 B.n191 585
R297 B.n193 B.n192 585
R298 B.n379 B.n378 585
R299 B.n378 B.n377 585
R300 B.n380 B.n190 585
R301 B.n190 B.n189 585
R302 B.n382 B.n381 585
R303 B.n383 B.n382 585
R304 B.n184 B.n183 585
R305 B.n185 B.n184 585
R306 B.n391 B.n390 585
R307 B.n390 B.n389 585
R308 B.n392 B.n182 585
R309 B.n182 B.n181 585
R310 B.n394 B.n393 585
R311 B.n395 B.n394 585
R312 B.n176 B.n175 585
R313 B.n177 B.n176 585
R314 B.n403 B.n402 585
R315 B.n402 B.n401 585
R316 B.n404 B.n174 585
R317 B.n174 B.n173 585
R318 B.n406 B.n405 585
R319 B.n407 B.n406 585
R320 B.n168 B.n167 585
R321 B.n169 B.n168 585
R322 B.n416 B.n415 585
R323 B.n415 B.n414 585
R324 B.n417 B.n166 585
R325 B.n413 B.n166 585
R326 B.n419 B.n418 585
R327 B.n420 B.n419 585
R328 B.n161 B.n160 585
R329 B.n162 B.n161 585
R330 B.n429 B.n428 585
R331 B.n428 B.n427 585
R332 B.n430 B.n159 585
R333 B.n159 B.n158 585
R334 B.n432 B.n431 585
R335 B.n433 B.n432 585
R336 B.n3 B.n0 585
R337 B.n4 B.n3 585
R338 B.n571 B.n1 585
R339 B.n572 B.n571 585
R340 B.n570 B.n569 585
R341 B.n570 B.n8 585
R342 B.n568 B.n9 585
R343 B.n12 B.n9 585
R344 B.n567 B.n566 585
R345 B.n566 B.n565 585
R346 B.n11 B.n10 585
R347 B.n564 B.n11 585
R348 B.n562 B.n561 585
R349 B.n563 B.n562 585
R350 B.n560 B.n16 585
R351 B.n19 B.n16 585
R352 B.n559 B.n558 585
R353 B.n558 B.n557 585
R354 B.n18 B.n17 585
R355 B.n556 B.n18 585
R356 B.n554 B.n553 585
R357 B.n555 B.n554 585
R358 B.n552 B.n24 585
R359 B.n24 B.n23 585
R360 B.n551 B.n550 585
R361 B.n550 B.n549 585
R362 B.n26 B.n25 585
R363 B.n548 B.n26 585
R364 B.n546 B.n545 585
R365 B.n547 B.n546 585
R366 B.n544 B.n31 585
R367 B.n31 B.n30 585
R368 B.n543 B.n542 585
R369 B.n542 B.n541 585
R370 B.n33 B.n32 585
R371 B.n540 B.n33 585
R372 B.n538 B.n537 585
R373 B.n539 B.n538 585
R374 B.n536 B.n38 585
R375 B.n38 B.n37 585
R376 B.n535 B.n534 585
R377 B.n534 B.n533 585
R378 B.n40 B.n39 585
R379 B.n532 B.n40 585
R380 B.n530 B.n529 585
R381 B.n531 B.n530 585
R382 B.n528 B.n45 585
R383 B.n45 B.n44 585
R384 B.n527 B.n526 585
R385 B.n526 B.n525 585
R386 B.n47 B.n46 585
R387 B.n524 B.n47 585
R388 B.n522 B.n521 585
R389 B.n523 B.n522 585
R390 B.n520 B.n52 585
R391 B.n52 B.n51 585
R392 B.n519 B.n518 585
R393 B.n518 B.n517 585
R394 B.n54 B.n53 585
R395 B.n516 B.n54 585
R396 B.n514 B.n513 585
R397 B.n515 B.n514 585
R398 B.n512 B.n59 585
R399 B.n59 B.n58 585
R400 B.n511 B.n510 585
R401 B.n510 B.n509 585
R402 B.n61 B.n60 585
R403 B.n508 B.n61 585
R404 B.n506 B.n505 585
R405 B.n507 B.n506 585
R406 B.n504 B.n66 585
R407 B.n66 B.n65 585
R408 B.n503 B.n502 585
R409 B.n502 B.n501 585
R410 B.n68 B.n67 585
R411 B.n500 B.n68 585
R412 B.n498 B.n497 585
R413 B.n499 B.n498 585
R414 B.n496 B.n73 585
R415 B.n73 B.n72 585
R416 B.n495 B.n494 585
R417 B.n494 B.n493 585
R418 B.n575 B.n574 585
R419 B.n573 B.n2 585
R420 B.n494 B.n75 444.452
R421 B.n491 B.n76 444.452
R422 B.n316 B.n234 444.452
R423 B.n318 B.n232 444.452
R424 B.n492 B.n91 256.663
R425 B.n492 B.n90 256.663
R426 B.n492 B.n89 256.663
R427 B.n492 B.n88 256.663
R428 B.n492 B.n87 256.663
R429 B.n492 B.n86 256.663
R430 B.n492 B.n85 256.663
R431 B.n492 B.n84 256.663
R432 B.n492 B.n83 256.663
R433 B.n492 B.n82 256.663
R434 B.n492 B.n81 256.663
R435 B.n492 B.n80 256.663
R436 B.n492 B.n79 256.663
R437 B.n492 B.n78 256.663
R438 B.n492 B.n77 256.663
R439 B.n251 B.n233 256.663
R440 B.n257 B.n233 256.663
R441 B.n259 B.n233 256.663
R442 B.n265 B.n233 256.663
R443 B.n267 B.n233 256.663
R444 B.n274 B.n233 256.663
R445 B.n276 B.n233 256.663
R446 B.n282 B.n233 256.663
R447 B.n284 B.n233 256.663
R448 B.n293 B.n233 256.663
R449 B.n295 B.n233 256.663
R450 B.n301 B.n233 256.663
R451 B.n303 B.n233 256.663
R452 B.n309 B.n233 256.663
R453 B.n311 B.n233 256.663
R454 B.n577 B.n576 256.663
R455 B.n96 B.t4 209.476
R456 B.n93 B.t15 209.476
R457 B.n288 B.t12 209.476
R458 B.n245 B.t8 209.476
R459 B.n317 B.n233 192.522
R460 B.n493 B.n492 192.522
R461 B.n93 B.t16 177.418
R462 B.n288 B.t14 177.418
R463 B.n96 B.t6 177.417
R464 B.n245 B.t11 177.417
R465 B.n100 B.n99 163.367
R466 B.n104 B.n103 163.367
R467 B.n108 B.n107 163.367
R468 B.n112 B.n111 163.367
R469 B.n116 B.n115 163.367
R470 B.n121 B.n120 163.367
R471 B.n125 B.n124 163.367
R472 B.n129 B.n128 163.367
R473 B.n133 B.n132 163.367
R474 B.n137 B.n136 163.367
R475 B.n141 B.n140 163.367
R476 B.n145 B.n144 163.367
R477 B.n149 B.n148 163.367
R478 B.n153 B.n152 163.367
R479 B.n491 B.n92 163.367
R480 B.n316 B.n228 163.367
R481 B.n324 B.n228 163.367
R482 B.n324 B.n226 163.367
R483 B.n328 B.n226 163.367
R484 B.n328 B.n220 163.367
R485 B.n336 B.n220 163.367
R486 B.n336 B.n218 163.367
R487 B.n340 B.n218 163.367
R488 B.n340 B.n212 163.367
R489 B.n348 B.n212 163.367
R490 B.n348 B.n210 163.367
R491 B.n352 B.n210 163.367
R492 B.n352 B.n204 163.367
R493 B.n360 B.n204 163.367
R494 B.n360 B.n202 163.367
R495 B.n364 B.n202 163.367
R496 B.n364 B.n196 163.367
R497 B.n372 B.n196 163.367
R498 B.n372 B.n194 163.367
R499 B.n376 B.n194 163.367
R500 B.n376 B.n188 163.367
R501 B.n384 B.n188 163.367
R502 B.n384 B.n186 163.367
R503 B.n388 B.n186 163.367
R504 B.n388 B.n180 163.367
R505 B.n396 B.n180 163.367
R506 B.n396 B.n178 163.367
R507 B.n400 B.n178 163.367
R508 B.n400 B.n172 163.367
R509 B.n408 B.n172 163.367
R510 B.n408 B.n170 163.367
R511 B.n412 B.n170 163.367
R512 B.n412 B.n165 163.367
R513 B.n421 B.n165 163.367
R514 B.n421 B.n163 163.367
R515 B.n426 B.n163 163.367
R516 B.n426 B.n157 163.367
R517 B.n434 B.n157 163.367
R518 B.n435 B.n434 163.367
R519 B.n435 B.n5 163.367
R520 B.n6 B.n5 163.367
R521 B.n7 B.n6 163.367
R522 B.n441 B.n7 163.367
R523 B.n442 B.n441 163.367
R524 B.n442 B.n13 163.367
R525 B.n14 B.n13 163.367
R526 B.n15 B.n14 163.367
R527 B.n447 B.n15 163.367
R528 B.n447 B.n20 163.367
R529 B.n21 B.n20 163.367
R530 B.n22 B.n21 163.367
R531 B.n452 B.n22 163.367
R532 B.n452 B.n27 163.367
R533 B.n28 B.n27 163.367
R534 B.n29 B.n28 163.367
R535 B.n457 B.n29 163.367
R536 B.n457 B.n34 163.367
R537 B.n35 B.n34 163.367
R538 B.n36 B.n35 163.367
R539 B.n462 B.n36 163.367
R540 B.n462 B.n41 163.367
R541 B.n42 B.n41 163.367
R542 B.n43 B.n42 163.367
R543 B.n467 B.n43 163.367
R544 B.n467 B.n48 163.367
R545 B.n49 B.n48 163.367
R546 B.n50 B.n49 163.367
R547 B.n472 B.n50 163.367
R548 B.n472 B.n55 163.367
R549 B.n56 B.n55 163.367
R550 B.n57 B.n56 163.367
R551 B.n477 B.n57 163.367
R552 B.n477 B.n62 163.367
R553 B.n63 B.n62 163.367
R554 B.n64 B.n63 163.367
R555 B.n482 B.n64 163.367
R556 B.n482 B.n69 163.367
R557 B.n70 B.n69 163.367
R558 B.n71 B.n70 163.367
R559 B.n487 B.n71 163.367
R560 B.n487 B.n76 163.367
R561 B.n252 B.n250 163.367
R562 B.n256 B.n250 163.367
R563 B.n260 B.n258 163.367
R564 B.n264 B.n248 163.367
R565 B.n268 B.n266 163.367
R566 B.n273 B.n244 163.367
R567 B.n277 B.n275 163.367
R568 B.n281 B.n242 163.367
R569 B.n285 B.n283 163.367
R570 B.n292 B.n240 163.367
R571 B.n296 B.n294 163.367
R572 B.n300 B.n238 163.367
R573 B.n304 B.n302 163.367
R574 B.n308 B.n236 163.367
R575 B.n312 B.n310 163.367
R576 B.n318 B.n230 163.367
R577 B.n322 B.n230 163.367
R578 B.n322 B.n224 163.367
R579 B.n330 B.n224 163.367
R580 B.n330 B.n222 163.367
R581 B.n334 B.n222 163.367
R582 B.n334 B.n216 163.367
R583 B.n342 B.n216 163.367
R584 B.n342 B.n214 163.367
R585 B.n346 B.n214 163.367
R586 B.n346 B.n208 163.367
R587 B.n354 B.n208 163.367
R588 B.n354 B.n206 163.367
R589 B.n358 B.n206 163.367
R590 B.n358 B.n200 163.367
R591 B.n366 B.n200 163.367
R592 B.n366 B.n198 163.367
R593 B.n370 B.n198 163.367
R594 B.n370 B.n192 163.367
R595 B.n378 B.n192 163.367
R596 B.n378 B.n190 163.367
R597 B.n382 B.n190 163.367
R598 B.n382 B.n184 163.367
R599 B.n390 B.n184 163.367
R600 B.n390 B.n182 163.367
R601 B.n394 B.n182 163.367
R602 B.n394 B.n176 163.367
R603 B.n402 B.n176 163.367
R604 B.n402 B.n174 163.367
R605 B.n406 B.n174 163.367
R606 B.n406 B.n168 163.367
R607 B.n415 B.n168 163.367
R608 B.n415 B.n166 163.367
R609 B.n419 B.n166 163.367
R610 B.n419 B.n161 163.367
R611 B.n428 B.n161 163.367
R612 B.n428 B.n159 163.367
R613 B.n432 B.n159 163.367
R614 B.n432 B.n3 163.367
R615 B.n575 B.n3 163.367
R616 B.n571 B.n2 163.367
R617 B.n571 B.n570 163.367
R618 B.n570 B.n9 163.367
R619 B.n566 B.n9 163.367
R620 B.n566 B.n11 163.367
R621 B.n562 B.n11 163.367
R622 B.n562 B.n16 163.367
R623 B.n558 B.n16 163.367
R624 B.n558 B.n18 163.367
R625 B.n554 B.n18 163.367
R626 B.n554 B.n24 163.367
R627 B.n550 B.n24 163.367
R628 B.n550 B.n26 163.367
R629 B.n546 B.n26 163.367
R630 B.n546 B.n31 163.367
R631 B.n542 B.n31 163.367
R632 B.n542 B.n33 163.367
R633 B.n538 B.n33 163.367
R634 B.n538 B.n38 163.367
R635 B.n534 B.n38 163.367
R636 B.n534 B.n40 163.367
R637 B.n530 B.n40 163.367
R638 B.n530 B.n45 163.367
R639 B.n526 B.n45 163.367
R640 B.n526 B.n47 163.367
R641 B.n522 B.n47 163.367
R642 B.n522 B.n52 163.367
R643 B.n518 B.n52 163.367
R644 B.n518 B.n54 163.367
R645 B.n514 B.n54 163.367
R646 B.n514 B.n59 163.367
R647 B.n510 B.n59 163.367
R648 B.n510 B.n61 163.367
R649 B.n506 B.n61 163.367
R650 B.n506 B.n66 163.367
R651 B.n502 B.n66 163.367
R652 B.n502 B.n68 163.367
R653 B.n498 B.n68 163.367
R654 B.n498 B.n73 163.367
R655 B.n494 B.n73 163.367
R656 B.n317 B.n229 111.892
R657 B.n323 B.n229 111.892
R658 B.n323 B.n225 111.892
R659 B.n329 B.n225 111.892
R660 B.n329 B.n221 111.892
R661 B.n335 B.n221 111.892
R662 B.n335 B.n217 111.892
R663 B.n341 B.n217 111.892
R664 B.n347 B.n213 111.892
R665 B.n347 B.n209 111.892
R666 B.n353 B.n209 111.892
R667 B.n353 B.n205 111.892
R668 B.n359 B.n205 111.892
R669 B.n359 B.n201 111.892
R670 B.n365 B.n201 111.892
R671 B.n365 B.n197 111.892
R672 B.n371 B.n197 111.892
R673 B.n371 B.n193 111.892
R674 B.n377 B.n193 111.892
R675 B.n377 B.n189 111.892
R676 B.n383 B.n189 111.892
R677 B.n389 B.n185 111.892
R678 B.n389 B.n181 111.892
R679 B.n395 B.n181 111.892
R680 B.n395 B.n177 111.892
R681 B.n401 B.n177 111.892
R682 B.n401 B.n173 111.892
R683 B.n407 B.n173 111.892
R684 B.n407 B.n169 111.892
R685 B.n414 B.n169 111.892
R686 B.n414 B.n413 111.892
R687 B.n420 B.n162 111.892
R688 B.n427 B.n162 111.892
R689 B.n427 B.n158 111.892
R690 B.n433 B.n158 111.892
R691 B.n433 B.n4 111.892
R692 B.n574 B.n4 111.892
R693 B.n574 B.n573 111.892
R694 B.n573 B.n572 111.892
R695 B.n572 B.n8 111.892
R696 B.n12 B.n8 111.892
R697 B.n565 B.n12 111.892
R698 B.n565 B.n564 111.892
R699 B.n564 B.n563 111.892
R700 B.n557 B.n19 111.892
R701 B.n557 B.n556 111.892
R702 B.n556 B.n555 111.892
R703 B.n555 B.n23 111.892
R704 B.n549 B.n23 111.892
R705 B.n549 B.n548 111.892
R706 B.n548 B.n547 111.892
R707 B.n547 B.n30 111.892
R708 B.n541 B.n30 111.892
R709 B.n541 B.n540 111.892
R710 B.n539 B.n37 111.892
R711 B.n533 B.n37 111.892
R712 B.n533 B.n532 111.892
R713 B.n532 B.n531 111.892
R714 B.n531 B.n44 111.892
R715 B.n525 B.n44 111.892
R716 B.n525 B.n524 111.892
R717 B.n524 B.n523 111.892
R718 B.n523 B.n51 111.892
R719 B.n517 B.n51 111.892
R720 B.n517 B.n516 111.892
R721 B.n516 B.n515 111.892
R722 B.n515 B.n58 111.892
R723 B.n509 B.n508 111.892
R724 B.n508 B.n507 111.892
R725 B.n507 B.n65 111.892
R726 B.n501 B.n65 111.892
R727 B.n501 B.n500 111.892
R728 B.n500 B.n499 111.892
R729 B.n499 B.n72 111.892
R730 B.n493 B.n72 111.892
R731 B.n94 B.t17 106.436
R732 B.n289 B.t13 106.436
R733 B.n97 B.t7 106.436
R734 B.n246 B.t10 106.436
R735 B.n341 B.t9 87.2107
R736 B.n509 B.t5 87.2107
R737 B.n383 B.t1 83.9197
R738 B.t0 B.n539 83.9197
R739 B.n77 B.n75 71.676
R740 B.n100 B.n78 71.676
R741 B.n104 B.n79 71.676
R742 B.n108 B.n80 71.676
R743 B.n112 B.n81 71.676
R744 B.n116 B.n82 71.676
R745 B.n121 B.n83 71.676
R746 B.n125 B.n84 71.676
R747 B.n129 B.n85 71.676
R748 B.n133 B.n86 71.676
R749 B.n137 B.n87 71.676
R750 B.n141 B.n88 71.676
R751 B.n145 B.n89 71.676
R752 B.n149 B.n90 71.676
R753 B.n153 B.n91 71.676
R754 B.n92 B.n91 71.676
R755 B.n152 B.n90 71.676
R756 B.n148 B.n89 71.676
R757 B.n144 B.n88 71.676
R758 B.n140 B.n87 71.676
R759 B.n136 B.n86 71.676
R760 B.n132 B.n85 71.676
R761 B.n128 B.n84 71.676
R762 B.n124 B.n83 71.676
R763 B.n120 B.n82 71.676
R764 B.n115 B.n81 71.676
R765 B.n111 B.n80 71.676
R766 B.n107 B.n79 71.676
R767 B.n103 B.n78 71.676
R768 B.n99 B.n77 71.676
R769 B.n251 B.n232 71.676
R770 B.n257 B.n256 71.676
R771 B.n260 B.n259 71.676
R772 B.n265 B.n264 71.676
R773 B.n268 B.n267 71.676
R774 B.n274 B.n273 71.676
R775 B.n277 B.n276 71.676
R776 B.n282 B.n281 71.676
R777 B.n285 B.n284 71.676
R778 B.n293 B.n292 71.676
R779 B.n296 B.n295 71.676
R780 B.n301 B.n300 71.676
R781 B.n304 B.n303 71.676
R782 B.n309 B.n308 71.676
R783 B.n312 B.n311 71.676
R784 B.n252 B.n251 71.676
R785 B.n258 B.n257 71.676
R786 B.n259 B.n248 71.676
R787 B.n266 B.n265 71.676
R788 B.n267 B.n244 71.676
R789 B.n275 B.n274 71.676
R790 B.n276 B.n242 71.676
R791 B.n283 B.n282 71.676
R792 B.n284 B.n240 71.676
R793 B.n294 B.n293 71.676
R794 B.n295 B.n238 71.676
R795 B.n302 B.n301 71.676
R796 B.n303 B.n236 71.676
R797 B.n310 B.n309 71.676
R798 B.n311 B.n234 71.676
R799 B.n576 B.n575 71.676
R800 B.n576 B.n2 71.676
R801 B.n97 B.n96 70.9823
R802 B.n94 B.n93 70.9823
R803 B.n289 B.n288 70.9823
R804 B.n246 B.n245 70.9823
R805 B.n118 B.n97 59.5399
R806 B.n95 B.n94 59.5399
R807 B.n290 B.n289 59.5399
R808 B.n271 B.n246 59.5399
R809 B.n413 B.t3 57.5921
R810 B.n19 B.t2 57.5921
R811 B.n420 B.t3 54.3012
R812 B.n563 B.t2 54.3012
R813 B.n490 B.n489 28.8785
R814 B.n319 B.n231 28.8785
R815 B.n315 B.n314 28.8785
R816 B.n495 B.n74 28.8785
R817 B.t1 B.n185 27.9736
R818 B.n540 B.t0 27.9736
R819 B.t9 B.n213 24.6826
R820 B.t5 B.n58 24.6826
R821 B B.n577 18.0485
R822 B.n320 B.n319 10.6151
R823 B.n321 B.n320 10.6151
R824 B.n321 B.n223 10.6151
R825 B.n331 B.n223 10.6151
R826 B.n332 B.n331 10.6151
R827 B.n333 B.n332 10.6151
R828 B.n333 B.n215 10.6151
R829 B.n343 B.n215 10.6151
R830 B.n344 B.n343 10.6151
R831 B.n345 B.n344 10.6151
R832 B.n345 B.n207 10.6151
R833 B.n355 B.n207 10.6151
R834 B.n356 B.n355 10.6151
R835 B.n357 B.n356 10.6151
R836 B.n357 B.n199 10.6151
R837 B.n367 B.n199 10.6151
R838 B.n368 B.n367 10.6151
R839 B.n369 B.n368 10.6151
R840 B.n369 B.n191 10.6151
R841 B.n379 B.n191 10.6151
R842 B.n380 B.n379 10.6151
R843 B.n381 B.n380 10.6151
R844 B.n381 B.n183 10.6151
R845 B.n391 B.n183 10.6151
R846 B.n392 B.n391 10.6151
R847 B.n393 B.n392 10.6151
R848 B.n393 B.n175 10.6151
R849 B.n403 B.n175 10.6151
R850 B.n404 B.n403 10.6151
R851 B.n405 B.n404 10.6151
R852 B.n405 B.n167 10.6151
R853 B.n416 B.n167 10.6151
R854 B.n417 B.n416 10.6151
R855 B.n418 B.n417 10.6151
R856 B.n418 B.n160 10.6151
R857 B.n429 B.n160 10.6151
R858 B.n430 B.n429 10.6151
R859 B.n431 B.n430 10.6151
R860 B.n431 B.n0 10.6151
R861 B.n253 B.n231 10.6151
R862 B.n254 B.n253 10.6151
R863 B.n255 B.n254 10.6151
R864 B.n255 B.n249 10.6151
R865 B.n261 B.n249 10.6151
R866 B.n262 B.n261 10.6151
R867 B.n263 B.n262 10.6151
R868 B.n263 B.n247 10.6151
R869 B.n269 B.n247 10.6151
R870 B.n270 B.n269 10.6151
R871 B.n272 B.n243 10.6151
R872 B.n278 B.n243 10.6151
R873 B.n279 B.n278 10.6151
R874 B.n280 B.n279 10.6151
R875 B.n280 B.n241 10.6151
R876 B.n286 B.n241 10.6151
R877 B.n287 B.n286 10.6151
R878 B.n291 B.n287 10.6151
R879 B.n297 B.n239 10.6151
R880 B.n298 B.n297 10.6151
R881 B.n299 B.n298 10.6151
R882 B.n299 B.n237 10.6151
R883 B.n305 B.n237 10.6151
R884 B.n306 B.n305 10.6151
R885 B.n307 B.n306 10.6151
R886 B.n307 B.n235 10.6151
R887 B.n313 B.n235 10.6151
R888 B.n314 B.n313 10.6151
R889 B.n315 B.n227 10.6151
R890 B.n325 B.n227 10.6151
R891 B.n326 B.n325 10.6151
R892 B.n327 B.n326 10.6151
R893 B.n327 B.n219 10.6151
R894 B.n337 B.n219 10.6151
R895 B.n338 B.n337 10.6151
R896 B.n339 B.n338 10.6151
R897 B.n339 B.n211 10.6151
R898 B.n349 B.n211 10.6151
R899 B.n350 B.n349 10.6151
R900 B.n351 B.n350 10.6151
R901 B.n351 B.n203 10.6151
R902 B.n361 B.n203 10.6151
R903 B.n362 B.n361 10.6151
R904 B.n363 B.n362 10.6151
R905 B.n363 B.n195 10.6151
R906 B.n373 B.n195 10.6151
R907 B.n374 B.n373 10.6151
R908 B.n375 B.n374 10.6151
R909 B.n375 B.n187 10.6151
R910 B.n385 B.n187 10.6151
R911 B.n386 B.n385 10.6151
R912 B.n387 B.n386 10.6151
R913 B.n387 B.n179 10.6151
R914 B.n397 B.n179 10.6151
R915 B.n398 B.n397 10.6151
R916 B.n399 B.n398 10.6151
R917 B.n399 B.n171 10.6151
R918 B.n409 B.n171 10.6151
R919 B.n410 B.n409 10.6151
R920 B.n411 B.n410 10.6151
R921 B.n411 B.n164 10.6151
R922 B.n422 B.n164 10.6151
R923 B.n423 B.n422 10.6151
R924 B.n425 B.n423 10.6151
R925 B.n425 B.n424 10.6151
R926 B.n424 B.n156 10.6151
R927 B.n436 B.n156 10.6151
R928 B.n437 B.n436 10.6151
R929 B.n438 B.n437 10.6151
R930 B.n439 B.n438 10.6151
R931 B.n440 B.n439 10.6151
R932 B.n443 B.n440 10.6151
R933 B.n444 B.n443 10.6151
R934 B.n445 B.n444 10.6151
R935 B.n446 B.n445 10.6151
R936 B.n448 B.n446 10.6151
R937 B.n449 B.n448 10.6151
R938 B.n450 B.n449 10.6151
R939 B.n451 B.n450 10.6151
R940 B.n453 B.n451 10.6151
R941 B.n454 B.n453 10.6151
R942 B.n455 B.n454 10.6151
R943 B.n456 B.n455 10.6151
R944 B.n458 B.n456 10.6151
R945 B.n459 B.n458 10.6151
R946 B.n460 B.n459 10.6151
R947 B.n461 B.n460 10.6151
R948 B.n463 B.n461 10.6151
R949 B.n464 B.n463 10.6151
R950 B.n465 B.n464 10.6151
R951 B.n466 B.n465 10.6151
R952 B.n468 B.n466 10.6151
R953 B.n469 B.n468 10.6151
R954 B.n470 B.n469 10.6151
R955 B.n471 B.n470 10.6151
R956 B.n473 B.n471 10.6151
R957 B.n474 B.n473 10.6151
R958 B.n475 B.n474 10.6151
R959 B.n476 B.n475 10.6151
R960 B.n478 B.n476 10.6151
R961 B.n479 B.n478 10.6151
R962 B.n480 B.n479 10.6151
R963 B.n481 B.n480 10.6151
R964 B.n483 B.n481 10.6151
R965 B.n484 B.n483 10.6151
R966 B.n485 B.n484 10.6151
R967 B.n486 B.n485 10.6151
R968 B.n488 B.n486 10.6151
R969 B.n489 B.n488 10.6151
R970 B.n569 B.n1 10.6151
R971 B.n569 B.n568 10.6151
R972 B.n568 B.n567 10.6151
R973 B.n567 B.n10 10.6151
R974 B.n561 B.n10 10.6151
R975 B.n561 B.n560 10.6151
R976 B.n560 B.n559 10.6151
R977 B.n559 B.n17 10.6151
R978 B.n553 B.n17 10.6151
R979 B.n553 B.n552 10.6151
R980 B.n552 B.n551 10.6151
R981 B.n551 B.n25 10.6151
R982 B.n545 B.n25 10.6151
R983 B.n545 B.n544 10.6151
R984 B.n544 B.n543 10.6151
R985 B.n543 B.n32 10.6151
R986 B.n537 B.n32 10.6151
R987 B.n537 B.n536 10.6151
R988 B.n536 B.n535 10.6151
R989 B.n535 B.n39 10.6151
R990 B.n529 B.n39 10.6151
R991 B.n529 B.n528 10.6151
R992 B.n528 B.n527 10.6151
R993 B.n527 B.n46 10.6151
R994 B.n521 B.n46 10.6151
R995 B.n521 B.n520 10.6151
R996 B.n520 B.n519 10.6151
R997 B.n519 B.n53 10.6151
R998 B.n513 B.n53 10.6151
R999 B.n513 B.n512 10.6151
R1000 B.n512 B.n511 10.6151
R1001 B.n511 B.n60 10.6151
R1002 B.n505 B.n60 10.6151
R1003 B.n505 B.n504 10.6151
R1004 B.n504 B.n503 10.6151
R1005 B.n503 B.n67 10.6151
R1006 B.n497 B.n67 10.6151
R1007 B.n497 B.n496 10.6151
R1008 B.n496 B.n495 10.6151
R1009 B.n98 B.n74 10.6151
R1010 B.n101 B.n98 10.6151
R1011 B.n102 B.n101 10.6151
R1012 B.n105 B.n102 10.6151
R1013 B.n106 B.n105 10.6151
R1014 B.n109 B.n106 10.6151
R1015 B.n110 B.n109 10.6151
R1016 B.n113 B.n110 10.6151
R1017 B.n114 B.n113 10.6151
R1018 B.n117 B.n114 10.6151
R1019 B.n122 B.n119 10.6151
R1020 B.n123 B.n122 10.6151
R1021 B.n126 B.n123 10.6151
R1022 B.n127 B.n126 10.6151
R1023 B.n130 B.n127 10.6151
R1024 B.n131 B.n130 10.6151
R1025 B.n134 B.n131 10.6151
R1026 B.n135 B.n134 10.6151
R1027 B.n139 B.n138 10.6151
R1028 B.n142 B.n139 10.6151
R1029 B.n143 B.n142 10.6151
R1030 B.n146 B.n143 10.6151
R1031 B.n147 B.n146 10.6151
R1032 B.n150 B.n147 10.6151
R1033 B.n151 B.n150 10.6151
R1034 B.n154 B.n151 10.6151
R1035 B.n155 B.n154 10.6151
R1036 B.n490 B.n155 10.6151
R1037 B.n577 B.n0 8.11757
R1038 B.n577 B.n1 8.11757
R1039 B.n272 B.n271 6.5566
R1040 B.n291 B.n290 6.5566
R1041 B.n119 B.n118 6.5566
R1042 B.n135 B.n95 6.5566
R1043 B.n271 B.n270 4.05904
R1044 B.n290 B.n239 4.05904
R1045 B.n118 B.n117 4.05904
R1046 B.n138 B.n95 4.05904
R1047 VP.n17 VP.n16 161.3
R1048 VP.n15 VP.n1 161.3
R1049 VP.n14 VP.n13 161.3
R1050 VP.n12 VP.n2 161.3
R1051 VP.n11 VP.n10 161.3
R1052 VP.n9 VP.n3 161.3
R1053 VP.n8 VP.n7 161.3
R1054 VP.n6 VP.n4 73.9192
R1055 VP.n18 VP.n0 73.9192
R1056 VP.n5 VP.t1 45.2077
R1057 VP.n5 VP.t3 44.0818
R1058 VP.n6 VP.n5 43.0652
R1059 VP.n10 VP.n2 40.4934
R1060 VP.n14 VP.n2 40.4934
R1061 VP.n9 VP.n8 24.4675
R1062 VP.n10 VP.n9 24.4675
R1063 VP.n15 VP.n14 24.4675
R1064 VP.n16 VP.n15 24.4675
R1065 VP.n8 VP.n4 16.1487
R1066 VP.n16 VP.n0 16.1487
R1067 VP.n4 VP.t0 10.205
R1068 VP.n0 VP.t2 10.205
R1069 VP.n7 VP.n6 0.354971
R1070 VP.n18 VP.n17 0.354971
R1071 VP VP.n18 0.26696
R1072 VP.n7 VP.n3 0.189894
R1073 VP.n11 VP.n3 0.189894
R1074 VP.n12 VP.n11 0.189894
R1075 VP.n13 VP.n12 0.189894
R1076 VP.n13 VP.n1 0.189894
R1077 VP.n17 VP.n1 0.189894
R1078 VDD1 VDD1.n1 150.739
R1079 VDD1 VDD1.n0 115.876
R1080 VDD1.n0 VDD1.t2 14.0431
R1081 VDD1.n0 VDD1.t0 14.0431
R1082 VDD1.n1 VDD1.t3 14.0431
R1083 VDD1.n1 VDD1.t1 14.0431
C0 VP VTAIL 1.70051f
C1 VN VDD1 0.155938f
C2 VDD2 VTAIL 3.34201f
C3 VN VTAIL 1.6864f
C4 VTAIL VDD1 3.28291f
C5 VP VDD2 0.448283f
C6 VN VP 4.76353f
C7 VP VDD1 1.1714f
C8 VN VDD2 0.881425f
C9 VDD2 VDD1 1.19788f
C10 VDD2 B 3.314627f
C11 VDD1 B 6.06943f
C12 VTAIL B 3.535685f
C13 VN B 10.883071f
C14 VP B 9.49571f
C15 VDD1.t2 B 0.025755f
C16 VDD1.t0 B 0.025755f
C17 VDD1.n0 B 0.151371f
C18 VDD1.t3 B 0.025755f
C19 VDD1.t1 B 0.025755f
C20 VDD1.n1 B 0.358252f
C21 VP.t2 B 0.228391f
C22 VP.n0 B 0.212991f
C23 VP.n1 B 0.022731f
C24 VP.n2 B 0.018376f
C25 VP.n3 B 0.022731f
C26 VP.t0 B 0.228391f
C27 VP.n4 B 0.212991f
C28 VP.t1 B 0.456275f
C29 VP.t3 B 0.448304f
C30 VP.n5 B 1.42461f
C31 VP.n6 B 1.03454f
C32 VP.n7 B 0.036687f
C33 VP.n8 B 0.035253f
C34 VP.n9 B 0.042364f
C35 VP.n10 B 0.045177f
C36 VP.n11 B 0.022731f
C37 VP.n12 B 0.022731f
C38 VP.n13 B 0.022731f
C39 VP.n14 B 0.045177f
C40 VP.n15 B 0.042364f
C41 VP.n16 B 0.035253f
C42 VP.n17 B 0.036687f
C43 VP.n18 B 0.053882f
C44 VTAIL.t4 B 0.158047f
C45 VTAIL.n0 B 0.292369f
C46 VTAIL.t3 B 0.158047f
C47 VTAIL.n1 B 0.394408f
C48 VTAIL.t1 B 0.158047f
C49 VTAIL.n2 B 0.939497f
C50 VTAIL.t7 B 0.158048f
C51 VTAIL.n3 B 0.939497f
C52 VTAIL.t5 B 0.158048f
C53 VTAIL.n4 B 0.394408f
C54 VTAIL.t2 B 0.158048f
C55 VTAIL.n5 B 0.394408f
C56 VTAIL.t0 B 0.158047f
C57 VTAIL.n6 B 0.939497f
C58 VTAIL.t6 B 0.158047f
C59 VTAIL.n7 B 0.829642f
C60 VDD2.t1 B 0.026439f
C61 VDD2.t3 B 0.026439f
C62 VDD2.n0 B 0.354358f
C63 VDD2.t0 B 0.026439f
C64 VDD2.t2 B 0.026439f
C65 VDD2.n1 B 0.155184f
C66 VDD2.n2 B 2.43836f
C67 VN.t1 B 0.44534f
C68 VN.t3 B 0.453258f
C69 VN.n0 B 0.314558f
C70 VN.t0 B 0.44534f
C71 VN.t2 B 0.453258f
C72 VN.n1 B 1.42486f
.ends

