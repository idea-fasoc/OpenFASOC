* NGSPICE file created from diff_pair_sample_1688.ext - technology: sky130A

.subckt diff_pair_sample_1688 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=0 ps=0 w=15.46 l=3.54
X1 VDD1.t5 VP.t0 VTAIL.t6 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=6.0294 ps=31.7 w=15.46 l=3.54
X2 B.t8 B.t6 B.t7 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=0 ps=0 w=15.46 l=3.54
X3 VTAIL.t1 VN.t0 VDD2.t5 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=2.5509 ps=15.79 w=15.46 l=3.54
X4 VTAIL.t10 VP.t1 VDD1.t4 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=2.5509 ps=15.79 w=15.46 l=3.54
X5 VDD2.t4 VN.t1 VTAIL.t5 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=2.5509 ps=15.79 w=15.46 l=3.54
X6 VDD1.t3 VP.t2 VTAIL.t8 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=2.5509 ps=15.79 w=15.46 l=3.54
X7 VDD2.t3 VN.t2 VTAIL.t0 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=6.0294 ps=31.7 w=15.46 l=3.54
X8 VTAIL.t2 VN.t3 VDD2.t2 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=2.5509 ps=15.79 w=15.46 l=3.54
X9 VDD1.t2 VP.t3 VTAIL.t7 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=6.0294 ps=31.7 w=15.46 l=3.54
X10 B.t5 B.t3 B.t4 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=0 ps=0 w=15.46 l=3.54
X11 VTAIL.t11 VP.t4 VDD1.t1 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=2.5509 ps=15.79 w=15.46 l=3.54
X12 VDD1.t0 VP.t5 VTAIL.t9 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=2.5509 ps=15.79 w=15.46 l=3.54
X13 VDD2.t1 VN.t4 VTAIL.t3 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=2.5509 pd=15.79 as=6.0294 ps=31.7 w=15.46 l=3.54
X14 B.t2 B.t0 B.t1 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=0 ps=0 w=15.46 l=3.54
X15 VDD2.t0 VN.t5 VTAIL.t4 w_n4066_n4060# sky130_fd_pr__pfet_01v8 ad=6.0294 pd=31.7 as=2.5509 ps=15.79 w=15.46 l=3.54
R0 B.n479 B.n144 585
R1 B.n478 B.n477 585
R2 B.n476 B.n145 585
R3 B.n475 B.n474 585
R4 B.n473 B.n146 585
R5 B.n472 B.n471 585
R6 B.n470 B.n147 585
R7 B.n469 B.n468 585
R8 B.n467 B.n148 585
R9 B.n466 B.n465 585
R10 B.n464 B.n149 585
R11 B.n463 B.n462 585
R12 B.n461 B.n150 585
R13 B.n460 B.n459 585
R14 B.n458 B.n151 585
R15 B.n457 B.n456 585
R16 B.n455 B.n152 585
R17 B.n454 B.n453 585
R18 B.n452 B.n153 585
R19 B.n451 B.n450 585
R20 B.n449 B.n154 585
R21 B.n448 B.n447 585
R22 B.n446 B.n155 585
R23 B.n445 B.n444 585
R24 B.n443 B.n156 585
R25 B.n442 B.n441 585
R26 B.n440 B.n157 585
R27 B.n439 B.n438 585
R28 B.n437 B.n158 585
R29 B.n436 B.n435 585
R30 B.n434 B.n159 585
R31 B.n433 B.n432 585
R32 B.n431 B.n160 585
R33 B.n430 B.n429 585
R34 B.n428 B.n161 585
R35 B.n427 B.n426 585
R36 B.n425 B.n162 585
R37 B.n424 B.n423 585
R38 B.n422 B.n163 585
R39 B.n421 B.n420 585
R40 B.n419 B.n164 585
R41 B.n418 B.n417 585
R42 B.n416 B.n165 585
R43 B.n415 B.n414 585
R44 B.n413 B.n166 585
R45 B.n412 B.n411 585
R46 B.n410 B.n167 585
R47 B.n409 B.n408 585
R48 B.n407 B.n168 585
R49 B.n406 B.n405 585
R50 B.n404 B.n169 585
R51 B.n403 B.n402 585
R52 B.n400 B.n170 585
R53 B.n399 B.n398 585
R54 B.n397 B.n173 585
R55 B.n396 B.n395 585
R56 B.n394 B.n174 585
R57 B.n393 B.n392 585
R58 B.n391 B.n175 585
R59 B.n390 B.n389 585
R60 B.n388 B.n176 585
R61 B.n386 B.n385 585
R62 B.n384 B.n179 585
R63 B.n383 B.n382 585
R64 B.n381 B.n180 585
R65 B.n380 B.n379 585
R66 B.n378 B.n181 585
R67 B.n377 B.n376 585
R68 B.n375 B.n182 585
R69 B.n374 B.n373 585
R70 B.n372 B.n183 585
R71 B.n371 B.n370 585
R72 B.n369 B.n184 585
R73 B.n368 B.n367 585
R74 B.n366 B.n185 585
R75 B.n365 B.n364 585
R76 B.n363 B.n186 585
R77 B.n362 B.n361 585
R78 B.n360 B.n187 585
R79 B.n359 B.n358 585
R80 B.n357 B.n188 585
R81 B.n356 B.n355 585
R82 B.n354 B.n189 585
R83 B.n353 B.n352 585
R84 B.n351 B.n190 585
R85 B.n350 B.n349 585
R86 B.n348 B.n191 585
R87 B.n347 B.n346 585
R88 B.n345 B.n192 585
R89 B.n344 B.n343 585
R90 B.n342 B.n193 585
R91 B.n341 B.n340 585
R92 B.n339 B.n194 585
R93 B.n338 B.n337 585
R94 B.n336 B.n195 585
R95 B.n335 B.n334 585
R96 B.n333 B.n196 585
R97 B.n332 B.n331 585
R98 B.n330 B.n197 585
R99 B.n329 B.n328 585
R100 B.n327 B.n198 585
R101 B.n326 B.n325 585
R102 B.n324 B.n199 585
R103 B.n323 B.n322 585
R104 B.n321 B.n200 585
R105 B.n320 B.n319 585
R106 B.n318 B.n201 585
R107 B.n317 B.n316 585
R108 B.n315 B.n202 585
R109 B.n314 B.n313 585
R110 B.n312 B.n203 585
R111 B.n311 B.n310 585
R112 B.n309 B.n204 585
R113 B.n481 B.n480 585
R114 B.n482 B.n143 585
R115 B.n484 B.n483 585
R116 B.n485 B.n142 585
R117 B.n487 B.n486 585
R118 B.n488 B.n141 585
R119 B.n490 B.n489 585
R120 B.n491 B.n140 585
R121 B.n493 B.n492 585
R122 B.n494 B.n139 585
R123 B.n496 B.n495 585
R124 B.n497 B.n138 585
R125 B.n499 B.n498 585
R126 B.n500 B.n137 585
R127 B.n502 B.n501 585
R128 B.n503 B.n136 585
R129 B.n505 B.n504 585
R130 B.n506 B.n135 585
R131 B.n508 B.n507 585
R132 B.n509 B.n134 585
R133 B.n511 B.n510 585
R134 B.n512 B.n133 585
R135 B.n514 B.n513 585
R136 B.n515 B.n132 585
R137 B.n517 B.n516 585
R138 B.n518 B.n131 585
R139 B.n520 B.n519 585
R140 B.n521 B.n130 585
R141 B.n523 B.n522 585
R142 B.n524 B.n129 585
R143 B.n526 B.n525 585
R144 B.n527 B.n128 585
R145 B.n529 B.n528 585
R146 B.n530 B.n127 585
R147 B.n532 B.n531 585
R148 B.n533 B.n126 585
R149 B.n535 B.n534 585
R150 B.n536 B.n125 585
R151 B.n538 B.n537 585
R152 B.n539 B.n124 585
R153 B.n541 B.n540 585
R154 B.n542 B.n123 585
R155 B.n544 B.n543 585
R156 B.n545 B.n122 585
R157 B.n547 B.n546 585
R158 B.n548 B.n121 585
R159 B.n550 B.n549 585
R160 B.n551 B.n120 585
R161 B.n553 B.n552 585
R162 B.n554 B.n119 585
R163 B.n556 B.n555 585
R164 B.n557 B.n118 585
R165 B.n559 B.n558 585
R166 B.n560 B.n117 585
R167 B.n562 B.n561 585
R168 B.n563 B.n116 585
R169 B.n565 B.n564 585
R170 B.n566 B.n115 585
R171 B.n568 B.n567 585
R172 B.n569 B.n114 585
R173 B.n571 B.n570 585
R174 B.n572 B.n113 585
R175 B.n574 B.n573 585
R176 B.n575 B.n112 585
R177 B.n577 B.n576 585
R178 B.n578 B.n111 585
R179 B.n580 B.n579 585
R180 B.n581 B.n110 585
R181 B.n583 B.n582 585
R182 B.n584 B.n109 585
R183 B.n586 B.n585 585
R184 B.n587 B.n108 585
R185 B.n589 B.n588 585
R186 B.n590 B.n107 585
R187 B.n592 B.n591 585
R188 B.n593 B.n106 585
R189 B.n595 B.n594 585
R190 B.n596 B.n105 585
R191 B.n598 B.n597 585
R192 B.n599 B.n104 585
R193 B.n601 B.n600 585
R194 B.n602 B.n103 585
R195 B.n604 B.n603 585
R196 B.n605 B.n102 585
R197 B.n607 B.n606 585
R198 B.n608 B.n101 585
R199 B.n610 B.n609 585
R200 B.n611 B.n100 585
R201 B.n613 B.n612 585
R202 B.n614 B.n99 585
R203 B.n616 B.n615 585
R204 B.n617 B.n98 585
R205 B.n619 B.n618 585
R206 B.n620 B.n97 585
R207 B.n622 B.n621 585
R208 B.n623 B.n96 585
R209 B.n625 B.n624 585
R210 B.n626 B.n95 585
R211 B.n628 B.n627 585
R212 B.n629 B.n94 585
R213 B.n631 B.n630 585
R214 B.n632 B.n93 585
R215 B.n634 B.n633 585
R216 B.n635 B.n92 585
R217 B.n637 B.n636 585
R218 B.n638 B.n91 585
R219 B.n640 B.n639 585
R220 B.n641 B.n90 585
R221 B.n812 B.n811 585
R222 B.n810 B.n29 585
R223 B.n809 B.n808 585
R224 B.n807 B.n30 585
R225 B.n806 B.n805 585
R226 B.n804 B.n31 585
R227 B.n803 B.n802 585
R228 B.n801 B.n32 585
R229 B.n800 B.n799 585
R230 B.n798 B.n33 585
R231 B.n797 B.n796 585
R232 B.n795 B.n34 585
R233 B.n794 B.n793 585
R234 B.n792 B.n35 585
R235 B.n791 B.n790 585
R236 B.n789 B.n36 585
R237 B.n788 B.n787 585
R238 B.n786 B.n37 585
R239 B.n785 B.n784 585
R240 B.n783 B.n38 585
R241 B.n782 B.n781 585
R242 B.n780 B.n39 585
R243 B.n779 B.n778 585
R244 B.n777 B.n40 585
R245 B.n776 B.n775 585
R246 B.n774 B.n41 585
R247 B.n773 B.n772 585
R248 B.n771 B.n42 585
R249 B.n770 B.n769 585
R250 B.n768 B.n43 585
R251 B.n767 B.n766 585
R252 B.n765 B.n44 585
R253 B.n764 B.n763 585
R254 B.n762 B.n45 585
R255 B.n761 B.n760 585
R256 B.n759 B.n46 585
R257 B.n758 B.n757 585
R258 B.n756 B.n47 585
R259 B.n755 B.n754 585
R260 B.n753 B.n48 585
R261 B.n752 B.n751 585
R262 B.n750 B.n49 585
R263 B.n749 B.n748 585
R264 B.n747 B.n50 585
R265 B.n746 B.n745 585
R266 B.n744 B.n51 585
R267 B.n743 B.n742 585
R268 B.n741 B.n52 585
R269 B.n740 B.n739 585
R270 B.n738 B.n53 585
R271 B.n737 B.n736 585
R272 B.n735 B.n54 585
R273 B.n734 B.n733 585
R274 B.n732 B.n55 585
R275 B.n731 B.n730 585
R276 B.n729 B.n59 585
R277 B.n728 B.n727 585
R278 B.n726 B.n60 585
R279 B.n725 B.n724 585
R280 B.n723 B.n61 585
R281 B.n722 B.n721 585
R282 B.n719 B.n62 585
R283 B.n718 B.n717 585
R284 B.n716 B.n65 585
R285 B.n715 B.n714 585
R286 B.n713 B.n66 585
R287 B.n712 B.n711 585
R288 B.n710 B.n67 585
R289 B.n709 B.n708 585
R290 B.n707 B.n68 585
R291 B.n706 B.n705 585
R292 B.n704 B.n69 585
R293 B.n703 B.n702 585
R294 B.n701 B.n70 585
R295 B.n700 B.n699 585
R296 B.n698 B.n71 585
R297 B.n697 B.n696 585
R298 B.n695 B.n72 585
R299 B.n694 B.n693 585
R300 B.n692 B.n73 585
R301 B.n691 B.n690 585
R302 B.n689 B.n74 585
R303 B.n688 B.n687 585
R304 B.n686 B.n75 585
R305 B.n685 B.n684 585
R306 B.n683 B.n76 585
R307 B.n682 B.n681 585
R308 B.n680 B.n77 585
R309 B.n679 B.n678 585
R310 B.n677 B.n78 585
R311 B.n676 B.n675 585
R312 B.n674 B.n79 585
R313 B.n673 B.n672 585
R314 B.n671 B.n80 585
R315 B.n670 B.n669 585
R316 B.n668 B.n81 585
R317 B.n667 B.n666 585
R318 B.n665 B.n82 585
R319 B.n664 B.n663 585
R320 B.n662 B.n83 585
R321 B.n661 B.n660 585
R322 B.n659 B.n84 585
R323 B.n658 B.n657 585
R324 B.n656 B.n85 585
R325 B.n655 B.n654 585
R326 B.n653 B.n86 585
R327 B.n652 B.n651 585
R328 B.n650 B.n87 585
R329 B.n649 B.n648 585
R330 B.n647 B.n88 585
R331 B.n646 B.n645 585
R332 B.n644 B.n89 585
R333 B.n643 B.n642 585
R334 B.n813 B.n28 585
R335 B.n815 B.n814 585
R336 B.n816 B.n27 585
R337 B.n818 B.n817 585
R338 B.n819 B.n26 585
R339 B.n821 B.n820 585
R340 B.n822 B.n25 585
R341 B.n824 B.n823 585
R342 B.n825 B.n24 585
R343 B.n827 B.n826 585
R344 B.n828 B.n23 585
R345 B.n830 B.n829 585
R346 B.n831 B.n22 585
R347 B.n833 B.n832 585
R348 B.n834 B.n21 585
R349 B.n836 B.n835 585
R350 B.n837 B.n20 585
R351 B.n839 B.n838 585
R352 B.n840 B.n19 585
R353 B.n842 B.n841 585
R354 B.n843 B.n18 585
R355 B.n845 B.n844 585
R356 B.n846 B.n17 585
R357 B.n848 B.n847 585
R358 B.n849 B.n16 585
R359 B.n851 B.n850 585
R360 B.n852 B.n15 585
R361 B.n854 B.n853 585
R362 B.n855 B.n14 585
R363 B.n857 B.n856 585
R364 B.n858 B.n13 585
R365 B.n860 B.n859 585
R366 B.n861 B.n12 585
R367 B.n863 B.n862 585
R368 B.n864 B.n11 585
R369 B.n866 B.n865 585
R370 B.n867 B.n10 585
R371 B.n869 B.n868 585
R372 B.n870 B.n9 585
R373 B.n872 B.n871 585
R374 B.n873 B.n8 585
R375 B.n875 B.n874 585
R376 B.n876 B.n7 585
R377 B.n878 B.n877 585
R378 B.n879 B.n6 585
R379 B.n881 B.n880 585
R380 B.n882 B.n5 585
R381 B.n884 B.n883 585
R382 B.n885 B.n4 585
R383 B.n887 B.n886 585
R384 B.n888 B.n3 585
R385 B.n890 B.n889 585
R386 B.n891 B.n0 585
R387 B.n2 B.n1 585
R388 B.n231 B.n230 585
R389 B.n233 B.n232 585
R390 B.n234 B.n229 585
R391 B.n236 B.n235 585
R392 B.n237 B.n228 585
R393 B.n239 B.n238 585
R394 B.n240 B.n227 585
R395 B.n242 B.n241 585
R396 B.n243 B.n226 585
R397 B.n245 B.n244 585
R398 B.n246 B.n225 585
R399 B.n248 B.n247 585
R400 B.n249 B.n224 585
R401 B.n251 B.n250 585
R402 B.n252 B.n223 585
R403 B.n254 B.n253 585
R404 B.n255 B.n222 585
R405 B.n257 B.n256 585
R406 B.n258 B.n221 585
R407 B.n260 B.n259 585
R408 B.n261 B.n220 585
R409 B.n263 B.n262 585
R410 B.n264 B.n219 585
R411 B.n266 B.n265 585
R412 B.n267 B.n218 585
R413 B.n269 B.n268 585
R414 B.n270 B.n217 585
R415 B.n272 B.n271 585
R416 B.n273 B.n216 585
R417 B.n275 B.n274 585
R418 B.n276 B.n215 585
R419 B.n278 B.n277 585
R420 B.n279 B.n214 585
R421 B.n281 B.n280 585
R422 B.n282 B.n213 585
R423 B.n284 B.n283 585
R424 B.n285 B.n212 585
R425 B.n287 B.n286 585
R426 B.n288 B.n211 585
R427 B.n290 B.n289 585
R428 B.n291 B.n210 585
R429 B.n293 B.n292 585
R430 B.n294 B.n209 585
R431 B.n296 B.n295 585
R432 B.n297 B.n208 585
R433 B.n299 B.n298 585
R434 B.n300 B.n207 585
R435 B.n302 B.n301 585
R436 B.n303 B.n206 585
R437 B.n305 B.n304 585
R438 B.n306 B.n205 585
R439 B.n308 B.n307 585
R440 B.n307 B.n204 535.745
R441 B.n481 B.n144 535.745
R442 B.n643 B.n90 535.745
R443 B.n813 B.n812 535.745
R444 B.n171 B.t7 512.986
R445 B.n63 B.t11 512.986
R446 B.n177 B.t4 512.986
R447 B.n56 B.t2 512.986
R448 B.n172 B.t8 437.933
R449 B.n64 B.t10 437.933
R450 B.n178 B.t5 437.932
R451 B.n57 B.t1 437.932
R452 B.n177 B.t3 314.38
R453 B.n171 B.t6 314.38
R454 B.n63 B.t9 314.38
R455 B.n56 B.t0 314.38
R456 B.n893 B.n892 256.663
R457 B.n892 B.n891 235.042
R458 B.n892 B.n2 235.042
R459 B.n311 B.n204 163.367
R460 B.n312 B.n311 163.367
R461 B.n313 B.n312 163.367
R462 B.n313 B.n202 163.367
R463 B.n317 B.n202 163.367
R464 B.n318 B.n317 163.367
R465 B.n319 B.n318 163.367
R466 B.n319 B.n200 163.367
R467 B.n323 B.n200 163.367
R468 B.n324 B.n323 163.367
R469 B.n325 B.n324 163.367
R470 B.n325 B.n198 163.367
R471 B.n329 B.n198 163.367
R472 B.n330 B.n329 163.367
R473 B.n331 B.n330 163.367
R474 B.n331 B.n196 163.367
R475 B.n335 B.n196 163.367
R476 B.n336 B.n335 163.367
R477 B.n337 B.n336 163.367
R478 B.n337 B.n194 163.367
R479 B.n341 B.n194 163.367
R480 B.n342 B.n341 163.367
R481 B.n343 B.n342 163.367
R482 B.n343 B.n192 163.367
R483 B.n347 B.n192 163.367
R484 B.n348 B.n347 163.367
R485 B.n349 B.n348 163.367
R486 B.n349 B.n190 163.367
R487 B.n353 B.n190 163.367
R488 B.n354 B.n353 163.367
R489 B.n355 B.n354 163.367
R490 B.n355 B.n188 163.367
R491 B.n359 B.n188 163.367
R492 B.n360 B.n359 163.367
R493 B.n361 B.n360 163.367
R494 B.n361 B.n186 163.367
R495 B.n365 B.n186 163.367
R496 B.n366 B.n365 163.367
R497 B.n367 B.n366 163.367
R498 B.n367 B.n184 163.367
R499 B.n371 B.n184 163.367
R500 B.n372 B.n371 163.367
R501 B.n373 B.n372 163.367
R502 B.n373 B.n182 163.367
R503 B.n377 B.n182 163.367
R504 B.n378 B.n377 163.367
R505 B.n379 B.n378 163.367
R506 B.n379 B.n180 163.367
R507 B.n383 B.n180 163.367
R508 B.n384 B.n383 163.367
R509 B.n385 B.n384 163.367
R510 B.n385 B.n176 163.367
R511 B.n390 B.n176 163.367
R512 B.n391 B.n390 163.367
R513 B.n392 B.n391 163.367
R514 B.n392 B.n174 163.367
R515 B.n396 B.n174 163.367
R516 B.n397 B.n396 163.367
R517 B.n398 B.n397 163.367
R518 B.n398 B.n170 163.367
R519 B.n403 B.n170 163.367
R520 B.n404 B.n403 163.367
R521 B.n405 B.n404 163.367
R522 B.n405 B.n168 163.367
R523 B.n409 B.n168 163.367
R524 B.n410 B.n409 163.367
R525 B.n411 B.n410 163.367
R526 B.n411 B.n166 163.367
R527 B.n415 B.n166 163.367
R528 B.n416 B.n415 163.367
R529 B.n417 B.n416 163.367
R530 B.n417 B.n164 163.367
R531 B.n421 B.n164 163.367
R532 B.n422 B.n421 163.367
R533 B.n423 B.n422 163.367
R534 B.n423 B.n162 163.367
R535 B.n427 B.n162 163.367
R536 B.n428 B.n427 163.367
R537 B.n429 B.n428 163.367
R538 B.n429 B.n160 163.367
R539 B.n433 B.n160 163.367
R540 B.n434 B.n433 163.367
R541 B.n435 B.n434 163.367
R542 B.n435 B.n158 163.367
R543 B.n439 B.n158 163.367
R544 B.n440 B.n439 163.367
R545 B.n441 B.n440 163.367
R546 B.n441 B.n156 163.367
R547 B.n445 B.n156 163.367
R548 B.n446 B.n445 163.367
R549 B.n447 B.n446 163.367
R550 B.n447 B.n154 163.367
R551 B.n451 B.n154 163.367
R552 B.n452 B.n451 163.367
R553 B.n453 B.n452 163.367
R554 B.n453 B.n152 163.367
R555 B.n457 B.n152 163.367
R556 B.n458 B.n457 163.367
R557 B.n459 B.n458 163.367
R558 B.n459 B.n150 163.367
R559 B.n463 B.n150 163.367
R560 B.n464 B.n463 163.367
R561 B.n465 B.n464 163.367
R562 B.n465 B.n148 163.367
R563 B.n469 B.n148 163.367
R564 B.n470 B.n469 163.367
R565 B.n471 B.n470 163.367
R566 B.n471 B.n146 163.367
R567 B.n475 B.n146 163.367
R568 B.n476 B.n475 163.367
R569 B.n477 B.n476 163.367
R570 B.n477 B.n144 163.367
R571 B.n639 B.n90 163.367
R572 B.n639 B.n638 163.367
R573 B.n638 B.n637 163.367
R574 B.n637 B.n92 163.367
R575 B.n633 B.n92 163.367
R576 B.n633 B.n632 163.367
R577 B.n632 B.n631 163.367
R578 B.n631 B.n94 163.367
R579 B.n627 B.n94 163.367
R580 B.n627 B.n626 163.367
R581 B.n626 B.n625 163.367
R582 B.n625 B.n96 163.367
R583 B.n621 B.n96 163.367
R584 B.n621 B.n620 163.367
R585 B.n620 B.n619 163.367
R586 B.n619 B.n98 163.367
R587 B.n615 B.n98 163.367
R588 B.n615 B.n614 163.367
R589 B.n614 B.n613 163.367
R590 B.n613 B.n100 163.367
R591 B.n609 B.n100 163.367
R592 B.n609 B.n608 163.367
R593 B.n608 B.n607 163.367
R594 B.n607 B.n102 163.367
R595 B.n603 B.n102 163.367
R596 B.n603 B.n602 163.367
R597 B.n602 B.n601 163.367
R598 B.n601 B.n104 163.367
R599 B.n597 B.n104 163.367
R600 B.n597 B.n596 163.367
R601 B.n596 B.n595 163.367
R602 B.n595 B.n106 163.367
R603 B.n591 B.n106 163.367
R604 B.n591 B.n590 163.367
R605 B.n590 B.n589 163.367
R606 B.n589 B.n108 163.367
R607 B.n585 B.n108 163.367
R608 B.n585 B.n584 163.367
R609 B.n584 B.n583 163.367
R610 B.n583 B.n110 163.367
R611 B.n579 B.n110 163.367
R612 B.n579 B.n578 163.367
R613 B.n578 B.n577 163.367
R614 B.n577 B.n112 163.367
R615 B.n573 B.n112 163.367
R616 B.n573 B.n572 163.367
R617 B.n572 B.n571 163.367
R618 B.n571 B.n114 163.367
R619 B.n567 B.n114 163.367
R620 B.n567 B.n566 163.367
R621 B.n566 B.n565 163.367
R622 B.n565 B.n116 163.367
R623 B.n561 B.n116 163.367
R624 B.n561 B.n560 163.367
R625 B.n560 B.n559 163.367
R626 B.n559 B.n118 163.367
R627 B.n555 B.n118 163.367
R628 B.n555 B.n554 163.367
R629 B.n554 B.n553 163.367
R630 B.n553 B.n120 163.367
R631 B.n549 B.n120 163.367
R632 B.n549 B.n548 163.367
R633 B.n548 B.n547 163.367
R634 B.n547 B.n122 163.367
R635 B.n543 B.n122 163.367
R636 B.n543 B.n542 163.367
R637 B.n542 B.n541 163.367
R638 B.n541 B.n124 163.367
R639 B.n537 B.n124 163.367
R640 B.n537 B.n536 163.367
R641 B.n536 B.n535 163.367
R642 B.n535 B.n126 163.367
R643 B.n531 B.n126 163.367
R644 B.n531 B.n530 163.367
R645 B.n530 B.n529 163.367
R646 B.n529 B.n128 163.367
R647 B.n525 B.n128 163.367
R648 B.n525 B.n524 163.367
R649 B.n524 B.n523 163.367
R650 B.n523 B.n130 163.367
R651 B.n519 B.n130 163.367
R652 B.n519 B.n518 163.367
R653 B.n518 B.n517 163.367
R654 B.n517 B.n132 163.367
R655 B.n513 B.n132 163.367
R656 B.n513 B.n512 163.367
R657 B.n512 B.n511 163.367
R658 B.n511 B.n134 163.367
R659 B.n507 B.n134 163.367
R660 B.n507 B.n506 163.367
R661 B.n506 B.n505 163.367
R662 B.n505 B.n136 163.367
R663 B.n501 B.n136 163.367
R664 B.n501 B.n500 163.367
R665 B.n500 B.n499 163.367
R666 B.n499 B.n138 163.367
R667 B.n495 B.n138 163.367
R668 B.n495 B.n494 163.367
R669 B.n494 B.n493 163.367
R670 B.n493 B.n140 163.367
R671 B.n489 B.n140 163.367
R672 B.n489 B.n488 163.367
R673 B.n488 B.n487 163.367
R674 B.n487 B.n142 163.367
R675 B.n483 B.n142 163.367
R676 B.n483 B.n482 163.367
R677 B.n482 B.n481 163.367
R678 B.n812 B.n29 163.367
R679 B.n808 B.n29 163.367
R680 B.n808 B.n807 163.367
R681 B.n807 B.n806 163.367
R682 B.n806 B.n31 163.367
R683 B.n802 B.n31 163.367
R684 B.n802 B.n801 163.367
R685 B.n801 B.n800 163.367
R686 B.n800 B.n33 163.367
R687 B.n796 B.n33 163.367
R688 B.n796 B.n795 163.367
R689 B.n795 B.n794 163.367
R690 B.n794 B.n35 163.367
R691 B.n790 B.n35 163.367
R692 B.n790 B.n789 163.367
R693 B.n789 B.n788 163.367
R694 B.n788 B.n37 163.367
R695 B.n784 B.n37 163.367
R696 B.n784 B.n783 163.367
R697 B.n783 B.n782 163.367
R698 B.n782 B.n39 163.367
R699 B.n778 B.n39 163.367
R700 B.n778 B.n777 163.367
R701 B.n777 B.n776 163.367
R702 B.n776 B.n41 163.367
R703 B.n772 B.n41 163.367
R704 B.n772 B.n771 163.367
R705 B.n771 B.n770 163.367
R706 B.n770 B.n43 163.367
R707 B.n766 B.n43 163.367
R708 B.n766 B.n765 163.367
R709 B.n765 B.n764 163.367
R710 B.n764 B.n45 163.367
R711 B.n760 B.n45 163.367
R712 B.n760 B.n759 163.367
R713 B.n759 B.n758 163.367
R714 B.n758 B.n47 163.367
R715 B.n754 B.n47 163.367
R716 B.n754 B.n753 163.367
R717 B.n753 B.n752 163.367
R718 B.n752 B.n49 163.367
R719 B.n748 B.n49 163.367
R720 B.n748 B.n747 163.367
R721 B.n747 B.n746 163.367
R722 B.n746 B.n51 163.367
R723 B.n742 B.n51 163.367
R724 B.n742 B.n741 163.367
R725 B.n741 B.n740 163.367
R726 B.n740 B.n53 163.367
R727 B.n736 B.n53 163.367
R728 B.n736 B.n735 163.367
R729 B.n735 B.n734 163.367
R730 B.n734 B.n55 163.367
R731 B.n730 B.n55 163.367
R732 B.n730 B.n729 163.367
R733 B.n729 B.n728 163.367
R734 B.n728 B.n60 163.367
R735 B.n724 B.n60 163.367
R736 B.n724 B.n723 163.367
R737 B.n723 B.n722 163.367
R738 B.n722 B.n62 163.367
R739 B.n717 B.n62 163.367
R740 B.n717 B.n716 163.367
R741 B.n716 B.n715 163.367
R742 B.n715 B.n66 163.367
R743 B.n711 B.n66 163.367
R744 B.n711 B.n710 163.367
R745 B.n710 B.n709 163.367
R746 B.n709 B.n68 163.367
R747 B.n705 B.n68 163.367
R748 B.n705 B.n704 163.367
R749 B.n704 B.n703 163.367
R750 B.n703 B.n70 163.367
R751 B.n699 B.n70 163.367
R752 B.n699 B.n698 163.367
R753 B.n698 B.n697 163.367
R754 B.n697 B.n72 163.367
R755 B.n693 B.n72 163.367
R756 B.n693 B.n692 163.367
R757 B.n692 B.n691 163.367
R758 B.n691 B.n74 163.367
R759 B.n687 B.n74 163.367
R760 B.n687 B.n686 163.367
R761 B.n686 B.n685 163.367
R762 B.n685 B.n76 163.367
R763 B.n681 B.n76 163.367
R764 B.n681 B.n680 163.367
R765 B.n680 B.n679 163.367
R766 B.n679 B.n78 163.367
R767 B.n675 B.n78 163.367
R768 B.n675 B.n674 163.367
R769 B.n674 B.n673 163.367
R770 B.n673 B.n80 163.367
R771 B.n669 B.n80 163.367
R772 B.n669 B.n668 163.367
R773 B.n668 B.n667 163.367
R774 B.n667 B.n82 163.367
R775 B.n663 B.n82 163.367
R776 B.n663 B.n662 163.367
R777 B.n662 B.n661 163.367
R778 B.n661 B.n84 163.367
R779 B.n657 B.n84 163.367
R780 B.n657 B.n656 163.367
R781 B.n656 B.n655 163.367
R782 B.n655 B.n86 163.367
R783 B.n651 B.n86 163.367
R784 B.n651 B.n650 163.367
R785 B.n650 B.n649 163.367
R786 B.n649 B.n88 163.367
R787 B.n645 B.n88 163.367
R788 B.n645 B.n644 163.367
R789 B.n644 B.n643 163.367
R790 B.n814 B.n813 163.367
R791 B.n814 B.n27 163.367
R792 B.n818 B.n27 163.367
R793 B.n819 B.n818 163.367
R794 B.n820 B.n819 163.367
R795 B.n820 B.n25 163.367
R796 B.n824 B.n25 163.367
R797 B.n825 B.n824 163.367
R798 B.n826 B.n825 163.367
R799 B.n826 B.n23 163.367
R800 B.n830 B.n23 163.367
R801 B.n831 B.n830 163.367
R802 B.n832 B.n831 163.367
R803 B.n832 B.n21 163.367
R804 B.n836 B.n21 163.367
R805 B.n837 B.n836 163.367
R806 B.n838 B.n837 163.367
R807 B.n838 B.n19 163.367
R808 B.n842 B.n19 163.367
R809 B.n843 B.n842 163.367
R810 B.n844 B.n843 163.367
R811 B.n844 B.n17 163.367
R812 B.n848 B.n17 163.367
R813 B.n849 B.n848 163.367
R814 B.n850 B.n849 163.367
R815 B.n850 B.n15 163.367
R816 B.n854 B.n15 163.367
R817 B.n855 B.n854 163.367
R818 B.n856 B.n855 163.367
R819 B.n856 B.n13 163.367
R820 B.n860 B.n13 163.367
R821 B.n861 B.n860 163.367
R822 B.n862 B.n861 163.367
R823 B.n862 B.n11 163.367
R824 B.n866 B.n11 163.367
R825 B.n867 B.n866 163.367
R826 B.n868 B.n867 163.367
R827 B.n868 B.n9 163.367
R828 B.n872 B.n9 163.367
R829 B.n873 B.n872 163.367
R830 B.n874 B.n873 163.367
R831 B.n874 B.n7 163.367
R832 B.n878 B.n7 163.367
R833 B.n879 B.n878 163.367
R834 B.n880 B.n879 163.367
R835 B.n880 B.n5 163.367
R836 B.n884 B.n5 163.367
R837 B.n885 B.n884 163.367
R838 B.n886 B.n885 163.367
R839 B.n886 B.n3 163.367
R840 B.n890 B.n3 163.367
R841 B.n891 B.n890 163.367
R842 B.n230 B.n2 163.367
R843 B.n233 B.n230 163.367
R844 B.n234 B.n233 163.367
R845 B.n235 B.n234 163.367
R846 B.n235 B.n228 163.367
R847 B.n239 B.n228 163.367
R848 B.n240 B.n239 163.367
R849 B.n241 B.n240 163.367
R850 B.n241 B.n226 163.367
R851 B.n245 B.n226 163.367
R852 B.n246 B.n245 163.367
R853 B.n247 B.n246 163.367
R854 B.n247 B.n224 163.367
R855 B.n251 B.n224 163.367
R856 B.n252 B.n251 163.367
R857 B.n253 B.n252 163.367
R858 B.n253 B.n222 163.367
R859 B.n257 B.n222 163.367
R860 B.n258 B.n257 163.367
R861 B.n259 B.n258 163.367
R862 B.n259 B.n220 163.367
R863 B.n263 B.n220 163.367
R864 B.n264 B.n263 163.367
R865 B.n265 B.n264 163.367
R866 B.n265 B.n218 163.367
R867 B.n269 B.n218 163.367
R868 B.n270 B.n269 163.367
R869 B.n271 B.n270 163.367
R870 B.n271 B.n216 163.367
R871 B.n275 B.n216 163.367
R872 B.n276 B.n275 163.367
R873 B.n277 B.n276 163.367
R874 B.n277 B.n214 163.367
R875 B.n281 B.n214 163.367
R876 B.n282 B.n281 163.367
R877 B.n283 B.n282 163.367
R878 B.n283 B.n212 163.367
R879 B.n287 B.n212 163.367
R880 B.n288 B.n287 163.367
R881 B.n289 B.n288 163.367
R882 B.n289 B.n210 163.367
R883 B.n293 B.n210 163.367
R884 B.n294 B.n293 163.367
R885 B.n295 B.n294 163.367
R886 B.n295 B.n208 163.367
R887 B.n299 B.n208 163.367
R888 B.n300 B.n299 163.367
R889 B.n301 B.n300 163.367
R890 B.n301 B.n206 163.367
R891 B.n305 B.n206 163.367
R892 B.n306 B.n305 163.367
R893 B.n307 B.n306 163.367
R894 B.n178 B.n177 75.0551
R895 B.n172 B.n171 75.0551
R896 B.n64 B.n63 75.0551
R897 B.n57 B.n56 75.0551
R898 B.n387 B.n178 59.5399
R899 B.n401 B.n172 59.5399
R900 B.n720 B.n64 59.5399
R901 B.n58 B.n57 59.5399
R902 B.n811 B.n28 34.8103
R903 B.n642 B.n641 34.8103
R904 B.n480 B.n479 34.8103
R905 B.n309 B.n308 34.8103
R906 B B.n893 18.0485
R907 B.n815 B.n28 10.6151
R908 B.n816 B.n815 10.6151
R909 B.n817 B.n816 10.6151
R910 B.n817 B.n26 10.6151
R911 B.n821 B.n26 10.6151
R912 B.n822 B.n821 10.6151
R913 B.n823 B.n822 10.6151
R914 B.n823 B.n24 10.6151
R915 B.n827 B.n24 10.6151
R916 B.n828 B.n827 10.6151
R917 B.n829 B.n828 10.6151
R918 B.n829 B.n22 10.6151
R919 B.n833 B.n22 10.6151
R920 B.n834 B.n833 10.6151
R921 B.n835 B.n834 10.6151
R922 B.n835 B.n20 10.6151
R923 B.n839 B.n20 10.6151
R924 B.n840 B.n839 10.6151
R925 B.n841 B.n840 10.6151
R926 B.n841 B.n18 10.6151
R927 B.n845 B.n18 10.6151
R928 B.n846 B.n845 10.6151
R929 B.n847 B.n846 10.6151
R930 B.n847 B.n16 10.6151
R931 B.n851 B.n16 10.6151
R932 B.n852 B.n851 10.6151
R933 B.n853 B.n852 10.6151
R934 B.n853 B.n14 10.6151
R935 B.n857 B.n14 10.6151
R936 B.n858 B.n857 10.6151
R937 B.n859 B.n858 10.6151
R938 B.n859 B.n12 10.6151
R939 B.n863 B.n12 10.6151
R940 B.n864 B.n863 10.6151
R941 B.n865 B.n864 10.6151
R942 B.n865 B.n10 10.6151
R943 B.n869 B.n10 10.6151
R944 B.n870 B.n869 10.6151
R945 B.n871 B.n870 10.6151
R946 B.n871 B.n8 10.6151
R947 B.n875 B.n8 10.6151
R948 B.n876 B.n875 10.6151
R949 B.n877 B.n876 10.6151
R950 B.n877 B.n6 10.6151
R951 B.n881 B.n6 10.6151
R952 B.n882 B.n881 10.6151
R953 B.n883 B.n882 10.6151
R954 B.n883 B.n4 10.6151
R955 B.n887 B.n4 10.6151
R956 B.n888 B.n887 10.6151
R957 B.n889 B.n888 10.6151
R958 B.n889 B.n0 10.6151
R959 B.n811 B.n810 10.6151
R960 B.n810 B.n809 10.6151
R961 B.n809 B.n30 10.6151
R962 B.n805 B.n30 10.6151
R963 B.n805 B.n804 10.6151
R964 B.n804 B.n803 10.6151
R965 B.n803 B.n32 10.6151
R966 B.n799 B.n32 10.6151
R967 B.n799 B.n798 10.6151
R968 B.n798 B.n797 10.6151
R969 B.n797 B.n34 10.6151
R970 B.n793 B.n34 10.6151
R971 B.n793 B.n792 10.6151
R972 B.n792 B.n791 10.6151
R973 B.n791 B.n36 10.6151
R974 B.n787 B.n36 10.6151
R975 B.n787 B.n786 10.6151
R976 B.n786 B.n785 10.6151
R977 B.n785 B.n38 10.6151
R978 B.n781 B.n38 10.6151
R979 B.n781 B.n780 10.6151
R980 B.n780 B.n779 10.6151
R981 B.n779 B.n40 10.6151
R982 B.n775 B.n40 10.6151
R983 B.n775 B.n774 10.6151
R984 B.n774 B.n773 10.6151
R985 B.n773 B.n42 10.6151
R986 B.n769 B.n42 10.6151
R987 B.n769 B.n768 10.6151
R988 B.n768 B.n767 10.6151
R989 B.n767 B.n44 10.6151
R990 B.n763 B.n44 10.6151
R991 B.n763 B.n762 10.6151
R992 B.n762 B.n761 10.6151
R993 B.n761 B.n46 10.6151
R994 B.n757 B.n46 10.6151
R995 B.n757 B.n756 10.6151
R996 B.n756 B.n755 10.6151
R997 B.n755 B.n48 10.6151
R998 B.n751 B.n48 10.6151
R999 B.n751 B.n750 10.6151
R1000 B.n750 B.n749 10.6151
R1001 B.n749 B.n50 10.6151
R1002 B.n745 B.n50 10.6151
R1003 B.n745 B.n744 10.6151
R1004 B.n744 B.n743 10.6151
R1005 B.n743 B.n52 10.6151
R1006 B.n739 B.n52 10.6151
R1007 B.n739 B.n738 10.6151
R1008 B.n738 B.n737 10.6151
R1009 B.n737 B.n54 10.6151
R1010 B.n733 B.n732 10.6151
R1011 B.n732 B.n731 10.6151
R1012 B.n731 B.n59 10.6151
R1013 B.n727 B.n59 10.6151
R1014 B.n727 B.n726 10.6151
R1015 B.n726 B.n725 10.6151
R1016 B.n725 B.n61 10.6151
R1017 B.n721 B.n61 10.6151
R1018 B.n719 B.n718 10.6151
R1019 B.n718 B.n65 10.6151
R1020 B.n714 B.n65 10.6151
R1021 B.n714 B.n713 10.6151
R1022 B.n713 B.n712 10.6151
R1023 B.n712 B.n67 10.6151
R1024 B.n708 B.n67 10.6151
R1025 B.n708 B.n707 10.6151
R1026 B.n707 B.n706 10.6151
R1027 B.n706 B.n69 10.6151
R1028 B.n702 B.n69 10.6151
R1029 B.n702 B.n701 10.6151
R1030 B.n701 B.n700 10.6151
R1031 B.n700 B.n71 10.6151
R1032 B.n696 B.n71 10.6151
R1033 B.n696 B.n695 10.6151
R1034 B.n695 B.n694 10.6151
R1035 B.n694 B.n73 10.6151
R1036 B.n690 B.n73 10.6151
R1037 B.n690 B.n689 10.6151
R1038 B.n689 B.n688 10.6151
R1039 B.n688 B.n75 10.6151
R1040 B.n684 B.n75 10.6151
R1041 B.n684 B.n683 10.6151
R1042 B.n683 B.n682 10.6151
R1043 B.n682 B.n77 10.6151
R1044 B.n678 B.n77 10.6151
R1045 B.n678 B.n677 10.6151
R1046 B.n677 B.n676 10.6151
R1047 B.n676 B.n79 10.6151
R1048 B.n672 B.n79 10.6151
R1049 B.n672 B.n671 10.6151
R1050 B.n671 B.n670 10.6151
R1051 B.n670 B.n81 10.6151
R1052 B.n666 B.n81 10.6151
R1053 B.n666 B.n665 10.6151
R1054 B.n665 B.n664 10.6151
R1055 B.n664 B.n83 10.6151
R1056 B.n660 B.n83 10.6151
R1057 B.n660 B.n659 10.6151
R1058 B.n659 B.n658 10.6151
R1059 B.n658 B.n85 10.6151
R1060 B.n654 B.n85 10.6151
R1061 B.n654 B.n653 10.6151
R1062 B.n653 B.n652 10.6151
R1063 B.n652 B.n87 10.6151
R1064 B.n648 B.n87 10.6151
R1065 B.n648 B.n647 10.6151
R1066 B.n647 B.n646 10.6151
R1067 B.n646 B.n89 10.6151
R1068 B.n642 B.n89 10.6151
R1069 B.n641 B.n640 10.6151
R1070 B.n640 B.n91 10.6151
R1071 B.n636 B.n91 10.6151
R1072 B.n636 B.n635 10.6151
R1073 B.n635 B.n634 10.6151
R1074 B.n634 B.n93 10.6151
R1075 B.n630 B.n93 10.6151
R1076 B.n630 B.n629 10.6151
R1077 B.n629 B.n628 10.6151
R1078 B.n628 B.n95 10.6151
R1079 B.n624 B.n95 10.6151
R1080 B.n624 B.n623 10.6151
R1081 B.n623 B.n622 10.6151
R1082 B.n622 B.n97 10.6151
R1083 B.n618 B.n97 10.6151
R1084 B.n618 B.n617 10.6151
R1085 B.n617 B.n616 10.6151
R1086 B.n616 B.n99 10.6151
R1087 B.n612 B.n99 10.6151
R1088 B.n612 B.n611 10.6151
R1089 B.n611 B.n610 10.6151
R1090 B.n610 B.n101 10.6151
R1091 B.n606 B.n101 10.6151
R1092 B.n606 B.n605 10.6151
R1093 B.n605 B.n604 10.6151
R1094 B.n604 B.n103 10.6151
R1095 B.n600 B.n103 10.6151
R1096 B.n600 B.n599 10.6151
R1097 B.n599 B.n598 10.6151
R1098 B.n598 B.n105 10.6151
R1099 B.n594 B.n105 10.6151
R1100 B.n594 B.n593 10.6151
R1101 B.n593 B.n592 10.6151
R1102 B.n592 B.n107 10.6151
R1103 B.n588 B.n107 10.6151
R1104 B.n588 B.n587 10.6151
R1105 B.n587 B.n586 10.6151
R1106 B.n586 B.n109 10.6151
R1107 B.n582 B.n109 10.6151
R1108 B.n582 B.n581 10.6151
R1109 B.n581 B.n580 10.6151
R1110 B.n580 B.n111 10.6151
R1111 B.n576 B.n111 10.6151
R1112 B.n576 B.n575 10.6151
R1113 B.n575 B.n574 10.6151
R1114 B.n574 B.n113 10.6151
R1115 B.n570 B.n113 10.6151
R1116 B.n570 B.n569 10.6151
R1117 B.n569 B.n568 10.6151
R1118 B.n568 B.n115 10.6151
R1119 B.n564 B.n115 10.6151
R1120 B.n564 B.n563 10.6151
R1121 B.n563 B.n562 10.6151
R1122 B.n562 B.n117 10.6151
R1123 B.n558 B.n117 10.6151
R1124 B.n558 B.n557 10.6151
R1125 B.n557 B.n556 10.6151
R1126 B.n556 B.n119 10.6151
R1127 B.n552 B.n119 10.6151
R1128 B.n552 B.n551 10.6151
R1129 B.n551 B.n550 10.6151
R1130 B.n550 B.n121 10.6151
R1131 B.n546 B.n121 10.6151
R1132 B.n546 B.n545 10.6151
R1133 B.n545 B.n544 10.6151
R1134 B.n544 B.n123 10.6151
R1135 B.n540 B.n123 10.6151
R1136 B.n540 B.n539 10.6151
R1137 B.n539 B.n538 10.6151
R1138 B.n538 B.n125 10.6151
R1139 B.n534 B.n125 10.6151
R1140 B.n534 B.n533 10.6151
R1141 B.n533 B.n532 10.6151
R1142 B.n532 B.n127 10.6151
R1143 B.n528 B.n127 10.6151
R1144 B.n528 B.n527 10.6151
R1145 B.n527 B.n526 10.6151
R1146 B.n526 B.n129 10.6151
R1147 B.n522 B.n129 10.6151
R1148 B.n522 B.n521 10.6151
R1149 B.n521 B.n520 10.6151
R1150 B.n520 B.n131 10.6151
R1151 B.n516 B.n131 10.6151
R1152 B.n516 B.n515 10.6151
R1153 B.n515 B.n514 10.6151
R1154 B.n514 B.n133 10.6151
R1155 B.n510 B.n133 10.6151
R1156 B.n510 B.n509 10.6151
R1157 B.n509 B.n508 10.6151
R1158 B.n508 B.n135 10.6151
R1159 B.n504 B.n135 10.6151
R1160 B.n504 B.n503 10.6151
R1161 B.n503 B.n502 10.6151
R1162 B.n502 B.n137 10.6151
R1163 B.n498 B.n137 10.6151
R1164 B.n498 B.n497 10.6151
R1165 B.n497 B.n496 10.6151
R1166 B.n496 B.n139 10.6151
R1167 B.n492 B.n139 10.6151
R1168 B.n492 B.n491 10.6151
R1169 B.n491 B.n490 10.6151
R1170 B.n490 B.n141 10.6151
R1171 B.n486 B.n141 10.6151
R1172 B.n486 B.n485 10.6151
R1173 B.n485 B.n484 10.6151
R1174 B.n484 B.n143 10.6151
R1175 B.n480 B.n143 10.6151
R1176 B.n231 B.n1 10.6151
R1177 B.n232 B.n231 10.6151
R1178 B.n232 B.n229 10.6151
R1179 B.n236 B.n229 10.6151
R1180 B.n237 B.n236 10.6151
R1181 B.n238 B.n237 10.6151
R1182 B.n238 B.n227 10.6151
R1183 B.n242 B.n227 10.6151
R1184 B.n243 B.n242 10.6151
R1185 B.n244 B.n243 10.6151
R1186 B.n244 B.n225 10.6151
R1187 B.n248 B.n225 10.6151
R1188 B.n249 B.n248 10.6151
R1189 B.n250 B.n249 10.6151
R1190 B.n250 B.n223 10.6151
R1191 B.n254 B.n223 10.6151
R1192 B.n255 B.n254 10.6151
R1193 B.n256 B.n255 10.6151
R1194 B.n256 B.n221 10.6151
R1195 B.n260 B.n221 10.6151
R1196 B.n261 B.n260 10.6151
R1197 B.n262 B.n261 10.6151
R1198 B.n262 B.n219 10.6151
R1199 B.n266 B.n219 10.6151
R1200 B.n267 B.n266 10.6151
R1201 B.n268 B.n267 10.6151
R1202 B.n268 B.n217 10.6151
R1203 B.n272 B.n217 10.6151
R1204 B.n273 B.n272 10.6151
R1205 B.n274 B.n273 10.6151
R1206 B.n274 B.n215 10.6151
R1207 B.n278 B.n215 10.6151
R1208 B.n279 B.n278 10.6151
R1209 B.n280 B.n279 10.6151
R1210 B.n280 B.n213 10.6151
R1211 B.n284 B.n213 10.6151
R1212 B.n285 B.n284 10.6151
R1213 B.n286 B.n285 10.6151
R1214 B.n286 B.n211 10.6151
R1215 B.n290 B.n211 10.6151
R1216 B.n291 B.n290 10.6151
R1217 B.n292 B.n291 10.6151
R1218 B.n292 B.n209 10.6151
R1219 B.n296 B.n209 10.6151
R1220 B.n297 B.n296 10.6151
R1221 B.n298 B.n297 10.6151
R1222 B.n298 B.n207 10.6151
R1223 B.n302 B.n207 10.6151
R1224 B.n303 B.n302 10.6151
R1225 B.n304 B.n303 10.6151
R1226 B.n304 B.n205 10.6151
R1227 B.n308 B.n205 10.6151
R1228 B.n310 B.n309 10.6151
R1229 B.n310 B.n203 10.6151
R1230 B.n314 B.n203 10.6151
R1231 B.n315 B.n314 10.6151
R1232 B.n316 B.n315 10.6151
R1233 B.n316 B.n201 10.6151
R1234 B.n320 B.n201 10.6151
R1235 B.n321 B.n320 10.6151
R1236 B.n322 B.n321 10.6151
R1237 B.n322 B.n199 10.6151
R1238 B.n326 B.n199 10.6151
R1239 B.n327 B.n326 10.6151
R1240 B.n328 B.n327 10.6151
R1241 B.n328 B.n197 10.6151
R1242 B.n332 B.n197 10.6151
R1243 B.n333 B.n332 10.6151
R1244 B.n334 B.n333 10.6151
R1245 B.n334 B.n195 10.6151
R1246 B.n338 B.n195 10.6151
R1247 B.n339 B.n338 10.6151
R1248 B.n340 B.n339 10.6151
R1249 B.n340 B.n193 10.6151
R1250 B.n344 B.n193 10.6151
R1251 B.n345 B.n344 10.6151
R1252 B.n346 B.n345 10.6151
R1253 B.n346 B.n191 10.6151
R1254 B.n350 B.n191 10.6151
R1255 B.n351 B.n350 10.6151
R1256 B.n352 B.n351 10.6151
R1257 B.n352 B.n189 10.6151
R1258 B.n356 B.n189 10.6151
R1259 B.n357 B.n356 10.6151
R1260 B.n358 B.n357 10.6151
R1261 B.n358 B.n187 10.6151
R1262 B.n362 B.n187 10.6151
R1263 B.n363 B.n362 10.6151
R1264 B.n364 B.n363 10.6151
R1265 B.n364 B.n185 10.6151
R1266 B.n368 B.n185 10.6151
R1267 B.n369 B.n368 10.6151
R1268 B.n370 B.n369 10.6151
R1269 B.n370 B.n183 10.6151
R1270 B.n374 B.n183 10.6151
R1271 B.n375 B.n374 10.6151
R1272 B.n376 B.n375 10.6151
R1273 B.n376 B.n181 10.6151
R1274 B.n380 B.n181 10.6151
R1275 B.n381 B.n380 10.6151
R1276 B.n382 B.n381 10.6151
R1277 B.n382 B.n179 10.6151
R1278 B.n386 B.n179 10.6151
R1279 B.n389 B.n388 10.6151
R1280 B.n389 B.n175 10.6151
R1281 B.n393 B.n175 10.6151
R1282 B.n394 B.n393 10.6151
R1283 B.n395 B.n394 10.6151
R1284 B.n395 B.n173 10.6151
R1285 B.n399 B.n173 10.6151
R1286 B.n400 B.n399 10.6151
R1287 B.n402 B.n169 10.6151
R1288 B.n406 B.n169 10.6151
R1289 B.n407 B.n406 10.6151
R1290 B.n408 B.n407 10.6151
R1291 B.n408 B.n167 10.6151
R1292 B.n412 B.n167 10.6151
R1293 B.n413 B.n412 10.6151
R1294 B.n414 B.n413 10.6151
R1295 B.n414 B.n165 10.6151
R1296 B.n418 B.n165 10.6151
R1297 B.n419 B.n418 10.6151
R1298 B.n420 B.n419 10.6151
R1299 B.n420 B.n163 10.6151
R1300 B.n424 B.n163 10.6151
R1301 B.n425 B.n424 10.6151
R1302 B.n426 B.n425 10.6151
R1303 B.n426 B.n161 10.6151
R1304 B.n430 B.n161 10.6151
R1305 B.n431 B.n430 10.6151
R1306 B.n432 B.n431 10.6151
R1307 B.n432 B.n159 10.6151
R1308 B.n436 B.n159 10.6151
R1309 B.n437 B.n436 10.6151
R1310 B.n438 B.n437 10.6151
R1311 B.n438 B.n157 10.6151
R1312 B.n442 B.n157 10.6151
R1313 B.n443 B.n442 10.6151
R1314 B.n444 B.n443 10.6151
R1315 B.n444 B.n155 10.6151
R1316 B.n448 B.n155 10.6151
R1317 B.n449 B.n448 10.6151
R1318 B.n450 B.n449 10.6151
R1319 B.n450 B.n153 10.6151
R1320 B.n454 B.n153 10.6151
R1321 B.n455 B.n454 10.6151
R1322 B.n456 B.n455 10.6151
R1323 B.n456 B.n151 10.6151
R1324 B.n460 B.n151 10.6151
R1325 B.n461 B.n460 10.6151
R1326 B.n462 B.n461 10.6151
R1327 B.n462 B.n149 10.6151
R1328 B.n466 B.n149 10.6151
R1329 B.n467 B.n466 10.6151
R1330 B.n468 B.n467 10.6151
R1331 B.n468 B.n147 10.6151
R1332 B.n472 B.n147 10.6151
R1333 B.n473 B.n472 10.6151
R1334 B.n474 B.n473 10.6151
R1335 B.n474 B.n145 10.6151
R1336 B.n478 B.n145 10.6151
R1337 B.n479 B.n478 10.6151
R1338 B.n893 B.n0 8.11757
R1339 B.n893 B.n1 8.11757
R1340 B.n733 B.n58 6.5566
R1341 B.n721 B.n720 6.5566
R1342 B.n388 B.n387 6.5566
R1343 B.n401 B.n400 6.5566
R1344 B.n58 B.n54 4.05904
R1345 B.n720 B.n719 4.05904
R1346 B.n387 B.n386 4.05904
R1347 B.n402 B.n401 4.05904
R1348 VP.n16 VP.n13 161.3
R1349 VP.n18 VP.n17 161.3
R1350 VP.n19 VP.n12 161.3
R1351 VP.n21 VP.n20 161.3
R1352 VP.n22 VP.n11 161.3
R1353 VP.n24 VP.n23 161.3
R1354 VP.n25 VP.n10 161.3
R1355 VP.n27 VP.n26 161.3
R1356 VP.n55 VP.n54 161.3
R1357 VP.n53 VP.n1 161.3
R1358 VP.n52 VP.n51 161.3
R1359 VP.n50 VP.n2 161.3
R1360 VP.n49 VP.n48 161.3
R1361 VP.n47 VP.n3 161.3
R1362 VP.n46 VP.n45 161.3
R1363 VP.n44 VP.n4 161.3
R1364 VP.n43 VP.n42 161.3
R1365 VP.n40 VP.n5 161.3
R1366 VP.n39 VP.n38 161.3
R1367 VP.n37 VP.n6 161.3
R1368 VP.n36 VP.n35 161.3
R1369 VP.n34 VP.n7 161.3
R1370 VP.n33 VP.n32 161.3
R1371 VP.n31 VP.n8 161.3
R1372 VP.n15 VP.t5 137.962
R1373 VP.n29 VP.t2 105.251
R1374 VP.n41 VP.t1 105.251
R1375 VP.n0 VP.t3 105.251
R1376 VP.n9 VP.t0 105.251
R1377 VP.n14 VP.t4 105.251
R1378 VP.n30 VP.n29 84.3435
R1379 VP.n56 VP.n0 84.3435
R1380 VP.n28 VP.n9 84.3435
R1381 VP.n15 VP.n14 62.4068
R1382 VP.n35 VP.n6 56.5617
R1383 VP.n48 VP.n2 56.5617
R1384 VP.n20 VP.n11 56.5617
R1385 VP.n30 VP.n28 55.0185
R1386 VP.n33 VP.n8 24.5923
R1387 VP.n34 VP.n33 24.5923
R1388 VP.n35 VP.n34 24.5923
R1389 VP.n39 VP.n6 24.5923
R1390 VP.n40 VP.n39 24.5923
R1391 VP.n42 VP.n40 24.5923
R1392 VP.n46 VP.n4 24.5923
R1393 VP.n47 VP.n46 24.5923
R1394 VP.n48 VP.n47 24.5923
R1395 VP.n52 VP.n2 24.5923
R1396 VP.n53 VP.n52 24.5923
R1397 VP.n54 VP.n53 24.5923
R1398 VP.n24 VP.n11 24.5923
R1399 VP.n25 VP.n24 24.5923
R1400 VP.n26 VP.n25 24.5923
R1401 VP.n18 VP.n13 24.5923
R1402 VP.n19 VP.n18 24.5923
R1403 VP.n20 VP.n19 24.5923
R1404 VP.n42 VP.n41 12.2964
R1405 VP.n41 VP.n4 12.2964
R1406 VP.n14 VP.n13 12.2964
R1407 VP.n29 VP.n8 5.90254
R1408 VP.n54 VP.n0 5.90254
R1409 VP.n26 VP.n9 5.90254
R1410 VP.n16 VP.n15 3.27861
R1411 VP.n28 VP.n27 0.354861
R1412 VP.n31 VP.n30 0.354861
R1413 VP.n56 VP.n55 0.354861
R1414 VP VP.n56 0.267071
R1415 VP.n17 VP.n16 0.189894
R1416 VP.n17 VP.n12 0.189894
R1417 VP.n21 VP.n12 0.189894
R1418 VP.n22 VP.n21 0.189894
R1419 VP.n23 VP.n22 0.189894
R1420 VP.n23 VP.n10 0.189894
R1421 VP.n27 VP.n10 0.189894
R1422 VP.n32 VP.n31 0.189894
R1423 VP.n32 VP.n7 0.189894
R1424 VP.n36 VP.n7 0.189894
R1425 VP.n37 VP.n36 0.189894
R1426 VP.n38 VP.n37 0.189894
R1427 VP.n38 VP.n5 0.189894
R1428 VP.n43 VP.n5 0.189894
R1429 VP.n44 VP.n43 0.189894
R1430 VP.n45 VP.n44 0.189894
R1431 VP.n45 VP.n3 0.189894
R1432 VP.n49 VP.n3 0.189894
R1433 VP.n50 VP.n49 0.189894
R1434 VP.n51 VP.n50 0.189894
R1435 VP.n51 VP.n1 0.189894
R1436 VP.n55 VP.n1 0.189894
R1437 VTAIL.n346 VTAIL.n266 756.745
R1438 VTAIL.n82 VTAIL.n2 756.745
R1439 VTAIL.n260 VTAIL.n180 756.745
R1440 VTAIL.n172 VTAIL.n92 756.745
R1441 VTAIL.n295 VTAIL.n294 585
R1442 VTAIL.n297 VTAIL.n296 585
R1443 VTAIL.n290 VTAIL.n289 585
R1444 VTAIL.n303 VTAIL.n302 585
R1445 VTAIL.n305 VTAIL.n304 585
R1446 VTAIL.n286 VTAIL.n285 585
R1447 VTAIL.n311 VTAIL.n310 585
R1448 VTAIL.n313 VTAIL.n312 585
R1449 VTAIL.n282 VTAIL.n281 585
R1450 VTAIL.n319 VTAIL.n318 585
R1451 VTAIL.n321 VTAIL.n320 585
R1452 VTAIL.n278 VTAIL.n277 585
R1453 VTAIL.n327 VTAIL.n326 585
R1454 VTAIL.n329 VTAIL.n328 585
R1455 VTAIL.n274 VTAIL.n273 585
R1456 VTAIL.n336 VTAIL.n335 585
R1457 VTAIL.n337 VTAIL.n272 585
R1458 VTAIL.n339 VTAIL.n338 585
R1459 VTAIL.n270 VTAIL.n269 585
R1460 VTAIL.n345 VTAIL.n344 585
R1461 VTAIL.n347 VTAIL.n346 585
R1462 VTAIL.n31 VTAIL.n30 585
R1463 VTAIL.n33 VTAIL.n32 585
R1464 VTAIL.n26 VTAIL.n25 585
R1465 VTAIL.n39 VTAIL.n38 585
R1466 VTAIL.n41 VTAIL.n40 585
R1467 VTAIL.n22 VTAIL.n21 585
R1468 VTAIL.n47 VTAIL.n46 585
R1469 VTAIL.n49 VTAIL.n48 585
R1470 VTAIL.n18 VTAIL.n17 585
R1471 VTAIL.n55 VTAIL.n54 585
R1472 VTAIL.n57 VTAIL.n56 585
R1473 VTAIL.n14 VTAIL.n13 585
R1474 VTAIL.n63 VTAIL.n62 585
R1475 VTAIL.n65 VTAIL.n64 585
R1476 VTAIL.n10 VTAIL.n9 585
R1477 VTAIL.n72 VTAIL.n71 585
R1478 VTAIL.n73 VTAIL.n8 585
R1479 VTAIL.n75 VTAIL.n74 585
R1480 VTAIL.n6 VTAIL.n5 585
R1481 VTAIL.n81 VTAIL.n80 585
R1482 VTAIL.n83 VTAIL.n82 585
R1483 VTAIL.n261 VTAIL.n260 585
R1484 VTAIL.n259 VTAIL.n258 585
R1485 VTAIL.n184 VTAIL.n183 585
R1486 VTAIL.n188 VTAIL.n186 585
R1487 VTAIL.n253 VTAIL.n252 585
R1488 VTAIL.n251 VTAIL.n250 585
R1489 VTAIL.n190 VTAIL.n189 585
R1490 VTAIL.n245 VTAIL.n244 585
R1491 VTAIL.n243 VTAIL.n242 585
R1492 VTAIL.n194 VTAIL.n193 585
R1493 VTAIL.n237 VTAIL.n236 585
R1494 VTAIL.n235 VTAIL.n234 585
R1495 VTAIL.n198 VTAIL.n197 585
R1496 VTAIL.n229 VTAIL.n228 585
R1497 VTAIL.n227 VTAIL.n226 585
R1498 VTAIL.n202 VTAIL.n201 585
R1499 VTAIL.n221 VTAIL.n220 585
R1500 VTAIL.n219 VTAIL.n218 585
R1501 VTAIL.n206 VTAIL.n205 585
R1502 VTAIL.n213 VTAIL.n212 585
R1503 VTAIL.n211 VTAIL.n210 585
R1504 VTAIL.n173 VTAIL.n172 585
R1505 VTAIL.n171 VTAIL.n170 585
R1506 VTAIL.n96 VTAIL.n95 585
R1507 VTAIL.n100 VTAIL.n98 585
R1508 VTAIL.n165 VTAIL.n164 585
R1509 VTAIL.n163 VTAIL.n162 585
R1510 VTAIL.n102 VTAIL.n101 585
R1511 VTAIL.n157 VTAIL.n156 585
R1512 VTAIL.n155 VTAIL.n154 585
R1513 VTAIL.n106 VTAIL.n105 585
R1514 VTAIL.n149 VTAIL.n148 585
R1515 VTAIL.n147 VTAIL.n146 585
R1516 VTAIL.n110 VTAIL.n109 585
R1517 VTAIL.n141 VTAIL.n140 585
R1518 VTAIL.n139 VTAIL.n138 585
R1519 VTAIL.n114 VTAIL.n113 585
R1520 VTAIL.n133 VTAIL.n132 585
R1521 VTAIL.n131 VTAIL.n130 585
R1522 VTAIL.n118 VTAIL.n117 585
R1523 VTAIL.n125 VTAIL.n124 585
R1524 VTAIL.n123 VTAIL.n122 585
R1525 VTAIL.n293 VTAIL.t3 327.466
R1526 VTAIL.n29 VTAIL.t7 327.466
R1527 VTAIL.n209 VTAIL.t6 327.466
R1528 VTAIL.n121 VTAIL.t0 327.466
R1529 VTAIL.n296 VTAIL.n295 171.744
R1530 VTAIL.n296 VTAIL.n289 171.744
R1531 VTAIL.n303 VTAIL.n289 171.744
R1532 VTAIL.n304 VTAIL.n303 171.744
R1533 VTAIL.n304 VTAIL.n285 171.744
R1534 VTAIL.n311 VTAIL.n285 171.744
R1535 VTAIL.n312 VTAIL.n311 171.744
R1536 VTAIL.n312 VTAIL.n281 171.744
R1537 VTAIL.n319 VTAIL.n281 171.744
R1538 VTAIL.n320 VTAIL.n319 171.744
R1539 VTAIL.n320 VTAIL.n277 171.744
R1540 VTAIL.n327 VTAIL.n277 171.744
R1541 VTAIL.n328 VTAIL.n327 171.744
R1542 VTAIL.n328 VTAIL.n273 171.744
R1543 VTAIL.n336 VTAIL.n273 171.744
R1544 VTAIL.n337 VTAIL.n336 171.744
R1545 VTAIL.n338 VTAIL.n337 171.744
R1546 VTAIL.n338 VTAIL.n269 171.744
R1547 VTAIL.n345 VTAIL.n269 171.744
R1548 VTAIL.n346 VTAIL.n345 171.744
R1549 VTAIL.n32 VTAIL.n31 171.744
R1550 VTAIL.n32 VTAIL.n25 171.744
R1551 VTAIL.n39 VTAIL.n25 171.744
R1552 VTAIL.n40 VTAIL.n39 171.744
R1553 VTAIL.n40 VTAIL.n21 171.744
R1554 VTAIL.n47 VTAIL.n21 171.744
R1555 VTAIL.n48 VTAIL.n47 171.744
R1556 VTAIL.n48 VTAIL.n17 171.744
R1557 VTAIL.n55 VTAIL.n17 171.744
R1558 VTAIL.n56 VTAIL.n55 171.744
R1559 VTAIL.n56 VTAIL.n13 171.744
R1560 VTAIL.n63 VTAIL.n13 171.744
R1561 VTAIL.n64 VTAIL.n63 171.744
R1562 VTAIL.n64 VTAIL.n9 171.744
R1563 VTAIL.n72 VTAIL.n9 171.744
R1564 VTAIL.n73 VTAIL.n72 171.744
R1565 VTAIL.n74 VTAIL.n73 171.744
R1566 VTAIL.n74 VTAIL.n5 171.744
R1567 VTAIL.n81 VTAIL.n5 171.744
R1568 VTAIL.n82 VTAIL.n81 171.744
R1569 VTAIL.n260 VTAIL.n259 171.744
R1570 VTAIL.n259 VTAIL.n183 171.744
R1571 VTAIL.n188 VTAIL.n183 171.744
R1572 VTAIL.n252 VTAIL.n188 171.744
R1573 VTAIL.n252 VTAIL.n251 171.744
R1574 VTAIL.n251 VTAIL.n189 171.744
R1575 VTAIL.n244 VTAIL.n189 171.744
R1576 VTAIL.n244 VTAIL.n243 171.744
R1577 VTAIL.n243 VTAIL.n193 171.744
R1578 VTAIL.n236 VTAIL.n193 171.744
R1579 VTAIL.n236 VTAIL.n235 171.744
R1580 VTAIL.n235 VTAIL.n197 171.744
R1581 VTAIL.n228 VTAIL.n197 171.744
R1582 VTAIL.n228 VTAIL.n227 171.744
R1583 VTAIL.n227 VTAIL.n201 171.744
R1584 VTAIL.n220 VTAIL.n201 171.744
R1585 VTAIL.n220 VTAIL.n219 171.744
R1586 VTAIL.n219 VTAIL.n205 171.744
R1587 VTAIL.n212 VTAIL.n205 171.744
R1588 VTAIL.n212 VTAIL.n211 171.744
R1589 VTAIL.n172 VTAIL.n171 171.744
R1590 VTAIL.n171 VTAIL.n95 171.744
R1591 VTAIL.n100 VTAIL.n95 171.744
R1592 VTAIL.n164 VTAIL.n100 171.744
R1593 VTAIL.n164 VTAIL.n163 171.744
R1594 VTAIL.n163 VTAIL.n101 171.744
R1595 VTAIL.n156 VTAIL.n101 171.744
R1596 VTAIL.n156 VTAIL.n155 171.744
R1597 VTAIL.n155 VTAIL.n105 171.744
R1598 VTAIL.n148 VTAIL.n105 171.744
R1599 VTAIL.n148 VTAIL.n147 171.744
R1600 VTAIL.n147 VTAIL.n109 171.744
R1601 VTAIL.n140 VTAIL.n109 171.744
R1602 VTAIL.n140 VTAIL.n139 171.744
R1603 VTAIL.n139 VTAIL.n113 171.744
R1604 VTAIL.n132 VTAIL.n113 171.744
R1605 VTAIL.n132 VTAIL.n131 171.744
R1606 VTAIL.n131 VTAIL.n117 171.744
R1607 VTAIL.n124 VTAIL.n117 171.744
R1608 VTAIL.n124 VTAIL.n123 171.744
R1609 VTAIL.n295 VTAIL.t3 85.8723
R1610 VTAIL.n31 VTAIL.t7 85.8723
R1611 VTAIL.n211 VTAIL.t6 85.8723
R1612 VTAIL.n123 VTAIL.t0 85.8723
R1613 VTAIL.n179 VTAIL.n178 55.5188
R1614 VTAIL.n91 VTAIL.n90 55.5188
R1615 VTAIL.n1 VTAIL.n0 55.5186
R1616 VTAIL.n89 VTAIL.n88 55.5186
R1617 VTAIL.n351 VTAIL.n350 34.1247
R1618 VTAIL.n87 VTAIL.n86 34.1247
R1619 VTAIL.n265 VTAIL.n264 34.1247
R1620 VTAIL.n177 VTAIL.n176 34.1247
R1621 VTAIL.n91 VTAIL.n89 32.3669
R1622 VTAIL.n351 VTAIL.n265 29.0307
R1623 VTAIL.n294 VTAIL.n293 16.3895
R1624 VTAIL.n30 VTAIL.n29 16.3895
R1625 VTAIL.n210 VTAIL.n209 16.3895
R1626 VTAIL.n122 VTAIL.n121 16.3895
R1627 VTAIL.n339 VTAIL.n270 13.1884
R1628 VTAIL.n75 VTAIL.n6 13.1884
R1629 VTAIL.n186 VTAIL.n184 13.1884
R1630 VTAIL.n98 VTAIL.n96 13.1884
R1631 VTAIL.n297 VTAIL.n292 12.8005
R1632 VTAIL.n340 VTAIL.n272 12.8005
R1633 VTAIL.n344 VTAIL.n343 12.8005
R1634 VTAIL.n33 VTAIL.n28 12.8005
R1635 VTAIL.n76 VTAIL.n8 12.8005
R1636 VTAIL.n80 VTAIL.n79 12.8005
R1637 VTAIL.n258 VTAIL.n257 12.8005
R1638 VTAIL.n254 VTAIL.n253 12.8005
R1639 VTAIL.n213 VTAIL.n208 12.8005
R1640 VTAIL.n170 VTAIL.n169 12.8005
R1641 VTAIL.n166 VTAIL.n165 12.8005
R1642 VTAIL.n125 VTAIL.n120 12.8005
R1643 VTAIL.n298 VTAIL.n290 12.0247
R1644 VTAIL.n335 VTAIL.n334 12.0247
R1645 VTAIL.n347 VTAIL.n268 12.0247
R1646 VTAIL.n34 VTAIL.n26 12.0247
R1647 VTAIL.n71 VTAIL.n70 12.0247
R1648 VTAIL.n83 VTAIL.n4 12.0247
R1649 VTAIL.n261 VTAIL.n182 12.0247
R1650 VTAIL.n250 VTAIL.n187 12.0247
R1651 VTAIL.n214 VTAIL.n206 12.0247
R1652 VTAIL.n173 VTAIL.n94 12.0247
R1653 VTAIL.n162 VTAIL.n99 12.0247
R1654 VTAIL.n126 VTAIL.n118 12.0247
R1655 VTAIL.n302 VTAIL.n301 11.249
R1656 VTAIL.n333 VTAIL.n274 11.249
R1657 VTAIL.n348 VTAIL.n266 11.249
R1658 VTAIL.n38 VTAIL.n37 11.249
R1659 VTAIL.n69 VTAIL.n10 11.249
R1660 VTAIL.n84 VTAIL.n2 11.249
R1661 VTAIL.n262 VTAIL.n180 11.249
R1662 VTAIL.n249 VTAIL.n190 11.249
R1663 VTAIL.n218 VTAIL.n217 11.249
R1664 VTAIL.n174 VTAIL.n92 11.249
R1665 VTAIL.n161 VTAIL.n102 11.249
R1666 VTAIL.n130 VTAIL.n129 11.249
R1667 VTAIL.n305 VTAIL.n288 10.4732
R1668 VTAIL.n330 VTAIL.n329 10.4732
R1669 VTAIL.n41 VTAIL.n24 10.4732
R1670 VTAIL.n66 VTAIL.n65 10.4732
R1671 VTAIL.n246 VTAIL.n245 10.4732
R1672 VTAIL.n221 VTAIL.n204 10.4732
R1673 VTAIL.n158 VTAIL.n157 10.4732
R1674 VTAIL.n133 VTAIL.n116 10.4732
R1675 VTAIL.n306 VTAIL.n286 9.69747
R1676 VTAIL.n326 VTAIL.n276 9.69747
R1677 VTAIL.n42 VTAIL.n22 9.69747
R1678 VTAIL.n62 VTAIL.n12 9.69747
R1679 VTAIL.n242 VTAIL.n192 9.69747
R1680 VTAIL.n222 VTAIL.n202 9.69747
R1681 VTAIL.n154 VTAIL.n104 9.69747
R1682 VTAIL.n134 VTAIL.n114 9.69747
R1683 VTAIL.n350 VTAIL.n349 9.45567
R1684 VTAIL.n86 VTAIL.n85 9.45567
R1685 VTAIL.n264 VTAIL.n263 9.45567
R1686 VTAIL.n176 VTAIL.n175 9.45567
R1687 VTAIL.n349 VTAIL.n348 9.3005
R1688 VTAIL.n268 VTAIL.n267 9.3005
R1689 VTAIL.n343 VTAIL.n342 9.3005
R1690 VTAIL.n315 VTAIL.n314 9.3005
R1691 VTAIL.n284 VTAIL.n283 9.3005
R1692 VTAIL.n309 VTAIL.n308 9.3005
R1693 VTAIL.n307 VTAIL.n306 9.3005
R1694 VTAIL.n288 VTAIL.n287 9.3005
R1695 VTAIL.n301 VTAIL.n300 9.3005
R1696 VTAIL.n299 VTAIL.n298 9.3005
R1697 VTAIL.n292 VTAIL.n291 9.3005
R1698 VTAIL.n317 VTAIL.n316 9.3005
R1699 VTAIL.n280 VTAIL.n279 9.3005
R1700 VTAIL.n323 VTAIL.n322 9.3005
R1701 VTAIL.n325 VTAIL.n324 9.3005
R1702 VTAIL.n276 VTAIL.n275 9.3005
R1703 VTAIL.n331 VTAIL.n330 9.3005
R1704 VTAIL.n333 VTAIL.n332 9.3005
R1705 VTAIL.n334 VTAIL.n271 9.3005
R1706 VTAIL.n341 VTAIL.n340 9.3005
R1707 VTAIL.n85 VTAIL.n84 9.3005
R1708 VTAIL.n4 VTAIL.n3 9.3005
R1709 VTAIL.n79 VTAIL.n78 9.3005
R1710 VTAIL.n51 VTAIL.n50 9.3005
R1711 VTAIL.n20 VTAIL.n19 9.3005
R1712 VTAIL.n45 VTAIL.n44 9.3005
R1713 VTAIL.n43 VTAIL.n42 9.3005
R1714 VTAIL.n24 VTAIL.n23 9.3005
R1715 VTAIL.n37 VTAIL.n36 9.3005
R1716 VTAIL.n35 VTAIL.n34 9.3005
R1717 VTAIL.n28 VTAIL.n27 9.3005
R1718 VTAIL.n53 VTAIL.n52 9.3005
R1719 VTAIL.n16 VTAIL.n15 9.3005
R1720 VTAIL.n59 VTAIL.n58 9.3005
R1721 VTAIL.n61 VTAIL.n60 9.3005
R1722 VTAIL.n12 VTAIL.n11 9.3005
R1723 VTAIL.n67 VTAIL.n66 9.3005
R1724 VTAIL.n69 VTAIL.n68 9.3005
R1725 VTAIL.n70 VTAIL.n7 9.3005
R1726 VTAIL.n77 VTAIL.n76 9.3005
R1727 VTAIL.n196 VTAIL.n195 9.3005
R1728 VTAIL.n239 VTAIL.n238 9.3005
R1729 VTAIL.n241 VTAIL.n240 9.3005
R1730 VTAIL.n192 VTAIL.n191 9.3005
R1731 VTAIL.n247 VTAIL.n246 9.3005
R1732 VTAIL.n249 VTAIL.n248 9.3005
R1733 VTAIL.n187 VTAIL.n185 9.3005
R1734 VTAIL.n255 VTAIL.n254 9.3005
R1735 VTAIL.n263 VTAIL.n262 9.3005
R1736 VTAIL.n182 VTAIL.n181 9.3005
R1737 VTAIL.n257 VTAIL.n256 9.3005
R1738 VTAIL.n233 VTAIL.n232 9.3005
R1739 VTAIL.n231 VTAIL.n230 9.3005
R1740 VTAIL.n200 VTAIL.n199 9.3005
R1741 VTAIL.n225 VTAIL.n224 9.3005
R1742 VTAIL.n223 VTAIL.n222 9.3005
R1743 VTAIL.n204 VTAIL.n203 9.3005
R1744 VTAIL.n217 VTAIL.n216 9.3005
R1745 VTAIL.n215 VTAIL.n214 9.3005
R1746 VTAIL.n208 VTAIL.n207 9.3005
R1747 VTAIL.n108 VTAIL.n107 9.3005
R1748 VTAIL.n151 VTAIL.n150 9.3005
R1749 VTAIL.n153 VTAIL.n152 9.3005
R1750 VTAIL.n104 VTAIL.n103 9.3005
R1751 VTAIL.n159 VTAIL.n158 9.3005
R1752 VTAIL.n161 VTAIL.n160 9.3005
R1753 VTAIL.n99 VTAIL.n97 9.3005
R1754 VTAIL.n167 VTAIL.n166 9.3005
R1755 VTAIL.n175 VTAIL.n174 9.3005
R1756 VTAIL.n94 VTAIL.n93 9.3005
R1757 VTAIL.n169 VTAIL.n168 9.3005
R1758 VTAIL.n145 VTAIL.n144 9.3005
R1759 VTAIL.n143 VTAIL.n142 9.3005
R1760 VTAIL.n112 VTAIL.n111 9.3005
R1761 VTAIL.n137 VTAIL.n136 9.3005
R1762 VTAIL.n135 VTAIL.n134 9.3005
R1763 VTAIL.n116 VTAIL.n115 9.3005
R1764 VTAIL.n129 VTAIL.n128 9.3005
R1765 VTAIL.n127 VTAIL.n126 9.3005
R1766 VTAIL.n120 VTAIL.n119 9.3005
R1767 VTAIL.n310 VTAIL.n309 8.92171
R1768 VTAIL.n325 VTAIL.n278 8.92171
R1769 VTAIL.n46 VTAIL.n45 8.92171
R1770 VTAIL.n61 VTAIL.n14 8.92171
R1771 VTAIL.n241 VTAIL.n194 8.92171
R1772 VTAIL.n226 VTAIL.n225 8.92171
R1773 VTAIL.n153 VTAIL.n106 8.92171
R1774 VTAIL.n138 VTAIL.n137 8.92171
R1775 VTAIL.n313 VTAIL.n284 8.14595
R1776 VTAIL.n322 VTAIL.n321 8.14595
R1777 VTAIL.n49 VTAIL.n20 8.14595
R1778 VTAIL.n58 VTAIL.n57 8.14595
R1779 VTAIL.n238 VTAIL.n237 8.14595
R1780 VTAIL.n229 VTAIL.n200 8.14595
R1781 VTAIL.n150 VTAIL.n149 8.14595
R1782 VTAIL.n141 VTAIL.n112 8.14595
R1783 VTAIL.n314 VTAIL.n282 7.3702
R1784 VTAIL.n318 VTAIL.n280 7.3702
R1785 VTAIL.n50 VTAIL.n18 7.3702
R1786 VTAIL.n54 VTAIL.n16 7.3702
R1787 VTAIL.n234 VTAIL.n196 7.3702
R1788 VTAIL.n230 VTAIL.n198 7.3702
R1789 VTAIL.n146 VTAIL.n108 7.3702
R1790 VTAIL.n142 VTAIL.n110 7.3702
R1791 VTAIL.n317 VTAIL.n282 6.59444
R1792 VTAIL.n318 VTAIL.n317 6.59444
R1793 VTAIL.n53 VTAIL.n18 6.59444
R1794 VTAIL.n54 VTAIL.n53 6.59444
R1795 VTAIL.n234 VTAIL.n233 6.59444
R1796 VTAIL.n233 VTAIL.n198 6.59444
R1797 VTAIL.n146 VTAIL.n145 6.59444
R1798 VTAIL.n145 VTAIL.n110 6.59444
R1799 VTAIL.n314 VTAIL.n313 5.81868
R1800 VTAIL.n321 VTAIL.n280 5.81868
R1801 VTAIL.n50 VTAIL.n49 5.81868
R1802 VTAIL.n57 VTAIL.n16 5.81868
R1803 VTAIL.n237 VTAIL.n196 5.81868
R1804 VTAIL.n230 VTAIL.n229 5.81868
R1805 VTAIL.n149 VTAIL.n108 5.81868
R1806 VTAIL.n142 VTAIL.n141 5.81868
R1807 VTAIL.n310 VTAIL.n284 5.04292
R1808 VTAIL.n322 VTAIL.n278 5.04292
R1809 VTAIL.n46 VTAIL.n20 5.04292
R1810 VTAIL.n58 VTAIL.n14 5.04292
R1811 VTAIL.n238 VTAIL.n194 5.04292
R1812 VTAIL.n226 VTAIL.n200 5.04292
R1813 VTAIL.n150 VTAIL.n106 5.04292
R1814 VTAIL.n138 VTAIL.n112 5.04292
R1815 VTAIL.n309 VTAIL.n286 4.26717
R1816 VTAIL.n326 VTAIL.n325 4.26717
R1817 VTAIL.n45 VTAIL.n22 4.26717
R1818 VTAIL.n62 VTAIL.n61 4.26717
R1819 VTAIL.n242 VTAIL.n241 4.26717
R1820 VTAIL.n225 VTAIL.n202 4.26717
R1821 VTAIL.n154 VTAIL.n153 4.26717
R1822 VTAIL.n137 VTAIL.n114 4.26717
R1823 VTAIL.n293 VTAIL.n291 3.70982
R1824 VTAIL.n29 VTAIL.n27 3.70982
R1825 VTAIL.n209 VTAIL.n207 3.70982
R1826 VTAIL.n121 VTAIL.n119 3.70982
R1827 VTAIL.n306 VTAIL.n305 3.49141
R1828 VTAIL.n329 VTAIL.n276 3.49141
R1829 VTAIL.n42 VTAIL.n41 3.49141
R1830 VTAIL.n65 VTAIL.n12 3.49141
R1831 VTAIL.n245 VTAIL.n192 3.49141
R1832 VTAIL.n222 VTAIL.n221 3.49141
R1833 VTAIL.n157 VTAIL.n104 3.49141
R1834 VTAIL.n134 VTAIL.n133 3.49141
R1835 VTAIL.n177 VTAIL.n91 3.33671
R1836 VTAIL.n265 VTAIL.n179 3.33671
R1837 VTAIL.n89 VTAIL.n87 3.33671
R1838 VTAIL.n302 VTAIL.n288 2.71565
R1839 VTAIL.n330 VTAIL.n274 2.71565
R1840 VTAIL.n350 VTAIL.n266 2.71565
R1841 VTAIL.n38 VTAIL.n24 2.71565
R1842 VTAIL.n66 VTAIL.n10 2.71565
R1843 VTAIL.n86 VTAIL.n2 2.71565
R1844 VTAIL.n264 VTAIL.n180 2.71565
R1845 VTAIL.n246 VTAIL.n190 2.71565
R1846 VTAIL.n218 VTAIL.n204 2.71565
R1847 VTAIL.n176 VTAIL.n92 2.71565
R1848 VTAIL.n158 VTAIL.n102 2.71565
R1849 VTAIL.n130 VTAIL.n116 2.71565
R1850 VTAIL VTAIL.n351 2.44447
R1851 VTAIL.n179 VTAIL.n177 2.13843
R1852 VTAIL.n87 VTAIL.n1 2.13843
R1853 VTAIL.n0 VTAIL.t4 2.10302
R1854 VTAIL.n0 VTAIL.t1 2.10302
R1855 VTAIL.n88 VTAIL.t8 2.10302
R1856 VTAIL.n88 VTAIL.t10 2.10302
R1857 VTAIL.n178 VTAIL.t9 2.10302
R1858 VTAIL.n178 VTAIL.t11 2.10302
R1859 VTAIL.n90 VTAIL.t5 2.10302
R1860 VTAIL.n90 VTAIL.t2 2.10302
R1861 VTAIL.n301 VTAIL.n290 1.93989
R1862 VTAIL.n335 VTAIL.n333 1.93989
R1863 VTAIL.n348 VTAIL.n347 1.93989
R1864 VTAIL.n37 VTAIL.n26 1.93989
R1865 VTAIL.n71 VTAIL.n69 1.93989
R1866 VTAIL.n84 VTAIL.n83 1.93989
R1867 VTAIL.n262 VTAIL.n261 1.93989
R1868 VTAIL.n250 VTAIL.n249 1.93989
R1869 VTAIL.n217 VTAIL.n206 1.93989
R1870 VTAIL.n174 VTAIL.n173 1.93989
R1871 VTAIL.n162 VTAIL.n161 1.93989
R1872 VTAIL.n129 VTAIL.n118 1.93989
R1873 VTAIL.n298 VTAIL.n297 1.16414
R1874 VTAIL.n334 VTAIL.n272 1.16414
R1875 VTAIL.n344 VTAIL.n268 1.16414
R1876 VTAIL.n34 VTAIL.n33 1.16414
R1877 VTAIL.n70 VTAIL.n8 1.16414
R1878 VTAIL.n80 VTAIL.n4 1.16414
R1879 VTAIL.n258 VTAIL.n182 1.16414
R1880 VTAIL.n253 VTAIL.n187 1.16414
R1881 VTAIL.n214 VTAIL.n213 1.16414
R1882 VTAIL.n170 VTAIL.n94 1.16414
R1883 VTAIL.n165 VTAIL.n99 1.16414
R1884 VTAIL.n126 VTAIL.n125 1.16414
R1885 VTAIL VTAIL.n1 0.892741
R1886 VTAIL.n294 VTAIL.n292 0.388379
R1887 VTAIL.n340 VTAIL.n339 0.388379
R1888 VTAIL.n343 VTAIL.n270 0.388379
R1889 VTAIL.n30 VTAIL.n28 0.388379
R1890 VTAIL.n76 VTAIL.n75 0.388379
R1891 VTAIL.n79 VTAIL.n6 0.388379
R1892 VTAIL.n257 VTAIL.n184 0.388379
R1893 VTAIL.n254 VTAIL.n186 0.388379
R1894 VTAIL.n210 VTAIL.n208 0.388379
R1895 VTAIL.n169 VTAIL.n96 0.388379
R1896 VTAIL.n166 VTAIL.n98 0.388379
R1897 VTAIL.n122 VTAIL.n120 0.388379
R1898 VTAIL.n299 VTAIL.n291 0.155672
R1899 VTAIL.n300 VTAIL.n299 0.155672
R1900 VTAIL.n300 VTAIL.n287 0.155672
R1901 VTAIL.n307 VTAIL.n287 0.155672
R1902 VTAIL.n308 VTAIL.n307 0.155672
R1903 VTAIL.n308 VTAIL.n283 0.155672
R1904 VTAIL.n315 VTAIL.n283 0.155672
R1905 VTAIL.n316 VTAIL.n315 0.155672
R1906 VTAIL.n316 VTAIL.n279 0.155672
R1907 VTAIL.n323 VTAIL.n279 0.155672
R1908 VTAIL.n324 VTAIL.n323 0.155672
R1909 VTAIL.n324 VTAIL.n275 0.155672
R1910 VTAIL.n331 VTAIL.n275 0.155672
R1911 VTAIL.n332 VTAIL.n331 0.155672
R1912 VTAIL.n332 VTAIL.n271 0.155672
R1913 VTAIL.n341 VTAIL.n271 0.155672
R1914 VTAIL.n342 VTAIL.n341 0.155672
R1915 VTAIL.n342 VTAIL.n267 0.155672
R1916 VTAIL.n349 VTAIL.n267 0.155672
R1917 VTAIL.n35 VTAIL.n27 0.155672
R1918 VTAIL.n36 VTAIL.n35 0.155672
R1919 VTAIL.n36 VTAIL.n23 0.155672
R1920 VTAIL.n43 VTAIL.n23 0.155672
R1921 VTAIL.n44 VTAIL.n43 0.155672
R1922 VTAIL.n44 VTAIL.n19 0.155672
R1923 VTAIL.n51 VTAIL.n19 0.155672
R1924 VTAIL.n52 VTAIL.n51 0.155672
R1925 VTAIL.n52 VTAIL.n15 0.155672
R1926 VTAIL.n59 VTAIL.n15 0.155672
R1927 VTAIL.n60 VTAIL.n59 0.155672
R1928 VTAIL.n60 VTAIL.n11 0.155672
R1929 VTAIL.n67 VTAIL.n11 0.155672
R1930 VTAIL.n68 VTAIL.n67 0.155672
R1931 VTAIL.n68 VTAIL.n7 0.155672
R1932 VTAIL.n77 VTAIL.n7 0.155672
R1933 VTAIL.n78 VTAIL.n77 0.155672
R1934 VTAIL.n78 VTAIL.n3 0.155672
R1935 VTAIL.n85 VTAIL.n3 0.155672
R1936 VTAIL.n263 VTAIL.n181 0.155672
R1937 VTAIL.n256 VTAIL.n181 0.155672
R1938 VTAIL.n256 VTAIL.n255 0.155672
R1939 VTAIL.n255 VTAIL.n185 0.155672
R1940 VTAIL.n248 VTAIL.n185 0.155672
R1941 VTAIL.n248 VTAIL.n247 0.155672
R1942 VTAIL.n247 VTAIL.n191 0.155672
R1943 VTAIL.n240 VTAIL.n191 0.155672
R1944 VTAIL.n240 VTAIL.n239 0.155672
R1945 VTAIL.n239 VTAIL.n195 0.155672
R1946 VTAIL.n232 VTAIL.n195 0.155672
R1947 VTAIL.n232 VTAIL.n231 0.155672
R1948 VTAIL.n231 VTAIL.n199 0.155672
R1949 VTAIL.n224 VTAIL.n199 0.155672
R1950 VTAIL.n224 VTAIL.n223 0.155672
R1951 VTAIL.n223 VTAIL.n203 0.155672
R1952 VTAIL.n216 VTAIL.n203 0.155672
R1953 VTAIL.n216 VTAIL.n215 0.155672
R1954 VTAIL.n215 VTAIL.n207 0.155672
R1955 VTAIL.n175 VTAIL.n93 0.155672
R1956 VTAIL.n168 VTAIL.n93 0.155672
R1957 VTAIL.n168 VTAIL.n167 0.155672
R1958 VTAIL.n167 VTAIL.n97 0.155672
R1959 VTAIL.n160 VTAIL.n97 0.155672
R1960 VTAIL.n160 VTAIL.n159 0.155672
R1961 VTAIL.n159 VTAIL.n103 0.155672
R1962 VTAIL.n152 VTAIL.n103 0.155672
R1963 VTAIL.n152 VTAIL.n151 0.155672
R1964 VTAIL.n151 VTAIL.n107 0.155672
R1965 VTAIL.n144 VTAIL.n107 0.155672
R1966 VTAIL.n144 VTAIL.n143 0.155672
R1967 VTAIL.n143 VTAIL.n111 0.155672
R1968 VTAIL.n136 VTAIL.n111 0.155672
R1969 VTAIL.n136 VTAIL.n135 0.155672
R1970 VTAIL.n135 VTAIL.n115 0.155672
R1971 VTAIL.n128 VTAIL.n115 0.155672
R1972 VTAIL.n128 VTAIL.n127 0.155672
R1973 VTAIL.n127 VTAIL.n119 0.155672
R1974 VDD1.n80 VDD1.n0 756.745
R1975 VDD1.n165 VDD1.n85 756.745
R1976 VDD1.n81 VDD1.n80 585
R1977 VDD1.n79 VDD1.n78 585
R1978 VDD1.n4 VDD1.n3 585
R1979 VDD1.n8 VDD1.n6 585
R1980 VDD1.n73 VDD1.n72 585
R1981 VDD1.n71 VDD1.n70 585
R1982 VDD1.n10 VDD1.n9 585
R1983 VDD1.n65 VDD1.n64 585
R1984 VDD1.n63 VDD1.n62 585
R1985 VDD1.n14 VDD1.n13 585
R1986 VDD1.n57 VDD1.n56 585
R1987 VDD1.n55 VDD1.n54 585
R1988 VDD1.n18 VDD1.n17 585
R1989 VDD1.n49 VDD1.n48 585
R1990 VDD1.n47 VDD1.n46 585
R1991 VDD1.n22 VDD1.n21 585
R1992 VDD1.n41 VDD1.n40 585
R1993 VDD1.n39 VDD1.n38 585
R1994 VDD1.n26 VDD1.n25 585
R1995 VDD1.n33 VDD1.n32 585
R1996 VDD1.n31 VDD1.n30 585
R1997 VDD1.n114 VDD1.n113 585
R1998 VDD1.n116 VDD1.n115 585
R1999 VDD1.n109 VDD1.n108 585
R2000 VDD1.n122 VDD1.n121 585
R2001 VDD1.n124 VDD1.n123 585
R2002 VDD1.n105 VDD1.n104 585
R2003 VDD1.n130 VDD1.n129 585
R2004 VDD1.n132 VDD1.n131 585
R2005 VDD1.n101 VDD1.n100 585
R2006 VDD1.n138 VDD1.n137 585
R2007 VDD1.n140 VDD1.n139 585
R2008 VDD1.n97 VDD1.n96 585
R2009 VDD1.n146 VDD1.n145 585
R2010 VDD1.n148 VDD1.n147 585
R2011 VDD1.n93 VDD1.n92 585
R2012 VDD1.n155 VDD1.n154 585
R2013 VDD1.n156 VDD1.n91 585
R2014 VDD1.n158 VDD1.n157 585
R2015 VDD1.n89 VDD1.n88 585
R2016 VDD1.n164 VDD1.n163 585
R2017 VDD1.n166 VDD1.n165 585
R2018 VDD1.n29 VDD1.t0 327.466
R2019 VDD1.n112 VDD1.t3 327.466
R2020 VDD1.n80 VDD1.n79 171.744
R2021 VDD1.n79 VDD1.n3 171.744
R2022 VDD1.n8 VDD1.n3 171.744
R2023 VDD1.n72 VDD1.n8 171.744
R2024 VDD1.n72 VDD1.n71 171.744
R2025 VDD1.n71 VDD1.n9 171.744
R2026 VDD1.n64 VDD1.n9 171.744
R2027 VDD1.n64 VDD1.n63 171.744
R2028 VDD1.n63 VDD1.n13 171.744
R2029 VDD1.n56 VDD1.n13 171.744
R2030 VDD1.n56 VDD1.n55 171.744
R2031 VDD1.n55 VDD1.n17 171.744
R2032 VDD1.n48 VDD1.n17 171.744
R2033 VDD1.n48 VDD1.n47 171.744
R2034 VDD1.n47 VDD1.n21 171.744
R2035 VDD1.n40 VDD1.n21 171.744
R2036 VDD1.n40 VDD1.n39 171.744
R2037 VDD1.n39 VDD1.n25 171.744
R2038 VDD1.n32 VDD1.n25 171.744
R2039 VDD1.n32 VDD1.n31 171.744
R2040 VDD1.n115 VDD1.n114 171.744
R2041 VDD1.n115 VDD1.n108 171.744
R2042 VDD1.n122 VDD1.n108 171.744
R2043 VDD1.n123 VDD1.n122 171.744
R2044 VDD1.n123 VDD1.n104 171.744
R2045 VDD1.n130 VDD1.n104 171.744
R2046 VDD1.n131 VDD1.n130 171.744
R2047 VDD1.n131 VDD1.n100 171.744
R2048 VDD1.n138 VDD1.n100 171.744
R2049 VDD1.n139 VDD1.n138 171.744
R2050 VDD1.n139 VDD1.n96 171.744
R2051 VDD1.n146 VDD1.n96 171.744
R2052 VDD1.n147 VDD1.n146 171.744
R2053 VDD1.n147 VDD1.n92 171.744
R2054 VDD1.n155 VDD1.n92 171.744
R2055 VDD1.n156 VDD1.n155 171.744
R2056 VDD1.n157 VDD1.n156 171.744
R2057 VDD1.n157 VDD1.n88 171.744
R2058 VDD1.n164 VDD1.n88 171.744
R2059 VDD1.n165 VDD1.n164 171.744
R2060 VDD1.n31 VDD1.t0 85.8723
R2061 VDD1.n114 VDD1.t3 85.8723
R2062 VDD1.n171 VDD1.n170 72.9761
R2063 VDD1.n173 VDD1.n172 72.1974
R2064 VDD1 VDD1.n84 53.3639
R2065 VDD1.n171 VDD1.n169 53.2503
R2066 VDD1.n173 VDD1.n171 50.1367
R2067 VDD1.n30 VDD1.n29 16.3895
R2068 VDD1.n113 VDD1.n112 16.3895
R2069 VDD1.n6 VDD1.n4 13.1884
R2070 VDD1.n158 VDD1.n89 13.1884
R2071 VDD1.n78 VDD1.n77 12.8005
R2072 VDD1.n74 VDD1.n73 12.8005
R2073 VDD1.n33 VDD1.n28 12.8005
R2074 VDD1.n116 VDD1.n111 12.8005
R2075 VDD1.n159 VDD1.n91 12.8005
R2076 VDD1.n163 VDD1.n162 12.8005
R2077 VDD1.n81 VDD1.n2 12.0247
R2078 VDD1.n70 VDD1.n7 12.0247
R2079 VDD1.n34 VDD1.n26 12.0247
R2080 VDD1.n117 VDD1.n109 12.0247
R2081 VDD1.n154 VDD1.n153 12.0247
R2082 VDD1.n166 VDD1.n87 12.0247
R2083 VDD1.n82 VDD1.n0 11.249
R2084 VDD1.n69 VDD1.n10 11.249
R2085 VDD1.n38 VDD1.n37 11.249
R2086 VDD1.n121 VDD1.n120 11.249
R2087 VDD1.n152 VDD1.n93 11.249
R2088 VDD1.n167 VDD1.n85 11.249
R2089 VDD1.n66 VDD1.n65 10.4732
R2090 VDD1.n41 VDD1.n24 10.4732
R2091 VDD1.n124 VDD1.n107 10.4732
R2092 VDD1.n149 VDD1.n148 10.4732
R2093 VDD1.n62 VDD1.n12 9.69747
R2094 VDD1.n42 VDD1.n22 9.69747
R2095 VDD1.n125 VDD1.n105 9.69747
R2096 VDD1.n145 VDD1.n95 9.69747
R2097 VDD1.n84 VDD1.n83 9.45567
R2098 VDD1.n169 VDD1.n168 9.45567
R2099 VDD1.n16 VDD1.n15 9.3005
R2100 VDD1.n59 VDD1.n58 9.3005
R2101 VDD1.n61 VDD1.n60 9.3005
R2102 VDD1.n12 VDD1.n11 9.3005
R2103 VDD1.n67 VDD1.n66 9.3005
R2104 VDD1.n69 VDD1.n68 9.3005
R2105 VDD1.n7 VDD1.n5 9.3005
R2106 VDD1.n75 VDD1.n74 9.3005
R2107 VDD1.n83 VDD1.n82 9.3005
R2108 VDD1.n2 VDD1.n1 9.3005
R2109 VDD1.n77 VDD1.n76 9.3005
R2110 VDD1.n53 VDD1.n52 9.3005
R2111 VDD1.n51 VDD1.n50 9.3005
R2112 VDD1.n20 VDD1.n19 9.3005
R2113 VDD1.n45 VDD1.n44 9.3005
R2114 VDD1.n43 VDD1.n42 9.3005
R2115 VDD1.n24 VDD1.n23 9.3005
R2116 VDD1.n37 VDD1.n36 9.3005
R2117 VDD1.n35 VDD1.n34 9.3005
R2118 VDD1.n28 VDD1.n27 9.3005
R2119 VDD1.n168 VDD1.n167 9.3005
R2120 VDD1.n87 VDD1.n86 9.3005
R2121 VDD1.n162 VDD1.n161 9.3005
R2122 VDD1.n134 VDD1.n133 9.3005
R2123 VDD1.n103 VDD1.n102 9.3005
R2124 VDD1.n128 VDD1.n127 9.3005
R2125 VDD1.n126 VDD1.n125 9.3005
R2126 VDD1.n107 VDD1.n106 9.3005
R2127 VDD1.n120 VDD1.n119 9.3005
R2128 VDD1.n118 VDD1.n117 9.3005
R2129 VDD1.n111 VDD1.n110 9.3005
R2130 VDD1.n136 VDD1.n135 9.3005
R2131 VDD1.n99 VDD1.n98 9.3005
R2132 VDD1.n142 VDD1.n141 9.3005
R2133 VDD1.n144 VDD1.n143 9.3005
R2134 VDD1.n95 VDD1.n94 9.3005
R2135 VDD1.n150 VDD1.n149 9.3005
R2136 VDD1.n152 VDD1.n151 9.3005
R2137 VDD1.n153 VDD1.n90 9.3005
R2138 VDD1.n160 VDD1.n159 9.3005
R2139 VDD1.n61 VDD1.n14 8.92171
R2140 VDD1.n46 VDD1.n45 8.92171
R2141 VDD1.n129 VDD1.n128 8.92171
R2142 VDD1.n144 VDD1.n97 8.92171
R2143 VDD1.n58 VDD1.n57 8.14595
R2144 VDD1.n49 VDD1.n20 8.14595
R2145 VDD1.n132 VDD1.n103 8.14595
R2146 VDD1.n141 VDD1.n140 8.14595
R2147 VDD1.n54 VDD1.n16 7.3702
R2148 VDD1.n50 VDD1.n18 7.3702
R2149 VDD1.n133 VDD1.n101 7.3702
R2150 VDD1.n137 VDD1.n99 7.3702
R2151 VDD1.n54 VDD1.n53 6.59444
R2152 VDD1.n53 VDD1.n18 6.59444
R2153 VDD1.n136 VDD1.n101 6.59444
R2154 VDD1.n137 VDD1.n136 6.59444
R2155 VDD1.n57 VDD1.n16 5.81868
R2156 VDD1.n50 VDD1.n49 5.81868
R2157 VDD1.n133 VDD1.n132 5.81868
R2158 VDD1.n140 VDD1.n99 5.81868
R2159 VDD1.n58 VDD1.n14 5.04292
R2160 VDD1.n46 VDD1.n20 5.04292
R2161 VDD1.n129 VDD1.n103 5.04292
R2162 VDD1.n141 VDD1.n97 5.04292
R2163 VDD1.n62 VDD1.n61 4.26717
R2164 VDD1.n45 VDD1.n22 4.26717
R2165 VDD1.n128 VDD1.n105 4.26717
R2166 VDD1.n145 VDD1.n144 4.26717
R2167 VDD1.n29 VDD1.n27 3.70982
R2168 VDD1.n112 VDD1.n110 3.70982
R2169 VDD1.n65 VDD1.n12 3.49141
R2170 VDD1.n42 VDD1.n41 3.49141
R2171 VDD1.n125 VDD1.n124 3.49141
R2172 VDD1.n148 VDD1.n95 3.49141
R2173 VDD1.n84 VDD1.n0 2.71565
R2174 VDD1.n66 VDD1.n10 2.71565
R2175 VDD1.n38 VDD1.n24 2.71565
R2176 VDD1.n121 VDD1.n107 2.71565
R2177 VDD1.n149 VDD1.n93 2.71565
R2178 VDD1.n169 VDD1.n85 2.71565
R2179 VDD1.n172 VDD1.t1 2.10302
R2180 VDD1.n172 VDD1.t5 2.10302
R2181 VDD1.n170 VDD1.t4 2.10302
R2182 VDD1.n170 VDD1.t2 2.10302
R2183 VDD1.n82 VDD1.n81 1.93989
R2184 VDD1.n70 VDD1.n69 1.93989
R2185 VDD1.n37 VDD1.n26 1.93989
R2186 VDD1.n120 VDD1.n109 1.93989
R2187 VDD1.n154 VDD1.n152 1.93989
R2188 VDD1.n167 VDD1.n166 1.93989
R2189 VDD1.n78 VDD1.n2 1.16414
R2190 VDD1.n73 VDD1.n7 1.16414
R2191 VDD1.n34 VDD1.n33 1.16414
R2192 VDD1.n117 VDD1.n116 1.16414
R2193 VDD1.n153 VDD1.n91 1.16414
R2194 VDD1.n163 VDD1.n87 1.16414
R2195 VDD1 VDD1.n173 0.776362
R2196 VDD1.n77 VDD1.n4 0.388379
R2197 VDD1.n74 VDD1.n6 0.388379
R2198 VDD1.n30 VDD1.n28 0.388379
R2199 VDD1.n113 VDD1.n111 0.388379
R2200 VDD1.n159 VDD1.n158 0.388379
R2201 VDD1.n162 VDD1.n89 0.388379
R2202 VDD1.n83 VDD1.n1 0.155672
R2203 VDD1.n76 VDD1.n1 0.155672
R2204 VDD1.n76 VDD1.n75 0.155672
R2205 VDD1.n75 VDD1.n5 0.155672
R2206 VDD1.n68 VDD1.n5 0.155672
R2207 VDD1.n68 VDD1.n67 0.155672
R2208 VDD1.n67 VDD1.n11 0.155672
R2209 VDD1.n60 VDD1.n11 0.155672
R2210 VDD1.n60 VDD1.n59 0.155672
R2211 VDD1.n59 VDD1.n15 0.155672
R2212 VDD1.n52 VDD1.n15 0.155672
R2213 VDD1.n52 VDD1.n51 0.155672
R2214 VDD1.n51 VDD1.n19 0.155672
R2215 VDD1.n44 VDD1.n19 0.155672
R2216 VDD1.n44 VDD1.n43 0.155672
R2217 VDD1.n43 VDD1.n23 0.155672
R2218 VDD1.n36 VDD1.n23 0.155672
R2219 VDD1.n36 VDD1.n35 0.155672
R2220 VDD1.n35 VDD1.n27 0.155672
R2221 VDD1.n118 VDD1.n110 0.155672
R2222 VDD1.n119 VDD1.n118 0.155672
R2223 VDD1.n119 VDD1.n106 0.155672
R2224 VDD1.n126 VDD1.n106 0.155672
R2225 VDD1.n127 VDD1.n126 0.155672
R2226 VDD1.n127 VDD1.n102 0.155672
R2227 VDD1.n134 VDD1.n102 0.155672
R2228 VDD1.n135 VDD1.n134 0.155672
R2229 VDD1.n135 VDD1.n98 0.155672
R2230 VDD1.n142 VDD1.n98 0.155672
R2231 VDD1.n143 VDD1.n142 0.155672
R2232 VDD1.n143 VDD1.n94 0.155672
R2233 VDD1.n150 VDD1.n94 0.155672
R2234 VDD1.n151 VDD1.n150 0.155672
R2235 VDD1.n151 VDD1.n90 0.155672
R2236 VDD1.n160 VDD1.n90 0.155672
R2237 VDD1.n161 VDD1.n160 0.155672
R2238 VDD1.n161 VDD1.n86 0.155672
R2239 VDD1.n168 VDD1.n86 0.155672
R2240 VN.n38 VN.n37 161.3
R2241 VN.n36 VN.n21 161.3
R2242 VN.n35 VN.n34 161.3
R2243 VN.n33 VN.n22 161.3
R2244 VN.n32 VN.n31 161.3
R2245 VN.n30 VN.n23 161.3
R2246 VN.n29 VN.n28 161.3
R2247 VN.n27 VN.n24 161.3
R2248 VN.n18 VN.n17 161.3
R2249 VN.n16 VN.n1 161.3
R2250 VN.n15 VN.n14 161.3
R2251 VN.n13 VN.n2 161.3
R2252 VN.n12 VN.n11 161.3
R2253 VN.n10 VN.n3 161.3
R2254 VN.n9 VN.n8 161.3
R2255 VN.n7 VN.n4 161.3
R2256 VN.n26 VN.t2 137.962
R2257 VN.n6 VN.t5 137.962
R2258 VN.n5 VN.t0 105.251
R2259 VN.n0 VN.t4 105.251
R2260 VN.n25 VN.t3 105.251
R2261 VN.n20 VN.t1 105.251
R2262 VN.n19 VN.n0 84.3435
R2263 VN.n39 VN.n20 84.3435
R2264 VN.n6 VN.n5 62.4068
R2265 VN.n26 VN.n25 62.4068
R2266 VN.n11 VN.n2 56.5617
R2267 VN.n31 VN.n22 56.5617
R2268 VN VN.n39 55.1837
R2269 VN.n9 VN.n4 24.5923
R2270 VN.n10 VN.n9 24.5923
R2271 VN.n11 VN.n10 24.5923
R2272 VN.n15 VN.n2 24.5923
R2273 VN.n16 VN.n15 24.5923
R2274 VN.n17 VN.n16 24.5923
R2275 VN.n31 VN.n30 24.5923
R2276 VN.n30 VN.n29 24.5923
R2277 VN.n29 VN.n24 24.5923
R2278 VN.n37 VN.n36 24.5923
R2279 VN.n36 VN.n35 24.5923
R2280 VN.n35 VN.n22 24.5923
R2281 VN.n5 VN.n4 12.2964
R2282 VN.n25 VN.n24 12.2964
R2283 VN.n17 VN.n0 5.90254
R2284 VN.n37 VN.n20 5.90254
R2285 VN.n27 VN.n26 3.27862
R2286 VN.n7 VN.n6 3.27862
R2287 VN.n39 VN.n38 0.354861
R2288 VN.n19 VN.n18 0.354861
R2289 VN VN.n19 0.267071
R2290 VN.n38 VN.n21 0.189894
R2291 VN.n34 VN.n21 0.189894
R2292 VN.n34 VN.n33 0.189894
R2293 VN.n33 VN.n32 0.189894
R2294 VN.n32 VN.n23 0.189894
R2295 VN.n28 VN.n23 0.189894
R2296 VN.n28 VN.n27 0.189894
R2297 VN.n8 VN.n7 0.189894
R2298 VN.n8 VN.n3 0.189894
R2299 VN.n12 VN.n3 0.189894
R2300 VN.n13 VN.n12 0.189894
R2301 VN.n14 VN.n13 0.189894
R2302 VN.n14 VN.n1 0.189894
R2303 VN.n18 VN.n1 0.189894
R2304 VDD2.n167 VDD2.n87 756.745
R2305 VDD2.n80 VDD2.n0 756.745
R2306 VDD2.n168 VDD2.n167 585
R2307 VDD2.n166 VDD2.n165 585
R2308 VDD2.n91 VDD2.n90 585
R2309 VDD2.n95 VDD2.n93 585
R2310 VDD2.n160 VDD2.n159 585
R2311 VDD2.n158 VDD2.n157 585
R2312 VDD2.n97 VDD2.n96 585
R2313 VDD2.n152 VDD2.n151 585
R2314 VDD2.n150 VDD2.n149 585
R2315 VDD2.n101 VDD2.n100 585
R2316 VDD2.n144 VDD2.n143 585
R2317 VDD2.n142 VDD2.n141 585
R2318 VDD2.n105 VDD2.n104 585
R2319 VDD2.n136 VDD2.n135 585
R2320 VDD2.n134 VDD2.n133 585
R2321 VDD2.n109 VDD2.n108 585
R2322 VDD2.n128 VDD2.n127 585
R2323 VDD2.n126 VDD2.n125 585
R2324 VDD2.n113 VDD2.n112 585
R2325 VDD2.n120 VDD2.n119 585
R2326 VDD2.n118 VDD2.n117 585
R2327 VDD2.n29 VDD2.n28 585
R2328 VDD2.n31 VDD2.n30 585
R2329 VDD2.n24 VDD2.n23 585
R2330 VDD2.n37 VDD2.n36 585
R2331 VDD2.n39 VDD2.n38 585
R2332 VDD2.n20 VDD2.n19 585
R2333 VDD2.n45 VDD2.n44 585
R2334 VDD2.n47 VDD2.n46 585
R2335 VDD2.n16 VDD2.n15 585
R2336 VDD2.n53 VDD2.n52 585
R2337 VDD2.n55 VDD2.n54 585
R2338 VDD2.n12 VDD2.n11 585
R2339 VDD2.n61 VDD2.n60 585
R2340 VDD2.n63 VDD2.n62 585
R2341 VDD2.n8 VDD2.n7 585
R2342 VDD2.n70 VDD2.n69 585
R2343 VDD2.n71 VDD2.n6 585
R2344 VDD2.n73 VDD2.n72 585
R2345 VDD2.n4 VDD2.n3 585
R2346 VDD2.n79 VDD2.n78 585
R2347 VDD2.n81 VDD2.n80 585
R2348 VDD2.n116 VDD2.t4 327.466
R2349 VDD2.n27 VDD2.t0 327.466
R2350 VDD2.n167 VDD2.n166 171.744
R2351 VDD2.n166 VDD2.n90 171.744
R2352 VDD2.n95 VDD2.n90 171.744
R2353 VDD2.n159 VDD2.n95 171.744
R2354 VDD2.n159 VDD2.n158 171.744
R2355 VDD2.n158 VDD2.n96 171.744
R2356 VDD2.n151 VDD2.n96 171.744
R2357 VDD2.n151 VDD2.n150 171.744
R2358 VDD2.n150 VDD2.n100 171.744
R2359 VDD2.n143 VDD2.n100 171.744
R2360 VDD2.n143 VDD2.n142 171.744
R2361 VDD2.n142 VDD2.n104 171.744
R2362 VDD2.n135 VDD2.n104 171.744
R2363 VDD2.n135 VDD2.n134 171.744
R2364 VDD2.n134 VDD2.n108 171.744
R2365 VDD2.n127 VDD2.n108 171.744
R2366 VDD2.n127 VDD2.n126 171.744
R2367 VDD2.n126 VDD2.n112 171.744
R2368 VDD2.n119 VDD2.n112 171.744
R2369 VDD2.n119 VDD2.n118 171.744
R2370 VDD2.n30 VDD2.n29 171.744
R2371 VDD2.n30 VDD2.n23 171.744
R2372 VDD2.n37 VDD2.n23 171.744
R2373 VDD2.n38 VDD2.n37 171.744
R2374 VDD2.n38 VDD2.n19 171.744
R2375 VDD2.n45 VDD2.n19 171.744
R2376 VDD2.n46 VDD2.n45 171.744
R2377 VDD2.n46 VDD2.n15 171.744
R2378 VDD2.n53 VDD2.n15 171.744
R2379 VDD2.n54 VDD2.n53 171.744
R2380 VDD2.n54 VDD2.n11 171.744
R2381 VDD2.n61 VDD2.n11 171.744
R2382 VDD2.n62 VDD2.n61 171.744
R2383 VDD2.n62 VDD2.n7 171.744
R2384 VDD2.n70 VDD2.n7 171.744
R2385 VDD2.n71 VDD2.n70 171.744
R2386 VDD2.n72 VDD2.n71 171.744
R2387 VDD2.n72 VDD2.n3 171.744
R2388 VDD2.n79 VDD2.n3 171.744
R2389 VDD2.n80 VDD2.n79 171.744
R2390 VDD2.n118 VDD2.t4 85.8723
R2391 VDD2.n29 VDD2.t0 85.8723
R2392 VDD2.n86 VDD2.n85 72.9761
R2393 VDD2 VDD2.n173 72.9732
R2394 VDD2.n86 VDD2.n84 53.2503
R2395 VDD2.n172 VDD2.n171 50.8035
R2396 VDD2.n172 VDD2.n86 47.8856
R2397 VDD2.n117 VDD2.n116 16.3895
R2398 VDD2.n28 VDD2.n27 16.3895
R2399 VDD2.n93 VDD2.n91 13.1884
R2400 VDD2.n73 VDD2.n4 13.1884
R2401 VDD2.n165 VDD2.n164 12.8005
R2402 VDD2.n161 VDD2.n160 12.8005
R2403 VDD2.n120 VDD2.n115 12.8005
R2404 VDD2.n31 VDD2.n26 12.8005
R2405 VDD2.n74 VDD2.n6 12.8005
R2406 VDD2.n78 VDD2.n77 12.8005
R2407 VDD2.n168 VDD2.n89 12.0247
R2408 VDD2.n157 VDD2.n94 12.0247
R2409 VDD2.n121 VDD2.n113 12.0247
R2410 VDD2.n32 VDD2.n24 12.0247
R2411 VDD2.n69 VDD2.n68 12.0247
R2412 VDD2.n81 VDD2.n2 12.0247
R2413 VDD2.n169 VDD2.n87 11.249
R2414 VDD2.n156 VDD2.n97 11.249
R2415 VDD2.n125 VDD2.n124 11.249
R2416 VDD2.n36 VDD2.n35 11.249
R2417 VDD2.n67 VDD2.n8 11.249
R2418 VDD2.n82 VDD2.n0 11.249
R2419 VDD2.n153 VDD2.n152 10.4732
R2420 VDD2.n128 VDD2.n111 10.4732
R2421 VDD2.n39 VDD2.n22 10.4732
R2422 VDD2.n64 VDD2.n63 10.4732
R2423 VDD2.n149 VDD2.n99 9.69747
R2424 VDD2.n129 VDD2.n109 9.69747
R2425 VDD2.n40 VDD2.n20 9.69747
R2426 VDD2.n60 VDD2.n10 9.69747
R2427 VDD2.n171 VDD2.n170 9.45567
R2428 VDD2.n84 VDD2.n83 9.45567
R2429 VDD2.n103 VDD2.n102 9.3005
R2430 VDD2.n146 VDD2.n145 9.3005
R2431 VDD2.n148 VDD2.n147 9.3005
R2432 VDD2.n99 VDD2.n98 9.3005
R2433 VDD2.n154 VDD2.n153 9.3005
R2434 VDD2.n156 VDD2.n155 9.3005
R2435 VDD2.n94 VDD2.n92 9.3005
R2436 VDD2.n162 VDD2.n161 9.3005
R2437 VDD2.n170 VDD2.n169 9.3005
R2438 VDD2.n89 VDD2.n88 9.3005
R2439 VDD2.n164 VDD2.n163 9.3005
R2440 VDD2.n140 VDD2.n139 9.3005
R2441 VDD2.n138 VDD2.n137 9.3005
R2442 VDD2.n107 VDD2.n106 9.3005
R2443 VDD2.n132 VDD2.n131 9.3005
R2444 VDD2.n130 VDD2.n129 9.3005
R2445 VDD2.n111 VDD2.n110 9.3005
R2446 VDD2.n124 VDD2.n123 9.3005
R2447 VDD2.n122 VDD2.n121 9.3005
R2448 VDD2.n115 VDD2.n114 9.3005
R2449 VDD2.n83 VDD2.n82 9.3005
R2450 VDD2.n2 VDD2.n1 9.3005
R2451 VDD2.n77 VDD2.n76 9.3005
R2452 VDD2.n49 VDD2.n48 9.3005
R2453 VDD2.n18 VDD2.n17 9.3005
R2454 VDD2.n43 VDD2.n42 9.3005
R2455 VDD2.n41 VDD2.n40 9.3005
R2456 VDD2.n22 VDD2.n21 9.3005
R2457 VDD2.n35 VDD2.n34 9.3005
R2458 VDD2.n33 VDD2.n32 9.3005
R2459 VDD2.n26 VDD2.n25 9.3005
R2460 VDD2.n51 VDD2.n50 9.3005
R2461 VDD2.n14 VDD2.n13 9.3005
R2462 VDD2.n57 VDD2.n56 9.3005
R2463 VDD2.n59 VDD2.n58 9.3005
R2464 VDD2.n10 VDD2.n9 9.3005
R2465 VDD2.n65 VDD2.n64 9.3005
R2466 VDD2.n67 VDD2.n66 9.3005
R2467 VDD2.n68 VDD2.n5 9.3005
R2468 VDD2.n75 VDD2.n74 9.3005
R2469 VDD2.n148 VDD2.n101 8.92171
R2470 VDD2.n133 VDD2.n132 8.92171
R2471 VDD2.n44 VDD2.n43 8.92171
R2472 VDD2.n59 VDD2.n12 8.92171
R2473 VDD2.n145 VDD2.n144 8.14595
R2474 VDD2.n136 VDD2.n107 8.14595
R2475 VDD2.n47 VDD2.n18 8.14595
R2476 VDD2.n56 VDD2.n55 8.14595
R2477 VDD2.n141 VDD2.n103 7.3702
R2478 VDD2.n137 VDD2.n105 7.3702
R2479 VDD2.n48 VDD2.n16 7.3702
R2480 VDD2.n52 VDD2.n14 7.3702
R2481 VDD2.n141 VDD2.n140 6.59444
R2482 VDD2.n140 VDD2.n105 6.59444
R2483 VDD2.n51 VDD2.n16 6.59444
R2484 VDD2.n52 VDD2.n51 6.59444
R2485 VDD2.n144 VDD2.n103 5.81868
R2486 VDD2.n137 VDD2.n136 5.81868
R2487 VDD2.n48 VDD2.n47 5.81868
R2488 VDD2.n55 VDD2.n14 5.81868
R2489 VDD2.n145 VDD2.n101 5.04292
R2490 VDD2.n133 VDD2.n107 5.04292
R2491 VDD2.n44 VDD2.n18 5.04292
R2492 VDD2.n56 VDD2.n12 5.04292
R2493 VDD2.n149 VDD2.n148 4.26717
R2494 VDD2.n132 VDD2.n109 4.26717
R2495 VDD2.n43 VDD2.n20 4.26717
R2496 VDD2.n60 VDD2.n59 4.26717
R2497 VDD2.n116 VDD2.n114 3.70982
R2498 VDD2.n27 VDD2.n25 3.70982
R2499 VDD2.n152 VDD2.n99 3.49141
R2500 VDD2.n129 VDD2.n128 3.49141
R2501 VDD2.n40 VDD2.n39 3.49141
R2502 VDD2.n63 VDD2.n10 3.49141
R2503 VDD2.n171 VDD2.n87 2.71565
R2504 VDD2.n153 VDD2.n97 2.71565
R2505 VDD2.n125 VDD2.n111 2.71565
R2506 VDD2.n36 VDD2.n22 2.71565
R2507 VDD2.n64 VDD2.n8 2.71565
R2508 VDD2.n84 VDD2.n0 2.71565
R2509 VDD2 VDD2.n172 2.56084
R2510 VDD2.n173 VDD2.t2 2.10302
R2511 VDD2.n173 VDD2.t3 2.10302
R2512 VDD2.n85 VDD2.t5 2.10302
R2513 VDD2.n85 VDD2.t1 2.10302
R2514 VDD2.n169 VDD2.n168 1.93989
R2515 VDD2.n157 VDD2.n156 1.93989
R2516 VDD2.n124 VDD2.n113 1.93989
R2517 VDD2.n35 VDD2.n24 1.93989
R2518 VDD2.n69 VDD2.n67 1.93989
R2519 VDD2.n82 VDD2.n81 1.93989
R2520 VDD2.n165 VDD2.n89 1.16414
R2521 VDD2.n160 VDD2.n94 1.16414
R2522 VDD2.n121 VDD2.n120 1.16414
R2523 VDD2.n32 VDD2.n31 1.16414
R2524 VDD2.n68 VDD2.n6 1.16414
R2525 VDD2.n78 VDD2.n2 1.16414
R2526 VDD2.n164 VDD2.n91 0.388379
R2527 VDD2.n161 VDD2.n93 0.388379
R2528 VDD2.n117 VDD2.n115 0.388379
R2529 VDD2.n28 VDD2.n26 0.388379
R2530 VDD2.n74 VDD2.n73 0.388379
R2531 VDD2.n77 VDD2.n4 0.388379
R2532 VDD2.n170 VDD2.n88 0.155672
R2533 VDD2.n163 VDD2.n88 0.155672
R2534 VDD2.n163 VDD2.n162 0.155672
R2535 VDD2.n162 VDD2.n92 0.155672
R2536 VDD2.n155 VDD2.n92 0.155672
R2537 VDD2.n155 VDD2.n154 0.155672
R2538 VDD2.n154 VDD2.n98 0.155672
R2539 VDD2.n147 VDD2.n98 0.155672
R2540 VDD2.n147 VDD2.n146 0.155672
R2541 VDD2.n146 VDD2.n102 0.155672
R2542 VDD2.n139 VDD2.n102 0.155672
R2543 VDD2.n139 VDD2.n138 0.155672
R2544 VDD2.n138 VDD2.n106 0.155672
R2545 VDD2.n131 VDD2.n106 0.155672
R2546 VDD2.n131 VDD2.n130 0.155672
R2547 VDD2.n130 VDD2.n110 0.155672
R2548 VDD2.n123 VDD2.n110 0.155672
R2549 VDD2.n123 VDD2.n122 0.155672
R2550 VDD2.n122 VDD2.n114 0.155672
R2551 VDD2.n33 VDD2.n25 0.155672
R2552 VDD2.n34 VDD2.n33 0.155672
R2553 VDD2.n34 VDD2.n21 0.155672
R2554 VDD2.n41 VDD2.n21 0.155672
R2555 VDD2.n42 VDD2.n41 0.155672
R2556 VDD2.n42 VDD2.n17 0.155672
R2557 VDD2.n49 VDD2.n17 0.155672
R2558 VDD2.n50 VDD2.n49 0.155672
R2559 VDD2.n50 VDD2.n13 0.155672
R2560 VDD2.n57 VDD2.n13 0.155672
R2561 VDD2.n58 VDD2.n57 0.155672
R2562 VDD2.n58 VDD2.n9 0.155672
R2563 VDD2.n65 VDD2.n9 0.155672
R2564 VDD2.n66 VDD2.n65 0.155672
R2565 VDD2.n66 VDD2.n5 0.155672
R2566 VDD2.n75 VDD2.n5 0.155672
R2567 VDD2.n76 VDD2.n75 0.155672
R2568 VDD2.n76 VDD2.n1 0.155672
R2569 VDD2.n83 VDD2.n1 0.155672
C0 VP VTAIL 9.23715f
C1 VTAIL w_n4066_n4060# 3.52972f
C2 VDD1 VDD2 1.77469f
C3 B VN 1.41075f
C4 VP VDD1 9.3833f
C5 VDD1 w_n4066_n4060# 2.75764f
C6 B VTAIL 4.86502f
C7 VP VDD2 0.538677f
C8 VDD2 w_n4066_n4060# 2.87276f
C9 VN VTAIL 9.22289f
C10 B VDD1 2.61623f
C11 VP w_n4066_n4060# 8.51722f
C12 B VDD2 2.71287f
C13 VN VDD1 0.152453f
C14 VN VDD2 9.00059f
C15 B VP 2.29753f
C16 B w_n4066_n4060# 11.944401f
C17 VTAIL VDD1 9.16501f
C18 VP VN 8.47802f
C19 VN w_n4066_n4060# 7.98892f
C20 VTAIL VDD2 9.22237f
C21 VDD2 VSUBS 2.23345f
C22 VDD1 VSUBS 2.245789f
C23 VTAIL VSUBS 1.49153f
C24 VN VSUBS 6.86953f
C25 VP VSUBS 3.790312f
C26 B VSUBS 5.858046f
C27 w_n4066_n4060# VSUBS 0.20234p
C28 VDD2.n0 VSUBS 0.029595f
C29 VDD2.n1 VSUBS 0.027681f
C30 VDD2.n2 VSUBS 0.014874f
C31 VDD2.n3 VSUBS 0.035157f
C32 VDD2.n4 VSUBS 0.015312f
C33 VDD2.n5 VSUBS 0.027681f
C34 VDD2.n6 VSUBS 0.015749f
C35 VDD2.n7 VSUBS 0.035157f
C36 VDD2.n8 VSUBS 0.015749f
C37 VDD2.n9 VSUBS 0.027681f
C38 VDD2.n10 VSUBS 0.014874f
C39 VDD2.n11 VSUBS 0.035157f
C40 VDD2.n12 VSUBS 0.015749f
C41 VDD2.n13 VSUBS 0.027681f
C42 VDD2.n14 VSUBS 0.014874f
C43 VDD2.n15 VSUBS 0.035157f
C44 VDD2.n16 VSUBS 0.015749f
C45 VDD2.n17 VSUBS 0.027681f
C46 VDD2.n18 VSUBS 0.014874f
C47 VDD2.n19 VSUBS 0.035157f
C48 VDD2.n20 VSUBS 0.015749f
C49 VDD2.n21 VSUBS 0.027681f
C50 VDD2.n22 VSUBS 0.014874f
C51 VDD2.n23 VSUBS 0.035157f
C52 VDD2.n24 VSUBS 0.015749f
C53 VDD2.n25 VSUBS 1.82526f
C54 VDD2.n26 VSUBS 0.014874f
C55 VDD2.t0 VSUBS 0.075297f
C56 VDD2.n27 VSUBS 0.198879f
C57 VDD2.n28 VSUBS 0.022365f
C58 VDD2.n29 VSUBS 0.026368f
C59 VDD2.n30 VSUBS 0.035157f
C60 VDD2.n31 VSUBS 0.015749f
C61 VDD2.n32 VSUBS 0.014874f
C62 VDD2.n33 VSUBS 0.027681f
C63 VDD2.n34 VSUBS 0.027681f
C64 VDD2.n35 VSUBS 0.014874f
C65 VDD2.n36 VSUBS 0.015749f
C66 VDD2.n37 VSUBS 0.035157f
C67 VDD2.n38 VSUBS 0.035157f
C68 VDD2.n39 VSUBS 0.015749f
C69 VDD2.n40 VSUBS 0.014874f
C70 VDD2.n41 VSUBS 0.027681f
C71 VDD2.n42 VSUBS 0.027681f
C72 VDD2.n43 VSUBS 0.014874f
C73 VDD2.n44 VSUBS 0.015749f
C74 VDD2.n45 VSUBS 0.035157f
C75 VDD2.n46 VSUBS 0.035157f
C76 VDD2.n47 VSUBS 0.015749f
C77 VDD2.n48 VSUBS 0.014874f
C78 VDD2.n49 VSUBS 0.027681f
C79 VDD2.n50 VSUBS 0.027681f
C80 VDD2.n51 VSUBS 0.014874f
C81 VDD2.n52 VSUBS 0.015749f
C82 VDD2.n53 VSUBS 0.035157f
C83 VDD2.n54 VSUBS 0.035157f
C84 VDD2.n55 VSUBS 0.015749f
C85 VDD2.n56 VSUBS 0.014874f
C86 VDD2.n57 VSUBS 0.027681f
C87 VDD2.n58 VSUBS 0.027681f
C88 VDD2.n59 VSUBS 0.014874f
C89 VDD2.n60 VSUBS 0.015749f
C90 VDD2.n61 VSUBS 0.035157f
C91 VDD2.n62 VSUBS 0.035157f
C92 VDD2.n63 VSUBS 0.015749f
C93 VDD2.n64 VSUBS 0.014874f
C94 VDD2.n65 VSUBS 0.027681f
C95 VDD2.n66 VSUBS 0.027681f
C96 VDD2.n67 VSUBS 0.014874f
C97 VDD2.n68 VSUBS 0.014874f
C98 VDD2.n69 VSUBS 0.015749f
C99 VDD2.n70 VSUBS 0.035157f
C100 VDD2.n71 VSUBS 0.035157f
C101 VDD2.n72 VSUBS 0.035157f
C102 VDD2.n73 VSUBS 0.015312f
C103 VDD2.n74 VSUBS 0.014874f
C104 VDD2.n75 VSUBS 0.027681f
C105 VDD2.n76 VSUBS 0.027681f
C106 VDD2.n77 VSUBS 0.014874f
C107 VDD2.n78 VSUBS 0.015749f
C108 VDD2.n79 VSUBS 0.035157f
C109 VDD2.n80 VSUBS 0.08232f
C110 VDD2.n81 VSUBS 0.015749f
C111 VDD2.n82 VSUBS 0.014874f
C112 VDD2.n83 VSUBS 0.067763f
C113 VDD2.n84 VSUBS 0.073061f
C114 VDD2.t5 VSUBS 0.338171f
C115 VDD2.t1 VSUBS 0.338171f
C116 VDD2.n85 VSUBS 2.77285f
C117 VDD2.n86 VSUBS 3.95059f
C118 VDD2.n87 VSUBS 0.029595f
C119 VDD2.n88 VSUBS 0.027681f
C120 VDD2.n89 VSUBS 0.014874f
C121 VDD2.n90 VSUBS 0.035157f
C122 VDD2.n91 VSUBS 0.015312f
C123 VDD2.n92 VSUBS 0.027681f
C124 VDD2.n93 VSUBS 0.015312f
C125 VDD2.n94 VSUBS 0.014874f
C126 VDD2.n95 VSUBS 0.035157f
C127 VDD2.n96 VSUBS 0.035157f
C128 VDD2.n97 VSUBS 0.015749f
C129 VDD2.n98 VSUBS 0.027681f
C130 VDD2.n99 VSUBS 0.014874f
C131 VDD2.n100 VSUBS 0.035157f
C132 VDD2.n101 VSUBS 0.015749f
C133 VDD2.n102 VSUBS 0.027681f
C134 VDD2.n103 VSUBS 0.014874f
C135 VDD2.n104 VSUBS 0.035157f
C136 VDD2.n105 VSUBS 0.015749f
C137 VDD2.n106 VSUBS 0.027681f
C138 VDD2.n107 VSUBS 0.014874f
C139 VDD2.n108 VSUBS 0.035157f
C140 VDD2.n109 VSUBS 0.015749f
C141 VDD2.n110 VSUBS 0.027681f
C142 VDD2.n111 VSUBS 0.014874f
C143 VDD2.n112 VSUBS 0.035157f
C144 VDD2.n113 VSUBS 0.015749f
C145 VDD2.n114 VSUBS 1.82526f
C146 VDD2.n115 VSUBS 0.014874f
C147 VDD2.t4 VSUBS 0.075297f
C148 VDD2.n116 VSUBS 0.198879f
C149 VDD2.n117 VSUBS 0.022365f
C150 VDD2.n118 VSUBS 0.026368f
C151 VDD2.n119 VSUBS 0.035157f
C152 VDD2.n120 VSUBS 0.015749f
C153 VDD2.n121 VSUBS 0.014874f
C154 VDD2.n122 VSUBS 0.027681f
C155 VDD2.n123 VSUBS 0.027681f
C156 VDD2.n124 VSUBS 0.014874f
C157 VDD2.n125 VSUBS 0.015749f
C158 VDD2.n126 VSUBS 0.035157f
C159 VDD2.n127 VSUBS 0.035157f
C160 VDD2.n128 VSUBS 0.015749f
C161 VDD2.n129 VSUBS 0.014874f
C162 VDD2.n130 VSUBS 0.027681f
C163 VDD2.n131 VSUBS 0.027681f
C164 VDD2.n132 VSUBS 0.014874f
C165 VDD2.n133 VSUBS 0.015749f
C166 VDD2.n134 VSUBS 0.035157f
C167 VDD2.n135 VSUBS 0.035157f
C168 VDD2.n136 VSUBS 0.015749f
C169 VDD2.n137 VSUBS 0.014874f
C170 VDD2.n138 VSUBS 0.027681f
C171 VDD2.n139 VSUBS 0.027681f
C172 VDD2.n140 VSUBS 0.014874f
C173 VDD2.n141 VSUBS 0.015749f
C174 VDD2.n142 VSUBS 0.035157f
C175 VDD2.n143 VSUBS 0.035157f
C176 VDD2.n144 VSUBS 0.015749f
C177 VDD2.n145 VSUBS 0.014874f
C178 VDD2.n146 VSUBS 0.027681f
C179 VDD2.n147 VSUBS 0.027681f
C180 VDD2.n148 VSUBS 0.014874f
C181 VDD2.n149 VSUBS 0.015749f
C182 VDD2.n150 VSUBS 0.035157f
C183 VDD2.n151 VSUBS 0.035157f
C184 VDD2.n152 VSUBS 0.015749f
C185 VDD2.n153 VSUBS 0.014874f
C186 VDD2.n154 VSUBS 0.027681f
C187 VDD2.n155 VSUBS 0.027681f
C188 VDD2.n156 VSUBS 0.014874f
C189 VDD2.n157 VSUBS 0.015749f
C190 VDD2.n158 VSUBS 0.035157f
C191 VDD2.n159 VSUBS 0.035157f
C192 VDD2.n160 VSUBS 0.015749f
C193 VDD2.n161 VSUBS 0.014874f
C194 VDD2.n162 VSUBS 0.027681f
C195 VDD2.n163 VSUBS 0.027681f
C196 VDD2.n164 VSUBS 0.014874f
C197 VDD2.n165 VSUBS 0.015749f
C198 VDD2.n166 VSUBS 0.035157f
C199 VDD2.n167 VSUBS 0.08232f
C200 VDD2.n168 VSUBS 0.015749f
C201 VDD2.n169 VSUBS 0.014874f
C202 VDD2.n170 VSUBS 0.067763f
C203 VDD2.n171 VSUBS 0.060472f
C204 VDD2.n172 VSUBS 3.41531f
C205 VDD2.t2 VSUBS 0.338171f
C206 VDD2.t3 VSUBS 0.338171f
C207 VDD2.n173 VSUBS 2.77281f
C208 VN.t4 VSUBS 3.57714f
C209 VN.n0 VSUBS 1.32725f
C210 VN.n1 VSUBS 0.023837f
C211 VN.n2 VSUBS 0.038937f
C212 VN.n3 VSUBS 0.023837f
C213 VN.n4 VSUBS 0.033292f
C214 VN.t0 VSUBS 3.57714f
C215 VN.n5 VSUBS 1.32206f
C216 VN.t5 VSUBS 3.91318f
C217 VN.n6 VSUBS 1.26269f
C218 VN.n7 VSUBS 0.296936f
C219 VN.n8 VSUBS 0.023837f
C220 VN.n9 VSUBS 0.044203f
C221 VN.n10 VSUBS 0.044203f
C222 VN.n11 VSUBS 0.030364f
C223 VN.n12 VSUBS 0.023837f
C224 VN.n13 VSUBS 0.023837f
C225 VN.n14 VSUBS 0.023837f
C226 VN.n15 VSUBS 0.044203f
C227 VN.n16 VSUBS 0.044203f
C228 VN.n17 VSUBS 0.027618f
C229 VN.n18 VSUBS 0.038466f
C230 VN.n19 VSUBS 0.067652f
C231 VN.t1 VSUBS 3.57714f
C232 VN.n20 VSUBS 1.32725f
C233 VN.n21 VSUBS 0.023837f
C234 VN.n22 VSUBS 0.038937f
C235 VN.n23 VSUBS 0.023837f
C236 VN.n24 VSUBS 0.033292f
C237 VN.t2 VSUBS 3.91318f
C238 VN.t3 VSUBS 3.57714f
C239 VN.n25 VSUBS 1.32206f
C240 VN.n26 VSUBS 1.26269f
C241 VN.n27 VSUBS 0.296936f
C242 VN.n28 VSUBS 0.023837f
C243 VN.n29 VSUBS 0.044203f
C244 VN.n30 VSUBS 0.044203f
C245 VN.n31 VSUBS 0.030364f
C246 VN.n32 VSUBS 0.023837f
C247 VN.n33 VSUBS 0.023837f
C248 VN.n34 VSUBS 0.023837f
C249 VN.n35 VSUBS 0.044203f
C250 VN.n36 VSUBS 0.044203f
C251 VN.n37 VSUBS 0.027618f
C252 VN.n38 VSUBS 0.038466f
C253 VN.n39 VSUBS 1.57f
C254 VDD1.n0 VSUBS 0.029716f
C255 VDD1.n1 VSUBS 0.027794f
C256 VDD1.n2 VSUBS 0.014935f
C257 VDD1.n3 VSUBS 0.035301f
C258 VDD1.n4 VSUBS 0.015374f
C259 VDD1.n5 VSUBS 0.027794f
C260 VDD1.n6 VSUBS 0.015374f
C261 VDD1.n7 VSUBS 0.014935f
C262 VDD1.n8 VSUBS 0.035301f
C263 VDD1.n9 VSUBS 0.035301f
C264 VDD1.n10 VSUBS 0.015814f
C265 VDD1.n11 VSUBS 0.027794f
C266 VDD1.n12 VSUBS 0.014935f
C267 VDD1.n13 VSUBS 0.035301f
C268 VDD1.n14 VSUBS 0.015814f
C269 VDD1.n15 VSUBS 0.027794f
C270 VDD1.n16 VSUBS 0.014935f
C271 VDD1.n17 VSUBS 0.035301f
C272 VDD1.n18 VSUBS 0.015814f
C273 VDD1.n19 VSUBS 0.027794f
C274 VDD1.n20 VSUBS 0.014935f
C275 VDD1.n21 VSUBS 0.035301f
C276 VDD1.n22 VSUBS 0.015814f
C277 VDD1.n23 VSUBS 0.027794f
C278 VDD1.n24 VSUBS 0.014935f
C279 VDD1.n25 VSUBS 0.035301f
C280 VDD1.n26 VSUBS 0.015814f
C281 VDD1.n27 VSUBS 1.83272f
C282 VDD1.n28 VSUBS 0.014935f
C283 VDD1.t0 VSUBS 0.075605f
C284 VDD1.n29 VSUBS 0.199692f
C285 VDD1.n30 VSUBS 0.022457f
C286 VDD1.n31 VSUBS 0.026476f
C287 VDD1.n32 VSUBS 0.035301f
C288 VDD1.n33 VSUBS 0.015814f
C289 VDD1.n34 VSUBS 0.014935f
C290 VDD1.n35 VSUBS 0.027794f
C291 VDD1.n36 VSUBS 0.027794f
C292 VDD1.n37 VSUBS 0.014935f
C293 VDD1.n38 VSUBS 0.015814f
C294 VDD1.n39 VSUBS 0.035301f
C295 VDD1.n40 VSUBS 0.035301f
C296 VDD1.n41 VSUBS 0.015814f
C297 VDD1.n42 VSUBS 0.014935f
C298 VDD1.n43 VSUBS 0.027794f
C299 VDD1.n44 VSUBS 0.027794f
C300 VDD1.n45 VSUBS 0.014935f
C301 VDD1.n46 VSUBS 0.015814f
C302 VDD1.n47 VSUBS 0.035301f
C303 VDD1.n48 VSUBS 0.035301f
C304 VDD1.n49 VSUBS 0.015814f
C305 VDD1.n50 VSUBS 0.014935f
C306 VDD1.n51 VSUBS 0.027794f
C307 VDD1.n52 VSUBS 0.027794f
C308 VDD1.n53 VSUBS 0.014935f
C309 VDD1.n54 VSUBS 0.015814f
C310 VDD1.n55 VSUBS 0.035301f
C311 VDD1.n56 VSUBS 0.035301f
C312 VDD1.n57 VSUBS 0.015814f
C313 VDD1.n58 VSUBS 0.014935f
C314 VDD1.n59 VSUBS 0.027794f
C315 VDD1.n60 VSUBS 0.027794f
C316 VDD1.n61 VSUBS 0.014935f
C317 VDD1.n62 VSUBS 0.015814f
C318 VDD1.n63 VSUBS 0.035301f
C319 VDD1.n64 VSUBS 0.035301f
C320 VDD1.n65 VSUBS 0.015814f
C321 VDD1.n66 VSUBS 0.014935f
C322 VDD1.n67 VSUBS 0.027794f
C323 VDD1.n68 VSUBS 0.027794f
C324 VDD1.n69 VSUBS 0.014935f
C325 VDD1.n70 VSUBS 0.015814f
C326 VDD1.n71 VSUBS 0.035301f
C327 VDD1.n72 VSUBS 0.035301f
C328 VDD1.n73 VSUBS 0.015814f
C329 VDD1.n74 VSUBS 0.014935f
C330 VDD1.n75 VSUBS 0.027794f
C331 VDD1.n76 VSUBS 0.027794f
C332 VDD1.n77 VSUBS 0.014935f
C333 VDD1.n78 VSUBS 0.015814f
C334 VDD1.n79 VSUBS 0.035301f
C335 VDD1.n80 VSUBS 0.082657f
C336 VDD1.n81 VSUBS 0.015814f
C337 VDD1.n82 VSUBS 0.014935f
C338 VDD1.n83 VSUBS 0.068041f
C339 VDD1.n84 VSUBS 0.074393f
C340 VDD1.n85 VSUBS 0.029716f
C341 VDD1.n86 VSUBS 0.027794f
C342 VDD1.n87 VSUBS 0.014935f
C343 VDD1.n88 VSUBS 0.035301f
C344 VDD1.n89 VSUBS 0.015374f
C345 VDD1.n90 VSUBS 0.027794f
C346 VDD1.n91 VSUBS 0.015814f
C347 VDD1.n92 VSUBS 0.035301f
C348 VDD1.n93 VSUBS 0.015814f
C349 VDD1.n94 VSUBS 0.027794f
C350 VDD1.n95 VSUBS 0.014935f
C351 VDD1.n96 VSUBS 0.035301f
C352 VDD1.n97 VSUBS 0.015814f
C353 VDD1.n98 VSUBS 0.027794f
C354 VDD1.n99 VSUBS 0.014935f
C355 VDD1.n100 VSUBS 0.035301f
C356 VDD1.n101 VSUBS 0.015814f
C357 VDD1.n102 VSUBS 0.027794f
C358 VDD1.n103 VSUBS 0.014935f
C359 VDD1.n104 VSUBS 0.035301f
C360 VDD1.n105 VSUBS 0.015814f
C361 VDD1.n106 VSUBS 0.027794f
C362 VDD1.n107 VSUBS 0.014935f
C363 VDD1.n108 VSUBS 0.035301f
C364 VDD1.n109 VSUBS 0.015814f
C365 VDD1.n110 VSUBS 1.83272f
C366 VDD1.n111 VSUBS 0.014935f
C367 VDD1.t3 VSUBS 0.075605f
C368 VDD1.n112 VSUBS 0.199692f
C369 VDD1.n113 VSUBS 0.022457f
C370 VDD1.n114 VSUBS 0.026476f
C371 VDD1.n115 VSUBS 0.035301f
C372 VDD1.n116 VSUBS 0.015814f
C373 VDD1.n117 VSUBS 0.014935f
C374 VDD1.n118 VSUBS 0.027794f
C375 VDD1.n119 VSUBS 0.027794f
C376 VDD1.n120 VSUBS 0.014935f
C377 VDD1.n121 VSUBS 0.015814f
C378 VDD1.n122 VSUBS 0.035301f
C379 VDD1.n123 VSUBS 0.035301f
C380 VDD1.n124 VSUBS 0.015814f
C381 VDD1.n125 VSUBS 0.014935f
C382 VDD1.n126 VSUBS 0.027794f
C383 VDD1.n127 VSUBS 0.027794f
C384 VDD1.n128 VSUBS 0.014935f
C385 VDD1.n129 VSUBS 0.015814f
C386 VDD1.n130 VSUBS 0.035301f
C387 VDD1.n131 VSUBS 0.035301f
C388 VDD1.n132 VSUBS 0.015814f
C389 VDD1.n133 VSUBS 0.014935f
C390 VDD1.n134 VSUBS 0.027794f
C391 VDD1.n135 VSUBS 0.027794f
C392 VDD1.n136 VSUBS 0.014935f
C393 VDD1.n137 VSUBS 0.015814f
C394 VDD1.n138 VSUBS 0.035301f
C395 VDD1.n139 VSUBS 0.035301f
C396 VDD1.n140 VSUBS 0.015814f
C397 VDD1.n141 VSUBS 0.014935f
C398 VDD1.n142 VSUBS 0.027794f
C399 VDD1.n143 VSUBS 0.027794f
C400 VDD1.n144 VSUBS 0.014935f
C401 VDD1.n145 VSUBS 0.015814f
C402 VDD1.n146 VSUBS 0.035301f
C403 VDD1.n147 VSUBS 0.035301f
C404 VDD1.n148 VSUBS 0.015814f
C405 VDD1.n149 VSUBS 0.014935f
C406 VDD1.n150 VSUBS 0.027794f
C407 VDD1.n151 VSUBS 0.027794f
C408 VDD1.n152 VSUBS 0.014935f
C409 VDD1.n153 VSUBS 0.014935f
C410 VDD1.n154 VSUBS 0.015814f
C411 VDD1.n155 VSUBS 0.035301f
C412 VDD1.n156 VSUBS 0.035301f
C413 VDD1.n157 VSUBS 0.035301f
C414 VDD1.n158 VSUBS 0.015374f
C415 VDD1.n159 VSUBS 0.014935f
C416 VDD1.n160 VSUBS 0.027794f
C417 VDD1.n161 VSUBS 0.027794f
C418 VDD1.n162 VSUBS 0.014935f
C419 VDD1.n163 VSUBS 0.015814f
C420 VDD1.n164 VSUBS 0.035301f
C421 VDD1.n165 VSUBS 0.082657f
C422 VDD1.n166 VSUBS 0.015814f
C423 VDD1.n167 VSUBS 0.014935f
C424 VDD1.n168 VSUBS 0.068041f
C425 VDD1.n169 VSUBS 0.073359f
C426 VDD1.t4 VSUBS 0.339554f
C427 VDD1.t2 VSUBS 0.339554f
C428 VDD1.n170 VSUBS 2.78419f
C429 VDD1.n171 VSUBS 4.13576f
C430 VDD1.t1 VSUBS 0.339554f
C431 VDD1.t5 VSUBS 0.339554f
C432 VDD1.n172 VSUBS 2.77451f
C433 VDD1.n173 VSUBS 3.98453f
C434 VTAIL.t4 VSUBS 0.350689f
C435 VTAIL.t1 VSUBS 0.350689f
C436 VTAIL.n0 VSUBS 2.70358f
C437 VTAIL.n1 VSUBS 0.947577f
C438 VTAIL.n2 VSUBS 0.030691f
C439 VTAIL.n3 VSUBS 0.028705f
C440 VTAIL.n4 VSUBS 0.015425f
C441 VTAIL.n5 VSUBS 0.036459f
C442 VTAIL.n6 VSUBS 0.015879f
C443 VTAIL.n7 VSUBS 0.028705f
C444 VTAIL.n8 VSUBS 0.016332f
C445 VTAIL.n9 VSUBS 0.036459f
C446 VTAIL.n10 VSUBS 0.016332f
C447 VTAIL.n11 VSUBS 0.028705f
C448 VTAIL.n12 VSUBS 0.015425f
C449 VTAIL.n13 VSUBS 0.036459f
C450 VTAIL.n14 VSUBS 0.016332f
C451 VTAIL.n15 VSUBS 0.028705f
C452 VTAIL.n16 VSUBS 0.015425f
C453 VTAIL.n17 VSUBS 0.036459f
C454 VTAIL.n18 VSUBS 0.016332f
C455 VTAIL.n19 VSUBS 0.028705f
C456 VTAIL.n20 VSUBS 0.015425f
C457 VTAIL.n21 VSUBS 0.036459f
C458 VTAIL.n22 VSUBS 0.016332f
C459 VTAIL.n23 VSUBS 0.028705f
C460 VTAIL.n24 VSUBS 0.015425f
C461 VTAIL.n25 VSUBS 0.036459f
C462 VTAIL.n26 VSUBS 0.016332f
C463 VTAIL.n27 VSUBS 1.89282f
C464 VTAIL.n28 VSUBS 0.015425f
C465 VTAIL.t7 VSUBS 0.078084f
C466 VTAIL.n29 VSUBS 0.206241f
C467 VTAIL.n30 VSUBS 0.023193f
C468 VTAIL.n31 VSUBS 0.027344f
C469 VTAIL.n32 VSUBS 0.036459f
C470 VTAIL.n33 VSUBS 0.016332f
C471 VTAIL.n34 VSUBS 0.015425f
C472 VTAIL.n35 VSUBS 0.028705f
C473 VTAIL.n36 VSUBS 0.028705f
C474 VTAIL.n37 VSUBS 0.015425f
C475 VTAIL.n38 VSUBS 0.016332f
C476 VTAIL.n39 VSUBS 0.036459f
C477 VTAIL.n40 VSUBS 0.036459f
C478 VTAIL.n41 VSUBS 0.016332f
C479 VTAIL.n42 VSUBS 0.015425f
C480 VTAIL.n43 VSUBS 0.028705f
C481 VTAIL.n44 VSUBS 0.028705f
C482 VTAIL.n45 VSUBS 0.015425f
C483 VTAIL.n46 VSUBS 0.016332f
C484 VTAIL.n47 VSUBS 0.036459f
C485 VTAIL.n48 VSUBS 0.036459f
C486 VTAIL.n49 VSUBS 0.016332f
C487 VTAIL.n50 VSUBS 0.015425f
C488 VTAIL.n51 VSUBS 0.028705f
C489 VTAIL.n52 VSUBS 0.028705f
C490 VTAIL.n53 VSUBS 0.015425f
C491 VTAIL.n54 VSUBS 0.016332f
C492 VTAIL.n55 VSUBS 0.036459f
C493 VTAIL.n56 VSUBS 0.036459f
C494 VTAIL.n57 VSUBS 0.016332f
C495 VTAIL.n58 VSUBS 0.015425f
C496 VTAIL.n59 VSUBS 0.028705f
C497 VTAIL.n60 VSUBS 0.028705f
C498 VTAIL.n61 VSUBS 0.015425f
C499 VTAIL.n62 VSUBS 0.016332f
C500 VTAIL.n63 VSUBS 0.036459f
C501 VTAIL.n64 VSUBS 0.036459f
C502 VTAIL.n65 VSUBS 0.016332f
C503 VTAIL.n66 VSUBS 0.015425f
C504 VTAIL.n67 VSUBS 0.028705f
C505 VTAIL.n68 VSUBS 0.028705f
C506 VTAIL.n69 VSUBS 0.015425f
C507 VTAIL.n70 VSUBS 0.015425f
C508 VTAIL.n71 VSUBS 0.016332f
C509 VTAIL.n72 VSUBS 0.036459f
C510 VTAIL.n73 VSUBS 0.036459f
C511 VTAIL.n74 VSUBS 0.036459f
C512 VTAIL.n75 VSUBS 0.015879f
C513 VTAIL.n76 VSUBS 0.015425f
C514 VTAIL.n77 VSUBS 0.028705f
C515 VTAIL.n78 VSUBS 0.028705f
C516 VTAIL.n79 VSUBS 0.015425f
C517 VTAIL.n80 VSUBS 0.016332f
C518 VTAIL.n81 VSUBS 0.036459f
C519 VTAIL.n82 VSUBS 0.085367f
C520 VTAIL.n83 VSUBS 0.016332f
C521 VTAIL.n84 VSUBS 0.015425f
C522 VTAIL.n85 VSUBS 0.070272f
C523 VTAIL.n86 VSUBS 0.042919f
C524 VTAIL.n87 VSUBS 0.533059f
C525 VTAIL.t8 VSUBS 0.350689f
C526 VTAIL.t10 VSUBS 0.350689f
C527 VTAIL.n88 VSUBS 2.70358f
C528 VTAIL.n89 VSUBS 3.21569f
C529 VTAIL.t5 VSUBS 0.350689f
C530 VTAIL.t2 VSUBS 0.350689f
C531 VTAIL.n90 VSUBS 2.7036f
C532 VTAIL.n91 VSUBS 3.21568f
C533 VTAIL.n92 VSUBS 0.030691f
C534 VTAIL.n93 VSUBS 0.028705f
C535 VTAIL.n94 VSUBS 0.015425f
C536 VTAIL.n95 VSUBS 0.036459f
C537 VTAIL.n96 VSUBS 0.015879f
C538 VTAIL.n97 VSUBS 0.028705f
C539 VTAIL.n98 VSUBS 0.015879f
C540 VTAIL.n99 VSUBS 0.015425f
C541 VTAIL.n100 VSUBS 0.036459f
C542 VTAIL.n101 VSUBS 0.036459f
C543 VTAIL.n102 VSUBS 0.016332f
C544 VTAIL.n103 VSUBS 0.028705f
C545 VTAIL.n104 VSUBS 0.015425f
C546 VTAIL.n105 VSUBS 0.036459f
C547 VTAIL.n106 VSUBS 0.016332f
C548 VTAIL.n107 VSUBS 0.028705f
C549 VTAIL.n108 VSUBS 0.015425f
C550 VTAIL.n109 VSUBS 0.036459f
C551 VTAIL.n110 VSUBS 0.016332f
C552 VTAIL.n111 VSUBS 0.028705f
C553 VTAIL.n112 VSUBS 0.015425f
C554 VTAIL.n113 VSUBS 0.036459f
C555 VTAIL.n114 VSUBS 0.016332f
C556 VTAIL.n115 VSUBS 0.028705f
C557 VTAIL.n116 VSUBS 0.015425f
C558 VTAIL.n117 VSUBS 0.036459f
C559 VTAIL.n118 VSUBS 0.016332f
C560 VTAIL.n119 VSUBS 1.89282f
C561 VTAIL.n120 VSUBS 0.015425f
C562 VTAIL.t0 VSUBS 0.078084f
C563 VTAIL.n121 VSUBS 0.206241f
C564 VTAIL.n122 VSUBS 0.023193f
C565 VTAIL.n123 VSUBS 0.027344f
C566 VTAIL.n124 VSUBS 0.036459f
C567 VTAIL.n125 VSUBS 0.016332f
C568 VTAIL.n126 VSUBS 0.015425f
C569 VTAIL.n127 VSUBS 0.028705f
C570 VTAIL.n128 VSUBS 0.028705f
C571 VTAIL.n129 VSUBS 0.015425f
C572 VTAIL.n130 VSUBS 0.016332f
C573 VTAIL.n131 VSUBS 0.036459f
C574 VTAIL.n132 VSUBS 0.036459f
C575 VTAIL.n133 VSUBS 0.016332f
C576 VTAIL.n134 VSUBS 0.015425f
C577 VTAIL.n135 VSUBS 0.028705f
C578 VTAIL.n136 VSUBS 0.028705f
C579 VTAIL.n137 VSUBS 0.015425f
C580 VTAIL.n138 VSUBS 0.016332f
C581 VTAIL.n139 VSUBS 0.036459f
C582 VTAIL.n140 VSUBS 0.036459f
C583 VTAIL.n141 VSUBS 0.016332f
C584 VTAIL.n142 VSUBS 0.015425f
C585 VTAIL.n143 VSUBS 0.028705f
C586 VTAIL.n144 VSUBS 0.028705f
C587 VTAIL.n145 VSUBS 0.015425f
C588 VTAIL.n146 VSUBS 0.016332f
C589 VTAIL.n147 VSUBS 0.036459f
C590 VTAIL.n148 VSUBS 0.036459f
C591 VTAIL.n149 VSUBS 0.016332f
C592 VTAIL.n150 VSUBS 0.015425f
C593 VTAIL.n151 VSUBS 0.028705f
C594 VTAIL.n152 VSUBS 0.028705f
C595 VTAIL.n153 VSUBS 0.015425f
C596 VTAIL.n154 VSUBS 0.016332f
C597 VTAIL.n155 VSUBS 0.036459f
C598 VTAIL.n156 VSUBS 0.036459f
C599 VTAIL.n157 VSUBS 0.016332f
C600 VTAIL.n158 VSUBS 0.015425f
C601 VTAIL.n159 VSUBS 0.028705f
C602 VTAIL.n160 VSUBS 0.028705f
C603 VTAIL.n161 VSUBS 0.015425f
C604 VTAIL.n162 VSUBS 0.016332f
C605 VTAIL.n163 VSUBS 0.036459f
C606 VTAIL.n164 VSUBS 0.036459f
C607 VTAIL.n165 VSUBS 0.016332f
C608 VTAIL.n166 VSUBS 0.015425f
C609 VTAIL.n167 VSUBS 0.028705f
C610 VTAIL.n168 VSUBS 0.028705f
C611 VTAIL.n169 VSUBS 0.015425f
C612 VTAIL.n170 VSUBS 0.016332f
C613 VTAIL.n171 VSUBS 0.036459f
C614 VTAIL.n172 VSUBS 0.085367f
C615 VTAIL.n173 VSUBS 0.016332f
C616 VTAIL.n174 VSUBS 0.015425f
C617 VTAIL.n175 VSUBS 0.070272f
C618 VTAIL.n176 VSUBS 0.042919f
C619 VTAIL.n177 VSUBS 0.533059f
C620 VTAIL.t9 VSUBS 0.350689f
C621 VTAIL.t11 VSUBS 0.350689f
C622 VTAIL.n178 VSUBS 2.7036f
C623 VTAIL.n179 VSUBS 1.17361f
C624 VTAIL.n180 VSUBS 0.030691f
C625 VTAIL.n181 VSUBS 0.028705f
C626 VTAIL.n182 VSUBS 0.015425f
C627 VTAIL.n183 VSUBS 0.036459f
C628 VTAIL.n184 VSUBS 0.015879f
C629 VTAIL.n185 VSUBS 0.028705f
C630 VTAIL.n186 VSUBS 0.015879f
C631 VTAIL.n187 VSUBS 0.015425f
C632 VTAIL.n188 VSUBS 0.036459f
C633 VTAIL.n189 VSUBS 0.036459f
C634 VTAIL.n190 VSUBS 0.016332f
C635 VTAIL.n191 VSUBS 0.028705f
C636 VTAIL.n192 VSUBS 0.015425f
C637 VTAIL.n193 VSUBS 0.036459f
C638 VTAIL.n194 VSUBS 0.016332f
C639 VTAIL.n195 VSUBS 0.028705f
C640 VTAIL.n196 VSUBS 0.015425f
C641 VTAIL.n197 VSUBS 0.036459f
C642 VTAIL.n198 VSUBS 0.016332f
C643 VTAIL.n199 VSUBS 0.028705f
C644 VTAIL.n200 VSUBS 0.015425f
C645 VTAIL.n201 VSUBS 0.036459f
C646 VTAIL.n202 VSUBS 0.016332f
C647 VTAIL.n203 VSUBS 0.028705f
C648 VTAIL.n204 VSUBS 0.015425f
C649 VTAIL.n205 VSUBS 0.036459f
C650 VTAIL.n206 VSUBS 0.016332f
C651 VTAIL.n207 VSUBS 1.89282f
C652 VTAIL.n208 VSUBS 0.015425f
C653 VTAIL.t6 VSUBS 0.078084f
C654 VTAIL.n209 VSUBS 0.206241f
C655 VTAIL.n210 VSUBS 0.023193f
C656 VTAIL.n211 VSUBS 0.027344f
C657 VTAIL.n212 VSUBS 0.036459f
C658 VTAIL.n213 VSUBS 0.016332f
C659 VTAIL.n214 VSUBS 0.015425f
C660 VTAIL.n215 VSUBS 0.028705f
C661 VTAIL.n216 VSUBS 0.028705f
C662 VTAIL.n217 VSUBS 0.015425f
C663 VTAIL.n218 VSUBS 0.016332f
C664 VTAIL.n219 VSUBS 0.036459f
C665 VTAIL.n220 VSUBS 0.036459f
C666 VTAIL.n221 VSUBS 0.016332f
C667 VTAIL.n222 VSUBS 0.015425f
C668 VTAIL.n223 VSUBS 0.028705f
C669 VTAIL.n224 VSUBS 0.028705f
C670 VTAIL.n225 VSUBS 0.015425f
C671 VTAIL.n226 VSUBS 0.016332f
C672 VTAIL.n227 VSUBS 0.036459f
C673 VTAIL.n228 VSUBS 0.036459f
C674 VTAIL.n229 VSUBS 0.016332f
C675 VTAIL.n230 VSUBS 0.015425f
C676 VTAIL.n231 VSUBS 0.028705f
C677 VTAIL.n232 VSUBS 0.028705f
C678 VTAIL.n233 VSUBS 0.015425f
C679 VTAIL.n234 VSUBS 0.016332f
C680 VTAIL.n235 VSUBS 0.036459f
C681 VTAIL.n236 VSUBS 0.036459f
C682 VTAIL.n237 VSUBS 0.016332f
C683 VTAIL.n238 VSUBS 0.015425f
C684 VTAIL.n239 VSUBS 0.028705f
C685 VTAIL.n240 VSUBS 0.028705f
C686 VTAIL.n241 VSUBS 0.015425f
C687 VTAIL.n242 VSUBS 0.016332f
C688 VTAIL.n243 VSUBS 0.036459f
C689 VTAIL.n244 VSUBS 0.036459f
C690 VTAIL.n245 VSUBS 0.016332f
C691 VTAIL.n246 VSUBS 0.015425f
C692 VTAIL.n247 VSUBS 0.028705f
C693 VTAIL.n248 VSUBS 0.028705f
C694 VTAIL.n249 VSUBS 0.015425f
C695 VTAIL.n250 VSUBS 0.016332f
C696 VTAIL.n251 VSUBS 0.036459f
C697 VTAIL.n252 VSUBS 0.036459f
C698 VTAIL.n253 VSUBS 0.016332f
C699 VTAIL.n254 VSUBS 0.015425f
C700 VTAIL.n255 VSUBS 0.028705f
C701 VTAIL.n256 VSUBS 0.028705f
C702 VTAIL.n257 VSUBS 0.015425f
C703 VTAIL.n258 VSUBS 0.016332f
C704 VTAIL.n259 VSUBS 0.036459f
C705 VTAIL.n260 VSUBS 0.085367f
C706 VTAIL.n261 VSUBS 0.016332f
C707 VTAIL.n262 VSUBS 0.015425f
C708 VTAIL.n263 VSUBS 0.070272f
C709 VTAIL.n264 VSUBS 0.042919f
C710 VTAIL.n265 VSUBS 2.26654f
C711 VTAIL.n266 VSUBS 0.030691f
C712 VTAIL.n267 VSUBS 0.028705f
C713 VTAIL.n268 VSUBS 0.015425f
C714 VTAIL.n269 VSUBS 0.036459f
C715 VTAIL.n270 VSUBS 0.015879f
C716 VTAIL.n271 VSUBS 0.028705f
C717 VTAIL.n272 VSUBS 0.016332f
C718 VTAIL.n273 VSUBS 0.036459f
C719 VTAIL.n274 VSUBS 0.016332f
C720 VTAIL.n275 VSUBS 0.028705f
C721 VTAIL.n276 VSUBS 0.015425f
C722 VTAIL.n277 VSUBS 0.036459f
C723 VTAIL.n278 VSUBS 0.016332f
C724 VTAIL.n279 VSUBS 0.028705f
C725 VTAIL.n280 VSUBS 0.015425f
C726 VTAIL.n281 VSUBS 0.036459f
C727 VTAIL.n282 VSUBS 0.016332f
C728 VTAIL.n283 VSUBS 0.028705f
C729 VTAIL.n284 VSUBS 0.015425f
C730 VTAIL.n285 VSUBS 0.036459f
C731 VTAIL.n286 VSUBS 0.016332f
C732 VTAIL.n287 VSUBS 0.028705f
C733 VTAIL.n288 VSUBS 0.015425f
C734 VTAIL.n289 VSUBS 0.036459f
C735 VTAIL.n290 VSUBS 0.016332f
C736 VTAIL.n291 VSUBS 1.89282f
C737 VTAIL.n292 VSUBS 0.015425f
C738 VTAIL.t3 VSUBS 0.078084f
C739 VTAIL.n293 VSUBS 0.206241f
C740 VTAIL.n294 VSUBS 0.023193f
C741 VTAIL.n295 VSUBS 0.027344f
C742 VTAIL.n296 VSUBS 0.036459f
C743 VTAIL.n297 VSUBS 0.016332f
C744 VTAIL.n298 VSUBS 0.015425f
C745 VTAIL.n299 VSUBS 0.028705f
C746 VTAIL.n300 VSUBS 0.028705f
C747 VTAIL.n301 VSUBS 0.015425f
C748 VTAIL.n302 VSUBS 0.016332f
C749 VTAIL.n303 VSUBS 0.036459f
C750 VTAIL.n304 VSUBS 0.036459f
C751 VTAIL.n305 VSUBS 0.016332f
C752 VTAIL.n306 VSUBS 0.015425f
C753 VTAIL.n307 VSUBS 0.028705f
C754 VTAIL.n308 VSUBS 0.028705f
C755 VTAIL.n309 VSUBS 0.015425f
C756 VTAIL.n310 VSUBS 0.016332f
C757 VTAIL.n311 VSUBS 0.036459f
C758 VTAIL.n312 VSUBS 0.036459f
C759 VTAIL.n313 VSUBS 0.016332f
C760 VTAIL.n314 VSUBS 0.015425f
C761 VTAIL.n315 VSUBS 0.028705f
C762 VTAIL.n316 VSUBS 0.028705f
C763 VTAIL.n317 VSUBS 0.015425f
C764 VTAIL.n318 VSUBS 0.016332f
C765 VTAIL.n319 VSUBS 0.036459f
C766 VTAIL.n320 VSUBS 0.036459f
C767 VTAIL.n321 VSUBS 0.016332f
C768 VTAIL.n322 VSUBS 0.015425f
C769 VTAIL.n323 VSUBS 0.028705f
C770 VTAIL.n324 VSUBS 0.028705f
C771 VTAIL.n325 VSUBS 0.015425f
C772 VTAIL.n326 VSUBS 0.016332f
C773 VTAIL.n327 VSUBS 0.036459f
C774 VTAIL.n328 VSUBS 0.036459f
C775 VTAIL.n329 VSUBS 0.016332f
C776 VTAIL.n330 VSUBS 0.015425f
C777 VTAIL.n331 VSUBS 0.028705f
C778 VTAIL.n332 VSUBS 0.028705f
C779 VTAIL.n333 VSUBS 0.015425f
C780 VTAIL.n334 VSUBS 0.015425f
C781 VTAIL.n335 VSUBS 0.016332f
C782 VTAIL.n336 VSUBS 0.036459f
C783 VTAIL.n337 VSUBS 0.036459f
C784 VTAIL.n338 VSUBS 0.036459f
C785 VTAIL.n339 VSUBS 0.015879f
C786 VTAIL.n340 VSUBS 0.015425f
C787 VTAIL.n341 VSUBS 0.028705f
C788 VTAIL.n342 VSUBS 0.028705f
C789 VTAIL.n343 VSUBS 0.015425f
C790 VTAIL.n344 VSUBS 0.016332f
C791 VTAIL.n345 VSUBS 0.036459f
C792 VTAIL.n346 VSUBS 0.085367f
C793 VTAIL.n347 VSUBS 0.016332f
C794 VTAIL.n348 VSUBS 0.015425f
C795 VTAIL.n349 VSUBS 0.070272f
C796 VTAIL.n350 VSUBS 0.042919f
C797 VTAIL.n351 VSUBS 2.18402f
C798 VP.t3 VSUBS 3.91079f
C799 VP.n0 VSUBS 1.45104f
C800 VP.n1 VSUBS 0.02606f
C801 VP.n2 VSUBS 0.042569f
C802 VP.n3 VSUBS 0.02606f
C803 VP.n4 VSUBS 0.036397f
C804 VP.n5 VSUBS 0.02606f
C805 VP.n6 VSUBS 0.033196f
C806 VP.n7 VSUBS 0.02606f
C807 VP.n8 VSUBS 0.030195f
C808 VP.t0 VSUBS 3.91079f
C809 VP.n9 VSUBS 1.45104f
C810 VP.n10 VSUBS 0.02606f
C811 VP.n11 VSUBS 0.042569f
C812 VP.n12 VSUBS 0.02606f
C813 VP.n13 VSUBS 0.036397f
C814 VP.t5 VSUBS 4.27818f
C815 VP.t4 VSUBS 3.91079f
C816 VP.n14 VSUBS 1.44537f
C817 VP.n15 VSUBS 1.38047f
C818 VP.n16 VSUBS 0.324633f
C819 VP.n17 VSUBS 0.02606f
C820 VP.n18 VSUBS 0.048326f
C821 VP.n19 VSUBS 0.048326f
C822 VP.n20 VSUBS 0.033196f
C823 VP.n21 VSUBS 0.02606f
C824 VP.n22 VSUBS 0.02606f
C825 VP.n23 VSUBS 0.02606f
C826 VP.n24 VSUBS 0.048326f
C827 VP.n25 VSUBS 0.048326f
C828 VP.n26 VSUBS 0.030195f
C829 VP.n27 VSUBS 0.042054f
C830 VP.n28 VSUBS 1.70611f
C831 VP.t2 VSUBS 3.91079f
C832 VP.n29 VSUBS 1.45104f
C833 VP.n30 VSUBS 1.72319f
C834 VP.n31 VSUBS 0.042054f
C835 VP.n32 VSUBS 0.02606f
C836 VP.n33 VSUBS 0.048326f
C837 VP.n34 VSUBS 0.048326f
C838 VP.n35 VSUBS 0.042569f
C839 VP.n36 VSUBS 0.02606f
C840 VP.n37 VSUBS 0.02606f
C841 VP.n38 VSUBS 0.02606f
C842 VP.n39 VSUBS 0.048326f
C843 VP.n40 VSUBS 0.048326f
C844 VP.t1 VSUBS 3.91079f
C845 VP.n41 VSUBS 1.35618f
C846 VP.n42 VSUBS 0.036397f
C847 VP.n43 VSUBS 0.02606f
C848 VP.n44 VSUBS 0.02606f
C849 VP.n45 VSUBS 0.02606f
C850 VP.n46 VSUBS 0.048326f
C851 VP.n47 VSUBS 0.048326f
C852 VP.n48 VSUBS 0.033196f
C853 VP.n49 VSUBS 0.02606f
C854 VP.n50 VSUBS 0.02606f
C855 VP.n51 VSUBS 0.02606f
C856 VP.n52 VSUBS 0.048326f
C857 VP.n53 VSUBS 0.048326f
C858 VP.n54 VSUBS 0.030195f
C859 VP.n55 VSUBS 0.042054f
C860 VP.n56 VSUBS 0.073963f
C861 B.n0 VSUBS 0.006773f
C862 B.n1 VSUBS 0.006773f
C863 B.n2 VSUBS 0.010017f
C864 B.n3 VSUBS 0.007676f
C865 B.n4 VSUBS 0.007676f
C866 B.n5 VSUBS 0.007676f
C867 B.n6 VSUBS 0.007676f
C868 B.n7 VSUBS 0.007676f
C869 B.n8 VSUBS 0.007676f
C870 B.n9 VSUBS 0.007676f
C871 B.n10 VSUBS 0.007676f
C872 B.n11 VSUBS 0.007676f
C873 B.n12 VSUBS 0.007676f
C874 B.n13 VSUBS 0.007676f
C875 B.n14 VSUBS 0.007676f
C876 B.n15 VSUBS 0.007676f
C877 B.n16 VSUBS 0.007676f
C878 B.n17 VSUBS 0.007676f
C879 B.n18 VSUBS 0.007676f
C880 B.n19 VSUBS 0.007676f
C881 B.n20 VSUBS 0.007676f
C882 B.n21 VSUBS 0.007676f
C883 B.n22 VSUBS 0.007676f
C884 B.n23 VSUBS 0.007676f
C885 B.n24 VSUBS 0.007676f
C886 B.n25 VSUBS 0.007676f
C887 B.n26 VSUBS 0.007676f
C888 B.n27 VSUBS 0.007676f
C889 B.n28 VSUBS 0.018293f
C890 B.n29 VSUBS 0.007676f
C891 B.n30 VSUBS 0.007676f
C892 B.n31 VSUBS 0.007676f
C893 B.n32 VSUBS 0.007676f
C894 B.n33 VSUBS 0.007676f
C895 B.n34 VSUBS 0.007676f
C896 B.n35 VSUBS 0.007676f
C897 B.n36 VSUBS 0.007676f
C898 B.n37 VSUBS 0.007676f
C899 B.n38 VSUBS 0.007676f
C900 B.n39 VSUBS 0.007676f
C901 B.n40 VSUBS 0.007676f
C902 B.n41 VSUBS 0.007676f
C903 B.n42 VSUBS 0.007676f
C904 B.n43 VSUBS 0.007676f
C905 B.n44 VSUBS 0.007676f
C906 B.n45 VSUBS 0.007676f
C907 B.n46 VSUBS 0.007676f
C908 B.n47 VSUBS 0.007676f
C909 B.n48 VSUBS 0.007676f
C910 B.n49 VSUBS 0.007676f
C911 B.n50 VSUBS 0.007676f
C912 B.n51 VSUBS 0.007676f
C913 B.n52 VSUBS 0.007676f
C914 B.n53 VSUBS 0.007676f
C915 B.n54 VSUBS 0.005306f
C916 B.n55 VSUBS 0.007676f
C917 B.t1 VSUBS 0.318453f
C918 B.t2 VSUBS 0.365216f
C919 B.t0 VSUBS 2.74739f
C920 B.n56 VSUBS 0.580296f
C921 B.n57 VSUBS 0.330568f
C922 B.n58 VSUBS 0.017785f
C923 B.n59 VSUBS 0.007676f
C924 B.n60 VSUBS 0.007676f
C925 B.n61 VSUBS 0.007676f
C926 B.n62 VSUBS 0.007676f
C927 B.t10 VSUBS 0.318457f
C928 B.t11 VSUBS 0.36522f
C929 B.t9 VSUBS 2.74739f
C930 B.n63 VSUBS 0.580293f
C931 B.n64 VSUBS 0.330564f
C932 B.n65 VSUBS 0.007676f
C933 B.n66 VSUBS 0.007676f
C934 B.n67 VSUBS 0.007676f
C935 B.n68 VSUBS 0.007676f
C936 B.n69 VSUBS 0.007676f
C937 B.n70 VSUBS 0.007676f
C938 B.n71 VSUBS 0.007676f
C939 B.n72 VSUBS 0.007676f
C940 B.n73 VSUBS 0.007676f
C941 B.n74 VSUBS 0.007676f
C942 B.n75 VSUBS 0.007676f
C943 B.n76 VSUBS 0.007676f
C944 B.n77 VSUBS 0.007676f
C945 B.n78 VSUBS 0.007676f
C946 B.n79 VSUBS 0.007676f
C947 B.n80 VSUBS 0.007676f
C948 B.n81 VSUBS 0.007676f
C949 B.n82 VSUBS 0.007676f
C950 B.n83 VSUBS 0.007676f
C951 B.n84 VSUBS 0.007676f
C952 B.n85 VSUBS 0.007676f
C953 B.n86 VSUBS 0.007676f
C954 B.n87 VSUBS 0.007676f
C955 B.n88 VSUBS 0.007676f
C956 B.n89 VSUBS 0.007676f
C957 B.n90 VSUBS 0.018293f
C958 B.n91 VSUBS 0.007676f
C959 B.n92 VSUBS 0.007676f
C960 B.n93 VSUBS 0.007676f
C961 B.n94 VSUBS 0.007676f
C962 B.n95 VSUBS 0.007676f
C963 B.n96 VSUBS 0.007676f
C964 B.n97 VSUBS 0.007676f
C965 B.n98 VSUBS 0.007676f
C966 B.n99 VSUBS 0.007676f
C967 B.n100 VSUBS 0.007676f
C968 B.n101 VSUBS 0.007676f
C969 B.n102 VSUBS 0.007676f
C970 B.n103 VSUBS 0.007676f
C971 B.n104 VSUBS 0.007676f
C972 B.n105 VSUBS 0.007676f
C973 B.n106 VSUBS 0.007676f
C974 B.n107 VSUBS 0.007676f
C975 B.n108 VSUBS 0.007676f
C976 B.n109 VSUBS 0.007676f
C977 B.n110 VSUBS 0.007676f
C978 B.n111 VSUBS 0.007676f
C979 B.n112 VSUBS 0.007676f
C980 B.n113 VSUBS 0.007676f
C981 B.n114 VSUBS 0.007676f
C982 B.n115 VSUBS 0.007676f
C983 B.n116 VSUBS 0.007676f
C984 B.n117 VSUBS 0.007676f
C985 B.n118 VSUBS 0.007676f
C986 B.n119 VSUBS 0.007676f
C987 B.n120 VSUBS 0.007676f
C988 B.n121 VSUBS 0.007676f
C989 B.n122 VSUBS 0.007676f
C990 B.n123 VSUBS 0.007676f
C991 B.n124 VSUBS 0.007676f
C992 B.n125 VSUBS 0.007676f
C993 B.n126 VSUBS 0.007676f
C994 B.n127 VSUBS 0.007676f
C995 B.n128 VSUBS 0.007676f
C996 B.n129 VSUBS 0.007676f
C997 B.n130 VSUBS 0.007676f
C998 B.n131 VSUBS 0.007676f
C999 B.n132 VSUBS 0.007676f
C1000 B.n133 VSUBS 0.007676f
C1001 B.n134 VSUBS 0.007676f
C1002 B.n135 VSUBS 0.007676f
C1003 B.n136 VSUBS 0.007676f
C1004 B.n137 VSUBS 0.007676f
C1005 B.n138 VSUBS 0.007676f
C1006 B.n139 VSUBS 0.007676f
C1007 B.n140 VSUBS 0.007676f
C1008 B.n141 VSUBS 0.007676f
C1009 B.n142 VSUBS 0.007676f
C1010 B.n143 VSUBS 0.007676f
C1011 B.n144 VSUBS 0.019185f
C1012 B.n145 VSUBS 0.007676f
C1013 B.n146 VSUBS 0.007676f
C1014 B.n147 VSUBS 0.007676f
C1015 B.n148 VSUBS 0.007676f
C1016 B.n149 VSUBS 0.007676f
C1017 B.n150 VSUBS 0.007676f
C1018 B.n151 VSUBS 0.007676f
C1019 B.n152 VSUBS 0.007676f
C1020 B.n153 VSUBS 0.007676f
C1021 B.n154 VSUBS 0.007676f
C1022 B.n155 VSUBS 0.007676f
C1023 B.n156 VSUBS 0.007676f
C1024 B.n157 VSUBS 0.007676f
C1025 B.n158 VSUBS 0.007676f
C1026 B.n159 VSUBS 0.007676f
C1027 B.n160 VSUBS 0.007676f
C1028 B.n161 VSUBS 0.007676f
C1029 B.n162 VSUBS 0.007676f
C1030 B.n163 VSUBS 0.007676f
C1031 B.n164 VSUBS 0.007676f
C1032 B.n165 VSUBS 0.007676f
C1033 B.n166 VSUBS 0.007676f
C1034 B.n167 VSUBS 0.007676f
C1035 B.n168 VSUBS 0.007676f
C1036 B.n169 VSUBS 0.007676f
C1037 B.n170 VSUBS 0.007676f
C1038 B.t8 VSUBS 0.318457f
C1039 B.t7 VSUBS 0.36522f
C1040 B.t6 VSUBS 2.74739f
C1041 B.n171 VSUBS 0.580293f
C1042 B.n172 VSUBS 0.330564f
C1043 B.n173 VSUBS 0.007676f
C1044 B.n174 VSUBS 0.007676f
C1045 B.n175 VSUBS 0.007676f
C1046 B.n176 VSUBS 0.007676f
C1047 B.t5 VSUBS 0.318453f
C1048 B.t4 VSUBS 0.365216f
C1049 B.t3 VSUBS 2.74739f
C1050 B.n177 VSUBS 0.580296f
C1051 B.n178 VSUBS 0.330568f
C1052 B.n179 VSUBS 0.007676f
C1053 B.n180 VSUBS 0.007676f
C1054 B.n181 VSUBS 0.007676f
C1055 B.n182 VSUBS 0.007676f
C1056 B.n183 VSUBS 0.007676f
C1057 B.n184 VSUBS 0.007676f
C1058 B.n185 VSUBS 0.007676f
C1059 B.n186 VSUBS 0.007676f
C1060 B.n187 VSUBS 0.007676f
C1061 B.n188 VSUBS 0.007676f
C1062 B.n189 VSUBS 0.007676f
C1063 B.n190 VSUBS 0.007676f
C1064 B.n191 VSUBS 0.007676f
C1065 B.n192 VSUBS 0.007676f
C1066 B.n193 VSUBS 0.007676f
C1067 B.n194 VSUBS 0.007676f
C1068 B.n195 VSUBS 0.007676f
C1069 B.n196 VSUBS 0.007676f
C1070 B.n197 VSUBS 0.007676f
C1071 B.n198 VSUBS 0.007676f
C1072 B.n199 VSUBS 0.007676f
C1073 B.n200 VSUBS 0.007676f
C1074 B.n201 VSUBS 0.007676f
C1075 B.n202 VSUBS 0.007676f
C1076 B.n203 VSUBS 0.007676f
C1077 B.n204 VSUBS 0.019185f
C1078 B.n205 VSUBS 0.007676f
C1079 B.n206 VSUBS 0.007676f
C1080 B.n207 VSUBS 0.007676f
C1081 B.n208 VSUBS 0.007676f
C1082 B.n209 VSUBS 0.007676f
C1083 B.n210 VSUBS 0.007676f
C1084 B.n211 VSUBS 0.007676f
C1085 B.n212 VSUBS 0.007676f
C1086 B.n213 VSUBS 0.007676f
C1087 B.n214 VSUBS 0.007676f
C1088 B.n215 VSUBS 0.007676f
C1089 B.n216 VSUBS 0.007676f
C1090 B.n217 VSUBS 0.007676f
C1091 B.n218 VSUBS 0.007676f
C1092 B.n219 VSUBS 0.007676f
C1093 B.n220 VSUBS 0.007676f
C1094 B.n221 VSUBS 0.007676f
C1095 B.n222 VSUBS 0.007676f
C1096 B.n223 VSUBS 0.007676f
C1097 B.n224 VSUBS 0.007676f
C1098 B.n225 VSUBS 0.007676f
C1099 B.n226 VSUBS 0.007676f
C1100 B.n227 VSUBS 0.007676f
C1101 B.n228 VSUBS 0.007676f
C1102 B.n229 VSUBS 0.007676f
C1103 B.n230 VSUBS 0.007676f
C1104 B.n231 VSUBS 0.007676f
C1105 B.n232 VSUBS 0.007676f
C1106 B.n233 VSUBS 0.007676f
C1107 B.n234 VSUBS 0.007676f
C1108 B.n235 VSUBS 0.007676f
C1109 B.n236 VSUBS 0.007676f
C1110 B.n237 VSUBS 0.007676f
C1111 B.n238 VSUBS 0.007676f
C1112 B.n239 VSUBS 0.007676f
C1113 B.n240 VSUBS 0.007676f
C1114 B.n241 VSUBS 0.007676f
C1115 B.n242 VSUBS 0.007676f
C1116 B.n243 VSUBS 0.007676f
C1117 B.n244 VSUBS 0.007676f
C1118 B.n245 VSUBS 0.007676f
C1119 B.n246 VSUBS 0.007676f
C1120 B.n247 VSUBS 0.007676f
C1121 B.n248 VSUBS 0.007676f
C1122 B.n249 VSUBS 0.007676f
C1123 B.n250 VSUBS 0.007676f
C1124 B.n251 VSUBS 0.007676f
C1125 B.n252 VSUBS 0.007676f
C1126 B.n253 VSUBS 0.007676f
C1127 B.n254 VSUBS 0.007676f
C1128 B.n255 VSUBS 0.007676f
C1129 B.n256 VSUBS 0.007676f
C1130 B.n257 VSUBS 0.007676f
C1131 B.n258 VSUBS 0.007676f
C1132 B.n259 VSUBS 0.007676f
C1133 B.n260 VSUBS 0.007676f
C1134 B.n261 VSUBS 0.007676f
C1135 B.n262 VSUBS 0.007676f
C1136 B.n263 VSUBS 0.007676f
C1137 B.n264 VSUBS 0.007676f
C1138 B.n265 VSUBS 0.007676f
C1139 B.n266 VSUBS 0.007676f
C1140 B.n267 VSUBS 0.007676f
C1141 B.n268 VSUBS 0.007676f
C1142 B.n269 VSUBS 0.007676f
C1143 B.n270 VSUBS 0.007676f
C1144 B.n271 VSUBS 0.007676f
C1145 B.n272 VSUBS 0.007676f
C1146 B.n273 VSUBS 0.007676f
C1147 B.n274 VSUBS 0.007676f
C1148 B.n275 VSUBS 0.007676f
C1149 B.n276 VSUBS 0.007676f
C1150 B.n277 VSUBS 0.007676f
C1151 B.n278 VSUBS 0.007676f
C1152 B.n279 VSUBS 0.007676f
C1153 B.n280 VSUBS 0.007676f
C1154 B.n281 VSUBS 0.007676f
C1155 B.n282 VSUBS 0.007676f
C1156 B.n283 VSUBS 0.007676f
C1157 B.n284 VSUBS 0.007676f
C1158 B.n285 VSUBS 0.007676f
C1159 B.n286 VSUBS 0.007676f
C1160 B.n287 VSUBS 0.007676f
C1161 B.n288 VSUBS 0.007676f
C1162 B.n289 VSUBS 0.007676f
C1163 B.n290 VSUBS 0.007676f
C1164 B.n291 VSUBS 0.007676f
C1165 B.n292 VSUBS 0.007676f
C1166 B.n293 VSUBS 0.007676f
C1167 B.n294 VSUBS 0.007676f
C1168 B.n295 VSUBS 0.007676f
C1169 B.n296 VSUBS 0.007676f
C1170 B.n297 VSUBS 0.007676f
C1171 B.n298 VSUBS 0.007676f
C1172 B.n299 VSUBS 0.007676f
C1173 B.n300 VSUBS 0.007676f
C1174 B.n301 VSUBS 0.007676f
C1175 B.n302 VSUBS 0.007676f
C1176 B.n303 VSUBS 0.007676f
C1177 B.n304 VSUBS 0.007676f
C1178 B.n305 VSUBS 0.007676f
C1179 B.n306 VSUBS 0.007676f
C1180 B.n307 VSUBS 0.018293f
C1181 B.n308 VSUBS 0.018293f
C1182 B.n309 VSUBS 0.019185f
C1183 B.n310 VSUBS 0.007676f
C1184 B.n311 VSUBS 0.007676f
C1185 B.n312 VSUBS 0.007676f
C1186 B.n313 VSUBS 0.007676f
C1187 B.n314 VSUBS 0.007676f
C1188 B.n315 VSUBS 0.007676f
C1189 B.n316 VSUBS 0.007676f
C1190 B.n317 VSUBS 0.007676f
C1191 B.n318 VSUBS 0.007676f
C1192 B.n319 VSUBS 0.007676f
C1193 B.n320 VSUBS 0.007676f
C1194 B.n321 VSUBS 0.007676f
C1195 B.n322 VSUBS 0.007676f
C1196 B.n323 VSUBS 0.007676f
C1197 B.n324 VSUBS 0.007676f
C1198 B.n325 VSUBS 0.007676f
C1199 B.n326 VSUBS 0.007676f
C1200 B.n327 VSUBS 0.007676f
C1201 B.n328 VSUBS 0.007676f
C1202 B.n329 VSUBS 0.007676f
C1203 B.n330 VSUBS 0.007676f
C1204 B.n331 VSUBS 0.007676f
C1205 B.n332 VSUBS 0.007676f
C1206 B.n333 VSUBS 0.007676f
C1207 B.n334 VSUBS 0.007676f
C1208 B.n335 VSUBS 0.007676f
C1209 B.n336 VSUBS 0.007676f
C1210 B.n337 VSUBS 0.007676f
C1211 B.n338 VSUBS 0.007676f
C1212 B.n339 VSUBS 0.007676f
C1213 B.n340 VSUBS 0.007676f
C1214 B.n341 VSUBS 0.007676f
C1215 B.n342 VSUBS 0.007676f
C1216 B.n343 VSUBS 0.007676f
C1217 B.n344 VSUBS 0.007676f
C1218 B.n345 VSUBS 0.007676f
C1219 B.n346 VSUBS 0.007676f
C1220 B.n347 VSUBS 0.007676f
C1221 B.n348 VSUBS 0.007676f
C1222 B.n349 VSUBS 0.007676f
C1223 B.n350 VSUBS 0.007676f
C1224 B.n351 VSUBS 0.007676f
C1225 B.n352 VSUBS 0.007676f
C1226 B.n353 VSUBS 0.007676f
C1227 B.n354 VSUBS 0.007676f
C1228 B.n355 VSUBS 0.007676f
C1229 B.n356 VSUBS 0.007676f
C1230 B.n357 VSUBS 0.007676f
C1231 B.n358 VSUBS 0.007676f
C1232 B.n359 VSUBS 0.007676f
C1233 B.n360 VSUBS 0.007676f
C1234 B.n361 VSUBS 0.007676f
C1235 B.n362 VSUBS 0.007676f
C1236 B.n363 VSUBS 0.007676f
C1237 B.n364 VSUBS 0.007676f
C1238 B.n365 VSUBS 0.007676f
C1239 B.n366 VSUBS 0.007676f
C1240 B.n367 VSUBS 0.007676f
C1241 B.n368 VSUBS 0.007676f
C1242 B.n369 VSUBS 0.007676f
C1243 B.n370 VSUBS 0.007676f
C1244 B.n371 VSUBS 0.007676f
C1245 B.n372 VSUBS 0.007676f
C1246 B.n373 VSUBS 0.007676f
C1247 B.n374 VSUBS 0.007676f
C1248 B.n375 VSUBS 0.007676f
C1249 B.n376 VSUBS 0.007676f
C1250 B.n377 VSUBS 0.007676f
C1251 B.n378 VSUBS 0.007676f
C1252 B.n379 VSUBS 0.007676f
C1253 B.n380 VSUBS 0.007676f
C1254 B.n381 VSUBS 0.007676f
C1255 B.n382 VSUBS 0.007676f
C1256 B.n383 VSUBS 0.007676f
C1257 B.n384 VSUBS 0.007676f
C1258 B.n385 VSUBS 0.007676f
C1259 B.n386 VSUBS 0.005306f
C1260 B.n387 VSUBS 0.017785f
C1261 B.n388 VSUBS 0.006209f
C1262 B.n389 VSUBS 0.007676f
C1263 B.n390 VSUBS 0.007676f
C1264 B.n391 VSUBS 0.007676f
C1265 B.n392 VSUBS 0.007676f
C1266 B.n393 VSUBS 0.007676f
C1267 B.n394 VSUBS 0.007676f
C1268 B.n395 VSUBS 0.007676f
C1269 B.n396 VSUBS 0.007676f
C1270 B.n397 VSUBS 0.007676f
C1271 B.n398 VSUBS 0.007676f
C1272 B.n399 VSUBS 0.007676f
C1273 B.n400 VSUBS 0.006209f
C1274 B.n401 VSUBS 0.017785f
C1275 B.n402 VSUBS 0.005306f
C1276 B.n403 VSUBS 0.007676f
C1277 B.n404 VSUBS 0.007676f
C1278 B.n405 VSUBS 0.007676f
C1279 B.n406 VSUBS 0.007676f
C1280 B.n407 VSUBS 0.007676f
C1281 B.n408 VSUBS 0.007676f
C1282 B.n409 VSUBS 0.007676f
C1283 B.n410 VSUBS 0.007676f
C1284 B.n411 VSUBS 0.007676f
C1285 B.n412 VSUBS 0.007676f
C1286 B.n413 VSUBS 0.007676f
C1287 B.n414 VSUBS 0.007676f
C1288 B.n415 VSUBS 0.007676f
C1289 B.n416 VSUBS 0.007676f
C1290 B.n417 VSUBS 0.007676f
C1291 B.n418 VSUBS 0.007676f
C1292 B.n419 VSUBS 0.007676f
C1293 B.n420 VSUBS 0.007676f
C1294 B.n421 VSUBS 0.007676f
C1295 B.n422 VSUBS 0.007676f
C1296 B.n423 VSUBS 0.007676f
C1297 B.n424 VSUBS 0.007676f
C1298 B.n425 VSUBS 0.007676f
C1299 B.n426 VSUBS 0.007676f
C1300 B.n427 VSUBS 0.007676f
C1301 B.n428 VSUBS 0.007676f
C1302 B.n429 VSUBS 0.007676f
C1303 B.n430 VSUBS 0.007676f
C1304 B.n431 VSUBS 0.007676f
C1305 B.n432 VSUBS 0.007676f
C1306 B.n433 VSUBS 0.007676f
C1307 B.n434 VSUBS 0.007676f
C1308 B.n435 VSUBS 0.007676f
C1309 B.n436 VSUBS 0.007676f
C1310 B.n437 VSUBS 0.007676f
C1311 B.n438 VSUBS 0.007676f
C1312 B.n439 VSUBS 0.007676f
C1313 B.n440 VSUBS 0.007676f
C1314 B.n441 VSUBS 0.007676f
C1315 B.n442 VSUBS 0.007676f
C1316 B.n443 VSUBS 0.007676f
C1317 B.n444 VSUBS 0.007676f
C1318 B.n445 VSUBS 0.007676f
C1319 B.n446 VSUBS 0.007676f
C1320 B.n447 VSUBS 0.007676f
C1321 B.n448 VSUBS 0.007676f
C1322 B.n449 VSUBS 0.007676f
C1323 B.n450 VSUBS 0.007676f
C1324 B.n451 VSUBS 0.007676f
C1325 B.n452 VSUBS 0.007676f
C1326 B.n453 VSUBS 0.007676f
C1327 B.n454 VSUBS 0.007676f
C1328 B.n455 VSUBS 0.007676f
C1329 B.n456 VSUBS 0.007676f
C1330 B.n457 VSUBS 0.007676f
C1331 B.n458 VSUBS 0.007676f
C1332 B.n459 VSUBS 0.007676f
C1333 B.n460 VSUBS 0.007676f
C1334 B.n461 VSUBS 0.007676f
C1335 B.n462 VSUBS 0.007676f
C1336 B.n463 VSUBS 0.007676f
C1337 B.n464 VSUBS 0.007676f
C1338 B.n465 VSUBS 0.007676f
C1339 B.n466 VSUBS 0.007676f
C1340 B.n467 VSUBS 0.007676f
C1341 B.n468 VSUBS 0.007676f
C1342 B.n469 VSUBS 0.007676f
C1343 B.n470 VSUBS 0.007676f
C1344 B.n471 VSUBS 0.007676f
C1345 B.n472 VSUBS 0.007676f
C1346 B.n473 VSUBS 0.007676f
C1347 B.n474 VSUBS 0.007676f
C1348 B.n475 VSUBS 0.007676f
C1349 B.n476 VSUBS 0.007676f
C1350 B.n477 VSUBS 0.007676f
C1351 B.n478 VSUBS 0.007676f
C1352 B.n479 VSUBS 0.018334f
C1353 B.n480 VSUBS 0.019144f
C1354 B.n481 VSUBS 0.018293f
C1355 B.n482 VSUBS 0.007676f
C1356 B.n483 VSUBS 0.007676f
C1357 B.n484 VSUBS 0.007676f
C1358 B.n485 VSUBS 0.007676f
C1359 B.n486 VSUBS 0.007676f
C1360 B.n487 VSUBS 0.007676f
C1361 B.n488 VSUBS 0.007676f
C1362 B.n489 VSUBS 0.007676f
C1363 B.n490 VSUBS 0.007676f
C1364 B.n491 VSUBS 0.007676f
C1365 B.n492 VSUBS 0.007676f
C1366 B.n493 VSUBS 0.007676f
C1367 B.n494 VSUBS 0.007676f
C1368 B.n495 VSUBS 0.007676f
C1369 B.n496 VSUBS 0.007676f
C1370 B.n497 VSUBS 0.007676f
C1371 B.n498 VSUBS 0.007676f
C1372 B.n499 VSUBS 0.007676f
C1373 B.n500 VSUBS 0.007676f
C1374 B.n501 VSUBS 0.007676f
C1375 B.n502 VSUBS 0.007676f
C1376 B.n503 VSUBS 0.007676f
C1377 B.n504 VSUBS 0.007676f
C1378 B.n505 VSUBS 0.007676f
C1379 B.n506 VSUBS 0.007676f
C1380 B.n507 VSUBS 0.007676f
C1381 B.n508 VSUBS 0.007676f
C1382 B.n509 VSUBS 0.007676f
C1383 B.n510 VSUBS 0.007676f
C1384 B.n511 VSUBS 0.007676f
C1385 B.n512 VSUBS 0.007676f
C1386 B.n513 VSUBS 0.007676f
C1387 B.n514 VSUBS 0.007676f
C1388 B.n515 VSUBS 0.007676f
C1389 B.n516 VSUBS 0.007676f
C1390 B.n517 VSUBS 0.007676f
C1391 B.n518 VSUBS 0.007676f
C1392 B.n519 VSUBS 0.007676f
C1393 B.n520 VSUBS 0.007676f
C1394 B.n521 VSUBS 0.007676f
C1395 B.n522 VSUBS 0.007676f
C1396 B.n523 VSUBS 0.007676f
C1397 B.n524 VSUBS 0.007676f
C1398 B.n525 VSUBS 0.007676f
C1399 B.n526 VSUBS 0.007676f
C1400 B.n527 VSUBS 0.007676f
C1401 B.n528 VSUBS 0.007676f
C1402 B.n529 VSUBS 0.007676f
C1403 B.n530 VSUBS 0.007676f
C1404 B.n531 VSUBS 0.007676f
C1405 B.n532 VSUBS 0.007676f
C1406 B.n533 VSUBS 0.007676f
C1407 B.n534 VSUBS 0.007676f
C1408 B.n535 VSUBS 0.007676f
C1409 B.n536 VSUBS 0.007676f
C1410 B.n537 VSUBS 0.007676f
C1411 B.n538 VSUBS 0.007676f
C1412 B.n539 VSUBS 0.007676f
C1413 B.n540 VSUBS 0.007676f
C1414 B.n541 VSUBS 0.007676f
C1415 B.n542 VSUBS 0.007676f
C1416 B.n543 VSUBS 0.007676f
C1417 B.n544 VSUBS 0.007676f
C1418 B.n545 VSUBS 0.007676f
C1419 B.n546 VSUBS 0.007676f
C1420 B.n547 VSUBS 0.007676f
C1421 B.n548 VSUBS 0.007676f
C1422 B.n549 VSUBS 0.007676f
C1423 B.n550 VSUBS 0.007676f
C1424 B.n551 VSUBS 0.007676f
C1425 B.n552 VSUBS 0.007676f
C1426 B.n553 VSUBS 0.007676f
C1427 B.n554 VSUBS 0.007676f
C1428 B.n555 VSUBS 0.007676f
C1429 B.n556 VSUBS 0.007676f
C1430 B.n557 VSUBS 0.007676f
C1431 B.n558 VSUBS 0.007676f
C1432 B.n559 VSUBS 0.007676f
C1433 B.n560 VSUBS 0.007676f
C1434 B.n561 VSUBS 0.007676f
C1435 B.n562 VSUBS 0.007676f
C1436 B.n563 VSUBS 0.007676f
C1437 B.n564 VSUBS 0.007676f
C1438 B.n565 VSUBS 0.007676f
C1439 B.n566 VSUBS 0.007676f
C1440 B.n567 VSUBS 0.007676f
C1441 B.n568 VSUBS 0.007676f
C1442 B.n569 VSUBS 0.007676f
C1443 B.n570 VSUBS 0.007676f
C1444 B.n571 VSUBS 0.007676f
C1445 B.n572 VSUBS 0.007676f
C1446 B.n573 VSUBS 0.007676f
C1447 B.n574 VSUBS 0.007676f
C1448 B.n575 VSUBS 0.007676f
C1449 B.n576 VSUBS 0.007676f
C1450 B.n577 VSUBS 0.007676f
C1451 B.n578 VSUBS 0.007676f
C1452 B.n579 VSUBS 0.007676f
C1453 B.n580 VSUBS 0.007676f
C1454 B.n581 VSUBS 0.007676f
C1455 B.n582 VSUBS 0.007676f
C1456 B.n583 VSUBS 0.007676f
C1457 B.n584 VSUBS 0.007676f
C1458 B.n585 VSUBS 0.007676f
C1459 B.n586 VSUBS 0.007676f
C1460 B.n587 VSUBS 0.007676f
C1461 B.n588 VSUBS 0.007676f
C1462 B.n589 VSUBS 0.007676f
C1463 B.n590 VSUBS 0.007676f
C1464 B.n591 VSUBS 0.007676f
C1465 B.n592 VSUBS 0.007676f
C1466 B.n593 VSUBS 0.007676f
C1467 B.n594 VSUBS 0.007676f
C1468 B.n595 VSUBS 0.007676f
C1469 B.n596 VSUBS 0.007676f
C1470 B.n597 VSUBS 0.007676f
C1471 B.n598 VSUBS 0.007676f
C1472 B.n599 VSUBS 0.007676f
C1473 B.n600 VSUBS 0.007676f
C1474 B.n601 VSUBS 0.007676f
C1475 B.n602 VSUBS 0.007676f
C1476 B.n603 VSUBS 0.007676f
C1477 B.n604 VSUBS 0.007676f
C1478 B.n605 VSUBS 0.007676f
C1479 B.n606 VSUBS 0.007676f
C1480 B.n607 VSUBS 0.007676f
C1481 B.n608 VSUBS 0.007676f
C1482 B.n609 VSUBS 0.007676f
C1483 B.n610 VSUBS 0.007676f
C1484 B.n611 VSUBS 0.007676f
C1485 B.n612 VSUBS 0.007676f
C1486 B.n613 VSUBS 0.007676f
C1487 B.n614 VSUBS 0.007676f
C1488 B.n615 VSUBS 0.007676f
C1489 B.n616 VSUBS 0.007676f
C1490 B.n617 VSUBS 0.007676f
C1491 B.n618 VSUBS 0.007676f
C1492 B.n619 VSUBS 0.007676f
C1493 B.n620 VSUBS 0.007676f
C1494 B.n621 VSUBS 0.007676f
C1495 B.n622 VSUBS 0.007676f
C1496 B.n623 VSUBS 0.007676f
C1497 B.n624 VSUBS 0.007676f
C1498 B.n625 VSUBS 0.007676f
C1499 B.n626 VSUBS 0.007676f
C1500 B.n627 VSUBS 0.007676f
C1501 B.n628 VSUBS 0.007676f
C1502 B.n629 VSUBS 0.007676f
C1503 B.n630 VSUBS 0.007676f
C1504 B.n631 VSUBS 0.007676f
C1505 B.n632 VSUBS 0.007676f
C1506 B.n633 VSUBS 0.007676f
C1507 B.n634 VSUBS 0.007676f
C1508 B.n635 VSUBS 0.007676f
C1509 B.n636 VSUBS 0.007676f
C1510 B.n637 VSUBS 0.007676f
C1511 B.n638 VSUBS 0.007676f
C1512 B.n639 VSUBS 0.007676f
C1513 B.n640 VSUBS 0.007676f
C1514 B.n641 VSUBS 0.018293f
C1515 B.n642 VSUBS 0.019185f
C1516 B.n643 VSUBS 0.019185f
C1517 B.n644 VSUBS 0.007676f
C1518 B.n645 VSUBS 0.007676f
C1519 B.n646 VSUBS 0.007676f
C1520 B.n647 VSUBS 0.007676f
C1521 B.n648 VSUBS 0.007676f
C1522 B.n649 VSUBS 0.007676f
C1523 B.n650 VSUBS 0.007676f
C1524 B.n651 VSUBS 0.007676f
C1525 B.n652 VSUBS 0.007676f
C1526 B.n653 VSUBS 0.007676f
C1527 B.n654 VSUBS 0.007676f
C1528 B.n655 VSUBS 0.007676f
C1529 B.n656 VSUBS 0.007676f
C1530 B.n657 VSUBS 0.007676f
C1531 B.n658 VSUBS 0.007676f
C1532 B.n659 VSUBS 0.007676f
C1533 B.n660 VSUBS 0.007676f
C1534 B.n661 VSUBS 0.007676f
C1535 B.n662 VSUBS 0.007676f
C1536 B.n663 VSUBS 0.007676f
C1537 B.n664 VSUBS 0.007676f
C1538 B.n665 VSUBS 0.007676f
C1539 B.n666 VSUBS 0.007676f
C1540 B.n667 VSUBS 0.007676f
C1541 B.n668 VSUBS 0.007676f
C1542 B.n669 VSUBS 0.007676f
C1543 B.n670 VSUBS 0.007676f
C1544 B.n671 VSUBS 0.007676f
C1545 B.n672 VSUBS 0.007676f
C1546 B.n673 VSUBS 0.007676f
C1547 B.n674 VSUBS 0.007676f
C1548 B.n675 VSUBS 0.007676f
C1549 B.n676 VSUBS 0.007676f
C1550 B.n677 VSUBS 0.007676f
C1551 B.n678 VSUBS 0.007676f
C1552 B.n679 VSUBS 0.007676f
C1553 B.n680 VSUBS 0.007676f
C1554 B.n681 VSUBS 0.007676f
C1555 B.n682 VSUBS 0.007676f
C1556 B.n683 VSUBS 0.007676f
C1557 B.n684 VSUBS 0.007676f
C1558 B.n685 VSUBS 0.007676f
C1559 B.n686 VSUBS 0.007676f
C1560 B.n687 VSUBS 0.007676f
C1561 B.n688 VSUBS 0.007676f
C1562 B.n689 VSUBS 0.007676f
C1563 B.n690 VSUBS 0.007676f
C1564 B.n691 VSUBS 0.007676f
C1565 B.n692 VSUBS 0.007676f
C1566 B.n693 VSUBS 0.007676f
C1567 B.n694 VSUBS 0.007676f
C1568 B.n695 VSUBS 0.007676f
C1569 B.n696 VSUBS 0.007676f
C1570 B.n697 VSUBS 0.007676f
C1571 B.n698 VSUBS 0.007676f
C1572 B.n699 VSUBS 0.007676f
C1573 B.n700 VSUBS 0.007676f
C1574 B.n701 VSUBS 0.007676f
C1575 B.n702 VSUBS 0.007676f
C1576 B.n703 VSUBS 0.007676f
C1577 B.n704 VSUBS 0.007676f
C1578 B.n705 VSUBS 0.007676f
C1579 B.n706 VSUBS 0.007676f
C1580 B.n707 VSUBS 0.007676f
C1581 B.n708 VSUBS 0.007676f
C1582 B.n709 VSUBS 0.007676f
C1583 B.n710 VSUBS 0.007676f
C1584 B.n711 VSUBS 0.007676f
C1585 B.n712 VSUBS 0.007676f
C1586 B.n713 VSUBS 0.007676f
C1587 B.n714 VSUBS 0.007676f
C1588 B.n715 VSUBS 0.007676f
C1589 B.n716 VSUBS 0.007676f
C1590 B.n717 VSUBS 0.007676f
C1591 B.n718 VSUBS 0.007676f
C1592 B.n719 VSUBS 0.005306f
C1593 B.n720 VSUBS 0.017785f
C1594 B.n721 VSUBS 0.006209f
C1595 B.n722 VSUBS 0.007676f
C1596 B.n723 VSUBS 0.007676f
C1597 B.n724 VSUBS 0.007676f
C1598 B.n725 VSUBS 0.007676f
C1599 B.n726 VSUBS 0.007676f
C1600 B.n727 VSUBS 0.007676f
C1601 B.n728 VSUBS 0.007676f
C1602 B.n729 VSUBS 0.007676f
C1603 B.n730 VSUBS 0.007676f
C1604 B.n731 VSUBS 0.007676f
C1605 B.n732 VSUBS 0.007676f
C1606 B.n733 VSUBS 0.006209f
C1607 B.n734 VSUBS 0.007676f
C1608 B.n735 VSUBS 0.007676f
C1609 B.n736 VSUBS 0.007676f
C1610 B.n737 VSUBS 0.007676f
C1611 B.n738 VSUBS 0.007676f
C1612 B.n739 VSUBS 0.007676f
C1613 B.n740 VSUBS 0.007676f
C1614 B.n741 VSUBS 0.007676f
C1615 B.n742 VSUBS 0.007676f
C1616 B.n743 VSUBS 0.007676f
C1617 B.n744 VSUBS 0.007676f
C1618 B.n745 VSUBS 0.007676f
C1619 B.n746 VSUBS 0.007676f
C1620 B.n747 VSUBS 0.007676f
C1621 B.n748 VSUBS 0.007676f
C1622 B.n749 VSUBS 0.007676f
C1623 B.n750 VSUBS 0.007676f
C1624 B.n751 VSUBS 0.007676f
C1625 B.n752 VSUBS 0.007676f
C1626 B.n753 VSUBS 0.007676f
C1627 B.n754 VSUBS 0.007676f
C1628 B.n755 VSUBS 0.007676f
C1629 B.n756 VSUBS 0.007676f
C1630 B.n757 VSUBS 0.007676f
C1631 B.n758 VSUBS 0.007676f
C1632 B.n759 VSUBS 0.007676f
C1633 B.n760 VSUBS 0.007676f
C1634 B.n761 VSUBS 0.007676f
C1635 B.n762 VSUBS 0.007676f
C1636 B.n763 VSUBS 0.007676f
C1637 B.n764 VSUBS 0.007676f
C1638 B.n765 VSUBS 0.007676f
C1639 B.n766 VSUBS 0.007676f
C1640 B.n767 VSUBS 0.007676f
C1641 B.n768 VSUBS 0.007676f
C1642 B.n769 VSUBS 0.007676f
C1643 B.n770 VSUBS 0.007676f
C1644 B.n771 VSUBS 0.007676f
C1645 B.n772 VSUBS 0.007676f
C1646 B.n773 VSUBS 0.007676f
C1647 B.n774 VSUBS 0.007676f
C1648 B.n775 VSUBS 0.007676f
C1649 B.n776 VSUBS 0.007676f
C1650 B.n777 VSUBS 0.007676f
C1651 B.n778 VSUBS 0.007676f
C1652 B.n779 VSUBS 0.007676f
C1653 B.n780 VSUBS 0.007676f
C1654 B.n781 VSUBS 0.007676f
C1655 B.n782 VSUBS 0.007676f
C1656 B.n783 VSUBS 0.007676f
C1657 B.n784 VSUBS 0.007676f
C1658 B.n785 VSUBS 0.007676f
C1659 B.n786 VSUBS 0.007676f
C1660 B.n787 VSUBS 0.007676f
C1661 B.n788 VSUBS 0.007676f
C1662 B.n789 VSUBS 0.007676f
C1663 B.n790 VSUBS 0.007676f
C1664 B.n791 VSUBS 0.007676f
C1665 B.n792 VSUBS 0.007676f
C1666 B.n793 VSUBS 0.007676f
C1667 B.n794 VSUBS 0.007676f
C1668 B.n795 VSUBS 0.007676f
C1669 B.n796 VSUBS 0.007676f
C1670 B.n797 VSUBS 0.007676f
C1671 B.n798 VSUBS 0.007676f
C1672 B.n799 VSUBS 0.007676f
C1673 B.n800 VSUBS 0.007676f
C1674 B.n801 VSUBS 0.007676f
C1675 B.n802 VSUBS 0.007676f
C1676 B.n803 VSUBS 0.007676f
C1677 B.n804 VSUBS 0.007676f
C1678 B.n805 VSUBS 0.007676f
C1679 B.n806 VSUBS 0.007676f
C1680 B.n807 VSUBS 0.007676f
C1681 B.n808 VSUBS 0.007676f
C1682 B.n809 VSUBS 0.007676f
C1683 B.n810 VSUBS 0.007676f
C1684 B.n811 VSUBS 0.019185f
C1685 B.n812 VSUBS 0.019185f
C1686 B.n813 VSUBS 0.018293f
C1687 B.n814 VSUBS 0.007676f
C1688 B.n815 VSUBS 0.007676f
C1689 B.n816 VSUBS 0.007676f
C1690 B.n817 VSUBS 0.007676f
C1691 B.n818 VSUBS 0.007676f
C1692 B.n819 VSUBS 0.007676f
C1693 B.n820 VSUBS 0.007676f
C1694 B.n821 VSUBS 0.007676f
C1695 B.n822 VSUBS 0.007676f
C1696 B.n823 VSUBS 0.007676f
C1697 B.n824 VSUBS 0.007676f
C1698 B.n825 VSUBS 0.007676f
C1699 B.n826 VSUBS 0.007676f
C1700 B.n827 VSUBS 0.007676f
C1701 B.n828 VSUBS 0.007676f
C1702 B.n829 VSUBS 0.007676f
C1703 B.n830 VSUBS 0.007676f
C1704 B.n831 VSUBS 0.007676f
C1705 B.n832 VSUBS 0.007676f
C1706 B.n833 VSUBS 0.007676f
C1707 B.n834 VSUBS 0.007676f
C1708 B.n835 VSUBS 0.007676f
C1709 B.n836 VSUBS 0.007676f
C1710 B.n837 VSUBS 0.007676f
C1711 B.n838 VSUBS 0.007676f
C1712 B.n839 VSUBS 0.007676f
C1713 B.n840 VSUBS 0.007676f
C1714 B.n841 VSUBS 0.007676f
C1715 B.n842 VSUBS 0.007676f
C1716 B.n843 VSUBS 0.007676f
C1717 B.n844 VSUBS 0.007676f
C1718 B.n845 VSUBS 0.007676f
C1719 B.n846 VSUBS 0.007676f
C1720 B.n847 VSUBS 0.007676f
C1721 B.n848 VSUBS 0.007676f
C1722 B.n849 VSUBS 0.007676f
C1723 B.n850 VSUBS 0.007676f
C1724 B.n851 VSUBS 0.007676f
C1725 B.n852 VSUBS 0.007676f
C1726 B.n853 VSUBS 0.007676f
C1727 B.n854 VSUBS 0.007676f
C1728 B.n855 VSUBS 0.007676f
C1729 B.n856 VSUBS 0.007676f
C1730 B.n857 VSUBS 0.007676f
C1731 B.n858 VSUBS 0.007676f
C1732 B.n859 VSUBS 0.007676f
C1733 B.n860 VSUBS 0.007676f
C1734 B.n861 VSUBS 0.007676f
C1735 B.n862 VSUBS 0.007676f
C1736 B.n863 VSUBS 0.007676f
C1737 B.n864 VSUBS 0.007676f
C1738 B.n865 VSUBS 0.007676f
C1739 B.n866 VSUBS 0.007676f
C1740 B.n867 VSUBS 0.007676f
C1741 B.n868 VSUBS 0.007676f
C1742 B.n869 VSUBS 0.007676f
C1743 B.n870 VSUBS 0.007676f
C1744 B.n871 VSUBS 0.007676f
C1745 B.n872 VSUBS 0.007676f
C1746 B.n873 VSUBS 0.007676f
C1747 B.n874 VSUBS 0.007676f
C1748 B.n875 VSUBS 0.007676f
C1749 B.n876 VSUBS 0.007676f
C1750 B.n877 VSUBS 0.007676f
C1751 B.n878 VSUBS 0.007676f
C1752 B.n879 VSUBS 0.007676f
C1753 B.n880 VSUBS 0.007676f
C1754 B.n881 VSUBS 0.007676f
C1755 B.n882 VSUBS 0.007676f
C1756 B.n883 VSUBS 0.007676f
C1757 B.n884 VSUBS 0.007676f
C1758 B.n885 VSUBS 0.007676f
C1759 B.n886 VSUBS 0.007676f
C1760 B.n887 VSUBS 0.007676f
C1761 B.n888 VSUBS 0.007676f
C1762 B.n889 VSUBS 0.007676f
C1763 B.n890 VSUBS 0.007676f
C1764 B.n891 VSUBS 0.010017f
C1765 B.n892 VSUBS 0.010671f
C1766 B.n893 VSUBS 0.02122f
.ends

