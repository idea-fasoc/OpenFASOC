* NGSPICE file created from diff_pair_sample_0399.ext - technology: sky130A

.subckt diff_pair_sample_0399 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X1 VTAIL.t18 VP.t1 VDD1.t8 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X2 VDD2.t9 VN.t0 VTAIL.t7 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=2.53935 ps=15.72 w=15.39 l=1.63
X3 VTAIL.t15 VP.t2 VDD1.t7 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X4 B.t11 B.t9 B.t10 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=0 ps=0 w=15.39 l=1.63
X5 VDD1.t6 VP.t3 VTAIL.t19 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=2.53935 ps=15.72 w=15.39 l=1.63
X6 B.t8 B.t6 B.t7 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=0 ps=0 w=15.39 l=1.63
X7 VDD2.t8 VN.t1 VTAIL.t5 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=2.53935 ps=15.72 w=15.39 l=1.63
X8 VDD2.t7 VN.t2 VTAIL.t8 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X9 B.t5 B.t3 B.t4 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=0 ps=0 w=15.39 l=1.63
X10 VDD1.t5 VP.t4 VTAIL.t14 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=6.0021 ps=31.56 w=15.39 l=1.63
X11 VTAIL.t16 VP.t5 VDD1.t4 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X12 VDD2.t6 VN.t3 VTAIL.t9 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=6.0021 ps=31.56 w=15.39 l=1.63
X13 VDD1.t3 VP.t6 VTAIL.t13 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=6.0021 ps=31.56 w=15.39 l=1.63
X14 VDD2.t5 VN.t4 VTAIL.t4 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X15 VTAIL.t2 VN.t5 VDD2.t4 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X16 VDD1.t2 VP.t7 VTAIL.t12 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X17 VTAIL.t3 VN.t6 VDD2.t3 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X18 VTAIL.t17 VP.t8 VDD1.t1 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X19 VTAIL.t0 VN.t7 VDD2.t2 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X20 B.t2 B.t0 B.t1 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=0 ps=0 w=15.39 l=1.63
X21 VTAIL.t1 VN.t8 VDD2.t1 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=2.53935 ps=15.72 w=15.39 l=1.63
X22 VDD1.t0 VP.t9 VTAIL.t10 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=6.0021 pd=31.56 as=2.53935 ps=15.72 w=15.39 l=1.63
X23 VDD2.t0 VN.t9 VTAIL.t6 w_n3322_n4046# sky130_fd_pr__pfet_01v8 ad=2.53935 pd=15.72 as=6.0021 ps=31.56 w=15.39 l=1.63
R0 VP.n14 VP.t9 260.39
R1 VP.n39 VP.t3 227.546
R2 VP.n46 VP.t2 227.546
R3 VP.n53 VP.t0 227.546
R4 VP.n60 VP.t8 227.546
R5 VP.n67 VP.t6 227.546
R6 VP.n36 VP.t4 227.546
R7 VP.n29 VP.t1 227.546
R8 VP.n22 VP.t7 227.546
R9 VP.n15 VP.t5 227.546
R10 VP.n39 VP.n38 177.448
R11 VP.n68 VP.n67 177.448
R12 VP.n37 VP.n36 177.448
R13 VP.n17 VP.n16 161.3
R14 VP.n18 VP.n13 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n12 161.3
R17 VP.n24 VP.n23 161.3
R18 VP.n25 VP.n11 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n28 VP.n10 161.3
R21 VP.n31 VP.n30 161.3
R22 VP.n32 VP.n9 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n35 VP.n8 161.3
R25 VP.n66 VP.n0 161.3
R26 VP.n65 VP.n64 161.3
R27 VP.n63 VP.n1 161.3
R28 VP.n62 VP.n61 161.3
R29 VP.n59 VP.n2 161.3
R30 VP.n58 VP.n57 161.3
R31 VP.n56 VP.n3 161.3
R32 VP.n55 VP.n54 161.3
R33 VP.n52 VP.n4 161.3
R34 VP.n51 VP.n50 161.3
R35 VP.n49 VP.n5 161.3
R36 VP.n48 VP.n47 161.3
R37 VP.n45 VP.n6 161.3
R38 VP.n44 VP.n43 161.3
R39 VP.n42 VP.n7 161.3
R40 VP.n41 VP.n40 161.3
R41 VP.n44 VP.n7 56.5193
R42 VP.n51 VP.n5 56.5193
R43 VP.n58 VP.n3 56.5193
R44 VP.n65 VP.n1 56.5193
R45 VP.n34 VP.n9 56.5193
R46 VP.n27 VP.n11 56.5193
R47 VP.n20 VP.n13 56.5193
R48 VP.n15 VP.n14 55.9298
R49 VP.n38 VP.n37 50.3414
R50 VP.n40 VP.n7 24.4675
R51 VP.n45 VP.n44 24.4675
R52 VP.n47 VP.n5 24.4675
R53 VP.n52 VP.n51 24.4675
R54 VP.n54 VP.n3 24.4675
R55 VP.n59 VP.n58 24.4675
R56 VP.n61 VP.n1 24.4675
R57 VP.n66 VP.n65 24.4675
R58 VP.n35 VP.n34 24.4675
R59 VP.n28 VP.n27 24.4675
R60 VP.n30 VP.n9 24.4675
R61 VP.n21 VP.n20 24.4675
R62 VP.n23 VP.n11 24.4675
R63 VP.n16 VP.n13 24.4675
R64 VP.n17 VP.n14 17.9509
R65 VP.n46 VP.n45 14.1914
R66 VP.n61 VP.n60 14.1914
R67 VP.n30 VP.n29 14.1914
R68 VP.n53 VP.n52 12.234
R69 VP.n54 VP.n53 12.234
R70 VP.n22 VP.n21 12.234
R71 VP.n23 VP.n22 12.234
R72 VP.n47 VP.n46 10.2766
R73 VP.n60 VP.n59 10.2766
R74 VP.n29 VP.n28 10.2766
R75 VP.n16 VP.n15 10.2766
R76 VP.n40 VP.n39 8.31928
R77 VP.n67 VP.n66 8.31928
R78 VP.n36 VP.n35 8.31928
R79 VP.n18 VP.n17 0.189894
R80 VP.n19 VP.n18 0.189894
R81 VP.n19 VP.n12 0.189894
R82 VP.n24 VP.n12 0.189894
R83 VP.n25 VP.n24 0.189894
R84 VP.n26 VP.n25 0.189894
R85 VP.n26 VP.n10 0.189894
R86 VP.n31 VP.n10 0.189894
R87 VP.n32 VP.n31 0.189894
R88 VP.n33 VP.n32 0.189894
R89 VP.n33 VP.n8 0.189894
R90 VP.n37 VP.n8 0.189894
R91 VP.n41 VP.n38 0.189894
R92 VP.n42 VP.n41 0.189894
R93 VP.n43 VP.n42 0.189894
R94 VP.n43 VP.n6 0.189894
R95 VP.n48 VP.n6 0.189894
R96 VP.n49 VP.n48 0.189894
R97 VP.n50 VP.n49 0.189894
R98 VP.n50 VP.n4 0.189894
R99 VP.n55 VP.n4 0.189894
R100 VP.n56 VP.n55 0.189894
R101 VP.n57 VP.n56 0.189894
R102 VP.n57 VP.n2 0.189894
R103 VP.n62 VP.n2 0.189894
R104 VP.n63 VP.n62 0.189894
R105 VP.n64 VP.n63 0.189894
R106 VP.n64 VP.n0 0.189894
R107 VP.n68 VP.n0 0.189894
R108 VP VP.n68 0.0516364
R109 VTAIL.n352 VTAIL.n272 756.745
R110 VTAIL.n82 VTAIL.n2 756.745
R111 VTAIL.n266 VTAIL.n186 756.745
R112 VTAIL.n176 VTAIL.n96 756.745
R113 VTAIL.n301 VTAIL.n300 585
R114 VTAIL.n303 VTAIL.n302 585
R115 VTAIL.n296 VTAIL.n295 585
R116 VTAIL.n309 VTAIL.n308 585
R117 VTAIL.n311 VTAIL.n310 585
R118 VTAIL.n292 VTAIL.n291 585
R119 VTAIL.n317 VTAIL.n316 585
R120 VTAIL.n319 VTAIL.n318 585
R121 VTAIL.n288 VTAIL.n287 585
R122 VTAIL.n325 VTAIL.n324 585
R123 VTAIL.n327 VTAIL.n326 585
R124 VTAIL.n284 VTAIL.n283 585
R125 VTAIL.n333 VTAIL.n332 585
R126 VTAIL.n335 VTAIL.n334 585
R127 VTAIL.n280 VTAIL.n279 585
R128 VTAIL.n342 VTAIL.n341 585
R129 VTAIL.n343 VTAIL.n278 585
R130 VTAIL.n345 VTAIL.n344 585
R131 VTAIL.n276 VTAIL.n275 585
R132 VTAIL.n351 VTAIL.n350 585
R133 VTAIL.n353 VTAIL.n352 585
R134 VTAIL.n31 VTAIL.n30 585
R135 VTAIL.n33 VTAIL.n32 585
R136 VTAIL.n26 VTAIL.n25 585
R137 VTAIL.n39 VTAIL.n38 585
R138 VTAIL.n41 VTAIL.n40 585
R139 VTAIL.n22 VTAIL.n21 585
R140 VTAIL.n47 VTAIL.n46 585
R141 VTAIL.n49 VTAIL.n48 585
R142 VTAIL.n18 VTAIL.n17 585
R143 VTAIL.n55 VTAIL.n54 585
R144 VTAIL.n57 VTAIL.n56 585
R145 VTAIL.n14 VTAIL.n13 585
R146 VTAIL.n63 VTAIL.n62 585
R147 VTAIL.n65 VTAIL.n64 585
R148 VTAIL.n10 VTAIL.n9 585
R149 VTAIL.n72 VTAIL.n71 585
R150 VTAIL.n73 VTAIL.n8 585
R151 VTAIL.n75 VTAIL.n74 585
R152 VTAIL.n6 VTAIL.n5 585
R153 VTAIL.n81 VTAIL.n80 585
R154 VTAIL.n83 VTAIL.n82 585
R155 VTAIL.n267 VTAIL.n266 585
R156 VTAIL.n265 VTAIL.n264 585
R157 VTAIL.n190 VTAIL.n189 585
R158 VTAIL.n194 VTAIL.n192 585
R159 VTAIL.n259 VTAIL.n258 585
R160 VTAIL.n257 VTAIL.n256 585
R161 VTAIL.n196 VTAIL.n195 585
R162 VTAIL.n251 VTAIL.n250 585
R163 VTAIL.n249 VTAIL.n248 585
R164 VTAIL.n200 VTAIL.n199 585
R165 VTAIL.n243 VTAIL.n242 585
R166 VTAIL.n241 VTAIL.n240 585
R167 VTAIL.n204 VTAIL.n203 585
R168 VTAIL.n235 VTAIL.n234 585
R169 VTAIL.n233 VTAIL.n232 585
R170 VTAIL.n208 VTAIL.n207 585
R171 VTAIL.n227 VTAIL.n226 585
R172 VTAIL.n225 VTAIL.n224 585
R173 VTAIL.n212 VTAIL.n211 585
R174 VTAIL.n219 VTAIL.n218 585
R175 VTAIL.n217 VTAIL.n216 585
R176 VTAIL.n177 VTAIL.n176 585
R177 VTAIL.n175 VTAIL.n174 585
R178 VTAIL.n100 VTAIL.n99 585
R179 VTAIL.n104 VTAIL.n102 585
R180 VTAIL.n169 VTAIL.n168 585
R181 VTAIL.n167 VTAIL.n166 585
R182 VTAIL.n106 VTAIL.n105 585
R183 VTAIL.n161 VTAIL.n160 585
R184 VTAIL.n159 VTAIL.n158 585
R185 VTAIL.n110 VTAIL.n109 585
R186 VTAIL.n153 VTAIL.n152 585
R187 VTAIL.n151 VTAIL.n150 585
R188 VTAIL.n114 VTAIL.n113 585
R189 VTAIL.n145 VTAIL.n144 585
R190 VTAIL.n143 VTAIL.n142 585
R191 VTAIL.n118 VTAIL.n117 585
R192 VTAIL.n137 VTAIL.n136 585
R193 VTAIL.n135 VTAIL.n134 585
R194 VTAIL.n122 VTAIL.n121 585
R195 VTAIL.n129 VTAIL.n128 585
R196 VTAIL.n127 VTAIL.n126 585
R197 VTAIL.n299 VTAIL.t6 327.466
R198 VTAIL.n29 VTAIL.t13 327.466
R199 VTAIL.n215 VTAIL.t14 327.466
R200 VTAIL.n125 VTAIL.t9 327.466
R201 VTAIL.n302 VTAIL.n301 171.744
R202 VTAIL.n302 VTAIL.n295 171.744
R203 VTAIL.n309 VTAIL.n295 171.744
R204 VTAIL.n310 VTAIL.n309 171.744
R205 VTAIL.n310 VTAIL.n291 171.744
R206 VTAIL.n317 VTAIL.n291 171.744
R207 VTAIL.n318 VTAIL.n317 171.744
R208 VTAIL.n318 VTAIL.n287 171.744
R209 VTAIL.n325 VTAIL.n287 171.744
R210 VTAIL.n326 VTAIL.n325 171.744
R211 VTAIL.n326 VTAIL.n283 171.744
R212 VTAIL.n333 VTAIL.n283 171.744
R213 VTAIL.n334 VTAIL.n333 171.744
R214 VTAIL.n334 VTAIL.n279 171.744
R215 VTAIL.n342 VTAIL.n279 171.744
R216 VTAIL.n343 VTAIL.n342 171.744
R217 VTAIL.n344 VTAIL.n343 171.744
R218 VTAIL.n344 VTAIL.n275 171.744
R219 VTAIL.n351 VTAIL.n275 171.744
R220 VTAIL.n352 VTAIL.n351 171.744
R221 VTAIL.n32 VTAIL.n31 171.744
R222 VTAIL.n32 VTAIL.n25 171.744
R223 VTAIL.n39 VTAIL.n25 171.744
R224 VTAIL.n40 VTAIL.n39 171.744
R225 VTAIL.n40 VTAIL.n21 171.744
R226 VTAIL.n47 VTAIL.n21 171.744
R227 VTAIL.n48 VTAIL.n47 171.744
R228 VTAIL.n48 VTAIL.n17 171.744
R229 VTAIL.n55 VTAIL.n17 171.744
R230 VTAIL.n56 VTAIL.n55 171.744
R231 VTAIL.n56 VTAIL.n13 171.744
R232 VTAIL.n63 VTAIL.n13 171.744
R233 VTAIL.n64 VTAIL.n63 171.744
R234 VTAIL.n64 VTAIL.n9 171.744
R235 VTAIL.n72 VTAIL.n9 171.744
R236 VTAIL.n73 VTAIL.n72 171.744
R237 VTAIL.n74 VTAIL.n73 171.744
R238 VTAIL.n74 VTAIL.n5 171.744
R239 VTAIL.n81 VTAIL.n5 171.744
R240 VTAIL.n82 VTAIL.n81 171.744
R241 VTAIL.n266 VTAIL.n265 171.744
R242 VTAIL.n265 VTAIL.n189 171.744
R243 VTAIL.n194 VTAIL.n189 171.744
R244 VTAIL.n258 VTAIL.n194 171.744
R245 VTAIL.n258 VTAIL.n257 171.744
R246 VTAIL.n257 VTAIL.n195 171.744
R247 VTAIL.n250 VTAIL.n195 171.744
R248 VTAIL.n250 VTAIL.n249 171.744
R249 VTAIL.n249 VTAIL.n199 171.744
R250 VTAIL.n242 VTAIL.n199 171.744
R251 VTAIL.n242 VTAIL.n241 171.744
R252 VTAIL.n241 VTAIL.n203 171.744
R253 VTAIL.n234 VTAIL.n203 171.744
R254 VTAIL.n234 VTAIL.n233 171.744
R255 VTAIL.n233 VTAIL.n207 171.744
R256 VTAIL.n226 VTAIL.n207 171.744
R257 VTAIL.n226 VTAIL.n225 171.744
R258 VTAIL.n225 VTAIL.n211 171.744
R259 VTAIL.n218 VTAIL.n211 171.744
R260 VTAIL.n218 VTAIL.n217 171.744
R261 VTAIL.n176 VTAIL.n175 171.744
R262 VTAIL.n175 VTAIL.n99 171.744
R263 VTAIL.n104 VTAIL.n99 171.744
R264 VTAIL.n168 VTAIL.n104 171.744
R265 VTAIL.n168 VTAIL.n167 171.744
R266 VTAIL.n167 VTAIL.n105 171.744
R267 VTAIL.n160 VTAIL.n105 171.744
R268 VTAIL.n160 VTAIL.n159 171.744
R269 VTAIL.n159 VTAIL.n109 171.744
R270 VTAIL.n152 VTAIL.n109 171.744
R271 VTAIL.n152 VTAIL.n151 171.744
R272 VTAIL.n151 VTAIL.n113 171.744
R273 VTAIL.n144 VTAIL.n113 171.744
R274 VTAIL.n144 VTAIL.n143 171.744
R275 VTAIL.n143 VTAIL.n117 171.744
R276 VTAIL.n136 VTAIL.n117 171.744
R277 VTAIL.n136 VTAIL.n135 171.744
R278 VTAIL.n135 VTAIL.n121 171.744
R279 VTAIL.n128 VTAIL.n121 171.744
R280 VTAIL.n128 VTAIL.n127 171.744
R281 VTAIL.n301 VTAIL.t6 85.8723
R282 VTAIL.n31 VTAIL.t13 85.8723
R283 VTAIL.n217 VTAIL.t14 85.8723
R284 VTAIL.n127 VTAIL.t9 85.8723
R285 VTAIL.n185 VTAIL.n184 54.1612
R286 VTAIL.n183 VTAIL.n182 54.1612
R287 VTAIL.n95 VTAIL.n94 54.1612
R288 VTAIL.n93 VTAIL.n92 54.1612
R289 VTAIL.n359 VTAIL.n358 54.161
R290 VTAIL.n1 VTAIL.n0 54.161
R291 VTAIL.n89 VTAIL.n88 54.161
R292 VTAIL.n91 VTAIL.n90 54.161
R293 VTAIL.n357 VTAIL.n356 32.7672
R294 VTAIL.n87 VTAIL.n86 32.7672
R295 VTAIL.n271 VTAIL.n270 32.7672
R296 VTAIL.n181 VTAIL.n180 32.7672
R297 VTAIL.n93 VTAIL.n91 29.0134
R298 VTAIL.n357 VTAIL.n271 27.3238
R299 VTAIL.n300 VTAIL.n299 16.3895
R300 VTAIL.n30 VTAIL.n29 16.3895
R301 VTAIL.n216 VTAIL.n215 16.3895
R302 VTAIL.n126 VTAIL.n125 16.3895
R303 VTAIL.n345 VTAIL.n276 13.1884
R304 VTAIL.n75 VTAIL.n6 13.1884
R305 VTAIL.n192 VTAIL.n190 13.1884
R306 VTAIL.n102 VTAIL.n100 13.1884
R307 VTAIL.n303 VTAIL.n298 12.8005
R308 VTAIL.n346 VTAIL.n278 12.8005
R309 VTAIL.n350 VTAIL.n349 12.8005
R310 VTAIL.n33 VTAIL.n28 12.8005
R311 VTAIL.n76 VTAIL.n8 12.8005
R312 VTAIL.n80 VTAIL.n79 12.8005
R313 VTAIL.n264 VTAIL.n263 12.8005
R314 VTAIL.n260 VTAIL.n259 12.8005
R315 VTAIL.n219 VTAIL.n214 12.8005
R316 VTAIL.n174 VTAIL.n173 12.8005
R317 VTAIL.n170 VTAIL.n169 12.8005
R318 VTAIL.n129 VTAIL.n124 12.8005
R319 VTAIL.n304 VTAIL.n296 12.0247
R320 VTAIL.n341 VTAIL.n340 12.0247
R321 VTAIL.n353 VTAIL.n274 12.0247
R322 VTAIL.n34 VTAIL.n26 12.0247
R323 VTAIL.n71 VTAIL.n70 12.0247
R324 VTAIL.n83 VTAIL.n4 12.0247
R325 VTAIL.n267 VTAIL.n188 12.0247
R326 VTAIL.n256 VTAIL.n193 12.0247
R327 VTAIL.n220 VTAIL.n212 12.0247
R328 VTAIL.n177 VTAIL.n98 12.0247
R329 VTAIL.n166 VTAIL.n103 12.0247
R330 VTAIL.n130 VTAIL.n122 12.0247
R331 VTAIL.n308 VTAIL.n307 11.249
R332 VTAIL.n339 VTAIL.n280 11.249
R333 VTAIL.n354 VTAIL.n272 11.249
R334 VTAIL.n38 VTAIL.n37 11.249
R335 VTAIL.n69 VTAIL.n10 11.249
R336 VTAIL.n84 VTAIL.n2 11.249
R337 VTAIL.n268 VTAIL.n186 11.249
R338 VTAIL.n255 VTAIL.n196 11.249
R339 VTAIL.n224 VTAIL.n223 11.249
R340 VTAIL.n178 VTAIL.n96 11.249
R341 VTAIL.n165 VTAIL.n106 11.249
R342 VTAIL.n134 VTAIL.n133 11.249
R343 VTAIL.n311 VTAIL.n294 10.4732
R344 VTAIL.n336 VTAIL.n335 10.4732
R345 VTAIL.n41 VTAIL.n24 10.4732
R346 VTAIL.n66 VTAIL.n65 10.4732
R347 VTAIL.n252 VTAIL.n251 10.4732
R348 VTAIL.n227 VTAIL.n210 10.4732
R349 VTAIL.n162 VTAIL.n161 10.4732
R350 VTAIL.n137 VTAIL.n120 10.4732
R351 VTAIL.n312 VTAIL.n292 9.69747
R352 VTAIL.n332 VTAIL.n282 9.69747
R353 VTAIL.n42 VTAIL.n22 9.69747
R354 VTAIL.n62 VTAIL.n12 9.69747
R355 VTAIL.n248 VTAIL.n198 9.69747
R356 VTAIL.n228 VTAIL.n208 9.69747
R357 VTAIL.n158 VTAIL.n108 9.69747
R358 VTAIL.n138 VTAIL.n118 9.69747
R359 VTAIL.n356 VTAIL.n355 9.45567
R360 VTAIL.n86 VTAIL.n85 9.45567
R361 VTAIL.n270 VTAIL.n269 9.45567
R362 VTAIL.n180 VTAIL.n179 9.45567
R363 VTAIL.n355 VTAIL.n354 9.3005
R364 VTAIL.n274 VTAIL.n273 9.3005
R365 VTAIL.n349 VTAIL.n348 9.3005
R366 VTAIL.n321 VTAIL.n320 9.3005
R367 VTAIL.n290 VTAIL.n289 9.3005
R368 VTAIL.n315 VTAIL.n314 9.3005
R369 VTAIL.n313 VTAIL.n312 9.3005
R370 VTAIL.n294 VTAIL.n293 9.3005
R371 VTAIL.n307 VTAIL.n306 9.3005
R372 VTAIL.n305 VTAIL.n304 9.3005
R373 VTAIL.n298 VTAIL.n297 9.3005
R374 VTAIL.n323 VTAIL.n322 9.3005
R375 VTAIL.n286 VTAIL.n285 9.3005
R376 VTAIL.n329 VTAIL.n328 9.3005
R377 VTAIL.n331 VTAIL.n330 9.3005
R378 VTAIL.n282 VTAIL.n281 9.3005
R379 VTAIL.n337 VTAIL.n336 9.3005
R380 VTAIL.n339 VTAIL.n338 9.3005
R381 VTAIL.n340 VTAIL.n277 9.3005
R382 VTAIL.n347 VTAIL.n346 9.3005
R383 VTAIL.n85 VTAIL.n84 9.3005
R384 VTAIL.n4 VTAIL.n3 9.3005
R385 VTAIL.n79 VTAIL.n78 9.3005
R386 VTAIL.n51 VTAIL.n50 9.3005
R387 VTAIL.n20 VTAIL.n19 9.3005
R388 VTAIL.n45 VTAIL.n44 9.3005
R389 VTAIL.n43 VTAIL.n42 9.3005
R390 VTAIL.n24 VTAIL.n23 9.3005
R391 VTAIL.n37 VTAIL.n36 9.3005
R392 VTAIL.n35 VTAIL.n34 9.3005
R393 VTAIL.n28 VTAIL.n27 9.3005
R394 VTAIL.n53 VTAIL.n52 9.3005
R395 VTAIL.n16 VTAIL.n15 9.3005
R396 VTAIL.n59 VTAIL.n58 9.3005
R397 VTAIL.n61 VTAIL.n60 9.3005
R398 VTAIL.n12 VTAIL.n11 9.3005
R399 VTAIL.n67 VTAIL.n66 9.3005
R400 VTAIL.n69 VTAIL.n68 9.3005
R401 VTAIL.n70 VTAIL.n7 9.3005
R402 VTAIL.n77 VTAIL.n76 9.3005
R403 VTAIL.n202 VTAIL.n201 9.3005
R404 VTAIL.n245 VTAIL.n244 9.3005
R405 VTAIL.n247 VTAIL.n246 9.3005
R406 VTAIL.n198 VTAIL.n197 9.3005
R407 VTAIL.n253 VTAIL.n252 9.3005
R408 VTAIL.n255 VTAIL.n254 9.3005
R409 VTAIL.n193 VTAIL.n191 9.3005
R410 VTAIL.n261 VTAIL.n260 9.3005
R411 VTAIL.n269 VTAIL.n268 9.3005
R412 VTAIL.n188 VTAIL.n187 9.3005
R413 VTAIL.n263 VTAIL.n262 9.3005
R414 VTAIL.n239 VTAIL.n238 9.3005
R415 VTAIL.n237 VTAIL.n236 9.3005
R416 VTAIL.n206 VTAIL.n205 9.3005
R417 VTAIL.n231 VTAIL.n230 9.3005
R418 VTAIL.n229 VTAIL.n228 9.3005
R419 VTAIL.n210 VTAIL.n209 9.3005
R420 VTAIL.n223 VTAIL.n222 9.3005
R421 VTAIL.n221 VTAIL.n220 9.3005
R422 VTAIL.n214 VTAIL.n213 9.3005
R423 VTAIL.n112 VTAIL.n111 9.3005
R424 VTAIL.n155 VTAIL.n154 9.3005
R425 VTAIL.n157 VTAIL.n156 9.3005
R426 VTAIL.n108 VTAIL.n107 9.3005
R427 VTAIL.n163 VTAIL.n162 9.3005
R428 VTAIL.n165 VTAIL.n164 9.3005
R429 VTAIL.n103 VTAIL.n101 9.3005
R430 VTAIL.n171 VTAIL.n170 9.3005
R431 VTAIL.n179 VTAIL.n178 9.3005
R432 VTAIL.n98 VTAIL.n97 9.3005
R433 VTAIL.n173 VTAIL.n172 9.3005
R434 VTAIL.n149 VTAIL.n148 9.3005
R435 VTAIL.n147 VTAIL.n146 9.3005
R436 VTAIL.n116 VTAIL.n115 9.3005
R437 VTAIL.n141 VTAIL.n140 9.3005
R438 VTAIL.n139 VTAIL.n138 9.3005
R439 VTAIL.n120 VTAIL.n119 9.3005
R440 VTAIL.n133 VTAIL.n132 9.3005
R441 VTAIL.n131 VTAIL.n130 9.3005
R442 VTAIL.n124 VTAIL.n123 9.3005
R443 VTAIL.n316 VTAIL.n315 8.92171
R444 VTAIL.n331 VTAIL.n284 8.92171
R445 VTAIL.n46 VTAIL.n45 8.92171
R446 VTAIL.n61 VTAIL.n14 8.92171
R447 VTAIL.n247 VTAIL.n200 8.92171
R448 VTAIL.n232 VTAIL.n231 8.92171
R449 VTAIL.n157 VTAIL.n110 8.92171
R450 VTAIL.n142 VTAIL.n141 8.92171
R451 VTAIL.n319 VTAIL.n290 8.14595
R452 VTAIL.n328 VTAIL.n327 8.14595
R453 VTAIL.n49 VTAIL.n20 8.14595
R454 VTAIL.n58 VTAIL.n57 8.14595
R455 VTAIL.n244 VTAIL.n243 8.14595
R456 VTAIL.n235 VTAIL.n206 8.14595
R457 VTAIL.n154 VTAIL.n153 8.14595
R458 VTAIL.n145 VTAIL.n116 8.14595
R459 VTAIL.n320 VTAIL.n288 7.3702
R460 VTAIL.n324 VTAIL.n286 7.3702
R461 VTAIL.n50 VTAIL.n18 7.3702
R462 VTAIL.n54 VTAIL.n16 7.3702
R463 VTAIL.n240 VTAIL.n202 7.3702
R464 VTAIL.n236 VTAIL.n204 7.3702
R465 VTAIL.n150 VTAIL.n112 7.3702
R466 VTAIL.n146 VTAIL.n114 7.3702
R467 VTAIL.n323 VTAIL.n288 6.59444
R468 VTAIL.n324 VTAIL.n323 6.59444
R469 VTAIL.n53 VTAIL.n18 6.59444
R470 VTAIL.n54 VTAIL.n53 6.59444
R471 VTAIL.n240 VTAIL.n239 6.59444
R472 VTAIL.n239 VTAIL.n204 6.59444
R473 VTAIL.n150 VTAIL.n149 6.59444
R474 VTAIL.n149 VTAIL.n114 6.59444
R475 VTAIL.n320 VTAIL.n319 5.81868
R476 VTAIL.n327 VTAIL.n286 5.81868
R477 VTAIL.n50 VTAIL.n49 5.81868
R478 VTAIL.n57 VTAIL.n16 5.81868
R479 VTAIL.n243 VTAIL.n202 5.81868
R480 VTAIL.n236 VTAIL.n235 5.81868
R481 VTAIL.n153 VTAIL.n112 5.81868
R482 VTAIL.n146 VTAIL.n145 5.81868
R483 VTAIL.n316 VTAIL.n290 5.04292
R484 VTAIL.n328 VTAIL.n284 5.04292
R485 VTAIL.n46 VTAIL.n20 5.04292
R486 VTAIL.n58 VTAIL.n14 5.04292
R487 VTAIL.n244 VTAIL.n200 5.04292
R488 VTAIL.n232 VTAIL.n206 5.04292
R489 VTAIL.n154 VTAIL.n110 5.04292
R490 VTAIL.n142 VTAIL.n116 5.04292
R491 VTAIL.n315 VTAIL.n292 4.26717
R492 VTAIL.n332 VTAIL.n331 4.26717
R493 VTAIL.n45 VTAIL.n22 4.26717
R494 VTAIL.n62 VTAIL.n61 4.26717
R495 VTAIL.n248 VTAIL.n247 4.26717
R496 VTAIL.n231 VTAIL.n208 4.26717
R497 VTAIL.n158 VTAIL.n157 4.26717
R498 VTAIL.n141 VTAIL.n118 4.26717
R499 VTAIL.n299 VTAIL.n297 3.70982
R500 VTAIL.n29 VTAIL.n27 3.70982
R501 VTAIL.n215 VTAIL.n213 3.70982
R502 VTAIL.n125 VTAIL.n123 3.70982
R503 VTAIL.n312 VTAIL.n311 3.49141
R504 VTAIL.n335 VTAIL.n282 3.49141
R505 VTAIL.n42 VTAIL.n41 3.49141
R506 VTAIL.n65 VTAIL.n12 3.49141
R507 VTAIL.n251 VTAIL.n198 3.49141
R508 VTAIL.n228 VTAIL.n227 3.49141
R509 VTAIL.n161 VTAIL.n108 3.49141
R510 VTAIL.n138 VTAIL.n137 3.49141
R511 VTAIL.n308 VTAIL.n294 2.71565
R512 VTAIL.n336 VTAIL.n280 2.71565
R513 VTAIL.n356 VTAIL.n272 2.71565
R514 VTAIL.n38 VTAIL.n24 2.71565
R515 VTAIL.n66 VTAIL.n10 2.71565
R516 VTAIL.n86 VTAIL.n2 2.71565
R517 VTAIL.n270 VTAIL.n186 2.71565
R518 VTAIL.n252 VTAIL.n196 2.71565
R519 VTAIL.n224 VTAIL.n210 2.71565
R520 VTAIL.n180 VTAIL.n96 2.71565
R521 VTAIL.n162 VTAIL.n106 2.71565
R522 VTAIL.n134 VTAIL.n120 2.71565
R523 VTAIL.n358 VTAIL.t4 2.11259
R524 VTAIL.n358 VTAIL.t0 2.11259
R525 VTAIL.n0 VTAIL.t5 2.11259
R526 VTAIL.n0 VTAIL.t2 2.11259
R527 VTAIL.n88 VTAIL.t11 2.11259
R528 VTAIL.n88 VTAIL.t17 2.11259
R529 VTAIL.n90 VTAIL.t19 2.11259
R530 VTAIL.n90 VTAIL.t15 2.11259
R531 VTAIL.n184 VTAIL.t12 2.11259
R532 VTAIL.n184 VTAIL.t18 2.11259
R533 VTAIL.n182 VTAIL.t10 2.11259
R534 VTAIL.n182 VTAIL.t16 2.11259
R535 VTAIL.n94 VTAIL.t8 2.11259
R536 VTAIL.n94 VTAIL.t1 2.11259
R537 VTAIL.n92 VTAIL.t7 2.11259
R538 VTAIL.n92 VTAIL.t3 2.11259
R539 VTAIL.n307 VTAIL.n296 1.93989
R540 VTAIL.n341 VTAIL.n339 1.93989
R541 VTAIL.n354 VTAIL.n353 1.93989
R542 VTAIL.n37 VTAIL.n26 1.93989
R543 VTAIL.n71 VTAIL.n69 1.93989
R544 VTAIL.n84 VTAIL.n83 1.93989
R545 VTAIL.n268 VTAIL.n267 1.93989
R546 VTAIL.n256 VTAIL.n255 1.93989
R547 VTAIL.n223 VTAIL.n212 1.93989
R548 VTAIL.n178 VTAIL.n177 1.93989
R549 VTAIL.n166 VTAIL.n165 1.93989
R550 VTAIL.n133 VTAIL.n122 1.93989
R551 VTAIL.n95 VTAIL.n93 1.69016
R552 VTAIL.n181 VTAIL.n95 1.69016
R553 VTAIL.n185 VTAIL.n183 1.69016
R554 VTAIL.n271 VTAIL.n185 1.69016
R555 VTAIL.n91 VTAIL.n89 1.69016
R556 VTAIL.n89 VTAIL.n87 1.69016
R557 VTAIL.n359 VTAIL.n357 1.69016
R558 VTAIL VTAIL.n1 1.32593
R559 VTAIL.n183 VTAIL.n181 1.31516
R560 VTAIL.n87 VTAIL.n1 1.31516
R561 VTAIL.n304 VTAIL.n303 1.16414
R562 VTAIL.n340 VTAIL.n278 1.16414
R563 VTAIL.n350 VTAIL.n274 1.16414
R564 VTAIL.n34 VTAIL.n33 1.16414
R565 VTAIL.n70 VTAIL.n8 1.16414
R566 VTAIL.n80 VTAIL.n4 1.16414
R567 VTAIL.n264 VTAIL.n188 1.16414
R568 VTAIL.n259 VTAIL.n193 1.16414
R569 VTAIL.n220 VTAIL.n219 1.16414
R570 VTAIL.n174 VTAIL.n98 1.16414
R571 VTAIL.n169 VTAIL.n103 1.16414
R572 VTAIL.n130 VTAIL.n129 1.16414
R573 VTAIL.n300 VTAIL.n298 0.388379
R574 VTAIL.n346 VTAIL.n345 0.388379
R575 VTAIL.n349 VTAIL.n276 0.388379
R576 VTAIL.n30 VTAIL.n28 0.388379
R577 VTAIL.n76 VTAIL.n75 0.388379
R578 VTAIL.n79 VTAIL.n6 0.388379
R579 VTAIL.n263 VTAIL.n190 0.388379
R580 VTAIL.n260 VTAIL.n192 0.388379
R581 VTAIL.n216 VTAIL.n214 0.388379
R582 VTAIL.n173 VTAIL.n100 0.388379
R583 VTAIL.n170 VTAIL.n102 0.388379
R584 VTAIL.n126 VTAIL.n124 0.388379
R585 VTAIL VTAIL.n359 0.364724
R586 VTAIL.n305 VTAIL.n297 0.155672
R587 VTAIL.n306 VTAIL.n305 0.155672
R588 VTAIL.n306 VTAIL.n293 0.155672
R589 VTAIL.n313 VTAIL.n293 0.155672
R590 VTAIL.n314 VTAIL.n313 0.155672
R591 VTAIL.n314 VTAIL.n289 0.155672
R592 VTAIL.n321 VTAIL.n289 0.155672
R593 VTAIL.n322 VTAIL.n321 0.155672
R594 VTAIL.n322 VTAIL.n285 0.155672
R595 VTAIL.n329 VTAIL.n285 0.155672
R596 VTAIL.n330 VTAIL.n329 0.155672
R597 VTAIL.n330 VTAIL.n281 0.155672
R598 VTAIL.n337 VTAIL.n281 0.155672
R599 VTAIL.n338 VTAIL.n337 0.155672
R600 VTAIL.n338 VTAIL.n277 0.155672
R601 VTAIL.n347 VTAIL.n277 0.155672
R602 VTAIL.n348 VTAIL.n347 0.155672
R603 VTAIL.n348 VTAIL.n273 0.155672
R604 VTAIL.n355 VTAIL.n273 0.155672
R605 VTAIL.n35 VTAIL.n27 0.155672
R606 VTAIL.n36 VTAIL.n35 0.155672
R607 VTAIL.n36 VTAIL.n23 0.155672
R608 VTAIL.n43 VTAIL.n23 0.155672
R609 VTAIL.n44 VTAIL.n43 0.155672
R610 VTAIL.n44 VTAIL.n19 0.155672
R611 VTAIL.n51 VTAIL.n19 0.155672
R612 VTAIL.n52 VTAIL.n51 0.155672
R613 VTAIL.n52 VTAIL.n15 0.155672
R614 VTAIL.n59 VTAIL.n15 0.155672
R615 VTAIL.n60 VTAIL.n59 0.155672
R616 VTAIL.n60 VTAIL.n11 0.155672
R617 VTAIL.n67 VTAIL.n11 0.155672
R618 VTAIL.n68 VTAIL.n67 0.155672
R619 VTAIL.n68 VTAIL.n7 0.155672
R620 VTAIL.n77 VTAIL.n7 0.155672
R621 VTAIL.n78 VTAIL.n77 0.155672
R622 VTAIL.n78 VTAIL.n3 0.155672
R623 VTAIL.n85 VTAIL.n3 0.155672
R624 VTAIL.n269 VTAIL.n187 0.155672
R625 VTAIL.n262 VTAIL.n187 0.155672
R626 VTAIL.n262 VTAIL.n261 0.155672
R627 VTAIL.n261 VTAIL.n191 0.155672
R628 VTAIL.n254 VTAIL.n191 0.155672
R629 VTAIL.n254 VTAIL.n253 0.155672
R630 VTAIL.n253 VTAIL.n197 0.155672
R631 VTAIL.n246 VTAIL.n197 0.155672
R632 VTAIL.n246 VTAIL.n245 0.155672
R633 VTAIL.n245 VTAIL.n201 0.155672
R634 VTAIL.n238 VTAIL.n201 0.155672
R635 VTAIL.n238 VTAIL.n237 0.155672
R636 VTAIL.n237 VTAIL.n205 0.155672
R637 VTAIL.n230 VTAIL.n205 0.155672
R638 VTAIL.n230 VTAIL.n229 0.155672
R639 VTAIL.n229 VTAIL.n209 0.155672
R640 VTAIL.n222 VTAIL.n209 0.155672
R641 VTAIL.n222 VTAIL.n221 0.155672
R642 VTAIL.n221 VTAIL.n213 0.155672
R643 VTAIL.n179 VTAIL.n97 0.155672
R644 VTAIL.n172 VTAIL.n97 0.155672
R645 VTAIL.n172 VTAIL.n171 0.155672
R646 VTAIL.n171 VTAIL.n101 0.155672
R647 VTAIL.n164 VTAIL.n101 0.155672
R648 VTAIL.n164 VTAIL.n163 0.155672
R649 VTAIL.n163 VTAIL.n107 0.155672
R650 VTAIL.n156 VTAIL.n107 0.155672
R651 VTAIL.n156 VTAIL.n155 0.155672
R652 VTAIL.n155 VTAIL.n111 0.155672
R653 VTAIL.n148 VTAIL.n111 0.155672
R654 VTAIL.n148 VTAIL.n147 0.155672
R655 VTAIL.n147 VTAIL.n115 0.155672
R656 VTAIL.n140 VTAIL.n115 0.155672
R657 VTAIL.n140 VTAIL.n139 0.155672
R658 VTAIL.n139 VTAIL.n119 0.155672
R659 VTAIL.n132 VTAIL.n119 0.155672
R660 VTAIL.n132 VTAIL.n131 0.155672
R661 VTAIL.n131 VTAIL.n123 0.155672
R662 VDD1.n80 VDD1.n0 756.745
R663 VDD1.n167 VDD1.n87 756.745
R664 VDD1.n81 VDD1.n80 585
R665 VDD1.n79 VDD1.n78 585
R666 VDD1.n4 VDD1.n3 585
R667 VDD1.n8 VDD1.n6 585
R668 VDD1.n73 VDD1.n72 585
R669 VDD1.n71 VDD1.n70 585
R670 VDD1.n10 VDD1.n9 585
R671 VDD1.n65 VDD1.n64 585
R672 VDD1.n63 VDD1.n62 585
R673 VDD1.n14 VDD1.n13 585
R674 VDD1.n57 VDD1.n56 585
R675 VDD1.n55 VDD1.n54 585
R676 VDD1.n18 VDD1.n17 585
R677 VDD1.n49 VDD1.n48 585
R678 VDD1.n47 VDD1.n46 585
R679 VDD1.n22 VDD1.n21 585
R680 VDD1.n41 VDD1.n40 585
R681 VDD1.n39 VDD1.n38 585
R682 VDD1.n26 VDD1.n25 585
R683 VDD1.n33 VDD1.n32 585
R684 VDD1.n31 VDD1.n30 585
R685 VDD1.n116 VDD1.n115 585
R686 VDD1.n118 VDD1.n117 585
R687 VDD1.n111 VDD1.n110 585
R688 VDD1.n124 VDD1.n123 585
R689 VDD1.n126 VDD1.n125 585
R690 VDD1.n107 VDD1.n106 585
R691 VDD1.n132 VDD1.n131 585
R692 VDD1.n134 VDD1.n133 585
R693 VDD1.n103 VDD1.n102 585
R694 VDD1.n140 VDD1.n139 585
R695 VDD1.n142 VDD1.n141 585
R696 VDD1.n99 VDD1.n98 585
R697 VDD1.n148 VDD1.n147 585
R698 VDD1.n150 VDD1.n149 585
R699 VDD1.n95 VDD1.n94 585
R700 VDD1.n157 VDD1.n156 585
R701 VDD1.n158 VDD1.n93 585
R702 VDD1.n160 VDD1.n159 585
R703 VDD1.n91 VDD1.n90 585
R704 VDD1.n166 VDD1.n165 585
R705 VDD1.n168 VDD1.n167 585
R706 VDD1.n29 VDD1.t0 327.466
R707 VDD1.n114 VDD1.t6 327.466
R708 VDD1.n80 VDD1.n79 171.744
R709 VDD1.n79 VDD1.n3 171.744
R710 VDD1.n8 VDD1.n3 171.744
R711 VDD1.n72 VDD1.n8 171.744
R712 VDD1.n72 VDD1.n71 171.744
R713 VDD1.n71 VDD1.n9 171.744
R714 VDD1.n64 VDD1.n9 171.744
R715 VDD1.n64 VDD1.n63 171.744
R716 VDD1.n63 VDD1.n13 171.744
R717 VDD1.n56 VDD1.n13 171.744
R718 VDD1.n56 VDD1.n55 171.744
R719 VDD1.n55 VDD1.n17 171.744
R720 VDD1.n48 VDD1.n17 171.744
R721 VDD1.n48 VDD1.n47 171.744
R722 VDD1.n47 VDD1.n21 171.744
R723 VDD1.n40 VDD1.n21 171.744
R724 VDD1.n40 VDD1.n39 171.744
R725 VDD1.n39 VDD1.n25 171.744
R726 VDD1.n32 VDD1.n25 171.744
R727 VDD1.n32 VDD1.n31 171.744
R728 VDD1.n117 VDD1.n116 171.744
R729 VDD1.n117 VDD1.n110 171.744
R730 VDD1.n124 VDD1.n110 171.744
R731 VDD1.n125 VDD1.n124 171.744
R732 VDD1.n125 VDD1.n106 171.744
R733 VDD1.n132 VDD1.n106 171.744
R734 VDD1.n133 VDD1.n132 171.744
R735 VDD1.n133 VDD1.n102 171.744
R736 VDD1.n140 VDD1.n102 171.744
R737 VDD1.n141 VDD1.n140 171.744
R738 VDD1.n141 VDD1.n98 171.744
R739 VDD1.n148 VDD1.n98 171.744
R740 VDD1.n149 VDD1.n148 171.744
R741 VDD1.n149 VDD1.n94 171.744
R742 VDD1.n157 VDD1.n94 171.744
R743 VDD1.n158 VDD1.n157 171.744
R744 VDD1.n159 VDD1.n158 171.744
R745 VDD1.n159 VDD1.n90 171.744
R746 VDD1.n166 VDD1.n90 171.744
R747 VDD1.n167 VDD1.n166 171.744
R748 VDD1.n31 VDD1.t0 85.8723
R749 VDD1.n116 VDD1.t6 85.8723
R750 VDD1.n175 VDD1.n174 72.0517
R751 VDD1.n86 VDD1.n85 70.84
R752 VDD1.n173 VDD1.n172 70.8398
R753 VDD1.n177 VDD1.n176 70.8398
R754 VDD1.n86 VDD1.n84 51.1356
R755 VDD1.n173 VDD1.n171 51.1356
R756 VDD1.n177 VDD1.n175 46.4362
R757 VDD1.n30 VDD1.n29 16.3895
R758 VDD1.n115 VDD1.n114 16.3895
R759 VDD1.n6 VDD1.n4 13.1884
R760 VDD1.n160 VDD1.n91 13.1884
R761 VDD1.n78 VDD1.n77 12.8005
R762 VDD1.n74 VDD1.n73 12.8005
R763 VDD1.n33 VDD1.n28 12.8005
R764 VDD1.n118 VDD1.n113 12.8005
R765 VDD1.n161 VDD1.n93 12.8005
R766 VDD1.n165 VDD1.n164 12.8005
R767 VDD1.n81 VDD1.n2 12.0247
R768 VDD1.n70 VDD1.n7 12.0247
R769 VDD1.n34 VDD1.n26 12.0247
R770 VDD1.n119 VDD1.n111 12.0247
R771 VDD1.n156 VDD1.n155 12.0247
R772 VDD1.n168 VDD1.n89 12.0247
R773 VDD1.n82 VDD1.n0 11.249
R774 VDD1.n69 VDD1.n10 11.249
R775 VDD1.n38 VDD1.n37 11.249
R776 VDD1.n123 VDD1.n122 11.249
R777 VDD1.n154 VDD1.n95 11.249
R778 VDD1.n169 VDD1.n87 11.249
R779 VDD1.n66 VDD1.n65 10.4732
R780 VDD1.n41 VDD1.n24 10.4732
R781 VDD1.n126 VDD1.n109 10.4732
R782 VDD1.n151 VDD1.n150 10.4732
R783 VDD1.n62 VDD1.n12 9.69747
R784 VDD1.n42 VDD1.n22 9.69747
R785 VDD1.n127 VDD1.n107 9.69747
R786 VDD1.n147 VDD1.n97 9.69747
R787 VDD1.n84 VDD1.n83 9.45567
R788 VDD1.n171 VDD1.n170 9.45567
R789 VDD1.n16 VDD1.n15 9.3005
R790 VDD1.n59 VDD1.n58 9.3005
R791 VDD1.n61 VDD1.n60 9.3005
R792 VDD1.n12 VDD1.n11 9.3005
R793 VDD1.n67 VDD1.n66 9.3005
R794 VDD1.n69 VDD1.n68 9.3005
R795 VDD1.n7 VDD1.n5 9.3005
R796 VDD1.n75 VDD1.n74 9.3005
R797 VDD1.n83 VDD1.n82 9.3005
R798 VDD1.n2 VDD1.n1 9.3005
R799 VDD1.n77 VDD1.n76 9.3005
R800 VDD1.n53 VDD1.n52 9.3005
R801 VDD1.n51 VDD1.n50 9.3005
R802 VDD1.n20 VDD1.n19 9.3005
R803 VDD1.n45 VDD1.n44 9.3005
R804 VDD1.n43 VDD1.n42 9.3005
R805 VDD1.n24 VDD1.n23 9.3005
R806 VDD1.n37 VDD1.n36 9.3005
R807 VDD1.n35 VDD1.n34 9.3005
R808 VDD1.n28 VDD1.n27 9.3005
R809 VDD1.n170 VDD1.n169 9.3005
R810 VDD1.n89 VDD1.n88 9.3005
R811 VDD1.n164 VDD1.n163 9.3005
R812 VDD1.n136 VDD1.n135 9.3005
R813 VDD1.n105 VDD1.n104 9.3005
R814 VDD1.n130 VDD1.n129 9.3005
R815 VDD1.n128 VDD1.n127 9.3005
R816 VDD1.n109 VDD1.n108 9.3005
R817 VDD1.n122 VDD1.n121 9.3005
R818 VDD1.n120 VDD1.n119 9.3005
R819 VDD1.n113 VDD1.n112 9.3005
R820 VDD1.n138 VDD1.n137 9.3005
R821 VDD1.n101 VDD1.n100 9.3005
R822 VDD1.n144 VDD1.n143 9.3005
R823 VDD1.n146 VDD1.n145 9.3005
R824 VDD1.n97 VDD1.n96 9.3005
R825 VDD1.n152 VDD1.n151 9.3005
R826 VDD1.n154 VDD1.n153 9.3005
R827 VDD1.n155 VDD1.n92 9.3005
R828 VDD1.n162 VDD1.n161 9.3005
R829 VDD1.n61 VDD1.n14 8.92171
R830 VDD1.n46 VDD1.n45 8.92171
R831 VDD1.n131 VDD1.n130 8.92171
R832 VDD1.n146 VDD1.n99 8.92171
R833 VDD1.n58 VDD1.n57 8.14595
R834 VDD1.n49 VDD1.n20 8.14595
R835 VDD1.n134 VDD1.n105 8.14595
R836 VDD1.n143 VDD1.n142 8.14595
R837 VDD1.n54 VDD1.n16 7.3702
R838 VDD1.n50 VDD1.n18 7.3702
R839 VDD1.n135 VDD1.n103 7.3702
R840 VDD1.n139 VDD1.n101 7.3702
R841 VDD1.n54 VDD1.n53 6.59444
R842 VDD1.n53 VDD1.n18 6.59444
R843 VDD1.n138 VDD1.n103 6.59444
R844 VDD1.n139 VDD1.n138 6.59444
R845 VDD1.n57 VDD1.n16 5.81868
R846 VDD1.n50 VDD1.n49 5.81868
R847 VDD1.n135 VDD1.n134 5.81868
R848 VDD1.n142 VDD1.n101 5.81868
R849 VDD1.n58 VDD1.n14 5.04292
R850 VDD1.n46 VDD1.n20 5.04292
R851 VDD1.n131 VDD1.n105 5.04292
R852 VDD1.n143 VDD1.n99 5.04292
R853 VDD1.n62 VDD1.n61 4.26717
R854 VDD1.n45 VDD1.n22 4.26717
R855 VDD1.n130 VDD1.n107 4.26717
R856 VDD1.n147 VDD1.n146 4.26717
R857 VDD1.n29 VDD1.n27 3.70982
R858 VDD1.n114 VDD1.n112 3.70982
R859 VDD1.n65 VDD1.n12 3.49141
R860 VDD1.n42 VDD1.n41 3.49141
R861 VDD1.n127 VDD1.n126 3.49141
R862 VDD1.n150 VDD1.n97 3.49141
R863 VDD1.n84 VDD1.n0 2.71565
R864 VDD1.n66 VDD1.n10 2.71565
R865 VDD1.n38 VDD1.n24 2.71565
R866 VDD1.n123 VDD1.n109 2.71565
R867 VDD1.n151 VDD1.n95 2.71565
R868 VDD1.n171 VDD1.n87 2.71565
R869 VDD1.n176 VDD1.t8 2.11259
R870 VDD1.n176 VDD1.t5 2.11259
R871 VDD1.n85 VDD1.t4 2.11259
R872 VDD1.n85 VDD1.t2 2.11259
R873 VDD1.n174 VDD1.t1 2.11259
R874 VDD1.n174 VDD1.t3 2.11259
R875 VDD1.n172 VDD1.t7 2.11259
R876 VDD1.n172 VDD1.t9 2.11259
R877 VDD1.n82 VDD1.n81 1.93989
R878 VDD1.n70 VDD1.n69 1.93989
R879 VDD1.n37 VDD1.n26 1.93989
R880 VDD1.n122 VDD1.n111 1.93989
R881 VDD1.n156 VDD1.n154 1.93989
R882 VDD1.n169 VDD1.n168 1.93989
R883 VDD1 VDD1.n177 1.20955
R884 VDD1.n78 VDD1.n2 1.16414
R885 VDD1.n73 VDD1.n7 1.16414
R886 VDD1.n34 VDD1.n33 1.16414
R887 VDD1.n119 VDD1.n118 1.16414
R888 VDD1.n155 VDD1.n93 1.16414
R889 VDD1.n165 VDD1.n89 1.16414
R890 VDD1 VDD1.n86 0.481103
R891 VDD1.n77 VDD1.n4 0.388379
R892 VDD1.n74 VDD1.n6 0.388379
R893 VDD1.n30 VDD1.n28 0.388379
R894 VDD1.n115 VDD1.n113 0.388379
R895 VDD1.n161 VDD1.n160 0.388379
R896 VDD1.n164 VDD1.n91 0.388379
R897 VDD1.n175 VDD1.n173 0.367568
R898 VDD1.n83 VDD1.n1 0.155672
R899 VDD1.n76 VDD1.n1 0.155672
R900 VDD1.n76 VDD1.n75 0.155672
R901 VDD1.n75 VDD1.n5 0.155672
R902 VDD1.n68 VDD1.n5 0.155672
R903 VDD1.n68 VDD1.n67 0.155672
R904 VDD1.n67 VDD1.n11 0.155672
R905 VDD1.n60 VDD1.n11 0.155672
R906 VDD1.n60 VDD1.n59 0.155672
R907 VDD1.n59 VDD1.n15 0.155672
R908 VDD1.n52 VDD1.n15 0.155672
R909 VDD1.n52 VDD1.n51 0.155672
R910 VDD1.n51 VDD1.n19 0.155672
R911 VDD1.n44 VDD1.n19 0.155672
R912 VDD1.n44 VDD1.n43 0.155672
R913 VDD1.n43 VDD1.n23 0.155672
R914 VDD1.n36 VDD1.n23 0.155672
R915 VDD1.n36 VDD1.n35 0.155672
R916 VDD1.n35 VDD1.n27 0.155672
R917 VDD1.n120 VDD1.n112 0.155672
R918 VDD1.n121 VDD1.n120 0.155672
R919 VDD1.n121 VDD1.n108 0.155672
R920 VDD1.n128 VDD1.n108 0.155672
R921 VDD1.n129 VDD1.n128 0.155672
R922 VDD1.n129 VDD1.n104 0.155672
R923 VDD1.n136 VDD1.n104 0.155672
R924 VDD1.n137 VDD1.n136 0.155672
R925 VDD1.n137 VDD1.n100 0.155672
R926 VDD1.n144 VDD1.n100 0.155672
R927 VDD1.n145 VDD1.n144 0.155672
R928 VDD1.n145 VDD1.n96 0.155672
R929 VDD1.n152 VDD1.n96 0.155672
R930 VDD1.n153 VDD1.n152 0.155672
R931 VDD1.n153 VDD1.n92 0.155672
R932 VDD1.n162 VDD1.n92 0.155672
R933 VDD1.n163 VDD1.n162 0.155672
R934 VDD1.n163 VDD1.n88 0.155672
R935 VDD1.n170 VDD1.n88 0.155672
R936 VN.n6 VN.t1 260.39
R937 VN.n36 VN.t3 260.39
R938 VN.n7 VN.t5 227.546
R939 VN.n14 VN.t4 227.546
R940 VN.n21 VN.t7 227.546
R941 VN.n28 VN.t9 227.546
R942 VN.n37 VN.t8 227.546
R943 VN.n44 VN.t2 227.546
R944 VN.n51 VN.t6 227.546
R945 VN.n58 VN.t0 227.546
R946 VN.n29 VN.n28 177.448
R947 VN.n59 VN.n58 177.448
R948 VN.n57 VN.n30 161.3
R949 VN.n56 VN.n55 161.3
R950 VN.n54 VN.n31 161.3
R951 VN.n53 VN.n52 161.3
R952 VN.n50 VN.n32 161.3
R953 VN.n49 VN.n48 161.3
R954 VN.n47 VN.n33 161.3
R955 VN.n46 VN.n45 161.3
R956 VN.n43 VN.n34 161.3
R957 VN.n42 VN.n41 161.3
R958 VN.n40 VN.n35 161.3
R959 VN.n39 VN.n38 161.3
R960 VN.n27 VN.n0 161.3
R961 VN.n26 VN.n25 161.3
R962 VN.n24 VN.n1 161.3
R963 VN.n23 VN.n22 161.3
R964 VN.n20 VN.n2 161.3
R965 VN.n19 VN.n18 161.3
R966 VN.n17 VN.n3 161.3
R967 VN.n16 VN.n15 161.3
R968 VN.n13 VN.n4 161.3
R969 VN.n12 VN.n11 161.3
R970 VN.n10 VN.n5 161.3
R971 VN.n9 VN.n8 161.3
R972 VN.n12 VN.n5 56.5193
R973 VN.n19 VN.n3 56.5193
R974 VN.n26 VN.n1 56.5193
R975 VN.n42 VN.n35 56.5193
R976 VN.n49 VN.n33 56.5193
R977 VN.n56 VN.n31 56.5193
R978 VN.n7 VN.n6 55.9298
R979 VN.n37 VN.n36 55.9298
R980 VN VN.n59 50.7221
R981 VN.n8 VN.n5 24.4675
R982 VN.n13 VN.n12 24.4675
R983 VN.n15 VN.n3 24.4675
R984 VN.n20 VN.n19 24.4675
R985 VN.n22 VN.n1 24.4675
R986 VN.n27 VN.n26 24.4675
R987 VN.n38 VN.n35 24.4675
R988 VN.n45 VN.n33 24.4675
R989 VN.n43 VN.n42 24.4675
R990 VN.n52 VN.n31 24.4675
R991 VN.n50 VN.n49 24.4675
R992 VN.n57 VN.n56 24.4675
R993 VN.n39 VN.n36 17.9509
R994 VN.n9 VN.n6 17.9509
R995 VN.n22 VN.n21 14.1914
R996 VN.n52 VN.n51 14.1914
R997 VN.n14 VN.n13 12.234
R998 VN.n15 VN.n14 12.234
R999 VN.n45 VN.n44 12.234
R1000 VN.n44 VN.n43 12.234
R1001 VN.n8 VN.n7 10.2766
R1002 VN.n21 VN.n20 10.2766
R1003 VN.n38 VN.n37 10.2766
R1004 VN.n51 VN.n50 10.2766
R1005 VN.n28 VN.n27 8.31928
R1006 VN.n58 VN.n57 8.31928
R1007 VN.n59 VN.n30 0.189894
R1008 VN.n55 VN.n30 0.189894
R1009 VN.n55 VN.n54 0.189894
R1010 VN.n54 VN.n53 0.189894
R1011 VN.n53 VN.n32 0.189894
R1012 VN.n48 VN.n32 0.189894
R1013 VN.n48 VN.n47 0.189894
R1014 VN.n47 VN.n46 0.189894
R1015 VN.n46 VN.n34 0.189894
R1016 VN.n41 VN.n34 0.189894
R1017 VN.n41 VN.n40 0.189894
R1018 VN.n40 VN.n39 0.189894
R1019 VN.n10 VN.n9 0.189894
R1020 VN.n11 VN.n10 0.189894
R1021 VN.n11 VN.n4 0.189894
R1022 VN.n16 VN.n4 0.189894
R1023 VN.n17 VN.n16 0.189894
R1024 VN.n18 VN.n17 0.189894
R1025 VN.n18 VN.n2 0.189894
R1026 VN.n23 VN.n2 0.189894
R1027 VN.n24 VN.n23 0.189894
R1028 VN.n25 VN.n24 0.189894
R1029 VN.n25 VN.n0 0.189894
R1030 VN.n29 VN.n0 0.189894
R1031 VN VN.n29 0.0516364
R1032 VDD2.n169 VDD2.n89 756.745
R1033 VDD2.n80 VDD2.n0 756.745
R1034 VDD2.n170 VDD2.n169 585
R1035 VDD2.n168 VDD2.n167 585
R1036 VDD2.n93 VDD2.n92 585
R1037 VDD2.n97 VDD2.n95 585
R1038 VDD2.n162 VDD2.n161 585
R1039 VDD2.n160 VDD2.n159 585
R1040 VDD2.n99 VDD2.n98 585
R1041 VDD2.n154 VDD2.n153 585
R1042 VDD2.n152 VDD2.n151 585
R1043 VDD2.n103 VDD2.n102 585
R1044 VDD2.n146 VDD2.n145 585
R1045 VDD2.n144 VDD2.n143 585
R1046 VDD2.n107 VDD2.n106 585
R1047 VDD2.n138 VDD2.n137 585
R1048 VDD2.n136 VDD2.n135 585
R1049 VDD2.n111 VDD2.n110 585
R1050 VDD2.n130 VDD2.n129 585
R1051 VDD2.n128 VDD2.n127 585
R1052 VDD2.n115 VDD2.n114 585
R1053 VDD2.n122 VDD2.n121 585
R1054 VDD2.n120 VDD2.n119 585
R1055 VDD2.n29 VDD2.n28 585
R1056 VDD2.n31 VDD2.n30 585
R1057 VDD2.n24 VDD2.n23 585
R1058 VDD2.n37 VDD2.n36 585
R1059 VDD2.n39 VDD2.n38 585
R1060 VDD2.n20 VDD2.n19 585
R1061 VDD2.n45 VDD2.n44 585
R1062 VDD2.n47 VDD2.n46 585
R1063 VDD2.n16 VDD2.n15 585
R1064 VDD2.n53 VDD2.n52 585
R1065 VDD2.n55 VDD2.n54 585
R1066 VDD2.n12 VDD2.n11 585
R1067 VDD2.n61 VDD2.n60 585
R1068 VDD2.n63 VDD2.n62 585
R1069 VDD2.n8 VDD2.n7 585
R1070 VDD2.n70 VDD2.n69 585
R1071 VDD2.n71 VDD2.n6 585
R1072 VDD2.n73 VDD2.n72 585
R1073 VDD2.n4 VDD2.n3 585
R1074 VDD2.n79 VDD2.n78 585
R1075 VDD2.n81 VDD2.n80 585
R1076 VDD2.n118 VDD2.t9 327.466
R1077 VDD2.n27 VDD2.t8 327.466
R1078 VDD2.n169 VDD2.n168 171.744
R1079 VDD2.n168 VDD2.n92 171.744
R1080 VDD2.n97 VDD2.n92 171.744
R1081 VDD2.n161 VDD2.n97 171.744
R1082 VDD2.n161 VDD2.n160 171.744
R1083 VDD2.n160 VDD2.n98 171.744
R1084 VDD2.n153 VDD2.n98 171.744
R1085 VDD2.n153 VDD2.n152 171.744
R1086 VDD2.n152 VDD2.n102 171.744
R1087 VDD2.n145 VDD2.n102 171.744
R1088 VDD2.n145 VDD2.n144 171.744
R1089 VDD2.n144 VDD2.n106 171.744
R1090 VDD2.n137 VDD2.n106 171.744
R1091 VDD2.n137 VDD2.n136 171.744
R1092 VDD2.n136 VDD2.n110 171.744
R1093 VDD2.n129 VDD2.n110 171.744
R1094 VDD2.n129 VDD2.n128 171.744
R1095 VDD2.n128 VDD2.n114 171.744
R1096 VDD2.n121 VDD2.n114 171.744
R1097 VDD2.n121 VDD2.n120 171.744
R1098 VDD2.n30 VDD2.n29 171.744
R1099 VDD2.n30 VDD2.n23 171.744
R1100 VDD2.n37 VDD2.n23 171.744
R1101 VDD2.n38 VDD2.n37 171.744
R1102 VDD2.n38 VDD2.n19 171.744
R1103 VDD2.n45 VDD2.n19 171.744
R1104 VDD2.n46 VDD2.n45 171.744
R1105 VDD2.n46 VDD2.n15 171.744
R1106 VDD2.n53 VDD2.n15 171.744
R1107 VDD2.n54 VDD2.n53 171.744
R1108 VDD2.n54 VDD2.n11 171.744
R1109 VDD2.n61 VDD2.n11 171.744
R1110 VDD2.n62 VDD2.n61 171.744
R1111 VDD2.n62 VDD2.n7 171.744
R1112 VDD2.n70 VDD2.n7 171.744
R1113 VDD2.n71 VDD2.n70 171.744
R1114 VDD2.n72 VDD2.n71 171.744
R1115 VDD2.n72 VDD2.n3 171.744
R1116 VDD2.n79 VDD2.n3 171.744
R1117 VDD2.n80 VDD2.n79 171.744
R1118 VDD2.n120 VDD2.t9 85.8723
R1119 VDD2.n29 VDD2.t8 85.8723
R1120 VDD2.n88 VDD2.n87 72.0517
R1121 VDD2 VDD2.n177 72.0488
R1122 VDD2.n176 VDD2.n175 70.84
R1123 VDD2.n86 VDD2.n85 70.8398
R1124 VDD2.n86 VDD2.n84 51.1356
R1125 VDD2.n174 VDD2.n173 49.446
R1126 VDD2.n174 VDD2.n88 45.0084
R1127 VDD2.n119 VDD2.n118 16.3895
R1128 VDD2.n28 VDD2.n27 16.3895
R1129 VDD2.n95 VDD2.n93 13.1884
R1130 VDD2.n73 VDD2.n4 13.1884
R1131 VDD2.n167 VDD2.n166 12.8005
R1132 VDD2.n163 VDD2.n162 12.8005
R1133 VDD2.n122 VDD2.n117 12.8005
R1134 VDD2.n31 VDD2.n26 12.8005
R1135 VDD2.n74 VDD2.n6 12.8005
R1136 VDD2.n78 VDD2.n77 12.8005
R1137 VDD2.n170 VDD2.n91 12.0247
R1138 VDD2.n159 VDD2.n96 12.0247
R1139 VDD2.n123 VDD2.n115 12.0247
R1140 VDD2.n32 VDD2.n24 12.0247
R1141 VDD2.n69 VDD2.n68 12.0247
R1142 VDD2.n81 VDD2.n2 12.0247
R1143 VDD2.n171 VDD2.n89 11.249
R1144 VDD2.n158 VDD2.n99 11.249
R1145 VDD2.n127 VDD2.n126 11.249
R1146 VDD2.n36 VDD2.n35 11.249
R1147 VDD2.n67 VDD2.n8 11.249
R1148 VDD2.n82 VDD2.n0 11.249
R1149 VDD2.n155 VDD2.n154 10.4732
R1150 VDD2.n130 VDD2.n113 10.4732
R1151 VDD2.n39 VDD2.n22 10.4732
R1152 VDD2.n64 VDD2.n63 10.4732
R1153 VDD2.n151 VDD2.n101 9.69747
R1154 VDD2.n131 VDD2.n111 9.69747
R1155 VDD2.n40 VDD2.n20 9.69747
R1156 VDD2.n60 VDD2.n10 9.69747
R1157 VDD2.n173 VDD2.n172 9.45567
R1158 VDD2.n84 VDD2.n83 9.45567
R1159 VDD2.n105 VDD2.n104 9.3005
R1160 VDD2.n148 VDD2.n147 9.3005
R1161 VDD2.n150 VDD2.n149 9.3005
R1162 VDD2.n101 VDD2.n100 9.3005
R1163 VDD2.n156 VDD2.n155 9.3005
R1164 VDD2.n158 VDD2.n157 9.3005
R1165 VDD2.n96 VDD2.n94 9.3005
R1166 VDD2.n164 VDD2.n163 9.3005
R1167 VDD2.n172 VDD2.n171 9.3005
R1168 VDD2.n91 VDD2.n90 9.3005
R1169 VDD2.n166 VDD2.n165 9.3005
R1170 VDD2.n142 VDD2.n141 9.3005
R1171 VDD2.n140 VDD2.n139 9.3005
R1172 VDD2.n109 VDD2.n108 9.3005
R1173 VDD2.n134 VDD2.n133 9.3005
R1174 VDD2.n132 VDD2.n131 9.3005
R1175 VDD2.n113 VDD2.n112 9.3005
R1176 VDD2.n126 VDD2.n125 9.3005
R1177 VDD2.n124 VDD2.n123 9.3005
R1178 VDD2.n117 VDD2.n116 9.3005
R1179 VDD2.n83 VDD2.n82 9.3005
R1180 VDD2.n2 VDD2.n1 9.3005
R1181 VDD2.n77 VDD2.n76 9.3005
R1182 VDD2.n49 VDD2.n48 9.3005
R1183 VDD2.n18 VDD2.n17 9.3005
R1184 VDD2.n43 VDD2.n42 9.3005
R1185 VDD2.n41 VDD2.n40 9.3005
R1186 VDD2.n22 VDD2.n21 9.3005
R1187 VDD2.n35 VDD2.n34 9.3005
R1188 VDD2.n33 VDD2.n32 9.3005
R1189 VDD2.n26 VDD2.n25 9.3005
R1190 VDD2.n51 VDD2.n50 9.3005
R1191 VDD2.n14 VDD2.n13 9.3005
R1192 VDD2.n57 VDD2.n56 9.3005
R1193 VDD2.n59 VDD2.n58 9.3005
R1194 VDD2.n10 VDD2.n9 9.3005
R1195 VDD2.n65 VDD2.n64 9.3005
R1196 VDD2.n67 VDD2.n66 9.3005
R1197 VDD2.n68 VDD2.n5 9.3005
R1198 VDD2.n75 VDD2.n74 9.3005
R1199 VDD2.n150 VDD2.n103 8.92171
R1200 VDD2.n135 VDD2.n134 8.92171
R1201 VDD2.n44 VDD2.n43 8.92171
R1202 VDD2.n59 VDD2.n12 8.92171
R1203 VDD2.n147 VDD2.n146 8.14595
R1204 VDD2.n138 VDD2.n109 8.14595
R1205 VDD2.n47 VDD2.n18 8.14595
R1206 VDD2.n56 VDD2.n55 8.14595
R1207 VDD2.n143 VDD2.n105 7.3702
R1208 VDD2.n139 VDD2.n107 7.3702
R1209 VDD2.n48 VDD2.n16 7.3702
R1210 VDD2.n52 VDD2.n14 7.3702
R1211 VDD2.n143 VDD2.n142 6.59444
R1212 VDD2.n142 VDD2.n107 6.59444
R1213 VDD2.n51 VDD2.n16 6.59444
R1214 VDD2.n52 VDD2.n51 6.59444
R1215 VDD2.n146 VDD2.n105 5.81868
R1216 VDD2.n139 VDD2.n138 5.81868
R1217 VDD2.n48 VDD2.n47 5.81868
R1218 VDD2.n55 VDD2.n14 5.81868
R1219 VDD2.n147 VDD2.n103 5.04292
R1220 VDD2.n135 VDD2.n109 5.04292
R1221 VDD2.n44 VDD2.n18 5.04292
R1222 VDD2.n56 VDD2.n12 5.04292
R1223 VDD2.n151 VDD2.n150 4.26717
R1224 VDD2.n134 VDD2.n111 4.26717
R1225 VDD2.n43 VDD2.n20 4.26717
R1226 VDD2.n60 VDD2.n59 4.26717
R1227 VDD2.n118 VDD2.n116 3.70982
R1228 VDD2.n27 VDD2.n25 3.70982
R1229 VDD2.n154 VDD2.n101 3.49141
R1230 VDD2.n131 VDD2.n130 3.49141
R1231 VDD2.n40 VDD2.n39 3.49141
R1232 VDD2.n63 VDD2.n10 3.49141
R1233 VDD2.n173 VDD2.n89 2.71565
R1234 VDD2.n155 VDD2.n99 2.71565
R1235 VDD2.n127 VDD2.n113 2.71565
R1236 VDD2.n36 VDD2.n22 2.71565
R1237 VDD2.n64 VDD2.n8 2.71565
R1238 VDD2.n84 VDD2.n0 2.71565
R1239 VDD2.n177 VDD2.t1 2.11259
R1240 VDD2.n177 VDD2.t6 2.11259
R1241 VDD2.n175 VDD2.t3 2.11259
R1242 VDD2.n175 VDD2.t7 2.11259
R1243 VDD2.n87 VDD2.t2 2.11259
R1244 VDD2.n87 VDD2.t0 2.11259
R1245 VDD2.n85 VDD2.t4 2.11259
R1246 VDD2.n85 VDD2.t5 2.11259
R1247 VDD2.n171 VDD2.n170 1.93989
R1248 VDD2.n159 VDD2.n158 1.93989
R1249 VDD2.n126 VDD2.n115 1.93989
R1250 VDD2.n35 VDD2.n24 1.93989
R1251 VDD2.n69 VDD2.n67 1.93989
R1252 VDD2.n82 VDD2.n81 1.93989
R1253 VDD2.n176 VDD2.n174 1.69016
R1254 VDD2.n167 VDD2.n91 1.16414
R1255 VDD2.n162 VDD2.n96 1.16414
R1256 VDD2.n123 VDD2.n122 1.16414
R1257 VDD2.n32 VDD2.n31 1.16414
R1258 VDD2.n68 VDD2.n6 1.16414
R1259 VDD2.n78 VDD2.n2 1.16414
R1260 VDD2 VDD2.n176 0.481103
R1261 VDD2.n166 VDD2.n93 0.388379
R1262 VDD2.n163 VDD2.n95 0.388379
R1263 VDD2.n119 VDD2.n117 0.388379
R1264 VDD2.n28 VDD2.n26 0.388379
R1265 VDD2.n74 VDD2.n73 0.388379
R1266 VDD2.n77 VDD2.n4 0.388379
R1267 VDD2.n88 VDD2.n86 0.367568
R1268 VDD2.n172 VDD2.n90 0.155672
R1269 VDD2.n165 VDD2.n90 0.155672
R1270 VDD2.n165 VDD2.n164 0.155672
R1271 VDD2.n164 VDD2.n94 0.155672
R1272 VDD2.n157 VDD2.n94 0.155672
R1273 VDD2.n157 VDD2.n156 0.155672
R1274 VDD2.n156 VDD2.n100 0.155672
R1275 VDD2.n149 VDD2.n100 0.155672
R1276 VDD2.n149 VDD2.n148 0.155672
R1277 VDD2.n148 VDD2.n104 0.155672
R1278 VDD2.n141 VDD2.n104 0.155672
R1279 VDD2.n141 VDD2.n140 0.155672
R1280 VDD2.n140 VDD2.n108 0.155672
R1281 VDD2.n133 VDD2.n108 0.155672
R1282 VDD2.n133 VDD2.n132 0.155672
R1283 VDD2.n132 VDD2.n112 0.155672
R1284 VDD2.n125 VDD2.n112 0.155672
R1285 VDD2.n125 VDD2.n124 0.155672
R1286 VDD2.n124 VDD2.n116 0.155672
R1287 VDD2.n33 VDD2.n25 0.155672
R1288 VDD2.n34 VDD2.n33 0.155672
R1289 VDD2.n34 VDD2.n21 0.155672
R1290 VDD2.n41 VDD2.n21 0.155672
R1291 VDD2.n42 VDD2.n41 0.155672
R1292 VDD2.n42 VDD2.n17 0.155672
R1293 VDD2.n49 VDD2.n17 0.155672
R1294 VDD2.n50 VDD2.n49 0.155672
R1295 VDD2.n50 VDD2.n13 0.155672
R1296 VDD2.n57 VDD2.n13 0.155672
R1297 VDD2.n58 VDD2.n57 0.155672
R1298 VDD2.n58 VDD2.n9 0.155672
R1299 VDD2.n65 VDD2.n9 0.155672
R1300 VDD2.n66 VDD2.n65 0.155672
R1301 VDD2.n66 VDD2.n5 0.155672
R1302 VDD2.n75 VDD2.n5 0.155672
R1303 VDD2.n76 VDD2.n75 0.155672
R1304 VDD2.n76 VDD2.n1 0.155672
R1305 VDD2.n83 VDD2.n1 0.155672
R1306 B.n440 B.n439 585
R1307 B.n438 B.n127 585
R1308 B.n437 B.n436 585
R1309 B.n435 B.n128 585
R1310 B.n434 B.n433 585
R1311 B.n432 B.n129 585
R1312 B.n431 B.n430 585
R1313 B.n429 B.n130 585
R1314 B.n428 B.n427 585
R1315 B.n426 B.n131 585
R1316 B.n425 B.n424 585
R1317 B.n423 B.n132 585
R1318 B.n422 B.n421 585
R1319 B.n420 B.n133 585
R1320 B.n419 B.n418 585
R1321 B.n417 B.n134 585
R1322 B.n416 B.n415 585
R1323 B.n414 B.n135 585
R1324 B.n413 B.n412 585
R1325 B.n411 B.n136 585
R1326 B.n410 B.n409 585
R1327 B.n408 B.n137 585
R1328 B.n407 B.n406 585
R1329 B.n405 B.n138 585
R1330 B.n404 B.n403 585
R1331 B.n402 B.n139 585
R1332 B.n401 B.n400 585
R1333 B.n399 B.n140 585
R1334 B.n398 B.n397 585
R1335 B.n396 B.n141 585
R1336 B.n395 B.n394 585
R1337 B.n393 B.n142 585
R1338 B.n392 B.n391 585
R1339 B.n390 B.n143 585
R1340 B.n389 B.n388 585
R1341 B.n387 B.n144 585
R1342 B.n386 B.n385 585
R1343 B.n384 B.n145 585
R1344 B.n383 B.n382 585
R1345 B.n381 B.n146 585
R1346 B.n380 B.n379 585
R1347 B.n378 B.n147 585
R1348 B.n377 B.n376 585
R1349 B.n375 B.n148 585
R1350 B.n374 B.n373 585
R1351 B.n372 B.n149 585
R1352 B.n371 B.n370 585
R1353 B.n369 B.n150 585
R1354 B.n368 B.n367 585
R1355 B.n366 B.n151 585
R1356 B.n365 B.n364 585
R1357 B.n363 B.n152 585
R1358 B.n362 B.n361 585
R1359 B.n357 B.n153 585
R1360 B.n356 B.n355 585
R1361 B.n354 B.n154 585
R1362 B.n353 B.n352 585
R1363 B.n351 B.n155 585
R1364 B.n350 B.n349 585
R1365 B.n348 B.n156 585
R1366 B.n347 B.n346 585
R1367 B.n344 B.n157 585
R1368 B.n343 B.n342 585
R1369 B.n341 B.n160 585
R1370 B.n340 B.n339 585
R1371 B.n338 B.n161 585
R1372 B.n337 B.n336 585
R1373 B.n335 B.n162 585
R1374 B.n334 B.n333 585
R1375 B.n332 B.n163 585
R1376 B.n331 B.n330 585
R1377 B.n329 B.n164 585
R1378 B.n328 B.n327 585
R1379 B.n326 B.n165 585
R1380 B.n325 B.n324 585
R1381 B.n323 B.n166 585
R1382 B.n322 B.n321 585
R1383 B.n320 B.n167 585
R1384 B.n319 B.n318 585
R1385 B.n317 B.n168 585
R1386 B.n316 B.n315 585
R1387 B.n314 B.n169 585
R1388 B.n313 B.n312 585
R1389 B.n311 B.n170 585
R1390 B.n310 B.n309 585
R1391 B.n308 B.n171 585
R1392 B.n307 B.n306 585
R1393 B.n305 B.n172 585
R1394 B.n304 B.n303 585
R1395 B.n302 B.n173 585
R1396 B.n301 B.n300 585
R1397 B.n299 B.n174 585
R1398 B.n298 B.n297 585
R1399 B.n296 B.n175 585
R1400 B.n295 B.n294 585
R1401 B.n293 B.n176 585
R1402 B.n292 B.n291 585
R1403 B.n290 B.n177 585
R1404 B.n289 B.n288 585
R1405 B.n287 B.n178 585
R1406 B.n286 B.n285 585
R1407 B.n284 B.n179 585
R1408 B.n283 B.n282 585
R1409 B.n281 B.n180 585
R1410 B.n280 B.n279 585
R1411 B.n278 B.n181 585
R1412 B.n277 B.n276 585
R1413 B.n275 B.n182 585
R1414 B.n274 B.n273 585
R1415 B.n272 B.n183 585
R1416 B.n271 B.n270 585
R1417 B.n269 B.n184 585
R1418 B.n268 B.n267 585
R1419 B.n441 B.n126 585
R1420 B.n443 B.n442 585
R1421 B.n444 B.n125 585
R1422 B.n446 B.n445 585
R1423 B.n447 B.n124 585
R1424 B.n449 B.n448 585
R1425 B.n450 B.n123 585
R1426 B.n452 B.n451 585
R1427 B.n453 B.n122 585
R1428 B.n455 B.n454 585
R1429 B.n456 B.n121 585
R1430 B.n458 B.n457 585
R1431 B.n459 B.n120 585
R1432 B.n461 B.n460 585
R1433 B.n462 B.n119 585
R1434 B.n464 B.n463 585
R1435 B.n465 B.n118 585
R1436 B.n467 B.n466 585
R1437 B.n468 B.n117 585
R1438 B.n470 B.n469 585
R1439 B.n471 B.n116 585
R1440 B.n473 B.n472 585
R1441 B.n474 B.n115 585
R1442 B.n476 B.n475 585
R1443 B.n477 B.n114 585
R1444 B.n479 B.n478 585
R1445 B.n480 B.n113 585
R1446 B.n482 B.n481 585
R1447 B.n483 B.n112 585
R1448 B.n485 B.n484 585
R1449 B.n486 B.n111 585
R1450 B.n488 B.n487 585
R1451 B.n489 B.n110 585
R1452 B.n491 B.n490 585
R1453 B.n492 B.n109 585
R1454 B.n494 B.n493 585
R1455 B.n495 B.n108 585
R1456 B.n497 B.n496 585
R1457 B.n498 B.n107 585
R1458 B.n500 B.n499 585
R1459 B.n501 B.n106 585
R1460 B.n503 B.n502 585
R1461 B.n504 B.n105 585
R1462 B.n506 B.n505 585
R1463 B.n507 B.n104 585
R1464 B.n509 B.n508 585
R1465 B.n510 B.n103 585
R1466 B.n512 B.n511 585
R1467 B.n513 B.n102 585
R1468 B.n515 B.n514 585
R1469 B.n516 B.n101 585
R1470 B.n518 B.n517 585
R1471 B.n519 B.n100 585
R1472 B.n521 B.n520 585
R1473 B.n522 B.n99 585
R1474 B.n524 B.n523 585
R1475 B.n525 B.n98 585
R1476 B.n527 B.n526 585
R1477 B.n528 B.n97 585
R1478 B.n530 B.n529 585
R1479 B.n531 B.n96 585
R1480 B.n533 B.n532 585
R1481 B.n534 B.n95 585
R1482 B.n536 B.n535 585
R1483 B.n537 B.n94 585
R1484 B.n539 B.n538 585
R1485 B.n540 B.n93 585
R1486 B.n542 B.n541 585
R1487 B.n543 B.n92 585
R1488 B.n545 B.n544 585
R1489 B.n546 B.n91 585
R1490 B.n548 B.n547 585
R1491 B.n549 B.n90 585
R1492 B.n551 B.n550 585
R1493 B.n552 B.n89 585
R1494 B.n554 B.n553 585
R1495 B.n555 B.n88 585
R1496 B.n557 B.n556 585
R1497 B.n558 B.n87 585
R1498 B.n560 B.n559 585
R1499 B.n561 B.n86 585
R1500 B.n563 B.n562 585
R1501 B.n564 B.n85 585
R1502 B.n566 B.n565 585
R1503 B.n567 B.n84 585
R1504 B.n569 B.n568 585
R1505 B.n740 B.n23 585
R1506 B.n739 B.n738 585
R1507 B.n737 B.n24 585
R1508 B.n736 B.n735 585
R1509 B.n734 B.n25 585
R1510 B.n733 B.n732 585
R1511 B.n731 B.n26 585
R1512 B.n730 B.n729 585
R1513 B.n728 B.n27 585
R1514 B.n727 B.n726 585
R1515 B.n725 B.n28 585
R1516 B.n724 B.n723 585
R1517 B.n722 B.n29 585
R1518 B.n721 B.n720 585
R1519 B.n719 B.n30 585
R1520 B.n718 B.n717 585
R1521 B.n716 B.n31 585
R1522 B.n715 B.n714 585
R1523 B.n713 B.n32 585
R1524 B.n712 B.n711 585
R1525 B.n710 B.n33 585
R1526 B.n709 B.n708 585
R1527 B.n707 B.n34 585
R1528 B.n706 B.n705 585
R1529 B.n704 B.n35 585
R1530 B.n703 B.n702 585
R1531 B.n701 B.n36 585
R1532 B.n700 B.n699 585
R1533 B.n698 B.n37 585
R1534 B.n697 B.n696 585
R1535 B.n695 B.n38 585
R1536 B.n694 B.n693 585
R1537 B.n692 B.n39 585
R1538 B.n691 B.n690 585
R1539 B.n689 B.n40 585
R1540 B.n688 B.n687 585
R1541 B.n686 B.n41 585
R1542 B.n685 B.n684 585
R1543 B.n683 B.n42 585
R1544 B.n682 B.n681 585
R1545 B.n680 B.n43 585
R1546 B.n679 B.n678 585
R1547 B.n677 B.n44 585
R1548 B.n676 B.n675 585
R1549 B.n674 B.n45 585
R1550 B.n673 B.n672 585
R1551 B.n671 B.n46 585
R1552 B.n670 B.n669 585
R1553 B.n668 B.n47 585
R1554 B.n667 B.n666 585
R1555 B.n665 B.n48 585
R1556 B.n664 B.n663 585
R1557 B.n661 B.n49 585
R1558 B.n660 B.n659 585
R1559 B.n658 B.n52 585
R1560 B.n657 B.n656 585
R1561 B.n655 B.n53 585
R1562 B.n654 B.n653 585
R1563 B.n652 B.n54 585
R1564 B.n651 B.n650 585
R1565 B.n649 B.n55 585
R1566 B.n647 B.n646 585
R1567 B.n645 B.n58 585
R1568 B.n644 B.n643 585
R1569 B.n642 B.n59 585
R1570 B.n641 B.n640 585
R1571 B.n639 B.n60 585
R1572 B.n638 B.n637 585
R1573 B.n636 B.n61 585
R1574 B.n635 B.n634 585
R1575 B.n633 B.n62 585
R1576 B.n632 B.n631 585
R1577 B.n630 B.n63 585
R1578 B.n629 B.n628 585
R1579 B.n627 B.n64 585
R1580 B.n626 B.n625 585
R1581 B.n624 B.n65 585
R1582 B.n623 B.n622 585
R1583 B.n621 B.n66 585
R1584 B.n620 B.n619 585
R1585 B.n618 B.n67 585
R1586 B.n617 B.n616 585
R1587 B.n615 B.n68 585
R1588 B.n614 B.n613 585
R1589 B.n612 B.n69 585
R1590 B.n611 B.n610 585
R1591 B.n609 B.n70 585
R1592 B.n608 B.n607 585
R1593 B.n606 B.n71 585
R1594 B.n605 B.n604 585
R1595 B.n603 B.n72 585
R1596 B.n602 B.n601 585
R1597 B.n600 B.n73 585
R1598 B.n599 B.n598 585
R1599 B.n597 B.n74 585
R1600 B.n596 B.n595 585
R1601 B.n594 B.n75 585
R1602 B.n593 B.n592 585
R1603 B.n591 B.n76 585
R1604 B.n590 B.n589 585
R1605 B.n588 B.n77 585
R1606 B.n587 B.n586 585
R1607 B.n585 B.n78 585
R1608 B.n584 B.n583 585
R1609 B.n582 B.n79 585
R1610 B.n581 B.n580 585
R1611 B.n579 B.n80 585
R1612 B.n578 B.n577 585
R1613 B.n576 B.n81 585
R1614 B.n575 B.n574 585
R1615 B.n573 B.n82 585
R1616 B.n572 B.n571 585
R1617 B.n570 B.n83 585
R1618 B.n742 B.n741 585
R1619 B.n743 B.n22 585
R1620 B.n745 B.n744 585
R1621 B.n746 B.n21 585
R1622 B.n748 B.n747 585
R1623 B.n749 B.n20 585
R1624 B.n751 B.n750 585
R1625 B.n752 B.n19 585
R1626 B.n754 B.n753 585
R1627 B.n755 B.n18 585
R1628 B.n757 B.n756 585
R1629 B.n758 B.n17 585
R1630 B.n760 B.n759 585
R1631 B.n761 B.n16 585
R1632 B.n763 B.n762 585
R1633 B.n764 B.n15 585
R1634 B.n766 B.n765 585
R1635 B.n767 B.n14 585
R1636 B.n769 B.n768 585
R1637 B.n770 B.n13 585
R1638 B.n772 B.n771 585
R1639 B.n773 B.n12 585
R1640 B.n775 B.n774 585
R1641 B.n776 B.n11 585
R1642 B.n778 B.n777 585
R1643 B.n779 B.n10 585
R1644 B.n781 B.n780 585
R1645 B.n782 B.n9 585
R1646 B.n784 B.n783 585
R1647 B.n785 B.n8 585
R1648 B.n787 B.n786 585
R1649 B.n788 B.n7 585
R1650 B.n790 B.n789 585
R1651 B.n791 B.n6 585
R1652 B.n793 B.n792 585
R1653 B.n794 B.n5 585
R1654 B.n796 B.n795 585
R1655 B.n797 B.n4 585
R1656 B.n799 B.n798 585
R1657 B.n800 B.n3 585
R1658 B.n802 B.n801 585
R1659 B.n803 B.n0 585
R1660 B.n2 B.n1 585
R1661 B.n206 B.n205 585
R1662 B.n208 B.n207 585
R1663 B.n209 B.n204 585
R1664 B.n211 B.n210 585
R1665 B.n212 B.n203 585
R1666 B.n214 B.n213 585
R1667 B.n215 B.n202 585
R1668 B.n217 B.n216 585
R1669 B.n218 B.n201 585
R1670 B.n220 B.n219 585
R1671 B.n221 B.n200 585
R1672 B.n223 B.n222 585
R1673 B.n224 B.n199 585
R1674 B.n226 B.n225 585
R1675 B.n227 B.n198 585
R1676 B.n229 B.n228 585
R1677 B.n230 B.n197 585
R1678 B.n232 B.n231 585
R1679 B.n233 B.n196 585
R1680 B.n235 B.n234 585
R1681 B.n236 B.n195 585
R1682 B.n238 B.n237 585
R1683 B.n239 B.n194 585
R1684 B.n241 B.n240 585
R1685 B.n242 B.n193 585
R1686 B.n244 B.n243 585
R1687 B.n245 B.n192 585
R1688 B.n247 B.n246 585
R1689 B.n248 B.n191 585
R1690 B.n250 B.n249 585
R1691 B.n251 B.n190 585
R1692 B.n253 B.n252 585
R1693 B.n254 B.n189 585
R1694 B.n256 B.n255 585
R1695 B.n257 B.n188 585
R1696 B.n259 B.n258 585
R1697 B.n260 B.n187 585
R1698 B.n262 B.n261 585
R1699 B.n263 B.n186 585
R1700 B.n265 B.n264 585
R1701 B.n266 B.n185 585
R1702 B.n268 B.n185 511.721
R1703 B.n441 B.n440 511.721
R1704 B.n568 B.n83 511.721
R1705 B.n742 B.n23 511.721
R1706 B.n358 B.t10 474.587
R1707 B.n56 B.t5 474.587
R1708 B.n158 B.t7 474.587
R1709 B.n50 B.t2 474.587
R1710 B.n359 B.t11 436.575
R1711 B.n57 B.t4 436.575
R1712 B.n159 B.t8 436.575
R1713 B.n51 B.t1 436.575
R1714 B.n158 B.t6 433.438
R1715 B.n358 B.t9 433.438
R1716 B.n56 B.t3 433.438
R1717 B.n50 B.t0 433.438
R1718 B.n805 B.n804 256.663
R1719 B.n804 B.n803 235.042
R1720 B.n804 B.n2 235.042
R1721 B.n269 B.n268 163.367
R1722 B.n270 B.n269 163.367
R1723 B.n270 B.n183 163.367
R1724 B.n274 B.n183 163.367
R1725 B.n275 B.n274 163.367
R1726 B.n276 B.n275 163.367
R1727 B.n276 B.n181 163.367
R1728 B.n280 B.n181 163.367
R1729 B.n281 B.n280 163.367
R1730 B.n282 B.n281 163.367
R1731 B.n282 B.n179 163.367
R1732 B.n286 B.n179 163.367
R1733 B.n287 B.n286 163.367
R1734 B.n288 B.n287 163.367
R1735 B.n288 B.n177 163.367
R1736 B.n292 B.n177 163.367
R1737 B.n293 B.n292 163.367
R1738 B.n294 B.n293 163.367
R1739 B.n294 B.n175 163.367
R1740 B.n298 B.n175 163.367
R1741 B.n299 B.n298 163.367
R1742 B.n300 B.n299 163.367
R1743 B.n300 B.n173 163.367
R1744 B.n304 B.n173 163.367
R1745 B.n305 B.n304 163.367
R1746 B.n306 B.n305 163.367
R1747 B.n306 B.n171 163.367
R1748 B.n310 B.n171 163.367
R1749 B.n311 B.n310 163.367
R1750 B.n312 B.n311 163.367
R1751 B.n312 B.n169 163.367
R1752 B.n316 B.n169 163.367
R1753 B.n317 B.n316 163.367
R1754 B.n318 B.n317 163.367
R1755 B.n318 B.n167 163.367
R1756 B.n322 B.n167 163.367
R1757 B.n323 B.n322 163.367
R1758 B.n324 B.n323 163.367
R1759 B.n324 B.n165 163.367
R1760 B.n328 B.n165 163.367
R1761 B.n329 B.n328 163.367
R1762 B.n330 B.n329 163.367
R1763 B.n330 B.n163 163.367
R1764 B.n334 B.n163 163.367
R1765 B.n335 B.n334 163.367
R1766 B.n336 B.n335 163.367
R1767 B.n336 B.n161 163.367
R1768 B.n340 B.n161 163.367
R1769 B.n341 B.n340 163.367
R1770 B.n342 B.n341 163.367
R1771 B.n342 B.n157 163.367
R1772 B.n347 B.n157 163.367
R1773 B.n348 B.n347 163.367
R1774 B.n349 B.n348 163.367
R1775 B.n349 B.n155 163.367
R1776 B.n353 B.n155 163.367
R1777 B.n354 B.n353 163.367
R1778 B.n355 B.n354 163.367
R1779 B.n355 B.n153 163.367
R1780 B.n362 B.n153 163.367
R1781 B.n363 B.n362 163.367
R1782 B.n364 B.n363 163.367
R1783 B.n364 B.n151 163.367
R1784 B.n368 B.n151 163.367
R1785 B.n369 B.n368 163.367
R1786 B.n370 B.n369 163.367
R1787 B.n370 B.n149 163.367
R1788 B.n374 B.n149 163.367
R1789 B.n375 B.n374 163.367
R1790 B.n376 B.n375 163.367
R1791 B.n376 B.n147 163.367
R1792 B.n380 B.n147 163.367
R1793 B.n381 B.n380 163.367
R1794 B.n382 B.n381 163.367
R1795 B.n382 B.n145 163.367
R1796 B.n386 B.n145 163.367
R1797 B.n387 B.n386 163.367
R1798 B.n388 B.n387 163.367
R1799 B.n388 B.n143 163.367
R1800 B.n392 B.n143 163.367
R1801 B.n393 B.n392 163.367
R1802 B.n394 B.n393 163.367
R1803 B.n394 B.n141 163.367
R1804 B.n398 B.n141 163.367
R1805 B.n399 B.n398 163.367
R1806 B.n400 B.n399 163.367
R1807 B.n400 B.n139 163.367
R1808 B.n404 B.n139 163.367
R1809 B.n405 B.n404 163.367
R1810 B.n406 B.n405 163.367
R1811 B.n406 B.n137 163.367
R1812 B.n410 B.n137 163.367
R1813 B.n411 B.n410 163.367
R1814 B.n412 B.n411 163.367
R1815 B.n412 B.n135 163.367
R1816 B.n416 B.n135 163.367
R1817 B.n417 B.n416 163.367
R1818 B.n418 B.n417 163.367
R1819 B.n418 B.n133 163.367
R1820 B.n422 B.n133 163.367
R1821 B.n423 B.n422 163.367
R1822 B.n424 B.n423 163.367
R1823 B.n424 B.n131 163.367
R1824 B.n428 B.n131 163.367
R1825 B.n429 B.n428 163.367
R1826 B.n430 B.n429 163.367
R1827 B.n430 B.n129 163.367
R1828 B.n434 B.n129 163.367
R1829 B.n435 B.n434 163.367
R1830 B.n436 B.n435 163.367
R1831 B.n436 B.n127 163.367
R1832 B.n440 B.n127 163.367
R1833 B.n568 B.n567 163.367
R1834 B.n567 B.n566 163.367
R1835 B.n566 B.n85 163.367
R1836 B.n562 B.n85 163.367
R1837 B.n562 B.n561 163.367
R1838 B.n561 B.n560 163.367
R1839 B.n560 B.n87 163.367
R1840 B.n556 B.n87 163.367
R1841 B.n556 B.n555 163.367
R1842 B.n555 B.n554 163.367
R1843 B.n554 B.n89 163.367
R1844 B.n550 B.n89 163.367
R1845 B.n550 B.n549 163.367
R1846 B.n549 B.n548 163.367
R1847 B.n548 B.n91 163.367
R1848 B.n544 B.n91 163.367
R1849 B.n544 B.n543 163.367
R1850 B.n543 B.n542 163.367
R1851 B.n542 B.n93 163.367
R1852 B.n538 B.n93 163.367
R1853 B.n538 B.n537 163.367
R1854 B.n537 B.n536 163.367
R1855 B.n536 B.n95 163.367
R1856 B.n532 B.n95 163.367
R1857 B.n532 B.n531 163.367
R1858 B.n531 B.n530 163.367
R1859 B.n530 B.n97 163.367
R1860 B.n526 B.n97 163.367
R1861 B.n526 B.n525 163.367
R1862 B.n525 B.n524 163.367
R1863 B.n524 B.n99 163.367
R1864 B.n520 B.n99 163.367
R1865 B.n520 B.n519 163.367
R1866 B.n519 B.n518 163.367
R1867 B.n518 B.n101 163.367
R1868 B.n514 B.n101 163.367
R1869 B.n514 B.n513 163.367
R1870 B.n513 B.n512 163.367
R1871 B.n512 B.n103 163.367
R1872 B.n508 B.n103 163.367
R1873 B.n508 B.n507 163.367
R1874 B.n507 B.n506 163.367
R1875 B.n506 B.n105 163.367
R1876 B.n502 B.n105 163.367
R1877 B.n502 B.n501 163.367
R1878 B.n501 B.n500 163.367
R1879 B.n500 B.n107 163.367
R1880 B.n496 B.n107 163.367
R1881 B.n496 B.n495 163.367
R1882 B.n495 B.n494 163.367
R1883 B.n494 B.n109 163.367
R1884 B.n490 B.n109 163.367
R1885 B.n490 B.n489 163.367
R1886 B.n489 B.n488 163.367
R1887 B.n488 B.n111 163.367
R1888 B.n484 B.n111 163.367
R1889 B.n484 B.n483 163.367
R1890 B.n483 B.n482 163.367
R1891 B.n482 B.n113 163.367
R1892 B.n478 B.n113 163.367
R1893 B.n478 B.n477 163.367
R1894 B.n477 B.n476 163.367
R1895 B.n476 B.n115 163.367
R1896 B.n472 B.n115 163.367
R1897 B.n472 B.n471 163.367
R1898 B.n471 B.n470 163.367
R1899 B.n470 B.n117 163.367
R1900 B.n466 B.n117 163.367
R1901 B.n466 B.n465 163.367
R1902 B.n465 B.n464 163.367
R1903 B.n464 B.n119 163.367
R1904 B.n460 B.n119 163.367
R1905 B.n460 B.n459 163.367
R1906 B.n459 B.n458 163.367
R1907 B.n458 B.n121 163.367
R1908 B.n454 B.n121 163.367
R1909 B.n454 B.n453 163.367
R1910 B.n453 B.n452 163.367
R1911 B.n452 B.n123 163.367
R1912 B.n448 B.n123 163.367
R1913 B.n448 B.n447 163.367
R1914 B.n447 B.n446 163.367
R1915 B.n446 B.n125 163.367
R1916 B.n442 B.n125 163.367
R1917 B.n442 B.n441 163.367
R1918 B.n738 B.n23 163.367
R1919 B.n738 B.n737 163.367
R1920 B.n737 B.n736 163.367
R1921 B.n736 B.n25 163.367
R1922 B.n732 B.n25 163.367
R1923 B.n732 B.n731 163.367
R1924 B.n731 B.n730 163.367
R1925 B.n730 B.n27 163.367
R1926 B.n726 B.n27 163.367
R1927 B.n726 B.n725 163.367
R1928 B.n725 B.n724 163.367
R1929 B.n724 B.n29 163.367
R1930 B.n720 B.n29 163.367
R1931 B.n720 B.n719 163.367
R1932 B.n719 B.n718 163.367
R1933 B.n718 B.n31 163.367
R1934 B.n714 B.n31 163.367
R1935 B.n714 B.n713 163.367
R1936 B.n713 B.n712 163.367
R1937 B.n712 B.n33 163.367
R1938 B.n708 B.n33 163.367
R1939 B.n708 B.n707 163.367
R1940 B.n707 B.n706 163.367
R1941 B.n706 B.n35 163.367
R1942 B.n702 B.n35 163.367
R1943 B.n702 B.n701 163.367
R1944 B.n701 B.n700 163.367
R1945 B.n700 B.n37 163.367
R1946 B.n696 B.n37 163.367
R1947 B.n696 B.n695 163.367
R1948 B.n695 B.n694 163.367
R1949 B.n694 B.n39 163.367
R1950 B.n690 B.n39 163.367
R1951 B.n690 B.n689 163.367
R1952 B.n689 B.n688 163.367
R1953 B.n688 B.n41 163.367
R1954 B.n684 B.n41 163.367
R1955 B.n684 B.n683 163.367
R1956 B.n683 B.n682 163.367
R1957 B.n682 B.n43 163.367
R1958 B.n678 B.n43 163.367
R1959 B.n678 B.n677 163.367
R1960 B.n677 B.n676 163.367
R1961 B.n676 B.n45 163.367
R1962 B.n672 B.n45 163.367
R1963 B.n672 B.n671 163.367
R1964 B.n671 B.n670 163.367
R1965 B.n670 B.n47 163.367
R1966 B.n666 B.n47 163.367
R1967 B.n666 B.n665 163.367
R1968 B.n665 B.n664 163.367
R1969 B.n664 B.n49 163.367
R1970 B.n659 B.n49 163.367
R1971 B.n659 B.n658 163.367
R1972 B.n658 B.n657 163.367
R1973 B.n657 B.n53 163.367
R1974 B.n653 B.n53 163.367
R1975 B.n653 B.n652 163.367
R1976 B.n652 B.n651 163.367
R1977 B.n651 B.n55 163.367
R1978 B.n646 B.n55 163.367
R1979 B.n646 B.n645 163.367
R1980 B.n645 B.n644 163.367
R1981 B.n644 B.n59 163.367
R1982 B.n640 B.n59 163.367
R1983 B.n640 B.n639 163.367
R1984 B.n639 B.n638 163.367
R1985 B.n638 B.n61 163.367
R1986 B.n634 B.n61 163.367
R1987 B.n634 B.n633 163.367
R1988 B.n633 B.n632 163.367
R1989 B.n632 B.n63 163.367
R1990 B.n628 B.n63 163.367
R1991 B.n628 B.n627 163.367
R1992 B.n627 B.n626 163.367
R1993 B.n626 B.n65 163.367
R1994 B.n622 B.n65 163.367
R1995 B.n622 B.n621 163.367
R1996 B.n621 B.n620 163.367
R1997 B.n620 B.n67 163.367
R1998 B.n616 B.n67 163.367
R1999 B.n616 B.n615 163.367
R2000 B.n615 B.n614 163.367
R2001 B.n614 B.n69 163.367
R2002 B.n610 B.n69 163.367
R2003 B.n610 B.n609 163.367
R2004 B.n609 B.n608 163.367
R2005 B.n608 B.n71 163.367
R2006 B.n604 B.n71 163.367
R2007 B.n604 B.n603 163.367
R2008 B.n603 B.n602 163.367
R2009 B.n602 B.n73 163.367
R2010 B.n598 B.n73 163.367
R2011 B.n598 B.n597 163.367
R2012 B.n597 B.n596 163.367
R2013 B.n596 B.n75 163.367
R2014 B.n592 B.n75 163.367
R2015 B.n592 B.n591 163.367
R2016 B.n591 B.n590 163.367
R2017 B.n590 B.n77 163.367
R2018 B.n586 B.n77 163.367
R2019 B.n586 B.n585 163.367
R2020 B.n585 B.n584 163.367
R2021 B.n584 B.n79 163.367
R2022 B.n580 B.n79 163.367
R2023 B.n580 B.n579 163.367
R2024 B.n579 B.n578 163.367
R2025 B.n578 B.n81 163.367
R2026 B.n574 B.n81 163.367
R2027 B.n574 B.n573 163.367
R2028 B.n573 B.n572 163.367
R2029 B.n572 B.n83 163.367
R2030 B.n743 B.n742 163.367
R2031 B.n744 B.n743 163.367
R2032 B.n744 B.n21 163.367
R2033 B.n748 B.n21 163.367
R2034 B.n749 B.n748 163.367
R2035 B.n750 B.n749 163.367
R2036 B.n750 B.n19 163.367
R2037 B.n754 B.n19 163.367
R2038 B.n755 B.n754 163.367
R2039 B.n756 B.n755 163.367
R2040 B.n756 B.n17 163.367
R2041 B.n760 B.n17 163.367
R2042 B.n761 B.n760 163.367
R2043 B.n762 B.n761 163.367
R2044 B.n762 B.n15 163.367
R2045 B.n766 B.n15 163.367
R2046 B.n767 B.n766 163.367
R2047 B.n768 B.n767 163.367
R2048 B.n768 B.n13 163.367
R2049 B.n772 B.n13 163.367
R2050 B.n773 B.n772 163.367
R2051 B.n774 B.n773 163.367
R2052 B.n774 B.n11 163.367
R2053 B.n778 B.n11 163.367
R2054 B.n779 B.n778 163.367
R2055 B.n780 B.n779 163.367
R2056 B.n780 B.n9 163.367
R2057 B.n784 B.n9 163.367
R2058 B.n785 B.n784 163.367
R2059 B.n786 B.n785 163.367
R2060 B.n786 B.n7 163.367
R2061 B.n790 B.n7 163.367
R2062 B.n791 B.n790 163.367
R2063 B.n792 B.n791 163.367
R2064 B.n792 B.n5 163.367
R2065 B.n796 B.n5 163.367
R2066 B.n797 B.n796 163.367
R2067 B.n798 B.n797 163.367
R2068 B.n798 B.n3 163.367
R2069 B.n802 B.n3 163.367
R2070 B.n803 B.n802 163.367
R2071 B.n205 B.n2 163.367
R2072 B.n208 B.n205 163.367
R2073 B.n209 B.n208 163.367
R2074 B.n210 B.n209 163.367
R2075 B.n210 B.n203 163.367
R2076 B.n214 B.n203 163.367
R2077 B.n215 B.n214 163.367
R2078 B.n216 B.n215 163.367
R2079 B.n216 B.n201 163.367
R2080 B.n220 B.n201 163.367
R2081 B.n221 B.n220 163.367
R2082 B.n222 B.n221 163.367
R2083 B.n222 B.n199 163.367
R2084 B.n226 B.n199 163.367
R2085 B.n227 B.n226 163.367
R2086 B.n228 B.n227 163.367
R2087 B.n228 B.n197 163.367
R2088 B.n232 B.n197 163.367
R2089 B.n233 B.n232 163.367
R2090 B.n234 B.n233 163.367
R2091 B.n234 B.n195 163.367
R2092 B.n238 B.n195 163.367
R2093 B.n239 B.n238 163.367
R2094 B.n240 B.n239 163.367
R2095 B.n240 B.n193 163.367
R2096 B.n244 B.n193 163.367
R2097 B.n245 B.n244 163.367
R2098 B.n246 B.n245 163.367
R2099 B.n246 B.n191 163.367
R2100 B.n250 B.n191 163.367
R2101 B.n251 B.n250 163.367
R2102 B.n252 B.n251 163.367
R2103 B.n252 B.n189 163.367
R2104 B.n256 B.n189 163.367
R2105 B.n257 B.n256 163.367
R2106 B.n258 B.n257 163.367
R2107 B.n258 B.n187 163.367
R2108 B.n262 B.n187 163.367
R2109 B.n263 B.n262 163.367
R2110 B.n264 B.n263 163.367
R2111 B.n264 B.n185 163.367
R2112 B.n345 B.n159 59.5399
R2113 B.n360 B.n359 59.5399
R2114 B.n648 B.n57 59.5399
R2115 B.n662 B.n51 59.5399
R2116 B.n159 B.n158 38.0126
R2117 B.n359 B.n358 38.0126
R2118 B.n57 B.n56 38.0126
R2119 B.n51 B.n50 38.0126
R2120 B.n741 B.n740 33.2493
R2121 B.n570 B.n569 33.2493
R2122 B.n439 B.n126 33.2493
R2123 B.n267 B.n266 33.2493
R2124 B B.n805 18.0485
R2125 B.n741 B.n22 10.6151
R2126 B.n745 B.n22 10.6151
R2127 B.n746 B.n745 10.6151
R2128 B.n747 B.n746 10.6151
R2129 B.n747 B.n20 10.6151
R2130 B.n751 B.n20 10.6151
R2131 B.n752 B.n751 10.6151
R2132 B.n753 B.n752 10.6151
R2133 B.n753 B.n18 10.6151
R2134 B.n757 B.n18 10.6151
R2135 B.n758 B.n757 10.6151
R2136 B.n759 B.n758 10.6151
R2137 B.n759 B.n16 10.6151
R2138 B.n763 B.n16 10.6151
R2139 B.n764 B.n763 10.6151
R2140 B.n765 B.n764 10.6151
R2141 B.n765 B.n14 10.6151
R2142 B.n769 B.n14 10.6151
R2143 B.n770 B.n769 10.6151
R2144 B.n771 B.n770 10.6151
R2145 B.n771 B.n12 10.6151
R2146 B.n775 B.n12 10.6151
R2147 B.n776 B.n775 10.6151
R2148 B.n777 B.n776 10.6151
R2149 B.n777 B.n10 10.6151
R2150 B.n781 B.n10 10.6151
R2151 B.n782 B.n781 10.6151
R2152 B.n783 B.n782 10.6151
R2153 B.n783 B.n8 10.6151
R2154 B.n787 B.n8 10.6151
R2155 B.n788 B.n787 10.6151
R2156 B.n789 B.n788 10.6151
R2157 B.n789 B.n6 10.6151
R2158 B.n793 B.n6 10.6151
R2159 B.n794 B.n793 10.6151
R2160 B.n795 B.n794 10.6151
R2161 B.n795 B.n4 10.6151
R2162 B.n799 B.n4 10.6151
R2163 B.n800 B.n799 10.6151
R2164 B.n801 B.n800 10.6151
R2165 B.n801 B.n0 10.6151
R2166 B.n740 B.n739 10.6151
R2167 B.n739 B.n24 10.6151
R2168 B.n735 B.n24 10.6151
R2169 B.n735 B.n734 10.6151
R2170 B.n734 B.n733 10.6151
R2171 B.n733 B.n26 10.6151
R2172 B.n729 B.n26 10.6151
R2173 B.n729 B.n728 10.6151
R2174 B.n728 B.n727 10.6151
R2175 B.n727 B.n28 10.6151
R2176 B.n723 B.n28 10.6151
R2177 B.n723 B.n722 10.6151
R2178 B.n722 B.n721 10.6151
R2179 B.n721 B.n30 10.6151
R2180 B.n717 B.n30 10.6151
R2181 B.n717 B.n716 10.6151
R2182 B.n716 B.n715 10.6151
R2183 B.n715 B.n32 10.6151
R2184 B.n711 B.n32 10.6151
R2185 B.n711 B.n710 10.6151
R2186 B.n710 B.n709 10.6151
R2187 B.n709 B.n34 10.6151
R2188 B.n705 B.n34 10.6151
R2189 B.n705 B.n704 10.6151
R2190 B.n704 B.n703 10.6151
R2191 B.n703 B.n36 10.6151
R2192 B.n699 B.n36 10.6151
R2193 B.n699 B.n698 10.6151
R2194 B.n698 B.n697 10.6151
R2195 B.n697 B.n38 10.6151
R2196 B.n693 B.n38 10.6151
R2197 B.n693 B.n692 10.6151
R2198 B.n692 B.n691 10.6151
R2199 B.n691 B.n40 10.6151
R2200 B.n687 B.n40 10.6151
R2201 B.n687 B.n686 10.6151
R2202 B.n686 B.n685 10.6151
R2203 B.n685 B.n42 10.6151
R2204 B.n681 B.n42 10.6151
R2205 B.n681 B.n680 10.6151
R2206 B.n680 B.n679 10.6151
R2207 B.n679 B.n44 10.6151
R2208 B.n675 B.n44 10.6151
R2209 B.n675 B.n674 10.6151
R2210 B.n674 B.n673 10.6151
R2211 B.n673 B.n46 10.6151
R2212 B.n669 B.n46 10.6151
R2213 B.n669 B.n668 10.6151
R2214 B.n668 B.n667 10.6151
R2215 B.n667 B.n48 10.6151
R2216 B.n663 B.n48 10.6151
R2217 B.n661 B.n660 10.6151
R2218 B.n660 B.n52 10.6151
R2219 B.n656 B.n52 10.6151
R2220 B.n656 B.n655 10.6151
R2221 B.n655 B.n654 10.6151
R2222 B.n654 B.n54 10.6151
R2223 B.n650 B.n54 10.6151
R2224 B.n650 B.n649 10.6151
R2225 B.n647 B.n58 10.6151
R2226 B.n643 B.n58 10.6151
R2227 B.n643 B.n642 10.6151
R2228 B.n642 B.n641 10.6151
R2229 B.n641 B.n60 10.6151
R2230 B.n637 B.n60 10.6151
R2231 B.n637 B.n636 10.6151
R2232 B.n636 B.n635 10.6151
R2233 B.n635 B.n62 10.6151
R2234 B.n631 B.n62 10.6151
R2235 B.n631 B.n630 10.6151
R2236 B.n630 B.n629 10.6151
R2237 B.n629 B.n64 10.6151
R2238 B.n625 B.n64 10.6151
R2239 B.n625 B.n624 10.6151
R2240 B.n624 B.n623 10.6151
R2241 B.n623 B.n66 10.6151
R2242 B.n619 B.n66 10.6151
R2243 B.n619 B.n618 10.6151
R2244 B.n618 B.n617 10.6151
R2245 B.n617 B.n68 10.6151
R2246 B.n613 B.n68 10.6151
R2247 B.n613 B.n612 10.6151
R2248 B.n612 B.n611 10.6151
R2249 B.n611 B.n70 10.6151
R2250 B.n607 B.n70 10.6151
R2251 B.n607 B.n606 10.6151
R2252 B.n606 B.n605 10.6151
R2253 B.n605 B.n72 10.6151
R2254 B.n601 B.n72 10.6151
R2255 B.n601 B.n600 10.6151
R2256 B.n600 B.n599 10.6151
R2257 B.n599 B.n74 10.6151
R2258 B.n595 B.n74 10.6151
R2259 B.n595 B.n594 10.6151
R2260 B.n594 B.n593 10.6151
R2261 B.n593 B.n76 10.6151
R2262 B.n589 B.n76 10.6151
R2263 B.n589 B.n588 10.6151
R2264 B.n588 B.n587 10.6151
R2265 B.n587 B.n78 10.6151
R2266 B.n583 B.n78 10.6151
R2267 B.n583 B.n582 10.6151
R2268 B.n582 B.n581 10.6151
R2269 B.n581 B.n80 10.6151
R2270 B.n577 B.n80 10.6151
R2271 B.n577 B.n576 10.6151
R2272 B.n576 B.n575 10.6151
R2273 B.n575 B.n82 10.6151
R2274 B.n571 B.n82 10.6151
R2275 B.n571 B.n570 10.6151
R2276 B.n569 B.n84 10.6151
R2277 B.n565 B.n84 10.6151
R2278 B.n565 B.n564 10.6151
R2279 B.n564 B.n563 10.6151
R2280 B.n563 B.n86 10.6151
R2281 B.n559 B.n86 10.6151
R2282 B.n559 B.n558 10.6151
R2283 B.n558 B.n557 10.6151
R2284 B.n557 B.n88 10.6151
R2285 B.n553 B.n88 10.6151
R2286 B.n553 B.n552 10.6151
R2287 B.n552 B.n551 10.6151
R2288 B.n551 B.n90 10.6151
R2289 B.n547 B.n90 10.6151
R2290 B.n547 B.n546 10.6151
R2291 B.n546 B.n545 10.6151
R2292 B.n545 B.n92 10.6151
R2293 B.n541 B.n92 10.6151
R2294 B.n541 B.n540 10.6151
R2295 B.n540 B.n539 10.6151
R2296 B.n539 B.n94 10.6151
R2297 B.n535 B.n94 10.6151
R2298 B.n535 B.n534 10.6151
R2299 B.n534 B.n533 10.6151
R2300 B.n533 B.n96 10.6151
R2301 B.n529 B.n96 10.6151
R2302 B.n529 B.n528 10.6151
R2303 B.n528 B.n527 10.6151
R2304 B.n527 B.n98 10.6151
R2305 B.n523 B.n98 10.6151
R2306 B.n523 B.n522 10.6151
R2307 B.n522 B.n521 10.6151
R2308 B.n521 B.n100 10.6151
R2309 B.n517 B.n100 10.6151
R2310 B.n517 B.n516 10.6151
R2311 B.n516 B.n515 10.6151
R2312 B.n515 B.n102 10.6151
R2313 B.n511 B.n102 10.6151
R2314 B.n511 B.n510 10.6151
R2315 B.n510 B.n509 10.6151
R2316 B.n509 B.n104 10.6151
R2317 B.n505 B.n104 10.6151
R2318 B.n505 B.n504 10.6151
R2319 B.n504 B.n503 10.6151
R2320 B.n503 B.n106 10.6151
R2321 B.n499 B.n106 10.6151
R2322 B.n499 B.n498 10.6151
R2323 B.n498 B.n497 10.6151
R2324 B.n497 B.n108 10.6151
R2325 B.n493 B.n108 10.6151
R2326 B.n493 B.n492 10.6151
R2327 B.n492 B.n491 10.6151
R2328 B.n491 B.n110 10.6151
R2329 B.n487 B.n110 10.6151
R2330 B.n487 B.n486 10.6151
R2331 B.n486 B.n485 10.6151
R2332 B.n485 B.n112 10.6151
R2333 B.n481 B.n112 10.6151
R2334 B.n481 B.n480 10.6151
R2335 B.n480 B.n479 10.6151
R2336 B.n479 B.n114 10.6151
R2337 B.n475 B.n114 10.6151
R2338 B.n475 B.n474 10.6151
R2339 B.n474 B.n473 10.6151
R2340 B.n473 B.n116 10.6151
R2341 B.n469 B.n116 10.6151
R2342 B.n469 B.n468 10.6151
R2343 B.n468 B.n467 10.6151
R2344 B.n467 B.n118 10.6151
R2345 B.n463 B.n118 10.6151
R2346 B.n463 B.n462 10.6151
R2347 B.n462 B.n461 10.6151
R2348 B.n461 B.n120 10.6151
R2349 B.n457 B.n120 10.6151
R2350 B.n457 B.n456 10.6151
R2351 B.n456 B.n455 10.6151
R2352 B.n455 B.n122 10.6151
R2353 B.n451 B.n122 10.6151
R2354 B.n451 B.n450 10.6151
R2355 B.n450 B.n449 10.6151
R2356 B.n449 B.n124 10.6151
R2357 B.n445 B.n124 10.6151
R2358 B.n445 B.n444 10.6151
R2359 B.n444 B.n443 10.6151
R2360 B.n443 B.n126 10.6151
R2361 B.n206 B.n1 10.6151
R2362 B.n207 B.n206 10.6151
R2363 B.n207 B.n204 10.6151
R2364 B.n211 B.n204 10.6151
R2365 B.n212 B.n211 10.6151
R2366 B.n213 B.n212 10.6151
R2367 B.n213 B.n202 10.6151
R2368 B.n217 B.n202 10.6151
R2369 B.n218 B.n217 10.6151
R2370 B.n219 B.n218 10.6151
R2371 B.n219 B.n200 10.6151
R2372 B.n223 B.n200 10.6151
R2373 B.n224 B.n223 10.6151
R2374 B.n225 B.n224 10.6151
R2375 B.n225 B.n198 10.6151
R2376 B.n229 B.n198 10.6151
R2377 B.n230 B.n229 10.6151
R2378 B.n231 B.n230 10.6151
R2379 B.n231 B.n196 10.6151
R2380 B.n235 B.n196 10.6151
R2381 B.n236 B.n235 10.6151
R2382 B.n237 B.n236 10.6151
R2383 B.n237 B.n194 10.6151
R2384 B.n241 B.n194 10.6151
R2385 B.n242 B.n241 10.6151
R2386 B.n243 B.n242 10.6151
R2387 B.n243 B.n192 10.6151
R2388 B.n247 B.n192 10.6151
R2389 B.n248 B.n247 10.6151
R2390 B.n249 B.n248 10.6151
R2391 B.n249 B.n190 10.6151
R2392 B.n253 B.n190 10.6151
R2393 B.n254 B.n253 10.6151
R2394 B.n255 B.n254 10.6151
R2395 B.n255 B.n188 10.6151
R2396 B.n259 B.n188 10.6151
R2397 B.n260 B.n259 10.6151
R2398 B.n261 B.n260 10.6151
R2399 B.n261 B.n186 10.6151
R2400 B.n265 B.n186 10.6151
R2401 B.n266 B.n265 10.6151
R2402 B.n267 B.n184 10.6151
R2403 B.n271 B.n184 10.6151
R2404 B.n272 B.n271 10.6151
R2405 B.n273 B.n272 10.6151
R2406 B.n273 B.n182 10.6151
R2407 B.n277 B.n182 10.6151
R2408 B.n278 B.n277 10.6151
R2409 B.n279 B.n278 10.6151
R2410 B.n279 B.n180 10.6151
R2411 B.n283 B.n180 10.6151
R2412 B.n284 B.n283 10.6151
R2413 B.n285 B.n284 10.6151
R2414 B.n285 B.n178 10.6151
R2415 B.n289 B.n178 10.6151
R2416 B.n290 B.n289 10.6151
R2417 B.n291 B.n290 10.6151
R2418 B.n291 B.n176 10.6151
R2419 B.n295 B.n176 10.6151
R2420 B.n296 B.n295 10.6151
R2421 B.n297 B.n296 10.6151
R2422 B.n297 B.n174 10.6151
R2423 B.n301 B.n174 10.6151
R2424 B.n302 B.n301 10.6151
R2425 B.n303 B.n302 10.6151
R2426 B.n303 B.n172 10.6151
R2427 B.n307 B.n172 10.6151
R2428 B.n308 B.n307 10.6151
R2429 B.n309 B.n308 10.6151
R2430 B.n309 B.n170 10.6151
R2431 B.n313 B.n170 10.6151
R2432 B.n314 B.n313 10.6151
R2433 B.n315 B.n314 10.6151
R2434 B.n315 B.n168 10.6151
R2435 B.n319 B.n168 10.6151
R2436 B.n320 B.n319 10.6151
R2437 B.n321 B.n320 10.6151
R2438 B.n321 B.n166 10.6151
R2439 B.n325 B.n166 10.6151
R2440 B.n326 B.n325 10.6151
R2441 B.n327 B.n326 10.6151
R2442 B.n327 B.n164 10.6151
R2443 B.n331 B.n164 10.6151
R2444 B.n332 B.n331 10.6151
R2445 B.n333 B.n332 10.6151
R2446 B.n333 B.n162 10.6151
R2447 B.n337 B.n162 10.6151
R2448 B.n338 B.n337 10.6151
R2449 B.n339 B.n338 10.6151
R2450 B.n339 B.n160 10.6151
R2451 B.n343 B.n160 10.6151
R2452 B.n344 B.n343 10.6151
R2453 B.n346 B.n156 10.6151
R2454 B.n350 B.n156 10.6151
R2455 B.n351 B.n350 10.6151
R2456 B.n352 B.n351 10.6151
R2457 B.n352 B.n154 10.6151
R2458 B.n356 B.n154 10.6151
R2459 B.n357 B.n356 10.6151
R2460 B.n361 B.n357 10.6151
R2461 B.n365 B.n152 10.6151
R2462 B.n366 B.n365 10.6151
R2463 B.n367 B.n366 10.6151
R2464 B.n367 B.n150 10.6151
R2465 B.n371 B.n150 10.6151
R2466 B.n372 B.n371 10.6151
R2467 B.n373 B.n372 10.6151
R2468 B.n373 B.n148 10.6151
R2469 B.n377 B.n148 10.6151
R2470 B.n378 B.n377 10.6151
R2471 B.n379 B.n378 10.6151
R2472 B.n379 B.n146 10.6151
R2473 B.n383 B.n146 10.6151
R2474 B.n384 B.n383 10.6151
R2475 B.n385 B.n384 10.6151
R2476 B.n385 B.n144 10.6151
R2477 B.n389 B.n144 10.6151
R2478 B.n390 B.n389 10.6151
R2479 B.n391 B.n390 10.6151
R2480 B.n391 B.n142 10.6151
R2481 B.n395 B.n142 10.6151
R2482 B.n396 B.n395 10.6151
R2483 B.n397 B.n396 10.6151
R2484 B.n397 B.n140 10.6151
R2485 B.n401 B.n140 10.6151
R2486 B.n402 B.n401 10.6151
R2487 B.n403 B.n402 10.6151
R2488 B.n403 B.n138 10.6151
R2489 B.n407 B.n138 10.6151
R2490 B.n408 B.n407 10.6151
R2491 B.n409 B.n408 10.6151
R2492 B.n409 B.n136 10.6151
R2493 B.n413 B.n136 10.6151
R2494 B.n414 B.n413 10.6151
R2495 B.n415 B.n414 10.6151
R2496 B.n415 B.n134 10.6151
R2497 B.n419 B.n134 10.6151
R2498 B.n420 B.n419 10.6151
R2499 B.n421 B.n420 10.6151
R2500 B.n421 B.n132 10.6151
R2501 B.n425 B.n132 10.6151
R2502 B.n426 B.n425 10.6151
R2503 B.n427 B.n426 10.6151
R2504 B.n427 B.n130 10.6151
R2505 B.n431 B.n130 10.6151
R2506 B.n432 B.n431 10.6151
R2507 B.n433 B.n432 10.6151
R2508 B.n433 B.n128 10.6151
R2509 B.n437 B.n128 10.6151
R2510 B.n438 B.n437 10.6151
R2511 B.n439 B.n438 10.6151
R2512 B.n805 B.n0 8.11757
R2513 B.n805 B.n1 8.11757
R2514 B.n662 B.n661 6.5566
R2515 B.n649 B.n648 6.5566
R2516 B.n346 B.n345 6.5566
R2517 B.n361 B.n360 6.5566
R2518 B.n663 B.n662 4.05904
R2519 B.n648 B.n647 4.05904
R2520 B.n345 B.n344 4.05904
R2521 B.n360 B.n152 4.05904
C0 VP VTAIL 12.1551f
C1 w_n3322_n4046# VTAIL 3.59092f
C2 VDD1 VN 0.151285f
C3 B VN 1.07634f
C4 VDD2 VN 12.0437f
C5 VDD1 VTAIL 12.745799f
C6 B VTAIL 3.97919f
C7 w_n3322_n4046# VP 7.2948f
C8 VDD2 VTAIL 12.7876f
C9 VN VTAIL 12.140599f
C10 VDD1 VP 12.348f
C11 w_n3322_n4046# VDD1 2.66216f
C12 B VP 1.79325f
C13 w_n3322_n4046# B 9.865821f
C14 VDD2 VP 0.460437f
C15 w_n3322_n4046# VDD2 2.7554f
C16 VDD1 B 2.3542f
C17 VP VN 7.59503f
C18 w_n3322_n4046# VN 6.86529f
C19 VDD1 VDD2 1.54522f
C20 VDD2 B 2.43434f
C21 VDD2 VSUBS 1.878988f
C22 VDD1 VSUBS 1.656003f
C23 VTAIL VSUBS 1.172281f
C24 VN VSUBS 6.30025f
C25 VP VSUBS 3.117728f
C26 B VSUBS 4.44977f
C27 w_n3322_n4046# VSUBS 0.164758p
C28 B.n0 VSUBS 0.007439f
C29 B.n1 VSUBS 0.007439f
C30 B.n2 VSUBS 0.011002f
C31 B.n3 VSUBS 0.008431f
C32 B.n4 VSUBS 0.008431f
C33 B.n5 VSUBS 0.008431f
C34 B.n6 VSUBS 0.008431f
C35 B.n7 VSUBS 0.008431f
C36 B.n8 VSUBS 0.008431f
C37 B.n9 VSUBS 0.008431f
C38 B.n10 VSUBS 0.008431f
C39 B.n11 VSUBS 0.008431f
C40 B.n12 VSUBS 0.008431f
C41 B.n13 VSUBS 0.008431f
C42 B.n14 VSUBS 0.008431f
C43 B.n15 VSUBS 0.008431f
C44 B.n16 VSUBS 0.008431f
C45 B.n17 VSUBS 0.008431f
C46 B.n18 VSUBS 0.008431f
C47 B.n19 VSUBS 0.008431f
C48 B.n20 VSUBS 0.008431f
C49 B.n21 VSUBS 0.008431f
C50 B.n22 VSUBS 0.008431f
C51 B.n23 VSUBS 0.02069f
C52 B.n24 VSUBS 0.008431f
C53 B.n25 VSUBS 0.008431f
C54 B.n26 VSUBS 0.008431f
C55 B.n27 VSUBS 0.008431f
C56 B.n28 VSUBS 0.008431f
C57 B.n29 VSUBS 0.008431f
C58 B.n30 VSUBS 0.008431f
C59 B.n31 VSUBS 0.008431f
C60 B.n32 VSUBS 0.008431f
C61 B.n33 VSUBS 0.008431f
C62 B.n34 VSUBS 0.008431f
C63 B.n35 VSUBS 0.008431f
C64 B.n36 VSUBS 0.008431f
C65 B.n37 VSUBS 0.008431f
C66 B.n38 VSUBS 0.008431f
C67 B.n39 VSUBS 0.008431f
C68 B.n40 VSUBS 0.008431f
C69 B.n41 VSUBS 0.008431f
C70 B.n42 VSUBS 0.008431f
C71 B.n43 VSUBS 0.008431f
C72 B.n44 VSUBS 0.008431f
C73 B.n45 VSUBS 0.008431f
C74 B.n46 VSUBS 0.008431f
C75 B.n47 VSUBS 0.008431f
C76 B.n48 VSUBS 0.008431f
C77 B.n49 VSUBS 0.008431f
C78 B.t1 VSUBS 0.347669f
C79 B.t2 VSUBS 0.374949f
C80 B.t0 VSUBS 1.3073f
C81 B.n50 VSUBS 0.54941f
C82 B.n51 VSUBS 0.352617f
C83 B.n52 VSUBS 0.008431f
C84 B.n53 VSUBS 0.008431f
C85 B.n54 VSUBS 0.008431f
C86 B.n55 VSUBS 0.008431f
C87 B.t4 VSUBS 0.347673f
C88 B.t5 VSUBS 0.374953f
C89 B.t3 VSUBS 1.3073f
C90 B.n56 VSUBS 0.549406f
C91 B.n57 VSUBS 0.352613f
C92 B.n58 VSUBS 0.008431f
C93 B.n59 VSUBS 0.008431f
C94 B.n60 VSUBS 0.008431f
C95 B.n61 VSUBS 0.008431f
C96 B.n62 VSUBS 0.008431f
C97 B.n63 VSUBS 0.008431f
C98 B.n64 VSUBS 0.008431f
C99 B.n65 VSUBS 0.008431f
C100 B.n66 VSUBS 0.008431f
C101 B.n67 VSUBS 0.008431f
C102 B.n68 VSUBS 0.008431f
C103 B.n69 VSUBS 0.008431f
C104 B.n70 VSUBS 0.008431f
C105 B.n71 VSUBS 0.008431f
C106 B.n72 VSUBS 0.008431f
C107 B.n73 VSUBS 0.008431f
C108 B.n74 VSUBS 0.008431f
C109 B.n75 VSUBS 0.008431f
C110 B.n76 VSUBS 0.008431f
C111 B.n77 VSUBS 0.008431f
C112 B.n78 VSUBS 0.008431f
C113 B.n79 VSUBS 0.008431f
C114 B.n80 VSUBS 0.008431f
C115 B.n81 VSUBS 0.008431f
C116 B.n82 VSUBS 0.008431f
C117 B.n83 VSUBS 0.02069f
C118 B.n84 VSUBS 0.008431f
C119 B.n85 VSUBS 0.008431f
C120 B.n86 VSUBS 0.008431f
C121 B.n87 VSUBS 0.008431f
C122 B.n88 VSUBS 0.008431f
C123 B.n89 VSUBS 0.008431f
C124 B.n90 VSUBS 0.008431f
C125 B.n91 VSUBS 0.008431f
C126 B.n92 VSUBS 0.008431f
C127 B.n93 VSUBS 0.008431f
C128 B.n94 VSUBS 0.008431f
C129 B.n95 VSUBS 0.008431f
C130 B.n96 VSUBS 0.008431f
C131 B.n97 VSUBS 0.008431f
C132 B.n98 VSUBS 0.008431f
C133 B.n99 VSUBS 0.008431f
C134 B.n100 VSUBS 0.008431f
C135 B.n101 VSUBS 0.008431f
C136 B.n102 VSUBS 0.008431f
C137 B.n103 VSUBS 0.008431f
C138 B.n104 VSUBS 0.008431f
C139 B.n105 VSUBS 0.008431f
C140 B.n106 VSUBS 0.008431f
C141 B.n107 VSUBS 0.008431f
C142 B.n108 VSUBS 0.008431f
C143 B.n109 VSUBS 0.008431f
C144 B.n110 VSUBS 0.008431f
C145 B.n111 VSUBS 0.008431f
C146 B.n112 VSUBS 0.008431f
C147 B.n113 VSUBS 0.008431f
C148 B.n114 VSUBS 0.008431f
C149 B.n115 VSUBS 0.008431f
C150 B.n116 VSUBS 0.008431f
C151 B.n117 VSUBS 0.008431f
C152 B.n118 VSUBS 0.008431f
C153 B.n119 VSUBS 0.008431f
C154 B.n120 VSUBS 0.008431f
C155 B.n121 VSUBS 0.008431f
C156 B.n122 VSUBS 0.008431f
C157 B.n123 VSUBS 0.008431f
C158 B.n124 VSUBS 0.008431f
C159 B.n125 VSUBS 0.008431f
C160 B.n126 VSUBS 0.020213f
C161 B.n127 VSUBS 0.008431f
C162 B.n128 VSUBS 0.008431f
C163 B.n129 VSUBS 0.008431f
C164 B.n130 VSUBS 0.008431f
C165 B.n131 VSUBS 0.008431f
C166 B.n132 VSUBS 0.008431f
C167 B.n133 VSUBS 0.008431f
C168 B.n134 VSUBS 0.008431f
C169 B.n135 VSUBS 0.008431f
C170 B.n136 VSUBS 0.008431f
C171 B.n137 VSUBS 0.008431f
C172 B.n138 VSUBS 0.008431f
C173 B.n139 VSUBS 0.008431f
C174 B.n140 VSUBS 0.008431f
C175 B.n141 VSUBS 0.008431f
C176 B.n142 VSUBS 0.008431f
C177 B.n143 VSUBS 0.008431f
C178 B.n144 VSUBS 0.008431f
C179 B.n145 VSUBS 0.008431f
C180 B.n146 VSUBS 0.008431f
C181 B.n147 VSUBS 0.008431f
C182 B.n148 VSUBS 0.008431f
C183 B.n149 VSUBS 0.008431f
C184 B.n150 VSUBS 0.008431f
C185 B.n151 VSUBS 0.008431f
C186 B.n152 VSUBS 0.005828f
C187 B.n153 VSUBS 0.008431f
C188 B.n154 VSUBS 0.008431f
C189 B.n155 VSUBS 0.008431f
C190 B.n156 VSUBS 0.008431f
C191 B.n157 VSUBS 0.008431f
C192 B.t8 VSUBS 0.347669f
C193 B.t7 VSUBS 0.374949f
C194 B.t6 VSUBS 1.3073f
C195 B.n158 VSUBS 0.54941f
C196 B.n159 VSUBS 0.352617f
C197 B.n160 VSUBS 0.008431f
C198 B.n161 VSUBS 0.008431f
C199 B.n162 VSUBS 0.008431f
C200 B.n163 VSUBS 0.008431f
C201 B.n164 VSUBS 0.008431f
C202 B.n165 VSUBS 0.008431f
C203 B.n166 VSUBS 0.008431f
C204 B.n167 VSUBS 0.008431f
C205 B.n168 VSUBS 0.008431f
C206 B.n169 VSUBS 0.008431f
C207 B.n170 VSUBS 0.008431f
C208 B.n171 VSUBS 0.008431f
C209 B.n172 VSUBS 0.008431f
C210 B.n173 VSUBS 0.008431f
C211 B.n174 VSUBS 0.008431f
C212 B.n175 VSUBS 0.008431f
C213 B.n176 VSUBS 0.008431f
C214 B.n177 VSUBS 0.008431f
C215 B.n178 VSUBS 0.008431f
C216 B.n179 VSUBS 0.008431f
C217 B.n180 VSUBS 0.008431f
C218 B.n181 VSUBS 0.008431f
C219 B.n182 VSUBS 0.008431f
C220 B.n183 VSUBS 0.008431f
C221 B.n184 VSUBS 0.008431f
C222 B.n185 VSUBS 0.019234f
C223 B.n186 VSUBS 0.008431f
C224 B.n187 VSUBS 0.008431f
C225 B.n188 VSUBS 0.008431f
C226 B.n189 VSUBS 0.008431f
C227 B.n190 VSUBS 0.008431f
C228 B.n191 VSUBS 0.008431f
C229 B.n192 VSUBS 0.008431f
C230 B.n193 VSUBS 0.008431f
C231 B.n194 VSUBS 0.008431f
C232 B.n195 VSUBS 0.008431f
C233 B.n196 VSUBS 0.008431f
C234 B.n197 VSUBS 0.008431f
C235 B.n198 VSUBS 0.008431f
C236 B.n199 VSUBS 0.008431f
C237 B.n200 VSUBS 0.008431f
C238 B.n201 VSUBS 0.008431f
C239 B.n202 VSUBS 0.008431f
C240 B.n203 VSUBS 0.008431f
C241 B.n204 VSUBS 0.008431f
C242 B.n205 VSUBS 0.008431f
C243 B.n206 VSUBS 0.008431f
C244 B.n207 VSUBS 0.008431f
C245 B.n208 VSUBS 0.008431f
C246 B.n209 VSUBS 0.008431f
C247 B.n210 VSUBS 0.008431f
C248 B.n211 VSUBS 0.008431f
C249 B.n212 VSUBS 0.008431f
C250 B.n213 VSUBS 0.008431f
C251 B.n214 VSUBS 0.008431f
C252 B.n215 VSUBS 0.008431f
C253 B.n216 VSUBS 0.008431f
C254 B.n217 VSUBS 0.008431f
C255 B.n218 VSUBS 0.008431f
C256 B.n219 VSUBS 0.008431f
C257 B.n220 VSUBS 0.008431f
C258 B.n221 VSUBS 0.008431f
C259 B.n222 VSUBS 0.008431f
C260 B.n223 VSUBS 0.008431f
C261 B.n224 VSUBS 0.008431f
C262 B.n225 VSUBS 0.008431f
C263 B.n226 VSUBS 0.008431f
C264 B.n227 VSUBS 0.008431f
C265 B.n228 VSUBS 0.008431f
C266 B.n229 VSUBS 0.008431f
C267 B.n230 VSUBS 0.008431f
C268 B.n231 VSUBS 0.008431f
C269 B.n232 VSUBS 0.008431f
C270 B.n233 VSUBS 0.008431f
C271 B.n234 VSUBS 0.008431f
C272 B.n235 VSUBS 0.008431f
C273 B.n236 VSUBS 0.008431f
C274 B.n237 VSUBS 0.008431f
C275 B.n238 VSUBS 0.008431f
C276 B.n239 VSUBS 0.008431f
C277 B.n240 VSUBS 0.008431f
C278 B.n241 VSUBS 0.008431f
C279 B.n242 VSUBS 0.008431f
C280 B.n243 VSUBS 0.008431f
C281 B.n244 VSUBS 0.008431f
C282 B.n245 VSUBS 0.008431f
C283 B.n246 VSUBS 0.008431f
C284 B.n247 VSUBS 0.008431f
C285 B.n248 VSUBS 0.008431f
C286 B.n249 VSUBS 0.008431f
C287 B.n250 VSUBS 0.008431f
C288 B.n251 VSUBS 0.008431f
C289 B.n252 VSUBS 0.008431f
C290 B.n253 VSUBS 0.008431f
C291 B.n254 VSUBS 0.008431f
C292 B.n255 VSUBS 0.008431f
C293 B.n256 VSUBS 0.008431f
C294 B.n257 VSUBS 0.008431f
C295 B.n258 VSUBS 0.008431f
C296 B.n259 VSUBS 0.008431f
C297 B.n260 VSUBS 0.008431f
C298 B.n261 VSUBS 0.008431f
C299 B.n262 VSUBS 0.008431f
C300 B.n263 VSUBS 0.008431f
C301 B.n264 VSUBS 0.008431f
C302 B.n265 VSUBS 0.008431f
C303 B.n266 VSUBS 0.019234f
C304 B.n267 VSUBS 0.02069f
C305 B.n268 VSUBS 0.02069f
C306 B.n269 VSUBS 0.008431f
C307 B.n270 VSUBS 0.008431f
C308 B.n271 VSUBS 0.008431f
C309 B.n272 VSUBS 0.008431f
C310 B.n273 VSUBS 0.008431f
C311 B.n274 VSUBS 0.008431f
C312 B.n275 VSUBS 0.008431f
C313 B.n276 VSUBS 0.008431f
C314 B.n277 VSUBS 0.008431f
C315 B.n278 VSUBS 0.008431f
C316 B.n279 VSUBS 0.008431f
C317 B.n280 VSUBS 0.008431f
C318 B.n281 VSUBS 0.008431f
C319 B.n282 VSUBS 0.008431f
C320 B.n283 VSUBS 0.008431f
C321 B.n284 VSUBS 0.008431f
C322 B.n285 VSUBS 0.008431f
C323 B.n286 VSUBS 0.008431f
C324 B.n287 VSUBS 0.008431f
C325 B.n288 VSUBS 0.008431f
C326 B.n289 VSUBS 0.008431f
C327 B.n290 VSUBS 0.008431f
C328 B.n291 VSUBS 0.008431f
C329 B.n292 VSUBS 0.008431f
C330 B.n293 VSUBS 0.008431f
C331 B.n294 VSUBS 0.008431f
C332 B.n295 VSUBS 0.008431f
C333 B.n296 VSUBS 0.008431f
C334 B.n297 VSUBS 0.008431f
C335 B.n298 VSUBS 0.008431f
C336 B.n299 VSUBS 0.008431f
C337 B.n300 VSUBS 0.008431f
C338 B.n301 VSUBS 0.008431f
C339 B.n302 VSUBS 0.008431f
C340 B.n303 VSUBS 0.008431f
C341 B.n304 VSUBS 0.008431f
C342 B.n305 VSUBS 0.008431f
C343 B.n306 VSUBS 0.008431f
C344 B.n307 VSUBS 0.008431f
C345 B.n308 VSUBS 0.008431f
C346 B.n309 VSUBS 0.008431f
C347 B.n310 VSUBS 0.008431f
C348 B.n311 VSUBS 0.008431f
C349 B.n312 VSUBS 0.008431f
C350 B.n313 VSUBS 0.008431f
C351 B.n314 VSUBS 0.008431f
C352 B.n315 VSUBS 0.008431f
C353 B.n316 VSUBS 0.008431f
C354 B.n317 VSUBS 0.008431f
C355 B.n318 VSUBS 0.008431f
C356 B.n319 VSUBS 0.008431f
C357 B.n320 VSUBS 0.008431f
C358 B.n321 VSUBS 0.008431f
C359 B.n322 VSUBS 0.008431f
C360 B.n323 VSUBS 0.008431f
C361 B.n324 VSUBS 0.008431f
C362 B.n325 VSUBS 0.008431f
C363 B.n326 VSUBS 0.008431f
C364 B.n327 VSUBS 0.008431f
C365 B.n328 VSUBS 0.008431f
C366 B.n329 VSUBS 0.008431f
C367 B.n330 VSUBS 0.008431f
C368 B.n331 VSUBS 0.008431f
C369 B.n332 VSUBS 0.008431f
C370 B.n333 VSUBS 0.008431f
C371 B.n334 VSUBS 0.008431f
C372 B.n335 VSUBS 0.008431f
C373 B.n336 VSUBS 0.008431f
C374 B.n337 VSUBS 0.008431f
C375 B.n338 VSUBS 0.008431f
C376 B.n339 VSUBS 0.008431f
C377 B.n340 VSUBS 0.008431f
C378 B.n341 VSUBS 0.008431f
C379 B.n342 VSUBS 0.008431f
C380 B.n343 VSUBS 0.008431f
C381 B.n344 VSUBS 0.005828f
C382 B.n345 VSUBS 0.019534f
C383 B.n346 VSUBS 0.006819f
C384 B.n347 VSUBS 0.008431f
C385 B.n348 VSUBS 0.008431f
C386 B.n349 VSUBS 0.008431f
C387 B.n350 VSUBS 0.008431f
C388 B.n351 VSUBS 0.008431f
C389 B.n352 VSUBS 0.008431f
C390 B.n353 VSUBS 0.008431f
C391 B.n354 VSUBS 0.008431f
C392 B.n355 VSUBS 0.008431f
C393 B.n356 VSUBS 0.008431f
C394 B.n357 VSUBS 0.008431f
C395 B.t11 VSUBS 0.347673f
C396 B.t10 VSUBS 0.374953f
C397 B.t9 VSUBS 1.3073f
C398 B.n358 VSUBS 0.549406f
C399 B.n359 VSUBS 0.352613f
C400 B.n360 VSUBS 0.019534f
C401 B.n361 VSUBS 0.006819f
C402 B.n362 VSUBS 0.008431f
C403 B.n363 VSUBS 0.008431f
C404 B.n364 VSUBS 0.008431f
C405 B.n365 VSUBS 0.008431f
C406 B.n366 VSUBS 0.008431f
C407 B.n367 VSUBS 0.008431f
C408 B.n368 VSUBS 0.008431f
C409 B.n369 VSUBS 0.008431f
C410 B.n370 VSUBS 0.008431f
C411 B.n371 VSUBS 0.008431f
C412 B.n372 VSUBS 0.008431f
C413 B.n373 VSUBS 0.008431f
C414 B.n374 VSUBS 0.008431f
C415 B.n375 VSUBS 0.008431f
C416 B.n376 VSUBS 0.008431f
C417 B.n377 VSUBS 0.008431f
C418 B.n378 VSUBS 0.008431f
C419 B.n379 VSUBS 0.008431f
C420 B.n380 VSUBS 0.008431f
C421 B.n381 VSUBS 0.008431f
C422 B.n382 VSUBS 0.008431f
C423 B.n383 VSUBS 0.008431f
C424 B.n384 VSUBS 0.008431f
C425 B.n385 VSUBS 0.008431f
C426 B.n386 VSUBS 0.008431f
C427 B.n387 VSUBS 0.008431f
C428 B.n388 VSUBS 0.008431f
C429 B.n389 VSUBS 0.008431f
C430 B.n390 VSUBS 0.008431f
C431 B.n391 VSUBS 0.008431f
C432 B.n392 VSUBS 0.008431f
C433 B.n393 VSUBS 0.008431f
C434 B.n394 VSUBS 0.008431f
C435 B.n395 VSUBS 0.008431f
C436 B.n396 VSUBS 0.008431f
C437 B.n397 VSUBS 0.008431f
C438 B.n398 VSUBS 0.008431f
C439 B.n399 VSUBS 0.008431f
C440 B.n400 VSUBS 0.008431f
C441 B.n401 VSUBS 0.008431f
C442 B.n402 VSUBS 0.008431f
C443 B.n403 VSUBS 0.008431f
C444 B.n404 VSUBS 0.008431f
C445 B.n405 VSUBS 0.008431f
C446 B.n406 VSUBS 0.008431f
C447 B.n407 VSUBS 0.008431f
C448 B.n408 VSUBS 0.008431f
C449 B.n409 VSUBS 0.008431f
C450 B.n410 VSUBS 0.008431f
C451 B.n411 VSUBS 0.008431f
C452 B.n412 VSUBS 0.008431f
C453 B.n413 VSUBS 0.008431f
C454 B.n414 VSUBS 0.008431f
C455 B.n415 VSUBS 0.008431f
C456 B.n416 VSUBS 0.008431f
C457 B.n417 VSUBS 0.008431f
C458 B.n418 VSUBS 0.008431f
C459 B.n419 VSUBS 0.008431f
C460 B.n420 VSUBS 0.008431f
C461 B.n421 VSUBS 0.008431f
C462 B.n422 VSUBS 0.008431f
C463 B.n423 VSUBS 0.008431f
C464 B.n424 VSUBS 0.008431f
C465 B.n425 VSUBS 0.008431f
C466 B.n426 VSUBS 0.008431f
C467 B.n427 VSUBS 0.008431f
C468 B.n428 VSUBS 0.008431f
C469 B.n429 VSUBS 0.008431f
C470 B.n430 VSUBS 0.008431f
C471 B.n431 VSUBS 0.008431f
C472 B.n432 VSUBS 0.008431f
C473 B.n433 VSUBS 0.008431f
C474 B.n434 VSUBS 0.008431f
C475 B.n435 VSUBS 0.008431f
C476 B.n436 VSUBS 0.008431f
C477 B.n437 VSUBS 0.008431f
C478 B.n438 VSUBS 0.008431f
C479 B.n439 VSUBS 0.019712f
C480 B.n440 VSUBS 0.02069f
C481 B.n441 VSUBS 0.019234f
C482 B.n442 VSUBS 0.008431f
C483 B.n443 VSUBS 0.008431f
C484 B.n444 VSUBS 0.008431f
C485 B.n445 VSUBS 0.008431f
C486 B.n446 VSUBS 0.008431f
C487 B.n447 VSUBS 0.008431f
C488 B.n448 VSUBS 0.008431f
C489 B.n449 VSUBS 0.008431f
C490 B.n450 VSUBS 0.008431f
C491 B.n451 VSUBS 0.008431f
C492 B.n452 VSUBS 0.008431f
C493 B.n453 VSUBS 0.008431f
C494 B.n454 VSUBS 0.008431f
C495 B.n455 VSUBS 0.008431f
C496 B.n456 VSUBS 0.008431f
C497 B.n457 VSUBS 0.008431f
C498 B.n458 VSUBS 0.008431f
C499 B.n459 VSUBS 0.008431f
C500 B.n460 VSUBS 0.008431f
C501 B.n461 VSUBS 0.008431f
C502 B.n462 VSUBS 0.008431f
C503 B.n463 VSUBS 0.008431f
C504 B.n464 VSUBS 0.008431f
C505 B.n465 VSUBS 0.008431f
C506 B.n466 VSUBS 0.008431f
C507 B.n467 VSUBS 0.008431f
C508 B.n468 VSUBS 0.008431f
C509 B.n469 VSUBS 0.008431f
C510 B.n470 VSUBS 0.008431f
C511 B.n471 VSUBS 0.008431f
C512 B.n472 VSUBS 0.008431f
C513 B.n473 VSUBS 0.008431f
C514 B.n474 VSUBS 0.008431f
C515 B.n475 VSUBS 0.008431f
C516 B.n476 VSUBS 0.008431f
C517 B.n477 VSUBS 0.008431f
C518 B.n478 VSUBS 0.008431f
C519 B.n479 VSUBS 0.008431f
C520 B.n480 VSUBS 0.008431f
C521 B.n481 VSUBS 0.008431f
C522 B.n482 VSUBS 0.008431f
C523 B.n483 VSUBS 0.008431f
C524 B.n484 VSUBS 0.008431f
C525 B.n485 VSUBS 0.008431f
C526 B.n486 VSUBS 0.008431f
C527 B.n487 VSUBS 0.008431f
C528 B.n488 VSUBS 0.008431f
C529 B.n489 VSUBS 0.008431f
C530 B.n490 VSUBS 0.008431f
C531 B.n491 VSUBS 0.008431f
C532 B.n492 VSUBS 0.008431f
C533 B.n493 VSUBS 0.008431f
C534 B.n494 VSUBS 0.008431f
C535 B.n495 VSUBS 0.008431f
C536 B.n496 VSUBS 0.008431f
C537 B.n497 VSUBS 0.008431f
C538 B.n498 VSUBS 0.008431f
C539 B.n499 VSUBS 0.008431f
C540 B.n500 VSUBS 0.008431f
C541 B.n501 VSUBS 0.008431f
C542 B.n502 VSUBS 0.008431f
C543 B.n503 VSUBS 0.008431f
C544 B.n504 VSUBS 0.008431f
C545 B.n505 VSUBS 0.008431f
C546 B.n506 VSUBS 0.008431f
C547 B.n507 VSUBS 0.008431f
C548 B.n508 VSUBS 0.008431f
C549 B.n509 VSUBS 0.008431f
C550 B.n510 VSUBS 0.008431f
C551 B.n511 VSUBS 0.008431f
C552 B.n512 VSUBS 0.008431f
C553 B.n513 VSUBS 0.008431f
C554 B.n514 VSUBS 0.008431f
C555 B.n515 VSUBS 0.008431f
C556 B.n516 VSUBS 0.008431f
C557 B.n517 VSUBS 0.008431f
C558 B.n518 VSUBS 0.008431f
C559 B.n519 VSUBS 0.008431f
C560 B.n520 VSUBS 0.008431f
C561 B.n521 VSUBS 0.008431f
C562 B.n522 VSUBS 0.008431f
C563 B.n523 VSUBS 0.008431f
C564 B.n524 VSUBS 0.008431f
C565 B.n525 VSUBS 0.008431f
C566 B.n526 VSUBS 0.008431f
C567 B.n527 VSUBS 0.008431f
C568 B.n528 VSUBS 0.008431f
C569 B.n529 VSUBS 0.008431f
C570 B.n530 VSUBS 0.008431f
C571 B.n531 VSUBS 0.008431f
C572 B.n532 VSUBS 0.008431f
C573 B.n533 VSUBS 0.008431f
C574 B.n534 VSUBS 0.008431f
C575 B.n535 VSUBS 0.008431f
C576 B.n536 VSUBS 0.008431f
C577 B.n537 VSUBS 0.008431f
C578 B.n538 VSUBS 0.008431f
C579 B.n539 VSUBS 0.008431f
C580 B.n540 VSUBS 0.008431f
C581 B.n541 VSUBS 0.008431f
C582 B.n542 VSUBS 0.008431f
C583 B.n543 VSUBS 0.008431f
C584 B.n544 VSUBS 0.008431f
C585 B.n545 VSUBS 0.008431f
C586 B.n546 VSUBS 0.008431f
C587 B.n547 VSUBS 0.008431f
C588 B.n548 VSUBS 0.008431f
C589 B.n549 VSUBS 0.008431f
C590 B.n550 VSUBS 0.008431f
C591 B.n551 VSUBS 0.008431f
C592 B.n552 VSUBS 0.008431f
C593 B.n553 VSUBS 0.008431f
C594 B.n554 VSUBS 0.008431f
C595 B.n555 VSUBS 0.008431f
C596 B.n556 VSUBS 0.008431f
C597 B.n557 VSUBS 0.008431f
C598 B.n558 VSUBS 0.008431f
C599 B.n559 VSUBS 0.008431f
C600 B.n560 VSUBS 0.008431f
C601 B.n561 VSUBS 0.008431f
C602 B.n562 VSUBS 0.008431f
C603 B.n563 VSUBS 0.008431f
C604 B.n564 VSUBS 0.008431f
C605 B.n565 VSUBS 0.008431f
C606 B.n566 VSUBS 0.008431f
C607 B.n567 VSUBS 0.008431f
C608 B.n568 VSUBS 0.019234f
C609 B.n569 VSUBS 0.019234f
C610 B.n570 VSUBS 0.02069f
C611 B.n571 VSUBS 0.008431f
C612 B.n572 VSUBS 0.008431f
C613 B.n573 VSUBS 0.008431f
C614 B.n574 VSUBS 0.008431f
C615 B.n575 VSUBS 0.008431f
C616 B.n576 VSUBS 0.008431f
C617 B.n577 VSUBS 0.008431f
C618 B.n578 VSUBS 0.008431f
C619 B.n579 VSUBS 0.008431f
C620 B.n580 VSUBS 0.008431f
C621 B.n581 VSUBS 0.008431f
C622 B.n582 VSUBS 0.008431f
C623 B.n583 VSUBS 0.008431f
C624 B.n584 VSUBS 0.008431f
C625 B.n585 VSUBS 0.008431f
C626 B.n586 VSUBS 0.008431f
C627 B.n587 VSUBS 0.008431f
C628 B.n588 VSUBS 0.008431f
C629 B.n589 VSUBS 0.008431f
C630 B.n590 VSUBS 0.008431f
C631 B.n591 VSUBS 0.008431f
C632 B.n592 VSUBS 0.008431f
C633 B.n593 VSUBS 0.008431f
C634 B.n594 VSUBS 0.008431f
C635 B.n595 VSUBS 0.008431f
C636 B.n596 VSUBS 0.008431f
C637 B.n597 VSUBS 0.008431f
C638 B.n598 VSUBS 0.008431f
C639 B.n599 VSUBS 0.008431f
C640 B.n600 VSUBS 0.008431f
C641 B.n601 VSUBS 0.008431f
C642 B.n602 VSUBS 0.008431f
C643 B.n603 VSUBS 0.008431f
C644 B.n604 VSUBS 0.008431f
C645 B.n605 VSUBS 0.008431f
C646 B.n606 VSUBS 0.008431f
C647 B.n607 VSUBS 0.008431f
C648 B.n608 VSUBS 0.008431f
C649 B.n609 VSUBS 0.008431f
C650 B.n610 VSUBS 0.008431f
C651 B.n611 VSUBS 0.008431f
C652 B.n612 VSUBS 0.008431f
C653 B.n613 VSUBS 0.008431f
C654 B.n614 VSUBS 0.008431f
C655 B.n615 VSUBS 0.008431f
C656 B.n616 VSUBS 0.008431f
C657 B.n617 VSUBS 0.008431f
C658 B.n618 VSUBS 0.008431f
C659 B.n619 VSUBS 0.008431f
C660 B.n620 VSUBS 0.008431f
C661 B.n621 VSUBS 0.008431f
C662 B.n622 VSUBS 0.008431f
C663 B.n623 VSUBS 0.008431f
C664 B.n624 VSUBS 0.008431f
C665 B.n625 VSUBS 0.008431f
C666 B.n626 VSUBS 0.008431f
C667 B.n627 VSUBS 0.008431f
C668 B.n628 VSUBS 0.008431f
C669 B.n629 VSUBS 0.008431f
C670 B.n630 VSUBS 0.008431f
C671 B.n631 VSUBS 0.008431f
C672 B.n632 VSUBS 0.008431f
C673 B.n633 VSUBS 0.008431f
C674 B.n634 VSUBS 0.008431f
C675 B.n635 VSUBS 0.008431f
C676 B.n636 VSUBS 0.008431f
C677 B.n637 VSUBS 0.008431f
C678 B.n638 VSUBS 0.008431f
C679 B.n639 VSUBS 0.008431f
C680 B.n640 VSUBS 0.008431f
C681 B.n641 VSUBS 0.008431f
C682 B.n642 VSUBS 0.008431f
C683 B.n643 VSUBS 0.008431f
C684 B.n644 VSUBS 0.008431f
C685 B.n645 VSUBS 0.008431f
C686 B.n646 VSUBS 0.008431f
C687 B.n647 VSUBS 0.005828f
C688 B.n648 VSUBS 0.019534f
C689 B.n649 VSUBS 0.006819f
C690 B.n650 VSUBS 0.008431f
C691 B.n651 VSUBS 0.008431f
C692 B.n652 VSUBS 0.008431f
C693 B.n653 VSUBS 0.008431f
C694 B.n654 VSUBS 0.008431f
C695 B.n655 VSUBS 0.008431f
C696 B.n656 VSUBS 0.008431f
C697 B.n657 VSUBS 0.008431f
C698 B.n658 VSUBS 0.008431f
C699 B.n659 VSUBS 0.008431f
C700 B.n660 VSUBS 0.008431f
C701 B.n661 VSUBS 0.006819f
C702 B.n662 VSUBS 0.019534f
C703 B.n663 VSUBS 0.005828f
C704 B.n664 VSUBS 0.008431f
C705 B.n665 VSUBS 0.008431f
C706 B.n666 VSUBS 0.008431f
C707 B.n667 VSUBS 0.008431f
C708 B.n668 VSUBS 0.008431f
C709 B.n669 VSUBS 0.008431f
C710 B.n670 VSUBS 0.008431f
C711 B.n671 VSUBS 0.008431f
C712 B.n672 VSUBS 0.008431f
C713 B.n673 VSUBS 0.008431f
C714 B.n674 VSUBS 0.008431f
C715 B.n675 VSUBS 0.008431f
C716 B.n676 VSUBS 0.008431f
C717 B.n677 VSUBS 0.008431f
C718 B.n678 VSUBS 0.008431f
C719 B.n679 VSUBS 0.008431f
C720 B.n680 VSUBS 0.008431f
C721 B.n681 VSUBS 0.008431f
C722 B.n682 VSUBS 0.008431f
C723 B.n683 VSUBS 0.008431f
C724 B.n684 VSUBS 0.008431f
C725 B.n685 VSUBS 0.008431f
C726 B.n686 VSUBS 0.008431f
C727 B.n687 VSUBS 0.008431f
C728 B.n688 VSUBS 0.008431f
C729 B.n689 VSUBS 0.008431f
C730 B.n690 VSUBS 0.008431f
C731 B.n691 VSUBS 0.008431f
C732 B.n692 VSUBS 0.008431f
C733 B.n693 VSUBS 0.008431f
C734 B.n694 VSUBS 0.008431f
C735 B.n695 VSUBS 0.008431f
C736 B.n696 VSUBS 0.008431f
C737 B.n697 VSUBS 0.008431f
C738 B.n698 VSUBS 0.008431f
C739 B.n699 VSUBS 0.008431f
C740 B.n700 VSUBS 0.008431f
C741 B.n701 VSUBS 0.008431f
C742 B.n702 VSUBS 0.008431f
C743 B.n703 VSUBS 0.008431f
C744 B.n704 VSUBS 0.008431f
C745 B.n705 VSUBS 0.008431f
C746 B.n706 VSUBS 0.008431f
C747 B.n707 VSUBS 0.008431f
C748 B.n708 VSUBS 0.008431f
C749 B.n709 VSUBS 0.008431f
C750 B.n710 VSUBS 0.008431f
C751 B.n711 VSUBS 0.008431f
C752 B.n712 VSUBS 0.008431f
C753 B.n713 VSUBS 0.008431f
C754 B.n714 VSUBS 0.008431f
C755 B.n715 VSUBS 0.008431f
C756 B.n716 VSUBS 0.008431f
C757 B.n717 VSUBS 0.008431f
C758 B.n718 VSUBS 0.008431f
C759 B.n719 VSUBS 0.008431f
C760 B.n720 VSUBS 0.008431f
C761 B.n721 VSUBS 0.008431f
C762 B.n722 VSUBS 0.008431f
C763 B.n723 VSUBS 0.008431f
C764 B.n724 VSUBS 0.008431f
C765 B.n725 VSUBS 0.008431f
C766 B.n726 VSUBS 0.008431f
C767 B.n727 VSUBS 0.008431f
C768 B.n728 VSUBS 0.008431f
C769 B.n729 VSUBS 0.008431f
C770 B.n730 VSUBS 0.008431f
C771 B.n731 VSUBS 0.008431f
C772 B.n732 VSUBS 0.008431f
C773 B.n733 VSUBS 0.008431f
C774 B.n734 VSUBS 0.008431f
C775 B.n735 VSUBS 0.008431f
C776 B.n736 VSUBS 0.008431f
C777 B.n737 VSUBS 0.008431f
C778 B.n738 VSUBS 0.008431f
C779 B.n739 VSUBS 0.008431f
C780 B.n740 VSUBS 0.02069f
C781 B.n741 VSUBS 0.019234f
C782 B.n742 VSUBS 0.019234f
C783 B.n743 VSUBS 0.008431f
C784 B.n744 VSUBS 0.008431f
C785 B.n745 VSUBS 0.008431f
C786 B.n746 VSUBS 0.008431f
C787 B.n747 VSUBS 0.008431f
C788 B.n748 VSUBS 0.008431f
C789 B.n749 VSUBS 0.008431f
C790 B.n750 VSUBS 0.008431f
C791 B.n751 VSUBS 0.008431f
C792 B.n752 VSUBS 0.008431f
C793 B.n753 VSUBS 0.008431f
C794 B.n754 VSUBS 0.008431f
C795 B.n755 VSUBS 0.008431f
C796 B.n756 VSUBS 0.008431f
C797 B.n757 VSUBS 0.008431f
C798 B.n758 VSUBS 0.008431f
C799 B.n759 VSUBS 0.008431f
C800 B.n760 VSUBS 0.008431f
C801 B.n761 VSUBS 0.008431f
C802 B.n762 VSUBS 0.008431f
C803 B.n763 VSUBS 0.008431f
C804 B.n764 VSUBS 0.008431f
C805 B.n765 VSUBS 0.008431f
C806 B.n766 VSUBS 0.008431f
C807 B.n767 VSUBS 0.008431f
C808 B.n768 VSUBS 0.008431f
C809 B.n769 VSUBS 0.008431f
C810 B.n770 VSUBS 0.008431f
C811 B.n771 VSUBS 0.008431f
C812 B.n772 VSUBS 0.008431f
C813 B.n773 VSUBS 0.008431f
C814 B.n774 VSUBS 0.008431f
C815 B.n775 VSUBS 0.008431f
C816 B.n776 VSUBS 0.008431f
C817 B.n777 VSUBS 0.008431f
C818 B.n778 VSUBS 0.008431f
C819 B.n779 VSUBS 0.008431f
C820 B.n780 VSUBS 0.008431f
C821 B.n781 VSUBS 0.008431f
C822 B.n782 VSUBS 0.008431f
C823 B.n783 VSUBS 0.008431f
C824 B.n784 VSUBS 0.008431f
C825 B.n785 VSUBS 0.008431f
C826 B.n786 VSUBS 0.008431f
C827 B.n787 VSUBS 0.008431f
C828 B.n788 VSUBS 0.008431f
C829 B.n789 VSUBS 0.008431f
C830 B.n790 VSUBS 0.008431f
C831 B.n791 VSUBS 0.008431f
C832 B.n792 VSUBS 0.008431f
C833 B.n793 VSUBS 0.008431f
C834 B.n794 VSUBS 0.008431f
C835 B.n795 VSUBS 0.008431f
C836 B.n796 VSUBS 0.008431f
C837 B.n797 VSUBS 0.008431f
C838 B.n798 VSUBS 0.008431f
C839 B.n799 VSUBS 0.008431f
C840 B.n800 VSUBS 0.008431f
C841 B.n801 VSUBS 0.008431f
C842 B.n802 VSUBS 0.008431f
C843 B.n803 VSUBS 0.011002f
C844 B.n804 VSUBS 0.01172f
C845 B.n805 VSUBS 0.023307f
C846 VDD2.n0 VSUBS 0.028f
C847 VDD2.n1 VSUBS 0.026936f
C848 VDD2.n2 VSUBS 0.014474f
C849 VDD2.n3 VSUBS 0.034211f
C850 VDD2.n4 VSUBS 0.0149f
C851 VDD2.n5 VSUBS 0.026936f
C852 VDD2.n6 VSUBS 0.015325f
C853 VDD2.n7 VSUBS 0.034211f
C854 VDD2.n8 VSUBS 0.015325f
C855 VDD2.n9 VSUBS 0.026936f
C856 VDD2.n10 VSUBS 0.014474f
C857 VDD2.n11 VSUBS 0.034211f
C858 VDD2.n12 VSUBS 0.015325f
C859 VDD2.n13 VSUBS 0.026936f
C860 VDD2.n14 VSUBS 0.014474f
C861 VDD2.n15 VSUBS 0.034211f
C862 VDD2.n16 VSUBS 0.015325f
C863 VDD2.n17 VSUBS 0.026936f
C864 VDD2.n18 VSUBS 0.014474f
C865 VDD2.n19 VSUBS 0.034211f
C866 VDD2.n20 VSUBS 0.015325f
C867 VDD2.n21 VSUBS 0.026936f
C868 VDD2.n22 VSUBS 0.014474f
C869 VDD2.n23 VSUBS 0.034211f
C870 VDD2.n24 VSUBS 0.015325f
C871 VDD2.n25 VSUBS 1.76759f
C872 VDD2.n26 VSUBS 0.014474f
C873 VDD2.t8 VSUBS 0.073266f
C874 VDD2.n27 VSUBS 0.192972f
C875 VDD2.n28 VSUBS 0.021764f
C876 VDD2.n29 VSUBS 0.025659f
C877 VDD2.n30 VSUBS 0.034211f
C878 VDD2.n31 VSUBS 0.015325f
C879 VDD2.n32 VSUBS 0.014474f
C880 VDD2.n33 VSUBS 0.026936f
C881 VDD2.n34 VSUBS 0.026936f
C882 VDD2.n35 VSUBS 0.014474f
C883 VDD2.n36 VSUBS 0.015325f
C884 VDD2.n37 VSUBS 0.034211f
C885 VDD2.n38 VSUBS 0.034211f
C886 VDD2.n39 VSUBS 0.015325f
C887 VDD2.n40 VSUBS 0.014474f
C888 VDD2.n41 VSUBS 0.026936f
C889 VDD2.n42 VSUBS 0.026936f
C890 VDD2.n43 VSUBS 0.014474f
C891 VDD2.n44 VSUBS 0.015325f
C892 VDD2.n45 VSUBS 0.034211f
C893 VDD2.n46 VSUBS 0.034211f
C894 VDD2.n47 VSUBS 0.015325f
C895 VDD2.n48 VSUBS 0.014474f
C896 VDD2.n49 VSUBS 0.026936f
C897 VDD2.n50 VSUBS 0.026936f
C898 VDD2.n51 VSUBS 0.014474f
C899 VDD2.n52 VSUBS 0.015325f
C900 VDD2.n53 VSUBS 0.034211f
C901 VDD2.n54 VSUBS 0.034211f
C902 VDD2.n55 VSUBS 0.015325f
C903 VDD2.n56 VSUBS 0.014474f
C904 VDD2.n57 VSUBS 0.026936f
C905 VDD2.n58 VSUBS 0.026936f
C906 VDD2.n59 VSUBS 0.014474f
C907 VDD2.n60 VSUBS 0.015325f
C908 VDD2.n61 VSUBS 0.034211f
C909 VDD2.n62 VSUBS 0.034211f
C910 VDD2.n63 VSUBS 0.015325f
C911 VDD2.n64 VSUBS 0.014474f
C912 VDD2.n65 VSUBS 0.026936f
C913 VDD2.n66 VSUBS 0.026936f
C914 VDD2.n67 VSUBS 0.014474f
C915 VDD2.n68 VSUBS 0.014474f
C916 VDD2.n69 VSUBS 0.015325f
C917 VDD2.n70 VSUBS 0.034211f
C918 VDD2.n71 VSUBS 0.034211f
C919 VDD2.n72 VSUBS 0.034211f
C920 VDD2.n73 VSUBS 0.0149f
C921 VDD2.n74 VSUBS 0.014474f
C922 VDD2.n75 VSUBS 0.026936f
C923 VDD2.n76 VSUBS 0.026936f
C924 VDD2.n77 VSUBS 0.014474f
C925 VDD2.n78 VSUBS 0.015325f
C926 VDD2.n79 VSUBS 0.034211f
C927 VDD2.n80 VSUBS 0.077383f
C928 VDD2.n81 VSUBS 0.015325f
C929 VDD2.n82 VSUBS 0.014474f
C930 VDD2.n83 VSUBS 0.063365f
C931 VDD2.n84 VSUBS 0.063878f
C932 VDD2.t4 VSUBS 0.327583f
C933 VDD2.t5 VSUBS 0.327583f
C934 VDD2.n85 VSUBS 2.66919f
C935 VDD2.n86 VSUBS 0.889125f
C936 VDD2.t2 VSUBS 0.327583f
C937 VDD2.t0 VSUBS 0.327583f
C938 VDD2.n87 VSUBS 2.68231f
C939 VDD2.n88 VSUBS 3.09892f
C940 VDD2.n89 VSUBS 0.028f
C941 VDD2.n90 VSUBS 0.026936f
C942 VDD2.n91 VSUBS 0.014474f
C943 VDD2.n92 VSUBS 0.034211f
C944 VDD2.n93 VSUBS 0.0149f
C945 VDD2.n94 VSUBS 0.026936f
C946 VDD2.n95 VSUBS 0.0149f
C947 VDD2.n96 VSUBS 0.014474f
C948 VDD2.n97 VSUBS 0.034211f
C949 VDD2.n98 VSUBS 0.034211f
C950 VDD2.n99 VSUBS 0.015325f
C951 VDD2.n100 VSUBS 0.026936f
C952 VDD2.n101 VSUBS 0.014474f
C953 VDD2.n102 VSUBS 0.034211f
C954 VDD2.n103 VSUBS 0.015325f
C955 VDD2.n104 VSUBS 0.026936f
C956 VDD2.n105 VSUBS 0.014474f
C957 VDD2.n106 VSUBS 0.034211f
C958 VDD2.n107 VSUBS 0.015325f
C959 VDD2.n108 VSUBS 0.026936f
C960 VDD2.n109 VSUBS 0.014474f
C961 VDD2.n110 VSUBS 0.034211f
C962 VDD2.n111 VSUBS 0.015325f
C963 VDD2.n112 VSUBS 0.026936f
C964 VDD2.n113 VSUBS 0.014474f
C965 VDD2.n114 VSUBS 0.034211f
C966 VDD2.n115 VSUBS 0.015325f
C967 VDD2.n116 VSUBS 1.76759f
C968 VDD2.n117 VSUBS 0.014474f
C969 VDD2.t9 VSUBS 0.073266f
C970 VDD2.n118 VSUBS 0.192972f
C971 VDD2.n119 VSUBS 0.021764f
C972 VDD2.n120 VSUBS 0.025659f
C973 VDD2.n121 VSUBS 0.034211f
C974 VDD2.n122 VSUBS 0.015325f
C975 VDD2.n123 VSUBS 0.014474f
C976 VDD2.n124 VSUBS 0.026936f
C977 VDD2.n125 VSUBS 0.026936f
C978 VDD2.n126 VSUBS 0.014474f
C979 VDD2.n127 VSUBS 0.015325f
C980 VDD2.n128 VSUBS 0.034211f
C981 VDD2.n129 VSUBS 0.034211f
C982 VDD2.n130 VSUBS 0.015325f
C983 VDD2.n131 VSUBS 0.014474f
C984 VDD2.n132 VSUBS 0.026936f
C985 VDD2.n133 VSUBS 0.026936f
C986 VDD2.n134 VSUBS 0.014474f
C987 VDD2.n135 VSUBS 0.015325f
C988 VDD2.n136 VSUBS 0.034211f
C989 VDD2.n137 VSUBS 0.034211f
C990 VDD2.n138 VSUBS 0.015325f
C991 VDD2.n139 VSUBS 0.014474f
C992 VDD2.n140 VSUBS 0.026936f
C993 VDD2.n141 VSUBS 0.026936f
C994 VDD2.n142 VSUBS 0.014474f
C995 VDD2.n143 VSUBS 0.015325f
C996 VDD2.n144 VSUBS 0.034211f
C997 VDD2.n145 VSUBS 0.034211f
C998 VDD2.n146 VSUBS 0.015325f
C999 VDD2.n147 VSUBS 0.014474f
C1000 VDD2.n148 VSUBS 0.026936f
C1001 VDD2.n149 VSUBS 0.026936f
C1002 VDD2.n150 VSUBS 0.014474f
C1003 VDD2.n151 VSUBS 0.015325f
C1004 VDD2.n152 VSUBS 0.034211f
C1005 VDD2.n153 VSUBS 0.034211f
C1006 VDD2.n154 VSUBS 0.015325f
C1007 VDD2.n155 VSUBS 0.014474f
C1008 VDD2.n156 VSUBS 0.026936f
C1009 VDD2.n157 VSUBS 0.026936f
C1010 VDD2.n158 VSUBS 0.014474f
C1011 VDD2.n159 VSUBS 0.015325f
C1012 VDD2.n160 VSUBS 0.034211f
C1013 VDD2.n161 VSUBS 0.034211f
C1014 VDD2.n162 VSUBS 0.015325f
C1015 VDD2.n163 VSUBS 0.014474f
C1016 VDD2.n164 VSUBS 0.026936f
C1017 VDD2.n165 VSUBS 0.026936f
C1018 VDD2.n166 VSUBS 0.014474f
C1019 VDD2.n167 VSUBS 0.015325f
C1020 VDD2.n168 VSUBS 0.034211f
C1021 VDD2.n169 VSUBS 0.077383f
C1022 VDD2.n170 VSUBS 0.015325f
C1023 VDD2.n171 VSUBS 0.014474f
C1024 VDD2.n172 VSUBS 0.063365f
C1025 VDD2.n173 VSUBS 0.057297f
C1026 VDD2.n174 VSUBS 2.99009f
C1027 VDD2.t3 VSUBS 0.327583f
C1028 VDD2.t7 VSUBS 0.327583f
C1029 VDD2.n175 VSUBS 2.66921f
C1030 VDD2.n176 VSUBS 0.704697f
C1031 VDD2.t1 VSUBS 0.327583f
C1032 VDD2.t6 VSUBS 0.327583f
C1033 VDD2.n177 VSUBS 2.68226f
C1034 VN.n0 VSUBS 0.034076f
C1035 VN.t9 VSUBS 2.3437f
C1036 VN.n1 VSUBS 0.044047f
C1037 VN.n2 VSUBS 0.034076f
C1038 VN.t7 VSUBS 2.3437f
C1039 VN.n3 VSUBS 0.047845f
C1040 VN.n4 VSUBS 0.034076f
C1041 VN.t4 VSUBS 2.3437f
C1042 VN.n5 VSUBS 0.051644f
C1043 VN.t1 VSUBS 2.46619f
C1044 VN.n6 VSUBS 0.913688f
C1045 VN.t5 VSUBS 2.3437f
C1046 VN.n7 VSUBS 0.894756f
C1047 VN.n8 VSUBS 0.045323f
C1048 VN.n9 VSUBS 0.218118f
C1049 VN.n10 VSUBS 0.034076f
C1050 VN.n11 VSUBS 0.034076f
C1051 VN.n12 VSUBS 0.047845f
C1052 VN.n13 VSUBS 0.047831f
C1053 VN.n14 VSUBS 0.829883f
C1054 VN.n15 VSUBS 0.047831f
C1055 VN.n16 VSUBS 0.034076f
C1056 VN.n17 VSUBS 0.034076f
C1057 VN.n18 VSUBS 0.034076f
C1058 VN.n19 VSUBS 0.051644f
C1059 VN.n20 VSUBS 0.045323f
C1060 VN.n21 VSUBS 0.829883f
C1061 VN.n22 VSUBS 0.05034f
C1062 VN.n23 VSUBS 0.034076f
C1063 VN.n24 VSUBS 0.034076f
C1064 VN.n25 VSUBS 0.034076f
C1065 VN.n26 VSUBS 0.055442f
C1066 VN.n27 VSUBS 0.042814f
C1067 VN.n28 VSUBS 0.904712f
C1068 VN.n29 VSUBS 0.033899f
C1069 VN.n30 VSUBS 0.034076f
C1070 VN.t0 VSUBS 2.3437f
C1071 VN.n31 VSUBS 0.044047f
C1072 VN.n32 VSUBS 0.034076f
C1073 VN.t6 VSUBS 2.3437f
C1074 VN.n33 VSUBS 0.047845f
C1075 VN.n34 VSUBS 0.034076f
C1076 VN.t2 VSUBS 2.3437f
C1077 VN.n35 VSUBS 0.051644f
C1078 VN.t3 VSUBS 2.46619f
C1079 VN.n36 VSUBS 0.913688f
C1080 VN.t8 VSUBS 2.3437f
C1081 VN.n37 VSUBS 0.894756f
C1082 VN.n38 VSUBS 0.045323f
C1083 VN.n39 VSUBS 0.218118f
C1084 VN.n40 VSUBS 0.034076f
C1085 VN.n41 VSUBS 0.034076f
C1086 VN.n42 VSUBS 0.047845f
C1087 VN.n43 VSUBS 0.047831f
C1088 VN.n44 VSUBS 0.829883f
C1089 VN.n45 VSUBS 0.047831f
C1090 VN.n46 VSUBS 0.034076f
C1091 VN.n47 VSUBS 0.034076f
C1092 VN.n48 VSUBS 0.034076f
C1093 VN.n49 VSUBS 0.051644f
C1094 VN.n50 VSUBS 0.045323f
C1095 VN.n51 VSUBS 0.829883f
C1096 VN.n52 VSUBS 0.05034f
C1097 VN.n53 VSUBS 0.034076f
C1098 VN.n54 VSUBS 0.034076f
C1099 VN.n55 VSUBS 0.034076f
C1100 VN.n56 VSUBS 0.055442f
C1101 VN.n57 VSUBS 0.042814f
C1102 VN.n58 VSUBS 0.904712f
C1103 VN.n59 VSUBS 1.90124f
C1104 VDD1.n0 VSUBS 0.028f
C1105 VDD1.n1 VSUBS 0.026936f
C1106 VDD1.n2 VSUBS 0.014474f
C1107 VDD1.n3 VSUBS 0.034212f
C1108 VDD1.n4 VSUBS 0.0149f
C1109 VDD1.n5 VSUBS 0.026936f
C1110 VDD1.n6 VSUBS 0.0149f
C1111 VDD1.n7 VSUBS 0.014474f
C1112 VDD1.n8 VSUBS 0.034212f
C1113 VDD1.n9 VSUBS 0.034212f
C1114 VDD1.n10 VSUBS 0.015326f
C1115 VDD1.n11 VSUBS 0.026936f
C1116 VDD1.n12 VSUBS 0.014474f
C1117 VDD1.n13 VSUBS 0.034212f
C1118 VDD1.n14 VSUBS 0.015326f
C1119 VDD1.n15 VSUBS 0.026936f
C1120 VDD1.n16 VSUBS 0.014474f
C1121 VDD1.n17 VSUBS 0.034212f
C1122 VDD1.n18 VSUBS 0.015326f
C1123 VDD1.n19 VSUBS 0.026936f
C1124 VDD1.n20 VSUBS 0.014474f
C1125 VDD1.n21 VSUBS 0.034212f
C1126 VDD1.n22 VSUBS 0.015326f
C1127 VDD1.n23 VSUBS 0.026936f
C1128 VDD1.n24 VSUBS 0.014474f
C1129 VDD1.n25 VSUBS 0.034212f
C1130 VDD1.n26 VSUBS 0.015326f
C1131 VDD1.n27 VSUBS 1.76762f
C1132 VDD1.n28 VSUBS 0.014474f
C1133 VDD1.t0 VSUBS 0.073267f
C1134 VDD1.n29 VSUBS 0.192975f
C1135 VDD1.n30 VSUBS 0.021764f
C1136 VDD1.n31 VSUBS 0.025659f
C1137 VDD1.n32 VSUBS 0.034212f
C1138 VDD1.n33 VSUBS 0.015326f
C1139 VDD1.n34 VSUBS 0.014474f
C1140 VDD1.n35 VSUBS 0.026936f
C1141 VDD1.n36 VSUBS 0.026936f
C1142 VDD1.n37 VSUBS 0.014474f
C1143 VDD1.n38 VSUBS 0.015326f
C1144 VDD1.n39 VSUBS 0.034212f
C1145 VDD1.n40 VSUBS 0.034212f
C1146 VDD1.n41 VSUBS 0.015326f
C1147 VDD1.n42 VSUBS 0.014474f
C1148 VDD1.n43 VSUBS 0.026936f
C1149 VDD1.n44 VSUBS 0.026936f
C1150 VDD1.n45 VSUBS 0.014474f
C1151 VDD1.n46 VSUBS 0.015326f
C1152 VDD1.n47 VSUBS 0.034212f
C1153 VDD1.n48 VSUBS 0.034212f
C1154 VDD1.n49 VSUBS 0.015326f
C1155 VDD1.n50 VSUBS 0.014474f
C1156 VDD1.n51 VSUBS 0.026936f
C1157 VDD1.n52 VSUBS 0.026936f
C1158 VDD1.n53 VSUBS 0.014474f
C1159 VDD1.n54 VSUBS 0.015326f
C1160 VDD1.n55 VSUBS 0.034212f
C1161 VDD1.n56 VSUBS 0.034212f
C1162 VDD1.n57 VSUBS 0.015326f
C1163 VDD1.n58 VSUBS 0.014474f
C1164 VDD1.n59 VSUBS 0.026936f
C1165 VDD1.n60 VSUBS 0.026936f
C1166 VDD1.n61 VSUBS 0.014474f
C1167 VDD1.n62 VSUBS 0.015326f
C1168 VDD1.n63 VSUBS 0.034212f
C1169 VDD1.n64 VSUBS 0.034212f
C1170 VDD1.n65 VSUBS 0.015326f
C1171 VDD1.n66 VSUBS 0.014474f
C1172 VDD1.n67 VSUBS 0.026936f
C1173 VDD1.n68 VSUBS 0.026936f
C1174 VDD1.n69 VSUBS 0.014474f
C1175 VDD1.n70 VSUBS 0.015326f
C1176 VDD1.n71 VSUBS 0.034212f
C1177 VDD1.n72 VSUBS 0.034212f
C1178 VDD1.n73 VSUBS 0.015326f
C1179 VDD1.n74 VSUBS 0.014474f
C1180 VDD1.n75 VSUBS 0.026936f
C1181 VDD1.n76 VSUBS 0.026936f
C1182 VDD1.n77 VSUBS 0.014474f
C1183 VDD1.n78 VSUBS 0.015326f
C1184 VDD1.n79 VSUBS 0.034212f
C1185 VDD1.n80 VSUBS 0.077384f
C1186 VDD1.n81 VSUBS 0.015326f
C1187 VDD1.n82 VSUBS 0.014474f
C1188 VDD1.n83 VSUBS 0.063366f
C1189 VDD1.n84 VSUBS 0.063879f
C1190 VDD1.t4 VSUBS 0.327588f
C1191 VDD1.t2 VSUBS 0.327588f
C1192 VDD1.n85 VSUBS 2.66925f
C1193 VDD1.n86 VSUBS 0.897281f
C1194 VDD1.n87 VSUBS 0.028f
C1195 VDD1.n88 VSUBS 0.026936f
C1196 VDD1.n89 VSUBS 0.014474f
C1197 VDD1.n90 VSUBS 0.034212f
C1198 VDD1.n91 VSUBS 0.0149f
C1199 VDD1.n92 VSUBS 0.026936f
C1200 VDD1.n93 VSUBS 0.015326f
C1201 VDD1.n94 VSUBS 0.034212f
C1202 VDD1.n95 VSUBS 0.015326f
C1203 VDD1.n96 VSUBS 0.026936f
C1204 VDD1.n97 VSUBS 0.014474f
C1205 VDD1.n98 VSUBS 0.034212f
C1206 VDD1.n99 VSUBS 0.015326f
C1207 VDD1.n100 VSUBS 0.026936f
C1208 VDD1.n101 VSUBS 0.014474f
C1209 VDD1.n102 VSUBS 0.034212f
C1210 VDD1.n103 VSUBS 0.015326f
C1211 VDD1.n104 VSUBS 0.026936f
C1212 VDD1.n105 VSUBS 0.014474f
C1213 VDD1.n106 VSUBS 0.034212f
C1214 VDD1.n107 VSUBS 0.015326f
C1215 VDD1.n108 VSUBS 0.026936f
C1216 VDD1.n109 VSUBS 0.014474f
C1217 VDD1.n110 VSUBS 0.034212f
C1218 VDD1.n111 VSUBS 0.015326f
C1219 VDD1.n112 VSUBS 1.76762f
C1220 VDD1.n113 VSUBS 0.014474f
C1221 VDD1.t6 VSUBS 0.073267f
C1222 VDD1.n114 VSUBS 0.192975f
C1223 VDD1.n115 VSUBS 0.021764f
C1224 VDD1.n116 VSUBS 0.025659f
C1225 VDD1.n117 VSUBS 0.034212f
C1226 VDD1.n118 VSUBS 0.015326f
C1227 VDD1.n119 VSUBS 0.014474f
C1228 VDD1.n120 VSUBS 0.026936f
C1229 VDD1.n121 VSUBS 0.026936f
C1230 VDD1.n122 VSUBS 0.014474f
C1231 VDD1.n123 VSUBS 0.015326f
C1232 VDD1.n124 VSUBS 0.034212f
C1233 VDD1.n125 VSUBS 0.034212f
C1234 VDD1.n126 VSUBS 0.015326f
C1235 VDD1.n127 VSUBS 0.014474f
C1236 VDD1.n128 VSUBS 0.026936f
C1237 VDD1.n129 VSUBS 0.026936f
C1238 VDD1.n130 VSUBS 0.014474f
C1239 VDD1.n131 VSUBS 0.015326f
C1240 VDD1.n132 VSUBS 0.034212f
C1241 VDD1.n133 VSUBS 0.034212f
C1242 VDD1.n134 VSUBS 0.015326f
C1243 VDD1.n135 VSUBS 0.014474f
C1244 VDD1.n136 VSUBS 0.026936f
C1245 VDD1.n137 VSUBS 0.026936f
C1246 VDD1.n138 VSUBS 0.014474f
C1247 VDD1.n139 VSUBS 0.015326f
C1248 VDD1.n140 VSUBS 0.034212f
C1249 VDD1.n141 VSUBS 0.034212f
C1250 VDD1.n142 VSUBS 0.015326f
C1251 VDD1.n143 VSUBS 0.014474f
C1252 VDD1.n144 VSUBS 0.026936f
C1253 VDD1.n145 VSUBS 0.026936f
C1254 VDD1.n146 VSUBS 0.014474f
C1255 VDD1.n147 VSUBS 0.015326f
C1256 VDD1.n148 VSUBS 0.034212f
C1257 VDD1.n149 VSUBS 0.034212f
C1258 VDD1.n150 VSUBS 0.015326f
C1259 VDD1.n151 VSUBS 0.014474f
C1260 VDD1.n152 VSUBS 0.026936f
C1261 VDD1.n153 VSUBS 0.026936f
C1262 VDD1.n154 VSUBS 0.014474f
C1263 VDD1.n155 VSUBS 0.014474f
C1264 VDD1.n156 VSUBS 0.015326f
C1265 VDD1.n157 VSUBS 0.034212f
C1266 VDD1.n158 VSUBS 0.034212f
C1267 VDD1.n159 VSUBS 0.034212f
C1268 VDD1.n160 VSUBS 0.0149f
C1269 VDD1.n161 VSUBS 0.014474f
C1270 VDD1.n162 VSUBS 0.026936f
C1271 VDD1.n163 VSUBS 0.026936f
C1272 VDD1.n164 VSUBS 0.014474f
C1273 VDD1.n165 VSUBS 0.015326f
C1274 VDD1.n166 VSUBS 0.034212f
C1275 VDD1.n167 VSUBS 0.077384f
C1276 VDD1.n168 VSUBS 0.015326f
C1277 VDD1.n169 VSUBS 0.014474f
C1278 VDD1.n170 VSUBS 0.063366f
C1279 VDD1.n171 VSUBS 0.063879f
C1280 VDD1.t7 VSUBS 0.327588f
C1281 VDD1.t9 VSUBS 0.327588f
C1282 VDD1.n172 VSUBS 2.66924f
C1283 VDD1.n173 VSUBS 0.88914f
C1284 VDD1.t1 VSUBS 0.327588f
C1285 VDD1.t3 VSUBS 0.327588f
C1286 VDD1.n174 VSUBS 2.68235f
C1287 VDD1.n175 VSUBS 3.20819f
C1288 VDD1.t8 VSUBS 0.327588f
C1289 VDD1.t5 VSUBS 0.327588f
C1290 VDD1.n176 VSUBS 2.66924f
C1291 VDD1.n177 VSUBS 3.56005f
C1292 VTAIL.t5 VSUBS 0.333661f
C1293 VTAIL.t2 VSUBS 0.333661f
C1294 VTAIL.n0 VSUBS 2.55837f
C1295 VTAIL.n1 VSUBS 0.88238f
C1296 VTAIL.n2 VSUBS 0.028519f
C1297 VTAIL.n3 VSUBS 0.027436f
C1298 VTAIL.n4 VSUBS 0.014743f
C1299 VTAIL.n5 VSUBS 0.034846f
C1300 VTAIL.n6 VSUBS 0.015176f
C1301 VTAIL.n7 VSUBS 0.027436f
C1302 VTAIL.n8 VSUBS 0.01561f
C1303 VTAIL.n9 VSUBS 0.034846f
C1304 VTAIL.n10 VSUBS 0.01561f
C1305 VTAIL.n11 VSUBS 0.027436f
C1306 VTAIL.n12 VSUBS 0.014743f
C1307 VTAIL.n13 VSUBS 0.034846f
C1308 VTAIL.n14 VSUBS 0.01561f
C1309 VTAIL.n15 VSUBS 0.027436f
C1310 VTAIL.n16 VSUBS 0.014743f
C1311 VTAIL.n17 VSUBS 0.034846f
C1312 VTAIL.n18 VSUBS 0.01561f
C1313 VTAIL.n19 VSUBS 0.027436f
C1314 VTAIL.n20 VSUBS 0.014743f
C1315 VTAIL.n21 VSUBS 0.034846f
C1316 VTAIL.n22 VSUBS 0.01561f
C1317 VTAIL.n23 VSUBS 0.027436f
C1318 VTAIL.n24 VSUBS 0.014743f
C1319 VTAIL.n25 VSUBS 0.034846f
C1320 VTAIL.n26 VSUBS 0.01561f
C1321 VTAIL.n27 VSUBS 1.80039f
C1322 VTAIL.n28 VSUBS 0.014743f
C1323 VTAIL.t13 VSUBS 0.074625f
C1324 VTAIL.n29 VSUBS 0.196552f
C1325 VTAIL.n30 VSUBS 0.022168f
C1326 VTAIL.n31 VSUBS 0.026135f
C1327 VTAIL.n32 VSUBS 0.034846f
C1328 VTAIL.n33 VSUBS 0.01561f
C1329 VTAIL.n34 VSUBS 0.014743f
C1330 VTAIL.n35 VSUBS 0.027436f
C1331 VTAIL.n36 VSUBS 0.027436f
C1332 VTAIL.n37 VSUBS 0.014743f
C1333 VTAIL.n38 VSUBS 0.01561f
C1334 VTAIL.n39 VSUBS 0.034846f
C1335 VTAIL.n40 VSUBS 0.034846f
C1336 VTAIL.n41 VSUBS 0.01561f
C1337 VTAIL.n42 VSUBS 0.014743f
C1338 VTAIL.n43 VSUBS 0.027436f
C1339 VTAIL.n44 VSUBS 0.027436f
C1340 VTAIL.n45 VSUBS 0.014743f
C1341 VTAIL.n46 VSUBS 0.01561f
C1342 VTAIL.n47 VSUBS 0.034846f
C1343 VTAIL.n48 VSUBS 0.034846f
C1344 VTAIL.n49 VSUBS 0.01561f
C1345 VTAIL.n50 VSUBS 0.014743f
C1346 VTAIL.n51 VSUBS 0.027436f
C1347 VTAIL.n52 VSUBS 0.027436f
C1348 VTAIL.n53 VSUBS 0.014743f
C1349 VTAIL.n54 VSUBS 0.01561f
C1350 VTAIL.n55 VSUBS 0.034846f
C1351 VTAIL.n56 VSUBS 0.034846f
C1352 VTAIL.n57 VSUBS 0.01561f
C1353 VTAIL.n58 VSUBS 0.014743f
C1354 VTAIL.n59 VSUBS 0.027436f
C1355 VTAIL.n60 VSUBS 0.027436f
C1356 VTAIL.n61 VSUBS 0.014743f
C1357 VTAIL.n62 VSUBS 0.01561f
C1358 VTAIL.n63 VSUBS 0.034846f
C1359 VTAIL.n64 VSUBS 0.034846f
C1360 VTAIL.n65 VSUBS 0.01561f
C1361 VTAIL.n66 VSUBS 0.014743f
C1362 VTAIL.n67 VSUBS 0.027436f
C1363 VTAIL.n68 VSUBS 0.027436f
C1364 VTAIL.n69 VSUBS 0.014743f
C1365 VTAIL.n70 VSUBS 0.014743f
C1366 VTAIL.n71 VSUBS 0.01561f
C1367 VTAIL.n72 VSUBS 0.034846f
C1368 VTAIL.n73 VSUBS 0.034846f
C1369 VTAIL.n74 VSUBS 0.034846f
C1370 VTAIL.n75 VSUBS 0.015176f
C1371 VTAIL.n76 VSUBS 0.014743f
C1372 VTAIL.n77 VSUBS 0.027436f
C1373 VTAIL.n78 VSUBS 0.027436f
C1374 VTAIL.n79 VSUBS 0.014743f
C1375 VTAIL.n80 VSUBS 0.01561f
C1376 VTAIL.n81 VSUBS 0.034846f
C1377 VTAIL.n82 VSUBS 0.078818f
C1378 VTAIL.n83 VSUBS 0.01561f
C1379 VTAIL.n84 VSUBS 0.014743f
C1380 VTAIL.n85 VSUBS 0.06454f
C1381 VTAIL.n86 VSUBS 0.039425f
C1382 VTAIL.n87 VSUBS 0.289658f
C1383 VTAIL.t11 VSUBS 0.333661f
C1384 VTAIL.t17 VSUBS 0.333661f
C1385 VTAIL.n88 VSUBS 2.55837f
C1386 VTAIL.n89 VSUBS 0.94773f
C1387 VTAIL.t19 VSUBS 0.333661f
C1388 VTAIL.t15 VSUBS 0.333661f
C1389 VTAIL.n90 VSUBS 2.55837f
C1390 VTAIL.n91 VSUBS 2.64265f
C1391 VTAIL.t7 VSUBS 0.333661f
C1392 VTAIL.t3 VSUBS 0.333661f
C1393 VTAIL.n92 VSUBS 2.55838f
C1394 VTAIL.n93 VSUBS 2.64263f
C1395 VTAIL.t8 VSUBS 0.333661f
C1396 VTAIL.t1 VSUBS 0.333661f
C1397 VTAIL.n94 VSUBS 2.55838f
C1398 VTAIL.n95 VSUBS 0.947713f
C1399 VTAIL.n96 VSUBS 0.028519f
C1400 VTAIL.n97 VSUBS 0.027436f
C1401 VTAIL.n98 VSUBS 0.014743f
C1402 VTAIL.n99 VSUBS 0.034846f
C1403 VTAIL.n100 VSUBS 0.015176f
C1404 VTAIL.n101 VSUBS 0.027436f
C1405 VTAIL.n102 VSUBS 0.015176f
C1406 VTAIL.n103 VSUBS 0.014743f
C1407 VTAIL.n104 VSUBS 0.034846f
C1408 VTAIL.n105 VSUBS 0.034846f
C1409 VTAIL.n106 VSUBS 0.01561f
C1410 VTAIL.n107 VSUBS 0.027436f
C1411 VTAIL.n108 VSUBS 0.014743f
C1412 VTAIL.n109 VSUBS 0.034846f
C1413 VTAIL.n110 VSUBS 0.01561f
C1414 VTAIL.n111 VSUBS 0.027436f
C1415 VTAIL.n112 VSUBS 0.014743f
C1416 VTAIL.n113 VSUBS 0.034846f
C1417 VTAIL.n114 VSUBS 0.01561f
C1418 VTAIL.n115 VSUBS 0.027436f
C1419 VTAIL.n116 VSUBS 0.014743f
C1420 VTAIL.n117 VSUBS 0.034846f
C1421 VTAIL.n118 VSUBS 0.01561f
C1422 VTAIL.n119 VSUBS 0.027436f
C1423 VTAIL.n120 VSUBS 0.014743f
C1424 VTAIL.n121 VSUBS 0.034846f
C1425 VTAIL.n122 VSUBS 0.01561f
C1426 VTAIL.n123 VSUBS 1.80039f
C1427 VTAIL.n124 VSUBS 0.014743f
C1428 VTAIL.t9 VSUBS 0.074625f
C1429 VTAIL.n125 VSUBS 0.196552f
C1430 VTAIL.n126 VSUBS 0.022168f
C1431 VTAIL.n127 VSUBS 0.026135f
C1432 VTAIL.n128 VSUBS 0.034846f
C1433 VTAIL.n129 VSUBS 0.01561f
C1434 VTAIL.n130 VSUBS 0.014743f
C1435 VTAIL.n131 VSUBS 0.027436f
C1436 VTAIL.n132 VSUBS 0.027436f
C1437 VTAIL.n133 VSUBS 0.014743f
C1438 VTAIL.n134 VSUBS 0.01561f
C1439 VTAIL.n135 VSUBS 0.034846f
C1440 VTAIL.n136 VSUBS 0.034846f
C1441 VTAIL.n137 VSUBS 0.01561f
C1442 VTAIL.n138 VSUBS 0.014743f
C1443 VTAIL.n139 VSUBS 0.027436f
C1444 VTAIL.n140 VSUBS 0.027436f
C1445 VTAIL.n141 VSUBS 0.014743f
C1446 VTAIL.n142 VSUBS 0.01561f
C1447 VTAIL.n143 VSUBS 0.034846f
C1448 VTAIL.n144 VSUBS 0.034846f
C1449 VTAIL.n145 VSUBS 0.01561f
C1450 VTAIL.n146 VSUBS 0.014743f
C1451 VTAIL.n147 VSUBS 0.027436f
C1452 VTAIL.n148 VSUBS 0.027436f
C1453 VTAIL.n149 VSUBS 0.014743f
C1454 VTAIL.n150 VSUBS 0.01561f
C1455 VTAIL.n151 VSUBS 0.034846f
C1456 VTAIL.n152 VSUBS 0.034846f
C1457 VTAIL.n153 VSUBS 0.01561f
C1458 VTAIL.n154 VSUBS 0.014743f
C1459 VTAIL.n155 VSUBS 0.027436f
C1460 VTAIL.n156 VSUBS 0.027436f
C1461 VTAIL.n157 VSUBS 0.014743f
C1462 VTAIL.n158 VSUBS 0.01561f
C1463 VTAIL.n159 VSUBS 0.034846f
C1464 VTAIL.n160 VSUBS 0.034846f
C1465 VTAIL.n161 VSUBS 0.01561f
C1466 VTAIL.n162 VSUBS 0.014743f
C1467 VTAIL.n163 VSUBS 0.027436f
C1468 VTAIL.n164 VSUBS 0.027436f
C1469 VTAIL.n165 VSUBS 0.014743f
C1470 VTAIL.n166 VSUBS 0.01561f
C1471 VTAIL.n167 VSUBS 0.034846f
C1472 VTAIL.n168 VSUBS 0.034846f
C1473 VTAIL.n169 VSUBS 0.01561f
C1474 VTAIL.n170 VSUBS 0.014743f
C1475 VTAIL.n171 VSUBS 0.027436f
C1476 VTAIL.n172 VSUBS 0.027436f
C1477 VTAIL.n173 VSUBS 0.014743f
C1478 VTAIL.n174 VSUBS 0.01561f
C1479 VTAIL.n175 VSUBS 0.034846f
C1480 VTAIL.n176 VSUBS 0.078818f
C1481 VTAIL.n177 VSUBS 0.01561f
C1482 VTAIL.n178 VSUBS 0.014743f
C1483 VTAIL.n179 VSUBS 0.06454f
C1484 VTAIL.n180 VSUBS 0.039425f
C1485 VTAIL.n181 VSUBS 0.289658f
C1486 VTAIL.t10 VSUBS 0.333661f
C1487 VTAIL.t16 VSUBS 0.333661f
C1488 VTAIL.n182 VSUBS 2.55838f
C1489 VTAIL.n183 VSUBS 0.914562f
C1490 VTAIL.t12 VSUBS 0.333661f
C1491 VTAIL.t18 VSUBS 0.333661f
C1492 VTAIL.n184 VSUBS 2.55838f
C1493 VTAIL.n185 VSUBS 0.947713f
C1494 VTAIL.n186 VSUBS 0.028519f
C1495 VTAIL.n187 VSUBS 0.027436f
C1496 VTAIL.n188 VSUBS 0.014743f
C1497 VTAIL.n189 VSUBS 0.034846f
C1498 VTAIL.n190 VSUBS 0.015176f
C1499 VTAIL.n191 VSUBS 0.027436f
C1500 VTAIL.n192 VSUBS 0.015176f
C1501 VTAIL.n193 VSUBS 0.014743f
C1502 VTAIL.n194 VSUBS 0.034846f
C1503 VTAIL.n195 VSUBS 0.034846f
C1504 VTAIL.n196 VSUBS 0.01561f
C1505 VTAIL.n197 VSUBS 0.027436f
C1506 VTAIL.n198 VSUBS 0.014743f
C1507 VTAIL.n199 VSUBS 0.034846f
C1508 VTAIL.n200 VSUBS 0.01561f
C1509 VTAIL.n201 VSUBS 0.027436f
C1510 VTAIL.n202 VSUBS 0.014743f
C1511 VTAIL.n203 VSUBS 0.034846f
C1512 VTAIL.n204 VSUBS 0.01561f
C1513 VTAIL.n205 VSUBS 0.027436f
C1514 VTAIL.n206 VSUBS 0.014743f
C1515 VTAIL.n207 VSUBS 0.034846f
C1516 VTAIL.n208 VSUBS 0.01561f
C1517 VTAIL.n209 VSUBS 0.027436f
C1518 VTAIL.n210 VSUBS 0.014743f
C1519 VTAIL.n211 VSUBS 0.034846f
C1520 VTAIL.n212 VSUBS 0.01561f
C1521 VTAIL.n213 VSUBS 1.80039f
C1522 VTAIL.n214 VSUBS 0.014743f
C1523 VTAIL.t14 VSUBS 0.074625f
C1524 VTAIL.n215 VSUBS 0.196552f
C1525 VTAIL.n216 VSUBS 0.022168f
C1526 VTAIL.n217 VSUBS 0.026135f
C1527 VTAIL.n218 VSUBS 0.034846f
C1528 VTAIL.n219 VSUBS 0.01561f
C1529 VTAIL.n220 VSUBS 0.014743f
C1530 VTAIL.n221 VSUBS 0.027436f
C1531 VTAIL.n222 VSUBS 0.027436f
C1532 VTAIL.n223 VSUBS 0.014743f
C1533 VTAIL.n224 VSUBS 0.01561f
C1534 VTAIL.n225 VSUBS 0.034846f
C1535 VTAIL.n226 VSUBS 0.034846f
C1536 VTAIL.n227 VSUBS 0.01561f
C1537 VTAIL.n228 VSUBS 0.014743f
C1538 VTAIL.n229 VSUBS 0.027436f
C1539 VTAIL.n230 VSUBS 0.027436f
C1540 VTAIL.n231 VSUBS 0.014743f
C1541 VTAIL.n232 VSUBS 0.01561f
C1542 VTAIL.n233 VSUBS 0.034846f
C1543 VTAIL.n234 VSUBS 0.034846f
C1544 VTAIL.n235 VSUBS 0.01561f
C1545 VTAIL.n236 VSUBS 0.014743f
C1546 VTAIL.n237 VSUBS 0.027436f
C1547 VTAIL.n238 VSUBS 0.027436f
C1548 VTAIL.n239 VSUBS 0.014743f
C1549 VTAIL.n240 VSUBS 0.01561f
C1550 VTAIL.n241 VSUBS 0.034846f
C1551 VTAIL.n242 VSUBS 0.034846f
C1552 VTAIL.n243 VSUBS 0.01561f
C1553 VTAIL.n244 VSUBS 0.014743f
C1554 VTAIL.n245 VSUBS 0.027436f
C1555 VTAIL.n246 VSUBS 0.027436f
C1556 VTAIL.n247 VSUBS 0.014743f
C1557 VTAIL.n248 VSUBS 0.01561f
C1558 VTAIL.n249 VSUBS 0.034846f
C1559 VTAIL.n250 VSUBS 0.034846f
C1560 VTAIL.n251 VSUBS 0.01561f
C1561 VTAIL.n252 VSUBS 0.014743f
C1562 VTAIL.n253 VSUBS 0.027436f
C1563 VTAIL.n254 VSUBS 0.027436f
C1564 VTAIL.n255 VSUBS 0.014743f
C1565 VTAIL.n256 VSUBS 0.01561f
C1566 VTAIL.n257 VSUBS 0.034846f
C1567 VTAIL.n258 VSUBS 0.034846f
C1568 VTAIL.n259 VSUBS 0.01561f
C1569 VTAIL.n260 VSUBS 0.014743f
C1570 VTAIL.n261 VSUBS 0.027436f
C1571 VTAIL.n262 VSUBS 0.027436f
C1572 VTAIL.n263 VSUBS 0.014743f
C1573 VTAIL.n264 VSUBS 0.01561f
C1574 VTAIL.n265 VSUBS 0.034846f
C1575 VTAIL.n266 VSUBS 0.078818f
C1576 VTAIL.n267 VSUBS 0.01561f
C1577 VTAIL.n268 VSUBS 0.014743f
C1578 VTAIL.n269 VSUBS 0.06454f
C1579 VTAIL.n270 VSUBS 0.039425f
C1580 VTAIL.n271 VSUBS 1.86836f
C1581 VTAIL.n272 VSUBS 0.028519f
C1582 VTAIL.n273 VSUBS 0.027436f
C1583 VTAIL.n274 VSUBS 0.014743f
C1584 VTAIL.n275 VSUBS 0.034846f
C1585 VTAIL.n276 VSUBS 0.015176f
C1586 VTAIL.n277 VSUBS 0.027436f
C1587 VTAIL.n278 VSUBS 0.01561f
C1588 VTAIL.n279 VSUBS 0.034846f
C1589 VTAIL.n280 VSUBS 0.01561f
C1590 VTAIL.n281 VSUBS 0.027436f
C1591 VTAIL.n282 VSUBS 0.014743f
C1592 VTAIL.n283 VSUBS 0.034846f
C1593 VTAIL.n284 VSUBS 0.01561f
C1594 VTAIL.n285 VSUBS 0.027436f
C1595 VTAIL.n286 VSUBS 0.014743f
C1596 VTAIL.n287 VSUBS 0.034846f
C1597 VTAIL.n288 VSUBS 0.01561f
C1598 VTAIL.n289 VSUBS 0.027436f
C1599 VTAIL.n290 VSUBS 0.014743f
C1600 VTAIL.n291 VSUBS 0.034846f
C1601 VTAIL.n292 VSUBS 0.01561f
C1602 VTAIL.n293 VSUBS 0.027436f
C1603 VTAIL.n294 VSUBS 0.014743f
C1604 VTAIL.n295 VSUBS 0.034846f
C1605 VTAIL.n296 VSUBS 0.01561f
C1606 VTAIL.n297 VSUBS 1.80039f
C1607 VTAIL.n298 VSUBS 0.014743f
C1608 VTAIL.t6 VSUBS 0.074625f
C1609 VTAIL.n299 VSUBS 0.196552f
C1610 VTAIL.n300 VSUBS 0.022168f
C1611 VTAIL.n301 VSUBS 0.026135f
C1612 VTAIL.n302 VSUBS 0.034846f
C1613 VTAIL.n303 VSUBS 0.01561f
C1614 VTAIL.n304 VSUBS 0.014743f
C1615 VTAIL.n305 VSUBS 0.027436f
C1616 VTAIL.n306 VSUBS 0.027436f
C1617 VTAIL.n307 VSUBS 0.014743f
C1618 VTAIL.n308 VSUBS 0.01561f
C1619 VTAIL.n309 VSUBS 0.034846f
C1620 VTAIL.n310 VSUBS 0.034846f
C1621 VTAIL.n311 VSUBS 0.01561f
C1622 VTAIL.n312 VSUBS 0.014743f
C1623 VTAIL.n313 VSUBS 0.027436f
C1624 VTAIL.n314 VSUBS 0.027436f
C1625 VTAIL.n315 VSUBS 0.014743f
C1626 VTAIL.n316 VSUBS 0.01561f
C1627 VTAIL.n317 VSUBS 0.034846f
C1628 VTAIL.n318 VSUBS 0.034846f
C1629 VTAIL.n319 VSUBS 0.01561f
C1630 VTAIL.n320 VSUBS 0.014743f
C1631 VTAIL.n321 VSUBS 0.027436f
C1632 VTAIL.n322 VSUBS 0.027436f
C1633 VTAIL.n323 VSUBS 0.014743f
C1634 VTAIL.n324 VSUBS 0.01561f
C1635 VTAIL.n325 VSUBS 0.034846f
C1636 VTAIL.n326 VSUBS 0.034846f
C1637 VTAIL.n327 VSUBS 0.01561f
C1638 VTAIL.n328 VSUBS 0.014743f
C1639 VTAIL.n329 VSUBS 0.027436f
C1640 VTAIL.n330 VSUBS 0.027436f
C1641 VTAIL.n331 VSUBS 0.014743f
C1642 VTAIL.n332 VSUBS 0.01561f
C1643 VTAIL.n333 VSUBS 0.034846f
C1644 VTAIL.n334 VSUBS 0.034846f
C1645 VTAIL.n335 VSUBS 0.01561f
C1646 VTAIL.n336 VSUBS 0.014743f
C1647 VTAIL.n337 VSUBS 0.027436f
C1648 VTAIL.n338 VSUBS 0.027436f
C1649 VTAIL.n339 VSUBS 0.014743f
C1650 VTAIL.n340 VSUBS 0.014743f
C1651 VTAIL.n341 VSUBS 0.01561f
C1652 VTAIL.n342 VSUBS 0.034846f
C1653 VTAIL.n343 VSUBS 0.034846f
C1654 VTAIL.n344 VSUBS 0.034846f
C1655 VTAIL.n345 VSUBS 0.015176f
C1656 VTAIL.n346 VSUBS 0.014743f
C1657 VTAIL.n347 VSUBS 0.027436f
C1658 VTAIL.n348 VSUBS 0.027436f
C1659 VTAIL.n349 VSUBS 0.014743f
C1660 VTAIL.n350 VSUBS 0.01561f
C1661 VTAIL.n351 VSUBS 0.034846f
C1662 VTAIL.n352 VSUBS 0.078818f
C1663 VTAIL.n353 VSUBS 0.01561f
C1664 VTAIL.n354 VSUBS 0.014743f
C1665 VTAIL.n355 VSUBS 0.06454f
C1666 VTAIL.n356 VSUBS 0.039425f
C1667 VTAIL.n357 VSUBS 1.86836f
C1668 VTAIL.t4 VSUBS 0.333661f
C1669 VTAIL.t0 VSUBS 0.333661f
C1670 VTAIL.n358 VSUBS 2.55837f
C1671 VTAIL.n359 VSUBS 0.830557f
C1672 VP.n0 VSUBS 0.034825f
C1673 VP.t6 VSUBS 2.39524f
C1674 VP.n1 VSUBS 0.045016f
C1675 VP.n2 VSUBS 0.034825f
C1676 VP.t8 VSUBS 2.39524f
C1677 VP.n3 VSUBS 0.048897f
C1678 VP.n4 VSUBS 0.034825f
C1679 VP.t0 VSUBS 2.39524f
C1680 VP.n5 VSUBS 0.052779f
C1681 VP.n6 VSUBS 0.034825f
C1682 VP.t2 VSUBS 2.39524f
C1683 VP.n7 VSUBS 0.056661f
C1684 VP.n8 VSUBS 0.034825f
C1685 VP.t4 VSUBS 2.39524f
C1686 VP.n9 VSUBS 0.045016f
C1687 VP.n10 VSUBS 0.034825f
C1688 VP.t1 VSUBS 2.39524f
C1689 VP.n11 VSUBS 0.048897f
C1690 VP.n12 VSUBS 0.034825f
C1691 VP.t7 VSUBS 2.39524f
C1692 VP.n13 VSUBS 0.052779f
C1693 VP.t9 VSUBS 2.52043f
C1694 VP.n14 VSUBS 0.933784f
C1695 VP.t5 VSUBS 2.39524f
C1696 VP.n15 VSUBS 0.914434f
C1697 VP.n16 VSUBS 0.04632f
C1698 VP.n17 VSUBS 0.222915f
C1699 VP.n18 VSUBS 0.034825f
C1700 VP.n19 VSUBS 0.034825f
C1701 VP.n20 VSUBS 0.048897f
C1702 VP.n21 VSUBS 0.048883f
C1703 VP.n22 VSUBS 0.848135f
C1704 VP.n23 VSUBS 0.048883f
C1705 VP.n24 VSUBS 0.034825f
C1706 VP.n25 VSUBS 0.034825f
C1707 VP.n26 VSUBS 0.034825f
C1708 VP.n27 VSUBS 0.052779f
C1709 VP.n28 VSUBS 0.04632f
C1710 VP.n29 VSUBS 0.848135f
C1711 VP.n30 VSUBS 0.051447f
C1712 VP.n31 VSUBS 0.034825f
C1713 VP.n32 VSUBS 0.034825f
C1714 VP.n33 VSUBS 0.034825f
C1715 VP.n34 VSUBS 0.056661f
C1716 VP.n35 VSUBS 0.043756f
C1717 VP.n36 VSUBS 0.92461f
C1718 VP.n37 VSUBS 1.92042f
C1719 VP.n38 VSUBS 1.94529f
C1720 VP.t3 VSUBS 2.39524f
C1721 VP.n39 VSUBS 0.92461f
C1722 VP.n40 VSUBS 0.043756f
C1723 VP.n41 VSUBS 0.034825f
C1724 VP.n42 VSUBS 0.034825f
C1725 VP.n43 VSUBS 0.034825f
C1726 VP.n44 VSUBS 0.045016f
C1727 VP.n45 VSUBS 0.051447f
C1728 VP.n46 VSUBS 0.848135f
C1729 VP.n47 VSUBS 0.04632f
C1730 VP.n48 VSUBS 0.034825f
C1731 VP.n49 VSUBS 0.034825f
C1732 VP.n50 VSUBS 0.034825f
C1733 VP.n51 VSUBS 0.048897f
C1734 VP.n52 VSUBS 0.048883f
C1735 VP.n53 VSUBS 0.848135f
C1736 VP.n54 VSUBS 0.048883f
C1737 VP.n55 VSUBS 0.034825f
C1738 VP.n56 VSUBS 0.034825f
C1739 VP.n57 VSUBS 0.034825f
C1740 VP.n58 VSUBS 0.052779f
C1741 VP.n59 VSUBS 0.04632f
C1742 VP.n60 VSUBS 0.848135f
C1743 VP.n61 VSUBS 0.051447f
C1744 VP.n62 VSUBS 0.034825f
C1745 VP.n63 VSUBS 0.034825f
C1746 VP.n64 VSUBS 0.034825f
C1747 VP.n65 VSUBS 0.056661f
C1748 VP.n66 VSUBS 0.043756f
C1749 VP.n67 VSUBS 0.92461f
C1750 VP.n68 VSUBS 0.034644f
.ends

