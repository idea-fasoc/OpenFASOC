* NGSPICE file created from diff_pair_sample_1629.ext - technology: sky130A

.subckt diff_pair_sample_1629 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=2.08
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=5.8422 ps=30.74 w=14.98 l=2.08
X2 VDD2.t0 VN.t1 VTAIL.t2 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=5.8422 ps=30.74 w=14.98 l=2.08
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=5.8422 ps=30.74 w=14.98 l=2.08
X4 B.t8 B.t6 B.t7 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=2.08
X5 B.t5 B.t3 B.t4 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=2.08
X6 B.t2 B.t0 B.t1 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=0 ps=0 w=14.98 l=2.08
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1934_n3964# sky130_fd_pr__pfet_01v8 ad=5.8422 pd=30.74 as=5.8422 ps=30.74 w=14.98 l=2.08
R0 B.n363 B.n362 585
R1 B.n361 B.n96 585
R2 B.n360 B.n359 585
R3 B.n358 B.n97 585
R4 B.n357 B.n356 585
R5 B.n355 B.n98 585
R6 B.n354 B.n353 585
R7 B.n352 B.n99 585
R8 B.n351 B.n350 585
R9 B.n349 B.n100 585
R10 B.n348 B.n347 585
R11 B.n346 B.n101 585
R12 B.n345 B.n344 585
R13 B.n343 B.n102 585
R14 B.n342 B.n341 585
R15 B.n340 B.n103 585
R16 B.n339 B.n338 585
R17 B.n337 B.n104 585
R18 B.n336 B.n335 585
R19 B.n334 B.n105 585
R20 B.n333 B.n332 585
R21 B.n331 B.n106 585
R22 B.n330 B.n329 585
R23 B.n328 B.n107 585
R24 B.n327 B.n326 585
R25 B.n325 B.n108 585
R26 B.n324 B.n323 585
R27 B.n322 B.n109 585
R28 B.n321 B.n320 585
R29 B.n319 B.n110 585
R30 B.n318 B.n317 585
R31 B.n316 B.n111 585
R32 B.n315 B.n314 585
R33 B.n313 B.n112 585
R34 B.n312 B.n311 585
R35 B.n310 B.n113 585
R36 B.n309 B.n308 585
R37 B.n307 B.n114 585
R38 B.n306 B.n305 585
R39 B.n304 B.n115 585
R40 B.n303 B.n302 585
R41 B.n301 B.n116 585
R42 B.n300 B.n299 585
R43 B.n298 B.n117 585
R44 B.n297 B.n296 585
R45 B.n295 B.n118 585
R46 B.n294 B.n293 585
R47 B.n292 B.n119 585
R48 B.n291 B.n290 585
R49 B.n289 B.n120 585
R50 B.n288 B.n287 585
R51 B.n283 B.n121 585
R52 B.n282 B.n281 585
R53 B.n280 B.n122 585
R54 B.n279 B.n278 585
R55 B.n277 B.n123 585
R56 B.n276 B.n275 585
R57 B.n274 B.n124 585
R58 B.n273 B.n272 585
R59 B.n271 B.n125 585
R60 B.n269 B.n268 585
R61 B.n267 B.n128 585
R62 B.n266 B.n265 585
R63 B.n264 B.n129 585
R64 B.n263 B.n262 585
R65 B.n261 B.n130 585
R66 B.n260 B.n259 585
R67 B.n258 B.n131 585
R68 B.n257 B.n256 585
R69 B.n255 B.n132 585
R70 B.n254 B.n253 585
R71 B.n252 B.n133 585
R72 B.n251 B.n250 585
R73 B.n249 B.n134 585
R74 B.n248 B.n247 585
R75 B.n246 B.n135 585
R76 B.n245 B.n244 585
R77 B.n243 B.n136 585
R78 B.n242 B.n241 585
R79 B.n240 B.n137 585
R80 B.n239 B.n238 585
R81 B.n237 B.n138 585
R82 B.n236 B.n235 585
R83 B.n234 B.n139 585
R84 B.n233 B.n232 585
R85 B.n231 B.n140 585
R86 B.n230 B.n229 585
R87 B.n228 B.n141 585
R88 B.n227 B.n226 585
R89 B.n225 B.n142 585
R90 B.n224 B.n223 585
R91 B.n222 B.n143 585
R92 B.n221 B.n220 585
R93 B.n219 B.n144 585
R94 B.n218 B.n217 585
R95 B.n216 B.n145 585
R96 B.n215 B.n214 585
R97 B.n213 B.n146 585
R98 B.n212 B.n211 585
R99 B.n210 B.n147 585
R100 B.n209 B.n208 585
R101 B.n207 B.n148 585
R102 B.n206 B.n205 585
R103 B.n204 B.n149 585
R104 B.n203 B.n202 585
R105 B.n201 B.n150 585
R106 B.n200 B.n199 585
R107 B.n198 B.n151 585
R108 B.n197 B.n196 585
R109 B.n195 B.n152 585
R110 B.n364 B.n95 585
R111 B.n366 B.n365 585
R112 B.n367 B.n94 585
R113 B.n369 B.n368 585
R114 B.n370 B.n93 585
R115 B.n372 B.n371 585
R116 B.n373 B.n92 585
R117 B.n375 B.n374 585
R118 B.n376 B.n91 585
R119 B.n378 B.n377 585
R120 B.n379 B.n90 585
R121 B.n381 B.n380 585
R122 B.n382 B.n89 585
R123 B.n384 B.n383 585
R124 B.n385 B.n88 585
R125 B.n387 B.n386 585
R126 B.n388 B.n87 585
R127 B.n390 B.n389 585
R128 B.n391 B.n86 585
R129 B.n393 B.n392 585
R130 B.n394 B.n85 585
R131 B.n396 B.n395 585
R132 B.n397 B.n84 585
R133 B.n399 B.n398 585
R134 B.n400 B.n83 585
R135 B.n402 B.n401 585
R136 B.n403 B.n82 585
R137 B.n405 B.n404 585
R138 B.n406 B.n81 585
R139 B.n408 B.n407 585
R140 B.n409 B.n80 585
R141 B.n411 B.n410 585
R142 B.n412 B.n79 585
R143 B.n414 B.n413 585
R144 B.n415 B.n78 585
R145 B.n417 B.n416 585
R146 B.n418 B.n77 585
R147 B.n420 B.n419 585
R148 B.n421 B.n76 585
R149 B.n423 B.n422 585
R150 B.n424 B.n75 585
R151 B.n426 B.n425 585
R152 B.n427 B.n74 585
R153 B.n429 B.n428 585
R154 B.n430 B.n73 585
R155 B.n432 B.n431 585
R156 B.n598 B.n13 585
R157 B.n597 B.n596 585
R158 B.n595 B.n14 585
R159 B.n594 B.n593 585
R160 B.n592 B.n15 585
R161 B.n591 B.n590 585
R162 B.n589 B.n16 585
R163 B.n588 B.n587 585
R164 B.n586 B.n17 585
R165 B.n585 B.n584 585
R166 B.n583 B.n18 585
R167 B.n582 B.n581 585
R168 B.n580 B.n19 585
R169 B.n579 B.n578 585
R170 B.n577 B.n20 585
R171 B.n576 B.n575 585
R172 B.n574 B.n21 585
R173 B.n573 B.n572 585
R174 B.n571 B.n22 585
R175 B.n570 B.n569 585
R176 B.n568 B.n23 585
R177 B.n567 B.n566 585
R178 B.n565 B.n24 585
R179 B.n564 B.n563 585
R180 B.n562 B.n25 585
R181 B.n561 B.n560 585
R182 B.n559 B.n26 585
R183 B.n558 B.n557 585
R184 B.n556 B.n27 585
R185 B.n555 B.n554 585
R186 B.n553 B.n28 585
R187 B.n552 B.n551 585
R188 B.n550 B.n29 585
R189 B.n549 B.n548 585
R190 B.n547 B.n30 585
R191 B.n546 B.n545 585
R192 B.n544 B.n31 585
R193 B.n543 B.n542 585
R194 B.n541 B.n32 585
R195 B.n540 B.n539 585
R196 B.n538 B.n33 585
R197 B.n537 B.n536 585
R198 B.n535 B.n34 585
R199 B.n534 B.n533 585
R200 B.n532 B.n35 585
R201 B.n531 B.n530 585
R202 B.n529 B.n36 585
R203 B.n528 B.n527 585
R204 B.n526 B.n37 585
R205 B.n525 B.n524 585
R206 B.n523 B.n522 585
R207 B.n521 B.n41 585
R208 B.n520 B.n519 585
R209 B.n518 B.n42 585
R210 B.n517 B.n516 585
R211 B.n515 B.n43 585
R212 B.n514 B.n513 585
R213 B.n512 B.n44 585
R214 B.n511 B.n510 585
R215 B.n509 B.n45 585
R216 B.n507 B.n506 585
R217 B.n505 B.n48 585
R218 B.n504 B.n503 585
R219 B.n502 B.n49 585
R220 B.n501 B.n500 585
R221 B.n499 B.n50 585
R222 B.n498 B.n497 585
R223 B.n496 B.n51 585
R224 B.n495 B.n494 585
R225 B.n493 B.n52 585
R226 B.n492 B.n491 585
R227 B.n490 B.n53 585
R228 B.n489 B.n488 585
R229 B.n487 B.n54 585
R230 B.n486 B.n485 585
R231 B.n484 B.n55 585
R232 B.n483 B.n482 585
R233 B.n481 B.n56 585
R234 B.n480 B.n479 585
R235 B.n478 B.n57 585
R236 B.n477 B.n476 585
R237 B.n475 B.n58 585
R238 B.n474 B.n473 585
R239 B.n472 B.n59 585
R240 B.n471 B.n470 585
R241 B.n469 B.n60 585
R242 B.n468 B.n467 585
R243 B.n466 B.n61 585
R244 B.n465 B.n464 585
R245 B.n463 B.n62 585
R246 B.n462 B.n461 585
R247 B.n460 B.n63 585
R248 B.n459 B.n458 585
R249 B.n457 B.n64 585
R250 B.n456 B.n455 585
R251 B.n454 B.n65 585
R252 B.n453 B.n452 585
R253 B.n451 B.n66 585
R254 B.n450 B.n449 585
R255 B.n448 B.n67 585
R256 B.n447 B.n446 585
R257 B.n445 B.n68 585
R258 B.n444 B.n443 585
R259 B.n442 B.n69 585
R260 B.n441 B.n440 585
R261 B.n439 B.n70 585
R262 B.n438 B.n437 585
R263 B.n436 B.n71 585
R264 B.n435 B.n434 585
R265 B.n433 B.n72 585
R266 B.n600 B.n599 585
R267 B.n601 B.n12 585
R268 B.n603 B.n602 585
R269 B.n604 B.n11 585
R270 B.n606 B.n605 585
R271 B.n607 B.n10 585
R272 B.n609 B.n608 585
R273 B.n610 B.n9 585
R274 B.n612 B.n611 585
R275 B.n613 B.n8 585
R276 B.n615 B.n614 585
R277 B.n616 B.n7 585
R278 B.n618 B.n617 585
R279 B.n619 B.n6 585
R280 B.n621 B.n620 585
R281 B.n622 B.n5 585
R282 B.n624 B.n623 585
R283 B.n625 B.n4 585
R284 B.n627 B.n626 585
R285 B.n628 B.n3 585
R286 B.n630 B.n629 585
R287 B.n631 B.n0 585
R288 B.n2 B.n1 585
R289 B.n164 B.n163 585
R290 B.n165 B.n162 585
R291 B.n167 B.n166 585
R292 B.n168 B.n161 585
R293 B.n170 B.n169 585
R294 B.n171 B.n160 585
R295 B.n173 B.n172 585
R296 B.n174 B.n159 585
R297 B.n176 B.n175 585
R298 B.n177 B.n158 585
R299 B.n179 B.n178 585
R300 B.n180 B.n157 585
R301 B.n182 B.n181 585
R302 B.n183 B.n156 585
R303 B.n185 B.n184 585
R304 B.n186 B.n155 585
R305 B.n188 B.n187 585
R306 B.n189 B.n154 585
R307 B.n191 B.n190 585
R308 B.n192 B.n153 585
R309 B.n194 B.n193 585
R310 B.n195 B.n194 492.5
R311 B.n362 B.n95 492.5
R312 B.n433 B.n432 492.5
R313 B.n600 B.n13 492.5
R314 B.n126 B.t3 380.666
R315 B.n284 B.t6 380.666
R316 B.n46 B.t0 380.666
R317 B.n38 B.t9 380.666
R318 B.n633 B.n632 256.663
R319 B.n632 B.n631 235.042
R320 B.n632 B.n2 235.042
R321 B.n196 B.n195 163.367
R322 B.n196 B.n151 163.367
R323 B.n200 B.n151 163.367
R324 B.n201 B.n200 163.367
R325 B.n202 B.n201 163.367
R326 B.n202 B.n149 163.367
R327 B.n206 B.n149 163.367
R328 B.n207 B.n206 163.367
R329 B.n208 B.n207 163.367
R330 B.n208 B.n147 163.367
R331 B.n212 B.n147 163.367
R332 B.n213 B.n212 163.367
R333 B.n214 B.n213 163.367
R334 B.n214 B.n145 163.367
R335 B.n218 B.n145 163.367
R336 B.n219 B.n218 163.367
R337 B.n220 B.n219 163.367
R338 B.n220 B.n143 163.367
R339 B.n224 B.n143 163.367
R340 B.n225 B.n224 163.367
R341 B.n226 B.n225 163.367
R342 B.n226 B.n141 163.367
R343 B.n230 B.n141 163.367
R344 B.n231 B.n230 163.367
R345 B.n232 B.n231 163.367
R346 B.n232 B.n139 163.367
R347 B.n236 B.n139 163.367
R348 B.n237 B.n236 163.367
R349 B.n238 B.n237 163.367
R350 B.n238 B.n137 163.367
R351 B.n242 B.n137 163.367
R352 B.n243 B.n242 163.367
R353 B.n244 B.n243 163.367
R354 B.n244 B.n135 163.367
R355 B.n248 B.n135 163.367
R356 B.n249 B.n248 163.367
R357 B.n250 B.n249 163.367
R358 B.n250 B.n133 163.367
R359 B.n254 B.n133 163.367
R360 B.n255 B.n254 163.367
R361 B.n256 B.n255 163.367
R362 B.n256 B.n131 163.367
R363 B.n260 B.n131 163.367
R364 B.n261 B.n260 163.367
R365 B.n262 B.n261 163.367
R366 B.n262 B.n129 163.367
R367 B.n266 B.n129 163.367
R368 B.n267 B.n266 163.367
R369 B.n268 B.n267 163.367
R370 B.n268 B.n125 163.367
R371 B.n273 B.n125 163.367
R372 B.n274 B.n273 163.367
R373 B.n275 B.n274 163.367
R374 B.n275 B.n123 163.367
R375 B.n279 B.n123 163.367
R376 B.n280 B.n279 163.367
R377 B.n281 B.n280 163.367
R378 B.n281 B.n121 163.367
R379 B.n288 B.n121 163.367
R380 B.n289 B.n288 163.367
R381 B.n290 B.n289 163.367
R382 B.n290 B.n119 163.367
R383 B.n294 B.n119 163.367
R384 B.n295 B.n294 163.367
R385 B.n296 B.n295 163.367
R386 B.n296 B.n117 163.367
R387 B.n300 B.n117 163.367
R388 B.n301 B.n300 163.367
R389 B.n302 B.n301 163.367
R390 B.n302 B.n115 163.367
R391 B.n306 B.n115 163.367
R392 B.n307 B.n306 163.367
R393 B.n308 B.n307 163.367
R394 B.n308 B.n113 163.367
R395 B.n312 B.n113 163.367
R396 B.n313 B.n312 163.367
R397 B.n314 B.n313 163.367
R398 B.n314 B.n111 163.367
R399 B.n318 B.n111 163.367
R400 B.n319 B.n318 163.367
R401 B.n320 B.n319 163.367
R402 B.n320 B.n109 163.367
R403 B.n324 B.n109 163.367
R404 B.n325 B.n324 163.367
R405 B.n326 B.n325 163.367
R406 B.n326 B.n107 163.367
R407 B.n330 B.n107 163.367
R408 B.n331 B.n330 163.367
R409 B.n332 B.n331 163.367
R410 B.n332 B.n105 163.367
R411 B.n336 B.n105 163.367
R412 B.n337 B.n336 163.367
R413 B.n338 B.n337 163.367
R414 B.n338 B.n103 163.367
R415 B.n342 B.n103 163.367
R416 B.n343 B.n342 163.367
R417 B.n344 B.n343 163.367
R418 B.n344 B.n101 163.367
R419 B.n348 B.n101 163.367
R420 B.n349 B.n348 163.367
R421 B.n350 B.n349 163.367
R422 B.n350 B.n99 163.367
R423 B.n354 B.n99 163.367
R424 B.n355 B.n354 163.367
R425 B.n356 B.n355 163.367
R426 B.n356 B.n97 163.367
R427 B.n360 B.n97 163.367
R428 B.n361 B.n360 163.367
R429 B.n362 B.n361 163.367
R430 B.n432 B.n73 163.367
R431 B.n428 B.n73 163.367
R432 B.n428 B.n427 163.367
R433 B.n427 B.n426 163.367
R434 B.n426 B.n75 163.367
R435 B.n422 B.n75 163.367
R436 B.n422 B.n421 163.367
R437 B.n421 B.n420 163.367
R438 B.n420 B.n77 163.367
R439 B.n416 B.n77 163.367
R440 B.n416 B.n415 163.367
R441 B.n415 B.n414 163.367
R442 B.n414 B.n79 163.367
R443 B.n410 B.n79 163.367
R444 B.n410 B.n409 163.367
R445 B.n409 B.n408 163.367
R446 B.n408 B.n81 163.367
R447 B.n404 B.n81 163.367
R448 B.n404 B.n403 163.367
R449 B.n403 B.n402 163.367
R450 B.n402 B.n83 163.367
R451 B.n398 B.n83 163.367
R452 B.n398 B.n397 163.367
R453 B.n397 B.n396 163.367
R454 B.n396 B.n85 163.367
R455 B.n392 B.n85 163.367
R456 B.n392 B.n391 163.367
R457 B.n391 B.n390 163.367
R458 B.n390 B.n87 163.367
R459 B.n386 B.n87 163.367
R460 B.n386 B.n385 163.367
R461 B.n385 B.n384 163.367
R462 B.n384 B.n89 163.367
R463 B.n380 B.n89 163.367
R464 B.n380 B.n379 163.367
R465 B.n379 B.n378 163.367
R466 B.n378 B.n91 163.367
R467 B.n374 B.n91 163.367
R468 B.n374 B.n373 163.367
R469 B.n373 B.n372 163.367
R470 B.n372 B.n93 163.367
R471 B.n368 B.n93 163.367
R472 B.n368 B.n367 163.367
R473 B.n367 B.n366 163.367
R474 B.n366 B.n95 163.367
R475 B.n596 B.n13 163.367
R476 B.n596 B.n595 163.367
R477 B.n595 B.n594 163.367
R478 B.n594 B.n15 163.367
R479 B.n590 B.n15 163.367
R480 B.n590 B.n589 163.367
R481 B.n589 B.n588 163.367
R482 B.n588 B.n17 163.367
R483 B.n584 B.n17 163.367
R484 B.n584 B.n583 163.367
R485 B.n583 B.n582 163.367
R486 B.n582 B.n19 163.367
R487 B.n578 B.n19 163.367
R488 B.n578 B.n577 163.367
R489 B.n577 B.n576 163.367
R490 B.n576 B.n21 163.367
R491 B.n572 B.n21 163.367
R492 B.n572 B.n571 163.367
R493 B.n571 B.n570 163.367
R494 B.n570 B.n23 163.367
R495 B.n566 B.n23 163.367
R496 B.n566 B.n565 163.367
R497 B.n565 B.n564 163.367
R498 B.n564 B.n25 163.367
R499 B.n560 B.n25 163.367
R500 B.n560 B.n559 163.367
R501 B.n559 B.n558 163.367
R502 B.n558 B.n27 163.367
R503 B.n554 B.n27 163.367
R504 B.n554 B.n553 163.367
R505 B.n553 B.n552 163.367
R506 B.n552 B.n29 163.367
R507 B.n548 B.n29 163.367
R508 B.n548 B.n547 163.367
R509 B.n547 B.n546 163.367
R510 B.n546 B.n31 163.367
R511 B.n542 B.n31 163.367
R512 B.n542 B.n541 163.367
R513 B.n541 B.n540 163.367
R514 B.n540 B.n33 163.367
R515 B.n536 B.n33 163.367
R516 B.n536 B.n535 163.367
R517 B.n535 B.n534 163.367
R518 B.n534 B.n35 163.367
R519 B.n530 B.n35 163.367
R520 B.n530 B.n529 163.367
R521 B.n529 B.n528 163.367
R522 B.n528 B.n37 163.367
R523 B.n524 B.n37 163.367
R524 B.n524 B.n523 163.367
R525 B.n523 B.n41 163.367
R526 B.n519 B.n41 163.367
R527 B.n519 B.n518 163.367
R528 B.n518 B.n517 163.367
R529 B.n517 B.n43 163.367
R530 B.n513 B.n43 163.367
R531 B.n513 B.n512 163.367
R532 B.n512 B.n511 163.367
R533 B.n511 B.n45 163.367
R534 B.n506 B.n45 163.367
R535 B.n506 B.n505 163.367
R536 B.n505 B.n504 163.367
R537 B.n504 B.n49 163.367
R538 B.n500 B.n49 163.367
R539 B.n500 B.n499 163.367
R540 B.n499 B.n498 163.367
R541 B.n498 B.n51 163.367
R542 B.n494 B.n51 163.367
R543 B.n494 B.n493 163.367
R544 B.n493 B.n492 163.367
R545 B.n492 B.n53 163.367
R546 B.n488 B.n53 163.367
R547 B.n488 B.n487 163.367
R548 B.n487 B.n486 163.367
R549 B.n486 B.n55 163.367
R550 B.n482 B.n55 163.367
R551 B.n482 B.n481 163.367
R552 B.n481 B.n480 163.367
R553 B.n480 B.n57 163.367
R554 B.n476 B.n57 163.367
R555 B.n476 B.n475 163.367
R556 B.n475 B.n474 163.367
R557 B.n474 B.n59 163.367
R558 B.n470 B.n59 163.367
R559 B.n470 B.n469 163.367
R560 B.n469 B.n468 163.367
R561 B.n468 B.n61 163.367
R562 B.n464 B.n61 163.367
R563 B.n464 B.n463 163.367
R564 B.n463 B.n462 163.367
R565 B.n462 B.n63 163.367
R566 B.n458 B.n63 163.367
R567 B.n458 B.n457 163.367
R568 B.n457 B.n456 163.367
R569 B.n456 B.n65 163.367
R570 B.n452 B.n65 163.367
R571 B.n452 B.n451 163.367
R572 B.n451 B.n450 163.367
R573 B.n450 B.n67 163.367
R574 B.n446 B.n67 163.367
R575 B.n446 B.n445 163.367
R576 B.n445 B.n444 163.367
R577 B.n444 B.n69 163.367
R578 B.n440 B.n69 163.367
R579 B.n440 B.n439 163.367
R580 B.n439 B.n438 163.367
R581 B.n438 B.n71 163.367
R582 B.n434 B.n71 163.367
R583 B.n434 B.n433 163.367
R584 B.n601 B.n600 163.367
R585 B.n602 B.n601 163.367
R586 B.n602 B.n11 163.367
R587 B.n606 B.n11 163.367
R588 B.n607 B.n606 163.367
R589 B.n608 B.n607 163.367
R590 B.n608 B.n9 163.367
R591 B.n612 B.n9 163.367
R592 B.n613 B.n612 163.367
R593 B.n614 B.n613 163.367
R594 B.n614 B.n7 163.367
R595 B.n618 B.n7 163.367
R596 B.n619 B.n618 163.367
R597 B.n620 B.n619 163.367
R598 B.n620 B.n5 163.367
R599 B.n624 B.n5 163.367
R600 B.n625 B.n624 163.367
R601 B.n626 B.n625 163.367
R602 B.n626 B.n3 163.367
R603 B.n630 B.n3 163.367
R604 B.n631 B.n630 163.367
R605 B.n164 B.n2 163.367
R606 B.n165 B.n164 163.367
R607 B.n166 B.n165 163.367
R608 B.n166 B.n161 163.367
R609 B.n170 B.n161 163.367
R610 B.n171 B.n170 163.367
R611 B.n172 B.n171 163.367
R612 B.n172 B.n159 163.367
R613 B.n176 B.n159 163.367
R614 B.n177 B.n176 163.367
R615 B.n178 B.n177 163.367
R616 B.n178 B.n157 163.367
R617 B.n182 B.n157 163.367
R618 B.n183 B.n182 163.367
R619 B.n184 B.n183 163.367
R620 B.n184 B.n155 163.367
R621 B.n188 B.n155 163.367
R622 B.n189 B.n188 163.367
R623 B.n190 B.n189 163.367
R624 B.n190 B.n153 163.367
R625 B.n194 B.n153 163.367
R626 B.n284 B.t7 153.691
R627 B.n46 B.t2 153.691
R628 B.n126 B.t4 153.673
R629 B.n38 B.t11 153.673
R630 B.n285 B.t8 106.953
R631 B.n47 B.t1 106.953
R632 B.n127 B.t5 106.933
R633 B.n39 B.t10 106.933
R634 B.n270 B.n127 59.5399
R635 B.n286 B.n285 59.5399
R636 B.n508 B.n47 59.5399
R637 B.n40 B.n39 59.5399
R638 B.n127 B.n126 46.7399
R639 B.n285 B.n284 46.7399
R640 B.n47 B.n46 46.7399
R641 B.n39 B.n38 46.7399
R642 B.n599 B.n598 32.0005
R643 B.n431 B.n72 32.0005
R644 B.n364 B.n363 32.0005
R645 B.n193 B.n152 32.0005
R646 B B.n633 18.0485
R647 B.n599 B.n12 10.6151
R648 B.n603 B.n12 10.6151
R649 B.n604 B.n603 10.6151
R650 B.n605 B.n604 10.6151
R651 B.n605 B.n10 10.6151
R652 B.n609 B.n10 10.6151
R653 B.n610 B.n609 10.6151
R654 B.n611 B.n610 10.6151
R655 B.n611 B.n8 10.6151
R656 B.n615 B.n8 10.6151
R657 B.n616 B.n615 10.6151
R658 B.n617 B.n616 10.6151
R659 B.n617 B.n6 10.6151
R660 B.n621 B.n6 10.6151
R661 B.n622 B.n621 10.6151
R662 B.n623 B.n622 10.6151
R663 B.n623 B.n4 10.6151
R664 B.n627 B.n4 10.6151
R665 B.n628 B.n627 10.6151
R666 B.n629 B.n628 10.6151
R667 B.n629 B.n0 10.6151
R668 B.n598 B.n597 10.6151
R669 B.n597 B.n14 10.6151
R670 B.n593 B.n14 10.6151
R671 B.n593 B.n592 10.6151
R672 B.n592 B.n591 10.6151
R673 B.n591 B.n16 10.6151
R674 B.n587 B.n16 10.6151
R675 B.n587 B.n586 10.6151
R676 B.n586 B.n585 10.6151
R677 B.n585 B.n18 10.6151
R678 B.n581 B.n18 10.6151
R679 B.n581 B.n580 10.6151
R680 B.n580 B.n579 10.6151
R681 B.n579 B.n20 10.6151
R682 B.n575 B.n20 10.6151
R683 B.n575 B.n574 10.6151
R684 B.n574 B.n573 10.6151
R685 B.n573 B.n22 10.6151
R686 B.n569 B.n22 10.6151
R687 B.n569 B.n568 10.6151
R688 B.n568 B.n567 10.6151
R689 B.n567 B.n24 10.6151
R690 B.n563 B.n24 10.6151
R691 B.n563 B.n562 10.6151
R692 B.n562 B.n561 10.6151
R693 B.n561 B.n26 10.6151
R694 B.n557 B.n26 10.6151
R695 B.n557 B.n556 10.6151
R696 B.n556 B.n555 10.6151
R697 B.n555 B.n28 10.6151
R698 B.n551 B.n28 10.6151
R699 B.n551 B.n550 10.6151
R700 B.n550 B.n549 10.6151
R701 B.n549 B.n30 10.6151
R702 B.n545 B.n30 10.6151
R703 B.n545 B.n544 10.6151
R704 B.n544 B.n543 10.6151
R705 B.n543 B.n32 10.6151
R706 B.n539 B.n32 10.6151
R707 B.n539 B.n538 10.6151
R708 B.n538 B.n537 10.6151
R709 B.n537 B.n34 10.6151
R710 B.n533 B.n34 10.6151
R711 B.n533 B.n532 10.6151
R712 B.n532 B.n531 10.6151
R713 B.n531 B.n36 10.6151
R714 B.n527 B.n36 10.6151
R715 B.n527 B.n526 10.6151
R716 B.n526 B.n525 10.6151
R717 B.n522 B.n521 10.6151
R718 B.n521 B.n520 10.6151
R719 B.n520 B.n42 10.6151
R720 B.n516 B.n42 10.6151
R721 B.n516 B.n515 10.6151
R722 B.n515 B.n514 10.6151
R723 B.n514 B.n44 10.6151
R724 B.n510 B.n44 10.6151
R725 B.n510 B.n509 10.6151
R726 B.n507 B.n48 10.6151
R727 B.n503 B.n48 10.6151
R728 B.n503 B.n502 10.6151
R729 B.n502 B.n501 10.6151
R730 B.n501 B.n50 10.6151
R731 B.n497 B.n50 10.6151
R732 B.n497 B.n496 10.6151
R733 B.n496 B.n495 10.6151
R734 B.n495 B.n52 10.6151
R735 B.n491 B.n52 10.6151
R736 B.n491 B.n490 10.6151
R737 B.n490 B.n489 10.6151
R738 B.n489 B.n54 10.6151
R739 B.n485 B.n54 10.6151
R740 B.n485 B.n484 10.6151
R741 B.n484 B.n483 10.6151
R742 B.n483 B.n56 10.6151
R743 B.n479 B.n56 10.6151
R744 B.n479 B.n478 10.6151
R745 B.n478 B.n477 10.6151
R746 B.n477 B.n58 10.6151
R747 B.n473 B.n58 10.6151
R748 B.n473 B.n472 10.6151
R749 B.n472 B.n471 10.6151
R750 B.n471 B.n60 10.6151
R751 B.n467 B.n60 10.6151
R752 B.n467 B.n466 10.6151
R753 B.n466 B.n465 10.6151
R754 B.n465 B.n62 10.6151
R755 B.n461 B.n62 10.6151
R756 B.n461 B.n460 10.6151
R757 B.n460 B.n459 10.6151
R758 B.n459 B.n64 10.6151
R759 B.n455 B.n64 10.6151
R760 B.n455 B.n454 10.6151
R761 B.n454 B.n453 10.6151
R762 B.n453 B.n66 10.6151
R763 B.n449 B.n66 10.6151
R764 B.n449 B.n448 10.6151
R765 B.n448 B.n447 10.6151
R766 B.n447 B.n68 10.6151
R767 B.n443 B.n68 10.6151
R768 B.n443 B.n442 10.6151
R769 B.n442 B.n441 10.6151
R770 B.n441 B.n70 10.6151
R771 B.n437 B.n70 10.6151
R772 B.n437 B.n436 10.6151
R773 B.n436 B.n435 10.6151
R774 B.n435 B.n72 10.6151
R775 B.n431 B.n430 10.6151
R776 B.n430 B.n429 10.6151
R777 B.n429 B.n74 10.6151
R778 B.n425 B.n74 10.6151
R779 B.n425 B.n424 10.6151
R780 B.n424 B.n423 10.6151
R781 B.n423 B.n76 10.6151
R782 B.n419 B.n76 10.6151
R783 B.n419 B.n418 10.6151
R784 B.n418 B.n417 10.6151
R785 B.n417 B.n78 10.6151
R786 B.n413 B.n78 10.6151
R787 B.n413 B.n412 10.6151
R788 B.n412 B.n411 10.6151
R789 B.n411 B.n80 10.6151
R790 B.n407 B.n80 10.6151
R791 B.n407 B.n406 10.6151
R792 B.n406 B.n405 10.6151
R793 B.n405 B.n82 10.6151
R794 B.n401 B.n82 10.6151
R795 B.n401 B.n400 10.6151
R796 B.n400 B.n399 10.6151
R797 B.n399 B.n84 10.6151
R798 B.n395 B.n84 10.6151
R799 B.n395 B.n394 10.6151
R800 B.n394 B.n393 10.6151
R801 B.n393 B.n86 10.6151
R802 B.n389 B.n86 10.6151
R803 B.n389 B.n388 10.6151
R804 B.n388 B.n387 10.6151
R805 B.n387 B.n88 10.6151
R806 B.n383 B.n88 10.6151
R807 B.n383 B.n382 10.6151
R808 B.n382 B.n381 10.6151
R809 B.n381 B.n90 10.6151
R810 B.n377 B.n90 10.6151
R811 B.n377 B.n376 10.6151
R812 B.n376 B.n375 10.6151
R813 B.n375 B.n92 10.6151
R814 B.n371 B.n92 10.6151
R815 B.n371 B.n370 10.6151
R816 B.n370 B.n369 10.6151
R817 B.n369 B.n94 10.6151
R818 B.n365 B.n94 10.6151
R819 B.n365 B.n364 10.6151
R820 B.n163 B.n1 10.6151
R821 B.n163 B.n162 10.6151
R822 B.n167 B.n162 10.6151
R823 B.n168 B.n167 10.6151
R824 B.n169 B.n168 10.6151
R825 B.n169 B.n160 10.6151
R826 B.n173 B.n160 10.6151
R827 B.n174 B.n173 10.6151
R828 B.n175 B.n174 10.6151
R829 B.n175 B.n158 10.6151
R830 B.n179 B.n158 10.6151
R831 B.n180 B.n179 10.6151
R832 B.n181 B.n180 10.6151
R833 B.n181 B.n156 10.6151
R834 B.n185 B.n156 10.6151
R835 B.n186 B.n185 10.6151
R836 B.n187 B.n186 10.6151
R837 B.n187 B.n154 10.6151
R838 B.n191 B.n154 10.6151
R839 B.n192 B.n191 10.6151
R840 B.n193 B.n192 10.6151
R841 B.n197 B.n152 10.6151
R842 B.n198 B.n197 10.6151
R843 B.n199 B.n198 10.6151
R844 B.n199 B.n150 10.6151
R845 B.n203 B.n150 10.6151
R846 B.n204 B.n203 10.6151
R847 B.n205 B.n204 10.6151
R848 B.n205 B.n148 10.6151
R849 B.n209 B.n148 10.6151
R850 B.n210 B.n209 10.6151
R851 B.n211 B.n210 10.6151
R852 B.n211 B.n146 10.6151
R853 B.n215 B.n146 10.6151
R854 B.n216 B.n215 10.6151
R855 B.n217 B.n216 10.6151
R856 B.n217 B.n144 10.6151
R857 B.n221 B.n144 10.6151
R858 B.n222 B.n221 10.6151
R859 B.n223 B.n222 10.6151
R860 B.n223 B.n142 10.6151
R861 B.n227 B.n142 10.6151
R862 B.n228 B.n227 10.6151
R863 B.n229 B.n228 10.6151
R864 B.n229 B.n140 10.6151
R865 B.n233 B.n140 10.6151
R866 B.n234 B.n233 10.6151
R867 B.n235 B.n234 10.6151
R868 B.n235 B.n138 10.6151
R869 B.n239 B.n138 10.6151
R870 B.n240 B.n239 10.6151
R871 B.n241 B.n240 10.6151
R872 B.n241 B.n136 10.6151
R873 B.n245 B.n136 10.6151
R874 B.n246 B.n245 10.6151
R875 B.n247 B.n246 10.6151
R876 B.n247 B.n134 10.6151
R877 B.n251 B.n134 10.6151
R878 B.n252 B.n251 10.6151
R879 B.n253 B.n252 10.6151
R880 B.n253 B.n132 10.6151
R881 B.n257 B.n132 10.6151
R882 B.n258 B.n257 10.6151
R883 B.n259 B.n258 10.6151
R884 B.n259 B.n130 10.6151
R885 B.n263 B.n130 10.6151
R886 B.n264 B.n263 10.6151
R887 B.n265 B.n264 10.6151
R888 B.n265 B.n128 10.6151
R889 B.n269 B.n128 10.6151
R890 B.n272 B.n271 10.6151
R891 B.n272 B.n124 10.6151
R892 B.n276 B.n124 10.6151
R893 B.n277 B.n276 10.6151
R894 B.n278 B.n277 10.6151
R895 B.n278 B.n122 10.6151
R896 B.n282 B.n122 10.6151
R897 B.n283 B.n282 10.6151
R898 B.n287 B.n283 10.6151
R899 B.n291 B.n120 10.6151
R900 B.n292 B.n291 10.6151
R901 B.n293 B.n292 10.6151
R902 B.n293 B.n118 10.6151
R903 B.n297 B.n118 10.6151
R904 B.n298 B.n297 10.6151
R905 B.n299 B.n298 10.6151
R906 B.n299 B.n116 10.6151
R907 B.n303 B.n116 10.6151
R908 B.n304 B.n303 10.6151
R909 B.n305 B.n304 10.6151
R910 B.n305 B.n114 10.6151
R911 B.n309 B.n114 10.6151
R912 B.n310 B.n309 10.6151
R913 B.n311 B.n310 10.6151
R914 B.n311 B.n112 10.6151
R915 B.n315 B.n112 10.6151
R916 B.n316 B.n315 10.6151
R917 B.n317 B.n316 10.6151
R918 B.n317 B.n110 10.6151
R919 B.n321 B.n110 10.6151
R920 B.n322 B.n321 10.6151
R921 B.n323 B.n322 10.6151
R922 B.n323 B.n108 10.6151
R923 B.n327 B.n108 10.6151
R924 B.n328 B.n327 10.6151
R925 B.n329 B.n328 10.6151
R926 B.n329 B.n106 10.6151
R927 B.n333 B.n106 10.6151
R928 B.n334 B.n333 10.6151
R929 B.n335 B.n334 10.6151
R930 B.n335 B.n104 10.6151
R931 B.n339 B.n104 10.6151
R932 B.n340 B.n339 10.6151
R933 B.n341 B.n340 10.6151
R934 B.n341 B.n102 10.6151
R935 B.n345 B.n102 10.6151
R936 B.n346 B.n345 10.6151
R937 B.n347 B.n346 10.6151
R938 B.n347 B.n100 10.6151
R939 B.n351 B.n100 10.6151
R940 B.n352 B.n351 10.6151
R941 B.n353 B.n352 10.6151
R942 B.n353 B.n98 10.6151
R943 B.n357 B.n98 10.6151
R944 B.n358 B.n357 10.6151
R945 B.n359 B.n358 10.6151
R946 B.n359 B.n96 10.6151
R947 B.n363 B.n96 10.6151
R948 B.n525 B.n40 9.36635
R949 B.n508 B.n507 9.36635
R950 B.n270 B.n269 9.36635
R951 B.n286 B.n120 9.36635
R952 B.n633 B.n0 8.11757
R953 B.n633 B.n1 8.11757
R954 B.n522 B.n40 1.24928
R955 B.n509 B.n508 1.24928
R956 B.n271 B.n270 1.24928
R957 B.n287 B.n286 1.24928
R958 VN VN.t1 278.178
R959 VN VN.t0 232.694
R960 VTAIL.n1 VTAIL.t2 55.6084
R961 VTAIL.n3 VTAIL.t3 55.6081
R962 VTAIL.n0 VTAIL.t1 55.6081
R963 VTAIL.n2 VTAIL.t0 55.6081
R964 VTAIL.n1 VTAIL.n0 29.4358
R965 VTAIL.n3 VTAIL.n2 27.3583
R966 VTAIL.n2 VTAIL.n1 1.50912
R967 VTAIL VTAIL.n0 1.04791
R968 VTAIL VTAIL.n3 0.461707
R969 VDD2.n0 VDD2.t1 113.016
R970 VDD2.n0 VDD2.t0 72.2869
R971 VDD2 VDD2.n0 0.578086
R972 VP.n0 VP.t1 277.988
R973 VP.n0 VP.t0 232.452
R974 VP VP.n0 0.241678
R975 VDD1 VDD1.t1 114.059
R976 VDD1 VDD1.t0 72.8645
C0 VTAIL VP 2.78557f
C1 VDD1 VDD2 0.613146f
C2 VTAIL VN 2.77118f
C3 B w_n1934_n3964# 9.08333f
C4 VN VP 5.75723f
C5 VTAIL w_n1934_n3964# 3.20738f
C6 VDD2 B 1.8919f
C7 VDD1 B 1.86643f
C8 w_n1934_n3964# VP 2.91775f
C9 VN w_n1934_n3964# 2.67252f
C10 VTAIL VDD2 5.88797f
C11 VTAIL VDD1 5.84234f
C12 VDD2 VP 0.311872f
C13 VDD1 VP 3.44122f
C14 VN VDD2 3.28103f
C15 VN VDD1 0.148217f
C16 VTAIL B 4.0776f
C17 B VP 1.40149f
C18 VDD2 w_n1934_n3964# 1.95201f
C19 VDD1 w_n1934_n3964# 1.93236f
C20 VN B 1.00041f
C21 VDD2 VSUBS 0.940346f
C22 VDD1 VSUBS 4.62703f
C23 VTAIL VSUBS 1.053977f
C24 VN VSUBS 8.36613f
C25 VP VSUBS 1.637656f
C26 B VSUBS 3.757024f
C27 w_n1934_n3964# VSUBS 94.0156f
C28 VDD1.t0 VSUBS 2.49187f
C29 VDD1.t1 VSUBS 3.14957f
C30 VP.t1 VSUBS 4.65289f
C31 VP.t0 VSUBS 4.10833f
C32 VP.n0 VSUBS 6.06279f
C33 VDD2.t1 VSUBS 3.14145f
C34 VDD2.t0 VSUBS 2.508f
C35 VDD2.n0 VSUBS 3.44527f
C36 VTAIL.t1 VSUBS 3.35568f
C37 VTAIL.n0 VSUBS 2.84726f
C38 VTAIL.t2 VSUBS 3.35568f
C39 VTAIL.n1 VSUBS 2.88953f
C40 VTAIL.t0 VSUBS 3.35568f
C41 VTAIL.n2 VSUBS 2.69911f
C42 VTAIL.t3 VSUBS 3.35568f
C43 VTAIL.n3 VSUBS 2.60311f
C44 VN.t0 VSUBS 4.01047f
C45 VN.t1 VSUBS 4.54559f
C46 B.n0 VSUBS 0.005278f
C47 B.n1 VSUBS 0.005278f
C48 B.n2 VSUBS 0.007806f
C49 B.n3 VSUBS 0.005982f
C50 B.n4 VSUBS 0.005982f
C51 B.n5 VSUBS 0.005982f
C52 B.n6 VSUBS 0.005982f
C53 B.n7 VSUBS 0.005982f
C54 B.n8 VSUBS 0.005982f
C55 B.n9 VSUBS 0.005982f
C56 B.n10 VSUBS 0.005982f
C57 B.n11 VSUBS 0.005982f
C58 B.n12 VSUBS 0.005982f
C59 B.n13 VSUBS 0.013926f
C60 B.n14 VSUBS 0.005982f
C61 B.n15 VSUBS 0.005982f
C62 B.n16 VSUBS 0.005982f
C63 B.n17 VSUBS 0.005982f
C64 B.n18 VSUBS 0.005982f
C65 B.n19 VSUBS 0.005982f
C66 B.n20 VSUBS 0.005982f
C67 B.n21 VSUBS 0.005982f
C68 B.n22 VSUBS 0.005982f
C69 B.n23 VSUBS 0.005982f
C70 B.n24 VSUBS 0.005982f
C71 B.n25 VSUBS 0.005982f
C72 B.n26 VSUBS 0.005982f
C73 B.n27 VSUBS 0.005982f
C74 B.n28 VSUBS 0.005982f
C75 B.n29 VSUBS 0.005982f
C76 B.n30 VSUBS 0.005982f
C77 B.n31 VSUBS 0.005982f
C78 B.n32 VSUBS 0.005982f
C79 B.n33 VSUBS 0.005982f
C80 B.n34 VSUBS 0.005982f
C81 B.n35 VSUBS 0.005982f
C82 B.n36 VSUBS 0.005982f
C83 B.n37 VSUBS 0.005982f
C84 B.t10 VSUBS 0.42609f
C85 B.t11 VSUBS 0.441653f
C86 B.t9 VSUBS 1.17618f
C87 B.n38 VSUBS 0.218285f
C88 B.n39 VSUBS 0.059702f
C89 B.n40 VSUBS 0.01386f
C90 B.n41 VSUBS 0.005982f
C91 B.n42 VSUBS 0.005982f
C92 B.n43 VSUBS 0.005982f
C93 B.n44 VSUBS 0.005982f
C94 B.n45 VSUBS 0.005982f
C95 B.t1 VSUBS 0.426077f
C96 B.t2 VSUBS 0.441642f
C97 B.t0 VSUBS 1.17618f
C98 B.n46 VSUBS 0.218295f
C99 B.n47 VSUBS 0.059715f
C100 B.n48 VSUBS 0.005982f
C101 B.n49 VSUBS 0.005982f
C102 B.n50 VSUBS 0.005982f
C103 B.n51 VSUBS 0.005982f
C104 B.n52 VSUBS 0.005982f
C105 B.n53 VSUBS 0.005982f
C106 B.n54 VSUBS 0.005982f
C107 B.n55 VSUBS 0.005982f
C108 B.n56 VSUBS 0.005982f
C109 B.n57 VSUBS 0.005982f
C110 B.n58 VSUBS 0.005982f
C111 B.n59 VSUBS 0.005982f
C112 B.n60 VSUBS 0.005982f
C113 B.n61 VSUBS 0.005982f
C114 B.n62 VSUBS 0.005982f
C115 B.n63 VSUBS 0.005982f
C116 B.n64 VSUBS 0.005982f
C117 B.n65 VSUBS 0.005982f
C118 B.n66 VSUBS 0.005982f
C119 B.n67 VSUBS 0.005982f
C120 B.n68 VSUBS 0.005982f
C121 B.n69 VSUBS 0.005982f
C122 B.n70 VSUBS 0.005982f
C123 B.n71 VSUBS 0.005982f
C124 B.n72 VSUBS 0.013926f
C125 B.n73 VSUBS 0.005982f
C126 B.n74 VSUBS 0.005982f
C127 B.n75 VSUBS 0.005982f
C128 B.n76 VSUBS 0.005982f
C129 B.n77 VSUBS 0.005982f
C130 B.n78 VSUBS 0.005982f
C131 B.n79 VSUBS 0.005982f
C132 B.n80 VSUBS 0.005982f
C133 B.n81 VSUBS 0.005982f
C134 B.n82 VSUBS 0.005982f
C135 B.n83 VSUBS 0.005982f
C136 B.n84 VSUBS 0.005982f
C137 B.n85 VSUBS 0.005982f
C138 B.n86 VSUBS 0.005982f
C139 B.n87 VSUBS 0.005982f
C140 B.n88 VSUBS 0.005982f
C141 B.n89 VSUBS 0.005982f
C142 B.n90 VSUBS 0.005982f
C143 B.n91 VSUBS 0.005982f
C144 B.n92 VSUBS 0.005982f
C145 B.n93 VSUBS 0.005982f
C146 B.n94 VSUBS 0.005982f
C147 B.n95 VSUBS 0.013697f
C148 B.n96 VSUBS 0.005982f
C149 B.n97 VSUBS 0.005982f
C150 B.n98 VSUBS 0.005982f
C151 B.n99 VSUBS 0.005982f
C152 B.n100 VSUBS 0.005982f
C153 B.n101 VSUBS 0.005982f
C154 B.n102 VSUBS 0.005982f
C155 B.n103 VSUBS 0.005982f
C156 B.n104 VSUBS 0.005982f
C157 B.n105 VSUBS 0.005982f
C158 B.n106 VSUBS 0.005982f
C159 B.n107 VSUBS 0.005982f
C160 B.n108 VSUBS 0.005982f
C161 B.n109 VSUBS 0.005982f
C162 B.n110 VSUBS 0.005982f
C163 B.n111 VSUBS 0.005982f
C164 B.n112 VSUBS 0.005982f
C165 B.n113 VSUBS 0.005982f
C166 B.n114 VSUBS 0.005982f
C167 B.n115 VSUBS 0.005982f
C168 B.n116 VSUBS 0.005982f
C169 B.n117 VSUBS 0.005982f
C170 B.n118 VSUBS 0.005982f
C171 B.n119 VSUBS 0.005982f
C172 B.n120 VSUBS 0.00563f
C173 B.n121 VSUBS 0.005982f
C174 B.n122 VSUBS 0.005982f
C175 B.n123 VSUBS 0.005982f
C176 B.n124 VSUBS 0.005982f
C177 B.n125 VSUBS 0.005982f
C178 B.t5 VSUBS 0.42609f
C179 B.t4 VSUBS 0.441653f
C180 B.t3 VSUBS 1.17618f
C181 B.n126 VSUBS 0.218285f
C182 B.n127 VSUBS 0.059702f
C183 B.n128 VSUBS 0.005982f
C184 B.n129 VSUBS 0.005982f
C185 B.n130 VSUBS 0.005982f
C186 B.n131 VSUBS 0.005982f
C187 B.n132 VSUBS 0.005982f
C188 B.n133 VSUBS 0.005982f
C189 B.n134 VSUBS 0.005982f
C190 B.n135 VSUBS 0.005982f
C191 B.n136 VSUBS 0.005982f
C192 B.n137 VSUBS 0.005982f
C193 B.n138 VSUBS 0.005982f
C194 B.n139 VSUBS 0.005982f
C195 B.n140 VSUBS 0.005982f
C196 B.n141 VSUBS 0.005982f
C197 B.n142 VSUBS 0.005982f
C198 B.n143 VSUBS 0.005982f
C199 B.n144 VSUBS 0.005982f
C200 B.n145 VSUBS 0.005982f
C201 B.n146 VSUBS 0.005982f
C202 B.n147 VSUBS 0.005982f
C203 B.n148 VSUBS 0.005982f
C204 B.n149 VSUBS 0.005982f
C205 B.n150 VSUBS 0.005982f
C206 B.n151 VSUBS 0.005982f
C207 B.n152 VSUBS 0.013926f
C208 B.n153 VSUBS 0.005982f
C209 B.n154 VSUBS 0.005982f
C210 B.n155 VSUBS 0.005982f
C211 B.n156 VSUBS 0.005982f
C212 B.n157 VSUBS 0.005982f
C213 B.n158 VSUBS 0.005982f
C214 B.n159 VSUBS 0.005982f
C215 B.n160 VSUBS 0.005982f
C216 B.n161 VSUBS 0.005982f
C217 B.n162 VSUBS 0.005982f
C218 B.n163 VSUBS 0.005982f
C219 B.n164 VSUBS 0.005982f
C220 B.n165 VSUBS 0.005982f
C221 B.n166 VSUBS 0.005982f
C222 B.n167 VSUBS 0.005982f
C223 B.n168 VSUBS 0.005982f
C224 B.n169 VSUBS 0.005982f
C225 B.n170 VSUBS 0.005982f
C226 B.n171 VSUBS 0.005982f
C227 B.n172 VSUBS 0.005982f
C228 B.n173 VSUBS 0.005982f
C229 B.n174 VSUBS 0.005982f
C230 B.n175 VSUBS 0.005982f
C231 B.n176 VSUBS 0.005982f
C232 B.n177 VSUBS 0.005982f
C233 B.n178 VSUBS 0.005982f
C234 B.n179 VSUBS 0.005982f
C235 B.n180 VSUBS 0.005982f
C236 B.n181 VSUBS 0.005982f
C237 B.n182 VSUBS 0.005982f
C238 B.n183 VSUBS 0.005982f
C239 B.n184 VSUBS 0.005982f
C240 B.n185 VSUBS 0.005982f
C241 B.n186 VSUBS 0.005982f
C242 B.n187 VSUBS 0.005982f
C243 B.n188 VSUBS 0.005982f
C244 B.n189 VSUBS 0.005982f
C245 B.n190 VSUBS 0.005982f
C246 B.n191 VSUBS 0.005982f
C247 B.n192 VSUBS 0.005982f
C248 B.n193 VSUBS 0.013697f
C249 B.n194 VSUBS 0.013697f
C250 B.n195 VSUBS 0.013926f
C251 B.n196 VSUBS 0.005982f
C252 B.n197 VSUBS 0.005982f
C253 B.n198 VSUBS 0.005982f
C254 B.n199 VSUBS 0.005982f
C255 B.n200 VSUBS 0.005982f
C256 B.n201 VSUBS 0.005982f
C257 B.n202 VSUBS 0.005982f
C258 B.n203 VSUBS 0.005982f
C259 B.n204 VSUBS 0.005982f
C260 B.n205 VSUBS 0.005982f
C261 B.n206 VSUBS 0.005982f
C262 B.n207 VSUBS 0.005982f
C263 B.n208 VSUBS 0.005982f
C264 B.n209 VSUBS 0.005982f
C265 B.n210 VSUBS 0.005982f
C266 B.n211 VSUBS 0.005982f
C267 B.n212 VSUBS 0.005982f
C268 B.n213 VSUBS 0.005982f
C269 B.n214 VSUBS 0.005982f
C270 B.n215 VSUBS 0.005982f
C271 B.n216 VSUBS 0.005982f
C272 B.n217 VSUBS 0.005982f
C273 B.n218 VSUBS 0.005982f
C274 B.n219 VSUBS 0.005982f
C275 B.n220 VSUBS 0.005982f
C276 B.n221 VSUBS 0.005982f
C277 B.n222 VSUBS 0.005982f
C278 B.n223 VSUBS 0.005982f
C279 B.n224 VSUBS 0.005982f
C280 B.n225 VSUBS 0.005982f
C281 B.n226 VSUBS 0.005982f
C282 B.n227 VSUBS 0.005982f
C283 B.n228 VSUBS 0.005982f
C284 B.n229 VSUBS 0.005982f
C285 B.n230 VSUBS 0.005982f
C286 B.n231 VSUBS 0.005982f
C287 B.n232 VSUBS 0.005982f
C288 B.n233 VSUBS 0.005982f
C289 B.n234 VSUBS 0.005982f
C290 B.n235 VSUBS 0.005982f
C291 B.n236 VSUBS 0.005982f
C292 B.n237 VSUBS 0.005982f
C293 B.n238 VSUBS 0.005982f
C294 B.n239 VSUBS 0.005982f
C295 B.n240 VSUBS 0.005982f
C296 B.n241 VSUBS 0.005982f
C297 B.n242 VSUBS 0.005982f
C298 B.n243 VSUBS 0.005982f
C299 B.n244 VSUBS 0.005982f
C300 B.n245 VSUBS 0.005982f
C301 B.n246 VSUBS 0.005982f
C302 B.n247 VSUBS 0.005982f
C303 B.n248 VSUBS 0.005982f
C304 B.n249 VSUBS 0.005982f
C305 B.n250 VSUBS 0.005982f
C306 B.n251 VSUBS 0.005982f
C307 B.n252 VSUBS 0.005982f
C308 B.n253 VSUBS 0.005982f
C309 B.n254 VSUBS 0.005982f
C310 B.n255 VSUBS 0.005982f
C311 B.n256 VSUBS 0.005982f
C312 B.n257 VSUBS 0.005982f
C313 B.n258 VSUBS 0.005982f
C314 B.n259 VSUBS 0.005982f
C315 B.n260 VSUBS 0.005982f
C316 B.n261 VSUBS 0.005982f
C317 B.n262 VSUBS 0.005982f
C318 B.n263 VSUBS 0.005982f
C319 B.n264 VSUBS 0.005982f
C320 B.n265 VSUBS 0.005982f
C321 B.n266 VSUBS 0.005982f
C322 B.n267 VSUBS 0.005982f
C323 B.n268 VSUBS 0.005982f
C324 B.n269 VSUBS 0.00563f
C325 B.n270 VSUBS 0.01386f
C326 B.n271 VSUBS 0.003343f
C327 B.n272 VSUBS 0.005982f
C328 B.n273 VSUBS 0.005982f
C329 B.n274 VSUBS 0.005982f
C330 B.n275 VSUBS 0.005982f
C331 B.n276 VSUBS 0.005982f
C332 B.n277 VSUBS 0.005982f
C333 B.n278 VSUBS 0.005982f
C334 B.n279 VSUBS 0.005982f
C335 B.n280 VSUBS 0.005982f
C336 B.n281 VSUBS 0.005982f
C337 B.n282 VSUBS 0.005982f
C338 B.n283 VSUBS 0.005982f
C339 B.t8 VSUBS 0.426077f
C340 B.t7 VSUBS 0.441642f
C341 B.t6 VSUBS 1.17618f
C342 B.n284 VSUBS 0.218295f
C343 B.n285 VSUBS 0.059715f
C344 B.n286 VSUBS 0.01386f
C345 B.n287 VSUBS 0.003343f
C346 B.n288 VSUBS 0.005982f
C347 B.n289 VSUBS 0.005982f
C348 B.n290 VSUBS 0.005982f
C349 B.n291 VSUBS 0.005982f
C350 B.n292 VSUBS 0.005982f
C351 B.n293 VSUBS 0.005982f
C352 B.n294 VSUBS 0.005982f
C353 B.n295 VSUBS 0.005982f
C354 B.n296 VSUBS 0.005982f
C355 B.n297 VSUBS 0.005982f
C356 B.n298 VSUBS 0.005982f
C357 B.n299 VSUBS 0.005982f
C358 B.n300 VSUBS 0.005982f
C359 B.n301 VSUBS 0.005982f
C360 B.n302 VSUBS 0.005982f
C361 B.n303 VSUBS 0.005982f
C362 B.n304 VSUBS 0.005982f
C363 B.n305 VSUBS 0.005982f
C364 B.n306 VSUBS 0.005982f
C365 B.n307 VSUBS 0.005982f
C366 B.n308 VSUBS 0.005982f
C367 B.n309 VSUBS 0.005982f
C368 B.n310 VSUBS 0.005982f
C369 B.n311 VSUBS 0.005982f
C370 B.n312 VSUBS 0.005982f
C371 B.n313 VSUBS 0.005982f
C372 B.n314 VSUBS 0.005982f
C373 B.n315 VSUBS 0.005982f
C374 B.n316 VSUBS 0.005982f
C375 B.n317 VSUBS 0.005982f
C376 B.n318 VSUBS 0.005982f
C377 B.n319 VSUBS 0.005982f
C378 B.n320 VSUBS 0.005982f
C379 B.n321 VSUBS 0.005982f
C380 B.n322 VSUBS 0.005982f
C381 B.n323 VSUBS 0.005982f
C382 B.n324 VSUBS 0.005982f
C383 B.n325 VSUBS 0.005982f
C384 B.n326 VSUBS 0.005982f
C385 B.n327 VSUBS 0.005982f
C386 B.n328 VSUBS 0.005982f
C387 B.n329 VSUBS 0.005982f
C388 B.n330 VSUBS 0.005982f
C389 B.n331 VSUBS 0.005982f
C390 B.n332 VSUBS 0.005982f
C391 B.n333 VSUBS 0.005982f
C392 B.n334 VSUBS 0.005982f
C393 B.n335 VSUBS 0.005982f
C394 B.n336 VSUBS 0.005982f
C395 B.n337 VSUBS 0.005982f
C396 B.n338 VSUBS 0.005982f
C397 B.n339 VSUBS 0.005982f
C398 B.n340 VSUBS 0.005982f
C399 B.n341 VSUBS 0.005982f
C400 B.n342 VSUBS 0.005982f
C401 B.n343 VSUBS 0.005982f
C402 B.n344 VSUBS 0.005982f
C403 B.n345 VSUBS 0.005982f
C404 B.n346 VSUBS 0.005982f
C405 B.n347 VSUBS 0.005982f
C406 B.n348 VSUBS 0.005982f
C407 B.n349 VSUBS 0.005982f
C408 B.n350 VSUBS 0.005982f
C409 B.n351 VSUBS 0.005982f
C410 B.n352 VSUBS 0.005982f
C411 B.n353 VSUBS 0.005982f
C412 B.n354 VSUBS 0.005982f
C413 B.n355 VSUBS 0.005982f
C414 B.n356 VSUBS 0.005982f
C415 B.n357 VSUBS 0.005982f
C416 B.n358 VSUBS 0.005982f
C417 B.n359 VSUBS 0.005982f
C418 B.n360 VSUBS 0.005982f
C419 B.n361 VSUBS 0.005982f
C420 B.n362 VSUBS 0.013926f
C421 B.n363 VSUBS 0.013205f
C422 B.n364 VSUBS 0.014419f
C423 B.n365 VSUBS 0.005982f
C424 B.n366 VSUBS 0.005982f
C425 B.n367 VSUBS 0.005982f
C426 B.n368 VSUBS 0.005982f
C427 B.n369 VSUBS 0.005982f
C428 B.n370 VSUBS 0.005982f
C429 B.n371 VSUBS 0.005982f
C430 B.n372 VSUBS 0.005982f
C431 B.n373 VSUBS 0.005982f
C432 B.n374 VSUBS 0.005982f
C433 B.n375 VSUBS 0.005982f
C434 B.n376 VSUBS 0.005982f
C435 B.n377 VSUBS 0.005982f
C436 B.n378 VSUBS 0.005982f
C437 B.n379 VSUBS 0.005982f
C438 B.n380 VSUBS 0.005982f
C439 B.n381 VSUBS 0.005982f
C440 B.n382 VSUBS 0.005982f
C441 B.n383 VSUBS 0.005982f
C442 B.n384 VSUBS 0.005982f
C443 B.n385 VSUBS 0.005982f
C444 B.n386 VSUBS 0.005982f
C445 B.n387 VSUBS 0.005982f
C446 B.n388 VSUBS 0.005982f
C447 B.n389 VSUBS 0.005982f
C448 B.n390 VSUBS 0.005982f
C449 B.n391 VSUBS 0.005982f
C450 B.n392 VSUBS 0.005982f
C451 B.n393 VSUBS 0.005982f
C452 B.n394 VSUBS 0.005982f
C453 B.n395 VSUBS 0.005982f
C454 B.n396 VSUBS 0.005982f
C455 B.n397 VSUBS 0.005982f
C456 B.n398 VSUBS 0.005982f
C457 B.n399 VSUBS 0.005982f
C458 B.n400 VSUBS 0.005982f
C459 B.n401 VSUBS 0.005982f
C460 B.n402 VSUBS 0.005982f
C461 B.n403 VSUBS 0.005982f
C462 B.n404 VSUBS 0.005982f
C463 B.n405 VSUBS 0.005982f
C464 B.n406 VSUBS 0.005982f
C465 B.n407 VSUBS 0.005982f
C466 B.n408 VSUBS 0.005982f
C467 B.n409 VSUBS 0.005982f
C468 B.n410 VSUBS 0.005982f
C469 B.n411 VSUBS 0.005982f
C470 B.n412 VSUBS 0.005982f
C471 B.n413 VSUBS 0.005982f
C472 B.n414 VSUBS 0.005982f
C473 B.n415 VSUBS 0.005982f
C474 B.n416 VSUBS 0.005982f
C475 B.n417 VSUBS 0.005982f
C476 B.n418 VSUBS 0.005982f
C477 B.n419 VSUBS 0.005982f
C478 B.n420 VSUBS 0.005982f
C479 B.n421 VSUBS 0.005982f
C480 B.n422 VSUBS 0.005982f
C481 B.n423 VSUBS 0.005982f
C482 B.n424 VSUBS 0.005982f
C483 B.n425 VSUBS 0.005982f
C484 B.n426 VSUBS 0.005982f
C485 B.n427 VSUBS 0.005982f
C486 B.n428 VSUBS 0.005982f
C487 B.n429 VSUBS 0.005982f
C488 B.n430 VSUBS 0.005982f
C489 B.n431 VSUBS 0.013697f
C490 B.n432 VSUBS 0.013697f
C491 B.n433 VSUBS 0.013926f
C492 B.n434 VSUBS 0.005982f
C493 B.n435 VSUBS 0.005982f
C494 B.n436 VSUBS 0.005982f
C495 B.n437 VSUBS 0.005982f
C496 B.n438 VSUBS 0.005982f
C497 B.n439 VSUBS 0.005982f
C498 B.n440 VSUBS 0.005982f
C499 B.n441 VSUBS 0.005982f
C500 B.n442 VSUBS 0.005982f
C501 B.n443 VSUBS 0.005982f
C502 B.n444 VSUBS 0.005982f
C503 B.n445 VSUBS 0.005982f
C504 B.n446 VSUBS 0.005982f
C505 B.n447 VSUBS 0.005982f
C506 B.n448 VSUBS 0.005982f
C507 B.n449 VSUBS 0.005982f
C508 B.n450 VSUBS 0.005982f
C509 B.n451 VSUBS 0.005982f
C510 B.n452 VSUBS 0.005982f
C511 B.n453 VSUBS 0.005982f
C512 B.n454 VSUBS 0.005982f
C513 B.n455 VSUBS 0.005982f
C514 B.n456 VSUBS 0.005982f
C515 B.n457 VSUBS 0.005982f
C516 B.n458 VSUBS 0.005982f
C517 B.n459 VSUBS 0.005982f
C518 B.n460 VSUBS 0.005982f
C519 B.n461 VSUBS 0.005982f
C520 B.n462 VSUBS 0.005982f
C521 B.n463 VSUBS 0.005982f
C522 B.n464 VSUBS 0.005982f
C523 B.n465 VSUBS 0.005982f
C524 B.n466 VSUBS 0.005982f
C525 B.n467 VSUBS 0.005982f
C526 B.n468 VSUBS 0.005982f
C527 B.n469 VSUBS 0.005982f
C528 B.n470 VSUBS 0.005982f
C529 B.n471 VSUBS 0.005982f
C530 B.n472 VSUBS 0.005982f
C531 B.n473 VSUBS 0.005982f
C532 B.n474 VSUBS 0.005982f
C533 B.n475 VSUBS 0.005982f
C534 B.n476 VSUBS 0.005982f
C535 B.n477 VSUBS 0.005982f
C536 B.n478 VSUBS 0.005982f
C537 B.n479 VSUBS 0.005982f
C538 B.n480 VSUBS 0.005982f
C539 B.n481 VSUBS 0.005982f
C540 B.n482 VSUBS 0.005982f
C541 B.n483 VSUBS 0.005982f
C542 B.n484 VSUBS 0.005982f
C543 B.n485 VSUBS 0.005982f
C544 B.n486 VSUBS 0.005982f
C545 B.n487 VSUBS 0.005982f
C546 B.n488 VSUBS 0.005982f
C547 B.n489 VSUBS 0.005982f
C548 B.n490 VSUBS 0.005982f
C549 B.n491 VSUBS 0.005982f
C550 B.n492 VSUBS 0.005982f
C551 B.n493 VSUBS 0.005982f
C552 B.n494 VSUBS 0.005982f
C553 B.n495 VSUBS 0.005982f
C554 B.n496 VSUBS 0.005982f
C555 B.n497 VSUBS 0.005982f
C556 B.n498 VSUBS 0.005982f
C557 B.n499 VSUBS 0.005982f
C558 B.n500 VSUBS 0.005982f
C559 B.n501 VSUBS 0.005982f
C560 B.n502 VSUBS 0.005982f
C561 B.n503 VSUBS 0.005982f
C562 B.n504 VSUBS 0.005982f
C563 B.n505 VSUBS 0.005982f
C564 B.n506 VSUBS 0.005982f
C565 B.n507 VSUBS 0.00563f
C566 B.n508 VSUBS 0.01386f
C567 B.n509 VSUBS 0.003343f
C568 B.n510 VSUBS 0.005982f
C569 B.n511 VSUBS 0.005982f
C570 B.n512 VSUBS 0.005982f
C571 B.n513 VSUBS 0.005982f
C572 B.n514 VSUBS 0.005982f
C573 B.n515 VSUBS 0.005982f
C574 B.n516 VSUBS 0.005982f
C575 B.n517 VSUBS 0.005982f
C576 B.n518 VSUBS 0.005982f
C577 B.n519 VSUBS 0.005982f
C578 B.n520 VSUBS 0.005982f
C579 B.n521 VSUBS 0.005982f
C580 B.n522 VSUBS 0.003343f
C581 B.n523 VSUBS 0.005982f
C582 B.n524 VSUBS 0.005982f
C583 B.n525 VSUBS 0.00563f
C584 B.n526 VSUBS 0.005982f
C585 B.n527 VSUBS 0.005982f
C586 B.n528 VSUBS 0.005982f
C587 B.n529 VSUBS 0.005982f
C588 B.n530 VSUBS 0.005982f
C589 B.n531 VSUBS 0.005982f
C590 B.n532 VSUBS 0.005982f
C591 B.n533 VSUBS 0.005982f
C592 B.n534 VSUBS 0.005982f
C593 B.n535 VSUBS 0.005982f
C594 B.n536 VSUBS 0.005982f
C595 B.n537 VSUBS 0.005982f
C596 B.n538 VSUBS 0.005982f
C597 B.n539 VSUBS 0.005982f
C598 B.n540 VSUBS 0.005982f
C599 B.n541 VSUBS 0.005982f
C600 B.n542 VSUBS 0.005982f
C601 B.n543 VSUBS 0.005982f
C602 B.n544 VSUBS 0.005982f
C603 B.n545 VSUBS 0.005982f
C604 B.n546 VSUBS 0.005982f
C605 B.n547 VSUBS 0.005982f
C606 B.n548 VSUBS 0.005982f
C607 B.n549 VSUBS 0.005982f
C608 B.n550 VSUBS 0.005982f
C609 B.n551 VSUBS 0.005982f
C610 B.n552 VSUBS 0.005982f
C611 B.n553 VSUBS 0.005982f
C612 B.n554 VSUBS 0.005982f
C613 B.n555 VSUBS 0.005982f
C614 B.n556 VSUBS 0.005982f
C615 B.n557 VSUBS 0.005982f
C616 B.n558 VSUBS 0.005982f
C617 B.n559 VSUBS 0.005982f
C618 B.n560 VSUBS 0.005982f
C619 B.n561 VSUBS 0.005982f
C620 B.n562 VSUBS 0.005982f
C621 B.n563 VSUBS 0.005982f
C622 B.n564 VSUBS 0.005982f
C623 B.n565 VSUBS 0.005982f
C624 B.n566 VSUBS 0.005982f
C625 B.n567 VSUBS 0.005982f
C626 B.n568 VSUBS 0.005982f
C627 B.n569 VSUBS 0.005982f
C628 B.n570 VSUBS 0.005982f
C629 B.n571 VSUBS 0.005982f
C630 B.n572 VSUBS 0.005982f
C631 B.n573 VSUBS 0.005982f
C632 B.n574 VSUBS 0.005982f
C633 B.n575 VSUBS 0.005982f
C634 B.n576 VSUBS 0.005982f
C635 B.n577 VSUBS 0.005982f
C636 B.n578 VSUBS 0.005982f
C637 B.n579 VSUBS 0.005982f
C638 B.n580 VSUBS 0.005982f
C639 B.n581 VSUBS 0.005982f
C640 B.n582 VSUBS 0.005982f
C641 B.n583 VSUBS 0.005982f
C642 B.n584 VSUBS 0.005982f
C643 B.n585 VSUBS 0.005982f
C644 B.n586 VSUBS 0.005982f
C645 B.n587 VSUBS 0.005982f
C646 B.n588 VSUBS 0.005982f
C647 B.n589 VSUBS 0.005982f
C648 B.n590 VSUBS 0.005982f
C649 B.n591 VSUBS 0.005982f
C650 B.n592 VSUBS 0.005982f
C651 B.n593 VSUBS 0.005982f
C652 B.n594 VSUBS 0.005982f
C653 B.n595 VSUBS 0.005982f
C654 B.n596 VSUBS 0.005982f
C655 B.n597 VSUBS 0.005982f
C656 B.n598 VSUBS 0.013926f
C657 B.n599 VSUBS 0.013697f
C658 B.n600 VSUBS 0.013697f
C659 B.n601 VSUBS 0.005982f
C660 B.n602 VSUBS 0.005982f
C661 B.n603 VSUBS 0.005982f
C662 B.n604 VSUBS 0.005982f
C663 B.n605 VSUBS 0.005982f
C664 B.n606 VSUBS 0.005982f
C665 B.n607 VSUBS 0.005982f
C666 B.n608 VSUBS 0.005982f
C667 B.n609 VSUBS 0.005982f
C668 B.n610 VSUBS 0.005982f
C669 B.n611 VSUBS 0.005982f
C670 B.n612 VSUBS 0.005982f
C671 B.n613 VSUBS 0.005982f
C672 B.n614 VSUBS 0.005982f
C673 B.n615 VSUBS 0.005982f
C674 B.n616 VSUBS 0.005982f
C675 B.n617 VSUBS 0.005982f
C676 B.n618 VSUBS 0.005982f
C677 B.n619 VSUBS 0.005982f
C678 B.n620 VSUBS 0.005982f
C679 B.n621 VSUBS 0.005982f
C680 B.n622 VSUBS 0.005982f
C681 B.n623 VSUBS 0.005982f
C682 B.n624 VSUBS 0.005982f
C683 B.n625 VSUBS 0.005982f
C684 B.n626 VSUBS 0.005982f
C685 B.n627 VSUBS 0.005982f
C686 B.n628 VSUBS 0.005982f
C687 B.n629 VSUBS 0.005982f
C688 B.n630 VSUBS 0.005982f
C689 B.n631 VSUBS 0.007806f
C690 B.n632 VSUBS 0.008316f
C691 B.n633 VSUBS 0.016537f
.ends

