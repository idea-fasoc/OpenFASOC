* NGSPICE file created from diff_pair_sample_1763.ext - technology: sky130A

.subckt diff_pair_sample_1763 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0 ps=0 w=1.02 l=0.66
X1 VDD2.t5 VN.t0 VTAIL.t8 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.3978 ps=2.82 w=1.02 l=0.66
X2 B.t8 B.t6 B.t7 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0 ps=0 w=1.02 l=0.66
X3 B.t5 B.t3 B.t4 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0 ps=0 w=1.02 l=0.66
X4 VDD2.t4 VN.t1 VTAIL.t3 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0.1683 ps=1.35 w=1.02 l=0.66
X5 VTAIL.t6 VN.t2 VDD2.t3 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.1683 ps=1.35 w=1.02 l=0.66
X6 VDD2.t2 VN.t3 VTAIL.t5 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.3978 ps=2.82 w=1.02 l=0.66
X7 VTAIL.t4 VN.t4 VDD2.t1 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.1683 ps=1.35 w=1.02 l=0.66
X8 VDD1.t5 VP.t0 VTAIL.t9 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0.1683 ps=1.35 w=1.02 l=0.66
X9 VDD2.t0 VN.t5 VTAIL.t7 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0.1683 ps=1.35 w=1.02 l=0.66
X10 B.t2 B.t0 B.t1 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0 ps=0 w=1.02 l=0.66
X11 VDD1.t4 VP.t1 VTAIL.t10 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.3978 pd=2.82 as=0.1683 ps=1.35 w=1.02 l=0.66
X12 VTAIL.t11 VP.t2 VDD1.t3 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.1683 ps=1.35 w=1.02 l=0.66
X13 VDD1.t2 VP.t3 VTAIL.t1 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.3978 ps=2.82 w=1.02 l=0.66
X14 VDD1.t1 VP.t4 VTAIL.t0 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.3978 ps=2.82 w=1.02 l=0.66
X15 VTAIL.t2 VP.t5 VDD1.t0 w_n1762_n1172# sky130_fd_pr__pfet_01v8 ad=0.1683 pd=1.35 as=0.1683 ps=1.35 w=1.02 l=0.66
R0 B.n147 B.n50 585
R1 B.n146 B.n145 585
R2 B.n144 B.n51 585
R3 B.n143 B.n142 585
R4 B.n141 B.n52 585
R5 B.n140 B.n139 585
R6 B.n138 B.n53 585
R7 B.n137 B.n136 585
R8 B.n135 B.n54 585
R9 B.n134 B.n133 585
R10 B.n129 B.n55 585
R11 B.n128 B.n127 585
R12 B.n126 B.n56 585
R13 B.n125 B.n124 585
R14 B.n123 B.n57 585
R15 B.n122 B.n121 585
R16 B.n120 B.n58 585
R17 B.n119 B.n118 585
R18 B.n117 B.n59 585
R19 B.n115 B.n114 585
R20 B.n113 B.n62 585
R21 B.n112 B.n111 585
R22 B.n110 B.n63 585
R23 B.n109 B.n108 585
R24 B.n107 B.n64 585
R25 B.n106 B.n105 585
R26 B.n104 B.n65 585
R27 B.n103 B.n102 585
R28 B.n149 B.n148 585
R29 B.n150 B.n49 585
R30 B.n152 B.n151 585
R31 B.n153 B.n48 585
R32 B.n155 B.n154 585
R33 B.n156 B.n47 585
R34 B.n158 B.n157 585
R35 B.n159 B.n46 585
R36 B.n161 B.n160 585
R37 B.n162 B.n45 585
R38 B.n164 B.n163 585
R39 B.n165 B.n44 585
R40 B.n167 B.n166 585
R41 B.n168 B.n43 585
R42 B.n170 B.n169 585
R43 B.n171 B.n42 585
R44 B.n173 B.n172 585
R45 B.n174 B.n41 585
R46 B.n176 B.n175 585
R47 B.n177 B.n40 585
R48 B.n179 B.n178 585
R49 B.n180 B.n39 585
R50 B.n182 B.n181 585
R51 B.n183 B.n38 585
R52 B.n185 B.n184 585
R53 B.n186 B.n37 585
R54 B.n188 B.n187 585
R55 B.n189 B.n36 585
R56 B.n191 B.n190 585
R57 B.n192 B.n35 585
R58 B.n194 B.n193 585
R59 B.n195 B.n34 585
R60 B.n197 B.n196 585
R61 B.n198 B.n33 585
R62 B.n200 B.n199 585
R63 B.n201 B.n32 585
R64 B.n203 B.n202 585
R65 B.n204 B.n31 585
R66 B.n206 B.n205 585
R67 B.n207 B.n30 585
R68 B.n251 B.n250 585
R69 B.n249 B.n12 585
R70 B.n248 B.n247 585
R71 B.n246 B.n13 585
R72 B.n245 B.n244 585
R73 B.n243 B.n14 585
R74 B.n242 B.n241 585
R75 B.n240 B.n15 585
R76 B.n239 B.n238 585
R77 B.n237 B.n236 585
R78 B.n235 B.n19 585
R79 B.n234 B.n233 585
R80 B.n232 B.n20 585
R81 B.n231 B.n230 585
R82 B.n229 B.n21 585
R83 B.n228 B.n227 585
R84 B.n226 B.n22 585
R85 B.n225 B.n224 585
R86 B.n223 B.n23 585
R87 B.n221 B.n220 585
R88 B.n219 B.n26 585
R89 B.n218 B.n217 585
R90 B.n216 B.n27 585
R91 B.n215 B.n214 585
R92 B.n213 B.n28 585
R93 B.n212 B.n211 585
R94 B.n210 B.n29 585
R95 B.n209 B.n208 585
R96 B.n252 B.n11 585
R97 B.n254 B.n253 585
R98 B.n255 B.n10 585
R99 B.n257 B.n256 585
R100 B.n258 B.n9 585
R101 B.n260 B.n259 585
R102 B.n261 B.n8 585
R103 B.n263 B.n262 585
R104 B.n264 B.n7 585
R105 B.n266 B.n265 585
R106 B.n267 B.n6 585
R107 B.n269 B.n268 585
R108 B.n270 B.n5 585
R109 B.n272 B.n271 585
R110 B.n273 B.n4 585
R111 B.n275 B.n274 585
R112 B.n276 B.n3 585
R113 B.n278 B.n277 585
R114 B.n279 B.n0 585
R115 B.n2 B.n1 585
R116 B.n76 B.n75 585
R117 B.n77 B.n74 585
R118 B.n79 B.n78 585
R119 B.n80 B.n73 585
R120 B.n82 B.n81 585
R121 B.n83 B.n72 585
R122 B.n85 B.n84 585
R123 B.n86 B.n71 585
R124 B.n88 B.n87 585
R125 B.n89 B.n70 585
R126 B.n91 B.n90 585
R127 B.n92 B.n69 585
R128 B.n94 B.n93 585
R129 B.n95 B.n68 585
R130 B.n97 B.n96 585
R131 B.n98 B.n67 585
R132 B.n100 B.n99 585
R133 B.n101 B.n66 585
R134 B.n102 B.n101 559.769
R135 B.n148 B.n147 559.769
R136 B.n208 B.n207 559.769
R137 B.n250 B.n11 559.769
R138 B.n60 B.t4 380.788
R139 B.n130 B.t1 380.788
R140 B.n24 B.t11 380.788
R141 B.n16 B.t8 380.788
R142 B.n61 B.t5 361.587
R143 B.n131 B.t2 361.587
R144 B.n25 B.t10 361.587
R145 B.n17 B.t7 361.587
R146 B.n281 B.n280 256.663
R147 B.n60 B.t3 240.732
R148 B.n130 B.t0 240.732
R149 B.n24 B.t9 240.732
R150 B.n16 B.t6 240.732
R151 B.n280 B.n279 235.042
R152 B.n280 B.n2 235.042
R153 B.n102 B.n65 163.367
R154 B.n106 B.n65 163.367
R155 B.n107 B.n106 163.367
R156 B.n108 B.n107 163.367
R157 B.n108 B.n63 163.367
R158 B.n112 B.n63 163.367
R159 B.n113 B.n112 163.367
R160 B.n114 B.n113 163.367
R161 B.n114 B.n59 163.367
R162 B.n119 B.n59 163.367
R163 B.n120 B.n119 163.367
R164 B.n121 B.n120 163.367
R165 B.n121 B.n57 163.367
R166 B.n125 B.n57 163.367
R167 B.n126 B.n125 163.367
R168 B.n127 B.n126 163.367
R169 B.n127 B.n55 163.367
R170 B.n134 B.n55 163.367
R171 B.n135 B.n134 163.367
R172 B.n136 B.n135 163.367
R173 B.n136 B.n53 163.367
R174 B.n140 B.n53 163.367
R175 B.n141 B.n140 163.367
R176 B.n142 B.n141 163.367
R177 B.n142 B.n51 163.367
R178 B.n146 B.n51 163.367
R179 B.n147 B.n146 163.367
R180 B.n207 B.n206 163.367
R181 B.n206 B.n31 163.367
R182 B.n202 B.n31 163.367
R183 B.n202 B.n201 163.367
R184 B.n201 B.n200 163.367
R185 B.n200 B.n33 163.367
R186 B.n196 B.n33 163.367
R187 B.n196 B.n195 163.367
R188 B.n195 B.n194 163.367
R189 B.n194 B.n35 163.367
R190 B.n190 B.n35 163.367
R191 B.n190 B.n189 163.367
R192 B.n189 B.n188 163.367
R193 B.n188 B.n37 163.367
R194 B.n184 B.n37 163.367
R195 B.n184 B.n183 163.367
R196 B.n183 B.n182 163.367
R197 B.n182 B.n39 163.367
R198 B.n178 B.n39 163.367
R199 B.n178 B.n177 163.367
R200 B.n177 B.n176 163.367
R201 B.n176 B.n41 163.367
R202 B.n172 B.n41 163.367
R203 B.n172 B.n171 163.367
R204 B.n171 B.n170 163.367
R205 B.n170 B.n43 163.367
R206 B.n166 B.n43 163.367
R207 B.n166 B.n165 163.367
R208 B.n165 B.n164 163.367
R209 B.n164 B.n45 163.367
R210 B.n160 B.n45 163.367
R211 B.n160 B.n159 163.367
R212 B.n159 B.n158 163.367
R213 B.n158 B.n47 163.367
R214 B.n154 B.n47 163.367
R215 B.n154 B.n153 163.367
R216 B.n153 B.n152 163.367
R217 B.n152 B.n49 163.367
R218 B.n148 B.n49 163.367
R219 B.n250 B.n249 163.367
R220 B.n249 B.n248 163.367
R221 B.n248 B.n13 163.367
R222 B.n244 B.n13 163.367
R223 B.n244 B.n243 163.367
R224 B.n243 B.n242 163.367
R225 B.n242 B.n15 163.367
R226 B.n238 B.n15 163.367
R227 B.n238 B.n237 163.367
R228 B.n237 B.n19 163.367
R229 B.n233 B.n19 163.367
R230 B.n233 B.n232 163.367
R231 B.n232 B.n231 163.367
R232 B.n231 B.n21 163.367
R233 B.n227 B.n21 163.367
R234 B.n227 B.n226 163.367
R235 B.n226 B.n225 163.367
R236 B.n225 B.n23 163.367
R237 B.n220 B.n23 163.367
R238 B.n220 B.n219 163.367
R239 B.n219 B.n218 163.367
R240 B.n218 B.n27 163.367
R241 B.n214 B.n27 163.367
R242 B.n214 B.n213 163.367
R243 B.n213 B.n212 163.367
R244 B.n212 B.n29 163.367
R245 B.n208 B.n29 163.367
R246 B.n254 B.n11 163.367
R247 B.n255 B.n254 163.367
R248 B.n256 B.n255 163.367
R249 B.n256 B.n9 163.367
R250 B.n260 B.n9 163.367
R251 B.n261 B.n260 163.367
R252 B.n262 B.n261 163.367
R253 B.n262 B.n7 163.367
R254 B.n266 B.n7 163.367
R255 B.n267 B.n266 163.367
R256 B.n268 B.n267 163.367
R257 B.n268 B.n5 163.367
R258 B.n272 B.n5 163.367
R259 B.n273 B.n272 163.367
R260 B.n274 B.n273 163.367
R261 B.n274 B.n3 163.367
R262 B.n278 B.n3 163.367
R263 B.n279 B.n278 163.367
R264 B.n76 B.n2 163.367
R265 B.n77 B.n76 163.367
R266 B.n78 B.n77 163.367
R267 B.n78 B.n73 163.367
R268 B.n82 B.n73 163.367
R269 B.n83 B.n82 163.367
R270 B.n84 B.n83 163.367
R271 B.n84 B.n71 163.367
R272 B.n88 B.n71 163.367
R273 B.n89 B.n88 163.367
R274 B.n90 B.n89 163.367
R275 B.n90 B.n69 163.367
R276 B.n94 B.n69 163.367
R277 B.n95 B.n94 163.367
R278 B.n96 B.n95 163.367
R279 B.n96 B.n67 163.367
R280 B.n100 B.n67 163.367
R281 B.n101 B.n100 163.367
R282 B.n116 B.n61 59.5399
R283 B.n132 B.n131 59.5399
R284 B.n222 B.n25 59.5399
R285 B.n18 B.n17 59.5399
R286 B.n149 B.n50 36.3712
R287 B.n252 B.n251 36.3712
R288 B.n209 B.n30 36.3712
R289 B.n103 B.n66 36.3712
R290 B.n61 B.n60 19.2005
R291 B.n131 B.n130 19.2005
R292 B.n25 B.n24 19.2005
R293 B.n17 B.n16 19.2005
R294 B B.n281 18.0485
R295 B.n253 B.n252 10.6151
R296 B.n253 B.n10 10.6151
R297 B.n257 B.n10 10.6151
R298 B.n258 B.n257 10.6151
R299 B.n259 B.n258 10.6151
R300 B.n259 B.n8 10.6151
R301 B.n263 B.n8 10.6151
R302 B.n264 B.n263 10.6151
R303 B.n265 B.n264 10.6151
R304 B.n265 B.n6 10.6151
R305 B.n269 B.n6 10.6151
R306 B.n270 B.n269 10.6151
R307 B.n271 B.n270 10.6151
R308 B.n271 B.n4 10.6151
R309 B.n275 B.n4 10.6151
R310 B.n276 B.n275 10.6151
R311 B.n277 B.n276 10.6151
R312 B.n277 B.n0 10.6151
R313 B.n251 B.n12 10.6151
R314 B.n247 B.n12 10.6151
R315 B.n247 B.n246 10.6151
R316 B.n246 B.n245 10.6151
R317 B.n245 B.n14 10.6151
R318 B.n241 B.n14 10.6151
R319 B.n241 B.n240 10.6151
R320 B.n240 B.n239 10.6151
R321 B.n236 B.n235 10.6151
R322 B.n235 B.n234 10.6151
R323 B.n234 B.n20 10.6151
R324 B.n230 B.n20 10.6151
R325 B.n230 B.n229 10.6151
R326 B.n229 B.n228 10.6151
R327 B.n228 B.n22 10.6151
R328 B.n224 B.n22 10.6151
R329 B.n224 B.n223 10.6151
R330 B.n221 B.n26 10.6151
R331 B.n217 B.n26 10.6151
R332 B.n217 B.n216 10.6151
R333 B.n216 B.n215 10.6151
R334 B.n215 B.n28 10.6151
R335 B.n211 B.n28 10.6151
R336 B.n211 B.n210 10.6151
R337 B.n210 B.n209 10.6151
R338 B.n205 B.n30 10.6151
R339 B.n205 B.n204 10.6151
R340 B.n204 B.n203 10.6151
R341 B.n203 B.n32 10.6151
R342 B.n199 B.n32 10.6151
R343 B.n199 B.n198 10.6151
R344 B.n198 B.n197 10.6151
R345 B.n197 B.n34 10.6151
R346 B.n193 B.n34 10.6151
R347 B.n193 B.n192 10.6151
R348 B.n192 B.n191 10.6151
R349 B.n191 B.n36 10.6151
R350 B.n187 B.n36 10.6151
R351 B.n187 B.n186 10.6151
R352 B.n186 B.n185 10.6151
R353 B.n185 B.n38 10.6151
R354 B.n181 B.n38 10.6151
R355 B.n181 B.n180 10.6151
R356 B.n180 B.n179 10.6151
R357 B.n179 B.n40 10.6151
R358 B.n175 B.n40 10.6151
R359 B.n175 B.n174 10.6151
R360 B.n174 B.n173 10.6151
R361 B.n173 B.n42 10.6151
R362 B.n169 B.n42 10.6151
R363 B.n169 B.n168 10.6151
R364 B.n168 B.n167 10.6151
R365 B.n167 B.n44 10.6151
R366 B.n163 B.n44 10.6151
R367 B.n163 B.n162 10.6151
R368 B.n162 B.n161 10.6151
R369 B.n161 B.n46 10.6151
R370 B.n157 B.n46 10.6151
R371 B.n157 B.n156 10.6151
R372 B.n156 B.n155 10.6151
R373 B.n155 B.n48 10.6151
R374 B.n151 B.n48 10.6151
R375 B.n151 B.n150 10.6151
R376 B.n150 B.n149 10.6151
R377 B.n75 B.n1 10.6151
R378 B.n75 B.n74 10.6151
R379 B.n79 B.n74 10.6151
R380 B.n80 B.n79 10.6151
R381 B.n81 B.n80 10.6151
R382 B.n81 B.n72 10.6151
R383 B.n85 B.n72 10.6151
R384 B.n86 B.n85 10.6151
R385 B.n87 B.n86 10.6151
R386 B.n87 B.n70 10.6151
R387 B.n91 B.n70 10.6151
R388 B.n92 B.n91 10.6151
R389 B.n93 B.n92 10.6151
R390 B.n93 B.n68 10.6151
R391 B.n97 B.n68 10.6151
R392 B.n98 B.n97 10.6151
R393 B.n99 B.n98 10.6151
R394 B.n99 B.n66 10.6151
R395 B.n104 B.n103 10.6151
R396 B.n105 B.n104 10.6151
R397 B.n105 B.n64 10.6151
R398 B.n109 B.n64 10.6151
R399 B.n110 B.n109 10.6151
R400 B.n111 B.n110 10.6151
R401 B.n111 B.n62 10.6151
R402 B.n115 B.n62 10.6151
R403 B.n118 B.n117 10.6151
R404 B.n118 B.n58 10.6151
R405 B.n122 B.n58 10.6151
R406 B.n123 B.n122 10.6151
R407 B.n124 B.n123 10.6151
R408 B.n124 B.n56 10.6151
R409 B.n128 B.n56 10.6151
R410 B.n129 B.n128 10.6151
R411 B.n133 B.n129 10.6151
R412 B.n137 B.n54 10.6151
R413 B.n138 B.n137 10.6151
R414 B.n139 B.n138 10.6151
R415 B.n139 B.n52 10.6151
R416 B.n143 B.n52 10.6151
R417 B.n144 B.n143 10.6151
R418 B.n145 B.n144 10.6151
R419 B.n145 B.n50 10.6151
R420 B.n239 B.n18 9.36635
R421 B.n222 B.n221 9.36635
R422 B.n116 B.n115 9.36635
R423 B.n132 B.n54 9.36635
R424 B.n281 B.n0 8.11757
R425 B.n281 B.n1 8.11757
R426 B.n236 B.n18 1.24928
R427 B.n223 B.n222 1.24928
R428 B.n117 B.n116 1.24928
R429 B.n133 B.n132 1.24928
R430 VN.n5 VN.n4 161.3
R431 VN.n11 VN.n10 161.3
R432 VN.n9 VN.n6 161.3
R433 VN.n3 VN.n0 161.3
R434 VN.n1 VN.t1 118.29
R435 VN.n7 VN.t3 118.29
R436 VN.n2 VN.t2 97.496
R437 VN.n4 VN.t0 97.496
R438 VN.n8 VN.t4 97.496
R439 VN.n10 VN.t5 97.496
R440 VN.n7 VN.n6 44.8515
R441 VN.n1 VN.n0 44.8515
R442 VN VN.n11 33.0668
R443 VN.n3 VN.n2 24.8308
R444 VN.n9 VN.n8 24.8308
R445 VN.n4 VN.n3 23.3702
R446 VN.n10 VN.n9 23.3702
R447 VN.n2 VN.n1 21.148
R448 VN.n8 VN.n7 21.148
R449 VN.n11 VN.n6 0.189894
R450 VN.n5 VN.n0 0.189894
R451 VN VN.n5 0.0516364
R452 VTAIL.n11 VTAIL.t8 370.971
R453 VTAIL.n2 VTAIL.t0 370.971
R454 VTAIL.n10 VTAIL.t1 370.971
R455 VTAIL.n7 VTAIL.t5 370.971
R456 VTAIL.n1 VTAIL.n0 328.034
R457 VTAIL.n4 VTAIL.n3 328.034
R458 VTAIL.n9 VTAIL.n8 328.033
R459 VTAIL.n6 VTAIL.n5 328.033
R460 VTAIL.n0 VTAIL.t3 31.8681
R461 VTAIL.n0 VTAIL.t6 31.8681
R462 VTAIL.n3 VTAIL.t9 31.8681
R463 VTAIL.n3 VTAIL.t2 31.8681
R464 VTAIL.n8 VTAIL.t10 31.8681
R465 VTAIL.n8 VTAIL.t11 31.8681
R466 VTAIL.n5 VTAIL.t7 31.8681
R467 VTAIL.n5 VTAIL.t4 31.8681
R468 VTAIL.n6 VTAIL.n4 14.9531
R469 VTAIL.n11 VTAIL.n10 14.0996
R470 VTAIL.n9 VTAIL.n7 0.897052
R471 VTAIL.n2 VTAIL.n1 0.897052
R472 VTAIL.n7 VTAIL.n6 0.853948
R473 VTAIL.n10 VTAIL.n9 0.853948
R474 VTAIL.n4 VTAIL.n2 0.853948
R475 VTAIL VTAIL.n11 0.582397
R476 VTAIL VTAIL.n1 0.272052
R477 VDD2.n1 VDD2.t4 388.235
R478 VDD2.n2 VDD2.t0 387.649
R479 VDD2.n1 VDD2.n0 344.87
R480 VDD2 VDD2.n3 344.868
R481 VDD2.n3 VDD2.t1 31.8681
R482 VDD2.n3 VDD2.t2 31.8681
R483 VDD2.n0 VDD2.t3 31.8681
R484 VDD2.n0 VDD2.t5 31.8681
R485 VDD2.n2 VDD2.n1 27.3683
R486 VDD2 VDD2.n2 0.698776
R487 VP.n15 VP.n14 161.3
R488 VP.n5 VP.n2 161.3
R489 VP.n7 VP.n6 161.3
R490 VP.n13 VP.n0 161.3
R491 VP.n12 VP.n11 161.3
R492 VP.n10 VP.n1 161.3
R493 VP.n9 VP.n8 161.3
R494 VP.n3 VP.t1 118.29
R495 VP.n8 VP.t0 97.496
R496 VP.n12 VP.t5 97.496
R497 VP.n14 VP.t4 97.496
R498 VP.n6 VP.t3 97.496
R499 VP.n4 VP.t2 97.496
R500 VP.n3 VP.n2 44.8515
R501 VP.n9 VP.n7 32.6861
R502 VP.n12 VP.n1 24.8308
R503 VP.n13 VP.n12 24.8308
R504 VP.n5 VP.n4 24.8308
R505 VP.n8 VP.n1 23.3702
R506 VP.n14 VP.n13 23.3702
R507 VP.n6 VP.n5 23.3702
R508 VP.n4 VP.n3 21.148
R509 VP.n7 VP.n2 0.189894
R510 VP.n10 VP.n9 0.189894
R511 VP.n11 VP.n10 0.189894
R512 VP.n11 VP.n0 0.189894
R513 VP.n15 VP.n0 0.189894
R514 VP VP.n15 0.0516364
R515 VDD1 VDD1.t4 388.349
R516 VDD1.n1 VDD1.t5 388.235
R517 VDD1.n1 VDD1.n0 344.87
R518 VDD1.n3 VDD1.n2 344.712
R519 VDD1.n2 VDD1.t3 31.8681
R520 VDD1.n2 VDD1.t2 31.8681
R521 VDD1.n0 VDD1.t0 31.8681
R522 VDD1.n0 VDD1.t1 31.8681
R523 VDD1.n3 VDD1.n1 28.378
R524 VDD1 VDD1.n3 0.155672
C0 VDD2 VDD1 0.691731f
C1 VP B 0.960135f
C2 VTAIL w_n1762_n1172# 1.10904f
C3 VTAIL VN 0.934528f
C4 VDD2 VTAIL 2.58706f
C5 w_n1762_n1172# B 3.90068f
C6 VN B 0.59982f
C7 VP w_n1762_n1172# 2.84335f
C8 VDD2 B 0.776648f
C9 VTAIL VDD1 2.54716f
C10 VP VN 3.02352f
C11 VDD2 VP 0.300895f
C12 VDD1 B 0.748335f
C13 VDD1 VP 0.81317f
C14 VN w_n1762_n1172# 2.62861f
C15 VDD2 w_n1762_n1172# 0.996447f
C16 VTAIL B 0.677552f
C17 VDD2 VN 0.669458f
C18 VTAIL VP 0.948678f
C19 VDD1 w_n1762_n1172# 0.974684f
C20 VDD1 VN 0.155324f
C21 VDD2 VSUBS 0.618112f
C22 VDD1 VSUBS 0.839163f
C23 VTAIL VSUBS 0.266764f
C24 VN VSUBS 3.28484f
C25 VP VSUBS 0.927329f
C26 B VSUBS 1.700013f
C27 w_n1762_n1172# VSUBS 26.6203f
C28 VDD1.t4 VSUBS 0.078265f
C29 VDD1.t5 VSUBS 0.078202f
C30 VDD1.t0 VSUBS 0.014282f
C31 VDD1.t1 VSUBS 0.014282f
C32 VDD1.n0 VSUBS 0.047371f
C33 VDD1.n1 VSUBS 1.00491f
C34 VDD1.t3 VSUBS 0.014282f
C35 VDD1.t2 VSUBS 0.014282f
C36 VDD1.n2 VSUBS 0.047278f
C37 VDD1.n3 VSUBS 0.949444f
C38 VP.n0 VSUBS 0.065046f
C39 VP.n1 VSUBS 0.01476f
C40 VP.n2 VSUBS 0.26453f
C41 VP.t3 VSUBS 0.148785f
C42 VP.t2 VSUBS 0.148785f
C43 VP.t1 VSUBS 0.174558f
C44 VP.n3 VSUBS 0.127245f
C45 VP.n4 VSUBS 0.153207f
C46 VP.n5 VSUBS 0.01476f
C47 VP.n6 VSUBS 0.141488f
C48 VP.n7 VSUBS 1.69098f
C49 VP.t0 VSUBS 0.148785f
C50 VP.n8 VSUBS 0.141488f
C51 VP.n9 VSUBS 1.76231f
C52 VP.n10 VSUBS 0.065046f
C53 VP.n11 VSUBS 0.065046f
C54 VP.t5 VSUBS 0.148785f
C55 VP.n12 VSUBS 0.148707f
C56 VP.n13 VSUBS 0.01476f
C57 VP.t4 VSUBS 0.148785f
C58 VP.n14 VSUBS 0.141488f
C59 VP.n15 VSUBS 0.050408f
C60 VDD2.t4 VSUBS 0.083516f
C61 VDD2.t3 VSUBS 0.015253f
C62 VDD2.t5 VSUBS 0.015253f
C63 VDD2.n0 VSUBS 0.05059f
C64 VDD2.n1 VSUBS 1.01989f
C65 VDD2.t0 VSUBS 0.083221f
C66 VDD2.n2 VSUBS 0.98733f
C67 VDD2.t1 VSUBS 0.015253f
C68 VDD2.t2 VSUBS 0.015253f
C69 VDD2.n3 VSUBS 0.050587f
C70 VTAIL.t3 VSUBS 0.02037f
C71 VTAIL.t6 VSUBS 0.02037f
C72 VTAIL.n0 VSUBS 0.05798f
C73 VTAIL.n1 VSUBS 0.260921f
C74 VTAIL.t0 VSUBS 0.102252f
C75 VTAIL.n2 VSUBS 0.319589f
C76 VTAIL.t9 VSUBS 0.02037f
C77 VTAIL.t2 VSUBS 0.02037f
C78 VTAIL.n3 VSUBS 0.05798f
C79 VTAIL.n4 VSUBS 0.789188f
C80 VTAIL.t7 VSUBS 0.02037f
C81 VTAIL.t4 VSUBS 0.02037f
C82 VTAIL.n5 VSUBS 0.05798f
C83 VTAIL.n6 VSUBS 0.789188f
C84 VTAIL.t5 VSUBS 0.102252f
C85 VTAIL.n7 VSUBS 0.319589f
C86 VTAIL.t10 VSUBS 0.02037f
C87 VTAIL.t11 VSUBS 0.02037f
C88 VTAIL.n8 VSUBS 0.05798f
C89 VTAIL.n9 VSUBS 0.308306f
C90 VTAIL.t1 VSUBS 0.102252f
C91 VTAIL.n10 VSUBS 0.730972f
C92 VTAIL.t8 VSUBS 0.102252f
C93 VTAIL.n11 VSUBS 0.708859f
C94 VN.n0 VSUBS 0.251444f
C95 VN.t1 VSUBS 0.165923f
C96 VN.n1 VSUBS 0.120951f
C97 VN.t2 VSUBS 0.141425f
C98 VN.n2 VSUBS 0.145628f
C99 VN.n3 VSUBS 0.01403f
C100 VN.t0 VSUBS 0.141425f
C101 VN.n4 VSUBS 0.134489f
C102 VN.n5 VSUBS 0.047915f
C103 VN.n6 VSUBS 0.251444f
C104 VN.t3 VSUBS 0.165923f
C105 VN.n7 VSUBS 0.120951f
C106 VN.t4 VSUBS 0.141425f
C107 VN.n8 VSUBS 0.145628f
C108 VN.n9 VSUBS 0.01403f
C109 VN.t5 VSUBS 0.141425f
C110 VN.n10 VSUBS 0.134489f
C111 VN.n11 VSUBS 1.64864f
C112 B.n0 VSUBS 0.00876f
C113 B.n1 VSUBS 0.00876f
C114 B.n2 VSUBS 0.012956f
C115 B.n3 VSUBS 0.009928f
C116 B.n4 VSUBS 0.009928f
C117 B.n5 VSUBS 0.009928f
C118 B.n6 VSUBS 0.009928f
C119 B.n7 VSUBS 0.009928f
C120 B.n8 VSUBS 0.009928f
C121 B.n9 VSUBS 0.009928f
C122 B.n10 VSUBS 0.009928f
C123 B.n11 VSUBS 0.024337f
C124 B.n12 VSUBS 0.009928f
C125 B.n13 VSUBS 0.009928f
C126 B.n14 VSUBS 0.009928f
C127 B.n15 VSUBS 0.009928f
C128 B.t7 VSUBS 0.027195f
C129 B.t8 VSUBS 0.029246f
C130 B.t6 VSUBS 0.048916f
C131 B.n16 VSUBS 0.057045f
C132 B.n17 VSUBS 0.054841f
C133 B.n18 VSUBS 0.023002f
C134 B.n19 VSUBS 0.009928f
C135 B.n20 VSUBS 0.009928f
C136 B.n21 VSUBS 0.009928f
C137 B.n22 VSUBS 0.009928f
C138 B.n23 VSUBS 0.009928f
C139 B.t10 VSUBS 0.027195f
C140 B.t11 VSUBS 0.029246f
C141 B.t9 VSUBS 0.048916f
C142 B.n24 VSUBS 0.057045f
C143 B.n25 VSUBS 0.054841f
C144 B.n26 VSUBS 0.009928f
C145 B.n27 VSUBS 0.009928f
C146 B.n28 VSUBS 0.009928f
C147 B.n29 VSUBS 0.009928f
C148 B.n30 VSUBS 0.024337f
C149 B.n31 VSUBS 0.009928f
C150 B.n32 VSUBS 0.009928f
C151 B.n33 VSUBS 0.009928f
C152 B.n34 VSUBS 0.009928f
C153 B.n35 VSUBS 0.009928f
C154 B.n36 VSUBS 0.009928f
C155 B.n37 VSUBS 0.009928f
C156 B.n38 VSUBS 0.009928f
C157 B.n39 VSUBS 0.009928f
C158 B.n40 VSUBS 0.009928f
C159 B.n41 VSUBS 0.009928f
C160 B.n42 VSUBS 0.009928f
C161 B.n43 VSUBS 0.009928f
C162 B.n44 VSUBS 0.009928f
C163 B.n45 VSUBS 0.009928f
C164 B.n46 VSUBS 0.009928f
C165 B.n47 VSUBS 0.009928f
C166 B.n48 VSUBS 0.009928f
C167 B.n49 VSUBS 0.009928f
C168 B.n50 VSUBS 0.024542f
C169 B.n51 VSUBS 0.009928f
C170 B.n52 VSUBS 0.009928f
C171 B.n53 VSUBS 0.009928f
C172 B.n54 VSUBS 0.009344f
C173 B.n55 VSUBS 0.009928f
C174 B.n56 VSUBS 0.009928f
C175 B.n57 VSUBS 0.009928f
C176 B.n58 VSUBS 0.009928f
C177 B.n59 VSUBS 0.009928f
C178 B.t5 VSUBS 0.027195f
C179 B.t4 VSUBS 0.029246f
C180 B.t3 VSUBS 0.048916f
C181 B.n60 VSUBS 0.057045f
C182 B.n61 VSUBS 0.054841f
C183 B.n62 VSUBS 0.009928f
C184 B.n63 VSUBS 0.009928f
C185 B.n64 VSUBS 0.009928f
C186 B.n65 VSUBS 0.009928f
C187 B.n66 VSUBS 0.024337f
C188 B.n67 VSUBS 0.009928f
C189 B.n68 VSUBS 0.009928f
C190 B.n69 VSUBS 0.009928f
C191 B.n70 VSUBS 0.009928f
C192 B.n71 VSUBS 0.009928f
C193 B.n72 VSUBS 0.009928f
C194 B.n73 VSUBS 0.009928f
C195 B.n74 VSUBS 0.009928f
C196 B.n75 VSUBS 0.009928f
C197 B.n76 VSUBS 0.009928f
C198 B.n77 VSUBS 0.009928f
C199 B.n78 VSUBS 0.009928f
C200 B.n79 VSUBS 0.009928f
C201 B.n80 VSUBS 0.009928f
C202 B.n81 VSUBS 0.009928f
C203 B.n82 VSUBS 0.009928f
C204 B.n83 VSUBS 0.009928f
C205 B.n84 VSUBS 0.009928f
C206 B.n85 VSUBS 0.009928f
C207 B.n86 VSUBS 0.009928f
C208 B.n87 VSUBS 0.009928f
C209 B.n88 VSUBS 0.009928f
C210 B.n89 VSUBS 0.009928f
C211 B.n90 VSUBS 0.009928f
C212 B.n91 VSUBS 0.009928f
C213 B.n92 VSUBS 0.009928f
C214 B.n93 VSUBS 0.009928f
C215 B.n94 VSUBS 0.009928f
C216 B.n95 VSUBS 0.009928f
C217 B.n96 VSUBS 0.009928f
C218 B.n97 VSUBS 0.009928f
C219 B.n98 VSUBS 0.009928f
C220 B.n99 VSUBS 0.009928f
C221 B.n100 VSUBS 0.009928f
C222 B.n101 VSUBS 0.024337f
C223 B.n102 VSUBS 0.025596f
C224 B.n103 VSUBS 0.025596f
C225 B.n104 VSUBS 0.009928f
C226 B.n105 VSUBS 0.009928f
C227 B.n106 VSUBS 0.009928f
C228 B.n107 VSUBS 0.009928f
C229 B.n108 VSUBS 0.009928f
C230 B.n109 VSUBS 0.009928f
C231 B.n110 VSUBS 0.009928f
C232 B.n111 VSUBS 0.009928f
C233 B.n112 VSUBS 0.009928f
C234 B.n113 VSUBS 0.009928f
C235 B.n114 VSUBS 0.009928f
C236 B.n115 VSUBS 0.009344f
C237 B.n116 VSUBS 0.023002f
C238 B.n117 VSUBS 0.005548f
C239 B.n118 VSUBS 0.009928f
C240 B.n119 VSUBS 0.009928f
C241 B.n120 VSUBS 0.009928f
C242 B.n121 VSUBS 0.009928f
C243 B.n122 VSUBS 0.009928f
C244 B.n123 VSUBS 0.009928f
C245 B.n124 VSUBS 0.009928f
C246 B.n125 VSUBS 0.009928f
C247 B.n126 VSUBS 0.009928f
C248 B.n127 VSUBS 0.009928f
C249 B.n128 VSUBS 0.009928f
C250 B.n129 VSUBS 0.009928f
C251 B.t2 VSUBS 0.027195f
C252 B.t1 VSUBS 0.029246f
C253 B.t0 VSUBS 0.048916f
C254 B.n130 VSUBS 0.057045f
C255 B.n131 VSUBS 0.054841f
C256 B.n132 VSUBS 0.023002f
C257 B.n133 VSUBS 0.005548f
C258 B.n134 VSUBS 0.009928f
C259 B.n135 VSUBS 0.009928f
C260 B.n136 VSUBS 0.009928f
C261 B.n137 VSUBS 0.009928f
C262 B.n138 VSUBS 0.009928f
C263 B.n139 VSUBS 0.009928f
C264 B.n140 VSUBS 0.009928f
C265 B.n141 VSUBS 0.009928f
C266 B.n142 VSUBS 0.009928f
C267 B.n143 VSUBS 0.009928f
C268 B.n144 VSUBS 0.009928f
C269 B.n145 VSUBS 0.009928f
C270 B.n146 VSUBS 0.009928f
C271 B.n147 VSUBS 0.025596f
C272 B.n148 VSUBS 0.024337f
C273 B.n149 VSUBS 0.02539f
C274 B.n150 VSUBS 0.009928f
C275 B.n151 VSUBS 0.009928f
C276 B.n152 VSUBS 0.009928f
C277 B.n153 VSUBS 0.009928f
C278 B.n154 VSUBS 0.009928f
C279 B.n155 VSUBS 0.009928f
C280 B.n156 VSUBS 0.009928f
C281 B.n157 VSUBS 0.009928f
C282 B.n158 VSUBS 0.009928f
C283 B.n159 VSUBS 0.009928f
C284 B.n160 VSUBS 0.009928f
C285 B.n161 VSUBS 0.009928f
C286 B.n162 VSUBS 0.009928f
C287 B.n163 VSUBS 0.009928f
C288 B.n164 VSUBS 0.009928f
C289 B.n165 VSUBS 0.009928f
C290 B.n166 VSUBS 0.009928f
C291 B.n167 VSUBS 0.009928f
C292 B.n168 VSUBS 0.009928f
C293 B.n169 VSUBS 0.009928f
C294 B.n170 VSUBS 0.009928f
C295 B.n171 VSUBS 0.009928f
C296 B.n172 VSUBS 0.009928f
C297 B.n173 VSUBS 0.009928f
C298 B.n174 VSUBS 0.009928f
C299 B.n175 VSUBS 0.009928f
C300 B.n176 VSUBS 0.009928f
C301 B.n177 VSUBS 0.009928f
C302 B.n178 VSUBS 0.009928f
C303 B.n179 VSUBS 0.009928f
C304 B.n180 VSUBS 0.009928f
C305 B.n181 VSUBS 0.009928f
C306 B.n182 VSUBS 0.009928f
C307 B.n183 VSUBS 0.009928f
C308 B.n184 VSUBS 0.009928f
C309 B.n185 VSUBS 0.009928f
C310 B.n186 VSUBS 0.009928f
C311 B.n187 VSUBS 0.009928f
C312 B.n188 VSUBS 0.009928f
C313 B.n189 VSUBS 0.009928f
C314 B.n190 VSUBS 0.009928f
C315 B.n191 VSUBS 0.009928f
C316 B.n192 VSUBS 0.009928f
C317 B.n193 VSUBS 0.009928f
C318 B.n194 VSUBS 0.009928f
C319 B.n195 VSUBS 0.009928f
C320 B.n196 VSUBS 0.009928f
C321 B.n197 VSUBS 0.009928f
C322 B.n198 VSUBS 0.009928f
C323 B.n199 VSUBS 0.009928f
C324 B.n200 VSUBS 0.009928f
C325 B.n201 VSUBS 0.009928f
C326 B.n202 VSUBS 0.009928f
C327 B.n203 VSUBS 0.009928f
C328 B.n204 VSUBS 0.009928f
C329 B.n205 VSUBS 0.009928f
C330 B.n206 VSUBS 0.009928f
C331 B.n207 VSUBS 0.024337f
C332 B.n208 VSUBS 0.025596f
C333 B.n209 VSUBS 0.025596f
C334 B.n210 VSUBS 0.009928f
C335 B.n211 VSUBS 0.009928f
C336 B.n212 VSUBS 0.009928f
C337 B.n213 VSUBS 0.009928f
C338 B.n214 VSUBS 0.009928f
C339 B.n215 VSUBS 0.009928f
C340 B.n216 VSUBS 0.009928f
C341 B.n217 VSUBS 0.009928f
C342 B.n218 VSUBS 0.009928f
C343 B.n219 VSUBS 0.009928f
C344 B.n220 VSUBS 0.009928f
C345 B.n221 VSUBS 0.009344f
C346 B.n222 VSUBS 0.023002f
C347 B.n223 VSUBS 0.005548f
C348 B.n224 VSUBS 0.009928f
C349 B.n225 VSUBS 0.009928f
C350 B.n226 VSUBS 0.009928f
C351 B.n227 VSUBS 0.009928f
C352 B.n228 VSUBS 0.009928f
C353 B.n229 VSUBS 0.009928f
C354 B.n230 VSUBS 0.009928f
C355 B.n231 VSUBS 0.009928f
C356 B.n232 VSUBS 0.009928f
C357 B.n233 VSUBS 0.009928f
C358 B.n234 VSUBS 0.009928f
C359 B.n235 VSUBS 0.009928f
C360 B.n236 VSUBS 0.005548f
C361 B.n237 VSUBS 0.009928f
C362 B.n238 VSUBS 0.009928f
C363 B.n239 VSUBS 0.009344f
C364 B.n240 VSUBS 0.009928f
C365 B.n241 VSUBS 0.009928f
C366 B.n242 VSUBS 0.009928f
C367 B.n243 VSUBS 0.009928f
C368 B.n244 VSUBS 0.009928f
C369 B.n245 VSUBS 0.009928f
C370 B.n246 VSUBS 0.009928f
C371 B.n247 VSUBS 0.009928f
C372 B.n248 VSUBS 0.009928f
C373 B.n249 VSUBS 0.009928f
C374 B.n250 VSUBS 0.025596f
C375 B.n251 VSUBS 0.025596f
C376 B.n252 VSUBS 0.024337f
C377 B.n253 VSUBS 0.009928f
C378 B.n254 VSUBS 0.009928f
C379 B.n255 VSUBS 0.009928f
C380 B.n256 VSUBS 0.009928f
C381 B.n257 VSUBS 0.009928f
C382 B.n258 VSUBS 0.009928f
C383 B.n259 VSUBS 0.009928f
C384 B.n260 VSUBS 0.009928f
C385 B.n261 VSUBS 0.009928f
C386 B.n262 VSUBS 0.009928f
C387 B.n263 VSUBS 0.009928f
C388 B.n264 VSUBS 0.009928f
C389 B.n265 VSUBS 0.009928f
C390 B.n266 VSUBS 0.009928f
C391 B.n267 VSUBS 0.009928f
C392 B.n268 VSUBS 0.009928f
C393 B.n269 VSUBS 0.009928f
C394 B.n270 VSUBS 0.009928f
C395 B.n271 VSUBS 0.009928f
C396 B.n272 VSUBS 0.009928f
C397 B.n273 VSUBS 0.009928f
C398 B.n274 VSUBS 0.009928f
C399 B.n275 VSUBS 0.009928f
C400 B.n276 VSUBS 0.009928f
C401 B.n277 VSUBS 0.009928f
C402 B.n278 VSUBS 0.009928f
C403 B.n279 VSUBS 0.012956f
C404 B.n280 VSUBS 0.013801f
C405 B.n281 VSUBS 0.027445f
.ends

