* NGSPICE file created from diff_pair_sample_0660.ext - technology: sky130A

.subckt diff_pair_sample_0660 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t2 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X1 VDD2.t9 VN.t0 VTAIL.t1 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0.83325 ps=5.38 w=5.05 l=0.71
X2 B.t11 B.t9 B.t10 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0 ps=0 w=5.05 l=0.71
X3 VDD2.t8 VN.t1 VTAIL.t5 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X4 VTAIL.t18 VP.t1 VDD1.t5 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X5 VTAIL.t6 VN.t2 VDD2.t7 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X6 VTAIL.t17 VP.t2 VDD1.t3 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X7 VTAIL.t3 VN.t3 VDD2.t6 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X8 VTAIL.t4 VN.t4 VDD2.t5 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X9 B.t8 B.t6 B.t7 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0 ps=0 w=5.05 l=0.71
X10 VDD2.t4 VN.t5 VTAIL.t7 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=1.9695 ps=10.88 w=5.05 l=0.71
X11 VDD1.t1 VP.t3 VTAIL.t16 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0.83325 ps=5.38 w=5.05 l=0.71
X12 VDD1.t0 VP.t4 VTAIL.t15 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0.83325 ps=5.38 w=5.05 l=0.71
X13 B.t5 B.t3 B.t4 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0 ps=0 w=5.05 l=0.71
X14 VDD1.t6 VP.t5 VTAIL.t14 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=1.9695 ps=10.88 w=5.05 l=0.71
X15 VDD2.t3 VN.t6 VTAIL.t0 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=1.9695 ps=10.88 w=5.05 l=0.71
X16 VTAIL.t13 VP.t6 VDD1.t4 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X17 VDD2.t2 VN.t7 VTAIL.t8 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X18 B.t2 B.t0 B.t1 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0 ps=0 w=5.05 l=0.71
X19 VDD2.t1 VN.t8 VTAIL.t9 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=1.9695 pd=10.88 as=0.83325 ps=5.38 w=5.05 l=0.71
X20 VDD1.t9 VP.t7 VTAIL.t12 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=1.9695 ps=10.88 w=5.05 l=0.71
X21 VTAIL.t2 VN.t9 VDD2.t0 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X22 VDD1.t8 VP.t8 VTAIL.t11 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
X23 VDD1.t7 VP.t9 VTAIL.t10 w_n2218_n1978# sky130_fd_pr__pfet_01v8 ad=0.83325 pd=5.38 as=0.83325 ps=5.38 w=5.05 l=0.71
R0 VP.n7 VP.t4 250.387
R1 VP.n18 VP.t3 227.083
R2 VP.n22 VP.t2 227.083
R3 VP.n24 VP.t9 227.083
R4 VP.n28 VP.t6 227.083
R5 VP.n30 VP.t5 227.083
R6 VP.n16 VP.t7 227.083
R7 VP.n14 VP.t0 227.083
R8 VP.n6 VP.t8 227.083
R9 VP.n8 VP.t1 227.083
R10 VP.n31 VP.n30 161.3
R11 VP.n10 VP.n9 161.3
R12 VP.n11 VP.n6 161.3
R13 VP.n13 VP.n12 161.3
R14 VP.n14 VP.n5 161.3
R15 VP.n15 VP.n4 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n29 VP.n0 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.n1 161.3
R20 VP.n25 VP.n24 161.3
R21 VP.n23 VP.n2 161.3
R22 VP.n22 VP.n21 161.3
R23 VP.n20 VP.n3 161.3
R24 VP.n19 VP.n18 161.3
R25 VP.n10 VP.n7 44.8907
R26 VP.n19 VP.n17 37.5914
R27 VP.n18 VP.n3 32.8641
R28 VP.n30 VP.n29 32.8641
R29 VP.n16 VP.n15 32.8641
R30 VP.n23 VP.n22 27.0217
R31 VP.n28 VP.n1 27.0217
R32 VP.n14 VP.n13 27.0217
R33 VP.n9 VP.n8 27.0217
R34 VP.n24 VP.n23 21.1793
R35 VP.n24 VP.n1 21.1793
R36 VP.n13 VP.n6 21.1793
R37 VP.n9 VP.n6 21.1793
R38 VP.n8 VP.n7 18.4104
R39 VP.n22 VP.n3 15.3369
R40 VP.n29 VP.n28 15.3369
R41 VP.n15 VP.n14 15.3369
R42 VP.n11 VP.n10 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n5 0.189894
R45 VP.n5 VP.n4 0.189894
R46 VP.n17 VP.n4 0.189894
R47 VP.n20 VP.n19 0.189894
R48 VP.n21 VP.n20 0.189894
R49 VP.n21 VP.n2 0.189894
R50 VP.n25 VP.n2 0.189894
R51 VP.n26 VP.n25 0.189894
R52 VP.n27 VP.n26 0.189894
R53 VP.n27 VP.n0 0.189894
R54 VP.n31 VP.n0 0.189894
R55 VP VP.n31 0.0516364
R56 VDD1.n1 VDD1.t0 110.296
R57 VDD1.n3 VDD1.t1 110.296
R58 VDD1.n5 VDD1.n4 103.579
R59 VDD1.n1 VDD1.n0 102.963
R60 VDD1.n7 VDD1.n6 102.962
R61 VDD1.n3 VDD1.n2 102.962
R62 VDD1.n7 VDD1.n5 33.3586
R63 VDD1.n6 VDD1.t2 6.43713
R64 VDD1.n6 VDD1.t9 6.43713
R65 VDD1.n0 VDD1.t5 6.43713
R66 VDD1.n0 VDD1.t8 6.43713
R67 VDD1.n4 VDD1.t4 6.43713
R68 VDD1.n4 VDD1.t6 6.43713
R69 VDD1.n2 VDD1.t3 6.43713
R70 VDD1.n2 VDD1.t7 6.43713
R71 VDD1 VDD1.n7 0.614724
R72 VDD1 VDD1.n1 0.282828
R73 VDD1.n5 VDD1.n3 0.169292
R74 VTAIL.n11 VTAIL.t0 92.7198
R75 VTAIL.n16 VTAIL.t12 92.7197
R76 VTAIL.n17 VTAIL.t7 92.7197
R77 VTAIL.n2 VTAIL.t14 92.7197
R78 VTAIL.n15 VTAIL.n14 86.2832
R79 VTAIL.n13 VTAIL.n12 86.2832
R80 VTAIL.n10 VTAIL.n9 86.2832
R81 VTAIL.n8 VTAIL.n7 86.2832
R82 VTAIL.n19 VTAIL.n18 86.283
R83 VTAIL.n1 VTAIL.n0 86.283
R84 VTAIL.n4 VTAIL.n3 86.283
R85 VTAIL.n6 VTAIL.n5 86.283
R86 VTAIL.n8 VTAIL.n6 18.5134
R87 VTAIL.n17 VTAIL.n16 17.6169
R88 VTAIL.n18 VTAIL.t8 6.43713
R89 VTAIL.n18 VTAIL.t6 6.43713
R90 VTAIL.n0 VTAIL.t1 6.43713
R91 VTAIL.n0 VTAIL.t3 6.43713
R92 VTAIL.n3 VTAIL.t10 6.43713
R93 VTAIL.n3 VTAIL.t13 6.43713
R94 VTAIL.n5 VTAIL.t16 6.43713
R95 VTAIL.n5 VTAIL.t17 6.43713
R96 VTAIL.n14 VTAIL.t11 6.43713
R97 VTAIL.n14 VTAIL.t19 6.43713
R98 VTAIL.n12 VTAIL.t15 6.43713
R99 VTAIL.n12 VTAIL.t18 6.43713
R100 VTAIL.n9 VTAIL.t5 6.43713
R101 VTAIL.n9 VTAIL.t4 6.43713
R102 VTAIL.n7 VTAIL.t9 6.43713
R103 VTAIL.n7 VTAIL.t2 6.43713
R104 VTAIL.n13 VTAIL.n11 0.918603
R105 VTAIL.n2 VTAIL.n1 0.918603
R106 VTAIL.n10 VTAIL.n8 0.897052
R107 VTAIL.n11 VTAIL.n10 0.897052
R108 VTAIL.n15 VTAIL.n13 0.897052
R109 VTAIL.n16 VTAIL.n15 0.897052
R110 VTAIL.n6 VTAIL.n4 0.897052
R111 VTAIL.n4 VTAIL.n2 0.897052
R112 VTAIL.n19 VTAIL.n17 0.897052
R113 VTAIL VTAIL.n1 0.731103
R114 VTAIL VTAIL.n19 0.166448
R115 VN.n3 VN.t0 250.387
R116 VN.n17 VN.t6 250.387
R117 VN.n4 VN.t3 227.083
R118 VN.n6 VN.t7 227.083
R119 VN.n10 VN.t2 227.083
R120 VN.n12 VN.t5 227.083
R121 VN.n18 VN.t4 227.083
R122 VN.n20 VN.t1 227.083
R123 VN.n24 VN.t9 227.083
R124 VN.n26 VN.t8 227.083
R125 VN.n13 VN.n12 161.3
R126 VN.n27 VN.n26 161.3
R127 VN.n25 VN.n14 161.3
R128 VN.n24 VN.n23 161.3
R129 VN.n22 VN.n15 161.3
R130 VN.n21 VN.n20 161.3
R131 VN.n19 VN.n16 161.3
R132 VN.n11 VN.n0 161.3
R133 VN.n10 VN.n9 161.3
R134 VN.n8 VN.n1 161.3
R135 VN.n7 VN.n6 161.3
R136 VN.n5 VN.n2 161.3
R137 VN.n17 VN.n16 44.8907
R138 VN.n3 VN.n2 44.8907
R139 VN VN.n27 37.9721
R140 VN.n12 VN.n11 32.8641
R141 VN.n26 VN.n25 32.8641
R142 VN.n5 VN.n4 27.0217
R143 VN.n10 VN.n1 27.0217
R144 VN.n19 VN.n18 27.0217
R145 VN.n24 VN.n15 27.0217
R146 VN.n6 VN.n5 21.1793
R147 VN.n6 VN.n1 21.1793
R148 VN.n20 VN.n19 21.1793
R149 VN.n20 VN.n15 21.1793
R150 VN.n4 VN.n3 18.4104
R151 VN.n18 VN.n17 18.4104
R152 VN.n11 VN.n10 15.3369
R153 VN.n25 VN.n24 15.3369
R154 VN.n27 VN.n14 0.189894
R155 VN.n23 VN.n14 0.189894
R156 VN.n23 VN.n22 0.189894
R157 VN.n22 VN.n21 0.189894
R158 VN.n21 VN.n16 0.189894
R159 VN.n7 VN.n2 0.189894
R160 VN.n8 VN.n7 0.189894
R161 VN.n9 VN.n8 0.189894
R162 VN.n9 VN.n0 0.189894
R163 VN.n13 VN.n0 0.189894
R164 VN VN.n13 0.0516364
R165 VDD2.n1 VDD2.t9 110.296
R166 VDD2.n4 VDD2.t1 109.398
R167 VDD2.n3 VDD2.n2 103.579
R168 VDD2 VDD2.n7 103.576
R169 VDD2.n6 VDD2.n5 102.963
R170 VDD2.n1 VDD2.n0 102.962
R171 VDD2.n4 VDD2.n3 32.3274
R172 VDD2.n7 VDD2.t5 6.43713
R173 VDD2.n7 VDD2.t3 6.43713
R174 VDD2.n5 VDD2.t0 6.43713
R175 VDD2.n5 VDD2.t8 6.43713
R176 VDD2.n2 VDD2.t7 6.43713
R177 VDD2.n2 VDD2.t4 6.43713
R178 VDD2.n0 VDD2.t6 6.43713
R179 VDD2.n0 VDD2.t2 6.43713
R180 VDD2.n6 VDD2.n4 0.897052
R181 VDD2 VDD2.n6 0.282828
R182 VDD2.n3 VDD2.n1 0.169292
R183 B.n232 B.n73 585
R184 B.n231 B.n230 585
R185 B.n229 B.n74 585
R186 B.n228 B.n227 585
R187 B.n226 B.n75 585
R188 B.n225 B.n224 585
R189 B.n223 B.n76 585
R190 B.n222 B.n221 585
R191 B.n220 B.n77 585
R192 B.n219 B.n218 585
R193 B.n217 B.n78 585
R194 B.n216 B.n215 585
R195 B.n214 B.n79 585
R196 B.n213 B.n212 585
R197 B.n211 B.n80 585
R198 B.n210 B.n209 585
R199 B.n208 B.n81 585
R200 B.n207 B.n206 585
R201 B.n205 B.n82 585
R202 B.n204 B.n203 585
R203 B.n202 B.n83 585
R204 B.n201 B.n200 585
R205 B.n196 B.n84 585
R206 B.n195 B.n194 585
R207 B.n193 B.n85 585
R208 B.n192 B.n191 585
R209 B.n190 B.n86 585
R210 B.n189 B.n188 585
R211 B.n187 B.n87 585
R212 B.n186 B.n185 585
R213 B.n184 B.n88 585
R214 B.n182 B.n181 585
R215 B.n180 B.n91 585
R216 B.n179 B.n178 585
R217 B.n177 B.n92 585
R218 B.n176 B.n175 585
R219 B.n174 B.n93 585
R220 B.n173 B.n172 585
R221 B.n171 B.n94 585
R222 B.n170 B.n169 585
R223 B.n168 B.n95 585
R224 B.n167 B.n166 585
R225 B.n165 B.n96 585
R226 B.n164 B.n163 585
R227 B.n162 B.n97 585
R228 B.n161 B.n160 585
R229 B.n159 B.n98 585
R230 B.n158 B.n157 585
R231 B.n156 B.n99 585
R232 B.n155 B.n154 585
R233 B.n153 B.n100 585
R234 B.n152 B.n151 585
R235 B.n234 B.n233 585
R236 B.n235 B.n72 585
R237 B.n237 B.n236 585
R238 B.n238 B.n71 585
R239 B.n240 B.n239 585
R240 B.n241 B.n70 585
R241 B.n243 B.n242 585
R242 B.n244 B.n69 585
R243 B.n246 B.n245 585
R244 B.n247 B.n68 585
R245 B.n249 B.n248 585
R246 B.n250 B.n67 585
R247 B.n252 B.n251 585
R248 B.n253 B.n66 585
R249 B.n255 B.n254 585
R250 B.n256 B.n65 585
R251 B.n258 B.n257 585
R252 B.n259 B.n64 585
R253 B.n261 B.n260 585
R254 B.n262 B.n63 585
R255 B.n264 B.n263 585
R256 B.n265 B.n62 585
R257 B.n267 B.n266 585
R258 B.n268 B.n61 585
R259 B.n270 B.n269 585
R260 B.n271 B.n60 585
R261 B.n273 B.n272 585
R262 B.n274 B.n59 585
R263 B.n276 B.n275 585
R264 B.n277 B.n58 585
R265 B.n279 B.n278 585
R266 B.n280 B.n57 585
R267 B.n282 B.n281 585
R268 B.n283 B.n56 585
R269 B.n285 B.n284 585
R270 B.n286 B.n55 585
R271 B.n288 B.n287 585
R272 B.n289 B.n54 585
R273 B.n291 B.n290 585
R274 B.n292 B.n53 585
R275 B.n294 B.n293 585
R276 B.n295 B.n52 585
R277 B.n297 B.n296 585
R278 B.n298 B.n51 585
R279 B.n300 B.n299 585
R280 B.n301 B.n50 585
R281 B.n303 B.n302 585
R282 B.n304 B.n49 585
R283 B.n306 B.n305 585
R284 B.n307 B.n48 585
R285 B.n309 B.n308 585
R286 B.n310 B.n47 585
R287 B.n312 B.n311 585
R288 B.n313 B.n46 585
R289 B.n392 B.n15 585
R290 B.n391 B.n390 585
R291 B.n389 B.n16 585
R292 B.n388 B.n387 585
R293 B.n386 B.n17 585
R294 B.n385 B.n384 585
R295 B.n383 B.n18 585
R296 B.n382 B.n381 585
R297 B.n380 B.n19 585
R298 B.n379 B.n378 585
R299 B.n377 B.n20 585
R300 B.n376 B.n375 585
R301 B.n374 B.n21 585
R302 B.n373 B.n372 585
R303 B.n371 B.n22 585
R304 B.n370 B.n369 585
R305 B.n368 B.n23 585
R306 B.n367 B.n366 585
R307 B.n365 B.n24 585
R308 B.n364 B.n363 585
R309 B.n362 B.n25 585
R310 B.n360 B.n359 585
R311 B.n358 B.n28 585
R312 B.n357 B.n356 585
R313 B.n355 B.n29 585
R314 B.n354 B.n353 585
R315 B.n352 B.n30 585
R316 B.n351 B.n350 585
R317 B.n349 B.n31 585
R318 B.n348 B.n347 585
R319 B.n346 B.n32 585
R320 B.n345 B.n344 585
R321 B.n343 B.n33 585
R322 B.n342 B.n341 585
R323 B.n340 B.n37 585
R324 B.n339 B.n338 585
R325 B.n337 B.n38 585
R326 B.n336 B.n335 585
R327 B.n334 B.n39 585
R328 B.n333 B.n332 585
R329 B.n331 B.n40 585
R330 B.n330 B.n329 585
R331 B.n328 B.n41 585
R332 B.n327 B.n326 585
R333 B.n325 B.n42 585
R334 B.n324 B.n323 585
R335 B.n322 B.n43 585
R336 B.n321 B.n320 585
R337 B.n319 B.n44 585
R338 B.n318 B.n317 585
R339 B.n316 B.n45 585
R340 B.n315 B.n314 585
R341 B.n394 B.n393 585
R342 B.n395 B.n14 585
R343 B.n397 B.n396 585
R344 B.n398 B.n13 585
R345 B.n400 B.n399 585
R346 B.n401 B.n12 585
R347 B.n403 B.n402 585
R348 B.n404 B.n11 585
R349 B.n406 B.n405 585
R350 B.n407 B.n10 585
R351 B.n409 B.n408 585
R352 B.n410 B.n9 585
R353 B.n412 B.n411 585
R354 B.n413 B.n8 585
R355 B.n415 B.n414 585
R356 B.n416 B.n7 585
R357 B.n418 B.n417 585
R358 B.n419 B.n6 585
R359 B.n421 B.n420 585
R360 B.n422 B.n5 585
R361 B.n424 B.n423 585
R362 B.n425 B.n4 585
R363 B.n427 B.n426 585
R364 B.n428 B.n3 585
R365 B.n430 B.n429 585
R366 B.n431 B.n0 585
R367 B.n2 B.n1 585
R368 B.n114 B.n113 585
R369 B.n116 B.n115 585
R370 B.n117 B.n112 585
R371 B.n119 B.n118 585
R372 B.n120 B.n111 585
R373 B.n122 B.n121 585
R374 B.n123 B.n110 585
R375 B.n125 B.n124 585
R376 B.n126 B.n109 585
R377 B.n128 B.n127 585
R378 B.n129 B.n108 585
R379 B.n131 B.n130 585
R380 B.n132 B.n107 585
R381 B.n134 B.n133 585
R382 B.n135 B.n106 585
R383 B.n137 B.n136 585
R384 B.n138 B.n105 585
R385 B.n140 B.n139 585
R386 B.n141 B.n104 585
R387 B.n143 B.n142 585
R388 B.n144 B.n103 585
R389 B.n146 B.n145 585
R390 B.n147 B.n102 585
R391 B.n149 B.n148 585
R392 B.n150 B.n101 585
R393 B.n151 B.n150 487.695
R394 B.n233 B.n232 487.695
R395 B.n315 B.n46 487.695
R396 B.n394 B.n15 487.695
R397 B.n89 B.t9 374.26
R398 B.n197 B.t3 374.26
R399 B.n34 B.t0 374.26
R400 B.n26 B.t6 374.26
R401 B.n433 B.n432 256.663
R402 B.n432 B.n431 235.042
R403 B.n432 B.n2 235.042
R404 B.n151 B.n100 163.367
R405 B.n155 B.n100 163.367
R406 B.n156 B.n155 163.367
R407 B.n157 B.n156 163.367
R408 B.n157 B.n98 163.367
R409 B.n161 B.n98 163.367
R410 B.n162 B.n161 163.367
R411 B.n163 B.n162 163.367
R412 B.n163 B.n96 163.367
R413 B.n167 B.n96 163.367
R414 B.n168 B.n167 163.367
R415 B.n169 B.n168 163.367
R416 B.n169 B.n94 163.367
R417 B.n173 B.n94 163.367
R418 B.n174 B.n173 163.367
R419 B.n175 B.n174 163.367
R420 B.n175 B.n92 163.367
R421 B.n179 B.n92 163.367
R422 B.n180 B.n179 163.367
R423 B.n181 B.n180 163.367
R424 B.n181 B.n88 163.367
R425 B.n186 B.n88 163.367
R426 B.n187 B.n186 163.367
R427 B.n188 B.n187 163.367
R428 B.n188 B.n86 163.367
R429 B.n192 B.n86 163.367
R430 B.n193 B.n192 163.367
R431 B.n194 B.n193 163.367
R432 B.n194 B.n84 163.367
R433 B.n201 B.n84 163.367
R434 B.n202 B.n201 163.367
R435 B.n203 B.n202 163.367
R436 B.n203 B.n82 163.367
R437 B.n207 B.n82 163.367
R438 B.n208 B.n207 163.367
R439 B.n209 B.n208 163.367
R440 B.n209 B.n80 163.367
R441 B.n213 B.n80 163.367
R442 B.n214 B.n213 163.367
R443 B.n215 B.n214 163.367
R444 B.n215 B.n78 163.367
R445 B.n219 B.n78 163.367
R446 B.n220 B.n219 163.367
R447 B.n221 B.n220 163.367
R448 B.n221 B.n76 163.367
R449 B.n225 B.n76 163.367
R450 B.n226 B.n225 163.367
R451 B.n227 B.n226 163.367
R452 B.n227 B.n74 163.367
R453 B.n231 B.n74 163.367
R454 B.n232 B.n231 163.367
R455 B.n311 B.n46 163.367
R456 B.n311 B.n310 163.367
R457 B.n310 B.n309 163.367
R458 B.n309 B.n48 163.367
R459 B.n305 B.n48 163.367
R460 B.n305 B.n304 163.367
R461 B.n304 B.n303 163.367
R462 B.n303 B.n50 163.367
R463 B.n299 B.n50 163.367
R464 B.n299 B.n298 163.367
R465 B.n298 B.n297 163.367
R466 B.n297 B.n52 163.367
R467 B.n293 B.n52 163.367
R468 B.n293 B.n292 163.367
R469 B.n292 B.n291 163.367
R470 B.n291 B.n54 163.367
R471 B.n287 B.n54 163.367
R472 B.n287 B.n286 163.367
R473 B.n286 B.n285 163.367
R474 B.n285 B.n56 163.367
R475 B.n281 B.n56 163.367
R476 B.n281 B.n280 163.367
R477 B.n280 B.n279 163.367
R478 B.n279 B.n58 163.367
R479 B.n275 B.n58 163.367
R480 B.n275 B.n274 163.367
R481 B.n274 B.n273 163.367
R482 B.n273 B.n60 163.367
R483 B.n269 B.n60 163.367
R484 B.n269 B.n268 163.367
R485 B.n268 B.n267 163.367
R486 B.n267 B.n62 163.367
R487 B.n263 B.n62 163.367
R488 B.n263 B.n262 163.367
R489 B.n262 B.n261 163.367
R490 B.n261 B.n64 163.367
R491 B.n257 B.n64 163.367
R492 B.n257 B.n256 163.367
R493 B.n256 B.n255 163.367
R494 B.n255 B.n66 163.367
R495 B.n251 B.n66 163.367
R496 B.n251 B.n250 163.367
R497 B.n250 B.n249 163.367
R498 B.n249 B.n68 163.367
R499 B.n245 B.n68 163.367
R500 B.n245 B.n244 163.367
R501 B.n244 B.n243 163.367
R502 B.n243 B.n70 163.367
R503 B.n239 B.n70 163.367
R504 B.n239 B.n238 163.367
R505 B.n238 B.n237 163.367
R506 B.n237 B.n72 163.367
R507 B.n233 B.n72 163.367
R508 B.n390 B.n15 163.367
R509 B.n390 B.n389 163.367
R510 B.n389 B.n388 163.367
R511 B.n388 B.n17 163.367
R512 B.n384 B.n17 163.367
R513 B.n384 B.n383 163.367
R514 B.n383 B.n382 163.367
R515 B.n382 B.n19 163.367
R516 B.n378 B.n19 163.367
R517 B.n378 B.n377 163.367
R518 B.n377 B.n376 163.367
R519 B.n376 B.n21 163.367
R520 B.n372 B.n21 163.367
R521 B.n372 B.n371 163.367
R522 B.n371 B.n370 163.367
R523 B.n370 B.n23 163.367
R524 B.n366 B.n23 163.367
R525 B.n366 B.n365 163.367
R526 B.n365 B.n364 163.367
R527 B.n364 B.n25 163.367
R528 B.n359 B.n25 163.367
R529 B.n359 B.n358 163.367
R530 B.n358 B.n357 163.367
R531 B.n357 B.n29 163.367
R532 B.n353 B.n29 163.367
R533 B.n353 B.n352 163.367
R534 B.n352 B.n351 163.367
R535 B.n351 B.n31 163.367
R536 B.n347 B.n31 163.367
R537 B.n347 B.n346 163.367
R538 B.n346 B.n345 163.367
R539 B.n345 B.n33 163.367
R540 B.n341 B.n33 163.367
R541 B.n341 B.n340 163.367
R542 B.n340 B.n339 163.367
R543 B.n339 B.n38 163.367
R544 B.n335 B.n38 163.367
R545 B.n335 B.n334 163.367
R546 B.n334 B.n333 163.367
R547 B.n333 B.n40 163.367
R548 B.n329 B.n40 163.367
R549 B.n329 B.n328 163.367
R550 B.n328 B.n327 163.367
R551 B.n327 B.n42 163.367
R552 B.n323 B.n42 163.367
R553 B.n323 B.n322 163.367
R554 B.n322 B.n321 163.367
R555 B.n321 B.n44 163.367
R556 B.n317 B.n44 163.367
R557 B.n317 B.n316 163.367
R558 B.n316 B.n315 163.367
R559 B.n395 B.n394 163.367
R560 B.n396 B.n395 163.367
R561 B.n396 B.n13 163.367
R562 B.n400 B.n13 163.367
R563 B.n401 B.n400 163.367
R564 B.n402 B.n401 163.367
R565 B.n402 B.n11 163.367
R566 B.n406 B.n11 163.367
R567 B.n407 B.n406 163.367
R568 B.n408 B.n407 163.367
R569 B.n408 B.n9 163.367
R570 B.n412 B.n9 163.367
R571 B.n413 B.n412 163.367
R572 B.n414 B.n413 163.367
R573 B.n414 B.n7 163.367
R574 B.n418 B.n7 163.367
R575 B.n419 B.n418 163.367
R576 B.n420 B.n419 163.367
R577 B.n420 B.n5 163.367
R578 B.n424 B.n5 163.367
R579 B.n425 B.n424 163.367
R580 B.n426 B.n425 163.367
R581 B.n426 B.n3 163.367
R582 B.n430 B.n3 163.367
R583 B.n431 B.n430 163.367
R584 B.n114 B.n2 163.367
R585 B.n115 B.n114 163.367
R586 B.n115 B.n112 163.367
R587 B.n119 B.n112 163.367
R588 B.n120 B.n119 163.367
R589 B.n121 B.n120 163.367
R590 B.n121 B.n110 163.367
R591 B.n125 B.n110 163.367
R592 B.n126 B.n125 163.367
R593 B.n127 B.n126 163.367
R594 B.n127 B.n108 163.367
R595 B.n131 B.n108 163.367
R596 B.n132 B.n131 163.367
R597 B.n133 B.n132 163.367
R598 B.n133 B.n106 163.367
R599 B.n137 B.n106 163.367
R600 B.n138 B.n137 163.367
R601 B.n139 B.n138 163.367
R602 B.n139 B.n104 163.367
R603 B.n143 B.n104 163.367
R604 B.n144 B.n143 163.367
R605 B.n145 B.n144 163.367
R606 B.n145 B.n102 163.367
R607 B.n149 B.n102 163.367
R608 B.n150 B.n149 163.367
R609 B.n197 B.t4 140.25
R610 B.n34 B.t2 140.25
R611 B.n89 B.t10 140.244
R612 B.n26 B.t8 140.244
R613 B.n198 B.t5 120.079
R614 B.n35 B.t1 120.079
R615 B.n90 B.t11 120.075
R616 B.n27 B.t7 120.075
R617 B.n183 B.n90 59.5399
R618 B.n199 B.n198 59.5399
R619 B.n36 B.n35 59.5399
R620 B.n361 B.n27 59.5399
R621 B.n393 B.n392 31.6883
R622 B.n314 B.n313 31.6883
R623 B.n234 B.n73 31.6883
R624 B.n152 B.n101 31.6883
R625 B.n90 B.n89 20.1702
R626 B.n198 B.n197 20.1702
R627 B.n35 B.n34 20.1702
R628 B.n27 B.n26 20.1702
R629 B B.n433 18.0485
R630 B.n393 B.n14 10.6151
R631 B.n397 B.n14 10.6151
R632 B.n398 B.n397 10.6151
R633 B.n399 B.n398 10.6151
R634 B.n399 B.n12 10.6151
R635 B.n403 B.n12 10.6151
R636 B.n404 B.n403 10.6151
R637 B.n405 B.n404 10.6151
R638 B.n405 B.n10 10.6151
R639 B.n409 B.n10 10.6151
R640 B.n410 B.n409 10.6151
R641 B.n411 B.n410 10.6151
R642 B.n411 B.n8 10.6151
R643 B.n415 B.n8 10.6151
R644 B.n416 B.n415 10.6151
R645 B.n417 B.n416 10.6151
R646 B.n417 B.n6 10.6151
R647 B.n421 B.n6 10.6151
R648 B.n422 B.n421 10.6151
R649 B.n423 B.n422 10.6151
R650 B.n423 B.n4 10.6151
R651 B.n427 B.n4 10.6151
R652 B.n428 B.n427 10.6151
R653 B.n429 B.n428 10.6151
R654 B.n429 B.n0 10.6151
R655 B.n392 B.n391 10.6151
R656 B.n391 B.n16 10.6151
R657 B.n387 B.n16 10.6151
R658 B.n387 B.n386 10.6151
R659 B.n386 B.n385 10.6151
R660 B.n385 B.n18 10.6151
R661 B.n381 B.n18 10.6151
R662 B.n381 B.n380 10.6151
R663 B.n380 B.n379 10.6151
R664 B.n379 B.n20 10.6151
R665 B.n375 B.n20 10.6151
R666 B.n375 B.n374 10.6151
R667 B.n374 B.n373 10.6151
R668 B.n373 B.n22 10.6151
R669 B.n369 B.n22 10.6151
R670 B.n369 B.n368 10.6151
R671 B.n368 B.n367 10.6151
R672 B.n367 B.n24 10.6151
R673 B.n363 B.n24 10.6151
R674 B.n363 B.n362 10.6151
R675 B.n360 B.n28 10.6151
R676 B.n356 B.n28 10.6151
R677 B.n356 B.n355 10.6151
R678 B.n355 B.n354 10.6151
R679 B.n354 B.n30 10.6151
R680 B.n350 B.n30 10.6151
R681 B.n350 B.n349 10.6151
R682 B.n349 B.n348 10.6151
R683 B.n348 B.n32 10.6151
R684 B.n344 B.n343 10.6151
R685 B.n343 B.n342 10.6151
R686 B.n342 B.n37 10.6151
R687 B.n338 B.n37 10.6151
R688 B.n338 B.n337 10.6151
R689 B.n337 B.n336 10.6151
R690 B.n336 B.n39 10.6151
R691 B.n332 B.n39 10.6151
R692 B.n332 B.n331 10.6151
R693 B.n331 B.n330 10.6151
R694 B.n330 B.n41 10.6151
R695 B.n326 B.n41 10.6151
R696 B.n326 B.n325 10.6151
R697 B.n325 B.n324 10.6151
R698 B.n324 B.n43 10.6151
R699 B.n320 B.n43 10.6151
R700 B.n320 B.n319 10.6151
R701 B.n319 B.n318 10.6151
R702 B.n318 B.n45 10.6151
R703 B.n314 B.n45 10.6151
R704 B.n313 B.n312 10.6151
R705 B.n312 B.n47 10.6151
R706 B.n308 B.n47 10.6151
R707 B.n308 B.n307 10.6151
R708 B.n307 B.n306 10.6151
R709 B.n306 B.n49 10.6151
R710 B.n302 B.n49 10.6151
R711 B.n302 B.n301 10.6151
R712 B.n301 B.n300 10.6151
R713 B.n300 B.n51 10.6151
R714 B.n296 B.n51 10.6151
R715 B.n296 B.n295 10.6151
R716 B.n295 B.n294 10.6151
R717 B.n294 B.n53 10.6151
R718 B.n290 B.n53 10.6151
R719 B.n290 B.n289 10.6151
R720 B.n289 B.n288 10.6151
R721 B.n288 B.n55 10.6151
R722 B.n284 B.n55 10.6151
R723 B.n284 B.n283 10.6151
R724 B.n283 B.n282 10.6151
R725 B.n282 B.n57 10.6151
R726 B.n278 B.n57 10.6151
R727 B.n278 B.n277 10.6151
R728 B.n277 B.n276 10.6151
R729 B.n276 B.n59 10.6151
R730 B.n272 B.n59 10.6151
R731 B.n272 B.n271 10.6151
R732 B.n271 B.n270 10.6151
R733 B.n270 B.n61 10.6151
R734 B.n266 B.n61 10.6151
R735 B.n266 B.n265 10.6151
R736 B.n265 B.n264 10.6151
R737 B.n264 B.n63 10.6151
R738 B.n260 B.n63 10.6151
R739 B.n260 B.n259 10.6151
R740 B.n259 B.n258 10.6151
R741 B.n258 B.n65 10.6151
R742 B.n254 B.n65 10.6151
R743 B.n254 B.n253 10.6151
R744 B.n253 B.n252 10.6151
R745 B.n252 B.n67 10.6151
R746 B.n248 B.n67 10.6151
R747 B.n248 B.n247 10.6151
R748 B.n247 B.n246 10.6151
R749 B.n246 B.n69 10.6151
R750 B.n242 B.n69 10.6151
R751 B.n242 B.n241 10.6151
R752 B.n241 B.n240 10.6151
R753 B.n240 B.n71 10.6151
R754 B.n236 B.n71 10.6151
R755 B.n236 B.n235 10.6151
R756 B.n235 B.n234 10.6151
R757 B.n113 B.n1 10.6151
R758 B.n116 B.n113 10.6151
R759 B.n117 B.n116 10.6151
R760 B.n118 B.n117 10.6151
R761 B.n118 B.n111 10.6151
R762 B.n122 B.n111 10.6151
R763 B.n123 B.n122 10.6151
R764 B.n124 B.n123 10.6151
R765 B.n124 B.n109 10.6151
R766 B.n128 B.n109 10.6151
R767 B.n129 B.n128 10.6151
R768 B.n130 B.n129 10.6151
R769 B.n130 B.n107 10.6151
R770 B.n134 B.n107 10.6151
R771 B.n135 B.n134 10.6151
R772 B.n136 B.n135 10.6151
R773 B.n136 B.n105 10.6151
R774 B.n140 B.n105 10.6151
R775 B.n141 B.n140 10.6151
R776 B.n142 B.n141 10.6151
R777 B.n142 B.n103 10.6151
R778 B.n146 B.n103 10.6151
R779 B.n147 B.n146 10.6151
R780 B.n148 B.n147 10.6151
R781 B.n148 B.n101 10.6151
R782 B.n153 B.n152 10.6151
R783 B.n154 B.n153 10.6151
R784 B.n154 B.n99 10.6151
R785 B.n158 B.n99 10.6151
R786 B.n159 B.n158 10.6151
R787 B.n160 B.n159 10.6151
R788 B.n160 B.n97 10.6151
R789 B.n164 B.n97 10.6151
R790 B.n165 B.n164 10.6151
R791 B.n166 B.n165 10.6151
R792 B.n166 B.n95 10.6151
R793 B.n170 B.n95 10.6151
R794 B.n171 B.n170 10.6151
R795 B.n172 B.n171 10.6151
R796 B.n172 B.n93 10.6151
R797 B.n176 B.n93 10.6151
R798 B.n177 B.n176 10.6151
R799 B.n178 B.n177 10.6151
R800 B.n178 B.n91 10.6151
R801 B.n182 B.n91 10.6151
R802 B.n185 B.n184 10.6151
R803 B.n185 B.n87 10.6151
R804 B.n189 B.n87 10.6151
R805 B.n190 B.n189 10.6151
R806 B.n191 B.n190 10.6151
R807 B.n191 B.n85 10.6151
R808 B.n195 B.n85 10.6151
R809 B.n196 B.n195 10.6151
R810 B.n200 B.n196 10.6151
R811 B.n204 B.n83 10.6151
R812 B.n205 B.n204 10.6151
R813 B.n206 B.n205 10.6151
R814 B.n206 B.n81 10.6151
R815 B.n210 B.n81 10.6151
R816 B.n211 B.n210 10.6151
R817 B.n212 B.n211 10.6151
R818 B.n212 B.n79 10.6151
R819 B.n216 B.n79 10.6151
R820 B.n217 B.n216 10.6151
R821 B.n218 B.n217 10.6151
R822 B.n218 B.n77 10.6151
R823 B.n222 B.n77 10.6151
R824 B.n223 B.n222 10.6151
R825 B.n224 B.n223 10.6151
R826 B.n224 B.n75 10.6151
R827 B.n228 B.n75 10.6151
R828 B.n229 B.n228 10.6151
R829 B.n230 B.n229 10.6151
R830 B.n230 B.n73 10.6151
R831 B.n362 B.n361 9.36635
R832 B.n344 B.n36 9.36635
R833 B.n183 B.n182 9.36635
R834 B.n199 B.n83 9.36635
R835 B.n433 B.n0 8.11757
R836 B.n433 B.n1 8.11757
R837 B.n361 B.n360 1.24928
R838 B.n36 B.n32 1.24928
R839 B.n184 B.n183 1.24928
R840 B.n200 B.n199 1.24928
C0 VDD2 VTAIL 7.44919f
C1 VDD2 VP 0.345558f
C2 VN w_n2218_n1978# 4.04356f
C3 VN B 0.727443f
C4 B w_n2218_n1978# 5.42344f
C5 VN VDD2 3.09531f
C6 VDD2 w_n2218_n1978# 1.57179f
C7 VDD2 B 1.24634f
C8 VDD1 VTAIL 7.411049f
C9 VDD1 VP 3.28572f
C10 VP VTAIL 3.29958f
C11 VN VDD1 0.148708f
C12 VDD1 w_n2218_n1978# 1.52694f
C13 VDD1 B 1.20163f
C14 VN VTAIL 3.28526f
C15 VN VP 4.32495f
C16 VTAIL w_n2218_n1978# 1.91669f
C17 VTAIL B 1.48916f
C18 VP w_n2218_n1978# 4.32641f
C19 VP B 1.19274f
C20 VDD1 VDD2 0.974489f
C21 VDD2 VSUBS 1.090333f
C22 VDD1 VSUBS 0.937658f
C23 VTAIL VSUBS 0.4099f
C24 VN VSUBS 4.42458f
C25 VP VSUBS 1.470065f
C26 B VSUBS 2.330262f
C27 w_n2218_n1978# VSUBS 54.961998f
C28 B.n0 VSUBS 0.006017f
C29 B.n1 VSUBS 0.006017f
C30 B.n2 VSUBS 0.008899f
C31 B.n3 VSUBS 0.006819f
C32 B.n4 VSUBS 0.006819f
C33 B.n5 VSUBS 0.006819f
C34 B.n6 VSUBS 0.006819f
C35 B.n7 VSUBS 0.006819f
C36 B.n8 VSUBS 0.006819f
C37 B.n9 VSUBS 0.006819f
C38 B.n10 VSUBS 0.006819f
C39 B.n11 VSUBS 0.006819f
C40 B.n12 VSUBS 0.006819f
C41 B.n13 VSUBS 0.006819f
C42 B.n14 VSUBS 0.006819f
C43 B.n15 VSUBS 0.01604f
C44 B.n16 VSUBS 0.006819f
C45 B.n17 VSUBS 0.006819f
C46 B.n18 VSUBS 0.006819f
C47 B.n19 VSUBS 0.006819f
C48 B.n20 VSUBS 0.006819f
C49 B.n21 VSUBS 0.006819f
C50 B.n22 VSUBS 0.006819f
C51 B.n23 VSUBS 0.006819f
C52 B.n24 VSUBS 0.006819f
C53 B.n25 VSUBS 0.006819f
C54 B.t7 VSUBS 0.13755f
C55 B.t8 VSUBS 0.144916f
C56 B.t6 VSUBS 0.153394f
C57 B.n26 VSUBS 0.079584f
C58 B.n27 VSUBS 0.060946f
C59 B.n28 VSUBS 0.006819f
C60 B.n29 VSUBS 0.006819f
C61 B.n30 VSUBS 0.006819f
C62 B.n31 VSUBS 0.006819f
C63 B.n32 VSUBS 0.003811f
C64 B.n33 VSUBS 0.006819f
C65 B.t1 VSUBS 0.13755f
C66 B.t2 VSUBS 0.144916f
C67 B.t0 VSUBS 0.153394f
C68 B.n34 VSUBS 0.079585f
C69 B.n35 VSUBS 0.060946f
C70 B.n36 VSUBS 0.0158f
C71 B.n37 VSUBS 0.006819f
C72 B.n38 VSUBS 0.006819f
C73 B.n39 VSUBS 0.006819f
C74 B.n40 VSUBS 0.006819f
C75 B.n41 VSUBS 0.006819f
C76 B.n42 VSUBS 0.006819f
C77 B.n43 VSUBS 0.006819f
C78 B.n44 VSUBS 0.006819f
C79 B.n45 VSUBS 0.006819f
C80 B.n46 VSUBS 0.01525f
C81 B.n47 VSUBS 0.006819f
C82 B.n48 VSUBS 0.006819f
C83 B.n49 VSUBS 0.006819f
C84 B.n50 VSUBS 0.006819f
C85 B.n51 VSUBS 0.006819f
C86 B.n52 VSUBS 0.006819f
C87 B.n53 VSUBS 0.006819f
C88 B.n54 VSUBS 0.006819f
C89 B.n55 VSUBS 0.006819f
C90 B.n56 VSUBS 0.006819f
C91 B.n57 VSUBS 0.006819f
C92 B.n58 VSUBS 0.006819f
C93 B.n59 VSUBS 0.006819f
C94 B.n60 VSUBS 0.006819f
C95 B.n61 VSUBS 0.006819f
C96 B.n62 VSUBS 0.006819f
C97 B.n63 VSUBS 0.006819f
C98 B.n64 VSUBS 0.006819f
C99 B.n65 VSUBS 0.006819f
C100 B.n66 VSUBS 0.006819f
C101 B.n67 VSUBS 0.006819f
C102 B.n68 VSUBS 0.006819f
C103 B.n69 VSUBS 0.006819f
C104 B.n70 VSUBS 0.006819f
C105 B.n71 VSUBS 0.006819f
C106 B.n72 VSUBS 0.006819f
C107 B.n73 VSUBS 0.015209f
C108 B.n74 VSUBS 0.006819f
C109 B.n75 VSUBS 0.006819f
C110 B.n76 VSUBS 0.006819f
C111 B.n77 VSUBS 0.006819f
C112 B.n78 VSUBS 0.006819f
C113 B.n79 VSUBS 0.006819f
C114 B.n80 VSUBS 0.006819f
C115 B.n81 VSUBS 0.006819f
C116 B.n82 VSUBS 0.006819f
C117 B.n83 VSUBS 0.006418f
C118 B.n84 VSUBS 0.006819f
C119 B.n85 VSUBS 0.006819f
C120 B.n86 VSUBS 0.006819f
C121 B.n87 VSUBS 0.006819f
C122 B.n88 VSUBS 0.006819f
C123 B.t11 VSUBS 0.13755f
C124 B.t10 VSUBS 0.144916f
C125 B.t9 VSUBS 0.153394f
C126 B.n89 VSUBS 0.079584f
C127 B.n90 VSUBS 0.060946f
C128 B.n91 VSUBS 0.006819f
C129 B.n92 VSUBS 0.006819f
C130 B.n93 VSUBS 0.006819f
C131 B.n94 VSUBS 0.006819f
C132 B.n95 VSUBS 0.006819f
C133 B.n96 VSUBS 0.006819f
C134 B.n97 VSUBS 0.006819f
C135 B.n98 VSUBS 0.006819f
C136 B.n99 VSUBS 0.006819f
C137 B.n100 VSUBS 0.006819f
C138 B.n101 VSUBS 0.01525f
C139 B.n102 VSUBS 0.006819f
C140 B.n103 VSUBS 0.006819f
C141 B.n104 VSUBS 0.006819f
C142 B.n105 VSUBS 0.006819f
C143 B.n106 VSUBS 0.006819f
C144 B.n107 VSUBS 0.006819f
C145 B.n108 VSUBS 0.006819f
C146 B.n109 VSUBS 0.006819f
C147 B.n110 VSUBS 0.006819f
C148 B.n111 VSUBS 0.006819f
C149 B.n112 VSUBS 0.006819f
C150 B.n113 VSUBS 0.006819f
C151 B.n114 VSUBS 0.006819f
C152 B.n115 VSUBS 0.006819f
C153 B.n116 VSUBS 0.006819f
C154 B.n117 VSUBS 0.006819f
C155 B.n118 VSUBS 0.006819f
C156 B.n119 VSUBS 0.006819f
C157 B.n120 VSUBS 0.006819f
C158 B.n121 VSUBS 0.006819f
C159 B.n122 VSUBS 0.006819f
C160 B.n123 VSUBS 0.006819f
C161 B.n124 VSUBS 0.006819f
C162 B.n125 VSUBS 0.006819f
C163 B.n126 VSUBS 0.006819f
C164 B.n127 VSUBS 0.006819f
C165 B.n128 VSUBS 0.006819f
C166 B.n129 VSUBS 0.006819f
C167 B.n130 VSUBS 0.006819f
C168 B.n131 VSUBS 0.006819f
C169 B.n132 VSUBS 0.006819f
C170 B.n133 VSUBS 0.006819f
C171 B.n134 VSUBS 0.006819f
C172 B.n135 VSUBS 0.006819f
C173 B.n136 VSUBS 0.006819f
C174 B.n137 VSUBS 0.006819f
C175 B.n138 VSUBS 0.006819f
C176 B.n139 VSUBS 0.006819f
C177 B.n140 VSUBS 0.006819f
C178 B.n141 VSUBS 0.006819f
C179 B.n142 VSUBS 0.006819f
C180 B.n143 VSUBS 0.006819f
C181 B.n144 VSUBS 0.006819f
C182 B.n145 VSUBS 0.006819f
C183 B.n146 VSUBS 0.006819f
C184 B.n147 VSUBS 0.006819f
C185 B.n148 VSUBS 0.006819f
C186 B.n149 VSUBS 0.006819f
C187 B.n150 VSUBS 0.01525f
C188 B.n151 VSUBS 0.01604f
C189 B.n152 VSUBS 0.01604f
C190 B.n153 VSUBS 0.006819f
C191 B.n154 VSUBS 0.006819f
C192 B.n155 VSUBS 0.006819f
C193 B.n156 VSUBS 0.006819f
C194 B.n157 VSUBS 0.006819f
C195 B.n158 VSUBS 0.006819f
C196 B.n159 VSUBS 0.006819f
C197 B.n160 VSUBS 0.006819f
C198 B.n161 VSUBS 0.006819f
C199 B.n162 VSUBS 0.006819f
C200 B.n163 VSUBS 0.006819f
C201 B.n164 VSUBS 0.006819f
C202 B.n165 VSUBS 0.006819f
C203 B.n166 VSUBS 0.006819f
C204 B.n167 VSUBS 0.006819f
C205 B.n168 VSUBS 0.006819f
C206 B.n169 VSUBS 0.006819f
C207 B.n170 VSUBS 0.006819f
C208 B.n171 VSUBS 0.006819f
C209 B.n172 VSUBS 0.006819f
C210 B.n173 VSUBS 0.006819f
C211 B.n174 VSUBS 0.006819f
C212 B.n175 VSUBS 0.006819f
C213 B.n176 VSUBS 0.006819f
C214 B.n177 VSUBS 0.006819f
C215 B.n178 VSUBS 0.006819f
C216 B.n179 VSUBS 0.006819f
C217 B.n180 VSUBS 0.006819f
C218 B.n181 VSUBS 0.006819f
C219 B.n182 VSUBS 0.006418f
C220 B.n183 VSUBS 0.0158f
C221 B.n184 VSUBS 0.003811f
C222 B.n185 VSUBS 0.006819f
C223 B.n186 VSUBS 0.006819f
C224 B.n187 VSUBS 0.006819f
C225 B.n188 VSUBS 0.006819f
C226 B.n189 VSUBS 0.006819f
C227 B.n190 VSUBS 0.006819f
C228 B.n191 VSUBS 0.006819f
C229 B.n192 VSUBS 0.006819f
C230 B.n193 VSUBS 0.006819f
C231 B.n194 VSUBS 0.006819f
C232 B.n195 VSUBS 0.006819f
C233 B.n196 VSUBS 0.006819f
C234 B.t5 VSUBS 0.13755f
C235 B.t4 VSUBS 0.144916f
C236 B.t3 VSUBS 0.153394f
C237 B.n197 VSUBS 0.079585f
C238 B.n198 VSUBS 0.060946f
C239 B.n199 VSUBS 0.0158f
C240 B.n200 VSUBS 0.003811f
C241 B.n201 VSUBS 0.006819f
C242 B.n202 VSUBS 0.006819f
C243 B.n203 VSUBS 0.006819f
C244 B.n204 VSUBS 0.006819f
C245 B.n205 VSUBS 0.006819f
C246 B.n206 VSUBS 0.006819f
C247 B.n207 VSUBS 0.006819f
C248 B.n208 VSUBS 0.006819f
C249 B.n209 VSUBS 0.006819f
C250 B.n210 VSUBS 0.006819f
C251 B.n211 VSUBS 0.006819f
C252 B.n212 VSUBS 0.006819f
C253 B.n213 VSUBS 0.006819f
C254 B.n214 VSUBS 0.006819f
C255 B.n215 VSUBS 0.006819f
C256 B.n216 VSUBS 0.006819f
C257 B.n217 VSUBS 0.006819f
C258 B.n218 VSUBS 0.006819f
C259 B.n219 VSUBS 0.006819f
C260 B.n220 VSUBS 0.006819f
C261 B.n221 VSUBS 0.006819f
C262 B.n222 VSUBS 0.006819f
C263 B.n223 VSUBS 0.006819f
C264 B.n224 VSUBS 0.006819f
C265 B.n225 VSUBS 0.006819f
C266 B.n226 VSUBS 0.006819f
C267 B.n227 VSUBS 0.006819f
C268 B.n228 VSUBS 0.006819f
C269 B.n229 VSUBS 0.006819f
C270 B.n230 VSUBS 0.006819f
C271 B.n231 VSUBS 0.006819f
C272 B.n232 VSUBS 0.01604f
C273 B.n233 VSUBS 0.01525f
C274 B.n234 VSUBS 0.01608f
C275 B.n235 VSUBS 0.006819f
C276 B.n236 VSUBS 0.006819f
C277 B.n237 VSUBS 0.006819f
C278 B.n238 VSUBS 0.006819f
C279 B.n239 VSUBS 0.006819f
C280 B.n240 VSUBS 0.006819f
C281 B.n241 VSUBS 0.006819f
C282 B.n242 VSUBS 0.006819f
C283 B.n243 VSUBS 0.006819f
C284 B.n244 VSUBS 0.006819f
C285 B.n245 VSUBS 0.006819f
C286 B.n246 VSUBS 0.006819f
C287 B.n247 VSUBS 0.006819f
C288 B.n248 VSUBS 0.006819f
C289 B.n249 VSUBS 0.006819f
C290 B.n250 VSUBS 0.006819f
C291 B.n251 VSUBS 0.006819f
C292 B.n252 VSUBS 0.006819f
C293 B.n253 VSUBS 0.006819f
C294 B.n254 VSUBS 0.006819f
C295 B.n255 VSUBS 0.006819f
C296 B.n256 VSUBS 0.006819f
C297 B.n257 VSUBS 0.006819f
C298 B.n258 VSUBS 0.006819f
C299 B.n259 VSUBS 0.006819f
C300 B.n260 VSUBS 0.006819f
C301 B.n261 VSUBS 0.006819f
C302 B.n262 VSUBS 0.006819f
C303 B.n263 VSUBS 0.006819f
C304 B.n264 VSUBS 0.006819f
C305 B.n265 VSUBS 0.006819f
C306 B.n266 VSUBS 0.006819f
C307 B.n267 VSUBS 0.006819f
C308 B.n268 VSUBS 0.006819f
C309 B.n269 VSUBS 0.006819f
C310 B.n270 VSUBS 0.006819f
C311 B.n271 VSUBS 0.006819f
C312 B.n272 VSUBS 0.006819f
C313 B.n273 VSUBS 0.006819f
C314 B.n274 VSUBS 0.006819f
C315 B.n275 VSUBS 0.006819f
C316 B.n276 VSUBS 0.006819f
C317 B.n277 VSUBS 0.006819f
C318 B.n278 VSUBS 0.006819f
C319 B.n279 VSUBS 0.006819f
C320 B.n280 VSUBS 0.006819f
C321 B.n281 VSUBS 0.006819f
C322 B.n282 VSUBS 0.006819f
C323 B.n283 VSUBS 0.006819f
C324 B.n284 VSUBS 0.006819f
C325 B.n285 VSUBS 0.006819f
C326 B.n286 VSUBS 0.006819f
C327 B.n287 VSUBS 0.006819f
C328 B.n288 VSUBS 0.006819f
C329 B.n289 VSUBS 0.006819f
C330 B.n290 VSUBS 0.006819f
C331 B.n291 VSUBS 0.006819f
C332 B.n292 VSUBS 0.006819f
C333 B.n293 VSUBS 0.006819f
C334 B.n294 VSUBS 0.006819f
C335 B.n295 VSUBS 0.006819f
C336 B.n296 VSUBS 0.006819f
C337 B.n297 VSUBS 0.006819f
C338 B.n298 VSUBS 0.006819f
C339 B.n299 VSUBS 0.006819f
C340 B.n300 VSUBS 0.006819f
C341 B.n301 VSUBS 0.006819f
C342 B.n302 VSUBS 0.006819f
C343 B.n303 VSUBS 0.006819f
C344 B.n304 VSUBS 0.006819f
C345 B.n305 VSUBS 0.006819f
C346 B.n306 VSUBS 0.006819f
C347 B.n307 VSUBS 0.006819f
C348 B.n308 VSUBS 0.006819f
C349 B.n309 VSUBS 0.006819f
C350 B.n310 VSUBS 0.006819f
C351 B.n311 VSUBS 0.006819f
C352 B.n312 VSUBS 0.006819f
C353 B.n313 VSUBS 0.01525f
C354 B.n314 VSUBS 0.01604f
C355 B.n315 VSUBS 0.01604f
C356 B.n316 VSUBS 0.006819f
C357 B.n317 VSUBS 0.006819f
C358 B.n318 VSUBS 0.006819f
C359 B.n319 VSUBS 0.006819f
C360 B.n320 VSUBS 0.006819f
C361 B.n321 VSUBS 0.006819f
C362 B.n322 VSUBS 0.006819f
C363 B.n323 VSUBS 0.006819f
C364 B.n324 VSUBS 0.006819f
C365 B.n325 VSUBS 0.006819f
C366 B.n326 VSUBS 0.006819f
C367 B.n327 VSUBS 0.006819f
C368 B.n328 VSUBS 0.006819f
C369 B.n329 VSUBS 0.006819f
C370 B.n330 VSUBS 0.006819f
C371 B.n331 VSUBS 0.006819f
C372 B.n332 VSUBS 0.006819f
C373 B.n333 VSUBS 0.006819f
C374 B.n334 VSUBS 0.006819f
C375 B.n335 VSUBS 0.006819f
C376 B.n336 VSUBS 0.006819f
C377 B.n337 VSUBS 0.006819f
C378 B.n338 VSUBS 0.006819f
C379 B.n339 VSUBS 0.006819f
C380 B.n340 VSUBS 0.006819f
C381 B.n341 VSUBS 0.006819f
C382 B.n342 VSUBS 0.006819f
C383 B.n343 VSUBS 0.006819f
C384 B.n344 VSUBS 0.006418f
C385 B.n345 VSUBS 0.006819f
C386 B.n346 VSUBS 0.006819f
C387 B.n347 VSUBS 0.006819f
C388 B.n348 VSUBS 0.006819f
C389 B.n349 VSUBS 0.006819f
C390 B.n350 VSUBS 0.006819f
C391 B.n351 VSUBS 0.006819f
C392 B.n352 VSUBS 0.006819f
C393 B.n353 VSUBS 0.006819f
C394 B.n354 VSUBS 0.006819f
C395 B.n355 VSUBS 0.006819f
C396 B.n356 VSUBS 0.006819f
C397 B.n357 VSUBS 0.006819f
C398 B.n358 VSUBS 0.006819f
C399 B.n359 VSUBS 0.006819f
C400 B.n360 VSUBS 0.003811f
C401 B.n361 VSUBS 0.0158f
C402 B.n362 VSUBS 0.006418f
C403 B.n363 VSUBS 0.006819f
C404 B.n364 VSUBS 0.006819f
C405 B.n365 VSUBS 0.006819f
C406 B.n366 VSUBS 0.006819f
C407 B.n367 VSUBS 0.006819f
C408 B.n368 VSUBS 0.006819f
C409 B.n369 VSUBS 0.006819f
C410 B.n370 VSUBS 0.006819f
C411 B.n371 VSUBS 0.006819f
C412 B.n372 VSUBS 0.006819f
C413 B.n373 VSUBS 0.006819f
C414 B.n374 VSUBS 0.006819f
C415 B.n375 VSUBS 0.006819f
C416 B.n376 VSUBS 0.006819f
C417 B.n377 VSUBS 0.006819f
C418 B.n378 VSUBS 0.006819f
C419 B.n379 VSUBS 0.006819f
C420 B.n380 VSUBS 0.006819f
C421 B.n381 VSUBS 0.006819f
C422 B.n382 VSUBS 0.006819f
C423 B.n383 VSUBS 0.006819f
C424 B.n384 VSUBS 0.006819f
C425 B.n385 VSUBS 0.006819f
C426 B.n386 VSUBS 0.006819f
C427 B.n387 VSUBS 0.006819f
C428 B.n388 VSUBS 0.006819f
C429 B.n389 VSUBS 0.006819f
C430 B.n390 VSUBS 0.006819f
C431 B.n391 VSUBS 0.006819f
C432 B.n392 VSUBS 0.01604f
C433 B.n393 VSUBS 0.01525f
C434 B.n394 VSUBS 0.01525f
C435 B.n395 VSUBS 0.006819f
C436 B.n396 VSUBS 0.006819f
C437 B.n397 VSUBS 0.006819f
C438 B.n398 VSUBS 0.006819f
C439 B.n399 VSUBS 0.006819f
C440 B.n400 VSUBS 0.006819f
C441 B.n401 VSUBS 0.006819f
C442 B.n402 VSUBS 0.006819f
C443 B.n403 VSUBS 0.006819f
C444 B.n404 VSUBS 0.006819f
C445 B.n405 VSUBS 0.006819f
C446 B.n406 VSUBS 0.006819f
C447 B.n407 VSUBS 0.006819f
C448 B.n408 VSUBS 0.006819f
C449 B.n409 VSUBS 0.006819f
C450 B.n410 VSUBS 0.006819f
C451 B.n411 VSUBS 0.006819f
C452 B.n412 VSUBS 0.006819f
C453 B.n413 VSUBS 0.006819f
C454 B.n414 VSUBS 0.006819f
C455 B.n415 VSUBS 0.006819f
C456 B.n416 VSUBS 0.006819f
C457 B.n417 VSUBS 0.006819f
C458 B.n418 VSUBS 0.006819f
C459 B.n419 VSUBS 0.006819f
C460 B.n420 VSUBS 0.006819f
C461 B.n421 VSUBS 0.006819f
C462 B.n422 VSUBS 0.006819f
C463 B.n423 VSUBS 0.006819f
C464 B.n424 VSUBS 0.006819f
C465 B.n425 VSUBS 0.006819f
C466 B.n426 VSUBS 0.006819f
C467 B.n427 VSUBS 0.006819f
C468 B.n428 VSUBS 0.006819f
C469 B.n429 VSUBS 0.006819f
C470 B.n430 VSUBS 0.006819f
C471 B.n431 VSUBS 0.008899f
C472 B.n432 VSUBS 0.00948f
C473 B.n433 VSUBS 0.018851f
C474 VDD2.t9 VSUBS 0.839166f
C475 VDD2.t6 VSUBS 0.097433f
C476 VDD2.t2 VSUBS 0.097433f
C477 VDD2.n0 VSUBS 0.61549f
C478 VDD2.n1 VSUBS 0.957037f
C479 VDD2.t7 VSUBS 0.097433f
C480 VDD2.t4 VSUBS 0.097433f
C481 VDD2.n2 VSUBS 0.61849f
C482 VDD2.n3 VSUBS 1.63472f
C483 VDD2.t1 VSUBS 0.835104f
C484 VDD2.n4 VSUBS 1.95013f
C485 VDD2.t0 VSUBS 0.097433f
C486 VDD2.t8 VSUBS 0.097433f
C487 VDD2.n5 VSUBS 0.615492f
C488 VDD2.n6 VSUBS 0.466469f
C489 VDD2.t5 VSUBS 0.097433f
C490 VDD2.t3 VSUBS 0.097433f
C491 VDD2.n7 VSUBS 0.618468f
C492 VN.n0 VSUBS 0.060228f
C493 VN.n1 VSUBS 0.013667f
C494 VN.n2 VSUBS 0.253399f
C495 VN.t0 VSUBS 0.659234f
C496 VN.n3 VSUBS 0.283066f
C497 VN.t3 VSUBS 0.630748f
C498 VN.n4 VSUBS 0.312521f
C499 VN.n5 VSUBS 0.013667f
C500 VN.t7 VSUBS 0.630748f
C501 VN.n6 VSUBS 0.305785f
C502 VN.n7 VSUBS 0.060228f
C503 VN.n8 VSUBS 0.060228f
C504 VN.n9 VSUBS 0.060228f
C505 VN.t2 VSUBS 0.630748f
C506 VN.n10 VSUBS 0.305785f
C507 VN.n11 VSUBS 0.013667f
C508 VN.t5 VSUBS 0.630748f
C509 VN.n12 VSUBS 0.303371f
C510 VN.n13 VSUBS 0.046674f
C511 VN.n14 VSUBS 0.060228f
C512 VN.n15 VSUBS 0.013667f
C513 VN.t9 VSUBS 0.630748f
C514 VN.n16 VSUBS 0.253399f
C515 VN.t6 VSUBS 0.659234f
C516 VN.n17 VSUBS 0.283066f
C517 VN.t4 VSUBS 0.630748f
C518 VN.n18 VSUBS 0.312521f
C519 VN.n19 VSUBS 0.013667f
C520 VN.t1 VSUBS 0.630748f
C521 VN.n20 VSUBS 0.305785f
C522 VN.n21 VSUBS 0.060228f
C523 VN.n22 VSUBS 0.060228f
C524 VN.n23 VSUBS 0.060228f
C525 VN.n24 VSUBS 0.305785f
C526 VN.n25 VSUBS 0.013667f
C527 VN.t8 VSUBS 0.630748f
C528 VN.n26 VSUBS 0.303371f
C529 VN.n27 VSUBS 2.09063f
C530 VTAIL.t1 VSUBS 0.111911f
C531 VTAIL.t3 VSUBS 0.111911f
C532 VTAIL.n0 VSUBS 0.625003f
C533 VTAIL.n1 VSUBS 0.622072f
C534 VTAIL.t14 VSUBS 0.873408f
C535 VTAIL.n2 VSUBS 0.693875f
C536 VTAIL.t10 VSUBS 0.111911f
C537 VTAIL.t13 VSUBS 0.111911f
C538 VTAIL.n3 VSUBS 0.625003f
C539 VTAIL.n4 VSUBS 0.635119f
C540 VTAIL.t16 VSUBS 0.111911f
C541 VTAIL.t17 VSUBS 0.111911f
C542 VTAIL.n5 VSUBS 0.625003f
C543 VTAIL.n6 VSUBS 1.49045f
C544 VTAIL.t9 VSUBS 0.111911f
C545 VTAIL.t2 VSUBS 0.111911f
C546 VTAIL.n7 VSUBS 0.625006f
C547 VTAIL.n8 VSUBS 1.49045f
C548 VTAIL.t5 VSUBS 0.111911f
C549 VTAIL.t4 VSUBS 0.111911f
C550 VTAIL.n9 VSUBS 0.625006f
C551 VTAIL.n10 VSUBS 0.635116f
C552 VTAIL.t0 VSUBS 0.873412f
C553 VTAIL.n11 VSUBS 0.69387f
C554 VTAIL.t15 VSUBS 0.111911f
C555 VTAIL.t18 VSUBS 0.111911f
C556 VTAIL.n12 VSUBS 0.625006f
C557 VTAIL.n13 VSUBS 0.637063f
C558 VTAIL.t11 VSUBS 0.111911f
C559 VTAIL.t19 VSUBS 0.111911f
C560 VTAIL.n14 VSUBS 0.625006f
C561 VTAIL.n15 VSUBS 0.635116f
C562 VTAIL.t12 VSUBS 0.873408f
C563 VTAIL.n16 VSUBS 1.46625f
C564 VTAIL.t7 VSUBS 0.873408f
C565 VTAIL.n17 VSUBS 1.46625f
C566 VTAIL.t8 VSUBS 0.111911f
C567 VTAIL.t6 VSUBS 0.111911f
C568 VTAIL.n18 VSUBS 0.625003f
C569 VTAIL.n19 VSUBS 0.569101f
C570 VDD1.t0 VSUBS 0.847872f
C571 VDD1.t5 VSUBS 0.098444f
C572 VDD1.t8 VSUBS 0.098444f
C573 VDD1.n0 VSUBS 0.621875f
C574 VDD1.n1 VSUBS 0.972592f
C575 VDD1.t1 VSUBS 0.847869f
C576 VDD1.t3 VSUBS 0.098444f
C577 VDD1.t7 VSUBS 0.098444f
C578 VDD1.n2 VSUBS 0.621872f
C579 VDD1.n3 VSUBS 0.966961f
C580 VDD1.t4 VSUBS 0.098444f
C581 VDD1.t6 VSUBS 0.098444f
C582 VDD1.n4 VSUBS 0.624903f
C583 VDD1.n5 VSUBS 1.72496f
C584 VDD1.t2 VSUBS 0.098444f
C585 VDD1.t9 VSUBS 0.098444f
C586 VDD1.n6 VSUBS 0.621872f
C587 VDD1.n7 VSUBS 1.99041f
C588 VP.n0 VSUBS 0.062637f
C589 VP.n1 VSUBS 0.014214f
C590 VP.n2 VSUBS 0.062637f
C591 VP.n3 VSUBS 0.014214f
C592 VP.n4 VSUBS 0.062637f
C593 VP.t7 VSUBS 0.65598f
C594 VP.t0 VSUBS 0.65598f
C595 VP.n5 VSUBS 0.062637f
C596 VP.t8 VSUBS 0.65598f
C597 VP.n6 VSUBS 0.318017f
C598 VP.t4 VSUBS 0.685606f
C599 VP.n7 VSUBS 0.29439f
C600 VP.t1 VSUBS 0.65598f
C601 VP.n8 VSUBS 0.325023f
C602 VP.n9 VSUBS 0.014214f
C603 VP.n10 VSUBS 0.263535f
C604 VP.n11 VSUBS 0.062637f
C605 VP.n12 VSUBS 0.062637f
C606 VP.n13 VSUBS 0.014214f
C607 VP.n14 VSUBS 0.318017f
C608 VP.n15 VSUBS 0.014214f
C609 VP.n16 VSUBS 0.315507f
C610 VP.n17 VSUBS 2.13285f
C611 VP.t3 VSUBS 0.65598f
C612 VP.n18 VSUBS 0.315507f
C613 VP.n19 VSUBS 2.19275f
C614 VP.n20 VSUBS 0.062637f
C615 VP.n21 VSUBS 0.062637f
C616 VP.t2 VSUBS 0.65598f
C617 VP.n22 VSUBS 0.318017f
C618 VP.n23 VSUBS 0.014214f
C619 VP.t9 VSUBS 0.65598f
C620 VP.n24 VSUBS 0.318017f
C621 VP.n25 VSUBS 0.062637f
C622 VP.n26 VSUBS 0.062637f
C623 VP.n27 VSUBS 0.062637f
C624 VP.t6 VSUBS 0.65598f
C625 VP.n28 VSUBS 0.318017f
C626 VP.n29 VSUBS 0.014214f
C627 VP.t5 VSUBS 0.65598f
C628 VP.n30 VSUBS 0.315507f
C629 VP.n31 VSUBS 0.048541f
.ends

