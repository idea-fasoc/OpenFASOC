* NGSPICE file created from diff_pair_sample_0374.ext - technology: sky130A

.subckt diff_pair_sample_0374 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=0 ps=0 w=9.2 l=3.07
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=3.588 ps=19.18 w=9.2 l=3.07
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=3.588 ps=19.18 w=9.2 l=3.07
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=0 ps=0 w=9.2 l=3.07
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=3.588 ps=19.18 w=9.2 l=3.07
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=3.588 ps=19.18 w=9.2 l=3.07
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=0 ps=0 w=9.2 l=3.07
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.588 pd=19.18 as=0 ps=0 w=9.2 l=3.07
R0 B.n616 B.n615 585
R1 B.n245 B.n92 585
R2 B.n244 B.n243 585
R3 B.n242 B.n241 585
R4 B.n240 B.n239 585
R5 B.n238 B.n237 585
R6 B.n236 B.n235 585
R7 B.n234 B.n233 585
R8 B.n232 B.n231 585
R9 B.n230 B.n229 585
R10 B.n228 B.n227 585
R11 B.n226 B.n225 585
R12 B.n224 B.n223 585
R13 B.n222 B.n221 585
R14 B.n220 B.n219 585
R15 B.n218 B.n217 585
R16 B.n216 B.n215 585
R17 B.n214 B.n213 585
R18 B.n212 B.n211 585
R19 B.n210 B.n209 585
R20 B.n208 B.n207 585
R21 B.n206 B.n205 585
R22 B.n204 B.n203 585
R23 B.n202 B.n201 585
R24 B.n200 B.n199 585
R25 B.n198 B.n197 585
R26 B.n196 B.n195 585
R27 B.n194 B.n193 585
R28 B.n192 B.n191 585
R29 B.n190 B.n189 585
R30 B.n188 B.n187 585
R31 B.n186 B.n185 585
R32 B.n184 B.n183 585
R33 B.n181 B.n180 585
R34 B.n179 B.n178 585
R35 B.n177 B.n176 585
R36 B.n175 B.n174 585
R37 B.n173 B.n172 585
R38 B.n171 B.n170 585
R39 B.n169 B.n168 585
R40 B.n167 B.n166 585
R41 B.n165 B.n164 585
R42 B.n163 B.n162 585
R43 B.n160 B.n159 585
R44 B.n158 B.n157 585
R45 B.n156 B.n155 585
R46 B.n154 B.n153 585
R47 B.n152 B.n151 585
R48 B.n150 B.n149 585
R49 B.n148 B.n147 585
R50 B.n146 B.n145 585
R51 B.n144 B.n143 585
R52 B.n142 B.n141 585
R53 B.n140 B.n139 585
R54 B.n138 B.n137 585
R55 B.n136 B.n135 585
R56 B.n134 B.n133 585
R57 B.n132 B.n131 585
R58 B.n130 B.n129 585
R59 B.n128 B.n127 585
R60 B.n126 B.n125 585
R61 B.n124 B.n123 585
R62 B.n122 B.n121 585
R63 B.n120 B.n119 585
R64 B.n118 B.n117 585
R65 B.n116 B.n115 585
R66 B.n114 B.n113 585
R67 B.n112 B.n111 585
R68 B.n110 B.n109 585
R69 B.n108 B.n107 585
R70 B.n106 B.n105 585
R71 B.n104 B.n103 585
R72 B.n102 B.n101 585
R73 B.n100 B.n99 585
R74 B.n98 B.n97 585
R75 B.n53 B.n52 585
R76 B.n614 B.n54 585
R77 B.n619 B.n54 585
R78 B.n613 B.n612 585
R79 B.n612 B.n50 585
R80 B.n611 B.n49 585
R81 B.n625 B.n49 585
R82 B.n610 B.n48 585
R83 B.n626 B.n48 585
R84 B.n609 B.n47 585
R85 B.n627 B.n47 585
R86 B.n608 B.n607 585
R87 B.n607 B.n43 585
R88 B.n606 B.n42 585
R89 B.n633 B.n42 585
R90 B.n605 B.n41 585
R91 B.n634 B.n41 585
R92 B.n604 B.n40 585
R93 B.n635 B.n40 585
R94 B.n603 B.n602 585
R95 B.n602 B.n36 585
R96 B.n601 B.n35 585
R97 B.n641 B.n35 585
R98 B.n600 B.n34 585
R99 B.n642 B.n34 585
R100 B.n599 B.n33 585
R101 B.n643 B.n33 585
R102 B.n598 B.n597 585
R103 B.n597 B.n29 585
R104 B.n596 B.n28 585
R105 B.n649 B.n28 585
R106 B.n595 B.n27 585
R107 B.n650 B.n27 585
R108 B.n594 B.n26 585
R109 B.n651 B.n26 585
R110 B.n593 B.n592 585
R111 B.n592 B.n22 585
R112 B.n591 B.n21 585
R113 B.n657 B.n21 585
R114 B.n590 B.n20 585
R115 B.n658 B.n20 585
R116 B.n589 B.n19 585
R117 B.n659 B.n19 585
R118 B.n588 B.n587 585
R119 B.n587 B.n18 585
R120 B.n586 B.n14 585
R121 B.n665 B.n14 585
R122 B.n585 B.n13 585
R123 B.n666 B.n13 585
R124 B.n584 B.n12 585
R125 B.n667 B.n12 585
R126 B.n583 B.n582 585
R127 B.n582 B.n8 585
R128 B.n581 B.n7 585
R129 B.n673 B.n7 585
R130 B.n580 B.n6 585
R131 B.n674 B.n6 585
R132 B.n579 B.n5 585
R133 B.n675 B.n5 585
R134 B.n578 B.n577 585
R135 B.n577 B.n4 585
R136 B.n576 B.n246 585
R137 B.n576 B.n575 585
R138 B.n566 B.n247 585
R139 B.n248 B.n247 585
R140 B.n568 B.n567 585
R141 B.n569 B.n568 585
R142 B.n565 B.n253 585
R143 B.n253 B.n252 585
R144 B.n564 B.n563 585
R145 B.n563 B.n562 585
R146 B.n255 B.n254 585
R147 B.n555 B.n255 585
R148 B.n554 B.n553 585
R149 B.n556 B.n554 585
R150 B.n552 B.n260 585
R151 B.n260 B.n259 585
R152 B.n551 B.n550 585
R153 B.n550 B.n549 585
R154 B.n262 B.n261 585
R155 B.n263 B.n262 585
R156 B.n542 B.n541 585
R157 B.n543 B.n542 585
R158 B.n540 B.n268 585
R159 B.n268 B.n267 585
R160 B.n539 B.n538 585
R161 B.n538 B.n537 585
R162 B.n270 B.n269 585
R163 B.n271 B.n270 585
R164 B.n530 B.n529 585
R165 B.n531 B.n530 585
R166 B.n528 B.n276 585
R167 B.n276 B.n275 585
R168 B.n527 B.n526 585
R169 B.n526 B.n525 585
R170 B.n278 B.n277 585
R171 B.n279 B.n278 585
R172 B.n518 B.n517 585
R173 B.n519 B.n518 585
R174 B.n516 B.n284 585
R175 B.n284 B.n283 585
R176 B.n515 B.n514 585
R177 B.n514 B.n513 585
R178 B.n286 B.n285 585
R179 B.n287 B.n286 585
R180 B.n506 B.n505 585
R181 B.n507 B.n506 585
R182 B.n504 B.n292 585
R183 B.n292 B.n291 585
R184 B.n503 B.n502 585
R185 B.n502 B.n501 585
R186 B.n294 B.n293 585
R187 B.n295 B.n294 585
R188 B.n494 B.n493 585
R189 B.n495 B.n494 585
R190 B.n298 B.n297 585
R191 B.n345 B.n344 585
R192 B.n346 B.n342 585
R193 B.n342 B.n299 585
R194 B.n348 B.n347 585
R195 B.n350 B.n341 585
R196 B.n353 B.n352 585
R197 B.n354 B.n340 585
R198 B.n356 B.n355 585
R199 B.n358 B.n339 585
R200 B.n361 B.n360 585
R201 B.n362 B.n338 585
R202 B.n364 B.n363 585
R203 B.n366 B.n337 585
R204 B.n369 B.n368 585
R205 B.n370 B.n336 585
R206 B.n372 B.n371 585
R207 B.n374 B.n335 585
R208 B.n377 B.n376 585
R209 B.n378 B.n334 585
R210 B.n380 B.n379 585
R211 B.n382 B.n333 585
R212 B.n385 B.n384 585
R213 B.n386 B.n332 585
R214 B.n388 B.n387 585
R215 B.n390 B.n331 585
R216 B.n393 B.n392 585
R217 B.n394 B.n330 585
R218 B.n396 B.n395 585
R219 B.n398 B.n329 585
R220 B.n401 B.n400 585
R221 B.n402 B.n328 585
R222 B.n404 B.n403 585
R223 B.n406 B.n327 585
R224 B.n409 B.n408 585
R225 B.n410 B.n323 585
R226 B.n412 B.n411 585
R227 B.n414 B.n322 585
R228 B.n417 B.n416 585
R229 B.n418 B.n321 585
R230 B.n420 B.n419 585
R231 B.n422 B.n320 585
R232 B.n425 B.n424 585
R233 B.n426 B.n317 585
R234 B.n429 B.n428 585
R235 B.n431 B.n316 585
R236 B.n434 B.n433 585
R237 B.n435 B.n315 585
R238 B.n437 B.n436 585
R239 B.n439 B.n314 585
R240 B.n442 B.n441 585
R241 B.n443 B.n313 585
R242 B.n445 B.n444 585
R243 B.n447 B.n312 585
R244 B.n450 B.n449 585
R245 B.n451 B.n311 585
R246 B.n453 B.n452 585
R247 B.n455 B.n310 585
R248 B.n458 B.n457 585
R249 B.n459 B.n309 585
R250 B.n461 B.n460 585
R251 B.n463 B.n308 585
R252 B.n466 B.n465 585
R253 B.n467 B.n307 585
R254 B.n469 B.n468 585
R255 B.n471 B.n306 585
R256 B.n474 B.n473 585
R257 B.n475 B.n305 585
R258 B.n477 B.n476 585
R259 B.n479 B.n304 585
R260 B.n482 B.n481 585
R261 B.n483 B.n303 585
R262 B.n485 B.n484 585
R263 B.n487 B.n302 585
R264 B.n488 B.n301 585
R265 B.n491 B.n490 585
R266 B.n492 B.n300 585
R267 B.n300 B.n299 585
R268 B.n497 B.n496 585
R269 B.n496 B.n495 585
R270 B.n498 B.n296 585
R271 B.n296 B.n295 585
R272 B.n500 B.n499 585
R273 B.n501 B.n500 585
R274 B.n290 B.n289 585
R275 B.n291 B.n290 585
R276 B.n509 B.n508 585
R277 B.n508 B.n507 585
R278 B.n510 B.n288 585
R279 B.n288 B.n287 585
R280 B.n512 B.n511 585
R281 B.n513 B.n512 585
R282 B.n282 B.n281 585
R283 B.n283 B.n282 585
R284 B.n521 B.n520 585
R285 B.n520 B.n519 585
R286 B.n522 B.n280 585
R287 B.n280 B.n279 585
R288 B.n524 B.n523 585
R289 B.n525 B.n524 585
R290 B.n274 B.n273 585
R291 B.n275 B.n274 585
R292 B.n533 B.n532 585
R293 B.n532 B.n531 585
R294 B.n534 B.n272 585
R295 B.n272 B.n271 585
R296 B.n536 B.n535 585
R297 B.n537 B.n536 585
R298 B.n266 B.n265 585
R299 B.n267 B.n266 585
R300 B.n545 B.n544 585
R301 B.n544 B.n543 585
R302 B.n546 B.n264 585
R303 B.n264 B.n263 585
R304 B.n548 B.n547 585
R305 B.n549 B.n548 585
R306 B.n258 B.n257 585
R307 B.n259 B.n258 585
R308 B.n558 B.n557 585
R309 B.n557 B.n556 585
R310 B.n559 B.n256 585
R311 B.n555 B.n256 585
R312 B.n561 B.n560 585
R313 B.n562 B.n561 585
R314 B.n251 B.n250 585
R315 B.n252 B.n251 585
R316 B.n571 B.n570 585
R317 B.n570 B.n569 585
R318 B.n572 B.n249 585
R319 B.n249 B.n248 585
R320 B.n574 B.n573 585
R321 B.n575 B.n574 585
R322 B.n2 B.n0 585
R323 B.n4 B.n2 585
R324 B.n3 B.n1 585
R325 B.n674 B.n3 585
R326 B.n672 B.n671 585
R327 B.n673 B.n672 585
R328 B.n670 B.n9 585
R329 B.n9 B.n8 585
R330 B.n669 B.n668 585
R331 B.n668 B.n667 585
R332 B.n11 B.n10 585
R333 B.n666 B.n11 585
R334 B.n664 B.n663 585
R335 B.n665 B.n664 585
R336 B.n662 B.n15 585
R337 B.n18 B.n15 585
R338 B.n661 B.n660 585
R339 B.n660 B.n659 585
R340 B.n17 B.n16 585
R341 B.n658 B.n17 585
R342 B.n656 B.n655 585
R343 B.n657 B.n656 585
R344 B.n654 B.n23 585
R345 B.n23 B.n22 585
R346 B.n653 B.n652 585
R347 B.n652 B.n651 585
R348 B.n25 B.n24 585
R349 B.n650 B.n25 585
R350 B.n648 B.n647 585
R351 B.n649 B.n648 585
R352 B.n646 B.n30 585
R353 B.n30 B.n29 585
R354 B.n645 B.n644 585
R355 B.n644 B.n643 585
R356 B.n32 B.n31 585
R357 B.n642 B.n32 585
R358 B.n640 B.n639 585
R359 B.n641 B.n640 585
R360 B.n638 B.n37 585
R361 B.n37 B.n36 585
R362 B.n637 B.n636 585
R363 B.n636 B.n635 585
R364 B.n39 B.n38 585
R365 B.n634 B.n39 585
R366 B.n632 B.n631 585
R367 B.n633 B.n632 585
R368 B.n630 B.n44 585
R369 B.n44 B.n43 585
R370 B.n629 B.n628 585
R371 B.n628 B.n627 585
R372 B.n46 B.n45 585
R373 B.n626 B.n46 585
R374 B.n624 B.n623 585
R375 B.n625 B.n624 585
R376 B.n622 B.n51 585
R377 B.n51 B.n50 585
R378 B.n621 B.n620 585
R379 B.n620 B.n619 585
R380 B.n677 B.n676 585
R381 B.n676 B.n675 585
R382 B.n496 B.n298 545.355
R383 B.n620 B.n53 545.355
R384 B.n494 B.n300 545.355
R385 B.n616 B.n54 545.355
R386 B.n318 B.t5 299.548
R387 B.n93 B.t11 299.548
R388 B.n324 B.t8 299.548
R389 B.n95 B.t14 299.548
R390 B.n318 B.t2 280.882
R391 B.n324 B.t6 280.882
R392 B.n95 B.t13 280.882
R393 B.n93 B.t9 280.882
R394 B.n618 B.n617 256.663
R395 B.n618 B.n91 256.663
R396 B.n618 B.n90 256.663
R397 B.n618 B.n89 256.663
R398 B.n618 B.n88 256.663
R399 B.n618 B.n87 256.663
R400 B.n618 B.n86 256.663
R401 B.n618 B.n85 256.663
R402 B.n618 B.n84 256.663
R403 B.n618 B.n83 256.663
R404 B.n618 B.n82 256.663
R405 B.n618 B.n81 256.663
R406 B.n618 B.n80 256.663
R407 B.n618 B.n79 256.663
R408 B.n618 B.n78 256.663
R409 B.n618 B.n77 256.663
R410 B.n618 B.n76 256.663
R411 B.n618 B.n75 256.663
R412 B.n618 B.n74 256.663
R413 B.n618 B.n73 256.663
R414 B.n618 B.n72 256.663
R415 B.n618 B.n71 256.663
R416 B.n618 B.n70 256.663
R417 B.n618 B.n69 256.663
R418 B.n618 B.n68 256.663
R419 B.n618 B.n67 256.663
R420 B.n618 B.n66 256.663
R421 B.n618 B.n65 256.663
R422 B.n618 B.n64 256.663
R423 B.n618 B.n63 256.663
R424 B.n618 B.n62 256.663
R425 B.n618 B.n61 256.663
R426 B.n618 B.n60 256.663
R427 B.n618 B.n59 256.663
R428 B.n618 B.n58 256.663
R429 B.n618 B.n57 256.663
R430 B.n618 B.n56 256.663
R431 B.n618 B.n55 256.663
R432 B.n343 B.n299 256.663
R433 B.n349 B.n299 256.663
R434 B.n351 B.n299 256.663
R435 B.n357 B.n299 256.663
R436 B.n359 B.n299 256.663
R437 B.n365 B.n299 256.663
R438 B.n367 B.n299 256.663
R439 B.n373 B.n299 256.663
R440 B.n375 B.n299 256.663
R441 B.n381 B.n299 256.663
R442 B.n383 B.n299 256.663
R443 B.n389 B.n299 256.663
R444 B.n391 B.n299 256.663
R445 B.n397 B.n299 256.663
R446 B.n399 B.n299 256.663
R447 B.n405 B.n299 256.663
R448 B.n407 B.n299 256.663
R449 B.n413 B.n299 256.663
R450 B.n415 B.n299 256.663
R451 B.n421 B.n299 256.663
R452 B.n423 B.n299 256.663
R453 B.n430 B.n299 256.663
R454 B.n432 B.n299 256.663
R455 B.n438 B.n299 256.663
R456 B.n440 B.n299 256.663
R457 B.n446 B.n299 256.663
R458 B.n448 B.n299 256.663
R459 B.n454 B.n299 256.663
R460 B.n456 B.n299 256.663
R461 B.n462 B.n299 256.663
R462 B.n464 B.n299 256.663
R463 B.n470 B.n299 256.663
R464 B.n472 B.n299 256.663
R465 B.n478 B.n299 256.663
R466 B.n480 B.n299 256.663
R467 B.n486 B.n299 256.663
R468 B.n489 B.n299 256.663
R469 B.n319 B.t4 233.608
R470 B.n94 B.t12 233.608
R471 B.n325 B.t7 233.608
R472 B.n96 B.t15 233.608
R473 B.n496 B.n296 163.367
R474 B.n500 B.n296 163.367
R475 B.n500 B.n290 163.367
R476 B.n508 B.n290 163.367
R477 B.n508 B.n288 163.367
R478 B.n512 B.n288 163.367
R479 B.n512 B.n282 163.367
R480 B.n520 B.n282 163.367
R481 B.n520 B.n280 163.367
R482 B.n524 B.n280 163.367
R483 B.n524 B.n274 163.367
R484 B.n532 B.n274 163.367
R485 B.n532 B.n272 163.367
R486 B.n536 B.n272 163.367
R487 B.n536 B.n266 163.367
R488 B.n544 B.n266 163.367
R489 B.n544 B.n264 163.367
R490 B.n548 B.n264 163.367
R491 B.n548 B.n258 163.367
R492 B.n557 B.n258 163.367
R493 B.n557 B.n256 163.367
R494 B.n561 B.n256 163.367
R495 B.n561 B.n251 163.367
R496 B.n570 B.n251 163.367
R497 B.n570 B.n249 163.367
R498 B.n574 B.n249 163.367
R499 B.n574 B.n2 163.367
R500 B.n676 B.n2 163.367
R501 B.n676 B.n3 163.367
R502 B.n672 B.n3 163.367
R503 B.n672 B.n9 163.367
R504 B.n668 B.n9 163.367
R505 B.n668 B.n11 163.367
R506 B.n664 B.n11 163.367
R507 B.n664 B.n15 163.367
R508 B.n660 B.n15 163.367
R509 B.n660 B.n17 163.367
R510 B.n656 B.n17 163.367
R511 B.n656 B.n23 163.367
R512 B.n652 B.n23 163.367
R513 B.n652 B.n25 163.367
R514 B.n648 B.n25 163.367
R515 B.n648 B.n30 163.367
R516 B.n644 B.n30 163.367
R517 B.n644 B.n32 163.367
R518 B.n640 B.n32 163.367
R519 B.n640 B.n37 163.367
R520 B.n636 B.n37 163.367
R521 B.n636 B.n39 163.367
R522 B.n632 B.n39 163.367
R523 B.n632 B.n44 163.367
R524 B.n628 B.n44 163.367
R525 B.n628 B.n46 163.367
R526 B.n624 B.n46 163.367
R527 B.n624 B.n51 163.367
R528 B.n620 B.n51 163.367
R529 B.n344 B.n342 163.367
R530 B.n348 B.n342 163.367
R531 B.n352 B.n350 163.367
R532 B.n356 B.n340 163.367
R533 B.n360 B.n358 163.367
R534 B.n364 B.n338 163.367
R535 B.n368 B.n366 163.367
R536 B.n372 B.n336 163.367
R537 B.n376 B.n374 163.367
R538 B.n380 B.n334 163.367
R539 B.n384 B.n382 163.367
R540 B.n388 B.n332 163.367
R541 B.n392 B.n390 163.367
R542 B.n396 B.n330 163.367
R543 B.n400 B.n398 163.367
R544 B.n404 B.n328 163.367
R545 B.n408 B.n406 163.367
R546 B.n412 B.n323 163.367
R547 B.n416 B.n414 163.367
R548 B.n420 B.n321 163.367
R549 B.n424 B.n422 163.367
R550 B.n429 B.n317 163.367
R551 B.n433 B.n431 163.367
R552 B.n437 B.n315 163.367
R553 B.n441 B.n439 163.367
R554 B.n445 B.n313 163.367
R555 B.n449 B.n447 163.367
R556 B.n453 B.n311 163.367
R557 B.n457 B.n455 163.367
R558 B.n461 B.n309 163.367
R559 B.n465 B.n463 163.367
R560 B.n469 B.n307 163.367
R561 B.n473 B.n471 163.367
R562 B.n477 B.n305 163.367
R563 B.n481 B.n479 163.367
R564 B.n485 B.n303 163.367
R565 B.n488 B.n487 163.367
R566 B.n490 B.n300 163.367
R567 B.n494 B.n294 163.367
R568 B.n502 B.n294 163.367
R569 B.n502 B.n292 163.367
R570 B.n506 B.n292 163.367
R571 B.n506 B.n286 163.367
R572 B.n514 B.n286 163.367
R573 B.n514 B.n284 163.367
R574 B.n518 B.n284 163.367
R575 B.n518 B.n278 163.367
R576 B.n526 B.n278 163.367
R577 B.n526 B.n276 163.367
R578 B.n530 B.n276 163.367
R579 B.n530 B.n270 163.367
R580 B.n538 B.n270 163.367
R581 B.n538 B.n268 163.367
R582 B.n542 B.n268 163.367
R583 B.n542 B.n262 163.367
R584 B.n550 B.n262 163.367
R585 B.n550 B.n260 163.367
R586 B.n554 B.n260 163.367
R587 B.n554 B.n255 163.367
R588 B.n563 B.n255 163.367
R589 B.n563 B.n253 163.367
R590 B.n568 B.n253 163.367
R591 B.n568 B.n247 163.367
R592 B.n576 B.n247 163.367
R593 B.n577 B.n576 163.367
R594 B.n577 B.n5 163.367
R595 B.n6 B.n5 163.367
R596 B.n7 B.n6 163.367
R597 B.n582 B.n7 163.367
R598 B.n582 B.n12 163.367
R599 B.n13 B.n12 163.367
R600 B.n14 B.n13 163.367
R601 B.n587 B.n14 163.367
R602 B.n587 B.n19 163.367
R603 B.n20 B.n19 163.367
R604 B.n21 B.n20 163.367
R605 B.n592 B.n21 163.367
R606 B.n592 B.n26 163.367
R607 B.n27 B.n26 163.367
R608 B.n28 B.n27 163.367
R609 B.n597 B.n28 163.367
R610 B.n597 B.n33 163.367
R611 B.n34 B.n33 163.367
R612 B.n35 B.n34 163.367
R613 B.n602 B.n35 163.367
R614 B.n602 B.n40 163.367
R615 B.n41 B.n40 163.367
R616 B.n42 B.n41 163.367
R617 B.n607 B.n42 163.367
R618 B.n607 B.n47 163.367
R619 B.n48 B.n47 163.367
R620 B.n49 B.n48 163.367
R621 B.n612 B.n49 163.367
R622 B.n612 B.n54 163.367
R623 B.n99 B.n98 163.367
R624 B.n103 B.n102 163.367
R625 B.n107 B.n106 163.367
R626 B.n111 B.n110 163.367
R627 B.n115 B.n114 163.367
R628 B.n119 B.n118 163.367
R629 B.n123 B.n122 163.367
R630 B.n127 B.n126 163.367
R631 B.n131 B.n130 163.367
R632 B.n135 B.n134 163.367
R633 B.n139 B.n138 163.367
R634 B.n143 B.n142 163.367
R635 B.n147 B.n146 163.367
R636 B.n151 B.n150 163.367
R637 B.n155 B.n154 163.367
R638 B.n159 B.n158 163.367
R639 B.n164 B.n163 163.367
R640 B.n168 B.n167 163.367
R641 B.n172 B.n171 163.367
R642 B.n176 B.n175 163.367
R643 B.n180 B.n179 163.367
R644 B.n185 B.n184 163.367
R645 B.n189 B.n188 163.367
R646 B.n193 B.n192 163.367
R647 B.n197 B.n196 163.367
R648 B.n201 B.n200 163.367
R649 B.n205 B.n204 163.367
R650 B.n209 B.n208 163.367
R651 B.n213 B.n212 163.367
R652 B.n217 B.n216 163.367
R653 B.n221 B.n220 163.367
R654 B.n225 B.n224 163.367
R655 B.n229 B.n228 163.367
R656 B.n233 B.n232 163.367
R657 B.n237 B.n236 163.367
R658 B.n241 B.n240 163.367
R659 B.n243 B.n92 163.367
R660 B.n495 B.n299 99.5515
R661 B.n619 B.n618 99.5515
R662 B.n343 B.n298 71.676
R663 B.n349 B.n348 71.676
R664 B.n352 B.n351 71.676
R665 B.n357 B.n356 71.676
R666 B.n360 B.n359 71.676
R667 B.n365 B.n364 71.676
R668 B.n368 B.n367 71.676
R669 B.n373 B.n372 71.676
R670 B.n376 B.n375 71.676
R671 B.n381 B.n380 71.676
R672 B.n384 B.n383 71.676
R673 B.n389 B.n388 71.676
R674 B.n392 B.n391 71.676
R675 B.n397 B.n396 71.676
R676 B.n400 B.n399 71.676
R677 B.n405 B.n404 71.676
R678 B.n408 B.n407 71.676
R679 B.n413 B.n412 71.676
R680 B.n416 B.n415 71.676
R681 B.n421 B.n420 71.676
R682 B.n424 B.n423 71.676
R683 B.n430 B.n429 71.676
R684 B.n433 B.n432 71.676
R685 B.n438 B.n437 71.676
R686 B.n441 B.n440 71.676
R687 B.n446 B.n445 71.676
R688 B.n449 B.n448 71.676
R689 B.n454 B.n453 71.676
R690 B.n457 B.n456 71.676
R691 B.n462 B.n461 71.676
R692 B.n465 B.n464 71.676
R693 B.n470 B.n469 71.676
R694 B.n473 B.n472 71.676
R695 B.n478 B.n477 71.676
R696 B.n481 B.n480 71.676
R697 B.n486 B.n485 71.676
R698 B.n489 B.n488 71.676
R699 B.n55 B.n53 71.676
R700 B.n99 B.n56 71.676
R701 B.n103 B.n57 71.676
R702 B.n107 B.n58 71.676
R703 B.n111 B.n59 71.676
R704 B.n115 B.n60 71.676
R705 B.n119 B.n61 71.676
R706 B.n123 B.n62 71.676
R707 B.n127 B.n63 71.676
R708 B.n131 B.n64 71.676
R709 B.n135 B.n65 71.676
R710 B.n139 B.n66 71.676
R711 B.n143 B.n67 71.676
R712 B.n147 B.n68 71.676
R713 B.n151 B.n69 71.676
R714 B.n155 B.n70 71.676
R715 B.n159 B.n71 71.676
R716 B.n164 B.n72 71.676
R717 B.n168 B.n73 71.676
R718 B.n172 B.n74 71.676
R719 B.n176 B.n75 71.676
R720 B.n180 B.n76 71.676
R721 B.n185 B.n77 71.676
R722 B.n189 B.n78 71.676
R723 B.n193 B.n79 71.676
R724 B.n197 B.n80 71.676
R725 B.n201 B.n81 71.676
R726 B.n205 B.n82 71.676
R727 B.n209 B.n83 71.676
R728 B.n213 B.n84 71.676
R729 B.n217 B.n85 71.676
R730 B.n221 B.n86 71.676
R731 B.n225 B.n87 71.676
R732 B.n229 B.n88 71.676
R733 B.n233 B.n89 71.676
R734 B.n237 B.n90 71.676
R735 B.n241 B.n91 71.676
R736 B.n617 B.n92 71.676
R737 B.n617 B.n616 71.676
R738 B.n243 B.n91 71.676
R739 B.n240 B.n90 71.676
R740 B.n236 B.n89 71.676
R741 B.n232 B.n88 71.676
R742 B.n228 B.n87 71.676
R743 B.n224 B.n86 71.676
R744 B.n220 B.n85 71.676
R745 B.n216 B.n84 71.676
R746 B.n212 B.n83 71.676
R747 B.n208 B.n82 71.676
R748 B.n204 B.n81 71.676
R749 B.n200 B.n80 71.676
R750 B.n196 B.n79 71.676
R751 B.n192 B.n78 71.676
R752 B.n188 B.n77 71.676
R753 B.n184 B.n76 71.676
R754 B.n179 B.n75 71.676
R755 B.n175 B.n74 71.676
R756 B.n171 B.n73 71.676
R757 B.n167 B.n72 71.676
R758 B.n163 B.n71 71.676
R759 B.n158 B.n70 71.676
R760 B.n154 B.n69 71.676
R761 B.n150 B.n68 71.676
R762 B.n146 B.n67 71.676
R763 B.n142 B.n66 71.676
R764 B.n138 B.n65 71.676
R765 B.n134 B.n64 71.676
R766 B.n130 B.n63 71.676
R767 B.n126 B.n62 71.676
R768 B.n122 B.n61 71.676
R769 B.n118 B.n60 71.676
R770 B.n114 B.n59 71.676
R771 B.n110 B.n58 71.676
R772 B.n106 B.n57 71.676
R773 B.n102 B.n56 71.676
R774 B.n98 B.n55 71.676
R775 B.n344 B.n343 71.676
R776 B.n350 B.n349 71.676
R777 B.n351 B.n340 71.676
R778 B.n358 B.n357 71.676
R779 B.n359 B.n338 71.676
R780 B.n366 B.n365 71.676
R781 B.n367 B.n336 71.676
R782 B.n374 B.n373 71.676
R783 B.n375 B.n334 71.676
R784 B.n382 B.n381 71.676
R785 B.n383 B.n332 71.676
R786 B.n390 B.n389 71.676
R787 B.n391 B.n330 71.676
R788 B.n398 B.n397 71.676
R789 B.n399 B.n328 71.676
R790 B.n406 B.n405 71.676
R791 B.n407 B.n323 71.676
R792 B.n414 B.n413 71.676
R793 B.n415 B.n321 71.676
R794 B.n422 B.n421 71.676
R795 B.n423 B.n317 71.676
R796 B.n431 B.n430 71.676
R797 B.n432 B.n315 71.676
R798 B.n439 B.n438 71.676
R799 B.n440 B.n313 71.676
R800 B.n447 B.n446 71.676
R801 B.n448 B.n311 71.676
R802 B.n455 B.n454 71.676
R803 B.n456 B.n309 71.676
R804 B.n463 B.n462 71.676
R805 B.n464 B.n307 71.676
R806 B.n471 B.n470 71.676
R807 B.n472 B.n305 71.676
R808 B.n479 B.n478 71.676
R809 B.n480 B.n303 71.676
R810 B.n487 B.n486 71.676
R811 B.n490 B.n489 71.676
R812 B.n319 B.n318 65.9399
R813 B.n325 B.n324 65.9399
R814 B.n96 B.n95 65.9399
R815 B.n94 B.n93 65.9399
R816 B.n427 B.n319 59.5399
R817 B.n326 B.n325 59.5399
R818 B.n161 B.n96 59.5399
R819 B.n182 B.n94 59.5399
R820 B.n495 B.n295 51.6758
R821 B.n501 B.n295 51.6758
R822 B.n501 B.n291 51.6758
R823 B.n507 B.n291 51.6758
R824 B.n507 B.n287 51.6758
R825 B.n513 B.n287 51.6758
R826 B.n513 B.n283 51.6758
R827 B.n519 B.n283 51.6758
R828 B.n525 B.n279 51.6758
R829 B.n525 B.n275 51.6758
R830 B.n531 B.n275 51.6758
R831 B.n531 B.n271 51.6758
R832 B.n537 B.n271 51.6758
R833 B.n537 B.n267 51.6758
R834 B.n543 B.n267 51.6758
R835 B.n543 B.n263 51.6758
R836 B.n549 B.n263 51.6758
R837 B.n549 B.n259 51.6758
R838 B.n556 B.n259 51.6758
R839 B.n556 B.n555 51.6758
R840 B.n562 B.n252 51.6758
R841 B.n569 B.n252 51.6758
R842 B.n569 B.n248 51.6758
R843 B.n575 B.n248 51.6758
R844 B.n575 B.n4 51.6758
R845 B.n675 B.n4 51.6758
R846 B.n675 B.n674 51.6758
R847 B.n674 B.n673 51.6758
R848 B.n673 B.n8 51.6758
R849 B.n667 B.n8 51.6758
R850 B.n667 B.n666 51.6758
R851 B.n666 B.n665 51.6758
R852 B.n659 B.n18 51.6758
R853 B.n659 B.n658 51.6758
R854 B.n658 B.n657 51.6758
R855 B.n657 B.n22 51.6758
R856 B.n651 B.n22 51.6758
R857 B.n651 B.n650 51.6758
R858 B.n650 B.n649 51.6758
R859 B.n649 B.n29 51.6758
R860 B.n643 B.n29 51.6758
R861 B.n643 B.n642 51.6758
R862 B.n642 B.n641 51.6758
R863 B.n641 B.n36 51.6758
R864 B.n635 B.n634 51.6758
R865 B.n634 B.n633 51.6758
R866 B.n633 B.n43 51.6758
R867 B.n627 B.n43 51.6758
R868 B.n627 B.n626 51.6758
R869 B.n626 B.n625 51.6758
R870 B.n625 B.n50 51.6758
R871 B.n619 B.n50 51.6758
R872 B.t3 B.n279 41.7967
R873 B.t10 B.n36 41.7967
R874 B.n621 B.n52 35.4346
R875 B.n493 B.n492 35.4346
R876 B.n497 B.n297 35.4346
R877 B.n615 B.n614 35.4346
R878 B.n562 B.t0 31.1577
R879 B.n665 B.t1 31.1577
R880 B.n555 B.t0 20.5186
R881 B.n18 B.t1 20.5186
R882 B B.n677 18.0485
R883 B.n97 B.n52 10.6151
R884 B.n100 B.n97 10.6151
R885 B.n101 B.n100 10.6151
R886 B.n104 B.n101 10.6151
R887 B.n105 B.n104 10.6151
R888 B.n108 B.n105 10.6151
R889 B.n109 B.n108 10.6151
R890 B.n112 B.n109 10.6151
R891 B.n113 B.n112 10.6151
R892 B.n116 B.n113 10.6151
R893 B.n117 B.n116 10.6151
R894 B.n120 B.n117 10.6151
R895 B.n121 B.n120 10.6151
R896 B.n124 B.n121 10.6151
R897 B.n125 B.n124 10.6151
R898 B.n128 B.n125 10.6151
R899 B.n129 B.n128 10.6151
R900 B.n132 B.n129 10.6151
R901 B.n133 B.n132 10.6151
R902 B.n136 B.n133 10.6151
R903 B.n137 B.n136 10.6151
R904 B.n140 B.n137 10.6151
R905 B.n141 B.n140 10.6151
R906 B.n144 B.n141 10.6151
R907 B.n145 B.n144 10.6151
R908 B.n148 B.n145 10.6151
R909 B.n149 B.n148 10.6151
R910 B.n152 B.n149 10.6151
R911 B.n153 B.n152 10.6151
R912 B.n156 B.n153 10.6151
R913 B.n157 B.n156 10.6151
R914 B.n160 B.n157 10.6151
R915 B.n165 B.n162 10.6151
R916 B.n166 B.n165 10.6151
R917 B.n169 B.n166 10.6151
R918 B.n170 B.n169 10.6151
R919 B.n173 B.n170 10.6151
R920 B.n174 B.n173 10.6151
R921 B.n177 B.n174 10.6151
R922 B.n178 B.n177 10.6151
R923 B.n181 B.n178 10.6151
R924 B.n186 B.n183 10.6151
R925 B.n187 B.n186 10.6151
R926 B.n190 B.n187 10.6151
R927 B.n191 B.n190 10.6151
R928 B.n194 B.n191 10.6151
R929 B.n195 B.n194 10.6151
R930 B.n198 B.n195 10.6151
R931 B.n199 B.n198 10.6151
R932 B.n202 B.n199 10.6151
R933 B.n203 B.n202 10.6151
R934 B.n206 B.n203 10.6151
R935 B.n207 B.n206 10.6151
R936 B.n210 B.n207 10.6151
R937 B.n211 B.n210 10.6151
R938 B.n214 B.n211 10.6151
R939 B.n215 B.n214 10.6151
R940 B.n218 B.n215 10.6151
R941 B.n219 B.n218 10.6151
R942 B.n222 B.n219 10.6151
R943 B.n223 B.n222 10.6151
R944 B.n226 B.n223 10.6151
R945 B.n227 B.n226 10.6151
R946 B.n230 B.n227 10.6151
R947 B.n231 B.n230 10.6151
R948 B.n234 B.n231 10.6151
R949 B.n235 B.n234 10.6151
R950 B.n238 B.n235 10.6151
R951 B.n239 B.n238 10.6151
R952 B.n242 B.n239 10.6151
R953 B.n244 B.n242 10.6151
R954 B.n245 B.n244 10.6151
R955 B.n615 B.n245 10.6151
R956 B.n493 B.n293 10.6151
R957 B.n503 B.n293 10.6151
R958 B.n504 B.n503 10.6151
R959 B.n505 B.n504 10.6151
R960 B.n505 B.n285 10.6151
R961 B.n515 B.n285 10.6151
R962 B.n516 B.n515 10.6151
R963 B.n517 B.n516 10.6151
R964 B.n517 B.n277 10.6151
R965 B.n527 B.n277 10.6151
R966 B.n528 B.n527 10.6151
R967 B.n529 B.n528 10.6151
R968 B.n529 B.n269 10.6151
R969 B.n539 B.n269 10.6151
R970 B.n540 B.n539 10.6151
R971 B.n541 B.n540 10.6151
R972 B.n541 B.n261 10.6151
R973 B.n551 B.n261 10.6151
R974 B.n552 B.n551 10.6151
R975 B.n553 B.n552 10.6151
R976 B.n553 B.n254 10.6151
R977 B.n564 B.n254 10.6151
R978 B.n565 B.n564 10.6151
R979 B.n567 B.n565 10.6151
R980 B.n567 B.n566 10.6151
R981 B.n566 B.n246 10.6151
R982 B.n578 B.n246 10.6151
R983 B.n579 B.n578 10.6151
R984 B.n580 B.n579 10.6151
R985 B.n581 B.n580 10.6151
R986 B.n583 B.n581 10.6151
R987 B.n584 B.n583 10.6151
R988 B.n585 B.n584 10.6151
R989 B.n586 B.n585 10.6151
R990 B.n588 B.n586 10.6151
R991 B.n589 B.n588 10.6151
R992 B.n590 B.n589 10.6151
R993 B.n591 B.n590 10.6151
R994 B.n593 B.n591 10.6151
R995 B.n594 B.n593 10.6151
R996 B.n595 B.n594 10.6151
R997 B.n596 B.n595 10.6151
R998 B.n598 B.n596 10.6151
R999 B.n599 B.n598 10.6151
R1000 B.n600 B.n599 10.6151
R1001 B.n601 B.n600 10.6151
R1002 B.n603 B.n601 10.6151
R1003 B.n604 B.n603 10.6151
R1004 B.n605 B.n604 10.6151
R1005 B.n606 B.n605 10.6151
R1006 B.n608 B.n606 10.6151
R1007 B.n609 B.n608 10.6151
R1008 B.n610 B.n609 10.6151
R1009 B.n611 B.n610 10.6151
R1010 B.n613 B.n611 10.6151
R1011 B.n614 B.n613 10.6151
R1012 B.n345 B.n297 10.6151
R1013 B.n346 B.n345 10.6151
R1014 B.n347 B.n346 10.6151
R1015 B.n347 B.n341 10.6151
R1016 B.n353 B.n341 10.6151
R1017 B.n354 B.n353 10.6151
R1018 B.n355 B.n354 10.6151
R1019 B.n355 B.n339 10.6151
R1020 B.n361 B.n339 10.6151
R1021 B.n362 B.n361 10.6151
R1022 B.n363 B.n362 10.6151
R1023 B.n363 B.n337 10.6151
R1024 B.n369 B.n337 10.6151
R1025 B.n370 B.n369 10.6151
R1026 B.n371 B.n370 10.6151
R1027 B.n371 B.n335 10.6151
R1028 B.n377 B.n335 10.6151
R1029 B.n378 B.n377 10.6151
R1030 B.n379 B.n378 10.6151
R1031 B.n379 B.n333 10.6151
R1032 B.n385 B.n333 10.6151
R1033 B.n386 B.n385 10.6151
R1034 B.n387 B.n386 10.6151
R1035 B.n387 B.n331 10.6151
R1036 B.n393 B.n331 10.6151
R1037 B.n394 B.n393 10.6151
R1038 B.n395 B.n394 10.6151
R1039 B.n395 B.n329 10.6151
R1040 B.n401 B.n329 10.6151
R1041 B.n402 B.n401 10.6151
R1042 B.n403 B.n402 10.6151
R1043 B.n403 B.n327 10.6151
R1044 B.n410 B.n409 10.6151
R1045 B.n411 B.n410 10.6151
R1046 B.n411 B.n322 10.6151
R1047 B.n417 B.n322 10.6151
R1048 B.n418 B.n417 10.6151
R1049 B.n419 B.n418 10.6151
R1050 B.n419 B.n320 10.6151
R1051 B.n425 B.n320 10.6151
R1052 B.n426 B.n425 10.6151
R1053 B.n428 B.n316 10.6151
R1054 B.n434 B.n316 10.6151
R1055 B.n435 B.n434 10.6151
R1056 B.n436 B.n435 10.6151
R1057 B.n436 B.n314 10.6151
R1058 B.n442 B.n314 10.6151
R1059 B.n443 B.n442 10.6151
R1060 B.n444 B.n443 10.6151
R1061 B.n444 B.n312 10.6151
R1062 B.n450 B.n312 10.6151
R1063 B.n451 B.n450 10.6151
R1064 B.n452 B.n451 10.6151
R1065 B.n452 B.n310 10.6151
R1066 B.n458 B.n310 10.6151
R1067 B.n459 B.n458 10.6151
R1068 B.n460 B.n459 10.6151
R1069 B.n460 B.n308 10.6151
R1070 B.n466 B.n308 10.6151
R1071 B.n467 B.n466 10.6151
R1072 B.n468 B.n467 10.6151
R1073 B.n468 B.n306 10.6151
R1074 B.n474 B.n306 10.6151
R1075 B.n475 B.n474 10.6151
R1076 B.n476 B.n475 10.6151
R1077 B.n476 B.n304 10.6151
R1078 B.n482 B.n304 10.6151
R1079 B.n483 B.n482 10.6151
R1080 B.n484 B.n483 10.6151
R1081 B.n484 B.n302 10.6151
R1082 B.n302 B.n301 10.6151
R1083 B.n491 B.n301 10.6151
R1084 B.n492 B.n491 10.6151
R1085 B.n498 B.n497 10.6151
R1086 B.n499 B.n498 10.6151
R1087 B.n499 B.n289 10.6151
R1088 B.n509 B.n289 10.6151
R1089 B.n510 B.n509 10.6151
R1090 B.n511 B.n510 10.6151
R1091 B.n511 B.n281 10.6151
R1092 B.n521 B.n281 10.6151
R1093 B.n522 B.n521 10.6151
R1094 B.n523 B.n522 10.6151
R1095 B.n523 B.n273 10.6151
R1096 B.n533 B.n273 10.6151
R1097 B.n534 B.n533 10.6151
R1098 B.n535 B.n534 10.6151
R1099 B.n535 B.n265 10.6151
R1100 B.n545 B.n265 10.6151
R1101 B.n546 B.n545 10.6151
R1102 B.n547 B.n546 10.6151
R1103 B.n547 B.n257 10.6151
R1104 B.n558 B.n257 10.6151
R1105 B.n559 B.n558 10.6151
R1106 B.n560 B.n559 10.6151
R1107 B.n560 B.n250 10.6151
R1108 B.n571 B.n250 10.6151
R1109 B.n572 B.n571 10.6151
R1110 B.n573 B.n572 10.6151
R1111 B.n573 B.n0 10.6151
R1112 B.n671 B.n1 10.6151
R1113 B.n671 B.n670 10.6151
R1114 B.n670 B.n669 10.6151
R1115 B.n669 B.n10 10.6151
R1116 B.n663 B.n10 10.6151
R1117 B.n663 B.n662 10.6151
R1118 B.n662 B.n661 10.6151
R1119 B.n661 B.n16 10.6151
R1120 B.n655 B.n16 10.6151
R1121 B.n655 B.n654 10.6151
R1122 B.n654 B.n653 10.6151
R1123 B.n653 B.n24 10.6151
R1124 B.n647 B.n24 10.6151
R1125 B.n647 B.n646 10.6151
R1126 B.n646 B.n645 10.6151
R1127 B.n645 B.n31 10.6151
R1128 B.n639 B.n31 10.6151
R1129 B.n639 B.n638 10.6151
R1130 B.n638 B.n637 10.6151
R1131 B.n637 B.n38 10.6151
R1132 B.n631 B.n38 10.6151
R1133 B.n631 B.n630 10.6151
R1134 B.n630 B.n629 10.6151
R1135 B.n629 B.n45 10.6151
R1136 B.n623 B.n45 10.6151
R1137 B.n623 B.n622 10.6151
R1138 B.n622 B.n621 10.6151
R1139 B.n519 B.t3 9.8796
R1140 B.n635 B.t10 9.8796
R1141 B.n161 B.n160 9.36635
R1142 B.n183 B.n182 9.36635
R1143 B.n327 B.n326 9.36635
R1144 B.n428 B.n427 9.36635
R1145 B.n677 B.n0 2.81026
R1146 B.n677 B.n1 2.81026
R1147 B.n162 B.n161 1.24928
R1148 B.n182 B.n181 1.24928
R1149 B.n409 B.n326 1.24928
R1150 B.n427 B.n426 1.24928
R1151 VP.n0 VP.t0 157.142
R1152 VP.n0 VP.t1 113.359
R1153 VP VP.n0 0.431812
R1154 VTAIL.n194 VTAIL.n150 289.615
R1155 VTAIL.n44 VTAIL.n0 289.615
R1156 VTAIL.n144 VTAIL.n100 289.615
R1157 VTAIL.n94 VTAIL.n50 289.615
R1158 VTAIL.n167 VTAIL.n166 185
R1159 VTAIL.n169 VTAIL.n168 185
R1160 VTAIL.n162 VTAIL.n161 185
R1161 VTAIL.n175 VTAIL.n174 185
R1162 VTAIL.n177 VTAIL.n176 185
R1163 VTAIL.n158 VTAIL.n157 185
R1164 VTAIL.n184 VTAIL.n183 185
R1165 VTAIL.n185 VTAIL.n156 185
R1166 VTAIL.n187 VTAIL.n186 185
R1167 VTAIL.n154 VTAIL.n153 185
R1168 VTAIL.n193 VTAIL.n192 185
R1169 VTAIL.n195 VTAIL.n194 185
R1170 VTAIL.n17 VTAIL.n16 185
R1171 VTAIL.n19 VTAIL.n18 185
R1172 VTAIL.n12 VTAIL.n11 185
R1173 VTAIL.n25 VTAIL.n24 185
R1174 VTAIL.n27 VTAIL.n26 185
R1175 VTAIL.n8 VTAIL.n7 185
R1176 VTAIL.n34 VTAIL.n33 185
R1177 VTAIL.n35 VTAIL.n6 185
R1178 VTAIL.n37 VTAIL.n36 185
R1179 VTAIL.n4 VTAIL.n3 185
R1180 VTAIL.n43 VTAIL.n42 185
R1181 VTAIL.n45 VTAIL.n44 185
R1182 VTAIL.n145 VTAIL.n144 185
R1183 VTAIL.n143 VTAIL.n142 185
R1184 VTAIL.n104 VTAIL.n103 185
R1185 VTAIL.n108 VTAIL.n106 185
R1186 VTAIL.n137 VTAIL.n136 185
R1187 VTAIL.n135 VTAIL.n134 185
R1188 VTAIL.n110 VTAIL.n109 185
R1189 VTAIL.n129 VTAIL.n128 185
R1190 VTAIL.n127 VTAIL.n126 185
R1191 VTAIL.n114 VTAIL.n113 185
R1192 VTAIL.n121 VTAIL.n120 185
R1193 VTAIL.n119 VTAIL.n118 185
R1194 VTAIL.n95 VTAIL.n94 185
R1195 VTAIL.n93 VTAIL.n92 185
R1196 VTAIL.n54 VTAIL.n53 185
R1197 VTAIL.n58 VTAIL.n56 185
R1198 VTAIL.n87 VTAIL.n86 185
R1199 VTAIL.n85 VTAIL.n84 185
R1200 VTAIL.n60 VTAIL.n59 185
R1201 VTAIL.n79 VTAIL.n78 185
R1202 VTAIL.n77 VTAIL.n76 185
R1203 VTAIL.n64 VTAIL.n63 185
R1204 VTAIL.n71 VTAIL.n70 185
R1205 VTAIL.n69 VTAIL.n68 185
R1206 VTAIL.n165 VTAIL.t1 149.524
R1207 VTAIL.n15 VTAIL.t2 149.524
R1208 VTAIL.n117 VTAIL.t3 149.524
R1209 VTAIL.n67 VTAIL.t0 149.524
R1210 VTAIL.n168 VTAIL.n167 104.615
R1211 VTAIL.n168 VTAIL.n161 104.615
R1212 VTAIL.n175 VTAIL.n161 104.615
R1213 VTAIL.n176 VTAIL.n175 104.615
R1214 VTAIL.n176 VTAIL.n157 104.615
R1215 VTAIL.n184 VTAIL.n157 104.615
R1216 VTAIL.n185 VTAIL.n184 104.615
R1217 VTAIL.n186 VTAIL.n185 104.615
R1218 VTAIL.n186 VTAIL.n153 104.615
R1219 VTAIL.n193 VTAIL.n153 104.615
R1220 VTAIL.n194 VTAIL.n193 104.615
R1221 VTAIL.n18 VTAIL.n17 104.615
R1222 VTAIL.n18 VTAIL.n11 104.615
R1223 VTAIL.n25 VTAIL.n11 104.615
R1224 VTAIL.n26 VTAIL.n25 104.615
R1225 VTAIL.n26 VTAIL.n7 104.615
R1226 VTAIL.n34 VTAIL.n7 104.615
R1227 VTAIL.n35 VTAIL.n34 104.615
R1228 VTAIL.n36 VTAIL.n35 104.615
R1229 VTAIL.n36 VTAIL.n3 104.615
R1230 VTAIL.n43 VTAIL.n3 104.615
R1231 VTAIL.n44 VTAIL.n43 104.615
R1232 VTAIL.n144 VTAIL.n143 104.615
R1233 VTAIL.n143 VTAIL.n103 104.615
R1234 VTAIL.n108 VTAIL.n103 104.615
R1235 VTAIL.n136 VTAIL.n108 104.615
R1236 VTAIL.n136 VTAIL.n135 104.615
R1237 VTAIL.n135 VTAIL.n109 104.615
R1238 VTAIL.n128 VTAIL.n109 104.615
R1239 VTAIL.n128 VTAIL.n127 104.615
R1240 VTAIL.n127 VTAIL.n113 104.615
R1241 VTAIL.n120 VTAIL.n113 104.615
R1242 VTAIL.n120 VTAIL.n119 104.615
R1243 VTAIL.n94 VTAIL.n93 104.615
R1244 VTAIL.n93 VTAIL.n53 104.615
R1245 VTAIL.n58 VTAIL.n53 104.615
R1246 VTAIL.n86 VTAIL.n58 104.615
R1247 VTAIL.n86 VTAIL.n85 104.615
R1248 VTAIL.n85 VTAIL.n59 104.615
R1249 VTAIL.n78 VTAIL.n59 104.615
R1250 VTAIL.n78 VTAIL.n77 104.615
R1251 VTAIL.n77 VTAIL.n63 104.615
R1252 VTAIL.n70 VTAIL.n63 104.615
R1253 VTAIL.n70 VTAIL.n69 104.615
R1254 VTAIL.n167 VTAIL.t1 52.3082
R1255 VTAIL.n17 VTAIL.t2 52.3082
R1256 VTAIL.n119 VTAIL.t3 52.3082
R1257 VTAIL.n69 VTAIL.t0 52.3082
R1258 VTAIL.n199 VTAIL.n198 31.4096
R1259 VTAIL.n49 VTAIL.n48 31.4096
R1260 VTAIL.n149 VTAIL.n148 31.4096
R1261 VTAIL.n99 VTAIL.n98 31.4096
R1262 VTAIL.n99 VTAIL.n49 26.16
R1263 VTAIL.n199 VTAIL.n149 23.2289
R1264 VTAIL.n187 VTAIL.n154 13.1884
R1265 VTAIL.n37 VTAIL.n4 13.1884
R1266 VTAIL.n106 VTAIL.n104 13.1884
R1267 VTAIL.n56 VTAIL.n54 13.1884
R1268 VTAIL.n188 VTAIL.n156 12.8005
R1269 VTAIL.n192 VTAIL.n191 12.8005
R1270 VTAIL.n38 VTAIL.n6 12.8005
R1271 VTAIL.n42 VTAIL.n41 12.8005
R1272 VTAIL.n142 VTAIL.n141 12.8005
R1273 VTAIL.n138 VTAIL.n137 12.8005
R1274 VTAIL.n92 VTAIL.n91 12.8005
R1275 VTAIL.n88 VTAIL.n87 12.8005
R1276 VTAIL.n183 VTAIL.n182 12.0247
R1277 VTAIL.n195 VTAIL.n152 12.0247
R1278 VTAIL.n33 VTAIL.n32 12.0247
R1279 VTAIL.n45 VTAIL.n2 12.0247
R1280 VTAIL.n145 VTAIL.n102 12.0247
R1281 VTAIL.n134 VTAIL.n107 12.0247
R1282 VTAIL.n95 VTAIL.n52 12.0247
R1283 VTAIL.n84 VTAIL.n57 12.0247
R1284 VTAIL.n181 VTAIL.n158 11.249
R1285 VTAIL.n196 VTAIL.n150 11.249
R1286 VTAIL.n31 VTAIL.n8 11.249
R1287 VTAIL.n46 VTAIL.n0 11.249
R1288 VTAIL.n146 VTAIL.n100 11.249
R1289 VTAIL.n133 VTAIL.n110 11.249
R1290 VTAIL.n96 VTAIL.n50 11.249
R1291 VTAIL.n83 VTAIL.n60 11.249
R1292 VTAIL.n178 VTAIL.n177 10.4732
R1293 VTAIL.n28 VTAIL.n27 10.4732
R1294 VTAIL.n130 VTAIL.n129 10.4732
R1295 VTAIL.n80 VTAIL.n79 10.4732
R1296 VTAIL.n166 VTAIL.n165 10.2747
R1297 VTAIL.n16 VTAIL.n15 10.2747
R1298 VTAIL.n118 VTAIL.n117 10.2747
R1299 VTAIL.n68 VTAIL.n67 10.2747
R1300 VTAIL.n174 VTAIL.n160 9.69747
R1301 VTAIL.n24 VTAIL.n10 9.69747
R1302 VTAIL.n126 VTAIL.n112 9.69747
R1303 VTAIL.n76 VTAIL.n62 9.69747
R1304 VTAIL.n198 VTAIL.n197 9.45567
R1305 VTAIL.n48 VTAIL.n47 9.45567
R1306 VTAIL.n148 VTAIL.n147 9.45567
R1307 VTAIL.n98 VTAIL.n97 9.45567
R1308 VTAIL.n197 VTAIL.n196 9.3005
R1309 VTAIL.n152 VTAIL.n151 9.3005
R1310 VTAIL.n191 VTAIL.n190 9.3005
R1311 VTAIL.n164 VTAIL.n163 9.3005
R1312 VTAIL.n171 VTAIL.n170 9.3005
R1313 VTAIL.n173 VTAIL.n172 9.3005
R1314 VTAIL.n160 VTAIL.n159 9.3005
R1315 VTAIL.n179 VTAIL.n178 9.3005
R1316 VTAIL.n181 VTAIL.n180 9.3005
R1317 VTAIL.n182 VTAIL.n155 9.3005
R1318 VTAIL.n189 VTAIL.n188 9.3005
R1319 VTAIL.n47 VTAIL.n46 9.3005
R1320 VTAIL.n2 VTAIL.n1 9.3005
R1321 VTAIL.n41 VTAIL.n40 9.3005
R1322 VTAIL.n14 VTAIL.n13 9.3005
R1323 VTAIL.n21 VTAIL.n20 9.3005
R1324 VTAIL.n23 VTAIL.n22 9.3005
R1325 VTAIL.n10 VTAIL.n9 9.3005
R1326 VTAIL.n29 VTAIL.n28 9.3005
R1327 VTAIL.n31 VTAIL.n30 9.3005
R1328 VTAIL.n32 VTAIL.n5 9.3005
R1329 VTAIL.n39 VTAIL.n38 9.3005
R1330 VTAIL.n116 VTAIL.n115 9.3005
R1331 VTAIL.n123 VTAIL.n122 9.3005
R1332 VTAIL.n125 VTAIL.n124 9.3005
R1333 VTAIL.n112 VTAIL.n111 9.3005
R1334 VTAIL.n131 VTAIL.n130 9.3005
R1335 VTAIL.n133 VTAIL.n132 9.3005
R1336 VTAIL.n107 VTAIL.n105 9.3005
R1337 VTAIL.n139 VTAIL.n138 9.3005
R1338 VTAIL.n147 VTAIL.n146 9.3005
R1339 VTAIL.n102 VTAIL.n101 9.3005
R1340 VTAIL.n141 VTAIL.n140 9.3005
R1341 VTAIL.n66 VTAIL.n65 9.3005
R1342 VTAIL.n73 VTAIL.n72 9.3005
R1343 VTAIL.n75 VTAIL.n74 9.3005
R1344 VTAIL.n62 VTAIL.n61 9.3005
R1345 VTAIL.n81 VTAIL.n80 9.3005
R1346 VTAIL.n83 VTAIL.n82 9.3005
R1347 VTAIL.n57 VTAIL.n55 9.3005
R1348 VTAIL.n89 VTAIL.n88 9.3005
R1349 VTAIL.n97 VTAIL.n96 9.3005
R1350 VTAIL.n52 VTAIL.n51 9.3005
R1351 VTAIL.n91 VTAIL.n90 9.3005
R1352 VTAIL.n173 VTAIL.n162 8.92171
R1353 VTAIL.n23 VTAIL.n12 8.92171
R1354 VTAIL.n125 VTAIL.n114 8.92171
R1355 VTAIL.n75 VTAIL.n64 8.92171
R1356 VTAIL.n170 VTAIL.n169 8.14595
R1357 VTAIL.n20 VTAIL.n19 8.14595
R1358 VTAIL.n122 VTAIL.n121 8.14595
R1359 VTAIL.n72 VTAIL.n71 8.14595
R1360 VTAIL.n166 VTAIL.n164 7.3702
R1361 VTAIL.n16 VTAIL.n14 7.3702
R1362 VTAIL.n118 VTAIL.n116 7.3702
R1363 VTAIL.n68 VTAIL.n66 7.3702
R1364 VTAIL.n169 VTAIL.n164 5.81868
R1365 VTAIL.n19 VTAIL.n14 5.81868
R1366 VTAIL.n121 VTAIL.n116 5.81868
R1367 VTAIL.n71 VTAIL.n66 5.81868
R1368 VTAIL.n170 VTAIL.n162 5.04292
R1369 VTAIL.n20 VTAIL.n12 5.04292
R1370 VTAIL.n122 VTAIL.n114 5.04292
R1371 VTAIL.n72 VTAIL.n64 5.04292
R1372 VTAIL.n174 VTAIL.n173 4.26717
R1373 VTAIL.n24 VTAIL.n23 4.26717
R1374 VTAIL.n126 VTAIL.n125 4.26717
R1375 VTAIL.n76 VTAIL.n75 4.26717
R1376 VTAIL.n177 VTAIL.n160 3.49141
R1377 VTAIL.n27 VTAIL.n10 3.49141
R1378 VTAIL.n129 VTAIL.n112 3.49141
R1379 VTAIL.n79 VTAIL.n62 3.49141
R1380 VTAIL.n165 VTAIL.n163 2.84303
R1381 VTAIL.n15 VTAIL.n13 2.84303
R1382 VTAIL.n117 VTAIL.n115 2.84303
R1383 VTAIL.n67 VTAIL.n65 2.84303
R1384 VTAIL.n178 VTAIL.n158 2.71565
R1385 VTAIL.n198 VTAIL.n150 2.71565
R1386 VTAIL.n28 VTAIL.n8 2.71565
R1387 VTAIL.n48 VTAIL.n0 2.71565
R1388 VTAIL.n148 VTAIL.n100 2.71565
R1389 VTAIL.n130 VTAIL.n110 2.71565
R1390 VTAIL.n98 VTAIL.n50 2.71565
R1391 VTAIL.n80 VTAIL.n60 2.71565
R1392 VTAIL.n183 VTAIL.n181 1.93989
R1393 VTAIL.n196 VTAIL.n195 1.93989
R1394 VTAIL.n33 VTAIL.n31 1.93989
R1395 VTAIL.n46 VTAIL.n45 1.93989
R1396 VTAIL.n146 VTAIL.n145 1.93989
R1397 VTAIL.n134 VTAIL.n133 1.93989
R1398 VTAIL.n96 VTAIL.n95 1.93989
R1399 VTAIL.n84 VTAIL.n83 1.93989
R1400 VTAIL.n149 VTAIL.n99 1.93584
R1401 VTAIL VTAIL.n49 1.26128
R1402 VTAIL.n182 VTAIL.n156 1.16414
R1403 VTAIL.n192 VTAIL.n152 1.16414
R1404 VTAIL.n32 VTAIL.n6 1.16414
R1405 VTAIL.n42 VTAIL.n2 1.16414
R1406 VTAIL.n142 VTAIL.n102 1.16414
R1407 VTAIL.n137 VTAIL.n107 1.16414
R1408 VTAIL.n92 VTAIL.n52 1.16414
R1409 VTAIL.n87 VTAIL.n57 1.16414
R1410 VTAIL VTAIL.n199 0.675069
R1411 VTAIL.n188 VTAIL.n187 0.388379
R1412 VTAIL.n191 VTAIL.n154 0.388379
R1413 VTAIL.n38 VTAIL.n37 0.388379
R1414 VTAIL.n41 VTAIL.n4 0.388379
R1415 VTAIL.n141 VTAIL.n104 0.388379
R1416 VTAIL.n138 VTAIL.n106 0.388379
R1417 VTAIL.n91 VTAIL.n54 0.388379
R1418 VTAIL.n88 VTAIL.n56 0.388379
R1419 VTAIL.n171 VTAIL.n163 0.155672
R1420 VTAIL.n172 VTAIL.n171 0.155672
R1421 VTAIL.n172 VTAIL.n159 0.155672
R1422 VTAIL.n179 VTAIL.n159 0.155672
R1423 VTAIL.n180 VTAIL.n179 0.155672
R1424 VTAIL.n180 VTAIL.n155 0.155672
R1425 VTAIL.n189 VTAIL.n155 0.155672
R1426 VTAIL.n190 VTAIL.n189 0.155672
R1427 VTAIL.n190 VTAIL.n151 0.155672
R1428 VTAIL.n197 VTAIL.n151 0.155672
R1429 VTAIL.n21 VTAIL.n13 0.155672
R1430 VTAIL.n22 VTAIL.n21 0.155672
R1431 VTAIL.n22 VTAIL.n9 0.155672
R1432 VTAIL.n29 VTAIL.n9 0.155672
R1433 VTAIL.n30 VTAIL.n29 0.155672
R1434 VTAIL.n30 VTAIL.n5 0.155672
R1435 VTAIL.n39 VTAIL.n5 0.155672
R1436 VTAIL.n40 VTAIL.n39 0.155672
R1437 VTAIL.n40 VTAIL.n1 0.155672
R1438 VTAIL.n47 VTAIL.n1 0.155672
R1439 VTAIL.n147 VTAIL.n101 0.155672
R1440 VTAIL.n140 VTAIL.n101 0.155672
R1441 VTAIL.n140 VTAIL.n139 0.155672
R1442 VTAIL.n139 VTAIL.n105 0.155672
R1443 VTAIL.n132 VTAIL.n105 0.155672
R1444 VTAIL.n132 VTAIL.n131 0.155672
R1445 VTAIL.n131 VTAIL.n111 0.155672
R1446 VTAIL.n124 VTAIL.n111 0.155672
R1447 VTAIL.n124 VTAIL.n123 0.155672
R1448 VTAIL.n123 VTAIL.n115 0.155672
R1449 VTAIL.n97 VTAIL.n51 0.155672
R1450 VTAIL.n90 VTAIL.n51 0.155672
R1451 VTAIL.n90 VTAIL.n89 0.155672
R1452 VTAIL.n89 VTAIL.n55 0.155672
R1453 VTAIL.n82 VTAIL.n55 0.155672
R1454 VTAIL.n82 VTAIL.n81 0.155672
R1455 VTAIL.n81 VTAIL.n61 0.155672
R1456 VTAIL.n74 VTAIL.n61 0.155672
R1457 VTAIL.n74 VTAIL.n73 0.155672
R1458 VTAIL.n73 VTAIL.n65 0.155672
R1459 VDD1.n44 VDD1.n0 289.615
R1460 VDD1.n93 VDD1.n49 289.615
R1461 VDD1.n45 VDD1.n44 185
R1462 VDD1.n43 VDD1.n42 185
R1463 VDD1.n4 VDD1.n3 185
R1464 VDD1.n8 VDD1.n6 185
R1465 VDD1.n37 VDD1.n36 185
R1466 VDD1.n35 VDD1.n34 185
R1467 VDD1.n10 VDD1.n9 185
R1468 VDD1.n29 VDD1.n28 185
R1469 VDD1.n27 VDD1.n26 185
R1470 VDD1.n14 VDD1.n13 185
R1471 VDD1.n21 VDD1.n20 185
R1472 VDD1.n19 VDD1.n18 185
R1473 VDD1.n66 VDD1.n65 185
R1474 VDD1.n68 VDD1.n67 185
R1475 VDD1.n61 VDD1.n60 185
R1476 VDD1.n74 VDD1.n73 185
R1477 VDD1.n76 VDD1.n75 185
R1478 VDD1.n57 VDD1.n56 185
R1479 VDD1.n83 VDD1.n82 185
R1480 VDD1.n84 VDD1.n55 185
R1481 VDD1.n86 VDD1.n85 185
R1482 VDD1.n53 VDD1.n52 185
R1483 VDD1.n92 VDD1.n91 185
R1484 VDD1.n94 VDD1.n93 185
R1485 VDD1.n17 VDD1.t1 149.524
R1486 VDD1.n64 VDD1.t0 149.524
R1487 VDD1.n44 VDD1.n43 104.615
R1488 VDD1.n43 VDD1.n3 104.615
R1489 VDD1.n8 VDD1.n3 104.615
R1490 VDD1.n36 VDD1.n8 104.615
R1491 VDD1.n36 VDD1.n35 104.615
R1492 VDD1.n35 VDD1.n9 104.615
R1493 VDD1.n28 VDD1.n9 104.615
R1494 VDD1.n28 VDD1.n27 104.615
R1495 VDD1.n27 VDD1.n13 104.615
R1496 VDD1.n20 VDD1.n13 104.615
R1497 VDD1.n20 VDD1.n19 104.615
R1498 VDD1.n67 VDD1.n66 104.615
R1499 VDD1.n67 VDD1.n60 104.615
R1500 VDD1.n74 VDD1.n60 104.615
R1501 VDD1.n75 VDD1.n74 104.615
R1502 VDD1.n75 VDD1.n56 104.615
R1503 VDD1.n83 VDD1.n56 104.615
R1504 VDD1.n84 VDD1.n83 104.615
R1505 VDD1.n85 VDD1.n84 104.615
R1506 VDD1.n85 VDD1.n52 104.615
R1507 VDD1.n92 VDD1.n52 104.615
R1508 VDD1.n93 VDD1.n92 104.615
R1509 VDD1 VDD1.n97 86.7985
R1510 VDD1.n19 VDD1.t1 52.3082
R1511 VDD1.n66 VDD1.t0 52.3082
R1512 VDD1 VDD1.n48 48.8793
R1513 VDD1.n6 VDD1.n4 13.1884
R1514 VDD1.n86 VDD1.n53 13.1884
R1515 VDD1.n42 VDD1.n41 12.8005
R1516 VDD1.n38 VDD1.n37 12.8005
R1517 VDD1.n87 VDD1.n55 12.8005
R1518 VDD1.n91 VDD1.n90 12.8005
R1519 VDD1.n45 VDD1.n2 12.0247
R1520 VDD1.n34 VDD1.n7 12.0247
R1521 VDD1.n82 VDD1.n81 12.0247
R1522 VDD1.n94 VDD1.n51 12.0247
R1523 VDD1.n46 VDD1.n0 11.249
R1524 VDD1.n33 VDD1.n10 11.249
R1525 VDD1.n80 VDD1.n57 11.249
R1526 VDD1.n95 VDD1.n49 11.249
R1527 VDD1.n30 VDD1.n29 10.4732
R1528 VDD1.n77 VDD1.n76 10.4732
R1529 VDD1.n18 VDD1.n17 10.2747
R1530 VDD1.n65 VDD1.n64 10.2747
R1531 VDD1.n26 VDD1.n12 9.69747
R1532 VDD1.n73 VDD1.n59 9.69747
R1533 VDD1.n48 VDD1.n47 9.45567
R1534 VDD1.n97 VDD1.n96 9.45567
R1535 VDD1.n16 VDD1.n15 9.3005
R1536 VDD1.n23 VDD1.n22 9.3005
R1537 VDD1.n25 VDD1.n24 9.3005
R1538 VDD1.n12 VDD1.n11 9.3005
R1539 VDD1.n31 VDD1.n30 9.3005
R1540 VDD1.n33 VDD1.n32 9.3005
R1541 VDD1.n7 VDD1.n5 9.3005
R1542 VDD1.n39 VDD1.n38 9.3005
R1543 VDD1.n47 VDD1.n46 9.3005
R1544 VDD1.n2 VDD1.n1 9.3005
R1545 VDD1.n41 VDD1.n40 9.3005
R1546 VDD1.n96 VDD1.n95 9.3005
R1547 VDD1.n51 VDD1.n50 9.3005
R1548 VDD1.n90 VDD1.n89 9.3005
R1549 VDD1.n63 VDD1.n62 9.3005
R1550 VDD1.n70 VDD1.n69 9.3005
R1551 VDD1.n72 VDD1.n71 9.3005
R1552 VDD1.n59 VDD1.n58 9.3005
R1553 VDD1.n78 VDD1.n77 9.3005
R1554 VDD1.n80 VDD1.n79 9.3005
R1555 VDD1.n81 VDD1.n54 9.3005
R1556 VDD1.n88 VDD1.n87 9.3005
R1557 VDD1.n25 VDD1.n14 8.92171
R1558 VDD1.n72 VDD1.n61 8.92171
R1559 VDD1.n22 VDD1.n21 8.14595
R1560 VDD1.n69 VDD1.n68 8.14595
R1561 VDD1.n18 VDD1.n16 7.3702
R1562 VDD1.n65 VDD1.n63 7.3702
R1563 VDD1.n21 VDD1.n16 5.81868
R1564 VDD1.n68 VDD1.n63 5.81868
R1565 VDD1.n22 VDD1.n14 5.04292
R1566 VDD1.n69 VDD1.n61 5.04292
R1567 VDD1.n26 VDD1.n25 4.26717
R1568 VDD1.n73 VDD1.n72 4.26717
R1569 VDD1.n29 VDD1.n12 3.49141
R1570 VDD1.n76 VDD1.n59 3.49141
R1571 VDD1.n17 VDD1.n15 2.84303
R1572 VDD1.n64 VDD1.n62 2.84303
R1573 VDD1.n48 VDD1.n0 2.71565
R1574 VDD1.n30 VDD1.n10 2.71565
R1575 VDD1.n77 VDD1.n57 2.71565
R1576 VDD1.n97 VDD1.n49 2.71565
R1577 VDD1.n46 VDD1.n45 1.93989
R1578 VDD1.n34 VDD1.n33 1.93989
R1579 VDD1.n82 VDD1.n80 1.93989
R1580 VDD1.n95 VDD1.n94 1.93989
R1581 VDD1.n42 VDD1.n2 1.16414
R1582 VDD1.n37 VDD1.n7 1.16414
R1583 VDD1.n81 VDD1.n55 1.16414
R1584 VDD1.n91 VDD1.n51 1.16414
R1585 VDD1.n41 VDD1.n4 0.388379
R1586 VDD1.n38 VDD1.n6 0.388379
R1587 VDD1.n87 VDD1.n86 0.388379
R1588 VDD1.n90 VDD1.n53 0.388379
R1589 VDD1.n47 VDD1.n1 0.155672
R1590 VDD1.n40 VDD1.n1 0.155672
R1591 VDD1.n40 VDD1.n39 0.155672
R1592 VDD1.n39 VDD1.n5 0.155672
R1593 VDD1.n32 VDD1.n5 0.155672
R1594 VDD1.n32 VDD1.n31 0.155672
R1595 VDD1.n31 VDD1.n11 0.155672
R1596 VDD1.n24 VDD1.n11 0.155672
R1597 VDD1.n24 VDD1.n23 0.155672
R1598 VDD1.n23 VDD1.n15 0.155672
R1599 VDD1.n70 VDD1.n62 0.155672
R1600 VDD1.n71 VDD1.n70 0.155672
R1601 VDD1.n71 VDD1.n58 0.155672
R1602 VDD1.n78 VDD1.n58 0.155672
R1603 VDD1.n79 VDD1.n78 0.155672
R1604 VDD1.n79 VDD1.n54 0.155672
R1605 VDD1.n88 VDD1.n54 0.155672
R1606 VDD1.n89 VDD1.n88 0.155672
R1607 VDD1.n89 VDD1.n50 0.155672
R1608 VDD1.n96 VDD1.n50 0.155672
R1609 VN VN.t1 157.143
R1610 VN VN.t0 113.791
R1611 VDD2.n93 VDD2.n49 289.615
R1612 VDD2.n44 VDD2.n0 289.615
R1613 VDD2.n94 VDD2.n93 185
R1614 VDD2.n92 VDD2.n91 185
R1615 VDD2.n53 VDD2.n52 185
R1616 VDD2.n57 VDD2.n55 185
R1617 VDD2.n86 VDD2.n85 185
R1618 VDD2.n84 VDD2.n83 185
R1619 VDD2.n59 VDD2.n58 185
R1620 VDD2.n78 VDD2.n77 185
R1621 VDD2.n76 VDD2.n75 185
R1622 VDD2.n63 VDD2.n62 185
R1623 VDD2.n70 VDD2.n69 185
R1624 VDD2.n68 VDD2.n67 185
R1625 VDD2.n17 VDD2.n16 185
R1626 VDD2.n19 VDD2.n18 185
R1627 VDD2.n12 VDD2.n11 185
R1628 VDD2.n25 VDD2.n24 185
R1629 VDD2.n27 VDD2.n26 185
R1630 VDD2.n8 VDD2.n7 185
R1631 VDD2.n34 VDD2.n33 185
R1632 VDD2.n35 VDD2.n6 185
R1633 VDD2.n37 VDD2.n36 185
R1634 VDD2.n4 VDD2.n3 185
R1635 VDD2.n43 VDD2.n42 185
R1636 VDD2.n45 VDD2.n44 185
R1637 VDD2.n66 VDD2.t0 149.524
R1638 VDD2.n15 VDD2.t1 149.524
R1639 VDD2.n93 VDD2.n92 104.615
R1640 VDD2.n92 VDD2.n52 104.615
R1641 VDD2.n57 VDD2.n52 104.615
R1642 VDD2.n85 VDD2.n57 104.615
R1643 VDD2.n85 VDD2.n84 104.615
R1644 VDD2.n84 VDD2.n58 104.615
R1645 VDD2.n77 VDD2.n58 104.615
R1646 VDD2.n77 VDD2.n76 104.615
R1647 VDD2.n76 VDD2.n62 104.615
R1648 VDD2.n69 VDD2.n62 104.615
R1649 VDD2.n69 VDD2.n68 104.615
R1650 VDD2.n18 VDD2.n17 104.615
R1651 VDD2.n18 VDD2.n11 104.615
R1652 VDD2.n25 VDD2.n11 104.615
R1653 VDD2.n26 VDD2.n25 104.615
R1654 VDD2.n26 VDD2.n7 104.615
R1655 VDD2.n34 VDD2.n7 104.615
R1656 VDD2.n35 VDD2.n34 104.615
R1657 VDD2.n36 VDD2.n35 104.615
R1658 VDD2.n36 VDD2.n3 104.615
R1659 VDD2.n43 VDD2.n3 104.615
R1660 VDD2.n44 VDD2.n43 104.615
R1661 VDD2.n98 VDD2.n48 85.5409
R1662 VDD2.n68 VDD2.t0 52.3082
R1663 VDD2.n17 VDD2.t1 52.3082
R1664 VDD2.n98 VDD2.n97 48.0884
R1665 VDD2.n55 VDD2.n53 13.1884
R1666 VDD2.n37 VDD2.n4 13.1884
R1667 VDD2.n91 VDD2.n90 12.8005
R1668 VDD2.n87 VDD2.n86 12.8005
R1669 VDD2.n38 VDD2.n6 12.8005
R1670 VDD2.n42 VDD2.n41 12.8005
R1671 VDD2.n94 VDD2.n51 12.0247
R1672 VDD2.n83 VDD2.n56 12.0247
R1673 VDD2.n33 VDD2.n32 12.0247
R1674 VDD2.n45 VDD2.n2 12.0247
R1675 VDD2.n95 VDD2.n49 11.249
R1676 VDD2.n82 VDD2.n59 11.249
R1677 VDD2.n31 VDD2.n8 11.249
R1678 VDD2.n46 VDD2.n0 11.249
R1679 VDD2.n79 VDD2.n78 10.4732
R1680 VDD2.n28 VDD2.n27 10.4732
R1681 VDD2.n67 VDD2.n66 10.2747
R1682 VDD2.n16 VDD2.n15 10.2747
R1683 VDD2.n75 VDD2.n61 9.69747
R1684 VDD2.n24 VDD2.n10 9.69747
R1685 VDD2.n97 VDD2.n96 9.45567
R1686 VDD2.n48 VDD2.n47 9.45567
R1687 VDD2.n65 VDD2.n64 9.3005
R1688 VDD2.n72 VDD2.n71 9.3005
R1689 VDD2.n74 VDD2.n73 9.3005
R1690 VDD2.n61 VDD2.n60 9.3005
R1691 VDD2.n80 VDD2.n79 9.3005
R1692 VDD2.n82 VDD2.n81 9.3005
R1693 VDD2.n56 VDD2.n54 9.3005
R1694 VDD2.n88 VDD2.n87 9.3005
R1695 VDD2.n96 VDD2.n95 9.3005
R1696 VDD2.n51 VDD2.n50 9.3005
R1697 VDD2.n90 VDD2.n89 9.3005
R1698 VDD2.n47 VDD2.n46 9.3005
R1699 VDD2.n2 VDD2.n1 9.3005
R1700 VDD2.n41 VDD2.n40 9.3005
R1701 VDD2.n14 VDD2.n13 9.3005
R1702 VDD2.n21 VDD2.n20 9.3005
R1703 VDD2.n23 VDD2.n22 9.3005
R1704 VDD2.n10 VDD2.n9 9.3005
R1705 VDD2.n29 VDD2.n28 9.3005
R1706 VDD2.n31 VDD2.n30 9.3005
R1707 VDD2.n32 VDD2.n5 9.3005
R1708 VDD2.n39 VDD2.n38 9.3005
R1709 VDD2.n74 VDD2.n63 8.92171
R1710 VDD2.n23 VDD2.n12 8.92171
R1711 VDD2.n71 VDD2.n70 8.14595
R1712 VDD2.n20 VDD2.n19 8.14595
R1713 VDD2.n67 VDD2.n65 7.3702
R1714 VDD2.n16 VDD2.n14 7.3702
R1715 VDD2.n70 VDD2.n65 5.81868
R1716 VDD2.n19 VDD2.n14 5.81868
R1717 VDD2.n71 VDD2.n63 5.04292
R1718 VDD2.n20 VDD2.n12 5.04292
R1719 VDD2.n75 VDD2.n74 4.26717
R1720 VDD2.n24 VDD2.n23 4.26717
R1721 VDD2.n78 VDD2.n61 3.49141
R1722 VDD2.n27 VDD2.n10 3.49141
R1723 VDD2.n66 VDD2.n64 2.84303
R1724 VDD2.n15 VDD2.n13 2.84303
R1725 VDD2.n97 VDD2.n49 2.71565
R1726 VDD2.n79 VDD2.n59 2.71565
R1727 VDD2.n28 VDD2.n8 2.71565
R1728 VDD2.n48 VDD2.n0 2.71565
R1729 VDD2.n95 VDD2.n94 1.93989
R1730 VDD2.n83 VDD2.n82 1.93989
R1731 VDD2.n33 VDD2.n31 1.93989
R1732 VDD2.n46 VDD2.n45 1.93989
R1733 VDD2.n91 VDD2.n51 1.16414
R1734 VDD2.n86 VDD2.n56 1.16414
R1735 VDD2.n32 VDD2.n6 1.16414
R1736 VDD2.n42 VDD2.n2 1.16414
R1737 VDD2 VDD2.n98 0.791448
R1738 VDD2.n90 VDD2.n53 0.388379
R1739 VDD2.n87 VDD2.n55 0.388379
R1740 VDD2.n38 VDD2.n37 0.388379
R1741 VDD2.n41 VDD2.n4 0.388379
R1742 VDD2.n96 VDD2.n50 0.155672
R1743 VDD2.n89 VDD2.n50 0.155672
R1744 VDD2.n89 VDD2.n88 0.155672
R1745 VDD2.n88 VDD2.n54 0.155672
R1746 VDD2.n81 VDD2.n54 0.155672
R1747 VDD2.n81 VDD2.n80 0.155672
R1748 VDD2.n80 VDD2.n60 0.155672
R1749 VDD2.n73 VDD2.n60 0.155672
R1750 VDD2.n73 VDD2.n72 0.155672
R1751 VDD2.n72 VDD2.n64 0.155672
R1752 VDD2.n21 VDD2.n13 0.155672
R1753 VDD2.n22 VDD2.n21 0.155672
R1754 VDD2.n22 VDD2.n9 0.155672
R1755 VDD2.n29 VDD2.n9 0.155672
R1756 VDD2.n30 VDD2.n29 0.155672
R1757 VDD2.n30 VDD2.n5 0.155672
R1758 VDD2.n39 VDD2.n5 0.155672
R1759 VDD2.n40 VDD2.n39 0.155672
R1760 VDD2.n40 VDD2.n1 0.155672
R1761 VDD2.n47 VDD2.n1 0.155672
C0 VDD2 VP 0.352943f
C1 VN VTAIL 2.07003f
C2 VDD1 VTAIL 4.42729f
C3 VN VDD1 0.148672f
C4 VP VTAIL 2.08425f
C5 VDD2 VTAIL 4.48205f
C6 VN VP 5.15177f
C7 VP VDD1 2.44308f
C8 VN VDD2 2.24071f
C9 VDD2 VDD1 0.731424f
C10 VDD2 B 4.093293f
C11 VDD1 B 6.691521f
C12 VTAIL B 6.451639f
C13 VN B 10.52514f
C14 VP B 6.789185f
C15 VDD2.n0 B 0.026117f
C16 VDD2.n1 B 0.020554f
C17 VDD2.n2 B 0.011045f
C18 VDD2.n3 B 0.026105f
C19 VDD2.n4 B 0.01137f
C20 VDD2.n5 B 0.020554f
C21 VDD2.n6 B 0.011694f
C22 VDD2.n7 B 0.026105f
C23 VDD2.n8 B 0.011694f
C24 VDD2.n9 B 0.020554f
C25 VDD2.n10 B 0.011045f
C26 VDD2.n11 B 0.026105f
C27 VDD2.n12 B 0.011694f
C28 VDD2.n13 B 0.780914f
C29 VDD2.n14 B 0.011045f
C30 VDD2.t1 B 0.043783f
C31 VDD2.n15 B 0.126099f
C32 VDD2.n16 B 0.018455f
C33 VDD2.n17 B 0.019579f
C34 VDD2.n18 B 0.026105f
C35 VDD2.n19 B 0.011694f
C36 VDD2.n20 B 0.011045f
C37 VDD2.n21 B 0.020554f
C38 VDD2.n22 B 0.020554f
C39 VDD2.n23 B 0.011045f
C40 VDD2.n24 B 0.011694f
C41 VDD2.n25 B 0.026105f
C42 VDD2.n26 B 0.026105f
C43 VDD2.n27 B 0.011694f
C44 VDD2.n28 B 0.011045f
C45 VDD2.n29 B 0.020554f
C46 VDD2.n30 B 0.020554f
C47 VDD2.n31 B 0.011045f
C48 VDD2.n32 B 0.011045f
C49 VDD2.n33 B 0.011694f
C50 VDD2.n34 B 0.026105f
C51 VDD2.n35 B 0.026105f
C52 VDD2.n36 B 0.026105f
C53 VDD2.n37 B 0.01137f
C54 VDD2.n38 B 0.011045f
C55 VDD2.n39 B 0.020554f
C56 VDD2.n40 B 0.020554f
C57 VDD2.n41 B 0.011045f
C58 VDD2.n42 B 0.011694f
C59 VDD2.n43 B 0.026105f
C60 VDD2.n44 B 0.051609f
C61 VDD2.n45 B 0.011694f
C62 VDD2.n46 B 0.011045f
C63 VDD2.n47 B 0.046386f
C64 VDD2.n48 B 0.550233f
C65 VDD2.n49 B 0.026117f
C66 VDD2.n50 B 0.020554f
C67 VDD2.n51 B 0.011045f
C68 VDD2.n52 B 0.026105f
C69 VDD2.n53 B 0.01137f
C70 VDD2.n54 B 0.020554f
C71 VDD2.n55 B 0.01137f
C72 VDD2.n56 B 0.011045f
C73 VDD2.n57 B 0.026105f
C74 VDD2.n58 B 0.026105f
C75 VDD2.n59 B 0.011694f
C76 VDD2.n60 B 0.020554f
C77 VDD2.n61 B 0.011045f
C78 VDD2.n62 B 0.026105f
C79 VDD2.n63 B 0.011694f
C80 VDD2.n64 B 0.780914f
C81 VDD2.n65 B 0.011045f
C82 VDD2.t0 B 0.043783f
C83 VDD2.n66 B 0.126099f
C84 VDD2.n67 B 0.018455f
C85 VDD2.n68 B 0.019579f
C86 VDD2.n69 B 0.026105f
C87 VDD2.n70 B 0.011694f
C88 VDD2.n71 B 0.011045f
C89 VDD2.n72 B 0.020554f
C90 VDD2.n73 B 0.020554f
C91 VDD2.n74 B 0.011045f
C92 VDD2.n75 B 0.011694f
C93 VDD2.n76 B 0.026105f
C94 VDD2.n77 B 0.026105f
C95 VDD2.n78 B 0.011694f
C96 VDD2.n79 B 0.011045f
C97 VDD2.n80 B 0.020554f
C98 VDD2.n81 B 0.020554f
C99 VDD2.n82 B 0.011045f
C100 VDD2.n83 B 0.011694f
C101 VDD2.n84 B 0.026105f
C102 VDD2.n85 B 0.026105f
C103 VDD2.n86 B 0.011694f
C104 VDD2.n87 B 0.011045f
C105 VDD2.n88 B 0.020554f
C106 VDD2.n89 B 0.020554f
C107 VDD2.n90 B 0.011045f
C108 VDD2.n91 B 0.011694f
C109 VDD2.n92 B 0.026105f
C110 VDD2.n93 B 0.051609f
C111 VDD2.n94 B 0.011694f
C112 VDD2.n95 B 0.011045f
C113 VDD2.n96 B 0.046386f
C114 VDD2.n97 B 0.042539f
C115 VDD2.n98 B 2.3403f
C116 VN.t0 B 2.60537f
C117 VN.t1 B 3.19368f
C118 VDD1.n0 B 0.026209f
C119 VDD1.n1 B 0.020627f
C120 VDD1.n2 B 0.011084f
C121 VDD1.n3 B 0.026198f
C122 VDD1.n4 B 0.01141f
C123 VDD1.n5 B 0.020627f
C124 VDD1.n6 B 0.01141f
C125 VDD1.n7 B 0.011084f
C126 VDD1.n8 B 0.026198f
C127 VDD1.n9 B 0.026198f
C128 VDD1.n10 B 0.011736f
C129 VDD1.n11 B 0.020627f
C130 VDD1.n12 B 0.011084f
C131 VDD1.n13 B 0.026198f
C132 VDD1.n14 B 0.011736f
C133 VDD1.n15 B 0.78369f
C134 VDD1.n16 B 0.011084f
C135 VDD1.t1 B 0.043939f
C136 VDD1.n17 B 0.126547f
C137 VDD1.n18 B 0.01852f
C138 VDD1.n19 B 0.019649f
C139 VDD1.n20 B 0.026198f
C140 VDD1.n21 B 0.011736f
C141 VDD1.n22 B 0.011084f
C142 VDD1.n23 B 0.020627f
C143 VDD1.n24 B 0.020627f
C144 VDD1.n25 B 0.011084f
C145 VDD1.n26 B 0.011736f
C146 VDD1.n27 B 0.026198f
C147 VDD1.n28 B 0.026198f
C148 VDD1.n29 B 0.011736f
C149 VDD1.n30 B 0.011084f
C150 VDD1.n31 B 0.020627f
C151 VDD1.n32 B 0.020627f
C152 VDD1.n33 B 0.011084f
C153 VDD1.n34 B 0.011736f
C154 VDD1.n35 B 0.026198f
C155 VDD1.n36 B 0.026198f
C156 VDD1.n37 B 0.011736f
C157 VDD1.n38 B 0.011084f
C158 VDD1.n39 B 0.020627f
C159 VDD1.n40 B 0.020627f
C160 VDD1.n41 B 0.011084f
C161 VDD1.n42 B 0.011736f
C162 VDD1.n43 B 0.026198f
C163 VDD1.n44 B 0.051793f
C164 VDD1.n45 B 0.011736f
C165 VDD1.n46 B 0.011084f
C166 VDD1.n47 B 0.04655f
C167 VDD1.n48 B 0.044174f
C168 VDD1.n49 B 0.026209f
C169 VDD1.n50 B 0.020627f
C170 VDD1.n51 B 0.011084f
C171 VDD1.n52 B 0.026198f
C172 VDD1.n53 B 0.01141f
C173 VDD1.n54 B 0.020627f
C174 VDD1.n55 B 0.011736f
C175 VDD1.n56 B 0.026198f
C176 VDD1.n57 B 0.011736f
C177 VDD1.n58 B 0.020627f
C178 VDD1.n59 B 0.011084f
C179 VDD1.n60 B 0.026198f
C180 VDD1.n61 B 0.011736f
C181 VDD1.n62 B 0.78369f
C182 VDD1.n63 B 0.011084f
C183 VDD1.t0 B 0.043939f
C184 VDD1.n64 B 0.126547f
C185 VDD1.n65 B 0.01852f
C186 VDD1.n66 B 0.019649f
C187 VDD1.n67 B 0.026198f
C188 VDD1.n68 B 0.011736f
C189 VDD1.n69 B 0.011084f
C190 VDD1.n70 B 0.020627f
C191 VDD1.n71 B 0.020627f
C192 VDD1.n72 B 0.011084f
C193 VDD1.n73 B 0.011736f
C194 VDD1.n74 B 0.026198f
C195 VDD1.n75 B 0.026198f
C196 VDD1.n76 B 0.011736f
C197 VDD1.n77 B 0.011084f
C198 VDD1.n78 B 0.020627f
C199 VDD1.n79 B 0.020627f
C200 VDD1.n80 B 0.011084f
C201 VDD1.n81 B 0.011084f
C202 VDD1.n82 B 0.011736f
C203 VDD1.n83 B 0.026198f
C204 VDD1.n84 B 0.026198f
C205 VDD1.n85 B 0.026198f
C206 VDD1.n86 B 0.01141f
C207 VDD1.n87 B 0.011084f
C208 VDD1.n88 B 0.020627f
C209 VDD1.n89 B 0.020627f
C210 VDD1.n90 B 0.011084f
C211 VDD1.n91 B 0.011736f
C212 VDD1.n92 B 0.026198f
C213 VDD1.n93 B 0.051793f
C214 VDD1.n94 B 0.011736f
C215 VDD1.n95 B 0.011084f
C216 VDD1.n96 B 0.04655f
C217 VDD1.n97 B 0.594236f
C218 VTAIL.n0 B 0.027792f
C219 VTAIL.n1 B 0.021872f
C220 VTAIL.n2 B 0.011753f
C221 VTAIL.n3 B 0.027781f
C222 VTAIL.n4 B 0.012099f
C223 VTAIL.n5 B 0.021872f
C224 VTAIL.n6 B 0.012445f
C225 VTAIL.n7 B 0.027781f
C226 VTAIL.n8 B 0.012445f
C227 VTAIL.n9 B 0.021872f
C228 VTAIL.n10 B 0.011753f
C229 VTAIL.n11 B 0.027781f
C230 VTAIL.n12 B 0.012445f
C231 VTAIL.n13 B 0.831022f
C232 VTAIL.n14 B 0.011753f
C233 VTAIL.t2 B 0.046592f
C234 VTAIL.n15 B 0.13419f
C235 VTAIL.n16 B 0.019639f
C236 VTAIL.n17 B 0.020836f
C237 VTAIL.n18 B 0.027781f
C238 VTAIL.n19 B 0.012445f
C239 VTAIL.n20 B 0.011753f
C240 VTAIL.n21 B 0.021872f
C241 VTAIL.n22 B 0.021872f
C242 VTAIL.n23 B 0.011753f
C243 VTAIL.n24 B 0.012445f
C244 VTAIL.n25 B 0.027781f
C245 VTAIL.n26 B 0.027781f
C246 VTAIL.n27 B 0.012445f
C247 VTAIL.n28 B 0.011753f
C248 VTAIL.n29 B 0.021872f
C249 VTAIL.n30 B 0.021872f
C250 VTAIL.n31 B 0.011753f
C251 VTAIL.n32 B 0.011753f
C252 VTAIL.n33 B 0.012445f
C253 VTAIL.n34 B 0.027781f
C254 VTAIL.n35 B 0.027781f
C255 VTAIL.n36 B 0.027781f
C256 VTAIL.n37 B 0.012099f
C257 VTAIL.n38 B 0.011753f
C258 VTAIL.n39 B 0.021872f
C259 VTAIL.n40 B 0.021872f
C260 VTAIL.n41 B 0.011753f
C261 VTAIL.n42 B 0.012445f
C262 VTAIL.n43 B 0.027781f
C263 VTAIL.n44 B 0.054921f
C264 VTAIL.n45 B 0.012445f
C265 VTAIL.n46 B 0.011753f
C266 VTAIL.n47 B 0.049362f
C267 VTAIL.n48 B 0.030157f
C268 VTAIL.n49 B 1.37609f
C269 VTAIL.n50 B 0.027792f
C270 VTAIL.n51 B 0.021872f
C271 VTAIL.n52 B 0.011753f
C272 VTAIL.n53 B 0.027781f
C273 VTAIL.n54 B 0.012099f
C274 VTAIL.n55 B 0.021872f
C275 VTAIL.n56 B 0.012099f
C276 VTAIL.n57 B 0.011753f
C277 VTAIL.n58 B 0.027781f
C278 VTAIL.n59 B 0.027781f
C279 VTAIL.n60 B 0.012445f
C280 VTAIL.n61 B 0.021872f
C281 VTAIL.n62 B 0.011753f
C282 VTAIL.n63 B 0.027781f
C283 VTAIL.n64 B 0.012445f
C284 VTAIL.n65 B 0.831022f
C285 VTAIL.n66 B 0.011753f
C286 VTAIL.t0 B 0.046592f
C287 VTAIL.n67 B 0.13419f
C288 VTAIL.n68 B 0.019639f
C289 VTAIL.n69 B 0.020836f
C290 VTAIL.n70 B 0.027781f
C291 VTAIL.n71 B 0.012445f
C292 VTAIL.n72 B 0.011753f
C293 VTAIL.n73 B 0.021872f
C294 VTAIL.n74 B 0.021872f
C295 VTAIL.n75 B 0.011753f
C296 VTAIL.n76 B 0.012445f
C297 VTAIL.n77 B 0.027781f
C298 VTAIL.n78 B 0.027781f
C299 VTAIL.n79 B 0.012445f
C300 VTAIL.n80 B 0.011753f
C301 VTAIL.n81 B 0.021872f
C302 VTAIL.n82 B 0.021872f
C303 VTAIL.n83 B 0.011753f
C304 VTAIL.n84 B 0.012445f
C305 VTAIL.n85 B 0.027781f
C306 VTAIL.n86 B 0.027781f
C307 VTAIL.n87 B 0.012445f
C308 VTAIL.n88 B 0.011753f
C309 VTAIL.n89 B 0.021872f
C310 VTAIL.n90 B 0.021872f
C311 VTAIL.n91 B 0.011753f
C312 VTAIL.n92 B 0.012445f
C313 VTAIL.n93 B 0.027781f
C314 VTAIL.n94 B 0.054921f
C315 VTAIL.n95 B 0.012445f
C316 VTAIL.n96 B 0.011753f
C317 VTAIL.n97 B 0.049362f
C318 VTAIL.n98 B 0.030157f
C319 VTAIL.n99 B 1.42363f
C320 VTAIL.n100 B 0.027792f
C321 VTAIL.n101 B 0.021872f
C322 VTAIL.n102 B 0.011753f
C323 VTAIL.n103 B 0.027781f
C324 VTAIL.n104 B 0.012099f
C325 VTAIL.n105 B 0.021872f
C326 VTAIL.n106 B 0.012099f
C327 VTAIL.n107 B 0.011753f
C328 VTAIL.n108 B 0.027781f
C329 VTAIL.n109 B 0.027781f
C330 VTAIL.n110 B 0.012445f
C331 VTAIL.n111 B 0.021872f
C332 VTAIL.n112 B 0.011753f
C333 VTAIL.n113 B 0.027781f
C334 VTAIL.n114 B 0.012445f
C335 VTAIL.n115 B 0.831022f
C336 VTAIL.n116 B 0.011753f
C337 VTAIL.t3 B 0.046592f
C338 VTAIL.n117 B 0.13419f
C339 VTAIL.n118 B 0.019639f
C340 VTAIL.n119 B 0.020836f
C341 VTAIL.n120 B 0.027781f
C342 VTAIL.n121 B 0.012445f
C343 VTAIL.n122 B 0.011753f
C344 VTAIL.n123 B 0.021872f
C345 VTAIL.n124 B 0.021872f
C346 VTAIL.n125 B 0.011753f
C347 VTAIL.n126 B 0.012445f
C348 VTAIL.n127 B 0.027781f
C349 VTAIL.n128 B 0.027781f
C350 VTAIL.n129 B 0.012445f
C351 VTAIL.n130 B 0.011753f
C352 VTAIL.n131 B 0.021872f
C353 VTAIL.n132 B 0.021872f
C354 VTAIL.n133 B 0.011753f
C355 VTAIL.n134 B 0.012445f
C356 VTAIL.n135 B 0.027781f
C357 VTAIL.n136 B 0.027781f
C358 VTAIL.n137 B 0.012445f
C359 VTAIL.n138 B 0.011753f
C360 VTAIL.n139 B 0.021872f
C361 VTAIL.n140 B 0.021872f
C362 VTAIL.n141 B 0.011753f
C363 VTAIL.n142 B 0.012445f
C364 VTAIL.n143 B 0.027781f
C365 VTAIL.n144 B 0.054921f
C366 VTAIL.n145 B 0.012445f
C367 VTAIL.n146 B 0.011753f
C368 VTAIL.n147 B 0.049362f
C369 VTAIL.n148 B 0.030157f
C370 VTAIL.n149 B 1.21706f
C371 VTAIL.n150 B 0.027792f
C372 VTAIL.n151 B 0.021872f
C373 VTAIL.n152 B 0.011753f
C374 VTAIL.n153 B 0.027781f
C375 VTAIL.n154 B 0.012099f
C376 VTAIL.n155 B 0.021872f
C377 VTAIL.n156 B 0.012445f
C378 VTAIL.n157 B 0.027781f
C379 VTAIL.n158 B 0.012445f
C380 VTAIL.n159 B 0.021872f
C381 VTAIL.n160 B 0.011753f
C382 VTAIL.n161 B 0.027781f
C383 VTAIL.n162 B 0.012445f
C384 VTAIL.n163 B 0.831022f
C385 VTAIL.n164 B 0.011753f
C386 VTAIL.t1 B 0.046592f
C387 VTAIL.n165 B 0.13419f
C388 VTAIL.n166 B 0.019639f
C389 VTAIL.n167 B 0.020836f
C390 VTAIL.n168 B 0.027781f
C391 VTAIL.n169 B 0.012445f
C392 VTAIL.n170 B 0.011753f
C393 VTAIL.n171 B 0.021872f
C394 VTAIL.n172 B 0.021872f
C395 VTAIL.n173 B 0.011753f
C396 VTAIL.n174 B 0.012445f
C397 VTAIL.n175 B 0.027781f
C398 VTAIL.n176 B 0.027781f
C399 VTAIL.n177 B 0.012445f
C400 VTAIL.n178 B 0.011753f
C401 VTAIL.n179 B 0.021872f
C402 VTAIL.n180 B 0.021872f
C403 VTAIL.n181 B 0.011753f
C404 VTAIL.n182 B 0.011753f
C405 VTAIL.n183 B 0.012445f
C406 VTAIL.n184 B 0.027781f
C407 VTAIL.n185 B 0.027781f
C408 VTAIL.n186 B 0.027781f
C409 VTAIL.n187 B 0.012099f
C410 VTAIL.n188 B 0.011753f
C411 VTAIL.n189 B 0.021872f
C412 VTAIL.n190 B 0.021872f
C413 VTAIL.n191 B 0.011753f
C414 VTAIL.n192 B 0.012445f
C415 VTAIL.n193 B 0.027781f
C416 VTAIL.n194 B 0.054921f
C417 VTAIL.n195 B 0.012445f
C418 VTAIL.n196 B 0.011753f
C419 VTAIL.n197 B 0.049362f
C420 VTAIL.n198 B 0.030157f
C421 VTAIL.n199 B 1.1282f
C422 VP.t1 B 2.66864f
C423 VP.t0 B 3.27296f
C424 VP.n0 B 3.6668f
.ends

