* NGSPICE file created from diff_pair_sample_0613.ext - technology: sky130A

.subckt diff_pair_sample_0613 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t7 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X1 VDD1.t6 VP.t1 VTAIL.t16 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=2.76
X2 VDD2.t9 VN.t0 VTAIL.t2 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=2.76
X3 VDD2.t8 VN.t1 VTAIL.t7 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X4 VDD2.t7 VN.t2 VTAIL.t0 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X5 VTAIL.t15 VP.t2 VDD1.t9 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X6 VTAIL.t14 VP.t3 VDD1.t8 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X7 VDD2.t6 VN.t3 VTAIL.t19 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=2.76
X8 VTAIL.t18 VN.t4 VDD2.t5 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X9 B.t11 B.t9 B.t10 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=2.76
X10 VDD1.t3 VP.t4 VTAIL.t13 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=2.76
X11 B.t8 B.t6 B.t7 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=2.76
X12 VDD2.t4 VN.t5 VTAIL.t6 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=2.76
X13 VTAIL.t4 VN.t6 VDD2.t3 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X14 VTAIL.t3 VN.t7 VDD2.t2 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X15 VDD1.t2 VP.t5 VTAIL.t12 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X16 VTAIL.t5 VN.t8 VDD2.t1 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X17 VDD1.t1 VP.t6 VTAIL.t11 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X18 B.t5 B.t3 B.t4 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=2.76
X19 B.t2 B.t0 B.t1 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=2.76
X20 VTAIL.t10 VP.t7 VDD1.t0 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=2.76
X21 VDD1.t5 VP.t8 VTAIL.t9 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=2.76
X22 VDD2.t0 VN.t9 VTAIL.t1 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=2.76
X23 VDD1.t4 VP.t9 VTAIL.t8 w_n4678_n3398# sky130_fd_pr__pfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=2.76
R0 VP.n25 VP.n22 161.3
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n21 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n20 161.3
R5 VP.n34 VP.n33 161.3
R6 VP.n35 VP.n19 161.3
R7 VP.n37 VP.n36 161.3
R8 VP.n38 VP.n18 161.3
R9 VP.n40 VP.n39 161.3
R10 VP.n41 VP.n17 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n45 VP.n16 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n48 VP.n15 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n51 VP.n14 161.3
R17 VP.n53 VP.n52 161.3
R18 VP.n95 VP.n94 161.3
R19 VP.n93 VP.n1 161.3
R20 VP.n92 VP.n91 161.3
R21 VP.n90 VP.n2 161.3
R22 VP.n89 VP.n88 161.3
R23 VP.n87 VP.n3 161.3
R24 VP.n85 VP.n84 161.3
R25 VP.n83 VP.n4 161.3
R26 VP.n82 VP.n81 161.3
R27 VP.n80 VP.n5 161.3
R28 VP.n79 VP.n78 161.3
R29 VP.n77 VP.n6 161.3
R30 VP.n76 VP.n75 161.3
R31 VP.n73 VP.n7 161.3
R32 VP.n72 VP.n71 161.3
R33 VP.n70 VP.n8 161.3
R34 VP.n69 VP.n68 161.3
R35 VP.n67 VP.n9 161.3
R36 VP.n65 VP.n64 161.3
R37 VP.n63 VP.n10 161.3
R38 VP.n62 VP.n61 161.3
R39 VP.n60 VP.n11 161.3
R40 VP.n59 VP.n58 161.3
R41 VP.n57 VP.n12 161.3
R42 VP.n23 VP.t8 137.976
R43 VP.n55 VP.t1 106.093
R44 VP.n66 VP.t2 106.093
R45 VP.n74 VP.t5 106.093
R46 VP.n86 VP.t0 106.093
R47 VP.n0 VP.t4 106.093
R48 VP.n13 VP.t9 106.093
R49 VP.n44 VP.t7 106.093
R50 VP.n32 VP.t6 106.093
R51 VP.n24 VP.t3 106.093
R52 VP.n56 VP.n55 69.0258
R53 VP.n96 VP.n0 69.0258
R54 VP.n54 VP.n13 69.0258
R55 VP.n24 VP.n23 56.938
R56 VP.n72 VP.n8 56.5193
R57 VP.n81 VP.n80 56.5193
R58 VP.n39 VP.n38 56.5193
R59 VP.n30 VP.n21 56.5193
R60 VP.n56 VP.n54 54.1774
R61 VP.n61 VP.n60 51.663
R62 VP.n92 VP.n2 51.663
R63 VP.n50 VP.n15 51.663
R64 VP.n60 VP.n59 29.3238
R65 VP.n93 VP.n92 29.3238
R66 VP.n51 VP.n50 29.3238
R67 VP.n59 VP.n12 24.4675
R68 VP.n61 VP.n10 24.4675
R69 VP.n65 VP.n10 24.4675
R70 VP.n68 VP.n67 24.4675
R71 VP.n68 VP.n8 24.4675
R72 VP.n73 VP.n72 24.4675
R73 VP.n75 VP.n73 24.4675
R74 VP.n79 VP.n6 24.4675
R75 VP.n80 VP.n79 24.4675
R76 VP.n81 VP.n4 24.4675
R77 VP.n85 VP.n4 24.4675
R78 VP.n88 VP.n87 24.4675
R79 VP.n88 VP.n2 24.4675
R80 VP.n94 VP.n93 24.4675
R81 VP.n52 VP.n51 24.4675
R82 VP.n39 VP.n17 24.4675
R83 VP.n43 VP.n17 24.4675
R84 VP.n46 VP.n45 24.4675
R85 VP.n46 VP.n15 24.4675
R86 VP.n31 VP.n30 24.4675
R87 VP.n33 VP.n31 24.4675
R88 VP.n37 VP.n19 24.4675
R89 VP.n38 VP.n37 24.4675
R90 VP.n26 VP.n25 24.4675
R91 VP.n26 VP.n21 24.4675
R92 VP.n55 VP.n12 21.0421
R93 VP.n94 VP.n0 21.0421
R94 VP.n52 VP.n13 21.0421
R95 VP.n67 VP.n66 16.6381
R96 VP.n86 VP.n85 16.6381
R97 VP.n44 VP.n43 16.6381
R98 VP.n25 VP.n24 16.6381
R99 VP.n75 VP.n74 12.234
R100 VP.n74 VP.n6 12.234
R101 VP.n33 VP.n32 12.234
R102 VP.n32 VP.n19 12.234
R103 VP.n66 VP.n65 7.82994
R104 VP.n87 VP.n86 7.82994
R105 VP.n45 VP.n44 7.82994
R106 VP.n23 VP.n22 5.4582
R107 VP.n54 VP.n53 0.354971
R108 VP.n57 VP.n56 0.354971
R109 VP.n96 VP.n95 0.354971
R110 VP VP.n96 0.26696
R111 VP.n27 VP.n22 0.189894
R112 VP.n28 VP.n27 0.189894
R113 VP.n29 VP.n28 0.189894
R114 VP.n29 VP.n20 0.189894
R115 VP.n34 VP.n20 0.189894
R116 VP.n35 VP.n34 0.189894
R117 VP.n36 VP.n35 0.189894
R118 VP.n36 VP.n18 0.189894
R119 VP.n40 VP.n18 0.189894
R120 VP.n41 VP.n40 0.189894
R121 VP.n42 VP.n41 0.189894
R122 VP.n42 VP.n16 0.189894
R123 VP.n47 VP.n16 0.189894
R124 VP.n48 VP.n47 0.189894
R125 VP.n49 VP.n48 0.189894
R126 VP.n49 VP.n14 0.189894
R127 VP.n53 VP.n14 0.189894
R128 VP.n58 VP.n57 0.189894
R129 VP.n58 VP.n11 0.189894
R130 VP.n62 VP.n11 0.189894
R131 VP.n63 VP.n62 0.189894
R132 VP.n64 VP.n63 0.189894
R133 VP.n64 VP.n9 0.189894
R134 VP.n69 VP.n9 0.189894
R135 VP.n70 VP.n69 0.189894
R136 VP.n71 VP.n70 0.189894
R137 VP.n71 VP.n7 0.189894
R138 VP.n76 VP.n7 0.189894
R139 VP.n77 VP.n76 0.189894
R140 VP.n78 VP.n77 0.189894
R141 VP.n78 VP.n5 0.189894
R142 VP.n82 VP.n5 0.189894
R143 VP.n83 VP.n82 0.189894
R144 VP.n84 VP.n83 0.189894
R145 VP.n84 VP.n3 0.189894
R146 VP.n89 VP.n3 0.189894
R147 VP.n90 VP.n89 0.189894
R148 VP.n91 VP.n90 0.189894
R149 VP.n91 VP.n1 0.189894
R150 VP.n95 VP.n1 0.189894
R151 VDD1.n60 VDD1.n0 756.745
R152 VDD1.n127 VDD1.n67 756.745
R153 VDD1.n61 VDD1.n60 585
R154 VDD1.n59 VDD1.n58 585
R155 VDD1.n4 VDD1.n3 585
R156 VDD1.n53 VDD1.n52 585
R157 VDD1.n51 VDD1.n50 585
R158 VDD1.n8 VDD1.n7 585
R159 VDD1.n45 VDD1.n44 585
R160 VDD1.n43 VDD1.n10 585
R161 VDD1.n42 VDD1.n41 585
R162 VDD1.n13 VDD1.n11 585
R163 VDD1.n36 VDD1.n35 585
R164 VDD1.n34 VDD1.n33 585
R165 VDD1.n17 VDD1.n16 585
R166 VDD1.n28 VDD1.n27 585
R167 VDD1.n26 VDD1.n25 585
R168 VDD1.n21 VDD1.n20 585
R169 VDD1.n87 VDD1.n86 585
R170 VDD1.n92 VDD1.n91 585
R171 VDD1.n94 VDD1.n93 585
R172 VDD1.n83 VDD1.n82 585
R173 VDD1.n100 VDD1.n99 585
R174 VDD1.n102 VDD1.n101 585
R175 VDD1.n79 VDD1.n78 585
R176 VDD1.n109 VDD1.n108 585
R177 VDD1.n110 VDD1.n77 585
R178 VDD1.n112 VDD1.n111 585
R179 VDD1.n75 VDD1.n74 585
R180 VDD1.n118 VDD1.n117 585
R181 VDD1.n120 VDD1.n119 585
R182 VDD1.n71 VDD1.n70 585
R183 VDD1.n126 VDD1.n125 585
R184 VDD1.n128 VDD1.n127 585
R185 VDD1.n22 VDD1.t5 329.036
R186 VDD1.n88 VDD1.t6 329.036
R187 VDD1.n60 VDD1.n59 171.744
R188 VDD1.n59 VDD1.n3 171.744
R189 VDD1.n52 VDD1.n3 171.744
R190 VDD1.n52 VDD1.n51 171.744
R191 VDD1.n51 VDD1.n7 171.744
R192 VDD1.n44 VDD1.n7 171.744
R193 VDD1.n44 VDD1.n43 171.744
R194 VDD1.n43 VDD1.n42 171.744
R195 VDD1.n42 VDD1.n11 171.744
R196 VDD1.n35 VDD1.n11 171.744
R197 VDD1.n35 VDD1.n34 171.744
R198 VDD1.n34 VDD1.n16 171.744
R199 VDD1.n27 VDD1.n16 171.744
R200 VDD1.n27 VDD1.n26 171.744
R201 VDD1.n26 VDD1.n20 171.744
R202 VDD1.n92 VDD1.n86 171.744
R203 VDD1.n93 VDD1.n92 171.744
R204 VDD1.n93 VDD1.n82 171.744
R205 VDD1.n100 VDD1.n82 171.744
R206 VDD1.n101 VDD1.n100 171.744
R207 VDD1.n101 VDD1.n78 171.744
R208 VDD1.n109 VDD1.n78 171.744
R209 VDD1.n110 VDD1.n109 171.744
R210 VDD1.n111 VDD1.n110 171.744
R211 VDD1.n111 VDD1.n74 171.744
R212 VDD1.n118 VDD1.n74 171.744
R213 VDD1.n119 VDD1.n118 171.744
R214 VDD1.n119 VDD1.n70 171.744
R215 VDD1.n126 VDD1.n70 171.744
R216 VDD1.n127 VDD1.n126 171.744
R217 VDD1.t5 VDD1.n20 85.8723
R218 VDD1.t6 VDD1.n86 85.8723
R219 VDD1.n135 VDD1.n134 76.3633
R220 VDD1.n66 VDD1.n65 74.421
R221 VDD1.n137 VDD1.n136 74.4208
R222 VDD1.n133 VDD1.n132 74.4208
R223 VDD1.n66 VDD1.n64 52.1097
R224 VDD1.n133 VDD1.n131 52.1097
R225 VDD1.n137 VDD1.n135 48.7574
R226 VDD1.n45 VDD1.n10 13.1884
R227 VDD1.n112 VDD1.n77 13.1884
R228 VDD1.n46 VDD1.n8 12.8005
R229 VDD1.n41 VDD1.n12 12.8005
R230 VDD1.n108 VDD1.n107 12.8005
R231 VDD1.n113 VDD1.n75 12.8005
R232 VDD1.n50 VDD1.n49 12.0247
R233 VDD1.n40 VDD1.n13 12.0247
R234 VDD1.n106 VDD1.n79 12.0247
R235 VDD1.n117 VDD1.n116 12.0247
R236 VDD1.n53 VDD1.n6 11.249
R237 VDD1.n37 VDD1.n36 11.249
R238 VDD1.n103 VDD1.n102 11.249
R239 VDD1.n120 VDD1.n73 11.249
R240 VDD1.n22 VDD1.n21 10.7239
R241 VDD1.n88 VDD1.n87 10.7239
R242 VDD1.n54 VDD1.n4 10.4732
R243 VDD1.n33 VDD1.n15 10.4732
R244 VDD1.n99 VDD1.n81 10.4732
R245 VDD1.n121 VDD1.n71 10.4732
R246 VDD1.n58 VDD1.n57 9.69747
R247 VDD1.n32 VDD1.n17 9.69747
R248 VDD1.n98 VDD1.n83 9.69747
R249 VDD1.n125 VDD1.n124 9.69747
R250 VDD1.n64 VDD1.n63 9.45567
R251 VDD1.n131 VDD1.n130 9.45567
R252 VDD1.n24 VDD1.n23 9.3005
R253 VDD1.n19 VDD1.n18 9.3005
R254 VDD1.n30 VDD1.n29 9.3005
R255 VDD1.n32 VDD1.n31 9.3005
R256 VDD1.n15 VDD1.n14 9.3005
R257 VDD1.n38 VDD1.n37 9.3005
R258 VDD1.n40 VDD1.n39 9.3005
R259 VDD1.n12 VDD1.n9 9.3005
R260 VDD1.n63 VDD1.n62 9.3005
R261 VDD1.n2 VDD1.n1 9.3005
R262 VDD1.n57 VDD1.n56 9.3005
R263 VDD1.n55 VDD1.n54 9.3005
R264 VDD1.n6 VDD1.n5 9.3005
R265 VDD1.n49 VDD1.n48 9.3005
R266 VDD1.n47 VDD1.n46 9.3005
R267 VDD1.n130 VDD1.n129 9.3005
R268 VDD1.n69 VDD1.n68 9.3005
R269 VDD1.n124 VDD1.n123 9.3005
R270 VDD1.n122 VDD1.n121 9.3005
R271 VDD1.n73 VDD1.n72 9.3005
R272 VDD1.n116 VDD1.n115 9.3005
R273 VDD1.n114 VDD1.n113 9.3005
R274 VDD1.n90 VDD1.n89 9.3005
R275 VDD1.n85 VDD1.n84 9.3005
R276 VDD1.n96 VDD1.n95 9.3005
R277 VDD1.n98 VDD1.n97 9.3005
R278 VDD1.n81 VDD1.n80 9.3005
R279 VDD1.n104 VDD1.n103 9.3005
R280 VDD1.n106 VDD1.n105 9.3005
R281 VDD1.n107 VDD1.n76 9.3005
R282 VDD1.n61 VDD1.n2 8.92171
R283 VDD1.n29 VDD1.n28 8.92171
R284 VDD1.n95 VDD1.n94 8.92171
R285 VDD1.n128 VDD1.n69 8.92171
R286 VDD1.n62 VDD1.n0 8.14595
R287 VDD1.n25 VDD1.n19 8.14595
R288 VDD1.n91 VDD1.n85 8.14595
R289 VDD1.n129 VDD1.n67 8.14595
R290 VDD1.n24 VDD1.n21 7.3702
R291 VDD1.n90 VDD1.n87 7.3702
R292 VDD1.n64 VDD1.n0 5.81868
R293 VDD1.n25 VDD1.n24 5.81868
R294 VDD1.n91 VDD1.n90 5.81868
R295 VDD1.n131 VDD1.n67 5.81868
R296 VDD1.n62 VDD1.n61 5.04292
R297 VDD1.n28 VDD1.n19 5.04292
R298 VDD1.n94 VDD1.n85 5.04292
R299 VDD1.n129 VDD1.n128 5.04292
R300 VDD1.n58 VDD1.n2 4.26717
R301 VDD1.n29 VDD1.n17 4.26717
R302 VDD1.n95 VDD1.n83 4.26717
R303 VDD1.n125 VDD1.n69 4.26717
R304 VDD1.n57 VDD1.n4 3.49141
R305 VDD1.n33 VDD1.n32 3.49141
R306 VDD1.n99 VDD1.n98 3.49141
R307 VDD1.n124 VDD1.n71 3.49141
R308 VDD1.n54 VDD1.n53 2.71565
R309 VDD1.n36 VDD1.n15 2.71565
R310 VDD1.n102 VDD1.n81 2.71565
R311 VDD1.n121 VDD1.n120 2.71565
R312 VDD1.n136 VDD1.t0 2.67581
R313 VDD1.n136 VDD1.t4 2.67581
R314 VDD1.n65 VDD1.t8 2.67581
R315 VDD1.n65 VDD1.t1 2.67581
R316 VDD1.n134 VDD1.t7 2.67581
R317 VDD1.n134 VDD1.t3 2.67581
R318 VDD1.n132 VDD1.t9 2.67581
R319 VDD1.n132 VDD1.t2 2.67581
R320 VDD1.n23 VDD1.n22 2.41282
R321 VDD1.n89 VDD1.n88 2.41282
R322 VDD1 VDD1.n137 1.94016
R323 VDD1.n50 VDD1.n6 1.93989
R324 VDD1.n37 VDD1.n13 1.93989
R325 VDD1.n103 VDD1.n79 1.93989
R326 VDD1.n117 VDD1.n73 1.93989
R327 VDD1.n49 VDD1.n8 1.16414
R328 VDD1.n41 VDD1.n40 1.16414
R329 VDD1.n108 VDD1.n106 1.16414
R330 VDD1.n116 VDD1.n75 1.16414
R331 VDD1 VDD1.n66 0.724638
R332 VDD1.n135 VDD1.n133 0.611102
R333 VDD1.n46 VDD1.n45 0.388379
R334 VDD1.n12 VDD1.n10 0.388379
R335 VDD1.n107 VDD1.n77 0.388379
R336 VDD1.n113 VDD1.n112 0.388379
R337 VDD1.n63 VDD1.n1 0.155672
R338 VDD1.n56 VDD1.n1 0.155672
R339 VDD1.n56 VDD1.n55 0.155672
R340 VDD1.n55 VDD1.n5 0.155672
R341 VDD1.n48 VDD1.n5 0.155672
R342 VDD1.n48 VDD1.n47 0.155672
R343 VDD1.n47 VDD1.n9 0.155672
R344 VDD1.n39 VDD1.n9 0.155672
R345 VDD1.n39 VDD1.n38 0.155672
R346 VDD1.n38 VDD1.n14 0.155672
R347 VDD1.n31 VDD1.n14 0.155672
R348 VDD1.n31 VDD1.n30 0.155672
R349 VDD1.n30 VDD1.n18 0.155672
R350 VDD1.n23 VDD1.n18 0.155672
R351 VDD1.n89 VDD1.n84 0.155672
R352 VDD1.n96 VDD1.n84 0.155672
R353 VDD1.n97 VDD1.n96 0.155672
R354 VDD1.n97 VDD1.n80 0.155672
R355 VDD1.n104 VDD1.n80 0.155672
R356 VDD1.n105 VDD1.n104 0.155672
R357 VDD1.n105 VDD1.n76 0.155672
R358 VDD1.n114 VDD1.n76 0.155672
R359 VDD1.n115 VDD1.n114 0.155672
R360 VDD1.n115 VDD1.n72 0.155672
R361 VDD1.n122 VDD1.n72 0.155672
R362 VDD1.n123 VDD1.n122 0.155672
R363 VDD1.n123 VDD1.n68 0.155672
R364 VDD1.n130 VDD1.n68 0.155672
R365 VTAIL.n272 VTAIL.n212 756.745
R366 VTAIL.n62 VTAIL.n2 756.745
R367 VTAIL.n206 VTAIL.n146 756.745
R368 VTAIL.n136 VTAIL.n76 756.745
R369 VTAIL.n232 VTAIL.n231 585
R370 VTAIL.n237 VTAIL.n236 585
R371 VTAIL.n239 VTAIL.n238 585
R372 VTAIL.n228 VTAIL.n227 585
R373 VTAIL.n245 VTAIL.n244 585
R374 VTAIL.n247 VTAIL.n246 585
R375 VTAIL.n224 VTAIL.n223 585
R376 VTAIL.n254 VTAIL.n253 585
R377 VTAIL.n255 VTAIL.n222 585
R378 VTAIL.n257 VTAIL.n256 585
R379 VTAIL.n220 VTAIL.n219 585
R380 VTAIL.n263 VTAIL.n262 585
R381 VTAIL.n265 VTAIL.n264 585
R382 VTAIL.n216 VTAIL.n215 585
R383 VTAIL.n271 VTAIL.n270 585
R384 VTAIL.n273 VTAIL.n272 585
R385 VTAIL.n22 VTAIL.n21 585
R386 VTAIL.n27 VTAIL.n26 585
R387 VTAIL.n29 VTAIL.n28 585
R388 VTAIL.n18 VTAIL.n17 585
R389 VTAIL.n35 VTAIL.n34 585
R390 VTAIL.n37 VTAIL.n36 585
R391 VTAIL.n14 VTAIL.n13 585
R392 VTAIL.n44 VTAIL.n43 585
R393 VTAIL.n45 VTAIL.n12 585
R394 VTAIL.n47 VTAIL.n46 585
R395 VTAIL.n10 VTAIL.n9 585
R396 VTAIL.n53 VTAIL.n52 585
R397 VTAIL.n55 VTAIL.n54 585
R398 VTAIL.n6 VTAIL.n5 585
R399 VTAIL.n61 VTAIL.n60 585
R400 VTAIL.n63 VTAIL.n62 585
R401 VTAIL.n207 VTAIL.n206 585
R402 VTAIL.n205 VTAIL.n204 585
R403 VTAIL.n150 VTAIL.n149 585
R404 VTAIL.n199 VTAIL.n198 585
R405 VTAIL.n197 VTAIL.n196 585
R406 VTAIL.n154 VTAIL.n153 585
R407 VTAIL.n191 VTAIL.n190 585
R408 VTAIL.n189 VTAIL.n156 585
R409 VTAIL.n188 VTAIL.n187 585
R410 VTAIL.n159 VTAIL.n157 585
R411 VTAIL.n182 VTAIL.n181 585
R412 VTAIL.n180 VTAIL.n179 585
R413 VTAIL.n163 VTAIL.n162 585
R414 VTAIL.n174 VTAIL.n173 585
R415 VTAIL.n172 VTAIL.n171 585
R416 VTAIL.n167 VTAIL.n166 585
R417 VTAIL.n137 VTAIL.n136 585
R418 VTAIL.n135 VTAIL.n134 585
R419 VTAIL.n80 VTAIL.n79 585
R420 VTAIL.n129 VTAIL.n128 585
R421 VTAIL.n127 VTAIL.n126 585
R422 VTAIL.n84 VTAIL.n83 585
R423 VTAIL.n121 VTAIL.n120 585
R424 VTAIL.n119 VTAIL.n86 585
R425 VTAIL.n118 VTAIL.n117 585
R426 VTAIL.n89 VTAIL.n87 585
R427 VTAIL.n112 VTAIL.n111 585
R428 VTAIL.n110 VTAIL.n109 585
R429 VTAIL.n93 VTAIL.n92 585
R430 VTAIL.n104 VTAIL.n103 585
R431 VTAIL.n102 VTAIL.n101 585
R432 VTAIL.n97 VTAIL.n96 585
R433 VTAIL.n233 VTAIL.t2 329.036
R434 VTAIL.n23 VTAIL.t13 329.036
R435 VTAIL.n168 VTAIL.t8 329.036
R436 VTAIL.n98 VTAIL.t19 329.036
R437 VTAIL.n237 VTAIL.n231 171.744
R438 VTAIL.n238 VTAIL.n237 171.744
R439 VTAIL.n238 VTAIL.n227 171.744
R440 VTAIL.n245 VTAIL.n227 171.744
R441 VTAIL.n246 VTAIL.n245 171.744
R442 VTAIL.n246 VTAIL.n223 171.744
R443 VTAIL.n254 VTAIL.n223 171.744
R444 VTAIL.n255 VTAIL.n254 171.744
R445 VTAIL.n256 VTAIL.n255 171.744
R446 VTAIL.n256 VTAIL.n219 171.744
R447 VTAIL.n263 VTAIL.n219 171.744
R448 VTAIL.n264 VTAIL.n263 171.744
R449 VTAIL.n264 VTAIL.n215 171.744
R450 VTAIL.n271 VTAIL.n215 171.744
R451 VTAIL.n272 VTAIL.n271 171.744
R452 VTAIL.n27 VTAIL.n21 171.744
R453 VTAIL.n28 VTAIL.n27 171.744
R454 VTAIL.n28 VTAIL.n17 171.744
R455 VTAIL.n35 VTAIL.n17 171.744
R456 VTAIL.n36 VTAIL.n35 171.744
R457 VTAIL.n36 VTAIL.n13 171.744
R458 VTAIL.n44 VTAIL.n13 171.744
R459 VTAIL.n45 VTAIL.n44 171.744
R460 VTAIL.n46 VTAIL.n45 171.744
R461 VTAIL.n46 VTAIL.n9 171.744
R462 VTAIL.n53 VTAIL.n9 171.744
R463 VTAIL.n54 VTAIL.n53 171.744
R464 VTAIL.n54 VTAIL.n5 171.744
R465 VTAIL.n61 VTAIL.n5 171.744
R466 VTAIL.n62 VTAIL.n61 171.744
R467 VTAIL.n206 VTAIL.n205 171.744
R468 VTAIL.n205 VTAIL.n149 171.744
R469 VTAIL.n198 VTAIL.n149 171.744
R470 VTAIL.n198 VTAIL.n197 171.744
R471 VTAIL.n197 VTAIL.n153 171.744
R472 VTAIL.n190 VTAIL.n153 171.744
R473 VTAIL.n190 VTAIL.n189 171.744
R474 VTAIL.n189 VTAIL.n188 171.744
R475 VTAIL.n188 VTAIL.n157 171.744
R476 VTAIL.n181 VTAIL.n157 171.744
R477 VTAIL.n181 VTAIL.n180 171.744
R478 VTAIL.n180 VTAIL.n162 171.744
R479 VTAIL.n173 VTAIL.n162 171.744
R480 VTAIL.n173 VTAIL.n172 171.744
R481 VTAIL.n172 VTAIL.n166 171.744
R482 VTAIL.n136 VTAIL.n135 171.744
R483 VTAIL.n135 VTAIL.n79 171.744
R484 VTAIL.n128 VTAIL.n79 171.744
R485 VTAIL.n128 VTAIL.n127 171.744
R486 VTAIL.n127 VTAIL.n83 171.744
R487 VTAIL.n120 VTAIL.n83 171.744
R488 VTAIL.n120 VTAIL.n119 171.744
R489 VTAIL.n119 VTAIL.n118 171.744
R490 VTAIL.n118 VTAIL.n87 171.744
R491 VTAIL.n111 VTAIL.n87 171.744
R492 VTAIL.n111 VTAIL.n110 171.744
R493 VTAIL.n110 VTAIL.n92 171.744
R494 VTAIL.n103 VTAIL.n92 171.744
R495 VTAIL.n103 VTAIL.n102 171.744
R496 VTAIL.n102 VTAIL.n96 171.744
R497 VTAIL.t2 VTAIL.n231 85.8723
R498 VTAIL.t13 VTAIL.n21 85.8723
R499 VTAIL.t8 VTAIL.n166 85.8723
R500 VTAIL.t19 VTAIL.n96 85.8723
R501 VTAIL.n145 VTAIL.n144 57.7422
R502 VTAIL.n143 VTAIL.n142 57.7422
R503 VTAIL.n75 VTAIL.n74 57.7422
R504 VTAIL.n73 VTAIL.n72 57.7422
R505 VTAIL.n279 VTAIL.n278 57.7421
R506 VTAIL.n1 VTAIL.n0 57.7421
R507 VTAIL.n69 VTAIL.n68 57.7421
R508 VTAIL.n71 VTAIL.n70 57.7421
R509 VTAIL.n277 VTAIL.n276 32.7672
R510 VTAIL.n67 VTAIL.n66 32.7672
R511 VTAIL.n211 VTAIL.n210 32.7672
R512 VTAIL.n141 VTAIL.n140 32.7672
R513 VTAIL.n73 VTAIL.n71 28.1686
R514 VTAIL.n277 VTAIL.n211 25.5048
R515 VTAIL.n257 VTAIL.n222 13.1884
R516 VTAIL.n47 VTAIL.n12 13.1884
R517 VTAIL.n191 VTAIL.n156 13.1884
R518 VTAIL.n121 VTAIL.n86 13.1884
R519 VTAIL.n253 VTAIL.n252 12.8005
R520 VTAIL.n258 VTAIL.n220 12.8005
R521 VTAIL.n43 VTAIL.n42 12.8005
R522 VTAIL.n48 VTAIL.n10 12.8005
R523 VTAIL.n192 VTAIL.n154 12.8005
R524 VTAIL.n187 VTAIL.n158 12.8005
R525 VTAIL.n122 VTAIL.n84 12.8005
R526 VTAIL.n117 VTAIL.n88 12.8005
R527 VTAIL.n251 VTAIL.n224 12.0247
R528 VTAIL.n262 VTAIL.n261 12.0247
R529 VTAIL.n41 VTAIL.n14 12.0247
R530 VTAIL.n52 VTAIL.n51 12.0247
R531 VTAIL.n196 VTAIL.n195 12.0247
R532 VTAIL.n186 VTAIL.n159 12.0247
R533 VTAIL.n126 VTAIL.n125 12.0247
R534 VTAIL.n116 VTAIL.n89 12.0247
R535 VTAIL.n248 VTAIL.n247 11.249
R536 VTAIL.n265 VTAIL.n218 11.249
R537 VTAIL.n38 VTAIL.n37 11.249
R538 VTAIL.n55 VTAIL.n8 11.249
R539 VTAIL.n199 VTAIL.n152 11.249
R540 VTAIL.n183 VTAIL.n182 11.249
R541 VTAIL.n129 VTAIL.n82 11.249
R542 VTAIL.n113 VTAIL.n112 11.249
R543 VTAIL.n233 VTAIL.n232 10.7239
R544 VTAIL.n23 VTAIL.n22 10.7239
R545 VTAIL.n168 VTAIL.n167 10.7239
R546 VTAIL.n98 VTAIL.n97 10.7239
R547 VTAIL.n244 VTAIL.n226 10.4732
R548 VTAIL.n266 VTAIL.n216 10.4732
R549 VTAIL.n34 VTAIL.n16 10.4732
R550 VTAIL.n56 VTAIL.n6 10.4732
R551 VTAIL.n200 VTAIL.n150 10.4732
R552 VTAIL.n179 VTAIL.n161 10.4732
R553 VTAIL.n130 VTAIL.n80 10.4732
R554 VTAIL.n109 VTAIL.n91 10.4732
R555 VTAIL.n243 VTAIL.n228 9.69747
R556 VTAIL.n270 VTAIL.n269 9.69747
R557 VTAIL.n33 VTAIL.n18 9.69747
R558 VTAIL.n60 VTAIL.n59 9.69747
R559 VTAIL.n204 VTAIL.n203 9.69747
R560 VTAIL.n178 VTAIL.n163 9.69747
R561 VTAIL.n134 VTAIL.n133 9.69747
R562 VTAIL.n108 VTAIL.n93 9.69747
R563 VTAIL.n276 VTAIL.n275 9.45567
R564 VTAIL.n66 VTAIL.n65 9.45567
R565 VTAIL.n210 VTAIL.n209 9.45567
R566 VTAIL.n140 VTAIL.n139 9.45567
R567 VTAIL.n275 VTAIL.n274 9.3005
R568 VTAIL.n214 VTAIL.n213 9.3005
R569 VTAIL.n269 VTAIL.n268 9.3005
R570 VTAIL.n267 VTAIL.n266 9.3005
R571 VTAIL.n218 VTAIL.n217 9.3005
R572 VTAIL.n261 VTAIL.n260 9.3005
R573 VTAIL.n259 VTAIL.n258 9.3005
R574 VTAIL.n235 VTAIL.n234 9.3005
R575 VTAIL.n230 VTAIL.n229 9.3005
R576 VTAIL.n241 VTAIL.n240 9.3005
R577 VTAIL.n243 VTAIL.n242 9.3005
R578 VTAIL.n226 VTAIL.n225 9.3005
R579 VTAIL.n249 VTAIL.n248 9.3005
R580 VTAIL.n251 VTAIL.n250 9.3005
R581 VTAIL.n252 VTAIL.n221 9.3005
R582 VTAIL.n65 VTAIL.n64 9.3005
R583 VTAIL.n4 VTAIL.n3 9.3005
R584 VTAIL.n59 VTAIL.n58 9.3005
R585 VTAIL.n57 VTAIL.n56 9.3005
R586 VTAIL.n8 VTAIL.n7 9.3005
R587 VTAIL.n51 VTAIL.n50 9.3005
R588 VTAIL.n49 VTAIL.n48 9.3005
R589 VTAIL.n25 VTAIL.n24 9.3005
R590 VTAIL.n20 VTAIL.n19 9.3005
R591 VTAIL.n31 VTAIL.n30 9.3005
R592 VTAIL.n33 VTAIL.n32 9.3005
R593 VTAIL.n16 VTAIL.n15 9.3005
R594 VTAIL.n39 VTAIL.n38 9.3005
R595 VTAIL.n41 VTAIL.n40 9.3005
R596 VTAIL.n42 VTAIL.n11 9.3005
R597 VTAIL.n170 VTAIL.n169 9.3005
R598 VTAIL.n165 VTAIL.n164 9.3005
R599 VTAIL.n176 VTAIL.n175 9.3005
R600 VTAIL.n178 VTAIL.n177 9.3005
R601 VTAIL.n161 VTAIL.n160 9.3005
R602 VTAIL.n184 VTAIL.n183 9.3005
R603 VTAIL.n186 VTAIL.n185 9.3005
R604 VTAIL.n158 VTAIL.n155 9.3005
R605 VTAIL.n209 VTAIL.n208 9.3005
R606 VTAIL.n148 VTAIL.n147 9.3005
R607 VTAIL.n203 VTAIL.n202 9.3005
R608 VTAIL.n201 VTAIL.n200 9.3005
R609 VTAIL.n152 VTAIL.n151 9.3005
R610 VTAIL.n195 VTAIL.n194 9.3005
R611 VTAIL.n193 VTAIL.n192 9.3005
R612 VTAIL.n100 VTAIL.n99 9.3005
R613 VTAIL.n95 VTAIL.n94 9.3005
R614 VTAIL.n106 VTAIL.n105 9.3005
R615 VTAIL.n108 VTAIL.n107 9.3005
R616 VTAIL.n91 VTAIL.n90 9.3005
R617 VTAIL.n114 VTAIL.n113 9.3005
R618 VTAIL.n116 VTAIL.n115 9.3005
R619 VTAIL.n88 VTAIL.n85 9.3005
R620 VTAIL.n139 VTAIL.n138 9.3005
R621 VTAIL.n78 VTAIL.n77 9.3005
R622 VTAIL.n133 VTAIL.n132 9.3005
R623 VTAIL.n131 VTAIL.n130 9.3005
R624 VTAIL.n82 VTAIL.n81 9.3005
R625 VTAIL.n125 VTAIL.n124 9.3005
R626 VTAIL.n123 VTAIL.n122 9.3005
R627 VTAIL.n240 VTAIL.n239 8.92171
R628 VTAIL.n273 VTAIL.n214 8.92171
R629 VTAIL.n30 VTAIL.n29 8.92171
R630 VTAIL.n63 VTAIL.n4 8.92171
R631 VTAIL.n207 VTAIL.n148 8.92171
R632 VTAIL.n175 VTAIL.n174 8.92171
R633 VTAIL.n137 VTAIL.n78 8.92171
R634 VTAIL.n105 VTAIL.n104 8.92171
R635 VTAIL.n236 VTAIL.n230 8.14595
R636 VTAIL.n274 VTAIL.n212 8.14595
R637 VTAIL.n26 VTAIL.n20 8.14595
R638 VTAIL.n64 VTAIL.n2 8.14595
R639 VTAIL.n208 VTAIL.n146 8.14595
R640 VTAIL.n171 VTAIL.n165 8.14595
R641 VTAIL.n138 VTAIL.n76 8.14595
R642 VTAIL.n101 VTAIL.n95 8.14595
R643 VTAIL.n235 VTAIL.n232 7.3702
R644 VTAIL.n25 VTAIL.n22 7.3702
R645 VTAIL.n170 VTAIL.n167 7.3702
R646 VTAIL.n100 VTAIL.n97 7.3702
R647 VTAIL.n236 VTAIL.n235 5.81868
R648 VTAIL.n276 VTAIL.n212 5.81868
R649 VTAIL.n26 VTAIL.n25 5.81868
R650 VTAIL.n66 VTAIL.n2 5.81868
R651 VTAIL.n210 VTAIL.n146 5.81868
R652 VTAIL.n171 VTAIL.n170 5.81868
R653 VTAIL.n140 VTAIL.n76 5.81868
R654 VTAIL.n101 VTAIL.n100 5.81868
R655 VTAIL.n239 VTAIL.n230 5.04292
R656 VTAIL.n274 VTAIL.n273 5.04292
R657 VTAIL.n29 VTAIL.n20 5.04292
R658 VTAIL.n64 VTAIL.n63 5.04292
R659 VTAIL.n208 VTAIL.n207 5.04292
R660 VTAIL.n174 VTAIL.n165 5.04292
R661 VTAIL.n138 VTAIL.n137 5.04292
R662 VTAIL.n104 VTAIL.n95 5.04292
R663 VTAIL.n240 VTAIL.n228 4.26717
R664 VTAIL.n270 VTAIL.n214 4.26717
R665 VTAIL.n30 VTAIL.n18 4.26717
R666 VTAIL.n60 VTAIL.n4 4.26717
R667 VTAIL.n204 VTAIL.n148 4.26717
R668 VTAIL.n175 VTAIL.n163 4.26717
R669 VTAIL.n134 VTAIL.n78 4.26717
R670 VTAIL.n105 VTAIL.n93 4.26717
R671 VTAIL.n244 VTAIL.n243 3.49141
R672 VTAIL.n269 VTAIL.n216 3.49141
R673 VTAIL.n34 VTAIL.n33 3.49141
R674 VTAIL.n59 VTAIL.n6 3.49141
R675 VTAIL.n203 VTAIL.n150 3.49141
R676 VTAIL.n179 VTAIL.n178 3.49141
R677 VTAIL.n133 VTAIL.n80 3.49141
R678 VTAIL.n109 VTAIL.n108 3.49141
R679 VTAIL.n247 VTAIL.n226 2.71565
R680 VTAIL.n266 VTAIL.n265 2.71565
R681 VTAIL.n37 VTAIL.n16 2.71565
R682 VTAIL.n56 VTAIL.n55 2.71565
R683 VTAIL.n200 VTAIL.n199 2.71565
R684 VTAIL.n182 VTAIL.n161 2.71565
R685 VTAIL.n130 VTAIL.n129 2.71565
R686 VTAIL.n112 VTAIL.n91 2.71565
R687 VTAIL.n278 VTAIL.t0 2.67581
R688 VTAIL.n278 VTAIL.t3 2.67581
R689 VTAIL.n0 VTAIL.t6 2.67581
R690 VTAIL.n0 VTAIL.t18 2.67581
R691 VTAIL.n68 VTAIL.t12 2.67581
R692 VTAIL.n68 VTAIL.t17 2.67581
R693 VTAIL.n70 VTAIL.t16 2.67581
R694 VTAIL.n70 VTAIL.t15 2.67581
R695 VTAIL.n144 VTAIL.t11 2.67581
R696 VTAIL.n144 VTAIL.t10 2.67581
R697 VTAIL.n142 VTAIL.t9 2.67581
R698 VTAIL.n142 VTAIL.t14 2.67581
R699 VTAIL.n74 VTAIL.t7 2.67581
R700 VTAIL.n74 VTAIL.t5 2.67581
R701 VTAIL.n72 VTAIL.t1 2.67581
R702 VTAIL.n72 VTAIL.t4 2.67581
R703 VTAIL.n75 VTAIL.n73 2.66429
R704 VTAIL.n141 VTAIL.n75 2.66429
R705 VTAIL.n145 VTAIL.n143 2.66429
R706 VTAIL.n211 VTAIL.n145 2.66429
R707 VTAIL.n71 VTAIL.n69 2.66429
R708 VTAIL.n69 VTAIL.n67 2.66429
R709 VTAIL.n279 VTAIL.n277 2.66429
R710 VTAIL.n169 VTAIL.n168 2.41282
R711 VTAIL.n99 VTAIL.n98 2.41282
R712 VTAIL.n234 VTAIL.n233 2.41282
R713 VTAIL.n24 VTAIL.n23 2.41282
R714 VTAIL VTAIL.n1 2.05653
R715 VTAIL.n248 VTAIL.n224 1.93989
R716 VTAIL.n262 VTAIL.n218 1.93989
R717 VTAIL.n38 VTAIL.n14 1.93989
R718 VTAIL.n52 VTAIL.n8 1.93989
R719 VTAIL.n196 VTAIL.n152 1.93989
R720 VTAIL.n183 VTAIL.n159 1.93989
R721 VTAIL.n126 VTAIL.n82 1.93989
R722 VTAIL.n113 VTAIL.n89 1.93989
R723 VTAIL.n143 VTAIL.n141 1.80222
R724 VTAIL.n67 VTAIL.n1 1.80222
R725 VTAIL.n253 VTAIL.n251 1.16414
R726 VTAIL.n261 VTAIL.n220 1.16414
R727 VTAIL.n43 VTAIL.n41 1.16414
R728 VTAIL.n51 VTAIL.n10 1.16414
R729 VTAIL.n195 VTAIL.n154 1.16414
R730 VTAIL.n187 VTAIL.n186 1.16414
R731 VTAIL.n125 VTAIL.n84 1.16414
R732 VTAIL.n117 VTAIL.n116 1.16414
R733 VTAIL VTAIL.n279 0.608259
R734 VTAIL.n252 VTAIL.n222 0.388379
R735 VTAIL.n258 VTAIL.n257 0.388379
R736 VTAIL.n42 VTAIL.n12 0.388379
R737 VTAIL.n48 VTAIL.n47 0.388379
R738 VTAIL.n192 VTAIL.n191 0.388379
R739 VTAIL.n158 VTAIL.n156 0.388379
R740 VTAIL.n122 VTAIL.n121 0.388379
R741 VTAIL.n88 VTAIL.n86 0.388379
R742 VTAIL.n234 VTAIL.n229 0.155672
R743 VTAIL.n241 VTAIL.n229 0.155672
R744 VTAIL.n242 VTAIL.n241 0.155672
R745 VTAIL.n242 VTAIL.n225 0.155672
R746 VTAIL.n249 VTAIL.n225 0.155672
R747 VTAIL.n250 VTAIL.n249 0.155672
R748 VTAIL.n250 VTAIL.n221 0.155672
R749 VTAIL.n259 VTAIL.n221 0.155672
R750 VTAIL.n260 VTAIL.n259 0.155672
R751 VTAIL.n260 VTAIL.n217 0.155672
R752 VTAIL.n267 VTAIL.n217 0.155672
R753 VTAIL.n268 VTAIL.n267 0.155672
R754 VTAIL.n268 VTAIL.n213 0.155672
R755 VTAIL.n275 VTAIL.n213 0.155672
R756 VTAIL.n24 VTAIL.n19 0.155672
R757 VTAIL.n31 VTAIL.n19 0.155672
R758 VTAIL.n32 VTAIL.n31 0.155672
R759 VTAIL.n32 VTAIL.n15 0.155672
R760 VTAIL.n39 VTAIL.n15 0.155672
R761 VTAIL.n40 VTAIL.n39 0.155672
R762 VTAIL.n40 VTAIL.n11 0.155672
R763 VTAIL.n49 VTAIL.n11 0.155672
R764 VTAIL.n50 VTAIL.n49 0.155672
R765 VTAIL.n50 VTAIL.n7 0.155672
R766 VTAIL.n57 VTAIL.n7 0.155672
R767 VTAIL.n58 VTAIL.n57 0.155672
R768 VTAIL.n58 VTAIL.n3 0.155672
R769 VTAIL.n65 VTAIL.n3 0.155672
R770 VTAIL.n209 VTAIL.n147 0.155672
R771 VTAIL.n202 VTAIL.n147 0.155672
R772 VTAIL.n202 VTAIL.n201 0.155672
R773 VTAIL.n201 VTAIL.n151 0.155672
R774 VTAIL.n194 VTAIL.n151 0.155672
R775 VTAIL.n194 VTAIL.n193 0.155672
R776 VTAIL.n193 VTAIL.n155 0.155672
R777 VTAIL.n185 VTAIL.n155 0.155672
R778 VTAIL.n185 VTAIL.n184 0.155672
R779 VTAIL.n184 VTAIL.n160 0.155672
R780 VTAIL.n177 VTAIL.n160 0.155672
R781 VTAIL.n177 VTAIL.n176 0.155672
R782 VTAIL.n176 VTAIL.n164 0.155672
R783 VTAIL.n169 VTAIL.n164 0.155672
R784 VTAIL.n139 VTAIL.n77 0.155672
R785 VTAIL.n132 VTAIL.n77 0.155672
R786 VTAIL.n132 VTAIL.n131 0.155672
R787 VTAIL.n131 VTAIL.n81 0.155672
R788 VTAIL.n124 VTAIL.n81 0.155672
R789 VTAIL.n124 VTAIL.n123 0.155672
R790 VTAIL.n123 VTAIL.n85 0.155672
R791 VTAIL.n115 VTAIL.n85 0.155672
R792 VTAIL.n115 VTAIL.n114 0.155672
R793 VTAIL.n114 VTAIL.n90 0.155672
R794 VTAIL.n107 VTAIL.n90 0.155672
R795 VTAIL.n107 VTAIL.n106 0.155672
R796 VTAIL.n106 VTAIL.n94 0.155672
R797 VTAIL.n99 VTAIL.n94 0.155672
R798 VN.n82 VN.n81 161.3
R799 VN.n80 VN.n43 161.3
R800 VN.n79 VN.n78 161.3
R801 VN.n77 VN.n44 161.3
R802 VN.n76 VN.n75 161.3
R803 VN.n74 VN.n45 161.3
R804 VN.n72 VN.n71 161.3
R805 VN.n70 VN.n46 161.3
R806 VN.n69 VN.n68 161.3
R807 VN.n67 VN.n47 161.3
R808 VN.n66 VN.n65 161.3
R809 VN.n64 VN.n48 161.3
R810 VN.n63 VN.n62 161.3
R811 VN.n61 VN.n49 161.3
R812 VN.n60 VN.n59 161.3
R813 VN.n58 VN.n51 161.3
R814 VN.n57 VN.n56 161.3
R815 VN.n55 VN.n52 161.3
R816 VN.n40 VN.n39 161.3
R817 VN.n38 VN.n1 161.3
R818 VN.n37 VN.n36 161.3
R819 VN.n35 VN.n2 161.3
R820 VN.n34 VN.n33 161.3
R821 VN.n32 VN.n3 161.3
R822 VN.n30 VN.n29 161.3
R823 VN.n28 VN.n4 161.3
R824 VN.n27 VN.n26 161.3
R825 VN.n25 VN.n5 161.3
R826 VN.n24 VN.n23 161.3
R827 VN.n22 VN.n6 161.3
R828 VN.n21 VN.n20 161.3
R829 VN.n18 VN.n7 161.3
R830 VN.n17 VN.n16 161.3
R831 VN.n15 VN.n8 161.3
R832 VN.n14 VN.n13 161.3
R833 VN.n12 VN.n9 161.3
R834 VN.n53 VN.t3 137.976
R835 VN.n10 VN.t5 137.976
R836 VN.n11 VN.t4 106.093
R837 VN.n19 VN.t2 106.093
R838 VN.n31 VN.t7 106.093
R839 VN.n0 VN.t0 106.093
R840 VN.n54 VN.t8 106.093
R841 VN.n50 VN.t1 106.093
R842 VN.n73 VN.t6 106.093
R843 VN.n42 VN.t9 106.093
R844 VN.n41 VN.n0 69.0258
R845 VN.n83 VN.n42 69.0258
R846 VN.n11 VN.n10 56.938
R847 VN.n54 VN.n53 56.938
R848 VN.n17 VN.n8 56.5193
R849 VN.n26 VN.n25 56.5193
R850 VN.n60 VN.n51 56.5193
R851 VN.n68 VN.n67 56.5193
R852 VN VN.n83 54.3427
R853 VN.n37 VN.n2 51.663
R854 VN.n79 VN.n44 51.663
R855 VN.n38 VN.n37 29.3238
R856 VN.n80 VN.n79 29.3238
R857 VN.n13 VN.n12 24.4675
R858 VN.n13 VN.n8 24.4675
R859 VN.n18 VN.n17 24.4675
R860 VN.n20 VN.n18 24.4675
R861 VN.n24 VN.n6 24.4675
R862 VN.n25 VN.n24 24.4675
R863 VN.n26 VN.n4 24.4675
R864 VN.n30 VN.n4 24.4675
R865 VN.n33 VN.n32 24.4675
R866 VN.n33 VN.n2 24.4675
R867 VN.n39 VN.n38 24.4675
R868 VN.n56 VN.n51 24.4675
R869 VN.n56 VN.n55 24.4675
R870 VN.n67 VN.n66 24.4675
R871 VN.n66 VN.n48 24.4675
R872 VN.n62 VN.n61 24.4675
R873 VN.n61 VN.n60 24.4675
R874 VN.n75 VN.n44 24.4675
R875 VN.n75 VN.n74 24.4675
R876 VN.n72 VN.n46 24.4675
R877 VN.n68 VN.n46 24.4675
R878 VN.n81 VN.n80 24.4675
R879 VN.n39 VN.n0 21.0421
R880 VN.n81 VN.n42 21.0421
R881 VN.n12 VN.n11 16.6381
R882 VN.n31 VN.n30 16.6381
R883 VN.n55 VN.n54 16.6381
R884 VN.n73 VN.n72 16.6381
R885 VN.n20 VN.n19 12.234
R886 VN.n19 VN.n6 12.234
R887 VN.n50 VN.n48 12.234
R888 VN.n62 VN.n50 12.234
R889 VN.n32 VN.n31 7.82994
R890 VN.n74 VN.n73 7.82994
R891 VN.n53 VN.n52 5.45824
R892 VN.n10 VN.n9 5.45823
R893 VN.n83 VN.n82 0.354971
R894 VN.n41 VN.n40 0.354971
R895 VN VN.n41 0.26696
R896 VN.n82 VN.n43 0.189894
R897 VN.n78 VN.n43 0.189894
R898 VN.n78 VN.n77 0.189894
R899 VN.n77 VN.n76 0.189894
R900 VN.n76 VN.n45 0.189894
R901 VN.n71 VN.n45 0.189894
R902 VN.n71 VN.n70 0.189894
R903 VN.n70 VN.n69 0.189894
R904 VN.n69 VN.n47 0.189894
R905 VN.n65 VN.n47 0.189894
R906 VN.n65 VN.n64 0.189894
R907 VN.n64 VN.n63 0.189894
R908 VN.n63 VN.n49 0.189894
R909 VN.n59 VN.n49 0.189894
R910 VN.n59 VN.n58 0.189894
R911 VN.n58 VN.n57 0.189894
R912 VN.n57 VN.n52 0.189894
R913 VN.n14 VN.n9 0.189894
R914 VN.n15 VN.n14 0.189894
R915 VN.n16 VN.n15 0.189894
R916 VN.n16 VN.n7 0.189894
R917 VN.n21 VN.n7 0.189894
R918 VN.n22 VN.n21 0.189894
R919 VN.n23 VN.n22 0.189894
R920 VN.n23 VN.n5 0.189894
R921 VN.n27 VN.n5 0.189894
R922 VN.n28 VN.n27 0.189894
R923 VN.n29 VN.n28 0.189894
R924 VN.n29 VN.n3 0.189894
R925 VN.n34 VN.n3 0.189894
R926 VN.n35 VN.n34 0.189894
R927 VN.n36 VN.n35 0.189894
R928 VN.n36 VN.n1 0.189894
R929 VN.n40 VN.n1 0.189894
R930 VDD2.n129 VDD2.n69 756.745
R931 VDD2.n60 VDD2.n0 756.745
R932 VDD2.n130 VDD2.n129 585
R933 VDD2.n128 VDD2.n127 585
R934 VDD2.n73 VDD2.n72 585
R935 VDD2.n122 VDD2.n121 585
R936 VDD2.n120 VDD2.n119 585
R937 VDD2.n77 VDD2.n76 585
R938 VDD2.n114 VDD2.n113 585
R939 VDD2.n112 VDD2.n79 585
R940 VDD2.n111 VDD2.n110 585
R941 VDD2.n82 VDD2.n80 585
R942 VDD2.n105 VDD2.n104 585
R943 VDD2.n103 VDD2.n102 585
R944 VDD2.n86 VDD2.n85 585
R945 VDD2.n97 VDD2.n96 585
R946 VDD2.n95 VDD2.n94 585
R947 VDD2.n90 VDD2.n89 585
R948 VDD2.n20 VDD2.n19 585
R949 VDD2.n25 VDD2.n24 585
R950 VDD2.n27 VDD2.n26 585
R951 VDD2.n16 VDD2.n15 585
R952 VDD2.n33 VDD2.n32 585
R953 VDD2.n35 VDD2.n34 585
R954 VDD2.n12 VDD2.n11 585
R955 VDD2.n42 VDD2.n41 585
R956 VDD2.n43 VDD2.n10 585
R957 VDD2.n45 VDD2.n44 585
R958 VDD2.n8 VDD2.n7 585
R959 VDD2.n51 VDD2.n50 585
R960 VDD2.n53 VDD2.n52 585
R961 VDD2.n4 VDD2.n3 585
R962 VDD2.n59 VDD2.n58 585
R963 VDD2.n61 VDD2.n60 585
R964 VDD2.n91 VDD2.t0 329.036
R965 VDD2.n21 VDD2.t4 329.036
R966 VDD2.n129 VDD2.n128 171.744
R967 VDD2.n128 VDD2.n72 171.744
R968 VDD2.n121 VDD2.n72 171.744
R969 VDD2.n121 VDD2.n120 171.744
R970 VDD2.n120 VDD2.n76 171.744
R971 VDD2.n113 VDD2.n76 171.744
R972 VDD2.n113 VDD2.n112 171.744
R973 VDD2.n112 VDD2.n111 171.744
R974 VDD2.n111 VDD2.n80 171.744
R975 VDD2.n104 VDD2.n80 171.744
R976 VDD2.n104 VDD2.n103 171.744
R977 VDD2.n103 VDD2.n85 171.744
R978 VDD2.n96 VDD2.n85 171.744
R979 VDD2.n96 VDD2.n95 171.744
R980 VDD2.n95 VDD2.n89 171.744
R981 VDD2.n25 VDD2.n19 171.744
R982 VDD2.n26 VDD2.n25 171.744
R983 VDD2.n26 VDD2.n15 171.744
R984 VDD2.n33 VDD2.n15 171.744
R985 VDD2.n34 VDD2.n33 171.744
R986 VDD2.n34 VDD2.n11 171.744
R987 VDD2.n42 VDD2.n11 171.744
R988 VDD2.n43 VDD2.n42 171.744
R989 VDD2.n44 VDD2.n43 171.744
R990 VDD2.n44 VDD2.n7 171.744
R991 VDD2.n51 VDD2.n7 171.744
R992 VDD2.n52 VDD2.n51 171.744
R993 VDD2.n52 VDD2.n3 171.744
R994 VDD2.n59 VDD2.n3 171.744
R995 VDD2.n60 VDD2.n59 171.744
R996 VDD2.t0 VDD2.n89 85.8723
R997 VDD2.t4 VDD2.n19 85.8723
R998 VDD2.n68 VDD2.n67 76.3633
R999 VDD2 VDD2.n137 76.3605
R1000 VDD2.n136 VDD2.n135 74.421
R1001 VDD2.n66 VDD2.n65 74.4208
R1002 VDD2.n66 VDD2.n64 52.1097
R1003 VDD2.n134 VDD2.n133 49.446
R1004 VDD2.n134 VDD2.n68 46.8424
R1005 VDD2.n114 VDD2.n79 13.1884
R1006 VDD2.n45 VDD2.n10 13.1884
R1007 VDD2.n115 VDD2.n77 12.8005
R1008 VDD2.n110 VDD2.n81 12.8005
R1009 VDD2.n41 VDD2.n40 12.8005
R1010 VDD2.n46 VDD2.n8 12.8005
R1011 VDD2.n119 VDD2.n118 12.0247
R1012 VDD2.n109 VDD2.n82 12.0247
R1013 VDD2.n39 VDD2.n12 12.0247
R1014 VDD2.n50 VDD2.n49 12.0247
R1015 VDD2.n122 VDD2.n75 11.249
R1016 VDD2.n106 VDD2.n105 11.249
R1017 VDD2.n36 VDD2.n35 11.249
R1018 VDD2.n53 VDD2.n6 11.249
R1019 VDD2.n91 VDD2.n90 10.7239
R1020 VDD2.n21 VDD2.n20 10.7239
R1021 VDD2.n123 VDD2.n73 10.4732
R1022 VDD2.n102 VDD2.n84 10.4732
R1023 VDD2.n32 VDD2.n14 10.4732
R1024 VDD2.n54 VDD2.n4 10.4732
R1025 VDD2.n127 VDD2.n126 9.69747
R1026 VDD2.n101 VDD2.n86 9.69747
R1027 VDD2.n31 VDD2.n16 9.69747
R1028 VDD2.n58 VDD2.n57 9.69747
R1029 VDD2.n133 VDD2.n132 9.45567
R1030 VDD2.n64 VDD2.n63 9.45567
R1031 VDD2.n93 VDD2.n92 9.3005
R1032 VDD2.n88 VDD2.n87 9.3005
R1033 VDD2.n99 VDD2.n98 9.3005
R1034 VDD2.n101 VDD2.n100 9.3005
R1035 VDD2.n84 VDD2.n83 9.3005
R1036 VDD2.n107 VDD2.n106 9.3005
R1037 VDD2.n109 VDD2.n108 9.3005
R1038 VDD2.n81 VDD2.n78 9.3005
R1039 VDD2.n132 VDD2.n131 9.3005
R1040 VDD2.n71 VDD2.n70 9.3005
R1041 VDD2.n126 VDD2.n125 9.3005
R1042 VDD2.n124 VDD2.n123 9.3005
R1043 VDD2.n75 VDD2.n74 9.3005
R1044 VDD2.n118 VDD2.n117 9.3005
R1045 VDD2.n116 VDD2.n115 9.3005
R1046 VDD2.n63 VDD2.n62 9.3005
R1047 VDD2.n2 VDD2.n1 9.3005
R1048 VDD2.n57 VDD2.n56 9.3005
R1049 VDD2.n55 VDD2.n54 9.3005
R1050 VDD2.n6 VDD2.n5 9.3005
R1051 VDD2.n49 VDD2.n48 9.3005
R1052 VDD2.n47 VDD2.n46 9.3005
R1053 VDD2.n23 VDD2.n22 9.3005
R1054 VDD2.n18 VDD2.n17 9.3005
R1055 VDD2.n29 VDD2.n28 9.3005
R1056 VDD2.n31 VDD2.n30 9.3005
R1057 VDD2.n14 VDD2.n13 9.3005
R1058 VDD2.n37 VDD2.n36 9.3005
R1059 VDD2.n39 VDD2.n38 9.3005
R1060 VDD2.n40 VDD2.n9 9.3005
R1061 VDD2.n130 VDD2.n71 8.92171
R1062 VDD2.n98 VDD2.n97 8.92171
R1063 VDD2.n28 VDD2.n27 8.92171
R1064 VDD2.n61 VDD2.n2 8.92171
R1065 VDD2.n131 VDD2.n69 8.14595
R1066 VDD2.n94 VDD2.n88 8.14595
R1067 VDD2.n24 VDD2.n18 8.14595
R1068 VDD2.n62 VDD2.n0 8.14595
R1069 VDD2.n93 VDD2.n90 7.3702
R1070 VDD2.n23 VDD2.n20 7.3702
R1071 VDD2.n133 VDD2.n69 5.81868
R1072 VDD2.n94 VDD2.n93 5.81868
R1073 VDD2.n24 VDD2.n23 5.81868
R1074 VDD2.n64 VDD2.n0 5.81868
R1075 VDD2.n131 VDD2.n130 5.04292
R1076 VDD2.n97 VDD2.n88 5.04292
R1077 VDD2.n27 VDD2.n18 5.04292
R1078 VDD2.n62 VDD2.n61 5.04292
R1079 VDD2.n127 VDD2.n71 4.26717
R1080 VDD2.n98 VDD2.n86 4.26717
R1081 VDD2.n28 VDD2.n16 4.26717
R1082 VDD2.n58 VDD2.n2 4.26717
R1083 VDD2.n126 VDD2.n73 3.49141
R1084 VDD2.n102 VDD2.n101 3.49141
R1085 VDD2.n32 VDD2.n31 3.49141
R1086 VDD2.n57 VDD2.n4 3.49141
R1087 VDD2.n123 VDD2.n122 2.71565
R1088 VDD2.n105 VDD2.n84 2.71565
R1089 VDD2.n35 VDD2.n14 2.71565
R1090 VDD2.n54 VDD2.n53 2.71565
R1091 VDD2.n137 VDD2.t1 2.67581
R1092 VDD2.n137 VDD2.t6 2.67581
R1093 VDD2.n135 VDD2.t3 2.67581
R1094 VDD2.n135 VDD2.t8 2.67581
R1095 VDD2.n67 VDD2.t2 2.67581
R1096 VDD2.n67 VDD2.t9 2.67581
R1097 VDD2.n65 VDD2.t5 2.67581
R1098 VDD2.n65 VDD2.t7 2.67581
R1099 VDD2.n136 VDD2.n134 2.66429
R1100 VDD2.n92 VDD2.n91 2.41282
R1101 VDD2.n22 VDD2.n21 2.41282
R1102 VDD2.n119 VDD2.n75 1.93989
R1103 VDD2.n106 VDD2.n82 1.93989
R1104 VDD2.n36 VDD2.n12 1.93989
R1105 VDD2.n50 VDD2.n6 1.93989
R1106 VDD2.n118 VDD2.n77 1.16414
R1107 VDD2.n110 VDD2.n109 1.16414
R1108 VDD2.n41 VDD2.n39 1.16414
R1109 VDD2.n49 VDD2.n8 1.16414
R1110 VDD2 VDD2.n136 0.724638
R1111 VDD2.n68 VDD2.n66 0.611102
R1112 VDD2.n115 VDD2.n114 0.388379
R1113 VDD2.n81 VDD2.n79 0.388379
R1114 VDD2.n40 VDD2.n10 0.388379
R1115 VDD2.n46 VDD2.n45 0.388379
R1116 VDD2.n132 VDD2.n70 0.155672
R1117 VDD2.n125 VDD2.n70 0.155672
R1118 VDD2.n125 VDD2.n124 0.155672
R1119 VDD2.n124 VDD2.n74 0.155672
R1120 VDD2.n117 VDD2.n74 0.155672
R1121 VDD2.n117 VDD2.n116 0.155672
R1122 VDD2.n116 VDD2.n78 0.155672
R1123 VDD2.n108 VDD2.n78 0.155672
R1124 VDD2.n108 VDD2.n107 0.155672
R1125 VDD2.n107 VDD2.n83 0.155672
R1126 VDD2.n100 VDD2.n83 0.155672
R1127 VDD2.n100 VDD2.n99 0.155672
R1128 VDD2.n99 VDD2.n87 0.155672
R1129 VDD2.n92 VDD2.n87 0.155672
R1130 VDD2.n22 VDD2.n17 0.155672
R1131 VDD2.n29 VDD2.n17 0.155672
R1132 VDD2.n30 VDD2.n29 0.155672
R1133 VDD2.n30 VDD2.n13 0.155672
R1134 VDD2.n37 VDD2.n13 0.155672
R1135 VDD2.n38 VDD2.n37 0.155672
R1136 VDD2.n38 VDD2.n9 0.155672
R1137 VDD2.n47 VDD2.n9 0.155672
R1138 VDD2.n48 VDD2.n47 0.155672
R1139 VDD2.n48 VDD2.n5 0.155672
R1140 VDD2.n55 VDD2.n5 0.155672
R1141 VDD2.n56 VDD2.n55 0.155672
R1142 VDD2.n56 VDD2.n1 0.155672
R1143 VDD2.n63 VDD2.n1 0.155672
R1144 B.n463 B.n462 585
R1145 B.n461 B.n148 585
R1146 B.n460 B.n459 585
R1147 B.n458 B.n149 585
R1148 B.n457 B.n456 585
R1149 B.n455 B.n150 585
R1150 B.n454 B.n453 585
R1151 B.n452 B.n151 585
R1152 B.n451 B.n450 585
R1153 B.n449 B.n152 585
R1154 B.n448 B.n447 585
R1155 B.n446 B.n153 585
R1156 B.n445 B.n444 585
R1157 B.n443 B.n154 585
R1158 B.n442 B.n441 585
R1159 B.n440 B.n155 585
R1160 B.n439 B.n438 585
R1161 B.n437 B.n156 585
R1162 B.n436 B.n435 585
R1163 B.n434 B.n157 585
R1164 B.n433 B.n432 585
R1165 B.n431 B.n158 585
R1166 B.n430 B.n429 585
R1167 B.n428 B.n159 585
R1168 B.n427 B.n426 585
R1169 B.n425 B.n160 585
R1170 B.n424 B.n423 585
R1171 B.n422 B.n161 585
R1172 B.n421 B.n420 585
R1173 B.n419 B.n162 585
R1174 B.n418 B.n417 585
R1175 B.n416 B.n163 585
R1176 B.n415 B.n414 585
R1177 B.n413 B.n164 585
R1178 B.n412 B.n411 585
R1179 B.n410 B.n165 585
R1180 B.n409 B.n408 585
R1181 B.n407 B.n166 585
R1182 B.n406 B.n405 585
R1183 B.n404 B.n167 585
R1184 B.n403 B.n402 585
R1185 B.n401 B.n168 585
R1186 B.n400 B.n399 585
R1187 B.n395 B.n169 585
R1188 B.n394 B.n393 585
R1189 B.n392 B.n170 585
R1190 B.n391 B.n390 585
R1191 B.n389 B.n171 585
R1192 B.n388 B.n387 585
R1193 B.n386 B.n172 585
R1194 B.n385 B.n384 585
R1195 B.n383 B.n173 585
R1196 B.n381 B.n380 585
R1197 B.n379 B.n176 585
R1198 B.n378 B.n377 585
R1199 B.n376 B.n177 585
R1200 B.n375 B.n374 585
R1201 B.n373 B.n178 585
R1202 B.n372 B.n371 585
R1203 B.n370 B.n179 585
R1204 B.n369 B.n368 585
R1205 B.n367 B.n180 585
R1206 B.n366 B.n365 585
R1207 B.n364 B.n181 585
R1208 B.n363 B.n362 585
R1209 B.n361 B.n182 585
R1210 B.n360 B.n359 585
R1211 B.n358 B.n183 585
R1212 B.n357 B.n356 585
R1213 B.n355 B.n184 585
R1214 B.n354 B.n353 585
R1215 B.n352 B.n185 585
R1216 B.n351 B.n350 585
R1217 B.n349 B.n186 585
R1218 B.n348 B.n347 585
R1219 B.n346 B.n187 585
R1220 B.n345 B.n344 585
R1221 B.n343 B.n188 585
R1222 B.n342 B.n341 585
R1223 B.n340 B.n189 585
R1224 B.n339 B.n338 585
R1225 B.n337 B.n190 585
R1226 B.n336 B.n335 585
R1227 B.n334 B.n191 585
R1228 B.n333 B.n332 585
R1229 B.n331 B.n192 585
R1230 B.n330 B.n329 585
R1231 B.n328 B.n193 585
R1232 B.n327 B.n326 585
R1233 B.n325 B.n194 585
R1234 B.n324 B.n323 585
R1235 B.n322 B.n195 585
R1236 B.n321 B.n320 585
R1237 B.n319 B.n196 585
R1238 B.n464 B.n147 585
R1239 B.n466 B.n465 585
R1240 B.n467 B.n146 585
R1241 B.n469 B.n468 585
R1242 B.n470 B.n145 585
R1243 B.n472 B.n471 585
R1244 B.n473 B.n144 585
R1245 B.n475 B.n474 585
R1246 B.n476 B.n143 585
R1247 B.n478 B.n477 585
R1248 B.n479 B.n142 585
R1249 B.n481 B.n480 585
R1250 B.n482 B.n141 585
R1251 B.n484 B.n483 585
R1252 B.n485 B.n140 585
R1253 B.n487 B.n486 585
R1254 B.n488 B.n139 585
R1255 B.n490 B.n489 585
R1256 B.n491 B.n138 585
R1257 B.n493 B.n492 585
R1258 B.n494 B.n137 585
R1259 B.n496 B.n495 585
R1260 B.n497 B.n136 585
R1261 B.n499 B.n498 585
R1262 B.n500 B.n135 585
R1263 B.n502 B.n501 585
R1264 B.n503 B.n134 585
R1265 B.n505 B.n504 585
R1266 B.n506 B.n133 585
R1267 B.n508 B.n507 585
R1268 B.n509 B.n132 585
R1269 B.n511 B.n510 585
R1270 B.n512 B.n131 585
R1271 B.n514 B.n513 585
R1272 B.n515 B.n130 585
R1273 B.n517 B.n516 585
R1274 B.n518 B.n129 585
R1275 B.n520 B.n519 585
R1276 B.n521 B.n128 585
R1277 B.n523 B.n522 585
R1278 B.n524 B.n127 585
R1279 B.n526 B.n525 585
R1280 B.n527 B.n126 585
R1281 B.n529 B.n528 585
R1282 B.n530 B.n125 585
R1283 B.n532 B.n531 585
R1284 B.n533 B.n124 585
R1285 B.n535 B.n534 585
R1286 B.n536 B.n123 585
R1287 B.n538 B.n537 585
R1288 B.n539 B.n122 585
R1289 B.n541 B.n540 585
R1290 B.n542 B.n121 585
R1291 B.n544 B.n543 585
R1292 B.n545 B.n120 585
R1293 B.n547 B.n546 585
R1294 B.n548 B.n119 585
R1295 B.n550 B.n549 585
R1296 B.n551 B.n118 585
R1297 B.n553 B.n552 585
R1298 B.n554 B.n117 585
R1299 B.n556 B.n555 585
R1300 B.n557 B.n116 585
R1301 B.n559 B.n558 585
R1302 B.n560 B.n115 585
R1303 B.n562 B.n561 585
R1304 B.n563 B.n114 585
R1305 B.n565 B.n564 585
R1306 B.n566 B.n113 585
R1307 B.n568 B.n567 585
R1308 B.n569 B.n112 585
R1309 B.n571 B.n570 585
R1310 B.n572 B.n111 585
R1311 B.n574 B.n573 585
R1312 B.n575 B.n110 585
R1313 B.n577 B.n576 585
R1314 B.n578 B.n109 585
R1315 B.n580 B.n579 585
R1316 B.n581 B.n108 585
R1317 B.n583 B.n582 585
R1318 B.n584 B.n107 585
R1319 B.n586 B.n585 585
R1320 B.n587 B.n106 585
R1321 B.n589 B.n588 585
R1322 B.n590 B.n105 585
R1323 B.n592 B.n591 585
R1324 B.n593 B.n104 585
R1325 B.n595 B.n594 585
R1326 B.n596 B.n103 585
R1327 B.n598 B.n597 585
R1328 B.n599 B.n102 585
R1329 B.n601 B.n600 585
R1330 B.n602 B.n101 585
R1331 B.n604 B.n603 585
R1332 B.n605 B.n100 585
R1333 B.n607 B.n606 585
R1334 B.n608 B.n99 585
R1335 B.n610 B.n609 585
R1336 B.n611 B.n98 585
R1337 B.n613 B.n612 585
R1338 B.n614 B.n97 585
R1339 B.n616 B.n615 585
R1340 B.n617 B.n96 585
R1341 B.n619 B.n618 585
R1342 B.n620 B.n95 585
R1343 B.n622 B.n621 585
R1344 B.n623 B.n94 585
R1345 B.n625 B.n624 585
R1346 B.n626 B.n93 585
R1347 B.n628 B.n627 585
R1348 B.n629 B.n92 585
R1349 B.n631 B.n630 585
R1350 B.n632 B.n91 585
R1351 B.n634 B.n633 585
R1352 B.n635 B.n90 585
R1353 B.n637 B.n636 585
R1354 B.n638 B.n89 585
R1355 B.n640 B.n639 585
R1356 B.n641 B.n88 585
R1357 B.n643 B.n642 585
R1358 B.n644 B.n87 585
R1359 B.n646 B.n645 585
R1360 B.n647 B.n86 585
R1361 B.n649 B.n648 585
R1362 B.n650 B.n85 585
R1363 B.n652 B.n651 585
R1364 B.n794 B.n33 585
R1365 B.n793 B.n792 585
R1366 B.n791 B.n34 585
R1367 B.n790 B.n789 585
R1368 B.n788 B.n35 585
R1369 B.n787 B.n786 585
R1370 B.n785 B.n36 585
R1371 B.n784 B.n783 585
R1372 B.n782 B.n37 585
R1373 B.n781 B.n780 585
R1374 B.n779 B.n38 585
R1375 B.n778 B.n777 585
R1376 B.n776 B.n39 585
R1377 B.n775 B.n774 585
R1378 B.n773 B.n40 585
R1379 B.n772 B.n771 585
R1380 B.n770 B.n41 585
R1381 B.n769 B.n768 585
R1382 B.n767 B.n42 585
R1383 B.n766 B.n765 585
R1384 B.n764 B.n43 585
R1385 B.n763 B.n762 585
R1386 B.n761 B.n44 585
R1387 B.n760 B.n759 585
R1388 B.n758 B.n45 585
R1389 B.n757 B.n756 585
R1390 B.n755 B.n46 585
R1391 B.n754 B.n753 585
R1392 B.n752 B.n47 585
R1393 B.n751 B.n750 585
R1394 B.n749 B.n48 585
R1395 B.n748 B.n747 585
R1396 B.n746 B.n49 585
R1397 B.n745 B.n744 585
R1398 B.n743 B.n50 585
R1399 B.n742 B.n741 585
R1400 B.n740 B.n51 585
R1401 B.n739 B.n738 585
R1402 B.n737 B.n52 585
R1403 B.n736 B.n735 585
R1404 B.n734 B.n53 585
R1405 B.n733 B.n732 585
R1406 B.n731 B.n730 585
R1407 B.n729 B.n57 585
R1408 B.n728 B.n727 585
R1409 B.n726 B.n58 585
R1410 B.n725 B.n724 585
R1411 B.n723 B.n59 585
R1412 B.n722 B.n721 585
R1413 B.n720 B.n60 585
R1414 B.n719 B.n718 585
R1415 B.n717 B.n61 585
R1416 B.n715 B.n714 585
R1417 B.n713 B.n64 585
R1418 B.n712 B.n711 585
R1419 B.n710 B.n65 585
R1420 B.n709 B.n708 585
R1421 B.n707 B.n66 585
R1422 B.n706 B.n705 585
R1423 B.n704 B.n67 585
R1424 B.n703 B.n702 585
R1425 B.n701 B.n68 585
R1426 B.n700 B.n699 585
R1427 B.n698 B.n69 585
R1428 B.n697 B.n696 585
R1429 B.n695 B.n70 585
R1430 B.n694 B.n693 585
R1431 B.n692 B.n71 585
R1432 B.n691 B.n690 585
R1433 B.n689 B.n72 585
R1434 B.n688 B.n687 585
R1435 B.n686 B.n73 585
R1436 B.n685 B.n684 585
R1437 B.n683 B.n74 585
R1438 B.n682 B.n681 585
R1439 B.n680 B.n75 585
R1440 B.n679 B.n678 585
R1441 B.n677 B.n76 585
R1442 B.n676 B.n675 585
R1443 B.n674 B.n77 585
R1444 B.n673 B.n672 585
R1445 B.n671 B.n78 585
R1446 B.n670 B.n669 585
R1447 B.n668 B.n79 585
R1448 B.n667 B.n666 585
R1449 B.n665 B.n80 585
R1450 B.n664 B.n663 585
R1451 B.n662 B.n81 585
R1452 B.n661 B.n660 585
R1453 B.n659 B.n82 585
R1454 B.n658 B.n657 585
R1455 B.n656 B.n83 585
R1456 B.n655 B.n654 585
R1457 B.n653 B.n84 585
R1458 B.n796 B.n795 585
R1459 B.n797 B.n32 585
R1460 B.n799 B.n798 585
R1461 B.n800 B.n31 585
R1462 B.n802 B.n801 585
R1463 B.n803 B.n30 585
R1464 B.n805 B.n804 585
R1465 B.n806 B.n29 585
R1466 B.n808 B.n807 585
R1467 B.n809 B.n28 585
R1468 B.n811 B.n810 585
R1469 B.n812 B.n27 585
R1470 B.n814 B.n813 585
R1471 B.n815 B.n26 585
R1472 B.n817 B.n816 585
R1473 B.n818 B.n25 585
R1474 B.n820 B.n819 585
R1475 B.n821 B.n24 585
R1476 B.n823 B.n822 585
R1477 B.n824 B.n23 585
R1478 B.n826 B.n825 585
R1479 B.n827 B.n22 585
R1480 B.n829 B.n828 585
R1481 B.n830 B.n21 585
R1482 B.n832 B.n831 585
R1483 B.n833 B.n20 585
R1484 B.n835 B.n834 585
R1485 B.n836 B.n19 585
R1486 B.n838 B.n837 585
R1487 B.n839 B.n18 585
R1488 B.n841 B.n840 585
R1489 B.n842 B.n17 585
R1490 B.n844 B.n843 585
R1491 B.n845 B.n16 585
R1492 B.n847 B.n846 585
R1493 B.n848 B.n15 585
R1494 B.n850 B.n849 585
R1495 B.n851 B.n14 585
R1496 B.n853 B.n852 585
R1497 B.n854 B.n13 585
R1498 B.n856 B.n855 585
R1499 B.n857 B.n12 585
R1500 B.n859 B.n858 585
R1501 B.n860 B.n11 585
R1502 B.n862 B.n861 585
R1503 B.n863 B.n10 585
R1504 B.n865 B.n864 585
R1505 B.n866 B.n9 585
R1506 B.n868 B.n867 585
R1507 B.n869 B.n8 585
R1508 B.n871 B.n870 585
R1509 B.n872 B.n7 585
R1510 B.n874 B.n873 585
R1511 B.n875 B.n6 585
R1512 B.n877 B.n876 585
R1513 B.n878 B.n5 585
R1514 B.n880 B.n879 585
R1515 B.n881 B.n4 585
R1516 B.n883 B.n882 585
R1517 B.n884 B.n3 585
R1518 B.n886 B.n885 585
R1519 B.n887 B.n0 585
R1520 B.n2 B.n1 585
R1521 B.n228 B.n227 585
R1522 B.n229 B.n226 585
R1523 B.n231 B.n230 585
R1524 B.n232 B.n225 585
R1525 B.n234 B.n233 585
R1526 B.n235 B.n224 585
R1527 B.n237 B.n236 585
R1528 B.n238 B.n223 585
R1529 B.n240 B.n239 585
R1530 B.n241 B.n222 585
R1531 B.n243 B.n242 585
R1532 B.n244 B.n221 585
R1533 B.n246 B.n245 585
R1534 B.n247 B.n220 585
R1535 B.n249 B.n248 585
R1536 B.n250 B.n219 585
R1537 B.n252 B.n251 585
R1538 B.n253 B.n218 585
R1539 B.n255 B.n254 585
R1540 B.n256 B.n217 585
R1541 B.n258 B.n257 585
R1542 B.n259 B.n216 585
R1543 B.n261 B.n260 585
R1544 B.n262 B.n215 585
R1545 B.n264 B.n263 585
R1546 B.n265 B.n214 585
R1547 B.n267 B.n266 585
R1548 B.n268 B.n213 585
R1549 B.n270 B.n269 585
R1550 B.n271 B.n212 585
R1551 B.n273 B.n272 585
R1552 B.n274 B.n211 585
R1553 B.n276 B.n275 585
R1554 B.n277 B.n210 585
R1555 B.n279 B.n278 585
R1556 B.n280 B.n209 585
R1557 B.n282 B.n281 585
R1558 B.n283 B.n208 585
R1559 B.n285 B.n284 585
R1560 B.n286 B.n207 585
R1561 B.n288 B.n287 585
R1562 B.n289 B.n206 585
R1563 B.n291 B.n290 585
R1564 B.n292 B.n205 585
R1565 B.n294 B.n293 585
R1566 B.n295 B.n204 585
R1567 B.n297 B.n296 585
R1568 B.n298 B.n203 585
R1569 B.n300 B.n299 585
R1570 B.n301 B.n202 585
R1571 B.n303 B.n302 585
R1572 B.n304 B.n201 585
R1573 B.n306 B.n305 585
R1574 B.n307 B.n200 585
R1575 B.n309 B.n308 585
R1576 B.n310 B.n199 585
R1577 B.n312 B.n311 585
R1578 B.n313 B.n198 585
R1579 B.n315 B.n314 585
R1580 B.n316 B.n197 585
R1581 B.n318 B.n317 585
R1582 B.n319 B.n318 497.305
R1583 B.n462 B.n147 497.305
R1584 B.n653 B.n652 497.305
R1585 B.n796 B.n33 497.305
R1586 B.n396 B.t1 438.366
R1587 B.n62 B.t11 438.366
R1588 B.n174 B.t4 438.366
R1589 B.n54 B.t8 438.366
R1590 B.n397 B.t2 378.44
R1591 B.n63 B.t10 378.44
R1592 B.n175 B.t5 378.44
R1593 B.n55 B.t7 378.44
R1594 B.n174 B.t3 314.368
R1595 B.n396 B.t0 314.368
R1596 B.n62 B.t9 314.368
R1597 B.n54 B.t6 314.368
R1598 B.n889 B.n888 256.663
R1599 B.n888 B.n887 235.042
R1600 B.n888 B.n2 235.042
R1601 B.n320 B.n319 163.367
R1602 B.n320 B.n195 163.367
R1603 B.n324 B.n195 163.367
R1604 B.n325 B.n324 163.367
R1605 B.n326 B.n325 163.367
R1606 B.n326 B.n193 163.367
R1607 B.n330 B.n193 163.367
R1608 B.n331 B.n330 163.367
R1609 B.n332 B.n331 163.367
R1610 B.n332 B.n191 163.367
R1611 B.n336 B.n191 163.367
R1612 B.n337 B.n336 163.367
R1613 B.n338 B.n337 163.367
R1614 B.n338 B.n189 163.367
R1615 B.n342 B.n189 163.367
R1616 B.n343 B.n342 163.367
R1617 B.n344 B.n343 163.367
R1618 B.n344 B.n187 163.367
R1619 B.n348 B.n187 163.367
R1620 B.n349 B.n348 163.367
R1621 B.n350 B.n349 163.367
R1622 B.n350 B.n185 163.367
R1623 B.n354 B.n185 163.367
R1624 B.n355 B.n354 163.367
R1625 B.n356 B.n355 163.367
R1626 B.n356 B.n183 163.367
R1627 B.n360 B.n183 163.367
R1628 B.n361 B.n360 163.367
R1629 B.n362 B.n361 163.367
R1630 B.n362 B.n181 163.367
R1631 B.n366 B.n181 163.367
R1632 B.n367 B.n366 163.367
R1633 B.n368 B.n367 163.367
R1634 B.n368 B.n179 163.367
R1635 B.n372 B.n179 163.367
R1636 B.n373 B.n372 163.367
R1637 B.n374 B.n373 163.367
R1638 B.n374 B.n177 163.367
R1639 B.n378 B.n177 163.367
R1640 B.n379 B.n378 163.367
R1641 B.n380 B.n379 163.367
R1642 B.n380 B.n173 163.367
R1643 B.n385 B.n173 163.367
R1644 B.n386 B.n385 163.367
R1645 B.n387 B.n386 163.367
R1646 B.n387 B.n171 163.367
R1647 B.n391 B.n171 163.367
R1648 B.n392 B.n391 163.367
R1649 B.n393 B.n392 163.367
R1650 B.n393 B.n169 163.367
R1651 B.n400 B.n169 163.367
R1652 B.n401 B.n400 163.367
R1653 B.n402 B.n401 163.367
R1654 B.n402 B.n167 163.367
R1655 B.n406 B.n167 163.367
R1656 B.n407 B.n406 163.367
R1657 B.n408 B.n407 163.367
R1658 B.n408 B.n165 163.367
R1659 B.n412 B.n165 163.367
R1660 B.n413 B.n412 163.367
R1661 B.n414 B.n413 163.367
R1662 B.n414 B.n163 163.367
R1663 B.n418 B.n163 163.367
R1664 B.n419 B.n418 163.367
R1665 B.n420 B.n419 163.367
R1666 B.n420 B.n161 163.367
R1667 B.n424 B.n161 163.367
R1668 B.n425 B.n424 163.367
R1669 B.n426 B.n425 163.367
R1670 B.n426 B.n159 163.367
R1671 B.n430 B.n159 163.367
R1672 B.n431 B.n430 163.367
R1673 B.n432 B.n431 163.367
R1674 B.n432 B.n157 163.367
R1675 B.n436 B.n157 163.367
R1676 B.n437 B.n436 163.367
R1677 B.n438 B.n437 163.367
R1678 B.n438 B.n155 163.367
R1679 B.n442 B.n155 163.367
R1680 B.n443 B.n442 163.367
R1681 B.n444 B.n443 163.367
R1682 B.n444 B.n153 163.367
R1683 B.n448 B.n153 163.367
R1684 B.n449 B.n448 163.367
R1685 B.n450 B.n449 163.367
R1686 B.n450 B.n151 163.367
R1687 B.n454 B.n151 163.367
R1688 B.n455 B.n454 163.367
R1689 B.n456 B.n455 163.367
R1690 B.n456 B.n149 163.367
R1691 B.n460 B.n149 163.367
R1692 B.n461 B.n460 163.367
R1693 B.n462 B.n461 163.367
R1694 B.n652 B.n85 163.367
R1695 B.n648 B.n85 163.367
R1696 B.n648 B.n647 163.367
R1697 B.n647 B.n646 163.367
R1698 B.n646 B.n87 163.367
R1699 B.n642 B.n87 163.367
R1700 B.n642 B.n641 163.367
R1701 B.n641 B.n640 163.367
R1702 B.n640 B.n89 163.367
R1703 B.n636 B.n89 163.367
R1704 B.n636 B.n635 163.367
R1705 B.n635 B.n634 163.367
R1706 B.n634 B.n91 163.367
R1707 B.n630 B.n91 163.367
R1708 B.n630 B.n629 163.367
R1709 B.n629 B.n628 163.367
R1710 B.n628 B.n93 163.367
R1711 B.n624 B.n93 163.367
R1712 B.n624 B.n623 163.367
R1713 B.n623 B.n622 163.367
R1714 B.n622 B.n95 163.367
R1715 B.n618 B.n95 163.367
R1716 B.n618 B.n617 163.367
R1717 B.n617 B.n616 163.367
R1718 B.n616 B.n97 163.367
R1719 B.n612 B.n97 163.367
R1720 B.n612 B.n611 163.367
R1721 B.n611 B.n610 163.367
R1722 B.n610 B.n99 163.367
R1723 B.n606 B.n99 163.367
R1724 B.n606 B.n605 163.367
R1725 B.n605 B.n604 163.367
R1726 B.n604 B.n101 163.367
R1727 B.n600 B.n101 163.367
R1728 B.n600 B.n599 163.367
R1729 B.n599 B.n598 163.367
R1730 B.n598 B.n103 163.367
R1731 B.n594 B.n103 163.367
R1732 B.n594 B.n593 163.367
R1733 B.n593 B.n592 163.367
R1734 B.n592 B.n105 163.367
R1735 B.n588 B.n105 163.367
R1736 B.n588 B.n587 163.367
R1737 B.n587 B.n586 163.367
R1738 B.n586 B.n107 163.367
R1739 B.n582 B.n107 163.367
R1740 B.n582 B.n581 163.367
R1741 B.n581 B.n580 163.367
R1742 B.n580 B.n109 163.367
R1743 B.n576 B.n109 163.367
R1744 B.n576 B.n575 163.367
R1745 B.n575 B.n574 163.367
R1746 B.n574 B.n111 163.367
R1747 B.n570 B.n111 163.367
R1748 B.n570 B.n569 163.367
R1749 B.n569 B.n568 163.367
R1750 B.n568 B.n113 163.367
R1751 B.n564 B.n113 163.367
R1752 B.n564 B.n563 163.367
R1753 B.n563 B.n562 163.367
R1754 B.n562 B.n115 163.367
R1755 B.n558 B.n115 163.367
R1756 B.n558 B.n557 163.367
R1757 B.n557 B.n556 163.367
R1758 B.n556 B.n117 163.367
R1759 B.n552 B.n117 163.367
R1760 B.n552 B.n551 163.367
R1761 B.n551 B.n550 163.367
R1762 B.n550 B.n119 163.367
R1763 B.n546 B.n119 163.367
R1764 B.n546 B.n545 163.367
R1765 B.n545 B.n544 163.367
R1766 B.n544 B.n121 163.367
R1767 B.n540 B.n121 163.367
R1768 B.n540 B.n539 163.367
R1769 B.n539 B.n538 163.367
R1770 B.n538 B.n123 163.367
R1771 B.n534 B.n123 163.367
R1772 B.n534 B.n533 163.367
R1773 B.n533 B.n532 163.367
R1774 B.n532 B.n125 163.367
R1775 B.n528 B.n125 163.367
R1776 B.n528 B.n527 163.367
R1777 B.n527 B.n526 163.367
R1778 B.n526 B.n127 163.367
R1779 B.n522 B.n127 163.367
R1780 B.n522 B.n521 163.367
R1781 B.n521 B.n520 163.367
R1782 B.n520 B.n129 163.367
R1783 B.n516 B.n129 163.367
R1784 B.n516 B.n515 163.367
R1785 B.n515 B.n514 163.367
R1786 B.n514 B.n131 163.367
R1787 B.n510 B.n131 163.367
R1788 B.n510 B.n509 163.367
R1789 B.n509 B.n508 163.367
R1790 B.n508 B.n133 163.367
R1791 B.n504 B.n133 163.367
R1792 B.n504 B.n503 163.367
R1793 B.n503 B.n502 163.367
R1794 B.n502 B.n135 163.367
R1795 B.n498 B.n135 163.367
R1796 B.n498 B.n497 163.367
R1797 B.n497 B.n496 163.367
R1798 B.n496 B.n137 163.367
R1799 B.n492 B.n137 163.367
R1800 B.n492 B.n491 163.367
R1801 B.n491 B.n490 163.367
R1802 B.n490 B.n139 163.367
R1803 B.n486 B.n139 163.367
R1804 B.n486 B.n485 163.367
R1805 B.n485 B.n484 163.367
R1806 B.n484 B.n141 163.367
R1807 B.n480 B.n141 163.367
R1808 B.n480 B.n479 163.367
R1809 B.n479 B.n478 163.367
R1810 B.n478 B.n143 163.367
R1811 B.n474 B.n143 163.367
R1812 B.n474 B.n473 163.367
R1813 B.n473 B.n472 163.367
R1814 B.n472 B.n145 163.367
R1815 B.n468 B.n145 163.367
R1816 B.n468 B.n467 163.367
R1817 B.n467 B.n466 163.367
R1818 B.n466 B.n147 163.367
R1819 B.n792 B.n33 163.367
R1820 B.n792 B.n791 163.367
R1821 B.n791 B.n790 163.367
R1822 B.n790 B.n35 163.367
R1823 B.n786 B.n35 163.367
R1824 B.n786 B.n785 163.367
R1825 B.n785 B.n784 163.367
R1826 B.n784 B.n37 163.367
R1827 B.n780 B.n37 163.367
R1828 B.n780 B.n779 163.367
R1829 B.n779 B.n778 163.367
R1830 B.n778 B.n39 163.367
R1831 B.n774 B.n39 163.367
R1832 B.n774 B.n773 163.367
R1833 B.n773 B.n772 163.367
R1834 B.n772 B.n41 163.367
R1835 B.n768 B.n41 163.367
R1836 B.n768 B.n767 163.367
R1837 B.n767 B.n766 163.367
R1838 B.n766 B.n43 163.367
R1839 B.n762 B.n43 163.367
R1840 B.n762 B.n761 163.367
R1841 B.n761 B.n760 163.367
R1842 B.n760 B.n45 163.367
R1843 B.n756 B.n45 163.367
R1844 B.n756 B.n755 163.367
R1845 B.n755 B.n754 163.367
R1846 B.n754 B.n47 163.367
R1847 B.n750 B.n47 163.367
R1848 B.n750 B.n749 163.367
R1849 B.n749 B.n748 163.367
R1850 B.n748 B.n49 163.367
R1851 B.n744 B.n49 163.367
R1852 B.n744 B.n743 163.367
R1853 B.n743 B.n742 163.367
R1854 B.n742 B.n51 163.367
R1855 B.n738 B.n51 163.367
R1856 B.n738 B.n737 163.367
R1857 B.n737 B.n736 163.367
R1858 B.n736 B.n53 163.367
R1859 B.n732 B.n53 163.367
R1860 B.n732 B.n731 163.367
R1861 B.n731 B.n57 163.367
R1862 B.n727 B.n57 163.367
R1863 B.n727 B.n726 163.367
R1864 B.n726 B.n725 163.367
R1865 B.n725 B.n59 163.367
R1866 B.n721 B.n59 163.367
R1867 B.n721 B.n720 163.367
R1868 B.n720 B.n719 163.367
R1869 B.n719 B.n61 163.367
R1870 B.n714 B.n61 163.367
R1871 B.n714 B.n713 163.367
R1872 B.n713 B.n712 163.367
R1873 B.n712 B.n65 163.367
R1874 B.n708 B.n65 163.367
R1875 B.n708 B.n707 163.367
R1876 B.n707 B.n706 163.367
R1877 B.n706 B.n67 163.367
R1878 B.n702 B.n67 163.367
R1879 B.n702 B.n701 163.367
R1880 B.n701 B.n700 163.367
R1881 B.n700 B.n69 163.367
R1882 B.n696 B.n69 163.367
R1883 B.n696 B.n695 163.367
R1884 B.n695 B.n694 163.367
R1885 B.n694 B.n71 163.367
R1886 B.n690 B.n71 163.367
R1887 B.n690 B.n689 163.367
R1888 B.n689 B.n688 163.367
R1889 B.n688 B.n73 163.367
R1890 B.n684 B.n73 163.367
R1891 B.n684 B.n683 163.367
R1892 B.n683 B.n682 163.367
R1893 B.n682 B.n75 163.367
R1894 B.n678 B.n75 163.367
R1895 B.n678 B.n677 163.367
R1896 B.n677 B.n676 163.367
R1897 B.n676 B.n77 163.367
R1898 B.n672 B.n77 163.367
R1899 B.n672 B.n671 163.367
R1900 B.n671 B.n670 163.367
R1901 B.n670 B.n79 163.367
R1902 B.n666 B.n79 163.367
R1903 B.n666 B.n665 163.367
R1904 B.n665 B.n664 163.367
R1905 B.n664 B.n81 163.367
R1906 B.n660 B.n81 163.367
R1907 B.n660 B.n659 163.367
R1908 B.n659 B.n658 163.367
R1909 B.n658 B.n83 163.367
R1910 B.n654 B.n83 163.367
R1911 B.n654 B.n653 163.367
R1912 B.n797 B.n796 163.367
R1913 B.n798 B.n797 163.367
R1914 B.n798 B.n31 163.367
R1915 B.n802 B.n31 163.367
R1916 B.n803 B.n802 163.367
R1917 B.n804 B.n803 163.367
R1918 B.n804 B.n29 163.367
R1919 B.n808 B.n29 163.367
R1920 B.n809 B.n808 163.367
R1921 B.n810 B.n809 163.367
R1922 B.n810 B.n27 163.367
R1923 B.n814 B.n27 163.367
R1924 B.n815 B.n814 163.367
R1925 B.n816 B.n815 163.367
R1926 B.n816 B.n25 163.367
R1927 B.n820 B.n25 163.367
R1928 B.n821 B.n820 163.367
R1929 B.n822 B.n821 163.367
R1930 B.n822 B.n23 163.367
R1931 B.n826 B.n23 163.367
R1932 B.n827 B.n826 163.367
R1933 B.n828 B.n827 163.367
R1934 B.n828 B.n21 163.367
R1935 B.n832 B.n21 163.367
R1936 B.n833 B.n832 163.367
R1937 B.n834 B.n833 163.367
R1938 B.n834 B.n19 163.367
R1939 B.n838 B.n19 163.367
R1940 B.n839 B.n838 163.367
R1941 B.n840 B.n839 163.367
R1942 B.n840 B.n17 163.367
R1943 B.n844 B.n17 163.367
R1944 B.n845 B.n844 163.367
R1945 B.n846 B.n845 163.367
R1946 B.n846 B.n15 163.367
R1947 B.n850 B.n15 163.367
R1948 B.n851 B.n850 163.367
R1949 B.n852 B.n851 163.367
R1950 B.n852 B.n13 163.367
R1951 B.n856 B.n13 163.367
R1952 B.n857 B.n856 163.367
R1953 B.n858 B.n857 163.367
R1954 B.n858 B.n11 163.367
R1955 B.n862 B.n11 163.367
R1956 B.n863 B.n862 163.367
R1957 B.n864 B.n863 163.367
R1958 B.n864 B.n9 163.367
R1959 B.n868 B.n9 163.367
R1960 B.n869 B.n868 163.367
R1961 B.n870 B.n869 163.367
R1962 B.n870 B.n7 163.367
R1963 B.n874 B.n7 163.367
R1964 B.n875 B.n874 163.367
R1965 B.n876 B.n875 163.367
R1966 B.n876 B.n5 163.367
R1967 B.n880 B.n5 163.367
R1968 B.n881 B.n880 163.367
R1969 B.n882 B.n881 163.367
R1970 B.n882 B.n3 163.367
R1971 B.n886 B.n3 163.367
R1972 B.n887 B.n886 163.367
R1973 B.n228 B.n2 163.367
R1974 B.n229 B.n228 163.367
R1975 B.n230 B.n229 163.367
R1976 B.n230 B.n225 163.367
R1977 B.n234 B.n225 163.367
R1978 B.n235 B.n234 163.367
R1979 B.n236 B.n235 163.367
R1980 B.n236 B.n223 163.367
R1981 B.n240 B.n223 163.367
R1982 B.n241 B.n240 163.367
R1983 B.n242 B.n241 163.367
R1984 B.n242 B.n221 163.367
R1985 B.n246 B.n221 163.367
R1986 B.n247 B.n246 163.367
R1987 B.n248 B.n247 163.367
R1988 B.n248 B.n219 163.367
R1989 B.n252 B.n219 163.367
R1990 B.n253 B.n252 163.367
R1991 B.n254 B.n253 163.367
R1992 B.n254 B.n217 163.367
R1993 B.n258 B.n217 163.367
R1994 B.n259 B.n258 163.367
R1995 B.n260 B.n259 163.367
R1996 B.n260 B.n215 163.367
R1997 B.n264 B.n215 163.367
R1998 B.n265 B.n264 163.367
R1999 B.n266 B.n265 163.367
R2000 B.n266 B.n213 163.367
R2001 B.n270 B.n213 163.367
R2002 B.n271 B.n270 163.367
R2003 B.n272 B.n271 163.367
R2004 B.n272 B.n211 163.367
R2005 B.n276 B.n211 163.367
R2006 B.n277 B.n276 163.367
R2007 B.n278 B.n277 163.367
R2008 B.n278 B.n209 163.367
R2009 B.n282 B.n209 163.367
R2010 B.n283 B.n282 163.367
R2011 B.n284 B.n283 163.367
R2012 B.n284 B.n207 163.367
R2013 B.n288 B.n207 163.367
R2014 B.n289 B.n288 163.367
R2015 B.n290 B.n289 163.367
R2016 B.n290 B.n205 163.367
R2017 B.n294 B.n205 163.367
R2018 B.n295 B.n294 163.367
R2019 B.n296 B.n295 163.367
R2020 B.n296 B.n203 163.367
R2021 B.n300 B.n203 163.367
R2022 B.n301 B.n300 163.367
R2023 B.n302 B.n301 163.367
R2024 B.n302 B.n201 163.367
R2025 B.n306 B.n201 163.367
R2026 B.n307 B.n306 163.367
R2027 B.n308 B.n307 163.367
R2028 B.n308 B.n199 163.367
R2029 B.n312 B.n199 163.367
R2030 B.n313 B.n312 163.367
R2031 B.n314 B.n313 163.367
R2032 B.n314 B.n197 163.367
R2033 B.n318 B.n197 163.367
R2034 B.n175 B.n174 59.9278
R2035 B.n397 B.n396 59.9278
R2036 B.n63 B.n62 59.9278
R2037 B.n55 B.n54 59.9278
R2038 B.n382 B.n175 59.5399
R2039 B.n398 B.n397 59.5399
R2040 B.n716 B.n63 59.5399
R2041 B.n56 B.n55 59.5399
R2042 B.n795 B.n794 32.3127
R2043 B.n651 B.n84 32.3127
R2044 B.n464 B.n463 32.3127
R2045 B.n317 B.n196 32.3127
R2046 B B.n889 18.0485
R2047 B.n795 B.n32 10.6151
R2048 B.n799 B.n32 10.6151
R2049 B.n800 B.n799 10.6151
R2050 B.n801 B.n800 10.6151
R2051 B.n801 B.n30 10.6151
R2052 B.n805 B.n30 10.6151
R2053 B.n806 B.n805 10.6151
R2054 B.n807 B.n806 10.6151
R2055 B.n807 B.n28 10.6151
R2056 B.n811 B.n28 10.6151
R2057 B.n812 B.n811 10.6151
R2058 B.n813 B.n812 10.6151
R2059 B.n813 B.n26 10.6151
R2060 B.n817 B.n26 10.6151
R2061 B.n818 B.n817 10.6151
R2062 B.n819 B.n818 10.6151
R2063 B.n819 B.n24 10.6151
R2064 B.n823 B.n24 10.6151
R2065 B.n824 B.n823 10.6151
R2066 B.n825 B.n824 10.6151
R2067 B.n825 B.n22 10.6151
R2068 B.n829 B.n22 10.6151
R2069 B.n830 B.n829 10.6151
R2070 B.n831 B.n830 10.6151
R2071 B.n831 B.n20 10.6151
R2072 B.n835 B.n20 10.6151
R2073 B.n836 B.n835 10.6151
R2074 B.n837 B.n836 10.6151
R2075 B.n837 B.n18 10.6151
R2076 B.n841 B.n18 10.6151
R2077 B.n842 B.n841 10.6151
R2078 B.n843 B.n842 10.6151
R2079 B.n843 B.n16 10.6151
R2080 B.n847 B.n16 10.6151
R2081 B.n848 B.n847 10.6151
R2082 B.n849 B.n848 10.6151
R2083 B.n849 B.n14 10.6151
R2084 B.n853 B.n14 10.6151
R2085 B.n854 B.n853 10.6151
R2086 B.n855 B.n854 10.6151
R2087 B.n855 B.n12 10.6151
R2088 B.n859 B.n12 10.6151
R2089 B.n860 B.n859 10.6151
R2090 B.n861 B.n860 10.6151
R2091 B.n861 B.n10 10.6151
R2092 B.n865 B.n10 10.6151
R2093 B.n866 B.n865 10.6151
R2094 B.n867 B.n866 10.6151
R2095 B.n867 B.n8 10.6151
R2096 B.n871 B.n8 10.6151
R2097 B.n872 B.n871 10.6151
R2098 B.n873 B.n872 10.6151
R2099 B.n873 B.n6 10.6151
R2100 B.n877 B.n6 10.6151
R2101 B.n878 B.n877 10.6151
R2102 B.n879 B.n878 10.6151
R2103 B.n879 B.n4 10.6151
R2104 B.n883 B.n4 10.6151
R2105 B.n884 B.n883 10.6151
R2106 B.n885 B.n884 10.6151
R2107 B.n885 B.n0 10.6151
R2108 B.n794 B.n793 10.6151
R2109 B.n793 B.n34 10.6151
R2110 B.n789 B.n34 10.6151
R2111 B.n789 B.n788 10.6151
R2112 B.n788 B.n787 10.6151
R2113 B.n787 B.n36 10.6151
R2114 B.n783 B.n36 10.6151
R2115 B.n783 B.n782 10.6151
R2116 B.n782 B.n781 10.6151
R2117 B.n781 B.n38 10.6151
R2118 B.n777 B.n38 10.6151
R2119 B.n777 B.n776 10.6151
R2120 B.n776 B.n775 10.6151
R2121 B.n775 B.n40 10.6151
R2122 B.n771 B.n40 10.6151
R2123 B.n771 B.n770 10.6151
R2124 B.n770 B.n769 10.6151
R2125 B.n769 B.n42 10.6151
R2126 B.n765 B.n42 10.6151
R2127 B.n765 B.n764 10.6151
R2128 B.n764 B.n763 10.6151
R2129 B.n763 B.n44 10.6151
R2130 B.n759 B.n44 10.6151
R2131 B.n759 B.n758 10.6151
R2132 B.n758 B.n757 10.6151
R2133 B.n757 B.n46 10.6151
R2134 B.n753 B.n46 10.6151
R2135 B.n753 B.n752 10.6151
R2136 B.n752 B.n751 10.6151
R2137 B.n751 B.n48 10.6151
R2138 B.n747 B.n48 10.6151
R2139 B.n747 B.n746 10.6151
R2140 B.n746 B.n745 10.6151
R2141 B.n745 B.n50 10.6151
R2142 B.n741 B.n50 10.6151
R2143 B.n741 B.n740 10.6151
R2144 B.n740 B.n739 10.6151
R2145 B.n739 B.n52 10.6151
R2146 B.n735 B.n52 10.6151
R2147 B.n735 B.n734 10.6151
R2148 B.n734 B.n733 10.6151
R2149 B.n730 B.n729 10.6151
R2150 B.n729 B.n728 10.6151
R2151 B.n728 B.n58 10.6151
R2152 B.n724 B.n58 10.6151
R2153 B.n724 B.n723 10.6151
R2154 B.n723 B.n722 10.6151
R2155 B.n722 B.n60 10.6151
R2156 B.n718 B.n60 10.6151
R2157 B.n718 B.n717 10.6151
R2158 B.n715 B.n64 10.6151
R2159 B.n711 B.n64 10.6151
R2160 B.n711 B.n710 10.6151
R2161 B.n710 B.n709 10.6151
R2162 B.n709 B.n66 10.6151
R2163 B.n705 B.n66 10.6151
R2164 B.n705 B.n704 10.6151
R2165 B.n704 B.n703 10.6151
R2166 B.n703 B.n68 10.6151
R2167 B.n699 B.n68 10.6151
R2168 B.n699 B.n698 10.6151
R2169 B.n698 B.n697 10.6151
R2170 B.n697 B.n70 10.6151
R2171 B.n693 B.n70 10.6151
R2172 B.n693 B.n692 10.6151
R2173 B.n692 B.n691 10.6151
R2174 B.n691 B.n72 10.6151
R2175 B.n687 B.n72 10.6151
R2176 B.n687 B.n686 10.6151
R2177 B.n686 B.n685 10.6151
R2178 B.n685 B.n74 10.6151
R2179 B.n681 B.n74 10.6151
R2180 B.n681 B.n680 10.6151
R2181 B.n680 B.n679 10.6151
R2182 B.n679 B.n76 10.6151
R2183 B.n675 B.n76 10.6151
R2184 B.n675 B.n674 10.6151
R2185 B.n674 B.n673 10.6151
R2186 B.n673 B.n78 10.6151
R2187 B.n669 B.n78 10.6151
R2188 B.n669 B.n668 10.6151
R2189 B.n668 B.n667 10.6151
R2190 B.n667 B.n80 10.6151
R2191 B.n663 B.n80 10.6151
R2192 B.n663 B.n662 10.6151
R2193 B.n662 B.n661 10.6151
R2194 B.n661 B.n82 10.6151
R2195 B.n657 B.n82 10.6151
R2196 B.n657 B.n656 10.6151
R2197 B.n656 B.n655 10.6151
R2198 B.n655 B.n84 10.6151
R2199 B.n651 B.n650 10.6151
R2200 B.n650 B.n649 10.6151
R2201 B.n649 B.n86 10.6151
R2202 B.n645 B.n86 10.6151
R2203 B.n645 B.n644 10.6151
R2204 B.n644 B.n643 10.6151
R2205 B.n643 B.n88 10.6151
R2206 B.n639 B.n88 10.6151
R2207 B.n639 B.n638 10.6151
R2208 B.n638 B.n637 10.6151
R2209 B.n637 B.n90 10.6151
R2210 B.n633 B.n90 10.6151
R2211 B.n633 B.n632 10.6151
R2212 B.n632 B.n631 10.6151
R2213 B.n631 B.n92 10.6151
R2214 B.n627 B.n92 10.6151
R2215 B.n627 B.n626 10.6151
R2216 B.n626 B.n625 10.6151
R2217 B.n625 B.n94 10.6151
R2218 B.n621 B.n94 10.6151
R2219 B.n621 B.n620 10.6151
R2220 B.n620 B.n619 10.6151
R2221 B.n619 B.n96 10.6151
R2222 B.n615 B.n96 10.6151
R2223 B.n615 B.n614 10.6151
R2224 B.n614 B.n613 10.6151
R2225 B.n613 B.n98 10.6151
R2226 B.n609 B.n98 10.6151
R2227 B.n609 B.n608 10.6151
R2228 B.n608 B.n607 10.6151
R2229 B.n607 B.n100 10.6151
R2230 B.n603 B.n100 10.6151
R2231 B.n603 B.n602 10.6151
R2232 B.n602 B.n601 10.6151
R2233 B.n601 B.n102 10.6151
R2234 B.n597 B.n102 10.6151
R2235 B.n597 B.n596 10.6151
R2236 B.n596 B.n595 10.6151
R2237 B.n595 B.n104 10.6151
R2238 B.n591 B.n104 10.6151
R2239 B.n591 B.n590 10.6151
R2240 B.n590 B.n589 10.6151
R2241 B.n589 B.n106 10.6151
R2242 B.n585 B.n106 10.6151
R2243 B.n585 B.n584 10.6151
R2244 B.n584 B.n583 10.6151
R2245 B.n583 B.n108 10.6151
R2246 B.n579 B.n108 10.6151
R2247 B.n579 B.n578 10.6151
R2248 B.n578 B.n577 10.6151
R2249 B.n577 B.n110 10.6151
R2250 B.n573 B.n110 10.6151
R2251 B.n573 B.n572 10.6151
R2252 B.n572 B.n571 10.6151
R2253 B.n571 B.n112 10.6151
R2254 B.n567 B.n112 10.6151
R2255 B.n567 B.n566 10.6151
R2256 B.n566 B.n565 10.6151
R2257 B.n565 B.n114 10.6151
R2258 B.n561 B.n114 10.6151
R2259 B.n561 B.n560 10.6151
R2260 B.n560 B.n559 10.6151
R2261 B.n559 B.n116 10.6151
R2262 B.n555 B.n116 10.6151
R2263 B.n555 B.n554 10.6151
R2264 B.n554 B.n553 10.6151
R2265 B.n553 B.n118 10.6151
R2266 B.n549 B.n118 10.6151
R2267 B.n549 B.n548 10.6151
R2268 B.n548 B.n547 10.6151
R2269 B.n547 B.n120 10.6151
R2270 B.n543 B.n120 10.6151
R2271 B.n543 B.n542 10.6151
R2272 B.n542 B.n541 10.6151
R2273 B.n541 B.n122 10.6151
R2274 B.n537 B.n122 10.6151
R2275 B.n537 B.n536 10.6151
R2276 B.n536 B.n535 10.6151
R2277 B.n535 B.n124 10.6151
R2278 B.n531 B.n124 10.6151
R2279 B.n531 B.n530 10.6151
R2280 B.n530 B.n529 10.6151
R2281 B.n529 B.n126 10.6151
R2282 B.n525 B.n126 10.6151
R2283 B.n525 B.n524 10.6151
R2284 B.n524 B.n523 10.6151
R2285 B.n523 B.n128 10.6151
R2286 B.n519 B.n128 10.6151
R2287 B.n519 B.n518 10.6151
R2288 B.n518 B.n517 10.6151
R2289 B.n517 B.n130 10.6151
R2290 B.n513 B.n130 10.6151
R2291 B.n513 B.n512 10.6151
R2292 B.n512 B.n511 10.6151
R2293 B.n511 B.n132 10.6151
R2294 B.n507 B.n132 10.6151
R2295 B.n507 B.n506 10.6151
R2296 B.n506 B.n505 10.6151
R2297 B.n505 B.n134 10.6151
R2298 B.n501 B.n134 10.6151
R2299 B.n501 B.n500 10.6151
R2300 B.n500 B.n499 10.6151
R2301 B.n499 B.n136 10.6151
R2302 B.n495 B.n136 10.6151
R2303 B.n495 B.n494 10.6151
R2304 B.n494 B.n493 10.6151
R2305 B.n493 B.n138 10.6151
R2306 B.n489 B.n138 10.6151
R2307 B.n489 B.n488 10.6151
R2308 B.n488 B.n487 10.6151
R2309 B.n487 B.n140 10.6151
R2310 B.n483 B.n140 10.6151
R2311 B.n483 B.n482 10.6151
R2312 B.n482 B.n481 10.6151
R2313 B.n481 B.n142 10.6151
R2314 B.n477 B.n142 10.6151
R2315 B.n477 B.n476 10.6151
R2316 B.n476 B.n475 10.6151
R2317 B.n475 B.n144 10.6151
R2318 B.n471 B.n144 10.6151
R2319 B.n471 B.n470 10.6151
R2320 B.n470 B.n469 10.6151
R2321 B.n469 B.n146 10.6151
R2322 B.n465 B.n146 10.6151
R2323 B.n465 B.n464 10.6151
R2324 B.n227 B.n1 10.6151
R2325 B.n227 B.n226 10.6151
R2326 B.n231 B.n226 10.6151
R2327 B.n232 B.n231 10.6151
R2328 B.n233 B.n232 10.6151
R2329 B.n233 B.n224 10.6151
R2330 B.n237 B.n224 10.6151
R2331 B.n238 B.n237 10.6151
R2332 B.n239 B.n238 10.6151
R2333 B.n239 B.n222 10.6151
R2334 B.n243 B.n222 10.6151
R2335 B.n244 B.n243 10.6151
R2336 B.n245 B.n244 10.6151
R2337 B.n245 B.n220 10.6151
R2338 B.n249 B.n220 10.6151
R2339 B.n250 B.n249 10.6151
R2340 B.n251 B.n250 10.6151
R2341 B.n251 B.n218 10.6151
R2342 B.n255 B.n218 10.6151
R2343 B.n256 B.n255 10.6151
R2344 B.n257 B.n256 10.6151
R2345 B.n257 B.n216 10.6151
R2346 B.n261 B.n216 10.6151
R2347 B.n262 B.n261 10.6151
R2348 B.n263 B.n262 10.6151
R2349 B.n263 B.n214 10.6151
R2350 B.n267 B.n214 10.6151
R2351 B.n268 B.n267 10.6151
R2352 B.n269 B.n268 10.6151
R2353 B.n269 B.n212 10.6151
R2354 B.n273 B.n212 10.6151
R2355 B.n274 B.n273 10.6151
R2356 B.n275 B.n274 10.6151
R2357 B.n275 B.n210 10.6151
R2358 B.n279 B.n210 10.6151
R2359 B.n280 B.n279 10.6151
R2360 B.n281 B.n280 10.6151
R2361 B.n281 B.n208 10.6151
R2362 B.n285 B.n208 10.6151
R2363 B.n286 B.n285 10.6151
R2364 B.n287 B.n286 10.6151
R2365 B.n287 B.n206 10.6151
R2366 B.n291 B.n206 10.6151
R2367 B.n292 B.n291 10.6151
R2368 B.n293 B.n292 10.6151
R2369 B.n293 B.n204 10.6151
R2370 B.n297 B.n204 10.6151
R2371 B.n298 B.n297 10.6151
R2372 B.n299 B.n298 10.6151
R2373 B.n299 B.n202 10.6151
R2374 B.n303 B.n202 10.6151
R2375 B.n304 B.n303 10.6151
R2376 B.n305 B.n304 10.6151
R2377 B.n305 B.n200 10.6151
R2378 B.n309 B.n200 10.6151
R2379 B.n310 B.n309 10.6151
R2380 B.n311 B.n310 10.6151
R2381 B.n311 B.n198 10.6151
R2382 B.n315 B.n198 10.6151
R2383 B.n316 B.n315 10.6151
R2384 B.n317 B.n316 10.6151
R2385 B.n321 B.n196 10.6151
R2386 B.n322 B.n321 10.6151
R2387 B.n323 B.n322 10.6151
R2388 B.n323 B.n194 10.6151
R2389 B.n327 B.n194 10.6151
R2390 B.n328 B.n327 10.6151
R2391 B.n329 B.n328 10.6151
R2392 B.n329 B.n192 10.6151
R2393 B.n333 B.n192 10.6151
R2394 B.n334 B.n333 10.6151
R2395 B.n335 B.n334 10.6151
R2396 B.n335 B.n190 10.6151
R2397 B.n339 B.n190 10.6151
R2398 B.n340 B.n339 10.6151
R2399 B.n341 B.n340 10.6151
R2400 B.n341 B.n188 10.6151
R2401 B.n345 B.n188 10.6151
R2402 B.n346 B.n345 10.6151
R2403 B.n347 B.n346 10.6151
R2404 B.n347 B.n186 10.6151
R2405 B.n351 B.n186 10.6151
R2406 B.n352 B.n351 10.6151
R2407 B.n353 B.n352 10.6151
R2408 B.n353 B.n184 10.6151
R2409 B.n357 B.n184 10.6151
R2410 B.n358 B.n357 10.6151
R2411 B.n359 B.n358 10.6151
R2412 B.n359 B.n182 10.6151
R2413 B.n363 B.n182 10.6151
R2414 B.n364 B.n363 10.6151
R2415 B.n365 B.n364 10.6151
R2416 B.n365 B.n180 10.6151
R2417 B.n369 B.n180 10.6151
R2418 B.n370 B.n369 10.6151
R2419 B.n371 B.n370 10.6151
R2420 B.n371 B.n178 10.6151
R2421 B.n375 B.n178 10.6151
R2422 B.n376 B.n375 10.6151
R2423 B.n377 B.n376 10.6151
R2424 B.n377 B.n176 10.6151
R2425 B.n381 B.n176 10.6151
R2426 B.n384 B.n383 10.6151
R2427 B.n384 B.n172 10.6151
R2428 B.n388 B.n172 10.6151
R2429 B.n389 B.n388 10.6151
R2430 B.n390 B.n389 10.6151
R2431 B.n390 B.n170 10.6151
R2432 B.n394 B.n170 10.6151
R2433 B.n395 B.n394 10.6151
R2434 B.n399 B.n395 10.6151
R2435 B.n403 B.n168 10.6151
R2436 B.n404 B.n403 10.6151
R2437 B.n405 B.n404 10.6151
R2438 B.n405 B.n166 10.6151
R2439 B.n409 B.n166 10.6151
R2440 B.n410 B.n409 10.6151
R2441 B.n411 B.n410 10.6151
R2442 B.n411 B.n164 10.6151
R2443 B.n415 B.n164 10.6151
R2444 B.n416 B.n415 10.6151
R2445 B.n417 B.n416 10.6151
R2446 B.n417 B.n162 10.6151
R2447 B.n421 B.n162 10.6151
R2448 B.n422 B.n421 10.6151
R2449 B.n423 B.n422 10.6151
R2450 B.n423 B.n160 10.6151
R2451 B.n427 B.n160 10.6151
R2452 B.n428 B.n427 10.6151
R2453 B.n429 B.n428 10.6151
R2454 B.n429 B.n158 10.6151
R2455 B.n433 B.n158 10.6151
R2456 B.n434 B.n433 10.6151
R2457 B.n435 B.n434 10.6151
R2458 B.n435 B.n156 10.6151
R2459 B.n439 B.n156 10.6151
R2460 B.n440 B.n439 10.6151
R2461 B.n441 B.n440 10.6151
R2462 B.n441 B.n154 10.6151
R2463 B.n445 B.n154 10.6151
R2464 B.n446 B.n445 10.6151
R2465 B.n447 B.n446 10.6151
R2466 B.n447 B.n152 10.6151
R2467 B.n451 B.n152 10.6151
R2468 B.n452 B.n451 10.6151
R2469 B.n453 B.n452 10.6151
R2470 B.n453 B.n150 10.6151
R2471 B.n457 B.n150 10.6151
R2472 B.n458 B.n457 10.6151
R2473 B.n459 B.n458 10.6151
R2474 B.n459 B.n148 10.6151
R2475 B.n463 B.n148 10.6151
R2476 B.n733 B.n56 9.36635
R2477 B.n716 B.n715 9.36635
R2478 B.n382 B.n381 9.36635
R2479 B.n398 B.n168 9.36635
R2480 B.n889 B.n0 8.11757
R2481 B.n889 B.n1 8.11757
R2482 B.n730 B.n56 1.24928
R2483 B.n717 B.n716 1.24928
R2484 B.n383 B.n382 1.24928
R2485 B.n399 B.n398 1.24928
C0 w_n4678_n3398# VTAIL 3.25647f
C1 VP VN 8.66743f
C2 VDD2 VN 10.918401f
C3 VN VTAIL 11.6205f
C4 w_n4678_n3398# B 10.8582f
C5 w_n4678_n3398# VDD1 2.86146f
C6 B VN 1.32578f
C7 VDD2 VP 0.604065f
C8 VN VDD1 0.15379f
C9 VP VTAIL 11.6348f
C10 VDD2 VTAIL 10.5531f
C11 B VP 2.35165f
C12 VDD2 B 2.67905f
C13 VP VDD1 11.364799f
C14 B VTAIL 3.83049f
C15 VDD2 VDD1 2.27905f
C16 VTAIL VDD1 10.501f
C17 w_n4678_n3398# VN 10.0675f
C18 B VDD1 2.55491f
C19 w_n4678_n3398# VP 10.677099f
C20 VDD2 w_n4678_n3398# 3.01333f
C21 VDD2 VSUBS 2.241229f
C22 VDD1 VSUBS 2.030916f
C23 VTAIL VSUBS 1.340368f
C24 VN VSUBS 7.95825f
C25 VP VSUBS 4.459489f
C26 B VSUBS 5.57923f
C27 w_n4678_n3398# VSUBS 0.195634p
C28 B.n0 VSUBS 0.008166f
C29 B.n1 VSUBS 0.008166f
C30 B.n2 VSUBS 0.012077f
C31 B.n3 VSUBS 0.009254f
C32 B.n4 VSUBS 0.009254f
C33 B.n5 VSUBS 0.009254f
C34 B.n6 VSUBS 0.009254f
C35 B.n7 VSUBS 0.009254f
C36 B.n8 VSUBS 0.009254f
C37 B.n9 VSUBS 0.009254f
C38 B.n10 VSUBS 0.009254f
C39 B.n11 VSUBS 0.009254f
C40 B.n12 VSUBS 0.009254f
C41 B.n13 VSUBS 0.009254f
C42 B.n14 VSUBS 0.009254f
C43 B.n15 VSUBS 0.009254f
C44 B.n16 VSUBS 0.009254f
C45 B.n17 VSUBS 0.009254f
C46 B.n18 VSUBS 0.009254f
C47 B.n19 VSUBS 0.009254f
C48 B.n20 VSUBS 0.009254f
C49 B.n21 VSUBS 0.009254f
C50 B.n22 VSUBS 0.009254f
C51 B.n23 VSUBS 0.009254f
C52 B.n24 VSUBS 0.009254f
C53 B.n25 VSUBS 0.009254f
C54 B.n26 VSUBS 0.009254f
C55 B.n27 VSUBS 0.009254f
C56 B.n28 VSUBS 0.009254f
C57 B.n29 VSUBS 0.009254f
C58 B.n30 VSUBS 0.009254f
C59 B.n31 VSUBS 0.009254f
C60 B.n32 VSUBS 0.009254f
C61 B.n33 VSUBS 0.022298f
C62 B.n34 VSUBS 0.009254f
C63 B.n35 VSUBS 0.009254f
C64 B.n36 VSUBS 0.009254f
C65 B.n37 VSUBS 0.009254f
C66 B.n38 VSUBS 0.009254f
C67 B.n39 VSUBS 0.009254f
C68 B.n40 VSUBS 0.009254f
C69 B.n41 VSUBS 0.009254f
C70 B.n42 VSUBS 0.009254f
C71 B.n43 VSUBS 0.009254f
C72 B.n44 VSUBS 0.009254f
C73 B.n45 VSUBS 0.009254f
C74 B.n46 VSUBS 0.009254f
C75 B.n47 VSUBS 0.009254f
C76 B.n48 VSUBS 0.009254f
C77 B.n49 VSUBS 0.009254f
C78 B.n50 VSUBS 0.009254f
C79 B.n51 VSUBS 0.009254f
C80 B.n52 VSUBS 0.009254f
C81 B.n53 VSUBS 0.009254f
C82 B.t7 VSUBS 0.283566f
C83 B.t8 VSUBS 0.327751f
C84 B.t6 VSUBS 2.02588f
C85 B.n54 VSUBS 0.52046f
C86 B.n55 VSUBS 0.336408f
C87 B.n56 VSUBS 0.021441f
C88 B.n57 VSUBS 0.009254f
C89 B.n58 VSUBS 0.009254f
C90 B.n59 VSUBS 0.009254f
C91 B.n60 VSUBS 0.009254f
C92 B.n61 VSUBS 0.009254f
C93 B.t10 VSUBS 0.28357f
C94 B.t11 VSUBS 0.327754f
C95 B.t9 VSUBS 2.02588f
C96 B.n62 VSUBS 0.520457f
C97 B.n63 VSUBS 0.336404f
C98 B.n64 VSUBS 0.009254f
C99 B.n65 VSUBS 0.009254f
C100 B.n66 VSUBS 0.009254f
C101 B.n67 VSUBS 0.009254f
C102 B.n68 VSUBS 0.009254f
C103 B.n69 VSUBS 0.009254f
C104 B.n70 VSUBS 0.009254f
C105 B.n71 VSUBS 0.009254f
C106 B.n72 VSUBS 0.009254f
C107 B.n73 VSUBS 0.009254f
C108 B.n74 VSUBS 0.009254f
C109 B.n75 VSUBS 0.009254f
C110 B.n76 VSUBS 0.009254f
C111 B.n77 VSUBS 0.009254f
C112 B.n78 VSUBS 0.009254f
C113 B.n79 VSUBS 0.009254f
C114 B.n80 VSUBS 0.009254f
C115 B.n81 VSUBS 0.009254f
C116 B.n82 VSUBS 0.009254f
C117 B.n83 VSUBS 0.009254f
C118 B.n84 VSUBS 0.022298f
C119 B.n85 VSUBS 0.009254f
C120 B.n86 VSUBS 0.009254f
C121 B.n87 VSUBS 0.009254f
C122 B.n88 VSUBS 0.009254f
C123 B.n89 VSUBS 0.009254f
C124 B.n90 VSUBS 0.009254f
C125 B.n91 VSUBS 0.009254f
C126 B.n92 VSUBS 0.009254f
C127 B.n93 VSUBS 0.009254f
C128 B.n94 VSUBS 0.009254f
C129 B.n95 VSUBS 0.009254f
C130 B.n96 VSUBS 0.009254f
C131 B.n97 VSUBS 0.009254f
C132 B.n98 VSUBS 0.009254f
C133 B.n99 VSUBS 0.009254f
C134 B.n100 VSUBS 0.009254f
C135 B.n101 VSUBS 0.009254f
C136 B.n102 VSUBS 0.009254f
C137 B.n103 VSUBS 0.009254f
C138 B.n104 VSUBS 0.009254f
C139 B.n105 VSUBS 0.009254f
C140 B.n106 VSUBS 0.009254f
C141 B.n107 VSUBS 0.009254f
C142 B.n108 VSUBS 0.009254f
C143 B.n109 VSUBS 0.009254f
C144 B.n110 VSUBS 0.009254f
C145 B.n111 VSUBS 0.009254f
C146 B.n112 VSUBS 0.009254f
C147 B.n113 VSUBS 0.009254f
C148 B.n114 VSUBS 0.009254f
C149 B.n115 VSUBS 0.009254f
C150 B.n116 VSUBS 0.009254f
C151 B.n117 VSUBS 0.009254f
C152 B.n118 VSUBS 0.009254f
C153 B.n119 VSUBS 0.009254f
C154 B.n120 VSUBS 0.009254f
C155 B.n121 VSUBS 0.009254f
C156 B.n122 VSUBS 0.009254f
C157 B.n123 VSUBS 0.009254f
C158 B.n124 VSUBS 0.009254f
C159 B.n125 VSUBS 0.009254f
C160 B.n126 VSUBS 0.009254f
C161 B.n127 VSUBS 0.009254f
C162 B.n128 VSUBS 0.009254f
C163 B.n129 VSUBS 0.009254f
C164 B.n130 VSUBS 0.009254f
C165 B.n131 VSUBS 0.009254f
C166 B.n132 VSUBS 0.009254f
C167 B.n133 VSUBS 0.009254f
C168 B.n134 VSUBS 0.009254f
C169 B.n135 VSUBS 0.009254f
C170 B.n136 VSUBS 0.009254f
C171 B.n137 VSUBS 0.009254f
C172 B.n138 VSUBS 0.009254f
C173 B.n139 VSUBS 0.009254f
C174 B.n140 VSUBS 0.009254f
C175 B.n141 VSUBS 0.009254f
C176 B.n142 VSUBS 0.009254f
C177 B.n143 VSUBS 0.009254f
C178 B.n144 VSUBS 0.009254f
C179 B.n145 VSUBS 0.009254f
C180 B.n146 VSUBS 0.009254f
C181 B.n147 VSUBS 0.020708f
C182 B.n148 VSUBS 0.009254f
C183 B.n149 VSUBS 0.009254f
C184 B.n150 VSUBS 0.009254f
C185 B.n151 VSUBS 0.009254f
C186 B.n152 VSUBS 0.009254f
C187 B.n153 VSUBS 0.009254f
C188 B.n154 VSUBS 0.009254f
C189 B.n155 VSUBS 0.009254f
C190 B.n156 VSUBS 0.009254f
C191 B.n157 VSUBS 0.009254f
C192 B.n158 VSUBS 0.009254f
C193 B.n159 VSUBS 0.009254f
C194 B.n160 VSUBS 0.009254f
C195 B.n161 VSUBS 0.009254f
C196 B.n162 VSUBS 0.009254f
C197 B.n163 VSUBS 0.009254f
C198 B.n164 VSUBS 0.009254f
C199 B.n165 VSUBS 0.009254f
C200 B.n166 VSUBS 0.009254f
C201 B.n167 VSUBS 0.009254f
C202 B.n168 VSUBS 0.00871f
C203 B.n169 VSUBS 0.009254f
C204 B.n170 VSUBS 0.009254f
C205 B.n171 VSUBS 0.009254f
C206 B.n172 VSUBS 0.009254f
C207 B.n173 VSUBS 0.009254f
C208 B.t5 VSUBS 0.283566f
C209 B.t4 VSUBS 0.327751f
C210 B.t3 VSUBS 2.02588f
C211 B.n174 VSUBS 0.52046f
C212 B.n175 VSUBS 0.336408f
C213 B.n176 VSUBS 0.009254f
C214 B.n177 VSUBS 0.009254f
C215 B.n178 VSUBS 0.009254f
C216 B.n179 VSUBS 0.009254f
C217 B.n180 VSUBS 0.009254f
C218 B.n181 VSUBS 0.009254f
C219 B.n182 VSUBS 0.009254f
C220 B.n183 VSUBS 0.009254f
C221 B.n184 VSUBS 0.009254f
C222 B.n185 VSUBS 0.009254f
C223 B.n186 VSUBS 0.009254f
C224 B.n187 VSUBS 0.009254f
C225 B.n188 VSUBS 0.009254f
C226 B.n189 VSUBS 0.009254f
C227 B.n190 VSUBS 0.009254f
C228 B.n191 VSUBS 0.009254f
C229 B.n192 VSUBS 0.009254f
C230 B.n193 VSUBS 0.009254f
C231 B.n194 VSUBS 0.009254f
C232 B.n195 VSUBS 0.009254f
C233 B.n196 VSUBS 0.022298f
C234 B.n197 VSUBS 0.009254f
C235 B.n198 VSUBS 0.009254f
C236 B.n199 VSUBS 0.009254f
C237 B.n200 VSUBS 0.009254f
C238 B.n201 VSUBS 0.009254f
C239 B.n202 VSUBS 0.009254f
C240 B.n203 VSUBS 0.009254f
C241 B.n204 VSUBS 0.009254f
C242 B.n205 VSUBS 0.009254f
C243 B.n206 VSUBS 0.009254f
C244 B.n207 VSUBS 0.009254f
C245 B.n208 VSUBS 0.009254f
C246 B.n209 VSUBS 0.009254f
C247 B.n210 VSUBS 0.009254f
C248 B.n211 VSUBS 0.009254f
C249 B.n212 VSUBS 0.009254f
C250 B.n213 VSUBS 0.009254f
C251 B.n214 VSUBS 0.009254f
C252 B.n215 VSUBS 0.009254f
C253 B.n216 VSUBS 0.009254f
C254 B.n217 VSUBS 0.009254f
C255 B.n218 VSUBS 0.009254f
C256 B.n219 VSUBS 0.009254f
C257 B.n220 VSUBS 0.009254f
C258 B.n221 VSUBS 0.009254f
C259 B.n222 VSUBS 0.009254f
C260 B.n223 VSUBS 0.009254f
C261 B.n224 VSUBS 0.009254f
C262 B.n225 VSUBS 0.009254f
C263 B.n226 VSUBS 0.009254f
C264 B.n227 VSUBS 0.009254f
C265 B.n228 VSUBS 0.009254f
C266 B.n229 VSUBS 0.009254f
C267 B.n230 VSUBS 0.009254f
C268 B.n231 VSUBS 0.009254f
C269 B.n232 VSUBS 0.009254f
C270 B.n233 VSUBS 0.009254f
C271 B.n234 VSUBS 0.009254f
C272 B.n235 VSUBS 0.009254f
C273 B.n236 VSUBS 0.009254f
C274 B.n237 VSUBS 0.009254f
C275 B.n238 VSUBS 0.009254f
C276 B.n239 VSUBS 0.009254f
C277 B.n240 VSUBS 0.009254f
C278 B.n241 VSUBS 0.009254f
C279 B.n242 VSUBS 0.009254f
C280 B.n243 VSUBS 0.009254f
C281 B.n244 VSUBS 0.009254f
C282 B.n245 VSUBS 0.009254f
C283 B.n246 VSUBS 0.009254f
C284 B.n247 VSUBS 0.009254f
C285 B.n248 VSUBS 0.009254f
C286 B.n249 VSUBS 0.009254f
C287 B.n250 VSUBS 0.009254f
C288 B.n251 VSUBS 0.009254f
C289 B.n252 VSUBS 0.009254f
C290 B.n253 VSUBS 0.009254f
C291 B.n254 VSUBS 0.009254f
C292 B.n255 VSUBS 0.009254f
C293 B.n256 VSUBS 0.009254f
C294 B.n257 VSUBS 0.009254f
C295 B.n258 VSUBS 0.009254f
C296 B.n259 VSUBS 0.009254f
C297 B.n260 VSUBS 0.009254f
C298 B.n261 VSUBS 0.009254f
C299 B.n262 VSUBS 0.009254f
C300 B.n263 VSUBS 0.009254f
C301 B.n264 VSUBS 0.009254f
C302 B.n265 VSUBS 0.009254f
C303 B.n266 VSUBS 0.009254f
C304 B.n267 VSUBS 0.009254f
C305 B.n268 VSUBS 0.009254f
C306 B.n269 VSUBS 0.009254f
C307 B.n270 VSUBS 0.009254f
C308 B.n271 VSUBS 0.009254f
C309 B.n272 VSUBS 0.009254f
C310 B.n273 VSUBS 0.009254f
C311 B.n274 VSUBS 0.009254f
C312 B.n275 VSUBS 0.009254f
C313 B.n276 VSUBS 0.009254f
C314 B.n277 VSUBS 0.009254f
C315 B.n278 VSUBS 0.009254f
C316 B.n279 VSUBS 0.009254f
C317 B.n280 VSUBS 0.009254f
C318 B.n281 VSUBS 0.009254f
C319 B.n282 VSUBS 0.009254f
C320 B.n283 VSUBS 0.009254f
C321 B.n284 VSUBS 0.009254f
C322 B.n285 VSUBS 0.009254f
C323 B.n286 VSUBS 0.009254f
C324 B.n287 VSUBS 0.009254f
C325 B.n288 VSUBS 0.009254f
C326 B.n289 VSUBS 0.009254f
C327 B.n290 VSUBS 0.009254f
C328 B.n291 VSUBS 0.009254f
C329 B.n292 VSUBS 0.009254f
C330 B.n293 VSUBS 0.009254f
C331 B.n294 VSUBS 0.009254f
C332 B.n295 VSUBS 0.009254f
C333 B.n296 VSUBS 0.009254f
C334 B.n297 VSUBS 0.009254f
C335 B.n298 VSUBS 0.009254f
C336 B.n299 VSUBS 0.009254f
C337 B.n300 VSUBS 0.009254f
C338 B.n301 VSUBS 0.009254f
C339 B.n302 VSUBS 0.009254f
C340 B.n303 VSUBS 0.009254f
C341 B.n304 VSUBS 0.009254f
C342 B.n305 VSUBS 0.009254f
C343 B.n306 VSUBS 0.009254f
C344 B.n307 VSUBS 0.009254f
C345 B.n308 VSUBS 0.009254f
C346 B.n309 VSUBS 0.009254f
C347 B.n310 VSUBS 0.009254f
C348 B.n311 VSUBS 0.009254f
C349 B.n312 VSUBS 0.009254f
C350 B.n313 VSUBS 0.009254f
C351 B.n314 VSUBS 0.009254f
C352 B.n315 VSUBS 0.009254f
C353 B.n316 VSUBS 0.009254f
C354 B.n317 VSUBS 0.020708f
C355 B.n318 VSUBS 0.020708f
C356 B.n319 VSUBS 0.022298f
C357 B.n320 VSUBS 0.009254f
C358 B.n321 VSUBS 0.009254f
C359 B.n322 VSUBS 0.009254f
C360 B.n323 VSUBS 0.009254f
C361 B.n324 VSUBS 0.009254f
C362 B.n325 VSUBS 0.009254f
C363 B.n326 VSUBS 0.009254f
C364 B.n327 VSUBS 0.009254f
C365 B.n328 VSUBS 0.009254f
C366 B.n329 VSUBS 0.009254f
C367 B.n330 VSUBS 0.009254f
C368 B.n331 VSUBS 0.009254f
C369 B.n332 VSUBS 0.009254f
C370 B.n333 VSUBS 0.009254f
C371 B.n334 VSUBS 0.009254f
C372 B.n335 VSUBS 0.009254f
C373 B.n336 VSUBS 0.009254f
C374 B.n337 VSUBS 0.009254f
C375 B.n338 VSUBS 0.009254f
C376 B.n339 VSUBS 0.009254f
C377 B.n340 VSUBS 0.009254f
C378 B.n341 VSUBS 0.009254f
C379 B.n342 VSUBS 0.009254f
C380 B.n343 VSUBS 0.009254f
C381 B.n344 VSUBS 0.009254f
C382 B.n345 VSUBS 0.009254f
C383 B.n346 VSUBS 0.009254f
C384 B.n347 VSUBS 0.009254f
C385 B.n348 VSUBS 0.009254f
C386 B.n349 VSUBS 0.009254f
C387 B.n350 VSUBS 0.009254f
C388 B.n351 VSUBS 0.009254f
C389 B.n352 VSUBS 0.009254f
C390 B.n353 VSUBS 0.009254f
C391 B.n354 VSUBS 0.009254f
C392 B.n355 VSUBS 0.009254f
C393 B.n356 VSUBS 0.009254f
C394 B.n357 VSUBS 0.009254f
C395 B.n358 VSUBS 0.009254f
C396 B.n359 VSUBS 0.009254f
C397 B.n360 VSUBS 0.009254f
C398 B.n361 VSUBS 0.009254f
C399 B.n362 VSUBS 0.009254f
C400 B.n363 VSUBS 0.009254f
C401 B.n364 VSUBS 0.009254f
C402 B.n365 VSUBS 0.009254f
C403 B.n366 VSUBS 0.009254f
C404 B.n367 VSUBS 0.009254f
C405 B.n368 VSUBS 0.009254f
C406 B.n369 VSUBS 0.009254f
C407 B.n370 VSUBS 0.009254f
C408 B.n371 VSUBS 0.009254f
C409 B.n372 VSUBS 0.009254f
C410 B.n373 VSUBS 0.009254f
C411 B.n374 VSUBS 0.009254f
C412 B.n375 VSUBS 0.009254f
C413 B.n376 VSUBS 0.009254f
C414 B.n377 VSUBS 0.009254f
C415 B.n378 VSUBS 0.009254f
C416 B.n379 VSUBS 0.009254f
C417 B.n380 VSUBS 0.009254f
C418 B.n381 VSUBS 0.00871f
C419 B.n382 VSUBS 0.021441f
C420 B.n383 VSUBS 0.005172f
C421 B.n384 VSUBS 0.009254f
C422 B.n385 VSUBS 0.009254f
C423 B.n386 VSUBS 0.009254f
C424 B.n387 VSUBS 0.009254f
C425 B.n388 VSUBS 0.009254f
C426 B.n389 VSUBS 0.009254f
C427 B.n390 VSUBS 0.009254f
C428 B.n391 VSUBS 0.009254f
C429 B.n392 VSUBS 0.009254f
C430 B.n393 VSUBS 0.009254f
C431 B.n394 VSUBS 0.009254f
C432 B.n395 VSUBS 0.009254f
C433 B.t2 VSUBS 0.28357f
C434 B.t1 VSUBS 0.327754f
C435 B.t0 VSUBS 2.02588f
C436 B.n396 VSUBS 0.520457f
C437 B.n397 VSUBS 0.336404f
C438 B.n398 VSUBS 0.021441f
C439 B.n399 VSUBS 0.005172f
C440 B.n400 VSUBS 0.009254f
C441 B.n401 VSUBS 0.009254f
C442 B.n402 VSUBS 0.009254f
C443 B.n403 VSUBS 0.009254f
C444 B.n404 VSUBS 0.009254f
C445 B.n405 VSUBS 0.009254f
C446 B.n406 VSUBS 0.009254f
C447 B.n407 VSUBS 0.009254f
C448 B.n408 VSUBS 0.009254f
C449 B.n409 VSUBS 0.009254f
C450 B.n410 VSUBS 0.009254f
C451 B.n411 VSUBS 0.009254f
C452 B.n412 VSUBS 0.009254f
C453 B.n413 VSUBS 0.009254f
C454 B.n414 VSUBS 0.009254f
C455 B.n415 VSUBS 0.009254f
C456 B.n416 VSUBS 0.009254f
C457 B.n417 VSUBS 0.009254f
C458 B.n418 VSUBS 0.009254f
C459 B.n419 VSUBS 0.009254f
C460 B.n420 VSUBS 0.009254f
C461 B.n421 VSUBS 0.009254f
C462 B.n422 VSUBS 0.009254f
C463 B.n423 VSUBS 0.009254f
C464 B.n424 VSUBS 0.009254f
C465 B.n425 VSUBS 0.009254f
C466 B.n426 VSUBS 0.009254f
C467 B.n427 VSUBS 0.009254f
C468 B.n428 VSUBS 0.009254f
C469 B.n429 VSUBS 0.009254f
C470 B.n430 VSUBS 0.009254f
C471 B.n431 VSUBS 0.009254f
C472 B.n432 VSUBS 0.009254f
C473 B.n433 VSUBS 0.009254f
C474 B.n434 VSUBS 0.009254f
C475 B.n435 VSUBS 0.009254f
C476 B.n436 VSUBS 0.009254f
C477 B.n437 VSUBS 0.009254f
C478 B.n438 VSUBS 0.009254f
C479 B.n439 VSUBS 0.009254f
C480 B.n440 VSUBS 0.009254f
C481 B.n441 VSUBS 0.009254f
C482 B.n442 VSUBS 0.009254f
C483 B.n443 VSUBS 0.009254f
C484 B.n444 VSUBS 0.009254f
C485 B.n445 VSUBS 0.009254f
C486 B.n446 VSUBS 0.009254f
C487 B.n447 VSUBS 0.009254f
C488 B.n448 VSUBS 0.009254f
C489 B.n449 VSUBS 0.009254f
C490 B.n450 VSUBS 0.009254f
C491 B.n451 VSUBS 0.009254f
C492 B.n452 VSUBS 0.009254f
C493 B.n453 VSUBS 0.009254f
C494 B.n454 VSUBS 0.009254f
C495 B.n455 VSUBS 0.009254f
C496 B.n456 VSUBS 0.009254f
C497 B.n457 VSUBS 0.009254f
C498 B.n458 VSUBS 0.009254f
C499 B.n459 VSUBS 0.009254f
C500 B.n460 VSUBS 0.009254f
C501 B.n461 VSUBS 0.009254f
C502 B.n462 VSUBS 0.022298f
C503 B.n463 VSUBS 0.021193f
C504 B.n464 VSUBS 0.021813f
C505 B.n465 VSUBS 0.009254f
C506 B.n466 VSUBS 0.009254f
C507 B.n467 VSUBS 0.009254f
C508 B.n468 VSUBS 0.009254f
C509 B.n469 VSUBS 0.009254f
C510 B.n470 VSUBS 0.009254f
C511 B.n471 VSUBS 0.009254f
C512 B.n472 VSUBS 0.009254f
C513 B.n473 VSUBS 0.009254f
C514 B.n474 VSUBS 0.009254f
C515 B.n475 VSUBS 0.009254f
C516 B.n476 VSUBS 0.009254f
C517 B.n477 VSUBS 0.009254f
C518 B.n478 VSUBS 0.009254f
C519 B.n479 VSUBS 0.009254f
C520 B.n480 VSUBS 0.009254f
C521 B.n481 VSUBS 0.009254f
C522 B.n482 VSUBS 0.009254f
C523 B.n483 VSUBS 0.009254f
C524 B.n484 VSUBS 0.009254f
C525 B.n485 VSUBS 0.009254f
C526 B.n486 VSUBS 0.009254f
C527 B.n487 VSUBS 0.009254f
C528 B.n488 VSUBS 0.009254f
C529 B.n489 VSUBS 0.009254f
C530 B.n490 VSUBS 0.009254f
C531 B.n491 VSUBS 0.009254f
C532 B.n492 VSUBS 0.009254f
C533 B.n493 VSUBS 0.009254f
C534 B.n494 VSUBS 0.009254f
C535 B.n495 VSUBS 0.009254f
C536 B.n496 VSUBS 0.009254f
C537 B.n497 VSUBS 0.009254f
C538 B.n498 VSUBS 0.009254f
C539 B.n499 VSUBS 0.009254f
C540 B.n500 VSUBS 0.009254f
C541 B.n501 VSUBS 0.009254f
C542 B.n502 VSUBS 0.009254f
C543 B.n503 VSUBS 0.009254f
C544 B.n504 VSUBS 0.009254f
C545 B.n505 VSUBS 0.009254f
C546 B.n506 VSUBS 0.009254f
C547 B.n507 VSUBS 0.009254f
C548 B.n508 VSUBS 0.009254f
C549 B.n509 VSUBS 0.009254f
C550 B.n510 VSUBS 0.009254f
C551 B.n511 VSUBS 0.009254f
C552 B.n512 VSUBS 0.009254f
C553 B.n513 VSUBS 0.009254f
C554 B.n514 VSUBS 0.009254f
C555 B.n515 VSUBS 0.009254f
C556 B.n516 VSUBS 0.009254f
C557 B.n517 VSUBS 0.009254f
C558 B.n518 VSUBS 0.009254f
C559 B.n519 VSUBS 0.009254f
C560 B.n520 VSUBS 0.009254f
C561 B.n521 VSUBS 0.009254f
C562 B.n522 VSUBS 0.009254f
C563 B.n523 VSUBS 0.009254f
C564 B.n524 VSUBS 0.009254f
C565 B.n525 VSUBS 0.009254f
C566 B.n526 VSUBS 0.009254f
C567 B.n527 VSUBS 0.009254f
C568 B.n528 VSUBS 0.009254f
C569 B.n529 VSUBS 0.009254f
C570 B.n530 VSUBS 0.009254f
C571 B.n531 VSUBS 0.009254f
C572 B.n532 VSUBS 0.009254f
C573 B.n533 VSUBS 0.009254f
C574 B.n534 VSUBS 0.009254f
C575 B.n535 VSUBS 0.009254f
C576 B.n536 VSUBS 0.009254f
C577 B.n537 VSUBS 0.009254f
C578 B.n538 VSUBS 0.009254f
C579 B.n539 VSUBS 0.009254f
C580 B.n540 VSUBS 0.009254f
C581 B.n541 VSUBS 0.009254f
C582 B.n542 VSUBS 0.009254f
C583 B.n543 VSUBS 0.009254f
C584 B.n544 VSUBS 0.009254f
C585 B.n545 VSUBS 0.009254f
C586 B.n546 VSUBS 0.009254f
C587 B.n547 VSUBS 0.009254f
C588 B.n548 VSUBS 0.009254f
C589 B.n549 VSUBS 0.009254f
C590 B.n550 VSUBS 0.009254f
C591 B.n551 VSUBS 0.009254f
C592 B.n552 VSUBS 0.009254f
C593 B.n553 VSUBS 0.009254f
C594 B.n554 VSUBS 0.009254f
C595 B.n555 VSUBS 0.009254f
C596 B.n556 VSUBS 0.009254f
C597 B.n557 VSUBS 0.009254f
C598 B.n558 VSUBS 0.009254f
C599 B.n559 VSUBS 0.009254f
C600 B.n560 VSUBS 0.009254f
C601 B.n561 VSUBS 0.009254f
C602 B.n562 VSUBS 0.009254f
C603 B.n563 VSUBS 0.009254f
C604 B.n564 VSUBS 0.009254f
C605 B.n565 VSUBS 0.009254f
C606 B.n566 VSUBS 0.009254f
C607 B.n567 VSUBS 0.009254f
C608 B.n568 VSUBS 0.009254f
C609 B.n569 VSUBS 0.009254f
C610 B.n570 VSUBS 0.009254f
C611 B.n571 VSUBS 0.009254f
C612 B.n572 VSUBS 0.009254f
C613 B.n573 VSUBS 0.009254f
C614 B.n574 VSUBS 0.009254f
C615 B.n575 VSUBS 0.009254f
C616 B.n576 VSUBS 0.009254f
C617 B.n577 VSUBS 0.009254f
C618 B.n578 VSUBS 0.009254f
C619 B.n579 VSUBS 0.009254f
C620 B.n580 VSUBS 0.009254f
C621 B.n581 VSUBS 0.009254f
C622 B.n582 VSUBS 0.009254f
C623 B.n583 VSUBS 0.009254f
C624 B.n584 VSUBS 0.009254f
C625 B.n585 VSUBS 0.009254f
C626 B.n586 VSUBS 0.009254f
C627 B.n587 VSUBS 0.009254f
C628 B.n588 VSUBS 0.009254f
C629 B.n589 VSUBS 0.009254f
C630 B.n590 VSUBS 0.009254f
C631 B.n591 VSUBS 0.009254f
C632 B.n592 VSUBS 0.009254f
C633 B.n593 VSUBS 0.009254f
C634 B.n594 VSUBS 0.009254f
C635 B.n595 VSUBS 0.009254f
C636 B.n596 VSUBS 0.009254f
C637 B.n597 VSUBS 0.009254f
C638 B.n598 VSUBS 0.009254f
C639 B.n599 VSUBS 0.009254f
C640 B.n600 VSUBS 0.009254f
C641 B.n601 VSUBS 0.009254f
C642 B.n602 VSUBS 0.009254f
C643 B.n603 VSUBS 0.009254f
C644 B.n604 VSUBS 0.009254f
C645 B.n605 VSUBS 0.009254f
C646 B.n606 VSUBS 0.009254f
C647 B.n607 VSUBS 0.009254f
C648 B.n608 VSUBS 0.009254f
C649 B.n609 VSUBS 0.009254f
C650 B.n610 VSUBS 0.009254f
C651 B.n611 VSUBS 0.009254f
C652 B.n612 VSUBS 0.009254f
C653 B.n613 VSUBS 0.009254f
C654 B.n614 VSUBS 0.009254f
C655 B.n615 VSUBS 0.009254f
C656 B.n616 VSUBS 0.009254f
C657 B.n617 VSUBS 0.009254f
C658 B.n618 VSUBS 0.009254f
C659 B.n619 VSUBS 0.009254f
C660 B.n620 VSUBS 0.009254f
C661 B.n621 VSUBS 0.009254f
C662 B.n622 VSUBS 0.009254f
C663 B.n623 VSUBS 0.009254f
C664 B.n624 VSUBS 0.009254f
C665 B.n625 VSUBS 0.009254f
C666 B.n626 VSUBS 0.009254f
C667 B.n627 VSUBS 0.009254f
C668 B.n628 VSUBS 0.009254f
C669 B.n629 VSUBS 0.009254f
C670 B.n630 VSUBS 0.009254f
C671 B.n631 VSUBS 0.009254f
C672 B.n632 VSUBS 0.009254f
C673 B.n633 VSUBS 0.009254f
C674 B.n634 VSUBS 0.009254f
C675 B.n635 VSUBS 0.009254f
C676 B.n636 VSUBS 0.009254f
C677 B.n637 VSUBS 0.009254f
C678 B.n638 VSUBS 0.009254f
C679 B.n639 VSUBS 0.009254f
C680 B.n640 VSUBS 0.009254f
C681 B.n641 VSUBS 0.009254f
C682 B.n642 VSUBS 0.009254f
C683 B.n643 VSUBS 0.009254f
C684 B.n644 VSUBS 0.009254f
C685 B.n645 VSUBS 0.009254f
C686 B.n646 VSUBS 0.009254f
C687 B.n647 VSUBS 0.009254f
C688 B.n648 VSUBS 0.009254f
C689 B.n649 VSUBS 0.009254f
C690 B.n650 VSUBS 0.009254f
C691 B.n651 VSUBS 0.020708f
C692 B.n652 VSUBS 0.020708f
C693 B.n653 VSUBS 0.022298f
C694 B.n654 VSUBS 0.009254f
C695 B.n655 VSUBS 0.009254f
C696 B.n656 VSUBS 0.009254f
C697 B.n657 VSUBS 0.009254f
C698 B.n658 VSUBS 0.009254f
C699 B.n659 VSUBS 0.009254f
C700 B.n660 VSUBS 0.009254f
C701 B.n661 VSUBS 0.009254f
C702 B.n662 VSUBS 0.009254f
C703 B.n663 VSUBS 0.009254f
C704 B.n664 VSUBS 0.009254f
C705 B.n665 VSUBS 0.009254f
C706 B.n666 VSUBS 0.009254f
C707 B.n667 VSUBS 0.009254f
C708 B.n668 VSUBS 0.009254f
C709 B.n669 VSUBS 0.009254f
C710 B.n670 VSUBS 0.009254f
C711 B.n671 VSUBS 0.009254f
C712 B.n672 VSUBS 0.009254f
C713 B.n673 VSUBS 0.009254f
C714 B.n674 VSUBS 0.009254f
C715 B.n675 VSUBS 0.009254f
C716 B.n676 VSUBS 0.009254f
C717 B.n677 VSUBS 0.009254f
C718 B.n678 VSUBS 0.009254f
C719 B.n679 VSUBS 0.009254f
C720 B.n680 VSUBS 0.009254f
C721 B.n681 VSUBS 0.009254f
C722 B.n682 VSUBS 0.009254f
C723 B.n683 VSUBS 0.009254f
C724 B.n684 VSUBS 0.009254f
C725 B.n685 VSUBS 0.009254f
C726 B.n686 VSUBS 0.009254f
C727 B.n687 VSUBS 0.009254f
C728 B.n688 VSUBS 0.009254f
C729 B.n689 VSUBS 0.009254f
C730 B.n690 VSUBS 0.009254f
C731 B.n691 VSUBS 0.009254f
C732 B.n692 VSUBS 0.009254f
C733 B.n693 VSUBS 0.009254f
C734 B.n694 VSUBS 0.009254f
C735 B.n695 VSUBS 0.009254f
C736 B.n696 VSUBS 0.009254f
C737 B.n697 VSUBS 0.009254f
C738 B.n698 VSUBS 0.009254f
C739 B.n699 VSUBS 0.009254f
C740 B.n700 VSUBS 0.009254f
C741 B.n701 VSUBS 0.009254f
C742 B.n702 VSUBS 0.009254f
C743 B.n703 VSUBS 0.009254f
C744 B.n704 VSUBS 0.009254f
C745 B.n705 VSUBS 0.009254f
C746 B.n706 VSUBS 0.009254f
C747 B.n707 VSUBS 0.009254f
C748 B.n708 VSUBS 0.009254f
C749 B.n709 VSUBS 0.009254f
C750 B.n710 VSUBS 0.009254f
C751 B.n711 VSUBS 0.009254f
C752 B.n712 VSUBS 0.009254f
C753 B.n713 VSUBS 0.009254f
C754 B.n714 VSUBS 0.009254f
C755 B.n715 VSUBS 0.00871f
C756 B.n716 VSUBS 0.021441f
C757 B.n717 VSUBS 0.005172f
C758 B.n718 VSUBS 0.009254f
C759 B.n719 VSUBS 0.009254f
C760 B.n720 VSUBS 0.009254f
C761 B.n721 VSUBS 0.009254f
C762 B.n722 VSUBS 0.009254f
C763 B.n723 VSUBS 0.009254f
C764 B.n724 VSUBS 0.009254f
C765 B.n725 VSUBS 0.009254f
C766 B.n726 VSUBS 0.009254f
C767 B.n727 VSUBS 0.009254f
C768 B.n728 VSUBS 0.009254f
C769 B.n729 VSUBS 0.009254f
C770 B.n730 VSUBS 0.005172f
C771 B.n731 VSUBS 0.009254f
C772 B.n732 VSUBS 0.009254f
C773 B.n733 VSUBS 0.00871f
C774 B.n734 VSUBS 0.009254f
C775 B.n735 VSUBS 0.009254f
C776 B.n736 VSUBS 0.009254f
C777 B.n737 VSUBS 0.009254f
C778 B.n738 VSUBS 0.009254f
C779 B.n739 VSUBS 0.009254f
C780 B.n740 VSUBS 0.009254f
C781 B.n741 VSUBS 0.009254f
C782 B.n742 VSUBS 0.009254f
C783 B.n743 VSUBS 0.009254f
C784 B.n744 VSUBS 0.009254f
C785 B.n745 VSUBS 0.009254f
C786 B.n746 VSUBS 0.009254f
C787 B.n747 VSUBS 0.009254f
C788 B.n748 VSUBS 0.009254f
C789 B.n749 VSUBS 0.009254f
C790 B.n750 VSUBS 0.009254f
C791 B.n751 VSUBS 0.009254f
C792 B.n752 VSUBS 0.009254f
C793 B.n753 VSUBS 0.009254f
C794 B.n754 VSUBS 0.009254f
C795 B.n755 VSUBS 0.009254f
C796 B.n756 VSUBS 0.009254f
C797 B.n757 VSUBS 0.009254f
C798 B.n758 VSUBS 0.009254f
C799 B.n759 VSUBS 0.009254f
C800 B.n760 VSUBS 0.009254f
C801 B.n761 VSUBS 0.009254f
C802 B.n762 VSUBS 0.009254f
C803 B.n763 VSUBS 0.009254f
C804 B.n764 VSUBS 0.009254f
C805 B.n765 VSUBS 0.009254f
C806 B.n766 VSUBS 0.009254f
C807 B.n767 VSUBS 0.009254f
C808 B.n768 VSUBS 0.009254f
C809 B.n769 VSUBS 0.009254f
C810 B.n770 VSUBS 0.009254f
C811 B.n771 VSUBS 0.009254f
C812 B.n772 VSUBS 0.009254f
C813 B.n773 VSUBS 0.009254f
C814 B.n774 VSUBS 0.009254f
C815 B.n775 VSUBS 0.009254f
C816 B.n776 VSUBS 0.009254f
C817 B.n777 VSUBS 0.009254f
C818 B.n778 VSUBS 0.009254f
C819 B.n779 VSUBS 0.009254f
C820 B.n780 VSUBS 0.009254f
C821 B.n781 VSUBS 0.009254f
C822 B.n782 VSUBS 0.009254f
C823 B.n783 VSUBS 0.009254f
C824 B.n784 VSUBS 0.009254f
C825 B.n785 VSUBS 0.009254f
C826 B.n786 VSUBS 0.009254f
C827 B.n787 VSUBS 0.009254f
C828 B.n788 VSUBS 0.009254f
C829 B.n789 VSUBS 0.009254f
C830 B.n790 VSUBS 0.009254f
C831 B.n791 VSUBS 0.009254f
C832 B.n792 VSUBS 0.009254f
C833 B.n793 VSUBS 0.009254f
C834 B.n794 VSUBS 0.022298f
C835 B.n795 VSUBS 0.020708f
C836 B.n796 VSUBS 0.020708f
C837 B.n797 VSUBS 0.009254f
C838 B.n798 VSUBS 0.009254f
C839 B.n799 VSUBS 0.009254f
C840 B.n800 VSUBS 0.009254f
C841 B.n801 VSUBS 0.009254f
C842 B.n802 VSUBS 0.009254f
C843 B.n803 VSUBS 0.009254f
C844 B.n804 VSUBS 0.009254f
C845 B.n805 VSUBS 0.009254f
C846 B.n806 VSUBS 0.009254f
C847 B.n807 VSUBS 0.009254f
C848 B.n808 VSUBS 0.009254f
C849 B.n809 VSUBS 0.009254f
C850 B.n810 VSUBS 0.009254f
C851 B.n811 VSUBS 0.009254f
C852 B.n812 VSUBS 0.009254f
C853 B.n813 VSUBS 0.009254f
C854 B.n814 VSUBS 0.009254f
C855 B.n815 VSUBS 0.009254f
C856 B.n816 VSUBS 0.009254f
C857 B.n817 VSUBS 0.009254f
C858 B.n818 VSUBS 0.009254f
C859 B.n819 VSUBS 0.009254f
C860 B.n820 VSUBS 0.009254f
C861 B.n821 VSUBS 0.009254f
C862 B.n822 VSUBS 0.009254f
C863 B.n823 VSUBS 0.009254f
C864 B.n824 VSUBS 0.009254f
C865 B.n825 VSUBS 0.009254f
C866 B.n826 VSUBS 0.009254f
C867 B.n827 VSUBS 0.009254f
C868 B.n828 VSUBS 0.009254f
C869 B.n829 VSUBS 0.009254f
C870 B.n830 VSUBS 0.009254f
C871 B.n831 VSUBS 0.009254f
C872 B.n832 VSUBS 0.009254f
C873 B.n833 VSUBS 0.009254f
C874 B.n834 VSUBS 0.009254f
C875 B.n835 VSUBS 0.009254f
C876 B.n836 VSUBS 0.009254f
C877 B.n837 VSUBS 0.009254f
C878 B.n838 VSUBS 0.009254f
C879 B.n839 VSUBS 0.009254f
C880 B.n840 VSUBS 0.009254f
C881 B.n841 VSUBS 0.009254f
C882 B.n842 VSUBS 0.009254f
C883 B.n843 VSUBS 0.009254f
C884 B.n844 VSUBS 0.009254f
C885 B.n845 VSUBS 0.009254f
C886 B.n846 VSUBS 0.009254f
C887 B.n847 VSUBS 0.009254f
C888 B.n848 VSUBS 0.009254f
C889 B.n849 VSUBS 0.009254f
C890 B.n850 VSUBS 0.009254f
C891 B.n851 VSUBS 0.009254f
C892 B.n852 VSUBS 0.009254f
C893 B.n853 VSUBS 0.009254f
C894 B.n854 VSUBS 0.009254f
C895 B.n855 VSUBS 0.009254f
C896 B.n856 VSUBS 0.009254f
C897 B.n857 VSUBS 0.009254f
C898 B.n858 VSUBS 0.009254f
C899 B.n859 VSUBS 0.009254f
C900 B.n860 VSUBS 0.009254f
C901 B.n861 VSUBS 0.009254f
C902 B.n862 VSUBS 0.009254f
C903 B.n863 VSUBS 0.009254f
C904 B.n864 VSUBS 0.009254f
C905 B.n865 VSUBS 0.009254f
C906 B.n866 VSUBS 0.009254f
C907 B.n867 VSUBS 0.009254f
C908 B.n868 VSUBS 0.009254f
C909 B.n869 VSUBS 0.009254f
C910 B.n870 VSUBS 0.009254f
C911 B.n871 VSUBS 0.009254f
C912 B.n872 VSUBS 0.009254f
C913 B.n873 VSUBS 0.009254f
C914 B.n874 VSUBS 0.009254f
C915 B.n875 VSUBS 0.009254f
C916 B.n876 VSUBS 0.009254f
C917 B.n877 VSUBS 0.009254f
C918 B.n878 VSUBS 0.009254f
C919 B.n879 VSUBS 0.009254f
C920 B.n880 VSUBS 0.009254f
C921 B.n881 VSUBS 0.009254f
C922 B.n882 VSUBS 0.009254f
C923 B.n883 VSUBS 0.009254f
C924 B.n884 VSUBS 0.009254f
C925 B.n885 VSUBS 0.009254f
C926 B.n886 VSUBS 0.009254f
C927 B.n887 VSUBS 0.012077f
C928 B.n888 VSUBS 0.012865f
C929 B.n889 VSUBS 0.025583f
C930 VDD2.n0 VSUBS 0.033457f
C931 VDD2.n1 VSUBS 0.030215f
C932 VDD2.n2 VSUBS 0.016236f
C933 VDD2.n3 VSUBS 0.038376f
C934 VDD2.n4 VSUBS 0.017191f
C935 VDD2.n5 VSUBS 0.030215f
C936 VDD2.n6 VSUBS 0.016236f
C937 VDD2.n7 VSUBS 0.038376f
C938 VDD2.n8 VSUBS 0.017191f
C939 VDD2.n9 VSUBS 0.030215f
C940 VDD2.n10 VSUBS 0.016713f
C941 VDD2.n11 VSUBS 0.038376f
C942 VDD2.n12 VSUBS 0.017191f
C943 VDD2.n13 VSUBS 0.030215f
C944 VDD2.n14 VSUBS 0.016236f
C945 VDD2.n15 VSUBS 0.038376f
C946 VDD2.n16 VSUBS 0.017191f
C947 VDD2.n17 VSUBS 0.030215f
C948 VDD2.n18 VSUBS 0.016236f
C949 VDD2.n19 VSUBS 0.028782f
C950 VDD2.n20 VSUBS 0.028869f
C951 VDD2.t4 VSUBS 0.082712f
C952 VDD2.n21 VSUBS 0.240008f
C953 VDD2.n22 VSUBS 1.5044f
C954 VDD2.n23 VSUBS 0.016236f
C955 VDD2.n24 VSUBS 0.017191f
C956 VDD2.n25 VSUBS 0.038376f
C957 VDD2.n26 VSUBS 0.038376f
C958 VDD2.n27 VSUBS 0.017191f
C959 VDD2.n28 VSUBS 0.016236f
C960 VDD2.n29 VSUBS 0.030215f
C961 VDD2.n30 VSUBS 0.030215f
C962 VDD2.n31 VSUBS 0.016236f
C963 VDD2.n32 VSUBS 0.017191f
C964 VDD2.n33 VSUBS 0.038376f
C965 VDD2.n34 VSUBS 0.038376f
C966 VDD2.n35 VSUBS 0.017191f
C967 VDD2.n36 VSUBS 0.016236f
C968 VDD2.n37 VSUBS 0.030215f
C969 VDD2.n38 VSUBS 0.030215f
C970 VDD2.n39 VSUBS 0.016236f
C971 VDD2.n40 VSUBS 0.016236f
C972 VDD2.n41 VSUBS 0.017191f
C973 VDD2.n42 VSUBS 0.038376f
C974 VDD2.n43 VSUBS 0.038376f
C975 VDD2.n44 VSUBS 0.038376f
C976 VDD2.n45 VSUBS 0.016713f
C977 VDD2.n46 VSUBS 0.016236f
C978 VDD2.n47 VSUBS 0.030215f
C979 VDD2.n48 VSUBS 0.030215f
C980 VDD2.n49 VSUBS 0.016236f
C981 VDD2.n50 VSUBS 0.017191f
C982 VDD2.n51 VSUBS 0.038376f
C983 VDD2.n52 VSUBS 0.038376f
C984 VDD2.n53 VSUBS 0.017191f
C985 VDD2.n54 VSUBS 0.016236f
C986 VDD2.n55 VSUBS 0.030215f
C987 VDD2.n56 VSUBS 0.030215f
C988 VDD2.n57 VSUBS 0.016236f
C989 VDD2.n58 VSUBS 0.017191f
C990 VDD2.n59 VSUBS 0.038376f
C991 VDD2.n60 VSUBS 0.093783f
C992 VDD2.n61 VSUBS 0.017191f
C993 VDD2.n62 VSUBS 0.016236f
C994 VDD2.n63 VSUBS 0.071078f
C995 VDD2.n64 VSUBS 0.08436f
C996 VDD2.t5 VSUBS 0.290099f
C997 VDD2.t7 VSUBS 0.290099f
C998 VDD2.n65 VSUBS 2.27043f
C999 VDD2.n66 VSUBS 1.18869f
C1000 VDD2.t2 VSUBS 0.290099f
C1001 VDD2.t9 VSUBS 0.290099f
C1002 VDD2.n67 VSUBS 2.29657f
C1003 VDD2.n68 VSUBS 3.93688f
C1004 VDD2.n69 VSUBS 0.033457f
C1005 VDD2.n70 VSUBS 0.030215f
C1006 VDD2.n71 VSUBS 0.016236f
C1007 VDD2.n72 VSUBS 0.038376f
C1008 VDD2.n73 VSUBS 0.017191f
C1009 VDD2.n74 VSUBS 0.030215f
C1010 VDD2.n75 VSUBS 0.016236f
C1011 VDD2.n76 VSUBS 0.038376f
C1012 VDD2.n77 VSUBS 0.017191f
C1013 VDD2.n78 VSUBS 0.030215f
C1014 VDD2.n79 VSUBS 0.016713f
C1015 VDD2.n80 VSUBS 0.038376f
C1016 VDD2.n81 VSUBS 0.016236f
C1017 VDD2.n82 VSUBS 0.017191f
C1018 VDD2.n83 VSUBS 0.030215f
C1019 VDD2.n84 VSUBS 0.016236f
C1020 VDD2.n85 VSUBS 0.038376f
C1021 VDD2.n86 VSUBS 0.017191f
C1022 VDD2.n87 VSUBS 0.030215f
C1023 VDD2.n88 VSUBS 0.016236f
C1024 VDD2.n89 VSUBS 0.028782f
C1025 VDD2.n90 VSUBS 0.028869f
C1026 VDD2.t0 VSUBS 0.082712f
C1027 VDD2.n91 VSUBS 0.240008f
C1028 VDD2.n92 VSUBS 1.5044f
C1029 VDD2.n93 VSUBS 0.016236f
C1030 VDD2.n94 VSUBS 0.017191f
C1031 VDD2.n95 VSUBS 0.038376f
C1032 VDD2.n96 VSUBS 0.038376f
C1033 VDD2.n97 VSUBS 0.017191f
C1034 VDD2.n98 VSUBS 0.016236f
C1035 VDD2.n99 VSUBS 0.030215f
C1036 VDD2.n100 VSUBS 0.030215f
C1037 VDD2.n101 VSUBS 0.016236f
C1038 VDD2.n102 VSUBS 0.017191f
C1039 VDD2.n103 VSUBS 0.038376f
C1040 VDD2.n104 VSUBS 0.038376f
C1041 VDD2.n105 VSUBS 0.017191f
C1042 VDD2.n106 VSUBS 0.016236f
C1043 VDD2.n107 VSUBS 0.030215f
C1044 VDD2.n108 VSUBS 0.030215f
C1045 VDD2.n109 VSUBS 0.016236f
C1046 VDD2.n110 VSUBS 0.017191f
C1047 VDD2.n111 VSUBS 0.038376f
C1048 VDD2.n112 VSUBS 0.038376f
C1049 VDD2.n113 VSUBS 0.038376f
C1050 VDD2.n114 VSUBS 0.016713f
C1051 VDD2.n115 VSUBS 0.016236f
C1052 VDD2.n116 VSUBS 0.030215f
C1053 VDD2.n117 VSUBS 0.030215f
C1054 VDD2.n118 VSUBS 0.016236f
C1055 VDD2.n119 VSUBS 0.017191f
C1056 VDD2.n120 VSUBS 0.038376f
C1057 VDD2.n121 VSUBS 0.038376f
C1058 VDD2.n122 VSUBS 0.017191f
C1059 VDD2.n123 VSUBS 0.016236f
C1060 VDD2.n124 VSUBS 0.030215f
C1061 VDD2.n125 VSUBS 0.030215f
C1062 VDD2.n126 VSUBS 0.016236f
C1063 VDD2.n127 VSUBS 0.017191f
C1064 VDD2.n128 VSUBS 0.038376f
C1065 VDD2.n129 VSUBS 0.093783f
C1066 VDD2.n130 VSUBS 0.017191f
C1067 VDD2.n131 VSUBS 0.016236f
C1068 VDD2.n132 VSUBS 0.071078f
C1069 VDD2.n133 VSUBS 0.068092f
C1070 VDD2.n134 VSUBS 3.58303f
C1071 VDD2.t3 VSUBS 0.290099f
C1072 VDD2.t8 VSUBS 0.290099f
C1073 VDD2.n135 VSUBS 2.27044f
C1074 VDD2.n136 VSUBS 0.896627f
C1075 VDD2.t1 VSUBS 0.290099f
C1076 VDD2.t6 VSUBS 0.290099f
C1077 VDD2.n137 VSUBS 2.29652f
C1078 VN.t0 VSUBS 2.4921f
C1079 VN.n0 VSUBS 0.981181f
C1080 VN.n1 VSUBS 0.027266f
C1081 VN.n2 VSUBS 0.049232f
C1082 VN.n3 VSUBS 0.027266f
C1083 VN.t7 VSUBS 2.4921f
C1084 VN.n4 VSUBS 0.050817f
C1085 VN.n5 VSUBS 0.027266f
C1086 VN.n6 VSUBS 0.038273f
C1087 VN.n7 VSUBS 0.027266f
C1088 VN.n8 VSUBS 0.036387f
C1089 VN.n9 VSUBS 0.286732f
C1090 VN.t4 VSUBS 2.4921f
C1091 VN.t5 VSUBS 2.73556f
C1092 VN.n10 VSUBS 0.935407f
C1093 VN.n11 VSUBS 0.96673f
C1094 VN.n12 VSUBS 0.042789f
C1095 VN.n13 VSUBS 0.050817f
C1096 VN.n14 VSUBS 0.027266f
C1097 VN.n15 VSUBS 0.027266f
C1098 VN.n16 VSUBS 0.027266f
C1099 VN.n17 VSUBS 0.043225f
C1100 VN.n18 VSUBS 0.050817f
C1101 VN.t2 VSUBS 2.4921f
C1102 VN.n19 VSUBS 0.879223f
C1103 VN.n20 VSUBS 0.038273f
C1104 VN.n21 VSUBS 0.027266f
C1105 VN.n22 VSUBS 0.027266f
C1106 VN.n23 VSUBS 0.027266f
C1107 VN.n24 VSUBS 0.050817f
C1108 VN.n25 VSUBS 0.043225f
C1109 VN.n26 VSUBS 0.036387f
C1110 VN.n27 VSUBS 0.027266f
C1111 VN.n28 VSUBS 0.027266f
C1112 VN.n29 VSUBS 0.027266f
C1113 VN.n30 VSUBS 0.042789f
C1114 VN.n31 VSUBS 0.879223f
C1115 VN.n32 VSUBS 0.033757f
C1116 VN.n33 VSUBS 0.050817f
C1117 VN.n34 VSUBS 0.027266f
C1118 VN.n35 VSUBS 0.027266f
C1119 VN.n36 VSUBS 0.027266f
C1120 VN.n37 VSUBS 0.027056f
C1121 VN.n38 VSUBS 0.054141f
C1122 VN.n39 VSUBS 0.047305f
C1123 VN.n40 VSUBS 0.044007f
C1124 VN.n41 VSUBS 0.053392f
C1125 VN.t9 VSUBS 2.4921f
C1126 VN.n42 VSUBS 0.981181f
C1127 VN.n43 VSUBS 0.027266f
C1128 VN.n44 VSUBS 0.049232f
C1129 VN.n45 VSUBS 0.027266f
C1130 VN.t6 VSUBS 2.4921f
C1131 VN.n46 VSUBS 0.050817f
C1132 VN.n47 VSUBS 0.027266f
C1133 VN.n48 VSUBS 0.038273f
C1134 VN.n49 VSUBS 0.027266f
C1135 VN.t1 VSUBS 2.4921f
C1136 VN.n50 VSUBS 0.879223f
C1137 VN.n51 VSUBS 0.036387f
C1138 VN.n52 VSUBS 0.286732f
C1139 VN.t8 VSUBS 2.4921f
C1140 VN.t3 VSUBS 2.73556f
C1141 VN.n53 VSUBS 0.935407f
C1142 VN.n54 VSUBS 0.96673f
C1143 VN.n55 VSUBS 0.042789f
C1144 VN.n56 VSUBS 0.050817f
C1145 VN.n57 VSUBS 0.027266f
C1146 VN.n58 VSUBS 0.027266f
C1147 VN.n59 VSUBS 0.027266f
C1148 VN.n60 VSUBS 0.043225f
C1149 VN.n61 VSUBS 0.050817f
C1150 VN.n62 VSUBS 0.038273f
C1151 VN.n63 VSUBS 0.027266f
C1152 VN.n64 VSUBS 0.027266f
C1153 VN.n65 VSUBS 0.027266f
C1154 VN.n66 VSUBS 0.050817f
C1155 VN.n67 VSUBS 0.043225f
C1156 VN.n68 VSUBS 0.036387f
C1157 VN.n69 VSUBS 0.027266f
C1158 VN.n70 VSUBS 0.027266f
C1159 VN.n71 VSUBS 0.027266f
C1160 VN.n72 VSUBS 0.042789f
C1161 VN.n73 VSUBS 0.879223f
C1162 VN.n74 VSUBS 0.033757f
C1163 VN.n75 VSUBS 0.050817f
C1164 VN.n76 VSUBS 0.027266f
C1165 VN.n77 VSUBS 0.027266f
C1166 VN.n78 VSUBS 0.027266f
C1167 VN.n79 VSUBS 0.027056f
C1168 VN.n80 VSUBS 0.054141f
C1169 VN.n81 VSUBS 0.047305f
C1170 VN.n82 VSUBS 0.044007f
C1171 VN.n83 VSUBS 1.733f
C1172 VTAIL.t6 VSUBS 0.278775f
C1173 VTAIL.t18 VSUBS 0.278775f
C1174 VTAIL.n0 VSUBS 2.02606f
C1175 VTAIL.n1 VSUBS 1.02186f
C1176 VTAIL.n2 VSUBS 0.032151f
C1177 VTAIL.n3 VSUBS 0.029035f
C1178 VTAIL.n4 VSUBS 0.015602f
C1179 VTAIL.n5 VSUBS 0.036878f
C1180 VTAIL.n6 VSUBS 0.01652f
C1181 VTAIL.n7 VSUBS 0.029035f
C1182 VTAIL.n8 VSUBS 0.015602f
C1183 VTAIL.n9 VSUBS 0.036878f
C1184 VTAIL.n10 VSUBS 0.01652f
C1185 VTAIL.n11 VSUBS 0.029035f
C1186 VTAIL.n12 VSUBS 0.016061f
C1187 VTAIL.n13 VSUBS 0.036878f
C1188 VTAIL.n14 VSUBS 0.01652f
C1189 VTAIL.n15 VSUBS 0.029035f
C1190 VTAIL.n16 VSUBS 0.015602f
C1191 VTAIL.n17 VSUBS 0.036878f
C1192 VTAIL.n18 VSUBS 0.01652f
C1193 VTAIL.n19 VSUBS 0.029035f
C1194 VTAIL.n20 VSUBS 0.015602f
C1195 VTAIL.n21 VSUBS 0.027659f
C1196 VTAIL.n22 VSUBS 0.027742f
C1197 VTAIL.t13 VSUBS 0.079483f
C1198 VTAIL.n23 VSUBS 0.230638f
C1199 VTAIL.n24 VSUBS 1.44567f
C1200 VTAIL.n25 VSUBS 0.015602f
C1201 VTAIL.n26 VSUBS 0.01652f
C1202 VTAIL.n27 VSUBS 0.036878f
C1203 VTAIL.n28 VSUBS 0.036878f
C1204 VTAIL.n29 VSUBS 0.01652f
C1205 VTAIL.n30 VSUBS 0.015602f
C1206 VTAIL.n31 VSUBS 0.029035f
C1207 VTAIL.n32 VSUBS 0.029035f
C1208 VTAIL.n33 VSUBS 0.015602f
C1209 VTAIL.n34 VSUBS 0.01652f
C1210 VTAIL.n35 VSUBS 0.036878f
C1211 VTAIL.n36 VSUBS 0.036878f
C1212 VTAIL.n37 VSUBS 0.01652f
C1213 VTAIL.n38 VSUBS 0.015602f
C1214 VTAIL.n39 VSUBS 0.029035f
C1215 VTAIL.n40 VSUBS 0.029035f
C1216 VTAIL.n41 VSUBS 0.015602f
C1217 VTAIL.n42 VSUBS 0.015602f
C1218 VTAIL.n43 VSUBS 0.01652f
C1219 VTAIL.n44 VSUBS 0.036878f
C1220 VTAIL.n45 VSUBS 0.036878f
C1221 VTAIL.n46 VSUBS 0.036878f
C1222 VTAIL.n47 VSUBS 0.016061f
C1223 VTAIL.n48 VSUBS 0.015602f
C1224 VTAIL.n49 VSUBS 0.029035f
C1225 VTAIL.n50 VSUBS 0.029035f
C1226 VTAIL.n51 VSUBS 0.015602f
C1227 VTAIL.n52 VSUBS 0.01652f
C1228 VTAIL.n53 VSUBS 0.036878f
C1229 VTAIL.n54 VSUBS 0.036878f
C1230 VTAIL.n55 VSUBS 0.01652f
C1231 VTAIL.n56 VSUBS 0.015602f
C1232 VTAIL.n57 VSUBS 0.029035f
C1233 VTAIL.n58 VSUBS 0.029035f
C1234 VTAIL.n59 VSUBS 0.015602f
C1235 VTAIL.n60 VSUBS 0.01652f
C1236 VTAIL.n61 VSUBS 0.036878f
C1237 VTAIL.n62 VSUBS 0.090122f
C1238 VTAIL.n63 VSUBS 0.01652f
C1239 VTAIL.n64 VSUBS 0.015602f
C1240 VTAIL.n65 VSUBS 0.068303f
C1241 VTAIL.n66 VSUBS 0.045395f
C1242 VTAIL.n67 VSUBS 0.443253f
C1243 VTAIL.t12 VSUBS 0.278775f
C1244 VTAIL.t17 VSUBS 0.278775f
C1245 VTAIL.n68 VSUBS 2.02606f
C1246 VTAIL.n69 VSUBS 1.15937f
C1247 VTAIL.t16 VSUBS 0.278775f
C1248 VTAIL.t15 VSUBS 0.278775f
C1249 VTAIL.n70 VSUBS 2.02606f
C1250 VTAIL.n71 VSUBS 2.78293f
C1251 VTAIL.t1 VSUBS 0.278775f
C1252 VTAIL.t4 VSUBS 0.278775f
C1253 VTAIL.n72 VSUBS 2.02608f
C1254 VTAIL.n73 VSUBS 2.78292f
C1255 VTAIL.t7 VSUBS 0.278775f
C1256 VTAIL.t5 VSUBS 0.278775f
C1257 VTAIL.n74 VSUBS 2.02608f
C1258 VTAIL.n75 VSUBS 1.15936f
C1259 VTAIL.n76 VSUBS 0.032151f
C1260 VTAIL.n77 VSUBS 0.029035f
C1261 VTAIL.n78 VSUBS 0.015602f
C1262 VTAIL.n79 VSUBS 0.036878f
C1263 VTAIL.n80 VSUBS 0.01652f
C1264 VTAIL.n81 VSUBS 0.029035f
C1265 VTAIL.n82 VSUBS 0.015602f
C1266 VTAIL.n83 VSUBS 0.036878f
C1267 VTAIL.n84 VSUBS 0.01652f
C1268 VTAIL.n85 VSUBS 0.029035f
C1269 VTAIL.n86 VSUBS 0.016061f
C1270 VTAIL.n87 VSUBS 0.036878f
C1271 VTAIL.n88 VSUBS 0.015602f
C1272 VTAIL.n89 VSUBS 0.01652f
C1273 VTAIL.n90 VSUBS 0.029035f
C1274 VTAIL.n91 VSUBS 0.015602f
C1275 VTAIL.n92 VSUBS 0.036878f
C1276 VTAIL.n93 VSUBS 0.01652f
C1277 VTAIL.n94 VSUBS 0.029035f
C1278 VTAIL.n95 VSUBS 0.015602f
C1279 VTAIL.n96 VSUBS 0.027659f
C1280 VTAIL.n97 VSUBS 0.027742f
C1281 VTAIL.t19 VSUBS 0.079483f
C1282 VTAIL.n98 VSUBS 0.230638f
C1283 VTAIL.n99 VSUBS 1.44567f
C1284 VTAIL.n100 VSUBS 0.015602f
C1285 VTAIL.n101 VSUBS 0.01652f
C1286 VTAIL.n102 VSUBS 0.036878f
C1287 VTAIL.n103 VSUBS 0.036878f
C1288 VTAIL.n104 VSUBS 0.01652f
C1289 VTAIL.n105 VSUBS 0.015602f
C1290 VTAIL.n106 VSUBS 0.029035f
C1291 VTAIL.n107 VSUBS 0.029035f
C1292 VTAIL.n108 VSUBS 0.015602f
C1293 VTAIL.n109 VSUBS 0.01652f
C1294 VTAIL.n110 VSUBS 0.036878f
C1295 VTAIL.n111 VSUBS 0.036878f
C1296 VTAIL.n112 VSUBS 0.01652f
C1297 VTAIL.n113 VSUBS 0.015602f
C1298 VTAIL.n114 VSUBS 0.029035f
C1299 VTAIL.n115 VSUBS 0.029035f
C1300 VTAIL.n116 VSUBS 0.015602f
C1301 VTAIL.n117 VSUBS 0.01652f
C1302 VTAIL.n118 VSUBS 0.036878f
C1303 VTAIL.n119 VSUBS 0.036878f
C1304 VTAIL.n120 VSUBS 0.036878f
C1305 VTAIL.n121 VSUBS 0.016061f
C1306 VTAIL.n122 VSUBS 0.015602f
C1307 VTAIL.n123 VSUBS 0.029035f
C1308 VTAIL.n124 VSUBS 0.029035f
C1309 VTAIL.n125 VSUBS 0.015602f
C1310 VTAIL.n126 VSUBS 0.01652f
C1311 VTAIL.n127 VSUBS 0.036878f
C1312 VTAIL.n128 VSUBS 0.036878f
C1313 VTAIL.n129 VSUBS 0.01652f
C1314 VTAIL.n130 VSUBS 0.015602f
C1315 VTAIL.n131 VSUBS 0.029035f
C1316 VTAIL.n132 VSUBS 0.029035f
C1317 VTAIL.n133 VSUBS 0.015602f
C1318 VTAIL.n134 VSUBS 0.01652f
C1319 VTAIL.n135 VSUBS 0.036878f
C1320 VTAIL.n136 VSUBS 0.090122f
C1321 VTAIL.n137 VSUBS 0.01652f
C1322 VTAIL.n138 VSUBS 0.015602f
C1323 VTAIL.n139 VSUBS 0.068303f
C1324 VTAIL.n140 VSUBS 0.045395f
C1325 VTAIL.n141 VSUBS 0.443253f
C1326 VTAIL.t9 VSUBS 0.278775f
C1327 VTAIL.t14 VSUBS 0.278775f
C1328 VTAIL.n142 VSUBS 2.02608f
C1329 VTAIL.n143 VSUBS 1.07871f
C1330 VTAIL.t11 VSUBS 0.278775f
C1331 VTAIL.t10 VSUBS 0.278775f
C1332 VTAIL.n144 VSUBS 2.02608f
C1333 VTAIL.n145 VSUBS 1.15936f
C1334 VTAIL.n146 VSUBS 0.032151f
C1335 VTAIL.n147 VSUBS 0.029035f
C1336 VTAIL.n148 VSUBS 0.015602f
C1337 VTAIL.n149 VSUBS 0.036878f
C1338 VTAIL.n150 VSUBS 0.01652f
C1339 VTAIL.n151 VSUBS 0.029035f
C1340 VTAIL.n152 VSUBS 0.015602f
C1341 VTAIL.n153 VSUBS 0.036878f
C1342 VTAIL.n154 VSUBS 0.01652f
C1343 VTAIL.n155 VSUBS 0.029035f
C1344 VTAIL.n156 VSUBS 0.016061f
C1345 VTAIL.n157 VSUBS 0.036878f
C1346 VTAIL.n158 VSUBS 0.015602f
C1347 VTAIL.n159 VSUBS 0.01652f
C1348 VTAIL.n160 VSUBS 0.029035f
C1349 VTAIL.n161 VSUBS 0.015602f
C1350 VTAIL.n162 VSUBS 0.036878f
C1351 VTAIL.n163 VSUBS 0.01652f
C1352 VTAIL.n164 VSUBS 0.029035f
C1353 VTAIL.n165 VSUBS 0.015602f
C1354 VTAIL.n166 VSUBS 0.027659f
C1355 VTAIL.n167 VSUBS 0.027742f
C1356 VTAIL.t8 VSUBS 0.079483f
C1357 VTAIL.n168 VSUBS 0.230638f
C1358 VTAIL.n169 VSUBS 1.44567f
C1359 VTAIL.n170 VSUBS 0.015602f
C1360 VTAIL.n171 VSUBS 0.01652f
C1361 VTAIL.n172 VSUBS 0.036878f
C1362 VTAIL.n173 VSUBS 0.036878f
C1363 VTAIL.n174 VSUBS 0.01652f
C1364 VTAIL.n175 VSUBS 0.015602f
C1365 VTAIL.n176 VSUBS 0.029035f
C1366 VTAIL.n177 VSUBS 0.029035f
C1367 VTAIL.n178 VSUBS 0.015602f
C1368 VTAIL.n179 VSUBS 0.01652f
C1369 VTAIL.n180 VSUBS 0.036878f
C1370 VTAIL.n181 VSUBS 0.036878f
C1371 VTAIL.n182 VSUBS 0.01652f
C1372 VTAIL.n183 VSUBS 0.015602f
C1373 VTAIL.n184 VSUBS 0.029035f
C1374 VTAIL.n185 VSUBS 0.029035f
C1375 VTAIL.n186 VSUBS 0.015602f
C1376 VTAIL.n187 VSUBS 0.01652f
C1377 VTAIL.n188 VSUBS 0.036878f
C1378 VTAIL.n189 VSUBS 0.036878f
C1379 VTAIL.n190 VSUBS 0.036878f
C1380 VTAIL.n191 VSUBS 0.016061f
C1381 VTAIL.n192 VSUBS 0.015602f
C1382 VTAIL.n193 VSUBS 0.029035f
C1383 VTAIL.n194 VSUBS 0.029035f
C1384 VTAIL.n195 VSUBS 0.015602f
C1385 VTAIL.n196 VSUBS 0.01652f
C1386 VTAIL.n197 VSUBS 0.036878f
C1387 VTAIL.n198 VSUBS 0.036878f
C1388 VTAIL.n199 VSUBS 0.01652f
C1389 VTAIL.n200 VSUBS 0.015602f
C1390 VTAIL.n201 VSUBS 0.029035f
C1391 VTAIL.n202 VSUBS 0.029035f
C1392 VTAIL.n203 VSUBS 0.015602f
C1393 VTAIL.n204 VSUBS 0.01652f
C1394 VTAIL.n205 VSUBS 0.036878f
C1395 VTAIL.n206 VSUBS 0.090122f
C1396 VTAIL.n207 VSUBS 0.01652f
C1397 VTAIL.n208 VSUBS 0.015602f
C1398 VTAIL.n209 VSUBS 0.068303f
C1399 VTAIL.n210 VSUBS 0.045395f
C1400 VTAIL.n211 VSUBS 1.89825f
C1401 VTAIL.n212 VSUBS 0.032151f
C1402 VTAIL.n213 VSUBS 0.029035f
C1403 VTAIL.n214 VSUBS 0.015602f
C1404 VTAIL.n215 VSUBS 0.036878f
C1405 VTAIL.n216 VSUBS 0.01652f
C1406 VTAIL.n217 VSUBS 0.029035f
C1407 VTAIL.n218 VSUBS 0.015602f
C1408 VTAIL.n219 VSUBS 0.036878f
C1409 VTAIL.n220 VSUBS 0.01652f
C1410 VTAIL.n221 VSUBS 0.029035f
C1411 VTAIL.n222 VSUBS 0.016061f
C1412 VTAIL.n223 VSUBS 0.036878f
C1413 VTAIL.n224 VSUBS 0.01652f
C1414 VTAIL.n225 VSUBS 0.029035f
C1415 VTAIL.n226 VSUBS 0.015602f
C1416 VTAIL.n227 VSUBS 0.036878f
C1417 VTAIL.n228 VSUBS 0.01652f
C1418 VTAIL.n229 VSUBS 0.029035f
C1419 VTAIL.n230 VSUBS 0.015602f
C1420 VTAIL.n231 VSUBS 0.027659f
C1421 VTAIL.n232 VSUBS 0.027742f
C1422 VTAIL.t2 VSUBS 0.079483f
C1423 VTAIL.n233 VSUBS 0.230638f
C1424 VTAIL.n234 VSUBS 1.44567f
C1425 VTAIL.n235 VSUBS 0.015602f
C1426 VTAIL.n236 VSUBS 0.01652f
C1427 VTAIL.n237 VSUBS 0.036878f
C1428 VTAIL.n238 VSUBS 0.036878f
C1429 VTAIL.n239 VSUBS 0.01652f
C1430 VTAIL.n240 VSUBS 0.015602f
C1431 VTAIL.n241 VSUBS 0.029035f
C1432 VTAIL.n242 VSUBS 0.029035f
C1433 VTAIL.n243 VSUBS 0.015602f
C1434 VTAIL.n244 VSUBS 0.01652f
C1435 VTAIL.n245 VSUBS 0.036878f
C1436 VTAIL.n246 VSUBS 0.036878f
C1437 VTAIL.n247 VSUBS 0.01652f
C1438 VTAIL.n248 VSUBS 0.015602f
C1439 VTAIL.n249 VSUBS 0.029035f
C1440 VTAIL.n250 VSUBS 0.029035f
C1441 VTAIL.n251 VSUBS 0.015602f
C1442 VTAIL.n252 VSUBS 0.015602f
C1443 VTAIL.n253 VSUBS 0.01652f
C1444 VTAIL.n254 VSUBS 0.036878f
C1445 VTAIL.n255 VSUBS 0.036878f
C1446 VTAIL.n256 VSUBS 0.036878f
C1447 VTAIL.n257 VSUBS 0.016061f
C1448 VTAIL.n258 VSUBS 0.015602f
C1449 VTAIL.n259 VSUBS 0.029035f
C1450 VTAIL.n260 VSUBS 0.029035f
C1451 VTAIL.n261 VSUBS 0.015602f
C1452 VTAIL.n262 VSUBS 0.01652f
C1453 VTAIL.n263 VSUBS 0.036878f
C1454 VTAIL.n264 VSUBS 0.036878f
C1455 VTAIL.n265 VSUBS 0.01652f
C1456 VTAIL.n266 VSUBS 0.015602f
C1457 VTAIL.n267 VSUBS 0.029035f
C1458 VTAIL.n268 VSUBS 0.029035f
C1459 VTAIL.n269 VSUBS 0.015602f
C1460 VTAIL.n270 VSUBS 0.01652f
C1461 VTAIL.n271 VSUBS 0.036878f
C1462 VTAIL.n272 VSUBS 0.090122f
C1463 VTAIL.n273 VSUBS 0.01652f
C1464 VTAIL.n274 VSUBS 0.015602f
C1465 VTAIL.n275 VSUBS 0.068303f
C1466 VTAIL.n276 VSUBS 0.045395f
C1467 VTAIL.n277 VSUBS 1.89825f
C1468 VTAIL.t0 VSUBS 0.278775f
C1469 VTAIL.t3 VSUBS 0.278775f
C1470 VTAIL.n278 VSUBS 2.02606f
C1471 VTAIL.n279 VSUBS 0.967016f
C1472 VDD1.n0 VSUBS 0.033557f
C1473 VDD1.n1 VSUBS 0.030305f
C1474 VDD1.n2 VSUBS 0.016284f
C1475 VDD1.n3 VSUBS 0.038491f
C1476 VDD1.n4 VSUBS 0.017242f
C1477 VDD1.n5 VSUBS 0.030305f
C1478 VDD1.n6 VSUBS 0.016284f
C1479 VDD1.n7 VSUBS 0.038491f
C1480 VDD1.n8 VSUBS 0.017242f
C1481 VDD1.n9 VSUBS 0.030305f
C1482 VDD1.n10 VSUBS 0.016763f
C1483 VDD1.n11 VSUBS 0.038491f
C1484 VDD1.n12 VSUBS 0.016284f
C1485 VDD1.n13 VSUBS 0.017242f
C1486 VDD1.n14 VSUBS 0.030305f
C1487 VDD1.n15 VSUBS 0.016284f
C1488 VDD1.n16 VSUBS 0.038491f
C1489 VDD1.n17 VSUBS 0.017242f
C1490 VDD1.n18 VSUBS 0.030305f
C1491 VDD1.n19 VSUBS 0.016284f
C1492 VDD1.n20 VSUBS 0.028868f
C1493 VDD1.n21 VSUBS 0.028955f
C1494 VDD1.t5 VSUBS 0.082959f
C1495 VDD1.n22 VSUBS 0.240724f
C1496 VDD1.n23 VSUBS 1.50889f
C1497 VDD1.n24 VSUBS 0.016284f
C1498 VDD1.n25 VSUBS 0.017242f
C1499 VDD1.n26 VSUBS 0.038491f
C1500 VDD1.n27 VSUBS 0.038491f
C1501 VDD1.n28 VSUBS 0.017242f
C1502 VDD1.n29 VSUBS 0.016284f
C1503 VDD1.n30 VSUBS 0.030305f
C1504 VDD1.n31 VSUBS 0.030305f
C1505 VDD1.n32 VSUBS 0.016284f
C1506 VDD1.n33 VSUBS 0.017242f
C1507 VDD1.n34 VSUBS 0.038491f
C1508 VDD1.n35 VSUBS 0.038491f
C1509 VDD1.n36 VSUBS 0.017242f
C1510 VDD1.n37 VSUBS 0.016284f
C1511 VDD1.n38 VSUBS 0.030305f
C1512 VDD1.n39 VSUBS 0.030305f
C1513 VDD1.n40 VSUBS 0.016284f
C1514 VDD1.n41 VSUBS 0.017242f
C1515 VDD1.n42 VSUBS 0.038491f
C1516 VDD1.n43 VSUBS 0.038491f
C1517 VDD1.n44 VSUBS 0.038491f
C1518 VDD1.n45 VSUBS 0.016763f
C1519 VDD1.n46 VSUBS 0.016284f
C1520 VDD1.n47 VSUBS 0.030305f
C1521 VDD1.n48 VSUBS 0.030305f
C1522 VDD1.n49 VSUBS 0.016284f
C1523 VDD1.n50 VSUBS 0.017242f
C1524 VDD1.n51 VSUBS 0.038491f
C1525 VDD1.n52 VSUBS 0.038491f
C1526 VDD1.n53 VSUBS 0.017242f
C1527 VDD1.n54 VSUBS 0.016284f
C1528 VDD1.n55 VSUBS 0.030305f
C1529 VDD1.n56 VSUBS 0.030305f
C1530 VDD1.n57 VSUBS 0.016284f
C1531 VDD1.n58 VSUBS 0.017242f
C1532 VDD1.n59 VSUBS 0.038491f
C1533 VDD1.n60 VSUBS 0.094063f
C1534 VDD1.n61 VSUBS 0.017242f
C1535 VDD1.n62 VSUBS 0.016284f
C1536 VDD1.n63 VSUBS 0.07129f
C1537 VDD1.n64 VSUBS 0.084612f
C1538 VDD1.t8 VSUBS 0.290965f
C1539 VDD1.t1 VSUBS 0.290965f
C1540 VDD1.n65 VSUBS 2.27721f
C1541 VDD1.n66 VSUBS 1.20217f
C1542 VDD1.n67 VSUBS 0.033557f
C1543 VDD1.n68 VSUBS 0.030305f
C1544 VDD1.n69 VSUBS 0.016284f
C1545 VDD1.n70 VSUBS 0.038491f
C1546 VDD1.n71 VSUBS 0.017242f
C1547 VDD1.n72 VSUBS 0.030305f
C1548 VDD1.n73 VSUBS 0.016284f
C1549 VDD1.n74 VSUBS 0.038491f
C1550 VDD1.n75 VSUBS 0.017242f
C1551 VDD1.n76 VSUBS 0.030305f
C1552 VDD1.n77 VSUBS 0.016763f
C1553 VDD1.n78 VSUBS 0.038491f
C1554 VDD1.n79 VSUBS 0.017242f
C1555 VDD1.n80 VSUBS 0.030305f
C1556 VDD1.n81 VSUBS 0.016284f
C1557 VDD1.n82 VSUBS 0.038491f
C1558 VDD1.n83 VSUBS 0.017242f
C1559 VDD1.n84 VSUBS 0.030305f
C1560 VDD1.n85 VSUBS 0.016284f
C1561 VDD1.n86 VSUBS 0.028868f
C1562 VDD1.n87 VSUBS 0.028955f
C1563 VDD1.t6 VSUBS 0.082959f
C1564 VDD1.n88 VSUBS 0.240724f
C1565 VDD1.n89 VSUBS 1.50889f
C1566 VDD1.n90 VSUBS 0.016284f
C1567 VDD1.n91 VSUBS 0.017242f
C1568 VDD1.n92 VSUBS 0.038491f
C1569 VDD1.n93 VSUBS 0.038491f
C1570 VDD1.n94 VSUBS 0.017242f
C1571 VDD1.n95 VSUBS 0.016284f
C1572 VDD1.n96 VSUBS 0.030305f
C1573 VDD1.n97 VSUBS 0.030305f
C1574 VDD1.n98 VSUBS 0.016284f
C1575 VDD1.n99 VSUBS 0.017242f
C1576 VDD1.n100 VSUBS 0.038491f
C1577 VDD1.n101 VSUBS 0.038491f
C1578 VDD1.n102 VSUBS 0.017242f
C1579 VDD1.n103 VSUBS 0.016284f
C1580 VDD1.n104 VSUBS 0.030305f
C1581 VDD1.n105 VSUBS 0.030305f
C1582 VDD1.n106 VSUBS 0.016284f
C1583 VDD1.n107 VSUBS 0.016284f
C1584 VDD1.n108 VSUBS 0.017242f
C1585 VDD1.n109 VSUBS 0.038491f
C1586 VDD1.n110 VSUBS 0.038491f
C1587 VDD1.n111 VSUBS 0.038491f
C1588 VDD1.n112 VSUBS 0.016763f
C1589 VDD1.n113 VSUBS 0.016284f
C1590 VDD1.n114 VSUBS 0.030305f
C1591 VDD1.n115 VSUBS 0.030305f
C1592 VDD1.n116 VSUBS 0.016284f
C1593 VDD1.n117 VSUBS 0.017242f
C1594 VDD1.n118 VSUBS 0.038491f
C1595 VDD1.n119 VSUBS 0.038491f
C1596 VDD1.n120 VSUBS 0.017242f
C1597 VDD1.n121 VSUBS 0.016284f
C1598 VDD1.n122 VSUBS 0.030305f
C1599 VDD1.n123 VSUBS 0.030305f
C1600 VDD1.n124 VSUBS 0.016284f
C1601 VDD1.n125 VSUBS 0.017242f
C1602 VDD1.n126 VSUBS 0.038491f
C1603 VDD1.n127 VSUBS 0.094063f
C1604 VDD1.n128 VSUBS 0.017242f
C1605 VDD1.n129 VSUBS 0.016284f
C1606 VDD1.n130 VSUBS 0.07129f
C1607 VDD1.n131 VSUBS 0.084612f
C1608 VDD1.t9 VSUBS 0.290965f
C1609 VDD1.t2 VSUBS 0.290965f
C1610 VDD1.n132 VSUBS 2.2772f
C1611 VDD1.n133 VSUBS 1.19224f
C1612 VDD1.t7 VSUBS 0.290965f
C1613 VDD1.t3 VSUBS 0.290965f
C1614 VDD1.n134 VSUBS 2.30343f
C1615 VDD1.n135 VSUBS 4.1056f
C1616 VDD1.t0 VSUBS 0.290965f
C1617 VDD1.t4 VSUBS 0.290965f
C1618 VDD1.n136 VSUBS 2.2772f
C1619 VDD1.n137 VSUBS 4.25972f
C1620 VP.t4 VSUBS 2.70581f
C1621 VP.n0 VSUBS 1.06532f
C1622 VP.n1 VSUBS 0.029604f
C1623 VP.n2 VSUBS 0.053454f
C1624 VP.n3 VSUBS 0.029604f
C1625 VP.t0 VSUBS 2.70581f
C1626 VP.n4 VSUBS 0.055175f
C1627 VP.n5 VSUBS 0.029604f
C1628 VP.n6 VSUBS 0.041555f
C1629 VP.n7 VSUBS 0.029604f
C1630 VP.n8 VSUBS 0.039507f
C1631 VP.n9 VSUBS 0.029604f
C1632 VP.t2 VSUBS 2.70581f
C1633 VP.n10 VSUBS 0.055175f
C1634 VP.n11 VSUBS 0.029604f
C1635 VP.n12 VSUBS 0.051361f
C1636 VP.t9 VSUBS 2.70581f
C1637 VP.n13 VSUBS 1.06532f
C1638 VP.n14 VSUBS 0.029604f
C1639 VP.n15 VSUBS 0.053454f
C1640 VP.n16 VSUBS 0.029604f
C1641 VP.t7 VSUBS 2.70581f
C1642 VP.n17 VSUBS 0.055175f
C1643 VP.n18 VSUBS 0.029604f
C1644 VP.n19 VSUBS 0.041555f
C1645 VP.n20 VSUBS 0.029604f
C1646 VP.n21 VSUBS 0.039507f
C1647 VP.n22 VSUBS 0.311321f
C1648 VP.t3 VSUBS 2.70581f
C1649 VP.t8 VSUBS 2.97014f
C1650 VP.n23 VSUBS 1.01562f
C1651 VP.n24 VSUBS 1.04963f
C1652 VP.n25 VSUBS 0.046458f
C1653 VP.n26 VSUBS 0.055175f
C1654 VP.n27 VSUBS 0.029604f
C1655 VP.n28 VSUBS 0.029604f
C1656 VP.n29 VSUBS 0.029604f
C1657 VP.n30 VSUBS 0.046932f
C1658 VP.n31 VSUBS 0.055175f
C1659 VP.t6 VSUBS 2.70581f
C1660 VP.n32 VSUBS 0.95462f
C1661 VP.n33 VSUBS 0.041555f
C1662 VP.n34 VSUBS 0.029604f
C1663 VP.n35 VSUBS 0.029604f
C1664 VP.n36 VSUBS 0.029604f
C1665 VP.n37 VSUBS 0.055175f
C1666 VP.n38 VSUBS 0.046932f
C1667 VP.n39 VSUBS 0.039507f
C1668 VP.n40 VSUBS 0.029604f
C1669 VP.n41 VSUBS 0.029604f
C1670 VP.n42 VSUBS 0.029604f
C1671 VP.n43 VSUBS 0.046458f
C1672 VP.n44 VSUBS 0.95462f
C1673 VP.n45 VSUBS 0.036651f
C1674 VP.n46 VSUBS 0.055175f
C1675 VP.n47 VSUBS 0.029604f
C1676 VP.n48 VSUBS 0.029604f
C1677 VP.n49 VSUBS 0.029604f
C1678 VP.n50 VSUBS 0.029376f
C1679 VP.n51 VSUBS 0.058784f
C1680 VP.n52 VSUBS 0.051361f
C1681 VP.n53 VSUBS 0.04778f
C1682 VP.n54 VSUBS 1.86981f
C1683 VP.t1 VSUBS 2.70581f
C1684 VP.n55 VSUBS 1.06532f
C1685 VP.n56 VSUBS 1.88945f
C1686 VP.n57 VSUBS 0.04778f
C1687 VP.n58 VSUBS 0.029604f
C1688 VP.n59 VSUBS 0.058784f
C1689 VP.n60 VSUBS 0.029376f
C1690 VP.n61 VSUBS 0.053454f
C1691 VP.n62 VSUBS 0.029604f
C1692 VP.n63 VSUBS 0.029604f
C1693 VP.n64 VSUBS 0.029604f
C1694 VP.n65 VSUBS 0.036651f
C1695 VP.n66 VSUBS 0.95462f
C1696 VP.n67 VSUBS 0.046458f
C1697 VP.n68 VSUBS 0.055175f
C1698 VP.n69 VSUBS 0.029604f
C1699 VP.n70 VSUBS 0.029604f
C1700 VP.n71 VSUBS 0.029604f
C1701 VP.n72 VSUBS 0.046932f
C1702 VP.n73 VSUBS 0.055175f
C1703 VP.t5 VSUBS 2.70581f
C1704 VP.n74 VSUBS 0.95462f
C1705 VP.n75 VSUBS 0.041555f
C1706 VP.n76 VSUBS 0.029604f
C1707 VP.n77 VSUBS 0.029604f
C1708 VP.n78 VSUBS 0.029604f
C1709 VP.n79 VSUBS 0.055175f
C1710 VP.n80 VSUBS 0.046932f
C1711 VP.n81 VSUBS 0.039507f
C1712 VP.n82 VSUBS 0.029604f
C1713 VP.n83 VSUBS 0.029604f
C1714 VP.n84 VSUBS 0.029604f
C1715 VP.n85 VSUBS 0.046458f
C1716 VP.n86 VSUBS 0.95462f
C1717 VP.n87 VSUBS 0.036651f
C1718 VP.n88 VSUBS 0.055175f
C1719 VP.n89 VSUBS 0.029604f
C1720 VP.n90 VSUBS 0.029604f
C1721 VP.n91 VSUBS 0.029604f
C1722 VP.n92 VSUBS 0.029376f
C1723 VP.n93 VSUBS 0.058784f
C1724 VP.n94 VSUBS 0.051361f
C1725 VP.n95 VSUBS 0.04778f
C1726 VP.n96 VSUBS 0.057971f
.ends

