* NGSPICE file created from diff_pair_sample_0484.ext - technology: sky130A

.subckt diff_pair_sample_0484 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.72
X1 VDD1.t5 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0.6633 ps=4.35 w=4.02 l=3.72
X2 VDD1.t4 VP.t1 VTAIL.t7 B.t19 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0.6633 ps=4.35 w=4.02 l=3.72
X3 VDD1.t3 VP.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=1.5678 ps=8.82 w=4.02 l=3.72
X4 VTAIL.t10 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=0.6633 ps=4.35 w=4.02 l=3.72
X5 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.72
X6 VTAIL.t9 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=0.6633 ps=4.35 w=4.02 l=3.72
X7 VDD2.t5 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0.6633 ps=4.35 w=4.02 l=3.72
X8 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=1.5678 ps=8.82 w=4.02 l=3.72
X9 VDD2.t3 VN.t2 VTAIL.t3 B.t19 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0.6633 ps=4.35 w=4.02 l=3.72
X10 VTAIL.t5 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=0.6633 ps=4.35 w=4.02 l=3.72
X11 VDD1.t0 VP.t5 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=1.5678 ps=8.82 w=4.02 l=3.72
X12 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.72
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.72
X14 VDD2.t1 VN.t4 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=1.5678 ps=8.82 w=4.02 l=3.72
X15 VTAIL.t0 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6633 pd=4.35 as=0.6633 ps=4.35 w=4.02 l=3.72
R0 B.n682 B.n681 585
R1 B.n217 B.n125 585
R2 B.n216 B.n215 585
R3 B.n214 B.n213 585
R4 B.n212 B.n211 585
R5 B.n210 B.n209 585
R6 B.n208 B.n207 585
R7 B.n206 B.n205 585
R8 B.n204 B.n203 585
R9 B.n202 B.n201 585
R10 B.n200 B.n199 585
R11 B.n198 B.n197 585
R12 B.n196 B.n195 585
R13 B.n194 B.n193 585
R14 B.n192 B.n191 585
R15 B.n190 B.n189 585
R16 B.n188 B.n187 585
R17 B.n186 B.n185 585
R18 B.n184 B.n183 585
R19 B.n182 B.n181 585
R20 B.n180 B.n179 585
R21 B.n178 B.n177 585
R22 B.n176 B.n175 585
R23 B.n174 B.n173 585
R24 B.n172 B.n171 585
R25 B.n170 B.n169 585
R26 B.n168 B.n167 585
R27 B.n166 B.n165 585
R28 B.n164 B.n163 585
R29 B.n162 B.n161 585
R30 B.n160 B.n159 585
R31 B.n158 B.n157 585
R32 B.n156 B.n155 585
R33 B.n154 B.n153 585
R34 B.n152 B.n151 585
R35 B.n150 B.n149 585
R36 B.n148 B.n147 585
R37 B.n146 B.n145 585
R38 B.n144 B.n143 585
R39 B.n142 B.n141 585
R40 B.n140 B.n139 585
R41 B.n138 B.n137 585
R42 B.n136 B.n135 585
R43 B.n134 B.n133 585
R44 B.n103 B.n102 585
R45 B.n687 B.n686 585
R46 B.n680 B.n126 585
R47 B.n126 B.n100 585
R48 B.n679 B.n99 585
R49 B.n691 B.n99 585
R50 B.n678 B.n98 585
R51 B.n692 B.n98 585
R52 B.n677 B.n97 585
R53 B.n693 B.n97 585
R54 B.n676 B.n675 585
R55 B.n675 B.n93 585
R56 B.n674 B.n92 585
R57 B.n699 B.n92 585
R58 B.n673 B.n91 585
R59 B.n700 B.n91 585
R60 B.n672 B.n90 585
R61 B.n701 B.n90 585
R62 B.n671 B.n670 585
R63 B.n670 B.n86 585
R64 B.n669 B.n85 585
R65 B.t10 B.n85 585
R66 B.n668 B.n84 585
R67 B.n707 B.n84 585
R68 B.n667 B.n83 585
R69 B.n708 B.n83 585
R70 B.n666 B.n665 585
R71 B.n665 B.n79 585
R72 B.n664 B.n78 585
R73 B.n714 B.n78 585
R74 B.n663 B.n77 585
R75 B.n715 B.n77 585
R76 B.n662 B.n76 585
R77 B.n716 B.n76 585
R78 B.n661 B.n660 585
R79 B.n660 B.n72 585
R80 B.n659 B.n71 585
R81 B.n722 B.n71 585
R82 B.n658 B.n70 585
R83 B.n723 B.n70 585
R84 B.n657 B.n69 585
R85 B.n724 B.n69 585
R86 B.n656 B.n655 585
R87 B.n655 B.n65 585
R88 B.n654 B.n64 585
R89 B.n730 B.n64 585
R90 B.n653 B.n63 585
R91 B.n731 B.n63 585
R92 B.n652 B.n62 585
R93 B.n732 B.n62 585
R94 B.n651 B.n650 585
R95 B.n650 B.n61 585
R96 B.n649 B.n57 585
R97 B.n738 B.n57 585
R98 B.n648 B.n56 585
R99 B.n739 B.n56 585
R100 B.n647 B.n55 585
R101 B.n740 B.n55 585
R102 B.n646 B.n645 585
R103 B.n645 B.n51 585
R104 B.n644 B.n50 585
R105 B.n746 B.n50 585
R106 B.n643 B.n49 585
R107 B.n747 B.n49 585
R108 B.n642 B.n48 585
R109 B.n748 B.n48 585
R110 B.n641 B.n640 585
R111 B.n640 B.n44 585
R112 B.n639 B.n43 585
R113 B.n754 B.n43 585
R114 B.n638 B.n42 585
R115 B.n755 B.n42 585
R116 B.n637 B.n41 585
R117 B.n756 B.n41 585
R118 B.n636 B.n635 585
R119 B.n635 B.n40 585
R120 B.n634 B.n36 585
R121 B.n762 B.n36 585
R122 B.n633 B.n35 585
R123 B.n763 B.n35 585
R124 B.n632 B.n34 585
R125 B.n764 B.n34 585
R126 B.n631 B.n630 585
R127 B.n630 B.n30 585
R128 B.n629 B.n29 585
R129 B.n770 B.n29 585
R130 B.n628 B.n28 585
R131 B.n771 B.n28 585
R132 B.n627 B.n27 585
R133 B.n772 B.n27 585
R134 B.n626 B.n625 585
R135 B.n625 B.n23 585
R136 B.n624 B.n22 585
R137 B.n778 B.n22 585
R138 B.n623 B.n21 585
R139 B.n779 B.n21 585
R140 B.n622 B.n20 585
R141 B.n780 B.n20 585
R142 B.n621 B.n620 585
R143 B.n620 B.n16 585
R144 B.n619 B.n15 585
R145 B.n786 B.n15 585
R146 B.n618 B.n14 585
R147 B.n787 B.n14 585
R148 B.n617 B.n13 585
R149 B.n788 B.n13 585
R150 B.n616 B.n615 585
R151 B.n615 B.n12 585
R152 B.n614 B.n613 585
R153 B.n614 B.n8 585
R154 B.n612 B.n7 585
R155 B.n795 B.n7 585
R156 B.n611 B.n6 585
R157 B.n796 B.n6 585
R158 B.n610 B.n5 585
R159 B.n797 B.n5 585
R160 B.n609 B.n608 585
R161 B.n608 B.n4 585
R162 B.n607 B.n218 585
R163 B.n607 B.n606 585
R164 B.n597 B.n219 585
R165 B.n220 B.n219 585
R166 B.n599 B.n598 585
R167 B.n600 B.n599 585
R168 B.n596 B.n225 585
R169 B.n225 B.n224 585
R170 B.n595 B.n594 585
R171 B.n594 B.n593 585
R172 B.n227 B.n226 585
R173 B.n228 B.n227 585
R174 B.n586 B.n585 585
R175 B.n587 B.n586 585
R176 B.n584 B.n233 585
R177 B.n233 B.n232 585
R178 B.n583 B.n582 585
R179 B.n582 B.n581 585
R180 B.n235 B.n234 585
R181 B.n236 B.n235 585
R182 B.n574 B.n573 585
R183 B.n575 B.n574 585
R184 B.n572 B.n241 585
R185 B.n241 B.n240 585
R186 B.n571 B.n570 585
R187 B.n570 B.n569 585
R188 B.n243 B.n242 585
R189 B.n244 B.n243 585
R190 B.n562 B.n561 585
R191 B.n563 B.n562 585
R192 B.n560 B.n249 585
R193 B.n249 B.n248 585
R194 B.n559 B.n558 585
R195 B.n558 B.n557 585
R196 B.n251 B.n250 585
R197 B.n550 B.n251 585
R198 B.n549 B.n548 585
R199 B.n551 B.n549 585
R200 B.n547 B.n256 585
R201 B.n256 B.n255 585
R202 B.n546 B.n545 585
R203 B.n545 B.n544 585
R204 B.n258 B.n257 585
R205 B.n259 B.n258 585
R206 B.n537 B.n536 585
R207 B.n538 B.n537 585
R208 B.n535 B.n264 585
R209 B.n264 B.n263 585
R210 B.n534 B.n533 585
R211 B.n533 B.n532 585
R212 B.n266 B.n265 585
R213 B.n267 B.n266 585
R214 B.n525 B.n524 585
R215 B.n526 B.n525 585
R216 B.n523 B.n272 585
R217 B.n272 B.n271 585
R218 B.n522 B.n521 585
R219 B.n521 B.n520 585
R220 B.n274 B.n273 585
R221 B.n513 B.n274 585
R222 B.n512 B.n511 585
R223 B.n514 B.n512 585
R224 B.n510 B.n279 585
R225 B.n279 B.n278 585
R226 B.n509 B.n508 585
R227 B.n508 B.n507 585
R228 B.n281 B.n280 585
R229 B.n282 B.n281 585
R230 B.n500 B.n499 585
R231 B.n501 B.n500 585
R232 B.n498 B.n287 585
R233 B.n287 B.n286 585
R234 B.n497 B.n496 585
R235 B.n496 B.n495 585
R236 B.n289 B.n288 585
R237 B.n290 B.n289 585
R238 B.n488 B.n487 585
R239 B.n489 B.n488 585
R240 B.n486 B.n295 585
R241 B.n295 B.n294 585
R242 B.n485 B.n484 585
R243 B.n484 B.n483 585
R244 B.n297 B.n296 585
R245 B.n298 B.n297 585
R246 B.n476 B.n475 585
R247 B.n477 B.n476 585
R248 B.n474 B.n303 585
R249 B.n303 B.n302 585
R250 B.n473 B.n472 585
R251 B.n472 B.t6 585
R252 B.n305 B.n304 585
R253 B.n306 B.n305 585
R254 B.n465 B.n464 585
R255 B.n466 B.n465 585
R256 B.n463 B.n311 585
R257 B.n311 B.n310 585
R258 B.n462 B.n461 585
R259 B.n461 B.n460 585
R260 B.n313 B.n312 585
R261 B.n314 B.n313 585
R262 B.n453 B.n452 585
R263 B.n454 B.n453 585
R264 B.n451 B.n319 585
R265 B.n319 B.n318 585
R266 B.n450 B.n449 585
R267 B.n449 B.n448 585
R268 B.n321 B.n320 585
R269 B.n322 B.n321 585
R270 B.n444 B.n443 585
R271 B.n325 B.n324 585
R272 B.n440 B.n439 585
R273 B.n441 B.n440 585
R274 B.n438 B.n348 585
R275 B.n437 B.n436 585
R276 B.n435 B.n434 585
R277 B.n433 B.n432 585
R278 B.n431 B.n430 585
R279 B.n429 B.n428 585
R280 B.n427 B.n426 585
R281 B.n425 B.n424 585
R282 B.n423 B.n422 585
R283 B.n421 B.n420 585
R284 B.n419 B.n418 585
R285 B.n417 B.n416 585
R286 B.n415 B.n414 585
R287 B.n413 B.n412 585
R288 B.n411 B.n410 585
R289 B.n408 B.n407 585
R290 B.n406 B.n405 585
R291 B.n404 B.n403 585
R292 B.n402 B.n401 585
R293 B.n400 B.n399 585
R294 B.n398 B.n397 585
R295 B.n396 B.n395 585
R296 B.n394 B.n393 585
R297 B.n392 B.n391 585
R298 B.n390 B.n389 585
R299 B.n387 B.n386 585
R300 B.n385 B.n384 585
R301 B.n383 B.n382 585
R302 B.n381 B.n380 585
R303 B.n379 B.n378 585
R304 B.n377 B.n376 585
R305 B.n375 B.n374 585
R306 B.n373 B.n372 585
R307 B.n371 B.n370 585
R308 B.n369 B.n368 585
R309 B.n367 B.n366 585
R310 B.n365 B.n364 585
R311 B.n363 B.n362 585
R312 B.n361 B.n360 585
R313 B.n359 B.n358 585
R314 B.n357 B.n356 585
R315 B.n355 B.n354 585
R316 B.n353 B.n347 585
R317 B.n441 B.n347 585
R318 B.n445 B.n323 585
R319 B.n323 B.n322 585
R320 B.n447 B.n446 585
R321 B.n448 B.n447 585
R322 B.n317 B.n316 585
R323 B.n318 B.n317 585
R324 B.n456 B.n455 585
R325 B.n455 B.n454 585
R326 B.n457 B.n315 585
R327 B.n315 B.n314 585
R328 B.n459 B.n458 585
R329 B.n460 B.n459 585
R330 B.n309 B.n308 585
R331 B.n310 B.n309 585
R332 B.n468 B.n467 585
R333 B.n467 B.n466 585
R334 B.n469 B.n307 585
R335 B.n307 B.n306 585
R336 B.n471 B.n470 585
R337 B.t6 B.n471 585
R338 B.n301 B.n300 585
R339 B.n302 B.n301 585
R340 B.n479 B.n478 585
R341 B.n478 B.n477 585
R342 B.n480 B.n299 585
R343 B.n299 B.n298 585
R344 B.n482 B.n481 585
R345 B.n483 B.n482 585
R346 B.n293 B.n292 585
R347 B.n294 B.n293 585
R348 B.n491 B.n490 585
R349 B.n490 B.n489 585
R350 B.n492 B.n291 585
R351 B.n291 B.n290 585
R352 B.n494 B.n493 585
R353 B.n495 B.n494 585
R354 B.n285 B.n284 585
R355 B.n286 B.n285 585
R356 B.n503 B.n502 585
R357 B.n502 B.n501 585
R358 B.n504 B.n283 585
R359 B.n283 B.n282 585
R360 B.n506 B.n505 585
R361 B.n507 B.n506 585
R362 B.n277 B.n276 585
R363 B.n278 B.n277 585
R364 B.n516 B.n515 585
R365 B.n515 B.n514 585
R366 B.n517 B.n275 585
R367 B.n513 B.n275 585
R368 B.n519 B.n518 585
R369 B.n520 B.n519 585
R370 B.n270 B.n269 585
R371 B.n271 B.n270 585
R372 B.n528 B.n527 585
R373 B.n527 B.n526 585
R374 B.n529 B.n268 585
R375 B.n268 B.n267 585
R376 B.n531 B.n530 585
R377 B.n532 B.n531 585
R378 B.n262 B.n261 585
R379 B.n263 B.n262 585
R380 B.n540 B.n539 585
R381 B.n539 B.n538 585
R382 B.n541 B.n260 585
R383 B.n260 B.n259 585
R384 B.n543 B.n542 585
R385 B.n544 B.n543 585
R386 B.n254 B.n253 585
R387 B.n255 B.n254 585
R388 B.n553 B.n552 585
R389 B.n552 B.n551 585
R390 B.n554 B.n252 585
R391 B.n550 B.n252 585
R392 B.n556 B.n555 585
R393 B.n557 B.n556 585
R394 B.n247 B.n246 585
R395 B.n248 B.n247 585
R396 B.n565 B.n564 585
R397 B.n564 B.n563 585
R398 B.n566 B.n245 585
R399 B.n245 B.n244 585
R400 B.n568 B.n567 585
R401 B.n569 B.n568 585
R402 B.n239 B.n238 585
R403 B.n240 B.n239 585
R404 B.n577 B.n576 585
R405 B.n576 B.n575 585
R406 B.n578 B.n237 585
R407 B.n237 B.n236 585
R408 B.n580 B.n579 585
R409 B.n581 B.n580 585
R410 B.n231 B.n230 585
R411 B.n232 B.n231 585
R412 B.n589 B.n588 585
R413 B.n588 B.n587 585
R414 B.n590 B.n229 585
R415 B.n229 B.n228 585
R416 B.n592 B.n591 585
R417 B.n593 B.n592 585
R418 B.n223 B.n222 585
R419 B.n224 B.n223 585
R420 B.n602 B.n601 585
R421 B.n601 B.n600 585
R422 B.n603 B.n221 585
R423 B.n221 B.n220 585
R424 B.n605 B.n604 585
R425 B.n606 B.n605 585
R426 B.n3 B.n0 585
R427 B.n4 B.n3 585
R428 B.n794 B.n1 585
R429 B.n795 B.n794 585
R430 B.n793 B.n792 585
R431 B.n793 B.n8 585
R432 B.n791 B.n9 585
R433 B.n12 B.n9 585
R434 B.n790 B.n789 585
R435 B.n789 B.n788 585
R436 B.n11 B.n10 585
R437 B.n787 B.n11 585
R438 B.n785 B.n784 585
R439 B.n786 B.n785 585
R440 B.n783 B.n17 585
R441 B.n17 B.n16 585
R442 B.n782 B.n781 585
R443 B.n781 B.n780 585
R444 B.n19 B.n18 585
R445 B.n779 B.n19 585
R446 B.n777 B.n776 585
R447 B.n778 B.n777 585
R448 B.n775 B.n24 585
R449 B.n24 B.n23 585
R450 B.n774 B.n773 585
R451 B.n773 B.n772 585
R452 B.n26 B.n25 585
R453 B.n771 B.n26 585
R454 B.n769 B.n768 585
R455 B.n770 B.n769 585
R456 B.n767 B.n31 585
R457 B.n31 B.n30 585
R458 B.n766 B.n765 585
R459 B.n765 B.n764 585
R460 B.n33 B.n32 585
R461 B.n763 B.n33 585
R462 B.n761 B.n760 585
R463 B.n762 B.n761 585
R464 B.n759 B.n37 585
R465 B.n40 B.n37 585
R466 B.n758 B.n757 585
R467 B.n757 B.n756 585
R468 B.n39 B.n38 585
R469 B.n755 B.n39 585
R470 B.n753 B.n752 585
R471 B.n754 B.n753 585
R472 B.n751 B.n45 585
R473 B.n45 B.n44 585
R474 B.n750 B.n749 585
R475 B.n749 B.n748 585
R476 B.n47 B.n46 585
R477 B.n747 B.n47 585
R478 B.n745 B.n744 585
R479 B.n746 B.n745 585
R480 B.n743 B.n52 585
R481 B.n52 B.n51 585
R482 B.n742 B.n741 585
R483 B.n741 B.n740 585
R484 B.n54 B.n53 585
R485 B.n739 B.n54 585
R486 B.n737 B.n736 585
R487 B.n738 B.n737 585
R488 B.n735 B.n58 585
R489 B.n61 B.n58 585
R490 B.n734 B.n733 585
R491 B.n733 B.n732 585
R492 B.n60 B.n59 585
R493 B.n731 B.n60 585
R494 B.n729 B.n728 585
R495 B.n730 B.n729 585
R496 B.n727 B.n66 585
R497 B.n66 B.n65 585
R498 B.n726 B.n725 585
R499 B.n725 B.n724 585
R500 B.n68 B.n67 585
R501 B.n723 B.n68 585
R502 B.n721 B.n720 585
R503 B.n722 B.n721 585
R504 B.n719 B.n73 585
R505 B.n73 B.n72 585
R506 B.n718 B.n717 585
R507 B.n717 B.n716 585
R508 B.n75 B.n74 585
R509 B.n715 B.n75 585
R510 B.n713 B.n712 585
R511 B.n714 B.n713 585
R512 B.n711 B.n80 585
R513 B.n80 B.n79 585
R514 B.n710 B.n709 585
R515 B.n709 B.n708 585
R516 B.n82 B.n81 585
R517 B.n707 B.n82 585
R518 B.n706 B.n705 585
R519 B.t10 B.n706 585
R520 B.n704 B.n87 585
R521 B.n87 B.n86 585
R522 B.n703 B.n702 585
R523 B.n702 B.n701 585
R524 B.n89 B.n88 585
R525 B.n700 B.n89 585
R526 B.n698 B.n697 585
R527 B.n699 B.n698 585
R528 B.n696 B.n94 585
R529 B.n94 B.n93 585
R530 B.n695 B.n694 585
R531 B.n694 B.n693 585
R532 B.n96 B.n95 585
R533 B.n692 B.n96 585
R534 B.n690 B.n689 585
R535 B.n691 B.n690 585
R536 B.n688 B.n101 585
R537 B.n101 B.n100 585
R538 B.n798 B.n797 585
R539 B.n796 B.n2 585
R540 B.n686 B.n101 530.939
R541 B.n682 B.n126 530.939
R542 B.n347 B.n321 530.939
R543 B.n443 B.n323 530.939
R544 B.n684 B.n683 256.663
R545 B.n684 B.n124 256.663
R546 B.n684 B.n123 256.663
R547 B.n684 B.n122 256.663
R548 B.n684 B.n121 256.663
R549 B.n684 B.n120 256.663
R550 B.n684 B.n119 256.663
R551 B.n684 B.n118 256.663
R552 B.n684 B.n117 256.663
R553 B.n684 B.n116 256.663
R554 B.n684 B.n115 256.663
R555 B.n684 B.n114 256.663
R556 B.n684 B.n113 256.663
R557 B.n684 B.n112 256.663
R558 B.n684 B.n111 256.663
R559 B.n684 B.n110 256.663
R560 B.n684 B.n109 256.663
R561 B.n684 B.n108 256.663
R562 B.n684 B.n107 256.663
R563 B.n684 B.n106 256.663
R564 B.n684 B.n105 256.663
R565 B.n684 B.n104 256.663
R566 B.n685 B.n684 256.663
R567 B.n442 B.n441 256.663
R568 B.n441 B.n326 256.663
R569 B.n441 B.n327 256.663
R570 B.n441 B.n328 256.663
R571 B.n441 B.n329 256.663
R572 B.n441 B.n330 256.663
R573 B.n441 B.n331 256.663
R574 B.n441 B.n332 256.663
R575 B.n441 B.n333 256.663
R576 B.n441 B.n334 256.663
R577 B.n441 B.n335 256.663
R578 B.n441 B.n336 256.663
R579 B.n441 B.n337 256.663
R580 B.n441 B.n338 256.663
R581 B.n441 B.n339 256.663
R582 B.n441 B.n340 256.663
R583 B.n441 B.n341 256.663
R584 B.n441 B.n342 256.663
R585 B.n441 B.n343 256.663
R586 B.n441 B.n344 256.663
R587 B.n441 B.n345 256.663
R588 B.n441 B.n346 256.663
R589 B.n800 B.n799 256.663
R590 B.n130 B.t13 235.325
R591 B.n127 B.t9 235.325
R592 B.n351 B.t5 235.325
R593 B.n349 B.t16 235.325
R594 B.n127 B.t11 224.194
R595 B.n351 B.t8 224.194
R596 B.n130 B.t14 224.194
R597 B.n349 B.t18 224.194
R598 B.n441 B.n322 166.864
R599 B.n684 B.n100 166.864
R600 B.n133 B.n103 163.367
R601 B.n137 B.n136 163.367
R602 B.n141 B.n140 163.367
R603 B.n145 B.n144 163.367
R604 B.n149 B.n148 163.367
R605 B.n153 B.n152 163.367
R606 B.n157 B.n156 163.367
R607 B.n161 B.n160 163.367
R608 B.n165 B.n164 163.367
R609 B.n169 B.n168 163.367
R610 B.n173 B.n172 163.367
R611 B.n177 B.n176 163.367
R612 B.n181 B.n180 163.367
R613 B.n185 B.n184 163.367
R614 B.n189 B.n188 163.367
R615 B.n193 B.n192 163.367
R616 B.n197 B.n196 163.367
R617 B.n201 B.n200 163.367
R618 B.n205 B.n204 163.367
R619 B.n209 B.n208 163.367
R620 B.n213 B.n212 163.367
R621 B.n215 B.n125 163.367
R622 B.n449 B.n321 163.367
R623 B.n449 B.n319 163.367
R624 B.n453 B.n319 163.367
R625 B.n453 B.n313 163.367
R626 B.n461 B.n313 163.367
R627 B.n461 B.n311 163.367
R628 B.n465 B.n311 163.367
R629 B.n465 B.n305 163.367
R630 B.n472 B.n305 163.367
R631 B.n472 B.n303 163.367
R632 B.n476 B.n303 163.367
R633 B.n476 B.n297 163.367
R634 B.n484 B.n297 163.367
R635 B.n484 B.n295 163.367
R636 B.n488 B.n295 163.367
R637 B.n488 B.n289 163.367
R638 B.n496 B.n289 163.367
R639 B.n496 B.n287 163.367
R640 B.n500 B.n287 163.367
R641 B.n500 B.n281 163.367
R642 B.n508 B.n281 163.367
R643 B.n508 B.n279 163.367
R644 B.n512 B.n279 163.367
R645 B.n512 B.n274 163.367
R646 B.n521 B.n274 163.367
R647 B.n521 B.n272 163.367
R648 B.n525 B.n272 163.367
R649 B.n525 B.n266 163.367
R650 B.n533 B.n266 163.367
R651 B.n533 B.n264 163.367
R652 B.n537 B.n264 163.367
R653 B.n537 B.n258 163.367
R654 B.n545 B.n258 163.367
R655 B.n545 B.n256 163.367
R656 B.n549 B.n256 163.367
R657 B.n549 B.n251 163.367
R658 B.n558 B.n251 163.367
R659 B.n558 B.n249 163.367
R660 B.n562 B.n249 163.367
R661 B.n562 B.n243 163.367
R662 B.n570 B.n243 163.367
R663 B.n570 B.n241 163.367
R664 B.n574 B.n241 163.367
R665 B.n574 B.n235 163.367
R666 B.n582 B.n235 163.367
R667 B.n582 B.n233 163.367
R668 B.n586 B.n233 163.367
R669 B.n586 B.n227 163.367
R670 B.n594 B.n227 163.367
R671 B.n594 B.n225 163.367
R672 B.n599 B.n225 163.367
R673 B.n599 B.n219 163.367
R674 B.n607 B.n219 163.367
R675 B.n608 B.n607 163.367
R676 B.n608 B.n5 163.367
R677 B.n6 B.n5 163.367
R678 B.n7 B.n6 163.367
R679 B.n614 B.n7 163.367
R680 B.n615 B.n614 163.367
R681 B.n615 B.n13 163.367
R682 B.n14 B.n13 163.367
R683 B.n15 B.n14 163.367
R684 B.n620 B.n15 163.367
R685 B.n620 B.n20 163.367
R686 B.n21 B.n20 163.367
R687 B.n22 B.n21 163.367
R688 B.n625 B.n22 163.367
R689 B.n625 B.n27 163.367
R690 B.n28 B.n27 163.367
R691 B.n29 B.n28 163.367
R692 B.n630 B.n29 163.367
R693 B.n630 B.n34 163.367
R694 B.n35 B.n34 163.367
R695 B.n36 B.n35 163.367
R696 B.n635 B.n36 163.367
R697 B.n635 B.n41 163.367
R698 B.n42 B.n41 163.367
R699 B.n43 B.n42 163.367
R700 B.n640 B.n43 163.367
R701 B.n640 B.n48 163.367
R702 B.n49 B.n48 163.367
R703 B.n50 B.n49 163.367
R704 B.n645 B.n50 163.367
R705 B.n645 B.n55 163.367
R706 B.n56 B.n55 163.367
R707 B.n57 B.n56 163.367
R708 B.n650 B.n57 163.367
R709 B.n650 B.n62 163.367
R710 B.n63 B.n62 163.367
R711 B.n64 B.n63 163.367
R712 B.n655 B.n64 163.367
R713 B.n655 B.n69 163.367
R714 B.n70 B.n69 163.367
R715 B.n71 B.n70 163.367
R716 B.n660 B.n71 163.367
R717 B.n660 B.n76 163.367
R718 B.n77 B.n76 163.367
R719 B.n78 B.n77 163.367
R720 B.n665 B.n78 163.367
R721 B.n665 B.n83 163.367
R722 B.n84 B.n83 163.367
R723 B.n85 B.n84 163.367
R724 B.n670 B.n85 163.367
R725 B.n670 B.n90 163.367
R726 B.n91 B.n90 163.367
R727 B.n92 B.n91 163.367
R728 B.n675 B.n92 163.367
R729 B.n675 B.n97 163.367
R730 B.n98 B.n97 163.367
R731 B.n99 B.n98 163.367
R732 B.n126 B.n99 163.367
R733 B.n440 B.n325 163.367
R734 B.n440 B.n348 163.367
R735 B.n436 B.n435 163.367
R736 B.n432 B.n431 163.367
R737 B.n428 B.n427 163.367
R738 B.n424 B.n423 163.367
R739 B.n420 B.n419 163.367
R740 B.n416 B.n415 163.367
R741 B.n412 B.n411 163.367
R742 B.n407 B.n406 163.367
R743 B.n403 B.n402 163.367
R744 B.n399 B.n398 163.367
R745 B.n395 B.n394 163.367
R746 B.n391 B.n390 163.367
R747 B.n386 B.n385 163.367
R748 B.n382 B.n381 163.367
R749 B.n378 B.n377 163.367
R750 B.n374 B.n373 163.367
R751 B.n370 B.n369 163.367
R752 B.n366 B.n365 163.367
R753 B.n362 B.n361 163.367
R754 B.n358 B.n357 163.367
R755 B.n354 B.n347 163.367
R756 B.n447 B.n323 163.367
R757 B.n447 B.n317 163.367
R758 B.n455 B.n317 163.367
R759 B.n455 B.n315 163.367
R760 B.n459 B.n315 163.367
R761 B.n459 B.n309 163.367
R762 B.n467 B.n309 163.367
R763 B.n467 B.n307 163.367
R764 B.n471 B.n307 163.367
R765 B.n471 B.n301 163.367
R766 B.n478 B.n301 163.367
R767 B.n478 B.n299 163.367
R768 B.n482 B.n299 163.367
R769 B.n482 B.n293 163.367
R770 B.n490 B.n293 163.367
R771 B.n490 B.n291 163.367
R772 B.n494 B.n291 163.367
R773 B.n494 B.n285 163.367
R774 B.n502 B.n285 163.367
R775 B.n502 B.n283 163.367
R776 B.n506 B.n283 163.367
R777 B.n506 B.n277 163.367
R778 B.n515 B.n277 163.367
R779 B.n515 B.n275 163.367
R780 B.n519 B.n275 163.367
R781 B.n519 B.n270 163.367
R782 B.n527 B.n270 163.367
R783 B.n527 B.n268 163.367
R784 B.n531 B.n268 163.367
R785 B.n531 B.n262 163.367
R786 B.n539 B.n262 163.367
R787 B.n539 B.n260 163.367
R788 B.n543 B.n260 163.367
R789 B.n543 B.n254 163.367
R790 B.n552 B.n254 163.367
R791 B.n552 B.n252 163.367
R792 B.n556 B.n252 163.367
R793 B.n556 B.n247 163.367
R794 B.n564 B.n247 163.367
R795 B.n564 B.n245 163.367
R796 B.n568 B.n245 163.367
R797 B.n568 B.n239 163.367
R798 B.n576 B.n239 163.367
R799 B.n576 B.n237 163.367
R800 B.n580 B.n237 163.367
R801 B.n580 B.n231 163.367
R802 B.n588 B.n231 163.367
R803 B.n588 B.n229 163.367
R804 B.n592 B.n229 163.367
R805 B.n592 B.n223 163.367
R806 B.n601 B.n223 163.367
R807 B.n601 B.n221 163.367
R808 B.n605 B.n221 163.367
R809 B.n605 B.n3 163.367
R810 B.n798 B.n3 163.367
R811 B.n794 B.n2 163.367
R812 B.n794 B.n793 163.367
R813 B.n793 B.n9 163.367
R814 B.n789 B.n9 163.367
R815 B.n789 B.n11 163.367
R816 B.n785 B.n11 163.367
R817 B.n785 B.n17 163.367
R818 B.n781 B.n17 163.367
R819 B.n781 B.n19 163.367
R820 B.n777 B.n19 163.367
R821 B.n777 B.n24 163.367
R822 B.n773 B.n24 163.367
R823 B.n773 B.n26 163.367
R824 B.n769 B.n26 163.367
R825 B.n769 B.n31 163.367
R826 B.n765 B.n31 163.367
R827 B.n765 B.n33 163.367
R828 B.n761 B.n33 163.367
R829 B.n761 B.n37 163.367
R830 B.n757 B.n37 163.367
R831 B.n757 B.n39 163.367
R832 B.n753 B.n39 163.367
R833 B.n753 B.n45 163.367
R834 B.n749 B.n45 163.367
R835 B.n749 B.n47 163.367
R836 B.n745 B.n47 163.367
R837 B.n745 B.n52 163.367
R838 B.n741 B.n52 163.367
R839 B.n741 B.n54 163.367
R840 B.n737 B.n54 163.367
R841 B.n737 B.n58 163.367
R842 B.n733 B.n58 163.367
R843 B.n733 B.n60 163.367
R844 B.n729 B.n60 163.367
R845 B.n729 B.n66 163.367
R846 B.n725 B.n66 163.367
R847 B.n725 B.n68 163.367
R848 B.n721 B.n68 163.367
R849 B.n721 B.n73 163.367
R850 B.n717 B.n73 163.367
R851 B.n717 B.n75 163.367
R852 B.n713 B.n75 163.367
R853 B.n713 B.n80 163.367
R854 B.n709 B.n80 163.367
R855 B.n709 B.n82 163.367
R856 B.n706 B.n82 163.367
R857 B.n706 B.n87 163.367
R858 B.n702 B.n87 163.367
R859 B.n702 B.n89 163.367
R860 B.n698 B.n89 163.367
R861 B.n698 B.n94 163.367
R862 B.n694 B.n94 163.367
R863 B.n694 B.n96 163.367
R864 B.n690 B.n96 163.367
R865 B.n690 B.n101 163.367
R866 B.n128 B.t12 145.649
R867 B.n352 B.t7 145.649
R868 B.n131 B.t15 145.649
R869 B.n350 B.t17 145.649
R870 B.n448 B.n322 80.4739
R871 B.n448 B.n318 80.4739
R872 B.n454 B.n318 80.4739
R873 B.n454 B.n314 80.4739
R874 B.n460 B.n314 80.4739
R875 B.n460 B.n310 80.4739
R876 B.n466 B.n310 80.4739
R877 B.n466 B.n306 80.4739
R878 B.t6 B.n306 80.4739
R879 B.t6 B.n302 80.4739
R880 B.n477 B.n302 80.4739
R881 B.n477 B.n298 80.4739
R882 B.n483 B.n298 80.4739
R883 B.n483 B.n294 80.4739
R884 B.n489 B.n294 80.4739
R885 B.n489 B.n290 80.4739
R886 B.n495 B.n290 80.4739
R887 B.n495 B.n286 80.4739
R888 B.n501 B.n286 80.4739
R889 B.n501 B.n282 80.4739
R890 B.n507 B.n282 80.4739
R891 B.n507 B.n278 80.4739
R892 B.n514 B.n278 80.4739
R893 B.n514 B.n513 80.4739
R894 B.n520 B.n271 80.4739
R895 B.n526 B.n271 80.4739
R896 B.n526 B.n267 80.4739
R897 B.n532 B.n267 80.4739
R898 B.n532 B.n263 80.4739
R899 B.n538 B.n263 80.4739
R900 B.n538 B.n259 80.4739
R901 B.n544 B.n259 80.4739
R902 B.n544 B.n255 80.4739
R903 B.n551 B.n255 80.4739
R904 B.n551 B.n550 80.4739
R905 B.n557 B.n248 80.4739
R906 B.n563 B.n248 80.4739
R907 B.n563 B.n244 80.4739
R908 B.n569 B.n244 80.4739
R909 B.n569 B.n240 80.4739
R910 B.n575 B.n240 80.4739
R911 B.n575 B.n236 80.4739
R912 B.n581 B.n236 80.4739
R913 B.n581 B.n232 80.4739
R914 B.n587 B.n232 80.4739
R915 B.n593 B.n228 80.4739
R916 B.n593 B.n224 80.4739
R917 B.n600 B.n224 80.4739
R918 B.n600 B.n220 80.4739
R919 B.n606 B.n220 80.4739
R920 B.n606 B.n4 80.4739
R921 B.n797 B.n4 80.4739
R922 B.n797 B.n796 80.4739
R923 B.n796 B.n795 80.4739
R924 B.n795 B.n8 80.4739
R925 B.n12 B.n8 80.4739
R926 B.n788 B.n12 80.4739
R927 B.n788 B.n787 80.4739
R928 B.n787 B.n786 80.4739
R929 B.n786 B.n16 80.4739
R930 B.n780 B.n779 80.4739
R931 B.n779 B.n778 80.4739
R932 B.n778 B.n23 80.4739
R933 B.n772 B.n23 80.4739
R934 B.n772 B.n771 80.4739
R935 B.n771 B.n770 80.4739
R936 B.n770 B.n30 80.4739
R937 B.n764 B.n30 80.4739
R938 B.n764 B.n763 80.4739
R939 B.n763 B.n762 80.4739
R940 B.n756 B.n40 80.4739
R941 B.n756 B.n755 80.4739
R942 B.n755 B.n754 80.4739
R943 B.n754 B.n44 80.4739
R944 B.n748 B.n44 80.4739
R945 B.n748 B.n747 80.4739
R946 B.n747 B.n746 80.4739
R947 B.n746 B.n51 80.4739
R948 B.n740 B.n51 80.4739
R949 B.n740 B.n739 80.4739
R950 B.n739 B.n738 80.4739
R951 B.n732 B.n61 80.4739
R952 B.n732 B.n731 80.4739
R953 B.n731 B.n730 80.4739
R954 B.n730 B.n65 80.4739
R955 B.n724 B.n65 80.4739
R956 B.n724 B.n723 80.4739
R957 B.n723 B.n722 80.4739
R958 B.n722 B.n72 80.4739
R959 B.n716 B.n72 80.4739
R960 B.n716 B.n715 80.4739
R961 B.n715 B.n714 80.4739
R962 B.n714 B.n79 80.4739
R963 B.n708 B.n79 80.4739
R964 B.n708 B.n707 80.4739
R965 B.n707 B.t10 80.4739
R966 B.t10 B.n86 80.4739
R967 B.n701 B.n86 80.4739
R968 B.n701 B.n700 80.4739
R969 B.n700 B.n699 80.4739
R970 B.n699 B.n93 80.4739
R971 B.n693 B.n93 80.4739
R972 B.n693 B.n692 80.4739
R973 B.n692 B.n691 80.4739
R974 B.n691 B.n100 80.4739
R975 B.n131 B.n130 78.546
R976 B.n128 B.n127 78.546
R977 B.n352 B.n351 78.546
R978 B.n350 B.n349 78.546
R979 B.n557 B.t3 78.107
R980 B.n762 B.t4 78.107
R981 B.n587 B.t1 75.7401
R982 B.n780 B.t19 75.7401
R983 B.n686 B.n685 71.676
R984 B.n133 B.n104 71.676
R985 B.n137 B.n105 71.676
R986 B.n141 B.n106 71.676
R987 B.n145 B.n107 71.676
R988 B.n149 B.n108 71.676
R989 B.n153 B.n109 71.676
R990 B.n157 B.n110 71.676
R991 B.n161 B.n111 71.676
R992 B.n165 B.n112 71.676
R993 B.n169 B.n113 71.676
R994 B.n173 B.n114 71.676
R995 B.n177 B.n115 71.676
R996 B.n181 B.n116 71.676
R997 B.n185 B.n117 71.676
R998 B.n189 B.n118 71.676
R999 B.n193 B.n119 71.676
R1000 B.n197 B.n120 71.676
R1001 B.n201 B.n121 71.676
R1002 B.n205 B.n122 71.676
R1003 B.n209 B.n123 71.676
R1004 B.n213 B.n124 71.676
R1005 B.n683 B.n125 71.676
R1006 B.n683 B.n682 71.676
R1007 B.n215 B.n124 71.676
R1008 B.n212 B.n123 71.676
R1009 B.n208 B.n122 71.676
R1010 B.n204 B.n121 71.676
R1011 B.n200 B.n120 71.676
R1012 B.n196 B.n119 71.676
R1013 B.n192 B.n118 71.676
R1014 B.n188 B.n117 71.676
R1015 B.n184 B.n116 71.676
R1016 B.n180 B.n115 71.676
R1017 B.n176 B.n114 71.676
R1018 B.n172 B.n113 71.676
R1019 B.n168 B.n112 71.676
R1020 B.n164 B.n111 71.676
R1021 B.n160 B.n110 71.676
R1022 B.n156 B.n109 71.676
R1023 B.n152 B.n108 71.676
R1024 B.n148 B.n107 71.676
R1025 B.n144 B.n106 71.676
R1026 B.n140 B.n105 71.676
R1027 B.n136 B.n104 71.676
R1028 B.n685 B.n103 71.676
R1029 B.n443 B.n442 71.676
R1030 B.n348 B.n326 71.676
R1031 B.n435 B.n327 71.676
R1032 B.n431 B.n328 71.676
R1033 B.n427 B.n329 71.676
R1034 B.n423 B.n330 71.676
R1035 B.n419 B.n331 71.676
R1036 B.n415 B.n332 71.676
R1037 B.n411 B.n333 71.676
R1038 B.n406 B.n334 71.676
R1039 B.n402 B.n335 71.676
R1040 B.n398 B.n336 71.676
R1041 B.n394 B.n337 71.676
R1042 B.n390 B.n338 71.676
R1043 B.n385 B.n339 71.676
R1044 B.n381 B.n340 71.676
R1045 B.n377 B.n341 71.676
R1046 B.n373 B.n342 71.676
R1047 B.n369 B.n343 71.676
R1048 B.n365 B.n344 71.676
R1049 B.n361 B.n345 71.676
R1050 B.n357 B.n346 71.676
R1051 B.n442 B.n325 71.676
R1052 B.n436 B.n326 71.676
R1053 B.n432 B.n327 71.676
R1054 B.n428 B.n328 71.676
R1055 B.n424 B.n329 71.676
R1056 B.n420 B.n330 71.676
R1057 B.n416 B.n331 71.676
R1058 B.n412 B.n332 71.676
R1059 B.n407 B.n333 71.676
R1060 B.n403 B.n334 71.676
R1061 B.n399 B.n335 71.676
R1062 B.n395 B.n336 71.676
R1063 B.n391 B.n337 71.676
R1064 B.n386 B.n338 71.676
R1065 B.n382 B.n339 71.676
R1066 B.n378 B.n340 71.676
R1067 B.n374 B.n341 71.676
R1068 B.n370 B.n342 71.676
R1069 B.n366 B.n343 71.676
R1070 B.n362 B.n344 71.676
R1071 B.n358 B.n345 71.676
R1072 B.n354 B.n346 71.676
R1073 B.n799 B.n798 71.676
R1074 B.n799 B.n2 71.676
R1075 B.n520 B.t0 71.0064
R1076 B.n738 B.t2 71.0064
R1077 B.n132 B.n131 59.5399
R1078 B.n129 B.n128 59.5399
R1079 B.n388 B.n352 59.5399
R1080 B.n409 B.n350 59.5399
R1081 B.n445 B.n444 34.4981
R1082 B.n353 B.n320 34.4981
R1083 B.n681 B.n680 34.4981
R1084 B.n688 B.n687 34.4981
R1085 B B.n800 18.0485
R1086 B.n446 B.n445 10.6151
R1087 B.n446 B.n316 10.6151
R1088 B.n456 B.n316 10.6151
R1089 B.n457 B.n456 10.6151
R1090 B.n458 B.n457 10.6151
R1091 B.n458 B.n308 10.6151
R1092 B.n468 B.n308 10.6151
R1093 B.n469 B.n468 10.6151
R1094 B.n470 B.n469 10.6151
R1095 B.n470 B.n300 10.6151
R1096 B.n479 B.n300 10.6151
R1097 B.n480 B.n479 10.6151
R1098 B.n481 B.n480 10.6151
R1099 B.n481 B.n292 10.6151
R1100 B.n491 B.n292 10.6151
R1101 B.n492 B.n491 10.6151
R1102 B.n493 B.n492 10.6151
R1103 B.n493 B.n284 10.6151
R1104 B.n503 B.n284 10.6151
R1105 B.n504 B.n503 10.6151
R1106 B.n505 B.n504 10.6151
R1107 B.n505 B.n276 10.6151
R1108 B.n516 B.n276 10.6151
R1109 B.n517 B.n516 10.6151
R1110 B.n518 B.n517 10.6151
R1111 B.n518 B.n269 10.6151
R1112 B.n528 B.n269 10.6151
R1113 B.n529 B.n528 10.6151
R1114 B.n530 B.n529 10.6151
R1115 B.n530 B.n261 10.6151
R1116 B.n540 B.n261 10.6151
R1117 B.n541 B.n540 10.6151
R1118 B.n542 B.n541 10.6151
R1119 B.n542 B.n253 10.6151
R1120 B.n553 B.n253 10.6151
R1121 B.n554 B.n553 10.6151
R1122 B.n555 B.n554 10.6151
R1123 B.n555 B.n246 10.6151
R1124 B.n565 B.n246 10.6151
R1125 B.n566 B.n565 10.6151
R1126 B.n567 B.n566 10.6151
R1127 B.n567 B.n238 10.6151
R1128 B.n577 B.n238 10.6151
R1129 B.n578 B.n577 10.6151
R1130 B.n579 B.n578 10.6151
R1131 B.n579 B.n230 10.6151
R1132 B.n589 B.n230 10.6151
R1133 B.n590 B.n589 10.6151
R1134 B.n591 B.n590 10.6151
R1135 B.n591 B.n222 10.6151
R1136 B.n602 B.n222 10.6151
R1137 B.n603 B.n602 10.6151
R1138 B.n604 B.n603 10.6151
R1139 B.n604 B.n0 10.6151
R1140 B.n444 B.n324 10.6151
R1141 B.n439 B.n324 10.6151
R1142 B.n439 B.n438 10.6151
R1143 B.n438 B.n437 10.6151
R1144 B.n437 B.n434 10.6151
R1145 B.n434 B.n433 10.6151
R1146 B.n433 B.n430 10.6151
R1147 B.n430 B.n429 10.6151
R1148 B.n429 B.n426 10.6151
R1149 B.n426 B.n425 10.6151
R1150 B.n425 B.n422 10.6151
R1151 B.n422 B.n421 10.6151
R1152 B.n421 B.n418 10.6151
R1153 B.n418 B.n417 10.6151
R1154 B.n417 B.n414 10.6151
R1155 B.n414 B.n413 10.6151
R1156 B.n413 B.n410 10.6151
R1157 B.n408 B.n405 10.6151
R1158 B.n405 B.n404 10.6151
R1159 B.n404 B.n401 10.6151
R1160 B.n401 B.n400 10.6151
R1161 B.n400 B.n397 10.6151
R1162 B.n397 B.n396 10.6151
R1163 B.n396 B.n393 10.6151
R1164 B.n393 B.n392 10.6151
R1165 B.n392 B.n389 10.6151
R1166 B.n387 B.n384 10.6151
R1167 B.n384 B.n383 10.6151
R1168 B.n383 B.n380 10.6151
R1169 B.n380 B.n379 10.6151
R1170 B.n379 B.n376 10.6151
R1171 B.n376 B.n375 10.6151
R1172 B.n375 B.n372 10.6151
R1173 B.n372 B.n371 10.6151
R1174 B.n371 B.n368 10.6151
R1175 B.n368 B.n367 10.6151
R1176 B.n367 B.n364 10.6151
R1177 B.n364 B.n363 10.6151
R1178 B.n363 B.n360 10.6151
R1179 B.n360 B.n359 10.6151
R1180 B.n359 B.n356 10.6151
R1181 B.n356 B.n355 10.6151
R1182 B.n355 B.n353 10.6151
R1183 B.n450 B.n320 10.6151
R1184 B.n451 B.n450 10.6151
R1185 B.n452 B.n451 10.6151
R1186 B.n452 B.n312 10.6151
R1187 B.n462 B.n312 10.6151
R1188 B.n463 B.n462 10.6151
R1189 B.n464 B.n463 10.6151
R1190 B.n464 B.n304 10.6151
R1191 B.n473 B.n304 10.6151
R1192 B.n474 B.n473 10.6151
R1193 B.n475 B.n474 10.6151
R1194 B.n475 B.n296 10.6151
R1195 B.n485 B.n296 10.6151
R1196 B.n486 B.n485 10.6151
R1197 B.n487 B.n486 10.6151
R1198 B.n487 B.n288 10.6151
R1199 B.n497 B.n288 10.6151
R1200 B.n498 B.n497 10.6151
R1201 B.n499 B.n498 10.6151
R1202 B.n499 B.n280 10.6151
R1203 B.n509 B.n280 10.6151
R1204 B.n510 B.n509 10.6151
R1205 B.n511 B.n510 10.6151
R1206 B.n511 B.n273 10.6151
R1207 B.n522 B.n273 10.6151
R1208 B.n523 B.n522 10.6151
R1209 B.n524 B.n523 10.6151
R1210 B.n524 B.n265 10.6151
R1211 B.n534 B.n265 10.6151
R1212 B.n535 B.n534 10.6151
R1213 B.n536 B.n535 10.6151
R1214 B.n536 B.n257 10.6151
R1215 B.n546 B.n257 10.6151
R1216 B.n547 B.n546 10.6151
R1217 B.n548 B.n547 10.6151
R1218 B.n548 B.n250 10.6151
R1219 B.n559 B.n250 10.6151
R1220 B.n560 B.n559 10.6151
R1221 B.n561 B.n560 10.6151
R1222 B.n561 B.n242 10.6151
R1223 B.n571 B.n242 10.6151
R1224 B.n572 B.n571 10.6151
R1225 B.n573 B.n572 10.6151
R1226 B.n573 B.n234 10.6151
R1227 B.n583 B.n234 10.6151
R1228 B.n584 B.n583 10.6151
R1229 B.n585 B.n584 10.6151
R1230 B.n585 B.n226 10.6151
R1231 B.n595 B.n226 10.6151
R1232 B.n596 B.n595 10.6151
R1233 B.n598 B.n596 10.6151
R1234 B.n598 B.n597 10.6151
R1235 B.n597 B.n218 10.6151
R1236 B.n609 B.n218 10.6151
R1237 B.n610 B.n609 10.6151
R1238 B.n611 B.n610 10.6151
R1239 B.n612 B.n611 10.6151
R1240 B.n613 B.n612 10.6151
R1241 B.n616 B.n613 10.6151
R1242 B.n617 B.n616 10.6151
R1243 B.n618 B.n617 10.6151
R1244 B.n619 B.n618 10.6151
R1245 B.n621 B.n619 10.6151
R1246 B.n622 B.n621 10.6151
R1247 B.n623 B.n622 10.6151
R1248 B.n624 B.n623 10.6151
R1249 B.n626 B.n624 10.6151
R1250 B.n627 B.n626 10.6151
R1251 B.n628 B.n627 10.6151
R1252 B.n629 B.n628 10.6151
R1253 B.n631 B.n629 10.6151
R1254 B.n632 B.n631 10.6151
R1255 B.n633 B.n632 10.6151
R1256 B.n634 B.n633 10.6151
R1257 B.n636 B.n634 10.6151
R1258 B.n637 B.n636 10.6151
R1259 B.n638 B.n637 10.6151
R1260 B.n639 B.n638 10.6151
R1261 B.n641 B.n639 10.6151
R1262 B.n642 B.n641 10.6151
R1263 B.n643 B.n642 10.6151
R1264 B.n644 B.n643 10.6151
R1265 B.n646 B.n644 10.6151
R1266 B.n647 B.n646 10.6151
R1267 B.n648 B.n647 10.6151
R1268 B.n649 B.n648 10.6151
R1269 B.n651 B.n649 10.6151
R1270 B.n652 B.n651 10.6151
R1271 B.n653 B.n652 10.6151
R1272 B.n654 B.n653 10.6151
R1273 B.n656 B.n654 10.6151
R1274 B.n657 B.n656 10.6151
R1275 B.n658 B.n657 10.6151
R1276 B.n659 B.n658 10.6151
R1277 B.n661 B.n659 10.6151
R1278 B.n662 B.n661 10.6151
R1279 B.n663 B.n662 10.6151
R1280 B.n664 B.n663 10.6151
R1281 B.n666 B.n664 10.6151
R1282 B.n667 B.n666 10.6151
R1283 B.n668 B.n667 10.6151
R1284 B.n669 B.n668 10.6151
R1285 B.n671 B.n669 10.6151
R1286 B.n672 B.n671 10.6151
R1287 B.n673 B.n672 10.6151
R1288 B.n674 B.n673 10.6151
R1289 B.n676 B.n674 10.6151
R1290 B.n677 B.n676 10.6151
R1291 B.n678 B.n677 10.6151
R1292 B.n679 B.n678 10.6151
R1293 B.n680 B.n679 10.6151
R1294 B.n792 B.n1 10.6151
R1295 B.n792 B.n791 10.6151
R1296 B.n791 B.n790 10.6151
R1297 B.n790 B.n10 10.6151
R1298 B.n784 B.n10 10.6151
R1299 B.n784 B.n783 10.6151
R1300 B.n783 B.n782 10.6151
R1301 B.n782 B.n18 10.6151
R1302 B.n776 B.n18 10.6151
R1303 B.n776 B.n775 10.6151
R1304 B.n775 B.n774 10.6151
R1305 B.n774 B.n25 10.6151
R1306 B.n768 B.n25 10.6151
R1307 B.n768 B.n767 10.6151
R1308 B.n767 B.n766 10.6151
R1309 B.n766 B.n32 10.6151
R1310 B.n760 B.n32 10.6151
R1311 B.n760 B.n759 10.6151
R1312 B.n759 B.n758 10.6151
R1313 B.n758 B.n38 10.6151
R1314 B.n752 B.n38 10.6151
R1315 B.n752 B.n751 10.6151
R1316 B.n751 B.n750 10.6151
R1317 B.n750 B.n46 10.6151
R1318 B.n744 B.n46 10.6151
R1319 B.n744 B.n743 10.6151
R1320 B.n743 B.n742 10.6151
R1321 B.n742 B.n53 10.6151
R1322 B.n736 B.n53 10.6151
R1323 B.n736 B.n735 10.6151
R1324 B.n735 B.n734 10.6151
R1325 B.n734 B.n59 10.6151
R1326 B.n728 B.n59 10.6151
R1327 B.n728 B.n727 10.6151
R1328 B.n727 B.n726 10.6151
R1329 B.n726 B.n67 10.6151
R1330 B.n720 B.n67 10.6151
R1331 B.n720 B.n719 10.6151
R1332 B.n719 B.n718 10.6151
R1333 B.n718 B.n74 10.6151
R1334 B.n712 B.n74 10.6151
R1335 B.n712 B.n711 10.6151
R1336 B.n711 B.n710 10.6151
R1337 B.n710 B.n81 10.6151
R1338 B.n705 B.n81 10.6151
R1339 B.n705 B.n704 10.6151
R1340 B.n704 B.n703 10.6151
R1341 B.n703 B.n88 10.6151
R1342 B.n697 B.n88 10.6151
R1343 B.n697 B.n696 10.6151
R1344 B.n696 B.n695 10.6151
R1345 B.n695 B.n95 10.6151
R1346 B.n689 B.n95 10.6151
R1347 B.n689 B.n688 10.6151
R1348 B.n687 B.n102 10.6151
R1349 B.n134 B.n102 10.6151
R1350 B.n135 B.n134 10.6151
R1351 B.n138 B.n135 10.6151
R1352 B.n139 B.n138 10.6151
R1353 B.n142 B.n139 10.6151
R1354 B.n143 B.n142 10.6151
R1355 B.n146 B.n143 10.6151
R1356 B.n147 B.n146 10.6151
R1357 B.n150 B.n147 10.6151
R1358 B.n151 B.n150 10.6151
R1359 B.n154 B.n151 10.6151
R1360 B.n155 B.n154 10.6151
R1361 B.n158 B.n155 10.6151
R1362 B.n159 B.n158 10.6151
R1363 B.n162 B.n159 10.6151
R1364 B.n163 B.n162 10.6151
R1365 B.n167 B.n166 10.6151
R1366 B.n170 B.n167 10.6151
R1367 B.n171 B.n170 10.6151
R1368 B.n174 B.n171 10.6151
R1369 B.n175 B.n174 10.6151
R1370 B.n178 B.n175 10.6151
R1371 B.n179 B.n178 10.6151
R1372 B.n182 B.n179 10.6151
R1373 B.n183 B.n182 10.6151
R1374 B.n187 B.n186 10.6151
R1375 B.n190 B.n187 10.6151
R1376 B.n191 B.n190 10.6151
R1377 B.n194 B.n191 10.6151
R1378 B.n195 B.n194 10.6151
R1379 B.n198 B.n195 10.6151
R1380 B.n199 B.n198 10.6151
R1381 B.n202 B.n199 10.6151
R1382 B.n203 B.n202 10.6151
R1383 B.n206 B.n203 10.6151
R1384 B.n207 B.n206 10.6151
R1385 B.n210 B.n207 10.6151
R1386 B.n211 B.n210 10.6151
R1387 B.n214 B.n211 10.6151
R1388 B.n216 B.n214 10.6151
R1389 B.n217 B.n216 10.6151
R1390 B.n681 B.n217 10.6151
R1391 B.n513 B.t0 9.46796
R1392 B.n61 B.t2 9.46796
R1393 B.n410 B.n409 9.36635
R1394 B.n388 B.n387 9.36635
R1395 B.n163 B.n132 9.36635
R1396 B.n186 B.n129 9.36635
R1397 B.n800 B.n0 8.11757
R1398 B.n800 B.n1 8.11757
R1399 B.t1 B.n228 4.73423
R1400 B.t19 B.n16 4.73423
R1401 B.n550 B.t3 2.36736
R1402 B.n40 B.t4 2.36736
R1403 B.n409 B.n408 1.24928
R1404 B.n389 B.n388 1.24928
R1405 B.n166 B.n132 1.24928
R1406 B.n183 B.n129 1.24928
R1407 VP.n16 VP.n13 161.3
R1408 VP.n18 VP.n17 161.3
R1409 VP.n19 VP.n12 161.3
R1410 VP.n21 VP.n20 161.3
R1411 VP.n22 VP.n11 161.3
R1412 VP.n24 VP.n23 161.3
R1413 VP.n25 VP.n10 161.3
R1414 VP.n27 VP.n26 161.3
R1415 VP.n56 VP.n55 161.3
R1416 VP.n54 VP.n1 161.3
R1417 VP.n53 VP.n52 161.3
R1418 VP.n51 VP.n2 161.3
R1419 VP.n50 VP.n49 161.3
R1420 VP.n48 VP.n3 161.3
R1421 VP.n47 VP.n46 161.3
R1422 VP.n45 VP.n4 161.3
R1423 VP.n44 VP.n43 161.3
R1424 VP.n42 VP.n5 161.3
R1425 VP.n41 VP.n40 161.3
R1426 VP.n39 VP.n6 161.3
R1427 VP.n38 VP.n37 161.3
R1428 VP.n36 VP.n7 161.3
R1429 VP.n35 VP.n34 161.3
R1430 VP.n33 VP.n8 161.3
R1431 VP.n32 VP.n31 161.3
R1432 VP.n30 VP.n29 87.7864
R1433 VP.n57 VP.n0 87.7864
R1434 VP.n28 VP.n9 87.7864
R1435 VP.n15 VP.t1 58.9142
R1436 VP.n15 VP.n14 50.5915
R1437 VP.n29 VP.n28 47.0488
R1438 VP.n37 VP.n36 42.999
R1439 VP.n49 VP.n2 42.999
R1440 VP.n20 VP.n11 42.999
R1441 VP.n37 VP.n6 38.1551
R1442 VP.n49 VP.n48 38.1551
R1443 VP.n20 VP.n19 38.1551
R1444 VP.n43 VP.t3 26.044
R1445 VP.n30 VP.t0 26.044
R1446 VP.n0 VP.t2 26.044
R1447 VP.n14 VP.t4 26.044
R1448 VP.n9 VP.t5 26.044
R1449 VP.n31 VP.n8 24.5923
R1450 VP.n35 VP.n8 24.5923
R1451 VP.n36 VP.n35 24.5923
R1452 VP.n41 VP.n6 24.5923
R1453 VP.n42 VP.n41 24.5923
R1454 VP.n43 VP.n42 24.5923
R1455 VP.n43 VP.n4 24.5923
R1456 VP.n47 VP.n4 24.5923
R1457 VP.n48 VP.n47 24.5923
R1458 VP.n53 VP.n2 24.5923
R1459 VP.n54 VP.n53 24.5923
R1460 VP.n55 VP.n54 24.5923
R1461 VP.n24 VP.n11 24.5923
R1462 VP.n25 VP.n24 24.5923
R1463 VP.n26 VP.n25 24.5923
R1464 VP.n14 VP.n13 24.5923
R1465 VP.n18 VP.n13 24.5923
R1466 VP.n19 VP.n18 24.5923
R1467 VP.n16 VP.n15 2.46239
R1468 VP.n31 VP.n30 2.45968
R1469 VP.n55 VP.n0 2.45968
R1470 VP.n26 VP.n9 2.45968
R1471 VP.n28 VP.n27 0.354861
R1472 VP.n32 VP.n29 0.354861
R1473 VP.n57 VP.n56 0.354861
R1474 VP VP.n57 0.267071
R1475 VP.n17 VP.n16 0.189894
R1476 VP.n17 VP.n12 0.189894
R1477 VP.n21 VP.n12 0.189894
R1478 VP.n22 VP.n21 0.189894
R1479 VP.n23 VP.n22 0.189894
R1480 VP.n23 VP.n10 0.189894
R1481 VP.n27 VP.n10 0.189894
R1482 VP.n33 VP.n32 0.189894
R1483 VP.n34 VP.n33 0.189894
R1484 VP.n34 VP.n7 0.189894
R1485 VP.n38 VP.n7 0.189894
R1486 VP.n39 VP.n38 0.189894
R1487 VP.n40 VP.n39 0.189894
R1488 VP.n40 VP.n5 0.189894
R1489 VP.n44 VP.n5 0.189894
R1490 VP.n45 VP.n44 0.189894
R1491 VP.n46 VP.n45 0.189894
R1492 VP.n46 VP.n3 0.189894
R1493 VP.n50 VP.n3 0.189894
R1494 VP.n51 VP.n50 0.189894
R1495 VP.n52 VP.n51 0.189894
R1496 VP.n52 VP.n1 0.189894
R1497 VP.n56 VP.n1 0.189894
R1498 VTAIL.n82 VTAIL.n68 289.615
R1499 VTAIL.n16 VTAIL.n2 289.615
R1500 VTAIL.n62 VTAIL.n48 289.615
R1501 VTAIL.n40 VTAIL.n26 289.615
R1502 VTAIL.n75 VTAIL.n74 185
R1503 VTAIL.n72 VTAIL.n71 185
R1504 VTAIL.n81 VTAIL.n80 185
R1505 VTAIL.n83 VTAIL.n82 185
R1506 VTAIL.n9 VTAIL.n8 185
R1507 VTAIL.n6 VTAIL.n5 185
R1508 VTAIL.n15 VTAIL.n14 185
R1509 VTAIL.n17 VTAIL.n16 185
R1510 VTAIL.n63 VTAIL.n62 185
R1511 VTAIL.n61 VTAIL.n60 185
R1512 VTAIL.n52 VTAIL.n51 185
R1513 VTAIL.n55 VTAIL.n54 185
R1514 VTAIL.n41 VTAIL.n40 185
R1515 VTAIL.n39 VTAIL.n38 185
R1516 VTAIL.n30 VTAIL.n29 185
R1517 VTAIL.n33 VTAIL.n32 185
R1518 VTAIL.t4 VTAIL.n73 147.888
R1519 VTAIL.t6 VTAIL.n7 147.888
R1520 VTAIL.t11 VTAIL.n53 147.888
R1521 VTAIL.t1 VTAIL.n31 147.888
R1522 VTAIL.n74 VTAIL.n71 104.615
R1523 VTAIL.n81 VTAIL.n71 104.615
R1524 VTAIL.n82 VTAIL.n81 104.615
R1525 VTAIL.n8 VTAIL.n5 104.615
R1526 VTAIL.n15 VTAIL.n5 104.615
R1527 VTAIL.n16 VTAIL.n15 104.615
R1528 VTAIL.n62 VTAIL.n61 104.615
R1529 VTAIL.n61 VTAIL.n51 104.615
R1530 VTAIL.n54 VTAIL.n51 104.615
R1531 VTAIL.n40 VTAIL.n39 104.615
R1532 VTAIL.n39 VTAIL.n29 104.615
R1533 VTAIL.n32 VTAIL.n29 104.615
R1534 VTAIL.n47 VTAIL.n46 60.2762
R1535 VTAIL.n25 VTAIL.n24 60.2762
R1536 VTAIL.n1 VTAIL.n0 60.2761
R1537 VTAIL.n23 VTAIL.n22 60.2761
R1538 VTAIL.n74 VTAIL.t4 52.3082
R1539 VTAIL.n8 VTAIL.t6 52.3082
R1540 VTAIL.n54 VTAIL.t11 52.3082
R1541 VTAIL.n32 VTAIL.t1 52.3082
R1542 VTAIL.n87 VTAIL.n86 35.6763
R1543 VTAIL.n21 VTAIL.n20 35.6763
R1544 VTAIL.n67 VTAIL.n66 35.6763
R1545 VTAIL.n45 VTAIL.n44 35.6763
R1546 VTAIL.n25 VTAIL.n23 22.8152
R1547 VTAIL.n87 VTAIL.n67 19.3238
R1548 VTAIL.n75 VTAIL.n73 15.6496
R1549 VTAIL.n9 VTAIL.n7 15.6496
R1550 VTAIL.n55 VTAIL.n53 15.6496
R1551 VTAIL.n33 VTAIL.n31 15.6496
R1552 VTAIL.n76 VTAIL.n72 12.8005
R1553 VTAIL.n10 VTAIL.n6 12.8005
R1554 VTAIL.n56 VTAIL.n52 12.8005
R1555 VTAIL.n34 VTAIL.n30 12.8005
R1556 VTAIL.n80 VTAIL.n79 12.0247
R1557 VTAIL.n14 VTAIL.n13 12.0247
R1558 VTAIL.n60 VTAIL.n59 12.0247
R1559 VTAIL.n38 VTAIL.n37 12.0247
R1560 VTAIL.n83 VTAIL.n70 11.249
R1561 VTAIL.n17 VTAIL.n4 11.249
R1562 VTAIL.n63 VTAIL.n50 11.249
R1563 VTAIL.n41 VTAIL.n28 11.249
R1564 VTAIL.n84 VTAIL.n68 10.4732
R1565 VTAIL.n18 VTAIL.n2 10.4732
R1566 VTAIL.n64 VTAIL.n48 10.4732
R1567 VTAIL.n42 VTAIL.n26 10.4732
R1568 VTAIL.n86 VTAIL.n85 9.45567
R1569 VTAIL.n20 VTAIL.n19 9.45567
R1570 VTAIL.n66 VTAIL.n65 9.45567
R1571 VTAIL.n44 VTAIL.n43 9.45567
R1572 VTAIL.n85 VTAIL.n84 9.3005
R1573 VTAIL.n70 VTAIL.n69 9.3005
R1574 VTAIL.n79 VTAIL.n78 9.3005
R1575 VTAIL.n77 VTAIL.n76 9.3005
R1576 VTAIL.n19 VTAIL.n18 9.3005
R1577 VTAIL.n4 VTAIL.n3 9.3005
R1578 VTAIL.n13 VTAIL.n12 9.3005
R1579 VTAIL.n11 VTAIL.n10 9.3005
R1580 VTAIL.n65 VTAIL.n64 9.3005
R1581 VTAIL.n50 VTAIL.n49 9.3005
R1582 VTAIL.n59 VTAIL.n58 9.3005
R1583 VTAIL.n57 VTAIL.n56 9.3005
R1584 VTAIL.n43 VTAIL.n42 9.3005
R1585 VTAIL.n28 VTAIL.n27 9.3005
R1586 VTAIL.n37 VTAIL.n36 9.3005
R1587 VTAIL.n35 VTAIL.n34 9.3005
R1588 VTAIL.n0 VTAIL.t3 4.92587
R1589 VTAIL.n0 VTAIL.t5 4.92587
R1590 VTAIL.n22 VTAIL.t8 4.92587
R1591 VTAIL.n22 VTAIL.t10 4.92587
R1592 VTAIL.n46 VTAIL.t7 4.92587
R1593 VTAIL.n46 VTAIL.t9 4.92587
R1594 VTAIL.n24 VTAIL.t2 4.92587
R1595 VTAIL.n24 VTAIL.t0 4.92587
R1596 VTAIL.n77 VTAIL.n73 4.40546
R1597 VTAIL.n11 VTAIL.n7 4.40546
R1598 VTAIL.n57 VTAIL.n53 4.40546
R1599 VTAIL.n35 VTAIL.n31 4.40546
R1600 VTAIL.n45 VTAIL.n25 3.49188
R1601 VTAIL.n67 VTAIL.n47 3.49188
R1602 VTAIL.n23 VTAIL.n21 3.49188
R1603 VTAIL.n86 VTAIL.n68 3.49141
R1604 VTAIL.n20 VTAIL.n2 3.49141
R1605 VTAIL.n66 VTAIL.n48 3.49141
R1606 VTAIL.n44 VTAIL.n26 3.49141
R1607 VTAIL.n84 VTAIL.n83 2.71565
R1608 VTAIL.n18 VTAIL.n17 2.71565
R1609 VTAIL.n64 VTAIL.n63 2.71565
R1610 VTAIL.n42 VTAIL.n41 2.71565
R1611 VTAIL VTAIL.n87 2.56084
R1612 VTAIL.n47 VTAIL.n45 2.21602
R1613 VTAIL.n21 VTAIL.n1 2.21602
R1614 VTAIL.n80 VTAIL.n70 1.93989
R1615 VTAIL.n14 VTAIL.n4 1.93989
R1616 VTAIL.n60 VTAIL.n50 1.93989
R1617 VTAIL.n38 VTAIL.n28 1.93989
R1618 VTAIL.n79 VTAIL.n72 1.16414
R1619 VTAIL.n13 VTAIL.n6 1.16414
R1620 VTAIL.n59 VTAIL.n52 1.16414
R1621 VTAIL.n37 VTAIL.n30 1.16414
R1622 VTAIL VTAIL.n1 0.931535
R1623 VTAIL.n76 VTAIL.n75 0.388379
R1624 VTAIL.n10 VTAIL.n9 0.388379
R1625 VTAIL.n56 VTAIL.n55 0.388379
R1626 VTAIL.n34 VTAIL.n33 0.388379
R1627 VTAIL.n78 VTAIL.n77 0.155672
R1628 VTAIL.n78 VTAIL.n69 0.155672
R1629 VTAIL.n85 VTAIL.n69 0.155672
R1630 VTAIL.n12 VTAIL.n11 0.155672
R1631 VTAIL.n12 VTAIL.n3 0.155672
R1632 VTAIL.n19 VTAIL.n3 0.155672
R1633 VTAIL.n65 VTAIL.n49 0.155672
R1634 VTAIL.n58 VTAIL.n49 0.155672
R1635 VTAIL.n58 VTAIL.n57 0.155672
R1636 VTAIL.n43 VTAIL.n27 0.155672
R1637 VTAIL.n36 VTAIL.n27 0.155672
R1638 VTAIL.n36 VTAIL.n35 0.155672
R1639 VDD1.n14 VDD1.n0 289.615
R1640 VDD1.n33 VDD1.n19 289.615
R1641 VDD1.n15 VDD1.n14 185
R1642 VDD1.n13 VDD1.n12 185
R1643 VDD1.n4 VDD1.n3 185
R1644 VDD1.n7 VDD1.n6 185
R1645 VDD1.n26 VDD1.n25 185
R1646 VDD1.n23 VDD1.n22 185
R1647 VDD1.n32 VDD1.n31 185
R1648 VDD1.n34 VDD1.n33 185
R1649 VDD1.t4 VDD1.n5 147.888
R1650 VDD1.t5 VDD1.n24 147.888
R1651 VDD1.n14 VDD1.n13 104.615
R1652 VDD1.n13 VDD1.n3 104.615
R1653 VDD1.n6 VDD1.n3 104.615
R1654 VDD1.n25 VDD1.n22 104.615
R1655 VDD1.n32 VDD1.n22 104.615
R1656 VDD1.n33 VDD1.n32 104.615
R1657 VDD1.n39 VDD1.n38 77.7724
R1658 VDD1.n41 VDD1.n40 76.9549
R1659 VDD1 VDD1.n18 55.0318
R1660 VDD1.n39 VDD1.n37 54.9182
R1661 VDD1.n6 VDD1.t4 52.3082
R1662 VDD1.n25 VDD1.t5 52.3082
R1663 VDD1.n41 VDD1.n39 40.8565
R1664 VDD1.n7 VDD1.n5 15.6496
R1665 VDD1.n26 VDD1.n24 15.6496
R1666 VDD1.n8 VDD1.n4 12.8005
R1667 VDD1.n27 VDD1.n23 12.8005
R1668 VDD1.n12 VDD1.n11 12.0247
R1669 VDD1.n31 VDD1.n30 12.0247
R1670 VDD1.n15 VDD1.n2 11.249
R1671 VDD1.n34 VDD1.n21 11.249
R1672 VDD1.n16 VDD1.n0 10.4732
R1673 VDD1.n35 VDD1.n19 10.4732
R1674 VDD1.n18 VDD1.n17 9.45567
R1675 VDD1.n37 VDD1.n36 9.45567
R1676 VDD1.n17 VDD1.n16 9.3005
R1677 VDD1.n2 VDD1.n1 9.3005
R1678 VDD1.n11 VDD1.n10 9.3005
R1679 VDD1.n9 VDD1.n8 9.3005
R1680 VDD1.n36 VDD1.n35 9.3005
R1681 VDD1.n21 VDD1.n20 9.3005
R1682 VDD1.n30 VDD1.n29 9.3005
R1683 VDD1.n28 VDD1.n27 9.3005
R1684 VDD1.n40 VDD1.t1 4.92587
R1685 VDD1.n40 VDD1.t0 4.92587
R1686 VDD1.n38 VDD1.t2 4.92587
R1687 VDD1.n38 VDD1.t3 4.92587
R1688 VDD1.n9 VDD1.n5 4.40546
R1689 VDD1.n28 VDD1.n24 4.40546
R1690 VDD1.n18 VDD1.n0 3.49141
R1691 VDD1.n37 VDD1.n19 3.49141
R1692 VDD1.n16 VDD1.n15 2.71565
R1693 VDD1.n35 VDD1.n34 2.71565
R1694 VDD1.n12 VDD1.n2 1.93989
R1695 VDD1.n31 VDD1.n21 1.93989
R1696 VDD1.n11 VDD1.n4 1.16414
R1697 VDD1.n30 VDD1.n23 1.16414
R1698 VDD1 VDD1.n41 0.815155
R1699 VDD1.n8 VDD1.n7 0.388379
R1700 VDD1.n27 VDD1.n26 0.388379
R1701 VDD1.n17 VDD1.n1 0.155672
R1702 VDD1.n10 VDD1.n1 0.155672
R1703 VDD1.n10 VDD1.n9 0.155672
R1704 VDD1.n29 VDD1.n28 0.155672
R1705 VDD1.n29 VDD1.n20 0.155672
R1706 VDD1.n36 VDD1.n20 0.155672
R1707 VN.n38 VN.n37 161.3
R1708 VN.n36 VN.n21 161.3
R1709 VN.n35 VN.n34 161.3
R1710 VN.n33 VN.n22 161.3
R1711 VN.n32 VN.n31 161.3
R1712 VN.n30 VN.n23 161.3
R1713 VN.n29 VN.n28 161.3
R1714 VN.n27 VN.n24 161.3
R1715 VN.n18 VN.n17 161.3
R1716 VN.n16 VN.n1 161.3
R1717 VN.n15 VN.n14 161.3
R1718 VN.n13 VN.n2 161.3
R1719 VN.n12 VN.n11 161.3
R1720 VN.n10 VN.n3 161.3
R1721 VN.n9 VN.n8 161.3
R1722 VN.n7 VN.n4 161.3
R1723 VN.n19 VN.n0 87.7864
R1724 VN.n39 VN.n20 87.7864
R1725 VN.n26 VN.t1 58.9143
R1726 VN.n6 VN.t2 58.9143
R1727 VN.n6 VN.n5 50.5915
R1728 VN.n26 VN.n25 50.5915
R1729 VN VN.n39 47.214
R1730 VN.n11 VN.n2 42.999
R1731 VN.n31 VN.n22 42.999
R1732 VN.n11 VN.n10 38.1551
R1733 VN.n31 VN.n30 38.1551
R1734 VN.n5 VN.t3 26.044
R1735 VN.n0 VN.t4 26.044
R1736 VN.n25 VN.t5 26.044
R1737 VN.n20 VN.t0 26.044
R1738 VN.n5 VN.n4 24.5923
R1739 VN.n9 VN.n4 24.5923
R1740 VN.n10 VN.n9 24.5923
R1741 VN.n15 VN.n2 24.5923
R1742 VN.n16 VN.n15 24.5923
R1743 VN.n17 VN.n16 24.5923
R1744 VN.n30 VN.n29 24.5923
R1745 VN.n29 VN.n24 24.5923
R1746 VN.n25 VN.n24 24.5923
R1747 VN.n37 VN.n36 24.5923
R1748 VN.n36 VN.n35 24.5923
R1749 VN.n35 VN.n22 24.5923
R1750 VN.n27 VN.n26 2.4624
R1751 VN.n7 VN.n6 2.4624
R1752 VN.n17 VN.n0 2.45968
R1753 VN.n37 VN.n20 2.45968
R1754 VN.n39 VN.n38 0.354861
R1755 VN.n19 VN.n18 0.354861
R1756 VN VN.n19 0.267071
R1757 VN.n38 VN.n21 0.189894
R1758 VN.n34 VN.n21 0.189894
R1759 VN.n34 VN.n33 0.189894
R1760 VN.n33 VN.n32 0.189894
R1761 VN.n32 VN.n23 0.189894
R1762 VN.n28 VN.n23 0.189894
R1763 VN.n28 VN.n27 0.189894
R1764 VN.n8 VN.n7 0.189894
R1765 VN.n8 VN.n3 0.189894
R1766 VN.n12 VN.n3 0.189894
R1767 VN.n13 VN.n12 0.189894
R1768 VN.n14 VN.n13 0.189894
R1769 VN.n14 VN.n1 0.189894
R1770 VN.n18 VN.n1 0.189894
R1771 VDD2.n35 VDD2.n21 289.615
R1772 VDD2.n14 VDD2.n0 289.615
R1773 VDD2.n36 VDD2.n35 185
R1774 VDD2.n34 VDD2.n33 185
R1775 VDD2.n25 VDD2.n24 185
R1776 VDD2.n28 VDD2.n27 185
R1777 VDD2.n7 VDD2.n6 185
R1778 VDD2.n4 VDD2.n3 185
R1779 VDD2.n13 VDD2.n12 185
R1780 VDD2.n15 VDD2.n14 185
R1781 VDD2.t5 VDD2.n26 147.888
R1782 VDD2.t3 VDD2.n5 147.888
R1783 VDD2.n35 VDD2.n34 104.615
R1784 VDD2.n34 VDD2.n24 104.615
R1785 VDD2.n27 VDD2.n24 104.615
R1786 VDD2.n6 VDD2.n3 104.615
R1787 VDD2.n13 VDD2.n3 104.615
R1788 VDD2.n14 VDD2.n13 104.615
R1789 VDD2.n20 VDD2.n19 77.7724
R1790 VDD2 VDD2.n41 77.7695
R1791 VDD2.n20 VDD2.n18 54.9182
R1792 VDD2.n40 VDD2.n39 52.355
R1793 VDD2.n27 VDD2.t5 52.3082
R1794 VDD2.n6 VDD2.t3 52.3082
R1795 VDD2.n40 VDD2.n20 38.5278
R1796 VDD2.n28 VDD2.n26 15.6496
R1797 VDD2.n7 VDD2.n5 15.6496
R1798 VDD2.n29 VDD2.n25 12.8005
R1799 VDD2.n8 VDD2.n4 12.8005
R1800 VDD2.n33 VDD2.n32 12.0247
R1801 VDD2.n12 VDD2.n11 12.0247
R1802 VDD2.n36 VDD2.n23 11.249
R1803 VDD2.n15 VDD2.n2 11.249
R1804 VDD2.n37 VDD2.n21 10.4732
R1805 VDD2.n16 VDD2.n0 10.4732
R1806 VDD2.n39 VDD2.n38 9.45567
R1807 VDD2.n18 VDD2.n17 9.45567
R1808 VDD2.n38 VDD2.n37 9.3005
R1809 VDD2.n23 VDD2.n22 9.3005
R1810 VDD2.n32 VDD2.n31 9.3005
R1811 VDD2.n30 VDD2.n29 9.3005
R1812 VDD2.n17 VDD2.n16 9.3005
R1813 VDD2.n2 VDD2.n1 9.3005
R1814 VDD2.n11 VDD2.n10 9.3005
R1815 VDD2.n9 VDD2.n8 9.3005
R1816 VDD2.n41 VDD2.t0 4.92587
R1817 VDD2.n41 VDD2.t4 4.92587
R1818 VDD2.n19 VDD2.t2 4.92587
R1819 VDD2.n19 VDD2.t1 4.92587
R1820 VDD2.n30 VDD2.n26 4.40546
R1821 VDD2.n9 VDD2.n5 4.40546
R1822 VDD2.n39 VDD2.n21 3.49141
R1823 VDD2.n18 VDD2.n0 3.49141
R1824 VDD2.n37 VDD2.n36 2.71565
R1825 VDD2.n16 VDD2.n15 2.71565
R1826 VDD2 VDD2.n40 2.67722
R1827 VDD2.n33 VDD2.n23 1.93989
R1828 VDD2.n12 VDD2.n2 1.93989
R1829 VDD2.n32 VDD2.n25 1.16414
R1830 VDD2.n11 VDD2.n4 1.16414
R1831 VDD2.n29 VDD2.n28 0.388379
R1832 VDD2.n8 VDD2.n7 0.388379
R1833 VDD2.n38 VDD2.n22 0.155672
R1834 VDD2.n31 VDD2.n22 0.155672
R1835 VDD2.n31 VDD2.n30 0.155672
R1836 VDD2.n10 VDD2.n9 0.155672
R1837 VDD2.n10 VDD2.n1 0.155672
R1838 VDD2.n17 VDD2.n1 0.155672
C0 VDD1 VTAIL 5.56677f
C1 VDD2 VP 0.557776f
C2 VDD2 VN 2.66301f
C3 VN VP 6.53928f
C4 VDD1 VDD2 1.84228f
C5 VDD1 VP 3.06141f
C6 VDD1 VN 0.156716f
C7 VDD2 VTAIL 5.62729f
C8 VTAIL VP 3.72234f
C9 VTAIL VN 3.70808f
C10 VDD2 B 5.42277f
C11 VDD1 B 5.616266f
C12 VTAIL B 4.81954f
C13 VN B 15.47746f
C14 VP B 14.106197f
C15 VDD2.n0 B 0.032182f
C16 VDD2.n1 B 0.022254f
C17 VDD2.n2 B 0.011959f
C18 VDD2.n3 B 0.028266f
C19 VDD2.n4 B 0.012662f
C20 VDD2.n5 B 0.086314f
C21 VDD2.t3 B 0.047107f
C22 VDD2.n6 B 0.021199f
C23 VDD2.n7 B 0.016636f
C24 VDD2.n8 B 0.011959f
C25 VDD2.n9 B 0.324322f
C26 VDD2.n10 B 0.022254f
C27 VDD2.n11 B 0.011959f
C28 VDD2.n12 B 0.012662f
C29 VDD2.n13 B 0.028266f
C30 VDD2.n14 B 0.062784f
C31 VDD2.n15 B 0.012662f
C32 VDD2.n16 B 0.011959f
C33 VDD2.n17 B 0.056913f
C34 VDD2.n18 B 0.061517f
C35 VDD2.t2 B 0.070696f
C36 VDD2.t1 B 0.070696f
C37 VDD2.n19 B 0.560589f
C38 VDD2.n20 B 2.37741f
C39 VDD2.n21 B 0.032182f
C40 VDD2.n22 B 0.022254f
C41 VDD2.n23 B 0.011959f
C42 VDD2.n24 B 0.028266f
C43 VDD2.n25 B 0.012662f
C44 VDD2.n26 B 0.086314f
C45 VDD2.t5 B 0.047107f
C46 VDD2.n27 B 0.021199f
C47 VDD2.n28 B 0.016636f
C48 VDD2.n29 B 0.011959f
C49 VDD2.n30 B 0.324322f
C50 VDD2.n31 B 0.022254f
C51 VDD2.n32 B 0.011959f
C52 VDD2.n33 B 0.012662f
C53 VDD2.n34 B 0.028266f
C54 VDD2.n35 B 0.062784f
C55 VDD2.n36 B 0.012662f
C56 VDD2.n37 B 0.011959f
C57 VDD2.n38 B 0.056913f
C58 VDD2.n39 B 0.050782f
C59 VDD2.n40 B 2.00086f
C60 VDD2.t0 B 0.070696f
C61 VDD2.t4 B 0.070696f
C62 VDD2.n41 B 0.560563f
C63 VN.t4 B 0.912898f
C64 VN.n0 B 0.439784f
C65 VN.n1 B 0.023752f
C66 VN.n2 B 0.04628f
C67 VN.n3 B 0.023752f
C68 VN.n4 B 0.044046f
C69 VN.t3 B 0.912898f
C70 VN.n5 B 0.450241f
C71 VN.t2 B 1.21399f
C72 VN.n6 B 0.446316f
C73 VN.n7 B 0.302873f
C74 VN.n8 B 0.023752f
C75 VN.n9 B 0.044046f
C76 VN.n10 B 0.047447f
C77 VN.n11 B 0.019374f
C78 VN.n12 B 0.023752f
C79 VN.n13 B 0.023752f
C80 VN.n14 B 0.023752f
C81 VN.n15 B 0.044046f
C82 VN.n16 B 0.044046f
C83 VN.n17 B 0.024476f
C84 VN.n18 B 0.03833f
C85 VN.n19 B 0.072103f
C86 VN.t0 B 0.912898f
C87 VN.n20 B 0.439784f
C88 VN.n21 B 0.023752f
C89 VN.n22 B 0.04628f
C90 VN.n23 B 0.023752f
C91 VN.n24 B 0.044046f
C92 VN.t1 B 1.21399f
C93 VN.t5 B 0.912898f
C94 VN.n25 B 0.450241f
C95 VN.n26 B 0.446316f
C96 VN.n27 B 0.302873f
C97 VN.n28 B 0.023752f
C98 VN.n29 B 0.044046f
C99 VN.n30 B 0.047447f
C100 VN.n31 B 0.019374f
C101 VN.n32 B 0.023752f
C102 VN.n33 B 0.023752f
C103 VN.n34 B 0.023752f
C104 VN.n35 B 0.044046f
C105 VN.n36 B 0.044046f
C106 VN.n37 B 0.024476f
C107 VN.n38 B 0.03833f
C108 VN.n39 B 1.26053f
C109 VDD1.n0 B 0.033402f
C110 VDD1.n1 B 0.023098f
C111 VDD1.n2 B 0.012412f
C112 VDD1.n3 B 0.029337f
C113 VDD1.n4 B 0.013142f
C114 VDD1.n5 B 0.089587f
C115 VDD1.t4 B 0.048893f
C116 VDD1.n6 B 0.022003f
C117 VDD1.n7 B 0.017267f
C118 VDD1.n8 B 0.012412f
C119 VDD1.n9 B 0.336618f
C120 VDD1.n10 B 0.023098f
C121 VDD1.n11 B 0.012412f
C122 VDD1.n12 B 0.013142f
C123 VDD1.n13 B 0.029337f
C124 VDD1.n14 B 0.065164f
C125 VDD1.n15 B 0.013142f
C126 VDD1.n16 B 0.012412f
C127 VDD1.n17 B 0.05907f
C128 VDD1.n18 B 0.064719f
C129 VDD1.n19 B 0.033402f
C130 VDD1.n20 B 0.023098f
C131 VDD1.n21 B 0.012412f
C132 VDD1.n22 B 0.029337f
C133 VDD1.n23 B 0.013142f
C134 VDD1.n24 B 0.089587f
C135 VDD1.t5 B 0.048893f
C136 VDD1.n25 B 0.022003f
C137 VDD1.n26 B 0.017267f
C138 VDD1.n27 B 0.012412f
C139 VDD1.n28 B 0.336618f
C140 VDD1.n29 B 0.023098f
C141 VDD1.n30 B 0.012412f
C142 VDD1.n31 B 0.013142f
C143 VDD1.n32 B 0.029337f
C144 VDD1.n33 B 0.065164f
C145 VDD1.n34 B 0.013142f
C146 VDD1.n35 B 0.012412f
C147 VDD1.n36 B 0.05907f
C148 VDD1.n37 B 0.063849f
C149 VDD1.t2 B 0.073377f
C150 VDD1.t3 B 0.073377f
C151 VDD1.n38 B 0.581843f
C152 VDD1.n39 B 2.60121f
C153 VDD1.t1 B 0.073377f
C154 VDD1.t0 B 0.073377f
C155 VDD1.n40 B 0.57647f
C156 VDD1.n41 B 2.2917f
C157 VTAIL.t3 B 0.099069f
C158 VTAIL.t5 B 0.099069f
C159 VTAIL.n0 B 0.712525f
C160 VTAIL.n1 B 0.583284f
C161 VTAIL.n2 B 0.045097f
C162 VTAIL.n3 B 0.031186f
C163 VTAIL.n4 B 0.016758f
C164 VTAIL.n5 B 0.03961f
C165 VTAIL.n6 B 0.017744f
C166 VTAIL.n7 B 0.120954f
C167 VTAIL.t6 B 0.066012f
C168 VTAIL.n8 B 0.029707f
C169 VTAIL.n9 B 0.023313f
C170 VTAIL.n10 B 0.016758f
C171 VTAIL.n11 B 0.45448f
C172 VTAIL.n12 B 0.031186f
C173 VTAIL.n13 B 0.016758f
C174 VTAIL.n14 B 0.017744f
C175 VTAIL.n15 B 0.03961f
C176 VTAIL.n16 B 0.087981f
C177 VTAIL.n17 B 0.017744f
C178 VTAIL.n18 B 0.016758f
C179 VTAIL.n19 B 0.079753f
C180 VTAIL.n20 B 0.049683f
C181 VTAIL.n21 B 0.604446f
C182 VTAIL.t8 B 0.099069f
C183 VTAIL.t10 B 0.099069f
C184 VTAIL.n22 B 0.712525f
C185 VTAIL.n23 B 2.09148f
C186 VTAIL.t2 B 0.099069f
C187 VTAIL.t0 B 0.099069f
C188 VTAIL.n24 B 0.71253f
C189 VTAIL.n25 B 2.09147f
C190 VTAIL.n26 B 0.045097f
C191 VTAIL.n27 B 0.031186f
C192 VTAIL.n28 B 0.016758f
C193 VTAIL.n29 B 0.03961f
C194 VTAIL.n30 B 0.017744f
C195 VTAIL.n31 B 0.120954f
C196 VTAIL.t1 B 0.066012f
C197 VTAIL.n32 B 0.029707f
C198 VTAIL.n33 B 0.023313f
C199 VTAIL.n34 B 0.016758f
C200 VTAIL.n35 B 0.45448f
C201 VTAIL.n36 B 0.031186f
C202 VTAIL.n37 B 0.016758f
C203 VTAIL.n38 B 0.017744f
C204 VTAIL.n39 B 0.03961f
C205 VTAIL.n40 B 0.087981f
C206 VTAIL.n41 B 0.017744f
C207 VTAIL.n42 B 0.016758f
C208 VTAIL.n43 B 0.079753f
C209 VTAIL.n44 B 0.049683f
C210 VTAIL.n45 B 0.604446f
C211 VTAIL.t7 B 0.099069f
C212 VTAIL.t9 B 0.099069f
C213 VTAIL.n46 B 0.71253f
C214 VTAIL.n47 B 0.840562f
C215 VTAIL.n48 B 0.045097f
C216 VTAIL.n49 B 0.031186f
C217 VTAIL.n50 B 0.016758f
C218 VTAIL.n51 B 0.03961f
C219 VTAIL.n52 B 0.017744f
C220 VTAIL.n53 B 0.120954f
C221 VTAIL.t11 B 0.066012f
C222 VTAIL.n54 B 0.029707f
C223 VTAIL.n55 B 0.023313f
C224 VTAIL.n56 B 0.016758f
C225 VTAIL.n57 B 0.45448f
C226 VTAIL.n58 B 0.031186f
C227 VTAIL.n59 B 0.016758f
C228 VTAIL.n60 B 0.017744f
C229 VTAIL.n61 B 0.03961f
C230 VTAIL.n62 B 0.087981f
C231 VTAIL.n63 B 0.017744f
C232 VTAIL.n64 B 0.016758f
C233 VTAIL.n65 B 0.079753f
C234 VTAIL.n66 B 0.049683f
C235 VTAIL.n67 B 1.50452f
C236 VTAIL.n68 B 0.045097f
C237 VTAIL.n69 B 0.031186f
C238 VTAIL.n70 B 0.016758f
C239 VTAIL.n71 B 0.03961f
C240 VTAIL.n72 B 0.017744f
C241 VTAIL.n73 B 0.120954f
C242 VTAIL.t4 B 0.066012f
C243 VTAIL.n74 B 0.029707f
C244 VTAIL.n75 B 0.023313f
C245 VTAIL.n76 B 0.016758f
C246 VTAIL.n77 B 0.45448f
C247 VTAIL.n78 B 0.031186f
C248 VTAIL.n79 B 0.016758f
C249 VTAIL.n80 B 0.017744f
C250 VTAIL.n81 B 0.03961f
C251 VTAIL.n82 B 0.087981f
C252 VTAIL.n83 B 0.017744f
C253 VTAIL.n84 B 0.016758f
C254 VTAIL.n85 B 0.079753f
C255 VTAIL.n86 B 0.049683f
C256 VTAIL.n87 B 1.41096f
C257 VP.t2 B 0.943647f
C258 VP.n0 B 0.454597f
C259 VP.n1 B 0.024552f
C260 VP.n2 B 0.047839f
C261 VP.n3 B 0.024552f
C262 VP.n4 B 0.04553f
C263 VP.n5 B 0.024552f
C264 VP.t3 B 0.943647f
C265 VP.n6 B 0.049045f
C266 VP.n7 B 0.024552f
C267 VP.n8 B 0.04553f
C268 VP.t5 B 0.943647f
C269 VP.n9 B 0.454597f
C270 VP.n10 B 0.024552f
C271 VP.n11 B 0.047839f
C272 VP.n12 B 0.024552f
C273 VP.n13 B 0.04553f
C274 VP.t1 B 1.25488f
C275 VP.t4 B 0.943647f
C276 VP.n14 B 0.465407f
C277 VP.n15 B 0.46135f
C278 VP.n16 B 0.313075f
C279 VP.n17 B 0.024552f
C280 VP.n18 B 0.04553f
C281 VP.n19 B 0.049045f
C282 VP.n20 B 0.020026f
C283 VP.n21 B 0.024552f
C284 VP.n22 B 0.024552f
C285 VP.n23 B 0.024552f
C286 VP.n24 B 0.04553f
C287 VP.n25 B 0.04553f
C288 VP.n26 B 0.025301f
C289 VP.n27 B 0.039621f
C290 VP.n28 B 1.29272f
C291 VP.n29 B 1.31154f
C292 VP.t0 B 0.943647f
C293 VP.n30 B 0.454597f
C294 VP.n31 B 0.025301f
C295 VP.n32 B 0.039621f
C296 VP.n33 B 0.024552f
C297 VP.n34 B 0.024552f
C298 VP.n35 B 0.04553f
C299 VP.n36 B 0.047839f
C300 VP.n37 B 0.020026f
C301 VP.n38 B 0.024552f
C302 VP.n39 B 0.024552f
C303 VP.n40 B 0.024552f
C304 VP.n41 B 0.04553f
C305 VP.n42 B 0.04553f
C306 VP.n43 B 0.388519f
C307 VP.n44 B 0.024552f
C308 VP.n45 B 0.024552f
C309 VP.n46 B 0.024552f
C310 VP.n47 B 0.04553f
C311 VP.n48 B 0.049045f
C312 VP.n49 B 0.020026f
C313 VP.n50 B 0.024552f
C314 VP.n51 B 0.024552f
C315 VP.n52 B 0.024552f
C316 VP.n53 B 0.04553f
C317 VP.n54 B 0.04553f
C318 VP.n55 B 0.025301f
C319 VP.n56 B 0.039621f
C320 VP.n57 B 0.074532f
.ends

