* NGSPICE file created from diff_pair_sample_0980.ext - technology: sky130A

.subckt diff_pair_sample_0980 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=5.7759 ps=30.4 w=14.81 l=0.6
X1 B.t11 B.t9 B.t10 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=0 ps=0 w=14.81 l=0.6
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=5.7759 ps=30.4 w=14.81 l=0.6
X3 B.t8 B.t6 B.t7 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=0 ps=0 w=14.81 l=0.6
X4 B.t5 B.t3 B.t4 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=0 ps=0 w=14.81 l=0.6
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=5.7759 ps=30.4 w=14.81 l=0.6
X6 B.t2 B.t0 B.t1 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=0 ps=0 w=14.81 l=0.6
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1342_n3934# sky130_fd_pr__pfet_01v8 ad=5.7759 pd=30.4 as=5.7759 ps=30.4 w=14.81 l=0.6
R0 VN VN.t1 863.919
R1 VN VN.t0 822.093
R2 VTAIL.n322 VTAIL.n246 756.745
R3 VTAIL.n76 VTAIL.n0 756.745
R4 VTAIL.n240 VTAIL.n164 756.745
R5 VTAIL.n158 VTAIL.n82 756.745
R6 VTAIL.n273 VTAIL.n272 585
R7 VTAIL.n270 VTAIL.n269 585
R8 VTAIL.n279 VTAIL.n278 585
R9 VTAIL.n281 VTAIL.n280 585
R10 VTAIL.n266 VTAIL.n265 585
R11 VTAIL.n287 VTAIL.n286 585
R12 VTAIL.n289 VTAIL.n288 585
R13 VTAIL.n262 VTAIL.n261 585
R14 VTAIL.n295 VTAIL.n294 585
R15 VTAIL.n297 VTAIL.n296 585
R16 VTAIL.n258 VTAIL.n257 585
R17 VTAIL.n303 VTAIL.n302 585
R18 VTAIL.n305 VTAIL.n304 585
R19 VTAIL.n254 VTAIL.n253 585
R20 VTAIL.n311 VTAIL.n310 585
R21 VTAIL.n314 VTAIL.n313 585
R22 VTAIL.n312 VTAIL.n250 585
R23 VTAIL.n319 VTAIL.n249 585
R24 VTAIL.n321 VTAIL.n320 585
R25 VTAIL.n323 VTAIL.n322 585
R26 VTAIL.n27 VTAIL.n26 585
R27 VTAIL.n24 VTAIL.n23 585
R28 VTAIL.n33 VTAIL.n32 585
R29 VTAIL.n35 VTAIL.n34 585
R30 VTAIL.n20 VTAIL.n19 585
R31 VTAIL.n41 VTAIL.n40 585
R32 VTAIL.n43 VTAIL.n42 585
R33 VTAIL.n16 VTAIL.n15 585
R34 VTAIL.n49 VTAIL.n48 585
R35 VTAIL.n51 VTAIL.n50 585
R36 VTAIL.n12 VTAIL.n11 585
R37 VTAIL.n57 VTAIL.n56 585
R38 VTAIL.n59 VTAIL.n58 585
R39 VTAIL.n8 VTAIL.n7 585
R40 VTAIL.n65 VTAIL.n64 585
R41 VTAIL.n68 VTAIL.n67 585
R42 VTAIL.n66 VTAIL.n4 585
R43 VTAIL.n73 VTAIL.n3 585
R44 VTAIL.n75 VTAIL.n74 585
R45 VTAIL.n77 VTAIL.n76 585
R46 VTAIL.n241 VTAIL.n240 585
R47 VTAIL.n239 VTAIL.n238 585
R48 VTAIL.n237 VTAIL.n167 585
R49 VTAIL.n171 VTAIL.n168 585
R50 VTAIL.n232 VTAIL.n231 585
R51 VTAIL.n230 VTAIL.n229 585
R52 VTAIL.n173 VTAIL.n172 585
R53 VTAIL.n224 VTAIL.n223 585
R54 VTAIL.n222 VTAIL.n221 585
R55 VTAIL.n177 VTAIL.n176 585
R56 VTAIL.n216 VTAIL.n215 585
R57 VTAIL.n214 VTAIL.n213 585
R58 VTAIL.n181 VTAIL.n180 585
R59 VTAIL.n208 VTAIL.n207 585
R60 VTAIL.n206 VTAIL.n205 585
R61 VTAIL.n185 VTAIL.n184 585
R62 VTAIL.n200 VTAIL.n199 585
R63 VTAIL.n198 VTAIL.n197 585
R64 VTAIL.n189 VTAIL.n188 585
R65 VTAIL.n192 VTAIL.n191 585
R66 VTAIL.n159 VTAIL.n158 585
R67 VTAIL.n157 VTAIL.n156 585
R68 VTAIL.n155 VTAIL.n85 585
R69 VTAIL.n89 VTAIL.n86 585
R70 VTAIL.n150 VTAIL.n149 585
R71 VTAIL.n148 VTAIL.n147 585
R72 VTAIL.n91 VTAIL.n90 585
R73 VTAIL.n142 VTAIL.n141 585
R74 VTAIL.n140 VTAIL.n139 585
R75 VTAIL.n95 VTAIL.n94 585
R76 VTAIL.n134 VTAIL.n133 585
R77 VTAIL.n132 VTAIL.n131 585
R78 VTAIL.n99 VTAIL.n98 585
R79 VTAIL.n126 VTAIL.n125 585
R80 VTAIL.n124 VTAIL.n123 585
R81 VTAIL.n103 VTAIL.n102 585
R82 VTAIL.n118 VTAIL.n117 585
R83 VTAIL.n116 VTAIL.n115 585
R84 VTAIL.n107 VTAIL.n106 585
R85 VTAIL.n110 VTAIL.n109 585
R86 VTAIL.t0 VTAIL.n190 327.466
R87 VTAIL.t3 VTAIL.n108 327.466
R88 VTAIL.t2 VTAIL.n271 327.466
R89 VTAIL.t1 VTAIL.n25 327.466
R90 VTAIL.n272 VTAIL.n269 171.744
R91 VTAIL.n279 VTAIL.n269 171.744
R92 VTAIL.n280 VTAIL.n279 171.744
R93 VTAIL.n280 VTAIL.n265 171.744
R94 VTAIL.n287 VTAIL.n265 171.744
R95 VTAIL.n288 VTAIL.n287 171.744
R96 VTAIL.n288 VTAIL.n261 171.744
R97 VTAIL.n295 VTAIL.n261 171.744
R98 VTAIL.n296 VTAIL.n295 171.744
R99 VTAIL.n296 VTAIL.n257 171.744
R100 VTAIL.n303 VTAIL.n257 171.744
R101 VTAIL.n304 VTAIL.n303 171.744
R102 VTAIL.n304 VTAIL.n253 171.744
R103 VTAIL.n311 VTAIL.n253 171.744
R104 VTAIL.n313 VTAIL.n311 171.744
R105 VTAIL.n313 VTAIL.n312 171.744
R106 VTAIL.n312 VTAIL.n249 171.744
R107 VTAIL.n321 VTAIL.n249 171.744
R108 VTAIL.n322 VTAIL.n321 171.744
R109 VTAIL.n26 VTAIL.n23 171.744
R110 VTAIL.n33 VTAIL.n23 171.744
R111 VTAIL.n34 VTAIL.n33 171.744
R112 VTAIL.n34 VTAIL.n19 171.744
R113 VTAIL.n41 VTAIL.n19 171.744
R114 VTAIL.n42 VTAIL.n41 171.744
R115 VTAIL.n42 VTAIL.n15 171.744
R116 VTAIL.n49 VTAIL.n15 171.744
R117 VTAIL.n50 VTAIL.n49 171.744
R118 VTAIL.n50 VTAIL.n11 171.744
R119 VTAIL.n57 VTAIL.n11 171.744
R120 VTAIL.n58 VTAIL.n57 171.744
R121 VTAIL.n58 VTAIL.n7 171.744
R122 VTAIL.n65 VTAIL.n7 171.744
R123 VTAIL.n67 VTAIL.n65 171.744
R124 VTAIL.n67 VTAIL.n66 171.744
R125 VTAIL.n66 VTAIL.n3 171.744
R126 VTAIL.n75 VTAIL.n3 171.744
R127 VTAIL.n76 VTAIL.n75 171.744
R128 VTAIL.n240 VTAIL.n239 171.744
R129 VTAIL.n239 VTAIL.n167 171.744
R130 VTAIL.n171 VTAIL.n167 171.744
R131 VTAIL.n231 VTAIL.n171 171.744
R132 VTAIL.n231 VTAIL.n230 171.744
R133 VTAIL.n230 VTAIL.n172 171.744
R134 VTAIL.n223 VTAIL.n172 171.744
R135 VTAIL.n223 VTAIL.n222 171.744
R136 VTAIL.n222 VTAIL.n176 171.744
R137 VTAIL.n215 VTAIL.n176 171.744
R138 VTAIL.n215 VTAIL.n214 171.744
R139 VTAIL.n214 VTAIL.n180 171.744
R140 VTAIL.n207 VTAIL.n180 171.744
R141 VTAIL.n207 VTAIL.n206 171.744
R142 VTAIL.n206 VTAIL.n184 171.744
R143 VTAIL.n199 VTAIL.n184 171.744
R144 VTAIL.n199 VTAIL.n198 171.744
R145 VTAIL.n198 VTAIL.n188 171.744
R146 VTAIL.n191 VTAIL.n188 171.744
R147 VTAIL.n158 VTAIL.n157 171.744
R148 VTAIL.n157 VTAIL.n85 171.744
R149 VTAIL.n89 VTAIL.n85 171.744
R150 VTAIL.n149 VTAIL.n89 171.744
R151 VTAIL.n149 VTAIL.n148 171.744
R152 VTAIL.n148 VTAIL.n90 171.744
R153 VTAIL.n141 VTAIL.n90 171.744
R154 VTAIL.n141 VTAIL.n140 171.744
R155 VTAIL.n140 VTAIL.n94 171.744
R156 VTAIL.n133 VTAIL.n94 171.744
R157 VTAIL.n133 VTAIL.n132 171.744
R158 VTAIL.n132 VTAIL.n98 171.744
R159 VTAIL.n125 VTAIL.n98 171.744
R160 VTAIL.n125 VTAIL.n124 171.744
R161 VTAIL.n124 VTAIL.n102 171.744
R162 VTAIL.n117 VTAIL.n102 171.744
R163 VTAIL.n117 VTAIL.n116 171.744
R164 VTAIL.n116 VTAIL.n106 171.744
R165 VTAIL.n109 VTAIL.n106 171.744
R166 VTAIL.n272 VTAIL.t2 85.8723
R167 VTAIL.n26 VTAIL.t1 85.8723
R168 VTAIL.n191 VTAIL.t0 85.8723
R169 VTAIL.n109 VTAIL.t3 85.8723
R170 VTAIL.n327 VTAIL.n326 35.4823
R171 VTAIL.n81 VTAIL.n80 35.4823
R172 VTAIL.n245 VTAIL.n244 35.4823
R173 VTAIL.n163 VTAIL.n162 35.4823
R174 VTAIL.n163 VTAIL.n81 26.7548
R175 VTAIL.n327 VTAIL.n245 25.9531
R176 VTAIL.n273 VTAIL.n271 16.3895
R177 VTAIL.n27 VTAIL.n25 16.3895
R178 VTAIL.n192 VTAIL.n190 16.3895
R179 VTAIL.n110 VTAIL.n108 16.3895
R180 VTAIL.n320 VTAIL.n319 13.1884
R181 VTAIL.n74 VTAIL.n73 13.1884
R182 VTAIL.n238 VTAIL.n237 13.1884
R183 VTAIL.n156 VTAIL.n155 13.1884
R184 VTAIL.n274 VTAIL.n270 12.8005
R185 VTAIL.n318 VTAIL.n250 12.8005
R186 VTAIL.n323 VTAIL.n248 12.8005
R187 VTAIL.n28 VTAIL.n24 12.8005
R188 VTAIL.n72 VTAIL.n4 12.8005
R189 VTAIL.n77 VTAIL.n2 12.8005
R190 VTAIL.n241 VTAIL.n166 12.8005
R191 VTAIL.n236 VTAIL.n168 12.8005
R192 VTAIL.n193 VTAIL.n189 12.8005
R193 VTAIL.n159 VTAIL.n84 12.8005
R194 VTAIL.n154 VTAIL.n86 12.8005
R195 VTAIL.n111 VTAIL.n107 12.8005
R196 VTAIL.n278 VTAIL.n277 12.0247
R197 VTAIL.n315 VTAIL.n314 12.0247
R198 VTAIL.n324 VTAIL.n246 12.0247
R199 VTAIL.n32 VTAIL.n31 12.0247
R200 VTAIL.n69 VTAIL.n68 12.0247
R201 VTAIL.n78 VTAIL.n0 12.0247
R202 VTAIL.n242 VTAIL.n164 12.0247
R203 VTAIL.n233 VTAIL.n232 12.0247
R204 VTAIL.n197 VTAIL.n196 12.0247
R205 VTAIL.n160 VTAIL.n82 12.0247
R206 VTAIL.n151 VTAIL.n150 12.0247
R207 VTAIL.n115 VTAIL.n114 12.0247
R208 VTAIL.n281 VTAIL.n268 11.249
R209 VTAIL.n310 VTAIL.n252 11.249
R210 VTAIL.n35 VTAIL.n22 11.249
R211 VTAIL.n64 VTAIL.n6 11.249
R212 VTAIL.n229 VTAIL.n170 11.249
R213 VTAIL.n200 VTAIL.n187 11.249
R214 VTAIL.n147 VTAIL.n88 11.249
R215 VTAIL.n118 VTAIL.n105 11.249
R216 VTAIL.n282 VTAIL.n266 10.4732
R217 VTAIL.n309 VTAIL.n254 10.4732
R218 VTAIL.n36 VTAIL.n20 10.4732
R219 VTAIL.n63 VTAIL.n8 10.4732
R220 VTAIL.n228 VTAIL.n173 10.4732
R221 VTAIL.n201 VTAIL.n185 10.4732
R222 VTAIL.n146 VTAIL.n91 10.4732
R223 VTAIL.n119 VTAIL.n103 10.4732
R224 VTAIL.n286 VTAIL.n285 9.69747
R225 VTAIL.n306 VTAIL.n305 9.69747
R226 VTAIL.n40 VTAIL.n39 9.69747
R227 VTAIL.n60 VTAIL.n59 9.69747
R228 VTAIL.n225 VTAIL.n224 9.69747
R229 VTAIL.n205 VTAIL.n204 9.69747
R230 VTAIL.n143 VTAIL.n142 9.69747
R231 VTAIL.n123 VTAIL.n122 9.69747
R232 VTAIL.n326 VTAIL.n325 9.45567
R233 VTAIL.n80 VTAIL.n79 9.45567
R234 VTAIL.n244 VTAIL.n243 9.45567
R235 VTAIL.n162 VTAIL.n161 9.45567
R236 VTAIL.n325 VTAIL.n324 9.3005
R237 VTAIL.n248 VTAIL.n247 9.3005
R238 VTAIL.n293 VTAIL.n292 9.3005
R239 VTAIL.n291 VTAIL.n290 9.3005
R240 VTAIL.n264 VTAIL.n263 9.3005
R241 VTAIL.n285 VTAIL.n284 9.3005
R242 VTAIL.n283 VTAIL.n282 9.3005
R243 VTAIL.n268 VTAIL.n267 9.3005
R244 VTAIL.n277 VTAIL.n276 9.3005
R245 VTAIL.n275 VTAIL.n274 9.3005
R246 VTAIL.n260 VTAIL.n259 9.3005
R247 VTAIL.n299 VTAIL.n298 9.3005
R248 VTAIL.n301 VTAIL.n300 9.3005
R249 VTAIL.n256 VTAIL.n255 9.3005
R250 VTAIL.n307 VTAIL.n306 9.3005
R251 VTAIL.n309 VTAIL.n308 9.3005
R252 VTAIL.n252 VTAIL.n251 9.3005
R253 VTAIL.n316 VTAIL.n315 9.3005
R254 VTAIL.n318 VTAIL.n317 9.3005
R255 VTAIL.n79 VTAIL.n78 9.3005
R256 VTAIL.n2 VTAIL.n1 9.3005
R257 VTAIL.n47 VTAIL.n46 9.3005
R258 VTAIL.n45 VTAIL.n44 9.3005
R259 VTAIL.n18 VTAIL.n17 9.3005
R260 VTAIL.n39 VTAIL.n38 9.3005
R261 VTAIL.n37 VTAIL.n36 9.3005
R262 VTAIL.n22 VTAIL.n21 9.3005
R263 VTAIL.n31 VTAIL.n30 9.3005
R264 VTAIL.n29 VTAIL.n28 9.3005
R265 VTAIL.n14 VTAIL.n13 9.3005
R266 VTAIL.n53 VTAIL.n52 9.3005
R267 VTAIL.n55 VTAIL.n54 9.3005
R268 VTAIL.n10 VTAIL.n9 9.3005
R269 VTAIL.n61 VTAIL.n60 9.3005
R270 VTAIL.n63 VTAIL.n62 9.3005
R271 VTAIL.n6 VTAIL.n5 9.3005
R272 VTAIL.n70 VTAIL.n69 9.3005
R273 VTAIL.n72 VTAIL.n71 9.3005
R274 VTAIL.n218 VTAIL.n217 9.3005
R275 VTAIL.n220 VTAIL.n219 9.3005
R276 VTAIL.n175 VTAIL.n174 9.3005
R277 VTAIL.n226 VTAIL.n225 9.3005
R278 VTAIL.n228 VTAIL.n227 9.3005
R279 VTAIL.n170 VTAIL.n169 9.3005
R280 VTAIL.n234 VTAIL.n233 9.3005
R281 VTAIL.n236 VTAIL.n235 9.3005
R282 VTAIL.n243 VTAIL.n242 9.3005
R283 VTAIL.n166 VTAIL.n165 9.3005
R284 VTAIL.n179 VTAIL.n178 9.3005
R285 VTAIL.n212 VTAIL.n211 9.3005
R286 VTAIL.n210 VTAIL.n209 9.3005
R287 VTAIL.n183 VTAIL.n182 9.3005
R288 VTAIL.n204 VTAIL.n203 9.3005
R289 VTAIL.n202 VTAIL.n201 9.3005
R290 VTAIL.n187 VTAIL.n186 9.3005
R291 VTAIL.n196 VTAIL.n195 9.3005
R292 VTAIL.n194 VTAIL.n193 9.3005
R293 VTAIL.n136 VTAIL.n135 9.3005
R294 VTAIL.n138 VTAIL.n137 9.3005
R295 VTAIL.n93 VTAIL.n92 9.3005
R296 VTAIL.n144 VTAIL.n143 9.3005
R297 VTAIL.n146 VTAIL.n145 9.3005
R298 VTAIL.n88 VTAIL.n87 9.3005
R299 VTAIL.n152 VTAIL.n151 9.3005
R300 VTAIL.n154 VTAIL.n153 9.3005
R301 VTAIL.n161 VTAIL.n160 9.3005
R302 VTAIL.n84 VTAIL.n83 9.3005
R303 VTAIL.n97 VTAIL.n96 9.3005
R304 VTAIL.n130 VTAIL.n129 9.3005
R305 VTAIL.n128 VTAIL.n127 9.3005
R306 VTAIL.n101 VTAIL.n100 9.3005
R307 VTAIL.n122 VTAIL.n121 9.3005
R308 VTAIL.n120 VTAIL.n119 9.3005
R309 VTAIL.n105 VTAIL.n104 9.3005
R310 VTAIL.n114 VTAIL.n113 9.3005
R311 VTAIL.n112 VTAIL.n111 9.3005
R312 VTAIL.n289 VTAIL.n264 8.92171
R313 VTAIL.n302 VTAIL.n256 8.92171
R314 VTAIL.n43 VTAIL.n18 8.92171
R315 VTAIL.n56 VTAIL.n10 8.92171
R316 VTAIL.n221 VTAIL.n175 8.92171
R317 VTAIL.n208 VTAIL.n183 8.92171
R318 VTAIL.n139 VTAIL.n93 8.92171
R319 VTAIL.n126 VTAIL.n101 8.92171
R320 VTAIL.n290 VTAIL.n262 8.14595
R321 VTAIL.n301 VTAIL.n258 8.14595
R322 VTAIL.n44 VTAIL.n16 8.14595
R323 VTAIL.n55 VTAIL.n12 8.14595
R324 VTAIL.n220 VTAIL.n177 8.14595
R325 VTAIL.n209 VTAIL.n181 8.14595
R326 VTAIL.n138 VTAIL.n95 8.14595
R327 VTAIL.n127 VTAIL.n99 8.14595
R328 VTAIL.n294 VTAIL.n293 7.3702
R329 VTAIL.n298 VTAIL.n297 7.3702
R330 VTAIL.n48 VTAIL.n47 7.3702
R331 VTAIL.n52 VTAIL.n51 7.3702
R332 VTAIL.n217 VTAIL.n216 7.3702
R333 VTAIL.n213 VTAIL.n212 7.3702
R334 VTAIL.n135 VTAIL.n134 7.3702
R335 VTAIL.n131 VTAIL.n130 7.3702
R336 VTAIL.n294 VTAIL.n260 6.59444
R337 VTAIL.n297 VTAIL.n260 6.59444
R338 VTAIL.n48 VTAIL.n14 6.59444
R339 VTAIL.n51 VTAIL.n14 6.59444
R340 VTAIL.n216 VTAIL.n179 6.59444
R341 VTAIL.n213 VTAIL.n179 6.59444
R342 VTAIL.n134 VTAIL.n97 6.59444
R343 VTAIL.n131 VTAIL.n97 6.59444
R344 VTAIL.n293 VTAIL.n262 5.81868
R345 VTAIL.n298 VTAIL.n258 5.81868
R346 VTAIL.n47 VTAIL.n16 5.81868
R347 VTAIL.n52 VTAIL.n12 5.81868
R348 VTAIL.n217 VTAIL.n177 5.81868
R349 VTAIL.n212 VTAIL.n181 5.81868
R350 VTAIL.n135 VTAIL.n95 5.81868
R351 VTAIL.n130 VTAIL.n99 5.81868
R352 VTAIL.n290 VTAIL.n289 5.04292
R353 VTAIL.n302 VTAIL.n301 5.04292
R354 VTAIL.n44 VTAIL.n43 5.04292
R355 VTAIL.n56 VTAIL.n55 5.04292
R356 VTAIL.n221 VTAIL.n220 5.04292
R357 VTAIL.n209 VTAIL.n208 5.04292
R358 VTAIL.n139 VTAIL.n138 5.04292
R359 VTAIL.n127 VTAIL.n126 5.04292
R360 VTAIL.n286 VTAIL.n264 4.26717
R361 VTAIL.n305 VTAIL.n256 4.26717
R362 VTAIL.n40 VTAIL.n18 4.26717
R363 VTAIL.n59 VTAIL.n10 4.26717
R364 VTAIL.n224 VTAIL.n175 4.26717
R365 VTAIL.n205 VTAIL.n183 4.26717
R366 VTAIL.n142 VTAIL.n93 4.26717
R367 VTAIL.n123 VTAIL.n101 4.26717
R368 VTAIL.n275 VTAIL.n271 3.70982
R369 VTAIL.n29 VTAIL.n25 3.70982
R370 VTAIL.n194 VTAIL.n190 3.70982
R371 VTAIL.n112 VTAIL.n108 3.70982
R372 VTAIL.n285 VTAIL.n266 3.49141
R373 VTAIL.n306 VTAIL.n254 3.49141
R374 VTAIL.n39 VTAIL.n20 3.49141
R375 VTAIL.n60 VTAIL.n8 3.49141
R376 VTAIL.n225 VTAIL.n173 3.49141
R377 VTAIL.n204 VTAIL.n185 3.49141
R378 VTAIL.n143 VTAIL.n91 3.49141
R379 VTAIL.n122 VTAIL.n103 3.49141
R380 VTAIL.n282 VTAIL.n281 2.71565
R381 VTAIL.n310 VTAIL.n309 2.71565
R382 VTAIL.n36 VTAIL.n35 2.71565
R383 VTAIL.n64 VTAIL.n63 2.71565
R384 VTAIL.n229 VTAIL.n228 2.71565
R385 VTAIL.n201 VTAIL.n200 2.71565
R386 VTAIL.n147 VTAIL.n146 2.71565
R387 VTAIL.n119 VTAIL.n118 2.71565
R388 VTAIL.n278 VTAIL.n268 1.93989
R389 VTAIL.n314 VTAIL.n252 1.93989
R390 VTAIL.n326 VTAIL.n246 1.93989
R391 VTAIL.n32 VTAIL.n22 1.93989
R392 VTAIL.n68 VTAIL.n6 1.93989
R393 VTAIL.n80 VTAIL.n0 1.93989
R394 VTAIL.n244 VTAIL.n164 1.93989
R395 VTAIL.n232 VTAIL.n170 1.93989
R396 VTAIL.n197 VTAIL.n187 1.93989
R397 VTAIL.n162 VTAIL.n82 1.93989
R398 VTAIL.n150 VTAIL.n88 1.93989
R399 VTAIL.n115 VTAIL.n105 1.93989
R400 VTAIL.n277 VTAIL.n270 1.16414
R401 VTAIL.n315 VTAIL.n250 1.16414
R402 VTAIL.n324 VTAIL.n323 1.16414
R403 VTAIL.n31 VTAIL.n24 1.16414
R404 VTAIL.n69 VTAIL.n4 1.16414
R405 VTAIL.n78 VTAIL.n77 1.16414
R406 VTAIL.n242 VTAIL.n241 1.16414
R407 VTAIL.n233 VTAIL.n168 1.16414
R408 VTAIL.n196 VTAIL.n189 1.16414
R409 VTAIL.n160 VTAIL.n159 1.16414
R410 VTAIL.n151 VTAIL.n86 1.16414
R411 VTAIL.n114 VTAIL.n107 1.16414
R412 VTAIL.n245 VTAIL.n163 0.87119
R413 VTAIL VTAIL.n81 0.728948
R414 VTAIL.n274 VTAIL.n273 0.388379
R415 VTAIL.n319 VTAIL.n318 0.388379
R416 VTAIL.n320 VTAIL.n248 0.388379
R417 VTAIL.n28 VTAIL.n27 0.388379
R418 VTAIL.n73 VTAIL.n72 0.388379
R419 VTAIL.n74 VTAIL.n2 0.388379
R420 VTAIL.n238 VTAIL.n166 0.388379
R421 VTAIL.n237 VTAIL.n236 0.388379
R422 VTAIL.n193 VTAIL.n192 0.388379
R423 VTAIL.n156 VTAIL.n84 0.388379
R424 VTAIL.n155 VTAIL.n154 0.388379
R425 VTAIL.n111 VTAIL.n110 0.388379
R426 VTAIL.n276 VTAIL.n275 0.155672
R427 VTAIL.n276 VTAIL.n267 0.155672
R428 VTAIL.n283 VTAIL.n267 0.155672
R429 VTAIL.n284 VTAIL.n283 0.155672
R430 VTAIL.n284 VTAIL.n263 0.155672
R431 VTAIL.n291 VTAIL.n263 0.155672
R432 VTAIL.n292 VTAIL.n291 0.155672
R433 VTAIL.n292 VTAIL.n259 0.155672
R434 VTAIL.n299 VTAIL.n259 0.155672
R435 VTAIL.n300 VTAIL.n299 0.155672
R436 VTAIL.n300 VTAIL.n255 0.155672
R437 VTAIL.n307 VTAIL.n255 0.155672
R438 VTAIL.n308 VTAIL.n307 0.155672
R439 VTAIL.n308 VTAIL.n251 0.155672
R440 VTAIL.n316 VTAIL.n251 0.155672
R441 VTAIL.n317 VTAIL.n316 0.155672
R442 VTAIL.n317 VTAIL.n247 0.155672
R443 VTAIL.n325 VTAIL.n247 0.155672
R444 VTAIL.n30 VTAIL.n29 0.155672
R445 VTAIL.n30 VTAIL.n21 0.155672
R446 VTAIL.n37 VTAIL.n21 0.155672
R447 VTAIL.n38 VTAIL.n37 0.155672
R448 VTAIL.n38 VTAIL.n17 0.155672
R449 VTAIL.n45 VTAIL.n17 0.155672
R450 VTAIL.n46 VTAIL.n45 0.155672
R451 VTAIL.n46 VTAIL.n13 0.155672
R452 VTAIL.n53 VTAIL.n13 0.155672
R453 VTAIL.n54 VTAIL.n53 0.155672
R454 VTAIL.n54 VTAIL.n9 0.155672
R455 VTAIL.n61 VTAIL.n9 0.155672
R456 VTAIL.n62 VTAIL.n61 0.155672
R457 VTAIL.n62 VTAIL.n5 0.155672
R458 VTAIL.n70 VTAIL.n5 0.155672
R459 VTAIL.n71 VTAIL.n70 0.155672
R460 VTAIL.n71 VTAIL.n1 0.155672
R461 VTAIL.n79 VTAIL.n1 0.155672
R462 VTAIL.n243 VTAIL.n165 0.155672
R463 VTAIL.n235 VTAIL.n165 0.155672
R464 VTAIL.n235 VTAIL.n234 0.155672
R465 VTAIL.n234 VTAIL.n169 0.155672
R466 VTAIL.n227 VTAIL.n169 0.155672
R467 VTAIL.n227 VTAIL.n226 0.155672
R468 VTAIL.n226 VTAIL.n174 0.155672
R469 VTAIL.n219 VTAIL.n174 0.155672
R470 VTAIL.n219 VTAIL.n218 0.155672
R471 VTAIL.n218 VTAIL.n178 0.155672
R472 VTAIL.n211 VTAIL.n178 0.155672
R473 VTAIL.n211 VTAIL.n210 0.155672
R474 VTAIL.n210 VTAIL.n182 0.155672
R475 VTAIL.n203 VTAIL.n182 0.155672
R476 VTAIL.n203 VTAIL.n202 0.155672
R477 VTAIL.n202 VTAIL.n186 0.155672
R478 VTAIL.n195 VTAIL.n186 0.155672
R479 VTAIL.n195 VTAIL.n194 0.155672
R480 VTAIL.n161 VTAIL.n83 0.155672
R481 VTAIL.n153 VTAIL.n83 0.155672
R482 VTAIL.n153 VTAIL.n152 0.155672
R483 VTAIL.n152 VTAIL.n87 0.155672
R484 VTAIL.n145 VTAIL.n87 0.155672
R485 VTAIL.n145 VTAIL.n144 0.155672
R486 VTAIL.n144 VTAIL.n92 0.155672
R487 VTAIL.n137 VTAIL.n92 0.155672
R488 VTAIL.n137 VTAIL.n136 0.155672
R489 VTAIL.n136 VTAIL.n96 0.155672
R490 VTAIL.n129 VTAIL.n96 0.155672
R491 VTAIL.n129 VTAIL.n128 0.155672
R492 VTAIL.n128 VTAIL.n100 0.155672
R493 VTAIL.n121 VTAIL.n100 0.155672
R494 VTAIL.n121 VTAIL.n120 0.155672
R495 VTAIL.n120 VTAIL.n104 0.155672
R496 VTAIL.n113 VTAIL.n104 0.155672
R497 VTAIL.n113 VTAIL.n112 0.155672
R498 VTAIL VTAIL.n327 0.142741
R499 VDD2.n157 VDD2.n81 756.745
R500 VDD2.n76 VDD2.n0 756.745
R501 VDD2.n158 VDD2.n157 585
R502 VDD2.n156 VDD2.n155 585
R503 VDD2.n154 VDD2.n84 585
R504 VDD2.n88 VDD2.n85 585
R505 VDD2.n149 VDD2.n148 585
R506 VDD2.n147 VDD2.n146 585
R507 VDD2.n90 VDD2.n89 585
R508 VDD2.n141 VDD2.n140 585
R509 VDD2.n139 VDD2.n138 585
R510 VDD2.n94 VDD2.n93 585
R511 VDD2.n133 VDD2.n132 585
R512 VDD2.n131 VDD2.n130 585
R513 VDD2.n98 VDD2.n97 585
R514 VDD2.n125 VDD2.n124 585
R515 VDD2.n123 VDD2.n122 585
R516 VDD2.n102 VDD2.n101 585
R517 VDD2.n117 VDD2.n116 585
R518 VDD2.n115 VDD2.n114 585
R519 VDD2.n106 VDD2.n105 585
R520 VDD2.n109 VDD2.n108 585
R521 VDD2.n27 VDD2.n26 585
R522 VDD2.n24 VDD2.n23 585
R523 VDD2.n33 VDD2.n32 585
R524 VDD2.n35 VDD2.n34 585
R525 VDD2.n20 VDD2.n19 585
R526 VDD2.n41 VDD2.n40 585
R527 VDD2.n43 VDD2.n42 585
R528 VDD2.n16 VDD2.n15 585
R529 VDD2.n49 VDD2.n48 585
R530 VDD2.n51 VDD2.n50 585
R531 VDD2.n12 VDD2.n11 585
R532 VDD2.n57 VDD2.n56 585
R533 VDD2.n59 VDD2.n58 585
R534 VDD2.n8 VDD2.n7 585
R535 VDD2.n65 VDD2.n64 585
R536 VDD2.n68 VDD2.n67 585
R537 VDD2.n66 VDD2.n4 585
R538 VDD2.n73 VDD2.n3 585
R539 VDD2.n75 VDD2.n74 585
R540 VDD2.n77 VDD2.n76 585
R541 VDD2.t0 VDD2.n107 327.466
R542 VDD2.t1 VDD2.n25 327.466
R543 VDD2.n157 VDD2.n156 171.744
R544 VDD2.n156 VDD2.n84 171.744
R545 VDD2.n88 VDD2.n84 171.744
R546 VDD2.n148 VDD2.n88 171.744
R547 VDD2.n148 VDD2.n147 171.744
R548 VDD2.n147 VDD2.n89 171.744
R549 VDD2.n140 VDD2.n89 171.744
R550 VDD2.n140 VDD2.n139 171.744
R551 VDD2.n139 VDD2.n93 171.744
R552 VDD2.n132 VDD2.n93 171.744
R553 VDD2.n132 VDD2.n131 171.744
R554 VDD2.n131 VDD2.n97 171.744
R555 VDD2.n124 VDD2.n97 171.744
R556 VDD2.n124 VDD2.n123 171.744
R557 VDD2.n123 VDD2.n101 171.744
R558 VDD2.n116 VDD2.n101 171.744
R559 VDD2.n116 VDD2.n115 171.744
R560 VDD2.n115 VDD2.n105 171.744
R561 VDD2.n108 VDD2.n105 171.744
R562 VDD2.n26 VDD2.n23 171.744
R563 VDD2.n33 VDD2.n23 171.744
R564 VDD2.n34 VDD2.n33 171.744
R565 VDD2.n34 VDD2.n19 171.744
R566 VDD2.n41 VDD2.n19 171.744
R567 VDD2.n42 VDD2.n41 171.744
R568 VDD2.n42 VDD2.n15 171.744
R569 VDD2.n49 VDD2.n15 171.744
R570 VDD2.n50 VDD2.n49 171.744
R571 VDD2.n50 VDD2.n11 171.744
R572 VDD2.n57 VDD2.n11 171.744
R573 VDD2.n58 VDD2.n57 171.744
R574 VDD2.n58 VDD2.n7 171.744
R575 VDD2.n65 VDD2.n7 171.744
R576 VDD2.n67 VDD2.n65 171.744
R577 VDD2.n67 VDD2.n66 171.744
R578 VDD2.n66 VDD2.n3 171.744
R579 VDD2.n75 VDD2.n3 171.744
R580 VDD2.n76 VDD2.n75 171.744
R581 VDD2.n162 VDD2.n80 90.2085
R582 VDD2.n108 VDD2.t0 85.8723
R583 VDD2.n26 VDD2.t1 85.8723
R584 VDD2.n162 VDD2.n161 52.1611
R585 VDD2.n109 VDD2.n107 16.3895
R586 VDD2.n27 VDD2.n25 16.3895
R587 VDD2.n155 VDD2.n154 13.1884
R588 VDD2.n74 VDD2.n73 13.1884
R589 VDD2.n158 VDD2.n83 12.8005
R590 VDD2.n153 VDD2.n85 12.8005
R591 VDD2.n110 VDD2.n106 12.8005
R592 VDD2.n28 VDD2.n24 12.8005
R593 VDD2.n72 VDD2.n4 12.8005
R594 VDD2.n77 VDD2.n2 12.8005
R595 VDD2.n159 VDD2.n81 12.0247
R596 VDD2.n150 VDD2.n149 12.0247
R597 VDD2.n114 VDD2.n113 12.0247
R598 VDD2.n32 VDD2.n31 12.0247
R599 VDD2.n69 VDD2.n68 12.0247
R600 VDD2.n78 VDD2.n0 12.0247
R601 VDD2.n146 VDD2.n87 11.249
R602 VDD2.n117 VDD2.n104 11.249
R603 VDD2.n35 VDD2.n22 11.249
R604 VDD2.n64 VDD2.n6 11.249
R605 VDD2.n145 VDD2.n90 10.4732
R606 VDD2.n118 VDD2.n102 10.4732
R607 VDD2.n36 VDD2.n20 10.4732
R608 VDD2.n63 VDD2.n8 10.4732
R609 VDD2.n142 VDD2.n141 9.69747
R610 VDD2.n122 VDD2.n121 9.69747
R611 VDD2.n40 VDD2.n39 9.69747
R612 VDD2.n60 VDD2.n59 9.69747
R613 VDD2.n161 VDD2.n160 9.45567
R614 VDD2.n80 VDD2.n79 9.45567
R615 VDD2.n135 VDD2.n134 9.3005
R616 VDD2.n137 VDD2.n136 9.3005
R617 VDD2.n92 VDD2.n91 9.3005
R618 VDD2.n143 VDD2.n142 9.3005
R619 VDD2.n145 VDD2.n144 9.3005
R620 VDD2.n87 VDD2.n86 9.3005
R621 VDD2.n151 VDD2.n150 9.3005
R622 VDD2.n153 VDD2.n152 9.3005
R623 VDD2.n160 VDD2.n159 9.3005
R624 VDD2.n83 VDD2.n82 9.3005
R625 VDD2.n96 VDD2.n95 9.3005
R626 VDD2.n129 VDD2.n128 9.3005
R627 VDD2.n127 VDD2.n126 9.3005
R628 VDD2.n100 VDD2.n99 9.3005
R629 VDD2.n121 VDD2.n120 9.3005
R630 VDD2.n119 VDD2.n118 9.3005
R631 VDD2.n104 VDD2.n103 9.3005
R632 VDD2.n113 VDD2.n112 9.3005
R633 VDD2.n111 VDD2.n110 9.3005
R634 VDD2.n79 VDD2.n78 9.3005
R635 VDD2.n2 VDD2.n1 9.3005
R636 VDD2.n47 VDD2.n46 9.3005
R637 VDD2.n45 VDD2.n44 9.3005
R638 VDD2.n18 VDD2.n17 9.3005
R639 VDD2.n39 VDD2.n38 9.3005
R640 VDD2.n37 VDD2.n36 9.3005
R641 VDD2.n22 VDD2.n21 9.3005
R642 VDD2.n31 VDD2.n30 9.3005
R643 VDD2.n29 VDD2.n28 9.3005
R644 VDD2.n14 VDD2.n13 9.3005
R645 VDD2.n53 VDD2.n52 9.3005
R646 VDD2.n55 VDD2.n54 9.3005
R647 VDD2.n10 VDD2.n9 9.3005
R648 VDD2.n61 VDD2.n60 9.3005
R649 VDD2.n63 VDD2.n62 9.3005
R650 VDD2.n6 VDD2.n5 9.3005
R651 VDD2.n70 VDD2.n69 9.3005
R652 VDD2.n72 VDD2.n71 9.3005
R653 VDD2.n138 VDD2.n92 8.92171
R654 VDD2.n125 VDD2.n100 8.92171
R655 VDD2.n43 VDD2.n18 8.92171
R656 VDD2.n56 VDD2.n10 8.92171
R657 VDD2.n137 VDD2.n94 8.14595
R658 VDD2.n126 VDD2.n98 8.14595
R659 VDD2.n44 VDD2.n16 8.14595
R660 VDD2.n55 VDD2.n12 8.14595
R661 VDD2.n134 VDD2.n133 7.3702
R662 VDD2.n130 VDD2.n129 7.3702
R663 VDD2.n48 VDD2.n47 7.3702
R664 VDD2.n52 VDD2.n51 7.3702
R665 VDD2.n133 VDD2.n96 6.59444
R666 VDD2.n130 VDD2.n96 6.59444
R667 VDD2.n48 VDD2.n14 6.59444
R668 VDD2.n51 VDD2.n14 6.59444
R669 VDD2.n134 VDD2.n94 5.81868
R670 VDD2.n129 VDD2.n98 5.81868
R671 VDD2.n47 VDD2.n16 5.81868
R672 VDD2.n52 VDD2.n12 5.81868
R673 VDD2.n138 VDD2.n137 5.04292
R674 VDD2.n126 VDD2.n125 5.04292
R675 VDD2.n44 VDD2.n43 5.04292
R676 VDD2.n56 VDD2.n55 5.04292
R677 VDD2.n141 VDD2.n92 4.26717
R678 VDD2.n122 VDD2.n100 4.26717
R679 VDD2.n40 VDD2.n18 4.26717
R680 VDD2.n59 VDD2.n10 4.26717
R681 VDD2.n111 VDD2.n107 3.70982
R682 VDD2.n29 VDD2.n25 3.70982
R683 VDD2.n142 VDD2.n90 3.49141
R684 VDD2.n121 VDD2.n102 3.49141
R685 VDD2.n39 VDD2.n20 3.49141
R686 VDD2.n60 VDD2.n8 3.49141
R687 VDD2.n146 VDD2.n145 2.71565
R688 VDD2.n118 VDD2.n117 2.71565
R689 VDD2.n36 VDD2.n35 2.71565
R690 VDD2.n64 VDD2.n63 2.71565
R691 VDD2.n161 VDD2.n81 1.93989
R692 VDD2.n149 VDD2.n87 1.93989
R693 VDD2.n114 VDD2.n104 1.93989
R694 VDD2.n32 VDD2.n22 1.93989
R695 VDD2.n68 VDD2.n6 1.93989
R696 VDD2.n80 VDD2.n0 1.93989
R697 VDD2.n159 VDD2.n158 1.16414
R698 VDD2.n150 VDD2.n85 1.16414
R699 VDD2.n113 VDD2.n106 1.16414
R700 VDD2.n31 VDD2.n24 1.16414
R701 VDD2.n69 VDD2.n4 1.16414
R702 VDD2.n78 VDD2.n77 1.16414
R703 VDD2.n155 VDD2.n83 0.388379
R704 VDD2.n154 VDD2.n153 0.388379
R705 VDD2.n110 VDD2.n109 0.388379
R706 VDD2.n28 VDD2.n27 0.388379
R707 VDD2.n73 VDD2.n72 0.388379
R708 VDD2.n74 VDD2.n2 0.388379
R709 VDD2 VDD2.n162 0.259121
R710 VDD2.n160 VDD2.n82 0.155672
R711 VDD2.n152 VDD2.n82 0.155672
R712 VDD2.n152 VDD2.n151 0.155672
R713 VDD2.n151 VDD2.n86 0.155672
R714 VDD2.n144 VDD2.n86 0.155672
R715 VDD2.n144 VDD2.n143 0.155672
R716 VDD2.n143 VDD2.n91 0.155672
R717 VDD2.n136 VDD2.n91 0.155672
R718 VDD2.n136 VDD2.n135 0.155672
R719 VDD2.n135 VDD2.n95 0.155672
R720 VDD2.n128 VDD2.n95 0.155672
R721 VDD2.n128 VDD2.n127 0.155672
R722 VDD2.n127 VDD2.n99 0.155672
R723 VDD2.n120 VDD2.n99 0.155672
R724 VDD2.n120 VDD2.n119 0.155672
R725 VDD2.n119 VDD2.n103 0.155672
R726 VDD2.n112 VDD2.n103 0.155672
R727 VDD2.n112 VDD2.n111 0.155672
R728 VDD2.n30 VDD2.n29 0.155672
R729 VDD2.n30 VDD2.n21 0.155672
R730 VDD2.n37 VDD2.n21 0.155672
R731 VDD2.n38 VDD2.n37 0.155672
R732 VDD2.n38 VDD2.n17 0.155672
R733 VDD2.n45 VDD2.n17 0.155672
R734 VDD2.n46 VDD2.n45 0.155672
R735 VDD2.n46 VDD2.n13 0.155672
R736 VDD2.n53 VDD2.n13 0.155672
R737 VDD2.n54 VDD2.n53 0.155672
R738 VDD2.n54 VDD2.n9 0.155672
R739 VDD2.n61 VDD2.n9 0.155672
R740 VDD2.n62 VDD2.n61 0.155672
R741 VDD2.n62 VDD2.n5 0.155672
R742 VDD2.n70 VDD2.n5 0.155672
R743 VDD2.n71 VDD2.n70 0.155672
R744 VDD2.n71 VDD2.n1 0.155672
R745 VDD2.n79 VDD2.n1 0.155672
R746 B.n112 B.t6 799.269
R747 B.n250 B.t3 799.269
R748 B.n40 B.t0 799.269
R749 B.n34 B.t9 799.269
R750 B.n329 B.n328 585
R751 B.n327 B.n82 585
R752 B.n326 B.n325 585
R753 B.n324 B.n83 585
R754 B.n323 B.n322 585
R755 B.n321 B.n84 585
R756 B.n320 B.n319 585
R757 B.n318 B.n85 585
R758 B.n317 B.n316 585
R759 B.n315 B.n86 585
R760 B.n314 B.n313 585
R761 B.n312 B.n87 585
R762 B.n311 B.n310 585
R763 B.n309 B.n88 585
R764 B.n308 B.n307 585
R765 B.n306 B.n89 585
R766 B.n305 B.n304 585
R767 B.n303 B.n90 585
R768 B.n302 B.n301 585
R769 B.n300 B.n91 585
R770 B.n299 B.n298 585
R771 B.n297 B.n92 585
R772 B.n296 B.n295 585
R773 B.n294 B.n93 585
R774 B.n293 B.n292 585
R775 B.n291 B.n94 585
R776 B.n290 B.n289 585
R777 B.n288 B.n95 585
R778 B.n287 B.n286 585
R779 B.n285 B.n96 585
R780 B.n284 B.n283 585
R781 B.n282 B.n97 585
R782 B.n281 B.n280 585
R783 B.n279 B.n98 585
R784 B.n278 B.n277 585
R785 B.n276 B.n99 585
R786 B.n275 B.n274 585
R787 B.n273 B.n100 585
R788 B.n272 B.n271 585
R789 B.n270 B.n101 585
R790 B.n269 B.n268 585
R791 B.n267 B.n102 585
R792 B.n266 B.n265 585
R793 B.n264 B.n103 585
R794 B.n263 B.n262 585
R795 B.n261 B.n104 585
R796 B.n260 B.n259 585
R797 B.n258 B.n105 585
R798 B.n257 B.n256 585
R799 B.n255 B.n106 585
R800 B.n254 B.n253 585
R801 B.n249 B.n107 585
R802 B.n248 B.n247 585
R803 B.n246 B.n108 585
R804 B.n245 B.n244 585
R805 B.n243 B.n109 585
R806 B.n242 B.n241 585
R807 B.n240 B.n110 585
R808 B.n239 B.n238 585
R809 B.n236 B.n111 585
R810 B.n235 B.n234 585
R811 B.n233 B.n114 585
R812 B.n232 B.n231 585
R813 B.n230 B.n115 585
R814 B.n229 B.n228 585
R815 B.n227 B.n116 585
R816 B.n226 B.n225 585
R817 B.n224 B.n117 585
R818 B.n223 B.n222 585
R819 B.n221 B.n118 585
R820 B.n220 B.n219 585
R821 B.n218 B.n119 585
R822 B.n217 B.n216 585
R823 B.n215 B.n120 585
R824 B.n214 B.n213 585
R825 B.n212 B.n121 585
R826 B.n211 B.n210 585
R827 B.n209 B.n122 585
R828 B.n208 B.n207 585
R829 B.n206 B.n123 585
R830 B.n205 B.n204 585
R831 B.n203 B.n124 585
R832 B.n202 B.n201 585
R833 B.n200 B.n125 585
R834 B.n199 B.n198 585
R835 B.n197 B.n126 585
R836 B.n196 B.n195 585
R837 B.n194 B.n127 585
R838 B.n193 B.n192 585
R839 B.n191 B.n128 585
R840 B.n190 B.n189 585
R841 B.n188 B.n129 585
R842 B.n187 B.n186 585
R843 B.n185 B.n130 585
R844 B.n184 B.n183 585
R845 B.n182 B.n131 585
R846 B.n181 B.n180 585
R847 B.n179 B.n132 585
R848 B.n178 B.n177 585
R849 B.n176 B.n133 585
R850 B.n175 B.n174 585
R851 B.n173 B.n134 585
R852 B.n172 B.n171 585
R853 B.n170 B.n135 585
R854 B.n169 B.n168 585
R855 B.n167 B.n136 585
R856 B.n166 B.n165 585
R857 B.n164 B.n137 585
R858 B.n163 B.n162 585
R859 B.n330 B.n81 585
R860 B.n332 B.n331 585
R861 B.n333 B.n80 585
R862 B.n335 B.n334 585
R863 B.n336 B.n79 585
R864 B.n338 B.n337 585
R865 B.n339 B.n78 585
R866 B.n341 B.n340 585
R867 B.n342 B.n77 585
R868 B.n344 B.n343 585
R869 B.n345 B.n76 585
R870 B.n347 B.n346 585
R871 B.n348 B.n75 585
R872 B.n350 B.n349 585
R873 B.n351 B.n74 585
R874 B.n353 B.n352 585
R875 B.n354 B.n73 585
R876 B.n356 B.n355 585
R877 B.n357 B.n72 585
R878 B.n359 B.n358 585
R879 B.n360 B.n71 585
R880 B.n362 B.n361 585
R881 B.n363 B.n70 585
R882 B.n365 B.n364 585
R883 B.n366 B.n69 585
R884 B.n368 B.n367 585
R885 B.n369 B.n68 585
R886 B.n371 B.n370 585
R887 B.n536 B.n535 585
R888 B.n534 B.n9 585
R889 B.n533 B.n532 585
R890 B.n531 B.n10 585
R891 B.n530 B.n529 585
R892 B.n528 B.n11 585
R893 B.n527 B.n526 585
R894 B.n525 B.n12 585
R895 B.n524 B.n523 585
R896 B.n522 B.n13 585
R897 B.n521 B.n520 585
R898 B.n519 B.n14 585
R899 B.n518 B.n517 585
R900 B.n516 B.n15 585
R901 B.n515 B.n514 585
R902 B.n513 B.n16 585
R903 B.n512 B.n511 585
R904 B.n510 B.n17 585
R905 B.n509 B.n508 585
R906 B.n507 B.n18 585
R907 B.n506 B.n505 585
R908 B.n504 B.n19 585
R909 B.n503 B.n502 585
R910 B.n501 B.n20 585
R911 B.n500 B.n499 585
R912 B.n498 B.n21 585
R913 B.n497 B.n496 585
R914 B.n495 B.n22 585
R915 B.n494 B.n493 585
R916 B.n492 B.n23 585
R917 B.n491 B.n490 585
R918 B.n489 B.n24 585
R919 B.n488 B.n487 585
R920 B.n486 B.n25 585
R921 B.n485 B.n484 585
R922 B.n483 B.n26 585
R923 B.n482 B.n481 585
R924 B.n480 B.n27 585
R925 B.n479 B.n478 585
R926 B.n477 B.n28 585
R927 B.n476 B.n475 585
R928 B.n474 B.n29 585
R929 B.n473 B.n472 585
R930 B.n471 B.n30 585
R931 B.n470 B.n469 585
R932 B.n468 B.n31 585
R933 B.n467 B.n466 585
R934 B.n465 B.n32 585
R935 B.n464 B.n463 585
R936 B.n462 B.n33 585
R937 B.n460 B.n459 585
R938 B.n458 B.n36 585
R939 B.n457 B.n456 585
R940 B.n455 B.n37 585
R941 B.n454 B.n453 585
R942 B.n452 B.n38 585
R943 B.n451 B.n450 585
R944 B.n449 B.n39 585
R945 B.n448 B.n447 585
R946 B.n446 B.n445 585
R947 B.n444 B.n43 585
R948 B.n443 B.n442 585
R949 B.n441 B.n44 585
R950 B.n440 B.n439 585
R951 B.n438 B.n45 585
R952 B.n437 B.n436 585
R953 B.n435 B.n46 585
R954 B.n434 B.n433 585
R955 B.n432 B.n47 585
R956 B.n431 B.n430 585
R957 B.n429 B.n48 585
R958 B.n428 B.n427 585
R959 B.n426 B.n49 585
R960 B.n425 B.n424 585
R961 B.n423 B.n50 585
R962 B.n422 B.n421 585
R963 B.n420 B.n51 585
R964 B.n419 B.n418 585
R965 B.n417 B.n52 585
R966 B.n416 B.n415 585
R967 B.n414 B.n53 585
R968 B.n413 B.n412 585
R969 B.n411 B.n54 585
R970 B.n410 B.n409 585
R971 B.n408 B.n55 585
R972 B.n407 B.n406 585
R973 B.n405 B.n56 585
R974 B.n404 B.n403 585
R975 B.n402 B.n57 585
R976 B.n401 B.n400 585
R977 B.n399 B.n58 585
R978 B.n398 B.n397 585
R979 B.n396 B.n59 585
R980 B.n395 B.n394 585
R981 B.n393 B.n60 585
R982 B.n392 B.n391 585
R983 B.n390 B.n61 585
R984 B.n389 B.n388 585
R985 B.n387 B.n62 585
R986 B.n386 B.n385 585
R987 B.n384 B.n63 585
R988 B.n383 B.n382 585
R989 B.n381 B.n64 585
R990 B.n380 B.n379 585
R991 B.n378 B.n65 585
R992 B.n377 B.n376 585
R993 B.n375 B.n66 585
R994 B.n374 B.n373 585
R995 B.n372 B.n67 585
R996 B.n537 B.n8 585
R997 B.n539 B.n538 585
R998 B.n540 B.n7 585
R999 B.n542 B.n541 585
R1000 B.n543 B.n6 585
R1001 B.n545 B.n544 585
R1002 B.n546 B.n5 585
R1003 B.n548 B.n547 585
R1004 B.n549 B.n4 585
R1005 B.n551 B.n550 585
R1006 B.n552 B.n3 585
R1007 B.n554 B.n553 585
R1008 B.n555 B.n0 585
R1009 B.n2 B.n1 585
R1010 B.n145 B.n144 585
R1011 B.n146 B.n143 585
R1012 B.n148 B.n147 585
R1013 B.n149 B.n142 585
R1014 B.n151 B.n150 585
R1015 B.n152 B.n141 585
R1016 B.n154 B.n153 585
R1017 B.n155 B.n140 585
R1018 B.n157 B.n156 585
R1019 B.n158 B.n139 585
R1020 B.n160 B.n159 585
R1021 B.n161 B.n138 585
R1022 B.n162 B.n161 550.159
R1023 B.n328 B.n81 550.159
R1024 B.n370 B.n67 550.159
R1025 B.n537 B.n536 550.159
R1026 B.n250 B.t4 444.303
R1027 B.n40 B.t2 444.303
R1028 B.n112 B.t7 444.301
R1029 B.n34 B.t11 444.301
R1030 B.n251 B.t5 426.265
R1031 B.n41 B.t1 426.265
R1032 B.n113 B.t8 426.265
R1033 B.n35 B.t10 426.265
R1034 B.n557 B.n556 256.663
R1035 B.n556 B.n555 235.042
R1036 B.n556 B.n2 235.042
R1037 B.n162 B.n137 163.367
R1038 B.n166 B.n137 163.367
R1039 B.n167 B.n166 163.367
R1040 B.n168 B.n167 163.367
R1041 B.n168 B.n135 163.367
R1042 B.n172 B.n135 163.367
R1043 B.n173 B.n172 163.367
R1044 B.n174 B.n173 163.367
R1045 B.n174 B.n133 163.367
R1046 B.n178 B.n133 163.367
R1047 B.n179 B.n178 163.367
R1048 B.n180 B.n179 163.367
R1049 B.n180 B.n131 163.367
R1050 B.n184 B.n131 163.367
R1051 B.n185 B.n184 163.367
R1052 B.n186 B.n185 163.367
R1053 B.n186 B.n129 163.367
R1054 B.n190 B.n129 163.367
R1055 B.n191 B.n190 163.367
R1056 B.n192 B.n191 163.367
R1057 B.n192 B.n127 163.367
R1058 B.n196 B.n127 163.367
R1059 B.n197 B.n196 163.367
R1060 B.n198 B.n197 163.367
R1061 B.n198 B.n125 163.367
R1062 B.n202 B.n125 163.367
R1063 B.n203 B.n202 163.367
R1064 B.n204 B.n203 163.367
R1065 B.n204 B.n123 163.367
R1066 B.n208 B.n123 163.367
R1067 B.n209 B.n208 163.367
R1068 B.n210 B.n209 163.367
R1069 B.n210 B.n121 163.367
R1070 B.n214 B.n121 163.367
R1071 B.n215 B.n214 163.367
R1072 B.n216 B.n215 163.367
R1073 B.n216 B.n119 163.367
R1074 B.n220 B.n119 163.367
R1075 B.n221 B.n220 163.367
R1076 B.n222 B.n221 163.367
R1077 B.n222 B.n117 163.367
R1078 B.n226 B.n117 163.367
R1079 B.n227 B.n226 163.367
R1080 B.n228 B.n227 163.367
R1081 B.n228 B.n115 163.367
R1082 B.n232 B.n115 163.367
R1083 B.n233 B.n232 163.367
R1084 B.n234 B.n233 163.367
R1085 B.n234 B.n111 163.367
R1086 B.n239 B.n111 163.367
R1087 B.n240 B.n239 163.367
R1088 B.n241 B.n240 163.367
R1089 B.n241 B.n109 163.367
R1090 B.n245 B.n109 163.367
R1091 B.n246 B.n245 163.367
R1092 B.n247 B.n246 163.367
R1093 B.n247 B.n107 163.367
R1094 B.n254 B.n107 163.367
R1095 B.n255 B.n254 163.367
R1096 B.n256 B.n255 163.367
R1097 B.n256 B.n105 163.367
R1098 B.n260 B.n105 163.367
R1099 B.n261 B.n260 163.367
R1100 B.n262 B.n261 163.367
R1101 B.n262 B.n103 163.367
R1102 B.n266 B.n103 163.367
R1103 B.n267 B.n266 163.367
R1104 B.n268 B.n267 163.367
R1105 B.n268 B.n101 163.367
R1106 B.n272 B.n101 163.367
R1107 B.n273 B.n272 163.367
R1108 B.n274 B.n273 163.367
R1109 B.n274 B.n99 163.367
R1110 B.n278 B.n99 163.367
R1111 B.n279 B.n278 163.367
R1112 B.n280 B.n279 163.367
R1113 B.n280 B.n97 163.367
R1114 B.n284 B.n97 163.367
R1115 B.n285 B.n284 163.367
R1116 B.n286 B.n285 163.367
R1117 B.n286 B.n95 163.367
R1118 B.n290 B.n95 163.367
R1119 B.n291 B.n290 163.367
R1120 B.n292 B.n291 163.367
R1121 B.n292 B.n93 163.367
R1122 B.n296 B.n93 163.367
R1123 B.n297 B.n296 163.367
R1124 B.n298 B.n297 163.367
R1125 B.n298 B.n91 163.367
R1126 B.n302 B.n91 163.367
R1127 B.n303 B.n302 163.367
R1128 B.n304 B.n303 163.367
R1129 B.n304 B.n89 163.367
R1130 B.n308 B.n89 163.367
R1131 B.n309 B.n308 163.367
R1132 B.n310 B.n309 163.367
R1133 B.n310 B.n87 163.367
R1134 B.n314 B.n87 163.367
R1135 B.n315 B.n314 163.367
R1136 B.n316 B.n315 163.367
R1137 B.n316 B.n85 163.367
R1138 B.n320 B.n85 163.367
R1139 B.n321 B.n320 163.367
R1140 B.n322 B.n321 163.367
R1141 B.n322 B.n83 163.367
R1142 B.n326 B.n83 163.367
R1143 B.n327 B.n326 163.367
R1144 B.n328 B.n327 163.367
R1145 B.n370 B.n369 163.367
R1146 B.n369 B.n368 163.367
R1147 B.n368 B.n69 163.367
R1148 B.n364 B.n69 163.367
R1149 B.n364 B.n363 163.367
R1150 B.n363 B.n362 163.367
R1151 B.n362 B.n71 163.367
R1152 B.n358 B.n71 163.367
R1153 B.n358 B.n357 163.367
R1154 B.n357 B.n356 163.367
R1155 B.n356 B.n73 163.367
R1156 B.n352 B.n73 163.367
R1157 B.n352 B.n351 163.367
R1158 B.n351 B.n350 163.367
R1159 B.n350 B.n75 163.367
R1160 B.n346 B.n75 163.367
R1161 B.n346 B.n345 163.367
R1162 B.n345 B.n344 163.367
R1163 B.n344 B.n77 163.367
R1164 B.n340 B.n77 163.367
R1165 B.n340 B.n339 163.367
R1166 B.n339 B.n338 163.367
R1167 B.n338 B.n79 163.367
R1168 B.n334 B.n79 163.367
R1169 B.n334 B.n333 163.367
R1170 B.n333 B.n332 163.367
R1171 B.n332 B.n81 163.367
R1172 B.n536 B.n9 163.367
R1173 B.n532 B.n9 163.367
R1174 B.n532 B.n531 163.367
R1175 B.n531 B.n530 163.367
R1176 B.n530 B.n11 163.367
R1177 B.n526 B.n11 163.367
R1178 B.n526 B.n525 163.367
R1179 B.n525 B.n524 163.367
R1180 B.n524 B.n13 163.367
R1181 B.n520 B.n13 163.367
R1182 B.n520 B.n519 163.367
R1183 B.n519 B.n518 163.367
R1184 B.n518 B.n15 163.367
R1185 B.n514 B.n15 163.367
R1186 B.n514 B.n513 163.367
R1187 B.n513 B.n512 163.367
R1188 B.n512 B.n17 163.367
R1189 B.n508 B.n17 163.367
R1190 B.n508 B.n507 163.367
R1191 B.n507 B.n506 163.367
R1192 B.n506 B.n19 163.367
R1193 B.n502 B.n19 163.367
R1194 B.n502 B.n501 163.367
R1195 B.n501 B.n500 163.367
R1196 B.n500 B.n21 163.367
R1197 B.n496 B.n21 163.367
R1198 B.n496 B.n495 163.367
R1199 B.n495 B.n494 163.367
R1200 B.n494 B.n23 163.367
R1201 B.n490 B.n23 163.367
R1202 B.n490 B.n489 163.367
R1203 B.n489 B.n488 163.367
R1204 B.n488 B.n25 163.367
R1205 B.n484 B.n25 163.367
R1206 B.n484 B.n483 163.367
R1207 B.n483 B.n482 163.367
R1208 B.n482 B.n27 163.367
R1209 B.n478 B.n27 163.367
R1210 B.n478 B.n477 163.367
R1211 B.n477 B.n476 163.367
R1212 B.n476 B.n29 163.367
R1213 B.n472 B.n29 163.367
R1214 B.n472 B.n471 163.367
R1215 B.n471 B.n470 163.367
R1216 B.n470 B.n31 163.367
R1217 B.n466 B.n31 163.367
R1218 B.n466 B.n465 163.367
R1219 B.n465 B.n464 163.367
R1220 B.n464 B.n33 163.367
R1221 B.n459 B.n33 163.367
R1222 B.n459 B.n458 163.367
R1223 B.n458 B.n457 163.367
R1224 B.n457 B.n37 163.367
R1225 B.n453 B.n37 163.367
R1226 B.n453 B.n452 163.367
R1227 B.n452 B.n451 163.367
R1228 B.n451 B.n39 163.367
R1229 B.n447 B.n39 163.367
R1230 B.n447 B.n446 163.367
R1231 B.n446 B.n43 163.367
R1232 B.n442 B.n43 163.367
R1233 B.n442 B.n441 163.367
R1234 B.n441 B.n440 163.367
R1235 B.n440 B.n45 163.367
R1236 B.n436 B.n45 163.367
R1237 B.n436 B.n435 163.367
R1238 B.n435 B.n434 163.367
R1239 B.n434 B.n47 163.367
R1240 B.n430 B.n47 163.367
R1241 B.n430 B.n429 163.367
R1242 B.n429 B.n428 163.367
R1243 B.n428 B.n49 163.367
R1244 B.n424 B.n49 163.367
R1245 B.n424 B.n423 163.367
R1246 B.n423 B.n422 163.367
R1247 B.n422 B.n51 163.367
R1248 B.n418 B.n51 163.367
R1249 B.n418 B.n417 163.367
R1250 B.n417 B.n416 163.367
R1251 B.n416 B.n53 163.367
R1252 B.n412 B.n53 163.367
R1253 B.n412 B.n411 163.367
R1254 B.n411 B.n410 163.367
R1255 B.n410 B.n55 163.367
R1256 B.n406 B.n55 163.367
R1257 B.n406 B.n405 163.367
R1258 B.n405 B.n404 163.367
R1259 B.n404 B.n57 163.367
R1260 B.n400 B.n57 163.367
R1261 B.n400 B.n399 163.367
R1262 B.n399 B.n398 163.367
R1263 B.n398 B.n59 163.367
R1264 B.n394 B.n59 163.367
R1265 B.n394 B.n393 163.367
R1266 B.n393 B.n392 163.367
R1267 B.n392 B.n61 163.367
R1268 B.n388 B.n61 163.367
R1269 B.n388 B.n387 163.367
R1270 B.n387 B.n386 163.367
R1271 B.n386 B.n63 163.367
R1272 B.n382 B.n63 163.367
R1273 B.n382 B.n381 163.367
R1274 B.n381 B.n380 163.367
R1275 B.n380 B.n65 163.367
R1276 B.n376 B.n65 163.367
R1277 B.n376 B.n375 163.367
R1278 B.n375 B.n374 163.367
R1279 B.n374 B.n67 163.367
R1280 B.n538 B.n537 163.367
R1281 B.n538 B.n7 163.367
R1282 B.n542 B.n7 163.367
R1283 B.n543 B.n542 163.367
R1284 B.n544 B.n543 163.367
R1285 B.n544 B.n5 163.367
R1286 B.n548 B.n5 163.367
R1287 B.n549 B.n548 163.367
R1288 B.n550 B.n549 163.367
R1289 B.n550 B.n3 163.367
R1290 B.n554 B.n3 163.367
R1291 B.n555 B.n554 163.367
R1292 B.n144 B.n2 163.367
R1293 B.n144 B.n143 163.367
R1294 B.n148 B.n143 163.367
R1295 B.n149 B.n148 163.367
R1296 B.n150 B.n149 163.367
R1297 B.n150 B.n141 163.367
R1298 B.n154 B.n141 163.367
R1299 B.n155 B.n154 163.367
R1300 B.n156 B.n155 163.367
R1301 B.n156 B.n139 163.367
R1302 B.n160 B.n139 163.367
R1303 B.n161 B.n160 163.367
R1304 B.n237 B.n113 59.5399
R1305 B.n252 B.n251 59.5399
R1306 B.n42 B.n41 59.5399
R1307 B.n461 B.n35 59.5399
R1308 B.n535 B.n8 35.7468
R1309 B.n372 B.n371 35.7468
R1310 B.n163 B.n138 35.7468
R1311 B.n330 B.n329 35.7468
R1312 B B.n557 18.0485
R1313 B.n113 B.n112 18.0369
R1314 B.n251 B.n250 18.0369
R1315 B.n41 B.n40 18.0369
R1316 B.n35 B.n34 18.0369
R1317 B.n539 B.n8 10.6151
R1318 B.n540 B.n539 10.6151
R1319 B.n541 B.n540 10.6151
R1320 B.n541 B.n6 10.6151
R1321 B.n545 B.n6 10.6151
R1322 B.n546 B.n545 10.6151
R1323 B.n547 B.n546 10.6151
R1324 B.n547 B.n4 10.6151
R1325 B.n551 B.n4 10.6151
R1326 B.n552 B.n551 10.6151
R1327 B.n553 B.n552 10.6151
R1328 B.n553 B.n0 10.6151
R1329 B.n535 B.n534 10.6151
R1330 B.n534 B.n533 10.6151
R1331 B.n533 B.n10 10.6151
R1332 B.n529 B.n10 10.6151
R1333 B.n529 B.n528 10.6151
R1334 B.n528 B.n527 10.6151
R1335 B.n527 B.n12 10.6151
R1336 B.n523 B.n12 10.6151
R1337 B.n523 B.n522 10.6151
R1338 B.n522 B.n521 10.6151
R1339 B.n521 B.n14 10.6151
R1340 B.n517 B.n14 10.6151
R1341 B.n517 B.n516 10.6151
R1342 B.n516 B.n515 10.6151
R1343 B.n515 B.n16 10.6151
R1344 B.n511 B.n16 10.6151
R1345 B.n511 B.n510 10.6151
R1346 B.n510 B.n509 10.6151
R1347 B.n509 B.n18 10.6151
R1348 B.n505 B.n18 10.6151
R1349 B.n505 B.n504 10.6151
R1350 B.n504 B.n503 10.6151
R1351 B.n503 B.n20 10.6151
R1352 B.n499 B.n20 10.6151
R1353 B.n499 B.n498 10.6151
R1354 B.n498 B.n497 10.6151
R1355 B.n497 B.n22 10.6151
R1356 B.n493 B.n22 10.6151
R1357 B.n493 B.n492 10.6151
R1358 B.n492 B.n491 10.6151
R1359 B.n491 B.n24 10.6151
R1360 B.n487 B.n24 10.6151
R1361 B.n487 B.n486 10.6151
R1362 B.n486 B.n485 10.6151
R1363 B.n485 B.n26 10.6151
R1364 B.n481 B.n26 10.6151
R1365 B.n481 B.n480 10.6151
R1366 B.n480 B.n479 10.6151
R1367 B.n479 B.n28 10.6151
R1368 B.n475 B.n28 10.6151
R1369 B.n475 B.n474 10.6151
R1370 B.n474 B.n473 10.6151
R1371 B.n473 B.n30 10.6151
R1372 B.n469 B.n30 10.6151
R1373 B.n469 B.n468 10.6151
R1374 B.n468 B.n467 10.6151
R1375 B.n467 B.n32 10.6151
R1376 B.n463 B.n32 10.6151
R1377 B.n463 B.n462 10.6151
R1378 B.n460 B.n36 10.6151
R1379 B.n456 B.n36 10.6151
R1380 B.n456 B.n455 10.6151
R1381 B.n455 B.n454 10.6151
R1382 B.n454 B.n38 10.6151
R1383 B.n450 B.n38 10.6151
R1384 B.n450 B.n449 10.6151
R1385 B.n449 B.n448 10.6151
R1386 B.n445 B.n444 10.6151
R1387 B.n444 B.n443 10.6151
R1388 B.n443 B.n44 10.6151
R1389 B.n439 B.n44 10.6151
R1390 B.n439 B.n438 10.6151
R1391 B.n438 B.n437 10.6151
R1392 B.n437 B.n46 10.6151
R1393 B.n433 B.n46 10.6151
R1394 B.n433 B.n432 10.6151
R1395 B.n432 B.n431 10.6151
R1396 B.n431 B.n48 10.6151
R1397 B.n427 B.n48 10.6151
R1398 B.n427 B.n426 10.6151
R1399 B.n426 B.n425 10.6151
R1400 B.n425 B.n50 10.6151
R1401 B.n421 B.n50 10.6151
R1402 B.n421 B.n420 10.6151
R1403 B.n420 B.n419 10.6151
R1404 B.n419 B.n52 10.6151
R1405 B.n415 B.n52 10.6151
R1406 B.n415 B.n414 10.6151
R1407 B.n414 B.n413 10.6151
R1408 B.n413 B.n54 10.6151
R1409 B.n409 B.n54 10.6151
R1410 B.n409 B.n408 10.6151
R1411 B.n408 B.n407 10.6151
R1412 B.n407 B.n56 10.6151
R1413 B.n403 B.n56 10.6151
R1414 B.n403 B.n402 10.6151
R1415 B.n402 B.n401 10.6151
R1416 B.n401 B.n58 10.6151
R1417 B.n397 B.n58 10.6151
R1418 B.n397 B.n396 10.6151
R1419 B.n396 B.n395 10.6151
R1420 B.n395 B.n60 10.6151
R1421 B.n391 B.n60 10.6151
R1422 B.n391 B.n390 10.6151
R1423 B.n390 B.n389 10.6151
R1424 B.n389 B.n62 10.6151
R1425 B.n385 B.n62 10.6151
R1426 B.n385 B.n384 10.6151
R1427 B.n384 B.n383 10.6151
R1428 B.n383 B.n64 10.6151
R1429 B.n379 B.n64 10.6151
R1430 B.n379 B.n378 10.6151
R1431 B.n378 B.n377 10.6151
R1432 B.n377 B.n66 10.6151
R1433 B.n373 B.n66 10.6151
R1434 B.n373 B.n372 10.6151
R1435 B.n371 B.n68 10.6151
R1436 B.n367 B.n68 10.6151
R1437 B.n367 B.n366 10.6151
R1438 B.n366 B.n365 10.6151
R1439 B.n365 B.n70 10.6151
R1440 B.n361 B.n70 10.6151
R1441 B.n361 B.n360 10.6151
R1442 B.n360 B.n359 10.6151
R1443 B.n359 B.n72 10.6151
R1444 B.n355 B.n72 10.6151
R1445 B.n355 B.n354 10.6151
R1446 B.n354 B.n353 10.6151
R1447 B.n353 B.n74 10.6151
R1448 B.n349 B.n74 10.6151
R1449 B.n349 B.n348 10.6151
R1450 B.n348 B.n347 10.6151
R1451 B.n347 B.n76 10.6151
R1452 B.n343 B.n76 10.6151
R1453 B.n343 B.n342 10.6151
R1454 B.n342 B.n341 10.6151
R1455 B.n341 B.n78 10.6151
R1456 B.n337 B.n78 10.6151
R1457 B.n337 B.n336 10.6151
R1458 B.n336 B.n335 10.6151
R1459 B.n335 B.n80 10.6151
R1460 B.n331 B.n80 10.6151
R1461 B.n331 B.n330 10.6151
R1462 B.n145 B.n1 10.6151
R1463 B.n146 B.n145 10.6151
R1464 B.n147 B.n146 10.6151
R1465 B.n147 B.n142 10.6151
R1466 B.n151 B.n142 10.6151
R1467 B.n152 B.n151 10.6151
R1468 B.n153 B.n152 10.6151
R1469 B.n153 B.n140 10.6151
R1470 B.n157 B.n140 10.6151
R1471 B.n158 B.n157 10.6151
R1472 B.n159 B.n158 10.6151
R1473 B.n159 B.n138 10.6151
R1474 B.n164 B.n163 10.6151
R1475 B.n165 B.n164 10.6151
R1476 B.n165 B.n136 10.6151
R1477 B.n169 B.n136 10.6151
R1478 B.n170 B.n169 10.6151
R1479 B.n171 B.n170 10.6151
R1480 B.n171 B.n134 10.6151
R1481 B.n175 B.n134 10.6151
R1482 B.n176 B.n175 10.6151
R1483 B.n177 B.n176 10.6151
R1484 B.n177 B.n132 10.6151
R1485 B.n181 B.n132 10.6151
R1486 B.n182 B.n181 10.6151
R1487 B.n183 B.n182 10.6151
R1488 B.n183 B.n130 10.6151
R1489 B.n187 B.n130 10.6151
R1490 B.n188 B.n187 10.6151
R1491 B.n189 B.n188 10.6151
R1492 B.n189 B.n128 10.6151
R1493 B.n193 B.n128 10.6151
R1494 B.n194 B.n193 10.6151
R1495 B.n195 B.n194 10.6151
R1496 B.n195 B.n126 10.6151
R1497 B.n199 B.n126 10.6151
R1498 B.n200 B.n199 10.6151
R1499 B.n201 B.n200 10.6151
R1500 B.n201 B.n124 10.6151
R1501 B.n205 B.n124 10.6151
R1502 B.n206 B.n205 10.6151
R1503 B.n207 B.n206 10.6151
R1504 B.n207 B.n122 10.6151
R1505 B.n211 B.n122 10.6151
R1506 B.n212 B.n211 10.6151
R1507 B.n213 B.n212 10.6151
R1508 B.n213 B.n120 10.6151
R1509 B.n217 B.n120 10.6151
R1510 B.n218 B.n217 10.6151
R1511 B.n219 B.n218 10.6151
R1512 B.n219 B.n118 10.6151
R1513 B.n223 B.n118 10.6151
R1514 B.n224 B.n223 10.6151
R1515 B.n225 B.n224 10.6151
R1516 B.n225 B.n116 10.6151
R1517 B.n229 B.n116 10.6151
R1518 B.n230 B.n229 10.6151
R1519 B.n231 B.n230 10.6151
R1520 B.n231 B.n114 10.6151
R1521 B.n235 B.n114 10.6151
R1522 B.n236 B.n235 10.6151
R1523 B.n238 B.n110 10.6151
R1524 B.n242 B.n110 10.6151
R1525 B.n243 B.n242 10.6151
R1526 B.n244 B.n243 10.6151
R1527 B.n244 B.n108 10.6151
R1528 B.n248 B.n108 10.6151
R1529 B.n249 B.n248 10.6151
R1530 B.n253 B.n249 10.6151
R1531 B.n257 B.n106 10.6151
R1532 B.n258 B.n257 10.6151
R1533 B.n259 B.n258 10.6151
R1534 B.n259 B.n104 10.6151
R1535 B.n263 B.n104 10.6151
R1536 B.n264 B.n263 10.6151
R1537 B.n265 B.n264 10.6151
R1538 B.n265 B.n102 10.6151
R1539 B.n269 B.n102 10.6151
R1540 B.n270 B.n269 10.6151
R1541 B.n271 B.n270 10.6151
R1542 B.n271 B.n100 10.6151
R1543 B.n275 B.n100 10.6151
R1544 B.n276 B.n275 10.6151
R1545 B.n277 B.n276 10.6151
R1546 B.n277 B.n98 10.6151
R1547 B.n281 B.n98 10.6151
R1548 B.n282 B.n281 10.6151
R1549 B.n283 B.n282 10.6151
R1550 B.n283 B.n96 10.6151
R1551 B.n287 B.n96 10.6151
R1552 B.n288 B.n287 10.6151
R1553 B.n289 B.n288 10.6151
R1554 B.n289 B.n94 10.6151
R1555 B.n293 B.n94 10.6151
R1556 B.n294 B.n293 10.6151
R1557 B.n295 B.n294 10.6151
R1558 B.n295 B.n92 10.6151
R1559 B.n299 B.n92 10.6151
R1560 B.n300 B.n299 10.6151
R1561 B.n301 B.n300 10.6151
R1562 B.n301 B.n90 10.6151
R1563 B.n305 B.n90 10.6151
R1564 B.n306 B.n305 10.6151
R1565 B.n307 B.n306 10.6151
R1566 B.n307 B.n88 10.6151
R1567 B.n311 B.n88 10.6151
R1568 B.n312 B.n311 10.6151
R1569 B.n313 B.n312 10.6151
R1570 B.n313 B.n86 10.6151
R1571 B.n317 B.n86 10.6151
R1572 B.n318 B.n317 10.6151
R1573 B.n319 B.n318 10.6151
R1574 B.n319 B.n84 10.6151
R1575 B.n323 B.n84 10.6151
R1576 B.n324 B.n323 10.6151
R1577 B.n325 B.n324 10.6151
R1578 B.n325 B.n82 10.6151
R1579 B.n329 B.n82 10.6151
R1580 B.n557 B.n0 8.11757
R1581 B.n557 B.n1 8.11757
R1582 B.n461 B.n460 7.18099
R1583 B.n448 B.n42 7.18099
R1584 B.n238 B.n237 7.18099
R1585 B.n253 B.n252 7.18099
R1586 B.n462 B.n461 3.43465
R1587 B.n445 B.n42 3.43465
R1588 B.n237 B.n236 3.43465
R1589 B.n252 B.n106 3.43465
R1590 VP.n0 VP.t1 863.538
R1591 VP.n0 VP.t0 822.043
R1592 VP VP.n0 0.0516364
R1593 VDD1.n76 VDD1.n0 756.745
R1594 VDD1.n157 VDD1.n81 756.745
R1595 VDD1.n77 VDD1.n76 585
R1596 VDD1.n75 VDD1.n74 585
R1597 VDD1.n73 VDD1.n3 585
R1598 VDD1.n7 VDD1.n4 585
R1599 VDD1.n68 VDD1.n67 585
R1600 VDD1.n66 VDD1.n65 585
R1601 VDD1.n9 VDD1.n8 585
R1602 VDD1.n60 VDD1.n59 585
R1603 VDD1.n58 VDD1.n57 585
R1604 VDD1.n13 VDD1.n12 585
R1605 VDD1.n52 VDD1.n51 585
R1606 VDD1.n50 VDD1.n49 585
R1607 VDD1.n17 VDD1.n16 585
R1608 VDD1.n44 VDD1.n43 585
R1609 VDD1.n42 VDD1.n41 585
R1610 VDD1.n21 VDD1.n20 585
R1611 VDD1.n36 VDD1.n35 585
R1612 VDD1.n34 VDD1.n33 585
R1613 VDD1.n25 VDD1.n24 585
R1614 VDD1.n28 VDD1.n27 585
R1615 VDD1.n108 VDD1.n107 585
R1616 VDD1.n105 VDD1.n104 585
R1617 VDD1.n114 VDD1.n113 585
R1618 VDD1.n116 VDD1.n115 585
R1619 VDD1.n101 VDD1.n100 585
R1620 VDD1.n122 VDD1.n121 585
R1621 VDD1.n124 VDD1.n123 585
R1622 VDD1.n97 VDD1.n96 585
R1623 VDD1.n130 VDD1.n129 585
R1624 VDD1.n132 VDD1.n131 585
R1625 VDD1.n93 VDD1.n92 585
R1626 VDD1.n138 VDD1.n137 585
R1627 VDD1.n140 VDD1.n139 585
R1628 VDD1.n89 VDD1.n88 585
R1629 VDD1.n146 VDD1.n145 585
R1630 VDD1.n149 VDD1.n148 585
R1631 VDD1.n147 VDD1.n85 585
R1632 VDD1.n154 VDD1.n84 585
R1633 VDD1.n156 VDD1.n155 585
R1634 VDD1.n158 VDD1.n157 585
R1635 VDD1.t0 VDD1.n26 327.466
R1636 VDD1.t1 VDD1.n106 327.466
R1637 VDD1.n76 VDD1.n75 171.744
R1638 VDD1.n75 VDD1.n3 171.744
R1639 VDD1.n7 VDD1.n3 171.744
R1640 VDD1.n67 VDD1.n7 171.744
R1641 VDD1.n67 VDD1.n66 171.744
R1642 VDD1.n66 VDD1.n8 171.744
R1643 VDD1.n59 VDD1.n8 171.744
R1644 VDD1.n59 VDD1.n58 171.744
R1645 VDD1.n58 VDD1.n12 171.744
R1646 VDD1.n51 VDD1.n12 171.744
R1647 VDD1.n51 VDD1.n50 171.744
R1648 VDD1.n50 VDD1.n16 171.744
R1649 VDD1.n43 VDD1.n16 171.744
R1650 VDD1.n43 VDD1.n42 171.744
R1651 VDD1.n42 VDD1.n20 171.744
R1652 VDD1.n35 VDD1.n20 171.744
R1653 VDD1.n35 VDD1.n34 171.744
R1654 VDD1.n34 VDD1.n24 171.744
R1655 VDD1.n27 VDD1.n24 171.744
R1656 VDD1.n107 VDD1.n104 171.744
R1657 VDD1.n114 VDD1.n104 171.744
R1658 VDD1.n115 VDD1.n114 171.744
R1659 VDD1.n115 VDD1.n100 171.744
R1660 VDD1.n122 VDD1.n100 171.744
R1661 VDD1.n123 VDD1.n122 171.744
R1662 VDD1.n123 VDD1.n96 171.744
R1663 VDD1.n130 VDD1.n96 171.744
R1664 VDD1.n131 VDD1.n130 171.744
R1665 VDD1.n131 VDD1.n92 171.744
R1666 VDD1.n138 VDD1.n92 171.744
R1667 VDD1.n139 VDD1.n138 171.744
R1668 VDD1.n139 VDD1.n88 171.744
R1669 VDD1.n146 VDD1.n88 171.744
R1670 VDD1.n148 VDD1.n146 171.744
R1671 VDD1.n148 VDD1.n147 171.744
R1672 VDD1.n147 VDD1.n84 171.744
R1673 VDD1.n156 VDD1.n84 171.744
R1674 VDD1.n157 VDD1.n156 171.744
R1675 VDD1 VDD1.n161 90.9337
R1676 VDD1.n27 VDD1.t0 85.8723
R1677 VDD1.n107 VDD1.t1 85.8723
R1678 VDD1 VDD1.n80 52.4197
R1679 VDD1.n28 VDD1.n26 16.3895
R1680 VDD1.n108 VDD1.n106 16.3895
R1681 VDD1.n74 VDD1.n73 13.1884
R1682 VDD1.n155 VDD1.n154 13.1884
R1683 VDD1.n77 VDD1.n2 12.8005
R1684 VDD1.n72 VDD1.n4 12.8005
R1685 VDD1.n29 VDD1.n25 12.8005
R1686 VDD1.n109 VDD1.n105 12.8005
R1687 VDD1.n153 VDD1.n85 12.8005
R1688 VDD1.n158 VDD1.n83 12.8005
R1689 VDD1.n78 VDD1.n0 12.0247
R1690 VDD1.n69 VDD1.n68 12.0247
R1691 VDD1.n33 VDD1.n32 12.0247
R1692 VDD1.n113 VDD1.n112 12.0247
R1693 VDD1.n150 VDD1.n149 12.0247
R1694 VDD1.n159 VDD1.n81 12.0247
R1695 VDD1.n65 VDD1.n6 11.249
R1696 VDD1.n36 VDD1.n23 11.249
R1697 VDD1.n116 VDD1.n103 11.249
R1698 VDD1.n145 VDD1.n87 11.249
R1699 VDD1.n64 VDD1.n9 10.4732
R1700 VDD1.n37 VDD1.n21 10.4732
R1701 VDD1.n117 VDD1.n101 10.4732
R1702 VDD1.n144 VDD1.n89 10.4732
R1703 VDD1.n61 VDD1.n60 9.69747
R1704 VDD1.n41 VDD1.n40 9.69747
R1705 VDD1.n121 VDD1.n120 9.69747
R1706 VDD1.n141 VDD1.n140 9.69747
R1707 VDD1.n80 VDD1.n79 9.45567
R1708 VDD1.n161 VDD1.n160 9.45567
R1709 VDD1.n54 VDD1.n53 9.3005
R1710 VDD1.n56 VDD1.n55 9.3005
R1711 VDD1.n11 VDD1.n10 9.3005
R1712 VDD1.n62 VDD1.n61 9.3005
R1713 VDD1.n64 VDD1.n63 9.3005
R1714 VDD1.n6 VDD1.n5 9.3005
R1715 VDD1.n70 VDD1.n69 9.3005
R1716 VDD1.n72 VDD1.n71 9.3005
R1717 VDD1.n79 VDD1.n78 9.3005
R1718 VDD1.n2 VDD1.n1 9.3005
R1719 VDD1.n15 VDD1.n14 9.3005
R1720 VDD1.n48 VDD1.n47 9.3005
R1721 VDD1.n46 VDD1.n45 9.3005
R1722 VDD1.n19 VDD1.n18 9.3005
R1723 VDD1.n40 VDD1.n39 9.3005
R1724 VDD1.n38 VDD1.n37 9.3005
R1725 VDD1.n23 VDD1.n22 9.3005
R1726 VDD1.n32 VDD1.n31 9.3005
R1727 VDD1.n30 VDD1.n29 9.3005
R1728 VDD1.n160 VDD1.n159 9.3005
R1729 VDD1.n83 VDD1.n82 9.3005
R1730 VDD1.n128 VDD1.n127 9.3005
R1731 VDD1.n126 VDD1.n125 9.3005
R1732 VDD1.n99 VDD1.n98 9.3005
R1733 VDD1.n120 VDD1.n119 9.3005
R1734 VDD1.n118 VDD1.n117 9.3005
R1735 VDD1.n103 VDD1.n102 9.3005
R1736 VDD1.n112 VDD1.n111 9.3005
R1737 VDD1.n110 VDD1.n109 9.3005
R1738 VDD1.n95 VDD1.n94 9.3005
R1739 VDD1.n134 VDD1.n133 9.3005
R1740 VDD1.n136 VDD1.n135 9.3005
R1741 VDD1.n91 VDD1.n90 9.3005
R1742 VDD1.n142 VDD1.n141 9.3005
R1743 VDD1.n144 VDD1.n143 9.3005
R1744 VDD1.n87 VDD1.n86 9.3005
R1745 VDD1.n151 VDD1.n150 9.3005
R1746 VDD1.n153 VDD1.n152 9.3005
R1747 VDD1.n57 VDD1.n11 8.92171
R1748 VDD1.n44 VDD1.n19 8.92171
R1749 VDD1.n124 VDD1.n99 8.92171
R1750 VDD1.n137 VDD1.n91 8.92171
R1751 VDD1.n56 VDD1.n13 8.14595
R1752 VDD1.n45 VDD1.n17 8.14595
R1753 VDD1.n125 VDD1.n97 8.14595
R1754 VDD1.n136 VDD1.n93 8.14595
R1755 VDD1.n53 VDD1.n52 7.3702
R1756 VDD1.n49 VDD1.n48 7.3702
R1757 VDD1.n129 VDD1.n128 7.3702
R1758 VDD1.n133 VDD1.n132 7.3702
R1759 VDD1.n52 VDD1.n15 6.59444
R1760 VDD1.n49 VDD1.n15 6.59444
R1761 VDD1.n129 VDD1.n95 6.59444
R1762 VDD1.n132 VDD1.n95 6.59444
R1763 VDD1.n53 VDD1.n13 5.81868
R1764 VDD1.n48 VDD1.n17 5.81868
R1765 VDD1.n128 VDD1.n97 5.81868
R1766 VDD1.n133 VDD1.n93 5.81868
R1767 VDD1.n57 VDD1.n56 5.04292
R1768 VDD1.n45 VDD1.n44 5.04292
R1769 VDD1.n125 VDD1.n124 5.04292
R1770 VDD1.n137 VDD1.n136 5.04292
R1771 VDD1.n60 VDD1.n11 4.26717
R1772 VDD1.n41 VDD1.n19 4.26717
R1773 VDD1.n121 VDD1.n99 4.26717
R1774 VDD1.n140 VDD1.n91 4.26717
R1775 VDD1.n30 VDD1.n26 3.70982
R1776 VDD1.n110 VDD1.n106 3.70982
R1777 VDD1.n61 VDD1.n9 3.49141
R1778 VDD1.n40 VDD1.n21 3.49141
R1779 VDD1.n120 VDD1.n101 3.49141
R1780 VDD1.n141 VDD1.n89 3.49141
R1781 VDD1.n65 VDD1.n64 2.71565
R1782 VDD1.n37 VDD1.n36 2.71565
R1783 VDD1.n117 VDD1.n116 2.71565
R1784 VDD1.n145 VDD1.n144 2.71565
R1785 VDD1.n80 VDD1.n0 1.93989
R1786 VDD1.n68 VDD1.n6 1.93989
R1787 VDD1.n33 VDD1.n23 1.93989
R1788 VDD1.n113 VDD1.n103 1.93989
R1789 VDD1.n149 VDD1.n87 1.93989
R1790 VDD1.n161 VDD1.n81 1.93989
R1791 VDD1.n78 VDD1.n77 1.16414
R1792 VDD1.n69 VDD1.n4 1.16414
R1793 VDD1.n32 VDD1.n25 1.16414
R1794 VDD1.n112 VDD1.n105 1.16414
R1795 VDD1.n150 VDD1.n85 1.16414
R1796 VDD1.n159 VDD1.n158 1.16414
R1797 VDD1.n74 VDD1.n2 0.388379
R1798 VDD1.n73 VDD1.n72 0.388379
R1799 VDD1.n29 VDD1.n28 0.388379
R1800 VDD1.n109 VDD1.n108 0.388379
R1801 VDD1.n154 VDD1.n153 0.388379
R1802 VDD1.n155 VDD1.n83 0.388379
R1803 VDD1.n79 VDD1.n1 0.155672
R1804 VDD1.n71 VDD1.n1 0.155672
R1805 VDD1.n71 VDD1.n70 0.155672
R1806 VDD1.n70 VDD1.n5 0.155672
R1807 VDD1.n63 VDD1.n5 0.155672
R1808 VDD1.n63 VDD1.n62 0.155672
R1809 VDD1.n62 VDD1.n10 0.155672
R1810 VDD1.n55 VDD1.n10 0.155672
R1811 VDD1.n55 VDD1.n54 0.155672
R1812 VDD1.n54 VDD1.n14 0.155672
R1813 VDD1.n47 VDD1.n14 0.155672
R1814 VDD1.n47 VDD1.n46 0.155672
R1815 VDD1.n46 VDD1.n18 0.155672
R1816 VDD1.n39 VDD1.n18 0.155672
R1817 VDD1.n39 VDD1.n38 0.155672
R1818 VDD1.n38 VDD1.n22 0.155672
R1819 VDD1.n31 VDD1.n22 0.155672
R1820 VDD1.n31 VDD1.n30 0.155672
R1821 VDD1.n111 VDD1.n110 0.155672
R1822 VDD1.n111 VDD1.n102 0.155672
R1823 VDD1.n118 VDD1.n102 0.155672
R1824 VDD1.n119 VDD1.n118 0.155672
R1825 VDD1.n119 VDD1.n98 0.155672
R1826 VDD1.n126 VDD1.n98 0.155672
R1827 VDD1.n127 VDD1.n126 0.155672
R1828 VDD1.n127 VDD1.n94 0.155672
R1829 VDD1.n134 VDD1.n94 0.155672
R1830 VDD1.n135 VDD1.n134 0.155672
R1831 VDD1.n135 VDD1.n90 0.155672
R1832 VDD1.n142 VDD1.n90 0.155672
R1833 VDD1.n143 VDD1.n142 0.155672
R1834 VDD1.n143 VDD1.n86 0.155672
R1835 VDD1.n151 VDD1.n86 0.155672
R1836 VDD1.n152 VDD1.n151 0.155672
R1837 VDD1.n152 VDD1.n82 0.155672
R1838 VDD1.n160 VDD1.n82 0.155672
C0 VDD2 VTAIL 6.96875f
C1 VDD2 VP 0.251294f
C2 w_n1342_n3934# VDD1 1.76982f
C3 VN w_n1342_n3934# 1.73933f
C4 VDD2 VDD1 0.453552f
C5 VDD2 VN 2.26225f
C6 B VTAIL 3.18303f
C7 B VP 1.00905f
C8 VDD2 w_n1342_n3934# 1.77346f
C9 B VDD1 1.6f
C10 VP VTAIL 1.62609f
C11 B VN 0.743122f
C12 VTAIL VDD1 6.93765f
C13 VP VDD1 2.35947f
C14 VN VTAIL 1.61133f
C15 VN VP 5.03691f
C16 B w_n1342_n3934# 7.43937f
C17 B VDD2 1.61383f
C18 VN VDD1 0.148543f
C19 VTAIL w_n1342_n3934# 3.40801f
C20 VP w_n1342_n3934# 1.90596f
C21 VDD2 VSUBS 0.838184f
C22 VDD1 VSUBS 3.564634f
C23 VTAIL VSUBS 0.840031f
C24 VN VSUBS 6.29698f
C25 VP VSUBS 1.18553f
C26 B VSUBS 2.661087f
C27 w_n1342_n3934# VSUBS 64.754196f
C28 VDD1.n0 VSUBS 0.022939f
C29 VDD1.n1 VSUBS 0.021203f
C30 VDD1.n2 VSUBS 0.011394f
C31 VDD1.n3 VSUBS 0.02693f
C32 VDD1.n4 VSUBS 0.012064f
C33 VDD1.n5 VSUBS 0.021203f
C34 VDD1.n6 VSUBS 0.011394f
C35 VDD1.n7 VSUBS 0.02693f
C36 VDD1.n8 VSUBS 0.02693f
C37 VDD1.n9 VSUBS 0.012064f
C38 VDD1.n10 VSUBS 0.021203f
C39 VDD1.n11 VSUBS 0.011394f
C40 VDD1.n12 VSUBS 0.02693f
C41 VDD1.n13 VSUBS 0.012064f
C42 VDD1.n14 VSUBS 0.021203f
C43 VDD1.n15 VSUBS 0.011394f
C44 VDD1.n16 VSUBS 0.02693f
C45 VDD1.n17 VSUBS 0.012064f
C46 VDD1.n18 VSUBS 0.021203f
C47 VDD1.n19 VSUBS 0.011394f
C48 VDD1.n20 VSUBS 0.02693f
C49 VDD1.n21 VSUBS 0.012064f
C50 VDD1.n22 VSUBS 0.021203f
C51 VDD1.n23 VSUBS 0.011394f
C52 VDD1.n24 VSUBS 0.02693f
C53 VDD1.n25 VSUBS 0.012064f
C54 VDD1.n26 VSUBS 0.148274f
C55 VDD1.t0 VSUBS 0.057642f
C56 VDD1.n27 VSUBS 0.020198f
C57 VDD1.n28 VSUBS 0.017132f
C58 VDD1.n29 VSUBS 0.011394f
C59 VDD1.n30 VSUBS 1.33556f
C60 VDD1.n31 VSUBS 0.021203f
C61 VDD1.n32 VSUBS 0.011394f
C62 VDD1.n33 VSUBS 0.012064f
C63 VDD1.n34 VSUBS 0.02693f
C64 VDD1.n35 VSUBS 0.02693f
C65 VDD1.n36 VSUBS 0.012064f
C66 VDD1.n37 VSUBS 0.011394f
C67 VDD1.n38 VSUBS 0.021203f
C68 VDD1.n39 VSUBS 0.021203f
C69 VDD1.n40 VSUBS 0.011394f
C70 VDD1.n41 VSUBS 0.012064f
C71 VDD1.n42 VSUBS 0.02693f
C72 VDD1.n43 VSUBS 0.02693f
C73 VDD1.n44 VSUBS 0.012064f
C74 VDD1.n45 VSUBS 0.011394f
C75 VDD1.n46 VSUBS 0.021203f
C76 VDD1.n47 VSUBS 0.021203f
C77 VDD1.n48 VSUBS 0.011394f
C78 VDD1.n49 VSUBS 0.012064f
C79 VDD1.n50 VSUBS 0.02693f
C80 VDD1.n51 VSUBS 0.02693f
C81 VDD1.n52 VSUBS 0.012064f
C82 VDD1.n53 VSUBS 0.011394f
C83 VDD1.n54 VSUBS 0.021203f
C84 VDD1.n55 VSUBS 0.021203f
C85 VDD1.n56 VSUBS 0.011394f
C86 VDD1.n57 VSUBS 0.012064f
C87 VDD1.n58 VSUBS 0.02693f
C88 VDD1.n59 VSUBS 0.02693f
C89 VDD1.n60 VSUBS 0.012064f
C90 VDD1.n61 VSUBS 0.011394f
C91 VDD1.n62 VSUBS 0.021203f
C92 VDD1.n63 VSUBS 0.021203f
C93 VDD1.n64 VSUBS 0.011394f
C94 VDD1.n65 VSUBS 0.012064f
C95 VDD1.n66 VSUBS 0.02693f
C96 VDD1.n67 VSUBS 0.02693f
C97 VDD1.n68 VSUBS 0.012064f
C98 VDD1.n69 VSUBS 0.011394f
C99 VDD1.n70 VSUBS 0.021203f
C100 VDD1.n71 VSUBS 0.021203f
C101 VDD1.n72 VSUBS 0.011394f
C102 VDD1.n73 VSUBS 0.011729f
C103 VDD1.n74 VSUBS 0.011729f
C104 VDD1.n75 VSUBS 0.02693f
C105 VDD1.n76 VSUBS 0.063975f
C106 VDD1.n77 VSUBS 0.012064f
C107 VDD1.n78 VSUBS 0.011394f
C108 VDD1.n79 VSUBS 0.053934f
C109 VDD1.n80 VSUBS 0.047171f
C110 VDD1.n81 VSUBS 0.022939f
C111 VDD1.n82 VSUBS 0.021203f
C112 VDD1.n83 VSUBS 0.011394f
C113 VDD1.n84 VSUBS 0.02693f
C114 VDD1.n85 VSUBS 0.012064f
C115 VDD1.n86 VSUBS 0.021203f
C116 VDD1.n87 VSUBS 0.011394f
C117 VDD1.n88 VSUBS 0.02693f
C118 VDD1.n89 VSUBS 0.012064f
C119 VDD1.n90 VSUBS 0.021203f
C120 VDD1.n91 VSUBS 0.011394f
C121 VDD1.n92 VSUBS 0.02693f
C122 VDD1.n93 VSUBS 0.012064f
C123 VDD1.n94 VSUBS 0.021203f
C124 VDD1.n95 VSUBS 0.011394f
C125 VDD1.n96 VSUBS 0.02693f
C126 VDD1.n97 VSUBS 0.012064f
C127 VDD1.n98 VSUBS 0.021203f
C128 VDD1.n99 VSUBS 0.011394f
C129 VDD1.n100 VSUBS 0.02693f
C130 VDD1.n101 VSUBS 0.012064f
C131 VDD1.n102 VSUBS 0.021203f
C132 VDD1.n103 VSUBS 0.011394f
C133 VDD1.n104 VSUBS 0.02693f
C134 VDD1.n105 VSUBS 0.012064f
C135 VDD1.n106 VSUBS 0.148274f
C136 VDD1.t1 VSUBS 0.057642f
C137 VDD1.n107 VSUBS 0.020198f
C138 VDD1.n108 VSUBS 0.017132f
C139 VDD1.n109 VSUBS 0.011394f
C140 VDD1.n110 VSUBS 1.33556f
C141 VDD1.n111 VSUBS 0.021203f
C142 VDD1.n112 VSUBS 0.011394f
C143 VDD1.n113 VSUBS 0.012064f
C144 VDD1.n114 VSUBS 0.02693f
C145 VDD1.n115 VSUBS 0.02693f
C146 VDD1.n116 VSUBS 0.012064f
C147 VDD1.n117 VSUBS 0.011394f
C148 VDD1.n118 VSUBS 0.021203f
C149 VDD1.n119 VSUBS 0.021203f
C150 VDD1.n120 VSUBS 0.011394f
C151 VDD1.n121 VSUBS 0.012064f
C152 VDD1.n122 VSUBS 0.02693f
C153 VDD1.n123 VSUBS 0.02693f
C154 VDD1.n124 VSUBS 0.012064f
C155 VDD1.n125 VSUBS 0.011394f
C156 VDD1.n126 VSUBS 0.021203f
C157 VDD1.n127 VSUBS 0.021203f
C158 VDD1.n128 VSUBS 0.011394f
C159 VDD1.n129 VSUBS 0.012064f
C160 VDD1.n130 VSUBS 0.02693f
C161 VDD1.n131 VSUBS 0.02693f
C162 VDD1.n132 VSUBS 0.012064f
C163 VDD1.n133 VSUBS 0.011394f
C164 VDD1.n134 VSUBS 0.021203f
C165 VDD1.n135 VSUBS 0.021203f
C166 VDD1.n136 VSUBS 0.011394f
C167 VDD1.n137 VSUBS 0.012064f
C168 VDD1.n138 VSUBS 0.02693f
C169 VDD1.n139 VSUBS 0.02693f
C170 VDD1.n140 VSUBS 0.012064f
C171 VDD1.n141 VSUBS 0.011394f
C172 VDD1.n142 VSUBS 0.021203f
C173 VDD1.n143 VSUBS 0.021203f
C174 VDD1.n144 VSUBS 0.011394f
C175 VDD1.n145 VSUBS 0.012064f
C176 VDD1.n146 VSUBS 0.02693f
C177 VDD1.n147 VSUBS 0.02693f
C178 VDD1.n148 VSUBS 0.02693f
C179 VDD1.n149 VSUBS 0.012064f
C180 VDD1.n150 VSUBS 0.011394f
C181 VDD1.n151 VSUBS 0.021203f
C182 VDD1.n152 VSUBS 0.021203f
C183 VDD1.n153 VSUBS 0.011394f
C184 VDD1.n154 VSUBS 0.011729f
C185 VDD1.n155 VSUBS 0.011729f
C186 VDD1.n156 VSUBS 0.02693f
C187 VDD1.n157 VSUBS 0.063975f
C188 VDD1.n158 VSUBS 0.012064f
C189 VDD1.n159 VSUBS 0.011394f
C190 VDD1.n160 VSUBS 0.053934f
C191 VDD1.n161 VSUBS 0.606122f
C192 VP.t1 VSUBS 1.43788f
C193 VP.t0 VSUBS 1.32477f
C194 VP.n0 VSUBS 4.62336f
C195 B.n0 VSUBS 0.006349f
C196 B.n1 VSUBS 0.006349f
C197 B.n2 VSUBS 0.009389f
C198 B.n3 VSUBS 0.007195f
C199 B.n4 VSUBS 0.007195f
C200 B.n5 VSUBS 0.007195f
C201 B.n6 VSUBS 0.007195f
C202 B.n7 VSUBS 0.007195f
C203 B.n8 VSUBS 0.017607f
C204 B.n9 VSUBS 0.007195f
C205 B.n10 VSUBS 0.007195f
C206 B.n11 VSUBS 0.007195f
C207 B.n12 VSUBS 0.007195f
C208 B.n13 VSUBS 0.007195f
C209 B.n14 VSUBS 0.007195f
C210 B.n15 VSUBS 0.007195f
C211 B.n16 VSUBS 0.007195f
C212 B.n17 VSUBS 0.007195f
C213 B.n18 VSUBS 0.007195f
C214 B.n19 VSUBS 0.007195f
C215 B.n20 VSUBS 0.007195f
C216 B.n21 VSUBS 0.007195f
C217 B.n22 VSUBS 0.007195f
C218 B.n23 VSUBS 0.007195f
C219 B.n24 VSUBS 0.007195f
C220 B.n25 VSUBS 0.007195f
C221 B.n26 VSUBS 0.007195f
C222 B.n27 VSUBS 0.007195f
C223 B.n28 VSUBS 0.007195f
C224 B.n29 VSUBS 0.007195f
C225 B.n30 VSUBS 0.007195f
C226 B.n31 VSUBS 0.007195f
C227 B.n32 VSUBS 0.007195f
C228 B.n33 VSUBS 0.007195f
C229 B.t10 VSUBS 0.282875f
C230 B.t11 VSUBS 0.294181f
C231 B.t9 VSUBS 0.368555f
C232 B.n34 VSUBS 0.370843f
C233 B.n35 VSUBS 0.288787f
C234 B.n36 VSUBS 0.007195f
C235 B.n37 VSUBS 0.007195f
C236 B.n38 VSUBS 0.007195f
C237 B.n39 VSUBS 0.007195f
C238 B.t1 VSUBS 0.282878f
C239 B.t2 VSUBS 0.294185f
C240 B.t0 VSUBS 0.368555f
C241 B.n40 VSUBS 0.37084f
C242 B.n41 VSUBS 0.288783f
C243 B.n42 VSUBS 0.01667f
C244 B.n43 VSUBS 0.007195f
C245 B.n44 VSUBS 0.007195f
C246 B.n45 VSUBS 0.007195f
C247 B.n46 VSUBS 0.007195f
C248 B.n47 VSUBS 0.007195f
C249 B.n48 VSUBS 0.007195f
C250 B.n49 VSUBS 0.007195f
C251 B.n50 VSUBS 0.007195f
C252 B.n51 VSUBS 0.007195f
C253 B.n52 VSUBS 0.007195f
C254 B.n53 VSUBS 0.007195f
C255 B.n54 VSUBS 0.007195f
C256 B.n55 VSUBS 0.007195f
C257 B.n56 VSUBS 0.007195f
C258 B.n57 VSUBS 0.007195f
C259 B.n58 VSUBS 0.007195f
C260 B.n59 VSUBS 0.007195f
C261 B.n60 VSUBS 0.007195f
C262 B.n61 VSUBS 0.007195f
C263 B.n62 VSUBS 0.007195f
C264 B.n63 VSUBS 0.007195f
C265 B.n64 VSUBS 0.007195f
C266 B.n65 VSUBS 0.007195f
C267 B.n66 VSUBS 0.007195f
C268 B.n67 VSUBS 0.018156f
C269 B.n68 VSUBS 0.007195f
C270 B.n69 VSUBS 0.007195f
C271 B.n70 VSUBS 0.007195f
C272 B.n71 VSUBS 0.007195f
C273 B.n72 VSUBS 0.007195f
C274 B.n73 VSUBS 0.007195f
C275 B.n74 VSUBS 0.007195f
C276 B.n75 VSUBS 0.007195f
C277 B.n76 VSUBS 0.007195f
C278 B.n77 VSUBS 0.007195f
C279 B.n78 VSUBS 0.007195f
C280 B.n79 VSUBS 0.007195f
C281 B.n80 VSUBS 0.007195f
C282 B.n81 VSUBS 0.017607f
C283 B.n82 VSUBS 0.007195f
C284 B.n83 VSUBS 0.007195f
C285 B.n84 VSUBS 0.007195f
C286 B.n85 VSUBS 0.007195f
C287 B.n86 VSUBS 0.007195f
C288 B.n87 VSUBS 0.007195f
C289 B.n88 VSUBS 0.007195f
C290 B.n89 VSUBS 0.007195f
C291 B.n90 VSUBS 0.007195f
C292 B.n91 VSUBS 0.007195f
C293 B.n92 VSUBS 0.007195f
C294 B.n93 VSUBS 0.007195f
C295 B.n94 VSUBS 0.007195f
C296 B.n95 VSUBS 0.007195f
C297 B.n96 VSUBS 0.007195f
C298 B.n97 VSUBS 0.007195f
C299 B.n98 VSUBS 0.007195f
C300 B.n99 VSUBS 0.007195f
C301 B.n100 VSUBS 0.007195f
C302 B.n101 VSUBS 0.007195f
C303 B.n102 VSUBS 0.007195f
C304 B.n103 VSUBS 0.007195f
C305 B.n104 VSUBS 0.007195f
C306 B.n105 VSUBS 0.007195f
C307 B.n106 VSUBS 0.004761f
C308 B.n107 VSUBS 0.007195f
C309 B.n108 VSUBS 0.007195f
C310 B.n109 VSUBS 0.007195f
C311 B.n110 VSUBS 0.007195f
C312 B.n111 VSUBS 0.007195f
C313 B.t8 VSUBS 0.282875f
C314 B.t7 VSUBS 0.294181f
C315 B.t6 VSUBS 0.368555f
C316 B.n112 VSUBS 0.370843f
C317 B.n113 VSUBS 0.288787f
C318 B.n114 VSUBS 0.007195f
C319 B.n115 VSUBS 0.007195f
C320 B.n116 VSUBS 0.007195f
C321 B.n117 VSUBS 0.007195f
C322 B.n118 VSUBS 0.007195f
C323 B.n119 VSUBS 0.007195f
C324 B.n120 VSUBS 0.007195f
C325 B.n121 VSUBS 0.007195f
C326 B.n122 VSUBS 0.007195f
C327 B.n123 VSUBS 0.007195f
C328 B.n124 VSUBS 0.007195f
C329 B.n125 VSUBS 0.007195f
C330 B.n126 VSUBS 0.007195f
C331 B.n127 VSUBS 0.007195f
C332 B.n128 VSUBS 0.007195f
C333 B.n129 VSUBS 0.007195f
C334 B.n130 VSUBS 0.007195f
C335 B.n131 VSUBS 0.007195f
C336 B.n132 VSUBS 0.007195f
C337 B.n133 VSUBS 0.007195f
C338 B.n134 VSUBS 0.007195f
C339 B.n135 VSUBS 0.007195f
C340 B.n136 VSUBS 0.007195f
C341 B.n137 VSUBS 0.007195f
C342 B.n138 VSUBS 0.017607f
C343 B.n139 VSUBS 0.007195f
C344 B.n140 VSUBS 0.007195f
C345 B.n141 VSUBS 0.007195f
C346 B.n142 VSUBS 0.007195f
C347 B.n143 VSUBS 0.007195f
C348 B.n144 VSUBS 0.007195f
C349 B.n145 VSUBS 0.007195f
C350 B.n146 VSUBS 0.007195f
C351 B.n147 VSUBS 0.007195f
C352 B.n148 VSUBS 0.007195f
C353 B.n149 VSUBS 0.007195f
C354 B.n150 VSUBS 0.007195f
C355 B.n151 VSUBS 0.007195f
C356 B.n152 VSUBS 0.007195f
C357 B.n153 VSUBS 0.007195f
C358 B.n154 VSUBS 0.007195f
C359 B.n155 VSUBS 0.007195f
C360 B.n156 VSUBS 0.007195f
C361 B.n157 VSUBS 0.007195f
C362 B.n158 VSUBS 0.007195f
C363 B.n159 VSUBS 0.007195f
C364 B.n160 VSUBS 0.007195f
C365 B.n161 VSUBS 0.017607f
C366 B.n162 VSUBS 0.018156f
C367 B.n163 VSUBS 0.018156f
C368 B.n164 VSUBS 0.007195f
C369 B.n165 VSUBS 0.007195f
C370 B.n166 VSUBS 0.007195f
C371 B.n167 VSUBS 0.007195f
C372 B.n168 VSUBS 0.007195f
C373 B.n169 VSUBS 0.007195f
C374 B.n170 VSUBS 0.007195f
C375 B.n171 VSUBS 0.007195f
C376 B.n172 VSUBS 0.007195f
C377 B.n173 VSUBS 0.007195f
C378 B.n174 VSUBS 0.007195f
C379 B.n175 VSUBS 0.007195f
C380 B.n176 VSUBS 0.007195f
C381 B.n177 VSUBS 0.007195f
C382 B.n178 VSUBS 0.007195f
C383 B.n179 VSUBS 0.007195f
C384 B.n180 VSUBS 0.007195f
C385 B.n181 VSUBS 0.007195f
C386 B.n182 VSUBS 0.007195f
C387 B.n183 VSUBS 0.007195f
C388 B.n184 VSUBS 0.007195f
C389 B.n185 VSUBS 0.007195f
C390 B.n186 VSUBS 0.007195f
C391 B.n187 VSUBS 0.007195f
C392 B.n188 VSUBS 0.007195f
C393 B.n189 VSUBS 0.007195f
C394 B.n190 VSUBS 0.007195f
C395 B.n191 VSUBS 0.007195f
C396 B.n192 VSUBS 0.007195f
C397 B.n193 VSUBS 0.007195f
C398 B.n194 VSUBS 0.007195f
C399 B.n195 VSUBS 0.007195f
C400 B.n196 VSUBS 0.007195f
C401 B.n197 VSUBS 0.007195f
C402 B.n198 VSUBS 0.007195f
C403 B.n199 VSUBS 0.007195f
C404 B.n200 VSUBS 0.007195f
C405 B.n201 VSUBS 0.007195f
C406 B.n202 VSUBS 0.007195f
C407 B.n203 VSUBS 0.007195f
C408 B.n204 VSUBS 0.007195f
C409 B.n205 VSUBS 0.007195f
C410 B.n206 VSUBS 0.007195f
C411 B.n207 VSUBS 0.007195f
C412 B.n208 VSUBS 0.007195f
C413 B.n209 VSUBS 0.007195f
C414 B.n210 VSUBS 0.007195f
C415 B.n211 VSUBS 0.007195f
C416 B.n212 VSUBS 0.007195f
C417 B.n213 VSUBS 0.007195f
C418 B.n214 VSUBS 0.007195f
C419 B.n215 VSUBS 0.007195f
C420 B.n216 VSUBS 0.007195f
C421 B.n217 VSUBS 0.007195f
C422 B.n218 VSUBS 0.007195f
C423 B.n219 VSUBS 0.007195f
C424 B.n220 VSUBS 0.007195f
C425 B.n221 VSUBS 0.007195f
C426 B.n222 VSUBS 0.007195f
C427 B.n223 VSUBS 0.007195f
C428 B.n224 VSUBS 0.007195f
C429 B.n225 VSUBS 0.007195f
C430 B.n226 VSUBS 0.007195f
C431 B.n227 VSUBS 0.007195f
C432 B.n228 VSUBS 0.007195f
C433 B.n229 VSUBS 0.007195f
C434 B.n230 VSUBS 0.007195f
C435 B.n231 VSUBS 0.007195f
C436 B.n232 VSUBS 0.007195f
C437 B.n233 VSUBS 0.007195f
C438 B.n234 VSUBS 0.007195f
C439 B.n235 VSUBS 0.007195f
C440 B.n236 VSUBS 0.004761f
C441 B.n237 VSUBS 0.01667f
C442 B.n238 VSUBS 0.006031f
C443 B.n239 VSUBS 0.007195f
C444 B.n240 VSUBS 0.007195f
C445 B.n241 VSUBS 0.007195f
C446 B.n242 VSUBS 0.007195f
C447 B.n243 VSUBS 0.007195f
C448 B.n244 VSUBS 0.007195f
C449 B.n245 VSUBS 0.007195f
C450 B.n246 VSUBS 0.007195f
C451 B.n247 VSUBS 0.007195f
C452 B.n248 VSUBS 0.007195f
C453 B.n249 VSUBS 0.007195f
C454 B.t5 VSUBS 0.282878f
C455 B.t4 VSUBS 0.294185f
C456 B.t3 VSUBS 0.368555f
C457 B.n250 VSUBS 0.37084f
C458 B.n251 VSUBS 0.288783f
C459 B.n252 VSUBS 0.01667f
C460 B.n253 VSUBS 0.006031f
C461 B.n254 VSUBS 0.007195f
C462 B.n255 VSUBS 0.007195f
C463 B.n256 VSUBS 0.007195f
C464 B.n257 VSUBS 0.007195f
C465 B.n258 VSUBS 0.007195f
C466 B.n259 VSUBS 0.007195f
C467 B.n260 VSUBS 0.007195f
C468 B.n261 VSUBS 0.007195f
C469 B.n262 VSUBS 0.007195f
C470 B.n263 VSUBS 0.007195f
C471 B.n264 VSUBS 0.007195f
C472 B.n265 VSUBS 0.007195f
C473 B.n266 VSUBS 0.007195f
C474 B.n267 VSUBS 0.007195f
C475 B.n268 VSUBS 0.007195f
C476 B.n269 VSUBS 0.007195f
C477 B.n270 VSUBS 0.007195f
C478 B.n271 VSUBS 0.007195f
C479 B.n272 VSUBS 0.007195f
C480 B.n273 VSUBS 0.007195f
C481 B.n274 VSUBS 0.007195f
C482 B.n275 VSUBS 0.007195f
C483 B.n276 VSUBS 0.007195f
C484 B.n277 VSUBS 0.007195f
C485 B.n278 VSUBS 0.007195f
C486 B.n279 VSUBS 0.007195f
C487 B.n280 VSUBS 0.007195f
C488 B.n281 VSUBS 0.007195f
C489 B.n282 VSUBS 0.007195f
C490 B.n283 VSUBS 0.007195f
C491 B.n284 VSUBS 0.007195f
C492 B.n285 VSUBS 0.007195f
C493 B.n286 VSUBS 0.007195f
C494 B.n287 VSUBS 0.007195f
C495 B.n288 VSUBS 0.007195f
C496 B.n289 VSUBS 0.007195f
C497 B.n290 VSUBS 0.007195f
C498 B.n291 VSUBS 0.007195f
C499 B.n292 VSUBS 0.007195f
C500 B.n293 VSUBS 0.007195f
C501 B.n294 VSUBS 0.007195f
C502 B.n295 VSUBS 0.007195f
C503 B.n296 VSUBS 0.007195f
C504 B.n297 VSUBS 0.007195f
C505 B.n298 VSUBS 0.007195f
C506 B.n299 VSUBS 0.007195f
C507 B.n300 VSUBS 0.007195f
C508 B.n301 VSUBS 0.007195f
C509 B.n302 VSUBS 0.007195f
C510 B.n303 VSUBS 0.007195f
C511 B.n304 VSUBS 0.007195f
C512 B.n305 VSUBS 0.007195f
C513 B.n306 VSUBS 0.007195f
C514 B.n307 VSUBS 0.007195f
C515 B.n308 VSUBS 0.007195f
C516 B.n309 VSUBS 0.007195f
C517 B.n310 VSUBS 0.007195f
C518 B.n311 VSUBS 0.007195f
C519 B.n312 VSUBS 0.007195f
C520 B.n313 VSUBS 0.007195f
C521 B.n314 VSUBS 0.007195f
C522 B.n315 VSUBS 0.007195f
C523 B.n316 VSUBS 0.007195f
C524 B.n317 VSUBS 0.007195f
C525 B.n318 VSUBS 0.007195f
C526 B.n319 VSUBS 0.007195f
C527 B.n320 VSUBS 0.007195f
C528 B.n321 VSUBS 0.007195f
C529 B.n322 VSUBS 0.007195f
C530 B.n323 VSUBS 0.007195f
C531 B.n324 VSUBS 0.007195f
C532 B.n325 VSUBS 0.007195f
C533 B.n326 VSUBS 0.007195f
C534 B.n327 VSUBS 0.007195f
C535 B.n328 VSUBS 0.018156f
C536 B.n329 VSUBS 0.01738f
C537 B.n330 VSUBS 0.018384f
C538 B.n331 VSUBS 0.007195f
C539 B.n332 VSUBS 0.007195f
C540 B.n333 VSUBS 0.007195f
C541 B.n334 VSUBS 0.007195f
C542 B.n335 VSUBS 0.007195f
C543 B.n336 VSUBS 0.007195f
C544 B.n337 VSUBS 0.007195f
C545 B.n338 VSUBS 0.007195f
C546 B.n339 VSUBS 0.007195f
C547 B.n340 VSUBS 0.007195f
C548 B.n341 VSUBS 0.007195f
C549 B.n342 VSUBS 0.007195f
C550 B.n343 VSUBS 0.007195f
C551 B.n344 VSUBS 0.007195f
C552 B.n345 VSUBS 0.007195f
C553 B.n346 VSUBS 0.007195f
C554 B.n347 VSUBS 0.007195f
C555 B.n348 VSUBS 0.007195f
C556 B.n349 VSUBS 0.007195f
C557 B.n350 VSUBS 0.007195f
C558 B.n351 VSUBS 0.007195f
C559 B.n352 VSUBS 0.007195f
C560 B.n353 VSUBS 0.007195f
C561 B.n354 VSUBS 0.007195f
C562 B.n355 VSUBS 0.007195f
C563 B.n356 VSUBS 0.007195f
C564 B.n357 VSUBS 0.007195f
C565 B.n358 VSUBS 0.007195f
C566 B.n359 VSUBS 0.007195f
C567 B.n360 VSUBS 0.007195f
C568 B.n361 VSUBS 0.007195f
C569 B.n362 VSUBS 0.007195f
C570 B.n363 VSUBS 0.007195f
C571 B.n364 VSUBS 0.007195f
C572 B.n365 VSUBS 0.007195f
C573 B.n366 VSUBS 0.007195f
C574 B.n367 VSUBS 0.007195f
C575 B.n368 VSUBS 0.007195f
C576 B.n369 VSUBS 0.007195f
C577 B.n370 VSUBS 0.017607f
C578 B.n371 VSUBS 0.017607f
C579 B.n372 VSUBS 0.018156f
C580 B.n373 VSUBS 0.007195f
C581 B.n374 VSUBS 0.007195f
C582 B.n375 VSUBS 0.007195f
C583 B.n376 VSUBS 0.007195f
C584 B.n377 VSUBS 0.007195f
C585 B.n378 VSUBS 0.007195f
C586 B.n379 VSUBS 0.007195f
C587 B.n380 VSUBS 0.007195f
C588 B.n381 VSUBS 0.007195f
C589 B.n382 VSUBS 0.007195f
C590 B.n383 VSUBS 0.007195f
C591 B.n384 VSUBS 0.007195f
C592 B.n385 VSUBS 0.007195f
C593 B.n386 VSUBS 0.007195f
C594 B.n387 VSUBS 0.007195f
C595 B.n388 VSUBS 0.007195f
C596 B.n389 VSUBS 0.007195f
C597 B.n390 VSUBS 0.007195f
C598 B.n391 VSUBS 0.007195f
C599 B.n392 VSUBS 0.007195f
C600 B.n393 VSUBS 0.007195f
C601 B.n394 VSUBS 0.007195f
C602 B.n395 VSUBS 0.007195f
C603 B.n396 VSUBS 0.007195f
C604 B.n397 VSUBS 0.007195f
C605 B.n398 VSUBS 0.007195f
C606 B.n399 VSUBS 0.007195f
C607 B.n400 VSUBS 0.007195f
C608 B.n401 VSUBS 0.007195f
C609 B.n402 VSUBS 0.007195f
C610 B.n403 VSUBS 0.007195f
C611 B.n404 VSUBS 0.007195f
C612 B.n405 VSUBS 0.007195f
C613 B.n406 VSUBS 0.007195f
C614 B.n407 VSUBS 0.007195f
C615 B.n408 VSUBS 0.007195f
C616 B.n409 VSUBS 0.007195f
C617 B.n410 VSUBS 0.007195f
C618 B.n411 VSUBS 0.007195f
C619 B.n412 VSUBS 0.007195f
C620 B.n413 VSUBS 0.007195f
C621 B.n414 VSUBS 0.007195f
C622 B.n415 VSUBS 0.007195f
C623 B.n416 VSUBS 0.007195f
C624 B.n417 VSUBS 0.007195f
C625 B.n418 VSUBS 0.007195f
C626 B.n419 VSUBS 0.007195f
C627 B.n420 VSUBS 0.007195f
C628 B.n421 VSUBS 0.007195f
C629 B.n422 VSUBS 0.007195f
C630 B.n423 VSUBS 0.007195f
C631 B.n424 VSUBS 0.007195f
C632 B.n425 VSUBS 0.007195f
C633 B.n426 VSUBS 0.007195f
C634 B.n427 VSUBS 0.007195f
C635 B.n428 VSUBS 0.007195f
C636 B.n429 VSUBS 0.007195f
C637 B.n430 VSUBS 0.007195f
C638 B.n431 VSUBS 0.007195f
C639 B.n432 VSUBS 0.007195f
C640 B.n433 VSUBS 0.007195f
C641 B.n434 VSUBS 0.007195f
C642 B.n435 VSUBS 0.007195f
C643 B.n436 VSUBS 0.007195f
C644 B.n437 VSUBS 0.007195f
C645 B.n438 VSUBS 0.007195f
C646 B.n439 VSUBS 0.007195f
C647 B.n440 VSUBS 0.007195f
C648 B.n441 VSUBS 0.007195f
C649 B.n442 VSUBS 0.007195f
C650 B.n443 VSUBS 0.007195f
C651 B.n444 VSUBS 0.007195f
C652 B.n445 VSUBS 0.004761f
C653 B.n446 VSUBS 0.007195f
C654 B.n447 VSUBS 0.007195f
C655 B.n448 VSUBS 0.006031f
C656 B.n449 VSUBS 0.007195f
C657 B.n450 VSUBS 0.007195f
C658 B.n451 VSUBS 0.007195f
C659 B.n452 VSUBS 0.007195f
C660 B.n453 VSUBS 0.007195f
C661 B.n454 VSUBS 0.007195f
C662 B.n455 VSUBS 0.007195f
C663 B.n456 VSUBS 0.007195f
C664 B.n457 VSUBS 0.007195f
C665 B.n458 VSUBS 0.007195f
C666 B.n459 VSUBS 0.007195f
C667 B.n460 VSUBS 0.006031f
C668 B.n461 VSUBS 0.01667f
C669 B.n462 VSUBS 0.004761f
C670 B.n463 VSUBS 0.007195f
C671 B.n464 VSUBS 0.007195f
C672 B.n465 VSUBS 0.007195f
C673 B.n466 VSUBS 0.007195f
C674 B.n467 VSUBS 0.007195f
C675 B.n468 VSUBS 0.007195f
C676 B.n469 VSUBS 0.007195f
C677 B.n470 VSUBS 0.007195f
C678 B.n471 VSUBS 0.007195f
C679 B.n472 VSUBS 0.007195f
C680 B.n473 VSUBS 0.007195f
C681 B.n474 VSUBS 0.007195f
C682 B.n475 VSUBS 0.007195f
C683 B.n476 VSUBS 0.007195f
C684 B.n477 VSUBS 0.007195f
C685 B.n478 VSUBS 0.007195f
C686 B.n479 VSUBS 0.007195f
C687 B.n480 VSUBS 0.007195f
C688 B.n481 VSUBS 0.007195f
C689 B.n482 VSUBS 0.007195f
C690 B.n483 VSUBS 0.007195f
C691 B.n484 VSUBS 0.007195f
C692 B.n485 VSUBS 0.007195f
C693 B.n486 VSUBS 0.007195f
C694 B.n487 VSUBS 0.007195f
C695 B.n488 VSUBS 0.007195f
C696 B.n489 VSUBS 0.007195f
C697 B.n490 VSUBS 0.007195f
C698 B.n491 VSUBS 0.007195f
C699 B.n492 VSUBS 0.007195f
C700 B.n493 VSUBS 0.007195f
C701 B.n494 VSUBS 0.007195f
C702 B.n495 VSUBS 0.007195f
C703 B.n496 VSUBS 0.007195f
C704 B.n497 VSUBS 0.007195f
C705 B.n498 VSUBS 0.007195f
C706 B.n499 VSUBS 0.007195f
C707 B.n500 VSUBS 0.007195f
C708 B.n501 VSUBS 0.007195f
C709 B.n502 VSUBS 0.007195f
C710 B.n503 VSUBS 0.007195f
C711 B.n504 VSUBS 0.007195f
C712 B.n505 VSUBS 0.007195f
C713 B.n506 VSUBS 0.007195f
C714 B.n507 VSUBS 0.007195f
C715 B.n508 VSUBS 0.007195f
C716 B.n509 VSUBS 0.007195f
C717 B.n510 VSUBS 0.007195f
C718 B.n511 VSUBS 0.007195f
C719 B.n512 VSUBS 0.007195f
C720 B.n513 VSUBS 0.007195f
C721 B.n514 VSUBS 0.007195f
C722 B.n515 VSUBS 0.007195f
C723 B.n516 VSUBS 0.007195f
C724 B.n517 VSUBS 0.007195f
C725 B.n518 VSUBS 0.007195f
C726 B.n519 VSUBS 0.007195f
C727 B.n520 VSUBS 0.007195f
C728 B.n521 VSUBS 0.007195f
C729 B.n522 VSUBS 0.007195f
C730 B.n523 VSUBS 0.007195f
C731 B.n524 VSUBS 0.007195f
C732 B.n525 VSUBS 0.007195f
C733 B.n526 VSUBS 0.007195f
C734 B.n527 VSUBS 0.007195f
C735 B.n528 VSUBS 0.007195f
C736 B.n529 VSUBS 0.007195f
C737 B.n530 VSUBS 0.007195f
C738 B.n531 VSUBS 0.007195f
C739 B.n532 VSUBS 0.007195f
C740 B.n533 VSUBS 0.007195f
C741 B.n534 VSUBS 0.007195f
C742 B.n535 VSUBS 0.018156f
C743 B.n536 VSUBS 0.018156f
C744 B.n537 VSUBS 0.017607f
C745 B.n538 VSUBS 0.007195f
C746 B.n539 VSUBS 0.007195f
C747 B.n540 VSUBS 0.007195f
C748 B.n541 VSUBS 0.007195f
C749 B.n542 VSUBS 0.007195f
C750 B.n543 VSUBS 0.007195f
C751 B.n544 VSUBS 0.007195f
C752 B.n545 VSUBS 0.007195f
C753 B.n546 VSUBS 0.007195f
C754 B.n547 VSUBS 0.007195f
C755 B.n548 VSUBS 0.007195f
C756 B.n549 VSUBS 0.007195f
C757 B.n550 VSUBS 0.007195f
C758 B.n551 VSUBS 0.007195f
C759 B.n552 VSUBS 0.007195f
C760 B.n553 VSUBS 0.007195f
C761 B.n554 VSUBS 0.007195f
C762 B.n555 VSUBS 0.009389f
C763 B.n556 VSUBS 0.010002f
C764 B.n557 VSUBS 0.019889f
C765 VDD2.n0 VSUBS 0.023134f
C766 VDD2.n1 VSUBS 0.021383f
C767 VDD2.n2 VSUBS 0.01149f
C768 VDD2.n3 VSUBS 0.027159f
C769 VDD2.n4 VSUBS 0.012166f
C770 VDD2.n5 VSUBS 0.021383f
C771 VDD2.n6 VSUBS 0.01149f
C772 VDD2.n7 VSUBS 0.027159f
C773 VDD2.n8 VSUBS 0.012166f
C774 VDD2.n9 VSUBS 0.021383f
C775 VDD2.n10 VSUBS 0.01149f
C776 VDD2.n11 VSUBS 0.027159f
C777 VDD2.n12 VSUBS 0.012166f
C778 VDD2.n13 VSUBS 0.021383f
C779 VDD2.n14 VSUBS 0.01149f
C780 VDD2.n15 VSUBS 0.027159f
C781 VDD2.n16 VSUBS 0.012166f
C782 VDD2.n17 VSUBS 0.021383f
C783 VDD2.n18 VSUBS 0.01149f
C784 VDD2.n19 VSUBS 0.027159f
C785 VDD2.n20 VSUBS 0.012166f
C786 VDD2.n21 VSUBS 0.021383f
C787 VDD2.n22 VSUBS 0.01149f
C788 VDD2.n23 VSUBS 0.027159f
C789 VDD2.n24 VSUBS 0.012166f
C790 VDD2.n25 VSUBS 0.149533f
C791 VDD2.t1 VSUBS 0.058132f
C792 VDD2.n26 VSUBS 0.020369f
C793 VDD2.n27 VSUBS 0.017277f
C794 VDD2.n28 VSUBS 0.01149f
C795 VDD2.n29 VSUBS 1.3469f
C796 VDD2.n30 VSUBS 0.021383f
C797 VDD2.n31 VSUBS 0.01149f
C798 VDD2.n32 VSUBS 0.012166f
C799 VDD2.n33 VSUBS 0.027159f
C800 VDD2.n34 VSUBS 0.027159f
C801 VDD2.n35 VSUBS 0.012166f
C802 VDD2.n36 VSUBS 0.01149f
C803 VDD2.n37 VSUBS 0.021383f
C804 VDD2.n38 VSUBS 0.021383f
C805 VDD2.n39 VSUBS 0.01149f
C806 VDD2.n40 VSUBS 0.012166f
C807 VDD2.n41 VSUBS 0.027159f
C808 VDD2.n42 VSUBS 0.027159f
C809 VDD2.n43 VSUBS 0.012166f
C810 VDD2.n44 VSUBS 0.01149f
C811 VDD2.n45 VSUBS 0.021383f
C812 VDD2.n46 VSUBS 0.021383f
C813 VDD2.n47 VSUBS 0.01149f
C814 VDD2.n48 VSUBS 0.012166f
C815 VDD2.n49 VSUBS 0.027159f
C816 VDD2.n50 VSUBS 0.027159f
C817 VDD2.n51 VSUBS 0.012166f
C818 VDD2.n52 VSUBS 0.01149f
C819 VDD2.n53 VSUBS 0.021383f
C820 VDD2.n54 VSUBS 0.021383f
C821 VDD2.n55 VSUBS 0.01149f
C822 VDD2.n56 VSUBS 0.012166f
C823 VDD2.n57 VSUBS 0.027159f
C824 VDD2.n58 VSUBS 0.027159f
C825 VDD2.n59 VSUBS 0.012166f
C826 VDD2.n60 VSUBS 0.01149f
C827 VDD2.n61 VSUBS 0.021383f
C828 VDD2.n62 VSUBS 0.021383f
C829 VDD2.n63 VSUBS 0.01149f
C830 VDD2.n64 VSUBS 0.012166f
C831 VDD2.n65 VSUBS 0.027159f
C832 VDD2.n66 VSUBS 0.027159f
C833 VDD2.n67 VSUBS 0.027159f
C834 VDD2.n68 VSUBS 0.012166f
C835 VDD2.n69 VSUBS 0.01149f
C836 VDD2.n70 VSUBS 0.021383f
C837 VDD2.n71 VSUBS 0.021383f
C838 VDD2.n72 VSUBS 0.01149f
C839 VDD2.n73 VSUBS 0.011828f
C840 VDD2.n74 VSUBS 0.011828f
C841 VDD2.n75 VSUBS 0.027159f
C842 VDD2.n76 VSUBS 0.064518f
C843 VDD2.n77 VSUBS 0.012166f
C844 VDD2.n78 VSUBS 0.01149f
C845 VDD2.n79 VSUBS 0.054392f
C846 VDD2.n80 VSUBS 0.583013f
C847 VDD2.n81 VSUBS 0.023134f
C848 VDD2.n82 VSUBS 0.021383f
C849 VDD2.n83 VSUBS 0.01149f
C850 VDD2.n84 VSUBS 0.027159f
C851 VDD2.n85 VSUBS 0.012166f
C852 VDD2.n86 VSUBS 0.021383f
C853 VDD2.n87 VSUBS 0.01149f
C854 VDD2.n88 VSUBS 0.027159f
C855 VDD2.n89 VSUBS 0.027159f
C856 VDD2.n90 VSUBS 0.012166f
C857 VDD2.n91 VSUBS 0.021383f
C858 VDD2.n92 VSUBS 0.01149f
C859 VDD2.n93 VSUBS 0.027159f
C860 VDD2.n94 VSUBS 0.012166f
C861 VDD2.n95 VSUBS 0.021383f
C862 VDD2.n96 VSUBS 0.01149f
C863 VDD2.n97 VSUBS 0.027159f
C864 VDD2.n98 VSUBS 0.012166f
C865 VDD2.n99 VSUBS 0.021383f
C866 VDD2.n100 VSUBS 0.01149f
C867 VDD2.n101 VSUBS 0.027159f
C868 VDD2.n102 VSUBS 0.012166f
C869 VDD2.n103 VSUBS 0.021383f
C870 VDD2.n104 VSUBS 0.01149f
C871 VDD2.n105 VSUBS 0.027159f
C872 VDD2.n106 VSUBS 0.012166f
C873 VDD2.n107 VSUBS 0.149533f
C874 VDD2.t0 VSUBS 0.058132f
C875 VDD2.n108 VSUBS 0.020369f
C876 VDD2.n109 VSUBS 0.017277f
C877 VDD2.n110 VSUBS 0.01149f
C878 VDD2.n111 VSUBS 1.3469f
C879 VDD2.n112 VSUBS 0.021383f
C880 VDD2.n113 VSUBS 0.01149f
C881 VDD2.n114 VSUBS 0.012166f
C882 VDD2.n115 VSUBS 0.027159f
C883 VDD2.n116 VSUBS 0.027159f
C884 VDD2.n117 VSUBS 0.012166f
C885 VDD2.n118 VSUBS 0.01149f
C886 VDD2.n119 VSUBS 0.021383f
C887 VDD2.n120 VSUBS 0.021383f
C888 VDD2.n121 VSUBS 0.01149f
C889 VDD2.n122 VSUBS 0.012166f
C890 VDD2.n123 VSUBS 0.027159f
C891 VDD2.n124 VSUBS 0.027159f
C892 VDD2.n125 VSUBS 0.012166f
C893 VDD2.n126 VSUBS 0.01149f
C894 VDD2.n127 VSUBS 0.021383f
C895 VDD2.n128 VSUBS 0.021383f
C896 VDD2.n129 VSUBS 0.01149f
C897 VDD2.n130 VSUBS 0.012166f
C898 VDD2.n131 VSUBS 0.027159f
C899 VDD2.n132 VSUBS 0.027159f
C900 VDD2.n133 VSUBS 0.012166f
C901 VDD2.n134 VSUBS 0.01149f
C902 VDD2.n135 VSUBS 0.021383f
C903 VDD2.n136 VSUBS 0.021383f
C904 VDD2.n137 VSUBS 0.01149f
C905 VDD2.n138 VSUBS 0.012166f
C906 VDD2.n139 VSUBS 0.027159f
C907 VDD2.n140 VSUBS 0.027159f
C908 VDD2.n141 VSUBS 0.012166f
C909 VDD2.n142 VSUBS 0.01149f
C910 VDD2.n143 VSUBS 0.021383f
C911 VDD2.n144 VSUBS 0.021383f
C912 VDD2.n145 VSUBS 0.01149f
C913 VDD2.n146 VSUBS 0.012166f
C914 VDD2.n147 VSUBS 0.027159f
C915 VDD2.n148 VSUBS 0.027159f
C916 VDD2.n149 VSUBS 0.012166f
C917 VDD2.n150 VSUBS 0.01149f
C918 VDD2.n151 VSUBS 0.021383f
C919 VDD2.n152 VSUBS 0.021383f
C920 VDD2.n153 VSUBS 0.01149f
C921 VDD2.n154 VSUBS 0.011828f
C922 VDD2.n155 VSUBS 0.011828f
C923 VDD2.n156 VSUBS 0.027159f
C924 VDD2.n157 VSUBS 0.064518f
C925 VDD2.n158 VSUBS 0.012166f
C926 VDD2.n159 VSUBS 0.01149f
C927 VDD2.n160 VSUBS 0.054392f
C928 VDD2.n161 VSUBS 0.047266f
C929 VDD2.n162 VSUBS 2.55283f
C930 VTAIL.n0 VSUBS 0.026926f
C931 VTAIL.n1 VSUBS 0.024888f
C932 VTAIL.n2 VSUBS 0.013374f
C933 VTAIL.n3 VSUBS 0.031611f
C934 VTAIL.n4 VSUBS 0.01416f
C935 VTAIL.n5 VSUBS 0.024888f
C936 VTAIL.n6 VSUBS 0.013374f
C937 VTAIL.n7 VSUBS 0.031611f
C938 VTAIL.n8 VSUBS 0.01416f
C939 VTAIL.n9 VSUBS 0.024888f
C940 VTAIL.n10 VSUBS 0.013374f
C941 VTAIL.n11 VSUBS 0.031611f
C942 VTAIL.n12 VSUBS 0.01416f
C943 VTAIL.n13 VSUBS 0.024888f
C944 VTAIL.n14 VSUBS 0.013374f
C945 VTAIL.n15 VSUBS 0.031611f
C946 VTAIL.n16 VSUBS 0.01416f
C947 VTAIL.n17 VSUBS 0.024888f
C948 VTAIL.n18 VSUBS 0.013374f
C949 VTAIL.n19 VSUBS 0.031611f
C950 VTAIL.n20 VSUBS 0.01416f
C951 VTAIL.n21 VSUBS 0.024888f
C952 VTAIL.n22 VSUBS 0.013374f
C953 VTAIL.n23 VSUBS 0.031611f
C954 VTAIL.n24 VSUBS 0.01416f
C955 VTAIL.n25 VSUBS 0.174046f
C956 VTAIL.t1 VSUBS 0.067661f
C957 VTAIL.n26 VSUBS 0.023708f
C958 VTAIL.n27 VSUBS 0.020109f
C959 VTAIL.n28 VSUBS 0.013374f
C960 VTAIL.n29 VSUBS 1.56769f
C961 VTAIL.n30 VSUBS 0.024888f
C962 VTAIL.n31 VSUBS 0.013374f
C963 VTAIL.n32 VSUBS 0.01416f
C964 VTAIL.n33 VSUBS 0.031611f
C965 VTAIL.n34 VSUBS 0.031611f
C966 VTAIL.n35 VSUBS 0.01416f
C967 VTAIL.n36 VSUBS 0.013374f
C968 VTAIL.n37 VSUBS 0.024888f
C969 VTAIL.n38 VSUBS 0.024888f
C970 VTAIL.n39 VSUBS 0.013374f
C971 VTAIL.n40 VSUBS 0.01416f
C972 VTAIL.n41 VSUBS 0.031611f
C973 VTAIL.n42 VSUBS 0.031611f
C974 VTAIL.n43 VSUBS 0.01416f
C975 VTAIL.n44 VSUBS 0.013374f
C976 VTAIL.n45 VSUBS 0.024888f
C977 VTAIL.n46 VSUBS 0.024888f
C978 VTAIL.n47 VSUBS 0.013374f
C979 VTAIL.n48 VSUBS 0.01416f
C980 VTAIL.n49 VSUBS 0.031611f
C981 VTAIL.n50 VSUBS 0.031611f
C982 VTAIL.n51 VSUBS 0.01416f
C983 VTAIL.n52 VSUBS 0.013374f
C984 VTAIL.n53 VSUBS 0.024888f
C985 VTAIL.n54 VSUBS 0.024888f
C986 VTAIL.n55 VSUBS 0.013374f
C987 VTAIL.n56 VSUBS 0.01416f
C988 VTAIL.n57 VSUBS 0.031611f
C989 VTAIL.n58 VSUBS 0.031611f
C990 VTAIL.n59 VSUBS 0.01416f
C991 VTAIL.n60 VSUBS 0.013374f
C992 VTAIL.n61 VSUBS 0.024888f
C993 VTAIL.n62 VSUBS 0.024888f
C994 VTAIL.n63 VSUBS 0.013374f
C995 VTAIL.n64 VSUBS 0.01416f
C996 VTAIL.n65 VSUBS 0.031611f
C997 VTAIL.n66 VSUBS 0.031611f
C998 VTAIL.n67 VSUBS 0.031611f
C999 VTAIL.n68 VSUBS 0.01416f
C1000 VTAIL.n69 VSUBS 0.013374f
C1001 VTAIL.n70 VSUBS 0.024888f
C1002 VTAIL.n71 VSUBS 0.024888f
C1003 VTAIL.n72 VSUBS 0.013374f
C1004 VTAIL.n73 VSUBS 0.013767f
C1005 VTAIL.n74 VSUBS 0.013767f
C1006 VTAIL.n75 VSUBS 0.031611f
C1007 VTAIL.n76 VSUBS 0.075094f
C1008 VTAIL.n77 VSUBS 0.01416f
C1009 VTAIL.n78 VSUBS 0.013374f
C1010 VTAIL.n79 VSUBS 0.063308f
C1011 VTAIL.n80 VSUBS 0.037871f
C1012 VTAIL.n81 VSUBS 1.57486f
C1013 VTAIL.n82 VSUBS 0.026926f
C1014 VTAIL.n83 VSUBS 0.024888f
C1015 VTAIL.n84 VSUBS 0.013374f
C1016 VTAIL.n85 VSUBS 0.031611f
C1017 VTAIL.n86 VSUBS 0.01416f
C1018 VTAIL.n87 VSUBS 0.024888f
C1019 VTAIL.n88 VSUBS 0.013374f
C1020 VTAIL.n89 VSUBS 0.031611f
C1021 VTAIL.n90 VSUBS 0.031611f
C1022 VTAIL.n91 VSUBS 0.01416f
C1023 VTAIL.n92 VSUBS 0.024888f
C1024 VTAIL.n93 VSUBS 0.013374f
C1025 VTAIL.n94 VSUBS 0.031611f
C1026 VTAIL.n95 VSUBS 0.01416f
C1027 VTAIL.n96 VSUBS 0.024888f
C1028 VTAIL.n97 VSUBS 0.013374f
C1029 VTAIL.n98 VSUBS 0.031611f
C1030 VTAIL.n99 VSUBS 0.01416f
C1031 VTAIL.n100 VSUBS 0.024888f
C1032 VTAIL.n101 VSUBS 0.013374f
C1033 VTAIL.n102 VSUBS 0.031611f
C1034 VTAIL.n103 VSUBS 0.01416f
C1035 VTAIL.n104 VSUBS 0.024888f
C1036 VTAIL.n105 VSUBS 0.013374f
C1037 VTAIL.n106 VSUBS 0.031611f
C1038 VTAIL.n107 VSUBS 0.01416f
C1039 VTAIL.n108 VSUBS 0.174046f
C1040 VTAIL.t3 VSUBS 0.067661f
C1041 VTAIL.n109 VSUBS 0.023708f
C1042 VTAIL.n110 VSUBS 0.020109f
C1043 VTAIL.n111 VSUBS 0.013374f
C1044 VTAIL.n112 VSUBS 1.56769f
C1045 VTAIL.n113 VSUBS 0.024888f
C1046 VTAIL.n114 VSUBS 0.013374f
C1047 VTAIL.n115 VSUBS 0.01416f
C1048 VTAIL.n116 VSUBS 0.031611f
C1049 VTAIL.n117 VSUBS 0.031611f
C1050 VTAIL.n118 VSUBS 0.01416f
C1051 VTAIL.n119 VSUBS 0.013374f
C1052 VTAIL.n120 VSUBS 0.024888f
C1053 VTAIL.n121 VSUBS 0.024888f
C1054 VTAIL.n122 VSUBS 0.013374f
C1055 VTAIL.n123 VSUBS 0.01416f
C1056 VTAIL.n124 VSUBS 0.031611f
C1057 VTAIL.n125 VSUBS 0.031611f
C1058 VTAIL.n126 VSUBS 0.01416f
C1059 VTAIL.n127 VSUBS 0.013374f
C1060 VTAIL.n128 VSUBS 0.024888f
C1061 VTAIL.n129 VSUBS 0.024888f
C1062 VTAIL.n130 VSUBS 0.013374f
C1063 VTAIL.n131 VSUBS 0.01416f
C1064 VTAIL.n132 VSUBS 0.031611f
C1065 VTAIL.n133 VSUBS 0.031611f
C1066 VTAIL.n134 VSUBS 0.01416f
C1067 VTAIL.n135 VSUBS 0.013374f
C1068 VTAIL.n136 VSUBS 0.024888f
C1069 VTAIL.n137 VSUBS 0.024888f
C1070 VTAIL.n138 VSUBS 0.013374f
C1071 VTAIL.n139 VSUBS 0.01416f
C1072 VTAIL.n140 VSUBS 0.031611f
C1073 VTAIL.n141 VSUBS 0.031611f
C1074 VTAIL.n142 VSUBS 0.01416f
C1075 VTAIL.n143 VSUBS 0.013374f
C1076 VTAIL.n144 VSUBS 0.024888f
C1077 VTAIL.n145 VSUBS 0.024888f
C1078 VTAIL.n146 VSUBS 0.013374f
C1079 VTAIL.n147 VSUBS 0.01416f
C1080 VTAIL.n148 VSUBS 0.031611f
C1081 VTAIL.n149 VSUBS 0.031611f
C1082 VTAIL.n150 VSUBS 0.01416f
C1083 VTAIL.n151 VSUBS 0.013374f
C1084 VTAIL.n152 VSUBS 0.024888f
C1085 VTAIL.n153 VSUBS 0.024888f
C1086 VTAIL.n154 VSUBS 0.013374f
C1087 VTAIL.n155 VSUBS 0.013767f
C1088 VTAIL.n156 VSUBS 0.013767f
C1089 VTAIL.n157 VSUBS 0.031611f
C1090 VTAIL.n158 VSUBS 0.075094f
C1091 VTAIL.n159 VSUBS 0.01416f
C1092 VTAIL.n160 VSUBS 0.013374f
C1093 VTAIL.n161 VSUBS 0.063308f
C1094 VTAIL.n162 VSUBS 0.037871f
C1095 VTAIL.n163 VSUBS 1.58627f
C1096 VTAIL.n164 VSUBS 0.026926f
C1097 VTAIL.n165 VSUBS 0.024888f
C1098 VTAIL.n166 VSUBS 0.013374f
C1099 VTAIL.n167 VSUBS 0.031611f
C1100 VTAIL.n168 VSUBS 0.01416f
C1101 VTAIL.n169 VSUBS 0.024888f
C1102 VTAIL.n170 VSUBS 0.013374f
C1103 VTAIL.n171 VSUBS 0.031611f
C1104 VTAIL.n172 VSUBS 0.031611f
C1105 VTAIL.n173 VSUBS 0.01416f
C1106 VTAIL.n174 VSUBS 0.024888f
C1107 VTAIL.n175 VSUBS 0.013374f
C1108 VTAIL.n176 VSUBS 0.031611f
C1109 VTAIL.n177 VSUBS 0.01416f
C1110 VTAIL.n178 VSUBS 0.024888f
C1111 VTAIL.n179 VSUBS 0.013374f
C1112 VTAIL.n180 VSUBS 0.031611f
C1113 VTAIL.n181 VSUBS 0.01416f
C1114 VTAIL.n182 VSUBS 0.024888f
C1115 VTAIL.n183 VSUBS 0.013374f
C1116 VTAIL.n184 VSUBS 0.031611f
C1117 VTAIL.n185 VSUBS 0.01416f
C1118 VTAIL.n186 VSUBS 0.024888f
C1119 VTAIL.n187 VSUBS 0.013374f
C1120 VTAIL.n188 VSUBS 0.031611f
C1121 VTAIL.n189 VSUBS 0.01416f
C1122 VTAIL.n190 VSUBS 0.174046f
C1123 VTAIL.t0 VSUBS 0.067661f
C1124 VTAIL.n191 VSUBS 0.023708f
C1125 VTAIL.n192 VSUBS 0.020109f
C1126 VTAIL.n193 VSUBS 0.013374f
C1127 VTAIL.n194 VSUBS 1.56769f
C1128 VTAIL.n195 VSUBS 0.024888f
C1129 VTAIL.n196 VSUBS 0.013374f
C1130 VTAIL.n197 VSUBS 0.01416f
C1131 VTAIL.n198 VSUBS 0.031611f
C1132 VTAIL.n199 VSUBS 0.031611f
C1133 VTAIL.n200 VSUBS 0.01416f
C1134 VTAIL.n201 VSUBS 0.013374f
C1135 VTAIL.n202 VSUBS 0.024888f
C1136 VTAIL.n203 VSUBS 0.024888f
C1137 VTAIL.n204 VSUBS 0.013374f
C1138 VTAIL.n205 VSUBS 0.01416f
C1139 VTAIL.n206 VSUBS 0.031611f
C1140 VTAIL.n207 VSUBS 0.031611f
C1141 VTAIL.n208 VSUBS 0.01416f
C1142 VTAIL.n209 VSUBS 0.013374f
C1143 VTAIL.n210 VSUBS 0.024888f
C1144 VTAIL.n211 VSUBS 0.024888f
C1145 VTAIL.n212 VSUBS 0.013374f
C1146 VTAIL.n213 VSUBS 0.01416f
C1147 VTAIL.n214 VSUBS 0.031611f
C1148 VTAIL.n215 VSUBS 0.031611f
C1149 VTAIL.n216 VSUBS 0.01416f
C1150 VTAIL.n217 VSUBS 0.013374f
C1151 VTAIL.n218 VSUBS 0.024888f
C1152 VTAIL.n219 VSUBS 0.024888f
C1153 VTAIL.n220 VSUBS 0.013374f
C1154 VTAIL.n221 VSUBS 0.01416f
C1155 VTAIL.n222 VSUBS 0.031611f
C1156 VTAIL.n223 VSUBS 0.031611f
C1157 VTAIL.n224 VSUBS 0.01416f
C1158 VTAIL.n225 VSUBS 0.013374f
C1159 VTAIL.n226 VSUBS 0.024888f
C1160 VTAIL.n227 VSUBS 0.024888f
C1161 VTAIL.n228 VSUBS 0.013374f
C1162 VTAIL.n229 VSUBS 0.01416f
C1163 VTAIL.n230 VSUBS 0.031611f
C1164 VTAIL.n231 VSUBS 0.031611f
C1165 VTAIL.n232 VSUBS 0.01416f
C1166 VTAIL.n233 VSUBS 0.013374f
C1167 VTAIL.n234 VSUBS 0.024888f
C1168 VTAIL.n235 VSUBS 0.024888f
C1169 VTAIL.n236 VSUBS 0.013374f
C1170 VTAIL.n237 VSUBS 0.013767f
C1171 VTAIL.n238 VSUBS 0.013767f
C1172 VTAIL.n239 VSUBS 0.031611f
C1173 VTAIL.n240 VSUBS 0.075094f
C1174 VTAIL.n241 VSUBS 0.01416f
C1175 VTAIL.n242 VSUBS 0.013374f
C1176 VTAIL.n243 VSUBS 0.063308f
C1177 VTAIL.n244 VSUBS 0.037871f
C1178 VTAIL.n245 VSUBS 1.52198f
C1179 VTAIL.n246 VSUBS 0.026926f
C1180 VTAIL.n247 VSUBS 0.024888f
C1181 VTAIL.n248 VSUBS 0.013374f
C1182 VTAIL.n249 VSUBS 0.031611f
C1183 VTAIL.n250 VSUBS 0.01416f
C1184 VTAIL.n251 VSUBS 0.024888f
C1185 VTAIL.n252 VSUBS 0.013374f
C1186 VTAIL.n253 VSUBS 0.031611f
C1187 VTAIL.n254 VSUBS 0.01416f
C1188 VTAIL.n255 VSUBS 0.024888f
C1189 VTAIL.n256 VSUBS 0.013374f
C1190 VTAIL.n257 VSUBS 0.031611f
C1191 VTAIL.n258 VSUBS 0.01416f
C1192 VTAIL.n259 VSUBS 0.024888f
C1193 VTAIL.n260 VSUBS 0.013374f
C1194 VTAIL.n261 VSUBS 0.031611f
C1195 VTAIL.n262 VSUBS 0.01416f
C1196 VTAIL.n263 VSUBS 0.024888f
C1197 VTAIL.n264 VSUBS 0.013374f
C1198 VTAIL.n265 VSUBS 0.031611f
C1199 VTAIL.n266 VSUBS 0.01416f
C1200 VTAIL.n267 VSUBS 0.024888f
C1201 VTAIL.n268 VSUBS 0.013374f
C1202 VTAIL.n269 VSUBS 0.031611f
C1203 VTAIL.n270 VSUBS 0.01416f
C1204 VTAIL.n271 VSUBS 0.174046f
C1205 VTAIL.t2 VSUBS 0.067661f
C1206 VTAIL.n272 VSUBS 0.023708f
C1207 VTAIL.n273 VSUBS 0.020109f
C1208 VTAIL.n274 VSUBS 0.013374f
C1209 VTAIL.n275 VSUBS 1.56769f
C1210 VTAIL.n276 VSUBS 0.024888f
C1211 VTAIL.n277 VSUBS 0.013374f
C1212 VTAIL.n278 VSUBS 0.01416f
C1213 VTAIL.n279 VSUBS 0.031611f
C1214 VTAIL.n280 VSUBS 0.031611f
C1215 VTAIL.n281 VSUBS 0.01416f
C1216 VTAIL.n282 VSUBS 0.013374f
C1217 VTAIL.n283 VSUBS 0.024888f
C1218 VTAIL.n284 VSUBS 0.024888f
C1219 VTAIL.n285 VSUBS 0.013374f
C1220 VTAIL.n286 VSUBS 0.01416f
C1221 VTAIL.n287 VSUBS 0.031611f
C1222 VTAIL.n288 VSUBS 0.031611f
C1223 VTAIL.n289 VSUBS 0.01416f
C1224 VTAIL.n290 VSUBS 0.013374f
C1225 VTAIL.n291 VSUBS 0.024888f
C1226 VTAIL.n292 VSUBS 0.024888f
C1227 VTAIL.n293 VSUBS 0.013374f
C1228 VTAIL.n294 VSUBS 0.01416f
C1229 VTAIL.n295 VSUBS 0.031611f
C1230 VTAIL.n296 VSUBS 0.031611f
C1231 VTAIL.n297 VSUBS 0.01416f
C1232 VTAIL.n298 VSUBS 0.013374f
C1233 VTAIL.n299 VSUBS 0.024888f
C1234 VTAIL.n300 VSUBS 0.024888f
C1235 VTAIL.n301 VSUBS 0.013374f
C1236 VTAIL.n302 VSUBS 0.01416f
C1237 VTAIL.n303 VSUBS 0.031611f
C1238 VTAIL.n304 VSUBS 0.031611f
C1239 VTAIL.n305 VSUBS 0.01416f
C1240 VTAIL.n306 VSUBS 0.013374f
C1241 VTAIL.n307 VSUBS 0.024888f
C1242 VTAIL.n308 VSUBS 0.024888f
C1243 VTAIL.n309 VSUBS 0.013374f
C1244 VTAIL.n310 VSUBS 0.01416f
C1245 VTAIL.n311 VSUBS 0.031611f
C1246 VTAIL.n312 VSUBS 0.031611f
C1247 VTAIL.n313 VSUBS 0.031611f
C1248 VTAIL.n314 VSUBS 0.01416f
C1249 VTAIL.n315 VSUBS 0.013374f
C1250 VTAIL.n316 VSUBS 0.024888f
C1251 VTAIL.n317 VSUBS 0.024888f
C1252 VTAIL.n318 VSUBS 0.013374f
C1253 VTAIL.n319 VSUBS 0.013767f
C1254 VTAIL.n320 VSUBS 0.013767f
C1255 VTAIL.n321 VSUBS 0.031611f
C1256 VTAIL.n322 VSUBS 0.075094f
C1257 VTAIL.n323 VSUBS 0.01416f
C1258 VTAIL.n324 VSUBS 0.013374f
C1259 VTAIL.n325 VSUBS 0.063308f
C1260 VTAIL.n326 VSUBS 0.037871f
C1261 VTAIL.n327 VSUBS 1.46356f
C1262 VN.t0 VSUBS 1.29489f
C1263 VN.t1 VSUBS 1.4079f
.ends

