* NGSPICE file created from diff_pair_sample_0512.ext - technology: sky130A

.subckt diff_pair_sample_0512 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=0 ps=0 w=13.66 l=2.35
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=0 ps=0 w=13.66 l=2.35
X2 VDD2.t3 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2539 pd=13.99 as=5.3274 ps=28.1 w=13.66 l=2.35
X3 VTAIL.t4 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=2.2539 ps=13.99 w=13.66 l=2.35
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=0 ps=0 w=13.66 l=2.35
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=0 ps=0 w=13.66 l=2.35
X6 VTAIL.t5 VN.t2 VDD2.t1 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=2.2539 ps=13.99 w=13.66 l=2.35
X7 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2539 pd=13.99 as=5.3274 ps=28.1 w=13.66 l=2.35
X8 VDD1.t2 VP.t1 VTAIL.t3 B.t17 sky130_fd_pr__nfet_01v8 ad=2.2539 pd=13.99 as=5.3274 ps=28.1 w=13.66 l=2.35
X9 VTAIL.t2 VP.t2 VDD1.t1 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=2.2539 ps=13.99 w=13.66 l=2.35
X10 VDD2.t0 VN.t3 VTAIL.t7 B.t17 sky130_fd_pr__nfet_01v8 ad=2.2539 pd=13.99 as=5.3274 ps=28.1 w=13.66 l=2.35
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3274 pd=28.1 as=2.2539 ps=13.99 w=13.66 l=2.35
R0 B.n777 B.n776 585
R1 B.n778 B.n777 585
R2 B.n318 B.n112 585
R3 B.n317 B.n316 585
R4 B.n315 B.n314 585
R5 B.n313 B.n312 585
R6 B.n311 B.n310 585
R7 B.n309 B.n308 585
R8 B.n307 B.n306 585
R9 B.n305 B.n304 585
R10 B.n303 B.n302 585
R11 B.n301 B.n300 585
R12 B.n299 B.n298 585
R13 B.n297 B.n296 585
R14 B.n295 B.n294 585
R15 B.n293 B.n292 585
R16 B.n291 B.n290 585
R17 B.n289 B.n288 585
R18 B.n287 B.n286 585
R19 B.n285 B.n284 585
R20 B.n283 B.n282 585
R21 B.n281 B.n280 585
R22 B.n279 B.n278 585
R23 B.n277 B.n276 585
R24 B.n275 B.n274 585
R25 B.n273 B.n272 585
R26 B.n271 B.n270 585
R27 B.n269 B.n268 585
R28 B.n267 B.n266 585
R29 B.n265 B.n264 585
R30 B.n263 B.n262 585
R31 B.n261 B.n260 585
R32 B.n259 B.n258 585
R33 B.n257 B.n256 585
R34 B.n255 B.n254 585
R35 B.n253 B.n252 585
R36 B.n251 B.n250 585
R37 B.n249 B.n248 585
R38 B.n247 B.n246 585
R39 B.n245 B.n244 585
R40 B.n243 B.n242 585
R41 B.n241 B.n240 585
R42 B.n239 B.n238 585
R43 B.n237 B.n236 585
R44 B.n235 B.n234 585
R45 B.n233 B.n232 585
R46 B.n231 B.n230 585
R47 B.n229 B.n228 585
R48 B.n227 B.n226 585
R49 B.n225 B.n224 585
R50 B.n223 B.n222 585
R51 B.n221 B.n220 585
R52 B.n219 B.n218 585
R53 B.n217 B.n216 585
R54 B.n215 B.n214 585
R55 B.n213 B.n212 585
R56 B.n211 B.n210 585
R57 B.n208 B.n207 585
R58 B.n206 B.n205 585
R59 B.n204 B.n203 585
R60 B.n202 B.n201 585
R61 B.n200 B.n199 585
R62 B.n198 B.n197 585
R63 B.n196 B.n195 585
R64 B.n194 B.n193 585
R65 B.n192 B.n191 585
R66 B.n190 B.n189 585
R67 B.n188 B.n187 585
R68 B.n186 B.n185 585
R69 B.n184 B.n183 585
R70 B.n182 B.n181 585
R71 B.n180 B.n179 585
R72 B.n178 B.n177 585
R73 B.n176 B.n175 585
R74 B.n174 B.n173 585
R75 B.n172 B.n171 585
R76 B.n170 B.n169 585
R77 B.n168 B.n167 585
R78 B.n166 B.n165 585
R79 B.n164 B.n163 585
R80 B.n162 B.n161 585
R81 B.n160 B.n159 585
R82 B.n158 B.n157 585
R83 B.n156 B.n155 585
R84 B.n154 B.n153 585
R85 B.n152 B.n151 585
R86 B.n150 B.n149 585
R87 B.n148 B.n147 585
R88 B.n146 B.n145 585
R89 B.n144 B.n143 585
R90 B.n142 B.n141 585
R91 B.n140 B.n139 585
R92 B.n138 B.n137 585
R93 B.n136 B.n135 585
R94 B.n134 B.n133 585
R95 B.n132 B.n131 585
R96 B.n130 B.n129 585
R97 B.n128 B.n127 585
R98 B.n126 B.n125 585
R99 B.n124 B.n123 585
R100 B.n122 B.n121 585
R101 B.n120 B.n119 585
R102 B.n61 B.n60 585
R103 B.n781 B.n780 585
R104 B.n775 B.n113 585
R105 B.n113 B.n58 585
R106 B.n774 B.n57 585
R107 B.n785 B.n57 585
R108 B.n773 B.n56 585
R109 B.n786 B.n56 585
R110 B.n772 B.n55 585
R111 B.n787 B.n55 585
R112 B.n771 B.n770 585
R113 B.n770 B.n51 585
R114 B.n769 B.n50 585
R115 B.n793 B.n50 585
R116 B.n768 B.n49 585
R117 B.n794 B.n49 585
R118 B.n767 B.n48 585
R119 B.n795 B.n48 585
R120 B.n766 B.n765 585
R121 B.n765 B.n44 585
R122 B.n764 B.n43 585
R123 B.n801 B.n43 585
R124 B.n763 B.n42 585
R125 B.n802 B.n42 585
R126 B.n762 B.n41 585
R127 B.n803 B.n41 585
R128 B.n761 B.n760 585
R129 B.n760 B.n37 585
R130 B.n759 B.n36 585
R131 B.n809 B.n36 585
R132 B.n758 B.n35 585
R133 B.n810 B.n35 585
R134 B.n757 B.n34 585
R135 B.n811 B.n34 585
R136 B.n756 B.n755 585
R137 B.n755 B.n30 585
R138 B.n754 B.n29 585
R139 B.n817 B.n29 585
R140 B.n753 B.n28 585
R141 B.n818 B.n28 585
R142 B.n752 B.n27 585
R143 B.n819 B.n27 585
R144 B.n751 B.n750 585
R145 B.n750 B.n23 585
R146 B.n749 B.n22 585
R147 B.n825 B.n22 585
R148 B.n748 B.n21 585
R149 B.n826 B.n21 585
R150 B.n747 B.n20 585
R151 B.n827 B.n20 585
R152 B.n746 B.n745 585
R153 B.n745 B.n16 585
R154 B.n744 B.n15 585
R155 B.n833 B.n15 585
R156 B.n743 B.n14 585
R157 B.n834 B.n14 585
R158 B.n742 B.n13 585
R159 B.n835 B.n13 585
R160 B.n741 B.n740 585
R161 B.n740 B.n12 585
R162 B.n739 B.n738 585
R163 B.n739 B.n8 585
R164 B.n737 B.n7 585
R165 B.n842 B.n7 585
R166 B.n736 B.n6 585
R167 B.n843 B.n6 585
R168 B.n735 B.n5 585
R169 B.n844 B.n5 585
R170 B.n734 B.n733 585
R171 B.n733 B.n4 585
R172 B.n732 B.n319 585
R173 B.n732 B.n731 585
R174 B.n722 B.n320 585
R175 B.n321 B.n320 585
R176 B.n724 B.n723 585
R177 B.n725 B.n724 585
R178 B.n721 B.n326 585
R179 B.n326 B.n325 585
R180 B.n720 B.n719 585
R181 B.n719 B.n718 585
R182 B.n328 B.n327 585
R183 B.n329 B.n328 585
R184 B.n711 B.n710 585
R185 B.n712 B.n711 585
R186 B.n709 B.n334 585
R187 B.n334 B.n333 585
R188 B.n708 B.n707 585
R189 B.n707 B.n706 585
R190 B.n336 B.n335 585
R191 B.n337 B.n336 585
R192 B.n699 B.n698 585
R193 B.n700 B.n699 585
R194 B.n697 B.n341 585
R195 B.n345 B.n341 585
R196 B.n696 B.n695 585
R197 B.n695 B.n694 585
R198 B.n343 B.n342 585
R199 B.n344 B.n343 585
R200 B.n687 B.n686 585
R201 B.n688 B.n687 585
R202 B.n685 B.n350 585
R203 B.n350 B.n349 585
R204 B.n684 B.n683 585
R205 B.n683 B.n682 585
R206 B.n352 B.n351 585
R207 B.n353 B.n352 585
R208 B.n675 B.n674 585
R209 B.n676 B.n675 585
R210 B.n673 B.n358 585
R211 B.n358 B.n357 585
R212 B.n672 B.n671 585
R213 B.n671 B.n670 585
R214 B.n360 B.n359 585
R215 B.n361 B.n360 585
R216 B.n663 B.n662 585
R217 B.n664 B.n663 585
R218 B.n661 B.n365 585
R219 B.n369 B.n365 585
R220 B.n660 B.n659 585
R221 B.n659 B.n658 585
R222 B.n367 B.n366 585
R223 B.n368 B.n367 585
R224 B.n651 B.n650 585
R225 B.n652 B.n651 585
R226 B.n649 B.n374 585
R227 B.n374 B.n373 585
R228 B.n648 B.n647 585
R229 B.n647 B.n646 585
R230 B.n376 B.n375 585
R231 B.n377 B.n376 585
R232 B.n642 B.n641 585
R233 B.n380 B.n379 585
R234 B.n638 B.n637 585
R235 B.n639 B.n638 585
R236 B.n636 B.n431 585
R237 B.n635 B.n634 585
R238 B.n633 B.n632 585
R239 B.n631 B.n630 585
R240 B.n629 B.n628 585
R241 B.n627 B.n626 585
R242 B.n625 B.n624 585
R243 B.n623 B.n622 585
R244 B.n621 B.n620 585
R245 B.n619 B.n618 585
R246 B.n617 B.n616 585
R247 B.n615 B.n614 585
R248 B.n613 B.n612 585
R249 B.n611 B.n610 585
R250 B.n609 B.n608 585
R251 B.n607 B.n606 585
R252 B.n605 B.n604 585
R253 B.n603 B.n602 585
R254 B.n601 B.n600 585
R255 B.n599 B.n598 585
R256 B.n597 B.n596 585
R257 B.n595 B.n594 585
R258 B.n593 B.n592 585
R259 B.n591 B.n590 585
R260 B.n589 B.n588 585
R261 B.n587 B.n586 585
R262 B.n585 B.n584 585
R263 B.n583 B.n582 585
R264 B.n581 B.n580 585
R265 B.n579 B.n578 585
R266 B.n577 B.n576 585
R267 B.n575 B.n574 585
R268 B.n573 B.n572 585
R269 B.n571 B.n570 585
R270 B.n569 B.n568 585
R271 B.n567 B.n566 585
R272 B.n565 B.n564 585
R273 B.n563 B.n562 585
R274 B.n561 B.n560 585
R275 B.n559 B.n558 585
R276 B.n557 B.n556 585
R277 B.n555 B.n554 585
R278 B.n553 B.n552 585
R279 B.n551 B.n550 585
R280 B.n549 B.n548 585
R281 B.n547 B.n546 585
R282 B.n545 B.n544 585
R283 B.n543 B.n542 585
R284 B.n541 B.n540 585
R285 B.n539 B.n538 585
R286 B.n537 B.n536 585
R287 B.n535 B.n534 585
R288 B.n533 B.n532 585
R289 B.n530 B.n529 585
R290 B.n528 B.n527 585
R291 B.n526 B.n525 585
R292 B.n524 B.n523 585
R293 B.n522 B.n521 585
R294 B.n520 B.n519 585
R295 B.n518 B.n517 585
R296 B.n516 B.n515 585
R297 B.n514 B.n513 585
R298 B.n512 B.n511 585
R299 B.n510 B.n509 585
R300 B.n508 B.n507 585
R301 B.n506 B.n505 585
R302 B.n504 B.n503 585
R303 B.n502 B.n501 585
R304 B.n500 B.n499 585
R305 B.n498 B.n497 585
R306 B.n496 B.n495 585
R307 B.n494 B.n493 585
R308 B.n492 B.n491 585
R309 B.n490 B.n489 585
R310 B.n488 B.n487 585
R311 B.n486 B.n485 585
R312 B.n484 B.n483 585
R313 B.n482 B.n481 585
R314 B.n480 B.n479 585
R315 B.n478 B.n477 585
R316 B.n476 B.n475 585
R317 B.n474 B.n473 585
R318 B.n472 B.n471 585
R319 B.n470 B.n469 585
R320 B.n468 B.n467 585
R321 B.n466 B.n465 585
R322 B.n464 B.n463 585
R323 B.n462 B.n461 585
R324 B.n460 B.n459 585
R325 B.n458 B.n457 585
R326 B.n456 B.n455 585
R327 B.n454 B.n453 585
R328 B.n452 B.n451 585
R329 B.n450 B.n449 585
R330 B.n448 B.n447 585
R331 B.n446 B.n445 585
R332 B.n444 B.n443 585
R333 B.n442 B.n441 585
R334 B.n440 B.n439 585
R335 B.n438 B.n437 585
R336 B.n643 B.n378 585
R337 B.n378 B.n377 585
R338 B.n645 B.n644 585
R339 B.n646 B.n645 585
R340 B.n372 B.n371 585
R341 B.n373 B.n372 585
R342 B.n654 B.n653 585
R343 B.n653 B.n652 585
R344 B.n655 B.n370 585
R345 B.n370 B.n368 585
R346 B.n657 B.n656 585
R347 B.n658 B.n657 585
R348 B.n364 B.n363 585
R349 B.n369 B.n364 585
R350 B.n666 B.n665 585
R351 B.n665 B.n664 585
R352 B.n667 B.n362 585
R353 B.n362 B.n361 585
R354 B.n669 B.n668 585
R355 B.n670 B.n669 585
R356 B.n356 B.n355 585
R357 B.n357 B.n356 585
R358 B.n678 B.n677 585
R359 B.n677 B.n676 585
R360 B.n679 B.n354 585
R361 B.n354 B.n353 585
R362 B.n681 B.n680 585
R363 B.n682 B.n681 585
R364 B.n348 B.n347 585
R365 B.n349 B.n348 585
R366 B.n690 B.n689 585
R367 B.n689 B.n688 585
R368 B.n691 B.n346 585
R369 B.n346 B.n344 585
R370 B.n693 B.n692 585
R371 B.n694 B.n693 585
R372 B.n340 B.n339 585
R373 B.n345 B.n340 585
R374 B.n702 B.n701 585
R375 B.n701 B.n700 585
R376 B.n703 B.n338 585
R377 B.n338 B.n337 585
R378 B.n705 B.n704 585
R379 B.n706 B.n705 585
R380 B.n332 B.n331 585
R381 B.n333 B.n332 585
R382 B.n714 B.n713 585
R383 B.n713 B.n712 585
R384 B.n715 B.n330 585
R385 B.n330 B.n329 585
R386 B.n717 B.n716 585
R387 B.n718 B.n717 585
R388 B.n324 B.n323 585
R389 B.n325 B.n324 585
R390 B.n727 B.n726 585
R391 B.n726 B.n725 585
R392 B.n728 B.n322 585
R393 B.n322 B.n321 585
R394 B.n730 B.n729 585
R395 B.n731 B.n730 585
R396 B.n3 B.n0 585
R397 B.n4 B.n3 585
R398 B.n841 B.n1 585
R399 B.n842 B.n841 585
R400 B.n840 B.n839 585
R401 B.n840 B.n8 585
R402 B.n838 B.n9 585
R403 B.n12 B.n9 585
R404 B.n837 B.n836 585
R405 B.n836 B.n835 585
R406 B.n11 B.n10 585
R407 B.n834 B.n11 585
R408 B.n832 B.n831 585
R409 B.n833 B.n832 585
R410 B.n830 B.n17 585
R411 B.n17 B.n16 585
R412 B.n829 B.n828 585
R413 B.n828 B.n827 585
R414 B.n19 B.n18 585
R415 B.n826 B.n19 585
R416 B.n824 B.n823 585
R417 B.n825 B.n824 585
R418 B.n822 B.n24 585
R419 B.n24 B.n23 585
R420 B.n821 B.n820 585
R421 B.n820 B.n819 585
R422 B.n26 B.n25 585
R423 B.n818 B.n26 585
R424 B.n816 B.n815 585
R425 B.n817 B.n816 585
R426 B.n814 B.n31 585
R427 B.n31 B.n30 585
R428 B.n813 B.n812 585
R429 B.n812 B.n811 585
R430 B.n33 B.n32 585
R431 B.n810 B.n33 585
R432 B.n808 B.n807 585
R433 B.n809 B.n808 585
R434 B.n806 B.n38 585
R435 B.n38 B.n37 585
R436 B.n805 B.n804 585
R437 B.n804 B.n803 585
R438 B.n40 B.n39 585
R439 B.n802 B.n40 585
R440 B.n800 B.n799 585
R441 B.n801 B.n800 585
R442 B.n798 B.n45 585
R443 B.n45 B.n44 585
R444 B.n797 B.n796 585
R445 B.n796 B.n795 585
R446 B.n47 B.n46 585
R447 B.n794 B.n47 585
R448 B.n792 B.n791 585
R449 B.n793 B.n792 585
R450 B.n790 B.n52 585
R451 B.n52 B.n51 585
R452 B.n789 B.n788 585
R453 B.n788 B.n787 585
R454 B.n54 B.n53 585
R455 B.n786 B.n54 585
R456 B.n784 B.n783 585
R457 B.n785 B.n784 585
R458 B.n782 B.n59 585
R459 B.n59 B.n58 585
R460 B.n845 B.n844 585
R461 B.n843 B.n2 585
R462 B.n780 B.n59 506.916
R463 B.n777 B.n113 506.916
R464 B.n437 B.n376 506.916
R465 B.n641 B.n378 506.916
R466 B.n117 B.t13 347.724
R467 B.n114 B.t6 347.724
R468 B.n435 B.t2 347.724
R469 B.n432 B.t10 347.724
R470 B.n778 B.n111 256.663
R471 B.n778 B.n110 256.663
R472 B.n778 B.n109 256.663
R473 B.n778 B.n108 256.663
R474 B.n778 B.n107 256.663
R475 B.n778 B.n106 256.663
R476 B.n778 B.n105 256.663
R477 B.n778 B.n104 256.663
R478 B.n778 B.n103 256.663
R479 B.n778 B.n102 256.663
R480 B.n778 B.n101 256.663
R481 B.n778 B.n100 256.663
R482 B.n778 B.n99 256.663
R483 B.n778 B.n98 256.663
R484 B.n778 B.n97 256.663
R485 B.n778 B.n96 256.663
R486 B.n778 B.n95 256.663
R487 B.n778 B.n94 256.663
R488 B.n778 B.n93 256.663
R489 B.n778 B.n92 256.663
R490 B.n778 B.n91 256.663
R491 B.n778 B.n90 256.663
R492 B.n778 B.n89 256.663
R493 B.n778 B.n88 256.663
R494 B.n778 B.n87 256.663
R495 B.n778 B.n86 256.663
R496 B.n778 B.n85 256.663
R497 B.n778 B.n84 256.663
R498 B.n778 B.n83 256.663
R499 B.n778 B.n82 256.663
R500 B.n778 B.n81 256.663
R501 B.n778 B.n80 256.663
R502 B.n778 B.n79 256.663
R503 B.n778 B.n78 256.663
R504 B.n778 B.n77 256.663
R505 B.n778 B.n76 256.663
R506 B.n778 B.n75 256.663
R507 B.n778 B.n74 256.663
R508 B.n778 B.n73 256.663
R509 B.n778 B.n72 256.663
R510 B.n778 B.n71 256.663
R511 B.n778 B.n70 256.663
R512 B.n778 B.n69 256.663
R513 B.n778 B.n68 256.663
R514 B.n778 B.n67 256.663
R515 B.n778 B.n66 256.663
R516 B.n778 B.n65 256.663
R517 B.n778 B.n64 256.663
R518 B.n778 B.n63 256.663
R519 B.n778 B.n62 256.663
R520 B.n779 B.n778 256.663
R521 B.n640 B.n639 256.663
R522 B.n639 B.n381 256.663
R523 B.n639 B.n382 256.663
R524 B.n639 B.n383 256.663
R525 B.n639 B.n384 256.663
R526 B.n639 B.n385 256.663
R527 B.n639 B.n386 256.663
R528 B.n639 B.n387 256.663
R529 B.n639 B.n388 256.663
R530 B.n639 B.n389 256.663
R531 B.n639 B.n390 256.663
R532 B.n639 B.n391 256.663
R533 B.n639 B.n392 256.663
R534 B.n639 B.n393 256.663
R535 B.n639 B.n394 256.663
R536 B.n639 B.n395 256.663
R537 B.n639 B.n396 256.663
R538 B.n639 B.n397 256.663
R539 B.n639 B.n398 256.663
R540 B.n639 B.n399 256.663
R541 B.n639 B.n400 256.663
R542 B.n639 B.n401 256.663
R543 B.n639 B.n402 256.663
R544 B.n639 B.n403 256.663
R545 B.n639 B.n404 256.663
R546 B.n639 B.n405 256.663
R547 B.n639 B.n406 256.663
R548 B.n639 B.n407 256.663
R549 B.n639 B.n408 256.663
R550 B.n639 B.n409 256.663
R551 B.n639 B.n410 256.663
R552 B.n639 B.n411 256.663
R553 B.n639 B.n412 256.663
R554 B.n639 B.n413 256.663
R555 B.n639 B.n414 256.663
R556 B.n639 B.n415 256.663
R557 B.n639 B.n416 256.663
R558 B.n639 B.n417 256.663
R559 B.n639 B.n418 256.663
R560 B.n639 B.n419 256.663
R561 B.n639 B.n420 256.663
R562 B.n639 B.n421 256.663
R563 B.n639 B.n422 256.663
R564 B.n639 B.n423 256.663
R565 B.n639 B.n424 256.663
R566 B.n639 B.n425 256.663
R567 B.n639 B.n426 256.663
R568 B.n639 B.n427 256.663
R569 B.n639 B.n428 256.663
R570 B.n639 B.n429 256.663
R571 B.n639 B.n430 256.663
R572 B.n847 B.n846 256.663
R573 B.n119 B.n61 163.367
R574 B.n123 B.n122 163.367
R575 B.n127 B.n126 163.367
R576 B.n131 B.n130 163.367
R577 B.n135 B.n134 163.367
R578 B.n139 B.n138 163.367
R579 B.n143 B.n142 163.367
R580 B.n147 B.n146 163.367
R581 B.n151 B.n150 163.367
R582 B.n155 B.n154 163.367
R583 B.n159 B.n158 163.367
R584 B.n163 B.n162 163.367
R585 B.n167 B.n166 163.367
R586 B.n171 B.n170 163.367
R587 B.n175 B.n174 163.367
R588 B.n179 B.n178 163.367
R589 B.n183 B.n182 163.367
R590 B.n187 B.n186 163.367
R591 B.n191 B.n190 163.367
R592 B.n195 B.n194 163.367
R593 B.n199 B.n198 163.367
R594 B.n203 B.n202 163.367
R595 B.n207 B.n206 163.367
R596 B.n212 B.n211 163.367
R597 B.n216 B.n215 163.367
R598 B.n220 B.n219 163.367
R599 B.n224 B.n223 163.367
R600 B.n228 B.n227 163.367
R601 B.n232 B.n231 163.367
R602 B.n236 B.n235 163.367
R603 B.n240 B.n239 163.367
R604 B.n244 B.n243 163.367
R605 B.n248 B.n247 163.367
R606 B.n252 B.n251 163.367
R607 B.n256 B.n255 163.367
R608 B.n260 B.n259 163.367
R609 B.n264 B.n263 163.367
R610 B.n268 B.n267 163.367
R611 B.n272 B.n271 163.367
R612 B.n276 B.n275 163.367
R613 B.n280 B.n279 163.367
R614 B.n284 B.n283 163.367
R615 B.n288 B.n287 163.367
R616 B.n292 B.n291 163.367
R617 B.n296 B.n295 163.367
R618 B.n300 B.n299 163.367
R619 B.n304 B.n303 163.367
R620 B.n308 B.n307 163.367
R621 B.n312 B.n311 163.367
R622 B.n316 B.n315 163.367
R623 B.n777 B.n112 163.367
R624 B.n647 B.n376 163.367
R625 B.n647 B.n374 163.367
R626 B.n651 B.n374 163.367
R627 B.n651 B.n367 163.367
R628 B.n659 B.n367 163.367
R629 B.n659 B.n365 163.367
R630 B.n663 B.n365 163.367
R631 B.n663 B.n360 163.367
R632 B.n671 B.n360 163.367
R633 B.n671 B.n358 163.367
R634 B.n675 B.n358 163.367
R635 B.n675 B.n352 163.367
R636 B.n683 B.n352 163.367
R637 B.n683 B.n350 163.367
R638 B.n687 B.n350 163.367
R639 B.n687 B.n343 163.367
R640 B.n695 B.n343 163.367
R641 B.n695 B.n341 163.367
R642 B.n699 B.n341 163.367
R643 B.n699 B.n336 163.367
R644 B.n707 B.n336 163.367
R645 B.n707 B.n334 163.367
R646 B.n711 B.n334 163.367
R647 B.n711 B.n328 163.367
R648 B.n719 B.n328 163.367
R649 B.n719 B.n326 163.367
R650 B.n724 B.n326 163.367
R651 B.n724 B.n320 163.367
R652 B.n732 B.n320 163.367
R653 B.n733 B.n732 163.367
R654 B.n733 B.n5 163.367
R655 B.n6 B.n5 163.367
R656 B.n7 B.n6 163.367
R657 B.n739 B.n7 163.367
R658 B.n740 B.n739 163.367
R659 B.n740 B.n13 163.367
R660 B.n14 B.n13 163.367
R661 B.n15 B.n14 163.367
R662 B.n745 B.n15 163.367
R663 B.n745 B.n20 163.367
R664 B.n21 B.n20 163.367
R665 B.n22 B.n21 163.367
R666 B.n750 B.n22 163.367
R667 B.n750 B.n27 163.367
R668 B.n28 B.n27 163.367
R669 B.n29 B.n28 163.367
R670 B.n755 B.n29 163.367
R671 B.n755 B.n34 163.367
R672 B.n35 B.n34 163.367
R673 B.n36 B.n35 163.367
R674 B.n760 B.n36 163.367
R675 B.n760 B.n41 163.367
R676 B.n42 B.n41 163.367
R677 B.n43 B.n42 163.367
R678 B.n765 B.n43 163.367
R679 B.n765 B.n48 163.367
R680 B.n49 B.n48 163.367
R681 B.n50 B.n49 163.367
R682 B.n770 B.n50 163.367
R683 B.n770 B.n55 163.367
R684 B.n56 B.n55 163.367
R685 B.n57 B.n56 163.367
R686 B.n113 B.n57 163.367
R687 B.n638 B.n380 163.367
R688 B.n638 B.n431 163.367
R689 B.n634 B.n633 163.367
R690 B.n630 B.n629 163.367
R691 B.n626 B.n625 163.367
R692 B.n622 B.n621 163.367
R693 B.n618 B.n617 163.367
R694 B.n614 B.n613 163.367
R695 B.n610 B.n609 163.367
R696 B.n606 B.n605 163.367
R697 B.n602 B.n601 163.367
R698 B.n598 B.n597 163.367
R699 B.n594 B.n593 163.367
R700 B.n590 B.n589 163.367
R701 B.n586 B.n585 163.367
R702 B.n582 B.n581 163.367
R703 B.n578 B.n577 163.367
R704 B.n574 B.n573 163.367
R705 B.n570 B.n569 163.367
R706 B.n566 B.n565 163.367
R707 B.n562 B.n561 163.367
R708 B.n558 B.n557 163.367
R709 B.n554 B.n553 163.367
R710 B.n550 B.n549 163.367
R711 B.n546 B.n545 163.367
R712 B.n542 B.n541 163.367
R713 B.n538 B.n537 163.367
R714 B.n534 B.n533 163.367
R715 B.n529 B.n528 163.367
R716 B.n525 B.n524 163.367
R717 B.n521 B.n520 163.367
R718 B.n517 B.n516 163.367
R719 B.n513 B.n512 163.367
R720 B.n509 B.n508 163.367
R721 B.n505 B.n504 163.367
R722 B.n501 B.n500 163.367
R723 B.n497 B.n496 163.367
R724 B.n493 B.n492 163.367
R725 B.n489 B.n488 163.367
R726 B.n485 B.n484 163.367
R727 B.n481 B.n480 163.367
R728 B.n477 B.n476 163.367
R729 B.n473 B.n472 163.367
R730 B.n469 B.n468 163.367
R731 B.n465 B.n464 163.367
R732 B.n461 B.n460 163.367
R733 B.n457 B.n456 163.367
R734 B.n453 B.n452 163.367
R735 B.n449 B.n448 163.367
R736 B.n445 B.n444 163.367
R737 B.n441 B.n440 163.367
R738 B.n645 B.n378 163.367
R739 B.n645 B.n372 163.367
R740 B.n653 B.n372 163.367
R741 B.n653 B.n370 163.367
R742 B.n657 B.n370 163.367
R743 B.n657 B.n364 163.367
R744 B.n665 B.n364 163.367
R745 B.n665 B.n362 163.367
R746 B.n669 B.n362 163.367
R747 B.n669 B.n356 163.367
R748 B.n677 B.n356 163.367
R749 B.n677 B.n354 163.367
R750 B.n681 B.n354 163.367
R751 B.n681 B.n348 163.367
R752 B.n689 B.n348 163.367
R753 B.n689 B.n346 163.367
R754 B.n693 B.n346 163.367
R755 B.n693 B.n340 163.367
R756 B.n701 B.n340 163.367
R757 B.n701 B.n338 163.367
R758 B.n705 B.n338 163.367
R759 B.n705 B.n332 163.367
R760 B.n713 B.n332 163.367
R761 B.n713 B.n330 163.367
R762 B.n717 B.n330 163.367
R763 B.n717 B.n324 163.367
R764 B.n726 B.n324 163.367
R765 B.n726 B.n322 163.367
R766 B.n730 B.n322 163.367
R767 B.n730 B.n3 163.367
R768 B.n845 B.n3 163.367
R769 B.n841 B.n2 163.367
R770 B.n841 B.n840 163.367
R771 B.n840 B.n9 163.367
R772 B.n836 B.n9 163.367
R773 B.n836 B.n11 163.367
R774 B.n832 B.n11 163.367
R775 B.n832 B.n17 163.367
R776 B.n828 B.n17 163.367
R777 B.n828 B.n19 163.367
R778 B.n824 B.n19 163.367
R779 B.n824 B.n24 163.367
R780 B.n820 B.n24 163.367
R781 B.n820 B.n26 163.367
R782 B.n816 B.n26 163.367
R783 B.n816 B.n31 163.367
R784 B.n812 B.n31 163.367
R785 B.n812 B.n33 163.367
R786 B.n808 B.n33 163.367
R787 B.n808 B.n38 163.367
R788 B.n804 B.n38 163.367
R789 B.n804 B.n40 163.367
R790 B.n800 B.n40 163.367
R791 B.n800 B.n45 163.367
R792 B.n796 B.n45 163.367
R793 B.n796 B.n47 163.367
R794 B.n792 B.n47 163.367
R795 B.n792 B.n52 163.367
R796 B.n788 B.n52 163.367
R797 B.n788 B.n54 163.367
R798 B.n784 B.n54 163.367
R799 B.n784 B.n59 163.367
R800 B.n114 B.t8 120.731
R801 B.n435 B.t5 120.731
R802 B.n117 B.t14 120.713
R803 B.n432 B.t12 120.713
R804 B.n639 B.n377 81.9123
R805 B.n778 B.n58 81.9123
R806 B.n780 B.n779 71.676
R807 B.n119 B.n62 71.676
R808 B.n123 B.n63 71.676
R809 B.n127 B.n64 71.676
R810 B.n131 B.n65 71.676
R811 B.n135 B.n66 71.676
R812 B.n139 B.n67 71.676
R813 B.n143 B.n68 71.676
R814 B.n147 B.n69 71.676
R815 B.n151 B.n70 71.676
R816 B.n155 B.n71 71.676
R817 B.n159 B.n72 71.676
R818 B.n163 B.n73 71.676
R819 B.n167 B.n74 71.676
R820 B.n171 B.n75 71.676
R821 B.n175 B.n76 71.676
R822 B.n179 B.n77 71.676
R823 B.n183 B.n78 71.676
R824 B.n187 B.n79 71.676
R825 B.n191 B.n80 71.676
R826 B.n195 B.n81 71.676
R827 B.n199 B.n82 71.676
R828 B.n203 B.n83 71.676
R829 B.n207 B.n84 71.676
R830 B.n212 B.n85 71.676
R831 B.n216 B.n86 71.676
R832 B.n220 B.n87 71.676
R833 B.n224 B.n88 71.676
R834 B.n228 B.n89 71.676
R835 B.n232 B.n90 71.676
R836 B.n236 B.n91 71.676
R837 B.n240 B.n92 71.676
R838 B.n244 B.n93 71.676
R839 B.n248 B.n94 71.676
R840 B.n252 B.n95 71.676
R841 B.n256 B.n96 71.676
R842 B.n260 B.n97 71.676
R843 B.n264 B.n98 71.676
R844 B.n268 B.n99 71.676
R845 B.n272 B.n100 71.676
R846 B.n276 B.n101 71.676
R847 B.n280 B.n102 71.676
R848 B.n284 B.n103 71.676
R849 B.n288 B.n104 71.676
R850 B.n292 B.n105 71.676
R851 B.n296 B.n106 71.676
R852 B.n300 B.n107 71.676
R853 B.n304 B.n108 71.676
R854 B.n308 B.n109 71.676
R855 B.n312 B.n110 71.676
R856 B.n316 B.n111 71.676
R857 B.n112 B.n111 71.676
R858 B.n315 B.n110 71.676
R859 B.n311 B.n109 71.676
R860 B.n307 B.n108 71.676
R861 B.n303 B.n107 71.676
R862 B.n299 B.n106 71.676
R863 B.n295 B.n105 71.676
R864 B.n291 B.n104 71.676
R865 B.n287 B.n103 71.676
R866 B.n283 B.n102 71.676
R867 B.n279 B.n101 71.676
R868 B.n275 B.n100 71.676
R869 B.n271 B.n99 71.676
R870 B.n267 B.n98 71.676
R871 B.n263 B.n97 71.676
R872 B.n259 B.n96 71.676
R873 B.n255 B.n95 71.676
R874 B.n251 B.n94 71.676
R875 B.n247 B.n93 71.676
R876 B.n243 B.n92 71.676
R877 B.n239 B.n91 71.676
R878 B.n235 B.n90 71.676
R879 B.n231 B.n89 71.676
R880 B.n227 B.n88 71.676
R881 B.n223 B.n87 71.676
R882 B.n219 B.n86 71.676
R883 B.n215 B.n85 71.676
R884 B.n211 B.n84 71.676
R885 B.n206 B.n83 71.676
R886 B.n202 B.n82 71.676
R887 B.n198 B.n81 71.676
R888 B.n194 B.n80 71.676
R889 B.n190 B.n79 71.676
R890 B.n186 B.n78 71.676
R891 B.n182 B.n77 71.676
R892 B.n178 B.n76 71.676
R893 B.n174 B.n75 71.676
R894 B.n170 B.n74 71.676
R895 B.n166 B.n73 71.676
R896 B.n162 B.n72 71.676
R897 B.n158 B.n71 71.676
R898 B.n154 B.n70 71.676
R899 B.n150 B.n69 71.676
R900 B.n146 B.n68 71.676
R901 B.n142 B.n67 71.676
R902 B.n138 B.n66 71.676
R903 B.n134 B.n65 71.676
R904 B.n130 B.n64 71.676
R905 B.n126 B.n63 71.676
R906 B.n122 B.n62 71.676
R907 B.n779 B.n61 71.676
R908 B.n641 B.n640 71.676
R909 B.n431 B.n381 71.676
R910 B.n633 B.n382 71.676
R911 B.n629 B.n383 71.676
R912 B.n625 B.n384 71.676
R913 B.n621 B.n385 71.676
R914 B.n617 B.n386 71.676
R915 B.n613 B.n387 71.676
R916 B.n609 B.n388 71.676
R917 B.n605 B.n389 71.676
R918 B.n601 B.n390 71.676
R919 B.n597 B.n391 71.676
R920 B.n593 B.n392 71.676
R921 B.n589 B.n393 71.676
R922 B.n585 B.n394 71.676
R923 B.n581 B.n395 71.676
R924 B.n577 B.n396 71.676
R925 B.n573 B.n397 71.676
R926 B.n569 B.n398 71.676
R927 B.n565 B.n399 71.676
R928 B.n561 B.n400 71.676
R929 B.n557 B.n401 71.676
R930 B.n553 B.n402 71.676
R931 B.n549 B.n403 71.676
R932 B.n545 B.n404 71.676
R933 B.n541 B.n405 71.676
R934 B.n537 B.n406 71.676
R935 B.n533 B.n407 71.676
R936 B.n528 B.n408 71.676
R937 B.n524 B.n409 71.676
R938 B.n520 B.n410 71.676
R939 B.n516 B.n411 71.676
R940 B.n512 B.n412 71.676
R941 B.n508 B.n413 71.676
R942 B.n504 B.n414 71.676
R943 B.n500 B.n415 71.676
R944 B.n496 B.n416 71.676
R945 B.n492 B.n417 71.676
R946 B.n488 B.n418 71.676
R947 B.n484 B.n419 71.676
R948 B.n480 B.n420 71.676
R949 B.n476 B.n421 71.676
R950 B.n472 B.n422 71.676
R951 B.n468 B.n423 71.676
R952 B.n464 B.n424 71.676
R953 B.n460 B.n425 71.676
R954 B.n456 B.n426 71.676
R955 B.n452 B.n427 71.676
R956 B.n448 B.n428 71.676
R957 B.n444 B.n429 71.676
R958 B.n440 B.n430 71.676
R959 B.n640 B.n380 71.676
R960 B.n634 B.n381 71.676
R961 B.n630 B.n382 71.676
R962 B.n626 B.n383 71.676
R963 B.n622 B.n384 71.676
R964 B.n618 B.n385 71.676
R965 B.n614 B.n386 71.676
R966 B.n610 B.n387 71.676
R967 B.n606 B.n388 71.676
R968 B.n602 B.n389 71.676
R969 B.n598 B.n390 71.676
R970 B.n594 B.n391 71.676
R971 B.n590 B.n392 71.676
R972 B.n586 B.n393 71.676
R973 B.n582 B.n394 71.676
R974 B.n578 B.n395 71.676
R975 B.n574 B.n396 71.676
R976 B.n570 B.n397 71.676
R977 B.n566 B.n398 71.676
R978 B.n562 B.n399 71.676
R979 B.n558 B.n400 71.676
R980 B.n554 B.n401 71.676
R981 B.n550 B.n402 71.676
R982 B.n546 B.n403 71.676
R983 B.n542 B.n404 71.676
R984 B.n538 B.n405 71.676
R985 B.n534 B.n406 71.676
R986 B.n529 B.n407 71.676
R987 B.n525 B.n408 71.676
R988 B.n521 B.n409 71.676
R989 B.n517 B.n410 71.676
R990 B.n513 B.n411 71.676
R991 B.n509 B.n412 71.676
R992 B.n505 B.n413 71.676
R993 B.n501 B.n414 71.676
R994 B.n497 B.n415 71.676
R995 B.n493 B.n416 71.676
R996 B.n489 B.n417 71.676
R997 B.n485 B.n418 71.676
R998 B.n481 B.n419 71.676
R999 B.n477 B.n420 71.676
R1000 B.n473 B.n421 71.676
R1001 B.n469 B.n422 71.676
R1002 B.n465 B.n423 71.676
R1003 B.n461 B.n424 71.676
R1004 B.n457 B.n425 71.676
R1005 B.n453 B.n426 71.676
R1006 B.n449 B.n427 71.676
R1007 B.n445 B.n428 71.676
R1008 B.n441 B.n429 71.676
R1009 B.n437 B.n430 71.676
R1010 B.n846 B.n845 71.676
R1011 B.n846 B.n2 71.676
R1012 B.n115 B.t9 68.7555
R1013 B.n436 B.t4 68.7555
R1014 B.n118 B.t15 68.7378
R1015 B.n433 B.t11 68.7378
R1016 B.n209 B.n118 59.5399
R1017 B.n116 B.n115 59.5399
R1018 B.n531 B.n436 59.5399
R1019 B.n434 B.n433 59.5399
R1020 B.n118 B.n117 51.9763
R1021 B.n115 B.n114 51.9763
R1022 B.n436 B.n435 51.9763
R1023 B.n433 B.n432 51.9763
R1024 B.n646 B.n377 39.5041
R1025 B.n646 B.n373 39.5041
R1026 B.n652 B.n373 39.5041
R1027 B.n652 B.n368 39.5041
R1028 B.n658 B.n368 39.5041
R1029 B.n658 B.n369 39.5041
R1030 B.n664 B.n361 39.5041
R1031 B.n670 B.n361 39.5041
R1032 B.n670 B.n357 39.5041
R1033 B.n676 B.n357 39.5041
R1034 B.n676 B.n353 39.5041
R1035 B.n682 B.n353 39.5041
R1036 B.n682 B.n349 39.5041
R1037 B.n688 B.n349 39.5041
R1038 B.n688 B.n344 39.5041
R1039 B.n694 B.n344 39.5041
R1040 B.n694 B.n345 39.5041
R1041 B.n700 B.n337 39.5041
R1042 B.n706 B.n337 39.5041
R1043 B.n706 B.n333 39.5041
R1044 B.n712 B.n333 39.5041
R1045 B.n712 B.n329 39.5041
R1046 B.n718 B.n329 39.5041
R1047 B.n725 B.n325 39.5041
R1048 B.n725 B.n321 39.5041
R1049 B.n731 B.n321 39.5041
R1050 B.n731 B.n4 39.5041
R1051 B.n844 B.n4 39.5041
R1052 B.n844 B.n843 39.5041
R1053 B.n843 B.n842 39.5041
R1054 B.n842 B.n8 39.5041
R1055 B.n12 B.n8 39.5041
R1056 B.n835 B.n12 39.5041
R1057 B.n835 B.n834 39.5041
R1058 B.n833 B.n16 39.5041
R1059 B.n827 B.n16 39.5041
R1060 B.n827 B.n826 39.5041
R1061 B.n826 B.n825 39.5041
R1062 B.n825 B.n23 39.5041
R1063 B.n819 B.n23 39.5041
R1064 B.n818 B.n817 39.5041
R1065 B.n817 B.n30 39.5041
R1066 B.n811 B.n30 39.5041
R1067 B.n811 B.n810 39.5041
R1068 B.n810 B.n809 39.5041
R1069 B.n809 B.n37 39.5041
R1070 B.n803 B.n37 39.5041
R1071 B.n803 B.n802 39.5041
R1072 B.n802 B.n801 39.5041
R1073 B.n801 B.n44 39.5041
R1074 B.n795 B.n44 39.5041
R1075 B.n794 B.n793 39.5041
R1076 B.n793 B.n51 39.5041
R1077 B.n787 B.n51 39.5041
R1078 B.n787 B.n786 39.5041
R1079 B.n786 B.n785 39.5041
R1080 B.n785 B.n58 39.5041
R1081 B.n369 B.t3 38.9231
R1082 B.t7 B.n794 38.9231
R1083 B.n718 B.t17 37.7613
R1084 B.t0 B.n833 37.7613
R1085 B.n700 B.t16 36.5994
R1086 B.n819 B.t1 36.5994
R1087 B.n643 B.n642 32.9371
R1088 B.n438 B.n375 32.9371
R1089 B.n776 B.n775 32.9371
R1090 B.n782 B.n781 32.9371
R1091 B B.n847 18.0485
R1092 B.n644 B.n643 10.6151
R1093 B.n644 B.n371 10.6151
R1094 B.n654 B.n371 10.6151
R1095 B.n655 B.n654 10.6151
R1096 B.n656 B.n655 10.6151
R1097 B.n656 B.n363 10.6151
R1098 B.n666 B.n363 10.6151
R1099 B.n667 B.n666 10.6151
R1100 B.n668 B.n667 10.6151
R1101 B.n668 B.n355 10.6151
R1102 B.n678 B.n355 10.6151
R1103 B.n679 B.n678 10.6151
R1104 B.n680 B.n679 10.6151
R1105 B.n680 B.n347 10.6151
R1106 B.n690 B.n347 10.6151
R1107 B.n691 B.n690 10.6151
R1108 B.n692 B.n691 10.6151
R1109 B.n692 B.n339 10.6151
R1110 B.n702 B.n339 10.6151
R1111 B.n703 B.n702 10.6151
R1112 B.n704 B.n703 10.6151
R1113 B.n704 B.n331 10.6151
R1114 B.n714 B.n331 10.6151
R1115 B.n715 B.n714 10.6151
R1116 B.n716 B.n715 10.6151
R1117 B.n716 B.n323 10.6151
R1118 B.n727 B.n323 10.6151
R1119 B.n728 B.n727 10.6151
R1120 B.n729 B.n728 10.6151
R1121 B.n729 B.n0 10.6151
R1122 B.n642 B.n379 10.6151
R1123 B.n637 B.n379 10.6151
R1124 B.n637 B.n636 10.6151
R1125 B.n636 B.n635 10.6151
R1126 B.n635 B.n632 10.6151
R1127 B.n632 B.n631 10.6151
R1128 B.n631 B.n628 10.6151
R1129 B.n628 B.n627 10.6151
R1130 B.n627 B.n624 10.6151
R1131 B.n624 B.n623 10.6151
R1132 B.n623 B.n620 10.6151
R1133 B.n620 B.n619 10.6151
R1134 B.n619 B.n616 10.6151
R1135 B.n616 B.n615 10.6151
R1136 B.n615 B.n612 10.6151
R1137 B.n612 B.n611 10.6151
R1138 B.n611 B.n608 10.6151
R1139 B.n608 B.n607 10.6151
R1140 B.n607 B.n604 10.6151
R1141 B.n604 B.n603 10.6151
R1142 B.n603 B.n600 10.6151
R1143 B.n600 B.n599 10.6151
R1144 B.n599 B.n596 10.6151
R1145 B.n596 B.n595 10.6151
R1146 B.n595 B.n592 10.6151
R1147 B.n592 B.n591 10.6151
R1148 B.n591 B.n588 10.6151
R1149 B.n588 B.n587 10.6151
R1150 B.n587 B.n584 10.6151
R1151 B.n584 B.n583 10.6151
R1152 B.n583 B.n580 10.6151
R1153 B.n580 B.n579 10.6151
R1154 B.n579 B.n576 10.6151
R1155 B.n576 B.n575 10.6151
R1156 B.n575 B.n572 10.6151
R1157 B.n572 B.n571 10.6151
R1158 B.n571 B.n568 10.6151
R1159 B.n568 B.n567 10.6151
R1160 B.n567 B.n564 10.6151
R1161 B.n564 B.n563 10.6151
R1162 B.n563 B.n560 10.6151
R1163 B.n560 B.n559 10.6151
R1164 B.n559 B.n556 10.6151
R1165 B.n556 B.n555 10.6151
R1166 B.n555 B.n552 10.6151
R1167 B.n552 B.n551 10.6151
R1168 B.n548 B.n547 10.6151
R1169 B.n547 B.n544 10.6151
R1170 B.n544 B.n543 10.6151
R1171 B.n543 B.n540 10.6151
R1172 B.n540 B.n539 10.6151
R1173 B.n539 B.n536 10.6151
R1174 B.n536 B.n535 10.6151
R1175 B.n535 B.n532 10.6151
R1176 B.n530 B.n527 10.6151
R1177 B.n527 B.n526 10.6151
R1178 B.n526 B.n523 10.6151
R1179 B.n523 B.n522 10.6151
R1180 B.n522 B.n519 10.6151
R1181 B.n519 B.n518 10.6151
R1182 B.n518 B.n515 10.6151
R1183 B.n515 B.n514 10.6151
R1184 B.n514 B.n511 10.6151
R1185 B.n511 B.n510 10.6151
R1186 B.n510 B.n507 10.6151
R1187 B.n507 B.n506 10.6151
R1188 B.n506 B.n503 10.6151
R1189 B.n503 B.n502 10.6151
R1190 B.n502 B.n499 10.6151
R1191 B.n499 B.n498 10.6151
R1192 B.n498 B.n495 10.6151
R1193 B.n495 B.n494 10.6151
R1194 B.n494 B.n491 10.6151
R1195 B.n491 B.n490 10.6151
R1196 B.n490 B.n487 10.6151
R1197 B.n487 B.n486 10.6151
R1198 B.n486 B.n483 10.6151
R1199 B.n483 B.n482 10.6151
R1200 B.n482 B.n479 10.6151
R1201 B.n479 B.n478 10.6151
R1202 B.n478 B.n475 10.6151
R1203 B.n475 B.n474 10.6151
R1204 B.n474 B.n471 10.6151
R1205 B.n471 B.n470 10.6151
R1206 B.n470 B.n467 10.6151
R1207 B.n467 B.n466 10.6151
R1208 B.n466 B.n463 10.6151
R1209 B.n463 B.n462 10.6151
R1210 B.n462 B.n459 10.6151
R1211 B.n459 B.n458 10.6151
R1212 B.n458 B.n455 10.6151
R1213 B.n455 B.n454 10.6151
R1214 B.n454 B.n451 10.6151
R1215 B.n451 B.n450 10.6151
R1216 B.n450 B.n447 10.6151
R1217 B.n447 B.n446 10.6151
R1218 B.n446 B.n443 10.6151
R1219 B.n443 B.n442 10.6151
R1220 B.n442 B.n439 10.6151
R1221 B.n439 B.n438 10.6151
R1222 B.n648 B.n375 10.6151
R1223 B.n649 B.n648 10.6151
R1224 B.n650 B.n649 10.6151
R1225 B.n650 B.n366 10.6151
R1226 B.n660 B.n366 10.6151
R1227 B.n661 B.n660 10.6151
R1228 B.n662 B.n661 10.6151
R1229 B.n662 B.n359 10.6151
R1230 B.n672 B.n359 10.6151
R1231 B.n673 B.n672 10.6151
R1232 B.n674 B.n673 10.6151
R1233 B.n674 B.n351 10.6151
R1234 B.n684 B.n351 10.6151
R1235 B.n685 B.n684 10.6151
R1236 B.n686 B.n685 10.6151
R1237 B.n686 B.n342 10.6151
R1238 B.n696 B.n342 10.6151
R1239 B.n697 B.n696 10.6151
R1240 B.n698 B.n697 10.6151
R1241 B.n698 B.n335 10.6151
R1242 B.n708 B.n335 10.6151
R1243 B.n709 B.n708 10.6151
R1244 B.n710 B.n709 10.6151
R1245 B.n710 B.n327 10.6151
R1246 B.n720 B.n327 10.6151
R1247 B.n721 B.n720 10.6151
R1248 B.n723 B.n721 10.6151
R1249 B.n723 B.n722 10.6151
R1250 B.n722 B.n319 10.6151
R1251 B.n734 B.n319 10.6151
R1252 B.n735 B.n734 10.6151
R1253 B.n736 B.n735 10.6151
R1254 B.n737 B.n736 10.6151
R1255 B.n738 B.n737 10.6151
R1256 B.n741 B.n738 10.6151
R1257 B.n742 B.n741 10.6151
R1258 B.n743 B.n742 10.6151
R1259 B.n744 B.n743 10.6151
R1260 B.n746 B.n744 10.6151
R1261 B.n747 B.n746 10.6151
R1262 B.n748 B.n747 10.6151
R1263 B.n749 B.n748 10.6151
R1264 B.n751 B.n749 10.6151
R1265 B.n752 B.n751 10.6151
R1266 B.n753 B.n752 10.6151
R1267 B.n754 B.n753 10.6151
R1268 B.n756 B.n754 10.6151
R1269 B.n757 B.n756 10.6151
R1270 B.n758 B.n757 10.6151
R1271 B.n759 B.n758 10.6151
R1272 B.n761 B.n759 10.6151
R1273 B.n762 B.n761 10.6151
R1274 B.n763 B.n762 10.6151
R1275 B.n764 B.n763 10.6151
R1276 B.n766 B.n764 10.6151
R1277 B.n767 B.n766 10.6151
R1278 B.n768 B.n767 10.6151
R1279 B.n769 B.n768 10.6151
R1280 B.n771 B.n769 10.6151
R1281 B.n772 B.n771 10.6151
R1282 B.n773 B.n772 10.6151
R1283 B.n774 B.n773 10.6151
R1284 B.n775 B.n774 10.6151
R1285 B.n839 B.n1 10.6151
R1286 B.n839 B.n838 10.6151
R1287 B.n838 B.n837 10.6151
R1288 B.n837 B.n10 10.6151
R1289 B.n831 B.n10 10.6151
R1290 B.n831 B.n830 10.6151
R1291 B.n830 B.n829 10.6151
R1292 B.n829 B.n18 10.6151
R1293 B.n823 B.n18 10.6151
R1294 B.n823 B.n822 10.6151
R1295 B.n822 B.n821 10.6151
R1296 B.n821 B.n25 10.6151
R1297 B.n815 B.n25 10.6151
R1298 B.n815 B.n814 10.6151
R1299 B.n814 B.n813 10.6151
R1300 B.n813 B.n32 10.6151
R1301 B.n807 B.n32 10.6151
R1302 B.n807 B.n806 10.6151
R1303 B.n806 B.n805 10.6151
R1304 B.n805 B.n39 10.6151
R1305 B.n799 B.n39 10.6151
R1306 B.n799 B.n798 10.6151
R1307 B.n798 B.n797 10.6151
R1308 B.n797 B.n46 10.6151
R1309 B.n791 B.n46 10.6151
R1310 B.n791 B.n790 10.6151
R1311 B.n790 B.n789 10.6151
R1312 B.n789 B.n53 10.6151
R1313 B.n783 B.n53 10.6151
R1314 B.n783 B.n782 10.6151
R1315 B.n781 B.n60 10.6151
R1316 B.n120 B.n60 10.6151
R1317 B.n121 B.n120 10.6151
R1318 B.n124 B.n121 10.6151
R1319 B.n125 B.n124 10.6151
R1320 B.n128 B.n125 10.6151
R1321 B.n129 B.n128 10.6151
R1322 B.n132 B.n129 10.6151
R1323 B.n133 B.n132 10.6151
R1324 B.n136 B.n133 10.6151
R1325 B.n137 B.n136 10.6151
R1326 B.n140 B.n137 10.6151
R1327 B.n141 B.n140 10.6151
R1328 B.n144 B.n141 10.6151
R1329 B.n145 B.n144 10.6151
R1330 B.n148 B.n145 10.6151
R1331 B.n149 B.n148 10.6151
R1332 B.n152 B.n149 10.6151
R1333 B.n153 B.n152 10.6151
R1334 B.n156 B.n153 10.6151
R1335 B.n157 B.n156 10.6151
R1336 B.n160 B.n157 10.6151
R1337 B.n161 B.n160 10.6151
R1338 B.n164 B.n161 10.6151
R1339 B.n165 B.n164 10.6151
R1340 B.n168 B.n165 10.6151
R1341 B.n169 B.n168 10.6151
R1342 B.n172 B.n169 10.6151
R1343 B.n173 B.n172 10.6151
R1344 B.n176 B.n173 10.6151
R1345 B.n177 B.n176 10.6151
R1346 B.n180 B.n177 10.6151
R1347 B.n181 B.n180 10.6151
R1348 B.n184 B.n181 10.6151
R1349 B.n185 B.n184 10.6151
R1350 B.n188 B.n185 10.6151
R1351 B.n189 B.n188 10.6151
R1352 B.n192 B.n189 10.6151
R1353 B.n193 B.n192 10.6151
R1354 B.n196 B.n193 10.6151
R1355 B.n197 B.n196 10.6151
R1356 B.n200 B.n197 10.6151
R1357 B.n201 B.n200 10.6151
R1358 B.n204 B.n201 10.6151
R1359 B.n205 B.n204 10.6151
R1360 B.n208 B.n205 10.6151
R1361 B.n213 B.n210 10.6151
R1362 B.n214 B.n213 10.6151
R1363 B.n217 B.n214 10.6151
R1364 B.n218 B.n217 10.6151
R1365 B.n221 B.n218 10.6151
R1366 B.n222 B.n221 10.6151
R1367 B.n225 B.n222 10.6151
R1368 B.n226 B.n225 10.6151
R1369 B.n230 B.n229 10.6151
R1370 B.n233 B.n230 10.6151
R1371 B.n234 B.n233 10.6151
R1372 B.n237 B.n234 10.6151
R1373 B.n238 B.n237 10.6151
R1374 B.n241 B.n238 10.6151
R1375 B.n242 B.n241 10.6151
R1376 B.n245 B.n242 10.6151
R1377 B.n246 B.n245 10.6151
R1378 B.n249 B.n246 10.6151
R1379 B.n250 B.n249 10.6151
R1380 B.n253 B.n250 10.6151
R1381 B.n254 B.n253 10.6151
R1382 B.n257 B.n254 10.6151
R1383 B.n258 B.n257 10.6151
R1384 B.n261 B.n258 10.6151
R1385 B.n262 B.n261 10.6151
R1386 B.n265 B.n262 10.6151
R1387 B.n266 B.n265 10.6151
R1388 B.n269 B.n266 10.6151
R1389 B.n270 B.n269 10.6151
R1390 B.n273 B.n270 10.6151
R1391 B.n274 B.n273 10.6151
R1392 B.n277 B.n274 10.6151
R1393 B.n278 B.n277 10.6151
R1394 B.n281 B.n278 10.6151
R1395 B.n282 B.n281 10.6151
R1396 B.n285 B.n282 10.6151
R1397 B.n286 B.n285 10.6151
R1398 B.n289 B.n286 10.6151
R1399 B.n290 B.n289 10.6151
R1400 B.n293 B.n290 10.6151
R1401 B.n294 B.n293 10.6151
R1402 B.n297 B.n294 10.6151
R1403 B.n298 B.n297 10.6151
R1404 B.n301 B.n298 10.6151
R1405 B.n302 B.n301 10.6151
R1406 B.n305 B.n302 10.6151
R1407 B.n306 B.n305 10.6151
R1408 B.n309 B.n306 10.6151
R1409 B.n310 B.n309 10.6151
R1410 B.n313 B.n310 10.6151
R1411 B.n314 B.n313 10.6151
R1412 B.n317 B.n314 10.6151
R1413 B.n318 B.n317 10.6151
R1414 B.n776 B.n318 10.6151
R1415 B.n847 B.n0 8.11757
R1416 B.n847 B.n1 8.11757
R1417 B.n548 B.n434 6.5566
R1418 B.n532 B.n531 6.5566
R1419 B.n210 B.n209 6.5566
R1420 B.n226 B.n116 6.5566
R1421 B.n551 B.n434 4.05904
R1422 B.n531 B.n530 4.05904
R1423 B.n209 B.n208 4.05904
R1424 B.n229 B.n116 4.05904
R1425 B.n345 B.t16 2.90517
R1426 B.t1 B.n818 2.90517
R1427 B.t17 B.n325 1.7433
R1428 B.n834 B.t0 1.7433
R1429 B.n664 B.t3 0.581435
R1430 B.n795 B.t7 0.581435
R1431 VN.n0 VN.t1 176.812
R1432 VN.n1 VN.t3 176.812
R1433 VN.n0 VN.t0 176.15
R1434 VN.n1 VN.t2 176.15
R1435 VN VN.n1 52.5283
R1436 VN VN.n0 5.41845
R1437 VTAIL.n5 VTAIL.t0 47.7772
R1438 VTAIL.n4 VTAIL.t7 47.7772
R1439 VTAIL.n3 VTAIL.t5 47.7772
R1440 VTAIL.n7 VTAIL.t6 47.777
R1441 VTAIL.n0 VTAIL.t4 47.777
R1442 VTAIL.n1 VTAIL.t3 47.777
R1443 VTAIL.n2 VTAIL.t2 47.777
R1444 VTAIL.n6 VTAIL.t1 47.777
R1445 VTAIL.n7 VTAIL.n6 26.4531
R1446 VTAIL.n3 VTAIL.n2 26.4531
R1447 VTAIL.n4 VTAIL.n3 2.31084
R1448 VTAIL.n6 VTAIL.n5 2.31084
R1449 VTAIL.n2 VTAIL.n1 2.31084
R1450 VTAIL VTAIL.n0 1.21386
R1451 VTAIL VTAIL.n7 1.09748
R1452 VTAIL.n5 VTAIL.n4 0.470328
R1453 VTAIL.n1 VTAIL.n0 0.470328
R1454 VDD2.n2 VDD2.n0 105.428
R1455 VDD2.n2 VDD2.n1 63.0063
R1456 VDD2.n1 VDD2.t1 1.44999
R1457 VDD2.n1 VDD2.t0 1.44999
R1458 VDD2.n0 VDD2.t2 1.44999
R1459 VDD2.n0 VDD2.t3 1.44999
R1460 VDD2 VDD2.n2 0.0586897
R1461 VP.n3 VP.t3 176.812
R1462 VP.n3 VP.t0 176.15
R1463 VP.n12 VP.n0 161.3
R1464 VP.n11 VP.n10 161.3
R1465 VP.n9 VP.n1 161.3
R1466 VP.n8 VP.n7 161.3
R1467 VP.n6 VP.n2 161.3
R1468 VP.n5 VP.t2 140.089
R1469 VP.n13 VP.t1 140.089
R1470 VP.n5 VP.n4 94.1858
R1471 VP.n14 VP.n13 94.1858
R1472 VP.n4 VP.n3 52.2495
R1473 VP.n7 VP.n1 40.577
R1474 VP.n11 VP.n1 40.577
R1475 VP.n7 VP.n6 24.5923
R1476 VP.n12 VP.n11 24.5923
R1477 VP.n6 VP.n5 16.7229
R1478 VP.n13 VP.n12 16.7229
R1479 VP.n4 VP.n2 0.278335
R1480 VP.n14 VP.n0 0.278335
R1481 VP.n8 VP.n2 0.189894
R1482 VP.n9 VP.n8 0.189894
R1483 VP.n10 VP.n9 0.189894
R1484 VP.n10 VP.n0 0.189894
R1485 VP VP.n14 0.153485
R1486 VDD1 VDD1.n1 105.953
R1487 VDD1 VDD1.n0 63.0645
R1488 VDD1.n0 VDD1.t0 1.44999
R1489 VDD1.n0 VDD1.t3 1.44999
R1490 VDD1.n1 VDD1.t1 1.44999
R1491 VDD1.n1 VDD1.t2 1.44999
C0 VN VDD2 5.26684f
C1 VP VDD2 0.378562f
C2 VDD1 VTAIL 5.78892f
C3 VP VN 6.31257f
C4 VDD1 VDD2 0.969641f
C5 VTAIL VDD2 5.84145f
C6 VDD1 VN 0.148939f
C7 VDD1 VP 5.49579f
C8 VN VTAIL 5.06522f
C9 VP VTAIL 5.07933f
C10 VDD2 B 3.744837f
C11 VDD1 B 7.97347f
C12 VTAIL B 10.925116f
C13 VN B 10.37064f
C14 VP B 8.514333f
C15 VDD1.t0 B 0.290319f
C16 VDD1.t3 B 0.290319f
C17 VDD1.n0 B 2.615f
C18 VDD1.t1 B 0.290319f
C19 VDD1.t2 B 0.290319f
C20 VDD1.n1 B 3.35233f
C21 VP.n0 B 0.035802f
C22 VP.t1 B 2.38351f
C23 VP.n1 B 0.021934f
C24 VP.n2 B 0.035802f
C25 VP.t2 B 2.38351f
C26 VP.t0 B 2.58813f
C27 VP.t3 B 2.59181f
C28 VP.n3 B 3.09993f
C29 VP.n4 B 1.55106f
C30 VP.n5 B 0.9309f
C31 VP.n6 B 0.042405f
C32 VP.n7 B 0.053691f
C33 VP.n8 B 0.027157f
C34 VP.n9 B 0.027157f
C35 VP.n10 B 0.027157f
C36 VP.n11 B 0.053691f
C37 VP.n12 B 0.042405f
C38 VP.n13 B 0.9309f
C39 VP.n14 B 0.037296f
C40 VDD2.t2 B 0.28771f
C41 VDD2.t3 B 0.28771f
C42 VDD2.n0 B 3.29555f
C43 VDD2.t1 B 0.28771f
C44 VDD2.t0 B 0.28771f
C45 VDD2.n1 B 2.5911f
C46 VDD2.n2 B 3.85835f
C47 VTAIL.t4 B 1.91837f
C48 VTAIL.n0 B 0.292556f
C49 VTAIL.t3 B 1.91837f
C50 VTAIL.n1 B 0.348876f
C51 VTAIL.t2 B 1.91837f
C52 VTAIL.n2 B 1.26439f
C53 VTAIL.t5 B 1.91837f
C54 VTAIL.n3 B 1.26439f
C55 VTAIL.t7 B 1.91837f
C56 VTAIL.n4 B 0.348874f
C57 VTAIL.t0 B 1.91837f
C58 VTAIL.n5 B 0.348874f
C59 VTAIL.t1 B 1.91837f
C60 VTAIL.n6 B 1.26439f
C61 VTAIL.t6 B 1.91837f
C62 VTAIL.n7 B 1.2021f
C63 VN.t1 B 2.55537f
C64 VN.t0 B 2.55174f
C65 VN.n0 B 1.65818f
C66 VN.t3 B 2.55537f
C67 VN.t2 B 2.55174f
C68 VN.n1 B 3.07025f
.ends

