* NGSPICE file created from diff_pair_sample_0949.ext - technology: sky130A

.subckt diff_pair_sample_0949 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5311 pd=15.67 as=5.9826 ps=31.46 w=15.34 l=3.7
X1 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5311 pd=15.67 as=5.9826 ps=31.46 w=15.34 l=3.7
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.7
X3 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=2.5311 ps=15.67 w=15.34 l=3.7
X4 VTAIL.t4 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=2.5311 ps=15.67 w=15.34 l=3.7
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.7
X6 VTAIL.t6 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=2.5311 ps=15.67 w=15.34 l=3.7
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.7
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=0 ps=0 w=15.34 l=3.7
X9 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5311 pd=15.67 as=5.9826 ps=31.46 w=15.34 l=3.7
X10 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9826 pd=31.46 as=2.5311 ps=15.67 w=15.34 l=3.7
X11 VDD1.t0 VP.t3 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5311 pd=15.67 as=5.9826 ps=31.46 w=15.34 l=3.7
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n5 VP.t1 133.264
R10 VP.n5 VP.t0 131.939
R11 VP.n7 VP.t2 99.9178
R12 VP.n0 VP.t3 99.9178
R13 VP.n7 VP.n6 89.5078
R14 VP.n22 VP.n0 89.5078
R15 VP.n6 VP.n5 54.1237
R16 VP.n14 VP.n13 40.577
R17 VP.n14 VP.n2 40.577
R18 VP.n8 VP.n4 24.5923
R19 VP.n12 VP.n4 24.5923
R20 VP.n13 VP.n12 24.5923
R21 VP.n18 VP.n2 24.5923
R22 VP.n19 VP.n18 24.5923
R23 VP.n20 VP.n19 24.5923
R24 VP.n8 VP.n7 0.738255
R25 VP.n20 VP.n0 0.738255
R26 VP.n9 VP.n6 0.354861
R27 VP.n22 VP.n21 0.354861
R28 VP VP.n22 0.267071
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VTAIL.n682 VTAIL.n602 289.615
R38 VTAIL.n80 VTAIL.n0 289.615
R39 VTAIL.n166 VTAIL.n86 289.615
R40 VTAIL.n252 VTAIL.n172 289.615
R41 VTAIL.n596 VTAIL.n516 289.615
R42 VTAIL.n510 VTAIL.n430 289.615
R43 VTAIL.n424 VTAIL.n344 289.615
R44 VTAIL.n338 VTAIL.n258 289.615
R45 VTAIL.n631 VTAIL.n630 185
R46 VTAIL.n633 VTAIL.n632 185
R47 VTAIL.n626 VTAIL.n625 185
R48 VTAIL.n639 VTAIL.n638 185
R49 VTAIL.n641 VTAIL.n640 185
R50 VTAIL.n622 VTAIL.n621 185
R51 VTAIL.n647 VTAIL.n646 185
R52 VTAIL.n649 VTAIL.n648 185
R53 VTAIL.n618 VTAIL.n617 185
R54 VTAIL.n655 VTAIL.n654 185
R55 VTAIL.n657 VTAIL.n656 185
R56 VTAIL.n614 VTAIL.n613 185
R57 VTAIL.n663 VTAIL.n662 185
R58 VTAIL.n665 VTAIL.n664 185
R59 VTAIL.n610 VTAIL.n609 185
R60 VTAIL.n672 VTAIL.n671 185
R61 VTAIL.n673 VTAIL.n608 185
R62 VTAIL.n675 VTAIL.n674 185
R63 VTAIL.n606 VTAIL.n605 185
R64 VTAIL.n681 VTAIL.n680 185
R65 VTAIL.n683 VTAIL.n682 185
R66 VTAIL.n29 VTAIL.n28 185
R67 VTAIL.n31 VTAIL.n30 185
R68 VTAIL.n24 VTAIL.n23 185
R69 VTAIL.n37 VTAIL.n36 185
R70 VTAIL.n39 VTAIL.n38 185
R71 VTAIL.n20 VTAIL.n19 185
R72 VTAIL.n45 VTAIL.n44 185
R73 VTAIL.n47 VTAIL.n46 185
R74 VTAIL.n16 VTAIL.n15 185
R75 VTAIL.n53 VTAIL.n52 185
R76 VTAIL.n55 VTAIL.n54 185
R77 VTAIL.n12 VTAIL.n11 185
R78 VTAIL.n61 VTAIL.n60 185
R79 VTAIL.n63 VTAIL.n62 185
R80 VTAIL.n8 VTAIL.n7 185
R81 VTAIL.n70 VTAIL.n69 185
R82 VTAIL.n71 VTAIL.n6 185
R83 VTAIL.n73 VTAIL.n72 185
R84 VTAIL.n4 VTAIL.n3 185
R85 VTAIL.n79 VTAIL.n78 185
R86 VTAIL.n81 VTAIL.n80 185
R87 VTAIL.n115 VTAIL.n114 185
R88 VTAIL.n117 VTAIL.n116 185
R89 VTAIL.n110 VTAIL.n109 185
R90 VTAIL.n123 VTAIL.n122 185
R91 VTAIL.n125 VTAIL.n124 185
R92 VTAIL.n106 VTAIL.n105 185
R93 VTAIL.n131 VTAIL.n130 185
R94 VTAIL.n133 VTAIL.n132 185
R95 VTAIL.n102 VTAIL.n101 185
R96 VTAIL.n139 VTAIL.n138 185
R97 VTAIL.n141 VTAIL.n140 185
R98 VTAIL.n98 VTAIL.n97 185
R99 VTAIL.n147 VTAIL.n146 185
R100 VTAIL.n149 VTAIL.n148 185
R101 VTAIL.n94 VTAIL.n93 185
R102 VTAIL.n156 VTAIL.n155 185
R103 VTAIL.n157 VTAIL.n92 185
R104 VTAIL.n159 VTAIL.n158 185
R105 VTAIL.n90 VTAIL.n89 185
R106 VTAIL.n165 VTAIL.n164 185
R107 VTAIL.n167 VTAIL.n166 185
R108 VTAIL.n201 VTAIL.n200 185
R109 VTAIL.n203 VTAIL.n202 185
R110 VTAIL.n196 VTAIL.n195 185
R111 VTAIL.n209 VTAIL.n208 185
R112 VTAIL.n211 VTAIL.n210 185
R113 VTAIL.n192 VTAIL.n191 185
R114 VTAIL.n217 VTAIL.n216 185
R115 VTAIL.n219 VTAIL.n218 185
R116 VTAIL.n188 VTAIL.n187 185
R117 VTAIL.n225 VTAIL.n224 185
R118 VTAIL.n227 VTAIL.n226 185
R119 VTAIL.n184 VTAIL.n183 185
R120 VTAIL.n233 VTAIL.n232 185
R121 VTAIL.n235 VTAIL.n234 185
R122 VTAIL.n180 VTAIL.n179 185
R123 VTAIL.n242 VTAIL.n241 185
R124 VTAIL.n243 VTAIL.n178 185
R125 VTAIL.n245 VTAIL.n244 185
R126 VTAIL.n176 VTAIL.n175 185
R127 VTAIL.n251 VTAIL.n250 185
R128 VTAIL.n253 VTAIL.n252 185
R129 VTAIL.n597 VTAIL.n596 185
R130 VTAIL.n595 VTAIL.n594 185
R131 VTAIL.n520 VTAIL.n519 185
R132 VTAIL.n524 VTAIL.n522 185
R133 VTAIL.n589 VTAIL.n588 185
R134 VTAIL.n587 VTAIL.n586 185
R135 VTAIL.n526 VTAIL.n525 185
R136 VTAIL.n581 VTAIL.n580 185
R137 VTAIL.n579 VTAIL.n578 185
R138 VTAIL.n530 VTAIL.n529 185
R139 VTAIL.n573 VTAIL.n572 185
R140 VTAIL.n571 VTAIL.n570 185
R141 VTAIL.n534 VTAIL.n533 185
R142 VTAIL.n565 VTAIL.n564 185
R143 VTAIL.n563 VTAIL.n562 185
R144 VTAIL.n538 VTAIL.n537 185
R145 VTAIL.n557 VTAIL.n556 185
R146 VTAIL.n555 VTAIL.n554 185
R147 VTAIL.n542 VTAIL.n541 185
R148 VTAIL.n549 VTAIL.n548 185
R149 VTAIL.n547 VTAIL.n546 185
R150 VTAIL.n511 VTAIL.n510 185
R151 VTAIL.n509 VTAIL.n508 185
R152 VTAIL.n434 VTAIL.n433 185
R153 VTAIL.n438 VTAIL.n436 185
R154 VTAIL.n503 VTAIL.n502 185
R155 VTAIL.n501 VTAIL.n500 185
R156 VTAIL.n440 VTAIL.n439 185
R157 VTAIL.n495 VTAIL.n494 185
R158 VTAIL.n493 VTAIL.n492 185
R159 VTAIL.n444 VTAIL.n443 185
R160 VTAIL.n487 VTAIL.n486 185
R161 VTAIL.n485 VTAIL.n484 185
R162 VTAIL.n448 VTAIL.n447 185
R163 VTAIL.n479 VTAIL.n478 185
R164 VTAIL.n477 VTAIL.n476 185
R165 VTAIL.n452 VTAIL.n451 185
R166 VTAIL.n471 VTAIL.n470 185
R167 VTAIL.n469 VTAIL.n468 185
R168 VTAIL.n456 VTAIL.n455 185
R169 VTAIL.n463 VTAIL.n462 185
R170 VTAIL.n461 VTAIL.n460 185
R171 VTAIL.n425 VTAIL.n424 185
R172 VTAIL.n423 VTAIL.n422 185
R173 VTAIL.n348 VTAIL.n347 185
R174 VTAIL.n352 VTAIL.n350 185
R175 VTAIL.n417 VTAIL.n416 185
R176 VTAIL.n415 VTAIL.n414 185
R177 VTAIL.n354 VTAIL.n353 185
R178 VTAIL.n409 VTAIL.n408 185
R179 VTAIL.n407 VTAIL.n406 185
R180 VTAIL.n358 VTAIL.n357 185
R181 VTAIL.n401 VTAIL.n400 185
R182 VTAIL.n399 VTAIL.n398 185
R183 VTAIL.n362 VTAIL.n361 185
R184 VTAIL.n393 VTAIL.n392 185
R185 VTAIL.n391 VTAIL.n390 185
R186 VTAIL.n366 VTAIL.n365 185
R187 VTAIL.n385 VTAIL.n384 185
R188 VTAIL.n383 VTAIL.n382 185
R189 VTAIL.n370 VTAIL.n369 185
R190 VTAIL.n377 VTAIL.n376 185
R191 VTAIL.n375 VTAIL.n374 185
R192 VTAIL.n339 VTAIL.n338 185
R193 VTAIL.n337 VTAIL.n336 185
R194 VTAIL.n262 VTAIL.n261 185
R195 VTAIL.n266 VTAIL.n264 185
R196 VTAIL.n331 VTAIL.n330 185
R197 VTAIL.n329 VTAIL.n328 185
R198 VTAIL.n268 VTAIL.n267 185
R199 VTAIL.n323 VTAIL.n322 185
R200 VTAIL.n321 VTAIL.n320 185
R201 VTAIL.n272 VTAIL.n271 185
R202 VTAIL.n315 VTAIL.n314 185
R203 VTAIL.n313 VTAIL.n312 185
R204 VTAIL.n276 VTAIL.n275 185
R205 VTAIL.n307 VTAIL.n306 185
R206 VTAIL.n305 VTAIL.n304 185
R207 VTAIL.n280 VTAIL.n279 185
R208 VTAIL.n299 VTAIL.n298 185
R209 VTAIL.n297 VTAIL.n296 185
R210 VTAIL.n284 VTAIL.n283 185
R211 VTAIL.n291 VTAIL.n290 185
R212 VTAIL.n289 VTAIL.n288 185
R213 VTAIL.n629 VTAIL.t0 147.659
R214 VTAIL.n27 VTAIL.t3 147.659
R215 VTAIL.n113 VTAIL.t5 147.659
R216 VTAIL.n199 VTAIL.t6 147.659
R217 VTAIL.n545 VTAIL.t7 147.659
R218 VTAIL.n459 VTAIL.t4 147.659
R219 VTAIL.n373 VTAIL.t2 147.659
R220 VTAIL.n287 VTAIL.t1 147.659
R221 VTAIL.n632 VTAIL.n631 104.615
R222 VTAIL.n632 VTAIL.n625 104.615
R223 VTAIL.n639 VTAIL.n625 104.615
R224 VTAIL.n640 VTAIL.n639 104.615
R225 VTAIL.n640 VTAIL.n621 104.615
R226 VTAIL.n647 VTAIL.n621 104.615
R227 VTAIL.n648 VTAIL.n647 104.615
R228 VTAIL.n648 VTAIL.n617 104.615
R229 VTAIL.n655 VTAIL.n617 104.615
R230 VTAIL.n656 VTAIL.n655 104.615
R231 VTAIL.n656 VTAIL.n613 104.615
R232 VTAIL.n663 VTAIL.n613 104.615
R233 VTAIL.n664 VTAIL.n663 104.615
R234 VTAIL.n664 VTAIL.n609 104.615
R235 VTAIL.n672 VTAIL.n609 104.615
R236 VTAIL.n673 VTAIL.n672 104.615
R237 VTAIL.n674 VTAIL.n673 104.615
R238 VTAIL.n674 VTAIL.n605 104.615
R239 VTAIL.n681 VTAIL.n605 104.615
R240 VTAIL.n682 VTAIL.n681 104.615
R241 VTAIL.n30 VTAIL.n29 104.615
R242 VTAIL.n30 VTAIL.n23 104.615
R243 VTAIL.n37 VTAIL.n23 104.615
R244 VTAIL.n38 VTAIL.n37 104.615
R245 VTAIL.n38 VTAIL.n19 104.615
R246 VTAIL.n45 VTAIL.n19 104.615
R247 VTAIL.n46 VTAIL.n45 104.615
R248 VTAIL.n46 VTAIL.n15 104.615
R249 VTAIL.n53 VTAIL.n15 104.615
R250 VTAIL.n54 VTAIL.n53 104.615
R251 VTAIL.n54 VTAIL.n11 104.615
R252 VTAIL.n61 VTAIL.n11 104.615
R253 VTAIL.n62 VTAIL.n61 104.615
R254 VTAIL.n62 VTAIL.n7 104.615
R255 VTAIL.n70 VTAIL.n7 104.615
R256 VTAIL.n71 VTAIL.n70 104.615
R257 VTAIL.n72 VTAIL.n71 104.615
R258 VTAIL.n72 VTAIL.n3 104.615
R259 VTAIL.n79 VTAIL.n3 104.615
R260 VTAIL.n80 VTAIL.n79 104.615
R261 VTAIL.n116 VTAIL.n115 104.615
R262 VTAIL.n116 VTAIL.n109 104.615
R263 VTAIL.n123 VTAIL.n109 104.615
R264 VTAIL.n124 VTAIL.n123 104.615
R265 VTAIL.n124 VTAIL.n105 104.615
R266 VTAIL.n131 VTAIL.n105 104.615
R267 VTAIL.n132 VTAIL.n131 104.615
R268 VTAIL.n132 VTAIL.n101 104.615
R269 VTAIL.n139 VTAIL.n101 104.615
R270 VTAIL.n140 VTAIL.n139 104.615
R271 VTAIL.n140 VTAIL.n97 104.615
R272 VTAIL.n147 VTAIL.n97 104.615
R273 VTAIL.n148 VTAIL.n147 104.615
R274 VTAIL.n148 VTAIL.n93 104.615
R275 VTAIL.n156 VTAIL.n93 104.615
R276 VTAIL.n157 VTAIL.n156 104.615
R277 VTAIL.n158 VTAIL.n157 104.615
R278 VTAIL.n158 VTAIL.n89 104.615
R279 VTAIL.n165 VTAIL.n89 104.615
R280 VTAIL.n166 VTAIL.n165 104.615
R281 VTAIL.n202 VTAIL.n201 104.615
R282 VTAIL.n202 VTAIL.n195 104.615
R283 VTAIL.n209 VTAIL.n195 104.615
R284 VTAIL.n210 VTAIL.n209 104.615
R285 VTAIL.n210 VTAIL.n191 104.615
R286 VTAIL.n217 VTAIL.n191 104.615
R287 VTAIL.n218 VTAIL.n217 104.615
R288 VTAIL.n218 VTAIL.n187 104.615
R289 VTAIL.n225 VTAIL.n187 104.615
R290 VTAIL.n226 VTAIL.n225 104.615
R291 VTAIL.n226 VTAIL.n183 104.615
R292 VTAIL.n233 VTAIL.n183 104.615
R293 VTAIL.n234 VTAIL.n233 104.615
R294 VTAIL.n234 VTAIL.n179 104.615
R295 VTAIL.n242 VTAIL.n179 104.615
R296 VTAIL.n243 VTAIL.n242 104.615
R297 VTAIL.n244 VTAIL.n243 104.615
R298 VTAIL.n244 VTAIL.n175 104.615
R299 VTAIL.n251 VTAIL.n175 104.615
R300 VTAIL.n252 VTAIL.n251 104.615
R301 VTAIL.n596 VTAIL.n595 104.615
R302 VTAIL.n595 VTAIL.n519 104.615
R303 VTAIL.n524 VTAIL.n519 104.615
R304 VTAIL.n588 VTAIL.n524 104.615
R305 VTAIL.n588 VTAIL.n587 104.615
R306 VTAIL.n587 VTAIL.n525 104.615
R307 VTAIL.n580 VTAIL.n525 104.615
R308 VTAIL.n580 VTAIL.n579 104.615
R309 VTAIL.n579 VTAIL.n529 104.615
R310 VTAIL.n572 VTAIL.n529 104.615
R311 VTAIL.n572 VTAIL.n571 104.615
R312 VTAIL.n571 VTAIL.n533 104.615
R313 VTAIL.n564 VTAIL.n533 104.615
R314 VTAIL.n564 VTAIL.n563 104.615
R315 VTAIL.n563 VTAIL.n537 104.615
R316 VTAIL.n556 VTAIL.n537 104.615
R317 VTAIL.n556 VTAIL.n555 104.615
R318 VTAIL.n555 VTAIL.n541 104.615
R319 VTAIL.n548 VTAIL.n541 104.615
R320 VTAIL.n548 VTAIL.n547 104.615
R321 VTAIL.n510 VTAIL.n509 104.615
R322 VTAIL.n509 VTAIL.n433 104.615
R323 VTAIL.n438 VTAIL.n433 104.615
R324 VTAIL.n502 VTAIL.n438 104.615
R325 VTAIL.n502 VTAIL.n501 104.615
R326 VTAIL.n501 VTAIL.n439 104.615
R327 VTAIL.n494 VTAIL.n439 104.615
R328 VTAIL.n494 VTAIL.n493 104.615
R329 VTAIL.n493 VTAIL.n443 104.615
R330 VTAIL.n486 VTAIL.n443 104.615
R331 VTAIL.n486 VTAIL.n485 104.615
R332 VTAIL.n485 VTAIL.n447 104.615
R333 VTAIL.n478 VTAIL.n447 104.615
R334 VTAIL.n478 VTAIL.n477 104.615
R335 VTAIL.n477 VTAIL.n451 104.615
R336 VTAIL.n470 VTAIL.n451 104.615
R337 VTAIL.n470 VTAIL.n469 104.615
R338 VTAIL.n469 VTAIL.n455 104.615
R339 VTAIL.n462 VTAIL.n455 104.615
R340 VTAIL.n462 VTAIL.n461 104.615
R341 VTAIL.n424 VTAIL.n423 104.615
R342 VTAIL.n423 VTAIL.n347 104.615
R343 VTAIL.n352 VTAIL.n347 104.615
R344 VTAIL.n416 VTAIL.n352 104.615
R345 VTAIL.n416 VTAIL.n415 104.615
R346 VTAIL.n415 VTAIL.n353 104.615
R347 VTAIL.n408 VTAIL.n353 104.615
R348 VTAIL.n408 VTAIL.n407 104.615
R349 VTAIL.n407 VTAIL.n357 104.615
R350 VTAIL.n400 VTAIL.n357 104.615
R351 VTAIL.n400 VTAIL.n399 104.615
R352 VTAIL.n399 VTAIL.n361 104.615
R353 VTAIL.n392 VTAIL.n361 104.615
R354 VTAIL.n392 VTAIL.n391 104.615
R355 VTAIL.n391 VTAIL.n365 104.615
R356 VTAIL.n384 VTAIL.n365 104.615
R357 VTAIL.n384 VTAIL.n383 104.615
R358 VTAIL.n383 VTAIL.n369 104.615
R359 VTAIL.n376 VTAIL.n369 104.615
R360 VTAIL.n376 VTAIL.n375 104.615
R361 VTAIL.n338 VTAIL.n337 104.615
R362 VTAIL.n337 VTAIL.n261 104.615
R363 VTAIL.n266 VTAIL.n261 104.615
R364 VTAIL.n330 VTAIL.n266 104.615
R365 VTAIL.n330 VTAIL.n329 104.615
R366 VTAIL.n329 VTAIL.n267 104.615
R367 VTAIL.n322 VTAIL.n267 104.615
R368 VTAIL.n322 VTAIL.n321 104.615
R369 VTAIL.n321 VTAIL.n271 104.615
R370 VTAIL.n314 VTAIL.n271 104.615
R371 VTAIL.n314 VTAIL.n313 104.615
R372 VTAIL.n313 VTAIL.n275 104.615
R373 VTAIL.n306 VTAIL.n275 104.615
R374 VTAIL.n306 VTAIL.n305 104.615
R375 VTAIL.n305 VTAIL.n279 104.615
R376 VTAIL.n298 VTAIL.n279 104.615
R377 VTAIL.n298 VTAIL.n297 104.615
R378 VTAIL.n297 VTAIL.n283 104.615
R379 VTAIL.n290 VTAIL.n283 104.615
R380 VTAIL.n290 VTAIL.n289 104.615
R381 VTAIL.n631 VTAIL.t0 52.3082
R382 VTAIL.n29 VTAIL.t3 52.3082
R383 VTAIL.n115 VTAIL.t5 52.3082
R384 VTAIL.n201 VTAIL.t6 52.3082
R385 VTAIL.n547 VTAIL.t7 52.3082
R386 VTAIL.n461 VTAIL.t4 52.3082
R387 VTAIL.n375 VTAIL.t2 52.3082
R388 VTAIL.n289 VTAIL.t1 52.3082
R389 VTAIL.n687 VTAIL.n686 31.7975
R390 VTAIL.n85 VTAIL.n84 31.7975
R391 VTAIL.n171 VTAIL.n170 31.7975
R392 VTAIL.n257 VTAIL.n256 31.7975
R393 VTAIL.n601 VTAIL.n600 31.7975
R394 VTAIL.n515 VTAIL.n514 31.7975
R395 VTAIL.n429 VTAIL.n428 31.7975
R396 VTAIL.n343 VTAIL.n342 31.7975
R397 VTAIL.n687 VTAIL.n601 29.0652
R398 VTAIL.n343 VTAIL.n257 29.0652
R399 VTAIL.n630 VTAIL.n629 15.6677
R400 VTAIL.n28 VTAIL.n27 15.6677
R401 VTAIL.n114 VTAIL.n113 15.6677
R402 VTAIL.n200 VTAIL.n199 15.6677
R403 VTAIL.n546 VTAIL.n545 15.6677
R404 VTAIL.n460 VTAIL.n459 15.6677
R405 VTAIL.n374 VTAIL.n373 15.6677
R406 VTAIL.n288 VTAIL.n287 15.6677
R407 VTAIL.n675 VTAIL.n606 13.1884
R408 VTAIL.n73 VTAIL.n4 13.1884
R409 VTAIL.n159 VTAIL.n90 13.1884
R410 VTAIL.n245 VTAIL.n176 13.1884
R411 VTAIL.n522 VTAIL.n520 13.1884
R412 VTAIL.n436 VTAIL.n434 13.1884
R413 VTAIL.n350 VTAIL.n348 13.1884
R414 VTAIL.n264 VTAIL.n262 13.1884
R415 VTAIL.n633 VTAIL.n628 12.8005
R416 VTAIL.n676 VTAIL.n608 12.8005
R417 VTAIL.n680 VTAIL.n679 12.8005
R418 VTAIL.n31 VTAIL.n26 12.8005
R419 VTAIL.n74 VTAIL.n6 12.8005
R420 VTAIL.n78 VTAIL.n77 12.8005
R421 VTAIL.n117 VTAIL.n112 12.8005
R422 VTAIL.n160 VTAIL.n92 12.8005
R423 VTAIL.n164 VTAIL.n163 12.8005
R424 VTAIL.n203 VTAIL.n198 12.8005
R425 VTAIL.n246 VTAIL.n178 12.8005
R426 VTAIL.n250 VTAIL.n249 12.8005
R427 VTAIL.n594 VTAIL.n593 12.8005
R428 VTAIL.n590 VTAIL.n589 12.8005
R429 VTAIL.n549 VTAIL.n544 12.8005
R430 VTAIL.n508 VTAIL.n507 12.8005
R431 VTAIL.n504 VTAIL.n503 12.8005
R432 VTAIL.n463 VTAIL.n458 12.8005
R433 VTAIL.n422 VTAIL.n421 12.8005
R434 VTAIL.n418 VTAIL.n417 12.8005
R435 VTAIL.n377 VTAIL.n372 12.8005
R436 VTAIL.n336 VTAIL.n335 12.8005
R437 VTAIL.n332 VTAIL.n331 12.8005
R438 VTAIL.n291 VTAIL.n286 12.8005
R439 VTAIL.n634 VTAIL.n626 12.0247
R440 VTAIL.n671 VTAIL.n670 12.0247
R441 VTAIL.n683 VTAIL.n604 12.0247
R442 VTAIL.n32 VTAIL.n24 12.0247
R443 VTAIL.n69 VTAIL.n68 12.0247
R444 VTAIL.n81 VTAIL.n2 12.0247
R445 VTAIL.n118 VTAIL.n110 12.0247
R446 VTAIL.n155 VTAIL.n154 12.0247
R447 VTAIL.n167 VTAIL.n88 12.0247
R448 VTAIL.n204 VTAIL.n196 12.0247
R449 VTAIL.n241 VTAIL.n240 12.0247
R450 VTAIL.n253 VTAIL.n174 12.0247
R451 VTAIL.n597 VTAIL.n518 12.0247
R452 VTAIL.n586 VTAIL.n523 12.0247
R453 VTAIL.n550 VTAIL.n542 12.0247
R454 VTAIL.n511 VTAIL.n432 12.0247
R455 VTAIL.n500 VTAIL.n437 12.0247
R456 VTAIL.n464 VTAIL.n456 12.0247
R457 VTAIL.n425 VTAIL.n346 12.0247
R458 VTAIL.n414 VTAIL.n351 12.0247
R459 VTAIL.n378 VTAIL.n370 12.0247
R460 VTAIL.n339 VTAIL.n260 12.0247
R461 VTAIL.n328 VTAIL.n265 12.0247
R462 VTAIL.n292 VTAIL.n284 12.0247
R463 VTAIL.n638 VTAIL.n637 11.249
R464 VTAIL.n669 VTAIL.n610 11.249
R465 VTAIL.n684 VTAIL.n602 11.249
R466 VTAIL.n36 VTAIL.n35 11.249
R467 VTAIL.n67 VTAIL.n8 11.249
R468 VTAIL.n82 VTAIL.n0 11.249
R469 VTAIL.n122 VTAIL.n121 11.249
R470 VTAIL.n153 VTAIL.n94 11.249
R471 VTAIL.n168 VTAIL.n86 11.249
R472 VTAIL.n208 VTAIL.n207 11.249
R473 VTAIL.n239 VTAIL.n180 11.249
R474 VTAIL.n254 VTAIL.n172 11.249
R475 VTAIL.n598 VTAIL.n516 11.249
R476 VTAIL.n585 VTAIL.n526 11.249
R477 VTAIL.n554 VTAIL.n553 11.249
R478 VTAIL.n512 VTAIL.n430 11.249
R479 VTAIL.n499 VTAIL.n440 11.249
R480 VTAIL.n468 VTAIL.n467 11.249
R481 VTAIL.n426 VTAIL.n344 11.249
R482 VTAIL.n413 VTAIL.n354 11.249
R483 VTAIL.n382 VTAIL.n381 11.249
R484 VTAIL.n340 VTAIL.n258 11.249
R485 VTAIL.n327 VTAIL.n268 11.249
R486 VTAIL.n296 VTAIL.n295 11.249
R487 VTAIL.n641 VTAIL.n624 10.4732
R488 VTAIL.n666 VTAIL.n665 10.4732
R489 VTAIL.n39 VTAIL.n22 10.4732
R490 VTAIL.n64 VTAIL.n63 10.4732
R491 VTAIL.n125 VTAIL.n108 10.4732
R492 VTAIL.n150 VTAIL.n149 10.4732
R493 VTAIL.n211 VTAIL.n194 10.4732
R494 VTAIL.n236 VTAIL.n235 10.4732
R495 VTAIL.n582 VTAIL.n581 10.4732
R496 VTAIL.n557 VTAIL.n540 10.4732
R497 VTAIL.n496 VTAIL.n495 10.4732
R498 VTAIL.n471 VTAIL.n454 10.4732
R499 VTAIL.n410 VTAIL.n409 10.4732
R500 VTAIL.n385 VTAIL.n368 10.4732
R501 VTAIL.n324 VTAIL.n323 10.4732
R502 VTAIL.n299 VTAIL.n282 10.4732
R503 VTAIL.n642 VTAIL.n622 9.69747
R504 VTAIL.n662 VTAIL.n612 9.69747
R505 VTAIL.n40 VTAIL.n20 9.69747
R506 VTAIL.n60 VTAIL.n10 9.69747
R507 VTAIL.n126 VTAIL.n106 9.69747
R508 VTAIL.n146 VTAIL.n96 9.69747
R509 VTAIL.n212 VTAIL.n192 9.69747
R510 VTAIL.n232 VTAIL.n182 9.69747
R511 VTAIL.n578 VTAIL.n528 9.69747
R512 VTAIL.n558 VTAIL.n538 9.69747
R513 VTAIL.n492 VTAIL.n442 9.69747
R514 VTAIL.n472 VTAIL.n452 9.69747
R515 VTAIL.n406 VTAIL.n356 9.69747
R516 VTAIL.n386 VTAIL.n366 9.69747
R517 VTAIL.n320 VTAIL.n270 9.69747
R518 VTAIL.n300 VTAIL.n280 9.69747
R519 VTAIL.n686 VTAIL.n685 9.45567
R520 VTAIL.n84 VTAIL.n83 9.45567
R521 VTAIL.n170 VTAIL.n169 9.45567
R522 VTAIL.n256 VTAIL.n255 9.45567
R523 VTAIL.n600 VTAIL.n599 9.45567
R524 VTAIL.n514 VTAIL.n513 9.45567
R525 VTAIL.n428 VTAIL.n427 9.45567
R526 VTAIL.n342 VTAIL.n341 9.45567
R527 VTAIL.n685 VTAIL.n684 9.3005
R528 VTAIL.n604 VTAIL.n603 9.3005
R529 VTAIL.n679 VTAIL.n678 9.3005
R530 VTAIL.n651 VTAIL.n650 9.3005
R531 VTAIL.n620 VTAIL.n619 9.3005
R532 VTAIL.n645 VTAIL.n644 9.3005
R533 VTAIL.n643 VTAIL.n642 9.3005
R534 VTAIL.n624 VTAIL.n623 9.3005
R535 VTAIL.n637 VTAIL.n636 9.3005
R536 VTAIL.n635 VTAIL.n634 9.3005
R537 VTAIL.n628 VTAIL.n627 9.3005
R538 VTAIL.n653 VTAIL.n652 9.3005
R539 VTAIL.n616 VTAIL.n615 9.3005
R540 VTAIL.n659 VTAIL.n658 9.3005
R541 VTAIL.n661 VTAIL.n660 9.3005
R542 VTAIL.n612 VTAIL.n611 9.3005
R543 VTAIL.n667 VTAIL.n666 9.3005
R544 VTAIL.n669 VTAIL.n668 9.3005
R545 VTAIL.n670 VTAIL.n607 9.3005
R546 VTAIL.n677 VTAIL.n676 9.3005
R547 VTAIL.n83 VTAIL.n82 9.3005
R548 VTAIL.n2 VTAIL.n1 9.3005
R549 VTAIL.n77 VTAIL.n76 9.3005
R550 VTAIL.n49 VTAIL.n48 9.3005
R551 VTAIL.n18 VTAIL.n17 9.3005
R552 VTAIL.n43 VTAIL.n42 9.3005
R553 VTAIL.n41 VTAIL.n40 9.3005
R554 VTAIL.n22 VTAIL.n21 9.3005
R555 VTAIL.n35 VTAIL.n34 9.3005
R556 VTAIL.n33 VTAIL.n32 9.3005
R557 VTAIL.n26 VTAIL.n25 9.3005
R558 VTAIL.n51 VTAIL.n50 9.3005
R559 VTAIL.n14 VTAIL.n13 9.3005
R560 VTAIL.n57 VTAIL.n56 9.3005
R561 VTAIL.n59 VTAIL.n58 9.3005
R562 VTAIL.n10 VTAIL.n9 9.3005
R563 VTAIL.n65 VTAIL.n64 9.3005
R564 VTAIL.n67 VTAIL.n66 9.3005
R565 VTAIL.n68 VTAIL.n5 9.3005
R566 VTAIL.n75 VTAIL.n74 9.3005
R567 VTAIL.n169 VTAIL.n168 9.3005
R568 VTAIL.n88 VTAIL.n87 9.3005
R569 VTAIL.n163 VTAIL.n162 9.3005
R570 VTAIL.n135 VTAIL.n134 9.3005
R571 VTAIL.n104 VTAIL.n103 9.3005
R572 VTAIL.n129 VTAIL.n128 9.3005
R573 VTAIL.n127 VTAIL.n126 9.3005
R574 VTAIL.n108 VTAIL.n107 9.3005
R575 VTAIL.n121 VTAIL.n120 9.3005
R576 VTAIL.n119 VTAIL.n118 9.3005
R577 VTAIL.n112 VTAIL.n111 9.3005
R578 VTAIL.n137 VTAIL.n136 9.3005
R579 VTAIL.n100 VTAIL.n99 9.3005
R580 VTAIL.n143 VTAIL.n142 9.3005
R581 VTAIL.n145 VTAIL.n144 9.3005
R582 VTAIL.n96 VTAIL.n95 9.3005
R583 VTAIL.n151 VTAIL.n150 9.3005
R584 VTAIL.n153 VTAIL.n152 9.3005
R585 VTAIL.n154 VTAIL.n91 9.3005
R586 VTAIL.n161 VTAIL.n160 9.3005
R587 VTAIL.n255 VTAIL.n254 9.3005
R588 VTAIL.n174 VTAIL.n173 9.3005
R589 VTAIL.n249 VTAIL.n248 9.3005
R590 VTAIL.n221 VTAIL.n220 9.3005
R591 VTAIL.n190 VTAIL.n189 9.3005
R592 VTAIL.n215 VTAIL.n214 9.3005
R593 VTAIL.n213 VTAIL.n212 9.3005
R594 VTAIL.n194 VTAIL.n193 9.3005
R595 VTAIL.n207 VTAIL.n206 9.3005
R596 VTAIL.n205 VTAIL.n204 9.3005
R597 VTAIL.n198 VTAIL.n197 9.3005
R598 VTAIL.n223 VTAIL.n222 9.3005
R599 VTAIL.n186 VTAIL.n185 9.3005
R600 VTAIL.n229 VTAIL.n228 9.3005
R601 VTAIL.n231 VTAIL.n230 9.3005
R602 VTAIL.n182 VTAIL.n181 9.3005
R603 VTAIL.n237 VTAIL.n236 9.3005
R604 VTAIL.n239 VTAIL.n238 9.3005
R605 VTAIL.n240 VTAIL.n177 9.3005
R606 VTAIL.n247 VTAIL.n246 9.3005
R607 VTAIL.n532 VTAIL.n531 9.3005
R608 VTAIL.n575 VTAIL.n574 9.3005
R609 VTAIL.n577 VTAIL.n576 9.3005
R610 VTAIL.n528 VTAIL.n527 9.3005
R611 VTAIL.n583 VTAIL.n582 9.3005
R612 VTAIL.n585 VTAIL.n584 9.3005
R613 VTAIL.n523 VTAIL.n521 9.3005
R614 VTAIL.n591 VTAIL.n590 9.3005
R615 VTAIL.n599 VTAIL.n598 9.3005
R616 VTAIL.n518 VTAIL.n517 9.3005
R617 VTAIL.n593 VTAIL.n592 9.3005
R618 VTAIL.n569 VTAIL.n568 9.3005
R619 VTAIL.n567 VTAIL.n566 9.3005
R620 VTAIL.n536 VTAIL.n535 9.3005
R621 VTAIL.n561 VTAIL.n560 9.3005
R622 VTAIL.n559 VTAIL.n558 9.3005
R623 VTAIL.n540 VTAIL.n539 9.3005
R624 VTAIL.n553 VTAIL.n552 9.3005
R625 VTAIL.n551 VTAIL.n550 9.3005
R626 VTAIL.n544 VTAIL.n543 9.3005
R627 VTAIL.n446 VTAIL.n445 9.3005
R628 VTAIL.n489 VTAIL.n488 9.3005
R629 VTAIL.n491 VTAIL.n490 9.3005
R630 VTAIL.n442 VTAIL.n441 9.3005
R631 VTAIL.n497 VTAIL.n496 9.3005
R632 VTAIL.n499 VTAIL.n498 9.3005
R633 VTAIL.n437 VTAIL.n435 9.3005
R634 VTAIL.n505 VTAIL.n504 9.3005
R635 VTAIL.n513 VTAIL.n512 9.3005
R636 VTAIL.n432 VTAIL.n431 9.3005
R637 VTAIL.n507 VTAIL.n506 9.3005
R638 VTAIL.n483 VTAIL.n482 9.3005
R639 VTAIL.n481 VTAIL.n480 9.3005
R640 VTAIL.n450 VTAIL.n449 9.3005
R641 VTAIL.n475 VTAIL.n474 9.3005
R642 VTAIL.n473 VTAIL.n472 9.3005
R643 VTAIL.n454 VTAIL.n453 9.3005
R644 VTAIL.n467 VTAIL.n466 9.3005
R645 VTAIL.n465 VTAIL.n464 9.3005
R646 VTAIL.n458 VTAIL.n457 9.3005
R647 VTAIL.n360 VTAIL.n359 9.3005
R648 VTAIL.n403 VTAIL.n402 9.3005
R649 VTAIL.n405 VTAIL.n404 9.3005
R650 VTAIL.n356 VTAIL.n355 9.3005
R651 VTAIL.n411 VTAIL.n410 9.3005
R652 VTAIL.n413 VTAIL.n412 9.3005
R653 VTAIL.n351 VTAIL.n349 9.3005
R654 VTAIL.n419 VTAIL.n418 9.3005
R655 VTAIL.n427 VTAIL.n426 9.3005
R656 VTAIL.n346 VTAIL.n345 9.3005
R657 VTAIL.n421 VTAIL.n420 9.3005
R658 VTAIL.n397 VTAIL.n396 9.3005
R659 VTAIL.n395 VTAIL.n394 9.3005
R660 VTAIL.n364 VTAIL.n363 9.3005
R661 VTAIL.n389 VTAIL.n388 9.3005
R662 VTAIL.n387 VTAIL.n386 9.3005
R663 VTAIL.n368 VTAIL.n367 9.3005
R664 VTAIL.n381 VTAIL.n380 9.3005
R665 VTAIL.n379 VTAIL.n378 9.3005
R666 VTAIL.n372 VTAIL.n371 9.3005
R667 VTAIL.n274 VTAIL.n273 9.3005
R668 VTAIL.n317 VTAIL.n316 9.3005
R669 VTAIL.n319 VTAIL.n318 9.3005
R670 VTAIL.n270 VTAIL.n269 9.3005
R671 VTAIL.n325 VTAIL.n324 9.3005
R672 VTAIL.n327 VTAIL.n326 9.3005
R673 VTAIL.n265 VTAIL.n263 9.3005
R674 VTAIL.n333 VTAIL.n332 9.3005
R675 VTAIL.n341 VTAIL.n340 9.3005
R676 VTAIL.n260 VTAIL.n259 9.3005
R677 VTAIL.n335 VTAIL.n334 9.3005
R678 VTAIL.n311 VTAIL.n310 9.3005
R679 VTAIL.n309 VTAIL.n308 9.3005
R680 VTAIL.n278 VTAIL.n277 9.3005
R681 VTAIL.n303 VTAIL.n302 9.3005
R682 VTAIL.n301 VTAIL.n300 9.3005
R683 VTAIL.n282 VTAIL.n281 9.3005
R684 VTAIL.n295 VTAIL.n294 9.3005
R685 VTAIL.n293 VTAIL.n292 9.3005
R686 VTAIL.n286 VTAIL.n285 9.3005
R687 VTAIL.n646 VTAIL.n645 8.92171
R688 VTAIL.n661 VTAIL.n614 8.92171
R689 VTAIL.n44 VTAIL.n43 8.92171
R690 VTAIL.n59 VTAIL.n12 8.92171
R691 VTAIL.n130 VTAIL.n129 8.92171
R692 VTAIL.n145 VTAIL.n98 8.92171
R693 VTAIL.n216 VTAIL.n215 8.92171
R694 VTAIL.n231 VTAIL.n184 8.92171
R695 VTAIL.n577 VTAIL.n530 8.92171
R696 VTAIL.n562 VTAIL.n561 8.92171
R697 VTAIL.n491 VTAIL.n444 8.92171
R698 VTAIL.n476 VTAIL.n475 8.92171
R699 VTAIL.n405 VTAIL.n358 8.92171
R700 VTAIL.n390 VTAIL.n389 8.92171
R701 VTAIL.n319 VTAIL.n272 8.92171
R702 VTAIL.n304 VTAIL.n303 8.92171
R703 VTAIL.n649 VTAIL.n620 8.14595
R704 VTAIL.n658 VTAIL.n657 8.14595
R705 VTAIL.n47 VTAIL.n18 8.14595
R706 VTAIL.n56 VTAIL.n55 8.14595
R707 VTAIL.n133 VTAIL.n104 8.14595
R708 VTAIL.n142 VTAIL.n141 8.14595
R709 VTAIL.n219 VTAIL.n190 8.14595
R710 VTAIL.n228 VTAIL.n227 8.14595
R711 VTAIL.n574 VTAIL.n573 8.14595
R712 VTAIL.n565 VTAIL.n536 8.14595
R713 VTAIL.n488 VTAIL.n487 8.14595
R714 VTAIL.n479 VTAIL.n450 8.14595
R715 VTAIL.n402 VTAIL.n401 8.14595
R716 VTAIL.n393 VTAIL.n364 8.14595
R717 VTAIL.n316 VTAIL.n315 8.14595
R718 VTAIL.n307 VTAIL.n278 8.14595
R719 VTAIL.n650 VTAIL.n618 7.3702
R720 VTAIL.n654 VTAIL.n616 7.3702
R721 VTAIL.n48 VTAIL.n16 7.3702
R722 VTAIL.n52 VTAIL.n14 7.3702
R723 VTAIL.n134 VTAIL.n102 7.3702
R724 VTAIL.n138 VTAIL.n100 7.3702
R725 VTAIL.n220 VTAIL.n188 7.3702
R726 VTAIL.n224 VTAIL.n186 7.3702
R727 VTAIL.n570 VTAIL.n532 7.3702
R728 VTAIL.n566 VTAIL.n534 7.3702
R729 VTAIL.n484 VTAIL.n446 7.3702
R730 VTAIL.n480 VTAIL.n448 7.3702
R731 VTAIL.n398 VTAIL.n360 7.3702
R732 VTAIL.n394 VTAIL.n362 7.3702
R733 VTAIL.n312 VTAIL.n274 7.3702
R734 VTAIL.n308 VTAIL.n276 7.3702
R735 VTAIL.n653 VTAIL.n618 6.59444
R736 VTAIL.n654 VTAIL.n653 6.59444
R737 VTAIL.n51 VTAIL.n16 6.59444
R738 VTAIL.n52 VTAIL.n51 6.59444
R739 VTAIL.n137 VTAIL.n102 6.59444
R740 VTAIL.n138 VTAIL.n137 6.59444
R741 VTAIL.n223 VTAIL.n188 6.59444
R742 VTAIL.n224 VTAIL.n223 6.59444
R743 VTAIL.n570 VTAIL.n569 6.59444
R744 VTAIL.n569 VTAIL.n534 6.59444
R745 VTAIL.n484 VTAIL.n483 6.59444
R746 VTAIL.n483 VTAIL.n448 6.59444
R747 VTAIL.n398 VTAIL.n397 6.59444
R748 VTAIL.n397 VTAIL.n362 6.59444
R749 VTAIL.n312 VTAIL.n311 6.59444
R750 VTAIL.n311 VTAIL.n276 6.59444
R751 VTAIL.n650 VTAIL.n649 5.81868
R752 VTAIL.n657 VTAIL.n616 5.81868
R753 VTAIL.n48 VTAIL.n47 5.81868
R754 VTAIL.n55 VTAIL.n14 5.81868
R755 VTAIL.n134 VTAIL.n133 5.81868
R756 VTAIL.n141 VTAIL.n100 5.81868
R757 VTAIL.n220 VTAIL.n219 5.81868
R758 VTAIL.n227 VTAIL.n186 5.81868
R759 VTAIL.n573 VTAIL.n532 5.81868
R760 VTAIL.n566 VTAIL.n565 5.81868
R761 VTAIL.n487 VTAIL.n446 5.81868
R762 VTAIL.n480 VTAIL.n479 5.81868
R763 VTAIL.n401 VTAIL.n360 5.81868
R764 VTAIL.n394 VTAIL.n393 5.81868
R765 VTAIL.n315 VTAIL.n274 5.81868
R766 VTAIL.n308 VTAIL.n307 5.81868
R767 VTAIL.n646 VTAIL.n620 5.04292
R768 VTAIL.n658 VTAIL.n614 5.04292
R769 VTAIL.n44 VTAIL.n18 5.04292
R770 VTAIL.n56 VTAIL.n12 5.04292
R771 VTAIL.n130 VTAIL.n104 5.04292
R772 VTAIL.n142 VTAIL.n98 5.04292
R773 VTAIL.n216 VTAIL.n190 5.04292
R774 VTAIL.n228 VTAIL.n184 5.04292
R775 VTAIL.n574 VTAIL.n530 5.04292
R776 VTAIL.n562 VTAIL.n536 5.04292
R777 VTAIL.n488 VTAIL.n444 5.04292
R778 VTAIL.n476 VTAIL.n450 5.04292
R779 VTAIL.n402 VTAIL.n358 5.04292
R780 VTAIL.n390 VTAIL.n364 5.04292
R781 VTAIL.n316 VTAIL.n272 5.04292
R782 VTAIL.n304 VTAIL.n278 5.04292
R783 VTAIL.n629 VTAIL.n627 4.38563
R784 VTAIL.n27 VTAIL.n25 4.38563
R785 VTAIL.n113 VTAIL.n111 4.38563
R786 VTAIL.n199 VTAIL.n197 4.38563
R787 VTAIL.n545 VTAIL.n543 4.38563
R788 VTAIL.n459 VTAIL.n457 4.38563
R789 VTAIL.n373 VTAIL.n371 4.38563
R790 VTAIL.n287 VTAIL.n285 4.38563
R791 VTAIL.n645 VTAIL.n622 4.26717
R792 VTAIL.n662 VTAIL.n661 4.26717
R793 VTAIL.n43 VTAIL.n20 4.26717
R794 VTAIL.n60 VTAIL.n59 4.26717
R795 VTAIL.n129 VTAIL.n106 4.26717
R796 VTAIL.n146 VTAIL.n145 4.26717
R797 VTAIL.n215 VTAIL.n192 4.26717
R798 VTAIL.n232 VTAIL.n231 4.26717
R799 VTAIL.n578 VTAIL.n577 4.26717
R800 VTAIL.n561 VTAIL.n538 4.26717
R801 VTAIL.n492 VTAIL.n491 4.26717
R802 VTAIL.n475 VTAIL.n452 4.26717
R803 VTAIL.n406 VTAIL.n405 4.26717
R804 VTAIL.n389 VTAIL.n366 4.26717
R805 VTAIL.n320 VTAIL.n319 4.26717
R806 VTAIL.n303 VTAIL.n280 4.26717
R807 VTAIL.n642 VTAIL.n641 3.49141
R808 VTAIL.n665 VTAIL.n612 3.49141
R809 VTAIL.n40 VTAIL.n39 3.49141
R810 VTAIL.n63 VTAIL.n10 3.49141
R811 VTAIL.n126 VTAIL.n125 3.49141
R812 VTAIL.n149 VTAIL.n96 3.49141
R813 VTAIL.n212 VTAIL.n211 3.49141
R814 VTAIL.n235 VTAIL.n182 3.49141
R815 VTAIL.n581 VTAIL.n528 3.49141
R816 VTAIL.n558 VTAIL.n557 3.49141
R817 VTAIL.n495 VTAIL.n442 3.49141
R818 VTAIL.n472 VTAIL.n471 3.49141
R819 VTAIL.n409 VTAIL.n356 3.49141
R820 VTAIL.n386 VTAIL.n385 3.49141
R821 VTAIL.n323 VTAIL.n270 3.49141
R822 VTAIL.n300 VTAIL.n299 3.49141
R823 VTAIL.n429 VTAIL.n343 3.47464
R824 VTAIL.n601 VTAIL.n515 3.47464
R825 VTAIL.n257 VTAIL.n171 3.47464
R826 VTAIL.n638 VTAIL.n624 2.71565
R827 VTAIL.n666 VTAIL.n610 2.71565
R828 VTAIL.n686 VTAIL.n602 2.71565
R829 VTAIL.n36 VTAIL.n22 2.71565
R830 VTAIL.n64 VTAIL.n8 2.71565
R831 VTAIL.n84 VTAIL.n0 2.71565
R832 VTAIL.n122 VTAIL.n108 2.71565
R833 VTAIL.n150 VTAIL.n94 2.71565
R834 VTAIL.n170 VTAIL.n86 2.71565
R835 VTAIL.n208 VTAIL.n194 2.71565
R836 VTAIL.n236 VTAIL.n180 2.71565
R837 VTAIL.n256 VTAIL.n172 2.71565
R838 VTAIL.n600 VTAIL.n516 2.71565
R839 VTAIL.n582 VTAIL.n526 2.71565
R840 VTAIL.n554 VTAIL.n540 2.71565
R841 VTAIL.n514 VTAIL.n430 2.71565
R842 VTAIL.n496 VTAIL.n440 2.71565
R843 VTAIL.n468 VTAIL.n454 2.71565
R844 VTAIL.n428 VTAIL.n344 2.71565
R845 VTAIL.n410 VTAIL.n354 2.71565
R846 VTAIL.n382 VTAIL.n368 2.71565
R847 VTAIL.n342 VTAIL.n258 2.71565
R848 VTAIL.n324 VTAIL.n268 2.71565
R849 VTAIL.n296 VTAIL.n282 2.71565
R850 VTAIL.n637 VTAIL.n626 1.93989
R851 VTAIL.n671 VTAIL.n669 1.93989
R852 VTAIL.n684 VTAIL.n683 1.93989
R853 VTAIL.n35 VTAIL.n24 1.93989
R854 VTAIL.n69 VTAIL.n67 1.93989
R855 VTAIL.n82 VTAIL.n81 1.93989
R856 VTAIL.n121 VTAIL.n110 1.93989
R857 VTAIL.n155 VTAIL.n153 1.93989
R858 VTAIL.n168 VTAIL.n167 1.93989
R859 VTAIL.n207 VTAIL.n196 1.93989
R860 VTAIL.n241 VTAIL.n239 1.93989
R861 VTAIL.n254 VTAIL.n253 1.93989
R862 VTAIL.n598 VTAIL.n597 1.93989
R863 VTAIL.n586 VTAIL.n585 1.93989
R864 VTAIL.n553 VTAIL.n542 1.93989
R865 VTAIL.n512 VTAIL.n511 1.93989
R866 VTAIL.n500 VTAIL.n499 1.93989
R867 VTAIL.n467 VTAIL.n456 1.93989
R868 VTAIL.n426 VTAIL.n425 1.93989
R869 VTAIL.n414 VTAIL.n413 1.93989
R870 VTAIL.n381 VTAIL.n370 1.93989
R871 VTAIL.n340 VTAIL.n339 1.93989
R872 VTAIL.n328 VTAIL.n327 1.93989
R873 VTAIL.n295 VTAIL.n284 1.93989
R874 VTAIL VTAIL.n85 1.79576
R875 VTAIL VTAIL.n687 1.67938
R876 VTAIL.n634 VTAIL.n633 1.16414
R877 VTAIL.n670 VTAIL.n608 1.16414
R878 VTAIL.n680 VTAIL.n604 1.16414
R879 VTAIL.n32 VTAIL.n31 1.16414
R880 VTAIL.n68 VTAIL.n6 1.16414
R881 VTAIL.n78 VTAIL.n2 1.16414
R882 VTAIL.n118 VTAIL.n117 1.16414
R883 VTAIL.n154 VTAIL.n92 1.16414
R884 VTAIL.n164 VTAIL.n88 1.16414
R885 VTAIL.n204 VTAIL.n203 1.16414
R886 VTAIL.n240 VTAIL.n178 1.16414
R887 VTAIL.n250 VTAIL.n174 1.16414
R888 VTAIL.n594 VTAIL.n518 1.16414
R889 VTAIL.n589 VTAIL.n523 1.16414
R890 VTAIL.n550 VTAIL.n549 1.16414
R891 VTAIL.n508 VTAIL.n432 1.16414
R892 VTAIL.n503 VTAIL.n437 1.16414
R893 VTAIL.n464 VTAIL.n463 1.16414
R894 VTAIL.n422 VTAIL.n346 1.16414
R895 VTAIL.n417 VTAIL.n351 1.16414
R896 VTAIL.n378 VTAIL.n377 1.16414
R897 VTAIL.n336 VTAIL.n260 1.16414
R898 VTAIL.n331 VTAIL.n265 1.16414
R899 VTAIL.n292 VTAIL.n291 1.16414
R900 VTAIL.n515 VTAIL.n429 0.470328
R901 VTAIL.n171 VTAIL.n85 0.470328
R902 VTAIL.n630 VTAIL.n628 0.388379
R903 VTAIL.n676 VTAIL.n675 0.388379
R904 VTAIL.n679 VTAIL.n606 0.388379
R905 VTAIL.n28 VTAIL.n26 0.388379
R906 VTAIL.n74 VTAIL.n73 0.388379
R907 VTAIL.n77 VTAIL.n4 0.388379
R908 VTAIL.n114 VTAIL.n112 0.388379
R909 VTAIL.n160 VTAIL.n159 0.388379
R910 VTAIL.n163 VTAIL.n90 0.388379
R911 VTAIL.n200 VTAIL.n198 0.388379
R912 VTAIL.n246 VTAIL.n245 0.388379
R913 VTAIL.n249 VTAIL.n176 0.388379
R914 VTAIL.n593 VTAIL.n520 0.388379
R915 VTAIL.n590 VTAIL.n522 0.388379
R916 VTAIL.n546 VTAIL.n544 0.388379
R917 VTAIL.n507 VTAIL.n434 0.388379
R918 VTAIL.n504 VTAIL.n436 0.388379
R919 VTAIL.n460 VTAIL.n458 0.388379
R920 VTAIL.n421 VTAIL.n348 0.388379
R921 VTAIL.n418 VTAIL.n350 0.388379
R922 VTAIL.n374 VTAIL.n372 0.388379
R923 VTAIL.n335 VTAIL.n262 0.388379
R924 VTAIL.n332 VTAIL.n264 0.388379
R925 VTAIL.n288 VTAIL.n286 0.388379
R926 VTAIL.n635 VTAIL.n627 0.155672
R927 VTAIL.n636 VTAIL.n635 0.155672
R928 VTAIL.n636 VTAIL.n623 0.155672
R929 VTAIL.n643 VTAIL.n623 0.155672
R930 VTAIL.n644 VTAIL.n643 0.155672
R931 VTAIL.n644 VTAIL.n619 0.155672
R932 VTAIL.n651 VTAIL.n619 0.155672
R933 VTAIL.n652 VTAIL.n651 0.155672
R934 VTAIL.n652 VTAIL.n615 0.155672
R935 VTAIL.n659 VTAIL.n615 0.155672
R936 VTAIL.n660 VTAIL.n659 0.155672
R937 VTAIL.n660 VTAIL.n611 0.155672
R938 VTAIL.n667 VTAIL.n611 0.155672
R939 VTAIL.n668 VTAIL.n667 0.155672
R940 VTAIL.n668 VTAIL.n607 0.155672
R941 VTAIL.n677 VTAIL.n607 0.155672
R942 VTAIL.n678 VTAIL.n677 0.155672
R943 VTAIL.n678 VTAIL.n603 0.155672
R944 VTAIL.n685 VTAIL.n603 0.155672
R945 VTAIL.n33 VTAIL.n25 0.155672
R946 VTAIL.n34 VTAIL.n33 0.155672
R947 VTAIL.n34 VTAIL.n21 0.155672
R948 VTAIL.n41 VTAIL.n21 0.155672
R949 VTAIL.n42 VTAIL.n41 0.155672
R950 VTAIL.n42 VTAIL.n17 0.155672
R951 VTAIL.n49 VTAIL.n17 0.155672
R952 VTAIL.n50 VTAIL.n49 0.155672
R953 VTAIL.n50 VTAIL.n13 0.155672
R954 VTAIL.n57 VTAIL.n13 0.155672
R955 VTAIL.n58 VTAIL.n57 0.155672
R956 VTAIL.n58 VTAIL.n9 0.155672
R957 VTAIL.n65 VTAIL.n9 0.155672
R958 VTAIL.n66 VTAIL.n65 0.155672
R959 VTAIL.n66 VTAIL.n5 0.155672
R960 VTAIL.n75 VTAIL.n5 0.155672
R961 VTAIL.n76 VTAIL.n75 0.155672
R962 VTAIL.n76 VTAIL.n1 0.155672
R963 VTAIL.n83 VTAIL.n1 0.155672
R964 VTAIL.n119 VTAIL.n111 0.155672
R965 VTAIL.n120 VTAIL.n119 0.155672
R966 VTAIL.n120 VTAIL.n107 0.155672
R967 VTAIL.n127 VTAIL.n107 0.155672
R968 VTAIL.n128 VTAIL.n127 0.155672
R969 VTAIL.n128 VTAIL.n103 0.155672
R970 VTAIL.n135 VTAIL.n103 0.155672
R971 VTAIL.n136 VTAIL.n135 0.155672
R972 VTAIL.n136 VTAIL.n99 0.155672
R973 VTAIL.n143 VTAIL.n99 0.155672
R974 VTAIL.n144 VTAIL.n143 0.155672
R975 VTAIL.n144 VTAIL.n95 0.155672
R976 VTAIL.n151 VTAIL.n95 0.155672
R977 VTAIL.n152 VTAIL.n151 0.155672
R978 VTAIL.n152 VTAIL.n91 0.155672
R979 VTAIL.n161 VTAIL.n91 0.155672
R980 VTAIL.n162 VTAIL.n161 0.155672
R981 VTAIL.n162 VTAIL.n87 0.155672
R982 VTAIL.n169 VTAIL.n87 0.155672
R983 VTAIL.n205 VTAIL.n197 0.155672
R984 VTAIL.n206 VTAIL.n205 0.155672
R985 VTAIL.n206 VTAIL.n193 0.155672
R986 VTAIL.n213 VTAIL.n193 0.155672
R987 VTAIL.n214 VTAIL.n213 0.155672
R988 VTAIL.n214 VTAIL.n189 0.155672
R989 VTAIL.n221 VTAIL.n189 0.155672
R990 VTAIL.n222 VTAIL.n221 0.155672
R991 VTAIL.n222 VTAIL.n185 0.155672
R992 VTAIL.n229 VTAIL.n185 0.155672
R993 VTAIL.n230 VTAIL.n229 0.155672
R994 VTAIL.n230 VTAIL.n181 0.155672
R995 VTAIL.n237 VTAIL.n181 0.155672
R996 VTAIL.n238 VTAIL.n237 0.155672
R997 VTAIL.n238 VTAIL.n177 0.155672
R998 VTAIL.n247 VTAIL.n177 0.155672
R999 VTAIL.n248 VTAIL.n247 0.155672
R1000 VTAIL.n248 VTAIL.n173 0.155672
R1001 VTAIL.n255 VTAIL.n173 0.155672
R1002 VTAIL.n599 VTAIL.n517 0.155672
R1003 VTAIL.n592 VTAIL.n517 0.155672
R1004 VTAIL.n592 VTAIL.n591 0.155672
R1005 VTAIL.n591 VTAIL.n521 0.155672
R1006 VTAIL.n584 VTAIL.n521 0.155672
R1007 VTAIL.n584 VTAIL.n583 0.155672
R1008 VTAIL.n583 VTAIL.n527 0.155672
R1009 VTAIL.n576 VTAIL.n527 0.155672
R1010 VTAIL.n576 VTAIL.n575 0.155672
R1011 VTAIL.n575 VTAIL.n531 0.155672
R1012 VTAIL.n568 VTAIL.n531 0.155672
R1013 VTAIL.n568 VTAIL.n567 0.155672
R1014 VTAIL.n567 VTAIL.n535 0.155672
R1015 VTAIL.n560 VTAIL.n535 0.155672
R1016 VTAIL.n560 VTAIL.n559 0.155672
R1017 VTAIL.n559 VTAIL.n539 0.155672
R1018 VTAIL.n552 VTAIL.n539 0.155672
R1019 VTAIL.n552 VTAIL.n551 0.155672
R1020 VTAIL.n551 VTAIL.n543 0.155672
R1021 VTAIL.n513 VTAIL.n431 0.155672
R1022 VTAIL.n506 VTAIL.n431 0.155672
R1023 VTAIL.n506 VTAIL.n505 0.155672
R1024 VTAIL.n505 VTAIL.n435 0.155672
R1025 VTAIL.n498 VTAIL.n435 0.155672
R1026 VTAIL.n498 VTAIL.n497 0.155672
R1027 VTAIL.n497 VTAIL.n441 0.155672
R1028 VTAIL.n490 VTAIL.n441 0.155672
R1029 VTAIL.n490 VTAIL.n489 0.155672
R1030 VTAIL.n489 VTAIL.n445 0.155672
R1031 VTAIL.n482 VTAIL.n445 0.155672
R1032 VTAIL.n482 VTAIL.n481 0.155672
R1033 VTAIL.n481 VTAIL.n449 0.155672
R1034 VTAIL.n474 VTAIL.n449 0.155672
R1035 VTAIL.n474 VTAIL.n473 0.155672
R1036 VTAIL.n473 VTAIL.n453 0.155672
R1037 VTAIL.n466 VTAIL.n453 0.155672
R1038 VTAIL.n466 VTAIL.n465 0.155672
R1039 VTAIL.n465 VTAIL.n457 0.155672
R1040 VTAIL.n427 VTAIL.n345 0.155672
R1041 VTAIL.n420 VTAIL.n345 0.155672
R1042 VTAIL.n420 VTAIL.n419 0.155672
R1043 VTAIL.n419 VTAIL.n349 0.155672
R1044 VTAIL.n412 VTAIL.n349 0.155672
R1045 VTAIL.n412 VTAIL.n411 0.155672
R1046 VTAIL.n411 VTAIL.n355 0.155672
R1047 VTAIL.n404 VTAIL.n355 0.155672
R1048 VTAIL.n404 VTAIL.n403 0.155672
R1049 VTAIL.n403 VTAIL.n359 0.155672
R1050 VTAIL.n396 VTAIL.n359 0.155672
R1051 VTAIL.n396 VTAIL.n395 0.155672
R1052 VTAIL.n395 VTAIL.n363 0.155672
R1053 VTAIL.n388 VTAIL.n363 0.155672
R1054 VTAIL.n388 VTAIL.n387 0.155672
R1055 VTAIL.n387 VTAIL.n367 0.155672
R1056 VTAIL.n380 VTAIL.n367 0.155672
R1057 VTAIL.n380 VTAIL.n379 0.155672
R1058 VTAIL.n379 VTAIL.n371 0.155672
R1059 VTAIL.n341 VTAIL.n259 0.155672
R1060 VTAIL.n334 VTAIL.n259 0.155672
R1061 VTAIL.n334 VTAIL.n333 0.155672
R1062 VTAIL.n333 VTAIL.n263 0.155672
R1063 VTAIL.n326 VTAIL.n263 0.155672
R1064 VTAIL.n326 VTAIL.n325 0.155672
R1065 VTAIL.n325 VTAIL.n269 0.155672
R1066 VTAIL.n318 VTAIL.n269 0.155672
R1067 VTAIL.n318 VTAIL.n317 0.155672
R1068 VTAIL.n317 VTAIL.n273 0.155672
R1069 VTAIL.n310 VTAIL.n273 0.155672
R1070 VTAIL.n310 VTAIL.n309 0.155672
R1071 VTAIL.n309 VTAIL.n277 0.155672
R1072 VTAIL.n302 VTAIL.n277 0.155672
R1073 VTAIL.n302 VTAIL.n301 0.155672
R1074 VTAIL.n301 VTAIL.n281 0.155672
R1075 VTAIL.n294 VTAIL.n281 0.155672
R1076 VTAIL.n294 VTAIL.n293 0.155672
R1077 VTAIL.n293 VTAIL.n285 0.155672
R1078 VDD1 VDD1.n1 108.341
R1079 VDD1 VDD1.n0 60.5127
R1080 VDD1.n0 VDD1.t2 1.29124
R1081 VDD1.n0 VDD1.t3 1.29124
R1082 VDD1.n1 VDD1.t1 1.29124
R1083 VDD1.n1 VDD1.t0 1.29124
R1084 B.n917 B.n916 585
R1085 B.n361 B.n137 585
R1086 B.n360 B.n359 585
R1087 B.n358 B.n357 585
R1088 B.n356 B.n355 585
R1089 B.n354 B.n353 585
R1090 B.n352 B.n351 585
R1091 B.n350 B.n349 585
R1092 B.n348 B.n347 585
R1093 B.n346 B.n345 585
R1094 B.n344 B.n343 585
R1095 B.n342 B.n341 585
R1096 B.n340 B.n339 585
R1097 B.n338 B.n337 585
R1098 B.n336 B.n335 585
R1099 B.n334 B.n333 585
R1100 B.n332 B.n331 585
R1101 B.n330 B.n329 585
R1102 B.n328 B.n327 585
R1103 B.n326 B.n325 585
R1104 B.n324 B.n323 585
R1105 B.n322 B.n321 585
R1106 B.n320 B.n319 585
R1107 B.n318 B.n317 585
R1108 B.n316 B.n315 585
R1109 B.n314 B.n313 585
R1110 B.n312 B.n311 585
R1111 B.n310 B.n309 585
R1112 B.n308 B.n307 585
R1113 B.n306 B.n305 585
R1114 B.n304 B.n303 585
R1115 B.n302 B.n301 585
R1116 B.n300 B.n299 585
R1117 B.n298 B.n297 585
R1118 B.n296 B.n295 585
R1119 B.n294 B.n293 585
R1120 B.n292 B.n291 585
R1121 B.n290 B.n289 585
R1122 B.n288 B.n287 585
R1123 B.n286 B.n285 585
R1124 B.n284 B.n283 585
R1125 B.n282 B.n281 585
R1126 B.n280 B.n279 585
R1127 B.n278 B.n277 585
R1128 B.n276 B.n275 585
R1129 B.n274 B.n273 585
R1130 B.n272 B.n271 585
R1131 B.n270 B.n269 585
R1132 B.n268 B.n267 585
R1133 B.n266 B.n265 585
R1134 B.n264 B.n263 585
R1135 B.n261 B.n260 585
R1136 B.n259 B.n258 585
R1137 B.n257 B.n256 585
R1138 B.n255 B.n254 585
R1139 B.n253 B.n252 585
R1140 B.n251 B.n250 585
R1141 B.n249 B.n248 585
R1142 B.n247 B.n246 585
R1143 B.n245 B.n244 585
R1144 B.n243 B.n242 585
R1145 B.n240 B.n239 585
R1146 B.n238 B.n237 585
R1147 B.n236 B.n235 585
R1148 B.n234 B.n233 585
R1149 B.n232 B.n231 585
R1150 B.n230 B.n229 585
R1151 B.n228 B.n227 585
R1152 B.n226 B.n225 585
R1153 B.n224 B.n223 585
R1154 B.n222 B.n221 585
R1155 B.n220 B.n219 585
R1156 B.n218 B.n217 585
R1157 B.n216 B.n215 585
R1158 B.n214 B.n213 585
R1159 B.n212 B.n211 585
R1160 B.n210 B.n209 585
R1161 B.n208 B.n207 585
R1162 B.n206 B.n205 585
R1163 B.n204 B.n203 585
R1164 B.n202 B.n201 585
R1165 B.n200 B.n199 585
R1166 B.n198 B.n197 585
R1167 B.n196 B.n195 585
R1168 B.n194 B.n193 585
R1169 B.n192 B.n191 585
R1170 B.n190 B.n189 585
R1171 B.n188 B.n187 585
R1172 B.n186 B.n185 585
R1173 B.n184 B.n183 585
R1174 B.n182 B.n181 585
R1175 B.n180 B.n179 585
R1176 B.n178 B.n177 585
R1177 B.n176 B.n175 585
R1178 B.n174 B.n173 585
R1179 B.n172 B.n171 585
R1180 B.n170 B.n169 585
R1181 B.n168 B.n167 585
R1182 B.n166 B.n165 585
R1183 B.n164 B.n163 585
R1184 B.n162 B.n161 585
R1185 B.n160 B.n159 585
R1186 B.n158 B.n157 585
R1187 B.n156 B.n155 585
R1188 B.n154 B.n153 585
R1189 B.n152 B.n151 585
R1190 B.n150 B.n149 585
R1191 B.n148 B.n147 585
R1192 B.n146 B.n145 585
R1193 B.n144 B.n143 585
R1194 B.n82 B.n81 585
R1195 B.n922 B.n921 585
R1196 B.n915 B.n138 585
R1197 B.n138 B.n79 585
R1198 B.n914 B.n78 585
R1199 B.n926 B.n78 585
R1200 B.n913 B.n77 585
R1201 B.n927 B.n77 585
R1202 B.n912 B.n76 585
R1203 B.n928 B.n76 585
R1204 B.n911 B.n910 585
R1205 B.n910 B.n72 585
R1206 B.n909 B.n71 585
R1207 B.n934 B.n71 585
R1208 B.n908 B.n70 585
R1209 B.n935 B.n70 585
R1210 B.n907 B.n69 585
R1211 B.n936 B.n69 585
R1212 B.n906 B.n905 585
R1213 B.n905 B.n65 585
R1214 B.n904 B.n64 585
R1215 B.n942 B.n64 585
R1216 B.n903 B.n63 585
R1217 B.n943 B.n63 585
R1218 B.n902 B.n62 585
R1219 B.n944 B.n62 585
R1220 B.n901 B.n900 585
R1221 B.n900 B.n58 585
R1222 B.n899 B.n57 585
R1223 B.n950 B.n57 585
R1224 B.n898 B.n56 585
R1225 B.n951 B.n56 585
R1226 B.n897 B.n55 585
R1227 B.n952 B.n55 585
R1228 B.n896 B.n895 585
R1229 B.n895 B.n51 585
R1230 B.n894 B.n50 585
R1231 B.n958 B.n50 585
R1232 B.n893 B.n49 585
R1233 B.n959 B.n49 585
R1234 B.n892 B.n48 585
R1235 B.n960 B.n48 585
R1236 B.n891 B.n890 585
R1237 B.n890 B.n44 585
R1238 B.n889 B.n43 585
R1239 B.n966 B.n43 585
R1240 B.n888 B.n42 585
R1241 B.n967 B.n42 585
R1242 B.n887 B.n41 585
R1243 B.n968 B.n41 585
R1244 B.n886 B.n885 585
R1245 B.n885 B.n40 585
R1246 B.n884 B.n36 585
R1247 B.n974 B.n36 585
R1248 B.n883 B.n35 585
R1249 B.n975 B.n35 585
R1250 B.n882 B.n34 585
R1251 B.n976 B.n34 585
R1252 B.n881 B.n880 585
R1253 B.n880 B.n30 585
R1254 B.n879 B.n29 585
R1255 B.n982 B.n29 585
R1256 B.n878 B.n28 585
R1257 B.n983 B.n28 585
R1258 B.n877 B.n27 585
R1259 B.n984 B.n27 585
R1260 B.n876 B.n875 585
R1261 B.n875 B.n23 585
R1262 B.n874 B.n22 585
R1263 B.n990 B.n22 585
R1264 B.n873 B.n21 585
R1265 B.n991 B.n21 585
R1266 B.n872 B.n20 585
R1267 B.n992 B.n20 585
R1268 B.n871 B.n870 585
R1269 B.n870 B.n16 585
R1270 B.n869 B.n15 585
R1271 B.n998 B.n15 585
R1272 B.n868 B.n14 585
R1273 B.n999 B.n14 585
R1274 B.n867 B.n13 585
R1275 B.n1000 B.n13 585
R1276 B.n866 B.n865 585
R1277 B.n865 B.n12 585
R1278 B.n864 B.n863 585
R1279 B.n864 B.n8 585
R1280 B.n862 B.n7 585
R1281 B.n1007 B.n7 585
R1282 B.n861 B.n6 585
R1283 B.n1008 B.n6 585
R1284 B.n860 B.n5 585
R1285 B.n1009 B.n5 585
R1286 B.n859 B.n858 585
R1287 B.n858 B.n4 585
R1288 B.n857 B.n362 585
R1289 B.n857 B.n856 585
R1290 B.n847 B.n363 585
R1291 B.n364 B.n363 585
R1292 B.n849 B.n848 585
R1293 B.n850 B.n849 585
R1294 B.n846 B.n369 585
R1295 B.n369 B.n368 585
R1296 B.n845 B.n844 585
R1297 B.n844 B.n843 585
R1298 B.n371 B.n370 585
R1299 B.n372 B.n371 585
R1300 B.n836 B.n835 585
R1301 B.n837 B.n836 585
R1302 B.n834 B.n377 585
R1303 B.n377 B.n376 585
R1304 B.n833 B.n832 585
R1305 B.n832 B.n831 585
R1306 B.n379 B.n378 585
R1307 B.n380 B.n379 585
R1308 B.n824 B.n823 585
R1309 B.n825 B.n824 585
R1310 B.n822 B.n385 585
R1311 B.n385 B.n384 585
R1312 B.n821 B.n820 585
R1313 B.n820 B.n819 585
R1314 B.n387 B.n386 585
R1315 B.n388 B.n387 585
R1316 B.n812 B.n811 585
R1317 B.n813 B.n812 585
R1318 B.n810 B.n393 585
R1319 B.n393 B.n392 585
R1320 B.n809 B.n808 585
R1321 B.n808 B.n807 585
R1322 B.n395 B.n394 585
R1323 B.n800 B.n395 585
R1324 B.n799 B.n798 585
R1325 B.n801 B.n799 585
R1326 B.n797 B.n400 585
R1327 B.n400 B.n399 585
R1328 B.n796 B.n795 585
R1329 B.n795 B.n794 585
R1330 B.n402 B.n401 585
R1331 B.n403 B.n402 585
R1332 B.n787 B.n786 585
R1333 B.n788 B.n787 585
R1334 B.n785 B.n408 585
R1335 B.n408 B.n407 585
R1336 B.n784 B.n783 585
R1337 B.n783 B.n782 585
R1338 B.n410 B.n409 585
R1339 B.n411 B.n410 585
R1340 B.n775 B.n774 585
R1341 B.n776 B.n775 585
R1342 B.n773 B.n416 585
R1343 B.n416 B.n415 585
R1344 B.n772 B.n771 585
R1345 B.n771 B.n770 585
R1346 B.n418 B.n417 585
R1347 B.n419 B.n418 585
R1348 B.n763 B.n762 585
R1349 B.n764 B.n763 585
R1350 B.n761 B.n424 585
R1351 B.n424 B.n423 585
R1352 B.n760 B.n759 585
R1353 B.n759 B.n758 585
R1354 B.n426 B.n425 585
R1355 B.n427 B.n426 585
R1356 B.n751 B.n750 585
R1357 B.n752 B.n751 585
R1358 B.n749 B.n432 585
R1359 B.n432 B.n431 585
R1360 B.n748 B.n747 585
R1361 B.n747 B.n746 585
R1362 B.n434 B.n433 585
R1363 B.n435 B.n434 585
R1364 B.n739 B.n738 585
R1365 B.n740 B.n739 585
R1366 B.n737 B.n440 585
R1367 B.n440 B.n439 585
R1368 B.n736 B.n735 585
R1369 B.n735 B.n734 585
R1370 B.n442 B.n441 585
R1371 B.n443 B.n442 585
R1372 B.n730 B.n729 585
R1373 B.n446 B.n445 585
R1374 B.n726 B.n725 585
R1375 B.n727 B.n726 585
R1376 B.n724 B.n502 585
R1377 B.n723 B.n722 585
R1378 B.n721 B.n720 585
R1379 B.n719 B.n718 585
R1380 B.n717 B.n716 585
R1381 B.n715 B.n714 585
R1382 B.n713 B.n712 585
R1383 B.n711 B.n710 585
R1384 B.n709 B.n708 585
R1385 B.n707 B.n706 585
R1386 B.n705 B.n704 585
R1387 B.n703 B.n702 585
R1388 B.n701 B.n700 585
R1389 B.n699 B.n698 585
R1390 B.n697 B.n696 585
R1391 B.n695 B.n694 585
R1392 B.n693 B.n692 585
R1393 B.n691 B.n690 585
R1394 B.n689 B.n688 585
R1395 B.n687 B.n686 585
R1396 B.n685 B.n684 585
R1397 B.n683 B.n682 585
R1398 B.n681 B.n680 585
R1399 B.n679 B.n678 585
R1400 B.n677 B.n676 585
R1401 B.n675 B.n674 585
R1402 B.n673 B.n672 585
R1403 B.n671 B.n670 585
R1404 B.n669 B.n668 585
R1405 B.n667 B.n666 585
R1406 B.n665 B.n664 585
R1407 B.n663 B.n662 585
R1408 B.n661 B.n660 585
R1409 B.n659 B.n658 585
R1410 B.n657 B.n656 585
R1411 B.n655 B.n654 585
R1412 B.n653 B.n652 585
R1413 B.n651 B.n650 585
R1414 B.n649 B.n648 585
R1415 B.n647 B.n646 585
R1416 B.n645 B.n644 585
R1417 B.n643 B.n642 585
R1418 B.n641 B.n640 585
R1419 B.n639 B.n638 585
R1420 B.n637 B.n636 585
R1421 B.n635 B.n634 585
R1422 B.n633 B.n632 585
R1423 B.n631 B.n630 585
R1424 B.n629 B.n628 585
R1425 B.n627 B.n626 585
R1426 B.n625 B.n624 585
R1427 B.n623 B.n622 585
R1428 B.n621 B.n620 585
R1429 B.n619 B.n618 585
R1430 B.n617 B.n616 585
R1431 B.n615 B.n614 585
R1432 B.n613 B.n612 585
R1433 B.n611 B.n610 585
R1434 B.n609 B.n608 585
R1435 B.n607 B.n606 585
R1436 B.n605 B.n604 585
R1437 B.n603 B.n602 585
R1438 B.n601 B.n600 585
R1439 B.n599 B.n598 585
R1440 B.n597 B.n596 585
R1441 B.n595 B.n594 585
R1442 B.n593 B.n592 585
R1443 B.n591 B.n590 585
R1444 B.n589 B.n588 585
R1445 B.n587 B.n586 585
R1446 B.n585 B.n584 585
R1447 B.n583 B.n582 585
R1448 B.n581 B.n580 585
R1449 B.n579 B.n578 585
R1450 B.n577 B.n576 585
R1451 B.n575 B.n574 585
R1452 B.n573 B.n572 585
R1453 B.n571 B.n570 585
R1454 B.n569 B.n568 585
R1455 B.n567 B.n566 585
R1456 B.n565 B.n564 585
R1457 B.n563 B.n562 585
R1458 B.n561 B.n560 585
R1459 B.n559 B.n558 585
R1460 B.n557 B.n556 585
R1461 B.n555 B.n554 585
R1462 B.n553 B.n552 585
R1463 B.n551 B.n550 585
R1464 B.n549 B.n548 585
R1465 B.n547 B.n546 585
R1466 B.n545 B.n544 585
R1467 B.n543 B.n542 585
R1468 B.n541 B.n540 585
R1469 B.n539 B.n538 585
R1470 B.n537 B.n536 585
R1471 B.n535 B.n534 585
R1472 B.n533 B.n532 585
R1473 B.n531 B.n530 585
R1474 B.n529 B.n528 585
R1475 B.n527 B.n526 585
R1476 B.n525 B.n524 585
R1477 B.n523 B.n522 585
R1478 B.n521 B.n520 585
R1479 B.n519 B.n518 585
R1480 B.n517 B.n516 585
R1481 B.n515 B.n514 585
R1482 B.n513 B.n512 585
R1483 B.n511 B.n510 585
R1484 B.n509 B.n501 585
R1485 B.n727 B.n501 585
R1486 B.n731 B.n444 585
R1487 B.n444 B.n443 585
R1488 B.n733 B.n732 585
R1489 B.n734 B.n733 585
R1490 B.n438 B.n437 585
R1491 B.n439 B.n438 585
R1492 B.n742 B.n741 585
R1493 B.n741 B.n740 585
R1494 B.n743 B.n436 585
R1495 B.n436 B.n435 585
R1496 B.n745 B.n744 585
R1497 B.n746 B.n745 585
R1498 B.n430 B.n429 585
R1499 B.n431 B.n430 585
R1500 B.n754 B.n753 585
R1501 B.n753 B.n752 585
R1502 B.n755 B.n428 585
R1503 B.n428 B.n427 585
R1504 B.n757 B.n756 585
R1505 B.n758 B.n757 585
R1506 B.n422 B.n421 585
R1507 B.n423 B.n422 585
R1508 B.n766 B.n765 585
R1509 B.n765 B.n764 585
R1510 B.n767 B.n420 585
R1511 B.n420 B.n419 585
R1512 B.n769 B.n768 585
R1513 B.n770 B.n769 585
R1514 B.n414 B.n413 585
R1515 B.n415 B.n414 585
R1516 B.n778 B.n777 585
R1517 B.n777 B.n776 585
R1518 B.n779 B.n412 585
R1519 B.n412 B.n411 585
R1520 B.n781 B.n780 585
R1521 B.n782 B.n781 585
R1522 B.n406 B.n405 585
R1523 B.n407 B.n406 585
R1524 B.n790 B.n789 585
R1525 B.n789 B.n788 585
R1526 B.n791 B.n404 585
R1527 B.n404 B.n403 585
R1528 B.n793 B.n792 585
R1529 B.n794 B.n793 585
R1530 B.n398 B.n397 585
R1531 B.n399 B.n398 585
R1532 B.n803 B.n802 585
R1533 B.n802 B.n801 585
R1534 B.n804 B.n396 585
R1535 B.n800 B.n396 585
R1536 B.n806 B.n805 585
R1537 B.n807 B.n806 585
R1538 B.n391 B.n390 585
R1539 B.n392 B.n391 585
R1540 B.n815 B.n814 585
R1541 B.n814 B.n813 585
R1542 B.n816 B.n389 585
R1543 B.n389 B.n388 585
R1544 B.n818 B.n817 585
R1545 B.n819 B.n818 585
R1546 B.n383 B.n382 585
R1547 B.n384 B.n383 585
R1548 B.n827 B.n826 585
R1549 B.n826 B.n825 585
R1550 B.n828 B.n381 585
R1551 B.n381 B.n380 585
R1552 B.n830 B.n829 585
R1553 B.n831 B.n830 585
R1554 B.n375 B.n374 585
R1555 B.n376 B.n375 585
R1556 B.n839 B.n838 585
R1557 B.n838 B.n837 585
R1558 B.n840 B.n373 585
R1559 B.n373 B.n372 585
R1560 B.n842 B.n841 585
R1561 B.n843 B.n842 585
R1562 B.n367 B.n366 585
R1563 B.n368 B.n367 585
R1564 B.n852 B.n851 585
R1565 B.n851 B.n850 585
R1566 B.n853 B.n365 585
R1567 B.n365 B.n364 585
R1568 B.n855 B.n854 585
R1569 B.n856 B.n855 585
R1570 B.n3 B.n0 585
R1571 B.n4 B.n3 585
R1572 B.n1006 B.n1 585
R1573 B.n1007 B.n1006 585
R1574 B.n1005 B.n1004 585
R1575 B.n1005 B.n8 585
R1576 B.n1003 B.n9 585
R1577 B.n12 B.n9 585
R1578 B.n1002 B.n1001 585
R1579 B.n1001 B.n1000 585
R1580 B.n11 B.n10 585
R1581 B.n999 B.n11 585
R1582 B.n997 B.n996 585
R1583 B.n998 B.n997 585
R1584 B.n995 B.n17 585
R1585 B.n17 B.n16 585
R1586 B.n994 B.n993 585
R1587 B.n993 B.n992 585
R1588 B.n19 B.n18 585
R1589 B.n991 B.n19 585
R1590 B.n989 B.n988 585
R1591 B.n990 B.n989 585
R1592 B.n987 B.n24 585
R1593 B.n24 B.n23 585
R1594 B.n986 B.n985 585
R1595 B.n985 B.n984 585
R1596 B.n26 B.n25 585
R1597 B.n983 B.n26 585
R1598 B.n981 B.n980 585
R1599 B.n982 B.n981 585
R1600 B.n979 B.n31 585
R1601 B.n31 B.n30 585
R1602 B.n978 B.n977 585
R1603 B.n977 B.n976 585
R1604 B.n33 B.n32 585
R1605 B.n975 B.n33 585
R1606 B.n973 B.n972 585
R1607 B.n974 B.n973 585
R1608 B.n971 B.n37 585
R1609 B.n40 B.n37 585
R1610 B.n970 B.n969 585
R1611 B.n969 B.n968 585
R1612 B.n39 B.n38 585
R1613 B.n967 B.n39 585
R1614 B.n965 B.n964 585
R1615 B.n966 B.n965 585
R1616 B.n963 B.n45 585
R1617 B.n45 B.n44 585
R1618 B.n962 B.n961 585
R1619 B.n961 B.n960 585
R1620 B.n47 B.n46 585
R1621 B.n959 B.n47 585
R1622 B.n957 B.n956 585
R1623 B.n958 B.n957 585
R1624 B.n955 B.n52 585
R1625 B.n52 B.n51 585
R1626 B.n954 B.n953 585
R1627 B.n953 B.n952 585
R1628 B.n54 B.n53 585
R1629 B.n951 B.n54 585
R1630 B.n949 B.n948 585
R1631 B.n950 B.n949 585
R1632 B.n947 B.n59 585
R1633 B.n59 B.n58 585
R1634 B.n946 B.n945 585
R1635 B.n945 B.n944 585
R1636 B.n61 B.n60 585
R1637 B.n943 B.n61 585
R1638 B.n941 B.n940 585
R1639 B.n942 B.n941 585
R1640 B.n939 B.n66 585
R1641 B.n66 B.n65 585
R1642 B.n938 B.n937 585
R1643 B.n937 B.n936 585
R1644 B.n68 B.n67 585
R1645 B.n935 B.n68 585
R1646 B.n933 B.n932 585
R1647 B.n934 B.n933 585
R1648 B.n931 B.n73 585
R1649 B.n73 B.n72 585
R1650 B.n930 B.n929 585
R1651 B.n929 B.n928 585
R1652 B.n75 B.n74 585
R1653 B.n927 B.n75 585
R1654 B.n925 B.n924 585
R1655 B.n926 B.n925 585
R1656 B.n923 B.n80 585
R1657 B.n80 B.n79 585
R1658 B.n1010 B.n1009 585
R1659 B.n1008 B.n2 585
R1660 B.n921 B.n80 564.573
R1661 B.n917 B.n138 564.573
R1662 B.n501 B.n442 564.573
R1663 B.n729 B.n444 564.573
R1664 B.n139 B.t10 417.565
R1665 B.n506 B.t14 417.565
R1666 B.n141 B.t16 417.565
R1667 B.n503 B.t7 417.565
R1668 B.n140 B.t11 339.406
R1669 B.n507 B.t13 339.406
R1670 B.n142 B.t17 339.406
R1671 B.n504 B.t6 339.406
R1672 B.n141 B.t15 309.182
R1673 B.n139 B.t8 309.182
R1674 B.n506 B.t12 309.182
R1675 B.n503 B.t4 309.182
R1676 B.n919 B.n918 256.663
R1677 B.n919 B.n136 256.663
R1678 B.n919 B.n135 256.663
R1679 B.n919 B.n134 256.663
R1680 B.n919 B.n133 256.663
R1681 B.n919 B.n132 256.663
R1682 B.n919 B.n131 256.663
R1683 B.n919 B.n130 256.663
R1684 B.n919 B.n129 256.663
R1685 B.n919 B.n128 256.663
R1686 B.n919 B.n127 256.663
R1687 B.n919 B.n126 256.663
R1688 B.n919 B.n125 256.663
R1689 B.n919 B.n124 256.663
R1690 B.n919 B.n123 256.663
R1691 B.n919 B.n122 256.663
R1692 B.n919 B.n121 256.663
R1693 B.n919 B.n120 256.663
R1694 B.n919 B.n119 256.663
R1695 B.n919 B.n118 256.663
R1696 B.n919 B.n117 256.663
R1697 B.n919 B.n116 256.663
R1698 B.n919 B.n115 256.663
R1699 B.n919 B.n114 256.663
R1700 B.n919 B.n113 256.663
R1701 B.n919 B.n112 256.663
R1702 B.n919 B.n111 256.663
R1703 B.n919 B.n110 256.663
R1704 B.n919 B.n109 256.663
R1705 B.n919 B.n108 256.663
R1706 B.n919 B.n107 256.663
R1707 B.n919 B.n106 256.663
R1708 B.n919 B.n105 256.663
R1709 B.n919 B.n104 256.663
R1710 B.n919 B.n103 256.663
R1711 B.n919 B.n102 256.663
R1712 B.n919 B.n101 256.663
R1713 B.n919 B.n100 256.663
R1714 B.n919 B.n99 256.663
R1715 B.n919 B.n98 256.663
R1716 B.n919 B.n97 256.663
R1717 B.n919 B.n96 256.663
R1718 B.n919 B.n95 256.663
R1719 B.n919 B.n94 256.663
R1720 B.n919 B.n93 256.663
R1721 B.n919 B.n92 256.663
R1722 B.n919 B.n91 256.663
R1723 B.n919 B.n90 256.663
R1724 B.n919 B.n89 256.663
R1725 B.n919 B.n88 256.663
R1726 B.n919 B.n87 256.663
R1727 B.n919 B.n86 256.663
R1728 B.n919 B.n85 256.663
R1729 B.n919 B.n84 256.663
R1730 B.n919 B.n83 256.663
R1731 B.n920 B.n919 256.663
R1732 B.n728 B.n727 256.663
R1733 B.n727 B.n447 256.663
R1734 B.n727 B.n448 256.663
R1735 B.n727 B.n449 256.663
R1736 B.n727 B.n450 256.663
R1737 B.n727 B.n451 256.663
R1738 B.n727 B.n452 256.663
R1739 B.n727 B.n453 256.663
R1740 B.n727 B.n454 256.663
R1741 B.n727 B.n455 256.663
R1742 B.n727 B.n456 256.663
R1743 B.n727 B.n457 256.663
R1744 B.n727 B.n458 256.663
R1745 B.n727 B.n459 256.663
R1746 B.n727 B.n460 256.663
R1747 B.n727 B.n461 256.663
R1748 B.n727 B.n462 256.663
R1749 B.n727 B.n463 256.663
R1750 B.n727 B.n464 256.663
R1751 B.n727 B.n465 256.663
R1752 B.n727 B.n466 256.663
R1753 B.n727 B.n467 256.663
R1754 B.n727 B.n468 256.663
R1755 B.n727 B.n469 256.663
R1756 B.n727 B.n470 256.663
R1757 B.n727 B.n471 256.663
R1758 B.n727 B.n472 256.663
R1759 B.n727 B.n473 256.663
R1760 B.n727 B.n474 256.663
R1761 B.n727 B.n475 256.663
R1762 B.n727 B.n476 256.663
R1763 B.n727 B.n477 256.663
R1764 B.n727 B.n478 256.663
R1765 B.n727 B.n479 256.663
R1766 B.n727 B.n480 256.663
R1767 B.n727 B.n481 256.663
R1768 B.n727 B.n482 256.663
R1769 B.n727 B.n483 256.663
R1770 B.n727 B.n484 256.663
R1771 B.n727 B.n485 256.663
R1772 B.n727 B.n486 256.663
R1773 B.n727 B.n487 256.663
R1774 B.n727 B.n488 256.663
R1775 B.n727 B.n489 256.663
R1776 B.n727 B.n490 256.663
R1777 B.n727 B.n491 256.663
R1778 B.n727 B.n492 256.663
R1779 B.n727 B.n493 256.663
R1780 B.n727 B.n494 256.663
R1781 B.n727 B.n495 256.663
R1782 B.n727 B.n496 256.663
R1783 B.n727 B.n497 256.663
R1784 B.n727 B.n498 256.663
R1785 B.n727 B.n499 256.663
R1786 B.n727 B.n500 256.663
R1787 B.n1012 B.n1011 256.663
R1788 B.n143 B.n82 163.367
R1789 B.n147 B.n146 163.367
R1790 B.n151 B.n150 163.367
R1791 B.n155 B.n154 163.367
R1792 B.n159 B.n158 163.367
R1793 B.n163 B.n162 163.367
R1794 B.n167 B.n166 163.367
R1795 B.n171 B.n170 163.367
R1796 B.n175 B.n174 163.367
R1797 B.n179 B.n178 163.367
R1798 B.n183 B.n182 163.367
R1799 B.n187 B.n186 163.367
R1800 B.n191 B.n190 163.367
R1801 B.n195 B.n194 163.367
R1802 B.n199 B.n198 163.367
R1803 B.n203 B.n202 163.367
R1804 B.n207 B.n206 163.367
R1805 B.n211 B.n210 163.367
R1806 B.n215 B.n214 163.367
R1807 B.n219 B.n218 163.367
R1808 B.n223 B.n222 163.367
R1809 B.n227 B.n226 163.367
R1810 B.n231 B.n230 163.367
R1811 B.n235 B.n234 163.367
R1812 B.n239 B.n238 163.367
R1813 B.n244 B.n243 163.367
R1814 B.n248 B.n247 163.367
R1815 B.n252 B.n251 163.367
R1816 B.n256 B.n255 163.367
R1817 B.n260 B.n259 163.367
R1818 B.n265 B.n264 163.367
R1819 B.n269 B.n268 163.367
R1820 B.n273 B.n272 163.367
R1821 B.n277 B.n276 163.367
R1822 B.n281 B.n280 163.367
R1823 B.n285 B.n284 163.367
R1824 B.n289 B.n288 163.367
R1825 B.n293 B.n292 163.367
R1826 B.n297 B.n296 163.367
R1827 B.n301 B.n300 163.367
R1828 B.n305 B.n304 163.367
R1829 B.n309 B.n308 163.367
R1830 B.n313 B.n312 163.367
R1831 B.n317 B.n316 163.367
R1832 B.n321 B.n320 163.367
R1833 B.n325 B.n324 163.367
R1834 B.n329 B.n328 163.367
R1835 B.n333 B.n332 163.367
R1836 B.n337 B.n336 163.367
R1837 B.n341 B.n340 163.367
R1838 B.n345 B.n344 163.367
R1839 B.n349 B.n348 163.367
R1840 B.n353 B.n352 163.367
R1841 B.n357 B.n356 163.367
R1842 B.n359 B.n137 163.367
R1843 B.n735 B.n442 163.367
R1844 B.n735 B.n440 163.367
R1845 B.n739 B.n440 163.367
R1846 B.n739 B.n434 163.367
R1847 B.n747 B.n434 163.367
R1848 B.n747 B.n432 163.367
R1849 B.n751 B.n432 163.367
R1850 B.n751 B.n426 163.367
R1851 B.n759 B.n426 163.367
R1852 B.n759 B.n424 163.367
R1853 B.n763 B.n424 163.367
R1854 B.n763 B.n418 163.367
R1855 B.n771 B.n418 163.367
R1856 B.n771 B.n416 163.367
R1857 B.n775 B.n416 163.367
R1858 B.n775 B.n410 163.367
R1859 B.n783 B.n410 163.367
R1860 B.n783 B.n408 163.367
R1861 B.n787 B.n408 163.367
R1862 B.n787 B.n402 163.367
R1863 B.n795 B.n402 163.367
R1864 B.n795 B.n400 163.367
R1865 B.n799 B.n400 163.367
R1866 B.n799 B.n395 163.367
R1867 B.n808 B.n395 163.367
R1868 B.n808 B.n393 163.367
R1869 B.n812 B.n393 163.367
R1870 B.n812 B.n387 163.367
R1871 B.n820 B.n387 163.367
R1872 B.n820 B.n385 163.367
R1873 B.n824 B.n385 163.367
R1874 B.n824 B.n379 163.367
R1875 B.n832 B.n379 163.367
R1876 B.n832 B.n377 163.367
R1877 B.n836 B.n377 163.367
R1878 B.n836 B.n371 163.367
R1879 B.n844 B.n371 163.367
R1880 B.n844 B.n369 163.367
R1881 B.n849 B.n369 163.367
R1882 B.n849 B.n363 163.367
R1883 B.n857 B.n363 163.367
R1884 B.n858 B.n857 163.367
R1885 B.n858 B.n5 163.367
R1886 B.n6 B.n5 163.367
R1887 B.n7 B.n6 163.367
R1888 B.n864 B.n7 163.367
R1889 B.n865 B.n864 163.367
R1890 B.n865 B.n13 163.367
R1891 B.n14 B.n13 163.367
R1892 B.n15 B.n14 163.367
R1893 B.n870 B.n15 163.367
R1894 B.n870 B.n20 163.367
R1895 B.n21 B.n20 163.367
R1896 B.n22 B.n21 163.367
R1897 B.n875 B.n22 163.367
R1898 B.n875 B.n27 163.367
R1899 B.n28 B.n27 163.367
R1900 B.n29 B.n28 163.367
R1901 B.n880 B.n29 163.367
R1902 B.n880 B.n34 163.367
R1903 B.n35 B.n34 163.367
R1904 B.n36 B.n35 163.367
R1905 B.n885 B.n36 163.367
R1906 B.n885 B.n41 163.367
R1907 B.n42 B.n41 163.367
R1908 B.n43 B.n42 163.367
R1909 B.n890 B.n43 163.367
R1910 B.n890 B.n48 163.367
R1911 B.n49 B.n48 163.367
R1912 B.n50 B.n49 163.367
R1913 B.n895 B.n50 163.367
R1914 B.n895 B.n55 163.367
R1915 B.n56 B.n55 163.367
R1916 B.n57 B.n56 163.367
R1917 B.n900 B.n57 163.367
R1918 B.n900 B.n62 163.367
R1919 B.n63 B.n62 163.367
R1920 B.n64 B.n63 163.367
R1921 B.n905 B.n64 163.367
R1922 B.n905 B.n69 163.367
R1923 B.n70 B.n69 163.367
R1924 B.n71 B.n70 163.367
R1925 B.n910 B.n71 163.367
R1926 B.n910 B.n76 163.367
R1927 B.n77 B.n76 163.367
R1928 B.n78 B.n77 163.367
R1929 B.n138 B.n78 163.367
R1930 B.n726 B.n446 163.367
R1931 B.n726 B.n502 163.367
R1932 B.n722 B.n721 163.367
R1933 B.n718 B.n717 163.367
R1934 B.n714 B.n713 163.367
R1935 B.n710 B.n709 163.367
R1936 B.n706 B.n705 163.367
R1937 B.n702 B.n701 163.367
R1938 B.n698 B.n697 163.367
R1939 B.n694 B.n693 163.367
R1940 B.n690 B.n689 163.367
R1941 B.n686 B.n685 163.367
R1942 B.n682 B.n681 163.367
R1943 B.n678 B.n677 163.367
R1944 B.n674 B.n673 163.367
R1945 B.n670 B.n669 163.367
R1946 B.n666 B.n665 163.367
R1947 B.n662 B.n661 163.367
R1948 B.n658 B.n657 163.367
R1949 B.n654 B.n653 163.367
R1950 B.n650 B.n649 163.367
R1951 B.n646 B.n645 163.367
R1952 B.n642 B.n641 163.367
R1953 B.n638 B.n637 163.367
R1954 B.n634 B.n633 163.367
R1955 B.n630 B.n629 163.367
R1956 B.n626 B.n625 163.367
R1957 B.n622 B.n621 163.367
R1958 B.n618 B.n617 163.367
R1959 B.n614 B.n613 163.367
R1960 B.n610 B.n609 163.367
R1961 B.n606 B.n605 163.367
R1962 B.n602 B.n601 163.367
R1963 B.n598 B.n597 163.367
R1964 B.n594 B.n593 163.367
R1965 B.n590 B.n589 163.367
R1966 B.n586 B.n585 163.367
R1967 B.n582 B.n581 163.367
R1968 B.n578 B.n577 163.367
R1969 B.n574 B.n573 163.367
R1970 B.n570 B.n569 163.367
R1971 B.n566 B.n565 163.367
R1972 B.n562 B.n561 163.367
R1973 B.n558 B.n557 163.367
R1974 B.n554 B.n553 163.367
R1975 B.n550 B.n549 163.367
R1976 B.n546 B.n545 163.367
R1977 B.n542 B.n541 163.367
R1978 B.n538 B.n537 163.367
R1979 B.n534 B.n533 163.367
R1980 B.n530 B.n529 163.367
R1981 B.n526 B.n525 163.367
R1982 B.n522 B.n521 163.367
R1983 B.n518 B.n517 163.367
R1984 B.n514 B.n513 163.367
R1985 B.n510 B.n501 163.367
R1986 B.n733 B.n444 163.367
R1987 B.n733 B.n438 163.367
R1988 B.n741 B.n438 163.367
R1989 B.n741 B.n436 163.367
R1990 B.n745 B.n436 163.367
R1991 B.n745 B.n430 163.367
R1992 B.n753 B.n430 163.367
R1993 B.n753 B.n428 163.367
R1994 B.n757 B.n428 163.367
R1995 B.n757 B.n422 163.367
R1996 B.n765 B.n422 163.367
R1997 B.n765 B.n420 163.367
R1998 B.n769 B.n420 163.367
R1999 B.n769 B.n414 163.367
R2000 B.n777 B.n414 163.367
R2001 B.n777 B.n412 163.367
R2002 B.n781 B.n412 163.367
R2003 B.n781 B.n406 163.367
R2004 B.n789 B.n406 163.367
R2005 B.n789 B.n404 163.367
R2006 B.n793 B.n404 163.367
R2007 B.n793 B.n398 163.367
R2008 B.n802 B.n398 163.367
R2009 B.n802 B.n396 163.367
R2010 B.n806 B.n396 163.367
R2011 B.n806 B.n391 163.367
R2012 B.n814 B.n391 163.367
R2013 B.n814 B.n389 163.367
R2014 B.n818 B.n389 163.367
R2015 B.n818 B.n383 163.367
R2016 B.n826 B.n383 163.367
R2017 B.n826 B.n381 163.367
R2018 B.n830 B.n381 163.367
R2019 B.n830 B.n375 163.367
R2020 B.n838 B.n375 163.367
R2021 B.n838 B.n373 163.367
R2022 B.n842 B.n373 163.367
R2023 B.n842 B.n367 163.367
R2024 B.n851 B.n367 163.367
R2025 B.n851 B.n365 163.367
R2026 B.n855 B.n365 163.367
R2027 B.n855 B.n3 163.367
R2028 B.n1010 B.n3 163.367
R2029 B.n1006 B.n2 163.367
R2030 B.n1006 B.n1005 163.367
R2031 B.n1005 B.n9 163.367
R2032 B.n1001 B.n9 163.367
R2033 B.n1001 B.n11 163.367
R2034 B.n997 B.n11 163.367
R2035 B.n997 B.n17 163.367
R2036 B.n993 B.n17 163.367
R2037 B.n993 B.n19 163.367
R2038 B.n989 B.n19 163.367
R2039 B.n989 B.n24 163.367
R2040 B.n985 B.n24 163.367
R2041 B.n985 B.n26 163.367
R2042 B.n981 B.n26 163.367
R2043 B.n981 B.n31 163.367
R2044 B.n977 B.n31 163.367
R2045 B.n977 B.n33 163.367
R2046 B.n973 B.n33 163.367
R2047 B.n973 B.n37 163.367
R2048 B.n969 B.n37 163.367
R2049 B.n969 B.n39 163.367
R2050 B.n965 B.n39 163.367
R2051 B.n965 B.n45 163.367
R2052 B.n961 B.n45 163.367
R2053 B.n961 B.n47 163.367
R2054 B.n957 B.n47 163.367
R2055 B.n957 B.n52 163.367
R2056 B.n953 B.n52 163.367
R2057 B.n953 B.n54 163.367
R2058 B.n949 B.n54 163.367
R2059 B.n949 B.n59 163.367
R2060 B.n945 B.n59 163.367
R2061 B.n945 B.n61 163.367
R2062 B.n941 B.n61 163.367
R2063 B.n941 B.n66 163.367
R2064 B.n937 B.n66 163.367
R2065 B.n937 B.n68 163.367
R2066 B.n933 B.n68 163.367
R2067 B.n933 B.n73 163.367
R2068 B.n929 B.n73 163.367
R2069 B.n929 B.n75 163.367
R2070 B.n925 B.n75 163.367
R2071 B.n925 B.n80 163.367
R2072 B.n142 B.n141 78.1581
R2073 B.n140 B.n139 78.1581
R2074 B.n507 B.n506 78.1581
R2075 B.n504 B.n503 78.1581
R2076 B.n727 B.n443 72.0354
R2077 B.n919 B.n79 72.0354
R2078 B.n921 B.n920 71.676
R2079 B.n143 B.n83 71.676
R2080 B.n147 B.n84 71.676
R2081 B.n151 B.n85 71.676
R2082 B.n155 B.n86 71.676
R2083 B.n159 B.n87 71.676
R2084 B.n163 B.n88 71.676
R2085 B.n167 B.n89 71.676
R2086 B.n171 B.n90 71.676
R2087 B.n175 B.n91 71.676
R2088 B.n179 B.n92 71.676
R2089 B.n183 B.n93 71.676
R2090 B.n187 B.n94 71.676
R2091 B.n191 B.n95 71.676
R2092 B.n195 B.n96 71.676
R2093 B.n199 B.n97 71.676
R2094 B.n203 B.n98 71.676
R2095 B.n207 B.n99 71.676
R2096 B.n211 B.n100 71.676
R2097 B.n215 B.n101 71.676
R2098 B.n219 B.n102 71.676
R2099 B.n223 B.n103 71.676
R2100 B.n227 B.n104 71.676
R2101 B.n231 B.n105 71.676
R2102 B.n235 B.n106 71.676
R2103 B.n239 B.n107 71.676
R2104 B.n244 B.n108 71.676
R2105 B.n248 B.n109 71.676
R2106 B.n252 B.n110 71.676
R2107 B.n256 B.n111 71.676
R2108 B.n260 B.n112 71.676
R2109 B.n265 B.n113 71.676
R2110 B.n269 B.n114 71.676
R2111 B.n273 B.n115 71.676
R2112 B.n277 B.n116 71.676
R2113 B.n281 B.n117 71.676
R2114 B.n285 B.n118 71.676
R2115 B.n289 B.n119 71.676
R2116 B.n293 B.n120 71.676
R2117 B.n297 B.n121 71.676
R2118 B.n301 B.n122 71.676
R2119 B.n305 B.n123 71.676
R2120 B.n309 B.n124 71.676
R2121 B.n313 B.n125 71.676
R2122 B.n317 B.n126 71.676
R2123 B.n321 B.n127 71.676
R2124 B.n325 B.n128 71.676
R2125 B.n329 B.n129 71.676
R2126 B.n333 B.n130 71.676
R2127 B.n337 B.n131 71.676
R2128 B.n341 B.n132 71.676
R2129 B.n345 B.n133 71.676
R2130 B.n349 B.n134 71.676
R2131 B.n353 B.n135 71.676
R2132 B.n357 B.n136 71.676
R2133 B.n918 B.n137 71.676
R2134 B.n918 B.n917 71.676
R2135 B.n359 B.n136 71.676
R2136 B.n356 B.n135 71.676
R2137 B.n352 B.n134 71.676
R2138 B.n348 B.n133 71.676
R2139 B.n344 B.n132 71.676
R2140 B.n340 B.n131 71.676
R2141 B.n336 B.n130 71.676
R2142 B.n332 B.n129 71.676
R2143 B.n328 B.n128 71.676
R2144 B.n324 B.n127 71.676
R2145 B.n320 B.n126 71.676
R2146 B.n316 B.n125 71.676
R2147 B.n312 B.n124 71.676
R2148 B.n308 B.n123 71.676
R2149 B.n304 B.n122 71.676
R2150 B.n300 B.n121 71.676
R2151 B.n296 B.n120 71.676
R2152 B.n292 B.n119 71.676
R2153 B.n288 B.n118 71.676
R2154 B.n284 B.n117 71.676
R2155 B.n280 B.n116 71.676
R2156 B.n276 B.n115 71.676
R2157 B.n272 B.n114 71.676
R2158 B.n268 B.n113 71.676
R2159 B.n264 B.n112 71.676
R2160 B.n259 B.n111 71.676
R2161 B.n255 B.n110 71.676
R2162 B.n251 B.n109 71.676
R2163 B.n247 B.n108 71.676
R2164 B.n243 B.n107 71.676
R2165 B.n238 B.n106 71.676
R2166 B.n234 B.n105 71.676
R2167 B.n230 B.n104 71.676
R2168 B.n226 B.n103 71.676
R2169 B.n222 B.n102 71.676
R2170 B.n218 B.n101 71.676
R2171 B.n214 B.n100 71.676
R2172 B.n210 B.n99 71.676
R2173 B.n206 B.n98 71.676
R2174 B.n202 B.n97 71.676
R2175 B.n198 B.n96 71.676
R2176 B.n194 B.n95 71.676
R2177 B.n190 B.n94 71.676
R2178 B.n186 B.n93 71.676
R2179 B.n182 B.n92 71.676
R2180 B.n178 B.n91 71.676
R2181 B.n174 B.n90 71.676
R2182 B.n170 B.n89 71.676
R2183 B.n166 B.n88 71.676
R2184 B.n162 B.n87 71.676
R2185 B.n158 B.n86 71.676
R2186 B.n154 B.n85 71.676
R2187 B.n150 B.n84 71.676
R2188 B.n146 B.n83 71.676
R2189 B.n920 B.n82 71.676
R2190 B.n729 B.n728 71.676
R2191 B.n502 B.n447 71.676
R2192 B.n721 B.n448 71.676
R2193 B.n717 B.n449 71.676
R2194 B.n713 B.n450 71.676
R2195 B.n709 B.n451 71.676
R2196 B.n705 B.n452 71.676
R2197 B.n701 B.n453 71.676
R2198 B.n697 B.n454 71.676
R2199 B.n693 B.n455 71.676
R2200 B.n689 B.n456 71.676
R2201 B.n685 B.n457 71.676
R2202 B.n681 B.n458 71.676
R2203 B.n677 B.n459 71.676
R2204 B.n673 B.n460 71.676
R2205 B.n669 B.n461 71.676
R2206 B.n665 B.n462 71.676
R2207 B.n661 B.n463 71.676
R2208 B.n657 B.n464 71.676
R2209 B.n653 B.n465 71.676
R2210 B.n649 B.n466 71.676
R2211 B.n645 B.n467 71.676
R2212 B.n641 B.n468 71.676
R2213 B.n637 B.n469 71.676
R2214 B.n633 B.n470 71.676
R2215 B.n629 B.n471 71.676
R2216 B.n625 B.n472 71.676
R2217 B.n621 B.n473 71.676
R2218 B.n617 B.n474 71.676
R2219 B.n613 B.n475 71.676
R2220 B.n609 B.n476 71.676
R2221 B.n605 B.n477 71.676
R2222 B.n601 B.n478 71.676
R2223 B.n597 B.n479 71.676
R2224 B.n593 B.n480 71.676
R2225 B.n589 B.n481 71.676
R2226 B.n585 B.n482 71.676
R2227 B.n581 B.n483 71.676
R2228 B.n577 B.n484 71.676
R2229 B.n573 B.n485 71.676
R2230 B.n569 B.n486 71.676
R2231 B.n565 B.n487 71.676
R2232 B.n561 B.n488 71.676
R2233 B.n557 B.n489 71.676
R2234 B.n553 B.n490 71.676
R2235 B.n549 B.n491 71.676
R2236 B.n545 B.n492 71.676
R2237 B.n541 B.n493 71.676
R2238 B.n537 B.n494 71.676
R2239 B.n533 B.n495 71.676
R2240 B.n529 B.n496 71.676
R2241 B.n525 B.n497 71.676
R2242 B.n521 B.n498 71.676
R2243 B.n517 B.n499 71.676
R2244 B.n513 B.n500 71.676
R2245 B.n728 B.n446 71.676
R2246 B.n722 B.n447 71.676
R2247 B.n718 B.n448 71.676
R2248 B.n714 B.n449 71.676
R2249 B.n710 B.n450 71.676
R2250 B.n706 B.n451 71.676
R2251 B.n702 B.n452 71.676
R2252 B.n698 B.n453 71.676
R2253 B.n694 B.n454 71.676
R2254 B.n690 B.n455 71.676
R2255 B.n686 B.n456 71.676
R2256 B.n682 B.n457 71.676
R2257 B.n678 B.n458 71.676
R2258 B.n674 B.n459 71.676
R2259 B.n670 B.n460 71.676
R2260 B.n666 B.n461 71.676
R2261 B.n662 B.n462 71.676
R2262 B.n658 B.n463 71.676
R2263 B.n654 B.n464 71.676
R2264 B.n650 B.n465 71.676
R2265 B.n646 B.n466 71.676
R2266 B.n642 B.n467 71.676
R2267 B.n638 B.n468 71.676
R2268 B.n634 B.n469 71.676
R2269 B.n630 B.n470 71.676
R2270 B.n626 B.n471 71.676
R2271 B.n622 B.n472 71.676
R2272 B.n618 B.n473 71.676
R2273 B.n614 B.n474 71.676
R2274 B.n610 B.n475 71.676
R2275 B.n606 B.n476 71.676
R2276 B.n602 B.n477 71.676
R2277 B.n598 B.n478 71.676
R2278 B.n594 B.n479 71.676
R2279 B.n590 B.n480 71.676
R2280 B.n586 B.n481 71.676
R2281 B.n582 B.n482 71.676
R2282 B.n578 B.n483 71.676
R2283 B.n574 B.n484 71.676
R2284 B.n570 B.n485 71.676
R2285 B.n566 B.n486 71.676
R2286 B.n562 B.n487 71.676
R2287 B.n558 B.n488 71.676
R2288 B.n554 B.n489 71.676
R2289 B.n550 B.n490 71.676
R2290 B.n546 B.n491 71.676
R2291 B.n542 B.n492 71.676
R2292 B.n538 B.n493 71.676
R2293 B.n534 B.n494 71.676
R2294 B.n530 B.n495 71.676
R2295 B.n526 B.n496 71.676
R2296 B.n522 B.n497 71.676
R2297 B.n518 B.n498 71.676
R2298 B.n514 B.n499 71.676
R2299 B.n510 B.n500 71.676
R2300 B.n1011 B.n1010 71.676
R2301 B.n1011 B.n2 71.676
R2302 B.n241 B.n142 59.5399
R2303 B.n262 B.n140 59.5399
R2304 B.n508 B.n507 59.5399
R2305 B.n505 B.n504 59.5399
R2306 B.n731 B.n730 36.6834
R2307 B.n509 B.n441 36.6834
R2308 B.n916 B.n915 36.6834
R2309 B.n923 B.n922 36.6834
R2310 B.n734 B.n443 36.2848
R2311 B.n734 B.n439 36.2848
R2312 B.n740 B.n439 36.2848
R2313 B.n740 B.n435 36.2848
R2314 B.n746 B.n435 36.2848
R2315 B.n746 B.n431 36.2848
R2316 B.n752 B.n431 36.2848
R2317 B.n752 B.n427 36.2848
R2318 B.n758 B.n427 36.2848
R2319 B.n764 B.n423 36.2848
R2320 B.n764 B.n419 36.2848
R2321 B.n770 B.n419 36.2848
R2322 B.n770 B.n415 36.2848
R2323 B.n776 B.n415 36.2848
R2324 B.n776 B.n411 36.2848
R2325 B.n782 B.n411 36.2848
R2326 B.n782 B.n407 36.2848
R2327 B.n788 B.n407 36.2848
R2328 B.n788 B.n403 36.2848
R2329 B.n794 B.n403 36.2848
R2330 B.n794 B.n399 36.2848
R2331 B.n801 B.n399 36.2848
R2332 B.n801 B.n800 36.2848
R2333 B.n807 B.n392 36.2848
R2334 B.n813 B.n392 36.2848
R2335 B.n813 B.n388 36.2848
R2336 B.n819 B.n388 36.2848
R2337 B.n819 B.n384 36.2848
R2338 B.n825 B.n384 36.2848
R2339 B.n825 B.n380 36.2848
R2340 B.n831 B.n380 36.2848
R2341 B.n831 B.n376 36.2848
R2342 B.n837 B.n376 36.2848
R2343 B.n843 B.n372 36.2848
R2344 B.n843 B.n368 36.2848
R2345 B.n850 B.n368 36.2848
R2346 B.n850 B.n364 36.2848
R2347 B.n856 B.n364 36.2848
R2348 B.n856 B.n4 36.2848
R2349 B.n1009 B.n4 36.2848
R2350 B.n1009 B.n1008 36.2848
R2351 B.n1008 B.n1007 36.2848
R2352 B.n1007 B.n8 36.2848
R2353 B.n12 B.n8 36.2848
R2354 B.n1000 B.n12 36.2848
R2355 B.n1000 B.n999 36.2848
R2356 B.n999 B.n998 36.2848
R2357 B.n998 B.n16 36.2848
R2358 B.n992 B.n991 36.2848
R2359 B.n991 B.n990 36.2848
R2360 B.n990 B.n23 36.2848
R2361 B.n984 B.n23 36.2848
R2362 B.n984 B.n983 36.2848
R2363 B.n983 B.n982 36.2848
R2364 B.n982 B.n30 36.2848
R2365 B.n976 B.n30 36.2848
R2366 B.n976 B.n975 36.2848
R2367 B.n975 B.n974 36.2848
R2368 B.n968 B.n40 36.2848
R2369 B.n968 B.n967 36.2848
R2370 B.n967 B.n966 36.2848
R2371 B.n966 B.n44 36.2848
R2372 B.n960 B.n44 36.2848
R2373 B.n960 B.n959 36.2848
R2374 B.n959 B.n958 36.2848
R2375 B.n958 B.n51 36.2848
R2376 B.n952 B.n51 36.2848
R2377 B.n952 B.n951 36.2848
R2378 B.n951 B.n950 36.2848
R2379 B.n950 B.n58 36.2848
R2380 B.n944 B.n58 36.2848
R2381 B.n944 B.n943 36.2848
R2382 B.n942 B.n65 36.2848
R2383 B.n936 B.n65 36.2848
R2384 B.n936 B.n935 36.2848
R2385 B.n935 B.n934 36.2848
R2386 B.n934 B.n72 36.2848
R2387 B.n928 B.n72 36.2848
R2388 B.n928 B.n927 36.2848
R2389 B.n927 B.n926 36.2848
R2390 B.n926 B.n79 36.2848
R2391 B.n837 B.t2 35.2176
R2392 B.n992 B.t3 35.2176
R2393 B.t5 B.n423 34.1504
R2394 B.n943 B.t9 34.1504
R2395 B.n807 B.t1 32.016
R2396 B.n974 B.t0 32.016
R2397 B B.n1012 18.0485
R2398 B.n732 B.n731 10.6151
R2399 B.n732 B.n437 10.6151
R2400 B.n742 B.n437 10.6151
R2401 B.n743 B.n742 10.6151
R2402 B.n744 B.n743 10.6151
R2403 B.n744 B.n429 10.6151
R2404 B.n754 B.n429 10.6151
R2405 B.n755 B.n754 10.6151
R2406 B.n756 B.n755 10.6151
R2407 B.n756 B.n421 10.6151
R2408 B.n766 B.n421 10.6151
R2409 B.n767 B.n766 10.6151
R2410 B.n768 B.n767 10.6151
R2411 B.n768 B.n413 10.6151
R2412 B.n778 B.n413 10.6151
R2413 B.n779 B.n778 10.6151
R2414 B.n780 B.n779 10.6151
R2415 B.n780 B.n405 10.6151
R2416 B.n790 B.n405 10.6151
R2417 B.n791 B.n790 10.6151
R2418 B.n792 B.n791 10.6151
R2419 B.n792 B.n397 10.6151
R2420 B.n803 B.n397 10.6151
R2421 B.n804 B.n803 10.6151
R2422 B.n805 B.n804 10.6151
R2423 B.n805 B.n390 10.6151
R2424 B.n815 B.n390 10.6151
R2425 B.n816 B.n815 10.6151
R2426 B.n817 B.n816 10.6151
R2427 B.n817 B.n382 10.6151
R2428 B.n827 B.n382 10.6151
R2429 B.n828 B.n827 10.6151
R2430 B.n829 B.n828 10.6151
R2431 B.n829 B.n374 10.6151
R2432 B.n839 B.n374 10.6151
R2433 B.n840 B.n839 10.6151
R2434 B.n841 B.n840 10.6151
R2435 B.n841 B.n366 10.6151
R2436 B.n852 B.n366 10.6151
R2437 B.n853 B.n852 10.6151
R2438 B.n854 B.n853 10.6151
R2439 B.n854 B.n0 10.6151
R2440 B.n730 B.n445 10.6151
R2441 B.n725 B.n445 10.6151
R2442 B.n725 B.n724 10.6151
R2443 B.n724 B.n723 10.6151
R2444 B.n723 B.n720 10.6151
R2445 B.n720 B.n719 10.6151
R2446 B.n719 B.n716 10.6151
R2447 B.n716 B.n715 10.6151
R2448 B.n715 B.n712 10.6151
R2449 B.n712 B.n711 10.6151
R2450 B.n711 B.n708 10.6151
R2451 B.n708 B.n707 10.6151
R2452 B.n707 B.n704 10.6151
R2453 B.n704 B.n703 10.6151
R2454 B.n703 B.n700 10.6151
R2455 B.n700 B.n699 10.6151
R2456 B.n699 B.n696 10.6151
R2457 B.n696 B.n695 10.6151
R2458 B.n695 B.n692 10.6151
R2459 B.n692 B.n691 10.6151
R2460 B.n691 B.n688 10.6151
R2461 B.n688 B.n687 10.6151
R2462 B.n687 B.n684 10.6151
R2463 B.n684 B.n683 10.6151
R2464 B.n683 B.n680 10.6151
R2465 B.n680 B.n679 10.6151
R2466 B.n679 B.n676 10.6151
R2467 B.n676 B.n675 10.6151
R2468 B.n675 B.n672 10.6151
R2469 B.n672 B.n671 10.6151
R2470 B.n671 B.n668 10.6151
R2471 B.n668 B.n667 10.6151
R2472 B.n667 B.n664 10.6151
R2473 B.n664 B.n663 10.6151
R2474 B.n663 B.n660 10.6151
R2475 B.n660 B.n659 10.6151
R2476 B.n659 B.n656 10.6151
R2477 B.n656 B.n655 10.6151
R2478 B.n655 B.n652 10.6151
R2479 B.n652 B.n651 10.6151
R2480 B.n651 B.n648 10.6151
R2481 B.n648 B.n647 10.6151
R2482 B.n647 B.n644 10.6151
R2483 B.n644 B.n643 10.6151
R2484 B.n643 B.n640 10.6151
R2485 B.n640 B.n639 10.6151
R2486 B.n639 B.n636 10.6151
R2487 B.n636 B.n635 10.6151
R2488 B.n635 B.n632 10.6151
R2489 B.n632 B.n631 10.6151
R2490 B.n628 B.n627 10.6151
R2491 B.n627 B.n624 10.6151
R2492 B.n624 B.n623 10.6151
R2493 B.n623 B.n620 10.6151
R2494 B.n620 B.n619 10.6151
R2495 B.n619 B.n616 10.6151
R2496 B.n616 B.n615 10.6151
R2497 B.n615 B.n612 10.6151
R2498 B.n612 B.n611 10.6151
R2499 B.n608 B.n607 10.6151
R2500 B.n607 B.n604 10.6151
R2501 B.n604 B.n603 10.6151
R2502 B.n603 B.n600 10.6151
R2503 B.n600 B.n599 10.6151
R2504 B.n599 B.n596 10.6151
R2505 B.n596 B.n595 10.6151
R2506 B.n595 B.n592 10.6151
R2507 B.n592 B.n591 10.6151
R2508 B.n591 B.n588 10.6151
R2509 B.n588 B.n587 10.6151
R2510 B.n587 B.n584 10.6151
R2511 B.n584 B.n583 10.6151
R2512 B.n583 B.n580 10.6151
R2513 B.n580 B.n579 10.6151
R2514 B.n579 B.n576 10.6151
R2515 B.n576 B.n575 10.6151
R2516 B.n575 B.n572 10.6151
R2517 B.n572 B.n571 10.6151
R2518 B.n571 B.n568 10.6151
R2519 B.n568 B.n567 10.6151
R2520 B.n567 B.n564 10.6151
R2521 B.n564 B.n563 10.6151
R2522 B.n563 B.n560 10.6151
R2523 B.n560 B.n559 10.6151
R2524 B.n559 B.n556 10.6151
R2525 B.n556 B.n555 10.6151
R2526 B.n555 B.n552 10.6151
R2527 B.n552 B.n551 10.6151
R2528 B.n551 B.n548 10.6151
R2529 B.n548 B.n547 10.6151
R2530 B.n547 B.n544 10.6151
R2531 B.n544 B.n543 10.6151
R2532 B.n543 B.n540 10.6151
R2533 B.n540 B.n539 10.6151
R2534 B.n539 B.n536 10.6151
R2535 B.n536 B.n535 10.6151
R2536 B.n535 B.n532 10.6151
R2537 B.n532 B.n531 10.6151
R2538 B.n531 B.n528 10.6151
R2539 B.n528 B.n527 10.6151
R2540 B.n527 B.n524 10.6151
R2541 B.n524 B.n523 10.6151
R2542 B.n523 B.n520 10.6151
R2543 B.n520 B.n519 10.6151
R2544 B.n519 B.n516 10.6151
R2545 B.n516 B.n515 10.6151
R2546 B.n515 B.n512 10.6151
R2547 B.n512 B.n511 10.6151
R2548 B.n511 B.n509 10.6151
R2549 B.n736 B.n441 10.6151
R2550 B.n737 B.n736 10.6151
R2551 B.n738 B.n737 10.6151
R2552 B.n738 B.n433 10.6151
R2553 B.n748 B.n433 10.6151
R2554 B.n749 B.n748 10.6151
R2555 B.n750 B.n749 10.6151
R2556 B.n750 B.n425 10.6151
R2557 B.n760 B.n425 10.6151
R2558 B.n761 B.n760 10.6151
R2559 B.n762 B.n761 10.6151
R2560 B.n762 B.n417 10.6151
R2561 B.n772 B.n417 10.6151
R2562 B.n773 B.n772 10.6151
R2563 B.n774 B.n773 10.6151
R2564 B.n774 B.n409 10.6151
R2565 B.n784 B.n409 10.6151
R2566 B.n785 B.n784 10.6151
R2567 B.n786 B.n785 10.6151
R2568 B.n786 B.n401 10.6151
R2569 B.n796 B.n401 10.6151
R2570 B.n797 B.n796 10.6151
R2571 B.n798 B.n797 10.6151
R2572 B.n798 B.n394 10.6151
R2573 B.n809 B.n394 10.6151
R2574 B.n810 B.n809 10.6151
R2575 B.n811 B.n810 10.6151
R2576 B.n811 B.n386 10.6151
R2577 B.n821 B.n386 10.6151
R2578 B.n822 B.n821 10.6151
R2579 B.n823 B.n822 10.6151
R2580 B.n823 B.n378 10.6151
R2581 B.n833 B.n378 10.6151
R2582 B.n834 B.n833 10.6151
R2583 B.n835 B.n834 10.6151
R2584 B.n835 B.n370 10.6151
R2585 B.n845 B.n370 10.6151
R2586 B.n846 B.n845 10.6151
R2587 B.n848 B.n846 10.6151
R2588 B.n848 B.n847 10.6151
R2589 B.n847 B.n362 10.6151
R2590 B.n859 B.n362 10.6151
R2591 B.n860 B.n859 10.6151
R2592 B.n861 B.n860 10.6151
R2593 B.n862 B.n861 10.6151
R2594 B.n863 B.n862 10.6151
R2595 B.n866 B.n863 10.6151
R2596 B.n867 B.n866 10.6151
R2597 B.n868 B.n867 10.6151
R2598 B.n869 B.n868 10.6151
R2599 B.n871 B.n869 10.6151
R2600 B.n872 B.n871 10.6151
R2601 B.n873 B.n872 10.6151
R2602 B.n874 B.n873 10.6151
R2603 B.n876 B.n874 10.6151
R2604 B.n877 B.n876 10.6151
R2605 B.n878 B.n877 10.6151
R2606 B.n879 B.n878 10.6151
R2607 B.n881 B.n879 10.6151
R2608 B.n882 B.n881 10.6151
R2609 B.n883 B.n882 10.6151
R2610 B.n884 B.n883 10.6151
R2611 B.n886 B.n884 10.6151
R2612 B.n887 B.n886 10.6151
R2613 B.n888 B.n887 10.6151
R2614 B.n889 B.n888 10.6151
R2615 B.n891 B.n889 10.6151
R2616 B.n892 B.n891 10.6151
R2617 B.n893 B.n892 10.6151
R2618 B.n894 B.n893 10.6151
R2619 B.n896 B.n894 10.6151
R2620 B.n897 B.n896 10.6151
R2621 B.n898 B.n897 10.6151
R2622 B.n899 B.n898 10.6151
R2623 B.n901 B.n899 10.6151
R2624 B.n902 B.n901 10.6151
R2625 B.n903 B.n902 10.6151
R2626 B.n904 B.n903 10.6151
R2627 B.n906 B.n904 10.6151
R2628 B.n907 B.n906 10.6151
R2629 B.n908 B.n907 10.6151
R2630 B.n909 B.n908 10.6151
R2631 B.n911 B.n909 10.6151
R2632 B.n912 B.n911 10.6151
R2633 B.n913 B.n912 10.6151
R2634 B.n914 B.n913 10.6151
R2635 B.n915 B.n914 10.6151
R2636 B.n1004 B.n1 10.6151
R2637 B.n1004 B.n1003 10.6151
R2638 B.n1003 B.n1002 10.6151
R2639 B.n1002 B.n10 10.6151
R2640 B.n996 B.n10 10.6151
R2641 B.n996 B.n995 10.6151
R2642 B.n995 B.n994 10.6151
R2643 B.n994 B.n18 10.6151
R2644 B.n988 B.n18 10.6151
R2645 B.n988 B.n987 10.6151
R2646 B.n987 B.n986 10.6151
R2647 B.n986 B.n25 10.6151
R2648 B.n980 B.n25 10.6151
R2649 B.n980 B.n979 10.6151
R2650 B.n979 B.n978 10.6151
R2651 B.n978 B.n32 10.6151
R2652 B.n972 B.n32 10.6151
R2653 B.n972 B.n971 10.6151
R2654 B.n971 B.n970 10.6151
R2655 B.n970 B.n38 10.6151
R2656 B.n964 B.n38 10.6151
R2657 B.n964 B.n963 10.6151
R2658 B.n963 B.n962 10.6151
R2659 B.n962 B.n46 10.6151
R2660 B.n956 B.n46 10.6151
R2661 B.n956 B.n955 10.6151
R2662 B.n955 B.n954 10.6151
R2663 B.n954 B.n53 10.6151
R2664 B.n948 B.n53 10.6151
R2665 B.n948 B.n947 10.6151
R2666 B.n947 B.n946 10.6151
R2667 B.n946 B.n60 10.6151
R2668 B.n940 B.n60 10.6151
R2669 B.n940 B.n939 10.6151
R2670 B.n939 B.n938 10.6151
R2671 B.n938 B.n67 10.6151
R2672 B.n932 B.n67 10.6151
R2673 B.n932 B.n931 10.6151
R2674 B.n931 B.n930 10.6151
R2675 B.n930 B.n74 10.6151
R2676 B.n924 B.n74 10.6151
R2677 B.n924 B.n923 10.6151
R2678 B.n922 B.n81 10.6151
R2679 B.n144 B.n81 10.6151
R2680 B.n145 B.n144 10.6151
R2681 B.n148 B.n145 10.6151
R2682 B.n149 B.n148 10.6151
R2683 B.n152 B.n149 10.6151
R2684 B.n153 B.n152 10.6151
R2685 B.n156 B.n153 10.6151
R2686 B.n157 B.n156 10.6151
R2687 B.n160 B.n157 10.6151
R2688 B.n161 B.n160 10.6151
R2689 B.n164 B.n161 10.6151
R2690 B.n165 B.n164 10.6151
R2691 B.n168 B.n165 10.6151
R2692 B.n169 B.n168 10.6151
R2693 B.n172 B.n169 10.6151
R2694 B.n173 B.n172 10.6151
R2695 B.n176 B.n173 10.6151
R2696 B.n177 B.n176 10.6151
R2697 B.n180 B.n177 10.6151
R2698 B.n181 B.n180 10.6151
R2699 B.n184 B.n181 10.6151
R2700 B.n185 B.n184 10.6151
R2701 B.n188 B.n185 10.6151
R2702 B.n189 B.n188 10.6151
R2703 B.n192 B.n189 10.6151
R2704 B.n193 B.n192 10.6151
R2705 B.n196 B.n193 10.6151
R2706 B.n197 B.n196 10.6151
R2707 B.n200 B.n197 10.6151
R2708 B.n201 B.n200 10.6151
R2709 B.n204 B.n201 10.6151
R2710 B.n205 B.n204 10.6151
R2711 B.n208 B.n205 10.6151
R2712 B.n209 B.n208 10.6151
R2713 B.n212 B.n209 10.6151
R2714 B.n213 B.n212 10.6151
R2715 B.n216 B.n213 10.6151
R2716 B.n217 B.n216 10.6151
R2717 B.n220 B.n217 10.6151
R2718 B.n221 B.n220 10.6151
R2719 B.n224 B.n221 10.6151
R2720 B.n225 B.n224 10.6151
R2721 B.n228 B.n225 10.6151
R2722 B.n229 B.n228 10.6151
R2723 B.n232 B.n229 10.6151
R2724 B.n233 B.n232 10.6151
R2725 B.n236 B.n233 10.6151
R2726 B.n237 B.n236 10.6151
R2727 B.n240 B.n237 10.6151
R2728 B.n245 B.n242 10.6151
R2729 B.n246 B.n245 10.6151
R2730 B.n249 B.n246 10.6151
R2731 B.n250 B.n249 10.6151
R2732 B.n253 B.n250 10.6151
R2733 B.n254 B.n253 10.6151
R2734 B.n257 B.n254 10.6151
R2735 B.n258 B.n257 10.6151
R2736 B.n261 B.n258 10.6151
R2737 B.n266 B.n263 10.6151
R2738 B.n267 B.n266 10.6151
R2739 B.n270 B.n267 10.6151
R2740 B.n271 B.n270 10.6151
R2741 B.n274 B.n271 10.6151
R2742 B.n275 B.n274 10.6151
R2743 B.n278 B.n275 10.6151
R2744 B.n279 B.n278 10.6151
R2745 B.n282 B.n279 10.6151
R2746 B.n283 B.n282 10.6151
R2747 B.n286 B.n283 10.6151
R2748 B.n287 B.n286 10.6151
R2749 B.n290 B.n287 10.6151
R2750 B.n291 B.n290 10.6151
R2751 B.n294 B.n291 10.6151
R2752 B.n295 B.n294 10.6151
R2753 B.n298 B.n295 10.6151
R2754 B.n299 B.n298 10.6151
R2755 B.n302 B.n299 10.6151
R2756 B.n303 B.n302 10.6151
R2757 B.n306 B.n303 10.6151
R2758 B.n307 B.n306 10.6151
R2759 B.n310 B.n307 10.6151
R2760 B.n311 B.n310 10.6151
R2761 B.n314 B.n311 10.6151
R2762 B.n315 B.n314 10.6151
R2763 B.n318 B.n315 10.6151
R2764 B.n319 B.n318 10.6151
R2765 B.n322 B.n319 10.6151
R2766 B.n323 B.n322 10.6151
R2767 B.n326 B.n323 10.6151
R2768 B.n327 B.n326 10.6151
R2769 B.n330 B.n327 10.6151
R2770 B.n331 B.n330 10.6151
R2771 B.n334 B.n331 10.6151
R2772 B.n335 B.n334 10.6151
R2773 B.n338 B.n335 10.6151
R2774 B.n339 B.n338 10.6151
R2775 B.n342 B.n339 10.6151
R2776 B.n343 B.n342 10.6151
R2777 B.n346 B.n343 10.6151
R2778 B.n347 B.n346 10.6151
R2779 B.n350 B.n347 10.6151
R2780 B.n351 B.n350 10.6151
R2781 B.n354 B.n351 10.6151
R2782 B.n355 B.n354 10.6151
R2783 B.n358 B.n355 10.6151
R2784 B.n360 B.n358 10.6151
R2785 B.n361 B.n360 10.6151
R2786 B.n916 B.n361 10.6151
R2787 B.n631 B.n505 9.36635
R2788 B.n608 B.n508 9.36635
R2789 B.n241 B.n240 9.36635
R2790 B.n263 B.n262 9.36635
R2791 B.n1012 B.n0 8.11757
R2792 B.n1012 B.n1 8.11757
R2793 B.n800 B.t1 4.26924
R2794 B.n40 B.t0 4.26924
R2795 B.n758 B.t5 2.13487
R2796 B.t9 B.n942 2.13487
R2797 B.n628 B.n505 1.24928
R2798 B.n611 B.n508 1.24928
R2799 B.n242 B.n241 1.24928
R2800 B.n262 B.n261 1.24928
R2801 B.t2 B.n372 1.06768
R2802 B.t3 B.n16 1.06768
R2803 VN.n1 VN.t2 133.266
R2804 VN.n0 VN.t3 133.266
R2805 VN.n0 VN.t0 131.939
R2806 VN.n1 VN.t1 131.939
R2807 VN VN.n1 54.2889
R2808 VN VN.n0 1.92908
R2809 VDD2.n2 VDD2.n0 107.816
R2810 VDD2.n2 VDD2.n1 60.4545
R2811 VDD2.n1 VDD2.t2 1.29124
R2812 VDD2.n1 VDD2.t1 1.29124
R2813 VDD2.n0 VDD2.t0 1.29124
R2814 VDD2.n0 VDD2.t3 1.29124
R2815 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 6.47393f
C1 VN VP 7.60106f
C2 VDD1 VDD2 1.2916f
C3 VTAIL VP 6.248971f
C4 VDD1 VP 6.63779f
C5 VN VTAIL 6.23487f
C6 VDD2 VP 0.464488f
C7 VDD1 VN 0.150182f
C8 VDD1 VTAIL 6.41235f
C9 VDD2 VN 6.3245f
C10 VDD2 B 4.646266f
C11 VDD1 B 9.494009f
C12 VTAIL B 12.708332f
C13 VN B 13.08293f
C14 VP B 11.505142f
C15 VDD2.t0 B 0.326579f
C16 VDD2.t3 B 0.326579f
C17 VDD2.n0 B 3.82494f
C18 VDD2.t2 B 0.326579f
C19 VDD2.t1 B 0.326579f
C20 VDD2.n1 B 2.95439f
C21 VDD2.n2 B 4.40697f
C22 VN.t0 B 3.30861f
C23 VN.t3 B 3.32013f
C24 VN.n0 B 2.02256f
C25 VN.t1 B 3.30861f
C26 VN.t2 B 3.32013f
C27 VN.n1 B 3.36513f
C28 VDD1.t2 B 0.329123f
C29 VDD1.t3 B 0.329123f
C30 VDD1.n0 B 2.97793f
C31 VDD1.t1 B 0.329123f
C32 VDD1.t0 B 0.329123f
C33 VDD1.n1 B 3.88366f
C34 VTAIL.n0 B 0.020801f
C35 VTAIL.n1 B 0.016198f
C36 VTAIL.n2 B 0.008704f
C37 VTAIL.n3 B 0.020574f
C38 VTAIL.n4 B 0.00896f
C39 VTAIL.n5 B 0.016198f
C40 VTAIL.n6 B 0.009216f
C41 VTAIL.n7 B 0.020574f
C42 VTAIL.n8 B 0.009216f
C43 VTAIL.n9 B 0.016198f
C44 VTAIL.n10 B 0.008704f
C45 VTAIL.n11 B 0.020574f
C46 VTAIL.n12 B 0.009216f
C47 VTAIL.n13 B 0.016198f
C48 VTAIL.n14 B 0.008704f
C49 VTAIL.n15 B 0.020574f
C50 VTAIL.n16 B 0.009216f
C51 VTAIL.n17 B 0.016198f
C52 VTAIL.n18 B 0.008704f
C53 VTAIL.n19 B 0.020574f
C54 VTAIL.n20 B 0.009216f
C55 VTAIL.n21 B 0.016198f
C56 VTAIL.n22 B 0.008704f
C57 VTAIL.n23 B 0.020574f
C58 VTAIL.n24 B 0.009216f
C59 VTAIL.n25 B 1.07913f
C60 VTAIL.n26 B 0.008704f
C61 VTAIL.t3 B 0.033943f
C62 VTAIL.n27 B 0.10703f
C63 VTAIL.n28 B 0.012154f
C64 VTAIL.n29 B 0.01543f
C65 VTAIL.n30 B 0.020574f
C66 VTAIL.n31 B 0.009216f
C67 VTAIL.n32 B 0.008704f
C68 VTAIL.n33 B 0.016198f
C69 VTAIL.n34 B 0.016198f
C70 VTAIL.n35 B 0.008704f
C71 VTAIL.n36 B 0.009216f
C72 VTAIL.n37 B 0.020574f
C73 VTAIL.n38 B 0.020574f
C74 VTAIL.n39 B 0.009216f
C75 VTAIL.n40 B 0.008704f
C76 VTAIL.n41 B 0.016198f
C77 VTAIL.n42 B 0.016198f
C78 VTAIL.n43 B 0.008704f
C79 VTAIL.n44 B 0.009216f
C80 VTAIL.n45 B 0.020574f
C81 VTAIL.n46 B 0.020574f
C82 VTAIL.n47 B 0.009216f
C83 VTAIL.n48 B 0.008704f
C84 VTAIL.n49 B 0.016198f
C85 VTAIL.n50 B 0.016198f
C86 VTAIL.n51 B 0.008704f
C87 VTAIL.n52 B 0.009216f
C88 VTAIL.n53 B 0.020574f
C89 VTAIL.n54 B 0.020574f
C90 VTAIL.n55 B 0.009216f
C91 VTAIL.n56 B 0.008704f
C92 VTAIL.n57 B 0.016198f
C93 VTAIL.n58 B 0.016198f
C94 VTAIL.n59 B 0.008704f
C95 VTAIL.n60 B 0.009216f
C96 VTAIL.n61 B 0.020574f
C97 VTAIL.n62 B 0.020574f
C98 VTAIL.n63 B 0.009216f
C99 VTAIL.n64 B 0.008704f
C100 VTAIL.n65 B 0.016198f
C101 VTAIL.n66 B 0.016198f
C102 VTAIL.n67 B 0.008704f
C103 VTAIL.n68 B 0.008704f
C104 VTAIL.n69 B 0.009216f
C105 VTAIL.n70 B 0.020574f
C106 VTAIL.n71 B 0.020574f
C107 VTAIL.n72 B 0.020574f
C108 VTAIL.n73 B 0.00896f
C109 VTAIL.n74 B 0.008704f
C110 VTAIL.n75 B 0.016198f
C111 VTAIL.n76 B 0.016198f
C112 VTAIL.n77 B 0.008704f
C113 VTAIL.n78 B 0.009216f
C114 VTAIL.n79 B 0.020574f
C115 VTAIL.n80 B 0.04106f
C116 VTAIL.n81 B 0.009216f
C117 VTAIL.n82 B 0.008704f
C118 VTAIL.n83 B 0.036999f
C119 VTAIL.n84 B 0.022604f
C120 VTAIL.n85 B 0.13181f
C121 VTAIL.n86 B 0.020801f
C122 VTAIL.n87 B 0.016198f
C123 VTAIL.n88 B 0.008704f
C124 VTAIL.n89 B 0.020574f
C125 VTAIL.n90 B 0.00896f
C126 VTAIL.n91 B 0.016198f
C127 VTAIL.n92 B 0.009216f
C128 VTAIL.n93 B 0.020574f
C129 VTAIL.n94 B 0.009216f
C130 VTAIL.n95 B 0.016198f
C131 VTAIL.n96 B 0.008704f
C132 VTAIL.n97 B 0.020574f
C133 VTAIL.n98 B 0.009216f
C134 VTAIL.n99 B 0.016198f
C135 VTAIL.n100 B 0.008704f
C136 VTAIL.n101 B 0.020574f
C137 VTAIL.n102 B 0.009216f
C138 VTAIL.n103 B 0.016198f
C139 VTAIL.n104 B 0.008704f
C140 VTAIL.n105 B 0.020574f
C141 VTAIL.n106 B 0.009216f
C142 VTAIL.n107 B 0.016198f
C143 VTAIL.n108 B 0.008704f
C144 VTAIL.n109 B 0.020574f
C145 VTAIL.n110 B 0.009216f
C146 VTAIL.n111 B 1.07913f
C147 VTAIL.n112 B 0.008704f
C148 VTAIL.t5 B 0.033943f
C149 VTAIL.n113 B 0.10703f
C150 VTAIL.n114 B 0.012154f
C151 VTAIL.n115 B 0.01543f
C152 VTAIL.n116 B 0.020574f
C153 VTAIL.n117 B 0.009216f
C154 VTAIL.n118 B 0.008704f
C155 VTAIL.n119 B 0.016198f
C156 VTAIL.n120 B 0.016198f
C157 VTAIL.n121 B 0.008704f
C158 VTAIL.n122 B 0.009216f
C159 VTAIL.n123 B 0.020574f
C160 VTAIL.n124 B 0.020574f
C161 VTAIL.n125 B 0.009216f
C162 VTAIL.n126 B 0.008704f
C163 VTAIL.n127 B 0.016198f
C164 VTAIL.n128 B 0.016198f
C165 VTAIL.n129 B 0.008704f
C166 VTAIL.n130 B 0.009216f
C167 VTAIL.n131 B 0.020574f
C168 VTAIL.n132 B 0.020574f
C169 VTAIL.n133 B 0.009216f
C170 VTAIL.n134 B 0.008704f
C171 VTAIL.n135 B 0.016198f
C172 VTAIL.n136 B 0.016198f
C173 VTAIL.n137 B 0.008704f
C174 VTAIL.n138 B 0.009216f
C175 VTAIL.n139 B 0.020574f
C176 VTAIL.n140 B 0.020574f
C177 VTAIL.n141 B 0.009216f
C178 VTAIL.n142 B 0.008704f
C179 VTAIL.n143 B 0.016198f
C180 VTAIL.n144 B 0.016198f
C181 VTAIL.n145 B 0.008704f
C182 VTAIL.n146 B 0.009216f
C183 VTAIL.n147 B 0.020574f
C184 VTAIL.n148 B 0.020574f
C185 VTAIL.n149 B 0.009216f
C186 VTAIL.n150 B 0.008704f
C187 VTAIL.n151 B 0.016198f
C188 VTAIL.n152 B 0.016198f
C189 VTAIL.n153 B 0.008704f
C190 VTAIL.n154 B 0.008704f
C191 VTAIL.n155 B 0.009216f
C192 VTAIL.n156 B 0.020574f
C193 VTAIL.n157 B 0.020574f
C194 VTAIL.n158 B 0.020574f
C195 VTAIL.n159 B 0.00896f
C196 VTAIL.n160 B 0.008704f
C197 VTAIL.n161 B 0.016198f
C198 VTAIL.n162 B 0.016198f
C199 VTAIL.n163 B 0.008704f
C200 VTAIL.n164 B 0.009216f
C201 VTAIL.n165 B 0.020574f
C202 VTAIL.n166 B 0.04106f
C203 VTAIL.n167 B 0.009216f
C204 VTAIL.n168 B 0.008704f
C205 VTAIL.n169 B 0.036999f
C206 VTAIL.n170 B 0.022604f
C207 VTAIL.n171 B 0.219439f
C208 VTAIL.n172 B 0.020801f
C209 VTAIL.n173 B 0.016198f
C210 VTAIL.n174 B 0.008704f
C211 VTAIL.n175 B 0.020574f
C212 VTAIL.n176 B 0.00896f
C213 VTAIL.n177 B 0.016198f
C214 VTAIL.n178 B 0.009216f
C215 VTAIL.n179 B 0.020574f
C216 VTAIL.n180 B 0.009216f
C217 VTAIL.n181 B 0.016198f
C218 VTAIL.n182 B 0.008704f
C219 VTAIL.n183 B 0.020574f
C220 VTAIL.n184 B 0.009216f
C221 VTAIL.n185 B 0.016198f
C222 VTAIL.n186 B 0.008704f
C223 VTAIL.n187 B 0.020574f
C224 VTAIL.n188 B 0.009216f
C225 VTAIL.n189 B 0.016198f
C226 VTAIL.n190 B 0.008704f
C227 VTAIL.n191 B 0.020574f
C228 VTAIL.n192 B 0.009216f
C229 VTAIL.n193 B 0.016198f
C230 VTAIL.n194 B 0.008704f
C231 VTAIL.n195 B 0.020574f
C232 VTAIL.n196 B 0.009216f
C233 VTAIL.n197 B 1.07913f
C234 VTAIL.n198 B 0.008704f
C235 VTAIL.t6 B 0.033943f
C236 VTAIL.n199 B 0.10703f
C237 VTAIL.n200 B 0.012154f
C238 VTAIL.n201 B 0.01543f
C239 VTAIL.n202 B 0.020574f
C240 VTAIL.n203 B 0.009216f
C241 VTAIL.n204 B 0.008704f
C242 VTAIL.n205 B 0.016198f
C243 VTAIL.n206 B 0.016198f
C244 VTAIL.n207 B 0.008704f
C245 VTAIL.n208 B 0.009216f
C246 VTAIL.n209 B 0.020574f
C247 VTAIL.n210 B 0.020574f
C248 VTAIL.n211 B 0.009216f
C249 VTAIL.n212 B 0.008704f
C250 VTAIL.n213 B 0.016198f
C251 VTAIL.n214 B 0.016198f
C252 VTAIL.n215 B 0.008704f
C253 VTAIL.n216 B 0.009216f
C254 VTAIL.n217 B 0.020574f
C255 VTAIL.n218 B 0.020574f
C256 VTAIL.n219 B 0.009216f
C257 VTAIL.n220 B 0.008704f
C258 VTAIL.n221 B 0.016198f
C259 VTAIL.n222 B 0.016198f
C260 VTAIL.n223 B 0.008704f
C261 VTAIL.n224 B 0.009216f
C262 VTAIL.n225 B 0.020574f
C263 VTAIL.n226 B 0.020574f
C264 VTAIL.n227 B 0.009216f
C265 VTAIL.n228 B 0.008704f
C266 VTAIL.n229 B 0.016198f
C267 VTAIL.n230 B 0.016198f
C268 VTAIL.n231 B 0.008704f
C269 VTAIL.n232 B 0.009216f
C270 VTAIL.n233 B 0.020574f
C271 VTAIL.n234 B 0.020574f
C272 VTAIL.n235 B 0.009216f
C273 VTAIL.n236 B 0.008704f
C274 VTAIL.n237 B 0.016198f
C275 VTAIL.n238 B 0.016198f
C276 VTAIL.n239 B 0.008704f
C277 VTAIL.n240 B 0.008704f
C278 VTAIL.n241 B 0.009216f
C279 VTAIL.n242 B 0.020574f
C280 VTAIL.n243 B 0.020574f
C281 VTAIL.n244 B 0.020574f
C282 VTAIL.n245 B 0.00896f
C283 VTAIL.n246 B 0.008704f
C284 VTAIL.n247 B 0.016198f
C285 VTAIL.n248 B 0.016198f
C286 VTAIL.n249 B 0.008704f
C287 VTAIL.n250 B 0.009216f
C288 VTAIL.n251 B 0.020574f
C289 VTAIL.n252 B 0.04106f
C290 VTAIL.n253 B 0.009216f
C291 VTAIL.n254 B 0.008704f
C292 VTAIL.n255 B 0.036999f
C293 VTAIL.n256 B 0.022604f
C294 VTAIL.n257 B 1.28652f
C295 VTAIL.n258 B 0.020801f
C296 VTAIL.n259 B 0.016198f
C297 VTAIL.n260 B 0.008704f
C298 VTAIL.n261 B 0.020574f
C299 VTAIL.n262 B 0.00896f
C300 VTAIL.n263 B 0.016198f
C301 VTAIL.n264 B 0.00896f
C302 VTAIL.n265 B 0.008704f
C303 VTAIL.n266 B 0.020574f
C304 VTAIL.n267 B 0.020574f
C305 VTAIL.n268 B 0.009216f
C306 VTAIL.n269 B 0.016198f
C307 VTAIL.n270 B 0.008704f
C308 VTAIL.n271 B 0.020574f
C309 VTAIL.n272 B 0.009216f
C310 VTAIL.n273 B 0.016198f
C311 VTAIL.n274 B 0.008704f
C312 VTAIL.n275 B 0.020574f
C313 VTAIL.n276 B 0.009216f
C314 VTAIL.n277 B 0.016198f
C315 VTAIL.n278 B 0.008704f
C316 VTAIL.n279 B 0.020574f
C317 VTAIL.n280 B 0.009216f
C318 VTAIL.n281 B 0.016198f
C319 VTAIL.n282 B 0.008704f
C320 VTAIL.n283 B 0.020574f
C321 VTAIL.n284 B 0.009216f
C322 VTAIL.n285 B 1.07913f
C323 VTAIL.n286 B 0.008704f
C324 VTAIL.t1 B 0.033943f
C325 VTAIL.n287 B 0.10703f
C326 VTAIL.n288 B 0.012154f
C327 VTAIL.n289 B 0.01543f
C328 VTAIL.n290 B 0.020574f
C329 VTAIL.n291 B 0.009216f
C330 VTAIL.n292 B 0.008704f
C331 VTAIL.n293 B 0.016198f
C332 VTAIL.n294 B 0.016198f
C333 VTAIL.n295 B 0.008704f
C334 VTAIL.n296 B 0.009216f
C335 VTAIL.n297 B 0.020574f
C336 VTAIL.n298 B 0.020574f
C337 VTAIL.n299 B 0.009216f
C338 VTAIL.n300 B 0.008704f
C339 VTAIL.n301 B 0.016198f
C340 VTAIL.n302 B 0.016198f
C341 VTAIL.n303 B 0.008704f
C342 VTAIL.n304 B 0.009216f
C343 VTAIL.n305 B 0.020574f
C344 VTAIL.n306 B 0.020574f
C345 VTAIL.n307 B 0.009216f
C346 VTAIL.n308 B 0.008704f
C347 VTAIL.n309 B 0.016198f
C348 VTAIL.n310 B 0.016198f
C349 VTAIL.n311 B 0.008704f
C350 VTAIL.n312 B 0.009216f
C351 VTAIL.n313 B 0.020574f
C352 VTAIL.n314 B 0.020574f
C353 VTAIL.n315 B 0.009216f
C354 VTAIL.n316 B 0.008704f
C355 VTAIL.n317 B 0.016198f
C356 VTAIL.n318 B 0.016198f
C357 VTAIL.n319 B 0.008704f
C358 VTAIL.n320 B 0.009216f
C359 VTAIL.n321 B 0.020574f
C360 VTAIL.n322 B 0.020574f
C361 VTAIL.n323 B 0.009216f
C362 VTAIL.n324 B 0.008704f
C363 VTAIL.n325 B 0.016198f
C364 VTAIL.n326 B 0.016198f
C365 VTAIL.n327 B 0.008704f
C366 VTAIL.n328 B 0.009216f
C367 VTAIL.n329 B 0.020574f
C368 VTAIL.n330 B 0.020574f
C369 VTAIL.n331 B 0.009216f
C370 VTAIL.n332 B 0.008704f
C371 VTAIL.n333 B 0.016198f
C372 VTAIL.n334 B 0.016198f
C373 VTAIL.n335 B 0.008704f
C374 VTAIL.n336 B 0.009216f
C375 VTAIL.n337 B 0.020574f
C376 VTAIL.n338 B 0.04106f
C377 VTAIL.n339 B 0.009216f
C378 VTAIL.n340 B 0.008704f
C379 VTAIL.n341 B 0.036999f
C380 VTAIL.n342 B 0.022604f
C381 VTAIL.n343 B 1.28652f
C382 VTAIL.n344 B 0.020801f
C383 VTAIL.n345 B 0.016198f
C384 VTAIL.n346 B 0.008704f
C385 VTAIL.n347 B 0.020574f
C386 VTAIL.n348 B 0.00896f
C387 VTAIL.n349 B 0.016198f
C388 VTAIL.n350 B 0.00896f
C389 VTAIL.n351 B 0.008704f
C390 VTAIL.n352 B 0.020574f
C391 VTAIL.n353 B 0.020574f
C392 VTAIL.n354 B 0.009216f
C393 VTAIL.n355 B 0.016198f
C394 VTAIL.n356 B 0.008704f
C395 VTAIL.n357 B 0.020574f
C396 VTAIL.n358 B 0.009216f
C397 VTAIL.n359 B 0.016198f
C398 VTAIL.n360 B 0.008704f
C399 VTAIL.n361 B 0.020574f
C400 VTAIL.n362 B 0.009216f
C401 VTAIL.n363 B 0.016198f
C402 VTAIL.n364 B 0.008704f
C403 VTAIL.n365 B 0.020574f
C404 VTAIL.n366 B 0.009216f
C405 VTAIL.n367 B 0.016198f
C406 VTAIL.n368 B 0.008704f
C407 VTAIL.n369 B 0.020574f
C408 VTAIL.n370 B 0.009216f
C409 VTAIL.n371 B 1.07913f
C410 VTAIL.n372 B 0.008704f
C411 VTAIL.t2 B 0.033943f
C412 VTAIL.n373 B 0.10703f
C413 VTAIL.n374 B 0.012154f
C414 VTAIL.n375 B 0.01543f
C415 VTAIL.n376 B 0.020574f
C416 VTAIL.n377 B 0.009216f
C417 VTAIL.n378 B 0.008704f
C418 VTAIL.n379 B 0.016198f
C419 VTAIL.n380 B 0.016198f
C420 VTAIL.n381 B 0.008704f
C421 VTAIL.n382 B 0.009216f
C422 VTAIL.n383 B 0.020574f
C423 VTAIL.n384 B 0.020574f
C424 VTAIL.n385 B 0.009216f
C425 VTAIL.n386 B 0.008704f
C426 VTAIL.n387 B 0.016198f
C427 VTAIL.n388 B 0.016198f
C428 VTAIL.n389 B 0.008704f
C429 VTAIL.n390 B 0.009216f
C430 VTAIL.n391 B 0.020574f
C431 VTAIL.n392 B 0.020574f
C432 VTAIL.n393 B 0.009216f
C433 VTAIL.n394 B 0.008704f
C434 VTAIL.n395 B 0.016198f
C435 VTAIL.n396 B 0.016198f
C436 VTAIL.n397 B 0.008704f
C437 VTAIL.n398 B 0.009216f
C438 VTAIL.n399 B 0.020574f
C439 VTAIL.n400 B 0.020574f
C440 VTAIL.n401 B 0.009216f
C441 VTAIL.n402 B 0.008704f
C442 VTAIL.n403 B 0.016198f
C443 VTAIL.n404 B 0.016198f
C444 VTAIL.n405 B 0.008704f
C445 VTAIL.n406 B 0.009216f
C446 VTAIL.n407 B 0.020574f
C447 VTAIL.n408 B 0.020574f
C448 VTAIL.n409 B 0.009216f
C449 VTAIL.n410 B 0.008704f
C450 VTAIL.n411 B 0.016198f
C451 VTAIL.n412 B 0.016198f
C452 VTAIL.n413 B 0.008704f
C453 VTAIL.n414 B 0.009216f
C454 VTAIL.n415 B 0.020574f
C455 VTAIL.n416 B 0.020574f
C456 VTAIL.n417 B 0.009216f
C457 VTAIL.n418 B 0.008704f
C458 VTAIL.n419 B 0.016198f
C459 VTAIL.n420 B 0.016198f
C460 VTAIL.n421 B 0.008704f
C461 VTAIL.n422 B 0.009216f
C462 VTAIL.n423 B 0.020574f
C463 VTAIL.n424 B 0.04106f
C464 VTAIL.n425 B 0.009216f
C465 VTAIL.n426 B 0.008704f
C466 VTAIL.n427 B 0.036999f
C467 VTAIL.n428 B 0.022604f
C468 VTAIL.n429 B 0.219439f
C469 VTAIL.n430 B 0.020801f
C470 VTAIL.n431 B 0.016198f
C471 VTAIL.n432 B 0.008704f
C472 VTAIL.n433 B 0.020574f
C473 VTAIL.n434 B 0.00896f
C474 VTAIL.n435 B 0.016198f
C475 VTAIL.n436 B 0.00896f
C476 VTAIL.n437 B 0.008704f
C477 VTAIL.n438 B 0.020574f
C478 VTAIL.n439 B 0.020574f
C479 VTAIL.n440 B 0.009216f
C480 VTAIL.n441 B 0.016198f
C481 VTAIL.n442 B 0.008704f
C482 VTAIL.n443 B 0.020574f
C483 VTAIL.n444 B 0.009216f
C484 VTAIL.n445 B 0.016198f
C485 VTAIL.n446 B 0.008704f
C486 VTAIL.n447 B 0.020574f
C487 VTAIL.n448 B 0.009216f
C488 VTAIL.n449 B 0.016198f
C489 VTAIL.n450 B 0.008704f
C490 VTAIL.n451 B 0.020574f
C491 VTAIL.n452 B 0.009216f
C492 VTAIL.n453 B 0.016198f
C493 VTAIL.n454 B 0.008704f
C494 VTAIL.n455 B 0.020574f
C495 VTAIL.n456 B 0.009216f
C496 VTAIL.n457 B 1.07913f
C497 VTAIL.n458 B 0.008704f
C498 VTAIL.t4 B 0.033943f
C499 VTAIL.n459 B 0.10703f
C500 VTAIL.n460 B 0.012154f
C501 VTAIL.n461 B 0.01543f
C502 VTAIL.n462 B 0.020574f
C503 VTAIL.n463 B 0.009216f
C504 VTAIL.n464 B 0.008704f
C505 VTAIL.n465 B 0.016198f
C506 VTAIL.n466 B 0.016198f
C507 VTAIL.n467 B 0.008704f
C508 VTAIL.n468 B 0.009216f
C509 VTAIL.n469 B 0.020574f
C510 VTAIL.n470 B 0.020574f
C511 VTAIL.n471 B 0.009216f
C512 VTAIL.n472 B 0.008704f
C513 VTAIL.n473 B 0.016198f
C514 VTAIL.n474 B 0.016198f
C515 VTAIL.n475 B 0.008704f
C516 VTAIL.n476 B 0.009216f
C517 VTAIL.n477 B 0.020574f
C518 VTAIL.n478 B 0.020574f
C519 VTAIL.n479 B 0.009216f
C520 VTAIL.n480 B 0.008704f
C521 VTAIL.n481 B 0.016198f
C522 VTAIL.n482 B 0.016198f
C523 VTAIL.n483 B 0.008704f
C524 VTAIL.n484 B 0.009216f
C525 VTAIL.n485 B 0.020574f
C526 VTAIL.n486 B 0.020574f
C527 VTAIL.n487 B 0.009216f
C528 VTAIL.n488 B 0.008704f
C529 VTAIL.n489 B 0.016198f
C530 VTAIL.n490 B 0.016198f
C531 VTAIL.n491 B 0.008704f
C532 VTAIL.n492 B 0.009216f
C533 VTAIL.n493 B 0.020574f
C534 VTAIL.n494 B 0.020574f
C535 VTAIL.n495 B 0.009216f
C536 VTAIL.n496 B 0.008704f
C537 VTAIL.n497 B 0.016198f
C538 VTAIL.n498 B 0.016198f
C539 VTAIL.n499 B 0.008704f
C540 VTAIL.n500 B 0.009216f
C541 VTAIL.n501 B 0.020574f
C542 VTAIL.n502 B 0.020574f
C543 VTAIL.n503 B 0.009216f
C544 VTAIL.n504 B 0.008704f
C545 VTAIL.n505 B 0.016198f
C546 VTAIL.n506 B 0.016198f
C547 VTAIL.n507 B 0.008704f
C548 VTAIL.n508 B 0.009216f
C549 VTAIL.n509 B 0.020574f
C550 VTAIL.n510 B 0.04106f
C551 VTAIL.n511 B 0.009216f
C552 VTAIL.n512 B 0.008704f
C553 VTAIL.n513 B 0.036999f
C554 VTAIL.n514 B 0.022604f
C555 VTAIL.n515 B 0.219439f
C556 VTAIL.n516 B 0.020801f
C557 VTAIL.n517 B 0.016198f
C558 VTAIL.n518 B 0.008704f
C559 VTAIL.n519 B 0.020574f
C560 VTAIL.n520 B 0.00896f
C561 VTAIL.n521 B 0.016198f
C562 VTAIL.n522 B 0.00896f
C563 VTAIL.n523 B 0.008704f
C564 VTAIL.n524 B 0.020574f
C565 VTAIL.n525 B 0.020574f
C566 VTAIL.n526 B 0.009216f
C567 VTAIL.n527 B 0.016198f
C568 VTAIL.n528 B 0.008704f
C569 VTAIL.n529 B 0.020574f
C570 VTAIL.n530 B 0.009216f
C571 VTAIL.n531 B 0.016198f
C572 VTAIL.n532 B 0.008704f
C573 VTAIL.n533 B 0.020574f
C574 VTAIL.n534 B 0.009216f
C575 VTAIL.n535 B 0.016198f
C576 VTAIL.n536 B 0.008704f
C577 VTAIL.n537 B 0.020574f
C578 VTAIL.n538 B 0.009216f
C579 VTAIL.n539 B 0.016198f
C580 VTAIL.n540 B 0.008704f
C581 VTAIL.n541 B 0.020574f
C582 VTAIL.n542 B 0.009216f
C583 VTAIL.n543 B 1.07913f
C584 VTAIL.n544 B 0.008704f
C585 VTAIL.t7 B 0.033943f
C586 VTAIL.n545 B 0.10703f
C587 VTAIL.n546 B 0.012154f
C588 VTAIL.n547 B 0.01543f
C589 VTAIL.n548 B 0.020574f
C590 VTAIL.n549 B 0.009216f
C591 VTAIL.n550 B 0.008704f
C592 VTAIL.n551 B 0.016198f
C593 VTAIL.n552 B 0.016198f
C594 VTAIL.n553 B 0.008704f
C595 VTAIL.n554 B 0.009216f
C596 VTAIL.n555 B 0.020574f
C597 VTAIL.n556 B 0.020574f
C598 VTAIL.n557 B 0.009216f
C599 VTAIL.n558 B 0.008704f
C600 VTAIL.n559 B 0.016198f
C601 VTAIL.n560 B 0.016198f
C602 VTAIL.n561 B 0.008704f
C603 VTAIL.n562 B 0.009216f
C604 VTAIL.n563 B 0.020574f
C605 VTAIL.n564 B 0.020574f
C606 VTAIL.n565 B 0.009216f
C607 VTAIL.n566 B 0.008704f
C608 VTAIL.n567 B 0.016198f
C609 VTAIL.n568 B 0.016198f
C610 VTAIL.n569 B 0.008704f
C611 VTAIL.n570 B 0.009216f
C612 VTAIL.n571 B 0.020574f
C613 VTAIL.n572 B 0.020574f
C614 VTAIL.n573 B 0.009216f
C615 VTAIL.n574 B 0.008704f
C616 VTAIL.n575 B 0.016198f
C617 VTAIL.n576 B 0.016198f
C618 VTAIL.n577 B 0.008704f
C619 VTAIL.n578 B 0.009216f
C620 VTAIL.n579 B 0.020574f
C621 VTAIL.n580 B 0.020574f
C622 VTAIL.n581 B 0.009216f
C623 VTAIL.n582 B 0.008704f
C624 VTAIL.n583 B 0.016198f
C625 VTAIL.n584 B 0.016198f
C626 VTAIL.n585 B 0.008704f
C627 VTAIL.n586 B 0.009216f
C628 VTAIL.n587 B 0.020574f
C629 VTAIL.n588 B 0.020574f
C630 VTAIL.n589 B 0.009216f
C631 VTAIL.n590 B 0.008704f
C632 VTAIL.n591 B 0.016198f
C633 VTAIL.n592 B 0.016198f
C634 VTAIL.n593 B 0.008704f
C635 VTAIL.n594 B 0.009216f
C636 VTAIL.n595 B 0.020574f
C637 VTAIL.n596 B 0.04106f
C638 VTAIL.n597 B 0.009216f
C639 VTAIL.n598 B 0.008704f
C640 VTAIL.n599 B 0.036999f
C641 VTAIL.n600 B 0.022604f
C642 VTAIL.n601 B 1.28652f
C643 VTAIL.n602 B 0.020801f
C644 VTAIL.n603 B 0.016198f
C645 VTAIL.n604 B 0.008704f
C646 VTAIL.n605 B 0.020574f
C647 VTAIL.n606 B 0.00896f
C648 VTAIL.n607 B 0.016198f
C649 VTAIL.n608 B 0.009216f
C650 VTAIL.n609 B 0.020574f
C651 VTAIL.n610 B 0.009216f
C652 VTAIL.n611 B 0.016198f
C653 VTAIL.n612 B 0.008704f
C654 VTAIL.n613 B 0.020574f
C655 VTAIL.n614 B 0.009216f
C656 VTAIL.n615 B 0.016198f
C657 VTAIL.n616 B 0.008704f
C658 VTAIL.n617 B 0.020574f
C659 VTAIL.n618 B 0.009216f
C660 VTAIL.n619 B 0.016198f
C661 VTAIL.n620 B 0.008704f
C662 VTAIL.n621 B 0.020574f
C663 VTAIL.n622 B 0.009216f
C664 VTAIL.n623 B 0.016198f
C665 VTAIL.n624 B 0.008704f
C666 VTAIL.n625 B 0.020574f
C667 VTAIL.n626 B 0.009216f
C668 VTAIL.n627 B 1.07913f
C669 VTAIL.n628 B 0.008704f
C670 VTAIL.t0 B 0.033943f
C671 VTAIL.n629 B 0.10703f
C672 VTAIL.n630 B 0.012154f
C673 VTAIL.n631 B 0.01543f
C674 VTAIL.n632 B 0.020574f
C675 VTAIL.n633 B 0.009216f
C676 VTAIL.n634 B 0.008704f
C677 VTAIL.n635 B 0.016198f
C678 VTAIL.n636 B 0.016198f
C679 VTAIL.n637 B 0.008704f
C680 VTAIL.n638 B 0.009216f
C681 VTAIL.n639 B 0.020574f
C682 VTAIL.n640 B 0.020574f
C683 VTAIL.n641 B 0.009216f
C684 VTAIL.n642 B 0.008704f
C685 VTAIL.n643 B 0.016198f
C686 VTAIL.n644 B 0.016198f
C687 VTAIL.n645 B 0.008704f
C688 VTAIL.n646 B 0.009216f
C689 VTAIL.n647 B 0.020574f
C690 VTAIL.n648 B 0.020574f
C691 VTAIL.n649 B 0.009216f
C692 VTAIL.n650 B 0.008704f
C693 VTAIL.n651 B 0.016198f
C694 VTAIL.n652 B 0.016198f
C695 VTAIL.n653 B 0.008704f
C696 VTAIL.n654 B 0.009216f
C697 VTAIL.n655 B 0.020574f
C698 VTAIL.n656 B 0.020574f
C699 VTAIL.n657 B 0.009216f
C700 VTAIL.n658 B 0.008704f
C701 VTAIL.n659 B 0.016198f
C702 VTAIL.n660 B 0.016198f
C703 VTAIL.n661 B 0.008704f
C704 VTAIL.n662 B 0.009216f
C705 VTAIL.n663 B 0.020574f
C706 VTAIL.n664 B 0.020574f
C707 VTAIL.n665 B 0.009216f
C708 VTAIL.n666 B 0.008704f
C709 VTAIL.n667 B 0.016198f
C710 VTAIL.n668 B 0.016198f
C711 VTAIL.n669 B 0.008704f
C712 VTAIL.n670 B 0.008704f
C713 VTAIL.n671 B 0.009216f
C714 VTAIL.n672 B 0.020574f
C715 VTAIL.n673 B 0.020574f
C716 VTAIL.n674 B 0.020574f
C717 VTAIL.n675 B 0.00896f
C718 VTAIL.n676 B 0.008704f
C719 VTAIL.n677 B 0.016198f
C720 VTAIL.n678 B 0.016198f
C721 VTAIL.n679 B 0.008704f
C722 VTAIL.n680 B 0.009216f
C723 VTAIL.n681 B 0.020574f
C724 VTAIL.n682 B 0.04106f
C725 VTAIL.n683 B 0.009216f
C726 VTAIL.n684 B 0.008704f
C727 VTAIL.n685 B 0.036999f
C728 VTAIL.n686 B 0.022604f
C729 VTAIL.n687 B 1.19281f
C730 VP.t3 B 3.0683f
C731 VP.n0 B 1.13306f
C732 VP.n1 B 0.019718f
C733 VP.n2 B 0.038984f
C734 VP.n3 B 0.019718f
C735 VP.n4 B 0.036566f
C736 VP.t1 B 3.37426f
C737 VP.t0 B 3.36256f
C738 VP.n5 B 3.41217f
C739 VP.n6 B 1.27058f
C740 VP.t2 B 3.0683f
C741 VP.n7 B 1.13306f
C742 VP.n8 B 0.019056f
C743 VP.n9 B 0.03182f
C744 VP.n10 B 0.019718f
C745 VP.n11 B 0.019718f
C746 VP.n12 B 0.036566f
C747 VP.n13 B 0.038984f
C748 VP.n14 B 0.015926f
C749 VP.n15 B 0.019718f
C750 VP.n16 B 0.019718f
C751 VP.n17 B 0.019718f
C752 VP.n18 B 0.036566f
C753 VP.n19 B 0.036566f
C754 VP.n20 B 0.019056f
C755 VP.n21 B 0.03182f
C756 VP.n22 B 0.060545f
.ends

