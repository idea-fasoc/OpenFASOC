* NGSPICE file created from diff_pair_sample_1484.ext - technology: sky130A

.subckt diff_pair_sample_1484 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=3.5646 ps=19.06 w=9.14 l=0.4
X1 B.t11 B.t9 B.t10 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=0 ps=0 w=9.14 l=0.4
X2 B.t8 B.t6 B.t7 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=0 ps=0 w=9.14 l=0.4
X3 B.t5 B.t3 B.t4 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=0 ps=0 w=9.14 l=0.4
X4 VDD2.t1 VN.t0 VTAIL.t0 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=3.5646 ps=19.06 w=9.14 l=0.4
X5 B.t2 B.t0 B.t1 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=0 ps=0 w=9.14 l=0.4
X6 VDD2.t0 VN.t1 VTAIL.t1 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=3.5646 ps=19.06 w=9.14 l=0.4
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n1262_n2800# sky130_fd_pr__pfet_01v8 ad=3.5646 pd=19.06 as=3.5646 ps=19.06 w=9.14 l=0.4
R0 VP.n0 VP.t1 848.068
R1 VP.n0 VP.t0 811.399
R2 VP VP.n0 0.0516364
R3 VTAIL.n2 VTAIL.t3 64.7354
R4 VTAIL.n1 VTAIL.t1 64.7353
R5 VTAIL.n3 VTAIL.t0 64.7352
R6 VTAIL.n0 VTAIL.t2 64.7352
R7 VTAIL.n1 VTAIL.n0 21.5221
R8 VTAIL.n3 VTAIL.n2 20.8927
R9 VTAIL.n2 VTAIL.n1 0.784983
R10 VTAIL VTAIL.n0 0.685845
R11 VTAIL VTAIL.n3 0.0996379
R12 VDD1 VDD1.t1 114.91
R13 VDD1 VDD1.t0 81.6297
R14 B.n174 B.t9 760.106
R15 B.n81 B.t0 760.106
R16 B.n33 B.t3 760.106
R17 B.n26 B.t6 760.106
R18 B.n243 B.n64 585
R19 B.n242 B.n241 585
R20 B.n240 B.n65 585
R21 B.n239 B.n238 585
R22 B.n237 B.n66 585
R23 B.n236 B.n235 585
R24 B.n234 B.n67 585
R25 B.n233 B.n232 585
R26 B.n231 B.n68 585
R27 B.n230 B.n229 585
R28 B.n228 B.n69 585
R29 B.n227 B.n226 585
R30 B.n225 B.n70 585
R31 B.n224 B.n223 585
R32 B.n222 B.n71 585
R33 B.n221 B.n220 585
R34 B.n219 B.n72 585
R35 B.n218 B.n217 585
R36 B.n216 B.n73 585
R37 B.n215 B.n214 585
R38 B.n213 B.n74 585
R39 B.n212 B.n211 585
R40 B.n210 B.n75 585
R41 B.n209 B.n208 585
R42 B.n207 B.n76 585
R43 B.n206 B.n205 585
R44 B.n204 B.n77 585
R45 B.n203 B.n202 585
R46 B.n201 B.n78 585
R47 B.n200 B.n199 585
R48 B.n198 B.n79 585
R49 B.n197 B.n196 585
R50 B.n195 B.n80 585
R51 B.n193 B.n192 585
R52 B.n191 B.n83 585
R53 B.n190 B.n189 585
R54 B.n188 B.n84 585
R55 B.n187 B.n186 585
R56 B.n185 B.n85 585
R57 B.n184 B.n183 585
R58 B.n182 B.n86 585
R59 B.n181 B.n180 585
R60 B.n179 B.n87 585
R61 B.n178 B.n177 585
R62 B.n173 B.n88 585
R63 B.n172 B.n171 585
R64 B.n170 B.n89 585
R65 B.n169 B.n168 585
R66 B.n167 B.n90 585
R67 B.n166 B.n165 585
R68 B.n164 B.n91 585
R69 B.n163 B.n162 585
R70 B.n161 B.n92 585
R71 B.n160 B.n159 585
R72 B.n158 B.n93 585
R73 B.n157 B.n156 585
R74 B.n155 B.n94 585
R75 B.n154 B.n153 585
R76 B.n152 B.n95 585
R77 B.n151 B.n150 585
R78 B.n149 B.n96 585
R79 B.n148 B.n147 585
R80 B.n146 B.n97 585
R81 B.n145 B.n144 585
R82 B.n143 B.n98 585
R83 B.n142 B.n141 585
R84 B.n140 B.n99 585
R85 B.n139 B.n138 585
R86 B.n137 B.n100 585
R87 B.n136 B.n135 585
R88 B.n134 B.n101 585
R89 B.n133 B.n132 585
R90 B.n131 B.n102 585
R91 B.n130 B.n129 585
R92 B.n128 B.n103 585
R93 B.n127 B.n126 585
R94 B.n245 B.n244 585
R95 B.n246 B.n63 585
R96 B.n248 B.n247 585
R97 B.n249 B.n62 585
R98 B.n251 B.n250 585
R99 B.n252 B.n61 585
R100 B.n254 B.n253 585
R101 B.n255 B.n60 585
R102 B.n257 B.n256 585
R103 B.n258 B.n59 585
R104 B.n260 B.n259 585
R105 B.n261 B.n58 585
R106 B.n263 B.n262 585
R107 B.n264 B.n57 585
R108 B.n266 B.n265 585
R109 B.n267 B.n56 585
R110 B.n269 B.n268 585
R111 B.n270 B.n55 585
R112 B.n272 B.n271 585
R113 B.n273 B.n54 585
R114 B.n275 B.n274 585
R115 B.n276 B.n53 585
R116 B.n278 B.n277 585
R117 B.n279 B.n52 585
R118 B.n281 B.n280 585
R119 B.n282 B.n51 585
R120 B.n397 B.n8 585
R121 B.n396 B.n395 585
R122 B.n394 B.n9 585
R123 B.n393 B.n392 585
R124 B.n391 B.n10 585
R125 B.n390 B.n389 585
R126 B.n388 B.n11 585
R127 B.n387 B.n386 585
R128 B.n385 B.n12 585
R129 B.n384 B.n383 585
R130 B.n382 B.n13 585
R131 B.n381 B.n380 585
R132 B.n379 B.n14 585
R133 B.n378 B.n377 585
R134 B.n376 B.n15 585
R135 B.n375 B.n374 585
R136 B.n373 B.n16 585
R137 B.n372 B.n371 585
R138 B.n370 B.n17 585
R139 B.n369 B.n368 585
R140 B.n367 B.n18 585
R141 B.n366 B.n365 585
R142 B.n364 B.n19 585
R143 B.n363 B.n362 585
R144 B.n361 B.n20 585
R145 B.n360 B.n359 585
R146 B.n358 B.n21 585
R147 B.n357 B.n356 585
R148 B.n355 B.n22 585
R149 B.n354 B.n353 585
R150 B.n352 B.n23 585
R151 B.n351 B.n350 585
R152 B.n349 B.n24 585
R153 B.n348 B.n347 585
R154 B.n346 B.n25 585
R155 B.n345 B.n344 585
R156 B.n343 B.n29 585
R157 B.n342 B.n341 585
R158 B.n340 B.n30 585
R159 B.n339 B.n338 585
R160 B.n337 B.n31 585
R161 B.n336 B.n335 585
R162 B.n334 B.n32 585
R163 B.n332 B.n331 585
R164 B.n330 B.n35 585
R165 B.n329 B.n328 585
R166 B.n327 B.n36 585
R167 B.n326 B.n325 585
R168 B.n324 B.n37 585
R169 B.n323 B.n322 585
R170 B.n321 B.n38 585
R171 B.n320 B.n319 585
R172 B.n318 B.n39 585
R173 B.n317 B.n316 585
R174 B.n315 B.n40 585
R175 B.n314 B.n313 585
R176 B.n312 B.n41 585
R177 B.n311 B.n310 585
R178 B.n309 B.n42 585
R179 B.n308 B.n307 585
R180 B.n306 B.n43 585
R181 B.n305 B.n304 585
R182 B.n303 B.n44 585
R183 B.n302 B.n301 585
R184 B.n300 B.n45 585
R185 B.n299 B.n298 585
R186 B.n297 B.n46 585
R187 B.n296 B.n295 585
R188 B.n294 B.n47 585
R189 B.n293 B.n292 585
R190 B.n291 B.n48 585
R191 B.n290 B.n289 585
R192 B.n288 B.n49 585
R193 B.n287 B.n286 585
R194 B.n285 B.n50 585
R195 B.n284 B.n283 585
R196 B.n399 B.n398 585
R197 B.n400 B.n7 585
R198 B.n402 B.n401 585
R199 B.n403 B.n6 585
R200 B.n405 B.n404 585
R201 B.n406 B.n5 585
R202 B.n408 B.n407 585
R203 B.n409 B.n4 585
R204 B.n411 B.n410 585
R205 B.n412 B.n3 585
R206 B.n414 B.n413 585
R207 B.n415 B.n0 585
R208 B.n2 B.n1 585
R209 B.n110 B.n109 585
R210 B.n112 B.n111 585
R211 B.n113 B.n108 585
R212 B.n115 B.n114 585
R213 B.n116 B.n107 585
R214 B.n118 B.n117 585
R215 B.n119 B.n106 585
R216 B.n121 B.n120 585
R217 B.n122 B.n105 585
R218 B.n124 B.n123 585
R219 B.n125 B.n104 585
R220 B.n127 B.n104 492.5
R221 B.n245 B.n64 492.5
R222 B.n283 B.n282 492.5
R223 B.n398 B.n397 492.5
R224 B.n417 B.n416 256.663
R225 B.n416 B.n415 235.042
R226 B.n416 B.n2 235.042
R227 B.n128 B.n127 163.367
R228 B.n129 B.n128 163.367
R229 B.n129 B.n102 163.367
R230 B.n133 B.n102 163.367
R231 B.n134 B.n133 163.367
R232 B.n135 B.n134 163.367
R233 B.n135 B.n100 163.367
R234 B.n139 B.n100 163.367
R235 B.n140 B.n139 163.367
R236 B.n141 B.n140 163.367
R237 B.n141 B.n98 163.367
R238 B.n145 B.n98 163.367
R239 B.n146 B.n145 163.367
R240 B.n147 B.n146 163.367
R241 B.n147 B.n96 163.367
R242 B.n151 B.n96 163.367
R243 B.n152 B.n151 163.367
R244 B.n153 B.n152 163.367
R245 B.n153 B.n94 163.367
R246 B.n157 B.n94 163.367
R247 B.n158 B.n157 163.367
R248 B.n159 B.n158 163.367
R249 B.n159 B.n92 163.367
R250 B.n163 B.n92 163.367
R251 B.n164 B.n163 163.367
R252 B.n165 B.n164 163.367
R253 B.n165 B.n90 163.367
R254 B.n169 B.n90 163.367
R255 B.n170 B.n169 163.367
R256 B.n171 B.n170 163.367
R257 B.n171 B.n88 163.367
R258 B.n178 B.n88 163.367
R259 B.n179 B.n178 163.367
R260 B.n180 B.n179 163.367
R261 B.n180 B.n86 163.367
R262 B.n184 B.n86 163.367
R263 B.n185 B.n184 163.367
R264 B.n186 B.n185 163.367
R265 B.n186 B.n84 163.367
R266 B.n190 B.n84 163.367
R267 B.n191 B.n190 163.367
R268 B.n192 B.n191 163.367
R269 B.n192 B.n80 163.367
R270 B.n197 B.n80 163.367
R271 B.n198 B.n197 163.367
R272 B.n199 B.n198 163.367
R273 B.n199 B.n78 163.367
R274 B.n203 B.n78 163.367
R275 B.n204 B.n203 163.367
R276 B.n205 B.n204 163.367
R277 B.n205 B.n76 163.367
R278 B.n209 B.n76 163.367
R279 B.n210 B.n209 163.367
R280 B.n211 B.n210 163.367
R281 B.n211 B.n74 163.367
R282 B.n215 B.n74 163.367
R283 B.n216 B.n215 163.367
R284 B.n217 B.n216 163.367
R285 B.n217 B.n72 163.367
R286 B.n221 B.n72 163.367
R287 B.n222 B.n221 163.367
R288 B.n223 B.n222 163.367
R289 B.n223 B.n70 163.367
R290 B.n227 B.n70 163.367
R291 B.n228 B.n227 163.367
R292 B.n229 B.n228 163.367
R293 B.n229 B.n68 163.367
R294 B.n233 B.n68 163.367
R295 B.n234 B.n233 163.367
R296 B.n235 B.n234 163.367
R297 B.n235 B.n66 163.367
R298 B.n239 B.n66 163.367
R299 B.n240 B.n239 163.367
R300 B.n241 B.n240 163.367
R301 B.n241 B.n64 163.367
R302 B.n282 B.n281 163.367
R303 B.n281 B.n52 163.367
R304 B.n277 B.n52 163.367
R305 B.n277 B.n276 163.367
R306 B.n276 B.n275 163.367
R307 B.n275 B.n54 163.367
R308 B.n271 B.n54 163.367
R309 B.n271 B.n270 163.367
R310 B.n270 B.n269 163.367
R311 B.n269 B.n56 163.367
R312 B.n265 B.n56 163.367
R313 B.n265 B.n264 163.367
R314 B.n264 B.n263 163.367
R315 B.n263 B.n58 163.367
R316 B.n259 B.n58 163.367
R317 B.n259 B.n258 163.367
R318 B.n258 B.n257 163.367
R319 B.n257 B.n60 163.367
R320 B.n253 B.n60 163.367
R321 B.n253 B.n252 163.367
R322 B.n252 B.n251 163.367
R323 B.n251 B.n62 163.367
R324 B.n247 B.n62 163.367
R325 B.n247 B.n246 163.367
R326 B.n246 B.n245 163.367
R327 B.n397 B.n396 163.367
R328 B.n396 B.n9 163.367
R329 B.n392 B.n9 163.367
R330 B.n392 B.n391 163.367
R331 B.n391 B.n390 163.367
R332 B.n390 B.n11 163.367
R333 B.n386 B.n11 163.367
R334 B.n386 B.n385 163.367
R335 B.n385 B.n384 163.367
R336 B.n384 B.n13 163.367
R337 B.n380 B.n13 163.367
R338 B.n380 B.n379 163.367
R339 B.n379 B.n378 163.367
R340 B.n378 B.n15 163.367
R341 B.n374 B.n15 163.367
R342 B.n374 B.n373 163.367
R343 B.n373 B.n372 163.367
R344 B.n372 B.n17 163.367
R345 B.n368 B.n17 163.367
R346 B.n368 B.n367 163.367
R347 B.n367 B.n366 163.367
R348 B.n366 B.n19 163.367
R349 B.n362 B.n19 163.367
R350 B.n362 B.n361 163.367
R351 B.n361 B.n360 163.367
R352 B.n360 B.n21 163.367
R353 B.n356 B.n21 163.367
R354 B.n356 B.n355 163.367
R355 B.n355 B.n354 163.367
R356 B.n354 B.n23 163.367
R357 B.n350 B.n23 163.367
R358 B.n350 B.n349 163.367
R359 B.n349 B.n348 163.367
R360 B.n348 B.n25 163.367
R361 B.n344 B.n25 163.367
R362 B.n344 B.n343 163.367
R363 B.n343 B.n342 163.367
R364 B.n342 B.n30 163.367
R365 B.n338 B.n30 163.367
R366 B.n338 B.n337 163.367
R367 B.n337 B.n336 163.367
R368 B.n336 B.n32 163.367
R369 B.n331 B.n32 163.367
R370 B.n331 B.n330 163.367
R371 B.n330 B.n329 163.367
R372 B.n329 B.n36 163.367
R373 B.n325 B.n36 163.367
R374 B.n325 B.n324 163.367
R375 B.n324 B.n323 163.367
R376 B.n323 B.n38 163.367
R377 B.n319 B.n38 163.367
R378 B.n319 B.n318 163.367
R379 B.n318 B.n317 163.367
R380 B.n317 B.n40 163.367
R381 B.n313 B.n40 163.367
R382 B.n313 B.n312 163.367
R383 B.n312 B.n311 163.367
R384 B.n311 B.n42 163.367
R385 B.n307 B.n42 163.367
R386 B.n307 B.n306 163.367
R387 B.n306 B.n305 163.367
R388 B.n305 B.n44 163.367
R389 B.n301 B.n44 163.367
R390 B.n301 B.n300 163.367
R391 B.n300 B.n299 163.367
R392 B.n299 B.n46 163.367
R393 B.n295 B.n46 163.367
R394 B.n295 B.n294 163.367
R395 B.n294 B.n293 163.367
R396 B.n293 B.n48 163.367
R397 B.n289 B.n48 163.367
R398 B.n289 B.n288 163.367
R399 B.n288 B.n287 163.367
R400 B.n287 B.n50 163.367
R401 B.n283 B.n50 163.367
R402 B.n398 B.n7 163.367
R403 B.n402 B.n7 163.367
R404 B.n403 B.n402 163.367
R405 B.n404 B.n403 163.367
R406 B.n404 B.n5 163.367
R407 B.n408 B.n5 163.367
R408 B.n409 B.n408 163.367
R409 B.n410 B.n409 163.367
R410 B.n410 B.n3 163.367
R411 B.n414 B.n3 163.367
R412 B.n415 B.n414 163.367
R413 B.n110 B.n2 163.367
R414 B.n111 B.n110 163.367
R415 B.n111 B.n108 163.367
R416 B.n115 B.n108 163.367
R417 B.n116 B.n115 163.367
R418 B.n117 B.n116 163.367
R419 B.n117 B.n106 163.367
R420 B.n121 B.n106 163.367
R421 B.n122 B.n121 163.367
R422 B.n123 B.n122 163.367
R423 B.n123 B.n104 163.367
R424 B.n81 B.t1 128.014
R425 B.n33 B.t5 128.014
R426 B.n174 B.t10 128.005
R427 B.n26 B.t8 128.005
R428 B.n82 B.t2 113.858
R429 B.n34 B.t4 113.858
R430 B.n175 B.t11 113.847
R431 B.n27 B.t7 113.847
R432 B.n176 B.n175 59.5399
R433 B.n194 B.n82 59.5399
R434 B.n333 B.n34 59.5399
R435 B.n28 B.n27 59.5399
R436 B.n399 B.n8 32.0005
R437 B.n284 B.n51 32.0005
R438 B.n244 B.n243 32.0005
R439 B.n126 B.n125 32.0005
R440 B B.n417 18.0485
R441 B.n175 B.n174 14.1581
R442 B.n82 B.n81 14.1581
R443 B.n34 B.n33 14.1581
R444 B.n27 B.n26 14.1581
R445 B.n400 B.n399 10.6151
R446 B.n401 B.n400 10.6151
R447 B.n401 B.n6 10.6151
R448 B.n405 B.n6 10.6151
R449 B.n406 B.n405 10.6151
R450 B.n407 B.n406 10.6151
R451 B.n407 B.n4 10.6151
R452 B.n411 B.n4 10.6151
R453 B.n412 B.n411 10.6151
R454 B.n413 B.n412 10.6151
R455 B.n413 B.n0 10.6151
R456 B.n395 B.n8 10.6151
R457 B.n395 B.n394 10.6151
R458 B.n394 B.n393 10.6151
R459 B.n393 B.n10 10.6151
R460 B.n389 B.n10 10.6151
R461 B.n389 B.n388 10.6151
R462 B.n388 B.n387 10.6151
R463 B.n387 B.n12 10.6151
R464 B.n383 B.n12 10.6151
R465 B.n383 B.n382 10.6151
R466 B.n382 B.n381 10.6151
R467 B.n381 B.n14 10.6151
R468 B.n377 B.n14 10.6151
R469 B.n377 B.n376 10.6151
R470 B.n376 B.n375 10.6151
R471 B.n375 B.n16 10.6151
R472 B.n371 B.n16 10.6151
R473 B.n371 B.n370 10.6151
R474 B.n370 B.n369 10.6151
R475 B.n369 B.n18 10.6151
R476 B.n365 B.n18 10.6151
R477 B.n365 B.n364 10.6151
R478 B.n364 B.n363 10.6151
R479 B.n363 B.n20 10.6151
R480 B.n359 B.n20 10.6151
R481 B.n359 B.n358 10.6151
R482 B.n358 B.n357 10.6151
R483 B.n357 B.n22 10.6151
R484 B.n353 B.n22 10.6151
R485 B.n353 B.n352 10.6151
R486 B.n352 B.n351 10.6151
R487 B.n351 B.n24 10.6151
R488 B.n347 B.n346 10.6151
R489 B.n346 B.n345 10.6151
R490 B.n345 B.n29 10.6151
R491 B.n341 B.n29 10.6151
R492 B.n341 B.n340 10.6151
R493 B.n340 B.n339 10.6151
R494 B.n339 B.n31 10.6151
R495 B.n335 B.n31 10.6151
R496 B.n335 B.n334 10.6151
R497 B.n332 B.n35 10.6151
R498 B.n328 B.n35 10.6151
R499 B.n328 B.n327 10.6151
R500 B.n327 B.n326 10.6151
R501 B.n326 B.n37 10.6151
R502 B.n322 B.n37 10.6151
R503 B.n322 B.n321 10.6151
R504 B.n321 B.n320 10.6151
R505 B.n320 B.n39 10.6151
R506 B.n316 B.n39 10.6151
R507 B.n316 B.n315 10.6151
R508 B.n315 B.n314 10.6151
R509 B.n314 B.n41 10.6151
R510 B.n310 B.n41 10.6151
R511 B.n310 B.n309 10.6151
R512 B.n309 B.n308 10.6151
R513 B.n308 B.n43 10.6151
R514 B.n304 B.n43 10.6151
R515 B.n304 B.n303 10.6151
R516 B.n303 B.n302 10.6151
R517 B.n302 B.n45 10.6151
R518 B.n298 B.n45 10.6151
R519 B.n298 B.n297 10.6151
R520 B.n297 B.n296 10.6151
R521 B.n296 B.n47 10.6151
R522 B.n292 B.n47 10.6151
R523 B.n292 B.n291 10.6151
R524 B.n291 B.n290 10.6151
R525 B.n290 B.n49 10.6151
R526 B.n286 B.n49 10.6151
R527 B.n286 B.n285 10.6151
R528 B.n285 B.n284 10.6151
R529 B.n280 B.n51 10.6151
R530 B.n280 B.n279 10.6151
R531 B.n279 B.n278 10.6151
R532 B.n278 B.n53 10.6151
R533 B.n274 B.n53 10.6151
R534 B.n274 B.n273 10.6151
R535 B.n273 B.n272 10.6151
R536 B.n272 B.n55 10.6151
R537 B.n268 B.n55 10.6151
R538 B.n268 B.n267 10.6151
R539 B.n267 B.n266 10.6151
R540 B.n266 B.n57 10.6151
R541 B.n262 B.n57 10.6151
R542 B.n262 B.n261 10.6151
R543 B.n261 B.n260 10.6151
R544 B.n260 B.n59 10.6151
R545 B.n256 B.n59 10.6151
R546 B.n256 B.n255 10.6151
R547 B.n255 B.n254 10.6151
R548 B.n254 B.n61 10.6151
R549 B.n250 B.n61 10.6151
R550 B.n250 B.n249 10.6151
R551 B.n249 B.n248 10.6151
R552 B.n248 B.n63 10.6151
R553 B.n244 B.n63 10.6151
R554 B.n109 B.n1 10.6151
R555 B.n112 B.n109 10.6151
R556 B.n113 B.n112 10.6151
R557 B.n114 B.n113 10.6151
R558 B.n114 B.n107 10.6151
R559 B.n118 B.n107 10.6151
R560 B.n119 B.n118 10.6151
R561 B.n120 B.n119 10.6151
R562 B.n120 B.n105 10.6151
R563 B.n124 B.n105 10.6151
R564 B.n125 B.n124 10.6151
R565 B.n126 B.n103 10.6151
R566 B.n130 B.n103 10.6151
R567 B.n131 B.n130 10.6151
R568 B.n132 B.n131 10.6151
R569 B.n132 B.n101 10.6151
R570 B.n136 B.n101 10.6151
R571 B.n137 B.n136 10.6151
R572 B.n138 B.n137 10.6151
R573 B.n138 B.n99 10.6151
R574 B.n142 B.n99 10.6151
R575 B.n143 B.n142 10.6151
R576 B.n144 B.n143 10.6151
R577 B.n144 B.n97 10.6151
R578 B.n148 B.n97 10.6151
R579 B.n149 B.n148 10.6151
R580 B.n150 B.n149 10.6151
R581 B.n150 B.n95 10.6151
R582 B.n154 B.n95 10.6151
R583 B.n155 B.n154 10.6151
R584 B.n156 B.n155 10.6151
R585 B.n156 B.n93 10.6151
R586 B.n160 B.n93 10.6151
R587 B.n161 B.n160 10.6151
R588 B.n162 B.n161 10.6151
R589 B.n162 B.n91 10.6151
R590 B.n166 B.n91 10.6151
R591 B.n167 B.n166 10.6151
R592 B.n168 B.n167 10.6151
R593 B.n168 B.n89 10.6151
R594 B.n172 B.n89 10.6151
R595 B.n173 B.n172 10.6151
R596 B.n177 B.n173 10.6151
R597 B.n181 B.n87 10.6151
R598 B.n182 B.n181 10.6151
R599 B.n183 B.n182 10.6151
R600 B.n183 B.n85 10.6151
R601 B.n187 B.n85 10.6151
R602 B.n188 B.n187 10.6151
R603 B.n189 B.n188 10.6151
R604 B.n189 B.n83 10.6151
R605 B.n193 B.n83 10.6151
R606 B.n196 B.n195 10.6151
R607 B.n196 B.n79 10.6151
R608 B.n200 B.n79 10.6151
R609 B.n201 B.n200 10.6151
R610 B.n202 B.n201 10.6151
R611 B.n202 B.n77 10.6151
R612 B.n206 B.n77 10.6151
R613 B.n207 B.n206 10.6151
R614 B.n208 B.n207 10.6151
R615 B.n208 B.n75 10.6151
R616 B.n212 B.n75 10.6151
R617 B.n213 B.n212 10.6151
R618 B.n214 B.n213 10.6151
R619 B.n214 B.n73 10.6151
R620 B.n218 B.n73 10.6151
R621 B.n219 B.n218 10.6151
R622 B.n220 B.n219 10.6151
R623 B.n220 B.n71 10.6151
R624 B.n224 B.n71 10.6151
R625 B.n225 B.n224 10.6151
R626 B.n226 B.n225 10.6151
R627 B.n226 B.n69 10.6151
R628 B.n230 B.n69 10.6151
R629 B.n231 B.n230 10.6151
R630 B.n232 B.n231 10.6151
R631 B.n232 B.n67 10.6151
R632 B.n236 B.n67 10.6151
R633 B.n237 B.n236 10.6151
R634 B.n238 B.n237 10.6151
R635 B.n238 B.n65 10.6151
R636 B.n242 B.n65 10.6151
R637 B.n243 B.n242 10.6151
R638 B.n28 B.n24 8.74196
R639 B.n333 B.n332 8.74196
R640 B.n177 B.n176 8.74196
R641 B.n195 B.n194 8.74196
R642 B.n417 B.n0 8.11757
R643 B.n417 B.n1 8.11757
R644 B.n347 B.n28 1.87367
R645 B.n334 B.n333 1.87367
R646 B.n176 B.n87 1.87367
R647 B.n194 B.n193 1.87367
R648 VN VN.t1 848.449
R649 VN VN.t0 811.449
R650 VDD2.n0 VDD2.t1 114.228
R651 VDD2.n0 VDD2.t0 81.4141
R652 VDD2 VDD2.n0 0.216017
C0 VDD2 VDD1 0.434099f
C1 VDD1 w_n1262_n2800# 1.32624f
C2 VDD2 B 1.16861f
C3 B w_n1262_n2800# 5.63331f
C4 VDD2 VTAIL 5.22084f
C5 VTAIL w_n1262_n2800# 2.49283f
C6 VDD1 VN 0.148119f
C7 VN B 0.639739f
C8 VTAIL VN 0.849979f
C9 VDD1 B 1.15609f
C10 VDD2 VP 0.24174f
C11 VP w_n1262_n2800# 1.66915f
C12 VTAIL VDD1 5.18843f
C13 VTAIL B 2.04769f
C14 VN VP 3.89833f
C15 VDD2 w_n1262_n2800# 1.3279f
C16 VDD1 VP 1.36866f
C17 VDD2 VN 1.27879f
C18 VP B 0.887402f
C19 VN w_n1262_n2800# 1.51314f
C20 VTAIL VP 0.86455f
C21 VDD2 VSUBS 0.62624f
C22 VDD1 VSUBS 3.128521f
C23 VTAIL VSUBS 0.236907f
C24 VN VSUBS 4.32808f
C25 VP VSUBS 0.915094f
C26 B VSUBS 2.035697f
C27 w_n1262_n2800# VSUBS 43.7207f
C28 VDD2.t1 VSUBS 1.57509f
C29 VDD2.t0 VSUBS 1.24467f
C30 VDD2.n0 VSUBS 2.34924f
C31 VN.t0 VSUBS 0.456456f
C32 VN.t1 VSUBS 0.520728f
C33 B.n0 VSUBS 0.007102f
C34 B.n1 VSUBS 0.007102f
C35 B.n2 VSUBS 0.010504f
C36 B.n3 VSUBS 0.008049f
C37 B.n4 VSUBS 0.008049f
C38 B.n5 VSUBS 0.008049f
C39 B.n6 VSUBS 0.008049f
C40 B.n7 VSUBS 0.008049f
C41 B.n8 VSUBS 0.018928f
C42 B.n9 VSUBS 0.008049f
C43 B.n10 VSUBS 0.008049f
C44 B.n11 VSUBS 0.008049f
C45 B.n12 VSUBS 0.008049f
C46 B.n13 VSUBS 0.008049f
C47 B.n14 VSUBS 0.008049f
C48 B.n15 VSUBS 0.008049f
C49 B.n16 VSUBS 0.008049f
C50 B.n17 VSUBS 0.008049f
C51 B.n18 VSUBS 0.008049f
C52 B.n19 VSUBS 0.008049f
C53 B.n20 VSUBS 0.008049f
C54 B.n21 VSUBS 0.008049f
C55 B.n22 VSUBS 0.008049f
C56 B.n23 VSUBS 0.008049f
C57 B.n24 VSUBS 0.007339f
C58 B.n25 VSUBS 0.008049f
C59 B.t7 VSUBS 0.331025f
C60 B.t8 VSUBS 0.337701f
C61 B.t6 VSUBS 0.169881f
C62 B.n26 VSUBS 0.108148f
C63 B.n27 VSUBS 0.071836f
C64 B.n28 VSUBS 0.018649f
C65 B.n29 VSUBS 0.008049f
C66 B.n30 VSUBS 0.008049f
C67 B.n31 VSUBS 0.008049f
C68 B.n32 VSUBS 0.008049f
C69 B.t4 VSUBS 0.331022f
C70 B.t5 VSUBS 0.337697f
C71 B.t3 VSUBS 0.169881f
C72 B.n33 VSUBS 0.108151f
C73 B.n34 VSUBS 0.071839f
C74 B.n35 VSUBS 0.008049f
C75 B.n36 VSUBS 0.008049f
C76 B.n37 VSUBS 0.008049f
C77 B.n38 VSUBS 0.008049f
C78 B.n39 VSUBS 0.008049f
C79 B.n40 VSUBS 0.008049f
C80 B.n41 VSUBS 0.008049f
C81 B.n42 VSUBS 0.008049f
C82 B.n43 VSUBS 0.008049f
C83 B.n44 VSUBS 0.008049f
C84 B.n45 VSUBS 0.008049f
C85 B.n46 VSUBS 0.008049f
C86 B.n47 VSUBS 0.008049f
C87 B.n48 VSUBS 0.008049f
C88 B.n49 VSUBS 0.008049f
C89 B.n50 VSUBS 0.008049f
C90 B.n51 VSUBS 0.018241f
C91 B.n52 VSUBS 0.008049f
C92 B.n53 VSUBS 0.008049f
C93 B.n54 VSUBS 0.008049f
C94 B.n55 VSUBS 0.008049f
C95 B.n56 VSUBS 0.008049f
C96 B.n57 VSUBS 0.008049f
C97 B.n58 VSUBS 0.008049f
C98 B.n59 VSUBS 0.008049f
C99 B.n60 VSUBS 0.008049f
C100 B.n61 VSUBS 0.008049f
C101 B.n62 VSUBS 0.008049f
C102 B.n63 VSUBS 0.008049f
C103 B.n64 VSUBS 0.018928f
C104 B.n65 VSUBS 0.008049f
C105 B.n66 VSUBS 0.008049f
C106 B.n67 VSUBS 0.008049f
C107 B.n68 VSUBS 0.008049f
C108 B.n69 VSUBS 0.008049f
C109 B.n70 VSUBS 0.008049f
C110 B.n71 VSUBS 0.008049f
C111 B.n72 VSUBS 0.008049f
C112 B.n73 VSUBS 0.008049f
C113 B.n74 VSUBS 0.008049f
C114 B.n75 VSUBS 0.008049f
C115 B.n76 VSUBS 0.008049f
C116 B.n77 VSUBS 0.008049f
C117 B.n78 VSUBS 0.008049f
C118 B.n79 VSUBS 0.008049f
C119 B.n80 VSUBS 0.008049f
C120 B.t2 VSUBS 0.331022f
C121 B.t1 VSUBS 0.337697f
C122 B.t0 VSUBS 0.169881f
C123 B.n81 VSUBS 0.108151f
C124 B.n82 VSUBS 0.071839f
C125 B.n83 VSUBS 0.008049f
C126 B.n84 VSUBS 0.008049f
C127 B.n85 VSUBS 0.008049f
C128 B.n86 VSUBS 0.008049f
C129 B.n87 VSUBS 0.004735f
C130 B.n88 VSUBS 0.008049f
C131 B.n89 VSUBS 0.008049f
C132 B.n90 VSUBS 0.008049f
C133 B.n91 VSUBS 0.008049f
C134 B.n92 VSUBS 0.008049f
C135 B.n93 VSUBS 0.008049f
C136 B.n94 VSUBS 0.008049f
C137 B.n95 VSUBS 0.008049f
C138 B.n96 VSUBS 0.008049f
C139 B.n97 VSUBS 0.008049f
C140 B.n98 VSUBS 0.008049f
C141 B.n99 VSUBS 0.008049f
C142 B.n100 VSUBS 0.008049f
C143 B.n101 VSUBS 0.008049f
C144 B.n102 VSUBS 0.008049f
C145 B.n103 VSUBS 0.008049f
C146 B.n104 VSUBS 0.018241f
C147 B.n105 VSUBS 0.008049f
C148 B.n106 VSUBS 0.008049f
C149 B.n107 VSUBS 0.008049f
C150 B.n108 VSUBS 0.008049f
C151 B.n109 VSUBS 0.008049f
C152 B.n110 VSUBS 0.008049f
C153 B.n111 VSUBS 0.008049f
C154 B.n112 VSUBS 0.008049f
C155 B.n113 VSUBS 0.008049f
C156 B.n114 VSUBS 0.008049f
C157 B.n115 VSUBS 0.008049f
C158 B.n116 VSUBS 0.008049f
C159 B.n117 VSUBS 0.008049f
C160 B.n118 VSUBS 0.008049f
C161 B.n119 VSUBS 0.008049f
C162 B.n120 VSUBS 0.008049f
C163 B.n121 VSUBS 0.008049f
C164 B.n122 VSUBS 0.008049f
C165 B.n123 VSUBS 0.008049f
C166 B.n124 VSUBS 0.008049f
C167 B.n125 VSUBS 0.018241f
C168 B.n126 VSUBS 0.018928f
C169 B.n127 VSUBS 0.018928f
C170 B.n128 VSUBS 0.008049f
C171 B.n129 VSUBS 0.008049f
C172 B.n130 VSUBS 0.008049f
C173 B.n131 VSUBS 0.008049f
C174 B.n132 VSUBS 0.008049f
C175 B.n133 VSUBS 0.008049f
C176 B.n134 VSUBS 0.008049f
C177 B.n135 VSUBS 0.008049f
C178 B.n136 VSUBS 0.008049f
C179 B.n137 VSUBS 0.008049f
C180 B.n138 VSUBS 0.008049f
C181 B.n139 VSUBS 0.008049f
C182 B.n140 VSUBS 0.008049f
C183 B.n141 VSUBS 0.008049f
C184 B.n142 VSUBS 0.008049f
C185 B.n143 VSUBS 0.008049f
C186 B.n144 VSUBS 0.008049f
C187 B.n145 VSUBS 0.008049f
C188 B.n146 VSUBS 0.008049f
C189 B.n147 VSUBS 0.008049f
C190 B.n148 VSUBS 0.008049f
C191 B.n149 VSUBS 0.008049f
C192 B.n150 VSUBS 0.008049f
C193 B.n151 VSUBS 0.008049f
C194 B.n152 VSUBS 0.008049f
C195 B.n153 VSUBS 0.008049f
C196 B.n154 VSUBS 0.008049f
C197 B.n155 VSUBS 0.008049f
C198 B.n156 VSUBS 0.008049f
C199 B.n157 VSUBS 0.008049f
C200 B.n158 VSUBS 0.008049f
C201 B.n159 VSUBS 0.008049f
C202 B.n160 VSUBS 0.008049f
C203 B.n161 VSUBS 0.008049f
C204 B.n162 VSUBS 0.008049f
C205 B.n163 VSUBS 0.008049f
C206 B.n164 VSUBS 0.008049f
C207 B.n165 VSUBS 0.008049f
C208 B.n166 VSUBS 0.008049f
C209 B.n167 VSUBS 0.008049f
C210 B.n168 VSUBS 0.008049f
C211 B.n169 VSUBS 0.008049f
C212 B.n170 VSUBS 0.008049f
C213 B.n171 VSUBS 0.008049f
C214 B.n172 VSUBS 0.008049f
C215 B.n173 VSUBS 0.008049f
C216 B.t11 VSUBS 0.331025f
C217 B.t10 VSUBS 0.337701f
C218 B.t9 VSUBS 0.169881f
C219 B.n174 VSUBS 0.108148f
C220 B.n175 VSUBS 0.071836f
C221 B.n176 VSUBS 0.018649f
C222 B.n177 VSUBS 0.007339f
C223 B.n178 VSUBS 0.008049f
C224 B.n179 VSUBS 0.008049f
C225 B.n180 VSUBS 0.008049f
C226 B.n181 VSUBS 0.008049f
C227 B.n182 VSUBS 0.008049f
C228 B.n183 VSUBS 0.008049f
C229 B.n184 VSUBS 0.008049f
C230 B.n185 VSUBS 0.008049f
C231 B.n186 VSUBS 0.008049f
C232 B.n187 VSUBS 0.008049f
C233 B.n188 VSUBS 0.008049f
C234 B.n189 VSUBS 0.008049f
C235 B.n190 VSUBS 0.008049f
C236 B.n191 VSUBS 0.008049f
C237 B.n192 VSUBS 0.008049f
C238 B.n193 VSUBS 0.004735f
C239 B.n194 VSUBS 0.018649f
C240 B.n195 VSUBS 0.007339f
C241 B.n196 VSUBS 0.008049f
C242 B.n197 VSUBS 0.008049f
C243 B.n198 VSUBS 0.008049f
C244 B.n199 VSUBS 0.008049f
C245 B.n200 VSUBS 0.008049f
C246 B.n201 VSUBS 0.008049f
C247 B.n202 VSUBS 0.008049f
C248 B.n203 VSUBS 0.008049f
C249 B.n204 VSUBS 0.008049f
C250 B.n205 VSUBS 0.008049f
C251 B.n206 VSUBS 0.008049f
C252 B.n207 VSUBS 0.008049f
C253 B.n208 VSUBS 0.008049f
C254 B.n209 VSUBS 0.008049f
C255 B.n210 VSUBS 0.008049f
C256 B.n211 VSUBS 0.008049f
C257 B.n212 VSUBS 0.008049f
C258 B.n213 VSUBS 0.008049f
C259 B.n214 VSUBS 0.008049f
C260 B.n215 VSUBS 0.008049f
C261 B.n216 VSUBS 0.008049f
C262 B.n217 VSUBS 0.008049f
C263 B.n218 VSUBS 0.008049f
C264 B.n219 VSUBS 0.008049f
C265 B.n220 VSUBS 0.008049f
C266 B.n221 VSUBS 0.008049f
C267 B.n222 VSUBS 0.008049f
C268 B.n223 VSUBS 0.008049f
C269 B.n224 VSUBS 0.008049f
C270 B.n225 VSUBS 0.008049f
C271 B.n226 VSUBS 0.008049f
C272 B.n227 VSUBS 0.008049f
C273 B.n228 VSUBS 0.008049f
C274 B.n229 VSUBS 0.008049f
C275 B.n230 VSUBS 0.008049f
C276 B.n231 VSUBS 0.008049f
C277 B.n232 VSUBS 0.008049f
C278 B.n233 VSUBS 0.008049f
C279 B.n234 VSUBS 0.008049f
C280 B.n235 VSUBS 0.008049f
C281 B.n236 VSUBS 0.008049f
C282 B.n237 VSUBS 0.008049f
C283 B.n238 VSUBS 0.008049f
C284 B.n239 VSUBS 0.008049f
C285 B.n240 VSUBS 0.008049f
C286 B.n241 VSUBS 0.008049f
C287 B.n242 VSUBS 0.008049f
C288 B.n243 VSUBS 0.017957f
C289 B.n244 VSUBS 0.019212f
C290 B.n245 VSUBS 0.018241f
C291 B.n246 VSUBS 0.008049f
C292 B.n247 VSUBS 0.008049f
C293 B.n248 VSUBS 0.008049f
C294 B.n249 VSUBS 0.008049f
C295 B.n250 VSUBS 0.008049f
C296 B.n251 VSUBS 0.008049f
C297 B.n252 VSUBS 0.008049f
C298 B.n253 VSUBS 0.008049f
C299 B.n254 VSUBS 0.008049f
C300 B.n255 VSUBS 0.008049f
C301 B.n256 VSUBS 0.008049f
C302 B.n257 VSUBS 0.008049f
C303 B.n258 VSUBS 0.008049f
C304 B.n259 VSUBS 0.008049f
C305 B.n260 VSUBS 0.008049f
C306 B.n261 VSUBS 0.008049f
C307 B.n262 VSUBS 0.008049f
C308 B.n263 VSUBS 0.008049f
C309 B.n264 VSUBS 0.008049f
C310 B.n265 VSUBS 0.008049f
C311 B.n266 VSUBS 0.008049f
C312 B.n267 VSUBS 0.008049f
C313 B.n268 VSUBS 0.008049f
C314 B.n269 VSUBS 0.008049f
C315 B.n270 VSUBS 0.008049f
C316 B.n271 VSUBS 0.008049f
C317 B.n272 VSUBS 0.008049f
C318 B.n273 VSUBS 0.008049f
C319 B.n274 VSUBS 0.008049f
C320 B.n275 VSUBS 0.008049f
C321 B.n276 VSUBS 0.008049f
C322 B.n277 VSUBS 0.008049f
C323 B.n278 VSUBS 0.008049f
C324 B.n279 VSUBS 0.008049f
C325 B.n280 VSUBS 0.008049f
C326 B.n281 VSUBS 0.008049f
C327 B.n282 VSUBS 0.018241f
C328 B.n283 VSUBS 0.018928f
C329 B.n284 VSUBS 0.018928f
C330 B.n285 VSUBS 0.008049f
C331 B.n286 VSUBS 0.008049f
C332 B.n287 VSUBS 0.008049f
C333 B.n288 VSUBS 0.008049f
C334 B.n289 VSUBS 0.008049f
C335 B.n290 VSUBS 0.008049f
C336 B.n291 VSUBS 0.008049f
C337 B.n292 VSUBS 0.008049f
C338 B.n293 VSUBS 0.008049f
C339 B.n294 VSUBS 0.008049f
C340 B.n295 VSUBS 0.008049f
C341 B.n296 VSUBS 0.008049f
C342 B.n297 VSUBS 0.008049f
C343 B.n298 VSUBS 0.008049f
C344 B.n299 VSUBS 0.008049f
C345 B.n300 VSUBS 0.008049f
C346 B.n301 VSUBS 0.008049f
C347 B.n302 VSUBS 0.008049f
C348 B.n303 VSUBS 0.008049f
C349 B.n304 VSUBS 0.008049f
C350 B.n305 VSUBS 0.008049f
C351 B.n306 VSUBS 0.008049f
C352 B.n307 VSUBS 0.008049f
C353 B.n308 VSUBS 0.008049f
C354 B.n309 VSUBS 0.008049f
C355 B.n310 VSUBS 0.008049f
C356 B.n311 VSUBS 0.008049f
C357 B.n312 VSUBS 0.008049f
C358 B.n313 VSUBS 0.008049f
C359 B.n314 VSUBS 0.008049f
C360 B.n315 VSUBS 0.008049f
C361 B.n316 VSUBS 0.008049f
C362 B.n317 VSUBS 0.008049f
C363 B.n318 VSUBS 0.008049f
C364 B.n319 VSUBS 0.008049f
C365 B.n320 VSUBS 0.008049f
C366 B.n321 VSUBS 0.008049f
C367 B.n322 VSUBS 0.008049f
C368 B.n323 VSUBS 0.008049f
C369 B.n324 VSUBS 0.008049f
C370 B.n325 VSUBS 0.008049f
C371 B.n326 VSUBS 0.008049f
C372 B.n327 VSUBS 0.008049f
C373 B.n328 VSUBS 0.008049f
C374 B.n329 VSUBS 0.008049f
C375 B.n330 VSUBS 0.008049f
C376 B.n331 VSUBS 0.008049f
C377 B.n332 VSUBS 0.007339f
C378 B.n333 VSUBS 0.018649f
C379 B.n334 VSUBS 0.004735f
C380 B.n335 VSUBS 0.008049f
C381 B.n336 VSUBS 0.008049f
C382 B.n337 VSUBS 0.008049f
C383 B.n338 VSUBS 0.008049f
C384 B.n339 VSUBS 0.008049f
C385 B.n340 VSUBS 0.008049f
C386 B.n341 VSUBS 0.008049f
C387 B.n342 VSUBS 0.008049f
C388 B.n343 VSUBS 0.008049f
C389 B.n344 VSUBS 0.008049f
C390 B.n345 VSUBS 0.008049f
C391 B.n346 VSUBS 0.008049f
C392 B.n347 VSUBS 0.004735f
C393 B.n348 VSUBS 0.008049f
C394 B.n349 VSUBS 0.008049f
C395 B.n350 VSUBS 0.008049f
C396 B.n351 VSUBS 0.008049f
C397 B.n352 VSUBS 0.008049f
C398 B.n353 VSUBS 0.008049f
C399 B.n354 VSUBS 0.008049f
C400 B.n355 VSUBS 0.008049f
C401 B.n356 VSUBS 0.008049f
C402 B.n357 VSUBS 0.008049f
C403 B.n358 VSUBS 0.008049f
C404 B.n359 VSUBS 0.008049f
C405 B.n360 VSUBS 0.008049f
C406 B.n361 VSUBS 0.008049f
C407 B.n362 VSUBS 0.008049f
C408 B.n363 VSUBS 0.008049f
C409 B.n364 VSUBS 0.008049f
C410 B.n365 VSUBS 0.008049f
C411 B.n366 VSUBS 0.008049f
C412 B.n367 VSUBS 0.008049f
C413 B.n368 VSUBS 0.008049f
C414 B.n369 VSUBS 0.008049f
C415 B.n370 VSUBS 0.008049f
C416 B.n371 VSUBS 0.008049f
C417 B.n372 VSUBS 0.008049f
C418 B.n373 VSUBS 0.008049f
C419 B.n374 VSUBS 0.008049f
C420 B.n375 VSUBS 0.008049f
C421 B.n376 VSUBS 0.008049f
C422 B.n377 VSUBS 0.008049f
C423 B.n378 VSUBS 0.008049f
C424 B.n379 VSUBS 0.008049f
C425 B.n380 VSUBS 0.008049f
C426 B.n381 VSUBS 0.008049f
C427 B.n382 VSUBS 0.008049f
C428 B.n383 VSUBS 0.008049f
C429 B.n384 VSUBS 0.008049f
C430 B.n385 VSUBS 0.008049f
C431 B.n386 VSUBS 0.008049f
C432 B.n387 VSUBS 0.008049f
C433 B.n388 VSUBS 0.008049f
C434 B.n389 VSUBS 0.008049f
C435 B.n390 VSUBS 0.008049f
C436 B.n391 VSUBS 0.008049f
C437 B.n392 VSUBS 0.008049f
C438 B.n393 VSUBS 0.008049f
C439 B.n394 VSUBS 0.008049f
C440 B.n395 VSUBS 0.008049f
C441 B.n396 VSUBS 0.008049f
C442 B.n397 VSUBS 0.018928f
C443 B.n398 VSUBS 0.018241f
C444 B.n399 VSUBS 0.018241f
C445 B.n400 VSUBS 0.008049f
C446 B.n401 VSUBS 0.008049f
C447 B.n402 VSUBS 0.008049f
C448 B.n403 VSUBS 0.008049f
C449 B.n404 VSUBS 0.008049f
C450 B.n405 VSUBS 0.008049f
C451 B.n406 VSUBS 0.008049f
C452 B.n407 VSUBS 0.008049f
C453 B.n408 VSUBS 0.008049f
C454 B.n409 VSUBS 0.008049f
C455 B.n410 VSUBS 0.008049f
C456 B.n411 VSUBS 0.008049f
C457 B.n412 VSUBS 0.008049f
C458 B.n413 VSUBS 0.008049f
C459 B.n414 VSUBS 0.008049f
C460 B.n415 VSUBS 0.010504f
C461 B.n416 VSUBS 0.011189f
C462 B.n417 VSUBS 0.022251f
C463 VDD1.t0 VSUBS 1.23012f
C464 VDD1.t1 VSUBS 1.57229f
C465 VTAIL.t2 VSUBS 1.78404f
C466 VTAIL.n0 VSUBS 1.96024f
C467 VTAIL.t1 VSUBS 1.78405f
C468 VTAIL.n1 VSUBS 1.96909f
C469 VTAIL.t3 VSUBS 1.78405f
C470 VTAIL.n2 VSUBS 1.91281f
C471 VTAIL.t0 VSUBS 1.78404f
C472 VTAIL.n3 VSUBS 1.85153f
C473 VP.t1 VSUBS 0.526581f
C474 VP.t0 VSUBS 0.463163f
C475 VP.n0 VSUBS 2.90359f
.ends

