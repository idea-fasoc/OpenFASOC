* NGSPICE file created from diff_pair_sample_1010.ext - technology: sky130A

.subckt diff_pair_sample_1010 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=3.2472 ps=20.01 w=19.68 l=2.18
X1 VDD1.t4 VP.t1 VTAIL.t7 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=7.6752 ps=40.14 w=19.68 l=2.18
X2 VTAIL.t8 VP.t2 VDD1.t3 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=3.2472 ps=20.01 w=19.68 l=2.18
X3 VDD2.t5 VN.t0 VTAIL.t2 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=3.2472 ps=20.01 w=19.68 l=2.18
X4 VTAIL.t9 VP.t3 VDD1.t2 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=3.2472 ps=20.01 w=19.68 l=2.18
X5 VTAIL.t3 VN.t1 VDD2.t4 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=3.2472 ps=20.01 w=19.68 l=2.18
X6 VDD2.t3 VN.t2 VTAIL.t5 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=7.6752 ps=40.14 w=19.68 l=2.18
X7 VDD1.t1 VP.t4 VTAIL.t11 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=7.6752 ps=40.14 w=19.68 l=2.18
X8 VDD1.t0 VP.t5 VTAIL.t10 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=3.2472 ps=20.01 w=19.68 l=2.18
X9 VDD2.t2 VN.t3 VTAIL.t4 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=7.6752 ps=40.14 w=19.68 l=2.18
X10 B.t11 B.t9 B.t10 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=0 ps=0 w=19.68 l=2.18
X11 B.t8 B.t6 B.t7 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=0 ps=0 w=19.68 l=2.18
X12 B.t5 B.t3 B.t4 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=0 ps=0 w=19.68 l=2.18
X13 VTAIL.t1 VN.t4 VDD2.t1 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=3.2472 pd=20.01 as=3.2472 ps=20.01 w=19.68 l=2.18
X14 VDD2.t0 VN.t5 VTAIL.t0 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=3.2472 ps=20.01 w=19.68 l=2.18
X15 B.t2 B.t0 B.t1 w_n2978_n4904# sky130_fd_pr__pfet_01v8 ad=7.6752 pd=40.14 as=0 ps=0 w=19.68 l=2.18
R0 VP.n9 VP.t5 249.788
R1 VP.n5 VP.t0 217.564
R2 VP.n29 VP.t3 217.564
R3 VP.n37 VP.t4 217.564
R4 VP.n18 VP.t1 217.564
R5 VP.n10 VP.t2 217.564
R6 VP.n11 VP.n8 161.3
R7 VP.n13 VP.n12 161.3
R8 VP.n14 VP.n7 161.3
R9 VP.n16 VP.n15 161.3
R10 VP.n17 VP.n6 161.3
R11 VP.n36 VP.n0 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n1 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n2 161.3
R16 VP.n28 VP.n27 161.3
R17 VP.n26 VP.n3 161.3
R18 VP.n25 VP.n24 161.3
R19 VP.n23 VP.n4 161.3
R20 VP.n22 VP.n21 161.3
R21 VP.n20 VP.n5 98.1205
R22 VP.n38 VP.n37 98.1205
R23 VP.n19 VP.n18 98.1205
R24 VP.n10 VP.n9 59.417
R25 VP.n20 VP.n19 52.8065
R26 VP.n24 VP.n23 41.0614
R27 VP.n35 VP.n1 41.0614
R28 VP.n16 VP.n7 41.0614
R29 VP.n24 VP.n3 40.0926
R30 VP.n31 VP.n1 40.0926
R31 VP.n12 VP.n7 40.0926
R32 VP.n23 VP.n22 24.5923
R33 VP.n28 VP.n3 24.5923
R34 VP.n31 VP.n30 24.5923
R35 VP.n36 VP.n35 24.5923
R36 VP.n17 VP.n16 24.5923
R37 VP.n12 VP.n11 24.5923
R38 VP.n22 VP.n5 12.7883
R39 VP.n37 VP.n36 12.7883
R40 VP.n18 VP.n17 12.7883
R41 VP.n29 VP.n28 12.2964
R42 VP.n30 VP.n29 12.2964
R43 VP.n11 VP.n10 12.2964
R44 VP.n9 VP.n8 9.65766
R45 VP.n19 VP.n6 0.278335
R46 VP.n21 VP.n20 0.278335
R47 VP.n38 VP.n0 0.278335
R48 VP.n13 VP.n8 0.189894
R49 VP.n14 VP.n13 0.189894
R50 VP.n15 VP.n14 0.189894
R51 VP.n15 VP.n6 0.189894
R52 VP.n21 VP.n4 0.189894
R53 VP.n25 VP.n4 0.189894
R54 VP.n26 VP.n25 0.189894
R55 VP.n27 VP.n26 0.189894
R56 VP.n27 VP.n2 0.189894
R57 VP.n32 VP.n2 0.189894
R58 VP.n33 VP.n32 0.189894
R59 VP.n34 VP.n33 0.189894
R60 VP.n34 VP.n0 0.189894
R61 VP VP.n38 0.153485
R62 VTAIL.n442 VTAIL.n338 756.745
R63 VTAIL.n106 VTAIL.n2 756.745
R64 VTAIL.n332 VTAIL.n228 756.745
R65 VTAIL.n220 VTAIL.n116 756.745
R66 VTAIL.n375 VTAIL.n374 585
R67 VTAIL.n377 VTAIL.n376 585
R68 VTAIL.n370 VTAIL.n369 585
R69 VTAIL.n383 VTAIL.n382 585
R70 VTAIL.n385 VTAIL.n384 585
R71 VTAIL.n366 VTAIL.n365 585
R72 VTAIL.n391 VTAIL.n390 585
R73 VTAIL.n393 VTAIL.n392 585
R74 VTAIL.n362 VTAIL.n361 585
R75 VTAIL.n399 VTAIL.n398 585
R76 VTAIL.n401 VTAIL.n400 585
R77 VTAIL.n358 VTAIL.n357 585
R78 VTAIL.n407 VTAIL.n406 585
R79 VTAIL.n409 VTAIL.n408 585
R80 VTAIL.n354 VTAIL.n353 585
R81 VTAIL.n416 VTAIL.n415 585
R82 VTAIL.n417 VTAIL.n352 585
R83 VTAIL.n419 VTAIL.n418 585
R84 VTAIL.n350 VTAIL.n349 585
R85 VTAIL.n425 VTAIL.n424 585
R86 VTAIL.n427 VTAIL.n426 585
R87 VTAIL.n346 VTAIL.n345 585
R88 VTAIL.n433 VTAIL.n432 585
R89 VTAIL.n435 VTAIL.n434 585
R90 VTAIL.n342 VTAIL.n341 585
R91 VTAIL.n441 VTAIL.n440 585
R92 VTAIL.n443 VTAIL.n442 585
R93 VTAIL.n39 VTAIL.n38 585
R94 VTAIL.n41 VTAIL.n40 585
R95 VTAIL.n34 VTAIL.n33 585
R96 VTAIL.n47 VTAIL.n46 585
R97 VTAIL.n49 VTAIL.n48 585
R98 VTAIL.n30 VTAIL.n29 585
R99 VTAIL.n55 VTAIL.n54 585
R100 VTAIL.n57 VTAIL.n56 585
R101 VTAIL.n26 VTAIL.n25 585
R102 VTAIL.n63 VTAIL.n62 585
R103 VTAIL.n65 VTAIL.n64 585
R104 VTAIL.n22 VTAIL.n21 585
R105 VTAIL.n71 VTAIL.n70 585
R106 VTAIL.n73 VTAIL.n72 585
R107 VTAIL.n18 VTAIL.n17 585
R108 VTAIL.n80 VTAIL.n79 585
R109 VTAIL.n81 VTAIL.n16 585
R110 VTAIL.n83 VTAIL.n82 585
R111 VTAIL.n14 VTAIL.n13 585
R112 VTAIL.n89 VTAIL.n88 585
R113 VTAIL.n91 VTAIL.n90 585
R114 VTAIL.n10 VTAIL.n9 585
R115 VTAIL.n97 VTAIL.n96 585
R116 VTAIL.n99 VTAIL.n98 585
R117 VTAIL.n6 VTAIL.n5 585
R118 VTAIL.n105 VTAIL.n104 585
R119 VTAIL.n107 VTAIL.n106 585
R120 VTAIL.n333 VTAIL.n332 585
R121 VTAIL.n331 VTAIL.n330 585
R122 VTAIL.n232 VTAIL.n231 585
R123 VTAIL.n325 VTAIL.n324 585
R124 VTAIL.n323 VTAIL.n322 585
R125 VTAIL.n236 VTAIL.n235 585
R126 VTAIL.n317 VTAIL.n316 585
R127 VTAIL.n315 VTAIL.n314 585
R128 VTAIL.n240 VTAIL.n239 585
R129 VTAIL.n244 VTAIL.n242 585
R130 VTAIL.n309 VTAIL.n308 585
R131 VTAIL.n307 VTAIL.n306 585
R132 VTAIL.n246 VTAIL.n245 585
R133 VTAIL.n301 VTAIL.n300 585
R134 VTAIL.n299 VTAIL.n298 585
R135 VTAIL.n250 VTAIL.n249 585
R136 VTAIL.n293 VTAIL.n292 585
R137 VTAIL.n291 VTAIL.n290 585
R138 VTAIL.n254 VTAIL.n253 585
R139 VTAIL.n285 VTAIL.n284 585
R140 VTAIL.n283 VTAIL.n282 585
R141 VTAIL.n258 VTAIL.n257 585
R142 VTAIL.n277 VTAIL.n276 585
R143 VTAIL.n275 VTAIL.n274 585
R144 VTAIL.n262 VTAIL.n261 585
R145 VTAIL.n269 VTAIL.n268 585
R146 VTAIL.n267 VTAIL.n266 585
R147 VTAIL.n221 VTAIL.n220 585
R148 VTAIL.n219 VTAIL.n218 585
R149 VTAIL.n120 VTAIL.n119 585
R150 VTAIL.n213 VTAIL.n212 585
R151 VTAIL.n211 VTAIL.n210 585
R152 VTAIL.n124 VTAIL.n123 585
R153 VTAIL.n205 VTAIL.n204 585
R154 VTAIL.n203 VTAIL.n202 585
R155 VTAIL.n128 VTAIL.n127 585
R156 VTAIL.n132 VTAIL.n130 585
R157 VTAIL.n197 VTAIL.n196 585
R158 VTAIL.n195 VTAIL.n194 585
R159 VTAIL.n134 VTAIL.n133 585
R160 VTAIL.n189 VTAIL.n188 585
R161 VTAIL.n187 VTAIL.n186 585
R162 VTAIL.n138 VTAIL.n137 585
R163 VTAIL.n181 VTAIL.n180 585
R164 VTAIL.n179 VTAIL.n178 585
R165 VTAIL.n142 VTAIL.n141 585
R166 VTAIL.n173 VTAIL.n172 585
R167 VTAIL.n171 VTAIL.n170 585
R168 VTAIL.n146 VTAIL.n145 585
R169 VTAIL.n165 VTAIL.n164 585
R170 VTAIL.n163 VTAIL.n162 585
R171 VTAIL.n150 VTAIL.n149 585
R172 VTAIL.n157 VTAIL.n156 585
R173 VTAIL.n155 VTAIL.n154 585
R174 VTAIL.n373 VTAIL.t5 327.466
R175 VTAIL.n37 VTAIL.t11 327.466
R176 VTAIL.n265 VTAIL.t7 327.466
R177 VTAIL.n153 VTAIL.t4 327.466
R178 VTAIL.n376 VTAIL.n375 171.744
R179 VTAIL.n376 VTAIL.n369 171.744
R180 VTAIL.n383 VTAIL.n369 171.744
R181 VTAIL.n384 VTAIL.n383 171.744
R182 VTAIL.n384 VTAIL.n365 171.744
R183 VTAIL.n391 VTAIL.n365 171.744
R184 VTAIL.n392 VTAIL.n391 171.744
R185 VTAIL.n392 VTAIL.n361 171.744
R186 VTAIL.n399 VTAIL.n361 171.744
R187 VTAIL.n400 VTAIL.n399 171.744
R188 VTAIL.n400 VTAIL.n357 171.744
R189 VTAIL.n407 VTAIL.n357 171.744
R190 VTAIL.n408 VTAIL.n407 171.744
R191 VTAIL.n408 VTAIL.n353 171.744
R192 VTAIL.n416 VTAIL.n353 171.744
R193 VTAIL.n417 VTAIL.n416 171.744
R194 VTAIL.n418 VTAIL.n417 171.744
R195 VTAIL.n418 VTAIL.n349 171.744
R196 VTAIL.n425 VTAIL.n349 171.744
R197 VTAIL.n426 VTAIL.n425 171.744
R198 VTAIL.n426 VTAIL.n345 171.744
R199 VTAIL.n433 VTAIL.n345 171.744
R200 VTAIL.n434 VTAIL.n433 171.744
R201 VTAIL.n434 VTAIL.n341 171.744
R202 VTAIL.n441 VTAIL.n341 171.744
R203 VTAIL.n442 VTAIL.n441 171.744
R204 VTAIL.n40 VTAIL.n39 171.744
R205 VTAIL.n40 VTAIL.n33 171.744
R206 VTAIL.n47 VTAIL.n33 171.744
R207 VTAIL.n48 VTAIL.n47 171.744
R208 VTAIL.n48 VTAIL.n29 171.744
R209 VTAIL.n55 VTAIL.n29 171.744
R210 VTAIL.n56 VTAIL.n55 171.744
R211 VTAIL.n56 VTAIL.n25 171.744
R212 VTAIL.n63 VTAIL.n25 171.744
R213 VTAIL.n64 VTAIL.n63 171.744
R214 VTAIL.n64 VTAIL.n21 171.744
R215 VTAIL.n71 VTAIL.n21 171.744
R216 VTAIL.n72 VTAIL.n71 171.744
R217 VTAIL.n72 VTAIL.n17 171.744
R218 VTAIL.n80 VTAIL.n17 171.744
R219 VTAIL.n81 VTAIL.n80 171.744
R220 VTAIL.n82 VTAIL.n81 171.744
R221 VTAIL.n82 VTAIL.n13 171.744
R222 VTAIL.n89 VTAIL.n13 171.744
R223 VTAIL.n90 VTAIL.n89 171.744
R224 VTAIL.n90 VTAIL.n9 171.744
R225 VTAIL.n97 VTAIL.n9 171.744
R226 VTAIL.n98 VTAIL.n97 171.744
R227 VTAIL.n98 VTAIL.n5 171.744
R228 VTAIL.n105 VTAIL.n5 171.744
R229 VTAIL.n106 VTAIL.n105 171.744
R230 VTAIL.n332 VTAIL.n331 171.744
R231 VTAIL.n331 VTAIL.n231 171.744
R232 VTAIL.n324 VTAIL.n231 171.744
R233 VTAIL.n324 VTAIL.n323 171.744
R234 VTAIL.n323 VTAIL.n235 171.744
R235 VTAIL.n316 VTAIL.n235 171.744
R236 VTAIL.n316 VTAIL.n315 171.744
R237 VTAIL.n315 VTAIL.n239 171.744
R238 VTAIL.n244 VTAIL.n239 171.744
R239 VTAIL.n308 VTAIL.n244 171.744
R240 VTAIL.n308 VTAIL.n307 171.744
R241 VTAIL.n307 VTAIL.n245 171.744
R242 VTAIL.n300 VTAIL.n245 171.744
R243 VTAIL.n300 VTAIL.n299 171.744
R244 VTAIL.n299 VTAIL.n249 171.744
R245 VTAIL.n292 VTAIL.n249 171.744
R246 VTAIL.n292 VTAIL.n291 171.744
R247 VTAIL.n291 VTAIL.n253 171.744
R248 VTAIL.n284 VTAIL.n253 171.744
R249 VTAIL.n284 VTAIL.n283 171.744
R250 VTAIL.n283 VTAIL.n257 171.744
R251 VTAIL.n276 VTAIL.n257 171.744
R252 VTAIL.n276 VTAIL.n275 171.744
R253 VTAIL.n275 VTAIL.n261 171.744
R254 VTAIL.n268 VTAIL.n261 171.744
R255 VTAIL.n268 VTAIL.n267 171.744
R256 VTAIL.n220 VTAIL.n219 171.744
R257 VTAIL.n219 VTAIL.n119 171.744
R258 VTAIL.n212 VTAIL.n119 171.744
R259 VTAIL.n212 VTAIL.n211 171.744
R260 VTAIL.n211 VTAIL.n123 171.744
R261 VTAIL.n204 VTAIL.n123 171.744
R262 VTAIL.n204 VTAIL.n203 171.744
R263 VTAIL.n203 VTAIL.n127 171.744
R264 VTAIL.n132 VTAIL.n127 171.744
R265 VTAIL.n196 VTAIL.n132 171.744
R266 VTAIL.n196 VTAIL.n195 171.744
R267 VTAIL.n195 VTAIL.n133 171.744
R268 VTAIL.n188 VTAIL.n133 171.744
R269 VTAIL.n188 VTAIL.n187 171.744
R270 VTAIL.n187 VTAIL.n137 171.744
R271 VTAIL.n180 VTAIL.n137 171.744
R272 VTAIL.n180 VTAIL.n179 171.744
R273 VTAIL.n179 VTAIL.n141 171.744
R274 VTAIL.n172 VTAIL.n141 171.744
R275 VTAIL.n172 VTAIL.n171 171.744
R276 VTAIL.n171 VTAIL.n145 171.744
R277 VTAIL.n164 VTAIL.n145 171.744
R278 VTAIL.n164 VTAIL.n163 171.744
R279 VTAIL.n163 VTAIL.n149 171.744
R280 VTAIL.n156 VTAIL.n149 171.744
R281 VTAIL.n156 VTAIL.n155 171.744
R282 VTAIL.n375 VTAIL.t5 85.8723
R283 VTAIL.n39 VTAIL.t11 85.8723
R284 VTAIL.n267 VTAIL.t7 85.8723
R285 VTAIL.n155 VTAIL.t4 85.8723
R286 VTAIL.n227 VTAIL.n226 51.431
R287 VTAIL.n115 VTAIL.n114 51.431
R288 VTAIL.n1 VTAIL.n0 51.4308
R289 VTAIL.n113 VTAIL.n112 51.4308
R290 VTAIL.n115 VTAIL.n113 33.66
R291 VTAIL.n447 VTAIL.n446 32.1853
R292 VTAIL.n111 VTAIL.n110 32.1853
R293 VTAIL.n337 VTAIL.n336 32.1853
R294 VTAIL.n225 VTAIL.n224 32.1853
R295 VTAIL.n447 VTAIL.n337 31.4962
R296 VTAIL.n374 VTAIL.n373 16.3895
R297 VTAIL.n38 VTAIL.n37 16.3895
R298 VTAIL.n266 VTAIL.n265 16.3895
R299 VTAIL.n154 VTAIL.n153 16.3895
R300 VTAIL.n419 VTAIL.n350 13.1884
R301 VTAIL.n83 VTAIL.n14 13.1884
R302 VTAIL.n242 VTAIL.n240 13.1884
R303 VTAIL.n130 VTAIL.n128 13.1884
R304 VTAIL.n377 VTAIL.n372 12.8005
R305 VTAIL.n420 VTAIL.n352 12.8005
R306 VTAIL.n424 VTAIL.n423 12.8005
R307 VTAIL.n41 VTAIL.n36 12.8005
R308 VTAIL.n84 VTAIL.n16 12.8005
R309 VTAIL.n88 VTAIL.n87 12.8005
R310 VTAIL.n314 VTAIL.n313 12.8005
R311 VTAIL.n310 VTAIL.n309 12.8005
R312 VTAIL.n269 VTAIL.n264 12.8005
R313 VTAIL.n202 VTAIL.n201 12.8005
R314 VTAIL.n198 VTAIL.n197 12.8005
R315 VTAIL.n157 VTAIL.n152 12.8005
R316 VTAIL.n378 VTAIL.n370 12.0247
R317 VTAIL.n415 VTAIL.n414 12.0247
R318 VTAIL.n427 VTAIL.n348 12.0247
R319 VTAIL.n42 VTAIL.n34 12.0247
R320 VTAIL.n79 VTAIL.n78 12.0247
R321 VTAIL.n91 VTAIL.n12 12.0247
R322 VTAIL.n317 VTAIL.n238 12.0247
R323 VTAIL.n306 VTAIL.n243 12.0247
R324 VTAIL.n270 VTAIL.n262 12.0247
R325 VTAIL.n205 VTAIL.n126 12.0247
R326 VTAIL.n194 VTAIL.n131 12.0247
R327 VTAIL.n158 VTAIL.n150 12.0247
R328 VTAIL.n382 VTAIL.n381 11.249
R329 VTAIL.n413 VTAIL.n354 11.249
R330 VTAIL.n428 VTAIL.n346 11.249
R331 VTAIL.n46 VTAIL.n45 11.249
R332 VTAIL.n77 VTAIL.n18 11.249
R333 VTAIL.n92 VTAIL.n10 11.249
R334 VTAIL.n318 VTAIL.n236 11.249
R335 VTAIL.n305 VTAIL.n246 11.249
R336 VTAIL.n274 VTAIL.n273 11.249
R337 VTAIL.n206 VTAIL.n124 11.249
R338 VTAIL.n193 VTAIL.n134 11.249
R339 VTAIL.n162 VTAIL.n161 11.249
R340 VTAIL.n385 VTAIL.n368 10.4732
R341 VTAIL.n410 VTAIL.n409 10.4732
R342 VTAIL.n432 VTAIL.n431 10.4732
R343 VTAIL.n49 VTAIL.n32 10.4732
R344 VTAIL.n74 VTAIL.n73 10.4732
R345 VTAIL.n96 VTAIL.n95 10.4732
R346 VTAIL.n322 VTAIL.n321 10.4732
R347 VTAIL.n302 VTAIL.n301 10.4732
R348 VTAIL.n277 VTAIL.n260 10.4732
R349 VTAIL.n210 VTAIL.n209 10.4732
R350 VTAIL.n190 VTAIL.n189 10.4732
R351 VTAIL.n165 VTAIL.n148 10.4732
R352 VTAIL.n386 VTAIL.n366 9.69747
R353 VTAIL.n406 VTAIL.n356 9.69747
R354 VTAIL.n435 VTAIL.n344 9.69747
R355 VTAIL.n50 VTAIL.n30 9.69747
R356 VTAIL.n70 VTAIL.n20 9.69747
R357 VTAIL.n99 VTAIL.n8 9.69747
R358 VTAIL.n325 VTAIL.n234 9.69747
R359 VTAIL.n298 VTAIL.n248 9.69747
R360 VTAIL.n278 VTAIL.n258 9.69747
R361 VTAIL.n213 VTAIL.n122 9.69747
R362 VTAIL.n186 VTAIL.n136 9.69747
R363 VTAIL.n166 VTAIL.n146 9.69747
R364 VTAIL.n446 VTAIL.n445 9.45567
R365 VTAIL.n110 VTAIL.n109 9.45567
R366 VTAIL.n336 VTAIL.n335 9.45567
R367 VTAIL.n224 VTAIL.n223 9.45567
R368 VTAIL.n445 VTAIL.n444 9.3005
R369 VTAIL.n439 VTAIL.n438 9.3005
R370 VTAIL.n437 VTAIL.n436 9.3005
R371 VTAIL.n344 VTAIL.n343 9.3005
R372 VTAIL.n431 VTAIL.n430 9.3005
R373 VTAIL.n429 VTAIL.n428 9.3005
R374 VTAIL.n348 VTAIL.n347 9.3005
R375 VTAIL.n423 VTAIL.n422 9.3005
R376 VTAIL.n395 VTAIL.n394 9.3005
R377 VTAIL.n364 VTAIL.n363 9.3005
R378 VTAIL.n389 VTAIL.n388 9.3005
R379 VTAIL.n387 VTAIL.n386 9.3005
R380 VTAIL.n368 VTAIL.n367 9.3005
R381 VTAIL.n381 VTAIL.n380 9.3005
R382 VTAIL.n379 VTAIL.n378 9.3005
R383 VTAIL.n372 VTAIL.n371 9.3005
R384 VTAIL.n397 VTAIL.n396 9.3005
R385 VTAIL.n360 VTAIL.n359 9.3005
R386 VTAIL.n403 VTAIL.n402 9.3005
R387 VTAIL.n405 VTAIL.n404 9.3005
R388 VTAIL.n356 VTAIL.n355 9.3005
R389 VTAIL.n411 VTAIL.n410 9.3005
R390 VTAIL.n413 VTAIL.n412 9.3005
R391 VTAIL.n414 VTAIL.n351 9.3005
R392 VTAIL.n421 VTAIL.n420 9.3005
R393 VTAIL.n340 VTAIL.n339 9.3005
R394 VTAIL.n109 VTAIL.n108 9.3005
R395 VTAIL.n103 VTAIL.n102 9.3005
R396 VTAIL.n101 VTAIL.n100 9.3005
R397 VTAIL.n8 VTAIL.n7 9.3005
R398 VTAIL.n95 VTAIL.n94 9.3005
R399 VTAIL.n93 VTAIL.n92 9.3005
R400 VTAIL.n12 VTAIL.n11 9.3005
R401 VTAIL.n87 VTAIL.n86 9.3005
R402 VTAIL.n59 VTAIL.n58 9.3005
R403 VTAIL.n28 VTAIL.n27 9.3005
R404 VTAIL.n53 VTAIL.n52 9.3005
R405 VTAIL.n51 VTAIL.n50 9.3005
R406 VTAIL.n32 VTAIL.n31 9.3005
R407 VTAIL.n45 VTAIL.n44 9.3005
R408 VTAIL.n43 VTAIL.n42 9.3005
R409 VTAIL.n36 VTAIL.n35 9.3005
R410 VTAIL.n61 VTAIL.n60 9.3005
R411 VTAIL.n24 VTAIL.n23 9.3005
R412 VTAIL.n67 VTAIL.n66 9.3005
R413 VTAIL.n69 VTAIL.n68 9.3005
R414 VTAIL.n20 VTAIL.n19 9.3005
R415 VTAIL.n75 VTAIL.n74 9.3005
R416 VTAIL.n77 VTAIL.n76 9.3005
R417 VTAIL.n78 VTAIL.n15 9.3005
R418 VTAIL.n85 VTAIL.n84 9.3005
R419 VTAIL.n4 VTAIL.n3 9.3005
R420 VTAIL.n252 VTAIL.n251 9.3005
R421 VTAIL.n295 VTAIL.n294 9.3005
R422 VTAIL.n297 VTAIL.n296 9.3005
R423 VTAIL.n248 VTAIL.n247 9.3005
R424 VTAIL.n303 VTAIL.n302 9.3005
R425 VTAIL.n305 VTAIL.n304 9.3005
R426 VTAIL.n243 VTAIL.n241 9.3005
R427 VTAIL.n311 VTAIL.n310 9.3005
R428 VTAIL.n335 VTAIL.n334 9.3005
R429 VTAIL.n230 VTAIL.n229 9.3005
R430 VTAIL.n329 VTAIL.n328 9.3005
R431 VTAIL.n327 VTAIL.n326 9.3005
R432 VTAIL.n234 VTAIL.n233 9.3005
R433 VTAIL.n321 VTAIL.n320 9.3005
R434 VTAIL.n319 VTAIL.n318 9.3005
R435 VTAIL.n238 VTAIL.n237 9.3005
R436 VTAIL.n313 VTAIL.n312 9.3005
R437 VTAIL.n289 VTAIL.n288 9.3005
R438 VTAIL.n287 VTAIL.n286 9.3005
R439 VTAIL.n256 VTAIL.n255 9.3005
R440 VTAIL.n281 VTAIL.n280 9.3005
R441 VTAIL.n279 VTAIL.n278 9.3005
R442 VTAIL.n260 VTAIL.n259 9.3005
R443 VTAIL.n273 VTAIL.n272 9.3005
R444 VTAIL.n271 VTAIL.n270 9.3005
R445 VTAIL.n264 VTAIL.n263 9.3005
R446 VTAIL.n140 VTAIL.n139 9.3005
R447 VTAIL.n183 VTAIL.n182 9.3005
R448 VTAIL.n185 VTAIL.n184 9.3005
R449 VTAIL.n136 VTAIL.n135 9.3005
R450 VTAIL.n191 VTAIL.n190 9.3005
R451 VTAIL.n193 VTAIL.n192 9.3005
R452 VTAIL.n131 VTAIL.n129 9.3005
R453 VTAIL.n199 VTAIL.n198 9.3005
R454 VTAIL.n223 VTAIL.n222 9.3005
R455 VTAIL.n118 VTAIL.n117 9.3005
R456 VTAIL.n217 VTAIL.n216 9.3005
R457 VTAIL.n215 VTAIL.n214 9.3005
R458 VTAIL.n122 VTAIL.n121 9.3005
R459 VTAIL.n209 VTAIL.n208 9.3005
R460 VTAIL.n207 VTAIL.n206 9.3005
R461 VTAIL.n126 VTAIL.n125 9.3005
R462 VTAIL.n201 VTAIL.n200 9.3005
R463 VTAIL.n177 VTAIL.n176 9.3005
R464 VTAIL.n175 VTAIL.n174 9.3005
R465 VTAIL.n144 VTAIL.n143 9.3005
R466 VTAIL.n169 VTAIL.n168 9.3005
R467 VTAIL.n167 VTAIL.n166 9.3005
R468 VTAIL.n148 VTAIL.n147 9.3005
R469 VTAIL.n161 VTAIL.n160 9.3005
R470 VTAIL.n159 VTAIL.n158 9.3005
R471 VTAIL.n152 VTAIL.n151 9.3005
R472 VTAIL.n390 VTAIL.n389 8.92171
R473 VTAIL.n405 VTAIL.n358 8.92171
R474 VTAIL.n436 VTAIL.n342 8.92171
R475 VTAIL.n54 VTAIL.n53 8.92171
R476 VTAIL.n69 VTAIL.n22 8.92171
R477 VTAIL.n100 VTAIL.n6 8.92171
R478 VTAIL.n326 VTAIL.n232 8.92171
R479 VTAIL.n297 VTAIL.n250 8.92171
R480 VTAIL.n282 VTAIL.n281 8.92171
R481 VTAIL.n214 VTAIL.n120 8.92171
R482 VTAIL.n185 VTAIL.n138 8.92171
R483 VTAIL.n170 VTAIL.n169 8.92171
R484 VTAIL.n393 VTAIL.n364 8.14595
R485 VTAIL.n402 VTAIL.n401 8.14595
R486 VTAIL.n440 VTAIL.n439 8.14595
R487 VTAIL.n57 VTAIL.n28 8.14595
R488 VTAIL.n66 VTAIL.n65 8.14595
R489 VTAIL.n104 VTAIL.n103 8.14595
R490 VTAIL.n330 VTAIL.n329 8.14595
R491 VTAIL.n294 VTAIL.n293 8.14595
R492 VTAIL.n285 VTAIL.n256 8.14595
R493 VTAIL.n218 VTAIL.n217 8.14595
R494 VTAIL.n182 VTAIL.n181 8.14595
R495 VTAIL.n173 VTAIL.n144 8.14595
R496 VTAIL.n394 VTAIL.n362 7.3702
R497 VTAIL.n398 VTAIL.n360 7.3702
R498 VTAIL.n443 VTAIL.n340 7.3702
R499 VTAIL.n446 VTAIL.n338 7.3702
R500 VTAIL.n58 VTAIL.n26 7.3702
R501 VTAIL.n62 VTAIL.n24 7.3702
R502 VTAIL.n107 VTAIL.n4 7.3702
R503 VTAIL.n110 VTAIL.n2 7.3702
R504 VTAIL.n336 VTAIL.n228 7.3702
R505 VTAIL.n333 VTAIL.n230 7.3702
R506 VTAIL.n290 VTAIL.n252 7.3702
R507 VTAIL.n286 VTAIL.n254 7.3702
R508 VTAIL.n224 VTAIL.n116 7.3702
R509 VTAIL.n221 VTAIL.n118 7.3702
R510 VTAIL.n178 VTAIL.n140 7.3702
R511 VTAIL.n174 VTAIL.n142 7.3702
R512 VTAIL.n397 VTAIL.n362 6.59444
R513 VTAIL.n398 VTAIL.n397 6.59444
R514 VTAIL.n444 VTAIL.n443 6.59444
R515 VTAIL.n444 VTAIL.n338 6.59444
R516 VTAIL.n61 VTAIL.n26 6.59444
R517 VTAIL.n62 VTAIL.n61 6.59444
R518 VTAIL.n108 VTAIL.n107 6.59444
R519 VTAIL.n108 VTAIL.n2 6.59444
R520 VTAIL.n334 VTAIL.n228 6.59444
R521 VTAIL.n334 VTAIL.n333 6.59444
R522 VTAIL.n290 VTAIL.n289 6.59444
R523 VTAIL.n289 VTAIL.n254 6.59444
R524 VTAIL.n222 VTAIL.n116 6.59444
R525 VTAIL.n222 VTAIL.n221 6.59444
R526 VTAIL.n178 VTAIL.n177 6.59444
R527 VTAIL.n177 VTAIL.n142 6.59444
R528 VTAIL.n394 VTAIL.n393 5.81868
R529 VTAIL.n401 VTAIL.n360 5.81868
R530 VTAIL.n440 VTAIL.n340 5.81868
R531 VTAIL.n58 VTAIL.n57 5.81868
R532 VTAIL.n65 VTAIL.n24 5.81868
R533 VTAIL.n104 VTAIL.n4 5.81868
R534 VTAIL.n330 VTAIL.n230 5.81868
R535 VTAIL.n293 VTAIL.n252 5.81868
R536 VTAIL.n286 VTAIL.n285 5.81868
R537 VTAIL.n218 VTAIL.n118 5.81868
R538 VTAIL.n181 VTAIL.n140 5.81868
R539 VTAIL.n174 VTAIL.n173 5.81868
R540 VTAIL.n390 VTAIL.n364 5.04292
R541 VTAIL.n402 VTAIL.n358 5.04292
R542 VTAIL.n439 VTAIL.n342 5.04292
R543 VTAIL.n54 VTAIL.n28 5.04292
R544 VTAIL.n66 VTAIL.n22 5.04292
R545 VTAIL.n103 VTAIL.n6 5.04292
R546 VTAIL.n329 VTAIL.n232 5.04292
R547 VTAIL.n294 VTAIL.n250 5.04292
R548 VTAIL.n282 VTAIL.n256 5.04292
R549 VTAIL.n217 VTAIL.n120 5.04292
R550 VTAIL.n182 VTAIL.n138 5.04292
R551 VTAIL.n170 VTAIL.n144 5.04292
R552 VTAIL.n389 VTAIL.n366 4.26717
R553 VTAIL.n406 VTAIL.n405 4.26717
R554 VTAIL.n436 VTAIL.n435 4.26717
R555 VTAIL.n53 VTAIL.n30 4.26717
R556 VTAIL.n70 VTAIL.n69 4.26717
R557 VTAIL.n100 VTAIL.n99 4.26717
R558 VTAIL.n326 VTAIL.n325 4.26717
R559 VTAIL.n298 VTAIL.n297 4.26717
R560 VTAIL.n281 VTAIL.n258 4.26717
R561 VTAIL.n214 VTAIL.n213 4.26717
R562 VTAIL.n186 VTAIL.n185 4.26717
R563 VTAIL.n169 VTAIL.n146 4.26717
R564 VTAIL.n373 VTAIL.n371 3.70982
R565 VTAIL.n37 VTAIL.n35 3.70982
R566 VTAIL.n265 VTAIL.n263 3.70982
R567 VTAIL.n153 VTAIL.n151 3.70982
R568 VTAIL.n386 VTAIL.n385 3.49141
R569 VTAIL.n409 VTAIL.n356 3.49141
R570 VTAIL.n432 VTAIL.n344 3.49141
R571 VTAIL.n50 VTAIL.n49 3.49141
R572 VTAIL.n73 VTAIL.n20 3.49141
R573 VTAIL.n96 VTAIL.n8 3.49141
R574 VTAIL.n322 VTAIL.n234 3.49141
R575 VTAIL.n301 VTAIL.n248 3.49141
R576 VTAIL.n278 VTAIL.n277 3.49141
R577 VTAIL.n210 VTAIL.n122 3.49141
R578 VTAIL.n189 VTAIL.n136 3.49141
R579 VTAIL.n166 VTAIL.n165 3.49141
R580 VTAIL.n382 VTAIL.n368 2.71565
R581 VTAIL.n410 VTAIL.n354 2.71565
R582 VTAIL.n431 VTAIL.n346 2.71565
R583 VTAIL.n46 VTAIL.n32 2.71565
R584 VTAIL.n74 VTAIL.n18 2.71565
R585 VTAIL.n95 VTAIL.n10 2.71565
R586 VTAIL.n321 VTAIL.n236 2.71565
R587 VTAIL.n302 VTAIL.n246 2.71565
R588 VTAIL.n274 VTAIL.n260 2.71565
R589 VTAIL.n209 VTAIL.n124 2.71565
R590 VTAIL.n190 VTAIL.n134 2.71565
R591 VTAIL.n162 VTAIL.n148 2.71565
R592 VTAIL.n225 VTAIL.n115 2.16429
R593 VTAIL.n337 VTAIL.n227 2.16429
R594 VTAIL.n113 VTAIL.n111 2.16429
R595 VTAIL.n381 VTAIL.n370 1.93989
R596 VTAIL.n415 VTAIL.n413 1.93989
R597 VTAIL.n428 VTAIL.n427 1.93989
R598 VTAIL.n45 VTAIL.n34 1.93989
R599 VTAIL.n79 VTAIL.n77 1.93989
R600 VTAIL.n92 VTAIL.n91 1.93989
R601 VTAIL.n318 VTAIL.n317 1.93989
R602 VTAIL.n306 VTAIL.n305 1.93989
R603 VTAIL.n273 VTAIL.n262 1.93989
R604 VTAIL.n206 VTAIL.n205 1.93989
R605 VTAIL.n194 VTAIL.n193 1.93989
R606 VTAIL.n161 VTAIL.n150 1.93989
R607 VTAIL.n0 VTAIL.t0 1.65218
R608 VTAIL.n0 VTAIL.t1 1.65218
R609 VTAIL.n112 VTAIL.t6 1.65218
R610 VTAIL.n112 VTAIL.t9 1.65218
R611 VTAIL.n226 VTAIL.t10 1.65218
R612 VTAIL.n226 VTAIL.t8 1.65218
R613 VTAIL.n114 VTAIL.t2 1.65218
R614 VTAIL.n114 VTAIL.t3 1.65218
R615 VTAIL VTAIL.n447 1.56516
R616 VTAIL.n227 VTAIL.n225 1.55222
R617 VTAIL.n111 VTAIL.n1 1.55222
R618 VTAIL.n378 VTAIL.n377 1.16414
R619 VTAIL.n414 VTAIL.n352 1.16414
R620 VTAIL.n424 VTAIL.n348 1.16414
R621 VTAIL.n42 VTAIL.n41 1.16414
R622 VTAIL.n78 VTAIL.n16 1.16414
R623 VTAIL.n88 VTAIL.n12 1.16414
R624 VTAIL.n314 VTAIL.n238 1.16414
R625 VTAIL.n309 VTAIL.n243 1.16414
R626 VTAIL.n270 VTAIL.n269 1.16414
R627 VTAIL.n202 VTAIL.n126 1.16414
R628 VTAIL.n197 VTAIL.n131 1.16414
R629 VTAIL.n158 VTAIL.n157 1.16414
R630 VTAIL VTAIL.n1 0.599638
R631 VTAIL.n374 VTAIL.n372 0.388379
R632 VTAIL.n420 VTAIL.n419 0.388379
R633 VTAIL.n423 VTAIL.n350 0.388379
R634 VTAIL.n38 VTAIL.n36 0.388379
R635 VTAIL.n84 VTAIL.n83 0.388379
R636 VTAIL.n87 VTAIL.n14 0.388379
R637 VTAIL.n313 VTAIL.n240 0.388379
R638 VTAIL.n310 VTAIL.n242 0.388379
R639 VTAIL.n266 VTAIL.n264 0.388379
R640 VTAIL.n201 VTAIL.n128 0.388379
R641 VTAIL.n198 VTAIL.n130 0.388379
R642 VTAIL.n154 VTAIL.n152 0.388379
R643 VTAIL.n379 VTAIL.n371 0.155672
R644 VTAIL.n380 VTAIL.n379 0.155672
R645 VTAIL.n380 VTAIL.n367 0.155672
R646 VTAIL.n387 VTAIL.n367 0.155672
R647 VTAIL.n388 VTAIL.n387 0.155672
R648 VTAIL.n388 VTAIL.n363 0.155672
R649 VTAIL.n395 VTAIL.n363 0.155672
R650 VTAIL.n396 VTAIL.n395 0.155672
R651 VTAIL.n396 VTAIL.n359 0.155672
R652 VTAIL.n403 VTAIL.n359 0.155672
R653 VTAIL.n404 VTAIL.n403 0.155672
R654 VTAIL.n404 VTAIL.n355 0.155672
R655 VTAIL.n411 VTAIL.n355 0.155672
R656 VTAIL.n412 VTAIL.n411 0.155672
R657 VTAIL.n412 VTAIL.n351 0.155672
R658 VTAIL.n421 VTAIL.n351 0.155672
R659 VTAIL.n422 VTAIL.n421 0.155672
R660 VTAIL.n422 VTAIL.n347 0.155672
R661 VTAIL.n429 VTAIL.n347 0.155672
R662 VTAIL.n430 VTAIL.n429 0.155672
R663 VTAIL.n430 VTAIL.n343 0.155672
R664 VTAIL.n437 VTAIL.n343 0.155672
R665 VTAIL.n438 VTAIL.n437 0.155672
R666 VTAIL.n438 VTAIL.n339 0.155672
R667 VTAIL.n445 VTAIL.n339 0.155672
R668 VTAIL.n43 VTAIL.n35 0.155672
R669 VTAIL.n44 VTAIL.n43 0.155672
R670 VTAIL.n44 VTAIL.n31 0.155672
R671 VTAIL.n51 VTAIL.n31 0.155672
R672 VTAIL.n52 VTAIL.n51 0.155672
R673 VTAIL.n52 VTAIL.n27 0.155672
R674 VTAIL.n59 VTAIL.n27 0.155672
R675 VTAIL.n60 VTAIL.n59 0.155672
R676 VTAIL.n60 VTAIL.n23 0.155672
R677 VTAIL.n67 VTAIL.n23 0.155672
R678 VTAIL.n68 VTAIL.n67 0.155672
R679 VTAIL.n68 VTAIL.n19 0.155672
R680 VTAIL.n75 VTAIL.n19 0.155672
R681 VTAIL.n76 VTAIL.n75 0.155672
R682 VTAIL.n76 VTAIL.n15 0.155672
R683 VTAIL.n85 VTAIL.n15 0.155672
R684 VTAIL.n86 VTAIL.n85 0.155672
R685 VTAIL.n86 VTAIL.n11 0.155672
R686 VTAIL.n93 VTAIL.n11 0.155672
R687 VTAIL.n94 VTAIL.n93 0.155672
R688 VTAIL.n94 VTAIL.n7 0.155672
R689 VTAIL.n101 VTAIL.n7 0.155672
R690 VTAIL.n102 VTAIL.n101 0.155672
R691 VTAIL.n102 VTAIL.n3 0.155672
R692 VTAIL.n109 VTAIL.n3 0.155672
R693 VTAIL.n335 VTAIL.n229 0.155672
R694 VTAIL.n328 VTAIL.n229 0.155672
R695 VTAIL.n328 VTAIL.n327 0.155672
R696 VTAIL.n327 VTAIL.n233 0.155672
R697 VTAIL.n320 VTAIL.n233 0.155672
R698 VTAIL.n320 VTAIL.n319 0.155672
R699 VTAIL.n319 VTAIL.n237 0.155672
R700 VTAIL.n312 VTAIL.n237 0.155672
R701 VTAIL.n312 VTAIL.n311 0.155672
R702 VTAIL.n311 VTAIL.n241 0.155672
R703 VTAIL.n304 VTAIL.n241 0.155672
R704 VTAIL.n304 VTAIL.n303 0.155672
R705 VTAIL.n303 VTAIL.n247 0.155672
R706 VTAIL.n296 VTAIL.n247 0.155672
R707 VTAIL.n296 VTAIL.n295 0.155672
R708 VTAIL.n295 VTAIL.n251 0.155672
R709 VTAIL.n288 VTAIL.n251 0.155672
R710 VTAIL.n288 VTAIL.n287 0.155672
R711 VTAIL.n287 VTAIL.n255 0.155672
R712 VTAIL.n280 VTAIL.n255 0.155672
R713 VTAIL.n280 VTAIL.n279 0.155672
R714 VTAIL.n279 VTAIL.n259 0.155672
R715 VTAIL.n272 VTAIL.n259 0.155672
R716 VTAIL.n272 VTAIL.n271 0.155672
R717 VTAIL.n271 VTAIL.n263 0.155672
R718 VTAIL.n223 VTAIL.n117 0.155672
R719 VTAIL.n216 VTAIL.n117 0.155672
R720 VTAIL.n216 VTAIL.n215 0.155672
R721 VTAIL.n215 VTAIL.n121 0.155672
R722 VTAIL.n208 VTAIL.n121 0.155672
R723 VTAIL.n208 VTAIL.n207 0.155672
R724 VTAIL.n207 VTAIL.n125 0.155672
R725 VTAIL.n200 VTAIL.n125 0.155672
R726 VTAIL.n200 VTAIL.n199 0.155672
R727 VTAIL.n199 VTAIL.n129 0.155672
R728 VTAIL.n192 VTAIL.n129 0.155672
R729 VTAIL.n192 VTAIL.n191 0.155672
R730 VTAIL.n191 VTAIL.n135 0.155672
R731 VTAIL.n184 VTAIL.n135 0.155672
R732 VTAIL.n184 VTAIL.n183 0.155672
R733 VTAIL.n183 VTAIL.n139 0.155672
R734 VTAIL.n176 VTAIL.n139 0.155672
R735 VTAIL.n176 VTAIL.n175 0.155672
R736 VTAIL.n175 VTAIL.n143 0.155672
R737 VTAIL.n168 VTAIL.n143 0.155672
R738 VTAIL.n168 VTAIL.n167 0.155672
R739 VTAIL.n167 VTAIL.n147 0.155672
R740 VTAIL.n160 VTAIL.n147 0.155672
R741 VTAIL.n160 VTAIL.n159 0.155672
R742 VTAIL.n159 VTAIL.n151 0.155672
R743 VDD1.n104 VDD1.n0 756.745
R744 VDD1.n213 VDD1.n109 756.745
R745 VDD1.n105 VDD1.n104 585
R746 VDD1.n103 VDD1.n102 585
R747 VDD1.n4 VDD1.n3 585
R748 VDD1.n97 VDD1.n96 585
R749 VDD1.n95 VDD1.n94 585
R750 VDD1.n8 VDD1.n7 585
R751 VDD1.n89 VDD1.n88 585
R752 VDD1.n87 VDD1.n86 585
R753 VDD1.n12 VDD1.n11 585
R754 VDD1.n16 VDD1.n14 585
R755 VDD1.n81 VDD1.n80 585
R756 VDD1.n79 VDD1.n78 585
R757 VDD1.n18 VDD1.n17 585
R758 VDD1.n73 VDD1.n72 585
R759 VDD1.n71 VDD1.n70 585
R760 VDD1.n22 VDD1.n21 585
R761 VDD1.n65 VDD1.n64 585
R762 VDD1.n63 VDD1.n62 585
R763 VDD1.n26 VDD1.n25 585
R764 VDD1.n57 VDD1.n56 585
R765 VDD1.n55 VDD1.n54 585
R766 VDD1.n30 VDD1.n29 585
R767 VDD1.n49 VDD1.n48 585
R768 VDD1.n47 VDD1.n46 585
R769 VDD1.n34 VDD1.n33 585
R770 VDD1.n41 VDD1.n40 585
R771 VDD1.n39 VDD1.n38 585
R772 VDD1.n146 VDD1.n145 585
R773 VDD1.n148 VDD1.n147 585
R774 VDD1.n141 VDD1.n140 585
R775 VDD1.n154 VDD1.n153 585
R776 VDD1.n156 VDD1.n155 585
R777 VDD1.n137 VDD1.n136 585
R778 VDD1.n162 VDD1.n161 585
R779 VDD1.n164 VDD1.n163 585
R780 VDD1.n133 VDD1.n132 585
R781 VDD1.n170 VDD1.n169 585
R782 VDD1.n172 VDD1.n171 585
R783 VDD1.n129 VDD1.n128 585
R784 VDD1.n178 VDD1.n177 585
R785 VDD1.n180 VDD1.n179 585
R786 VDD1.n125 VDD1.n124 585
R787 VDD1.n187 VDD1.n186 585
R788 VDD1.n188 VDD1.n123 585
R789 VDD1.n190 VDD1.n189 585
R790 VDD1.n121 VDD1.n120 585
R791 VDD1.n196 VDD1.n195 585
R792 VDD1.n198 VDD1.n197 585
R793 VDD1.n117 VDD1.n116 585
R794 VDD1.n204 VDD1.n203 585
R795 VDD1.n206 VDD1.n205 585
R796 VDD1.n113 VDD1.n112 585
R797 VDD1.n212 VDD1.n211 585
R798 VDD1.n214 VDD1.n213 585
R799 VDD1.n37 VDD1.t0 327.466
R800 VDD1.n144 VDD1.t5 327.466
R801 VDD1.n104 VDD1.n103 171.744
R802 VDD1.n103 VDD1.n3 171.744
R803 VDD1.n96 VDD1.n3 171.744
R804 VDD1.n96 VDD1.n95 171.744
R805 VDD1.n95 VDD1.n7 171.744
R806 VDD1.n88 VDD1.n7 171.744
R807 VDD1.n88 VDD1.n87 171.744
R808 VDD1.n87 VDD1.n11 171.744
R809 VDD1.n16 VDD1.n11 171.744
R810 VDD1.n80 VDD1.n16 171.744
R811 VDD1.n80 VDD1.n79 171.744
R812 VDD1.n79 VDD1.n17 171.744
R813 VDD1.n72 VDD1.n17 171.744
R814 VDD1.n72 VDD1.n71 171.744
R815 VDD1.n71 VDD1.n21 171.744
R816 VDD1.n64 VDD1.n21 171.744
R817 VDD1.n64 VDD1.n63 171.744
R818 VDD1.n63 VDD1.n25 171.744
R819 VDD1.n56 VDD1.n25 171.744
R820 VDD1.n56 VDD1.n55 171.744
R821 VDD1.n55 VDD1.n29 171.744
R822 VDD1.n48 VDD1.n29 171.744
R823 VDD1.n48 VDD1.n47 171.744
R824 VDD1.n47 VDD1.n33 171.744
R825 VDD1.n40 VDD1.n33 171.744
R826 VDD1.n40 VDD1.n39 171.744
R827 VDD1.n147 VDD1.n146 171.744
R828 VDD1.n147 VDD1.n140 171.744
R829 VDD1.n154 VDD1.n140 171.744
R830 VDD1.n155 VDD1.n154 171.744
R831 VDD1.n155 VDD1.n136 171.744
R832 VDD1.n162 VDD1.n136 171.744
R833 VDD1.n163 VDD1.n162 171.744
R834 VDD1.n163 VDD1.n132 171.744
R835 VDD1.n170 VDD1.n132 171.744
R836 VDD1.n171 VDD1.n170 171.744
R837 VDD1.n171 VDD1.n128 171.744
R838 VDD1.n178 VDD1.n128 171.744
R839 VDD1.n179 VDD1.n178 171.744
R840 VDD1.n179 VDD1.n124 171.744
R841 VDD1.n187 VDD1.n124 171.744
R842 VDD1.n188 VDD1.n187 171.744
R843 VDD1.n189 VDD1.n188 171.744
R844 VDD1.n189 VDD1.n120 171.744
R845 VDD1.n196 VDD1.n120 171.744
R846 VDD1.n197 VDD1.n196 171.744
R847 VDD1.n197 VDD1.n116 171.744
R848 VDD1.n204 VDD1.n116 171.744
R849 VDD1.n205 VDD1.n204 171.744
R850 VDD1.n205 VDD1.n112 171.744
R851 VDD1.n212 VDD1.n112 171.744
R852 VDD1.n213 VDD1.n212 171.744
R853 VDD1.n39 VDD1.t0 85.8723
R854 VDD1.n146 VDD1.t5 85.8723
R855 VDD1.n219 VDD1.n218 68.5952
R856 VDD1.n221 VDD1.n220 68.1096
R857 VDD1 VDD1.n108 50.5452
R858 VDD1.n219 VDD1.n217 50.4316
R859 VDD1.n221 VDD1.n219 49.378
R860 VDD1.n38 VDD1.n37 16.3895
R861 VDD1.n145 VDD1.n144 16.3895
R862 VDD1.n14 VDD1.n12 13.1884
R863 VDD1.n190 VDD1.n121 13.1884
R864 VDD1.n86 VDD1.n85 12.8005
R865 VDD1.n82 VDD1.n81 12.8005
R866 VDD1.n41 VDD1.n36 12.8005
R867 VDD1.n148 VDD1.n143 12.8005
R868 VDD1.n191 VDD1.n123 12.8005
R869 VDD1.n195 VDD1.n194 12.8005
R870 VDD1.n89 VDD1.n10 12.0247
R871 VDD1.n78 VDD1.n15 12.0247
R872 VDD1.n42 VDD1.n34 12.0247
R873 VDD1.n149 VDD1.n141 12.0247
R874 VDD1.n186 VDD1.n185 12.0247
R875 VDD1.n198 VDD1.n119 12.0247
R876 VDD1.n90 VDD1.n8 11.249
R877 VDD1.n77 VDD1.n18 11.249
R878 VDD1.n46 VDD1.n45 11.249
R879 VDD1.n153 VDD1.n152 11.249
R880 VDD1.n184 VDD1.n125 11.249
R881 VDD1.n199 VDD1.n117 11.249
R882 VDD1.n94 VDD1.n93 10.4732
R883 VDD1.n74 VDD1.n73 10.4732
R884 VDD1.n49 VDD1.n32 10.4732
R885 VDD1.n156 VDD1.n139 10.4732
R886 VDD1.n181 VDD1.n180 10.4732
R887 VDD1.n203 VDD1.n202 10.4732
R888 VDD1.n97 VDD1.n6 9.69747
R889 VDD1.n70 VDD1.n20 9.69747
R890 VDD1.n50 VDD1.n30 9.69747
R891 VDD1.n157 VDD1.n137 9.69747
R892 VDD1.n177 VDD1.n127 9.69747
R893 VDD1.n206 VDD1.n115 9.69747
R894 VDD1.n108 VDD1.n107 9.45567
R895 VDD1.n217 VDD1.n216 9.45567
R896 VDD1.n24 VDD1.n23 9.3005
R897 VDD1.n67 VDD1.n66 9.3005
R898 VDD1.n69 VDD1.n68 9.3005
R899 VDD1.n20 VDD1.n19 9.3005
R900 VDD1.n75 VDD1.n74 9.3005
R901 VDD1.n77 VDD1.n76 9.3005
R902 VDD1.n15 VDD1.n13 9.3005
R903 VDD1.n83 VDD1.n82 9.3005
R904 VDD1.n107 VDD1.n106 9.3005
R905 VDD1.n2 VDD1.n1 9.3005
R906 VDD1.n101 VDD1.n100 9.3005
R907 VDD1.n99 VDD1.n98 9.3005
R908 VDD1.n6 VDD1.n5 9.3005
R909 VDD1.n93 VDD1.n92 9.3005
R910 VDD1.n91 VDD1.n90 9.3005
R911 VDD1.n10 VDD1.n9 9.3005
R912 VDD1.n85 VDD1.n84 9.3005
R913 VDD1.n61 VDD1.n60 9.3005
R914 VDD1.n59 VDD1.n58 9.3005
R915 VDD1.n28 VDD1.n27 9.3005
R916 VDD1.n53 VDD1.n52 9.3005
R917 VDD1.n51 VDD1.n50 9.3005
R918 VDD1.n32 VDD1.n31 9.3005
R919 VDD1.n45 VDD1.n44 9.3005
R920 VDD1.n43 VDD1.n42 9.3005
R921 VDD1.n36 VDD1.n35 9.3005
R922 VDD1.n216 VDD1.n215 9.3005
R923 VDD1.n210 VDD1.n209 9.3005
R924 VDD1.n208 VDD1.n207 9.3005
R925 VDD1.n115 VDD1.n114 9.3005
R926 VDD1.n202 VDD1.n201 9.3005
R927 VDD1.n200 VDD1.n199 9.3005
R928 VDD1.n119 VDD1.n118 9.3005
R929 VDD1.n194 VDD1.n193 9.3005
R930 VDD1.n166 VDD1.n165 9.3005
R931 VDD1.n135 VDD1.n134 9.3005
R932 VDD1.n160 VDD1.n159 9.3005
R933 VDD1.n158 VDD1.n157 9.3005
R934 VDD1.n139 VDD1.n138 9.3005
R935 VDD1.n152 VDD1.n151 9.3005
R936 VDD1.n150 VDD1.n149 9.3005
R937 VDD1.n143 VDD1.n142 9.3005
R938 VDD1.n168 VDD1.n167 9.3005
R939 VDD1.n131 VDD1.n130 9.3005
R940 VDD1.n174 VDD1.n173 9.3005
R941 VDD1.n176 VDD1.n175 9.3005
R942 VDD1.n127 VDD1.n126 9.3005
R943 VDD1.n182 VDD1.n181 9.3005
R944 VDD1.n184 VDD1.n183 9.3005
R945 VDD1.n185 VDD1.n122 9.3005
R946 VDD1.n192 VDD1.n191 9.3005
R947 VDD1.n111 VDD1.n110 9.3005
R948 VDD1.n98 VDD1.n4 8.92171
R949 VDD1.n69 VDD1.n22 8.92171
R950 VDD1.n54 VDD1.n53 8.92171
R951 VDD1.n161 VDD1.n160 8.92171
R952 VDD1.n176 VDD1.n129 8.92171
R953 VDD1.n207 VDD1.n113 8.92171
R954 VDD1.n102 VDD1.n101 8.14595
R955 VDD1.n66 VDD1.n65 8.14595
R956 VDD1.n57 VDD1.n28 8.14595
R957 VDD1.n164 VDD1.n135 8.14595
R958 VDD1.n173 VDD1.n172 8.14595
R959 VDD1.n211 VDD1.n210 8.14595
R960 VDD1.n108 VDD1.n0 7.3702
R961 VDD1.n105 VDD1.n2 7.3702
R962 VDD1.n62 VDD1.n24 7.3702
R963 VDD1.n58 VDD1.n26 7.3702
R964 VDD1.n165 VDD1.n133 7.3702
R965 VDD1.n169 VDD1.n131 7.3702
R966 VDD1.n214 VDD1.n111 7.3702
R967 VDD1.n217 VDD1.n109 7.3702
R968 VDD1.n106 VDD1.n0 6.59444
R969 VDD1.n106 VDD1.n105 6.59444
R970 VDD1.n62 VDD1.n61 6.59444
R971 VDD1.n61 VDD1.n26 6.59444
R972 VDD1.n168 VDD1.n133 6.59444
R973 VDD1.n169 VDD1.n168 6.59444
R974 VDD1.n215 VDD1.n214 6.59444
R975 VDD1.n215 VDD1.n109 6.59444
R976 VDD1.n102 VDD1.n2 5.81868
R977 VDD1.n65 VDD1.n24 5.81868
R978 VDD1.n58 VDD1.n57 5.81868
R979 VDD1.n165 VDD1.n164 5.81868
R980 VDD1.n172 VDD1.n131 5.81868
R981 VDD1.n211 VDD1.n111 5.81868
R982 VDD1.n101 VDD1.n4 5.04292
R983 VDD1.n66 VDD1.n22 5.04292
R984 VDD1.n54 VDD1.n28 5.04292
R985 VDD1.n161 VDD1.n135 5.04292
R986 VDD1.n173 VDD1.n129 5.04292
R987 VDD1.n210 VDD1.n113 5.04292
R988 VDD1.n98 VDD1.n97 4.26717
R989 VDD1.n70 VDD1.n69 4.26717
R990 VDD1.n53 VDD1.n30 4.26717
R991 VDD1.n160 VDD1.n137 4.26717
R992 VDD1.n177 VDD1.n176 4.26717
R993 VDD1.n207 VDD1.n206 4.26717
R994 VDD1.n37 VDD1.n35 3.70982
R995 VDD1.n144 VDD1.n142 3.70982
R996 VDD1.n94 VDD1.n6 3.49141
R997 VDD1.n73 VDD1.n20 3.49141
R998 VDD1.n50 VDD1.n49 3.49141
R999 VDD1.n157 VDD1.n156 3.49141
R1000 VDD1.n180 VDD1.n127 3.49141
R1001 VDD1.n203 VDD1.n115 3.49141
R1002 VDD1.n93 VDD1.n8 2.71565
R1003 VDD1.n74 VDD1.n18 2.71565
R1004 VDD1.n46 VDD1.n32 2.71565
R1005 VDD1.n153 VDD1.n139 2.71565
R1006 VDD1.n181 VDD1.n125 2.71565
R1007 VDD1.n202 VDD1.n117 2.71565
R1008 VDD1.n90 VDD1.n89 1.93989
R1009 VDD1.n78 VDD1.n77 1.93989
R1010 VDD1.n45 VDD1.n34 1.93989
R1011 VDD1.n152 VDD1.n141 1.93989
R1012 VDD1.n186 VDD1.n184 1.93989
R1013 VDD1.n199 VDD1.n198 1.93989
R1014 VDD1.n220 VDD1.t3 1.65218
R1015 VDD1.n220 VDD1.t4 1.65218
R1016 VDD1.n218 VDD1.t2 1.65218
R1017 VDD1.n218 VDD1.t1 1.65218
R1018 VDD1.n86 VDD1.n10 1.16414
R1019 VDD1.n81 VDD1.n15 1.16414
R1020 VDD1.n42 VDD1.n41 1.16414
R1021 VDD1.n149 VDD1.n148 1.16414
R1022 VDD1.n185 VDD1.n123 1.16414
R1023 VDD1.n195 VDD1.n119 1.16414
R1024 VDD1 VDD1.n221 0.483259
R1025 VDD1.n85 VDD1.n12 0.388379
R1026 VDD1.n82 VDD1.n14 0.388379
R1027 VDD1.n38 VDD1.n36 0.388379
R1028 VDD1.n145 VDD1.n143 0.388379
R1029 VDD1.n191 VDD1.n190 0.388379
R1030 VDD1.n194 VDD1.n121 0.388379
R1031 VDD1.n107 VDD1.n1 0.155672
R1032 VDD1.n100 VDD1.n1 0.155672
R1033 VDD1.n100 VDD1.n99 0.155672
R1034 VDD1.n99 VDD1.n5 0.155672
R1035 VDD1.n92 VDD1.n5 0.155672
R1036 VDD1.n92 VDD1.n91 0.155672
R1037 VDD1.n91 VDD1.n9 0.155672
R1038 VDD1.n84 VDD1.n9 0.155672
R1039 VDD1.n84 VDD1.n83 0.155672
R1040 VDD1.n83 VDD1.n13 0.155672
R1041 VDD1.n76 VDD1.n13 0.155672
R1042 VDD1.n76 VDD1.n75 0.155672
R1043 VDD1.n75 VDD1.n19 0.155672
R1044 VDD1.n68 VDD1.n19 0.155672
R1045 VDD1.n68 VDD1.n67 0.155672
R1046 VDD1.n67 VDD1.n23 0.155672
R1047 VDD1.n60 VDD1.n23 0.155672
R1048 VDD1.n60 VDD1.n59 0.155672
R1049 VDD1.n59 VDD1.n27 0.155672
R1050 VDD1.n52 VDD1.n27 0.155672
R1051 VDD1.n52 VDD1.n51 0.155672
R1052 VDD1.n51 VDD1.n31 0.155672
R1053 VDD1.n44 VDD1.n31 0.155672
R1054 VDD1.n44 VDD1.n43 0.155672
R1055 VDD1.n43 VDD1.n35 0.155672
R1056 VDD1.n150 VDD1.n142 0.155672
R1057 VDD1.n151 VDD1.n150 0.155672
R1058 VDD1.n151 VDD1.n138 0.155672
R1059 VDD1.n158 VDD1.n138 0.155672
R1060 VDD1.n159 VDD1.n158 0.155672
R1061 VDD1.n159 VDD1.n134 0.155672
R1062 VDD1.n166 VDD1.n134 0.155672
R1063 VDD1.n167 VDD1.n166 0.155672
R1064 VDD1.n167 VDD1.n130 0.155672
R1065 VDD1.n174 VDD1.n130 0.155672
R1066 VDD1.n175 VDD1.n174 0.155672
R1067 VDD1.n175 VDD1.n126 0.155672
R1068 VDD1.n182 VDD1.n126 0.155672
R1069 VDD1.n183 VDD1.n182 0.155672
R1070 VDD1.n183 VDD1.n122 0.155672
R1071 VDD1.n192 VDD1.n122 0.155672
R1072 VDD1.n193 VDD1.n192 0.155672
R1073 VDD1.n193 VDD1.n118 0.155672
R1074 VDD1.n200 VDD1.n118 0.155672
R1075 VDD1.n201 VDD1.n200 0.155672
R1076 VDD1.n201 VDD1.n114 0.155672
R1077 VDD1.n208 VDD1.n114 0.155672
R1078 VDD1.n209 VDD1.n208 0.155672
R1079 VDD1.n209 VDD1.n110 0.155672
R1080 VDD1.n216 VDD1.n110 0.155672
R1081 VN.n3 VN.t5 249.788
R1082 VN.n17 VN.t3 249.788
R1083 VN.n4 VN.t4 217.564
R1084 VN.n12 VN.t2 217.564
R1085 VN.n18 VN.t1 217.564
R1086 VN.n26 VN.t0 217.564
R1087 VN.n25 VN.n14 161.3
R1088 VN.n24 VN.n23 161.3
R1089 VN.n22 VN.n15 161.3
R1090 VN.n21 VN.n20 161.3
R1091 VN.n19 VN.n16 161.3
R1092 VN.n11 VN.n0 161.3
R1093 VN.n10 VN.n9 161.3
R1094 VN.n8 VN.n1 161.3
R1095 VN.n7 VN.n6 161.3
R1096 VN.n5 VN.n2 161.3
R1097 VN.n13 VN.n12 98.1205
R1098 VN.n27 VN.n26 98.1205
R1099 VN.n4 VN.n3 59.417
R1100 VN.n18 VN.n17 59.417
R1101 VN VN.n27 53.0853
R1102 VN.n10 VN.n1 41.0614
R1103 VN.n24 VN.n15 41.0614
R1104 VN.n6 VN.n1 40.0926
R1105 VN.n20 VN.n15 40.0926
R1106 VN.n6 VN.n5 24.5923
R1107 VN.n11 VN.n10 24.5923
R1108 VN.n20 VN.n19 24.5923
R1109 VN.n25 VN.n24 24.5923
R1110 VN.n12 VN.n11 12.7883
R1111 VN.n26 VN.n25 12.7883
R1112 VN.n5 VN.n4 12.2964
R1113 VN.n19 VN.n18 12.2964
R1114 VN.n17 VN.n16 9.65766
R1115 VN.n3 VN.n2 9.65766
R1116 VN.n27 VN.n14 0.278335
R1117 VN.n13 VN.n0 0.278335
R1118 VN.n23 VN.n14 0.189894
R1119 VN.n23 VN.n22 0.189894
R1120 VN.n22 VN.n21 0.189894
R1121 VN.n21 VN.n16 0.189894
R1122 VN.n7 VN.n2 0.189894
R1123 VN.n8 VN.n7 0.189894
R1124 VN.n9 VN.n8 0.189894
R1125 VN.n9 VN.n0 0.189894
R1126 VN VN.n13 0.153485
R1127 VDD2.n215 VDD2.n111 756.745
R1128 VDD2.n104 VDD2.n0 756.745
R1129 VDD2.n216 VDD2.n215 585
R1130 VDD2.n214 VDD2.n213 585
R1131 VDD2.n115 VDD2.n114 585
R1132 VDD2.n208 VDD2.n207 585
R1133 VDD2.n206 VDD2.n205 585
R1134 VDD2.n119 VDD2.n118 585
R1135 VDD2.n200 VDD2.n199 585
R1136 VDD2.n198 VDD2.n197 585
R1137 VDD2.n123 VDD2.n122 585
R1138 VDD2.n127 VDD2.n125 585
R1139 VDD2.n192 VDD2.n191 585
R1140 VDD2.n190 VDD2.n189 585
R1141 VDD2.n129 VDD2.n128 585
R1142 VDD2.n184 VDD2.n183 585
R1143 VDD2.n182 VDD2.n181 585
R1144 VDD2.n133 VDD2.n132 585
R1145 VDD2.n176 VDD2.n175 585
R1146 VDD2.n174 VDD2.n173 585
R1147 VDD2.n137 VDD2.n136 585
R1148 VDD2.n168 VDD2.n167 585
R1149 VDD2.n166 VDD2.n165 585
R1150 VDD2.n141 VDD2.n140 585
R1151 VDD2.n160 VDD2.n159 585
R1152 VDD2.n158 VDD2.n157 585
R1153 VDD2.n145 VDD2.n144 585
R1154 VDD2.n152 VDD2.n151 585
R1155 VDD2.n150 VDD2.n149 585
R1156 VDD2.n37 VDD2.n36 585
R1157 VDD2.n39 VDD2.n38 585
R1158 VDD2.n32 VDD2.n31 585
R1159 VDD2.n45 VDD2.n44 585
R1160 VDD2.n47 VDD2.n46 585
R1161 VDD2.n28 VDD2.n27 585
R1162 VDD2.n53 VDD2.n52 585
R1163 VDD2.n55 VDD2.n54 585
R1164 VDD2.n24 VDD2.n23 585
R1165 VDD2.n61 VDD2.n60 585
R1166 VDD2.n63 VDD2.n62 585
R1167 VDD2.n20 VDD2.n19 585
R1168 VDD2.n69 VDD2.n68 585
R1169 VDD2.n71 VDD2.n70 585
R1170 VDD2.n16 VDD2.n15 585
R1171 VDD2.n78 VDD2.n77 585
R1172 VDD2.n79 VDD2.n14 585
R1173 VDD2.n81 VDD2.n80 585
R1174 VDD2.n12 VDD2.n11 585
R1175 VDD2.n87 VDD2.n86 585
R1176 VDD2.n89 VDD2.n88 585
R1177 VDD2.n8 VDD2.n7 585
R1178 VDD2.n95 VDD2.n94 585
R1179 VDD2.n97 VDD2.n96 585
R1180 VDD2.n4 VDD2.n3 585
R1181 VDD2.n103 VDD2.n102 585
R1182 VDD2.n105 VDD2.n104 585
R1183 VDD2.n148 VDD2.t5 327.466
R1184 VDD2.n35 VDD2.t0 327.466
R1185 VDD2.n215 VDD2.n214 171.744
R1186 VDD2.n214 VDD2.n114 171.744
R1187 VDD2.n207 VDD2.n114 171.744
R1188 VDD2.n207 VDD2.n206 171.744
R1189 VDD2.n206 VDD2.n118 171.744
R1190 VDD2.n199 VDD2.n118 171.744
R1191 VDD2.n199 VDD2.n198 171.744
R1192 VDD2.n198 VDD2.n122 171.744
R1193 VDD2.n127 VDD2.n122 171.744
R1194 VDD2.n191 VDD2.n127 171.744
R1195 VDD2.n191 VDD2.n190 171.744
R1196 VDD2.n190 VDD2.n128 171.744
R1197 VDD2.n183 VDD2.n128 171.744
R1198 VDD2.n183 VDD2.n182 171.744
R1199 VDD2.n182 VDD2.n132 171.744
R1200 VDD2.n175 VDD2.n132 171.744
R1201 VDD2.n175 VDD2.n174 171.744
R1202 VDD2.n174 VDD2.n136 171.744
R1203 VDD2.n167 VDD2.n136 171.744
R1204 VDD2.n167 VDD2.n166 171.744
R1205 VDD2.n166 VDD2.n140 171.744
R1206 VDD2.n159 VDD2.n140 171.744
R1207 VDD2.n159 VDD2.n158 171.744
R1208 VDD2.n158 VDD2.n144 171.744
R1209 VDD2.n151 VDD2.n144 171.744
R1210 VDD2.n151 VDD2.n150 171.744
R1211 VDD2.n38 VDD2.n37 171.744
R1212 VDD2.n38 VDD2.n31 171.744
R1213 VDD2.n45 VDD2.n31 171.744
R1214 VDD2.n46 VDD2.n45 171.744
R1215 VDD2.n46 VDD2.n27 171.744
R1216 VDD2.n53 VDD2.n27 171.744
R1217 VDD2.n54 VDD2.n53 171.744
R1218 VDD2.n54 VDD2.n23 171.744
R1219 VDD2.n61 VDD2.n23 171.744
R1220 VDD2.n62 VDD2.n61 171.744
R1221 VDD2.n62 VDD2.n19 171.744
R1222 VDD2.n69 VDD2.n19 171.744
R1223 VDD2.n70 VDD2.n69 171.744
R1224 VDD2.n70 VDD2.n15 171.744
R1225 VDD2.n78 VDD2.n15 171.744
R1226 VDD2.n79 VDD2.n78 171.744
R1227 VDD2.n80 VDD2.n79 171.744
R1228 VDD2.n80 VDD2.n11 171.744
R1229 VDD2.n87 VDD2.n11 171.744
R1230 VDD2.n88 VDD2.n87 171.744
R1231 VDD2.n88 VDD2.n7 171.744
R1232 VDD2.n95 VDD2.n7 171.744
R1233 VDD2.n96 VDD2.n95 171.744
R1234 VDD2.n96 VDD2.n3 171.744
R1235 VDD2.n103 VDD2.n3 171.744
R1236 VDD2.n104 VDD2.n103 171.744
R1237 VDD2.n150 VDD2.t5 85.8723
R1238 VDD2.n37 VDD2.t0 85.8723
R1239 VDD2.n110 VDD2.n109 68.5952
R1240 VDD2 VDD2.n221 68.5923
R1241 VDD2.n110 VDD2.n108 50.4316
R1242 VDD2.n220 VDD2.n219 48.8641
R1243 VDD2.n220 VDD2.n110 47.7131
R1244 VDD2.n149 VDD2.n148 16.3895
R1245 VDD2.n36 VDD2.n35 16.3895
R1246 VDD2.n125 VDD2.n123 13.1884
R1247 VDD2.n81 VDD2.n12 13.1884
R1248 VDD2.n197 VDD2.n196 12.8005
R1249 VDD2.n193 VDD2.n192 12.8005
R1250 VDD2.n152 VDD2.n147 12.8005
R1251 VDD2.n39 VDD2.n34 12.8005
R1252 VDD2.n82 VDD2.n14 12.8005
R1253 VDD2.n86 VDD2.n85 12.8005
R1254 VDD2.n200 VDD2.n121 12.0247
R1255 VDD2.n189 VDD2.n126 12.0247
R1256 VDD2.n153 VDD2.n145 12.0247
R1257 VDD2.n40 VDD2.n32 12.0247
R1258 VDD2.n77 VDD2.n76 12.0247
R1259 VDD2.n89 VDD2.n10 12.0247
R1260 VDD2.n201 VDD2.n119 11.249
R1261 VDD2.n188 VDD2.n129 11.249
R1262 VDD2.n157 VDD2.n156 11.249
R1263 VDD2.n44 VDD2.n43 11.249
R1264 VDD2.n75 VDD2.n16 11.249
R1265 VDD2.n90 VDD2.n8 11.249
R1266 VDD2.n205 VDD2.n204 10.4732
R1267 VDD2.n185 VDD2.n184 10.4732
R1268 VDD2.n160 VDD2.n143 10.4732
R1269 VDD2.n47 VDD2.n30 10.4732
R1270 VDD2.n72 VDD2.n71 10.4732
R1271 VDD2.n94 VDD2.n93 10.4732
R1272 VDD2.n208 VDD2.n117 9.69747
R1273 VDD2.n181 VDD2.n131 9.69747
R1274 VDD2.n161 VDD2.n141 9.69747
R1275 VDD2.n48 VDD2.n28 9.69747
R1276 VDD2.n68 VDD2.n18 9.69747
R1277 VDD2.n97 VDD2.n6 9.69747
R1278 VDD2.n219 VDD2.n218 9.45567
R1279 VDD2.n108 VDD2.n107 9.45567
R1280 VDD2.n135 VDD2.n134 9.3005
R1281 VDD2.n178 VDD2.n177 9.3005
R1282 VDD2.n180 VDD2.n179 9.3005
R1283 VDD2.n131 VDD2.n130 9.3005
R1284 VDD2.n186 VDD2.n185 9.3005
R1285 VDD2.n188 VDD2.n187 9.3005
R1286 VDD2.n126 VDD2.n124 9.3005
R1287 VDD2.n194 VDD2.n193 9.3005
R1288 VDD2.n218 VDD2.n217 9.3005
R1289 VDD2.n113 VDD2.n112 9.3005
R1290 VDD2.n212 VDD2.n211 9.3005
R1291 VDD2.n210 VDD2.n209 9.3005
R1292 VDD2.n117 VDD2.n116 9.3005
R1293 VDD2.n204 VDD2.n203 9.3005
R1294 VDD2.n202 VDD2.n201 9.3005
R1295 VDD2.n121 VDD2.n120 9.3005
R1296 VDD2.n196 VDD2.n195 9.3005
R1297 VDD2.n172 VDD2.n171 9.3005
R1298 VDD2.n170 VDD2.n169 9.3005
R1299 VDD2.n139 VDD2.n138 9.3005
R1300 VDD2.n164 VDD2.n163 9.3005
R1301 VDD2.n162 VDD2.n161 9.3005
R1302 VDD2.n143 VDD2.n142 9.3005
R1303 VDD2.n156 VDD2.n155 9.3005
R1304 VDD2.n154 VDD2.n153 9.3005
R1305 VDD2.n147 VDD2.n146 9.3005
R1306 VDD2.n107 VDD2.n106 9.3005
R1307 VDD2.n101 VDD2.n100 9.3005
R1308 VDD2.n99 VDD2.n98 9.3005
R1309 VDD2.n6 VDD2.n5 9.3005
R1310 VDD2.n93 VDD2.n92 9.3005
R1311 VDD2.n91 VDD2.n90 9.3005
R1312 VDD2.n10 VDD2.n9 9.3005
R1313 VDD2.n85 VDD2.n84 9.3005
R1314 VDD2.n57 VDD2.n56 9.3005
R1315 VDD2.n26 VDD2.n25 9.3005
R1316 VDD2.n51 VDD2.n50 9.3005
R1317 VDD2.n49 VDD2.n48 9.3005
R1318 VDD2.n30 VDD2.n29 9.3005
R1319 VDD2.n43 VDD2.n42 9.3005
R1320 VDD2.n41 VDD2.n40 9.3005
R1321 VDD2.n34 VDD2.n33 9.3005
R1322 VDD2.n59 VDD2.n58 9.3005
R1323 VDD2.n22 VDD2.n21 9.3005
R1324 VDD2.n65 VDD2.n64 9.3005
R1325 VDD2.n67 VDD2.n66 9.3005
R1326 VDD2.n18 VDD2.n17 9.3005
R1327 VDD2.n73 VDD2.n72 9.3005
R1328 VDD2.n75 VDD2.n74 9.3005
R1329 VDD2.n76 VDD2.n13 9.3005
R1330 VDD2.n83 VDD2.n82 9.3005
R1331 VDD2.n2 VDD2.n1 9.3005
R1332 VDD2.n209 VDD2.n115 8.92171
R1333 VDD2.n180 VDD2.n133 8.92171
R1334 VDD2.n165 VDD2.n164 8.92171
R1335 VDD2.n52 VDD2.n51 8.92171
R1336 VDD2.n67 VDD2.n20 8.92171
R1337 VDD2.n98 VDD2.n4 8.92171
R1338 VDD2.n213 VDD2.n212 8.14595
R1339 VDD2.n177 VDD2.n176 8.14595
R1340 VDD2.n168 VDD2.n139 8.14595
R1341 VDD2.n55 VDD2.n26 8.14595
R1342 VDD2.n64 VDD2.n63 8.14595
R1343 VDD2.n102 VDD2.n101 8.14595
R1344 VDD2.n219 VDD2.n111 7.3702
R1345 VDD2.n216 VDD2.n113 7.3702
R1346 VDD2.n173 VDD2.n135 7.3702
R1347 VDD2.n169 VDD2.n137 7.3702
R1348 VDD2.n56 VDD2.n24 7.3702
R1349 VDD2.n60 VDD2.n22 7.3702
R1350 VDD2.n105 VDD2.n2 7.3702
R1351 VDD2.n108 VDD2.n0 7.3702
R1352 VDD2.n217 VDD2.n111 6.59444
R1353 VDD2.n217 VDD2.n216 6.59444
R1354 VDD2.n173 VDD2.n172 6.59444
R1355 VDD2.n172 VDD2.n137 6.59444
R1356 VDD2.n59 VDD2.n24 6.59444
R1357 VDD2.n60 VDD2.n59 6.59444
R1358 VDD2.n106 VDD2.n105 6.59444
R1359 VDD2.n106 VDD2.n0 6.59444
R1360 VDD2.n213 VDD2.n113 5.81868
R1361 VDD2.n176 VDD2.n135 5.81868
R1362 VDD2.n169 VDD2.n168 5.81868
R1363 VDD2.n56 VDD2.n55 5.81868
R1364 VDD2.n63 VDD2.n22 5.81868
R1365 VDD2.n102 VDD2.n2 5.81868
R1366 VDD2.n212 VDD2.n115 5.04292
R1367 VDD2.n177 VDD2.n133 5.04292
R1368 VDD2.n165 VDD2.n139 5.04292
R1369 VDD2.n52 VDD2.n26 5.04292
R1370 VDD2.n64 VDD2.n20 5.04292
R1371 VDD2.n101 VDD2.n4 5.04292
R1372 VDD2.n209 VDD2.n208 4.26717
R1373 VDD2.n181 VDD2.n180 4.26717
R1374 VDD2.n164 VDD2.n141 4.26717
R1375 VDD2.n51 VDD2.n28 4.26717
R1376 VDD2.n68 VDD2.n67 4.26717
R1377 VDD2.n98 VDD2.n97 4.26717
R1378 VDD2.n148 VDD2.n146 3.70982
R1379 VDD2.n35 VDD2.n33 3.70982
R1380 VDD2.n205 VDD2.n117 3.49141
R1381 VDD2.n184 VDD2.n131 3.49141
R1382 VDD2.n161 VDD2.n160 3.49141
R1383 VDD2.n48 VDD2.n47 3.49141
R1384 VDD2.n71 VDD2.n18 3.49141
R1385 VDD2.n94 VDD2.n6 3.49141
R1386 VDD2.n204 VDD2.n119 2.71565
R1387 VDD2.n185 VDD2.n129 2.71565
R1388 VDD2.n157 VDD2.n143 2.71565
R1389 VDD2.n44 VDD2.n30 2.71565
R1390 VDD2.n72 VDD2.n16 2.71565
R1391 VDD2.n93 VDD2.n8 2.71565
R1392 VDD2.n201 VDD2.n200 1.93989
R1393 VDD2.n189 VDD2.n188 1.93989
R1394 VDD2.n156 VDD2.n145 1.93989
R1395 VDD2.n43 VDD2.n32 1.93989
R1396 VDD2.n77 VDD2.n75 1.93989
R1397 VDD2.n90 VDD2.n89 1.93989
R1398 VDD2 VDD2.n220 1.68153
R1399 VDD2.n221 VDD2.t4 1.65218
R1400 VDD2.n221 VDD2.t2 1.65218
R1401 VDD2.n109 VDD2.t1 1.65218
R1402 VDD2.n109 VDD2.t3 1.65218
R1403 VDD2.n197 VDD2.n121 1.16414
R1404 VDD2.n192 VDD2.n126 1.16414
R1405 VDD2.n153 VDD2.n152 1.16414
R1406 VDD2.n40 VDD2.n39 1.16414
R1407 VDD2.n76 VDD2.n14 1.16414
R1408 VDD2.n86 VDD2.n10 1.16414
R1409 VDD2.n196 VDD2.n123 0.388379
R1410 VDD2.n193 VDD2.n125 0.388379
R1411 VDD2.n149 VDD2.n147 0.388379
R1412 VDD2.n36 VDD2.n34 0.388379
R1413 VDD2.n82 VDD2.n81 0.388379
R1414 VDD2.n85 VDD2.n12 0.388379
R1415 VDD2.n218 VDD2.n112 0.155672
R1416 VDD2.n211 VDD2.n112 0.155672
R1417 VDD2.n211 VDD2.n210 0.155672
R1418 VDD2.n210 VDD2.n116 0.155672
R1419 VDD2.n203 VDD2.n116 0.155672
R1420 VDD2.n203 VDD2.n202 0.155672
R1421 VDD2.n202 VDD2.n120 0.155672
R1422 VDD2.n195 VDD2.n120 0.155672
R1423 VDD2.n195 VDD2.n194 0.155672
R1424 VDD2.n194 VDD2.n124 0.155672
R1425 VDD2.n187 VDD2.n124 0.155672
R1426 VDD2.n187 VDD2.n186 0.155672
R1427 VDD2.n186 VDD2.n130 0.155672
R1428 VDD2.n179 VDD2.n130 0.155672
R1429 VDD2.n179 VDD2.n178 0.155672
R1430 VDD2.n178 VDD2.n134 0.155672
R1431 VDD2.n171 VDD2.n134 0.155672
R1432 VDD2.n171 VDD2.n170 0.155672
R1433 VDD2.n170 VDD2.n138 0.155672
R1434 VDD2.n163 VDD2.n138 0.155672
R1435 VDD2.n163 VDD2.n162 0.155672
R1436 VDD2.n162 VDD2.n142 0.155672
R1437 VDD2.n155 VDD2.n142 0.155672
R1438 VDD2.n155 VDD2.n154 0.155672
R1439 VDD2.n154 VDD2.n146 0.155672
R1440 VDD2.n41 VDD2.n33 0.155672
R1441 VDD2.n42 VDD2.n41 0.155672
R1442 VDD2.n42 VDD2.n29 0.155672
R1443 VDD2.n49 VDD2.n29 0.155672
R1444 VDD2.n50 VDD2.n49 0.155672
R1445 VDD2.n50 VDD2.n25 0.155672
R1446 VDD2.n57 VDD2.n25 0.155672
R1447 VDD2.n58 VDD2.n57 0.155672
R1448 VDD2.n58 VDD2.n21 0.155672
R1449 VDD2.n65 VDD2.n21 0.155672
R1450 VDD2.n66 VDD2.n65 0.155672
R1451 VDD2.n66 VDD2.n17 0.155672
R1452 VDD2.n73 VDD2.n17 0.155672
R1453 VDD2.n74 VDD2.n73 0.155672
R1454 VDD2.n74 VDD2.n13 0.155672
R1455 VDD2.n83 VDD2.n13 0.155672
R1456 VDD2.n84 VDD2.n83 0.155672
R1457 VDD2.n84 VDD2.n9 0.155672
R1458 VDD2.n91 VDD2.n9 0.155672
R1459 VDD2.n92 VDD2.n91 0.155672
R1460 VDD2.n92 VDD2.n5 0.155672
R1461 VDD2.n99 VDD2.n5 0.155672
R1462 VDD2.n100 VDD2.n99 0.155672
R1463 VDD2.n100 VDD2.n1 0.155672
R1464 VDD2.n107 VDD2.n1 0.155672
R1465 B.n486 B.n485 585
R1466 B.n484 B.n133 585
R1467 B.n483 B.n482 585
R1468 B.n481 B.n134 585
R1469 B.n480 B.n479 585
R1470 B.n478 B.n135 585
R1471 B.n477 B.n476 585
R1472 B.n475 B.n136 585
R1473 B.n474 B.n473 585
R1474 B.n472 B.n137 585
R1475 B.n471 B.n470 585
R1476 B.n469 B.n138 585
R1477 B.n468 B.n467 585
R1478 B.n466 B.n139 585
R1479 B.n465 B.n464 585
R1480 B.n463 B.n140 585
R1481 B.n462 B.n461 585
R1482 B.n460 B.n141 585
R1483 B.n459 B.n458 585
R1484 B.n457 B.n142 585
R1485 B.n456 B.n455 585
R1486 B.n454 B.n143 585
R1487 B.n453 B.n452 585
R1488 B.n451 B.n144 585
R1489 B.n450 B.n449 585
R1490 B.n448 B.n145 585
R1491 B.n447 B.n446 585
R1492 B.n445 B.n146 585
R1493 B.n444 B.n443 585
R1494 B.n442 B.n147 585
R1495 B.n441 B.n440 585
R1496 B.n439 B.n148 585
R1497 B.n438 B.n437 585
R1498 B.n436 B.n149 585
R1499 B.n435 B.n434 585
R1500 B.n433 B.n150 585
R1501 B.n432 B.n431 585
R1502 B.n430 B.n151 585
R1503 B.n429 B.n428 585
R1504 B.n427 B.n152 585
R1505 B.n426 B.n425 585
R1506 B.n424 B.n153 585
R1507 B.n423 B.n422 585
R1508 B.n421 B.n154 585
R1509 B.n420 B.n419 585
R1510 B.n418 B.n155 585
R1511 B.n417 B.n416 585
R1512 B.n415 B.n156 585
R1513 B.n414 B.n413 585
R1514 B.n412 B.n157 585
R1515 B.n411 B.n410 585
R1516 B.n409 B.n158 585
R1517 B.n408 B.n407 585
R1518 B.n406 B.n159 585
R1519 B.n405 B.n404 585
R1520 B.n403 B.n160 585
R1521 B.n402 B.n401 585
R1522 B.n400 B.n161 585
R1523 B.n399 B.n398 585
R1524 B.n397 B.n162 585
R1525 B.n396 B.n395 585
R1526 B.n394 B.n163 585
R1527 B.n393 B.n392 585
R1528 B.n391 B.n164 585
R1529 B.n389 B.n388 585
R1530 B.n387 B.n167 585
R1531 B.n386 B.n385 585
R1532 B.n384 B.n168 585
R1533 B.n383 B.n382 585
R1534 B.n381 B.n169 585
R1535 B.n380 B.n379 585
R1536 B.n378 B.n170 585
R1537 B.n377 B.n376 585
R1538 B.n375 B.n171 585
R1539 B.n374 B.n373 585
R1540 B.n369 B.n172 585
R1541 B.n368 B.n367 585
R1542 B.n366 B.n173 585
R1543 B.n365 B.n364 585
R1544 B.n363 B.n174 585
R1545 B.n362 B.n361 585
R1546 B.n360 B.n175 585
R1547 B.n359 B.n358 585
R1548 B.n357 B.n176 585
R1549 B.n356 B.n355 585
R1550 B.n354 B.n177 585
R1551 B.n353 B.n352 585
R1552 B.n351 B.n178 585
R1553 B.n350 B.n349 585
R1554 B.n348 B.n179 585
R1555 B.n347 B.n346 585
R1556 B.n345 B.n180 585
R1557 B.n344 B.n343 585
R1558 B.n342 B.n181 585
R1559 B.n341 B.n340 585
R1560 B.n339 B.n182 585
R1561 B.n338 B.n337 585
R1562 B.n336 B.n183 585
R1563 B.n335 B.n334 585
R1564 B.n333 B.n184 585
R1565 B.n332 B.n331 585
R1566 B.n330 B.n185 585
R1567 B.n329 B.n328 585
R1568 B.n327 B.n186 585
R1569 B.n326 B.n325 585
R1570 B.n324 B.n187 585
R1571 B.n323 B.n322 585
R1572 B.n321 B.n188 585
R1573 B.n320 B.n319 585
R1574 B.n318 B.n189 585
R1575 B.n317 B.n316 585
R1576 B.n315 B.n190 585
R1577 B.n314 B.n313 585
R1578 B.n312 B.n191 585
R1579 B.n311 B.n310 585
R1580 B.n309 B.n192 585
R1581 B.n308 B.n307 585
R1582 B.n306 B.n193 585
R1583 B.n305 B.n304 585
R1584 B.n303 B.n194 585
R1585 B.n302 B.n301 585
R1586 B.n300 B.n195 585
R1587 B.n299 B.n298 585
R1588 B.n297 B.n196 585
R1589 B.n296 B.n295 585
R1590 B.n294 B.n197 585
R1591 B.n293 B.n292 585
R1592 B.n291 B.n198 585
R1593 B.n290 B.n289 585
R1594 B.n288 B.n199 585
R1595 B.n287 B.n286 585
R1596 B.n285 B.n200 585
R1597 B.n284 B.n283 585
R1598 B.n282 B.n201 585
R1599 B.n281 B.n280 585
R1600 B.n279 B.n202 585
R1601 B.n278 B.n277 585
R1602 B.n276 B.n203 585
R1603 B.n487 B.n132 585
R1604 B.n489 B.n488 585
R1605 B.n490 B.n131 585
R1606 B.n492 B.n491 585
R1607 B.n493 B.n130 585
R1608 B.n495 B.n494 585
R1609 B.n496 B.n129 585
R1610 B.n498 B.n497 585
R1611 B.n499 B.n128 585
R1612 B.n501 B.n500 585
R1613 B.n502 B.n127 585
R1614 B.n504 B.n503 585
R1615 B.n505 B.n126 585
R1616 B.n507 B.n506 585
R1617 B.n508 B.n125 585
R1618 B.n510 B.n509 585
R1619 B.n511 B.n124 585
R1620 B.n513 B.n512 585
R1621 B.n514 B.n123 585
R1622 B.n516 B.n515 585
R1623 B.n517 B.n122 585
R1624 B.n519 B.n518 585
R1625 B.n520 B.n121 585
R1626 B.n522 B.n521 585
R1627 B.n523 B.n120 585
R1628 B.n525 B.n524 585
R1629 B.n526 B.n119 585
R1630 B.n528 B.n527 585
R1631 B.n529 B.n118 585
R1632 B.n531 B.n530 585
R1633 B.n532 B.n117 585
R1634 B.n534 B.n533 585
R1635 B.n535 B.n116 585
R1636 B.n537 B.n536 585
R1637 B.n538 B.n115 585
R1638 B.n540 B.n539 585
R1639 B.n541 B.n114 585
R1640 B.n543 B.n542 585
R1641 B.n544 B.n113 585
R1642 B.n546 B.n545 585
R1643 B.n547 B.n112 585
R1644 B.n549 B.n548 585
R1645 B.n550 B.n111 585
R1646 B.n552 B.n551 585
R1647 B.n553 B.n110 585
R1648 B.n555 B.n554 585
R1649 B.n556 B.n109 585
R1650 B.n558 B.n557 585
R1651 B.n559 B.n108 585
R1652 B.n561 B.n560 585
R1653 B.n562 B.n107 585
R1654 B.n564 B.n563 585
R1655 B.n565 B.n106 585
R1656 B.n567 B.n566 585
R1657 B.n568 B.n105 585
R1658 B.n570 B.n569 585
R1659 B.n571 B.n104 585
R1660 B.n573 B.n572 585
R1661 B.n574 B.n103 585
R1662 B.n576 B.n575 585
R1663 B.n577 B.n102 585
R1664 B.n579 B.n578 585
R1665 B.n580 B.n101 585
R1666 B.n582 B.n581 585
R1667 B.n583 B.n100 585
R1668 B.n585 B.n584 585
R1669 B.n586 B.n99 585
R1670 B.n588 B.n587 585
R1671 B.n589 B.n98 585
R1672 B.n591 B.n590 585
R1673 B.n592 B.n97 585
R1674 B.n594 B.n593 585
R1675 B.n595 B.n96 585
R1676 B.n597 B.n596 585
R1677 B.n598 B.n95 585
R1678 B.n600 B.n599 585
R1679 B.n808 B.n807 585
R1680 B.n806 B.n21 585
R1681 B.n805 B.n804 585
R1682 B.n803 B.n22 585
R1683 B.n802 B.n801 585
R1684 B.n800 B.n23 585
R1685 B.n799 B.n798 585
R1686 B.n797 B.n24 585
R1687 B.n796 B.n795 585
R1688 B.n794 B.n25 585
R1689 B.n793 B.n792 585
R1690 B.n791 B.n26 585
R1691 B.n790 B.n789 585
R1692 B.n788 B.n27 585
R1693 B.n787 B.n786 585
R1694 B.n785 B.n28 585
R1695 B.n784 B.n783 585
R1696 B.n782 B.n29 585
R1697 B.n781 B.n780 585
R1698 B.n779 B.n30 585
R1699 B.n778 B.n777 585
R1700 B.n776 B.n31 585
R1701 B.n775 B.n774 585
R1702 B.n773 B.n32 585
R1703 B.n772 B.n771 585
R1704 B.n770 B.n33 585
R1705 B.n769 B.n768 585
R1706 B.n767 B.n34 585
R1707 B.n766 B.n765 585
R1708 B.n764 B.n35 585
R1709 B.n763 B.n762 585
R1710 B.n761 B.n36 585
R1711 B.n760 B.n759 585
R1712 B.n758 B.n37 585
R1713 B.n757 B.n756 585
R1714 B.n755 B.n38 585
R1715 B.n754 B.n753 585
R1716 B.n752 B.n39 585
R1717 B.n751 B.n750 585
R1718 B.n749 B.n40 585
R1719 B.n748 B.n747 585
R1720 B.n746 B.n41 585
R1721 B.n745 B.n744 585
R1722 B.n743 B.n42 585
R1723 B.n742 B.n741 585
R1724 B.n740 B.n43 585
R1725 B.n739 B.n738 585
R1726 B.n737 B.n44 585
R1727 B.n736 B.n735 585
R1728 B.n734 B.n45 585
R1729 B.n733 B.n732 585
R1730 B.n731 B.n46 585
R1731 B.n730 B.n729 585
R1732 B.n728 B.n47 585
R1733 B.n727 B.n726 585
R1734 B.n725 B.n48 585
R1735 B.n724 B.n723 585
R1736 B.n722 B.n49 585
R1737 B.n721 B.n720 585
R1738 B.n719 B.n50 585
R1739 B.n718 B.n717 585
R1740 B.n716 B.n51 585
R1741 B.n715 B.n714 585
R1742 B.n713 B.n52 585
R1743 B.n712 B.n711 585
R1744 B.n710 B.n53 585
R1745 B.n709 B.n708 585
R1746 B.n707 B.n57 585
R1747 B.n706 B.n705 585
R1748 B.n704 B.n58 585
R1749 B.n703 B.n702 585
R1750 B.n701 B.n59 585
R1751 B.n700 B.n699 585
R1752 B.n698 B.n60 585
R1753 B.n696 B.n695 585
R1754 B.n694 B.n63 585
R1755 B.n693 B.n692 585
R1756 B.n691 B.n64 585
R1757 B.n690 B.n689 585
R1758 B.n688 B.n65 585
R1759 B.n687 B.n686 585
R1760 B.n685 B.n66 585
R1761 B.n684 B.n683 585
R1762 B.n682 B.n67 585
R1763 B.n681 B.n680 585
R1764 B.n679 B.n68 585
R1765 B.n678 B.n677 585
R1766 B.n676 B.n69 585
R1767 B.n675 B.n674 585
R1768 B.n673 B.n70 585
R1769 B.n672 B.n671 585
R1770 B.n670 B.n71 585
R1771 B.n669 B.n668 585
R1772 B.n667 B.n72 585
R1773 B.n666 B.n665 585
R1774 B.n664 B.n73 585
R1775 B.n663 B.n662 585
R1776 B.n661 B.n74 585
R1777 B.n660 B.n659 585
R1778 B.n658 B.n75 585
R1779 B.n657 B.n656 585
R1780 B.n655 B.n76 585
R1781 B.n654 B.n653 585
R1782 B.n652 B.n77 585
R1783 B.n651 B.n650 585
R1784 B.n649 B.n78 585
R1785 B.n648 B.n647 585
R1786 B.n646 B.n79 585
R1787 B.n645 B.n644 585
R1788 B.n643 B.n80 585
R1789 B.n642 B.n641 585
R1790 B.n640 B.n81 585
R1791 B.n639 B.n638 585
R1792 B.n637 B.n82 585
R1793 B.n636 B.n635 585
R1794 B.n634 B.n83 585
R1795 B.n633 B.n632 585
R1796 B.n631 B.n84 585
R1797 B.n630 B.n629 585
R1798 B.n628 B.n85 585
R1799 B.n627 B.n626 585
R1800 B.n625 B.n86 585
R1801 B.n624 B.n623 585
R1802 B.n622 B.n87 585
R1803 B.n621 B.n620 585
R1804 B.n619 B.n88 585
R1805 B.n618 B.n617 585
R1806 B.n616 B.n89 585
R1807 B.n615 B.n614 585
R1808 B.n613 B.n90 585
R1809 B.n612 B.n611 585
R1810 B.n610 B.n91 585
R1811 B.n609 B.n608 585
R1812 B.n607 B.n92 585
R1813 B.n606 B.n605 585
R1814 B.n604 B.n93 585
R1815 B.n603 B.n602 585
R1816 B.n601 B.n94 585
R1817 B.n809 B.n20 585
R1818 B.n811 B.n810 585
R1819 B.n812 B.n19 585
R1820 B.n814 B.n813 585
R1821 B.n815 B.n18 585
R1822 B.n817 B.n816 585
R1823 B.n818 B.n17 585
R1824 B.n820 B.n819 585
R1825 B.n821 B.n16 585
R1826 B.n823 B.n822 585
R1827 B.n824 B.n15 585
R1828 B.n826 B.n825 585
R1829 B.n827 B.n14 585
R1830 B.n829 B.n828 585
R1831 B.n830 B.n13 585
R1832 B.n832 B.n831 585
R1833 B.n833 B.n12 585
R1834 B.n835 B.n834 585
R1835 B.n836 B.n11 585
R1836 B.n838 B.n837 585
R1837 B.n839 B.n10 585
R1838 B.n841 B.n840 585
R1839 B.n842 B.n9 585
R1840 B.n844 B.n843 585
R1841 B.n845 B.n8 585
R1842 B.n847 B.n846 585
R1843 B.n848 B.n7 585
R1844 B.n850 B.n849 585
R1845 B.n851 B.n6 585
R1846 B.n853 B.n852 585
R1847 B.n854 B.n5 585
R1848 B.n856 B.n855 585
R1849 B.n857 B.n4 585
R1850 B.n859 B.n858 585
R1851 B.n860 B.n3 585
R1852 B.n862 B.n861 585
R1853 B.n863 B.n0 585
R1854 B.n2 B.n1 585
R1855 B.n222 B.n221 585
R1856 B.n224 B.n223 585
R1857 B.n225 B.n220 585
R1858 B.n227 B.n226 585
R1859 B.n228 B.n219 585
R1860 B.n230 B.n229 585
R1861 B.n231 B.n218 585
R1862 B.n233 B.n232 585
R1863 B.n234 B.n217 585
R1864 B.n236 B.n235 585
R1865 B.n237 B.n216 585
R1866 B.n239 B.n238 585
R1867 B.n240 B.n215 585
R1868 B.n242 B.n241 585
R1869 B.n243 B.n214 585
R1870 B.n245 B.n244 585
R1871 B.n246 B.n213 585
R1872 B.n248 B.n247 585
R1873 B.n249 B.n212 585
R1874 B.n251 B.n250 585
R1875 B.n252 B.n211 585
R1876 B.n254 B.n253 585
R1877 B.n255 B.n210 585
R1878 B.n257 B.n256 585
R1879 B.n258 B.n209 585
R1880 B.n260 B.n259 585
R1881 B.n261 B.n208 585
R1882 B.n263 B.n262 585
R1883 B.n264 B.n207 585
R1884 B.n266 B.n265 585
R1885 B.n267 B.n206 585
R1886 B.n269 B.n268 585
R1887 B.n270 B.n205 585
R1888 B.n272 B.n271 585
R1889 B.n273 B.n204 585
R1890 B.n275 B.n274 585
R1891 B.n165 B.t7 562.816
R1892 B.n61 B.t2 562.816
R1893 B.n370 B.t10 562.816
R1894 B.n54 B.t5 562.816
R1895 B.n276 B.n275 521.33
R1896 B.n485 B.n132 521.33
R1897 B.n599 B.n94 521.33
R1898 B.n809 B.n808 521.33
R1899 B.n166 B.t8 514.138
R1900 B.n62 B.t1 514.138
R1901 B.n371 B.t11 514.136
R1902 B.n55 B.t4 514.136
R1903 B.n370 B.t9 424.875
R1904 B.n165 B.t6 424.875
R1905 B.n61 B.t0 424.875
R1906 B.n54 B.t3 424.875
R1907 B.n865 B.n864 256.663
R1908 B.n864 B.n863 235.042
R1909 B.n864 B.n2 235.042
R1910 B.n277 B.n276 163.367
R1911 B.n277 B.n202 163.367
R1912 B.n281 B.n202 163.367
R1913 B.n282 B.n281 163.367
R1914 B.n283 B.n282 163.367
R1915 B.n283 B.n200 163.367
R1916 B.n287 B.n200 163.367
R1917 B.n288 B.n287 163.367
R1918 B.n289 B.n288 163.367
R1919 B.n289 B.n198 163.367
R1920 B.n293 B.n198 163.367
R1921 B.n294 B.n293 163.367
R1922 B.n295 B.n294 163.367
R1923 B.n295 B.n196 163.367
R1924 B.n299 B.n196 163.367
R1925 B.n300 B.n299 163.367
R1926 B.n301 B.n300 163.367
R1927 B.n301 B.n194 163.367
R1928 B.n305 B.n194 163.367
R1929 B.n306 B.n305 163.367
R1930 B.n307 B.n306 163.367
R1931 B.n307 B.n192 163.367
R1932 B.n311 B.n192 163.367
R1933 B.n312 B.n311 163.367
R1934 B.n313 B.n312 163.367
R1935 B.n313 B.n190 163.367
R1936 B.n317 B.n190 163.367
R1937 B.n318 B.n317 163.367
R1938 B.n319 B.n318 163.367
R1939 B.n319 B.n188 163.367
R1940 B.n323 B.n188 163.367
R1941 B.n324 B.n323 163.367
R1942 B.n325 B.n324 163.367
R1943 B.n325 B.n186 163.367
R1944 B.n329 B.n186 163.367
R1945 B.n330 B.n329 163.367
R1946 B.n331 B.n330 163.367
R1947 B.n331 B.n184 163.367
R1948 B.n335 B.n184 163.367
R1949 B.n336 B.n335 163.367
R1950 B.n337 B.n336 163.367
R1951 B.n337 B.n182 163.367
R1952 B.n341 B.n182 163.367
R1953 B.n342 B.n341 163.367
R1954 B.n343 B.n342 163.367
R1955 B.n343 B.n180 163.367
R1956 B.n347 B.n180 163.367
R1957 B.n348 B.n347 163.367
R1958 B.n349 B.n348 163.367
R1959 B.n349 B.n178 163.367
R1960 B.n353 B.n178 163.367
R1961 B.n354 B.n353 163.367
R1962 B.n355 B.n354 163.367
R1963 B.n355 B.n176 163.367
R1964 B.n359 B.n176 163.367
R1965 B.n360 B.n359 163.367
R1966 B.n361 B.n360 163.367
R1967 B.n361 B.n174 163.367
R1968 B.n365 B.n174 163.367
R1969 B.n366 B.n365 163.367
R1970 B.n367 B.n366 163.367
R1971 B.n367 B.n172 163.367
R1972 B.n374 B.n172 163.367
R1973 B.n375 B.n374 163.367
R1974 B.n376 B.n375 163.367
R1975 B.n376 B.n170 163.367
R1976 B.n380 B.n170 163.367
R1977 B.n381 B.n380 163.367
R1978 B.n382 B.n381 163.367
R1979 B.n382 B.n168 163.367
R1980 B.n386 B.n168 163.367
R1981 B.n387 B.n386 163.367
R1982 B.n388 B.n387 163.367
R1983 B.n388 B.n164 163.367
R1984 B.n393 B.n164 163.367
R1985 B.n394 B.n393 163.367
R1986 B.n395 B.n394 163.367
R1987 B.n395 B.n162 163.367
R1988 B.n399 B.n162 163.367
R1989 B.n400 B.n399 163.367
R1990 B.n401 B.n400 163.367
R1991 B.n401 B.n160 163.367
R1992 B.n405 B.n160 163.367
R1993 B.n406 B.n405 163.367
R1994 B.n407 B.n406 163.367
R1995 B.n407 B.n158 163.367
R1996 B.n411 B.n158 163.367
R1997 B.n412 B.n411 163.367
R1998 B.n413 B.n412 163.367
R1999 B.n413 B.n156 163.367
R2000 B.n417 B.n156 163.367
R2001 B.n418 B.n417 163.367
R2002 B.n419 B.n418 163.367
R2003 B.n419 B.n154 163.367
R2004 B.n423 B.n154 163.367
R2005 B.n424 B.n423 163.367
R2006 B.n425 B.n424 163.367
R2007 B.n425 B.n152 163.367
R2008 B.n429 B.n152 163.367
R2009 B.n430 B.n429 163.367
R2010 B.n431 B.n430 163.367
R2011 B.n431 B.n150 163.367
R2012 B.n435 B.n150 163.367
R2013 B.n436 B.n435 163.367
R2014 B.n437 B.n436 163.367
R2015 B.n437 B.n148 163.367
R2016 B.n441 B.n148 163.367
R2017 B.n442 B.n441 163.367
R2018 B.n443 B.n442 163.367
R2019 B.n443 B.n146 163.367
R2020 B.n447 B.n146 163.367
R2021 B.n448 B.n447 163.367
R2022 B.n449 B.n448 163.367
R2023 B.n449 B.n144 163.367
R2024 B.n453 B.n144 163.367
R2025 B.n454 B.n453 163.367
R2026 B.n455 B.n454 163.367
R2027 B.n455 B.n142 163.367
R2028 B.n459 B.n142 163.367
R2029 B.n460 B.n459 163.367
R2030 B.n461 B.n460 163.367
R2031 B.n461 B.n140 163.367
R2032 B.n465 B.n140 163.367
R2033 B.n466 B.n465 163.367
R2034 B.n467 B.n466 163.367
R2035 B.n467 B.n138 163.367
R2036 B.n471 B.n138 163.367
R2037 B.n472 B.n471 163.367
R2038 B.n473 B.n472 163.367
R2039 B.n473 B.n136 163.367
R2040 B.n477 B.n136 163.367
R2041 B.n478 B.n477 163.367
R2042 B.n479 B.n478 163.367
R2043 B.n479 B.n134 163.367
R2044 B.n483 B.n134 163.367
R2045 B.n484 B.n483 163.367
R2046 B.n485 B.n484 163.367
R2047 B.n599 B.n598 163.367
R2048 B.n598 B.n597 163.367
R2049 B.n597 B.n96 163.367
R2050 B.n593 B.n96 163.367
R2051 B.n593 B.n592 163.367
R2052 B.n592 B.n591 163.367
R2053 B.n591 B.n98 163.367
R2054 B.n587 B.n98 163.367
R2055 B.n587 B.n586 163.367
R2056 B.n586 B.n585 163.367
R2057 B.n585 B.n100 163.367
R2058 B.n581 B.n100 163.367
R2059 B.n581 B.n580 163.367
R2060 B.n580 B.n579 163.367
R2061 B.n579 B.n102 163.367
R2062 B.n575 B.n102 163.367
R2063 B.n575 B.n574 163.367
R2064 B.n574 B.n573 163.367
R2065 B.n573 B.n104 163.367
R2066 B.n569 B.n104 163.367
R2067 B.n569 B.n568 163.367
R2068 B.n568 B.n567 163.367
R2069 B.n567 B.n106 163.367
R2070 B.n563 B.n106 163.367
R2071 B.n563 B.n562 163.367
R2072 B.n562 B.n561 163.367
R2073 B.n561 B.n108 163.367
R2074 B.n557 B.n108 163.367
R2075 B.n557 B.n556 163.367
R2076 B.n556 B.n555 163.367
R2077 B.n555 B.n110 163.367
R2078 B.n551 B.n110 163.367
R2079 B.n551 B.n550 163.367
R2080 B.n550 B.n549 163.367
R2081 B.n549 B.n112 163.367
R2082 B.n545 B.n112 163.367
R2083 B.n545 B.n544 163.367
R2084 B.n544 B.n543 163.367
R2085 B.n543 B.n114 163.367
R2086 B.n539 B.n114 163.367
R2087 B.n539 B.n538 163.367
R2088 B.n538 B.n537 163.367
R2089 B.n537 B.n116 163.367
R2090 B.n533 B.n116 163.367
R2091 B.n533 B.n532 163.367
R2092 B.n532 B.n531 163.367
R2093 B.n531 B.n118 163.367
R2094 B.n527 B.n118 163.367
R2095 B.n527 B.n526 163.367
R2096 B.n526 B.n525 163.367
R2097 B.n525 B.n120 163.367
R2098 B.n521 B.n120 163.367
R2099 B.n521 B.n520 163.367
R2100 B.n520 B.n519 163.367
R2101 B.n519 B.n122 163.367
R2102 B.n515 B.n122 163.367
R2103 B.n515 B.n514 163.367
R2104 B.n514 B.n513 163.367
R2105 B.n513 B.n124 163.367
R2106 B.n509 B.n124 163.367
R2107 B.n509 B.n508 163.367
R2108 B.n508 B.n507 163.367
R2109 B.n507 B.n126 163.367
R2110 B.n503 B.n126 163.367
R2111 B.n503 B.n502 163.367
R2112 B.n502 B.n501 163.367
R2113 B.n501 B.n128 163.367
R2114 B.n497 B.n128 163.367
R2115 B.n497 B.n496 163.367
R2116 B.n496 B.n495 163.367
R2117 B.n495 B.n130 163.367
R2118 B.n491 B.n130 163.367
R2119 B.n491 B.n490 163.367
R2120 B.n490 B.n489 163.367
R2121 B.n489 B.n132 163.367
R2122 B.n808 B.n21 163.367
R2123 B.n804 B.n21 163.367
R2124 B.n804 B.n803 163.367
R2125 B.n803 B.n802 163.367
R2126 B.n802 B.n23 163.367
R2127 B.n798 B.n23 163.367
R2128 B.n798 B.n797 163.367
R2129 B.n797 B.n796 163.367
R2130 B.n796 B.n25 163.367
R2131 B.n792 B.n25 163.367
R2132 B.n792 B.n791 163.367
R2133 B.n791 B.n790 163.367
R2134 B.n790 B.n27 163.367
R2135 B.n786 B.n27 163.367
R2136 B.n786 B.n785 163.367
R2137 B.n785 B.n784 163.367
R2138 B.n784 B.n29 163.367
R2139 B.n780 B.n29 163.367
R2140 B.n780 B.n779 163.367
R2141 B.n779 B.n778 163.367
R2142 B.n778 B.n31 163.367
R2143 B.n774 B.n31 163.367
R2144 B.n774 B.n773 163.367
R2145 B.n773 B.n772 163.367
R2146 B.n772 B.n33 163.367
R2147 B.n768 B.n33 163.367
R2148 B.n768 B.n767 163.367
R2149 B.n767 B.n766 163.367
R2150 B.n766 B.n35 163.367
R2151 B.n762 B.n35 163.367
R2152 B.n762 B.n761 163.367
R2153 B.n761 B.n760 163.367
R2154 B.n760 B.n37 163.367
R2155 B.n756 B.n37 163.367
R2156 B.n756 B.n755 163.367
R2157 B.n755 B.n754 163.367
R2158 B.n754 B.n39 163.367
R2159 B.n750 B.n39 163.367
R2160 B.n750 B.n749 163.367
R2161 B.n749 B.n748 163.367
R2162 B.n748 B.n41 163.367
R2163 B.n744 B.n41 163.367
R2164 B.n744 B.n743 163.367
R2165 B.n743 B.n742 163.367
R2166 B.n742 B.n43 163.367
R2167 B.n738 B.n43 163.367
R2168 B.n738 B.n737 163.367
R2169 B.n737 B.n736 163.367
R2170 B.n736 B.n45 163.367
R2171 B.n732 B.n45 163.367
R2172 B.n732 B.n731 163.367
R2173 B.n731 B.n730 163.367
R2174 B.n730 B.n47 163.367
R2175 B.n726 B.n47 163.367
R2176 B.n726 B.n725 163.367
R2177 B.n725 B.n724 163.367
R2178 B.n724 B.n49 163.367
R2179 B.n720 B.n49 163.367
R2180 B.n720 B.n719 163.367
R2181 B.n719 B.n718 163.367
R2182 B.n718 B.n51 163.367
R2183 B.n714 B.n51 163.367
R2184 B.n714 B.n713 163.367
R2185 B.n713 B.n712 163.367
R2186 B.n712 B.n53 163.367
R2187 B.n708 B.n53 163.367
R2188 B.n708 B.n707 163.367
R2189 B.n707 B.n706 163.367
R2190 B.n706 B.n58 163.367
R2191 B.n702 B.n58 163.367
R2192 B.n702 B.n701 163.367
R2193 B.n701 B.n700 163.367
R2194 B.n700 B.n60 163.367
R2195 B.n695 B.n60 163.367
R2196 B.n695 B.n694 163.367
R2197 B.n694 B.n693 163.367
R2198 B.n693 B.n64 163.367
R2199 B.n689 B.n64 163.367
R2200 B.n689 B.n688 163.367
R2201 B.n688 B.n687 163.367
R2202 B.n687 B.n66 163.367
R2203 B.n683 B.n66 163.367
R2204 B.n683 B.n682 163.367
R2205 B.n682 B.n681 163.367
R2206 B.n681 B.n68 163.367
R2207 B.n677 B.n68 163.367
R2208 B.n677 B.n676 163.367
R2209 B.n676 B.n675 163.367
R2210 B.n675 B.n70 163.367
R2211 B.n671 B.n70 163.367
R2212 B.n671 B.n670 163.367
R2213 B.n670 B.n669 163.367
R2214 B.n669 B.n72 163.367
R2215 B.n665 B.n72 163.367
R2216 B.n665 B.n664 163.367
R2217 B.n664 B.n663 163.367
R2218 B.n663 B.n74 163.367
R2219 B.n659 B.n74 163.367
R2220 B.n659 B.n658 163.367
R2221 B.n658 B.n657 163.367
R2222 B.n657 B.n76 163.367
R2223 B.n653 B.n76 163.367
R2224 B.n653 B.n652 163.367
R2225 B.n652 B.n651 163.367
R2226 B.n651 B.n78 163.367
R2227 B.n647 B.n78 163.367
R2228 B.n647 B.n646 163.367
R2229 B.n646 B.n645 163.367
R2230 B.n645 B.n80 163.367
R2231 B.n641 B.n80 163.367
R2232 B.n641 B.n640 163.367
R2233 B.n640 B.n639 163.367
R2234 B.n639 B.n82 163.367
R2235 B.n635 B.n82 163.367
R2236 B.n635 B.n634 163.367
R2237 B.n634 B.n633 163.367
R2238 B.n633 B.n84 163.367
R2239 B.n629 B.n84 163.367
R2240 B.n629 B.n628 163.367
R2241 B.n628 B.n627 163.367
R2242 B.n627 B.n86 163.367
R2243 B.n623 B.n86 163.367
R2244 B.n623 B.n622 163.367
R2245 B.n622 B.n621 163.367
R2246 B.n621 B.n88 163.367
R2247 B.n617 B.n88 163.367
R2248 B.n617 B.n616 163.367
R2249 B.n616 B.n615 163.367
R2250 B.n615 B.n90 163.367
R2251 B.n611 B.n90 163.367
R2252 B.n611 B.n610 163.367
R2253 B.n610 B.n609 163.367
R2254 B.n609 B.n92 163.367
R2255 B.n605 B.n92 163.367
R2256 B.n605 B.n604 163.367
R2257 B.n604 B.n603 163.367
R2258 B.n603 B.n94 163.367
R2259 B.n810 B.n809 163.367
R2260 B.n810 B.n19 163.367
R2261 B.n814 B.n19 163.367
R2262 B.n815 B.n814 163.367
R2263 B.n816 B.n815 163.367
R2264 B.n816 B.n17 163.367
R2265 B.n820 B.n17 163.367
R2266 B.n821 B.n820 163.367
R2267 B.n822 B.n821 163.367
R2268 B.n822 B.n15 163.367
R2269 B.n826 B.n15 163.367
R2270 B.n827 B.n826 163.367
R2271 B.n828 B.n827 163.367
R2272 B.n828 B.n13 163.367
R2273 B.n832 B.n13 163.367
R2274 B.n833 B.n832 163.367
R2275 B.n834 B.n833 163.367
R2276 B.n834 B.n11 163.367
R2277 B.n838 B.n11 163.367
R2278 B.n839 B.n838 163.367
R2279 B.n840 B.n839 163.367
R2280 B.n840 B.n9 163.367
R2281 B.n844 B.n9 163.367
R2282 B.n845 B.n844 163.367
R2283 B.n846 B.n845 163.367
R2284 B.n846 B.n7 163.367
R2285 B.n850 B.n7 163.367
R2286 B.n851 B.n850 163.367
R2287 B.n852 B.n851 163.367
R2288 B.n852 B.n5 163.367
R2289 B.n856 B.n5 163.367
R2290 B.n857 B.n856 163.367
R2291 B.n858 B.n857 163.367
R2292 B.n858 B.n3 163.367
R2293 B.n862 B.n3 163.367
R2294 B.n863 B.n862 163.367
R2295 B.n222 B.n2 163.367
R2296 B.n223 B.n222 163.367
R2297 B.n223 B.n220 163.367
R2298 B.n227 B.n220 163.367
R2299 B.n228 B.n227 163.367
R2300 B.n229 B.n228 163.367
R2301 B.n229 B.n218 163.367
R2302 B.n233 B.n218 163.367
R2303 B.n234 B.n233 163.367
R2304 B.n235 B.n234 163.367
R2305 B.n235 B.n216 163.367
R2306 B.n239 B.n216 163.367
R2307 B.n240 B.n239 163.367
R2308 B.n241 B.n240 163.367
R2309 B.n241 B.n214 163.367
R2310 B.n245 B.n214 163.367
R2311 B.n246 B.n245 163.367
R2312 B.n247 B.n246 163.367
R2313 B.n247 B.n212 163.367
R2314 B.n251 B.n212 163.367
R2315 B.n252 B.n251 163.367
R2316 B.n253 B.n252 163.367
R2317 B.n253 B.n210 163.367
R2318 B.n257 B.n210 163.367
R2319 B.n258 B.n257 163.367
R2320 B.n259 B.n258 163.367
R2321 B.n259 B.n208 163.367
R2322 B.n263 B.n208 163.367
R2323 B.n264 B.n263 163.367
R2324 B.n265 B.n264 163.367
R2325 B.n265 B.n206 163.367
R2326 B.n269 B.n206 163.367
R2327 B.n270 B.n269 163.367
R2328 B.n271 B.n270 163.367
R2329 B.n271 B.n204 163.367
R2330 B.n275 B.n204 163.367
R2331 B.n372 B.n371 59.5399
R2332 B.n390 B.n166 59.5399
R2333 B.n697 B.n62 59.5399
R2334 B.n56 B.n55 59.5399
R2335 B.n371 B.n370 48.6793
R2336 B.n166 B.n165 48.6793
R2337 B.n62 B.n61 48.6793
R2338 B.n55 B.n54 48.6793
R2339 B.n807 B.n20 33.8737
R2340 B.n601 B.n600 33.8737
R2341 B.n487 B.n486 33.8737
R2342 B.n274 B.n203 33.8737
R2343 B B.n865 18.0485
R2344 B.n811 B.n20 10.6151
R2345 B.n812 B.n811 10.6151
R2346 B.n813 B.n812 10.6151
R2347 B.n813 B.n18 10.6151
R2348 B.n817 B.n18 10.6151
R2349 B.n818 B.n817 10.6151
R2350 B.n819 B.n818 10.6151
R2351 B.n819 B.n16 10.6151
R2352 B.n823 B.n16 10.6151
R2353 B.n824 B.n823 10.6151
R2354 B.n825 B.n824 10.6151
R2355 B.n825 B.n14 10.6151
R2356 B.n829 B.n14 10.6151
R2357 B.n830 B.n829 10.6151
R2358 B.n831 B.n830 10.6151
R2359 B.n831 B.n12 10.6151
R2360 B.n835 B.n12 10.6151
R2361 B.n836 B.n835 10.6151
R2362 B.n837 B.n836 10.6151
R2363 B.n837 B.n10 10.6151
R2364 B.n841 B.n10 10.6151
R2365 B.n842 B.n841 10.6151
R2366 B.n843 B.n842 10.6151
R2367 B.n843 B.n8 10.6151
R2368 B.n847 B.n8 10.6151
R2369 B.n848 B.n847 10.6151
R2370 B.n849 B.n848 10.6151
R2371 B.n849 B.n6 10.6151
R2372 B.n853 B.n6 10.6151
R2373 B.n854 B.n853 10.6151
R2374 B.n855 B.n854 10.6151
R2375 B.n855 B.n4 10.6151
R2376 B.n859 B.n4 10.6151
R2377 B.n860 B.n859 10.6151
R2378 B.n861 B.n860 10.6151
R2379 B.n861 B.n0 10.6151
R2380 B.n807 B.n806 10.6151
R2381 B.n806 B.n805 10.6151
R2382 B.n805 B.n22 10.6151
R2383 B.n801 B.n22 10.6151
R2384 B.n801 B.n800 10.6151
R2385 B.n800 B.n799 10.6151
R2386 B.n799 B.n24 10.6151
R2387 B.n795 B.n24 10.6151
R2388 B.n795 B.n794 10.6151
R2389 B.n794 B.n793 10.6151
R2390 B.n793 B.n26 10.6151
R2391 B.n789 B.n26 10.6151
R2392 B.n789 B.n788 10.6151
R2393 B.n788 B.n787 10.6151
R2394 B.n787 B.n28 10.6151
R2395 B.n783 B.n28 10.6151
R2396 B.n783 B.n782 10.6151
R2397 B.n782 B.n781 10.6151
R2398 B.n781 B.n30 10.6151
R2399 B.n777 B.n30 10.6151
R2400 B.n777 B.n776 10.6151
R2401 B.n776 B.n775 10.6151
R2402 B.n775 B.n32 10.6151
R2403 B.n771 B.n32 10.6151
R2404 B.n771 B.n770 10.6151
R2405 B.n770 B.n769 10.6151
R2406 B.n769 B.n34 10.6151
R2407 B.n765 B.n34 10.6151
R2408 B.n765 B.n764 10.6151
R2409 B.n764 B.n763 10.6151
R2410 B.n763 B.n36 10.6151
R2411 B.n759 B.n36 10.6151
R2412 B.n759 B.n758 10.6151
R2413 B.n758 B.n757 10.6151
R2414 B.n757 B.n38 10.6151
R2415 B.n753 B.n38 10.6151
R2416 B.n753 B.n752 10.6151
R2417 B.n752 B.n751 10.6151
R2418 B.n751 B.n40 10.6151
R2419 B.n747 B.n40 10.6151
R2420 B.n747 B.n746 10.6151
R2421 B.n746 B.n745 10.6151
R2422 B.n745 B.n42 10.6151
R2423 B.n741 B.n42 10.6151
R2424 B.n741 B.n740 10.6151
R2425 B.n740 B.n739 10.6151
R2426 B.n739 B.n44 10.6151
R2427 B.n735 B.n44 10.6151
R2428 B.n735 B.n734 10.6151
R2429 B.n734 B.n733 10.6151
R2430 B.n733 B.n46 10.6151
R2431 B.n729 B.n46 10.6151
R2432 B.n729 B.n728 10.6151
R2433 B.n728 B.n727 10.6151
R2434 B.n727 B.n48 10.6151
R2435 B.n723 B.n48 10.6151
R2436 B.n723 B.n722 10.6151
R2437 B.n722 B.n721 10.6151
R2438 B.n721 B.n50 10.6151
R2439 B.n717 B.n50 10.6151
R2440 B.n717 B.n716 10.6151
R2441 B.n716 B.n715 10.6151
R2442 B.n715 B.n52 10.6151
R2443 B.n711 B.n710 10.6151
R2444 B.n710 B.n709 10.6151
R2445 B.n709 B.n57 10.6151
R2446 B.n705 B.n57 10.6151
R2447 B.n705 B.n704 10.6151
R2448 B.n704 B.n703 10.6151
R2449 B.n703 B.n59 10.6151
R2450 B.n699 B.n59 10.6151
R2451 B.n699 B.n698 10.6151
R2452 B.n696 B.n63 10.6151
R2453 B.n692 B.n63 10.6151
R2454 B.n692 B.n691 10.6151
R2455 B.n691 B.n690 10.6151
R2456 B.n690 B.n65 10.6151
R2457 B.n686 B.n65 10.6151
R2458 B.n686 B.n685 10.6151
R2459 B.n685 B.n684 10.6151
R2460 B.n684 B.n67 10.6151
R2461 B.n680 B.n67 10.6151
R2462 B.n680 B.n679 10.6151
R2463 B.n679 B.n678 10.6151
R2464 B.n678 B.n69 10.6151
R2465 B.n674 B.n69 10.6151
R2466 B.n674 B.n673 10.6151
R2467 B.n673 B.n672 10.6151
R2468 B.n672 B.n71 10.6151
R2469 B.n668 B.n71 10.6151
R2470 B.n668 B.n667 10.6151
R2471 B.n667 B.n666 10.6151
R2472 B.n666 B.n73 10.6151
R2473 B.n662 B.n73 10.6151
R2474 B.n662 B.n661 10.6151
R2475 B.n661 B.n660 10.6151
R2476 B.n660 B.n75 10.6151
R2477 B.n656 B.n75 10.6151
R2478 B.n656 B.n655 10.6151
R2479 B.n655 B.n654 10.6151
R2480 B.n654 B.n77 10.6151
R2481 B.n650 B.n77 10.6151
R2482 B.n650 B.n649 10.6151
R2483 B.n649 B.n648 10.6151
R2484 B.n648 B.n79 10.6151
R2485 B.n644 B.n79 10.6151
R2486 B.n644 B.n643 10.6151
R2487 B.n643 B.n642 10.6151
R2488 B.n642 B.n81 10.6151
R2489 B.n638 B.n81 10.6151
R2490 B.n638 B.n637 10.6151
R2491 B.n637 B.n636 10.6151
R2492 B.n636 B.n83 10.6151
R2493 B.n632 B.n83 10.6151
R2494 B.n632 B.n631 10.6151
R2495 B.n631 B.n630 10.6151
R2496 B.n630 B.n85 10.6151
R2497 B.n626 B.n85 10.6151
R2498 B.n626 B.n625 10.6151
R2499 B.n625 B.n624 10.6151
R2500 B.n624 B.n87 10.6151
R2501 B.n620 B.n87 10.6151
R2502 B.n620 B.n619 10.6151
R2503 B.n619 B.n618 10.6151
R2504 B.n618 B.n89 10.6151
R2505 B.n614 B.n89 10.6151
R2506 B.n614 B.n613 10.6151
R2507 B.n613 B.n612 10.6151
R2508 B.n612 B.n91 10.6151
R2509 B.n608 B.n91 10.6151
R2510 B.n608 B.n607 10.6151
R2511 B.n607 B.n606 10.6151
R2512 B.n606 B.n93 10.6151
R2513 B.n602 B.n93 10.6151
R2514 B.n602 B.n601 10.6151
R2515 B.n600 B.n95 10.6151
R2516 B.n596 B.n95 10.6151
R2517 B.n596 B.n595 10.6151
R2518 B.n595 B.n594 10.6151
R2519 B.n594 B.n97 10.6151
R2520 B.n590 B.n97 10.6151
R2521 B.n590 B.n589 10.6151
R2522 B.n589 B.n588 10.6151
R2523 B.n588 B.n99 10.6151
R2524 B.n584 B.n99 10.6151
R2525 B.n584 B.n583 10.6151
R2526 B.n583 B.n582 10.6151
R2527 B.n582 B.n101 10.6151
R2528 B.n578 B.n101 10.6151
R2529 B.n578 B.n577 10.6151
R2530 B.n577 B.n576 10.6151
R2531 B.n576 B.n103 10.6151
R2532 B.n572 B.n103 10.6151
R2533 B.n572 B.n571 10.6151
R2534 B.n571 B.n570 10.6151
R2535 B.n570 B.n105 10.6151
R2536 B.n566 B.n105 10.6151
R2537 B.n566 B.n565 10.6151
R2538 B.n565 B.n564 10.6151
R2539 B.n564 B.n107 10.6151
R2540 B.n560 B.n107 10.6151
R2541 B.n560 B.n559 10.6151
R2542 B.n559 B.n558 10.6151
R2543 B.n558 B.n109 10.6151
R2544 B.n554 B.n109 10.6151
R2545 B.n554 B.n553 10.6151
R2546 B.n553 B.n552 10.6151
R2547 B.n552 B.n111 10.6151
R2548 B.n548 B.n111 10.6151
R2549 B.n548 B.n547 10.6151
R2550 B.n547 B.n546 10.6151
R2551 B.n546 B.n113 10.6151
R2552 B.n542 B.n113 10.6151
R2553 B.n542 B.n541 10.6151
R2554 B.n541 B.n540 10.6151
R2555 B.n540 B.n115 10.6151
R2556 B.n536 B.n115 10.6151
R2557 B.n536 B.n535 10.6151
R2558 B.n535 B.n534 10.6151
R2559 B.n534 B.n117 10.6151
R2560 B.n530 B.n117 10.6151
R2561 B.n530 B.n529 10.6151
R2562 B.n529 B.n528 10.6151
R2563 B.n528 B.n119 10.6151
R2564 B.n524 B.n119 10.6151
R2565 B.n524 B.n523 10.6151
R2566 B.n523 B.n522 10.6151
R2567 B.n522 B.n121 10.6151
R2568 B.n518 B.n121 10.6151
R2569 B.n518 B.n517 10.6151
R2570 B.n517 B.n516 10.6151
R2571 B.n516 B.n123 10.6151
R2572 B.n512 B.n123 10.6151
R2573 B.n512 B.n511 10.6151
R2574 B.n511 B.n510 10.6151
R2575 B.n510 B.n125 10.6151
R2576 B.n506 B.n125 10.6151
R2577 B.n506 B.n505 10.6151
R2578 B.n505 B.n504 10.6151
R2579 B.n504 B.n127 10.6151
R2580 B.n500 B.n127 10.6151
R2581 B.n500 B.n499 10.6151
R2582 B.n499 B.n498 10.6151
R2583 B.n498 B.n129 10.6151
R2584 B.n494 B.n129 10.6151
R2585 B.n494 B.n493 10.6151
R2586 B.n493 B.n492 10.6151
R2587 B.n492 B.n131 10.6151
R2588 B.n488 B.n131 10.6151
R2589 B.n488 B.n487 10.6151
R2590 B.n221 B.n1 10.6151
R2591 B.n224 B.n221 10.6151
R2592 B.n225 B.n224 10.6151
R2593 B.n226 B.n225 10.6151
R2594 B.n226 B.n219 10.6151
R2595 B.n230 B.n219 10.6151
R2596 B.n231 B.n230 10.6151
R2597 B.n232 B.n231 10.6151
R2598 B.n232 B.n217 10.6151
R2599 B.n236 B.n217 10.6151
R2600 B.n237 B.n236 10.6151
R2601 B.n238 B.n237 10.6151
R2602 B.n238 B.n215 10.6151
R2603 B.n242 B.n215 10.6151
R2604 B.n243 B.n242 10.6151
R2605 B.n244 B.n243 10.6151
R2606 B.n244 B.n213 10.6151
R2607 B.n248 B.n213 10.6151
R2608 B.n249 B.n248 10.6151
R2609 B.n250 B.n249 10.6151
R2610 B.n250 B.n211 10.6151
R2611 B.n254 B.n211 10.6151
R2612 B.n255 B.n254 10.6151
R2613 B.n256 B.n255 10.6151
R2614 B.n256 B.n209 10.6151
R2615 B.n260 B.n209 10.6151
R2616 B.n261 B.n260 10.6151
R2617 B.n262 B.n261 10.6151
R2618 B.n262 B.n207 10.6151
R2619 B.n266 B.n207 10.6151
R2620 B.n267 B.n266 10.6151
R2621 B.n268 B.n267 10.6151
R2622 B.n268 B.n205 10.6151
R2623 B.n272 B.n205 10.6151
R2624 B.n273 B.n272 10.6151
R2625 B.n274 B.n273 10.6151
R2626 B.n278 B.n203 10.6151
R2627 B.n279 B.n278 10.6151
R2628 B.n280 B.n279 10.6151
R2629 B.n280 B.n201 10.6151
R2630 B.n284 B.n201 10.6151
R2631 B.n285 B.n284 10.6151
R2632 B.n286 B.n285 10.6151
R2633 B.n286 B.n199 10.6151
R2634 B.n290 B.n199 10.6151
R2635 B.n291 B.n290 10.6151
R2636 B.n292 B.n291 10.6151
R2637 B.n292 B.n197 10.6151
R2638 B.n296 B.n197 10.6151
R2639 B.n297 B.n296 10.6151
R2640 B.n298 B.n297 10.6151
R2641 B.n298 B.n195 10.6151
R2642 B.n302 B.n195 10.6151
R2643 B.n303 B.n302 10.6151
R2644 B.n304 B.n303 10.6151
R2645 B.n304 B.n193 10.6151
R2646 B.n308 B.n193 10.6151
R2647 B.n309 B.n308 10.6151
R2648 B.n310 B.n309 10.6151
R2649 B.n310 B.n191 10.6151
R2650 B.n314 B.n191 10.6151
R2651 B.n315 B.n314 10.6151
R2652 B.n316 B.n315 10.6151
R2653 B.n316 B.n189 10.6151
R2654 B.n320 B.n189 10.6151
R2655 B.n321 B.n320 10.6151
R2656 B.n322 B.n321 10.6151
R2657 B.n322 B.n187 10.6151
R2658 B.n326 B.n187 10.6151
R2659 B.n327 B.n326 10.6151
R2660 B.n328 B.n327 10.6151
R2661 B.n328 B.n185 10.6151
R2662 B.n332 B.n185 10.6151
R2663 B.n333 B.n332 10.6151
R2664 B.n334 B.n333 10.6151
R2665 B.n334 B.n183 10.6151
R2666 B.n338 B.n183 10.6151
R2667 B.n339 B.n338 10.6151
R2668 B.n340 B.n339 10.6151
R2669 B.n340 B.n181 10.6151
R2670 B.n344 B.n181 10.6151
R2671 B.n345 B.n344 10.6151
R2672 B.n346 B.n345 10.6151
R2673 B.n346 B.n179 10.6151
R2674 B.n350 B.n179 10.6151
R2675 B.n351 B.n350 10.6151
R2676 B.n352 B.n351 10.6151
R2677 B.n352 B.n177 10.6151
R2678 B.n356 B.n177 10.6151
R2679 B.n357 B.n356 10.6151
R2680 B.n358 B.n357 10.6151
R2681 B.n358 B.n175 10.6151
R2682 B.n362 B.n175 10.6151
R2683 B.n363 B.n362 10.6151
R2684 B.n364 B.n363 10.6151
R2685 B.n364 B.n173 10.6151
R2686 B.n368 B.n173 10.6151
R2687 B.n369 B.n368 10.6151
R2688 B.n373 B.n369 10.6151
R2689 B.n377 B.n171 10.6151
R2690 B.n378 B.n377 10.6151
R2691 B.n379 B.n378 10.6151
R2692 B.n379 B.n169 10.6151
R2693 B.n383 B.n169 10.6151
R2694 B.n384 B.n383 10.6151
R2695 B.n385 B.n384 10.6151
R2696 B.n385 B.n167 10.6151
R2697 B.n389 B.n167 10.6151
R2698 B.n392 B.n391 10.6151
R2699 B.n392 B.n163 10.6151
R2700 B.n396 B.n163 10.6151
R2701 B.n397 B.n396 10.6151
R2702 B.n398 B.n397 10.6151
R2703 B.n398 B.n161 10.6151
R2704 B.n402 B.n161 10.6151
R2705 B.n403 B.n402 10.6151
R2706 B.n404 B.n403 10.6151
R2707 B.n404 B.n159 10.6151
R2708 B.n408 B.n159 10.6151
R2709 B.n409 B.n408 10.6151
R2710 B.n410 B.n409 10.6151
R2711 B.n410 B.n157 10.6151
R2712 B.n414 B.n157 10.6151
R2713 B.n415 B.n414 10.6151
R2714 B.n416 B.n415 10.6151
R2715 B.n416 B.n155 10.6151
R2716 B.n420 B.n155 10.6151
R2717 B.n421 B.n420 10.6151
R2718 B.n422 B.n421 10.6151
R2719 B.n422 B.n153 10.6151
R2720 B.n426 B.n153 10.6151
R2721 B.n427 B.n426 10.6151
R2722 B.n428 B.n427 10.6151
R2723 B.n428 B.n151 10.6151
R2724 B.n432 B.n151 10.6151
R2725 B.n433 B.n432 10.6151
R2726 B.n434 B.n433 10.6151
R2727 B.n434 B.n149 10.6151
R2728 B.n438 B.n149 10.6151
R2729 B.n439 B.n438 10.6151
R2730 B.n440 B.n439 10.6151
R2731 B.n440 B.n147 10.6151
R2732 B.n444 B.n147 10.6151
R2733 B.n445 B.n444 10.6151
R2734 B.n446 B.n445 10.6151
R2735 B.n446 B.n145 10.6151
R2736 B.n450 B.n145 10.6151
R2737 B.n451 B.n450 10.6151
R2738 B.n452 B.n451 10.6151
R2739 B.n452 B.n143 10.6151
R2740 B.n456 B.n143 10.6151
R2741 B.n457 B.n456 10.6151
R2742 B.n458 B.n457 10.6151
R2743 B.n458 B.n141 10.6151
R2744 B.n462 B.n141 10.6151
R2745 B.n463 B.n462 10.6151
R2746 B.n464 B.n463 10.6151
R2747 B.n464 B.n139 10.6151
R2748 B.n468 B.n139 10.6151
R2749 B.n469 B.n468 10.6151
R2750 B.n470 B.n469 10.6151
R2751 B.n470 B.n137 10.6151
R2752 B.n474 B.n137 10.6151
R2753 B.n475 B.n474 10.6151
R2754 B.n476 B.n475 10.6151
R2755 B.n476 B.n135 10.6151
R2756 B.n480 B.n135 10.6151
R2757 B.n481 B.n480 10.6151
R2758 B.n482 B.n481 10.6151
R2759 B.n482 B.n133 10.6151
R2760 B.n486 B.n133 10.6151
R2761 B.n56 B.n52 9.36635
R2762 B.n697 B.n696 9.36635
R2763 B.n373 B.n372 9.36635
R2764 B.n391 B.n390 9.36635
R2765 B.n865 B.n0 8.11757
R2766 B.n865 B.n1 8.11757
R2767 B.n711 B.n56 1.24928
R2768 B.n698 B.n697 1.24928
R2769 B.n372 B.n171 1.24928
R2770 B.n390 B.n389 1.24928
C0 w_n2978_n4904# VDD2 2.79596f
C1 VP VDD2 0.423548f
C2 w_n2978_n4904# VP 6.07493f
C3 VN VDD2 10.4005f
C4 w_n2978_n4904# VN 5.69109f
C5 VTAIL VDD1 10.6901f
C6 VDD1 B 2.58205f
C7 VP VN 7.939899f
C8 VTAIL B 5.18116f
C9 VDD1 VDD2 1.24299f
C10 VDD1 w_n2978_n4904# 2.72427f
C11 VDD1 VP 10.6689f
C12 VTAIL VDD2 10.735499f
C13 B VDD2 2.64607f
C14 VTAIL w_n2978_n4904# 4.02529f
C15 w_n2978_n4904# B 11.2488f
C16 VDD1 VN 0.150283f
C17 VTAIL VP 10.1449f
C18 B VP 1.81087f
C19 VTAIL VN 10.1305f
C20 B VN 1.17212f
C21 VDD2 VSUBS 2.032634f
C22 VDD1 VSUBS 1.908061f
C23 VTAIL VSUBS 1.393761f
C24 VN VSUBS 5.81783f
C25 VP VSUBS 2.89023f
C26 B VSUBS 4.870359f
C27 w_n2978_n4904# VSUBS 0.178358p
C28 B.n0 VSUBS 0.006413f
C29 B.n1 VSUBS 0.006413f
C30 B.n2 VSUBS 0.009484f
C31 B.n3 VSUBS 0.007268f
C32 B.n4 VSUBS 0.007268f
C33 B.n5 VSUBS 0.007268f
C34 B.n6 VSUBS 0.007268f
C35 B.n7 VSUBS 0.007268f
C36 B.n8 VSUBS 0.007268f
C37 B.n9 VSUBS 0.007268f
C38 B.n10 VSUBS 0.007268f
C39 B.n11 VSUBS 0.007268f
C40 B.n12 VSUBS 0.007268f
C41 B.n13 VSUBS 0.007268f
C42 B.n14 VSUBS 0.007268f
C43 B.n15 VSUBS 0.007268f
C44 B.n16 VSUBS 0.007268f
C45 B.n17 VSUBS 0.007268f
C46 B.n18 VSUBS 0.007268f
C47 B.n19 VSUBS 0.007268f
C48 B.n20 VSUBS 0.016926f
C49 B.n21 VSUBS 0.007268f
C50 B.n22 VSUBS 0.007268f
C51 B.n23 VSUBS 0.007268f
C52 B.n24 VSUBS 0.007268f
C53 B.n25 VSUBS 0.007268f
C54 B.n26 VSUBS 0.007268f
C55 B.n27 VSUBS 0.007268f
C56 B.n28 VSUBS 0.007268f
C57 B.n29 VSUBS 0.007268f
C58 B.n30 VSUBS 0.007268f
C59 B.n31 VSUBS 0.007268f
C60 B.n32 VSUBS 0.007268f
C61 B.n33 VSUBS 0.007268f
C62 B.n34 VSUBS 0.007268f
C63 B.n35 VSUBS 0.007268f
C64 B.n36 VSUBS 0.007268f
C65 B.n37 VSUBS 0.007268f
C66 B.n38 VSUBS 0.007268f
C67 B.n39 VSUBS 0.007268f
C68 B.n40 VSUBS 0.007268f
C69 B.n41 VSUBS 0.007268f
C70 B.n42 VSUBS 0.007268f
C71 B.n43 VSUBS 0.007268f
C72 B.n44 VSUBS 0.007268f
C73 B.n45 VSUBS 0.007268f
C74 B.n46 VSUBS 0.007268f
C75 B.n47 VSUBS 0.007268f
C76 B.n48 VSUBS 0.007268f
C77 B.n49 VSUBS 0.007268f
C78 B.n50 VSUBS 0.007268f
C79 B.n51 VSUBS 0.007268f
C80 B.n52 VSUBS 0.00684f
C81 B.n53 VSUBS 0.007268f
C82 B.t4 VSUBS 0.407171f
C83 B.t5 VSUBS 0.437399f
C84 B.t3 VSUBS 1.9376f
C85 B.n54 VSUBS 0.645634f
C86 B.n55 VSUBS 0.359858f
C87 B.n56 VSUBS 0.016838f
C88 B.n57 VSUBS 0.007268f
C89 B.n58 VSUBS 0.007268f
C90 B.n59 VSUBS 0.007268f
C91 B.n60 VSUBS 0.007268f
C92 B.t1 VSUBS 0.407174f
C93 B.t2 VSUBS 0.437402f
C94 B.t0 VSUBS 1.9376f
C95 B.n61 VSUBS 0.645631f
C96 B.n62 VSUBS 0.359854f
C97 B.n63 VSUBS 0.007268f
C98 B.n64 VSUBS 0.007268f
C99 B.n65 VSUBS 0.007268f
C100 B.n66 VSUBS 0.007268f
C101 B.n67 VSUBS 0.007268f
C102 B.n68 VSUBS 0.007268f
C103 B.n69 VSUBS 0.007268f
C104 B.n70 VSUBS 0.007268f
C105 B.n71 VSUBS 0.007268f
C106 B.n72 VSUBS 0.007268f
C107 B.n73 VSUBS 0.007268f
C108 B.n74 VSUBS 0.007268f
C109 B.n75 VSUBS 0.007268f
C110 B.n76 VSUBS 0.007268f
C111 B.n77 VSUBS 0.007268f
C112 B.n78 VSUBS 0.007268f
C113 B.n79 VSUBS 0.007268f
C114 B.n80 VSUBS 0.007268f
C115 B.n81 VSUBS 0.007268f
C116 B.n82 VSUBS 0.007268f
C117 B.n83 VSUBS 0.007268f
C118 B.n84 VSUBS 0.007268f
C119 B.n85 VSUBS 0.007268f
C120 B.n86 VSUBS 0.007268f
C121 B.n87 VSUBS 0.007268f
C122 B.n88 VSUBS 0.007268f
C123 B.n89 VSUBS 0.007268f
C124 B.n90 VSUBS 0.007268f
C125 B.n91 VSUBS 0.007268f
C126 B.n92 VSUBS 0.007268f
C127 B.n93 VSUBS 0.007268f
C128 B.n94 VSUBS 0.017916f
C129 B.n95 VSUBS 0.007268f
C130 B.n96 VSUBS 0.007268f
C131 B.n97 VSUBS 0.007268f
C132 B.n98 VSUBS 0.007268f
C133 B.n99 VSUBS 0.007268f
C134 B.n100 VSUBS 0.007268f
C135 B.n101 VSUBS 0.007268f
C136 B.n102 VSUBS 0.007268f
C137 B.n103 VSUBS 0.007268f
C138 B.n104 VSUBS 0.007268f
C139 B.n105 VSUBS 0.007268f
C140 B.n106 VSUBS 0.007268f
C141 B.n107 VSUBS 0.007268f
C142 B.n108 VSUBS 0.007268f
C143 B.n109 VSUBS 0.007268f
C144 B.n110 VSUBS 0.007268f
C145 B.n111 VSUBS 0.007268f
C146 B.n112 VSUBS 0.007268f
C147 B.n113 VSUBS 0.007268f
C148 B.n114 VSUBS 0.007268f
C149 B.n115 VSUBS 0.007268f
C150 B.n116 VSUBS 0.007268f
C151 B.n117 VSUBS 0.007268f
C152 B.n118 VSUBS 0.007268f
C153 B.n119 VSUBS 0.007268f
C154 B.n120 VSUBS 0.007268f
C155 B.n121 VSUBS 0.007268f
C156 B.n122 VSUBS 0.007268f
C157 B.n123 VSUBS 0.007268f
C158 B.n124 VSUBS 0.007268f
C159 B.n125 VSUBS 0.007268f
C160 B.n126 VSUBS 0.007268f
C161 B.n127 VSUBS 0.007268f
C162 B.n128 VSUBS 0.007268f
C163 B.n129 VSUBS 0.007268f
C164 B.n130 VSUBS 0.007268f
C165 B.n131 VSUBS 0.007268f
C166 B.n132 VSUBS 0.016926f
C167 B.n133 VSUBS 0.007268f
C168 B.n134 VSUBS 0.007268f
C169 B.n135 VSUBS 0.007268f
C170 B.n136 VSUBS 0.007268f
C171 B.n137 VSUBS 0.007268f
C172 B.n138 VSUBS 0.007268f
C173 B.n139 VSUBS 0.007268f
C174 B.n140 VSUBS 0.007268f
C175 B.n141 VSUBS 0.007268f
C176 B.n142 VSUBS 0.007268f
C177 B.n143 VSUBS 0.007268f
C178 B.n144 VSUBS 0.007268f
C179 B.n145 VSUBS 0.007268f
C180 B.n146 VSUBS 0.007268f
C181 B.n147 VSUBS 0.007268f
C182 B.n148 VSUBS 0.007268f
C183 B.n149 VSUBS 0.007268f
C184 B.n150 VSUBS 0.007268f
C185 B.n151 VSUBS 0.007268f
C186 B.n152 VSUBS 0.007268f
C187 B.n153 VSUBS 0.007268f
C188 B.n154 VSUBS 0.007268f
C189 B.n155 VSUBS 0.007268f
C190 B.n156 VSUBS 0.007268f
C191 B.n157 VSUBS 0.007268f
C192 B.n158 VSUBS 0.007268f
C193 B.n159 VSUBS 0.007268f
C194 B.n160 VSUBS 0.007268f
C195 B.n161 VSUBS 0.007268f
C196 B.n162 VSUBS 0.007268f
C197 B.n163 VSUBS 0.007268f
C198 B.n164 VSUBS 0.007268f
C199 B.t8 VSUBS 0.407174f
C200 B.t7 VSUBS 0.437402f
C201 B.t6 VSUBS 1.9376f
C202 B.n165 VSUBS 0.645631f
C203 B.n166 VSUBS 0.359854f
C204 B.n167 VSUBS 0.007268f
C205 B.n168 VSUBS 0.007268f
C206 B.n169 VSUBS 0.007268f
C207 B.n170 VSUBS 0.007268f
C208 B.n171 VSUBS 0.004061f
C209 B.n172 VSUBS 0.007268f
C210 B.n173 VSUBS 0.007268f
C211 B.n174 VSUBS 0.007268f
C212 B.n175 VSUBS 0.007268f
C213 B.n176 VSUBS 0.007268f
C214 B.n177 VSUBS 0.007268f
C215 B.n178 VSUBS 0.007268f
C216 B.n179 VSUBS 0.007268f
C217 B.n180 VSUBS 0.007268f
C218 B.n181 VSUBS 0.007268f
C219 B.n182 VSUBS 0.007268f
C220 B.n183 VSUBS 0.007268f
C221 B.n184 VSUBS 0.007268f
C222 B.n185 VSUBS 0.007268f
C223 B.n186 VSUBS 0.007268f
C224 B.n187 VSUBS 0.007268f
C225 B.n188 VSUBS 0.007268f
C226 B.n189 VSUBS 0.007268f
C227 B.n190 VSUBS 0.007268f
C228 B.n191 VSUBS 0.007268f
C229 B.n192 VSUBS 0.007268f
C230 B.n193 VSUBS 0.007268f
C231 B.n194 VSUBS 0.007268f
C232 B.n195 VSUBS 0.007268f
C233 B.n196 VSUBS 0.007268f
C234 B.n197 VSUBS 0.007268f
C235 B.n198 VSUBS 0.007268f
C236 B.n199 VSUBS 0.007268f
C237 B.n200 VSUBS 0.007268f
C238 B.n201 VSUBS 0.007268f
C239 B.n202 VSUBS 0.007268f
C240 B.n203 VSUBS 0.017916f
C241 B.n204 VSUBS 0.007268f
C242 B.n205 VSUBS 0.007268f
C243 B.n206 VSUBS 0.007268f
C244 B.n207 VSUBS 0.007268f
C245 B.n208 VSUBS 0.007268f
C246 B.n209 VSUBS 0.007268f
C247 B.n210 VSUBS 0.007268f
C248 B.n211 VSUBS 0.007268f
C249 B.n212 VSUBS 0.007268f
C250 B.n213 VSUBS 0.007268f
C251 B.n214 VSUBS 0.007268f
C252 B.n215 VSUBS 0.007268f
C253 B.n216 VSUBS 0.007268f
C254 B.n217 VSUBS 0.007268f
C255 B.n218 VSUBS 0.007268f
C256 B.n219 VSUBS 0.007268f
C257 B.n220 VSUBS 0.007268f
C258 B.n221 VSUBS 0.007268f
C259 B.n222 VSUBS 0.007268f
C260 B.n223 VSUBS 0.007268f
C261 B.n224 VSUBS 0.007268f
C262 B.n225 VSUBS 0.007268f
C263 B.n226 VSUBS 0.007268f
C264 B.n227 VSUBS 0.007268f
C265 B.n228 VSUBS 0.007268f
C266 B.n229 VSUBS 0.007268f
C267 B.n230 VSUBS 0.007268f
C268 B.n231 VSUBS 0.007268f
C269 B.n232 VSUBS 0.007268f
C270 B.n233 VSUBS 0.007268f
C271 B.n234 VSUBS 0.007268f
C272 B.n235 VSUBS 0.007268f
C273 B.n236 VSUBS 0.007268f
C274 B.n237 VSUBS 0.007268f
C275 B.n238 VSUBS 0.007268f
C276 B.n239 VSUBS 0.007268f
C277 B.n240 VSUBS 0.007268f
C278 B.n241 VSUBS 0.007268f
C279 B.n242 VSUBS 0.007268f
C280 B.n243 VSUBS 0.007268f
C281 B.n244 VSUBS 0.007268f
C282 B.n245 VSUBS 0.007268f
C283 B.n246 VSUBS 0.007268f
C284 B.n247 VSUBS 0.007268f
C285 B.n248 VSUBS 0.007268f
C286 B.n249 VSUBS 0.007268f
C287 B.n250 VSUBS 0.007268f
C288 B.n251 VSUBS 0.007268f
C289 B.n252 VSUBS 0.007268f
C290 B.n253 VSUBS 0.007268f
C291 B.n254 VSUBS 0.007268f
C292 B.n255 VSUBS 0.007268f
C293 B.n256 VSUBS 0.007268f
C294 B.n257 VSUBS 0.007268f
C295 B.n258 VSUBS 0.007268f
C296 B.n259 VSUBS 0.007268f
C297 B.n260 VSUBS 0.007268f
C298 B.n261 VSUBS 0.007268f
C299 B.n262 VSUBS 0.007268f
C300 B.n263 VSUBS 0.007268f
C301 B.n264 VSUBS 0.007268f
C302 B.n265 VSUBS 0.007268f
C303 B.n266 VSUBS 0.007268f
C304 B.n267 VSUBS 0.007268f
C305 B.n268 VSUBS 0.007268f
C306 B.n269 VSUBS 0.007268f
C307 B.n270 VSUBS 0.007268f
C308 B.n271 VSUBS 0.007268f
C309 B.n272 VSUBS 0.007268f
C310 B.n273 VSUBS 0.007268f
C311 B.n274 VSUBS 0.016926f
C312 B.n275 VSUBS 0.016926f
C313 B.n276 VSUBS 0.017916f
C314 B.n277 VSUBS 0.007268f
C315 B.n278 VSUBS 0.007268f
C316 B.n279 VSUBS 0.007268f
C317 B.n280 VSUBS 0.007268f
C318 B.n281 VSUBS 0.007268f
C319 B.n282 VSUBS 0.007268f
C320 B.n283 VSUBS 0.007268f
C321 B.n284 VSUBS 0.007268f
C322 B.n285 VSUBS 0.007268f
C323 B.n286 VSUBS 0.007268f
C324 B.n287 VSUBS 0.007268f
C325 B.n288 VSUBS 0.007268f
C326 B.n289 VSUBS 0.007268f
C327 B.n290 VSUBS 0.007268f
C328 B.n291 VSUBS 0.007268f
C329 B.n292 VSUBS 0.007268f
C330 B.n293 VSUBS 0.007268f
C331 B.n294 VSUBS 0.007268f
C332 B.n295 VSUBS 0.007268f
C333 B.n296 VSUBS 0.007268f
C334 B.n297 VSUBS 0.007268f
C335 B.n298 VSUBS 0.007268f
C336 B.n299 VSUBS 0.007268f
C337 B.n300 VSUBS 0.007268f
C338 B.n301 VSUBS 0.007268f
C339 B.n302 VSUBS 0.007268f
C340 B.n303 VSUBS 0.007268f
C341 B.n304 VSUBS 0.007268f
C342 B.n305 VSUBS 0.007268f
C343 B.n306 VSUBS 0.007268f
C344 B.n307 VSUBS 0.007268f
C345 B.n308 VSUBS 0.007268f
C346 B.n309 VSUBS 0.007268f
C347 B.n310 VSUBS 0.007268f
C348 B.n311 VSUBS 0.007268f
C349 B.n312 VSUBS 0.007268f
C350 B.n313 VSUBS 0.007268f
C351 B.n314 VSUBS 0.007268f
C352 B.n315 VSUBS 0.007268f
C353 B.n316 VSUBS 0.007268f
C354 B.n317 VSUBS 0.007268f
C355 B.n318 VSUBS 0.007268f
C356 B.n319 VSUBS 0.007268f
C357 B.n320 VSUBS 0.007268f
C358 B.n321 VSUBS 0.007268f
C359 B.n322 VSUBS 0.007268f
C360 B.n323 VSUBS 0.007268f
C361 B.n324 VSUBS 0.007268f
C362 B.n325 VSUBS 0.007268f
C363 B.n326 VSUBS 0.007268f
C364 B.n327 VSUBS 0.007268f
C365 B.n328 VSUBS 0.007268f
C366 B.n329 VSUBS 0.007268f
C367 B.n330 VSUBS 0.007268f
C368 B.n331 VSUBS 0.007268f
C369 B.n332 VSUBS 0.007268f
C370 B.n333 VSUBS 0.007268f
C371 B.n334 VSUBS 0.007268f
C372 B.n335 VSUBS 0.007268f
C373 B.n336 VSUBS 0.007268f
C374 B.n337 VSUBS 0.007268f
C375 B.n338 VSUBS 0.007268f
C376 B.n339 VSUBS 0.007268f
C377 B.n340 VSUBS 0.007268f
C378 B.n341 VSUBS 0.007268f
C379 B.n342 VSUBS 0.007268f
C380 B.n343 VSUBS 0.007268f
C381 B.n344 VSUBS 0.007268f
C382 B.n345 VSUBS 0.007268f
C383 B.n346 VSUBS 0.007268f
C384 B.n347 VSUBS 0.007268f
C385 B.n348 VSUBS 0.007268f
C386 B.n349 VSUBS 0.007268f
C387 B.n350 VSUBS 0.007268f
C388 B.n351 VSUBS 0.007268f
C389 B.n352 VSUBS 0.007268f
C390 B.n353 VSUBS 0.007268f
C391 B.n354 VSUBS 0.007268f
C392 B.n355 VSUBS 0.007268f
C393 B.n356 VSUBS 0.007268f
C394 B.n357 VSUBS 0.007268f
C395 B.n358 VSUBS 0.007268f
C396 B.n359 VSUBS 0.007268f
C397 B.n360 VSUBS 0.007268f
C398 B.n361 VSUBS 0.007268f
C399 B.n362 VSUBS 0.007268f
C400 B.n363 VSUBS 0.007268f
C401 B.n364 VSUBS 0.007268f
C402 B.n365 VSUBS 0.007268f
C403 B.n366 VSUBS 0.007268f
C404 B.n367 VSUBS 0.007268f
C405 B.n368 VSUBS 0.007268f
C406 B.n369 VSUBS 0.007268f
C407 B.t11 VSUBS 0.407171f
C408 B.t10 VSUBS 0.437399f
C409 B.t9 VSUBS 1.9376f
C410 B.n370 VSUBS 0.645634f
C411 B.n371 VSUBS 0.359858f
C412 B.n372 VSUBS 0.016838f
C413 B.n373 VSUBS 0.00684f
C414 B.n374 VSUBS 0.007268f
C415 B.n375 VSUBS 0.007268f
C416 B.n376 VSUBS 0.007268f
C417 B.n377 VSUBS 0.007268f
C418 B.n378 VSUBS 0.007268f
C419 B.n379 VSUBS 0.007268f
C420 B.n380 VSUBS 0.007268f
C421 B.n381 VSUBS 0.007268f
C422 B.n382 VSUBS 0.007268f
C423 B.n383 VSUBS 0.007268f
C424 B.n384 VSUBS 0.007268f
C425 B.n385 VSUBS 0.007268f
C426 B.n386 VSUBS 0.007268f
C427 B.n387 VSUBS 0.007268f
C428 B.n388 VSUBS 0.007268f
C429 B.n389 VSUBS 0.004061f
C430 B.n390 VSUBS 0.016838f
C431 B.n391 VSUBS 0.00684f
C432 B.n392 VSUBS 0.007268f
C433 B.n393 VSUBS 0.007268f
C434 B.n394 VSUBS 0.007268f
C435 B.n395 VSUBS 0.007268f
C436 B.n396 VSUBS 0.007268f
C437 B.n397 VSUBS 0.007268f
C438 B.n398 VSUBS 0.007268f
C439 B.n399 VSUBS 0.007268f
C440 B.n400 VSUBS 0.007268f
C441 B.n401 VSUBS 0.007268f
C442 B.n402 VSUBS 0.007268f
C443 B.n403 VSUBS 0.007268f
C444 B.n404 VSUBS 0.007268f
C445 B.n405 VSUBS 0.007268f
C446 B.n406 VSUBS 0.007268f
C447 B.n407 VSUBS 0.007268f
C448 B.n408 VSUBS 0.007268f
C449 B.n409 VSUBS 0.007268f
C450 B.n410 VSUBS 0.007268f
C451 B.n411 VSUBS 0.007268f
C452 B.n412 VSUBS 0.007268f
C453 B.n413 VSUBS 0.007268f
C454 B.n414 VSUBS 0.007268f
C455 B.n415 VSUBS 0.007268f
C456 B.n416 VSUBS 0.007268f
C457 B.n417 VSUBS 0.007268f
C458 B.n418 VSUBS 0.007268f
C459 B.n419 VSUBS 0.007268f
C460 B.n420 VSUBS 0.007268f
C461 B.n421 VSUBS 0.007268f
C462 B.n422 VSUBS 0.007268f
C463 B.n423 VSUBS 0.007268f
C464 B.n424 VSUBS 0.007268f
C465 B.n425 VSUBS 0.007268f
C466 B.n426 VSUBS 0.007268f
C467 B.n427 VSUBS 0.007268f
C468 B.n428 VSUBS 0.007268f
C469 B.n429 VSUBS 0.007268f
C470 B.n430 VSUBS 0.007268f
C471 B.n431 VSUBS 0.007268f
C472 B.n432 VSUBS 0.007268f
C473 B.n433 VSUBS 0.007268f
C474 B.n434 VSUBS 0.007268f
C475 B.n435 VSUBS 0.007268f
C476 B.n436 VSUBS 0.007268f
C477 B.n437 VSUBS 0.007268f
C478 B.n438 VSUBS 0.007268f
C479 B.n439 VSUBS 0.007268f
C480 B.n440 VSUBS 0.007268f
C481 B.n441 VSUBS 0.007268f
C482 B.n442 VSUBS 0.007268f
C483 B.n443 VSUBS 0.007268f
C484 B.n444 VSUBS 0.007268f
C485 B.n445 VSUBS 0.007268f
C486 B.n446 VSUBS 0.007268f
C487 B.n447 VSUBS 0.007268f
C488 B.n448 VSUBS 0.007268f
C489 B.n449 VSUBS 0.007268f
C490 B.n450 VSUBS 0.007268f
C491 B.n451 VSUBS 0.007268f
C492 B.n452 VSUBS 0.007268f
C493 B.n453 VSUBS 0.007268f
C494 B.n454 VSUBS 0.007268f
C495 B.n455 VSUBS 0.007268f
C496 B.n456 VSUBS 0.007268f
C497 B.n457 VSUBS 0.007268f
C498 B.n458 VSUBS 0.007268f
C499 B.n459 VSUBS 0.007268f
C500 B.n460 VSUBS 0.007268f
C501 B.n461 VSUBS 0.007268f
C502 B.n462 VSUBS 0.007268f
C503 B.n463 VSUBS 0.007268f
C504 B.n464 VSUBS 0.007268f
C505 B.n465 VSUBS 0.007268f
C506 B.n466 VSUBS 0.007268f
C507 B.n467 VSUBS 0.007268f
C508 B.n468 VSUBS 0.007268f
C509 B.n469 VSUBS 0.007268f
C510 B.n470 VSUBS 0.007268f
C511 B.n471 VSUBS 0.007268f
C512 B.n472 VSUBS 0.007268f
C513 B.n473 VSUBS 0.007268f
C514 B.n474 VSUBS 0.007268f
C515 B.n475 VSUBS 0.007268f
C516 B.n476 VSUBS 0.007268f
C517 B.n477 VSUBS 0.007268f
C518 B.n478 VSUBS 0.007268f
C519 B.n479 VSUBS 0.007268f
C520 B.n480 VSUBS 0.007268f
C521 B.n481 VSUBS 0.007268f
C522 B.n482 VSUBS 0.007268f
C523 B.n483 VSUBS 0.007268f
C524 B.n484 VSUBS 0.007268f
C525 B.n485 VSUBS 0.017916f
C526 B.n486 VSUBS 0.017088f
C527 B.n487 VSUBS 0.017754f
C528 B.n488 VSUBS 0.007268f
C529 B.n489 VSUBS 0.007268f
C530 B.n490 VSUBS 0.007268f
C531 B.n491 VSUBS 0.007268f
C532 B.n492 VSUBS 0.007268f
C533 B.n493 VSUBS 0.007268f
C534 B.n494 VSUBS 0.007268f
C535 B.n495 VSUBS 0.007268f
C536 B.n496 VSUBS 0.007268f
C537 B.n497 VSUBS 0.007268f
C538 B.n498 VSUBS 0.007268f
C539 B.n499 VSUBS 0.007268f
C540 B.n500 VSUBS 0.007268f
C541 B.n501 VSUBS 0.007268f
C542 B.n502 VSUBS 0.007268f
C543 B.n503 VSUBS 0.007268f
C544 B.n504 VSUBS 0.007268f
C545 B.n505 VSUBS 0.007268f
C546 B.n506 VSUBS 0.007268f
C547 B.n507 VSUBS 0.007268f
C548 B.n508 VSUBS 0.007268f
C549 B.n509 VSUBS 0.007268f
C550 B.n510 VSUBS 0.007268f
C551 B.n511 VSUBS 0.007268f
C552 B.n512 VSUBS 0.007268f
C553 B.n513 VSUBS 0.007268f
C554 B.n514 VSUBS 0.007268f
C555 B.n515 VSUBS 0.007268f
C556 B.n516 VSUBS 0.007268f
C557 B.n517 VSUBS 0.007268f
C558 B.n518 VSUBS 0.007268f
C559 B.n519 VSUBS 0.007268f
C560 B.n520 VSUBS 0.007268f
C561 B.n521 VSUBS 0.007268f
C562 B.n522 VSUBS 0.007268f
C563 B.n523 VSUBS 0.007268f
C564 B.n524 VSUBS 0.007268f
C565 B.n525 VSUBS 0.007268f
C566 B.n526 VSUBS 0.007268f
C567 B.n527 VSUBS 0.007268f
C568 B.n528 VSUBS 0.007268f
C569 B.n529 VSUBS 0.007268f
C570 B.n530 VSUBS 0.007268f
C571 B.n531 VSUBS 0.007268f
C572 B.n532 VSUBS 0.007268f
C573 B.n533 VSUBS 0.007268f
C574 B.n534 VSUBS 0.007268f
C575 B.n535 VSUBS 0.007268f
C576 B.n536 VSUBS 0.007268f
C577 B.n537 VSUBS 0.007268f
C578 B.n538 VSUBS 0.007268f
C579 B.n539 VSUBS 0.007268f
C580 B.n540 VSUBS 0.007268f
C581 B.n541 VSUBS 0.007268f
C582 B.n542 VSUBS 0.007268f
C583 B.n543 VSUBS 0.007268f
C584 B.n544 VSUBS 0.007268f
C585 B.n545 VSUBS 0.007268f
C586 B.n546 VSUBS 0.007268f
C587 B.n547 VSUBS 0.007268f
C588 B.n548 VSUBS 0.007268f
C589 B.n549 VSUBS 0.007268f
C590 B.n550 VSUBS 0.007268f
C591 B.n551 VSUBS 0.007268f
C592 B.n552 VSUBS 0.007268f
C593 B.n553 VSUBS 0.007268f
C594 B.n554 VSUBS 0.007268f
C595 B.n555 VSUBS 0.007268f
C596 B.n556 VSUBS 0.007268f
C597 B.n557 VSUBS 0.007268f
C598 B.n558 VSUBS 0.007268f
C599 B.n559 VSUBS 0.007268f
C600 B.n560 VSUBS 0.007268f
C601 B.n561 VSUBS 0.007268f
C602 B.n562 VSUBS 0.007268f
C603 B.n563 VSUBS 0.007268f
C604 B.n564 VSUBS 0.007268f
C605 B.n565 VSUBS 0.007268f
C606 B.n566 VSUBS 0.007268f
C607 B.n567 VSUBS 0.007268f
C608 B.n568 VSUBS 0.007268f
C609 B.n569 VSUBS 0.007268f
C610 B.n570 VSUBS 0.007268f
C611 B.n571 VSUBS 0.007268f
C612 B.n572 VSUBS 0.007268f
C613 B.n573 VSUBS 0.007268f
C614 B.n574 VSUBS 0.007268f
C615 B.n575 VSUBS 0.007268f
C616 B.n576 VSUBS 0.007268f
C617 B.n577 VSUBS 0.007268f
C618 B.n578 VSUBS 0.007268f
C619 B.n579 VSUBS 0.007268f
C620 B.n580 VSUBS 0.007268f
C621 B.n581 VSUBS 0.007268f
C622 B.n582 VSUBS 0.007268f
C623 B.n583 VSUBS 0.007268f
C624 B.n584 VSUBS 0.007268f
C625 B.n585 VSUBS 0.007268f
C626 B.n586 VSUBS 0.007268f
C627 B.n587 VSUBS 0.007268f
C628 B.n588 VSUBS 0.007268f
C629 B.n589 VSUBS 0.007268f
C630 B.n590 VSUBS 0.007268f
C631 B.n591 VSUBS 0.007268f
C632 B.n592 VSUBS 0.007268f
C633 B.n593 VSUBS 0.007268f
C634 B.n594 VSUBS 0.007268f
C635 B.n595 VSUBS 0.007268f
C636 B.n596 VSUBS 0.007268f
C637 B.n597 VSUBS 0.007268f
C638 B.n598 VSUBS 0.007268f
C639 B.n599 VSUBS 0.016926f
C640 B.n600 VSUBS 0.016926f
C641 B.n601 VSUBS 0.017916f
C642 B.n602 VSUBS 0.007268f
C643 B.n603 VSUBS 0.007268f
C644 B.n604 VSUBS 0.007268f
C645 B.n605 VSUBS 0.007268f
C646 B.n606 VSUBS 0.007268f
C647 B.n607 VSUBS 0.007268f
C648 B.n608 VSUBS 0.007268f
C649 B.n609 VSUBS 0.007268f
C650 B.n610 VSUBS 0.007268f
C651 B.n611 VSUBS 0.007268f
C652 B.n612 VSUBS 0.007268f
C653 B.n613 VSUBS 0.007268f
C654 B.n614 VSUBS 0.007268f
C655 B.n615 VSUBS 0.007268f
C656 B.n616 VSUBS 0.007268f
C657 B.n617 VSUBS 0.007268f
C658 B.n618 VSUBS 0.007268f
C659 B.n619 VSUBS 0.007268f
C660 B.n620 VSUBS 0.007268f
C661 B.n621 VSUBS 0.007268f
C662 B.n622 VSUBS 0.007268f
C663 B.n623 VSUBS 0.007268f
C664 B.n624 VSUBS 0.007268f
C665 B.n625 VSUBS 0.007268f
C666 B.n626 VSUBS 0.007268f
C667 B.n627 VSUBS 0.007268f
C668 B.n628 VSUBS 0.007268f
C669 B.n629 VSUBS 0.007268f
C670 B.n630 VSUBS 0.007268f
C671 B.n631 VSUBS 0.007268f
C672 B.n632 VSUBS 0.007268f
C673 B.n633 VSUBS 0.007268f
C674 B.n634 VSUBS 0.007268f
C675 B.n635 VSUBS 0.007268f
C676 B.n636 VSUBS 0.007268f
C677 B.n637 VSUBS 0.007268f
C678 B.n638 VSUBS 0.007268f
C679 B.n639 VSUBS 0.007268f
C680 B.n640 VSUBS 0.007268f
C681 B.n641 VSUBS 0.007268f
C682 B.n642 VSUBS 0.007268f
C683 B.n643 VSUBS 0.007268f
C684 B.n644 VSUBS 0.007268f
C685 B.n645 VSUBS 0.007268f
C686 B.n646 VSUBS 0.007268f
C687 B.n647 VSUBS 0.007268f
C688 B.n648 VSUBS 0.007268f
C689 B.n649 VSUBS 0.007268f
C690 B.n650 VSUBS 0.007268f
C691 B.n651 VSUBS 0.007268f
C692 B.n652 VSUBS 0.007268f
C693 B.n653 VSUBS 0.007268f
C694 B.n654 VSUBS 0.007268f
C695 B.n655 VSUBS 0.007268f
C696 B.n656 VSUBS 0.007268f
C697 B.n657 VSUBS 0.007268f
C698 B.n658 VSUBS 0.007268f
C699 B.n659 VSUBS 0.007268f
C700 B.n660 VSUBS 0.007268f
C701 B.n661 VSUBS 0.007268f
C702 B.n662 VSUBS 0.007268f
C703 B.n663 VSUBS 0.007268f
C704 B.n664 VSUBS 0.007268f
C705 B.n665 VSUBS 0.007268f
C706 B.n666 VSUBS 0.007268f
C707 B.n667 VSUBS 0.007268f
C708 B.n668 VSUBS 0.007268f
C709 B.n669 VSUBS 0.007268f
C710 B.n670 VSUBS 0.007268f
C711 B.n671 VSUBS 0.007268f
C712 B.n672 VSUBS 0.007268f
C713 B.n673 VSUBS 0.007268f
C714 B.n674 VSUBS 0.007268f
C715 B.n675 VSUBS 0.007268f
C716 B.n676 VSUBS 0.007268f
C717 B.n677 VSUBS 0.007268f
C718 B.n678 VSUBS 0.007268f
C719 B.n679 VSUBS 0.007268f
C720 B.n680 VSUBS 0.007268f
C721 B.n681 VSUBS 0.007268f
C722 B.n682 VSUBS 0.007268f
C723 B.n683 VSUBS 0.007268f
C724 B.n684 VSUBS 0.007268f
C725 B.n685 VSUBS 0.007268f
C726 B.n686 VSUBS 0.007268f
C727 B.n687 VSUBS 0.007268f
C728 B.n688 VSUBS 0.007268f
C729 B.n689 VSUBS 0.007268f
C730 B.n690 VSUBS 0.007268f
C731 B.n691 VSUBS 0.007268f
C732 B.n692 VSUBS 0.007268f
C733 B.n693 VSUBS 0.007268f
C734 B.n694 VSUBS 0.007268f
C735 B.n695 VSUBS 0.007268f
C736 B.n696 VSUBS 0.00684f
C737 B.n697 VSUBS 0.016838f
C738 B.n698 VSUBS 0.004061f
C739 B.n699 VSUBS 0.007268f
C740 B.n700 VSUBS 0.007268f
C741 B.n701 VSUBS 0.007268f
C742 B.n702 VSUBS 0.007268f
C743 B.n703 VSUBS 0.007268f
C744 B.n704 VSUBS 0.007268f
C745 B.n705 VSUBS 0.007268f
C746 B.n706 VSUBS 0.007268f
C747 B.n707 VSUBS 0.007268f
C748 B.n708 VSUBS 0.007268f
C749 B.n709 VSUBS 0.007268f
C750 B.n710 VSUBS 0.007268f
C751 B.n711 VSUBS 0.004061f
C752 B.n712 VSUBS 0.007268f
C753 B.n713 VSUBS 0.007268f
C754 B.n714 VSUBS 0.007268f
C755 B.n715 VSUBS 0.007268f
C756 B.n716 VSUBS 0.007268f
C757 B.n717 VSUBS 0.007268f
C758 B.n718 VSUBS 0.007268f
C759 B.n719 VSUBS 0.007268f
C760 B.n720 VSUBS 0.007268f
C761 B.n721 VSUBS 0.007268f
C762 B.n722 VSUBS 0.007268f
C763 B.n723 VSUBS 0.007268f
C764 B.n724 VSUBS 0.007268f
C765 B.n725 VSUBS 0.007268f
C766 B.n726 VSUBS 0.007268f
C767 B.n727 VSUBS 0.007268f
C768 B.n728 VSUBS 0.007268f
C769 B.n729 VSUBS 0.007268f
C770 B.n730 VSUBS 0.007268f
C771 B.n731 VSUBS 0.007268f
C772 B.n732 VSUBS 0.007268f
C773 B.n733 VSUBS 0.007268f
C774 B.n734 VSUBS 0.007268f
C775 B.n735 VSUBS 0.007268f
C776 B.n736 VSUBS 0.007268f
C777 B.n737 VSUBS 0.007268f
C778 B.n738 VSUBS 0.007268f
C779 B.n739 VSUBS 0.007268f
C780 B.n740 VSUBS 0.007268f
C781 B.n741 VSUBS 0.007268f
C782 B.n742 VSUBS 0.007268f
C783 B.n743 VSUBS 0.007268f
C784 B.n744 VSUBS 0.007268f
C785 B.n745 VSUBS 0.007268f
C786 B.n746 VSUBS 0.007268f
C787 B.n747 VSUBS 0.007268f
C788 B.n748 VSUBS 0.007268f
C789 B.n749 VSUBS 0.007268f
C790 B.n750 VSUBS 0.007268f
C791 B.n751 VSUBS 0.007268f
C792 B.n752 VSUBS 0.007268f
C793 B.n753 VSUBS 0.007268f
C794 B.n754 VSUBS 0.007268f
C795 B.n755 VSUBS 0.007268f
C796 B.n756 VSUBS 0.007268f
C797 B.n757 VSUBS 0.007268f
C798 B.n758 VSUBS 0.007268f
C799 B.n759 VSUBS 0.007268f
C800 B.n760 VSUBS 0.007268f
C801 B.n761 VSUBS 0.007268f
C802 B.n762 VSUBS 0.007268f
C803 B.n763 VSUBS 0.007268f
C804 B.n764 VSUBS 0.007268f
C805 B.n765 VSUBS 0.007268f
C806 B.n766 VSUBS 0.007268f
C807 B.n767 VSUBS 0.007268f
C808 B.n768 VSUBS 0.007268f
C809 B.n769 VSUBS 0.007268f
C810 B.n770 VSUBS 0.007268f
C811 B.n771 VSUBS 0.007268f
C812 B.n772 VSUBS 0.007268f
C813 B.n773 VSUBS 0.007268f
C814 B.n774 VSUBS 0.007268f
C815 B.n775 VSUBS 0.007268f
C816 B.n776 VSUBS 0.007268f
C817 B.n777 VSUBS 0.007268f
C818 B.n778 VSUBS 0.007268f
C819 B.n779 VSUBS 0.007268f
C820 B.n780 VSUBS 0.007268f
C821 B.n781 VSUBS 0.007268f
C822 B.n782 VSUBS 0.007268f
C823 B.n783 VSUBS 0.007268f
C824 B.n784 VSUBS 0.007268f
C825 B.n785 VSUBS 0.007268f
C826 B.n786 VSUBS 0.007268f
C827 B.n787 VSUBS 0.007268f
C828 B.n788 VSUBS 0.007268f
C829 B.n789 VSUBS 0.007268f
C830 B.n790 VSUBS 0.007268f
C831 B.n791 VSUBS 0.007268f
C832 B.n792 VSUBS 0.007268f
C833 B.n793 VSUBS 0.007268f
C834 B.n794 VSUBS 0.007268f
C835 B.n795 VSUBS 0.007268f
C836 B.n796 VSUBS 0.007268f
C837 B.n797 VSUBS 0.007268f
C838 B.n798 VSUBS 0.007268f
C839 B.n799 VSUBS 0.007268f
C840 B.n800 VSUBS 0.007268f
C841 B.n801 VSUBS 0.007268f
C842 B.n802 VSUBS 0.007268f
C843 B.n803 VSUBS 0.007268f
C844 B.n804 VSUBS 0.007268f
C845 B.n805 VSUBS 0.007268f
C846 B.n806 VSUBS 0.007268f
C847 B.n807 VSUBS 0.017916f
C848 B.n808 VSUBS 0.017916f
C849 B.n809 VSUBS 0.016926f
C850 B.n810 VSUBS 0.007268f
C851 B.n811 VSUBS 0.007268f
C852 B.n812 VSUBS 0.007268f
C853 B.n813 VSUBS 0.007268f
C854 B.n814 VSUBS 0.007268f
C855 B.n815 VSUBS 0.007268f
C856 B.n816 VSUBS 0.007268f
C857 B.n817 VSUBS 0.007268f
C858 B.n818 VSUBS 0.007268f
C859 B.n819 VSUBS 0.007268f
C860 B.n820 VSUBS 0.007268f
C861 B.n821 VSUBS 0.007268f
C862 B.n822 VSUBS 0.007268f
C863 B.n823 VSUBS 0.007268f
C864 B.n824 VSUBS 0.007268f
C865 B.n825 VSUBS 0.007268f
C866 B.n826 VSUBS 0.007268f
C867 B.n827 VSUBS 0.007268f
C868 B.n828 VSUBS 0.007268f
C869 B.n829 VSUBS 0.007268f
C870 B.n830 VSUBS 0.007268f
C871 B.n831 VSUBS 0.007268f
C872 B.n832 VSUBS 0.007268f
C873 B.n833 VSUBS 0.007268f
C874 B.n834 VSUBS 0.007268f
C875 B.n835 VSUBS 0.007268f
C876 B.n836 VSUBS 0.007268f
C877 B.n837 VSUBS 0.007268f
C878 B.n838 VSUBS 0.007268f
C879 B.n839 VSUBS 0.007268f
C880 B.n840 VSUBS 0.007268f
C881 B.n841 VSUBS 0.007268f
C882 B.n842 VSUBS 0.007268f
C883 B.n843 VSUBS 0.007268f
C884 B.n844 VSUBS 0.007268f
C885 B.n845 VSUBS 0.007268f
C886 B.n846 VSUBS 0.007268f
C887 B.n847 VSUBS 0.007268f
C888 B.n848 VSUBS 0.007268f
C889 B.n849 VSUBS 0.007268f
C890 B.n850 VSUBS 0.007268f
C891 B.n851 VSUBS 0.007268f
C892 B.n852 VSUBS 0.007268f
C893 B.n853 VSUBS 0.007268f
C894 B.n854 VSUBS 0.007268f
C895 B.n855 VSUBS 0.007268f
C896 B.n856 VSUBS 0.007268f
C897 B.n857 VSUBS 0.007268f
C898 B.n858 VSUBS 0.007268f
C899 B.n859 VSUBS 0.007268f
C900 B.n860 VSUBS 0.007268f
C901 B.n861 VSUBS 0.007268f
C902 B.n862 VSUBS 0.007268f
C903 B.n863 VSUBS 0.009484f
C904 B.n864 VSUBS 0.010103f
C905 B.n865 VSUBS 0.02009f
C906 VDD2.n0 VSUBS 0.030071f
C907 VDD2.n1 VSUBS 0.026647f
C908 VDD2.n2 VSUBS 0.014319f
C909 VDD2.n3 VSUBS 0.033845f
C910 VDD2.n4 VSUBS 0.015161f
C911 VDD2.n5 VSUBS 0.026647f
C912 VDD2.n6 VSUBS 0.014319f
C913 VDD2.n7 VSUBS 0.033845f
C914 VDD2.n8 VSUBS 0.015161f
C915 VDD2.n9 VSUBS 0.026647f
C916 VDD2.n10 VSUBS 0.014319f
C917 VDD2.n11 VSUBS 0.033845f
C918 VDD2.n12 VSUBS 0.01474f
C919 VDD2.n13 VSUBS 0.026647f
C920 VDD2.n14 VSUBS 0.015161f
C921 VDD2.n15 VSUBS 0.033845f
C922 VDD2.n16 VSUBS 0.015161f
C923 VDD2.n17 VSUBS 0.026647f
C924 VDD2.n18 VSUBS 0.014319f
C925 VDD2.n19 VSUBS 0.033845f
C926 VDD2.n20 VSUBS 0.015161f
C927 VDD2.n21 VSUBS 0.026647f
C928 VDD2.n22 VSUBS 0.014319f
C929 VDD2.n23 VSUBS 0.033845f
C930 VDD2.n24 VSUBS 0.015161f
C931 VDD2.n25 VSUBS 0.026647f
C932 VDD2.n26 VSUBS 0.014319f
C933 VDD2.n27 VSUBS 0.033845f
C934 VDD2.n28 VSUBS 0.015161f
C935 VDD2.n29 VSUBS 0.026647f
C936 VDD2.n30 VSUBS 0.014319f
C937 VDD2.n31 VSUBS 0.033845f
C938 VDD2.n32 VSUBS 0.015161f
C939 VDD2.n33 VSUBS 2.2676f
C940 VDD2.n34 VSUBS 0.014319f
C941 VDD2.t0 VSUBS 0.072765f
C942 VDD2.n35 VSUBS 0.224621f
C943 VDD2.n36 VSUBS 0.02153f
C944 VDD2.n37 VSUBS 0.025384f
C945 VDD2.n38 VSUBS 0.033845f
C946 VDD2.n39 VSUBS 0.015161f
C947 VDD2.n40 VSUBS 0.014319f
C948 VDD2.n41 VSUBS 0.026647f
C949 VDD2.n42 VSUBS 0.026647f
C950 VDD2.n43 VSUBS 0.014319f
C951 VDD2.n44 VSUBS 0.015161f
C952 VDD2.n45 VSUBS 0.033845f
C953 VDD2.n46 VSUBS 0.033845f
C954 VDD2.n47 VSUBS 0.015161f
C955 VDD2.n48 VSUBS 0.014319f
C956 VDD2.n49 VSUBS 0.026647f
C957 VDD2.n50 VSUBS 0.026647f
C958 VDD2.n51 VSUBS 0.014319f
C959 VDD2.n52 VSUBS 0.015161f
C960 VDD2.n53 VSUBS 0.033845f
C961 VDD2.n54 VSUBS 0.033845f
C962 VDD2.n55 VSUBS 0.015161f
C963 VDD2.n56 VSUBS 0.014319f
C964 VDD2.n57 VSUBS 0.026647f
C965 VDD2.n58 VSUBS 0.026647f
C966 VDD2.n59 VSUBS 0.014319f
C967 VDD2.n60 VSUBS 0.015161f
C968 VDD2.n61 VSUBS 0.033845f
C969 VDD2.n62 VSUBS 0.033845f
C970 VDD2.n63 VSUBS 0.015161f
C971 VDD2.n64 VSUBS 0.014319f
C972 VDD2.n65 VSUBS 0.026647f
C973 VDD2.n66 VSUBS 0.026647f
C974 VDD2.n67 VSUBS 0.014319f
C975 VDD2.n68 VSUBS 0.015161f
C976 VDD2.n69 VSUBS 0.033845f
C977 VDD2.n70 VSUBS 0.033845f
C978 VDD2.n71 VSUBS 0.015161f
C979 VDD2.n72 VSUBS 0.014319f
C980 VDD2.n73 VSUBS 0.026647f
C981 VDD2.n74 VSUBS 0.026647f
C982 VDD2.n75 VSUBS 0.014319f
C983 VDD2.n76 VSUBS 0.014319f
C984 VDD2.n77 VSUBS 0.015161f
C985 VDD2.n78 VSUBS 0.033845f
C986 VDD2.n79 VSUBS 0.033845f
C987 VDD2.n80 VSUBS 0.033845f
C988 VDD2.n81 VSUBS 0.01474f
C989 VDD2.n82 VSUBS 0.014319f
C990 VDD2.n83 VSUBS 0.026647f
C991 VDD2.n84 VSUBS 0.026647f
C992 VDD2.n85 VSUBS 0.014319f
C993 VDD2.n86 VSUBS 0.015161f
C994 VDD2.n87 VSUBS 0.033845f
C995 VDD2.n88 VSUBS 0.033845f
C996 VDD2.n89 VSUBS 0.015161f
C997 VDD2.n90 VSUBS 0.014319f
C998 VDD2.n91 VSUBS 0.026647f
C999 VDD2.n92 VSUBS 0.026647f
C1000 VDD2.n93 VSUBS 0.014319f
C1001 VDD2.n94 VSUBS 0.015161f
C1002 VDD2.n95 VSUBS 0.033845f
C1003 VDD2.n96 VSUBS 0.033845f
C1004 VDD2.n97 VSUBS 0.015161f
C1005 VDD2.n98 VSUBS 0.014319f
C1006 VDD2.n99 VSUBS 0.026647f
C1007 VDD2.n100 VSUBS 0.026647f
C1008 VDD2.n101 VSUBS 0.014319f
C1009 VDD2.n102 VSUBS 0.015161f
C1010 VDD2.n103 VSUBS 0.033845f
C1011 VDD2.n104 VSUBS 0.084633f
C1012 VDD2.n105 VSUBS 0.015161f
C1013 VDD2.n106 VSUBS 0.014319f
C1014 VDD2.n107 VSUBS 0.061593f
C1015 VDD2.n108 VSUBS 0.06687f
C1016 VDD2.t1 VSUBS 0.414406f
C1017 VDD2.t3 VSUBS 0.414406f
C1018 VDD2.n109 VSUBS 3.48317f
C1019 VDD2.n110 VSUBS 3.48491f
C1020 VDD2.n111 VSUBS 0.030071f
C1021 VDD2.n112 VSUBS 0.026647f
C1022 VDD2.n113 VSUBS 0.014319f
C1023 VDD2.n114 VSUBS 0.033845f
C1024 VDD2.n115 VSUBS 0.015161f
C1025 VDD2.n116 VSUBS 0.026647f
C1026 VDD2.n117 VSUBS 0.014319f
C1027 VDD2.n118 VSUBS 0.033845f
C1028 VDD2.n119 VSUBS 0.015161f
C1029 VDD2.n120 VSUBS 0.026647f
C1030 VDD2.n121 VSUBS 0.014319f
C1031 VDD2.n122 VSUBS 0.033845f
C1032 VDD2.n123 VSUBS 0.01474f
C1033 VDD2.n124 VSUBS 0.026647f
C1034 VDD2.n125 VSUBS 0.01474f
C1035 VDD2.n126 VSUBS 0.014319f
C1036 VDD2.n127 VSUBS 0.033845f
C1037 VDD2.n128 VSUBS 0.033845f
C1038 VDD2.n129 VSUBS 0.015161f
C1039 VDD2.n130 VSUBS 0.026647f
C1040 VDD2.n131 VSUBS 0.014319f
C1041 VDD2.n132 VSUBS 0.033845f
C1042 VDD2.n133 VSUBS 0.015161f
C1043 VDD2.n134 VSUBS 0.026647f
C1044 VDD2.n135 VSUBS 0.014319f
C1045 VDD2.n136 VSUBS 0.033845f
C1046 VDD2.n137 VSUBS 0.015161f
C1047 VDD2.n138 VSUBS 0.026647f
C1048 VDD2.n139 VSUBS 0.014319f
C1049 VDD2.n140 VSUBS 0.033845f
C1050 VDD2.n141 VSUBS 0.015161f
C1051 VDD2.n142 VSUBS 0.026647f
C1052 VDD2.n143 VSUBS 0.014319f
C1053 VDD2.n144 VSUBS 0.033845f
C1054 VDD2.n145 VSUBS 0.015161f
C1055 VDD2.n146 VSUBS 2.2676f
C1056 VDD2.n147 VSUBS 0.014319f
C1057 VDD2.t5 VSUBS 0.072765f
C1058 VDD2.n148 VSUBS 0.224621f
C1059 VDD2.n149 VSUBS 0.02153f
C1060 VDD2.n150 VSUBS 0.025384f
C1061 VDD2.n151 VSUBS 0.033845f
C1062 VDD2.n152 VSUBS 0.015161f
C1063 VDD2.n153 VSUBS 0.014319f
C1064 VDD2.n154 VSUBS 0.026647f
C1065 VDD2.n155 VSUBS 0.026647f
C1066 VDD2.n156 VSUBS 0.014319f
C1067 VDD2.n157 VSUBS 0.015161f
C1068 VDD2.n158 VSUBS 0.033845f
C1069 VDD2.n159 VSUBS 0.033845f
C1070 VDD2.n160 VSUBS 0.015161f
C1071 VDD2.n161 VSUBS 0.014319f
C1072 VDD2.n162 VSUBS 0.026647f
C1073 VDD2.n163 VSUBS 0.026647f
C1074 VDD2.n164 VSUBS 0.014319f
C1075 VDD2.n165 VSUBS 0.015161f
C1076 VDD2.n166 VSUBS 0.033845f
C1077 VDD2.n167 VSUBS 0.033845f
C1078 VDD2.n168 VSUBS 0.015161f
C1079 VDD2.n169 VSUBS 0.014319f
C1080 VDD2.n170 VSUBS 0.026647f
C1081 VDD2.n171 VSUBS 0.026647f
C1082 VDD2.n172 VSUBS 0.014319f
C1083 VDD2.n173 VSUBS 0.015161f
C1084 VDD2.n174 VSUBS 0.033845f
C1085 VDD2.n175 VSUBS 0.033845f
C1086 VDD2.n176 VSUBS 0.015161f
C1087 VDD2.n177 VSUBS 0.014319f
C1088 VDD2.n178 VSUBS 0.026647f
C1089 VDD2.n179 VSUBS 0.026647f
C1090 VDD2.n180 VSUBS 0.014319f
C1091 VDD2.n181 VSUBS 0.015161f
C1092 VDD2.n182 VSUBS 0.033845f
C1093 VDD2.n183 VSUBS 0.033845f
C1094 VDD2.n184 VSUBS 0.015161f
C1095 VDD2.n185 VSUBS 0.014319f
C1096 VDD2.n186 VSUBS 0.026647f
C1097 VDD2.n187 VSUBS 0.026647f
C1098 VDD2.n188 VSUBS 0.014319f
C1099 VDD2.n189 VSUBS 0.015161f
C1100 VDD2.n190 VSUBS 0.033845f
C1101 VDD2.n191 VSUBS 0.033845f
C1102 VDD2.n192 VSUBS 0.015161f
C1103 VDD2.n193 VSUBS 0.014319f
C1104 VDD2.n194 VSUBS 0.026647f
C1105 VDD2.n195 VSUBS 0.026647f
C1106 VDD2.n196 VSUBS 0.014319f
C1107 VDD2.n197 VSUBS 0.015161f
C1108 VDD2.n198 VSUBS 0.033845f
C1109 VDD2.n199 VSUBS 0.033845f
C1110 VDD2.n200 VSUBS 0.015161f
C1111 VDD2.n201 VSUBS 0.014319f
C1112 VDD2.n202 VSUBS 0.026647f
C1113 VDD2.n203 VSUBS 0.026647f
C1114 VDD2.n204 VSUBS 0.014319f
C1115 VDD2.n205 VSUBS 0.015161f
C1116 VDD2.n206 VSUBS 0.033845f
C1117 VDD2.n207 VSUBS 0.033845f
C1118 VDD2.n208 VSUBS 0.015161f
C1119 VDD2.n209 VSUBS 0.014319f
C1120 VDD2.n210 VSUBS 0.026647f
C1121 VDD2.n211 VSUBS 0.026647f
C1122 VDD2.n212 VSUBS 0.014319f
C1123 VDD2.n213 VSUBS 0.015161f
C1124 VDD2.n214 VSUBS 0.033845f
C1125 VDD2.n215 VSUBS 0.084633f
C1126 VDD2.n216 VSUBS 0.015161f
C1127 VDD2.n217 VSUBS 0.014319f
C1128 VDD2.n218 VSUBS 0.061593f
C1129 VDD2.n219 VSUBS 0.06108f
C1130 VDD2.n220 VSUBS 3.2327f
C1131 VDD2.t4 VSUBS 0.414406f
C1132 VDD2.t2 VSUBS 0.414406f
C1133 VDD2.n221 VSUBS 3.48312f
C1134 VN.n0 VSUBS 0.039248f
C1135 VN.t2 VSUBS 3.51884f
C1136 VN.n1 VSUBS 0.024055f
C1137 VN.n2 VSUBS 0.252683f
C1138 VN.t4 VSUBS 3.51884f
C1139 VN.t5 VSUBS 3.69649f
C1140 VN.n3 VSUBS 1.28861f
C1141 VN.n4 VSUBS 1.29634f
C1142 VN.n5 VSUBS 0.041581f
C1143 VN.n6 VSUBS 0.059001f
C1144 VN.n7 VSUBS 0.029771f
C1145 VN.n8 VSUBS 0.029771f
C1146 VN.n9 VSUBS 0.029771f
C1147 VN.n10 VSUBS 0.058706f
C1148 VN.n11 VSUBS 0.042126f
C1149 VN.n12 VSUBS 1.30697f
C1150 VN.n13 VSUBS 0.042767f
C1151 VN.n14 VSUBS 0.039248f
C1152 VN.t0 VSUBS 3.51884f
C1153 VN.n15 VSUBS 0.024055f
C1154 VN.n16 VSUBS 0.252683f
C1155 VN.t1 VSUBS 3.51884f
C1156 VN.t3 VSUBS 3.69649f
C1157 VN.n17 VSUBS 1.28861f
C1158 VN.n18 VSUBS 1.29634f
C1159 VN.n19 VSUBS 0.041581f
C1160 VN.n20 VSUBS 0.059001f
C1161 VN.n21 VSUBS 0.029771f
C1162 VN.n22 VSUBS 0.029771f
C1163 VN.n23 VSUBS 0.029771f
C1164 VN.n24 VSUBS 0.058706f
C1165 VN.n25 VSUBS 0.042126f
C1166 VN.n26 VSUBS 1.30697f
C1167 VN.n27 VSUBS 1.80197f
C1168 VDD1.n0 VSUBS 0.030186f
C1169 VDD1.n1 VSUBS 0.026749f
C1170 VDD1.n2 VSUBS 0.014374f
C1171 VDD1.n3 VSUBS 0.033974f
C1172 VDD1.n4 VSUBS 0.015219f
C1173 VDD1.n5 VSUBS 0.026749f
C1174 VDD1.n6 VSUBS 0.014374f
C1175 VDD1.n7 VSUBS 0.033974f
C1176 VDD1.n8 VSUBS 0.015219f
C1177 VDD1.n9 VSUBS 0.026749f
C1178 VDD1.n10 VSUBS 0.014374f
C1179 VDD1.n11 VSUBS 0.033974f
C1180 VDD1.n12 VSUBS 0.014796f
C1181 VDD1.n13 VSUBS 0.026749f
C1182 VDD1.n14 VSUBS 0.014796f
C1183 VDD1.n15 VSUBS 0.014374f
C1184 VDD1.n16 VSUBS 0.033974f
C1185 VDD1.n17 VSUBS 0.033974f
C1186 VDD1.n18 VSUBS 0.015219f
C1187 VDD1.n19 VSUBS 0.026749f
C1188 VDD1.n20 VSUBS 0.014374f
C1189 VDD1.n21 VSUBS 0.033974f
C1190 VDD1.n22 VSUBS 0.015219f
C1191 VDD1.n23 VSUBS 0.026749f
C1192 VDD1.n24 VSUBS 0.014374f
C1193 VDD1.n25 VSUBS 0.033974f
C1194 VDD1.n26 VSUBS 0.015219f
C1195 VDD1.n27 VSUBS 0.026749f
C1196 VDD1.n28 VSUBS 0.014374f
C1197 VDD1.n29 VSUBS 0.033974f
C1198 VDD1.n30 VSUBS 0.015219f
C1199 VDD1.n31 VSUBS 0.026749f
C1200 VDD1.n32 VSUBS 0.014374f
C1201 VDD1.n33 VSUBS 0.033974f
C1202 VDD1.n34 VSUBS 0.015219f
C1203 VDD1.n35 VSUBS 2.27626f
C1204 VDD1.n36 VSUBS 0.014374f
C1205 VDD1.t0 VSUBS 0.073043f
C1206 VDD1.n37 VSUBS 0.225479f
C1207 VDD1.n38 VSUBS 0.021613f
C1208 VDD1.n39 VSUBS 0.02548f
C1209 VDD1.n40 VSUBS 0.033974f
C1210 VDD1.n41 VSUBS 0.015219f
C1211 VDD1.n42 VSUBS 0.014374f
C1212 VDD1.n43 VSUBS 0.026749f
C1213 VDD1.n44 VSUBS 0.026749f
C1214 VDD1.n45 VSUBS 0.014374f
C1215 VDD1.n46 VSUBS 0.015219f
C1216 VDD1.n47 VSUBS 0.033974f
C1217 VDD1.n48 VSUBS 0.033974f
C1218 VDD1.n49 VSUBS 0.015219f
C1219 VDD1.n50 VSUBS 0.014374f
C1220 VDD1.n51 VSUBS 0.026749f
C1221 VDD1.n52 VSUBS 0.026749f
C1222 VDD1.n53 VSUBS 0.014374f
C1223 VDD1.n54 VSUBS 0.015219f
C1224 VDD1.n55 VSUBS 0.033974f
C1225 VDD1.n56 VSUBS 0.033974f
C1226 VDD1.n57 VSUBS 0.015219f
C1227 VDD1.n58 VSUBS 0.014374f
C1228 VDD1.n59 VSUBS 0.026749f
C1229 VDD1.n60 VSUBS 0.026749f
C1230 VDD1.n61 VSUBS 0.014374f
C1231 VDD1.n62 VSUBS 0.015219f
C1232 VDD1.n63 VSUBS 0.033974f
C1233 VDD1.n64 VSUBS 0.033974f
C1234 VDD1.n65 VSUBS 0.015219f
C1235 VDD1.n66 VSUBS 0.014374f
C1236 VDD1.n67 VSUBS 0.026749f
C1237 VDD1.n68 VSUBS 0.026749f
C1238 VDD1.n69 VSUBS 0.014374f
C1239 VDD1.n70 VSUBS 0.015219f
C1240 VDD1.n71 VSUBS 0.033974f
C1241 VDD1.n72 VSUBS 0.033974f
C1242 VDD1.n73 VSUBS 0.015219f
C1243 VDD1.n74 VSUBS 0.014374f
C1244 VDD1.n75 VSUBS 0.026749f
C1245 VDD1.n76 VSUBS 0.026749f
C1246 VDD1.n77 VSUBS 0.014374f
C1247 VDD1.n78 VSUBS 0.015219f
C1248 VDD1.n79 VSUBS 0.033974f
C1249 VDD1.n80 VSUBS 0.033974f
C1250 VDD1.n81 VSUBS 0.015219f
C1251 VDD1.n82 VSUBS 0.014374f
C1252 VDD1.n83 VSUBS 0.026749f
C1253 VDD1.n84 VSUBS 0.026749f
C1254 VDD1.n85 VSUBS 0.014374f
C1255 VDD1.n86 VSUBS 0.015219f
C1256 VDD1.n87 VSUBS 0.033974f
C1257 VDD1.n88 VSUBS 0.033974f
C1258 VDD1.n89 VSUBS 0.015219f
C1259 VDD1.n90 VSUBS 0.014374f
C1260 VDD1.n91 VSUBS 0.026749f
C1261 VDD1.n92 VSUBS 0.026749f
C1262 VDD1.n93 VSUBS 0.014374f
C1263 VDD1.n94 VSUBS 0.015219f
C1264 VDD1.n95 VSUBS 0.033974f
C1265 VDD1.n96 VSUBS 0.033974f
C1266 VDD1.n97 VSUBS 0.015219f
C1267 VDD1.n98 VSUBS 0.014374f
C1268 VDD1.n99 VSUBS 0.026749f
C1269 VDD1.n100 VSUBS 0.026749f
C1270 VDD1.n101 VSUBS 0.014374f
C1271 VDD1.n102 VSUBS 0.015219f
C1272 VDD1.n103 VSUBS 0.033974f
C1273 VDD1.n104 VSUBS 0.084956f
C1274 VDD1.n105 VSUBS 0.015219f
C1275 VDD1.n106 VSUBS 0.014374f
C1276 VDD1.n107 VSUBS 0.061828f
C1277 VDD1.n108 VSUBS 0.067845f
C1278 VDD1.n109 VSUBS 0.030186f
C1279 VDD1.n110 VSUBS 0.026749f
C1280 VDD1.n111 VSUBS 0.014374f
C1281 VDD1.n112 VSUBS 0.033974f
C1282 VDD1.n113 VSUBS 0.015219f
C1283 VDD1.n114 VSUBS 0.026749f
C1284 VDD1.n115 VSUBS 0.014374f
C1285 VDD1.n116 VSUBS 0.033974f
C1286 VDD1.n117 VSUBS 0.015219f
C1287 VDD1.n118 VSUBS 0.026749f
C1288 VDD1.n119 VSUBS 0.014374f
C1289 VDD1.n120 VSUBS 0.033974f
C1290 VDD1.n121 VSUBS 0.014796f
C1291 VDD1.n122 VSUBS 0.026749f
C1292 VDD1.n123 VSUBS 0.015219f
C1293 VDD1.n124 VSUBS 0.033974f
C1294 VDD1.n125 VSUBS 0.015219f
C1295 VDD1.n126 VSUBS 0.026749f
C1296 VDD1.n127 VSUBS 0.014374f
C1297 VDD1.n128 VSUBS 0.033974f
C1298 VDD1.n129 VSUBS 0.015219f
C1299 VDD1.n130 VSUBS 0.026749f
C1300 VDD1.n131 VSUBS 0.014374f
C1301 VDD1.n132 VSUBS 0.033974f
C1302 VDD1.n133 VSUBS 0.015219f
C1303 VDD1.n134 VSUBS 0.026749f
C1304 VDD1.n135 VSUBS 0.014374f
C1305 VDD1.n136 VSUBS 0.033974f
C1306 VDD1.n137 VSUBS 0.015219f
C1307 VDD1.n138 VSUBS 0.026749f
C1308 VDD1.n139 VSUBS 0.014374f
C1309 VDD1.n140 VSUBS 0.033974f
C1310 VDD1.n141 VSUBS 0.015219f
C1311 VDD1.n142 VSUBS 2.27626f
C1312 VDD1.n143 VSUBS 0.014374f
C1313 VDD1.t5 VSUBS 0.073043f
C1314 VDD1.n144 VSUBS 0.225479f
C1315 VDD1.n145 VSUBS 0.021613f
C1316 VDD1.n146 VSUBS 0.02548f
C1317 VDD1.n147 VSUBS 0.033974f
C1318 VDD1.n148 VSUBS 0.015219f
C1319 VDD1.n149 VSUBS 0.014374f
C1320 VDD1.n150 VSUBS 0.026749f
C1321 VDD1.n151 VSUBS 0.026749f
C1322 VDD1.n152 VSUBS 0.014374f
C1323 VDD1.n153 VSUBS 0.015219f
C1324 VDD1.n154 VSUBS 0.033974f
C1325 VDD1.n155 VSUBS 0.033974f
C1326 VDD1.n156 VSUBS 0.015219f
C1327 VDD1.n157 VSUBS 0.014374f
C1328 VDD1.n158 VSUBS 0.026749f
C1329 VDD1.n159 VSUBS 0.026749f
C1330 VDD1.n160 VSUBS 0.014374f
C1331 VDD1.n161 VSUBS 0.015219f
C1332 VDD1.n162 VSUBS 0.033974f
C1333 VDD1.n163 VSUBS 0.033974f
C1334 VDD1.n164 VSUBS 0.015219f
C1335 VDD1.n165 VSUBS 0.014374f
C1336 VDD1.n166 VSUBS 0.026749f
C1337 VDD1.n167 VSUBS 0.026749f
C1338 VDD1.n168 VSUBS 0.014374f
C1339 VDD1.n169 VSUBS 0.015219f
C1340 VDD1.n170 VSUBS 0.033974f
C1341 VDD1.n171 VSUBS 0.033974f
C1342 VDD1.n172 VSUBS 0.015219f
C1343 VDD1.n173 VSUBS 0.014374f
C1344 VDD1.n174 VSUBS 0.026749f
C1345 VDD1.n175 VSUBS 0.026749f
C1346 VDD1.n176 VSUBS 0.014374f
C1347 VDD1.n177 VSUBS 0.015219f
C1348 VDD1.n178 VSUBS 0.033974f
C1349 VDD1.n179 VSUBS 0.033974f
C1350 VDD1.n180 VSUBS 0.015219f
C1351 VDD1.n181 VSUBS 0.014374f
C1352 VDD1.n182 VSUBS 0.026749f
C1353 VDD1.n183 VSUBS 0.026749f
C1354 VDD1.n184 VSUBS 0.014374f
C1355 VDD1.n185 VSUBS 0.014374f
C1356 VDD1.n186 VSUBS 0.015219f
C1357 VDD1.n187 VSUBS 0.033974f
C1358 VDD1.n188 VSUBS 0.033974f
C1359 VDD1.n189 VSUBS 0.033974f
C1360 VDD1.n190 VSUBS 0.014796f
C1361 VDD1.n191 VSUBS 0.014374f
C1362 VDD1.n192 VSUBS 0.026749f
C1363 VDD1.n193 VSUBS 0.026749f
C1364 VDD1.n194 VSUBS 0.014374f
C1365 VDD1.n195 VSUBS 0.015219f
C1366 VDD1.n196 VSUBS 0.033974f
C1367 VDD1.n197 VSUBS 0.033974f
C1368 VDD1.n198 VSUBS 0.015219f
C1369 VDD1.n199 VSUBS 0.014374f
C1370 VDD1.n200 VSUBS 0.026749f
C1371 VDD1.n201 VSUBS 0.026749f
C1372 VDD1.n202 VSUBS 0.014374f
C1373 VDD1.n203 VSUBS 0.015219f
C1374 VDD1.n204 VSUBS 0.033974f
C1375 VDD1.n205 VSUBS 0.033974f
C1376 VDD1.n206 VSUBS 0.015219f
C1377 VDD1.n207 VSUBS 0.014374f
C1378 VDD1.n208 VSUBS 0.026749f
C1379 VDD1.n209 VSUBS 0.026749f
C1380 VDD1.n210 VSUBS 0.014374f
C1381 VDD1.n211 VSUBS 0.015219f
C1382 VDD1.n212 VSUBS 0.033974f
C1383 VDD1.n213 VSUBS 0.084956f
C1384 VDD1.n214 VSUBS 0.015219f
C1385 VDD1.n215 VSUBS 0.014374f
C1386 VDD1.n216 VSUBS 0.061828f
C1387 VDD1.n217 VSUBS 0.067126f
C1388 VDD1.t2 VSUBS 0.415988f
C1389 VDD1.t1 VSUBS 0.415988f
C1390 VDD1.n218 VSUBS 3.49647f
C1391 VDD1.n219 VSUBS 3.6241f
C1392 VDD1.t3 VSUBS 0.415988f
C1393 VDD1.t4 VSUBS 0.415988f
C1394 VDD1.n220 VSUBS 3.49098f
C1395 VDD1.n221 VSUBS 3.79573f
C1396 VTAIL.t0 VSUBS 0.420679f
C1397 VTAIL.t1 VSUBS 0.420679f
C1398 VTAIL.n0 VSUBS 3.35647f
C1399 VTAIL.n1 VSUBS 0.865899f
C1400 VTAIL.n2 VSUBS 0.030527f
C1401 VTAIL.n3 VSUBS 0.02705f
C1402 VTAIL.n4 VSUBS 0.014536f
C1403 VTAIL.n5 VSUBS 0.034357f
C1404 VTAIL.n6 VSUBS 0.015391f
C1405 VTAIL.n7 VSUBS 0.02705f
C1406 VTAIL.n8 VSUBS 0.014536f
C1407 VTAIL.n9 VSUBS 0.034357f
C1408 VTAIL.n10 VSUBS 0.015391f
C1409 VTAIL.n11 VSUBS 0.02705f
C1410 VTAIL.n12 VSUBS 0.014536f
C1411 VTAIL.n13 VSUBS 0.034357f
C1412 VTAIL.n14 VSUBS 0.014963f
C1413 VTAIL.n15 VSUBS 0.02705f
C1414 VTAIL.n16 VSUBS 0.015391f
C1415 VTAIL.n17 VSUBS 0.034357f
C1416 VTAIL.n18 VSUBS 0.015391f
C1417 VTAIL.n19 VSUBS 0.02705f
C1418 VTAIL.n20 VSUBS 0.014536f
C1419 VTAIL.n21 VSUBS 0.034357f
C1420 VTAIL.n22 VSUBS 0.015391f
C1421 VTAIL.n23 VSUBS 0.02705f
C1422 VTAIL.n24 VSUBS 0.014536f
C1423 VTAIL.n25 VSUBS 0.034357f
C1424 VTAIL.n26 VSUBS 0.015391f
C1425 VTAIL.n27 VSUBS 0.02705f
C1426 VTAIL.n28 VSUBS 0.014536f
C1427 VTAIL.n29 VSUBS 0.034357f
C1428 VTAIL.n30 VSUBS 0.015391f
C1429 VTAIL.n31 VSUBS 0.02705f
C1430 VTAIL.n32 VSUBS 0.014536f
C1431 VTAIL.n33 VSUBS 0.034357f
C1432 VTAIL.n34 VSUBS 0.015391f
C1433 VTAIL.n35 VSUBS 2.30193f
C1434 VTAIL.n36 VSUBS 0.014536f
C1435 VTAIL.t11 VSUBS 0.073866f
C1436 VTAIL.n37 VSUBS 0.228022f
C1437 VTAIL.n38 VSUBS 0.021856f
C1438 VTAIL.n39 VSUBS 0.025768f
C1439 VTAIL.n40 VSUBS 0.034357f
C1440 VTAIL.n41 VSUBS 0.015391f
C1441 VTAIL.n42 VSUBS 0.014536f
C1442 VTAIL.n43 VSUBS 0.02705f
C1443 VTAIL.n44 VSUBS 0.02705f
C1444 VTAIL.n45 VSUBS 0.014536f
C1445 VTAIL.n46 VSUBS 0.015391f
C1446 VTAIL.n47 VSUBS 0.034357f
C1447 VTAIL.n48 VSUBS 0.034357f
C1448 VTAIL.n49 VSUBS 0.015391f
C1449 VTAIL.n50 VSUBS 0.014536f
C1450 VTAIL.n51 VSUBS 0.02705f
C1451 VTAIL.n52 VSUBS 0.02705f
C1452 VTAIL.n53 VSUBS 0.014536f
C1453 VTAIL.n54 VSUBS 0.015391f
C1454 VTAIL.n55 VSUBS 0.034357f
C1455 VTAIL.n56 VSUBS 0.034357f
C1456 VTAIL.n57 VSUBS 0.015391f
C1457 VTAIL.n58 VSUBS 0.014536f
C1458 VTAIL.n59 VSUBS 0.02705f
C1459 VTAIL.n60 VSUBS 0.02705f
C1460 VTAIL.n61 VSUBS 0.014536f
C1461 VTAIL.n62 VSUBS 0.015391f
C1462 VTAIL.n63 VSUBS 0.034357f
C1463 VTAIL.n64 VSUBS 0.034357f
C1464 VTAIL.n65 VSUBS 0.015391f
C1465 VTAIL.n66 VSUBS 0.014536f
C1466 VTAIL.n67 VSUBS 0.02705f
C1467 VTAIL.n68 VSUBS 0.02705f
C1468 VTAIL.n69 VSUBS 0.014536f
C1469 VTAIL.n70 VSUBS 0.015391f
C1470 VTAIL.n71 VSUBS 0.034357f
C1471 VTAIL.n72 VSUBS 0.034357f
C1472 VTAIL.n73 VSUBS 0.015391f
C1473 VTAIL.n74 VSUBS 0.014536f
C1474 VTAIL.n75 VSUBS 0.02705f
C1475 VTAIL.n76 VSUBS 0.02705f
C1476 VTAIL.n77 VSUBS 0.014536f
C1477 VTAIL.n78 VSUBS 0.014536f
C1478 VTAIL.n79 VSUBS 0.015391f
C1479 VTAIL.n80 VSUBS 0.034357f
C1480 VTAIL.n81 VSUBS 0.034357f
C1481 VTAIL.n82 VSUBS 0.034357f
C1482 VTAIL.n83 VSUBS 0.014963f
C1483 VTAIL.n84 VSUBS 0.014536f
C1484 VTAIL.n85 VSUBS 0.02705f
C1485 VTAIL.n86 VSUBS 0.02705f
C1486 VTAIL.n87 VSUBS 0.014536f
C1487 VTAIL.n88 VSUBS 0.015391f
C1488 VTAIL.n89 VSUBS 0.034357f
C1489 VTAIL.n90 VSUBS 0.034357f
C1490 VTAIL.n91 VSUBS 0.015391f
C1491 VTAIL.n92 VSUBS 0.014536f
C1492 VTAIL.n93 VSUBS 0.02705f
C1493 VTAIL.n94 VSUBS 0.02705f
C1494 VTAIL.n95 VSUBS 0.014536f
C1495 VTAIL.n96 VSUBS 0.015391f
C1496 VTAIL.n97 VSUBS 0.034357f
C1497 VTAIL.n98 VSUBS 0.034357f
C1498 VTAIL.n99 VSUBS 0.015391f
C1499 VTAIL.n100 VSUBS 0.014536f
C1500 VTAIL.n101 VSUBS 0.02705f
C1501 VTAIL.n102 VSUBS 0.02705f
C1502 VTAIL.n103 VSUBS 0.014536f
C1503 VTAIL.n104 VSUBS 0.015391f
C1504 VTAIL.n105 VSUBS 0.034357f
C1505 VTAIL.n106 VSUBS 0.085914f
C1506 VTAIL.n107 VSUBS 0.015391f
C1507 VTAIL.n108 VSUBS 0.014536f
C1508 VTAIL.n109 VSUBS 0.062526f
C1509 VTAIL.n110 VSUBS 0.043327f
C1510 VTAIL.n111 VSUBS 0.346955f
C1511 VTAIL.t6 VSUBS 0.420679f
C1512 VTAIL.t9 VSUBS 0.420679f
C1513 VTAIL.n112 VSUBS 3.35647f
C1514 VTAIL.n113 VSUBS 3.09043f
C1515 VTAIL.t2 VSUBS 0.420679f
C1516 VTAIL.t3 VSUBS 0.420679f
C1517 VTAIL.n114 VSUBS 3.35649f
C1518 VTAIL.n115 VSUBS 3.09041f
C1519 VTAIL.n116 VSUBS 0.030527f
C1520 VTAIL.n117 VSUBS 0.02705f
C1521 VTAIL.n118 VSUBS 0.014536f
C1522 VTAIL.n119 VSUBS 0.034357f
C1523 VTAIL.n120 VSUBS 0.015391f
C1524 VTAIL.n121 VSUBS 0.02705f
C1525 VTAIL.n122 VSUBS 0.014536f
C1526 VTAIL.n123 VSUBS 0.034357f
C1527 VTAIL.n124 VSUBS 0.015391f
C1528 VTAIL.n125 VSUBS 0.02705f
C1529 VTAIL.n126 VSUBS 0.014536f
C1530 VTAIL.n127 VSUBS 0.034357f
C1531 VTAIL.n128 VSUBS 0.014963f
C1532 VTAIL.n129 VSUBS 0.02705f
C1533 VTAIL.n130 VSUBS 0.014963f
C1534 VTAIL.n131 VSUBS 0.014536f
C1535 VTAIL.n132 VSUBS 0.034357f
C1536 VTAIL.n133 VSUBS 0.034357f
C1537 VTAIL.n134 VSUBS 0.015391f
C1538 VTAIL.n135 VSUBS 0.02705f
C1539 VTAIL.n136 VSUBS 0.014536f
C1540 VTAIL.n137 VSUBS 0.034357f
C1541 VTAIL.n138 VSUBS 0.015391f
C1542 VTAIL.n139 VSUBS 0.02705f
C1543 VTAIL.n140 VSUBS 0.014536f
C1544 VTAIL.n141 VSUBS 0.034357f
C1545 VTAIL.n142 VSUBS 0.015391f
C1546 VTAIL.n143 VSUBS 0.02705f
C1547 VTAIL.n144 VSUBS 0.014536f
C1548 VTAIL.n145 VSUBS 0.034357f
C1549 VTAIL.n146 VSUBS 0.015391f
C1550 VTAIL.n147 VSUBS 0.02705f
C1551 VTAIL.n148 VSUBS 0.014536f
C1552 VTAIL.n149 VSUBS 0.034357f
C1553 VTAIL.n150 VSUBS 0.015391f
C1554 VTAIL.n151 VSUBS 2.30193f
C1555 VTAIL.n152 VSUBS 0.014536f
C1556 VTAIL.t4 VSUBS 0.073866f
C1557 VTAIL.n153 VSUBS 0.228022f
C1558 VTAIL.n154 VSUBS 0.021856f
C1559 VTAIL.n155 VSUBS 0.025768f
C1560 VTAIL.n156 VSUBS 0.034357f
C1561 VTAIL.n157 VSUBS 0.015391f
C1562 VTAIL.n158 VSUBS 0.014536f
C1563 VTAIL.n159 VSUBS 0.02705f
C1564 VTAIL.n160 VSUBS 0.02705f
C1565 VTAIL.n161 VSUBS 0.014536f
C1566 VTAIL.n162 VSUBS 0.015391f
C1567 VTAIL.n163 VSUBS 0.034357f
C1568 VTAIL.n164 VSUBS 0.034357f
C1569 VTAIL.n165 VSUBS 0.015391f
C1570 VTAIL.n166 VSUBS 0.014536f
C1571 VTAIL.n167 VSUBS 0.02705f
C1572 VTAIL.n168 VSUBS 0.02705f
C1573 VTAIL.n169 VSUBS 0.014536f
C1574 VTAIL.n170 VSUBS 0.015391f
C1575 VTAIL.n171 VSUBS 0.034357f
C1576 VTAIL.n172 VSUBS 0.034357f
C1577 VTAIL.n173 VSUBS 0.015391f
C1578 VTAIL.n174 VSUBS 0.014536f
C1579 VTAIL.n175 VSUBS 0.02705f
C1580 VTAIL.n176 VSUBS 0.02705f
C1581 VTAIL.n177 VSUBS 0.014536f
C1582 VTAIL.n178 VSUBS 0.015391f
C1583 VTAIL.n179 VSUBS 0.034357f
C1584 VTAIL.n180 VSUBS 0.034357f
C1585 VTAIL.n181 VSUBS 0.015391f
C1586 VTAIL.n182 VSUBS 0.014536f
C1587 VTAIL.n183 VSUBS 0.02705f
C1588 VTAIL.n184 VSUBS 0.02705f
C1589 VTAIL.n185 VSUBS 0.014536f
C1590 VTAIL.n186 VSUBS 0.015391f
C1591 VTAIL.n187 VSUBS 0.034357f
C1592 VTAIL.n188 VSUBS 0.034357f
C1593 VTAIL.n189 VSUBS 0.015391f
C1594 VTAIL.n190 VSUBS 0.014536f
C1595 VTAIL.n191 VSUBS 0.02705f
C1596 VTAIL.n192 VSUBS 0.02705f
C1597 VTAIL.n193 VSUBS 0.014536f
C1598 VTAIL.n194 VSUBS 0.015391f
C1599 VTAIL.n195 VSUBS 0.034357f
C1600 VTAIL.n196 VSUBS 0.034357f
C1601 VTAIL.n197 VSUBS 0.015391f
C1602 VTAIL.n198 VSUBS 0.014536f
C1603 VTAIL.n199 VSUBS 0.02705f
C1604 VTAIL.n200 VSUBS 0.02705f
C1605 VTAIL.n201 VSUBS 0.014536f
C1606 VTAIL.n202 VSUBS 0.015391f
C1607 VTAIL.n203 VSUBS 0.034357f
C1608 VTAIL.n204 VSUBS 0.034357f
C1609 VTAIL.n205 VSUBS 0.015391f
C1610 VTAIL.n206 VSUBS 0.014536f
C1611 VTAIL.n207 VSUBS 0.02705f
C1612 VTAIL.n208 VSUBS 0.02705f
C1613 VTAIL.n209 VSUBS 0.014536f
C1614 VTAIL.n210 VSUBS 0.015391f
C1615 VTAIL.n211 VSUBS 0.034357f
C1616 VTAIL.n212 VSUBS 0.034357f
C1617 VTAIL.n213 VSUBS 0.015391f
C1618 VTAIL.n214 VSUBS 0.014536f
C1619 VTAIL.n215 VSUBS 0.02705f
C1620 VTAIL.n216 VSUBS 0.02705f
C1621 VTAIL.n217 VSUBS 0.014536f
C1622 VTAIL.n218 VSUBS 0.015391f
C1623 VTAIL.n219 VSUBS 0.034357f
C1624 VTAIL.n220 VSUBS 0.085914f
C1625 VTAIL.n221 VSUBS 0.015391f
C1626 VTAIL.n222 VSUBS 0.014536f
C1627 VTAIL.n223 VSUBS 0.062526f
C1628 VTAIL.n224 VSUBS 0.043327f
C1629 VTAIL.n225 VSUBS 0.346955f
C1630 VTAIL.t10 VSUBS 0.420679f
C1631 VTAIL.t8 VSUBS 0.420679f
C1632 VTAIL.n226 VSUBS 3.35649f
C1633 VTAIL.n227 VSUBS 1.00226f
C1634 VTAIL.n228 VSUBS 0.030527f
C1635 VTAIL.n229 VSUBS 0.02705f
C1636 VTAIL.n230 VSUBS 0.014536f
C1637 VTAIL.n231 VSUBS 0.034357f
C1638 VTAIL.n232 VSUBS 0.015391f
C1639 VTAIL.n233 VSUBS 0.02705f
C1640 VTAIL.n234 VSUBS 0.014536f
C1641 VTAIL.n235 VSUBS 0.034357f
C1642 VTAIL.n236 VSUBS 0.015391f
C1643 VTAIL.n237 VSUBS 0.02705f
C1644 VTAIL.n238 VSUBS 0.014536f
C1645 VTAIL.n239 VSUBS 0.034357f
C1646 VTAIL.n240 VSUBS 0.014963f
C1647 VTAIL.n241 VSUBS 0.02705f
C1648 VTAIL.n242 VSUBS 0.014963f
C1649 VTAIL.n243 VSUBS 0.014536f
C1650 VTAIL.n244 VSUBS 0.034357f
C1651 VTAIL.n245 VSUBS 0.034357f
C1652 VTAIL.n246 VSUBS 0.015391f
C1653 VTAIL.n247 VSUBS 0.02705f
C1654 VTAIL.n248 VSUBS 0.014536f
C1655 VTAIL.n249 VSUBS 0.034357f
C1656 VTAIL.n250 VSUBS 0.015391f
C1657 VTAIL.n251 VSUBS 0.02705f
C1658 VTAIL.n252 VSUBS 0.014536f
C1659 VTAIL.n253 VSUBS 0.034357f
C1660 VTAIL.n254 VSUBS 0.015391f
C1661 VTAIL.n255 VSUBS 0.02705f
C1662 VTAIL.n256 VSUBS 0.014536f
C1663 VTAIL.n257 VSUBS 0.034357f
C1664 VTAIL.n258 VSUBS 0.015391f
C1665 VTAIL.n259 VSUBS 0.02705f
C1666 VTAIL.n260 VSUBS 0.014536f
C1667 VTAIL.n261 VSUBS 0.034357f
C1668 VTAIL.n262 VSUBS 0.015391f
C1669 VTAIL.n263 VSUBS 2.30193f
C1670 VTAIL.n264 VSUBS 0.014536f
C1671 VTAIL.t7 VSUBS 0.073866f
C1672 VTAIL.n265 VSUBS 0.228022f
C1673 VTAIL.n266 VSUBS 0.021856f
C1674 VTAIL.n267 VSUBS 0.025768f
C1675 VTAIL.n268 VSUBS 0.034357f
C1676 VTAIL.n269 VSUBS 0.015391f
C1677 VTAIL.n270 VSUBS 0.014536f
C1678 VTAIL.n271 VSUBS 0.02705f
C1679 VTAIL.n272 VSUBS 0.02705f
C1680 VTAIL.n273 VSUBS 0.014536f
C1681 VTAIL.n274 VSUBS 0.015391f
C1682 VTAIL.n275 VSUBS 0.034357f
C1683 VTAIL.n276 VSUBS 0.034357f
C1684 VTAIL.n277 VSUBS 0.015391f
C1685 VTAIL.n278 VSUBS 0.014536f
C1686 VTAIL.n279 VSUBS 0.02705f
C1687 VTAIL.n280 VSUBS 0.02705f
C1688 VTAIL.n281 VSUBS 0.014536f
C1689 VTAIL.n282 VSUBS 0.015391f
C1690 VTAIL.n283 VSUBS 0.034357f
C1691 VTAIL.n284 VSUBS 0.034357f
C1692 VTAIL.n285 VSUBS 0.015391f
C1693 VTAIL.n286 VSUBS 0.014536f
C1694 VTAIL.n287 VSUBS 0.02705f
C1695 VTAIL.n288 VSUBS 0.02705f
C1696 VTAIL.n289 VSUBS 0.014536f
C1697 VTAIL.n290 VSUBS 0.015391f
C1698 VTAIL.n291 VSUBS 0.034357f
C1699 VTAIL.n292 VSUBS 0.034357f
C1700 VTAIL.n293 VSUBS 0.015391f
C1701 VTAIL.n294 VSUBS 0.014536f
C1702 VTAIL.n295 VSUBS 0.02705f
C1703 VTAIL.n296 VSUBS 0.02705f
C1704 VTAIL.n297 VSUBS 0.014536f
C1705 VTAIL.n298 VSUBS 0.015391f
C1706 VTAIL.n299 VSUBS 0.034357f
C1707 VTAIL.n300 VSUBS 0.034357f
C1708 VTAIL.n301 VSUBS 0.015391f
C1709 VTAIL.n302 VSUBS 0.014536f
C1710 VTAIL.n303 VSUBS 0.02705f
C1711 VTAIL.n304 VSUBS 0.02705f
C1712 VTAIL.n305 VSUBS 0.014536f
C1713 VTAIL.n306 VSUBS 0.015391f
C1714 VTAIL.n307 VSUBS 0.034357f
C1715 VTAIL.n308 VSUBS 0.034357f
C1716 VTAIL.n309 VSUBS 0.015391f
C1717 VTAIL.n310 VSUBS 0.014536f
C1718 VTAIL.n311 VSUBS 0.02705f
C1719 VTAIL.n312 VSUBS 0.02705f
C1720 VTAIL.n313 VSUBS 0.014536f
C1721 VTAIL.n314 VSUBS 0.015391f
C1722 VTAIL.n315 VSUBS 0.034357f
C1723 VTAIL.n316 VSUBS 0.034357f
C1724 VTAIL.n317 VSUBS 0.015391f
C1725 VTAIL.n318 VSUBS 0.014536f
C1726 VTAIL.n319 VSUBS 0.02705f
C1727 VTAIL.n320 VSUBS 0.02705f
C1728 VTAIL.n321 VSUBS 0.014536f
C1729 VTAIL.n322 VSUBS 0.015391f
C1730 VTAIL.n323 VSUBS 0.034357f
C1731 VTAIL.n324 VSUBS 0.034357f
C1732 VTAIL.n325 VSUBS 0.015391f
C1733 VTAIL.n326 VSUBS 0.014536f
C1734 VTAIL.n327 VSUBS 0.02705f
C1735 VTAIL.n328 VSUBS 0.02705f
C1736 VTAIL.n329 VSUBS 0.014536f
C1737 VTAIL.n330 VSUBS 0.015391f
C1738 VTAIL.n331 VSUBS 0.034357f
C1739 VTAIL.n332 VSUBS 0.085914f
C1740 VTAIL.n333 VSUBS 0.015391f
C1741 VTAIL.n334 VSUBS 0.014536f
C1742 VTAIL.n335 VSUBS 0.062526f
C1743 VTAIL.n336 VSUBS 0.043327f
C1744 VTAIL.n337 VSUBS 2.2465f
C1745 VTAIL.n338 VSUBS 0.030527f
C1746 VTAIL.n339 VSUBS 0.02705f
C1747 VTAIL.n340 VSUBS 0.014536f
C1748 VTAIL.n341 VSUBS 0.034357f
C1749 VTAIL.n342 VSUBS 0.015391f
C1750 VTAIL.n343 VSUBS 0.02705f
C1751 VTAIL.n344 VSUBS 0.014536f
C1752 VTAIL.n345 VSUBS 0.034357f
C1753 VTAIL.n346 VSUBS 0.015391f
C1754 VTAIL.n347 VSUBS 0.02705f
C1755 VTAIL.n348 VSUBS 0.014536f
C1756 VTAIL.n349 VSUBS 0.034357f
C1757 VTAIL.n350 VSUBS 0.014963f
C1758 VTAIL.n351 VSUBS 0.02705f
C1759 VTAIL.n352 VSUBS 0.015391f
C1760 VTAIL.n353 VSUBS 0.034357f
C1761 VTAIL.n354 VSUBS 0.015391f
C1762 VTAIL.n355 VSUBS 0.02705f
C1763 VTAIL.n356 VSUBS 0.014536f
C1764 VTAIL.n357 VSUBS 0.034357f
C1765 VTAIL.n358 VSUBS 0.015391f
C1766 VTAIL.n359 VSUBS 0.02705f
C1767 VTAIL.n360 VSUBS 0.014536f
C1768 VTAIL.n361 VSUBS 0.034357f
C1769 VTAIL.n362 VSUBS 0.015391f
C1770 VTAIL.n363 VSUBS 0.02705f
C1771 VTAIL.n364 VSUBS 0.014536f
C1772 VTAIL.n365 VSUBS 0.034357f
C1773 VTAIL.n366 VSUBS 0.015391f
C1774 VTAIL.n367 VSUBS 0.02705f
C1775 VTAIL.n368 VSUBS 0.014536f
C1776 VTAIL.n369 VSUBS 0.034357f
C1777 VTAIL.n370 VSUBS 0.015391f
C1778 VTAIL.n371 VSUBS 2.30193f
C1779 VTAIL.n372 VSUBS 0.014536f
C1780 VTAIL.t5 VSUBS 0.073866f
C1781 VTAIL.n373 VSUBS 0.228022f
C1782 VTAIL.n374 VSUBS 0.021856f
C1783 VTAIL.n375 VSUBS 0.025768f
C1784 VTAIL.n376 VSUBS 0.034357f
C1785 VTAIL.n377 VSUBS 0.015391f
C1786 VTAIL.n378 VSUBS 0.014536f
C1787 VTAIL.n379 VSUBS 0.02705f
C1788 VTAIL.n380 VSUBS 0.02705f
C1789 VTAIL.n381 VSUBS 0.014536f
C1790 VTAIL.n382 VSUBS 0.015391f
C1791 VTAIL.n383 VSUBS 0.034357f
C1792 VTAIL.n384 VSUBS 0.034357f
C1793 VTAIL.n385 VSUBS 0.015391f
C1794 VTAIL.n386 VSUBS 0.014536f
C1795 VTAIL.n387 VSUBS 0.02705f
C1796 VTAIL.n388 VSUBS 0.02705f
C1797 VTAIL.n389 VSUBS 0.014536f
C1798 VTAIL.n390 VSUBS 0.015391f
C1799 VTAIL.n391 VSUBS 0.034357f
C1800 VTAIL.n392 VSUBS 0.034357f
C1801 VTAIL.n393 VSUBS 0.015391f
C1802 VTAIL.n394 VSUBS 0.014536f
C1803 VTAIL.n395 VSUBS 0.02705f
C1804 VTAIL.n396 VSUBS 0.02705f
C1805 VTAIL.n397 VSUBS 0.014536f
C1806 VTAIL.n398 VSUBS 0.015391f
C1807 VTAIL.n399 VSUBS 0.034357f
C1808 VTAIL.n400 VSUBS 0.034357f
C1809 VTAIL.n401 VSUBS 0.015391f
C1810 VTAIL.n402 VSUBS 0.014536f
C1811 VTAIL.n403 VSUBS 0.02705f
C1812 VTAIL.n404 VSUBS 0.02705f
C1813 VTAIL.n405 VSUBS 0.014536f
C1814 VTAIL.n406 VSUBS 0.015391f
C1815 VTAIL.n407 VSUBS 0.034357f
C1816 VTAIL.n408 VSUBS 0.034357f
C1817 VTAIL.n409 VSUBS 0.015391f
C1818 VTAIL.n410 VSUBS 0.014536f
C1819 VTAIL.n411 VSUBS 0.02705f
C1820 VTAIL.n412 VSUBS 0.02705f
C1821 VTAIL.n413 VSUBS 0.014536f
C1822 VTAIL.n414 VSUBS 0.014536f
C1823 VTAIL.n415 VSUBS 0.015391f
C1824 VTAIL.n416 VSUBS 0.034357f
C1825 VTAIL.n417 VSUBS 0.034357f
C1826 VTAIL.n418 VSUBS 0.034357f
C1827 VTAIL.n419 VSUBS 0.014963f
C1828 VTAIL.n420 VSUBS 0.014536f
C1829 VTAIL.n421 VSUBS 0.02705f
C1830 VTAIL.n422 VSUBS 0.02705f
C1831 VTAIL.n423 VSUBS 0.014536f
C1832 VTAIL.n424 VSUBS 0.015391f
C1833 VTAIL.n425 VSUBS 0.034357f
C1834 VTAIL.n426 VSUBS 0.034357f
C1835 VTAIL.n427 VSUBS 0.015391f
C1836 VTAIL.n428 VSUBS 0.014536f
C1837 VTAIL.n429 VSUBS 0.02705f
C1838 VTAIL.n430 VSUBS 0.02705f
C1839 VTAIL.n431 VSUBS 0.014536f
C1840 VTAIL.n432 VSUBS 0.015391f
C1841 VTAIL.n433 VSUBS 0.034357f
C1842 VTAIL.n434 VSUBS 0.034357f
C1843 VTAIL.n435 VSUBS 0.015391f
C1844 VTAIL.n436 VSUBS 0.014536f
C1845 VTAIL.n437 VSUBS 0.02705f
C1846 VTAIL.n438 VSUBS 0.02705f
C1847 VTAIL.n439 VSUBS 0.014536f
C1848 VTAIL.n440 VSUBS 0.015391f
C1849 VTAIL.n441 VSUBS 0.034357f
C1850 VTAIL.n442 VSUBS 0.085914f
C1851 VTAIL.n443 VSUBS 0.015391f
C1852 VTAIL.n444 VSUBS 0.014536f
C1853 VTAIL.n445 VSUBS 0.062526f
C1854 VTAIL.n446 VSUBS 0.043327f
C1855 VTAIL.n447 VSUBS 2.19428f
C1856 VP.n0 VSUBS 0.040103f
C1857 VP.t4 VSUBS 3.59549f
C1858 VP.n1 VSUBS 0.024579f
C1859 VP.n2 VSUBS 0.03042f
C1860 VP.t3 VSUBS 3.59549f
C1861 VP.n3 VSUBS 0.060286f
C1862 VP.n4 VSUBS 0.03042f
C1863 VP.t0 VSUBS 3.59549f
C1864 VP.n5 VSUBS 1.33544f
C1865 VP.n6 VSUBS 0.040103f
C1866 VP.t1 VSUBS 3.59549f
C1867 VP.n7 VSUBS 0.024579f
C1868 VP.n8 VSUBS 0.258187f
C1869 VP.t2 VSUBS 3.59549f
C1870 VP.t5 VSUBS 3.777f
C1871 VP.n9 VSUBS 1.31668f
C1872 VP.n10 VSUBS 1.32458f
C1873 VP.n11 VSUBS 0.042486f
C1874 VP.n12 VSUBS 0.060286f
C1875 VP.n13 VSUBS 0.03042f
C1876 VP.n14 VSUBS 0.03042f
C1877 VP.n15 VSUBS 0.03042f
C1878 VP.n16 VSUBS 0.059985f
C1879 VP.n17 VSUBS 0.043043f
C1880 VP.n18 VSUBS 1.33544f
C1881 VP.n19 VSUBS 1.82501f
C1882 VP.n20 VSUBS 1.84578f
C1883 VP.n21 VSUBS 0.040103f
C1884 VP.n22 VSUBS 0.043043f
C1885 VP.n23 VSUBS 0.059985f
C1886 VP.n24 VSUBS 0.024579f
C1887 VP.n25 VSUBS 0.03042f
C1888 VP.n26 VSUBS 0.03042f
C1889 VP.n27 VSUBS 0.03042f
C1890 VP.n28 VSUBS 0.042486f
C1891 VP.n29 VSUBS 1.24699f
C1892 VP.n30 VSUBS 0.042486f
C1893 VP.n31 VSUBS 0.060286f
C1894 VP.n32 VSUBS 0.03042f
C1895 VP.n33 VSUBS 0.03042f
C1896 VP.n34 VSUBS 0.03042f
C1897 VP.n35 VSUBS 0.059985f
C1898 VP.n36 VSUBS 0.043043f
C1899 VP.n37 VSUBS 1.33544f
C1900 VP.n38 VSUBS 0.043699f
.ends

