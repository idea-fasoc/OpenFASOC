* NGSPICE file created from diff_pair_sample_1647.ext - technology: sky130A

.subckt diff_pair_sample_1647 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X1 VTAIL.t1 VP.t0 VDD1.t9 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X2 B.t11 B.t9 B.t10 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0 ps=0 w=5.4 l=1.34
X3 VTAIL.t3 VP.t1 VDD1.t8 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X4 VDD1.t7 VP.t2 VTAIL.t4 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=2.106 ps=11.58 w=5.4 l=1.34
X5 VDD2.t0 VN.t1 VTAIL.t18 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X6 VDD1.t6 VP.t3 VTAIL.t5 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=2.106 ps=11.58 w=5.4 l=1.34
X7 VDD1.t5 VP.t4 VTAIL.t2 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0.891 ps=5.73 w=5.4 l=1.34
X8 VTAIL.t17 VN.t2 VDD2.t6 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X9 VDD2.t1 VN.t3 VTAIL.t16 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=2.106 ps=11.58 w=5.4 l=1.34
X10 VTAIL.t15 VN.t4 VDD2.t2 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X11 B.t8 B.t6 B.t7 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0 ps=0 w=5.4 l=1.34
X12 B.t5 B.t3 B.t4 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0 ps=0 w=5.4 l=1.34
X13 B.t2 B.t0 B.t1 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0 ps=0 w=5.4 l=1.34
X14 VTAIL.t9 VP.t5 VDD1.t4 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X15 VDD2.t8 VN.t5 VTAIL.t14 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X16 VDD2.t7 VN.t6 VTAIL.t13 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0.891 ps=5.73 w=5.4 l=1.34
X17 VDD1.t3 VP.t6 VTAIL.t0 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X18 VDD2.t9 VN.t7 VTAIL.t12 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=2.106 ps=11.58 w=5.4 l=1.34
X19 VTAIL.t8 VP.t7 VDD1.t2 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X20 VDD1.t1 VP.t8 VTAIL.t7 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0.891 ps=5.73 w=5.4 l=1.34
X21 VTAIL.t11 VN.t8 VDD2.t4 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
X22 VDD2.t5 VN.t9 VTAIL.t10 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=2.106 pd=11.58 as=0.891 ps=5.73 w=5.4 l=1.34
X23 VDD1.t0 VP.t9 VTAIL.t6 w_n2974_n2048# sky130_fd_pr__pfet_01v8 ad=0.891 pd=5.73 as=0.891 ps=5.73 w=5.4 l=1.34
R0 VN.n24 VN.n23 169.169
R1 VN.n49 VN.n48 169.169
R2 VN.n47 VN.n25 161.3
R3 VN.n46 VN.n45 161.3
R4 VN.n44 VN.n26 161.3
R5 VN.n43 VN.n42 161.3
R6 VN.n41 VN.n27 161.3
R7 VN.n40 VN.n39 161.3
R8 VN.n38 VN.n29 161.3
R9 VN.n37 VN.n36 161.3
R10 VN.n35 VN.n30 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n22 VN.n0 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n19 VN.n1 161.3
R15 VN.n18 VN.n17 161.3
R16 VN.n15 VN.n2 161.3
R17 VN.n14 VN.n13 161.3
R18 VN.n12 VN.n3 161.3
R19 VN.n11 VN.n10 161.3
R20 VN.n9 VN.n4 161.3
R21 VN.n8 VN.n7 161.3
R22 VN.n6 VN.t6 129.502
R23 VN.n32 VN.t3 129.502
R24 VN.n3 VN.t1 97.1199
R25 VN.n5 VN.t2 97.1199
R26 VN.n16 VN.t0 97.1199
R27 VN.n23 VN.t7 97.1199
R28 VN.n29 VN.t5 97.1199
R29 VN.n31 VN.t4 97.1199
R30 VN.n28 VN.t8 97.1199
R31 VN.n48 VN.t9 97.1199
R32 VN.n10 VN.n9 56.5617
R33 VN.n15 VN.n14 56.5617
R34 VN.n36 VN.n35 56.5617
R35 VN.n41 VN.n40 56.5617
R36 VN.n6 VN.n5 56.0469
R37 VN.n32 VN.n31 56.0469
R38 VN VN.n49 41.635
R39 VN.n22 VN.n21 41.0614
R40 VN.n47 VN.n46 41.0614
R41 VN.n21 VN.n1 40.0926
R42 VN.n46 VN.n26 40.0926
R43 VN.n33 VN.n32 26.3169
R44 VN.n7 VN.n6 26.3169
R45 VN.n9 VN.n8 24.5923
R46 VN.n10 VN.n3 24.5923
R47 VN.n14 VN.n3 24.5923
R48 VN.n17 VN.n15 24.5923
R49 VN.n35 VN.n34 24.5923
R50 VN.n40 VN.n29 24.5923
R51 VN.n36 VN.n29 24.5923
R52 VN.n42 VN.n41 24.5923
R53 VN.n23 VN.n22 16.7229
R54 VN.n48 VN.n47 16.7229
R55 VN.n16 VN.n1 16.2311
R56 VN.n28 VN.n26 16.2311
R57 VN.n8 VN.n5 8.36172
R58 VN.n17 VN.n16 8.36172
R59 VN.n34 VN.n31 8.36172
R60 VN.n42 VN.n28 8.36172
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n30 0.189894
R70 VN.n33 VN.n30 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n11 VN.n4 0.189894
R73 VN.n12 VN.n11 0.189894
R74 VN.n13 VN.n12 0.189894
R75 VN.n13 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VDD2.n53 VDD2.n31 756.745
R83 VDD2.n22 VDD2.n0 756.745
R84 VDD2.n54 VDD2.n53 585
R85 VDD2.n52 VDD2.n51 585
R86 VDD2.n35 VDD2.n34 585
R87 VDD2.n46 VDD2.n45 585
R88 VDD2.n44 VDD2.n43 585
R89 VDD2.n39 VDD2.n38 585
R90 VDD2.n8 VDD2.n7 585
R91 VDD2.n13 VDD2.n12 585
R92 VDD2.n15 VDD2.n14 585
R93 VDD2.n4 VDD2.n3 585
R94 VDD2.n21 VDD2.n20 585
R95 VDD2.n23 VDD2.n22 585
R96 VDD2.n40 VDD2.t5 327.856
R97 VDD2.n9 VDD2.t7 327.856
R98 VDD2.n53 VDD2.n52 171.744
R99 VDD2.n52 VDD2.n34 171.744
R100 VDD2.n45 VDD2.n34 171.744
R101 VDD2.n45 VDD2.n44 171.744
R102 VDD2.n44 VDD2.n38 171.744
R103 VDD2.n13 VDD2.n7 171.744
R104 VDD2.n14 VDD2.n13 171.744
R105 VDD2.n14 VDD2.n3 171.744
R106 VDD2.n21 VDD2.n3 171.744
R107 VDD2.n22 VDD2.n21 171.744
R108 VDD2.n30 VDD2.n29 100.683
R109 VDD2 VDD2.n61 100.68
R110 VDD2.n60 VDD2.n59 99.6582
R111 VDD2.n28 VDD2.n27 99.658
R112 VDD2.t5 VDD2.n38 85.8723
R113 VDD2.t7 VDD2.n7 85.8723
R114 VDD2.n28 VDD2.n26 52.6311
R115 VDD2.n58 VDD2.n57 51.1914
R116 VDD2.n58 VDD2.n30 35.2088
R117 VDD2.n40 VDD2.n39 16.381
R118 VDD2.n9 VDD2.n8 16.381
R119 VDD2.n43 VDD2.n42 12.8005
R120 VDD2.n12 VDD2.n11 12.8005
R121 VDD2.n46 VDD2.n37 12.0247
R122 VDD2.n15 VDD2.n6 12.0247
R123 VDD2.n47 VDD2.n35 11.249
R124 VDD2.n16 VDD2.n4 11.249
R125 VDD2.n51 VDD2.n50 10.4732
R126 VDD2.n20 VDD2.n19 10.4732
R127 VDD2.n54 VDD2.n33 9.69747
R128 VDD2.n23 VDD2.n2 9.69747
R129 VDD2.n57 VDD2.n56 9.45567
R130 VDD2.n26 VDD2.n25 9.45567
R131 VDD2.n56 VDD2.n55 9.3005
R132 VDD2.n33 VDD2.n32 9.3005
R133 VDD2.n50 VDD2.n49 9.3005
R134 VDD2.n48 VDD2.n47 9.3005
R135 VDD2.n37 VDD2.n36 9.3005
R136 VDD2.n42 VDD2.n41 9.3005
R137 VDD2.n25 VDD2.n24 9.3005
R138 VDD2.n2 VDD2.n1 9.3005
R139 VDD2.n19 VDD2.n18 9.3005
R140 VDD2.n17 VDD2.n16 9.3005
R141 VDD2.n6 VDD2.n5 9.3005
R142 VDD2.n11 VDD2.n10 9.3005
R143 VDD2.n55 VDD2.n31 8.92171
R144 VDD2.n24 VDD2.n0 8.92171
R145 VDD2.n61 VDD2.t2 6.01994
R146 VDD2.n61 VDD2.t1 6.01994
R147 VDD2.n59 VDD2.t4 6.01994
R148 VDD2.n59 VDD2.t8 6.01994
R149 VDD2.n29 VDD2.t3 6.01994
R150 VDD2.n29 VDD2.t9 6.01994
R151 VDD2.n27 VDD2.t6 6.01994
R152 VDD2.n27 VDD2.t0 6.01994
R153 VDD2.n57 VDD2.n31 5.04292
R154 VDD2.n26 VDD2.n0 5.04292
R155 VDD2.n55 VDD2.n54 4.26717
R156 VDD2.n24 VDD2.n23 4.26717
R157 VDD2.n41 VDD2.n40 3.71853
R158 VDD2.n10 VDD2.n9 3.71853
R159 VDD2.n51 VDD2.n33 3.49141
R160 VDD2.n20 VDD2.n2 3.49141
R161 VDD2.n50 VDD2.n35 2.71565
R162 VDD2.n19 VDD2.n4 2.71565
R163 VDD2.n47 VDD2.n46 1.93989
R164 VDD2.n16 VDD2.n15 1.93989
R165 VDD2.n60 VDD2.n58 1.44016
R166 VDD2.n43 VDD2.n37 1.16414
R167 VDD2.n12 VDD2.n6 1.16414
R168 VDD2 VDD2.n60 0.418603
R169 VDD2.n42 VDD2.n39 0.388379
R170 VDD2.n11 VDD2.n8 0.388379
R171 VDD2.n30 VDD2.n28 0.305068
R172 VDD2.n56 VDD2.n32 0.155672
R173 VDD2.n49 VDD2.n32 0.155672
R174 VDD2.n49 VDD2.n48 0.155672
R175 VDD2.n48 VDD2.n36 0.155672
R176 VDD2.n41 VDD2.n36 0.155672
R177 VDD2.n10 VDD2.n5 0.155672
R178 VDD2.n17 VDD2.n5 0.155672
R179 VDD2.n18 VDD2.n17 0.155672
R180 VDD2.n18 VDD2.n1 0.155672
R181 VDD2.n25 VDD2.n1 0.155672
R182 VTAIL.n120 VTAIL.n98 756.745
R183 VTAIL.n24 VTAIL.n2 756.745
R184 VTAIL.n92 VTAIL.n70 756.745
R185 VTAIL.n60 VTAIL.n38 756.745
R186 VTAIL.n106 VTAIL.n105 585
R187 VTAIL.n111 VTAIL.n110 585
R188 VTAIL.n113 VTAIL.n112 585
R189 VTAIL.n102 VTAIL.n101 585
R190 VTAIL.n119 VTAIL.n118 585
R191 VTAIL.n121 VTAIL.n120 585
R192 VTAIL.n10 VTAIL.n9 585
R193 VTAIL.n15 VTAIL.n14 585
R194 VTAIL.n17 VTAIL.n16 585
R195 VTAIL.n6 VTAIL.n5 585
R196 VTAIL.n23 VTAIL.n22 585
R197 VTAIL.n25 VTAIL.n24 585
R198 VTAIL.n93 VTAIL.n92 585
R199 VTAIL.n91 VTAIL.n90 585
R200 VTAIL.n74 VTAIL.n73 585
R201 VTAIL.n85 VTAIL.n84 585
R202 VTAIL.n83 VTAIL.n82 585
R203 VTAIL.n78 VTAIL.n77 585
R204 VTAIL.n61 VTAIL.n60 585
R205 VTAIL.n59 VTAIL.n58 585
R206 VTAIL.n42 VTAIL.n41 585
R207 VTAIL.n53 VTAIL.n52 585
R208 VTAIL.n51 VTAIL.n50 585
R209 VTAIL.n46 VTAIL.n45 585
R210 VTAIL.n107 VTAIL.t12 327.856
R211 VTAIL.n11 VTAIL.t5 327.856
R212 VTAIL.n79 VTAIL.t4 327.856
R213 VTAIL.n47 VTAIL.t16 327.856
R214 VTAIL.n111 VTAIL.n105 171.744
R215 VTAIL.n112 VTAIL.n111 171.744
R216 VTAIL.n112 VTAIL.n101 171.744
R217 VTAIL.n119 VTAIL.n101 171.744
R218 VTAIL.n120 VTAIL.n119 171.744
R219 VTAIL.n15 VTAIL.n9 171.744
R220 VTAIL.n16 VTAIL.n15 171.744
R221 VTAIL.n16 VTAIL.n5 171.744
R222 VTAIL.n23 VTAIL.n5 171.744
R223 VTAIL.n24 VTAIL.n23 171.744
R224 VTAIL.n92 VTAIL.n91 171.744
R225 VTAIL.n91 VTAIL.n73 171.744
R226 VTAIL.n84 VTAIL.n73 171.744
R227 VTAIL.n84 VTAIL.n83 171.744
R228 VTAIL.n83 VTAIL.n77 171.744
R229 VTAIL.n60 VTAIL.n59 171.744
R230 VTAIL.n59 VTAIL.n41 171.744
R231 VTAIL.n52 VTAIL.n41 171.744
R232 VTAIL.n52 VTAIL.n51 171.744
R233 VTAIL.n51 VTAIL.n45 171.744
R234 VTAIL.t12 VTAIL.n105 85.8723
R235 VTAIL.t5 VTAIL.n9 85.8723
R236 VTAIL.t4 VTAIL.n77 85.8723
R237 VTAIL.t16 VTAIL.n45 85.8723
R238 VTAIL.n69 VTAIL.n68 82.9794
R239 VTAIL.n67 VTAIL.n66 82.9794
R240 VTAIL.n37 VTAIL.n36 82.9794
R241 VTAIL.n35 VTAIL.n34 82.9794
R242 VTAIL.n127 VTAIL.n126 82.9793
R243 VTAIL.n1 VTAIL.n0 82.9793
R244 VTAIL.n31 VTAIL.n30 82.9793
R245 VTAIL.n33 VTAIL.n32 82.9793
R246 VTAIL.n125 VTAIL.n124 34.5126
R247 VTAIL.n29 VTAIL.n28 34.5126
R248 VTAIL.n97 VTAIL.n96 34.5126
R249 VTAIL.n65 VTAIL.n64 34.5126
R250 VTAIL.n35 VTAIL.n33 19.9014
R251 VTAIL.n125 VTAIL.n97 18.4617
R252 VTAIL.n107 VTAIL.n106 16.381
R253 VTAIL.n11 VTAIL.n10 16.381
R254 VTAIL.n79 VTAIL.n78 16.381
R255 VTAIL.n47 VTAIL.n46 16.381
R256 VTAIL.n110 VTAIL.n109 12.8005
R257 VTAIL.n14 VTAIL.n13 12.8005
R258 VTAIL.n82 VTAIL.n81 12.8005
R259 VTAIL.n50 VTAIL.n49 12.8005
R260 VTAIL.n113 VTAIL.n104 12.0247
R261 VTAIL.n17 VTAIL.n8 12.0247
R262 VTAIL.n85 VTAIL.n76 12.0247
R263 VTAIL.n53 VTAIL.n44 12.0247
R264 VTAIL.n114 VTAIL.n102 11.249
R265 VTAIL.n18 VTAIL.n6 11.249
R266 VTAIL.n86 VTAIL.n74 11.249
R267 VTAIL.n54 VTAIL.n42 11.249
R268 VTAIL.n118 VTAIL.n117 10.4732
R269 VTAIL.n22 VTAIL.n21 10.4732
R270 VTAIL.n90 VTAIL.n89 10.4732
R271 VTAIL.n58 VTAIL.n57 10.4732
R272 VTAIL.n121 VTAIL.n100 9.69747
R273 VTAIL.n25 VTAIL.n4 9.69747
R274 VTAIL.n93 VTAIL.n72 9.69747
R275 VTAIL.n61 VTAIL.n40 9.69747
R276 VTAIL.n124 VTAIL.n123 9.45567
R277 VTAIL.n28 VTAIL.n27 9.45567
R278 VTAIL.n96 VTAIL.n95 9.45567
R279 VTAIL.n64 VTAIL.n63 9.45567
R280 VTAIL.n123 VTAIL.n122 9.3005
R281 VTAIL.n100 VTAIL.n99 9.3005
R282 VTAIL.n117 VTAIL.n116 9.3005
R283 VTAIL.n115 VTAIL.n114 9.3005
R284 VTAIL.n104 VTAIL.n103 9.3005
R285 VTAIL.n109 VTAIL.n108 9.3005
R286 VTAIL.n27 VTAIL.n26 9.3005
R287 VTAIL.n4 VTAIL.n3 9.3005
R288 VTAIL.n21 VTAIL.n20 9.3005
R289 VTAIL.n19 VTAIL.n18 9.3005
R290 VTAIL.n8 VTAIL.n7 9.3005
R291 VTAIL.n13 VTAIL.n12 9.3005
R292 VTAIL.n95 VTAIL.n94 9.3005
R293 VTAIL.n72 VTAIL.n71 9.3005
R294 VTAIL.n89 VTAIL.n88 9.3005
R295 VTAIL.n87 VTAIL.n86 9.3005
R296 VTAIL.n76 VTAIL.n75 9.3005
R297 VTAIL.n81 VTAIL.n80 9.3005
R298 VTAIL.n63 VTAIL.n62 9.3005
R299 VTAIL.n40 VTAIL.n39 9.3005
R300 VTAIL.n57 VTAIL.n56 9.3005
R301 VTAIL.n55 VTAIL.n54 9.3005
R302 VTAIL.n44 VTAIL.n43 9.3005
R303 VTAIL.n49 VTAIL.n48 9.3005
R304 VTAIL.n122 VTAIL.n98 8.92171
R305 VTAIL.n26 VTAIL.n2 8.92171
R306 VTAIL.n94 VTAIL.n70 8.92171
R307 VTAIL.n62 VTAIL.n38 8.92171
R308 VTAIL.n126 VTAIL.t18 6.01994
R309 VTAIL.n126 VTAIL.t19 6.01994
R310 VTAIL.n0 VTAIL.t13 6.01994
R311 VTAIL.n0 VTAIL.t17 6.01994
R312 VTAIL.n30 VTAIL.t6 6.01994
R313 VTAIL.n30 VTAIL.t1 6.01994
R314 VTAIL.n32 VTAIL.t2 6.01994
R315 VTAIL.n32 VTAIL.t9 6.01994
R316 VTAIL.n68 VTAIL.t0 6.01994
R317 VTAIL.n68 VTAIL.t3 6.01994
R318 VTAIL.n66 VTAIL.t7 6.01994
R319 VTAIL.n66 VTAIL.t8 6.01994
R320 VTAIL.n36 VTAIL.t14 6.01994
R321 VTAIL.n36 VTAIL.t15 6.01994
R322 VTAIL.n34 VTAIL.t10 6.01994
R323 VTAIL.n34 VTAIL.t11 6.01994
R324 VTAIL.n124 VTAIL.n98 5.04292
R325 VTAIL.n28 VTAIL.n2 5.04292
R326 VTAIL.n96 VTAIL.n70 5.04292
R327 VTAIL.n64 VTAIL.n38 5.04292
R328 VTAIL.n122 VTAIL.n121 4.26717
R329 VTAIL.n26 VTAIL.n25 4.26717
R330 VTAIL.n94 VTAIL.n93 4.26717
R331 VTAIL.n62 VTAIL.n61 4.26717
R332 VTAIL.n80 VTAIL.n79 3.71853
R333 VTAIL.n48 VTAIL.n47 3.71853
R334 VTAIL.n108 VTAIL.n107 3.71853
R335 VTAIL.n12 VTAIL.n11 3.71853
R336 VTAIL.n118 VTAIL.n100 3.49141
R337 VTAIL.n22 VTAIL.n4 3.49141
R338 VTAIL.n90 VTAIL.n72 3.49141
R339 VTAIL.n58 VTAIL.n40 3.49141
R340 VTAIL.n117 VTAIL.n102 2.71565
R341 VTAIL.n21 VTAIL.n6 2.71565
R342 VTAIL.n89 VTAIL.n74 2.71565
R343 VTAIL.n57 VTAIL.n42 2.71565
R344 VTAIL.n114 VTAIL.n113 1.93989
R345 VTAIL.n18 VTAIL.n17 1.93989
R346 VTAIL.n86 VTAIL.n85 1.93989
R347 VTAIL.n54 VTAIL.n53 1.93989
R348 VTAIL.n37 VTAIL.n35 1.44016
R349 VTAIL.n65 VTAIL.n37 1.44016
R350 VTAIL.n69 VTAIL.n67 1.44016
R351 VTAIL.n97 VTAIL.n69 1.44016
R352 VTAIL.n33 VTAIL.n31 1.44016
R353 VTAIL.n31 VTAIL.n29 1.44016
R354 VTAIL.n127 VTAIL.n125 1.44016
R355 VTAIL.n67 VTAIL.n65 1.19016
R356 VTAIL.n29 VTAIL.n1 1.19016
R357 VTAIL.n110 VTAIL.n104 1.16414
R358 VTAIL.n14 VTAIL.n8 1.16414
R359 VTAIL.n82 VTAIL.n76 1.16414
R360 VTAIL.n50 VTAIL.n44 1.16414
R361 VTAIL VTAIL.n1 1.13843
R362 VTAIL.n109 VTAIL.n106 0.388379
R363 VTAIL.n13 VTAIL.n10 0.388379
R364 VTAIL.n81 VTAIL.n78 0.388379
R365 VTAIL.n49 VTAIL.n46 0.388379
R366 VTAIL VTAIL.n127 0.302224
R367 VTAIL.n108 VTAIL.n103 0.155672
R368 VTAIL.n115 VTAIL.n103 0.155672
R369 VTAIL.n116 VTAIL.n115 0.155672
R370 VTAIL.n116 VTAIL.n99 0.155672
R371 VTAIL.n123 VTAIL.n99 0.155672
R372 VTAIL.n12 VTAIL.n7 0.155672
R373 VTAIL.n19 VTAIL.n7 0.155672
R374 VTAIL.n20 VTAIL.n19 0.155672
R375 VTAIL.n20 VTAIL.n3 0.155672
R376 VTAIL.n27 VTAIL.n3 0.155672
R377 VTAIL.n95 VTAIL.n71 0.155672
R378 VTAIL.n88 VTAIL.n71 0.155672
R379 VTAIL.n88 VTAIL.n87 0.155672
R380 VTAIL.n87 VTAIL.n75 0.155672
R381 VTAIL.n80 VTAIL.n75 0.155672
R382 VTAIL.n63 VTAIL.n39 0.155672
R383 VTAIL.n56 VTAIL.n39 0.155672
R384 VTAIL.n56 VTAIL.n55 0.155672
R385 VTAIL.n55 VTAIL.n43 0.155672
R386 VTAIL.n48 VTAIL.n43 0.155672
R387 VP.n33 VP.n7 169.169
R388 VP.n56 VP.n55 169.169
R389 VP.n32 VP.n31 169.169
R390 VP.n16 VP.n15 161.3
R391 VP.n17 VP.n12 161.3
R392 VP.n19 VP.n18 161.3
R393 VP.n20 VP.n11 161.3
R394 VP.n22 VP.n21 161.3
R395 VP.n23 VP.n10 161.3
R396 VP.n26 VP.n25 161.3
R397 VP.n27 VP.n9 161.3
R398 VP.n29 VP.n28 161.3
R399 VP.n30 VP.n8 161.3
R400 VP.n54 VP.n0 161.3
R401 VP.n53 VP.n52 161.3
R402 VP.n51 VP.n1 161.3
R403 VP.n50 VP.n49 161.3
R404 VP.n47 VP.n2 161.3
R405 VP.n46 VP.n45 161.3
R406 VP.n44 VP.n3 161.3
R407 VP.n43 VP.n42 161.3
R408 VP.n41 VP.n4 161.3
R409 VP.n40 VP.n39 161.3
R410 VP.n38 VP.n37 161.3
R411 VP.n36 VP.n6 161.3
R412 VP.n35 VP.n34 161.3
R413 VP.n14 VP.t8 129.502
R414 VP.n3 VP.t9 97.1199
R415 VP.n7 VP.t4 97.1199
R416 VP.n5 VP.t5 97.1199
R417 VP.n48 VP.t0 97.1199
R418 VP.n55 VP.t3 97.1199
R419 VP.n11 VP.t6 97.1199
R420 VP.n31 VP.t2 97.1199
R421 VP.n24 VP.t1 97.1199
R422 VP.n13 VP.t7 97.1199
R423 VP.n42 VP.n41 56.5617
R424 VP.n47 VP.n46 56.5617
R425 VP.n23 VP.n22 56.5617
R426 VP.n18 VP.n17 56.5617
R427 VP.n14 VP.n13 56.047
R428 VP.n33 VP.n32 41.2543
R429 VP.n36 VP.n35 41.0614
R430 VP.n54 VP.n53 41.0614
R431 VP.n30 VP.n29 41.0614
R432 VP.n37 VP.n36 40.0926
R433 VP.n53 VP.n1 40.0926
R434 VP.n29 VP.n9 40.0926
R435 VP.n15 VP.n14 26.3169
R436 VP.n41 VP.n40 24.5923
R437 VP.n42 VP.n3 24.5923
R438 VP.n46 VP.n3 24.5923
R439 VP.n49 VP.n47 24.5923
R440 VP.n25 VP.n23 24.5923
R441 VP.n18 VP.n11 24.5923
R442 VP.n22 VP.n11 24.5923
R443 VP.n17 VP.n16 24.5923
R444 VP.n35 VP.n7 16.7229
R445 VP.n55 VP.n54 16.7229
R446 VP.n31 VP.n30 16.7229
R447 VP.n37 VP.n5 16.2311
R448 VP.n48 VP.n1 16.2311
R449 VP.n24 VP.n9 16.2311
R450 VP.n40 VP.n5 8.36172
R451 VP.n49 VP.n48 8.36172
R452 VP.n25 VP.n24 8.36172
R453 VP.n16 VP.n13 8.36172
R454 VP.n15 VP.n12 0.189894
R455 VP.n19 VP.n12 0.189894
R456 VP.n20 VP.n19 0.189894
R457 VP.n21 VP.n20 0.189894
R458 VP.n21 VP.n10 0.189894
R459 VP.n26 VP.n10 0.189894
R460 VP.n27 VP.n26 0.189894
R461 VP.n28 VP.n27 0.189894
R462 VP.n28 VP.n8 0.189894
R463 VP.n32 VP.n8 0.189894
R464 VP.n34 VP.n33 0.189894
R465 VP.n34 VP.n6 0.189894
R466 VP.n38 VP.n6 0.189894
R467 VP.n39 VP.n38 0.189894
R468 VP.n39 VP.n4 0.189894
R469 VP.n43 VP.n4 0.189894
R470 VP.n44 VP.n43 0.189894
R471 VP.n45 VP.n44 0.189894
R472 VP.n45 VP.n2 0.189894
R473 VP.n50 VP.n2 0.189894
R474 VP.n51 VP.n50 0.189894
R475 VP.n52 VP.n51 0.189894
R476 VP.n52 VP.n0 0.189894
R477 VP.n56 VP.n0 0.189894
R478 VP VP.n56 0.0516364
R479 VDD1.n22 VDD1.n0 756.745
R480 VDD1.n51 VDD1.n29 756.745
R481 VDD1.n23 VDD1.n22 585
R482 VDD1.n21 VDD1.n20 585
R483 VDD1.n4 VDD1.n3 585
R484 VDD1.n15 VDD1.n14 585
R485 VDD1.n13 VDD1.n12 585
R486 VDD1.n8 VDD1.n7 585
R487 VDD1.n37 VDD1.n36 585
R488 VDD1.n42 VDD1.n41 585
R489 VDD1.n44 VDD1.n43 585
R490 VDD1.n33 VDD1.n32 585
R491 VDD1.n50 VDD1.n49 585
R492 VDD1.n52 VDD1.n51 585
R493 VDD1.n9 VDD1.t1 327.856
R494 VDD1.n38 VDD1.t5 327.856
R495 VDD1.n22 VDD1.n21 171.744
R496 VDD1.n21 VDD1.n3 171.744
R497 VDD1.n14 VDD1.n3 171.744
R498 VDD1.n14 VDD1.n13 171.744
R499 VDD1.n13 VDD1.n7 171.744
R500 VDD1.n42 VDD1.n36 171.744
R501 VDD1.n43 VDD1.n42 171.744
R502 VDD1.n43 VDD1.n32 171.744
R503 VDD1.n50 VDD1.n32 171.744
R504 VDD1.n51 VDD1.n50 171.744
R505 VDD1.n59 VDD1.n58 100.683
R506 VDD1.n28 VDD1.n27 99.6582
R507 VDD1.n57 VDD1.n56 99.658
R508 VDD1.n61 VDD1.n60 99.658
R509 VDD1.t1 VDD1.n7 85.8723
R510 VDD1.t5 VDD1.n36 85.8723
R511 VDD1.n28 VDD1.n26 52.6311
R512 VDD1.n57 VDD1.n55 52.6311
R513 VDD1.n61 VDD1.n59 36.5117
R514 VDD1.n9 VDD1.n8 16.381
R515 VDD1.n38 VDD1.n37 16.381
R516 VDD1.n12 VDD1.n11 12.8005
R517 VDD1.n41 VDD1.n40 12.8005
R518 VDD1.n15 VDD1.n6 12.0247
R519 VDD1.n44 VDD1.n35 12.0247
R520 VDD1.n16 VDD1.n4 11.249
R521 VDD1.n45 VDD1.n33 11.249
R522 VDD1.n20 VDD1.n19 10.4732
R523 VDD1.n49 VDD1.n48 10.4732
R524 VDD1.n23 VDD1.n2 9.69747
R525 VDD1.n52 VDD1.n31 9.69747
R526 VDD1.n26 VDD1.n25 9.45567
R527 VDD1.n55 VDD1.n54 9.45567
R528 VDD1.n25 VDD1.n24 9.3005
R529 VDD1.n2 VDD1.n1 9.3005
R530 VDD1.n19 VDD1.n18 9.3005
R531 VDD1.n17 VDD1.n16 9.3005
R532 VDD1.n6 VDD1.n5 9.3005
R533 VDD1.n11 VDD1.n10 9.3005
R534 VDD1.n54 VDD1.n53 9.3005
R535 VDD1.n31 VDD1.n30 9.3005
R536 VDD1.n48 VDD1.n47 9.3005
R537 VDD1.n46 VDD1.n45 9.3005
R538 VDD1.n35 VDD1.n34 9.3005
R539 VDD1.n40 VDD1.n39 9.3005
R540 VDD1.n24 VDD1.n0 8.92171
R541 VDD1.n53 VDD1.n29 8.92171
R542 VDD1.n60 VDD1.t8 6.01994
R543 VDD1.n60 VDD1.t7 6.01994
R544 VDD1.n27 VDD1.t2 6.01994
R545 VDD1.n27 VDD1.t3 6.01994
R546 VDD1.n58 VDD1.t9 6.01994
R547 VDD1.n58 VDD1.t6 6.01994
R548 VDD1.n56 VDD1.t4 6.01994
R549 VDD1.n56 VDD1.t0 6.01994
R550 VDD1.n26 VDD1.n0 5.04292
R551 VDD1.n55 VDD1.n29 5.04292
R552 VDD1.n24 VDD1.n23 4.26717
R553 VDD1.n53 VDD1.n52 4.26717
R554 VDD1.n10 VDD1.n9 3.71853
R555 VDD1.n39 VDD1.n38 3.71853
R556 VDD1.n20 VDD1.n2 3.49141
R557 VDD1.n49 VDD1.n31 3.49141
R558 VDD1.n19 VDD1.n4 2.71565
R559 VDD1.n48 VDD1.n33 2.71565
R560 VDD1.n16 VDD1.n15 1.93989
R561 VDD1.n45 VDD1.n44 1.93989
R562 VDD1.n12 VDD1.n6 1.16414
R563 VDD1.n41 VDD1.n35 1.16414
R564 VDD1 VDD1.n61 1.02205
R565 VDD1 VDD1.n28 0.418603
R566 VDD1.n11 VDD1.n8 0.388379
R567 VDD1.n40 VDD1.n37 0.388379
R568 VDD1.n59 VDD1.n57 0.305068
R569 VDD1.n25 VDD1.n1 0.155672
R570 VDD1.n18 VDD1.n1 0.155672
R571 VDD1.n18 VDD1.n17 0.155672
R572 VDD1.n17 VDD1.n5 0.155672
R573 VDD1.n10 VDD1.n5 0.155672
R574 VDD1.n39 VDD1.n34 0.155672
R575 VDD1.n46 VDD1.n34 0.155672
R576 VDD1.n47 VDD1.n46 0.155672
R577 VDD1.n47 VDD1.n30 0.155672
R578 VDD1.n54 VDD1.n30 0.155672
R579 B.n276 B.n275 585
R580 B.n274 B.n91 585
R581 B.n273 B.n272 585
R582 B.n271 B.n92 585
R583 B.n270 B.n269 585
R584 B.n268 B.n93 585
R585 B.n267 B.n266 585
R586 B.n265 B.n94 585
R587 B.n264 B.n263 585
R588 B.n262 B.n95 585
R589 B.n261 B.n260 585
R590 B.n259 B.n96 585
R591 B.n258 B.n257 585
R592 B.n256 B.n97 585
R593 B.n255 B.n254 585
R594 B.n253 B.n98 585
R595 B.n252 B.n251 585
R596 B.n250 B.n99 585
R597 B.n249 B.n248 585
R598 B.n247 B.n100 585
R599 B.n246 B.n245 585
R600 B.n244 B.n101 585
R601 B.n243 B.n242 585
R602 B.n238 B.n102 585
R603 B.n237 B.n236 585
R604 B.n235 B.n103 585
R605 B.n234 B.n233 585
R606 B.n232 B.n104 585
R607 B.n231 B.n230 585
R608 B.n229 B.n105 585
R609 B.n228 B.n227 585
R610 B.n226 B.n106 585
R611 B.n224 B.n223 585
R612 B.n222 B.n109 585
R613 B.n221 B.n220 585
R614 B.n219 B.n110 585
R615 B.n218 B.n217 585
R616 B.n216 B.n111 585
R617 B.n215 B.n214 585
R618 B.n213 B.n112 585
R619 B.n212 B.n211 585
R620 B.n210 B.n113 585
R621 B.n209 B.n208 585
R622 B.n207 B.n114 585
R623 B.n206 B.n205 585
R624 B.n204 B.n115 585
R625 B.n203 B.n202 585
R626 B.n201 B.n116 585
R627 B.n200 B.n199 585
R628 B.n198 B.n117 585
R629 B.n197 B.n196 585
R630 B.n195 B.n118 585
R631 B.n194 B.n193 585
R632 B.n192 B.n119 585
R633 B.n277 B.n90 585
R634 B.n279 B.n278 585
R635 B.n280 B.n89 585
R636 B.n282 B.n281 585
R637 B.n283 B.n88 585
R638 B.n285 B.n284 585
R639 B.n286 B.n87 585
R640 B.n288 B.n287 585
R641 B.n289 B.n86 585
R642 B.n291 B.n290 585
R643 B.n292 B.n85 585
R644 B.n294 B.n293 585
R645 B.n295 B.n84 585
R646 B.n297 B.n296 585
R647 B.n298 B.n83 585
R648 B.n300 B.n299 585
R649 B.n301 B.n82 585
R650 B.n303 B.n302 585
R651 B.n304 B.n81 585
R652 B.n306 B.n305 585
R653 B.n307 B.n80 585
R654 B.n309 B.n308 585
R655 B.n310 B.n79 585
R656 B.n312 B.n311 585
R657 B.n313 B.n78 585
R658 B.n315 B.n314 585
R659 B.n316 B.n77 585
R660 B.n318 B.n317 585
R661 B.n319 B.n76 585
R662 B.n321 B.n320 585
R663 B.n322 B.n75 585
R664 B.n324 B.n323 585
R665 B.n325 B.n74 585
R666 B.n327 B.n326 585
R667 B.n328 B.n73 585
R668 B.n330 B.n329 585
R669 B.n331 B.n72 585
R670 B.n333 B.n332 585
R671 B.n334 B.n71 585
R672 B.n336 B.n335 585
R673 B.n337 B.n70 585
R674 B.n339 B.n338 585
R675 B.n340 B.n69 585
R676 B.n342 B.n341 585
R677 B.n343 B.n68 585
R678 B.n345 B.n344 585
R679 B.n346 B.n67 585
R680 B.n348 B.n347 585
R681 B.n349 B.n66 585
R682 B.n351 B.n350 585
R683 B.n352 B.n65 585
R684 B.n354 B.n353 585
R685 B.n355 B.n64 585
R686 B.n357 B.n356 585
R687 B.n358 B.n63 585
R688 B.n360 B.n359 585
R689 B.n361 B.n62 585
R690 B.n363 B.n362 585
R691 B.n364 B.n61 585
R692 B.n366 B.n365 585
R693 B.n367 B.n60 585
R694 B.n369 B.n368 585
R695 B.n370 B.n59 585
R696 B.n372 B.n371 585
R697 B.n373 B.n58 585
R698 B.n375 B.n374 585
R699 B.n376 B.n57 585
R700 B.n378 B.n377 585
R701 B.n379 B.n56 585
R702 B.n381 B.n380 585
R703 B.n382 B.n55 585
R704 B.n384 B.n383 585
R705 B.n385 B.n54 585
R706 B.n387 B.n386 585
R707 B.n388 B.n53 585
R708 B.n390 B.n389 585
R709 B.n472 B.n471 585
R710 B.n470 B.n21 585
R711 B.n469 B.n468 585
R712 B.n467 B.n22 585
R713 B.n466 B.n465 585
R714 B.n464 B.n23 585
R715 B.n463 B.n462 585
R716 B.n461 B.n24 585
R717 B.n460 B.n459 585
R718 B.n458 B.n25 585
R719 B.n457 B.n456 585
R720 B.n455 B.n26 585
R721 B.n454 B.n453 585
R722 B.n452 B.n27 585
R723 B.n451 B.n450 585
R724 B.n449 B.n28 585
R725 B.n448 B.n447 585
R726 B.n446 B.n29 585
R727 B.n445 B.n444 585
R728 B.n443 B.n30 585
R729 B.n442 B.n441 585
R730 B.n440 B.n31 585
R731 B.n438 B.n437 585
R732 B.n436 B.n34 585
R733 B.n435 B.n434 585
R734 B.n433 B.n35 585
R735 B.n432 B.n431 585
R736 B.n430 B.n36 585
R737 B.n429 B.n428 585
R738 B.n427 B.n37 585
R739 B.n426 B.n425 585
R740 B.n424 B.n38 585
R741 B.n423 B.n422 585
R742 B.n421 B.n39 585
R743 B.n420 B.n419 585
R744 B.n418 B.n43 585
R745 B.n417 B.n416 585
R746 B.n415 B.n44 585
R747 B.n414 B.n413 585
R748 B.n412 B.n45 585
R749 B.n411 B.n410 585
R750 B.n409 B.n46 585
R751 B.n408 B.n407 585
R752 B.n406 B.n47 585
R753 B.n405 B.n404 585
R754 B.n403 B.n48 585
R755 B.n402 B.n401 585
R756 B.n400 B.n49 585
R757 B.n399 B.n398 585
R758 B.n397 B.n50 585
R759 B.n396 B.n395 585
R760 B.n394 B.n51 585
R761 B.n393 B.n392 585
R762 B.n391 B.n52 585
R763 B.n473 B.n20 585
R764 B.n475 B.n474 585
R765 B.n476 B.n19 585
R766 B.n478 B.n477 585
R767 B.n479 B.n18 585
R768 B.n481 B.n480 585
R769 B.n482 B.n17 585
R770 B.n484 B.n483 585
R771 B.n485 B.n16 585
R772 B.n487 B.n486 585
R773 B.n488 B.n15 585
R774 B.n490 B.n489 585
R775 B.n491 B.n14 585
R776 B.n493 B.n492 585
R777 B.n494 B.n13 585
R778 B.n496 B.n495 585
R779 B.n497 B.n12 585
R780 B.n499 B.n498 585
R781 B.n500 B.n11 585
R782 B.n502 B.n501 585
R783 B.n503 B.n10 585
R784 B.n505 B.n504 585
R785 B.n506 B.n9 585
R786 B.n508 B.n507 585
R787 B.n509 B.n8 585
R788 B.n511 B.n510 585
R789 B.n512 B.n7 585
R790 B.n514 B.n513 585
R791 B.n515 B.n6 585
R792 B.n517 B.n516 585
R793 B.n518 B.n5 585
R794 B.n520 B.n519 585
R795 B.n521 B.n4 585
R796 B.n523 B.n522 585
R797 B.n524 B.n3 585
R798 B.n526 B.n525 585
R799 B.n527 B.n0 585
R800 B.n2 B.n1 585
R801 B.n138 B.n137 585
R802 B.n140 B.n139 585
R803 B.n141 B.n136 585
R804 B.n143 B.n142 585
R805 B.n144 B.n135 585
R806 B.n146 B.n145 585
R807 B.n147 B.n134 585
R808 B.n149 B.n148 585
R809 B.n150 B.n133 585
R810 B.n152 B.n151 585
R811 B.n153 B.n132 585
R812 B.n155 B.n154 585
R813 B.n156 B.n131 585
R814 B.n158 B.n157 585
R815 B.n159 B.n130 585
R816 B.n161 B.n160 585
R817 B.n162 B.n129 585
R818 B.n164 B.n163 585
R819 B.n165 B.n128 585
R820 B.n167 B.n166 585
R821 B.n168 B.n127 585
R822 B.n170 B.n169 585
R823 B.n171 B.n126 585
R824 B.n173 B.n172 585
R825 B.n174 B.n125 585
R826 B.n176 B.n175 585
R827 B.n177 B.n124 585
R828 B.n179 B.n178 585
R829 B.n180 B.n123 585
R830 B.n182 B.n181 585
R831 B.n183 B.n122 585
R832 B.n185 B.n184 585
R833 B.n186 B.n121 585
R834 B.n188 B.n187 585
R835 B.n189 B.n120 585
R836 B.n191 B.n190 585
R837 B.n192 B.n191 511.721
R838 B.n275 B.n90 511.721
R839 B.n389 B.n52 511.721
R840 B.n473 B.n472 511.721
R841 B.n107 B.t0 301.909
R842 B.n239 B.t3 301.909
R843 B.n40 B.t9 301.909
R844 B.n32 B.t6 301.909
R845 B.n239 B.t4 290.363
R846 B.n40 B.t11 290.363
R847 B.n107 B.t1 290.363
R848 B.n32 B.t8 290.363
R849 B.n240 B.t5 257.976
R850 B.n41 B.t10 257.976
R851 B.n108 B.t2 257.976
R852 B.n33 B.t7 257.976
R853 B.n529 B.n528 256.663
R854 B.n528 B.n527 235.042
R855 B.n528 B.n2 235.042
R856 B.n193 B.n192 163.367
R857 B.n193 B.n118 163.367
R858 B.n197 B.n118 163.367
R859 B.n198 B.n197 163.367
R860 B.n199 B.n198 163.367
R861 B.n199 B.n116 163.367
R862 B.n203 B.n116 163.367
R863 B.n204 B.n203 163.367
R864 B.n205 B.n204 163.367
R865 B.n205 B.n114 163.367
R866 B.n209 B.n114 163.367
R867 B.n210 B.n209 163.367
R868 B.n211 B.n210 163.367
R869 B.n211 B.n112 163.367
R870 B.n215 B.n112 163.367
R871 B.n216 B.n215 163.367
R872 B.n217 B.n216 163.367
R873 B.n217 B.n110 163.367
R874 B.n221 B.n110 163.367
R875 B.n222 B.n221 163.367
R876 B.n223 B.n222 163.367
R877 B.n223 B.n106 163.367
R878 B.n228 B.n106 163.367
R879 B.n229 B.n228 163.367
R880 B.n230 B.n229 163.367
R881 B.n230 B.n104 163.367
R882 B.n234 B.n104 163.367
R883 B.n235 B.n234 163.367
R884 B.n236 B.n235 163.367
R885 B.n236 B.n102 163.367
R886 B.n243 B.n102 163.367
R887 B.n244 B.n243 163.367
R888 B.n245 B.n244 163.367
R889 B.n245 B.n100 163.367
R890 B.n249 B.n100 163.367
R891 B.n250 B.n249 163.367
R892 B.n251 B.n250 163.367
R893 B.n251 B.n98 163.367
R894 B.n255 B.n98 163.367
R895 B.n256 B.n255 163.367
R896 B.n257 B.n256 163.367
R897 B.n257 B.n96 163.367
R898 B.n261 B.n96 163.367
R899 B.n262 B.n261 163.367
R900 B.n263 B.n262 163.367
R901 B.n263 B.n94 163.367
R902 B.n267 B.n94 163.367
R903 B.n268 B.n267 163.367
R904 B.n269 B.n268 163.367
R905 B.n269 B.n92 163.367
R906 B.n273 B.n92 163.367
R907 B.n274 B.n273 163.367
R908 B.n275 B.n274 163.367
R909 B.n389 B.n388 163.367
R910 B.n388 B.n387 163.367
R911 B.n387 B.n54 163.367
R912 B.n383 B.n54 163.367
R913 B.n383 B.n382 163.367
R914 B.n382 B.n381 163.367
R915 B.n381 B.n56 163.367
R916 B.n377 B.n56 163.367
R917 B.n377 B.n376 163.367
R918 B.n376 B.n375 163.367
R919 B.n375 B.n58 163.367
R920 B.n371 B.n58 163.367
R921 B.n371 B.n370 163.367
R922 B.n370 B.n369 163.367
R923 B.n369 B.n60 163.367
R924 B.n365 B.n60 163.367
R925 B.n365 B.n364 163.367
R926 B.n364 B.n363 163.367
R927 B.n363 B.n62 163.367
R928 B.n359 B.n62 163.367
R929 B.n359 B.n358 163.367
R930 B.n358 B.n357 163.367
R931 B.n357 B.n64 163.367
R932 B.n353 B.n64 163.367
R933 B.n353 B.n352 163.367
R934 B.n352 B.n351 163.367
R935 B.n351 B.n66 163.367
R936 B.n347 B.n66 163.367
R937 B.n347 B.n346 163.367
R938 B.n346 B.n345 163.367
R939 B.n345 B.n68 163.367
R940 B.n341 B.n68 163.367
R941 B.n341 B.n340 163.367
R942 B.n340 B.n339 163.367
R943 B.n339 B.n70 163.367
R944 B.n335 B.n70 163.367
R945 B.n335 B.n334 163.367
R946 B.n334 B.n333 163.367
R947 B.n333 B.n72 163.367
R948 B.n329 B.n72 163.367
R949 B.n329 B.n328 163.367
R950 B.n328 B.n327 163.367
R951 B.n327 B.n74 163.367
R952 B.n323 B.n74 163.367
R953 B.n323 B.n322 163.367
R954 B.n322 B.n321 163.367
R955 B.n321 B.n76 163.367
R956 B.n317 B.n76 163.367
R957 B.n317 B.n316 163.367
R958 B.n316 B.n315 163.367
R959 B.n315 B.n78 163.367
R960 B.n311 B.n78 163.367
R961 B.n311 B.n310 163.367
R962 B.n310 B.n309 163.367
R963 B.n309 B.n80 163.367
R964 B.n305 B.n80 163.367
R965 B.n305 B.n304 163.367
R966 B.n304 B.n303 163.367
R967 B.n303 B.n82 163.367
R968 B.n299 B.n82 163.367
R969 B.n299 B.n298 163.367
R970 B.n298 B.n297 163.367
R971 B.n297 B.n84 163.367
R972 B.n293 B.n84 163.367
R973 B.n293 B.n292 163.367
R974 B.n292 B.n291 163.367
R975 B.n291 B.n86 163.367
R976 B.n287 B.n86 163.367
R977 B.n287 B.n286 163.367
R978 B.n286 B.n285 163.367
R979 B.n285 B.n88 163.367
R980 B.n281 B.n88 163.367
R981 B.n281 B.n280 163.367
R982 B.n280 B.n279 163.367
R983 B.n279 B.n90 163.367
R984 B.n472 B.n21 163.367
R985 B.n468 B.n21 163.367
R986 B.n468 B.n467 163.367
R987 B.n467 B.n466 163.367
R988 B.n466 B.n23 163.367
R989 B.n462 B.n23 163.367
R990 B.n462 B.n461 163.367
R991 B.n461 B.n460 163.367
R992 B.n460 B.n25 163.367
R993 B.n456 B.n25 163.367
R994 B.n456 B.n455 163.367
R995 B.n455 B.n454 163.367
R996 B.n454 B.n27 163.367
R997 B.n450 B.n27 163.367
R998 B.n450 B.n449 163.367
R999 B.n449 B.n448 163.367
R1000 B.n448 B.n29 163.367
R1001 B.n444 B.n29 163.367
R1002 B.n444 B.n443 163.367
R1003 B.n443 B.n442 163.367
R1004 B.n442 B.n31 163.367
R1005 B.n437 B.n31 163.367
R1006 B.n437 B.n436 163.367
R1007 B.n436 B.n435 163.367
R1008 B.n435 B.n35 163.367
R1009 B.n431 B.n35 163.367
R1010 B.n431 B.n430 163.367
R1011 B.n430 B.n429 163.367
R1012 B.n429 B.n37 163.367
R1013 B.n425 B.n37 163.367
R1014 B.n425 B.n424 163.367
R1015 B.n424 B.n423 163.367
R1016 B.n423 B.n39 163.367
R1017 B.n419 B.n39 163.367
R1018 B.n419 B.n418 163.367
R1019 B.n418 B.n417 163.367
R1020 B.n417 B.n44 163.367
R1021 B.n413 B.n44 163.367
R1022 B.n413 B.n412 163.367
R1023 B.n412 B.n411 163.367
R1024 B.n411 B.n46 163.367
R1025 B.n407 B.n46 163.367
R1026 B.n407 B.n406 163.367
R1027 B.n406 B.n405 163.367
R1028 B.n405 B.n48 163.367
R1029 B.n401 B.n48 163.367
R1030 B.n401 B.n400 163.367
R1031 B.n400 B.n399 163.367
R1032 B.n399 B.n50 163.367
R1033 B.n395 B.n50 163.367
R1034 B.n395 B.n394 163.367
R1035 B.n394 B.n393 163.367
R1036 B.n393 B.n52 163.367
R1037 B.n474 B.n473 163.367
R1038 B.n474 B.n19 163.367
R1039 B.n478 B.n19 163.367
R1040 B.n479 B.n478 163.367
R1041 B.n480 B.n479 163.367
R1042 B.n480 B.n17 163.367
R1043 B.n484 B.n17 163.367
R1044 B.n485 B.n484 163.367
R1045 B.n486 B.n485 163.367
R1046 B.n486 B.n15 163.367
R1047 B.n490 B.n15 163.367
R1048 B.n491 B.n490 163.367
R1049 B.n492 B.n491 163.367
R1050 B.n492 B.n13 163.367
R1051 B.n496 B.n13 163.367
R1052 B.n497 B.n496 163.367
R1053 B.n498 B.n497 163.367
R1054 B.n498 B.n11 163.367
R1055 B.n502 B.n11 163.367
R1056 B.n503 B.n502 163.367
R1057 B.n504 B.n503 163.367
R1058 B.n504 B.n9 163.367
R1059 B.n508 B.n9 163.367
R1060 B.n509 B.n508 163.367
R1061 B.n510 B.n509 163.367
R1062 B.n510 B.n7 163.367
R1063 B.n514 B.n7 163.367
R1064 B.n515 B.n514 163.367
R1065 B.n516 B.n515 163.367
R1066 B.n516 B.n5 163.367
R1067 B.n520 B.n5 163.367
R1068 B.n521 B.n520 163.367
R1069 B.n522 B.n521 163.367
R1070 B.n522 B.n3 163.367
R1071 B.n526 B.n3 163.367
R1072 B.n527 B.n526 163.367
R1073 B.n138 B.n2 163.367
R1074 B.n139 B.n138 163.367
R1075 B.n139 B.n136 163.367
R1076 B.n143 B.n136 163.367
R1077 B.n144 B.n143 163.367
R1078 B.n145 B.n144 163.367
R1079 B.n145 B.n134 163.367
R1080 B.n149 B.n134 163.367
R1081 B.n150 B.n149 163.367
R1082 B.n151 B.n150 163.367
R1083 B.n151 B.n132 163.367
R1084 B.n155 B.n132 163.367
R1085 B.n156 B.n155 163.367
R1086 B.n157 B.n156 163.367
R1087 B.n157 B.n130 163.367
R1088 B.n161 B.n130 163.367
R1089 B.n162 B.n161 163.367
R1090 B.n163 B.n162 163.367
R1091 B.n163 B.n128 163.367
R1092 B.n167 B.n128 163.367
R1093 B.n168 B.n167 163.367
R1094 B.n169 B.n168 163.367
R1095 B.n169 B.n126 163.367
R1096 B.n173 B.n126 163.367
R1097 B.n174 B.n173 163.367
R1098 B.n175 B.n174 163.367
R1099 B.n175 B.n124 163.367
R1100 B.n179 B.n124 163.367
R1101 B.n180 B.n179 163.367
R1102 B.n181 B.n180 163.367
R1103 B.n181 B.n122 163.367
R1104 B.n185 B.n122 163.367
R1105 B.n186 B.n185 163.367
R1106 B.n187 B.n186 163.367
R1107 B.n187 B.n120 163.367
R1108 B.n191 B.n120 163.367
R1109 B.n225 B.n108 59.5399
R1110 B.n241 B.n240 59.5399
R1111 B.n42 B.n41 59.5399
R1112 B.n439 B.n33 59.5399
R1113 B.n471 B.n20 33.2493
R1114 B.n391 B.n390 33.2493
R1115 B.n277 B.n276 33.2493
R1116 B.n190 B.n119 33.2493
R1117 B.n108 B.n107 32.3884
R1118 B.n240 B.n239 32.3884
R1119 B.n41 B.n40 32.3884
R1120 B.n33 B.n32 32.3884
R1121 B B.n529 18.0485
R1122 B.n475 B.n20 10.6151
R1123 B.n476 B.n475 10.6151
R1124 B.n477 B.n476 10.6151
R1125 B.n477 B.n18 10.6151
R1126 B.n481 B.n18 10.6151
R1127 B.n482 B.n481 10.6151
R1128 B.n483 B.n482 10.6151
R1129 B.n483 B.n16 10.6151
R1130 B.n487 B.n16 10.6151
R1131 B.n488 B.n487 10.6151
R1132 B.n489 B.n488 10.6151
R1133 B.n489 B.n14 10.6151
R1134 B.n493 B.n14 10.6151
R1135 B.n494 B.n493 10.6151
R1136 B.n495 B.n494 10.6151
R1137 B.n495 B.n12 10.6151
R1138 B.n499 B.n12 10.6151
R1139 B.n500 B.n499 10.6151
R1140 B.n501 B.n500 10.6151
R1141 B.n501 B.n10 10.6151
R1142 B.n505 B.n10 10.6151
R1143 B.n506 B.n505 10.6151
R1144 B.n507 B.n506 10.6151
R1145 B.n507 B.n8 10.6151
R1146 B.n511 B.n8 10.6151
R1147 B.n512 B.n511 10.6151
R1148 B.n513 B.n512 10.6151
R1149 B.n513 B.n6 10.6151
R1150 B.n517 B.n6 10.6151
R1151 B.n518 B.n517 10.6151
R1152 B.n519 B.n518 10.6151
R1153 B.n519 B.n4 10.6151
R1154 B.n523 B.n4 10.6151
R1155 B.n524 B.n523 10.6151
R1156 B.n525 B.n524 10.6151
R1157 B.n525 B.n0 10.6151
R1158 B.n471 B.n470 10.6151
R1159 B.n470 B.n469 10.6151
R1160 B.n469 B.n22 10.6151
R1161 B.n465 B.n22 10.6151
R1162 B.n465 B.n464 10.6151
R1163 B.n464 B.n463 10.6151
R1164 B.n463 B.n24 10.6151
R1165 B.n459 B.n24 10.6151
R1166 B.n459 B.n458 10.6151
R1167 B.n458 B.n457 10.6151
R1168 B.n457 B.n26 10.6151
R1169 B.n453 B.n26 10.6151
R1170 B.n453 B.n452 10.6151
R1171 B.n452 B.n451 10.6151
R1172 B.n451 B.n28 10.6151
R1173 B.n447 B.n28 10.6151
R1174 B.n447 B.n446 10.6151
R1175 B.n446 B.n445 10.6151
R1176 B.n445 B.n30 10.6151
R1177 B.n441 B.n30 10.6151
R1178 B.n441 B.n440 10.6151
R1179 B.n438 B.n34 10.6151
R1180 B.n434 B.n34 10.6151
R1181 B.n434 B.n433 10.6151
R1182 B.n433 B.n432 10.6151
R1183 B.n432 B.n36 10.6151
R1184 B.n428 B.n36 10.6151
R1185 B.n428 B.n427 10.6151
R1186 B.n427 B.n426 10.6151
R1187 B.n426 B.n38 10.6151
R1188 B.n422 B.n421 10.6151
R1189 B.n421 B.n420 10.6151
R1190 B.n420 B.n43 10.6151
R1191 B.n416 B.n43 10.6151
R1192 B.n416 B.n415 10.6151
R1193 B.n415 B.n414 10.6151
R1194 B.n414 B.n45 10.6151
R1195 B.n410 B.n45 10.6151
R1196 B.n410 B.n409 10.6151
R1197 B.n409 B.n408 10.6151
R1198 B.n408 B.n47 10.6151
R1199 B.n404 B.n47 10.6151
R1200 B.n404 B.n403 10.6151
R1201 B.n403 B.n402 10.6151
R1202 B.n402 B.n49 10.6151
R1203 B.n398 B.n49 10.6151
R1204 B.n398 B.n397 10.6151
R1205 B.n397 B.n396 10.6151
R1206 B.n396 B.n51 10.6151
R1207 B.n392 B.n51 10.6151
R1208 B.n392 B.n391 10.6151
R1209 B.n390 B.n53 10.6151
R1210 B.n386 B.n53 10.6151
R1211 B.n386 B.n385 10.6151
R1212 B.n385 B.n384 10.6151
R1213 B.n384 B.n55 10.6151
R1214 B.n380 B.n55 10.6151
R1215 B.n380 B.n379 10.6151
R1216 B.n379 B.n378 10.6151
R1217 B.n378 B.n57 10.6151
R1218 B.n374 B.n57 10.6151
R1219 B.n374 B.n373 10.6151
R1220 B.n373 B.n372 10.6151
R1221 B.n372 B.n59 10.6151
R1222 B.n368 B.n59 10.6151
R1223 B.n368 B.n367 10.6151
R1224 B.n367 B.n366 10.6151
R1225 B.n366 B.n61 10.6151
R1226 B.n362 B.n61 10.6151
R1227 B.n362 B.n361 10.6151
R1228 B.n361 B.n360 10.6151
R1229 B.n360 B.n63 10.6151
R1230 B.n356 B.n63 10.6151
R1231 B.n356 B.n355 10.6151
R1232 B.n355 B.n354 10.6151
R1233 B.n354 B.n65 10.6151
R1234 B.n350 B.n65 10.6151
R1235 B.n350 B.n349 10.6151
R1236 B.n349 B.n348 10.6151
R1237 B.n348 B.n67 10.6151
R1238 B.n344 B.n67 10.6151
R1239 B.n344 B.n343 10.6151
R1240 B.n343 B.n342 10.6151
R1241 B.n342 B.n69 10.6151
R1242 B.n338 B.n69 10.6151
R1243 B.n338 B.n337 10.6151
R1244 B.n337 B.n336 10.6151
R1245 B.n336 B.n71 10.6151
R1246 B.n332 B.n71 10.6151
R1247 B.n332 B.n331 10.6151
R1248 B.n331 B.n330 10.6151
R1249 B.n330 B.n73 10.6151
R1250 B.n326 B.n73 10.6151
R1251 B.n326 B.n325 10.6151
R1252 B.n325 B.n324 10.6151
R1253 B.n324 B.n75 10.6151
R1254 B.n320 B.n75 10.6151
R1255 B.n320 B.n319 10.6151
R1256 B.n319 B.n318 10.6151
R1257 B.n318 B.n77 10.6151
R1258 B.n314 B.n77 10.6151
R1259 B.n314 B.n313 10.6151
R1260 B.n313 B.n312 10.6151
R1261 B.n312 B.n79 10.6151
R1262 B.n308 B.n79 10.6151
R1263 B.n308 B.n307 10.6151
R1264 B.n307 B.n306 10.6151
R1265 B.n306 B.n81 10.6151
R1266 B.n302 B.n81 10.6151
R1267 B.n302 B.n301 10.6151
R1268 B.n301 B.n300 10.6151
R1269 B.n300 B.n83 10.6151
R1270 B.n296 B.n83 10.6151
R1271 B.n296 B.n295 10.6151
R1272 B.n295 B.n294 10.6151
R1273 B.n294 B.n85 10.6151
R1274 B.n290 B.n85 10.6151
R1275 B.n290 B.n289 10.6151
R1276 B.n289 B.n288 10.6151
R1277 B.n288 B.n87 10.6151
R1278 B.n284 B.n87 10.6151
R1279 B.n284 B.n283 10.6151
R1280 B.n283 B.n282 10.6151
R1281 B.n282 B.n89 10.6151
R1282 B.n278 B.n89 10.6151
R1283 B.n278 B.n277 10.6151
R1284 B.n137 B.n1 10.6151
R1285 B.n140 B.n137 10.6151
R1286 B.n141 B.n140 10.6151
R1287 B.n142 B.n141 10.6151
R1288 B.n142 B.n135 10.6151
R1289 B.n146 B.n135 10.6151
R1290 B.n147 B.n146 10.6151
R1291 B.n148 B.n147 10.6151
R1292 B.n148 B.n133 10.6151
R1293 B.n152 B.n133 10.6151
R1294 B.n153 B.n152 10.6151
R1295 B.n154 B.n153 10.6151
R1296 B.n154 B.n131 10.6151
R1297 B.n158 B.n131 10.6151
R1298 B.n159 B.n158 10.6151
R1299 B.n160 B.n159 10.6151
R1300 B.n160 B.n129 10.6151
R1301 B.n164 B.n129 10.6151
R1302 B.n165 B.n164 10.6151
R1303 B.n166 B.n165 10.6151
R1304 B.n166 B.n127 10.6151
R1305 B.n170 B.n127 10.6151
R1306 B.n171 B.n170 10.6151
R1307 B.n172 B.n171 10.6151
R1308 B.n172 B.n125 10.6151
R1309 B.n176 B.n125 10.6151
R1310 B.n177 B.n176 10.6151
R1311 B.n178 B.n177 10.6151
R1312 B.n178 B.n123 10.6151
R1313 B.n182 B.n123 10.6151
R1314 B.n183 B.n182 10.6151
R1315 B.n184 B.n183 10.6151
R1316 B.n184 B.n121 10.6151
R1317 B.n188 B.n121 10.6151
R1318 B.n189 B.n188 10.6151
R1319 B.n190 B.n189 10.6151
R1320 B.n194 B.n119 10.6151
R1321 B.n195 B.n194 10.6151
R1322 B.n196 B.n195 10.6151
R1323 B.n196 B.n117 10.6151
R1324 B.n200 B.n117 10.6151
R1325 B.n201 B.n200 10.6151
R1326 B.n202 B.n201 10.6151
R1327 B.n202 B.n115 10.6151
R1328 B.n206 B.n115 10.6151
R1329 B.n207 B.n206 10.6151
R1330 B.n208 B.n207 10.6151
R1331 B.n208 B.n113 10.6151
R1332 B.n212 B.n113 10.6151
R1333 B.n213 B.n212 10.6151
R1334 B.n214 B.n213 10.6151
R1335 B.n214 B.n111 10.6151
R1336 B.n218 B.n111 10.6151
R1337 B.n219 B.n218 10.6151
R1338 B.n220 B.n219 10.6151
R1339 B.n220 B.n109 10.6151
R1340 B.n224 B.n109 10.6151
R1341 B.n227 B.n226 10.6151
R1342 B.n227 B.n105 10.6151
R1343 B.n231 B.n105 10.6151
R1344 B.n232 B.n231 10.6151
R1345 B.n233 B.n232 10.6151
R1346 B.n233 B.n103 10.6151
R1347 B.n237 B.n103 10.6151
R1348 B.n238 B.n237 10.6151
R1349 B.n242 B.n238 10.6151
R1350 B.n246 B.n101 10.6151
R1351 B.n247 B.n246 10.6151
R1352 B.n248 B.n247 10.6151
R1353 B.n248 B.n99 10.6151
R1354 B.n252 B.n99 10.6151
R1355 B.n253 B.n252 10.6151
R1356 B.n254 B.n253 10.6151
R1357 B.n254 B.n97 10.6151
R1358 B.n258 B.n97 10.6151
R1359 B.n259 B.n258 10.6151
R1360 B.n260 B.n259 10.6151
R1361 B.n260 B.n95 10.6151
R1362 B.n264 B.n95 10.6151
R1363 B.n265 B.n264 10.6151
R1364 B.n266 B.n265 10.6151
R1365 B.n266 B.n93 10.6151
R1366 B.n270 B.n93 10.6151
R1367 B.n271 B.n270 10.6151
R1368 B.n272 B.n271 10.6151
R1369 B.n272 B.n91 10.6151
R1370 B.n276 B.n91 10.6151
R1371 B.n440 B.n439 9.36635
R1372 B.n422 B.n42 9.36635
R1373 B.n225 B.n224 9.36635
R1374 B.n241 B.n101 9.36635
R1375 B.n529 B.n0 8.11757
R1376 B.n529 B.n1 8.11757
R1377 B.n439 B.n438 1.24928
R1378 B.n42 B.n38 1.24928
R1379 B.n226 B.n225 1.24928
R1380 B.n242 B.n241 1.24928
C0 VTAIL VDD1 6.86248f
C1 VTAIL w_n2974_n2048# 2.07239f
C2 VDD2 B 1.54481f
C3 VTAIL VP 4.79147f
C4 VDD1 VN 0.15065f
C5 VN w_n2974_n2048# 5.84776f
C6 VN VP 5.31187f
C7 VDD1 VDD2 1.353f
C8 VDD1 B 1.47582f
C9 VDD2 w_n2974_n2048# 1.90685f
C10 VDD2 VP 0.426286f
C11 B w_n2974_n2048# 6.58347f
C12 B VP 1.52094f
C13 VTAIL VN 4.77721f
C14 VDD1 w_n2974_n2048# 1.82899f
C15 VDD1 VP 4.54353f
C16 w_n2974_n2048# VP 6.23103f
C17 VTAIL VDD2 6.90555f
C18 VTAIL B 1.80888f
C19 VDD2 VN 4.27423f
C20 B VN 0.883333f
C21 VDD2 VSUBS 1.280742f
C22 VDD1 VSUBS 1.218332f
C23 VTAIL VSUBS 0.51152f
C24 VN VSUBS 5.35147f
C25 VP VSUBS 2.247269f
C26 B VSUBS 3.148838f
C27 w_n2974_n2048# VSUBS 76.1939f
C28 B.n0 VSUBS 0.005742f
C29 B.n1 VSUBS 0.005742f
C30 B.n2 VSUBS 0.008492f
C31 B.n3 VSUBS 0.006508f
C32 B.n4 VSUBS 0.006508f
C33 B.n5 VSUBS 0.006508f
C34 B.n6 VSUBS 0.006508f
C35 B.n7 VSUBS 0.006508f
C36 B.n8 VSUBS 0.006508f
C37 B.n9 VSUBS 0.006508f
C38 B.n10 VSUBS 0.006508f
C39 B.n11 VSUBS 0.006508f
C40 B.n12 VSUBS 0.006508f
C41 B.n13 VSUBS 0.006508f
C42 B.n14 VSUBS 0.006508f
C43 B.n15 VSUBS 0.006508f
C44 B.n16 VSUBS 0.006508f
C45 B.n17 VSUBS 0.006508f
C46 B.n18 VSUBS 0.006508f
C47 B.n19 VSUBS 0.006508f
C48 B.n20 VSUBS 0.014993f
C49 B.n21 VSUBS 0.006508f
C50 B.n22 VSUBS 0.006508f
C51 B.n23 VSUBS 0.006508f
C52 B.n24 VSUBS 0.006508f
C53 B.n25 VSUBS 0.006508f
C54 B.n26 VSUBS 0.006508f
C55 B.n27 VSUBS 0.006508f
C56 B.n28 VSUBS 0.006508f
C57 B.n29 VSUBS 0.006508f
C58 B.n30 VSUBS 0.006508f
C59 B.n31 VSUBS 0.006508f
C60 B.t7 VSUBS 0.073916f
C61 B.t8 VSUBS 0.087347f
C62 B.t6 VSUBS 0.308f
C63 B.n32 VSUBS 0.154722f
C64 B.n33 VSUBS 0.129692f
C65 B.n34 VSUBS 0.006508f
C66 B.n35 VSUBS 0.006508f
C67 B.n36 VSUBS 0.006508f
C68 B.n37 VSUBS 0.006508f
C69 B.n38 VSUBS 0.003637f
C70 B.n39 VSUBS 0.006508f
C71 B.t10 VSUBS 0.073917f
C72 B.t11 VSUBS 0.087348f
C73 B.t9 VSUBS 0.308f
C74 B.n40 VSUBS 0.154721f
C75 B.n41 VSUBS 0.129691f
C76 B.n42 VSUBS 0.015077f
C77 B.n43 VSUBS 0.006508f
C78 B.n44 VSUBS 0.006508f
C79 B.n45 VSUBS 0.006508f
C80 B.n46 VSUBS 0.006508f
C81 B.n47 VSUBS 0.006508f
C82 B.n48 VSUBS 0.006508f
C83 B.n49 VSUBS 0.006508f
C84 B.n50 VSUBS 0.006508f
C85 B.n51 VSUBS 0.006508f
C86 B.n52 VSUBS 0.015822f
C87 B.n53 VSUBS 0.006508f
C88 B.n54 VSUBS 0.006508f
C89 B.n55 VSUBS 0.006508f
C90 B.n56 VSUBS 0.006508f
C91 B.n57 VSUBS 0.006508f
C92 B.n58 VSUBS 0.006508f
C93 B.n59 VSUBS 0.006508f
C94 B.n60 VSUBS 0.006508f
C95 B.n61 VSUBS 0.006508f
C96 B.n62 VSUBS 0.006508f
C97 B.n63 VSUBS 0.006508f
C98 B.n64 VSUBS 0.006508f
C99 B.n65 VSUBS 0.006508f
C100 B.n66 VSUBS 0.006508f
C101 B.n67 VSUBS 0.006508f
C102 B.n68 VSUBS 0.006508f
C103 B.n69 VSUBS 0.006508f
C104 B.n70 VSUBS 0.006508f
C105 B.n71 VSUBS 0.006508f
C106 B.n72 VSUBS 0.006508f
C107 B.n73 VSUBS 0.006508f
C108 B.n74 VSUBS 0.006508f
C109 B.n75 VSUBS 0.006508f
C110 B.n76 VSUBS 0.006508f
C111 B.n77 VSUBS 0.006508f
C112 B.n78 VSUBS 0.006508f
C113 B.n79 VSUBS 0.006508f
C114 B.n80 VSUBS 0.006508f
C115 B.n81 VSUBS 0.006508f
C116 B.n82 VSUBS 0.006508f
C117 B.n83 VSUBS 0.006508f
C118 B.n84 VSUBS 0.006508f
C119 B.n85 VSUBS 0.006508f
C120 B.n86 VSUBS 0.006508f
C121 B.n87 VSUBS 0.006508f
C122 B.n88 VSUBS 0.006508f
C123 B.n89 VSUBS 0.006508f
C124 B.n90 VSUBS 0.014993f
C125 B.n91 VSUBS 0.006508f
C126 B.n92 VSUBS 0.006508f
C127 B.n93 VSUBS 0.006508f
C128 B.n94 VSUBS 0.006508f
C129 B.n95 VSUBS 0.006508f
C130 B.n96 VSUBS 0.006508f
C131 B.n97 VSUBS 0.006508f
C132 B.n98 VSUBS 0.006508f
C133 B.n99 VSUBS 0.006508f
C134 B.n100 VSUBS 0.006508f
C135 B.n101 VSUBS 0.006125f
C136 B.n102 VSUBS 0.006508f
C137 B.n103 VSUBS 0.006508f
C138 B.n104 VSUBS 0.006508f
C139 B.n105 VSUBS 0.006508f
C140 B.n106 VSUBS 0.006508f
C141 B.t2 VSUBS 0.073916f
C142 B.t1 VSUBS 0.087347f
C143 B.t0 VSUBS 0.308f
C144 B.n107 VSUBS 0.154722f
C145 B.n108 VSUBS 0.129692f
C146 B.n109 VSUBS 0.006508f
C147 B.n110 VSUBS 0.006508f
C148 B.n111 VSUBS 0.006508f
C149 B.n112 VSUBS 0.006508f
C150 B.n113 VSUBS 0.006508f
C151 B.n114 VSUBS 0.006508f
C152 B.n115 VSUBS 0.006508f
C153 B.n116 VSUBS 0.006508f
C154 B.n117 VSUBS 0.006508f
C155 B.n118 VSUBS 0.006508f
C156 B.n119 VSUBS 0.015822f
C157 B.n120 VSUBS 0.006508f
C158 B.n121 VSUBS 0.006508f
C159 B.n122 VSUBS 0.006508f
C160 B.n123 VSUBS 0.006508f
C161 B.n124 VSUBS 0.006508f
C162 B.n125 VSUBS 0.006508f
C163 B.n126 VSUBS 0.006508f
C164 B.n127 VSUBS 0.006508f
C165 B.n128 VSUBS 0.006508f
C166 B.n129 VSUBS 0.006508f
C167 B.n130 VSUBS 0.006508f
C168 B.n131 VSUBS 0.006508f
C169 B.n132 VSUBS 0.006508f
C170 B.n133 VSUBS 0.006508f
C171 B.n134 VSUBS 0.006508f
C172 B.n135 VSUBS 0.006508f
C173 B.n136 VSUBS 0.006508f
C174 B.n137 VSUBS 0.006508f
C175 B.n138 VSUBS 0.006508f
C176 B.n139 VSUBS 0.006508f
C177 B.n140 VSUBS 0.006508f
C178 B.n141 VSUBS 0.006508f
C179 B.n142 VSUBS 0.006508f
C180 B.n143 VSUBS 0.006508f
C181 B.n144 VSUBS 0.006508f
C182 B.n145 VSUBS 0.006508f
C183 B.n146 VSUBS 0.006508f
C184 B.n147 VSUBS 0.006508f
C185 B.n148 VSUBS 0.006508f
C186 B.n149 VSUBS 0.006508f
C187 B.n150 VSUBS 0.006508f
C188 B.n151 VSUBS 0.006508f
C189 B.n152 VSUBS 0.006508f
C190 B.n153 VSUBS 0.006508f
C191 B.n154 VSUBS 0.006508f
C192 B.n155 VSUBS 0.006508f
C193 B.n156 VSUBS 0.006508f
C194 B.n157 VSUBS 0.006508f
C195 B.n158 VSUBS 0.006508f
C196 B.n159 VSUBS 0.006508f
C197 B.n160 VSUBS 0.006508f
C198 B.n161 VSUBS 0.006508f
C199 B.n162 VSUBS 0.006508f
C200 B.n163 VSUBS 0.006508f
C201 B.n164 VSUBS 0.006508f
C202 B.n165 VSUBS 0.006508f
C203 B.n166 VSUBS 0.006508f
C204 B.n167 VSUBS 0.006508f
C205 B.n168 VSUBS 0.006508f
C206 B.n169 VSUBS 0.006508f
C207 B.n170 VSUBS 0.006508f
C208 B.n171 VSUBS 0.006508f
C209 B.n172 VSUBS 0.006508f
C210 B.n173 VSUBS 0.006508f
C211 B.n174 VSUBS 0.006508f
C212 B.n175 VSUBS 0.006508f
C213 B.n176 VSUBS 0.006508f
C214 B.n177 VSUBS 0.006508f
C215 B.n178 VSUBS 0.006508f
C216 B.n179 VSUBS 0.006508f
C217 B.n180 VSUBS 0.006508f
C218 B.n181 VSUBS 0.006508f
C219 B.n182 VSUBS 0.006508f
C220 B.n183 VSUBS 0.006508f
C221 B.n184 VSUBS 0.006508f
C222 B.n185 VSUBS 0.006508f
C223 B.n186 VSUBS 0.006508f
C224 B.n187 VSUBS 0.006508f
C225 B.n188 VSUBS 0.006508f
C226 B.n189 VSUBS 0.006508f
C227 B.n190 VSUBS 0.014993f
C228 B.n191 VSUBS 0.014993f
C229 B.n192 VSUBS 0.015822f
C230 B.n193 VSUBS 0.006508f
C231 B.n194 VSUBS 0.006508f
C232 B.n195 VSUBS 0.006508f
C233 B.n196 VSUBS 0.006508f
C234 B.n197 VSUBS 0.006508f
C235 B.n198 VSUBS 0.006508f
C236 B.n199 VSUBS 0.006508f
C237 B.n200 VSUBS 0.006508f
C238 B.n201 VSUBS 0.006508f
C239 B.n202 VSUBS 0.006508f
C240 B.n203 VSUBS 0.006508f
C241 B.n204 VSUBS 0.006508f
C242 B.n205 VSUBS 0.006508f
C243 B.n206 VSUBS 0.006508f
C244 B.n207 VSUBS 0.006508f
C245 B.n208 VSUBS 0.006508f
C246 B.n209 VSUBS 0.006508f
C247 B.n210 VSUBS 0.006508f
C248 B.n211 VSUBS 0.006508f
C249 B.n212 VSUBS 0.006508f
C250 B.n213 VSUBS 0.006508f
C251 B.n214 VSUBS 0.006508f
C252 B.n215 VSUBS 0.006508f
C253 B.n216 VSUBS 0.006508f
C254 B.n217 VSUBS 0.006508f
C255 B.n218 VSUBS 0.006508f
C256 B.n219 VSUBS 0.006508f
C257 B.n220 VSUBS 0.006508f
C258 B.n221 VSUBS 0.006508f
C259 B.n222 VSUBS 0.006508f
C260 B.n223 VSUBS 0.006508f
C261 B.n224 VSUBS 0.006125f
C262 B.n225 VSUBS 0.015077f
C263 B.n226 VSUBS 0.003637f
C264 B.n227 VSUBS 0.006508f
C265 B.n228 VSUBS 0.006508f
C266 B.n229 VSUBS 0.006508f
C267 B.n230 VSUBS 0.006508f
C268 B.n231 VSUBS 0.006508f
C269 B.n232 VSUBS 0.006508f
C270 B.n233 VSUBS 0.006508f
C271 B.n234 VSUBS 0.006508f
C272 B.n235 VSUBS 0.006508f
C273 B.n236 VSUBS 0.006508f
C274 B.n237 VSUBS 0.006508f
C275 B.n238 VSUBS 0.006508f
C276 B.t5 VSUBS 0.073917f
C277 B.t4 VSUBS 0.087348f
C278 B.t3 VSUBS 0.308f
C279 B.n239 VSUBS 0.154721f
C280 B.n240 VSUBS 0.129691f
C281 B.n241 VSUBS 0.015077f
C282 B.n242 VSUBS 0.003637f
C283 B.n243 VSUBS 0.006508f
C284 B.n244 VSUBS 0.006508f
C285 B.n245 VSUBS 0.006508f
C286 B.n246 VSUBS 0.006508f
C287 B.n247 VSUBS 0.006508f
C288 B.n248 VSUBS 0.006508f
C289 B.n249 VSUBS 0.006508f
C290 B.n250 VSUBS 0.006508f
C291 B.n251 VSUBS 0.006508f
C292 B.n252 VSUBS 0.006508f
C293 B.n253 VSUBS 0.006508f
C294 B.n254 VSUBS 0.006508f
C295 B.n255 VSUBS 0.006508f
C296 B.n256 VSUBS 0.006508f
C297 B.n257 VSUBS 0.006508f
C298 B.n258 VSUBS 0.006508f
C299 B.n259 VSUBS 0.006508f
C300 B.n260 VSUBS 0.006508f
C301 B.n261 VSUBS 0.006508f
C302 B.n262 VSUBS 0.006508f
C303 B.n263 VSUBS 0.006508f
C304 B.n264 VSUBS 0.006508f
C305 B.n265 VSUBS 0.006508f
C306 B.n266 VSUBS 0.006508f
C307 B.n267 VSUBS 0.006508f
C308 B.n268 VSUBS 0.006508f
C309 B.n269 VSUBS 0.006508f
C310 B.n270 VSUBS 0.006508f
C311 B.n271 VSUBS 0.006508f
C312 B.n272 VSUBS 0.006508f
C313 B.n273 VSUBS 0.006508f
C314 B.n274 VSUBS 0.006508f
C315 B.n275 VSUBS 0.015822f
C316 B.n276 VSUBS 0.015067f
C317 B.n277 VSUBS 0.015748f
C318 B.n278 VSUBS 0.006508f
C319 B.n279 VSUBS 0.006508f
C320 B.n280 VSUBS 0.006508f
C321 B.n281 VSUBS 0.006508f
C322 B.n282 VSUBS 0.006508f
C323 B.n283 VSUBS 0.006508f
C324 B.n284 VSUBS 0.006508f
C325 B.n285 VSUBS 0.006508f
C326 B.n286 VSUBS 0.006508f
C327 B.n287 VSUBS 0.006508f
C328 B.n288 VSUBS 0.006508f
C329 B.n289 VSUBS 0.006508f
C330 B.n290 VSUBS 0.006508f
C331 B.n291 VSUBS 0.006508f
C332 B.n292 VSUBS 0.006508f
C333 B.n293 VSUBS 0.006508f
C334 B.n294 VSUBS 0.006508f
C335 B.n295 VSUBS 0.006508f
C336 B.n296 VSUBS 0.006508f
C337 B.n297 VSUBS 0.006508f
C338 B.n298 VSUBS 0.006508f
C339 B.n299 VSUBS 0.006508f
C340 B.n300 VSUBS 0.006508f
C341 B.n301 VSUBS 0.006508f
C342 B.n302 VSUBS 0.006508f
C343 B.n303 VSUBS 0.006508f
C344 B.n304 VSUBS 0.006508f
C345 B.n305 VSUBS 0.006508f
C346 B.n306 VSUBS 0.006508f
C347 B.n307 VSUBS 0.006508f
C348 B.n308 VSUBS 0.006508f
C349 B.n309 VSUBS 0.006508f
C350 B.n310 VSUBS 0.006508f
C351 B.n311 VSUBS 0.006508f
C352 B.n312 VSUBS 0.006508f
C353 B.n313 VSUBS 0.006508f
C354 B.n314 VSUBS 0.006508f
C355 B.n315 VSUBS 0.006508f
C356 B.n316 VSUBS 0.006508f
C357 B.n317 VSUBS 0.006508f
C358 B.n318 VSUBS 0.006508f
C359 B.n319 VSUBS 0.006508f
C360 B.n320 VSUBS 0.006508f
C361 B.n321 VSUBS 0.006508f
C362 B.n322 VSUBS 0.006508f
C363 B.n323 VSUBS 0.006508f
C364 B.n324 VSUBS 0.006508f
C365 B.n325 VSUBS 0.006508f
C366 B.n326 VSUBS 0.006508f
C367 B.n327 VSUBS 0.006508f
C368 B.n328 VSUBS 0.006508f
C369 B.n329 VSUBS 0.006508f
C370 B.n330 VSUBS 0.006508f
C371 B.n331 VSUBS 0.006508f
C372 B.n332 VSUBS 0.006508f
C373 B.n333 VSUBS 0.006508f
C374 B.n334 VSUBS 0.006508f
C375 B.n335 VSUBS 0.006508f
C376 B.n336 VSUBS 0.006508f
C377 B.n337 VSUBS 0.006508f
C378 B.n338 VSUBS 0.006508f
C379 B.n339 VSUBS 0.006508f
C380 B.n340 VSUBS 0.006508f
C381 B.n341 VSUBS 0.006508f
C382 B.n342 VSUBS 0.006508f
C383 B.n343 VSUBS 0.006508f
C384 B.n344 VSUBS 0.006508f
C385 B.n345 VSUBS 0.006508f
C386 B.n346 VSUBS 0.006508f
C387 B.n347 VSUBS 0.006508f
C388 B.n348 VSUBS 0.006508f
C389 B.n349 VSUBS 0.006508f
C390 B.n350 VSUBS 0.006508f
C391 B.n351 VSUBS 0.006508f
C392 B.n352 VSUBS 0.006508f
C393 B.n353 VSUBS 0.006508f
C394 B.n354 VSUBS 0.006508f
C395 B.n355 VSUBS 0.006508f
C396 B.n356 VSUBS 0.006508f
C397 B.n357 VSUBS 0.006508f
C398 B.n358 VSUBS 0.006508f
C399 B.n359 VSUBS 0.006508f
C400 B.n360 VSUBS 0.006508f
C401 B.n361 VSUBS 0.006508f
C402 B.n362 VSUBS 0.006508f
C403 B.n363 VSUBS 0.006508f
C404 B.n364 VSUBS 0.006508f
C405 B.n365 VSUBS 0.006508f
C406 B.n366 VSUBS 0.006508f
C407 B.n367 VSUBS 0.006508f
C408 B.n368 VSUBS 0.006508f
C409 B.n369 VSUBS 0.006508f
C410 B.n370 VSUBS 0.006508f
C411 B.n371 VSUBS 0.006508f
C412 B.n372 VSUBS 0.006508f
C413 B.n373 VSUBS 0.006508f
C414 B.n374 VSUBS 0.006508f
C415 B.n375 VSUBS 0.006508f
C416 B.n376 VSUBS 0.006508f
C417 B.n377 VSUBS 0.006508f
C418 B.n378 VSUBS 0.006508f
C419 B.n379 VSUBS 0.006508f
C420 B.n380 VSUBS 0.006508f
C421 B.n381 VSUBS 0.006508f
C422 B.n382 VSUBS 0.006508f
C423 B.n383 VSUBS 0.006508f
C424 B.n384 VSUBS 0.006508f
C425 B.n385 VSUBS 0.006508f
C426 B.n386 VSUBS 0.006508f
C427 B.n387 VSUBS 0.006508f
C428 B.n388 VSUBS 0.006508f
C429 B.n389 VSUBS 0.014993f
C430 B.n390 VSUBS 0.014993f
C431 B.n391 VSUBS 0.015822f
C432 B.n392 VSUBS 0.006508f
C433 B.n393 VSUBS 0.006508f
C434 B.n394 VSUBS 0.006508f
C435 B.n395 VSUBS 0.006508f
C436 B.n396 VSUBS 0.006508f
C437 B.n397 VSUBS 0.006508f
C438 B.n398 VSUBS 0.006508f
C439 B.n399 VSUBS 0.006508f
C440 B.n400 VSUBS 0.006508f
C441 B.n401 VSUBS 0.006508f
C442 B.n402 VSUBS 0.006508f
C443 B.n403 VSUBS 0.006508f
C444 B.n404 VSUBS 0.006508f
C445 B.n405 VSUBS 0.006508f
C446 B.n406 VSUBS 0.006508f
C447 B.n407 VSUBS 0.006508f
C448 B.n408 VSUBS 0.006508f
C449 B.n409 VSUBS 0.006508f
C450 B.n410 VSUBS 0.006508f
C451 B.n411 VSUBS 0.006508f
C452 B.n412 VSUBS 0.006508f
C453 B.n413 VSUBS 0.006508f
C454 B.n414 VSUBS 0.006508f
C455 B.n415 VSUBS 0.006508f
C456 B.n416 VSUBS 0.006508f
C457 B.n417 VSUBS 0.006508f
C458 B.n418 VSUBS 0.006508f
C459 B.n419 VSUBS 0.006508f
C460 B.n420 VSUBS 0.006508f
C461 B.n421 VSUBS 0.006508f
C462 B.n422 VSUBS 0.006125f
C463 B.n423 VSUBS 0.006508f
C464 B.n424 VSUBS 0.006508f
C465 B.n425 VSUBS 0.006508f
C466 B.n426 VSUBS 0.006508f
C467 B.n427 VSUBS 0.006508f
C468 B.n428 VSUBS 0.006508f
C469 B.n429 VSUBS 0.006508f
C470 B.n430 VSUBS 0.006508f
C471 B.n431 VSUBS 0.006508f
C472 B.n432 VSUBS 0.006508f
C473 B.n433 VSUBS 0.006508f
C474 B.n434 VSUBS 0.006508f
C475 B.n435 VSUBS 0.006508f
C476 B.n436 VSUBS 0.006508f
C477 B.n437 VSUBS 0.006508f
C478 B.n438 VSUBS 0.003637f
C479 B.n439 VSUBS 0.015077f
C480 B.n440 VSUBS 0.006125f
C481 B.n441 VSUBS 0.006508f
C482 B.n442 VSUBS 0.006508f
C483 B.n443 VSUBS 0.006508f
C484 B.n444 VSUBS 0.006508f
C485 B.n445 VSUBS 0.006508f
C486 B.n446 VSUBS 0.006508f
C487 B.n447 VSUBS 0.006508f
C488 B.n448 VSUBS 0.006508f
C489 B.n449 VSUBS 0.006508f
C490 B.n450 VSUBS 0.006508f
C491 B.n451 VSUBS 0.006508f
C492 B.n452 VSUBS 0.006508f
C493 B.n453 VSUBS 0.006508f
C494 B.n454 VSUBS 0.006508f
C495 B.n455 VSUBS 0.006508f
C496 B.n456 VSUBS 0.006508f
C497 B.n457 VSUBS 0.006508f
C498 B.n458 VSUBS 0.006508f
C499 B.n459 VSUBS 0.006508f
C500 B.n460 VSUBS 0.006508f
C501 B.n461 VSUBS 0.006508f
C502 B.n462 VSUBS 0.006508f
C503 B.n463 VSUBS 0.006508f
C504 B.n464 VSUBS 0.006508f
C505 B.n465 VSUBS 0.006508f
C506 B.n466 VSUBS 0.006508f
C507 B.n467 VSUBS 0.006508f
C508 B.n468 VSUBS 0.006508f
C509 B.n469 VSUBS 0.006508f
C510 B.n470 VSUBS 0.006508f
C511 B.n471 VSUBS 0.015822f
C512 B.n472 VSUBS 0.015822f
C513 B.n473 VSUBS 0.014993f
C514 B.n474 VSUBS 0.006508f
C515 B.n475 VSUBS 0.006508f
C516 B.n476 VSUBS 0.006508f
C517 B.n477 VSUBS 0.006508f
C518 B.n478 VSUBS 0.006508f
C519 B.n479 VSUBS 0.006508f
C520 B.n480 VSUBS 0.006508f
C521 B.n481 VSUBS 0.006508f
C522 B.n482 VSUBS 0.006508f
C523 B.n483 VSUBS 0.006508f
C524 B.n484 VSUBS 0.006508f
C525 B.n485 VSUBS 0.006508f
C526 B.n486 VSUBS 0.006508f
C527 B.n487 VSUBS 0.006508f
C528 B.n488 VSUBS 0.006508f
C529 B.n489 VSUBS 0.006508f
C530 B.n490 VSUBS 0.006508f
C531 B.n491 VSUBS 0.006508f
C532 B.n492 VSUBS 0.006508f
C533 B.n493 VSUBS 0.006508f
C534 B.n494 VSUBS 0.006508f
C535 B.n495 VSUBS 0.006508f
C536 B.n496 VSUBS 0.006508f
C537 B.n497 VSUBS 0.006508f
C538 B.n498 VSUBS 0.006508f
C539 B.n499 VSUBS 0.006508f
C540 B.n500 VSUBS 0.006508f
C541 B.n501 VSUBS 0.006508f
C542 B.n502 VSUBS 0.006508f
C543 B.n503 VSUBS 0.006508f
C544 B.n504 VSUBS 0.006508f
C545 B.n505 VSUBS 0.006508f
C546 B.n506 VSUBS 0.006508f
C547 B.n507 VSUBS 0.006508f
C548 B.n508 VSUBS 0.006508f
C549 B.n509 VSUBS 0.006508f
C550 B.n510 VSUBS 0.006508f
C551 B.n511 VSUBS 0.006508f
C552 B.n512 VSUBS 0.006508f
C553 B.n513 VSUBS 0.006508f
C554 B.n514 VSUBS 0.006508f
C555 B.n515 VSUBS 0.006508f
C556 B.n516 VSUBS 0.006508f
C557 B.n517 VSUBS 0.006508f
C558 B.n518 VSUBS 0.006508f
C559 B.n519 VSUBS 0.006508f
C560 B.n520 VSUBS 0.006508f
C561 B.n521 VSUBS 0.006508f
C562 B.n522 VSUBS 0.006508f
C563 B.n523 VSUBS 0.006508f
C564 B.n524 VSUBS 0.006508f
C565 B.n525 VSUBS 0.006508f
C566 B.n526 VSUBS 0.006508f
C567 B.n527 VSUBS 0.008492f
C568 B.n528 VSUBS 0.009046f
C569 B.n529 VSUBS 0.017989f
C570 VDD1.n0 VSUBS 0.026291f
C571 VDD1.n1 VSUBS 0.023297f
C572 VDD1.n2 VSUBS 0.012519f
C573 VDD1.n3 VSUBS 0.02959f
C574 VDD1.n4 VSUBS 0.013255f
C575 VDD1.n5 VSUBS 0.023297f
C576 VDD1.n6 VSUBS 0.012519f
C577 VDD1.n7 VSUBS 0.022192f
C578 VDD1.n8 VSUBS 0.018796f
C579 VDD1.t1 VSUBS 0.064067f
C580 VDD1.n9 VSUBS 0.099429f
C581 VDD1.n10 VSUBS 0.469824f
C582 VDD1.n11 VSUBS 0.012519f
C583 VDD1.n12 VSUBS 0.013255f
C584 VDD1.n13 VSUBS 0.02959f
C585 VDD1.n14 VSUBS 0.02959f
C586 VDD1.n15 VSUBS 0.013255f
C587 VDD1.n16 VSUBS 0.012519f
C588 VDD1.n17 VSUBS 0.023297f
C589 VDD1.n18 VSUBS 0.023297f
C590 VDD1.n19 VSUBS 0.012519f
C591 VDD1.n20 VSUBS 0.013255f
C592 VDD1.n21 VSUBS 0.02959f
C593 VDD1.n22 VSUBS 0.073993f
C594 VDD1.n23 VSUBS 0.013255f
C595 VDD1.n24 VSUBS 0.012519f
C596 VDD1.n25 VSUBS 0.057669f
C597 VDD1.n26 VSUBS 0.05773f
C598 VDD1.t2 VSUBS 0.099414f
C599 VDD1.t3 VSUBS 0.099414f
C600 VDD1.n27 VSUBS 0.640893f
C601 VDD1.n28 VSUBS 0.654661f
C602 VDD1.n29 VSUBS 0.026291f
C603 VDD1.n30 VSUBS 0.023297f
C604 VDD1.n31 VSUBS 0.012519f
C605 VDD1.n32 VSUBS 0.02959f
C606 VDD1.n33 VSUBS 0.013255f
C607 VDD1.n34 VSUBS 0.023297f
C608 VDD1.n35 VSUBS 0.012519f
C609 VDD1.n36 VSUBS 0.022192f
C610 VDD1.n37 VSUBS 0.018796f
C611 VDD1.t5 VSUBS 0.064067f
C612 VDD1.n38 VSUBS 0.099429f
C613 VDD1.n39 VSUBS 0.469824f
C614 VDD1.n40 VSUBS 0.012519f
C615 VDD1.n41 VSUBS 0.013255f
C616 VDD1.n42 VSUBS 0.02959f
C617 VDD1.n43 VSUBS 0.02959f
C618 VDD1.n44 VSUBS 0.013255f
C619 VDD1.n45 VSUBS 0.012519f
C620 VDD1.n46 VSUBS 0.023297f
C621 VDD1.n47 VSUBS 0.023297f
C622 VDD1.n48 VSUBS 0.012519f
C623 VDD1.n49 VSUBS 0.013255f
C624 VDD1.n50 VSUBS 0.02959f
C625 VDD1.n51 VSUBS 0.073993f
C626 VDD1.n52 VSUBS 0.013255f
C627 VDD1.n53 VSUBS 0.012519f
C628 VDD1.n54 VSUBS 0.057669f
C629 VDD1.n55 VSUBS 0.05773f
C630 VDD1.t4 VSUBS 0.099414f
C631 VDD1.t0 VSUBS 0.099414f
C632 VDD1.n56 VSUBS 0.64089f
C633 VDD1.n57 VSUBS 0.647915f
C634 VDD1.t9 VSUBS 0.099414f
C635 VDD1.t6 VSUBS 0.099414f
C636 VDD1.n58 VSUBS 0.64658f
C637 VDD1.n59 VSUBS 1.97791f
C638 VDD1.t8 VSUBS 0.099414f
C639 VDD1.t7 VSUBS 0.099414f
C640 VDD1.n60 VSUBS 0.64089f
C641 VDD1.n61 VSUBS 2.16102f
C642 VP.n0 VSUBS 0.049463f
C643 VP.t3 VSUBS 0.941127f
C644 VP.n1 VSUBS 0.082631f
C645 VP.n2 VSUBS 0.049463f
C646 VP.t9 VSUBS 0.941127f
C647 VP.n3 VSUBS 0.426072f
C648 VP.n4 VSUBS 0.049463f
C649 VP.t5 VSUBS 0.941127f
C650 VP.n5 VSUBS 0.37963f
C651 VP.n6 VSUBS 0.049463f
C652 VP.t4 VSUBS 0.941127f
C653 VP.n7 VSUBS 0.482631f
C654 VP.n8 VSUBS 0.049463f
C655 VP.t2 VSUBS 0.941127f
C656 VP.n9 VSUBS 0.082631f
C657 VP.n10 VSUBS 0.049463f
C658 VP.t6 VSUBS 0.941127f
C659 VP.n11 VSUBS 0.426072f
C660 VP.n12 VSUBS 0.049463f
C661 VP.t7 VSUBS 0.941127f
C662 VP.n13 VSUBS 0.453619f
C663 VP.t8 VSUBS 1.07768f
C664 VP.n14 VSUBS 0.480388f
C665 VP.n15 VSUBS 0.265542f
C666 VP.n16 VSUBS 0.061838f
C667 VP.n17 VSUBS 0.06027f
C668 VP.n18 VSUBS 0.083534f
C669 VP.n19 VSUBS 0.049463f
C670 VP.n20 VSUBS 0.049463f
C671 VP.n21 VSUBS 0.049463f
C672 VP.n22 VSUBS 0.083534f
C673 VP.n23 VSUBS 0.06027f
C674 VP.t1 VSUBS 0.941127f
C675 VP.n24 VSUBS 0.37963f
C676 VP.n25 VSUBS 0.061838f
C677 VP.n26 VSUBS 0.049463f
C678 VP.n27 VSUBS 0.049463f
C679 VP.n28 VSUBS 0.049463f
C680 VP.n29 VSUBS 0.039965f
C681 VP.n30 VSUBS 0.083046f
C682 VP.n31 VSUBS 0.482631f
C683 VP.n32 VSUBS 1.98622f
C684 VP.n33 VSUBS 2.02945f
C685 VP.n34 VSUBS 0.049463f
C686 VP.n35 VSUBS 0.083046f
C687 VP.n36 VSUBS 0.039965f
C688 VP.n37 VSUBS 0.082631f
C689 VP.n38 VSUBS 0.049463f
C690 VP.n39 VSUBS 0.049463f
C691 VP.n40 VSUBS 0.061838f
C692 VP.n41 VSUBS 0.06027f
C693 VP.n42 VSUBS 0.083534f
C694 VP.n43 VSUBS 0.049463f
C695 VP.n44 VSUBS 0.049463f
C696 VP.n45 VSUBS 0.049463f
C697 VP.n46 VSUBS 0.083534f
C698 VP.n47 VSUBS 0.06027f
C699 VP.t0 VSUBS 0.941127f
C700 VP.n48 VSUBS 0.37963f
C701 VP.n49 VSUBS 0.061838f
C702 VP.n50 VSUBS 0.049463f
C703 VP.n51 VSUBS 0.049463f
C704 VP.n52 VSUBS 0.049463f
C705 VP.n53 VSUBS 0.039965f
C706 VP.n54 VSUBS 0.083046f
C707 VP.n55 VSUBS 0.482631f
C708 VP.n56 VSUBS 0.043357f
C709 VTAIL.t13 VSUBS 0.128317f
C710 VTAIL.t17 VSUBS 0.128317f
C711 VTAIL.n0 VSUBS 0.733846f
C712 VTAIL.n1 VSUBS 0.748275f
C713 VTAIL.n2 VSUBS 0.033935f
C714 VTAIL.n3 VSUBS 0.03007f
C715 VTAIL.n4 VSUBS 0.016158f
C716 VTAIL.n5 VSUBS 0.038192f
C717 VTAIL.n6 VSUBS 0.017109f
C718 VTAIL.n7 VSUBS 0.03007f
C719 VTAIL.n8 VSUBS 0.016158f
C720 VTAIL.n9 VSUBS 0.028644f
C721 VTAIL.n10 VSUBS 0.02426f
C722 VTAIL.t5 VSUBS 0.082693f
C723 VTAIL.n11 VSUBS 0.128336f
C724 VTAIL.n12 VSUBS 0.606415f
C725 VTAIL.n13 VSUBS 0.016158f
C726 VTAIL.n14 VSUBS 0.017109f
C727 VTAIL.n15 VSUBS 0.038192f
C728 VTAIL.n16 VSUBS 0.038192f
C729 VTAIL.n17 VSUBS 0.017109f
C730 VTAIL.n18 VSUBS 0.016158f
C731 VTAIL.n19 VSUBS 0.03007f
C732 VTAIL.n20 VSUBS 0.03007f
C733 VTAIL.n21 VSUBS 0.016158f
C734 VTAIL.n22 VSUBS 0.017109f
C735 VTAIL.n23 VSUBS 0.038192f
C736 VTAIL.n24 VSUBS 0.095505f
C737 VTAIL.n25 VSUBS 0.017109f
C738 VTAIL.n26 VSUBS 0.016158f
C739 VTAIL.n27 VSUBS 0.074435f
C740 VTAIL.n28 VSUBS 0.048311f
C741 VTAIL.n29 VSUBS 0.28323f
C742 VTAIL.t6 VSUBS 0.128317f
C743 VTAIL.t1 VSUBS 0.128317f
C744 VTAIL.n30 VSUBS 0.733846f
C745 VTAIL.n31 VSUBS 0.801733f
C746 VTAIL.t2 VSUBS 0.128317f
C747 VTAIL.t9 VSUBS 0.128317f
C748 VTAIL.n32 VSUBS 0.733846f
C749 VTAIL.n33 VSUBS 1.80074f
C750 VTAIL.t10 VSUBS 0.128317f
C751 VTAIL.t11 VSUBS 0.128317f
C752 VTAIL.n34 VSUBS 0.733851f
C753 VTAIL.n35 VSUBS 1.80074f
C754 VTAIL.t14 VSUBS 0.128317f
C755 VTAIL.t15 VSUBS 0.128317f
C756 VTAIL.n36 VSUBS 0.733851f
C757 VTAIL.n37 VSUBS 0.801728f
C758 VTAIL.n38 VSUBS 0.033935f
C759 VTAIL.n39 VSUBS 0.03007f
C760 VTAIL.n40 VSUBS 0.016158f
C761 VTAIL.n41 VSUBS 0.038192f
C762 VTAIL.n42 VSUBS 0.017109f
C763 VTAIL.n43 VSUBS 0.03007f
C764 VTAIL.n44 VSUBS 0.016158f
C765 VTAIL.n45 VSUBS 0.028644f
C766 VTAIL.n46 VSUBS 0.02426f
C767 VTAIL.t16 VSUBS 0.082693f
C768 VTAIL.n47 VSUBS 0.128336f
C769 VTAIL.n48 VSUBS 0.606415f
C770 VTAIL.n49 VSUBS 0.016158f
C771 VTAIL.n50 VSUBS 0.017109f
C772 VTAIL.n51 VSUBS 0.038192f
C773 VTAIL.n52 VSUBS 0.038192f
C774 VTAIL.n53 VSUBS 0.017109f
C775 VTAIL.n54 VSUBS 0.016158f
C776 VTAIL.n55 VSUBS 0.03007f
C777 VTAIL.n56 VSUBS 0.03007f
C778 VTAIL.n57 VSUBS 0.016158f
C779 VTAIL.n58 VSUBS 0.017109f
C780 VTAIL.n59 VSUBS 0.038192f
C781 VTAIL.n60 VSUBS 0.095505f
C782 VTAIL.n61 VSUBS 0.017109f
C783 VTAIL.n62 VSUBS 0.016158f
C784 VTAIL.n63 VSUBS 0.074435f
C785 VTAIL.n64 VSUBS 0.048311f
C786 VTAIL.n65 VSUBS 0.28323f
C787 VTAIL.t7 VSUBS 0.128317f
C788 VTAIL.t8 VSUBS 0.128317f
C789 VTAIL.n66 VSUBS 0.733851f
C790 VTAIL.n67 VSUBS 0.777505f
C791 VTAIL.t0 VSUBS 0.128317f
C792 VTAIL.t3 VSUBS 0.128317f
C793 VTAIL.n68 VSUBS 0.733851f
C794 VTAIL.n69 VSUBS 0.801728f
C795 VTAIL.n70 VSUBS 0.033935f
C796 VTAIL.n71 VSUBS 0.03007f
C797 VTAIL.n72 VSUBS 0.016158f
C798 VTAIL.n73 VSUBS 0.038192f
C799 VTAIL.n74 VSUBS 0.017109f
C800 VTAIL.n75 VSUBS 0.03007f
C801 VTAIL.n76 VSUBS 0.016158f
C802 VTAIL.n77 VSUBS 0.028644f
C803 VTAIL.n78 VSUBS 0.02426f
C804 VTAIL.t4 VSUBS 0.082693f
C805 VTAIL.n79 VSUBS 0.128336f
C806 VTAIL.n80 VSUBS 0.606415f
C807 VTAIL.n81 VSUBS 0.016158f
C808 VTAIL.n82 VSUBS 0.017109f
C809 VTAIL.n83 VSUBS 0.038192f
C810 VTAIL.n84 VSUBS 0.038192f
C811 VTAIL.n85 VSUBS 0.017109f
C812 VTAIL.n86 VSUBS 0.016158f
C813 VTAIL.n87 VSUBS 0.03007f
C814 VTAIL.n88 VSUBS 0.03007f
C815 VTAIL.n89 VSUBS 0.016158f
C816 VTAIL.n90 VSUBS 0.017109f
C817 VTAIL.n91 VSUBS 0.038192f
C818 VTAIL.n92 VSUBS 0.095505f
C819 VTAIL.n93 VSUBS 0.017109f
C820 VTAIL.n94 VSUBS 0.016158f
C821 VTAIL.n95 VSUBS 0.074435f
C822 VTAIL.n96 VSUBS 0.048311f
C823 VTAIL.n97 VSUBS 1.16697f
C824 VTAIL.n98 VSUBS 0.033935f
C825 VTAIL.n99 VSUBS 0.03007f
C826 VTAIL.n100 VSUBS 0.016158f
C827 VTAIL.n101 VSUBS 0.038192f
C828 VTAIL.n102 VSUBS 0.017109f
C829 VTAIL.n103 VSUBS 0.03007f
C830 VTAIL.n104 VSUBS 0.016158f
C831 VTAIL.n105 VSUBS 0.028644f
C832 VTAIL.n106 VSUBS 0.02426f
C833 VTAIL.t12 VSUBS 0.082693f
C834 VTAIL.n107 VSUBS 0.128336f
C835 VTAIL.n108 VSUBS 0.606415f
C836 VTAIL.n109 VSUBS 0.016158f
C837 VTAIL.n110 VSUBS 0.017109f
C838 VTAIL.n111 VSUBS 0.038192f
C839 VTAIL.n112 VSUBS 0.038192f
C840 VTAIL.n113 VSUBS 0.017109f
C841 VTAIL.n114 VSUBS 0.016158f
C842 VTAIL.n115 VSUBS 0.03007f
C843 VTAIL.n116 VSUBS 0.03007f
C844 VTAIL.n117 VSUBS 0.016158f
C845 VTAIL.n118 VSUBS 0.017109f
C846 VTAIL.n119 VSUBS 0.038192f
C847 VTAIL.n120 VSUBS 0.095505f
C848 VTAIL.n121 VSUBS 0.017109f
C849 VTAIL.n122 VSUBS 0.016158f
C850 VTAIL.n123 VSUBS 0.074435f
C851 VTAIL.n124 VSUBS 0.048311f
C852 VTAIL.n125 VSUBS 1.16697f
C853 VTAIL.t18 VSUBS 0.128317f
C854 VTAIL.t19 VSUBS 0.128317f
C855 VTAIL.n126 VSUBS 0.733846f
C856 VTAIL.n127 VSUBS 0.691476f
C857 VDD2.n0 VSUBS 0.026026f
C858 VDD2.n1 VSUBS 0.023062f
C859 VDD2.n2 VSUBS 0.012393f
C860 VDD2.n3 VSUBS 0.029292f
C861 VDD2.n4 VSUBS 0.013122f
C862 VDD2.n5 VSUBS 0.023062f
C863 VDD2.n6 VSUBS 0.012393f
C864 VDD2.n7 VSUBS 0.021969f
C865 VDD2.n8 VSUBS 0.018606f
C866 VDD2.t7 VSUBS 0.063422f
C867 VDD2.n9 VSUBS 0.098428f
C868 VDD2.n10 VSUBS 0.465092f
C869 VDD2.n11 VSUBS 0.012393f
C870 VDD2.n12 VSUBS 0.013122f
C871 VDD2.n13 VSUBS 0.029292f
C872 VDD2.n14 VSUBS 0.029292f
C873 VDD2.n15 VSUBS 0.013122f
C874 VDD2.n16 VSUBS 0.012393f
C875 VDD2.n17 VSUBS 0.023062f
C876 VDD2.n18 VSUBS 0.023062f
C877 VDD2.n19 VSUBS 0.012393f
C878 VDD2.n20 VSUBS 0.013122f
C879 VDD2.n21 VSUBS 0.029292f
C880 VDD2.n22 VSUBS 0.073248f
C881 VDD2.n23 VSUBS 0.013122f
C882 VDD2.n24 VSUBS 0.012393f
C883 VDD2.n25 VSUBS 0.057088f
C884 VDD2.n26 VSUBS 0.057149f
C885 VDD2.t6 VSUBS 0.098413f
C886 VDD2.t0 VSUBS 0.098413f
C887 VDD2.n27 VSUBS 0.634435f
C888 VDD2.n28 VSUBS 0.641389f
C889 VDD2.t3 VSUBS 0.098413f
C890 VDD2.t9 VSUBS 0.098413f
C891 VDD2.n29 VSUBS 0.640068f
C892 VDD2.n30 VSUBS 1.87635f
C893 VDD2.n31 VSUBS 0.026026f
C894 VDD2.n32 VSUBS 0.023062f
C895 VDD2.n33 VSUBS 0.012393f
C896 VDD2.n34 VSUBS 0.029292f
C897 VDD2.n35 VSUBS 0.013122f
C898 VDD2.n36 VSUBS 0.023062f
C899 VDD2.n37 VSUBS 0.012393f
C900 VDD2.n38 VSUBS 0.021969f
C901 VDD2.n39 VSUBS 0.018606f
C902 VDD2.t5 VSUBS 0.063422f
C903 VDD2.n40 VSUBS 0.098428f
C904 VDD2.n41 VSUBS 0.465092f
C905 VDD2.n42 VSUBS 0.012393f
C906 VDD2.n43 VSUBS 0.013122f
C907 VDD2.n44 VSUBS 0.029292f
C908 VDD2.n45 VSUBS 0.029292f
C909 VDD2.n46 VSUBS 0.013122f
C910 VDD2.n47 VSUBS 0.012393f
C911 VDD2.n48 VSUBS 0.023062f
C912 VDD2.n49 VSUBS 0.023062f
C913 VDD2.n50 VSUBS 0.012393f
C914 VDD2.n51 VSUBS 0.013122f
C915 VDD2.n52 VSUBS 0.029292f
C916 VDD2.n53 VSUBS 0.073248f
C917 VDD2.n54 VSUBS 0.013122f
C918 VDD2.n55 VSUBS 0.012393f
C919 VDD2.n56 VSUBS 0.057088f
C920 VDD2.n57 VSUBS 0.052949f
C921 VDD2.n58 VSUBS 1.73642f
C922 VDD2.t4 VSUBS 0.098413f
C923 VDD2.t8 VSUBS 0.098413f
C924 VDD2.n59 VSUBS 0.634438f
C925 VDD2.n60 VSUBS 0.498711f
C926 VDD2.t2 VSUBS 0.098413f
C927 VDD2.t1 VSUBS 0.098413f
C928 VDD2.n61 VSUBS 0.640045f
C929 VN.n0 VSUBS 0.047876f
C930 VN.t7 VSUBS 0.910934f
C931 VN.n1 VSUBS 0.07998f
C932 VN.n2 VSUBS 0.047876f
C933 VN.t1 VSUBS 0.910934f
C934 VN.n3 VSUBS 0.412403f
C935 VN.n4 VSUBS 0.047876f
C936 VN.t2 VSUBS 0.910934f
C937 VN.n5 VSUBS 0.439066f
C938 VN.t6 VSUBS 1.04311f
C939 VN.n6 VSUBS 0.464976f
C940 VN.n7 VSUBS 0.257023f
C941 VN.n8 VSUBS 0.059854f
C942 VN.n9 VSUBS 0.058336f
C943 VN.n10 VSUBS 0.080855f
C944 VN.n11 VSUBS 0.047876f
C945 VN.n12 VSUBS 0.047876f
C946 VN.n13 VSUBS 0.047876f
C947 VN.n14 VSUBS 0.080855f
C948 VN.n15 VSUBS 0.058336f
C949 VN.t0 VSUBS 0.910934f
C950 VN.n16 VSUBS 0.367451f
C951 VN.n17 VSUBS 0.059854f
C952 VN.n18 VSUBS 0.047876f
C953 VN.n19 VSUBS 0.047876f
C954 VN.n20 VSUBS 0.047876f
C955 VN.n21 VSUBS 0.038683f
C956 VN.n22 VSUBS 0.080382f
C957 VN.n23 VSUBS 0.467147f
C958 VN.n24 VSUBS 0.041966f
C959 VN.n25 VSUBS 0.047876f
C960 VN.t9 VSUBS 0.910934f
C961 VN.n26 VSUBS 0.07998f
C962 VN.n27 VSUBS 0.047876f
C963 VN.t8 VSUBS 0.910934f
C964 VN.n28 VSUBS 0.367451f
C965 VN.t5 VSUBS 0.910934f
C966 VN.n29 VSUBS 0.412403f
C967 VN.n30 VSUBS 0.047876f
C968 VN.t4 VSUBS 0.910934f
C969 VN.n31 VSUBS 0.439066f
C970 VN.t3 VSUBS 1.04311f
C971 VN.n32 VSUBS 0.464976f
C972 VN.n33 VSUBS 0.257023f
C973 VN.n34 VSUBS 0.059854f
C974 VN.n35 VSUBS 0.058336f
C975 VN.n36 VSUBS 0.080855f
C976 VN.n37 VSUBS 0.047876f
C977 VN.n38 VSUBS 0.047876f
C978 VN.n39 VSUBS 0.047876f
C979 VN.n40 VSUBS 0.080855f
C980 VN.n41 VSUBS 0.058336f
C981 VN.n42 VSUBS 0.059854f
C982 VN.n43 VSUBS 0.047876f
C983 VN.n44 VSUBS 0.047876f
C984 VN.n45 VSUBS 0.047876f
C985 VN.n46 VSUBS 0.038683f
C986 VN.n47 VSUBS 0.080382f
C987 VN.n48 VSUBS 0.467147f
C988 VN.n49 VSUBS 1.95397f
.ends

