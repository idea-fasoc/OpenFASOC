* NGSPICE file created from diff_pair_sample_0101.ext - technology: sky130A

.subckt diff_pair_sample_0101 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.4992 ps=3.34 w=1.28 l=2.73
X1 VTAIL.t3 VN.t0 VDD2.t3 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0.2112 ps=1.61 w=1.28 l=2.73
X2 B.t11 B.t9 B.t10 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0 ps=0 w=1.28 l=2.73
X3 VDD2.t2 VN.t1 VTAIL.t2 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.4992 ps=3.34 w=1.28 l=2.73
X4 VTAIL.t6 VP.t1 VDD1.t2 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0.2112 ps=1.61 w=1.28 l=2.73
X5 B.t8 B.t6 B.t7 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0 ps=0 w=1.28 l=2.73
X6 VTAIL.t1 VN.t2 VDD2.t1 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0.2112 ps=1.61 w=1.28 l=2.73
X7 B.t5 B.t3 B.t4 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0 ps=0 w=1.28 l=2.73
X8 VTAIL.t5 VP.t2 VDD1.t1 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0.2112 ps=1.61 w=1.28 l=2.73
X9 VDD1.t0 VP.t3 VTAIL.t4 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.4992 ps=3.34 w=1.28 l=2.73
X10 VDD2.t0 VN.t3 VTAIL.t0 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.2112 pd=1.61 as=0.4992 ps=3.34 w=1.28 l=2.73
X11 B.t2 B.t0 B.t1 w_n2806_n1224# sky130_fd_pr__pfet_01v8 ad=0.4992 pd=3.34 as=0 ps=0 w=1.28 l=2.73
R0 VP.n16 VP.n0 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n13 VP.n1 161.3
R3 VP.n12 VP.n11 161.3
R4 VP.n10 VP.n2 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n3 161.3
R7 VP.n6 VP.n5 109.433
R8 VP.n18 VP.n17 109.433
R9 VP.n4 VP.t2 45.6769
R10 VP.n4 VP.t0 44.8002
R11 VP.n6 VP.n4 42.1102
R12 VP.n11 VP.n10 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n9 VP.n3 24.5923
R15 VP.n10 VP.n9 24.5923
R16 VP.n15 VP.n1 24.5923
R17 VP.n16 VP.n15 24.5923
R18 VP.n5 VP.t1 11.3001
R19 VP.n17 VP.t3 11.3001
R20 VP.n5 VP.n3 1.47601
R21 VP.n17 VP.n16 1.47601
R22 VP.n7 VP.n6 0.278335
R23 VP.n18 VP.n0 0.278335
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153485
R31 VTAIL.n5 VTAIL.t5 372.7
R32 VTAIL.n4 VTAIL.t2 372.7
R33 VTAIL.n3 VTAIL.t1 372.7
R34 VTAIL.n7 VTAIL.t0 372.7
R35 VTAIL.n0 VTAIL.t3 372.7
R36 VTAIL.n1 VTAIL.t4 372.7
R37 VTAIL.n2 VTAIL.t6 372.7
R38 VTAIL.n6 VTAIL.t7 372.7
R39 VTAIL.n7 VTAIL.n6 16.1083
R40 VTAIL.n3 VTAIL.n2 16.1083
R41 VTAIL.n4 VTAIL.n3 2.63843
R42 VTAIL.n6 VTAIL.n5 2.63843
R43 VTAIL.n2 VTAIL.n1 2.63843
R44 VTAIL VTAIL.n0 1.37766
R45 VTAIL VTAIL.n7 1.26128
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 VDD1 VDD1.n1 379.699
R49 VDD1 VDD1.n0 346.5
R50 VDD1.n0 VDD1.t1 25.395
R51 VDD1.n0 VDD1.t3 25.395
R52 VDD1.n1 VDD1.t2 25.395
R53 VDD1.n1 VDD1.t0 25.395
R54 VN.n0 VN.t0 45.6769
R55 VN.n1 VN.t1 45.6769
R56 VN.n0 VN.t3 44.8002
R57 VN.n1 VN.t2 44.8002
R58 VN VN.n1 42.3891
R59 VN VN.n0 3.59742
R60 VDD2.n2 VDD2.n0 379.173
R61 VDD2.n2 VDD2.n1 346.442
R62 VDD2.n1 VDD2.t1 25.395
R63 VDD2.n1 VDD2.t2 25.395
R64 VDD2.n0 VDD2.t3 25.395
R65 VDD2.n0 VDD2.t0 25.395
R66 VDD2 VDD2.n2 0.0586897
R67 B.n316 B.n39 585
R68 B.n318 B.n317 585
R69 B.n319 B.n38 585
R70 B.n321 B.n320 585
R71 B.n322 B.n37 585
R72 B.n324 B.n323 585
R73 B.n325 B.n36 585
R74 B.n327 B.n326 585
R75 B.n328 B.n35 585
R76 B.n330 B.n329 585
R77 B.n332 B.n32 585
R78 B.n334 B.n333 585
R79 B.n335 B.n31 585
R80 B.n337 B.n336 585
R81 B.n338 B.n30 585
R82 B.n340 B.n339 585
R83 B.n341 B.n29 585
R84 B.n343 B.n342 585
R85 B.n344 B.n25 585
R86 B.n346 B.n345 585
R87 B.n347 B.n24 585
R88 B.n349 B.n348 585
R89 B.n350 B.n23 585
R90 B.n352 B.n351 585
R91 B.n353 B.n22 585
R92 B.n355 B.n354 585
R93 B.n356 B.n21 585
R94 B.n358 B.n357 585
R95 B.n359 B.n20 585
R96 B.n361 B.n360 585
R97 B.n315 B.n314 585
R98 B.n313 B.n40 585
R99 B.n312 B.n311 585
R100 B.n310 B.n41 585
R101 B.n309 B.n308 585
R102 B.n307 B.n42 585
R103 B.n306 B.n305 585
R104 B.n304 B.n43 585
R105 B.n303 B.n302 585
R106 B.n301 B.n44 585
R107 B.n300 B.n299 585
R108 B.n298 B.n45 585
R109 B.n297 B.n296 585
R110 B.n295 B.n46 585
R111 B.n294 B.n293 585
R112 B.n292 B.n47 585
R113 B.n291 B.n290 585
R114 B.n289 B.n48 585
R115 B.n288 B.n287 585
R116 B.n286 B.n49 585
R117 B.n285 B.n284 585
R118 B.n283 B.n50 585
R119 B.n282 B.n281 585
R120 B.n280 B.n51 585
R121 B.n279 B.n278 585
R122 B.n277 B.n52 585
R123 B.n276 B.n275 585
R124 B.n274 B.n53 585
R125 B.n273 B.n272 585
R126 B.n271 B.n54 585
R127 B.n270 B.n269 585
R128 B.n268 B.n55 585
R129 B.n267 B.n266 585
R130 B.n265 B.n56 585
R131 B.n264 B.n263 585
R132 B.n262 B.n57 585
R133 B.n261 B.n260 585
R134 B.n259 B.n58 585
R135 B.n258 B.n257 585
R136 B.n256 B.n59 585
R137 B.n255 B.n254 585
R138 B.n253 B.n60 585
R139 B.n252 B.n251 585
R140 B.n250 B.n61 585
R141 B.n249 B.n248 585
R142 B.n247 B.n62 585
R143 B.n246 B.n245 585
R144 B.n244 B.n63 585
R145 B.n243 B.n242 585
R146 B.n241 B.n64 585
R147 B.n240 B.n239 585
R148 B.n238 B.n65 585
R149 B.n237 B.n236 585
R150 B.n235 B.n66 585
R151 B.n234 B.n233 585
R152 B.n232 B.n67 585
R153 B.n231 B.n230 585
R154 B.n229 B.n68 585
R155 B.n228 B.n227 585
R156 B.n226 B.n69 585
R157 B.n225 B.n224 585
R158 B.n223 B.n70 585
R159 B.n222 B.n221 585
R160 B.n220 B.n71 585
R161 B.n219 B.n218 585
R162 B.n217 B.n72 585
R163 B.n216 B.n215 585
R164 B.n214 B.n73 585
R165 B.n213 B.n212 585
R166 B.n211 B.n74 585
R167 B.n210 B.n209 585
R168 B.n163 B.n94 585
R169 B.n165 B.n164 585
R170 B.n166 B.n93 585
R171 B.n168 B.n167 585
R172 B.n169 B.n92 585
R173 B.n171 B.n170 585
R174 B.n172 B.n91 585
R175 B.n174 B.n173 585
R176 B.n175 B.n90 585
R177 B.n177 B.n176 585
R178 B.n179 B.n178 585
R179 B.n180 B.n86 585
R180 B.n182 B.n181 585
R181 B.n183 B.n85 585
R182 B.n185 B.n184 585
R183 B.n186 B.n84 585
R184 B.n188 B.n187 585
R185 B.n189 B.n83 585
R186 B.n191 B.n190 585
R187 B.n192 B.n80 585
R188 B.n195 B.n194 585
R189 B.n196 B.n79 585
R190 B.n198 B.n197 585
R191 B.n199 B.n78 585
R192 B.n201 B.n200 585
R193 B.n202 B.n77 585
R194 B.n204 B.n203 585
R195 B.n205 B.n76 585
R196 B.n207 B.n206 585
R197 B.n208 B.n75 585
R198 B.n162 B.n161 585
R199 B.n160 B.n95 585
R200 B.n159 B.n158 585
R201 B.n157 B.n96 585
R202 B.n156 B.n155 585
R203 B.n154 B.n97 585
R204 B.n153 B.n152 585
R205 B.n151 B.n98 585
R206 B.n150 B.n149 585
R207 B.n148 B.n99 585
R208 B.n147 B.n146 585
R209 B.n145 B.n100 585
R210 B.n144 B.n143 585
R211 B.n142 B.n101 585
R212 B.n141 B.n140 585
R213 B.n139 B.n102 585
R214 B.n138 B.n137 585
R215 B.n136 B.n103 585
R216 B.n135 B.n134 585
R217 B.n133 B.n104 585
R218 B.n132 B.n131 585
R219 B.n130 B.n105 585
R220 B.n129 B.n128 585
R221 B.n127 B.n106 585
R222 B.n126 B.n125 585
R223 B.n124 B.n107 585
R224 B.n123 B.n122 585
R225 B.n121 B.n108 585
R226 B.n120 B.n119 585
R227 B.n118 B.n109 585
R228 B.n117 B.n116 585
R229 B.n115 B.n110 585
R230 B.n114 B.n113 585
R231 B.n112 B.n111 585
R232 B.n2 B.n0 585
R233 B.n413 B.n1 585
R234 B.n412 B.n411 585
R235 B.n410 B.n3 585
R236 B.n409 B.n408 585
R237 B.n407 B.n4 585
R238 B.n406 B.n405 585
R239 B.n404 B.n5 585
R240 B.n403 B.n402 585
R241 B.n401 B.n6 585
R242 B.n400 B.n399 585
R243 B.n398 B.n7 585
R244 B.n397 B.n396 585
R245 B.n395 B.n8 585
R246 B.n394 B.n393 585
R247 B.n392 B.n9 585
R248 B.n391 B.n390 585
R249 B.n389 B.n10 585
R250 B.n388 B.n387 585
R251 B.n386 B.n11 585
R252 B.n385 B.n384 585
R253 B.n383 B.n12 585
R254 B.n382 B.n381 585
R255 B.n380 B.n13 585
R256 B.n379 B.n378 585
R257 B.n377 B.n14 585
R258 B.n376 B.n375 585
R259 B.n374 B.n15 585
R260 B.n373 B.n372 585
R261 B.n371 B.n16 585
R262 B.n370 B.n369 585
R263 B.n368 B.n17 585
R264 B.n367 B.n366 585
R265 B.n365 B.n18 585
R266 B.n364 B.n363 585
R267 B.n362 B.n19 585
R268 B.n415 B.n414 585
R269 B.n161 B.n94 497.305
R270 B.n360 B.n19 497.305
R271 B.n209 B.n208 497.305
R272 B.n316 B.n315 497.305
R273 B.n81 B.t5 425.974
R274 B.n87 B.t8 425.974
R275 B.n26 B.t1 425.974
R276 B.n33 B.t10 425.974
R277 B.n82 B.t4 366.63
R278 B.n88 B.t7 366.63
R279 B.n27 B.t2 366.63
R280 B.n34 B.t11 366.63
R281 B.n81 B.t3 208.933
R282 B.n87 B.t6 208.933
R283 B.n26 B.t0 208.933
R284 B.n33 B.t9 208.933
R285 B.n161 B.n160 163.367
R286 B.n160 B.n159 163.367
R287 B.n159 B.n96 163.367
R288 B.n155 B.n96 163.367
R289 B.n155 B.n154 163.367
R290 B.n154 B.n153 163.367
R291 B.n153 B.n98 163.367
R292 B.n149 B.n98 163.367
R293 B.n149 B.n148 163.367
R294 B.n148 B.n147 163.367
R295 B.n147 B.n100 163.367
R296 B.n143 B.n100 163.367
R297 B.n143 B.n142 163.367
R298 B.n142 B.n141 163.367
R299 B.n141 B.n102 163.367
R300 B.n137 B.n102 163.367
R301 B.n137 B.n136 163.367
R302 B.n136 B.n135 163.367
R303 B.n135 B.n104 163.367
R304 B.n131 B.n104 163.367
R305 B.n131 B.n130 163.367
R306 B.n130 B.n129 163.367
R307 B.n129 B.n106 163.367
R308 B.n125 B.n106 163.367
R309 B.n125 B.n124 163.367
R310 B.n124 B.n123 163.367
R311 B.n123 B.n108 163.367
R312 B.n119 B.n108 163.367
R313 B.n119 B.n118 163.367
R314 B.n118 B.n117 163.367
R315 B.n117 B.n110 163.367
R316 B.n113 B.n110 163.367
R317 B.n113 B.n112 163.367
R318 B.n112 B.n2 163.367
R319 B.n414 B.n2 163.367
R320 B.n414 B.n413 163.367
R321 B.n413 B.n412 163.367
R322 B.n412 B.n3 163.367
R323 B.n408 B.n3 163.367
R324 B.n408 B.n407 163.367
R325 B.n407 B.n406 163.367
R326 B.n406 B.n5 163.367
R327 B.n402 B.n5 163.367
R328 B.n402 B.n401 163.367
R329 B.n401 B.n400 163.367
R330 B.n400 B.n7 163.367
R331 B.n396 B.n7 163.367
R332 B.n396 B.n395 163.367
R333 B.n395 B.n394 163.367
R334 B.n394 B.n9 163.367
R335 B.n390 B.n9 163.367
R336 B.n390 B.n389 163.367
R337 B.n389 B.n388 163.367
R338 B.n388 B.n11 163.367
R339 B.n384 B.n11 163.367
R340 B.n384 B.n383 163.367
R341 B.n383 B.n382 163.367
R342 B.n382 B.n13 163.367
R343 B.n378 B.n13 163.367
R344 B.n378 B.n377 163.367
R345 B.n377 B.n376 163.367
R346 B.n376 B.n15 163.367
R347 B.n372 B.n15 163.367
R348 B.n372 B.n371 163.367
R349 B.n371 B.n370 163.367
R350 B.n370 B.n17 163.367
R351 B.n366 B.n17 163.367
R352 B.n366 B.n365 163.367
R353 B.n365 B.n364 163.367
R354 B.n364 B.n19 163.367
R355 B.n165 B.n94 163.367
R356 B.n166 B.n165 163.367
R357 B.n167 B.n166 163.367
R358 B.n167 B.n92 163.367
R359 B.n171 B.n92 163.367
R360 B.n172 B.n171 163.367
R361 B.n173 B.n172 163.367
R362 B.n173 B.n90 163.367
R363 B.n177 B.n90 163.367
R364 B.n178 B.n177 163.367
R365 B.n178 B.n86 163.367
R366 B.n182 B.n86 163.367
R367 B.n183 B.n182 163.367
R368 B.n184 B.n183 163.367
R369 B.n184 B.n84 163.367
R370 B.n188 B.n84 163.367
R371 B.n189 B.n188 163.367
R372 B.n190 B.n189 163.367
R373 B.n190 B.n80 163.367
R374 B.n195 B.n80 163.367
R375 B.n196 B.n195 163.367
R376 B.n197 B.n196 163.367
R377 B.n197 B.n78 163.367
R378 B.n201 B.n78 163.367
R379 B.n202 B.n201 163.367
R380 B.n203 B.n202 163.367
R381 B.n203 B.n76 163.367
R382 B.n207 B.n76 163.367
R383 B.n208 B.n207 163.367
R384 B.n209 B.n74 163.367
R385 B.n213 B.n74 163.367
R386 B.n214 B.n213 163.367
R387 B.n215 B.n214 163.367
R388 B.n215 B.n72 163.367
R389 B.n219 B.n72 163.367
R390 B.n220 B.n219 163.367
R391 B.n221 B.n220 163.367
R392 B.n221 B.n70 163.367
R393 B.n225 B.n70 163.367
R394 B.n226 B.n225 163.367
R395 B.n227 B.n226 163.367
R396 B.n227 B.n68 163.367
R397 B.n231 B.n68 163.367
R398 B.n232 B.n231 163.367
R399 B.n233 B.n232 163.367
R400 B.n233 B.n66 163.367
R401 B.n237 B.n66 163.367
R402 B.n238 B.n237 163.367
R403 B.n239 B.n238 163.367
R404 B.n239 B.n64 163.367
R405 B.n243 B.n64 163.367
R406 B.n244 B.n243 163.367
R407 B.n245 B.n244 163.367
R408 B.n245 B.n62 163.367
R409 B.n249 B.n62 163.367
R410 B.n250 B.n249 163.367
R411 B.n251 B.n250 163.367
R412 B.n251 B.n60 163.367
R413 B.n255 B.n60 163.367
R414 B.n256 B.n255 163.367
R415 B.n257 B.n256 163.367
R416 B.n257 B.n58 163.367
R417 B.n261 B.n58 163.367
R418 B.n262 B.n261 163.367
R419 B.n263 B.n262 163.367
R420 B.n263 B.n56 163.367
R421 B.n267 B.n56 163.367
R422 B.n268 B.n267 163.367
R423 B.n269 B.n268 163.367
R424 B.n269 B.n54 163.367
R425 B.n273 B.n54 163.367
R426 B.n274 B.n273 163.367
R427 B.n275 B.n274 163.367
R428 B.n275 B.n52 163.367
R429 B.n279 B.n52 163.367
R430 B.n280 B.n279 163.367
R431 B.n281 B.n280 163.367
R432 B.n281 B.n50 163.367
R433 B.n285 B.n50 163.367
R434 B.n286 B.n285 163.367
R435 B.n287 B.n286 163.367
R436 B.n287 B.n48 163.367
R437 B.n291 B.n48 163.367
R438 B.n292 B.n291 163.367
R439 B.n293 B.n292 163.367
R440 B.n293 B.n46 163.367
R441 B.n297 B.n46 163.367
R442 B.n298 B.n297 163.367
R443 B.n299 B.n298 163.367
R444 B.n299 B.n44 163.367
R445 B.n303 B.n44 163.367
R446 B.n304 B.n303 163.367
R447 B.n305 B.n304 163.367
R448 B.n305 B.n42 163.367
R449 B.n309 B.n42 163.367
R450 B.n310 B.n309 163.367
R451 B.n311 B.n310 163.367
R452 B.n311 B.n40 163.367
R453 B.n315 B.n40 163.367
R454 B.n360 B.n359 163.367
R455 B.n359 B.n358 163.367
R456 B.n358 B.n21 163.367
R457 B.n354 B.n21 163.367
R458 B.n354 B.n353 163.367
R459 B.n353 B.n352 163.367
R460 B.n352 B.n23 163.367
R461 B.n348 B.n23 163.367
R462 B.n348 B.n347 163.367
R463 B.n347 B.n346 163.367
R464 B.n346 B.n25 163.367
R465 B.n342 B.n25 163.367
R466 B.n342 B.n341 163.367
R467 B.n341 B.n340 163.367
R468 B.n340 B.n30 163.367
R469 B.n336 B.n30 163.367
R470 B.n336 B.n335 163.367
R471 B.n335 B.n334 163.367
R472 B.n334 B.n32 163.367
R473 B.n329 B.n32 163.367
R474 B.n329 B.n328 163.367
R475 B.n328 B.n327 163.367
R476 B.n327 B.n36 163.367
R477 B.n323 B.n36 163.367
R478 B.n323 B.n322 163.367
R479 B.n322 B.n321 163.367
R480 B.n321 B.n38 163.367
R481 B.n317 B.n38 163.367
R482 B.n317 B.n316 163.367
R483 B.n193 B.n82 59.5399
R484 B.n89 B.n88 59.5399
R485 B.n28 B.n27 59.5399
R486 B.n331 B.n34 59.5399
R487 B.n82 B.n81 59.346
R488 B.n88 B.n87 59.346
R489 B.n27 B.n26 59.346
R490 B.n34 B.n33 59.346
R491 B.n362 B.n361 32.3127
R492 B.n314 B.n39 32.3127
R493 B.n210 B.n75 32.3127
R494 B.n163 B.n162 32.3127
R495 B B.n415 18.0485
R496 B.n361 B.n20 10.6151
R497 B.n357 B.n20 10.6151
R498 B.n357 B.n356 10.6151
R499 B.n356 B.n355 10.6151
R500 B.n355 B.n22 10.6151
R501 B.n351 B.n22 10.6151
R502 B.n351 B.n350 10.6151
R503 B.n350 B.n349 10.6151
R504 B.n349 B.n24 10.6151
R505 B.n345 B.n344 10.6151
R506 B.n344 B.n343 10.6151
R507 B.n343 B.n29 10.6151
R508 B.n339 B.n29 10.6151
R509 B.n339 B.n338 10.6151
R510 B.n338 B.n337 10.6151
R511 B.n337 B.n31 10.6151
R512 B.n333 B.n31 10.6151
R513 B.n333 B.n332 10.6151
R514 B.n330 B.n35 10.6151
R515 B.n326 B.n35 10.6151
R516 B.n326 B.n325 10.6151
R517 B.n325 B.n324 10.6151
R518 B.n324 B.n37 10.6151
R519 B.n320 B.n37 10.6151
R520 B.n320 B.n319 10.6151
R521 B.n319 B.n318 10.6151
R522 B.n318 B.n39 10.6151
R523 B.n211 B.n210 10.6151
R524 B.n212 B.n211 10.6151
R525 B.n212 B.n73 10.6151
R526 B.n216 B.n73 10.6151
R527 B.n217 B.n216 10.6151
R528 B.n218 B.n217 10.6151
R529 B.n218 B.n71 10.6151
R530 B.n222 B.n71 10.6151
R531 B.n223 B.n222 10.6151
R532 B.n224 B.n223 10.6151
R533 B.n224 B.n69 10.6151
R534 B.n228 B.n69 10.6151
R535 B.n229 B.n228 10.6151
R536 B.n230 B.n229 10.6151
R537 B.n230 B.n67 10.6151
R538 B.n234 B.n67 10.6151
R539 B.n235 B.n234 10.6151
R540 B.n236 B.n235 10.6151
R541 B.n236 B.n65 10.6151
R542 B.n240 B.n65 10.6151
R543 B.n241 B.n240 10.6151
R544 B.n242 B.n241 10.6151
R545 B.n242 B.n63 10.6151
R546 B.n246 B.n63 10.6151
R547 B.n247 B.n246 10.6151
R548 B.n248 B.n247 10.6151
R549 B.n248 B.n61 10.6151
R550 B.n252 B.n61 10.6151
R551 B.n253 B.n252 10.6151
R552 B.n254 B.n253 10.6151
R553 B.n254 B.n59 10.6151
R554 B.n258 B.n59 10.6151
R555 B.n259 B.n258 10.6151
R556 B.n260 B.n259 10.6151
R557 B.n260 B.n57 10.6151
R558 B.n264 B.n57 10.6151
R559 B.n265 B.n264 10.6151
R560 B.n266 B.n265 10.6151
R561 B.n266 B.n55 10.6151
R562 B.n270 B.n55 10.6151
R563 B.n271 B.n270 10.6151
R564 B.n272 B.n271 10.6151
R565 B.n272 B.n53 10.6151
R566 B.n276 B.n53 10.6151
R567 B.n277 B.n276 10.6151
R568 B.n278 B.n277 10.6151
R569 B.n278 B.n51 10.6151
R570 B.n282 B.n51 10.6151
R571 B.n283 B.n282 10.6151
R572 B.n284 B.n283 10.6151
R573 B.n284 B.n49 10.6151
R574 B.n288 B.n49 10.6151
R575 B.n289 B.n288 10.6151
R576 B.n290 B.n289 10.6151
R577 B.n290 B.n47 10.6151
R578 B.n294 B.n47 10.6151
R579 B.n295 B.n294 10.6151
R580 B.n296 B.n295 10.6151
R581 B.n296 B.n45 10.6151
R582 B.n300 B.n45 10.6151
R583 B.n301 B.n300 10.6151
R584 B.n302 B.n301 10.6151
R585 B.n302 B.n43 10.6151
R586 B.n306 B.n43 10.6151
R587 B.n307 B.n306 10.6151
R588 B.n308 B.n307 10.6151
R589 B.n308 B.n41 10.6151
R590 B.n312 B.n41 10.6151
R591 B.n313 B.n312 10.6151
R592 B.n314 B.n313 10.6151
R593 B.n164 B.n163 10.6151
R594 B.n164 B.n93 10.6151
R595 B.n168 B.n93 10.6151
R596 B.n169 B.n168 10.6151
R597 B.n170 B.n169 10.6151
R598 B.n170 B.n91 10.6151
R599 B.n174 B.n91 10.6151
R600 B.n175 B.n174 10.6151
R601 B.n176 B.n175 10.6151
R602 B.n180 B.n179 10.6151
R603 B.n181 B.n180 10.6151
R604 B.n181 B.n85 10.6151
R605 B.n185 B.n85 10.6151
R606 B.n186 B.n185 10.6151
R607 B.n187 B.n186 10.6151
R608 B.n187 B.n83 10.6151
R609 B.n191 B.n83 10.6151
R610 B.n192 B.n191 10.6151
R611 B.n194 B.n79 10.6151
R612 B.n198 B.n79 10.6151
R613 B.n199 B.n198 10.6151
R614 B.n200 B.n199 10.6151
R615 B.n200 B.n77 10.6151
R616 B.n204 B.n77 10.6151
R617 B.n205 B.n204 10.6151
R618 B.n206 B.n205 10.6151
R619 B.n206 B.n75 10.6151
R620 B.n162 B.n95 10.6151
R621 B.n158 B.n95 10.6151
R622 B.n158 B.n157 10.6151
R623 B.n157 B.n156 10.6151
R624 B.n156 B.n97 10.6151
R625 B.n152 B.n97 10.6151
R626 B.n152 B.n151 10.6151
R627 B.n151 B.n150 10.6151
R628 B.n150 B.n99 10.6151
R629 B.n146 B.n99 10.6151
R630 B.n146 B.n145 10.6151
R631 B.n145 B.n144 10.6151
R632 B.n144 B.n101 10.6151
R633 B.n140 B.n101 10.6151
R634 B.n140 B.n139 10.6151
R635 B.n139 B.n138 10.6151
R636 B.n138 B.n103 10.6151
R637 B.n134 B.n103 10.6151
R638 B.n134 B.n133 10.6151
R639 B.n133 B.n132 10.6151
R640 B.n132 B.n105 10.6151
R641 B.n128 B.n105 10.6151
R642 B.n128 B.n127 10.6151
R643 B.n127 B.n126 10.6151
R644 B.n126 B.n107 10.6151
R645 B.n122 B.n107 10.6151
R646 B.n122 B.n121 10.6151
R647 B.n121 B.n120 10.6151
R648 B.n120 B.n109 10.6151
R649 B.n116 B.n109 10.6151
R650 B.n116 B.n115 10.6151
R651 B.n115 B.n114 10.6151
R652 B.n114 B.n111 10.6151
R653 B.n111 B.n0 10.6151
R654 B.n411 B.n1 10.6151
R655 B.n411 B.n410 10.6151
R656 B.n410 B.n409 10.6151
R657 B.n409 B.n4 10.6151
R658 B.n405 B.n4 10.6151
R659 B.n405 B.n404 10.6151
R660 B.n404 B.n403 10.6151
R661 B.n403 B.n6 10.6151
R662 B.n399 B.n6 10.6151
R663 B.n399 B.n398 10.6151
R664 B.n398 B.n397 10.6151
R665 B.n397 B.n8 10.6151
R666 B.n393 B.n8 10.6151
R667 B.n393 B.n392 10.6151
R668 B.n392 B.n391 10.6151
R669 B.n391 B.n10 10.6151
R670 B.n387 B.n10 10.6151
R671 B.n387 B.n386 10.6151
R672 B.n386 B.n385 10.6151
R673 B.n385 B.n12 10.6151
R674 B.n381 B.n12 10.6151
R675 B.n381 B.n380 10.6151
R676 B.n380 B.n379 10.6151
R677 B.n379 B.n14 10.6151
R678 B.n375 B.n14 10.6151
R679 B.n375 B.n374 10.6151
R680 B.n374 B.n373 10.6151
R681 B.n373 B.n16 10.6151
R682 B.n369 B.n16 10.6151
R683 B.n369 B.n368 10.6151
R684 B.n368 B.n367 10.6151
R685 B.n367 B.n18 10.6151
R686 B.n363 B.n18 10.6151
R687 B.n363 B.n362 10.6151
R688 B.n28 B.n24 9.36635
R689 B.n331 B.n330 9.36635
R690 B.n176 B.n89 9.36635
R691 B.n194 B.n193 9.36635
R692 B.n415 B.n0 2.81026
R693 B.n415 B.n1 2.81026
R694 B.n345 B.n28 1.24928
R695 B.n332 B.n331 1.24928
R696 B.n179 B.n89 1.24928
R697 B.n193 B.n192 1.24928
C0 VDD1 w_n2806_n1224# 1.18034f
C1 VTAIL VN 1.48361f
C2 VTAIL VP 1.49771f
C3 VDD1 VDD2 1.05217f
C4 B VTAIL 1.31221f
C5 VDD2 w_n2806_n1224# 1.23838f
C6 VDD1 VN 0.155899f
C7 VN w_n2806_n1224# 4.56028f
C8 VDD1 VP 1.06156f
C9 B VDD1 0.994334f
C10 VP w_n2806_n1224# 4.9145f
C11 B w_n2806_n1224# 6.45648f
C12 VDD2 VN 0.809042f
C13 VDD2 VP 0.410611f
C14 B VDD2 1.04918f
C15 VP VN 4.30616f
C16 B VN 0.963149f
C17 B VP 1.56182f
C18 VDD1 VTAIL 2.92685f
C19 VTAIL w_n2806_n1224# 1.50963f
C20 VDD2 VTAIL 2.98192f
C21 VDD2 VSUBS 0.682099f
C22 VDD1 VSUBS 3.460555f
C23 VTAIL VSUBS 0.406266f
C24 VN VSUBS 5.4497f
C25 VP VSUBS 1.779926f
C26 B VSUBS 3.286642f
C27 w_n2806_n1224# VSUBS 44.144f
C28 B.n0 VSUBS 0.006493f
C29 B.n1 VSUBS 0.006493f
C30 B.n2 VSUBS 0.010268f
C31 B.n3 VSUBS 0.010268f
C32 B.n4 VSUBS 0.010268f
C33 B.n5 VSUBS 0.010268f
C34 B.n6 VSUBS 0.010268f
C35 B.n7 VSUBS 0.010268f
C36 B.n8 VSUBS 0.010268f
C37 B.n9 VSUBS 0.010268f
C38 B.n10 VSUBS 0.010268f
C39 B.n11 VSUBS 0.010268f
C40 B.n12 VSUBS 0.010268f
C41 B.n13 VSUBS 0.010268f
C42 B.n14 VSUBS 0.010268f
C43 B.n15 VSUBS 0.010268f
C44 B.n16 VSUBS 0.010268f
C45 B.n17 VSUBS 0.010268f
C46 B.n18 VSUBS 0.010268f
C47 B.n19 VSUBS 0.023034f
C48 B.n20 VSUBS 0.010268f
C49 B.n21 VSUBS 0.010268f
C50 B.n22 VSUBS 0.010268f
C51 B.n23 VSUBS 0.010268f
C52 B.n24 VSUBS 0.009664f
C53 B.n25 VSUBS 0.010268f
C54 B.t2 VSUBS 0.035478f
C55 B.t1 VSUBS 0.043988f
C56 B.t0 VSUBS 0.259189f
C57 B.n26 VSUBS 0.095976f
C58 B.n27 VSUBS 0.075729f
C59 B.n28 VSUBS 0.023789f
C60 B.n29 VSUBS 0.010268f
C61 B.n30 VSUBS 0.010268f
C62 B.n31 VSUBS 0.010268f
C63 B.n32 VSUBS 0.010268f
C64 B.t11 VSUBS 0.035478f
C65 B.t10 VSUBS 0.043988f
C66 B.t9 VSUBS 0.259189f
C67 B.n33 VSUBS 0.095976f
C68 B.n34 VSUBS 0.075729f
C69 B.n35 VSUBS 0.010268f
C70 B.n36 VSUBS 0.010268f
C71 B.n37 VSUBS 0.010268f
C72 B.n38 VSUBS 0.010268f
C73 B.n39 VSUBS 0.023453f
C74 B.n40 VSUBS 0.010268f
C75 B.n41 VSUBS 0.010268f
C76 B.n42 VSUBS 0.010268f
C77 B.n43 VSUBS 0.010268f
C78 B.n44 VSUBS 0.010268f
C79 B.n45 VSUBS 0.010268f
C80 B.n46 VSUBS 0.010268f
C81 B.n47 VSUBS 0.010268f
C82 B.n48 VSUBS 0.010268f
C83 B.n49 VSUBS 0.010268f
C84 B.n50 VSUBS 0.010268f
C85 B.n51 VSUBS 0.010268f
C86 B.n52 VSUBS 0.010268f
C87 B.n53 VSUBS 0.010268f
C88 B.n54 VSUBS 0.010268f
C89 B.n55 VSUBS 0.010268f
C90 B.n56 VSUBS 0.010268f
C91 B.n57 VSUBS 0.010268f
C92 B.n58 VSUBS 0.010268f
C93 B.n59 VSUBS 0.010268f
C94 B.n60 VSUBS 0.010268f
C95 B.n61 VSUBS 0.010268f
C96 B.n62 VSUBS 0.010268f
C97 B.n63 VSUBS 0.010268f
C98 B.n64 VSUBS 0.010268f
C99 B.n65 VSUBS 0.010268f
C100 B.n66 VSUBS 0.010268f
C101 B.n67 VSUBS 0.010268f
C102 B.n68 VSUBS 0.010268f
C103 B.n69 VSUBS 0.010268f
C104 B.n70 VSUBS 0.010268f
C105 B.n71 VSUBS 0.010268f
C106 B.n72 VSUBS 0.010268f
C107 B.n73 VSUBS 0.010268f
C108 B.n74 VSUBS 0.010268f
C109 B.n75 VSUBS 0.024679f
C110 B.n76 VSUBS 0.010268f
C111 B.n77 VSUBS 0.010268f
C112 B.n78 VSUBS 0.010268f
C113 B.n79 VSUBS 0.010268f
C114 B.n80 VSUBS 0.010268f
C115 B.t4 VSUBS 0.035478f
C116 B.t5 VSUBS 0.043988f
C117 B.t3 VSUBS 0.259189f
C118 B.n81 VSUBS 0.095976f
C119 B.n82 VSUBS 0.075729f
C120 B.n83 VSUBS 0.010268f
C121 B.n84 VSUBS 0.010268f
C122 B.n85 VSUBS 0.010268f
C123 B.n86 VSUBS 0.010268f
C124 B.t7 VSUBS 0.035478f
C125 B.t8 VSUBS 0.043988f
C126 B.t6 VSUBS 0.259189f
C127 B.n87 VSUBS 0.095976f
C128 B.n88 VSUBS 0.075729f
C129 B.n89 VSUBS 0.023789f
C130 B.n90 VSUBS 0.010268f
C131 B.n91 VSUBS 0.010268f
C132 B.n92 VSUBS 0.010268f
C133 B.n93 VSUBS 0.010268f
C134 B.n94 VSUBS 0.024679f
C135 B.n95 VSUBS 0.010268f
C136 B.n96 VSUBS 0.010268f
C137 B.n97 VSUBS 0.010268f
C138 B.n98 VSUBS 0.010268f
C139 B.n99 VSUBS 0.010268f
C140 B.n100 VSUBS 0.010268f
C141 B.n101 VSUBS 0.010268f
C142 B.n102 VSUBS 0.010268f
C143 B.n103 VSUBS 0.010268f
C144 B.n104 VSUBS 0.010268f
C145 B.n105 VSUBS 0.010268f
C146 B.n106 VSUBS 0.010268f
C147 B.n107 VSUBS 0.010268f
C148 B.n108 VSUBS 0.010268f
C149 B.n109 VSUBS 0.010268f
C150 B.n110 VSUBS 0.010268f
C151 B.n111 VSUBS 0.010268f
C152 B.n112 VSUBS 0.010268f
C153 B.n113 VSUBS 0.010268f
C154 B.n114 VSUBS 0.010268f
C155 B.n115 VSUBS 0.010268f
C156 B.n116 VSUBS 0.010268f
C157 B.n117 VSUBS 0.010268f
C158 B.n118 VSUBS 0.010268f
C159 B.n119 VSUBS 0.010268f
C160 B.n120 VSUBS 0.010268f
C161 B.n121 VSUBS 0.010268f
C162 B.n122 VSUBS 0.010268f
C163 B.n123 VSUBS 0.010268f
C164 B.n124 VSUBS 0.010268f
C165 B.n125 VSUBS 0.010268f
C166 B.n126 VSUBS 0.010268f
C167 B.n127 VSUBS 0.010268f
C168 B.n128 VSUBS 0.010268f
C169 B.n129 VSUBS 0.010268f
C170 B.n130 VSUBS 0.010268f
C171 B.n131 VSUBS 0.010268f
C172 B.n132 VSUBS 0.010268f
C173 B.n133 VSUBS 0.010268f
C174 B.n134 VSUBS 0.010268f
C175 B.n135 VSUBS 0.010268f
C176 B.n136 VSUBS 0.010268f
C177 B.n137 VSUBS 0.010268f
C178 B.n138 VSUBS 0.010268f
C179 B.n139 VSUBS 0.010268f
C180 B.n140 VSUBS 0.010268f
C181 B.n141 VSUBS 0.010268f
C182 B.n142 VSUBS 0.010268f
C183 B.n143 VSUBS 0.010268f
C184 B.n144 VSUBS 0.010268f
C185 B.n145 VSUBS 0.010268f
C186 B.n146 VSUBS 0.010268f
C187 B.n147 VSUBS 0.010268f
C188 B.n148 VSUBS 0.010268f
C189 B.n149 VSUBS 0.010268f
C190 B.n150 VSUBS 0.010268f
C191 B.n151 VSUBS 0.010268f
C192 B.n152 VSUBS 0.010268f
C193 B.n153 VSUBS 0.010268f
C194 B.n154 VSUBS 0.010268f
C195 B.n155 VSUBS 0.010268f
C196 B.n156 VSUBS 0.010268f
C197 B.n157 VSUBS 0.010268f
C198 B.n158 VSUBS 0.010268f
C199 B.n159 VSUBS 0.010268f
C200 B.n160 VSUBS 0.010268f
C201 B.n161 VSUBS 0.023034f
C202 B.n162 VSUBS 0.023034f
C203 B.n163 VSUBS 0.024679f
C204 B.n164 VSUBS 0.010268f
C205 B.n165 VSUBS 0.010268f
C206 B.n166 VSUBS 0.010268f
C207 B.n167 VSUBS 0.010268f
C208 B.n168 VSUBS 0.010268f
C209 B.n169 VSUBS 0.010268f
C210 B.n170 VSUBS 0.010268f
C211 B.n171 VSUBS 0.010268f
C212 B.n172 VSUBS 0.010268f
C213 B.n173 VSUBS 0.010268f
C214 B.n174 VSUBS 0.010268f
C215 B.n175 VSUBS 0.010268f
C216 B.n176 VSUBS 0.009664f
C217 B.n177 VSUBS 0.010268f
C218 B.n178 VSUBS 0.010268f
C219 B.n179 VSUBS 0.005738f
C220 B.n180 VSUBS 0.010268f
C221 B.n181 VSUBS 0.010268f
C222 B.n182 VSUBS 0.010268f
C223 B.n183 VSUBS 0.010268f
C224 B.n184 VSUBS 0.010268f
C225 B.n185 VSUBS 0.010268f
C226 B.n186 VSUBS 0.010268f
C227 B.n187 VSUBS 0.010268f
C228 B.n188 VSUBS 0.010268f
C229 B.n189 VSUBS 0.010268f
C230 B.n190 VSUBS 0.010268f
C231 B.n191 VSUBS 0.010268f
C232 B.n192 VSUBS 0.005738f
C233 B.n193 VSUBS 0.023789f
C234 B.n194 VSUBS 0.009664f
C235 B.n195 VSUBS 0.010268f
C236 B.n196 VSUBS 0.010268f
C237 B.n197 VSUBS 0.010268f
C238 B.n198 VSUBS 0.010268f
C239 B.n199 VSUBS 0.010268f
C240 B.n200 VSUBS 0.010268f
C241 B.n201 VSUBS 0.010268f
C242 B.n202 VSUBS 0.010268f
C243 B.n203 VSUBS 0.010268f
C244 B.n204 VSUBS 0.010268f
C245 B.n205 VSUBS 0.010268f
C246 B.n206 VSUBS 0.010268f
C247 B.n207 VSUBS 0.010268f
C248 B.n208 VSUBS 0.024679f
C249 B.n209 VSUBS 0.023034f
C250 B.n210 VSUBS 0.023034f
C251 B.n211 VSUBS 0.010268f
C252 B.n212 VSUBS 0.010268f
C253 B.n213 VSUBS 0.010268f
C254 B.n214 VSUBS 0.010268f
C255 B.n215 VSUBS 0.010268f
C256 B.n216 VSUBS 0.010268f
C257 B.n217 VSUBS 0.010268f
C258 B.n218 VSUBS 0.010268f
C259 B.n219 VSUBS 0.010268f
C260 B.n220 VSUBS 0.010268f
C261 B.n221 VSUBS 0.010268f
C262 B.n222 VSUBS 0.010268f
C263 B.n223 VSUBS 0.010268f
C264 B.n224 VSUBS 0.010268f
C265 B.n225 VSUBS 0.010268f
C266 B.n226 VSUBS 0.010268f
C267 B.n227 VSUBS 0.010268f
C268 B.n228 VSUBS 0.010268f
C269 B.n229 VSUBS 0.010268f
C270 B.n230 VSUBS 0.010268f
C271 B.n231 VSUBS 0.010268f
C272 B.n232 VSUBS 0.010268f
C273 B.n233 VSUBS 0.010268f
C274 B.n234 VSUBS 0.010268f
C275 B.n235 VSUBS 0.010268f
C276 B.n236 VSUBS 0.010268f
C277 B.n237 VSUBS 0.010268f
C278 B.n238 VSUBS 0.010268f
C279 B.n239 VSUBS 0.010268f
C280 B.n240 VSUBS 0.010268f
C281 B.n241 VSUBS 0.010268f
C282 B.n242 VSUBS 0.010268f
C283 B.n243 VSUBS 0.010268f
C284 B.n244 VSUBS 0.010268f
C285 B.n245 VSUBS 0.010268f
C286 B.n246 VSUBS 0.010268f
C287 B.n247 VSUBS 0.010268f
C288 B.n248 VSUBS 0.010268f
C289 B.n249 VSUBS 0.010268f
C290 B.n250 VSUBS 0.010268f
C291 B.n251 VSUBS 0.010268f
C292 B.n252 VSUBS 0.010268f
C293 B.n253 VSUBS 0.010268f
C294 B.n254 VSUBS 0.010268f
C295 B.n255 VSUBS 0.010268f
C296 B.n256 VSUBS 0.010268f
C297 B.n257 VSUBS 0.010268f
C298 B.n258 VSUBS 0.010268f
C299 B.n259 VSUBS 0.010268f
C300 B.n260 VSUBS 0.010268f
C301 B.n261 VSUBS 0.010268f
C302 B.n262 VSUBS 0.010268f
C303 B.n263 VSUBS 0.010268f
C304 B.n264 VSUBS 0.010268f
C305 B.n265 VSUBS 0.010268f
C306 B.n266 VSUBS 0.010268f
C307 B.n267 VSUBS 0.010268f
C308 B.n268 VSUBS 0.010268f
C309 B.n269 VSUBS 0.010268f
C310 B.n270 VSUBS 0.010268f
C311 B.n271 VSUBS 0.010268f
C312 B.n272 VSUBS 0.010268f
C313 B.n273 VSUBS 0.010268f
C314 B.n274 VSUBS 0.010268f
C315 B.n275 VSUBS 0.010268f
C316 B.n276 VSUBS 0.010268f
C317 B.n277 VSUBS 0.010268f
C318 B.n278 VSUBS 0.010268f
C319 B.n279 VSUBS 0.010268f
C320 B.n280 VSUBS 0.010268f
C321 B.n281 VSUBS 0.010268f
C322 B.n282 VSUBS 0.010268f
C323 B.n283 VSUBS 0.010268f
C324 B.n284 VSUBS 0.010268f
C325 B.n285 VSUBS 0.010268f
C326 B.n286 VSUBS 0.010268f
C327 B.n287 VSUBS 0.010268f
C328 B.n288 VSUBS 0.010268f
C329 B.n289 VSUBS 0.010268f
C330 B.n290 VSUBS 0.010268f
C331 B.n291 VSUBS 0.010268f
C332 B.n292 VSUBS 0.010268f
C333 B.n293 VSUBS 0.010268f
C334 B.n294 VSUBS 0.010268f
C335 B.n295 VSUBS 0.010268f
C336 B.n296 VSUBS 0.010268f
C337 B.n297 VSUBS 0.010268f
C338 B.n298 VSUBS 0.010268f
C339 B.n299 VSUBS 0.010268f
C340 B.n300 VSUBS 0.010268f
C341 B.n301 VSUBS 0.010268f
C342 B.n302 VSUBS 0.010268f
C343 B.n303 VSUBS 0.010268f
C344 B.n304 VSUBS 0.010268f
C345 B.n305 VSUBS 0.010268f
C346 B.n306 VSUBS 0.010268f
C347 B.n307 VSUBS 0.010268f
C348 B.n308 VSUBS 0.010268f
C349 B.n309 VSUBS 0.010268f
C350 B.n310 VSUBS 0.010268f
C351 B.n311 VSUBS 0.010268f
C352 B.n312 VSUBS 0.010268f
C353 B.n313 VSUBS 0.010268f
C354 B.n314 VSUBS 0.024261f
C355 B.n315 VSUBS 0.023034f
C356 B.n316 VSUBS 0.024679f
C357 B.n317 VSUBS 0.010268f
C358 B.n318 VSUBS 0.010268f
C359 B.n319 VSUBS 0.010268f
C360 B.n320 VSUBS 0.010268f
C361 B.n321 VSUBS 0.010268f
C362 B.n322 VSUBS 0.010268f
C363 B.n323 VSUBS 0.010268f
C364 B.n324 VSUBS 0.010268f
C365 B.n325 VSUBS 0.010268f
C366 B.n326 VSUBS 0.010268f
C367 B.n327 VSUBS 0.010268f
C368 B.n328 VSUBS 0.010268f
C369 B.n329 VSUBS 0.010268f
C370 B.n330 VSUBS 0.009664f
C371 B.n331 VSUBS 0.023789f
C372 B.n332 VSUBS 0.005738f
C373 B.n333 VSUBS 0.010268f
C374 B.n334 VSUBS 0.010268f
C375 B.n335 VSUBS 0.010268f
C376 B.n336 VSUBS 0.010268f
C377 B.n337 VSUBS 0.010268f
C378 B.n338 VSUBS 0.010268f
C379 B.n339 VSUBS 0.010268f
C380 B.n340 VSUBS 0.010268f
C381 B.n341 VSUBS 0.010268f
C382 B.n342 VSUBS 0.010268f
C383 B.n343 VSUBS 0.010268f
C384 B.n344 VSUBS 0.010268f
C385 B.n345 VSUBS 0.005738f
C386 B.n346 VSUBS 0.010268f
C387 B.n347 VSUBS 0.010268f
C388 B.n348 VSUBS 0.010268f
C389 B.n349 VSUBS 0.010268f
C390 B.n350 VSUBS 0.010268f
C391 B.n351 VSUBS 0.010268f
C392 B.n352 VSUBS 0.010268f
C393 B.n353 VSUBS 0.010268f
C394 B.n354 VSUBS 0.010268f
C395 B.n355 VSUBS 0.010268f
C396 B.n356 VSUBS 0.010268f
C397 B.n357 VSUBS 0.010268f
C398 B.n358 VSUBS 0.010268f
C399 B.n359 VSUBS 0.010268f
C400 B.n360 VSUBS 0.024679f
C401 B.n361 VSUBS 0.024679f
C402 B.n362 VSUBS 0.023034f
C403 B.n363 VSUBS 0.010268f
C404 B.n364 VSUBS 0.010268f
C405 B.n365 VSUBS 0.010268f
C406 B.n366 VSUBS 0.010268f
C407 B.n367 VSUBS 0.010268f
C408 B.n368 VSUBS 0.010268f
C409 B.n369 VSUBS 0.010268f
C410 B.n370 VSUBS 0.010268f
C411 B.n371 VSUBS 0.010268f
C412 B.n372 VSUBS 0.010268f
C413 B.n373 VSUBS 0.010268f
C414 B.n374 VSUBS 0.010268f
C415 B.n375 VSUBS 0.010268f
C416 B.n376 VSUBS 0.010268f
C417 B.n377 VSUBS 0.010268f
C418 B.n378 VSUBS 0.010268f
C419 B.n379 VSUBS 0.010268f
C420 B.n380 VSUBS 0.010268f
C421 B.n381 VSUBS 0.010268f
C422 B.n382 VSUBS 0.010268f
C423 B.n383 VSUBS 0.010268f
C424 B.n384 VSUBS 0.010268f
C425 B.n385 VSUBS 0.010268f
C426 B.n386 VSUBS 0.010268f
C427 B.n387 VSUBS 0.010268f
C428 B.n388 VSUBS 0.010268f
C429 B.n389 VSUBS 0.010268f
C430 B.n390 VSUBS 0.010268f
C431 B.n391 VSUBS 0.010268f
C432 B.n392 VSUBS 0.010268f
C433 B.n393 VSUBS 0.010268f
C434 B.n394 VSUBS 0.010268f
C435 B.n395 VSUBS 0.010268f
C436 B.n396 VSUBS 0.010268f
C437 B.n397 VSUBS 0.010268f
C438 B.n398 VSUBS 0.010268f
C439 B.n399 VSUBS 0.010268f
C440 B.n400 VSUBS 0.010268f
C441 B.n401 VSUBS 0.010268f
C442 B.n402 VSUBS 0.010268f
C443 B.n403 VSUBS 0.010268f
C444 B.n404 VSUBS 0.010268f
C445 B.n405 VSUBS 0.010268f
C446 B.n406 VSUBS 0.010268f
C447 B.n407 VSUBS 0.010268f
C448 B.n408 VSUBS 0.010268f
C449 B.n409 VSUBS 0.010268f
C450 B.n410 VSUBS 0.010268f
C451 B.n411 VSUBS 0.010268f
C452 B.n412 VSUBS 0.010268f
C453 B.n413 VSUBS 0.010268f
C454 B.n414 VSUBS 0.010268f
C455 B.n415 VSUBS 0.023249f
C456 VDD2.t3 VSUBS 0.023772f
C457 VDD2.t0 VSUBS 0.023772f
C458 VDD2.n0 VSUBS 0.153474f
C459 VDD2.t1 VSUBS 0.023772f
C460 VDD2.t2 VSUBS 0.023772f
C461 VDD2.n1 VSUBS 0.077748f
C462 VDD2.n2 VSUBS 2.46887f
C463 VN.t0 VSUBS 0.776794f
C464 VN.t3 VSUBS 0.765951f
C465 VN.n0 VSUBS 0.517099f
C466 VN.t1 VSUBS 0.776794f
C467 VN.t2 VSUBS 0.765951f
C468 VN.n1 VSUBS 2.68306f
C469 VDD1.t1 VSUBS 0.022333f
C470 VDD1.t3 VSUBS 0.022333f
C471 VDD1.n0 VSUBS 0.073109f
C472 VDD1.t2 VSUBS 0.022333f
C473 VDD1.t0 VSUBS 0.022333f
C474 VDD1.n1 VSUBS 0.149147f
C475 VTAIL.t3 VSUBS 0.104549f
C476 VTAIL.n0 VSUBS 0.299319f
C477 VTAIL.t4 VSUBS 0.104549f
C478 VTAIL.n1 VSUBS 0.383372f
C479 VTAIL.t6 VSUBS 0.104549f
C480 VTAIL.n2 VSUBS 0.88253f
C481 VTAIL.t1 VSUBS 0.104549f
C482 VTAIL.n3 VSUBS 0.88253f
C483 VTAIL.t2 VSUBS 0.104549f
C484 VTAIL.n4 VSUBS 0.383372f
C485 VTAIL.t5 VSUBS 0.104549f
C486 VTAIL.n5 VSUBS 0.383372f
C487 VTAIL.t7 VSUBS 0.104549f
C488 VTAIL.n6 VSUBS 0.88253f
C489 VTAIL.t0 VSUBS 0.104549f
C490 VTAIL.n7 VSUBS 0.790718f
C491 VP.n0 VSUBS 0.06907f
C492 VP.t3 VSUBS 0.379463f
C493 VP.n1 VSUBS 0.103581f
C494 VP.n2 VSUBS 0.052393f
C495 VP.n3 VSUBS 0.052071f
C496 VP.t0 VSUBS 0.798108f
C497 VP.t2 VSUBS 0.809406f
C498 VP.n4 VSUBS 2.76731f
C499 VP.t1 VSUBS 0.379463f
C500 VP.n5 VSUBS 0.378889f
C501 VP.n6 VSUBS 2.20361f
C502 VP.n7 VSUBS 0.06907f
C503 VP.n8 VSUBS 0.052393f
C504 VP.n9 VSUBS 0.097157f
C505 VP.n10 VSUBS 0.103581f
C506 VP.n11 VSUBS 0.042316f
C507 VP.n12 VSUBS 0.052393f
C508 VP.n13 VSUBS 0.052393f
C509 VP.n14 VSUBS 0.052393f
C510 VP.n15 VSUBS 0.097157f
C511 VP.n16 VSUBS 0.052071f
C512 VP.n17 VSUBS 0.378889f
C513 VP.n18 VSUBS 0.097635f
.ends

