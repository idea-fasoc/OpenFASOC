* NGSPICE file created from diff_pair_sample_1719.ext - technology: sky130A

.subckt diff_pair_sample_1719 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=1.69455 ps=10.6 w=10.27 l=2.08
X1 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=1.69455 ps=10.6 w=10.27 l=2.08
X2 VDD2.t3 VN.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.69455 pd=10.6 as=4.0053 ps=21.32 w=10.27 l=2.08
X3 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=0 ps=0 w=10.27 l=2.08
X4 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.69455 pd=10.6 as=4.0053 ps=21.32 w=10.27 l=2.08
X5 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=1.69455 ps=10.6 w=10.27 l=2.08
X6 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=0 ps=0 w=10.27 l=2.08
X7 VDD2.t1 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.69455 pd=10.6 as=4.0053 ps=21.32 w=10.27 l=2.08
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=0 ps=0 w=10.27 l=2.08
X9 VTAIL.t4 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=1.69455 ps=10.6 w=10.27 l=2.08
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0053 pd=21.32 as=0 ps=0 w=10.27 l=2.08
X11 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.69455 pd=10.6 as=4.0053 ps=21.32 w=10.27 l=2.08
R0 VN.n0 VN.t3 155.004
R1 VN.n1 VN.t2 155.004
R2 VN.n0 VN.t1 154.458
R3 VN.n1 VN.t0 154.458
R4 VN VN.n1 50.6874
R5 VN VN.n0 6.97905
R6 VDD2.n2 VDD2.n0 100.314
R7 VDD2.n2 VDD2.n1 61.5131
R8 VDD2.n1 VDD2.t2 1.92845
R9 VDD2.n1 VDD2.t1 1.92845
R10 VDD2.n0 VDD2.t0 1.92845
R11 VDD2.n0 VDD2.t3 1.92845
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t3 46.7625
R14 VTAIL.n4 VTAIL.t5 46.7625
R15 VTAIL.n3 VTAIL.t7 46.7625
R16 VTAIL.n7 VTAIL.t6 46.7622
R17 VTAIL.n0 VTAIL.t4 46.7622
R18 VTAIL.n1 VTAIL.t0 46.7622
R19 VTAIL.n2 VTAIL.t1 46.7622
R20 VTAIL.n6 VTAIL.t2 46.7622
R21 VTAIL.n7 VTAIL.n6 23.2979
R22 VTAIL.n3 VTAIL.n2 23.2979
R23 VTAIL.n4 VTAIL.n3 2.07809
R24 VTAIL.n6 VTAIL.n5 2.07809
R25 VTAIL.n2 VTAIL.n1 2.07809
R26 VTAIL VTAIL.n0 1.09748
R27 VTAIL VTAIL.n7 0.981103
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n664 B.n663 585
R31 B.n665 B.n664 585
R32 B.n267 B.n98 585
R33 B.n266 B.n265 585
R34 B.n264 B.n263 585
R35 B.n262 B.n261 585
R36 B.n260 B.n259 585
R37 B.n258 B.n257 585
R38 B.n256 B.n255 585
R39 B.n254 B.n253 585
R40 B.n252 B.n251 585
R41 B.n250 B.n249 585
R42 B.n248 B.n247 585
R43 B.n246 B.n245 585
R44 B.n244 B.n243 585
R45 B.n242 B.n241 585
R46 B.n240 B.n239 585
R47 B.n238 B.n237 585
R48 B.n236 B.n235 585
R49 B.n234 B.n233 585
R50 B.n232 B.n231 585
R51 B.n230 B.n229 585
R52 B.n228 B.n227 585
R53 B.n226 B.n225 585
R54 B.n224 B.n223 585
R55 B.n222 B.n221 585
R56 B.n220 B.n219 585
R57 B.n218 B.n217 585
R58 B.n216 B.n215 585
R59 B.n214 B.n213 585
R60 B.n212 B.n211 585
R61 B.n210 B.n209 585
R62 B.n208 B.n207 585
R63 B.n206 B.n205 585
R64 B.n204 B.n203 585
R65 B.n202 B.n201 585
R66 B.n200 B.n199 585
R67 B.n198 B.n197 585
R68 B.n196 B.n195 585
R69 B.n194 B.n193 585
R70 B.n192 B.n191 585
R71 B.n190 B.n189 585
R72 B.n188 B.n187 585
R73 B.n186 B.n185 585
R74 B.n184 B.n183 585
R75 B.n182 B.n181 585
R76 B.n180 B.n179 585
R77 B.n177 B.n176 585
R78 B.n175 B.n174 585
R79 B.n173 B.n172 585
R80 B.n171 B.n170 585
R81 B.n169 B.n168 585
R82 B.n167 B.n166 585
R83 B.n165 B.n164 585
R84 B.n163 B.n162 585
R85 B.n161 B.n160 585
R86 B.n159 B.n158 585
R87 B.n157 B.n156 585
R88 B.n155 B.n154 585
R89 B.n153 B.n152 585
R90 B.n151 B.n150 585
R91 B.n149 B.n148 585
R92 B.n147 B.n146 585
R93 B.n145 B.n144 585
R94 B.n143 B.n142 585
R95 B.n141 B.n140 585
R96 B.n139 B.n138 585
R97 B.n137 B.n136 585
R98 B.n135 B.n134 585
R99 B.n133 B.n132 585
R100 B.n131 B.n130 585
R101 B.n129 B.n128 585
R102 B.n127 B.n126 585
R103 B.n125 B.n124 585
R104 B.n123 B.n122 585
R105 B.n121 B.n120 585
R106 B.n119 B.n118 585
R107 B.n117 B.n116 585
R108 B.n115 B.n114 585
R109 B.n113 B.n112 585
R110 B.n111 B.n110 585
R111 B.n109 B.n108 585
R112 B.n107 B.n106 585
R113 B.n105 B.n104 585
R114 B.n662 B.n56 585
R115 B.n666 B.n56 585
R116 B.n661 B.n55 585
R117 B.n667 B.n55 585
R118 B.n660 B.n659 585
R119 B.n659 B.n51 585
R120 B.n658 B.n50 585
R121 B.n673 B.n50 585
R122 B.n657 B.n49 585
R123 B.n674 B.n49 585
R124 B.n656 B.n48 585
R125 B.n675 B.n48 585
R126 B.n655 B.n654 585
R127 B.n654 B.n47 585
R128 B.n653 B.n43 585
R129 B.n681 B.n43 585
R130 B.n652 B.n42 585
R131 B.n682 B.n42 585
R132 B.n651 B.n41 585
R133 B.n683 B.n41 585
R134 B.n650 B.n649 585
R135 B.n649 B.n37 585
R136 B.n648 B.n36 585
R137 B.n689 B.n36 585
R138 B.n647 B.n35 585
R139 B.n690 B.n35 585
R140 B.n646 B.n34 585
R141 B.n691 B.n34 585
R142 B.n645 B.n644 585
R143 B.n644 B.n30 585
R144 B.n643 B.n29 585
R145 B.n697 B.n29 585
R146 B.n642 B.n28 585
R147 B.n698 B.n28 585
R148 B.n641 B.n27 585
R149 B.n699 B.n27 585
R150 B.n640 B.n639 585
R151 B.n639 B.n23 585
R152 B.n638 B.n22 585
R153 B.n705 B.n22 585
R154 B.n637 B.n21 585
R155 B.n706 B.n21 585
R156 B.n636 B.n20 585
R157 B.n707 B.n20 585
R158 B.n635 B.n634 585
R159 B.n634 B.n16 585
R160 B.n633 B.n15 585
R161 B.n713 B.n15 585
R162 B.n632 B.n14 585
R163 B.n714 B.n14 585
R164 B.n631 B.n13 585
R165 B.n715 B.n13 585
R166 B.n630 B.n629 585
R167 B.n629 B.n12 585
R168 B.n628 B.n627 585
R169 B.n628 B.n8 585
R170 B.n626 B.n7 585
R171 B.n722 B.n7 585
R172 B.n625 B.n6 585
R173 B.n723 B.n6 585
R174 B.n624 B.n5 585
R175 B.n724 B.n5 585
R176 B.n623 B.n622 585
R177 B.n622 B.n4 585
R178 B.n621 B.n268 585
R179 B.n621 B.n620 585
R180 B.n611 B.n269 585
R181 B.n270 B.n269 585
R182 B.n613 B.n612 585
R183 B.n614 B.n613 585
R184 B.n610 B.n274 585
R185 B.n278 B.n274 585
R186 B.n609 B.n608 585
R187 B.n608 B.n607 585
R188 B.n276 B.n275 585
R189 B.n277 B.n276 585
R190 B.n600 B.n599 585
R191 B.n601 B.n600 585
R192 B.n598 B.n283 585
R193 B.n283 B.n282 585
R194 B.n597 B.n596 585
R195 B.n596 B.n595 585
R196 B.n285 B.n284 585
R197 B.n286 B.n285 585
R198 B.n588 B.n587 585
R199 B.n589 B.n588 585
R200 B.n586 B.n291 585
R201 B.n291 B.n290 585
R202 B.n585 B.n584 585
R203 B.n584 B.n583 585
R204 B.n293 B.n292 585
R205 B.n294 B.n293 585
R206 B.n576 B.n575 585
R207 B.n577 B.n576 585
R208 B.n574 B.n299 585
R209 B.n299 B.n298 585
R210 B.n573 B.n572 585
R211 B.n572 B.n571 585
R212 B.n301 B.n300 585
R213 B.n302 B.n301 585
R214 B.n564 B.n563 585
R215 B.n565 B.n564 585
R216 B.n562 B.n307 585
R217 B.n307 B.n306 585
R218 B.n561 B.n560 585
R219 B.n560 B.n559 585
R220 B.n309 B.n308 585
R221 B.n552 B.n309 585
R222 B.n551 B.n550 585
R223 B.n553 B.n551 585
R224 B.n549 B.n314 585
R225 B.n314 B.n313 585
R226 B.n548 B.n547 585
R227 B.n547 B.n546 585
R228 B.n316 B.n315 585
R229 B.n317 B.n316 585
R230 B.n539 B.n538 585
R231 B.n540 B.n539 585
R232 B.n537 B.n322 585
R233 B.n322 B.n321 585
R234 B.n531 B.n530 585
R235 B.n529 B.n365 585
R236 B.n528 B.n364 585
R237 B.n533 B.n364 585
R238 B.n527 B.n526 585
R239 B.n525 B.n524 585
R240 B.n523 B.n522 585
R241 B.n521 B.n520 585
R242 B.n519 B.n518 585
R243 B.n517 B.n516 585
R244 B.n515 B.n514 585
R245 B.n513 B.n512 585
R246 B.n511 B.n510 585
R247 B.n509 B.n508 585
R248 B.n507 B.n506 585
R249 B.n505 B.n504 585
R250 B.n503 B.n502 585
R251 B.n501 B.n500 585
R252 B.n499 B.n498 585
R253 B.n497 B.n496 585
R254 B.n495 B.n494 585
R255 B.n493 B.n492 585
R256 B.n491 B.n490 585
R257 B.n489 B.n488 585
R258 B.n487 B.n486 585
R259 B.n485 B.n484 585
R260 B.n483 B.n482 585
R261 B.n481 B.n480 585
R262 B.n479 B.n478 585
R263 B.n477 B.n476 585
R264 B.n475 B.n474 585
R265 B.n473 B.n472 585
R266 B.n471 B.n470 585
R267 B.n469 B.n468 585
R268 B.n467 B.n466 585
R269 B.n465 B.n464 585
R270 B.n463 B.n462 585
R271 B.n461 B.n460 585
R272 B.n459 B.n458 585
R273 B.n457 B.n456 585
R274 B.n455 B.n454 585
R275 B.n453 B.n452 585
R276 B.n451 B.n450 585
R277 B.n449 B.n448 585
R278 B.n447 B.n446 585
R279 B.n445 B.n444 585
R280 B.n443 B.n442 585
R281 B.n440 B.n439 585
R282 B.n438 B.n437 585
R283 B.n436 B.n435 585
R284 B.n434 B.n433 585
R285 B.n432 B.n431 585
R286 B.n430 B.n429 585
R287 B.n428 B.n427 585
R288 B.n426 B.n425 585
R289 B.n424 B.n423 585
R290 B.n422 B.n421 585
R291 B.n420 B.n419 585
R292 B.n418 B.n417 585
R293 B.n416 B.n415 585
R294 B.n414 B.n413 585
R295 B.n412 B.n411 585
R296 B.n410 B.n409 585
R297 B.n408 B.n407 585
R298 B.n406 B.n405 585
R299 B.n404 B.n403 585
R300 B.n402 B.n401 585
R301 B.n400 B.n399 585
R302 B.n398 B.n397 585
R303 B.n396 B.n395 585
R304 B.n394 B.n393 585
R305 B.n392 B.n391 585
R306 B.n390 B.n389 585
R307 B.n388 B.n387 585
R308 B.n386 B.n385 585
R309 B.n384 B.n383 585
R310 B.n382 B.n381 585
R311 B.n380 B.n379 585
R312 B.n378 B.n377 585
R313 B.n376 B.n375 585
R314 B.n374 B.n373 585
R315 B.n372 B.n371 585
R316 B.n324 B.n323 585
R317 B.n536 B.n535 585
R318 B.n320 B.n319 585
R319 B.n321 B.n320 585
R320 B.n542 B.n541 585
R321 B.n541 B.n540 585
R322 B.n543 B.n318 585
R323 B.n318 B.n317 585
R324 B.n545 B.n544 585
R325 B.n546 B.n545 585
R326 B.n312 B.n311 585
R327 B.n313 B.n312 585
R328 B.n555 B.n554 585
R329 B.n554 B.n553 585
R330 B.n556 B.n310 585
R331 B.n552 B.n310 585
R332 B.n558 B.n557 585
R333 B.n559 B.n558 585
R334 B.n305 B.n304 585
R335 B.n306 B.n305 585
R336 B.n567 B.n566 585
R337 B.n566 B.n565 585
R338 B.n568 B.n303 585
R339 B.n303 B.n302 585
R340 B.n570 B.n569 585
R341 B.n571 B.n570 585
R342 B.n297 B.n296 585
R343 B.n298 B.n297 585
R344 B.n579 B.n578 585
R345 B.n578 B.n577 585
R346 B.n580 B.n295 585
R347 B.n295 B.n294 585
R348 B.n582 B.n581 585
R349 B.n583 B.n582 585
R350 B.n289 B.n288 585
R351 B.n290 B.n289 585
R352 B.n591 B.n590 585
R353 B.n590 B.n589 585
R354 B.n592 B.n287 585
R355 B.n287 B.n286 585
R356 B.n594 B.n593 585
R357 B.n595 B.n594 585
R358 B.n281 B.n280 585
R359 B.n282 B.n281 585
R360 B.n603 B.n602 585
R361 B.n602 B.n601 585
R362 B.n604 B.n279 585
R363 B.n279 B.n277 585
R364 B.n606 B.n605 585
R365 B.n607 B.n606 585
R366 B.n273 B.n272 585
R367 B.n278 B.n273 585
R368 B.n616 B.n615 585
R369 B.n615 B.n614 585
R370 B.n617 B.n271 585
R371 B.n271 B.n270 585
R372 B.n619 B.n618 585
R373 B.n620 B.n619 585
R374 B.n3 B.n0 585
R375 B.n4 B.n3 585
R376 B.n721 B.n1 585
R377 B.n722 B.n721 585
R378 B.n720 B.n719 585
R379 B.n720 B.n8 585
R380 B.n718 B.n9 585
R381 B.n12 B.n9 585
R382 B.n717 B.n716 585
R383 B.n716 B.n715 585
R384 B.n11 B.n10 585
R385 B.n714 B.n11 585
R386 B.n712 B.n711 585
R387 B.n713 B.n712 585
R388 B.n710 B.n17 585
R389 B.n17 B.n16 585
R390 B.n709 B.n708 585
R391 B.n708 B.n707 585
R392 B.n19 B.n18 585
R393 B.n706 B.n19 585
R394 B.n704 B.n703 585
R395 B.n705 B.n704 585
R396 B.n702 B.n24 585
R397 B.n24 B.n23 585
R398 B.n701 B.n700 585
R399 B.n700 B.n699 585
R400 B.n26 B.n25 585
R401 B.n698 B.n26 585
R402 B.n696 B.n695 585
R403 B.n697 B.n696 585
R404 B.n694 B.n31 585
R405 B.n31 B.n30 585
R406 B.n693 B.n692 585
R407 B.n692 B.n691 585
R408 B.n33 B.n32 585
R409 B.n690 B.n33 585
R410 B.n688 B.n687 585
R411 B.n689 B.n688 585
R412 B.n686 B.n38 585
R413 B.n38 B.n37 585
R414 B.n685 B.n684 585
R415 B.n684 B.n683 585
R416 B.n40 B.n39 585
R417 B.n682 B.n40 585
R418 B.n680 B.n679 585
R419 B.n681 B.n680 585
R420 B.n678 B.n44 585
R421 B.n47 B.n44 585
R422 B.n677 B.n676 585
R423 B.n676 B.n675 585
R424 B.n46 B.n45 585
R425 B.n674 B.n46 585
R426 B.n672 B.n671 585
R427 B.n673 B.n672 585
R428 B.n670 B.n52 585
R429 B.n52 B.n51 585
R430 B.n669 B.n668 585
R431 B.n668 B.n667 585
R432 B.n54 B.n53 585
R433 B.n666 B.n54 585
R434 B.n725 B.n724 585
R435 B.n723 B.n2 585
R436 B.n104 B.n54 449.257
R437 B.n664 B.n56 449.257
R438 B.n535 B.n322 449.257
R439 B.n531 B.n320 449.257
R440 B.n102 B.t15 326.094
R441 B.n99 B.t8 326.094
R442 B.n369 B.t12 326.094
R443 B.n366 B.t4 326.094
R444 B.n665 B.n97 256.663
R445 B.n665 B.n96 256.663
R446 B.n665 B.n95 256.663
R447 B.n665 B.n94 256.663
R448 B.n665 B.n93 256.663
R449 B.n665 B.n92 256.663
R450 B.n665 B.n91 256.663
R451 B.n665 B.n90 256.663
R452 B.n665 B.n89 256.663
R453 B.n665 B.n88 256.663
R454 B.n665 B.n87 256.663
R455 B.n665 B.n86 256.663
R456 B.n665 B.n85 256.663
R457 B.n665 B.n84 256.663
R458 B.n665 B.n83 256.663
R459 B.n665 B.n82 256.663
R460 B.n665 B.n81 256.663
R461 B.n665 B.n80 256.663
R462 B.n665 B.n79 256.663
R463 B.n665 B.n78 256.663
R464 B.n665 B.n77 256.663
R465 B.n665 B.n76 256.663
R466 B.n665 B.n75 256.663
R467 B.n665 B.n74 256.663
R468 B.n665 B.n73 256.663
R469 B.n665 B.n72 256.663
R470 B.n665 B.n71 256.663
R471 B.n665 B.n70 256.663
R472 B.n665 B.n69 256.663
R473 B.n665 B.n68 256.663
R474 B.n665 B.n67 256.663
R475 B.n665 B.n66 256.663
R476 B.n665 B.n65 256.663
R477 B.n665 B.n64 256.663
R478 B.n665 B.n63 256.663
R479 B.n665 B.n62 256.663
R480 B.n665 B.n61 256.663
R481 B.n665 B.n60 256.663
R482 B.n665 B.n59 256.663
R483 B.n665 B.n58 256.663
R484 B.n665 B.n57 256.663
R485 B.n533 B.n532 256.663
R486 B.n533 B.n325 256.663
R487 B.n533 B.n326 256.663
R488 B.n533 B.n327 256.663
R489 B.n533 B.n328 256.663
R490 B.n533 B.n329 256.663
R491 B.n533 B.n330 256.663
R492 B.n533 B.n331 256.663
R493 B.n533 B.n332 256.663
R494 B.n533 B.n333 256.663
R495 B.n533 B.n334 256.663
R496 B.n533 B.n335 256.663
R497 B.n533 B.n336 256.663
R498 B.n533 B.n337 256.663
R499 B.n533 B.n338 256.663
R500 B.n533 B.n339 256.663
R501 B.n533 B.n340 256.663
R502 B.n533 B.n341 256.663
R503 B.n533 B.n342 256.663
R504 B.n533 B.n343 256.663
R505 B.n533 B.n344 256.663
R506 B.n533 B.n345 256.663
R507 B.n533 B.n346 256.663
R508 B.n533 B.n347 256.663
R509 B.n533 B.n348 256.663
R510 B.n533 B.n349 256.663
R511 B.n533 B.n350 256.663
R512 B.n533 B.n351 256.663
R513 B.n533 B.n352 256.663
R514 B.n533 B.n353 256.663
R515 B.n533 B.n354 256.663
R516 B.n533 B.n355 256.663
R517 B.n533 B.n356 256.663
R518 B.n533 B.n357 256.663
R519 B.n533 B.n358 256.663
R520 B.n533 B.n359 256.663
R521 B.n533 B.n360 256.663
R522 B.n533 B.n361 256.663
R523 B.n533 B.n362 256.663
R524 B.n533 B.n363 256.663
R525 B.n534 B.n533 256.663
R526 B.n727 B.n726 256.663
R527 B.n108 B.n107 163.367
R528 B.n112 B.n111 163.367
R529 B.n116 B.n115 163.367
R530 B.n120 B.n119 163.367
R531 B.n124 B.n123 163.367
R532 B.n128 B.n127 163.367
R533 B.n132 B.n131 163.367
R534 B.n136 B.n135 163.367
R535 B.n140 B.n139 163.367
R536 B.n144 B.n143 163.367
R537 B.n148 B.n147 163.367
R538 B.n152 B.n151 163.367
R539 B.n156 B.n155 163.367
R540 B.n160 B.n159 163.367
R541 B.n164 B.n163 163.367
R542 B.n168 B.n167 163.367
R543 B.n172 B.n171 163.367
R544 B.n176 B.n175 163.367
R545 B.n181 B.n180 163.367
R546 B.n185 B.n184 163.367
R547 B.n189 B.n188 163.367
R548 B.n193 B.n192 163.367
R549 B.n197 B.n196 163.367
R550 B.n201 B.n200 163.367
R551 B.n205 B.n204 163.367
R552 B.n209 B.n208 163.367
R553 B.n213 B.n212 163.367
R554 B.n217 B.n216 163.367
R555 B.n221 B.n220 163.367
R556 B.n225 B.n224 163.367
R557 B.n229 B.n228 163.367
R558 B.n233 B.n232 163.367
R559 B.n237 B.n236 163.367
R560 B.n241 B.n240 163.367
R561 B.n245 B.n244 163.367
R562 B.n249 B.n248 163.367
R563 B.n253 B.n252 163.367
R564 B.n257 B.n256 163.367
R565 B.n261 B.n260 163.367
R566 B.n265 B.n264 163.367
R567 B.n664 B.n98 163.367
R568 B.n539 B.n322 163.367
R569 B.n539 B.n316 163.367
R570 B.n547 B.n316 163.367
R571 B.n547 B.n314 163.367
R572 B.n551 B.n314 163.367
R573 B.n551 B.n309 163.367
R574 B.n560 B.n309 163.367
R575 B.n560 B.n307 163.367
R576 B.n564 B.n307 163.367
R577 B.n564 B.n301 163.367
R578 B.n572 B.n301 163.367
R579 B.n572 B.n299 163.367
R580 B.n576 B.n299 163.367
R581 B.n576 B.n293 163.367
R582 B.n584 B.n293 163.367
R583 B.n584 B.n291 163.367
R584 B.n588 B.n291 163.367
R585 B.n588 B.n285 163.367
R586 B.n596 B.n285 163.367
R587 B.n596 B.n283 163.367
R588 B.n600 B.n283 163.367
R589 B.n600 B.n276 163.367
R590 B.n608 B.n276 163.367
R591 B.n608 B.n274 163.367
R592 B.n613 B.n274 163.367
R593 B.n613 B.n269 163.367
R594 B.n621 B.n269 163.367
R595 B.n622 B.n621 163.367
R596 B.n622 B.n5 163.367
R597 B.n6 B.n5 163.367
R598 B.n7 B.n6 163.367
R599 B.n628 B.n7 163.367
R600 B.n629 B.n628 163.367
R601 B.n629 B.n13 163.367
R602 B.n14 B.n13 163.367
R603 B.n15 B.n14 163.367
R604 B.n634 B.n15 163.367
R605 B.n634 B.n20 163.367
R606 B.n21 B.n20 163.367
R607 B.n22 B.n21 163.367
R608 B.n639 B.n22 163.367
R609 B.n639 B.n27 163.367
R610 B.n28 B.n27 163.367
R611 B.n29 B.n28 163.367
R612 B.n644 B.n29 163.367
R613 B.n644 B.n34 163.367
R614 B.n35 B.n34 163.367
R615 B.n36 B.n35 163.367
R616 B.n649 B.n36 163.367
R617 B.n649 B.n41 163.367
R618 B.n42 B.n41 163.367
R619 B.n43 B.n42 163.367
R620 B.n654 B.n43 163.367
R621 B.n654 B.n48 163.367
R622 B.n49 B.n48 163.367
R623 B.n50 B.n49 163.367
R624 B.n659 B.n50 163.367
R625 B.n659 B.n55 163.367
R626 B.n56 B.n55 163.367
R627 B.n365 B.n364 163.367
R628 B.n526 B.n364 163.367
R629 B.n524 B.n523 163.367
R630 B.n520 B.n519 163.367
R631 B.n516 B.n515 163.367
R632 B.n512 B.n511 163.367
R633 B.n508 B.n507 163.367
R634 B.n504 B.n503 163.367
R635 B.n500 B.n499 163.367
R636 B.n496 B.n495 163.367
R637 B.n492 B.n491 163.367
R638 B.n488 B.n487 163.367
R639 B.n484 B.n483 163.367
R640 B.n480 B.n479 163.367
R641 B.n476 B.n475 163.367
R642 B.n472 B.n471 163.367
R643 B.n468 B.n467 163.367
R644 B.n464 B.n463 163.367
R645 B.n460 B.n459 163.367
R646 B.n456 B.n455 163.367
R647 B.n452 B.n451 163.367
R648 B.n448 B.n447 163.367
R649 B.n444 B.n443 163.367
R650 B.n439 B.n438 163.367
R651 B.n435 B.n434 163.367
R652 B.n431 B.n430 163.367
R653 B.n427 B.n426 163.367
R654 B.n423 B.n422 163.367
R655 B.n419 B.n418 163.367
R656 B.n415 B.n414 163.367
R657 B.n411 B.n410 163.367
R658 B.n407 B.n406 163.367
R659 B.n403 B.n402 163.367
R660 B.n399 B.n398 163.367
R661 B.n395 B.n394 163.367
R662 B.n391 B.n390 163.367
R663 B.n387 B.n386 163.367
R664 B.n383 B.n382 163.367
R665 B.n379 B.n378 163.367
R666 B.n375 B.n374 163.367
R667 B.n371 B.n324 163.367
R668 B.n541 B.n320 163.367
R669 B.n541 B.n318 163.367
R670 B.n545 B.n318 163.367
R671 B.n545 B.n312 163.367
R672 B.n554 B.n312 163.367
R673 B.n554 B.n310 163.367
R674 B.n558 B.n310 163.367
R675 B.n558 B.n305 163.367
R676 B.n566 B.n305 163.367
R677 B.n566 B.n303 163.367
R678 B.n570 B.n303 163.367
R679 B.n570 B.n297 163.367
R680 B.n578 B.n297 163.367
R681 B.n578 B.n295 163.367
R682 B.n582 B.n295 163.367
R683 B.n582 B.n289 163.367
R684 B.n590 B.n289 163.367
R685 B.n590 B.n287 163.367
R686 B.n594 B.n287 163.367
R687 B.n594 B.n281 163.367
R688 B.n602 B.n281 163.367
R689 B.n602 B.n279 163.367
R690 B.n606 B.n279 163.367
R691 B.n606 B.n273 163.367
R692 B.n615 B.n273 163.367
R693 B.n615 B.n271 163.367
R694 B.n619 B.n271 163.367
R695 B.n619 B.n3 163.367
R696 B.n725 B.n3 163.367
R697 B.n721 B.n2 163.367
R698 B.n721 B.n720 163.367
R699 B.n720 B.n9 163.367
R700 B.n716 B.n9 163.367
R701 B.n716 B.n11 163.367
R702 B.n712 B.n11 163.367
R703 B.n712 B.n17 163.367
R704 B.n708 B.n17 163.367
R705 B.n708 B.n19 163.367
R706 B.n704 B.n19 163.367
R707 B.n704 B.n24 163.367
R708 B.n700 B.n24 163.367
R709 B.n700 B.n26 163.367
R710 B.n696 B.n26 163.367
R711 B.n696 B.n31 163.367
R712 B.n692 B.n31 163.367
R713 B.n692 B.n33 163.367
R714 B.n688 B.n33 163.367
R715 B.n688 B.n38 163.367
R716 B.n684 B.n38 163.367
R717 B.n684 B.n40 163.367
R718 B.n680 B.n40 163.367
R719 B.n680 B.n44 163.367
R720 B.n676 B.n44 163.367
R721 B.n676 B.n46 163.367
R722 B.n672 B.n46 163.367
R723 B.n672 B.n52 163.367
R724 B.n668 B.n52 163.367
R725 B.n668 B.n54 163.367
R726 B.n99 B.t10 116.162
R727 B.n369 B.t14 116.162
R728 B.n102 B.t16 116.15
R729 B.n366 B.t7 116.15
R730 B.n533 B.n321 81.3771
R731 B.n666 B.n665 81.3771
R732 B.n104 B.n57 71.676
R733 B.n108 B.n58 71.676
R734 B.n112 B.n59 71.676
R735 B.n116 B.n60 71.676
R736 B.n120 B.n61 71.676
R737 B.n124 B.n62 71.676
R738 B.n128 B.n63 71.676
R739 B.n132 B.n64 71.676
R740 B.n136 B.n65 71.676
R741 B.n140 B.n66 71.676
R742 B.n144 B.n67 71.676
R743 B.n148 B.n68 71.676
R744 B.n152 B.n69 71.676
R745 B.n156 B.n70 71.676
R746 B.n160 B.n71 71.676
R747 B.n164 B.n72 71.676
R748 B.n168 B.n73 71.676
R749 B.n172 B.n74 71.676
R750 B.n176 B.n75 71.676
R751 B.n181 B.n76 71.676
R752 B.n185 B.n77 71.676
R753 B.n189 B.n78 71.676
R754 B.n193 B.n79 71.676
R755 B.n197 B.n80 71.676
R756 B.n201 B.n81 71.676
R757 B.n205 B.n82 71.676
R758 B.n209 B.n83 71.676
R759 B.n213 B.n84 71.676
R760 B.n217 B.n85 71.676
R761 B.n221 B.n86 71.676
R762 B.n225 B.n87 71.676
R763 B.n229 B.n88 71.676
R764 B.n233 B.n89 71.676
R765 B.n237 B.n90 71.676
R766 B.n241 B.n91 71.676
R767 B.n245 B.n92 71.676
R768 B.n249 B.n93 71.676
R769 B.n253 B.n94 71.676
R770 B.n257 B.n95 71.676
R771 B.n261 B.n96 71.676
R772 B.n265 B.n97 71.676
R773 B.n98 B.n97 71.676
R774 B.n264 B.n96 71.676
R775 B.n260 B.n95 71.676
R776 B.n256 B.n94 71.676
R777 B.n252 B.n93 71.676
R778 B.n248 B.n92 71.676
R779 B.n244 B.n91 71.676
R780 B.n240 B.n90 71.676
R781 B.n236 B.n89 71.676
R782 B.n232 B.n88 71.676
R783 B.n228 B.n87 71.676
R784 B.n224 B.n86 71.676
R785 B.n220 B.n85 71.676
R786 B.n216 B.n84 71.676
R787 B.n212 B.n83 71.676
R788 B.n208 B.n82 71.676
R789 B.n204 B.n81 71.676
R790 B.n200 B.n80 71.676
R791 B.n196 B.n79 71.676
R792 B.n192 B.n78 71.676
R793 B.n188 B.n77 71.676
R794 B.n184 B.n76 71.676
R795 B.n180 B.n75 71.676
R796 B.n175 B.n74 71.676
R797 B.n171 B.n73 71.676
R798 B.n167 B.n72 71.676
R799 B.n163 B.n71 71.676
R800 B.n159 B.n70 71.676
R801 B.n155 B.n69 71.676
R802 B.n151 B.n68 71.676
R803 B.n147 B.n67 71.676
R804 B.n143 B.n66 71.676
R805 B.n139 B.n65 71.676
R806 B.n135 B.n64 71.676
R807 B.n131 B.n63 71.676
R808 B.n127 B.n62 71.676
R809 B.n123 B.n61 71.676
R810 B.n119 B.n60 71.676
R811 B.n115 B.n59 71.676
R812 B.n111 B.n58 71.676
R813 B.n107 B.n57 71.676
R814 B.n532 B.n531 71.676
R815 B.n526 B.n325 71.676
R816 B.n523 B.n326 71.676
R817 B.n519 B.n327 71.676
R818 B.n515 B.n328 71.676
R819 B.n511 B.n329 71.676
R820 B.n507 B.n330 71.676
R821 B.n503 B.n331 71.676
R822 B.n499 B.n332 71.676
R823 B.n495 B.n333 71.676
R824 B.n491 B.n334 71.676
R825 B.n487 B.n335 71.676
R826 B.n483 B.n336 71.676
R827 B.n479 B.n337 71.676
R828 B.n475 B.n338 71.676
R829 B.n471 B.n339 71.676
R830 B.n467 B.n340 71.676
R831 B.n463 B.n341 71.676
R832 B.n459 B.n342 71.676
R833 B.n455 B.n343 71.676
R834 B.n451 B.n344 71.676
R835 B.n447 B.n345 71.676
R836 B.n443 B.n346 71.676
R837 B.n438 B.n347 71.676
R838 B.n434 B.n348 71.676
R839 B.n430 B.n349 71.676
R840 B.n426 B.n350 71.676
R841 B.n422 B.n351 71.676
R842 B.n418 B.n352 71.676
R843 B.n414 B.n353 71.676
R844 B.n410 B.n354 71.676
R845 B.n406 B.n355 71.676
R846 B.n402 B.n356 71.676
R847 B.n398 B.n357 71.676
R848 B.n394 B.n358 71.676
R849 B.n390 B.n359 71.676
R850 B.n386 B.n360 71.676
R851 B.n382 B.n361 71.676
R852 B.n378 B.n362 71.676
R853 B.n374 B.n363 71.676
R854 B.n534 B.n324 71.676
R855 B.n532 B.n365 71.676
R856 B.n524 B.n325 71.676
R857 B.n520 B.n326 71.676
R858 B.n516 B.n327 71.676
R859 B.n512 B.n328 71.676
R860 B.n508 B.n329 71.676
R861 B.n504 B.n330 71.676
R862 B.n500 B.n331 71.676
R863 B.n496 B.n332 71.676
R864 B.n492 B.n333 71.676
R865 B.n488 B.n334 71.676
R866 B.n484 B.n335 71.676
R867 B.n480 B.n336 71.676
R868 B.n476 B.n337 71.676
R869 B.n472 B.n338 71.676
R870 B.n468 B.n339 71.676
R871 B.n464 B.n340 71.676
R872 B.n460 B.n341 71.676
R873 B.n456 B.n342 71.676
R874 B.n452 B.n343 71.676
R875 B.n448 B.n344 71.676
R876 B.n444 B.n345 71.676
R877 B.n439 B.n346 71.676
R878 B.n435 B.n347 71.676
R879 B.n431 B.n348 71.676
R880 B.n427 B.n349 71.676
R881 B.n423 B.n350 71.676
R882 B.n419 B.n351 71.676
R883 B.n415 B.n352 71.676
R884 B.n411 B.n353 71.676
R885 B.n407 B.n354 71.676
R886 B.n403 B.n355 71.676
R887 B.n399 B.n356 71.676
R888 B.n395 B.n357 71.676
R889 B.n391 B.n358 71.676
R890 B.n387 B.n359 71.676
R891 B.n383 B.n360 71.676
R892 B.n379 B.n361 71.676
R893 B.n375 B.n362 71.676
R894 B.n371 B.n363 71.676
R895 B.n535 B.n534 71.676
R896 B.n726 B.n725 71.676
R897 B.n726 B.n2 71.676
R898 B.n100 B.t11 69.4229
R899 B.n370 B.t13 69.4229
R900 B.n103 B.t17 69.4102
R901 B.n367 B.t6 69.4102
R902 B.n178 B.n103 59.5399
R903 B.n101 B.n100 59.5399
R904 B.n441 B.n370 59.5399
R905 B.n368 B.n367 59.5399
R906 B.n540 B.n321 48.1189
R907 B.n540 B.n317 48.1189
R908 B.n546 B.n317 48.1189
R909 B.n546 B.n313 48.1189
R910 B.n553 B.n313 48.1189
R911 B.n553 B.n552 48.1189
R912 B.n559 B.n306 48.1189
R913 B.n565 B.n306 48.1189
R914 B.n565 B.n302 48.1189
R915 B.n571 B.n302 48.1189
R916 B.n571 B.n298 48.1189
R917 B.n577 B.n298 48.1189
R918 B.n577 B.n294 48.1189
R919 B.n583 B.n294 48.1189
R920 B.n583 B.n290 48.1189
R921 B.n589 B.n290 48.1189
R922 B.n595 B.n286 48.1189
R923 B.n595 B.n282 48.1189
R924 B.n601 B.n282 48.1189
R925 B.n601 B.n277 48.1189
R926 B.n607 B.n277 48.1189
R927 B.n607 B.n278 48.1189
R928 B.n614 B.n270 48.1189
R929 B.n620 B.n270 48.1189
R930 B.n620 B.n4 48.1189
R931 B.n724 B.n4 48.1189
R932 B.n724 B.n723 48.1189
R933 B.n723 B.n722 48.1189
R934 B.n722 B.n8 48.1189
R935 B.n12 B.n8 48.1189
R936 B.n715 B.n12 48.1189
R937 B.n714 B.n713 48.1189
R938 B.n713 B.n16 48.1189
R939 B.n707 B.n16 48.1189
R940 B.n707 B.n706 48.1189
R941 B.n706 B.n705 48.1189
R942 B.n705 B.n23 48.1189
R943 B.n699 B.n698 48.1189
R944 B.n698 B.n697 48.1189
R945 B.n697 B.n30 48.1189
R946 B.n691 B.n30 48.1189
R947 B.n691 B.n690 48.1189
R948 B.n690 B.n689 48.1189
R949 B.n689 B.n37 48.1189
R950 B.n683 B.n37 48.1189
R951 B.n683 B.n682 48.1189
R952 B.n682 B.n681 48.1189
R953 B.n675 B.n47 48.1189
R954 B.n675 B.n674 48.1189
R955 B.n674 B.n673 48.1189
R956 B.n673 B.n51 48.1189
R957 B.n667 B.n51 48.1189
R958 B.n667 B.n666 48.1189
R959 B.n103 B.n102 46.7399
R960 B.n100 B.n99 46.7399
R961 B.n370 B.n369 46.7399
R962 B.n367 B.n366 46.7399
R963 B.n552 B.t5 46.7036
R964 B.n47 B.t9 46.7036
R965 B.t1 B.n286 35.3817
R966 B.t2 B.n23 35.3817
R967 B.n614 B.t0 31.1359
R968 B.n715 B.t3 31.1359
R969 B.n530 B.n319 29.1907
R970 B.n537 B.n536 29.1907
R971 B.n663 B.n662 29.1907
R972 B.n105 B.n53 29.1907
R973 B B.n727 18.0485
R974 B.n278 B.t0 16.9835
R975 B.t3 B.n714 16.9835
R976 B.n589 B.t1 12.7377
R977 B.n699 B.t2 12.7377
R978 B.n542 B.n319 10.6151
R979 B.n543 B.n542 10.6151
R980 B.n544 B.n543 10.6151
R981 B.n544 B.n311 10.6151
R982 B.n555 B.n311 10.6151
R983 B.n556 B.n555 10.6151
R984 B.n557 B.n556 10.6151
R985 B.n557 B.n304 10.6151
R986 B.n567 B.n304 10.6151
R987 B.n568 B.n567 10.6151
R988 B.n569 B.n568 10.6151
R989 B.n569 B.n296 10.6151
R990 B.n579 B.n296 10.6151
R991 B.n580 B.n579 10.6151
R992 B.n581 B.n580 10.6151
R993 B.n581 B.n288 10.6151
R994 B.n591 B.n288 10.6151
R995 B.n592 B.n591 10.6151
R996 B.n593 B.n592 10.6151
R997 B.n593 B.n280 10.6151
R998 B.n603 B.n280 10.6151
R999 B.n604 B.n603 10.6151
R1000 B.n605 B.n604 10.6151
R1001 B.n605 B.n272 10.6151
R1002 B.n616 B.n272 10.6151
R1003 B.n617 B.n616 10.6151
R1004 B.n618 B.n617 10.6151
R1005 B.n618 B.n0 10.6151
R1006 B.n530 B.n529 10.6151
R1007 B.n529 B.n528 10.6151
R1008 B.n528 B.n527 10.6151
R1009 B.n527 B.n525 10.6151
R1010 B.n525 B.n522 10.6151
R1011 B.n522 B.n521 10.6151
R1012 B.n521 B.n518 10.6151
R1013 B.n518 B.n517 10.6151
R1014 B.n517 B.n514 10.6151
R1015 B.n514 B.n513 10.6151
R1016 B.n513 B.n510 10.6151
R1017 B.n510 B.n509 10.6151
R1018 B.n509 B.n506 10.6151
R1019 B.n506 B.n505 10.6151
R1020 B.n505 B.n502 10.6151
R1021 B.n502 B.n501 10.6151
R1022 B.n501 B.n498 10.6151
R1023 B.n498 B.n497 10.6151
R1024 B.n497 B.n494 10.6151
R1025 B.n494 B.n493 10.6151
R1026 B.n493 B.n490 10.6151
R1027 B.n490 B.n489 10.6151
R1028 B.n489 B.n486 10.6151
R1029 B.n486 B.n485 10.6151
R1030 B.n485 B.n482 10.6151
R1031 B.n482 B.n481 10.6151
R1032 B.n481 B.n478 10.6151
R1033 B.n478 B.n477 10.6151
R1034 B.n477 B.n474 10.6151
R1035 B.n474 B.n473 10.6151
R1036 B.n473 B.n470 10.6151
R1037 B.n470 B.n469 10.6151
R1038 B.n469 B.n466 10.6151
R1039 B.n466 B.n465 10.6151
R1040 B.n465 B.n462 10.6151
R1041 B.n462 B.n461 10.6151
R1042 B.n458 B.n457 10.6151
R1043 B.n457 B.n454 10.6151
R1044 B.n454 B.n453 10.6151
R1045 B.n453 B.n450 10.6151
R1046 B.n450 B.n449 10.6151
R1047 B.n449 B.n446 10.6151
R1048 B.n446 B.n445 10.6151
R1049 B.n445 B.n442 10.6151
R1050 B.n440 B.n437 10.6151
R1051 B.n437 B.n436 10.6151
R1052 B.n436 B.n433 10.6151
R1053 B.n433 B.n432 10.6151
R1054 B.n432 B.n429 10.6151
R1055 B.n429 B.n428 10.6151
R1056 B.n428 B.n425 10.6151
R1057 B.n425 B.n424 10.6151
R1058 B.n424 B.n421 10.6151
R1059 B.n421 B.n420 10.6151
R1060 B.n420 B.n417 10.6151
R1061 B.n417 B.n416 10.6151
R1062 B.n416 B.n413 10.6151
R1063 B.n413 B.n412 10.6151
R1064 B.n412 B.n409 10.6151
R1065 B.n409 B.n408 10.6151
R1066 B.n408 B.n405 10.6151
R1067 B.n405 B.n404 10.6151
R1068 B.n404 B.n401 10.6151
R1069 B.n401 B.n400 10.6151
R1070 B.n400 B.n397 10.6151
R1071 B.n397 B.n396 10.6151
R1072 B.n396 B.n393 10.6151
R1073 B.n393 B.n392 10.6151
R1074 B.n392 B.n389 10.6151
R1075 B.n389 B.n388 10.6151
R1076 B.n388 B.n385 10.6151
R1077 B.n385 B.n384 10.6151
R1078 B.n384 B.n381 10.6151
R1079 B.n381 B.n380 10.6151
R1080 B.n380 B.n377 10.6151
R1081 B.n377 B.n376 10.6151
R1082 B.n376 B.n373 10.6151
R1083 B.n373 B.n372 10.6151
R1084 B.n372 B.n323 10.6151
R1085 B.n536 B.n323 10.6151
R1086 B.n538 B.n537 10.6151
R1087 B.n538 B.n315 10.6151
R1088 B.n548 B.n315 10.6151
R1089 B.n549 B.n548 10.6151
R1090 B.n550 B.n549 10.6151
R1091 B.n550 B.n308 10.6151
R1092 B.n561 B.n308 10.6151
R1093 B.n562 B.n561 10.6151
R1094 B.n563 B.n562 10.6151
R1095 B.n563 B.n300 10.6151
R1096 B.n573 B.n300 10.6151
R1097 B.n574 B.n573 10.6151
R1098 B.n575 B.n574 10.6151
R1099 B.n575 B.n292 10.6151
R1100 B.n585 B.n292 10.6151
R1101 B.n586 B.n585 10.6151
R1102 B.n587 B.n586 10.6151
R1103 B.n587 B.n284 10.6151
R1104 B.n597 B.n284 10.6151
R1105 B.n598 B.n597 10.6151
R1106 B.n599 B.n598 10.6151
R1107 B.n599 B.n275 10.6151
R1108 B.n609 B.n275 10.6151
R1109 B.n610 B.n609 10.6151
R1110 B.n612 B.n610 10.6151
R1111 B.n612 B.n611 10.6151
R1112 B.n611 B.n268 10.6151
R1113 B.n623 B.n268 10.6151
R1114 B.n624 B.n623 10.6151
R1115 B.n625 B.n624 10.6151
R1116 B.n626 B.n625 10.6151
R1117 B.n627 B.n626 10.6151
R1118 B.n630 B.n627 10.6151
R1119 B.n631 B.n630 10.6151
R1120 B.n632 B.n631 10.6151
R1121 B.n633 B.n632 10.6151
R1122 B.n635 B.n633 10.6151
R1123 B.n636 B.n635 10.6151
R1124 B.n637 B.n636 10.6151
R1125 B.n638 B.n637 10.6151
R1126 B.n640 B.n638 10.6151
R1127 B.n641 B.n640 10.6151
R1128 B.n642 B.n641 10.6151
R1129 B.n643 B.n642 10.6151
R1130 B.n645 B.n643 10.6151
R1131 B.n646 B.n645 10.6151
R1132 B.n647 B.n646 10.6151
R1133 B.n648 B.n647 10.6151
R1134 B.n650 B.n648 10.6151
R1135 B.n651 B.n650 10.6151
R1136 B.n652 B.n651 10.6151
R1137 B.n653 B.n652 10.6151
R1138 B.n655 B.n653 10.6151
R1139 B.n656 B.n655 10.6151
R1140 B.n657 B.n656 10.6151
R1141 B.n658 B.n657 10.6151
R1142 B.n660 B.n658 10.6151
R1143 B.n661 B.n660 10.6151
R1144 B.n662 B.n661 10.6151
R1145 B.n719 B.n1 10.6151
R1146 B.n719 B.n718 10.6151
R1147 B.n718 B.n717 10.6151
R1148 B.n717 B.n10 10.6151
R1149 B.n711 B.n10 10.6151
R1150 B.n711 B.n710 10.6151
R1151 B.n710 B.n709 10.6151
R1152 B.n709 B.n18 10.6151
R1153 B.n703 B.n18 10.6151
R1154 B.n703 B.n702 10.6151
R1155 B.n702 B.n701 10.6151
R1156 B.n701 B.n25 10.6151
R1157 B.n695 B.n25 10.6151
R1158 B.n695 B.n694 10.6151
R1159 B.n694 B.n693 10.6151
R1160 B.n693 B.n32 10.6151
R1161 B.n687 B.n32 10.6151
R1162 B.n687 B.n686 10.6151
R1163 B.n686 B.n685 10.6151
R1164 B.n685 B.n39 10.6151
R1165 B.n679 B.n39 10.6151
R1166 B.n679 B.n678 10.6151
R1167 B.n678 B.n677 10.6151
R1168 B.n677 B.n45 10.6151
R1169 B.n671 B.n45 10.6151
R1170 B.n671 B.n670 10.6151
R1171 B.n670 B.n669 10.6151
R1172 B.n669 B.n53 10.6151
R1173 B.n106 B.n105 10.6151
R1174 B.n109 B.n106 10.6151
R1175 B.n110 B.n109 10.6151
R1176 B.n113 B.n110 10.6151
R1177 B.n114 B.n113 10.6151
R1178 B.n117 B.n114 10.6151
R1179 B.n118 B.n117 10.6151
R1180 B.n121 B.n118 10.6151
R1181 B.n122 B.n121 10.6151
R1182 B.n125 B.n122 10.6151
R1183 B.n126 B.n125 10.6151
R1184 B.n129 B.n126 10.6151
R1185 B.n130 B.n129 10.6151
R1186 B.n133 B.n130 10.6151
R1187 B.n134 B.n133 10.6151
R1188 B.n137 B.n134 10.6151
R1189 B.n138 B.n137 10.6151
R1190 B.n141 B.n138 10.6151
R1191 B.n142 B.n141 10.6151
R1192 B.n145 B.n142 10.6151
R1193 B.n146 B.n145 10.6151
R1194 B.n149 B.n146 10.6151
R1195 B.n150 B.n149 10.6151
R1196 B.n153 B.n150 10.6151
R1197 B.n154 B.n153 10.6151
R1198 B.n157 B.n154 10.6151
R1199 B.n158 B.n157 10.6151
R1200 B.n161 B.n158 10.6151
R1201 B.n162 B.n161 10.6151
R1202 B.n165 B.n162 10.6151
R1203 B.n166 B.n165 10.6151
R1204 B.n169 B.n166 10.6151
R1205 B.n170 B.n169 10.6151
R1206 B.n173 B.n170 10.6151
R1207 B.n174 B.n173 10.6151
R1208 B.n177 B.n174 10.6151
R1209 B.n182 B.n179 10.6151
R1210 B.n183 B.n182 10.6151
R1211 B.n186 B.n183 10.6151
R1212 B.n187 B.n186 10.6151
R1213 B.n190 B.n187 10.6151
R1214 B.n191 B.n190 10.6151
R1215 B.n194 B.n191 10.6151
R1216 B.n195 B.n194 10.6151
R1217 B.n199 B.n198 10.6151
R1218 B.n202 B.n199 10.6151
R1219 B.n203 B.n202 10.6151
R1220 B.n206 B.n203 10.6151
R1221 B.n207 B.n206 10.6151
R1222 B.n210 B.n207 10.6151
R1223 B.n211 B.n210 10.6151
R1224 B.n214 B.n211 10.6151
R1225 B.n215 B.n214 10.6151
R1226 B.n218 B.n215 10.6151
R1227 B.n219 B.n218 10.6151
R1228 B.n222 B.n219 10.6151
R1229 B.n223 B.n222 10.6151
R1230 B.n226 B.n223 10.6151
R1231 B.n227 B.n226 10.6151
R1232 B.n230 B.n227 10.6151
R1233 B.n231 B.n230 10.6151
R1234 B.n234 B.n231 10.6151
R1235 B.n235 B.n234 10.6151
R1236 B.n238 B.n235 10.6151
R1237 B.n239 B.n238 10.6151
R1238 B.n242 B.n239 10.6151
R1239 B.n243 B.n242 10.6151
R1240 B.n246 B.n243 10.6151
R1241 B.n247 B.n246 10.6151
R1242 B.n250 B.n247 10.6151
R1243 B.n251 B.n250 10.6151
R1244 B.n254 B.n251 10.6151
R1245 B.n255 B.n254 10.6151
R1246 B.n258 B.n255 10.6151
R1247 B.n259 B.n258 10.6151
R1248 B.n262 B.n259 10.6151
R1249 B.n263 B.n262 10.6151
R1250 B.n266 B.n263 10.6151
R1251 B.n267 B.n266 10.6151
R1252 B.n663 B.n267 10.6151
R1253 B.n727 B.n0 8.11757
R1254 B.n727 B.n1 8.11757
R1255 B.n458 B.n368 6.5566
R1256 B.n442 B.n441 6.5566
R1257 B.n179 B.n178 6.5566
R1258 B.n195 B.n101 6.5566
R1259 B.n461 B.n368 4.05904
R1260 B.n441 B.n440 4.05904
R1261 B.n178 B.n177 4.05904
R1262 B.n198 B.n101 4.05904
R1263 B.n559 B.t5 1.41575
R1264 B.n681 B.t9 1.41575
R1265 VP.n10 VP.n0 161.3
R1266 VP.n9 VP.n8 161.3
R1267 VP.n7 VP.n1 161.3
R1268 VP.n6 VP.n5 161.3
R1269 VP.n2 VP.t0 155.004
R1270 VP.n2 VP.t1 154.458
R1271 VP.n4 VP.t2 118.995
R1272 VP.n11 VP.t3 118.995
R1273 VP.n4 VP.n3 88.4915
R1274 VP.n12 VP.n11 88.4915
R1275 VP.n9 VP.n1 56.5193
R1276 VP.n3 VP.n2 50.4085
R1277 VP.n5 VP.n1 24.4675
R1278 VP.n10 VP.n9 24.4675
R1279 VP.n5 VP.n4 22.2655
R1280 VP.n11 VP.n10 22.2655
R1281 VP.n6 VP.n3 0.278367
R1282 VP.n12 VP.n0 0.278367
R1283 VP.n7 VP.n6 0.189894
R1284 VP.n8 VP.n7 0.189894
R1285 VP.n8 VP.n0 0.189894
R1286 VP VP.n12 0.153454
R1287 VDD1 VDD1.n1 100.838
R1288 VDD1 VDD1.n0 61.5713
R1289 VDD1.n0 VDD1.t3 1.92845
R1290 VDD1.n0 VDD1.t2 1.92845
R1291 VDD1.n1 VDD1.t1 1.92845
R1292 VDD1.n1 VDD1.t0 1.92845
C0 VTAIL VP 3.85976f
C1 VDD2 VP 0.361344f
C2 VDD1 VTAIL 4.92488f
C3 VDD1 VDD2 0.903829f
C4 VDD2 VTAIL 4.9756f
C5 VN VP 5.49454f
C6 VDD1 VN 0.148657f
C7 VDD1 VP 4.14203f
C8 VN VTAIL 3.84566f
C9 VN VDD2 3.92995f
C10 VDD2 B 3.33779f
C11 VDD1 B 7.08073f
C12 VTAIL B 8.742281f
C13 VN B 9.577499f
C14 VP B 7.715846f
C15 VDD1.t3 B 0.217466f
C16 VDD1.t2 B 0.217466f
C17 VDD1.n0 B 1.91771f
C18 VDD1.t1 B 0.217466f
C19 VDD1.t0 B 0.217466f
C20 VDD1.n1 B 2.53143f
C21 VP.n0 B 0.039923f
C22 VP.t3 B 1.75394f
C23 VP.n1 B 0.044205f
C24 VP.t1 B 1.93705f
C25 VP.t0 B 1.93983f
C26 VP.n2 B 2.64951f
C27 VP.n3 B 1.58871f
C28 VP.t2 B 1.75394f
C29 VP.n4 B 0.73333f
C30 VP.n5 B 0.053927f
C31 VP.n6 B 0.039923f
C32 VP.n7 B 0.030281f
C33 VP.n8 B 0.030281f
C34 VP.n9 B 0.044205f
C35 VP.n10 B 0.053927f
C36 VP.n11 B 0.73333f
C37 VP.n12 B 0.034755f
C38 VTAIL.t4 B 1.45061f
C39 VTAIL.n0 B 0.303962f
C40 VTAIL.t0 B 1.45061f
C41 VTAIL.n1 B 0.356467f
C42 VTAIL.t1 B 1.45061f
C43 VTAIL.n2 B 1.14232f
C44 VTAIL.t7 B 1.45061f
C45 VTAIL.n3 B 1.14231f
C46 VTAIL.t5 B 1.45061f
C47 VTAIL.n4 B 0.356463f
C48 VTAIL.t3 B 1.45061f
C49 VTAIL.n5 B 0.356463f
C50 VTAIL.t2 B 1.45061f
C51 VTAIL.n6 B 1.14232f
C52 VTAIL.t6 B 1.45061f
C53 VTAIL.n7 B 1.08358f
C54 VDD2.t0 B 0.21744f
C55 VDD2.t3 B 0.21744f
C56 VDD2.n0 B 2.50532f
C57 VDD2.t2 B 0.21744f
C58 VDD2.t1 B 0.21744f
C59 VDD2.n1 B 1.91709f
C60 VDD2.n2 B 3.4227f
C61 VN.t3 B 1.89076f
C62 VN.t1 B 1.88805f
C63 VN.n0 B 1.27371f
C64 VN.t2 B 1.89076f
C65 VN.t0 B 1.88805f
C66 VN.n1 B 2.59766f
.ends

