* NGSPICE file created from diff_pair_sample_1623.ext - technology: sky130A

.subckt diff_pair_sample_1623 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=6.7704 ps=35.5 w=17.36 l=0.63
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=0 ps=0 w=17.36 l=0.63
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=0 ps=0 w=17.36 l=0.63
X3 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=6.7704 ps=35.5 w=17.36 l=0.63
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=0 ps=0 w=17.36 l=0.63
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=6.7704 ps=35.5 w=17.36 l=0.63
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=0 ps=0 w=17.36 l=0.63
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7704 pd=35.5 as=6.7704 ps=35.5 w=17.36 l=0.63
R0 VN VN.t0 931.631
R1 VN VN.t1 887.794
R2 VTAIL.n382 VTAIL.n381 289.615
R3 VTAIL.n94 VTAIL.n93 289.615
R4 VTAIL.n286 VTAIL.n285 289.615
R5 VTAIL.n190 VTAIL.n189 289.615
R6 VTAIL.n318 VTAIL.n317 185
R7 VTAIL.n323 VTAIL.n322 185
R8 VTAIL.n325 VTAIL.n324 185
R9 VTAIL.n314 VTAIL.n313 185
R10 VTAIL.n331 VTAIL.n330 185
R11 VTAIL.n333 VTAIL.n332 185
R12 VTAIL.n310 VTAIL.n309 185
R13 VTAIL.n340 VTAIL.n339 185
R14 VTAIL.n341 VTAIL.n308 185
R15 VTAIL.n343 VTAIL.n342 185
R16 VTAIL.n306 VTAIL.n305 185
R17 VTAIL.n349 VTAIL.n348 185
R18 VTAIL.n351 VTAIL.n350 185
R19 VTAIL.n302 VTAIL.n301 185
R20 VTAIL.n357 VTAIL.n356 185
R21 VTAIL.n359 VTAIL.n358 185
R22 VTAIL.n298 VTAIL.n297 185
R23 VTAIL.n365 VTAIL.n364 185
R24 VTAIL.n367 VTAIL.n366 185
R25 VTAIL.n294 VTAIL.n293 185
R26 VTAIL.n373 VTAIL.n372 185
R27 VTAIL.n375 VTAIL.n374 185
R28 VTAIL.n290 VTAIL.n289 185
R29 VTAIL.n381 VTAIL.n380 185
R30 VTAIL.n30 VTAIL.n29 185
R31 VTAIL.n35 VTAIL.n34 185
R32 VTAIL.n37 VTAIL.n36 185
R33 VTAIL.n26 VTAIL.n25 185
R34 VTAIL.n43 VTAIL.n42 185
R35 VTAIL.n45 VTAIL.n44 185
R36 VTAIL.n22 VTAIL.n21 185
R37 VTAIL.n52 VTAIL.n51 185
R38 VTAIL.n53 VTAIL.n20 185
R39 VTAIL.n55 VTAIL.n54 185
R40 VTAIL.n18 VTAIL.n17 185
R41 VTAIL.n61 VTAIL.n60 185
R42 VTAIL.n63 VTAIL.n62 185
R43 VTAIL.n14 VTAIL.n13 185
R44 VTAIL.n69 VTAIL.n68 185
R45 VTAIL.n71 VTAIL.n70 185
R46 VTAIL.n10 VTAIL.n9 185
R47 VTAIL.n77 VTAIL.n76 185
R48 VTAIL.n79 VTAIL.n78 185
R49 VTAIL.n6 VTAIL.n5 185
R50 VTAIL.n85 VTAIL.n84 185
R51 VTAIL.n87 VTAIL.n86 185
R52 VTAIL.n2 VTAIL.n1 185
R53 VTAIL.n93 VTAIL.n92 185
R54 VTAIL.n285 VTAIL.n284 185
R55 VTAIL.n194 VTAIL.n193 185
R56 VTAIL.n279 VTAIL.n278 185
R57 VTAIL.n277 VTAIL.n276 185
R58 VTAIL.n198 VTAIL.n197 185
R59 VTAIL.n271 VTAIL.n270 185
R60 VTAIL.n269 VTAIL.n268 185
R61 VTAIL.n202 VTAIL.n201 185
R62 VTAIL.n263 VTAIL.n262 185
R63 VTAIL.n261 VTAIL.n260 185
R64 VTAIL.n206 VTAIL.n205 185
R65 VTAIL.n255 VTAIL.n254 185
R66 VTAIL.n253 VTAIL.n252 185
R67 VTAIL.n210 VTAIL.n209 185
R68 VTAIL.n247 VTAIL.n246 185
R69 VTAIL.n245 VTAIL.n212 185
R70 VTAIL.n244 VTAIL.n243 185
R71 VTAIL.n215 VTAIL.n213 185
R72 VTAIL.n238 VTAIL.n237 185
R73 VTAIL.n236 VTAIL.n235 185
R74 VTAIL.n219 VTAIL.n218 185
R75 VTAIL.n230 VTAIL.n229 185
R76 VTAIL.n228 VTAIL.n227 185
R77 VTAIL.n223 VTAIL.n222 185
R78 VTAIL.n189 VTAIL.n188 185
R79 VTAIL.n98 VTAIL.n97 185
R80 VTAIL.n183 VTAIL.n182 185
R81 VTAIL.n181 VTAIL.n180 185
R82 VTAIL.n102 VTAIL.n101 185
R83 VTAIL.n175 VTAIL.n174 185
R84 VTAIL.n173 VTAIL.n172 185
R85 VTAIL.n106 VTAIL.n105 185
R86 VTAIL.n167 VTAIL.n166 185
R87 VTAIL.n165 VTAIL.n164 185
R88 VTAIL.n110 VTAIL.n109 185
R89 VTAIL.n159 VTAIL.n158 185
R90 VTAIL.n157 VTAIL.n156 185
R91 VTAIL.n114 VTAIL.n113 185
R92 VTAIL.n151 VTAIL.n150 185
R93 VTAIL.n149 VTAIL.n116 185
R94 VTAIL.n148 VTAIL.n147 185
R95 VTAIL.n119 VTAIL.n117 185
R96 VTAIL.n142 VTAIL.n141 185
R97 VTAIL.n140 VTAIL.n139 185
R98 VTAIL.n123 VTAIL.n122 185
R99 VTAIL.n134 VTAIL.n133 185
R100 VTAIL.n132 VTAIL.n131 185
R101 VTAIL.n127 VTAIL.n126 185
R102 VTAIL.n319 VTAIL.t3 149.524
R103 VTAIL.n31 VTAIL.t1 149.524
R104 VTAIL.n224 VTAIL.t0 149.524
R105 VTAIL.n128 VTAIL.t2 149.524
R106 VTAIL.n323 VTAIL.n317 104.615
R107 VTAIL.n324 VTAIL.n323 104.615
R108 VTAIL.n324 VTAIL.n313 104.615
R109 VTAIL.n331 VTAIL.n313 104.615
R110 VTAIL.n332 VTAIL.n331 104.615
R111 VTAIL.n332 VTAIL.n309 104.615
R112 VTAIL.n340 VTAIL.n309 104.615
R113 VTAIL.n341 VTAIL.n340 104.615
R114 VTAIL.n342 VTAIL.n341 104.615
R115 VTAIL.n342 VTAIL.n305 104.615
R116 VTAIL.n349 VTAIL.n305 104.615
R117 VTAIL.n350 VTAIL.n349 104.615
R118 VTAIL.n350 VTAIL.n301 104.615
R119 VTAIL.n357 VTAIL.n301 104.615
R120 VTAIL.n358 VTAIL.n357 104.615
R121 VTAIL.n358 VTAIL.n297 104.615
R122 VTAIL.n365 VTAIL.n297 104.615
R123 VTAIL.n366 VTAIL.n365 104.615
R124 VTAIL.n366 VTAIL.n293 104.615
R125 VTAIL.n373 VTAIL.n293 104.615
R126 VTAIL.n374 VTAIL.n373 104.615
R127 VTAIL.n374 VTAIL.n289 104.615
R128 VTAIL.n381 VTAIL.n289 104.615
R129 VTAIL.n35 VTAIL.n29 104.615
R130 VTAIL.n36 VTAIL.n35 104.615
R131 VTAIL.n36 VTAIL.n25 104.615
R132 VTAIL.n43 VTAIL.n25 104.615
R133 VTAIL.n44 VTAIL.n43 104.615
R134 VTAIL.n44 VTAIL.n21 104.615
R135 VTAIL.n52 VTAIL.n21 104.615
R136 VTAIL.n53 VTAIL.n52 104.615
R137 VTAIL.n54 VTAIL.n53 104.615
R138 VTAIL.n54 VTAIL.n17 104.615
R139 VTAIL.n61 VTAIL.n17 104.615
R140 VTAIL.n62 VTAIL.n61 104.615
R141 VTAIL.n62 VTAIL.n13 104.615
R142 VTAIL.n69 VTAIL.n13 104.615
R143 VTAIL.n70 VTAIL.n69 104.615
R144 VTAIL.n70 VTAIL.n9 104.615
R145 VTAIL.n77 VTAIL.n9 104.615
R146 VTAIL.n78 VTAIL.n77 104.615
R147 VTAIL.n78 VTAIL.n5 104.615
R148 VTAIL.n85 VTAIL.n5 104.615
R149 VTAIL.n86 VTAIL.n85 104.615
R150 VTAIL.n86 VTAIL.n1 104.615
R151 VTAIL.n93 VTAIL.n1 104.615
R152 VTAIL.n285 VTAIL.n193 104.615
R153 VTAIL.n278 VTAIL.n193 104.615
R154 VTAIL.n278 VTAIL.n277 104.615
R155 VTAIL.n277 VTAIL.n197 104.615
R156 VTAIL.n270 VTAIL.n197 104.615
R157 VTAIL.n270 VTAIL.n269 104.615
R158 VTAIL.n269 VTAIL.n201 104.615
R159 VTAIL.n262 VTAIL.n201 104.615
R160 VTAIL.n262 VTAIL.n261 104.615
R161 VTAIL.n261 VTAIL.n205 104.615
R162 VTAIL.n254 VTAIL.n205 104.615
R163 VTAIL.n254 VTAIL.n253 104.615
R164 VTAIL.n253 VTAIL.n209 104.615
R165 VTAIL.n246 VTAIL.n209 104.615
R166 VTAIL.n246 VTAIL.n245 104.615
R167 VTAIL.n245 VTAIL.n244 104.615
R168 VTAIL.n244 VTAIL.n213 104.615
R169 VTAIL.n237 VTAIL.n213 104.615
R170 VTAIL.n237 VTAIL.n236 104.615
R171 VTAIL.n236 VTAIL.n218 104.615
R172 VTAIL.n229 VTAIL.n218 104.615
R173 VTAIL.n229 VTAIL.n228 104.615
R174 VTAIL.n228 VTAIL.n222 104.615
R175 VTAIL.n189 VTAIL.n97 104.615
R176 VTAIL.n182 VTAIL.n97 104.615
R177 VTAIL.n182 VTAIL.n181 104.615
R178 VTAIL.n181 VTAIL.n101 104.615
R179 VTAIL.n174 VTAIL.n101 104.615
R180 VTAIL.n174 VTAIL.n173 104.615
R181 VTAIL.n173 VTAIL.n105 104.615
R182 VTAIL.n166 VTAIL.n105 104.615
R183 VTAIL.n166 VTAIL.n165 104.615
R184 VTAIL.n165 VTAIL.n109 104.615
R185 VTAIL.n158 VTAIL.n109 104.615
R186 VTAIL.n158 VTAIL.n157 104.615
R187 VTAIL.n157 VTAIL.n113 104.615
R188 VTAIL.n150 VTAIL.n113 104.615
R189 VTAIL.n150 VTAIL.n149 104.615
R190 VTAIL.n149 VTAIL.n148 104.615
R191 VTAIL.n148 VTAIL.n117 104.615
R192 VTAIL.n141 VTAIL.n117 104.615
R193 VTAIL.n141 VTAIL.n140 104.615
R194 VTAIL.n140 VTAIL.n122 104.615
R195 VTAIL.n133 VTAIL.n122 104.615
R196 VTAIL.n133 VTAIL.n132 104.615
R197 VTAIL.n132 VTAIL.n126 104.615
R198 VTAIL.t3 VTAIL.n317 52.3082
R199 VTAIL.t1 VTAIL.n29 52.3082
R200 VTAIL.t0 VTAIL.n222 52.3082
R201 VTAIL.t2 VTAIL.n126 52.3082
R202 VTAIL.n383 VTAIL.n382 34.1247
R203 VTAIL.n95 VTAIL.n94 34.1247
R204 VTAIL.n287 VTAIL.n286 34.1247
R205 VTAIL.n191 VTAIL.n190 34.1247
R206 VTAIL.n191 VTAIL.n95 29.0048
R207 VTAIL.n383 VTAIL.n287 28.1772
R208 VTAIL.n343 VTAIL.n308 13.1884
R209 VTAIL.n55 VTAIL.n20 13.1884
R210 VTAIL.n247 VTAIL.n212 13.1884
R211 VTAIL.n151 VTAIL.n116 13.1884
R212 VTAIL.n339 VTAIL.n338 12.8005
R213 VTAIL.n344 VTAIL.n306 12.8005
R214 VTAIL.n51 VTAIL.n50 12.8005
R215 VTAIL.n56 VTAIL.n18 12.8005
R216 VTAIL.n248 VTAIL.n210 12.8005
R217 VTAIL.n243 VTAIL.n214 12.8005
R218 VTAIL.n152 VTAIL.n114 12.8005
R219 VTAIL.n147 VTAIL.n118 12.8005
R220 VTAIL.n337 VTAIL.n310 12.0247
R221 VTAIL.n348 VTAIL.n347 12.0247
R222 VTAIL.n49 VTAIL.n22 12.0247
R223 VTAIL.n60 VTAIL.n59 12.0247
R224 VTAIL.n252 VTAIL.n251 12.0247
R225 VTAIL.n242 VTAIL.n215 12.0247
R226 VTAIL.n156 VTAIL.n155 12.0247
R227 VTAIL.n146 VTAIL.n119 12.0247
R228 VTAIL.n334 VTAIL.n333 11.249
R229 VTAIL.n351 VTAIL.n304 11.249
R230 VTAIL.n380 VTAIL.n288 11.249
R231 VTAIL.n46 VTAIL.n45 11.249
R232 VTAIL.n63 VTAIL.n16 11.249
R233 VTAIL.n92 VTAIL.n0 11.249
R234 VTAIL.n284 VTAIL.n192 11.249
R235 VTAIL.n255 VTAIL.n208 11.249
R236 VTAIL.n239 VTAIL.n238 11.249
R237 VTAIL.n188 VTAIL.n96 11.249
R238 VTAIL.n159 VTAIL.n112 11.249
R239 VTAIL.n143 VTAIL.n142 11.249
R240 VTAIL.n330 VTAIL.n312 10.4732
R241 VTAIL.n352 VTAIL.n302 10.4732
R242 VTAIL.n379 VTAIL.n290 10.4732
R243 VTAIL.n42 VTAIL.n24 10.4732
R244 VTAIL.n64 VTAIL.n14 10.4732
R245 VTAIL.n91 VTAIL.n2 10.4732
R246 VTAIL.n283 VTAIL.n194 10.4732
R247 VTAIL.n256 VTAIL.n206 10.4732
R248 VTAIL.n235 VTAIL.n217 10.4732
R249 VTAIL.n187 VTAIL.n98 10.4732
R250 VTAIL.n160 VTAIL.n110 10.4732
R251 VTAIL.n139 VTAIL.n121 10.4732
R252 VTAIL.n319 VTAIL.n318 10.2747
R253 VTAIL.n31 VTAIL.n30 10.2747
R254 VTAIL.n224 VTAIL.n223 10.2747
R255 VTAIL.n128 VTAIL.n127 10.2747
R256 VTAIL.n329 VTAIL.n314 9.69747
R257 VTAIL.n356 VTAIL.n355 9.69747
R258 VTAIL.n376 VTAIL.n375 9.69747
R259 VTAIL.n41 VTAIL.n26 9.69747
R260 VTAIL.n68 VTAIL.n67 9.69747
R261 VTAIL.n88 VTAIL.n87 9.69747
R262 VTAIL.n280 VTAIL.n279 9.69747
R263 VTAIL.n260 VTAIL.n259 9.69747
R264 VTAIL.n234 VTAIL.n219 9.69747
R265 VTAIL.n184 VTAIL.n183 9.69747
R266 VTAIL.n164 VTAIL.n163 9.69747
R267 VTAIL.n138 VTAIL.n123 9.69747
R268 VTAIL.n378 VTAIL.n288 9.45567
R269 VTAIL.n90 VTAIL.n0 9.45567
R270 VTAIL.n282 VTAIL.n192 9.45567
R271 VTAIL.n186 VTAIL.n96 9.45567
R272 VTAIL.n296 VTAIL.n295 9.3005
R273 VTAIL.n369 VTAIL.n368 9.3005
R274 VTAIL.n371 VTAIL.n370 9.3005
R275 VTAIL.n292 VTAIL.n291 9.3005
R276 VTAIL.n377 VTAIL.n376 9.3005
R277 VTAIL.n379 VTAIL.n378 9.3005
R278 VTAIL.n361 VTAIL.n360 9.3005
R279 VTAIL.n300 VTAIL.n299 9.3005
R280 VTAIL.n355 VTAIL.n354 9.3005
R281 VTAIL.n353 VTAIL.n352 9.3005
R282 VTAIL.n304 VTAIL.n303 9.3005
R283 VTAIL.n347 VTAIL.n346 9.3005
R284 VTAIL.n345 VTAIL.n344 9.3005
R285 VTAIL.n321 VTAIL.n320 9.3005
R286 VTAIL.n316 VTAIL.n315 9.3005
R287 VTAIL.n327 VTAIL.n326 9.3005
R288 VTAIL.n329 VTAIL.n328 9.3005
R289 VTAIL.n312 VTAIL.n311 9.3005
R290 VTAIL.n335 VTAIL.n334 9.3005
R291 VTAIL.n337 VTAIL.n336 9.3005
R292 VTAIL.n338 VTAIL.n307 9.3005
R293 VTAIL.n363 VTAIL.n362 9.3005
R294 VTAIL.n8 VTAIL.n7 9.3005
R295 VTAIL.n81 VTAIL.n80 9.3005
R296 VTAIL.n83 VTAIL.n82 9.3005
R297 VTAIL.n4 VTAIL.n3 9.3005
R298 VTAIL.n89 VTAIL.n88 9.3005
R299 VTAIL.n91 VTAIL.n90 9.3005
R300 VTAIL.n73 VTAIL.n72 9.3005
R301 VTAIL.n12 VTAIL.n11 9.3005
R302 VTAIL.n67 VTAIL.n66 9.3005
R303 VTAIL.n65 VTAIL.n64 9.3005
R304 VTAIL.n16 VTAIL.n15 9.3005
R305 VTAIL.n59 VTAIL.n58 9.3005
R306 VTAIL.n57 VTAIL.n56 9.3005
R307 VTAIL.n33 VTAIL.n32 9.3005
R308 VTAIL.n28 VTAIL.n27 9.3005
R309 VTAIL.n39 VTAIL.n38 9.3005
R310 VTAIL.n41 VTAIL.n40 9.3005
R311 VTAIL.n24 VTAIL.n23 9.3005
R312 VTAIL.n47 VTAIL.n46 9.3005
R313 VTAIL.n49 VTAIL.n48 9.3005
R314 VTAIL.n50 VTAIL.n19 9.3005
R315 VTAIL.n75 VTAIL.n74 9.3005
R316 VTAIL.n283 VTAIL.n282 9.3005
R317 VTAIL.n281 VTAIL.n280 9.3005
R318 VTAIL.n196 VTAIL.n195 9.3005
R319 VTAIL.n275 VTAIL.n274 9.3005
R320 VTAIL.n273 VTAIL.n272 9.3005
R321 VTAIL.n200 VTAIL.n199 9.3005
R322 VTAIL.n267 VTAIL.n266 9.3005
R323 VTAIL.n265 VTAIL.n264 9.3005
R324 VTAIL.n204 VTAIL.n203 9.3005
R325 VTAIL.n259 VTAIL.n258 9.3005
R326 VTAIL.n257 VTAIL.n256 9.3005
R327 VTAIL.n208 VTAIL.n207 9.3005
R328 VTAIL.n251 VTAIL.n250 9.3005
R329 VTAIL.n249 VTAIL.n248 9.3005
R330 VTAIL.n214 VTAIL.n211 9.3005
R331 VTAIL.n242 VTAIL.n241 9.3005
R332 VTAIL.n240 VTAIL.n239 9.3005
R333 VTAIL.n217 VTAIL.n216 9.3005
R334 VTAIL.n234 VTAIL.n233 9.3005
R335 VTAIL.n232 VTAIL.n231 9.3005
R336 VTAIL.n221 VTAIL.n220 9.3005
R337 VTAIL.n226 VTAIL.n225 9.3005
R338 VTAIL.n130 VTAIL.n129 9.3005
R339 VTAIL.n125 VTAIL.n124 9.3005
R340 VTAIL.n136 VTAIL.n135 9.3005
R341 VTAIL.n138 VTAIL.n137 9.3005
R342 VTAIL.n121 VTAIL.n120 9.3005
R343 VTAIL.n144 VTAIL.n143 9.3005
R344 VTAIL.n146 VTAIL.n145 9.3005
R345 VTAIL.n118 VTAIL.n115 9.3005
R346 VTAIL.n177 VTAIL.n176 9.3005
R347 VTAIL.n179 VTAIL.n178 9.3005
R348 VTAIL.n100 VTAIL.n99 9.3005
R349 VTAIL.n185 VTAIL.n184 9.3005
R350 VTAIL.n187 VTAIL.n186 9.3005
R351 VTAIL.n104 VTAIL.n103 9.3005
R352 VTAIL.n171 VTAIL.n170 9.3005
R353 VTAIL.n169 VTAIL.n168 9.3005
R354 VTAIL.n108 VTAIL.n107 9.3005
R355 VTAIL.n163 VTAIL.n162 9.3005
R356 VTAIL.n161 VTAIL.n160 9.3005
R357 VTAIL.n112 VTAIL.n111 9.3005
R358 VTAIL.n155 VTAIL.n154 9.3005
R359 VTAIL.n153 VTAIL.n152 9.3005
R360 VTAIL.n326 VTAIL.n325 8.92171
R361 VTAIL.n359 VTAIL.n300 8.92171
R362 VTAIL.n372 VTAIL.n292 8.92171
R363 VTAIL.n38 VTAIL.n37 8.92171
R364 VTAIL.n71 VTAIL.n12 8.92171
R365 VTAIL.n84 VTAIL.n4 8.92171
R366 VTAIL.n276 VTAIL.n196 8.92171
R367 VTAIL.n263 VTAIL.n204 8.92171
R368 VTAIL.n231 VTAIL.n230 8.92171
R369 VTAIL.n180 VTAIL.n100 8.92171
R370 VTAIL.n167 VTAIL.n108 8.92171
R371 VTAIL.n135 VTAIL.n134 8.92171
R372 VTAIL.n322 VTAIL.n316 8.14595
R373 VTAIL.n360 VTAIL.n298 8.14595
R374 VTAIL.n371 VTAIL.n294 8.14595
R375 VTAIL.n34 VTAIL.n28 8.14595
R376 VTAIL.n72 VTAIL.n10 8.14595
R377 VTAIL.n83 VTAIL.n6 8.14595
R378 VTAIL.n275 VTAIL.n198 8.14595
R379 VTAIL.n264 VTAIL.n202 8.14595
R380 VTAIL.n227 VTAIL.n221 8.14595
R381 VTAIL.n179 VTAIL.n102 8.14595
R382 VTAIL.n168 VTAIL.n106 8.14595
R383 VTAIL.n131 VTAIL.n125 8.14595
R384 VTAIL.n321 VTAIL.n318 7.3702
R385 VTAIL.n364 VTAIL.n363 7.3702
R386 VTAIL.n368 VTAIL.n367 7.3702
R387 VTAIL.n33 VTAIL.n30 7.3702
R388 VTAIL.n76 VTAIL.n75 7.3702
R389 VTAIL.n80 VTAIL.n79 7.3702
R390 VTAIL.n272 VTAIL.n271 7.3702
R391 VTAIL.n268 VTAIL.n267 7.3702
R392 VTAIL.n226 VTAIL.n223 7.3702
R393 VTAIL.n176 VTAIL.n175 7.3702
R394 VTAIL.n172 VTAIL.n171 7.3702
R395 VTAIL.n130 VTAIL.n127 7.3702
R396 VTAIL.n364 VTAIL.n296 6.59444
R397 VTAIL.n367 VTAIL.n296 6.59444
R398 VTAIL.n76 VTAIL.n8 6.59444
R399 VTAIL.n79 VTAIL.n8 6.59444
R400 VTAIL.n271 VTAIL.n200 6.59444
R401 VTAIL.n268 VTAIL.n200 6.59444
R402 VTAIL.n175 VTAIL.n104 6.59444
R403 VTAIL.n172 VTAIL.n104 6.59444
R404 VTAIL.n322 VTAIL.n321 5.81868
R405 VTAIL.n363 VTAIL.n298 5.81868
R406 VTAIL.n368 VTAIL.n294 5.81868
R407 VTAIL.n34 VTAIL.n33 5.81868
R408 VTAIL.n75 VTAIL.n10 5.81868
R409 VTAIL.n80 VTAIL.n6 5.81868
R410 VTAIL.n272 VTAIL.n198 5.81868
R411 VTAIL.n267 VTAIL.n202 5.81868
R412 VTAIL.n227 VTAIL.n226 5.81868
R413 VTAIL.n176 VTAIL.n102 5.81868
R414 VTAIL.n171 VTAIL.n106 5.81868
R415 VTAIL.n131 VTAIL.n130 5.81868
R416 VTAIL.n325 VTAIL.n316 5.04292
R417 VTAIL.n360 VTAIL.n359 5.04292
R418 VTAIL.n372 VTAIL.n371 5.04292
R419 VTAIL.n37 VTAIL.n28 5.04292
R420 VTAIL.n72 VTAIL.n71 5.04292
R421 VTAIL.n84 VTAIL.n83 5.04292
R422 VTAIL.n276 VTAIL.n275 5.04292
R423 VTAIL.n264 VTAIL.n263 5.04292
R424 VTAIL.n230 VTAIL.n221 5.04292
R425 VTAIL.n180 VTAIL.n179 5.04292
R426 VTAIL.n168 VTAIL.n167 5.04292
R427 VTAIL.n134 VTAIL.n125 5.04292
R428 VTAIL.n326 VTAIL.n314 4.26717
R429 VTAIL.n356 VTAIL.n300 4.26717
R430 VTAIL.n375 VTAIL.n292 4.26717
R431 VTAIL.n38 VTAIL.n26 4.26717
R432 VTAIL.n68 VTAIL.n12 4.26717
R433 VTAIL.n87 VTAIL.n4 4.26717
R434 VTAIL.n279 VTAIL.n196 4.26717
R435 VTAIL.n260 VTAIL.n204 4.26717
R436 VTAIL.n231 VTAIL.n219 4.26717
R437 VTAIL.n183 VTAIL.n100 4.26717
R438 VTAIL.n164 VTAIL.n108 4.26717
R439 VTAIL.n135 VTAIL.n123 4.26717
R440 VTAIL.n330 VTAIL.n329 3.49141
R441 VTAIL.n355 VTAIL.n302 3.49141
R442 VTAIL.n376 VTAIL.n290 3.49141
R443 VTAIL.n42 VTAIL.n41 3.49141
R444 VTAIL.n67 VTAIL.n14 3.49141
R445 VTAIL.n88 VTAIL.n2 3.49141
R446 VTAIL.n280 VTAIL.n194 3.49141
R447 VTAIL.n259 VTAIL.n206 3.49141
R448 VTAIL.n235 VTAIL.n234 3.49141
R449 VTAIL.n184 VTAIL.n98 3.49141
R450 VTAIL.n163 VTAIL.n110 3.49141
R451 VTAIL.n139 VTAIL.n138 3.49141
R452 VTAIL.n320 VTAIL.n319 2.84303
R453 VTAIL.n32 VTAIL.n31 2.84303
R454 VTAIL.n225 VTAIL.n224 2.84303
R455 VTAIL.n129 VTAIL.n128 2.84303
R456 VTAIL.n333 VTAIL.n312 2.71565
R457 VTAIL.n352 VTAIL.n351 2.71565
R458 VTAIL.n380 VTAIL.n379 2.71565
R459 VTAIL.n45 VTAIL.n24 2.71565
R460 VTAIL.n64 VTAIL.n63 2.71565
R461 VTAIL.n92 VTAIL.n91 2.71565
R462 VTAIL.n284 VTAIL.n283 2.71565
R463 VTAIL.n256 VTAIL.n255 2.71565
R464 VTAIL.n238 VTAIL.n217 2.71565
R465 VTAIL.n188 VTAIL.n187 2.71565
R466 VTAIL.n160 VTAIL.n159 2.71565
R467 VTAIL.n142 VTAIL.n121 2.71565
R468 VTAIL.n334 VTAIL.n310 1.93989
R469 VTAIL.n348 VTAIL.n304 1.93989
R470 VTAIL.n382 VTAIL.n288 1.93989
R471 VTAIL.n46 VTAIL.n22 1.93989
R472 VTAIL.n60 VTAIL.n16 1.93989
R473 VTAIL.n94 VTAIL.n0 1.93989
R474 VTAIL.n286 VTAIL.n192 1.93989
R475 VTAIL.n252 VTAIL.n208 1.93989
R476 VTAIL.n239 VTAIL.n215 1.93989
R477 VTAIL.n190 VTAIL.n96 1.93989
R478 VTAIL.n156 VTAIL.n112 1.93989
R479 VTAIL.n143 VTAIL.n119 1.93989
R480 VTAIL.n339 VTAIL.n337 1.16414
R481 VTAIL.n347 VTAIL.n306 1.16414
R482 VTAIL.n51 VTAIL.n49 1.16414
R483 VTAIL.n59 VTAIL.n18 1.16414
R484 VTAIL.n251 VTAIL.n210 1.16414
R485 VTAIL.n243 VTAIL.n242 1.16414
R486 VTAIL.n155 VTAIL.n114 1.16414
R487 VTAIL.n147 VTAIL.n146 1.16414
R488 VTAIL.n287 VTAIL.n191 0.884121
R489 VTAIL VTAIL.n95 0.735414
R490 VTAIL.n338 VTAIL.n308 0.388379
R491 VTAIL.n344 VTAIL.n343 0.388379
R492 VTAIL.n50 VTAIL.n20 0.388379
R493 VTAIL.n56 VTAIL.n55 0.388379
R494 VTAIL.n248 VTAIL.n247 0.388379
R495 VTAIL.n214 VTAIL.n212 0.388379
R496 VTAIL.n152 VTAIL.n151 0.388379
R497 VTAIL.n118 VTAIL.n116 0.388379
R498 VTAIL.n320 VTAIL.n315 0.155672
R499 VTAIL.n327 VTAIL.n315 0.155672
R500 VTAIL.n328 VTAIL.n327 0.155672
R501 VTAIL.n328 VTAIL.n311 0.155672
R502 VTAIL.n335 VTAIL.n311 0.155672
R503 VTAIL.n336 VTAIL.n335 0.155672
R504 VTAIL.n336 VTAIL.n307 0.155672
R505 VTAIL.n345 VTAIL.n307 0.155672
R506 VTAIL.n346 VTAIL.n345 0.155672
R507 VTAIL.n346 VTAIL.n303 0.155672
R508 VTAIL.n353 VTAIL.n303 0.155672
R509 VTAIL.n354 VTAIL.n353 0.155672
R510 VTAIL.n354 VTAIL.n299 0.155672
R511 VTAIL.n361 VTAIL.n299 0.155672
R512 VTAIL.n362 VTAIL.n361 0.155672
R513 VTAIL.n362 VTAIL.n295 0.155672
R514 VTAIL.n369 VTAIL.n295 0.155672
R515 VTAIL.n370 VTAIL.n369 0.155672
R516 VTAIL.n370 VTAIL.n291 0.155672
R517 VTAIL.n377 VTAIL.n291 0.155672
R518 VTAIL.n378 VTAIL.n377 0.155672
R519 VTAIL.n32 VTAIL.n27 0.155672
R520 VTAIL.n39 VTAIL.n27 0.155672
R521 VTAIL.n40 VTAIL.n39 0.155672
R522 VTAIL.n40 VTAIL.n23 0.155672
R523 VTAIL.n47 VTAIL.n23 0.155672
R524 VTAIL.n48 VTAIL.n47 0.155672
R525 VTAIL.n48 VTAIL.n19 0.155672
R526 VTAIL.n57 VTAIL.n19 0.155672
R527 VTAIL.n58 VTAIL.n57 0.155672
R528 VTAIL.n58 VTAIL.n15 0.155672
R529 VTAIL.n65 VTAIL.n15 0.155672
R530 VTAIL.n66 VTAIL.n65 0.155672
R531 VTAIL.n66 VTAIL.n11 0.155672
R532 VTAIL.n73 VTAIL.n11 0.155672
R533 VTAIL.n74 VTAIL.n73 0.155672
R534 VTAIL.n74 VTAIL.n7 0.155672
R535 VTAIL.n81 VTAIL.n7 0.155672
R536 VTAIL.n82 VTAIL.n81 0.155672
R537 VTAIL.n82 VTAIL.n3 0.155672
R538 VTAIL.n89 VTAIL.n3 0.155672
R539 VTAIL.n90 VTAIL.n89 0.155672
R540 VTAIL.n282 VTAIL.n281 0.155672
R541 VTAIL.n281 VTAIL.n195 0.155672
R542 VTAIL.n274 VTAIL.n195 0.155672
R543 VTAIL.n274 VTAIL.n273 0.155672
R544 VTAIL.n273 VTAIL.n199 0.155672
R545 VTAIL.n266 VTAIL.n199 0.155672
R546 VTAIL.n266 VTAIL.n265 0.155672
R547 VTAIL.n265 VTAIL.n203 0.155672
R548 VTAIL.n258 VTAIL.n203 0.155672
R549 VTAIL.n258 VTAIL.n257 0.155672
R550 VTAIL.n257 VTAIL.n207 0.155672
R551 VTAIL.n250 VTAIL.n207 0.155672
R552 VTAIL.n250 VTAIL.n249 0.155672
R553 VTAIL.n249 VTAIL.n211 0.155672
R554 VTAIL.n241 VTAIL.n211 0.155672
R555 VTAIL.n241 VTAIL.n240 0.155672
R556 VTAIL.n240 VTAIL.n216 0.155672
R557 VTAIL.n233 VTAIL.n216 0.155672
R558 VTAIL.n233 VTAIL.n232 0.155672
R559 VTAIL.n232 VTAIL.n220 0.155672
R560 VTAIL.n225 VTAIL.n220 0.155672
R561 VTAIL.n186 VTAIL.n185 0.155672
R562 VTAIL.n185 VTAIL.n99 0.155672
R563 VTAIL.n178 VTAIL.n99 0.155672
R564 VTAIL.n178 VTAIL.n177 0.155672
R565 VTAIL.n177 VTAIL.n103 0.155672
R566 VTAIL.n170 VTAIL.n103 0.155672
R567 VTAIL.n170 VTAIL.n169 0.155672
R568 VTAIL.n169 VTAIL.n107 0.155672
R569 VTAIL.n162 VTAIL.n107 0.155672
R570 VTAIL.n162 VTAIL.n161 0.155672
R571 VTAIL.n161 VTAIL.n111 0.155672
R572 VTAIL.n154 VTAIL.n111 0.155672
R573 VTAIL.n154 VTAIL.n153 0.155672
R574 VTAIL.n153 VTAIL.n115 0.155672
R575 VTAIL.n145 VTAIL.n115 0.155672
R576 VTAIL.n145 VTAIL.n144 0.155672
R577 VTAIL.n144 VTAIL.n120 0.155672
R578 VTAIL.n137 VTAIL.n120 0.155672
R579 VTAIL.n137 VTAIL.n136 0.155672
R580 VTAIL.n136 VTAIL.n124 0.155672
R581 VTAIL.n129 VTAIL.n124 0.155672
R582 VTAIL VTAIL.n383 0.149207
R583 VDD2.n189 VDD2.n188 289.615
R584 VDD2.n94 VDD2.n93 289.615
R585 VDD2.n188 VDD2.n187 185
R586 VDD2.n97 VDD2.n96 185
R587 VDD2.n182 VDD2.n181 185
R588 VDD2.n180 VDD2.n179 185
R589 VDD2.n101 VDD2.n100 185
R590 VDD2.n174 VDD2.n173 185
R591 VDD2.n172 VDD2.n171 185
R592 VDD2.n105 VDD2.n104 185
R593 VDD2.n166 VDD2.n165 185
R594 VDD2.n164 VDD2.n163 185
R595 VDD2.n109 VDD2.n108 185
R596 VDD2.n158 VDD2.n157 185
R597 VDD2.n156 VDD2.n155 185
R598 VDD2.n113 VDD2.n112 185
R599 VDD2.n150 VDD2.n149 185
R600 VDD2.n148 VDD2.n115 185
R601 VDD2.n147 VDD2.n146 185
R602 VDD2.n118 VDD2.n116 185
R603 VDD2.n141 VDD2.n140 185
R604 VDD2.n139 VDD2.n138 185
R605 VDD2.n122 VDD2.n121 185
R606 VDD2.n133 VDD2.n132 185
R607 VDD2.n131 VDD2.n130 185
R608 VDD2.n126 VDD2.n125 185
R609 VDD2.n30 VDD2.n29 185
R610 VDD2.n35 VDD2.n34 185
R611 VDD2.n37 VDD2.n36 185
R612 VDD2.n26 VDD2.n25 185
R613 VDD2.n43 VDD2.n42 185
R614 VDD2.n45 VDD2.n44 185
R615 VDD2.n22 VDD2.n21 185
R616 VDD2.n52 VDD2.n51 185
R617 VDD2.n53 VDD2.n20 185
R618 VDD2.n55 VDD2.n54 185
R619 VDD2.n18 VDD2.n17 185
R620 VDD2.n61 VDD2.n60 185
R621 VDD2.n63 VDD2.n62 185
R622 VDD2.n14 VDD2.n13 185
R623 VDD2.n69 VDD2.n68 185
R624 VDD2.n71 VDD2.n70 185
R625 VDD2.n10 VDD2.n9 185
R626 VDD2.n77 VDD2.n76 185
R627 VDD2.n79 VDD2.n78 185
R628 VDD2.n6 VDD2.n5 185
R629 VDD2.n85 VDD2.n84 185
R630 VDD2.n87 VDD2.n86 185
R631 VDD2.n2 VDD2.n1 185
R632 VDD2.n93 VDD2.n92 185
R633 VDD2.n127 VDD2.t1 149.524
R634 VDD2.n31 VDD2.t0 149.524
R635 VDD2.n188 VDD2.n96 104.615
R636 VDD2.n181 VDD2.n96 104.615
R637 VDD2.n181 VDD2.n180 104.615
R638 VDD2.n180 VDD2.n100 104.615
R639 VDD2.n173 VDD2.n100 104.615
R640 VDD2.n173 VDD2.n172 104.615
R641 VDD2.n172 VDD2.n104 104.615
R642 VDD2.n165 VDD2.n104 104.615
R643 VDD2.n165 VDD2.n164 104.615
R644 VDD2.n164 VDD2.n108 104.615
R645 VDD2.n157 VDD2.n108 104.615
R646 VDD2.n157 VDD2.n156 104.615
R647 VDD2.n156 VDD2.n112 104.615
R648 VDD2.n149 VDD2.n112 104.615
R649 VDD2.n149 VDD2.n148 104.615
R650 VDD2.n148 VDD2.n147 104.615
R651 VDD2.n147 VDD2.n116 104.615
R652 VDD2.n140 VDD2.n116 104.615
R653 VDD2.n140 VDD2.n139 104.615
R654 VDD2.n139 VDD2.n121 104.615
R655 VDD2.n132 VDD2.n121 104.615
R656 VDD2.n132 VDD2.n131 104.615
R657 VDD2.n131 VDD2.n125 104.615
R658 VDD2.n35 VDD2.n29 104.615
R659 VDD2.n36 VDD2.n35 104.615
R660 VDD2.n36 VDD2.n25 104.615
R661 VDD2.n43 VDD2.n25 104.615
R662 VDD2.n44 VDD2.n43 104.615
R663 VDD2.n44 VDD2.n21 104.615
R664 VDD2.n52 VDD2.n21 104.615
R665 VDD2.n53 VDD2.n52 104.615
R666 VDD2.n54 VDD2.n53 104.615
R667 VDD2.n54 VDD2.n17 104.615
R668 VDD2.n61 VDD2.n17 104.615
R669 VDD2.n62 VDD2.n61 104.615
R670 VDD2.n62 VDD2.n13 104.615
R671 VDD2.n69 VDD2.n13 104.615
R672 VDD2.n70 VDD2.n69 104.615
R673 VDD2.n70 VDD2.n9 104.615
R674 VDD2.n77 VDD2.n9 104.615
R675 VDD2.n78 VDD2.n77 104.615
R676 VDD2.n78 VDD2.n5 104.615
R677 VDD2.n85 VDD2.n5 104.615
R678 VDD2.n86 VDD2.n85 104.615
R679 VDD2.n86 VDD2.n1 104.615
R680 VDD2.n93 VDD2.n1 104.615
R681 VDD2.n190 VDD2.n94 91.1009
R682 VDD2.t1 VDD2.n125 52.3082
R683 VDD2.t0 VDD2.n29 52.3082
R684 VDD2.n190 VDD2.n189 50.8035
R685 VDD2.n150 VDD2.n115 13.1884
R686 VDD2.n55 VDD2.n20 13.1884
R687 VDD2.n151 VDD2.n113 12.8005
R688 VDD2.n146 VDD2.n117 12.8005
R689 VDD2.n51 VDD2.n50 12.8005
R690 VDD2.n56 VDD2.n18 12.8005
R691 VDD2.n155 VDD2.n154 12.0247
R692 VDD2.n145 VDD2.n118 12.0247
R693 VDD2.n49 VDD2.n22 12.0247
R694 VDD2.n60 VDD2.n59 12.0247
R695 VDD2.n187 VDD2.n95 11.249
R696 VDD2.n158 VDD2.n111 11.249
R697 VDD2.n142 VDD2.n141 11.249
R698 VDD2.n46 VDD2.n45 11.249
R699 VDD2.n63 VDD2.n16 11.249
R700 VDD2.n92 VDD2.n0 11.249
R701 VDD2.n186 VDD2.n97 10.4732
R702 VDD2.n159 VDD2.n109 10.4732
R703 VDD2.n138 VDD2.n120 10.4732
R704 VDD2.n42 VDD2.n24 10.4732
R705 VDD2.n64 VDD2.n14 10.4732
R706 VDD2.n91 VDD2.n2 10.4732
R707 VDD2.n127 VDD2.n126 10.2747
R708 VDD2.n31 VDD2.n30 10.2747
R709 VDD2.n183 VDD2.n182 9.69747
R710 VDD2.n163 VDD2.n162 9.69747
R711 VDD2.n137 VDD2.n122 9.69747
R712 VDD2.n41 VDD2.n26 9.69747
R713 VDD2.n68 VDD2.n67 9.69747
R714 VDD2.n88 VDD2.n87 9.69747
R715 VDD2.n185 VDD2.n95 9.45567
R716 VDD2.n90 VDD2.n0 9.45567
R717 VDD2.n186 VDD2.n185 9.3005
R718 VDD2.n184 VDD2.n183 9.3005
R719 VDD2.n99 VDD2.n98 9.3005
R720 VDD2.n178 VDD2.n177 9.3005
R721 VDD2.n176 VDD2.n175 9.3005
R722 VDD2.n103 VDD2.n102 9.3005
R723 VDD2.n170 VDD2.n169 9.3005
R724 VDD2.n168 VDD2.n167 9.3005
R725 VDD2.n107 VDD2.n106 9.3005
R726 VDD2.n162 VDD2.n161 9.3005
R727 VDD2.n160 VDD2.n159 9.3005
R728 VDD2.n111 VDD2.n110 9.3005
R729 VDD2.n154 VDD2.n153 9.3005
R730 VDD2.n152 VDD2.n151 9.3005
R731 VDD2.n117 VDD2.n114 9.3005
R732 VDD2.n145 VDD2.n144 9.3005
R733 VDD2.n143 VDD2.n142 9.3005
R734 VDD2.n120 VDD2.n119 9.3005
R735 VDD2.n137 VDD2.n136 9.3005
R736 VDD2.n135 VDD2.n134 9.3005
R737 VDD2.n124 VDD2.n123 9.3005
R738 VDD2.n129 VDD2.n128 9.3005
R739 VDD2.n8 VDD2.n7 9.3005
R740 VDD2.n81 VDD2.n80 9.3005
R741 VDD2.n83 VDD2.n82 9.3005
R742 VDD2.n4 VDD2.n3 9.3005
R743 VDD2.n89 VDD2.n88 9.3005
R744 VDD2.n91 VDD2.n90 9.3005
R745 VDD2.n73 VDD2.n72 9.3005
R746 VDD2.n12 VDD2.n11 9.3005
R747 VDD2.n67 VDD2.n66 9.3005
R748 VDD2.n65 VDD2.n64 9.3005
R749 VDD2.n16 VDD2.n15 9.3005
R750 VDD2.n59 VDD2.n58 9.3005
R751 VDD2.n57 VDD2.n56 9.3005
R752 VDD2.n33 VDD2.n32 9.3005
R753 VDD2.n28 VDD2.n27 9.3005
R754 VDD2.n39 VDD2.n38 9.3005
R755 VDD2.n41 VDD2.n40 9.3005
R756 VDD2.n24 VDD2.n23 9.3005
R757 VDD2.n47 VDD2.n46 9.3005
R758 VDD2.n49 VDD2.n48 9.3005
R759 VDD2.n50 VDD2.n19 9.3005
R760 VDD2.n75 VDD2.n74 9.3005
R761 VDD2.n179 VDD2.n99 8.92171
R762 VDD2.n166 VDD2.n107 8.92171
R763 VDD2.n134 VDD2.n133 8.92171
R764 VDD2.n38 VDD2.n37 8.92171
R765 VDD2.n71 VDD2.n12 8.92171
R766 VDD2.n84 VDD2.n4 8.92171
R767 VDD2.n178 VDD2.n101 8.14595
R768 VDD2.n167 VDD2.n105 8.14595
R769 VDD2.n130 VDD2.n124 8.14595
R770 VDD2.n34 VDD2.n28 8.14595
R771 VDD2.n72 VDD2.n10 8.14595
R772 VDD2.n83 VDD2.n6 8.14595
R773 VDD2.n175 VDD2.n174 7.3702
R774 VDD2.n171 VDD2.n170 7.3702
R775 VDD2.n129 VDD2.n126 7.3702
R776 VDD2.n33 VDD2.n30 7.3702
R777 VDD2.n76 VDD2.n75 7.3702
R778 VDD2.n80 VDD2.n79 7.3702
R779 VDD2.n174 VDD2.n103 6.59444
R780 VDD2.n171 VDD2.n103 6.59444
R781 VDD2.n76 VDD2.n8 6.59444
R782 VDD2.n79 VDD2.n8 6.59444
R783 VDD2.n175 VDD2.n101 5.81868
R784 VDD2.n170 VDD2.n105 5.81868
R785 VDD2.n130 VDD2.n129 5.81868
R786 VDD2.n34 VDD2.n33 5.81868
R787 VDD2.n75 VDD2.n10 5.81868
R788 VDD2.n80 VDD2.n6 5.81868
R789 VDD2.n179 VDD2.n178 5.04292
R790 VDD2.n167 VDD2.n166 5.04292
R791 VDD2.n133 VDD2.n124 5.04292
R792 VDD2.n37 VDD2.n28 5.04292
R793 VDD2.n72 VDD2.n71 5.04292
R794 VDD2.n84 VDD2.n83 5.04292
R795 VDD2.n182 VDD2.n99 4.26717
R796 VDD2.n163 VDD2.n107 4.26717
R797 VDD2.n134 VDD2.n122 4.26717
R798 VDD2.n38 VDD2.n26 4.26717
R799 VDD2.n68 VDD2.n12 4.26717
R800 VDD2.n87 VDD2.n4 4.26717
R801 VDD2.n183 VDD2.n97 3.49141
R802 VDD2.n162 VDD2.n109 3.49141
R803 VDD2.n138 VDD2.n137 3.49141
R804 VDD2.n42 VDD2.n41 3.49141
R805 VDD2.n67 VDD2.n14 3.49141
R806 VDD2.n88 VDD2.n2 3.49141
R807 VDD2.n128 VDD2.n127 2.84303
R808 VDD2.n32 VDD2.n31 2.84303
R809 VDD2.n187 VDD2.n186 2.71565
R810 VDD2.n159 VDD2.n158 2.71565
R811 VDD2.n141 VDD2.n120 2.71565
R812 VDD2.n45 VDD2.n24 2.71565
R813 VDD2.n64 VDD2.n63 2.71565
R814 VDD2.n92 VDD2.n91 2.71565
R815 VDD2.n189 VDD2.n95 1.93989
R816 VDD2.n155 VDD2.n111 1.93989
R817 VDD2.n142 VDD2.n118 1.93989
R818 VDD2.n46 VDD2.n22 1.93989
R819 VDD2.n60 VDD2.n16 1.93989
R820 VDD2.n94 VDD2.n0 1.93989
R821 VDD2.n154 VDD2.n113 1.16414
R822 VDD2.n146 VDD2.n145 1.16414
R823 VDD2.n51 VDD2.n49 1.16414
R824 VDD2.n59 VDD2.n18 1.16414
R825 VDD2.n151 VDD2.n150 0.388379
R826 VDD2.n117 VDD2.n115 0.388379
R827 VDD2.n50 VDD2.n20 0.388379
R828 VDD2.n56 VDD2.n55 0.388379
R829 VDD2 VDD2.n190 0.265586
R830 VDD2.n185 VDD2.n184 0.155672
R831 VDD2.n184 VDD2.n98 0.155672
R832 VDD2.n177 VDD2.n98 0.155672
R833 VDD2.n177 VDD2.n176 0.155672
R834 VDD2.n176 VDD2.n102 0.155672
R835 VDD2.n169 VDD2.n102 0.155672
R836 VDD2.n169 VDD2.n168 0.155672
R837 VDD2.n168 VDD2.n106 0.155672
R838 VDD2.n161 VDD2.n106 0.155672
R839 VDD2.n161 VDD2.n160 0.155672
R840 VDD2.n160 VDD2.n110 0.155672
R841 VDD2.n153 VDD2.n110 0.155672
R842 VDD2.n153 VDD2.n152 0.155672
R843 VDD2.n152 VDD2.n114 0.155672
R844 VDD2.n144 VDD2.n114 0.155672
R845 VDD2.n144 VDD2.n143 0.155672
R846 VDD2.n143 VDD2.n119 0.155672
R847 VDD2.n136 VDD2.n119 0.155672
R848 VDD2.n136 VDD2.n135 0.155672
R849 VDD2.n135 VDD2.n123 0.155672
R850 VDD2.n128 VDD2.n123 0.155672
R851 VDD2.n32 VDD2.n27 0.155672
R852 VDD2.n39 VDD2.n27 0.155672
R853 VDD2.n40 VDD2.n39 0.155672
R854 VDD2.n40 VDD2.n23 0.155672
R855 VDD2.n47 VDD2.n23 0.155672
R856 VDD2.n48 VDD2.n47 0.155672
R857 VDD2.n48 VDD2.n19 0.155672
R858 VDD2.n57 VDD2.n19 0.155672
R859 VDD2.n58 VDD2.n57 0.155672
R860 VDD2.n58 VDD2.n15 0.155672
R861 VDD2.n65 VDD2.n15 0.155672
R862 VDD2.n66 VDD2.n65 0.155672
R863 VDD2.n66 VDD2.n11 0.155672
R864 VDD2.n73 VDD2.n11 0.155672
R865 VDD2.n74 VDD2.n73 0.155672
R866 VDD2.n74 VDD2.n7 0.155672
R867 VDD2.n81 VDD2.n7 0.155672
R868 VDD2.n82 VDD2.n81 0.155672
R869 VDD2.n82 VDD2.n3 0.155672
R870 VDD2.n89 VDD2.n3 0.155672
R871 VDD2.n90 VDD2.n89 0.155672
R872 B.n93 B.t2 868.01
R873 B.n91 B.t13 868.01
R874 B.n432 B.t10 868.01
R875 B.n429 B.t6 868.01
R876 B.n740 B.n739 585
R877 B.n341 B.n90 585
R878 B.n340 B.n339 585
R879 B.n338 B.n337 585
R880 B.n336 B.n335 585
R881 B.n334 B.n333 585
R882 B.n332 B.n331 585
R883 B.n330 B.n329 585
R884 B.n328 B.n327 585
R885 B.n326 B.n325 585
R886 B.n324 B.n323 585
R887 B.n322 B.n321 585
R888 B.n320 B.n319 585
R889 B.n318 B.n317 585
R890 B.n316 B.n315 585
R891 B.n314 B.n313 585
R892 B.n312 B.n311 585
R893 B.n310 B.n309 585
R894 B.n308 B.n307 585
R895 B.n306 B.n305 585
R896 B.n304 B.n303 585
R897 B.n302 B.n301 585
R898 B.n300 B.n299 585
R899 B.n298 B.n297 585
R900 B.n296 B.n295 585
R901 B.n294 B.n293 585
R902 B.n292 B.n291 585
R903 B.n290 B.n289 585
R904 B.n288 B.n287 585
R905 B.n286 B.n285 585
R906 B.n284 B.n283 585
R907 B.n282 B.n281 585
R908 B.n280 B.n279 585
R909 B.n278 B.n277 585
R910 B.n276 B.n275 585
R911 B.n274 B.n273 585
R912 B.n272 B.n271 585
R913 B.n270 B.n269 585
R914 B.n268 B.n267 585
R915 B.n266 B.n265 585
R916 B.n264 B.n263 585
R917 B.n262 B.n261 585
R918 B.n260 B.n259 585
R919 B.n258 B.n257 585
R920 B.n256 B.n255 585
R921 B.n254 B.n253 585
R922 B.n252 B.n251 585
R923 B.n250 B.n249 585
R924 B.n248 B.n247 585
R925 B.n246 B.n245 585
R926 B.n244 B.n243 585
R927 B.n242 B.n241 585
R928 B.n240 B.n239 585
R929 B.n238 B.n237 585
R930 B.n236 B.n235 585
R931 B.n234 B.n233 585
R932 B.n232 B.n231 585
R933 B.n229 B.n228 585
R934 B.n227 B.n226 585
R935 B.n225 B.n224 585
R936 B.n223 B.n222 585
R937 B.n221 B.n220 585
R938 B.n219 B.n218 585
R939 B.n217 B.n216 585
R940 B.n215 B.n214 585
R941 B.n213 B.n212 585
R942 B.n211 B.n210 585
R943 B.n208 B.n207 585
R944 B.n206 B.n205 585
R945 B.n204 B.n203 585
R946 B.n202 B.n201 585
R947 B.n200 B.n199 585
R948 B.n198 B.n197 585
R949 B.n196 B.n195 585
R950 B.n194 B.n193 585
R951 B.n192 B.n191 585
R952 B.n190 B.n189 585
R953 B.n188 B.n187 585
R954 B.n186 B.n185 585
R955 B.n184 B.n183 585
R956 B.n182 B.n181 585
R957 B.n180 B.n179 585
R958 B.n178 B.n177 585
R959 B.n176 B.n175 585
R960 B.n174 B.n173 585
R961 B.n172 B.n171 585
R962 B.n170 B.n169 585
R963 B.n168 B.n167 585
R964 B.n166 B.n165 585
R965 B.n164 B.n163 585
R966 B.n162 B.n161 585
R967 B.n160 B.n159 585
R968 B.n158 B.n157 585
R969 B.n156 B.n155 585
R970 B.n154 B.n153 585
R971 B.n152 B.n151 585
R972 B.n150 B.n149 585
R973 B.n148 B.n147 585
R974 B.n146 B.n145 585
R975 B.n144 B.n143 585
R976 B.n142 B.n141 585
R977 B.n140 B.n139 585
R978 B.n138 B.n137 585
R979 B.n136 B.n135 585
R980 B.n134 B.n133 585
R981 B.n132 B.n131 585
R982 B.n130 B.n129 585
R983 B.n128 B.n127 585
R984 B.n126 B.n125 585
R985 B.n124 B.n123 585
R986 B.n122 B.n121 585
R987 B.n120 B.n119 585
R988 B.n118 B.n117 585
R989 B.n116 B.n115 585
R990 B.n114 B.n113 585
R991 B.n112 B.n111 585
R992 B.n110 B.n109 585
R993 B.n108 B.n107 585
R994 B.n106 B.n105 585
R995 B.n104 B.n103 585
R996 B.n102 B.n101 585
R997 B.n100 B.n99 585
R998 B.n98 B.n97 585
R999 B.n96 B.n95 585
R1000 B.n738 B.n28 585
R1001 B.n743 B.n28 585
R1002 B.n737 B.n27 585
R1003 B.n744 B.n27 585
R1004 B.n736 B.n735 585
R1005 B.n735 B.n23 585
R1006 B.n734 B.n22 585
R1007 B.n750 B.n22 585
R1008 B.n733 B.n21 585
R1009 B.n751 B.n21 585
R1010 B.n732 B.n20 585
R1011 B.n752 B.n20 585
R1012 B.n731 B.n730 585
R1013 B.n730 B.n16 585
R1014 B.n729 B.n15 585
R1015 B.n758 B.n15 585
R1016 B.n728 B.n14 585
R1017 B.n759 B.n14 585
R1018 B.n727 B.n13 585
R1019 B.n760 B.n13 585
R1020 B.n726 B.n725 585
R1021 B.n725 B.n12 585
R1022 B.n724 B.n723 585
R1023 B.n724 B.n8 585
R1024 B.n722 B.n7 585
R1025 B.n767 B.n7 585
R1026 B.n721 B.n6 585
R1027 B.n768 B.n6 585
R1028 B.n720 B.n5 585
R1029 B.n769 B.n5 585
R1030 B.n719 B.n718 585
R1031 B.n718 B.n4 585
R1032 B.n717 B.n342 585
R1033 B.n717 B.n716 585
R1034 B.n706 B.n343 585
R1035 B.n709 B.n343 585
R1036 B.n708 B.n707 585
R1037 B.n710 B.n708 585
R1038 B.n705 B.n348 585
R1039 B.n348 B.n347 585
R1040 B.n704 B.n703 585
R1041 B.n703 B.n702 585
R1042 B.n350 B.n349 585
R1043 B.n351 B.n350 585
R1044 B.n695 B.n694 585
R1045 B.n696 B.n695 585
R1046 B.n693 B.n355 585
R1047 B.n359 B.n355 585
R1048 B.n692 B.n691 585
R1049 B.n691 B.n690 585
R1050 B.n357 B.n356 585
R1051 B.n358 B.n357 585
R1052 B.n683 B.n682 585
R1053 B.n684 B.n683 585
R1054 B.n681 B.n364 585
R1055 B.n364 B.n363 585
R1056 B.n676 B.n675 585
R1057 B.n674 B.n428 585
R1058 B.n673 B.n427 585
R1059 B.n678 B.n427 585
R1060 B.n672 B.n671 585
R1061 B.n670 B.n669 585
R1062 B.n668 B.n667 585
R1063 B.n666 B.n665 585
R1064 B.n664 B.n663 585
R1065 B.n662 B.n661 585
R1066 B.n660 B.n659 585
R1067 B.n658 B.n657 585
R1068 B.n656 B.n655 585
R1069 B.n654 B.n653 585
R1070 B.n652 B.n651 585
R1071 B.n650 B.n649 585
R1072 B.n648 B.n647 585
R1073 B.n646 B.n645 585
R1074 B.n644 B.n643 585
R1075 B.n642 B.n641 585
R1076 B.n640 B.n639 585
R1077 B.n638 B.n637 585
R1078 B.n636 B.n635 585
R1079 B.n634 B.n633 585
R1080 B.n632 B.n631 585
R1081 B.n630 B.n629 585
R1082 B.n628 B.n627 585
R1083 B.n626 B.n625 585
R1084 B.n624 B.n623 585
R1085 B.n622 B.n621 585
R1086 B.n620 B.n619 585
R1087 B.n618 B.n617 585
R1088 B.n616 B.n615 585
R1089 B.n614 B.n613 585
R1090 B.n612 B.n611 585
R1091 B.n610 B.n609 585
R1092 B.n608 B.n607 585
R1093 B.n606 B.n605 585
R1094 B.n604 B.n603 585
R1095 B.n602 B.n601 585
R1096 B.n600 B.n599 585
R1097 B.n598 B.n597 585
R1098 B.n596 B.n595 585
R1099 B.n594 B.n593 585
R1100 B.n592 B.n591 585
R1101 B.n590 B.n589 585
R1102 B.n588 B.n587 585
R1103 B.n586 B.n585 585
R1104 B.n584 B.n583 585
R1105 B.n582 B.n581 585
R1106 B.n580 B.n579 585
R1107 B.n578 B.n577 585
R1108 B.n576 B.n575 585
R1109 B.n574 B.n573 585
R1110 B.n572 B.n571 585
R1111 B.n570 B.n569 585
R1112 B.n568 B.n567 585
R1113 B.n566 B.n565 585
R1114 B.n564 B.n563 585
R1115 B.n562 B.n561 585
R1116 B.n560 B.n559 585
R1117 B.n558 B.n557 585
R1118 B.n556 B.n555 585
R1119 B.n554 B.n553 585
R1120 B.n552 B.n551 585
R1121 B.n550 B.n549 585
R1122 B.n548 B.n547 585
R1123 B.n546 B.n545 585
R1124 B.n544 B.n543 585
R1125 B.n542 B.n541 585
R1126 B.n540 B.n539 585
R1127 B.n538 B.n537 585
R1128 B.n536 B.n535 585
R1129 B.n534 B.n533 585
R1130 B.n532 B.n531 585
R1131 B.n530 B.n529 585
R1132 B.n528 B.n527 585
R1133 B.n526 B.n525 585
R1134 B.n524 B.n523 585
R1135 B.n522 B.n521 585
R1136 B.n520 B.n519 585
R1137 B.n518 B.n517 585
R1138 B.n516 B.n515 585
R1139 B.n514 B.n513 585
R1140 B.n512 B.n511 585
R1141 B.n510 B.n509 585
R1142 B.n508 B.n507 585
R1143 B.n506 B.n505 585
R1144 B.n504 B.n503 585
R1145 B.n502 B.n501 585
R1146 B.n500 B.n499 585
R1147 B.n498 B.n497 585
R1148 B.n496 B.n495 585
R1149 B.n494 B.n493 585
R1150 B.n492 B.n491 585
R1151 B.n490 B.n489 585
R1152 B.n488 B.n487 585
R1153 B.n486 B.n485 585
R1154 B.n484 B.n483 585
R1155 B.n482 B.n481 585
R1156 B.n480 B.n479 585
R1157 B.n478 B.n477 585
R1158 B.n476 B.n475 585
R1159 B.n474 B.n473 585
R1160 B.n472 B.n471 585
R1161 B.n470 B.n469 585
R1162 B.n468 B.n467 585
R1163 B.n466 B.n465 585
R1164 B.n464 B.n463 585
R1165 B.n462 B.n461 585
R1166 B.n460 B.n459 585
R1167 B.n458 B.n457 585
R1168 B.n456 B.n455 585
R1169 B.n454 B.n453 585
R1170 B.n452 B.n451 585
R1171 B.n450 B.n449 585
R1172 B.n448 B.n447 585
R1173 B.n446 B.n445 585
R1174 B.n444 B.n443 585
R1175 B.n442 B.n441 585
R1176 B.n440 B.n439 585
R1177 B.n438 B.n437 585
R1178 B.n436 B.n435 585
R1179 B.n366 B.n365 585
R1180 B.n680 B.n679 585
R1181 B.n679 B.n678 585
R1182 B.n362 B.n361 585
R1183 B.n363 B.n362 585
R1184 B.n686 B.n685 585
R1185 B.n685 B.n684 585
R1186 B.n687 B.n360 585
R1187 B.n360 B.n358 585
R1188 B.n689 B.n688 585
R1189 B.n690 B.n689 585
R1190 B.n354 B.n353 585
R1191 B.n359 B.n354 585
R1192 B.n698 B.n697 585
R1193 B.n697 B.n696 585
R1194 B.n699 B.n352 585
R1195 B.n352 B.n351 585
R1196 B.n701 B.n700 585
R1197 B.n702 B.n701 585
R1198 B.n346 B.n345 585
R1199 B.n347 B.n346 585
R1200 B.n712 B.n711 585
R1201 B.n711 B.n710 585
R1202 B.n713 B.n344 585
R1203 B.n709 B.n344 585
R1204 B.n715 B.n714 585
R1205 B.n716 B.n715 585
R1206 B.n3 B.n0 585
R1207 B.n4 B.n3 585
R1208 B.n766 B.n1 585
R1209 B.n767 B.n766 585
R1210 B.n765 B.n764 585
R1211 B.n765 B.n8 585
R1212 B.n763 B.n9 585
R1213 B.n12 B.n9 585
R1214 B.n762 B.n761 585
R1215 B.n761 B.n760 585
R1216 B.n11 B.n10 585
R1217 B.n759 B.n11 585
R1218 B.n757 B.n756 585
R1219 B.n758 B.n757 585
R1220 B.n755 B.n17 585
R1221 B.n17 B.n16 585
R1222 B.n754 B.n753 585
R1223 B.n753 B.n752 585
R1224 B.n19 B.n18 585
R1225 B.n751 B.n19 585
R1226 B.n749 B.n748 585
R1227 B.n750 B.n749 585
R1228 B.n747 B.n24 585
R1229 B.n24 B.n23 585
R1230 B.n746 B.n745 585
R1231 B.n745 B.n744 585
R1232 B.n26 B.n25 585
R1233 B.n743 B.n26 585
R1234 B.n770 B.n769 585
R1235 B.n768 B.n2 585
R1236 B.n95 B.n26 578.989
R1237 B.n740 B.n28 578.989
R1238 B.n679 B.n364 578.989
R1239 B.n676 B.n362 578.989
R1240 B.n91 B.t14 392.774
R1241 B.n432 B.t12 392.774
R1242 B.n93 B.t4 392.774
R1243 B.n429 B.t9 392.774
R1244 B.n92 B.t15 374.156
R1245 B.n433 B.t11 374.156
R1246 B.n94 B.t5 374.156
R1247 B.n430 B.t8 374.156
R1248 B.n742 B.n741 256.663
R1249 B.n742 B.n89 256.663
R1250 B.n742 B.n88 256.663
R1251 B.n742 B.n87 256.663
R1252 B.n742 B.n86 256.663
R1253 B.n742 B.n85 256.663
R1254 B.n742 B.n84 256.663
R1255 B.n742 B.n83 256.663
R1256 B.n742 B.n82 256.663
R1257 B.n742 B.n81 256.663
R1258 B.n742 B.n80 256.663
R1259 B.n742 B.n79 256.663
R1260 B.n742 B.n78 256.663
R1261 B.n742 B.n77 256.663
R1262 B.n742 B.n76 256.663
R1263 B.n742 B.n75 256.663
R1264 B.n742 B.n74 256.663
R1265 B.n742 B.n73 256.663
R1266 B.n742 B.n72 256.663
R1267 B.n742 B.n71 256.663
R1268 B.n742 B.n70 256.663
R1269 B.n742 B.n69 256.663
R1270 B.n742 B.n68 256.663
R1271 B.n742 B.n67 256.663
R1272 B.n742 B.n66 256.663
R1273 B.n742 B.n65 256.663
R1274 B.n742 B.n64 256.663
R1275 B.n742 B.n63 256.663
R1276 B.n742 B.n62 256.663
R1277 B.n742 B.n61 256.663
R1278 B.n742 B.n60 256.663
R1279 B.n742 B.n59 256.663
R1280 B.n742 B.n58 256.663
R1281 B.n742 B.n57 256.663
R1282 B.n742 B.n56 256.663
R1283 B.n742 B.n55 256.663
R1284 B.n742 B.n54 256.663
R1285 B.n742 B.n53 256.663
R1286 B.n742 B.n52 256.663
R1287 B.n742 B.n51 256.663
R1288 B.n742 B.n50 256.663
R1289 B.n742 B.n49 256.663
R1290 B.n742 B.n48 256.663
R1291 B.n742 B.n47 256.663
R1292 B.n742 B.n46 256.663
R1293 B.n742 B.n45 256.663
R1294 B.n742 B.n44 256.663
R1295 B.n742 B.n43 256.663
R1296 B.n742 B.n42 256.663
R1297 B.n742 B.n41 256.663
R1298 B.n742 B.n40 256.663
R1299 B.n742 B.n39 256.663
R1300 B.n742 B.n38 256.663
R1301 B.n742 B.n37 256.663
R1302 B.n742 B.n36 256.663
R1303 B.n742 B.n35 256.663
R1304 B.n742 B.n34 256.663
R1305 B.n742 B.n33 256.663
R1306 B.n742 B.n32 256.663
R1307 B.n742 B.n31 256.663
R1308 B.n742 B.n30 256.663
R1309 B.n742 B.n29 256.663
R1310 B.n678 B.n677 256.663
R1311 B.n678 B.n367 256.663
R1312 B.n678 B.n368 256.663
R1313 B.n678 B.n369 256.663
R1314 B.n678 B.n370 256.663
R1315 B.n678 B.n371 256.663
R1316 B.n678 B.n372 256.663
R1317 B.n678 B.n373 256.663
R1318 B.n678 B.n374 256.663
R1319 B.n678 B.n375 256.663
R1320 B.n678 B.n376 256.663
R1321 B.n678 B.n377 256.663
R1322 B.n678 B.n378 256.663
R1323 B.n678 B.n379 256.663
R1324 B.n678 B.n380 256.663
R1325 B.n678 B.n381 256.663
R1326 B.n678 B.n382 256.663
R1327 B.n678 B.n383 256.663
R1328 B.n678 B.n384 256.663
R1329 B.n678 B.n385 256.663
R1330 B.n678 B.n386 256.663
R1331 B.n678 B.n387 256.663
R1332 B.n678 B.n388 256.663
R1333 B.n678 B.n389 256.663
R1334 B.n678 B.n390 256.663
R1335 B.n678 B.n391 256.663
R1336 B.n678 B.n392 256.663
R1337 B.n678 B.n393 256.663
R1338 B.n678 B.n394 256.663
R1339 B.n678 B.n395 256.663
R1340 B.n678 B.n396 256.663
R1341 B.n678 B.n397 256.663
R1342 B.n678 B.n398 256.663
R1343 B.n678 B.n399 256.663
R1344 B.n678 B.n400 256.663
R1345 B.n678 B.n401 256.663
R1346 B.n678 B.n402 256.663
R1347 B.n678 B.n403 256.663
R1348 B.n678 B.n404 256.663
R1349 B.n678 B.n405 256.663
R1350 B.n678 B.n406 256.663
R1351 B.n678 B.n407 256.663
R1352 B.n678 B.n408 256.663
R1353 B.n678 B.n409 256.663
R1354 B.n678 B.n410 256.663
R1355 B.n678 B.n411 256.663
R1356 B.n678 B.n412 256.663
R1357 B.n678 B.n413 256.663
R1358 B.n678 B.n414 256.663
R1359 B.n678 B.n415 256.663
R1360 B.n678 B.n416 256.663
R1361 B.n678 B.n417 256.663
R1362 B.n678 B.n418 256.663
R1363 B.n678 B.n419 256.663
R1364 B.n678 B.n420 256.663
R1365 B.n678 B.n421 256.663
R1366 B.n678 B.n422 256.663
R1367 B.n678 B.n423 256.663
R1368 B.n678 B.n424 256.663
R1369 B.n678 B.n425 256.663
R1370 B.n678 B.n426 256.663
R1371 B.n772 B.n771 256.663
R1372 B.n99 B.n98 163.367
R1373 B.n103 B.n102 163.367
R1374 B.n107 B.n106 163.367
R1375 B.n111 B.n110 163.367
R1376 B.n115 B.n114 163.367
R1377 B.n119 B.n118 163.367
R1378 B.n123 B.n122 163.367
R1379 B.n127 B.n126 163.367
R1380 B.n131 B.n130 163.367
R1381 B.n135 B.n134 163.367
R1382 B.n139 B.n138 163.367
R1383 B.n143 B.n142 163.367
R1384 B.n147 B.n146 163.367
R1385 B.n151 B.n150 163.367
R1386 B.n155 B.n154 163.367
R1387 B.n159 B.n158 163.367
R1388 B.n163 B.n162 163.367
R1389 B.n167 B.n166 163.367
R1390 B.n171 B.n170 163.367
R1391 B.n175 B.n174 163.367
R1392 B.n179 B.n178 163.367
R1393 B.n183 B.n182 163.367
R1394 B.n187 B.n186 163.367
R1395 B.n191 B.n190 163.367
R1396 B.n195 B.n194 163.367
R1397 B.n199 B.n198 163.367
R1398 B.n203 B.n202 163.367
R1399 B.n207 B.n206 163.367
R1400 B.n212 B.n211 163.367
R1401 B.n216 B.n215 163.367
R1402 B.n220 B.n219 163.367
R1403 B.n224 B.n223 163.367
R1404 B.n228 B.n227 163.367
R1405 B.n233 B.n232 163.367
R1406 B.n237 B.n236 163.367
R1407 B.n241 B.n240 163.367
R1408 B.n245 B.n244 163.367
R1409 B.n249 B.n248 163.367
R1410 B.n253 B.n252 163.367
R1411 B.n257 B.n256 163.367
R1412 B.n261 B.n260 163.367
R1413 B.n265 B.n264 163.367
R1414 B.n269 B.n268 163.367
R1415 B.n273 B.n272 163.367
R1416 B.n277 B.n276 163.367
R1417 B.n281 B.n280 163.367
R1418 B.n285 B.n284 163.367
R1419 B.n289 B.n288 163.367
R1420 B.n293 B.n292 163.367
R1421 B.n297 B.n296 163.367
R1422 B.n301 B.n300 163.367
R1423 B.n305 B.n304 163.367
R1424 B.n309 B.n308 163.367
R1425 B.n313 B.n312 163.367
R1426 B.n317 B.n316 163.367
R1427 B.n321 B.n320 163.367
R1428 B.n325 B.n324 163.367
R1429 B.n329 B.n328 163.367
R1430 B.n333 B.n332 163.367
R1431 B.n337 B.n336 163.367
R1432 B.n339 B.n90 163.367
R1433 B.n683 B.n364 163.367
R1434 B.n683 B.n357 163.367
R1435 B.n691 B.n357 163.367
R1436 B.n691 B.n355 163.367
R1437 B.n695 B.n355 163.367
R1438 B.n695 B.n350 163.367
R1439 B.n703 B.n350 163.367
R1440 B.n703 B.n348 163.367
R1441 B.n708 B.n348 163.367
R1442 B.n708 B.n343 163.367
R1443 B.n717 B.n343 163.367
R1444 B.n718 B.n717 163.367
R1445 B.n718 B.n5 163.367
R1446 B.n6 B.n5 163.367
R1447 B.n7 B.n6 163.367
R1448 B.n724 B.n7 163.367
R1449 B.n725 B.n724 163.367
R1450 B.n725 B.n13 163.367
R1451 B.n14 B.n13 163.367
R1452 B.n15 B.n14 163.367
R1453 B.n730 B.n15 163.367
R1454 B.n730 B.n20 163.367
R1455 B.n21 B.n20 163.367
R1456 B.n22 B.n21 163.367
R1457 B.n735 B.n22 163.367
R1458 B.n735 B.n27 163.367
R1459 B.n28 B.n27 163.367
R1460 B.n428 B.n427 163.367
R1461 B.n671 B.n427 163.367
R1462 B.n669 B.n668 163.367
R1463 B.n665 B.n664 163.367
R1464 B.n661 B.n660 163.367
R1465 B.n657 B.n656 163.367
R1466 B.n653 B.n652 163.367
R1467 B.n649 B.n648 163.367
R1468 B.n645 B.n644 163.367
R1469 B.n641 B.n640 163.367
R1470 B.n637 B.n636 163.367
R1471 B.n633 B.n632 163.367
R1472 B.n629 B.n628 163.367
R1473 B.n625 B.n624 163.367
R1474 B.n621 B.n620 163.367
R1475 B.n617 B.n616 163.367
R1476 B.n613 B.n612 163.367
R1477 B.n609 B.n608 163.367
R1478 B.n605 B.n604 163.367
R1479 B.n601 B.n600 163.367
R1480 B.n597 B.n596 163.367
R1481 B.n593 B.n592 163.367
R1482 B.n589 B.n588 163.367
R1483 B.n585 B.n584 163.367
R1484 B.n581 B.n580 163.367
R1485 B.n577 B.n576 163.367
R1486 B.n573 B.n572 163.367
R1487 B.n569 B.n568 163.367
R1488 B.n565 B.n564 163.367
R1489 B.n561 B.n560 163.367
R1490 B.n557 B.n556 163.367
R1491 B.n553 B.n552 163.367
R1492 B.n549 B.n548 163.367
R1493 B.n545 B.n544 163.367
R1494 B.n541 B.n540 163.367
R1495 B.n537 B.n536 163.367
R1496 B.n533 B.n532 163.367
R1497 B.n529 B.n528 163.367
R1498 B.n525 B.n524 163.367
R1499 B.n521 B.n520 163.367
R1500 B.n517 B.n516 163.367
R1501 B.n513 B.n512 163.367
R1502 B.n509 B.n508 163.367
R1503 B.n505 B.n504 163.367
R1504 B.n501 B.n500 163.367
R1505 B.n497 B.n496 163.367
R1506 B.n493 B.n492 163.367
R1507 B.n489 B.n488 163.367
R1508 B.n485 B.n484 163.367
R1509 B.n481 B.n480 163.367
R1510 B.n477 B.n476 163.367
R1511 B.n473 B.n472 163.367
R1512 B.n469 B.n468 163.367
R1513 B.n465 B.n464 163.367
R1514 B.n461 B.n460 163.367
R1515 B.n457 B.n456 163.367
R1516 B.n453 B.n452 163.367
R1517 B.n449 B.n448 163.367
R1518 B.n445 B.n444 163.367
R1519 B.n441 B.n440 163.367
R1520 B.n437 B.n436 163.367
R1521 B.n679 B.n366 163.367
R1522 B.n685 B.n362 163.367
R1523 B.n685 B.n360 163.367
R1524 B.n689 B.n360 163.367
R1525 B.n689 B.n354 163.367
R1526 B.n697 B.n354 163.367
R1527 B.n697 B.n352 163.367
R1528 B.n701 B.n352 163.367
R1529 B.n701 B.n346 163.367
R1530 B.n711 B.n346 163.367
R1531 B.n711 B.n344 163.367
R1532 B.n715 B.n344 163.367
R1533 B.n715 B.n3 163.367
R1534 B.n770 B.n3 163.367
R1535 B.n766 B.n2 163.367
R1536 B.n766 B.n765 163.367
R1537 B.n765 B.n9 163.367
R1538 B.n761 B.n9 163.367
R1539 B.n761 B.n11 163.367
R1540 B.n757 B.n11 163.367
R1541 B.n757 B.n17 163.367
R1542 B.n753 B.n17 163.367
R1543 B.n753 B.n19 163.367
R1544 B.n749 B.n19 163.367
R1545 B.n749 B.n24 163.367
R1546 B.n745 B.n24 163.367
R1547 B.n745 B.n26 163.367
R1548 B.n95 B.n29 71.676
R1549 B.n99 B.n30 71.676
R1550 B.n103 B.n31 71.676
R1551 B.n107 B.n32 71.676
R1552 B.n111 B.n33 71.676
R1553 B.n115 B.n34 71.676
R1554 B.n119 B.n35 71.676
R1555 B.n123 B.n36 71.676
R1556 B.n127 B.n37 71.676
R1557 B.n131 B.n38 71.676
R1558 B.n135 B.n39 71.676
R1559 B.n139 B.n40 71.676
R1560 B.n143 B.n41 71.676
R1561 B.n147 B.n42 71.676
R1562 B.n151 B.n43 71.676
R1563 B.n155 B.n44 71.676
R1564 B.n159 B.n45 71.676
R1565 B.n163 B.n46 71.676
R1566 B.n167 B.n47 71.676
R1567 B.n171 B.n48 71.676
R1568 B.n175 B.n49 71.676
R1569 B.n179 B.n50 71.676
R1570 B.n183 B.n51 71.676
R1571 B.n187 B.n52 71.676
R1572 B.n191 B.n53 71.676
R1573 B.n195 B.n54 71.676
R1574 B.n199 B.n55 71.676
R1575 B.n203 B.n56 71.676
R1576 B.n207 B.n57 71.676
R1577 B.n212 B.n58 71.676
R1578 B.n216 B.n59 71.676
R1579 B.n220 B.n60 71.676
R1580 B.n224 B.n61 71.676
R1581 B.n228 B.n62 71.676
R1582 B.n233 B.n63 71.676
R1583 B.n237 B.n64 71.676
R1584 B.n241 B.n65 71.676
R1585 B.n245 B.n66 71.676
R1586 B.n249 B.n67 71.676
R1587 B.n253 B.n68 71.676
R1588 B.n257 B.n69 71.676
R1589 B.n261 B.n70 71.676
R1590 B.n265 B.n71 71.676
R1591 B.n269 B.n72 71.676
R1592 B.n273 B.n73 71.676
R1593 B.n277 B.n74 71.676
R1594 B.n281 B.n75 71.676
R1595 B.n285 B.n76 71.676
R1596 B.n289 B.n77 71.676
R1597 B.n293 B.n78 71.676
R1598 B.n297 B.n79 71.676
R1599 B.n301 B.n80 71.676
R1600 B.n305 B.n81 71.676
R1601 B.n309 B.n82 71.676
R1602 B.n313 B.n83 71.676
R1603 B.n317 B.n84 71.676
R1604 B.n321 B.n85 71.676
R1605 B.n325 B.n86 71.676
R1606 B.n329 B.n87 71.676
R1607 B.n333 B.n88 71.676
R1608 B.n337 B.n89 71.676
R1609 B.n741 B.n90 71.676
R1610 B.n741 B.n740 71.676
R1611 B.n339 B.n89 71.676
R1612 B.n336 B.n88 71.676
R1613 B.n332 B.n87 71.676
R1614 B.n328 B.n86 71.676
R1615 B.n324 B.n85 71.676
R1616 B.n320 B.n84 71.676
R1617 B.n316 B.n83 71.676
R1618 B.n312 B.n82 71.676
R1619 B.n308 B.n81 71.676
R1620 B.n304 B.n80 71.676
R1621 B.n300 B.n79 71.676
R1622 B.n296 B.n78 71.676
R1623 B.n292 B.n77 71.676
R1624 B.n288 B.n76 71.676
R1625 B.n284 B.n75 71.676
R1626 B.n280 B.n74 71.676
R1627 B.n276 B.n73 71.676
R1628 B.n272 B.n72 71.676
R1629 B.n268 B.n71 71.676
R1630 B.n264 B.n70 71.676
R1631 B.n260 B.n69 71.676
R1632 B.n256 B.n68 71.676
R1633 B.n252 B.n67 71.676
R1634 B.n248 B.n66 71.676
R1635 B.n244 B.n65 71.676
R1636 B.n240 B.n64 71.676
R1637 B.n236 B.n63 71.676
R1638 B.n232 B.n62 71.676
R1639 B.n227 B.n61 71.676
R1640 B.n223 B.n60 71.676
R1641 B.n219 B.n59 71.676
R1642 B.n215 B.n58 71.676
R1643 B.n211 B.n57 71.676
R1644 B.n206 B.n56 71.676
R1645 B.n202 B.n55 71.676
R1646 B.n198 B.n54 71.676
R1647 B.n194 B.n53 71.676
R1648 B.n190 B.n52 71.676
R1649 B.n186 B.n51 71.676
R1650 B.n182 B.n50 71.676
R1651 B.n178 B.n49 71.676
R1652 B.n174 B.n48 71.676
R1653 B.n170 B.n47 71.676
R1654 B.n166 B.n46 71.676
R1655 B.n162 B.n45 71.676
R1656 B.n158 B.n44 71.676
R1657 B.n154 B.n43 71.676
R1658 B.n150 B.n42 71.676
R1659 B.n146 B.n41 71.676
R1660 B.n142 B.n40 71.676
R1661 B.n138 B.n39 71.676
R1662 B.n134 B.n38 71.676
R1663 B.n130 B.n37 71.676
R1664 B.n126 B.n36 71.676
R1665 B.n122 B.n35 71.676
R1666 B.n118 B.n34 71.676
R1667 B.n114 B.n33 71.676
R1668 B.n110 B.n32 71.676
R1669 B.n106 B.n31 71.676
R1670 B.n102 B.n30 71.676
R1671 B.n98 B.n29 71.676
R1672 B.n677 B.n676 71.676
R1673 B.n671 B.n367 71.676
R1674 B.n668 B.n368 71.676
R1675 B.n664 B.n369 71.676
R1676 B.n660 B.n370 71.676
R1677 B.n656 B.n371 71.676
R1678 B.n652 B.n372 71.676
R1679 B.n648 B.n373 71.676
R1680 B.n644 B.n374 71.676
R1681 B.n640 B.n375 71.676
R1682 B.n636 B.n376 71.676
R1683 B.n632 B.n377 71.676
R1684 B.n628 B.n378 71.676
R1685 B.n624 B.n379 71.676
R1686 B.n620 B.n380 71.676
R1687 B.n616 B.n381 71.676
R1688 B.n612 B.n382 71.676
R1689 B.n608 B.n383 71.676
R1690 B.n604 B.n384 71.676
R1691 B.n600 B.n385 71.676
R1692 B.n596 B.n386 71.676
R1693 B.n592 B.n387 71.676
R1694 B.n588 B.n388 71.676
R1695 B.n584 B.n389 71.676
R1696 B.n580 B.n390 71.676
R1697 B.n576 B.n391 71.676
R1698 B.n572 B.n392 71.676
R1699 B.n568 B.n393 71.676
R1700 B.n564 B.n394 71.676
R1701 B.n560 B.n395 71.676
R1702 B.n556 B.n396 71.676
R1703 B.n552 B.n397 71.676
R1704 B.n548 B.n398 71.676
R1705 B.n544 B.n399 71.676
R1706 B.n540 B.n400 71.676
R1707 B.n536 B.n401 71.676
R1708 B.n532 B.n402 71.676
R1709 B.n528 B.n403 71.676
R1710 B.n524 B.n404 71.676
R1711 B.n520 B.n405 71.676
R1712 B.n516 B.n406 71.676
R1713 B.n512 B.n407 71.676
R1714 B.n508 B.n408 71.676
R1715 B.n504 B.n409 71.676
R1716 B.n500 B.n410 71.676
R1717 B.n496 B.n411 71.676
R1718 B.n492 B.n412 71.676
R1719 B.n488 B.n413 71.676
R1720 B.n484 B.n414 71.676
R1721 B.n480 B.n415 71.676
R1722 B.n476 B.n416 71.676
R1723 B.n472 B.n417 71.676
R1724 B.n468 B.n418 71.676
R1725 B.n464 B.n419 71.676
R1726 B.n460 B.n420 71.676
R1727 B.n456 B.n421 71.676
R1728 B.n452 B.n422 71.676
R1729 B.n448 B.n423 71.676
R1730 B.n444 B.n424 71.676
R1731 B.n440 B.n425 71.676
R1732 B.n436 B.n426 71.676
R1733 B.n677 B.n428 71.676
R1734 B.n669 B.n367 71.676
R1735 B.n665 B.n368 71.676
R1736 B.n661 B.n369 71.676
R1737 B.n657 B.n370 71.676
R1738 B.n653 B.n371 71.676
R1739 B.n649 B.n372 71.676
R1740 B.n645 B.n373 71.676
R1741 B.n641 B.n374 71.676
R1742 B.n637 B.n375 71.676
R1743 B.n633 B.n376 71.676
R1744 B.n629 B.n377 71.676
R1745 B.n625 B.n378 71.676
R1746 B.n621 B.n379 71.676
R1747 B.n617 B.n380 71.676
R1748 B.n613 B.n381 71.676
R1749 B.n609 B.n382 71.676
R1750 B.n605 B.n383 71.676
R1751 B.n601 B.n384 71.676
R1752 B.n597 B.n385 71.676
R1753 B.n593 B.n386 71.676
R1754 B.n589 B.n387 71.676
R1755 B.n585 B.n388 71.676
R1756 B.n581 B.n389 71.676
R1757 B.n577 B.n390 71.676
R1758 B.n573 B.n391 71.676
R1759 B.n569 B.n392 71.676
R1760 B.n565 B.n393 71.676
R1761 B.n561 B.n394 71.676
R1762 B.n557 B.n395 71.676
R1763 B.n553 B.n396 71.676
R1764 B.n549 B.n397 71.676
R1765 B.n545 B.n398 71.676
R1766 B.n541 B.n399 71.676
R1767 B.n537 B.n400 71.676
R1768 B.n533 B.n401 71.676
R1769 B.n529 B.n402 71.676
R1770 B.n525 B.n403 71.676
R1771 B.n521 B.n404 71.676
R1772 B.n517 B.n405 71.676
R1773 B.n513 B.n406 71.676
R1774 B.n509 B.n407 71.676
R1775 B.n505 B.n408 71.676
R1776 B.n501 B.n409 71.676
R1777 B.n497 B.n410 71.676
R1778 B.n493 B.n411 71.676
R1779 B.n489 B.n412 71.676
R1780 B.n485 B.n413 71.676
R1781 B.n481 B.n414 71.676
R1782 B.n477 B.n415 71.676
R1783 B.n473 B.n416 71.676
R1784 B.n469 B.n417 71.676
R1785 B.n465 B.n418 71.676
R1786 B.n461 B.n419 71.676
R1787 B.n457 B.n420 71.676
R1788 B.n453 B.n421 71.676
R1789 B.n449 B.n422 71.676
R1790 B.n445 B.n423 71.676
R1791 B.n441 B.n424 71.676
R1792 B.n437 B.n425 71.676
R1793 B.n426 B.n366 71.676
R1794 B.n771 B.n770 71.676
R1795 B.n771 B.n2 71.676
R1796 B.n678 B.n363 68.4622
R1797 B.n743 B.n742 68.4622
R1798 B.n209 B.n94 59.5399
R1799 B.n230 B.n92 59.5399
R1800 B.n434 B.n433 59.5399
R1801 B.n431 B.n430 59.5399
R1802 B.n675 B.n361 37.62
R1803 B.n681 B.n680 37.62
R1804 B.n739 B.n738 37.62
R1805 B.n96 B.n25 37.62
R1806 B.n684 B.n363 33.0175
R1807 B.n684 B.n358 33.0175
R1808 B.n690 B.n358 33.0175
R1809 B.n690 B.n359 33.0175
R1810 B.n696 B.n351 33.0175
R1811 B.n702 B.n351 33.0175
R1812 B.n702 B.n347 33.0175
R1813 B.n710 B.n347 33.0175
R1814 B.n710 B.n709 33.0175
R1815 B.n716 B.n4 33.0175
R1816 B.n769 B.n4 33.0175
R1817 B.n769 B.n768 33.0175
R1818 B.n768 B.n767 33.0175
R1819 B.n767 B.n8 33.0175
R1820 B.n760 B.n12 33.0175
R1821 B.n760 B.n759 33.0175
R1822 B.n759 B.n758 33.0175
R1823 B.n758 B.n16 33.0175
R1824 B.n752 B.n16 33.0175
R1825 B.n751 B.n750 33.0175
R1826 B.n750 B.n23 33.0175
R1827 B.n744 B.n23 33.0175
R1828 B.n744 B.n743 33.0175
R1829 B.n94 B.n93 18.6187
R1830 B.n92 B.n91 18.6187
R1831 B.n433 B.n432 18.6187
R1832 B.n430 B.n429 18.6187
R1833 B B.n772 18.0485
R1834 B.n696 B.t7 17.9656
R1835 B.n752 B.t3 17.9656
R1836 B.n716 B.t1 16.9945
R1837 B.t0 B.n8 16.9945
R1838 B.n709 B.t1 16.0235
R1839 B.n12 B.t0 16.0235
R1840 B.n359 B.t7 15.0524
R1841 B.t3 B.n751 15.0524
R1842 B.n686 B.n361 10.6151
R1843 B.n687 B.n686 10.6151
R1844 B.n688 B.n687 10.6151
R1845 B.n688 B.n353 10.6151
R1846 B.n698 B.n353 10.6151
R1847 B.n699 B.n698 10.6151
R1848 B.n700 B.n699 10.6151
R1849 B.n700 B.n345 10.6151
R1850 B.n712 B.n345 10.6151
R1851 B.n713 B.n712 10.6151
R1852 B.n714 B.n713 10.6151
R1853 B.n714 B.n0 10.6151
R1854 B.n675 B.n674 10.6151
R1855 B.n674 B.n673 10.6151
R1856 B.n673 B.n672 10.6151
R1857 B.n672 B.n670 10.6151
R1858 B.n670 B.n667 10.6151
R1859 B.n667 B.n666 10.6151
R1860 B.n666 B.n663 10.6151
R1861 B.n663 B.n662 10.6151
R1862 B.n662 B.n659 10.6151
R1863 B.n659 B.n658 10.6151
R1864 B.n658 B.n655 10.6151
R1865 B.n655 B.n654 10.6151
R1866 B.n654 B.n651 10.6151
R1867 B.n651 B.n650 10.6151
R1868 B.n650 B.n647 10.6151
R1869 B.n647 B.n646 10.6151
R1870 B.n646 B.n643 10.6151
R1871 B.n643 B.n642 10.6151
R1872 B.n642 B.n639 10.6151
R1873 B.n639 B.n638 10.6151
R1874 B.n638 B.n635 10.6151
R1875 B.n635 B.n634 10.6151
R1876 B.n634 B.n631 10.6151
R1877 B.n631 B.n630 10.6151
R1878 B.n630 B.n627 10.6151
R1879 B.n627 B.n626 10.6151
R1880 B.n626 B.n623 10.6151
R1881 B.n623 B.n622 10.6151
R1882 B.n622 B.n619 10.6151
R1883 B.n619 B.n618 10.6151
R1884 B.n618 B.n615 10.6151
R1885 B.n615 B.n614 10.6151
R1886 B.n614 B.n611 10.6151
R1887 B.n611 B.n610 10.6151
R1888 B.n610 B.n607 10.6151
R1889 B.n607 B.n606 10.6151
R1890 B.n606 B.n603 10.6151
R1891 B.n603 B.n602 10.6151
R1892 B.n602 B.n599 10.6151
R1893 B.n599 B.n598 10.6151
R1894 B.n598 B.n595 10.6151
R1895 B.n595 B.n594 10.6151
R1896 B.n594 B.n591 10.6151
R1897 B.n591 B.n590 10.6151
R1898 B.n590 B.n587 10.6151
R1899 B.n587 B.n586 10.6151
R1900 B.n586 B.n583 10.6151
R1901 B.n583 B.n582 10.6151
R1902 B.n582 B.n579 10.6151
R1903 B.n579 B.n578 10.6151
R1904 B.n578 B.n575 10.6151
R1905 B.n575 B.n574 10.6151
R1906 B.n574 B.n571 10.6151
R1907 B.n571 B.n570 10.6151
R1908 B.n570 B.n567 10.6151
R1909 B.n567 B.n566 10.6151
R1910 B.n563 B.n562 10.6151
R1911 B.n562 B.n559 10.6151
R1912 B.n559 B.n558 10.6151
R1913 B.n558 B.n555 10.6151
R1914 B.n555 B.n554 10.6151
R1915 B.n554 B.n551 10.6151
R1916 B.n551 B.n550 10.6151
R1917 B.n550 B.n547 10.6151
R1918 B.n547 B.n546 10.6151
R1919 B.n543 B.n542 10.6151
R1920 B.n542 B.n539 10.6151
R1921 B.n539 B.n538 10.6151
R1922 B.n538 B.n535 10.6151
R1923 B.n535 B.n534 10.6151
R1924 B.n534 B.n531 10.6151
R1925 B.n531 B.n530 10.6151
R1926 B.n530 B.n527 10.6151
R1927 B.n527 B.n526 10.6151
R1928 B.n526 B.n523 10.6151
R1929 B.n523 B.n522 10.6151
R1930 B.n522 B.n519 10.6151
R1931 B.n519 B.n518 10.6151
R1932 B.n518 B.n515 10.6151
R1933 B.n515 B.n514 10.6151
R1934 B.n514 B.n511 10.6151
R1935 B.n511 B.n510 10.6151
R1936 B.n510 B.n507 10.6151
R1937 B.n507 B.n506 10.6151
R1938 B.n506 B.n503 10.6151
R1939 B.n503 B.n502 10.6151
R1940 B.n502 B.n499 10.6151
R1941 B.n499 B.n498 10.6151
R1942 B.n498 B.n495 10.6151
R1943 B.n495 B.n494 10.6151
R1944 B.n494 B.n491 10.6151
R1945 B.n491 B.n490 10.6151
R1946 B.n490 B.n487 10.6151
R1947 B.n487 B.n486 10.6151
R1948 B.n486 B.n483 10.6151
R1949 B.n483 B.n482 10.6151
R1950 B.n482 B.n479 10.6151
R1951 B.n479 B.n478 10.6151
R1952 B.n478 B.n475 10.6151
R1953 B.n475 B.n474 10.6151
R1954 B.n474 B.n471 10.6151
R1955 B.n471 B.n470 10.6151
R1956 B.n470 B.n467 10.6151
R1957 B.n467 B.n466 10.6151
R1958 B.n466 B.n463 10.6151
R1959 B.n463 B.n462 10.6151
R1960 B.n462 B.n459 10.6151
R1961 B.n459 B.n458 10.6151
R1962 B.n458 B.n455 10.6151
R1963 B.n455 B.n454 10.6151
R1964 B.n454 B.n451 10.6151
R1965 B.n451 B.n450 10.6151
R1966 B.n450 B.n447 10.6151
R1967 B.n447 B.n446 10.6151
R1968 B.n446 B.n443 10.6151
R1969 B.n443 B.n442 10.6151
R1970 B.n442 B.n439 10.6151
R1971 B.n439 B.n438 10.6151
R1972 B.n438 B.n435 10.6151
R1973 B.n435 B.n365 10.6151
R1974 B.n680 B.n365 10.6151
R1975 B.n682 B.n681 10.6151
R1976 B.n682 B.n356 10.6151
R1977 B.n692 B.n356 10.6151
R1978 B.n693 B.n692 10.6151
R1979 B.n694 B.n693 10.6151
R1980 B.n694 B.n349 10.6151
R1981 B.n704 B.n349 10.6151
R1982 B.n705 B.n704 10.6151
R1983 B.n707 B.n705 10.6151
R1984 B.n707 B.n706 10.6151
R1985 B.n706 B.n342 10.6151
R1986 B.n719 B.n342 10.6151
R1987 B.n720 B.n719 10.6151
R1988 B.n721 B.n720 10.6151
R1989 B.n722 B.n721 10.6151
R1990 B.n723 B.n722 10.6151
R1991 B.n726 B.n723 10.6151
R1992 B.n727 B.n726 10.6151
R1993 B.n728 B.n727 10.6151
R1994 B.n729 B.n728 10.6151
R1995 B.n731 B.n729 10.6151
R1996 B.n732 B.n731 10.6151
R1997 B.n733 B.n732 10.6151
R1998 B.n734 B.n733 10.6151
R1999 B.n736 B.n734 10.6151
R2000 B.n737 B.n736 10.6151
R2001 B.n738 B.n737 10.6151
R2002 B.n764 B.n1 10.6151
R2003 B.n764 B.n763 10.6151
R2004 B.n763 B.n762 10.6151
R2005 B.n762 B.n10 10.6151
R2006 B.n756 B.n10 10.6151
R2007 B.n756 B.n755 10.6151
R2008 B.n755 B.n754 10.6151
R2009 B.n754 B.n18 10.6151
R2010 B.n748 B.n18 10.6151
R2011 B.n748 B.n747 10.6151
R2012 B.n747 B.n746 10.6151
R2013 B.n746 B.n25 10.6151
R2014 B.n97 B.n96 10.6151
R2015 B.n100 B.n97 10.6151
R2016 B.n101 B.n100 10.6151
R2017 B.n104 B.n101 10.6151
R2018 B.n105 B.n104 10.6151
R2019 B.n108 B.n105 10.6151
R2020 B.n109 B.n108 10.6151
R2021 B.n112 B.n109 10.6151
R2022 B.n113 B.n112 10.6151
R2023 B.n116 B.n113 10.6151
R2024 B.n117 B.n116 10.6151
R2025 B.n120 B.n117 10.6151
R2026 B.n121 B.n120 10.6151
R2027 B.n124 B.n121 10.6151
R2028 B.n125 B.n124 10.6151
R2029 B.n128 B.n125 10.6151
R2030 B.n129 B.n128 10.6151
R2031 B.n132 B.n129 10.6151
R2032 B.n133 B.n132 10.6151
R2033 B.n136 B.n133 10.6151
R2034 B.n137 B.n136 10.6151
R2035 B.n140 B.n137 10.6151
R2036 B.n141 B.n140 10.6151
R2037 B.n144 B.n141 10.6151
R2038 B.n145 B.n144 10.6151
R2039 B.n148 B.n145 10.6151
R2040 B.n149 B.n148 10.6151
R2041 B.n152 B.n149 10.6151
R2042 B.n153 B.n152 10.6151
R2043 B.n156 B.n153 10.6151
R2044 B.n157 B.n156 10.6151
R2045 B.n160 B.n157 10.6151
R2046 B.n161 B.n160 10.6151
R2047 B.n164 B.n161 10.6151
R2048 B.n165 B.n164 10.6151
R2049 B.n168 B.n165 10.6151
R2050 B.n169 B.n168 10.6151
R2051 B.n172 B.n169 10.6151
R2052 B.n173 B.n172 10.6151
R2053 B.n176 B.n173 10.6151
R2054 B.n177 B.n176 10.6151
R2055 B.n180 B.n177 10.6151
R2056 B.n181 B.n180 10.6151
R2057 B.n184 B.n181 10.6151
R2058 B.n185 B.n184 10.6151
R2059 B.n188 B.n185 10.6151
R2060 B.n189 B.n188 10.6151
R2061 B.n192 B.n189 10.6151
R2062 B.n193 B.n192 10.6151
R2063 B.n196 B.n193 10.6151
R2064 B.n197 B.n196 10.6151
R2065 B.n200 B.n197 10.6151
R2066 B.n201 B.n200 10.6151
R2067 B.n204 B.n201 10.6151
R2068 B.n205 B.n204 10.6151
R2069 B.n208 B.n205 10.6151
R2070 B.n213 B.n210 10.6151
R2071 B.n214 B.n213 10.6151
R2072 B.n217 B.n214 10.6151
R2073 B.n218 B.n217 10.6151
R2074 B.n221 B.n218 10.6151
R2075 B.n222 B.n221 10.6151
R2076 B.n225 B.n222 10.6151
R2077 B.n226 B.n225 10.6151
R2078 B.n229 B.n226 10.6151
R2079 B.n234 B.n231 10.6151
R2080 B.n235 B.n234 10.6151
R2081 B.n238 B.n235 10.6151
R2082 B.n239 B.n238 10.6151
R2083 B.n242 B.n239 10.6151
R2084 B.n243 B.n242 10.6151
R2085 B.n246 B.n243 10.6151
R2086 B.n247 B.n246 10.6151
R2087 B.n250 B.n247 10.6151
R2088 B.n251 B.n250 10.6151
R2089 B.n254 B.n251 10.6151
R2090 B.n255 B.n254 10.6151
R2091 B.n258 B.n255 10.6151
R2092 B.n259 B.n258 10.6151
R2093 B.n262 B.n259 10.6151
R2094 B.n263 B.n262 10.6151
R2095 B.n266 B.n263 10.6151
R2096 B.n267 B.n266 10.6151
R2097 B.n270 B.n267 10.6151
R2098 B.n271 B.n270 10.6151
R2099 B.n274 B.n271 10.6151
R2100 B.n275 B.n274 10.6151
R2101 B.n278 B.n275 10.6151
R2102 B.n279 B.n278 10.6151
R2103 B.n282 B.n279 10.6151
R2104 B.n283 B.n282 10.6151
R2105 B.n286 B.n283 10.6151
R2106 B.n287 B.n286 10.6151
R2107 B.n290 B.n287 10.6151
R2108 B.n291 B.n290 10.6151
R2109 B.n294 B.n291 10.6151
R2110 B.n295 B.n294 10.6151
R2111 B.n298 B.n295 10.6151
R2112 B.n299 B.n298 10.6151
R2113 B.n302 B.n299 10.6151
R2114 B.n303 B.n302 10.6151
R2115 B.n306 B.n303 10.6151
R2116 B.n307 B.n306 10.6151
R2117 B.n310 B.n307 10.6151
R2118 B.n311 B.n310 10.6151
R2119 B.n314 B.n311 10.6151
R2120 B.n315 B.n314 10.6151
R2121 B.n318 B.n315 10.6151
R2122 B.n319 B.n318 10.6151
R2123 B.n322 B.n319 10.6151
R2124 B.n323 B.n322 10.6151
R2125 B.n326 B.n323 10.6151
R2126 B.n327 B.n326 10.6151
R2127 B.n330 B.n327 10.6151
R2128 B.n331 B.n330 10.6151
R2129 B.n334 B.n331 10.6151
R2130 B.n335 B.n334 10.6151
R2131 B.n338 B.n335 10.6151
R2132 B.n340 B.n338 10.6151
R2133 B.n341 B.n340 10.6151
R2134 B.n739 B.n341 10.6151
R2135 B.n566 B.n431 8.74196
R2136 B.n543 B.n434 8.74196
R2137 B.n209 B.n208 8.74196
R2138 B.n231 B.n230 8.74196
R2139 B.n772 B.n0 8.11757
R2140 B.n772 B.n1 8.11757
R2141 B.n563 B.n431 1.87367
R2142 B.n546 B.n434 1.87367
R2143 B.n210 B.n209 1.87367
R2144 B.n230 B.n229 1.87367
R2145 VP.n0 VP.t0 931.25
R2146 VP.n0 VP.t1 887.744
R2147 VP VP.n0 0.0516364
R2148 VDD1.n94 VDD1.n93 289.615
R2149 VDD1.n189 VDD1.n188 289.615
R2150 VDD1.n93 VDD1.n92 185
R2151 VDD1.n2 VDD1.n1 185
R2152 VDD1.n87 VDD1.n86 185
R2153 VDD1.n85 VDD1.n84 185
R2154 VDD1.n6 VDD1.n5 185
R2155 VDD1.n79 VDD1.n78 185
R2156 VDD1.n77 VDD1.n76 185
R2157 VDD1.n10 VDD1.n9 185
R2158 VDD1.n71 VDD1.n70 185
R2159 VDD1.n69 VDD1.n68 185
R2160 VDD1.n14 VDD1.n13 185
R2161 VDD1.n63 VDD1.n62 185
R2162 VDD1.n61 VDD1.n60 185
R2163 VDD1.n18 VDD1.n17 185
R2164 VDD1.n55 VDD1.n54 185
R2165 VDD1.n53 VDD1.n20 185
R2166 VDD1.n52 VDD1.n51 185
R2167 VDD1.n23 VDD1.n21 185
R2168 VDD1.n46 VDD1.n45 185
R2169 VDD1.n44 VDD1.n43 185
R2170 VDD1.n27 VDD1.n26 185
R2171 VDD1.n38 VDD1.n37 185
R2172 VDD1.n36 VDD1.n35 185
R2173 VDD1.n31 VDD1.n30 185
R2174 VDD1.n125 VDD1.n124 185
R2175 VDD1.n130 VDD1.n129 185
R2176 VDD1.n132 VDD1.n131 185
R2177 VDD1.n121 VDD1.n120 185
R2178 VDD1.n138 VDD1.n137 185
R2179 VDD1.n140 VDD1.n139 185
R2180 VDD1.n117 VDD1.n116 185
R2181 VDD1.n147 VDD1.n146 185
R2182 VDD1.n148 VDD1.n115 185
R2183 VDD1.n150 VDD1.n149 185
R2184 VDD1.n113 VDD1.n112 185
R2185 VDD1.n156 VDD1.n155 185
R2186 VDD1.n158 VDD1.n157 185
R2187 VDD1.n109 VDD1.n108 185
R2188 VDD1.n164 VDD1.n163 185
R2189 VDD1.n166 VDD1.n165 185
R2190 VDD1.n105 VDD1.n104 185
R2191 VDD1.n172 VDD1.n171 185
R2192 VDD1.n174 VDD1.n173 185
R2193 VDD1.n101 VDD1.n100 185
R2194 VDD1.n180 VDD1.n179 185
R2195 VDD1.n182 VDD1.n181 185
R2196 VDD1.n97 VDD1.n96 185
R2197 VDD1.n188 VDD1.n187 185
R2198 VDD1.n32 VDD1.t1 149.524
R2199 VDD1.n126 VDD1.t0 149.524
R2200 VDD1.n93 VDD1.n1 104.615
R2201 VDD1.n86 VDD1.n1 104.615
R2202 VDD1.n86 VDD1.n85 104.615
R2203 VDD1.n85 VDD1.n5 104.615
R2204 VDD1.n78 VDD1.n5 104.615
R2205 VDD1.n78 VDD1.n77 104.615
R2206 VDD1.n77 VDD1.n9 104.615
R2207 VDD1.n70 VDD1.n9 104.615
R2208 VDD1.n70 VDD1.n69 104.615
R2209 VDD1.n69 VDD1.n13 104.615
R2210 VDD1.n62 VDD1.n13 104.615
R2211 VDD1.n62 VDD1.n61 104.615
R2212 VDD1.n61 VDD1.n17 104.615
R2213 VDD1.n54 VDD1.n17 104.615
R2214 VDD1.n54 VDD1.n53 104.615
R2215 VDD1.n53 VDD1.n52 104.615
R2216 VDD1.n52 VDD1.n21 104.615
R2217 VDD1.n45 VDD1.n21 104.615
R2218 VDD1.n45 VDD1.n44 104.615
R2219 VDD1.n44 VDD1.n26 104.615
R2220 VDD1.n37 VDD1.n26 104.615
R2221 VDD1.n37 VDD1.n36 104.615
R2222 VDD1.n36 VDD1.n30 104.615
R2223 VDD1.n130 VDD1.n124 104.615
R2224 VDD1.n131 VDD1.n130 104.615
R2225 VDD1.n131 VDD1.n120 104.615
R2226 VDD1.n138 VDD1.n120 104.615
R2227 VDD1.n139 VDD1.n138 104.615
R2228 VDD1.n139 VDD1.n116 104.615
R2229 VDD1.n147 VDD1.n116 104.615
R2230 VDD1.n148 VDD1.n147 104.615
R2231 VDD1.n149 VDD1.n148 104.615
R2232 VDD1.n149 VDD1.n112 104.615
R2233 VDD1.n156 VDD1.n112 104.615
R2234 VDD1.n157 VDD1.n156 104.615
R2235 VDD1.n157 VDD1.n108 104.615
R2236 VDD1.n164 VDD1.n108 104.615
R2237 VDD1.n165 VDD1.n164 104.615
R2238 VDD1.n165 VDD1.n104 104.615
R2239 VDD1.n172 VDD1.n104 104.615
R2240 VDD1.n173 VDD1.n172 104.615
R2241 VDD1.n173 VDD1.n100 104.615
R2242 VDD1.n180 VDD1.n100 104.615
R2243 VDD1.n181 VDD1.n180 104.615
R2244 VDD1.n181 VDD1.n96 104.615
R2245 VDD1.n188 VDD1.n96 104.615
R2246 VDD1 VDD1.n189 91.8326
R2247 VDD1.t1 VDD1.n30 52.3082
R2248 VDD1.t0 VDD1.n124 52.3082
R2249 VDD1 VDD1.n94 51.0686
R2250 VDD1.n55 VDD1.n20 13.1884
R2251 VDD1.n150 VDD1.n115 13.1884
R2252 VDD1.n56 VDD1.n18 12.8005
R2253 VDD1.n51 VDD1.n22 12.8005
R2254 VDD1.n146 VDD1.n145 12.8005
R2255 VDD1.n151 VDD1.n113 12.8005
R2256 VDD1.n60 VDD1.n59 12.0247
R2257 VDD1.n50 VDD1.n23 12.0247
R2258 VDD1.n144 VDD1.n117 12.0247
R2259 VDD1.n155 VDD1.n154 12.0247
R2260 VDD1.n92 VDD1.n0 11.249
R2261 VDD1.n63 VDD1.n16 11.249
R2262 VDD1.n47 VDD1.n46 11.249
R2263 VDD1.n141 VDD1.n140 11.249
R2264 VDD1.n158 VDD1.n111 11.249
R2265 VDD1.n187 VDD1.n95 11.249
R2266 VDD1.n91 VDD1.n2 10.4732
R2267 VDD1.n64 VDD1.n14 10.4732
R2268 VDD1.n43 VDD1.n25 10.4732
R2269 VDD1.n137 VDD1.n119 10.4732
R2270 VDD1.n159 VDD1.n109 10.4732
R2271 VDD1.n186 VDD1.n97 10.4732
R2272 VDD1.n32 VDD1.n31 10.2747
R2273 VDD1.n126 VDD1.n125 10.2747
R2274 VDD1.n88 VDD1.n87 9.69747
R2275 VDD1.n68 VDD1.n67 9.69747
R2276 VDD1.n42 VDD1.n27 9.69747
R2277 VDD1.n136 VDD1.n121 9.69747
R2278 VDD1.n163 VDD1.n162 9.69747
R2279 VDD1.n183 VDD1.n182 9.69747
R2280 VDD1.n90 VDD1.n0 9.45567
R2281 VDD1.n185 VDD1.n95 9.45567
R2282 VDD1.n91 VDD1.n90 9.3005
R2283 VDD1.n89 VDD1.n88 9.3005
R2284 VDD1.n4 VDD1.n3 9.3005
R2285 VDD1.n83 VDD1.n82 9.3005
R2286 VDD1.n81 VDD1.n80 9.3005
R2287 VDD1.n8 VDD1.n7 9.3005
R2288 VDD1.n75 VDD1.n74 9.3005
R2289 VDD1.n73 VDD1.n72 9.3005
R2290 VDD1.n12 VDD1.n11 9.3005
R2291 VDD1.n67 VDD1.n66 9.3005
R2292 VDD1.n65 VDD1.n64 9.3005
R2293 VDD1.n16 VDD1.n15 9.3005
R2294 VDD1.n59 VDD1.n58 9.3005
R2295 VDD1.n57 VDD1.n56 9.3005
R2296 VDD1.n22 VDD1.n19 9.3005
R2297 VDD1.n50 VDD1.n49 9.3005
R2298 VDD1.n48 VDD1.n47 9.3005
R2299 VDD1.n25 VDD1.n24 9.3005
R2300 VDD1.n42 VDD1.n41 9.3005
R2301 VDD1.n40 VDD1.n39 9.3005
R2302 VDD1.n29 VDD1.n28 9.3005
R2303 VDD1.n34 VDD1.n33 9.3005
R2304 VDD1.n103 VDD1.n102 9.3005
R2305 VDD1.n176 VDD1.n175 9.3005
R2306 VDD1.n178 VDD1.n177 9.3005
R2307 VDD1.n99 VDD1.n98 9.3005
R2308 VDD1.n184 VDD1.n183 9.3005
R2309 VDD1.n186 VDD1.n185 9.3005
R2310 VDD1.n168 VDD1.n167 9.3005
R2311 VDD1.n107 VDD1.n106 9.3005
R2312 VDD1.n162 VDD1.n161 9.3005
R2313 VDD1.n160 VDD1.n159 9.3005
R2314 VDD1.n111 VDD1.n110 9.3005
R2315 VDD1.n154 VDD1.n153 9.3005
R2316 VDD1.n152 VDD1.n151 9.3005
R2317 VDD1.n128 VDD1.n127 9.3005
R2318 VDD1.n123 VDD1.n122 9.3005
R2319 VDD1.n134 VDD1.n133 9.3005
R2320 VDD1.n136 VDD1.n135 9.3005
R2321 VDD1.n119 VDD1.n118 9.3005
R2322 VDD1.n142 VDD1.n141 9.3005
R2323 VDD1.n144 VDD1.n143 9.3005
R2324 VDD1.n145 VDD1.n114 9.3005
R2325 VDD1.n170 VDD1.n169 9.3005
R2326 VDD1.n84 VDD1.n4 8.92171
R2327 VDD1.n71 VDD1.n12 8.92171
R2328 VDD1.n39 VDD1.n38 8.92171
R2329 VDD1.n133 VDD1.n132 8.92171
R2330 VDD1.n166 VDD1.n107 8.92171
R2331 VDD1.n179 VDD1.n99 8.92171
R2332 VDD1.n83 VDD1.n6 8.14595
R2333 VDD1.n72 VDD1.n10 8.14595
R2334 VDD1.n35 VDD1.n29 8.14595
R2335 VDD1.n129 VDD1.n123 8.14595
R2336 VDD1.n167 VDD1.n105 8.14595
R2337 VDD1.n178 VDD1.n101 8.14595
R2338 VDD1.n80 VDD1.n79 7.3702
R2339 VDD1.n76 VDD1.n75 7.3702
R2340 VDD1.n34 VDD1.n31 7.3702
R2341 VDD1.n128 VDD1.n125 7.3702
R2342 VDD1.n171 VDD1.n170 7.3702
R2343 VDD1.n175 VDD1.n174 7.3702
R2344 VDD1.n79 VDD1.n8 6.59444
R2345 VDD1.n76 VDD1.n8 6.59444
R2346 VDD1.n171 VDD1.n103 6.59444
R2347 VDD1.n174 VDD1.n103 6.59444
R2348 VDD1.n80 VDD1.n6 5.81868
R2349 VDD1.n75 VDD1.n10 5.81868
R2350 VDD1.n35 VDD1.n34 5.81868
R2351 VDD1.n129 VDD1.n128 5.81868
R2352 VDD1.n170 VDD1.n105 5.81868
R2353 VDD1.n175 VDD1.n101 5.81868
R2354 VDD1.n84 VDD1.n83 5.04292
R2355 VDD1.n72 VDD1.n71 5.04292
R2356 VDD1.n38 VDD1.n29 5.04292
R2357 VDD1.n132 VDD1.n123 5.04292
R2358 VDD1.n167 VDD1.n166 5.04292
R2359 VDD1.n179 VDD1.n178 5.04292
R2360 VDD1.n87 VDD1.n4 4.26717
R2361 VDD1.n68 VDD1.n12 4.26717
R2362 VDD1.n39 VDD1.n27 4.26717
R2363 VDD1.n133 VDD1.n121 4.26717
R2364 VDD1.n163 VDD1.n107 4.26717
R2365 VDD1.n182 VDD1.n99 4.26717
R2366 VDD1.n88 VDD1.n2 3.49141
R2367 VDD1.n67 VDD1.n14 3.49141
R2368 VDD1.n43 VDD1.n42 3.49141
R2369 VDD1.n137 VDD1.n136 3.49141
R2370 VDD1.n162 VDD1.n109 3.49141
R2371 VDD1.n183 VDD1.n97 3.49141
R2372 VDD1.n33 VDD1.n32 2.84303
R2373 VDD1.n127 VDD1.n126 2.84303
R2374 VDD1.n92 VDD1.n91 2.71565
R2375 VDD1.n64 VDD1.n63 2.71565
R2376 VDD1.n46 VDD1.n25 2.71565
R2377 VDD1.n140 VDD1.n119 2.71565
R2378 VDD1.n159 VDD1.n158 2.71565
R2379 VDD1.n187 VDD1.n186 2.71565
R2380 VDD1.n94 VDD1.n0 1.93989
R2381 VDD1.n60 VDD1.n16 1.93989
R2382 VDD1.n47 VDD1.n23 1.93989
R2383 VDD1.n141 VDD1.n117 1.93989
R2384 VDD1.n155 VDD1.n111 1.93989
R2385 VDD1.n189 VDD1.n95 1.93989
R2386 VDD1.n59 VDD1.n18 1.16414
R2387 VDD1.n51 VDD1.n50 1.16414
R2388 VDD1.n146 VDD1.n144 1.16414
R2389 VDD1.n154 VDD1.n113 1.16414
R2390 VDD1.n56 VDD1.n55 0.388379
R2391 VDD1.n22 VDD1.n20 0.388379
R2392 VDD1.n145 VDD1.n115 0.388379
R2393 VDD1.n151 VDD1.n150 0.388379
R2394 VDD1.n90 VDD1.n89 0.155672
R2395 VDD1.n89 VDD1.n3 0.155672
R2396 VDD1.n82 VDD1.n3 0.155672
R2397 VDD1.n82 VDD1.n81 0.155672
R2398 VDD1.n81 VDD1.n7 0.155672
R2399 VDD1.n74 VDD1.n7 0.155672
R2400 VDD1.n74 VDD1.n73 0.155672
R2401 VDD1.n73 VDD1.n11 0.155672
R2402 VDD1.n66 VDD1.n11 0.155672
R2403 VDD1.n66 VDD1.n65 0.155672
R2404 VDD1.n65 VDD1.n15 0.155672
R2405 VDD1.n58 VDD1.n15 0.155672
R2406 VDD1.n58 VDD1.n57 0.155672
R2407 VDD1.n57 VDD1.n19 0.155672
R2408 VDD1.n49 VDD1.n19 0.155672
R2409 VDD1.n49 VDD1.n48 0.155672
R2410 VDD1.n48 VDD1.n24 0.155672
R2411 VDD1.n41 VDD1.n24 0.155672
R2412 VDD1.n41 VDD1.n40 0.155672
R2413 VDD1.n40 VDD1.n28 0.155672
R2414 VDD1.n33 VDD1.n28 0.155672
R2415 VDD1.n127 VDD1.n122 0.155672
R2416 VDD1.n134 VDD1.n122 0.155672
R2417 VDD1.n135 VDD1.n134 0.155672
R2418 VDD1.n135 VDD1.n118 0.155672
R2419 VDD1.n142 VDD1.n118 0.155672
R2420 VDD1.n143 VDD1.n142 0.155672
R2421 VDD1.n143 VDD1.n114 0.155672
R2422 VDD1.n152 VDD1.n114 0.155672
R2423 VDD1.n153 VDD1.n152 0.155672
R2424 VDD1.n153 VDD1.n110 0.155672
R2425 VDD1.n160 VDD1.n110 0.155672
R2426 VDD1.n161 VDD1.n160 0.155672
R2427 VDD1.n161 VDD1.n106 0.155672
R2428 VDD1.n168 VDD1.n106 0.155672
R2429 VDD1.n169 VDD1.n168 0.155672
R2430 VDD1.n169 VDD1.n102 0.155672
R2431 VDD1.n176 VDD1.n102 0.155672
R2432 VDD1.n177 VDD1.n176 0.155672
R2433 VDD1.n177 VDD1.n98 0.155672
R2434 VDD1.n184 VDD1.n98 0.155672
R2435 VDD1.n185 VDD1.n184 0.155672
C0 VN VDD2 2.66123f
C1 VDD1 VDD2 0.457065f
C2 VP VDD2 0.253265f
C3 VTAIL VDD2 7.8596f
C4 VN VDD1 0.14889f
C5 VN VP 5.52065f
C6 VN VTAIL 1.90133f
C7 VP VDD1 2.75923f
C8 VTAIL VDD1 7.82962f
C9 VTAIL VP 1.91619f
C10 VDD2 B 4.695606f
C11 VDD1 B 7.60832f
C12 VTAIL B 8.394836f
C13 VN B 9.370231f
C14 VP B 4.310434f
C15 VDD1.n0 B 0.011893f
C16 VDD1.n1 B 0.026792f
C17 VDD1.n2 B 0.012002f
C18 VDD1.n3 B 0.021095f
C19 VDD1.n4 B 0.011335f
C20 VDD1.n5 B 0.026792f
C21 VDD1.n6 B 0.012002f
C22 VDD1.n7 B 0.021095f
C23 VDD1.n8 B 0.011335f
C24 VDD1.n9 B 0.026792f
C25 VDD1.n10 B 0.012002f
C26 VDD1.n11 B 0.021095f
C27 VDD1.n12 B 0.011335f
C28 VDD1.n13 B 0.026792f
C29 VDD1.n14 B 0.012002f
C30 VDD1.n15 B 0.021095f
C31 VDD1.n16 B 0.011335f
C32 VDD1.n17 B 0.026792f
C33 VDD1.n18 B 0.012002f
C34 VDD1.n19 B 0.021095f
C35 VDD1.n20 B 0.011669f
C36 VDD1.n21 B 0.026792f
C37 VDD1.n22 B 0.011335f
C38 VDD1.n23 B 0.012002f
C39 VDD1.n24 B 0.021095f
C40 VDD1.n25 B 0.011335f
C41 VDD1.n26 B 0.026792f
C42 VDD1.n27 B 0.012002f
C43 VDD1.n28 B 0.021095f
C44 VDD1.n29 B 0.011335f
C45 VDD1.n30 B 0.020094f
C46 VDD1.n31 B 0.01894f
C47 VDD1.t1 B 0.04586f
C48 VDD1.n32 B 0.195498f
C49 VDD1.n33 B 1.56709f
C50 VDD1.n34 B 0.011335f
C51 VDD1.n35 B 0.012002f
C52 VDD1.n36 B 0.026792f
C53 VDD1.n37 B 0.026792f
C54 VDD1.n38 B 0.012002f
C55 VDD1.n39 B 0.011335f
C56 VDD1.n40 B 0.021095f
C57 VDD1.n41 B 0.021095f
C58 VDD1.n42 B 0.011335f
C59 VDD1.n43 B 0.012002f
C60 VDD1.n44 B 0.026792f
C61 VDD1.n45 B 0.026792f
C62 VDD1.n46 B 0.012002f
C63 VDD1.n47 B 0.011335f
C64 VDD1.n48 B 0.021095f
C65 VDD1.n49 B 0.021095f
C66 VDD1.n50 B 0.011335f
C67 VDD1.n51 B 0.012002f
C68 VDD1.n52 B 0.026792f
C69 VDD1.n53 B 0.026792f
C70 VDD1.n54 B 0.026792f
C71 VDD1.n55 B 0.011669f
C72 VDD1.n56 B 0.011335f
C73 VDD1.n57 B 0.021095f
C74 VDD1.n58 B 0.021095f
C75 VDD1.n59 B 0.011335f
C76 VDD1.n60 B 0.012002f
C77 VDD1.n61 B 0.026792f
C78 VDD1.n62 B 0.026792f
C79 VDD1.n63 B 0.012002f
C80 VDD1.n64 B 0.011335f
C81 VDD1.n65 B 0.021095f
C82 VDD1.n66 B 0.021095f
C83 VDD1.n67 B 0.011335f
C84 VDD1.n68 B 0.012002f
C85 VDD1.n69 B 0.026792f
C86 VDD1.n70 B 0.026792f
C87 VDD1.n71 B 0.012002f
C88 VDD1.n72 B 0.011335f
C89 VDD1.n73 B 0.021095f
C90 VDD1.n74 B 0.021095f
C91 VDD1.n75 B 0.011335f
C92 VDD1.n76 B 0.012002f
C93 VDD1.n77 B 0.026792f
C94 VDD1.n78 B 0.026792f
C95 VDD1.n79 B 0.012002f
C96 VDD1.n80 B 0.011335f
C97 VDD1.n81 B 0.021095f
C98 VDD1.n82 B 0.021095f
C99 VDD1.n83 B 0.011335f
C100 VDD1.n84 B 0.012002f
C101 VDD1.n85 B 0.026792f
C102 VDD1.n86 B 0.026792f
C103 VDD1.n87 B 0.012002f
C104 VDD1.n88 B 0.011335f
C105 VDD1.n89 B 0.021095f
C106 VDD1.n90 B 0.054522f
C107 VDD1.n91 B 0.011335f
C108 VDD1.n92 B 0.012002f
C109 VDD1.n93 B 0.052968f
C110 VDD1.n94 B 0.060022f
C111 VDD1.n95 B 0.011893f
C112 VDD1.n96 B 0.026792f
C113 VDD1.n97 B 0.012002f
C114 VDD1.n98 B 0.021095f
C115 VDD1.n99 B 0.011335f
C116 VDD1.n100 B 0.026792f
C117 VDD1.n101 B 0.012002f
C118 VDD1.n102 B 0.021095f
C119 VDD1.n103 B 0.011335f
C120 VDD1.n104 B 0.026792f
C121 VDD1.n105 B 0.012002f
C122 VDD1.n106 B 0.021095f
C123 VDD1.n107 B 0.011335f
C124 VDD1.n108 B 0.026792f
C125 VDD1.n109 B 0.012002f
C126 VDD1.n110 B 0.021095f
C127 VDD1.n111 B 0.011335f
C128 VDD1.n112 B 0.026792f
C129 VDD1.n113 B 0.012002f
C130 VDD1.n114 B 0.021095f
C131 VDD1.n115 B 0.011669f
C132 VDD1.n116 B 0.026792f
C133 VDD1.n117 B 0.012002f
C134 VDD1.n118 B 0.021095f
C135 VDD1.n119 B 0.011335f
C136 VDD1.n120 B 0.026792f
C137 VDD1.n121 B 0.012002f
C138 VDD1.n122 B 0.021095f
C139 VDD1.n123 B 0.011335f
C140 VDD1.n124 B 0.020094f
C141 VDD1.n125 B 0.01894f
C142 VDD1.t0 B 0.04586f
C143 VDD1.n126 B 0.195498f
C144 VDD1.n127 B 1.56709f
C145 VDD1.n128 B 0.011335f
C146 VDD1.n129 B 0.012002f
C147 VDD1.n130 B 0.026792f
C148 VDD1.n131 B 0.026792f
C149 VDD1.n132 B 0.012002f
C150 VDD1.n133 B 0.011335f
C151 VDD1.n134 B 0.021095f
C152 VDD1.n135 B 0.021095f
C153 VDD1.n136 B 0.011335f
C154 VDD1.n137 B 0.012002f
C155 VDD1.n138 B 0.026792f
C156 VDD1.n139 B 0.026792f
C157 VDD1.n140 B 0.012002f
C158 VDD1.n141 B 0.011335f
C159 VDD1.n142 B 0.021095f
C160 VDD1.n143 B 0.021095f
C161 VDD1.n144 B 0.011335f
C162 VDD1.n145 B 0.011335f
C163 VDD1.n146 B 0.012002f
C164 VDD1.n147 B 0.026792f
C165 VDD1.n148 B 0.026792f
C166 VDD1.n149 B 0.026792f
C167 VDD1.n150 B 0.011669f
C168 VDD1.n151 B 0.011335f
C169 VDD1.n152 B 0.021095f
C170 VDD1.n153 B 0.021095f
C171 VDD1.n154 B 0.011335f
C172 VDD1.n155 B 0.012002f
C173 VDD1.n156 B 0.026792f
C174 VDD1.n157 B 0.026792f
C175 VDD1.n158 B 0.012002f
C176 VDD1.n159 B 0.011335f
C177 VDD1.n160 B 0.021095f
C178 VDD1.n161 B 0.021095f
C179 VDD1.n162 B 0.011335f
C180 VDD1.n163 B 0.012002f
C181 VDD1.n164 B 0.026792f
C182 VDD1.n165 B 0.026792f
C183 VDD1.n166 B 0.012002f
C184 VDD1.n167 B 0.011335f
C185 VDD1.n168 B 0.021095f
C186 VDD1.n169 B 0.021095f
C187 VDD1.n170 B 0.011335f
C188 VDD1.n171 B 0.012002f
C189 VDD1.n172 B 0.026792f
C190 VDD1.n173 B 0.026792f
C191 VDD1.n174 B 0.012002f
C192 VDD1.n175 B 0.011335f
C193 VDD1.n176 B 0.021095f
C194 VDD1.n177 B 0.021095f
C195 VDD1.n178 B 0.011335f
C196 VDD1.n179 B 0.012002f
C197 VDD1.n180 B 0.026792f
C198 VDD1.n181 B 0.026792f
C199 VDD1.n182 B 0.012002f
C200 VDD1.n183 B 0.011335f
C201 VDD1.n184 B 0.021095f
C202 VDD1.n185 B 0.054522f
C203 VDD1.n186 B 0.011335f
C204 VDD1.n187 B 0.012002f
C205 VDD1.n188 B 0.052968f
C206 VDD1.n189 B 0.703295f
C207 VP.t0 B 1.70192f
C208 VP.t1 B 1.58292f
C209 VP.n0 B 5.00058f
C210 VDD2.n0 B 0.011981f
C211 VDD2.n1 B 0.026991f
C212 VDD2.n2 B 0.012091f
C213 VDD2.n3 B 0.021251f
C214 VDD2.n4 B 0.011419f
C215 VDD2.n5 B 0.026991f
C216 VDD2.n6 B 0.012091f
C217 VDD2.n7 B 0.021251f
C218 VDD2.n8 B 0.011419f
C219 VDD2.n9 B 0.026991f
C220 VDD2.n10 B 0.012091f
C221 VDD2.n11 B 0.021251f
C222 VDD2.n12 B 0.011419f
C223 VDD2.n13 B 0.026991f
C224 VDD2.n14 B 0.012091f
C225 VDD2.n15 B 0.021251f
C226 VDD2.n16 B 0.011419f
C227 VDD2.n17 B 0.026991f
C228 VDD2.n18 B 0.012091f
C229 VDD2.n19 B 0.021251f
C230 VDD2.n20 B 0.011755f
C231 VDD2.n21 B 0.026991f
C232 VDD2.n22 B 0.012091f
C233 VDD2.n23 B 0.021251f
C234 VDD2.n24 B 0.011419f
C235 VDD2.n25 B 0.026991f
C236 VDD2.n26 B 0.012091f
C237 VDD2.n27 B 0.021251f
C238 VDD2.n28 B 0.011419f
C239 VDD2.n29 B 0.020243f
C240 VDD2.n30 B 0.01908f
C241 VDD2.t0 B 0.046199f
C242 VDD2.n31 B 0.196945f
C243 VDD2.n32 B 1.57869f
C244 VDD2.n33 B 0.011419f
C245 VDD2.n34 B 0.012091f
C246 VDD2.n35 B 0.026991f
C247 VDD2.n36 B 0.026991f
C248 VDD2.n37 B 0.012091f
C249 VDD2.n38 B 0.011419f
C250 VDD2.n39 B 0.021251f
C251 VDD2.n40 B 0.021251f
C252 VDD2.n41 B 0.011419f
C253 VDD2.n42 B 0.012091f
C254 VDD2.n43 B 0.026991f
C255 VDD2.n44 B 0.026991f
C256 VDD2.n45 B 0.012091f
C257 VDD2.n46 B 0.011419f
C258 VDD2.n47 B 0.021251f
C259 VDD2.n48 B 0.021251f
C260 VDD2.n49 B 0.011419f
C261 VDD2.n50 B 0.011419f
C262 VDD2.n51 B 0.012091f
C263 VDD2.n52 B 0.026991f
C264 VDD2.n53 B 0.026991f
C265 VDD2.n54 B 0.026991f
C266 VDD2.n55 B 0.011755f
C267 VDD2.n56 B 0.011419f
C268 VDD2.n57 B 0.021251f
C269 VDD2.n58 B 0.021251f
C270 VDD2.n59 B 0.011419f
C271 VDD2.n60 B 0.012091f
C272 VDD2.n61 B 0.026991f
C273 VDD2.n62 B 0.026991f
C274 VDD2.n63 B 0.012091f
C275 VDD2.n64 B 0.011419f
C276 VDD2.n65 B 0.021251f
C277 VDD2.n66 B 0.021251f
C278 VDD2.n67 B 0.011419f
C279 VDD2.n68 B 0.012091f
C280 VDD2.n69 B 0.026991f
C281 VDD2.n70 B 0.026991f
C282 VDD2.n71 B 0.012091f
C283 VDD2.n72 B 0.011419f
C284 VDD2.n73 B 0.021251f
C285 VDD2.n74 B 0.021251f
C286 VDD2.n75 B 0.011419f
C287 VDD2.n76 B 0.012091f
C288 VDD2.n77 B 0.026991f
C289 VDD2.n78 B 0.026991f
C290 VDD2.n79 B 0.012091f
C291 VDD2.n80 B 0.011419f
C292 VDD2.n81 B 0.021251f
C293 VDD2.n82 B 0.021251f
C294 VDD2.n83 B 0.011419f
C295 VDD2.n84 B 0.012091f
C296 VDD2.n85 B 0.026991f
C297 VDD2.n86 B 0.026991f
C298 VDD2.n87 B 0.012091f
C299 VDD2.n88 B 0.011419f
C300 VDD2.n89 B 0.021251f
C301 VDD2.n90 B 0.054926f
C302 VDD2.n91 B 0.011419f
C303 VDD2.n92 B 0.012091f
C304 VDD2.n93 B 0.05336f
C305 VDD2.n94 B 0.678795f
C306 VDD2.n95 B 0.011981f
C307 VDD2.n96 B 0.026991f
C308 VDD2.n97 B 0.012091f
C309 VDD2.n98 B 0.021251f
C310 VDD2.n99 B 0.011419f
C311 VDD2.n100 B 0.026991f
C312 VDD2.n101 B 0.012091f
C313 VDD2.n102 B 0.021251f
C314 VDD2.n103 B 0.011419f
C315 VDD2.n104 B 0.026991f
C316 VDD2.n105 B 0.012091f
C317 VDD2.n106 B 0.021251f
C318 VDD2.n107 B 0.011419f
C319 VDD2.n108 B 0.026991f
C320 VDD2.n109 B 0.012091f
C321 VDD2.n110 B 0.021251f
C322 VDD2.n111 B 0.011419f
C323 VDD2.n112 B 0.026991f
C324 VDD2.n113 B 0.012091f
C325 VDD2.n114 B 0.021251f
C326 VDD2.n115 B 0.011755f
C327 VDD2.n116 B 0.026991f
C328 VDD2.n117 B 0.011419f
C329 VDD2.n118 B 0.012091f
C330 VDD2.n119 B 0.021251f
C331 VDD2.n120 B 0.011419f
C332 VDD2.n121 B 0.026991f
C333 VDD2.n122 B 0.012091f
C334 VDD2.n123 B 0.021251f
C335 VDD2.n124 B 0.011419f
C336 VDD2.n125 B 0.020243f
C337 VDD2.n126 B 0.01908f
C338 VDD2.t1 B 0.046199f
C339 VDD2.n127 B 0.196945f
C340 VDD2.n128 B 1.57869f
C341 VDD2.n129 B 0.011419f
C342 VDD2.n130 B 0.012091f
C343 VDD2.n131 B 0.026991f
C344 VDD2.n132 B 0.026991f
C345 VDD2.n133 B 0.012091f
C346 VDD2.n134 B 0.011419f
C347 VDD2.n135 B 0.021251f
C348 VDD2.n136 B 0.021251f
C349 VDD2.n137 B 0.011419f
C350 VDD2.n138 B 0.012091f
C351 VDD2.n139 B 0.026991f
C352 VDD2.n140 B 0.026991f
C353 VDD2.n141 B 0.012091f
C354 VDD2.n142 B 0.011419f
C355 VDD2.n143 B 0.021251f
C356 VDD2.n144 B 0.021251f
C357 VDD2.n145 B 0.011419f
C358 VDD2.n146 B 0.012091f
C359 VDD2.n147 B 0.026991f
C360 VDD2.n148 B 0.026991f
C361 VDD2.n149 B 0.026991f
C362 VDD2.n150 B 0.011755f
C363 VDD2.n151 B 0.011419f
C364 VDD2.n152 B 0.021251f
C365 VDD2.n153 B 0.021251f
C366 VDD2.n154 B 0.011419f
C367 VDD2.n155 B 0.012091f
C368 VDD2.n156 B 0.026991f
C369 VDD2.n157 B 0.026991f
C370 VDD2.n158 B 0.012091f
C371 VDD2.n159 B 0.011419f
C372 VDD2.n160 B 0.021251f
C373 VDD2.n161 B 0.021251f
C374 VDD2.n162 B 0.011419f
C375 VDD2.n163 B 0.012091f
C376 VDD2.n164 B 0.026991f
C377 VDD2.n165 B 0.026991f
C378 VDD2.n166 B 0.012091f
C379 VDD2.n167 B 0.011419f
C380 VDD2.n168 B 0.021251f
C381 VDD2.n169 B 0.021251f
C382 VDD2.n170 B 0.011419f
C383 VDD2.n171 B 0.012091f
C384 VDD2.n172 B 0.026991f
C385 VDD2.n173 B 0.026991f
C386 VDD2.n174 B 0.012091f
C387 VDD2.n175 B 0.011419f
C388 VDD2.n176 B 0.021251f
C389 VDD2.n177 B 0.021251f
C390 VDD2.n178 B 0.011419f
C391 VDD2.n179 B 0.012091f
C392 VDD2.n180 B 0.026991f
C393 VDD2.n181 B 0.026991f
C394 VDD2.n182 B 0.012091f
C395 VDD2.n183 B 0.011419f
C396 VDD2.n184 B 0.021251f
C397 VDD2.n185 B 0.054926f
C398 VDD2.n186 B 0.011419f
C399 VDD2.n187 B 0.012091f
C400 VDD2.n188 B 0.05336f
C401 VDD2.n189 B 0.060151f
C402 VDD2.n190 B 2.7562f
C403 VTAIL.n0 B 0.009304f
C404 VTAIL.n1 B 0.02096f
C405 VTAIL.n2 B 0.009389f
C406 VTAIL.n3 B 0.016503f
C407 VTAIL.n4 B 0.008868f
C408 VTAIL.n5 B 0.02096f
C409 VTAIL.n6 B 0.009389f
C410 VTAIL.n7 B 0.016503f
C411 VTAIL.n8 B 0.008868f
C412 VTAIL.n9 B 0.02096f
C413 VTAIL.n10 B 0.009389f
C414 VTAIL.n11 B 0.016503f
C415 VTAIL.n12 B 0.008868f
C416 VTAIL.n13 B 0.02096f
C417 VTAIL.n14 B 0.009389f
C418 VTAIL.n15 B 0.016503f
C419 VTAIL.n16 B 0.008868f
C420 VTAIL.n17 B 0.02096f
C421 VTAIL.n18 B 0.009389f
C422 VTAIL.n19 B 0.016503f
C423 VTAIL.n20 B 0.009129f
C424 VTAIL.n21 B 0.02096f
C425 VTAIL.n22 B 0.009389f
C426 VTAIL.n23 B 0.016503f
C427 VTAIL.n24 B 0.008868f
C428 VTAIL.n25 B 0.02096f
C429 VTAIL.n26 B 0.009389f
C430 VTAIL.n27 B 0.016503f
C431 VTAIL.n28 B 0.008868f
C432 VTAIL.n29 B 0.01572f
C433 VTAIL.n30 B 0.014817f
C434 VTAIL.t1 B 0.035877f
C435 VTAIL.n31 B 0.152941f
C436 VTAIL.n32 B 1.22596f
C437 VTAIL.n33 B 0.008868f
C438 VTAIL.n34 B 0.009389f
C439 VTAIL.n35 B 0.02096f
C440 VTAIL.n36 B 0.02096f
C441 VTAIL.n37 B 0.009389f
C442 VTAIL.n38 B 0.008868f
C443 VTAIL.n39 B 0.016503f
C444 VTAIL.n40 B 0.016503f
C445 VTAIL.n41 B 0.008868f
C446 VTAIL.n42 B 0.009389f
C447 VTAIL.n43 B 0.02096f
C448 VTAIL.n44 B 0.02096f
C449 VTAIL.n45 B 0.009389f
C450 VTAIL.n46 B 0.008868f
C451 VTAIL.n47 B 0.016503f
C452 VTAIL.n48 B 0.016503f
C453 VTAIL.n49 B 0.008868f
C454 VTAIL.n50 B 0.008868f
C455 VTAIL.n51 B 0.009389f
C456 VTAIL.n52 B 0.02096f
C457 VTAIL.n53 B 0.02096f
C458 VTAIL.n54 B 0.02096f
C459 VTAIL.n55 B 0.009129f
C460 VTAIL.n56 B 0.008868f
C461 VTAIL.n57 B 0.016503f
C462 VTAIL.n58 B 0.016503f
C463 VTAIL.n59 B 0.008868f
C464 VTAIL.n60 B 0.009389f
C465 VTAIL.n61 B 0.02096f
C466 VTAIL.n62 B 0.02096f
C467 VTAIL.n63 B 0.009389f
C468 VTAIL.n64 B 0.008868f
C469 VTAIL.n65 B 0.016503f
C470 VTAIL.n66 B 0.016503f
C471 VTAIL.n67 B 0.008868f
C472 VTAIL.n68 B 0.009389f
C473 VTAIL.n69 B 0.02096f
C474 VTAIL.n70 B 0.02096f
C475 VTAIL.n71 B 0.009389f
C476 VTAIL.n72 B 0.008868f
C477 VTAIL.n73 B 0.016503f
C478 VTAIL.n74 B 0.016503f
C479 VTAIL.n75 B 0.008868f
C480 VTAIL.n76 B 0.009389f
C481 VTAIL.n77 B 0.02096f
C482 VTAIL.n78 B 0.02096f
C483 VTAIL.n79 B 0.009389f
C484 VTAIL.n80 B 0.008868f
C485 VTAIL.n81 B 0.016503f
C486 VTAIL.n82 B 0.016503f
C487 VTAIL.n83 B 0.008868f
C488 VTAIL.n84 B 0.009389f
C489 VTAIL.n85 B 0.02096f
C490 VTAIL.n86 B 0.02096f
C491 VTAIL.n87 B 0.009389f
C492 VTAIL.n88 B 0.008868f
C493 VTAIL.n89 B 0.016503f
C494 VTAIL.n90 B 0.042654f
C495 VTAIL.n91 B 0.008868f
C496 VTAIL.n92 B 0.009389f
C497 VTAIL.n93 B 0.041437f
C498 VTAIL.n94 B 0.035334f
C499 VTAIL.n95 B 1.16334f
C500 VTAIL.n96 B 0.009304f
C501 VTAIL.n97 B 0.02096f
C502 VTAIL.n98 B 0.009389f
C503 VTAIL.n99 B 0.016503f
C504 VTAIL.n100 B 0.008868f
C505 VTAIL.n101 B 0.02096f
C506 VTAIL.n102 B 0.009389f
C507 VTAIL.n103 B 0.016503f
C508 VTAIL.n104 B 0.008868f
C509 VTAIL.n105 B 0.02096f
C510 VTAIL.n106 B 0.009389f
C511 VTAIL.n107 B 0.016503f
C512 VTAIL.n108 B 0.008868f
C513 VTAIL.n109 B 0.02096f
C514 VTAIL.n110 B 0.009389f
C515 VTAIL.n111 B 0.016503f
C516 VTAIL.n112 B 0.008868f
C517 VTAIL.n113 B 0.02096f
C518 VTAIL.n114 B 0.009389f
C519 VTAIL.n115 B 0.016503f
C520 VTAIL.n116 B 0.009129f
C521 VTAIL.n117 B 0.02096f
C522 VTAIL.n118 B 0.008868f
C523 VTAIL.n119 B 0.009389f
C524 VTAIL.n120 B 0.016503f
C525 VTAIL.n121 B 0.008868f
C526 VTAIL.n122 B 0.02096f
C527 VTAIL.n123 B 0.009389f
C528 VTAIL.n124 B 0.016503f
C529 VTAIL.n125 B 0.008868f
C530 VTAIL.n126 B 0.01572f
C531 VTAIL.n127 B 0.014817f
C532 VTAIL.t2 B 0.035877f
C533 VTAIL.n128 B 0.152941f
C534 VTAIL.n129 B 1.22596f
C535 VTAIL.n130 B 0.008868f
C536 VTAIL.n131 B 0.009389f
C537 VTAIL.n132 B 0.02096f
C538 VTAIL.n133 B 0.02096f
C539 VTAIL.n134 B 0.009389f
C540 VTAIL.n135 B 0.008868f
C541 VTAIL.n136 B 0.016503f
C542 VTAIL.n137 B 0.016503f
C543 VTAIL.n138 B 0.008868f
C544 VTAIL.n139 B 0.009389f
C545 VTAIL.n140 B 0.02096f
C546 VTAIL.n141 B 0.02096f
C547 VTAIL.n142 B 0.009389f
C548 VTAIL.n143 B 0.008868f
C549 VTAIL.n144 B 0.016503f
C550 VTAIL.n145 B 0.016503f
C551 VTAIL.n146 B 0.008868f
C552 VTAIL.n147 B 0.009389f
C553 VTAIL.n148 B 0.02096f
C554 VTAIL.n149 B 0.02096f
C555 VTAIL.n150 B 0.02096f
C556 VTAIL.n151 B 0.009129f
C557 VTAIL.n152 B 0.008868f
C558 VTAIL.n153 B 0.016503f
C559 VTAIL.n154 B 0.016503f
C560 VTAIL.n155 B 0.008868f
C561 VTAIL.n156 B 0.009389f
C562 VTAIL.n157 B 0.02096f
C563 VTAIL.n158 B 0.02096f
C564 VTAIL.n159 B 0.009389f
C565 VTAIL.n160 B 0.008868f
C566 VTAIL.n161 B 0.016503f
C567 VTAIL.n162 B 0.016503f
C568 VTAIL.n163 B 0.008868f
C569 VTAIL.n164 B 0.009389f
C570 VTAIL.n165 B 0.02096f
C571 VTAIL.n166 B 0.02096f
C572 VTAIL.n167 B 0.009389f
C573 VTAIL.n168 B 0.008868f
C574 VTAIL.n169 B 0.016503f
C575 VTAIL.n170 B 0.016503f
C576 VTAIL.n171 B 0.008868f
C577 VTAIL.n172 B 0.009389f
C578 VTAIL.n173 B 0.02096f
C579 VTAIL.n174 B 0.02096f
C580 VTAIL.n175 B 0.009389f
C581 VTAIL.n176 B 0.008868f
C582 VTAIL.n177 B 0.016503f
C583 VTAIL.n178 B 0.016503f
C584 VTAIL.n179 B 0.008868f
C585 VTAIL.n180 B 0.009389f
C586 VTAIL.n181 B 0.02096f
C587 VTAIL.n182 B 0.02096f
C588 VTAIL.n183 B 0.009389f
C589 VTAIL.n184 B 0.008868f
C590 VTAIL.n185 B 0.016503f
C591 VTAIL.n186 B 0.042654f
C592 VTAIL.n187 B 0.008868f
C593 VTAIL.n188 B 0.009389f
C594 VTAIL.n189 B 0.041437f
C595 VTAIL.n190 B 0.035334f
C596 VTAIL.n191 B 1.17125f
C597 VTAIL.n192 B 0.009304f
C598 VTAIL.n193 B 0.02096f
C599 VTAIL.n194 B 0.009389f
C600 VTAIL.n195 B 0.016503f
C601 VTAIL.n196 B 0.008868f
C602 VTAIL.n197 B 0.02096f
C603 VTAIL.n198 B 0.009389f
C604 VTAIL.n199 B 0.016503f
C605 VTAIL.n200 B 0.008868f
C606 VTAIL.n201 B 0.02096f
C607 VTAIL.n202 B 0.009389f
C608 VTAIL.n203 B 0.016503f
C609 VTAIL.n204 B 0.008868f
C610 VTAIL.n205 B 0.02096f
C611 VTAIL.n206 B 0.009389f
C612 VTAIL.n207 B 0.016503f
C613 VTAIL.n208 B 0.008868f
C614 VTAIL.n209 B 0.02096f
C615 VTAIL.n210 B 0.009389f
C616 VTAIL.n211 B 0.016503f
C617 VTAIL.n212 B 0.009129f
C618 VTAIL.n213 B 0.02096f
C619 VTAIL.n214 B 0.008868f
C620 VTAIL.n215 B 0.009389f
C621 VTAIL.n216 B 0.016503f
C622 VTAIL.n217 B 0.008868f
C623 VTAIL.n218 B 0.02096f
C624 VTAIL.n219 B 0.009389f
C625 VTAIL.n220 B 0.016503f
C626 VTAIL.n221 B 0.008868f
C627 VTAIL.n222 B 0.01572f
C628 VTAIL.n223 B 0.014817f
C629 VTAIL.t0 B 0.035877f
C630 VTAIL.n224 B 0.152941f
C631 VTAIL.n225 B 1.22596f
C632 VTAIL.n226 B 0.008868f
C633 VTAIL.n227 B 0.009389f
C634 VTAIL.n228 B 0.02096f
C635 VTAIL.n229 B 0.02096f
C636 VTAIL.n230 B 0.009389f
C637 VTAIL.n231 B 0.008868f
C638 VTAIL.n232 B 0.016503f
C639 VTAIL.n233 B 0.016503f
C640 VTAIL.n234 B 0.008868f
C641 VTAIL.n235 B 0.009389f
C642 VTAIL.n236 B 0.02096f
C643 VTAIL.n237 B 0.02096f
C644 VTAIL.n238 B 0.009389f
C645 VTAIL.n239 B 0.008868f
C646 VTAIL.n240 B 0.016503f
C647 VTAIL.n241 B 0.016503f
C648 VTAIL.n242 B 0.008868f
C649 VTAIL.n243 B 0.009389f
C650 VTAIL.n244 B 0.02096f
C651 VTAIL.n245 B 0.02096f
C652 VTAIL.n246 B 0.02096f
C653 VTAIL.n247 B 0.009129f
C654 VTAIL.n248 B 0.008868f
C655 VTAIL.n249 B 0.016503f
C656 VTAIL.n250 B 0.016503f
C657 VTAIL.n251 B 0.008868f
C658 VTAIL.n252 B 0.009389f
C659 VTAIL.n253 B 0.02096f
C660 VTAIL.n254 B 0.02096f
C661 VTAIL.n255 B 0.009389f
C662 VTAIL.n256 B 0.008868f
C663 VTAIL.n257 B 0.016503f
C664 VTAIL.n258 B 0.016503f
C665 VTAIL.n259 B 0.008868f
C666 VTAIL.n260 B 0.009389f
C667 VTAIL.n261 B 0.02096f
C668 VTAIL.n262 B 0.02096f
C669 VTAIL.n263 B 0.009389f
C670 VTAIL.n264 B 0.008868f
C671 VTAIL.n265 B 0.016503f
C672 VTAIL.n266 B 0.016503f
C673 VTAIL.n267 B 0.008868f
C674 VTAIL.n268 B 0.009389f
C675 VTAIL.n269 B 0.02096f
C676 VTAIL.n270 B 0.02096f
C677 VTAIL.n271 B 0.009389f
C678 VTAIL.n272 B 0.008868f
C679 VTAIL.n273 B 0.016503f
C680 VTAIL.n274 B 0.016503f
C681 VTAIL.n275 B 0.008868f
C682 VTAIL.n276 B 0.009389f
C683 VTAIL.n277 B 0.02096f
C684 VTAIL.n278 B 0.02096f
C685 VTAIL.n279 B 0.009389f
C686 VTAIL.n280 B 0.008868f
C687 VTAIL.n281 B 0.016503f
C688 VTAIL.n282 B 0.042654f
C689 VTAIL.n283 B 0.008868f
C690 VTAIL.n284 B 0.009389f
C691 VTAIL.n285 B 0.041437f
C692 VTAIL.n286 B 0.035334f
C693 VTAIL.n287 B 1.12724f
C694 VTAIL.n288 B 0.009304f
C695 VTAIL.n289 B 0.02096f
C696 VTAIL.n290 B 0.009389f
C697 VTAIL.n291 B 0.016503f
C698 VTAIL.n292 B 0.008868f
C699 VTAIL.n293 B 0.02096f
C700 VTAIL.n294 B 0.009389f
C701 VTAIL.n295 B 0.016503f
C702 VTAIL.n296 B 0.008868f
C703 VTAIL.n297 B 0.02096f
C704 VTAIL.n298 B 0.009389f
C705 VTAIL.n299 B 0.016503f
C706 VTAIL.n300 B 0.008868f
C707 VTAIL.n301 B 0.02096f
C708 VTAIL.n302 B 0.009389f
C709 VTAIL.n303 B 0.016503f
C710 VTAIL.n304 B 0.008868f
C711 VTAIL.n305 B 0.02096f
C712 VTAIL.n306 B 0.009389f
C713 VTAIL.n307 B 0.016503f
C714 VTAIL.n308 B 0.009129f
C715 VTAIL.n309 B 0.02096f
C716 VTAIL.n310 B 0.009389f
C717 VTAIL.n311 B 0.016503f
C718 VTAIL.n312 B 0.008868f
C719 VTAIL.n313 B 0.02096f
C720 VTAIL.n314 B 0.009389f
C721 VTAIL.n315 B 0.016503f
C722 VTAIL.n316 B 0.008868f
C723 VTAIL.n317 B 0.01572f
C724 VTAIL.n318 B 0.014817f
C725 VTAIL.t3 B 0.035877f
C726 VTAIL.n319 B 0.152941f
C727 VTAIL.n320 B 1.22596f
C728 VTAIL.n321 B 0.008868f
C729 VTAIL.n322 B 0.009389f
C730 VTAIL.n323 B 0.02096f
C731 VTAIL.n324 B 0.02096f
C732 VTAIL.n325 B 0.009389f
C733 VTAIL.n326 B 0.008868f
C734 VTAIL.n327 B 0.016503f
C735 VTAIL.n328 B 0.016503f
C736 VTAIL.n329 B 0.008868f
C737 VTAIL.n330 B 0.009389f
C738 VTAIL.n331 B 0.02096f
C739 VTAIL.n332 B 0.02096f
C740 VTAIL.n333 B 0.009389f
C741 VTAIL.n334 B 0.008868f
C742 VTAIL.n335 B 0.016503f
C743 VTAIL.n336 B 0.016503f
C744 VTAIL.n337 B 0.008868f
C745 VTAIL.n338 B 0.008868f
C746 VTAIL.n339 B 0.009389f
C747 VTAIL.n340 B 0.02096f
C748 VTAIL.n341 B 0.02096f
C749 VTAIL.n342 B 0.02096f
C750 VTAIL.n343 B 0.009129f
C751 VTAIL.n344 B 0.008868f
C752 VTAIL.n345 B 0.016503f
C753 VTAIL.n346 B 0.016503f
C754 VTAIL.n347 B 0.008868f
C755 VTAIL.n348 B 0.009389f
C756 VTAIL.n349 B 0.02096f
C757 VTAIL.n350 B 0.02096f
C758 VTAIL.n351 B 0.009389f
C759 VTAIL.n352 B 0.008868f
C760 VTAIL.n353 B 0.016503f
C761 VTAIL.n354 B 0.016503f
C762 VTAIL.n355 B 0.008868f
C763 VTAIL.n356 B 0.009389f
C764 VTAIL.n357 B 0.02096f
C765 VTAIL.n358 B 0.02096f
C766 VTAIL.n359 B 0.009389f
C767 VTAIL.n360 B 0.008868f
C768 VTAIL.n361 B 0.016503f
C769 VTAIL.n362 B 0.016503f
C770 VTAIL.n363 B 0.008868f
C771 VTAIL.n364 B 0.009389f
C772 VTAIL.n365 B 0.02096f
C773 VTAIL.n366 B 0.02096f
C774 VTAIL.n367 B 0.009389f
C775 VTAIL.n368 B 0.008868f
C776 VTAIL.n369 B 0.016503f
C777 VTAIL.n370 B 0.016503f
C778 VTAIL.n371 B 0.008868f
C779 VTAIL.n372 B 0.009389f
C780 VTAIL.n373 B 0.02096f
C781 VTAIL.n374 B 0.02096f
C782 VTAIL.n375 B 0.009389f
C783 VTAIL.n376 B 0.008868f
C784 VTAIL.n377 B 0.016503f
C785 VTAIL.n378 B 0.042654f
C786 VTAIL.n379 B 0.008868f
C787 VTAIL.n380 B 0.009389f
C788 VTAIL.n381 B 0.041437f
C789 VTAIL.n382 B 0.035334f
C790 VTAIL.n383 B 1.08816f
C791 VN.t1 B 1.55132f
C792 VN.t0 B 1.67033f
.ends

