* NGSPICE file created from diff_pair_sample_1096.ext - technology: sky130A

.subckt diff_pair_sample_1096 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0.44055 ps=3 w=2.67 l=2.62
X1 B.t11 B.t9 B.t10 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0 ps=0 w=2.67 l=2.62
X2 VDD1.t7 VP.t1 VTAIL.t14 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=1.0413 ps=6.12 w=2.67 l=2.62
X3 VDD2.t7 VN.t0 VTAIL.t3 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X4 VDD2.t6 VN.t1 VTAIL.t5 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=1.0413 ps=6.12 w=2.67 l=2.62
X5 VTAIL.t4 VN.t2 VDD2.t5 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0.44055 ps=3 w=2.67 l=2.62
X6 VDD1.t4 VP.t2 VTAIL.t13 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X7 VDD2.t4 VN.t3 VTAIL.t7 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=1.0413 ps=6.12 w=2.67 l=2.62
X8 VTAIL.t12 VP.t3 VDD1.t0 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0.44055 ps=3 w=2.67 l=2.62
X9 VDD2.t3 VN.t4 VTAIL.t2 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X10 VDD1.t1 VP.t4 VTAIL.t11 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X11 B.t8 B.t6 B.t7 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0 ps=0 w=2.67 l=2.62
X12 B.t5 B.t3 B.t4 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0 ps=0 w=2.67 l=2.62
X13 VTAIL.t10 VP.t5 VDD1.t2 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X14 B.t2 B.t0 B.t1 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0 ps=0 w=2.67 l=2.62
X15 VTAIL.t9 VP.t6 VDD1.t5 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X16 VTAIL.t1 VN.t5 VDD2.t2 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
X17 VTAIL.t0 VN.t6 VDD2.t1 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=1.0413 pd=6.12 as=0.44055 ps=3 w=2.67 l=2.62
X18 VDD1.t6 VP.t7 VTAIL.t8 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=1.0413 ps=6.12 w=2.67 l=2.62
X19 VTAIL.t6 VN.t7 VDD2.t0 w_n3920_n1502# sky130_fd_pr__pfet_01v8 ad=0.44055 pd=3 as=0.44055 ps=3 w=2.67 l=2.62
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n12 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n33 VP.n11 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n36 VP.n10 161.3
R12 VP.n68 VP.n0 161.3
R13 VP.n67 VP.n66 161.3
R14 VP.n65 VP.n1 161.3
R15 VP.n64 VP.n63 161.3
R16 VP.n62 VP.n2 161.3
R17 VP.n61 VP.n60 161.3
R18 VP.n59 VP.n58 161.3
R19 VP.n57 VP.n4 161.3
R20 VP.n56 VP.n55 161.3
R21 VP.n54 VP.n5 161.3
R22 VP.n53 VP.n52 161.3
R23 VP.n51 VP.n6 161.3
R24 VP.n49 VP.n48 161.3
R25 VP.n47 VP.n7 161.3
R26 VP.n46 VP.n45 161.3
R27 VP.n44 VP.n8 161.3
R28 VP.n43 VP.n42 161.3
R29 VP.n41 VP.n9 161.3
R30 VP.n40 VP.n39 102.192
R31 VP.n70 VP.n69 102.192
R32 VP.n38 VP.n37 102.192
R33 VP.n18 VP.n17 61.3525
R34 VP.n17 VP.t0 57.7507
R35 VP.n45 VP.n44 56.5193
R36 VP.n56 VP.n5 56.5193
R37 VP.n63 VP.n1 56.5193
R38 VP.n31 VP.n11 56.5193
R39 VP.n24 VP.n15 56.5193
R40 VP.n40 VP.n38 43.9238
R41 VP.n39 VP.t3 24.5604
R42 VP.n50 VP.t4 24.5604
R43 VP.n3 VP.t5 24.5604
R44 VP.n69 VP.t7 24.5604
R45 VP.n37 VP.t1 24.5604
R46 VP.n13 VP.t6 24.5604
R47 VP.n18 VP.t2 24.5604
R48 VP.n43 VP.n9 24.4675
R49 VP.n44 VP.n43 24.4675
R50 VP.n45 VP.n7 24.4675
R51 VP.n49 VP.n7 24.4675
R52 VP.n52 VP.n51 24.4675
R53 VP.n52 VP.n5 24.4675
R54 VP.n57 VP.n56 24.4675
R55 VP.n58 VP.n57 24.4675
R56 VP.n62 VP.n61 24.4675
R57 VP.n63 VP.n62 24.4675
R58 VP.n67 VP.n1 24.4675
R59 VP.n68 VP.n67 24.4675
R60 VP.n35 VP.n11 24.4675
R61 VP.n36 VP.n35 24.4675
R62 VP.n25 VP.n24 24.4675
R63 VP.n26 VP.n25 24.4675
R64 VP.n30 VP.n29 24.4675
R65 VP.n31 VP.n30 24.4675
R66 VP.n20 VP.n19 24.4675
R67 VP.n20 VP.n15 24.4675
R68 VP.n50 VP.n49 13.4574
R69 VP.n61 VP.n3 13.4574
R70 VP.n29 VP.n13 13.4574
R71 VP.n51 VP.n50 11.0107
R72 VP.n58 VP.n3 11.0107
R73 VP.n26 VP.n13 11.0107
R74 VP.n19 VP.n18 11.0107
R75 VP.n39 VP.n9 8.56395
R76 VP.n69 VP.n68 8.56395
R77 VP.n37 VP.n36 8.56395
R78 VP.n17 VP.n16 6.94033
R79 VP.n38 VP.n10 0.278367
R80 VP.n41 VP.n40 0.278367
R81 VP.n70 VP.n0 0.278367
R82 VP.n21 VP.n16 0.189894
R83 VP.n22 VP.n21 0.189894
R84 VP.n23 VP.n22 0.189894
R85 VP.n23 VP.n14 0.189894
R86 VP.n27 VP.n14 0.189894
R87 VP.n28 VP.n27 0.189894
R88 VP.n28 VP.n12 0.189894
R89 VP.n32 VP.n12 0.189894
R90 VP.n33 VP.n32 0.189894
R91 VP.n34 VP.n33 0.189894
R92 VP.n34 VP.n10 0.189894
R93 VP.n42 VP.n41 0.189894
R94 VP.n42 VP.n8 0.189894
R95 VP.n46 VP.n8 0.189894
R96 VP.n47 VP.n46 0.189894
R97 VP.n48 VP.n47 0.189894
R98 VP.n48 VP.n6 0.189894
R99 VP.n53 VP.n6 0.189894
R100 VP.n54 VP.n53 0.189894
R101 VP.n55 VP.n54 0.189894
R102 VP.n55 VP.n4 0.189894
R103 VP.n59 VP.n4 0.189894
R104 VP.n60 VP.n59 0.189894
R105 VP.n60 VP.n2 0.189894
R106 VP.n64 VP.n2 0.189894
R107 VP.n65 VP.n64 0.189894
R108 VP.n66 VP.n65 0.189894
R109 VP.n66 VP.n0 0.189894
R110 VP VP.n70 0.153454
R111 VDD1 VDD1.n0 152.714
R112 VDD1.n3 VDD1.n2 152.6
R113 VDD1.n3 VDD1.n1 152.6
R114 VDD1.n5 VDD1.n4 151.383
R115 VDD1.n5 VDD1.n3 38.044
R116 VDD1.n4 VDD1.t5 12.1747
R117 VDD1.n4 VDD1.t7 12.1747
R118 VDD1.n0 VDD1.t3 12.1747
R119 VDD1.n0 VDD1.t4 12.1747
R120 VDD1.n2 VDD1.t2 12.1747
R121 VDD1.n2 VDD1.t6 12.1747
R122 VDD1.n1 VDD1.t0 12.1747
R123 VDD1.n1 VDD1.t1 12.1747
R124 VDD1 VDD1.n5 1.21386
R125 VTAIL.n98 VTAIL.n92 756.745
R126 VTAIL.n8 VTAIL.n2 756.745
R127 VTAIL.n20 VTAIL.n14 756.745
R128 VTAIL.n34 VTAIL.n28 756.745
R129 VTAIL.n86 VTAIL.n80 756.745
R130 VTAIL.n72 VTAIL.n66 756.745
R131 VTAIL.n60 VTAIL.n54 756.745
R132 VTAIL.n46 VTAIL.n40 756.745
R133 VTAIL.n97 VTAIL.n96 585
R134 VTAIL.n99 VTAIL.n98 585
R135 VTAIL.n7 VTAIL.n6 585
R136 VTAIL.n9 VTAIL.n8 585
R137 VTAIL.n19 VTAIL.n18 585
R138 VTAIL.n21 VTAIL.n20 585
R139 VTAIL.n33 VTAIL.n32 585
R140 VTAIL.n35 VTAIL.n34 585
R141 VTAIL.n87 VTAIL.n86 585
R142 VTAIL.n85 VTAIL.n84 585
R143 VTAIL.n73 VTAIL.n72 585
R144 VTAIL.n71 VTAIL.n70 585
R145 VTAIL.n61 VTAIL.n60 585
R146 VTAIL.n59 VTAIL.n58 585
R147 VTAIL.n47 VTAIL.n46 585
R148 VTAIL.n45 VTAIL.n44 585
R149 VTAIL.n95 VTAIL.t5 357.269
R150 VTAIL.n5 VTAIL.t4 357.269
R151 VTAIL.n17 VTAIL.t8 357.269
R152 VTAIL.n31 VTAIL.t12 357.269
R153 VTAIL.n83 VTAIL.t14 357.269
R154 VTAIL.n69 VTAIL.t15 357.269
R155 VTAIL.n57 VTAIL.t7 357.269
R156 VTAIL.n43 VTAIL.t0 357.269
R157 VTAIL.n98 VTAIL.n97 171.744
R158 VTAIL.n8 VTAIL.n7 171.744
R159 VTAIL.n20 VTAIL.n19 171.744
R160 VTAIL.n34 VTAIL.n33 171.744
R161 VTAIL.n86 VTAIL.n85 171.744
R162 VTAIL.n72 VTAIL.n71 171.744
R163 VTAIL.n60 VTAIL.n59 171.744
R164 VTAIL.n46 VTAIL.n45 171.744
R165 VTAIL.n1 VTAIL.n0 134.704
R166 VTAIL.n27 VTAIL.n26 134.704
R167 VTAIL.n79 VTAIL.n78 134.704
R168 VTAIL.n53 VTAIL.n52 134.704
R169 VTAIL.n97 VTAIL.t5 85.8723
R170 VTAIL.n7 VTAIL.t4 85.8723
R171 VTAIL.n19 VTAIL.t8 85.8723
R172 VTAIL.n33 VTAIL.t12 85.8723
R173 VTAIL.n85 VTAIL.t14 85.8723
R174 VTAIL.n71 VTAIL.t15 85.8723
R175 VTAIL.n59 VTAIL.t7 85.8723
R176 VTAIL.n45 VTAIL.t0 85.8723
R177 VTAIL.n103 VTAIL.n102 30.4399
R178 VTAIL.n13 VTAIL.n12 30.4399
R179 VTAIL.n25 VTAIL.n24 30.4399
R180 VTAIL.n39 VTAIL.n38 30.4399
R181 VTAIL.n91 VTAIL.n90 30.4399
R182 VTAIL.n77 VTAIL.n76 30.4399
R183 VTAIL.n65 VTAIL.n64 30.4399
R184 VTAIL.n51 VTAIL.n50 30.4399
R185 VTAIL.n103 VTAIL.n91 17.2117
R186 VTAIL.n51 VTAIL.n39 17.2117
R187 VTAIL.n0 VTAIL.t3 12.1747
R188 VTAIL.n0 VTAIL.t6 12.1747
R189 VTAIL.n26 VTAIL.t11 12.1747
R190 VTAIL.n26 VTAIL.t10 12.1747
R191 VTAIL.n78 VTAIL.t13 12.1747
R192 VTAIL.n78 VTAIL.t9 12.1747
R193 VTAIL.n52 VTAIL.t2 12.1747
R194 VTAIL.n52 VTAIL.t1 12.1747
R195 VTAIL.n96 VTAIL.n95 10.3978
R196 VTAIL.n6 VTAIL.n5 10.3978
R197 VTAIL.n18 VTAIL.n17 10.3978
R198 VTAIL.n32 VTAIL.n31 10.3978
R199 VTAIL.n84 VTAIL.n83 10.3978
R200 VTAIL.n70 VTAIL.n69 10.3978
R201 VTAIL.n58 VTAIL.n57 10.3978
R202 VTAIL.n44 VTAIL.n43 10.3978
R203 VTAIL.n102 VTAIL.n101 9.45567
R204 VTAIL.n12 VTAIL.n11 9.45567
R205 VTAIL.n24 VTAIL.n23 9.45567
R206 VTAIL.n38 VTAIL.n37 9.45567
R207 VTAIL.n90 VTAIL.n89 9.45567
R208 VTAIL.n76 VTAIL.n75 9.45567
R209 VTAIL.n64 VTAIL.n63 9.45567
R210 VTAIL.n50 VTAIL.n49 9.45567
R211 VTAIL.n94 VTAIL.n93 9.3005
R212 VTAIL.n101 VTAIL.n100 9.3005
R213 VTAIL.n4 VTAIL.n3 9.3005
R214 VTAIL.n11 VTAIL.n10 9.3005
R215 VTAIL.n16 VTAIL.n15 9.3005
R216 VTAIL.n23 VTAIL.n22 9.3005
R217 VTAIL.n30 VTAIL.n29 9.3005
R218 VTAIL.n37 VTAIL.n36 9.3005
R219 VTAIL.n82 VTAIL.n81 9.3005
R220 VTAIL.n89 VTAIL.n88 9.3005
R221 VTAIL.n75 VTAIL.n74 9.3005
R222 VTAIL.n68 VTAIL.n67 9.3005
R223 VTAIL.n63 VTAIL.n62 9.3005
R224 VTAIL.n56 VTAIL.n55 9.3005
R225 VTAIL.n49 VTAIL.n48 9.3005
R226 VTAIL.n42 VTAIL.n41 9.3005
R227 VTAIL.n102 VTAIL.n92 8.92171
R228 VTAIL.n12 VTAIL.n2 8.92171
R229 VTAIL.n24 VTAIL.n14 8.92171
R230 VTAIL.n38 VTAIL.n28 8.92171
R231 VTAIL.n90 VTAIL.n80 8.92171
R232 VTAIL.n76 VTAIL.n66 8.92171
R233 VTAIL.n64 VTAIL.n54 8.92171
R234 VTAIL.n50 VTAIL.n40 8.92171
R235 VTAIL.n100 VTAIL.n99 8.14595
R236 VTAIL.n10 VTAIL.n9 8.14595
R237 VTAIL.n22 VTAIL.n21 8.14595
R238 VTAIL.n36 VTAIL.n35 8.14595
R239 VTAIL.n88 VTAIL.n87 8.14595
R240 VTAIL.n74 VTAIL.n73 8.14595
R241 VTAIL.n62 VTAIL.n61 8.14595
R242 VTAIL.n48 VTAIL.n47 8.14595
R243 VTAIL.n96 VTAIL.n94 7.3702
R244 VTAIL.n6 VTAIL.n4 7.3702
R245 VTAIL.n18 VTAIL.n16 7.3702
R246 VTAIL.n32 VTAIL.n30 7.3702
R247 VTAIL.n84 VTAIL.n82 7.3702
R248 VTAIL.n70 VTAIL.n68 7.3702
R249 VTAIL.n58 VTAIL.n56 7.3702
R250 VTAIL.n44 VTAIL.n42 7.3702
R251 VTAIL.n99 VTAIL.n94 5.81868
R252 VTAIL.n9 VTAIL.n4 5.81868
R253 VTAIL.n21 VTAIL.n16 5.81868
R254 VTAIL.n35 VTAIL.n30 5.81868
R255 VTAIL.n87 VTAIL.n82 5.81868
R256 VTAIL.n73 VTAIL.n68 5.81868
R257 VTAIL.n61 VTAIL.n56 5.81868
R258 VTAIL.n47 VTAIL.n42 5.81868
R259 VTAIL.n100 VTAIL.n92 5.04292
R260 VTAIL.n10 VTAIL.n2 5.04292
R261 VTAIL.n22 VTAIL.n14 5.04292
R262 VTAIL.n36 VTAIL.n28 5.04292
R263 VTAIL.n88 VTAIL.n80 5.04292
R264 VTAIL.n74 VTAIL.n66 5.04292
R265 VTAIL.n62 VTAIL.n54 5.04292
R266 VTAIL.n48 VTAIL.n40 5.04292
R267 VTAIL.n95 VTAIL.n93 2.74506
R268 VTAIL.n5 VTAIL.n3 2.74506
R269 VTAIL.n17 VTAIL.n15 2.74506
R270 VTAIL.n31 VTAIL.n29 2.74506
R271 VTAIL.n83 VTAIL.n81 2.74506
R272 VTAIL.n69 VTAIL.n67 2.74506
R273 VTAIL.n57 VTAIL.n55 2.74506
R274 VTAIL.n43 VTAIL.n41 2.74506
R275 VTAIL.n53 VTAIL.n51 2.5436
R276 VTAIL.n65 VTAIL.n53 2.5436
R277 VTAIL.n79 VTAIL.n77 2.5436
R278 VTAIL.n91 VTAIL.n79 2.5436
R279 VTAIL.n39 VTAIL.n27 2.5436
R280 VTAIL.n27 VTAIL.n25 2.5436
R281 VTAIL.n13 VTAIL.n1 2.5436
R282 VTAIL VTAIL.n103 2.48541
R283 VTAIL.n77 VTAIL.n65 0.470328
R284 VTAIL.n25 VTAIL.n13 0.470328
R285 VTAIL.n101 VTAIL.n93 0.155672
R286 VTAIL.n11 VTAIL.n3 0.155672
R287 VTAIL.n23 VTAIL.n15 0.155672
R288 VTAIL.n37 VTAIL.n29 0.155672
R289 VTAIL.n89 VTAIL.n81 0.155672
R290 VTAIL.n75 VTAIL.n67 0.155672
R291 VTAIL.n63 VTAIL.n55 0.155672
R292 VTAIL.n49 VTAIL.n41 0.155672
R293 VTAIL VTAIL.n1 0.0586897
R294 B.n285 B.n284 585
R295 B.n283 B.n104 585
R296 B.n282 B.n281 585
R297 B.n280 B.n105 585
R298 B.n279 B.n278 585
R299 B.n277 B.n106 585
R300 B.n276 B.n275 585
R301 B.n274 B.n107 585
R302 B.n273 B.n272 585
R303 B.n271 B.n108 585
R304 B.n270 B.n269 585
R305 B.n268 B.n109 585
R306 B.n267 B.n266 585
R307 B.n265 B.n110 585
R308 B.n263 B.n262 585
R309 B.n261 B.n113 585
R310 B.n260 B.n259 585
R311 B.n258 B.n114 585
R312 B.n257 B.n256 585
R313 B.n255 B.n115 585
R314 B.n254 B.n253 585
R315 B.n252 B.n116 585
R316 B.n251 B.n250 585
R317 B.n249 B.n117 585
R318 B.n248 B.n247 585
R319 B.n243 B.n118 585
R320 B.n242 B.n241 585
R321 B.n240 B.n119 585
R322 B.n239 B.n238 585
R323 B.n237 B.n120 585
R324 B.n236 B.n235 585
R325 B.n234 B.n121 585
R326 B.n233 B.n232 585
R327 B.n231 B.n122 585
R328 B.n230 B.n229 585
R329 B.n228 B.n123 585
R330 B.n227 B.n226 585
R331 B.n225 B.n124 585
R332 B.n286 B.n103 585
R333 B.n288 B.n287 585
R334 B.n289 B.n102 585
R335 B.n291 B.n290 585
R336 B.n292 B.n101 585
R337 B.n294 B.n293 585
R338 B.n295 B.n100 585
R339 B.n297 B.n296 585
R340 B.n298 B.n99 585
R341 B.n300 B.n299 585
R342 B.n301 B.n98 585
R343 B.n303 B.n302 585
R344 B.n304 B.n97 585
R345 B.n306 B.n305 585
R346 B.n307 B.n96 585
R347 B.n309 B.n308 585
R348 B.n310 B.n95 585
R349 B.n312 B.n311 585
R350 B.n313 B.n94 585
R351 B.n315 B.n314 585
R352 B.n316 B.n93 585
R353 B.n318 B.n317 585
R354 B.n319 B.n92 585
R355 B.n321 B.n320 585
R356 B.n322 B.n91 585
R357 B.n324 B.n323 585
R358 B.n325 B.n90 585
R359 B.n327 B.n326 585
R360 B.n328 B.n89 585
R361 B.n330 B.n329 585
R362 B.n331 B.n88 585
R363 B.n333 B.n332 585
R364 B.n334 B.n87 585
R365 B.n336 B.n335 585
R366 B.n337 B.n86 585
R367 B.n339 B.n338 585
R368 B.n340 B.n85 585
R369 B.n342 B.n341 585
R370 B.n343 B.n84 585
R371 B.n345 B.n344 585
R372 B.n346 B.n83 585
R373 B.n348 B.n347 585
R374 B.n349 B.n82 585
R375 B.n351 B.n350 585
R376 B.n352 B.n81 585
R377 B.n354 B.n353 585
R378 B.n355 B.n80 585
R379 B.n357 B.n356 585
R380 B.n358 B.n79 585
R381 B.n360 B.n359 585
R382 B.n361 B.n78 585
R383 B.n363 B.n362 585
R384 B.n364 B.n77 585
R385 B.n366 B.n365 585
R386 B.n367 B.n76 585
R387 B.n369 B.n368 585
R388 B.n370 B.n75 585
R389 B.n372 B.n371 585
R390 B.n373 B.n74 585
R391 B.n375 B.n374 585
R392 B.n376 B.n73 585
R393 B.n378 B.n377 585
R394 B.n379 B.n72 585
R395 B.n381 B.n380 585
R396 B.n382 B.n71 585
R397 B.n384 B.n383 585
R398 B.n385 B.n70 585
R399 B.n387 B.n386 585
R400 B.n388 B.n69 585
R401 B.n390 B.n389 585
R402 B.n391 B.n68 585
R403 B.n393 B.n392 585
R404 B.n394 B.n67 585
R405 B.n396 B.n395 585
R406 B.n397 B.n66 585
R407 B.n399 B.n398 585
R408 B.n400 B.n65 585
R409 B.n402 B.n401 585
R410 B.n403 B.n64 585
R411 B.n405 B.n404 585
R412 B.n406 B.n63 585
R413 B.n408 B.n407 585
R414 B.n409 B.n62 585
R415 B.n411 B.n410 585
R416 B.n412 B.n61 585
R417 B.n414 B.n413 585
R418 B.n415 B.n60 585
R419 B.n417 B.n416 585
R420 B.n418 B.n59 585
R421 B.n420 B.n419 585
R422 B.n421 B.n58 585
R423 B.n423 B.n422 585
R424 B.n424 B.n57 585
R425 B.n426 B.n425 585
R426 B.n427 B.n56 585
R427 B.n429 B.n428 585
R428 B.n430 B.n55 585
R429 B.n432 B.n431 585
R430 B.n433 B.n54 585
R431 B.n435 B.n434 585
R432 B.n436 B.n53 585
R433 B.n438 B.n437 585
R434 B.n439 B.n52 585
R435 B.n441 B.n440 585
R436 B.n499 B.n498 585
R437 B.n497 B.n28 585
R438 B.n496 B.n495 585
R439 B.n494 B.n29 585
R440 B.n493 B.n492 585
R441 B.n491 B.n30 585
R442 B.n490 B.n489 585
R443 B.n488 B.n31 585
R444 B.n487 B.n486 585
R445 B.n485 B.n32 585
R446 B.n484 B.n483 585
R447 B.n482 B.n33 585
R448 B.n481 B.n480 585
R449 B.n479 B.n34 585
R450 B.n478 B.n477 585
R451 B.n476 B.n35 585
R452 B.n475 B.n474 585
R453 B.n473 B.n39 585
R454 B.n472 B.n471 585
R455 B.n470 B.n40 585
R456 B.n469 B.n468 585
R457 B.n467 B.n41 585
R458 B.n466 B.n465 585
R459 B.n464 B.n42 585
R460 B.n462 B.n461 585
R461 B.n460 B.n45 585
R462 B.n459 B.n458 585
R463 B.n457 B.n46 585
R464 B.n456 B.n455 585
R465 B.n454 B.n47 585
R466 B.n453 B.n452 585
R467 B.n451 B.n48 585
R468 B.n450 B.n449 585
R469 B.n448 B.n49 585
R470 B.n447 B.n446 585
R471 B.n445 B.n50 585
R472 B.n444 B.n443 585
R473 B.n442 B.n51 585
R474 B.n500 B.n27 585
R475 B.n502 B.n501 585
R476 B.n503 B.n26 585
R477 B.n505 B.n504 585
R478 B.n506 B.n25 585
R479 B.n508 B.n507 585
R480 B.n509 B.n24 585
R481 B.n511 B.n510 585
R482 B.n512 B.n23 585
R483 B.n514 B.n513 585
R484 B.n515 B.n22 585
R485 B.n517 B.n516 585
R486 B.n518 B.n21 585
R487 B.n520 B.n519 585
R488 B.n521 B.n20 585
R489 B.n523 B.n522 585
R490 B.n524 B.n19 585
R491 B.n526 B.n525 585
R492 B.n527 B.n18 585
R493 B.n529 B.n528 585
R494 B.n530 B.n17 585
R495 B.n532 B.n531 585
R496 B.n533 B.n16 585
R497 B.n535 B.n534 585
R498 B.n536 B.n15 585
R499 B.n538 B.n537 585
R500 B.n539 B.n14 585
R501 B.n541 B.n540 585
R502 B.n542 B.n13 585
R503 B.n544 B.n543 585
R504 B.n545 B.n12 585
R505 B.n547 B.n546 585
R506 B.n548 B.n11 585
R507 B.n550 B.n549 585
R508 B.n551 B.n10 585
R509 B.n553 B.n552 585
R510 B.n554 B.n9 585
R511 B.n556 B.n555 585
R512 B.n557 B.n8 585
R513 B.n559 B.n558 585
R514 B.n560 B.n7 585
R515 B.n562 B.n561 585
R516 B.n563 B.n6 585
R517 B.n565 B.n564 585
R518 B.n566 B.n5 585
R519 B.n568 B.n567 585
R520 B.n569 B.n4 585
R521 B.n571 B.n570 585
R522 B.n572 B.n3 585
R523 B.n574 B.n573 585
R524 B.n575 B.n0 585
R525 B.n2 B.n1 585
R526 B.n150 B.n149 585
R527 B.n152 B.n151 585
R528 B.n153 B.n148 585
R529 B.n155 B.n154 585
R530 B.n156 B.n147 585
R531 B.n158 B.n157 585
R532 B.n159 B.n146 585
R533 B.n161 B.n160 585
R534 B.n162 B.n145 585
R535 B.n164 B.n163 585
R536 B.n165 B.n144 585
R537 B.n167 B.n166 585
R538 B.n168 B.n143 585
R539 B.n170 B.n169 585
R540 B.n171 B.n142 585
R541 B.n173 B.n172 585
R542 B.n174 B.n141 585
R543 B.n176 B.n175 585
R544 B.n177 B.n140 585
R545 B.n179 B.n178 585
R546 B.n180 B.n139 585
R547 B.n182 B.n181 585
R548 B.n183 B.n138 585
R549 B.n185 B.n184 585
R550 B.n186 B.n137 585
R551 B.n188 B.n187 585
R552 B.n189 B.n136 585
R553 B.n191 B.n190 585
R554 B.n192 B.n135 585
R555 B.n194 B.n193 585
R556 B.n195 B.n134 585
R557 B.n197 B.n196 585
R558 B.n198 B.n133 585
R559 B.n200 B.n199 585
R560 B.n201 B.n132 585
R561 B.n203 B.n202 585
R562 B.n204 B.n131 585
R563 B.n206 B.n205 585
R564 B.n207 B.n130 585
R565 B.n209 B.n208 585
R566 B.n210 B.n129 585
R567 B.n212 B.n211 585
R568 B.n213 B.n128 585
R569 B.n215 B.n214 585
R570 B.n216 B.n127 585
R571 B.n218 B.n217 585
R572 B.n219 B.n126 585
R573 B.n221 B.n220 585
R574 B.n222 B.n125 585
R575 B.n224 B.n223 585
R576 B.n223 B.n124 492.5
R577 B.n286 B.n285 492.5
R578 B.n442 B.n441 492.5
R579 B.n498 B.n27 492.5
R580 B.n111 B.t4 284.76
R581 B.n43 B.t11 284.76
R582 B.n244 B.t1 284.76
R583 B.n36 B.t8 284.76
R584 B.n577 B.n576 256.663
R585 B.n576 B.n575 235.042
R586 B.n576 B.n2 235.042
R587 B.n244 B.t0 232.637
R588 B.n111 B.t3 232.637
R589 B.n43 B.t9 232.637
R590 B.n36 B.t6 232.637
R591 B.n112 B.t5 227.548
R592 B.n44 B.t10 227.548
R593 B.n245 B.t2 227.548
R594 B.n37 B.t7 227.548
R595 B.n227 B.n124 163.367
R596 B.n228 B.n227 163.367
R597 B.n229 B.n228 163.367
R598 B.n229 B.n122 163.367
R599 B.n233 B.n122 163.367
R600 B.n234 B.n233 163.367
R601 B.n235 B.n234 163.367
R602 B.n235 B.n120 163.367
R603 B.n239 B.n120 163.367
R604 B.n240 B.n239 163.367
R605 B.n241 B.n240 163.367
R606 B.n241 B.n118 163.367
R607 B.n248 B.n118 163.367
R608 B.n249 B.n248 163.367
R609 B.n250 B.n249 163.367
R610 B.n250 B.n116 163.367
R611 B.n254 B.n116 163.367
R612 B.n255 B.n254 163.367
R613 B.n256 B.n255 163.367
R614 B.n256 B.n114 163.367
R615 B.n260 B.n114 163.367
R616 B.n261 B.n260 163.367
R617 B.n262 B.n261 163.367
R618 B.n262 B.n110 163.367
R619 B.n267 B.n110 163.367
R620 B.n268 B.n267 163.367
R621 B.n269 B.n268 163.367
R622 B.n269 B.n108 163.367
R623 B.n273 B.n108 163.367
R624 B.n274 B.n273 163.367
R625 B.n275 B.n274 163.367
R626 B.n275 B.n106 163.367
R627 B.n279 B.n106 163.367
R628 B.n280 B.n279 163.367
R629 B.n281 B.n280 163.367
R630 B.n281 B.n104 163.367
R631 B.n285 B.n104 163.367
R632 B.n441 B.n52 163.367
R633 B.n437 B.n52 163.367
R634 B.n437 B.n436 163.367
R635 B.n436 B.n435 163.367
R636 B.n435 B.n54 163.367
R637 B.n431 B.n54 163.367
R638 B.n431 B.n430 163.367
R639 B.n430 B.n429 163.367
R640 B.n429 B.n56 163.367
R641 B.n425 B.n56 163.367
R642 B.n425 B.n424 163.367
R643 B.n424 B.n423 163.367
R644 B.n423 B.n58 163.367
R645 B.n419 B.n58 163.367
R646 B.n419 B.n418 163.367
R647 B.n418 B.n417 163.367
R648 B.n417 B.n60 163.367
R649 B.n413 B.n60 163.367
R650 B.n413 B.n412 163.367
R651 B.n412 B.n411 163.367
R652 B.n411 B.n62 163.367
R653 B.n407 B.n62 163.367
R654 B.n407 B.n406 163.367
R655 B.n406 B.n405 163.367
R656 B.n405 B.n64 163.367
R657 B.n401 B.n64 163.367
R658 B.n401 B.n400 163.367
R659 B.n400 B.n399 163.367
R660 B.n399 B.n66 163.367
R661 B.n395 B.n66 163.367
R662 B.n395 B.n394 163.367
R663 B.n394 B.n393 163.367
R664 B.n393 B.n68 163.367
R665 B.n389 B.n68 163.367
R666 B.n389 B.n388 163.367
R667 B.n388 B.n387 163.367
R668 B.n387 B.n70 163.367
R669 B.n383 B.n70 163.367
R670 B.n383 B.n382 163.367
R671 B.n382 B.n381 163.367
R672 B.n381 B.n72 163.367
R673 B.n377 B.n72 163.367
R674 B.n377 B.n376 163.367
R675 B.n376 B.n375 163.367
R676 B.n375 B.n74 163.367
R677 B.n371 B.n74 163.367
R678 B.n371 B.n370 163.367
R679 B.n370 B.n369 163.367
R680 B.n369 B.n76 163.367
R681 B.n365 B.n76 163.367
R682 B.n365 B.n364 163.367
R683 B.n364 B.n363 163.367
R684 B.n363 B.n78 163.367
R685 B.n359 B.n78 163.367
R686 B.n359 B.n358 163.367
R687 B.n358 B.n357 163.367
R688 B.n357 B.n80 163.367
R689 B.n353 B.n80 163.367
R690 B.n353 B.n352 163.367
R691 B.n352 B.n351 163.367
R692 B.n351 B.n82 163.367
R693 B.n347 B.n82 163.367
R694 B.n347 B.n346 163.367
R695 B.n346 B.n345 163.367
R696 B.n345 B.n84 163.367
R697 B.n341 B.n84 163.367
R698 B.n341 B.n340 163.367
R699 B.n340 B.n339 163.367
R700 B.n339 B.n86 163.367
R701 B.n335 B.n86 163.367
R702 B.n335 B.n334 163.367
R703 B.n334 B.n333 163.367
R704 B.n333 B.n88 163.367
R705 B.n329 B.n88 163.367
R706 B.n329 B.n328 163.367
R707 B.n328 B.n327 163.367
R708 B.n327 B.n90 163.367
R709 B.n323 B.n90 163.367
R710 B.n323 B.n322 163.367
R711 B.n322 B.n321 163.367
R712 B.n321 B.n92 163.367
R713 B.n317 B.n92 163.367
R714 B.n317 B.n316 163.367
R715 B.n316 B.n315 163.367
R716 B.n315 B.n94 163.367
R717 B.n311 B.n94 163.367
R718 B.n311 B.n310 163.367
R719 B.n310 B.n309 163.367
R720 B.n309 B.n96 163.367
R721 B.n305 B.n96 163.367
R722 B.n305 B.n304 163.367
R723 B.n304 B.n303 163.367
R724 B.n303 B.n98 163.367
R725 B.n299 B.n98 163.367
R726 B.n299 B.n298 163.367
R727 B.n298 B.n297 163.367
R728 B.n297 B.n100 163.367
R729 B.n293 B.n100 163.367
R730 B.n293 B.n292 163.367
R731 B.n292 B.n291 163.367
R732 B.n291 B.n102 163.367
R733 B.n287 B.n102 163.367
R734 B.n287 B.n286 163.367
R735 B.n498 B.n497 163.367
R736 B.n497 B.n496 163.367
R737 B.n496 B.n29 163.367
R738 B.n492 B.n29 163.367
R739 B.n492 B.n491 163.367
R740 B.n491 B.n490 163.367
R741 B.n490 B.n31 163.367
R742 B.n486 B.n31 163.367
R743 B.n486 B.n485 163.367
R744 B.n485 B.n484 163.367
R745 B.n484 B.n33 163.367
R746 B.n480 B.n33 163.367
R747 B.n480 B.n479 163.367
R748 B.n479 B.n478 163.367
R749 B.n478 B.n35 163.367
R750 B.n474 B.n35 163.367
R751 B.n474 B.n473 163.367
R752 B.n473 B.n472 163.367
R753 B.n472 B.n40 163.367
R754 B.n468 B.n40 163.367
R755 B.n468 B.n467 163.367
R756 B.n467 B.n466 163.367
R757 B.n466 B.n42 163.367
R758 B.n461 B.n42 163.367
R759 B.n461 B.n460 163.367
R760 B.n460 B.n459 163.367
R761 B.n459 B.n46 163.367
R762 B.n455 B.n46 163.367
R763 B.n455 B.n454 163.367
R764 B.n454 B.n453 163.367
R765 B.n453 B.n48 163.367
R766 B.n449 B.n48 163.367
R767 B.n449 B.n448 163.367
R768 B.n448 B.n447 163.367
R769 B.n447 B.n50 163.367
R770 B.n443 B.n50 163.367
R771 B.n443 B.n442 163.367
R772 B.n502 B.n27 163.367
R773 B.n503 B.n502 163.367
R774 B.n504 B.n503 163.367
R775 B.n504 B.n25 163.367
R776 B.n508 B.n25 163.367
R777 B.n509 B.n508 163.367
R778 B.n510 B.n509 163.367
R779 B.n510 B.n23 163.367
R780 B.n514 B.n23 163.367
R781 B.n515 B.n514 163.367
R782 B.n516 B.n515 163.367
R783 B.n516 B.n21 163.367
R784 B.n520 B.n21 163.367
R785 B.n521 B.n520 163.367
R786 B.n522 B.n521 163.367
R787 B.n522 B.n19 163.367
R788 B.n526 B.n19 163.367
R789 B.n527 B.n526 163.367
R790 B.n528 B.n527 163.367
R791 B.n528 B.n17 163.367
R792 B.n532 B.n17 163.367
R793 B.n533 B.n532 163.367
R794 B.n534 B.n533 163.367
R795 B.n534 B.n15 163.367
R796 B.n538 B.n15 163.367
R797 B.n539 B.n538 163.367
R798 B.n540 B.n539 163.367
R799 B.n540 B.n13 163.367
R800 B.n544 B.n13 163.367
R801 B.n545 B.n544 163.367
R802 B.n546 B.n545 163.367
R803 B.n546 B.n11 163.367
R804 B.n550 B.n11 163.367
R805 B.n551 B.n550 163.367
R806 B.n552 B.n551 163.367
R807 B.n552 B.n9 163.367
R808 B.n556 B.n9 163.367
R809 B.n557 B.n556 163.367
R810 B.n558 B.n557 163.367
R811 B.n558 B.n7 163.367
R812 B.n562 B.n7 163.367
R813 B.n563 B.n562 163.367
R814 B.n564 B.n563 163.367
R815 B.n564 B.n5 163.367
R816 B.n568 B.n5 163.367
R817 B.n569 B.n568 163.367
R818 B.n570 B.n569 163.367
R819 B.n570 B.n3 163.367
R820 B.n574 B.n3 163.367
R821 B.n575 B.n574 163.367
R822 B.n150 B.n2 163.367
R823 B.n151 B.n150 163.367
R824 B.n151 B.n148 163.367
R825 B.n155 B.n148 163.367
R826 B.n156 B.n155 163.367
R827 B.n157 B.n156 163.367
R828 B.n157 B.n146 163.367
R829 B.n161 B.n146 163.367
R830 B.n162 B.n161 163.367
R831 B.n163 B.n162 163.367
R832 B.n163 B.n144 163.367
R833 B.n167 B.n144 163.367
R834 B.n168 B.n167 163.367
R835 B.n169 B.n168 163.367
R836 B.n169 B.n142 163.367
R837 B.n173 B.n142 163.367
R838 B.n174 B.n173 163.367
R839 B.n175 B.n174 163.367
R840 B.n175 B.n140 163.367
R841 B.n179 B.n140 163.367
R842 B.n180 B.n179 163.367
R843 B.n181 B.n180 163.367
R844 B.n181 B.n138 163.367
R845 B.n185 B.n138 163.367
R846 B.n186 B.n185 163.367
R847 B.n187 B.n186 163.367
R848 B.n187 B.n136 163.367
R849 B.n191 B.n136 163.367
R850 B.n192 B.n191 163.367
R851 B.n193 B.n192 163.367
R852 B.n193 B.n134 163.367
R853 B.n197 B.n134 163.367
R854 B.n198 B.n197 163.367
R855 B.n199 B.n198 163.367
R856 B.n199 B.n132 163.367
R857 B.n203 B.n132 163.367
R858 B.n204 B.n203 163.367
R859 B.n205 B.n204 163.367
R860 B.n205 B.n130 163.367
R861 B.n209 B.n130 163.367
R862 B.n210 B.n209 163.367
R863 B.n211 B.n210 163.367
R864 B.n211 B.n128 163.367
R865 B.n215 B.n128 163.367
R866 B.n216 B.n215 163.367
R867 B.n217 B.n216 163.367
R868 B.n217 B.n126 163.367
R869 B.n221 B.n126 163.367
R870 B.n222 B.n221 163.367
R871 B.n223 B.n222 163.367
R872 B.n246 B.n245 59.5399
R873 B.n264 B.n112 59.5399
R874 B.n463 B.n44 59.5399
R875 B.n38 B.n37 59.5399
R876 B.n245 B.n244 57.2126
R877 B.n112 B.n111 57.2126
R878 B.n44 B.n43 57.2126
R879 B.n37 B.n36 57.2126
R880 B.n500 B.n499 32.0005
R881 B.n440 B.n51 32.0005
R882 B.n284 B.n103 32.0005
R883 B.n225 B.n224 32.0005
R884 B B.n577 18.0485
R885 B.n501 B.n500 10.6151
R886 B.n501 B.n26 10.6151
R887 B.n505 B.n26 10.6151
R888 B.n506 B.n505 10.6151
R889 B.n507 B.n506 10.6151
R890 B.n507 B.n24 10.6151
R891 B.n511 B.n24 10.6151
R892 B.n512 B.n511 10.6151
R893 B.n513 B.n512 10.6151
R894 B.n513 B.n22 10.6151
R895 B.n517 B.n22 10.6151
R896 B.n518 B.n517 10.6151
R897 B.n519 B.n518 10.6151
R898 B.n519 B.n20 10.6151
R899 B.n523 B.n20 10.6151
R900 B.n524 B.n523 10.6151
R901 B.n525 B.n524 10.6151
R902 B.n525 B.n18 10.6151
R903 B.n529 B.n18 10.6151
R904 B.n530 B.n529 10.6151
R905 B.n531 B.n530 10.6151
R906 B.n531 B.n16 10.6151
R907 B.n535 B.n16 10.6151
R908 B.n536 B.n535 10.6151
R909 B.n537 B.n536 10.6151
R910 B.n537 B.n14 10.6151
R911 B.n541 B.n14 10.6151
R912 B.n542 B.n541 10.6151
R913 B.n543 B.n542 10.6151
R914 B.n543 B.n12 10.6151
R915 B.n547 B.n12 10.6151
R916 B.n548 B.n547 10.6151
R917 B.n549 B.n548 10.6151
R918 B.n549 B.n10 10.6151
R919 B.n553 B.n10 10.6151
R920 B.n554 B.n553 10.6151
R921 B.n555 B.n554 10.6151
R922 B.n555 B.n8 10.6151
R923 B.n559 B.n8 10.6151
R924 B.n560 B.n559 10.6151
R925 B.n561 B.n560 10.6151
R926 B.n561 B.n6 10.6151
R927 B.n565 B.n6 10.6151
R928 B.n566 B.n565 10.6151
R929 B.n567 B.n566 10.6151
R930 B.n567 B.n4 10.6151
R931 B.n571 B.n4 10.6151
R932 B.n572 B.n571 10.6151
R933 B.n573 B.n572 10.6151
R934 B.n573 B.n0 10.6151
R935 B.n499 B.n28 10.6151
R936 B.n495 B.n28 10.6151
R937 B.n495 B.n494 10.6151
R938 B.n494 B.n493 10.6151
R939 B.n493 B.n30 10.6151
R940 B.n489 B.n30 10.6151
R941 B.n489 B.n488 10.6151
R942 B.n488 B.n487 10.6151
R943 B.n487 B.n32 10.6151
R944 B.n483 B.n32 10.6151
R945 B.n483 B.n482 10.6151
R946 B.n482 B.n481 10.6151
R947 B.n481 B.n34 10.6151
R948 B.n477 B.n476 10.6151
R949 B.n476 B.n475 10.6151
R950 B.n475 B.n39 10.6151
R951 B.n471 B.n39 10.6151
R952 B.n471 B.n470 10.6151
R953 B.n470 B.n469 10.6151
R954 B.n469 B.n41 10.6151
R955 B.n465 B.n41 10.6151
R956 B.n465 B.n464 10.6151
R957 B.n462 B.n45 10.6151
R958 B.n458 B.n45 10.6151
R959 B.n458 B.n457 10.6151
R960 B.n457 B.n456 10.6151
R961 B.n456 B.n47 10.6151
R962 B.n452 B.n47 10.6151
R963 B.n452 B.n451 10.6151
R964 B.n451 B.n450 10.6151
R965 B.n450 B.n49 10.6151
R966 B.n446 B.n49 10.6151
R967 B.n446 B.n445 10.6151
R968 B.n445 B.n444 10.6151
R969 B.n444 B.n51 10.6151
R970 B.n440 B.n439 10.6151
R971 B.n439 B.n438 10.6151
R972 B.n438 B.n53 10.6151
R973 B.n434 B.n53 10.6151
R974 B.n434 B.n433 10.6151
R975 B.n433 B.n432 10.6151
R976 B.n432 B.n55 10.6151
R977 B.n428 B.n55 10.6151
R978 B.n428 B.n427 10.6151
R979 B.n427 B.n426 10.6151
R980 B.n426 B.n57 10.6151
R981 B.n422 B.n57 10.6151
R982 B.n422 B.n421 10.6151
R983 B.n421 B.n420 10.6151
R984 B.n420 B.n59 10.6151
R985 B.n416 B.n59 10.6151
R986 B.n416 B.n415 10.6151
R987 B.n415 B.n414 10.6151
R988 B.n414 B.n61 10.6151
R989 B.n410 B.n61 10.6151
R990 B.n410 B.n409 10.6151
R991 B.n409 B.n408 10.6151
R992 B.n408 B.n63 10.6151
R993 B.n404 B.n63 10.6151
R994 B.n404 B.n403 10.6151
R995 B.n403 B.n402 10.6151
R996 B.n402 B.n65 10.6151
R997 B.n398 B.n65 10.6151
R998 B.n398 B.n397 10.6151
R999 B.n397 B.n396 10.6151
R1000 B.n396 B.n67 10.6151
R1001 B.n392 B.n67 10.6151
R1002 B.n392 B.n391 10.6151
R1003 B.n391 B.n390 10.6151
R1004 B.n390 B.n69 10.6151
R1005 B.n386 B.n69 10.6151
R1006 B.n386 B.n385 10.6151
R1007 B.n385 B.n384 10.6151
R1008 B.n384 B.n71 10.6151
R1009 B.n380 B.n71 10.6151
R1010 B.n380 B.n379 10.6151
R1011 B.n379 B.n378 10.6151
R1012 B.n378 B.n73 10.6151
R1013 B.n374 B.n73 10.6151
R1014 B.n374 B.n373 10.6151
R1015 B.n373 B.n372 10.6151
R1016 B.n372 B.n75 10.6151
R1017 B.n368 B.n75 10.6151
R1018 B.n368 B.n367 10.6151
R1019 B.n367 B.n366 10.6151
R1020 B.n366 B.n77 10.6151
R1021 B.n362 B.n77 10.6151
R1022 B.n362 B.n361 10.6151
R1023 B.n361 B.n360 10.6151
R1024 B.n360 B.n79 10.6151
R1025 B.n356 B.n79 10.6151
R1026 B.n356 B.n355 10.6151
R1027 B.n355 B.n354 10.6151
R1028 B.n354 B.n81 10.6151
R1029 B.n350 B.n81 10.6151
R1030 B.n350 B.n349 10.6151
R1031 B.n349 B.n348 10.6151
R1032 B.n348 B.n83 10.6151
R1033 B.n344 B.n83 10.6151
R1034 B.n344 B.n343 10.6151
R1035 B.n343 B.n342 10.6151
R1036 B.n342 B.n85 10.6151
R1037 B.n338 B.n85 10.6151
R1038 B.n338 B.n337 10.6151
R1039 B.n337 B.n336 10.6151
R1040 B.n336 B.n87 10.6151
R1041 B.n332 B.n87 10.6151
R1042 B.n332 B.n331 10.6151
R1043 B.n331 B.n330 10.6151
R1044 B.n330 B.n89 10.6151
R1045 B.n326 B.n89 10.6151
R1046 B.n326 B.n325 10.6151
R1047 B.n325 B.n324 10.6151
R1048 B.n324 B.n91 10.6151
R1049 B.n320 B.n91 10.6151
R1050 B.n320 B.n319 10.6151
R1051 B.n319 B.n318 10.6151
R1052 B.n318 B.n93 10.6151
R1053 B.n314 B.n93 10.6151
R1054 B.n314 B.n313 10.6151
R1055 B.n313 B.n312 10.6151
R1056 B.n312 B.n95 10.6151
R1057 B.n308 B.n95 10.6151
R1058 B.n308 B.n307 10.6151
R1059 B.n307 B.n306 10.6151
R1060 B.n306 B.n97 10.6151
R1061 B.n302 B.n97 10.6151
R1062 B.n302 B.n301 10.6151
R1063 B.n301 B.n300 10.6151
R1064 B.n300 B.n99 10.6151
R1065 B.n296 B.n99 10.6151
R1066 B.n296 B.n295 10.6151
R1067 B.n295 B.n294 10.6151
R1068 B.n294 B.n101 10.6151
R1069 B.n290 B.n101 10.6151
R1070 B.n290 B.n289 10.6151
R1071 B.n289 B.n288 10.6151
R1072 B.n288 B.n103 10.6151
R1073 B.n149 B.n1 10.6151
R1074 B.n152 B.n149 10.6151
R1075 B.n153 B.n152 10.6151
R1076 B.n154 B.n153 10.6151
R1077 B.n154 B.n147 10.6151
R1078 B.n158 B.n147 10.6151
R1079 B.n159 B.n158 10.6151
R1080 B.n160 B.n159 10.6151
R1081 B.n160 B.n145 10.6151
R1082 B.n164 B.n145 10.6151
R1083 B.n165 B.n164 10.6151
R1084 B.n166 B.n165 10.6151
R1085 B.n166 B.n143 10.6151
R1086 B.n170 B.n143 10.6151
R1087 B.n171 B.n170 10.6151
R1088 B.n172 B.n171 10.6151
R1089 B.n172 B.n141 10.6151
R1090 B.n176 B.n141 10.6151
R1091 B.n177 B.n176 10.6151
R1092 B.n178 B.n177 10.6151
R1093 B.n178 B.n139 10.6151
R1094 B.n182 B.n139 10.6151
R1095 B.n183 B.n182 10.6151
R1096 B.n184 B.n183 10.6151
R1097 B.n184 B.n137 10.6151
R1098 B.n188 B.n137 10.6151
R1099 B.n189 B.n188 10.6151
R1100 B.n190 B.n189 10.6151
R1101 B.n190 B.n135 10.6151
R1102 B.n194 B.n135 10.6151
R1103 B.n195 B.n194 10.6151
R1104 B.n196 B.n195 10.6151
R1105 B.n196 B.n133 10.6151
R1106 B.n200 B.n133 10.6151
R1107 B.n201 B.n200 10.6151
R1108 B.n202 B.n201 10.6151
R1109 B.n202 B.n131 10.6151
R1110 B.n206 B.n131 10.6151
R1111 B.n207 B.n206 10.6151
R1112 B.n208 B.n207 10.6151
R1113 B.n208 B.n129 10.6151
R1114 B.n212 B.n129 10.6151
R1115 B.n213 B.n212 10.6151
R1116 B.n214 B.n213 10.6151
R1117 B.n214 B.n127 10.6151
R1118 B.n218 B.n127 10.6151
R1119 B.n219 B.n218 10.6151
R1120 B.n220 B.n219 10.6151
R1121 B.n220 B.n125 10.6151
R1122 B.n224 B.n125 10.6151
R1123 B.n226 B.n225 10.6151
R1124 B.n226 B.n123 10.6151
R1125 B.n230 B.n123 10.6151
R1126 B.n231 B.n230 10.6151
R1127 B.n232 B.n231 10.6151
R1128 B.n232 B.n121 10.6151
R1129 B.n236 B.n121 10.6151
R1130 B.n237 B.n236 10.6151
R1131 B.n238 B.n237 10.6151
R1132 B.n238 B.n119 10.6151
R1133 B.n242 B.n119 10.6151
R1134 B.n243 B.n242 10.6151
R1135 B.n247 B.n243 10.6151
R1136 B.n251 B.n117 10.6151
R1137 B.n252 B.n251 10.6151
R1138 B.n253 B.n252 10.6151
R1139 B.n253 B.n115 10.6151
R1140 B.n257 B.n115 10.6151
R1141 B.n258 B.n257 10.6151
R1142 B.n259 B.n258 10.6151
R1143 B.n259 B.n113 10.6151
R1144 B.n263 B.n113 10.6151
R1145 B.n266 B.n265 10.6151
R1146 B.n266 B.n109 10.6151
R1147 B.n270 B.n109 10.6151
R1148 B.n271 B.n270 10.6151
R1149 B.n272 B.n271 10.6151
R1150 B.n272 B.n107 10.6151
R1151 B.n276 B.n107 10.6151
R1152 B.n277 B.n276 10.6151
R1153 B.n278 B.n277 10.6151
R1154 B.n278 B.n105 10.6151
R1155 B.n282 B.n105 10.6151
R1156 B.n283 B.n282 10.6151
R1157 B.n284 B.n283 10.6151
R1158 B.n38 B.n34 9.36635
R1159 B.n463 B.n462 9.36635
R1160 B.n247 B.n246 9.36635
R1161 B.n265 B.n264 9.36635
R1162 B.n577 B.n0 8.11757
R1163 B.n577 B.n1 8.11757
R1164 B.n477 B.n38 1.24928
R1165 B.n464 B.n463 1.24928
R1166 B.n246 B.n117 1.24928
R1167 B.n264 B.n263 1.24928
R1168 VN.n55 VN.n29 161.3
R1169 VN.n54 VN.n53 161.3
R1170 VN.n52 VN.n30 161.3
R1171 VN.n51 VN.n50 161.3
R1172 VN.n49 VN.n31 161.3
R1173 VN.n48 VN.n47 161.3
R1174 VN.n46 VN.n45 161.3
R1175 VN.n44 VN.n33 161.3
R1176 VN.n43 VN.n42 161.3
R1177 VN.n41 VN.n34 161.3
R1178 VN.n40 VN.n39 161.3
R1179 VN.n38 VN.n35 161.3
R1180 VN.n26 VN.n0 161.3
R1181 VN.n25 VN.n24 161.3
R1182 VN.n23 VN.n1 161.3
R1183 VN.n22 VN.n21 161.3
R1184 VN.n20 VN.n2 161.3
R1185 VN.n19 VN.n18 161.3
R1186 VN.n17 VN.n16 161.3
R1187 VN.n15 VN.n4 161.3
R1188 VN.n14 VN.n13 161.3
R1189 VN.n12 VN.n5 161.3
R1190 VN.n11 VN.n10 161.3
R1191 VN.n9 VN.n6 161.3
R1192 VN.n28 VN.n27 102.192
R1193 VN.n57 VN.n56 102.192
R1194 VN.n8 VN.n7 61.3525
R1195 VN.n37 VN.n36 61.3525
R1196 VN.n7 VN.t2 57.7507
R1197 VN.n36 VN.t3 57.7507
R1198 VN.n14 VN.n5 56.5193
R1199 VN.n21 VN.n1 56.5193
R1200 VN.n43 VN.n34 56.5193
R1201 VN.n50 VN.n30 56.5193
R1202 VN VN.n57 44.2027
R1203 VN.n8 VN.t0 24.5604
R1204 VN.n3 VN.t7 24.5604
R1205 VN.n27 VN.t1 24.5604
R1206 VN.n37 VN.t5 24.5604
R1207 VN.n32 VN.t4 24.5604
R1208 VN.n56 VN.t6 24.5604
R1209 VN.n10 VN.n9 24.4675
R1210 VN.n10 VN.n5 24.4675
R1211 VN.n15 VN.n14 24.4675
R1212 VN.n16 VN.n15 24.4675
R1213 VN.n20 VN.n19 24.4675
R1214 VN.n21 VN.n20 24.4675
R1215 VN.n25 VN.n1 24.4675
R1216 VN.n26 VN.n25 24.4675
R1217 VN.n39 VN.n34 24.4675
R1218 VN.n39 VN.n38 24.4675
R1219 VN.n50 VN.n49 24.4675
R1220 VN.n49 VN.n48 24.4675
R1221 VN.n45 VN.n44 24.4675
R1222 VN.n44 VN.n43 24.4675
R1223 VN.n55 VN.n54 24.4675
R1224 VN.n54 VN.n30 24.4675
R1225 VN.n19 VN.n3 13.4574
R1226 VN.n48 VN.n32 13.4574
R1227 VN.n9 VN.n8 11.0107
R1228 VN.n16 VN.n3 11.0107
R1229 VN.n38 VN.n37 11.0107
R1230 VN.n45 VN.n32 11.0107
R1231 VN.n27 VN.n26 8.56395
R1232 VN.n56 VN.n55 8.56395
R1233 VN.n36 VN.n35 6.94033
R1234 VN.n7 VN.n6 6.94033
R1235 VN.n57 VN.n29 0.278367
R1236 VN.n28 VN.n0 0.278367
R1237 VN.n53 VN.n29 0.189894
R1238 VN.n53 VN.n52 0.189894
R1239 VN.n52 VN.n51 0.189894
R1240 VN.n51 VN.n31 0.189894
R1241 VN.n47 VN.n31 0.189894
R1242 VN.n47 VN.n46 0.189894
R1243 VN.n46 VN.n33 0.189894
R1244 VN.n42 VN.n33 0.189894
R1245 VN.n42 VN.n41 0.189894
R1246 VN.n41 VN.n40 0.189894
R1247 VN.n40 VN.n35 0.189894
R1248 VN.n11 VN.n6 0.189894
R1249 VN.n12 VN.n11 0.189894
R1250 VN.n13 VN.n12 0.189894
R1251 VN.n13 VN.n4 0.189894
R1252 VN.n17 VN.n4 0.189894
R1253 VN.n18 VN.n17 0.189894
R1254 VN.n18 VN.n2 0.189894
R1255 VN.n22 VN.n2 0.189894
R1256 VN.n23 VN.n22 0.189894
R1257 VN.n24 VN.n23 0.189894
R1258 VN.n24 VN.n0 0.189894
R1259 VN VN.n28 0.153454
R1260 VDD2.n2 VDD2.n1 152.6
R1261 VDD2.n2 VDD2.n0 152.6
R1262 VDD2 VDD2.n5 152.596
R1263 VDD2.n4 VDD2.n3 151.383
R1264 VDD2.n4 VDD2.n2 37.461
R1265 VDD2.n5 VDD2.t2 12.1747
R1266 VDD2.n5 VDD2.t4 12.1747
R1267 VDD2.n3 VDD2.t1 12.1747
R1268 VDD2.n3 VDD2.t3 12.1747
R1269 VDD2.n1 VDD2.t0 12.1747
R1270 VDD2.n1 VDD2.t6 12.1747
R1271 VDD2.n0 VDD2.t5 12.1747
R1272 VDD2.n0 VDD2.t7 12.1747
R1273 VDD2 VDD2.n4 1.33024
C0 VP VN 5.96555f
C1 VP w_n3920_n1502# 8.31962f
C2 B VDD2 1.4992f
C3 VP VTAIL 3.37032f
C4 VP VDD2 0.528037f
C5 VN VDD1 0.157077f
C6 w_n3920_n1502# VDD1 1.7101f
C7 VTAIL VDD1 4.95551f
C8 w_n3920_n1502# VN 7.81356f
C9 B VP 1.98411f
C10 VTAIL VN 3.35622f
C11 w_n3920_n1502# VTAIL 2.08592f
C12 VDD2 VDD1 1.78853f
C13 VDD2 VN 2.28706f
C14 w_n3920_n1502# VDD2 1.82506f
C15 B VDD1 1.4023f
C16 VDD2 VTAIL 5.01006f
C17 B VN 1.13134f
C18 B w_n3920_n1502# 7.56714f
C19 B VTAIL 1.85501f
C20 VP VDD1 2.65547f
C21 VDD2 VSUBS 1.415172f
C22 VDD1 VSUBS 2.092003f
C23 VTAIL VSUBS 0.58581f
C24 VN VSUBS 6.70914f
C25 VP VSUBS 3.008925f
C26 B VSUBS 3.983136f
C27 w_n3920_n1502# VSUBS 74.7466f
C28 VDD2.t5 VSUBS 0.05097f
C29 VDD2.t7 VSUBS 0.05097f
C30 VDD2.n0 VSUBS 0.248658f
C31 VDD2.t0 VSUBS 0.05097f
C32 VDD2.t6 VSUBS 0.05097f
C33 VDD2.n1 VSUBS 0.248658f
C34 VDD2.n2 VSUBS 2.84525f
C35 VDD2.t1 VSUBS 0.05097f
C36 VDD2.t3 VSUBS 0.05097f
C37 VDD2.n3 VSUBS 0.243833f
C38 VDD2.n4 VSUBS 2.25929f
C39 VDD2.t2 VSUBS 0.05097f
C40 VDD2.t4 VSUBS 0.05097f
C41 VDD2.n5 VSUBS 0.248642f
C42 VN.n0 VSUBS 0.063771f
C43 VN.t1 VSUBS 0.829875f
C44 VN.n1 VSUBS 0.07735f
C45 VN.n2 VSUBS 0.04837f
C46 VN.t7 VSUBS 0.829875f
C47 VN.n3 VSUBS 0.360589f
C48 VN.n4 VSUBS 0.04837f
C49 VN.n5 VSUBS 0.070611f
C50 VN.n6 VSUBS 0.468504f
C51 VN.t0 VSUBS 0.829875f
C52 VN.t2 VSUBS 1.2097f
C53 VN.n7 VSUBS 0.48323f
C54 VN.n8 VSUBS 0.498377f
C55 VN.n9 VSUBS 0.065668f
C56 VN.n10 VSUBS 0.090149f
C57 VN.n11 VSUBS 0.04837f
C58 VN.n12 VSUBS 0.04837f
C59 VN.n13 VSUBS 0.04837f
C60 VN.n14 VSUBS 0.070611f
C61 VN.n15 VSUBS 0.090149f
C62 VN.n16 VSUBS 0.065668f
C63 VN.n17 VSUBS 0.04837f
C64 VN.n18 VSUBS 0.04837f
C65 VN.n19 VSUBS 0.070119f
C66 VN.n20 VSUBS 0.090149f
C67 VN.n21 VSUBS 0.063872f
C68 VN.n22 VSUBS 0.04837f
C69 VN.n23 VSUBS 0.04837f
C70 VN.n24 VSUBS 0.04837f
C71 VN.n25 VSUBS 0.090149f
C72 VN.n26 VSUBS 0.061217f
C73 VN.n27 VSUBS 0.520321f
C74 VN.n28 VSUBS 0.080752f
C75 VN.n29 VSUBS 0.063771f
C76 VN.t6 VSUBS 0.829875f
C77 VN.n30 VSUBS 0.07735f
C78 VN.n31 VSUBS 0.04837f
C79 VN.t4 VSUBS 0.829875f
C80 VN.n32 VSUBS 0.360589f
C81 VN.n33 VSUBS 0.04837f
C82 VN.n34 VSUBS 0.070611f
C83 VN.n35 VSUBS 0.468504f
C84 VN.t5 VSUBS 0.829875f
C85 VN.t3 VSUBS 1.2097f
C86 VN.n36 VSUBS 0.48323f
C87 VN.n37 VSUBS 0.498377f
C88 VN.n38 VSUBS 0.065668f
C89 VN.n39 VSUBS 0.090149f
C90 VN.n40 VSUBS 0.04837f
C91 VN.n41 VSUBS 0.04837f
C92 VN.n42 VSUBS 0.04837f
C93 VN.n43 VSUBS 0.070611f
C94 VN.n44 VSUBS 0.090149f
C95 VN.n45 VSUBS 0.065668f
C96 VN.n46 VSUBS 0.04837f
C97 VN.n47 VSUBS 0.04837f
C98 VN.n48 VSUBS 0.070119f
C99 VN.n49 VSUBS 0.090149f
C100 VN.n50 VSUBS 0.063872f
C101 VN.n51 VSUBS 0.04837f
C102 VN.n52 VSUBS 0.04837f
C103 VN.n53 VSUBS 0.04837f
C104 VN.n54 VSUBS 0.090149f
C105 VN.n55 VSUBS 0.061217f
C106 VN.n56 VSUBS 0.520321f
C107 VN.n57 VSUBS 2.23924f
C108 B.n0 VSUBS 0.007032f
C109 B.n1 VSUBS 0.007032f
C110 B.n2 VSUBS 0.010399f
C111 B.n3 VSUBS 0.007969f
C112 B.n4 VSUBS 0.007969f
C113 B.n5 VSUBS 0.007969f
C114 B.n6 VSUBS 0.007969f
C115 B.n7 VSUBS 0.007969f
C116 B.n8 VSUBS 0.007969f
C117 B.n9 VSUBS 0.007969f
C118 B.n10 VSUBS 0.007969f
C119 B.n11 VSUBS 0.007969f
C120 B.n12 VSUBS 0.007969f
C121 B.n13 VSUBS 0.007969f
C122 B.n14 VSUBS 0.007969f
C123 B.n15 VSUBS 0.007969f
C124 B.n16 VSUBS 0.007969f
C125 B.n17 VSUBS 0.007969f
C126 B.n18 VSUBS 0.007969f
C127 B.n19 VSUBS 0.007969f
C128 B.n20 VSUBS 0.007969f
C129 B.n21 VSUBS 0.007969f
C130 B.n22 VSUBS 0.007969f
C131 B.n23 VSUBS 0.007969f
C132 B.n24 VSUBS 0.007969f
C133 B.n25 VSUBS 0.007969f
C134 B.n26 VSUBS 0.007969f
C135 B.n27 VSUBS 0.017919f
C136 B.n28 VSUBS 0.007969f
C137 B.n29 VSUBS 0.007969f
C138 B.n30 VSUBS 0.007969f
C139 B.n31 VSUBS 0.007969f
C140 B.n32 VSUBS 0.007969f
C141 B.n33 VSUBS 0.007969f
C142 B.n34 VSUBS 0.0075f
C143 B.n35 VSUBS 0.007969f
C144 B.t7 VSUBS 0.047402f
C145 B.t8 VSUBS 0.064327f
C146 B.t6 VSUBS 0.388846f
C147 B.n36 VSUBS 0.112429f
C148 B.n37 VSUBS 0.095605f
C149 B.n38 VSUBS 0.018464f
C150 B.n39 VSUBS 0.007969f
C151 B.n40 VSUBS 0.007969f
C152 B.n41 VSUBS 0.007969f
C153 B.n42 VSUBS 0.007969f
C154 B.t10 VSUBS 0.047402f
C155 B.t11 VSUBS 0.064327f
C156 B.t9 VSUBS 0.388846f
C157 B.n43 VSUBS 0.112428f
C158 B.n44 VSUBS 0.095605f
C159 B.n45 VSUBS 0.007969f
C160 B.n46 VSUBS 0.007969f
C161 B.n47 VSUBS 0.007969f
C162 B.n48 VSUBS 0.007969f
C163 B.n49 VSUBS 0.007969f
C164 B.n50 VSUBS 0.007969f
C165 B.n51 VSUBS 0.01888f
C166 B.n52 VSUBS 0.007969f
C167 B.n53 VSUBS 0.007969f
C168 B.n54 VSUBS 0.007969f
C169 B.n55 VSUBS 0.007969f
C170 B.n56 VSUBS 0.007969f
C171 B.n57 VSUBS 0.007969f
C172 B.n58 VSUBS 0.007969f
C173 B.n59 VSUBS 0.007969f
C174 B.n60 VSUBS 0.007969f
C175 B.n61 VSUBS 0.007969f
C176 B.n62 VSUBS 0.007969f
C177 B.n63 VSUBS 0.007969f
C178 B.n64 VSUBS 0.007969f
C179 B.n65 VSUBS 0.007969f
C180 B.n66 VSUBS 0.007969f
C181 B.n67 VSUBS 0.007969f
C182 B.n68 VSUBS 0.007969f
C183 B.n69 VSUBS 0.007969f
C184 B.n70 VSUBS 0.007969f
C185 B.n71 VSUBS 0.007969f
C186 B.n72 VSUBS 0.007969f
C187 B.n73 VSUBS 0.007969f
C188 B.n74 VSUBS 0.007969f
C189 B.n75 VSUBS 0.007969f
C190 B.n76 VSUBS 0.007969f
C191 B.n77 VSUBS 0.007969f
C192 B.n78 VSUBS 0.007969f
C193 B.n79 VSUBS 0.007969f
C194 B.n80 VSUBS 0.007969f
C195 B.n81 VSUBS 0.007969f
C196 B.n82 VSUBS 0.007969f
C197 B.n83 VSUBS 0.007969f
C198 B.n84 VSUBS 0.007969f
C199 B.n85 VSUBS 0.007969f
C200 B.n86 VSUBS 0.007969f
C201 B.n87 VSUBS 0.007969f
C202 B.n88 VSUBS 0.007969f
C203 B.n89 VSUBS 0.007969f
C204 B.n90 VSUBS 0.007969f
C205 B.n91 VSUBS 0.007969f
C206 B.n92 VSUBS 0.007969f
C207 B.n93 VSUBS 0.007969f
C208 B.n94 VSUBS 0.007969f
C209 B.n95 VSUBS 0.007969f
C210 B.n96 VSUBS 0.007969f
C211 B.n97 VSUBS 0.007969f
C212 B.n98 VSUBS 0.007969f
C213 B.n99 VSUBS 0.007969f
C214 B.n100 VSUBS 0.007969f
C215 B.n101 VSUBS 0.007969f
C216 B.n102 VSUBS 0.007969f
C217 B.n103 VSUBS 0.01888f
C218 B.n104 VSUBS 0.007969f
C219 B.n105 VSUBS 0.007969f
C220 B.n106 VSUBS 0.007969f
C221 B.n107 VSUBS 0.007969f
C222 B.n108 VSUBS 0.007969f
C223 B.n109 VSUBS 0.007969f
C224 B.n110 VSUBS 0.007969f
C225 B.t5 VSUBS 0.047402f
C226 B.t4 VSUBS 0.064327f
C227 B.t3 VSUBS 0.388846f
C228 B.n111 VSUBS 0.112428f
C229 B.n112 VSUBS 0.095605f
C230 B.n113 VSUBS 0.007969f
C231 B.n114 VSUBS 0.007969f
C232 B.n115 VSUBS 0.007969f
C233 B.n116 VSUBS 0.007969f
C234 B.n117 VSUBS 0.004453f
C235 B.n118 VSUBS 0.007969f
C236 B.n119 VSUBS 0.007969f
C237 B.n120 VSUBS 0.007969f
C238 B.n121 VSUBS 0.007969f
C239 B.n122 VSUBS 0.007969f
C240 B.n123 VSUBS 0.007969f
C241 B.n124 VSUBS 0.01888f
C242 B.n125 VSUBS 0.007969f
C243 B.n126 VSUBS 0.007969f
C244 B.n127 VSUBS 0.007969f
C245 B.n128 VSUBS 0.007969f
C246 B.n129 VSUBS 0.007969f
C247 B.n130 VSUBS 0.007969f
C248 B.n131 VSUBS 0.007969f
C249 B.n132 VSUBS 0.007969f
C250 B.n133 VSUBS 0.007969f
C251 B.n134 VSUBS 0.007969f
C252 B.n135 VSUBS 0.007969f
C253 B.n136 VSUBS 0.007969f
C254 B.n137 VSUBS 0.007969f
C255 B.n138 VSUBS 0.007969f
C256 B.n139 VSUBS 0.007969f
C257 B.n140 VSUBS 0.007969f
C258 B.n141 VSUBS 0.007969f
C259 B.n142 VSUBS 0.007969f
C260 B.n143 VSUBS 0.007969f
C261 B.n144 VSUBS 0.007969f
C262 B.n145 VSUBS 0.007969f
C263 B.n146 VSUBS 0.007969f
C264 B.n147 VSUBS 0.007969f
C265 B.n148 VSUBS 0.007969f
C266 B.n149 VSUBS 0.007969f
C267 B.n150 VSUBS 0.007969f
C268 B.n151 VSUBS 0.007969f
C269 B.n152 VSUBS 0.007969f
C270 B.n153 VSUBS 0.007969f
C271 B.n154 VSUBS 0.007969f
C272 B.n155 VSUBS 0.007969f
C273 B.n156 VSUBS 0.007969f
C274 B.n157 VSUBS 0.007969f
C275 B.n158 VSUBS 0.007969f
C276 B.n159 VSUBS 0.007969f
C277 B.n160 VSUBS 0.007969f
C278 B.n161 VSUBS 0.007969f
C279 B.n162 VSUBS 0.007969f
C280 B.n163 VSUBS 0.007969f
C281 B.n164 VSUBS 0.007969f
C282 B.n165 VSUBS 0.007969f
C283 B.n166 VSUBS 0.007969f
C284 B.n167 VSUBS 0.007969f
C285 B.n168 VSUBS 0.007969f
C286 B.n169 VSUBS 0.007969f
C287 B.n170 VSUBS 0.007969f
C288 B.n171 VSUBS 0.007969f
C289 B.n172 VSUBS 0.007969f
C290 B.n173 VSUBS 0.007969f
C291 B.n174 VSUBS 0.007969f
C292 B.n175 VSUBS 0.007969f
C293 B.n176 VSUBS 0.007969f
C294 B.n177 VSUBS 0.007969f
C295 B.n178 VSUBS 0.007969f
C296 B.n179 VSUBS 0.007969f
C297 B.n180 VSUBS 0.007969f
C298 B.n181 VSUBS 0.007969f
C299 B.n182 VSUBS 0.007969f
C300 B.n183 VSUBS 0.007969f
C301 B.n184 VSUBS 0.007969f
C302 B.n185 VSUBS 0.007969f
C303 B.n186 VSUBS 0.007969f
C304 B.n187 VSUBS 0.007969f
C305 B.n188 VSUBS 0.007969f
C306 B.n189 VSUBS 0.007969f
C307 B.n190 VSUBS 0.007969f
C308 B.n191 VSUBS 0.007969f
C309 B.n192 VSUBS 0.007969f
C310 B.n193 VSUBS 0.007969f
C311 B.n194 VSUBS 0.007969f
C312 B.n195 VSUBS 0.007969f
C313 B.n196 VSUBS 0.007969f
C314 B.n197 VSUBS 0.007969f
C315 B.n198 VSUBS 0.007969f
C316 B.n199 VSUBS 0.007969f
C317 B.n200 VSUBS 0.007969f
C318 B.n201 VSUBS 0.007969f
C319 B.n202 VSUBS 0.007969f
C320 B.n203 VSUBS 0.007969f
C321 B.n204 VSUBS 0.007969f
C322 B.n205 VSUBS 0.007969f
C323 B.n206 VSUBS 0.007969f
C324 B.n207 VSUBS 0.007969f
C325 B.n208 VSUBS 0.007969f
C326 B.n209 VSUBS 0.007969f
C327 B.n210 VSUBS 0.007969f
C328 B.n211 VSUBS 0.007969f
C329 B.n212 VSUBS 0.007969f
C330 B.n213 VSUBS 0.007969f
C331 B.n214 VSUBS 0.007969f
C332 B.n215 VSUBS 0.007969f
C333 B.n216 VSUBS 0.007969f
C334 B.n217 VSUBS 0.007969f
C335 B.n218 VSUBS 0.007969f
C336 B.n219 VSUBS 0.007969f
C337 B.n220 VSUBS 0.007969f
C338 B.n221 VSUBS 0.007969f
C339 B.n222 VSUBS 0.007969f
C340 B.n223 VSUBS 0.017919f
C341 B.n224 VSUBS 0.017919f
C342 B.n225 VSUBS 0.01888f
C343 B.n226 VSUBS 0.007969f
C344 B.n227 VSUBS 0.007969f
C345 B.n228 VSUBS 0.007969f
C346 B.n229 VSUBS 0.007969f
C347 B.n230 VSUBS 0.007969f
C348 B.n231 VSUBS 0.007969f
C349 B.n232 VSUBS 0.007969f
C350 B.n233 VSUBS 0.007969f
C351 B.n234 VSUBS 0.007969f
C352 B.n235 VSUBS 0.007969f
C353 B.n236 VSUBS 0.007969f
C354 B.n237 VSUBS 0.007969f
C355 B.n238 VSUBS 0.007969f
C356 B.n239 VSUBS 0.007969f
C357 B.n240 VSUBS 0.007969f
C358 B.n241 VSUBS 0.007969f
C359 B.n242 VSUBS 0.007969f
C360 B.n243 VSUBS 0.007969f
C361 B.t2 VSUBS 0.047402f
C362 B.t1 VSUBS 0.064327f
C363 B.t0 VSUBS 0.388846f
C364 B.n244 VSUBS 0.112429f
C365 B.n245 VSUBS 0.095605f
C366 B.n246 VSUBS 0.018464f
C367 B.n247 VSUBS 0.0075f
C368 B.n248 VSUBS 0.007969f
C369 B.n249 VSUBS 0.007969f
C370 B.n250 VSUBS 0.007969f
C371 B.n251 VSUBS 0.007969f
C372 B.n252 VSUBS 0.007969f
C373 B.n253 VSUBS 0.007969f
C374 B.n254 VSUBS 0.007969f
C375 B.n255 VSUBS 0.007969f
C376 B.n256 VSUBS 0.007969f
C377 B.n257 VSUBS 0.007969f
C378 B.n258 VSUBS 0.007969f
C379 B.n259 VSUBS 0.007969f
C380 B.n260 VSUBS 0.007969f
C381 B.n261 VSUBS 0.007969f
C382 B.n262 VSUBS 0.007969f
C383 B.n263 VSUBS 0.004453f
C384 B.n264 VSUBS 0.018464f
C385 B.n265 VSUBS 0.0075f
C386 B.n266 VSUBS 0.007969f
C387 B.n267 VSUBS 0.007969f
C388 B.n268 VSUBS 0.007969f
C389 B.n269 VSUBS 0.007969f
C390 B.n270 VSUBS 0.007969f
C391 B.n271 VSUBS 0.007969f
C392 B.n272 VSUBS 0.007969f
C393 B.n273 VSUBS 0.007969f
C394 B.n274 VSUBS 0.007969f
C395 B.n275 VSUBS 0.007969f
C396 B.n276 VSUBS 0.007969f
C397 B.n277 VSUBS 0.007969f
C398 B.n278 VSUBS 0.007969f
C399 B.n279 VSUBS 0.007969f
C400 B.n280 VSUBS 0.007969f
C401 B.n281 VSUBS 0.007969f
C402 B.n282 VSUBS 0.007969f
C403 B.n283 VSUBS 0.007969f
C404 B.n284 VSUBS 0.017919f
C405 B.n285 VSUBS 0.01888f
C406 B.n286 VSUBS 0.017919f
C407 B.n287 VSUBS 0.007969f
C408 B.n288 VSUBS 0.007969f
C409 B.n289 VSUBS 0.007969f
C410 B.n290 VSUBS 0.007969f
C411 B.n291 VSUBS 0.007969f
C412 B.n292 VSUBS 0.007969f
C413 B.n293 VSUBS 0.007969f
C414 B.n294 VSUBS 0.007969f
C415 B.n295 VSUBS 0.007969f
C416 B.n296 VSUBS 0.007969f
C417 B.n297 VSUBS 0.007969f
C418 B.n298 VSUBS 0.007969f
C419 B.n299 VSUBS 0.007969f
C420 B.n300 VSUBS 0.007969f
C421 B.n301 VSUBS 0.007969f
C422 B.n302 VSUBS 0.007969f
C423 B.n303 VSUBS 0.007969f
C424 B.n304 VSUBS 0.007969f
C425 B.n305 VSUBS 0.007969f
C426 B.n306 VSUBS 0.007969f
C427 B.n307 VSUBS 0.007969f
C428 B.n308 VSUBS 0.007969f
C429 B.n309 VSUBS 0.007969f
C430 B.n310 VSUBS 0.007969f
C431 B.n311 VSUBS 0.007969f
C432 B.n312 VSUBS 0.007969f
C433 B.n313 VSUBS 0.007969f
C434 B.n314 VSUBS 0.007969f
C435 B.n315 VSUBS 0.007969f
C436 B.n316 VSUBS 0.007969f
C437 B.n317 VSUBS 0.007969f
C438 B.n318 VSUBS 0.007969f
C439 B.n319 VSUBS 0.007969f
C440 B.n320 VSUBS 0.007969f
C441 B.n321 VSUBS 0.007969f
C442 B.n322 VSUBS 0.007969f
C443 B.n323 VSUBS 0.007969f
C444 B.n324 VSUBS 0.007969f
C445 B.n325 VSUBS 0.007969f
C446 B.n326 VSUBS 0.007969f
C447 B.n327 VSUBS 0.007969f
C448 B.n328 VSUBS 0.007969f
C449 B.n329 VSUBS 0.007969f
C450 B.n330 VSUBS 0.007969f
C451 B.n331 VSUBS 0.007969f
C452 B.n332 VSUBS 0.007969f
C453 B.n333 VSUBS 0.007969f
C454 B.n334 VSUBS 0.007969f
C455 B.n335 VSUBS 0.007969f
C456 B.n336 VSUBS 0.007969f
C457 B.n337 VSUBS 0.007969f
C458 B.n338 VSUBS 0.007969f
C459 B.n339 VSUBS 0.007969f
C460 B.n340 VSUBS 0.007969f
C461 B.n341 VSUBS 0.007969f
C462 B.n342 VSUBS 0.007969f
C463 B.n343 VSUBS 0.007969f
C464 B.n344 VSUBS 0.007969f
C465 B.n345 VSUBS 0.007969f
C466 B.n346 VSUBS 0.007969f
C467 B.n347 VSUBS 0.007969f
C468 B.n348 VSUBS 0.007969f
C469 B.n349 VSUBS 0.007969f
C470 B.n350 VSUBS 0.007969f
C471 B.n351 VSUBS 0.007969f
C472 B.n352 VSUBS 0.007969f
C473 B.n353 VSUBS 0.007969f
C474 B.n354 VSUBS 0.007969f
C475 B.n355 VSUBS 0.007969f
C476 B.n356 VSUBS 0.007969f
C477 B.n357 VSUBS 0.007969f
C478 B.n358 VSUBS 0.007969f
C479 B.n359 VSUBS 0.007969f
C480 B.n360 VSUBS 0.007969f
C481 B.n361 VSUBS 0.007969f
C482 B.n362 VSUBS 0.007969f
C483 B.n363 VSUBS 0.007969f
C484 B.n364 VSUBS 0.007969f
C485 B.n365 VSUBS 0.007969f
C486 B.n366 VSUBS 0.007969f
C487 B.n367 VSUBS 0.007969f
C488 B.n368 VSUBS 0.007969f
C489 B.n369 VSUBS 0.007969f
C490 B.n370 VSUBS 0.007969f
C491 B.n371 VSUBS 0.007969f
C492 B.n372 VSUBS 0.007969f
C493 B.n373 VSUBS 0.007969f
C494 B.n374 VSUBS 0.007969f
C495 B.n375 VSUBS 0.007969f
C496 B.n376 VSUBS 0.007969f
C497 B.n377 VSUBS 0.007969f
C498 B.n378 VSUBS 0.007969f
C499 B.n379 VSUBS 0.007969f
C500 B.n380 VSUBS 0.007969f
C501 B.n381 VSUBS 0.007969f
C502 B.n382 VSUBS 0.007969f
C503 B.n383 VSUBS 0.007969f
C504 B.n384 VSUBS 0.007969f
C505 B.n385 VSUBS 0.007969f
C506 B.n386 VSUBS 0.007969f
C507 B.n387 VSUBS 0.007969f
C508 B.n388 VSUBS 0.007969f
C509 B.n389 VSUBS 0.007969f
C510 B.n390 VSUBS 0.007969f
C511 B.n391 VSUBS 0.007969f
C512 B.n392 VSUBS 0.007969f
C513 B.n393 VSUBS 0.007969f
C514 B.n394 VSUBS 0.007969f
C515 B.n395 VSUBS 0.007969f
C516 B.n396 VSUBS 0.007969f
C517 B.n397 VSUBS 0.007969f
C518 B.n398 VSUBS 0.007969f
C519 B.n399 VSUBS 0.007969f
C520 B.n400 VSUBS 0.007969f
C521 B.n401 VSUBS 0.007969f
C522 B.n402 VSUBS 0.007969f
C523 B.n403 VSUBS 0.007969f
C524 B.n404 VSUBS 0.007969f
C525 B.n405 VSUBS 0.007969f
C526 B.n406 VSUBS 0.007969f
C527 B.n407 VSUBS 0.007969f
C528 B.n408 VSUBS 0.007969f
C529 B.n409 VSUBS 0.007969f
C530 B.n410 VSUBS 0.007969f
C531 B.n411 VSUBS 0.007969f
C532 B.n412 VSUBS 0.007969f
C533 B.n413 VSUBS 0.007969f
C534 B.n414 VSUBS 0.007969f
C535 B.n415 VSUBS 0.007969f
C536 B.n416 VSUBS 0.007969f
C537 B.n417 VSUBS 0.007969f
C538 B.n418 VSUBS 0.007969f
C539 B.n419 VSUBS 0.007969f
C540 B.n420 VSUBS 0.007969f
C541 B.n421 VSUBS 0.007969f
C542 B.n422 VSUBS 0.007969f
C543 B.n423 VSUBS 0.007969f
C544 B.n424 VSUBS 0.007969f
C545 B.n425 VSUBS 0.007969f
C546 B.n426 VSUBS 0.007969f
C547 B.n427 VSUBS 0.007969f
C548 B.n428 VSUBS 0.007969f
C549 B.n429 VSUBS 0.007969f
C550 B.n430 VSUBS 0.007969f
C551 B.n431 VSUBS 0.007969f
C552 B.n432 VSUBS 0.007969f
C553 B.n433 VSUBS 0.007969f
C554 B.n434 VSUBS 0.007969f
C555 B.n435 VSUBS 0.007969f
C556 B.n436 VSUBS 0.007969f
C557 B.n437 VSUBS 0.007969f
C558 B.n438 VSUBS 0.007969f
C559 B.n439 VSUBS 0.007969f
C560 B.n440 VSUBS 0.017919f
C561 B.n441 VSUBS 0.017919f
C562 B.n442 VSUBS 0.01888f
C563 B.n443 VSUBS 0.007969f
C564 B.n444 VSUBS 0.007969f
C565 B.n445 VSUBS 0.007969f
C566 B.n446 VSUBS 0.007969f
C567 B.n447 VSUBS 0.007969f
C568 B.n448 VSUBS 0.007969f
C569 B.n449 VSUBS 0.007969f
C570 B.n450 VSUBS 0.007969f
C571 B.n451 VSUBS 0.007969f
C572 B.n452 VSUBS 0.007969f
C573 B.n453 VSUBS 0.007969f
C574 B.n454 VSUBS 0.007969f
C575 B.n455 VSUBS 0.007969f
C576 B.n456 VSUBS 0.007969f
C577 B.n457 VSUBS 0.007969f
C578 B.n458 VSUBS 0.007969f
C579 B.n459 VSUBS 0.007969f
C580 B.n460 VSUBS 0.007969f
C581 B.n461 VSUBS 0.007969f
C582 B.n462 VSUBS 0.0075f
C583 B.n463 VSUBS 0.018464f
C584 B.n464 VSUBS 0.004453f
C585 B.n465 VSUBS 0.007969f
C586 B.n466 VSUBS 0.007969f
C587 B.n467 VSUBS 0.007969f
C588 B.n468 VSUBS 0.007969f
C589 B.n469 VSUBS 0.007969f
C590 B.n470 VSUBS 0.007969f
C591 B.n471 VSUBS 0.007969f
C592 B.n472 VSUBS 0.007969f
C593 B.n473 VSUBS 0.007969f
C594 B.n474 VSUBS 0.007969f
C595 B.n475 VSUBS 0.007969f
C596 B.n476 VSUBS 0.007969f
C597 B.n477 VSUBS 0.004453f
C598 B.n478 VSUBS 0.007969f
C599 B.n479 VSUBS 0.007969f
C600 B.n480 VSUBS 0.007969f
C601 B.n481 VSUBS 0.007969f
C602 B.n482 VSUBS 0.007969f
C603 B.n483 VSUBS 0.007969f
C604 B.n484 VSUBS 0.007969f
C605 B.n485 VSUBS 0.007969f
C606 B.n486 VSUBS 0.007969f
C607 B.n487 VSUBS 0.007969f
C608 B.n488 VSUBS 0.007969f
C609 B.n489 VSUBS 0.007969f
C610 B.n490 VSUBS 0.007969f
C611 B.n491 VSUBS 0.007969f
C612 B.n492 VSUBS 0.007969f
C613 B.n493 VSUBS 0.007969f
C614 B.n494 VSUBS 0.007969f
C615 B.n495 VSUBS 0.007969f
C616 B.n496 VSUBS 0.007969f
C617 B.n497 VSUBS 0.007969f
C618 B.n498 VSUBS 0.01888f
C619 B.n499 VSUBS 0.01888f
C620 B.n500 VSUBS 0.017919f
C621 B.n501 VSUBS 0.007969f
C622 B.n502 VSUBS 0.007969f
C623 B.n503 VSUBS 0.007969f
C624 B.n504 VSUBS 0.007969f
C625 B.n505 VSUBS 0.007969f
C626 B.n506 VSUBS 0.007969f
C627 B.n507 VSUBS 0.007969f
C628 B.n508 VSUBS 0.007969f
C629 B.n509 VSUBS 0.007969f
C630 B.n510 VSUBS 0.007969f
C631 B.n511 VSUBS 0.007969f
C632 B.n512 VSUBS 0.007969f
C633 B.n513 VSUBS 0.007969f
C634 B.n514 VSUBS 0.007969f
C635 B.n515 VSUBS 0.007969f
C636 B.n516 VSUBS 0.007969f
C637 B.n517 VSUBS 0.007969f
C638 B.n518 VSUBS 0.007969f
C639 B.n519 VSUBS 0.007969f
C640 B.n520 VSUBS 0.007969f
C641 B.n521 VSUBS 0.007969f
C642 B.n522 VSUBS 0.007969f
C643 B.n523 VSUBS 0.007969f
C644 B.n524 VSUBS 0.007969f
C645 B.n525 VSUBS 0.007969f
C646 B.n526 VSUBS 0.007969f
C647 B.n527 VSUBS 0.007969f
C648 B.n528 VSUBS 0.007969f
C649 B.n529 VSUBS 0.007969f
C650 B.n530 VSUBS 0.007969f
C651 B.n531 VSUBS 0.007969f
C652 B.n532 VSUBS 0.007969f
C653 B.n533 VSUBS 0.007969f
C654 B.n534 VSUBS 0.007969f
C655 B.n535 VSUBS 0.007969f
C656 B.n536 VSUBS 0.007969f
C657 B.n537 VSUBS 0.007969f
C658 B.n538 VSUBS 0.007969f
C659 B.n539 VSUBS 0.007969f
C660 B.n540 VSUBS 0.007969f
C661 B.n541 VSUBS 0.007969f
C662 B.n542 VSUBS 0.007969f
C663 B.n543 VSUBS 0.007969f
C664 B.n544 VSUBS 0.007969f
C665 B.n545 VSUBS 0.007969f
C666 B.n546 VSUBS 0.007969f
C667 B.n547 VSUBS 0.007969f
C668 B.n548 VSUBS 0.007969f
C669 B.n549 VSUBS 0.007969f
C670 B.n550 VSUBS 0.007969f
C671 B.n551 VSUBS 0.007969f
C672 B.n552 VSUBS 0.007969f
C673 B.n553 VSUBS 0.007969f
C674 B.n554 VSUBS 0.007969f
C675 B.n555 VSUBS 0.007969f
C676 B.n556 VSUBS 0.007969f
C677 B.n557 VSUBS 0.007969f
C678 B.n558 VSUBS 0.007969f
C679 B.n559 VSUBS 0.007969f
C680 B.n560 VSUBS 0.007969f
C681 B.n561 VSUBS 0.007969f
C682 B.n562 VSUBS 0.007969f
C683 B.n563 VSUBS 0.007969f
C684 B.n564 VSUBS 0.007969f
C685 B.n565 VSUBS 0.007969f
C686 B.n566 VSUBS 0.007969f
C687 B.n567 VSUBS 0.007969f
C688 B.n568 VSUBS 0.007969f
C689 B.n569 VSUBS 0.007969f
C690 B.n570 VSUBS 0.007969f
C691 B.n571 VSUBS 0.007969f
C692 B.n572 VSUBS 0.007969f
C693 B.n573 VSUBS 0.007969f
C694 B.n574 VSUBS 0.007969f
C695 B.n575 VSUBS 0.010399f
C696 B.n576 VSUBS 0.011078f
C697 B.n577 VSUBS 0.022029f
C698 VTAIL.t3 VSUBS 0.069716f
C699 VTAIL.t6 VSUBS 0.069716f
C700 VTAIL.n0 VSUBS 0.283038f
C701 VTAIL.n1 VSUBS 0.696442f
C702 VTAIL.n2 VSUBS 0.037148f
C703 VTAIL.n3 VSUBS 0.268488f
C704 VTAIL.n4 VSUBS 0.017755f
C705 VTAIL.t4 VSUBS 0.098138f
C706 VTAIL.n5 VSUBS 0.118091f
C707 VTAIL.n6 VSUBS 0.029761f
C708 VTAIL.n7 VSUBS 0.031475f
C709 VTAIL.n8 VSUBS 0.104467f
C710 VTAIL.n9 VSUBS 0.0188f
C711 VTAIL.n10 VSUBS 0.017755f
C712 VTAIL.n11 VSUBS 0.072313f
C713 VTAIL.n12 VSUBS 0.052535f
C714 VTAIL.n13 VSUBS 0.346714f
C715 VTAIL.n14 VSUBS 0.037148f
C716 VTAIL.n15 VSUBS 0.268488f
C717 VTAIL.n16 VSUBS 0.017755f
C718 VTAIL.t8 VSUBS 0.098138f
C719 VTAIL.n17 VSUBS 0.118091f
C720 VTAIL.n18 VSUBS 0.029761f
C721 VTAIL.n19 VSUBS 0.031475f
C722 VTAIL.n20 VSUBS 0.104467f
C723 VTAIL.n21 VSUBS 0.0188f
C724 VTAIL.n22 VSUBS 0.017755f
C725 VTAIL.n23 VSUBS 0.072313f
C726 VTAIL.n24 VSUBS 0.052535f
C727 VTAIL.n25 VSUBS 0.346714f
C728 VTAIL.t11 VSUBS 0.069716f
C729 VTAIL.t10 VSUBS 0.069716f
C730 VTAIL.n26 VSUBS 0.283038f
C731 VTAIL.n27 VSUBS 0.961008f
C732 VTAIL.n28 VSUBS 0.037148f
C733 VTAIL.n29 VSUBS 0.268488f
C734 VTAIL.n30 VSUBS 0.017755f
C735 VTAIL.t12 VSUBS 0.098138f
C736 VTAIL.n31 VSUBS 0.118091f
C737 VTAIL.n32 VSUBS 0.029761f
C738 VTAIL.n33 VSUBS 0.031475f
C739 VTAIL.n34 VSUBS 0.104467f
C740 VTAIL.n35 VSUBS 0.0188f
C741 VTAIL.n36 VSUBS 0.017755f
C742 VTAIL.n37 VSUBS 0.072313f
C743 VTAIL.n38 VSUBS 0.052535f
C744 VTAIL.n39 VSUBS 1.26135f
C745 VTAIL.n40 VSUBS 0.037148f
C746 VTAIL.n41 VSUBS 0.268488f
C747 VTAIL.n42 VSUBS 0.017755f
C748 VTAIL.t0 VSUBS 0.098138f
C749 VTAIL.n43 VSUBS 0.118091f
C750 VTAIL.n44 VSUBS 0.029761f
C751 VTAIL.n45 VSUBS 0.031475f
C752 VTAIL.n46 VSUBS 0.104467f
C753 VTAIL.n47 VSUBS 0.0188f
C754 VTAIL.n48 VSUBS 0.017755f
C755 VTAIL.n49 VSUBS 0.072313f
C756 VTAIL.n50 VSUBS 0.052535f
C757 VTAIL.n51 VSUBS 1.26135f
C758 VTAIL.t2 VSUBS 0.069716f
C759 VTAIL.t1 VSUBS 0.069716f
C760 VTAIL.n52 VSUBS 0.28304f
C761 VTAIL.n53 VSUBS 0.961007f
C762 VTAIL.n54 VSUBS 0.037148f
C763 VTAIL.n55 VSUBS 0.268488f
C764 VTAIL.n56 VSUBS 0.017755f
C765 VTAIL.t7 VSUBS 0.098138f
C766 VTAIL.n57 VSUBS 0.118091f
C767 VTAIL.n58 VSUBS 0.029761f
C768 VTAIL.n59 VSUBS 0.031475f
C769 VTAIL.n60 VSUBS 0.104467f
C770 VTAIL.n61 VSUBS 0.0188f
C771 VTAIL.n62 VSUBS 0.017755f
C772 VTAIL.n63 VSUBS 0.072313f
C773 VTAIL.n64 VSUBS 0.052535f
C774 VTAIL.n65 VSUBS 0.346714f
C775 VTAIL.n66 VSUBS 0.037148f
C776 VTAIL.n67 VSUBS 0.268488f
C777 VTAIL.n68 VSUBS 0.017755f
C778 VTAIL.t15 VSUBS 0.098138f
C779 VTAIL.n69 VSUBS 0.118091f
C780 VTAIL.n70 VSUBS 0.029761f
C781 VTAIL.n71 VSUBS 0.031475f
C782 VTAIL.n72 VSUBS 0.104467f
C783 VTAIL.n73 VSUBS 0.0188f
C784 VTAIL.n74 VSUBS 0.017755f
C785 VTAIL.n75 VSUBS 0.072313f
C786 VTAIL.n76 VSUBS 0.052535f
C787 VTAIL.n77 VSUBS 0.346714f
C788 VTAIL.t13 VSUBS 0.069716f
C789 VTAIL.t9 VSUBS 0.069716f
C790 VTAIL.n78 VSUBS 0.28304f
C791 VTAIL.n79 VSUBS 0.961007f
C792 VTAIL.n80 VSUBS 0.037148f
C793 VTAIL.n81 VSUBS 0.268488f
C794 VTAIL.n82 VSUBS 0.017755f
C795 VTAIL.t14 VSUBS 0.098138f
C796 VTAIL.n83 VSUBS 0.118091f
C797 VTAIL.n84 VSUBS 0.029761f
C798 VTAIL.n85 VSUBS 0.031475f
C799 VTAIL.n86 VSUBS 0.104467f
C800 VTAIL.n87 VSUBS 0.0188f
C801 VTAIL.n88 VSUBS 0.017755f
C802 VTAIL.n89 VSUBS 0.072313f
C803 VTAIL.n90 VSUBS 0.052535f
C804 VTAIL.n91 VSUBS 1.26135f
C805 VTAIL.n92 VSUBS 0.037148f
C806 VTAIL.n93 VSUBS 0.268488f
C807 VTAIL.n94 VSUBS 0.017755f
C808 VTAIL.t5 VSUBS 0.098138f
C809 VTAIL.n95 VSUBS 0.118091f
C810 VTAIL.n96 VSUBS 0.029761f
C811 VTAIL.n97 VSUBS 0.031475f
C812 VTAIL.n98 VSUBS 0.104467f
C813 VTAIL.n99 VSUBS 0.0188f
C814 VTAIL.n100 VSUBS 0.017755f
C815 VTAIL.n101 VSUBS 0.072313f
C816 VTAIL.n102 VSUBS 0.052535f
C817 VTAIL.n103 VSUBS 1.25516f
C818 VDD1.t3 VSUBS 0.053114f
C819 VDD1.t4 VSUBS 0.053114f
C820 VDD1.n0 VSUBS 0.259658f
C821 VDD1.t0 VSUBS 0.053114f
C822 VDD1.t1 VSUBS 0.053114f
C823 VDD1.n1 VSUBS 0.259116f
C824 VDD1.t2 VSUBS 0.053114f
C825 VDD1.t6 VSUBS 0.053114f
C826 VDD1.n2 VSUBS 0.259116f
C827 VDD1.n3 VSUBS 3.01756f
C828 VDD1.t5 VSUBS 0.053114f
C829 VDD1.t7 VSUBS 0.053114f
C830 VDD1.n4 VSUBS 0.254088f
C831 VDD1.n5 VSUBS 2.38522f
C832 VP.n0 VSUBS 0.066947f
C833 VP.t7 VSUBS 0.871215f
C834 VP.n1 VSUBS 0.081204f
C835 VP.n2 VSUBS 0.050779f
C836 VP.t5 VSUBS 0.871215f
C837 VP.n3 VSUBS 0.378552f
C838 VP.n4 VSUBS 0.050779f
C839 VP.n5 VSUBS 0.074129f
C840 VP.n6 VSUBS 0.050779f
C841 VP.t4 VSUBS 0.871215f
C842 VP.n7 VSUBS 0.09464f
C843 VP.n8 VSUBS 0.050779f
C844 VP.n9 VSUBS 0.064267f
C845 VP.n10 VSUBS 0.066947f
C846 VP.t1 VSUBS 0.871215f
C847 VP.n11 VSUBS 0.081204f
C848 VP.n12 VSUBS 0.050779f
C849 VP.t6 VSUBS 0.871215f
C850 VP.n13 VSUBS 0.378552f
C851 VP.n14 VSUBS 0.050779f
C852 VP.n15 VSUBS 0.074129f
C853 VP.n16 VSUBS 0.491843f
C854 VP.t2 VSUBS 0.871215f
C855 VP.t0 VSUBS 1.26996f
C856 VP.n17 VSUBS 0.507302f
C857 VP.n18 VSUBS 0.523203f
C858 VP.n19 VSUBS 0.068939f
C859 VP.n20 VSUBS 0.09464f
C860 VP.n21 VSUBS 0.050779f
C861 VP.n22 VSUBS 0.050779f
C862 VP.n23 VSUBS 0.050779f
C863 VP.n24 VSUBS 0.074129f
C864 VP.n25 VSUBS 0.09464f
C865 VP.n26 VSUBS 0.068939f
C866 VP.n27 VSUBS 0.050779f
C867 VP.n28 VSUBS 0.050779f
C868 VP.n29 VSUBS 0.073612f
C869 VP.n30 VSUBS 0.09464f
C870 VP.n31 VSUBS 0.067053f
C871 VP.n32 VSUBS 0.050779f
C872 VP.n33 VSUBS 0.050779f
C873 VP.n34 VSUBS 0.050779f
C874 VP.n35 VSUBS 0.09464f
C875 VP.n36 VSUBS 0.064267f
C876 VP.n37 VSUBS 0.546241f
C877 VP.n38 VSUBS 2.32291f
C878 VP.t3 VSUBS 0.871215f
C879 VP.n39 VSUBS 0.546241f
C880 VP.n40 VSUBS 2.36447f
C881 VP.n41 VSUBS 0.066947f
C882 VP.n42 VSUBS 0.050779f
C883 VP.n43 VSUBS 0.09464f
C884 VP.n44 VSUBS 0.081204f
C885 VP.n45 VSUBS 0.067053f
C886 VP.n46 VSUBS 0.050779f
C887 VP.n47 VSUBS 0.050779f
C888 VP.n48 VSUBS 0.050779f
C889 VP.n49 VSUBS 0.073612f
C890 VP.n50 VSUBS 0.378552f
C891 VP.n51 VSUBS 0.068939f
C892 VP.n52 VSUBS 0.09464f
C893 VP.n53 VSUBS 0.050779f
C894 VP.n54 VSUBS 0.050779f
C895 VP.n55 VSUBS 0.050779f
C896 VP.n56 VSUBS 0.074129f
C897 VP.n57 VSUBS 0.09464f
C898 VP.n58 VSUBS 0.068939f
C899 VP.n59 VSUBS 0.050779f
C900 VP.n60 VSUBS 0.050779f
C901 VP.n61 VSUBS 0.073612f
C902 VP.n62 VSUBS 0.09464f
C903 VP.n63 VSUBS 0.067053f
C904 VP.n64 VSUBS 0.050779f
C905 VP.n65 VSUBS 0.050779f
C906 VP.n66 VSUBS 0.050779f
C907 VP.n67 VSUBS 0.09464f
C908 VP.n68 VSUBS 0.064267f
C909 VP.n69 VSUBS 0.546241f
C910 VP.n70 VSUBS 0.084775f
.ends

