* NGSPICE file created from diff_pair_sample_1299.ext - technology: sky130A

.subckt diff_pair_sample_1299 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=0 ps=0 w=9.04 l=2.55
X1 B.t8 B.t6 B.t7 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=0 ps=0 w=9.04 l=2.55
X2 VDD2.t3 VN.t0 VTAIL.t5 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=1.4916 pd=9.37 as=3.5256 ps=18.86 w=9.04 l=2.55
X3 VDD1.t3 VP.t0 VTAIL.t0 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=1.4916 pd=9.37 as=3.5256 ps=18.86 w=9.04 l=2.55
X4 VDD2.t2 VN.t1 VTAIL.t6 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=1.4916 pd=9.37 as=3.5256 ps=18.86 w=9.04 l=2.55
X5 VTAIL.t4 VN.t2 VDD2.t1 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=1.4916 ps=9.37 w=9.04 l=2.55
X6 VDD1.t2 VP.t1 VTAIL.t1 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=1.4916 pd=9.37 as=3.5256 ps=18.86 w=9.04 l=2.55
X7 VTAIL.t3 VP.t2 VDD1.t1 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=1.4916 ps=9.37 w=9.04 l=2.55
X8 B.t5 B.t3 B.t4 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=0 ps=0 w=9.04 l=2.55
X9 VTAIL.t2 VP.t3 VDD1.t0 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=1.4916 ps=9.37 w=9.04 l=2.55
X10 B.t2 B.t0 B.t1 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=0 ps=0 w=9.04 l=2.55
X11 VTAIL.t7 VN.t3 VDD2.t0 w_n2698_n2776# sky130_fd_pr__pfet_01v8 ad=3.5256 pd=18.86 as=1.4916 ps=9.37 w=9.04 l=2.55
R0 B.n313 B.n94 585
R1 B.n312 B.n311 585
R2 B.n310 B.n95 585
R3 B.n309 B.n308 585
R4 B.n307 B.n96 585
R5 B.n306 B.n305 585
R6 B.n304 B.n97 585
R7 B.n303 B.n302 585
R8 B.n301 B.n98 585
R9 B.n300 B.n299 585
R10 B.n298 B.n99 585
R11 B.n297 B.n296 585
R12 B.n295 B.n100 585
R13 B.n294 B.n293 585
R14 B.n292 B.n101 585
R15 B.n291 B.n290 585
R16 B.n289 B.n102 585
R17 B.n288 B.n287 585
R18 B.n286 B.n103 585
R19 B.n285 B.n284 585
R20 B.n283 B.n104 585
R21 B.n282 B.n281 585
R22 B.n280 B.n105 585
R23 B.n279 B.n278 585
R24 B.n277 B.n106 585
R25 B.n276 B.n275 585
R26 B.n274 B.n107 585
R27 B.n273 B.n272 585
R28 B.n271 B.n108 585
R29 B.n270 B.n269 585
R30 B.n268 B.n109 585
R31 B.n267 B.n266 585
R32 B.n265 B.n110 585
R33 B.n264 B.n263 585
R34 B.n259 B.n111 585
R35 B.n258 B.n257 585
R36 B.n256 B.n112 585
R37 B.n255 B.n254 585
R38 B.n253 B.n113 585
R39 B.n252 B.n251 585
R40 B.n250 B.n114 585
R41 B.n249 B.n248 585
R42 B.n246 B.n115 585
R43 B.n245 B.n244 585
R44 B.n243 B.n118 585
R45 B.n242 B.n241 585
R46 B.n240 B.n119 585
R47 B.n239 B.n238 585
R48 B.n237 B.n120 585
R49 B.n236 B.n235 585
R50 B.n234 B.n121 585
R51 B.n233 B.n232 585
R52 B.n231 B.n122 585
R53 B.n230 B.n229 585
R54 B.n228 B.n123 585
R55 B.n227 B.n226 585
R56 B.n225 B.n124 585
R57 B.n224 B.n223 585
R58 B.n222 B.n125 585
R59 B.n221 B.n220 585
R60 B.n219 B.n126 585
R61 B.n218 B.n217 585
R62 B.n216 B.n127 585
R63 B.n215 B.n214 585
R64 B.n213 B.n128 585
R65 B.n212 B.n211 585
R66 B.n210 B.n129 585
R67 B.n209 B.n208 585
R68 B.n207 B.n130 585
R69 B.n206 B.n205 585
R70 B.n204 B.n131 585
R71 B.n203 B.n202 585
R72 B.n201 B.n132 585
R73 B.n200 B.n199 585
R74 B.n198 B.n133 585
R75 B.n315 B.n314 585
R76 B.n316 B.n93 585
R77 B.n318 B.n317 585
R78 B.n319 B.n92 585
R79 B.n321 B.n320 585
R80 B.n322 B.n91 585
R81 B.n324 B.n323 585
R82 B.n325 B.n90 585
R83 B.n327 B.n326 585
R84 B.n328 B.n89 585
R85 B.n330 B.n329 585
R86 B.n331 B.n88 585
R87 B.n333 B.n332 585
R88 B.n334 B.n87 585
R89 B.n336 B.n335 585
R90 B.n337 B.n86 585
R91 B.n339 B.n338 585
R92 B.n340 B.n85 585
R93 B.n342 B.n341 585
R94 B.n343 B.n84 585
R95 B.n345 B.n344 585
R96 B.n346 B.n83 585
R97 B.n348 B.n347 585
R98 B.n349 B.n82 585
R99 B.n351 B.n350 585
R100 B.n352 B.n81 585
R101 B.n354 B.n353 585
R102 B.n355 B.n80 585
R103 B.n357 B.n356 585
R104 B.n358 B.n79 585
R105 B.n360 B.n359 585
R106 B.n361 B.n78 585
R107 B.n363 B.n362 585
R108 B.n364 B.n77 585
R109 B.n366 B.n365 585
R110 B.n367 B.n76 585
R111 B.n369 B.n368 585
R112 B.n370 B.n75 585
R113 B.n372 B.n371 585
R114 B.n373 B.n74 585
R115 B.n375 B.n374 585
R116 B.n376 B.n73 585
R117 B.n378 B.n377 585
R118 B.n379 B.n72 585
R119 B.n381 B.n380 585
R120 B.n382 B.n71 585
R121 B.n384 B.n383 585
R122 B.n385 B.n70 585
R123 B.n387 B.n386 585
R124 B.n388 B.n69 585
R125 B.n390 B.n389 585
R126 B.n391 B.n68 585
R127 B.n393 B.n392 585
R128 B.n394 B.n67 585
R129 B.n396 B.n395 585
R130 B.n397 B.n66 585
R131 B.n399 B.n398 585
R132 B.n400 B.n65 585
R133 B.n402 B.n401 585
R134 B.n403 B.n64 585
R135 B.n405 B.n404 585
R136 B.n406 B.n63 585
R137 B.n408 B.n407 585
R138 B.n409 B.n62 585
R139 B.n411 B.n410 585
R140 B.n412 B.n61 585
R141 B.n414 B.n413 585
R142 B.n415 B.n60 585
R143 B.n530 B.n529 585
R144 B.n528 B.n19 585
R145 B.n527 B.n526 585
R146 B.n525 B.n20 585
R147 B.n524 B.n523 585
R148 B.n522 B.n21 585
R149 B.n521 B.n520 585
R150 B.n519 B.n22 585
R151 B.n518 B.n517 585
R152 B.n516 B.n23 585
R153 B.n515 B.n514 585
R154 B.n513 B.n24 585
R155 B.n512 B.n511 585
R156 B.n510 B.n25 585
R157 B.n509 B.n508 585
R158 B.n507 B.n26 585
R159 B.n506 B.n505 585
R160 B.n504 B.n27 585
R161 B.n503 B.n502 585
R162 B.n501 B.n28 585
R163 B.n500 B.n499 585
R164 B.n498 B.n29 585
R165 B.n497 B.n496 585
R166 B.n495 B.n30 585
R167 B.n494 B.n493 585
R168 B.n492 B.n31 585
R169 B.n491 B.n490 585
R170 B.n489 B.n32 585
R171 B.n488 B.n487 585
R172 B.n486 B.n33 585
R173 B.n485 B.n484 585
R174 B.n483 B.n34 585
R175 B.n482 B.n481 585
R176 B.n479 B.n35 585
R177 B.n478 B.n477 585
R178 B.n476 B.n38 585
R179 B.n475 B.n474 585
R180 B.n473 B.n39 585
R181 B.n472 B.n471 585
R182 B.n470 B.n40 585
R183 B.n469 B.n468 585
R184 B.n467 B.n41 585
R185 B.n465 B.n464 585
R186 B.n463 B.n44 585
R187 B.n462 B.n461 585
R188 B.n460 B.n45 585
R189 B.n459 B.n458 585
R190 B.n457 B.n46 585
R191 B.n456 B.n455 585
R192 B.n454 B.n47 585
R193 B.n453 B.n452 585
R194 B.n451 B.n48 585
R195 B.n450 B.n449 585
R196 B.n448 B.n49 585
R197 B.n447 B.n446 585
R198 B.n445 B.n50 585
R199 B.n444 B.n443 585
R200 B.n442 B.n51 585
R201 B.n441 B.n440 585
R202 B.n439 B.n52 585
R203 B.n438 B.n437 585
R204 B.n436 B.n53 585
R205 B.n435 B.n434 585
R206 B.n433 B.n54 585
R207 B.n432 B.n431 585
R208 B.n430 B.n55 585
R209 B.n429 B.n428 585
R210 B.n427 B.n56 585
R211 B.n426 B.n425 585
R212 B.n424 B.n57 585
R213 B.n423 B.n422 585
R214 B.n421 B.n58 585
R215 B.n420 B.n419 585
R216 B.n418 B.n59 585
R217 B.n417 B.n416 585
R218 B.n531 B.n18 585
R219 B.n533 B.n532 585
R220 B.n534 B.n17 585
R221 B.n536 B.n535 585
R222 B.n537 B.n16 585
R223 B.n539 B.n538 585
R224 B.n540 B.n15 585
R225 B.n542 B.n541 585
R226 B.n543 B.n14 585
R227 B.n545 B.n544 585
R228 B.n546 B.n13 585
R229 B.n548 B.n547 585
R230 B.n549 B.n12 585
R231 B.n551 B.n550 585
R232 B.n552 B.n11 585
R233 B.n554 B.n553 585
R234 B.n555 B.n10 585
R235 B.n557 B.n556 585
R236 B.n558 B.n9 585
R237 B.n560 B.n559 585
R238 B.n561 B.n8 585
R239 B.n563 B.n562 585
R240 B.n564 B.n7 585
R241 B.n566 B.n565 585
R242 B.n567 B.n6 585
R243 B.n569 B.n568 585
R244 B.n570 B.n5 585
R245 B.n572 B.n571 585
R246 B.n573 B.n4 585
R247 B.n575 B.n574 585
R248 B.n576 B.n3 585
R249 B.n578 B.n577 585
R250 B.n579 B.n0 585
R251 B.n2 B.n1 585
R252 B.n150 B.n149 585
R253 B.n152 B.n151 585
R254 B.n153 B.n148 585
R255 B.n155 B.n154 585
R256 B.n156 B.n147 585
R257 B.n158 B.n157 585
R258 B.n159 B.n146 585
R259 B.n161 B.n160 585
R260 B.n162 B.n145 585
R261 B.n164 B.n163 585
R262 B.n165 B.n144 585
R263 B.n167 B.n166 585
R264 B.n168 B.n143 585
R265 B.n170 B.n169 585
R266 B.n171 B.n142 585
R267 B.n173 B.n172 585
R268 B.n174 B.n141 585
R269 B.n176 B.n175 585
R270 B.n177 B.n140 585
R271 B.n179 B.n178 585
R272 B.n180 B.n139 585
R273 B.n182 B.n181 585
R274 B.n183 B.n138 585
R275 B.n185 B.n184 585
R276 B.n186 B.n137 585
R277 B.n188 B.n187 585
R278 B.n189 B.n136 585
R279 B.n191 B.n190 585
R280 B.n192 B.n135 585
R281 B.n194 B.n193 585
R282 B.n195 B.n134 585
R283 B.n197 B.n196 585
R284 B.n196 B.n133 535.745
R285 B.n314 B.n313 535.745
R286 B.n416 B.n415 535.745
R287 B.n531 B.n530 535.745
R288 B.n116 B.t0 293.408
R289 B.n260 B.t6 293.408
R290 B.n42 B.t3 293.408
R291 B.n36 B.t9 293.408
R292 B.n581 B.n580 256.663
R293 B.n580 B.n579 235.042
R294 B.n580 B.n2 235.042
R295 B.n260 B.t7 167.811
R296 B.n42 B.t5 167.811
R297 B.n116 B.t1 167.802
R298 B.n36 B.t11 167.802
R299 B.n200 B.n133 163.367
R300 B.n201 B.n200 163.367
R301 B.n202 B.n201 163.367
R302 B.n202 B.n131 163.367
R303 B.n206 B.n131 163.367
R304 B.n207 B.n206 163.367
R305 B.n208 B.n207 163.367
R306 B.n208 B.n129 163.367
R307 B.n212 B.n129 163.367
R308 B.n213 B.n212 163.367
R309 B.n214 B.n213 163.367
R310 B.n214 B.n127 163.367
R311 B.n218 B.n127 163.367
R312 B.n219 B.n218 163.367
R313 B.n220 B.n219 163.367
R314 B.n220 B.n125 163.367
R315 B.n224 B.n125 163.367
R316 B.n225 B.n224 163.367
R317 B.n226 B.n225 163.367
R318 B.n226 B.n123 163.367
R319 B.n230 B.n123 163.367
R320 B.n231 B.n230 163.367
R321 B.n232 B.n231 163.367
R322 B.n232 B.n121 163.367
R323 B.n236 B.n121 163.367
R324 B.n237 B.n236 163.367
R325 B.n238 B.n237 163.367
R326 B.n238 B.n119 163.367
R327 B.n242 B.n119 163.367
R328 B.n243 B.n242 163.367
R329 B.n244 B.n243 163.367
R330 B.n244 B.n115 163.367
R331 B.n249 B.n115 163.367
R332 B.n250 B.n249 163.367
R333 B.n251 B.n250 163.367
R334 B.n251 B.n113 163.367
R335 B.n255 B.n113 163.367
R336 B.n256 B.n255 163.367
R337 B.n257 B.n256 163.367
R338 B.n257 B.n111 163.367
R339 B.n264 B.n111 163.367
R340 B.n265 B.n264 163.367
R341 B.n266 B.n265 163.367
R342 B.n266 B.n109 163.367
R343 B.n270 B.n109 163.367
R344 B.n271 B.n270 163.367
R345 B.n272 B.n271 163.367
R346 B.n272 B.n107 163.367
R347 B.n276 B.n107 163.367
R348 B.n277 B.n276 163.367
R349 B.n278 B.n277 163.367
R350 B.n278 B.n105 163.367
R351 B.n282 B.n105 163.367
R352 B.n283 B.n282 163.367
R353 B.n284 B.n283 163.367
R354 B.n284 B.n103 163.367
R355 B.n288 B.n103 163.367
R356 B.n289 B.n288 163.367
R357 B.n290 B.n289 163.367
R358 B.n290 B.n101 163.367
R359 B.n294 B.n101 163.367
R360 B.n295 B.n294 163.367
R361 B.n296 B.n295 163.367
R362 B.n296 B.n99 163.367
R363 B.n300 B.n99 163.367
R364 B.n301 B.n300 163.367
R365 B.n302 B.n301 163.367
R366 B.n302 B.n97 163.367
R367 B.n306 B.n97 163.367
R368 B.n307 B.n306 163.367
R369 B.n308 B.n307 163.367
R370 B.n308 B.n95 163.367
R371 B.n312 B.n95 163.367
R372 B.n313 B.n312 163.367
R373 B.n415 B.n414 163.367
R374 B.n414 B.n61 163.367
R375 B.n410 B.n61 163.367
R376 B.n410 B.n409 163.367
R377 B.n409 B.n408 163.367
R378 B.n408 B.n63 163.367
R379 B.n404 B.n63 163.367
R380 B.n404 B.n403 163.367
R381 B.n403 B.n402 163.367
R382 B.n402 B.n65 163.367
R383 B.n398 B.n65 163.367
R384 B.n398 B.n397 163.367
R385 B.n397 B.n396 163.367
R386 B.n396 B.n67 163.367
R387 B.n392 B.n67 163.367
R388 B.n392 B.n391 163.367
R389 B.n391 B.n390 163.367
R390 B.n390 B.n69 163.367
R391 B.n386 B.n69 163.367
R392 B.n386 B.n385 163.367
R393 B.n385 B.n384 163.367
R394 B.n384 B.n71 163.367
R395 B.n380 B.n71 163.367
R396 B.n380 B.n379 163.367
R397 B.n379 B.n378 163.367
R398 B.n378 B.n73 163.367
R399 B.n374 B.n73 163.367
R400 B.n374 B.n373 163.367
R401 B.n373 B.n372 163.367
R402 B.n372 B.n75 163.367
R403 B.n368 B.n75 163.367
R404 B.n368 B.n367 163.367
R405 B.n367 B.n366 163.367
R406 B.n366 B.n77 163.367
R407 B.n362 B.n77 163.367
R408 B.n362 B.n361 163.367
R409 B.n361 B.n360 163.367
R410 B.n360 B.n79 163.367
R411 B.n356 B.n79 163.367
R412 B.n356 B.n355 163.367
R413 B.n355 B.n354 163.367
R414 B.n354 B.n81 163.367
R415 B.n350 B.n81 163.367
R416 B.n350 B.n349 163.367
R417 B.n349 B.n348 163.367
R418 B.n348 B.n83 163.367
R419 B.n344 B.n83 163.367
R420 B.n344 B.n343 163.367
R421 B.n343 B.n342 163.367
R422 B.n342 B.n85 163.367
R423 B.n338 B.n85 163.367
R424 B.n338 B.n337 163.367
R425 B.n337 B.n336 163.367
R426 B.n336 B.n87 163.367
R427 B.n332 B.n87 163.367
R428 B.n332 B.n331 163.367
R429 B.n331 B.n330 163.367
R430 B.n330 B.n89 163.367
R431 B.n326 B.n89 163.367
R432 B.n326 B.n325 163.367
R433 B.n325 B.n324 163.367
R434 B.n324 B.n91 163.367
R435 B.n320 B.n91 163.367
R436 B.n320 B.n319 163.367
R437 B.n319 B.n318 163.367
R438 B.n318 B.n93 163.367
R439 B.n314 B.n93 163.367
R440 B.n530 B.n19 163.367
R441 B.n526 B.n19 163.367
R442 B.n526 B.n525 163.367
R443 B.n525 B.n524 163.367
R444 B.n524 B.n21 163.367
R445 B.n520 B.n21 163.367
R446 B.n520 B.n519 163.367
R447 B.n519 B.n518 163.367
R448 B.n518 B.n23 163.367
R449 B.n514 B.n23 163.367
R450 B.n514 B.n513 163.367
R451 B.n513 B.n512 163.367
R452 B.n512 B.n25 163.367
R453 B.n508 B.n25 163.367
R454 B.n508 B.n507 163.367
R455 B.n507 B.n506 163.367
R456 B.n506 B.n27 163.367
R457 B.n502 B.n27 163.367
R458 B.n502 B.n501 163.367
R459 B.n501 B.n500 163.367
R460 B.n500 B.n29 163.367
R461 B.n496 B.n29 163.367
R462 B.n496 B.n495 163.367
R463 B.n495 B.n494 163.367
R464 B.n494 B.n31 163.367
R465 B.n490 B.n31 163.367
R466 B.n490 B.n489 163.367
R467 B.n489 B.n488 163.367
R468 B.n488 B.n33 163.367
R469 B.n484 B.n33 163.367
R470 B.n484 B.n483 163.367
R471 B.n483 B.n482 163.367
R472 B.n482 B.n35 163.367
R473 B.n477 B.n35 163.367
R474 B.n477 B.n476 163.367
R475 B.n476 B.n475 163.367
R476 B.n475 B.n39 163.367
R477 B.n471 B.n39 163.367
R478 B.n471 B.n470 163.367
R479 B.n470 B.n469 163.367
R480 B.n469 B.n41 163.367
R481 B.n464 B.n41 163.367
R482 B.n464 B.n463 163.367
R483 B.n463 B.n462 163.367
R484 B.n462 B.n45 163.367
R485 B.n458 B.n45 163.367
R486 B.n458 B.n457 163.367
R487 B.n457 B.n456 163.367
R488 B.n456 B.n47 163.367
R489 B.n452 B.n47 163.367
R490 B.n452 B.n451 163.367
R491 B.n451 B.n450 163.367
R492 B.n450 B.n49 163.367
R493 B.n446 B.n49 163.367
R494 B.n446 B.n445 163.367
R495 B.n445 B.n444 163.367
R496 B.n444 B.n51 163.367
R497 B.n440 B.n51 163.367
R498 B.n440 B.n439 163.367
R499 B.n439 B.n438 163.367
R500 B.n438 B.n53 163.367
R501 B.n434 B.n53 163.367
R502 B.n434 B.n433 163.367
R503 B.n433 B.n432 163.367
R504 B.n432 B.n55 163.367
R505 B.n428 B.n55 163.367
R506 B.n428 B.n427 163.367
R507 B.n427 B.n426 163.367
R508 B.n426 B.n57 163.367
R509 B.n422 B.n57 163.367
R510 B.n422 B.n421 163.367
R511 B.n421 B.n420 163.367
R512 B.n420 B.n59 163.367
R513 B.n416 B.n59 163.367
R514 B.n532 B.n531 163.367
R515 B.n532 B.n17 163.367
R516 B.n536 B.n17 163.367
R517 B.n537 B.n536 163.367
R518 B.n538 B.n537 163.367
R519 B.n538 B.n15 163.367
R520 B.n542 B.n15 163.367
R521 B.n543 B.n542 163.367
R522 B.n544 B.n543 163.367
R523 B.n544 B.n13 163.367
R524 B.n548 B.n13 163.367
R525 B.n549 B.n548 163.367
R526 B.n550 B.n549 163.367
R527 B.n550 B.n11 163.367
R528 B.n554 B.n11 163.367
R529 B.n555 B.n554 163.367
R530 B.n556 B.n555 163.367
R531 B.n556 B.n9 163.367
R532 B.n560 B.n9 163.367
R533 B.n561 B.n560 163.367
R534 B.n562 B.n561 163.367
R535 B.n562 B.n7 163.367
R536 B.n566 B.n7 163.367
R537 B.n567 B.n566 163.367
R538 B.n568 B.n567 163.367
R539 B.n568 B.n5 163.367
R540 B.n572 B.n5 163.367
R541 B.n573 B.n572 163.367
R542 B.n574 B.n573 163.367
R543 B.n574 B.n3 163.367
R544 B.n578 B.n3 163.367
R545 B.n579 B.n578 163.367
R546 B.n149 B.n2 163.367
R547 B.n152 B.n149 163.367
R548 B.n153 B.n152 163.367
R549 B.n154 B.n153 163.367
R550 B.n154 B.n147 163.367
R551 B.n158 B.n147 163.367
R552 B.n159 B.n158 163.367
R553 B.n160 B.n159 163.367
R554 B.n160 B.n145 163.367
R555 B.n164 B.n145 163.367
R556 B.n165 B.n164 163.367
R557 B.n166 B.n165 163.367
R558 B.n166 B.n143 163.367
R559 B.n170 B.n143 163.367
R560 B.n171 B.n170 163.367
R561 B.n172 B.n171 163.367
R562 B.n172 B.n141 163.367
R563 B.n176 B.n141 163.367
R564 B.n177 B.n176 163.367
R565 B.n178 B.n177 163.367
R566 B.n178 B.n139 163.367
R567 B.n182 B.n139 163.367
R568 B.n183 B.n182 163.367
R569 B.n184 B.n183 163.367
R570 B.n184 B.n137 163.367
R571 B.n188 B.n137 163.367
R572 B.n189 B.n188 163.367
R573 B.n190 B.n189 163.367
R574 B.n190 B.n135 163.367
R575 B.n194 B.n135 163.367
R576 B.n195 B.n194 163.367
R577 B.n196 B.n195 163.367
R578 B.n261 B.t8 111.957
R579 B.n43 B.t4 111.957
R580 B.n117 B.t2 111.947
R581 B.n37 B.t10 111.947
R582 B.n247 B.n117 59.5399
R583 B.n262 B.n261 59.5399
R584 B.n466 B.n43 59.5399
R585 B.n480 B.n37 59.5399
R586 B.n117 B.n116 55.855
R587 B.n261 B.n260 55.855
R588 B.n43 B.n42 55.855
R589 B.n37 B.n36 55.855
R590 B.n529 B.n18 34.8103
R591 B.n417 B.n60 34.8103
R592 B.n315 B.n94 34.8103
R593 B.n198 B.n197 34.8103
R594 B B.n581 18.0485
R595 B.n533 B.n18 10.6151
R596 B.n534 B.n533 10.6151
R597 B.n535 B.n534 10.6151
R598 B.n535 B.n16 10.6151
R599 B.n539 B.n16 10.6151
R600 B.n540 B.n539 10.6151
R601 B.n541 B.n540 10.6151
R602 B.n541 B.n14 10.6151
R603 B.n545 B.n14 10.6151
R604 B.n546 B.n545 10.6151
R605 B.n547 B.n546 10.6151
R606 B.n547 B.n12 10.6151
R607 B.n551 B.n12 10.6151
R608 B.n552 B.n551 10.6151
R609 B.n553 B.n552 10.6151
R610 B.n553 B.n10 10.6151
R611 B.n557 B.n10 10.6151
R612 B.n558 B.n557 10.6151
R613 B.n559 B.n558 10.6151
R614 B.n559 B.n8 10.6151
R615 B.n563 B.n8 10.6151
R616 B.n564 B.n563 10.6151
R617 B.n565 B.n564 10.6151
R618 B.n565 B.n6 10.6151
R619 B.n569 B.n6 10.6151
R620 B.n570 B.n569 10.6151
R621 B.n571 B.n570 10.6151
R622 B.n571 B.n4 10.6151
R623 B.n575 B.n4 10.6151
R624 B.n576 B.n575 10.6151
R625 B.n577 B.n576 10.6151
R626 B.n577 B.n0 10.6151
R627 B.n529 B.n528 10.6151
R628 B.n528 B.n527 10.6151
R629 B.n527 B.n20 10.6151
R630 B.n523 B.n20 10.6151
R631 B.n523 B.n522 10.6151
R632 B.n522 B.n521 10.6151
R633 B.n521 B.n22 10.6151
R634 B.n517 B.n22 10.6151
R635 B.n517 B.n516 10.6151
R636 B.n516 B.n515 10.6151
R637 B.n515 B.n24 10.6151
R638 B.n511 B.n24 10.6151
R639 B.n511 B.n510 10.6151
R640 B.n510 B.n509 10.6151
R641 B.n509 B.n26 10.6151
R642 B.n505 B.n26 10.6151
R643 B.n505 B.n504 10.6151
R644 B.n504 B.n503 10.6151
R645 B.n503 B.n28 10.6151
R646 B.n499 B.n28 10.6151
R647 B.n499 B.n498 10.6151
R648 B.n498 B.n497 10.6151
R649 B.n497 B.n30 10.6151
R650 B.n493 B.n30 10.6151
R651 B.n493 B.n492 10.6151
R652 B.n492 B.n491 10.6151
R653 B.n491 B.n32 10.6151
R654 B.n487 B.n32 10.6151
R655 B.n487 B.n486 10.6151
R656 B.n486 B.n485 10.6151
R657 B.n485 B.n34 10.6151
R658 B.n481 B.n34 10.6151
R659 B.n479 B.n478 10.6151
R660 B.n478 B.n38 10.6151
R661 B.n474 B.n38 10.6151
R662 B.n474 B.n473 10.6151
R663 B.n473 B.n472 10.6151
R664 B.n472 B.n40 10.6151
R665 B.n468 B.n40 10.6151
R666 B.n468 B.n467 10.6151
R667 B.n465 B.n44 10.6151
R668 B.n461 B.n44 10.6151
R669 B.n461 B.n460 10.6151
R670 B.n460 B.n459 10.6151
R671 B.n459 B.n46 10.6151
R672 B.n455 B.n46 10.6151
R673 B.n455 B.n454 10.6151
R674 B.n454 B.n453 10.6151
R675 B.n453 B.n48 10.6151
R676 B.n449 B.n48 10.6151
R677 B.n449 B.n448 10.6151
R678 B.n448 B.n447 10.6151
R679 B.n447 B.n50 10.6151
R680 B.n443 B.n50 10.6151
R681 B.n443 B.n442 10.6151
R682 B.n442 B.n441 10.6151
R683 B.n441 B.n52 10.6151
R684 B.n437 B.n52 10.6151
R685 B.n437 B.n436 10.6151
R686 B.n436 B.n435 10.6151
R687 B.n435 B.n54 10.6151
R688 B.n431 B.n54 10.6151
R689 B.n431 B.n430 10.6151
R690 B.n430 B.n429 10.6151
R691 B.n429 B.n56 10.6151
R692 B.n425 B.n56 10.6151
R693 B.n425 B.n424 10.6151
R694 B.n424 B.n423 10.6151
R695 B.n423 B.n58 10.6151
R696 B.n419 B.n58 10.6151
R697 B.n419 B.n418 10.6151
R698 B.n418 B.n417 10.6151
R699 B.n413 B.n60 10.6151
R700 B.n413 B.n412 10.6151
R701 B.n412 B.n411 10.6151
R702 B.n411 B.n62 10.6151
R703 B.n407 B.n62 10.6151
R704 B.n407 B.n406 10.6151
R705 B.n406 B.n405 10.6151
R706 B.n405 B.n64 10.6151
R707 B.n401 B.n64 10.6151
R708 B.n401 B.n400 10.6151
R709 B.n400 B.n399 10.6151
R710 B.n399 B.n66 10.6151
R711 B.n395 B.n66 10.6151
R712 B.n395 B.n394 10.6151
R713 B.n394 B.n393 10.6151
R714 B.n393 B.n68 10.6151
R715 B.n389 B.n68 10.6151
R716 B.n389 B.n388 10.6151
R717 B.n388 B.n387 10.6151
R718 B.n387 B.n70 10.6151
R719 B.n383 B.n70 10.6151
R720 B.n383 B.n382 10.6151
R721 B.n382 B.n381 10.6151
R722 B.n381 B.n72 10.6151
R723 B.n377 B.n72 10.6151
R724 B.n377 B.n376 10.6151
R725 B.n376 B.n375 10.6151
R726 B.n375 B.n74 10.6151
R727 B.n371 B.n74 10.6151
R728 B.n371 B.n370 10.6151
R729 B.n370 B.n369 10.6151
R730 B.n369 B.n76 10.6151
R731 B.n365 B.n76 10.6151
R732 B.n365 B.n364 10.6151
R733 B.n364 B.n363 10.6151
R734 B.n363 B.n78 10.6151
R735 B.n359 B.n78 10.6151
R736 B.n359 B.n358 10.6151
R737 B.n358 B.n357 10.6151
R738 B.n357 B.n80 10.6151
R739 B.n353 B.n80 10.6151
R740 B.n353 B.n352 10.6151
R741 B.n352 B.n351 10.6151
R742 B.n351 B.n82 10.6151
R743 B.n347 B.n82 10.6151
R744 B.n347 B.n346 10.6151
R745 B.n346 B.n345 10.6151
R746 B.n345 B.n84 10.6151
R747 B.n341 B.n84 10.6151
R748 B.n341 B.n340 10.6151
R749 B.n340 B.n339 10.6151
R750 B.n339 B.n86 10.6151
R751 B.n335 B.n86 10.6151
R752 B.n335 B.n334 10.6151
R753 B.n334 B.n333 10.6151
R754 B.n333 B.n88 10.6151
R755 B.n329 B.n88 10.6151
R756 B.n329 B.n328 10.6151
R757 B.n328 B.n327 10.6151
R758 B.n327 B.n90 10.6151
R759 B.n323 B.n90 10.6151
R760 B.n323 B.n322 10.6151
R761 B.n322 B.n321 10.6151
R762 B.n321 B.n92 10.6151
R763 B.n317 B.n92 10.6151
R764 B.n317 B.n316 10.6151
R765 B.n316 B.n315 10.6151
R766 B.n150 B.n1 10.6151
R767 B.n151 B.n150 10.6151
R768 B.n151 B.n148 10.6151
R769 B.n155 B.n148 10.6151
R770 B.n156 B.n155 10.6151
R771 B.n157 B.n156 10.6151
R772 B.n157 B.n146 10.6151
R773 B.n161 B.n146 10.6151
R774 B.n162 B.n161 10.6151
R775 B.n163 B.n162 10.6151
R776 B.n163 B.n144 10.6151
R777 B.n167 B.n144 10.6151
R778 B.n168 B.n167 10.6151
R779 B.n169 B.n168 10.6151
R780 B.n169 B.n142 10.6151
R781 B.n173 B.n142 10.6151
R782 B.n174 B.n173 10.6151
R783 B.n175 B.n174 10.6151
R784 B.n175 B.n140 10.6151
R785 B.n179 B.n140 10.6151
R786 B.n180 B.n179 10.6151
R787 B.n181 B.n180 10.6151
R788 B.n181 B.n138 10.6151
R789 B.n185 B.n138 10.6151
R790 B.n186 B.n185 10.6151
R791 B.n187 B.n186 10.6151
R792 B.n187 B.n136 10.6151
R793 B.n191 B.n136 10.6151
R794 B.n192 B.n191 10.6151
R795 B.n193 B.n192 10.6151
R796 B.n193 B.n134 10.6151
R797 B.n197 B.n134 10.6151
R798 B.n199 B.n198 10.6151
R799 B.n199 B.n132 10.6151
R800 B.n203 B.n132 10.6151
R801 B.n204 B.n203 10.6151
R802 B.n205 B.n204 10.6151
R803 B.n205 B.n130 10.6151
R804 B.n209 B.n130 10.6151
R805 B.n210 B.n209 10.6151
R806 B.n211 B.n210 10.6151
R807 B.n211 B.n128 10.6151
R808 B.n215 B.n128 10.6151
R809 B.n216 B.n215 10.6151
R810 B.n217 B.n216 10.6151
R811 B.n217 B.n126 10.6151
R812 B.n221 B.n126 10.6151
R813 B.n222 B.n221 10.6151
R814 B.n223 B.n222 10.6151
R815 B.n223 B.n124 10.6151
R816 B.n227 B.n124 10.6151
R817 B.n228 B.n227 10.6151
R818 B.n229 B.n228 10.6151
R819 B.n229 B.n122 10.6151
R820 B.n233 B.n122 10.6151
R821 B.n234 B.n233 10.6151
R822 B.n235 B.n234 10.6151
R823 B.n235 B.n120 10.6151
R824 B.n239 B.n120 10.6151
R825 B.n240 B.n239 10.6151
R826 B.n241 B.n240 10.6151
R827 B.n241 B.n118 10.6151
R828 B.n245 B.n118 10.6151
R829 B.n246 B.n245 10.6151
R830 B.n248 B.n114 10.6151
R831 B.n252 B.n114 10.6151
R832 B.n253 B.n252 10.6151
R833 B.n254 B.n253 10.6151
R834 B.n254 B.n112 10.6151
R835 B.n258 B.n112 10.6151
R836 B.n259 B.n258 10.6151
R837 B.n263 B.n259 10.6151
R838 B.n267 B.n110 10.6151
R839 B.n268 B.n267 10.6151
R840 B.n269 B.n268 10.6151
R841 B.n269 B.n108 10.6151
R842 B.n273 B.n108 10.6151
R843 B.n274 B.n273 10.6151
R844 B.n275 B.n274 10.6151
R845 B.n275 B.n106 10.6151
R846 B.n279 B.n106 10.6151
R847 B.n280 B.n279 10.6151
R848 B.n281 B.n280 10.6151
R849 B.n281 B.n104 10.6151
R850 B.n285 B.n104 10.6151
R851 B.n286 B.n285 10.6151
R852 B.n287 B.n286 10.6151
R853 B.n287 B.n102 10.6151
R854 B.n291 B.n102 10.6151
R855 B.n292 B.n291 10.6151
R856 B.n293 B.n292 10.6151
R857 B.n293 B.n100 10.6151
R858 B.n297 B.n100 10.6151
R859 B.n298 B.n297 10.6151
R860 B.n299 B.n298 10.6151
R861 B.n299 B.n98 10.6151
R862 B.n303 B.n98 10.6151
R863 B.n304 B.n303 10.6151
R864 B.n305 B.n304 10.6151
R865 B.n305 B.n96 10.6151
R866 B.n309 B.n96 10.6151
R867 B.n310 B.n309 10.6151
R868 B.n311 B.n310 10.6151
R869 B.n311 B.n94 10.6151
R870 B.n581 B.n0 8.11757
R871 B.n581 B.n1 8.11757
R872 B.n480 B.n479 6.5566
R873 B.n467 B.n466 6.5566
R874 B.n248 B.n247 6.5566
R875 B.n263 B.n262 6.5566
R876 B.n481 B.n480 4.05904
R877 B.n466 B.n465 4.05904
R878 B.n247 B.n246 4.05904
R879 B.n262 B.n110 4.05904
R880 VN.n0 VN.t3 121.337
R881 VN.n1 VN.t1 121.337
R882 VN.n0 VN.t0 120.569
R883 VN.n1 VN.t2 120.569
R884 VN VN.n1 48.594
R885 VN VN.n0 4.41597
R886 VTAIL.n5 VTAIL.t3 69.4255
R887 VTAIL.n4 VTAIL.t6 69.4255
R888 VTAIL.n3 VTAIL.t4 69.4255
R889 VTAIL.n6 VTAIL.t1 69.4252
R890 VTAIL.n7 VTAIL.t5 69.4252
R891 VTAIL.n0 VTAIL.t7 69.4252
R892 VTAIL.n1 VTAIL.t0 69.4252
R893 VTAIL.n2 VTAIL.t2 69.4252
R894 VTAIL.n7 VTAIL.n6 22.6427
R895 VTAIL.n3 VTAIL.n2 22.6427
R896 VTAIL.n4 VTAIL.n3 2.48326
R897 VTAIL.n6 VTAIL.n5 2.48326
R898 VTAIL.n2 VTAIL.n1 2.48326
R899 VTAIL VTAIL.n0 1.30007
R900 VTAIL VTAIL.n7 1.18369
R901 VTAIL.n5 VTAIL.n4 0.470328
R902 VTAIL.n1 VTAIL.n0 0.470328
R903 VDD2.n2 VDD2.n0 121.465
R904 VDD2.n2 VDD2.n1 82.5084
R905 VDD2.n1 VDD2.t1 3.59619
R906 VDD2.n1 VDD2.t2 3.59619
R907 VDD2.n0 VDD2.t0 3.59619
R908 VDD2.n0 VDD2.t3 3.59619
R909 VDD2 VDD2.n2 0.0586897
R910 VP.n14 VP.n0 161.3
R911 VP.n13 VP.n12 161.3
R912 VP.n11 VP.n1 161.3
R913 VP.n10 VP.n9 161.3
R914 VP.n8 VP.n2 161.3
R915 VP.n7 VP.n6 161.3
R916 VP.n4 VP.t2 121.337
R917 VP.n4 VP.t1 120.569
R918 VP.n5 VP.n3 101.564
R919 VP.n16 VP.n15 101.564
R920 VP.n3 VP.t3 85.4374
R921 VP.n15 VP.t0 85.4374
R922 VP.n9 VP.n1 56.5617
R923 VP.n5 VP.n4 48.3152
R924 VP.n8 VP.n7 24.5923
R925 VP.n9 VP.n8 24.5923
R926 VP.n13 VP.n1 24.5923
R927 VP.n14 VP.n13 24.5923
R928 VP.n7 VP.n3 9.3454
R929 VP.n15 VP.n14 9.3454
R930 VP.n6 VP.n5 0.278335
R931 VP.n16 VP.n0 0.278335
R932 VP.n6 VP.n2 0.189894
R933 VP.n10 VP.n2 0.189894
R934 VP.n11 VP.n10 0.189894
R935 VP.n12 VP.n11 0.189894
R936 VP.n12 VP.n0 0.189894
R937 VP VP.n16 0.153485
R938 VDD1 VDD1.n1 121.99
R939 VDD1 VDD1.n0 82.5666
R940 VDD1.n0 VDD1.t1 3.59619
R941 VDD1.n0 VDD1.t2 3.59619
R942 VDD1.n1 VDD1.t0 3.59619
R943 VDD1.n1 VDD1.t3 3.59619
C0 w_n2698_n2776# B 8.35516f
C1 VP VDD1 3.88128f
C2 VP VTAIL 3.6903f
C3 w_n2698_n2776# VDD2 1.42213f
C4 VN VDD1 0.149423f
C5 VN VTAIL 3.6762f
C6 B VDD1 1.17214f
C7 B VTAIL 3.95543f
C8 VP VN 5.60275f
C9 VDD2 VDD1 1.0102f
C10 VDD2 VTAIL 4.74438f
C11 VP B 1.64326f
C12 w_n2698_n2776# VDD1 1.3671f
C13 w_n2698_n2776# VTAIL 3.30846f
C14 VP VDD2 0.391592f
C15 VN B 1.06813f
C16 VP w_n2698_n2776# 4.84435f
C17 VDD2 VN 3.63984f
C18 VTAIL VDD1 4.69051f
C19 w_n2698_n2776# VN 4.49763f
C20 VDD2 B 1.22344f
C21 VDD2 VSUBS 0.871963f
C22 VDD1 VSUBS 5.33768f
C23 VTAIL VSUBS 1.070261f
C24 VN VSUBS 5.35749f
C25 VP VSUBS 2.150437f
C26 B VSUBS 3.984545f
C27 w_n2698_n2776# VSUBS 92.692505f
C28 VDD1.t1 VSUBS 0.196165f
C29 VDD1.t2 VSUBS 0.196165f
C30 VDD1.n0 VSUBS 1.46083f
C31 VDD1.t0 VSUBS 0.196165f
C32 VDD1.t3 VSUBS 0.196165f
C33 VDD1.n1 VSUBS 2.04681f
C34 VP.n0 VSUBS 0.049272f
C35 VP.t0 VSUBS 2.32546f
C36 VP.n1 VSUBS 0.05433f
C37 VP.n2 VSUBS 0.037375f
C38 VP.t3 VSUBS 2.32546f
C39 VP.n3 VSUBS 0.959707f
C40 VP.t1 VSUBS 2.63719f
C41 VP.t2 VSUBS 2.64382f
C42 VP.n4 VSUBS 3.52328f
C43 VP.n5 VSUBS 1.92674f
C44 VP.n6 VSUBS 0.049272f
C45 VP.n7 VSUBS 0.048094f
C46 VP.n8 VSUBS 0.069308f
C47 VP.n9 VSUBS 0.05433f
C48 VP.n10 VSUBS 0.037375f
C49 VP.n11 VSUBS 0.037375f
C50 VP.n12 VSUBS 0.037375f
C51 VP.n13 VSUBS 0.069308f
C52 VP.n14 VSUBS 0.048094f
C53 VP.n15 VSUBS 0.959707f
C54 VP.n16 VSUBS 0.060839f
C55 VDD2.t0 VSUBS 0.191582f
C56 VDD2.t3 VSUBS 0.191582f
C57 VDD2.n0 VSUBS 1.97659f
C58 VDD2.t1 VSUBS 0.191582f
C59 VDD2.t2 VSUBS 0.191582f
C60 VDD2.n1 VSUBS 1.42621f
C61 VDD2.n2 VSUBS 3.91055f
C62 VTAIL.t7 VSUBS 1.62544f
C63 VTAIL.n0 VSUBS 0.728326f
C64 VTAIL.t0 VSUBS 1.62544f
C65 VTAIL.n1 VSUBS 0.823445f
C66 VTAIL.t2 VSUBS 1.62544f
C67 VTAIL.n2 VSUBS 1.95067f
C68 VTAIL.t4 VSUBS 1.62545f
C69 VTAIL.n3 VSUBS 1.95067f
C70 VTAIL.t6 VSUBS 1.62545f
C71 VTAIL.n4 VSUBS 0.82344f
C72 VTAIL.t3 VSUBS 1.62545f
C73 VTAIL.n5 VSUBS 0.82344f
C74 VTAIL.t1 VSUBS 1.62544f
C75 VTAIL.n6 VSUBS 1.95067f
C76 VTAIL.t5 VSUBS 1.62544f
C77 VTAIL.n7 VSUBS 1.8462f
C78 VN.t3 VSUBS 2.54826f
C79 VN.t0 VSUBS 2.54186f
C80 VN.n0 VSUBS 1.61178f
C81 VN.t1 VSUBS 2.54826f
C82 VN.t2 VSUBS 2.54186f
C83 VN.n1 VSUBS 3.41496f
C84 B.n0 VSUBS 0.006501f
C85 B.n1 VSUBS 0.006501f
C86 B.n2 VSUBS 0.009614f
C87 B.n3 VSUBS 0.007367f
C88 B.n4 VSUBS 0.007367f
C89 B.n5 VSUBS 0.007367f
C90 B.n6 VSUBS 0.007367f
C91 B.n7 VSUBS 0.007367f
C92 B.n8 VSUBS 0.007367f
C93 B.n9 VSUBS 0.007367f
C94 B.n10 VSUBS 0.007367f
C95 B.n11 VSUBS 0.007367f
C96 B.n12 VSUBS 0.007367f
C97 B.n13 VSUBS 0.007367f
C98 B.n14 VSUBS 0.007367f
C99 B.n15 VSUBS 0.007367f
C100 B.n16 VSUBS 0.007367f
C101 B.n17 VSUBS 0.007367f
C102 B.n18 VSUBS 0.017716f
C103 B.n19 VSUBS 0.007367f
C104 B.n20 VSUBS 0.007367f
C105 B.n21 VSUBS 0.007367f
C106 B.n22 VSUBS 0.007367f
C107 B.n23 VSUBS 0.007367f
C108 B.n24 VSUBS 0.007367f
C109 B.n25 VSUBS 0.007367f
C110 B.n26 VSUBS 0.007367f
C111 B.n27 VSUBS 0.007367f
C112 B.n28 VSUBS 0.007367f
C113 B.n29 VSUBS 0.007367f
C114 B.n30 VSUBS 0.007367f
C115 B.n31 VSUBS 0.007367f
C116 B.n32 VSUBS 0.007367f
C117 B.n33 VSUBS 0.007367f
C118 B.n34 VSUBS 0.007367f
C119 B.n35 VSUBS 0.007367f
C120 B.t10 VSUBS 0.299224f
C121 B.t11 VSUBS 0.320717f
C122 B.t9 VSUBS 1.12236f
C123 B.n36 VSUBS 0.169909f
C124 B.n37 VSUBS 0.075077f
C125 B.n38 VSUBS 0.007367f
C126 B.n39 VSUBS 0.007367f
C127 B.n40 VSUBS 0.007367f
C128 B.n41 VSUBS 0.007367f
C129 B.t4 VSUBS 0.299221f
C130 B.t5 VSUBS 0.320714f
C131 B.t3 VSUBS 1.12236f
C132 B.n42 VSUBS 0.169912f
C133 B.n43 VSUBS 0.07508f
C134 B.n44 VSUBS 0.007367f
C135 B.n45 VSUBS 0.007367f
C136 B.n46 VSUBS 0.007367f
C137 B.n47 VSUBS 0.007367f
C138 B.n48 VSUBS 0.007367f
C139 B.n49 VSUBS 0.007367f
C140 B.n50 VSUBS 0.007367f
C141 B.n51 VSUBS 0.007367f
C142 B.n52 VSUBS 0.007367f
C143 B.n53 VSUBS 0.007367f
C144 B.n54 VSUBS 0.007367f
C145 B.n55 VSUBS 0.007367f
C146 B.n56 VSUBS 0.007367f
C147 B.n57 VSUBS 0.007367f
C148 B.n58 VSUBS 0.007367f
C149 B.n59 VSUBS 0.007367f
C150 B.n60 VSUBS 0.017716f
C151 B.n61 VSUBS 0.007367f
C152 B.n62 VSUBS 0.007367f
C153 B.n63 VSUBS 0.007367f
C154 B.n64 VSUBS 0.007367f
C155 B.n65 VSUBS 0.007367f
C156 B.n66 VSUBS 0.007367f
C157 B.n67 VSUBS 0.007367f
C158 B.n68 VSUBS 0.007367f
C159 B.n69 VSUBS 0.007367f
C160 B.n70 VSUBS 0.007367f
C161 B.n71 VSUBS 0.007367f
C162 B.n72 VSUBS 0.007367f
C163 B.n73 VSUBS 0.007367f
C164 B.n74 VSUBS 0.007367f
C165 B.n75 VSUBS 0.007367f
C166 B.n76 VSUBS 0.007367f
C167 B.n77 VSUBS 0.007367f
C168 B.n78 VSUBS 0.007367f
C169 B.n79 VSUBS 0.007367f
C170 B.n80 VSUBS 0.007367f
C171 B.n81 VSUBS 0.007367f
C172 B.n82 VSUBS 0.007367f
C173 B.n83 VSUBS 0.007367f
C174 B.n84 VSUBS 0.007367f
C175 B.n85 VSUBS 0.007367f
C176 B.n86 VSUBS 0.007367f
C177 B.n87 VSUBS 0.007367f
C178 B.n88 VSUBS 0.007367f
C179 B.n89 VSUBS 0.007367f
C180 B.n90 VSUBS 0.007367f
C181 B.n91 VSUBS 0.007367f
C182 B.n92 VSUBS 0.007367f
C183 B.n93 VSUBS 0.007367f
C184 B.n94 VSUBS 0.017438f
C185 B.n95 VSUBS 0.007367f
C186 B.n96 VSUBS 0.007367f
C187 B.n97 VSUBS 0.007367f
C188 B.n98 VSUBS 0.007367f
C189 B.n99 VSUBS 0.007367f
C190 B.n100 VSUBS 0.007367f
C191 B.n101 VSUBS 0.007367f
C192 B.n102 VSUBS 0.007367f
C193 B.n103 VSUBS 0.007367f
C194 B.n104 VSUBS 0.007367f
C195 B.n105 VSUBS 0.007367f
C196 B.n106 VSUBS 0.007367f
C197 B.n107 VSUBS 0.007367f
C198 B.n108 VSUBS 0.007367f
C199 B.n109 VSUBS 0.007367f
C200 B.n110 VSUBS 0.005092f
C201 B.n111 VSUBS 0.007367f
C202 B.n112 VSUBS 0.007367f
C203 B.n113 VSUBS 0.007367f
C204 B.n114 VSUBS 0.007367f
C205 B.n115 VSUBS 0.007367f
C206 B.t2 VSUBS 0.299224f
C207 B.t1 VSUBS 0.320717f
C208 B.t0 VSUBS 1.12236f
C209 B.n116 VSUBS 0.169909f
C210 B.n117 VSUBS 0.075077f
C211 B.n118 VSUBS 0.007367f
C212 B.n119 VSUBS 0.007367f
C213 B.n120 VSUBS 0.007367f
C214 B.n121 VSUBS 0.007367f
C215 B.n122 VSUBS 0.007367f
C216 B.n123 VSUBS 0.007367f
C217 B.n124 VSUBS 0.007367f
C218 B.n125 VSUBS 0.007367f
C219 B.n126 VSUBS 0.007367f
C220 B.n127 VSUBS 0.007367f
C221 B.n128 VSUBS 0.007367f
C222 B.n129 VSUBS 0.007367f
C223 B.n130 VSUBS 0.007367f
C224 B.n131 VSUBS 0.007367f
C225 B.n132 VSUBS 0.007367f
C226 B.n133 VSUBS 0.018254f
C227 B.n134 VSUBS 0.007367f
C228 B.n135 VSUBS 0.007367f
C229 B.n136 VSUBS 0.007367f
C230 B.n137 VSUBS 0.007367f
C231 B.n138 VSUBS 0.007367f
C232 B.n139 VSUBS 0.007367f
C233 B.n140 VSUBS 0.007367f
C234 B.n141 VSUBS 0.007367f
C235 B.n142 VSUBS 0.007367f
C236 B.n143 VSUBS 0.007367f
C237 B.n144 VSUBS 0.007367f
C238 B.n145 VSUBS 0.007367f
C239 B.n146 VSUBS 0.007367f
C240 B.n147 VSUBS 0.007367f
C241 B.n148 VSUBS 0.007367f
C242 B.n149 VSUBS 0.007367f
C243 B.n150 VSUBS 0.007367f
C244 B.n151 VSUBS 0.007367f
C245 B.n152 VSUBS 0.007367f
C246 B.n153 VSUBS 0.007367f
C247 B.n154 VSUBS 0.007367f
C248 B.n155 VSUBS 0.007367f
C249 B.n156 VSUBS 0.007367f
C250 B.n157 VSUBS 0.007367f
C251 B.n158 VSUBS 0.007367f
C252 B.n159 VSUBS 0.007367f
C253 B.n160 VSUBS 0.007367f
C254 B.n161 VSUBS 0.007367f
C255 B.n162 VSUBS 0.007367f
C256 B.n163 VSUBS 0.007367f
C257 B.n164 VSUBS 0.007367f
C258 B.n165 VSUBS 0.007367f
C259 B.n166 VSUBS 0.007367f
C260 B.n167 VSUBS 0.007367f
C261 B.n168 VSUBS 0.007367f
C262 B.n169 VSUBS 0.007367f
C263 B.n170 VSUBS 0.007367f
C264 B.n171 VSUBS 0.007367f
C265 B.n172 VSUBS 0.007367f
C266 B.n173 VSUBS 0.007367f
C267 B.n174 VSUBS 0.007367f
C268 B.n175 VSUBS 0.007367f
C269 B.n176 VSUBS 0.007367f
C270 B.n177 VSUBS 0.007367f
C271 B.n178 VSUBS 0.007367f
C272 B.n179 VSUBS 0.007367f
C273 B.n180 VSUBS 0.007367f
C274 B.n181 VSUBS 0.007367f
C275 B.n182 VSUBS 0.007367f
C276 B.n183 VSUBS 0.007367f
C277 B.n184 VSUBS 0.007367f
C278 B.n185 VSUBS 0.007367f
C279 B.n186 VSUBS 0.007367f
C280 B.n187 VSUBS 0.007367f
C281 B.n188 VSUBS 0.007367f
C282 B.n189 VSUBS 0.007367f
C283 B.n190 VSUBS 0.007367f
C284 B.n191 VSUBS 0.007367f
C285 B.n192 VSUBS 0.007367f
C286 B.n193 VSUBS 0.007367f
C287 B.n194 VSUBS 0.007367f
C288 B.n195 VSUBS 0.007367f
C289 B.n196 VSUBS 0.017716f
C290 B.n197 VSUBS 0.017716f
C291 B.n198 VSUBS 0.018254f
C292 B.n199 VSUBS 0.007367f
C293 B.n200 VSUBS 0.007367f
C294 B.n201 VSUBS 0.007367f
C295 B.n202 VSUBS 0.007367f
C296 B.n203 VSUBS 0.007367f
C297 B.n204 VSUBS 0.007367f
C298 B.n205 VSUBS 0.007367f
C299 B.n206 VSUBS 0.007367f
C300 B.n207 VSUBS 0.007367f
C301 B.n208 VSUBS 0.007367f
C302 B.n209 VSUBS 0.007367f
C303 B.n210 VSUBS 0.007367f
C304 B.n211 VSUBS 0.007367f
C305 B.n212 VSUBS 0.007367f
C306 B.n213 VSUBS 0.007367f
C307 B.n214 VSUBS 0.007367f
C308 B.n215 VSUBS 0.007367f
C309 B.n216 VSUBS 0.007367f
C310 B.n217 VSUBS 0.007367f
C311 B.n218 VSUBS 0.007367f
C312 B.n219 VSUBS 0.007367f
C313 B.n220 VSUBS 0.007367f
C314 B.n221 VSUBS 0.007367f
C315 B.n222 VSUBS 0.007367f
C316 B.n223 VSUBS 0.007367f
C317 B.n224 VSUBS 0.007367f
C318 B.n225 VSUBS 0.007367f
C319 B.n226 VSUBS 0.007367f
C320 B.n227 VSUBS 0.007367f
C321 B.n228 VSUBS 0.007367f
C322 B.n229 VSUBS 0.007367f
C323 B.n230 VSUBS 0.007367f
C324 B.n231 VSUBS 0.007367f
C325 B.n232 VSUBS 0.007367f
C326 B.n233 VSUBS 0.007367f
C327 B.n234 VSUBS 0.007367f
C328 B.n235 VSUBS 0.007367f
C329 B.n236 VSUBS 0.007367f
C330 B.n237 VSUBS 0.007367f
C331 B.n238 VSUBS 0.007367f
C332 B.n239 VSUBS 0.007367f
C333 B.n240 VSUBS 0.007367f
C334 B.n241 VSUBS 0.007367f
C335 B.n242 VSUBS 0.007367f
C336 B.n243 VSUBS 0.007367f
C337 B.n244 VSUBS 0.007367f
C338 B.n245 VSUBS 0.007367f
C339 B.n246 VSUBS 0.005092f
C340 B.n247 VSUBS 0.01707f
C341 B.n248 VSUBS 0.005959f
C342 B.n249 VSUBS 0.007367f
C343 B.n250 VSUBS 0.007367f
C344 B.n251 VSUBS 0.007367f
C345 B.n252 VSUBS 0.007367f
C346 B.n253 VSUBS 0.007367f
C347 B.n254 VSUBS 0.007367f
C348 B.n255 VSUBS 0.007367f
C349 B.n256 VSUBS 0.007367f
C350 B.n257 VSUBS 0.007367f
C351 B.n258 VSUBS 0.007367f
C352 B.n259 VSUBS 0.007367f
C353 B.t8 VSUBS 0.299221f
C354 B.t7 VSUBS 0.320714f
C355 B.t6 VSUBS 1.12236f
C356 B.n260 VSUBS 0.169912f
C357 B.n261 VSUBS 0.07508f
C358 B.n262 VSUBS 0.01707f
C359 B.n263 VSUBS 0.005959f
C360 B.n264 VSUBS 0.007367f
C361 B.n265 VSUBS 0.007367f
C362 B.n266 VSUBS 0.007367f
C363 B.n267 VSUBS 0.007367f
C364 B.n268 VSUBS 0.007367f
C365 B.n269 VSUBS 0.007367f
C366 B.n270 VSUBS 0.007367f
C367 B.n271 VSUBS 0.007367f
C368 B.n272 VSUBS 0.007367f
C369 B.n273 VSUBS 0.007367f
C370 B.n274 VSUBS 0.007367f
C371 B.n275 VSUBS 0.007367f
C372 B.n276 VSUBS 0.007367f
C373 B.n277 VSUBS 0.007367f
C374 B.n278 VSUBS 0.007367f
C375 B.n279 VSUBS 0.007367f
C376 B.n280 VSUBS 0.007367f
C377 B.n281 VSUBS 0.007367f
C378 B.n282 VSUBS 0.007367f
C379 B.n283 VSUBS 0.007367f
C380 B.n284 VSUBS 0.007367f
C381 B.n285 VSUBS 0.007367f
C382 B.n286 VSUBS 0.007367f
C383 B.n287 VSUBS 0.007367f
C384 B.n288 VSUBS 0.007367f
C385 B.n289 VSUBS 0.007367f
C386 B.n290 VSUBS 0.007367f
C387 B.n291 VSUBS 0.007367f
C388 B.n292 VSUBS 0.007367f
C389 B.n293 VSUBS 0.007367f
C390 B.n294 VSUBS 0.007367f
C391 B.n295 VSUBS 0.007367f
C392 B.n296 VSUBS 0.007367f
C393 B.n297 VSUBS 0.007367f
C394 B.n298 VSUBS 0.007367f
C395 B.n299 VSUBS 0.007367f
C396 B.n300 VSUBS 0.007367f
C397 B.n301 VSUBS 0.007367f
C398 B.n302 VSUBS 0.007367f
C399 B.n303 VSUBS 0.007367f
C400 B.n304 VSUBS 0.007367f
C401 B.n305 VSUBS 0.007367f
C402 B.n306 VSUBS 0.007367f
C403 B.n307 VSUBS 0.007367f
C404 B.n308 VSUBS 0.007367f
C405 B.n309 VSUBS 0.007367f
C406 B.n310 VSUBS 0.007367f
C407 B.n311 VSUBS 0.007367f
C408 B.n312 VSUBS 0.007367f
C409 B.n313 VSUBS 0.018254f
C410 B.n314 VSUBS 0.017716f
C411 B.n315 VSUBS 0.018533f
C412 B.n316 VSUBS 0.007367f
C413 B.n317 VSUBS 0.007367f
C414 B.n318 VSUBS 0.007367f
C415 B.n319 VSUBS 0.007367f
C416 B.n320 VSUBS 0.007367f
C417 B.n321 VSUBS 0.007367f
C418 B.n322 VSUBS 0.007367f
C419 B.n323 VSUBS 0.007367f
C420 B.n324 VSUBS 0.007367f
C421 B.n325 VSUBS 0.007367f
C422 B.n326 VSUBS 0.007367f
C423 B.n327 VSUBS 0.007367f
C424 B.n328 VSUBS 0.007367f
C425 B.n329 VSUBS 0.007367f
C426 B.n330 VSUBS 0.007367f
C427 B.n331 VSUBS 0.007367f
C428 B.n332 VSUBS 0.007367f
C429 B.n333 VSUBS 0.007367f
C430 B.n334 VSUBS 0.007367f
C431 B.n335 VSUBS 0.007367f
C432 B.n336 VSUBS 0.007367f
C433 B.n337 VSUBS 0.007367f
C434 B.n338 VSUBS 0.007367f
C435 B.n339 VSUBS 0.007367f
C436 B.n340 VSUBS 0.007367f
C437 B.n341 VSUBS 0.007367f
C438 B.n342 VSUBS 0.007367f
C439 B.n343 VSUBS 0.007367f
C440 B.n344 VSUBS 0.007367f
C441 B.n345 VSUBS 0.007367f
C442 B.n346 VSUBS 0.007367f
C443 B.n347 VSUBS 0.007367f
C444 B.n348 VSUBS 0.007367f
C445 B.n349 VSUBS 0.007367f
C446 B.n350 VSUBS 0.007367f
C447 B.n351 VSUBS 0.007367f
C448 B.n352 VSUBS 0.007367f
C449 B.n353 VSUBS 0.007367f
C450 B.n354 VSUBS 0.007367f
C451 B.n355 VSUBS 0.007367f
C452 B.n356 VSUBS 0.007367f
C453 B.n357 VSUBS 0.007367f
C454 B.n358 VSUBS 0.007367f
C455 B.n359 VSUBS 0.007367f
C456 B.n360 VSUBS 0.007367f
C457 B.n361 VSUBS 0.007367f
C458 B.n362 VSUBS 0.007367f
C459 B.n363 VSUBS 0.007367f
C460 B.n364 VSUBS 0.007367f
C461 B.n365 VSUBS 0.007367f
C462 B.n366 VSUBS 0.007367f
C463 B.n367 VSUBS 0.007367f
C464 B.n368 VSUBS 0.007367f
C465 B.n369 VSUBS 0.007367f
C466 B.n370 VSUBS 0.007367f
C467 B.n371 VSUBS 0.007367f
C468 B.n372 VSUBS 0.007367f
C469 B.n373 VSUBS 0.007367f
C470 B.n374 VSUBS 0.007367f
C471 B.n375 VSUBS 0.007367f
C472 B.n376 VSUBS 0.007367f
C473 B.n377 VSUBS 0.007367f
C474 B.n378 VSUBS 0.007367f
C475 B.n379 VSUBS 0.007367f
C476 B.n380 VSUBS 0.007367f
C477 B.n381 VSUBS 0.007367f
C478 B.n382 VSUBS 0.007367f
C479 B.n383 VSUBS 0.007367f
C480 B.n384 VSUBS 0.007367f
C481 B.n385 VSUBS 0.007367f
C482 B.n386 VSUBS 0.007367f
C483 B.n387 VSUBS 0.007367f
C484 B.n388 VSUBS 0.007367f
C485 B.n389 VSUBS 0.007367f
C486 B.n390 VSUBS 0.007367f
C487 B.n391 VSUBS 0.007367f
C488 B.n392 VSUBS 0.007367f
C489 B.n393 VSUBS 0.007367f
C490 B.n394 VSUBS 0.007367f
C491 B.n395 VSUBS 0.007367f
C492 B.n396 VSUBS 0.007367f
C493 B.n397 VSUBS 0.007367f
C494 B.n398 VSUBS 0.007367f
C495 B.n399 VSUBS 0.007367f
C496 B.n400 VSUBS 0.007367f
C497 B.n401 VSUBS 0.007367f
C498 B.n402 VSUBS 0.007367f
C499 B.n403 VSUBS 0.007367f
C500 B.n404 VSUBS 0.007367f
C501 B.n405 VSUBS 0.007367f
C502 B.n406 VSUBS 0.007367f
C503 B.n407 VSUBS 0.007367f
C504 B.n408 VSUBS 0.007367f
C505 B.n409 VSUBS 0.007367f
C506 B.n410 VSUBS 0.007367f
C507 B.n411 VSUBS 0.007367f
C508 B.n412 VSUBS 0.007367f
C509 B.n413 VSUBS 0.007367f
C510 B.n414 VSUBS 0.007367f
C511 B.n415 VSUBS 0.017716f
C512 B.n416 VSUBS 0.018254f
C513 B.n417 VSUBS 0.018254f
C514 B.n418 VSUBS 0.007367f
C515 B.n419 VSUBS 0.007367f
C516 B.n420 VSUBS 0.007367f
C517 B.n421 VSUBS 0.007367f
C518 B.n422 VSUBS 0.007367f
C519 B.n423 VSUBS 0.007367f
C520 B.n424 VSUBS 0.007367f
C521 B.n425 VSUBS 0.007367f
C522 B.n426 VSUBS 0.007367f
C523 B.n427 VSUBS 0.007367f
C524 B.n428 VSUBS 0.007367f
C525 B.n429 VSUBS 0.007367f
C526 B.n430 VSUBS 0.007367f
C527 B.n431 VSUBS 0.007367f
C528 B.n432 VSUBS 0.007367f
C529 B.n433 VSUBS 0.007367f
C530 B.n434 VSUBS 0.007367f
C531 B.n435 VSUBS 0.007367f
C532 B.n436 VSUBS 0.007367f
C533 B.n437 VSUBS 0.007367f
C534 B.n438 VSUBS 0.007367f
C535 B.n439 VSUBS 0.007367f
C536 B.n440 VSUBS 0.007367f
C537 B.n441 VSUBS 0.007367f
C538 B.n442 VSUBS 0.007367f
C539 B.n443 VSUBS 0.007367f
C540 B.n444 VSUBS 0.007367f
C541 B.n445 VSUBS 0.007367f
C542 B.n446 VSUBS 0.007367f
C543 B.n447 VSUBS 0.007367f
C544 B.n448 VSUBS 0.007367f
C545 B.n449 VSUBS 0.007367f
C546 B.n450 VSUBS 0.007367f
C547 B.n451 VSUBS 0.007367f
C548 B.n452 VSUBS 0.007367f
C549 B.n453 VSUBS 0.007367f
C550 B.n454 VSUBS 0.007367f
C551 B.n455 VSUBS 0.007367f
C552 B.n456 VSUBS 0.007367f
C553 B.n457 VSUBS 0.007367f
C554 B.n458 VSUBS 0.007367f
C555 B.n459 VSUBS 0.007367f
C556 B.n460 VSUBS 0.007367f
C557 B.n461 VSUBS 0.007367f
C558 B.n462 VSUBS 0.007367f
C559 B.n463 VSUBS 0.007367f
C560 B.n464 VSUBS 0.007367f
C561 B.n465 VSUBS 0.005092f
C562 B.n466 VSUBS 0.01707f
C563 B.n467 VSUBS 0.005959f
C564 B.n468 VSUBS 0.007367f
C565 B.n469 VSUBS 0.007367f
C566 B.n470 VSUBS 0.007367f
C567 B.n471 VSUBS 0.007367f
C568 B.n472 VSUBS 0.007367f
C569 B.n473 VSUBS 0.007367f
C570 B.n474 VSUBS 0.007367f
C571 B.n475 VSUBS 0.007367f
C572 B.n476 VSUBS 0.007367f
C573 B.n477 VSUBS 0.007367f
C574 B.n478 VSUBS 0.007367f
C575 B.n479 VSUBS 0.005959f
C576 B.n480 VSUBS 0.01707f
C577 B.n481 VSUBS 0.005092f
C578 B.n482 VSUBS 0.007367f
C579 B.n483 VSUBS 0.007367f
C580 B.n484 VSUBS 0.007367f
C581 B.n485 VSUBS 0.007367f
C582 B.n486 VSUBS 0.007367f
C583 B.n487 VSUBS 0.007367f
C584 B.n488 VSUBS 0.007367f
C585 B.n489 VSUBS 0.007367f
C586 B.n490 VSUBS 0.007367f
C587 B.n491 VSUBS 0.007367f
C588 B.n492 VSUBS 0.007367f
C589 B.n493 VSUBS 0.007367f
C590 B.n494 VSUBS 0.007367f
C591 B.n495 VSUBS 0.007367f
C592 B.n496 VSUBS 0.007367f
C593 B.n497 VSUBS 0.007367f
C594 B.n498 VSUBS 0.007367f
C595 B.n499 VSUBS 0.007367f
C596 B.n500 VSUBS 0.007367f
C597 B.n501 VSUBS 0.007367f
C598 B.n502 VSUBS 0.007367f
C599 B.n503 VSUBS 0.007367f
C600 B.n504 VSUBS 0.007367f
C601 B.n505 VSUBS 0.007367f
C602 B.n506 VSUBS 0.007367f
C603 B.n507 VSUBS 0.007367f
C604 B.n508 VSUBS 0.007367f
C605 B.n509 VSUBS 0.007367f
C606 B.n510 VSUBS 0.007367f
C607 B.n511 VSUBS 0.007367f
C608 B.n512 VSUBS 0.007367f
C609 B.n513 VSUBS 0.007367f
C610 B.n514 VSUBS 0.007367f
C611 B.n515 VSUBS 0.007367f
C612 B.n516 VSUBS 0.007367f
C613 B.n517 VSUBS 0.007367f
C614 B.n518 VSUBS 0.007367f
C615 B.n519 VSUBS 0.007367f
C616 B.n520 VSUBS 0.007367f
C617 B.n521 VSUBS 0.007367f
C618 B.n522 VSUBS 0.007367f
C619 B.n523 VSUBS 0.007367f
C620 B.n524 VSUBS 0.007367f
C621 B.n525 VSUBS 0.007367f
C622 B.n526 VSUBS 0.007367f
C623 B.n527 VSUBS 0.007367f
C624 B.n528 VSUBS 0.007367f
C625 B.n529 VSUBS 0.018254f
C626 B.n530 VSUBS 0.018254f
C627 B.n531 VSUBS 0.017716f
C628 B.n532 VSUBS 0.007367f
C629 B.n533 VSUBS 0.007367f
C630 B.n534 VSUBS 0.007367f
C631 B.n535 VSUBS 0.007367f
C632 B.n536 VSUBS 0.007367f
C633 B.n537 VSUBS 0.007367f
C634 B.n538 VSUBS 0.007367f
C635 B.n539 VSUBS 0.007367f
C636 B.n540 VSUBS 0.007367f
C637 B.n541 VSUBS 0.007367f
C638 B.n542 VSUBS 0.007367f
C639 B.n543 VSUBS 0.007367f
C640 B.n544 VSUBS 0.007367f
C641 B.n545 VSUBS 0.007367f
C642 B.n546 VSUBS 0.007367f
C643 B.n547 VSUBS 0.007367f
C644 B.n548 VSUBS 0.007367f
C645 B.n549 VSUBS 0.007367f
C646 B.n550 VSUBS 0.007367f
C647 B.n551 VSUBS 0.007367f
C648 B.n552 VSUBS 0.007367f
C649 B.n553 VSUBS 0.007367f
C650 B.n554 VSUBS 0.007367f
C651 B.n555 VSUBS 0.007367f
C652 B.n556 VSUBS 0.007367f
C653 B.n557 VSUBS 0.007367f
C654 B.n558 VSUBS 0.007367f
C655 B.n559 VSUBS 0.007367f
C656 B.n560 VSUBS 0.007367f
C657 B.n561 VSUBS 0.007367f
C658 B.n562 VSUBS 0.007367f
C659 B.n563 VSUBS 0.007367f
C660 B.n564 VSUBS 0.007367f
C661 B.n565 VSUBS 0.007367f
C662 B.n566 VSUBS 0.007367f
C663 B.n567 VSUBS 0.007367f
C664 B.n568 VSUBS 0.007367f
C665 B.n569 VSUBS 0.007367f
C666 B.n570 VSUBS 0.007367f
C667 B.n571 VSUBS 0.007367f
C668 B.n572 VSUBS 0.007367f
C669 B.n573 VSUBS 0.007367f
C670 B.n574 VSUBS 0.007367f
C671 B.n575 VSUBS 0.007367f
C672 B.n576 VSUBS 0.007367f
C673 B.n577 VSUBS 0.007367f
C674 B.n578 VSUBS 0.007367f
C675 B.n579 VSUBS 0.009614f
C676 B.n580 VSUBS 0.010242f
C677 B.n581 VSUBS 0.020366f
.ends

