* NGSPICE file created from diff_pair_sample_1779.ext - technology: sky130A

.subckt diff_pair_sample_1779 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0.9042 ps=5.81 w=5.48 l=1.21
X1 VDD1.t4 VP.t1 VTAIL.t10 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=2.1372 ps=11.74 w=5.48 l=1.21
X2 VDD2.t5 VN.t0 VTAIL.t3 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=2.1372 ps=11.74 w=5.48 l=1.21
X3 VDD1.t3 VP.t2 VTAIL.t11 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=2.1372 ps=11.74 w=5.48 l=1.21
X4 B.t11 B.t9 B.t10 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0 ps=0 w=5.48 l=1.21
X5 VTAIL.t7 VP.t3 VDD1.t2 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=0.9042 ps=5.81 w=5.48 l=1.21
X6 VDD2.t4 VN.t1 VTAIL.t5 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=2.1372 ps=11.74 w=5.48 l=1.21
X7 VDD2.t3 VN.t2 VTAIL.t0 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0.9042 ps=5.81 w=5.48 l=1.21
X8 B.t8 B.t6 B.t7 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0 ps=0 w=5.48 l=1.21
X9 VTAIL.t9 VP.t4 VDD1.t1 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=0.9042 ps=5.81 w=5.48 l=1.21
X10 B.t5 B.t3 B.t4 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0 ps=0 w=5.48 l=1.21
X11 B.t2 B.t0 B.t1 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0 ps=0 w=5.48 l=1.21
X12 VDD1.t0 VP.t5 VTAIL.t8 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0.9042 ps=5.81 w=5.48 l=1.21
X13 VDD2.t2 VN.t3 VTAIL.t1 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=2.1372 pd=11.74 as=0.9042 ps=5.81 w=5.48 l=1.21
X14 VTAIL.t2 VN.t4 VDD2.t1 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=0.9042 ps=5.81 w=5.48 l=1.21
X15 VTAIL.t4 VN.t5 VDD2.t0 w_n2202_n2064# sky130_fd_pr__pfet_01v8 ad=0.9042 pd=5.81 as=0.9042 ps=5.81 w=5.48 l=1.21
R0 VP.n14 VP.n3 171.63
R1 VP.n26 VP.n25 171.63
R2 VP.n13 VP.n12 171.63
R3 VP.n8 VP.n5 161.3
R4 VP.n10 VP.n9 161.3
R5 VP.n11 VP.n4 161.3
R6 VP.n24 VP.n0 161.3
R7 VP.n23 VP.n22 161.3
R8 VP.n21 VP.n1 161.3
R9 VP.n20 VP.n19 161.3
R10 VP.n17 VP.n2 161.3
R11 VP.n16 VP.n15 161.3
R12 VP.n7 VP.t0 140.554
R13 VP.n3 VP.t5 109.147
R14 VP.n18 VP.t3 109.147
R15 VP.n25 VP.t2 109.147
R16 VP.n12 VP.t1 109.147
R17 VP.n6 VP.t4 109.147
R18 VP.n7 VP.n6 51.4185
R19 VP.n17 VP.n16 42.5146
R20 VP.n24 VP.n23 42.5146
R21 VP.n11 VP.n10 42.5146
R22 VP.n19 VP.n17 38.6395
R23 VP.n23 VP.n1 38.6395
R24 VP.n10 VP.n5 38.6395
R25 VP.n14 VP.n13 38.205
R26 VP.n8 VP.n7 26.6589
R27 VP.n16 VP.n3 14.2638
R28 VP.n25 VP.n24 14.2638
R29 VP.n12 VP.n11 14.2638
R30 VP.n19 VP.n18 12.2964
R31 VP.n18 VP.n1 12.2964
R32 VP.n6 VP.n5 12.2964
R33 VP.n9 VP.n8 0.189894
R34 VP.n9 VP.n4 0.189894
R35 VP.n13 VP.n4 0.189894
R36 VP.n15 VP.n14 0.189894
R37 VP.n15 VP.n2 0.189894
R38 VP.n20 VP.n2 0.189894
R39 VP.n21 VP.n20 0.189894
R40 VP.n22 VP.n21 0.189894
R41 VP.n22 VP.n0 0.189894
R42 VP.n26 VP.n0 0.189894
R43 VP VP.n26 0.0516364
R44 VTAIL.n7 VTAIL.t5 87.0253
R45 VTAIL.n10 VTAIL.t10 87.0243
R46 VTAIL.n11 VTAIL.t3 87.0243
R47 VTAIL.n2 VTAIL.t11 87.0243
R48 VTAIL.n9 VTAIL.n8 81.0937
R49 VTAIL.n6 VTAIL.n5 81.0937
R50 VTAIL.n1 VTAIL.n0 81.0936
R51 VTAIL.n4 VTAIL.n3 81.0936
R52 VTAIL.n6 VTAIL.n4 19.7462
R53 VTAIL.n11 VTAIL.n10 18.4186
R54 VTAIL.n0 VTAIL.t1 5.93207
R55 VTAIL.n0 VTAIL.t2 5.93207
R56 VTAIL.n3 VTAIL.t8 5.93207
R57 VTAIL.n3 VTAIL.t7 5.93207
R58 VTAIL.n8 VTAIL.t6 5.93207
R59 VTAIL.n8 VTAIL.t9 5.93207
R60 VTAIL.n5 VTAIL.t0 5.93207
R61 VTAIL.n5 VTAIL.t4 5.93207
R62 VTAIL.n7 VTAIL.n6 1.32809
R63 VTAIL.n10 VTAIL.n9 1.32809
R64 VTAIL.n4 VTAIL.n2 1.32809
R65 VTAIL.n9 VTAIL.n7 1.13412
R66 VTAIL.n2 VTAIL.n1 1.13412
R67 VTAIL VTAIL.n11 0.938
R68 VTAIL VTAIL.n1 0.390586
R69 VDD1 VDD1.t5 104.757
R70 VDD1.n1 VDD1.t0 104.644
R71 VDD1.n1 VDD1.n0 98.0489
R72 VDD1.n3 VDD1.n2 97.7715
R73 VDD1.n3 VDD1.n1 34.0009
R74 VDD1.n2 VDD1.t1 5.93207
R75 VDD1.n2 VDD1.t4 5.93207
R76 VDD1.n0 VDD1.t2 5.93207
R77 VDD1.n0 VDD1.t3 5.93207
R78 VDD1 VDD1.n3 0.274207
R79 VN.n9 VN.n8 171.63
R80 VN.n19 VN.n18 171.63
R81 VN.n17 VN.n10 161.3
R82 VN.n16 VN.n15 161.3
R83 VN.n14 VN.n11 161.3
R84 VN.n7 VN.n0 161.3
R85 VN.n6 VN.n5 161.3
R86 VN.n4 VN.n1 161.3
R87 VN.n3 VN.t3 140.554
R88 VN.n13 VN.t1 140.554
R89 VN.n2 VN.t4 109.147
R90 VN.n8 VN.t0 109.147
R91 VN.n12 VN.t5 109.147
R92 VN.n18 VN.t2 109.147
R93 VN.n3 VN.n2 51.4185
R94 VN.n13 VN.n12 51.4185
R95 VN.n7 VN.n6 42.5146
R96 VN.n17 VN.n16 42.5146
R97 VN.n6 VN.n1 38.6395
R98 VN.n16 VN.n11 38.6395
R99 VN VN.n19 38.5857
R100 VN.n14 VN.n13 26.6589
R101 VN.n4 VN.n3 26.6589
R102 VN.n8 VN.n7 14.2638
R103 VN.n18 VN.n17 14.2638
R104 VN.n2 VN.n1 12.2964
R105 VN.n12 VN.n11 12.2964
R106 VN.n19 VN.n10 0.189894
R107 VN.n15 VN.n10 0.189894
R108 VN.n15 VN.n14 0.189894
R109 VN.n5 VN.n4 0.189894
R110 VN.n5 VN.n0 0.189894
R111 VN.n9 VN.n0 0.189894
R112 VN VN.n9 0.0516364
R113 VDD2.n1 VDD2.t2 104.644
R114 VDD2.n2 VDD2.t3 103.704
R115 VDD2.n1 VDD2.n0 98.0489
R116 VDD2 VDD2.n3 98.0452
R117 VDD2.n2 VDD2.n1 32.7541
R118 VDD2.n3 VDD2.t0 5.93207
R119 VDD2.n3 VDD2.t4 5.93207
R120 VDD2.n0 VDD2.t1 5.93207
R121 VDD2.n0 VDD2.t5 5.93207
R122 VDD2 VDD2.n2 1.05438
R123 B.n317 B.n46 585
R124 B.n319 B.n318 585
R125 B.n320 B.n45 585
R126 B.n322 B.n321 585
R127 B.n323 B.n44 585
R128 B.n325 B.n324 585
R129 B.n326 B.n43 585
R130 B.n328 B.n327 585
R131 B.n329 B.n42 585
R132 B.n331 B.n330 585
R133 B.n332 B.n41 585
R134 B.n334 B.n333 585
R135 B.n335 B.n40 585
R136 B.n337 B.n336 585
R137 B.n338 B.n39 585
R138 B.n340 B.n339 585
R139 B.n341 B.n38 585
R140 B.n343 B.n342 585
R141 B.n344 B.n37 585
R142 B.n346 B.n345 585
R143 B.n347 B.n36 585
R144 B.n349 B.n348 585
R145 B.n351 B.n33 585
R146 B.n353 B.n352 585
R147 B.n354 B.n32 585
R148 B.n356 B.n355 585
R149 B.n357 B.n31 585
R150 B.n359 B.n358 585
R151 B.n360 B.n30 585
R152 B.n362 B.n361 585
R153 B.n363 B.n29 585
R154 B.n365 B.n364 585
R155 B.n367 B.n366 585
R156 B.n368 B.n25 585
R157 B.n370 B.n369 585
R158 B.n371 B.n24 585
R159 B.n373 B.n372 585
R160 B.n374 B.n23 585
R161 B.n376 B.n375 585
R162 B.n377 B.n22 585
R163 B.n379 B.n378 585
R164 B.n380 B.n21 585
R165 B.n382 B.n381 585
R166 B.n383 B.n20 585
R167 B.n385 B.n384 585
R168 B.n386 B.n19 585
R169 B.n388 B.n387 585
R170 B.n389 B.n18 585
R171 B.n391 B.n390 585
R172 B.n392 B.n17 585
R173 B.n394 B.n393 585
R174 B.n395 B.n16 585
R175 B.n397 B.n396 585
R176 B.n398 B.n15 585
R177 B.n316 B.n315 585
R178 B.n314 B.n47 585
R179 B.n313 B.n312 585
R180 B.n311 B.n48 585
R181 B.n310 B.n309 585
R182 B.n308 B.n49 585
R183 B.n307 B.n306 585
R184 B.n305 B.n50 585
R185 B.n304 B.n303 585
R186 B.n302 B.n51 585
R187 B.n301 B.n300 585
R188 B.n299 B.n52 585
R189 B.n298 B.n297 585
R190 B.n296 B.n53 585
R191 B.n295 B.n294 585
R192 B.n293 B.n54 585
R193 B.n292 B.n291 585
R194 B.n290 B.n55 585
R195 B.n289 B.n288 585
R196 B.n287 B.n56 585
R197 B.n286 B.n285 585
R198 B.n284 B.n57 585
R199 B.n283 B.n282 585
R200 B.n281 B.n58 585
R201 B.n280 B.n279 585
R202 B.n278 B.n59 585
R203 B.n277 B.n276 585
R204 B.n275 B.n60 585
R205 B.n274 B.n273 585
R206 B.n272 B.n61 585
R207 B.n271 B.n270 585
R208 B.n269 B.n62 585
R209 B.n268 B.n267 585
R210 B.n266 B.n63 585
R211 B.n265 B.n264 585
R212 B.n263 B.n64 585
R213 B.n262 B.n261 585
R214 B.n260 B.n65 585
R215 B.n259 B.n258 585
R216 B.n257 B.n66 585
R217 B.n256 B.n255 585
R218 B.n254 B.n67 585
R219 B.n253 B.n252 585
R220 B.n251 B.n68 585
R221 B.n250 B.n249 585
R222 B.n248 B.n69 585
R223 B.n247 B.n246 585
R224 B.n245 B.n70 585
R225 B.n244 B.n243 585
R226 B.n242 B.n71 585
R227 B.n241 B.n240 585
R228 B.n239 B.n72 585
R229 B.n238 B.n237 585
R230 B.n155 B.n104 585
R231 B.n157 B.n156 585
R232 B.n158 B.n103 585
R233 B.n160 B.n159 585
R234 B.n161 B.n102 585
R235 B.n163 B.n162 585
R236 B.n164 B.n101 585
R237 B.n166 B.n165 585
R238 B.n167 B.n100 585
R239 B.n169 B.n168 585
R240 B.n170 B.n99 585
R241 B.n172 B.n171 585
R242 B.n173 B.n98 585
R243 B.n175 B.n174 585
R244 B.n176 B.n97 585
R245 B.n178 B.n177 585
R246 B.n179 B.n96 585
R247 B.n181 B.n180 585
R248 B.n182 B.n95 585
R249 B.n184 B.n183 585
R250 B.n185 B.n94 585
R251 B.n187 B.n186 585
R252 B.n189 B.n91 585
R253 B.n191 B.n190 585
R254 B.n192 B.n90 585
R255 B.n194 B.n193 585
R256 B.n195 B.n89 585
R257 B.n197 B.n196 585
R258 B.n198 B.n88 585
R259 B.n200 B.n199 585
R260 B.n201 B.n87 585
R261 B.n203 B.n202 585
R262 B.n205 B.n204 585
R263 B.n206 B.n83 585
R264 B.n208 B.n207 585
R265 B.n209 B.n82 585
R266 B.n211 B.n210 585
R267 B.n212 B.n81 585
R268 B.n214 B.n213 585
R269 B.n215 B.n80 585
R270 B.n217 B.n216 585
R271 B.n218 B.n79 585
R272 B.n220 B.n219 585
R273 B.n221 B.n78 585
R274 B.n223 B.n222 585
R275 B.n224 B.n77 585
R276 B.n226 B.n225 585
R277 B.n227 B.n76 585
R278 B.n229 B.n228 585
R279 B.n230 B.n75 585
R280 B.n232 B.n231 585
R281 B.n233 B.n74 585
R282 B.n235 B.n234 585
R283 B.n236 B.n73 585
R284 B.n154 B.n153 585
R285 B.n152 B.n105 585
R286 B.n151 B.n150 585
R287 B.n149 B.n106 585
R288 B.n148 B.n147 585
R289 B.n146 B.n107 585
R290 B.n145 B.n144 585
R291 B.n143 B.n108 585
R292 B.n142 B.n141 585
R293 B.n140 B.n109 585
R294 B.n139 B.n138 585
R295 B.n137 B.n110 585
R296 B.n136 B.n135 585
R297 B.n134 B.n111 585
R298 B.n133 B.n132 585
R299 B.n131 B.n112 585
R300 B.n130 B.n129 585
R301 B.n128 B.n113 585
R302 B.n127 B.n126 585
R303 B.n125 B.n114 585
R304 B.n124 B.n123 585
R305 B.n122 B.n115 585
R306 B.n121 B.n120 585
R307 B.n119 B.n116 585
R308 B.n118 B.n117 585
R309 B.n2 B.n0 585
R310 B.n437 B.n1 585
R311 B.n436 B.n435 585
R312 B.n434 B.n3 585
R313 B.n433 B.n432 585
R314 B.n431 B.n4 585
R315 B.n430 B.n429 585
R316 B.n428 B.n5 585
R317 B.n427 B.n426 585
R318 B.n425 B.n6 585
R319 B.n424 B.n423 585
R320 B.n422 B.n7 585
R321 B.n421 B.n420 585
R322 B.n419 B.n8 585
R323 B.n418 B.n417 585
R324 B.n416 B.n9 585
R325 B.n415 B.n414 585
R326 B.n413 B.n10 585
R327 B.n412 B.n411 585
R328 B.n410 B.n11 585
R329 B.n409 B.n408 585
R330 B.n407 B.n12 585
R331 B.n406 B.n405 585
R332 B.n404 B.n13 585
R333 B.n403 B.n402 585
R334 B.n401 B.n14 585
R335 B.n400 B.n399 585
R336 B.n439 B.n438 585
R337 B.n155 B.n154 574.183
R338 B.n400 B.n15 574.183
R339 B.n238 B.n73 574.183
R340 B.n317 B.n316 574.183
R341 B.n84 B.t6 313.317
R342 B.n92 B.t0 313.317
R343 B.n26 B.t9 313.317
R344 B.n34 B.t3 313.317
R345 B.n154 B.n105 163.367
R346 B.n150 B.n105 163.367
R347 B.n150 B.n149 163.367
R348 B.n149 B.n148 163.367
R349 B.n148 B.n107 163.367
R350 B.n144 B.n107 163.367
R351 B.n144 B.n143 163.367
R352 B.n143 B.n142 163.367
R353 B.n142 B.n109 163.367
R354 B.n138 B.n109 163.367
R355 B.n138 B.n137 163.367
R356 B.n137 B.n136 163.367
R357 B.n136 B.n111 163.367
R358 B.n132 B.n111 163.367
R359 B.n132 B.n131 163.367
R360 B.n131 B.n130 163.367
R361 B.n130 B.n113 163.367
R362 B.n126 B.n113 163.367
R363 B.n126 B.n125 163.367
R364 B.n125 B.n124 163.367
R365 B.n124 B.n115 163.367
R366 B.n120 B.n115 163.367
R367 B.n120 B.n119 163.367
R368 B.n119 B.n118 163.367
R369 B.n118 B.n2 163.367
R370 B.n438 B.n2 163.367
R371 B.n438 B.n437 163.367
R372 B.n437 B.n436 163.367
R373 B.n436 B.n3 163.367
R374 B.n432 B.n3 163.367
R375 B.n432 B.n431 163.367
R376 B.n431 B.n430 163.367
R377 B.n430 B.n5 163.367
R378 B.n426 B.n5 163.367
R379 B.n426 B.n425 163.367
R380 B.n425 B.n424 163.367
R381 B.n424 B.n7 163.367
R382 B.n420 B.n7 163.367
R383 B.n420 B.n419 163.367
R384 B.n419 B.n418 163.367
R385 B.n418 B.n9 163.367
R386 B.n414 B.n9 163.367
R387 B.n414 B.n413 163.367
R388 B.n413 B.n412 163.367
R389 B.n412 B.n11 163.367
R390 B.n408 B.n11 163.367
R391 B.n408 B.n407 163.367
R392 B.n407 B.n406 163.367
R393 B.n406 B.n13 163.367
R394 B.n402 B.n13 163.367
R395 B.n402 B.n401 163.367
R396 B.n401 B.n400 163.367
R397 B.n156 B.n155 163.367
R398 B.n156 B.n103 163.367
R399 B.n160 B.n103 163.367
R400 B.n161 B.n160 163.367
R401 B.n162 B.n161 163.367
R402 B.n162 B.n101 163.367
R403 B.n166 B.n101 163.367
R404 B.n167 B.n166 163.367
R405 B.n168 B.n167 163.367
R406 B.n168 B.n99 163.367
R407 B.n172 B.n99 163.367
R408 B.n173 B.n172 163.367
R409 B.n174 B.n173 163.367
R410 B.n174 B.n97 163.367
R411 B.n178 B.n97 163.367
R412 B.n179 B.n178 163.367
R413 B.n180 B.n179 163.367
R414 B.n180 B.n95 163.367
R415 B.n184 B.n95 163.367
R416 B.n185 B.n184 163.367
R417 B.n186 B.n185 163.367
R418 B.n186 B.n91 163.367
R419 B.n191 B.n91 163.367
R420 B.n192 B.n191 163.367
R421 B.n193 B.n192 163.367
R422 B.n193 B.n89 163.367
R423 B.n197 B.n89 163.367
R424 B.n198 B.n197 163.367
R425 B.n199 B.n198 163.367
R426 B.n199 B.n87 163.367
R427 B.n203 B.n87 163.367
R428 B.n204 B.n203 163.367
R429 B.n204 B.n83 163.367
R430 B.n208 B.n83 163.367
R431 B.n209 B.n208 163.367
R432 B.n210 B.n209 163.367
R433 B.n210 B.n81 163.367
R434 B.n214 B.n81 163.367
R435 B.n215 B.n214 163.367
R436 B.n216 B.n215 163.367
R437 B.n216 B.n79 163.367
R438 B.n220 B.n79 163.367
R439 B.n221 B.n220 163.367
R440 B.n222 B.n221 163.367
R441 B.n222 B.n77 163.367
R442 B.n226 B.n77 163.367
R443 B.n227 B.n226 163.367
R444 B.n228 B.n227 163.367
R445 B.n228 B.n75 163.367
R446 B.n232 B.n75 163.367
R447 B.n233 B.n232 163.367
R448 B.n234 B.n233 163.367
R449 B.n234 B.n73 163.367
R450 B.n239 B.n238 163.367
R451 B.n240 B.n239 163.367
R452 B.n240 B.n71 163.367
R453 B.n244 B.n71 163.367
R454 B.n245 B.n244 163.367
R455 B.n246 B.n245 163.367
R456 B.n246 B.n69 163.367
R457 B.n250 B.n69 163.367
R458 B.n251 B.n250 163.367
R459 B.n252 B.n251 163.367
R460 B.n252 B.n67 163.367
R461 B.n256 B.n67 163.367
R462 B.n257 B.n256 163.367
R463 B.n258 B.n257 163.367
R464 B.n258 B.n65 163.367
R465 B.n262 B.n65 163.367
R466 B.n263 B.n262 163.367
R467 B.n264 B.n263 163.367
R468 B.n264 B.n63 163.367
R469 B.n268 B.n63 163.367
R470 B.n269 B.n268 163.367
R471 B.n270 B.n269 163.367
R472 B.n270 B.n61 163.367
R473 B.n274 B.n61 163.367
R474 B.n275 B.n274 163.367
R475 B.n276 B.n275 163.367
R476 B.n276 B.n59 163.367
R477 B.n280 B.n59 163.367
R478 B.n281 B.n280 163.367
R479 B.n282 B.n281 163.367
R480 B.n282 B.n57 163.367
R481 B.n286 B.n57 163.367
R482 B.n287 B.n286 163.367
R483 B.n288 B.n287 163.367
R484 B.n288 B.n55 163.367
R485 B.n292 B.n55 163.367
R486 B.n293 B.n292 163.367
R487 B.n294 B.n293 163.367
R488 B.n294 B.n53 163.367
R489 B.n298 B.n53 163.367
R490 B.n299 B.n298 163.367
R491 B.n300 B.n299 163.367
R492 B.n300 B.n51 163.367
R493 B.n304 B.n51 163.367
R494 B.n305 B.n304 163.367
R495 B.n306 B.n305 163.367
R496 B.n306 B.n49 163.367
R497 B.n310 B.n49 163.367
R498 B.n311 B.n310 163.367
R499 B.n312 B.n311 163.367
R500 B.n312 B.n47 163.367
R501 B.n316 B.n47 163.367
R502 B.n396 B.n15 163.367
R503 B.n396 B.n395 163.367
R504 B.n395 B.n394 163.367
R505 B.n394 B.n17 163.367
R506 B.n390 B.n17 163.367
R507 B.n390 B.n389 163.367
R508 B.n389 B.n388 163.367
R509 B.n388 B.n19 163.367
R510 B.n384 B.n19 163.367
R511 B.n384 B.n383 163.367
R512 B.n383 B.n382 163.367
R513 B.n382 B.n21 163.367
R514 B.n378 B.n21 163.367
R515 B.n378 B.n377 163.367
R516 B.n377 B.n376 163.367
R517 B.n376 B.n23 163.367
R518 B.n372 B.n23 163.367
R519 B.n372 B.n371 163.367
R520 B.n371 B.n370 163.367
R521 B.n370 B.n25 163.367
R522 B.n366 B.n25 163.367
R523 B.n366 B.n365 163.367
R524 B.n365 B.n29 163.367
R525 B.n361 B.n29 163.367
R526 B.n361 B.n360 163.367
R527 B.n360 B.n359 163.367
R528 B.n359 B.n31 163.367
R529 B.n355 B.n31 163.367
R530 B.n355 B.n354 163.367
R531 B.n354 B.n353 163.367
R532 B.n353 B.n33 163.367
R533 B.n348 B.n33 163.367
R534 B.n348 B.n347 163.367
R535 B.n347 B.n346 163.367
R536 B.n346 B.n37 163.367
R537 B.n342 B.n37 163.367
R538 B.n342 B.n341 163.367
R539 B.n341 B.n340 163.367
R540 B.n340 B.n39 163.367
R541 B.n336 B.n39 163.367
R542 B.n336 B.n335 163.367
R543 B.n335 B.n334 163.367
R544 B.n334 B.n41 163.367
R545 B.n330 B.n41 163.367
R546 B.n330 B.n329 163.367
R547 B.n329 B.n328 163.367
R548 B.n328 B.n43 163.367
R549 B.n324 B.n43 163.367
R550 B.n324 B.n323 163.367
R551 B.n323 B.n322 163.367
R552 B.n322 B.n45 163.367
R553 B.n318 B.n45 163.367
R554 B.n318 B.n317 163.367
R555 B.n84 B.t8 142.934
R556 B.n34 B.t4 142.934
R557 B.n92 B.t2 142.928
R558 B.n26 B.t10 142.928
R559 B.n85 B.t7 113.067
R560 B.n35 B.t5 113.067
R561 B.n93 B.t1 113.061
R562 B.n27 B.t11 113.061
R563 B.n86 B.n85 59.5399
R564 B.n188 B.n93 59.5399
R565 B.n28 B.n27 59.5399
R566 B.n350 B.n35 59.5399
R567 B.n399 B.n398 37.3078
R568 B.n315 B.n46 37.3078
R569 B.n237 B.n236 37.3078
R570 B.n153 B.n104 37.3078
R571 B.n85 B.n84 29.8672
R572 B.n93 B.n92 29.8672
R573 B.n27 B.n26 29.8672
R574 B.n35 B.n34 29.8672
R575 B B.n439 18.0485
R576 B.n398 B.n397 10.6151
R577 B.n397 B.n16 10.6151
R578 B.n393 B.n16 10.6151
R579 B.n393 B.n392 10.6151
R580 B.n392 B.n391 10.6151
R581 B.n391 B.n18 10.6151
R582 B.n387 B.n18 10.6151
R583 B.n387 B.n386 10.6151
R584 B.n386 B.n385 10.6151
R585 B.n385 B.n20 10.6151
R586 B.n381 B.n20 10.6151
R587 B.n381 B.n380 10.6151
R588 B.n380 B.n379 10.6151
R589 B.n379 B.n22 10.6151
R590 B.n375 B.n22 10.6151
R591 B.n375 B.n374 10.6151
R592 B.n374 B.n373 10.6151
R593 B.n373 B.n24 10.6151
R594 B.n369 B.n24 10.6151
R595 B.n369 B.n368 10.6151
R596 B.n368 B.n367 10.6151
R597 B.n364 B.n363 10.6151
R598 B.n363 B.n362 10.6151
R599 B.n362 B.n30 10.6151
R600 B.n358 B.n30 10.6151
R601 B.n358 B.n357 10.6151
R602 B.n357 B.n356 10.6151
R603 B.n356 B.n32 10.6151
R604 B.n352 B.n32 10.6151
R605 B.n352 B.n351 10.6151
R606 B.n349 B.n36 10.6151
R607 B.n345 B.n36 10.6151
R608 B.n345 B.n344 10.6151
R609 B.n344 B.n343 10.6151
R610 B.n343 B.n38 10.6151
R611 B.n339 B.n38 10.6151
R612 B.n339 B.n338 10.6151
R613 B.n338 B.n337 10.6151
R614 B.n337 B.n40 10.6151
R615 B.n333 B.n40 10.6151
R616 B.n333 B.n332 10.6151
R617 B.n332 B.n331 10.6151
R618 B.n331 B.n42 10.6151
R619 B.n327 B.n42 10.6151
R620 B.n327 B.n326 10.6151
R621 B.n326 B.n325 10.6151
R622 B.n325 B.n44 10.6151
R623 B.n321 B.n44 10.6151
R624 B.n321 B.n320 10.6151
R625 B.n320 B.n319 10.6151
R626 B.n319 B.n46 10.6151
R627 B.n237 B.n72 10.6151
R628 B.n241 B.n72 10.6151
R629 B.n242 B.n241 10.6151
R630 B.n243 B.n242 10.6151
R631 B.n243 B.n70 10.6151
R632 B.n247 B.n70 10.6151
R633 B.n248 B.n247 10.6151
R634 B.n249 B.n248 10.6151
R635 B.n249 B.n68 10.6151
R636 B.n253 B.n68 10.6151
R637 B.n254 B.n253 10.6151
R638 B.n255 B.n254 10.6151
R639 B.n255 B.n66 10.6151
R640 B.n259 B.n66 10.6151
R641 B.n260 B.n259 10.6151
R642 B.n261 B.n260 10.6151
R643 B.n261 B.n64 10.6151
R644 B.n265 B.n64 10.6151
R645 B.n266 B.n265 10.6151
R646 B.n267 B.n266 10.6151
R647 B.n267 B.n62 10.6151
R648 B.n271 B.n62 10.6151
R649 B.n272 B.n271 10.6151
R650 B.n273 B.n272 10.6151
R651 B.n273 B.n60 10.6151
R652 B.n277 B.n60 10.6151
R653 B.n278 B.n277 10.6151
R654 B.n279 B.n278 10.6151
R655 B.n279 B.n58 10.6151
R656 B.n283 B.n58 10.6151
R657 B.n284 B.n283 10.6151
R658 B.n285 B.n284 10.6151
R659 B.n285 B.n56 10.6151
R660 B.n289 B.n56 10.6151
R661 B.n290 B.n289 10.6151
R662 B.n291 B.n290 10.6151
R663 B.n291 B.n54 10.6151
R664 B.n295 B.n54 10.6151
R665 B.n296 B.n295 10.6151
R666 B.n297 B.n296 10.6151
R667 B.n297 B.n52 10.6151
R668 B.n301 B.n52 10.6151
R669 B.n302 B.n301 10.6151
R670 B.n303 B.n302 10.6151
R671 B.n303 B.n50 10.6151
R672 B.n307 B.n50 10.6151
R673 B.n308 B.n307 10.6151
R674 B.n309 B.n308 10.6151
R675 B.n309 B.n48 10.6151
R676 B.n313 B.n48 10.6151
R677 B.n314 B.n313 10.6151
R678 B.n315 B.n314 10.6151
R679 B.n157 B.n104 10.6151
R680 B.n158 B.n157 10.6151
R681 B.n159 B.n158 10.6151
R682 B.n159 B.n102 10.6151
R683 B.n163 B.n102 10.6151
R684 B.n164 B.n163 10.6151
R685 B.n165 B.n164 10.6151
R686 B.n165 B.n100 10.6151
R687 B.n169 B.n100 10.6151
R688 B.n170 B.n169 10.6151
R689 B.n171 B.n170 10.6151
R690 B.n171 B.n98 10.6151
R691 B.n175 B.n98 10.6151
R692 B.n176 B.n175 10.6151
R693 B.n177 B.n176 10.6151
R694 B.n177 B.n96 10.6151
R695 B.n181 B.n96 10.6151
R696 B.n182 B.n181 10.6151
R697 B.n183 B.n182 10.6151
R698 B.n183 B.n94 10.6151
R699 B.n187 B.n94 10.6151
R700 B.n190 B.n189 10.6151
R701 B.n190 B.n90 10.6151
R702 B.n194 B.n90 10.6151
R703 B.n195 B.n194 10.6151
R704 B.n196 B.n195 10.6151
R705 B.n196 B.n88 10.6151
R706 B.n200 B.n88 10.6151
R707 B.n201 B.n200 10.6151
R708 B.n202 B.n201 10.6151
R709 B.n206 B.n205 10.6151
R710 B.n207 B.n206 10.6151
R711 B.n207 B.n82 10.6151
R712 B.n211 B.n82 10.6151
R713 B.n212 B.n211 10.6151
R714 B.n213 B.n212 10.6151
R715 B.n213 B.n80 10.6151
R716 B.n217 B.n80 10.6151
R717 B.n218 B.n217 10.6151
R718 B.n219 B.n218 10.6151
R719 B.n219 B.n78 10.6151
R720 B.n223 B.n78 10.6151
R721 B.n224 B.n223 10.6151
R722 B.n225 B.n224 10.6151
R723 B.n225 B.n76 10.6151
R724 B.n229 B.n76 10.6151
R725 B.n230 B.n229 10.6151
R726 B.n231 B.n230 10.6151
R727 B.n231 B.n74 10.6151
R728 B.n235 B.n74 10.6151
R729 B.n236 B.n235 10.6151
R730 B.n153 B.n152 10.6151
R731 B.n152 B.n151 10.6151
R732 B.n151 B.n106 10.6151
R733 B.n147 B.n106 10.6151
R734 B.n147 B.n146 10.6151
R735 B.n146 B.n145 10.6151
R736 B.n145 B.n108 10.6151
R737 B.n141 B.n108 10.6151
R738 B.n141 B.n140 10.6151
R739 B.n140 B.n139 10.6151
R740 B.n139 B.n110 10.6151
R741 B.n135 B.n110 10.6151
R742 B.n135 B.n134 10.6151
R743 B.n134 B.n133 10.6151
R744 B.n133 B.n112 10.6151
R745 B.n129 B.n112 10.6151
R746 B.n129 B.n128 10.6151
R747 B.n128 B.n127 10.6151
R748 B.n127 B.n114 10.6151
R749 B.n123 B.n114 10.6151
R750 B.n123 B.n122 10.6151
R751 B.n122 B.n121 10.6151
R752 B.n121 B.n116 10.6151
R753 B.n117 B.n116 10.6151
R754 B.n117 B.n0 10.6151
R755 B.n435 B.n1 10.6151
R756 B.n435 B.n434 10.6151
R757 B.n434 B.n433 10.6151
R758 B.n433 B.n4 10.6151
R759 B.n429 B.n4 10.6151
R760 B.n429 B.n428 10.6151
R761 B.n428 B.n427 10.6151
R762 B.n427 B.n6 10.6151
R763 B.n423 B.n6 10.6151
R764 B.n423 B.n422 10.6151
R765 B.n422 B.n421 10.6151
R766 B.n421 B.n8 10.6151
R767 B.n417 B.n8 10.6151
R768 B.n417 B.n416 10.6151
R769 B.n416 B.n415 10.6151
R770 B.n415 B.n10 10.6151
R771 B.n411 B.n10 10.6151
R772 B.n411 B.n410 10.6151
R773 B.n410 B.n409 10.6151
R774 B.n409 B.n12 10.6151
R775 B.n405 B.n12 10.6151
R776 B.n405 B.n404 10.6151
R777 B.n404 B.n403 10.6151
R778 B.n403 B.n14 10.6151
R779 B.n399 B.n14 10.6151
R780 B.n367 B.n28 9.36635
R781 B.n350 B.n349 9.36635
R782 B.n188 B.n187 9.36635
R783 B.n205 B.n86 9.36635
R784 B.n439 B.n0 2.81026
R785 B.n439 B.n1 2.81026
R786 B.n364 B.n28 1.24928
R787 B.n351 B.n350 1.24928
R788 B.n189 B.n188 1.24928
R789 B.n202 B.n86 1.24928
C0 VTAIL VDD2 5.09201f
C1 VP VDD2 0.343785f
C2 VTAIL VP 2.88873f
C3 w_n2202_n2064# VDD2 1.51217f
C4 B VDD1 1.22181f
C5 w_n2202_n2064# VTAIL 1.91066f
C6 B VN 0.795136f
C7 VDD1 VN 0.14897f
C8 w_n2202_n2064# VP 3.99764f
C9 B VDD2 1.26291f
C10 VDD1 VDD2 0.895556f
C11 VTAIL B 1.74791f
C12 VTAIL VDD1 5.05011f
C13 VN VDD2 2.69802f
C14 VP B 1.25699f
C15 VP VDD1 2.88692f
C16 VTAIL VN 2.87445f
C17 VP VN 4.36668f
C18 w_n2202_n2064# B 5.93422f
C19 w_n2202_n2064# VDD1 1.47215f
C20 w_n2202_n2064# VN 3.71683f
C21 VDD2 VSUBS 1.093276f
C22 VDD1 VSUBS 1.429951f
C23 VTAIL VSUBS 0.48278f
C24 VN VSUBS 4.27644f
C25 VP VSUBS 1.513461f
C26 B VSUBS 2.622048f
C27 w_n2202_n2064# VSUBS 56.838f
C28 B.n0 VSUBS 0.0041f
C29 B.n1 VSUBS 0.0041f
C30 B.n2 VSUBS 0.006484f
C31 B.n3 VSUBS 0.006484f
C32 B.n4 VSUBS 0.006484f
C33 B.n5 VSUBS 0.006484f
C34 B.n6 VSUBS 0.006484f
C35 B.n7 VSUBS 0.006484f
C36 B.n8 VSUBS 0.006484f
C37 B.n9 VSUBS 0.006484f
C38 B.n10 VSUBS 0.006484f
C39 B.n11 VSUBS 0.006484f
C40 B.n12 VSUBS 0.006484f
C41 B.n13 VSUBS 0.006484f
C42 B.n14 VSUBS 0.006484f
C43 B.n15 VSUBS 0.01691f
C44 B.n16 VSUBS 0.006484f
C45 B.n17 VSUBS 0.006484f
C46 B.n18 VSUBS 0.006484f
C47 B.n19 VSUBS 0.006484f
C48 B.n20 VSUBS 0.006484f
C49 B.n21 VSUBS 0.006484f
C50 B.n22 VSUBS 0.006484f
C51 B.n23 VSUBS 0.006484f
C52 B.n24 VSUBS 0.006484f
C53 B.n25 VSUBS 0.006484f
C54 B.t11 VSUBS 0.145175f
C55 B.t10 VSUBS 0.155753f
C56 B.t9 VSUBS 0.278976f
C57 B.n26 VSUBS 0.086358f
C58 B.n27 VSUBS 0.059868f
C59 B.n28 VSUBS 0.015022f
C60 B.n29 VSUBS 0.006484f
C61 B.n30 VSUBS 0.006484f
C62 B.n31 VSUBS 0.006484f
C63 B.n32 VSUBS 0.006484f
C64 B.n33 VSUBS 0.006484f
C65 B.t5 VSUBS 0.145175f
C66 B.t4 VSUBS 0.155752f
C67 B.t3 VSUBS 0.278976f
C68 B.n34 VSUBS 0.086359f
C69 B.n35 VSUBS 0.059868f
C70 B.n36 VSUBS 0.006484f
C71 B.n37 VSUBS 0.006484f
C72 B.n38 VSUBS 0.006484f
C73 B.n39 VSUBS 0.006484f
C74 B.n40 VSUBS 0.006484f
C75 B.n41 VSUBS 0.006484f
C76 B.n42 VSUBS 0.006484f
C77 B.n43 VSUBS 0.006484f
C78 B.n44 VSUBS 0.006484f
C79 B.n45 VSUBS 0.006484f
C80 B.n46 VSUBS 0.016239f
C81 B.n47 VSUBS 0.006484f
C82 B.n48 VSUBS 0.006484f
C83 B.n49 VSUBS 0.006484f
C84 B.n50 VSUBS 0.006484f
C85 B.n51 VSUBS 0.006484f
C86 B.n52 VSUBS 0.006484f
C87 B.n53 VSUBS 0.006484f
C88 B.n54 VSUBS 0.006484f
C89 B.n55 VSUBS 0.006484f
C90 B.n56 VSUBS 0.006484f
C91 B.n57 VSUBS 0.006484f
C92 B.n58 VSUBS 0.006484f
C93 B.n59 VSUBS 0.006484f
C94 B.n60 VSUBS 0.006484f
C95 B.n61 VSUBS 0.006484f
C96 B.n62 VSUBS 0.006484f
C97 B.n63 VSUBS 0.006484f
C98 B.n64 VSUBS 0.006484f
C99 B.n65 VSUBS 0.006484f
C100 B.n66 VSUBS 0.006484f
C101 B.n67 VSUBS 0.006484f
C102 B.n68 VSUBS 0.006484f
C103 B.n69 VSUBS 0.006484f
C104 B.n70 VSUBS 0.006484f
C105 B.n71 VSUBS 0.006484f
C106 B.n72 VSUBS 0.006484f
C107 B.n73 VSUBS 0.01691f
C108 B.n74 VSUBS 0.006484f
C109 B.n75 VSUBS 0.006484f
C110 B.n76 VSUBS 0.006484f
C111 B.n77 VSUBS 0.006484f
C112 B.n78 VSUBS 0.006484f
C113 B.n79 VSUBS 0.006484f
C114 B.n80 VSUBS 0.006484f
C115 B.n81 VSUBS 0.006484f
C116 B.n82 VSUBS 0.006484f
C117 B.n83 VSUBS 0.006484f
C118 B.t7 VSUBS 0.145175f
C119 B.t8 VSUBS 0.155752f
C120 B.t6 VSUBS 0.278976f
C121 B.n84 VSUBS 0.086359f
C122 B.n85 VSUBS 0.059868f
C123 B.n86 VSUBS 0.015022f
C124 B.n87 VSUBS 0.006484f
C125 B.n88 VSUBS 0.006484f
C126 B.n89 VSUBS 0.006484f
C127 B.n90 VSUBS 0.006484f
C128 B.n91 VSUBS 0.006484f
C129 B.t1 VSUBS 0.145175f
C130 B.t2 VSUBS 0.155753f
C131 B.t0 VSUBS 0.278976f
C132 B.n92 VSUBS 0.086358f
C133 B.n93 VSUBS 0.059868f
C134 B.n94 VSUBS 0.006484f
C135 B.n95 VSUBS 0.006484f
C136 B.n96 VSUBS 0.006484f
C137 B.n97 VSUBS 0.006484f
C138 B.n98 VSUBS 0.006484f
C139 B.n99 VSUBS 0.006484f
C140 B.n100 VSUBS 0.006484f
C141 B.n101 VSUBS 0.006484f
C142 B.n102 VSUBS 0.006484f
C143 B.n103 VSUBS 0.006484f
C144 B.n104 VSUBS 0.01691f
C145 B.n105 VSUBS 0.006484f
C146 B.n106 VSUBS 0.006484f
C147 B.n107 VSUBS 0.006484f
C148 B.n108 VSUBS 0.006484f
C149 B.n109 VSUBS 0.006484f
C150 B.n110 VSUBS 0.006484f
C151 B.n111 VSUBS 0.006484f
C152 B.n112 VSUBS 0.006484f
C153 B.n113 VSUBS 0.006484f
C154 B.n114 VSUBS 0.006484f
C155 B.n115 VSUBS 0.006484f
C156 B.n116 VSUBS 0.006484f
C157 B.n117 VSUBS 0.006484f
C158 B.n118 VSUBS 0.006484f
C159 B.n119 VSUBS 0.006484f
C160 B.n120 VSUBS 0.006484f
C161 B.n121 VSUBS 0.006484f
C162 B.n122 VSUBS 0.006484f
C163 B.n123 VSUBS 0.006484f
C164 B.n124 VSUBS 0.006484f
C165 B.n125 VSUBS 0.006484f
C166 B.n126 VSUBS 0.006484f
C167 B.n127 VSUBS 0.006484f
C168 B.n128 VSUBS 0.006484f
C169 B.n129 VSUBS 0.006484f
C170 B.n130 VSUBS 0.006484f
C171 B.n131 VSUBS 0.006484f
C172 B.n132 VSUBS 0.006484f
C173 B.n133 VSUBS 0.006484f
C174 B.n134 VSUBS 0.006484f
C175 B.n135 VSUBS 0.006484f
C176 B.n136 VSUBS 0.006484f
C177 B.n137 VSUBS 0.006484f
C178 B.n138 VSUBS 0.006484f
C179 B.n139 VSUBS 0.006484f
C180 B.n140 VSUBS 0.006484f
C181 B.n141 VSUBS 0.006484f
C182 B.n142 VSUBS 0.006484f
C183 B.n143 VSUBS 0.006484f
C184 B.n144 VSUBS 0.006484f
C185 B.n145 VSUBS 0.006484f
C186 B.n146 VSUBS 0.006484f
C187 B.n147 VSUBS 0.006484f
C188 B.n148 VSUBS 0.006484f
C189 B.n149 VSUBS 0.006484f
C190 B.n150 VSUBS 0.006484f
C191 B.n151 VSUBS 0.006484f
C192 B.n152 VSUBS 0.006484f
C193 B.n153 VSUBS 0.016272f
C194 B.n154 VSUBS 0.016272f
C195 B.n155 VSUBS 0.01691f
C196 B.n156 VSUBS 0.006484f
C197 B.n157 VSUBS 0.006484f
C198 B.n158 VSUBS 0.006484f
C199 B.n159 VSUBS 0.006484f
C200 B.n160 VSUBS 0.006484f
C201 B.n161 VSUBS 0.006484f
C202 B.n162 VSUBS 0.006484f
C203 B.n163 VSUBS 0.006484f
C204 B.n164 VSUBS 0.006484f
C205 B.n165 VSUBS 0.006484f
C206 B.n166 VSUBS 0.006484f
C207 B.n167 VSUBS 0.006484f
C208 B.n168 VSUBS 0.006484f
C209 B.n169 VSUBS 0.006484f
C210 B.n170 VSUBS 0.006484f
C211 B.n171 VSUBS 0.006484f
C212 B.n172 VSUBS 0.006484f
C213 B.n173 VSUBS 0.006484f
C214 B.n174 VSUBS 0.006484f
C215 B.n175 VSUBS 0.006484f
C216 B.n176 VSUBS 0.006484f
C217 B.n177 VSUBS 0.006484f
C218 B.n178 VSUBS 0.006484f
C219 B.n179 VSUBS 0.006484f
C220 B.n180 VSUBS 0.006484f
C221 B.n181 VSUBS 0.006484f
C222 B.n182 VSUBS 0.006484f
C223 B.n183 VSUBS 0.006484f
C224 B.n184 VSUBS 0.006484f
C225 B.n185 VSUBS 0.006484f
C226 B.n186 VSUBS 0.006484f
C227 B.n187 VSUBS 0.006102f
C228 B.n188 VSUBS 0.015022f
C229 B.n189 VSUBS 0.003623f
C230 B.n190 VSUBS 0.006484f
C231 B.n191 VSUBS 0.006484f
C232 B.n192 VSUBS 0.006484f
C233 B.n193 VSUBS 0.006484f
C234 B.n194 VSUBS 0.006484f
C235 B.n195 VSUBS 0.006484f
C236 B.n196 VSUBS 0.006484f
C237 B.n197 VSUBS 0.006484f
C238 B.n198 VSUBS 0.006484f
C239 B.n199 VSUBS 0.006484f
C240 B.n200 VSUBS 0.006484f
C241 B.n201 VSUBS 0.006484f
C242 B.n202 VSUBS 0.003623f
C243 B.n203 VSUBS 0.006484f
C244 B.n204 VSUBS 0.006484f
C245 B.n205 VSUBS 0.006102f
C246 B.n206 VSUBS 0.006484f
C247 B.n207 VSUBS 0.006484f
C248 B.n208 VSUBS 0.006484f
C249 B.n209 VSUBS 0.006484f
C250 B.n210 VSUBS 0.006484f
C251 B.n211 VSUBS 0.006484f
C252 B.n212 VSUBS 0.006484f
C253 B.n213 VSUBS 0.006484f
C254 B.n214 VSUBS 0.006484f
C255 B.n215 VSUBS 0.006484f
C256 B.n216 VSUBS 0.006484f
C257 B.n217 VSUBS 0.006484f
C258 B.n218 VSUBS 0.006484f
C259 B.n219 VSUBS 0.006484f
C260 B.n220 VSUBS 0.006484f
C261 B.n221 VSUBS 0.006484f
C262 B.n222 VSUBS 0.006484f
C263 B.n223 VSUBS 0.006484f
C264 B.n224 VSUBS 0.006484f
C265 B.n225 VSUBS 0.006484f
C266 B.n226 VSUBS 0.006484f
C267 B.n227 VSUBS 0.006484f
C268 B.n228 VSUBS 0.006484f
C269 B.n229 VSUBS 0.006484f
C270 B.n230 VSUBS 0.006484f
C271 B.n231 VSUBS 0.006484f
C272 B.n232 VSUBS 0.006484f
C273 B.n233 VSUBS 0.006484f
C274 B.n234 VSUBS 0.006484f
C275 B.n235 VSUBS 0.006484f
C276 B.n236 VSUBS 0.01691f
C277 B.n237 VSUBS 0.016272f
C278 B.n238 VSUBS 0.016272f
C279 B.n239 VSUBS 0.006484f
C280 B.n240 VSUBS 0.006484f
C281 B.n241 VSUBS 0.006484f
C282 B.n242 VSUBS 0.006484f
C283 B.n243 VSUBS 0.006484f
C284 B.n244 VSUBS 0.006484f
C285 B.n245 VSUBS 0.006484f
C286 B.n246 VSUBS 0.006484f
C287 B.n247 VSUBS 0.006484f
C288 B.n248 VSUBS 0.006484f
C289 B.n249 VSUBS 0.006484f
C290 B.n250 VSUBS 0.006484f
C291 B.n251 VSUBS 0.006484f
C292 B.n252 VSUBS 0.006484f
C293 B.n253 VSUBS 0.006484f
C294 B.n254 VSUBS 0.006484f
C295 B.n255 VSUBS 0.006484f
C296 B.n256 VSUBS 0.006484f
C297 B.n257 VSUBS 0.006484f
C298 B.n258 VSUBS 0.006484f
C299 B.n259 VSUBS 0.006484f
C300 B.n260 VSUBS 0.006484f
C301 B.n261 VSUBS 0.006484f
C302 B.n262 VSUBS 0.006484f
C303 B.n263 VSUBS 0.006484f
C304 B.n264 VSUBS 0.006484f
C305 B.n265 VSUBS 0.006484f
C306 B.n266 VSUBS 0.006484f
C307 B.n267 VSUBS 0.006484f
C308 B.n268 VSUBS 0.006484f
C309 B.n269 VSUBS 0.006484f
C310 B.n270 VSUBS 0.006484f
C311 B.n271 VSUBS 0.006484f
C312 B.n272 VSUBS 0.006484f
C313 B.n273 VSUBS 0.006484f
C314 B.n274 VSUBS 0.006484f
C315 B.n275 VSUBS 0.006484f
C316 B.n276 VSUBS 0.006484f
C317 B.n277 VSUBS 0.006484f
C318 B.n278 VSUBS 0.006484f
C319 B.n279 VSUBS 0.006484f
C320 B.n280 VSUBS 0.006484f
C321 B.n281 VSUBS 0.006484f
C322 B.n282 VSUBS 0.006484f
C323 B.n283 VSUBS 0.006484f
C324 B.n284 VSUBS 0.006484f
C325 B.n285 VSUBS 0.006484f
C326 B.n286 VSUBS 0.006484f
C327 B.n287 VSUBS 0.006484f
C328 B.n288 VSUBS 0.006484f
C329 B.n289 VSUBS 0.006484f
C330 B.n290 VSUBS 0.006484f
C331 B.n291 VSUBS 0.006484f
C332 B.n292 VSUBS 0.006484f
C333 B.n293 VSUBS 0.006484f
C334 B.n294 VSUBS 0.006484f
C335 B.n295 VSUBS 0.006484f
C336 B.n296 VSUBS 0.006484f
C337 B.n297 VSUBS 0.006484f
C338 B.n298 VSUBS 0.006484f
C339 B.n299 VSUBS 0.006484f
C340 B.n300 VSUBS 0.006484f
C341 B.n301 VSUBS 0.006484f
C342 B.n302 VSUBS 0.006484f
C343 B.n303 VSUBS 0.006484f
C344 B.n304 VSUBS 0.006484f
C345 B.n305 VSUBS 0.006484f
C346 B.n306 VSUBS 0.006484f
C347 B.n307 VSUBS 0.006484f
C348 B.n308 VSUBS 0.006484f
C349 B.n309 VSUBS 0.006484f
C350 B.n310 VSUBS 0.006484f
C351 B.n311 VSUBS 0.006484f
C352 B.n312 VSUBS 0.006484f
C353 B.n313 VSUBS 0.006484f
C354 B.n314 VSUBS 0.006484f
C355 B.n315 VSUBS 0.016942f
C356 B.n316 VSUBS 0.016272f
C357 B.n317 VSUBS 0.01691f
C358 B.n318 VSUBS 0.006484f
C359 B.n319 VSUBS 0.006484f
C360 B.n320 VSUBS 0.006484f
C361 B.n321 VSUBS 0.006484f
C362 B.n322 VSUBS 0.006484f
C363 B.n323 VSUBS 0.006484f
C364 B.n324 VSUBS 0.006484f
C365 B.n325 VSUBS 0.006484f
C366 B.n326 VSUBS 0.006484f
C367 B.n327 VSUBS 0.006484f
C368 B.n328 VSUBS 0.006484f
C369 B.n329 VSUBS 0.006484f
C370 B.n330 VSUBS 0.006484f
C371 B.n331 VSUBS 0.006484f
C372 B.n332 VSUBS 0.006484f
C373 B.n333 VSUBS 0.006484f
C374 B.n334 VSUBS 0.006484f
C375 B.n335 VSUBS 0.006484f
C376 B.n336 VSUBS 0.006484f
C377 B.n337 VSUBS 0.006484f
C378 B.n338 VSUBS 0.006484f
C379 B.n339 VSUBS 0.006484f
C380 B.n340 VSUBS 0.006484f
C381 B.n341 VSUBS 0.006484f
C382 B.n342 VSUBS 0.006484f
C383 B.n343 VSUBS 0.006484f
C384 B.n344 VSUBS 0.006484f
C385 B.n345 VSUBS 0.006484f
C386 B.n346 VSUBS 0.006484f
C387 B.n347 VSUBS 0.006484f
C388 B.n348 VSUBS 0.006484f
C389 B.n349 VSUBS 0.006102f
C390 B.n350 VSUBS 0.015022f
C391 B.n351 VSUBS 0.003623f
C392 B.n352 VSUBS 0.006484f
C393 B.n353 VSUBS 0.006484f
C394 B.n354 VSUBS 0.006484f
C395 B.n355 VSUBS 0.006484f
C396 B.n356 VSUBS 0.006484f
C397 B.n357 VSUBS 0.006484f
C398 B.n358 VSUBS 0.006484f
C399 B.n359 VSUBS 0.006484f
C400 B.n360 VSUBS 0.006484f
C401 B.n361 VSUBS 0.006484f
C402 B.n362 VSUBS 0.006484f
C403 B.n363 VSUBS 0.006484f
C404 B.n364 VSUBS 0.003623f
C405 B.n365 VSUBS 0.006484f
C406 B.n366 VSUBS 0.006484f
C407 B.n367 VSUBS 0.006102f
C408 B.n368 VSUBS 0.006484f
C409 B.n369 VSUBS 0.006484f
C410 B.n370 VSUBS 0.006484f
C411 B.n371 VSUBS 0.006484f
C412 B.n372 VSUBS 0.006484f
C413 B.n373 VSUBS 0.006484f
C414 B.n374 VSUBS 0.006484f
C415 B.n375 VSUBS 0.006484f
C416 B.n376 VSUBS 0.006484f
C417 B.n377 VSUBS 0.006484f
C418 B.n378 VSUBS 0.006484f
C419 B.n379 VSUBS 0.006484f
C420 B.n380 VSUBS 0.006484f
C421 B.n381 VSUBS 0.006484f
C422 B.n382 VSUBS 0.006484f
C423 B.n383 VSUBS 0.006484f
C424 B.n384 VSUBS 0.006484f
C425 B.n385 VSUBS 0.006484f
C426 B.n386 VSUBS 0.006484f
C427 B.n387 VSUBS 0.006484f
C428 B.n388 VSUBS 0.006484f
C429 B.n389 VSUBS 0.006484f
C430 B.n390 VSUBS 0.006484f
C431 B.n391 VSUBS 0.006484f
C432 B.n392 VSUBS 0.006484f
C433 B.n393 VSUBS 0.006484f
C434 B.n394 VSUBS 0.006484f
C435 B.n395 VSUBS 0.006484f
C436 B.n396 VSUBS 0.006484f
C437 B.n397 VSUBS 0.006484f
C438 B.n398 VSUBS 0.01691f
C439 B.n399 VSUBS 0.016272f
C440 B.n400 VSUBS 0.016272f
C441 B.n401 VSUBS 0.006484f
C442 B.n402 VSUBS 0.006484f
C443 B.n403 VSUBS 0.006484f
C444 B.n404 VSUBS 0.006484f
C445 B.n405 VSUBS 0.006484f
C446 B.n406 VSUBS 0.006484f
C447 B.n407 VSUBS 0.006484f
C448 B.n408 VSUBS 0.006484f
C449 B.n409 VSUBS 0.006484f
C450 B.n410 VSUBS 0.006484f
C451 B.n411 VSUBS 0.006484f
C452 B.n412 VSUBS 0.006484f
C453 B.n413 VSUBS 0.006484f
C454 B.n414 VSUBS 0.006484f
C455 B.n415 VSUBS 0.006484f
C456 B.n416 VSUBS 0.006484f
C457 B.n417 VSUBS 0.006484f
C458 B.n418 VSUBS 0.006484f
C459 B.n419 VSUBS 0.006484f
C460 B.n420 VSUBS 0.006484f
C461 B.n421 VSUBS 0.006484f
C462 B.n422 VSUBS 0.006484f
C463 B.n423 VSUBS 0.006484f
C464 B.n424 VSUBS 0.006484f
C465 B.n425 VSUBS 0.006484f
C466 B.n426 VSUBS 0.006484f
C467 B.n427 VSUBS 0.006484f
C468 B.n428 VSUBS 0.006484f
C469 B.n429 VSUBS 0.006484f
C470 B.n430 VSUBS 0.006484f
C471 B.n431 VSUBS 0.006484f
C472 B.n432 VSUBS 0.006484f
C473 B.n433 VSUBS 0.006484f
C474 B.n434 VSUBS 0.006484f
C475 B.n435 VSUBS 0.006484f
C476 B.n436 VSUBS 0.006484f
C477 B.n437 VSUBS 0.006484f
C478 B.n438 VSUBS 0.006484f
C479 B.n439 VSUBS 0.014681f
C480 VDD2.t2 VSUBS 0.862977f
C481 VDD2.t1 VSUBS 0.096857f
C482 VDD2.t5 VSUBS 0.096857f
C483 VDD2.n0 VSUBS 0.642213f
C484 VDD2.n1 VSUBS 2.01012f
C485 VDD2.t3 VSUBS 0.858835f
C486 VDD2.n2 VSUBS 1.83982f
C487 VDD2.t0 VSUBS 0.096857f
C488 VDD2.t4 VSUBS 0.096857f
C489 VDD2.n3 VSUBS 0.642192f
C490 VN.n0 VSUBS 0.053248f
C491 VN.t0 VSUBS 0.9293f
C492 VN.n1 VSUBS 0.081813f
C493 VN.t3 VSUBS 1.04975f
C494 VN.t4 VSUBS 0.9293f
C495 VN.n2 VSUBS 0.458006f
C496 VN.n3 VSUBS 0.482928f
C497 VN.n4 VSUBS 0.278981f
C498 VN.n5 VSUBS 0.053248f
C499 VN.n6 VSUBS 0.043279f
C500 VN.n7 VSUBS 0.083613f
C501 VN.n8 VSUBS 0.471378f
C502 VN.n9 VSUBS 0.047208f
C503 VN.n10 VSUBS 0.053248f
C504 VN.t2 VSUBS 0.9293f
C505 VN.n11 VSUBS 0.081813f
C506 VN.t1 VSUBS 1.04975f
C507 VN.t5 VSUBS 0.9293f
C508 VN.n12 VSUBS 0.458006f
C509 VN.n13 VSUBS 0.482928f
C510 VN.n14 VSUBS 0.278981f
C511 VN.n15 VSUBS 0.053248f
C512 VN.n16 VSUBS 0.043279f
C513 VN.n17 VSUBS 0.083613f
C514 VN.n18 VSUBS 0.471378f
C515 VN.n19 VSUBS 1.90778f
C516 VDD1.t5 VSUBS 0.876411f
C517 VDD1.t0 VSUBS 0.875829f
C518 VDD1.t2 VSUBS 0.098299f
C519 VDD1.t3 VSUBS 0.098299f
C520 VDD1.n0 VSUBS 0.651777f
C521 VDD1.n1 VSUBS 2.11745f
C522 VDD1.t1 VSUBS 0.098299f
C523 VDD1.t4 VSUBS 0.098299f
C524 VDD1.n2 VSUBS 0.650447f
C525 VDD1.n3 VSUBS 1.86679f
C526 VTAIL.t1 VSUBS 0.11345f
C527 VTAIL.t2 VSUBS 0.11345f
C528 VTAIL.n0 VSUBS 0.670388f
C529 VTAIL.n1 VSUBS 0.568782f
C530 VTAIL.t11 VSUBS 0.920747f
C531 VTAIL.n2 VSUBS 0.706972f
C532 VTAIL.t8 VSUBS 0.11345f
C533 VTAIL.t7 VSUBS 0.11345f
C534 VTAIL.n3 VSUBS 0.670388f
C535 VTAIL.n4 VSUBS 1.53103f
C536 VTAIL.t0 VSUBS 0.11345f
C537 VTAIL.t4 VSUBS 0.11345f
C538 VTAIL.n5 VSUBS 0.670392f
C539 VTAIL.n6 VSUBS 1.53102f
C540 VTAIL.t5 VSUBS 0.92075f
C541 VTAIL.n7 VSUBS 0.706968f
C542 VTAIL.t6 VSUBS 0.11345f
C543 VTAIL.t9 VSUBS 0.11345f
C544 VTAIL.n8 VSUBS 0.670392f
C545 VTAIL.n9 VSUBS 0.647918f
C546 VTAIL.t10 VSUBS 0.920743f
C547 VTAIL.n10 VSUBS 1.47801f
C548 VTAIL.t3 VSUBS 0.920747f
C549 VTAIL.n11 VSUBS 1.44508f
C550 VP.n0 VSUBS 0.055495f
C551 VP.t2 VSUBS 0.968508f
C552 VP.n1 VSUBS 0.085265f
C553 VP.n2 VSUBS 0.055495f
C554 VP.t5 VSUBS 0.968508f
C555 VP.n3 VSUBS 0.491265f
C556 VP.n4 VSUBS 0.055495f
C557 VP.t1 VSUBS 0.968508f
C558 VP.n5 VSUBS 0.085265f
C559 VP.t0 VSUBS 1.09404f
C560 VP.t4 VSUBS 0.968508f
C561 VP.n6 VSUBS 0.47733f
C562 VP.n7 VSUBS 0.503303f
C563 VP.n8 VSUBS 0.290752f
C564 VP.n9 VSUBS 0.055495f
C565 VP.n10 VSUBS 0.045105f
C566 VP.n11 VSUBS 0.08714f
C567 VP.n12 VSUBS 0.491265f
C568 VP.n13 VSUBS 1.95162f
C569 VP.n14 VSUBS 2.00398f
C570 VP.n15 VSUBS 0.055495f
C571 VP.n16 VSUBS 0.08714f
C572 VP.n17 VSUBS 0.045105f
C573 VP.t3 VSUBS 0.968508f
C574 VP.n18 VSUBS 0.394549f
C575 VP.n19 VSUBS 0.085265f
C576 VP.n20 VSUBS 0.055495f
C577 VP.n21 VSUBS 0.055495f
C578 VP.n22 VSUBS 0.055495f
C579 VP.n23 VSUBS 0.045105f
C580 VP.n24 VSUBS 0.08714f
C581 VP.n25 VSUBS 0.491265f
C582 VP.n26 VSUBS 0.049199f
.ends

