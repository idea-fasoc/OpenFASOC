* NGSPICE file created from diff_pair_sample_1393.ext - technology: sky130A

.subckt diff_pair_sample_1393 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t14 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=2.9568 ps=18.25 w=17.92 l=3.44
X1 VDD1.t9 VP.t0 VTAIL.t7 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X2 VDD1.t8 VP.t1 VTAIL.t4 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=2.9568 ps=18.25 w=17.92 l=3.44
X3 VDD1.t7 VP.t2 VTAIL.t9 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=2.9568 ps=18.25 w=17.92 l=3.44
X4 VTAIL.t6 VP.t3 VDD1.t6 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X5 B.t11 B.t9 B.t10 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=0 ps=0 w=17.92 l=3.44
X6 VTAIL.t3 VP.t4 VDD1.t5 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X7 VDD1.t4 VP.t5 VTAIL.t1 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=6.9888 ps=36.62 w=17.92 l=3.44
X8 VDD1.t3 VP.t6 VTAIL.t2 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=6.9888 ps=36.62 w=17.92 l=3.44
X9 VTAIL.t5 VP.t7 VDD1.t2 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X10 VDD2.t8 VN.t1 VTAIL.t12 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=6.9888 ps=36.62 w=17.92 l=3.44
X11 VDD2.t7 VN.t2 VTAIL.t11 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X12 VTAIL.t17 VN.t3 VDD2.t6 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X13 B.t8 B.t6 B.t7 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=0 ps=0 w=17.92 l=3.44
X14 VTAIL.t16 VN.t4 VDD2.t5 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X15 VDD1.t1 VP.t8 VTAIL.t0 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X16 VTAIL.t19 VN.t5 VDD2.t4 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X17 VTAIL.t18 VN.t6 VDD2.t3 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X18 VDD2.t2 VN.t7 VTAIL.t10 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=6.9888 ps=36.62 w=17.92 l=3.44
X19 VTAIL.t8 VP.t9 VDD1.t0 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X20 VDD2.t1 VN.t8 VTAIL.t15 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=2.9568 ps=18.25 w=17.92 l=3.44
X21 B.t5 B.t3 B.t4 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=0 ps=0 w=17.92 l=3.44
X22 VDD2.t0 VN.t9 VTAIL.t13 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=2.9568 pd=18.25 as=2.9568 ps=18.25 w=17.92 l=3.44
X23 B.t2 B.t0 B.t1 w_n5494_n4552# sky130_fd_pr__pfet_01v8 ad=6.9888 pd=36.62 as=0 ps=0 w=17.92 l=3.44
R0 VN.n102 VN.n101 161.3
R1 VN.n100 VN.n53 161.3
R2 VN.n99 VN.n98 161.3
R3 VN.n97 VN.n54 161.3
R4 VN.n96 VN.n95 161.3
R5 VN.n94 VN.n55 161.3
R6 VN.n93 VN.n92 161.3
R7 VN.n91 VN.n90 161.3
R8 VN.n89 VN.n57 161.3
R9 VN.n88 VN.n87 161.3
R10 VN.n86 VN.n58 161.3
R11 VN.n85 VN.n84 161.3
R12 VN.n83 VN.n59 161.3
R13 VN.n82 VN.n81 161.3
R14 VN.n80 VN.n60 161.3
R15 VN.n79 VN.n78 161.3
R16 VN.n77 VN.n61 161.3
R17 VN.n76 VN.n75 161.3
R18 VN.n74 VN.n63 161.3
R19 VN.n73 VN.n72 161.3
R20 VN.n71 VN.n64 161.3
R21 VN.n70 VN.n69 161.3
R22 VN.n68 VN.n65 161.3
R23 VN.n50 VN.n49 161.3
R24 VN.n48 VN.n1 161.3
R25 VN.n47 VN.n46 161.3
R26 VN.n45 VN.n2 161.3
R27 VN.n44 VN.n43 161.3
R28 VN.n42 VN.n3 161.3
R29 VN.n41 VN.n40 161.3
R30 VN.n39 VN.n38 161.3
R31 VN.n37 VN.n5 161.3
R32 VN.n36 VN.n35 161.3
R33 VN.n34 VN.n6 161.3
R34 VN.n33 VN.n32 161.3
R35 VN.n31 VN.n7 161.3
R36 VN.n30 VN.n29 161.3
R37 VN.n28 VN.n8 161.3
R38 VN.n27 VN.n26 161.3
R39 VN.n24 VN.n9 161.3
R40 VN.n23 VN.n22 161.3
R41 VN.n21 VN.n10 161.3
R42 VN.n20 VN.n19 161.3
R43 VN.n18 VN.n11 161.3
R44 VN.n17 VN.n16 161.3
R45 VN.n15 VN.n12 161.3
R46 VN.n67 VN.t1 158.196
R47 VN.n14 VN.t0 158.196
R48 VN.n13 VN.t4 125.544
R49 VN.n25 VN.t9 125.544
R50 VN.n4 VN.t3 125.544
R51 VN.n0 VN.t7 125.544
R52 VN.n66 VN.t5 125.544
R53 VN.n62 VN.t2 125.544
R54 VN.n56 VN.t6 125.544
R55 VN.n52 VN.t8 125.544
R56 VN.n51 VN.n0 75.7718
R57 VN.n103 VN.n52 75.7718
R58 VN.n67 VN.n66 73.5205
R59 VN.n14 VN.n13 73.5205
R60 VN VN.n103 62.4714
R61 VN.n19 VN.n10 53.5561
R62 VN.n32 VN.n6 53.5561
R63 VN.n72 VN.n63 53.5561
R64 VN.n84 VN.n58 53.5561
R65 VN.n43 VN.n2 49.6611
R66 VN.n95 VN.n54 49.6611
R67 VN.n47 VN.n2 31.1601
R68 VN.n99 VN.n54 31.1601
R69 VN.n23 VN.n10 27.2651
R70 VN.n32 VN.n31 27.2651
R71 VN.n76 VN.n63 27.2651
R72 VN.n84 VN.n83 27.2651
R73 VN.n17 VN.n12 24.3439
R74 VN.n18 VN.n17 24.3439
R75 VN.n19 VN.n18 24.3439
R76 VN.n24 VN.n23 24.3439
R77 VN.n26 VN.n24 24.3439
R78 VN.n30 VN.n8 24.3439
R79 VN.n31 VN.n30 24.3439
R80 VN.n36 VN.n6 24.3439
R81 VN.n37 VN.n36 24.3439
R82 VN.n38 VN.n37 24.3439
R83 VN.n42 VN.n41 24.3439
R84 VN.n43 VN.n42 24.3439
R85 VN.n48 VN.n47 24.3439
R86 VN.n49 VN.n48 24.3439
R87 VN.n72 VN.n71 24.3439
R88 VN.n71 VN.n70 24.3439
R89 VN.n70 VN.n65 24.3439
R90 VN.n83 VN.n82 24.3439
R91 VN.n82 VN.n60 24.3439
R92 VN.n78 VN.n77 24.3439
R93 VN.n77 VN.n76 24.3439
R94 VN.n95 VN.n94 24.3439
R95 VN.n94 VN.n93 24.3439
R96 VN.n90 VN.n89 24.3439
R97 VN.n89 VN.n88 24.3439
R98 VN.n88 VN.n58 24.3439
R99 VN.n101 VN.n100 24.3439
R100 VN.n100 VN.n99 24.3439
R101 VN.n41 VN.n4 23.3702
R102 VN.n93 VN.n56 23.3702
R103 VN.n49 VN.n0 14.1197
R104 VN.n101 VN.n52 14.1197
R105 VN.n26 VN.n25 12.1722
R106 VN.n25 VN.n8 12.1722
R107 VN.n62 VN.n60 12.1722
R108 VN.n78 VN.n62 12.1722
R109 VN.n68 VN.n67 4.21324
R110 VN.n15 VN.n14 4.21323
R111 VN.n13 VN.n12 0.974237
R112 VN.n38 VN.n4 0.974237
R113 VN.n66 VN.n65 0.974237
R114 VN.n90 VN.n56 0.974237
R115 VN.n103 VN.n102 0.355081
R116 VN.n51 VN.n50 0.355081
R117 VN VN.n51 0.26685
R118 VN.n102 VN.n53 0.189894
R119 VN.n98 VN.n53 0.189894
R120 VN.n98 VN.n97 0.189894
R121 VN.n97 VN.n96 0.189894
R122 VN.n96 VN.n55 0.189894
R123 VN.n92 VN.n55 0.189894
R124 VN.n92 VN.n91 0.189894
R125 VN.n91 VN.n57 0.189894
R126 VN.n87 VN.n57 0.189894
R127 VN.n87 VN.n86 0.189894
R128 VN.n86 VN.n85 0.189894
R129 VN.n85 VN.n59 0.189894
R130 VN.n81 VN.n59 0.189894
R131 VN.n81 VN.n80 0.189894
R132 VN.n80 VN.n79 0.189894
R133 VN.n79 VN.n61 0.189894
R134 VN.n75 VN.n61 0.189894
R135 VN.n75 VN.n74 0.189894
R136 VN.n74 VN.n73 0.189894
R137 VN.n73 VN.n64 0.189894
R138 VN.n69 VN.n64 0.189894
R139 VN.n69 VN.n68 0.189894
R140 VN.n16 VN.n15 0.189894
R141 VN.n16 VN.n11 0.189894
R142 VN.n20 VN.n11 0.189894
R143 VN.n21 VN.n20 0.189894
R144 VN.n22 VN.n21 0.189894
R145 VN.n22 VN.n9 0.189894
R146 VN.n27 VN.n9 0.189894
R147 VN.n28 VN.n27 0.189894
R148 VN.n29 VN.n28 0.189894
R149 VN.n29 VN.n7 0.189894
R150 VN.n33 VN.n7 0.189894
R151 VN.n34 VN.n33 0.189894
R152 VN.n35 VN.n34 0.189894
R153 VN.n35 VN.n5 0.189894
R154 VN.n39 VN.n5 0.189894
R155 VN.n40 VN.n39 0.189894
R156 VN.n40 VN.n3 0.189894
R157 VN.n44 VN.n3 0.189894
R158 VN.n45 VN.n44 0.189894
R159 VN.n46 VN.n45 0.189894
R160 VN.n46 VN.n1 0.189894
R161 VN.n50 VN.n1 0.189894
R162 VTAIL.n11 VTAIL.t12 54.7616
R163 VTAIL.n17 VTAIL.t10 54.7613
R164 VTAIL.n2 VTAIL.t1 54.7613
R165 VTAIL.n16 VTAIL.t2 54.7613
R166 VTAIL.n15 VTAIL.n14 52.9477
R167 VTAIL.n13 VTAIL.n12 52.9477
R168 VTAIL.n10 VTAIL.n9 52.9477
R169 VTAIL.n8 VTAIL.n7 52.9477
R170 VTAIL.n19 VTAIL.n18 52.9474
R171 VTAIL.n1 VTAIL.n0 52.9474
R172 VTAIL.n4 VTAIL.n3 52.9474
R173 VTAIL.n6 VTAIL.n5 52.9474
R174 VTAIL.n8 VTAIL.n6 34.3152
R175 VTAIL.n17 VTAIL.n16 31.0652
R176 VTAIL.n10 VTAIL.n8 3.2505
R177 VTAIL.n11 VTAIL.n10 3.2505
R178 VTAIL.n15 VTAIL.n13 3.2505
R179 VTAIL.n16 VTAIL.n15 3.2505
R180 VTAIL.n6 VTAIL.n4 3.2505
R181 VTAIL.n4 VTAIL.n2 3.2505
R182 VTAIL.n19 VTAIL.n17 3.2505
R183 VTAIL VTAIL.n1 2.49619
R184 VTAIL.n13 VTAIL.n11 2.09533
R185 VTAIL.n2 VTAIL.n1 2.09533
R186 VTAIL.n18 VTAIL.t13 1.8144
R187 VTAIL.n18 VTAIL.t17 1.8144
R188 VTAIL.n0 VTAIL.t14 1.8144
R189 VTAIL.n0 VTAIL.t16 1.8144
R190 VTAIL.n3 VTAIL.t7 1.8144
R191 VTAIL.n3 VTAIL.t6 1.8144
R192 VTAIL.n5 VTAIL.t4 1.8144
R193 VTAIL.n5 VTAIL.t3 1.8144
R194 VTAIL.n14 VTAIL.t0 1.8144
R195 VTAIL.n14 VTAIL.t8 1.8144
R196 VTAIL.n12 VTAIL.t9 1.8144
R197 VTAIL.n12 VTAIL.t5 1.8144
R198 VTAIL.n9 VTAIL.t11 1.8144
R199 VTAIL.n9 VTAIL.t19 1.8144
R200 VTAIL.n7 VTAIL.t15 1.8144
R201 VTAIL.n7 VTAIL.t18 1.8144
R202 VTAIL VTAIL.n19 0.75481
R203 VDD2.n1 VDD2.t9 74.6901
R204 VDD2.n3 VDD2.n2 72.0084
R205 VDD2 VDD2.n7 72.0056
R206 VDD2.n4 VDD2.t1 71.4403
R207 VDD2.n6 VDD2.n5 69.6265
R208 VDD2.n1 VDD2.n0 69.6262
R209 VDD2.n4 VDD2.n3 54.6011
R210 VDD2.n6 VDD2.n4 3.2505
R211 VDD2.n7 VDD2.t4 1.8144
R212 VDD2.n7 VDD2.t8 1.8144
R213 VDD2.n5 VDD2.t3 1.8144
R214 VDD2.n5 VDD2.t7 1.8144
R215 VDD2.n2 VDD2.t6 1.8144
R216 VDD2.n2 VDD2.t2 1.8144
R217 VDD2.n0 VDD2.t5 1.8144
R218 VDD2.n0 VDD2.t0 1.8144
R219 VDD2 VDD2.n6 0.87119
R220 VDD2.n3 VDD2.n1 0.757654
R221 VP.n32 VP.n29 161.3
R222 VP.n34 VP.n33 161.3
R223 VP.n35 VP.n28 161.3
R224 VP.n37 VP.n36 161.3
R225 VP.n38 VP.n27 161.3
R226 VP.n40 VP.n39 161.3
R227 VP.n41 VP.n26 161.3
R228 VP.n44 VP.n43 161.3
R229 VP.n45 VP.n25 161.3
R230 VP.n47 VP.n46 161.3
R231 VP.n48 VP.n24 161.3
R232 VP.n50 VP.n49 161.3
R233 VP.n51 VP.n23 161.3
R234 VP.n53 VP.n52 161.3
R235 VP.n54 VP.n22 161.3
R236 VP.n56 VP.n55 161.3
R237 VP.n58 VP.n57 161.3
R238 VP.n59 VP.n20 161.3
R239 VP.n61 VP.n60 161.3
R240 VP.n62 VP.n19 161.3
R241 VP.n64 VP.n63 161.3
R242 VP.n65 VP.n18 161.3
R243 VP.n67 VP.n66 161.3
R244 VP.n117 VP.n116 161.3
R245 VP.n115 VP.n1 161.3
R246 VP.n114 VP.n113 161.3
R247 VP.n112 VP.n2 161.3
R248 VP.n111 VP.n110 161.3
R249 VP.n109 VP.n3 161.3
R250 VP.n108 VP.n107 161.3
R251 VP.n106 VP.n105 161.3
R252 VP.n104 VP.n5 161.3
R253 VP.n103 VP.n102 161.3
R254 VP.n101 VP.n6 161.3
R255 VP.n100 VP.n99 161.3
R256 VP.n98 VP.n7 161.3
R257 VP.n97 VP.n96 161.3
R258 VP.n95 VP.n8 161.3
R259 VP.n94 VP.n93 161.3
R260 VP.n91 VP.n9 161.3
R261 VP.n90 VP.n89 161.3
R262 VP.n88 VP.n10 161.3
R263 VP.n87 VP.n86 161.3
R264 VP.n85 VP.n11 161.3
R265 VP.n84 VP.n83 161.3
R266 VP.n82 VP.n12 161.3
R267 VP.n81 VP.n80 161.3
R268 VP.n78 VP.n13 161.3
R269 VP.n77 VP.n76 161.3
R270 VP.n75 VP.n14 161.3
R271 VP.n74 VP.n73 161.3
R272 VP.n72 VP.n15 161.3
R273 VP.n71 VP.n70 161.3
R274 VP.n31 VP.t2 158.196
R275 VP.n16 VP.t1 125.544
R276 VP.n79 VP.t4 125.544
R277 VP.n92 VP.t0 125.544
R278 VP.n4 VP.t3 125.544
R279 VP.n0 VP.t5 125.544
R280 VP.n17 VP.t6 125.544
R281 VP.n21 VP.t9 125.544
R282 VP.n42 VP.t8 125.544
R283 VP.n30 VP.t7 125.544
R284 VP.n69 VP.n16 75.7718
R285 VP.n118 VP.n0 75.7718
R286 VP.n68 VP.n17 75.7718
R287 VP.n31 VP.n30 73.5206
R288 VP.n69 VP.n68 62.3059
R289 VP.n86 VP.n10 53.5561
R290 VP.n99 VP.n6 53.5561
R291 VP.n49 VP.n23 53.5561
R292 VP.n36 VP.n27 53.5561
R293 VP.n77 VP.n14 49.6611
R294 VP.n110 VP.n2 49.6611
R295 VP.n60 VP.n19 49.6611
R296 VP.n73 VP.n14 31.1601
R297 VP.n114 VP.n2 31.1601
R298 VP.n64 VP.n19 31.1601
R299 VP.n90 VP.n10 27.2651
R300 VP.n99 VP.n98 27.2651
R301 VP.n49 VP.n48 27.2651
R302 VP.n40 VP.n27 27.2651
R303 VP.n72 VP.n71 24.3439
R304 VP.n73 VP.n72 24.3439
R305 VP.n78 VP.n77 24.3439
R306 VP.n80 VP.n78 24.3439
R307 VP.n84 VP.n12 24.3439
R308 VP.n85 VP.n84 24.3439
R309 VP.n86 VP.n85 24.3439
R310 VP.n91 VP.n90 24.3439
R311 VP.n93 VP.n91 24.3439
R312 VP.n97 VP.n8 24.3439
R313 VP.n98 VP.n97 24.3439
R314 VP.n103 VP.n6 24.3439
R315 VP.n104 VP.n103 24.3439
R316 VP.n105 VP.n104 24.3439
R317 VP.n109 VP.n108 24.3439
R318 VP.n110 VP.n109 24.3439
R319 VP.n115 VP.n114 24.3439
R320 VP.n116 VP.n115 24.3439
R321 VP.n65 VP.n64 24.3439
R322 VP.n66 VP.n65 24.3439
R323 VP.n53 VP.n23 24.3439
R324 VP.n54 VP.n53 24.3439
R325 VP.n55 VP.n54 24.3439
R326 VP.n59 VP.n58 24.3439
R327 VP.n60 VP.n59 24.3439
R328 VP.n41 VP.n40 24.3439
R329 VP.n43 VP.n41 24.3439
R330 VP.n47 VP.n25 24.3439
R331 VP.n48 VP.n47 24.3439
R332 VP.n34 VP.n29 24.3439
R333 VP.n35 VP.n34 24.3439
R334 VP.n36 VP.n35 24.3439
R335 VP.n80 VP.n79 23.3702
R336 VP.n108 VP.n4 23.3702
R337 VP.n58 VP.n21 23.3702
R338 VP.n71 VP.n16 14.1197
R339 VP.n116 VP.n0 14.1197
R340 VP.n66 VP.n17 14.1197
R341 VP.n93 VP.n92 12.1722
R342 VP.n92 VP.n8 12.1722
R343 VP.n43 VP.n42 12.1722
R344 VP.n42 VP.n25 12.1722
R345 VP.n32 VP.n31 4.21321
R346 VP.n79 VP.n12 0.974237
R347 VP.n105 VP.n4 0.974237
R348 VP.n55 VP.n21 0.974237
R349 VP.n30 VP.n29 0.974237
R350 VP.n68 VP.n67 0.355081
R351 VP.n70 VP.n69 0.355081
R352 VP.n118 VP.n117 0.355081
R353 VP VP.n118 0.26685
R354 VP.n33 VP.n32 0.189894
R355 VP.n33 VP.n28 0.189894
R356 VP.n37 VP.n28 0.189894
R357 VP.n38 VP.n37 0.189894
R358 VP.n39 VP.n38 0.189894
R359 VP.n39 VP.n26 0.189894
R360 VP.n44 VP.n26 0.189894
R361 VP.n45 VP.n44 0.189894
R362 VP.n46 VP.n45 0.189894
R363 VP.n46 VP.n24 0.189894
R364 VP.n50 VP.n24 0.189894
R365 VP.n51 VP.n50 0.189894
R366 VP.n52 VP.n51 0.189894
R367 VP.n52 VP.n22 0.189894
R368 VP.n56 VP.n22 0.189894
R369 VP.n57 VP.n56 0.189894
R370 VP.n57 VP.n20 0.189894
R371 VP.n61 VP.n20 0.189894
R372 VP.n62 VP.n61 0.189894
R373 VP.n63 VP.n62 0.189894
R374 VP.n63 VP.n18 0.189894
R375 VP.n67 VP.n18 0.189894
R376 VP.n70 VP.n15 0.189894
R377 VP.n74 VP.n15 0.189894
R378 VP.n75 VP.n74 0.189894
R379 VP.n76 VP.n75 0.189894
R380 VP.n76 VP.n13 0.189894
R381 VP.n81 VP.n13 0.189894
R382 VP.n82 VP.n81 0.189894
R383 VP.n83 VP.n82 0.189894
R384 VP.n83 VP.n11 0.189894
R385 VP.n87 VP.n11 0.189894
R386 VP.n88 VP.n87 0.189894
R387 VP.n89 VP.n88 0.189894
R388 VP.n89 VP.n9 0.189894
R389 VP.n94 VP.n9 0.189894
R390 VP.n95 VP.n94 0.189894
R391 VP.n96 VP.n95 0.189894
R392 VP.n96 VP.n7 0.189894
R393 VP.n100 VP.n7 0.189894
R394 VP.n101 VP.n100 0.189894
R395 VP.n102 VP.n101 0.189894
R396 VP.n102 VP.n5 0.189894
R397 VP.n106 VP.n5 0.189894
R398 VP.n107 VP.n106 0.189894
R399 VP.n107 VP.n3 0.189894
R400 VP.n111 VP.n3 0.189894
R401 VP.n112 VP.n111 0.189894
R402 VP.n113 VP.n112 0.189894
R403 VP.n113 VP.n1 0.189894
R404 VP.n117 VP.n1 0.189894
R405 VDD1.n1 VDD1.t7 74.6903
R406 VDD1.n3 VDD1.t8 74.6901
R407 VDD1.n5 VDD1.n4 72.0084
R408 VDD1.n1 VDD1.n0 69.6265
R409 VDD1.n7 VDD1.n6 69.6262
R410 VDD1.n3 VDD1.n2 69.6262
R411 VDD1.n7 VDD1.n5 56.8091
R412 VDD1 VDD1.n7 2.37981
R413 VDD1.n6 VDD1.t0 1.8144
R414 VDD1.n6 VDD1.t3 1.8144
R415 VDD1.n0 VDD1.t2 1.8144
R416 VDD1.n0 VDD1.t1 1.8144
R417 VDD1.n4 VDD1.t6 1.8144
R418 VDD1.n4 VDD1.t4 1.8144
R419 VDD1.n2 VDD1.t5 1.8144
R420 VDD1.n2 VDD1.t9 1.8144
R421 VDD1 VDD1.n1 0.87119
R422 VDD1.n5 VDD1.n3 0.757654
R423 B.n590 B.n183 585
R424 B.n589 B.n588 585
R425 B.n587 B.n184 585
R426 B.n586 B.n585 585
R427 B.n584 B.n185 585
R428 B.n583 B.n582 585
R429 B.n581 B.n186 585
R430 B.n580 B.n579 585
R431 B.n578 B.n187 585
R432 B.n577 B.n576 585
R433 B.n575 B.n188 585
R434 B.n574 B.n573 585
R435 B.n572 B.n189 585
R436 B.n571 B.n570 585
R437 B.n569 B.n190 585
R438 B.n568 B.n567 585
R439 B.n566 B.n191 585
R440 B.n565 B.n564 585
R441 B.n563 B.n192 585
R442 B.n562 B.n561 585
R443 B.n560 B.n193 585
R444 B.n559 B.n558 585
R445 B.n557 B.n194 585
R446 B.n556 B.n555 585
R447 B.n554 B.n195 585
R448 B.n553 B.n552 585
R449 B.n551 B.n196 585
R450 B.n550 B.n549 585
R451 B.n548 B.n197 585
R452 B.n547 B.n546 585
R453 B.n545 B.n198 585
R454 B.n544 B.n543 585
R455 B.n542 B.n199 585
R456 B.n541 B.n540 585
R457 B.n539 B.n200 585
R458 B.n538 B.n537 585
R459 B.n536 B.n201 585
R460 B.n535 B.n534 585
R461 B.n533 B.n202 585
R462 B.n532 B.n531 585
R463 B.n530 B.n203 585
R464 B.n529 B.n528 585
R465 B.n527 B.n204 585
R466 B.n526 B.n525 585
R467 B.n524 B.n205 585
R468 B.n523 B.n522 585
R469 B.n521 B.n206 585
R470 B.n520 B.n519 585
R471 B.n518 B.n207 585
R472 B.n517 B.n516 585
R473 B.n515 B.n208 585
R474 B.n514 B.n513 585
R475 B.n512 B.n209 585
R476 B.n511 B.n510 585
R477 B.n509 B.n210 585
R478 B.n508 B.n507 585
R479 B.n506 B.n211 585
R480 B.n505 B.n504 585
R481 B.n503 B.n212 585
R482 B.n501 B.n500 585
R483 B.n499 B.n215 585
R484 B.n498 B.n497 585
R485 B.n496 B.n216 585
R486 B.n495 B.n494 585
R487 B.n493 B.n217 585
R488 B.n492 B.n491 585
R489 B.n490 B.n218 585
R490 B.n489 B.n488 585
R491 B.n487 B.n219 585
R492 B.n486 B.n485 585
R493 B.n481 B.n220 585
R494 B.n480 B.n479 585
R495 B.n478 B.n221 585
R496 B.n477 B.n476 585
R497 B.n475 B.n222 585
R498 B.n474 B.n473 585
R499 B.n472 B.n223 585
R500 B.n471 B.n470 585
R501 B.n469 B.n224 585
R502 B.n468 B.n467 585
R503 B.n466 B.n225 585
R504 B.n465 B.n464 585
R505 B.n463 B.n226 585
R506 B.n462 B.n461 585
R507 B.n460 B.n227 585
R508 B.n459 B.n458 585
R509 B.n457 B.n228 585
R510 B.n456 B.n455 585
R511 B.n454 B.n229 585
R512 B.n453 B.n452 585
R513 B.n451 B.n230 585
R514 B.n450 B.n449 585
R515 B.n448 B.n231 585
R516 B.n447 B.n446 585
R517 B.n445 B.n232 585
R518 B.n444 B.n443 585
R519 B.n442 B.n233 585
R520 B.n441 B.n440 585
R521 B.n439 B.n234 585
R522 B.n438 B.n437 585
R523 B.n436 B.n235 585
R524 B.n435 B.n434 585
R525 B.n433 B.n236 585
R526 B.n432 B.n431 585
R527 B.n430 B.n237 585
R528 B.n429 B.n428 585
R529 B.n427 B.n238 585
R530 B.n426 B.n425 585
R531 B.n424 B.n239 585
R532 B.n423 B.n422 585
R533 B.n421 B.n240 585
R534 B.n420 B.n419 585
R535 B.n418 B.n241 585
R536 B.n417 B.n416 585
R537 B.n415 B.n242 585
R538 B.n414 B.n413 585
R539 B.n412 B.n243 585
R540 B.n411 B.n410 585
R541 B.n409 B.n244 585
R542 B.n408 B.n407 585
R543 B.n406 B.n245 585
R544 B.n405 B.n404 585
R545 B.n403 B.n246 585
R546 B.n402 B.n401 585
R547 B.n400 B.n247 585
R548 B.n399 B.n398 585
R549 B.n397 B.n248 585
R550 B.n396 B.n395 585
R551 B.n592 B.n591 585
R552 B.n593 B.n182 585
R553 B.n595 B.n594 585
R554 B.n596 B.n181 585
R555 B.n598 B.n597 585
R556 B.n599 B.n180 585
R557 B.n601 B.n600 585
R558 B.n602 B.n179 585
R559 B.n604 B.n603 585
R560 B.n605 B.n178 585
R561 B.n607 B.n606 585
R562 B.n608 B.n177 585
R563 B.n610 B.n609 585
R564 B.n611 B.n176 585
R565 B.n613 B.n612 585
R566 B.n614 B.n175 585
R567 B.n616 B.n615 585
R568 B.n617 B.n174 585
R569 B.n619 B.n618 585
R570 B.n620 B.n173 585
R571 B.n622 B.n621 585
R572 B.n623 B.n172 585
R573 B.n625 B.n624 585
R574 B.n626 B.n171 585
R575 B.n628 B.n627 585
R576 B.n629 B.n170 585
R577 B.n631 B.n630 585
R578 B.n632 B.n169 585
R579 B.n634 B.n633 585
R580 B.n635 B.n168 585
R581 B.n637 B.n636 585
R582 B.n638 B.n167 585
R583 B.n640 B.n639 585
R584 B.n641 B.n166 585
R585 B.n643 B.n642 585
R586 B.n644 B.n165 585
R587 B.n646 B.n645 585
R588 B.n647 B.n164 585
R589 B.n649 B.n648 585
R590 B.n650 B.n163 585
R591 B.n652 B.n651 585
R592 B.n653 B.n162 585
R593 B.n655 B.n654 585
R594 B.n656 B.n161 585
R595 B.n658 B.n657 585
R596 B.n659 B.n160 585
R597 B.n661 B.n660 585
R598 B.n662 B.n159 585
R599 B.n664 B.n663 585
R600 B.n665 B.n158 585
R601 B.n667 B.n666 585
R602 B.n668 B.n157 585
R603 B.n670 B.n669 585
R604 B.n671 B.n156 585
R605 B.n673 B.n672 585
R606 B.n674 B.n155 585
R607 B.n676 B.n675 585
R608 B.n677 B.n154 585
R609 B.n679 B.n678 585
R610 B.n680 B.n153 585
R611 B.n682 B.n681 585
R612 B.n683 B.n152 585
R613 B.n685 B.n684 585
R614 B.n686 B.n151 585
R615 B.n688 B.n687 585
R616 B.n689 B.n150 585
R617 B.n691 B.n690 585
R618 B.n692 B.n149 585
R619 B.n694 B.n693 585
R620 B.n695 B.n148 585
R621 B.n697 B.n696 585
R622 B.n698 B.n147 585
R623 B.n700 B.n699 585
R624 B.n701 B.n146 585
R625 B.n703 B.n702 585
R626 B.n704 B.n145 585
R627 B.n706 B.n705 585
R628 B.n707 B.n144 585
R629 B.n709 B.n708 585
R630 B.n710 B.n143 585
R631 B.n712 B.n711 585
R632 B.n713 B.n142 585
R633 B.n715 B.n714 585
R634 B.n716 B.n141 585
R635 B.n718 B.n717 585
R636 B.n719 B.n140 585
R637 B.n721 B.n720 585
R638 B.n722 B.n139 585
R639 B.n724 B.n723 585
R640 B.n725 B.n138 585
R641 B.n727 B.n726 585
R642 B.n728 B.n137 585
R643 B.n730 B.n729 585
R644 B.n731 B.n136 585
R645 B.n733 B.n732 585
R646 B.n734 B.n135 585
R647 B.n736 B.n735 585
R648 B.n737 B.n134 585
R649 B.n739 B.n738 585
R650 B.n740 B.n133 585
R651 B.n742 B.n741 585
R652 B.n743 B.n132 585
R653 B.n745 B.n744 585
R654 B.n746 B.n131 585
R655 B.n748 B.n747 585
R656 B.n749 B.n130 585
R657 B.n751 B.n750 585
R658 B.n752 B.n129 585
R659 B.n754 B.n753 585
R660 B.n755 B.n128 585
R661 B.n757 B.n756 585
R662 B.n758 B.n127 585
R663 B.n760 B.n759 585
R664 B.n761 B.n126 585
R665 B.n763 B.n762 585
R666 B.n764 B.n125 585
R667 B.n766 B.n765 585
R668 B.n767 B.n124 585
R669 B.n769 B.n768 585
R670 B.n770 B.n123 585
R671 B.n772 B.n771 585
R672 B.n773 B.n122 585
R673 B.n775 B.n774 585
R674 B.n776 B.n121 585
R675 B.n778 B.n777 585
R676 B.n779 B.n120 585
R677 B.n781 B.n780 585
R678 B.n782 B.n119 585
R679 B.n784 B.n783 585
R680 B.n785 B.n118 585
R681 B.n787 B.n786 585
R682 B.n788 B.n117 585
R683 B.n790 B.n789 585
R684 B.n791 B.n116 585
R685 B.n793 B.n792 585
R686 B.n794 B.n115 585
R687 B.n796 B.n795 585
R688 B.n797 B.n114 585
R689 B.n799 B.n798 585
R690 B.n800 B.n113 585
R691 B.n802 B.n801 585
R692 B.n803 B.n112 585
R693 B.n805 B.n804 585
R694 B.n806 B.n111 585
R695 B.n808 B.n807 585
R696 B.n809 B.n110 585
R697 B.n811 B.n810 585
R698 B.n812 B.n109 585
R699 B.n814 B.n813 585
R700 B.n815 B.n108 585
R701 B.n1008 B.n39 585
R702 B.n1007 B.n1006 585
R703 B.n1005 B.n40 585
R704 B.n1004 B.n1003 585
R705 B.n1002 B.n41 585
R706 B.n1001 B.n1000 585
R707 B.n999 B.n42 585
R708 B.n998 B.n997 585
R709 B.n996 B.n43 585
R710 B.n995 B.n994 585
R711 B.n993 B.n44 585
R712 B.n992 B.n991 585
R713 B.n990 B.n45 585
R714 B.n989 B.n988 585
R715 B.n987 B.n46 585
R716 B.n986 B.n985 585
R717 B.n984 B.n47 585
R718 B.n983 B.n982 585
R719 B.n981 B.n48 585
R720 B.n980 B.n979 585
R721 B.n978 B.n49 585
R722 B.n977 B.n976 585
R723 B.n975 B.n50 585
R724 B.n974 B.n973 585
R725 B.n972 B.n51 585
R726 B.n971 B.n970 585
R727 B.n969 B.n52 585
R728 B.n968 B.n967 585
R729 B.n966 B.n53 585
R730 B.n965 B.n964 585
R731 B.n963 B.n54 585
R732 B.n962 B.n961 585
R733 B.n960 B.n55 585
R734 B.n959 B.n958 585
R735 B.n957 B.n56 585
R736 B.n956 B.n955 585
R737 B.n954 B.n57 585
R738 B.n953 B.n952 585
R739 B.n951 B.n58 585
R740 B.n950 B.n949 585
R741 B.n948 B.n59 585
R742 B.n947 B.n946 585
R743 B.n945 B.n60 585
R744 B.n944 B.n943 585
R745 B.n942 B.n61 585
R746 B.n941 B.n940 585
R747 B.n939 B.n62 585
R748 B.n938 B.n937 585
R749 B.n936 B.n63 585
R750 B.n935 B.n934 585
R751 B.n933 B.n64 585
R752 B.n932 B.n931 585
R753 B.n930 B.n65 585
R754 B.n929 B.n928 585
R755 B.n927 B.n66 585
R756 B.n926 B.n925 585
R757 B.n924 B.n67 585
R758 B.n923 B.n922 585
R759 B.n921 B.n68 585
R760 B.n920 B.n919 585
R761 B.n918 B.n69 585
R762 B.n917 B.n916 585
R763 B.n915 B.n73 585
R764 B.n914 B.n913 585
R765 B.n912 B.n74 585
R766 B.n911 B.n910 585
R767 B.n909 B.n75 585
R768 B.n908 B.n907 585
R769 B.n906 B.n76 585
R770 B.n904 B.n903 585
R771 B.n902 B.n79 585
R772 B.n901 B.n900 585
R773 B.n899 B.n80 585
R774 B.n898 B.n897 585
R775 B.n896 B.n81 585
R776 B.n895 B.n894 585
R777 B.n893 B.n82 585
R778 B.n892 B.n891 585
R779 B.n890 B.n83 585
R780 B.n889 B.n888 585
R781 B.n887 B.n84 585
R782 B.n886 B.n885 585
R783 B.n884 B.n85 585
R784 B.n883 B.n882 585
R785 B.n881 B.n86 585
R786 B.n880 B.n879 585
R787 B.n878 B.n87 585
R788 B.n877 B.n876 585
R789 B.n875 B.n88 585
R790 B.n874 B.n873 585
R791 B.n872 B.n89 585
R792 B.n871 B.n870 585
R793 B.n869 B.n90 585
R794 B.n868 B.n867 585
R795 B.n866 B.n91 585
R796 B.n865 B.n864 585
R797 B.n863 B.n92 585
R798 B.n862 B.n861 585
R799 B.n860 B.n93 585
R800 B.n859 B.n858 585
R801 B.n857 B.n94 585
R802 B.n856 B.n855 585
R803 B.n854 B.n95 585
R804 B.n853 B.n852 585
R805 B.n851 B.n96 585
R806 B.n850 B.n849 585
R807 B.n848 B.n97 585
R808 B.n847 B.n846 585
R809 B.n845 B.n98 585
R810 B.n844 B.n843 585
R811 B.n842 B.n99 585
R812 B.n841 B.n840 585
R813 B.n839 B.n100 585
R814 B.n838 B.n837 585
R815 B.n836 B.n101 585
R816 B.n835 B.n834 585
R817 B.n833 B.n102 585
R818 B.n832 B.n831 585
R819 B.n830 B.n103 585
R820 B.n829 B.n828 585
R821 B.n827 B.n104 585
R822 B.n826 B.n825 585
R823 B.n824 B.n105 585
R824 B.n823 B.n822 585
R825 B.n821 B.n106 585
R826 B.n820 B.n819 585
R827 B.n818 B.n107 585
R828 B.n817 B.n816 585
R829 B.n1010 B.n1009 585
R830 B.n1011 B.n38 585
R831 B.n1013 B.n1012 585
R832 B.n1014 B.n37 585
R833 B.n1016 B.n1015 585
R834 B.n1017 B.n36 585
R835 B.n1019 B.n1018 585
R836 B.n1020 B.n35 585
R837 B.n1022 B.n1021 585
R838 B.n1023 B.n34 585
R839 B.n1025 B.n1024 585
R840 B.n1026 B.n33 585
R841 B.n1028 B.n1027 585
R842 B.n1029 B.n32 585
R843 B.n1031 B.n1030 585
R844 B.n1032 B.n31 585
R845 B.n1034 B.n1033 585
R846 B.n1035 B.n30 585
R847 B.n1037 B.n1036 585
R848 B.n1038 B.n29 585
R849 B.n1040 B.n1039 585
R850 B.n1041 B.n28 585
R851 B.n1043 B.n1042 585
R852 B.n1044 B.n27 585
R853 B.n1046 B.n1045 585
R854 B.n1047 B.n26 585
R855 B.n1049 B.n1048 585
R856 B.n1050 B.n25 585
R857 B.n1052 B.n1051 585
R858 B.n1053 B.n24 585
R859 B.n1055 B.n1054 585
R860 B.n1056 B.n23 585
R861 B.n1058 B.n1057 585
R862 B.n1059 B.n22 585
R863 B.n1061 B.n1060 585
R864 B.n1062 B.n21 585
R865 B.n1064 B.n1063 585
R866 B.n1065 B.n20 585
R867 B.n1067 B.n1066 585
R868 B.n1068 B.n19 585
R869 B.n1070 B.n1069 585
R870 B.n1071 B.n18 585
R871 B.n1073 B.n1072 585
R872 B.n1074 B.n17 585
R873 B.n1076 B.n1075 585
R874 B.n1077 B.n16 585
R875 B.n1079 B.n1078 585
R876 B.n1080 B.n15 585
R877 B.n1082 B.n1081 585
R878 B.n1083 B.n14 585
R879 B.n1085 B.n1084 585
R880 B.n1086 B.n13 585
R881 B.n1088 B.n1087 585
R882 B.n1089 B.n12 585
R883 B.n1091 B.n1090 585
R884 B.n1092 B.n11 585
R885 B.n1094 B.n1093 585
R886 B.n1095 B.n10 585
R887 B.n1097 B.n1096 585
R888 B.n1098 B.n9 585
R889 B.n1100 B.n1099 585
R890 B.n1101 B.n8 585
R891 B.n1103 B.n1102 585
R892 B.n1104 B.n7 585
R893 B.n1106 B.n1105 585
R894 B.n1107 B.n6 585
R895 B.n1109 B.n1108 585
R896 B.n1110 B.n5 585
R897 B.n1112 B.n1111 585
R898 B.n1113 B.n4 585
R899 B.n1115 B.n1114 585
R900 B.n1116 B.n3 585
R901 B.n1118 B.n1117 585
R902 B.n1119 B.n0 585
R903 B.n2 B.n1 585
R904 B.n286 B.n285 585
R905 B.n288 B.n287 585
R906 B.n289 B.n284 585
R907 B.n291 B.n290 585
R908 B.n292 B.n283 585
R909 B.n294 B.n293 585
R910 B.n295 B.n282 585
R911 B.n297 B.n296 585
R912 B.n298 B.n281 585
R913 B.n300 B.n299 585
R914 B.n301 B.n280 585
R915 B.n303 B.n302 585
R916 B.n304 B.n279 585
R917 B.n306 B.n305 585
R918 B.n307 B.n278 585
R919 B.n309 B.n308 585
R920 B.n310 B.n277 585
R921 B.n312 B.n311 585
R922 B.n313 B.n276 585
R923 B.n315 B.n314 585
R924 B.n316 B.n275 585
R925 B.n318 B.n317 585
R926 B.n319 B.n274 585
R927 B.n321 B.n320 585
R928 B.n322 B.n273 585
R929 B.n324 B.n323 585
R930 B.n325 B.n272 585
R931 B.n327 B.n326 585
R932 B.n328 B.n271 585
R933 B.n330 B.n329 585
R934 B.n331 B.n270 585
R935 B.n333 B.n332 585
R936 B.n334 B.n269 585
R937 B.n336 B.n335 585
R938 B.n337 B.n268 585
R939 B.n339 B.n338 585
R940 B.n340 B.n267 585
R941 B.n342 B.n341 585
R942 B.n343 B.n266 585
R943 B.n345 B.n344 585
R944 B.n346 B.n265 585
R945 B.n348 B.n347 585
R946 B.n349 B.n264 585
R947 B.n351 B.n350 585
R948 B.n352 B.n263 585
R949 B.n354 B.n353 585
R950 B.n355 B.n262 585
R951 B.n357 B.n356 585
R952 B.n358 B.n261 585
R953 B.n360 B.n359 585
R954 B.n361 B.n260 585
R955 B.n363 B.n362 585
R956 B.n364 B.n259 585
R957 B.n366 B.n365 585
R958 B.n367 B.n258 585
R959 B.n369 B.n368 585
R960 B.n370 B.n257 585
R961 B.n372 B.n371 585
R962 B.n373 B.n256 585
R963 B.n375 B.n374 585
R964 B.n376 B.n255 585
R965 B.n378 B.n377 585
R966 B.n379 B.n254 585
R967 B.n381 B.n380 585
R968 B.n382 B.n253 585
R969 B.n384 B.n383 585
R970 B.n385 B.n252 585
R971 B.n387 B.n386 585
R972 B.n388 B.n251 585
R973 B.n390 B.n389 585
R974 B.n391 B.n250 585
R975 B.n393 B.n392 585
R976 B.n394 B.n249 585
R977 B.n395 B.n394 492.5
R978 B.n591 B.n590 492.5
R979 B.n817 B.n108 492.5
R980 B.n1010 B.n39 492.5
R981 B.n482 B.t9 334.584
R982 B.n213 B.t3 334.584
R983 B.n77 B.t0 334.584
R984 B.n70 B.t6 334.584
R985 B.n1121 B.n1120 256.663
R986 B.n1120 B.n1119 235.042
R987 B.n1120 B.n2 235.042
R988 B.n213 B.t4 183.982
R989 B.n77 B.t2 183.982
R990 B.n482 B.t10 183.958
R991 B.n70 B.t8 183.958
R992 B.n395 B.n248 163.367
R993 B.n399 B.n248 163.367
R994 B.n400 B.n399 163.367
R995 B.n401 B.n400 163.367
R996 B.n401 B.n246 163.367
R997 B.n405 B.n246 163.367
R998 B.n406 B.n405 163.367
R999 B.n407 B.n406 163.367
R1000 B.n407 B.n244 163.367
R1001 B.n411 B.n244 163.367
R1002 B.n412 B.n411 163.367
R1003 B.n413 B.n412 163.367
R1004 B.n413 B.n242 163.367
R1005 B.n417 B.n242 163.367
R1006 B.n418 B.n417 163.367
R1007 B.n419 B.n418 163.367
R1008 B.n419 B.n240 163.367
R1009 B.n423 B.n240 163.367
R1010 B.n424 B.n423 163.367
R1011 B.n425 B.n424 163.367
R1012 B.n425 B.n238 163.367
R1013 B.n429 B.n238 163.367
R1014 B.n430 B.n429 163.367
R1015 B.n431 B.n430 163.367
R1016 B.n431 B.n236 163.367
R1017 B.n435 B.n236 163.367
R1018 B.n436 B.n435 163.367
R1019 B.n437 B.n436 163.367
R1020 B.n437 B.n234 163.367
R1021 B.n441 B.n234 163.367
R1022 B.n442 B.n441 163.367
R1023 B.n443 B.n442 163.367
R1024 B.n443 B.n232 163.367
R1025 B.n447 B.n232 163.367
R1026 B.n448 B.n447 163.367
R1027 B.n449 B.n448 163.367
R1028 B.n449 B.n230 163.367
R1029 B.n453 B.n230 163.367
R1030 B.n454 B.n453 163.367
R1031 B.n455 B.n454 163.367
R1032 B.n455 B.n228 163.367
R1033 B.n459 B.n228 163.367
R1034 B.n460 B.n459 163.367
R1035 B.n461 B.n460 163.367
R1036 B.n461 B.n226 163.367
R1037 B.n465 B.n226 163.367
R1038 B.n466 B.n465 163.367
R1039 B.n467 B.n466 163.367
R1040 B.n467 B.n224 163.367
R1041 B.n471 B.n224 163.367
R1042 B.n472 B.n471 163.367
R1043 B.n473 B.n472 163.367
R1044 B.n473 B.n222 163.367
R1045 B.n477 B.n222 163.367
R1046 B.n478 B.n477 163.367
R1047 B.n479 B.n478 163.367
R1048 B.n479 B.n220 163.367
R1049 B.n486 B.n220 163.367
R1050 B.n487 B.n486 163.367
R1051 B.n488 B.n487 163.367
R1052 B.n488 B.n218 163.367
R1053 B.n492 B.n218 163.367
R1054 B.n493 B.n492 163.367
R1055 B.n494 B.n493 163.367
R1056 B.n494 B.n216 163.367
R1057 B.n498 B.n216 163.367
R1058 B.n499 B.n498 163.367
R1059 B.n500 B.n499 163.367
R1060 B.n500 B.n212 163.367
R1061 B.n505 B.n212 163.367
R1062 B.n506 B.n505 163.367
R1063 B.n507 B.n506 163.367
R1064 B.n507 B.n210 163.367
R1065 B.n511 B.n210 163.367
R1066 B.n512 B.n511 163.367
R1067 B.n513 B.n512 163.367
R1068 B.n513 B.n208 163.367
R1069 B.n517 B.n208 163.367
R1070 B.n518 B.n517 163.367
R1071 B.n519 B.n518 163.367
R1072 B.n519 B.n206 163.367
R1073 B.n523 B.n206 163.367
R1074 B.n524 B.n523 163.367
R1075 B.n525 B.n524 163.367
R1076 B.n525 B.n204 163.367
R1077 B.n529 B.n204 163.367
R1078 B.n530 B.n529 163.367
R1079 B.n531 B.n530 163.367
R1080 B.n531 B.n202 163.367
R1081 B.n535 B.n202 163.367
R1082 B.n536 B.n535 163.367
R1083 B.n537 B.n536 163.367
R1084 B.n537 B.n200 163.367
R1085 B.n541 B.n200 163.367
R1086 B.n542 B.n541 163.367
R1087 B.n543 B.n542 163.367
R1088 B.n543 B.n198 163.367
R1089 B.n547 B.n198 163.367
R1090 B.n548 B.n547 163.367
R1091 B.n549 B.n548 163.367
R1092 B.n549 B.n196 163.367
R1093 B.n553 B.n196 163.367
R1094 B.n554 B.n553 163.367
R1095 B.n555 B.n554 163.367
R1096 B.n555 B.n194 163.367
R1097 B.n559 B.n194 163.367
R1098 B.n560 B.n559 163.367
R1099 B.n561 B.n560 163.367
R1100 B.n561 B.n192 163.367
R1101 B.n565 B.n192 163.367
R1102 B.n566 B.n565 163.367
R1103 B.n567 B.n566 163.367
R1104 B.n567 B.n190 163.367
R1105 B.n571 B.n190 163.367
R1106 B.n572 B.n571 163.367
R1107 B.n573 B.n572 163.367
R1108 B.n573 B.n188 163.367
R1109 B.n577 B.n188 163.367
R1110 B.n578 B.n577 163.367
R1111 B.n579 B.n578 163.367
R1112 B.n579 B.n186 163.367
R1113 B.n583 B.n186 163.367
R1114 B.n584 B.n583 163.367
R1115 B.n585 B.n584 163.367
R1116 B.n585 B.n184 163.367
R1117 B.n589 B.n184 163.367
R1118 B.n590 B.n589 163.367
R1119 B.n813 B.n108 163.367
R1120 B.n813 B.n812 163.367
R1121 B.n812 B.n811 163.367
R1122 B.n811 B.n110 163.367
R1123 B.n807 B.n110 163.367
R1124 B.n807 B.n806 163.367
R1125 B.n806 B.n805 163.367
R1126 B.n805 B.n112 163.367
R1127 B.n801 B.n112 163.367
R1128 B.n801 B.n800 163.367
R1129 B.n800 B.n799 163.367
R1130 B.n799 B.n114 163.367
R1131 B.n795 B.n114 163.367
R1132 B.n795 B.n794 163.367
R1133 B.n794 B.n793 163.367
R1134 B.n793 B.n116 163.367
R1135 B.n789 B.n116 163.367
R1136 B.n789 B.n788 163.367
R1137 B.n788 B.n787 163.367
R1138 B.n787 B.n118 163.367
R1139 B.n783 B.n118 163.367
R1140 B.n783 B.n782 163.367
R1141 B.n782 B.n781 163.367
R1142 B.n781 B.n120 163.367
R1143 B.n777 B.n120 163.367
R1144 B.n777 B.n776 163.367
R1145 B.n776 B.n775 163.367
R1146 B.n775 B.n122 163.367
R1147 B.n771 B.n122 163.367
R1148 B.n771 B.n770 163.367
R1149 B.n770 B.n769 163.367
R1150 B.n769 B.n124 163.367
R1151 B.n765 B.n124 163.367
R1152 B.n765 B.n764 163.367
R1153 B.n764 B.n763 163.367
R1154 B.n763 B.n126 163.367
R1155 B.n759 B.n126 163.367
R1156 B.n759 B.n758 163.367
R1157 B.n758 B.n757 163.367
R1158 B.n757 B.n128 163.367
R1159 B.n753 B.n128 163.367
R1160 B.n753 B.n752 163.367
R1161 B.n752 B.n751 163.367
R1162 B.n751 B.n130 163.367
R1163 B.n747 B.n130 163.367
R1164 B.n747 B.n746 163.367
R1165 B.n746 B.n745 163.367
R1166 B.n745 B.n132 163.367
R1167 B.n741 B.n132 163.367
R1168 B.n741 B.n740 163.367
R1169 B.n740 B.n739 163.367
R1170 B.n739 B.n134 163.367
R1171 B.n735 B.n134 163.367
R1172 B.n735 B.n734 163.367
R1173 B.n734 B.n733 163.367
R1174 B.n733 B.n136 163.367
R1175 B.n729 B.n136 163.367
R1176 B.n729 B.n728 163.367
R1177 B.n728 B.n727 163.367
R1178 B.n727 B.n138 163.367
R1179 B.n723 B.n138 163.367
R1180 B.n723 B.n722 163.367
R1181 B.n722 B.n721 163.367
R1182 B.n721 B.n140 163.367
R1183 B.n717 B.n140 163.367
R1184 B.n717 B.n716 163.367
R1185 B.n716 B.n715 163.367
R1186 B.n715 B.n142 163.367
R1187 B.n711 B.n142 163.367
R1188 B.n711 B.n710 163.367
R1189 B.n710 B.n709 163.367
R1190 B.n709 B.n144 163.367
R1191 B.n705 B.n144 163.367
R1192 B.n705 B.n704 163.367
R1193 B.n704 B.n703 163.367
R1194 B.n703 B.n146 163.367
R1195 B.n699 B.n146 163.367
R1196 B.n699 B.n698 163.367
R1197 B.n698 B.n697 163.367
R1198 B.n697 B.n148 163.367
R1199 B.n693 B.n148 163.367
R1200 B.n693 B.n692 163.367
R1201 B.n692 B.n691 163.367
R1202 B.n691 B.n150 163.367
R1203 B.n687 B.n150 163.367
R1204 B.n687 B.n686 163.367
R1205 B.n686 B.n685 163.367
R1206 B.n685 B.n152 163.367
R1207 B.n681 B.n152 163.367
R1208 B.n681 B.n680 163.367
R1209 B.n680 B.n679 163.367
R1210 B.n679 B.n154 163.367
R1211 B.n675 B.n154 163.367
R1212 B.n675 B.n674 163.367
R1213 B.n674 B.n673 163.367
R1214 B.n673 B.n156 163.367
R1215 B.n669 B.n156 163.367
R1216 B.n669 B.n668 163.367
R1217 B.n668 B.n667 163.367
R1218 B.n667 B.n158 163.367
R1219 B.n663 B.n158 163.367
R1220 B.n663 B.n662 163.367
R1221 B.n662 B.n661 163.367
R1222 B.n661 B.n160 163.367
R1223 B.n657 B.n160 163.367
R1224 B.n657 B.n656 163.367
R1225 B.n656 B.n655 163.367
R1226 B.n655 B.n162 163.367
R1227 B.n651 B.n162 163.367
R1228 B.n651 B.n650 163.367
R1229 B.n650 B.n649 163.367
R1230 B.n649 B.n164 163.367
R1231 B.n645 B.n164 163.367
R1232 B.n645 B.n644 163.367
R1233 B.n644 B.n643 163.367
R1234 B.n643 B.n166 163.367
R1235 B.n639 B.n166 163.367
R1236 B.n639 B.n638 163.367
R1237 B.n638 B.n637 163.367
R1238 B.n637 B.n168 163.367
R1239 B.n633 B.n168 163.367
R1240 B.n633 B.n632 163.367
R1241 B.n632 B.n631 163.367
R1242 B.n631 B.n170 163.367
R1243 B.n627 B.n170 163.367
R1244 B.n627 B.n626 163.367
R1245 B.n626 B.n625 163.367
R1246 B.n625 B.n172 163.367
R1247 B.n621 B.n172 163.367
R1248 B.n621 B.n620 163.367
R1249 B.n620 B.n619 163.367
R1250 B.n619 B.n174 163.367
R1251 B.n615 B.n174 163.367
R1252 B.n615 B.n614 163.367
R1253 B.n614 B.n613 163.367
R1254 B.n613 B.n176 163.367
R1255 B.n609 B.n176 163.367
R1256 B.n609 B.n608 163.367
R1257 B.n608 B.n607 163.367
R1258 B.n607 B.n178 163.367
R1259 B.n603 B.n178 163.367
R1260 B.n603 B.n602 163.367
R1261 B.n602 B.n601 163.367
R1262 B.n601 B.n180 163.367
R1263 B.n597 B.n180 163.367
R1264 B.n597 B.n596 163.367
R1265 B.n596 B.n595 163.367
R1266 B.n595 B.n182 163.367
R1267 B.n591 B.n182 163.367
R1268 B.n1006 B.n39 163.367
R1269 B.n1006 B.n1005 163.367
R1270 B.n1005 B.n1004 163.367
R1271 B.n1004 B.n41 163.367
R1272 B.n1000 B.n41 163.367
R1273 B.n1000 B.n999 163.367
R1274 B.n999 B.n998 163.367
R1275 B.n998 B.n43 163.367
R1276 B.n994 B.n43 163.367
R1277 B.n994 B.n993 163.367
R1278 B.n993 B.n992 163.367
R1279 B.n992 B.n45 163.367
R1280 B.n988 B.n45 163.367
R1281 B.n988 B.n987 163.367
R1282 B.n987 B.n986 163.367
R1283 B.n986 B.n47 163.367
R1284 B.n982 B.n47 163.367
R1285 B.n982 B.n981 163.367
R1286 B.n981 B.n980 163.367
R1287 B.n980 B.n49 163.367
R1288 B.n976 B.n49 163.367
R1289 B.n976 B.n975 163.367
R1290 B.n975 B.n974 163.367
R1291 B.n974 B.n51 163.367
R1292 B.n970 B.n51 163.367
R1293 B.n970 B.n969 163.367
R1294 B.n969 B.n968 163.367
R1295 B.n968 B.n53 163.367
R1296 B.n964 B.n53 163.367
R1297 B.n964 B.n963 163.367
R1298 B.n963 B.n962 163.367
R1299 B.n962 B.n55 163.367
R1300 B.n958 B.n55 163.367
R1301 B.n958 B.n957 163.367
R1302 B.n957 B.n956 163.367
R1303 B.n956 B.n57 163.367
R1304 B.n952 B.n57 163.367
R1305 B.n952 B.n951 163.367
R1306 B.n951 B.n950 163.367
R1307 B.n950 B.n59 163.367
R1308 B.n946 B.n59 163.367
R1309 B.n946 B.n945 163.367
R1310 B.n945 B.n944 163.367
R1311 B.n944 B.n61 163.367
R1312 B.n940 B.n61 163.367
R1313 B.n940 B.n939 163.367
R1314 B.n939 B.n938 163.367
R1315 B.n938 B.n63 163.367
R1316 B.n934 B.n63 163.367
R1317 B.n934 B.n933 163.367
R1318 B.n933 B.n932 163.367
R1319 B.n932 B.n65 163.367
R1320 B.n928 B.n65 163.367
R1321 B.n928 B.n927 163.367
R1322 B.n927 B.n926 163.367
R1323 B.n926 B.n67 163.367
R1324 B.n922 B.n67 163.367
R1325 B.n922 B.n921 163.367
R1326 B.n921 B.n920 163.367
R1327 B.n920 B.n69 163.367
R1328 B.n916 B.n69 163.367
R1329 B.n916 B.n915 163.367
R1330 B.n915 B.n914 163.367
R1331 B.n914 B.n74 163.367
R1332 B.n910 B.n74 163.367
R1333 B.n910 B.n909 163.367
R1334 B.n909 B.n908 163.367
R1335 B.n908 B.n76 163.367
R1336 B.n903 B.n76 163.367
R1337 B.n903 B.n902 163.367
R1338 B.n902 B.n901 163.367
R1339 B.n901 B.n80 163.367
R1340 B.n897 B.n80 163.367
R1341 B.n897 B.n896 163.367
R1342 B.n896 B.n895 163.367
R1343 B.n895 B.n82 163.367
R1344 B.n891 B.n82 163.367
R1345 B.n891 B.n890 163.367
R1346 B.n890 B.n889 163.367
R1347 B.n889 B.n84 163.367
R1348 B.n885 B.n84 163.367
R1349 B.n885 B.n884 163.367
R1350 B.n884 B.n883 163.367
R1351 B.n883 B.n86 163.367
R1352 B.n879 B.n86 163.367
R1353 B.n879 B.n878 163.367
R1354 B.n878 B.n877 163.367
R1355 B.n877 B.n88 163.367
R1356 B.n873 B.n88 163.367
R1357 B.n873 B.n872 163.367
R1358 B.n872 B.n871 163.367
R1359 B.n871 B.n90 163.367
R1360 B.n867 B.n90 163.367
R1361 B.n867 B.n866 163.367
R1362 B.n866 B.n865 163.367
R1363 B.n865 B.n92 163.367
R1364 B.n861 B.n92 163.367
R1365 B.n861 B.n860 163.367
R1366 B.n860 B.n859 163.367
R1367 B.n859 B.n94 163.367
R1368 B.n855 B.n94 163.367
R1369 B.n855 B.n854 163.367
R1370 B.n854 B.n853 163.367
R1371 B.n853 B.n96 163.367
R1372 B.n849 B.n96 163.367
R1373 B.n849 B.n848 163.367
R1374 B.n848 B.n847 163.367
R1375 B.n847 B.n98 163.367
R1376 B.n843 B.n98 163.367
R1377 B.n843 B.n842 163.367
R1378 B.n842 B.n841 163.367
R1379 B.n841 B.n100 163.367
R1380 B.n837 B.n100 163.367
R1381 B.n837 B.n836 163.367
R1382 B.n836 B.n835 163.367
R1383 B.n835 B.n102 163.367
R1384 B.n831 B.n102 163.367
R1385 B.n831 B.n830 163.367
R1386 B.n830 B.n829 163.367
R1387 B.n829 B.n104 163.367
R1388 B.n825 B.n104 163.367
R1389 B.n825 B.n824 163.367
R1390 B.n824 B.n823 163.367
R1391 B.n823 B.n106 163.367
R1392 B.n819 B.n106 163.367
R1393 B.n819 B.n818 163.367
R1394 B.n818 B.n817 163.367
R1395 B.n1011 B.n1010 163.367
R1396 B.n1012 B.n1011 163.367
R1397 B.n1012 B.n37 163.367
R1398 B.n1016 B.n37 163.367
R1399 B.n1017 B.n1016 163.367
R1400 B.n1018 B.n1017 163.367
R1401 B.n1018 B.n35 163.367
R1402 B.n1022 B.n35 163.367
R1403 B.n1023 B.n1022 163.367
R1404 B.n1024 B.n1023 163.367
R1405 B.n1024 B.n33 163.367
R1406 B.n1028 B.n33 163.367
R1407 B.n1029 B.n1028 163.367
R1408 B.n1030 B.n1029 163.367
R1409 B.n1030 B.n31 163.367
R1410 B.n1034 B.n31 163.367
R1411 B.n1035 B.n1034 163.367
R1412 B.n1036 B.n1035 163.367
R1413 B.n1036 B.n29 163.367
R1414 B.n1040 B.n29 163.367
R1415 B.n1041 B.n1040 163.367
R1416 B.n1042 B.n1041 163.367
R1417 B.n1042 B.n27 163.367
R1418 B.n1046 B.n27 163.367
R1419 B.n1047 B.n1046 163.367
R1420 B.n1048 B.n1047 163.367
R1421 B.n1048 B.n25 163.367
R1422 B.n1052 B.n25 163.367
R1423 B.n1053 B.n1052 163.367
R1424 B.n1054 B.n1053 163.367
R1425 B.n1054 B.n23 163.367
R1426 B.n1058 B.n23 163.367
R1427 B.n1059 B.n1058 163.367
R1428 B.n1060 B.n1059 163.367
R1429 B.n1060 B.n21 163.367
R1430 B.n1064 B.n21 163.367
R1431 B.n1065 B.n1064 163.367
R1432 B.n1066 B.n1065 163.367
R1433 B.n1066 B.n19 163.367
R1434 B.n1070 B.n19 163.367
R1435 B.n1071 B.n1070 163.367
R1436 B.n1072 B.n1071 163.367
R1437 B.n1072 B.n17 163.367
R1438 B.n1076 B.n17 163.367
R1439 B.n1077 B.n1076 163.367
R1440 B.n1078 B.n1077 163.367
R1441 B.n1078 B.n15 163.367
R1442 B.n1082 B.n15 163.367
R1443 B.n1083 B.n1082 163.367
R1444 B.n1084 B.n1083 163.367
R1445 B.n1084 B.n13 163.367
R1446 B.n1088 B.n13 163.367
R1447 B.n1089 B.n1088 163.367
R1448 B.n1090 B.n1089 163.367
R1449 B.n1090 B.n11 163.367
R1450 B.n1094 B.n11 163.367
R1451 B.n1095 B.n1094 163.367
R1452 B.n1096 B.n1095 163.367
R1453 B.n1096 B.n9 163.367
R1454 B.n1100 B.n9 163.367
R1455 B.n1101 B.n1100 163.367
R1456 B.n1102 B.n1101 163.367
R1457 B.n1102 B.n7 163.367
R1458 B.n1106 B.n7 163.367
R1459 B.n1107 B.n1106 163.367
R1460 B.n1108 B.n1107 163.367
R1461 B.n1108 B.n5 163.367
R1462 B.n1112 B.n5 163.367
R1463 B.n1113 B.n1112 163.367
R1464 B.n1114 B.n1113 163.367
R1465 B.n1114 B.n3 163.367
R1466 B.n1118 B.n3 163.367
R1467 B.n1119 B.n1118 163.367
R1468 B.n286 B.n2 163.367
R1469 B.n287 B.n286 163.367
R1470 B.n287 B.n284 163.367
R1471 B.n291 B.n284 163.367
R1472 B.n292 B.n291 163.367
R1473 B.n293 B.n292 163.367
R1474 B.n293 B.n282 163.367
R1475 B.n297 B.n282 163.367
R1476 B.n298 B.n297 163.367
R1477 B.n299 B.n298 163.367
R1478 B.n299 B.n280 163.367
R1479 B.n303 B.n280 163.367
R1480 B.n304 B.n303 163.367
R1481 B.n305 B.n304 163.367
R1482 B.n305 B.n278 163.367
R1483 B.n309 B.n278 163.367
R1484 B.n310 B.n309 163.367
R1485 B.n311 B.n310 163.367
R1486 B.n311 B.n276 163.367
R1487 B.n315 B.n276 163.367
R1488 B.n316 B.n315 163.367
R1489 B.n317 B.n316 163.367
R1490 B.n317 B.n274 163.367
R1491 B.n321 B.n274 163.367
R1492 B.n322 B.n321 163.367
R1493 B.n323 B.n322 163.367
R1494 B.n323 B.n272 163.367
R1495 B.n327 B.n272 163.367
R1496 B.n328 B.n327 163.367
R1497 B.n329 B.n328 163.367
R1498 B.n329 B.n270 163.367
R1499 B.n333 B.n270 163.367
R1500 B.n334 B.n333 163.367
R1501 B.n335 B.n334 163.367
R1502 B.n335 B.n268 163.367
R1503 B.n339 B.n268 163.367
R1504 B.n340 B.n339 163.367
R1505 B.n341 B.n340 163.367
R1506 B.n341 B.n266 163.367
R1507 B.n345 B.n266 163.367
R1508 B.n346 B.n345 163.367
R1509 B.n347 B.n346 163.367
R1510 B.n347 B.n264 163.367
R1511 B.n351 B.n264 163.367
R1512 B.n352 B.n351 163.367
R1513 B.n353 B.n352 163.367
R1514 B.n353 B.n262 163.367
R1515 B.n357 B.n262 163.367
R1516 B.n358 B.n357 163.367
R1517 B.n359 B.n358 163.367
R1518 B.n359 B.n260 163.367
R1519 B.n363 B.n260 163.367
R1520 B.n364 B.n363 163.367
R1521 B.n365 B.n364 163.367
R1522 B.n365 B.n258 163.367
R1523 B.n369 B.n258 163.367
R1524 B.n370 B.n369 163.367
R1525 B.n371 B.n370 163.367
R1526 B.n371 B.n256 163.367
R1527 B.n375 B.n256 163.367
R1528 B.n376 B.n375 163.367
R1529 B.n377 B.n376 163.367
R1530 B.n377 B.n254 163.367
R1531 B.n381 B.n254 163.367
R1532 B.n382 B.n381 163.367
R1533 B.n383 B.n382 163.367
R1534 B.n383 B.n252 163.367
R1535 B.n387 B.n252 163.367
R1536 B.n388 B.n387 163.367
R1537 B.n389 B.n388 163.367
R1538 B.n389 B.n250 163.367
R1539 B.n393 B.n250 163.367
R1540 B.n394 B.n393 163.367
R1541 B.n214 B.t5 110.867
R1542 B.n78 B.t1 110.867
R1543 B.n483 B.t11 110.844
R1544 B.n71 B.t7 110.844
R1545 B.n483 B.n482 73.1157
R1546 B.n214 B.n213 73.1157
R1547 B.n78 B.n77 73.1157
R1548 B.n71 B.n70 73.1157
R1549 B.n484 B.n483 59.5399
R1550 B.n502 B.n214 59.5399
R1551 B.n905 B.n78 59.5399
R1552 B.n72 B.n71 59.5399
R1553 B.n1009 B.n1008 32.0005
R1554 B.n816 B.n815 32.0005
R1555 B.n592 B.n183 32.0005
R1556 B.n396 B.n249 32.0005
R1557 B B.n1121 18.0485
R1558 B.n1009 B.n38 10.6151
R1559 B.n1013 B.n38 10.6151
R1560 B.n1014 B.n1013 10.6151
R1561 B.n1015 B.n1014 10.6151
R1562 B.n1015 B.n36 10.6151
R1563 B.n1019 B.n36 10.6151
R1564 B.n1020 B.n1019 10.6151
R1565 B.n1021 B.n1020 10.6151
R1566 B.n1021 B.n34 10.6151
R1567 B.n1025 B.n34 10.6151
R1568 B.n1026 B.n1025 10.6151
R1569 B.n1027 B.n1026 10.6151
R1570 B.n1027 B.n32 10.6151
R1571 B.n1031 B.n32 10.6151
R1572 B.n1032 B.n1031 10.6151
R1573 B.n1033 B.n1032 10.6151
R1574 B.n1033 B.n30 10.6151
R1575 B.n1037 B.n30 10.6151
R1576 B.n1038 B.n1037 10.6151
R1577 B.n1039 B.n1038 10.6151
R1578 B.n1039 B.n28 10.6151
R1579 B.n1043 B.n28 10.6151
R1580 B.n1044 B.n1043 10.6151
R1581 B.n1045 B.n1044 10.6151
R1582 B.n1045 B.n26 10.6151
R1583 B.n1049 B.n26 10.6151
R1584 B.n1050 B.n1049 10.6151
R1585 B.n1051 B.n1050 10.6151
R1586 B.n1051 B.n24 10.6151
R1587 B.n1055 B.n24 10.6151
R1588 B.n1056 B.n1055 10.6151
R1589 B.n1057 B.n1056 10.6151
R1590 B.n1057 B.n22 10.6151
R1591 B.n1061 B.n22 10.6151
R1592 B.n1062 B.n1061 10.6151
R1593 B.n1063 B.n1062 10.6151
R1594 B.n1063 B.n20 10.6151
R1595 B.n1067 B.n20 10.6151
R1596 B.n1068 B.n1067 10.6151
R1597 B.n1069 B.n1068 10.6151
R1598 B.n1069 B.n18 10.6151
R1599 B.n1073 B.n18 10.6151
R1600 B.n1074 B.n1073 10.6151
R1601 B.n1075 B.n1074 10.6151
R1602 B.n1075 B.n16 10.6151
R1603 B.n1079 B.n16 10.6151
R1604 B.n1080 B.n1079 10.6151
R1605 B.n1081 B.n1080 10.6151
R1606 B.n1081 B.n14 10.6151
R1607 B.n1085 B.n14 10.6151
R1608 B.n1086 B.n1085 10.6151
R1609 B.n1087 B.n1086 10.6151
R1610 B.n1087 B.n12 10.6151
R1611 B.n1091 B.n12 10.6151
R1612 B.n1092 B.n1091 10.6151
R1613 B.n1093 B.n1092 10.6151
R1614 B.n1093 B.n10 10.6151
R1615 B.n1097 B.n10 10.6151
R1616 B.n1098 B.n1097 10.6151
R1617 B.n1099 B.n1098 10.6151
R1618 B.n1099 B.n8 10.6151
R1619 B.n1103 B.n8 10.6151
R1620 B.n1104 B.n1103 10.6151
R1621 B.n1105 B.n1104 10.6151
R1622 B.n1105 B.n6 10.6151
R1623 B.n1109 B.n6 10.6151
R1624 B.n1110 B.n1109 10.6151
R1625 B.n1111 B.n1110 10.6151
R1626 B.n1111 B.n4 10.6151
R1627 B.n1115 B.n4 10.6151
R1628 B.n1116 B.n1115 10.6151
R1629 B.n1117 B.n1116 10.6151
R1630 B.n1117 B.n0 10.6151
R1631 B.n1008 B.n1007 10.6151
R1632 B.n1007 B.n40 10.6151
R1633 B.n1003 B.n40 10.6151
R1634 B.n1003 B.n1002 10.6151
R1635 B.n1002 B.n1001 10.6151
R1636 B.n1001 B.n42 10.6151
R1637 B.n997 B.n42 10.6151
R1638 B.n997 B.n996 10.6151
R1639 B.n996 B.n995 10.6151
R1640 B.n995 B.n44 10.6151
R1641 B.n991 B.n44 10.6151
R1642 B.n991 B.n990 10.6151
R1643 B.n990 B.n989 10.6151
R1644 B.n989 B.n46 10.6151
R1645 B.n985 B.n46 10.6151
R1646 B.n985 B.n984 10.6151
R1647 B.n984 B.n983 10.6151
R1648 B.n983 B.n48 10.6151
R1649 B.n979 B.n48 10.6151
R1650 B.n979 B.n978 10.6151
R1651 B.n978 B.n977 10.6151
R1652 B.n977 B.n50 10.6151
R1653 B.n973 B.n50 10.6151
R1654 B.n973 B.n972 10.6151
R1655 B.n972 B.n971 10.6151
R1656 B.n971 B.n52 10.6151
R1657 B.n967 B.n52 10.6151
R1658 B.n967 B.n966 10.6151
R1659 B.n966 B.n965 10.6151
R1660 B.n965 B.n54 10.6151
R1661 B.n961 B.n54 10.6151
R1662 B.n961 B.n960 10.6151
R1663 B.n960 B.n959 10.6151
R1664 B.n959 B.n56 10.6151
R1665 B.n955 B.n56 10.6151
R1666 B.n955 B.n954 10.6151
R1667 B.n954 B.n953 10.6151
R1668 B.n953 B.n58 10.6151
R1669 B.n949 B.n58 10.6151
R1670 B.n949 B.n948 10.6151
R1671 B.n948 B.n947 10.6151
R1672 B.n947 B.n60 10.6151
R1673 B.n943 B.n60 10.6151
R1674 B.n943 B.n942 10.6151
R1675 B.n942 B.n941 10.6151
R1676 B.n941 B.n62 10.6151
R1677 B.n937 B.n62 10.6151
R1678 B.n937 B.n936 10.6151
R1679 B.n936 B.n935 10.6151
R1680 B.n935 B.n64 10.6151
R1681 B.n931 B.n64 10.6151
R1682 B.n931 B.n930 10.6151
R1683 B.n930 B.n929 10.6151
R1684 B.n929 B.n66 10.6151
R1685 B.n925 B.n66 10.6151
R1686 B.n925 B.n924 10.6151
R1687 B.n924 B.n923 10.6151
R1688 B.n923 B.n68 10.6151
R1689 B.n919 B.n918 10.6151
R1690 B.n918 B.n917 10.6151
R1691 B.n917 B.n73 10.6151
R1692 B.n913 B.n73 10.6151
R1693 B.n913 B.n912 10.6151
R1694 B.n912 B.n911 10.6151
R1695 B.n911 B.n75 10.6151
R1696 B.n907 B.n75 10.6151
R1697 B.n907 B.n906 10.6151
R1698 B.n904 B.n79 10.6151
R1699 B.n900 B.n79 10.6151
R1700 B.n900 B.n899 10.6151
R1701 B.n899 B.n898 10.6151
R1702 B.n898 B.n81 10.6151
R1703 B.n894 B.n81 10.6151
R1704 B.n894 B.n893 10.6151
R1705 B.n893 B.n892 10.6151
R1706 B.n892 B.n83 10.6151
R1707 B.n888 B.n83 10.6151
R1708 B.n888 B.n887 10.6151
R1709 B.n887 B.n886 10.6151
R1710 B.n886 B.n85 10.6151
R1711 B.n882 B.n85 10.6151
R1712 B.n882 B.n881 10.6151
R1713 B.n881 B.n880 10.6151
R1714 B.n880 B.n87 10.6151
R1715 B.n876 B.n87 10.6151
R1716 B.n876 B.n875 10.6151
R1717 B.n875 B.n874 10.6151
R1718 B.n874 B.n89 10.6151
R1719 B.n870 B.n89 10.6151
R1720 B.n870 B.n869 10.6151
R1721 B.n869 B.n868 10.6151
R1722 B.n868 B.n91 10.6151
R1723 B.n864 B.n91 10.6151
R1724 B.n864 B.n863 10.6151
R1725 B.n863 B.n862 10.6151
R1726 B.n862 B.n93 10.6151
R1727 B.n858 B.n93 10.6151
R1728 B.n858 B.n857 10.6151
R1729 B.n857 B.n856 10.6151
R1730 B.n856 B.n95 10.6151
R1731 B.n852 B.n95 10.6151
R1732 B.n852 B.n851 10.6151
R1733 B.n851 B.n850 10.6151
R1734 B.n850 B.n97 10.6151
R1735 B.n846 B.n97 10.6151
R1736 B.n846 B.n845 10.6151
R1737 B.n845 B.n844 10.6151
R1738 B.n844 B.n99 10.6151
R1739 B.n840 B.n99 10.6151
R1740 B.n840 B.n839 10.6151
R1741 B.n839 B.n838 10.6151
R1742 B.n838 B.n101 10.6151
R1743 B.n834 B.n101 10.6151
R1744 B.n834 B.n833 10.6151
R1745 B.n833 B.n832 10.6151
R1746 B.n832 B.n103 10.6151
R1747 B.n828 B.n103 10.6151
R1748 B.n828 B.n827 10.6151
R1749 B.n827 B.n826 10.6151
R1750 B.n826 B.n105 10.6151
R1751 B.n822 B.n105 10.6151
R1752 B.n822 B.n821 10.6151
R1753 B.n821 B.n820 10.6151
R1754 B.n820 B.n107 10.6151
R1755 B.n816 B.n107 10.6151
R1756 B.n815 B.n814 10.6151
R1757 B.n814 B.n109 10.6151
R1758 B.n810 B.n109 10.6151
R1759 B.n810 B.n809 10.6151
R1760 B.n809 B.n808 10.6151
R1761 B.n808 B.n111 10.6151
R1762 B.n804 B.n111 10.6151
R1763 B.n804 B.n803 10.6151
R1764 B.n803 B.n802 10.6151
R1765 B.n802 B.n113 10.6151
R1766 B.n798 B.n113 10.6151
R1767 B.n798 B.n797 10.6151
R1768 B.n797 B.n796 10.6151
R1769 B.n796 B.n115 10.6151
R1770 B.n792 B.n115 10.6151
R1771 B.n792 B.n791 10.6151
R1772 B.n791 B.n790 10.6151
R1773 B.n790 B.n117 10.6151
R1774 B.n786 B.n117 10.6151
R1775 B.n786 B.n785 10.6151
R1776 B.n785 B.n784 10.6151
R1777 B.n784 B.n119 10.6151
R1778 B.n780 B.n119 10.6151
R1779 B.n780 B.n779 10.6151
R1780 B.n779 B.n778 10.6151
R1781 B.n778 B.n121 10.6151
R1782 B.n774 B.n121 10.6151
R1783 B.n774 B.n773 10.6151
R1784 B.n773 B.n772 10.6151
R1785 B.n772 B.n123 10.6151
R1786 B.n768 B.n123 10.6151
R1787 B.n768 B.n767 10.6151
R1788 B.n767 B.n766 10.6151
R1789 B.n766 B.n125 10.6151
R1790 B.n762 B.n125 10.6151
R1791 B.n762 B.n761 10.6151
R1792 B.n761 B.n760 10.6151
R1793 B.n760 B.n127 10.6151
R1794 B.n756 B.n127 10.6151
R1795 B.n756 B.n755 10.6151
R1796 B.n755 B.n754 10.6151
R1797 B.n754 B.n129 10.6151
R1798 B.n750 B.n129 10.6151
R1799 B.n750 B.n749 10.6151
R1800 B.n749 B.n748 10.6151
R1801 B.n748 B.n131 10.6151
R1802 B.n744 B.n131 10.6151
R1803 B.n744 B.n743 10.6151
R1804 B.n743 B.n742 10.6151
R1805 B.n742 B.n133 10.6151
R1806 B.n738 B.n133 10.6151
R1807 B.n738 B.n737 10.6151
R1808 B.n737 B.n736 10.6151
R1809 B.n736 B.n135 10.6151
R1810 B.n732 B.n135 10.6151
R1811 B.n732 B.n731 10.6151
R1812 B.n731 B.n730 10.6151
R1813 B.n730 B.n137 10.6151
R1814 B.n726 B.n137 10.6151
R1815 B.n726 B.n725 10.6151
R1816 B.n725 B.n724 10.6151
R1817 B.n724 B.n139 10.6151
R1818 B.n720 B.n139 10.6151
R1819 B.n720 B.n719 10.6151
R1820 B.n719 B.n718 10.6151
R1821 B.n718 B.n141 10.6151
R1822 B.n714 B.n141 10.6151
R1823 B.n714 B.n713 10.6151
R1824 B.n713 B.n712 10.6151
R1825 B.n712 B.n143 10.6151
R1826 B.n708 B.n143 10.6151
R1827 B.n708 B.n707 10.6151
R1828 B.n707 B.n706 10.6151
R1829 B.n706 B.n145 10.6151
R1830 B.n702 B.n145 10.6151
R1831 B.n702 B.n701 10.6151
R1832 B.n701 B.n700 10.6151
R1833 B.n700 B.n147 10.6151
R1834 B.n696 B.n147 10.6151
R1835 B.n696 B.n695 10.6151
R1836 B.n695 B.n694 10.6151
R1837 B.n694 B.n149 10.6151
R1838 B.n690 B.n149 10.6151
R1839 B.n690 B.n689 10.6151
R1840 B.n689 B.n688 10.6151
R1841 B.n688 B.n151 10.6151
R1842 B.n684 B.n151 10.6151
R1843 B.n684 B.n683 10.6151
R1844 B.n683 B.n682 10.6151
R1845 B.n682 B.n153 10.6151
R1846 B.n678 B.n153 10.6151
R1847 B.n678 B.n677 10.6151
R1848 B.n677 B.n676 10.6151
R1849 B.n676 B.n155 10.6151
R1850 B.n672 B.n155 10.6151
R1851 B.n672 B.n671 10.6151
R1852 B.n671 B.n670 10.6151
R1853 B.n670 B.n157 10.6151
R1854 B.n666 B.n157 10.6151
R1855 B.n666 B.n665 10.6151
R1856 B.n665 B.n664 10.6151
R1857 B.n664 B.n159 10.6151
R1858 B.n660 B.n159 10.6151
R1859 B.n660 B.n659 10.6151
R1860 B.n659 B.n658 10.6151
R1861 B.n658 B.n161 10.6151
R1862 B.n654 B.n161 10.6151
R1863 B.n654 B.n653 10.6151
R1864 B.n653 B.n652 10.6151
R1865 B.n652 B.n163 10.6151
R1866 B.n648 B.n163 10.6151
R1867 B.n648 B.n647 10.6151
R1868 B.n647 B.n646 10.6151
R1869 B.n646 B.n165 10.6151
R1870 B.n642 B.n165 10.6151
R1871 B.n642 B.n641 10.6151
R1872 B.n641 B.n640 10.6151
R1873 B.n640 B.n167 10.6151
R1874 B.n636 B.n167 10.6151
R1875 B.n636 B.n635 10.6151
R1876 B.n635 B.n634 10.6151
R1877 B.n634 B.n169 10.6151
R1878 B.n630 B.n169 10.6151
R1879 B.n630 B.n629 10.6151
R1880 B.n629 B.n628 10.6151
R1881 B.n628 B.n171 10.6151
R1882 B.n624 B.n171 10.6151
R1883 B.n624 B.n623 10.6151
R1884 B.n623 B.n622 10.6151
R1885 B.n622 B.n173 10.6151
R1886 B.n618 B.n173 10.6151
R1887 B.n618 B.n617 10.6151
R1888 B.n617 B.n616 10.6151
R1889 B.n616 B.n175 10.6151
R1890 B.n612 B.n175 10.6151
R1891 B.n612 B.n611 10.6151
R1892 B.n611 B.n610 10.6151
R1893 B.n610 B.n177 10.6151
R1894 B.n606 B.n177 10.6151
R1895 B.n606 B.n605 10.6151
R1896 B.n605 B.n604 10.6151
R1897 B.n604 B.n179 10.6151
R1898 B.n600 B.n179 10.6151
R1899 B.n600 B.n599 10.6151
R1900 B.n599 B.n598 10.6151
R1901 B.n598 B.n181 10.6151
R1902 B.n594 B.n181 10.6151
R1903 B.n594 B.n593 10.6151
R1904 B.n593 B.n592 10.6151
R1905 B.n285 B.n1 10.6151
R1906 B.n288 B.n285 10.6151
R1907 B.n289 B.n288 10.6151
R1908 B.n290 B.n289 10.6151
R1909 B.n290 B.n283 10.6151
R1910 B.n294 B.n283 10.6151
R1911 B.n295 B.n294 10.6151
R1912 B.n296 B.n295 10.6151
R1913 B.n296 B.n281 10.6151
R1914 B.n300 B.n281 10.6151
R1915 B.n301 B.n300 10.6151
R1916 B.n302 B.n301 10.6151
R1917 B.n302 B.n279 10.6151
R1918 B.n306 B.n279 10.6151
R1919 B.n307 B.n306 10.6151
R1920 B.n308 B.n307 10.6151
R1921 B.n308 B.n277 10.6151
R1922 B.n312 B.n277 10.6151
R1923 B.n313 B.n312 10.6151
R1924 B.n314 B.n313 10.6151
R1925 B.n314 B.n275 10.6151
R1926 B.n318 B.n275 10.6151
R1927 B.n319 B.n318 10.6151
R1928 B.n320 B.n319 10.6151
R1929 B.n320 B.n273 10.6151
R1930 B.n324 B.n273 10.6151
R1931 B.n325 B.n324 10.6151
R1932 B.n326 B.n325 10.6151
R1933 B.n326 B.n271 10.6151
R1934 B.n330 B.n271 10.6151
R1935 B.n331 B.n330 10.6151
R1936 B.n332 B.n331 10.6151
R1937 B.n332 B.n269 10.6151
R1938 B.n336 B.n269 10.6151
R1939 B.n337 B.n336 10.6151
R1940 B.n338 B.n337 10.6151
R1941 B.n338 B.n267 10.6151
R1942 B.n342 B.n267 10.6151
R1943 B.n343 B.n342 10.6151
R1944 B.n344 B.n343 10.6151
R1945 B.n344 B.n265 10.6151
R1946 B.n348 B.n265 10.6151
R1947 B.n349 B.n348 10.6151
R1948 B.n350 B.n349 10.6151
R1949 B.n350 B.n263 10.6151
R1950 B.n354 B.n263 10.6151
R1951 B.n355 B.n354 10.6151
R1952 B.n356 B.n355 10.6151
R1953 B.n356 B.n261 10.6151
R1954 B.n360 B.n261 10.6151
R1955 B.n361 B.n360 10.6151
R1956 B.n362 B.n361 10.6151
R1957 B.n362 B.n259 10.6151
R1958 B.n366 B.n259 10.6151
R1959 B.n367 B.n366 10.6151
R1960 B.n368 B.n367 10.6151
R1961 B.n368 B.n257 10.6151
R1962 B.n372 B.n257 10.6151
R1963 B.n373 B.n372 10.6151
R1964 B.n374 B.n373 10.6151
R1965 B.n374 B.n255 10.6151
R1966 B.n378 B.n255 10.6151
R1967 B.n379 B.n378 10.6151
R1968 B.n380 B.n379 10.6151
R1969 B.n380 B.n253 10.6151
R1970 B.n384 B.n253 10.6151
R1971 B.n385 B.n384 10.6151
R1972 B.n386 B.n385 10.6151
R1973 B.n386 B.n251 10.6151
R1974 B.n390 B.n251 10.6151
R1975 B.n391 B.n390 10.6151
R1976 B.n392 B.n391 10.6151
R1977 B.n392 B.n249 10.6151
R1978 B.n397 B.n396 10.6151
R1979 B.n398 B.n397 10.6151
R1980 B.n398 B.n247 10.6151
R1981 B.n402 B.n247 10.6151
R1982 B.n403 B.n402 10.6151
R1983 B.n404 B.n403 10.6151
R1984 B.n404 B.n245 10.6151
R1985 B.n408 B.n245 10.6151
R1986 B.n409 B.n408 10.6151
R1987 B.n410 B.n409 10.6151
R1988 B.n410 B.n243 10.6151
R1989 B.n414 B.n243 10.6151
R1990 B.n415 B.n414 10.6151
R1991 B.n416 B.n415 10.6151
R1992 B.n416 B.n241 10.6151
R1993 B.n420 B.n241 10.6151
R1994 B.n421 B.n420 10.6151
R1995 B.n422 B.n421 10.6151
R1996 B.n422 B.n239 10.6151
R1997 B.n426 B.n239 10.6151
R1998 B.n427 B.n426 10.6151
R1999 B.n428 B.n427 10.6151
R2000 B.n428 B.n237 10.6151
R2001 B.n432 B.n237 10.6151
R2002 B.n433 B.n432 10.6151
R2003 B.n434 B.n433 10.6151
R2004 B.n434 B.n235 10.6151
R2005 B.n438 B.n235 10.6151
R2006 B.n439 B.n438 10.6151
R2007 B.n440 B.n439 10.6151
R2008 B.n440 B.n233 10.6151
R2009 B.n444 B.n233 10.6151
R2010 B.n445 B.n444 10.6151
R2011 B.n446 B.n445 10.6151
R2012 B.n446 B.n231 10.6151
R2013 B.n450 B.n231 10.6151
R2014 B.n451 B.n450 10.6151
R2015 B.n452 B.n451 10.6151
R2016 B.n452 B.n229 10.6151
R2017 B.n456 B.n229 10.6151
R2018 B.n457 B.n456 10.6151
R2019 B.n458 B.n457 10.6151
R2020 B.n458 B.n227 10.6151
R2021 B.n462 B.n227 10.6151
R2022 B.n463 B.n462 10.6151
R2023 B.n464 B.n463 10.6151
R2024 B.n464 B.n225 10.6151
R2025 B.n468 B.n225 10.6151
R2026 B.n469 B.n468 10.6151
R2027 B.n470 B.n469 10.6151
R2028 B.n470 B.n223 10.6151
R2029 B.n474 B.n223 10.6151
R2030 B.n475 B.n474 10.6151
R2031 B.n476 B.n475 10.6151
R2032 B.n476 B.n221 10.6151
R2033 B.n480 B.n221 10.6151
R2034 B.n481 B.n480 10.6151
R2035 B.n485 B.n481 10.6151
R2036 B.n489 B.n219 10.6151
R2037 B.n490 B.n489 10.6151
R2038 B.n491 B.n490 10.6151
R2039 B.n491 B.n217 10.6151
R2040 B.n495 B.n217 10.6151
R2041 B.n496 B.n495 10.6151
R2042 B.n497 B.n496 10.6151
R2043 B.n497 B.n215 10.6151
R2044 B.n501 B.n215 10.6151
R2045 B.n504 B.n503 10.6151
R2046 B.n504 B.n211 10.6151
R2047 B.n508 B.n211 10.6151
R2048 B.n509 B.n508 10.6151
R2049 B.n510 B.n509 10.6151
R2050 B.n510 B.n209 10.6151
R2051 B.n514 B.n209 10.6151
R2052 B.n515 B.n514 10.6151
R2053 B.n516 B.n515 10.6151
R2054 B.n516 B.n207 10.6151
R2055 B.n520 B.n207 10.6151
R2056 B.n521 B.n520 10.6151
R2057 B.n522 B.n521 10.6151
R2058 B.n522 B.n205 10.6151
R2059 B.n526 B.n205 10.6151
R2060 B.n527 B.n526 10.6151
R2061 B.n528 B.n527 10.6151
R2062 B.n528 B.n203 10.6151
R2063 B.n532 B.n203 10.6151
R2064 B.n533 B.n532 10.6151
R2065 B.n534 B.n533 10.6151
R2066 B.n534 B.n201 10.6151
R2067 B.n538 B.n201 10.6151
R2068 B.n539 B.n538 10.6151
R2069 B.n540 B.n539 10.6151
R2070 B.n540 B.n199 10.6151
R2071 B.n544 B.n199 10.6151
R2072 B.n545 B.n544 10.6151
R2073 B.n546 B.n545 10.6151
R2074 B.n546 B.n197 10.6151
R2075 B.n550 B.n197 10.6151
R2076 B.n551 B.n550 10.6151
R2077 B.n552 B.n551 10.6151
R2078 B.n552 B.n195 10.6151
R2079 B.n556 B.n195 10.6151
R2080 B.n557 B.n556 10.6151
R2081 B.n558 B.n557 10.6151
R2082 B.n558 B.n193 10.6151
R2083 B.n562 B.n193 10.6151
R2084 B.n563 B.n562 10.6151
R2085 B.n564 B.n563 10.6151
R2086 B.n564 B.n191 10.6151
R2087 B.n568 B.n191 10.6151
R2088 B.n569 B.n568 10.6151
R2089 B.n570 B.n569 10.6151
R2090 B.n570 B.n189 10.6151
R2091 B.n574 B.n189 10.6151
R2092 B.n575 B.n574 10.6151
R2093 B.n576 B.n575 10.6151
R2094 B.n576 B.n187 10.6151
R2095 B.n580 B.n187 10.6151
R2096 B.n581 B.n580 10.6151
R2097 B.n582 B.n581 10.6151
R2098 B.n582 B.n185 10.6151
R2099 B.n586 B.n185 10.6151
R2100 B.n587 B.n586 10.6151
R2101 B.n588 B.n587 10.6151
R2102 B.n588 B.n183 10.6151
R2103 B.n72 B.n68 9.36635
R2104 B.n905 B.n904 9.36635
R2105 B.n485 B.n484 9.36635
R2106 B.n503 B.n502 9.36635
R2107 B.n1121 B.n0 8.11757
R2108 B.n1121 B.n1 8.11757
R2109 B.n919 B.n72 1.24928
R2110 B.n906 B.n905 1.24928
R2111 B.n484 B.n219 1.24928
R2112 B.n502 B.n501 1.24928
C0 VDD1 w_n5494_n4552# 3.51327f
C1 VTAIL VDD1 13.157499f
C2 B VN 1.56208f
C3 VN VP 10.740701f
C4 VN VDD2 16.470499f
C5 B w_n5494_n4552# 13.6187f
C6 w_n5494_n4552# VP 12.8468f
C7 VTAIL B 5.44714f
C8 VTAIL VP 17.2089f
C9 w_n5494_n4552# VDD2 3.70048f
C10 VTAIL VDD2 13.213799f
C11 VDD1 B 3.28301f
C12 VN w_n5494_n4552# 12.128901f
C13 VDD1 VP 17.0016f
C14 VTAIL VN 17.1946f
C15 VDD1 VDD2 2.72196f
C16 VTAIL w_n5494_n4552# 4.13629f
C17 B VP 2.77387f
C18 VDD1 VN 0.154927f
C19 B VDD2 3.43363f
C20 VDD2 VP 0.690779f
C21 VDD2 VSUBS 2.58153f
C22 VDD1 VSUBS 2.455104f
C23 VTAIL VSUBS 1.70142f
C24 VN VSUBS 9.27621f
C25 VP VSUBS 5.527499f
C26 B VSUBS 6.907479f
C27 w_n5494_n4552# VSUBS 0.30584p
C28 B.n0 VSUBS 0.00679f
C29 B.n1 VSUBS 0.00679f
C30 B.n2 VSUBS 0.010042f
C31 B.n3 VSUBS 0.007695f
C32 B.n4 VSUBS 0.007695f
C33 B.n5 VSUBS 0.007695f
C34 B.n6 VSUBS 0.007695f
C35 B.n7 VSUBS 0.007695f
C36 B.n8 VSUBS 0.007695f
C37 B.n9 VSUBS 0.007695f
C38 B.n10 VSUBS 0.007695f
C39 B.n11 VSUBS 0.007695f
C40 B.n12 VSUBS 0.007695f
C41 B.n13 VSUBS 0.007695f
C42 B.n14 VSUBS 0.007695f
C43 B.n15 VSUBS 0.007695f
C44 B.n16 VSUBS 0.007695f
C45 B.n17 VSUBS 0.007695f
C46 B.n18 VSUBS 0.007695f
C47 B.n19 VSUBS 0.007695f
C48 B.n20 VSUBS 0.007695f
C49 B.n21 VSUBS 0.007695f
C50 B.n22 VSUBS 0.007695f
C51 B.n23 VSUBS 0.007695f
C52 B.n24 VSUBS 0.007695f
C53 B.n25 VSUBS 0.007695f
C54 B.n26 VSUBS 0.007695f
C55 B.n27 VSUBS 0.007695f
C56 B.n28 VSUBS 0.007695f
C57 B.n29 VSUBS 0.007695f
C58 B.n30 VSUBS 0.007695f
C59 B.n31 VSUBS 0.007695f
C60 B.n32 VSUBS 0.007695f
C61 B.n33 VSUBS 0.007695f
C62 B.n34 VSUBS 0.007695f
C63 B.n35 VSUBS 0.007695f
C64 B.n36 VSUBS 0.007695f
C65 B.n37 VSUBS 0.007695f
C66 B.n38 VSUBS 0.007695f
C67 B.n39 VSUBS 0.018457f
C68 B.n40 VSUBS 0.007695f
C69 B.n41 VSUBS 0.007695f
C70 B.n42 VSUBS 0.007695f
C71 B.n43 VSUBS 0.007695f
C72 B.n44 VSUBS 0.007695f
C73 B.n45 VSUBS 0.007695f
C74 B.n46 VSUBS 0.007695f
C75 B.n47 VSUBS 0.007695f
C76 B.n48 VSUBS 0.007695f
C77 B.n49 VSUBS 0.007695f
C78 B.n50 VSUBS 0.007695f
C79 B.n51 VSUBS 0.007695f
C80 B.n52 VSUBS 0.007695f
C81 B.n53 VSUBS 0.007695f
C82 B.n54 VSUBS 0.007695f
C83 B.n55 VSUBS 0.007695f
C84 B.n56 VSUBS 0.007695f
C85 B.n57 VSUBS 0.007695f
C86 B.n58 VSUBS 0.007695f
C87 B.n59 VSUBS 0.007695f
C88 B.n60 VSUBS 0.007695f
C89 B.n61 VSUBS 0.007695f
C90 B.n62 VSUBS 0.007695f
C91 B.n63 VSUBS 0.007695f
C92 B.n64 VSUBS 0.007695f
C93 B.n65 VSUBS 0.007695f
C94 B.n66 VSUBS 0.007695f
C95 B.n67 VSUBS 0.007695f
C96 B.n68 VSUBS 0.007242f
C97 B.n69 VSUBS 0.007695f
C98 B.t7 VSUBS 0.664853f
C99 B.t8 VSUBS 0.693509f
C100 B.t6 VSUBS 3.06798f
C101 B.n70 VSUBS 0.418657f
C102 B.n71 VSUBS 0.083075f
C103 B.n72 VSUBS 0.017828f
C104 B.n73 VSUBS 0.007695f
C105 B.n74 VSUBS 0.007695f
C106 B.n75 VSUBS 0.007695f
C107 B.n76 VSUBS 0.007695f
C108 B.t1 VSUBS 0.664829f
C109 B.t2 VSUBS 0.693491f
C110 B.t0 VSUBS 3.06798f
C111 B.n77 VSUBS 0.418675f
C112 B.n78 VSUBS 0.083099f
C113 B.n79 VSUBS 0.007695f
C114 B.n80 VSUBS 0.007695f
C115 B.n81 VSUBS 0.007695f
C116 B.n82 VSUBS 0.007695f
C117 B.n83 VSUBS 0.007695f
C118 B.n84 VSUBS 0.007695f
C119 B.n85 VSUBS 0.007695f
C120 B.n86 VSUBS 0.007695f
C121 B.n87 VSUBS 0.007695f
C122 B.n88 VSUBS 0.007695f
C123 B.n89 VSUBS 0.007695f
C124 B.n90 VSUBS 0.007695f
C125 B.n91 VSUBS 0.007695f
C126 B.n92 VSUBS 0.007695f
C127 B.n93 VSUBS 0.007695f
C128 B.n94 VSUBS 0.007695f
C129 B.n95 VSUBS 0.007695f
C130 B.n96 VSUBS 0.007695f
C131 B.n97 VSUBS 0.007695f
C132 B.n98 VSUBS 0.007695f
C133 B.n99 VSUBS 0.007695f
C134 B.n100 VSUBS 0.007695f
C135 B.n101 VSUBS 0.007695f
C136 B.n102 VSUBS 0.007695f
C137 B.n103 VSUBS 0.007695f
C138 B.n104 VSUBS 0.007695f
C139 B.n105 VSUBS 0.007695f
C140 B.n106 VSUBS 0.007695f
C141 B.n107 VSUBS 0.007695f
C142 B.n108 VSUBS 0.017076f
C143 B.n109 VSUBS 0.007695f
C144 B.n110 VSUBS 0.007695f
C145 B.n111 VSUBS 0.007695f
C146 B.n112 VSUBS 0.007695f
C147 B.n113 VSUBS 0.007695f
C148 B.n114 VSUBS 0.007695f
C149 B.n115 VSUBS 0.007695f
C150 B.n116 VSUBS 0.007695f
C151 B.n117 VSUBS 0.007695f
C152 B.n118 VSUBS 0.007695f
C153 B.n119 VSUBS 0.007695f
C154 B.n120 VSUBS 0.007695f
C155 B.n121 VSUBS 0.007695f
C156 B.n122 VSUBS 0.007695f
C157 B.n123 VSUBS 0.007695f
C158 B.n124 VSUBS 0.007695f
C159 B.n125 VSUBS 0.007695f
C160 B.n126 VSUBS 0.007695f
C161 B.n127 VSUBS 0.007695f
C162 B.n128 VSUBS 0.007695f
C163 B.n129 VSUBS 0.007695f
C164 B.n130 VSUBS 0.007695f
C165 B.n131 VSUBS 0.007695f
C166 B.n132 VSUBS 0.007695f
C167 B.n133 VSUBS 0.007695f
C168 B.n134 VSUBS 0.007695f
C169 B.n135 VSUBS 0.007695f
C170 B.n136 VSUBS 0.007695f
C171 B.n137 VSUBS 0.007695f
C172 B.n138 VSUBS 0.007695f
C173 B.n139 VSUBS 0.007695f
C174 B.n140 VSUBS 0.007695f
C175 B.n141 VSUBS 0.007695f
C176 B.n142 VSUBS 0.007695f
C177 B.n143 VSUBS 0.007695f
C178 B.n144 VSUBS 0.007695f
C179 B.n145 VSUBS 0.007695f
C180 B.n146 VSUBS 0.007695f
C181 B.n147 VSUBS 0.007695f
C182 B.n148 VSUBS 0.007695f
C183 B.n149 VSUBS 0.007695f
C184 B.n150 VSUBS 0.007695f
C185 B.n151 VSUBS 0.007695f
C186 B.n152 VSUBS 0.007695f
C187 B.n153 VSUBS 0.007695f
C188 B.n154 VSUBS 0.007695f
C189 B.n155 VSUBS 0.007695f
C190 B.n156 VSUBS 0.007695f
C191 B.n157 VSUBS 0.007695f
C192 B.n158 VSUBS 0.007695f
C193 B.n159 VSUBS 0.007695f
C194 B.n160 VSUBS 0.007695f
C195 B.n161 VSUBS 0.007695f
C196 B.n162 VSUBS 0.007695f
C197 B.n163 VSUBS 0.007695f
C198 B.n164 VSUBS 0.007695f
C199 B.n165 VSUBS 0.007695f
C200 B.n166 VSUBS 0.007695f
C201 B.n167 VSUBS 0.007695f
C202 B.n168 VSUBS 0.007695f
C203 B.n169 VSUBS 0.007695f
C204 B.n170 VSUBS 0.007695f
C205 B.n171 VSUBS 0.007695f
C206 B.n172 VSUBS 0.007695f
C207 B.n173 VSUBS 0.007695f
C208 B.n174 VSUBS 0.007695f
C209 B.n175 VSUBS 0.007695f
C210 B.n176 VSUBS 0.007695f
C211 B.n177 VSUBS 0.007695f
C212 B.n178 VSUBS 0.007695f
C213 B.n179 VSUBS 0.007695f
C214 B.n180 VSUBS 0.007695f
C215 B.n181 VSUBS 0.007695f
C216 B.n182 VSUBS 0.007695f
C217 B.n183 VSUBS 0.017529f
C218 B.n184 VSUBS 0.007695f
C219 B.n185 VSUBS 0.007695f
C220 B.n186 VSUBS 0.007695f
C221 B.n187 VSUBS 0.007695f
C222 B.n188 VSUBS 0.007695f
C223 B.n189 VSUBS 0.007695f
C224 B.n190 VSUBS 0.007695f
C225 B.n191 VSUBS 0.007695f
C226 B.n192 VSUBS 0.007695f
C227 B.n193 VSUBS 0.007695f
C228 B.n194 VSUBS 0.007695f
C229 B.n195 VSUBS 0.007695f
C230 B.n196 VSUBS 0.007695f
C231 B.n197 VSUBS 0.007695f
C232 B.n198 VSUBS 0.007695f
C233 B.n199 VSUBS 0.007695f
C234 B.n200 VSUBS 0.007695f
C235 B.n201 VSUBS 0.007695f
C236 B.n202 VSUBS 0.007695f
C237 B.n203 VSUBS 0.007695f
C238 B.n204 VSUBS 0.007695f
C239 B.n205 VSUBS 0.007695f
C240 B.n206 VSUBS 0.007695f
C241 B.n207 VSUBS 0.007695f
C242 B.n208 VSUBS 0.007695f
C243 B.n209 VSUBS 0.007695f
C244 B.n210 VSUBS 0.007695f
C245 B.n211 VSUBS 0.007695f
C246 B.n212 VSUBS 0.007695f
C247 B.t5 VSUBS 0.664829f
C248 B.t4 VSUBS 0.693491f
C249 B.t3 VSUBS 3.06798f
C250 B.n213 VSUBS 0.418675f
C251 B.n214 VSUBS 0.083099f
C252 B.n215 VSUBS 0.007695f
C253 B.n216 VSUBS 0.007695f
C254 B.n217 VSUBS 0.007695f
C255 B.n218 VSUBS 0.007695f
C256 B.n219 VSUBS 0.0043f
C257 B.n220 VSUBS 0.007695f
C258 B.n221 VSUBS 0.007695f
C259 B.n222 VSUBS 0.007695f
C260 B.n223 VSUBS 0.007695f
C261 B.n224 VSUBS 0.007695f
C262 B.n225 VSUBS 0.007695f
C263 B.n226 VSUBS 0.007695f
C264 B.n227 VSUBS 0.007695f
C265 B.n228 VSUBS 0.007695f
C266 B.n229 VSUBS 0.007695f
C267 B.n230 VSUBS 0.007695f
C268 B.n231 VSUBS 0.007695f
C269 B.n232 VSUBS 0.007695f
C270 B.n233 VSUBS 0.007695f
C271 B.n234 VSUBS 0.007695f
C272 B.n235 VSUBS 0.007695f
C273 B.n236 VSUBS 0.007695f
C274 B.n237 VSUBS 0.007695f
C275 B.n238 VSUBS 0.007695f
C276 B.n239 VSUBS 0.007695f
C277 B.n240 VSUBS 0.007695f
C278 B.n241 VSUBS 0.007695f
C279 B.n242 VSUBS 0.007695f
C280 B.n243 VSUBS 0.007695f
C281 B.n244 VSUBS 0.007695f
C282 B.n245 VSUBS 0.007695f
C283 B.n246 VSUBS 0.007695f
C284 B.n247 VSUBS 0.007695f
C285 B.n248 VSUBS 0.007695f
C286 B.n249 VSUBS 0.017076f
C287 B.n250 VSUBS 0.007695f
C288 B.n251 VSUBS 0.007695f
C289 B.n252 VSUBS 0.007695f
C290 B.n253 VSUBS 0.007695f
C291 B.n254 VSUBS 0.007695f
C292 B.n255 VSUBS 0.007695f
C293 B.n256 VSUBS 0.007695f
C294 B.n257 VSUBS 0.007695f
C295 B.n258 VSUBS 0.007695f
C296 B.n259 VSUBS 0.007695f
C297 B.n260 VSUBS 0.007695f
C298 B.n261 VSUBS 0.007695f
C299 B.n262 VSUBS 0.007695f
C300 B.n263 VSUBS 0.007695f
C301 B.n264 VSUBS 0.007695f
C302 B.n265 VSUBS 0.007695f
C303 B.n266 VSUBS 0.007695f
C304 B.n267 VSUBS 0.007695f
C305 B.n268 VSUBS 0.007695f
C306 B.n269 VSUBS 0.007695f
C307 B.n270 VSUBS 0.007695f
C308 B.n271 VSUBS 0.007695f
C309 B.n272 VSUBS 0.007695f
C310 B.n273 VSUBS 0.007695f
C311 B.n274 VSUBS 0.007695f
C312 B.n275 VSUBS 0.007695f
C313 B.n276 VSUBS 0.007695f
C314 B.n277 VSUBS 0.007695f
C315 B.n278 VSUBS 0.007695f
C316 B.n279 VSUBS 0.007695f
C317 B.n280 VSUBS 0.007695f
C318 B.n281 VSUBS 0.007695f
C319 B.n282 VSUBS 0.007695f
C320 B.n283 VSUBS 0.007695f
C321 B.n284 VSUBS 0.007695f
C322 B.n285 VSUBS 0.007695f
C323 B.n286 VSUBS 0.007695f
C324 B.n287 VSUBS 0.007695f
C325 B.n288 VSUBS 0.007695f
C326 B.n289 VSUBS 0.007695f
C327 B.n290 VSUBS 0.007695f
C328 B.n291 VSUBS 0.007695f
C329 B.n292 VSUBS 0.007695f
C330 B.n293 VSUBS 0.007695f
C331 B.n294 VSUBS 0.007695f
C332 B.n295 VSUBS 0.007695f
C333 B.n296 VSUBS 0.007695f
C334 B.n297 VSUBS 0.007695f
C335 B.n298 VSUBS 0.007695f
C336 B.n299 VSUBS 0.007695f
C337 B.n300 VSUBS 0.007695f
C338 B.n301 VSUBS 0.007695f
C339 B.n302 VSUBS 0.007695f
C340 B.n303 VSUBS 0.007695f
C341 B.n304 VSUBS 0.007695f
C342 B.n305 VSUBS 0.007695f
C343 B.n306 VSUBS 0.007695f
C344 B.n307 VSUBS 0.007695f
C345 B.n308 VSUBS 0.007695f
C346 B.n309 VSUBS 0.007695f
C347 B.n310 VSUBS 0.007695f
C348 B.n311 VSUBS 0.007695f
C349 B.n312 VSUBS 0.007695f
C350 B.n313 VSUBS 0.007695f
C351 B.n314 VSUBS 0.007695f
C352 B.n315 VSUBS 0.007695f
C353 B.n316 VSUBS 0.007695f
C354 B.n317 VSUBS 0.007695f
C355 B.n318 VSUBS 0.007695f
C356 B.n319 VSUBS 0.007695f
C357 B.n320 VSUBS 0.007695f
C358 B.n321 VSUBS 0.007695f
C359 B.n322 VSUBS 0.007695f
C360 B.n323 VSUBS 0.007695f
C361 B.n324 VSUBS 0.007695f
C362 B.n325 VSUBS 0.007695f
C363 B.n326 VSUBS 0.007695f
C364 B.n327 VSUBS 0.007695f
C365 B.n328 VSUBS 0.007695f
C366 B.n329 VSUBS 0.007695f
C367 B.n330 VSUBS 0.007695f
C368 B.n331 VSUBS 0.007695f
C369 B.n332 VSUBS 0.007695f
C370 B.n333 VSUBS 0.007695f
C371 B.n334 VSUBS 0.007695f
C372 B.n335 VSUBS 0.007695f
C373 B.n336 VSUBS 0.007695f
C374 B.n337 VSUBS 0.007695f
C375 B.n338 VSUBS 0.007695f
C376 B.n339 VSUBS 0.007695f
C377 B.n340 VSUBS 0.007695f
C378 B.n341 VSUBS 0.007695f
C379 B.n342 VSUBS 0.007695f
C380 B.n343 VSUBS 0.007695f
C381 B.n344 VSUBS 0.007695f
C382 B.n345 VSUBS 0.007695f
C383 B.n346 VSUBS 0.007695f
C384 B.n347 VSUBS 0.007695f
C385 B.n348 VSUBS 0.007695f
C386 B.n349 VSUBS 0.007695f
C387 B.n350 VSUBS 0.007695f
C388 B.n351 VSUBS 0.007695f
C389 B.n352 VSUBS 0.007695f
C390 B.n353 VSUBS 0.007695f
C391 B.n354 VSUBS 0.007695f
C392 B.n355 VSUBS 0.007695f
C393 B.n356 VSUBS 0.007695f
C394 B.n357 VSUBS 0.007695f
C395 B.n358 VSUBS 0.007695f
C396 B.n359 VSUBS 0.007695f
C397 B.n360 VSUBS 0.007695f
C398 B.n361 VSUBS 0.007695f
C399 B.n362 VSUBS 0.007695f
C400 B.n363 VSUBS 0.007695f
C401 B.n364 VSUBS 0.007695f
C402 B.n365 VSUBS 0.007695f
C403 B.n366 VSUBS 0.007695f
C404 B.n367 VSUBS 0.007695f
C405 B.n368 VSUBS 0.007695f
C406 B.n369 VSUBS 0.007695f
C407 B.n370 VSUBS 0.007695f
C408 B.n371 VSUBS 0.007695f
C409 B.n372 VSUBS 0.007695f
C410 B.n373 VSUBS 0.007695f
C411 B.n374 VSUBS 0.007695f
C412 B.n375 VSUBS 0.007695f
C413 B.n376 VSUBS 0.007695f
C414 B.n377 VSUBS 0.007695f
C415 B.n378 VSUBS 0.007695f
C416 B.n379 VSUBS 0.007695f
C417 B.n380 VSUBS 0.007695f
C418 B.n381 VSUBS 0.007695f
C419 B.n382 VSUBS 0.007695f
C420 B.n383 VSUBS 0.007695f
C421 B.n384 VSUBS 0.007695f
C422 B.n385 VSUBS 0.007695f
C423 B.n386 VSUBS 0.007695f
C424 B.n387 VSUBS 0.007695f
C425 B.n388 VSUBS 0.007695f
C426 B.n389 VSUBS 0.007695f
C427 B.n390 VSUBS 0.007695f
C428 B.n391 VSUBS 0.007695f
C429 B.n392 VSUBS 0.007695f
C430 B.n393 VSUBS 0.007695f
C431 B.n394 VSUBS 0.017076f
C432 B.n395 VSUBS 0.018457f
C433 B.n396 VSUBS 0.018457f
C434 B.n397 VSUBS 0.007695f
C435 B.n398 VSUBS 0.007695f
C436 B.n399 VSUBS 0.007695f
C437 B.n400 VSUBS 0.007695f
C438 B.n401 VSUBS 0.007695f
C439 B.n402 VSUBS 0.007695f
C440 B.n403 VSUBS 0.007695f
C441 B.n404 VSUBS 0.007695f
C442 B.n405 VSUBS 0.007695f
C443 B.n406 VSUBS 0.007695f
C444 B.n407 VSUBS 0.007695f
C445 B.n408 VSUBS 0.007695f
C446 B.n409 VSUBS 0.007695f
C447 B.n410 VSUBS 0.007695f
C448 B.n411 VSUBS 0.007695f
C449 B.n412 VSUBS 0.007695f
C450 B.n413 VSUBS 0.007695f
C451 B.n414 VSUBS 0.007695f
C452 B.n415 VSUBS 0.007695f
C453 B.n416 VSUBS 0.007695f
C454 B.n417 VSUBS 0.007695f
C455 B.n418 VSUBS 0.007695f
C456 B.n419 VSUBS 0.007695f
C457 B.n420 VSUBS 0.007695f
C458 B.n421 VSUBS 0.007695f
C459 B.n422 VSUBS 0.007695f
C460 B.n423 VSUBS 0.007695f
C461 B.n424 VSUBS 0.007695f
C462 B.n425 VSUBS 0.007695f
C463 B.n426 VSUBS 0.007695f
C464 B.n427 VSUBS 0.007695f
C465 B.n428 VSUBS 0.007695f
C466 B.n429 VSUBS 0.007695f
C467 B.n430 VSUBS 0.007695f
C468 B.n431 VSUBS 0.007695f
C469 B.n432 VSUBS 0.007695f
C470 B.n433 VSUBS 0.007695f
C471 B.n434 VSUBS 0.007695f
C472 B.n435 VSUBS 0.007695f
C473 B.n436 VSUBS 0.007695f
C474 B.n437 VSUBS 0.007695f
C475 B.n438 VSUBS 0.007695f
C476 B.n439 VSUBS 0.007695f
C477 B.n440 VSUBS 0.007695f
C478 B.n441 VSUBS 0.007695f
C479 B.n442 VSUBS 0.007695f
C480 B.n443 VSUBS 0.007695f
C481 B.n444 VSUBS 0.007695f
C482 B.n445 VSUBS 0.007695f
C483 B.n446 VSUBS 0.007695f
C484 B.n447 VSUBS 0.007695f
C485 B.n448 VSUBS 0.007695f
C486 B.n449 VSUBS 0.007695f
C487 B.n450 VSUBS 0.007695f
C488 B.n451 VSUBS 0.007695f
C489 B.n452 VSUBS 0.007695f
C490 B.n453 VSUBS 0.007695f
C491 B.n454 VSUBS 0.007695f
C492 B.n455 VSUBS 0.007695f
C493 B.n456 VSUBS 0.007695f
C494 B.n457 VSUBS 0.007695f
C495 B.n458 VSUBS 0.007695f
C496 B.n459 VSUBS 0.007695f
C497 B.n460 VSUBS 0.007695f
C498 B.n461 VSUBS 0.007695f
C499 B.n462 VSUBS 0.007695f
C500 B.n463 VSUBS 0.007695f
C501 B.n464 VSUBS 0.007695f
C502 B.n465 VSUBS 0.007695f
C503 B.n466 VSUBS 0.007695f
C504 B.n467 VSUBS 0.007695f
C505 B.n468 VSUBS 0.007695f
C506 B.n469 VSUBS 0.007695f
C507 B.n470 VSUBS 0.007695f
C508 B.n471 VSUBS 0.007695f
C509 B.n472 VSUBS 0.007695f
C510 B.n473 VSUBS 0.007695f
C511 B.n474 VSUBS 0.007695f
C512 B.n475 VSUBS 0.007695f
C513 B.n476 VSUBS 0.007695f
C514 B.n477 VSUBS 0.007695f
C515 B.n478 VSUBS 0.007695f
C516 B.n479 VSUBS 0.007695f
C517 B.n480 VSUBS 0.007695f
C518 B.n481 VSUBS 0.007695f
C519 B.t11 VSUBS 0.664853f
C520 B.t10 VSUBS 0.693509f
C521 B.t9 VSUBS 3.06798f
C522 B.n482 VSUBS 0.418657f
C523 B.n483 VSUBS 0.083075f
C524 B.n484 VSUBS 0.017828f
C525 B.n485 VSUBS 0.007242f
C526 B.n486 VSUBS 0.007695f
C527 B.n487 VSUBS 0.007695f
C528 B.n488 VSUBS 0.007695f
C529 B.n489 VSUBS 0.007695f
C530 B.n490 VSUBS 0.007695f
C531 B.n491 VSUBS 0.007695f
C532 B.n492 VSUBS 0.007695f
C533 B.n493 VSUBS 0.007695f
C534 B.n494 VSUBS 0.007695f
C535 B.n495 VSUBS 0.007695f
C536 B.n496 VSUBS 0.007695f
C537 B.n497 VSUBS 0.007695f
C538 B.n498 VSUBS 0.007695f
C539 B.n499 VSUBS 0.007695f
C540 B.n500 VSUBS 0.007695f
C541 B.n501 VSUBS 0.0043f
C542 B.n502 VSUBS 0.017828f
C543 B.n503 VSUBS 0.007242f
C544 B.n504 VSUBS 0.007695f
C545 B.n505 VSUBS 0.007695f
C546 B.n506 VSUBS 0.007695f
C547 B.n507 VSUBS 0.007695f
C548 B.n508 VSUBS 0.007695f
C549 B.n509 VSUBS 0.007695f
C550 B.n510 VSUBS 0.007695f
C551 B.n511 VSUBS 0.007695f
C552 B.n512 VSUBS 0.007695f
C553 B.n513 VSUBS 0.007695f
C554 B.n514 VSUBS 0.007695f
C555 B.n515 VSUBS 0.007695f
C556 B.n516 VSUBS 0.007695f
C557 B.n517 VSUBS 0.007695f
C558 B.n518 VSUBS 0.007695f
C559 B.n519 VSUBS 0.007695f
C560 B.n520 VSUBS 0.007695f
C561 B.n521 VSUBS 0.007695f
C562 B.n522 VSUBS 0.007695f
C563 B.n523 VSUBS 0.007695f
C564 B.n524 VSUBS 0.007695f
C565 B.n525 VSUBS 0.007695f
C566 B.n526 VSUBS 0.007695f
C567 B.n527 VSUBS 0.007695f
C568 B.n528 VSUBS 0.007695f
C569 B.n529 VSUBS 0.007695f
C570 B.n530 VSUBS 0.007695f
C571 B.n531 VSUBS 0.007695f
C572 B.n532 VSUBS 0.007695f
C573 B.n533 VSUBS 0.007695f
C574 B.n534 VSUBS 0.007695f
C575 B.n535 VSUBS 0.007695f
C576 B.n536 VSUBS 0.007695f
C577 B.n537 VSUBS 0.007695f
C578 B.n538 VSUBS 0.007695f
C579 B.n539 VSUBS 0.007695f
C580 B.n540 VSUBS 0.007695f
C581 B.n541 VSUBS 0.007695f
C582 B.n542 VSUBS 0.007695f
C583 B.n543 VSUBS 0.007695f
C584 B.n544 VSUBS 0.007695f
C585 B.n545 VSUBS 0.007695f
C586 B.n546 VSUBS 0.007695f
C587 B.n547 VSUBS 0.007695f
C588 B.n548 VSUBS 0.007695f
C589 B.n549 VSUBS 0.007695f
C590 B.n550 VSUBS 0.007695f
C591 B.n551 VSUBS 0.007695f
C592 B.n552 VSUBS 0.007695f
C593 B.n553 VSUBS 0.007695f
C594 B.n554 VSUBS 0.007695f
C595 B.n555 VSUBS 0.007695f
C596 B.n556 VSUBS 0.007695f
C597 B.n557 VSUBS 0.007695f
C598 B.n558 VSUBS 0.007695f
C599 B.n559 VSUBS 0.007695f
C600 B.n560 VSUBS 0.007695f
C601 B.n561 VSUBS 0.007695f
C602 B.n562 VSUBS 0.007695f
C603 B.n563 VSUBS 0.007695f
C604 B.n564 VSUBS 0.007695f
C605 B.n565 VSUBS 0.007695f
C606 B.n566 VSUBS 0.007695f
C607 B.n567 VSUBS 0.007695f
C608 B.n568 VSUBS 0.007695f
C609 B.n569 VSUBS 0.007695f
C610 B.n570 VSUBS 0.007695f
C611 B.n571 VSUBS 0.007695f
C612 B.n572 VSUBS 0.007695f
C613 B.n573 VSUBS 0.007695f
C614 B.n574 VSUBS 0.007695f
C615 B.n575 VSUBS 0.007695f
C616 B.n576 VSUBS 0.007695f
C617 B.n577 VSUBS 0.007695f
C618 B.n578 VSUBS 0.007695f
C619 B.n579 VSUBS 0.007695f
C620 B.n580 VSUBS 0.007695f
C621 B.n581 VSUBS 0.007695f
C622 B.n582 VSUBS 0.007695f
C623 B.n583 VSUBS 0.007695f
C624 B.n584 VSUBS 0.007695f
C625 B.n585 VSUBS 0.007695f
C626 B.n586 VSUBS 0.007695f
C627 B.n587 VSUBS 0.007695f
C628 B.n588 VSUBS 0.007695f
C629 B.n589 VSUBS 0.007695f
C630 B.n590 VSUBS 0.018457f
C631 B.n591 VSUBS 0.017076f
C632 B.n592 VSUBS 0.018004f
C633 B.n593 VSUBS 0.007695f
C634 B.n594 VSUBS 0.007695f
C635 B.n595 VSUBS 0.007695f
C636 B.n596 VSUBS 0.007695f
C637 B.n597 VSUBS 0.007695f
C638 B.n598 VSUBS 0.007695f
C639 B.n599 VSUBS 0.007695f
C640 B.n600 VSUBS 0.007695f
C641 B.n601 VSUBS 0.007695f
C642 B.n602 VSUBS 0.007695f
C643 B.n603 VSUBS 0.007695f
C644 B.n604 VSUBS 0.007695f
C645 B.n605 VSUBS 0.007695f
C646 B.n606 VSUBS 0.007695f
C647 B.n607 VSUBS 0.007695f
C648 B.n608 VSUBS 0.007695f
C649 B.n609 VSUBS 0.007695f
C650 B.n610 VSUBS 0.007695f
C651 B.n611 VSUBS 0.007695f
C652 B.n612 VSUBS 0.007695f
C653 B.n613 VSUBS 0.007695f
C654 B.n614 VSUBS 0.007695f
C655 B.n615 VSUBS 0.007695f
C656 B.n616 VSUBS 0.007695f
C657 B.n617 VSUBS 0.007695f
C658 B.n618 VSUBS 0.007695f
C659 B.n619 VSUBS 0.007695f
C660 B.n620 VSUBS 0.007695f
C661 B.n621 VSUBS 0.007695f
C662 B.n622 VSUBS 0.007695f
C663 B.n623 VSUBS 0.007695f
C664 B.n624 VSUBS 0.007695f
C665 B.n625 VSUBS 0.007695f
C666 B.n626 VSUBS 0.007695f
C667 B.n627 VSUBS 0.007695f
C668 B.n628 VSUBS 0.007695f
C669 B.n629 VSUBS 0.007695f
C670 B.n630 VSUBS 0.007695f
C671 B.n631 VSUBS 0.007695f
C672 B.n632 VSUBS 0.007695f
C673 B.n633 VSUBS 0.007695f
C674 B.n634 VSUBS 0.007695f
C675 B.n635 VSUBS 0.007695f
C676 B.n636 VSUBS 0.007695f
C677 B.n637 VSUBS 0.007695f
C678 B.n638 VSUBS 0.007695f
C679 B.n639 VSUBS 0.007695f
C680 B.n640 VSUBS 0.007695f
C681 B.n641 VSUBS 0.007695f
C682 B.n642 VSUBS 0.007695f
C683 B.n643 VSUBS 0.007695f
C684 B.n644 VSUBS 0.007695f
C685 B.n645 VSUBS 0.007695f
C686 B.n646 VSUBS 0.007695f
C687 B.n647 VSUBS 0.007695f
C688 B.n648 VSUBS 0.007695f
C689 B.n649 VSUBS 0.007695f
C690 B.n650 VSUBS 0.007695f
C691 B.n651 VSUBS 0.007695f
C692 B.n652 VSUBS 0.007695f
C693 B.n653 VSUBS 0.007695f
C694 B.n654 VSUBS 0.007695f
C695 B.n655 VSUBS 0.007695f
C696 B.n656 VSUBS 0.007695f
C697 B.n657 VSUBS 0.007695f
C698 B.n658 VSUBS 0.007695f
C699 B.n659 VSUBS 0.007695f
C700 B.n660 VSUBS 0.007695f
C701 B.n661 VSUBS 0.007695f
C702 B.n662 VSUBS 0.007695f
C703 B.n663 VSUBS 0.007695f
C704 B.n664 VSUBS 0.007695f
C705 B.n665 VSUBS 0.007695f
C706 B.n666 VSUBS 0.007695f
C707 B.n667 VSUBS 0.007695f
C708 B.n668 VSUBS 0.007695f
C709 B.n669 VSUBS 0.007695f
C710 B.n670 VSUBS 0.007695f
C711 B.n671 VSUBS 0.007695f
C712 B.n672 VSUBS 0.007695f
C713 B.n673 VSUBS 0.007695f
C714 B.n674 VSUBS 0.007695f
C715 B.n675 VSUBS 0.007695f
C716 B.n676 VSUBS 0.007695f
C717 B.n677 VSUBS 0.007695f
C718 B.n678 VSUBS 0.007695f
C719 B.n679 VSUBS 0.007695f
C720 B.n680 VSUBS 0.007695f
C721 B.n681 VSUBS 0.007695f
C722 B.n682 VSUBS 0.007695f
C723 B.n683 VSUBS 0.007695f
C724 B.n684 VSUBS 0.007695f
C725 B.n685 VSUBS 0.007695f
C726 B.n686 VSUBS 0.007695f
C727 B.n687 VSUBS 0.007695f
C728 B.n688 VSUBS 0.007695f
C729 B.n689 VSUBS 0.007695f
C730 B.n690 VSUBS 0.007695f
C731 B.n691 VSUBS 0.007695f
C732 B.n692 VSUBS 0.007695f
C733 B.n693 VSUBS 0.007695f
C734 B.n694 VSUBS 0.007695f
C735 B.n695 VSUBS 0.007695f
C736 B.n696 VSUBS 0.007695f
C737 B.n697 VSUBS 0.007695f
C738 B.n698 VSUBS 0.007695f
C739 B.n699 VSUBS 0.007695f
C740 B.n700 VSUBS 0.007695f
C741 B.n701 VSUBS 0.007695f
C742 B.n702 VSUBS 0.007695f
C743 B.n703 VSUBS 0.007695f
C744 B.n704 VSUBS 0.007695f
C745 B.n705 VSUBS 0.007695f
C746 B.n706 VSUBS 0.007695f
C747 B.n707 VSUBS 0.007695f
C748 B.n708 VSUBS 0.007695f
C749 B.n709 VSUBS 0.007695f
C750 B.n710 VSUBS 0.007695f
C751 B.n711 VSUBS 0.007695f
C752 B.n712 VSUBS 0.007695f
C753 B.n713 VSUBS 0.007695f
C754 B.n714 VSUBS 0.007695f
C755 B.n715 VSUBS 0.007695f
C756 B.n716 VSUBS 0.007695f
C757 B.n717 VSUBS 0.007695f
C758 B.n718 VSUBS 0.007695f
C759 B.n719 VSUBS 0.007695f
C760 B.n720 VSUBS 0.007695f
C761 B.n721 VSUBS 0.007695f
C762 B.n722 VSUBS 0.007695f
C763 B.n723 VSUBS 0.007695f
C764 B.n724 VSUBS 0.007695f
C765 B.n725 VSUBS 0.007695f
C766 B.n726 VSUBS 0.007695f
C767 B.n727 VSUBS 0.007695f
C768 B.n728 VSUBS 0.007695f
C769 B.n729 VSUBS 0.007695f
C770 B.n730 VSUBS 0.007695f
C771 B.n731 VSUBS 0.007695f
C772 B.n732 VSUBS 0.007695f
C773 B.n733 VSUBS 0.007695f
C774 B.n734 VSUBS 0.007695f
C775 B.n735 VSUBS 0.007695f
C776 B.n736 VSUBS 0.007695f
C777 B.n737 VSUBS 0.007695f
C778 B.n738 VSUBS 0.007695f
C779 B.n739 VSUBS 0.007695f
C780 B.n740 VSUBS 0.007695f
C781 B.n741 VSUBS 0.007695f
C782 B.n742 VSUBS 0.007695f
C783 B.n743 VSUBS 0.007695f
C784 B.n744 VSUBS 0.007695f
C785 B.n745 VSUBS 0.007695f
C786 B.n746 VSUBS 0.007695f
C787 B.n747 VSUBS 0.007695f
C788 B.n748 VSUBS 0.007695f
C789 B.n749 VSUBS 0.007695f
C790 B.n750 VSUBS 0.007695f
C791 B.n751 VSUBS 0.007695f
C792 B.n752 VSUBS 0.007695f
C793 B.n753 VSUBS 0.007695f
C794 B.n754 VSUBS 0.007695f
C795 B.n755 VSUBS 0.007695f
C796 B.n756 VSUBS 0.007695f
C797 B.n757 VSUBS 0.007695f
C798 B.n758 VSUBS 0.007695f
C799 B.n759 VSUBS 0.007695f
C800 B.n760 VSUBS 0.007695f
C801 B.n761 VSUBS 0.007695f
C802 B.n762 VSUBS 0.007695f
C803 B.n763 VSUBS 0.007695f
C804 B.n764 VSUBS 0.007695f
C805 B.n765 VSUBS 0.007695f
C806 B.n766 VSUBS 0.007695f
C807 B.n767 VSUBS 0.007695f
C808 B.n768 VSUBS 0.007695f
C809 B.n769 VSUBS 0.007695f
C810 B.n770 VSUBS 0.007695f
C811 B.n771 VSUBS 0.007695f
C812 B.n772 VSUBS 0.007695f
C813 B.n773 VSUBS 0.007695f
C814 B.n774 VSUBS 0.007695f
C815 B.n775 VSUBS 0.007695f
C816 B.n776 VSUBS 0.007695f
C817 B.n777 VSUBS 0.007695f
C818 B.n778 VSUBS 0.007695f
C819 B.n779 VSUBS 0.007695f
C820 B.n780 VSUBS 0.007695f
C821 B.n781 VSUBS 0.007695f
C822 B.n782 VSUBS 0.007695f
C823 B.n783 VSUBS 0.007695f
C824 B.n784 VSUBS 0.007695f
C825 B.n785 VSUBS 0.007695f
C826 B.n786 VSUBS 0.007695f
C827 B.n787 VSUBS 0.007695f
C828 B.n788 VSUBS 0.007695f
C829 B.n789 VSUBS 0.007695f
C830 B.n790 VSUBS 0.007695f
C831 B.n791 VSUBS 0.007695f
C832 B.n792 VSUBS 0.007695f
C833 B.n793 VSUBS 0.007695f
C834 B.n794 VSUBS 0.007695f
C835 B.n795 VSUBS 0.007695f
C836 B.n796 VSUBS 0.007695f
C837 B.n797 VSUBS 0.007695f
C838 B.n798 VSUBS 0.007695f
C839 B.n799 VSUBS 0.007695f
C840 B.n800 VSUBS 0.007695f
C841 B.n801 VSUBS 0.007695f
C842 B.n802 VSUBS 0.007695f
C843 B.n803 VSUBS 0.007695f
C844 B.n804 VSUBS 0.007695f
C845 B.n805 VSUBS 0.007695f
C846 B.n806 VSUBS 0.007695f
C847 B.n807 VSUBS 0.007695f
C848 B.n808 VSUBS 0.007695f
C849 B.n809 VSUBS 0.007695f
C850 B.n810 VSUBS 0.007695f
C851 B.n811 VSUBS 0.007695f
C852 B.n812 VSUBS 0.007695f
C853 B.n813 VSUBS 0.007695f
C854 B.n814 VSUBS 0.007695f
C855 B.n815 VSUBS 0.017076f
C856 B.n816 VSUBS 0.018457f
C857 B.n817 VSUBS 0.018457f
C858 B.n818 VSUBS 0.007695f
C859 B.n819 VSUBS 0.007695f
C860 B.n820 VSUBS 0.007695f
C861 B.n821 VSUBS 0.007695f
C862 B.n822 VSUBS 0.007695f
C863 B.n823 VSUBS 0.007695f
C864 B.n824 VSUBS 0.007695f
C865 B.n825 VSUBS 0.007695f
C866 B.n826 VSUBS 0.007695f
C867 B.n827 VSUBS 0.007695f
C868 B.n828 VSUBS 0.007695f
C869 B.n829 VSUBS 0.007695f
C870 B.n830 VSUBS 0.007695f
C871 B.n831 VSUBS 0.007695f
C872 B.n832 VSUBS 0.007695f
C873 B.n833 VSUBS 0.007695f
C874 B.n834 VSUBS 0.007695f
C875 B.n835 VSUBS 0.007695f
C876 B.n836 VSUBS 0.007695f
C877 B.n837 VSUBS 0.007695f
C878 B.n838 VSUBS 0.007695f
C879 B.n839 VSUBS 0.007695f
C880 B.n840 VSUBS 0.007695f
C881 B.n841 VSUBS 0.007695f
C882 B.n842 VSUBS 0.007695f
C883 B.n843 VSUBS 0.007695f
C884 B.n844 VSUBS 0.007695f
C885 B.n845 VSUBS 0.007695f
C886 B.n846 VSUBS 0.007695f
C887 B.n847 VSUBS 0.007695f
C888 B.n848 VSUBS 0.007695f
C889 B.n849 VSUBS 0.007695f
C890 B.n850 VSUBS 0.007695f
C891 B.n851 VSUBS 0.007695f
C892 B.n852 VSUBS 0.007695f
C893 B.n853 VSUBS 0.007695f
C894 B.n854 VSUBS 0.007695f
C895 B.n855 VSUBS 0.007695f
C896 B.n856 VSUBS 0.007695f
C897 B.n857 VSUBS 0.007695f
C898 B.n858 VSUBS 0.007695f
C899 B.n859 VSUBS 0.007695f
C900 B.n860 VSUBS 0.007695f
C901 B.n861 VSUBS 0.007695f
C902 B.n862 VSUBS 0.007695f
C903 B.n863 VSUBS 0.007695f
C904 B.n864 VSUBS 0.007695f
C905 B.n865 VSUBS 0.007695f
C906 B.n866 VSUBS 0.007695f
C907 B.n867 VSUBS 0.007695f
C908 B.n868 VSUBS 0.007695f
C909 B.n869 VSUBS 0.007695f
C910 B.n870 VSUBS 0.007695f
C911 B.n871 VSUBS 0.007695f
C912 B.n872 VSUBS 0.007695f
C913 B.n873 VSUBS 0.007695f
C914 B.n874 VSUBS 0.007695f
C915 B.n875 VSUBS 0.007695f
C916 B.n876 VSUBS 0.007695f
C917 B.n877 VSUBS 0.007695f
C918 B.n878 VSUBS 0.007695f
C919 B.n879 VSUBS 0.007695f
C920 B.n880 VSUBS 0.007695f
C921 B.n881 VSUBS 0.007695f
C922 B.n882 VSUBS 0.007695f
C923 B.n883 VSUBS 0.007695f
C924 B.n884 VSUBS 0.007695f
C925 B.n885 VSUBS 0.007695f
C926 B.n886 VSUBS 0.007695f
C927 B.n887 VSUBS 0.007695f
C928 B.n888 VSUBS 0.007695f
C929 B.n889 VSUBS 0.007695f
C930 B.n890 VSUBS 0.007695f
C931 B.n891 VSUBS 0.007695f
C932 B.n892 VSUBS 0.007695f
C933 B.n893 VSUBS 0.007695f
C934 B.n894 VSUBS 0.007695f
C935 B.n895 VSUBS 0.007695f
C936 B.n896 VSUBS 0.007695f
C937 B.n897 VSUBS 0.007695f
C938 B.n898 VSUBS 0.007695f
C939 B.n899 VSUBS 0.007695f
C940 B.n900 VSUBS 0.007695f
C941 B.n901 VSUBS 0.007695f
C942 B.n902 VSUBS 0.007695f
C943 B.n903 VSUBS 0.007695f
C944 B.n904 VSUBS 0.007242f
C945 B.n905 VSUBS 0.017828f
C946 B.n906 VSUBS 0.0043f
C947 B.n907 VSUBS 0.007695f
C948 B.n908 VSUBS 0.007695f
C949 B.n909 VSUBS 0.007695f
C950 B.n910 VSUBS 0.007695f
C951 B.n911 VSUBS 0.007695f
C952 B.n912 VSUBS 0.007695f
C953 B.n913 VSUBS 0.007695f
C954 B.n914 VSUBS 0.007695f
C955 B.n915 VSUBS 0.007695f
C956 B.n916 VSUBS 0.007695f
C957 B.n917 VSUBS 0.007695f
C958 B.n918 VSUBS 0.007695f
C959 B.n919 VSUBS 0.0043f
C960 B.n920 VSUBS 0.007695f
C961 B.n921 VSUBS 0.007695f
C962 B.n922 VSUBS 0.007695f
C963 B.n923 VSUBS 0.007695f
C964 B.n924 VSUBS 0.007695f
C965 B.n925 VSUBS 0.007695f
C966 B.n926 VSUBS 0.007695f
C967 B.n927 VSUBS 0.007695f
C968 B.n928 VSUBS 0.007695f
C969 B.n929 VSUBS 0.007695f
C970 B.n930 VSUBS 0.007695f
C971 B.n931 VSUBS 0.007695f
C972 B.n932 VSUBS 0.007695f
C973 B.n933 VSUBS 0.007695f
C974 B.n934 VSUBS 0.007695f
C975 B.n935 VSUBS 0.007695f
C976 B.n936 VSUBS 0.007695f
C977 B.n937 VSUBS 0.007695f
C978 B.n938 VSUBS 0.007695f
C979 B.n939 VSUBS 0.007695f
C980 B.n940 VSUBS 0.007695f
C981 B.n941 VSUBS 0.007695f
C982 B.n942 VSUBS 0.007695f
C983 B.n943 VSUBS 0.007695f
C984 B.n944 VSUBS 0.007695f
C985 B.n945 VSUBS 0.007695f
C986 B.n946 VSUBS 0.007695f
C987 B.n947 VSUBS 0.007695f
C988 B.n948 VSUBS 0.007695f
C989 B.n949 VSUBS 0.007695f
C990 B.n950 VSUBS 0.007695f
C991 B.n951 VSUBS 0.007695f
C992 B.n952 VSUBS 0.007695f
C993 B.n953 VSUBS 0.007695f
C994 B.n954 VSUBS 0.007695f
C995 B.n955 VSUBS 0.007695f
C996 B.n956 VSUBS 0.007695f
C997 B.n957 VSUBS 0.007695f
C998 B.n958 VSUBS 0.007695f
C999 B.n959 VSUBS 0.007695f
C1000 B.n960 VSUBS 0.007695f
C1001 B.n961 VSUBS 0.007695f
C1002 B.n962 VSUBS 0.007695f
C1003 B.n963 VSUBS 0.007695f
C1004 B.n964 VSUBS 0.007695f
C1005 B.n965 VSUBS 0.007695f
C1006 B.n966 VSUBS 0.007695f
C1007 B.n967 VSUBS 0.007695f
C1008 B.n968 VSUBS 0.007695f
C1009 B.n969 VSUBS 0.007695f
C1010 B.n970 VSUBS 0.007695f
C1011 B.n971 VSUBS 0.007695f
C1012 B.n972 VSUBS 0.007695f
C1013 B.n973 VSUBS 0.007695f
C1014 B.n974 VSUBS 0.007695f
C1015 B.n975 VSUBS 0.007695f
C1016 B.n976 VSUBS 0.007695f
C1017 B.n977 VSUBS 0.007695f
C1018 B.n978 VSUBS 0.007695f
C1019 B.n979 VSUBS 0.007695f
C1020 B.n980 VSUBS 0.007695f
C1021 B.n981 VSUBS 0.007695f
C1022 B.n982 VSUBS 0.007695f
C1023 B.n983 VSUBS 0.007695f
C1024 B.n984 VSUBS 0.007695f
C1025 B.n985 VSUBS 0.007695f
C1026 B.n986 VSUBS 0.007695f
C1027 B.n987 VSUBS 0.007695f
C1028 B.n988 VSUBS 0.007695f
C1029 B.n989 VSUBS 0.007695f
C1030 B.n990 VSUBS 0.007695f
C1031 B.n991 VSUBS 0.007695f
C1032 B.n992 VSUBS 0.007695f
C1033 B.n993 VSUBS 0.007695f
C1034 B.n994 VSUBS 0.007695f
C1035 B.n995 VSUBS 0.007695f
C1036 B.n996 VSUBS 0.007695f
C1037 B.n997 VSUBS 0.007695f
C1038 B.n998 VSUBS 0.007695f
C1039 B.n999 VSUBS 0.007695f
C1040 B.n1000 VSUBS 0.007695f
C1041 B.n1001 VSUBS 0.007695f
C1042 B.n1002 VSUBS 0.007695f
C1043 B.n1003 VSUBS 0.007695f
C1044 B.n1004 VSUBS 0.007695f
C1045 B.n1005 VSUBS 0.007695f
C1046 B.n1006 VSUBS 0.007695f
C1047 B.n1007 VSUBS 0.007695f
C1048 B.n1008 VSUBS 0.018457f
C1049 B.n1009 VSUBS 0.017076f
C1050 B.n1010 VSUBS 0.017076f
C1051 B.n1011 VSUBS 0.007695f
C1052 B.n1012 VSUBS 0.007695f
C1053 B.n1013 VSUBS 0.007695f
C1054 B.n1014 VSUBS 0.007695f
C1055 B.n1015 VSUBS 0.007695f
C1056 B.n1016 VSUBS 0.007695f
C1057 B.n1017 VSUBS 0.007695f
C1058 B.n1018 VSUBS 0.007695f
C1059 B.n1019 VSUBS 0.007695f
C1060 B.n1020 VSUBS 0.007695f
C1061 B.n1021 VSUBS 0.007695f
C1062 B.n1022 VSUBS 0.007695f
C1063 B.n1023 VSUBS 0.007695f
C1064 B.n1024 VSUBS 0.007695f
C1065 B.n1025 VSUBS 0.007695f
C1066 B.n1026 VSUBS 0.007695f
C1067 B.n1027 VSUBS 0.007695f
C1068 B.n1028 VSUBS 0.007695f
C1069 B.n1029 VSUBS 0.007695f
C1070 B.n1030 VSUBS 0.007695f
C1071 B.n1031 VSUBS 0.007695f
C1072 B.n1032 VSUBS 0.007695f
C1073 B.n1033 VSUBS 0.007695f
C1074 B.n1034 VSUBS 0.007695f
C1075 B.n1035 VSUBS 0.007695f
C1076 B.n1036 VSUBS 0.007695f
C1077 B.n1037 VSUBS 0.007695f
C1078 B.n1038 VSUBS 0.007695f
C1079 B.n1039 VSUBS 0.007695f
C1080 B.n1040 VSUBS 0.007695f
C1081 B.n1041 VSUBS 0.007695f
C1082 B.n1042 VSUBS 0.007695f
C1083 B.n1043 VSUBS 0.007695f
C1084 B.n1044 VSUBS 0.007695f
C1085 B.n1045 VSUBS 0.007695f
C1086 B.n1046 VSUBS 0.007695f
C1087 B.n1047 VSUBS 0.007695f
C1088 B.n1048 VSUBS 0.007695f
C1089 B.n1049 VSUBS 0.007695f
C1090 B.n1050 VSUBS 0.007695f
C1091 B.n1051 VSUBS 0.007695f
C1092 B.n1052 VSUBS 0.007695f
C1093 B.n1053 VSUBS 0.007695f
C1094 B.n1054 VSUBS 0.007695f
C1095 B.n1055 VSUBS 0.007695f
C1096 B.n1056 VSUBS 0.007695f
C1097 B.n1057 VSUBS 0.007695f
C1098 B.n1058 VSUBS 0.007695f
C1099 B.n1059 VSUBS 0.007695f
C1100 B.n1060 VSUBS 0.007695f
C1101 B.n1061 VSUBS 0.007695f
C1102 B.n1062 VSUBS 0.007695f
C1103 B.n1063 VSUBS 0.007695f
C1104 B.n1064 VSUBS 0.007695f
C1105 B.n1065 VSUBS 0.007695f
C1106 B.n1066 VSUBS 0.007695f
C1107 B.n1067 VSUBS 0.007695f
C1108 B.n1068 VSUBS 0.007695f
C1109 B.n1069 VSUBS 0.007695f
C1110 B.n1070 VSUBS 0.007695f
C1111 B.n1071 VSUBS 0.007695f
C1112 B.n1072 VSUBS 0.007695f
C1113 B.n1073 VSUBS 0.007695f
C1114 B.n1074 VSUBS 0.007695f
C1115 B.n1075 VSUBS 0.007695f
C1116 B.n1076 VSUBS 0.007695f
C1117 B.n1077 VSUBS 0.007695f
C1118 B.n1078 VSUBS 0.007695f
C1119 B.n1079 VSUBS 0.007695f
C1120 B.n1080 VSUBS 0.007695f
C1121 B.n1081 VSUBS 0.007695f
C1122 B.n1082 VSUBS 0.007695f
C1123 B.n1083 VSUBS 0.007695f
C1124 B.n1084 VSUBS 0.007695f
C1125 B.n1085 VSUBS 0.007695f
C1126 B.n1086 VSUBS 0.007695f
C1127 B.n1087 VSUBS 0.007695f
C1128 B.n1088 VSUBS 0.007695f
C1129 B.n1089 VSUBS 0.007695f
C1130 B.n1090 VSUBS 0.007695f
C1131 B.n1091 VSUBS 0.007695f
C1132 B.n1092 VSUBS 0.007695f
C1133 B.n1093 VSUBS 0.007695f
C1134 B.n1094 VSUBS 0.007695f
C1135 B.n1095 VSUBS 0.007695f
C1136 B.n1096 VSUBS 0.007695f
C1137 B.n1097 VSUBS 0.007695f
C1138 B.n1098 VSUBS 0.007695f
C1139 B.n1099 VSUBS 0.007695f
C1140 B.n1100 VSUBS 0.007695f
C1141 B.n1101 VSUBS 0.007695f
C1142 B.n1102 VSUBS 0.007695f
C1143 B.n1103 VSUBS 0.007695f
C1144 B.n1104 VSUBS 0.007695f
C1145 B.n1105 VSUBS 0.007695f
C1146 B.n1106 VSUBS 0.007695f
C1147 B.n1107 VSUBS 0.007695f
C1148 B.n1108 VSUBS 0.007695f
C1149 B.n1109 VSUBS 0.007695f
C1150 B.n1110 VSUBS 0.007695f
C1151 B.n1111 VSUBS 0.007695f
C1152 B.n1112 VSUBS 0.007695f
C1153 B.n1113 VSUBS 0.007695f
C1154 B.n1114 VSUBS 0.007695f
C1155 B.n1115 VSUBS 0.007695f
C1156 B.n1116 VSUBS 0.007695f
C1157 B.n1117 VSUBS 0.007695f
C1158 B.n1118 VSUBS 0.007695f
C1159 B.n1119 VSUBS 0.010042f
C1160 B.n1120 VSUBS 0.010697f
C1161 B.n1121 VSUBS 0.021272f
C1162 VDD1.t7 VSUBS 4.46593f
C1163 VDD1.t2 VSUBS 0.410179f
C1164 VDD1.t1 VSUBS 0.410179f
C1165 VDD1.n0 VSUBS 3.40883f
C1166 VDD1.n1 VSUBS 1.89675f
C1167 VDD1.t8 VSUBS 4.46592f
C1168 VDD1.t5 VSUBS 0.410179f
C1169 VDD1.t9 VSUBS 0.410179f
C1170 VDD1.n2 VSUBS 3.40883f
C1171 VDD1.n3 VSUBS 1.88705f
C1172 VDD1.t6 VSUBS 0.410179f
C1173 VDD1.t4 VSUBS 0.410179f
C1174 VDD1.n4 VSUBS 3.4454f
C1175 VDD1.n5 VSUBS 4.802f
C1176 VDD1.t0 VSUBS 0.410179f
C1177 VDD1.t3 VSUBS 0.410179f
C1178 VDD1.n6 VSUBS 3.40882f
C1179 VDD1.n7 VSUBS 4.92569f
C1180 VP.t5 VSUBS 3.91168f
C1181 VP.n0 VSUBS 1.44412f
C1182 VP.n1 VSUBS 0.023072f
C1183 VP.n2 VSUBS 0.021513f
C1184 VP.n3 VSUBS 0.023072f
C1185 VP.t3 VSUBS 3.91168f
C1186 VP.n4 VSUBS 1.34995f
C1187 VP.n5 VSUBS 0.023072f
C1188 VP.n6 VSUBS 0.040888f
C1189 VP.n7 VSUBS 0.023072f
C1190 VP.n8 VSUBS 0.032547f
C1191 VP.n9 VSUBS 0.023072f
C1192 VP.n10 VSUBS 0.024755f
C1193 VP.n11 VSUBS 0.023072f
C1194 VP.n12 VSUBS 0.022732f
C1195 VP.n13 VSUBS 0.023072f
C1196 VP.n14 VSUBS 0.021513f
C1197 VP.n15 VSUBS 0.023072f
C1198 VP.t1 VSUBS 3.91168f
C1199 VP.n16 VSUBS 1.44412f
C1200 VP.t6 VSUBS 3.91168f
C1201 VP.n17 VSUBS 1.44412f
C1202 VP.n18 VSUBS 0.023072f
C1203 VP.n19 VSUBS 0.021513f
C1204 VP.n20 VSUBS 0.023072f
C1205 VP.t9 VSUBS 3.91168f
C1206 VP.n21 VSUBS 1.34995f
C1207 VP.n22 VSUBS 0.023072f
C1208 VP.n23 VSUBS 0.040888f
C1209 VP.n24 VSUBS 0.023072f
C1210 VP.n25 VSUBS 0.032547f
C1211 VP.n26 VSUBS 0.023072f
C1212 VP.n27 VSUBS 0.024755f
C1213 VP.n28 VSUBS 0.023072f
C1214 VP.n29 VSUBS 0.022732f
C1215 VP.t2 VSUBS 4.22528f
C1216 VP.t7 VSUBS 3.91168f
C1217 VP.n30 VSUBS 1.42079f
C1218 VP.n31 VSUBS 1.36445f
C1219 VP.n32 VSUBS 0.27561f
C1220 VP.n33 VSUBS 0.023072f
C1221 VP.n34 VSUBS 0.043215f
C1222 VP.n35 VSUBS 0.043215f
C1223 VP.n36 VSUBS 0.040888f
C1224 VP.n37 VSUBS 0.023072f
C1225 VP.n38 VSUBS 0.023072f
C1226 VP.n39 VSUBS 0.023072f
C1227 VP.n40 VSUBS 0.045227f
C1228 VP.n41 VSUBS 0.043215f
C1229 VP.t8 VSUBS 3.91168f
C1230 VP.n42 VSUBS 1.34995f
C1231 VP.n43 VSUBS 0.032547f
C1232 VP.n44 VSUBS 0.023072f
C1233 VP.n45 VSUBS 0.023072f
C1234 VP.n46 VSUBS 0.023072f
C1235 VP.n47 VSUBS 0.043215f
C1236 VP.n48 VSUBS 0.045227f
C1237 VP.n49 VSUBS 0.024755f
C1238 VP.n50 VSUBS 0.023072f
C1239 VP.n51 VSUBS 0.023072f
C1240 VP.n52 VSUBS 0.023072f
C1241 VP.n53 VSUBS 0.043215f
C1242 VP.n54 VSUBS 0.043215f
C1243 VP.n55 VSUBS 0.022732f
C1244 VP.n56 VSUBS 0.023072f
C1245 VP.n57 VSUBS 0.023072f
C1246 VP.n58 VSUBS 0.042362f
C1247 VP.n59 VSUBS 0.043215f
C1248 VP.n60 VSUBS 0.04278f
C1249 VP.n61 VSUBS 0.023072f
C1250 VP.n62 VSUBS 0.023072f
C1251 VP.n63 VSUBS 0.023072f
C1252 VP.n64 VSUBS 0.046576f
C1253 VP.n65 VSUBS 0.043215f
C1254 VP.n66 VSUBS 0.034254f
C1255 VP.n67 VSUBS 0.037243f
C1256 VP.n68 VSUBS 1.77922f
C1257 VP.n69 VSUBS 1.79249f
C1258 VP.n70 VSUBS 0.037243f
C1259 VP.n71 VSUBS 0.034254f
C1260 VP.n72 VSUBS 0.043215f
C1261 VP.n73 VSUBS 0.046576f
C1262 VP.n74 VSUBS 0.023072f
C1263 VP.n75 VSUBS 0.023072f
C1264 VP.n76 VSUBS 0.023072f
C1265 VP.n77 VSUBS 0.04278f
C1266 VP.n78 VSUBS 0.043215f
C1267 VP.t4 VSUBS 3.91168f
C1268 VP.n79 VSUBS 1.34995f
C1269 VP.n80 VSUBS 0.042362f
C1270 VP.n81 VSUBS 0.023072f
C1271 VP.n82 VSUBS 0.023072f
C1272 VP.n83 VSUBS 0.023072f
C1273 VP.n84 VSUBS 0.043215f
C1274 VP.n85 VSUBS 0.043215f
C1275 VP.n86 VSUBS 0.040888f
C1276 VP.n87 VSUBS 0.023072f
C1277 VP.n88 VSUBS 0.023072f
C1278 VP.n89 VSUBS 0.023072f
C1279 VP.n90 VSUBS 0.045227f
C1280 VP.n91 VSUBS 0.043215f
C1281 VP.t0 VSUBS 3.91168f
C1282 VP.n92 VSUBS 1.34995f
C1283 VP.n93 VSUBS 0.032547f
C1284 VP.n94 VSUBS 0.023072f
C1285 VP.n95 VSUBS 0.023072f
C1286 VP.n96 VSUBS 0.023072f
C1287 VP.n97 VSUBS 0.043215f
C1288 VP.n98 VSUBS 0.045227f
C1289 VP.n99 VSUBS 0.024755f
C1290 VP.n100 VSUBS 0.023072f
C1291 VP.n101 VSUBS 0.023072f
C1292 VP.n102 VSUBS 0.023072f
C1293 VP.n103 VSUBS 0.043215f
C1294 VP.n104 VSUBS 0.043215f
C1295 VP.n105 VSUBS 0.022732f
C1296 VP.n106 VSUBS 0.023072f
C1297 VP.n107 VSUBS 0.023072f
C1298 VP.n108 VSUBS 0.042362f
C1299 VP.n109 VSUBS 0.043215f
C1300 VP.n110 VSUBS 0.04278f
C1301 VP.n111 VSUBS 0.023072f
C1302 VP.n112 VSUBS 0.023072f
C1303 VP.n113 VSUBS 0.023072f
C1304 VP.n114 VSUBS 0.046576f
C1305 VP.n115 VSUBS 0.043215f
C1306 VP.n116 VSUBS 0.034254f
C1307 VP.n117 VSUBS 0.037243f
C1308 VP.n118 VSUBS 0.057687f
C1309 VDD2.t9 VSUBS 4.45543f
C1310 VDD2.t5 VSUBS 0.409216f
C1311 VDD2.t0 VSUBS 0.409216f
C1312 VDD2.n0 VSUBS 3.40082f
C1313 VDD2.n1 VSUBS 1.88262f
C1314 VDD2.t6 VSUBS 0.409216f
C1315 VDD2.t2 VSUBS 0.409216f
C1316 VDD2.n2 VSUBS 3.4373f
C1317 VDD2.n3 VSUBS 4.61489f
C1318 VDD2.t1 VSUBS 4.41257f
C1319 VDD2.n4 VSUBS 4.86596f
C1320 VDD2.t3 VSUBS 0.409216f
C1321 VDD2.t7 VSUBS 0.409216f
C1322 VDD2.n5 VSUBS 3.40083f
C1323 VDD2.n6 VSUBS 0.950148f
C1324 VDD2.t4 VSUBS 0.409216f
C1325 VDD2.t8 VSUBS 0.409216f
C1326 VDD2.n7 VSUBS 3.43723f
C1327 VTAIL.t14 VSUBS 0.394569f
C1328 VTAIL.t16 VSUBS 0.394569f
C1329 VTAIL.n0 VSUBS 3.10872f
C1330 VTAIL.n1 VSUBS 1.09084f
C1331 VTAIL.t1 VSUBS 4.05927f
C1332 VTAIL.n2 VSUBS 1.28411f
C1333 VTAIL.t7 VSUBS 0.394569f
C1334 VTAIL.t6 VSUBS 0.394569f
C1335 VTAIL.n3 VSUBS 3.10872f
C1336 VTAIL.n4 VSUBS 1.26227f
C1337 VTAIL.t4 VSUBS 0.394569f
C1338 VTAIL.t3 VSUBS 0.394569f
C1339 VTAIL.n5 VSUBS 3.10872f
C1340 VTAIL.n6 VSUBS 3.31952f
C1341 VTAIL.t15 VSUBS 0.394569f
C1342 VTAIL.t18 VSUBS 0.394569f
C1343 VTAIL.n7 VSUBS 3.10873f
C1344 VTAIL.n8 VSUBS 3.31952f
C1345 VTAIL.t11 VSUBS 0.394569f
C1346 VTAIL.t19 VSUBS 0.394569f
C1347 VTAIL.n9 VSUBS 3.10873f
C1348 VTAIL.n10 VSUBS 1.26227f
C1349 VTAIL.t12 VSUBS 4.05928f
C1350 VTAIL.n11 VSUBS 1.2841f
C1351 VTAIL.t9 VSUBS 0.394569f
C1352 VTAIL.t5 VSUBS 0.394569f
C1353 VTAIL.n12 VSUBS 3.10873f
C1354 VTAIL.n13 VSUBS 1.15855f
C1355 VTAIL.t0 VSUBS 0.394569f
C1356 VTAIL.t8 VSUBS 0.394569f
C1357 VTAIL.n14 VSUBS 3.10873f
C1358 VTAIL.n15 VSUBS 1.26227f
C1359 VTAIL.t2 VSUBS 4.05927f
C1360 VTAIL.n16 VSUBS 3.15328f
C1361 VTAIL.t10 VSUBS 4.05927f
C1362 VTAIL.n17 VSUBS 3.15328f
C1363 VTAIL.t13 VSUBS 0.394569f
C1364 VTAIL.t17 VSUBS 0.394569f
C1365 VTAIL.n18 VSUBS 3.10872f
C1366 VTAIL.n19 VSUBS 1.03821f
C1367 VN.t7 VSUBS 3.6511f
C1368 VN.n0 VSUBS 1.34792f
C1369 VN.n1 VSUBS 0.021535f
C1370 VN.n2 VSUBS 0.02008f
C1371 VN.n3 VSUBS 0.021535f
C1372 VN.t3 VSUBS 3.6511f
C1373 VN.n4 VSUBS 1.26002f
C1374 VN.n5 VSUBS 0.021535f
C1375 VN.n6 VSUBS 0.038164f
C1376 VN.n7 VSUBS 0.021535f
C1377 VN.n8 VSUBS 0.030379f
C1378 VN.n9 VSUBS 0.021535f
C1379 VN.n10 VSUBS 0.023106f
C1380 VN.n11 VSUBS 0.021535f
C1381 VN.n12 VSUBS 0.021218f
C1382 VN.t4 VSUBS 3.6511f
C1383 VN.n13 VSUBS 1.32615f
C1384 VN.t0 VSUBS 3.94381f
C1385 VN.n14 VSUBS 1.27356f
C1386 VN.n15 VSUBS 0.25725f
C1387 VN.n16 VSUBS 0.021535f
C1388 VN.n17 VSUBS 0.040337f
C1389 VN.n18 VSUBS 0.040337f
C1390 VN.n19 VSUBS 0.038164f
C1391 VN.n20 VSUBS 0.021535f
C1392 VN.n21 VSUBS 0.021535f
C1393 VN.n22 VSUBS 0.021535f
C1394 VN.n23 VSUBS 0.042214f
C1395 VN.n24 VSUBS 0.040337f
C1396 VN.t9 VSUBS 3.6511f
C1397 VN.n25 VSUBS 1.26002f
C1398 VN.n26 VSUBS 0.030379f
C1399 VN.n27 VSUBS 0.021535f
C1400 VN.n28 VSUBS 0.021535f
C1401 VN.n29 VSUBS 0.021535f
C1402 VN.n30 VSUBS 0.040337f
C1403 VN.n31 VSUBS 0.042214f
C1404 VN.n32 VSUBS 0.023106f
C1405 VN.n33 VSUBS 0.021535f
C1406 VN.n34 VSUBS 0.021535f
C1407 VN.n35 VSUBS 0.021535f
C1408 VN.n36 VSUBS 0.040337f
C1409 VN.n37 VSUBS 0.040337f
C1410 VN.n38 VSUBS 0.021218f
C1411 VN.n39 VSUBS 0.021535f
C1412 VN.n40 VSUBS 0.021535f
C1413 VN.n41 VSUBS 0.03954f
C1414 VN.n42 VSUBS 0.040337f
C1415 VN.n43 VSUBS 0.039931f
C1416 VN.n44 VSUBS 0.021535f
C1417 VN.n45 VSUBS 0.021535f
C1418 VN.n46 VSUBS 0.021535f
C1419 VN.n47 VSUBS 0.043473f
C1420 VN.n48 VSUBS 0.040337f
C1421 VN.n49 VSUBS 0.031972f
C1422 VN.n50 VSUBS 0.034762f
C1423 VN.n51 VSUBS 0.053844f
C1424 VN.t8 VSUBS 3.6511f
C1425 VN.n52 VSUBS 1.34792f
C1426 VN.n53 VSUBS 0.021535f
C1427 VN.n54 VSUBS 0.02008f
C1428 VN.n55 VSUBS 0.021535f
C1429 VN.t6 VSUBS 3.6511f
C1430 VN.n56 VSUBS 1.26002f
C1431 VN.n57 VSUBS 0.021535f
C1432 VN.n58 VSUBS 0.038164f
C1433 VN.n59 VSUBS 0.021535f
C1434 VN.n60 VSUBS 0.030379f
C1435 VN.n61 VSUBS 0.021535f
C1436 VN.t2 VSUBS 3.6511f
C1437 VN.n62 VSUBS 1.26002f
C1438 VN.n63 VSUBS 0.023106f
C1439 VN.n64 VSUBS 0.021535f
C1440 VN.n65 VSUBS 0.021218f
C1441 VN.t1 VSUBS 3.94381f
C1442 VN.t5 VSUBS 3.6511f
C1443 VN.n66 VSUBS 1.32615f
C1444 VN.n67 VSUBS 1.27356f
C1445 VN.n68 VSUBS 0.25725f
C1446 VN.n69 VSUBS 0.021535f
C1447 VN.n70 VSUBS 0.040337f
C1448 VN.n71 VSUBS 0.040337f
C1449 VN.n72 VSUBS 0.038164f
C1450 VN.n73 VSUBS 0.021535f
C1451 VN.n74 VSUBS 0.021535f
C1452 VN.n75 VSUBS 0.021535f
C1453 VN.n76 VSUBS 0.042214f
C1454 VN.n77 VSUBS 0.040337f
C1455 VN.n78 VSUBS 0.030379f
C1456 VN.n79 VSUBS 0.021535f
C1457 VN.n80 VSUBS 0.021535f
C1458 VN.n81 VSUBS 0.021535f
C1459 VN.n82 VSUBS 0.040337f
C1460 VN.n83 VSUBS 0.042214f
C1461 VN.n84 VSUBS 0.023106f
C1462 VN.n85 VSUBS 0.021535f
C1463 VN.n86 VSUBS 0.021535f
C1464 VN.n87 VSUBS 0.021535f
C1465 VN.n88 VSUBS 0.040337f
C1466 VN.n89 VSUBS 0.040337f
C1467 VN.n90 VSUBS 0.021218f
C1468 VN.n91 VSUBS 0.021535f
C1469 VN.n92 VSUBS 0.021535f
C1470 VN.n93 VSUBS 0.03954f
C1471 VN.n94 VSUBS 0.040337f
C1472 VN.n95 VSUBS 0.039931f
C1473 VN.n96 VSUBS 0.021535f
C1474 VN.n97 VSUBS 0.021535f
C1475 VN.n98 VSUBS 0.021535f
C1476 VN.n99 VSUBS 0.043473f
C1477 VN.n100 VSUBS 0.040337f
C1478 VN.n101 VSUBS 0.031972f
C1479 VN.n102 VSUBS 0.034762f
C1480 VN.n103 VSUBS 1.6689f
.ends

