* NGSPICE file created from diff_pair_sample_1043.ext - technology: sky130A

.subckt diff_pair_sample_1043 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=2.92
X1 B.t8 B.t6 B.t7 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=2.92
X2 VDD2.t1 VN.t0 VTAIL.t2 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=2.92
X3 B.t5 B.t3 B.t4 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=2.92
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=2.92
X5 B.t2 B.t0 B.t1 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=2.92
X6 VDD1.t1 VP.t0 VTAIL.t0 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=2.92
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n2270_n1410# sky130_fd_pr__pfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=2.92
R0 B.n276 B.n37 585
R1 B.n278 B.n277 585
R2 B.n279 B.n36 585
R3 B.n281 B.n280 585
R4 B.n282 B.n35 585
R5 B.n284 B.n283 585
R6 B.n285 B.n34 585
R7 B.n287 B.n286 585
R8 B.n288 B.n33 585
R9 B.n290 B.n289 585
R10 B.n291 B.n32 585
R11 B.n293 B.n292 585
R12 B.n294 B.n29 585
R13 B.n297 B.n296 585
R14 B.n298 B.n28 585
R15 B.n300 B.n299 585
R16 B.n301 B.n27 585
R17 B.n303 B.n302 585
R18 B.n304 B.n26 585
R19 B.n306 B.n305 585
R20 B.n307 B.n25 585
R21 B.n309 B.n308 585
R22 B.n311 B.n310 585
R23 B.n312 B.n21 585
R24 B.n314 B.n313 585
R25 B.n315 B.n20 585
R26 B.n317 B.n316 585
R27 B.n318 B.n19 585
R28 B.n320 B.n319 585
R29 B.n321 B.n18 585
R30 B.n323 B.n322 585
R31 B.n324 B.n17 585
R32 B.n326 B.n325 585
R33 B.n327 B.n16 585
R34 B.n329 B.n328 585
R35 B.n275 B.n274 585
R36 B.n273 B.n38 585
R37 B.n272 B.n271 585
R38 B.n270 B.n39 585
R39 B.n269 B.n268 585
R40 B.n267 B.n40 585
R41 B.n266 B.n265 585
R42 B.n264 B.n41 585
R43 B.n263 B.n262 585
R44 B.n261 B.n42 585
R45 B.n260 B.n259 585
R46 B.n258 B.n43 585
R47 B.n257 B.n256 585
R48 B.n255 B.n44 585
R49 B.n254 B.n253 585
R50 B.n252 B.n45 585
R51 B.n251 B.n250 585
R52 B.n249 B.n46 585
R53 B.n248 B.n247 585
R54 B.n246 B.n47 585
R55 B.n245 B.n244 585
R56 B.n243 B.n48 585
R57 B.n242 B.n241 585
R58 B.n240 B.n49 585
R59 B.n239 B.n238 585
R60 B.n237 B.n50 585
R61 B.n236 B.n235 585
R62 B.n234 B.n51 585
R63 B.n233 B.n232 585
R64 B.n231 B.n52 585
R65 B.n230 B.n229 585
R66 B.n228 B.n53 585
R67 B.n227 B.n226 585
R68 B.n225 B.n54 585
R69 B.n224 B.n223 585
R70 B.n222 B.n55 585
R71 B.n221 B.n220 585
R72 B.n219 B.n56 585
R73 B.n218 B.n217 585
R74 B.n216 B.n57 585
R75 B.n215 B.n214 585
R76 B.n213 B.n58 585
R77 B.n212 B.n211 585
R78 B.n210 B.n59 585
R79 B.n209 B.n208 585
R80 B.n207 B.n60 585
R81 B.n206 B.n205 585
R82 B.n204 B.n61 585
R83 B.n203 B.n202 585
R84 B.n201 B.n62 585
R85 B.n200 B.n199 585
R86 B.n198 B.n63 585
R87 B.n197 B.n196 585
R88 B.n195 B.n64 585
R89 B.n194 B.n193 585
R90 B.n140 B.n139 585
R91 B.n141 B.n86 585
R92 B.n143 B.n142 585
R93 B.n144 B.n85 585
R94 B.n146 B.n145 585
R95 B.n147 B.n84 585
R96 B.n149 B.n148 585
R97 B.n150 B.n83 585
R98 B.n152 B.n151 585
R99 B.n153 B.n82 585
R100 B.n155 B.n154 585
R101 B.n156 B.n81 585
R102 B.n158 B.n157 585
R103 B.n160 B.n159 585
R104 B.n161 B.n77 585
R105 B.n163 B.n162 585
R106 B.n164 B.n76 585
R107 B.n166 B.n165 585
R108 B.n167 B.n75 585
R109 B.n169 B.n168 585
R110 B.n170 B.n74 585
R111 B.n172 B.n171 585
R112 B.n174 B.n71 585
R113 B.n176 B.n175 585
R114 B.n177 B.n70 585
R115 B.n179 B.n178 585
R116 B.n180 B.n69 585
R117 B.n182 B.n181 585
R118 B.n183 B.n68 585
R119 B.n185 B.n184 585
R120 B.n186 B.n67 585
R121 B.n188 B.n187 585
R122 B.n189 B.n66 585
R123 B.n191 B.n190 585
R124 B.n192 B.n65 585
R125 B.n138 B.n87 585
R126 B.n137 B.n136 585
R127 B.n135 B.n88 585
R128 B.n134 B.n133 585
R129 B.n132 B.n89 585
R130 B.n131 B.n130 585
R131 B.n129 B.n90 585
R132 B.n128 B.n127 585
R133 B.n126 B.n91 585
R134 B.n125 B.n124 585
R135 B.n123 B.n92 585
R136 B.n122 B.n121 585
R137 B.n120 B.n93 585
R138 B.n119 B.n118 585
R139 B.n117 B.n94 585
R140 B.n116 B.n115 585
R141 B.n114 B.n95 585
R142 B.n113 B.n112 585
R143 B.n111 B.n96 585
R144 B.n110 B.n109 585
R145 B.n108 B.n97 585
R146 B.n107 B.n106 585
R147 B.n105 B.n98 585
R148 B.n104 B.n103 585
R149 B.n102 B.n99 585
R150 B.n101 B.n100 585
R151 B.n2 B.n0 585
R152 B.n369 B.n1 585
R153 B.n368 B.n367 585
R154 B.n366 B.n3 585
R155 B.n365 B.n364 585
R156 B.n363 B.n4 585
R157 B.n362 B.n361 585
R158 B.n360 B.n5 585
R159 B.n359 B.n358 585
R160 B.n357 B.n6 585
R161 B.n356 B.n355 585
R162 B.n354 B.n7 585
R163 B.n353 B.n352 585
R164 B.n351 B.n8 585
R165 B.n350 B.n349 585
R166 B.n348 B.n9 585
R167 B.n347 B.n346 585
R168 B.n345 B.n10 585
R169 B.n344 B.n343 585
R170 B.n342 B.n11 585
R171 B.n341 B.n340 585
R172 B.n339 B.n12 585
R173 B.n338 B.n337 585
R174 B.n336 B.n13 585
R175 B.n335 B.n334 585
R176 B.n333 B.n14 585
R177 B.n332 B.n331 585
R178 B.n330 B.n15 585
R179 B.n371 B.n370 585
R180 B.n140 B.n87 554.963
R181 B.n328 B.n15 554.963
R182 B.n194 B.n65 554.963
R183 B.n274 B.n37 554.963
R184 B.n72 B.t8 236.006
R185 B.n30 B.t1 236.006
R186 B.n78 B.t5 236.006
R187 B.n22 B.t10 236.006
R188 B.n72 B.t6 226.724
R189 B.n78 B.t3 226.724
R190 B.n22 B.t9 226.724
R191 B.n30 B.t0 226.724
R192 B.n73 B.t7 172.976
R193 B.n31 B.t2 172.976
R194 B.n79 B.t4 172.975
R195 B.n23 B.t11 172.975
R196 B.n136 B.n87 163.367
R197 B.n136 B.n135 163.367
R198 B.n135 B.n134 163.367
R199 B.n134 B.n89 163.367
R200 B.n130 B.n89 163.367
R201 B.n130 B.n129 163.367
R202 B.n129 B.n128 163.367
R203 B.n128 B.n91 163.367
R204 B.n124 B.n91 163.367
R205 B.n124 B.n123 163.367
R206 B.n123 B.n122 163.367
R207 B.n122 B.n93 163.367
R208 B.n118 B.n93 163.367
R209 B.n118 B.n117 163.367
R210 B.n117 B.n116 163.367
R211 B.n116 B.n95 163.367
R212 B.n112 B.n95 163.367
R213 B.n112 B.n111 163.367
R214 B.n111 B.n110 163.367
R215 B.n110 B.n97 163.367
R216 B.n106 B.n97 163.367
R217 B.n106 B.n105 163.367
R218 B.n105 B.n104 163.367
R219 B.n104 B.n99 163.367
R220 B.n100 B.n99 163.367
R221 B.n100 B.n2 163.367
R222 B.n370 B.n2 163.367
R223 B.n370 B.n369 163.367
R224 B.n369 B.n368 163.367
R225 B.n368 B.n3 163.367
R226 B.n364 B.n3 163.367
R227 B.n364 B.n363 163.367
R228 B.n363 B.n362 163.367
R229 B.n362 B.n5 163.367
R230 B.n358 B.n5 163.367
R231 B.n358 B.n357 163.367
R232 B.n357 B.n356 163.367
R233 B.n356 B.n7 163.367
R234 B.n352 B.n7 163.367
R235 B.n352 B.n351 163.367
R236 B.n351 B.n350 163.367
R237 B.n350 B.n9 163.367
R238 B.n346 B.n9 163.367
R239 B.n346 B.n345 163.367
R240 B.n345 B.n344 163.367
R241 B.n344 B.n11 163.367
R242 B.n340 B.n11 163.367
R243 B.n340 B.n339 163.367
R244 B.n339 B.n338 163.367
R245 B.n338 B.n13 163.367
R246 B.n334 B.n13 163.367
R247 B.n334 B.n333 163.367
R248 B.n333 B.n332 163.367
R249 B.n332 B.n15 163.367
R250 B.n141 B.n140 163.367
R251 B.n142 B.n141 163.367
R252 B.n142 B.n85 163.367
R253 B.n146 B.n85 163.367
R254 B.n147 B.n146 163.367
R255 B.n148 B.n147 163.367
R256 B.n148 B.n83 163.367
R257 B.n152 B.n83 163.367
R258 B.n153 B.n152 163.367
R259 B.n154 B.n153 163.367
R260 B.n154 B.n81 163.367
R261 B.n158 B.n81 163.367
R262 B.n159 B.n158 163.367
R263 B.n159 B.n77 163.367
R264 B.n163 B.n77 163.367
R265 B.n164 B.n163 163.367
R266 B.n165 B.n164 163.367
R267 B.n165 B.n75 163.367
R268 B.n169 B.n75 163.367
R269 B.n170 B.n169 163.367
R270 B.n171 B.n170 163.367
R271 B.n171 B.n71 163.367
R272 B.n176 B.n71 163.367
R273 B.n177 B.n176 163.367
R274 B.n178 B.n177 163.367
R275 B.n178 B.n69 163.367
R276 B.n182 B.n69 163.367
R277 B.n183 B.n182 163.367
R278 B.n184 B.n183 163.367
R279 B.n184 B.n67 163.367
R280 B.n188 B.n67 163.367
R281 B.n189 B.n188 163.367
R282 B.n190 B.n189 163.367
R283 B.n190 B.n65 163.367
R284 B.n195 B.n194 163.367
R285 B.n196 B.n195 163.367
R286 B.n196 B.n63 163.367
R287 B.n200 B.n63 163.367
R288 B.n201 B.n200 163.367
R289 B.n202 B.n201 163.367
R290 B.n202 B.n61 163.367
R291 B.n206 B.n61 163.367
R292 B.n207 B.n206 163.367
R293 B.n208 B.n207 163.367
R294 B.n208 B.n59 163.367
R295 B.n212 B.n59 163.367
R296 B.n213 B.n212 163.367
R297 B.n214 B.n213 163.367
R298 B.n214 B.n57 163.367
R299 B.n218 B.n57 163.367
R300 B.n219 B.n218 163.367
R301 B.n220 B.n219 163.367
R302 B.n220 B.n55 163.367
R303 B.n224 B.n55 163.367
R304 B.n225 B.n224 163.367
R305 B.n226 B.n225 163.367
R306 B.n226 B.n53 163.367
R307 B.n230 B.n53 163.367
R308 B.n231 B.n230 163.367
R309 B.n232 B.n231 163.367
R310 B.n232 B.n51 163.367
R311 B.n236 B.n51 163.367
R312 B.n237 B.n236 163.367
R313 B.n238 B.n237 163.367
R314 B.n238 B.n49 163.367
R315 B.n242 B.n49 163.367
R316 B.n243 B.n242 163.367
R317 B.n244 B.n243 163.367
R318 B.n244 B.n47 163.367
R319 B.n248 B.n47 163.367
R320 B.n249 B.n248 163.367
R321 B.n250 B.n249 163.367
R322 B.n250 B.n45 163.367
R323 B.n254 B.n45 163.367
R324 B.n255 B.n254 163.367
R325 B.n256 B.n255 163.367
R326 B.n256 B.n43 163.367
R327 B.n260 B.n43 163.367
R328 B.n261 B.n260 163.367
R329 B.n262 B.n261 163.367
R330 B.n262 B.n41 163.367
R331 B.n266 B.n41 163.367
R332 B.n267 B.n266 163.367
R333 B.n268 B.n267 163.367
R334 B.n268 B.n39 163.367
R335 B.n272 B.n39 163.367
R336 B.n273 B.n272 163.367
R337 B.n274 B.n273 163.367
R338 B.n328 B.n327 163.367
R339 B.n327 B.n326 163.367
R340 B.n326 B.n17 163.367
R341 B.n322 B.n17 163.367
R342 B.n322 B.n321 163.367
R343 B.n321 B.n320 163.367
R344 B.n320 B.n19 163.367
R345 B.n316 B.n19 163.367
R346 B.n316 B.n315 163.367
R347 B.n315 B.n314 163.367
R348 B.n314 B.n21 163.367
R349 B.n310 B.n21 163.367
R350 B.n310 B.n309 163.367
R351 B.n309 B.n25 163.367
R352 B.n305 B.n25 163.367
R353 B.n305 B.n304 163.367
R354 B.n304 B.n303 163.367
R355 B.n303 B.n27 163.367
R356 B.n299 B.n27 163.367
R357 B.n299 B.n298 163.367
R358 B.n298 B.n297 163.367
R359 B.n297 B.n29 163.367
R360 B.n292 B.n29 163.367
R361 B.n292 B.n291 163.367
R362 B.n291 B.n290 163.367
R363 B.n290 B.n33 163.367
R364 B.n286 B.n33 163.367
R365 B.n286 B.n285 163.367
R366 B.n285 B.n284 163.367
R367 B.n284 B.n35 163.367
R368 B.n280 B.n35 163.367
R369 B.n280 B.n279 163.367
R370 B.n279 B.n278 163.367
R371 B.n278 B.n37 163.367
R372 B.n73 B.n72 63.0308
R373 B.n79 B.n78 63.0308
R374 B.n23 B.n22 63.0308
R375 B.n31 B.n30 63.0308
R376 B.n173 B.n73 59.5399
R377 B.n80 B.n79 59.5399
R378 B.n24 B.n23 59.5399
R379 B.n295 B.n31 59.5399
R380 B.n276 B.n275 36.059
R381 B.n330 B.n329 36.059
R382 B.n193 B.n192 36.059
R383 B.n139 B.n138 36.059
R384 B B.n371 18.0485
R385 B.n329 B.n16 10.6151
R386 B.n325 B.n16 10.6151
R387 B.n325 B.n324 10.6151
R388 B.n324 B.n323 10.6151
R389 B.n323 B.n18 10.6151
R390 B.n319 B.n18 10.6151
R391 B.n319 B.n318 10.6151
R392 B.n318 B.n317 10.6151
R393 B.n317 B.n20 10.6151
R394 B.n313 B.n20 10.6151
R395 B.n313 B.n312 10.6151
R396 B.n312 B.n311 10.6151
R397 B.n308 B.n307 10.6151
R398 B.n307 B.n306 10.6151
R399 B.n306 B.n26 10.6151
R400 B.n302 B.n26 10.6151
R401 B.n302 B.n301 10.6151
R402 B.n301 B.n300 10.6151
R403 B.n300 B.n28 10.6151
R404 B.n296 B.n28 10.6151
R405 B.n294 B.n293 10.6151
R406 B.n293 B.n32 10.6151
R407 B.n289 B.n32 10.6151
R408 B.n289 B.n288 10.6151
R409 B.n288 B.n287 10.6151
R410 B.n287 B.n34 10.6151
R411 B.n283 B.n34 10.6151
R412 B.n283 B.n282 10.6151
R413 B.n282 B.n281 10.6151
R414 B.n281 B.n36 10.6151
R415 B.n277 B.n36 10.6151
R416 B.n277 B.n276 10.6151
R417 B.n193 B.n64 10.6151
R418 B.n197 B.n64 10.6151
R419 B.n198 B.n197 10.6151
R420 B.n199 B.n198 10.6151
R421 B.n199 B.n62 10.6151
R422 B.n203 B.n62 10.6151
R423 B.n204 B.n203 10.6151
R424 B.n205 B.n204 10.6151
R425 B.n205 B.n60 10.6151
R426 B.n209 B.n60 10.6151
R427 B.n210 B.n209 10.6151
R428 B.n211 B.n210 10.6151
R429 B.n211 B.n58 10.6151
R430 B.n215 B.n58 10.6151
R431 B.n216 B.n215 10.6151
R432 B.n217 B.n216 10.6151
R433 B.n217 B.n56 10.6151
R434 B.n221 B.n56 10.6151
R435 B.n222 B.n221 10.6151
R436 B.n223 B.n222 10.6151
R437 B.n223 B.n54 10.6151
R438 B.n227 B.n54 10.6151
R439 B.n228 B.n227 10.6151
R440 B.n229 B.n228 10.6151
R441 B.n229 B.n52 10.6151
R442 B.n233 B.n52 10.6151
R443 B.n234 B.n233 10.6151
R444 B.n235 B.n234 10.6151
R445 B.n235 B.n50 10.6151
R446 B.n239 B.n50 10.6151
R447 B.n240 B.n239 10.6151
R448 B.n241 B.n240 10.6151
R449 B.n241 B.n48 10.6151
R450 B.n245 B.n48 10.6151
R451 B.n246 B.n245 10.6151
R452 B.n247 B.n246 10.6151
R453 B.n247 B.n46 10.6151
R454 B.n251 B.n46 10.6151
R455 B.n252 B.n251 10.6151
R456 B.n253 B.n252 10.6151
R457 B.n253 B.n44 10.6151
R458 B.n257 B.n44 10.6151
R459 B.n258 B.n257 10.6151
R460 B.n259 B.n258 10.6151
R461 B.n259 B.n42 10.6151
R462 B.n263 B.n42 10.6151
R463 B.n264 B.n263 10.6151
R464 B.n265 B.n264 10.6151
R465 B.n265 B.n40 10.6151
R466 B.n269 B.n40 10.6151
R467 B.n270 B.n269 10.6151
R468 B.n271 B.n270 10.6151
R469 B.n271 B.n38 10.6151
R470 B.n275 B.n38 10.6151
R471 B.n139 B.n86 10.6151
R472 B.n143 B.n86 10.6151
R473 B.n144 B.n143 10.6151
R474 B.n145 B.n144 10.6151
R475 B.n145 B.n84 10.6151
R476 B.n149 B.n84 10.6151
R477 B.n150 B.n149 10.6151
R478 B.n151 B.n150 10.6151
R479 B.n151 B.n82 10.6151
R480 B.n155 B.n82 10.6151
R481 B.n156 B.n155 10.6151
R482 B.n157 B.n156 10.6151
R483 B.n161 B.n160 10.6151
R484 B.n162 B.n161 10.6151
R485 B.n162 B.n76 10.6151
R486 B.n166 B.n76 10.6151
R487 B.n167 B.n166 10.6151
R488 B.n168 B.n167 10.6151
R489 B.n168 B.n74 10.6151
R490 B.n172 B.n74 10.6151
R491 B.n175 B.n174 10.6151
R492 B.n175 B.n70 10.6151
R493 B.n179 B.n70 10.6151
R494 B.n180 B.n179 10.6151
R495 B.n181 B.n180 10.6151
R496 B.n181 B.n68 10.6151
R497 B.n185 B.n68 10.6151
R498 B.n186 B.n185 10.6151
R499 B.n187 B.n186 10.6151
R500 B.n187 B.n66 10.6151
R501 B.n191 B.n66 10.6151
R502 B.n192 B.n191 10.6151
R503 B.n138 B.n137 10.6151
R504 B.n137 B.n88 10.6151
R505 B.n133 B.n88 10.6151
R506 B.n133 B.n132 10.6151
R507 B.n132 B.n131 10.6151
R508 B.n131 B.n90 10.6151
R509 B.n127 B.n90 10.6151
R510 B.n127 B.n126 10.6151
R511 B.n126 B.n125 10.6151
R512 B.n125 B.n92 10.6151
R513 B.n121 B.n92 10.6151
R514 B.n121 B.n120 10.6151
R515 B.n120 B.n119 10.6151
R516 B.n119 B.n94 10.6151
R517 B.n115 B.n94 10.6151
R518 B.n115 B.n114 10.6151
R519 B.n114 B.n113 10.6151
R520 B.n113 B.n96 10.6151
R521 B.n109 B.n96 10.6151
R522 B.n109 B.n108 10.6151
R523 B.n108 B.n107 10.6151
R524 B.n107 B.n98 10.6151
R525 B.n103 B.n98 10.6151
R526 B.n103 B.n102 10.6151
R527 B.n102 B.n101 10.6151
R528 B.n101 B.n0 10.6151
R529 B.n367 B.n1 10.6151
R530 B.n367 B.n366 10.6151
R531 B.n366 B.n365 10.6151
R532 B.n365 B.n4 10.6151
R533 B.n361 B.n4 10.6151
R534 B.n361 B.n360 10.6151
R535 B.n360 B.n359 10.6151
R536 B.n359 B.n6 10.6151
R537 B.n355 B.n6 10.6151
R538 B.n355 B.n354 10.6151
R539 B.n354 B.n353 10.6151
R540 B.n353 B.n8 10.6151
R541 B.n349 B.n8 10.6151
R542 B.n349 B.n348 10.6151
R543 B.n348 B.n347 10.6151
R544 B.n347 B.n10 10.6151
R545 B.n343 B.n10 10.6151
R546 B.n343 B.n342 10.6151
R547 B.n342 B.n341 10.6151
R548 B.n341 B.n12 10.6151
R549 B.n337 B.n12 10.6151
R550 B.n337 B.n336 10.6151
R551 B.n336 B.n335 10.6151
R552 B.n335 B.n14 10.6151
R553 B.n331 B.n14 10.6151
R554 B.n331 B.n330 10.6151
R555 B.n308 B.n24 6.5566
R556 B.n296 B.n295 6.5566
R557 B.n160 B.n80 6.5566
R558 B.n173 B.n172 6.5566
R559 B.n311 B.n24 4.05904
R560 B.n295 B.n294 4.05904
R561 B.n157 B.n80 4.05904
R562 B.n174 B.n173 4.05904
R563 B.n371 B.n0 2.81026
R564 B.n371 B.n1 2.81026
R565 VN VN.t1 97.4267
R566 VN VN.t0 59.7676
R567 VTAIL.n3 VTAIL.t2 172.166
R568 VTAIL.n0 VTAIL.t1 172.166
R569 VTAIL.n2 VTAIL.t0 172.166
R570 VTAIL.n1 VTAIL.t3 172.166
R571 VTAIL.n1 VTAIL.n0 19.8755
R572 VTAIL.n3 VTAIL.n2 17.0738
R573 VTAIL.n2 VTAIL.n1 1.87119
R574 VTAIL VTAIL.n0 1.22895
R575 VTAIL VTAIL.n3 0.642741
R576 VDD2.n0 VDD2.t1 220.012
R577 VDD2.n0 VDD2.t0 188.845
R578 VDD2 VDD2.n0 0.759121
R579 VP.n0 VP.t0 97.425
R580 VP.n0 VP.t1 59.3363
R581 VP VP.n0 0.431811
R582 VDD1 VDD1.t0 221.238
R583 VDD1 VDD1.t1 189.603
C0 VN B 0.954017f
C1 VTAIL w_n2270_n1410# 1.35148f
C2 VDD2 VTAIL 2.63641f
C3 VN VP 3.79974f
C4 VDD1 w_n2270_n1410# 1.13536f
C5 VTAIL B 1.44566f
C6 VDD2 VDD1 0.712366f
C7 VTAIL VP 1.05603f
C8 VDD1 B 0.96848f
C9 VDD2 w_n2270_n1410# 1.1645f
C10 B w_n2270_n1410# 6.44075f
C11 VTAIL VN 1.04189f
C12 VDD1 VP 0.927568f
C13 VDD2 B 1.00177f
C14 VP w_n2270_n1410# 3.2471f
C15 VDD1 VN 0.15428f
C16 VDD2 VP 0.352508f
C17 VN w_n2270_n1410# 2.96114f
C18 VP B 1.43115f
C19 VDD2 VN 0.730923f
C20 VDD1 VTAIL 2.58131f
C21 VDD2 VSUBS 0.58115f
C22 VDD1 VSUBS 2.798261f
C23 VTAIL VSUBS 0.389643f
C24 VN VSUBS 5.61565f
C25 VP VSUBS 1.303614f
C26 B VSUBS 3.140985f
C27 w_n2270_n1410# VSUBS 40.7783f
C28 VDD1.t1 VSUBS 0.202923f
C29 VDD1.t0 VSUBS 0.333824f
C30 VP.t1 VSUBS 1.25428f
C31 VP.t0 VSUBS 2.12312f
C32 VP.n0 VSUBS 3.47897f
C33 VDD2.t1 VSUBS 0.329618f
C34 VDD2.t0 VSUBS 0.20689f
C35 VDD2.n0 VSUBS 1.94242f
C36 VTAIL.t1 VSUBS 0.226862f
C37 VTAIL.n0 VSUBS 1.12451f
C38 VTAIL.t3 VSUBS 0.226863f
C39 VTAIL.n1 VSUBS 1.168f
C40 VTAIL.t0 VSUBS 0.226862f
C41 VTAIL.n2 VSUBS 0.978274f
C42 VTAIL.t2 VSUBS 0.226862f
C43 VTAIL.n3 VSUBS 0.895086f
C44 VN.t0 VSUBS 1.20973f
C45 VN.t1 VSUBS 2.04756f
C46 B.n0 VSUBS 0.005644f
C47 B.n1 VSUBS 0.005644f
C48 B.n2 VSUBS 0.008926f
C49 B.n3 VSUBS 0.008926f
C50 B.n4 VSUBS 0.008926f
C51 B.n5 VSUBS 0.008926f
C52 B.n6 VSUBS 0.008926f
C53 B.n7 VSUBS 0.008926f
C54 B.n8 VSUBS 0.008926f
C55 B.n9 VSUBS 0.008926f
C56 B.n10 VSUBS 0.008926f
C57 B.n11 VSUBS 0.008926f
C58 B.n12 VSUBS 0.008926f
C59 B.n13 VSUBS 0.008926f
C60 B.n14 VSUBS 0.008926f
C61 B.n15 VSUBS 0.021767f
C62 B.n16 VSUBS 0.008926f
C63 B.n17 VSUBS 0.008926f
C64 B.n18 VSUBS 0.008926f
C65 B.n19 VSUBS 0.008926f
C66 B.n20 VSUBS 0.008926f
C67 B.n21 VSUBS 0.008926f
C68 B.t11 VSUBS 0.062187f
C69 B.t10 VSUBS 0.079717f
C70 B.t9 VSUBS 0.404995f
C71 B.n22 VSUBS 0.097626f
C72 B.n23 VSUBS 0.078367f
C73 B.n24 VSUBS 0.02068f
C74 B.n25 VSUBS 0.008926f
C75 B.n26 VSUBS 0.008926f
C76 B.n27 VSUBS 0.008926f
C77 B.n28 VSUBS 0.008926f
C78 B.n29 VSUBS 0.008926f
C79 B.t2 VSUBS 0.062187f
C80 B.t1 VSUBS 0.079717f
C81 B.t0 VSUBS 0.404995f
C82 B.n30 VSUBS 0.097626f
C83 B.n31 VSUBS 0.078367f
C84 B.n32 VSUBS 0.008926f
C85 B.n33 VSUBS 0.008926f
C86 B.n34 VSUBS 0.008926f
C87 B.n35 VSUBS 0.008926f
C88 B.n36 VSUBS 0.008926f
C89 B.n37 VSUBS 0.022862f
C90 B.n38 VSUBS 0.008926f
C91 B.n39 VSUBS 0.008926f
C92 B.n40 VSUBS 0.008926f
C93 B.n41 VSUBS 0.008926f
C94 B.n42 VSUBS 0.008926f
C95 B.n43 VSUBS 0.008926f
C96 B.n44 VSUBS 0.008926f
C97 B.n45 VSUBS 0.008926f
C98 B.n46 VSUBS 0.008926f
C99 B.n47 VSUBS 0.008926f
C100 B.n48 VSUBS 0.008926f
C101 B.n49 VSUBS 0.008926f
C102 B.n50 VSUBS 0.008926f
C103 B.n51 VSUBS 0.008926f
C104 B.n52 VSUBS 0.008926f
C105 B.n53 VSUBS 0.008926f
C106 B.n54 VSUBS 0.008926f
C107 B.n55 VSUBS 0.008926f
C108 B.n56 VSUBS 0.008926f
C109 B.n57 VSUBS 0.008926f
C110 B.n58 VSUBS 0.008926f
C111 B.n59 VSUBS 0.008926f
C112 B.n60 VSUBS 0.008926f
C113 B.n61 VSUBS 0.008926f
C114 B.n62 VSUBS 0.008926f
C115 B.n63 VSUBS 0.008926f
C116 B.n64 VSUBS 0.008926f
C117 B.n65 VSUBS 0.022862f
C118 B.n66 VSUBS 0.008926f
C119 B.n67 VSUBS 0.008926f
C120 B.n68 VSUBS 0.008926f
C121 B.n69 VSUBS 0.008926f
C122 B.n70 VSUBS 0.008926f
C123 B.n71 VSUBS 0.008926f
C124 B.t7 VSUBS 0.062187f
C125 B.t8 VSUBS 0.079717f
C126 B.t6 VSUBS 0.404995f
C127 B.n72 VSUBS 0.097626f
C128 B.n73 VSUBS 0.078367f
C129 B.n74 VSUBS 0.008926f
C130 B.n75 VSUBS 0.008926f
C131 B.n76 VSUBS 0.008926f
C132 B.n77 VSUBS 0.008926f
C133 B.t4 VSUBS 0.062187f
C134 B.t5 VSUBS 0.079717f
C135 B.t3 VSUBS 0.404995f
C136 B.n78 VSUBS 0.097626f
C137 B.n79 VSUBS 0.078367f
C138 B.n80 VSUBS 0.02068f
C139 B.n81 VSUBS 0.008926f
C140 B.n82 VSUBS 0.008926f
C141 B.n83 VSUBS 0.008926f
C142 B.n84 VSUBS 0.008926f
C143 B.n85 VSUBS 0.008926f
C144 B.n86 VSUBS 0.008926f
C145 B.n87 VSUBS 0.021767f
C146 B.n88 VSUBS 0.008926f
C147 B.n89 VSUBS 0.008926f
C148 B.n90 VSUBS 0.008926f
C149 B.n91 VSUBS 0.008926f
C150 B.n92 VSUBS 0.008926f
C151 B.n93 VSUBS 0.008926f
C152 B.n94 VSUBS 0.008926f
C153 B.n95 VSUBS 0.008926f
C154 B.n96 VSUBS 0.008926f
C155 B.n97 VSUBS 0.008926f
C156 B.n98 VSUBS 0.008926f
C157 B.n99 VSUBS 0.008926f
C158 B.n100 VSUBS 0.008926f
C159 B.n101 VSUBS 0.008926f
C160 B.n102 VSUBS 0.008926f
C161 B.n103 VSUBS 0.008926f
C162 B.n104 VSUBS 0.008926f
C163 B.n105 VSUBS 0.008926f
C164 B.n106 VSUBS 0.008926f
C165 B.n107 VSUBS 0.008926f
C166 B.n108 VSUBS 0.008926f
C167 B.n109 VSUBS 0.008926f
C168 B.n110 VSUBS 0.008926f
C169 B.n111 VSUBS 0.008926f
C170 B.n112 VSUBS 0.008926f
C171 B.n113 VSUBS 0.008926f
C172 B.n114 VSUBS 0.008926f
C173 B.n115 VSUBS 0.008926f
C174 B.n116 VSUBS 0.008926f
C175 B.n117 VSUBS 0.008926f
C176 B.n118 VSUBS 0.008926f
C177 B.n119 VSUBS 0.008926f
C178 B.n120 VSUBS 0.008926f
C179 B.n121 VSUBS 0.008926f
C180 B.n122 VSUBS 0.008926f
C181 B.n123 VSUBS 0.008926f
C182 B.n124 VSUBS 0.008926f
C183 B.n125 VSUBS 0.008926f
C184 B.n126 VSUBS 0.008926f
C185 B.n127 VSUBS 0.008926f
C186 B.n128 VSUBS 0.008926f
C187 B.n129 VSUBS 0.008926f
C188 B.n130 VSUBS 0.008926f
C189 B.n131 VSUBS 0.008926f
C190 B.n132 VSUBS 0.008926f
C191 B.n133 VSUBS 0.008926f
C192 B.n134 VSUBS 0.008926f
C193 B.n135 VSUBS 0.008926f
C194 B.n136 VSUBS 0.008926f
C195 B.n137 VSUBS 0.008926f
C196 B.n138 VSUBS 0.021767f
C197 B.n139 VSUBS 0.022862f
C198 B.n140 VSUBS 0.022862f
C199 B.n141 VSUBS 0.008926f
C200 B.n142 VSUBS 0.008926f
C201 B.n143 VSUBS 0.008926f
C202 B.n144 VSUBS 0.008926f
C203 B.n145 VSUBS 0.008926f
C204 B.n146 VSUBS 0.008926f
C205 B.n147 VSUBS 0.008926f
C206 B.n148 VSUBS 0.008926f
C207 B.n149 VSUBS 0.008926f
C208 B.n150 VSUBS 0.008926f
C209 B.n151 VSUBS 0.008926f
C210 B.n152 VSUBS 0.008926f
C211 B.n153 VSUBS 0.008926f
C212 B.n154 VSUBS 0.008926f
C213 B.n155 VSUBS 0.008926f
C214 B.n156 VSUBS 0.008926f
C215 B.n157 VSUBS 0.006169f
C216 B.n158 VSUBS 0.008926f
C217 B.n159 VSUBS 0.008926f
C218 B.n160 VSUBS 0.007219f
C219 B.n161 VSUBS 0.008926f
C220 B.n162 VSUBS 0.008926f
C221 B.n163 VSUBS 0.008926f
C222 B.n164 VSUBS 0.008926f
C223 B.n165 VSUBS 0.008926f
C224 B.n166 VSUBS 0.008926f
C225 B.n167 VSUBS 0.008926f
C226 B.n168 VSUBS 0.008926f
C227 B.n169 VSUBS 0.008926f
C228 B.n170 VSUBS 0.008926f
C229 B.n171 VSUBS 0.008926f
C230 B.n172 VSUBS 0.007219f
C231 B.n173 VSUBS 0.02068f
C232 B.n174 VSUBS 0.006169f
C233 B.n175 VSUBS 0.008926f
C234 B.n176 VSUBS 0.008926f
C235 B.n177 VSUBS 0.008926f
C236 B.n178 VSUBS 0.008926f
C237 B.n179 VSUBS 0.008926f
C238 B.n180 VSUBS 0.008926f
C239 B.n181 VSUBS 0.008926f
C240 B.n182 VSUBS 0.008926f
C241 B.n183 VSUBS 0.008926f
C242 B.n184 VSUBS 0.008926f
C243 B.n185 VSUBS 0.008926f
C244 B.n186 VSUBS 0.008926f
C245 B.n187 VSUBS 0.008926f
C246 B.n188 VSUBS 0.008926f
C247 B.n189 VSUBS 0.008926f
C248 B.n190 VSUBS 0.008926f
C249 B.n191 VSUBS 0.008926f
C250 B.n192 VSUBS 0.022862f
C251 B.n193 VSUBS 0.021767f
C252 B.n194 VSUBS 0.021767f
C253 B.n195 VSUBS 0.008926f
C254 B.n196 VSUBS 0.008926f
C255 B.n197 VSUBS 0.008926f
C256 B.n198 VSUBS 0.008926f
C257 B.n199 VSUBS 0.008926f
C258 B.n200 VSUBS 0.008926f
C259 B.n201 VSUBS 0.008926f
C260 B.n202 VSUBS 0.008926f
C261 B.n203 VSUBS 0.008926f
C262 B.n204 VSUBS 0.008926f
C263 B.n205 VSUBS 0.008926f
C264 B.n206 VSUBS 0.008926f
C265 B.n207 VSUBS 0.008926f
C266 B.n208 VSUBS 0.008926f
C267 B.n209 VSUBS 0.008926f
C268 B.n210 VSUBS 0.008926f
C269 B.n211 VSUBS 0.008926f
C270 B.n212 VSUBS 0.008926f
C271 B.n213 VSUBS 0.008926f
C272 B.n214 VSUBS 0.008926f
C273 B.n215 VSUBS 0.008926f
C274 B.n216 VSUBS 0.008926f
C275 B.n217 VSUBS 0.008926f
C276 B.n218 VSUBS 0.008926f
C277 B.n219 VSUBS 0.008926f
C278 B.n220 VSUBS 0.008926f
C279 B.n221 VSUBS 0.008926f
C280 B.n222 VSUBS 0.008926f
C281 B.n223 VSUBS 0.008926f
C282 B.n224 VSUBS 0.008926f
C283 B.n225 VSUBS 0.008926f
C284 B.n226 VSUBS 0.008926f
C285 B.n227 VSUBS 0.008926f
C286 B.n228 VSUBS 0.008926f
C287 B.n229 VSUBS 0.008926f
C288 B.n230 VSUBS 0.008926f
C289 B.n231 VSUBS 0.008926f
C290 B.n232 VSUBS 0.008926f
C291 B.n233 VSUBS 0.008926f
C292 B.n234 VSUBS 0.008926f
C293 B.n235 VSUBS 0.008926f
C294 B.n236 VSUBS 0.008926f
C295 B.n237 VSUBS 0.008926f
C296 B.n238 VSUBS 0.008926f
C297 B.n239 VSUBS 0.008926f
C298 B.n240 VSUBS 0.008926f
C299 B.n241 VSUBS 0.008926f
C300 B.n242 VSUBS 0.008926f
C301 B.n243 VSUBS 0.008926f
C302 B.n244 VSUBS 0.008926f
C303 B.n245 VSUBS 0.008926f
C304 B.n246 VSUBS 0.008926f
C305 B.n247 VSUBS 0.008926f
C306 B.n248 VSUBS 0.008926f
C307 B.n249 VSUBS 0.008926f
C308 B.n250 VSUBS 0.008926f
C309 B.n251 VSUBS 0.008926f
C310 B.n252 VSUBS 0.008926f
C311 B.n253 VSUBS 0.008926f
C312 B.n254 VSUBS 0.008926f
C313 B.n255 VSUBS 0.008926f
C314 B.n256 VSUBS 0.008926f
C315 B.n257 VSUBS 0.008926f
C316 B.n258 VSUBS 0.008926f
C317 B.n259 VSUBS 0.008926f
C318 B.n260 VSUBS 0.008926f
C319 B.n261 VSUBS 0.008926f
C320 B.n262 VSUBS 0.008926f
C321 B.n263 VSUBS 0.008926f
C322 B.n264 VSUBS 0.008926f
C323 B.n265 VSUBS 0.008926f
C324 B.n266 VSUBS 0.008926f
C325 B.n267 VSUBS 0.008926f
C326 B.n268 VSUBS 0.008926f
C327 B.n269 VSUBS 0.008926f
C328 B.n270 VSUBS 0.008926f
C329 B.n271 VSUBS 0.008926f
C330 B.n272 VSUBS 0.008926f
C331 B.n273 VSUBS 0.008926f
C332 B.n274 VSUBS 0.021767f
C333 B.n275 VSUBS 0.022722f
C334 B.n276 VSUBS 0.021907f
C335 B.n277 VSUBS 0.008926f
C336 B.n278 VSUBS 0.008926f
C337 B.n279 VSUBS 0.008926f
C338 B.n280 VSUBS 0.008926f
C339 B.n281 VSUBS 0.008926f
C340 B.n282 VSUBS 0.008926f
C341 B.n283 VSUBS 0.008926f
C342 B.n284 VSUBS 0.008926f
C343 B.n285 VSUBS 0.008926f
C344 B.n286 VSUBS 0.008926f
C345 B.n287 VSUBS 0.008926f
C346 B.n288 VSUBS 0.008926f
C347 B.n289 VSUBS 0.008926f
C348 B.n290 VSUBS 0.008926f
C349 B.n291 VSUBS 0.008926f
C350 B.n292 VSUBS 0.008926f
C351 B.n293 VSUBS 0.008926f
C352 B.n294 VSUBS 0.006169f
C353 B.n295 VSUBS 0.02068f
C354 B.n296 VSUBS 0.007219f
C355 B.n297 VSUBS 0.008926f
C356 B.n298 VSUBS 0.008926f
C357 B.n299 VSUBS 0.008926f
C358 B.n300 VSUBS 0.008926f
C359 B.n301 VSUBS 0.008926f
C360 B.n302 VSUBS 0.008926f
C361 B.n303 VSUBS 0.008926f
C362 B.n304 VSUBS 0.008926f
C363 B.n305 VSUBS 0.008926f
C364 B.n306 VSUBS 0.008926f
C365 B.n307 VSUBS 0.008926f
C366 B.n308 VSUBS 0.007219f
C367 B.n309 VSUBS 0.008926f
C368 B.n310 VSUBS 0.008926f
C369 B.n311 VSUBS 0.006169f
C370 B.n312 VSUBS 0.008926f
C371 B.n313 VSUBS 0.008926f
C372 B.n314 VSUBS 0.008926f
C373 B.n315 VSUBS 0.008926f
C374 B.n316 VSUBS 0.008926f
C375 B.n317 VSUBS 0.008926f
C376 B.n318 VSUBS 0.008926f
C377 B.n319 VSUBS 0.008926f
C378 B.n320 VSUBS 0.008926f
C379 B.n321 VSUBS 0.008926f
C380 B.n322 VSUBS 0.008926f
C381 B.n323 VSUBS 0.008926f
C382 B.n324 VSUBS 0.008926f
C383 B.n325 VSUBS 0.008926f
C384 B.n326 VSUBS 0.008926f
C385 B.n327 VSUBS 0.008926f
C386 B.n328 VSUBS 0.022862f
C387 B.n329 VSUBS 0.022862f
C388 B.n330 VSUBS 0.021767f
C389 B.n331 VSUBS 0.008926f
C390 B.n332 VSUBS 0.008926f
C391 B.n333 VSUBS 0.008926f
C392 B.n334 VSUBS 0.008926f
C393 B.n335 VSUBS 0.008926f
C394 B.n336 VSUBS 0.008926f
C395 B.n337 VSUBS 0.008926f
C396 B.n338 VSUBS 0.008926f
C397 B.n339 VSUBS 0.008926f
C398 B.n340 VSUBS 0.008926f
C399 B.n341 VSUBS 0.008926f
C400 B.n342 VSUBS 0.008926f
C401 B.n343 VSUBS 0.008926f
C402 B.n344 VSUBS 0.008926f
C403 B.n345 VSUBS 0.008926f
C404 B.n346 VSUBS 0.008926f
C405 B.n347 VSUBS 0.008926f
C406 B.n348 VSUBS 0.008926f
C407 B.n349 VSUBS 0.008926f
C408 B.n350 VSUBS 0.008926f
C409 B.n351 VSUBS 0.008926f
C410 B.n352 VSUBS 0.008926f
C411 B.n353 VSUBS 0.008926f
C412 B.n354 VSUBS 0.008926f
C413 B.n355 VSUBS 0.008926f
C414 B.n356 VSUBS 0.008926f
C415 B.n357 VSUBS 0.008926f
C416 B.n358 VSUBS 0.008926f
C417 B.n359 VSUBS 0.008926f
C418 B.n360 VSUBS 0.008926f
C419 B.n361 VSUBS 0.008926f
C420 B.n362 VSUBS 0.008926f
C421 B.n363 VSUBS 0.008926f
C422 B.n364 VSUBS 0.008926f
C423 B.n365 VSUBS 0.008926f
C424 B.n366 VSUBS 0.008926f
C425 B.n367 VSUBS 0.008926f
C426 B.n368 VSUBS 0.008926f
C427 B.n369 VSUBS 0.008926f
C428 B.n370 VSUBS 0.008926f
C429 B.n371 VSUBS 0.020211f
.ends

