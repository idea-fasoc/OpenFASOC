* NGSPICE file created from diff_pair_sample_0389.ext - technology: sky130A

.subckt diff_pair_sample_0389 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.92
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.92
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.92
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.92
X4 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.92
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.92
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.92
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.92
R0 B.n723 B.n722 585
R1 B.n724 B.n723 585
R2 B.n288 B.n107 585
R3 B.n287 B.n286 585
R4 B.n285 B.n284 585
R5 B.n283 B.n282 585
R6 B.n281 B.n280 585
R7 B.n279 B.n278 585
R8 B.n277 B.n276 585
R9 B.n275 B.n274 585
R10 B.n273 B.n272 585
R11 B.n271 B.n270 585
R12 B.n269 B.n268 585
R13 B.n267 B.n266 585
R14 B.n265 B.n264 585
R15 B.n263 B.n262 585
R16 B.n261 B.n260 585
R17 B.n259 B.n258 585
R18 B.n257 B.n256 585
R19 B.n255 B.n254 585
R20 B.n253 B.n252 585
R21 B.n251 B.n250 585
R22 B.n249 B.n248 585
R23 B.n247 B.n246 585
R24 B.n245 B.n244 585
R25 B.n243 B.n242 585
R26 B.n241 B.n240 585
R27 B.n239 B.n238 585
R28 B.n237 B.n236 585
R29 B.n235 B.n234 585
R30 B.n233 B.n232 585
R31 B.n231 B.n230 585
R32 B.n229 B.n228 585
R33 B.n227 B.n226 585
R34 B.n225 B.n224 585
R35 B.n223 B.n222 585
R36 B.n221 B.n220 585
R37 B.n219 B.n218 585
R38 B.n217 B.n216 585
R39 B.n215 B.n214 585
R40 B.n213 B.n212 585
R41 B.n210 B.n209 585
R42 B.n208 B.n207 585
R43 B.n206 B.n205 585
R44 B.n204 B.n203 585
R45 B.n202 B.n201 585
R46 B.n200 B.n199 585
R47 B.n198 B.n197 585
R48 B.n196 B.n195 585
R49 B.n194 B.n193 585
R50 B.n192 B.n191 585
R51 B.n190 B.n189 585
R52 B.n188 B.n187 585
R53 B.n186 B.n185 585
R54 B.n184 B.n183 585
R55 B.n182 B.n181 585
R56 B.n180 B.n179 585
R57 B.n178 B.n177 585
R58 B.n176 B.n175 585
R59 B.n174 B.n173 585
R60 B.n172 B.n171 585
R61 B.n170 B.n169 585
R62 B.n168 B.n167 585
R63 B.n166 B.n165 585
R64 B.n164 B.n163 585
R65 B.n162 B.n161 585
R66 B.n160 B.n159 585
R67 B.n158 B.n157 585
R68 B.n156 B.n155 585
R69 B.n154 B.n153 585
R70 B.n152 B.n151 585
R71 B.n150 B.n149 585
R72 B.n148 B.n147 585
R73 B.n146 B.n145 585
R74 B.n144 B.n143 585
R75 B.n142 B.n141 585
R76 B.n140 B.n139 585
R77 B.n138 B.n137 585
R78 B.n136 B.n135 585
R79 B.n134 B.n133 585
R80 B.n132 B.n131 585
R81 B.n130 B.n129 585
R82 B.n128 B.n127 585
R83 B.n126 B.n125 585
R84 B.n124 B.n123 585
R85 B.n122 B.n121 585
R86 B.n120 B.n119 585
R87 B.n118 B.n117 585
R88 B.n116 B.n115 585
R89 B.n114 B.n113 585
R90 B.n721 B.n62 585
R91 B.n725 B.n62 585
R92 B.n720 B.n61 585
R93 B.n726 B.n61 585
R94 B.n719 B.n718 585
R95 B.n718 B.n57 585
R96 B.n717 B.n56 585
R97 B.n732 B.n56 585
R98 B.n716 B.n55 585
R99 B.n733 B.n55 585
R100 B.n715 B.n54 585
R101 B.n734 B.n54 585
R102 B.n714 B.n713 585
R103 B.n713 B.n50 585
R104 B.n712 B.n49 585
R105 B.n740 B.n49 585
R106 B.n711 B.n48 585
R107 B.n741 B.n48 585
R108 B.n710 B.n47 585
R109 B.n742 B.n47 585
R110 B.n709 B.n708 585
R111 B.n708 B.n43 585
R112 B.n707 B.n42 585
R113 B.n748 B.n42 585
R114 B.n706 B.n41 585
R115 B.n749 B.n41 585
R116 B.n705 B.n40 585
R117 B.n750 B.n40 585
R118 B.n704 B.n703 585
R119 B.n703 B.n36 585
R120 B.n702 B.n35 585
R121 B.n756 B.n35 585
R122 B.n701 B.n34 585
R123 B.n757 B.n34 585
R124 B.n700 B.n33 585
R125 B.n758 B.n33 585
R126 B.n699 B.n698 585
R127 B.n698 B.n29 585
R128 B.n697 B.n28 585
R129 B.n764 B.n28 585
R130 B.n696 B.n27 585
R131 B.n765 B.n27 585
R132 B.n695 B.n26 585
R133 B.n766 B.n26 585
R134 B.n694 B.n693 585
R135 B.n693 B.n22 585
R136 B.n692 B.n21 585
R137 B.n772 B.n21 585
R138 B.n691 B.n20 585
R139 B.n773 B.n20 585
R140 B.n690 B.n19 585
R141 B.n774 B.n19 585
R142 B.n689 B.n688 585
R143 B.n688 B.n15 585
R144 B.n687 B.n14 585
R145 B.n780 B.n14 585
R146 B.n686 B.n13 585
R147 B.n781 B.n13 585
R148 B.n685 B.n12 585
R149 B.n782 B.n12 585
R150 B.n684 B.n683 585
R151 B.n683 B.n8 585
R152 B.n682 B.n7 585
R153 B.n788 B.n7 585
R154 B.n681 B.n6 585
R155 B.n789 B.n6 585
R156 B.n680 B.n5 585
R157 B.n790 B.n5 585
R158 B.n679 B.n678 585
R159 B.n678 B.n4 585
R160 B.n677 B.n289 585
R161 B.n677 B.n676 585
R162 B.n667 B.n290 585
R163 B.n291 B.n290 585
R164 B.n669 B.n668 585
R165 B.n670 B.n669 585
R166 B.n666 B.n296 585
R167 B.n296 B.n295 585
R168 B.n665 B.n664 585
R169 B.n664 B.n663 585
R170 B.n298 B.n297 585
R171 B.n299 B.n298 585
R172 B.n656 B.n655 585
R173 B.n657 B.n656 585
R174 B.n654 B.n304 585
R175 B.n304 B.n303 585
R176 B.n653 B.n652 585
R177 B.n652 B.n651 585
R178 B.n306 B.n305 585
R179 B.n307 B.n306 585
R180 B.n644 B.n643 585
R181 B.n645 B.n644 585
R182 B.n642 B.n312 585
R183 B.n312 B.n311 585
R184 B.n641 B.n640 585
R185 B.n640 B.n639 585
R186 B.n314 B.n313 585
R187 B.n315 B.n314 585
R188 B.n632 B.n631 585
R189 B.n633 B.n632 585
R190 B.n630 B.n320 585
R191 B.n320 B.n319 585
R192 B.n629 B.n628 585
R193 B.n628 B.n627 585
R194 B.n322 B.n321 585
R195 B.n323 B.n322 585
R196 B.n620 B.n619 585
R197 B.n621 B.n620 585
R198 B.n618 B.n328 585
R199 B.n328 B.n327 585
R200 B.n617 B.n616 585
R201 B.n616 B.n615 585
R202 B.n330 B.n329 585
R203 B.n331 B.n330 585
R204 B.n608 B.n607 585
R205 B.n609 B.n608 585
R206 B.n606 B.n336 585
R207 B.n336 B.n335 585
R208 B.n605 B.n604 585
R209 B.n604 B.n603 585
R210 B.n338 B.n337 585
R211 B.n339 B.n338 585
R212 B.n596 B.n595 585
R213 B.n597 B.n596 585
R214 B.n594 B.n344 585
R215 B.n344 B.n343 585
R216 B.n593 B.n592 585
R217 B.n592 B.n591 585
R218 B.n346 B.n345 585
R219 B.n347 B.n346 585
R220 B.n584 B.n583 585
R221 B.n585 B.n584 585
R222 B.n582 B.n352 585
R223 B.n352 B.n351 585
R224 B.n576 B.n575 585
R225 B.n574 B.n398 585
R226 B.n573 B.n397 585
R227 B.n578 B.n397 585
R228 B.n572 B.n571 585
R229 B.n570 B.n569 585
R230 B.n568 B.n567 585
R231 B.n566 B.n565 585
R232 B.n564 B.n563 585
R233 B.n562 B.n561 585
R234 B.n560 B.n559 585
R235 B.n558 B.n557 585
R236 B.n556 B.n555 585
R237 B.n554 B.n553 585
R238 B.n552 B.n551 585
R239 B.n550 B.n549 585
R240 B.n548 B.n547 585
R241 B.n546 B.n545 585
R242 B.n544 B.n543 585
R243 B.n542 B.n541 585
R244 B.n540 B.n539 585
R245 B.n538 B.n537 585
R246 B.n536 B.n535 585
R247 B.n534 B.n533 585
R248 B.n532 B.n531 585
R249 B.n530 B.n529 585
R250 B.n528 B.n527 585
R251 B.n526 B.n525 585
R252 B.n524 B.n523 585
R253 B.n522 B.n521 585
R254 B.n520 B.n519 585
R255 B.n518 B.n517 585
R256 B.n516 B.n515 585
R257 B.n514 B.n513 585
R258 B.n512 B.n511 585
R259 B.n510 B.n509 585
R260 B.n508 B.n507 585
R261 B.n506 B.n505 585
R262 B.n504 B.n503 585
R263 B.n502 B.n501 585
R264 B.n500 B.n499 585
R265 B.n497 B.n496 585
R266 B.n495 B.n494 585
R267 B.n493 B.n492 585
R268 B.n491 B.n490 585
R269 B.n489 B.n488 585
R270 B.n487 B.n486 585
R271 B.n485 B.n484 585
R272 B.n483 B.n482 585
R273 B.n481 B.n480 585
R274 B.n479 B.n478 585
R275 B.n477 B.n476 585
R276 B.n475 B.n474 585
R277 B.n473 B.n472 585
R278 B.n471 B.n470 585
R279 B.n469 B.n468 585
R280 B.n467 B.n466 585
R281 B.n465 B.n464 585
R282 B.n463 B.n462 585
R283 B.n461 B.n460 585
R284 B.n459 B.n458 585
R285 B.n457 B.n456 585
R286 B.n455 B.n454 585
R287 B.n453 B.n452 585
R288 B.n451 B.n450 585
R289 B.n449 B.n448 585
R290 B.n447 B.n446 585
R291 B.n445 B.n444 585
R292 B.n443 B.n442 585
R293 B.n441 B.n440 585
R294 B.n439 B.n438 585
R295 B.n437 B.n436 585
R296 B.n435 B.n434 585
R297 B.n433 B.n432 585
R298 B.n431 B.n430 585
R299 B.n429 B.n428 585
R300 B.n427 B.n426 585
R301 B.n425 B.n424 585
R302 B.n423 B.n422 585
R303 B.n421 B.n420 585
R304 B.n419 B.n418 585
R305 B.n417 B.n416 585
R306 B.n415 B.n414 585
R307 B.n413 B.n412 585
R308 B.n411 B.n410 585
R309 B.n409 B.n408 585
R310 B.n407 B.n406 585
R311 B.n405 B.n404 585
R312 B.n354 B.n353 585
R313 B.n581 B.n580 585
R314 B.n350 B.n349 585
R315 B.n351 B.n350 585
R316 B.n587 B.n586 585
R317 B.n586 B.n585 585
R318 B.n588 B.n348 585
R319 B.n348 B.n347 585
R320 B.n590 B.n589 585
R321 B.n591 B.n590 585
R322 B.n342 B.n341 585
R323 B.n343 B.n342 585
R324 B.n599 B.n598 585
R325 B.n598 B.n597 585
R326 B.n600 B.n340 585
R327 B.n340 B.n339 585
R328 B.n602 B.n601 585
R329 B.n603 B.n602 585
R330 B.n334 B.n333 585
R331 B.n335 B.n334 585
R332 B.n611 B.n610 585
R333 B.n610 B.n609 585
R334 B.n612 B.n332 585
R335 B.n332 B.n331 585
R336 B.n614 B.n613 585
R337 B.n615 B.n614 585
R338 B.n326 B.n325 585
R339 B.n327 B.n326 585
R340 B.n623 B.n622 585
R341 B.n622 B.n621 585
R342 B.n624 B.n324 585
R343 B.n324 B.n323 585
R344 B.n626 B.n625 585
R345 B.n627 B.n626 585
R346 B.n318 B.n317 585
R347 B.n319 B.n318 585
R348 B.n635 B.n634 585
R349 B.n634 B.n633 585
R350 B.n636 B.n316 585
R351 B.n316 B.n315 585
R352 B.n638 B.n637 585
R353 B.n639 B.n638 585
R354 B.n310 B.n309 585
R355 B.n311 B.n310 585
R356 B.n647 B.n646 585
R357 B.n646 B.n645 585
R358 B.n648 B.n308 585
R359 B.n308 B.n307 585
R360 B.n650 B.n649 585
R361 B.n651 B.n650 585
R362 B.n302 B.n301 585
R363 B.n303 B.n302 585
R364 B.n659 B.n658 585
R365 B.n658 B.n657 585
R366 B.n660 B.n300 585
R367 B.n300 B.n299 585
R368 B.n662 B.n661 585
R369 B.n663 B.n662 585
R370 B.n294 B.n293 585
R371 B.n295 B.n294 585
R372 B.n672 B.n671 585
R373 B.n671 B.n670 585
R374 B.n673 B.n292 585
R375 B.n292 B.n291 585
R376 B.n675 B.n674 585
R377 B.n676 B.n675 585
R378 B.n2 B.n0 585
R379 B.n4 B.n2 585
R380 B.n3 B.n1 585
R381 B.n789 B.n3 585
R382 B.n787 B.n786 585
R383 B.n788 B.n787 585
R384 B.n785 B.n9 585
R385 B.n9 B.n8 585
R386 B.n784 B.n783 585
R387 B.n783 B.n782 585
R388 B.n11 B.n10 585
R389 B.n781 B.n11 585
R390 B.n779 B.n778 585
R391 B.n780 B.n779 585
R392 B.n777 B.n16 585
R393 B.n16 B.n15 585
R394 B.n776 B.n775 585
R395 B.n775 B.n774 585
R396 B.n18 B.n17 585
R397 B.n773 B.n18 585
R398 B.n771 B.n770 585
R399 B.n772 B.n771 585
R400 B.n769 B.n23 585
R401 B.n23 B.n22 585
R402 B.n768 B.n767 585
R403 B.n767 B.n766 585
R404 B.n25 B.n24 585
R405 B.n765 B.n25 585
R406 B.n763 B.n762 585
R407 B.n764 B.n763 585
R408 B.n761 B.n30 585
R409 B.n30 B.n29 585
R410 B.n760 B.n759 585
R411 B.n759 B.n758 585
R412 B.n32 B.n31 585
R413 B.n757 B.n32 585
R414 B.n755 B.n754 585
R415 B.n756 B.n755 585
R416 B.n753 B.n37 585
R417 B.n37 B.n36 585
R418 B.n752 B.n751 585
R419 B.n751 B.n750 585
R420 B.n39 B.n38 585
R421 B.n749 B.n39 585
R422 B.n747 B.n746 585
R423 B.n748 B.n747 585
R424 B.n745 B.n44 585
R425 B.n44 B.n43 585
R426 B.n744 B.n743 585
R427 B.n743 B.n742 585
R428 B.n46 B.n45 585
R429 B.n741 B.n46 585
R430 B.n739 B.n738 585
R431 B.n740 B.n739 585
R432 B.n737 B.n51 585
R433 B.n51 B.n50 585
R434 B.n736 B.n735 585
R435 B.n735 B.n734 585
R436 B.n53 B.n52 585
R437 B.n733 B.n53 585
R438 B.n731 B.n730 585
R439 B.n732 B.n731 585
R440 B.n729 B.n58 585
R441 B.n58 B.n57 585
R442 B.n728 B.n727 585
R443 B.n727 B.n726 585
R444 B.n60 B.n59 585
R445 B.n725 B.n60 585
R446 B.n792 B.n791 585
R447 B.n791 B.n790 585
R448 B.n576 B.n350 511.721
R449 B.n113 B.n60 511.721
R450 B.n580 B.n352 511.721
R451 B.n723 B.n62 511.721
R452 B.n401 B.t8 353.108
R453 B.n108 B.t11 353.108
R454 B.n399 B.t5 353.108
R455 B.n110 B.t14 353.108
R456 B.n401 B.t6 279.152
R457 B.n399 B.t2 279.152
R458 B.n110 B.t13 279.152
R459 B.n108 B.t9 279.152
R460 B.n402 B.t7 270.683
R461 B.n109 B.t12 270.683
R462 B.n400 B.t4 270.683
R463 B.n111 B.t15 270.683
R464 B.n724 B.n106 256.663
R465 B.n724 B.n105 256.663
R466 B.n724 B.n104 256.663
R467 B.n724 B.n103 256.663
R468 B.n724 B.n102 256.663
R469 B.n724 B.n101 256.663
R470 B.n724 B.n100 256.663
R471 B.n724 B.n99 256.663
R472 B.n724 B.n98 256.663
R473 B.n724 B.n97 256.663
R474 B.n724 B.n96 256.663
R475 B.n724 B.n95 256.663
R476 B.n724 B.n94 256.663
R477 B.n724 B.n93 256.663
R478 B.n724 B.n92 256.663
R479 B.n724 B.n91 256.663
R480 B.n724 B.n90 256.663
R481 B.n724 B.n89 256.663
R482 B.n724 B.n88 256.663
R483 B.n724 B.n87 256.663
R484 B.n724 B.n86 256.663
R485 B.n724 B.n85 256.663
R486 B.n724 B.n84 256.663
R487 B.n724 B.n83 256.663
R488 B.n724 B.n82 256.663
R489 B.n724 B.n81 256.663
R490 B.n724 B.n80 256.663
R491 B.n724 B.n79 256.663
R492 B.n724 B.n78 256.663
R493 B.n724 B.n77 256.663
R494 B.n724 B.n76 256.663
R495 B.n724 B.n75 256.663
R496 B.n724 B.n74 256.663
R497 B.n724 B.n73 256.663
R498 B.n724 B.n72 256.663
R499 B.n724 B.n71 256.663
R500 B.n724 B.n70 256.663
R501 B.n724 B.n69 256.663
R502 B.n724 B.n68 256.663
R503 B.n724 B.n67 256.663
R504 B.n724 B.n66 256.663
R505 B.n724 B.n65 256.663
R506 B.n724 B.n64 256.663
R507 B.n724 B.n63 256.663
R508 B.n578 B.n577 256.663
R509 B.n578 B.n355 256.663
R510 B.n578 B.n356 256.663
R511 B.n578 B.n357 256.663
R512 B.n578 B.n358 256.663
R513 B.n578 B.n359 256.663
R514 B.n578 B.n360 256.663
R515 B.n578 B.n361 256.663
R516 B.n578 B.n362 256.663
R517 B.n578 B.n363 256.663
R518 B.n578 B.n364 256.663
R519 B.n578 B.n365 256.663
R520 B.n578 B.n366 256.663
R521 B.n578 B.n367 256.663
R522 B.n578 B.n368 256.663
R523 B.n578 B.n369 256.663
R524 B.n578 B.n370 256.663
R525 B.n578 B.n371 256.663
R526 B.n578 B.n372 256.663
R527 B.n578 B.n373 256.663
R528 B.n578 B.n374 256.663
R529 B.n578 B.n375 256.663
R530 B.n578 B.n376 256.663
R531 B.n578 B.n377 256.663
R532 B.n578 B.n378 256.663
R533 B.n578 B.n379 256.663
R534 B.n578 B.n380 256.663
R535 B.n578 B.n381 256.663
R536 B.n578 B.n382 256.663
R537 B.n578 B.n383 256.663
R538 B.n578 B.n384 256.663
R539 B.n578 B.n385 256.663
R540 B.n578 B.n386 256.663
R541 B.n578 B.n387 256.663
R542 B.n578 B.n388 256.663
R543 B.n578 B.n389 256.663
R544 B.n578 B.n390 256.663
R545 B.n578 B.n391 256.663
R546 B.n578 B.n392 256.663
R547 B.n578 B.n393 256.663
R548 B.n578 B.n394 256.663
R549 B.n578 B.n395 256.663
R550 B.n578 B.n396 256.663
R551 B.n579 B.n578 256.663
R552 B.n586 B.n350 163.367
R553 B.n586 B.n348 163.367
R554 B.n590 B.n348 163.367
R555 B.n590 B.n342 163.367
R556 B.n598 B.n342 163.367
R557 B.n598 B.n340 163.367
R558 B.n602 B.n340 163.367
R559 B.n602 B.n334 163.367
R560 B.n610 B.n334 163.367
R561 B.n610 B.n332 163.367
R562 B.n614 B.n332 163.367
R563 B.n614 B.n326 163.367
R564 B.n622 B.n326 163.367
R565 B.n622 B.n324 163.367
R566 B.n626 B.n324 163.367
R567 B.n626 B.n318 163.367
R568 B.n634 B.n318 163.367
R569 B.n634 B.n316 163.367
R570 B.n638 B.n316 163.367
R571 B.n638 B.n310 163.367
R572 B.n646 B.n310 163.367
R573 B.n646 B.n308 163.367
R574 B.n650 B.n308 163.367
R575 B.n650 B.n302 163.367
R576 B.n658 B.n302 163.367
R577 B.n658 B.n300 163.367
R578 B.n662 B.n300 163.367
R579 B.n662 B.n294 163.367
R580 B.n671 B.n294 163.367
R581 B.n671 B.n292 163.367
R582 B.n675 B.n292 163.367
R583 B.n675 B.n2 163.367
R584 B.n791 B.n2 163.367
R585 B.n791 B.n3 163.367
R586 B.n787 B.n3 163.367
R587 B.n787 B.n9 163.367
R588 B.n783 B.n9 163.367
R589 B.n783 B.n11 163.367
R590 B.n779 B.n11 163.367
R591 B.n779 B.n16 163.367
R592 B.n775 B.n16 163.367
R593 B.n775 B.n18 163.367
R594 B.n771 B.n18 163.367
R595 B.n771 B.n23 163.367
R596 B.n767 B.n23 163.367
R597 B.n767 B.n25 163.367
R598 B.n763 B.n25 163.367
R599 B.n763 B.n30 163.367
R600 B.n759 B.n30 163.367
R601 B.n759 B.n32 163.367
R602 B.n755 B.n32 163.367
R603 B.n755 B.n37 163.367
R604 B.n751 B.n37 163.367
R605 B.n751 B.n39 163.367
R606 B.n747 B.n39 163.367
R607 B.n747 B.n44 163.367
R608 B.n743 B.n44 163.367
R609 B.n743 B.n46 163.367
R610 B.n739 B.n46 163.367
R611 B.n739 B.n51 163.367
R612 B.n735 B.n51 163.367
R613 B.n735 B.n53 163.367
R614 B.n731 B.n53 163.367
R615 B.n731 B.n58 163.367
R616 B.n727 B.n58 163.367
R617 B.n727 B.n60 163.367
R618 B.n398 B.n397 163.367
R619 B.n571 B.n397 163.367
R620 B.n569 B.n568 163.367
R621 B.n565 B.n564 163.367
R622 B.n561 B.n560 163.367
R623 B.n557 B.n556 163.367
R624 B.n553 B.n552 163.367
R625 B.n549 B.n548 163.367
R626 B.n545 B.n544 163.367
R627 B.n541 B.n540 163.367
R628 B.n537 B.n536 163.367
R629 B.n533 B.n532 163.367
R630 B.n529 B.n528 163.367
R631 B.n525 B.n524 163.367
R632 B.n521 B.n520 163.367
R633 B.n517 B.n516 163.367
R634 B.n513 B.n512 163.367
R635 B.n509 B.n508 163.367
R636 B.n505 B.n504 163.367
R637 B.n501 B.n500 163.367
R638 B.n496 B.n495 163.367
R639 B.n492 B.n491 163.367
R640 B.n488 B.n487 163.367
R641 B.n484 B.n483 163.367
R642 B.n480 B.n479 163.367
R643 B.n476 B.n475 163.367
R644 B.n472 B.n471 163.367
R645 B.n468 B.n467 163.367
R646 B.n464 B.n463 163.367
R647 B.n460 B.n459 163.367
R648 B.n456 B.n455 163.367
R649 B.n452 B.n451 163.367
R650 B.n448 B.n447 163.367
R651 B.n444 B.n443 163.367
R652 B.n440 B.n439 163.367
R653 B.n436 B.n435 163.367
R654 B.n432 B.n431 163.367
R655 B.n428 B.n427 163.367
R656 B.n424 B.n423 163.367
R657 B.n420 B.n419 163.367
R658 B.n416 B.n415 163.367
R659 B.n412 B.n411 163.367
R660 B.n408 B.n407 163.367
R661 B.n404 B.n354 163.367
R662 B.n584 B.n352 163.367
R663 B.n584 B.n346 163.367
R664 B.n592 B.n346 163.367
R665 B.n592 B.n344 163.367
R666 B.n596 B.n344 163.367
R667 B.n596 B.n338 163.367
R668 B.n604 B.n338 163.367
R669 B.n604 B.n336 163.367
R670 B.n608 B.n336 163.367
R671 B.n608 B.n330 163.367
R672 B.n616 B.n330 163.367
R673 B.n616 B.n328 163.367
R674 B.n620 B.n328 163.367
R675 B.n620 B.n322 163.367
R676 B.n628 B.n322 163.367
R677 B.n628 B.n320 163.367
R678 B.n632 B.n320 163.367
R679 B.n632 B.n314 163.367
R680 B.n640 B.n314 163.367
R681 B.n640 B.n312 163.367
R682 B.n644 B.n312 163.367
R683 B.n644 B.n306 163.367
R684 B.n652 B.n306 163.367
R685 B.n652 B.n304 163.367
R686 B.n656 B.n304 163.367
R687 B.n656 B.n298 163.367
R688 B.n664 B.n298 163.367
R689 B.n664 B.n296 163.367
R690 B.n669 B.n296 163.367
R691 B.n669 B.n290 163.367
R692 B.n677 B.n290 163.367
R693 B.n678 B.n677 163.367
R694 B.n678 B.n5 163.367
R695 B.n6 B.n5 163.367
R696 B.n7 B.n6 163.367
R697 B.n683 B.n7 163.367
R698 B.n683 B.n12 163.367
R699 B.n13 B.n12 163.367
R700 B.n14 B.n13 163.367
R701 B.n688 B.n14 163.367
R702 B.n688 B.n19 163.367
R703 B.n20 B.n19 163.367
R704 B.n21 B.n20 163.367
R705 B.n693 B.n21 163.367
R706 B.n693 B.n26 163.367
R707 B.n27 B.n26 163.367
R708 B.n28 B.n27 163.367
R709 B.n698 B.n28 163.367
R710 B.n698 B.n33 163.367
R711 B.n34 B.n33 163.367
R712 B.n35 B.n34 163.367
R713 B.n703 B.n35 163.367
R714 B.n703 B.n40 163.367
R715 B.n41 B.n40 163.367
R716 B.n42 B.n41 163.367
R717 B.n708 B.n42 163.367
R718 B.n708 B.n47 163.367
R719 B.n48 B.n47 163.367
R720 B.n49 B.n48 163.367
R721 B.n713 B.n49 163.367
R722 B.n713 B.n54 163.367
R723 B.n55 B.n54 163.367
R724 B.n56 B.n55 163.367
R725 B.n718 B.n56 163.367
R726 B.n718 B.n61 163.367
R727 B.n62 B.n61 163.367
R728 B.n117 B.n116 163.367
R729 B.n121 B.n120 163.367
R730 B.n125 B.n124 163.367
R731 B.n129 B.n128 163.367
R732 B.n133 B.n132 163.367
R733 B.n137 B.n136 163.367
R734 B.n141 B.n140 163.367
R735 B.n145 B.n144 163.367
R736 B.n149 B.n148 163.367
R737 B.n153 B.n152 163.367
R738 B.n157 B.n156 163.367
R739 B.n161 B.n160 163.367
R740 B.n165 B.n164 163.367
R741 B.n169 B.n168 163.367
R742 B.n173 B.n172 163.367
R743 B.n177 B.n176 163.367
R744 B.n181 B.n180 163.367
R745 B.n185 B.n184 163.367
R746 B.n189 B.n188 163.367
R747 B.n193 B.n192 163.367
R748 B.n197 B.n196 163.367
R749 B.n201 B.n200 163.367
R750 B.n205 B.n204 163.367
R751 B.n209 B.n208 163.367
R752 B.n214 B.n213 163.367
R753 B.n218 B.n217 163.367
R754 B.n222 B.n221 163.367
R755 B.n226 B.n225 163.367
R756 B.n230 B.n229 163.367
R757 B.n234 B.n233 163.367
R758 B.n238 B.n237 163.367
R759 B.n242 B.n241 163.367
R760 B.n246 B.n245 163.367
R761 B.n250 B.n249 163.367
R762 B.n254 B.n253 163.367
R763 B.n258 B.n257 163.367
R764 B.n262 B.n261 163.367
R765 B.n266 B.n265 163.367
R766 B.n270 B.n269 163.367
R767 B.n274 B.n273 163.367
R768 B.n278 B.n277 163.367
R769 B.n282 B.n281 163.367
R770 B.n286 B.n285 163.367
R771 B.n723 B.n107 163.367
R772 B.n578 B.n351 86.7294
R773 B.n725 B.n724 86.7294
R774 B.n402 B.n401 82.4247
R775 B.n400 B.n399 82.4247
R776 B.n111 B.n110 82.4247
R777 B.n109 B.n108 82.4247
R778 B.n577 B.n576 71.676
R779 B.n571 B.n355 71.676
R780 B.n568 B.n356 71.676
R781 B.n564 B.n357 71.676
R782 B.n560 B.n358 71.676
R783 B.n556 B.n359 71.676
R784 B.n552 B.n360 71.676
R785 B.n548 B.n361 71.676
R786 B.n544 B.n362 71.676
R787 B.n540 B.n363 71.676
R788 B.n536 B.n364 71.676
R789 B.n532 B.n365 71.676
R790 B.n528 B.n366 71.676
R791 B.n524 B.n367 71.676
R792 B.n520 B.n368 71.676
R793 B.n516 B.n369 71.676
R794 B.n512 B.n370 71.676
R795 B.n508 B.n371 71.676
R796 B.n504 B.n372 71.676
R797 B.n500 B.n373 71.676
R798 B.n495 B.n374 71.676
R799 B.n491 B.n375 71.676
R800 B.n487 B.n376 71.676
R801 B.n483 B.n377 71.676
R802 B.n479 B.n378 71.676
R803 B.n475 B.n379 71.676
R804 B.n471 B.n380 71.676
R805 B.n467 B.n381 71.676
R806 B.n463 B.n382 71.676
R807 B.n459 B.n383 71.676
R808 B.n455 B.n384 71.676
R809 B.n451 B.n385 71.676
R810 B.n447 B.n386 71.676
R811 B.n443 B.n387 71.676
R812 B.n439 B.n388 71.676
R813 B.n435 B.n389 71.676
R814 B.n431 B.n390 71.676
R815 B.n427 B.n391 71.676
R816 B.n423 B.n392 71.676
R817 B.n419 B.n393 71.676
R818 B.n415 B.n394 71.676
R819 B.n411 B.n395 71.676
R820 B.n407 B.n396 71.676
R821 B.n579 B.n354 71.676
R822 B.n113 B.n63 71.676
R823 B.n117 B.n64 71.676
R824 B.n121 B.n65 71.676
R825 B.n125 B.n66 71.676
R826 B.n129 B.n67 71.676
R827 B.n133 B.n68 71.676
R828 B.n137 B.n69 71.676
R829 B.n141 B.n70 71.676
R830 B.n145 B.n71 71.676
R831 B.n149 B.n72 71.676
R832 B.n153 B.n73 71.676
R833 B.n157 B.n74 71.676
R834 B.n161 B.n75 71.676
R835 B.n165 B.n76 71.676
R836 B.n169 B.n77 71.676
R837 B.n173 B.n78 71.676
R838 B.n177 B.n79 71.676
R839 B.n181 B.n80 71.676
R840 B.n185 B.n81 71.676
R841 B.n189 B.n82 71.676
R842 B.n193 B.n83 71.676
R843 B.n197 B.n84 71.676
R844 B.n201 B.n85 71.676
R845 B.n205 B.n86 71.676
R846 B.n209 B.n87 71.676
R847 B.n214 B.n88 71.676
R848 B.n218 B.n89 71.676
R849 B.n222 B.n90 71.676
R850 B.n226 B.n91 71.676
R851 B.n230 B.n92 71.676
R852 B.n234 B.n93 71.676
R853 B.n238 B.n94 71.676
R854 B.n242 B.n95 71.676
R855 B.n246 B.n96 71.676
R856 B.n250 B.n97 71.676
R857 B.n254 B.n98 71.676
R858 B.n258 B.n99 71.676
R859 B.n262 B.n100 71.676
R860 B.n266 B.n101 71.676
R861 B.n270 B.n102 71.676
R862 B.n274 B.n103 71.676
R863 B.n278 B.n104 71.676
R864 B.n282 B.n105 71.676
R865 B.n286 B.n106 71.676
R866 B.n107 B.n106 71.676
R867 B.n285 B.n105 71.676
R868 B.n281 B.n104 71.676
R869 B.n277 B.n103 71.676
R870 B.n273 B.n102 71.676
R871 B.n269 B.n101 71.676
R872 B.n265 B.n100 71.676
R873 B.n261 B.n99 71.676
R874 B.n257 B.n98 71.676
R875 B.n253 B.n97 71.676
R876 B.n249 B.n96 71.676
R877 B.n245 B.n95 71.676
R878 B.n241 B.n94 71.676
R879 B.n237 B.n93 71.676
R880 B.n233 B.n92 71.676
R881 B.n229 B.n91 71.676
R882 B.n225 B.n90 71.676
R883 B.n221 B.n89 71.676
R884 B.n217 B.n88 71.676
R885 B.n213 B.n87 71.676
R886 B.n208 B.n86 71.676
R887 B.n204 B.n85 71.676
R888 B.n200 B.n84 71.676
R889 B.n196 B.n83 71.676
R890 B.n192 B.n82 71.676
R891 B.n188 B.n81 71.676
R892 B.n184 B.n80 71.676
R893 B.n180 B.n79 71.676
R894 B.n176 B.n78 71.676
R895 B.n172 B.n77 71.676
R896 B.n168 B.n76 71.676
R897 B.n164 B.n75 71.676
R898 B.n160 B.n74 71.676
R899 B.n156 B.n73 71.676
R900 B.n152 B.n72 71.676
R901 B.n148 B.n71 71.676
R902 B.n144 B.n70 71.676
R903 B.n140 B.n69 71.676
R904 B.n136 B.n68 71.676
R905 B.n132 B.n67 71.676
R906 B.n128 B.n66 71.676
R907 B.n124 B.n65 71.676
R908 B.n120 B.n64 71.676
R909 B.n116 B.n63 71.676
R910 B.n577 B.n398 71.676
R911 B.n569 B.n355 71.676
R912 B.n565 B.n356 71.676
R913 B.n561 B.n357 71.676
R914 B.n557 B.n358 71.676
R915 B.n553 B.n359 71.676
R916 B.n549 B.n360 71.676
R917 B.n545 B.n361 71.676
R918 B.n541 B.n362 71.676
R919 B.n537 B.n363 71.676
R920 B.n533 B.n364 71.676
R921 B.n529 B.n365 71.676
R922 B.n525 B.n366 71.676
R923 B.n521 B.n367 71.676
R924 B.n517 B.n368 71.676
R925 B.n513 B.n369 71.676
R926 B.n509 B.n370 71.676
R927 B.n505 B.n371 71.676
R928 B.n501 B.n372 71.676
R929 B.n496 B.n373 71.676
R930 B.n492 B.n374 71.676
R931 B.n488 B.n375 71.676
R932 B.n484 B.n376 71.676
R933 B.n480 B.n377 71.676
R934 B.n476 B.n378 71.676
R935 B.n472 B.n379 71.676
R936 B.n468 B.n380 71.676
R937 B.n464 B.n381 71.676
R938 B.n460 B.n382 71.676
R939 B.n456 B.n383 71.676
R940 B.n452 B.n384 71.676
R941 B.n448 B.n385 71.676
R942 B.n444 B.n386 71.676
R943 B.n440 B.n387 71.676
R944 B.n436 B.n388 71.676
R945 B.n432 B.n389 71.676
R946 B.n428 B.n390 71.676
R947 B.n424 B.n391 71.676
R948 B.n420 B.n392 71.676
R949 B.n416 B.n393 71.676
R950 B.n412 B.n394 71.676
R951 B.n408 B.n395 71.676
R952 B.n404 B.n396 71.676
R953 B.n580 B.n579 71.676
R954 B.n403 B.n402 59.5399
R955 B.n498 B.n400 59.5399
R956 B.n112 B.n111 59.5399
R957 B.n211 B.n109 59.5399
R958 B.n585 B.n351 45.0201
R959 B.n585 B.n347 45.0201
R960 B.n591 B.n347 45.0201
R961 B.n591 B.n343 45.0201
R962 B.n597 B.n343 45.0201
R963 B.n597 B.n339 45.0201
R964 B.n603 B.n339 45.0201
R965 B.n603 B.n335 45.0201
R966 B.n609 B.n335 45.0201
R967 B.n615 B.n331 45.0201
R968 B.n615 B.n327 45.0201
R969 B.n621 B.n327 45.0201
R970 B.n621 B.n323 45.0201
R971 B.n627 B.n323 45.0201
R972 B.n627 B.n319 45.0201
R973 B.n633 B.n319 45.0201
R974 B.n633 B.n315 45.0201
R975 B.n639 B.n315 45.0201
R976 B.n639 B.n311 45.0201
R977 B.n645 B.n311 45.0201
R978 B.n645 B.n307 45.0201
R979 B.n651 B.n307 45.0201
R980 B.n651 B.n303 45.0201
R981 B.n657 B.n303 45.0201
R982 B.n663 B.n299 45.0201
R983 B.n663 B.n295 45.0201
R984 B.n670 B.n295 45.0201
R985 B.n670 B.n291 45.0201
R986 B.n676 B.n291 45.0201
R987 B.n676 B.n4 45.0201
R988 B.n790 B.n4 45.0201
R989 B.n790 B.n789 45.0201
R990 B.n789 B.n788 45.0201
R991 B.n788 B.n8 45.0201
R992 B.n782 B.n8 45.0201
R993 B.n782 B.n781 45.0201
R994 B.n781 B.n780 45.0201
R995 B.n780 B.n15 45.0201
R996 B.n774 B.n773 45.0201
R997 B.n773 B.n772 45.0201
R998 B.n772 B.n22 45.0201
R999 B.n766 B.n22 45.0201
R1000 B.n766 B.n765 45.0201
R1001 B.n765 B.n764 45.0201
R1002 B.n764 B.n29 45.0201
R1003 B.n758 B.n29 45.0201
R1004 B.n758 B.n757 45.0201
R1005 B.n757 B.n756 45.0201
R1006 B.n756 B.n36 45.0201
R1007 B.n750 B.n36 45.0201
R1008 B.n750 B.n749 45.0201
R1009 B.n749 B.n748 45.0201
R1010 B.n748 B.n43 45.0201
R1011 B.n742 B.n741 45.0201
R1012 B.n741 B.n740 45.0201
R1013 B.n740 B.n50 45.0201
R1014 B.n734 B.n50 45.0201
R1015 B.n734 B.n733 45.0201
R1016 B.n733 B.n732 45.0201
R1017 B.n732 B.n57 45.0201
R1018 B.n726 B.n57 45.0201
R1019 B.n726 B.n725 45.0201
R1020 B.t0 B.n299 38.3995
R1021 B.t1 B.n15 38.3995
R1022 B.n114 B.n59 33.2493
R1023 B.n722 B.n721 33.2493
R1024 B.n582 B.n581 33.2493
R1025 B.n575 B.n349 33.2493
R1026 B.t3 B.n331 25.1585
R1027 B.t10 B.n43 25.1585
R1028 B.n609 B.t3 19.8621
R1029 B.n742 B.t10 19.8621
R1030 B B.n792 18.0485
R1031 B.n115 B.n114 10.6151
R1032 B.n118 B.n115 10.6151
R1033 B.n119 B.n118 10.6151
R1034 B.n122 B.n119 10.6151
R1035 B.n123 B.n122 10.6151
R1036 B.n126 B.n123 10.6151
R1037 B.n127 B.n126 10.6151
R1038 B.n130 B.n127 10.6151
R1039 B.n131 B.n130 10.6151
R1040 B.n134 B.n131 10.6151
R1041 B.n135 B.n134 10.6151
R1042 B.n138 B.n135 10.6151
R1043 B.n139 B.n138 10.6151
R1044 B.n142 B.n139 10.6151
R1045 B.n143 B.n142 10.6151
R1046 B.n146 B.n143 10.6151
R1047 B.n147 B.n146 10.6151
R1048 B.n150 B.n147 10.6151
R1049 B.n151 B.n150 10.6151
R1050 B.n154 B.n151 10.6151
R1051 B.n155 B.n154 10.6151
R1052 B.n158 B.n155 10.6151
R1053 B.n159 B.n158 10.6151
R1054 B.n162 B.n159 10.6151
R1055 B.n163 B.n162 10.6151
R1056 B.n166 B.n163 10.6151
R1057 B.n167 B.n166 10.6151
R1058 B.n170 B.n167 10.6151
R1059 B.n171 B.n170 10.6151
R1060 B.n174 B.n171 10.6151
R1061 B.n175 B.n174 10.6151
R1062 B.n178 B.n175 10.6151
R1063 B.n179 B.n178 10.6151
R1064 B.n182 B.n179 10.6151
R1065 B.n183 B.n182 10.6151
R1066 B.n186 B.n183 10.6151
R1067 B.n187 B.n186 10.6151
R1068 B.n190 B.n187 10.6151
R1069 B.n191 B.n190 10.6151
R1070 B.n195 B.n194 10.6151
R1071 B.n198 B.n195 10.6151
R1072 B.n199 B.n198 10.6151
R1073 B.n202 B.n199 10.6151
R1074 B.n203 B.n202 10.6151
R1075 B.n206 B.n203 10.6151
R1076 B.n207 B.n206 10.6151
R1077 B.n210 B.n207 10.6151
R1078 B.n215 B.n212 10.6151
R1079 B.n216 B.n215 10.6151
R1080 B.n219 B.n216 10.6151
R1081 B.n220 B.n219 10.6151
R1082 B.n223 B.n220 10.6151
R1083 B.n224 B.n223 10.6151
R1084 B.n227 B.n224 10.6151
R1085 B.n228 B.n227 10.6151
R1086 B.n231 B.n228 10.6151
R1087 B.n232 B.n231 10.6151
R1088 B.n235 B.n232 10.6151
R1089 B.n236 B.n235 10.6151
R1090 B.n239 B.n236 10.6151
R1091 B.n240 B.n239 10.6151
R1092 B.n243 B.n240 10.6151
R1093 B.n244 B.n243 10.6151
R1094 B.n247 B.n244 10.6151
R1095 B.n248 B.n247 10.6151
R1096 B.n251 B.n248 10.6151
R1097 B.n252 B.n251 10.6151
R1098 B.n255 B.n252 10.6151
R1099 B.n256 B.n255 10.6151
R1100 B.n259 B.n256 10.6151
R1101 B.n260 B.n259 10.6151
R1102 B.n263 B.n260 10.6151
R1103 B.n264 B.n263 10.6151
R1104 B.n267 B.n264 10.6151
R1105 B.n268 B.n267 10.6151
R1106 B.n271 B.n268 10.6151
R1107 B.n272 B.n271 10.6151
R1108 B.n275 B.n272 10.6151
R1109 B.n276 B.n275 10.6151
R1110 B.n279 B.n276 10.6151
R1111 B.n280 B.n279 10.6151
R1112 B.n283 B.n280 10.6151
R1113 B.n284 B.n283 10.6151
R1114 B.n287 B.n284 10.6151
R1115 B.n288 B.n287 10.6151
R1116 B.n722 B.n288 10.6151
R1117 B.n583 B.n582 10.6151
R1118 B.n583 B.n345 10.6151
R1119 B.n593 B.n345 10.6151
R1120 B.n594 B.n593 10.6151
R1121 B.n595 B.n594 10.6151
R1122 B.n595 B.n337 10.6151
R1123 B.n605 B.n337 10.6151
R1124 B.n606 B.n605 10.6151
R1125 B.n607 B.n606 10.6151
R1126 B.n607 B.n329 10.6151
R1127 B.n617 B.n329 10.6151
R1128 B.n618 B.n617 10.6151
R1129 B.n619 B.n618 10.6151
R1130 B.n619 B.n321 10.6151
R1131 B.n629 B.n321 10.6151
R1132 B.n630 B.n629 10.6151
R1133 B.n631 B.n630 10.6151
R1134 B.n631 B.n313 10.6151
R1135 B.n641 B.n313 10.6151
R1136 B.n642 B.n641 10.6151
R1137 B.n643 B.n642 10.6151
R1138 B.n643 B.n305 10.6151
R1139 B.n653 B.n305 10.6151
R1140 B.n654 B.n653 10.6151
R1141 B.n655 B.n654 10.6151
R1142 B.n655 B.n297 10.6151
R1143 B.n665 B.n297 10.6151
R1144 B.n666 B.n665 10.6151
R1145 B.n668 B.n666 10.6151
R1146 B.n668 B.n667 10.6151
R1147 B.n667 B.n289 10.6151
R1148 B.n679 B.n289 10.6151
R1149 B.n680 B.n679 10.6151
R1150 B.n681 B.n680 10.6151
R1151 B.n682 B.n681 10.6151
R1152 B.n684 B.n682 10.6151
R1153 B.n685 B.n684 10.6151
R1154 B.n686 B.n685 10.6151
R1155 B.n687 B.n686 10.6151
R1156 B.n689 B.n687 10.6151
R1157 B.n690 B.n689 10.6151
R1158 B.n691 B.n690 10.6151
R1159 B.n692 B.n691 10.6151
R1160 B.n694 B.n692 10.6151
R1161 B.n695 B.n694 10.6151
R1162 B.n696 B.n695 10.6151
R1163 B.n697 B.n696 10.6151
R1164 B.n699 B.n697 10.6151
R1165 B.n700 B.n699 10.6151
R1166 B.n701 B.n700 10.6151
R1167 B.n702 B.n701 10.6151
R1168 B.n704 B.n702 10.6151
R1169 B.n705 B.n704 10.6151
R1170 B.n706 B.n705 10.6151
R1171 B.n707 B.n706 10.6151
R1172 B.n709 B.n707 10.6151
R1173 B.n710 B.n709 10.6151
R1174 B.n711 B.n710 10.6151
R1175 B.n712 B.n711 10.6151
R1176 B.n714 B.n712 10.6151
R1177 B.n715 B.n714 10.6151
R1178 B.n716 B.n715 10.6151
R1179 B.n717 B.n716 10.6151
R1180 B.n719 B.n717 10.6151
R1181 B.n720 B.n719 10.6151
R1182 B.n721 B.n720 10.6151
R1183 B.n575 B.n574 10.6151
R1184 B.n574 B.n573 10.6151
R1185 B.n573 B.n572 10.6151
R1186 B.n572 B.n570 10.6151
R1187 B.n570 B.n567 10.6151
R1188 B.n567 B.n566 10.6151
R1189 B.n566 B.n563 10.6151
R1190 B.n563 B.n562 10.6151
R1191 B.n562 B.n559 10.6151
R1192 B.n559 B.n558 10.6151
R1193 B.n558 B.n555 10.6151
R1194 B.n555 B.n554 10.6151
R1195 B.n554 B.n551 10.6151
R1196 B.n551 B.n550 10.6151
R1197 B.n550 B.n547 10.6151
R1198 B.n547 B.n546 10.6151
R1199 B.n546 B.n543 10.6151
R1200 B.n543 B.n542 10.6151
R1201 B.n542 B.n539 10.6151
R1202 B.n539 B.n538 10.6151
R1203 B.n538 B.n535 10.6151
R1204 B.n535 B.n534 10.6151
R1205 B.n534 B.n531 10.6151
R1206 B.n531 B.n530 10.6151
R1207 B.n530 B.n527 10.6151
R1208 B.n527 B.n526 10.6151
R1209 B.n526 B.n523 10.6151
R1210 B.n523 B.n522 10.6151
R1211 B.n522 B.n519 10.6151
R1212 B.n519 B.n518 10.6151
R1213 B.n518 B.n515 10.6151
R1214 B.n515 B.n514 10.6151
R1215 B.n514 B.n511 10.6151
R1216 B.n511 B.n510 10.6151
R1217 B.n510 B.n507 10.6151
R1218 B.n507 B.n506 10.6151
R1219 B.n506 B.n503 10.6151
R1220 B.n503 B.n502 10.6151
R1221 B.n502 B.n499 10.6151
R1222 B.n497 B.n494 10.6151
R1223 B.n494 B.n493 10.6151
R1224 B.n493 B.n490 10.6151
R1225 B.n490 B.n489 10.6151
R1226 B.n489 B.n486 10.6151
R1227 B.n486 B.n485 10.6151
R1228 B.n485 B.n482 10.6151
R1229 B.n482 B.n481 10.6151
R1230 B.n478 B.n477 10.6151
R1231 B.n477 B.n474 10.6151
R1232 B.n474 B.n473 10.6151
R1233 B.n473 B.n470 10.6151
R1234 B.n470 B.n469 10.6151
R1235 B.n469 B.n466 10.6151
R1236 B.n466 B.n465 10.6151
R1237 B.n465 B.n462 10.6151
R1238 B.n462 B.n461 10.6151
R1239 B.n461 B.n458 10.6151
R1240 B.n458 B.n457 10.6151
R1241 B.n457 B.n454 10.6151
R1242 B.n454 B.n453 10.6151
R1243 B.n453 B.n450 10.6151
R1244 B.n450 B.n449 10.6151
R1245 B.n449 B.n446 10.6151
R1246 B.n446 B.n445 10.6151
R1247 B.n445 B.n442 10.6151
R1248 B.n442 B.n441 10.6151
R1249 B.n441 B.n438 10.6151
R1250 B.n438 B.n437 10.6151
R1251 B.n437 B.n434 10.6151
R1252 B.n434 B.n433 10.6151
R1253 B.n433 B.n430 10.6151
R1254 B.n430 B.n429 10.6151
R1255 B.n429 B.n426 10.6151
R1256 B.n426 B.n425 10.6151
R1257 B.n425 B.n422 10.6151
R1258 B.n422 B.n421 10.6151
R1259 B.n421 B.n418 10.6151
R1260 B.n418 B.n417 10.6151
R1261 B.n417 B.n414 10.6151
R1262 B.n414 B.n413 10.6151
R1263 B.n413 B.n410 10.6151
R1264 B.n410 B.n409 10.6151
R1265 B.n409 B.n406 10.6151
R1266 B.n406 B.n405 10.6151
R1267 B.n405 B.n353 10.6151
R1268 B.n581 B.n353 10.6151
R1269 B.n587 B.n349 10.6151
R1270 B.n588 B.n587 10.6151
R1271 B.n589 B.n588 10.6151
R1272 B.n589 B.n341 10.6151
R1273 B.n599 B.n341 10.6151
R1274 B.n600 B.n599 10.6151
R1275 B.n601 B.n600 10.6151
R1276 B.n601 B.n333 10.6151
R1277 B.n611 B.n333 10.6151
R1278 B.n612 B.n611 10.6151
R1279 B.n613 B.n612 10.6151
R1280 B.n613 B.n325 10.6151
R1281 B.n623 B.n325 10.6151
R1282 B.n624 B.n623 10.6151
R1283 B.n625 B.n624 10.6151
R1284 B.n625 B.n317 10.6151
R1285 B.n635 B.n317 10.6151
R1286 B.n636 B.n635 10.6151
R1287 B.n637 B.n636 10.6151
R1288 B.n637 B.n309 10.6151
R1289 B.n647 B.n309 10.6151
R1290 B.n648 B.n647 10.6151
R1291 B.n649 B.n648 10.6151
R1292 B.n649 B.n301 10.6151
R1293 B.n659 B.n301 10.6151
R1294 B.n660 B.n659 10.6151
R1295 B.n661 B.n660 10.6151
R1296 B.n661 B.n293 10.6151
R1297 B.n672 B.n293 10.6151
R1298 B.n673 B.n672 10.6151
R1299 B.n674 B.n673 10.6151
R1300 B.n674 B.n0 10.6151
R1301 B.n786 B.n1 10.6151
R1302 B.n786 B.n785 10.6151
R1303 B.n785 B.n784 10.6151
R1304 B.n784 B.n10 10.6151
R1305 B.n778 B.n10 10.6151
R1306 B.n778 B.n777 10.6151
R1307 B.n777 B.n776 10.6151
R1308 B.n776 B.n17 10.6151
R1309 B.n770 B.n17 10.6151
R1310 B.n770 B.n769 10.6151
R1311 B.n769 B.n768 10.6151
R1312 B.n768 B.n24 10.6151
R1313 B.n762 B.n24 10.6151
R1314 B.n762 B.n761 10.6151
R1315 B.n761 B.n760 10.6151
R1316 B.n760 B.n31 10.6151
R1317 B.n754 B.n31 10.6151
R1318 B.n754 B.n753 10.6151
R1319 B.n753 B.n752 10.6151
R1320 B.n752 B.n38 10.6151
R1321 B.n746 B.n38 10.6151
R1322 B.n746 B.n745 10.6151
R1323 B.n745 B.n744 10.6151
R1324 B.n744 B.n45 10.6151
R1325 B.n738 B.n45 10.6151
R1326 B.n738 B.n737 10.6151
R1327 B.n737 B.n736 10.6151
R1328 B.n736 B.n52 10.6151
R1329 B.n730 B.n52 10.6151
R1330 B.n730 B.n729 10.6151
R1331 B.n729 B.n728 10.6151
R1332 B.n728 B.n59 10.6151
R1333 B.n657 B.t0 6.62102
R1334 B.n774 B.t1 6.62102
R1335 B.n194 B.n112 6.5566
R1336 B.n211 B.n210 6.5566
R1337 B.n498 B.n497 6.5566
R1338 B.n481 B.n403 6.5566
R1339 B.n191 B.n112 4.05904
R1340 B.n212 B.n211 4.05904
R1341 B.n499 B.n498 4.05904
R1342 B.n478 B.n403 4.05904
R1343 B.n792 B.n0 2.81026
R1344 B.n792 B.n1 2.81026
R1345 VN VN.t1 152.28
R1346 VN VN.t0 105.43
R1347 VTAIL.n242 VTAIL.n186 289.615
R1348 VTAIL.n56 VTAIL.n0 289.615
R1349 VTAIL.n180 VTAIL.n124 289.615
R1350 VTAIL.n118 VTAIL.n62 289.615
R1351 VTAIL.n207 VTAIL.n206 185
R1352 VTAIL.n209 VTAIL.n208 185
R1353 VTAIL.n202 VTAIL.n201 185
R1354 VTAIL.n215 VTAIL.n214 185
R1355 VTAIL.n217 VTAIL.n216 185
R1356 VTAIL.n198 VTAIL.n197 185
R1357 VTAIL.n224 VTAIL.n223 185
R1358 VTAIL.n225 VTAIL.n196 185
R1359 VTAIL.n227 VTAIL.n226 185
R1360 VTAIL.n194 VTAIL.n193 185
R1361 VTAIL.n233 VTAIL.n232 185
R1362 VTAIL.n235 VTAIL.n234 185
R1363 VTAIL.n190 VTAIL.n189 185
R1364 VTAIL.n241 VTAIL.n240 185
R1365 VTAIL.n243 VTAIL.n242 185
R1366 VTAIL.n21 VTAIL.n20 185
R1367 VTAIL.n23 VTAIL.n22 185
R1368 VTAIL.n16 VTAIL.n15 185
R1369 VTAIL.n29 VTAIL.n28 185
R1370 VTAIL.n31 VTAIL.n30 185
R1371 VTAIL.n12 VTAIL.n11 185
R1372 VTAIL.n38 VTAIL.n37 185
R1373 VTAIL.n39 VTAIL.n10 185
R1374 VTAIL.n41 VTAIL.n40 185
R1375 VTAIL.n8 VTAIL.n7 185
R1376 VTAIL.n47 VTAIL.n46 185
R1377 VTAIL.n49 VTAIL.n48 185
R1378 VTAIL.n4 VTAIL.n3 185
R1379 VTAIL.n55 VTAIL.n54 185
R1380 VTAIL.n57 VTAIL.n56 185
R1381 VTAIL.n181 VTAIL.n180 185
R1382 VTAIL.n179 VTAIL.n178 185
R1383 VTAIL.n128 VTAIL.n127 185
R1384 VTAIL.n173 VTAIL.n172 185
R1385 VTAIL.n171 VTAIL.n170 185
R1386 VTAIL.n132 VTAIL.n131 185
R1387 VTAIL.n136 VTAIL.n134 185
R1388 VTAIL.n165 VTAIL.n164 185
R1389 VTAIL.n163 VTAIL.n162 185
R1390 VTAIL.n138 VTAIL.n137 185
R1391 VTAIL.n157 VTAIL.n156 185
R1392 VTAIL.n155 VTAIL.n154 185
R1393 VTAIL.n142 VTAIL.n141 185
R1394 VTAIL.n149 VTAIL.n148 185
R1395 VTAIL.n147 VTAIL.n146 185
R1396 VTAIL.n119 VTAIL.n118 185
R1397 VTAIL.n117 VTAIL.n116 185
R1398 VTAIL.n66 VTAIL.n65 185
R1399 VTAIL.n111 VTAIL.n110 185
R1400 VTAIL.n109 VTAIL.n108 185
R1401 VTAIL.n70 VTAIL.n69 185
R1402 VTAIL.n74 VTAIL.n72 185
R1403 VTAIL.n103 VTAIL.n102 185
R1404 VTAIL.n101 VTAIL.n100 185
R1405 VTAIL.n76 VTAIL.n75 185
R1406 VTAIL.n95 VTAIL.n94 185
R1407 VTAIL.n93 VTAIL.n92 185
R1408 VTAIL.n80 VTAIL.n79 185
R1409 VTAIL.n87 VTAIL.n86 185
R1410 VTAIL.n85 VTAIL.n84 185
R1411 VTAIL.n205 VTAIL.t1 149.524
R1412 VTAIL.n19 VTAIL.t0 149.524
R1413 VTAIL.n145 VTAIL.t3 149.524
R1414 VTAIL.n83 VTAIL.t2 149.524
R1415 VTAIL.n208 VTAIL.n207 104.615
R1416 VTAIL.n208 VTAIL.n201 104.615
R1417 VTAIL.n215 VTAIL.n201 104.615
R1418 VTAIL.n216 VTAIL.n215 104.615
R1419 VTAIL.n216 VTAIL.n197 104.615
R1420 VTAIL.n224 VTAIL.n197 104.615
R1421 VTAIL.n225 VTAIL.n224 104.615
R1422 VTAIL.n226 VTAIL.n225 104.615
R1423 VTAIL.n226 VTAIL.n193 104.615
R1424 VTAIL.n233 VTAIL.n193 104.615
R1425 VTAIL.n234 VTAIL.n233 104.615
R1426 VTAIL.n234 VTAIL.n189 104.615
R1427 VTAIL.n241 VTAIL.n189 104.615
R1428 VTAIL.n242 VTAIL.n241 104.615
R1429 VTAIL.n22 VTAIL.n21 104.615
R1430 VTAIL.n22 VTAIL.n15 104.615
R1431 VTAIL.n29 VTAIL.n15 104.615
R1432 VTAIL.n30 VTAIL.n29 104.615
R1433 VTAIL.n30 VTAIL.n11 104.615
R1434 VTAIL.n38 VTAIL.n11 104.615
R1435 VTAIL.n39 VTAIL.n38 104.615
R1436 VTAIL.n40 VTAIL.n39 104.615
R1437 VTAIL.n40 VTAIL.n7 104.615
R1438 VTAIL.n47 VTAIL.n7 104.615
R1439 VTAIL.n48 VTAIL.n47 104.615
R1440 VTAIL.n48 VTAIL.n3 104.615
R1441 VTAIL.n55 VTAIL.n3 104.615
R1442 VTAIL.n56 VTAIL.n55 104.615
R1443 VTAIL.n180 VTAIL.n179 104.615
R1444 VTAIL.n179 VTAIL.n127 104.615
R1445 VTAIL.n172 VTAIL.n127 104.615
R1446 VTAIL.n172 VTAIL.n171 104.615
R1447 VTAIL.n171 VTAIL.n131 104.615
R1448 VTAIL.n136 VTAIL.n131 104.615
R1449 VTAIL.n164 VTAIL.n136 104.615
R1450 VTAIL.n164 VTAIL.n163 104.615
R1451 VTAIL.n163 VTAIL.n137 104.615
R1452 VTAIL.n156 VTAIL.n137 104.615
R1453 VTAIL.n156 VTAIL.n155 104.615
R1454 VTAIL.n155 VTAIL.n141 104.615
R1455 VTAIL.n148 VTAIL.n141 104.615
R1456 VTAIL.n148 VTAIL.n147 104.615
R1457 VTAIL.n118 VTAIL.n117 104.615
R1458 VTAIL.n117 VTAIL.n65 104.615
R1459 VTAIL.n110 VTAIL.n65 104.615
R1460 VTAIL.n110 VTAIL.n109 104.615
R1461 VTAIL.n109 VTAIL.n69 104.615
R1462 VTAIL.n74 VTAIL.n69 104.615
R1463 VTAIL.n102 VTAIL.n74 104.615
R1464 VTAIL.n102 VTAIL.n101 104.615
R1465 VTAIL.n101 VTAIL.n75 104.615
R1466 VTAIL.n94 VTAIL.n75 104.615
R1467 VTAIL.n94 VTAIL.n93 104.615
R1468 VTAIL.n93 VTAIL.n79 104.615
R1469 VTAIL.n86 VTAIL.n79 104.615
R1470 VTAIL.n86 VTAIL.n85 104.615
R1471 VTAIL.n207 VTAIL.t1 52.3082
R1472 VTAIL.n21 VTAIL.t0 52.3082
R1473 VTAIL.n147 VTAIL.t3 52.3082
R1474 VTAIL.n85 VTAIL.t2 52.3082
R1475 VTAIL.n247 VTAIL.n246 31.0217
R1476 VTAIL.n61 VTAIL.n60 31.0217
R1477 VTAIL.n185 VTAIL.n184 31.0217
R1478 VTAIL.n123 VTAIL.n122 31.0217
R1479 VTAIL.n123 VTAIL.n61 29.4703
R1480 VTAIL.n247 VTAIL.n185 25.8065
R1481 VTAIL.n227 VTAIL.n194 13.1884
R1482 VTAIL.n41 VTAIL.n8 13.1884
R1483 VTAIL.n134 VTAIL.n132 13.1884
R1484 VTAIL.n72 VTAIL.n70 13.1884
R1485 VTAIL.n228 VTAIL.n196 12.8005
R1486 VTAIL.n232 VTAIL.n231 12.8005
R1487 VTAIL.n42 VTAIL.n10 12.8005
R1488 VTAIL.n46 VTAIL.n45 12.8005
R1489 VTAIL.n170 VTAIL.n169 12.8005
R1490 VTAIL.n166 VTAIL.n165 12.8005
R1491 VTAIL.n108 VTAIL.n107 12.8005
R1492 VTAIL.n104 VTAIL.n103 12.8005
R1493 VTAIL.n223 VTAIL.n222 12.0247
R1494 VTAIL.n235 VTAIL.n192 12.0247
R1495 VTAIL.n37 VTAIL.n36 12.0247
R1496 VTAIL.n49 VTAIL.n6 12.0247
R1497 VTAIL.n173 VTAIL.n130 12.0247
R1498 VTAIL.n162 VTAIL.n135 12.0247
R1499 VTAIL.n111 VTAIL.n68 12.0247
R1500 VTAIL.n100 VTAIL.n73 12.0247
R1501 VTAIL.n221 VTAIL.n198 11.249
R1502 VTAIL.n236 VTAIL.n190 11.249
R1503 VTAIL.n35 VTAIL.n12 11.249
R1504 VTAIL.n50 VTAIL.n4 11.249
R1505 VTAIL.n174 VTAIL.n128 11.249
R1506 VTAIL.n161 VTAIL.n138 11.249
R1507 VTAIL.n112 VTAIL.n66 11.249
R1508 VTAIL.n99 VTAIL.n76 11.249
R1509 VTAIL.n218 VTAIL.n217 10.4732
R1510 VTAIL.n240 VTAIL.n239 10.4732
R1511 VTAIL.n32 VTAIL.n31 10.4732
R1512 VTAIL.n54 VTAIL.n53 10.4732
R1513 VTAIL.n178 VTAIL.n177 10.4732
R1514 VTAIL.n158 VTAIL.n157 10.4732
R1515 VTAIL.n116 VTAIL.n115 10.4732
R1516 VTAIL.n96 VTAIL.n95 10.4732
R1517 VTAIL.n206 VTAIL.n205 10.2747
R1518 VTAIL.n20 VTAIL.n19 10.2747
R1519 VTAIL.n146 VTAIL.n145 10.2747
R1520 VTAIL.n84 VTAIL.n83 10.2747
R1521 VTAIL.n214 VTAIL.n200 9.69747
R1522 VTAIL.n243 VTAIL.n188 9.69747
R1523 VTAIL.n28 VTAIL.n14 9.69747
R1524 VTAIL.n57 VTAIL.n2 9.69747
R1525 VTAIL.n181 VTAIL.n126 9.69747
R1526 VTAIL.n154 VTAIL.n140 9.69747
R1527 VTAIL.n119 VTAIL.n64 9.69747
R1528 VTAIL.n92 VTAIL.n78 9.69747
R1529 VTAIL.n246 VTAIL.n245 9.45567
R1530 VTAIL.n60 VTAIL.n59 9.45567
R1531 VTAIL.n184 VTAIL.n183 9.45567
R1532 VTAIL.n122 VTAIL.n121 9.45567
R1533 VTAIL.n245 VTAIL.n244 9.3005
R1534 VTAIL.n188 VTAIL.n187 9.3005
R1535 VTAIL.n239 VTAIL.n238 9.3005
R1536 VTAIL.n237 VTAIL.n236 9.3005
R1537 VTAIL.n192 VTAIL.n191 9.3005
R1538 VTAIL.n231 VTAIL.n230 9.3005
R1539 VTAIL.n204 VTAIL.n203 9.3005
R1540 VTAIL.n211 VTAIL.n210 9.3005
R1541 VTAIL.n213 VTAIL.n212 9.3005
R1542 VTAIL.n200 VTAIL.n199 9.3005
R1543 VTAIL.n219 VTAIL.n218 9.3005
R1544 VTAIL.n221 VTAIL.n220 9.3005
R1545 VTAIL.n222 VTAIL.n195 9.3005
R1546 VTAIL.n229 VTAIL.n228 9.3005
R1547 VTAIL.n59 VTAIL.n58 9.3005
R1548 VTAIL.n2 VTAIL.n1 9.3005
R1549 VTAIL.n53 VTAIL.n52 9.3005
R1550 VTAIL.n51 VTAIL.n50 9.3005
R1551 VTAIL.n6 VTAIL.n5 9.3005
R1552 VTAIL.n45 VTAIL.n44 9.3005
R1553 VTAIL.n18 VTAIL.n17 9.3005
R1554 VTAIL.n25 VTAIL.n24 9.3005
R1555 VTAIL.n27 VTAIL.n26 9.3005
R1556 VTAIL.n14 VTAIL.n13 9.3005
R1557 VTAIL.n33 VTAIL.n32 9.3005
R1558 VTAIL.n35 VTAIL.n34 9.3005
R1559 VTAIL.n36 VTAIL.n9 9.3005
R1560 VTAIL.n43 VTAIL.n42 9.3005
R1561 VTAIL.n144 VTAIL.n143 9.3005
R1562 VTAIL.n151 VTAIL.n150 9.3005
R1563 VTAIL.n153 VTAIL.n152 9.3005
R1564 VTAIL.n140 VTAIL.n139 9.3005
R1565 VTAIL.n159 VTAIL.n158 9.3005
R1566 VTAIL.n161 VTAIL.n160 9.3005
R1567 VTAIL.n135 VTAIL.n133 9.3005
R1568 VTAIL.n167 VTAIL.n166 9.3005
R1569 VTAIL.n183 VTAIL.n182 9.3005
R1570 VTAIL.n126 VTAIL.n125 9.3005
R1571 VTAIL.n177 VTAIL.n176 9.3005
R1572 VTAIL.n175 VTAIL.n174 9.3005
R1573 VTAIL.n130 VTAIL.n129 9.3005
R1574 VTAIL.n169 VTAIL.n168 9.3005
R1575 VTAIL.n82 VTAIL.n81 9.3005
R1576 VTAIL.n89 VTAIL.n88 9.3005
R1577 VTAIL.n91 VTAIL.n90 9.3005
R1578 VTAIL.n78 VTAIL.n77 9.3005
R1579 VTAIL.n97 VTAIL.n96 9.3005
R1580 VTAIL.n99 VTAIL.n98 9.3005
R1581 VTAIL.n73 VTAIL.n71 9.3005
R1582 VTAIL.n105 VTAIL.n104 9.3005
R1583 VTAIL.n121 VTAIL.n120 9.3005
R1584 VTAIL.n64 VTAIL.n63 9.3005
R1585 VTAIL.n115 VTAIL.n114 9.3005
R1586 VTAIL.n113 VTAIL.n112 9.3005
R1587 VTAIL.n68 VTAIL.n67 9.3005
R1588 VTAIL.n107 VTAIL.n106 9.3005
R1589 VTAIL.n213 VTAIL.n202 8.92171
R1590 VTAIL.n244 VTAIL.n186 8.92171
R1591 VTAIL.n27 VTAIL.n16 8.92171
R1592 VTAIL.n58 VTAIL.n0 8.92171
R1593 VTAIL.n182 VTAIL.n124 8.92171
R1594 VTAIL.n153 VTAIL.n142 8.92171
R1595 VTAIL.n120 VTAIL.n62 8.92171
R1596 VTAIL.n91 VTAIL.n80 8.92171
R1597 VTAIL.n210 VTAIL.n209 8.14595
R1598 VTAIL.n24 VTAIL.n23 8.14595
R1599 VTAIL.n150 VTAIL.n149 8.14595
R1600 VTAIL.n88 VTAIL.n87 8.14595
R1601 VTAIL.n206 VTAIL.n204 7.3702
R1602 VTAIL.n20 VTAIL.n18 7.3702
R1603 VTAIL.n146 VTAIL.n144 7.3702
R1604 VTAIL.n84 VTAIL.n82 7.3702
R1605 VTAIL.n209 VTAIL.n204 5.81868
R1606 VTAIL.n23 VTAIL.n18 5.81868
R1607 VTAIL.n149 VTAIL.n144 5.81868
R1608 VTAIL.n87 VTAIL.n82 5.81868
R1609 VTAIL.n210 VTAIL.n202 5.04292
R1610 VTAIL.n246 VTAIL.n186 5.04292
R1611 VTAIL.n24 VTAIL.n16 5.04292
R1612 VTAIL.n60 VTAIL.n0 5.04292
R1613 VTAIL.n184 VTAIL.n124 5.04292
R1614 VTAIL.n150 VTAIL.n142 5.04292
R1615 VTAIL.n122 VTAIL.n62 5.04292
R1616 VTAIL.n88 VTAIL.n80 5.04292
R1617 VTAIL.n214 VTAIL.n213 4.26717
R1618 VTAIL.n244 VTAIL.n243 4.26717
R1619 VTAIL.n28 VTAIL.n27 4.26717
R1620 VTAIL.n58 VTAIL.n57 4.26717
R1621 VTAIL.n182 VTAIL.n181 4.26717
R1622 VTAIL.n154 VTAIL.n153 4.26717
R1623 VTAIL.n120 VTAIL.n119 4.26717
R1624 VTAIL.n92 VTAIL.n91 4.26717
R1625 VTAIL.n217 VTAIL.n200 3.49141
R1626 VTAIL.n240 VTAIL.n188 3.49141
R1627 VTAIL.n31 VTAIL.n14 3.49141
R1628 VTAIL.n54 VTAIL.n2 3.49141
R1629 VTAIL.n178 VTAIL.n126 3.49141
R1630 VTAIL.n157 VTAIL.n140 3.49141
R1631 VTAIL.n116 VTAIL.n64 3.49141
R1632 VTAIL.n95 VTAIL.n78 3.49141
R1633 VTAIL.n205 VTAIL.n203 2.84303
R1634 VTAIL.n19 VTAIL.n17 2.84303
R1635 VTAIL.n145 VTAIL.n143 2.84303
R1636 VTAIL.n83 VTAIL.n81 2.84303
R1637 VTAIL.n218 VTAIL.n198 2.71565
R1638 VTAIL.n239 VTAIL.n190 2.71565
R1639 VTAIL.n32 VTAIL.n12 2.71565
R1640 VTAIL.n53 VTAIL.n4 2.71565
R1641 VTAIL.n177 VTAIL.n128 2.71565
R1642 VTAIL.n158 VTAIL.n138 2.71565
R1643 VTAIL.n115 VTAIL.n66 2.71565
R1644 VTAIL.n96 VTAIL.n76 2.71565
R1645 VTAIL.n185 VTAIL.n123 2.30222
R1646 VTAIL.n223 VTAIL.n221 1.93989
R1647 VTAIL.n236 VTAIL.n235 1.93989
R1648 VTAIL.n37 VTAIL.n35 1.93989
R1649 VTAIL.n50 VTAIL.n49 1.93989
R1650 VTAIL.n174 VTAIL.n173 1.93989
R1651 VTAIL.n162 VTAIL.n161 1.93989
R1652 VTAIL.n112 VTAIL.n111 1.93989
R1653 VTAIL.n100 VTAIL.n99 1.93989
R1654 VTAIL VTAIL.n61 1.44447
R1655 VTAIL.n222 VTAIL.n196 1.16414
R1656 VTAIL.n232 VTAIL.n192 1.16414
R1657 VTAIL.n36 VTAIL.n10 1.16414
R1658 VTAIL.n46 VTAIL.n6 1.16414
R1659 VTAIL.n170 VTAIL.n130 1.16414
R1660 VTAIL.n165 VTAIL.n135 1.16414
R1661 VTAIL.n108 VTAIL.n68 1.16414
R1662 VTAIL.n103 VTAIL.n73 1.16414
R1663 VTAIL VTAIL.n247 0.858259
R1664 VTAIL.n228 VTAIL.n227 0.388379
R1665 VTAIL.n231 VTAIL.n194 0.388379
R1666 VTAIL.n42 VTAIL.n41 0.388379
R1667 VTAIL.n45 VTAIL.n8 0.388379
R1668 VTAIL.n169 VTAIL.n132 0.388379
R1669 VTAIL.n166 VTAIL.n134 0.388379
R1670 VTAIL.n107 VTAIL.n70 0.388379
R1671 VTAIL.n104 VTAIL.n72 0.388379
R1672 VTAIL.n211 VTAIL.n203 0.155672
R1673 VTAIL.n212 VTAIL.n211 0.155672
R1674 VTAIL.n212 VTAIL.n199 0.155672
R1675 VTAIL.n219 VTAIL.n199 0.155672
R1676 VTAIL.n220 VTAIL.n219 0.155672
R1677 VTAIL.n220 VTAIL.n195 0.155672
R1678 VTAIL.n229 VTAIL.n195 0.155672
R1679 VTAIL.n230 VTAIL.n229 0.155672
R1680 VTAIL.n230 VTAIL.n191 0.155672
R1681 VTAIL.n237 VTAIL.n191 0.155672
R1682 VTAIL.n238 VTAIL.n237 0.155672
R1683 VTAIL.n238 VTAIL.n187 0.155672
R1684 VTAIL.n245 VTAIL.n187 0.155672
R1685 VTAIL.n25 VTAIL.n17 0.155672
R1686 VTAIL.n26 VTAIL.n25 0.155672
R1687 VTAIL.n26 VTAIL.n13 0.155672
R1688 VTAIL.n33 VTAIL.n13 0.155672
R1689 VTAIL.n34 VTAIL.n33 0.155672
R1690 VTAIL.n34 VTAIL.n9 0.155672
R1691 VTAIL.n43 VTAIL.n9 0.155672
R1692 VTAIL.n44 VTAIL.n43 0.155672
R1693 VTAIL.n44 VTAIL.n5 0.155672
R1694 VTAIL.n51 VTAIL.n5 0.155672
R1695 VTAIL.n52 VTAIL.n51 0.155672
R1696 VTAIL.n52 VTAIL.n1 0.155672
R1697 VTAIL.n59 VTAIL.n1 0.155672
R1698 VTAIL.n183 VTAIL.n125 0.155672
R1699 VTAIL.n176 VTAIL.n125 0.155672
R1700 VTAIL.n176 VTAIL.n175 0.155672
R1701 VTAIL.n175 VTAIL.n129 0.155672
R1702 VTAIL.n168 VTAIL.n129 0.155672
R1703 VTAIL.n168 VTAIL.n167 0.155672
R1704 VTAIL.n167 VTAIL.n133 0.155672
R1705 VTAIL.n160 VTAIL.n133 0.155672
R1706 VTAIL.n160 VTAIL.n159 0.155672
R1707 VTAIL.n159 VTAIL.n139 0.155672
R1708 VTAIL.n152 VTAIL.n139 0.155672
R1709 VTAIL.n152 VTAIL.n151 0.155672
R1710 VTAIL.n151 VTAIL.n143 0.155672
R1711 VTAIL.n121 VTAIL.n63 0.155672
R1712 VTAIL.n114 VTAIL.n63 0.155672
R1713 VTAIL.n114 VTAIL.n113 0.155672
R1714 VTAIL.n113 VTAIL.n67 0.155672
R1715 VTAIL.n106 VTAIL.n67 0.155672
R1716 VTAIL.n106 VTAIL.n105 0.155672
R1717 VTAIL.n105 VTAIL.n71 0.155672
R1718 VTAIL.n98 VTAIL.n71 0.155672
R1719 VTAIL.n98 VTAIL.n97 0.155672
R1720 VTAIL.n97 VTAIL.n77 0.155672
R1721 VTAIL.n90 VTAIL.n77 0.155672
R1722 VTAIL.n90 VTAIL.n89 0.155672
R1723 VTAIL.n89 VTAIL.n81 0.155672
R1724 VDD2.n117 VDD2.n61 289.615
R1725 VDD2.n56 VDD2.n0 289.615
R1726 VDD2.n118 VDD2.n117 185
R1727 VDD2.n116 VDD2.n115 185
R1728 VDD2.n65 VDD2.n64 185
R1729 VDD2.n110 VDD2.n109 185
R1730 VDD2.n108 VDD2.n107 185
R1731 VDD2.n69 VDD2.n68 185
R1732 VDD2.n73 VDD2.n71 185
R1733 VDD2.n102 VDD2.n101 185
R1734 VDD2.n100 VDD2.n99 185
R1735 VDD2.n75 VDD2.n74 185
R1736 VDD2.n94 VDD2.n93 185
R1737 VDD2.n92 VDD2.n91 185
R1738 VDD2.n79 VDD2.n78 185
R1739 VDD2.n86 VDD2.n85 185
R1740 VDD2.n84 VDD2.n83 185
R1741 VDD2.n21 VDD2.n20 185
R1742 VDD2.n23 VDD2.n22 185
R1743 VDD2.n16 VDD2.n15 185
R1744 VDD2.n29 VDD2.n28 185
R1745 VDD2.n31 VDD2.n30 185
R1746 VDD2.n12 VDD2.n11 185
R1747 VDD2.n38 VDD2.n37 185
R1748 VDD2.n39 VDD2.n10 185
R1749 VDD2.n41 VDD2.n40 185
R1750 VDD2.n8 VDD2.n7 185
R1751 VDD2.n47 VDD2.n46 185
R1752 VDD2.n49 VDD2.n48 185
R1753 VDD2.n4 VDD2.n3 185
R1754 VDD2.n55 VDD2.n54 185
R1755 VDD2.n57 VDD2.n56 185
R1756 VDD2.n82 VDD2.t0 149.524
R1757 VDD2.n19 VDD2.t1 149.524
R1758 VDD2.n117 VDD2.n116 104.615
R1759 VDD2.n116 VDD2.n64 104.615
R1760 VDD2.n109 VDD2.n64 104.615
R1761 VDD2.n109 VDD2.n108 104.615
R1762 VDD2.n108 VDD2.n68 104.615
R1763 VDD2.n73 VDD2.n68 104.615
R1764 VDD2.n101 VDD2.n73 104.615
R1765 VDD2.n101 VDD2.n100 104.615
R1766 VDD2.n100 VDD2.n74 104.615
R1767 VDD2.n93 VDD2.n74 104.615
R1768 VDD2.n93 VDD2.n92 104.615
R1769 VDD2.n92 VDD2.n78 104.615
R1770 VDD2.n85 VDD2.n78 104.615
R1771 VDD2.n85 VDD2.n84 104.615
R1772 VDD2.n22 VDD2.n21 104.615
R1773 VDD2.n22 VDD2.n15 104.615
R1774 VDD2.n29 VDD2.n15 104.615
R1775 VDD2.n30 VDD2.n29 104.615
R1776 VDD2.n30 VDD2.n11 104.615
R1777 VDD2.n38 VDD2.n11 104.615
R1778 VDD2.n39 VDD2.n38 104.615
R1779 VDD2.n40 VDD2.n39 104.615
R1780 VDD2.n40 VDD2.n7 104.615
R1781 VDD2.n47 VDD2.n7 104.615
R1782 VDD2.n48 VDD2.n47 104.615
R1783 VDD2.n48 VDD2.n3 104.615
R1784 VDD2.n55 VDD2.n3 104.615
R1785 VDD2.n56 VDD2.n55 104.615
R1786 VDD2.n122 VDD2.n60 88.4634
R1787 VDD2.n84 VDD2.t0 52.3082
R1788 VDD2.n21 VDD2.t1 52.3082
R1789 VDD2.n122 VDD2.n121 47.7005
R1790 VDD2.n71 VDD2.n69 13.1884
R1791 VDD2.n41 VDD2.n8 13.1884
R1792 VDD2.n107 VDD2.n106 12.8005
R1793 VDD2.n103 VDD2.n102 12.8005
R1794 VDD2.n42 VDD2.n10 12.8005
R1795 VDD2.n46 VDD2.n45 12.8005
R1796 VDD2.n110 VDD2.n67 12.0247
R1797 VDD2.n99 VDD2.n72 12.0247
R1798 VDD2.n37 VDD2.n36 12.0247
R1799 VDD2.n49 VDD2.n6 12.0247
R1800 VDD2.n111 VDD2.n65 11.249
R1801 VDD2.n98 VDD2.n75 11.249
R1802 VDD2.n35 VDD2.n12 11.249
R1803 VDD2.n50 VDD2.n4 11.249
R1804 VDD2.n115 VDD2.n114 10.4732
R1805 VDD2.n95 VDD2.n94 10.4732
R1806 VDD2.n32 VDD2.n31 10.4732
R1807 VDD2.n54 VDD2.n53 10.4732
R1808 VDD2.n83 VDD2.n82 10.2747
R1809 VDD2.n20 VDD2.n19 10.2747
R1810 VDD2.n118 VDD2.n63 9.69747
R1811 VDD2.n91 VDD2.n77 9.69747
R1812 VDD2.n28 VDD2.n14 9.69747
R1813 VDD2.n57 VDD2.n2 9.69747
R1814 VDD2.n121 VDD2.n120 9.45567
R1815 VDD2.n60 VDD2.n59 9.45567
R1816 VDD2.n81 VDD2.n80 9.3005
R1817 VDD2.n88 VDD2.n87 9.3005
R1818 VDD2.n90 VDD2.n89 9.3005
R1819 VDD2.n77 VDD2.n76 9.3005
R1820 VDD2.n96 VDD2.n95 9.3005
R1821 VDD2.n98 VDD2.n97 9.3005
R1822 VDD2.n72 VDD2.n70 9.3005
R1823 VDD2.n104 VDD2.n103 9.3005
R1824 VDD2.n120 VDD2.n119 9.3005
R1825 VDD2.n63 VDD2.n62 9.3005
R1826 VDD2.n114 VDD2.n113 9.3005
R1827 VDD2.n112 VDD2.n111 9.3005
R1828 VDD2.n67 VDD2.n66 9.3005
R1829 VDD2.n106 VDD2.n105 9.3005
R1830 VDD2.n59 VDD2.n58 9.3005
R1831 VDD2.n2 VDD2.n1 9.3005
R1832 VDD2.n53 VDD2.n52 9.3005
R1833 VDD2.n51 VDD2.n50 9.3005
R1834 VDD2.n6 VDD2.n5 9.3005
R1835 VDD2.n45 VDD2.n44 9.3005
R1836 VDD2.n18 VDD2.n17 9.3005
R1837 VDD2.n25 VDD2.n24 9.3005
R1838 VDD2.n27 VDD2.n26 9.3005
R1839 VDD2.n14 VDD2.n13 9.3005
R1840 VDD2.n33 VDD2.n32 9.3005
R1841 VDD2.n35 VDD2.n34 9.3005
R1842 VDD2.n36 VDD2.n9 9.3005
R1843 VDD2.n43 VDD2.n42 9.3005
R1844 VDD2.n119 VDD2.n61 8.92171
R1845 VDD2.n90 VDD2.n79 8.92171
R1846 VDD2.n27 VDD2.n16 8.92171
R1847 VDD2.n58 VDD2.n0 8.92171
R1848 VDD2.n87 VDD2.n86 8.14595
R1849 VDD2.n24 VDD2.n23 8.14595
R1850 VDD2.n83 VDD2.n81 7.3702
R1851 VDD2.n20 VDD2.n18 7.3702
R1852 VDD2.n86 VDD2.n81 5.81868
R1853 VDD2.n23 VDD2.n18 5.81868
R1854 VDD2.n121 VDD2.n61 5.04292
R1855 VDD2.n87 VDD2.n79 5.04292
R1856 VDD2.n24 VDD2.n16 5.04292
R1857 VDD2.n60 VDD2.n0 5.04292
R1858 VDD2.n119 VDD2.n118 4.26717
R1859 VDD2.n91 VDD2.n90 4.26717
R1860 VDD2.n28 VDD2.n27 4.26717
R1861 VDD2.n58 VDD2.n57 4.26717
R1862 VDD2.n115 VDD2.n63 3.49141
R1863 VDD2.n94 VDD2.n77 3.49141
R1864 VDD2.n31 VDD2.n14 3.49141
R1865 VDD2.n54 VDD2.n2 3.49141
R1866 VDD2.n82 VDD2.n80 2.84303
R1867 VDD2.n19 VDD2.n17 2.84303
R1868 VDD2.n114 VDD2.n65 2.71565
R1869 VDD2.n95 VDD2.n75 2.71565
R1870 VDD2.n32 VDD2.n12 2.71565
R1871 VDD2.n53 VDD2.n4 2.71565
R1872 VDD2.n111 VDD2.n110 1.93989
R1873 VDD2.n99 VDD2.n98 1.93989
R1874 VDD2.n37 VDD2.n35 1.93989
R1875 VDD2.n50 VDD2.n49 1.93989
R1876 VDD2.n107 VDD2.n67 1.16414
R1877 VDD2.n102 VDD2.n72 1.16414
R1878 VDD2.n36 VDD2.n10 1.16414
R1879 VDD2.n46 VDD2.n6 1.16414
R1880 VDD2 VDD2.n122 0.974638
R1881 VDD2.n106 VDD2.n69 0.388379
R1882 VDD2.n103 VDD2.n71 0.388379
R1883 VDD2.n42 VDD2.n41 0.388379
R1884 VDD2.n45 VDD2.n8 0.388379
R1885 VDD2.n120 VDD2.n62 0.155672
R1886 VDD2.n113 VDD2.n62 0.155672
R1887 VDD2.n113 VDD2.n112 0.155672
R1888 VDD2.n112 VDD2.n66 0.155672
R1889 VDD2.n105 VDD2.n66 0.155672
R1890 VDD2.n105 VDD2.n104 0.155672
R1891 VDD2.n104 VDD2.n70 0.155672
R1892 VDD2.n97 VDD2.n70 0.155672
R1893 VDD2.n97 VDD2.n96 0.155672
R1894 VDD2.n96 VDD2.n76 0.155672
R1895 VDD2.n89 VDD2.n76 0.155672
R1896 VDD2.n89 VDD2.n88 0.155672
R1897 VDD2.n88 VDD2.n80 0.155672
R1898 VDD2.n25 VDD2.n17 0.155672
R1899 VDD2.n26 VDD2.n25 0.155672
R1900 VDD2.n26 VDD2.n13 0.155672
R1901 VDD2.n33 VDD2.n13 0.155672
R1902 VDD2.n34 VDD2.n33 0.155672
R1903 VDD2.n34 VDD2.n9 0.155672
R1904 VDD2.n43 VDD2.n9 0.155672
R1905 VDD2.n44 VDD2.n43 0.155672
R1906 VDD2.n44 VDD2.n5 0.155672
R1907 VDD2.n51 VDD2.n5 0.155672
R1908 VDD2.n52 VDD2.n51 0.155672
R1909 VDD2.n52 VDD2.n1 0.155672
R1910 VDD2.n59 VDD2.n1 0.155672
R1911 VP.n0 VP.t0 152.466
R1912 VP.n0 VP.t1 104.809
R1913 VP VP.n0 0.62124
R1914 VDD1.n56 VDD1.n0 289.615
R1915 VDD1.n117 VDD1.n61 289.615
R1916 VDD1.n57 VDD1.n56 185
R1917 VDD1.n55 VDD1.n54 185
R1918 VDD1.n4 VDD1.n3 185
R1919 VDD1.n49 VDD1.n48 185
R1920 VDD1.n47 VDD1.n46 185
R1921 VDD1.n8 VDD1.n7 185
R1922 VDD1.n12 VDD1.n10 185
R1923 VDD1.n41 VDD1.n40 185
R1924 VDD1.n39 VDD1.n38 185
R1925 VDD1.n14 VDD1.n13 185
R1926 VDD1.n33 VDD1.n32 185
R1927 VDD1.n31 VDD1.n30 185
R1928 VDD1.n18 VDD1.n17 185
R1929 VDD1.n25 VDD1.n24 185
R1930 VDD1.n23 VDD1.n22 185
R1931 VDD1.n82 VDD1.n81 185
R1932 VDD1.n84 VDD1.n83 185
R1933 VDD1.n77 VDD1.n76 185
R1934 VDD1.n90 VDD1.n89 185
R1935 VDD1.n92 VDD1.n91 185
R1936 VDD1.n73 VDD1.n72 185
R1937 VDD1.n99 VDD1.n98 185
R1938 VDD1.n100 VDD1.n71 185
R1939 VDD1.n102 VDD1.n101 185
R1940 VDD1.n69 VDD1.n68 185
R1941 VDD1.n108 VDD1.n107 185
R1942 VDD1.n110 VDD1.n109 185
R1943 VDD1.n65 VDD1.n64 185
R1944 VDD1.n116 VDD1.n115 185
R1945 VDD1.n118 VDD1.n117 185
R1946 VDD1.n21 VDD1.t1 149.524
R1947 VDD1.n80 VDD1.t0 149.524
R1948 VDD1.n56 VDD1.n55 104.615
R1949 VDD1.n55 VDD1.n3 104.615
R1950 VDD1.n48 VDD1.n3 104.615
R1951 VDD1.n48 VDD1.n47 104.615
R1952 VDD1.n47 VDD1.n7 104.615
R1953 VDD1.n12 VDD1.n7 104.615
R1954 VDD1.n40 VDD1.n12 104.615
R1955 VDD1.n40 VDD1.n39 104.615
R1956 VDD1.n39 VDD1.n13 104.615
R1957 VDD1.n32 VDD1.n13 104.615
R1958 VDD1.n32 VDD1.n31 104.615
R1959 VDD1.n31 VDD1.n17 104.615
R1960 VDD1.n24 VDD1.n17 104.615
R1961 VDD1.n24 VDD1.n23 104.615
R1962 VDD1.n83 VDD1.n82 104.615
R1963 VDD1.n83 VDD1.n76 104.615
R1964 VDD1.n90 VDD1.n76 104.615
R1965 VDD1.n91 VDD1.n90 104.615
R1966 VDD1.n91 VDD1.n72 104.615
R1967 VDD1.n99 VDD1.n72 104.615
R1968 VDD1.n100 VDD1.n99 104.615
R1969 VDD1.n101 VDD1.n100 104.615
R1970 VDD1.n101 VDD1.n68 104.615
R1971 VDD1.n108 VDD1.n68 104.615
R1972 VDD1.n109 VDD1.n108 104.615
R1973 VDD1.n109 VDD1.n64 104.615
R1974 VDD1.n116 VDD1.n64 104.615
R1975 VDD1.n117 VDD1.n116 104.615
R1976 VDD1 VDD1.n121 89.9042
R1977 VDD1.n23 VDD1.t1 52.3082
R1978 VDD1.n82 VDD1.t0 52.3082
R1979 VDD1 VDD1.n60 48.6746
R1980 VDD1.n10 VDD1.n8 13.1884
R1981 VDD1.n102 VDD1.n69 13.1884
R1982 VDD1.n46 VDD1.n45 12.8005
R1983 VDD1.n42 VDD1.n41 12.8005
R1984 VDD1.n103 VDD1.n71 12.8005
R1985 VDD1.n107 VDD1.n106 12.8005
R1986 VDD1.n49 VDD1.n6 12.0247
R1987 VDD1.n38 VDD1.n11 12.0247
R1988 VDD1.n98 VDD1.n97 12.0247
R1989 VDD1.n110 VDD1.n67 12.0247
R1990 VDD1.n50 VDD1.n4 11.249
R1991 VDD1.n37 VDD1.n14 11.249
R1992 VDD1.n96 VDD1.n73 11.249
R1993 VDD1.n111 VDD1.n65 11.249
R1994 VDD1.n54 VDD1.n53 10.4732
R1995 VDD1.n34 VDD1.n33 10.4732
R1996 VDD1.n93 VDD1.n92 10.4732
R1997 VDD1.n115 VDD1.n114 10.4732
R1998 VDD1.n22 VDD1.n21 10.2747
R1999 VDD1.n81 VDD1.n80 10.2747
R2000 VDD1.n57 VDD1.n2 9.69747
R2001 VDD1.n30 VDD1.n16 9.69747
R2002 VDD1.n89 VDD1.n75 9.69747
R2003 VDD1.n118 VDD1.n63 9.69747
R2004 VDD1.n60 VDD1.n59 9.45567
R2005 VDD1.n121 VDD1.n120 9.45567
R2006 VDD1.n20 VDD1.n19 9.3005
R2007 VDD1.n27 VDD1.n26 9.3005
R2008 VDD1.n29 VDD1.n28 9.3005
R2009 VDD1.n16 VDD1.n15 9.3005
R2010 VDD1.n35 VDD1.n34 9.3005
R2011 VDD1.n37 VDD1.n36 9.3005
R2012 VDD1.n11 VDD1.n9 9.3005
R2013 VDD1.n43 VDD1.n42 9.3005
R2014 VDD1.n59 VDD1.n58 9.3005
R2015 VDD1.n2 VDD1.n1 9.3005
R2016 VDD1.n53 VDD1.n52 9.3005
R2017 VDD1.n51 VDD1.n50 9.3005
R2018 VDD1.n6 VDD1.n5 9.3005
R2019 VDD1.n45 VDD1.n44 9.3005
R2020 VDD1.n120 VDD1.n119 9.3005
R2021 VDD1.n63 VDD1.n62 9.3005
R2022 VDD1.n114 VDD1.n113 9.3005
R2023 VDD1.n112 VDD1.n111 9.3005
R2024 VDD1.n67 VDD1.n66 9.3005
R2025 VDD1.n106 VDD1.n105 9.3005
R2026 VDD1.n79 VDD1.n78 9.3005
R2027 VDD1.n86 VDD1.n85 9.3005
R2028 VDD1.n88 VDD1.n87 9.3005
R2029 VDD1.n75 VDD1.n74 9.3005
R2030 VDD1.n94 VDD1.n93 9.3005
R2031 VDD1.n96 VDD1.n95 9.3005
R2032 VDD1.n97 VDD1.n70 9.3005
R2033 VDD1.n104 VDD1.n103 9.3005
R2034 VDD1.n58 VDD1.n0 8.92171
R2035 VDD1.n29 VDD1.n18 8.92171
R2036 VDD1.n88 VDD1.n77 8.92171
R2037 VDD1.n119 VDD1.n61 8.92171
R2038 VDD1.n26 VDD1.n25 8.14595
R2039 VDD1.n85 VDD1.n84 8.14595
R2040 VDD1.n22 VDD1.n20 7.3702
R2041 VDD1.n81 VDD1.n79 7.3702
R2042 VDD1.n25 VDD1.n20 5.81868
R2043 VDD1.n84 VDD1.n79 5.81868
R2044 VDD1.n60 VDD1.n0 5.04292
R2045 VDD1.n26 VDD1.n18 5.04292
R2046 VDD1.n85 VDD1.n77 5.04292
R2047 VDD1.n121 VDD1.n61 5.04292
R2048 VDD1.n58 VDD1.n57 4.26717
R2049 VDD1.n30 VDD1.n29 4.26717
R2050 VDD1.n89 VDD1.n88 4.26717
R2051 VDD1.n119 VDD1.n118 4.26717
R2052 VDD1.n54 VDD1.n2 3.49141
R2053 VDD1.n33 VDD1.n16 3.49141
R2054 VDD1.n92 VDD1.n75 3.49141
R2055 VDD1.n115 VDD1.n63 3.49141
R2056 VDD1.n21 VDD1.n19 2.84303
R2057 VDD1.n80 VDD1.n78 2.84303
R2058 VDD1.n53 VDD1.n4 2.71565
R2059 VDD1.n34 VDD1.n14 2.71565
R2060 VDD1.n93 VDD1.n73 2.71565
R2061 VDD1.n114 VDD1.n65 2.71565
R2062 VDD1.n50 VDD1.n49 1.93989
R2063 VDD1.n38 VDD1.n37 1.93989
R2064 VDD1.n98 VDD1.n96 1.93989
R2065 VDD1.n111 VDD1.n110 1.93989
R2066 VDD1.n46 VDD1.n6 1.16414
R2067 VDD1.n41 VDD1.n11 1.16414
R2068 VDD1.n97 VDD1.n71 1.16414
R2069 VDD1.n107 VDD1.n67 1.16414
R2070 VDD1.n45 VDD1.n8 0.388379
R2071 VDD1.n42 VDD1.n10 0.388379
R2072 VDD1.n103 VDD1.n102 0.388379
R2073 VDD1.n106 VDD1.n69 0.388379
R2074 VDD1.n59 VDD1.n1 0.155672
R2075 VDD1.n52 VDD1.n1 0.155672
R2076 VDD1.n52 VDD1.n51 0.155672
R2077 VDD1.n51 VDD1.n5 0.155672
R2078 VDD1.n44 VDD1.n5 0.155672
R2079 VDD1.n44 VDD1.n43 0.155672
R2080 VDD1.n43 VDD1.n9 0.155672
R2081 VDD1.n36 VDD1.n9 0.155672
R2082 VDD1.n36 VDD1.n35 0.155672
R2083 VDD1.n35 VDD1.n15 0.155672
R2084 VDD1.n28 VDD1.n15 0.155672
R2085 VDD1.n28 VDD1.n27 0.155672
R2086 VDD1.n27 VDD1.n19 0.155672
R2087 VDD1.n86 VDD1.n78 0.155672
R2088 VDD1.n87 VDD1.n86 0.155672
R2089 VDD1.n87 VDD1.n74 0.155672
R2090 VDD1.n94 VDD1.n74 0.155672
R2091 VDD1.n95 VDD1.n94 0.155672
R2092 VDD1.n95 VDD1.n70 0.155672
R2093 VDD1.n104 VDD1.n70 0.155672
R2094 VDD1.n105 VDD1.n104 0.155672
R2095 VDD1.n105 VDD1.n66 0.155672
R2096 VDD1.n112 VDD1.n66 0.155672
R2097 VDD1.n113 VDD1.n112 0.155672
R2098 VDD1.n113 VDD1.n62 0.155672
R2099 VDD1.n120 VDD1.n62 0.155672
C0 VN VTAIL 2.56252f
C1 VDD1 VDD2 0.823151f
C2 VDD1 VP 3.02106f
C3 VP VDD2 0.388213f
C4 VN VDD1 0.149063f
C5 VTAIL VDD1 5.18029f
C6 VN VDD2 2.78325f
C7 VN VP 5.94954f
C8 VTAIL VDD2 5.24088f
C9 VTAIL VP 2.57737f
C10 VDD2 B 4.790049f
C11 VDD1 B 7.748539f
C12 VTAIL B 7.708817f
C13 VN B 11.91788f
C14 VP B 7.995059f
C15 VDD1.n0 B 0.027878f
C16 VDD1.n1 B 0.020834f
C17 VDD1.n2 B 0.011195f
C18 VDD1.n3 B 0.026461f
C19 VDD1.n4 B 0.011854f
C20 VDD1.n5 B 0.020834f
C21 VDD1.n6 B 0.011195f
C22 VDD1.n7 B 0.026461f
C23 VDD1.n8 B 0.011524f
C24 VDD1.n9 B 0.020834f
C25 VDD1.n10 B 0.011524f
C26 VDD1.n11 B 0.011195f
C27 VDD1.n12 B 0.026461f
C28 VDD1.n13 B 0.026461f
C29 VDD1.n14 B 0.011854f
C30 VDD1.n15 B 0.020834f
C31 VDD1.n16 B 0.011195f
C32 VDD1.n17 B 0.026461f
C33 VDD1.n18 B 0.011854f
C34 VDD1.n19 B 0.989873f
C35 VDD1.n20 B 0.011195f
C36 VDD1.t1 B 0.044618f
C37 VDD1.n21 B 0.144931f
C38 VDD1.n22 B 0.018706f
C39 VDD1.n23 B 0.019846f
C40 VDD1.n24 B 0.026461f
C41 VDD1.n25 B 0.011854f
C42 VDD1.n26 B 0.011195f
C43 VDD1.n27 B 0.020834f
C44 VDD1.n28 B 0.020834f
C45 VDD1.n29 B 0.011195f
C46 VDD1.n30 B 0.011854f
C47 VDD1.n31 B 0.026461f
C48 VDD1.n32 B 0.026461f
C49 VDD1.n33 B 0.011854f
C50 VDD1.n34 B 0.011195f
C51 VDD1.n35 B 0.020834f
C52 VDD1.n36 B 0.020834f
C53 VDD1.n37 B 0.011195f
C54 VDD1.n38 B 0.011854f
C55 VDD1.n39 B 0.026461f
C56 VDD1.n40 B 0.026461f
C57 VDD1.n41 B 0.011854f
C58 VDD1.n42 B 0.011195f
C59 VDD1.n43 B 0.020834f
C60 VDD1.n44 B 0.020834f
C61 VDD1.n45 B 0.011195f
C62 VDD1.n46 B 0.011854f
C63 VDD1.n47 B 0.026461f
C64 VDD1.n48 B 0.026461f
C65 VDD1.n49 B 0.011854f
C66 VDD1.n50 B 0.011195f
C67 VDD1.n51 B 0.020834f
C68 VDD1.n52 B 0.020834f
C69 VDD1.n53 B 0.011195f
C70 VDD1.n54 B 0.011854f
C71 VDD1.n55 B 0.026461f
C72 VDD1.n56 B 0.054799f
C73 VDD1.n57 B 0.011854f
C74 VDD1.n58 B 0.011195f
C75 VDD1.n59 B 0.046449f
C76 VDD1.n60 B 0.046845f
C77 VDD1.n61 B 0.027878f
C78 VDD1.n62 B 0.020834f
C79 VDD1.n63 B 0.011195f
C80 VDD1.n64 B 0.026461f
C81 VDD1.n65 B 0.011854f
C82 VDD1.n66 B 0.020834f
C83 VDD1.n67 B 0.011195f
C84 VDD1.n68 B 0.026461f
C85 VDD1.n69 B 0.011524f
C86 VDD1.n70 B 0.020834f
C87 VDD1.n71 B 0.011854f
C88 VDD1.n72 B 0.026461f
C89 VDD1.n73 B 0.011854f
C90 VDD1.n74 B 0.020834f
C91 VDD1.n75 B 0.011195f
C92 VDD1.n76 B 0.026461f
C93 VDD1.n77 B 0.011854f
C94 VDD1.n78 B 0.989873f
C95 VDD1.n79 B 0.011195f
C96 VDD1.t0 B 0.044618f
C97 VDD1.n80 B 0.144931f
C98 VDD1.n81 B 0.018706f
C99 VDD1.n82 B 0.019846f
C100 VDD1.n83 B 0.026461f
C101 VDD1.n84 B 0.011854f
C102 VDD1.n85 B 0.011195f
C103 VDD1.n86 B 0.020834f
C104 VDD1.n87 B 0.020834f
C105 VDD1.n88 B 0.011195f
C106 VDD1.n89 B 0.011854f
C107 VDD1.n90 B 0.026461f
C108 VDD1.n91 B 0.026461f
C109 VDD1.n92 B 0.011854f
C110 VDD1.n93 B 0.011195f
C111 VDD1.n94 B 0.020834f
C112 VDD1.n95 B 0.020834f
C113 VDD1.n96 B 0.011195f
C114 VDD1.n97 B 0.011195f
C115 VDD1.n98 B 0.011854f
C116 VDD1.n99 B 0.026461f
C117 VDD1.n100 B 0.026461f
C118 VDD1.n101 B 0.026461f
C119 VDD1.n102 B 0.011524f
C120 VDD1.n103 B 0.011195f
C121 VDD1.n104 B 0.020834f
C122 VDD1.n105 B 0.020834f
C123 VDD1.n106 B 0.011195f
C124 VDD1.n107 B 0.011854f
C125 VDD1.n108 B 0.026461f
C126 VDD1.n109 B 0.026461f
C127 VDD1.n110 B 0.011854f
C128 VDD1.n111 B 0.011195f
C129 VDD1.n112 B 0.020834f
C130 VDD1.n113 B 0.020834f
C131 VDD1.n114 B 0.011195f
C132 VDD1.n115 B 0.011854f
C133 VDD1.n116 B 0.026461f
C134 VDD1.n117 B 0.054799f
C135 VDD1.n118 B 0.011854f
C136 VDD1.n119 B 0.011195f
C137 VDD1.n120 B 0.046449f
C138 VDD1.n121 B 0.722656f
C139 VP.t0 B 4.14117f
C140 VP.t1 B 3.41389f
C141 VP.n0 B 3.83594f
C142 VDD2.n0 B 0.027456f
C143 VDD2.n1 B 0.020518f
C144 VDD2.n2 B 0.011026f
C145 VDD2.n3 B 0.026061f
C146 VDD2.n4 B 0.011674f
C147 VDD2.n5 B 0.020518f
C148 VDD2.n6 B 0.011026f
C149 VDD2.n7 B 0.026061f
C150 VDD2.n8 B 0.01135f
C151 VDD2.n9 B 0.020518f
C152 VDD2.n10 B 0.011674f
C153 VDD2.n11 B 0.026061f
C154 VDD2.n12 B 0.011674f
C155 VDD2.n13 B 0.020518f
C156 VDD2.n14 B 0.011026f
C157 VDD2.n15 B 0.026061f
C158 VDD2.n16 B 0.011674f
C159 VDD2.n17 B 0.974878f
C160 VDD2.n18 B 0.011026f
C161 VDD2.t1 B 0.043942f
C162 VDD2.n19 B 0.142736f
C163 VDD2.n20 B 0.018423f
C164 VDD2.n21 B 0.019545f
C165 VDD2.n22 B 0.026061f
C166 VDD2.n23 B 0.011674f
C167 VDD2.n24 B 0.011026f
C168 VDD2.n25 B 0.020518f
C169 VDD2.n26 B 0.020518f
C170 VDD2.n27 B 0.011026f
C171 VDD2.n28 B 0.011674f
C172 VDD2.n29 B 0.026061f
C173 VDD2.n30 B 0.026061f
C174 VDD2.n31 B 0.011674f
C175 VDD2.n32 B 0.011026f
C176 VDD2.n33 B 0.020518f
C177 VDD2.n34 B 0.020518f
C178 VDD2.n35 B 0.011026f
C179 VDD2.n36 B 0.011026f
C180 VDD2.n37 B 0.011674f
C181 VDD2.n38 B 0.026061f
C182 VDD2.n39 B 0.026061f
C183 VDD2.n40 B 0.026061f
C184 VDD2.n41 B 0.01135f
C185 VDD2.n42 B 0.011026f
C186 VDD2.n43 B 0.020518f
C187 VDD2.n44 B 0.020518f
C188 VDD2.n45 B 0.011026f
C189 VDD2.n46 B 0.011674f
C190 VDD2.n47 B 0.026061f
C191 VDD2.n48 B 0.026061f
C192 VDD2.n49 B 0.011674f
C193 VDD2.n50 B 0.011026f
C194 VDD2.n51 B 0.020518f
C195 VDD2.n52 B 0.020518f
C196 VDD2.n53 B 0.011026f
C197 VDD2.n54 B 0.011674f
C198 VDD2.n55 B 0.026061f
C199 VDD2.n56 B 0.053969f
C200 VDD2.n57 B 0.011674f
C201 VDD2.n58 B 0.011026f
C202 VDD2.n59 B 0.045745f
C203 VDD2.n60 B 0.661573f
C204 VDD2.n61 B 0.027456f
C205 VDD2.n62 B 0.020518f
C206 VDD2.n63 B 0.011026f
C207 VDD2.n64 B 0.026061f
C208 VDD2.n65 B 0.011674f
C209 VDD2.n66 B 0.020518f
C210 VDD2.n67 B 0.011026f
C211 VDD2.n68 B 0.026061f
C212 VDD2.n69 B 0.01135f
C213 VDD2.n70 B 0.020518f
C214 VDD2.n71 B 0.01135f
C215 VDD2.n72 B 0.011026f
C216 VDD2.n73 B 0.026061f
C217 VDD2.n74 B 0.026061f
C218 VDD2.n75 B 0.011674f
C219 VDD2.n76 B 0.020518f
C220 VDD2.n77 B 0.011026f
C221 VDD2.n78 B 0.026061f
C222 VDD2.n79 B 0.011674f
C223 VDD2.n80 B 0.974878f
C224 VDD2.n81 B 0.011026f
C225 VDD2.t0 B 0.043942f
C226 VDD2.n82 B 0.142736f
C227 VDD2.n83 B 0.018423f
C228 VDD2.n84 B 0.019545f
C229 VDD2.n85 B 0.026061f
C230 VDD2.n86 B 0.011674f
C231 VDD2.n87 B 0.011026f
C232 VDD2.n88 B 0.020518f
C233 VDD2.n89 B 0.020518f
C234 VDD2.n90 B 0.011026f
C235 VDD2.n91 B 0.011674f
C236 VDD2.n92 B 0.026061f
C237 VDD2.n93 B 0.026061f
C238 VDD2.n94 B 0.011674f
C239 VDD2.n95 B 0.011026f
C240 VDD2.n96 B 0.020518f
C241 VDD2.n97 B 0.020518f
C242 VDD2.n98 B 0.011026f
C243 VDD2.n99 B 0.011674f
C244 VDD2.n100 B 0.026061f
C245 VDD2.n101 B 0.026061f
C246 VDD2.n102 B 0.011674f
C247 VDD2.n103 B 0.011026f
C248 VDD2.n104 B 0.020518f
C249 VDD2.n105 B 0.020518f
C250 VDD2.n106 B 0.011026f
C251 VDD2.n107 B 0.011674f
C252 VDD2.n108 B 0.026061f
C253 VDD2.n109 B 0.026061f
C254 VDD2.n110 B 0.011674f
C255 VDD2.n111 B 0.011026f
C256 VDD2.n112 B 0.020518f
C257 VDD2.n113 B 0.020518f
C258 VDD2.n114 B 0.011026f
C259 VDD2.n115 B 0.011674f
C260 VDD2.n116 B 0.026061f
C261 VDD2.n117 B 0.053969f
C262 VDD2.n118 B 0.011674f
C263 VDD2.n119 B 0.011026f
C264 VDD2.n120 B 0.045745f
C265 VDD2.n121 B 0.044075f
C266 VDD2.n122 B 2.65056f
C267 VTAIL.n0 B 0.028816f
C268 VTAIL.n1 B 0.021535f
C269 VTAIL.n2 B 0.011572f
C270 VTAIL.n3 B 0.027352f
C271 VTAIL.n4 B 0.012253f
C272 VTAIL.n5 B 0.021535f
C273 VTAIL.n6 B 0.011572f
C274 VTAIL.n7 B 0.027352f
C275 VTAIL.n8 B 0.011912f
C276 VTAIL.n9 B 0.021535f
C277 VTAIL.n10 B 0.012253f
C278 VTAIL.n11 B 0.027352f
C279 VTAIL.n12 B 0.012253f
C280 VTAIL.n13 B 0.021535f
C281 VTAIL.n14 B 0.011572f
C282 VTAIL.n15 B 0.027352f
C283 VTAIL.n16 B 0.012253f
C284 VTAIL.n17 B 1.02318f
C285 VTAIL.n18 B 0.011572f
C286 VTAIL.t0 B 0.046119f
C287 VTAIL.n19 B 0.149808f
C288 VTAIL.n20 B 0.019336f
C289 VTAIL.n21 B 0.020514f
C290 VTAIL.n22 B 0.027352f
C291 VTAIL.n23 B 0.012253f
C292 VTAIL.n24 B 0.011572f
C293 VTAIL.n25 B 0.021535f
C294 VTAIL.n26 B 0.021535f
C295 VTAIL.n27 B 0.011572f
C296 VTAIL.n28 B 0.012253f
C297 VTAIL.n29 B 0.027352f
C298 VTAIL.n30 B 0.027352f
C299 VTAIL.n31 B 0.012253f
C300 VTAIL.n32 B 0.011572f
C301 VTAIL.n33 B 0.021535f
C302 VTAIL.n34 B 0.021535f
C303 VTAIL.n35 B 0.011572f
C304 VTAIL.n36 B 0.011572f
C305 VTAIL.n37 B 0.012253f
C306 VTAIL.n38 B 0.027352f
C307 VTAIL.n39 B 0.027352f
C308 VTAIL.n40 B 0.027352f
C309 VTAIL.n41 B 0.011912f
C310 VTAIL.n42 B 0.011572f
C311 VTAIL.n43 B 0.021535f
C312 VTAIL.n44 B 0.021535f
C313 VTAIL.n45 B 0.011572f
C314 VTAIL.n46 B 0.012253f
C315 VTAIL.n47 B 0.027352f
C316 VTAIL.n48 B 0.027352f
C317 VTAIL.n49 B 0.012253f
C318 VTAIL.n50 B 0.011572f
C319 VTAIL.n51 B 0.021535f
C320 VTAIL.n52 B 0.021535f
C321 VTAIL.n53 B 0.011572f
C322 VTAIL.n54 B 0.012253f
C323 VTAIL.n55 B 0.027352f
C324 VTAIL.n56 B 0.056643f
C325 VTAIL.n57 B 0.012253f
C326 VTAIL.n58 B 0.011572f
C327 VTAIL.n59 B 0.048012f
C328 VTAIL.n60 B 0.031375f
C329 VTAIL.n61 B 1.59694f
C330 VTAIL.n62 B 0.028816f
C331 VTAIL.n63 B 0.021535f
C332 VTAIL.n64 B 0.011572f
C333 VTAIL.n65 B 0.027352f
C334 VTAIL.n66 B 0.012253f
C335 VTAIL.n67 B 0.021535f
C336 VTAIL.n68 B 0.011572f
C337 VTAIL.n69 B 0.027352f
C338 VTAIL.n70 B 0.011912f
C339 VTAIL.n71 B 0.021535f
C340 VTAIL.n72 B 0.011912f
C341 VTAIL.n73 B 0.011572f
C342 VTAIL.n74 B 0.027352f
C343 VTAIL.n75 B 0.027352f
C344 VTAIL.n76 B 0.012253f
C345 VTAIL.n77 B 0.021535f
C346 VTAIL.n78 B 0.011572f
C347 VTAIL.n79 B 0.027352f
C348 VTAIL.n80 B 0.012253f
C349 VTAIL.n81 B 1.02318f
C350 VTAIL.n82 B 0.011572f
C351 VTAIL.t2 B 0.046119f
C352 VTAIL.n83 B 0.149808f
C353 VTAIL.n84 B 0.019336f
C354 VTAIL.n85 B 0.020514f
C355 VTAIL.n86 B 0.027352f
C356 VTAIL.n87 B 0.012253f
C357 VTAIL.n88 B 0.011572f
C358 VTAIL.n89 B 0.021535f
C359 VTAIL.n90 B 0.021535f
C360 VTAIL.n91 B 0.011572f
C361 VTAIL.n92 B 0.012253f
C362 VTAIL.n93 B 0.027352f
C363 VTAIL.n94 B 0.027352f
C364 VTAIL.n95 B 0.012253f
C365 VTAIL.n96 B 0.011572f
C366 VTAIL.n97 B 0.021535f
C367 VTAIL.n98 B 0.021535f
C368 VTAIL.n99 B 0.011572f
C369 VTAIL.n100 B 0.012253f
C370 VTAIL.n101 B 0.027352f
C371 VTAIL.n102 B 0.027352f
C372 VTAIL.n103 B 0.012253f
C373 VTAIL.n104 B 0.011572f
C374 VTAIL.n105 B 0.021535f
C375 VTAIL.n106 B 0.021535f
C376 VTAIL.n107 B 0.011572f
C377 VTAIL.n108 B 0.012253f
C378 VTAIL.n109 B 0.027352f
C379 VTAIL.n110 B 0.027352f
C380 VTAIL.n111 B 0.012253f
C381 VTAIL.n112 B 0.011572f
C382 VTAIL.n113 B 0.021535f
C383 VTAIL.n114 B 0.021535f
C384 VTAIL.n115 B 0.011572f
C385 VTAIL.n116 B 0.012253f
C386 VTAIL.n117 B 0.027352f
C387 VTAIL.n118 B 0.056643f
C388 VTAIL.n119 B 0.012253f
C389 VTAIL.n120 B 0.011572f
C390 VTAIL.n121 B 0.048012f
C391 VTAIL.n122 B 0.031375f
C392 VTAIL.n123 B 1.65646f
C393 VTAIL.n124 B 0.028816f
C394 VTAIL.n125 B 0.021535f
C395 VTAIL.n126 B 0.011572f
C396 VTAIL.n127 B 0.027352f
C397 VTAIL.n128 B 0.012253f
C398 VTAIL.n129 B 0.021535f
C399 VTAIL.n130 B 0.011572f
C400 VTAIL.n131 B 0.027352f
C401 VTAIL.n132 B 0.011912f
C402 VTAIL.n133 B 0.021535f
C403 VTAIL.n134 B 0.011912f
C404 VTAIL.n135 B 0.011572f
C405 VTAIL.n136 B 0.027352f
C406 VTAIL.n137 B 0.027352f
C407 VTAIL.n138 B 0.012253f
C408 VTAIL.n139 B 0.021535f
C409 VTAIL.n140 B 0.011572f
C410 VTAIL.n141 B 0.027352f
C411 VTAIL.n142 B 0.012253f
C412 VTAIL.n143 B 1.02318f
C413 VTAIL.n144 B 0.011572f
C414 VTAIL.t3 B 0.046119f
C415 VTAIL.n145 B 0.149808f
C416 VTAIL.n146 B 0.019336f
C417 VTAIL.n147 B 0.020514f
C418 VTAIL.n148 B 0.027352f
C419 VTAIL.n149 B 0.012253f
C420 VTAIL.n150 B 0.011572f
C421 VTAIL.n151 B 0.021535f
C422 VTAIL.n152 B 0.021535f
C423 VTAIL.n153 B 0.011572f
C424 VTAIL.n154 B 0.012253f
C425 VTAIL.n155 B 0.027352f
C426 VTAIL.n156 B 0.027352f
C427 VTAIL.n157 B 0.012253f
C428 VTAIL.n158 B 0.011572f
C429 VTAIL.n159 B 0.021535f
C430 VTAIL.n160 B 0.021535f
C431 VTAIL.n161 B 0.011572f
C432 VTAIL.n162 B 0.012253f
C433 VTAIL.n163 B 0.027352f
C434 VTAIL.n164 B 0.027352f
C435 VTAIL.n165 B 0.012253f
C436 VTAIL.n166 B 0.011572f
C437 VTAIL.n167 B 0.021535f
C438 VTAIL.n168 B 0.021535f
C439 VTAIL.n169 B 0.011572f
C440 VTAIL.n170 B 0.012253f
C441 VTAIL.n171 B 0.027352f
C442 VTAIL.n172 B 0.027352f
C443 VTAIL.n173 B 0.012253f
C444 VTAIL.n174 B 0.011572f
C445 VTAIL.n175 B 0.021535f
C446 VTAIL.n176 B 0.021535f
C447 VTAIL.n177 B 0.011572f
C448 VTAIL.n178 B 0.012253f
C449 VTAIL.n179 B 0.027352f
C450 VTAIL.n180 B 0.056643f
C451 VTAIL.n181 B 0.012253f
C452 VTAIL.n182 B 0.011572f
C453 VTAIL.n183 B 0.048012f
C454 VTAIL.n184 B 0.031375f
C455 VTAIL.n185 B 1.40222f
C456 VTAIL.n186 B 0.028816f
C457 VTAIL.n187 B 0.021535f
C458 VTAIL.n188 B 0.011572f
C459 VTAIL.n189 B 0.027352f
C460 VTAIL.n190 B 0.012253f
C461 VTAIL.n191 B 0.021535f
C462 VTAIL.n192 B 0.011572f
C463 VTAIL.n193 B 0.027352f
C464 VTAIL.n194 B 0.011912f
C465 VTAIL.n195 B 0.021535f
C466 VTAIL.n196 B 0.012253f
C467 VTAIL.n197 B 0.027352f
C468 VTAIL.n198 B 0.012253f
C469 VTAIL.n199 B 0.021535f
C470 VTAIL.n200 B 0.011572f
C471 VTAIL.n201 B 0.027352f
C472 VTAIL.n202 B 0.012253f
C473 VTAIL.n203 B 1.02318f
C474 VTAIL.n204 B 0.011572f
C475 VTAIL.t1 B 0.046119f
C476 VTAIL.n205 B 0.149808f
C477 VTAIL.n206 B 0.019336f
C478 VTAIL.n207 B 0.020514f
C479 VTAIL.n208 B 0.027352f
C480 VTAIL.n209 B 0.012253f
C481 VTAIL.n210 B 0.011572f
C482 VTAIL.n211 B 0.021535f
C483 VTAIL.n212 B 0.021535f
C484 VTAIL.n213 B 0.011572f
C485 VTAIL.n214 B 0.012253f
C486 VTAIL.n215 B 0.027352f
C487 VTAIL.n216 B 0.027352f
C488 VTAIL.n217 B 0.012253f
C489 VTAIL.n218 B 0.011572f
C490 VTAIL.n219 B 0.021535f
C491 VTAIL.n220 B 0.021535f
C492 VTAIL.n221 B 0.011572f
C493 VTAIL.n222 B 0.011572f
C494 VTAIL.n223 B 0.012253f
C495 VTAIL.n224 B 0.027352f
C496 VTAIL.n225 B 0.027352f
C497 VTAIL.n226 B 0.027352f
C498 VTAIL.n227 B 0.011912f
C499 VTAIL.n228 B 0.011572f
C500 VTAIL.n229 B 0.021535f
C501 VTAIL.n230 B 0.021535f
C502 VTAIL.n231 B 0.011572f
C503 VTAIL.n232 B 0.012253f
C504 VTAIL.n233 B 0.027352f
C505 VTAIL.n234 B 0.027352f
C506 VTAIL.n235 B 0.012253f
C507 VTAIL.n236 B 0.011572f
C508 VTAIL.n237 B 0.021535f
C509 VTAIL.n238 B 0.021535f
C510 VTAIL.n239 B 0.011572f
C511 VTAIL.n240 B 0.012253f
C512 VTAIL.n241 B 0.027352f
C513 VTAIL.n242 B 0.056643f
C514 VTAIL.n243 B 0.012253f
C515 VTAIL.n244 B 0.011572f
C516 VTAIL.n245 B 0.048012f
C517 VTAIL.n246 B 0.031375f
C518 VTAIL.n247 B 1.30203f
C519 VN.t0 B 3.35042f
C520 VN.t1 B 4.05501f
.ends

