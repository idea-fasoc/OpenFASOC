* NGSPICE file created from diff_pair_sample_0986.ext - technology: sky130A

.subckt diff_pair_sample_0986 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=0 ps=0 w=6.23 l=1.65
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=2.4297 ps=13.24 w=6.23 l=1.65
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=0 ps=0 w=6.23 l=1.65
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=0 ps=0 w=6.23 l=1.65
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=2.4297 ps=13.24 w=6.23 l=1.65
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=0 ps=0 w=6.23 l=1.65
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=2.4297 ps=13.24 w=6.23 l=1.65
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4297 pd=13.24 as=2.4297 ps=13.24 w=6.23 l=1.65
R0 B.n461 B.n460 585
R1 B.n462 B.n461 585
R2 B.n187 B.n69 585
R3 B.n186 B.n185 585
R4 B.n184 B.n183 585
R5 B.n182 B.n181 585
R6 B.n180 B.n179 585
R7 B.n178 B.n177 585
R8 B.n176 B.n175 585
R9 B.n174 B.n173 585
R10 B.n172 B.n171 585
R11 B.n170 B.n169 585
R12 B.n168 B.n167 585
R13 B.n166 B.n165 585
R14 B.n164 B.n163 585
R15 B.n162 B.n161 585
R16 B.n160 B.n159 585
R17 B.n158 B.n157 585
R18 B.n156 B.n155 585
R19 B.n154 B.n153 585
R20 B.n152 B.n151 585
R21 B.n150 B.n149 585
R22 B.n148 B.n147 585
R23 B.n146 B.n145 585
R24 B.n144 B.n143 585
R25 B.n142 B.n141 585
R26 B.n140 B.n139 585
R27 B.n138 B.n137 585
R28 B.n136 B.n135 585
R29 B.n134 B.n133 585
R30 B.n132 B.n131 585
R31 B.n130 B.n129 585
R32 B.n128 B.n127 585
R33 B.n126 B.n125 585
R34 B.n124 B.n123 585
R35 B.n121 B.n120 585
R36 B.n119 B.n118 585
R37 B.n117 B.n116 585
R38 B.n115 B.n114 585
R39 B.n113 B.n112 585
R40 B.n111 B.n110 585
R41 B.n109 B.n108 585
R42 B.n107 B.n106 585
R43 B.n105 B.n104 585
R44 B.n103 B.n102 585
R45 B.n101 B.n100 585
R46 B.n99 B.n98 585
R47 B.n97 B.n96 585
R48 B.n95 B.n94 585
R49 B.n93 B.n92 585
R50 B.n91 B.n90 585
R51 B.n89 B.n88 585
R52 B.n87 B.n86 585
R53 B.n85 B.n84 585
R54 B.n83 B.n82 585
R55 B.n81 B.n80 585
R56 B.n79 B.n78 585
R57 B.n77 B.n76 585
R58 B.n40 B.n39 585
R59 B.n465 B.n464 585
R60 B.n459 B.n70 585
R61 B.n70 B.n37 585
R62 B.n458 B.n36 585
R63 B.n469 B.n36 585
R64 B.n457 B.n35 585
R65 B.n470 B.n35 585
R66 B.n456 B.n34 585
R67 B.n471 B.n34 585
R68 B.n455 B.n454 585
R69 B.n454 B.n30 585
R70 B.n453 B.n29 585
R71 B.n477 B.n29 585
R72 B.n452 B.n28 585
R73 B.n478 B.n28 585
R74 B.n451 B.n27 585
R75 B.n479 B.n27 585
R76 B.n450 B.n449 585
R77 B.n449 B.n23 585
R78 B.n448 B.n22 585
R79 B.n485 B.n22 585
R80 B.n447 B.n21 585
R81 B.n486 B.n21 585
R82 B.n446 B.n20 585
R83 B.n487 B.n20 585
R84 B.n445 B.n444 585
R85 B.n444 B.n16 585
R86 B.n443 B.n15 585
R87 B.n493 B.n15 585
R88 B.n442 B.n14 585
R89 B.n494 B.n14 585
R90 B.n441 B.n13 585
R91 B.n495 B.n13 585
R92 B.n440 B.n439 585
R93 B.n439 B.n12 585
R94 B.n438 B.n437 585
R95 B.n438 B.n8 585
R96 B.n436 B.n7 585
R97 B.n502 B.n7 585
R98 B.n435 B.n6 585
R99 B.n503 B.n6 585
R100 B.n434 B.n5 585
R101 B.n504 B.n5 585
R102 B.n433 B.n432 585
R103 B.n432 B.n4 585
R104 B.n431 B.n188 585
R105 B.n431 B.n430 585
R106 B.n421 B.n189 585
R107 B.n190 B.n189 585
R108 B.n423 B.n422 585
R109 B.n424 B.n423 585
R110 B.n420 B.n194 585
R111 B.n198 B.n194 585
R112 B.n419 B.n418 585
R113 B.n418 B.n417 585
R114 B.n196 B.n195 585
R115 B.n197 B.n196 585
R116 B.n410 B.n409 585
R117 B.n411 B.n410 585
R118 B.n408 B.n203 585
R119 B.n203 B.n202 585
R120 B.n407 B.n406 585
R121 B.n406 B.n405 585
R122 B.n205 B.n204 585
R123 B.n206 B.n205 585
R124 B.n398 B.n397 585
R125 B.n399 B.n398 585
R126 B.n396 B.n211 585
R127 B.n211 B.n210 585
R128 B.n395 B.n394 585
R129 B.n394 B.n393 585
R130 B.n213 B.n212 585
R131 B.n214 B.n213 585
R132 B.n386 B.n385 585
R133 B.n387 B.n386 585
R134 B.n384 B.n219 585
R135 B.n219 B.n218 585
R136 B.n383 B.n382 585
R137 B.n382 B.n381 585
R138 B.n221 B.n220 585
R139 B.n222 B.n221 585
R140 B.n377 B.n376 585
R141 B.n225 B.n224 585
R142 B.n373 B.n372 585
R143 B.n374 B.n373 585
R144 B.n371 B.n254 585
R145 B.n370 B.n369 585
R146 B.n368 B.n367 585
R147 B.n366 B.n365 585
R148 B.n364 B.n363 585
R149 B.n362 B.n361 585
R150 B.n360 B.n359 585
R151 B.n358 B.n357 585
R152 B.n356 B.n355 585
R153 B.n354 B.n353 585
R154 B.n352 B.n351 585
R155 B.n350 B.n349 585
R156 B.n348 B.n347 585
R157 B.n346 B.n345 585
R158 B.n344 B.n343 585
R159 B.n342 B.n341 585
R160 B.n340 B.n339 585
R161 B.n338 B.n337 585
R162 B.n336 B.n335 585
R163 B.n334 B.n333 585
R164 B.n332 B.n331 585
R165 B.n330 B.n329 585
R166 B.n328 B.n327 585
R167 B.n326 B.n325 585
R168 B.n324 B.n323 585
R169 B.n322 B.n321 585
R170 B.n320 B.n319 585
R171 B.n318 B.n317 585
R172 B.n316 B.n315 585
R173 B.n314 B.n313 585
R174 B.n312 B.n311 585
R175 B.n309 B.n308 585
R176 B.n307 B.n306 585
R177 B.n305 B.n304 585
R178 B.n303 B.n302 585
R179 B.n301 B.n300 585
R180 B.n299 B.n298 585
R181 B.n297 B.n296 585
R182 B.n295 B.n294 585
R183 B.n293 B.n292 585
R184 B.n291 B.n290 585
R185 B.n289 B.n288 585
R186 B.n287 B.n286 585
R187 B.n285 B.n284 585
R188 B.n283 B.n282 585
R189 B.n281 B.n280 585
R190 B.n279 B.n278 585
R191 B.n277 B.n276 585
R192 B.n275 B.n274 585
R193 B.n273 B.n272 585
R194 B.n271 B.n270 585
R195 B.n269 B.n268 585
R196 B.n267 B.n266 585
R197 B.n265 B.n264 585
R198 B.n263 B.n262 585
R199 B.n261 B.n260 585
R200 B.n378 B.n223 585
R201 B.n223 B.n222 585
R202 B.n380 B.n379 585
R203 B.n381 B.n380 585
R204 B.n217 B.n216 585
R205 B.n218 B.n217 585
R206 B.n389 B.n388 585
R207 B.n388 B.n387 585
R208 B.n390 B.n215 585
R209 B.n215 B.n214 585
R210 B.n392 B.n391 585
R211 B.n393 B.n392 585
R212 B.n209 B.n208 585
R213 B.n210 B.n209 585
R214 B.n401 B.n400 585
R215 B.n400 B.n399 585
R216 B.n402 B.n207 585
R217 B.n207 B.n206 585
R218 B.n404 B.n403 585
R219 B.n405 B.n404 585
R220 B.n201 B.n200 585
R221 B.n202 B.n201 585
R222 B.n413 B.n412 585
R223 B.n412 B.n411 585
R224 B.n414 B.n199 585
R225 B.n199 B.n197 585
R226 B.n416 B.n415 585
R227 B.n417 B.n416 585
R228 B.n193 B.n192 585
R229 B.n198 B.n193 585
R230 B.n426 B.n425 585
R231 B.n425 B.n424 585
R232 B.n427 B.n191 585
R233 B.n191 B.n190 585
R234 B.n429 B.n428 585
R235 B.n430 B.n429 585
R236 B.n3 B.n0 585
R237 B.n4 B.n3 585
R238 B.n501 B.n1 585
R239 B.n502 B.n501 585
R240 B.n500 B.n499 585
R241 B.n500 B.n8 585
R242 B.n498 B.n9 585
R243 B.n12 B.n9 585
R244 B.n497 B.n496 585
R245 B.n496 B.n495 585
R246 B.n11 B.n10 585
R247 B.n494 B.n11 585
R248 B.n492 B.n491 585
R249 B.n493 B.n492 585
R250 B.n490 B.n17 585
R251 B.n17 B.n16 585
R252 B.n489 B.n488 585
R253 B.n488 B.n487 585
R254 B.n19 B.n18 585
R255 B.n486 B.n19 585
R256 B.n484 B.n483 585
R257 B.n485 B.n484 585
R258 B.n482 B.n24 585
R259 B.n24 B.n23 585
R260 B.n481 B.n480 585
R261 B.n480 B.n479 585
R262 B.n26 B.n25 585
R263 B.n478 B.n26 585
R264 B.n476 B.n475 585
R265 B.n477 B.n476 585
R266 B.n474 B.n31 585
R267 B.n31 B.n30 585
R268 B.n473 B.n472 585
R269 B.n472 B.n471 585
R270 B.n33 B.n32 585
R271 B.n470 B.n33 585
R272 B.n468 B.n467 585
R273 B.n469 B.n468 585
R274 B.n466 B.n38 585
R275 B.n38 B.n37 585
R276 B.n505 B.n504 585
R277 B.n503 B.n2 585
R278 B.n464 B.n38 530.939
R279 B.n461 B.n70 530.939
R280 B.n260 B.n221 530.939
R281 B.n376 B.n223 530.939
R282 B.n74 B.t6 296.954
R283 B.n71 B.t2 296.954
R284 B.n258 B.t9 296.954
R285 B.n255 B.t13 296.954
R286 B.n462 B.n68 256.663
R287 B.n462 B.n67 256.663
R288 B.n462 B.n66 256.663
R289 B.n462 B.n65 256.663
R290 B.n462 B.n64 256.663
R291 B.n462 B.n63 256.663
R292 B.n462 B.n62 256.663
R293 B.n462 B.n61 256.663
R294 B.n462 B.n60 256.663
R295 B.n462 B.n59 256.663
R296 B.n462 B.n58 256.663
R297 B.n462 B.n57 256.663
R298 B.n462 B.n56 256.663
R299 B.n462 B.n55 256.663
R300 B.n462 B.n54 256.663
R301 B.n462 B.n53 256.663
R302 B.n462 B.n52 256.663
R303 B.n462 B.n51 256.663
R304 B.n462 B.n50 256.663
R305 B.n462 B.n49 256.663
R306 B.n462 B.n48 256.663
R307 B.n462 B.n47 256.663
R308 B.n462 B.n46 256.663
R309 B.n462 B.n45 256.663
R310 B.n462 B.n44 256.663
R311 B.n462 B.n43 256.663
R312 B.n462 B.n42 256.663
R313 B.n462 B.n41 256.663
R314 B.n463 B.n462 256.663
R315 B.n375 B.n374 256.663
R316 B.n374 B.n226 256.663
R317 B.n374 B.n227 256.663
R318 B.n374 B.n228 256.663
R319 B.n374 B.n229 256.663
R320 B.n374 B.n230 256.663
R321 B.n374 B.n231 256.663
R322 B.n374 B.n232 256.663
R323 B.n374 B.n233 256.663
R324 B.n374 B.n234 256.663
R325 B.n374 B.n235 256.663
R326 B.n374 B.n236 256.663
R327 B.n374 B.n237 256.663
R328 B.n374 B.n238 256.663
R329 B.n374 B.n239 256.663
R330 B.n374 B.n240 256.663
R331 B.n374 B.n241 256.663
R332 B.n374 B.n242 256.663
R333 B.n374 B.n243 256.663
R334 B.n374 B.n244 256.663
R335 B.n374 B.n245 256.663
R336 B.n374 B.n246 256.663
R337 B.n374 B.n247 256.663
R338 B.n374 B.n248 256.663
R339 B.n374 B.n249 256.663
R340 B.n374 B.n250 256.663
R341 B.n374 B.n251 256.663
R342 B.n374 B.n252 256.663
R343 B.n374 B.n253 256.663
R344 B.n507 B.n506 256.663
R345 B.n76 B.n40 163.367
R346 B.n80 B.n79 163.367
R347 B.n84 B.n83 163.367
R348 B.n88 B.n87 163.367
R349 B.n92 B.n91 163.367
R350 B.n96 B.n95 163.367
R351 B.n100 B.n99 163.367
R352 B.n104 B.n103 163.367
R353 B.n108 B.n107 163.367
R354 B.n112 B.n111 163.367
R355 B.n116 B.n115 163.367
R356 B.n120 B.n119 163.367
R357 B.n125 B.n124 163.367
R358 B.n129 B.n128 163.367
R359 B.n133 B.n132 163.367
R360 B.n137 B.n136 163.367
R361 B.n141 B.n140 163.367
R362 B.n145 B.n144 163.367
R363 B.n149 B.n148 163.367
R364 B.n153 B.n152 163.367
R365 B.n157 B.n156 163.367
R366 B.n161 B.n160 163.367
R367 B.n165 B.n164 163.367
R368 B.n169 B.n168 163.367
R369 B.n173 B.n172 163.367
R370 B.n177 B.n176 163.367
R371 B.n181 B.n180 163.367
R372 B.n185 B.n184 163.367
R373 B.n461 B.n69 163.367
R374 B.n382 B.n221 163.367
R375 B.n382 B.n219 163.367
R376 B.n386 B.n219 163.367
R377 B.n386 B.n213 163.367
R378 B.n394 B.n213 163.367
R379 B.n394 B.n211 163.367
R380 B.n398 B.n211 163.367
R381 B.n398 B.n205 163.367
R382 B.n406 B.n205 163.367
R383 B.n406 B.n203 163.367
R384 B.n410 B.n203 163.367
R385 B.n410 B.n196 163.367
R386 B.n418 B.n196 163.367
R387 B.n418 B.n194 163.367
R388 B.n423 B.n194 163.367
R389 B.n423 B.n189 163.367
R390 B.n431 B.n189 163.367
R391 B.n432 B.n431 163.367
R392 B.n432 B.n5 163.367
R393 B.n6 B.n5 163.367
R394 B.n7 B.n6 163.367
R395 B.n438 B.n7 163.367
R396 B.n439 B.n438 163.367
R397 B.n439 B.n13 163.367
R398 B.n14 B.n13 163.367
R399 B.n15 B.n14 163.367
R400 B.n444 B.n15 163.367
R401 B.n444 B.n20 163.367
R402 B.n21 B.n20 163.367
R403 B.n22 B.n21 163.367
R404 B.n449 B.n22 163.367
R405 B.n449 B.n27 163.367
R406 B.n28 B.n27 163.367
R407 B.n29 B.n28 163.367
R408 B.n454 B.n29 163.367
R409 B.n454 B.n34 163.367
R410 B.n35 B.n34 163.367
R411 B.n36 B.n35 163.367
R412 B.n70 B.n36 163.367
R413 B.n373 B.n225 163.367
R414 B.n373 B.n254 163.367
R415 B.n369 B.n368 163.367
R416 B.n365 B.n364 163.367
R417 B.n361 B.n360 163.367
R418 B.n357 B.n356 163.367
R419 B.n353 B.n352 163.367
R420 B.n349 B.n348 163.367
R421 B.n345 B.n344 163.367
R422 B.n341 B.n340 163.367
R423 B.n337 B.n336 163.367
R424 B.n333 B.n332 163.367
R425 B.n329 B.n328 163.367
R426 B.n325 B.n324 163.367
R427 B.n321 B.n320 163.367
R428 B.n317 B.n316 163.367
R429 B.n313 B.n312 163.367
R430 B.n308 B.n307 163.367
R431 B.n304 B.n303 163.367
R432 B.n300 B.n299 163.367
R433 B.n296 B.n295 163.367
R434 B.n292 B.n291 163.367
R435 B.n288 B.n287 163.367
R436 B.n284 B.n283 163.367
R437 B.n280 B.n279 163.367
R438 B.n276 B.n275 163.367
R439 B.n272 B.n271 163.367
R440 B.n268 B.n267 163.367
R441 B.n264 B.n263 163.367
R442 B.n380 B.n223 163.367
R443 B.n380 B.n217 163.367
R444 B.n388 B.n217 163.367
R445 B.n388 B.n215 163.367
R446 B.n392 B.n215 163.367
R447 B.n392 B.n209 163.367
R448 B.n400 B.n209 163.367
R449 B.n400 B.n207 163.367
R450 B.n404 B.n207 163.367
R451 B.n404 B.n201 163.367
R452 B.n412 B.n201 163.367
R453 B.n412 B.n199 163.367
R454 B.n416 B.n199 163.367
R455 B.n416 B.n193 163.367
R456 B.n425 B.n193 163.367
R457 B.n425 B.n191 163.367
R458 B.n429 B.n191 163.367
R459 B.n429 B.n3 163.367
R460 B.n505 B.n3 163.367
R461 B.n501 B.n2 163.367
R462 B.n501 B.n500 163.367
R463 B.n500 B.n9 163.367
R464 B.n496 B.n9 163.367
R465 B.n496 B.n11 163.367
R466 B.n492 B.n11 163.367
R467 B.n492 B.n17 163.367
R468 B.n488 B.n17 163.367
R469 B.n488 B.n19 163.367
R470 B.n484 B.n19 163.367
R471 B.n484 B.n24 163.367
R472 B.n480 B.n24 163.367
R473 B.n480 B.n26 163.367
R474 B.n476 B.n26 163.367
R475 B.n476 B.n31 163.367
R476 B.n472 B.n31 163.367
R477 B.n472 B.n33 163.367
R478 B.n468 B.n33 163.367
R479 B.n468 B.n38 163.367
R480 B.n374 B.n222 134.811
R481 B.n462 B.n37 134.811
R482 B.n71 B.t4 109.855
R483 B.n258 B.t12 109.855
R484 B.n74 B.t7 109.847
R485 B.n255 B.t15 109.847
R486 B.n464 B.n463 71.676
R487 B.n76 B.n41 71.676
R488 B.n80 B.n42 71.676
R489 B.n84 B.n43 71.676
R490 B.n88 B.n44 71.676
R491 B.n92 B.n45 71.676
R492 B.n96 B.n46 71.676
R493 B.n100 B.n47 71.676
R494 B.n104 B.n48 71.676
R495 B.n108 B.n49 71.676
R496 B.n112 B.n50 71.676
R497 B.n116 B.n51 71.676
R498 B.n120 B.n52 71.676
R499 B.n125 B.n53 71.676
R500 B.n129 B.n54 71.676
R501 B.n133 B.n55 71.676
R502 B.n137 B.n56 71.676
R503 B.n141 B.n57 71.676
R504 B.n145 B.n58 71.676
R505 B.n149 B.n59 71.676
R506 B.n153 B.n60 71.676
R507 B.n157 B.n61 71.676
R508 B.n161 B.n62 71.676
R509 B.n165 B.n63 71.676
R510 B.n169 B.n64 71.676
R511 B.n173 B.n65 71.676
R512 B.n177 B.n66 71.676
R513 B.n181 B.n67 71.676
R514 B.n185 B.n68 71.676
R515 B.n69 B.n68 71.676
R516 B.n184 B.n67 71.676
R517 B.n180 B.n66 71.676
R518 B.n176 B.n65 71.676
R519 B.n172 B.n64 71.676
R520 B.n168 B.n63 71.676
R521 B.n164 B.n62 71.676
R522 B.n160 B.n61 71.676
R523 B.n156 B.n60 71.676
R524 B.n152 B.n59 71.676
R525 B.n148 B.n58 71.676
R526 B.n144 B.n57 71.676
R527 B.n140 B.n56 71.676
R528 B.n136 B.n55 71.676
R529 B.n132 B.n54 71.676
R530 B.n128 B.n53 71.676
R531 B.n124 B.n52 71.676
R532 B.n119 B.n51 71.676
R533 B.n115 B.n50 71.676
R534 B.n111 B.n49 71.676
R535 B.n107 B.n48 71.676
R536 B.n103 B.n47 71.676
R537 B.n99 B.n46 71.676
R538 B.n95 B.n45 71.676
R539 B.n91 B.n44 71.676
R540 B.n87 B.n43 71.676
R541 B.n83 B.n42 71.676
R542 B.n79 B.n41 71.676
R543 B.n463 B.n40 71.676
R544 B.n376 B.n375 71.676
R545 B.n254 B.n226 71.676
R546 B.n368 B.n227 71.676
R547 B.n364 B.n228 71.676
R548 B.n360 B.n229 71.676
R549 B.n356 B.n230 71.676
R550 B.n352 B.n231 71.676
R551 B.n348 B.n232 71.676
R552 B.n344 B.n233 71.676
R553 B.n340 B.n234 71.676
R554 B.n336 B.n235 71.676
R555 B.n332 B.n236 71.676
R556 B.n328 B.n237 71.676
R557 B.n324 B.n238 71.676
R558 B.n320 B.n239 71.676
R559 B.n316 B.n240 71.676
R560 B.n312 B.n241 71.676
R561 B.n307 B.n242 71.676
R562 B.n303 B.n243 71.676
R563 B.n299 B.n244 71.676
R564 B.n295 B.n245 71.676
R565 B.n291 B.n246 71.676
R566 B.n287 B.n247 71.676
R567 B.n283 B.n248 71.676
R568 B.n279 B.n249 71.676
R569 B.n275 B.n250 71.676
R570 B.n271 B.n251 71.676
R571 B.n267 B.n252 71.676
R572 B.n263 B.n253 71.676
R573 B.n375 B.n225 71.676
R574 B.n369 B.n226 71.676
R575 B.n365 B.n227 71.676
R576 B.n361 B.n228 71.676
R577 B.n357 B.n229 71.676
R578 B.n353 B.n230 71.676
R579 B.n349 B.n231 71.676
R580 B.n345 B.n232 71.676
R581 B.n341 B.n233 71.676
R582 B.n337 B.n234 71.676
R583 B.n333 B.n235 71.676
R584 B.n329 B.n236 71.676
R585 B.n325 B.n237 71.676
R586 B.n321 B.n238 71.676
R587 B.n317 B.n239 71.676
R588 B.n313 B.n240 71.676
R589 B.n308 B.n241 71.676
R590 B.n304 B.n242 71.676
R591 B.n300 B.n243 71.676
R592 B.n296 B.n244 71.676
R593 B.n292 B.n245 71.676
R594 B.n288 B.n246 71.676
R595 B.n284 B.n247 71.676
R596 B.n280 B.n248 71.676
R597 B.n276 B.n249 71.676
R598 B.n272 B.n250 71.676
R599 B.n268 B.n251 71.676
R600 B.n264 B.n252 71.676
R601 B.n260 B.n253 71.676
R602 B.n506 B.n505 71.676
R603 B.n506 B.n2 71.676
R604 B.n72 B.t5 71.4546
R605 B.n259 B.t11 71.4546
R606 B.n75 B.t8 71.4479
R607 B.n256 B.t14 71.4479
R608 B.n381 B.n222 65.0157
R609 B.n381 B.n218 65.0157
R610 B.n387 B.n218 65.0157
R611 B.n387 B.n214 65.0157
R612 B.n393 B.n214 65.0157
R613 B.n399 B.n210 65.0157
R614 B.n399 B.n206 65.0157
R615 B.n405 B.n206 65.0157
R616 B.n405 B.n202 65.0157
R617 B.n411 B.n202 65.0157
R618 B.n411 B.n197 65.0157
R619 B.n417 B.n197 65.0157
R620 B.n417 B.n198 65.0157
R621 B.n424 B.n190 65.0157
R622 B.n430 B.n190 65.0157
R623 B.n430 B.n4 65.0157
R624 B.n504 B.n4 65.0157
R625 B.n504 B.n503 65.0157
R626 B.n503 B.n502 65.0157
R627 B.n502 B.n8 65.0157
R628 B.n12 B.n8 65.0157
R629 B.n495 B.n12 65.0157
R630 B.n494 B.n493 65.0157
R631 B.n493 B.n16 65.0157
R632 B.n487 B.n16 65.0157
R633 B.n487 B.n486 65.0157
R634 B.n486 B.n485 65.0157
R635 B.n485 B.n23 65.0157
R636 B.n479 B.n23 65.0157
R637 B.n479 B.n478 65.0157
R638 B.n477 B.n30 65.0157
R639 B.n471 B.n30 65.0157
R640 B.n471 B.n470 65.0157
R641 B.n470 B.n469 65.0157
R642 B.n469 B.n37 65.0157
R643 B.n198 B.t0 64.0596
R644 B.t1 B.n494 64.0596
R645 B.n393 B.t10 62.1474
R646 B.t3 B.n477 62.1474
R647 B.n122 B.n75 59.5399
R648 B.n73 B.n72 59.5399
R649 B.n310 B.n259 59.5399
R650 B.n257 B.n256 59.5399
R651 B.n75 B.n74 38.4005
R652 B.n72 B.n71 38.4005
R653 B.n259 B.n258 38.4005
R654 B.n256 B.n255 38.4005
R655 B.n378 B.n377 34.4981
R656 B.n261 B.n220 34.4981
R657 B.n460 B.n459 34.4981
R658 B.n466 B.n465 34.4981
R659 B B.n507 18.0485
R660 B.n379 B.n378 10.6151
R661 B.n379 B.n216 10.6151
R662 B.n389 B.n216 10.6151
R663 B.n390 B.n389 10.6151
R664 B.n391 B.n390 10.6151
R665 B.n391 B.n208 10.6151
R666 B.n401 B.n208 10.6151
R667 B.n402 B.n401 10.6151
R668 B.n403 B.n402 10.6151
R669 B.n403 B.n200 10.6151
R670 B.n413 B.n200 10.6151
R671 B.n414 B.n413 10.6151
R672 B.n415 B.n414 10.6151
R673 B.n415 B.n192 10.6151
R674 B.n426 B.n192 10.6151
R675 B.n427 B.n426 10.6151
R676 B.n428 B.n427 10.6151
R677 B.n428 B.n0 10.6151
R678 B.n377 B.n224 10.6151
R679 B.n372 B.n224 10.6151
R680 B.n372 B.n371 10.6151
R681 B.n371 B.n370 10.6151
R682 B.n370 B.n367 10.6151
R683 B.n367 B.n366 10.6151
R684 B.n366 B.n363 10.6151
R685 B.n363 B.n362 10.6151
R686 B.n362 B.n359 10.6151
R687 B.n359 B.n358 10.6151
R688 B.n358 B.n355 10.6151
R689 B.n355 B.n354 10.6151
R690 B.n354 B.n351 10.6151
R691 B.n351 B.n350 10.6151
R692 B.n350 B.n347 10.6151
R693 B.n347 B.n346 10.6151
R694 B.n346 B.n343 10.6151
R695 B.n343 B.n342 10.6151
R696 B.n342 B.n339 10.6151
R697 B.n339 B.n338 10.6151
R698 B.n338 B.n335 10.6151
R699 B.n335 B.n334 10.6151
R700 B.n334 B.n331 10.6151
R701 B.n331 B.n330 10.6151
R702 B.n327 B.n326 10.6151
R703 B.n326 B.n323 10.6151
R704 B.n323 B.n322 10.6151
R705 B.n322 B.n319 10.6151
R706 B.n319 B.n318 10.6151
R707 B.n318 B.n315 10.6151
R708 B.n315 B.n314 10.6151
R709 B.n314 B.n311 10.6151
R710 B.n309 B.n306 10.6151
R711 B.n306 B.n305 10.6151
R712 B.n305 B.n302 10.6151
R713 B.n302 B.n301 10.6151
R714 B.n301 B.n298 10.6151
R715 B.n298 B.n297 10.6151
R716 B.n297 B.n294 10.6151
R717 B.n294 B.n293 10.6151
R718 B.n293 B.n290 10.6151
R719 B.n290 B.n289 10.6151
R720 B.n289 B.n286 10.6151
R721 B.n286 B.n285 10.6151
R722 B.n285 B.n282 10.6151
R723 B.n282 B.n281 10.6151
R724 B.n281 B.n278 10.6151
R725 B.n278 B.n277 10.6151
R726 B.n277 B.n274 10.6151
R727 B.n274 B.n273 10.6151
R728 B.n273 B.n270 10.6151
R729 B.n270 B.n269 10.6151
R730 B.n269 B.n266 10.6151
R731 B.n266 B.n265 10.6151
R732 B.n265 B.n262 10.6151
R733 B.n262 B.n261 10.6151
R734 B.n383 B.n220 10.6151
R735 B.n384 B.n383 10.6151
R736 B.n385 B.n384 10.6151
R737 B.n385 B.n212 10.6151
R738 B.n395 B.n212 10.6151
R739 B.n396 B.n395 10.6151
R740 B.n397 B.n396 10.6151
R741 B.n397 B.n204 10.6151
R742 B.n407 B.n204 10.6151
R743 B.n408 B.n407 10.6151
R744 B.n409 B.n408 10.6151
R745 B.n409 B.n195 10.6151
R746 B.n419 B.n195 10.6151
R747 B.n420 B.n419 10.6151
R748 B.n422 B.n420 10.6151
R749 B.n422 B.n421 10.6151
R750 B.n421 B.n188 10.6151
R751 B.n433 B.n188 10.6151
R752 B.n434 B.n433 10.6151
R753 B.n435 B.n434 10.6151
R754 B.n436 B.n435 10.6151
R755 B.n437 B.n436 10.6151
R756 B.n440 B.n437 10.6151
R757 B.n441 B.n440 10.6151
R758 B.n442 B.n441 10.6151
R759 B.n443 B.n442 10.6151
R760 B.n445 B.n443 10.6151
R761 B.n446 B.n445 10.6151
R762 B.n447 B.n446 10.6151
R763 B.n448 B.n447 10.6151
R764 B.n450 B.n448 10.6151
R765 B.n451 B.n450 10.6151
R766 B.n452 B.n451 10.6151
R767 B.n453 B.n452 10.6151
R768 B.n455 B.n453 10.6151
R769 B.n456 B.n455 10.6151
R770 B.n457 B.n456 10.6151
R771 B.n458 B.n457 10.6151
R772 B.n459 B.n458 10.6151
R773 B.n499 B.n1 10.6151
R774 B.n499 B.n498 10.6151
R775 B.n498 B.n497 10.6151
R776 B.n497 B.n10 10.6151
R777 B.n491 B.n10 10.6151
R778 B.n491 B.n490 10.6151
R779 B.n490 B.n489 10.6151
R780 B.n489 B.n18 10.6151
R781 B.n483 B.n18 10.6151
R782 B.n483 B.n482 10.6151
R783 B.n482 B.n481 10.6151
R784 B.n481 B.n25 10.6151
R785 B.n475 B.n25 10.6151
R786 B.n475 B.n474 10.6151
R787 B.n474 B.n473 10.6151
R788 B.n473 B.n32 10.6151
R789 B.n467 B.n32 10.6151
R790 B.n467 B.n466 10.6151
R791 B.n465 B.n39 10.6151
R792 B.n77 B.n39 10.6151
R793 B.n78 B.n77 10.6151
R794 B.n81 B.n78 10.6151
R795 B.n82 B.n81 10.6151
R796 B.n85 B.n82 10.6151
R797 B.n86 B.n85 10.6151
R798 B.n89 B.n86 10.6151
R799 B.n90 B.n89 10.6151
R800 B.n93 B.n90 10.6151
R801 B.n94 B.n93 10.6151
R802 B.n97 B.n94 10.6151
R803 B.n98 B.n97 10.6151
R804 B.n101 B.n98 10.6151
R805 B.n102 B.n101 10.6151
R806 B.n105 B.n102 10.6151
R807 B.n106 B.n105 10.6151
R808 B.n109 B.n106 10.6151
R809 B.n110 B.n109 10.6151
R810 B.n113 B.n110 10.6151
R811 B.n114 B.n113 10.6151
R812 B.n117 B.n114 10.6151
R813 B.n118 B.n117 10.6151
R814 B.n121 B.n118 10.6151
R815 B.n126 B.n123 10.6151
R816 B.n127 B.n126 10.6151
R817 B.n130 B.n127 10.6151
R818 B.n131 B.n130 10.6151
R819 B.n134 B.n131 10.6151
R820 B.n135 B.n134 10.6151
R821 B.n138 B.n135 10.6151
R822 B.n139 B.n138 10.6151
R823 B.n143 B.n142 10.6151
R824 B.n146 B.n143 10.6151
R825 B.n147 B.n146 10.6151
R826 B.n150 B.n147 10.6151
R827 B.n151 B.n150 10.6151
R828 B.n154 B.n151 10.6151
R829 B.n155 B.n154 10.6151
R830 B.n158 B.n155 10.6151
R831 B.n159 B.n158 10.6151
R832 B.n162 B.n159 10.6151
R833 B.n163 B.n162 10.6151
R834 B.n166 B.n163 10.6151
R835 B.n167 B.n166 10.6151
R836 B.n170 B.n167 10.6151
R837 B.n171 B.n170 10.6151
R838 B.n174 B.n171 10.6151
R839 B.n175 B.n174 10.6151
R840 B.n178 B.n175 10.6151
R841 B.n179 B.n178 10.6151
R842 B.n182 B.n179 10.6151
R843 B.n183 B.n182 10.6151
R844 B.n186 B.n183 10.6151
R845 B.n187 B.n186 10.6151
R846 B.n460 B.n187 10.6151
R847 B.n507 B.n0 8.11757
R848 B.n507 B.n1 8.11757
R849 B.n327 B.n257 6.5566
R850 B.n311 B.n310 6.5566
R851 B.n123 B.n122 6.5566
R852 B.n139 B.n73 6.5566
R853 B.n330 B.n257 4.05904
R854 B.n310 B.n309 4.05904
R855 B.n122 B.n121 4.05904
R856 B.n142 B.n73 4.05904
R857 B.t10 B.n210 2.86882
R858 B.n478 B.t3 2.86882
R859 B.n424 B.t0 0.956606
R860 B.n495 B.t1 0.956606
R861 VP.n0 VP.t1 187.623
R862 VP.n0 VP.t0 149.857
R863 VP VP.n0 0.241678
R864 VTAIL.n1 VTAIL.t1 56.822
R865 VTAIL.n2 VTAIL.t2 56.8211
R866 VTAIL.n3 VTAIL.t0 56.821
R867 VTAIL.n0 VTAIL.t3 56.821
R868 VTAIL.n1 VTAIL.n0 21.1514
R869 VTAIL.n3 VTAIL.n2 19.4445
R870 VTAIL.n2 VTAIL.n1 1.32378
R871 VTAIL VTAIL.n0 0.955241
R872 VTAIL VTAIL.n3 0.369034
R873 VDD1 VDD1.t1 106.895
R874 VDD1 VDD1.t0 73.9848
R875 VN VN.t0 187.815
R876 VN VN.t1 150.099
R877 VDD2.n0 VDD2.t0 105.944
R878 VDD2.n0 VDD2.t1 73.4999
R879 VDD2 VDD2.n0 0.485414
C0 VTAIL VDD1 3.36553f
C1 VP VDD1 1.58909f
C2 VP VTAIL 1.37252f
C3 VDD2 VDD1 0.562087f
C4 VN VDD1 0.147686f
C5 VDD2 VTAIL 3.41038f
C6 VN VTAIL 1.35827f
C7 VP VDD2 0.292641f
C8 VN VP 3.94467f
C9 VN VDD2 1.44594f
C10 VDD2 B 3.028784f
C11 VDD1 B 4.78522f
C12 VTAIL B 4.441287f
C13 VN B 6.867401f
C14 VP B 4.740334f
C15 VDD2.t0 B 0.997665f
C16 VDD2.t1 B 0.768251f
C17 VDD2.n0 B 1.57109f
C18 VN.t1 B 0.810391f
C19 VN.t0 B 1.03691f
C20 VDD1.t0 B 0.757436f
C21 VDD1.t1 B 0.999433f
C22 VTAIL.t3 B 0.81203f
C23 VTAIL.n0 B 0.913302f
C24 VTAIL.t1 B 0.81203f
C25 VTAIL.n1 B 0.932554f
C26 VTAIL.t2 B 0.812026f
C27 VTAIL.n2 B 0.84339f
C28 VTAIL.t0 B 0.81203f
C29 VTAIL.n3 B 0.793512f
C30 VP.t1 B 1.0428f
C31 VP.t0 B 0.817117f
C32 VP.n0 B 2.00563f
.ends

