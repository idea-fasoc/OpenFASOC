* NGSPICE file created from diff_pair_sample_0539.ext - technology: sky130A

.subckt diff_pair_sample_0539 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=0 ps=0 w=9.26 l=3.52
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=3.6114 ps=19.3 w=9.26 l=3.52
X2 B.t8 B.t6 B.t7 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=0 ps=0 w=9.26 l=3.52
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=3.6114 ps=19.3 w=9.26 l=3.52
X4 B.t5 B.t3 B.t4 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=0 ps=0 w=9.26 l=3.52
X5 B.t2 B.t0 B.t1 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=0 ps=0 w=9.26 l=3.52
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=3.6114 ps=19.3 w=9.26 l=3.52
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n2510_n2820# sky130_fd_pr__pfet_01v8 ad=3.6114 pd=19.3 as=3.6114 ps=19.3 w=9.26 l=3.52
R0 B.n308 B.n91 585
R1 B.n307 B.n306 585
R2 B.n305 B.n92 585
R3 B.n304 B.n303 585
R4 B.n302 B.n93 585
R5 B.n301 B.n300 585
R6 B.n299 B.n94 585
R7 B.n298 B.n297 585
R8 B.n296 B.n95 585
R9 B.n295 B.n294 585
R10 B.n293 B.n96 585
R11 B.n292 B.n291 585
R12 B.n290 B.n97 585
R13 B.n289 B.n288 585
R14 B.n287 B.n98 585
R15 B.n286 B.n285 585
R16 B.n284 B.n99 585
R17 B.n283 B.n282 585
R18 B.n281 B.n100 585
R19 B.n280 B.n279 585
R20 B.n278 B.n101 585
R21 B.n277 B.n276 585
R22 B.n275 B.n102 585
R23 B.n274 B.n273 585
R24 B.n272 B.n103 585
R25 B.n271 B.n270 585
R26 B.n269 B.n104 585
R27 B.n268 B.n267 585
R28 B.n266 B.n105 585
R29 B.n265 B.n264 585
R30 B.n263 B.n106 585
R31 B.n262 B.n261 585
R32 B.n260 B.n107 585
R33 B.n259 B.n258 585
R34 B.n257 B.n256 585
R35 B.n255 B.n111 585
R36 B.n254 B.n253 585
R37 B.n252 B.n112 585
R38 B.n251 B.n250 585
R39 B.n249 B.n113 585
R40 B.n248 B.n247 585
R41 B.n246 B.n114 585
R42 B.n245 B.n244 585
R43 B.n242 B.n115 585
R44 B.n241 B.n240 585
R45 B.n239 B.n118 585
R46 B.n238 B.n237 585
R47 B.n236 B.n119 585
R48 B.n235 B.n234 585
R49 B.n233 B.n120 585
R50 B.n232 B.n231 585
R51 B.n230 B.n121 585
R52 B.n229 B.n228 585
R53 B.n227 B.n122 585
R54 B.n226 B.n225 585
R55 B.n224 B.n123 585
R56 B.n223 B.n222 585
R57 B.n221 B.n124 585
R58 B.n220 B.n219 585
R59 B.n218 B.n125 585
R60 B.n217 B.n216 585
R61 B.n215 B.n126 585
R62 B.n214 B.n213 585
R63 B.n212 B.n127 585
R64 B.n211 B.n210 585
R65 B.n209 B.n128 585
R66 B.n208 B.n207 585
R67 B.n206 B.n129 585
R68 B.n205 B.n204 585
R69 B.n203 B.n130 585
R70 B.n202 B.n201 585
R71 B.n200 B.n131 585
R72 B.n199 B.n198 585
R73 B.n197 B.n132 585
R74 B.n196 B.n195 585
R75 B.n194 B.n133 585
R76 B.n193 B.n192 585
R77 B.n310 B.n309 585
R78 B.n311 B.n90 585
R79 B.n313 B.n312 585
R80 B.n314 B.n89 585
R81 B.n316 B.n315 585
R82 B.n317 B.n88 585
R83 B.n319 B.n318 585
R84 B.n320 B.n87 585
R85 B.n322 B.n321 585
R86 B.n323 B.n86 585
R87 B.n325 B.n324 585
R88 B.n326 B.n85 585
R89 B.n328 B.n327 585
R90 B.n329 B.n84 585
R91 B.n331 B.n330 585
R92 B.n332 B.n83 585
R93 B.n334 B.n333 585
R94 B.n335 B.n82 585
R95 B.n337 B.n336 585
R96 B.n338 B.n81 585
R97 B.n340 B.n339 585
R98 B.n341 B.n80 585
R99 B.n343 B.n342 585
R100 B.n344 B.n79 585
R101 B.n346 B.n345 585
R102 B.n347 B.n78 585
R103 B.n349 B.n348 585
R104 B.n350 B.n77 585
R105 B.n352 B.n351 585
R106 B.n353 B.n76 585
R107 B.n355 B.n354 585
R108 B.n356 B.n75 585
R109 B.n358 B.n357 585
R110 B.n359 B.n74 585
R111 B.n361 B.n360 585
R112 B.n362 B.n73 585
R113 B.n364 B.n363 585
R114 B.n365 B.n72 585
R115 B.n367 B.n366 585
R116 B.n368 B.n71 585
R117 B.n370 B.n369 585
R118 B.n371 B.n70 585
R119 B.n373 B.n372 585
R120 B.n374 B.n69 585
R121 B.n376 B.n375 585
R122 B.n377 B.n68 585
R123 B.n379 B.n378 585
R124 B.n380 B.n67 585
R125 B.n382 B.n381 585
R126 B.n383 B.n66 585
R127 B.n385 B.n384 585
R128 B.n386 B.n65 585
R129 B.n388 B.n387 585
R130 B.n389 B.n64 585
R131 B.n391 B.n390 585
R132 B.n392 B.n63 585
R133 B.n394 B.n393 585
R134 B.n395 B.n62 585
R135 B.n397 B.n396 585
R136 B.n398 B.n61 585
R137 B.n400 B.n399 585
R138 B.n401 B.n60 585
R139 B.n518 B.n17 585
R140 B.n517 B.n516 585
R141 B.n515 B.n18 585
R142 B.n514 B.n513 585
R143 B.n512 B.n19 585
R144 B.n511 B.n510 585
R145 B.n509 B.n20 585
R146 B.n508 B.n507 585
R147 B.n506 B.n21 585
R148 B.n505 B.n504 585
R149 B.n503 B.n22 585
R150 B.n502 B.n501 585
R151 B.n500 B.n23 585
R152 B.n499 B.n498 585
R153 B.n497 B.n24 585
R154 B.n496 B.n495 585
R155 B.n494 B.n25 585
R156 B.n493 B.n492 585
R157 B.n491 B.n26 585
R158 B.n490 B.n489 585
R159 B.n488 B.n27 585
R160 B.n487 B.n486 585
R161 B.n485 B.n28 585
R162 B.n484 B.n483 585
R163 B.n482 B.n29 585
R164 B.n481 B.n480 585
R165 B.n479 B.n30 585
R166 B.n478 B.n477 585
R167 B.n476 B.n31 585
R168 B.n475 B.n474 585
R169 B.n473 B.n32 585
R170 B.n472 B.n471 585
R171 B.n470 B.n33 585
R172 B.n469 B.n468 585
R173 B.n467 B.n466 585
R174 B.n465 B.n37 585
R175 B.n464 B.n463 585
R176 B.n462 B.n38 585
R177 B.n461 B.n460 585
R178 B.n459 B.n39 585
R179 B.n458 B.n457 585
R180 B.n456 B.n40 585
R181 B.n455 B.n454 585
R182 B.n452 B.n41 585
R183 B.n451 B.n450 585
R184 B.n449 B.n44 585
R185 B.n448 B.n447 585
R186 B.n446 B.n45 585
R187 B.n445 B.n444 585
R188 B.n443 B.n46 585
R189 B.n442 B.n441 585
R190 B.n440 B.n47 585
R191 B.n439 B.n438 585
R192 B.n437 B.n48 585
R193 B.n436 B.n435 585
R194 B.n434 B.n49 585
R195 B.n433 B.n432 585
R196 B.n431 B.n50 585
R197 B.n430 B.n429 585
R198 B.n428 B.n51 585
R199 B.n427 B.n426 585
R200 B.n425 B.n52 585
R201 B.n424 B.n423 585
R202 B.n422 B.n53 585
R203 B.n421 B.n420 585
R204 B.n419 B.n54 585
R205 B.n418 B.n417 585
R206 B.n416 B.n55 585
R207 B.n415 B.n414 585
R208 B.n413 B.n56 585
R209 B.n412 B.n411 585
R210 B.n410 B.n57 585
R211 B.n409 B.n408 585
R212 B.n407 B.n58 585
R213 B.n406 B.n405 585
R214 B.n404 B.n59 585
R215 B.n403 B.n402 585
R216 B.n520 B.n519 585
R217 B.n521 B.n16 585
R218 B.n523 B.n522 585
R219 B.n524 B.n15 585
R220 B.n526 B.n525 585
R221 B.n527 B.n14 585
R222 B.n529 B.n528 585
R223 B.n530 B.n13 585
R224 B.n532 B.n531 585
R225 B.n533 B.n12 585
R226 B.n535 B.n534 585
R227 B.n536 B.n11 585
R228 B.n538 B.n537 585
R229 B.n539 B.n10 585
R230 B.n541 B.n540 585
R231 B.n542 B.n9 585
R232 B.n544 B.n543 585
R233 B.n545 B.n8 585
R234 B.n547 B.n546 585
R235 B.n548 B.n7 585
R236 B.n550 B.n549 585
R237 B.n551 B.n6 585
R238 B.n553 B.n552 585
R239 B.n554 B.n5 585
R240 B.n556 B.n555 585
R241 B.n557 B.n4 585
R242 B.n559 B.n558 585
R243 B.n560 B.n3 585
R244 B.n562 B.n561 585
R245 B.n563 B.n0 585
R246 B.n2 B.n1 585
R247 B.n149 B.n148 585
R248 B.n151 B.n150 585
R249 B.n152 B.n147 585
R250 B.n154 B.n153 585
R251 B.n155 B.n146 585
R252 B.n157 B.n156 585
R253 B.n158 B.n145 585
R254 B.n160 B.n159 585
R255 B.n161 B.n144 585
R256 B.n163 B.n162 585
R257 B.n164 B.n143 585
R258 B.n166 B.n165 585
R259 B.n167 B.n142 585
R260 B.n169 B.n168 585
R261 B.n170 B.n141 585
R262 B.n172 B.n171 585
R263 B.n173 B.n140 585
R264 B.n175 B.n174 585
R265 B.n176 B.n139 585
R266 B.n178 B.n177 585
R267 B.n179 B.n138 585
R268 B.n181 B.n180 585
R269 B.n182 B.n137 585
R270 B.n184 B.n183 585
R271 B.n185 B.n136 585
R272 B.n187 B.n186 585
R273 B.n188 B.n135 585
R274 B.n190 B.n189 585
R275 B.n191 B.n134 585
R276 B.n192 B.n191 516.524
R277 B.n310 B.n91 516.524
R278 B.n402 B.n401 516.524
R279 B.n520 B.n17 516.524
R280 B.n108 B.t1 400.846
R281 B.n42 B.t11 400.846
R282 B.n116 B.t4 400.846
R283 B.n34 B.t8 400.846
R284 B.n109 B.t2 326.178
R285 B.n43 B.t10 326.178
R286 B.n117 B.t5 326.178
R287 B.n35 B.t7 326.178
R288 B.n116 B.t3 272.512
R289 B.n108 B.t0 272.512
R290 B.n42 B.t9 272.512
R291 B.n34 B.t6 272.512
R292 B.n565 B.n564 256.663
R293 B.n564 B.n563 235.042
R294 B.n564 B.n2 235.042
R295 B.n192 B.n133 163.367
R296 B.n196 B.n133 163.367
R297 B.n197 B.n196 163.367
R298 B.n198 B.n197 163.367
R299 B.n198 B.n131 163.367
R300 B.n202 B.n131 163.367
R301 B.n203 B.n202 163.367
R302 B.n204 B.n203 163.367
R303 B.n204 B.n129 163.367
R304 B.n208 B.n129 163.367
R305 B.n209 B.n208 163.367
R306 B.n210 B.n209 163.367
R307 B.n210 B.n127 163.367
R308 B.n214 B.n127 163.367
R309 B.n215 B.n214 163.367
R310 B.n216 B.n215 163.367
R311 B.n216 B.n125 163.367
R312 B.n220 B.n125 163.367
R313 B.n221 B.n220 163.367
R314 B.n222 B.n221 163.367
R315 B.n222 B.n123 163.367
R316 B.n226 B.n123 163.367
R317 B.n227 B.n226 163.367
R318 B.n228 B.n227 163.367
R319 B.n228 B.n121 163.367
R320 B.n232 B.n121 163.367
R321 B.n233 B.n232 163.367
R322 B.n234 B.n233 163.367
R323 B.n234 B.n119 163.367
R324 B.n238 B.n119 163.367
R325 B.n239 B.n238 163.367
R326 B.n240 B.n239 163.367
R327 B.n240 B.n115 163.367
R328 B.n245 B.n115 163.367
R329 B.n246 B.n245 163.367
R330 B.n247 B.n246 163.367
R331 B.n247 B.n113 163.367
R332 B.n251 B.n113 163.367
R333 B.n252 B.n251 163.367
R334 B.n253 B.n252 163.367
R335 B.n253 B.n111 163.367
R336 B.n257 B.n111 163.367
R337 B.n258 B.n257 163.367
R338 B.n258 B.n107 163.367
R339 B.n262 B.n107 163.367
R340 B.n263 B.n262 163.367
R341 B.n264 B.n263 163.367
R342 B.n264 B.n105 163.367
R343 B.n268 B.n105 163.367
R344 B.n269 B.n268 163.367
R345 B.n270 B.n269 163.367
R346 B.n270 B.n103 163.367
R347 B.n274 B.n103 163.367
R348 B.n275 B.n274 163.367
R349 B.n276 B.n275 163.367
R350 B.n276 B.n101 163.367
R351 B.n280 B.n101 163.367
R352 B.n281 B.n280 163.367
R353 B.n282 B.n281 163.367
R354 B.n282 B.n99 163.367
R355 B.n286 B.n99 163.367
R356 B.n287 B.n286 163.367
R357 B.n288 B.n287 163.367
R358 B.n288 B.n97 163.367
R359 B.n292 B.n97 163.367
R360 B.n293 B.n292 163.367
R361 B.n294 B.n293 163.367
R362 B.n294 B.n95 163.367
R363 B.n298 B.n95 163.367
R364 B.n299 B.n298 163.367
R365 B.n300 B.n299 163.367
R366 B.n300 B.n93 163.367
R367 B.n304 B.n93 163.367
R368 B.n305 B.n304 163.367
R369 B.n306 B.n305 163.367
R370 B.n306 B.n91 163.367
R371 B.n401 B.n400 163.367
R372 B.n400 B.n61 163.367
R373 B.n396 B.n61 163.367
R374 B.n396 B.n395 163.367
R375 B.n395 B.n394 163.367
R376 B.n394 B.n63 163.367
R377 B.n390 B.n63 163.367
R378 B.n390 B.n389 163.367
R379 B.n389 B.n388 163.367
R380 B.n388 B.n65 163.367
R381 B.n384 B.n65 163.367
R382 B.n384 B.n383 163.367
R383 B.n383 B.n382 163.367
R384 B.n382 B.n67 163.367
R385 B.n378 B.n67 163.367
R386 B.n378 B.n377 163.367
R387 B.n377 B.n376 163.367
R388 B.n376 B.n69 163.367
R389 B.n372 B.n69 163.367
R390 B.n372 B.n371 163.367
R391 B.n371 B.n370 163.367
R392 B.n370 B.n71 163.367
R393 B.n366 B.n71 163.367
R394 B.n366 B.n365 163.367
R395 B.n365 B.n364 163.367
R396 B.n364 B.n73 163.367
R397 B.n360 B.n73 163.367
R398 B.n360 B.n359 163.367
R399 B.n359 B.n358 163.367
R400 B.n358 B.n75 163.367
R401 B.n354 B.n75 163.367
R402 B.n354 B.n353 163.367
R403 B.n353 B.n352 163.367
R404 B.n352 B.n77 163.367
R405 B.n348 B.n77 163.367
R406 B.n348 B.n347 163.367
R407 B.n347 B.n346 163.367
R408 B.n346 B.n79 163.367
R409 B.n342 B.n79 163.367
R410 B.n342 B.n341 163.367
R411 B.n341 B.n340 163.367
R412 B.n340 B.n81 163.367
R413 B.n336 B.n81 163.367
R414 B.n336 B.n335 163.367
R415 B.n335 B.n334 163.367
R416 B.n334 B.n83 163.367
R417 B.n330 B.n83 163.367
R418 B.n330 B.n329 163.367
R419 B.n329 B.n328 163.367
R420 B.n328 B.n85 163.367
R421 B.n324 B.n85 163.367
R422 B.n324 B.n323 163.367
R423 B.n323 B.n322 163.367
R424 B.n322 B.n87 163.367
R425 B.n318 B.n87 163.367
R426 B.n318 B.n317 163.367
R427 B.n317 B.n316 163.367
R428 B.n316 B.n89 163.367
R429 B.n312 B.n89 163.367
R430 B.n312 B.n311 163.367
R431 B.n311 B.n310 163.367
R432 B.n516 B.n17 163.367
R433 B.n516 B.n515 163.367
R434 B.n515 B.n514 163.367
R435 B.n514 B.n19 163.367
R436 B.n510 B.n19 163.367
R437 B.n510 B.n509 163.367
R438 B.n509 B.n508 163.367
R439 B.n508 B.n21 163.367
R440 B.n504 B.n21 163.367
R441 B.n504 B.n503 163.367
R442 B.n503 B.n502 163.367
R443 B.n502 B.n23 163.367
R444 B.n498 B.n23 163.367
R445 B.n498 B.n497 163.367
R446 B.n497 B.n496 163.367
R447 B.n496 B.n25 163.367
R448 B.n492 B.n25 163.367
R449 B.n492 B.n491 163.367
R450 B.n491 B.n490 163.367
R451 B.n490 B.n27 163.367
R452 B.n486 B.n27 163.367
R453 B.n486 B.n485 163.367
R454 B.n485 B.n484 163.367
R455 B.n484 B.n29 163.367
R456 B.n480 B.n29 163.367
R457 B.n480 B.n479 163.367
R458 B.n479 B.n478 163.367
R459 B.n478 B.n31 163.367
R460 B.n474 B.n31 163.367
R461 B.n474 B.n473 163.367
R462 B.n473 B.n472 163.367
R463 B.n472 B.n33 163.367
R464 B.n468 B.n33 163.367
R465 B.n468 B.n467 163.367
R466 B.n467 B.n37 163.367
R467 B.n463 B.n37 163.367
R468 B.n463 B.n462 163.367
R469 B.n462 B.n461 163.367
R470 B.n461 B.n39 163.367
R471 B.n457 B.n39 163.367
R472 B.n457 B.n456 163.367
R473 B.n456 B.n455 163.367
R474 B.n455 B.n41 163.367
R475 B.n450 B.n41 163.367
R476 B.n450 B.n449 163.367
R477 B.n449 B.n448 163.367
R478 B.n448 B.n45 163.367
R479 B.n444 B.n45 163.367
R480 B.n444 B.n443 163.367
R481 B.n443 B.n442 163.367
R482 B.n442 B.n47 163.367
R483 B.n438 B.n47 163.367
R484 B.n438 B.n437 163.367
R485 B.n437 B.n436 163.367
R486 B.n436 B.n49 163.367
R487 B.n432 B.n49 163.367
R488 B.n432 B.n431 163.367
R489 B.n431 B.n430 163.367
R490 B.n430 B.n51 163.367
R491 B.n426 B.n51 163.367
R492 B.n426 B.n425 163.367
R493 B.n425 B.n424 163.367
R494 B.n424 B.n53 163.367
R495 B.n420 B.n53 163.367
R496 B.n420 B.n419 163.367
R497 B.n419 B.n418 163.367
R498 B.n418 B.n55 163.367
R499 B.n414 B.n55 163.367
R500 B.n414 B.n413 163.367
R501 B.n413 B.n412 163.367
R502 B.n412 B.n57 163.367
R503 B.n408 B.n57 163.367
R504 B.n408 B.n407 163.367
R505 B.n407 B.n406 163.367
R506 B.n406 B.n59 163.367
R507 B.n402 B.n59 163.367
R508 B.n521 B.n520 163.367
R509 B.n522 B.n521 163.367
R510 B.n522 B.n15 163.367
R511 B.n526 B.n15 163.367
R512 B.n527 B.n526 163.367
R513 B.n528 B.n527 163.367
R514 B.n528 B.n13 163.367
R515 B.n532 B.n13 163.367
R516 B.n533 B.n532 163.367
R517 B.n534 B.n533 163.367
R518 B.n534 B.n11 163.367
R519 B.n538 B.n11 163.367
R520 B.n539 B.n538 163.367
R521 B.n540 B.n539 163.367
R522 B.n540 B.n9 163.367
R523 B.n544 B.n9 163.367
R524 B.n545 B.n544 163.367
R525 B.n546 B.n545 163.367
R526 B.n546 B.n7 163.367
R527 B.n550 B.n7 163.367
R528 B.n551 B.n550 163.367
R529 B.n552 B.n551 163.367
R530 B.n552 B.n5 163.367
R531 B.n556 B.n5 163.367
R532 B.n557 B.n556 163.367
R533 B.n558 B.n557 163.367
R534 B.n558 B.n3 163.367
R535 B.n562 B.n3 163.367
R536 B.n563 B.n562 163.367
R537 B.n149 B.n2 163.367
R538 B.n150 B.n149 163.367
R539 B.n150 B.n147 163.367
R540 B.n154 B.n147 163.367
R541 B.n155 B.n154 163.367
R542 B.n156 B.n155 163.367
R543 B.n156 B.n145 163.367
R544 B.n160 B.n145 163.367
R545 B.n161 B.n160 163.367
R546 B.n162 B.n161 163.367
R547 B.n162 B.n143 163.367
R548 B.n166 B.n143 163.367
R549 B.n167 B.n166 163.367
R550 B.n168 B.n167 163.367
R551 B.n168 B.n141 163.367
R552 B.n172 B.n141 163.367
R553 B.n173 B.n172 163.367
R554 B.n174 B.n173 163.367
R555 B.n174 B.n139 163.367
R556 B.n178 B.n139 163.367
R557 B.n179 B.n178 163.367
R558 B.n180 B.n179 163.367
R559 B.n180 B.n137 163.367
R560 B.n184 B.n137 163.367
R561 B.n185 B.n184 163.367
R562 B.n186 B.n185 163.367
R563 B.n186 B.n135 163.367
R564 B.n190 B.n135 163.367
R565 B.n191 B.n190 163.367
R566 B.n117 B.n116 74.6672
R567 B.n109 B.n108 74.6672
R568 B.n43 B.n42 74.6672
R569 B.n35 B.n34 74.6672
R570 B.n243 B.n117 59.5399
R571 B.n110 B.n109 59.5399
R572 B.n453 B.n43 59.5399
R573 B.n36 B.n35 59.5399
R574 B.n519 B.n518 33.5615
R575 B.n403 B.n60 33.5615
R576 B.n309 B.n308 33.5615
R577 B.n193 B.n134 33.5615
R578 B B.n565 18.0485
R579 B.n519 B.n16 10.6151
R580 B.n523 B.n16 10.6151
R581 B.n524 B.n523 10.6151
R582 B.n525 B.n524 10.6151
R583 B.n525 B.n14 10.6151
R584 B.n529 B.n14 10.6151
R585 B.n530 B.n529 10.6151
R586 B.n531 B.n530 10.6151
R587 B.n531 B.n12 10.6151
R588 B.n535 B.n12 10.6151
R589 B.n536 B.n535 10.6151
R590 B.n537 B.n536 10.6151
R591 B.n537 B.n10 10.6151
R592 B.n541 B.n10 10.6151
R593 B.n542 B.n541 10.6151
R594 B.n543 B.n542 10.6151
R595 B.n543 B.n8 10.6151
R596 B.n547 B.n8 10.6151
R597 B.n548 B.n547 10.6151
R598 B.n549 B.n548 10.6151
R599 B.n549 B.n6 10.6151
R600 B.n553 B.n6 10.6151
R601 B.n554 B.n553 10.6151
R602 B.n555 B.n554 10.6151
R603 B.n555 B.n4 10.6151
R604 B.n559 B.n4 10.6151
R605 B.n560 B.n559 10.6151
R606 B.n561 B.n560 10.6151
R607 B.n561 B.n0 10.6151
R608 B.n518 B.n517 10.6151
R609 B.n517 B.n18 10.6151
R610 B.n513 B.n18 10.6151
R611 B.n513 B.n512 10.6151
R612 B.n512 B.n511 10.6151
R613 B.n511 B.n20 10.6151
R614 B.n507 B.n20 10.6151
R615 B.n507 B.n506 10.6151
R616 B.n506 B.n505 10.6151
R617 B.n505 B.n22 10.6151
R618 B.n501 B.n22 10.6151
R619 B.n501 B.n500 10.6151
R620 B.n500 B.n499 10.6151
R621 B.n499 B.n24 10.6151
R622 B.n495 B.n24 10.6151
R623 B.n495 B.n494 10.6151
R624 B.n494 B.n493 10.6151
R625 B.n493 B.n26 10.6151
R626 B.n489 B.n26 10.6151
R627 B.n489 B.n488 10.6151
R628 B.n488 B.n487 10.6151
R629 B.n487 B.n28 10.6151
R630 B.n483 B.n28 10.6151
R631 B.n483 B.n482 10.6151
R632 B.n482 B.n481 10.6151
R633 B.n481 B.n30 10.6151
R634 B.n477 B.n30 10.6151
R635 B.n477 B.n476 10.6151
R636 B.n476 B.n475 10.6151
R637 B.n475 B.n32 10.6151
R638 B.n471 B.n32 10.6151
R639 B.n471 B.n470 10.6151
R640 B.n470 B.n469 10.6151
R641 B.n466 B.n465 10.6151
R642 B.n465 B.n464 10.6151
R643 B.n464 B.n38 10.6151
R644 B.n460 B.n38 10.6151
R645 B.n460 B.n459 10.6151
R646 B.n459 B.n458 10.6151
R647 B.n458 B.n40 10.6151
R648 B.n454 B.n40 10.6151
R649 B.n452 B.n451 10.6151
R650 B.n451 B.n44 10.6151
R651 B.n447 B.n44 10.6151
R652 B.n447 B.n446 10.6151
R653 B.n446 B.n445 10.6151
R654 B.n445 B.n46 10.6151
R655 B.n441 B.n46 10.6151
R656 B.n441 B.n440 10.6151
R657 B.n440 B.n439 10.6151
R658 B.n439 B.n48 10.6151
R659 B.n435 B.n48 10.6151
R660 B.n435 B.n434 10.6151
R661 B.n434 B.n433 10.6151
R662 B.n433 B.n50 10.6151
R663 B.n429 B.n50 10.6151
R664 B.n429 B.n428 10.6151
R665 B.n428 B.n427 10.6151
R666 B.n427 B.n52 10.6151
R667 B.n423 B.n52 10.6151
R668 B.n423 B.n422 10.6151
R669 B.n422 B.n421 10.6151
R670 B.n421 B.n54 10.6151
R671 B.n417 B.n54 10.6151
R672 B.n417 B.n416 10.6151
R673 B.n416 B.n415 10.6151
R674 B.n415 B.n56 10.6151
R675 B.n411 B.n56 10.6151
R676 B.n411 B.n410 10.6151
R677 B.n410 B.n409 10.6151
R678 B.n409 B.n58 10.6151
R679 B.n405 B.n58 10.6151
R680 B.n405 B.n404 10.6151
R681 B.n404 B.n403 10.6151
R682 B.n399 B.n60 10.6151
R683 B.n399 B.n398 10.6151
R684 B.n398 B.n397 10.6151
R685 B.n397 B.n62 10.6151
R686 B.n393 B.n62 10.6151
R687 B.n393 B.n392 10.6151
R688 B.n392 B.n391 10.6151
R689 B.n391 B.n64 10.6151
R690 B.n387 B.n64 10.6151
R691 B.n387 B.n386 10.6151
R692 B.n386 B.n385 10.6151
R693 B.n385 B.n66 10.6151
R694 B.n381 B.n66 10.6151
R695 B.n381 B.n380 10.6151
R696 B.n380 B.n379 10.6151
R697 B.n379 B.n68 10.6151
R698 B.n375 B.n68 10.6151
R699 B.n375 B.n374 10.6151
R700 B.n374 B.n373 10.6151
R701 B.n373 B.n70 10.6151
R702 B.n369 B.n70 10.6151
R703 B.n369 B.n368 10.6151
R704 B.n368 B.n367 10.6151
R705 B.n367 B.n72 10.6151
R706 B.n363 B.n72 10.6151
R707 B.n363 B.n362 10.6151
R708 B.n362 B.n361 10.6151
R709 B.n361 B.n74 10.6151
R710 B.n357 B.n74 10.6151
R711 B.n357 B.n356 10.6151
R712 B.n356 B.n355 10.6151
R713 B.n355 B.n76 10.6151
R714 B.n351 B.n76 10.6151
R715 B.n351 B.n350 10.6151
R716 B.n350 B.n349 10.6151
R717 B.n349 B.n78 10.6151
R718 B.n345 B.n78 10.6151
R719 B.n345 B.n344 10.6151
R720 B.n344 B.n343 10.6151
R721 B.n343 B.n80 10.6151
R722 B.n339 B.n80 10.6151
R723 B.n339 B.n338 10.6151
R724 B.n338 B.n337 10.6151
R725 B.n337 B.n82 10.6151
R726 B.n333 B.n82 10.6151
R727 B.n333 B.n332 10.6151
R728 B.n332 B.n331 10.6151
R729 B.n331 B.n84 10.6151
R730 B.n327 B.n84 10.6151
R731 B.n327 B.n326 10.6151
R732 B.n326 B.n325 10.6151
R733 B.n325 B.n86 10.6151
R734 B.n321 B.n86 10.6151
R735 B.n321 B.n320 10.6151
R736 B.n320 B.n319 10.6151
R737 B.n319 B.n88 10.6151
R738 B.n315 B.n88 10.6151
R739 B.n315 B.n314 10.6151
R740 B.n314 B.n313 10.6151
R741 B.n313 B.n90 10.6151
R742 B.n309 B.n90 10.6151
R743 B.n148 B.n1 10.6151
R744 B.n151 B.n148 10.6151
R745 B.n152 B.n151 10.6151
R746 B.n153 B.n152 10.6151
R747 B.n153 B.n146 10.6151
R748 B.n157 B.n146 10.6151
R749 B.n158 B.n157 10.6151
R750 B.n159 B.n158 10.6151
R751 B.n159 B.n144 10.6151
R752 B.n163 B.n144 10.6151
R753 B.n164 B.n163 10.6151
R754 B.n165 B.n164 10.6151
R755 B.n165 B.n142 10.6151
R756 B.n169 B.n142 10.6151
R757 B.n170 B.n169 10.6151
R758 B.n171 B.n170 10.6151
R759 B.n171 B.n140 10.6151
R760 B.n175 B.n140 10.6151
R761 B.n176 B.n175 10.6151
R762 B.n177 B.n176 10.6151
R763 B.n177 B.n138 10.6151
R764 B.n181 B.n138 10.6151
R765 B.n182 B.n181 10.6151
R766 B.n183 B.n182 10.6151
R767 B.n183 B.n136 10.6151
R768 B.n187 B.n136 10.6151
R769 B.n188 B.n187 10.6151
R770 B.n189 B.n188 10.6151
R771 B.n189 B.n134 10.6151
R772 B.n194 B.n193 10.6151
R773 B.n195 B.n194 10.6151
R774 B.n195 B.n132 10.6151
R775 B.n199 B.n132 10.6151
R776 B.n200 B.n199 10.6151
R777 B.n201 B.n200 10.6151
R778 B.n201 B.n130 10.6151
R779 B.n205 B.n130 10.6151
R780 B.n206 B.n205 10.6151
R781 B.n207 B.n206 10.6151
R782 B.n207 B.n128 10.6151
R783 B.n211 B.n128 10.6151
R784 B.n212 B.n211 10.6151
R785 B.n213 B.n212 10.6151
R786 B.n213 B.n126 10.6151
R787 B.n217 B.n126 10.6151
R788 B.n218 B.n217 10.6151
R789 B.n219 B.n218 10.6151
R790 B.n219 B.n124 10.6151
R791 B.n223 B.n124 10.6151
R792 B.n224 B.n223 10.6151
R793 B.n225 B.n224 10.6151
R794 B.n225 B.n122 10.6151
R795 B.n229 B.n122 10.6151
R796 B.n230 B.n229 10.6151
R797 B.n231 B.n230 10.6151
R798 B.n231 B.n120 10.6151
R799 B.n235 B.n120 10.6151
R800 B.n236 B.n235 10.6151
R801 B.n237 B.n236 10.6151
R802 B.n237 B.n118 10.6151
R803 B.n241 B.n118 10.6151
R804 B.n242 B.n241 10.6151
R805 B.n244 B.n114 10.6151
R806 B.n248 B.n114 10.6151
R807 B.n249 B.n248 10.6151
R808 B.n250 B.n249 10.6151
R809 B.n250 B.n112 10.6151
R810 B.n254 B.n112 10.6151
R811 B.n255 B.n254 10.6151
R812 B.n256 B.n255 10.6151
R813 B.n260 B.n259 10.6151
R814 B.n261 B.n260 10.6151
R815 B.n261 B.n106 10.6151
R816 B.n265 B.n106 10.6151
R817 B.n266 B.n265 10.6151
R818 B.n267 B.n266 10.6151
R819 B.n267 B.n104 10.6151
R820 B.n271 B.n104 10.6151
R821 B.n272 B.n271 10.6151
R822 B.n273 B.n272 10.6151
R823 B.n273 B.n102 10.6151
R824 B.n277 B.n102 10.6151
R825 B.n278 B.n277 10.6151
R826 B.n279 B.n278 10.6151
R827 B.n279 B.n100 10.6151
R828 B.n283 B.n100 10.6151
R829 B.n284 B.n283 10.6151
R830 B.n285 B.n284 10.6151
R831 B.n285 B.n98 10.6151
R832 B.n289 B.n98 10.6151
R833 B.n290 B.n289 10.6151
R834 B.n291 B.n290 10.6151
R835 B.n291 B.n96 10.6151
R836 B.n295 B.n96 10.6151
R837 B.n296 B.n295 10.6151
R838 B.n297 B.n296 10.6151
R839 B.n297 B.n94 10.6151
R840 B.n301 B.n94 10.6151
R841 B.n302 B.n301 10.6151
R842 B.n303 B.n302 10.6151
R843 B.n303 B.n92 10.6151
R844 B.n307 B.n92 10.6151
R845 B.n308 B.n307 10.6151
R846 B.n565 B.n0 8.11757
R847 B.n565 B.n1 8.11757
R848 B.n466 B.n36 6.5566
R849 B.n454 B.n453 6.5566
R850 B.n244 B.n243 6.5566
R851 B.n256 B.n110 6.5566
R852 B.n469 B.n36 4.05904
R853 B.n453 B.n452 4.05904
R854 B.n243 B.n242 4.05904
R855 B.n259 B.n110 4.05904
R856 VN VN.t0 147.173
R857 VN VN.t1 102.772
R858 VTAIL.n194 VTAIL.n150 756.745
R859 VTAIL.n44 VTAIL.n0 756.745
R860 VTAIL.n144 VTAIL.n100 756.745
R861 VTAIL.n94 VTAIL.n50 756.745
R862 VTAIL.n167 VTAIL.n166 585
R863 VTAIL.n169 VTAIL.n168 585
R864 VTAIL.n162 VTAIL.n161 585
R865 VTAIL.n175 VTAIL.n174 585
R866 VTAIL.n177 VTAIL.n176 585
R867 VTAIL.n158 VTAIL.n157 585
R868 VTAIL.n184 VTAIL.n183 585
R869 VTAIL.n185 VTAIL.n156 585
R870 VTAIL.n187 VTAIL.n186 585
R871 VTAIL.n154 VTAIL.n153 585
R872 VTAIL.n193 VTAIL.n192 585
R873 VTAIL.n195 VTAIL.n194 585
R874 VTAIL.n17 VTAIL.n16 585
R875 VTAIL.n19 VTAIL.n18 585
R876 VTAIL.n12 VTAIL.n11 585
R877 VTAIL.n25 VTAIL.n24 585
R878 VTAIL.n27 VTAIL.n26 585
R879 VTAIL.n8 VTAIL.n7 585
R880 VTAIL.n34 VTAIL.n33 585
R881 VTAIL.n35 VTAIL.n6 585
R882 VTAIL.n37 VTAIL.n36 585
R883 VTAIL.n4 VTAIL.n3 585
R884 VTAIL.n43 VTAIL.n42 585
R885 VTAIL.n45 VTAIL.n44 585
R886 VTAIL.n145 VTAIL.n144 585
R887 VTAIL.n143 VTAIL.n142 585
R888 VTAIL.n104 VTAIL.n103 585
R889 VTAIL.n108 VTAIL.n106 585
R890 VTAIL.n137 VTAIL.n136 585
R891 VTAIL.n135 VTAIL.n134 585
R892 VTAIL.n110 VTAIL.n109 585
R893 VTAIL.n129 VTAIL.n128 585
R894 VTAIL.n127 VTAIL.n126 585
R895 VTAIL.n114 VTAIL.n113 585
R896 VTAIL.n121 VTAIL.n120 585
R897 VTAIL.n119 VTAIL.n118 585
R898 VTAIL.n95 VTAIL.n94 585
R899 VTAIL.n93 VTAIL.n92 585
R900 VTAIL.n54 VTAIL.n53 585
R901 VTAIL.n58 VTAIL.n56 585
R902 VTAIL.n87 VTAIL.n86 585
R903 VTAIL.n85 VTAIL.n84 585
R904 VTAIL.n60 VTAIL.n59 585
R905 VTAIL.n79 VTAIL.n78 585
R906 VTAIL.n77 VTAIL.n76 585
R907 VTAIL.n64 VTAIL.n63 585
R908 VTAIL.n71 VTAIL.n70 585
R909 VTAIL.n69 VTAIL.n68 585
R910 VTAIL.n165 VTAIL.t2 329.038
R911 VTAIL.n15 VTAIL.t0 329.038
R912 VTAIL.n117 VTAIL.t1 329.038
R913 VTAIL.n67 VTAIL.t3 329.038
R914 VTAIL.n168 VTAIL.n167 171.744
R915 VTAIL.n168 VTAIL.n161 171.744
R916 VTAIL.n175 VTAIL.n161 171.744
R917 VTAIL.n176 VTAIL.n175 171.744
R918 VTAIL.n176 VTAIL.n157 171.744
R919 VTAIL.n184 VTAIL.n157 171.744
R920 VTAIL.n185 VTAIL.n184 171.744
R921 VTAIL.n186 VTAIL.n185 171.744
R922 VTAIL.n186 VTAIL.n153 171.744
R923 VTAIL.n193 VTAIL.n153 171.744
R924 VTAIL.n194 VTAIL.n193 171.744
R925 VTAIL.n18 VTAIL.n17 171.744
R926 VTAIL.n18 VTAIL.n11 171.744
R927 VTAIL.n25 VTAIL.n11 171.744
R928 VTAIL.n26 VTAIL.n25 171.744
R929 VTAIL.n26 VTAIL.n7 171.744
R930 VTAIL.n34 VTAIL.n7 171.744
R931 VTAIL.n35 VTAIL.n34 171.744
R932 VTAIL.n36 VTAIL.n35 171.744
R933 VTAIL.n36 VTAIL.n3 171.744
R934 VTAIL.n43 VTAIL.n3 171.744
R935 VTAIL.n44 VTAIL.n43 171.744
R936 VTAIL.n144 VTAIL.n143 171.744
R937 VTAIL.n143 VTAIL.n103 171.744
R938 VTAIL.n108 VTAIL.n103 171.744
R939 VTAIL.n136 VTAIL.n108 171.744
R940 VTAIL.n136 VTAIL.n135 171.744
R941 VTAIL.n135 VTAIL.n109 171.744
R942 VTAIL.n128 VTAIL.n109 171.744
R943 VTAIL.n128 VTAIL.n127 171.744
R944 VTAIL.n127 VTAIL.n113 171.744
R945 VTAIL.n120 VTAIL.n113 171.744
R946 VTAIL.n120 VTAIL.n119 171.744
R947 VTAIL.n94 VTAIL.n93 171.744
R948 VTAIL.n93 VTAIL.n53 171.744
R949 VTAIL.n58 VTAIL.n53 171.744
R950 VTAIL.n86 VTAIL.n58 171.744
R951 VTAIL.n86 VTAIL.n85 171.744
R952 VTAIL.n85 VTAIL.n59 171.744
R953 VTAIL.n78 VTAIL.n59 171.744
R954 VTAIL.n78 VTAIL.n77 171.744
R955 VTAIL.n77 VTAIL.n63 171.744
R956 VTAIL.n70 VTAIL.n63 171.744
R957 VTAIL.n70 VTAIL.n69 171.744
R958 VTAIL.n167 VTAIL.t2 85.8723
R959 VTAIL.n17 VTAIL.t0 85.8723
R960 VTAIL.n119 VTAIL.t1 85.8723
R961 VTAIL.n69 VTAIL.t3 85.8723
R962 VTAIL.n199 VTAIL.n198 32.5732
R963 VTAIL.n49 VTAIL.n48 32.5732
R964 VTAIL.n149 VTAIL.n148 32.5732
R965 VTAIL.n99 VTAIL.n98 32.5732
R966 VTAIL.n99 VTAIL.n49 26.9876
R967 VTAIL.n199 VTAIL.n149 23.6686
R968 VTAIL.n187 VTAIL.n154 13.1884
R969 VTAIL.n37 VTAIL.n4 13.1884
R970 VTAIL.n106 VTAIL.n104 13.1884
R971 VTAIL.n56 VTAIL.n54 13.1884
R972 VTAIL.n188 VTAIL.n156 12.8005
R973 VTAIL.n192 VTAIL.n191 12.8005
R974 VTAIL.n38 VTAIL.n6 12.8005
R975 VTAIL.n42 VTAIL.n41 12.8005
R976 VTAIL.n142 VTAIL.n141 12.8005
R977 VTAIL.n138 VTAIL.n137 12.8005
R978 VTAIL.n92 VTAIL.n91 12.8005
R979 VTAIL.n88 VTAIL.n87 12.8005
R980 VTAIL.n183 VTAIL.n182 12.0247
R981 VTAIL.n195 VTAIL.n152 12.0247
R982 VTAIL.n33 VTAIL.n32 12.0247
R983 VTAIL.n45 VTAIL.n2 12.0247
R984 VTAIL.n145 VTAIL.n102 12.0247
R985 VTAIL.n134 VTAIL.n107 12.0247
R986 VTAIL.n95 VTAIL.n52 12.0247
R987 VTAIL.n84 VTAIL.n57 12.0247
R988 VTAIL.n181 VTAIL.n158 11.249
R989 VTAIL.n196 VTAIL.n150 11.249
R990 VTAIL.n31 VTAIL.n8 11.249
R991 VTAIL.n46 VTAIL.n0 11.249
R992 VTAIL.n146 VTAIL.n100 11.249
R993 VTAIL.n133 VTAIL.n110 11.249
R994 VTAIL.n96 VTAIL.n50 11.249
R995 VTAIL.n83 VTAIL.n60 11.249
R996 VTAIL.n166 VTAIL.n165 10.7239
R997 VTAIL.n16 VTAIL.n15 10.7239
R998 VTAIL.n118 VTAIL.n117 10.7239
R999 VTAIL.n68 VTAIL.n67 10.7239
R1000 VTAIL.n178 VTAIL.n177 10.4732
R1001 VTAIL.n28 VTAIL.n27 10.4732
R1002 VTAIL.n130 VTAIL.n129 10.4732
R1003 VTAIL.n80 VTAIL.n79 10.4732
R1004 VTAIL.n174 VTAIL.n160 9.69747
R1005 VTAIL.n24 VTAIL.n10 9.69747
R1006 VTAIL.n126 VTAIL.n112 9.69747
R1007 VTAIL.n76 VTAIL.n62 9.69747
R1008 VTAIL.n198 VTAIL.n197 9.45567
R1009 VTAIL.n48 VTAIL.n47 9.45567
R1010 VTAIL.n148 VTAIL.n147 9.45567
R1011 VTAIL.n98 VTAIL.n97 9.45567
R1012 VTAIL.n197 VTAIL.n196 9.3005
R1013 VTAIL.n152 VTAIL.n151 9.3005
R1014 VTAIL.n191 VTAIL.n190 9.3005
R1015 VTAIL.n164 VTAIL.n163 9.3005
R1016 VTAIL.n171 VTAIL.n170 9.3005
R1017 VTAIL.n173 VTAIL.n172 9.3005
R1018 VTAIL.n160 VTAIL.n159 9.3005
R1019 VTAIL.n179 VTAIL.n178 9.3005
R1020 VTAIL.n181 VTAIL.n180 9.3005
R1021 VTAIL.n182 VTAIL.n155 9.3005
R1022 VTAIL.n189 VTAIL.n188 9.3005
R1023 VTAIL.n47 VTAIL.n46 9.3005
R1024 VTAIL.n2 VTAIL.n1 9.3005
R1025 VTAIL.n41 VTAIL.n40 9.3005
R1026 VTAIL.n14 VTAIL.n13 9.3005
R1027 VTAIL.n21 VTAIL.n20 9.3005
R1028 VTAIL.n23 VTAIL.n22 9.3005
R1029 VTAIL.n10 VTAIL.n9 9.3005
R1030 VTAIL.n29 VTAIL.n28 9.3005
R1031 VTAIL.n31 VTAIL.n30 9.3005
R1032 VTAIL.n32 VTAIL.n5 9.3005
R1033 VTAIL.n39 VTAIL.n38 9.3005
R1034 VTAIL.n116 VTAIL.n115 9.3005
R1035 VTAIL.n123 VTAIL.n122 9.3005
R1036 VTAIL.n125 VTAIL.n124 9.3005
R1037 VTAIL.n112 VTAIL.n111 9.3005
R1038 VTAIL.n131 VTAIL.n130 9.3005
R1039 VTAIL.n133 VTAIL.n132 9.3005
R1040 VTAIL.n107 VTAIL.n105 9.3005
R1041 VTAIL.n139 VTAIL.n138 9.3005
R1042 VTAIL.n147 VTAIL.n146 9.3005
R1043 VTAIL.n102 VTAIL.n101 9.3005
R1044 VTAIL.n141 VTAIL.n140 9.3005
R1045 VTAIL.n66 VTAIL.n65 9.3005
R1046 VTAIL.n73 VTAIL.n72 9.3005
R1047 VTAIL.n75 VTAIL.n74 9.3005
R1048 VTAIL.n62 VTAIL.n61 9.3005
R1049 VTAIL.n81 VTAIL.n80 9.3005
R1050 VTAIL.n83 VTAIL.n82 9.3005
R1051 VTAIL.n57 VTAIL.n55 9.3005
R1052 VTAIL.n89 VTAIL.n88 9.3005
R1053 VTAIL.n97 VTAIL.n96 9.3005
R1054 VTAIL.n52 VTAIL.n51 9.3005
R1055 VTAIL.n91 VTAIL.n90 9.3005
R1056 VTAIL.n173 VTAIL.n162 8.92171
R1057 VTAIL.n23 VTAIL.n12 8.92171
R1058 VTAIL.n125 VTAIL.n114 8.92171
R1059 VTAIL.n75 VTAIL.n64 8.92171
R1060 VTAIL.n170 VTAIL.n169 8.14595
R1061 VTAIL.n20 VTAIL.n19 8.14595
R1062 VTAIL.n122 VTAIL.n121 8.14595
R1063 VTAIL.n72 VTAIL.n71 8.14595
R1064 VTAIL.n166 VTAIL.n164 7.3702
R1065 VTAIL.n16 VTAIL.n14 7.3702
R1066 VTAIL.n118 VTAIL.n116 7.3702
R1067 VTAIL.n68 VTAIL.n66 7.3702
R1068 VTAIL.n169 VTAIL.n164 5.81868
R1069 VTAIL.n19 VTAIL.n14 5.81868
R1070 VTAIL.n121 VTAIL.n116 5.81868
R1071 VTAIL.n71 VTAIL.n66 5.81868
R1072 VTAIL.n170 VTAIL.n162 5.04292
R1073 VTAIL.n20 VTAIL.n12 5.04292
R1074 VTAIL.n122 VTAIL.n114 5.04292
R1075 VTAIL.n72 VTAIL.n64 5.04292
R1076 VTAIL.n174 VTAIL.n173 4.26717
R1077 VTAIL.n24 VTAIL.n23 4.26717
R1078 VTAIL.n126 VTAIL.n125 4.26717
R1079 VTAIL.n76 VTAIL.n75 4.26717
R1080 VTAIL.n177 VTAIL.n160 3.49141
R1081 VTAIL.n27 VTAIL.n10 3.49141
R1082 VTAIL.n129 VTAIL.n112 3.49141
R1083 VTAIL.n79 VTAIL.n62 3.49141
R1084 VTAIL.n178 VTAIL.n158 2.71565
R1085 VTAIL.n198 VTAIL.n150 2.71565
R1086 VTAIL.n28 VTAIL.n8 2.71565
R1087 VTAIL.n48 VTAIL.n0 2.71565
R1088 VTAIL.n148 VTAIL.n100 2.71565
R1089 VTAIL.n130 VTAIL.n110 2.71565
R1090 VTAIL.n98 VTAIL.n50 2.71565
R1091 VTAIL.n80 VTAIL.n60 2.71565
R1092 VTAIL.n165 VTAIL.n163 2.41283
R1093 VTAIL.n15 VTAIL.n13 2.41283
R1094 VTAIL.n117 VTAIL.n115 2.41283
R1095 VTAIL.n67 VTAIL.n65 2.41283
R1096 VTAIL.n149 VTAIL.n99 2.12981
R1097 VTAIL.n183 VTAIL.n181 1.93989
R1098 VTAIL.n196 VTAIL.n195 1.93989
R1099 VTAIL.n33 VTAIL.n31 1.93989
R1100 VTAIL.n46 VTAIL.n45 1.93989
R1101 VTAIL.n146 VTAIL.n145 1.93989
R1102 VTAIL.n134 VTAIL.n133 1.93989
R1103 VTAIL.n96 VTAIL.n95 1.93989
R1104 VTAIL.n84 VTAIL.n83 1.93989
R1105 VTAIL VTAIL.n49 1.35826
R1106 VTAIL.n182 VTAIL.n156 1.16414
R1107 VTAIL.n192 VTAIL.n152 1.16414
R1108 VTAIL.n32 VTAIL.n6 1.16414
R1109 VTAIL.n42 VTAIL.n2 1.16414
R1110 VTAIL.n142 VTAIL.n102 1.16414
R1111 VTAIL.n137 VTAIL.n107 1.16414
R1112 VTAIL.n92 VTAIL.n52 1.16414
R1113 VTAIL.n87 VTAIL.n57 1.16414
R1114 VTAIL VTAIL.n199 0.772052
R1115 VTAIL.n188 VTAIL.n187 0.388379
R1116 VTAIL.n191 VTAIL.n154 0.388379
R1117 VTAIL.n38 VTAIL.n37 0.388379
R1118 VTAIL.n41 VTAIL.n4 0.388379
R1119 VTAIL.n141 VTAIL.n104 0.388379
R1120 VTAIL.n138 VTAIL.n106 0.388379
R1121 VTAIL.n91 VTAIL.n54 0.388379
R1122 VTAIL.n88 VTAIL.n56 0.388379
R1123 VTAIL.n171 VTAIL.n163 0.155672
R1124 VTAIL.n172 VTAIL.n171 0.155672
R1125 VTAIL.n172 VTAIL.n159 0.155672
R1126 VTAIL.n179 VTAIL.n159 0.155672
R1127 VTAIL.n180 VTAIL.n179 0.155672
R1128 VTAIL.n180 VTAIL.n155 0.155672
R1129 VTAIL.n189 VTAIL.n155 0.155672
R1130 VTAIL.n190 VTAIL.n189 0.155672
R1131 VTAIL.n190 VTAIL.n151 0.155672
R1132 VTAIL.n197 VTAIL.n151 0.155672
R1133 VTAIL.n21 VTAIL.n13 0.155672
R1134 VTAIL.n22 VTAIL.n21 0.155672
R1135 VTAIL.n22 VTAIL.n9 0.155672
R1136 VTAIL.n29 VTAIL.n9 0.155672
R1137 VTAIL.n30 VTAIL.n29 0.155672
R1138 VTAIL.n30 VTAIL.n5 0.155672
R1139 VTAIL.n39 VTAIL.n5 0.155672
R1140 VTAIL.n40 VTAIL.n39 0.155672
R1141 VTAIL.n40 VTAIL.n1 0.155672
R1142 VTAIL.n47 VTAIL.n1 0.155672
R1143 VTAIL.n147 VTAIL.n101 0.155672
R1144 VTAIL.n140 VTAIL.n101 0.155672
R1145 VTAIL.n140 VTAIL.n139 0.155672
R1146 VTAIL.n139 VTAIL.n105 0.155672
R1147 VTAIL.n132 VTAIL.n105 0.155672
R1148 VTAIL.n132 VTAIL.n131 0.155672
R1149 VTAIL.n131 VTAIL.n111 0.155672
R1150 VTAIL.n124 VTAIL.n111 0.155672
R1151 VTAIL.n124 VTAIL.n123 0.155672
R1152 VTAIL.n123 VTAIL.n115 0.155672
R1153 VTAIL.n97 VTAIL.n51 0.155672
R1154 VTAIL.n90 VTAIL.n51 0.155672
R1155 VTAIL.n90 VTAIL.n89 0.155672
R1156 VTAIL.n89 VTAIL.n55 0.155672
R1157 VTAIL.n82 VTAIL.n55 0.155672
R1158 VTAIL.n82 VTAIL.n81 0.155672
R1159 VTAIL.n81 VTAIL.n61 0.155672
R1160 VTAIL.n74 VTAIL.n61 0.155672
R1161 VTAIL.n74 VTAIL.n73 0.155672
R1162 VTAIL.n73 VTAIL.n65 0.155672
R1163 VDD2.n93 VDD2.n49 756.745
R1164 VDD2.n44 VDD2.n0 756.745
R1165 VDD2.n94 VDD2.n93 585
R1166 VDD2.n92 VDD2.n91 585
R1167 VDD2.n53 VDD2.n52 585
R1168 VDD2.n57 VDD2.n55 585
R1169 VDD2.n86 VDD2.n85 585
R1170 VDD2.n84 VDD2.n83 585
R1171 VDD2.n59 VDD2.n58 585
R1172 VDD2.n78 VDD2.n77 585
R1173 VDD2.n76 VDD2.n75 585
R1174 VDD2.n63 VDD2.n62 585
R1175 VDD2.n70 VDD2.n69 585
R1176 VDD2.n68 VDD2.n67 585
R1177 VDD2.n17 VDD2.n16 585
R1178 VDD2.n19 VDD2.n18 585
R1179 VDD2.n12 VDD2.n11 585
R1180 VDD2.n25 VDD2.n24 585
R1181 VDD2.n27 VDD2.n26 585
R1182 VDD2.n8 VDD2.n7 585
R1183 VDD2.n34 VDD2.n33 585
R1184 VDD2.n35 VDD2.n6 585
R1185 VDD2.n37 VDD2.n36 585
R1186 VDD2.n4 VDD2.n3 585
R1187 VDD2.n43 VDD2.n42 585
R1188 VDD2.n45 VDD2.n44 585
R1189 VDD2.n66 VDD2.t1 329.038
R1190 VDD2.n15 VDD2.t0 329.038
R1191 VDD2.n93 VDD2.n92 171.744
R1192 VDD2.n92 VDD2.n52 171.744
R1193 VDD2.n57 VDD2.n52 171.744
R1194 VDD2.n85 VDD2.n57 171.744
R1195 VDD2.n85 VDD2.n84 171.744
R1196 VDD2.n84 VDD2.n58 171.744
R1197 VDD2.n77 VDD2.n58 171.744
R1198 VDD2.n77 VDD2.n76 171.744
R1199 VDD2.n76 VDD2.n62 171.744
R1200 VDD2.n69 VDD2.n62 171.744
R1201 VDD2.n69 VDD2.n68 171.744
R1202 VDD2.n18 VDD2.n17 171.744
R1203 VDD2.n18 VDD2.n11 171.744
R1204 VDD2.n25 VDD2.n11 171.744
R1205 VDD2.n26 VDD2.n25 171.744
R1206 VDD2.n26 VDD2.n7 171.744
R1207 VDD2.n34 VDD2.n7 171.744
R1208 VDD2.n35 VDD2.n34 171.744
R1209 VDD2.n36 VDD2.n35 171.744
R1210 VDD2.n36 VDD2.n3 171.744
R1211 VDD2.n43 VDD2.n3 171.744
R1212 VDD2.n44 VDD2.n43 171.744
R1213 VDD2.n98 VDD2.n48 87.5321
R1214 VDD2.n68 VDD2.t1 85.8723
R1215 VDD2.n17 VDD2.t0 85.8723
R1216 VDD2.n98 VDD2.n97 49.252
R1217 VDD2.n55 VDD2.n53 13.1884
R1218 VDD2.n37 VDD2.n4 13.1884
R1219 VDD2.n91 VDD2.n90 12.8005
R1220 VDD2.n87 VDD2.n86 12.8005
R1221 VDD2.n38 VDD2.n6 12.8005
R1222 VDD2.n42 VDD2.n41 12.8005
R1223 VDD2.n94 VDD2.n51 12.0247
R1224 VDD2.n83 VDD2.n56 12.0247
R1225 VDD2.n33 VDD2.n32 12.0247
R1226 VDD2.n45 VDD2.n2 12.0247
R1227 VDD2.n95 VDD2.n49 11.249
R1228 VDD2.n82 VDD2.n59 11.249
R1229 VDD2.n31 VDD2.n8 11.249
R1230 VDD2.n46 VDD2.n0 11.249
R1231 VDD2.n67 VDD2.n66 10.7239
R1232 VDD2.n16 VDD2.n15 10.7239
R1233 VDD2.n79 VDD2.n78 10.4732
R1234 VDD2.n28 VDD2.n27 10.4732
R1235 VDD2.n75 VDD2.n61 9.69747
R1236 VDD2.n24 VDD2.n10 9.69747
R1237 VDD2.n97 VDD2.n96 9.45567
R1238 VDD2.n48 VDD2.n47 9.45567
R1239 VDD2.n65 VDD2.n64 9.3005
R1240 VDD2.n72 VDD2.n71 9.3005
R1241 VDD2.n74 VDD2.n73 9.3005
R1242 VDD2.n61 VDD2.n60 9.3005
R1243 VDD2.n80 VDD2.n79 9.3005
R1244 VDD2.n82 VDD2.n81 9.3005
R1245 VDD2.n56 VDD2.n54 9.3005
R1246 VDD2.n88 VDD2.n87 9.3005
R1247 VDD2.n96 VDD2.n95 9.3005
R1248 VDD2.n51 VDD2.n50 9.3005
R1249 VDD2.n90 VDD2.n89 9.3005
R1250 VDD2.n47 VDD2.n46 9.3005
R1251 VDD2.n2 VDD2.n1 9.3005
R1252 VDD2.n41 VDD2.n40 9.3005
R1253 VDD2.n14 VDD2.n13 9.3005
R1254 VDD2.n21 VDD2.n20 9.3005
R1255 VDD2.n23 VDD2.n22 9.3005
R1256 VDD2.n10 VDD2.n9 9.3005
R1257 VDD2.n29 VDD2.n28 9.3005
R1258 VDD2.n31 VDD2.n30 9.3005
R1259 VDD2.n32 VDD2.n5 9.3005
R1260 VDD2.n39 VDD2.n38 9.3005
R1261 VDD2.n74 VDD2.n63 8.92171
R1262 VDD2.n23 VDD2.n12 8.92171
R1263 VDD2.n71 VDD2.n70 8.14595
R1264 VDD2.n20 VDD2.n19 8.14595
R1265 VDD2.n67 VDD2.n65 7.3702
R1266 VDD2.n16 VDD2.n14 7.3702
R1267 VDD2.n70 VDD2.n65 5.81868
R1268 VDD2.n19 VDD2.n14 5.81868
R1269 VDD2.n71 VDD2.n63 5.04292
R1270 VDD2.n20 VDD2.n12 5.04292
R1271 VDD2.n75 VDD2.n74 4.26717
R1272 VDD2.n24 VDD2.n23 4.26717
R1273 VDD2.n78 VDD2.n61 3.49141
R1274 VDD2.n27 VDD2.n10 3.49141
R1275 VDD2.n97 VDD2.n49 2.71565
R1276 VDD2.n79 VDD2.n59 2.71565
R1277 VDD2.n28 VDD2.n8 2.71565
R1278 VDD2.n48 VDD2.n0 2.71565
R1279 VDD2.n66 VDD2.n64 2.41283
R1280 VDD2.n15 VDD2.n13 2.41283
R1281 VDD2.n95 VDD2.n94 1.93989
R1282 VDD2.n83 VDD2.n82 1.93989
R1283 VDD2.n33 VDD2.n31 1.93989
R1284 VDD2.n46 VDD2.n45 1.93989
R1285 VDD2.n91 VDD2.n51 1.16414
R1286 VDD2.n86 VDD2.n56 1.16414
R1287 VDD2.n32 VDD2.n6 1.16414
R1288 VDD2.n42 VDD2.n2 1.16414
R1289 VDD2 VDD2.n98 0.888431
R1290 VDD2.n90 VDD2.n53 0.388379
R1291 VDD2.n87 VDD2.n55 0.388379
R1292 VDD2.n38 VDD2.n37 0.388379
R1293 VDD2.n41 VDD2.n4 0.388379
R1294 VDD2.n96 VDD2.n50 0.155672
R1295 VDD2.n89 VDD2.n50 0.155672
R1296 VDD2.n89 VDD2.n88 0.155672
R1297 VDD2.n88 VDD2.n54 0.155672
R1298 VDD2.n81 VDD2.n54 0.155672
R1299 VDD2.n81 VDD2.n80 0.155672
R1300 VDD2.n80 VDD2.n60 0.155672
R1301 VDD2.n73 VDD2.n60 0.155672
R1302 VDD2.n73 VDD2.n72 0.155672
R1303 VDD2.n72 VDD2.n64 0.155672
R1304 VDD2.n21 VDD2.n13 0.155672
R1305 VDD2.n22 VDD2.n21 0.155672
R1306 VDD2.n22 VDD2.n9 0.155672
R1307 VDD2.n29 VDD2.n9 0.155672
R1308 VDD2.n30 VDD2.n29 0.155672
R1309 VDD2.n30 VDD2.n5 0.155672
R1310 VDD2.n39 VDD2.n5 0.155672
R1311 VDD2.n40 VDD2.n39 0.155672
R1312 VDD2.n40 VDD2.n1 0.155672
R1313 VDD2.n47 VDD2.n1 0.155672
R1314 VP.n0 VP.t1 147.266
R1315 VP.n0 VP.t0 102.246
R1316 VP VP.n0 0.526373
R1317 VDD1.n44 VDD1.n0 756.745
R1318 VDD1.n93 VDD1.n49 756.745
R1319 VDD1.n45 VDD1.n44 585
R1320 VDD1.n43 VDD1.n42 585
R1321 VDD1.n4 VDD1.n3 585
R1322 VDD1.n8 VDD1.n6 585
R1323 VDD1.n37 VDD1.n36 585
R1324 VDD1.n35 VDD1.n34 585
R1325 VDD1.n10 VDD1.n9 585
R1326 VDD1.n29 VDD1.n28 585
R1327 VDD1.n27 VDD1.n26 585
R1328 VDD1.n14 VDD1.n13 585
R1329 VDD1.n21 VDD1.n20 585
R1330 VDD1.n19 VDD1.n18 585
R1331 VDD1.n66 VDD1.n65 585
R1332 VDD1.n68 VDD1.n67 585
R1333 VDD1.n61 VDD1.n60 585
R1334 VDD1.n74 VDD1.n73 585
R1335 VDD1.n76 VDD1.n75 585
R1336 VDD1.n57 VDD1.n56 585
R1337 VDD1.n83 VDD1.n82 585
R1338 VDD1.n84 VDD1.n55 585
R1339 VDD1.n86 VDD1.n85 585
R1340 VDD1.n53 VDD1.n52 585
R1341 VDD1.n92 VDD1.n91 585
R1342 VDD1.n94 VDD1.n93 585
R1343 VDD1.n17 VDD1.t0 329.038
R1344 VDD1.n64 VDD1.t1 329.038
R1345 VDD1.n44 VDD1.n43 171.744
R1346 VDD1.n43 VDD1.n3 171.744
R1347 VDD1.n8 VDD1.n3 171.744
R1348 VDD1.n36 VDD1.n8 171.744
R1349 VDD1.n36 VDD1.n35 171.744
R1350 VDD1.n35 VDD1.n9 171.744
R1351 VDD1.n28 VDD1.n9 171.744
R1352 VDD1.n28 VDD1.n27 171.744
R1353 VDD1.n27 VDD1.n13 171.744
R1354 VDD1.n20 VDD1.n13 171.744
R1355 VDD1.n20 VDD1.n19 171.744
R1356 VDD1.n67 VDD1.n66 171.744
R1357 VDD1.n67 VDD1.n60 171.744
R1358 VDD1.n74 VDD1.n60 171.744
R1359 VDD1.n75 VDD1.n74 171.744
R1360 VDD1.n75 VDD1.n56 171.744
R1361 VDD1.n83 VDD1.n56 171.744
R1362 VDD1.n84 VDD1.n83 171.744
R1363 VDD1.n85 VDD1.n84 171.744
R1364 VDD1.n85 VDD1.n52 171.744
R1365 VDD1.n92 VDD1.n52 171.744
R1366 VDD1.n93 VDD1.n92 171.744
R1367 VDD1 VDD1.n97 88.8867
R1368 VDD1.n19 VDD1.t0 85.8723
R1369 VDD1.n66 VDD1.t1 85.8723
R1370 VDD1 VDD1.n48 50.1399
R1371 VDD1.n6 VDD1.n4 13.1884
R1372 VDD1.n86 VDD1.n53 13.1884
R1373 VDD1.n42 VDD1.n41 12.8005
R1374 VDD1.n38 VDD1.n37 12.8005
R1375 VDD1.n87 VDD1.n55 12.8005
R1376 VDD1.n91 VDD1.n90 12.8005
R1377 VDD1.n45 VDD1.n2 12.0247
R1378 VDD1.n34 VDD1.n7 12.0247
R1379 VDD1.n82 VDD1.n81 12.0247
R1380 VDD1.n94 VDD1.n51 12.0247
R1381 VDD1.n46 VDD1.n0 11.249
R1382 VDD1.n33 VDD1.n10 11.249
R1383 VDD1.n80 VDD1.n57 11.249
R1384 VDD1.n95 VDD1.n49 11.249
R1385 VDD1.n18 VDD1.n17 10.7239
R1386 VDD1.n65 VDD1.n64 10.7239
R1387 VDD1.n30 VDD1.n29 10.4732
R1388 VDD1.n77 VDD1.n76 10.4732
R1389 VDD1.n26 VDD1.n12 9.69747
R1390 VDD1.n73 VDD1.n59 9.69747
R1391 VDD1.n48 VDD1.n47 9.45567
R1392 VDD1.n97 VDD1.n96 9.45567
R1393 VDD1.n16 VDD1.n15 9.3005
R1394 VDD1.n23 VDD1.n22 9.3005
R1395 VDD1.n25 VDD1.n24 9.3005
R1396 VDD1.n12 VDD1.n11 9.3005
R1397 VDD1.n31 VDD1.n30 9.3005
R1398 VDD1.n33 VDD1.n32 9.3005
R1399 VDD1.n7 VDD1.n5 9.3005
R1400 VDD1.n39 VDD1.n38 9.3005
R1401 VDD1.n47 VDD1.n46 9.3005
R1402 VDD1.n2 VDD1.n1 9.3005
R1403 VDD1.n41 VDD1.n40 9.3005
R1404 VDD1.n96 VDD1.n95 9.3005
R1405 VDD1.n51 VDD1.n50 9.3005
R1406 VDD1.n90 VDD1.n89 9.3005
R1407 VDD1.n63 VDD1.n62 9.3005
R1408 VDD1.n70 VDD1.n69 9.3005
R1409 VDD1.n72 VDD1.n71 9.3005
R1410 VDD1.n59 VDD1.n58 9.3005
R1411 VDD1.n78 VDD1.n77 9.3005
R1412 VDD1.n80 VDD1.n79 9.3005
R1413 VDD1.n81 VDD1.n54 9.3005
R1414 VDD1.n88 VDD1.n87 9.3005
R1415 VDD1.n25 VDD1.n14 8.92171
R1416 VDD1.n72 VDD1.n61 8.92171
R1417 VDD1.n22 VDD1.n21 8.14595
R1418 VDD1.n69 VDD1.n68 8.14595
R1419 VDD1.n18 VDD1.n16 7.3702
R1420 VDD1.n65 VDD1.n63 7.3702
R1421 VDD1.n21 VDD1.n16 5.81868
R1422 VDD1.n68 VDD1.n63 5.81868
R1423 VDD1.n22 VDD1.n14 5.04292
R1424 VDD1.n69 VDD1.n61 5.04292
R1425 VDD1.n26 VDD1.n25 4.26717
R1426 VDD1.n73 VDD1.n72 4.26717
R1427 VDD1.n29 VDD1.n12 3.49141
R1428 VDD1.n76 VDD1.n59 3.49141
R1429 VDD1.n48 VDD1.n0 2.71565
R1430 VDD1.n30 VDD1.n10 2.71565
R1431 VDD1.n77 VDD1.n57 2.71565
R1432 VDD1.n97 VDD1.n49 2.71565
R1433 VDD1.n17 VDD1.n15 2.41283
R1434 VDD1.n64 VDD1.n62 2.41283
R1435 VDD1.n46 VDD1.n45 1.93989
R1436 VDD1.n34 VDD1.n33 1.93989
R1437 VDD1.n82 VDD1.n80 1.93989
R1438 VDD1.n95 VDD1.n94 1.93989
R1439 VDD1.n42 VDD1.n2 1.16414
R1440 VDD1.n37 VDD1.n7 1.16414
R1441 VDD1.n81 VDD1.n55 1.16414
R1442 VDD1.n91 VDD1.n51 1.16414
R1443 VDD1.n41 VDD1.n4 0.388379
R1444 VDD1.n38 VDD1.n6 0.388379
R1445 VDD1.n87 VDD1.n86 0.388379
R1446 VDD1.n90 VDD1.n53 0.388379
R1447 VDD1.n47 VDD1.n1 0.155672
R1448 VDD1.n40 VDD1.n1 0.155672
R1449 VDD1.n40 VDD1.n39 0.155672
R1450 VDD1.n39 VDD1.n5 0.155672
R1451 VDD1.n32 VDD1.n5 0.155672
R1452 VDD1.n32 VDD1.n31 0.155672
R1453 VDD1.n31 VDD1.n11 0.155672
R1454 VDD1.n24 VDD1.n11 0.155672
R1455 VDD1.n24 VDD1.n23 0.155672
R1456 VDD1.n23 VDD1.n15 0.155672
R1457 VDD1.n70 VDD1.n62 0.155672
R1458 VDD1.n71 VDD1.n70 0.155672
R1459 VDD1.n71 VDD1.n58 0.155672
R1460 VDD1.n78 VDD1.n58 0.155672
R1461 VDD1.n79 VDD1.n78 0.155672
R1462 VDD1.n79 VDD1.n54 0.155672
R1463 VDD1.n88 VDD1.n54 0.155672
R1464 VDD1.n89 VDD1.n88 0.155672
R1465 VDD1.n89 VDD1.n50 0.155672
R1466 VDD1.n96 VDD1.n50 0.155672
C0 w_n2510_n2820# VDD1 1.69769f
C1 VP VN 5.37492f
C2 B VN 1.17691f
C3 VTAIL VDD2 4.61342f
C4 B VP 1.70951f
C5 VDD1 VN 0.148879f
C6 w_n2510_n2820# VDD2 1.73495f
C7 VDD1 VP 2.51325f
C8 B VDD1 1.60687f
C9 w_n2510_n2820# VTAIL 2.39691f
C10 VDD2 VN 2.29204f
C11 VP VDD2 0.371888f
C12 B VDD2 1.64515f
C13 VTAIL VN 2.14624f
C14 VTAIL VP 2.16044f
C15 B VTAIL 3.35084f
C16 VDD1 VDD2 0.774892f
C17 w_n2510_n2820# VN 3.49543f
C18 w_n2510_n2820# VP 3.81714f
C19 B w_n2510_n2820# 9.03462f
C20 VDD1 VTAIL 4.55539f
C21 VDD2 VSUBS 0.897865f
C22 VDD1 VSUBS 3.72461f
C23 VTAIL VSUBS 0.993851f
C24 VN VSUBS 7.63139f
C25 VP VSUBS 1.869541f
C26 B VSUBS 4.351936f
C27 w_n2510_n2820# VSUBS 87.5588f
C28 VDD1.n0 VSUBS 0.021825f
C29 VDD1.n1 VSUBS 0.021081f
C30 VDD1.n2 VSUBS 0.011328f
C31 VDD1.n3 VSUBS 0.026776f
C32 VDD1.n4 VSUBS 0.011661f
C33 VDD1.n5 VSUBS 0.021081f
C34 VDD1.n6 VSUBS 0.011661f
C35 VDD1.n7 VSUBS 0.011328f
C36 VDD1.n8 VSUBS 0.026776f
C37 VDD1.n9 VSUBS 0.026776f
C38 VDD1.n10 VSUBS 0.011995f
C39 VDD1.n11 VSUBS 0.021081f
C40 VDD1.n12 VSUBS 0.011328f
C41 VDD1.n13 VSUBS 0.026776f
C42 VDD1.n14 VSUBS 0.011995f
C43 VDD1.n15 VSUBS 0.782654f
C44 VDD1.n16 VSUBS 0.011328f
C45 VDD1.t0 VSUBS 0.05753f
C46 VDD1.n17 VSUBS 0.139933f
C47 VDD1.n18 VSUBS 0.020142f
C48 VDD1.n19 VSUBS 0.020082f
C49 VDD1.n20 VSUBS 0.026776f
C50 VDD1.n21 VSUBS 0.011995f
C51 VDD1.n22 VSUBS 0.011328f
C52 VDD1.n23 VSUBS 0.021081f
C53 VDD1.n24 VSUBS 0.021081f
C54 VDD1.n25 VSUBS 0.011328f
C55 VDD1.n26 VSUBS 0.011995f
C56 VDD1.n27 VSUBS 0.026776f
C57 VDD1.n28 VSUBS 0.026776f
C58 VDD1.n29 VSUBS 0.011995f
C59 VDD1.n30 VSUBS 0.011328f
C60 VDD1.n31 VSUBS 0.021081f
C61 VDD1.n32 VSUBS 0.021081f
C62 VDD1.n33 VSUBS 0.011328f
C63 VDD1.n34 VSUBS 0.011995f
C64 VDD1.n35 VSUBS 0.026776f
C65 VDD1.n36 VSUBS 0.026776f
C66 VDD1.n37 VSUBS 0.011995f
C67 VDD1.n38 VSUBS 0.011328f
C68 VDD1.n39 VSUBS 0.021081f
C69 VDD1.n40 VSUBS 0.021081f
C70 VDD1.n41 VSUBS 0.011328f
C71 VDD1.n42 VSUBS 0.011995f
C72 VDD1.n43 VSUBS 0.026776f
C73 VDD1.n44 VSUBS 0.06026f
C74 VDD1.n45 VSUBS 0.011995f
C75 VDD1.n46 VSUBS 0.011328f
C76 VDD1.n47 VSUBS 0.049305f
C77 VDD1.n48 VSUBS 0.046464f
C78 VDD1.n49 VSUBS 0.021825f
C79 VDD1.n50 VSUBS 0.021081f
C80 VDD1.n51 VSUBS 0.011328f
C81 VDD1.n52 VSUBS 0.026776f
C82 VDD1.n53 VSUBS 0.011661f
C83 VDD1.n54 VSUBS 0.021081f
C84 VDD1.n55 VSUBS 0.011995f
C85 VDD1.n56 VSUBS 0.026776f
C86 VDD1.n57 VSUBS 0.011995f
C87 VDD1.n58 VSUBS 0.021081f
C88 VDD1.n59 VSUBS 0.011328f
C89 VDD1.n60 VSUBS 0.026776f
C90 VDD1.n61 VSUBS 0.011995f
C91 VDD1.n62 VSUBS 0.782654f
C92 VDD1.n63 VSUBS 0.011328f
C93 VDD1.t1 VSUBS 0.05753f
C94 VDD1.n64 VSUBS 0.139933f
C95 VDD1.n65 VSUBS 0.020142f
C96 VDD1.n66 VSUBS 0.020082f
C97 VDD1.n67 VSUBS 0.026776f
C98 VDD1.n68 VSUBS 0.011995f
C99 VDD1.n69 VSUBS 0.011328f
C100 VDD1.n70 VSUBS 0.021081f
C101 VDD1.n71 VSUBS 0.021081f
C102 VDD1.n72 VSUBS 0.011328f
C103 VDD1.n73 VSUBS 0.011995f
C104 VDD1.n74 VSUBS 0.026776f
C105 VDD1.n75 VSUBS 0.026776f
C106 VDD1.n76 VSUBS 0.011995f
C107 VDD1.n77 VSUBS 0.011328f
C108 VDD1.n78 VSUBS 0.021081f
C109 VDD1.n79 VSUBS 0.021081f
C110 VDD1.n80 VSUBS 0.011328f
C111 VDD1.n81 VSUBS 0.011328f
C112 VDD1.n82 VSUBS 0.011995f
C113 VDD1.n83 VSUBS 0.026776f
C114 VDD1.n84 VSUBS 0.026776f
C115 VDD1.n85 VSUBS 0.026776f
C116 VDD1.n86 VSUBS 0.011661f
C117 VDD1.n87 VSUBS 0.011328f
C118 VDD1.n88 VSUBS 0.021081f
C119 VDD1.n89 VSUBS 0.021081f
C120 VDD1.n90 VSUBS 0.011328f
C121 VDD1.n91 VSUBS 0.011995f
C122 VDD1.n92 VSUBS 0.026776f
C123 VDD1.n93 VSUBS 0.06026f
C124 VDD1.n94 VSUBS 0.011995f
C125 VDD1.n95 VSUBS 0.011328f
C126 VDD1.n96 VSUBS 0.049305f
C127 VDD1.n97 VSUBS 0.630594f
C128 VP.t1 VSUBS 4.85192f
C129 VP.t0 VSUBS 3.93481f
C130 VP.n0 VSUBS 4.96978f
C131 VDD2.n0 VSUBS 0.021445f
C132 VDD2.n1 VSUBS 0.020715f
C133 VDD2.n2 VSUBS 0.011131f
C134 VDD2.n3 VSUBS 0.02631f
C135 VDD2.n4 VSUBS 0.011459f
C136 VDD2.n5 VSUBS 0.020715f
C137 VDD2.n6 VSUBS 0.011786f
C138 VDD2.n7 VSUBS 0.02631f
C139 VDD2.n8 VSUBS 0.011786f
C140 VDD2.n9 VSUBS 0.020715f
C141 VDD2.n10 VSUBS 0.011131f
C142 VDD2.n11 VSUBS 0.02631f
C143 VDD2.n12 VSUBS 0.011786f
C144 VDD2.n13 VSUBS 0.769041f
C145 VDD2.n14 VSUBS 0.011131f
C146 VDD2.t0 VSUBS 0.056529f
C147 VDD2.n15 VSUBS 0.137499f
C148 VDD2.n16 VSUBS 0.019792f
C149 VDD2.n17 VSUBS 0.019733f
C150 VDD2.n18 VSUBS 0.02631f
C151 VDD2.n19 VSUBS 0.011786f
C152 VDD2.n20 VSUBS 0.011131f
C153 VDD2.n21 VSUBS 0.020715f
C154 VDD2.n22 VSUBS 0.020715f
C155 VDD2.n23 VSUBS 0.011131f
C156 VDD2.n24 VSUBS 0.011786f
C157 VDD2.n25 VSUBS 0.02631f
C158 VDD2.n26 VSUBS 0.02631f
C159 VDD2.n27 VSUBS 0.011786f
C160 VDD2.n28 VSUBS 0.011131f
C161 VDD2.n29 VSUBS 0.020715f
C162 VDD2.n30 VSUBS 0.020715f
C163 VDD2.n31 VSUBS 0.011131f
C164 VDD2.n32 VSUBS 0.011131f
C165 VDD2.n33 VSUBS 0.011786f
C166 VDD2.n34 VSUBS 0.02631f
C167 VDD2.n35 VSUBS 0.02631f
C168 VDD2.n36 VSUBS 0.02631f
C169 VDD2.n37 VSUBS 0.011459f
C170 VDD2.n38 VSUBS 0.011131f
C171 VDD2.n39 VSUBS 0.020715f
C172 VDD2.n40 VSUBS 0.020715f
C173 VDD2.n41 VSUBS 0.011131f
C174 VDD2.n42 VSUBS 0.011786f
C175 VDD2.n43 VSUBS 0.02631f
C176 VDD2.n44 VSUBS 0.059212f
C177 VDD2.n45 VSUBS 0.011786f
C178 VDD2.n46 VSUBS 0.011131f
C179 VDD2.n47 VSUBS 0.048447f
C180 VDD2.n48 VSUBS 0.574519f
C181 VDD2.n49 VSUBS 0.021445f
C182 VDD2.n50 VSUBS 0.020715f
C183 VDD2.n51 VSUBS 0.011131f
C184 VDD2.n52 VSUBS 0.02631f
C185 VDD2.n53 VSUBS 0.011459f
C186 VDD2.n54 VSUBS 0.020715f
C187 VDD2.n55 VSUBS 0.011459f
C188 VDD2.n56 VSUBS 0.011131f
C189 VDD2.n57 VSUBS 0.02631f
C190 VDD2.n58 VSUBS 0.02631f
C191 VDD2.n59 VSUBS 0.011786f
C192 VDD2.n60 VSUBS 0.020715f
C193 VDD2.n61 VSUBS 0.011131f
C194 VDD2.n62 VSUBS 0.02631f
C195 VDD2.n63 VSUBS 0.011786f
C196 VDD2.n64 VSUBS 0.769041f
C197 VDD2.n65 VSUBS 0.011131f
C198 VDD2.t1 VSUBS 0.056529f
C199 VDD2.n66 VSUBS 0.137499f
C200 VDD2.n67 VSUBS 0.019792f
C201 VDD2.n68 VSUBS 0.019733f
C202 VDD2.n69 VSUBS 0.02631f
C203 VDD2.n70 VSUBS 0.011786f
C204 VDD2.n71 VSUBS 0.011131f
C205 VDD2.n72 VSUBS 0.020715f
C206 VDD2.n73 VSUBS 0.020715f
C207 VDD2.n74 VSUBS 0.011131f
C208 VDD2.n75 VSUBS 0.011786f
C209 VDD2.n76 VSUBS 0.02631f
C210 VDD2.n77 VSUBS 0.02631f
C211 VDD2.n78 VSUBS 0.011786f
C212 VDD2.n79 VSUBS 0.011131f
C213 VDD2.n80 VSUBS 0.020715f
C214 VDD2.n81 VSUBS 0.020715f
C215 VDD2.n82 VSUBS 0.011131f
C216 VDD2.n83 VSUBS 0.011786f
C217 VDD2.n84 VSUBS 0.02631f
C218 VDD2.n85 VSUBS 0.02631f
C219 VDD2.n86 VSUBS 0.011786f
C220 VDD2.n87 VSUBS 0.011131f
C221 VDD2.n88 VSUBS 0.020715f
C222 VDD2.n89 VSUBS 0.020715f
C223 VDD2.n90 VSUBS 0.011131f
C224 VDD2.n91 VSUBS 0.011786f
C225 VDD2.n92 VSUBS 0.02631f
C226 VDD2.n93 VSUBS 0.059212f
C227 VDD2.n94 VSUBS 0.011786f
C228 VDD2.n95 VSUBS 0.011131f
C229 VDD2.n96 VSUBS 0.048447f
C230 VDD2.n97 VSUBS 0.043894f
C231 VDD2.n98 VSUBS 2.44564f
C232 VTAIL.n0 VSUBS 0.032653f
C233 VTAIL.n1 VSUBS 0.03154f
C234 VTAIL.n2 VSUBS 0.016948f
C235 VTAIL.n3 VSUBS 0.04006f
C236 VTAIL.n4 VSUBS 0.017447f
C237 VTAIL.n5 VSUBS 0.03154f
C238 VTAIL.n6 VSUBS 0.017945f
C239 VTAIL.n7 VSUBS 0.04006f
C240 VTAIL.n8 VSUBS 0.017945f
C241 VTAIL.n9 VSUBS 0.03154f
C242 VTAIL.n10 VSUBS 0.016948f
C243 VTAIL.n11 VSUBS 0.04006f
C244 VTAIL.n12 VSUBS 0.017945f
C245 VTAIL.n13 VSUBS 1.17094f
C246 VTAIL.n14 VSUBS 0.016948f
C247 VTAIL.t0 VSUBS 0.086072f
C248 VTAIL.n15 VSUBS 0.209356f
C249 VTAIL.n16 VSUBS 0.030135f
C250 VTAIL.n17 VSUBS 0.030045f
C251 VTAIL.n18 VSUBS 0.04006f
C252 VTAIL.n19 VSUBS 0.017945f
C253 VTAIL.n20 VSUBS 0.016948f
C254 VTAIL.n21 VSUBS 0.03154f
C255 VTAIL.n22 VSUBS 0.03154f
C256 VTAIL.n23 VSUBS 0.016948f
C257 VTAIL.n24 VSUBS 0.017945f
C258 VTAIL.n25 VSUBS 0.04006f
C259 VTAIL.n26 VSUBS 0.04006f
C260 VTAIL.n27 VSUBS 0.017945f
C261 VTAIL.n28 VSUBS 0.016948f
C262 VTAIL.n29 VSUBS 0.03154f
C263 VTAIL.n30 VSUBS 0.03154f
C264 VTAIL.n31 VSUBS 0.016948f
C265 VTAIL.n32 VSUBS 0.016948f
C266 VTAIL.n33 VSUBS 0.017945f
C267 VTAIL.n34 VSUBS 0.04006f
C268 VTAIL.n35 VSUBS 0.04006f
C269 VTAIL.n36 VSUBS 0.04006f
C270 VTAIL.n37 VSUBS 0.017447f
C271 VTAIL.n38 VSUBS 0.016948f
C272 VTAIL.n39 VSUBS 0.03154f
C273 VTAIL.n40 VSUBS 0.03154f
C274 VTAIL.n41 VSUBS 0.016948f
C275 VTAIL.n42 VSUBS 0.017945f
C276 VTAIL.n43 VSUBS 0.04006f
C277 VTAIL.n44 VSUBS 0.090156f
C278 VTAIL.n45 VSUBS 0.017945f
C279 VTAIL.n46 VSUBS 0.016948f
C280 VTAIL.n47 VSUBS 0.073766f
C281 VTAIL.n48 VSUBS 0.045062f
C282 VTAIL.n49 VSUBS 2.07976f
C283 VTAIL.n50 VSUBS 0.032653f
C284 VTAIL.n51 VSUBS 0.03154f
C285 VTAIL.n52 VSUBS 0.016948f
C286 VTAIL.n53 VSUBS 0.04006f
C287 VTAIL.n54 VSUBS 0.017447f
C288 VTAIL.n55 VSUBS 0.03154f
C289 VTAIL.n56 VSUBS 0.017447f
C290 VTAIL.n57 VSUBS 0.016948f
C291 VTAIL.n58 VSUBS 0.04006f
C292 VTAIL.n59 VSUBS 0.04006f
C293 VTAIL.n60 VSUBS 0.017945f
C294 VTAIL.n61 VSUBS 0.03154f
C295 VTAIL.n62 VSUBS 0.016948f
C296 VTAIL.n63 VSUBS 0.04006f
C297 VTAIL.n64 VSUBS 0.017945f
C298 VTAIL.n65 VSUBS 1.17094f
C299 VTAIL.n66 VSUBS 0.016948f
C300 VTAIL.t3 VSUBS 0.086072f
C301 VTAIL.n67 VSUBS 0.209356f
C302 VTAIL.n68 VSUBS 0.030135f
C303 VTAIL.n69 VSUBS 0.030045f
C304 VTAIL.n70 VSUBS 0.04006f
C305 VTAIL.n71 VSUBS 0.017945f
C306 VTAIL.n72 VSUBS 0.016948f
C307 VTAIL.n73 VSUBS 0.03154f
C308 VTAIL.n74 VSUBS 0.03154f
C309 VTAIL.n75 VSUBS 0.016948f
C310 VTAIL.n76 VSUBS 0.017945f
C311 VTAIL.n77 VSUBS 0.04006f
C312 VTAIL.n78 VSUBS 0.04006f
C313 VTAIL.n79 VSUBS 0.017945f
C314 VTAIL.n80 VSUBS 0.016948f
C315 VTAIL.n81 VSUBS 0.03154f
C316 VTAIL.n82 VSUBS 0.03154f
C317 VTAIL.n83 VSUBS 0.016948f
C318 VTAIL.n84 VSUBS 0.017945f
C319 VTAIL.n85 VSUBS 0.04006f
C320 VTAIL.n86 VSUBS 0.04006f
C321 VTAIL.n87 VSUBS 0.017945f
C322 VTAIL.n88 VSUBS 0.016948f
C323 VTAIL.n89 VSUBS 0.03154f
C324 VTAIL.n90 VSUBS 0.03154f
C325 VTAIL.n91 VSUBS 0.016948f
C326 VTAIL.n92 VSUBS 0.017945f
C327 VTAIL.n93 VSUBS 0.04006f
C328 VTAIL.n94 VSUBS 0.090156f
C329 VTAIL.n95 VSUBS 0.017945f
C330 VTAIL.n96 VSUBS 0.016948f
C331 VTAIL.n97 VSUBS 0.073766f
C332 VTAIL.n98 VSUBS 0.045062f
C333 VTAIL.n99 VSUBS 2.15817f
C334 VTAIL.n100 VSUBS 0.032653f
C335 VTAIL.n101 VSUBS 0.03154f
C336 VTAIL.n102 VSUBS 0.016948f
C337 VTAIL.n103 VSUBS 0.04006f
C338 VTAIL.n104 VSUBS 0.017447f
C339 VTAIL.n105 VSUBS 0.03154f
C340 VTAIL.n106 VSUBS 0.017447f
C341 VTAIL.n107 VSUBS 0.016948f
C342 VTAIL.n108 VSUBS 0.04006f
C343 VTAIL.n109 VSUBS 0.04006f
C344 VTAIL.n110 VSUBS 0.017945f
C345 VTAIL.n111 VSUBS 0.03154f
C346 VTAIL.n112 VSUBS 0.016948f
C347 VTAIL.n113 VSUBS 0.04006f
C348 VTAIL.n114 VSUBS 0.017945f
C349 VTAIL.n115 VSUBS 1.17094f
C350 VTAIL.n116 VSUBS 0.016948f
C351 VTAIL.t1 VSUBS 0.086072f
C352 VTAIL.n117 VSUBS 0.209356f
C353 VTAIL.n118 VSUBS 0.030135f
C354 VTAIL.n119 VSUBS 0.030045f
C355 VTAIL.n120 VSUBS 0.04006f
C356 VTAIL.n121 VSUBS 0.017945f
C357 VTAIL.n122 VSUBS 0.016948f
C358 VTAIL.n123 VSUBS 0.03154f
C359 VTAIL.n124 VSUBS 0.03154f
C360 VTAIL.n125 VSUBS 0.016948f
C361 VTAIL.n126 VSUBS 0.017945f
C362 VTAIL.n127 VSUBS 0.04006f
C363 VTAIL.n128 VSUBS 0.04006f
C364 VTAIL.n129 VSUBS 0.017945f
C365 VTAIL.n130 VSUBS 0.016948f
C366 VTAIL.n131 VSUBS 0.03154f
C367 VTAIL.n132 VSUBS 0.03154f
C368 VTAIL.n133 VSUBS 0.016948f
C369 VTAIL.n134 VSUBS 0.017945f
C370 VTAIL.n135 VSUBS 0.04006f
C371 VTAIL.n136 VSUBS 0.04006f
C372 VTAIL.n137 VSUBS 0.017945f
C373 VTAIL.n138 VSUBS 0.016948f
C374 VTAIL.n139 VSUBS 0.03154f
C375 VTAIL.n140 VSUBS 0.03154f
C376 VTAIL.n141 VSUBS 0.016948f
C377 VTAIL.n142 VSUBS 0.017945f
C378 VTAIL.n143 VSUBS 0.04006f
C379 VTAIL.n144 VSUBS 0.090156f
C380 VTAIL.n145 VSUBS 0.017945f
C381 VTAIL.n146 VSUBS 0.016948f
C382 VTAIL.n147 VSUBS 0.073766f
C383 VTAIL.n148 VSUBS 0.045062f
C384 VTAIL.n149 VSUBS 1.82086f
C385 VTAIL.n150 VSUBS 0.032653f
C386 VTAIL.n151 VSUBS 0.03154f
C387 VTAIL.n152 VSUBS 0.016948f
C388 VTAIL.n153 VSUBS 0.04006f
C389 VTAIL.n154 VSUBS 0.017447f
C390 VTAIL.n155 VSUBS 0.03154f
C391 VTAIL.n156 VSUBS 0.017945f
C392 VTAIL.n157 VSUBS 0.04006f
C393 VTAIL.n158 VSUBS 0.017945f
C394 VTAIL.n159 VSUBS 0.03154f
C395 VTAIL.n160 VSUBS 0.016948f
C396 VTAIL.n161 VSUBS 0.04006f
C397 VTAIL.n162 VSUBS 0.017945f
C398 VTAIL.n163 VSUBS 1.17094f
C399 VTAIL.n164 VSUBS 0.016948f
C400 VTAIL.t2 VSUBS 0.086072f
C401 VTAIL.n165 VSUBS 0.209356f
C402 VTAIL.n166 VSUBS 0.030135f
C403 VTAIL.n167 VSUBS 0.030045f
C404 VTAIL.n168 VSUBS 0.04006f
C405 VTAIL.n169 VSUBS 0.017945f
C406 VTAIL.n170 VSUBS 0.016948f
C407 VTAIL.n171 VSUBS 0.03154f
C408 VTAIL.n172 VSUBS 0.03154f
C409 VTAIL.n173 VSUBS 0.016948f
C410 VTAIL.n174 VSUBS 0.017945f
C411 VTAIL.n175 VSUBS 0.04006f
C412 VTAIL.n176 VSUBS 0.04006f
C413 VTAIL.n177 VSUBS 0.017945f
C414 VTAIL.n178 VSUBS 0.016948f
C415 VTAIL.n179 VSUBS 0.03154f
C416 VTAIL.n180 VSUBS 0.03154f
C417 VTAIL.n181 VSUBS 0.016948f
C418 VTAIL.n182 VSUBS 0.016948f
C419 VTAIL.n183 VSUBS 0.017945f
C420 VTAIL.n184 VSUBS 0.04006f
C421 VTAIL.n185 VSUBS 0.04006f
C422 VTAIL.n186 VSUBS 0.04006f
C423 VTAIL.n187 VSUBS 0.017447f
C424 VTAIL.n188 VSUBS 0.016948f
C425 VTAIL.n189 VSUBS 0.03154f
C426 VTAIL.n190 VSUBS 0.03154f
C427 VTAIL.n191 VSUBS 0.016948f
C428 VTAIL.n192 VSUBS 0.017945f
C429 VTAIL.n193 VSUBS 0.04006f
C430 VTAIL.n194 VSUBS 0.090156f
C431 VTAIL.n195 VSUBS 0.017945f
C432 VTAIL.n196 VSUBS 0.016948f
C433 VTAIL.n197 VSUBS 0.073766f
C434 VTAIL.n198 VSUBS 0.045062f
C435 VTAIL.n199 VSUBS 1.68287f
C436 VN.t1 VSUBS 3.75632f
C437 VN.t0 VSUBS 4.62488f
C438 B.n0 VSUBS 0.005587f
C439 B.n1 VSUBS 0.005587f
C440 B.n2 VSUBS 0.008263f
C441 B.n3 VSUBS 0.006332f
C442 B.n4 VSUBS 0.006332f
C443 B.n5 VSUBS 0.006332f
C444 B.n6 VSUBS 0.006332f
C445 B.n7 VSUBS 0.006332f
C446 B.n8 VSUBS 0.006332f
C447 B.n9 VSUBS 0.006332f
C448 B.n10 VSUBS 0.006332f
C449 B.n11 VSUBS 0.006332f
C450 B.n12 VSUBS 0.006332f
C451 B.n13 VSUBS 0.006332f
C452 B.n14 VSUBS 0.006332f
C453 B.n15 VSUBS 0.006332f
C454 B.n16 VSUBS 0.006332f
C455 B.n17 VSUBS 0.01568f
C456 B.n18 VSUBS 0.006332f
C457 B.n19 VSUBS 0.006332f
C458 B.n20 VSUBS 0.006332f
C459 B.n21 VSUBS 0.006332f
C460 B.n22 VSUBS 0.006332f
C461 B.n23 VSUBS 0.006332f
C462 B.n24 VSUBS 0.006332f
C463 B.n25 VSUBS 0.006332f
C464 B.n26 VSUBS 0.006332f
C465 B.n27 VSUBS 0.006332f
C466 B.n28 VSUBS 0.006332f
C467 B.n29 VSUBS 0.006332f
C468 B.n30 VSUBS 0.006332f
C469 B.n31 VSUBS 0.006332f
C470 B.n32 VSUBS 0.006332f
C471 B.n33 VSUBS 0.006332f
C472 B.t7 VSUBS 0.137412f
C473 B.t8 VSUBS 0.172076f
C474 B.t6 VSUBS 1.38737f
C475 B.n34 VSUBS 0.278484f
C476 B.n35 VSUBS 0.195123f
C477 B.n36 VSUBS 0.014671f
C478 B.n37 VSUBS 0.006332f
C479 B.n38 VSUBS 0.006332f
C480 B.n39 VSUBS 0.006332f
C481 B.n40 VSUBS 0.006332f
C482 B.n41 VSUBS 0.006332f
C483 B.t10 VSUBS 0.137415f
C484 B.t11 VSUBS 0.172078f
C485 B.t9 VSUBS 1.38737f
C486 B.n42 VSUBS 0.278482f
C487 B.n43 VSUBS 0.195121f
C488 B.n44 VSUBS 0.006332f
C489 B.n45 VSUBS 0.006332f
C490 B.n46 VSUBS 0.006332f
C491 B.n47 VSUBS 0.006332f
C492 B.n48 VSUBS 0.006332f
C493 B.n49 VSUBS 0.006332f
C494 B.n50 VSUBS 0.006332f
C495 B.n51 VSUBS 0.006332f
C496 B.n52 VSUBS 0.006332f
C497 B.n53 VSUBS 0.006332f
C498 B.n54 VSUBS 0.006332f
C499 B.n55 VSUBS 0.006332f
C500 B.n56 VSUBS 0.006332f
C501 B.n57 VSUBS 0.006332f
C502 B.n58 VSUBS 0.006332f
C503 B.n59 VSUBS 0.006332f
C504 B.n60 VSUBS 0.014491f
C505 B.n61 VSUBS 0.006332f
C506 B.n62 VSUBS 0.006332f
C507 B.n63 VSUBS 0.006332f
C508 B.n64 VSUBS 0.006332f
C509 B.n65 VSUBS 0.006332f
C510 B.n66 VSUBS 0.006332f
C511 B.n67 VSUBS 0.006332f
C512 B.n68 VSUBS 0.006332f
C513 B.n69 VSUBS 0.006332f
C514 B.n70 VSUBS 0.006332f
C515 B.n71 VSUBS 0.006332f
C516 B.n72 VSUBS 0.006332f
C517 B.n73 VSUBS 0.006332f
C518 B.n74 VSUBS 0.006332f
C519 B.n75 VSUBS 0.006332f
C520 B.n76 VSUBS 0.006332f
C521 B.n77 VSUBS 0.006332f
C522 B.n78 VSUBS 0.006332f
C523 B.n79 VSUBS 0.006332f
C524 B.n80 VSUBS 0.006332f
C525 B.n81 VSUBS 0.006332f
C526 B.n82 VSUBS 0.006332f
C527 B.n83 VSUBS 0.006332f
C528 B.n84 VSUBS 0.006332f
C529 B.n85 VSUBS 0.006332f
C530 B.n86 VSUBS 0.006332f
C531 B.n87 VSUBS 0.006332f
C532 B.n88 VSUBS 0.006332f
C533 B.n89 VSUBS 0.006332f
C534 B.n90 VSUBS 0.006332f
C535 B.n91 VSUBS 0.01568f
C536 B.n92 VSUBS 0.006332f
C537 B.n93 VSUBS 0.006332f
C538 B.n94 VSUBS 0.006332f
C539 B.n95 VSUBS 0.006332f
C540 B.n96 VSUBS 0.006332f
C541 B.n97 VSUBS 0.006332f
C542 B.n98 VSUBS 0.006332f
C543 B.n99 VSUBS 0.006332f
C544 B.n100 VSUBS 0.006332f
C545 B.n101 VSUBS 0.006332f
C546 B.n102 VSUBS 0.006332f
C547 B.n103 VSUBS 0.006332f
C548 B.n104 VSUBS 0.006332f
C549 B.n105 VSUBS 0.006332f
C550 B.n106 VSUBS 0.006332f
C551 B.n107 VSUBS 0.006332f
C552 B.t2 VSUBS 0.137415f
C553 B.t1 VSUBS 0.172078f
C554 B.t0 VSUBS 1.38737f
C555 B.n108 VSUBS 0.278482f
C556 B.n109 VSUBS 0.195121f
C557 B.n110 VSUBS 0.014671f
C558 B.n111 VSUBS 0.006332f
C559 B.n112 VSUBS 0.006332f
C560 B.n113 VSUBS 0.006332f
C561 B.n114 VSUBS 0.006332f
C562 B.n115 VSUBS 0.006332f
C563 B.t5 VSUBS 0.137412f
C564 B.t4 VSUBS 0.172076f
C565 B.t3 VSUBS 1.38737f
C566 B.n116 VSUBS 0.278484f
C567 B.n117 VSUBS 0.195123f
C568 B.n118 VSUBS 0.006332f
C569 B.n119 VSUBS 0.006332f
C570 B.n120 VSUBS 0.006332f
C571 B.n121 VSUBS 0.006332f
C572 B.n122 VSUBS 0.006332f
C573 B.n123 VSUBS 0.006332f
C574 B.n124 VSUBS 0.006332f
C575 B.n125 VSUBS 0.006332f
C576 B.n126 VSUBS 0.006332f
C577 B.n127 VSUBS 0.006332f
C578 B.n128 VSUBS 0.006332f
C579 B.n129 VSUBS 0.006332f
C580 B.n130 VSUBS 0.006332f
C581 B.n131 VSUBS 0.006332f
C582 B.n132 VSUBS 0.006332f
C583 B.n133 VSUBS 0.006332f
C584 B.n134 VSUBS 0.014491f
C585 B.n135 VSUBS 0.006332f
C586 B.n136 VSUBS 0.006332f
C587 B.n137 VSUBS 0.006332f
C588 B.n138 VSUBS 0.006332f
C589 B.n139 VSUBS 0.006332f
C590 B.n140 VSUBS 0.006332f
C591 B.n141 VSUBS 0.006332f
C592 B.n142 VSUBS 0.006332f
C593 B.n143 VSUBS 0.006332f
C594 B.n144 VSUBS 0.006332f
C595 B.n145 VSUBS 0.006332f
C596 B.n146 VSUBS 0.006332f
C597 B.n147 VSUBS 0.006332f
C598 B.n148 VSUBS 0.006332f
C599 B.n149 VSUBS 0.006332f
C600 B.n150 VSUBS 0.006332f
C601 B.n151 VSUBS 0.006332f
C602 B.n152 VSUBS 0.006332f
C603 B.n153 VSUBS 0.006332f
C604 B.n154 VSUBS 0.006332f
C605 B.n155 VSUBS 0.006332f
C606 B.n156 VSUBS 0.006332f
C607 B.n157 VSUBS 0.006332f
C608 B.n158 VSUBS 0.006332f
C609 B.n159 VSUBS 0.006332f
C610 B.n160 VSUBS 0.006332f
C611 B.n161 VSUBS 0.006332f
C612 B.n162 VSUBS 0.006332f
C613 B.n163 VSUBS 0.006332f
C614 B.n164 VSUBS 0.006332f
C615 B.n165 VSUBS 0.006332f
C616 B.n166 VSUBS 0.006332f
C617 B.n167 VSUBS 0.006332f
C618 B.n168 VSUBS 0.006332f
C619 B.n169 VSUBS 0.006332f
C620 B.n170 VSUBS 0.006332f
C621 B.n171 VSUBS 0.006332f
C622 B.n172 VSUBS 0.006332f
C623 B.n173 VSUBS 0.006332f
C624 B.n174 VSUBS 0.006332f
C625 B.n175 VSUBS 0.006332f
C626 B.n176 VSUBS 0.006332f
C627 B.n177 VSUBS 0.006332f
C628 B.n178 VSUBS 0.006332f
C629 B.n179 VSUBS 0.006332f
C630 B.n180 VSUBS 0.006332f
C631 B.n181 VSUBS 0.006332f
C632 B.n182 VSUBS 0.006332f
C633 B.n183 VSUBS 0.006332f
C634 B.n184 VSUBS 0.006332f
C635 B.n185 VSUBS 0.006332f
C636 B.n186 VSUBS 0.006332f
C637 B.n187 VSUBS 0.006332f
C638 B.n188 VSUBS 0.006332f
C639 B.n189 VSUBS 0.006332f
C640 B.n190 VSUBS 0.006332f
C641 B.n191 VSUBS 0.014491f
C642 B.n192 VSUBS 0.01568f
C643 B.n193 VSUBS 0.01568f
C644 B.n194 VSUBS 0.006332f
C645 B.n195 VSUBS 0.006332f
C646 B.n196 VSUBS 0.006332f
C647 B.n197 VSUBS 0.006332f
C648 B.n198 VSUBS 0.006332f
C649 B.n199 VSUBS 0.006332f
C650 B.n200 VSUBS 0.006332f
C651 B.n201 VSUBS 0.006332f
C652 B.n202 VSUBS 0.006332f
C653 B.n203 VSUBS 0.006332f
C654 B.n204 VSUBS 0.006332f
C655 B.n205 VSUBS 0.006332f
C656 B.n206 VSUBS 0.006332f
C657 B.n207 VSUBS 0.006332f
C658 B.n208 VSUBS 0.006332f
C659 B.n209 VSUBS 0.006332f
C660 B.n210 VSUBS 0.006332f
C661 B.n211 VSUBS 0.006332f
C662 B.n212 VSUBS 0.006332f
C663 B.n213 VSUBS 0.006332f
C664 B.n214 VSUBS 0.006332f
C665 B.n215 VSUBS 0.006332f
C666 B.n216 VSUBS 0.006332f
C667 B.n217 VSUBS 0.006332f
C668 B.n218 VSUBS 0.006332f
C669 B.n219 VSUBS 0.006332f
C670 B.n220 VSUBS 0.006332f
C671 B.n221 VSUBS 0.006332f
C672 B.n222 VSUBS 0.006332f
C673 B.n223 VSUBS 0.006332f
C674 B.n224 VSUBS 0.006332f
C675 B.n225 VSUBS 0.006332f
C676 B.n226 VSUBS 0.006332f
C677 B.n227 VSUBS 0.006332f
C678 B.n228 VSUBS 0.006332f
C679 B.n229 VSUBS 0.006332f
C680 B.n230 VSUBS 0.006332f
C681 B.n231 VSUBS 0.006332f
C682 B.n232 VSUBS 0.006332f
C683 B.n233 VSUBS 0.006332f
C684 B.n234 VSUBS 0.006332f
C685 B.n235 VSUBS 0.006332f
C686 B.n236 VSUBS 0.006332f
C687 B.n237 VSUBS 0.006332f
C688 B.n238 VSUBS 0.006332f
C689 B.n239 VSUBS 0.006332f
C690 B.n240 VSUBS 0.006332f
C691 B.n241 VSUBS 0.006332f
C692 B.n242 VSUBS 0.004377f
C693 B.n243 VSUBS 0.014671f
C694 B.n244 VSUBS 0.005122f
C695 B.n245 VSUBS 0.006332f
C696 B.n246 VSUBS 0.006332f
C697 B.n247 VSUBS 0.006332f
C698 B.n248 VSUBS 0.006332f
C699 B.n249 VSUBS 0.006332f
C700 B.n250 VSUBS 0.006332f
C701 B.n251 VSUBS 0.006332f
C702 B.n252 VSUBS 0.006332f
C703 B.n253 VSUBS 0.006332f
C704 B.n254 VSUBS 0.006332f
C705 B.n255 VSUBS 0.006332f
C706 B.n256 VSUBS 0.005122f
C707 B.n257 VSUBS 0.006332f
C708 B.n258 VSUBS 0.006332f
C709 B.n259 VSUBS 0.004377f
C710 B.n260 VSUBS 0.006332f
C711 B.n261 VSUBS 0.006332f
C712 B.n262 VSUBS 0.006332f
C713 B.n263 VSUBS 0.006332f
C714 B.n264 VSUBS 0.006332f
C715 B.n265 VSUBS 0.006332f
C716 B.n266 VSUBS 0.006332f
C717 B.n267 VSUBS 0.006332f
C718 B.n268 VSUBS 0.006332f
C719 B.n269 VSUBS 0.006332f
C720 B.n270 VSUBS 0.006332f
C721 B.n271 VSUBS 0.006332f
C722 B.n272 VSUBS 0.006332f
C723 B.n273 VSUBS 0.006332f
C724 B.n274 VSUBS 0.006332f
C725 B.n275 VSUBS 0.006332f
C726 B.n276 VSUBS 0.006332f
C727 B.n277 VSUBS 0.006332f
C728 B.n278 VSUBS 0.006332f
C729 B.n279 VSUBS 0.006332f
C730 B.n280 VSUBS 0.006332f
C731 B.n281 VSUBS 0.006332f
C732 B.n282 VSUBS 0.006332f
C733 B.n283 VSUBS 0.006332f
C734 B.n284 VSUBS 0.006332f
C735 B.n285 VSUBS 0.006332f
C736 B.n286 VSUBS 0.006332f
C737 B.n287 VSUBS 0.006332f
C738 B.n288 VSUBS 0.006332f
C739 B.n289 VSUBS 0.006332f
C740 B.n290 VSUBS 0.006332f
C741 B.n291 VSUBS 0.006332f
C742 B.n292 VSUBS 0.006332f
C743 B.n293 VSUBS 0.006332f
C744 B.n294 VSUBS 0.006332f
C745 B.n295 VSUBS 0.006332f
C746 B.n296 VSUBS 0.006332f
C747 B.n297 VSUBS 0.006332f
C748 B.n298 VSUBS 0.006332f
C749 B.n299 VSUBS 0.006332f
C750 B.n300 VSUBS 0.006332f
C751 B.n301 VSUBS 0.006332f
C752 B.n302 VSUBS 0.006332f
C753 B.n303 VSUBS 0.006332f
C754 B.n304 VSUBS 0.006332f
C755 B.n305 VSUBS 0.006332f
C756 B.n306 VSUBS 0.006332f
C757 B.n307 VSUBS 0.006332f
C758 B.n308 VSUBS 0.014952f
C759 B.n309 VSUBS 0.015219f
C760 B.n310 VSUBS 0.014491f
C761 B.n311 VSUBS 0.006332f
C762 B.n312 VSUBS 0.006332f
C763 B.n313 VSUBS 0.006332f
C764 B.n314 VSUBS 0.006332f
C765 B.n315 VSUBS 0.006332f
C766 B.n316 VSUBS 0.006332f
C767 B.n317 VSUBS 0.006332f
C768 B.n318 VSUBS 0.006332f
C769 B.n319 VSUBS 0.006332f
C770 B.n320 VSUBS 0.006332f
C771 B.n321 VSUBS 0.006332f
C772 B.n322 VSUBS 0.006332f
C773 B.n323 VSUBS 0.006332f
C774 B.n324 VSUBS 0.006332f
C775 B.n325 VSUBS 0.006332f
C776 B.n326 VSUBS 0.006332f
C777 B.n327 VSUBS 0.006332f
C778 B.n328 VSUBS 0.006332f
C779 B.n329 VSUBS 0.006332f
C780 B.n330 VSUBS 0.006332f
C781 B.n331 VSUBS 0.006332f
C782 B.n332 VSUBS 0.006332f
C783 B.n333 VSUBS 0.006332f
C784 B.n334 VSUBS 0.006332f
C785 B.n335 VSUBS 0.006332f
C786 B.n336 VSUBS 0.006332f
C787 B.n337 VSUBS 0.006332f
C788 B.n338 VSUBS 0.006332f
C789 B.n339 VSUBS 0.006332f
C790 B.n340 VSUBS 0.006332f
C791 B.n341 VSUBS 0.006332f
C792 B.n342 VSUBS 0.006332f
C793 B.n343 VSUBS 0.006332f
C794 B.n344 VSUBS 0.006332f
C795 B.n345 VSUBS 0.006332f
C796 B.n346 VSUBS 0.006332f
C797 B.n347 VSUBS 0.006332f
C798 B.n348 VSUBS 0.006332f
C799 B.n349 VSUBS 0.006332f
C800 B.n350 VSUBS 0.006332f
C801 B.n351 VSUBS 0.006332f
C802 B.n352 VSUBS 0.006332f
C803 B.n353 VSUBS 0.006332f
C804 B.n354 VSUBS 0.006332f
C805 B.n355 VSUBS 0.006332f
C806 B.n356 VSUBS 0.006332f
C807 B.n357 VSUBS 0.006332f
C808 B.n358 VSUBS 0.006332f
C809 B.n359 VSUBS 0.006332f
C810 B.n360 VSUBS 0.006332f
C811 B.n361 VSUBS 0.006332f
C812 B.n362 VSUBS 0.006332f
C813 B.n363 VSUBS 0.006332f
C814 B.n364 VSUBS 0.006332f
C815 B.n365 VSUBS 0.006332f
C816 B.n366 VSUBS 0.006332f
C817 B.n367 VSUBS 0.006332f
C818 B.n368 VSUBS 0.006332f
C819 B.n369 VSUBS 0.006332f
C820 B.n370 VSUBS 0.006332f
C821 B.n371 VSUBS 0.006332f
C822 B.n372 VSUBS 0.006332f
C823 B.n373 VSUBS 0.006332f
C824 B.n374 VSUBS 0.006332f
C825 B.n375 VSUBS 0.006332f
C826 B.n376 VSUBS 0.006332f
C827 B.n377 VSUBS 0.006332f
C828 B.n378 VSUBS 0.006332f
C829 B.n379 VSUBS 0.006332f
C830 B.n380 VSUBS 0.006332f
C831 B.n381 VSUBS 0.006332f
C832 B.n382 VSUBS 0.006332f
C833 B.n383 VSUBS 0.006332f
C834 B.n384 VSUBS 0.006332f
C835 B.n385 VSUBS 0.006332f
C836 B.n386 VSUBS 0.006332f
C837 B.n387 VSUBS 0.006332f
C838 B.n388 VSUBS 0.006332f
C839 B.n389 VSUBS 0.006332f
C840 B.n390 VSUBS 0.006332f
C841 B.n391 VSUBS 0.006332f
C842 B.n392 VSUBS 0.006332f
C843 B.n393 VSUBS 0.006332f
C844 B.n394 VSUBS 0.006332f
C845 B.n395 VSUBS 0.006332f
C846 B.n396 VSUBS 0.006332f
C847 B.n397 VSUBS 0.006332f
C848 B.n398 VSUBS 0.006332f
C849 B.n399 VSUBS 0.006332f
C850 B.n400 VSUBS 0.006332f
C851 B.n401 VSUBS 0.014491f
C852 B.n402 VSUBS 0.01568f
C853 B.n403 VSUBS 0.01568f
C854 B.n404 VSUBS 0.006332f
C855 B.n405 VSUBS 0.006332f
C856 B.n406 VSUBS 0.006332f
C857 B.n407 VSUBS 0.006332f
C858 B.n408 VSUBS 0.006332f
C859 B.n409 VSUBS 0.006332f
C860 B.n410 VSUBS 0.006332f
C861 B.n411 VSUBS 0.006332f
C862 B.n412 VSUBS 0.006332f
C863 B.n413 VSUBS 0.006332f
C864 B.n414 VSUBS 0.006332f
C865 B.n415 VSUBS 0.006332f
C866 B.n416 VSUBS 0.006332f
C867 B.n417 VSUBS 0.006332f
C868 B.n418 VSUBS 0.006332f
C869 B.n419 VSUBS 0.006332f
C870 B.n420 VSUBS 0.006332f
C871 B.n421 VSUBS 0.006332f
C872 B.n422 VSUBS 0.006332f
C873 B.n423 VSUBS 0.006332f
C874 B.n424 VSUBS 0.006332f
C875 B.n425 VSUBS 0.006332f
C876 B.n426 VSUBS 0.006332f
C877 B.n427 VSUBS 0.006332f
C878 B.n428 VSUBS 0.006332f
C879 B.n429 VSUBS 0.006332f
C880 B.n430 VSUBS 0.006332f
C881 B.n431 VSUBS 0.006332f
C882 B.n432 VSUBS 0.006332f
C883 B.n433 VSUBS 0.006332f
C884 B.n434 VSUBS 0.006332f
C885 B.n435 VSUBS 0.006332f
C886 B.n436 VSUBS 0.006332f
C887 B.n437 VSUBS 0.006332f
C888 B.n438 VSUBS 0.006332f
C889 B.n439 VSUBS 0.006332f
C890 B.n440 VSUBS 0.006332f
C891 B.n441 VSUBS 0.006332f
C892 B.n442 VSUBS 0.006332f
C893 B.n443 VSUBS 0.006332f
C894 B.n444 VSUBS 0.006332f
C895 B.n445 VSUBS 0.006332f
C896 B.n446 VSUBS 0.006332f
C897 B.n447 VSUBS 0.006332f
C898 B.n448 VSUBS 0.006332f
C899 B.n449 VSUBS 0.006332f
C900 B.n450 VSUBS 0.006332f
C901 B.n451 VSUBS 0.006332f
C902 B.n452 VSUBS 0.004377f
C903 B.n453 VSUBS 0.014671f
C904 B.n454 VSUBS 0.005122f
C905 B.n455 VSUBS 0.006332f
C906 B.n456 VSUBS 0.006332f
C907 B.n457 VSUBS 0.006332f
C908 B.n458 VSUBS 0.006332f
C909 B.n459 VSUBS 0.006332f
C910 B.n460 VSUBS 0.006332f
C911 B.n461 VSUBS 0.006332f
C912 B.n462 VSUBS 0.006332f
C913 B.n463 VSUBS 0.006332f
C914 B.n464 VSUBS 0.006332f
C915 B.n465 VSUBS 0.006332f
C916 B.n466 VSUBS 0.005122f
C917 B.n467 VSUBS 0.006332f
C918 B.n468 VSUBS 0.006332f
C919 B.n469 VSUBS 0.004377f
C920 B.n470 VSUBS 0.006332f
C921 B.n471 VSUBS 0.006332f
C922 B.n472 VSUBS 0.006332f
C923 B.n473 VSUBS 0.006332f
C924 B.n474 VSUBS 0.006332f
C925 B.n475 VSUBS 0.006332f
C926 B.n476 VSUBS 0.006332f
C927 B.n477 VSUBS 0.006332f
C928 B.n478 VSUBS 0.006332f
C929 B.n479 VSUBS 0.006332f
C930 B.n480 VSUBS 0.006332f
C931 B.n481 VSUBS 0.006332f
C932 B.n482 VSUBS 0.006332f
C933 B.n483 VSUBS 0.006332f
C934 B.n484 VSUBS 0.006332f
C935 B.n485 VSUBS 0.006332f
C936 B.n486 VSUBS 0.006332f
C937 B.n487 VSUBS 0.006332f
C938 B.n488 VSUBS 0.006332f
C939 B.n489 VSUBS 0.006332f
C940 B.n490 VSUBS 0.006332f
C941 B.n491 VSUBS 0.006332f
C942 B.n492 VSUBS 0.006332f
C943 B.n493 VSUBS 0.006332f
C944 B.n494 VSUBS 0.006332f
C945 B.n495 VSUBS 0.006332f
C946 B.n496 VSUBS 0.006332f
C947 B.n497 VSUBS 0.006332f
C948 B.n498 VSUBS 0.006332f
C949 B.n499 VSUBS 0.006332f
C950 B.n500 VSUBS 0.006332f
C951 B.n501 VSUBS 0.006332f
C952 B.n502 VSUBS 0.006332f
C953 B.n503 VSUBS 0.006332f
C954 B.n504 VSUBS 0.006332f
C955 B.n505 VSUBS 0.006332f
C956 B.n506 VSUBS 0.006332f
C957 B.n507 VSUBS 0.006332f
C958 B.n508 VSUBS 0.006332f
C959 B.n509 VSUBS 0.006332f
C960 B.n510 VSUBS 0.006332f
C961 B.n511 VSUBS 0.006332f
C962 B.n512 VSUBS 0.006332f
C963 B.n513 VSUBS 0.006332f
C964 B.n514 VSUBS 0.006332f
C965 B.n515 VSUBS 0.006332f
C966 B.n516 VSUBS 0.006332f
C967 B.n517 VSUBS 0.006332f
C968 B.n518 VSUBS 0.01568f
C969 B.n519 VSUBS 0.014491f
C970 B.n520 VSUBS 0.014491f
C971 B.n521 VSUBS 0.006332f
C972 B.n522 VSUBS 0.006332f
C973 B.n523 VSUBS 0.006332f
C974 B.n524 VSUBS 0.006332f
C975 B.n525 VSUBS 0.006332f
C976 B.n526 VSUBS 0.006332f
C977 B.n527 VSUBS 0.006332f
C978 B.n528 VSUBS 0.006332f
C979 B.n529 VSUBS 0.006332f
C980 B.n530 VSUBS 0.006332f
C981 B.n531 VSUBS 0.006332f
C982 B.n532 VSUBS 0.006332f
C983 B.n533 VSUBS 0.006332f
C984 B.n534 VSUBS 0.006332f
C985 B.n535 VSUBS 0.006332f
C986 B.n536 VSUBS 0.006332f
C987 B.n537 VSUBS 0.006332f
C988 B.n538 VSUBS 0.006332f
C989 B.n539 VSUBS 0.006332f
C990 B.n540 VSUBS 0.006332f
C991 B.n541 VSUBS 0.006332f
C992 B.n542 VSUBS 0.006332f
C993 B.n543 VSUBS 0.006332f
C994 B.n544 VSUBS 0.006332f
C995 B.n545 VSUBS 0.006332f
C996 B.n546 VSUBS 0.006332f
C997 B.n547 VSUBS 0.006332f
C998 B.n548 VSUBS 0.006332f
C999 B.n549 VSUBS 0.006332f
C1000 B.n550 VSUBS 0.006332f
C1001 B.n551 VSUBS 0.006332f
C1002 B.n552 VSUBS 0.006332f
C1003 B.n553 VSUBS 0.006332f
C1004 B.n554 VSUBS 0.006332f
C1005 B.n555 VSUBS 0.006332f
C1006 B.n556 VSUBS 0.006332f
C1007 B.n557 VSUBS 0.006332f
C1008 B.n558 VSUBS 0.006332f
C1009 B.n559 VSUBS 0.006332f
C1010 B.n560 VSUBS 0.006332f
C1011 B.n561 VSUBS 0.006332f
C1012 B.n562 VSUBS 0.006332f
C1013 B.n563 VSUBS 0.008263f
C1014 B.n564 VSUBS 0.008802f
C1015 B.n565 VSUBS 0.017504f
.ends

