* NGSPICE file created from diff_pair_sample_0543.ext - technology: sky130A

.subckt diff_pair_sample_0543 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.38
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.38
X2 VTAIL.t2 VP.t1 VDD1.t4 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.38
X3 VTAIL.t11 VN.t1 VDD2.t4 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.38
X4 B.t11 B.t9 B.t10 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.38
X5 VDD2.t3 VN.t2 VTAIL.t10 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.38
X6 VDD2.t2 VN.t3 VTAIL.t7 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.38
X7 VDD1.t3 VP.t2 VTAIL.t4 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.38
X8 VDD2.t1 VN.t4 VTAIL.t8 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.38
X9 B.t8 B.t6 B.t7 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.38
X10 VDD1.t2 VP.t3 VTAIL.t0 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.38
X11 VTAIL.t9 VN.t5 VDD2.t0 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.38
X12 VTAIL.t1 VP.t4 VDD1.t1 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.38
X13 B.t5 B.t3 B.t4 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.38
X14 VDD1.t0 VP.t5 VTAIL.t3 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.38
X15 B.t2 B.t0 B.t1 w_n3938_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.38
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n17 VN.n0 79.7913
R15 VN.n35 VN.n18 79.7913
R16 VN.n23 VN.t3 68.3414
R17 VN.n5 VN.t4 68.3414
R18 VN.n9 VN.n2 54.5767
R19 VN.n27 VN.n20 54.5767
R20 VN.n5 VN.n4 50.1196
R21 VN.n23 VN.n22 50.1196
R22 VN VN.n35 46.5776
R23 VN.n4 VN.t1 34.8671
R24 VN.n0 VN.t0 34.8671
R25 VN.n22 VN.t5 34.8671
R26 VN.n18 VN.t2 34.8671
R27 VN.n13 VN.n2 26.41
R28 VN.n31 VN.n20 26.41
R29 VN.n7 VN.n4 24.4675
R30 VN.n8 VN.n7 24.4675
R31 VN.n9 VN.n8 24.4675
R32 VN.n14 VN.n13 24.4675
R33 VN.n15 VN.n14 24.4675
R34 VN.n27 VN.n26 24.4675
R35 VN.n26 VN.n25 24.4675
R36 VN.n25 VN.n22 24.4675
R37 VN.n33 VN.n32 24.4675
R38 VN.n32 VN.n31 24.4675
R39 VN.n15 VN.n0 10.2766
R40 VN.n33 VN.n18 10.2766
R41 VN.n24 VN.n23 3.14396
R42 VN.n6 VN.n5 3.14396
R43 VN.n35 VN.n34 0.354971
R44 VN.n17 VN.n16 0.354971
R45 VN VN.n17 0.26696
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VTAIL.n7 VTAIL.t7 89.8274
R59 VTAIL.n11 VTAIL.t6 89.8273
R60 VTAIL.n2 VTAIL.t3 89.8273
R61 VTAIL.n10 VTAIL.t4 89.8273
R62 VTAIL.n9 VTAIL.n8 83.1802
R63 VTAIL.n6 VTAIL.n5 83.1802
R64 VTAIL.n1 VTAIL.n0 83.18
R65 VTAIL.n4 VTAIL.n3 83.18
R66 VTAIL.n6 VTAIL.n4 22.9789
R67 VTAIL.n11 VTAIL.n10 19.7807
R68 VTAIL.n0 VTAIL.t8 6.64774
R69 VTAIL.n0 VTAIL.t11 6.64774
R70 VTAIL.n3 VTAIL.t0 6.64774
R71 VTAIL.n3 VTAIL.t1 6.64774
R72 VTAIL.n8 VTAIL.t5 6.64774
R73 VTAIL.n8 VTAIL.t2 6.64774
R74 VTAIL.n5 VTAIL.t10 6.64774
R75 VTAIL.n5 VTAIL.t9 6.64774
R76 VTAIL.n7 VTAIL.n6 3.19878
R77 VTAIL.n10 VTAIL.n9 3.19878
R78 VTAIL.n4 VTAIL.n2 3.19878
R79 VTAIL VTAIL.n11 2.34102
R80 VTAIL.n9 VTAIL.n7 2.06947
R81 VTAIL.n2 VTAIL.n1 2.06947
R82 VTAIL VTAIL.n1 0.858259
R83 VDD2.n1 VDD2.t1 108.85
R84 VDD2.n2 VDD2.t3 106.507
R85 VDD2.n1 VDD2.n0 100.603
R86 VDD2 VDD2.n3 100.6
R87 VDD2.n2 VDD2.n1 38.3252
R88 VDD2.n3 VDD2.t0 6.64774
R89 VDD2.n3 VDD2.t2 6.64774
R90 VDD2.n0 VDD2.t4 6.64774
R91 VDD2.n0 VDD2.t5 6.64774
R92 VDD2 VDD2.n2 2.4574
R93 VP.n16 VP.n15 161.3
R94 VP.n17 VP.n12 161.3
R95 VP.n19 VP.n18 161.3
R96 VP.n20 VP.n11 161.3
R97 VP.n22 VP.n21 161.3
R98 VP.n23 VP.n10 161.3
R99 VP.n25 VP.n24 161.3
R100 VP.n50 VP.n49 161.3
R101 VP.n48 VP.n1 161.3
R102 VP.n47 VP.n46 161.3
R103 VP.n45 VP.n2 161.3
R104 VP.n44 VP.n43 161.3
R105 VP.n42 VP.n3 161.3
R106 VP.n41 VP.n40 161.3
R107 VP.n39 VP.n4 161.3
R108 VP.n38 VP.n37 161.3
R109 VP.n36 VP.n5 161.3
R110 VP.n35 VP.n34 161.3
R111 VP.n33 VP.n6 161.3
R112 VP.n32 VP.n31 161.3
R113 VP.n30 VP.n7 161.3
R114 VP.n29 VP.n28 161.3
R115 VP.n27 VP.n8 79.7913
R116 VP.n51 VP.n0 79.7913
R117 VP.n26 VP.n9 79.7913
R118 VP.n14 VP.t0 68.3412
R119 VP.n35 VP.n6 54.5767
R120 VP.n43 VP.n2 54.5767
R121 VP.n18 VP.n11 54.5767
R122 VP.n14 VP.n13 50.1196
R123 VP.n27 VP.n26 46.4122
R124 VP.n4 VP.t4 34.8671
R125 VP.n8 VP.t3 34.8671
R126 VP.n0 VP.t5 34.8671
R127 VP.n13 VP.t1 34.8671
R128 VP.n9 VP.t2 34.8671
R129 VP.n31 VP.n6 26.41
R130 VP.n47 VP.n2 26.41
R131 VP.n22 VP.n11 26.41
R132 VP.n30 VP.n29 24.4675
R133 VP.n31 VP.n30 24.4675
R134 VP.n36 VP.n35 24.4675
R135 VP.n37 VP.n36 24.4675
R136 VP.n37 VP.n4 24.4675
R137 VP.n41 VP.n4 24.4675
R138 VP.n42 VP.n41 24.4675
R139 VP.n43 VP.n42 24.4675
R140 VP.n48 VP.n47 24.4675
R141 VP.n49 VP.n48 24.4675
R142 VP.n23 VP.n22 24.4675
R143 VP.n24 VP.n23 24.4675
R144 VP.n16 VP.n13 24.4675
R145 VP.n17 VP.n16 24.4675
R146 VP.n18 VP.n17 24.4675
R147 VP.n29 VP.n8 10.2766
R148 VP.n49 VP.n0 10.2766
R149 VP.n24 VP.n9 10.2766
R150 VP.n15 VP.n14 3.14395
R151 VP.n26 VP.n25 0.354971
R152 VP.n28 VP.n27 0.354971
R153 VP.n51 VP.n50 0.354971
R154 VP VP.n51 0.26696
R155 VP.n15 VP.n12 0.189894
R156 VP.n19 VP.n12 0.189894
R157 VP.n20 VP.n19 0.189894
R158 VP.n21 VP.n20 0.189894
R159 VP.n21 VP.n10 0.189894
R160 VP.n25 VP.n10 0.189894
R161 VP.n28 VP.n7 0.189894
R162 VP.n32 VP.n7 0.189894
R163 VP.n33 VP.n32 0.189894
R164 VP.n34 VP.n33 0.189894
R165 VP.n34 VP.n5 0.189894
R166 VP.n38 VP.n5 0.189894
R167 VP.n39 VP.n38 0.189894
R168 VP.n40 VP.n39 0.189894
R169 VP.n40 VP.n3 0.189894
R170 VP.n44 VP.n3 0.189894
R171 VP.n45 VP.n44 0.189894
R172 VP.n46 VP.n45 0.189894
R173 VP.n46 VP.n1 0.189894
R174 VP.n50 VP.n1 0.189894
R175 VDD1 VDD1.t5 108.963
R176 VDD1.n1 VDD1.t2 108.85
R177 VDD1.n1 VDD1.n0 100.603
R178 VDD1.n3 VDD1.n2 99.8588
R179 VDD1.n3 VDD1.n1 40.5074
R180 VDD1.n2 VDD1.t4 6.64774
R181 VDD1.n2 VDD1.t3 6.64774
R182 VDD1.n0 VDD1.t1 6.64774
R183 VDD1.n0 VDD1.t0 6.64774
R184 VDD1 VDD1.n3 0.741879
R185 B.n317 B.n316 585
R186 B.n315 B.n110 585
R187 B.n314 B.n313 585
R188 B.n312 B.n111 585
R189 B.n311 B.n310 585
R190 B.n309 B.n112 585
R191 B.n308 B.n307 585
R192 B.n306 B.n113 585
R193 B.n305 B.n304 585
R194 B.n303 B.n114 585
R195 B.n302 B.n301 585
R196 B.n300 B.n115 585
R197 B.n299 B.n298 585
R198 B.n297 B.n116 585
R199 B.n296 B.n295 585
R200 B.n294 B.n117 585
R201 B.n293 B.n292 585
R202 B.n291 B.n118 585
R203 B.n290 B.n289 585
R204 B.n288 B.n119 585
R205 B.n287 B.n286 585
R206 B.n285 B.n284 585
R207 B.n283 B.n123 585
R208 B.n282 B.n281 585
R209 B.n280 B.n124 585
R210 B.n279 B.n278 585
R211 B.n277 B.n125 585
R212 B.n276 B.n275 585
R213 B.n274 B.n126 585
R214 B.n273 B.n272 585
R215 B.n270 B.n127 585
R216 B.n269 B.n268 585
R217 B.n267 B.n130 585
R218 B.n266 B.n265 585
R219 B.n264 B.n131 585
R220 B.n263 B.n262 585
R221 B.n261 B.n132 585
R222 B.n260 B.n259 585
R223 B.n258 B.n133 585
R224 B.n257 B.n256 585
R225 B.n255 B.n134 585
R226 B.n254 B.n253 585
R227 B.n252 B.n135 585
R228 B.n251 B.n250 585
R229 B.n249 B.n136 585
R230 B.n248 B.n247 585
R231 B.n246 B.n137 585
R232 B.n245 B.n244 585
R233 B.n243 B.n138 585
R234 B.n242 B.n241 585
R235 B.n240 B.n139 585
R236 B.n318 B.n109 585
R237 B.n320 B.n319 585
R238 B.n321 B.n108 585
R239 B.n323 B.n322 585
R240 B.n324 B.n107 585
R241 B.n326 B.n325 585
R242 B.n327 B.n106 585
R243 B.n329 B.n328 585
R244 B.n330 B.n105 585
R245 B.n332 B.n331 585
R246 B.n333 B.n104 585
R247 B.n335 B.n334 585
R248 B.n336 B.n103 585
R249 B.n338 B.n337 585
R250 B.n339 B.n102 585
R251 B.n341 B.n340 585
R252 B.n342 B.n101 585
R253 B.n344 B.n343 585
R254 B.n345 B.n100 585
R255 B.n347 B.n346 585
R256 B.n348 B.n99 585
R257 B.n350 B.n349 585
R258 B.n351 B.n98 585
R259 B.n353 B.n352 585
R260 B.n354 B.n97 585
R261 B.n356 B.n355 585
R262 B.n357 B.n96 585
R263 B.n359 B.n358 585
R264 B.n360 B.n95 585
R265 B.n362 B.n361 585
R266 B.n363 B.n94 585
R267 B.n365 B.n364 585
R268 B.n366 B.n93 585
R269 B.n368 B.n367 585
R270 B.n369 B.n92 585
R271 B.n371 B.n370 585
R272 B.n372 B.n91 585
R273 B.n374 B.n373 585
R274 B.n375 B.n90 585
R275 B.n377 B.n376 585
R276 B.n378 B.n89 585
R277 B.n380 B.n379 585
R278 B.n381 B.n88 585
R279 B.n383 B.n382 585
R280 B.n384 B.n87 585
R281 B.n386 B.n385 585
R282 B.n387 B.n86 585
R283 B.n389 B.n388 585
R284 B.n390 B.n85 585
R285 B.n392 B.n391 585
R286 B.n393 B.n84 585
R287 B.n395 B.n394 585
R288 B.n396 B.n83 585
R289 B.n398 B.n397 585
R290 B.n399 B.n82 585
R291 B.n401 B.n400 585
R292 B.n402 B.n81 585
R293 B.n404 B.n403 585
R294 B.n405 B.n80 585
R295 B.n407 B.n406 585
R296 B.n408 B.n79 585
R297 B.n410 B.n409 585
R298 B.n411 B.n78 585
R299 B.n413 B.n412 585
R300 B.n414 B.n77 585
R301 B.n416 B.n415 585
R302 B.n417 B.n76 585
R303 B.n419 B.n418 585
R304 B.n420 B.n75 585
R305 B.n422 B.n421 585
R306 B.n423 B.n74 585
R307 B.n425 B.n424 585
R308 B.n426 B.n73 585
R309 B.n428 B.n427 585
R310 B.n429 B.n72 585
R311 B.n431 B.n430 585
R312 B.n432 B.n71 585
R313 B.n434 B.n433 585
R314 B.n435 B.n70 585
R315 B.n437 B.n436 585
R316 B.n438 B.n69 585
R317 B.n440 B.n439 585
R318 B.n441 B.n68 585
R319 B.n443 B.n442 585
R320 B.n444 B.n67 585
R321 B.n446 B.n445 585
R322 B.n447 B.n66 585
R323 B.n449 B.n448 585
R324 B.n450 B.n65 585
R325 B.n452 B.n451 585
R326 B.n453 B.n64 585
R327 B.n455 B.n454 585
R328 B.n456 B.n63 585
R329 B.n458 B.n457 585
R330 B.n459 B.n62 585
R331 B.n461 B.n460 585
R332 B.n462 B.n61 585
R333 B.n464 B.n463 585
R334 B.n465 B.n60 585
R335 B.n467 B.n466 585
R336 B.n468 B.n59 585
R337 B.n470 B.n469 585
R338 B.n471 B.n58 585
R339 B.n473 B.n472 585
R340 B.n551 B.n550 585
R341 B.n549 B.n28 585
R342 B.n548 B.n547 585
R343 B.n546 B.n29 585
R344 B.n545 B.n544 585
R345 B.n543 B.n30 585
R346 B.n542 B.n541 585
R347 B.n540 B.n31 585
R348 B.n539 B.n538 585
R349 B.n537 B.n32 585
R350 B.n536 B.n535 585
R351 B.n534 B.n33 585
R352 B.n533 B.n532 585
R353 B.n531 B.n34 585
R354 B.n530 B.n529 585
R355 B.n528 B.n35 585
R356 B.n527 B.n526 585
R357 B.n525 B.n36 585
R358 B.n524 B.n523 585
R359 B.n522 B.n37 585
R360 B.n521 B.n520 585
R361 B.n519 B.n518 585
R362 B.n517 B.n41 585
R363 B.n516 B.n515 585
R364 B.n514 B.n42 585
R365 B.n513 B.n512 585
R366 B.n511 B.n43 585
R367 B.n510 B.n509 585
R368 B.n508 B.n44 585
R369 B.n507 B.n506 585
R370 B.n504 B.n45 585
R371 B.n503 B.n502 585
R372 B.n501 B.n48 585
R373 B.n500 B.n499 585
R374 B.n498 B.n49 585
R375 B.n497 B.n496 585
R376 B.n495 B.n50 585
R377 B.n494 B.n493 585
R378 B.n492 B.n51 585
R379 B.n491 B.n490 585
R380 B.n489 B.n52 585
R381 B.n488 B.n487 585
R382 B.n486 B.n53 585
R383 B.n485 B.n484 585
R384 B.n483 B.n54 585
R385 B.n482 B.n481 585
R386 B.n480 B.n55 585
R387 B.n479 B.n478 585
R388 B.n477 B.n56 585
R389 B.n476 B.n475 585
R390 B.n474 B.n57 585
R391 B.n552 B.n27 585
R392 B.n554 B.n553 585
R393 B.n555 B.n26 585
R394 B.n557 B.n556 585
R395 B.n558 B.n25 585
R396 B.n560 B.n559 585
R397 B.n561 B.n24 585
R398 B.n563 B.n562 585
R399 B.n564 B.n23 585
R400 B.n566 B.n565 585
R401 B.n567 B.n22 585
R402 B.n569 B.n568 585
R403 B.n570 B.n21 585
R404 B.n572 B.n571 585
R405 B.n573 B.n20 585
R406 B.n575 B.n574 585
R407 B.n576 B.n19 585
R408 B.n578 B.n577 585
R409 B.n579 B.n18 585
R410 B.n581 B.n580 585
R411 B.n582 B.n17 585
R412 B.n584 B.n583 585
R413 B.n585 B.n16 585
R414 B.n587 B.n586 585
R415 B.n588 B.n15 585
R416 B.n590 B.n589 585
R417 B.n591 B.n14 585
R418 B.n593 B.n592 585
R419 B.n594 B.n13 585
R420 B.n596 B.n595 585
R421 B.n597 B.n12 585
R422 B.n599 B.n598 585
R423 B.n600 B.n11 585
R424 B.n602 B.n601 585
R425 B.n603 B.n10 585
R426 B.n605 B.n604 585
R427 B.n606 B.n9 585
R428 B.n608 B.n607 585
R429 B.n609 B.n8 585
R430 B.n611 B.n610 585
R431 B.n612 B.n7 585
R432 B.n614 B.n613 585
R433 B.n615 B.n6 585
R434 B.n617 B.n616 585
R435 B.n618 B.n5 585
R436 B.n620 B.n619 585
R437 B.n621 B.n4 585
R438 B.n623 B.n622 585
R439 B.n624 B.n3 585
R440 B.n626 B.n625 585
R441 B.n627 B.n0 585
R442 B.n2 B.n1 585
R443 B.n165 B.n164 585
R444 B.n167 B.n166 585
R445 B.n168 B.n163 585
R446 B.n170 B.n169 585
R447 B.n171 B.n162 585
R448 B.n173 B.n172 585
R449 B.n174 B.n161 585
R450 B.n176 B.n175 585
R451 B.n177 B.n160 585
R452 B.n179 B.n178 585
R453 B.n180 B.n159 585
R454 B.n182 B.n181 585
R455 B.n183 B.n158 585
R456 B.n185 B.n184 585
R457 B.n186 B.n157 585
R458 B.n188 B.n187 585
R459 B.n189 B.n156 585
R460 B.n191 B.n190 585
R461 B.n192 B.n155 585
R462 B.n194 B.n193 585
R463 B.n195 B.n154 585
R464 B.n197 B.n196 585
R465 B.n198 B.n153 585
R466 B.n200 B.n199 585
R467 B.n201 B.n152 585
R468 B.n203 B.n202 585
R469 B.n204 B.n151 585
R470 B.n206 B.n205 585
R471 B.n207 B.n150 585
R472 B.n209 B.n208 585
R473 B.n210 B.n149 585
R474 B.n212 B.n211 585
R475 B.n213 B.n148 585
R476 B.n215 B.n214 585
R477 B.n216 B.n147 585
R478 B.n218 B.n217 585
R479 B.n219 B.n146 585
R480 B.n221 B.n220 585
R481 B.n222 B.n145 585
R482 B.n224 B.n223 585
R483 B.n225 B.n144 585
R484 B.n227 B.n226 585
R485 B.n228 B.n143 585
R486 B.n230 B.n229 585
R487 B.n231 B.n142 585
R488 B.n233 B.n232 585
R489 B.n234 B.n141 585
R490 B.n236 B.n235 585
R491 B.n237 B.n140 585
R492 B.n239 B.n238 585
R493 B.n238 B.n139 540.549
R494 B.n316 B.n109 540.549
R495 B.n472 B.n57 540.549
R496 B.n550 B.n27 540.549
R497 B.n629 B.n628 256.663
R498 B.n128 B.t0 243.85
R499 B.n120 B.t6 243.85
R500 B.n46 B.t9 243.85
R501 B.n38 B.t3 243.85
R502 B.n628 B.n627 235.042
R503 B.n628 B.n2 235.042
R504 B.n120 B.t7 189.138
R505 B.n46 B.t11 189.138
R506 B.n128 B.t1 189.133
R507 B.n38 B.t5 189.133
R508 B.n242 B.n139 163.367
R509 B.n243 B.n242 163.367
R510 B.n244 B.n243 163.367
R511 B.n244 B.n137 163.367
R512 B.n248 B.n137 163.367
R513 B.n249 B.n248 163.367
R514 B.n250 B.n249 163.367
R515 B.n250 B.n135 163.367
R516 B.n254 B.n135 163.367
R517 B.n255 B.n254 163.367
R518 B.n256 B.n255 163.367
R519 B.n256 B.n133 163.367
R520 B.n260 B.n133 163.367
R521 B.n261 B.n260 163.367
R522 B.n262 B.n261 163.367
R523 B.n262 B.n131 163.367
R524 B.n266 B.n131 163.367
R525 B.n267 B.n266 163.367
R526 B.n268 B.n267 163.367
R527 B.n268 B.n127 163.367
R528 B.n273 B.n127 163.367
R529 B.n274 B.n273 163.367
R530 B.n275 B.n274 163.367
R531 B.n275 B.n125 163.367
R532 B.n279 B.n125 163.367
R533 B.n280 B.n279 163.367
R534 B.n281 B.n280 163.367
R535 B.n281 B.n123 163.367
R536 B.n285 B.n123 163.367
R537 B.n286 B.n285 163.367
R538 B.n286 B.n119 163.367
R539 B.n290 B.n119 163.367
R540 B.n291 B.n290 163.367
R541 B.n292 B.n291 163.367
R542 B.n292 B.n117 163.367
R543 B.n296 B.n117 163.367
R544 B.n297 B.n296 163.367
R545 B.n298 B.n297 163.367
R546 B.n298 B.n115 163.367
R547 B.n302 B.n115 163.367
R548 B.n303 B.n302 163.367
R549 B.n304 B.n303 163.367
R550 B.n304 B.n113 163.367
R551 B.n308 B.n113 163.367
R552 B.n309 B.n308 163.367
R553 B.n310 B.n309 163.367
R554 B.n310 B.n111 163.367
R555 B.n314 B.n111 163.367
R556 B.n315 B.n314 163.367
R557 B.n316 B.n315 163.367
R558 B.n472 B.n471 163.367
R559 B.n471 B.n470 163.367
R560 B.n470 B.n59 163.367
R561 B.n466 B.n59 163.367
R562 B.n466 B.n465 163.367
R563 B.n465 B.n464 163.367
R564 B.n464 B.n61 163.367
R565 B.n460 B.n61 163.367
R566 B.n460 B.n459 163.367
R567 B.n459 B.n458 163.367
R568 B.n458 B.n63 163.367
R569 B.n454 B.n63 163.367
R570 B.n454 B.n453 163.367
R571 B.n453 B.n452 163.367
R572 B.n452 B.n65 163.367
R573 B.n448 B.n65 163.367
R574 B.n448 B.n447 163.367
R575 B.n447 B.n446 163.367
R576 B.n446 B.n67 163.367
R577 B.n442 B.n67 163.367
R578 B.n442 B.n441 163.367
R579 B.n441 B.n440 163.367
R580 B.n440 B.n69 163.367
R581 B.n436 B.n69 163.367
R582 B.n436 B.n435 163.367
R583 B.n435 B.n434 163.367
R584 B.n434 B.n71 163.367
R585 B.n430 B.n71 163.367
R586 B.n430 B.n429 163.367
R587 B.n429 B.n428 163.367
R588 B.n428 B.n73 163.367
R589 B.n424 B.n73 163.367
R590 B.n424 B.n423 163.367
R591 B.n423 B.n422 163.367
R592 B.n422 B.n75 163.367
R593 B.n418 B.n75 163.367
R594 B.n418 B.n417 163.367
R595 B.n417 B.n416 163.367
R596 B.n416 B.n77 163.367
R597 B.n412 B.n77 163.367
R598 B.n412 B.n411 163.367
R599 B.n411 B.n410 163.367
R600 B.n410 B.n79 163.367
R601 B.n406 B.n79 163.367
R602 B.n406 B.n405 163.367
R603 B.n405 B.n404 163.367
R604 B.n404 B.n81 163.367
R605 B.n400 B.n81 163.367
R606 B.n400 B.n399 163.367
R607 B.n399 B.n398 163.367
R608 B.n398 B.n83 163.367
R609 B.n394 B.n83 163.367
R610 B.n394 B.n393 163.367
R611 B.n393 B.n392 163.367
R612 B.n392 B.n85 163.367
R613 B.n388 B.n85 163.367
R614 B.n388 B.n387 163.367
R615 B.n387 B.n386 163.367
R616 B.n386 B.n87 163.367
R617 B.n382 B.n87 163.367
R618 B.n382 B.n381 163.367
R619 B.n381 B.n380 163.367
R620 B.n380 B.n89 163.367
R621 B.n376 B.n89 163.367
R622 B.n376 B.n375 163.367
R623 B.n375 B.n374 163.367
R624 B.n374 B.n91 163.367
R625 B.n370 B.n91 163.367
R626 B.n370 B.n369 163.367
R627 B.n369 B.n368 163.367
R628 B.n368 B.n93 163.367
R629 B.n364 B.n93 163.367
R630 B.n364 B.n363 163.367
R631 B.n363 B.n362 163.367
R632 B.n362 B.n95 163.367
R633 B.n358 B.n95 163.367
R634 B.n358 B.n357 163.367
R635 B.n357 B.n356 163.367
R636 B.n356 B.n97 163.367
R637 B.n352 B.n97 163.367
R638 B.n352 B.n351 163.367
R639 B.n351 B.n350 163.367
R640 B.n350 B.n99 163.367
R641 B.n346 B.n99 163.367
R642 B.n346 B.n345 163.367
R643 B.n345 B.n344 163.367
R644 B.n344 B.n101 163.367
R645 B.n340 B.n101 163.367
R646 B.n340 B.n339 163.367
R647 B.n339 B.n338 163.367
R648 B.n338 B.n103 163.367
R649 B.n334 B.n103 163.367
R650 B.n334 B.n333 163.367
R651 B.n333 B.n332 163.367
R652 B.n332 B.n105 163.367
R653 B.n328 B.n105 163.367
R654 B.n328 B.n327 163.367
R655 B.n327 B.n326 163.367
R656 B.n326 B.n107 163.367
R657 B.n322 B.n107 163.367
R658 B.n322 B.n321 163.367
R659 B.n321 B.n320 163.367
R660 B.n320 B.n109 163.367
R661 B.n550 B.n549 163.367
R662 B.n549 B.n548 163.367
R663 B.n548 B.n29 163.367
R664 B.n544 B.n29 163.367
R665 B.n544 B.n543 163.367
R666 B.n543 B.n542 163.367
R667 B.n542 B.n31 163.367
R668 B.n538 B.n31 163.367
R669 B.n538 B.n537 163.367
R670 B.n537 B.n536 163.367
R671 B.n536 B.n33 163.367
R672 B.n532 B.n33 163.367
R673 B.n532 B.n531 163.367
R674 B.n531 B.n530 163.367
R675 B.n530 B.n35 163.367
R676 B.n526 B.n35 163.367
R677 B.n526 B.n525 163.367
R678 B.n525 B.n524 163.367
R679 B.n524 B.n37 163.367
R680 B.n520 B.n37 163.367
R681 B.n520 B.n519 163.367
R682 B.n519 B.n41 163.367
R683 B.n515 B.n41 163.367
R684 B.n515 B.n514 163.367
R685 B.n514 B.n513 163.367
R686 B.n513 B.n43 163.367
R687 B.n509 B.n43 163.367
R688 B.n509 B.n508 163.367
R689 B.n508 B.n507 163.367
R690 B.n507 B.n45 163.367
R691 B.n502 B.n45 163.367
R692 B.n502 B.n501 163.367
R693 B.n501 B.n500 163.367
R694 B.n500 B.n49 163.367
R695 B.n496 B.n49 163.367
R696 B.n496 B.n495 163.367
R697 B.n495 B.n494 163.367
R698 B.n494 B.n51 163.367
R699 B.n490 B.n51 163.367
R700 B.n490 B.n489 163.367
R701 B.n489 B.n488 163.367
R702 B.n488 B.n53 163.367
R703 B.n484 B.n53 163.367
R704 B.n484 B.n483 163.367
R705 B.n483 B.n482 163.367
R706 B.n482 B.n55 163.367
R707 B.n478 B.n55 163.367
R708 B.n478 B.n477 163.367
R709 B.n477 B.n476 163.367
R710 B.n476 B.n57 163.367
R711 B.n554 B.n27 163.367
R712 B.n555 B.n554 163.367
R713 B.n556 B.n555 163.367
R714 B.n556 B.n25 163.367
R715 B.n560 B.n25 163.367
R716 B.n561 B.n560 163.367
R717 B.n562 B.n561 163.367
R718 B.n562 B.n23 163.367
R719 B.n566 B.n23 163.367
R720 B.n567 B.n566 163.367
R721 B.n568 B.n567 163.367
R722 B.n568 B.n21 163.367
R723 B.n572 B.n21 163.367
R724 B.n573 B.n572 163.367
R725 B.n574 B.n573 163.367
R726 B.n574 B.n19 163.367
R727 B.n578 B.n19 163.367
R728 B.n579 B.n578 163.367
R729 B.n580 B.n579 163.367
R730 B.n580 B.n17 163.367
R731 B.n584 B.n17 163.367
R732 B.n585 B.n584 163.367
R733 B.n586 B.n585 163.367
R734 B.n586 B.n15 163.367
R735 B.n590 B.n15 163.367
R736 B.n591 B.n590 163.367
R737 B.n592 B.n591 163.367
R738 B.n592 B.n13 163.367
R739 B.n596 B.n13 163.367
R740 B.n597 B.n596 163.367
R741 B.n598 B.n597 163.367
R742 B.n598 B.n11 163.367
R743 B.n602 B.n11 163.367
R744 B.n603 B.n602 163.367
R745 B.n604 B.n603 163.367
R746 B.n604 B.n9 163.367
R747 B.n608 B.n9 163.367
R748 B.n609 B.n608 163.367
R749 B.n610 B.n609 163.367
R750 B.n610 B.n7 163.367
R751 B.n614 B.n7 163.367
R752 B.n615 B.n614 163.367
R753 B.n616 B.n615 163.367
R754 B.n616 B.n5 163.367
R755 B.n620 B.n5 163.367
R756 B.n621 B.n620 163.367
R757 B.n622 B.n621 163.367
R758 B.n622 B.n3 163.367
R759 B.n626 B.n3 163.367
R760 B.n627 B.n626 163.367
R761 B.n165 B.n2 163.367
R762 B.n166 B.n165 163.367
R763 B.n166 B.n163 163.367
R764 B.n170 B.n163 163.367
R765 B.n171 B.n170 163.367
R766 B.n172 B.n171 163.367
R767 B.n172 B.n161 163.367
R768 B.n176 B.n161 163.367
R769 B.n177 B.n176 163.367
R770 B.n178 B.n177 163.367
R771 B.n178 B.n159 163.367
R772 B.n182 B.n159 163.367
R773 B.n183 B.n182 163.367
R774 B.n184 B.n183 163.367
R775 B.n184 B.n157 163.367
R776 B.n188 B.n157 163.367
R777 B.n189 B.n188 163.367
R778 B.n190 B.n189 163.367
R779 B.n190 B.n155 163.367
R780 B.n194 B.n155 163.367
R781 B.n195 B.n194 163.367
R782 B.n196 B.n195 163.367
R783 B.n196 B.n153 163.367
R784 B.n200 B.n153 163.367
R785 B.n201 B.n200 163.367
R786 B.n202 B.n201 163.367
R787 B.n202 B.n151 163.367
R788 B.n206 B.n151 163.367
R789 B.n207 B.n206 163.367
R790 B.n208 B.n207 163.367
R791 B.n208 B.n149 163.367
R792 B.n212 B.n149 163.367
R793 B.n213 B.n212 163.367
R794 B.n214 B.n213 163.367
R795 B.n214 B.n147 163.367
R796 B.n218 B.n147 163.367
R797 B.n219 B.n218 163.367
R798 B.n220 B.n219 163.367
R799 B.n220 B.n145 163.367
R800 B.n224 B.n145 163.367
R801 B.n225 B.n224 163.367
R802 B.n226 B.n225 163.367
R803 B.n226 B.n143 163.367
R804 B.n230 B.n143 163.367
R805 B.n231 B.n230 163.367
R806 B.n232 B.n231 163.367
R807 B.n232 B.n141 163.367
R808 B.n236 B.n141 163.367
R809 B.n237 B.n236 163.367
R810 B.n238 B.n237 163.367
R811 B.n121 B.t8 117.186
R812 B.n47 B.t10 117.186
R813 B.n129 B.t2 117.183
R814 B.n39 B.t4 117.183
R815 B.n129 B.n128 71.952
R816 B.n121 B.n120 71.952
R817 B.n47 B.n46 71.952
R818 B.n39 B.n38 71.952
R819 B.n271 B.n129 59.5399
R820 B.n122 B.n121 59.5399
R821 B.n505 B.n47 59.5399
R822 B.n40 B.n39 59.5399
R823 B.n552 B.n551 35.1225
R824 B.n474 B.n473 35.1225
R825 B.n318 B.n317 35.1225
R826 B.n240 B.n239 35.1225
R827 B B.n629 18.0485
R828 B.n553 B.n552 10.6151
R829 B.n553 B.n26 10.6151
R830 B.n557 B.n26 10.6151
R831 B.n558 B.n557 10.6151
R832 B.n559 B.n558 10.6151
R833 B.n559 B.n24 10.6151
R834 B.n563 B.n24 10.6151
R835 B.n564 B.n563 10.6151
R836 B.n565 B.n564 10.6151
R837 B.n565 B.n22 10.6151
R838 B.n569 B.n22 10.6151
R839 B.n570 B.n569 10.6151
R840 B.n571 B.n570 10.6151
R841 B.n571 B.n20 10.6151
R842 B.n575 B.n20 10.6151
R843 B.n576 B.n575 10.6151
R844 B.n577 B.n576 10.6151
R845 B.n577 B.n18 10.6151
R846 B.n581 B.n18 10.6151
R847 B.n582 B.n581 10.6151
R848 B.n583 B.n582 10.6151
R849 B.n583 B.n16 10.6151
R850 B.n587 B.n16 10.6151
R851 B.n588 B.n587 10.6151
R852 B.n589 B.n588 10.6151
R853 B.n589 B.n14 10.6151
R854 B.n593 B.n14 10.6151
R855 B.n594 B.n593 10.6151
R856 B.n595 B.n594 10.6151
R857 B.n595 B.n12 10.6151
R858 B.n599 B.n12 10.6151
R859 B.n600 B.n599 10.6151
R860 B.n601 B.n600 10.6151
R861 B.n601 B.n10 10.6151
R862 B.n605 B.n10 10.6151
R863 B.n606 B.n605 10.6151
R864 B.n607 B.n606 10.6151
R865 B.n607 B.n8 10.6151
R866 B.n611 B.n8 10.6151
R867 B.n612 B.n611 10.6151
R868 B.n613 B.n612 10.6151
R869 B.n613 B.n6 10.6151
R870 B.n617 B.n6 10.6151
R871 B.n618 B.n617 10.6151
R872 B.n619 B.n618 10.6151
R873 B.n619 B.n4 10.6151
R874 B.n623 B.n4 10.6151
R875 B.n624 B.n623 10.6151
R876 B.n625 B.n624 10.6151
R877 B.n625 B.n0 10.6151
R878 B.n551 B.n28 10.6151
R879 B.n547 B.n28 10.6151
R880 B.n547 B.n546 10.6151
R881 B.n546 B.n545 10.6151
R882 B.n545 B.n30 10.6151
R883 B.n541 B.n30 10.6151
R884 B.n541 B.n540 10.6151
R885 B.n540 B.n539 10.6151
R886 B.n539 B.n32 10.6151
R887 B.n535 B.n32 10.6151
R888 B.n535 B.n534 10.6151
R889 B.n534 B.n533 10.6151
R890 B.n533 B.n34 10.6151
R891 B.n529 B.n34 10.6151
R892 B.n529 B.n528 10.6151
R893 B.n528 B.n527 10.6151
R894 B.n527 B.n36 10.6151
R895 B.n523 B.n36 10.6151
R896 B.n523 B.n522 10.6151
R897 B.n522 B.n521 10.6151
R898 B.n518 B.n517 10.6151
R899 B.n517 B.n516 10.6151
R900 B.n516 B.n42 10.6151
R901 B.n512 B.n42 10.6151
R902 B.n512 B.n511 10.6151
R903 B.n511 B.n510 10.6151
R904 B.n510 B.n44 10.6151
R905 B.n506 B.n44 10.6151
R906 B.n504 B.n503 10.6151
R907 B.n503 B.n48 10.6151
R908 B.n499 B.n48 10.6151
R909 B.n499 B.n498 10.6151
R910 B.n498 B.n497 10.6151
R911 B.n497 B.n50 10.6151
R912 B.n493 B.n50 10.6151
R913 B.n493 B.n492 10.6151
R914 B.n492 B.n491 10.6151
R915 B.n491 B.n52 10.6151
R916 B.n487 B.n52 10.6151
R917 B.n487 B.n486 10.6151
R918 B.n486 B.n485 10.6151
R919 B.n485 B.n54 10.6151
R920 B.n481 B.n54 10.6151
R921 B.n481 B.n480 10.6151
R922 B.n480 B.n479 10.6151
R923 B.n479 B.n56 10.6151
R924 B.n475 B.n56 10.6151
R925 B.n475 B.n474 10.6151
R926 B.n473 B.n58 10.6151
R927 B.n469 B.n58 10.6151
R928 B.n469 B.n468 10.6151
R929 B.n468 B.n467 10.6151
R930 B.n467 B.n60 10.6151
R931 B.n463 B.n60 10.6151
R932 B.n463 B.n462 10.6151
R933 B.n462 B.n461 10.6151
R934 B.n461 B.n62 10.6151
R935 B.n457 B.n62 10.6151
R936 B.n457 B.n456 10.6151
R937 B.n456 B.n455 10.6151
R938 B.n455 B.n64 10.6151
R939 B.n451 B.n64 10.6151
R940 B.n451 B.n450 10.6151
R941 B.n450 B.n449 10.6151
R942 B.n449 B.n66 10.6151
R943 B.n445 B.n66 10.6151
R944 B.n445 B.n444 10.6151
R945 B.n444 B.n443 10.6151
R946 B.n443 B.n68 10.6151
R947 B.n439 B.n68 10.6151
R948 B.n439 B.n438 10.6151
R949 B.n438 B.n437 10.6151
R950 B.n437 B.n70 10.6151
R951 B.n433 B.n70 10.6151
R952 B.n433 B.n432 10.6151
R953 B.n432 B.n431 10.6151
R954 B.n431 B.n72 10.6151
R955 B.n427 B.n72 10.6151
R956 B.n427 B.n426 10.6151
R957 B.n426 B.n425 10.6151
R958 B.n425 B.n74 10.6151
R959 B.n421 B.n74 10.6151
R960 B.n421 B.n420 10.6151
R961 B.n420 B.n419 10.6151
R962 B.n419 B.n76 10.6151
R963 B.n415 B.n76 10.6151
R964 B.n415 B.n414 10.6151
R965 B.n414 B.n413 10.6151
R966 B.n413 B.n78 10.6151
R967 B.n409 B.n78 10.6151
R968 B.n409 B.n408 10.6151
R969 B.n408 B.n407 10.6151
R970 B.n407 B.n80 10.6151
R971 B.n403 B.n80 10.6151
R972 B.n403 B.n402 10.6151
R973 B.n402 B.n401 10.6151
R974 B.n401 B.n82 10.6151
R975 B.n397 B.n82 10.6151
R976 B.n397 B.n396 10.6151
R977 B.n396 B.n395 10.6151
R978 B.n395 B.n84 10.6151
R979 B.n391 B.n84 10.6151
R980 B.n391 B.n390 10.6151
R981 B.n390 B.n389 10.6151
R982 B.n389 B.n86 10.6151
R983 B.n385 B.n86 10.6151
R984 B.n385 B.n384 10.6151
R985 B.n384 B.n383 10.6151
R986 B.n383 B.n88 10.6151
R987 B.n379 B.n88 10.6151
R988 B.n379 B.n378 10.6151
R989 B.n378 B.n377 10.6151
R990 B.n377 B.n90 10.6151
R991 B.n373 B.n90 10.6151
R992 B.n373 B.n372 10.6151
R993 B.n372 B.n371 10.6151
R994 B.n371 B.n92 10.6151
R995 B.n367 B.n92 10.6151
R996 B.n367 B.n366 10.6151
R997 B.n366 B.n365 10.6151
R998 B.n365 B.n94 10.6151
R999 B.n361 B.n94 10.6151
R1000 B.n361 B.n360 10.6151
R1001 B.n360 B.n359 10.6151
R1002 B.n359 B.n96 10.6151
R1003 B.n355 B.n96 10.6151
R1004 B.n355 B.n354 10.6151
R1005 B.n354 B.n353 10.6151
R1006 B.n353 B.n98 10.6151
R1007 B.n349 B.n98 10.6151
R1008 B.n349 B.n348 10.6151
R1009 B.n348 B.n347 10.6151
R1010 B.n347 B.n100 10.6151
R1011 B.n343 B.n100 10.6151
R1012 B.n343 B.n342 10.6151
R1013 B.n342 B.n341 10.6151
R1014 B.n341 B.n102 10.6151
R1015 B.n337 B.n102 10.6151
R1016 B.n337 B.n336 10.6151
R1017 B.n336 B.n335 10.6151
R1018 B.n335 B.n104 10.6151
R1019 B.n331 B.n104 10.6151
R1020 B.n331 B.n330 10.6151
R1021 B.n330 B.n329 10.6151
R1022 B.n329 B.n106 10.6151
R1023 B.n325 B.n106 10.6151
R1024 B.n325 B.n324 10.6151
R1025 B.n324 B.n323 10.6151
R1026 B.n323 B.n108 10.6151
R1027 B.n319 B.n108 10.6151
R1028 B.n319 B.n318 10.6151
R1029 B.n164 B.n1 10.6151
R1030 B.n167 B.n164 10.6151
R1031 B.n168 B.n167 10.6151
R1032 B.n169 B.n168 10.6151
R1033 B.n169 B.n162 10.6151
R1034 B.n173 B.n162 10.6151
R1035 B.n174 B.n173 10.6151
R1036 B.n175 B.n174 10.6151
R1037 B.n175 B.n160 10.6151
R1038 B.n179 B.n160 10.6151
R1039 B.n180 B.n179 10.6151
R1040 B.n181 B.n180 10.6151
R1041 B.n181 B.n158 10.6151
R1042 B.n185 B.n158 10.6151
R1043 B.n186 B.n185 10.6151
R1044 B.n187 B.n186 10.6151
R1045 B.n187 B.n156 10.6151
R1046 B.n191 B.n156 10.6151
R1047 B.n192 B.n191 10.6151
R1048 B.n193 B.n192 10.6151
R1049 B.n193 B.n154 10.6151
R1050 B.n197 B.n154 10.6151
R1051 B.n198 B.n197 10.6151
R1052 B.n199 B.n198 10.6151
R1053 B.n199 B.n152 10.6151
R1054 B.n203 B.n152 10.6151
R1055 B.n204 B.n203 10.6151
R1056 B.n205 B.n204 10.6151
R1057 B.n205 B.n150 10.6151
R1058 B.n209 B.n150 10.6151
R1059 B.n210 B.n209 10.6151
R1060 B.n211 B.n210 10.6151
R1061 B.n211 B.n148 10.6151
R1062 B.n215 B.n148 10.6151
R1063 B.n216 B.n215 10.6151
R1064 B.n217 B.n216 10.6151
R1065 B.n217 B.n146 10.6151
R1066 B.n221 B.n146 10.6151
R1067 B.n222 B.n221 10.6151
R1068 B.n223 B.n222 10.6151
R1069 B.n223 B.n144 10.6151
R1070 B.n227 B.n144 10.6151
R1071 B.n228 B.n227 10.6151
R1072 B.n229 B.n228 10.6151
R1073 B.n229 B.n142 10.6151
R1074 B.n233 B.n142 10.6151
R1075 B.n234 B.n233 10.6151
R1076 B.n235 B.n234 10.6151
R1077 B.n235 B.n140 10.6151
R1078 B.n239 B.n140 10.6151
R1079 B.n241 B.n240 10.6151
R1080 B.n241 B.n138 10.6151
R1081 B.n245 B.n138 10.6151
R1082 B.n246 B.n245 10.6151
R1083 B.n247 B.n246 10.6151
R1084 B.n247 B.n136 10.6151
R1085 B.n251 B.n136 10.6151
R1086 B.n252 B.n251 10.6151
R1087 B.n253 B.n252 10.6151
R1088 B.n253 B.n134 10.6151
R1089 B.n257 B.n134 10.6151
R1090 B.n258 B.n257 10.6151
R1091 B.n259 B.n258 10.6151
R1092 B.n259 B.n132 10.6151
R1093 B.n263 B.n132 10.6151
R1094 B.n264 B.n263 10.6151
R1095 B.n265 B.n264 10.6151
R1096 B.n265 B.n130 10.6151
R1097 B.n269 B.n130 10.6151
R1098 B.n270 B.n269 10.6151
R1099 B.n272 B.n126 10.6151
R1100 B.n276 B.n126 10.6151
R1101 B.n277 B.n276 10.6151
R1102 B.n278 B.n277 10.6151
R1103 B.n278 B.n124 10.6151
R1104 B.n282 B.n124 10.6151
R1105 B.n283 B.n282 10.6151
R1106 B.n284 B.n283 10.6151
R1107 B.n288 B.n287 10.6151
R1108 B.n289 B.n288 10.6151
R1109 B.n289 B.n118 10.6151
R1110 B.n293 B.n118 10.6151
R1111 B.n294 B.n293 10.6151
R1112 B.n295 B.n294 10.6151
R1113 B.n295 B.n116 10.6151
R1114 B.n299 B.n116 10.6151
R1115 B.n300 B.n299 10.6151
R1116 B.n301 B.n300 10.6151
R1117 B.n301 B.n114 10.6151
R1118 B.n305 B.n114 10.6151
R1119 B.n306 B.n305 10.6151
R1120 B.n307 B.n306 10.6151
R1121 B.n307 B.n112 10.6151
R1122 B.n311 B.n112 10.6151
R1123 B.n312 B.n311 10.6151
R1124 B.n313 B.n312 10.6151
R1125 B.n313 B.n110 10.6151
R1126 B.n317 B.n110 10.6151
R1127 B.n629 B.n0 8.11757
R1128 B.n629 B.n1 8.11757
R1129 B.n518 B.n40 6.5566
R1130 B.n506 B.n505 6.5566
R1131 B.n272 B.n271 6.5566
R1132 B.n284 B.n122 6.5566
R1133 B.n521 B.n40 4.05904
R1134 B.n505 B.n504 4.05904
R1135 B.n271 B.n270 4.05904
R1136 B.n287 B.n122 4.05904
C0 VDD2 VN 3.10161f
C1 VN B 1.27759f
C2 VDD2 VP 0.528355f
C3 w_n3938_n1946# VDD1 1.99287f
C4 B VP 2.13511f
C5 VN w_n3938_n1946# 7.53082f
C6 VDD2 VTAIL 5.67868f
C7 VN VDD1 0.155654f
C8 B VTAIL 2.29583f
C9 VP w_n3938_n1946# 8.042029f
C10 VP VDD1 3.47163f
C11 VDD2 B 1.81878f
C12 VN VP 6.37078f
C13 w_n3938_n1946# VTAIL 2.06523f
C14 VDD1 VTAIL 5.62067f
C15 VDD2 w_n3938_n1946# 2.10256f
C16 VDD2 VDD1 1.71097f
C17 B w_n3938_n1946# 8.77742f
C18 B VDD1 1.72585f
C19 VN VTAIL 3.9781f
C20 VP VTAIL 3.99226f
C21 VDD2 VSUBS 1.761227f
C22 VDD1 VSUBS 2.118421f
C23 VTAIL VSUBS 0.740588f
C24 VN VSUBS 6.37279f
C25 VP VSUBS 3.044908f
C26 B VSUBS 4.529469f
C27 w_n3938_n1946# VSUBS 96.071396f
C28 B.n0 VSUBS 0.008437f
C29 B.n1 VSUBS 0.008437f
C30 B.n2 VSUBS 0.012478f
C31 B.n3 VSUBS 0.009562f
C32 B.n4 VSUBS 0.009562f
C33 B.n5 VSUBS 0.009562f
C34 B.n6 VSUBS 0.009562f
C35 B.n7 VSUBS 0.009562f
C36 B.n8 VSUBS 0.009562f
C37 B.n9 VSUBS 0.009562f
C38 B.n10 VSUBS 0.009562f
C39 B.n11 VSUBS 0.009562f
C40 B.n12 VSUBS 0.009562f
C41 B.n13 VSUBS 0.009562f
C42 B.n14 VSUBS 0.009562f
C43 B.n15 VSUBS 0.009562f
C44 B.n16 VSUBS 0.009562f
C45 B.n17 VSUBS 0.009562f
C46 B.n18 VSUBS 0.009562f
C47 B.n19 VSUBS 0.009562f
C48 B.n20 VSUBS 0.009562f
C49 B.n21 VSUBS 0.009562f
C50 B.n22 VSUBS 0.009562f
C51 B.n23 VSUBS 0.009562f
C52 B.n24 VSUBS 0.009562f
C53 B.n25 VSUBS 0.009562f
C54 B.n26 VSUBS 0.009562f
C55 B.n27 VSUBS 0.022752f
C56 B.n28 VSUBS 0.009562f
C57 B.n29 VSUBS 0.009562f
C58 B.n30 VSUBS 0.009562f
C59 B.n31 VSUBS 0.009562f
C60 B.n32 VSUBS 0.009562f
C61 B.n33 VSUBS 0.009562f
C62 B.n34 VSUBS 0.009562f
C63 B.n35 VSUBS 0.009562f
C64 B.n36 VSUBS 0.009562f
C65 B.n37 VSUBS 0.009562f
C66 B.t4 VSUBS 0.185544f
C67 B.t5 VSUBS 0.218392f
C68 B.t3 VSUBS 1.08859f
C69 B.n38 VSUBS 0.148072f
C70 B.n39 VSUBS 0.099982f
C71 B.n40 VSUBS 0.022154f
C72 B.n41 VSUBS 0.009562f
C73 B.n42 VSUBS 0.009562f
C74 B.n43 VSUBS 0.009562f
C75 B.n44 VSUBS 0.009562f
C76 B.n45 VSUBS 0.009562f
C77 B.t10 VSUBS 0.185544f
C78 B.t11 VSUBS 0.218391f
C79 B.t9 VSUBS 1.08859f
C80 B.n46 VSUBS 0.148073f
C81 B.n47 VSUBS 0.099982f
C82 B.n48 VSUBS 0.009562f
C83 B.n49 VSUBS 0.009562f
C84 B.n50 VSUBS 0.009562f
C85 B.n51 VSUBS 0.009562f
C86 B.n52 VSUBS 0.009562f
C87 B.n53 VSUBS 0.009562f
C88 B.n54 VSUBS 0.009562f
C89 B.n55 VSUBS 0.009562f
C90 B.n56 VSUBS 0.009562f
C91 B.n57 VSUBS 0.024213f
C92 B.n58 VSUBS 0.009562f
C93 B.n59 VSUBS 0.009562f
C94 B.n60 VSUBS 0.009562f
C95 B.n61 VSUBS 0.009562f
C96 B.n62 VSUBS 0.009562f
C97 B.n63 VSUBS 0.009562f
C98 B.n64 VSUBS 0.009562f
C99 B.n65 VSUBS 0.009562f
C100 B.n66 VSUBS 0.009562f
C101 B.n67 VSUBS 0.009562f
C102 B.n68 VSUBS 0.009562f
C103 B.n69 VSUBS 0.009562f
C104 B.n70 VSUBS 0.009562f
C105 B.n71 VSUBS 0.009562f
C106 B.n72 VSUBS 0.009562f
C107 B.n73 VSUBS 0.009562f
C108 B.n74 VSUBS 0.009562f
C109 B.n75 VSUBS 0.009562f
C110 B.n76 VSUBS 0.009562f
C111 B.n77 VSUBS 0.009562f
C112 B.n78 VSUBS 0.009562f
C113 B.n79 VSUBS 0.009562f
C114 B.n80 VSUBS 0.009562f
C115 B.n81 VSUBS 0.009562f
C116 B.n82 VSUBS 0.009562f
C117 B.n83 VSUBS 0.009562f
C118 B.n84 VSUBS 0.009562f
C119 B.n85 VSUBS 0.009562f
C120 B.n86 VSUBS 0.009562f
C121 B.n87 VSUBS 0.009562f
C122 B.n88 VSUBS 0.009562f
C123 B.n89 VSUBS 0.009562f
C124 B.n90 VSUBS 0.009562f
C125 B.n91 VSUBS 0.009562f
C126 B.n92 VSUBS 0.009562f
C127 B.n93 VSUBS 0.009562f
C128 B.n94 VSUBS 0.009562f
C129 B.n95 VSUBS 0.009562f
C130 B.n96 VSUBS 0.009562f
C131 B.n97 VSUBS 0.009562f
C132 B.n98 VSUBS 0.009562f
C133 B.n99 VSUBS 0.009562f
C134 B.n100 VSUBS 0.009562f
C135 B.n101 VSUBS 0.009562f
C136 B.n102 VSUBS 0.009562f
C137 B.n103 VSUBS 0.009562f
C138 B.n104 VSUBS 0.009562f
C139 B.n105 VSUBS 0.009562f
C140 B.n106 VSUBS 0.009562f
C141 B.n107 VSUBS 0.009562f
C142 B.n108 VSUBS 0.009562f
C143 B.n109 VSUBS 0.022752f
C144 B.n110 VSUBS 0.009562f
C145 B.n111 VSUBS 0.009562f
C146 B.n112 VSUBS 0.009562f
C147 B.n113 VSUBS 0.009562f
C148 B.n114 VSUBS 0.009562f
C149 B.n115 VSUBS 0.009562f
C150 B.n116 VSUBS 0.009562f
C151 B.n117 VSUBS 0.009562f
C152 B.n118 VSUBS 0.009562f
C153 B.n119 VSUBS 0.009562f
C154 B.t8 VSUBS 0.185544f
C155 B.t7 VSUBS 0.218391f
C156 B.t6 VSUBS 1.08859f
C157 B.n120 VSUBS 0.148073f
C158 B.n121 VSUBS 0.099982f
C159 B.n122 VSUBS 0.022154f
C160 B.n123 VSUBS 0.009562f
C161 B.n124 VSUBS 0.009562f
C162 B.n125 VSUBS 0.009562f
C163 B.n126 VSUBS 0.009562f
C164 B.n127 VSUBS 0.009562f
C165 B.t2 VSUBS 0.185544f
C166 B.t1 VSUBS 0.218392f
C167 B.t0 VSUBS 1.08859f
C168 B.n128 VSUBS 0.148072f
C169 B.n129 VSUBS 0.099982f
C170 B.n130 VSUBS 0.009562f
C171 B.n131 VSUBS 0.009562f
C172 B.n132 VSUBS 0.009562f
C173 B.n133 VSUBS 0.009562f
C174 B.n134 VSUBS 0.009562f
C175 B.n135 VSUBS 0.009562f
C176 B.n136 VSUBS 0.009562f
C177 B.n137 VSUBS 0.009562f
C178 B.n138 VSUBS 0.009562f
C179 B.n139 VSUBS 0.024213f
C180 B.n140 VSUBS 0.009562f
C181 B.n141 VSUBS 0.009562f
C182 B.n142 VSUBS 0.009562f
C183 B.n143 VSUBS 0.009562f
C184 B.n144 VSUBS 0.009562f
C185 B.n145 VSUBS 0.009562f
C186 B.n146 VSUBS 0.009562f
C187 B.n147 VSUBS 0.009562f
C188 B.n148 VSUBS 0.009562f
C189 B.n149 VSUBS 0.009562f
C190 B.n150 VSUBS 0.009562f
C191 B.n151 VSUBS 0.009562f
C192 B.n152 VSUBS 0.009562f
C193 B.n153 VSUBS 0.009562f
C194 B.n154 VSUBS 0.009562f
C195 B.n155 VSUBS 0.009562f
C196 B.n156 VSUBS 0.009562f
C197 B.n157 VSUBS 0.009562f
C198 B.n158 VSUBS 0.009562f
C199 B.n159 VSUBS 0.009562f
C200 B.n160 VSUBS 0.009562f
C201 B.n161 VSUBS 0.009562f
C202 B.n162 VSUBS 0.009562f
C203 B.n163 VSUBS 0.009562f
C204 B.n164 VSUBS 0.009562f
C205 B.n165 VSUBS 0.009562f
C206 B.n166 VSUBS 0.009562f
C207 B.n167 VSUBS 0.009562f
C208 B.n168 VSUBS 0.009562f
C209 B.n169 VSUBS 0.009562f
C210 B.n170 VSUBS 0.009562f
C211 B.n171 VSUBS 0.009562f
C212 B.n172 VSUBS 0.009562f
C213 B.n173 VSUBS 0.009562f
C214 B.n174 VSUBS 0.009562f
C215 B.n175 VSUBS 0.009562f
C216 B.n176 VSUBS 0.009562f
C217 B.n177 VSUBS 0.009562f
C218 B.n178 VSUBS 0.009562f
C219 B.n179 VSUBS 0.009562f
C220 B.n180 VSUBS 0.009562f
C221 B.n181 VSUBS 0.009562f
C222 B.n182 VSUBS 0.009562f
C223 B.n183 VSUBS 0.009562f
C224 B.n184 VSUBS 0.009562f
C225 B.n185 VSUBS 0.009562f
C226 B.n186 VSUBS 0.009562f
C227 B.n187 VSUBS 0.009562f
C228 B.n188 VSUBS 0.009562f
C229 B.n189 VSUBS 0.009562f
C230 B.n190 VSUBS 0.009562f
C231 B.n191 VSUBS 0.009562f
C232 B.n192 VSUBS 0.009562f
C233 B.n193 VSUBS 0.009562f
C234 B.n194 VSUBS 0.009562f
C235 B.n195 VSUBS 0.009562f
C236 B.n196 VSUBS 0.009562f
C237 B.n197 VSUBS 0.009562f
C238 B.n198 VSUBS 0.009562f
C239 B.n199 VSUBS 0.009562f
C240 B.n200 VSUBS 0.009562f
C241 B.n201 VSUBS 0.009562f
C242 B.n202 VSUBS 0.009562f
C243 B.n203 VSUBS 0.009562f
C244 B.n204 VSUBS 0.009562f
C245 B.n205 VSUBS 0.009562f
C246 B.n206 VSUBS 0.009562f
C247 B.n207 VSUBS 0.009562f
C248 B.n208 VSUBS 0.009562f
C249 B.n209 VSUBS 0.009562f
C250 B.n210 VSUBS 0.009562f
C251 B.n211 VSUBS 0.009562f
C252 B.n212 VSUBS 0.009562f
C253 B.n213 VSUBS 0.009562f
C254 B.n214 VSUBS 0.009562f
C255 B.n215 VSUBS 0.009562f
C256 B.n216 VSUBS 0.009562f
C257 B.n217 VSUBS 0.009562f
C258 B.n218 VSUBS 0.009562f
C259 B.n219 VSUBS 0.009562f
C260 B.n220 VSUBS 0.009562f
C261 B.n221 VSUBS 0.009562f
C262 B.n222 VSUBS 0.009562f
C263 B.n223 VSUBS 0.009562f
C264 B.n224 VSUBS 0.009562f
C265 B.n225 VSUBS 0.009562f
C266 B.n226 VSUBS 0.009562f
C267 B.n227 VSUBS 0.009562f
C268 B.n228 VSUBS 0.009562f
C269 B.n229 VSUBS 0.009562f
C270 B.n230 VSUBS 0.009562f
C271 B.n231 VSUBS 0.009562f
C272 B.n232 VSUBS 0.009562f
C273 B.n233 VSUBS 0.009562f
C274 B.n234 VSUBS 0.009562f
C275 B.n235 VSUBS 0.009562f
C276 B.n236 VSUBS 0.009562f
C277 B.n237 VSUBS 0.009562f
C278 B.n238 VSUBS 0.022752f
C279 B.n239 VSUBS 0.022752f
C280 B.n240 VSUBS 0.024213f
C281 B.n241 VSUBS 0.009562f
C282 B.n242 VSUBS 0.009562f
C283 B.n243 VSUBS 0.009562f
C284 B.n244 VSUBS 0.009562f
C285 B.n245 VSUBS 0.009562f
C286 B.n246 VSUBS 0.009562f
C287 B.n247 VSUBS 0.009562f
C288 B.n248 VSUBS 0.009562f
C289 B.n249 VSUBS 0.009562f
C290 B.n250 VSUBS 0.009562f
C291 B.n251 VSUBS 0.009562f
C292 B.n252 VSUBS 0.009562f
C293 B.n253 VSUBS 0.009562f
C294 B.n254 VSUBS 0.009562f
C295 B.n255 VSUBS 0.009562f
C296 B.n256 VSUBS 0.009562f
C297 B.n257 VSUBS 0.009562f
C298 B.n258 VSUBS 0.009562f
C299 B.n259 VSUBS 0.009562f
C300 B.n260 VSUBS 0.009562f
C301 B.n261 VSUBS 0.009562f
C302 B.n262 VSUBS 0.009562f
C303 B.n263 VSUBS 0.009562f
C304 B.n264 VSUBS 0.009562f
C305 B.n265 VSUBS 0.009562f
C306 B.n266 VSUBS 0.009562f
C307 B.n267 VSUBS 0.009562f
C308 B.n268 VSUBS 0.009562f
C309 B.n269 VSUBS 0.009562f
C310 B.n270 VSUBS 0.006609f
C311 B.n271 VSUBS 0.022154f
C312 B.n272 VSUBS 0.007734f
C313 B.n273 VSUBS 0.009562f
C314 B.n274 VSUBS 0.009562f
C315 B.n275 VSUBS 0.009562f
C316 B.n276 VSUBS 0.009562f
C317 B.n277 VSUBS 0.009562f
C318 B.n278 VSUBS 0.009562f
C319 B.n279 VSUBS 0.009562f
C320 B.n280 VSUBS 0.009562f
C321 B.n281 VSUBS 0.009562f
C322 B.n282 VSUBS 0.009562f
C323 B.n283 VSUBS 0.009562f
C324 B.n284 VSUBS 0.007734f
C325 B.n285 VSUBS 0.009562f
C326 B.n286 VSUBS 0.009562f
C327 B.n287 VSUBS 0.006609f
C328 B.n288 VSUBS 0.009562f
C329 B.n289 VSUBS 0.009562f
C330 B.n290 VSUBS 0.009562f
C331 B.n291 VSUBS 0.009562f
C332 B.n292 VSUBS 0.009562f
C333 B.n293 VSUBS 0.009562f
C334 B.n294 VSUBS 0.009562f
C335 B.n295 VSUBS 0.009562f
C336 B.n296 VSUBS 0.009562f
C337 B.n297 VSUBS 0.009562f
C338 B.n298 VSUBS 0.009562f
C339 B.n299 VSUBS 0.009562f
C340 B.n300 VSUBS 0.009562f
C341 B.n301 VSUBS 0.009562f
C342 B.n302 VSUBS 0.009562f
C343 B.n303 VSUBS 0.009562f
C344 B.n304 VSUBS 0.009562f
C345 B.n305 VSUBS 0.009562f
C346 B.n306 VSUBS 0.009562f
C347 B.n307 VSUBS 0.009562f
C348 B.n308 VSUBS 0.009562f
C349 B.n309 VSUBS 0.009562f
C350 B.n310 VSUBS 0.009562f
C351 B.n311 VSUBS 0.009562f
C352 B.n312 VSUBS 0.009562f
C353 B.n313 VSUBS 0.009562f
C354 B.n314 VSUBS 0.009562f
C355 B.n315 VSUBS 0.009562f
C356 B.n316 VSUBS 0.024213f
C357 B.n317 VSUBS 0.023162f
C358 B.n318 VSUBS 0.023803f
C359 B.n319 VSUBS 0.009562f
C360 B.n320 VSUBS 0.009562f
C361 B.n321 VSUBS 0.009562f
C362 B.n322 VSUBS 0.009562f
C363 B.n323 VSUBS 0.009562f
C364 B.n324 VSUBS 0.009562f
C365 B.n325 VSUBS 0.009562f
C366 B.n326 VSUBS 0.009562f
C367 B.n327 VSUBS 0.009562f
C368 B.n328 VSUBS 0.009562f
C369 B.n329 VSUBS 0.009562f
C370 B.n330 VSUBS 0.009562f
C371 B.n331 VSUBS 0.009562f
C372 B.n332 VSUBS 0.009562f
C373 B.n333 VSUBS 0.009562f
C374 B.n334 VSUBS 0.009562f
C375 B.n335 VSUBS 0.009562f
C376 B.n336 VSUBS 0.009562f
C377 B.n337 VSUBS 0.009562f
C378 B.n338 VSUBS 0.009562f
C379 B.n339 VSUBS 0.009562f
C380 B.n340 VSUBS 0.009562f
C381 B.n341 VSUBS 0.009562f
C382 B.n342 VSUBS 0.009562f
C383 B.n343 VSUBS 0.009562f
C384 B.n344 VSUBS 0.009562f
C385 B.n345 VSUBS 0.009562f
C386 B.n346 VSUBS 0.009562f
C387 B.n347 VSUBS 0.009562f
C388 B.n348 VSUBS 0.009562f
C389 B.n349 VSUBS 0.009562f
C390 B.n350 VSUBS 0.009562f
C391 B.n351 VSUBS 0.009562f
C392 B.n352 VSUBS 0.009562f
C393 B.n353 VSUBS 0.009562f
C394 B.n354 VSUBS 0.009562f
C395 B.n355 VSUBS 0.009562f
C396 B.n356 VSUBS 0.009562f
C397 B.n357 VSUBS 0.009562f
C398 B.n358 VSUBS 0.009562f
C399 B.n359 VSUBS 0.009562f
C400 B.n360 VSUBS 0.009562f
C401 B.n361 VSUBS 0.009562f
C402 B.n362 VSUBS 0.009562f
C403 B.n363 VSUBS 0.009562f
C404 B.n364 VSUBS 0.009562f
C405 B.n365 VSUBS 0.009562f
C406 B.n366 VSUBS 0.009562f
C407 B.n367 VSUBS 0.009562f
C408 B.n368 VSUBS 0.009562f
C409 B.n369 VSUBS 0.009562f
C410 B.n370 VSUBS 0.009562f
C411 B.n371 VSUBS 0.009562f
C412 B.n372 VSUBS 0.009562f
C413 B.n373 VSUBS 0.009562f
C414 B.n374 VSUBS 0.009562f
C415 B.n375 VSUBS 0.009562f
C416 B.n376 VSUBS 0.009562f
C417 B.n377 VSUBS 0.009562f
C418 B.n378 VSUBS 0.009562f
C419 B.n379 VSUBS 0.009562f
C420 B.n380 VSUBS 0.009562f
C421 B.n381 VSUBS 0.009562f
C422 B.n382 VSUBS 0.009562f
C423 B.n383 VSUBS 0.009562f
C424 B.n384 VSUBS 0.009562f
C425 B.n385 VSUBS 0.009562f
C426 B.n386 VSUBS 0.009562f
C427 B.n387 VSUBS 0.009562f
C428 B.n388 VSUBS 0.009562f
C429 B.n389 VSUBS 0.009562f
C430 B.n390 VSUBS 0.009562f
C431 B.n391 VSUBS 0.009562f
C432 B.n392 VSUBS 0.009562f
C433 B.n393 VSUBS 0.009562f
C434 B.n394 VSUBS 0.009562f
C435 B.n395 VSUBS 0.009562f
C436 B.n396 VSUBS 0.009562f
C437 B.n397 VSUBS 0.009562f
C438 B.n398 VSUBS 0.009562f
C439 B.n399 VSUBS 0.009562f
C440 B.n400 VSUBS 0.009562f
C441 B.n401 VSUBS 0.009562f
C442 B.n402 VSUBS 0.009562f
C443 B.n403 VSUBS 0.009562f
C444 B.n404 VSUBS 0.009562f
C445 B.n405 VSUBS 0.009562f
C446 B.n406 VSUBS 0.009562f
C447 B.n407 VSUBS 0.009562f
C448 B.n408 VSUBS 0.009562f
C449 B.n409 VSUBS 0.009562f
C450 B.n410 VSUBS 0.009562f
C451 B.n411 VSUBS 0.009562f
C452 B.n412 VSUBS 0.009562f
C453 B.n413 VSUBS 0.009562f
C454 B.n414 VSUBS 0.009562f
C455 B.n415 VSUBS 0.009562f
C456 B.n416 VSUBS 0.009562f
C457 B.n417 VSUBS 0.009562f
C458 B.n418 VSUBS 0.009562f
C459 B.n419 VSUBS 0.009562f
C460 B.n420 VSUBS 0.009562f
C461 B.n421 VSUBS 0.009562f
C462 B.n422 VSUBS 0.009562f
C463 B.n423 VSUBS 0.009562f
C464 B.n424 VSUBS 0.009562f
C465 B.n425 VSUBS 0.009562f
C466 B.n426 VSUBS 0.009562f
C467 B.n427 VSUBS 0.009562f
C468 B.n428 VSUBS 0.009562f
C469 B.n429 VSUBS 0.009562f
C470 B.n430 VSUBS 0.009562f
C471 B.n431 VSUBS 0.009562f
C472 B.n432 VSUBS 0.009562f
C473 B.n433 VSUBS 0.009562f
C474 B.n434 VSUBS 0.009562f
C475 B.n435 VSUBS 0.009562f
C476 B.n436 VSUBS 0.009562f
C477 B.n437 VSUBS 0.009562f
C478 B.n438 VSUBS 0.009562f
C479 B.n439 VSUBS 0.009562f
C480 B.n440 VSUBS 0.009562f
C481 B.n441 VSUBS 0.009562f
C482 B.n442 VSUBS 0.009562f
C483 B.n443 VSUBS 0.009562f
C484 B.n444 VSUBS 0.009562f
C485 B.n445 VSUBS 0.009562f
C486 B.n446 VSUBS 0.009562f
C487 B.n447 VSUBS 0.009562f
C488 B.n448 VSUBS 0.009562f
C489 B.n449 VSUBS 0.009562f
C490 B.n450 VSUBS 0.009562f
C491 B.n451 VSUBS 0.009562f
C492 B.n452 VSUBS 0.009562f
C493 B.n453 VSUBS 0.009562f
C494 B.n454 VSUBS 0.009562f
C495 B.n455 VSUBS 0.009562f
C496 B.n456 VSUBS 0.009562f
C497 B.n457 VSUBS 0.009562f
C498 B.n458 VSUBS 0.009562f
C499 B.n459 VSUBS 0.009562f
C500 B.n460 VSUBS 0.009562f
C501 B.n461 VSUBS 0.009562f
C502 B.n462 VSUBS 0.009562f
C503 B.n463 VSUBS 0.009562f
C504 B.n464 VSUBS 0.009562f
C505 B.n465 VSUBS 0.009562f
C506 B.n466 VSUBS 0.009562f
C507 B.n467 VSUBS 0.009562f
C508 B.n468 VSUBS 0.009562f
C509 B.n469 VSUBS 0.009562f
C510 B.n470 VSUBS 0.009562f
C511 B.n471 VSUBS 0.009562f
C512 B.n472 VSUBS 0.022752f
C513 B.n473 VSUBS 0.022752f
C514 B.n474 VSUBS 0.024213f
C515 B.n475 VSUBS 0.009562f
C516 B.n476 VSUBS 0.009562f
C517 B.n477 VSUBS 0.009562f
C518 B.n478 VSUBS 0.009562f
C519 B.n479 VSUBS 0.009562f
C520 B.n480 VSUBS 0.009562f
C521 B.n481 VSUBS 0.009562f
C522 B.n482 VSUBS 0.009562f
C523 B.n483 VSUBS 0.009562f
C524 B.n484 VSUBS 0.009562f
C525 B.n485 VSUBS 0.009562f
C526 B.n486 VSUBS 0.009562f
C527 B.n487 VSUBS 0.009562f
C528 B.n488 VSUBS 0.009562f
C529 B.n489 VSUBS 0.009562f
C530 B.n490 VSUBS 0.009562f
C531 B.n491 VSUBS 0.009562f
C532 B.n492 VSUBS 0.009562f
C533 B.n493 VSUBS 0.009562f
C534 B.n494 VSUBS 0.009562f
C535 B.n495 VSUBS 0.009562f
C536 B.n496 VSUBS 0.009562f
C537 B.n497 VSUBS 0.009562f
C538 B.n498 VSUBS 0.009562f
C539 B.n499 VSUBS 0.009562f
C540 B.n500 VSUBS 0.009562f
C541 B.n501 VSUBS 0.009562f
C542 B.n502 VSUBS 0.009562f
C543 B.n503 VSUBS 0.009562f
C544 B.n504 VSUBS 0.006609f
C545 B.n505 VSUBS 0.022154f
C546 B.n506 VSUBS 0.007734f
C547 B.n507 VSUBS 0.009562f
C548 B.n508 VSUBS 0.009562f
C549 B.n509 VSUBS 0.009562f
C550 B.n510 VSUBS 0.009562f
C551 B.n511 VSUBS 0.009562f
C552 B.n512 VSUBS 0.009562f
C553 B.n513 VSUBS 0.009562f
C554 B.n514 VSUBS 0.009562f
C555 B.n515 VSUBS 0.009562f
C556 B.n516 VSUBS 0.009562f
C557 B.n517 VSUBS 0.009562f
C558 B.n518 VSUBS 0.007734f
C559 B.n519 VSUBS 0.009562f
C560 B.n520 VSUBS 0.009562f
C561 B.n521 VSUBS 0.006609f
C562 B.n522 VSUBS 0.009562f
C563 B.n523 VSUBS 0.009562f
C564 B.n524 VSUBS 0.009562f
C565 B.n525 VSUBS 0.009562f
C566 B.n526 VSUBS 0.009562f
C567 B.n527 VSUBS 0.009562f
C568 B.n528 VSUBS 0.009562f
C569 B.n529 VSUBS 0.009562f
C570 B.n530 VSUBS 0.009562f
C571 B.n531 VSUBS 0.009562f
C572 B.n532 VSUBS 0.009562f
C573 B.n533 VSUBS 0.009562f
C574 B.n534 VSUBS 0.009562f
C575 B.n535 VSUBS 0.009562f
C576 B.n536 VSUBS 0.009562f
C577 B.n537 VSUBS 0.009562f
C578 B.n538 VSUBS 0.009562f
C579 B.n539 VSUBS 0.009562f
C580 B.n540 VSUBS 0.009562f
C581 B.n541 VSUBS 0.009562f
C582 B.n542 VSUBS 0.009562f
C583 B.n543 VSUBS 0.009562f
C584 B.n544 VSUBS 0.009562f
C585 B.n545 VSUBS 0.009562f
C586 B.n546 VSUBS 0.009562f
C587 B.n547 VSUBS 0.009562f
C588 B.n548 VSUBS 0.009562f
C589 B.n549 VSUBS 0.009562f
C590 B.n550 VSUBS 0.024213f
C591 B.n551 VSUBS 0.024213f
C592 B.n552 VSUBS 0.022752f
C593 B.n553 VSUBS 0.009562f
C594 B.n554 VSUBS 0.009562f
C595 B.n555 VSUBS 0.009562f
C596 B.n556 VSUBS 0.009562f
C597 B.n557 VSUBS 0.009562f
C598 B.n558 VSUBS 0.009562f
C599 B.n559 VSUBS 0.009562f
C600 B.n560 VSUBS 0.009562f
C601 B.n561 VSUBS 0.009562f
C602 B.n562 VSUBS 0.009562f
C603 B.n563 VSUBS 0.009562f
C604 B.n564 VSUBS 0.009562f
C605 B.n565 VSUBS 0.009562f
C606 B.n566 VSUBS 0.009562f
C607 B.n567 VSUBS 0.009562f
C608 B.n568 VSUBS 0.009562f
C609 B.n569 VSUBS 0.009562f
C610 B.n570 VSUBS 0.009562f
C611 B.n571 VSUBS 0.009562f
C612 B.n572 VSUBS 0.009562f
C613 B.n573 VSUBS 0.009562f
C614 B.n574 VSUBS 0.009562f
C615 B.n575 VSUBS 0.009562f
C616 B.n576 VSUBS 0.009562f
C617 B.n577 VSUBS 0.009562f
C618 B.n578 VSUBS 0.009562f
C619 B.n579 VSUBS 0.009562f
C620 B.n580 VSUBS 0.009562f
C621 B.n581 VSUBS 0.009562f
C622 B.n582 VSUBS 0.009562f
C623 B.n583 VSUBS 0.009562f
C624 B.n584 VSUBS 0.009562f
C625 B.n585 VSUBS 0.009562f
C626 B.n586 VSUBS 0.009562f
C627 B.n587 VSUBS 0.009562f
C628 B.n588 VSUBS 0.009562f
C629 B.n589 VSUBS 0.009562f
C630 B.n590 VSUBS 0.009562f
C631 B.n591 VSUBS 0.009562f
C632 B.n592 VSUBS 0.009562f
C633 B.n593 VSUBS 0.009562f
C634 B.n594 VSUBS 0.009562f
C635 B.n595 VSUBS 0.009562f
C636 B.n596 VSUBS 0.009562f
C637 B.n597 VSUBS 0.009562f
C638 B.n598 VSUBS 0.009562f
C639 B.n599 VSUBS 0.009562f
C640 B.n600 VSUBS 0.009562f
C641 B.n601 VSUBS 0.009562f
C642 B.n602 VSUBS 0.009562f
C643 B.n603 VSUBS 0.009562f
C644 B.n604 VSUBS 0.009562f
C645 B.n605 VSUBS 0.009562f
C646 B.n606 VSUBS 0.009562f
C647 B.n607 VSUBS 0.009562f
C648 B.n608 VSUBS 0.009562f
C649 B.n609 VSUBS 0.009562f
C650 B.n610 VSUBS 0.009562f
C651 B.n611 VSUBS 0.009562f
C652 B.n612 VSUBS 0.009562f
C653 B.n613 VSUBS 0.009562f
C654 B.n614 VSUBS 0.009562f
C655 B.n615 VSUBS 0.009562f
C656 B.n616 VSUBS 0.009562f
C657 B.n617 VSUBS 0.009562f
C658 B.n618 VSUBS 0.009562f
C659 B.n619 VSUBS 0.009562f
C660 B.n620 VSUBS 0.009562f
C661 B.n621 VSUBS 0.009562f
C662 B.n622 VSUBS 0.009562f
C663 B.n623 VSUBS 0.009562f
C664 B.n624 VSUBS 0.009562f
C665 B.n625 VSUBS 0.009562f
C666 B.n626 VSUBS 0.009562f
C667 B.n627 VSUBS 0.012478f
C668 B.n628 VSUBS 0.013292f
C669 B.n629 VSUBS 0.026432f
C670 VDD1.t5 VSUBS 0.752706f
C671 VDD1.t2 VSUBS 0.751943f
C672 VDD1.t1 VSUBS 0.087398f
C673 VDD1.t0 VSUBS 0.087398f
C674 VDD1.n0 VSUBS 0.549526f
C675 VDD1.n1 VSUBS 2.97026f
C676 VDD1.t4 VSUBS 0.087398f
C677 VDD1.t3 VSUBS 0.087398f
C678 VDD1.n2 VSUBS 0.54478f
C679 VDD1.n3 VSUBS 2.38513f
C680 VP.t5 VSUBS 1.83147f
C681 VP.n0 VSUBS 0.853395f
C682 VP.n1 VSUBS 0.042432f
C683 VP.n2 VSUBS 0.047339f
C684 VP.n3 VSUBS 0.042432f
C685 VP.t4 VSUBS 1.83147f
C686 VP.n4 VSUBS 0.734231f
C687 VP.n5 VSUBS 0.042432f
C688 VP.n6 VSUBS 0.047339f
C689 VP.n7 VSUBS 0.042432f
C690 VP.t3 VSUBS 1.83147f
C691 VP.n8 VSUBS 0.853395f
C692 VP.t2 VSUBS 1.83147f
C693 VP.n9 VSUBS 0.853395f
C694 VP.n10 VSUBS 0.042432f
C695 VP.n11 VSUBS 0.047339f
C696 VP.n12 VSUBS 0.042432f
C697 VP.t1 VSUBS 1.83147f
C698 VP.n13 VSUBS 0.861397f
C699 VP.t0 VSUBS 2.32432f
C700 VP.n14 VSUBS 0.814204f
C701 VP.n15 VSUBS 0.517946f
C702 VP.n16 VSUBS 0.079083f
C703 VP.n17 VSUBS 0.079083f
C704 VP.n18 VSUBS 0.073913f
C705 VP.n19 VSUBS 0.042432f
C706 VP.n20 VSUBS 0.042432f
C707 VP.n21 VSUBS 0.042432f
C708 VP.n22 VSUBS 0.081725f
C709 VP.n23 VSUBS 0.079083f
C710 VP.n24 VSUBS 0.056437f
C711 VP.n25 VSUBS 0.068485f
C712 VP.n26 VSUBS 2.17207f
C713 VP.n27 VSUBS 2.20493f
C714 VP.n28 VSUBS 0.068485f
C715 VP.n29 VSUBS 0.056437f
C716 VP.n30 VSUBS 0.079083f
C717 VP.n31 VSUBS 0.081725f
C718 VP.n32 VSUBS 0.042432f
C719 VP.n33 VSUBS 0.042432f
C720 VP.n34 VSUBS 0.042432f
C721 VP.n35 VSUBS 0.073913f
C722 VP.n36 VSUBS 0.079083f
C723 VP.n37 VSUBS 0.079083f
C724 VP.n38 VSUBS 0.042432f
C725 VP.n39 VSUBS 0.042432f
C726 VP.n40 VSUBS 0.042432f
C727 VP.n41 VSUBS 0.079083f
C728 VP.n42 VSUBS 0.079083f
C729 VP.n43 VSUBS 0.073913f
C730 VP.n44 VSUBS 0.042432f
C731 VP.n45 VSUBS 0.042432f
C732 VP.n46 VSUBS 0.042432f
C733 VP.n47 VSUBS 0.081725f
C734 VP.n48 VSUBS 0.079083f
C735 VP.n49 VSUBS 0.056437f
C736 VP.n50 VSUBS 0.068485f
C737 VP.n51 VSUBS 0.111148f
C738 VDD2.t1 VSUBS 0.909024f
C739 VDD2.t4 VSUBS 0.105656f
C740 VDD2.t5 VSUBS 0.105656f
C741 VDD2.n0 VSUBS 0.664322f
C742 VDD2.n1 VSUBS 3.44089f
C743 VDD2.t3 VSUBS 0.894247f
C744 VDD2.n2 VSUBS 2.85411f
C745 VDD2.t0 VSUBS 0.105656f
C746 VDD2.t2 VSUBS 0.105656f
C747 VDD2.n3 VSUBS 0.664291f
C748 VTAIL.t8 VSUBS 0.13954f
C749 VTAIL.t11 VSUBS 0.13954f
C750 VTAIL.n0 VSUBS 0.760922f
C751 VTAIL.n1 VSUBS 0.950171f
C752 VTAIL.t3 VSUBS 1.06734f
C753 VTAIL.n2 VSUBS 1.29665f
C754 VTAIL.t0 VSUBS 0.13954f
C755 VTAIL.t1 VSUBS 0.13954f
C756 VTAIL.n3 VSUBS 0.760922f
C757 VTAIL.n4 VSUBS 2.70708f
C758 VTAIL.t10 VSUBS 0.13954f
C759 VTAIL.t9 VSUBS 0.13954f
C760 VTAIL.n5 VSUBS 0.760927f
C761 VTAIL.n6 VSUBS 2.70707f
C762 VTAIL.t7 VSUBS 1.06735f
C763 VTAIL.n7 VSUBS 1.29665f
C764 VTAIL.t5 VSUBS 0.13954f
C765 VTAIL.t2 VSUBS 0.13954f
C766 VTAIL.n8 VSUBS 0.760927f
C767 VTAIL.n9 VSUBS 1.2225f
C768 VTAIL.t4 VSUBS 1.06734f
C769 VTAIL.n10 VSUBS 2.40908f
C770 VTAIL.t6 VSUBS 1.06734f
C771 VTAIL.n11 VSUBS 2.30927f
C772 VN.t0 VSUBS 1.59856f
C773 VN.n0 VSUBS 0.744869f
C774 VN.n1 VSUBS 0.037036f
C775 VN.n2 VSUBS 0.041319f
C776 VN.n3 VSUBS 0.037036f
C777 VN.t1 VSUBS 1.59856f
C778 VN.n4 VSUBS 0.751853f
C779 VN.t4 VSUBS 2.02874f
C780 VN.n5 VSUBS 0.710661f
C781 VN.n6 VSUBS 0.452078f
C782 VN.n7 VSUBS 0.069026f
C783 VN.n8 VSUBS 0.069026f
C784 VN.n9 VSUBS 0.064514f
C785 VN.n10 VSUBS 0.037036f
C786 VN.n11 VSUBS 0.037036f
C787 VN.n12 VSUBS 0.037036f
C788 VN.n13 VSUBS 0.071332f
C789 VN.n14 VSUBS 0.069026f
C790 VN.n15 VSUBS 0.04926f
C791 VN.n16 VSUBS 0.059775f
C792 VN.n17 VSUBS 0.097013f
C793 VN.t2 VSUBS 1.59856f
C794 VN.n18 VSUBS 0.744869f
C795 VN.n19 VSUBS 0.037036f
C796 VN.n20 VSUBS 0.041319f
C797 VN.n21 VSUBS 0.037036f
C798 VN.t5 VSUBS 1.59856f
C799 VN.n22 VSUBS 0.751853f
C800 VN.t3 VSUBS 2.02874f
C801 VN.n23 VSUBS 0.710661f
C802 VN.n24 VSUBS 0.452078f
C803 VN.n25 VSUBS 0.069026f
C804 VN.n26 VSUBS 0.069026f
C805 VN.n27 VSUBS 0.064514f
C806 VN.n28 VSUBS 0.037036f
C807 VN.n29 VSUBS 0.037036f
C808 VN.n30 VSUBS 0.037036f
C809 VN.n31 VSUBS 0.071332f
C810 VN.n32 VSUBS 0.069026f
C811 VN.n33 VSUBS 0.04926f
C812 VN.n34 VSUBS 0.059775f
C813 VN.n35 VSUBS 1.91141f
.ends

