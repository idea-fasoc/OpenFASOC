* NGSPICE file created from diff_pair_sample_1214.ext - technology: sky130A

.subckt diff_pair_sample_1214 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t9 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X1 B.t11 B.t9 B.t10 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=0.97
X2 B.t8 B.t6 B.t7 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=0.97
X3 B.t5 B.t3 B.t4 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=0.97
X4 VTAIL.t6 VP.t0 VDD1.t9 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X5 VTAIL.t7 VP.t1 VDD1.t8 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X6 VDD2.t1 VN.t1 VTAIL.t16 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=2.3088 ps=12.62 w=5.92 l=0.97
X7 VDD2.t3 VN.t2 VTAIL.t15 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X8 B.t2 B.t0 B.t1 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0 ps=0 w=5.92 l=0.97
X9 VTAIL.t14 VN.t3 VDD2.t6 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X10 VDD2.t7 VN.t4 VTAIL.t13 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0.9768 ps=6.25 w=5.92 l=0.97
X11 VDD1.t7 VP.t2 VTAIL.t18 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0.9768 ps=6.25 w=5.92 l=0.97
X12 VTAIL.t19 VP.t3 VDD1.t6 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X13 VTAIL.t12 VN.t5 VDD2.t5 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X14 VTAIL.t11 VN.t6 VDD2.t4 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X15 VDD1.t5 VP.t4 VTAIL.t2 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=2.3088 ps=12.62 w=5.92 l=0.97
X16 VDD1.t4 VP.t5 VTAIL.t4 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=2.3088 ps=12.62 w=5.92 l=0.97
X17 VDD1.t3 VP.t6 VTAIL.t5 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X18 VDD1.t2 VP.t7 VTAIL.t1 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X19 VDD1.t1 VP.t8 VTAIL.t3 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0.9768 ps=6.25 w=5.92 l=0.97
X20 VTAIL.t0 VP.t9 VDD1.t0 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X21 VDD2.t8 VN.t7 VTAIL.t10 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=2.3088 pd=12.62 as=0.9768 ps=6.25 w=5.92 l=0.97
X22 VDD2.t0 VN.t8 VTAIL.t9 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=0.9768 ps=6.25 w=5.92 l=0.97
X23 VDD2.t2 VN.t9 VTAIL.t8 w_n2530_n2152# sky130_fd_pr__pfet_01v8 ad=0.9768 pd=6.25 as=2.3088 ps=12.62 w=5.92 l=0.97
R0 VN.n5 VN.t7 201.407
R1 VN.n25 VN.t1 201.407
R2 VN.n18 VN.t9 187.583
R3 VN.n38 VN.t4 187.583
R4 VN.n37 VN.n20 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n21 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n29 VN.n22 161.3
R9 VN.n28 VN.n27 161.3
R10 VN.n26 VN.n23 161.3
R11 VN.n17 VN.n0 161.3
R12 VN.n15 VN.n14 161.3
R13 VN.n13 VN.n1 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n9 VN.n2 161.3
R16 VN.n8 VN.n7 161.3
R17 VN.n6 VN.n3 161.3
R18 VN.n4 VN.t0 147.085
R19 VN.n10 VN.t8 147.085
R20 VN.n16 VN.t3 147.085
R21 VN.n24 VN.t5 147.085
R22 VN.n30 VN.t2 147.085
R23 VN.n36 VN.t6 147.085
R24 VN.n39 VN.n38 80.6037
R25 VN.n19 VN.n18 80.6037
R26 VN.n9 VN.n8 50.2647
R27 VN.n11 VN.n1 50.2647
R28 VN.n29 VN.n28 50.2647
R29 VN.n31 VN.n21 50.2647
R30 VN.n18 VN.n17 49.9219
R31 VN.n38 VN.n37 49.9219
R32 VN.n5 VN.n4 49.6998
R33 VN.n25 VN.n24 49.6998
R34 VN.n26 VN.n25 44.8559
R35 VN.n6 VN.n5 44.8559
R36 VN VN.n39 40.0294
R37 VN.n8 VN.n3 30.8893
R38 VN.n15 VN.n1 30.8893
R39 VN.n28 VN.n23 30.8893
R40 VN.n35 VN.n21 30.8893
R41 VN.n17 VN.n16 22.1332
R42 VN.n37 VN.n36 22.1332
R43 VN.n10 VN.n9 12.2964
R44 VN.n11 VN.n10 12.2964
R45 VN.n31 VN.n30 12.2964
R46 VN.n30 VN.n29 12.2964
R47 VN.n4 VN.n3 2.45968
R48 VN.n16 VN.n15 2.45968
R49 VN.n24 VN.n23 2.45968
R50 VN.n36 VN.n35 2.45968
R51 VN.n39 VN.n20 0.285035
R52 VN.n19 VN.n0 0.285035
R53 VN.n34 VN.n20 0.189894
R54 VN.n34 VN.n33 0.189894
R55 VN.n33 VN.n32 0.189894
R56 VN.n32 VN.n22 0.189894
R57 VN.n27 VN.n22 0.189894
R58 VN.n27 VN.n26 0.189894
R59 VN.n7 VN.n6 0.189894
R60 VN.n7 VN.n2 0.189894
R61 VN.n12 VN.n2 0.189894
R62 VN.n13 VN.n12 0.189894
R63 VN.n14 VN.n13 0.189894
R64 VN.n14 VN.n0 0.189894
R65 VN VN.n19 0.146778
R66 VDD2.n61 VDD2.n35 756.745
R67 VDD2.n26 VDD2.n0 756.745
R68 VDD2.n62 VDD2.n61 585
R69 VDD2.n60 VDD2.n59 585
R70 VDD2.n39 VDD2.n38 585
R71 VDD2.n54 VDD2.n53 585
R72 VDD2.n52 VDD2.n51 585
R73 VDD2.n43 VDD2.n42 585
R74 VDD2.n46 VDD2.n45 585
R75 VDD2.n11 VDD2.n10 585
R76 VDD2.n8 VDD2.n7 585
R77 VDD2.n17 VDD2.n16 585
R78 VDD2.n19 VDD2.n18 585
R79 VDD2.n4 VDD2.n3 585
R80 VDD2.n25 VDD2.n24 585
R81 VDD2.n27 VDD2.n26 585
R82 VDD2.t7 VDD2.n44 327.601
R83 VDD2.t8 VDD2.n9 327.601
R84 VDD2.n61 VDD2.n60 171.744
R85 VDD2.n60 VDD2.n38 171.744
R86 VDD2.n53 VDD2.n38 171.744
R87 VDD2.n53 VDD2.n52 171.744
R88 VDD2.n52 VDD2.n42 171.744
R89 VDD2.n45 VDD2.n42 171.744
R90 VDD2.n10 VDD2.n7 171.744
R91 VDD2.n17 VDD2.n7 171.744
R92 VDD2.n18 VDD2.n17 171.744
R93 VDD2.n18 VDD2.n3 171.744
R94 VDD2.n25 VDD2.n3 171.744
R95 VDD2.n26 VDD2.n25 171.744
R96 VDD2.n34 VDD2.n33 91.5278
R97 VDD2 VDD2.n69 91.5249
R98 VDD2.n68 VDD2.n67 90.7427
R99 VDD2.n32 VDD2.n31 90.7426
R100 VDD2.n45 VDD2.t7 85.8723
R101 VDD2.n10 VDD2.t8 85.8723
R102 VDD2.n32 VDD2.n30 48.4333
R103 VDD2.n66 VDD2.n65 47.3126
R104 VDD2.n66 VDD2.n34 34.142
R105 VDD2.n46 VDD2.n44 16.3865
R106 VDD2.n11 VDD2.n9 16.3865
R107 VDD2.n47 VDD2.n43 12.8005
R108 VDD2.n12 VDD2.n8 12.8005
R109 VDD2.n51 VDD2.n50 12.0247
R110 VDD2.n16 VDD2.n15 12.0247
R111 VDD2.n54 VDD2.n41 11.249
R112 VDD2.n19 VDD2.n6 11.249
R113 VDD2.n55 VDD2.n39 10.4732
R114 VDD2.n20 VDD2.n4 10.4732
R115 VDD2.n59 VDD2.n58 9.69747
R116 VDD2.n24 VDD2.n23 9.69747
R117 VDD2.n65 VDD2.n64 9.45567
R118 VDD2.n30 VDD2.n29 9.45567
R119 VDD2.n64 VDD2.n63 9.3005
R120 VDD2.n37 VDD2.n36 9.3005
R121 VDD2.n58 VDD2.n57 9.3005
R122 VDD2.n56 VDD2.n55 9.3005
R123 VDD2.n41 VDD2.n40 9.3005
R124 VDD2.n50 VDD2.n49 9.3005
R125 VDD2.n48 VDD2.n47 9.3005
R126 VDD2.n29 VDD2.n28 9.3005
R127 VDD2.n2 VDD2.n1 9.3005
R128 VDD2.n23 VDD2.n22 9.3005
R129 VDD2.n21 VDD2.n20 9.3005
R130 VDD2.n6 VDD2.n5 9.3005
R131 VDD2.n15 VDD2.n14 9.3005
R132 VDD2.n13 VDD2.n12 9.3005
R133 VDD2.n62 VDD2.n37 8.92171
R134 VDD2.n27 VDD2.n2 8.92171
R135 VDD2.n63 VDD2.n35 8.14595
R136 VDD2.n28 VDD2.n0 8.14595
R137 VDD2.n65 VDD2.n35 5.81868
R138 VDD2.n30 VDD2.n0 5.81868
R139 VDD2.n69 VDD2.t5 5.49121
R140 VDD2.n69 VDD2.t1 5.49121
R141 VDD2.n67 VDD2.t4 5.49121
R142 VDD2.n67 VDD2.t3 5.49121
R143 VDD2.n33 VDD2.t6 5.49121
R144 VDD2.n33 VDD2.t2 5.49121
R145 VDD2.n31 VDD2.t9 5.49121
R146 VDD2.n31 VDD2.t0 5.49121
R147 VDD2.n63 VDD2.n62 5.04292
R148 VDD2.n28 VDD2.n27 5.04292
R149 VDD2.n59 VDD2.n37 4.26717
R150 VDD2.n24 VDD2.n2 4.26717
R151 VDD2.n48 VDD2.n44 3.71286
R152 VDD2.n13 VDD2.n9 3.71286
R153 VDD2.n58 VDD2.n39 3.49141
R154 VDD2.n23 VDD2.n4 3.49141
R155 VDD2.n55 VDD2.n54 2.71565
R156 VDD2.n20 VDD2.n19 2.71565
R157 VDD2.n51 VDD2.n41 1.93989
R158 VDD2.n16 VDD2.n6 1.93989
R159 VDD2.n50 VDD2.n43 1.16414
R160 VDD2.n15 VDD2.n8 1.16414
R161 VDD2.n68 VDD2.n66 1.12119
R162 VDD2.n47 VDD2.n46 0.388379
R163 VDD2.n12 VDD2.n11 0.388379
R164 VDD2 VDD2.n68 0.338862
R165 VDD2.n34 VDD2.n32 0.225326
R166 VDD2.n64 VDD2.n36 0.155672
R167 VDD2.n57 VDD2.n36 0.155672
R168 VDD2.n57 VDD2.n56 0.155672
R169 VDD2.n56 VDD2.n40 0.155672
R170 VDD2.n49 VDD2.n40 0.155672
R171 VDD2.n49 VDD2.n48 0.155672
R172 VDD2.n14 VDD2.n13 0.155672
R173 VDD2.n14 VDD2.n5 0.155672
R174 VDD2.n21 VDD2.n5 0.155672
R175 VDD2.n22 VDD2.n21 0.155672
R176 VDD2.n22 VDD2.n1 0.155672
R177 VDD2.n29 VDD2.n1 0.155672
R178 VTAIL.n136 VTAIL.n110 756.745
R179 VTAIL.n28 VTAIL.n2 756.745
R180 VTAIL.n104 VTAIL.n78 756.745
R181 VTAIL.n68 VTAIL.n42 756.745
R182 VTAIL.n121 VTAIL.n120 585
R183 VTAIL.n118 VTAIL.n117 585
R184 VTAIL.n127 VTAIL.n126 585
R185 VTAIL.n129 VTAIL.n128 585
R186 VTAIL.n114 VTAIL.n113 585
R187 VTAIL.n135 VTAIL.n134 585
R188 VTAIL.n137 VTAIL.n136 585
R189 VTAIL.n13 VTAIL.n12 585
R190 VTAIL.n10 VTAIL.n9 585
R191 VTAIL.n19 VTAIL.n18 585
R192 VTAIL.n21 VTAIL.n20 585
R193 VTAIL.n6 VTAIL.n5 585
R194 VTAIL.n27 VTAIL.n26 585
R195 VTAIL.n29 VTAIL.n28 585
R196 VTAIL.n105 VTAIL.n104 585
R197 VTAIL.n103 VTAIL.n102 585
R198 VTAIL.n82 VTAIL.n81 585
R199 VTAIL.n97 VTAIL.n96 585
R200 VTAIL.n95 VTAIL.n94 585
R201 VTAIL.n86 VTAIL.n85 585
R202 VTAIL.n89 VTAIL.n88 585
R203 VTAIL.n69 VTAIL.n68 585
R204 VTAIL.n67 VTAIL.n66 585
R205 VTAIL.n46 VTAIL.n45 585
R206 VTAIL.n61 VTAIL.n60 585
R207 VTAIL.n59 VTAIL.n58 585
R208 VTAIL.n50 VTAIL.n49 585
R209 VTAIL.n53 VTAIL.n52 585
R210 VTAIL.t8 VTAIL.n119 327.601
R211 VTAIL.t4 VTAIL.n11 327.601
R212 VTAIL.t2 VTAIL.n87 327.601
R213 VTAIL.t16 VTAIL.n51 327.601
R214 VTAIL.n120 VTAIL.n117 171.744
R215 VTAIL.n127 VTAIL.n117 171.744
R216 VTAIL.n128 VTAIL.n127 171.744
R217 VTAIL.n128 VTAIL.n113 171.744
R218 VTAIL.n135 VTAIL.n113 171.744
R219 VTAIL.n136 VTAIL.n135 171.744
R220 VTAIL.n12 VTAIL.n9 171.744
R221 VTAIL.n19 VTAIL.n9 171.744
R222 VTAIL.n20 VTAIL.n19 171.744
R223 VTAIL.n20 VTAIL.n5 171.744
R224 VTAIL.n27 VTAIL.n5 171.744
R225 VTAIL.n28 VTAIL.n27 171.744
R226 VTAIL.n104 VTAIL.n103 171.744
R227 VTAIL.n103 VTAIL.n81 171.744
R228 VTAIL.n96 VTAIL.n81 171.744
R229 VTAIL.n96 VTAIL.n95 171.744
R230 VTAIL.n95 VTAIL.n85 171.744
R231 VTAIL.n88 VTAIL.n85 171.744
R232 VTAIL.n68 VTAIL.n67 171.744
R233 VTAIL.n67 VTAIL.n45 171.744
R234 VTAIL.n60 VTAIL.n45 171.744
R235 VTAIL.n60 VTAIL.n59 171.744
R236 VTAIL.n59 VTAIL.n49 171.744
R237 VTAIL.n52 VTAIL.n49 171.744
R238 VTAIL.n120 VTAIL.t8 85.8723
R239 VTAIL.n12 VTAIL.t4 85.8723
R240 VTAIL.n88 VTAIL.t2 85.8723
R241 VTAIL.n52 VTAIL.t16 85.8723
R242 VTAIL.n77 VTAIL.n76 74.064
R243 VTAIL.n75 VTAIL.n74 74.064
R244 VTAIL.n41 VTAIL.n40 74.064
R245 VTAIL.n39 VTAIL.n38 74.064
R246 VTAIL.n143 VTAIL.n142 74.0638
R247 VTAIL.n1 VTAIL.n0 74.0638
R248 VTAIL.n35 VTAIL.n34 74.0638
R249 VTAIL.n37 VTAIL.n36 74.0638
R250 VTAIL.n141 VTAIL.n140 30.6338
R251 VTAIL.n33 VTAIL.n32 30.6338
R252 VTAIL.n109 VTAIL.n108 30.6338
R253 VTAIL.n73 VTAIL.n72 30.6338
R254 VTAIL.n39 VTAIL.n37 19.7117
R255 VTAIL.n141 VTAIL.n109 18.591
R256 VTAIL.n121 VTAIL.n119 16.3865
R257 VTAIL.n13 VTAIL.n11 16.3865
R258 VTAIL.n89 VTAIL.n87 16.3865
R259 VTAIL.n53 VTAIL.n51 16.3865
R260 VTAIL.n122 VTAIL.n118 12.8005
R261 VTAIL.n14 VTAIL.n10 12.8005
R262 VTAIL.n90 VTAIL.n86 12.8005
R263 VTAIL.n54 VTAIL.n50 12.8005
R264 VTAIL.n126 VTAIL.n125 12.0247
R265 VTAIL.n18 VTAIL.n17 12.0247
R266 VTAIL.n94 VTAIL.n93 12.0247
R267 VTAIL.n58 VTAIL.n57 12.0247
R268 VTAIL.n129 VTAIL.n116 11.249
R269 VTAIL.n21 VTAIL.n8 11.249
R270 VTAIL.n97 VTAIL.n84 11.249
R271 VTAIL.n61 VTAIL.n48 11.249
R272 VTAIL.n130 VTAIL.n114 10.4732
R273 VTAIL.n22 VTAIL.n6 10.4732
R274 VTAIL.n98 VTAIL.n82 10.4732
R275 VTAIL.n62 VTAIL.n46 10.4732
R276 VTAIL.n134 VTAIL.n133 9.69747
R277 VTAIL.n26 VTAIL.n25 9.69747
R278 VTAIL.n102 VTAIL.n101 9.69747
R279 VTAIL.n66 VTAIL.n65 9.69747
R280 VTAIL.n140 VTAIL.n139 9.45567
R281 VTAIL.n32 VTAIL.n31 9.45567
R282 VTAIL.n108 VTAIL.n107 9.45567
R283 VTAIL.n72 VTAIL.n71 9.45567
R284 VTAIL.n139 VTAIL.n138 9.3005
R285 VTAIL.n112 VTAIL.n111 9.3005
R286 VTAIL.n133 VTAIL.n132 9.3005
R287 VTAIL.n131 VTAIL.n130 9.3005
R288 VTAIL.n116 VTAIL.n115 9.3005
R289 VTAIL.n125 VTAIL.n124 9.3005
R290 VTAIL.n123 VTAIL.n122 9.3005
R291 VTAIL.n31 VTAIL.n30 9.3005
R292 VTAIL.n4 VTAIL.n3 9.3005
R293 VTAIL.n25 VTAIL.n24 9.3005
R294 VTAIL.n23 VTAIL.n22 9.3005
R295 VTAIL.n8 VTAIL.n7 9.3005
R296 VTAIL.n17 VTAIL.n16 9.3005
R297 VTAIL.n15 VTAIL.n14 9.3005
R298 VTAIL.n107 VTAIL.n106 9.3005
R299 VTAIL.n80 VTAIL.n79 9.3005
R300 VTAIL.n101 VTAIL.n100 9.3005
R301 VTAIL.n99 VTAIL.n98 9.3005
R302 VTAIL.n84 VTAIL.n83 9.3005
R303 VTAIL.n93 VTAIL.n92 9.3005
R304 VTAIL.n91 VTAIL.n90 9.3005
R305 VTAIL.n71 VTAIL.n70 9.3005
R306 VTAIL.n44 VTAIL.n43 9.3005
R307 VTAIL.n65 VTAIL.n64 9.3005
R308 VTAIL.n63 VTAIL.n62 9.3005
R309 VTAIL.n48 VTAIL.n47 9.3005
R310 VTAIL.n57 VTAIL.n56 9.3005
R311 VTAIL.n55 VTAIL.n54 9.3005
R312 VTAIL.n137 VTAIL.n112 8.92171
R313 VTAIL.n29 VTAIL.n4 8.92171
R314 VTAIL.n105 VTAIL.n80 8.92171
R315 VTAIL.n69 VTAIL.n44 8.92171
R316 VTAIL.n138 VTAIL.n110 8.14595
R317 VTAIL.n30 VTAIL.n2 8.14595
R318 VTAIL.n106 VTAIL.n78 8.14595
R319 VTAIL.n70 VTAIL.n42 8.14595
R320 VTAIL.n140 VTAIL.n110 5.81868
R321 VTAIL.n32 VTAIL.n2 5.81868
R322 VTAIL.n108 VTAIL.n78 5.81868
R323 VTAIL.n72 VTAIL.n42 5.81868
R324 VTAIL.n142 VTAIL.t9 5.49121
R325 VTAIL.n142 VTAIL.t14 5.49121
R326 VTAIL.n0 VTAIL.t10 5.49121
R327 VTAIL.n0 VTAIL.t17 5.49121
R328 VTAIL.n34 VTAIL.t5 5.49121
R329 VTAIL.n34 VTAIL.t6 5.49121
R330 VTAIL.n36 VTAIL.t18 5.49121
R331 VTAIL.n36 VTAIL.t7 5.49121
R332 VTAIL.n76 VTAIL.t1 5.49121
R333 VTAIL.n76 VTAIL.t0 5.49121
R334 VTAIL.n74 VTAIL.t3 5.49121
R335 VTAIL.n74 VTAIL.t19 5.49121
R336 VTAIL.n40 VTAIL.t15 5.49121
R337 VTAIL.n40 VTAIL.t12 5.49121
R338 VTAIL.n38 VTAIL.t13 5.49121
R339 VTAIL.n38 VTAIL.t11 5.49121
R340 VTAIL.n138 VTAIL.n137 5.04292
R341 VTAIL.n30 VTAIL.n29 5.04292
R342 VTAIL.n106 VTAIL.n105 5.04292
R343 VTAIL.n70 VTAIL.n69 5.04292
R344 VTAIL.n134 VTAIL.n112 4.26717
R345 VTAIL.n26 VTAIL.n4 4.26717
R346 VTAIL.n102 VTAIL.n80 4.26717
R347 VTAIL.n66 VTAIL.n44 4.26717
R348 VTAIL.n91 VTAIL.n87 3.71286
R349 VTAIL.n55 VTAIL.n51 3.71286
R350 VTAIL.n123 VTAIL.n119 3.71286
R351 VTAIL.n15 VTAIL.n11 3.71286
R352 VTAIL.n133 VTAIL.n114 3.49141
R353 VTAIL.n25 VTAIL.n6 3.49141
R354 VTAIL.n101 VTAIL.n82 3.49141
R355 VTAIL.n65 VTAIL.n46 3.49141
R356 VTAIL.n130 VTAIL.n129 2.71565
R357 VTAIL.n22 VTAIL.n21 2.71565
R358 VTAIL.n98 VTAIL.n97 2.71565
R359 VTAIL.n62 VTAIL.n61 2.71565
R360 VTAIL.n126 VTAIL.n116 1.93989
R361 VTAIL.n18 VTAIL.n8 1.93989
R362 VTAIL.n94 VTAIL.n84 1.93989
R363 VTAIL.n58 VTAIL.n48 1.93989
R364 VTAIL.n125 VTAIL.n118 1.16414
R365 VTAIL.n17 VTAIL.n10 1.16414
R366 VTAIL.n93 VTAIL.n86 1.16414
R367 VTAIL.n57 VTAIL.n50 1.16414
R368 VTAIL.n41 VTAIL.n39 1.12119
R369 VTAIL.n73 VTAIL.n41 1.12119
R370 VTAIL.n77 VTAIL.n75 1.12119
R371 VTAIL.n109 VTAIL.n77 1.12119
R372 VTAIL.n37 VTAIL.n35 1.12119
R373 VTAIL.n35 VTAIL.n33 1.12119
R374 VTAIL.n143 VTAIL.n141 1.12119
R375 VTAIL.n75 VTAIL.n73 1.03067
R376 VTAIL.n33 VTAIL.n1 1.03067
R377 VTAIL VTAIL.n1 0.899207
R378 VTAIL.n122 VTAIL.n121 0.388379
R379 VTAIL.n14 VTAIL.n13 0.388379
R380 VTAIL.n90 VTAIL.n89 0.388379
R381 VTAIL.n54 VTAIL.n53 0.388379
R382 VTAIL VTAIL.n143 0.222483
R383 VTAIL.n124 VTAIL.n123 0.155672
R384 VTAIL.n124 VTAIL.n115 0.155672
R385 VTAIL.n131 VTAIL.n115 0.155672
R386 VTAIL.n132 VTAIL.n131 0.155672
R387 VTAIL.n132 VTAIL.n111 0.155672
R388 VTAIL.n139 VTAIL.n111 0.155672
R389 VTAIL.n16 VTAIL.n15 0.155672
R390 VTAIL.n16 VTAIL.n7 0.155672
R391 VTAIL.n23 VTAIL.n7 0.155672
R392 VTAIL.n24 VTAIL.n23 0.155672
R393 VTAIL.n24 VTAIL.n3 0.155672
R394 VTAIL.n31 VTAIL.n3 0.155672
R395 VTAIL.n107 VTAIL.n79 0.155672
R396 VTAIL.n100 VTAIL.n79 0.155672
R397 VTAIL.n100 VTAIL.n99 0.155672
R398 VTAIL.n99 VTAIL.n83 0.155672
R399 VTAIL.n92 VTAIL.n83 0.155672
R400 VTAIL.n92 VTAIL.n91 0.155672
R401 VTAIL.n71 VTAIL.n43 0.155672
R402 VTAIL.n64 VTAIL.n43 0.155672
R403 VTAIL.n64 VTAIL.n63 0.155672
R404 VTAIL.n63 VTAIL.n47 0.155672
R405 VTAIL.n56 VTAIL.n47 0.155672
R406 VTAIL.n56 VTAIL.n55 0.155672
R407 B.n357 B.n50 585
R408 B.n359 B.n358 585
R409 B.n360 B.n49 585
R410 B.n362 B.n361 585
R411 B.n363 B.n48 585
R412 B.n365 B.n364 585
R413 B.n366 B.n47 585
R414 B.n368 B.n367 585
R415 B.n369 B.n46 585
R416 B.n371 B.n370 585
R417 B.n372 B.n45 585
R418 B.n374 B.n373 585
R419 B.n375 B.n44 585
R420 B.n377 B.n376 585
R421 B.n378 B.n43 585
R422 B.n380 B.n379 585
R423 B.n381 B.n42 585
R424 B.n383 B.n382 585
R425 B.n384 B.n41 585
R426 B.n386 B.n385 585
R427 B.n387 B.n40 585
R428 B.n389 B.n388 585
R429 B.n390 B.n39 585
R430 B.n392 B.n391 585
R431 B.n394 B.n393 585
R432 B.n395 B.n35 585
R433 B.n397 B.n396 585
R434 B.n398 B.n34 585
R435 B.n400 B.n399 585
R436 B.n401 B.n33 585
R437 B.n403 B.n402 585
R438 B.n404 B.n32 585
R439 B.n406 B.n405 585
R440 B.n408 B.n29 585
R441 B.n410 B.n409 585
R442 B.n411 B.n28 585
R443 B.n413 B.n412 585
R444 B.n414 B.n27 585
R445 B.n416 B.n415 585
R446 B.n417 B.n26 585
R447 B.n419 B.n418 585
R448 B.n420 B.n25 585
R449 B.n422 B.n421 585
R450 B.n423 B.n24 585
R451 B.n425 B.n424 585
R452 B.n426 B.n23 585
R453 B.n428 B.n427 585
R454 B.n429 B.n22 585
R455 B.n431 B.n430 585
R456 B.n432 B.n21 585
R457 B.n434 B.n433 585
R458 B.n435 B.n20 585
R459 B.n437 B.n436 585
R460 B.n438 B.n19 585
R461 B.n440 B.n439 585
R462 B.n441 B.n18 585
R463 B.n443 B.n442 585
R464 B.n356 B.n355 585
R465 B.n354 B.n51 585
R466 B.n353 B.n352 585
R467 B.n351 B.n52 585
R468 B.n350 B.n349 585
R469 B.n348 B.n53 585
R470 B.n347 B.n346 585
R471 B.n345 B.n54 585
R472 B.n344 B.n343 585
R473 B.n342 B.n55 585
R474 B.n341 B.n340 585
R475 B.n339 B.n56 585
R476 B.n338 B.n337 585
R477 B.n336 B.n57 585
R478 B.n335 B.n334 585
R479 B.n333 B.n58 585
R480 B.n332 B.n331 585
R481 B.n330 B.n59 585
R482 B.n329 B.n328 585
R483 B.n327 B.n60 585
R484 B.n326 B.n325 585
R485 B.n324 B.n61 585
R486 B.n323 B.n322 585
R487 B.n321 B.n62 585
R488 B.n320 B.n319 585
R489 B.n318 B.n63 585
R490 B.n317 B.n316 585
R491 B.n315 B.n64 585
R492 B.n314 B.n313 585
R493 B.n312 B.n65 585
R494 B.n311 B.n310 585
R495 B.n309 B.n66 585
R496 B.n308 B.n307 585
R497 B.n306 B.n67 585
R498 B.n305 B.n304 585
R499 B.n303 B.n68 585
R500 B.n302 B.n301 585
R501 B.n300 B.n69 585
R502 B.n299 B.n298 585
R503 B.n297 B.n70 585
R504 B.n296 B.n295 585
R505 B.n294 B.n71 585
R506 B.n293 B.n292 585
R507 B.n291 B.n72 585
R508 B.n290 B.n289 585
R509 B.n288 B.n73 585
R510 B.n287 B.n286 585
R511 B.n285 B.n74 585
R512 B.n284 B.n283 585
R513 B.n282 B.n75 585
R514 B.n281 B.n280 585
R515 B.n279 B.n76 585
R516 B.n278 B.n277 585
R517 B.n276 B.n77 585
R518 B.n275 B.n274 585
R519 B.n273 B.n78 585
R520 B.n272 B.n271 585
R521 B.n270 B.n79 585
R522 B.n269 B.n268 585
R523 B.n267 B.n80 585
R524 B.n266 B.n265 585
R525 B.n264 B.n81 585
R526 B.n263 B.n262 585
R527 B.n176 B.n175 585
R528 B.n177 B.n114 585
R529 B.n179 B.n178 585
R530 B.n180 B.n113 585
R531 B.n182 B.n181 585
R532 B.n183 B.n112 585
R533 B.n185 B.n184 585
R534 B.n186 B.n111 585
R535 B.n188 B.n187 585
R536 B.n189 B.n110 585
R537 B.n191 B.n190 585
R538 B.n192 B.n109 585
R539 B.n194 B.n193 585
R540 B.n195 B.n108 585
R541 B.n197 B.n196 585
R542 B.n198 B.n107 585
R543 B.n200 B.n199 585
R544 B.n201 B.n106 585
R545 B.n203 B.n202 585
R546 B.n204 B.n105 585
R547 B.n206 B.n205 585
R548 B.n207 B.n104 585
R549 B.n209 B.n208 585
R550 B.n210 B.n101 585
R551 B.n213 B.n212 585
R552 B.n214 B.n100 585
R553 B.n216 B.n215 585
R554 B.n217 B.n99 585
R555 B.n219 B.n218 585
R556 B.n220 B.n98 585
R557 B.n222 B.n221 585
R558 B.n223 B.n97 585
R559 B.n225 B.n224 585
R560 B.n227 B.n226 585
R561 B.n228 B.n93 585
R562 B.n230 B.n229 585
R563 B.n231 B.n92 585
R564 B.n233 B.n232 585
R565 B.n234 B.n91 585
R566 B.n236 B.n235 585
R567 B.n237 B.n90 585
R568 B.n239 B.n238 585
R569 B.n240 B.n89 585
R570 B.n242 B.n241 585
R571 B.n243 B.n88 585
R572 B.n245 B.n244 585
R573 B.n246 B.n87 585
R574 B.n248 B.n247 585
R575 B.n249 B.n86 585
R576 B.n251 B.n250 585
R577 B.n252 B.n85 585
R578 B.n254 B.n253 585
R579 B.n255 B.n84 585
R580 B.n257 B.n256 585
R581 B.n258 B.n83 585
R582 B.n260 B.n259 585
R583 B.n261 B.n82 585
R584 B.n174 B.n115 585
R585 B.n173 B.n172 585
R586 B.n171 B.n116 585
R587 B.n170 B.n169 585
R588 B.n168 B.n117 585
R589 B.n167 B.n166 585
R590 B.n165 B.n118 585
R591 B.n164 B.n163 585
R592 B.n162 B.n119 585
R593 B.n161 B.n160 585
R594 B.n159 B.n120 585
R595 B.n158 B.n157 585
R596 B.n156 B.n121 585
R597 B.n155 B.n154 585
R598 B.n153 B.n122 585
R599 B.n152 B.n151 585
R600 B.n150 B.n123 585
R601 B.n149 B.n148 585
R602 B.n147 B.n124 585
R603 B.n146 B.n145 585
R604 B.n144 B.n125 585
R605 B.n143 B.n142 585
R606 B.n141 B.n126 585
R607 B.n140 B.n139 585
R608 B.n138 B.n127 585
R609 B.n137 B.n136 585
R610 B.n135 B.n128 585
R611 B.n134 B.n133 585
R612 B.n132 B.n129 585
R613 B.n131 B.n130 585
R614 B.n2 B.n0 585
R615 B.n489 B.n1 585
R616 B.n488 B.n487 585
R617 B.n486 B.n3 585
R618 B.n485 B.n484 585
R619 B.n483 B.n4 585
R620 B.n482 B.n481 585
R621 B.n480 B.n5 585
R622 B.n479 B.n478 585
R623 B.n477 B.n6 585
R624 B.n476 B.n475 585
R625 B.n474 B.n7 585
R626 B.n473 B.n472 585
R627 B.n471 B.n8 585
R628 B.n470 B.n469 585
R629 B.n468 B.n9 585
R630 B.n467 B.n466 585
R631 B.n465 B.n10 585
R632 B.n464 B.n463 585
R633 B.n462 B.n11 585
R634 B.n461 B.n460 585
R635 B.n459 B.n12 585
R636 B.n458 B.n457 585
R637 B.n456 B.n13 585
R638 B.n455 B.n454 585
R639 B.n453 B.n14 585
R640 B.n452 B.n451 585
R641 B.n450 B.n15 585
R642 B.n449 B.n448 585
R643 B.n447 B.n16 585
R644 B.n446 B.n445 585
R645 B.n444 B.n17 585
R646 B.n491 B.n490 585
R647 B.n176 B.n115 511.721
R648 B.n442 B.n17 511.721
R649 B.n262 B.n261 511.721
R650 B.n357 B.n356 511.721
R651 B.n94 B.t9 349.803
R652 B.n102 B.t6 349.803
R653 B.n30 B.t3 349.803
R654 B.n36 B.t0 349.803
R655 B.n94 B.t11 291.853
R656 B.n36 B.t1 291.853
R657 B.n102 B.t8 291.853
R658 B.n30 B.t4 291.853
R659 B.n95 B.t10 266.642
R660 B.n37 B.t2 266.642
R661 B.n103 B.t7 266.642
R662 B.n31 B.t5 266.642
R663 B.n172 B.n115 163.367
R664 B.n172 B.n171 163.367
R665 B.n171 B.n170 163.367
R666 B.n170 B.n117 163.367
R667 B.n166 B.n117 163.367
R668 B.n166 B.n165 163.367
R669 B.n165 B.n164 163.367
R670 B.n164 B.n119 163.367
R671 B.n160 B.n119 163.367
R672 B.n160 B.n159 163.367
R673 B.n159 B.n158 163.367
R674 B.n158 B.n121 163.367
R675 B.n154 B.n121 163.367
R676 B.n154 B.n153 163.367
R677 B.n153 B.n152 163.367
R678 B.n152 B.n123 163.367
R679 B.n148 B.n123 163.367
R680 B.n148 B.n147 163.367
R681 B.n147 B.n146 163.367
R682 B.n146 B.n125 163.367
R683 B.n142 B.n125 163.367
R684 B.n142 B.n141 163.367
R685 B.n141 B.n140 163.367
R686 B.n140 B.n127 163.367
R687 B.n136 B.n127 163.367
R688 B.n136 B.n135 163.367
R689 B.n135 B.n134 163.367
R690 B.n134 B.n129 163.367
R691 B.n130 B.n129 163.367
R692 B.n130 B.n2 163.367
R693 B.n490 B.n2 163.367
R694 B.n490 B.n489 163.367
R695 B.n489 B.n488 163.367
R696 B.n488 B.n3 163.367
R697 B.n484 B.n3 163.367
R698 B.n484 B.n483 163.367
R699 B.n483 B.n482 163.367
R700 B.n482 B.n5 163.367
R701 B.n478 B.n5 163.367
R702 B.n478 B.n477 163.367
R703 B.n477 B.n476 163.367
R704 B.n476 B.n7 163.367
R705 B.n472 B.n7 163.367
R706 B.n472 B.n471 163.367
R707 B.n471 B.n470 163.367
R708 B.n470 B.n9 163.367
R709 B.n466 B.n9 163.367
R710 B.n466 B.n465 163.367
R711 B.n465 B.n464 163.367
R712 B.n464 B.n11 163.367
R713 B.n460 B.n11 163.367
R714 B.n460 B.n459 163.367
R715 B.n459 B.n458 163.367
R716 B.n458 B.n13 163.367
R717 B.n454 B.n13 163.367
R718 B.n454 B.n453 163.367
R719 B.n453 B.n452 163.367
R720 B.n452 B.n15 163.367
R721 B.n448 B.n15 163.367
R722 B.n448 B.n447 163.367
R723 B.n447 B.n446 163.367
R724 B.n446 B.n17 163.367
R725 B.n177 B.n176 163.367
R726 B.n178 B.n177 163.367
R727 B.n178 B.n113 163.367
R728 B.n182 B.n113 163.367
R729 B.n183 B.n182 163.367
R730 B.n184 B.n183 163.367
R731 B.n184 B.n111 163.367
R732 B.n188 B.n111 163.367
R733 B.n189 B.n188 163.367
R734 B.n190 B.n189 163.367
R735 B.n190 B.n109 163.367
R736 B.n194 B.n109 163.367
R737 B.n195 B.n194 163.367
R738 B.n196 B.n195 163.367
R739 B.n196 B.n107 163.367
R740 B.n200 B.n107 163.367
R741 B.n201 B.n200 163.367
R742 B.n202 B.n201 163.367
R743 B.n202 B.n105 163.367
R744 B.n206 B.n105 163.367
R745 B.n207 B.n206 163.367
R746 B.n208 B.n207 163.367
R747 B.n208 B.n101 163.367
R748 B.n213 B.n101 163.367
R749 B.n214 B.n213 163.367
R750 B.n215 B.n214 163.367
R751 B.n215 B.n99 163.367
R752 B.n219 B.n99 163.367
R753 B.n220 B.n219 163.367
R754 B.n221 B.n220 163.367
R755 B.n221 B.n97 163.367
R756 B.n225 B.n97 163.367
R757 B.n226 B.n225 163.367
R758 B.n226 B.n93 163.367
R759 B.n230 B.n93 163.367
R760 B.n231 B.n230 163.367
R761 B.n232 B.n231 163.367
R762 B.n232 B.n91 163.367
R763 B.n236 B.n91 163.367
R764 B.n237 B.n236 163.367
R765 B.n238 B.n237 163.367
R766 B.n238 B.n89 163.367
R767 B.n242 B.n89 163.367
R768 B.n243 B.n242 163.367
R769 B.n244 B.n243 163.367
R770 B.n244 B.n87 163.367
R771 B.n248 B.n87 163.367
R772 B.n249 B.n248 163.367
R773 B.n250 B.n249 163.367
R774 B.n250 B.n85 163.367
R775 B.n254 B.n85 163.367
R776 B.n255 B.n254 163.367
R777 B.n256 B.n255 163.367
R778 B.n256 B.n83 163.367
R779 B.n260 B.n83 163.367
R780 B.n261 B.n260 163.367
R781 B.n262 B.n81 163.367
R782 B.n266 B.n81 163.367
R783 B.n267 B.n266 163.367
R784 B.n268 B.n267 163.367
R785 B.n268 B.n79 163.367
R786 B.n272 B.n79 163.367
R787 B.n273 B.n272 163.367
R788 B.n274 B.n273 163.367
R789 B.n274 B.n77 163.367
R790 B.n278 B.n77 163.367
R791 B.n279 B.n278 163.367
R792 B.n280 B.n279 163.367
R793 B.n280 B.n75 163.367
R794 B.n284 B.n75 163.367
R795 B.n285 B.n284 163.367
R796 B.n286 B.n285 163.367
R797 B.n286 B.n73 163.367
R798 B.n290 B.n73 163.367
R799 B.n291 B.n290 163.367
R800 B.n292 B.n291 163.367
R801 B.n292 B.n71 163.367
R802 B.n296 B.n71 163.367
R803 B.n297 B.n296 163.367
R804 B.n298 B.n297 163.367
R805 B.n298 B.n69 163.367
R806 B.n302 B.n69 163.367
R807 B.n303 B.n302 163.367
R808 B.n304 B.n303 163.367
R809 B.n304 B.n67 163.367
R810 B.n308 B.n67 163.367
R811 B.n309 B.n308 163.367
R812 B.n310 B.n309 163.367
R813 B.n310 B.n65 163.367
R814 B.n314 B.n65 163.367
R815 B.n315 B.n314 163.367
R816 B.n316 B.n315 163.367
R817 B.n316 B.n63 163.367
R818 B.n320 B.n63 163.367
R819 B.n321 B.n320 163.367
R820 B.n322 B.n321 163.367
R821 B.n322 B.n61 163.367
R822 B.n326 B.n61 163.367
R823 B.n327 B.n326 163.367
R824 B.n328 B.n327 163.367
R825 B.n328 B.n59 163.367
R826 B.n332 B.n59 163.367
R827 B.n333 B.n332 163.367
R828 B.n334 B.n333 163.367
R829 B.n334 B.n57 163.367
R830 B.n338 B.n57 163.367
R831 B.n339 B.n338 163.367
R832 B.n340 B.n339 163.367
R833 B.n340 B.n55 163.367
R834 B.n344 B.n55 163.367
R835 B.n345 B.n344 163.367
R836 B.n346 B.n345 163.367
R837 B.n346 B.n53 163.367
R838 B.n350 B.n53 163.367
R839 B.n351 B.n350 163.367
R840 B.n352 B.n351 163.367
R841 B.n352 B.n51 163.367
R842 B.n356 B.n51 163.367
R843 B.n442 B.n441 163.367
R844 B.n441 B.n440 163.367
R845 B.n440 B.n19 163.367
R846 B.n436 B.n19 163.367
R847 B.n436 B.n435 163.367
R848 B.n435 B.n434 163.367
R849 B.n434 B.n21 163.367
R850 B.n430 B.n21 163.367
R851 B.n430 B.n429 163.367
R852 B.n429 B.n428 163.367
R853 B.n428 B.n23 163.367
R854 B.n424 B.n23 163.367
R855 B.n424 B.n423 163.367
R856 B.n423 B.n422 163.367
R857 B.n422 B.n25 163.367
R858 B.n418 B.n25 163.367
R859 B.n418 B.n417 163.367
R860 B.n417 B.n416 163.367
R861 B.n416 B.n27 163.367
R862 B.n412 B.n27 163.367
R863 B.n412 B.n411 163.367
R864 B.n411 B.n410 163.367
R865 B.n410 B.n29 163.367
R866 B.n405 B.n29 163.367
R867 B.n405 B.n404 163.367
R868 B.n404 B.n403 163.367
R869 B.n403 B.n33 163.367
R870 B.n399 B.n33 163.367
R871 B.n399 B.n398 163.367
R872 B.n398 B.n397 163.367
R873 B.n397 B.n35 163.367
R874 B.n393 B.n35 163.367
R875 B.n393 B.n392 163.367
R876 B.n392 B.n39 163.367
R877 B.n388 B.n39 163.367
R878 B.n388 B.n387 163.367
R879 B.n387 B.n386 163.367
R880 B.n386 B.n41 163.367
R881 B.n382 B.n41 163.367
R882 B.n382 B.n381 163.367
R883 B.n381 B.n380 163.367
R884 B.n380 B.n43 163.367
R885 B.n376 B.n43 163.367
R886 B.n376 B.n375 163.367
R887 B.n375 B.n374 163.367
R888 B.n374 B.n45 163.367
R889 B.n370 B.n45 163.367
R890 B.n370 B.n369 163.367
R891 B.n369 B.n368 163.367
R892 B.n368 B.n47 163.367
R893 B.n364 B.n47 163.367
R894 B.n364 B.n363 163.367
R895 B.n363 B.n362 163.367
R896 B.n362 B.n49 163.367
R897 B.n358 B.n49 163.367
R898 B.n358 B.n357 163.367
R899 B.n96 B.n95 59.5399
R900 B.n211 B.n103 59.5399
R901 B.n407 B.n31 59.5399
R902 B.n38 B.n37 59.5399
R903 B.n444 B.n443 33.2493
R904 B.n355 B.n50 33.2493
R905 B.n263 B.n82 33.2493
R906 B.n175 B.n174 33.2493
R907 B.n95 B.n94 25.2126
R908 B.n103 B.n102 25.2126
R909 B.n31 B.n30 25.2126
R910 B.n37 B.n36 25.2126
R911 B B.n491 18.0485
R912 B.n443 B.n18 10.6151
R913 B.n439 B.n18 10.6151
R914 B.n439 B.n438 10.6151
R915 B.n438 B.n437 10.6151
R916 B.n437 B.n20 10.6151
R917 B.n433 B.n20 10.6151
R918 B.n433 B.n432 10.6151
R919 B.n432 B.n431 10.6151
R920 B.n431 B.n22 10.6151
R921 B.n427 B.n22 10.6151
R922 B.n427 B.n426 10.6151
R923 B.n426 B.n425 10.6151
R924 B.n425 B.n24 10.6151
R925 B.n421 B.n24 10.6151
R926 B.n421 B.n420 10.6151
R927 B.n420 B.n419 10.6151
R928 B.n419 B.n26 10.6151
R929 B.n415 B.n26 10.6151
R930 B.n415 B.n414 10.6151
R931 B.n414 B.n413 10.6151
R932 B.n413 B.n28 10.6151
R933 B.n409 B.n28 10.6151
R934 B.n409 B.n408 10.6151
R935 B.n406 B.n32 10.6151
R936 B.n402 B.n32 10.6151
R937 B.n402 B.n401 10.6151
R938 B.n401 B.n400 10.6151
R939 B.n400 B.n34 10.6151
R940 B.n396 B.n34 10.6151
R941 B.n396 B.n395 10.6151
R942 B.n395 B.n394 10.6151
R943 B.n391 B.n390 10.6151
R944 B.n390 B.n389 10.6151
R945 B.n389 B.n40 10.6151
R946 B.n385 B.n40 10.6151
R947 B.n385 B.n384 10.6151
R948 B.n384 B.n383 10.6151
R949 B.n383 B.n42 10.6151
R950 B.n379 B.n42 10.6151
R951 B.n379 B.n378 10.6151
R952 B.n378 B.n377 10.6151
R953 B.n377 B.n44 10.6151
R954 B.n373 B.n44 10.6151
R955 B.n373 B.n372 10.6151
R956 B.n372 B.n371 10.6151
R957 B.n371 B.n46 10.6151
R958 B.n367 B.n46 10.6151
R959 B.n367 B.n366 10.6151
R960 B.n366 B.n365 10.6151
R961 B.n365 B.n48 10.6151
R962 B.n361 B.n48 10.6151
R963 B.n361 B.n360 10.6151
R964 B.n360 B.n359 10.6151
R965 B.n359 B.n50 10.6151
R966 B.n264 B.n263 10.6151
R967 B.n265 B.n264 10.6151
R968 B.n265 B.n80 10.6151
R969 B.n269 B.n80 10.6151
R970 B.n270 B.n269 10.6151
R971 B.n271 B.n270 10.6151
R972 B.n271 B.n78 10.6151
R973 B.n275 B.n78 10.6151
R974 B.n276 B.n275 10.6151
R975 B.n277 B.n276 10.6151
R976 B.n277 B.n76 10.6151
R977 B.n281 B.n76 10.6151
R978 B.n282 B.n281 10.6151
R979 B.n283 B.n282 10.6151
R980 B.n283 B.n74 10.6151
R981 B.n287 B.n74 10.6151
R982 B.n288 B.n287 10.6151
R983 B.n289 B.n288 10.6151
R984 B.n289 B.n72 10.6151
R985 B.n293 B.n72 10.6151
R986 B.n294 B.n293 10.6151
R987 B.n295 B.n294 10.6151
R988 B.n295 B.n70 10.6151
R989 B.n299 B.n70 10.6151
R990 B.n300 B.n299 10.6151
R991 B.n301 B.n300 10.6151
R992 B.n301 B.n68 10.6151
R993 B.n305 B.n68 10.6151
R994 B.n306 B.n305 10.6151
R995 B.n307 B.n306 10.6151
R996 B.n307 B.n66 10.6151
R997 B.n311 B.n66 10.6151
R998 B.n312 B.n311 10.6151
R999 B.n313 B.n312 10.6151
R1000 B.n313 B.n64 10.6151
R1001 B.n317 B.n64 10.6151
R1002 B.n318 B.n317 10.6151
R1003 B.n319 B.n318 10.6151
R1004 B.n319 B.n62 10.6151
R1005 B.n323 B.n62 10.6151
R1006 B.n324 B.n323 10.6151
R1007 B.n325 B.n324 10.6151
R1008 B.n325 B.n60 10.6151
R1009 B.n329 B.n60 10.6151
R1010 B.n330 B.n329 10.6151
R1011 B.n331 B.n330 10.6151
R1012 B.n331 B.n58 10.6151
R1013 B.n335 B.n58 10.6151
R1014 B.n336 B.n335 10.6151
R1015 B.n337 B.n336 10.6151
R1016 B.n337 B.n56 10.6151
R1017 B.n341 B.n56 10.6151
R1018 B.n342 B.n341 10.6151
R1019 B.n343 B.n342 10.6151
R1020 B.n343 B.n54 10.6151
R1021 B.n347 B.n54 10.6151
R1022 B.n348 B.n347 10.6151
R1023 B.n349 B.n348 10.6151
R1024 B.n349 B.n52 10.6151
R1025 B.n353 B.n52 10.6151
R1026 B.n354 B.n353 10.6151
R1027 B.n355 B.n354 10.6151
R1028 B.n175 B.n114 10.6151
R1029 B.n179 B.n114 10.6151
R1030 B.n180 B.n179 10.6151
R1031 B.n181 B.n180 10.6151
R1032 B.n181 B.n112 10.6151
R1033 B.n185 B.n112 10.6151
R1034 B.n186 B.n185 10.6151
R1035 B.n187 B.n186 10.6151
R1036 B.n187 B.n110 10.6151
R1037 B.n191 B.n110 10.6151
R1038 B.n192 B.n191 10.6151
R1039 B.n193 B.n192 10.6151
R1040 B.n193 B.n108 10.6151
R1041 B.n197 B.n108 10.6151
R1042 B.n198 B.n197 10.6151
R1043 B.n199 B.n198 10.6151
R1044 B.n199 B.n106 10.6151
R1045 B.n203 B.n106 10.6151
R1046 B.n204 B.n203 10.6151
R1047 B.n205 B.n204 10.6151
R1048 B.n205 B.n104 10.6151
R1049 B.n209 B.n104 10.6151
R1050 B.n210 B.n209 10.6151
R1051 B.n212 B.n100 10.6151
R1052 B.n216 B.n100 10.6151
R1053 B.n217 B.n216 10.6151
R1054 B.n218 B.n217 10.6151
R1055 B.n218 B.n98 10.6151
R1056 B.n222 B.n98 10.6151
R1057 B.n223 B.n222 10.6151
R1058 B.n224 B.n223 10.6151
R1059 B.n228 B.n227 10.6151
R1060 B.n229 B.n228 10.6151
R1061 B.n229 B.n92 10.6151
R1062 B.n233 B.n92 10.6151
R1063 B.n234 B.n233 10.6151
R1064 B.n235 B.n234 10.6151
R1065 B.n235 B.n90 10.6151
R1066 B.n239 B.n90 10.6151
R1067 B.n240 B.n239 10.6151
R1068 B.n241 B.n240 10.6151
R1069 B.n241 B.n88 10.6151
R1070 B.n245 B.n88 10.6151
R1071 B.n246 B.n245 10.6151
R1072 B.n247 B.n246 10.6151
R1073 B.n247 B.n86 10.6151
R1074 B.n251 B.n86 10.6151
R1075 B.n252 B.n251 10.6151
R1076 B.n253 B.n252 10.6151
R1077 B.n253 B.n84 10.6151
R1078 B.n257 B.n84 10.6151
R1079 B.n258 B.n257 10.6151
R1080 B.n259 B.n258 10.6151
R1081 B.n259 B.n82 10.6151
R1082 B.n174 B.n173 10.6151
R1083 B.n173 B.n116 10.6151
R1084 B.n169 B.n116 10.6151
R1085 B.n169 B.n168 10.6151
R1086 B.n168 B.n167 10.6151
R1087 B.n167 B.n118 10.6151
R1088 B.n163 B.n118 10.6151
R1089 B.n163 B.n162 10.6151
R1090 B.n162 B.n161 10.6151
R1091 B.n161 B.n120 10.6151
R1092 B.n157 B.n120 10.6151
R1093 B.n157 B.n156 10.6151
R1094 B.n156 B.n155 10.6151
R1095 B.n155 B.n122 10.6151
R1096 B.n151 B.n122 10.6151
R1097 B.n151 B.n150 10.6151
R1098 B.n150 B.n149 10.6151
R1099 B.n149 B.n124 10.6151
R1100 B.n145 B.n124 10.6151
R1101 B.n145 B.n144 10.6151
R1102 B.n144 B.n143 10.6151
R1103 B.n143 B.n126 10.6151
R1104 B.n139 B.n126 10.6151
R1105 B.n139 B.n138 10.6151
R1106 B.n138 B.n137 10.6151
R1107 B.n137 B.n128 10.6151
R1108 B.n133 B.n128 10.6151
R1109 B.n133 B.n132 10.6151
R1110 B.n132 B.n131 10.6151
R1111 B.n131 B.n0 10.6151
R1112 B.n487 B.n1 10.6151
R1113 B.n487 B.n486 10.6151
R1114 B.n486 B.n485 10.6151
R1115 B.n485 B.n4 10.6151
R1116 B.n481 B.n4 10.6151
R1117 B.n481 B.n480 10.6151
R1118 B.n480 B.n479 10.6151
R1119 B.n479 B.n6 10.6151
R1120 B.n475 B.n6 10.6151
R1121 B.n475 B.n474 10.6151
R1122 B.n474 B.n473 10.6151
R1123 B.n473 B.n8 10.6151
R1124 B.n469 B.n8 10.6151
R1125 B.n469 B.n468 10.6151
R1126 B.n468 B.n467 10.6151
R1127 B.n467 B.n10 10.6151
R1128 B.n463 B.n10 10.6151
R1129 B.n463 B.n462 10.6151
R1130 B.n462 B.n461 10.6151
R1131 B.n461 B.n12 10.6151
R1132 B.n457 B.n12 10.6151
R1133 B.n457 B.n456 10.6151
R1134 B.n456 B.n455 10.6151
R1135 B.n455 B.n14 10.6151
R1136 B.n451 B.n14 10.6151
R1137 B.n451 B.n450 10.6151
R1138 B.n450 B.n449 10.6151
R1139 B.n449 B.n16 10.6151
R1140 B.n445 B.n16 10.6151
R1141 B.n445 B.n444 10.6151
R1142 B.n407 B.n406 6.5566
R1143 B.n394 B.n38 6.5566
R1144 B.n212 B.n211 6.5566
R1145 B.n224 B.n96 6.5566
R1146 B.n408 B.n407 4.05904
R1147 B.n391 B.n38 4.05904
R1148 B.n211 B.n210 4.05904
R1149 B.n227 B.n96 4.05904
R1150 B.n491 B.n0 2.81026
R1151 B.n491 B.n1 2.81026
R1152 VP.n9 VP.t8 201.407
R1153 VP.n25 VP.t2 187.583
R1154 VP.n41 VP.t5 187.583
R1155 VP.n22 VP.t4 187.583
R1156 VP.n10 VP.n7 161.3
R1157 VP.n12 VP.n11 161.3
R1158 VP.n13 VP.n6 161.3
R1159 VP.n16 VP.n15 161.3
R1160 VP.n17 VP.n5 161.3
R1161 VP.n19 VP.n18 161.3
R1162 VP.n21 VP.n4 161.3
R1163 VP.n40 VP.n0 161.3
R1164 VP.n38 VP.n37 161.3
R1165 VP.n36 VP.n1 161.3
R1166 VP.n35 VP.n34 161.3
R1167 VP.n32 VP.n2 161.3
R1168 VP.n31 VP.n30 161.3
R1169 VP.n29 VP.n3 161.3
R1170 VP.n28 VP.n27 161.3
R1171 VP.n26 VP.t1 147.085
R1172 VP.n33 VP.t6 147.085
R1173 VP.n39 VP.t0 147.085
R1174 VP.n20 VP.t9 147.085
R1175 VP.n14 VP.t7 147.085
R1176 VP.n8 VP.t3 147.085
R1177 VP.n23 VP.n22 80.6037
R1178 VP.n42 VP.n41 80.6037
R1179 VP.n25 VP.n24 80.6037
R1180 VP.n32 VP.n31 50.2647
R1181 VP.n34 VP.n1 50.2647
R1182 VP.n15 VP.n5 50.2647
R1183 VP.n13 VP.n12 50.2647
R1184 VP.n27 VP.n25 49.9219
R1185 VP.n41 VP.n40 49.9219
R1186 VP.n22 VP.n21 49.9219
R1187 VP.n9 VP.n8 49.6998
R1188 VP.n10 VP.n9 44.8559
R1189 VP.n24 VP.n23 39.7438
R1190 VP.n31 VP.n3 30.8893
R1191 VP.n38 VP.n1 30.8893
R1192 VP.n19 VP.n5 30.8893
R1193 VP.n12 VP.n7 30.8893
R1194 VP.n27 VP.n26 22.1332
R1195 VP.n40 VP.n39 22.1332
R1196 VP.n21 VP.n20 22.1332
R1197 VP.n33 VP.n32 12.2964
R1198 VP.n34 VP.n33 12.2964
R1199 VP.n14 VP.n13 12.2964
R1200 VP.n15 VP.n14 12.2964
R1201 VP.n26 VP.n3 2.45968
R1202 VP.n39 VP.n38 2.45968
R1203 VP.n20 VP.n19 2.45968
R1204 VP.n8 VP.n7 2.45968
R1205 VP.n23 VP.n4 0.285035
R1206 VP.n28 VP.n24 0.285035
R1207 VP.n42 VP.n0 0.285035
R1208 VP.n11 VP.n10 0.189894
R1209 VP.n11 VP.n6 0.189894
R1210 VP.n16 VP.n6 0.189894
R1211 VP.n17 VP.n16 0.189894
R1212 VP.n18 VP.n17 0.189894
R1213 VP.n18 VP.n4 0.189894
R1214 VP.n29 VP.n28 0.189894
R1215 VP.n30 VP.n29 0.189894
R1216 VP.n30 VP.n2 0.189894
R1217 VP.n35 VP.n2 0.189894
R1218 VP.n36 VP.n35 0.189894
R1219 VP.n37 VP.n36 0.189894
R1220 VP.n37 VP.n0 0.189894
R1221 VP VP.n42 0.146778
R1222 VDD1.n26 VDD1.n0 756.745
R1223 VDD1.n59 VDD1.n33 756.745
R1224 VDD1.n27 VDD1.n26 585
R1225 VDD1.n25 VDD1.n24 585
R1226 VDD1.n4 VDD1.n3 585
R1227 VDD1.n19 VDD1.n18 585
R1228 VDD1.n17 VDD1.n16 585
R1229 VDD1.n8 VDD1.n7 585
R1230 VDD1.n11 VDD1.n10 585
R1231 VDD1.n44 VDD1.n43 585
R1232 VDD1.n41 VDD1.n40 585
R1233 VDD1.n50 VDD1.n49 585
R1234 VDD1.n52 VDD1.n51 585
R1235 VDD1.n37 VDD1.n36 585
R1236 VDD1.n58 VDD1.n57 585
R1237 VDD1.n60 VDD1.n59 585
R1238 VDD1.t1 VDD1.n9 327.601
R1239 VDD1.t7 VDD1.n42 327.601
R1240 VDD1.n26 VDD1.n25 171.744
R1241 VDD1.n25 VDD1.n3 171.744
R1242 VDD1.n18 VDD1.n3 171.744
R1243 VDD1.n18 VDD1.n17 171.744
R1244 VDD1.n17 VDD1.n7 171.744
R1245 VDD1.n10 VDD1.n7 171.744
R1246 VDD1.n43 VDD1.n40 171.744
R1247 VDD1.n50 VDD1.n40 171.744
R1248 VDD1.n51 VDD1.n50 171.744
R1249 VDD1.n51 VDD1.n36 171.744
R1250 VDD1.n58 VDD1.n36 171.744
R1251 VDD1.n59 VDD1.n58 171.744
R1252 VDD1.n67 VDD1.n66 91.5278
R1253 VDD1.n32 VDD1.n31 90.7427
R1254 VDD1.n69 VDD1.n68 90.7426
R1255 VDD1.n65 VDD1.n64 90.7426
R1256 VDD1.n10 VDD1.t1 85.8723
R1257 VDD1.n43 VDD1.t7 85.8723
R1258 VDD1.n32 VDD1.n30 48.4333
R1259 VDD1.n65 VDD1.n63 48.4333
R1260 VDD1.n69 VDD1.n67 35.2854
R1261 VDD1.n11 VDD1.n9 16.3865
R1262 VDD1.n44 VDD1.n42 16.3865
R1263 VDD1.n12 VDD1.n8 12.8005
R1264 VDD1.n45 VDD1.n41 12.8005
R1265 VDD1.n16 VDD1.n15 12.0247
R1266 VDD1.n49 VDD1.n48 12.0247
R1267 VDD1.n19 VDD1.n6 11.249
R1268 VDD1.n52 VDD1.n39 11.249
R1269 VDD1.n20 VDD1.n4 10.4732
R1270 VDD1.n53 VDD1.n37 10.4732
R1271 VDD1.n24 VDD1.n23 9.69747
R1272 VDD1.n57 VDD1.n56 9.69747
R1273 VDD1.n30 VDD1.n29 9.45567
R1274 VDD1.n63 VDD1.n62 9.45567
R1275 VDD1.n29 VDD1.n28 9.3005
R1276 VDD1.n2 VDD1.n1 9.3005
R1277 VDD1.n23 VDD1.n22 9.3005
R1278 VDD1.n21 VDD1.n20 9.3005
R1279 VDD1.n6 VDD1.n5 9.3005
R1280 VDD1.n15 VDD1.n14 9.3005
R1281 VDD1.n13 VDD1.n12 9.3005
R1282 VDD1.n62 VDD1.n61 9.3005
R1283 VDD1.n35 VDD1.n34 9.3005
R1284 VDD1.n56 VDD1.n55 9.3005
R1285 VDD1.n54 VDD1.n53 9.3005
R1286 VDD1.n39 VDD1.n38 9.3005
R1287 VDD1.n48 VDD1.n47 9.3005
R1288 VDD1.n46 VDD1.n45 9.3005
R1289 VDD1.n27 VDD1.n2 8.92171
R1290 VDD1.n60 VDD1.n35 8.92171
R1291 VDD1.n28 VDD1.n0 8.14595
R1292 VDD1.n61 VDD1.n33 8.14595
R1293 VDD1.n30 VDD1.n0 5.81868
R1294 VDD1.n63 VDD1.n33 5.81868
R1295 VDD1.n68 VDD1.t0 5.49121
R1296 VDD1.n68 VDD1.t5 5.49121
R1297 VDD1.n31 VDD1.t6 5.49121
R1298 VDD1.n31 VDD1.t2 5.49121
R1299 VDD1.n66 VDD1.t9 5.49121
R1300 VDD1.n66 VDD1.t4 5.49121
R1301 VDD1.n64 VDD1.t8 5.49121
R1302 VDD1.n64 VDD1.t3 5.49121
R1303 VDD1.n28 VDD1.n27 5.04292
R1304 VDD1.n61 VDD1.n60 5.04292
R1305 VDD1.n24 VDD1.n2 4.26717
R1306 VDD1.n57 VDD1.n35 4.26717
R1307 VDD1.n13 VDD1.n9 3.71286
R1308 VDD1.n46 VDD1.n42 3.71286
R1309 VDD1.n23 VDD1.n4 3.49141
R1310 VDD1.n56 VDD1.n37 3.49141
R1311 VDD1.n20 VDD1.n19 2.71565
R1312 VDD1.n53 VDD1.n52 2.71565
R1313 VDD1.n16 VDD1.n6 1.93989
R1314 VDD1.n49 VDD1.n39 1.93989
R1315 VDD1.n15 VDD1.n8 1.16414
R1316 VDD1.n48 VDD1.n41 1.16414
R1317 VDD1 VDD1.n69 0.782828
R1318 VDD1.n12 VDD1.n11 0.388379
R1319 VDD1.n45 VDD1.n44 0.388379
R1320 VDD1 VDD1.n32 0.338862
R1321 VDD1.n67 VDD1.n65 0.225326
R1322 VDD1.n29 VDD1.n1 0.155672
R1323 VDD1.n22 VDD1.n1 0.155672
R1324 VDD1.n22 VDD1.n21 0.155672
R1325 VDD1.n21 VDD1.n5 0.155672
R1326 VDD1.n14 VDD1.n5 0.155672
R1327 VDD1.n14 VDD1.n13 0.155672
R1328 VDD1.n47 VDD1.n46 0.155672
R1329 VDD1.n47 VDD1.n38 0.155672
R1330 VDD1.n54 VDD1.n38 0.155672
R1331 VDD1.n55 VDD1.n54 0.155672
R1332 VDD1.n55 VDD1.n34 0.155672
R1333 VDD1.n62 VDD1.n34 0.155672
C0 VN VDD1 0.149975f
C1 VDD2 B 1.42392f
C2 w_n2530_n2152# VP 5.12809f
C3 VN B 0.796564f
C4 w_n2530_n2152# VTAIL 2.10336f
C5 w_n2530_n2152# VDD1 1.71302f
C6 VN VDD2 4.09663f
C7 VP VDD1 4.31952f
C8 VP VTAIL 4.39958f
C9 VDD1 VTAIL 7.58237f
C10 w_n2530_n2152# B 6.10623f
C11 VP B 1.33301f
C12 w_n2530_n2152# VDD2 1.77184f
C13 VTAIL B 1.76343f
C14 VDD1 B 1.36928f
C15 VP VDD2 0.375416f
C16 w_n2530_n2152# VN 4.80372f
C17 VDD2 VDD1 1.14095f
C18 VDD2 VTAIL 7.62224f
C19 VP VN 4.86886f
C20 VN VTAIL 4.38526f
C21 VDD2 VSUBS 1.194753f
C22 VDD1 VSUBS 1.062166f
C23 VTAIL VSUBS 0.481893f
C24 VN VSUBS 4.85271f
C25 VP VSUBS 1.853449f
C26 B VSUBS 2.828804f
C27 w_n2530_n2152# VSUBS 67.976f
C28 VDD1.n0 VSUBS 0.025186f
C29 VDD1.n1 VSUBS 0.023744f
C30 VDD1.n2 VSUBS 0.012759f
C31 VDD1.n3 VSUBS 0.030158f
C32 VDD1.n4 VSUBS 0.01351f
C33 VDD1.n5 VSUBS 0.023744f
C34 VDD1.n6 VSUBS 0.012759f
C35 VDD1.n7 VSUBS 0.030158f
C36 VDD1.n8 VSUBS 0.01351f
C37 VDD1.n9 VSUBS 0.104323f
C38 VDD1.t1 VSUBS 0.064605f
C39 VDD1.n10 VSUBS 0.022619f
C40 VDD1.n11 VSUBS 0.019175f
C41 VDD1.n12 VSUBS 0.012759f
C42 VDD1.n13 VSUBS 0.536263f
C43 VDD1.n14 VSUBS 0.023744f
C44 VDD1.n15 VSUBS 0.012759f
C45 VDD1.n16 VSUBS 0.01351f
C46 VDD1.n17 VSUBS 0.030158f
C47 VDD1.n18 VSUBS 0.030158f
C48 VDD1.n19 VSUBS 0.01351f
C49 VDD1.n20 VSUBS 0.012759f
C50 VDD1.n21 VSUBS 0.023744f
C51 VDD1.n22 VSUBS 0.023744f
C52 VDD1.n23 VSUBS 0.012759f
C53 VDD1.n24 VSUBS 0.01351f
C54 VDD1.n25 VSUBS 0.030158f
C55 VDD1.n26 VSUBS 0.069929f
C56 VDD1.n27 VSUBS 0.01351f
C57 VDD1.n28 VSUBS 0.012759f
C58 VDD1.n29 VSUBS 0.052289f
C59 VDD1.n30 VSUBS 0.054373f
C60 VDD1.t6 VSUBS 0.111081f
C61 VDD1.t2 VSUBS 0.111081f
C62 VDD1.n31 VSUBS 0.731017f
C63 VDD1.n32 VSUBS 0.624957f
C64 VDD1.n33 VSUBS 0.025186f
C65 VDD1.n34 VSUBS 0.023744f
C66 VDD1.n35 VSUBS 0.012759f
C67 VDD1.n36 VSUBS 0.030158f
C68 VDD1.n37 VSUBS 0.01351f
C69 VDD1.n38 VSUBS 0.023744f
C70 VDD1.n39 VSUBS 0.012759f
C71 VDD1.n40 VSUBS 0.030158f
C72 VDD1.n41 VSUBS 0.01351f
C73 VDD1.n42 VSUBS 0.104323f
C74 VDD1.t7 VSUBS 0.064605f
C75 VDD1.n43 VSUBS 0.022619f
C76 VDD1.n44 VSUBS 0.019175f
C77 VDD1.n45 VSUBS 0.012759f
C78 VDD1.n46 VSUBS 0.536264f
C79 VDD1.n47 VSUBS 0.023744f
C80 VDD1.n48 VSUBS 0.012759f
C81 VDD1.n49 VSUBS 0.01351f
C82 VDD1.n50 VSUBS 0.030158f
C83 VDD1.n51 VSUBS 0.030158f
C84 VDD1.n52 VSUBS 0.01351f
C85 VDD1.n53 VSUBS 0.012759f
C86 VDD1.n54 VSUBS 0.023744f
C87 VDD1.n55 VSUBS 0.023744f
C88 VDD1.n56 VSUBS 0.012759f
C89 VDD1.n57 VSUBS 0.01351f
C90 VDD1.n58 VSUBS 0.030158f
C91 VDD1.n59 VSUBS 0.069929f
C92 VDD1.n60 VSUBS 0.01351f
C93 VDD1.n61 VSUBS 0.012759f
C94 VDD1.n62 VSUBS 0.052289f
C95 VDD1.n63 VSUBS 0.054373f
C96 VDD1.t8 VSUBS 0.111081f
C97 VDD1.t3 VSUBS 0.111081f
C98 VDD1.n64 VSUBS 0.731013f
C99 VDD1.n65 VSUBS 0.618722f
C100 VDD1.t9 VSUBS 0.111081f
C101 VDD1.t4 VSUBS 0.111081f
C102 VDD1.n66 VSUBS 0.735666f
C103 VDD1.n67 VSUBS 1.86666f
C104 VDD1.t0 VSUBS 0.111081f
C105 VDD1.t5 VSUBS 0.111081f
C106 VDD1.n68 VSUBS 0.731013f
C107 VDD1.n69 VSUBS 2.10926f
C108 VP.n0 VSUBS 0.072854f
C109 VP.t0 VSUBS 0.829164f
C110 VP.n1 VSUBS 0.051478f
C111 VP.n2 VSUBS 0.054598f
C112 VP.t6 VSUBS 0.829164f
C113 VP.n3 VSUBS 0.063802f
C114 VP.n4 VSUBS 0.072854f
C115 VP.t4 VSUBS 0.909805f
C116 VP.t9 VSUBS 0.829164f
C117 VP.n5 VSUBS 0.051478f
C118 VP.n6 VSUBS 0.054598f
C119 VP.t7 VSUBS 0.829164f
C120 VP.n7 VSUBS 0.063802f
C121 VP.t3 VSUBS 0.829164f
C122 VP.n8 VSUBS 0.378287f
C123 VP.t8 VSUBS 0.93868f
C124 VP.n9 VSUBS 0.420967f
C125 VP.n10 VSUBS 0.22306f
C126 VP.n11 VSUBS 0.054598f
C127 VP.n12 VSUBS 0.051478f
C128 VP.n13 VSUBS 0.074723f
C129 VP.n14 VSUBS 0.342862f
C130 VP.n15 VSUBS 0.074723f
C131 VP.n16 VSUBS 0.054598f
C132 VP.n17 VSUBS 0.054598f
C133 VP.n18 VSUBS 0.054598f
C134 VP.n19 VSUBS 0.063802f
C135 VP.n20 VSUBS 0.342862f
C136 VP.n21 VSUBS 0.063868f
C137 VP.n22 VSUBS 0.420346f
C138 VP.n23 VSUBS 2.07116f
C139 VP.n24 VSUBS 2.12069f
C140 VP.t2 VSUBS 0.909805f
C141 VP.n25 VSUBS 0.420346f
C142 VP.t1 VSUBS 0.829164f
C143 VP.n26 VSUBS 0.342862f
C144 VP.n27 VSUBS 0.063868f
C145 VP.n28 VSUBS 0.072854f
C146 VP.n29 VSUBS 0.054598f
C147 VP.n30 VSUBS 0.054598f
C148 VP.n31 VSUBS 0.051478f
C149 VP.n32 VSUBS 0.074723f
C150 VP.n33 VSUBS 0.342862f
C151 VP.n34 VSUBS 0.074723f
C152 VP.n35 VSUBS 0.054598f
C153 VP.n36 VSUBS 0.054598f
C154 VP.n37 VSUBS 0.054598f
C155 VP.n38 VSUBS 0.063802f
C156 VP.n39 VSUBS 0.342862f
C157 VP.n40 VSUBS 0.063868f
C158 VP.t5 VSUBS 0.909805f
C159 VP.n41 VSUBS 0.420346f
C160 VP.n42 VSUBS 0.051133f
C161 B.n0 VSUBS 0.004063f
C162 B.n1 VSUBS 0.004063f
C163 B.n2 VSUBS 0.006426f
C164 B.n3 VSUBS 0.006426f
C165 B.n4 VSUBS 0.006426f
C166 B.n5 VSUBS 0.006426f
C167 B.n6 VSUBS 0.006426f
C168 B.n7 VSUBS 0.006426f
C169 B.n8 VSUBS 0.006426f
C170 B.n9 VSUBS 0.006426f
C171 B.n10 VSUBS 0.006426f
C172 B.n11 VSUBS 0.006426f
C173 B.n12 VSUBS 0.006426f
C174 B.n13 VSUBS 0.006426f
C175 B.n14 VSUBS 0.006426f
C176 B.n15 VSUBS 0.006426f
C177 B.n16 VSUBS 0.006426f
C178 B.n17 VSUBS 0.014841f
C179 B.n18 VSUBS 0.006426f
C180 B.n19 VSUBS 0.006426f
C181 B.n20 VSUBS 0.006426f
C182 B.n21 VSUBS 0.006426f
C183 B.n22 VSUBS 0.006426f
C184 B.n23 VSUBS 0.006426f
C185 B.n24 VSUBS 0.006426f
C186 B.n25 VSUBS 0.006426f
C187 B.n26 VSUBS 0.006426f
C188 B.n27 VSUBS 0.006426f
C189 B.n28 VSUBS 0.006426f
C190 B.n29 VSUBS 0.006426f
C191 B.t5 VSUBS 0.080724f
C192 B.t4 VSUBS 0.091696f
C193 B.t3 VSUBS 0.234274f
C194 B.n30 VSUBS 0.161359f
C195 B.n31 VSUBS 0.13617f
C196 B.n32 VSUBS 0.006426f
C197 B.n33 VSUBS 0.006426f
C198 B.n34 VSUBS 0.006426f
C199 B.n35 VSUBS 0.006426f
C200 B.t2 VSUBS 0.080726f
C201 B.t1 VSUBS 0.091697f
C202 B.t0 VSUBS 0.234274f
C203 B.n36 VSUBS 0.161358f
C204 B.n37 VSUBS 0.136168f
C205 B.n38 VSUBS 0.014887f
C206 B.n39 VSUBS 0.006426f
C207 B.n40 VSUBS 0.006426f
C208 B.n41 VSUBS 0.006426f
C209 B.n42 VSUBS 0.006426f
C210 B.n43 VSUBS 0.006426f
C211 B.n44 VSUBS 0.006426f
C212 B.n45 VSUBS 0.006426f
C213 B.n46 VSUBS 0.006426f
C214 B.n47 VSUBS 0.006426f
C215 B.n48 VSUBS 0.006426f
C216 B.n49 VSUBS 0.006426f
C217 B.n50 VSUBS 0.014841f
C218 B.n51 VSUBS 0.006426f
C219 B.n52 VSUBS 0.006426f
C220 B.n53 VSUBS 0.006426f
C221 B.n54 VSUBS 0.006426f
C222 B.n55 VSUBS 0.006426f
C223 B.n56 VSUBS 0.006426f
C224 B.n57 VSUBS 0.006426f
C225 B.n58 VSUBS 0.006426f
C226 B.n59 VSUBS 0.006426f
C227 B.n60 VSUBS 0.006426f
C228 B.n61 VSUBS 0.006426f
C229 B.n62 VSUBS 0.006426f
C230 B.n63 VSUBS 0.006426f
C231 B.n64 VSUBS 0.006426f
C232 B.n65 VSUBS 0.006426f
C233 B.n66 VSUBS 0.006426f
C234 B.n67 VSUBS 0.006426f
C235 B.n68 VSUBS 0.006426f
C236 B.n69 VSUBS 0.006426f
C237 B.n70 VSUBS 0.006426f
C238 B.n71 VSUBS 0.006426f
C239 B.n72 VSUBS 0.006426f
C240 B.n73 VSUBS 0.006426f
C241 B.n74 VSUBS 0.006426f
C242 B.n75 VSUBS 0.006426f
C243 B.n76 VSUBS 0.006426f
C244 B.n77 VSUBS 0.006426f
C245 B.n78 VSUBS 0.006426f
C246 B.n79 VSUBS 0.006426f
C247 B.n80 VSUBS 0.006426f
C248 B.n81 VSUBS 0.006426f
C249 B.n82 VSUBS 0.015586f
C250 B.n83 VSUBS 0.006426f
C251 B.n84 VSUBS 0.006426f
C252 B.n85 VSUBS 0.006426f
C253 B.n86 VSUBS 0.006426f
C254 B.n87 VSUBS 0.006426f
C255 B.n88 VSUBS 0.006426f
C256 B.n89 VSUBS 0.006426f
C257 B.n90 VSUBS 0.006426f
C258 B.n91 VSUBS 0.006426f
C259 B.n92 VSUBS 0.006426f
C260 B.n93 VSUBS 0.006426f
C261 B.t10 VSUBS 0.080726f
C262 B.t11 VSUBS 0.091697f
C263 B.t9 VSUBS 0.234274f
C264 B.n94 VSUBS 0.161358f
C265 B.n95 VSUBS 0.136168f
C266 B.n96 VSUBS 0.014887f
C267 B.n97 VSUBS 0.006426f
C268 B.n98 VSUBS 0.006426f
C269 B.n99 VSUBS 0.006426f
C270 B.n100 VSUBS 0.006426f
C271 B.n101 VSUBS 0.006426f
C272 B.t7 VSUBS 0.080724f
C273 B.t8 VSUBS 0.091696f
C274 B.t6 VSUBS 0.234274f
C275 B.n102 VSUBS 0.161359f
C276 B.n103 VSUBS 0.13617f
C277 B.n104 VSUBS 0.006426f
C278 B.n105 VSUBS 0.006426f
C279 B.n106 VSUBS 0.006426f
C280 B.n107 VSUBS 0.006426f
C281 B.n108 VSUBS 0.006426f
C282 B.n109 VSUBS 0.006426f
C283 B.n110 VSUBS 0.006426f
C284 B.n111 VSUBS 0.006426f
C285 B.n112 VSUBS 0.006426f
C286 B.n113 VSUBS 0.006426f
C287 B.n114 VSUBS 0.006426f
C288 B.n115 VSUBS 0.014841f
C289 B.n116 VSUBS 0.006426f
C290 B.n117 VSUBS 0.006426f
C291 B.n118 VSUBS 0.006426f
C292 B.n119 VSUBS 0.006426f
C293 B.n120 VSUBS 0.006426f
C294 B.n121 VSUBS 0.006426f
C295 B.n122 VSUBS 0.006426f
C296 B.n123 VSUBS 0.006426f
C297 B.n124 VSUBS 0.006426f
C298 B.n125 VSUBS 0.006426f
C299 B.n126 VSUBS 0.006426f
C300 B.n127 VSUBS 0.006426f
C301 B.n128 VSUBS 0.006426f
C302 B.n129 VSUBS 0.006426f
C303 B.n130 VSUBS 0.006426f
C304 B.n131 VSUBS 0.006426f
C305 B.n132 VSUBS 0.006426f
C306 B.n133 VSUBS 0.006426f
C307 B.n134 VSUBS 0.006426f
C308 B.n135 VSUBS 0.006426f
C309 B.n136 VSUBS 0.006426f
C310 B.n137 VSUBS 0.006426f
C311 B.n138 VSUBS 0.006426f
C312 B.n139 VSUBS 0.006426f
C313 B.n140 VSUBS 0.006426f
C314 B.n141 VSUBS 0.006426f
C315 B.n142 VSUBS 0.006426f
C316 B.n143 VSUBS 0.006426f
C317 B.n144 VSUBS 0.006426f
C318 B.n145 VSUBS 0.006426f
C319 B.n146 VSUBS 0.006426f
C320 B.n147 VSUBS 0.006426f
C321 B.n148 VSUBS 0.006426f
C322 B.n149 VSUBS 0.006426f
C323 B.n150 VSUBS 0.006426f
C324 B.n151 VSUBS 0.006426f
C325 B.n152 VSUBS 0.006426f
C326 B.n153 VSUBS 0.006426f
C327 B.n154 VSUBS 0.006426f
C328 B.n155 VSUBS 0.006426f
C329 B.n156 VSUBS 0.006426f
C330 B.n157 VSUBS 0.006426f
C331 B.n158 VSUBS 0.006426f
C332 B.n159 VSUBS 0.006426f
C333 B.n160 VSUBS 0.006426f
C334 B.n161 VSUBS 0.006426f
C335 B.n162 VSUBS 0.006426f
C336 B.n163 VSUBS 0.006426f
C337 B.n164 VSUBS 0.006426f
C338 B.n165 VSUBS 0.006426f
C339 B.n166 VSUBS 0.006426f
C340 B.n167 VSUBS 0.006426f
C341 B.n168 VSUBS 0.006426f
C342 B.n169 VSUBS 0.006426f
C343 B.n170 VSUBS 0.006426f
C344 B.n171 VSUBS 0.006426f
C345 B.n172 VSUBS 0.006426f
C346 B.n173 VSUBS 0.006426f
C347 B.n174 VSUBS 0.014841f
C348 B.n175 VSUBS 0.015586f
C349 B.n176 VSUBS 0.015586f
C350 B.n177 VSUBS 0.006426f
C351 B.n178 VSUBS 0.006426f
C352 B.n179 VSUBS 0.006426f
C353 B.n180 VSUBS 0.006426f
C354 B.n181 VSUBS 0.006426f
C355 B.n182 VSUBS 0.006426f
C356 B.n183 VSUBS 0.006426f
C357 B.n184 VSUBS 0.006426f
C358 B.n185 VSUBS 0.006426f
C359 B.n186 VSUBS 0.006426f
C360 B.n187 VSUBS 0.006426f
C361 B.n188 VSUBS 0.006426f
C362 B.n189 VSUBS 0.006426f
C363 B.n190 VSUBS 0.006426f
C364 B.n191 VSUBS 0.006426f
C365 B.n192 VSUBS 0.006426f
C366 B.n193 VSUBS 0.006426f
C367 B.n194 VSUBS 0.006426f
C368 B.n195 VSUBS 0.006426f
C369 B.n196 VSUBS 0.006426f
C370 B.n197 VSUBS 0.006426f
C371 B.n198 VSUBS 0.006426f
C372 B.n199 VSUBS 0.006426f
C373 B.n200 VSUBS 0.006426f
C374 B.n201 VSUBS 0.006426f
C375 B.n202 VSUBS 0.006426f
C376 B.n203 VSUBS 0.006426f
C377 B.n204 VSUBS 0.006426f
C378 B.n205 VSUBS 0.006426f
C379 B.n206 VSUBS 0.006426f
C380 B.n207 VSUBS 0.006426f
C381 B.n208 VSUBS 0.006426f
C382 B.n209 VSUBS 0.006426f
C383 B.n210 VSUBS 0.004441f
C384 B.n211 VSUBS 0.014887f
C385 B.n212 VSUBS 0.005197f
C386 B.n213 VSUBS 0.006426f
C387 B.n214 VSUBS 0.006426f
C388 B.n215 VSUBS 0.006426f
C389 B.n216 VSUBS 0.006426f
C390 B.n217 VSUBS 0.006426f
C391 B.n218 VSUBS 0.006426f
C392 B.n219 VSUBS 0.006426f
C393 B.n220 VSUBS 0.006426f
C394 B.n221 VSUBS 0.006426f
C395 B.n222 VSUBS 0.006426f
C396 B.n223 VSUBS 0.006426f
C397 B.n224 VSUBS 0.005197f
C398 B.n225 VSUBS 0.006426f
C399 B.n226 VSUBS 0.006426f
C400 B.n227 VSUBS 0.004441f
C401 B.n228 VSUBS 0.006426f
C402 B.n229 VSUBS 0.006426f
C403 B.n230 VSUBS 0.006426f
C404 B.n231 VSUBS 0.006426f
C405 B.n232 VSUBS 0.006426f
C406 B.n233 VSUBS 0.006426f
C407 B.n234 VSUBS 0.006426f
C408 B.n235 VSUBS 0.006426f
C409 B.n236 VSUBS 0.006426f
C410 B.n237 VSUBS 0.006426f
C411 B.n238 VSUBS 0.006426f
C412 B.n239 VSUBS 0.006426f
C413 B.n240 VSUBS 0.006426f
C414 B.n241 VSUBS 0.006426f
C415 B.n242 VSUBS 0.006426f
C416 B.n243 VSUBS 0.006426f
C417 B.n244 VSUBS 0.006426f
C418 B.n245 VSUBS 0.006426f
C419 B.n246 VSUBS 0.006426f
C420 B.n247 VSUBS 0.006426f
C421 B.n248 VSUBS 0.006426f
C422 B.n249 VSUBS 0.006426f
C423 B.n250 VSUBS 0.006426f
C424 B.n251 VSUBS 0.006426f
C425 B.n252 VSUBS 0.006426f
C426 B.n253 VSUBS 0.006426f
C427 B.n254 VSUBS 0.006426f
C428 B.n255 VSUBS 0.006426f
C429 B.n256 VSUBS 0.006426f
C430 B.n257 VSUBS 0.006426f
C431 B.n258 VSUBS 0.006426f
C432 B.n259 VSUBS 0.006426f
C433 B.n260 VSUBS 0.006426f
C434 B.n261 VSUBS 0.015586f
C435 B.n262 VSUBS 0.014841f
C436 B.n263 VSUBS 0.014841f
C437 B.n264 VSUBS 0.006426f
C438 B.n265 VSUBS 0.006426f
C439 B.n266 VSUBS 0.006426f
C440 B.n267 VSUBS 0.006426f
C441 B.n268 VSUBS 0.006426f
C442 B.n269 VSUBS 0.006426f
C443 B.n270 VSUBS 0.006426f
C444 B.n271 VSUBS 0.006426f
C445 B.n272 VSUBS 0.006426f
C446 B.n273 VSUBS 0.006426f
C447 B.n274 VSUBS 0.006426f
C448 B.n275 VSUBS 0.006426f
C449 B.n276 VSUBS 0.006426f
C450 B.n277 VSUBS 0.006426f
C451 B.n278 VSUBS 0.006426f
C452 B.n279 VSUBS 0.006426f
C453 B.n280 VSUBS 0.006426f
C454 B.n281 VSUBS 0.006426f
C455 B.n282 VSUBS 0.006426f
C456 B.n283 VSUBS 0.006426f
C457 B.n284 VSUBS 0.006426f
C458 B.n285 VSUBS 0.006426f
C459 B.n286 VSUBS 0.006426f
C460 B.n287 VSUBS 0.006426f
C461 B.n288 VSUBS 0.006426f
C462 B.n289 VSUBS 0.006426f
C463 B.n290 VSUBS 0.006426f
C464 B.n291 VSUBS 0.006426f
C465 B.n292 VSUBS 0.006426f
C466 B.n293 VSUBS 0.006426f
C467 B.n294 VSUBS 0.006426f
C468 B.n295 VSUBS 0.006426f
C469 B.n296 VSUBS 0.006426f
C470 B.n297 VSUBS 0.006426f
C471 B.n298 VSUBS 0.006426f
C472 B.n299 VSUBS 0.006426f
C473 B.n300 VSUBS 0.006426f
C474 B.n301 VSUBS 0.006426f
C475 B.n302 VSUBS 0.006426f
C476 B.n303 VSUBS 0.006426f
C477 B.n304 VSUBS 0.006426f
C478 B.n305 VSUBS 0.006426f
C479 B.n306 VSUBS 0.006426f
C480 B.n307 VSUBS 0.006426f
C481 B.n308 VSUBS 0.006426f
C482 B.n309 VSUBS 0.006426f
C483 B.n310 VSUBS 0.006426f
C484 B.n311 VSUBS 0.006426f
C485 B.n312 VSUBS 0.006426f
C486 B.n313 VSUBS 0.006426f
C487 B.n314 VSUBS 0.006426f
C488 B.n315 VSUBS 0.006426f
C489 B.n316 VSUBS 0.006426f
C490 B.n317 VSUBS 0.006426f
C491 B.n318 VSUBS 0.006426f
C492 B.n319 VSUBS 0.006426f
C493 B.n320 VSUBS 0.006426f
C494 B.n321 VSUBS 0.006426f
C495 B.n322 VSUBS 0.006426f
C496 B.n323 VSUBS 0.006426f
C497 B.n324 VSUBS 0.006426f
C498 B.n325 VSUBS 0.006426f
C499 B.n326 VSUBS 0.006426f
C500 B.n327 VSUBS 0.006426f
C501 B.n328 VSUBS 0.006426f
C502 B.n329 VSUBS 0.006426f
C503 B.n330 VSUBS 0.006426f
C504 B.n331 VSUBS 0.006426f
C505 B.n332 VSUBS 0.006426f
C506 B.n333 VSUBS 0.006426f
C507 B.n334 VSUBS 0.006426f
C508 B.n335 VSUBS 0.006426f
C509 B.n336 VSUBS 0.006426f
C510 B.n337 VSUBS 0.006426f
C511 B.n338 VSUBS 0.006426f
C512 B.n339 VSUBS 0.006426f
C513 B.n340 VSUBS 0.006426f
C514 B.n341 VSUBS 0.006426f
C515 B.n342 VSUBS 0.006426f
C516 B.n343 VSUBS 0.006426f
C517 B.n344 VSUBS 0.006426f
C518 B.n345 VSUBS 0.006426f
C519 B.n346 VSUBS 0.006426f
C520 B.n347 VSUBS 0.006426f
C521 B.n348 VSUBS 0.006426f
C522 B.n349 VSUBS 0.006426f
C523 B.n350 VSUBS 0.006426f
C524 B.n351 VSUBS 0.006426f
C525 B.n352 VSUBS 0.006426f
C526 B.n353 VSUBS 0.006426f
C527 B.n354 VSUBS 0.006426f
C528 B.n355 VSUBS 0.015586f
C529 B.n356 VSUBS 0.014841f
C530 B.n357 VSUBS 0.015586f
C531 B.n358 VSUBS 0.006426f
C532 B.n359 VSUBS 0.006426f
C533 B.n360 VSUBS 0.006426f
C534 B.n361 VSUBS 0.006426f
C535 B.n362 VSUBS 0.006426f
C536 B.n363 VSUBS 0.006426f
C537 B.n364 VSUBS 0.006426f
C538 B.n365 VSUBS 0.006426f
C539 B.n366 VSUBS 0.006426f
C540 B.n367 VSUBS 0.006426f
C541 B.n368 VSUBS 0.006426f
C542 B.n369 VSUBS 0.006426f
C543 B.n370 VSUBS 0.006426f
C544 B.n371 VSUBS 0.006426f
C545 B.n372 VSUBS 0.006426f
C546 B.n373 VSUBS 0.006426f
C547 B.n374 VSUBS 0.006426f
C548 B.n375 VSUBS 0.006426f
C549 B.n376 VSUBS 0.006426f
C550 B.n377 VSUBS 0.006426f
C551 B.n378 VSUBS 0.006426f
C552 B.n379 VSUBS 0.006426f
C553 B.n380 VSUBS 0.006426f
C554 B.n381 VSUBS 0.006426f
C555 B.n382 VSUBS 0.006426f
C556 B.n383 VSUBS 0.006426f
C557 B.n384 VSUBS 0.006426f
C558 B.n385 VSUBS 0.006426f
C559 B.n386 VSUBS 0.006426f
C560 B.n387 VSUBS 0.006426f
C561 B.n388 VSUBS 0.006426f
C562 B.n389 VSUBS 0.006426f
C563 B.n390 VSUBS 0.006426f
C564 B.n391 VSUBS 0.004441f
C565 B.n392 VSUBS 0.006426f
C566 B.n393 VSUBS 0.006426f
C567 B.n394 VSUBS 0.005197f
C568 B.n395 VSUBS 0.006426f
C569 B.n396 VSUBS 0.006426f
C570 B.n397 VSUBS 0.006426f
C571 B.n398 VSUBS 0.006426f
C572 B.n399 VSUBS 0.006426f
C573 B.n400 VSUBS 0.006426f
C574 B.n401 VSUBS 0.006426f
C575 B.n402 VSUBS 0.006426f
C576 B.n403 VSUBS 0.006426f
C577 B.n404 VSUBS 0.006426f
C578 B.n405 VSUBS 0.006426f
C579 B.n406 VSUBS 0.005197f
C580 B.n407 VSUBS 0.014887f
C581 B.n408 VSUBS 0.004441f
C582 B.n409 VSUBS 0.006426f
C583 B.n410 VSUBS 0.006426f
C584 B.n411 VSUBS 0.006426f
C585 B.n412 VSUBS 0.006426f
C586 B.n413 VSUBS 0.006426f
C587 B.n414 VSUBS 0.006426f
C588 B.n415 VSUBS 0.006426f
C589 B.n416 VSUBS 0.006426f
C590 B.n417 VSUBS 0.006426f
C591 B.n418 VSUBS 0.006426f
C592 B.n419 VSUBS 0.006426f
C593 B.n420 VSUBS 0.006426f
C594 B.n421 VSUBS 0.006426f
C595 B.n422 VSUBS 0.006426f
C596 B.n423 VSUBS 0.006426f
C597 B.n424 VSUBS 0.006426f
C598 B.n425 VSUBS 0.006426f
C599 B.n426 VSUBS 0.006426f
C600 B.n427 VSUBS 0.006426f
C601 B.n428 VSUBS 0.006426f
C602 B.n429 VSUBS 0.006426f
C603 B.n430 VSUBS 0.006426f
C604 B.n431 VSUBS 0.006426f
C605 B.n432 VSUBS 0.006426f
C606 B.n433 VSUBS 0.006426f
C607 B.n434 VSUBS 0.006426f
C608 B.n435 VSUBS 0.006426f
C609 B.n436 VSUBS 0.006426f
C610 B.n437 VSUBS 0.006426f
C611 B.n438 VSUBS 0.006426f
C612 B.n439 VSUBS 0.006426f
C613 B.n440 VSUBS 0.006426f
C614 B.n441 VSUBS 0.006426f
C615 B.n442 VSUBS 0.015586f
C616 B.n443 VSUBS 0.015586f
C617 B.n444 VSUBS 0.014841f
C618 B.n445 VSUBS 0.006426f
C619 B.n446 VSUBS 0.006426f
C620 B.n447 VSUBS 0.006426f
C621 B.n448 VSUBS 0.006426f
C622 B.n449 VSUBS 0.006426f
C623 B.n450 VSUBS 0.006426f
C624 B.n451 VSUBS 0.006426f
C625 B.n452 VSUBS 0.006426f
C626 B.n453 VSUBS 0.006426f
C627 B.n454 VSUBS 0.006426f
C628 B.n455 VSUBS 0.006426f
C629 B.n456 VSUBS 0.006426f
C630 B.n457 VSUBS 0.006426f
C631 B.n458 VSUBS 0.006426f
C632 B.n459 VSUBS 0.006426f
C633 B.n460 VSUBS 0.006426f
C634 B.n461 VSUBS 0.006426f
C635 B.n462 VSUBS 0.006426f
C636 B.n463 VSUBS 0.006426f
C637 B.n464 VSUBS 0.006426f
C638 B.n465 VSUBS 0.006426f
C639 B.n466 VSUBS 0.006426f
C640 B.n467 VSUBS 0.006426f
C641 B.n468 VSUBS 0.006426f
C642 B.n469 VSUBS 0.006426f
C643 B.n470 VSUBS 0.006426f
C644 B.n471 VSUBS 0.006426f
C645 B.n472 VSUBS 0.006426f
C646 B.n473 VSUBS 0.006426f
C647 B.n474 VSUBS 0.006426f
C648 B.n475 VSUBS 0.006426f
C649 B.n476 VSUBS 0.006426f
C650 B.n477 VSUBS 0.006426f
C651 B.n478 VSUBS 0.006426f
C652 B.n479 VSUBS 0.006426f
C653 B.n480 VSUBS 0.006426f
C654 B.n481 VSUBS 0.006426f
C655 B.n482 VSUBS 0.006426f
C656 B.n483 VSUBS 0.006426f
C657 B.n484 VSUBS 0.006426f
C658 B.n485 VSUBS 0.006426f
C659 B.n486 VSUBS 0.006426f
C660 B.n487 VSUBS 0.006426f
C661 B.n488 VSUBS 0.006426f
C662 B.n489 VSUBS 0.006426f
C663 B.n490 VSUBS 0.006426f
C664 B.n491 VSUBS 0.01455f
C665 VTAIL.t10 VSUBS 0.137639f
C666 VTAIL.t17 VSUBS 0.137639f
C667 VTAIL.n0 VSUBS 0.799243f
C668 VTAIL.n1 VSUBS 0.728147f
C669 VTAIL.n2 VSUBS 0.031207f
C670 VTAIL.n3 VSUBS 0.029422f
C671 VTAIL.n4 VSUBS 0.01581f
C672 VTAIL.n5 VSUBS 0.037369f
C673 VTAIL.n6 VSUBS 0.01674f
C674 VTAIL.n7 VSUBS 0.029422f
C675 VTAIL.n8 VSUBS 0.01581f
C676 VTAIL.n9 VSUBS 0.037369f
C677 VTAIL.n10 VSUBS 0.01674f
C678 VTAIL.n11 VSUBS 0.129266f
C679 VTAIL.t4 VSUBS 0.080051f
C680 VTAIL.n12 VSUBS 0.028027f
C681 VTAIL.n13 VSUBS 0.02376f
C682 VTAIL.n14 VSUBS 0.01581f
C683 VTAIL.n15 VSUBS 0.664478f
C684 VTAIL.n16 VSUBS 0.029422f
C685 VTAIL.n17 VSUBS 0.01581f
C686 VTAIL.n18 VSUBS 0.01674f
C687 VTAIL.n19 VSUBS 0.037369f
C688 VTAIL.n20 VSUBS 0.037369f
C689 VTAIL.n21 VSUBS 0.01674f
C690 VTAIL.n22 VSUBS 0.01581f
C691 VTAIL.n23 VSUBS 0.029422f
C692 VTAIL.n24 VSUBS 0.029422f
C693 VTAIL.n25 VSUBS 0.01581f
C694 VTAIL.n26 VSUBS 0.01674f
C695 VTAIL.n27 VSUBS 0.037369f
C696 VTAIL.n28 VSUBS 0.086648f
C697 VTAIL.n29 VSUBS 0.01674f
C698 VTAIL.n30 VSUBS 0.01581f
C699 VTAIL.n31 VSUBS 0.064791f
C700 VTAIL.n32 VSUBS 0.043304f
C701 VTAIL.n33 VSUBS 0.227223f
C702 VTAIL.t5 VSUBS 0.137639f
C703 VTAIL.t6 VSUBS 0.137639f
C704 VTAIL.n34 VSUBS 0.799243f
C705 VTAIL.n35 VSUBS 0.757773f
C706 VTAIL.t18 VSUBS 0.137639f
C707 VTAIL.t7 VSUBS 0.137639f
C708 VTAIL.n36 VSUBS 0.799243f
C709 VTAIL.n37 VSUBS 1.74749f
C710 VTAIL.t13 VSUBS 0.137639f
C711 VTAIL.t11 VSUBS 0.137639f
C712 VTAIL.n38 VSUBS 0.799249f
C713 VTAIL.n39 VSUBS 1.74749f
C714 VTAIL.t15 VSUBS 0.137639f
C715 VTAIL.t12 VSUBS 0.137639f
C716 VTAIL.n40 VSUBS 0.799249f
C717 VTAIL.n41 VSUBS 0.757767f
C718 VTAIL.n42 VSUBS 0.031207f
C719 VTAIL.n43 VSUBS 0.029422f
C720 VTAIL.n44 VSUBS 0.01581f
C721 VTAIL.n45 VSUBS 0.037369f
C722 VTAIL.n46 VSUBS 0.01674f
C723 VTAIL.n47 VSUBS 0.029422f
C724 VTAIL.n48 VSUBS 0.01581f
C725 VTAIL.n49 VSUBS 0.037369f
C726 VTAIL.n50 VSUBS 0.01674f
C727 VTAIL.n51 VSUBS 0.129266f
C728 VTAIL.t16 VSUBS 0.080051f
C729 VTAIL.n52 VSUBS 0.028027f
C730 VTAIL.n53 VSUBS 0.02376f
C731 VTAIL.n54 VSUBS 0.01581f
C732 VTAIL.n55 VSUBS 0.664478f
C733 VTAIL.n56 VSUBS 0.029422f
C734 VTAIL.n57 VSUBS 0.01581f
C735 VTAIL.n58 VSUBS 0.01674f
C736 VTAIL.n59 VSUBS 0.037369f
C737 VTAIL.n60 VSUBS 0.037369f
C738 VTAIL.n61 VSUBS 0.01674f
C739 VTAIL.n62 VSUBS 0.01581f
C740 VTAIL.n63 VSUBS 0.029422f
C741 VTAIL.n64 VSUBS 0.029422f
C742 VTAIL.n65 VSUBS 0.01581f
C743 VTAIL.n66 VSUBS 0.01674f
C744 VTAIL.n67 VSUBS 0.037369f
C745 VTAIL.n68 VSUBS 0.086648f
C746 VTAIL.n69 VSUBS 0.01674f
C747 VTAIL.n70 VSUBS 0.01581f
C748 VTAIL.n71 VSUBS 0.064791f
C749 VTAIL.n72 VSUBS 0.043304f
C750 VTAIL.n73 VSUBS 0.227223f
C751 VTAIL.t3 VSUBS 0.137639f
C752 VTAIL.t19 VSUBS 0.137639f
C753 VTAIL.n74 VSUBS 0.799249f
C754 VTAIL.n75 VSUBS 0.749186f
C755 VTAIL.t1 VSUBS 0.137639f
C756 VTAIL.t0 VSUBS 0.137639f
C757 VTAIL.n76 VSUBS 0.799249f
C758 VTAIL.n77 VSUBS 0.757767f
C759 VTAIL.n78 VSUBS 0.031207f
C760 VTAIL.n79 VSUBS 0.029422f
C761 VTAIL.n80 VSUBS 0.01581f
C762 VTAIL.n81 VSUBS 0.037369f
C763 VTAIL.n82 VSUBS 0.01674f
C764 VTAIL.n83 VSUBS 0.029422f
C765 VTAIL.n84 VSUBS 0.01581f
C766 VTAIL.n85 VSUBS 0.037369f
C767 VTAIL.n86 VSUBS 0.01674f
C768 VTAIL.n87 VSUBS 0.129266f
C769 VTAIL.t2 VSUBS 0.080051f
C770 VTAIL.n88 VSUBS 0.028027f
C771 VTAIL.n89 VSUBS 0.02376f
C772 VTAIL.n90 VSUBS 0.01581f
C773 VTAIL.n91 VSUBS 0.664478f
C774 VTAIL.n92 VSUBS 0.029422f
C775 VTAIL.n93 VSUBS 0.01581f
C776 VTAIL.n94 VSUBS 0.01674f
C777 VTAIL.n95 VSUBS 0.037369f
C778 VTAIL.n96 VSUBS 0.037369f
C779 VTAIL.n97 VSUBS 0.01674f
C780 VTAIL.n98 VSUBS 0.01581f
C781 VTAIL.n99 VSUBS 0.029422f
C782 VTAIL.n100 VSUBS 0.029422f
C783 VTAIL.n101 VSUBS 0.01581f
C784 VTAIL.n102 VSUBS 0.01674f
C785 VTAIL.n103 VSUBS 0.037369f
C786 VTAIL.n104 VSUBS 0.086648f
C787 VTAIL.n105 VSUBS 0.01674f
C788 VTAIL.n106 VSUBS 0.01581f
C789 VTAIL.n107 VSUBS 0.064791f
C790 VTAIL.n108 VSUBS 0.043304f
C791 VTAIL.n109 VSUBS 1.11928f
C792 VTAIL.n110 VSUBS 0.031207f
C793 VTAIL.n111 VSUBS 0.029422f
C794 VTAIL.n112 VSUBS 0.01581f
C795 VTAIL.n113 VSUBS 0.037369f
C796 VTAIL.n114 VSUBS 0.01674f
C797 VTAIL.n115 VSUBS 0.029422f
C798 VTAIL.n116 VSUBS 0.01581f
C799 VTAIL.n117 VSUBS 0.037369f
C800 VTAIL.n118 VSUBS 0.01674f
C801 VTAIL.n119 VSUBS 0.129266f
C802 VTAIL.t8 VSUBS 0.080051f
C803 VTAIL.n120 VSUBS 0.028027f
C804 VTAIL.n121 VSUBS 0.02376f
C805 VTAIL.n122 VSUBS 0.01581f
C806 VTAIL.n123 VSUBS 0.664478f
C807 VTAIL.n124 VSUBS 0.029422f
C808 VTAIL.n125 VSUBS 0.01581f
C809 VTAIL.n126 VSUBS 0.01674f
C810 VTAIL.n127 VSUBS 0.037369f
C811 VTAIL.n128 VSUBS 0.037369f
C812 VTAIL.n129 VSUBS 0.01674f
C813 VTAIL.n130 VSUBS 0.01581f
C814 VTAIL.n131 VSUBS 0.029422f
C815 VTAIL.n132 VSUBS 0.029422f
C816 VTAIL.n133 VSUBS 0.01581f
C817 VTAIL.n134 VSUBS 0.01674f
C818 VTAIL.n135 VSUBS 0.037369f
C819 VTAIL.n136 VSUBS 0.086648f
C820 VTAIL.n137 VSUBS 0.01674f
C821 VTAIL.n138 VSUBS 0.01581f
C822 VTAIL.n139 VSUBS 0.064791f
C823 VTAIL.n140 VSUBS 0.043304f
C824 VTAIL.n141 VSUBS 1.11928f
C825 VTAIL.t9 VSUBS 0.137639f
C826 VTAIL.t14 VSUBS 0.137639f
C827 VTAIL.n142 VSUBS 0.799243f
C828 VTAIL.n143 VSUBS 0.672573f
C829 VDD2.n0 VSUBS 0.024946f
C830 VDD2.n1 VSUBS 0.023519f
C831 VDD2.n2 VSUBS 0.012638f
C832 VDD2.n3 VSUBS 0.029872f
C833 VDD2.n4 VSUBS 0.013381f
C834 VDD2.n5 VSUBS 0.023519f
C835 VDD2.n6 VSUBS 0.012638f
C836 VDD2.n7 VSUBS 0.029872f
C837 VDD2.n8 VSUBS 0.013381f
C838 VDD2.n9 VSUBS 0.103331f
C839 VDD2.t8 VSUBS 0.063991f
C840 VDD2.n10 VSUBS 0.022404f
C841 VDD2.n11 VSUBS 0.018993f
C842 VDD2.n12 VSUBS 0.012638f
C843 VDD2.n13 VSUBS 0.531165f
C844 VDD2.n14 VSUBS 0.023519f
C845 VDD2.n15 VSUBS 0.012638f
C846 VDD2.n16 VSUBS 0.013381f
C847 VDD2.n17 VSUBS 0.029872f
C848 VDD2.n18 VSUBS 0.029872f
C849 VDD2.n19 VSUBS 0.013381f
C850 VDD2.n20 VSUBS 0.012638f
C851 VDD2.n21 VSUBS 0.023519f
C852 VDD2.n22 VSUBS 0.023519f
C853 VDD2.n23 VSUBS 0.012638f
C854 VDD2.n24 VSUBS 0.013381f
C855 VDD2.n25 VSUBS 0.029872f
C856 VDD2.n26 VSUBS 0.069264f
C857 VDD2.n27 VSUBS 0.013381f
C858 VDD2.n28 VSUBS 0.012638f
C859 VDD2.n29 VSUBS 0.051792f
C860 VDD2.n30 VSUBS 0.053856f
C861 VDD2.t9 VSUBS 0.110025f
C862 VDD2.t0 VSUBS 0.110025f
C863 VDD2.n31 VSUBS 0.724063f
C864 VDD2.n32 VSUBS 0.61284f
C865 VDD2.t6 VSUBS 0.110025f
C866 VDD2.t2 VSUBS 0.110025f
C867 VDD2.n33 VSUBS 0.728672f
C868 VDD2.n34 VSUBS 1.77325f
C869 VDD2.n35 VSUBS 0.024946f
C870 VDD2.n36 VSUBS 0.023519f
C871 VDD2.n37 VSUBS 0.012638f
C872 VDD2.n38 VSUBS 0.029872f
C873 VDD2.n39 VSUBS 0.013381f
C874 VDD2.n40 VSUBS 0.023519f
C875 VDD2.n41 VSUBS 0.012638f
C876 VDD2.n42 VSUBS 0.029872f
C877 VDD2.n43 VSUBS 0.013381f
C878 VDD2.n44 VSUBS 0.103331f
C879 VDD2.t7 VSUBS 0.063991f
C880 VDD2.n45 VSUBS 0.022404f
C881 VDD2.n46 VSUBS 0.018993f
C882 VDD2.n47 VSUBS 0.012638f
C883 VDD2.n48 VSUBS 0.531165f
C884 VDD2.n49 VSUBS 0.023519f
C885 VDD2.n50 VSUBS 0.012638f
C886 VDD2.n51 VSUBS 0.013381f
C887 VDD2.n52 VSUBS 0.029872f
C888 VDD2.n53 VSUBS 0.029872f
C889 VDD2.n54 VSUBS 0.013381f
C890 VDD2.n55 VSUBS 0.012638f
C891 VDD2.n56 VSUBS 0.023519f
C892 VDD2.n57 VSUBS 0.023519f
C893 VDD2.n58 VSUBS 0.012638f
C894 VDD2.n59 VSUBS 0.013381f
C895 VDD2.n60 VSUBS 0.029872f
C896 VDD2.n61 VSUBS 0.069264f
C897 VDD2.n62 VSUBS 0.013381f
C898 VDD2.n63 VSUBS 0.012638f
C899 VDD2.n64 VSUBS 0.051792f
C900 VDD2.n65 VSUBS 0.050877f
C901 VDD2.n66 VSUBS 1.67039f
C902 VDD2.t4 VSUBS 0.110025f
C903 VDD2.t3 VSUBS 0.110025f
C904 VDD2.n67 VSUBS 0.724067f
C905 VDD2.n68 VSUBS 0.493249f
C906 VDD2.t5 VSUBS 0.110025f
C907 VDD2.t1 VSUBS 0.110025f
C908 VDD2.n69 VSUBS 0.728648f
C909 VN.n0 VSUBS 0.070616f
C910 VN.t3 VSUBS 0.803695f
C911 VN.n1 VSUBS 0.049896f
C912 VN.n2 VSUBS 0.052921f
C913 VN.t8 VSUBS 0.803695f
C914 VN.n3 VSUBS 0.061842f
C915 VN.t7 VSUBS 0.909847f
C916 VN.t0 VSUBS 0.803695f
C917 VN.n4 VSUBS 0.366668f
C918 VN.n5 VSUBS 0.408037f
C919 VN.n6 VSUBS 0.216208f
C920 VN.n7 VSUBS 0.052921f
C921 VN.n8 VSUBS 0.049896f
C922 VN.n9 VSUBS 0.072428f
C923 VN.n10 VSUBS 0.33233f
C924 VN.n11 VSUBS 0.072428f
C925 VN.n12 VSUBS 0.052921f
C926 VN.n13 VSUBS 0.052921f
C927 VN.n14 VSUBS 0.052921f
C928 VN.n15 VSUBS 0.061842f
C929 VN.n16 VSUBS 0.33233f
C930 VN.n17 VSUBS 0.061906f
C931 VN.t9 VSUBS 0.881859f
C932 VN.n18 VSUBS 0.407434f
C933 VN.n19 VSUBS 0.049562f
C934 VN.n20 VSUBS 0.070616f
C935 VN.t6 VSUBS 0.803695f
C936 VN.n21 VSUBS 0.049896f
C937 VN.n22 VSUBS 0.052921f
C938 VN.t2 VSUBS 0.803695f
C939 VN.n23 VSUBS 0.061842f
C940 VN.t1 VSUBS 0.909847f
C941 VN.t5 VSUBS 0.803695f
C942 VN.n24 VSUBS 0.366668f
C943 VN.n25 VSUBS 0.408037f
C944 VN.n26 VSUBS 0.216208f
C945 VN.n27 VSUBS 0.052921f
C946 VN.n28 VSUBS 0.049896f
C947 VN.n29 VSUBS 0.072428f
C948 VN.n30 VSUBS 0.33233f
C949 VN.n31 VSUBS 0.072428f
C950 VN.n32 VSUBS 0.052921f
C951 VN.n33 VSUBS 0.052921f
C952 VN.n34 VSUBS 0.052921f
C953 VN.n35 VSUBS 0.061842f
C954 VN.n36 VSUBS 0.33233f
C955 VN.n37 VSUBS 0.061906f
C956 VN.t4 VSUBS 0.881859f
C957 VN.n38 VSUBS 0.407434f
C958 VN.n39 VSUBS 2.03753f
.ends

