* NGSPICE file created from diff_pair_sample_0657.ext - technology: sky130A

.subckt diff_pair_sample_0657 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=2.2968 ps=14.25 w=13.92 l=3.1
X1 VDD2.t9 VN.t0 VTAIL.t2 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=2.2968 ps=14.25 w=13.92 l=3.1
X2 VTAIL.t6 VN.t1 VDD2.t8 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X3 B.t11 B.t9 B.t10 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=0 ps=0 w=13.92 l=3.1
X4 VTAIL.t12 VP.t1 VDD1.t8 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X5 VTAIL.t18 VP.t2 VDD1.t7 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X6 VDD1.t6 VP.t3 VTAIL.t10 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=5.4288 ps=28.62 w=13.92 l=3.1
X7 B.t8 B.t6 B.t7 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=0 ps=0 w=13.92 l=3.1
X8 VTAIL.t17 VP.t4 VDD1.t5 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X9 VDD2.t7 VN.t2 VTAIL.t5 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=5.4288 ps=28.62 w=13.92 l=3.1
X10 VDD1.t4 VP.t5 VTAIL.t19 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X11 VDD2.t6 VN.t3 VTAIL.t9 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X12 B.t5 B.t3 B.t4 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=0 ps=0 w=13.92 l=3.1
X13 VDD2.t5 VN.t4 VTAIL.t4 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=5.4288 ps=28.62 w=13.92 l=3.1
X14 B.t2 B.t0 B.t1 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=0 ps=0 w=13.92 l=3.1
X15 VDD1.t3 VP.t6 VTAIL.t13 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X16 VTAIL.t7 VN.t5 VDD2.t4 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X17 VDD2.t3 VN.t6 VTAIL.t8 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X18 VDD1.t2 VP.t7 VTAIL.t14 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=5.4288 ps=28.62 w=13.92 l=3.1
X19 VTAIL.t3 VN.t7 VDD2.t2 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X20 VTAIL.t15 VP.t8 VDD1.t1 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
X21 VDD1.t0 VP.t9 VTAIL.t16 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=2.2968 ps=14.25 w=13.92 l=3.1
X22 VDD2.t1 VN.t8 VTAIL.t0 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=5.4288 pd=28.62 as=2.2968 ps=14.25 w=13.92 l=3.1
X23 VTAIL.t1 VN.t9 VDD2.t0 w_n5086_n3752# sky130_fd_pr__pfet_01v8 ad=2.2968 pd=14.25 as=2.2968 ps=14.25 w=13.92 l=3.1
R0 VP.n29 VP.n28 161.3
R1 VP.n30 VP.n25 161.3
R2 VP.n32 VP.n31 161.3
R3 VP.n33 VP.n24 161.3
R4 VP.n35 VP.n34 161.3
R5 VP.n36 VP.n23 161.3
R6 VP.n38 VP.n37 161.3
R7 VP.n39 VP.n22 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n42 VP.n21 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n45 VP.n20 161.3
R12 VP.n47 VP.n46 161.3
R13 VP.n49 VP.n48 161.3
R14 VP.n50 VP.n18 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n17 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n16 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n94 VP.n93 161.3
R27 VP.n92 VP.n91 161.3
R28 VP.n90 VP.n5 161.3
R29 VP.n89 VP.n88 161.3
R30 VP.n87 VP.n6 161.3
R31 VP.n86 VP.n85 161.3
R32 VP.n84 VP.n7 161.3
R33 VP.n83 VP.n82 161.3
R34 VP.n81 VP.n8 161.3
R35 VP.n80 VP.n79 161.3
R36 VP.n78 VP.n9 161.3
R37 VP.n77 VP.n76 161.3
R38 VP.n75 VP.n10 161.3
R39 VP.n74 VP.n73 161.3
R40 VP.n71 VP.n11 161.3
R41 VP.n70 VP.n69 161.3
R42 VP.n68 VP.n12 161.3
R43 VP.n67 VP.n66 161.3
R44 VP.n65 VP.n13 161.3
R45 VP.n64 VP.n63 161.3
R46 VP.n62 VP.n14 161.3
R47 VP.n26 VP.t0 141.593
R48 VP.n83 VP.t5 108.218
R49 VP.n60 VP.t9 108.218
R50 VP.n72 VP.t2 108.218
R51 VP.n4 VP.t8 108.218
R52 VP.n0 VP.t7 108.218
R53 VP.n38 VP.t6 108.218
R54 VP.n15 VP.t3 108.218
R55 VP.n19 VP.t1 108.218
R56 VP.n27 VP.t4 108.218
R57 VP.n61 VP.n60 72.5394
R58 VP.n104 VP.n0 72.5394
R59 VP.n59 VP.n15 72.5394
R60 VP.n61 VP.n59 57.3973
R61 VP.n78 VP.n77 56.5617
R62 VP.n44 VP.n21 56.5617
R63 VP.n89 VP.n6 56.5617
R64 VP.n33 VP.n32 56.5617
R65 VP.n66 VP.n65 54.6242
R66 VP.n100 VP.n2 54.6242
R67 VP.n55 VP.n17 54.6242
R68 VP.n27 VP.n26 52.9403
R69 VP.n66 VP.n12 26.5299
R70 VP.n96 VP.n2 26.5299
R71 VP.n51 VP.n17 26.5299
R72 VP.n64 VP.n14 24.5923
R73 VP.n65 VP.n64 24.5923
R74 VP.n70 VP.n12 24.5923
R75 VP.n71 VP.n70 24.5923
R76 VP.n73 VP.n10 24.5923
R77 VP.n77 VP.n10 24.5923
R78 VP.n79 VP.n78 24.5923
R79 VP.n79 VP.n8 24.5923
R80 VP.n83 VP.n8 24.5923
R81 VP.n84 VP.n83 24.5923
R82 VP.n85 VP.n84 24.5923
R83 VP.n85 VP.n6 24.5923
R84 VP.n90 VP.n89 24.5923
R85 VP.n91 VP.n90 24.5923
R86 VP.n95 VP.n94 24.5923
R87 VP.n96 VP.n95 24.5923
R88 VP.n101 VP.n100 24.5923
R89 VP.n102 VP.n101 24.5923
R90 VP.n56 VP.n55 24.5923
R91 VP.n57 VP.n56 24.5923
R92 VP.n45 VP.n44 24.5923
R93 VP.n46 VP.n45 24.5923
R94 VP.n50 VP.n49 24.5923
R95 VP.n51 VP.n50 24.5923
R96 VP.n34 VP.n33 24.5923
R97 VP.n34 VP.n23 24.5923
R98 VP.n38 VP.n23 24.5923
R99 VP.n39 VP.n38 24.5923
R100 VP.n40 VP.n39 24.5923
R101 VP.n40 VP.n21 24.5923
R102 VP.n28 VP.n25 24.5923
R103 VP.n32 VP.n25 24.5923
R104 VP.n73 VP.n72 21.1495
R105 VP.n91 VP.n4 21.1495
R106 VP.n46 VP.n19 21.1495
R107 VP.n28 VP.n27 21.1495
R108 VP.n60 VP.n14 17.7066
R109 VP.n102 VP.n0 17.7066
R110 VP.n57 VP.n15 17.7066
R111 VP.n29 VP.n26 4.01097
R112 VP.n72 VP.n71 3.44336
R113 VP.n94 VP.n4 3.44336
R114 VP.n49 VP.n19 3.44336
R115 VP.n59 VP.n58 0.354861
R116 VP.n62 VP.n61 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n30 VP.n29 0.189894
R120 VP.n31 VP.n30 0.189894
R121 VP.n31 VP.n24 0.189894
R122 VP.n35 VP.n24 0.189894
R123 VP.n36 VP.n35 0.189894
R124 VP.n37 VP.n36 0.189894
R125 VP.n37 VP.n22 0.189894
R126 VP.n41 VP.n22 0.189894
R127 VP.n42 VP.n41 0.189894
R128 VP.n43 VP.n42 0.189894
R129 VP.n43 VP.n20 0.189894
R130 VP.n47 VP.n20 0.189894
R131 VP.n48 VP.n47 0.189894
R132 VP.n48 VP.n18 0.189894
R133 VP.n52 VP.n18 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n16 0.189894
R137 VP.n58 VP.n16 0.189894
R138 VP.n63 VP.n62 0.189894
R139 VP.n63 VP.n13 0.189894
R140 VP.n67 VP.n13 0.189894
R141 VP.n68 VP.n67 0.189894
R142 VP.n69 VP.n68 0.189894
R143 VP.n69 VP.n11 0.189894
R144 VP.n74 VP.n11 0.189894
R145 VP.n75 VP.n74 0.189894
R146 VP.n76 VP.n75 0.189894
R147 VP.n76 VP.n9 0.189894
R148 VP.n80 VP.n9 0.189894
R149 VP.n81 VP.n80 0.189894
R150 VP.n82 VP.n81 0.189894
R151 VP.n82 VP.n7 0.189894
R152 VP.n86 VP.n7 0.189894
R153 VP.n87 VP.n86 0.189894
R154 VP.n88 VP.n87 0.189894
R155 VP.n88 VP.n5 0.189894
R156 VP.n92 VP.n5 0.189894
R157 VP.n93 VP.n92 0.189894
R158 VP.n93 VP.n3 0.189894
R159 VP.n97 VP.n3 0.189894
R160 VP.n98 VP.n97 0.189894
R161 VP.n99 VP.n98 0.189894
R162 VP.n99 VP.n1 0.189894
R163 VP.n103 VP.n1 0.189894
R164 VTAIL.n16 VTAIL.t10 57.6035
R165 VTAIL.n11 VTAIL.t5 57.6035
R166 VTAIL.n17 VTAIL.t4 57.6033
R167 VTAIL.n2 VTAIL.t14 57.6033
R168 VTAIL.n15 VTAIL.n14 55.2684
R169 VTAIL.n13 VTAIL.n12 55.2684
R170 VTAIL.n10 VTAIL.n9 55.2684
R171 VTAIL.n8 VTAIL.n7 55.2684
R172 VTAIL.n19 VTAIL.n18 55.2683
R173 VTAIL.n1 VTAIL.n0 55.2683
R174 VTAIL.n4 VTAIL.n3 55.2683
R175 VTAIL.n6 VTAIL.n5 55.2683
R176 VTAIL.n8 VTAIL.n6 30.2807
R177 VTAIL.n17 VTAIL.n16 27.3238
R178 VTAIL.n10 VTAIL.n8 2.9574
R179 VTAIL.n11 VTAIL.n10 2.9574
R180 VTAIL.n15 VTAIL.n13 2.9574
R181 VTAIL.n16 VTAIL.n15 2.9574
R182 VTAIL.n6 VTAIL.n4 2.9574
R183 VTAIL.n4 VTAIL.n2 2.9574
R184 VTAIL.n19 VTAIL.n17 2.9574
R185 VTAIL.n18 VTAIL.t8 2.33563
R186 VTAIL.n18 VTAIL.t3 2.33563
R187 VTAIL.n0 VTAIL.t2 2.33563
R188 VTAIL.n0 VTAIL.t6 2.33563
R189 VTAIL.n3 VTAIL.t19 2.33563
R190 VTAIL.n3 VTAIL.t15 2.33563
R191 VTAIL.n5 VTAIL.t16 2.33563
R192 VTAIL.n5 VTAIL.t18 2.33563
R193 VTAIL.n14 VTAIL.t13 2.33563
R194 VTAIL.n14 VTAIL.t12 2.33563
R195 VTAIL.n12 VTAIL.t11 2.33563
R196 VTAIL.n12 VTAIL.t17 2.33563
R197 VTAIL.n9 VTAIL.t9 2.33563
R198 VTAIL.n9 VTAIL.t1 2.33563
R199 VTAIL.n7 VTAIL.t0 2.33563
R200 VTAIL.n7 VTAIL.t7 2.33563
R201 VTAIL VTAIL.n1 2.27636
R202 VTAIL.n13 VTAIL.n11 1.94878
R203 VTAIL.n2 VTAIL.n1 1.94878
R204 VTAIL VTAIL.n19 0.681535
R205 VDD1.n1 VDD1.t9 77.2391
R206 VDD1.n3 VDD1.t0 77.239
R207 VDD1.n5 VDD1.n4 74.1094
R208 VDD1.n7 VDD1.n6 71.9472
R209 VDD1.n1 VDD1.n0 71.9472
R210 VDD1.n3 VDD1.n2 71.9471
R211 VDD1.n7 VDD1.n5 51.822
R212 VDD1.n6 VDD1.t8 2.33563
R213 VDD1.n6 VDD1.t6 2.33563
R214 VDD1.n0 VDD1.t5 2.33563
R215 VDD1.n0 VDD1.t3 2.33563
R216 VDD1.n4 VDD1.t1 2.33563
R217 VDD1.n4 VDD1.t2 2.33563
R218 VDD1.n2 VDD1.t7 2.33563
R219 VDD1.n2 VDD1.t4 2.33563
R220 VDD1 VDD1.n7 2.15998
R221 VDD1 VDD1.n1 0.797914
R222 VDD1.n5 VDD1.n3 0.684378
R223 VN.n88 VN.n87 161.3
R224 VN.n86 VN.n46 161.3
R225 VN.n85 VN.n84 161.3
R226 VN.n83 VN.n47 161.3
R227 VN.n82 VN.n81 161.3
R228 VN.n80 VN.n48 161.3
R229 VN.n79 VN.n78 161.3
R230 VN.n77 VN.n76 161.3
R231 VN.n75 VN.n50 161.3
R232 VN.n74 VN.n73 161.3
R233 VN.n72 VN.n51 161.3
R234 VN.n71 VN.n70 161.3
R235 VN.n69 VN.n52 161.3
R236 VN.n68 VN.n67 161.3
R237 VN.n66 VN.n53 161.3
R238 VN.n65 VN.n64 161.3
R239 VN.n63 VN.n54 161.3
R240 VN.n62 VN.n61 161.3
R241 VN.n60 VN.n55 161.3
R242 VN.n59 VN.n58 161.3
R243 VN.n43 VN.n42 161.3
R244 VN.n41 VN.n1 161.3
R245 VN.n40 VN.n39 161.3
R246 VN.n38 VN.n2 161.3
R247 VN.n37 VN.n36 161.3
R248 VN.n35 VN.n3 161.3
R249 VN.n34 VN.n33 161.3
R250 VN.n32 VN.n31 161.3
R251 VN.n30 VN.n5 161.3
R252 VN.n29 VN.n28 161.3
R253 VN.n27 VN.n6 161.3
R254 VN.n26 VN.n25 161.3
R255 VN.n24 VN.n7 161.3
R256 VN.n23 VN.n22 161.3
R257 VN.n21 VN.n8 161.3
R258 VN.n20 VN.n19 161.3
R259 VN.n18 VN.n9 161.3
R260 VN.n17 VN.n16 161.3
R261 VN.n15 VN.n10 161.3
R262 VN.n14 VN.n13 161.3
R263 VN.n56 VN.t2 141.593
R264 VN.n11 VN.t0 141.593
R265 VN.n23 VN.t6 108.218
R266 VN.n12 VN.t1 108.218
R267 VN.n4 VN.t7 108.218
R268 VN.n0 VN.t4 108.218
R269 VN.n68 VN.t3 108.218
R270 VN.n57 VN.t9 108.218
R271 VN.n49 VN.t5 108.218
R272 VN.n45 VN.t8 108.218
R273 VN.n44 VN.n0 72.5394
R274 VN.n89 VN.n45 72.5394
R275 VN VN.n89 57.5625
R276 VN.n18 VN.n17 56.5617
R277 VN.n63 VN.n62 56.5617
R278 VN.n29 VN.n6 56.5617
R279 VN.n74 VN.n51 56.5617
R280 VN.n40 VN.n2 54.6242
R281 VN.n85 VN.n47 54.6242
R282 VN.n12 VN.n11 52.9403
R283 VN.n57 VN.n56 52.9403
R284 VN.n36 VN.n2 26.5299
R285 VN.n81 VN.n47 26.5299
R286 VN.n13 VN.n10 24.5923
R287 VN.n17 VN.n10 24.5923
R288 VN.n19 VN.n18 24.5923
R289 VN.n19 VN.n8 24.5923
R290 VN.n23 VN.n8 24.5923
R291 VN.n24 VN.n23 24.5923
R292 VN.n25 VN.n24 24.5923
R293 VN.n25 VN.n6 24.5923
R294 VN.n30 VN.n29 24.5923
R295 VN.n31 VN.n30 24.5923
R296 VN.n35 VN.n34 24.5923
R297 VN.n36 VN.n35 24.5923
R298 VN.n41 VN.n40 24.5923
R299 VN.n42 VN.n41 24.5923
R300 VN.n62 VN.n55 24.5923
R301 VN.n58 VN.n55 24.5923
R302 VN.n70 VN.n51 24.5923
R303 VN.n70 VN.n69 24.5923
R304 VN.n69 VN.n68 24.5923
R305 VN.n68 VN.n53 24.5923
R306 VN.n64 VN.n53 24.5923
R307 VN.n64 VN.n63 24.5923
R308 VN.n81 VN.n80 24.5923
R309 VN.n80 VN.n79 24.5923
R310 VN.n76 VN.n75 24.5923
R311 VN.n75 VN.n74 24.5923
R312 VN.n87 VN.n86 24.5923
R313 VN.n86 VN.n85 24.5923
R314 VN.n13 VN.n12 21.1495
R315 VN.n31 VN.n4 21.1495
R316 VN.n58 VN.n57 21.1495
R317 VN.n76 VN.n49 21.1495
R318 VN.n42 VN.n0 17.7066
R319 VN.n87 VN.n45 17.7066
R320 VN.n59 VN.n56 4.011
R321 VN.n14 VN.n11 4.011
R322 VN.n34 VN.n4 3.44336
R323 VN.n79 VN.n49 3.44336
R324 VN.n89 VN.n88 0.354861
R325 VN.n44 VN.n43 0.354861
R326 VN VN.n44 0.267071
R327 VN.n88 VN.n46 0.189894
R328 VN.n84 VN.n46 0.189894
R329 VN.n84 VN.n83 0.189894
R330 VN.n83 VN.n82 0.189894
R331 VN.n82 VN.n48 0.189894
R332 VN.n78 VN.n48 0.189894
R333 VN.n78 VN.n77 0.189894
R334 VN.n77 VN.n50 0.189894
R335 VN.n73 VN.n50 0.189894
R336 VN.n73 VN.n72 0.189894
R337 VN.n72 VN.n71 0.189894
R338 VN.n71 VN.n52 0.189894
R339 VN.n67 VN.n52 0.189894
R340 VN.n67 VN.n66 0.189894
R341 VN.n66 VN.n65 0.189894
R342 VN.n65 VN.n54 0.189894
R343 VN.n61 VN.n54 0.189894
R344 VN.n61 VN.n60 0.189894
R345 VN.n60 VN.n59 0.189894
R346 VN.n15 VN.n14 0.189894
R347 VN.n16 VN.n15 0.189894
R348 VN.n16 VN.n9 0.189894
R349 VN.n20 VN.n9 0.189894
R350 VN.n21 VN.n20 0.189894
R351 VN.n22 VN.n21 0.189894
R352 VN.n22 VN.n7 0.189894
R353 VN.n26 VN.n7 0.189894
R354 VN.n27 VN.n26 0.189894
R355 VN.n28 VN.n27 0.189894
R356 VN.n28 VN.n5 0.189894
R357 VN.n32 VN.n5 0.189894
R358 VN.n33 VN.n32 0.189894
R359 VN.n33 VN.n3 0.189894
R360 VN.n37 VN.n3 0.189894
R361 VN.n38 VN.n37 0.189894
R362 VN.n39 VN.n38 0.189894
R363 VN.n39 VN.n1 0.189894
R364 VN.n43 VN.n1 0.189894
R365 VDD2.n1 VDD2.t9 77.239
R366 VDD2.n4 VDD2.t1 74.2823
R367 VDD2.n3 VDD2.n2 74.1094
R368 VDD2 VDD2.n7 74.1066
R369 VDD2.n6 VDD2.n5 71.9472
R370 VDD2.n1 VDD2.n0 71.9471
R371 VDD2.n4 VDD2.n3 49.7606
R372 VDD2.n6 VDD2.n4 2.9574
R373 VDD2.n7 VDD2.t0 2.33563
R374 VDD2.n7 VDD2.t7 2.33563
R375 VDD2.n5 VDD2.t4 2.33563
R376 VDD2.n5 VDD2.t6 2.33563
R377 VDD2.n2 VDD2.t2 2.33563
R378 VDD2.n2 VDD2.t5 2.33563
R379 VDD2.n0 VDD2.t8 2.33563
R380 VDD2.n0 VDD2.t3 2.33563
R381 VDD2 VDD2.n6 0.797914
R382 VDD2.n3 VDD2.n1 0.684378
R383 B.n509 B.n162 585
R384 B.n508 B.n507 585
R385 B.n506 B.n163 585
R386 B.n505 B.n504 585
R387 B.n503 B.n164 585
R388 B.n502 B.n501 585
R389 B.n500 B.n165 585
R390 B.n499 B.n498 585
R391 B.n497 B.n166 585
R392 B.n496 B.n495 585
R393 B.n494 B.n167 585
R394 B.n493 B.n492 585
R395 B.n491 B.n168 585
R396 B.n490 B.n489 585
R397 B.n488 B.n169 585
R398 B.n487 B.n486 585
R399 B.n485 B.n170 585
R400 B.n484 B.n483 585
R401 B.n482 B.n171 585
R402 B.n481 B.n480 585
R403 B.n479 B.n172 585
R404 B.n478 B.n477 585
R405 B.n476 B.n173 585
R406 B.n475 B.n474 585
R407 B.n473 B.n174 585
R408 B.n472 B.n471 585
R409 B.n470 B.n175 585
R410 B.n469 B.n468 585
R411 B.n467 B.n176 585
R412 B.n466 B.n465 585
R413 B.n464 B.n177 585
R414 B.n463 B.n462 585
R415 B.n461 B.n178 585
R416 B.n460 B.n459 585
R417 B.n458 B.n179 585
R418 B.n457 B.n456 585
R419 B.n455 B.n180 585
R420 B.n454 B.n453 585
R421 B.n452 B.n181 585
R422 B.n451 B.n450 585
R423 B.n449 B.n182 585
R424 B.n448 B.n447 585
R425 B.n446 B.n183 585
R426 B.n445 B.n444 585
R427 B.n443 B.n184 585
R428 B.n442 B.n441 585
R429 B.n440 B.n185 585
R430 B.n439 B.n438 585
R431 B.n434 B.n186 585
R432 B.n433 B.n432 585
R433 B.n431 B.n187 585
R434 B.n430 B.n429 585
R435 B.n428 B.n188 585
R436 B.n427 B.n426 585
R437 B.n425 B.n189 585
R438 B.n424 B.n423 585
R439 B.n422 B.n190 585
R440 B.n420 B.n419 585
R441 B.n418 B.n193 585
R442 B.n417 B.n416 585
R443 B.n415 B.n194 585
R444 B.n414 B.n413 585
R445 B.n412 B.n195 585
R446 B.n411 B.n410 585
R447 B.n409 B.n196 585
R448 B.n408 B.n407 585
R449 B.n406 B.n197 585
R450 B.n405 B.n404 585
R451 B.n403 B.n198 585
R452 B.n402 B.n401 585
R453 B.n400 B.n199 585
R454 B.n399 B.n398 585
R455 B.n397 B.n200 585
R456 B.n396 B.n395 585
R457 B.n394 B.n201 585
R458 B.n393 B.n392 585
R459 B.n391 B.n202 585
R460 B.n390 B.n389 585
R461 B.n388 B.n203 585
R462 B.n387 B.n386 585
R463 B.n385 B.n204 585
R464 B.n384 B.n383 585
R465 B.n382 B.n205 585
R466 B.n381 B.n380 585
R467 B.n379 B.n206 585
R468 B.n378 B.n377 585
R469 B.n376 B.n207 585
R470 B.n375 B.n374 585
R471 B.n373 B.n208 585
R472 B.n372 B.n371 585
R473 B.n370 B.n209 585
R474 B.n369 B.n368 585
R475 B.n367 B.n210 585
R476 B.n366 B.n365 585
R477 B.n364 B.n211 585
R478 B.n363 B.n362 585
R479 B.n361 B.n212 585
R480 B.n360 B.n359 585
R481 B.n358 B.n213 585
R482 B.n357 B.n356 585
R483 B.n355 B.n214 585
R484 B.n354 B.n353 585
R485 B.n352 B.n215 585
R486 B.n351 B.n350 585
R487 B.n511 B.n510 585
R488 B.n512 B.n161 585
R489 B.n514 B.n513 585
R490 B.n515 B.n160 585
R491 B.n517 B.n516 585
R492 B.n518 B.n159 585
R493 B.n520 B.n519 585
R494 B.n521 B.n158 585
R495 B.n523 B.n522 585
R496 B.n524 B.n157 585
R497 B.n526 B.n525 585
R498 B.n527 B.n156 585
R499 B.n529 B.n528 585
R500 B.n530 B.n155 585
R501 B.n532 B.n531 585
R502 B.n533 B.n154 585
R503 B.n535 B.n534 585
R504 B.n536 B.n153 585
R505 B.n538 B.n537 585
R506 B.n539 B.n152 585
R507 B.n541 B.n540 585
R508 B.n542 B.n151 585
R509 B.n544 B.n543 585
R510 B.n545 B.n150 585
R511 B.n547 B.n546 585
R512 B.n548 B.n149 585
R513 B.n550 B.n549 585
R514 B.n551 B.n148 585
R515 B.n553 B.n552 585
R516 B.n554 B.n147 585
R517 B.n556 B.n555 585
R518 B.n557 B.n146 585
R519 B.n559 B.n558 585
R520 B.n560 B.n145 585
R521 B.n562 B.n561 585
R522 B.n563 B.n144 585
R523 B.n565 B.n564 585
R524 B.n566 B.n143 585
R525 B.n568 B.n567 585
R526 B.n569 B.n142 585
R527 B.n571 B.n570 585
R528 B.n572 B.n141 585
R529 B.n574 B.n573 585
R530 B.n575 B.n140 585
R531 B.n577 B.n576 585
R532 B.n578 B.n139 585
R533 B.n580 B.n579 585
R534 B.n581 B.n138 585
R535 B.n583 B.n582 585
R536 B.n584 B.n137 585
R537 B.n586 B.n585 585
R538 B.n587 B.n136 585
R539 B.n589 B.n588 585
R540 B.n590 B.n135 585
R541 B.n592 B.n591 585
R542 B.n593 B.n134 585
R543 B.n595 B.n594 585
R544 B.n596 B.n133 585
R545 B.n598 B.n597 585
R546 B.n599 B.n132 585
R547 B.n601 B.n600 585
R548 B.n602 B.n131 585
R549 B.n604 B.n603 585
R550 B.n605 B.n130 585
R551 B.n607 B.n606 585
R552 B.n608 B.n129 585
R553 B.n610 B.n609 585
R554 B.n611 B.n128 585
R555 B.n613 B.n612 585
R556 B.n614 B.n127 585
R557 B.n616 B.n615 585
R558 B.n617 B.n126 585
R559 B.n619 B.n618 585
R560 B.n620 B.n125 585
R561 B.n622 B.n621 585
R562 B.n623 B.n124 585
R563 B.n625 B.n624 585
R564 B.n626 B.n123 585
R565 B.n628 B.n627 585
R566 B.n629 B.n122 585
R567 B.n631 B.n630 585
R568 B.n632 B.n121 585
R569 B.n634 B.n633 585
R570 B.n635 B.n120 585
R571 B.n637 B.n636 585
R572 B.n638 B.n119 585
R573 B.n640 B.n639 585
R574 B.n641 B.n118 585
R575 B.n643 B.n642 585
R576 B.n644 B.n117 585
R577 B.n646 B.n645 585
R578 B.n647 B.n116 585
R579 B.n649 B.n648 585
R580 B.n650 B.n115 585
R581 B.n652 B.n651 585
R582 B.n653 B.n114 585
R583 B.n655 B.n654 585
R584 B.n656 B.n113 585
R585 B.n658 B.n657 585
R586 B.n659 B.n112 585
R587 B.n661 B.n660 585
R588 B.n662 B.n111 585
R589 B.n664 B.n663 585
R590 B.n665 B.n110 585
R591 B.n667 B.n666 585
R592 B.n668 B.n109 585
R593 B.n670 B.n669 585
R594 B.n671 B.n108 585
R595 B.n673 B.n672 585
R596 B.n674 B.n107 585
R597 B.n676 B.n675 585
R598 B.n677 B.n106 585
R599 B.n679 B.n678 585
R600 B.n680 B.n105 585
R601 B.n682 B.n681 585
R602 B.n683 B.n104 585
R603 B.n685 B.n684 585
R604 B.n686 B.n103 585
R605 B.n688 B.n687 585
R606 B.n689 B.n102 585
R607 B.n691 B.n690 585
R608 B.n692 B.n101 585
R609 B.n694 B.n693 585
R610 B.n695 B.n100 585
R611 B.n697 B.n696 585
R612 B.n698 B.n99 585
R613 B.n700 B.n699 585
R614 B.n701 B.n98 585
R615 B.n703 B.n702 585
R616 B.n704 B.n97 585
R617 B.n706 B.n705 585
R618 B.n707 B.n96 585
R619 B.n709 B.n708 585
R620 B.n710 B.n95 585
R621 B.n712 B.n711 585
R622 B.n713 B.n94 585
R623 B.n715 B.n714 585
R624 B.n716 B.n93 585
R625 B.n873 B.n36 585
R626 B.n872 B.n871 585
R627 B.n870 B.n37 585
R628 B.n869 B.n868 585
R629 B.n867 B.n38 585
R630 B.n866 B.n865 585
R631 B.n864 B.n39 585
R632 B.n863 B.n862 585
R633 B.n861 B.n40 585
R634 B.n860 B.n859 585
R635 B.n858 B.n41 585
R636 B.n857 B.n856 585
R637 B.n855 B.n42 585
R638 B.n854 B.n853 585
R639 B.n852 B.n43 585
R640 B.n851 B.n850 585
R641 B.n849 B.n44 585
R642 B.n848 B.n847 585
R643 B.n846 B.n45 585
R644 B.n845 B.n844 585
R645 B.n843 B.n46 585
R646 B.n842 B.n841 585
R647 B.n840 B.n47 585
R648 B.n839 B.n838 585
R649 B.n837 B.n48 585
R650 B.n836 B.n835 585
R651 B.n834 B.n49 585
R652 B.n833 B.n832 585
R653 B.n831 B.n50 585
R654 B.n830 B.n829 585
R655 B.n828 B.n51 585
R656 B.n827 B.n826 585
R657 B.n825 B.n52 585
R658 B.n824 B.n823 585
R659 B.n822 B.n53 585
R660 B.n821 B.n820 585
R661 B.n819 B.n54 585
R662 B.n818 B.n817 585
R663 B.n816 B.n55 585
R664 B.n815 B.n814 585
R665 B.n813 B.n56 585
R666 B.n812 B.n811 585
R667 B.n810 B.n57 585
R668 B.n809 B.n808 585
R669 B.n807 B.n58 585
R670 B.n806 B.n805 585
R671 B.n804 B.n59 585
R672 B.n802 B.n801 585
R673 B.n800 B.n62 585
R674 B.n799 B.n798 585
R675 B.n797 B.n63 585
R676 B.n796 B.n795 585
R677 B.n794 B.n64 585
R678 B.n793 B.n792 585
R679 B.n791 B.n65 585
R680 B.n790 B.n789 585
R681 B.n788 B.n66 585
R682 B.n787 B.n786 585
R683 B.n785 B.n67 585
R684 B.n784 B.n783 585
R685 B.n782 B.n71 585
R686 B.n781 B.n780 585
R687 B.n779 B.n72 585
R688 B.n778 B.n777 585
R689 B.n776 B.n73 585
R690 B.n775 B.n774 585
R691 B.n773 B.n74 585
R692 B.n772 B.n771 585
R693 B.n770 B.n75 585
R694 B.n769 B.n768 585
R695 B.n767 B.n76 585
R696 B.n766 B.n765 585
R697 B.n764 B.n77 585
R698 B.n763 B.n762 585
R699 B.n761 B.n78 585
R700 B.n760 B.n759 585
R701 B.n758 B.n79 585
R702 B.n757 B.n756 585
R703 B.n755 B.n80 585
R704 B.n754 B.n753 585
R705 B.n752 B.n81 585
R706 B.n751 B.n750 585
R707 B.n749 B.n82 585
R708 B.n748 B.n747 585
R709 B.n746 B.n83 585
R710 B.n745 B.n744 585
R711 B.n743 B.n84 585
R712 B.n742 B.n741 585
R713 B.n740 B.n85 585
R714 B.n739 B.n738 585
R715 B.n737 B.n86 585
R716 B.n736 B.n735 585
R717 B.n734 B.n87 585
R718 B.n733 B.n732 585
R719 B.n731 B.n88 585
R720 B.n730 B.n729 585
R721 B.n728 B.n89 585
R722 B.n727 B.n726 585
R723 B.n725 B.n90 585
R724 B.n724 B.n723 585
R725 B.n722 B.n91 585
R726 B.n721 B.n720 585
R727 B.n719 B.n92 585
R728 B.n718 B.n717 585
R729 B.n875 B.n874 585
R730 B.n876 B.n35 585
R731 B.n878 B.n877 585
R732 B.n879 B.n34 585
R733 B.n881 B.n880 585
R734 B.n882 B.n33 585
R735 B.n884 B.n883 585
R736 B.n885 B.n32 585
R737 B.n887 B.n886 585
R738 B.n888 B.n31 585
R739 B.n890 B.n889 585
R740 B.n891 B.n30 585
R741 B.n893 B.n892 585
R742 B.n894 B.n29 585
R743 B.n896 B.n895 585
R744 B.n897 B.n28 585
R745 B.n899 B.n898 585
R746 B.n900 B.n27 585
R747 B.n902 B.n901 585
R748 B.n903 B.n26 585
R749 B.n905 B.n904 585
R750 B.n906 B.n25 585
R751 B.n908 B.n907 585
R752 B.n909 B.n24 585
R753 B.n911 B.n910 585
R754 B.n912 B.n23 585
R755 B.n914 B.n913 585
R756 B.n915 B.n22 585
R757 B.n917 B.n916 585
R758 B.n918 B.n21 585
R759 B.n920 B.n919 585
R760 B.n921 B.n20 585
R761 B.n923 B.n922 585
R762 B.n924 B.n19 585
R763 B.n926 B.n925 585
R764 B.n927 B.n18 585
R765 B.n929 B.n928 585
R766 B.n930 B.n17 585
R767 B.n932 B.n931 585
R768 B.n933 B.n16 585
R769 B.n935 B.n934 585
R770 B.n936 B.n15 585
R771 B.n938 B.n937 585
R772 B.n939 B.n14 585
R773 B.n941 B.n940 585
R774 B.n942 B.n13 585
R775 B.n944 B.n943 585
R776 B.n945 B.n12 585
R777 B.n947 B.n946 585
R778 B.n948 B.n11 585
R779 B.n950 B.n949 585
R780 B.n951 B.n10 585
R781 B.n953 B.n952 585
R782 B.n954 B.n9 585
R783 B.n956 B.n955 585
R784 B.n957 B.n8 585
R785 B.n959 B.n958 585
R786 B.n960 B.n7 585
R787 B.n962 B.n961 585
R788 B.n963 B.n6 585
R789 B.n965 B.n964 585
R790 B.n966 B.n5 585
R791 B.n968 B.n967 585
R792 B.n969 B.n4 585
R793 B.n971 B.n970 585
R794 B.n972 B.n3 585
R795 B.n974 B.n973 585
R796 B.n975 B.n0 585
R797 B.n2 B.n1 585
R798 B.n250 B.n249 585
R799 B.n252 B.n251 585
R800 B.n253 B.n248 585
R801 B.n255 B.n254 585
R802 B.n256 B.n247 585
R803 B.n258 B.n257 585
R804 B.n259 B.n246 585
R805 B.n261 B.n260 585
R806 B.n262 B.n245 585
R807 B.n264 B.n263 585
R808 B.n265 B.n244 585
R809 B.n267 B.n266 585
R810 B.n268 B.n243 585
R811 B.n270 B.n269 585
R812 B.n271 B.n242 585
R813 B.n273 B.n272 585
R814 B.n274 B.n241 585
R815 B.n276 B.n275 585
R816 B.n277 B.n240 585
R817 B.n279 B.n278 585
R818 B.n280 B.n239 585
R819 B.n282 B.n281 585
R820 B.n283 B.n238 585
R821 B.n285 B.n284 585
R822 B.n286 B.n237 585
R823 B.n288 B.n287 585
R824 B.n289 B.n236 585
R825 B.n291 B.n290 585
R826 B.n292 B.n235 585
R827 B.n294 B.n293 585
R828 B.n295 B.n234 585
R829 B.n297 B.n296 585
R830 B.n298 B.n233 585
R831 B.n300 B.n299 585
R832 B.n301 B.n232 585
R833 B.n303 B.n302 585
R834 B.n304 B.n231 585
R835 B.n306 B.n305 585
R836 B.n307 B.n230 585
R837 B.n309 B.n308 585
R838 B.n310 B.n229 585
R839 B.n312 B.n311 585
R840 B.n313 B.n228 585
R841 B.n315 B.n314 585
R842 B.n316 B.n227 585
R843 B.n318 B.n317 585
R844 B.n319 B.n226 585
R845 B.n321 B.n320 585
R846 B.n322 B.n225 585
R847 B.n324 B.n323 585
R848 B.n325 B.n224 585
R849 B.n327 B.n326 585
R850 B.n328 B.n223 585
R851 B.n330 B.n329 585
R852 B.n331 B.n222 585
R853 B.n333 B.n332 585
R854 B.n334 B.n221 585
R855 B.n336 B.n335 585
R856 B.n337 B.n220 585
R857 B.n339 B.n338 585
R858 B.n340 B.n219 585
R859 B.n342 B.n341 585
R860 B.n343 B.n218 585
R861 B.n345 B.n344 585
R862 B.n346 B.n217 585
R863 B.n348 B.n347 585
R864 B.n349 B.n216 585
R865 B.n351 B.n216 530.939
R866 B.n511 B.n162 530.939
R867 B.n717 B.n716 530.939
R868 B.n874 B.n873 530.939
R869 B.n191 B.t9 316.911
R870 B.n435 B.t6 316.911
R871 B.n68 B.t3 316.911
R872 B.n60 B.t0 316.911
R873 B.n977 B.n976 256.663
R874 B.n976 B.n975 235.042
R875 B.n976 B.n2 235.042
R876 B.n435 B.t7 179.456
R877 B.n68 B.t5 179.456
R878 B.n191 B.t10 179.439
R879 B.n60 B.t2 179.439
R880 B.n352 B.n351 163.367
R881 B.n353 B.n352 163.367
R882 B.n353 B.n214 163.367
R883 B.n357 B.n214 163.367
R884 B.n358 B.n357 163.367
R885 B.n359 B.n358 163.367
R886 B.n359 B.n212 163.367
R887 B.n363 B.n212 163.367
R888 B.n364 B.n363 163.367
R889 B.n365 B.n364 163.367
R890 B.n365 B.n210 163.367
R891 B.n369 B.n210 163.367
R892 B.n370 B.n369 163.367
R893 B.n371 B.n370 163.367
R894 B.n371 B.n208 163.367
R895 B.n375 B.n208 163.367
R896 B.n376 B.n375 163.367
R897 B.n377 B.n376 163.367
R898 B.n377 B.n206 163.367
R899 B.n381 B.n206 163.367
R900 B.n382 B.n381 163.367
R901 B.n383 B.n382 163.367
R902 B.n383 B.n204 163.367
R903 B.n387 B.n204 163.367
R904 B.n388 B.n387 163.367
R905 B.n389 B.n388 163.367
R906 B.n389 B.n202 163.367
R907 B.n393 B.n202 163.367
R908 B.n394 B.n393 163.367
R909 B.n395 B.n394 163.367
R910 B.n395 B.n200 163.367
R911 B.n399 B.n200 163.367
R912 B.n400 B.n399 163.367
R913 B.n401 B.n400 163.367
R914 B.n401 B.n198 163.367
R915 B.n405 B.n198 163.367
R916 B.n406 B.n405 163.367
R917 B.n407 B.n406 163.367
R918 B.n407 B.n196 163.367
R919 B.n411 B.n196 163.367
R920 B.n412 B.n411 163.367
R921 B.n413 B.n412 163.367
R922 B.n413 B.n194 163.367
R923 B.n417 B.n194 163.367
R924 B.n418 B.n417 163.367
R925 B.n419 B.n418 163.367
R926 B.n419 B.n190 163.367
R927 B.n424 B.n190 163.367
R928 B.n425 B.n424 163.367
R929 B.n426 B.n425 163.367
R930 B.n426 B.n188 163.367
R931 B.n430 B.n188 163.367
R932 B.n431 B.n430 163.367
R933 B.n432 B.n431 163.367
R934 B.n432 B.n186 163.367
R935 B.n439 B.n186 163.367
R936 B.n440 B.n439 163.367
R937 B.n441 B.n440 163.367
R938 B.n441 B.n184 163.367
R939 B.n445 B.n184 163.367
R940 B.n446 B.n445 163.367
R941 B.n447 B.n446 163.367
R942 B.n447 B.n182 163.367
R943 B.n451 B.n182 163.367
R944 B.n452 B.n451 163.367
R945 B.n453 B.n452 163.367
R946 B.n453 B.n180 163.367
R947 B.n457 B.n180 163.367
R948 B.n458 B.n457 163.367
R949 B.n459 B.n458 163.367
R950 B.n459 B.n178 163.367
R951 B.n463 B.n178 163.367
R952 B.n464 B.n463 163.367
R953 B.n465 B.n464 163.367
R954 B.n465 B.n176 163.367
R955 B.n469 B.n176 163.367
R956 B.n470 B.n469 163.367
R957 B.n471 B.n470 163.367
R958 B.n471 B.n174 163.367
R959 B.n475 B.n174 163.367
R960 B.n476 B.n475 163.367
R961 B.n477 B.n476 163.367
R962 B.n477 B.n172 163.367
R963 B.n481 B.n172 163.367
R964 B.n482 B.n481 163.367
R965 B.n483 B.n482 163.367
R966 B.n483 B.n170 163.367
R967 B.n487 B.n170 163.367
R968 B.n488 B.n487 163.367
R969 B.n489 B.n488 163.367
R970 B.n489 B.n168 163.367
R971 B.n493 B.n168 163.367
R972 B.n494 B.n493 163.367
R973 B.n495 B.n494 163.367
R974 B.n495 B.n166 163.367
R975 B.n499 B.n166 163.367
R976 B.n500 B.n499 163.367
R977 B.n501 B.n500 163.367
R978 B.n501 B.n164 163.367
R979 B.n505 B.n164 163.367
R980 B.n506 B.n505 163.367
R981 B.n507 B.n506 163.367
R982 B.n507 B.n162 163.367
R983 B.n716 B.n715 163.367
R984 B.n715 B.n94 163.367
R985 B.n711 B.n94 163.367
R986 B.n711 B.n710 163.367
R987 B.n710 B.n709 163.367
R988 B.n709 B.n96 163.367
R989 B.n705 B.n96 163.367
R990 B.n705 B.n704 163.367
R991 B.n704 B.n703 163.367
R992 B.n703 B.n98 163.367
R993 B.n699 B.n98 163.367
R994 B.n699 B.n698 163.367
R995 B.n698 B.n697 163.367
R996 B.n697 B.n100 163.367
R997 B.n693 B.n100 163.367
R998 B.n693 B.n692 163.367
R999 B.n692 B.n691 163.367
R1000 B.n691 B.n102 163.367
R1001 B.n687 B.n102 163.367
R1002 B.n687 B.n686 163.367
R1003 B.n686 B.n685 163.367
R1004 B.n685 B.n104 163.367
R1005 B.n681 B.n104 163.367
R1006 B.n681 B.n680 163.367
R1007 B.n680 B.n679 163.367
R1008 B.n679 B.n106 163.367
R1009 B.n675 B.n106 163.367
R1010 B.n675 B.n674 163.367
R1011 B.n674 B.n673 163.367
R1012 B.n673 B.n108 163.367
R1013 B.n669 B.n108 163.367
R1014 B.n669 B.n668 163.367
R1015 B.n668 B.n667 163.367
R1016 B.n667 B.n110 163.367
R1017 B.n663 B.n110 163.367
R1018 B.n663 B.n662 163.367
R1019 B.n662 B.n661 163.367
R1020 B.n661 B.n112 163.367
R1021 B.n657 B.n112 163.367
R1022 B.n657 B.n656 163.367
R1023 B.n656 B.n655 163.367
R1024 B.n655 B.n114 163.367
R1025 B.n651 B.n114 163.367
R1026 B.n651 B.n650 163.367
R1027 B.n650 B.n649 163.367
R1028 B.n649 B.n116 163.367
R1029 B.n645 B.n116 163.367
R1030 B.n645 B.n644 163.367
R1031 B.n644 B.n643 163.367
R1032 B.n643 B.n118 163.367
R1033 B.n639 B.n118 163.367
R1034 B.n639 B.n638 163.367
R1035 B.n638 B.n637 163.367
R1036 B.n637 B.n120 163.367
R1037 B.n633 B.n120 163.367
R1038 B.n633 B.n632 163.367
R1039 B.n632 B.n631 163.367
R1040 B.n631 B.n122 163.367
R1041 B.n627 B.n122 163.367
R1042 B.n627 B.n626 163.367
R1043 B.n626 B.n625 163.367
R1044 B.n625 B.n124 163.367
R1045 B.n621 B.n124 163.367
R1046 B.n621 B.n620 163.367
R1047 B.n620 B.n619 163.367
R1048 B.n619 B.n126 163.367
R1049 B.n615 B.n126 163.367
R1050 B.n615 B.n614 163.367
R1051 B.n614 B.n613 163.367
R1052 B.n613 B.n128 163.367
R1053 B.n609 B.n128 163.367
R1054 B.n609 B.n608 163.367
R1055 B.n608 B.n607 163.367
R1056 B.n607 B.n130 163.367
R1057 B.n603 B.n130 163.367
R1058 B.n603 B.n602 163.367
R1059 B.n602 B.n601 163.367
R1060 B.n601 B.n132 163.367
R1061 B.n597 B.n132 163.367
R1062 B.n597 B.n596 163.367
R1063 B.n596 B.n595 163.367
R1064 B.n595 B.n134 163.367
R1065 B.n591 B.n134 163.367
R1066 B.n591 B.n590 163.367
R1067 B.n590 B.n589 163.367
R1068 B.n589 B.n136 163.367
R1069 B.n585 B.n136 163.367
R1070 B.n585 B.n584 163.367
R1071 B.n584 B.n583 163.367
R1072 B.n583 B.n138 163.367
R1073 B.n579 B.n138 163.367
R1074 B.n579 B.n578 163.367
R1075 B.n578 B.n577 163.367
R1076 B.n577 B.n140 163.367
R1077 B.n573 B.n140 163.367
R1078 B.n573 B.n572 163.367
R1079 B.n572 B.n571 163.367
R1080 B.n571 B.n142 163.367
R1081 B.n567 B.n142 163.367
R1082 B.n567 B.n566 163.367
R1083 B.n566 B.n565 163.367
R1084 B.n565 B.n144 163.367
R1085 B.n561 B.n144 163.367
R1086 B.n561 B.n560 163.367
R1087 B.n560 B.n559 163.367
R1088 B.n559 B.n146 163.367
R1089 B.n555 B.n146 163.367
R1090 B.n555 B.n554 163.367
R1091 B.n554 B.n553 163.367
R1092 B.n553 B.n148 163.367
R1093 B.n549 B.n148 163.367
R1094 B.n549 B.n548 163.367
R1095 B.n548 B.n547 163.367
R1096 B.n547 B.n150 163.367
R1097 B.n543 B.n150 163.367
R1098 B.n543 B.n542 163.367
R1099 B.n542 B.n541 163.367
R1100 B.n541 B.n152 163.367
R1101 B.n537 B.n152 163.367
R1102 B.n537 B.n536 163.367
R1103 B.n536 B.n535 163.367
R1104 B.n535 B.n154 163.367
R1105 B.n531 B.n154 163.367
R1106 B.n531 B.n530 163.367
R1107 B.n530 B.n529 163.367
R1108 B.n529 B.n156 163.367
R1109 B.n525 B.n156 163.367
R1110 B.n525 B.n524 163.367
R1111 B.n524 B.n523 163.367
R1112 B.n523 B.n158 163.367
R1113 B.n519 B.n158 163.367
R1114 B.n519 B.n518 163.367
R1115 B.n518 B.n517 163.367
R1116 B.n517 B.n160 163.367
R1117 B.n513 B.n160 163.367
R1118 B.n513 B.n512 163.367
R1119 B.n512 B.n511 163.367
R1120 B.n873 B.n872 163.367
R1121 B.n872 B.n37 163.367
R1122 B.n868 B.n37 163.367
R1123 B.n868 B.n867 163.367
R1124 B.n867 B.n866 163.367
R1125 B.n866 B.n39 163.367
R1126 B.n862 B.n39 163.367
R1127 B.n862 B.n861 163.367
R1128 B.n861 B.n860 163.367
R1129 B.n860 B.n41 163.367
R1130 B.n856 B.n41 163.367
R1131 B.n856 B.n855 163.367
R1132 B.n855 B.n854 163.367
R1133 B.n854 B.n43 163.367
R1134 B.n850 B.n43 163.367
R1135 B.n850 B.n849 163.367
R1136 B.n849 B.n848 163.367
R1137 B.n848 B.n45 163.367
R1138 B.n844 B.n45 163.367
R1139 B.n844 B.n843 163.367
R1140 B.n843 B.n842 163.367
R1141 B.n842 B.n47 163.367
R1142 B.n838 B.n47 163.367
R1143 B.n838 B.n837 163.367
R1144 B.n837 B.n836 163.367
R1145 B.n836 B.n49 163.367
R1146 B.n832 B.n49 163.367
R1147 B.n832 B.n831 163.367
R1148 B.n831 B.n830 163.367
R1149 B.n830 B.n51 163.367
R1150 B.n826 B.n51 163.367
R1151 B.n826 B.n825 163.367
R1152 B.n825 B.n824 163.367
R1153 B.n824 B.n53 163.367
R1154 B.n820 B.n53 163.367
R1155 B.n820 B.n819 163.367
R1156 B.n819 B.n818 163.367
R1157 B.n818 B.n55 163.367
R1158 B.n814 B.n55 163.367
R1159 B.n814 B.n813 163.367
R1160 B.n813 B.n812 163.367
R1161 B.n812 B.n57 163.367
R1162 B.n808 B.n57 163.367
R1163 B.n808 B.n807 163.367
R1164 B.n807 B.n806 163.367
R1165 B.n806 B.n59 163.367
R1166 B.n801 B.n59 163.367
R1167 B.n801 B.n800 163.367
R1168 B.n800 B.n799 163.367
R1169 B.n799 B.n63 163.367
R1170 B.n795 B.n63 163.367
R1171 B.n795 B.n794 163.367
R1172 B.n794 B.n793 163.367
R1173 B.n793 B.n65 163.367
R1174 B.n789 B.n65 163.367
R1175 B.n789 B.n788 163.367
R1176 B.n788 B.n787 163.367
R1177 B.n787 B.n67 163.367
R1178 B.n783 B.n67 163.367
R1179 B.n783 B.n782 163.367
R1180 B.n782 B.n781 163.367
R1181 B.n781 B.n72 163.367
R1182 B.n777 B.n72 163.367
R1183 B.n777 B.n776 163.367
R1184 B.n776 B.n775 163.367
R1185 B.n775 B.n74 163.367
R1186 B.n771 B.n74 163.367
R1187 B.n771 B.n770 163.367
R1188 B.n770 B.n769 163.367
R1189 B.n769 B.n76 163.367
R1190 B.n765 B.n76 163.367
R1191 B.n765 B.n764 163.367
R1192 B.n764 B.n763 163.367
R1193 B.n763 B.n78 163.367
R1194 B.n759 B.n78 163.367
R1195 B.n759 B.n758 163.367
R1196 B.n758 B.n757 163.367
R1197 B.n757 B.n80 163.367
R1198 B.n753 B.n80 163.367
R1199 B.n753 B.n752 163.367
R1200 B.n752 B.n751 163.367
R1201 B.n751 B.n82 163.367
R1202 B.n747 B.n82 163.367
R1203 B.n747 B.n746 163.367
R1204 B.n746 B.n745 163.367
R1205 B.n745 B.n84 163.367
R1206 B.n741 B.n84 163.367
R1207 B.n741 B.n740 163.367
R1208 B.n740 B.n739 163.367
R1209 B.n739 B.n86 163.367
R1210 B.n735 B.n86 163.367
R1211 B.n735 B.n734 163.367
R1212 B.n734 B.n733 163.367
R1213 B.n733 B.n88 163.367
R1214 B.n729 B.n88 163.367
R1215 B.n729 B.n728 163.367
R1216 B.n728 B.n727 163.367
R1217 B.n727 B.n90 163.367
R1218 B.n723 B.n90 163.367
R1219 B.n723 B.n722 163.367
R1220 B.n722 B.n721 163.367
R1221 B.n721 B.n92 163.367
R1222 B.n717 B.n92 163.367
R1223 B.n874 B.n35 163.367
R1224 B.n878 B.n35 163.367
R1225 B.n879 B.n878 163.367
R1226 B.n880 B.n879 163.367
R1227 B.n880 B.n33 163.367
R1228 B.n884 B.n33 163.367
R1229 B.n885 B.n884 163.367
R1230 B.n886 B.n885 163.367
R1231 B.n886 B.n31 163.367
R1232 B.n890 B.n31 163.367
R1233 B.n891 B.n890 163.367
R1234 B.n892 B.n891 163.367
R1235 B.n892 B.n29 163.367
R1236 B.n896 B.n29 163.367
R1237 B.n897 B.n896 163.367
R1238 B.n898 B.n897 163.367
R1239 B.n898 B.n27 163.367
R1240 B.n902 B.n27 163.367
R1241 B.n903 B.n902 163.367
R1242 B.n904 B.n903 163.367
R1243 B.n904 B.n25 163.367
R1244 B.n908 B.n25 163.367
R1245 B.n909 B.n908 163.367
R1246 B.n910 B.n909 163.367
R1247 B.n910 B.n23 163.367
R1248 B.n914 B.n23 163.367
R1249 B.n915 B.n914 163.367
R1250 B.n916 B.n915 163.367
R1251 B.n916 B.n21 163.367
R1252 B.n920 B.n21 163.367
R1253 B.n921 B.n920 163.367
R1254 B.n922 B.n921 163.367
R1255 B.n922 B.n19 163.367
R1256 B.n926 B.n19 163.367
R1257 B.n927 B.n926 163.367
R1258 B.n928 B.n927 163.367
R1259 B.n928 B.n17 163.367
R1260 B.n932 B.n17 163.367
R1261 B.n933 B.n932 163.367
R1262 B.n934 B.n933 163.367
R1263 B.n934 B.n15 163.367
R1264 B.n938 B.n15 163.367
R1265 B.n939 B.n938 163.367
R1266 B.n940 B.n939 163.367
R1267 B.n940 B.n13 163.367
R1268 B.n944 B.n13 163.367
R1269 B.n945 B.n944 163.367
R1270 B.n946 B.n945 163.367
R1271 B.n946 B.n11 163.367
R1272 B.n950 B.n11 163.367
R1273 B.n951 B.n950 163.367
R1274 B.n952 B.n951 163.367
R1275 B.n952 B.n9 163.367
R1276 B.n956 B.n9 163.367
R1277 B.n957 B.n956 163.367
R1278 B.n958 B.n957 163.367
R1279 B.n958 B.n7 163.367
R1280 B.n962 B.n7 163.367
R1281 B.n963 B.n962 163.367
R1282 B.n964 B.n963 163.367
R1283 B.n964 B.n5 163.367
R1284 B.n968 B.n5 163.367
R1285 B.n969 B.n968 163.367
R1286 B.n970 B.n969 163.367
R1287 B.n970 B.n3 163.367
R1288 B.n974 B.n3 163.367
R1289 B.n975 B.n974 163.367
R1290 B.n250 B.n2 163.367
R1291 B.n251 B.n250 163.367
R1292 B.n251 B.n248 163.367
R1293 B.n255 B.n248 163.367
R1294 B.n256 B.n255 163.367
R1295 B.n257 B.n256 163.367
R1296 B.n257 B.n246 163.367
R1297 B.n261 B.n246 163.367
R1298 B.n262 B.n261 163.367
R1299 B.n263 B.n262 163.367
R1300 B.n263 B.n244 163.367
R1301 B.n267 B.n244 163.367
R1302 B.n268 B.n267 163.367
R1303 B.n269 B.n268 163.367
R1304 B.n269 B.n242 163.367
R1305 B.n273 B.n242 163.367
R1306 B.n274 B.n273 163.367
R1307 B.n275 B.n274 163.367
R1308 B.n275 B.n240 163.367
R1309 B.n279 B.n240 163.367
R1310 B.n280 B.n279 163.367
R1311 B.n281 B.n280 163.367
R1312 B.n281 B.n238 163.367
R1313 B.n285 B.n238 163.367
R1314 B.n286 B.n285 163.367
R1315 B.n287 B.n286 163.367
R1316 B.n287 B.n236 163.367
R1317 B.n291 B.n236 163.367
R1318 B.n292 B.n291 163.367
R1319 B.n293 B.n292 163.367
R1320 B.n293 B.n234 163.367
R1321 B.n297 B.n234 163.367
R1322 B.n298 B.n297 163.367
R1323 B.n299 B.n298 163.367
R1324 B.n299 B.n232 163.367
R1325 B.n303 B.n232 163.367
R1326 B.n304 B.n303 163.367
R1327 B.n305 B.n304 163.367
R1328 B.n305 B.n230 163.367
R1329 B.n309 B.n230 163.367
R1330 B.n310 B.n309 163.367
R1331 B.n311 B.n310 163.367
R1332 B.n311 B.n228 163.367
R1333 B.n315 B.n228 163.367
R1334 B.n316 B.n315 163.367
R1335 B.n317 B.n316 163.367
R1336 B.n317 B.n226 163.367
R1337 B.n321 B.n226 163.367
R1338 B.n322 B.n321 163.367
R1339 B.n323 B.n322 163.367
R1340 B.n323 B.n224 163.367
R1341 B.n327 B.n224 163.367
R1342 B.n328 B.n327 163.367
R1343 B.n329 B.n328 163.367
R1344 B.n329 B.n222 163.367
R1345 B.n333 B.n222 163.367
R1346 B.n334 B.n333 163.367
R1347 B.n335 B.n334 163.367
R1348 B.n335 B.n220 163.367
R1349 B.n339 B.n220 163.367
R1350 B.n340 B.n339 163.367
R1351 B.n341 B.n340 163.367
R1352 B.n341 B.n218 163.367
R1353 B.n345 B.n218 163.367
R1354 B.n346 B.n345 163.367
R1355 B.n347 B.n346 163.367
R1356 B.n347 B.n216 163.367
R1357 B.n436 B.t8 112.934
R1358 B.n69 B.t4 112.934
R1359 B.n192 B.t11 112.918
R1360 B.n61 B.t1 112.918
R1361 B.n192 B.n191 66.5217
R1362 B.n436 B.n435 66.5217
R1363 B.n69 B.n68 66.5217
R1364 B.n61 B.n60 66.5217
R1365 B.n421 B.n192 59.5399
R1366 B.n437 B.n436 59.5399
R1367 B.n70 B.n69 59.5399
R1368 B.n803 B.n61 59.5399
R1369 B.n875 B.n36 34.4981
R1370 B.n718 B.n93 34.4981
R1371 B.n510 B.n509 34.4981
R1372 B.n350 B.n349 34.4981
R1373 B B.n977 18.0485
R1374 B.n876 B.n875 10.6151
R1375 B.n877 B.n876 10.6151
R1376 B.n877 B.n34 10.6151
R1377 B.n881 B.n34 10.6151
R1378 B.n882 B.n881 10.6151
R1379 B.n883 B.n882 10.6151
R1380 B.n883 B.n32 10.6151
R1381 B.n887 B.n32 10.6151
R1382 B.n888 B.n887 10.6151
R1383 B.n889 B.n888 10.6151
R1384 B.n889 B.n30 10.6151
R1385 B.n893 B.n30 10.6151
R1386 B.n894 B.n893 10.6151
R1387 B.n895 B.n894 10.6151
R1388 B.n895 B.n28 10.6151
R1389 B.n899 B.n28 10.6151
R1390 B.n900 B.n899 10.6151
R1391 B.n901 B.n900 10.6151
R1392 B.n901 B.n26 10.6151
R1393 B.n905 B.n26 10.6151
R1394 B.n906 B.n905 10.6151
R1395 B.n907 B.n906 10.6151
R1396 B.n907 B.n24 10.6151
R1397 B.n911 B.n24 10.6151
R1398 B.n912 B.n911 10.6151
R1399 B.n913 B.n912 10.6151
R1400 B.n913 B.n22 10.6151
R1401 B.n917 B.n22 10.6151
R1402 B.n918 B.n917 10.6151
R1403 B.n919 B.n918 10.6151
R1404 B.n919 B.n20 10.6151
R1405 B.n923 B.n20 10.6151
R1406 B.n924 B.n923 10.6151
R1407 B.n925 B.n924 10.6151
R1408 B.n925 B.n18 10.6151
R1409 B.n929 B.n18 10.6151
R1410 B.n930 B.n929 10.6151
R1411 B.n931 B.n930 10.6151
R1412 B.n931 B.n16 10.6151
R1413 B.n935 B.n16 10.6151
R1414 B.n936 B.n935 10.6151
R1415 B.n937 B.n936 10.6151
R1416 B.n937 B.n14 10.6151
R1417 B.n941 B.n14 10.6151
R1418 B.n942 B.n941 10.6151
R1419 B.n943 B.n942 10.6151
R1420 B.n943 B.n12 10.6151
R1421 B.n947 B.n12 10.6151
R1422 B.n948 B.n947 10.6151
R1423 B.n949 B.n948 10.6151
R1424 B.n949 B.n10 10.6151
R1425 B.n953 B.n10 10.6151
R1426 B.n954 B.n953 10.6151
R1427 B.n955 B.n954 10.6151
R1428 B.n955 B.n8 10.6151
R1429 B.n959 B.n8 10.6151
R1430 B.n960 B.n959 10.6151
R1431 B.n961 B.n960 10.6151
R1432 B.n961 B.n6 10.6151
R1433 B.n965 B.n6 10.6151
R1434 B.n966 B.n965 10.6151
R1435 B.n967 B.n966 10.6151
R1436 B.n967 B.n4 10.6151
R1437 B.n971 B.n4 10.6151
R1438 B.n972 B.n971 10.6151
R1439 B.n973 B.n972 10.6151
R1440 B.n973 B.n0 10.6151
R1441 B.n871 B.n36 10.6151
R1442 B.n871 B.n870 10.6151
R1443 B.n870 B.n869 10.6151
R1444 B.n869 B.n38 10.6151
R1445 B.n865 B.n38 10.6151
R1446 B.n865 B.n864 10.6151
R1447 B.n864 B.n863 10.6151
R1448 B.n863 B.n40 10.6151
R1449 B.n859 B.n40 10.6151
R1450 B.n859 B.n858 10.6151
R1451 B.n858 B.n857 10.6151
R1452 B.n857 B.n42 10.6151
R1453 B.n853 B.n42 10.6151
R1454 B.n853 B.n852 10.6151
R1455 B.n852 B.n851 10.6151
R1456 B.n851 B.n44 10.6151
R1457 B.n847 B.n44 10.6151
R1458 B.n847 B.n846 10.6151
R1459 B.n846 B.n845 10.6151
R1460 B.n845 B.n46 10.6151
R1461 B.n841 B.n46 10.6151
R1462 B.n841 B.n840 10.6151
R1463 B.n840 B.n839 10.6151
R1464 B.n839 B.n48 10.6151
R1465 B.n835 B.n48 10.6151
R1466 B.n835 B.n834 10.6151
R1467 B.n834 B.n833 10.6151
R1468 B.n833 B.n50 10.6151
R1469 B.n829 B.n50 10.6151
R1470 B.n829 B.n828 10.6151
R1471 B.n828 B.n827 10.6151
R1472 B.n827 B.n52 10.6151
R1473 B.n823 B.n52 10.6151
R1474 B.n823 B.n822 10.6151
R1475 B.n822 B.n821 10.6151
R1476 B.n821 B.n54 10.6151
R1477 B.n817 B.n54 10.6151
R1478 B.n817 B.n816 10.6151
R1479 B.n816 B.n815 10.6151
R1480 B.n815 B.n56 10.6151
R1481 B.n811 B.n56 10.6151
R1482 B.n811 B.n810 10.6151
R1483 B.n810 B.n809 10.6151
R1484 B.n809 B.n58 10.6151
R1485 B.n805 B.n58 10.6151
R1486 B.n805 B.n804 10.6151
R1487 B.n802 B.n62 10.6151
R1488 B.n798 B.n62 10.6151
R1489 B.n798 B.n797 10.6151
R1490 B.n797 B.n796 10.6151
R1491 B.n796 B.n64 10.6151
R1492 B.n792 B.n64 10.6151
R1493 B.n792 B.n791 10.6151
R1494 B.n791 B.n790 10.6151
R1495 B.n790 B.n66 10.6151
R1496 B.n786 B.n785 10.6151
R1497 B.n785 B.n784 10.6151
R1498 B.n784 B.n71 10.6151
R1499 B.n780 B.n71 10.6151
R1500 B.n780 B.n779 10.6151
R1501 B.n779 B.n778 10.6151
R1502 B.n778 B.n73 10.6151
R1503 B.n774 B.n73 10.6151
R1504 B.n774 B.n773 10.6151
R1505 B.n773 B.n772 10.6151
R1506 B.n772 B.n75 10.6151
R1507 B.n768 B.n75 10.6151
R1508 B.n768 B.n767 10.6151
R1509 B.n767 B.n766 10.6151
R1510 B.n766 B.n77 10.6151
R1511 B.n762 B.n77 10.6151
R1512 B.n762 B.n761 10.6151
R1513 B.n761 B.n760 10.6151
R1514 B.n760 B.n79 10.6151
R1515 B.n756 B.n79 10.6151
R1516 B.n756 B.n755 10.6151
R1517 B.n755 B.n754 10.6151
R1518 B.n754 B.n81 10.6151
R1519 B.n750 B.n81 10.6151
R1520 B.n750 B.n749 10.6151
R1521 B.n749 B.n748 10.6151
R1522 B.n748 B.n83 10.6151
R1523 B.n744 B.n83 10.6151
R1524 B.n744 B.n743 10.6151
R1525 B.n743 B.n742 10.6151
R1526 B.n742 B.n85 10.6151
R1527 B.n738 B.n85 10.6151
R1528 B.n738 B.n737 10.6151
R1529 B.n737 B.n736 10.6151
R1530 B.n736 B.n87 10.6151
R1531 B.n732 B.n87 10.6151
R1532 B.n732 B.n731 10.6151
R1533 B.n731 B.n730 10.6151
R1534 B.n730 B.n89 10.6151
R1535 B.n726 B.n89 10.6151
R1536 B.n726 B.n725 10.6151
R1537 B.n725 B.n724 10.6151
R1538 B.n724 B.n91 10.6151
R1539 B.n720 B.n91 10.6151
R1540 B.n720 B.n719 10.6151
R1541 B.n719 B.n718 10.6151
R1542 B.n714 B.n93 10.6151
R1543 B.n714 B.n713 10.6151
R1544 B.n713 B.n712 10.6151
R1545 B.n712 B.n95 10.6151
R1546 B.n708 B.n95 10.6151
R1547 B.n708 B.n707 10.6151
R1548 B.n707 B.n706 10.6151
R1549 B.n706 B.n97 10.6151
R1550 B.n702 B.n97 10.6151
R1551 B.n702 B.n701 10.6151
R1552 B.n701 B.n700 10.6151
R1553 B.n700 B.n99 10.6151
R1554 B.n696 B.n99 10.6151
R1555 B.n696 B.n695 10.6151
R1556 B.n695 B.n694 10.6151
R1557 B.n694 B.n101 10.6151
R1558 B.n690 B.n101 10.6151
R1559 B.n690 B.n689 10.6151
R1560 B.n689 B.n688 10.6151
R1561 B.n688 B.n103 10.6151
R1562 B.n684 B.n103 10.6151
R1563 B.n684 B.n683 10.6151
R1564 B.n683 B.n682 10.6151
R1565 B.n682 B.n105 10.6151
R1566 B.n678 B.n105 10.6151
R1567 B.n678 B.n677 10.6151
R1568 B.n677 B.n676 10.6151
R1569 B.n676 B.n107 10.6151
R1570 B.n672 B.n107 10.6151
R1571 B.n672 B.n671 10.6151
R1572 B.n671 B.n670 10.6151
R1573 B.n670 B.n109 10.6151
R1574 B.n666 B.n109 10.6151
R1575 B.n666 B.n665 10.6151
R1576 B.n665 B.n664 10.6151
R1577 B.n664 B.n111 10.6151
R1578 B.n660 B.n111 10.6151
R1579 B.n660 B.n659 10.6151
R1580 B.n659 B.n658 10.6151
R1581 B.n658 B.n113 10.6151
R1582 B.n654 B.n113 10.6151
R1583 B.n654 B.n653 10.6151
R1584 B.n653 B.n652 10.6151
R1585 B.n652 B.n115 10.6151
R1586 B.n648 B.n115 10.6151
R1587 B.n648 B.n647 10.6151
R1588 B.n647 B.n646 10.6151
R1589 B.n646 B.n117 10.6151
R1590 B.n642 B.n117 10.6151
R1591 B.n642 B.n641 10.6151
R1592 B.n641 B.n640 10.6151
R1593 B.n640 B.n119 10.6151
R1594 B.n636 B.n119 10.6151
R1595 B.n636 B.n635 10.6151
R1596 B.n635 B.n634 10.6151
R1597 B.n634 B.n121 10.6151
R1598 B.n630 B.n121 10.6151
R1599 B.n630 B.n629 10.6151
R1600 B.n629 B.n628 10.6151
R1601 B.n628 B.n123 10.6151
R1602 B.n624 B.n123 10.6151
R1603 B.n624 B.n623 10.6151
R1604 B.n623 B.n622 10.6151
R1605 B.n622 B.n125 10.6151
R1606 B.n618 B.n125 10.6151
R1607 B.n618 B.n617 10.6151
R1608 B.n617 B.n616 10.6151
R1609 B.n616 B.n127 10.6151
R1610 B.n612 B.n127 10.6151
R1611 B.n612 B.n611 10.6151
R1612 B.n611 B.n610 10.6151
R1613 B.n610 B.n129 10.6151
R1614 B.n606 B.n129 10.6151
R1615 B.n606 B.n605 10.6151
R1616 B.n605 B.n604 10.6151
R1617 B.n604 B.n131 10.6151
R1618 B.n600 B.n131 10.6151
R1619 B.n600 B.n599 10.6151
R1620 B.n599 B.n598 10.6151
R1621 B.n598 B.n133 10.6151
R1622 B.n594 B.n133 10.6151
R1623 B.n594 B.n593 10.6151
R1624 B.n593 B.n592 10.6151
R1625 B.n592 B.n135 10.6151
R1626 B.n588 B.n135 10.6151
R1627 B.n588 B.n587 10.6151
R1628 B.n587 B.n586 10.6151
R1629 B.n586 B.n137 10.6151
R1630 B.n582 B.n137 10.6151
R1631 B.n582 B.n581 10.6151
R1632 B.n581 B.n580 10.6151
R1633 B.n580 B.n139 10.6151
R1634 B.n576 B.n139 10.6151
R1635 B.n576 B.n575 10.6151
R1636 B.n575 B.n574 10.6151
R1637 B.n574 B.n141 10.6151
R1638 B.n570 B.n141 10.6151
R1639 B.n570 B.n569 10.6151
R1640 B.n569 B.n568 10.6151
R1641 B.n568 B.n143 10.6151
R1642 B.n564 B.n143 10.6151
R1643 B.n564 B.n563 10.6151
R1644 B.n563 B.n562 10.6151
R1645 B.n562 B.n145 10.6151
R1646 B.n558 B.n145 10.6151
R1647 B.n558 B.n557 10.6151
R1648 B.n557 B.n556 10.6151
R1649 B.n556 B.n147 10.6151
R1650 B.n552 B.n147 10.6151
R1651 B.n552 B.n551 10.6151
R1652 B.n551 B.n550 10.6151
R1653 B.n550 B.n149 10.6151
R1654 B.n546 B.n149 10.6151
R1655 B.n546 B.n545 10.6151
R1656 B.n545 B.n544 10.6151
R1657 B.n544 B.n151 10.6151
R1658 B.n540 B.n151 10.6151
R1659 B.n540 B.n539 10.6151
R1660 B.n539 B.n538 10.6151
R1661 B.n538 B.n153 10.6151
R1662 B.n534 B.n153 10.6151
R1663 B.n534 B.n533 10.6151
R1664 B.n533 B.n532 10.6151
R1665 B.n532 B.n155 10.6151
R1666 B.n528 B.n155 10.6151
R1667 B.n528 B.n527 10.6151
R1668 B.n527 B.n526 10.6151
R1669 B.n526 B.n157 10.6151
R1670 B.n522 B.n157 10.6151
R1671 B.n522 B.n521 10.6151
R1672 B.n521 B.n520 10.6151
R1673 B.n520 B.n159 10.6151
R1674 B.n516 B.n159 10.6151
R1675 B.n516 B.n515 10.6151
R1676 B.n515 B.n514 10.6151
R1677 B.n514 B.n161 10.6151
R1678 B.n510 B.n161 10.6151
R1679 B.n249 B.n1 10.6151
R1680 B.n252 B.n249 10.6151
R1681 B.n253 B.n252 10.6151
R1682 B.n254 B.n253 10.6151
R1683 B.n254 B.n247 10.6151
R1684 B.n258 B.n247 10.6151
R1685 B.n259 B.n258 10.6151
R1686 B.n260 B.n259 10.6151
R1687 B.n260 B.n245 10.6151
R1688 B.n264 B.n245 10.6151
R1689 B.n265 B.n264 10.6151
R1690 B.n266 B.n265 10.6151
R1691 B.n266 B.n243 10.6151
R1692 B.n270 B.n243 10.6151
R1693 B.n271 B.n270 10.6151
R1694 B.n272 B.n271 10.6151
R1695 B.n272 B.n241 10.6151
R1696 B.n276 B.n241 10.6151
R1697 B.n277 B.n276 10.6151
R1698 B.n278 B.n277 10.6151
R1699 B.n278 B.n239 10.6151
R1700 B.n282 B.n239 10.6151
R1701 B.n283 B.n282 10.6151
R1702 B.n284 B.n283 10.6151
R1703 B.n284 B.n237 10.6151
R1704 B.n288 B.n237 10.6151
R1705 B.n289 B.n288 10.6151
R1706 B.n290 B.n289 10.6151
R1707 B.n290 B.n235 10.6151
R1708 B.n294 B.n235 10.6151
R1709 B.n295 B.n294 10.6151
R1710 B.n296 B.n295 10.6151
R1711 B.n296 B.n233 10.6151
R1712 B.n300 B.n233 10.6151
R1713 B.n301 B.n300 10.6151
R1714 B.n302 B.n301 10.6151
R1715 B.n302 B.n231 10.6151
R1716 B.n306 B.n231 10.6151
R1717 B.n307 B.n306 10.6151
R1718 B.n308 B.n307 10.6151
R1719 B.n308 B.n229 10.6151
R1720 B.n312 B.n229 10.6151
R1721 B.n313 B.n312 10.6151
R1722 B.n314 B.n313 10.6151
R1723 B.n314 B.n227 10.6151
R1724 B.n318 B.n227 10.6151
R1725 B.n319 B.n318 10.6151
R1726 B.n320 B.n319 10.6151
R1727 B.n320 B.n225 10.6151
R1728 B.n324 B.n225 10.6151
R1729 B.n325 B.n324 10.6151
R1730 B.n326 B.n325 10.6151
R1731 B.n326 B.n223 10.6151
R1732 B.n330 B.n223 10.6151
R1733 B.n331 B.n330 10.6151
R1734 B.n332 B.n331 10.6151
R1735 B.n332 B.n221 10.6151
R1736 B.n336 B.n221 10.6151
R1737 B.n337 B.n336 10.6151
R1738 B.n338 B.n337 10.6151
R1739 B.n338 B.n219 10.6151
R1740 B.n342 B.n219 10.6151
R1741 B.n343 B.n342 10.6151
R1742 B.n344 B.n343 10.6151
R1743 B.n344 B.n217 10.6151
R1744 B.n348 B.n217 10.6151
R1745 B.n349 B.n348 10.6151
R1746 B.n350 B.n215 10.6151
R1747 B.n354 B.n215 10.6151
R1748 B.n355 B.n354 10.6151
R1749 B.n356 B.n355 10.6151
R1750 B.n356 B.n213 10.6151
R1751 B.n360 B.n213 10.6151
R1752 B.n361 B.n360 10.6151
R1753 B.n362 B.n361 10.6151
R1754 B.n362 B.n211 10.6151
R1755 B.n366 B.n211 10.6151
R1756 B.n367 B.n366 10.6151
R1757 B.n368 B.n367 10.6151
R1758 B.n368 B.n209 10.6151
R1759 B.n372 B.n209 10.6151
R1760 B.n373 B.n372 10.6151
R1761 B.n374 B.n373 10.6151
R1762 B.n374 B.n207 10.6151
R1763 B.n378 B.n207 10.6151
R1764 B.n379 B.n378 10.6151
R1765 B.n380 B.n379 10.6151
R1766 B.n380 B.n205 10.6151
R1767 B.n384 B.n205 10.6151
R1768 B.n385 B.n384 10.6151
R1769 B.n386 B.n385 10.6151
R1770 B.n386 B.n203 10.6151
R1771 B.n390 B.n203 10.6151
R1772 B.n391 B.n390 10.6151
R1773 B.n392 B.n391 10.6151
R1774 B.n392 B.n201 10.6151
R1775 B.n396 B.n201 10.6151
R1776 B.n397 B.n396 10.6151
R1777 B.n398 B.n397 10.6151
R1778 B.n398 B.n199 10.6151
R1779 B.n402 B.n199 10.6151
R1780 B.n403 B.n402 10.6151
R1781 B.n404 B.n403 10.6151
R1782 B.n404 B.n197 10.6151
R1783 B.n408 B.n197 10.6151
R1784 B.n409 B.n408 10.6151
R1785 B.n410 B.n409 10.6151
R1786 B.n410 B.n195 10.6151
R1787 B.n414 B.n195 10.6151
R1788 B.n415 B.n414 10.6151
R1789 B.n416 B.n415 10.6151
R1790 B.n416 B.n193 10.6151
R1791 B.n420 B.n193 10.6151
R1792 B.n423 B.n422 10.6151
R1793 B.n423 B.n189 10.6151
R1794 B.n427 B.n189 10.6151
R1795 B.n428 B.n427 10.6151
R1796 B.n429 B.n428 10.6151
R1797 B.n429 B.n187 10.6151
R1798 B.n433 B.n187 10.6151
R1799 B.n434 B.n433 10.6151
R1800 B.n438 B.n434 10.6151
R1801 B.n442 B.n185 10.6151
R1802 B.n443 B.n442 10.6151
R1803 B.n444 B.n443 10.6151
R1804 B.n444 B.n183 10.6151
R1805 B.n448 B.n183 10.6151
R1806 B.n449 B.n448 10.6151
R1807 B.n450 B.n449 10.6151
R1808 B.n450 B.n181 10.6151
R1809 B.n454 B.n181 10.6151
R1810 B.n455 B.n454 10.6151
R1811 B.n456 B.n455 10.6151
R1812 B.n456 B.n179 10.6151
R1813 B.n460 B.n179 10.6151
R1814 B.n461 B.n460 10.6151
R1815 B.n462 B.n461 10.6151
R1816 B.n462 B.n177 10.6151
R1817 B.n466 B.n177 10.6151
R1818 B.n467 B.n466 10.6151
R1819 B.n468 B.n467 10.6151
R1820 B.n468 B.n175 10.6151
R1821 B.n472 B.n175 10.6151
R1822 B.n473 B.n472 10.6151
R1823 B.n474 B.n473 10.6151
R1824 B.n474 B.n173 10.6151
R1825 B.n478 B.n173 10.6151
R1826 B.n479 B.n478 10.6151
R1827 B.n480 B.n479 10.6151
R1828 B.n480 B.n171 10.6151
R1829 B.n484 B.n171 10.6151
R1830 B.n485 B.n484 10.6151
R1831 B.n486 B.n485 10.6151
R1832 B.n486 B.n169 10.6151
R1833 B.n490 B.n169 10.6151
R1834 B.n491 B.n490 10.6151
R1835 B.n492 B.n491 10.6151
R1836 B.n492 B.n167 10.6151
R1837 B.n496 B.n167 10.6151
R1838 B.n497 B.n496 10.6151
R1839 B.n498 B.n497 10.6151
R1840 B.n498 B.n165 10.6151
R1841 B.n502 B.n165 10.6151
R1842 B.n503 B.n502 10.6151
R1843 B.n504 B.n503 10.6151
R1844 B.n504 B.n163 10.6151
R1845 B.n508 B.n163 10.6151
R1846 B.n509 B.n508 10.6151
R1847 B.n804 B.n803 9.36635
R1848 B.n786 B.n70 9.36635
R1849 B.n421 B.n420 9.36635
R1850 B.n437 B.n185 9.36635
R1851 B.n977 B.n0 8.11757
R1852 B.n977 B.n1 8.11757
R1853 B.n803 B.n802 1.24928
R1854 B.n70 B.n66 1.24928
R1855 B.n422 B.n421 1.24928
R1856 B.n438 B.n437 1.24928
C0 VP VTAIL 13.4795f
C1 VTAIL w_n5086_n3752# 3.54873f
C2 VP VDD1 13.184f
C3 VDD1 w_n5086_n3752# 3.11307f
C4 VTAIL VDD1 11.385201f
C5 VDD2 B 2.96634f
C6 VN B 1.43724f
C7 VP B 2.55607f
C8 VDD2 VN 12.6952f
C9 w_n5086_n3752# B 11.9261f
C10 VDD2 VP 0.647957f
C11 VTAIL B 4.37308f
C12 VP VN 9.485661f
C13 VDD2 w_n5086_n3752# 3.28261f
C14 VN w_n5086_n3752# 11.0525f
C15 VDD1 B 2.82896f
C16 VDD2 VTAIL 11.439599f
C17 VN VTAIL 13.4652f
C18 VP w_n5086_n3752# 11.716299f
C19 VDD2 VDD1 2.50109f
C20 VN VDD1 0.154959f
C21 VDD2 VSUBS 2.39792f
C22 VDD1 VSUBS 2.213765f
C23 VTAIL VSUBS 1.490146f
C24 VN VSUBS 8.57845f
C25 VP VSUBS 4.954207f
C26 B VSUBS 6.14918f
C27 w_n5086_n3752# VSUBS 0.234302p
C28 B.n0 VSUBS 0.007614f
C29 B.n1 VSUBS 0.007614f
C30 B.n2 VSUBS 0.01126f
C31 B.n3 VSUBS 0.008629f
C32 B.n4 VSUBS 0.008629f
C33 B.n5 VSUBS 0.008629f
C34 B.n6 VSUBS 0.008629f
C35 B.n7 VSUBS 0.008629f
C36 B.n8 VSUBS 0.008629f
C37 B.n9 VSUBS 0.008629f
C38 B.n10 VSUBS 0.008629f
C39 B.n11 VSUBS 0.008629f
C40 B.n12 VSUBS 0.008629f
C41 B.n13 VSUBS 0.008629f
C42 B.n14 VSUBS 0.008629f
C43 B.n15 VSUBS 0.008629f
C44 B.n16 VSUBS 0.008629f
C45 B.n17 VSUBS 0.008629f
C46 B.n18 VSUBS 0.008629f
C47 B.n19 VSUBS 0.008629f
C48 B.n20 VSUBS 0.008629f
C49 B.n21 VSUBS 0.008629f
C50 B.n22 VSUBS 0.008629f
C51 B.n23 VSUBS 0.008629f
C52 B.n24 VSUBS 0.008629f
C53 B.n25 VSUBS 0.008629f
C54 B.n26 VSUBS 0.008629f
C55 B.n27 VSUBS 0.008629f
C56 B.n28 VSUBS 0.008629f
C57 B.n29 VSUBS 0.008629f
C58 B.n30 VSUBS 0.008629f
C59 B.n31 VSUBS 0.008629f
C60 B.n32 VSUBS 0.008629f
C61 B.n33 VSUBS 0.008629f
C62 B.n34 VSUBS 0.008629f
C63 B.n35 VSUBS 0.008629f
C64 B.n36 VSUBS 0.021468f
C65 B.n37 VSUBS 0.008629f
C66 B.n38 VSUBS 0.008629f
C67 B.n39 VSUBS 0.008629f
C68 B.n40 VSUBS 0.008629f
C69 B.n41 VSUBS 0.008629f
C70 B.n42 VSUBS 0.008629f
C71 B.n43 VSUBS 0.008629f
C72 B.n44 VSUBS 0.008629f
C73 B.n45 VSUBS 0.008629f
C74 B.n46 VSUBS 0.008629f
C75 B.n47 VSUBS 0.008629f
C76 B.n48 VSUBS 0.008629f
C77 B.n49 VSUBS 0.008629f
C78 B.n50 VSUBS 0.008629f
C79 B.n51 VSUBS 0.008629f
C80 B.n52 VSUBS 0.008629f
C81 B.n53 VSUBS 0.008629f
C82 B.n54 VSUBS 0.008629f
C83 B.n55 VSUBS 0.008629f
C84 B.n56 VSUBS 0.008629f
C85 B.n57 VSUBS 0.008629f
C86 B.n58 VSUBS 0.008629f
C87 B.n59 VSUBS 0.008629f
C88 B.t1 VSUBS 0.5675f
C89 B.t2 VSUBS 0.596746f
C90 B.t0 VSUBS 2.42936f
C91 B.n60 VSUBS 0.3332f
C92 B.n61 VSUBS 0.091196f
C93 B.n62 VSUBS 0.008629f
C94 B.n63 VSUBS 0.008629f
C95 B.n64 VSUBS 0.008629f
C96 B.n65 VSUBS 0.008629f
C97 B.n66 VSUBS 0.004822f
C98 B.n67 VSUBS 0.008629f
C99 B.t4 VSUBS 0.567487f
C100 B.t5 VSUBS 0.596734f
C101 B.t3 VSUBS 2.42936f
C102 B.n68 VSUBS 0.333211f
C103 B.n69 VSUBS 0.09121f
C104 B.n70 VSUBS 0.019992f
C105 B.n71 VSUBS 0.008629f
C106 B.n72 VSUBS 0.008629f
C107 B.n73 VSUBS 0.008629f
C108 B.n74 VSUBS 0.008629f
C109 B.n75 VSUBS 0.008629f
C110 B.n76 VSUBS 0.008629f
C111 B.n77 VSUBS 0.008629f
C112 B.n78 VSUBS 0.008629f
C113 B.n79 VSUBS 0.008629f
C114 B.n80 VSUBS 0.008629f
C115 B.n81 VSUBS 0.008629f
C116 B.n82 VSUBS 0.008629f
C117 B.n83 VSUBS 0.008629f
C118 B.n84 VSUBS 0.008629f
C119 B.n85 VSUBS 0.008629f
C120 B.n86 VSUBS 0.008629f
C121 B.n87 VSUBS 0.008629f
C122 B.n88 VSUBS 0.008629f
C123 B.n89 VSUBS 0.008629f
C124 B.n90 VSUBS 0.008629f
C125 B.n91 VSUBS 0.008629f
C126 B.n92 VSUBS 0.008629f
C127 B.n93 VSUBS 0.020408f
C128 B.n94 VSUBS 0.008629f
C129 B.n95 VSUBS 0.008629f
C130 B.n96 VSUBS 0.008629f
C131 B.n97 VSUBS 0.008629f
C132 B.n98 VSUBS 0.008629f
C133 B.n99 VSUBS 0.008629f
C134 B.n100 VSUBS 0.008629f
C135 B.n101 VSUBS 0.008629f
C136 B.n102 VSUBS 0.008629f
C137 B.n103 VSUBS 0.008629f
C138 B.n104 VSUBS 0.008629f
C139 B.n105 VSUBS 0.008629f
C140 B.n106 VSUBS 0.008629f
C141 B.n107 VSUBS 0.008629f
C142 B.n108 VSUBS 0.008629f
C143 B.n109 VSUBS 0.008629f
C144 B.n110 VSUBS 0.008629f
C145 B.n111 VSUBS 0.008629f
C146 B.n112 VSUBS 0.008629f
C147 B.n113 VSUBS 0.008629f
C148 B.n114 VSUBS 0.008629f
C149 B.n115 VSUBS 0.008629f
C150 B.n116 VSUBS 0.008629f
C151 B.n117 VSUBS 0.008629f
C152 B.n118 VSUBS 0.008629f
C153 B.n119 VSUBS 0.008629f
C154 B.n120 VSUBS 0.008629f
C155 B.n121 VSUBS 0.008629f
C156 B.n122 VSUBS 0.008629f
C157 B.n123 VSUBS 0.008629f
C158 B.n124 VSUBS 0.008629f
C159 B.n125 VSUBS 0.008629f
C160 B.n126 VSUBS 0.008629f
C161 B.n127 VSUBS 0.008629f
C162 B.n128 VSUBS 0.008629f
C163 B.n129 VSUBS 0.008629f
C164 B.n130 VSUBS 0.008629f
C165 B.n131 VSUBS 0.008629f
C166 B.n132 VSUBS 0.008629f
C167 B.n133 VSUBS 0.008629f
C168 B.n134 VSUBS 0.008629f
C169 B.n135 VSUBS 0.008629f
C170 B.n136 VSUBS 0.008629f
C171 B.n137 VSUBS 0.008629f
C172 B.n138 VSUBS 0.008629f
C173 B.n139 VSUBS 0.008629f
C174 B.n140 VSUBS 0.008629f
C175 B.n141 VSUBS 0.008629f
C176 B.n142 VSUBS 0.008629f
C177 B.n143 VSUBS 0.008629f
C178 B.n144 VSUBS 0.008629f
C179 B.n145 VSUBS 0.008629f
C180 B.n146 VSUBS 0.008629f
C181 B.n147 VSUBS 0.008629f
C182 B.n148 VSUBS 0.008629f
C183 B.n149 VSUBS 0.008629f
C184 B.n150 VSUBS 0.008629f
C185 B.n151 VSUBS 0.008629f
C186 B.n152 VSUBS 0.008629f
C187 B.n153 VSUBS 0.008629f
C188 B.n154 VSUBS 0.008629f
C189 B.n155 VSUBS 0.008629f
C190 B.n156 VSUBS 0.008629f
C191 B.n157 VSUBS 0.008629f
C192 B.n158 VSUBS 0.008629f
C193 B.n159 VSUBS 0.008629f
C194 B.n160 VSUBS 0.008629f
C195 B.n161 VSUBS 0.008629f
C196 B.n162 VSUBS 0.021468f
C197 B.n163 VSUBS 0.008629f
C198 B.n164 VSUBS 0.008629f
C199 B.n165 VSUBS 0.008629f
C200 B.n166 VSUBS 0.008629f
C201 B.n167 VSUBS 0.008629f
C202 B.n168 VSUBS 0.008629f
C203 B.n169 VSUBS 0.008629f
C204 B.n170 VSUBS 0.008629f
C205 B.n171 VSUBS 0.008629f
C206 B.n172 VSUBS 0.008629f
C207 B.n173 VSUBS 0.008629f
C208 B.n174 VSUBS 0.008629f
C209 B.n175 VSUBS 0.008629f
C210 B.n176 VSUBS 0.008629f
C211 B.n177 VSUBS 0.008629f
C212 B.n178 VSUBS 0.008629f
C213 B.n179 VSUBS 0.008629f
C214 B.n180 VSUBS 0.008629f
C215 B.n181 VSUBS 0.008629f
C216 B.n182 VSUBS 0.008629f
C217 B.n183 VSUBS 0.008629f
C218 B.n184 VSUBS 0.008629f
C219 B.n185 VSUBS 0.008121f
C220 B.n186 VSUBS 0.008629f
C221 B.n187 VSUBS 0.008629f
C222 B.n188 VSUBS 0.008629f
C223 B.n189 VSUBS 0.008629f
C224 B.n190 VSUBS 0.008629f
C225 B.t11 VSUBS 0.5675f
C226 B.t10 VSUBS 0.596746f
C227 B.t9 VSUBS 2.42936f
C228 B.n191 VSUBS 0.3332f
C229 B.n192 VSUBS 0.091196f
C230 B.n193 VSUBS 0.008629f
C231 B.n194 VSUBS 0.008629f
C232 B.n195 VSUBS 0.008629f
C233 B.n196 VSUBS 0.008629f
C234 B.n197 VSUBS 0.008629f
C235 B.n198 VSUBS 0.008629f
C236 B.n199 VSUBS 0.008629f
C237 B.n200 VSUBS 0.008629f
C238 B.n201 VSUBS 0.008629f
C239 B.n202 VSUBS 0.008629f
C240 B.n203 VSUBS 0.008629f
C241 B.n204 VSUBS 0.008629f
C242 B.n205 VSUBS 0.008629f
C243 B.n206 VSUBS 0.008629f
C244 B.n207 VSUBS 0.008629f
C245 B.n208 VSUBS 0.008629f
C246 B.n209 VSUBS 0.008629f
C247 B.n210 VSUBS 0.008629f
C248 B.n211 VSUBS 0.008629f
C249 B.n212 VSUBS 0.008629f
C250 B.n213 VSUBS 0.008629f
C251 B.n214 VSUBS 0.008629f
C252 B.n215 VSUBS 0.008629f
C253 B.n216 VSUBS 0.020408f
C254 B.n217 VSUBS 0.008629f
C255 B.n218 VSUBS 0.008629f
C256 B.n219 VSUBS 0.008629f
C257 B.n220 VSUBS 0.008629f
C258 B.n221 VSUBS 0.008629f
C259 B.n222 VSUBS 0.008629f
C260 B.n223 VSUBS 0.008629f
C261 B.n224 VSUBS 0.008629f
C262 B.n225 VSUBS 0.008629f
C263 B.n226 VSUBS 0.008629f
C264 B.n227 VSUBS 0.008629f
C265 B.n228 VSUBS 0.008629f
C266 B.n229 VSUBS 0.008629f
C267 B.n230 VSUBS 0.008629f
C268 B.n231 VSUBS 0.008629f
C269 B.n232 VSUBS 0.008629f
C270 B.n233 VSUBS 0.008629f
C271 B.n234 VSUBS 0.008629f
C272 B.n235 VSUBS 0.008629f
C273 B.n236 VSUBS 0.008629f
C274 B.n237 VSUBS 0.008629f
C275 B.n238 VSUBS 0.008629f
C276 B.n239 VSUBS 0.008629f
C277 B.n240 VSUBS 0.008629f
C278 B.n241 VSUBS 0.008629f
C279 B.n242 VSUBS 0.008629f
C280 B.n243 VSUBS 0.008629f
C281 B.n244 VSUBS 0.008629f
C282 B.n245 VSUBS 0.008629f
C283 B.n246 VSUBS 0.008629f
C284 B.n247 VSUBS 0.008629f
C285 B.n248 VSUBS 0.008629f
C286 B.n249 VSUBS 0.008629f
C287 B.n250 VSUBS 0.008629f
C288 B.n251 VSUBS 0.008629f
C289 B.n252 VSUBS 0.008629f
C290 B.n253 VSUBS 0.008629f
C291 B.n254 VSUBS 0.008629f
C292 B.n255 VSUBS 0.008629f
C293 B.n256 VSUBS 0.008629f
C294 B.n257 VSUBS 0.008629f
C295 B.n258 VSUBS 0.008629f
C296 B.n259 VSUBS 0.008629f
C297 B.n260 VSUBS 0.008629f
C298 B.n261 VSUBS 0.008629f
C299 B.n262 VSUBS 0.008629f
C300 B.n263 VSUBS 0.008629f
C301 B.n264 VSUBS 0.008629f
C302 B.n265 VSUBS 0.008629f
C303 B.n266 VSUBS 0.008629f
C304 B.n267 VSUBS 0.008629f
C305 B.n268 VSUBS 0.008629f
C306 B.n269 VSUBS 0.008629f
C307 B.n270 VSUBS 0.008629f
C308 B.n271 VSUBS 0.008629f
C309 B.n272 VSUBS 0.008629f
C310 B.n273 VSUBS 0.008629f
C311 B.n274 VSUBS 0.008629f
C312 B.n275 VSUBS 0.008629f
C313 B.n276 VSUBS 0.008629f
C314 B.n277 VSUBS 0.008629f
C315 B.n278 VSUBS 0.008629f
C316 B.n279 VSUBS 0.008629f
C317 B.n280 VSUBS 0.008629f
C318 B.n281 VSUBS 0.008629f
C319 B.n282 VSUBS 0.008629f
C320 B.n283 VSUBS 0.008629f
C321 B.n284 VSUBS 0.008629f
C322 B.n285 VSUBS 0.008629f
C323 B.n286 VSUBS 0.008629f
C324 B.n287 VSUBS 0.008629f
C325 B.n288 VSUBS 0.008629f
C326 B.n289 VSUBS 0.008629f
C327 B.n290 VSUBS 0.008629f
C328 B.n291 VSUBS 0.008629f
C329 B.n292 VSUBS 0.008629f
C330 B.n293 VSUBS 0.008629f
C331 B.n294 VSUBS 0.008629f
C332 B.n295 VSUBS 0.008629f
C333 B.n296 VSUBS 0.008629f
C334 B.n297 VSUBS 0.008629f
C335 B.n298 VSUBS 0.008629f
C336 B.n299 VSUBS 0.008629f
C337 B.n300 VSUBS 0.008629f
C338 B.n301 VSUBS 0.008629f
C339 B.n302 VSUBS 0.008629f
C340 B.n303 VSUBS 0.008629f
C341 B.n304 VSUBS 0.008629f
C342 B.n305 VSUBS 0.008629f
C343 B.n306 VSUBS 0.008629f
C344 B.n307 VSUBS 0.008629f
C345 B.n308 VSUBS 0.008629f
C346 B.n309 VSUBS 0.008629f
C347 B.n310 VSUBS 0.008629f
C348 B.n311 VSUBS 0.008629f
C349 B.n312 VSUBS 0.008629f
C350 B.n313 VSUBS 0.008629f
C351 B.n314 VSUBS 0.008629f
C352 B.n315 VSUBS 0.008629f
C353 B.n316 VSUBS 0.008629f
C354 B.n317 VSUBS 0.008629f
C355 B.n318 VSUBS 0.008629f
C356 B.n319 VSUBS 0.008629f
C357 B.n320 VSUBS 0.008629f
C358 B.n321 VSUBS 0.008629f
C359 B.n322 VSUBS 0.008629f
C360 B.n323 VSUBS 0.008629f
C361 B.n324 VSUBS 0.008629f
C362 B.n325 VSUBS 0.008629f
C363 B.n326 VSUBS 0.008629f
C364 B.n327 VSUBS 0.008629f
C365 B.n328 VSUBS 0.008629f
C366 B.n329 VSUBS 0.008629f
C367 B.n330 VSUBS 0.008629f
C368 B.n331 VSUBS 0.008629f
C369 B.n332 VSUBS 0.008629f
C370 B.n333 VSUBS 0.008629f
C371 B.n334 VSUBS 0.008629f
C372 B.n335 VSUBS 0.008629f
C373 B.n336 VSUBS 0.008629f
C374 B.n337 VSUBS 0.008629f
C375 B.n338 VSUBS 0.008629f
C376 B.n339 VSUBS 0.008629f
C377 B.n340 VSUBS 0.008629f
C378 B.n341 VSUBS 0.008629f
C379 B.n342 VSUBS 0.008629f
C380 B.n343 VSUBS 0.008629f
C381 B.n344 VSUBS 0.008629f
C382 B.n345 VSUBS 0.008629f
C383 B.n346 VSUBS 0.008629f
C384 B.n347 VSUBS 0.008629f
C385 B.n348 VSUBS 0.008629f
C386 B.n349 VSUBS 0.020408f
C387 B.n350 VSUBS 0.021468f
C388 B.n351 VSUBS 0.021468f
C389 B.n352 VSUBS 0.008629f
C390 B.n353 VSUBS 0.008629f
C391 B.n354 VSUBS 0.008629f
C392 B.n355 VSUBS 0.008629f
C393 B.n356 VSUBS 0.008629f
C394 B.n357 VSUBS 0.008629f
C395 B.n358 VSUBS 0.008629f
C396 B.n359 VSUBS 0.008629f
C397 B.n360 VSUBS 0.008629f
C398 B.n361 VSUBS 0.008629f
C399 B.n362 VSUBS 0.008629f
C400 B.n363 VSUBS 0.008629f
C401 B.n364 VSUBS 0.008629f
C402 B.n365 VSUBS 0.008629f
C403 B.n366 VSUBS 0.008629f
C404 B.n367 VSUBS 0.008629f
C405 B.n368 VSUBS 0.008629f
C406 B.n369 VSUBS 0.008629f
C407 B.n370 VSUBS 0.008629f
C408 B.n371 VSUBS 0.008629f
C409 B.n372 VSUBS 0.008629f
C410 B.n373 VSUBS 0.008629f
C411 B.n374 VSUBS 0.008629f
C412 B.n375 VSUBS 0.008629f
C413 B.n376 VSUBS 0.008629f
C414 B.n377 VSUBS 0.008629f
C415 B.n378 VSUBS 0.008629f
C416 B.n379 VSUBS 0.008629f
C417 B.n380 VSUBS 0.008629f
C418 B.n381 VSUBS 0.008629f
C419 B.n382 VSUBS 0.008629f
C420 B.n383 VSUBS 0.008629f
C421 B.n384 VSUBS 0.008629f
C422 B.n385 VSUBS 0.008629f
C423 B.n386 VSUBS 0.008629f
C424 B.n387 VSUBS 0.008629f
C425 B.n388 VSUBS 0.008629f
C426 B.n389 VSUBS 0.008629f
C427 B.n390 VSUBS 0.008629f
C428 B.n391 VSUBS 0.008629f
C429 B.n392 VSUBS 0.008629f
C430 B.n393 VSUBS 0.008629f
C431 B.n394 VSUBS 0.008629f
C432 B.n395 VSUBS 0.008629f
C433 B.n396 VSUBS 0.008629f
C434 B.n397 VSUBS 0.008629f
C435 B.n398 VSUBS 0.008629f
C436 B.n399 VSUBS 0.008629f
C437 B.n400 VSUBS 0.008629f
C438 B.n401 VSUBS 0.008629f
C439 B.n402 VSUBS 0.008629f
C440 B.n403 VSUBS 0.008629f
C441 B.n404 VSUBS 0.008629f
C442 B.n405 VSUBS 0.008629f
C443 B.n406 VSUBS 0.008629f
C444 B.n407 VSUBS 0.008629f
C445 B.n408 VSUBS 0.008629f
C446 B.n409 VSUBS 0.008629f
C447 B.n410 VSUBS 0.008629f
C448 B.n411 VSUBS 0.008629f
C449 B.n412 VSUBS 0.008629f
C450 B.n413 VSUBS 0.008629f
C451 B.n414 VSUBS 0.008629f
C452 B.n415 VSUBS 0.008629f
C453 B.n416 VSUBS 0.008629f
C454 B.n417 VSUBS 0.008629f
C455 B.n418 VSUBS 0.008629f
C456 B.n419 VSUBS 0.008629f
C457 B.n420 VSUBS 0.008121f
C458 B.n421 VSUBS 0.019992f
C459 B.n422 VSUBS 0.004822f
C460 B.n423 VSUBS 0.008629f
C461 B.n424 VSUBS 0.008629f
C462 B.n425 VSUBS 0.008629f
C463 B.n426 VSUBS 0.008629f
C464 B.n427 VSUBS 0.008629f
C465 B.n428 VSUBS 0.008629f
C466 B.n429 VSUBS 0.008629f
C467 B.n430 VSUBS 0.008629f
C468 B.n431 VSUBS 0.008629f
C469 B.n432 VSUBS 0.008629f
C470 B.n433 VSUBS 0.008629f
C471 B.n434 VSUBS 0.008629f
C472 B.t8 VSUBS 0.567487f
C473 B.t7 VSUBS 0.596734f
C474 B.t6 VSUBS 2.42936f
C475 B.n435 VSUBS 0.333211f
C476 B.n436 VSUBS 0.09121f
C477 B.n437 VSUBS 0.019992f
C478 B.n438 VSUBS 0.004822f
C479 B.n439 VSUBS 0.008629f
C480 B.n440 VSUBS 0.008629f
C481 B.n441 VSUBS 0.008629f
C482 B.n442 VSUBS 0.008629f
C483 B.n443 VSUBS 0.008629f
C484 B.n444 VSUBS 0.008629f
C485 B.n445 VSUBS 0.008629f
C486 B.n446 VSUBS 0.008629f
C487 B.n447 VSUBS 0.008629f
C488 B.n448 VSUBS 0.008629f
C489 B.n449 VSUBS 0.008629f
C490 B.n450 VSUBS 0.008629f
C491 B.n451 VSUBS 0.008629f
C492 B.n452 VSUBS 0.008629f
C493 B.n453 VSUBS 0.008629f
C494 B.n454 VSUBS 0.008629f
C495 B.n455 VSUBS 0.008629f
C496 B.n456 VSUBS 0.008629f
C497 B.n457 VSUBS 0.008629f
C498 B.n458 VSUBS 0.008629f
C499 B.n459 VSUBS 0.008629f
C500 B.n460 VSUBS 0.008629f
C501 B.n461 VSUBS 0.008629f
C502 B.n462 VSUBS 0.008629f
C503 B.n463 VSUBS 0.008629f
C504 B.n464 VSUBS 0.008629f
C505 B.n465 VSUBS 0.008629f
C506 B.n466 VSUBS 0.008629f
C507 B.n467 VSUBS 0.008629f
C508 B.n468 VSUBS 0.008629f
C509 B.n469 VSUBS 0.008629f
C510 B.n470 VSUBS 0.008629f
C511 B.n471 VSUBS 0.008629f
C512 B.n472 VSUBS 0.008629f
C513 B.n473 VSUBS 0.008629f
C514 B.n474 VSUBS 0.008629f
C515 B.n475 VSUBS 0.008629f
C516 B.n476 VSUBS 0.008629f
C517 B.n477 VSUBS 0.008629f
C518 B.n478 VSUBS 0.008629f
C519 B.n479 VSUBS 0.008629f
C520 B.n480 VSUBS 0.008629f
C521 B.n481 VSUBS 0.008629f
C522 B.n482 VSUBS 0.008629f
C523 B.n483 VSUBS 0.008629f
C524 B.n484 VSUBS 0.008629f
C525 B.n485 VSUBS 0.008629f
C526 B.n486 VSUBS 0.008629f
C527 B.n487 VSUBS 0.008629f
C528 B.n488 VSUBS 0.008629f
C529 B.n489 VSUBS 0.008629f
C530 B.n490 VSUBS 0.008629f
C531 B.n491 VSUBS 0.008629f
C532 B.n492 VSUBS 0.008629f
C533 B.n493 VSUBS 0.008629f
C534 B.n494 VSUBS 0.008629f
C535 B.n495 VSUBS 0.008629f
C536 B.n496 VSUBS 0.008629f
C537 B.n497 VSUBS 0.008629f
C538 B.n498 VSUBS 0.008629f
C539 B.n499 VSUBS 0.008629f
C540 B.n500 VSUBS 0.008629f
C541 B.n501 VSUBS 0.008629f
C542 B.n502 VSUBS 0.008629f
C543 B.n503 VSUBS 0.008629f
C544 B.n504 VSUBS 0.008629f
C545 B.n505 VSUBS 0.008629f
C546 B.n506 VSUBS 0.008629f
C547 B.n507 VSUBS 0.008629f
C548 B.n508 VSUBS 0.008629f
C549 B.n509 VSUBS 0.020502f
C550 B.n510 VSUBS 0.021374f
C551 B.n511 VSUBS 0.020408f
C552 B.n512 VSUBS 0.008629f
C553 B.n513 VSUBS 0.008629f
C554 B.n514 VSUBS 0.008629f
C555 B.n515 VSUBS 0.008629f
C556 B.n516 VSUBS 0.008629f
C557 B.n517 VSUBS 0.008629f
C558 B.n518 VSUBS 0.008629f
C559 B.n519 VSUBS 0.008629f
C560 B.n520 VSUBS 0.008629f
C561 B.n521 VSUBS 0.008629f
C562 B.n522 VSUBS 0.008629f
C563 B.n523 VSUBS 0.008629f
C564 B.n524 VSUBS 0.008629f
C565 B.n525 VSUBS 0.008629f
C566 B.n526 VSUBS 0.008629f
C567 B.n527 VSUBS 0.008629f
C568 B.n528 VSUBS 0.008629f
C569 B.n529 VSUBS 0.008629f
C570 B.n530 VSUBS 0.008629f
C571 B.n531 VSUBS 0.008629f
C572 B.n532 VSUBS 0.008629f
C573 B.n533 VSUBS 0.008629f
C574 B.n534 VSUBS 0.008629f
C575 B.n535 VSUBS 0.008629f
C576 B.n536 VSUBS 0.008629f
C577 B.n537 VSUBS 0.008629f
C578 B.n538 VSUBS 0.008629f
C579 B.n539 VSUBS 0.008629f
C580 B.n540 VSUBS 0.008629f
C581 B.n541 VSUBS 0.008629f
C582 B.n542 VSUBS 0.008629f
C583 B.n543 VSUBS 0.008629f
C584 B.n544 VSUBS 0.008629f
C585 B.n545 VSUBS 0.008629f
C586 B.n546 VSUBS 0.008629f
C587 B.n547 VSUBS 0.008629f
C588 B.n548 VSUBS 0.008629f
C589 B.n549 VSUBS 0.008629f
C590 B.n550 VSUBS 0.008629f
C591 B.n551 VSUBS 0.008629f
C592 B.n552 VSUBS 0.008629f
C593 B.n553 VSUBS 0.008629f
C594 B.n554 VSUBS 0.008629f
C595 B.n555 VSUBS 0.008629f
C596 B.n556 VSUBS 0.008629f
C597 B.n557 VSUBS 0.008629f
C598 B.n558 VSUBS 0.008629f
C599 B.n559 VSUBS 0.008629f
C600 B.n560 VSUBS 0.008629f
C601 B.n561 VSUBS 0.008629f
C602 B.n562 VSUBS 0.008629f
C603 B.n563 VSUBS 0.008629f
C604 B.n564 VSUBS 0.008629f
C605 B.n565 VSUBS 0.008629f
C606 B.n566 VSUBS 0.008629f
C607 B.n567 VSUBS 0.008629f
C608 B.n568 VSUBS 0.008629f
C609 B.n569 VSUBS 0.008629f
C610 B.n570 VSUBS 0.008629f
C611 B.n571 VSUBS 0.008629f
C612 B.n572 VSUBS 0.008629f
C613 B.n573 VSUBS 0.008629f
C614 B.n574 VSUBS 0.008629f
C615 B.n575 VSUBS 0.008629f
C616 B.n576 VSUBS 0.008629f
C617 B.n577 VSUBS 0.008629f
C618 B.n578 VSUBS 0.008629f
C619 B.n579 VSUBS 0.008629f
C620 B.n580 VSUBS 0.008629f
C621 B.n581 VSUBS 0.008629f
C622 B.n582 VSUBS 0.008629f
C623 B.n583 VSUBS 0.008629f
C624 B.n584 VSUBS 0.008629f
C625 B.n585 VSUBS 0.008629f
C626 B.n586 VSUBS 0.008629f
C627 B.n587 VSUBS 0.008629f
C628 B.n588 VSUBS 0.008629f
C629 B.n589 VSUBS 0.008629f
C630 B.n590 VSUBS 0.008629f
C631 B.n591 VSUBS 0.008629f
C632 B.n592 VSUBS 0.008629f
C633 B.n593 VSUBS 0.008629f
C634 B.n594 VSUBS 0.008629f
C635 B.n595 VSUBS 0.008629f
C636 B.n596 VSUBS 0.008629f
C637 B.n597 VSUBS 0.008629f
C638 B.n598 VSUBS 0.008629f
C639 B.n599 VSUBS 0.008629f
C640 B.n600 VSUBS 0.008629f
C641 B.n601 VSUBS 0.008629f
C642 B.n602 VSUBS 0.008629f
C643 B.n603 VSUBS 0.008629f
C644 B.n604 VSUBS 0.008629f
C645 B.n605 VSUBS 0.008629f
C646 B.n606 VSUBS 0.008629f
C647 B.n607 VSUBS 0.008629f
C648 B.n608 VSUBS 0.008629f
C649 B.n609 VSUBS 0.008629f
C650 B.n610 VSUBS 0.008629f
C651 B.n611 VSUBS 0.008629f
C652 B.n612 VSUBS 0.008629f
C653 B.n613 VSUBS 0.008629f
C654 B.n614 VSUBS 0.008629f
C655 B.n615 VSUBS 0.008629f
C656 B.n616 VSUBS 0.008629f
C657 B.n617 VSUBS 0.008629f
C658 B.n618 VSUBS 0.008629f
C659 B.n619 VSUBS 0.008629f
C660 B.n620 VSUBS 0.008629f
C661 B.n621 VSUBS 0.008629f
C662 B.n622 VSUBS 0.008629f
C663 B.n623 VSUBS 0.008629f
C664 B.n624 VSUBS 0.008629f
C665 B.n625 VSUBS 0.008629f
C666 B.n626 VSUBS 0.008629f
C667 B.n627 VSUBS 0.008629f
C668 B.n628 VSUBS 0.008629f
C669 B.n629 VSUBS 0.008629f
C670 B.n630 VSUBS 0.008629f
C671 B.n631 VSUBS 0.008629f
C672 B.n632 VSUBS 0.008629f
C673 B.n633 VSUBS 0.008629f
C674 B.n634 VSUBS 0.008629f
C675 B.n635 VSUBS 0.008629f
C676 B.n636 VSUBS 0.008629f
C677 B.n637 VSUBS 0.008629f
C678 B.n638 VSUBS 0.008629f
C679 B.n639 VSUBS 0.008629f
C680 B.n640 VSUBS 0.008629f
C681 B.n641 VSUBS 0.008629f
C682 B.n642 VSUBS 0.008629f
C683 B.n643 VSUBS 0.008629f
C684 B.n644 VSUBS 0.008629f
C685 B.n645 VSUBS 0.008629f
C686 B.n646 VSUBS 0.008629f
C687 B.n647 VSUBS 0.008629f
C688 B.n648 VSUBS 0.008629f
C689 B.n649 VSUBS 0.008629f
C690 B.n650 VSUBS 0.008629f
C691 B.n651 VSUBS 0.008629f
C692 B.n652 VSUBS 0.008629f
C693 B.n653 VSUBS 0.008629f
C694 B.n654 VSUBS 0.008629f
C695 B.n655 VSUBS 0.008629f
C696 B.n656 VSUBS 0.008629f
C697 B.n657 VSUBS 0.008629f
C698 B.n658 VSUBS 0.008629f
C699 B.n659 VSUBS 0.008629f
C700 B.n660 VSUBS 0.008629f
C701 B.n661 VSUBS 0.008629f
C702 B.n662 VSUBS 0.008629f
C703 B.n663 VSUBS 0.008629f
C704 B.n664 VSUBS 0.008629f
C705 B.n665 VSUBS 0.008629f
C706 B.n666 VSUBS 0.008629f
C707 B.n667 VSUBS 0.008629f
C708 B.n668 VSUBS 0.008629f
C709 B.n669 VSUBS 0.008629f
C710 B.n670 VSUBS 0.008629f
C711 B.n671 VSUBS 0.008629f
C712 B.n672 VSUBS 0.008629f
C713 B.n673 VSUBS 0.008629f
C714 B.n674 VSUBS 0.008629f
C715 B.n675 VSUBS 0.008629f
C716 B.n676 VSUBS 0.008629f
C717 B.n677 VSUBS 0.008629f
C718 B.n678 VSUBS 0.008629f
C719 B.n679 VSUBS 0.008629f
C720 B.n680 VSUBS 0.008629f
C721 B.n681 VSUBS 0.008629f
C722 B.n682 VSUBS 0.008629f
C723 B.n683 VSUBS 0.008629f
C724 B.n684 VSUBS 0.008629f
C725 B.n685 VSUBS 0.008629f
C726 B.n686 VSUBS 0.008629f
C727 B.n687 VSUBS 0.008629f
C728 B.n688 VSUBS 0.008629f
C729 B.n689 VSUBS 0.008629f
C730 B.n690 VSUBS 0.008629f
C731 B.n691 VSUBS 0.008629f
C732 B.n692 VSUBS 0.008629f
C733 B.n693 VSUBS 0.008629f
C734 B.n694 VSUBS 0.008629f
C735 B.n695 VSUBS 0.008629f
C736 B.n696 VSUBS 0.008629f
C737 B.n697 VSUBS 0.008629f
C738 B.n698 VSUBS 0.008629f
C739 B.n699 VSUBS 0.008629f
C740 B.n700 VSUBS 0.008629f
C741 B.n701 VSUBS 0.008629f
C742 B.n702 VSUBS 0.008629f
C743 B.n703 VSUBS 0.008629f
C744 B.n704 VSUBS 0.008629f
C745 B.n705 VSUBS 0.008629f
C746 B.n706 VSUBS 0.008629f
C747 B.n707 VSUBS 0.008629f
C748 B.n708 VSUBS 0.008629f
C749 B.n709 VSUBS 0.008629f
C750 B.n710 VSUBS 0.008629f
C751 B.n711 VSUBS 0.008629f
C752 B.n712 VSUBS 0.008629f
C753 B.n713 VSUBS 0.008629f
C754 B.n714 VSUBS 0.008629f
C755 B.n715 VSUBS 0.008629f
C756 B.n716 VSUBS 0.020408f
C757 B.n717 VSUBS 0.021468f
C758 B.n718 VSUBS 0.021468f
C759 B.n719 VSUBS 0.008629f
C760 B.n720 VSUBS 0.008629f
C761 B.n721 VSUBS 0.008629f
C762 B.n722 VSUBS 0.008629f
C763 B.n723 VSUBS 0.008629f
C764 B.n724 VSUBS 0.008629f
C765 B.n725 VSUBS 0.008629f
C766 B.n726 VSUBS 0.008629f
C767 B.n727 VSUBS 0.008629f
C768 B.n728 VSUBS 0.008629f
C769 B.n729 VSUBS 0.008629f
C770 B.n730 VSUBS 0.008629f
C771 B.n731 VSUBS 0.008629f
C772 B.n732 VSUBS 0.008629f
C773 B.n733 VSUBS 0.008629f
C774 B.n734 VSUBS 0.008629f
C775 B.n735 VSUBS 0.008629f
C776 B.n736 VSUBS 0.008629f
C777 B.n737 VSUBS 0.008629f
C778 B.n738 VSUBS 0.008629f
C779 B.n739 VSUBS 0.008629f
C780 B.n740 VSUBS 0.008629f
C781 B.n741 VSUBS 0.008629f
C782 B.n742 VSUBS 0.008629f
C783 B.n743 VSUBS 0.008629f
C784 B.n744 VSUBS 0.008629f
C785 B.n745 VSUBS 0.008629f
C786 B.n746 VSUBS 0.008629f
C787 B.n747 VSUBS 0.008629f
C788 B.n748 VSUBS 0.008629f
C789 B.n749 VSUBS 0.008629f
C790 B.n750 VSUBS 0.008629f
C791 B.n751 VSUBS 0.008629f
C792 B.n752 VSUBS 0.008629f
C793 B.n753 VSUBS 0.008629f
C794 B.n754 VSUBS 0.008629f
C795 B.n755 VSUBS 0.008629f
C796 B.n756 VSUBS 0.008629f
C797 B.n757 VSUBS 0.008629f
C798 B.n758 VSUBS 0.008629f
C799 B.n759 VSUBS 0.008629f
C800 B.n760 VSUBS 0.008629f
C801 B.n761 VSUBS 0.008629f
C802 B.n762 VSUBS 0.008629f
C803 B.n763 VSUBS 0.008629f
C804 B.n764 VSUBS 0.008629f
C805 B.n765 VSUBS 0.008629f
C806 B.n766 VSUBS 0.008629f
C807 B.n767 VSUBS 0.008629f
C808 B.n768 VSUBS 0.008629f
C809 B.n769 VSUBS 0.008629f
C810 B.n770 VSUBS 0.008629f
C811 B.n771 VSUBS 0.008629f
C812 B.n772 VSUBS 0.008629f
C813 B.n773 VSUBS 0.008629f
C814 B.n774 VSUBS 0.008629f
C815 B.n775 VSUBS 0.008629f
C816 B.n776 VSUBS 0.008629f
C817 B.n777 VSUBS 0.008629f
C818 B.n778 VSUBS 0.008629f
C819 B.n779 VSUBS 0.008629f
C820 B.n780 VSUBS 0.008629f
C821 B.n781 VSUBS 0.008629f
C822 B.n782 VSUBS 0.008629f
C823 B.n783 VSUBS 0.008629f
C824 B.n784 VSUBS 0.008629f
C825 B.n785 VSUBS 0.008629f
C826 B.n786 VSUBS 0.008121f
C827 B.n787 VSUBS 0.008629f
C828 B.n788 VSUBS 0.008629f
C829 B.n789 VSUBS 0.008629f
C830 B.n790 VSUBS 0.008629f
C831 B.n791 VSUBS 0.008629f
C832 B.n792 VSUBS 0.008629f
C833 B.n793 VSUBS 0.008629f
C834 B.n794 VSUBS 0.008629f
C835 B.n795 VSUBS 0.008629f
C836 B.n796 VSUBS 0.008629f
C837 B.n797 VSUBS 0.008629f
C838 B.n798 VSUBS 0.008629f
C839 B.n799 VSUBS 0.008629f
C840 B.n800 VSUBS 0.008629f
C841 B.n801 VSUBS 0.008629f
C842 B.n802 VSUBS 0.004822f
C843 B.n803 VSUBS 0.019992f
C844 B.n804 VSUBS 0.008121f
C845 B.n805 VSUBS 0.008629f
C846 B.n806 VSUBS 0.008629f
C847 B.n807 VSUBS 0.008629f
C848 B.n808 VSUBS 0.008629f
C849 B.n809 VSUBS 0.008629f
C850 B.n810 VSUBS 0.008629f
C851 B.n811 VSUBS 0.008629f
C852 B.n812 VSUBS 0.008629f
C853 B.n813 VSUBS 0.008629f
C854 B.n814 VSUBS 0.008629f
C855 B.n815 VSUBS 0.008629f
C856 B.n816 VSUBS 0.008629f
C857 B.n817 VSUBS 0.008629f
C858 B.n818 VSUBS 0.008629f
C859 B.n819 VSUBS 0.008629f
C860 B.n820 VSUBS 0.008629f
C861 B.n821 VSUBS 0.008629f
C862 B.n822 VSUBS 0.008629f
C863 B.n823 VSUBS 0.008629f
C864 B.n824 VSUBS 0.008629f
C865 B.n825 VSUBS 0.008629f
C866 B.n826 VSUBS 0.008629f
C867 B.n827 VSUBS 0.008629f
C868 B.n828 VSUBS 0.008629f
C869 B.n829 VSUBS 0.008629f
C870 B.n830 VSUBS 0.008629f
C871 B.n831 VSUBS 0.008629f
C872 B.n832 VSUBS 0.008629f
C873 B.n833 VSUBS 0.008629f
C874 B.n834 VSUBS 0.008629f
C875 B.n835 VSUBS 0.008629f
C876 B.n836 VSUBS 0.008629f
C877 B.n837 VSUBS 0.008629f
C878 B.n838 VSUBS 0.008629f
C879 B.n839 VSUBS 0.008629f
C880 B.n840 VSUBS 0.008629f
C881 B.n841 VSUBS 0.008629f
C882 B.n842 VSUBS 0.008629f
C883 B.n843 VSUBS 0.008629f
C884 B.n844 VSUBS 0.008629f
C885 B.n845 VSUBS 0.008629f
C886 B.n846 VSUBS 0.008629f
C887 B.n847 VSUBS 0.008629f
C888 B.n848 VSUBS 0.008629f
C889 B.n849 VSUBS 0.008629f
C890 B.n850 VSUBS 0.008629f
C891 B.n851 VSUBS 0.008629f
C892 B.n852 VSUBS 0.008629f
C893 B.n853 VSUBS 0.008629f
C894 B.n854 VSUBS 0.008629f
C895 B.n855 VSUBS 0.008629f
C896 B.n856 VSUBS 0.008629f
C897 B.n857 VSUBS 0.008629f
C898 B.n858 VSUBS 0.008629f
C899 B.n859 VSUBS 0.008629f
C900 B.n860 VSUBS 0.008629f
C901 B.n861 VSUBS 0.008629f
C902 B.n862 VSUBS 0.008629f
C903 B.n863 VSUBS 0.008629f
C904 B.n864 VSUBS 0.008629f
C905 B.n865 VSUBS 0.008629f
C906 B.n866 VSUBS 0.008629f
C907 B.n867 VSUBS 0.008629f
C908 B.n868 VSUBS 0.008629f
C909 B.n869 VSUBS 0.008629f
C910 B.n870 VSUBS 0.008629f
C911 B.n871 VSUBS 0.008629f
C912 B.n872 VSUBS 0.008629f
C913 B.n873 VSUBS 0.021468f
C914 B.n874 VSUBS 0.020408f
C915 B.n875 VSUBS 0.020408f
C916 B.n876 VSUBS 0.008629f
C917 B.n877 VSUBS 0.008629f
C918 B.n878 VSUBS 0.008629f
C919 B.n879 VSUBS 0.008629f
C920 B.n880 VSUBS 0.008629f
C921 B.n881 VSUBS 0.008629f
C922 B.n882 VSUBS 0.008629f
C923 B.n883 VSUBS 0.008629f
C924 B.n884 VSUBS 0.008629f
C925 B.n885 VSUBS 0.008629f
C926 B.n886 VSUBS 0.008629f
C927 B.n887 VSUBS 0.008629f
C928 B.n888 VSUBS 0.008629f
C929 B.n889 VSUBS 0.008629f
C930 B.n890 VSUBS 0.008629f
C931 B.n891 VSUBS 0.008629f
C932 B.n892 VSUBS 0.008629f
C933 B.n893 VSUBS 0.008629f
C934 B.n894 VSUBS 0.008629f
C935 B.n895 VSUBS 0.008629f
C936 B.n896 VSUBS 0.008629f
C937 B.n897 VSUBS 0.008629f
C938 B.n898 VSUBS 0.008629f
C939 B.n899 VSUBS 0.008629f
C940 B.n900 VSUBS 0.008629f
C941 B.n901 VSUBS 0.008629f
C942 B.n902 VSUBS 0.008629f
C943 B.n903 VSUBS 0.008629f
C944 B.n904 VSUBS 0.008629f
C945 B.n905 VSUBS 0.008629f
C946 B.n906 VSUBS 0.008629f
C947 B.n907 VSUBS 0.008629f
C948 B.n908 VSUBS 0.008629f
C949 B.n909 VSUBS 0.008629f
C950 B.n910 VSUBS 0.008629f
C951 B.n911 VSUBS 0.008629f
C952 B.n912 VSUBS 0.008629f
C953 B.n913 VSUBS 0.008629f
C954 B.n914 VSUBS 0.008629f
C955 B.n915 VSUBS 0.008629f
C956 B.n916 VSUBS 0.008629f
C957 B.n917 VSUBS 0.008629f
C958 B.n918 VSUBS 0.008629f
C959 B.n919 VSUBS 0.008629f
C960 B.n920 VSUBS 0.008629f
C961 B.n921 VSUBS 0.008629f
C962 B.n922 VSUBS 0.008629f
C963 B.n923 VSUBS 0.008629f
C964 B.n924 VSUBS 0.008629f
C965 B.n925 VSUBS 0.008629f
C966 B.n926 VSUBS 0.008629f
C967 B.n927 VSUBS 0.008629f
C968 B.n928 VSUBS 0.008629f
C969 B.n929 VSUBS 0.008629f
C970 B.n930 VSUBS 0.008629f
C971 B.n931 VSUBS 0.008629f
C972 B.n932 VSUBS 0.008629f
C973 B.n933 VSUBS 0.008629f
C974 B.n934 VSUBS 0.008629f
C975 B.n935 VSUBS 0.008629f
C976 B.n936 VSUBS 0.008629f
C977 B.n937 VSUBS 0.008629f
C978 B.n938 VSUBS 0.008629f
C979 B.n939 VSUBS 0.008629f
C980 B.n940 VSUBS 0.008629f
C981 B.n941 VSUBS 0.008629f
C982 B.n942 VSUBS 0.008629f
C983 B.n943 VSUBS 0.008629f
C984 B.n944 VSUBS 0.008629f
C985 B.n945 VSUBS 0.008629f
C986 B.n946 VSUBS 0.008629f
C987 B.n947 VSUBS 0.008629f
C988 B.n948 VSUBS 0.008629f
C989 B.n949 VSUBS 0.008629f
C990 B.n950 VSUBS 0.008629f
C991 B.n951 VSUBS 0.008629f
C992 B.n952 VSUBS 0.008629f
C993 B.n953 VSUBS 0.008629f
C994 B.n954 VSUBS 0.008629f
C995 B.n955 VSUBS 0.008629f
C996 B.n956 VSUBS 0.008629f
C997 B.n957 VSUBS 0.008629f
C998 B.n958 VSUBS 0.008629f
C999 B.n959 VSUBS 0.008629f
C1000 B.n960 VSUBS 0.008629f
C1001 B.n961 VSUBS 0.008629f
C1002 B.n962 VSUBS 0.008629f
C1003 B.n963 VSUBS 0.008629f
C1004 B.n964 VSUBS 0.008629f
C1005 B.n965 VSUBS 0.008629f
C1006 B.n966 VSUBS 0.008629f
C1007 B.n967 VSUBS 0.008629f
C1008 B.n968 VSUBS 0.008629f
C1009 B.n969 VSUBS 0.008629f
C1010 B.n970 VSUBS 0.008629f
C1011 B.n971 VSUBS 0.008629f
C1012 B.n972 VSUBS 0.008629f
C1013 B.n973 VSUBS 0.008629f
C1014 B.n974 VSUBS 0.008629f
C1015 B.n975 VSUBS 0.01126f
C1016 B.n976 VSUBS 0.011995f
C1017 B.n977 VSUBS 0.023853f
C1018 VDD2.t9 VSUBS 3.45247f
C1019 VDD2.t8 VSUBS 0.328024f
C1020 VDD2.t3 VSUBS 0.328024f
C1021 VDD2.n0 VSUBS 2.62083f
C1022 VDD2.n1 VSUBS 1.86246f
C1023 VDD2.t2 VSUBS 0.328024f
C1024 VDD2.t5 VSUBS 0.328024f
C1025 VDD2.n2 VSUBS 2.65236f
C1026 VDD2.n3 VSUBS 4.24355f
C1027 VDD2.t1 VSUBS 3.41525f
C1028 VDD2.n4 VSUBS 4.48623f
C1029 VDD2.t4 VSUBS 0.328024f
C1030 VDD2.t6 VSUBS 0.328024f
C1031 VDD2.n5 VSUBS 2.62083f
C1032 VDD2.n6 VSUBS 0.936991f
C1033 VDD2.t0 VSUBS 0.328024f
C1034 VDD2.t7 VSUBS 0.328024f
C1035 VDD2.n7 VSUBS 2.6523f
C1036 VN.t4 VSUBS 2.90784f
C1037 VN.n0 VSUBS 1.11119f
C1038 VN.n1 VSUBS 0.024635f
C1039 VN.n2 VSUBS 0.027399f
C1040 VN.n3 VSUBS 0.024635f
C1041 VN.t7 VSUBS 2.90784f
C1042 VN.n4 VSUBS 1.01561f
C1043 VN.n5 VSUBS 0.024635f
C1044 VN.n6 VSUBS 0.033425f
C1045 VN.n7 VSUBS 0.024635f
C1046 VN.t6 VSUBS 2.90784f
C1047 VN.n8 VSUBS 0.045684f
C1048 VN.n9 VSUBS 0.024635f
C1049 VN.n10 VSUBS 0.045684f
C1050 VN.t0 VSUBS 3.1877f
C1051 VN.n11 VSUBS 1.05131f
C1052 VN.t1 VSUBS 2.90784f
C1053 VN.n12 VSUBS 1.10342f
C1054 VN.n13 VSUBS 0.042526f
C1055 VN.n14 VSUBS 0.282061f
C1056 VN.n15 VSUBS 0.024635f
C1057 VN.n16 VSUBS 0.024635f
C1058 VN.n17 VSUBS 0.038197f
C1059 VN.n18 VSUBS 0.033425f
C1060 VN.n19 VSUBS 0.045684f
C1061 VN.n20 VSUBS 0.024635f
C1062 VN.n21 VSUBS 0.024635f
C1063 VN.n22 VSUBS 0.024635f
C1064 VN.n23 VSUBS 1.03874f
C1065 VN.n24 VSUBS 0.045684f
C1066 VN.n25 VSUBS 0.045684f
C1067 VN.n26 VSUBS 0.024635f
C1068 VN.n27 VSUBS 0.024635f
C1069 VN.n28 VSUBS 0.024635f
C1070 VN.n29 VSUBS 0.038197f
C1071 VN.n30 VSUBS 0.045684f
C1072 VN.n31 VSUBS 0.042526f
C1073 VN.n32 VSUBS 0.024635f
C1074 VN.n33 VSUBS 0.024635f
C1075 VN.n34 VSUBS 0.026288f
C1076 VN.n35 VSUBS 0.045684f
C1077 VN.n36 VSUBS 0.047199f
C1078 VN.n37 VSUBS 0.024635f
C1079 VN.n38 VSUBS 0.024635f
C1080 VN.n39 VSUBS 0.024635f
C1081 VN.n40 VSUBS 0.042708f
C1082 VN.n41 VSUBS 0.045684f
C1083 VN.n42 VSUBS 0.039369f
C1084 VN.n43 VSUBS 0.039754f
C1085 VN.n44 VSUBS 0.054659f
C1086 VN.t8 VSUBS 2.90784f
C1087 VN.n45 VSUBS 1.11119f
C1088 VN.n46 VSUBS 0.024635f
C1089 VN.n47 VSUBS 0.027399f
C1090 VN.n48 VSUBS 0.024635f
C1091 VN.t5 VSUBS 2.90784f
C1092 VN.n49 VSUBS 1.01561f
C1093 VN.n50 VSUBS 0.024635f
C1094 VN.n51 VSUBS 0.033425f
C1095 VN.n52 VSUBS 0.024635f
C1096 VN.t3 VSUBS 2.90784f
C1097 VN.n53 VSUBS 0.045684f
C1098 VN.n54 VSUBS 0.024635f
C1099 VN.n55 VSUBS 0.045684f
C1100 VN.t2 VSUBS 3.1877f
C1101 VN.n56 VSUBS 1.05131f
C1102 VN.t9 VSUBS 2.90784f
C1103 VN.n57 VSUBS 1.10342f
C1104 VN.n58 VSUBS 0.042526f
C1105 VN.n59 VSUBS 0.282061f
C1106 VN.n60 VSUBS 0.024635f
C1107 VN.n61 VSUBS 0.024635f
C1108 VN.n62 VSUBS 0.038197f
C1109 VN.n63 VSUBS 0.033425f
C1110 VN.n64 VSUBS 0.045684f
C1111 VN.n65 VSUBS 0.024635f
C1112 VN.n66 VSUBS 0.024635f
C1113 VN.n67 VSUBS 0.024635f
C1114 VN.n68 VSUBS 1.03874f
C1115 VN.n69 VSUBS 0.045684f
C1116 VN.n70 VSUBS 0.045684f
C1117 VN.n71 VSUBS 0.024635f
C1118 VN.n72 VSUBS 0.024635f
C1119 VN.n73 VSUBS 0.024635f
C1120 VN.n74 VSUBS 0.038197f
C1121 VN.n75 VSUBS 0.045684f
C1122 VN.n76 VSUBS 0.042526f
C1123 VN.n77 VSUBS 0.024635f
C1124 VN.n78 VSUBS 0.024635f
C1125 VN.n79 VSUBS 0.026288f
C1126 VN.n80 VSUBS 0.045684f
C1127 VN.n81 VSUBS 0.047199f
C1128 VN.n82 VSUBS 0.024635f
C1129 VN.n83 VSUBS 0.024635f
C1130 VN.n84 VSUBS 0.024635f
C1131 VN.n85 VSUBS 0.042708f
C1132 VN.n86 VSUBS 0.045684f
C1133 VN.n87 VSUBS 0.039369f
C1134 VN.n88 VSUBS 0.039754f
C1135 VN.n89 VSUBS 1.70325f
C1136 VDD1.t9 VSUBS 3.45142f
C1137 VDD1.t5 VSUBS 0.327924f
C1138 VDD1.t3 VSUBS 0.327924f
C1139 VDD1.n0 VSUBS 2.62003f
C1140 VDD1.n1 VSUBS 1.87176f
C1141 VDD1.t0 VSUBS 3.45141f
C1142 VDD1.t7 VSUBS 0.327924f
C1143 VDD1.t4 VSUBS 0.327924f
C1144 VDD1.n2 VSUBS 2.62002f
C1145 VDD1.n3 VSUBS 1.86188f
C1146 VDD1.t1 VSUBS 0.327924f
C1147 VDD1.t2 VSUBS 0.327924f
C1148 VDD1.n4 VSUBS 2.65154f
C1149 VDD1.n5 VSUBS 4.40923f
C1150 VDD1.t8 VSUBS 0.327924f
C1151 VDD1.t6 VSUBS 0.327924f
C1152 VDD1.n6 VSUBS 2.62003f
C1153 VDD1.n7 VSUBS 4.53525f
C1154 VTAIL.t2 VSUBS 0.315779f
C1155 VTAIL.t6 VSUBS 0.315779f
C1156 VTAIL.n0 VSUBS 2.35723f
C1157 VTAIL.n1 VSUBS 1.07222f
C1158 VTAIL.t14 VSUBS 3.10077f
C1159 VTAIL.n2 VSUBS 1.25289f
C1160 VTAIL.t19 VSUBS 0.315779f
C1161 VTAIL.t15 VSUBS 0.315779f
C1162 VTAIL.n3 VSUBS 2.35723f
C1163 VTAIL.n4 VSUBS 1.22851f
C1164 VTAIL.t16 VSUBS 0.315779f
C1165 VTAIL.t18 VSUBS 0.315779f
C1166 VTAIL.n5 VSUBS 2.35723f
C1167 VTAIL.n6 VSUBS 3.00199f
C1168 VTAIL.t0 VSUBS 0.315779f
C1169 VTAIL.t7 VSUBS 0.315779f
C1170 VTAIL.n7 VSUBS 2.35724f
C1171 VTAIL.n8 VSUBS 3.00199f
C1172 VTAIL.t9 VSUBS 0.315779f
C1173 VTAIL.t1 VSUBS 0.315779f
C1174 VTAIL.n9 VSUBS 2.35724f
C1175 VTAIL.n10 VSUBS 1.22851f
C1176 VTAIL.t5 VSUBS 3.10079f
C1177 VTAIL.n11 VSUBS 1.25287f
C1178 VTAIL.t11 VSUBS 0.315779f
C1179 VTAIL.t17 VSUBS 0.315779f
C1180 VTAIL.n12 VSUBS 2.35724f
C1181 VTAIL.n13 VSUBS 1.13521f
C1182 VTAIL.t13 VSUBS 0.315779f
C1183 VTAIL.t12 VSUBS 0.315779f
C1184 VTAIL.n14 VSUBS 2.35724f
C1185 VTAIL.n15 VSUBS 1.22851f
C1186 VTAIL.t10 VSUBS 3.10079f
C1187 VTAIL.n16 VSUBS 2.84614f
C1188 VTAIL.t4 VSUBS 3.10077f
C1189 VTAIL.n17 VSUBS 2.84616f
C1190 VTAIL.t8 VSUBS 0.315779f
C1191 VTAIL.t3 VSUBS 0.315779f
C1192 VTAIL.n18 VSUBS 2.35723f
C1193 VTAIL.n19 VSUBS 1.01799f
C1194 VP.t7 VSUBS 3.14006f
C1195 VP.n0 VSUBS 1.19993f
C1196 VP.n1 VSUBS 0.026603f
C1197 VP.n2 VSUBS 0.029587f
C1198 VP.n3 VSUBS 0.026603f
C1199 VP.t8 VSUBS 3.14006f
C1200 VP.n4 VSUBS 1.09672f
C1201 VP.n5 VSUBS 0.026603f
C1202 VP.n6 VSUBS 0.036095f
C1203 VP.n7 VSUBS 0.026603f
C1204 VP.t5 VSUBS 3.14006f
C1205 VP.n8 VSUBS 0.049332f
C1206 VP.n9 VSUBS 0.026603f
C1207 VP.n10 VSUBS 0.049332f
C1208 VP.n11 VSUBS 0.026603f
C1209 VP.t2 VSUBS 3.14006f
C1210 VP.n12 VSUBS 0.050968f
C1211 VP.n13 VSUBS 0.026603f
C1212 VP.n14 VSUBS 0.042513f
C1213 VP.t3 VSUBS 3.14006f
C1214 VP.n15 VSUBS 1.19993f
C1215 VP.n16 VSUBS 0.026603f
C1216 VP.n17 VSUBS 0.029587f
C1217 VP.n18 VSUBS 0.026603f
C1218 VP.t1 VSUBS 3.14006f
C1219 VP.n19 VSUBS 1.09672f
C1220 VP.n20 VSUBS 0.026603f
C1221 VP.n21 VSUBS 0.036095f
C1222 VP.n22 VSUBS 0.026603f
C1223 VP.t6 VSUBS 3.14006f
C1224 VP.n23 VSUBS 0.049332f
C1225 VP.n24 VSUBS 0.026603f
C1226 VP.n25 VSUBS 0.049332f
C1227 VP.t0 VSUBS 3.44227f
C1228 VP.n26 VSUBS 1.13527f
C1229 VP.t4 VSUBS 3.14006f
C1230 VP.n27 VSUBS 1.19154f
C1231 VP.n28 VSUBS 0.045922f
C1232 VP.n29 VSUBS 0.304586f
C1233 VP.n30 VSUBS 0.026603f
C1234 VP.n31 VSUBS 0.026603f
C1235 VP.n32 VSUBS 0.041247f
C1236 VP.n33 VSUBS 0.036095f
C1237 VP.n34 VSUBS 0.049332f
C1238 VP.n35 VSUBS 0.026603f
C1239 VP.n36 VSUBS 0.026603f
C1240 VP.n37 VSUBS 0.026603f
C1241 VP.n38 VSUBS 1.1217f
C1242 VP.n39 VSUBS 0.049332f
C1243 VP.n40 VSUBS 0.049332f
C1244 VP.n41 VSUBS 0.026603f
C1245 VP.n42 VSUBS 0.026603f
C1246 VP.n43 VSUBS 0.026603f
C1247 VP.n44 VSUBS 0.041247f
C1248 VP.n45 VSUBS 0.049332f
C1249 VP.n46 VSUBS 0.045922f
C1250 VP.n47 VSUBS 0.026603f
C1251 VP.n48 VSUBS 0.026603f
C1252 VP.n49 VSUBS 0.028388f
C1253 VP.n50 VSUBS 0.049332f
C1254 VP.n51 VSUBS 0.050968f
C1255 VP.n52 VSUBS 0.026603f
C1256 VP.n53 VSUBS 0.026603f
C1257 VP.n54 VSUBS 0.026603f
C1258 VP.n55 VSUBS 0.046118f
C1259 VP.n56 VSUBS 0.049332f
C1260 VP.n57 VSUBS 0.042513f
C1261 VP.n58 VSUBS 0.042929f
C1262 VP.n59 VSUBS 1.82887f
C1263 VP.t9 VSUBS 3.14006f
C1264 VP.n60 VSUBS 1.19993f
C1265 VP.n61 VSUBS 1.84558f
C1266 VP.n62 VSUBS 0.042929f
C1267 VP.n63 VSUBS 0.026603f
C1268 VP.n64 VSUBS 0.049332f
C1269 VP.n65 VSUBS 0.046118f
C1270 VP.n66 VSUBS 0.029587f
C1271 VP.n67 VSUBS 0.026603f
C1272 VP.n68 VSUBS 0.026603f
C1273 VP.n69 VSUBS 0.026603f
C1274 VP.n70 VSUBS 0.049332f
C1275 VP.n71 VSUBS 0.028388f
C1276 VP.n72 VSUBS 1.09672f
C1277 VP.n73 VSUBS 0.045922f
C1278 VP.n74 VSUBS 0.026603f
C1279 VP.n75 VSUBS 0.026603f
C1280 VP.n76 VSUBS 0.026603f
C1281 VP.n77 VSUBS 0.041247f
C1282 VP.n78 VSUBS 0.036095f
C1283 VP.n79 VSUBS 0.049332f
C1284 VP.n80 VSUBS 0.026603f
C1285 VP.n81 VSUBS 0.026603f
C1286 VP.n82 VSUBS 0.026603f
C1287 VP.n83 VSUBS 1.1217f
C1288 VP.n84 VSUBS 0.049332f
C1289 VP.n85 VSUBS 0.049332f
C1290 VP.n86 VSUBS 0.026603f
C1291 VP.n87 VSUBS 0.026603f
C1292 VP.n88 VSUBS 0.026603f
C1293 VP.n89 VSUBS 0.041247f
C1294 VP.n90 VSUBS 0.049332f
C1295 VP.n91 VSUBS 0.045922f
C1296 VP.n92 VSUBS 0.026603f
C1297 VP.n93 VSUBS 0.026603f
C1298 VP.n94 VSUBS 0.028388f
C1299 VP.n95 VSUBS 0.049332f
C1300 VP.n96 VSUBS 0.050968f
C1301 VP.n97 VSUBS 0.026603f
C1302 VP.n98 VSUBS 0.026603f
C1303 VP.n99 VSUBS 0.026603f
C1304 VP.n100 VSUBS 0.046118f
C1305 VP.n101 VSUBS 0.049332f
C1306 VP.n102 VSUBS 0.042513f
C1307 VP.n103 VSUBS 0.042929f
C1308 VP.n104 VSUBS 0.059024f
.ends

