* NGSPICE file created from diff_pair_sample_1004.ext - technology: sky130A

.subckt diff_pair_sample_1004 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X1 VDD2.t8 VN.t1 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=1.7655 ps=11.03 w=10.7 l=2.74
X2 VTAIL.t1 VP.t0 VDD1.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X3 B.t22 B.t20 B.t21 B.t14 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=2.74
X4 VTAIL.t5 VP.t1 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X5 VTAIL.t18 VN.t2 VDD2.t7 B.t23 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X6 VDD1.t7 VP.t2 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=4.173 ps=22.18 w=10.7 l=2.74
X7 VTAIL.t19 VP.t3 VDD1.t6 B.t23 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X8 B.t19 B.t17 B.t18 B.t10 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=2.74
X9 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=1.7655 ps=11.03 w=10.7 l=2.74
X10 VDD2.t6 VN.t3 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=4.173 ps=22.18 w=10.7 l=2.74
X11 VTAIL.t9 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X12 VDD2.t4 VN.t5 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=4.173 ps=22.18 w=10.7 l=2.74
X13 VDD1.t4 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=4.173 ps=22.18 w=10.7 l=2.74
X14 VTAIL.t11 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X15 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=2.74
X16 VDD2.t2 VN.t7 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=1.7655 ps=11.03 w=10.7 l=2.74
X17 VDD1.t3 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=1.7655 ps=11.03 w=10.7 l=2.74
X18 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=2.74
X19 VTAIL.t13 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X20 VDD1.t2 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X21 VDD2.t0 VN.t9 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X22 VDD1.t1 VP.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
X23 VTAIL.t3 VP.t9 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7655 pd=11.03 as=1.7655 ps=11.03 w=10.7 l=2.74
R0 VN.n83 VN.n43 161.3
R1 VN.n82 VN.n81 161.3
R2 VN.n80 VN.n44 161.3
R3 VN.n79 VN.n78 161.3
R4 VN.n77 VN.n45 161.3
R5 VN.n76 VN.n75 161.3
R6 VN.n74 VN.n73 161.3
R7 VN.n72 VN.n47 161.3
R8 VN.n71 VN.n70 161.3
R9 VN.n69 VN.n48 161.3
R10 VN.n68 VN.n67 161.3
R11 VN.n66 VN.n49 161.3
R12 VN.n65 VN.n64 161.3
R13 VN.n63 VN.n50 161.3
R14 VN.n62 VN.n61 161.3
R15 VN.n60 VN.n51 161.3
R16 VN.n59 VN.n58 161.3
R17 VN.n57 VN.n52 161.3
R18 VN.n56 VN.n55 161.3
R19 VN.n40 VN.n0 161.3
R20 VN.n39 VN.n38 161.3
R21 VN.n37 VN.n1 161.3
R22 VN.n36 VN.n35 161.3
R23 VN.n34 VN.n2 161.3
R24 VN.n33 VN.n32 161.3
R25 VN.n31 VN.n30 161.3
R26 VN.n29 VN.n4 161.3
R27 VN.n28 VN.n27 161.3
R28 VN.n26 VN.n5 161.3
R29 VN.n25 VN.n24 161.3
R30 VN.n23 VN.n6 161.3
R31 VN.n22 VN.n21 161.3
R32 VN.n20 VN.n7 161.3
R33 VN.n19 VN.n18 161.3
R34 VN.n17 VN.n8 161.3
R35 VN.n16 VN.n15 161.3
R36 VN.n14 VN.n9 161.3
R37 VN.n13 VN.n12 161.3
R38 VN.n10 VN.t7 126.767
R39 VN.n53 VN.t5 126.767
R40 VN.n42 VN.n41 104.022
R41 VN.n85 VN.n84 104.022
R42 VN.n22 VN.t9 94.1136
R43 VN.n11 VN.t8 94.1136
R44 VN.n3 VN.t4 94.1136
R45 VN.n41 VN.t3 94.1136
R46 VN.n65 VN.t0 94.1136
R47 VN.n54 VN.t2 94.1136
R48 VN.n46 VN.t6 94.1136
R49 VN.n84 VN.t1 94.1136
R50 VN.n11 VN.n10 69.6937
R51 VN.n54 VN.n53 69.6937
R52 VN VN.n85 53.1762
R53 VN.n35 VN.n1 50.7491
R54 VN.n78 VN.n44 50.7491
R55 VN.n17 VN.n16 43.9677
R56 VN.n28 VN.n5 43.9677
R57 VN.n60 VN.n59 43.9677
R58 VN.n71 VN.n48 43.9677
R59 VN.n18 VN.n17 37.1863
R60 VN.n24 VN.n5 37.1863
R61 VN.n61 VN.n60 37.1863
R62 VN.n67 VN.n48 37.1863
R63 VN.n35 VN.n34 30.405
R64 VN.n78 VN.n77 30.405
R65 VN.n12 VN.n9 24.5923
R66 VN.n16 VN.n9 24.5923
R67 VN.n18 VN.n7 24.5923
R68 VN.n22 VN.n7 24.5923
R69 VN.n23 VN.n22 24.5923
R70 VN.n24 VN.n23 24.5923
R71 VN.n29 VN.n28 24.5923
R72 VN.n30 VN.n29 24.5923
R73 VN.n34 VN.n33 24.5923
R74 VN.n39 VN.n1 24.5923
R75 VN.n40 VN.n39 24.5923
R76 VN.n59 VN.n52 24.5923
R77 VN.n55 VN.n52 24.5923
R78 VN.n67 VN.n66 24.5923
R79 VN.n66 VN.n65 24.5923
R80 VN.n65 VN.n50 24.5923
R81 VN.n61 VN.n50 24.5923
R82 VN.n77 VN.n76 24.5923
R83 VN.n73 VN.n72 24.5923
R84 VN.n72 VN.n71 24.5923
R85 VN.n83 VN.n82 24.5923
R86 VN.n82 VN.n44 24.5923
R87 VN.n33 VN.n3 21.1495
R88 VN.n76 VN.n46 21.1495
R89 VN.n56 VN.n53 7.0306
R90 VN.n13 VN.n10 7.0306
R91 VN.n41 VN.n40 6.88621
R92 VN.n84 VN.n83 6.88621
R93 VN.n12 VN.n11 3.44336
R94 VN.n30 VN.n3 3.44336
R95 VN.n55 VN.n54 3.44336
R96 VN.n73 VN.n46 3.44336
R97 VN.n85 VN.n43 0.278335
R98 VN.n42 VN.n0 0.278335
R99 VN.n81 VN.n43 0.189894
R100 VN.n81 VN.n80 0.189894
R101 VN.n80 VN.n79 0.189894
R102 VN.n79 VN.n45 0.189894
R103 VN.n75 VN.n45 0.189894
R104 VN.n75 VN.n74 0.189894
R105 VN.n74 VN.n47 0.189894
R106 VN.n70 VN.n47 0.189894
R107 VN.n70 VN.n69 0.189894
R108 VN.n69 VN.n68 0.189894
R109 VN.n68 VN.n49 0.189894
R110 VN.n64 VN.n49 0.189894
R111 VN.n64 VN.n63 0.189894
R112 VN.n63 VN.n62 0.189894
R113 VN.n62 VN.n51 0.189894
R114 VN.n58 VN.n51 0.189894
R115 VN.n58 VN.n57 0.189894
R116 VN.n57 VN.n56 0.189894
R117 VN.n14 VN.n13 0.189894
R118 VN.n15 VN.n14 0.189894
R119 VN.n15 VN.n8 0.189894
R120 VN.n19 VN.n8 0.189894
R121 VN.n20 VN.n19 0.189894
R122 VN.n21 VN.n20 0.189894
R123 VN.n21 VN.n6 0.189894
R124 VN.n25 VN.n6 0.189894
R125 VN.n26 VN.n25 0.189894
R126 VN.n27 VN.n26 0.189894
R127 VN.n27 VN.n4 0.189894
R128 VN.n31 VN.n4 0.189894
R129 VN.n32 VN.n31 0.189894
R130 VN.n32 VN.n2 0.189894
R131 VN.n36 VN.n2 0.189894
R132 VN.n37 VN.n36 0.189894
R133 VN.n38 VN.n37 0.189894
R134 VN.n38 VN.n0 0.189894
R135 VN VN.n42 0.153485
R136 VTAIL.n240 VTAIL.n188 289.615
R137 VTAIL.n54 VTAIL.n2 289.615
R138 VTAIL.n182 VTAIL.n130 289.615
R139 VTAIL.n120 VTAIL.n68 289.615
R140 VTAIL.n207 VTAIL.n206 185
R141 VTAIL.n204 VTAIL.n203 185
R142 VTAIL.n213 VTAIL.n212 185
R143 VTAIL.n215 VTAIL.n214 185
R144 VTAIL.n200 VTAIL.n199 185
R145 VTAIL.n221 VTAIL.n220 185
R146 VTAIL.n224 VTAIL.n223 185
R147 VTAIL.n222 VTAIL.n196 185
R148 VTAIL.n229 VTAIL.n195 185
R149 VTAIL.n231 VTAIL.n230 185
R150 VTAIL.n233 VTAIL.n232 185
R151 VTAIL.n192 VTAIL.n191 185
R152 VTAIL.n239 VTAIL.n238 185
R153 VTAIL.n241 VTAIL.n240 185
R154 VTAIL.n21 VTAIL.n20 185
R155 VTAIL.n18 VTAIL.n17 185
R156 VTAIL.n27 VTAIL.n26 185
R157 VTAIL.n29 VTAIL.n28 185
R158 VTAIL.n14 VTAIL.n13 185
R159 VTAIL.n35 VTAIL.n34 185
R160 VTAIL.n38 VTAIL.n37 185
R161 VTAIL.n36 VTAIL.n10 185
R162 VTAIL.n43 VTAIL.n9 185
R163 VTAIL.n45 VTAIL.n44 185
R164 VTAIL.n47 VTAIL.n46 185
R165 VTAIL.n6 VTAIL.n5 185
R166 VTAIL.n53 VTAIL.n52 185
R167 VTAIL.n55 VTAIL.n54 185
R168 VTAIL.n183 VTAIL.n182 185
R169 VTAIL.n181 VTAIL.n180 185
R170 VTAIL.n134 VTAIL.n133 185
R171 VTAIL.n175 VTAIL.n174 185
R172 VTAIL.n173 VTAIL.n172 185
R173 VTAIL.n171 VTAIL.n137 185
R174 VTAIL.n141 VTAIL.n138 185
R175 VTAIL.n166 VTAIL.n165 185
R176 VTAIL.n164 VTAIL.n163 185
R177 VTAIL.n143 VTAIL.n142 185
R178 VTAIL.n158 VTAIL.n157 185
R179 VTAIL.n156 VTAIL.n155 185
R180 VTAIL.n147 VTAIL.n146 185
R181 VTAIL.n150 VTAIL.n149 185
R182 VTAIL.n121 VTAIL.n120 185
R183 VTAIL.n119 VTAIL.n118 185
R184 VTAIL.n72 VTAIL.n71 185
R185 VTAIL.n113 VTAIL.n112 185
R186 VTAIL.n111 VTAIL.n110 185
R187 VTAIL.n109 VTAIL.n75 185
R188 VTAIL.n79 VTAIL.n76 185
R189 VTAIL.n104 VTAIL.n103 185
R190 VTAIL.n102 VTAIL.n101 185
R191 VTAIL.n81 VTAIL.n80 185
R192 VTAIL.n96 VTAIL.n95 185
R193 VTAIL.n94 VTAIL.n93 185
R194 VTAIL.n85 VTAIL.n84 185
R195 VTAIL.n88 VTAIL.n87 185
R196 VTAIL.t14 VTAIL.n205 149.524
R197 VTAIL.t8 VTAIL.n19 149.524
R198 VTAIL.t0 VTAIL.n148 149.524
R199 VTAIL.t16 VTAIL.n86 149.524
R200 VTAIL.n206 VTAIL.n203 104.615
R201 VTAIL.n213 VTAIL.n203 104.615
R202 VTAIL.n214 VTAIL.n213 104.615
R203 VTAIL.n214 VTAIL.n199 104.615
R204 VTAIL.n221 VTAIL.n199 104.615
R205 VTAIL.n223 VTAIL.n221 104.615
R206 VTAIL.n223 VTAIL.n222 104.615
R207 VTAIL.n222 VTAIL.n195 104.615
R208 VTAIL.n231 VTAIL.n195 104.615
R209 VTAIL.n232 VTAIL.n231 104.615
R210 VTAIL.n232 VTAIL.n191 104.615
R211 VTAIL.n239 VTAIL.n191 104.615
R212 VTAIL.n240 VTAIL.n239 104.615
R213 VTAIL.n20 VTAIL.n17 104.615
R214 VTAIL.n27 VTAIL.n17 104.615
R215 VTAIL.n28 VTAIL.n27 104.615
R216 VTAIL.n28 VTAIL.n13 104.615
R217 VTAIL.n35 VTAIL.n13 104.615
R218 VTAIL.n37 VTAIL.n35 104.615
R219 VTAIL.n37 VTAIL.n36 104.615
R220 VTAIL.n36 VTAIL.n9 104.615
R221 VTAIL.n45 VTAIL.n9 104.615
R222 VTAIL.n46 VTAIL.n45 104.615
R223 VTAIL.n46 VTAIL.n5 104.615
R224 VTAIL.n53 VTAIL.n5 104.615
R225 VTAIL.n54 VTAIL.n53 104.615
R226 VTAIL.n182 VTAIL.n181 104.615
R227 VTAIL.n181 VTAIL.n133 104.615
R228 VTAIL.n174 VTAIL.n133 104.615
R229 VTAIL.n174 VTAIL.n173 104.615
R230 VTAIL.n173 VTAIL.n137 104.615
R231 VTAIL.n141 VTAIL.n137 104.615
R232 VTAIL.n165 VTAIL.n141 104.615
R233 VTAIL.n165 VTAIL.n164 104.615
R234 VTAIL.n164 VTAIL.n142 104.615
R235 VTAIL.n157 VTAIL.n142 104.615
R236 VTAIL.n157 VTAIL.n156 104.615
R237 VTAIL.n156 VTAIL.n146 104.615
R238 VTAIL.n149 VTAIL.n146 104.615
R239 VTAIL.n120 VTAIL.n119 104.615
R240 VTAIL.n119 VTAIL.n71 104.615
R241 VTAIL.n112 VTAIL.n71 104.615
R242 VTAIL.n112 VTAIL.n111 104.615
R243 VTAIL.n111 VTAIL.n75 104.615
R244 VTAIL.n79 VTAIL.n75 104.615
R245 VTAIL.n103 VTAIL.n79 104.615
R246 VTAIL.n103 VTAIL.n102 104.615
R247 VTAIL.n102 VTAIL.n80 104.615
R248 VTAIL.n95 VTAIL.n80 104.615
R249 VTAIL.n95 VTAIL.n94 104.615
R250 VTAIL.n94 VTAIL.n84 104.615
R251 VTAIL.n87 VTAIL.n84 104.615
R252 VTAIL.n206 VTAIL.t14 52.3082
R253 VTAIL.n20 VTAIL.t8 52.3082
R254 VTAIL.n149 VTAIL.t0 52.3082
R255 VTAIL.n87 VTAIL.t16 52.3082
R256 VTAIL.n129 VTAIL.n128 46.0494
R257 VTAIL.n127 VTAIL.n126 46.0494
R258 VTAIL.n67 VTAIL.n66 46.0494
R259 VTAIL.n65 VTAIL.n64 46.0494
R260 VTAIL.n247 VTAIL.n246 46.0492
R261 VTAIL.n1 VTAIL.n0 46.0492
R262 VTAIL.n61 VTAIL.n60 46.0492
R263 VTAIL.n63 VTAIL.n62 46.0492
R264 VTAIL.n245 VTAIL.n244 32.5732
R265 VTAIL.n59 VTAIL.n58 32.5732
R266 VTAIL.n187 VTAIL.n186 32.5732
R267 VTAIL.n125 VTAIL.n124 32.5732
R268 VTAIL.n65 VTAIL.n63 26.8841
R269 VTAIL.n245 VTAIL.n187 24.2376
R270 VTAIL.n230 VTAIL.n229 13.1884
R271 VTAIL.n44 VTAIL.n43 13.1884
R272 VTAIL.n172 VTAIL.n171 13.1884
R273 VTAIL.n110 VTAIL.n109 13.1884
R274 VTAIL.n228 VTAIL.n196 12.8005
R275 VTAIL.n233 VTAIL.n194 12.8005
R276 VTAIL.n42 VTAIL.n10 12.8005
R277 VTAIL.n47 VTAIL.n8 12.8005
R278 VTAIL.n175 VTAIL.n136 12.8005
R279 VTAIL.n170 VTAIL.n138 12.8005
R280 VTAIL.n113 VTAIL.n74 12.8005
R281 VTAIL.n108 VTAIL.n76 12.8005
R282 VTAIL.n225 VTAIL.n224 12.0247
R283 VTAIL.n234 VTAIL.n192 12.0247
R284 VTAIL.n39 VTAIL.n38 12.0247
R285 VTAIL.n48 VTAIL.n6 12.0247
R286 VTAIL.n176 VTAIL.n134 12.0247
R287 VTAIL.n167 VTAIL.n166 12.0247
R288 VTAIL.n114 VTAIL.n72 12.0247
R289 VTAIL.n105 VTAIL.n104 12.0247
R290 VTAIL.n220 VTAIL.n198 11.249
R291 VTAIL.n238 VTAIL.n237 11.249
R292 VTAIL.n34 VTAIL.n12 11.249
R293 VTAIL.n52 VTAIL.n51 11.249
R294 VTAIL.n180 VTAIL.n179 11.249
R295 VTAIL.n163 VTAIL.n140 11.249
R296 VTAIL.n118 VTAIL.n117 11.249
R297 VTAIL.n101 VTAIL.n78 11.249
R298 VTAIL.n219 VTAIL.n200 10.4732
R299 VTAIL.n241 VTAIL.n190 10.4732
R300 VTAIL.n33 VTAIL.n14 10.4732
R301 VTAIL.n55 VTAIL.n4 10.4732
R302 VTAIL.n183 VTAIL.n132 10.4732
R303 VTAIL.n162 VTAIL.n143 10.4732
R304 VTAIL.n121 VTAIL.n70 10.4732
R305 VTAIL.n100 VTAIL.n81 10.4732
R306 VTAIL.n207 VTAIL.n205 10.2747
R307 VTAIL.n21 VTAIL.n19 10.2747
R308 VTAIL.n150 VTAIL.n148 10.2747
R309 VTAIL.n88 VTAIL.n86 10.2747
R310 VTAIL.n216 VTAIL.n215 9.69747
R311 VTAIL.n242 VTAIL.n188 9.69747
R312 VTAIL.n30 VTAIL.n29 9.69747
R313 VTAIL.n56 VTAIL.n2 9.69747
R314 VTAIL.n184 VTAIL.n130 9.69747
R315 VTAIL.n159 VTAIL.n158 9.69747
R316 VTAIL.n122 VTAIL.n68 9.69747
R317 VTAIL.n97 VTAIL.n96 9.69747
R318 VTAIL.n244 VTAIL.n243 9.45567
R319 VTAIL.n58 VTAIL.n57 9.45567
R320 VTAIL.n186 VTAIL.n185 9.45567
R321 VTAIL.n124 VTAIL.n123 9.45567
R322 VTAIL.n243 VTAIL.n242 9.3005
R323 VTAIL.n190 VTAIL.n189 9.3005
R324 VTAIL.n237 VTAIL.n236 9.3005
R325 VTAIL.n235 VTAIL.n234 9.3005
R326 VTAIL.n194 VTAIL.n193 9.3005
R327 VTAIL.n209 VTAIL.n208 9.3005
R328 VTAIL.n211 VTAIL.n210 9.3005
R329 VTAIL.n202 VTAIL.n201 9.3005
R330 VTAIL.n217 VTAIL.n216 9.3005
R331 VTAIL.n219 VTAIL.n218 9.3005
R332 VTAIL.n198 VTAIL.n197 9.3005
R333 VTAIL.n226 VTAIL.n225 9.3005
R334 VTAIL.n228 VTAIL.n227 9.3005
R335 VTAIL.n57 VTAIL.n56 9.3005
R336 VTAIL.n4 VTAIL.n3 9.3005
R337 VTAIL.n51 VTAIL.n50 9.3005
R338 VTAIL.n49 VTAIL.n48 9.3005
R339 VTAIL.n8 VTAIL.n7 9.3005
R340 VTAIL.n23 VTAIL.n22 9.3005
R341 VTAIL.n25 VTAIL.n24 9.3005
R342 VTAIL.n16 VTAIL.n15 9.3005
R343 VTAIL.n31 VTAIL.n30 9.3005
R344 VTAIL.n33 VTAIL.n32 9.3005
R345 VTAIL.n12 VTAIL.n11 9.3005
R346 VTAIL.n40 VTAIL.n39 9.3005
R347 VTAIL.n42 VTAIL.n41 9.3005
R348 VTAIL.n152 VTAIL.n151 9.3005
R349 VTAIL.n154 VTAIL.n153 9.3005
R350 VTAIL.n145 VTAIL.n144 9.3005
R351 VTAIL.n160 VTAIL.n159 9.3005
R352 VTAIL.n162 VTAIL.n161 9.3005
R353 VTAIL.n140 VTAIL.n139 9.3005
R354 VTAIL.n168 VTAIL.n167 9.3005
R355 VTAIL.n170 VTAIL.n169 9.3005
R356 VTAIL.n185 VTAIL.n184 9.3005
R357 VTAIL.n132 VTAIL.n131 9.3005
R358 VTAIL.n179 VTAIL.n178 9.3005
R359 VTAIL.n177 VTAIL.n176 9.3005
R360 VTAIL.n136 VTAIL.n135 9.3005
R361 VTAIL.n90 VTAIL.n89 9.3005
R362 VTAIL.n92 VTAIL.n91 9.3005
R363 VTAIL.n83 VTAIL.n82 9.3005
R364 VTAIL.n98 VTAIL.n97 9.3005
R365 VTAIL.n100 VTAIL.n99 9.3005
R366 VTAIL.n78 VTAIL.n77 9.3005
R367 VTAIL.n106 VTAIL.n105 9.3005
R368 VTAIL.n108 VTAIL.n107 9.3005
R369 VTAIL.n123 VTAIL.n122 9.3005
R370 VTAIL.n70 VTAIL.n69 9.3005
R371 VTAIL.n117 VTAIL.n116 9.3005
R372 VTAIL.n115 VTAIL.n114 9.3005
R373 VTAIL.n74 VTAIL.n73 9.3005
R374 VTAIL.n212 VTAIL.n202 8.92171
R375 VTAIL.n26 VTAIL.n16 8.92171
R376 VTAIL.n155 VTAIL.n145 8.92171
R377 VTAIL.n93 VTAIL.n83 8.92171
R378 VTAIL.n211 VTAIL.n204 8.14595
R379 VTAIL.n25 VTAIL.n18 8.14595
R380 VTAIL.n154 VTAIL.n147 8.14595
R381 VTAIL.n92 VTAIL.n85 8.14595
R382 VTAIL.n208 VTAIL.n207 7.3702
R383 VTAIL.n22 VTAIL.n21 7.3702
R384 VTAIL.n151 VTAIL.n150 7.3702
R385 VTAIL.n89 VTAIL.n88 7.3702
R386 VTAIL.n208 VTAIL.n204 5.81868
R387 VTAIL.n22 VTAIL.n18 5.81868
R388 VTAIL.n151 VTAIL.n147 5.81868
R389 VTAIL.n89 VTAIL.n85 5.81868
R390 VTAIL.n212 VTAIL.n211 5.04292
R391 VTAIL.n26 VTAIL.n25 5.04292
R392 VTAIL.n155 VTAIL.n154 5.04292
R393 VTAIL.n93 VTAIL.n92 5.04292
R394 VTAIL.n215 VTAIL.n202 4.26717
R395 VTAIL.n244 VTAIL.n188 4.26717
R396 VTAIL.n29 VTAIL.n16 4.26717
R397 VTAIL.n58 VTAIL.n2 4.26717
R398 VTAIL.n186 VTAIL.n130 4.26717
R399 VTAIL.n158 VTAIL.n145 4.26717
R400 VTAIL.n124 VTAIL.n68 4.26717
R401 VTAIL.n96 VTAIL.n83 4.26717
R402 VTAIL.n216 VTAIL.n200 3.49141
R403 VTAIL.n242 VTAIL.n241 3.49141
R404 VTAIL.n30 VTAIL.n14 3.49141
R405 VTAIL.n56 VTAIL.n55 3.49141
R406 VTAIL.n184 VTAIL.n183 3.49141
R407 VTAIL.n159 VTAIL.n143 3.49141
R408 VTAIL.n122 VTAIL.n121 3.49141
R409 VTAIL.n97 VTAIL.n81 3.49141
R410 VTAIL.n209 VTAIL.n205 2.84303
R411 VTAIL.n23 VTAIL.n19 2.84303
R412 VTAIL.n152 VTAIL.n148 2.84303
R413 VTAIL.n90 VTAIL.n86 2.84303
R414 VTAIL.n220 VTAIL.n219 2.71565
R415 VTAIL.n238 VTAIL.n190 2.71565
R416 VTAIL.n34 VTAIL.n33 2.71565
R417 VTAIL.n52 VTAIL.n4 2.71565
R418 VTAIL.n180 VTAIL.n132 2.71565
R419 VTAIL.n163 VTAIL.n162 2.71565
R420 VTAIL.n118 VTAIL.n70 2.71565
R421 VTAIL.n101 VTAIL.n100 2.71565
R422 VTAIL.n67 VTAIL.n65 2.64705
R423 VTAIL.n125 VTAIL.n67 2.64705
R424 VTAIL.n129 VTAIL.n127 2.64705
R425 VTAIL.n187 VTAIL.n129 2.64705
R426 VTAIL.n63 VTAIL.n61 2.64705
R427 VTAIL.n61 VTAIL.n59 2.64705
R428 VTAIL.n247 VTAIL.n245 2.64705
R429 VTAIL VTAIL.n1 2.0436
R430 VTAIL.n224 VTAIL.n198 1.93989
R431 VTAIL.n237 VTAIL.n192 1.93989
R432 VTAIL.n38 VTAIL.n12 1.93989
R433 VTAIL.n51 VTAIL.n6 1.93989
R434 VTAIL.n179 VTAIL.n134 1.93989
R435 VTAIL.n166 VTAIL.n140 1.93989
R436 VTAIL.n117 VTAIL.n72 1.93989
R437 VTAIL.n104 VTAIL.n78 1.93989
R438 VTAIL.n246 VTAIL.t15 1.85097
R439 VTAIL.n246 VTAIL.t9 1.85097
R440 VTAIL.n0 VTAIL.t10 1.85097
R441 VTAIL.n0 VTAIL.t13 1.85097
R442 VTAIL.n60 VTAIL.t7 1.85097
R443 VTAIL.n60 VTAIL.t19 1.85097
R444 VTAIL.n62 VTAIL.t6 1.85097
R445 VTAIL.n62 VTAIL.t3 1.85097
R446 VTAIL.n128 VTAIL.t2 1.85097
R447 VTAIL.n128 VTAIL.t5 1.85097
R448 VTAIL.n126 VTAIL.t4 1.85097
R449 VTAIL.n126 VTAIL.t1 1.85097
R450 VTAIL.n66 VTAIL.t17 1.85097
R451 VTAIL.n66 VTAIL.t18 1.85097
R452 VTAIL.n64 VTAIL.t12 1.85097
R453 VTAIL.n64 VTAIL.t11 1.85097
R454 VTAIL.n127 VTAIL.n125 1.7936
R455 VTAIL.n59 VTAIL.n1 1.7936
R456 VTAIL.n225 VTAIL.n196 1.16414
R457 VTAIL.n234 VTAIL.n233 1.16414
R458 VTAIL.n39 VTAIL.n10 1.16414
R459 VTAIL.n48 VTAIL.n47 1.16414
R460 VTAIL.n176 VTAIL.n175 1.16414
R461 VTAIL.n167 VTAIL.n138 1.16414
R462 VTAIL.n114 VTAIL.n113 1.16414
R463 VTAIL.n105 VTAIL.n76 1.16414
R464 VTAIL VTAIL.n247 0.603948
R465 VTAIL.n229 VTAIL.n228 0.388379
R466 VTAIL.n230 VTAIL.n194 0.388379
R467 VTAIL.n43 VTAIL.n42 0.388379
R468 VTAIL.n44 VTAIL.n8 0.388379
R469 VTAIL.n172 VTAIL.n136 0.388379
R470 VTAIL.n171 VTAIL.n170 0.388379
R471 VTAIL.n110 VTAIL.n74 0.388379
R472 VTAIL.n109 VTAIL.n108 0.388379
R473 VTAIL.n210 VTAIL.n209 0.155672
R474 VTAIL.n210 VTAIL.n201 0.155672
R475 VTAIL.n217 VTAIL.n201 0.155672
R476 VTAIL.n218 VTAIL.n217 0.155672
R477 VTAIL.n218 VTAIL.n197 0.155672
R478 VTAIL.n226 VTAIL.n197 0.155672
R479 VTAIL.n227 VTAIL.n226 0.155672
R480 VTAIL.n227 VTAIL.n193 0.155672
R481 VTAIL.n235 VTAIL.n193 0.155672
R482 VTAIL.n236 VTAIL.n235 0.155672
R483 VTAIL.n236 VTAIL.n189 0.155672
R484 VTAIL.n243 VTAIL.n189 0.155672
R485 VTAIL.n24 VTAIL.n23 0.155672
R486 VTAIL.n24 VTAIL.n15 0.155672
R487 VTAIL.n31 VTAIL.n15 0.155672
R488 VTAIL.n32 VTAIL.n31 0.155672
R489 VTAIL.n32 VTAIL.n11 0.155672
R490 VTAIL.n40 VTAIL.n11 0.155672
R491 VTAIL.n41 VTAIL.n40 0.155672
R492 VTAIL.n41 VTAIL.n7 0.155672
R493 VTAIL.n49 VTAIL.n7 0.155672
R494 VTAIL.n50 VTAIL.n49 0.155672
R495 VTAIL.n50 VTAIL.n3 0.155672
R496 VTAIL.n57 VTAIL.n3 0.155672
R497 VTAIL.n185 VTAIL.n131 0.155672
R498 VTAIL.n178 VTAIL.n131 0.155672
R499 VTAIL.n178 VTAIL.n177 0.155672
R500 VTAIL.n177 VTAIL.n135 0.155672
R501 VTAIL.n169 VTAIL.n135 0.155672
R502 VTAIL.n169 VTAIL.n168 0.155672
R503 VTAIL.n168 VTAIL.n139 0.155672
R504 VTAIL.n161 VTAIL.n139 0.155672
R505 VTAIL.n161 VTAIL.n160 0.155672
R506 VTAIL.n160 VTAIL.n144 0.155672
R507 VTAIL.n153 VTAIL.n144 0.155672
R508 VTAIL.n153 VTAIL.n152 0.155672
R509 VTAIL.n123 VTAIL.n69 0.155672
R510 VTAIL.n116 VTAIL.n69 0.155672
R511 VTAIL.n116 VTAIL.n115 0.155672
R512 VTAIL.n115 VTAIL.n73 0.155672
R513 VTAIL.n107 VTAIL.n73 0.155672
R514 VTAIL.n107 VTAIL.n106 0.155672
R515 VTAIL.n106 VTAIL.n77 0.155672
R516 VTAIL.n99 VTAIL.n77 0.155672
R517 VTAIL.n99 VTAIL.n98 0.155672
R518 VTAIL.n98 VTAIL.n82 0.155672
R519 VTAIL.n91 VTAIL.n82 0.155672
R520 VTAIL.n91 VTAIL.n90 0.155672
R521 VDD2.n113 VDD2.n61 289.615
R522 VDD2.n52 VDD2.n0 289.615
R523 VDD2.n114 VDD2.n113 185
R524 VDD2.n112 VDD2.n111 185
R525 VDD2.n65 VDD2.n64 185
R526 VDD2.n106 VDD2.n105 185
R527 VDD2.n104 VDD2.n103 185
R528 VDD2.n102 VDD2.n68 185
R529 VDD2.n72 VDD2.n69 185
R530 VDD2.n97 VDD2.n96 185
R531 VDD2.n95 VDD2.n94 185
R532 VDD2.n74 VDD2.n73 185
R533 VDD2.n89 VDD2.n88 185
R534 VDD2.n87 VDD2.n86 185
R535 VDD2.n78 VDD2.n77 185
R536 VDD2.n81 VDD2.n80 185
R537 VDD2.n19 VDD2.n18 185
R538 VDD2.n16 VDD2.n15 185
R539 VDD2.n25 VDD2.n24 185
R540 VDD2.n27 VDD2.n26 185
R541 VDD2.n12 VDD2.n11 185
R542 VDD2.n33 VDD2.n32 185
R543 VDD2.n36 VDD2.n35 185
R544 VDD2.n34 VDD2.n8 185
R545 VDD2.n41 VDD2.n7 185
R546 VDD2.n43 VDD2.n42 185
R547 VDD2.n45 VDD2.n44 185
R548 VDD2.n4 VDD2.n3 185
R549 VDD2.n51 VDD2.n50 185
R550 VDD2.n53 VDD2.n52 185
R551 VDD2.t8 VDD2.n79 149.524
R552 VDD2.t2 VDD2.n17 149.524
R553 VDD2.n113 VDD2.n112 104.615
R554 VDD2.n112 VDD2.n64 104.615
R555 VDD2.n105 VDD2.n64 104.615
R556 VDD2.n105 VDD2.n104 104.615
R557 VDD2.n104 VDD2.n68 104.615
R558 VDD2.n72 VDD2.n68 104.615
R559 VDD2.n96 VDD2.n72 104.615
R560 VDD2.n96 VDD2.n95 104.615
R561 VDD2.n95 VDD2.n73 104.615
R562 VDD2.n88 VDD2.n73 104.615
R563 VDD2.n88 VDD2.n87 104.615
R564 VDD2.n87 VDD2.n77 104.615
R565 VDD2.n80 VDD2.n77 104.615
R566 VDD2.n18 VDD2.n15 104.615
R567 VDD2.n25 VDD2.n15 104.615
R568 VDD2.n26 VDD2.n25 104.615
R569 VDD2.n26 VDD2.n11 104.615
R570 VDD2.n33 VDD2.n11 104.615
R571 VDD2.n35 VDD2.n33 104.615
R572 VDD2.n35 VDD2.n34 104.615
R573 VDD2.n34 VDD2.n7 104.615
R574 VDD2.n43 VDD2.n7 104.615
R575 VDD2.n44 VDD2.n43 104.615
R576 VDD2.n44 VDD2.n3 104.615
R577 VDD2.n51 VDD2.n3 104.615
R578 VDD2.n52 VDD2.n51 104.615
R579 VDD2.n60 VDD2.n59 64.6576
R580 VDD2 VDD2.n121 64.6547
R581 VDD2.n120 VDD2.n119 62.7282
R582 VDD2.n58 VDD2.n57 62.728
R583 VDD2.n80 VDD2.t8 52.3082
R584 VDD2.n18 VDD2.t2 52.3082
R585 VDD2.n58 VDD2.n56 51.8986
R586 VDD2.n118 VDD2.n117 49.252
R587 VDD2.n118 VDD2.n60 45.5106
R588 VDD2.n103 VDD2.n102 13.1884
R589 VDD2.n42 VDD2.n41 13.1884
R590 VDD2.n106 VDD2.n67 12.8005
R591 VDD2.n101 VDD2.n69 12.8005
R592 VDD2.n40 VDD2.n8 12.8005
R593 VDD2.n45 VDD2.n6 12.8005
R594 VDD2.n107 VDD2.n65 12.0247
R595 VDD2.n98 VDD2.n97 12.0247
R596 VDD2.n37 VDD2.n36 12.0247
R597 VDD2.n46 VDD2.n4 12.0247
R598 VDD2.n111 VDD2.n110 11.249
R599 VDD2.n94 VDD2.n71 11.249
R600 VDD2.n32 VDD2.n10 11.249
R601 VDD2.n50 VDD2.n49 11.249
R602 VDD2.n114 VDD2.n63 10.4732
R603 VDD2.n93 VDD2.n74 10.4732
R604 VDD2.n31 VDD2.n12 10.4732
R605 VDD2.n53 VDD2.n2 10.4732
R606 VDD2.n81 VDD2.n79 10.2747
R607 VDD2.n19 VDD2.n17 10.2747
R608 VDD2.n115 VDD2.n61 9.69747
R609 VDD2.n90 VDD2.n89 9.69747
R610 VDD2.n28 VDD2.n27 9.69747
R611 VDD2.n54 VDD2.n0 9.69747
R612 VDD2.n117 VDD2.n116 9.45567
R613 VDD2.n56 VDD2.n55 9.45567
R614 VDD2.n83 VDD2.n82 9.3005
R615 VDD2.n85 VDD2.n84 9.3005
R616 VDD2.n76 VDD2.n75 9.3005
R617 VDD2.n91 VDD2.n90 9.3005
R618 VDD2.n93 VDD2.n92 9.3005
R619 VDD2.n71 VDD2.n70 9.3005
R620 VDD2.n99 VDD2.n98 9.3005
R621 VDD2.n101 VDD2.n100 9.3005
R622 VDD2.n116 VDD2.n115 9.3005
R623 VDD2.n63 VDD2.n62 9.3005
R624 VDD2.n110 VDD2.n109 9.3005
R625 VDD2.n108 VDD2.n107 9.3005
R626 VDD2.n67 VDD2.n66 9.3005
R627 VDD2.n55 VDD2.n54 9.3005
R628 VDD2.n2 VDD2.n1 9.3005
R629 VDD2.n49 VDD2.n48 9.3005
R630 VDD2.n47 VDD2.n46 9.3005
R631 VDD2.n6 VDD2.n5 9.3005
R632 VDD2.n21 VDD2.n20 9.3005
R633 VDD2.n23 VDD2.n22 9.3005
R634 VDD2.n14 VDD2.n13 9.3005
R635 VDD2.n29 VDD2.n28 9.3005
R636 VDD2.n31 VDD2.n30 9.3005
R637 VDD2.n10 VDD2.n9 9.3005
R638 VDD2.n38 VDD2.n37 9.3005
R639 VDD2.n40 VDD2.n39 9.3005
R640 VDD2.n86 VDD2.n76 8.92171
R641 VDD2.n24 VDD2.n14 8.92171
R642 VDD2.n85 VDD2.n78 8.14595
R643 VDD2.n23 VDD2.n16 8.14595
R644 VDD2.n82 VDD2.n81 7.3702
R645 VDD2.n20 VDD2.n19 7.3702
R646 VDD2.n82 VDD2.n78 5.81868
R647 VDD2.n20 VDD2.n16 5.81868
R648 VDD2.n86 VDD2.n85 5.04292
R649 VDD2.n24 VDD2.n23 5.04292
R650 VDD2.n117 VDD2.n61 4.26717
R651 VDD2.n89 VDD2.n76 4.26717
R652 VDD2.n27 VDD2.n14 4.26717
R653 VDD2.n56 VDD2.n0 4.26717
R654 VDD2.n115 VDD2.n114 3.49141
R655 VDD2.n90 VDD2.n74 3.49141
R656 VDD2.n28 VDD2.n12 3.49141
R657 VDD2.n54 VDD2.n53 3.49141
R658 VDD2.n83 VDD2.n79 2.84303
R659 VDD2.n21 VDD2.n17 2.84303
R660 VDD2.n111 VDD2.n63 2.71565
R661 VDD2.n94 VDD2.n93 2.71565
R662 VDD2.n32 VDD2.n31 2.71565
R663 VDD2.n50 VDD2.n2 2.71565
R664 VDD2.n120 VDD2.n118 2.64705
R665 VDD2.n110 VDD2.n65 1.93989
R666 VDD2.n97 VDD2.n71 1.93989
R667 VDD2.n36 VDD2.n10 1.93989
R668 VDD2.n49 VDD2.n4 1.93989
R669 VDD2.n121 VDD2.t7 1.85097
R670 VDD2.n121 VDD2.t4 1.85097
R671 VDD2.n119 VDD2.t3 1.85097
R672 VDD2.n119 VDD2.t9 1.85097
R673 VDD2.n59 VDD2.t5 1.85097
R674 VDD2.n59 VDD2.t6 1.85097
R675 VDD2.n57 VDD2.t1 1.85097
R676 VDD2.n57 VDD2.t0 1.85097
R677 VDD2.n107 VDD2.n106 1.16414
R678 VDD2.n98 VDD2.n69 1.16414
R679 VDD2.n37 VDD2.n8 1.16414
R680 VDD2.n46 VDD2.n45 1.16414
R681 VDD2 VDD2.n120 0.720328
R682 VDD2.n60 VDD2.n58 0.606792
R683 VDD2.n103 VDD2.n67 0.388379
R684 VDD2.n102 VDD2.n101 0.388379
R685 VDD2.n41 VDD2.n40 0.388379
R686 VDD2.n42 VDD2.n6 0.388379
R687 VDD2.n116 VDD2.n62 0.155672
R688 VDD2.n109 VDD2.n62 0.155672
R689 VDD2.n109 VDD2.n108 0.155672
R690 VDD2.n108 VDD2.n66 0.155672
R691 VDD2.n100 VDD2.n66 0.155672
R692 VDD2.n100 VDD2.n99 0.155672
R693 VDD2.n99 VDD2.n70 0.155672
R694 VDD2.n92 VDD2.n70 0.155672
R695 VDD2.n92 VDD2.n91 0.155672
R696 VDD2.n91 VDD2.n75 0.155672
R697 VDD2.n84 VDD2.n75 0.155672
R698 VDD2.n84 VDD2.n83 0.155672
R699 VDD2.n22 VDD2.n21 0.155672
R700 VDD2.n22 VDD2.n13 0.155672
R701 VDD2.n29 VDD2.n13 0.155672
R702 VDD2.n30 VDD2.n29 0.155672
R703 VDD2.n30 VDD2.n9 0.155672
R704 VDD2.n38 VDD2.n9 0.155672
R705 VDD2.n39 VDD2.n38 0.155672
R706 VDD2.n39 VDD2.n5 0.155672
R707 VDD2.n47 VDD2.n5 0.155672
R708 VDD2.n48 VDD2.n47 0.155672
R709 VDD2.n48 VDD2.n1 0.155672
R710 VDD2.n55 VDD2.n1 0.155672
R711 B.n766 B.n765 585
R712 B.n766 B.n113 585
R713 B.n769 B.n768 585
R714 B.n770 B.n160 585
R715 B.n772 B.n771 585
R716 B.n774 B.n159 585
R717 B.n777 B.n776 585
R718 B.n778 B.n158 585
R719 B.n780 B.n779 585
R720 B.n782 B.n157 585
R721 B.n785 B.n784 585
R722 B.n786 B.n156 585
R723 B.n788 B.n787 585
R724 B.n790 B.n155 585
R725 B.n793 B.n792 585
R726 B.n794 B.n154 585
R727 B.n796 B.n795 585
R728 B.n798 B.n153 585
R729 B.n801 B.n800 585
R730 B.n802 B.n152 585
R731 B.n804 B.n803 585
R732 B.n806 B.n151 585
R733 B.n809 B.n808 585
R734 B.n810 B.n150 585
R735 B.n812 B.n811 585
R736 B.n814 B.n149 585
R737 B.n817 B.n816 585
R738 B.n818 B.n148 585
R739 B.n820 B.n819 585
R740 B.n822 B.n147 585
R741 B.n825 B.n824 585
R742 B.n826 B.n146 585
R743 B.n828 B.n827 585
R744 B.n830 B.n145 585
R745 B.n833 B.n832 585
R746 B.n834 B.n144 585
R747 B.n836 B.n835 585
R748 B.n838 B.n143 585
R749 B.n841 B.n840 585
R750 B.n843 B.n140 585
R751 B.n845 B.n844 585
R752 B.n847 B.n139 585
R753 B.n850 B.n849 585
R754 B.n851 B.n138 585
R755 B.n853 B.n852 585
R756 B.n855 B.n137 585
R757 B.n857 B.n856 585
R758 B.n859 B.n858 585
R759 B.n862 B.n861 585
R760 B.n863 B.n132 585
R761 B.n865 B.n864 585
R762 B.n867 B.n131 585
R763 B.n870 B.n869 585
R764 B.n871 B.n130 585
R765 B.n873 B.n872 585
R766 B.n875 B.n129 585
R767 B.n878 B.n877 585
R768 B.n879 B.n128 585
R769 B.n881 B.n880 585
R770 B.n883 B.n127 585
R771 B.n886 B.n885 585
R772 B.n887 B.n126 585
R773 B.n889 B.n888 585
R774 B.n891 B.n125 585
R775 B.n894 B.n893 585
R776 B.n895 B.n124 585
R777 B.n897 B.n896 585
R778 B.n899 B.n123 585
R779 B.n902 B.n901 585
R780 B.n903 B.n122 585
R781 B.n905 B.n904 585
R782 B.n907 B.n121 585
R783 B.n910 B.n909 585
R784 B.n911 B.n120 585
R785 B.n913 B.n912 585
R786 B.n915 B.n119 585
R787 B.n918 B.n917 585
R788 B.n919 B.n118 585
R789 B.n921 B.n920 585
R790 B.n923 B.n117 585
R791 B.n926 B.n925 585
R792 B.n927 B.n116 585
R793 B.n929 B.n928 585
R794 B.n931 B.n115 585
R795 B.n934 B.n933 585
R796 B.n935 B.n114 585
R797 B.n764 B.n112 585
R798 B.n938 B.n112 585
R799 B.n763 B.n111 585
R800 B.n939 B.n111 585
R801 B.n762 B.n110 585
R802 B.n940 B.n110 585
R803 B.n761 B.n760 585
R804 B.n760 B.n106 585
R805 B.n759 B.n105 585
R806 B.n946 B.n105 585
R807 B.n758 B.n104 585
R808 B.n947 B.n104 585
R809 B.n757 B.n103 585
R810 B.n948 B.n103 585
R811 B.n756 B.n755 585
R812 B.n755 B.n102 585
R813 B.n754 B.n98 585
R814 B.n954 B.n98 585
R815 B.n753 B.n97 585
R816 B.n955 B.n97 585
R817 B.n752 B.n96 585
R818 B.n956 B.n96 585
R819 B.n751 B.n750 585
R820 B.n750 B.n92 585
R821 B.n749 B.n91 585
R822 B.n962 B.n91 585
R823 B.n748 B.n90 585
R824 B.n963 B.n90 585
R825 B.n747 B.n89 585
R826 B.n964 B.n89 585
R827 B.n746 B.n745 585
R828 B.n745 B.n85 585
R829 B.n744 B.n84 585
R830 B.n970 B.n84 585
R831 B.n743 B.n83 585
R832 B.n971 B.n83 585
R833 B.n742 B.n82 585
R834 B.n972 B.n82 585
R835 B.n741 B.n740 585
R836 B.n740 B.n81 585
R837 B.n739 B.n77 585
R838 B.n978 B.n77 585
R839 B.n738 B.n76 585
R840 B.n979 B.n76 585
R841 B.n737 B.n75 585
R842 B.n980 B.n75 585
R843 B.n736 B.n735 585
R844 B.n735 B.n71 585
R845 B.n734 B.n70 585
R846 B.n986 B.n70 585
R847 B.n733 B.n69 585
R848 B.n987 B.n69 585
R849 B.n732 B.n68 585
R850 B.n988 B.n68 585
R851 B.n731 B.n730 585
R852 B.n730 B.n64 585
R853 B.n729 B.n63 585
R854 B.n994 B.n63 585
R855 B.n728 B.n62 585
R856 B.n995 B.n62 585
R857 B.n727 B.n61 585
R858 B.n996 B.n61 585
R859 B.n726 B.n725 585
R860 B.n725 B.n57 585
R861 B.n724 B.n56 585
R862 B.n1002 B.n56 585
R863 B.n723 B.n55 585
R864 B.n1003 B.n55 585
R865 B.n722 B.n54 585
R866 B.n1004 B.n54 585
R867 B.n721 B.n720 585
R868 B.n720 B.n50 585
R869 B.n719 B.n49 585
R870 B.n1010 B.n49 585
R871 B.n718 B.n48 585
R872 B.n1011 B.n48 585
R873 B.n717 B.n47 585
R874 B.n1012 B.n47 585
R875 B.n716 B.n715 585
R876 B.n715 B.n43 585
R877 B.n714 B.n42 585
R878 B.n1018 B.n42 585
R879 B.n713 B.n41 585
R880 B.n1019 B.n41 585
R881 B.n712 B.n40 585
R882 B.n1020 B.n40 585
R883 B.n711 B.n710 585
R884 B.n710 B.n36 585
R885 B.n709 B.n35 585
R886 B.n1026 B.n35 585
R887 B.n708 B.n34 585
R888 B.n1027 B.n34 585
R889 B.n707 B.n33 585
R890 B.n1028 B.n33 585
R891 B.n706 B.n705 585
R892 B.n705 B.n29 585
R893 B.n704 B.n28 585
R894 B.n1034 B.n28 585
R895 B.n703 B.n27 585
R896 B.n1035 B.n27 585
R897 B.n702 B.n26 585
R898 B.n1036 B.n26 585
R899 B.n701 B.n700 585
R900 B.n700 B.n22 585
R901 B.n699 B.n21 585
R902 B.n1042 B.n21 585
R903 B.n698 B.n20 585
R904 B.n1043 B.n20 585
R905 B.n697 B.n19 585
R906 B.n1044 B.n19 585
R907 B.n696 B.n695 585
R908 B.n695 B.n18 585
R909 B.n694 B.n14 585
R910 B.n1050 B.n14 585
R911 B.n693 B.n13 585
R912 B.n1051 B.n13 585
R913 B.n692 B.n12 585
R914 B.n1052 B.n12 585
R915 B.n691 B.n690 585
R916 B.n690 B.n8 585
R917 B.n689 B.n7 585
R918 B.n1058 B.n7 585
R919 B.n688 B.n6 585
R920 B.n1059 B.n6 585
R921 B.n687 B.n5 585
R922 B.n1060 B.n5 585
R923 B.n686 B.n685 585
R924 B.n685 B.n4 585
R925 B.n684 B.n161 585
R926 B.n684 B.n683 585
R927 B.n674 B.n162 585
R928 B.n163 B.n162 585
R929 B.n676 B.n675 585
R930 B.n677 B.n676 585
R931 B.n673 B.n168 585
R932 B.n168 B.n167 585
R933 B.n672 B.n671 585
R934 B.n671 B.n670 585
R935 B.n170 B.n169 585
R936 B.n663 B.n170 585
R937 B.n662 B.n661 585
R938 B.n664 B.n662 585
R939 B.n660 B.n175 585
R940 B.n175 B.n174 585
R941 B.n659 B.n658 585
R942 B.n658 B.n657 585
R943 B.n177 B.n176 585
R944 B.n178 B.n177 585
R945 B.n650 B.n649 585
R946 B.n651 B.n650 585
R947 B.n648 B.n183 585
R948 B.n183 B.n182 585
R949 B.n647 B.n646 585
R950 B.n646 B.n645 585
R951 B.n185 B.n184 585
R952 B.n186 B.n185 585
R953 B.n638 B.n637 585
R954 B.n639 B.n638 585
R955 B.n636 B.n191 585
R956 B.n191 B.n190 585
R957 B.n635 B.n634 585
R958 B.n634 B.n633 585
R959 B.n193 B.n192 585
R960 B.n194 B.n193 585
R961 B.n626 B.n625 585
R962 B.n627 B.n626 585
R963 B.n624 B.n199 585
R964 B.n199 B.n198 585
R965 B.n623 B.n622 585
R966 B.n622 B.n621 585
R967 B.n201 B.n200 585
R968 B.n202 B.n201 585
R969 B.n614 B.n613 585
R970 B.n615 B.n614 585
R971 B.n612 B.n206 585
R972 B.n210 B.n206 585
R973 B.n611 B.n610 585
R974 B.n610 B.n609 585
R975 B.n208 B.n207 585
R976 B.n209 B.n208 585
R977 B.n602 B.n601 585
R978 B.n603 B.n602 585
R979 B.n600 B.n215 585
R980 B.n215 B.n214 585
R981 B.n599 B.n598 585
R982 B.n598 B.n597 585
R983 B.n217 B.n216 585
R984 B.n218 B.n217 585
R985 B.n590 B.n589 585
R986 B.n591 B.n590 585
R987 B.n588 B.n223 585
R988 B.n223 B.n222 585
R989 B.n587 B.n586 585
R990 B.n586 B.n585 585
R991 B.n225 B.n224 585
R992 B.n226 B.n225 585
R993 B.n578 B.n577 585
R994 B.n579 B.n578 585
R995 B.n576 B.n231 585
R996 B.n231 B.n230 585
R997 B.n575 B.n574 585
R998 B.n574 B.n573 585
R999 B.n233 B.n232 585
R1000 B.n234 B.n233 585
R1001 B.n566 B.n565 585
R1002 B.n567 B.n566 585
R1003 B.n564 B.n239 585
R1004 B.n239 B.n238 585
R1005 B.n563 B.n562 585
R1006 B.n562 B.n561 585
R1007 B.n241 B.n240 585
R1008 B.n554 B.n241 585
R1009 B.n553 B.n552 585
R1010 B.n555 B.n553 585
R1011 B.n551 B.n246 585
R1012 B.n246 B.n245 585
R1013 B.n550 B.n549 585
R1014 B.n549 B.n548 585
R1015 B.n248 B.n247 585
R1016 B.n249 B.n248 585
R1017 B.n541 B.n540 585
R1018 B.n542 B.n541 585
R1019 B.n539 B.n254 585
R1020 B.n254 B.n253 585
R1021 B.n538 B.n537 585
R1022 B.n537 B.n536 585
R1023 B.n256 B.n255 585
R1024 B.n257 B.n256 585
R1025 B.n529 B.n528 585
R1026 B.n530 B.n529 585
R1027 B.n527 B.n262 585
R1028 B.n262 B.n261 585
R1029 B.n526 B.n525 585
R1030 B.n525 B.n524 585
R1031 B.n264 B.n263 585
R1032 B.n517 B.n264 585
R1033 B.n516 B.n515 585
R1034 B.n518 B.n516 585
R1035 B.n514 B.n269 585
R1036 B.n269 B.n268 585
R1037 B.n513 B.n512 585
R1038 B.n512 B.n511 585
R1039 B.n271 B.n270 585
R1040 B.n272 B.n271 585
R1041 B.n504 B.n503 585
R1042 B.n505 B.n504 585
R1043 B.n502 B.n277 585
R1044 B.n277 B.n276 585
R1045 B.n501 B.n500 585
R1046 B.n500 B.n499 585
R1047 B.n496 B.n281 585
R1048 B.n495 B.n494 585
R1049 B.n492 B.n282 585
R1050 B.n492 B.n280 585
R1051 B.n491 B.n490 585
R1052 B.n489 B.n488 585
R1053 B.n487 B.n284 585
R1054 B.n485 B.n484 585
R1055 B.n483 B.n285 585
R1056 B.n482 B.n481 585
R1057 B.n479 B.n286 585
R1058 B.n477 B.n476 585
R1059 B.n475 B.n287 585
R1060 B.n474 B.n473 585
R1061 B.n471 B.n288 585
R1062 B.n469 B.n468 585
R1063 B.n467 B.n289 585
R1064 B.n466 B.n465 585
R1065 B.n463 B.n290 585
R1066 B.n461 B.n460 585
R1067 B.n459 B.n291 585
R1068 B.n458 B.n457 585
R1069 B.n455 B.n292 585
R1070 B.n453 B.n452 585
R1071 B.n451 B.n293 585
R1072 B.n450 B.n449 585
R1073 B.n447 B.n294 585
R1074 B.n445 B.n444 585
R1075 B.n443 B.n295 585
R1076 B.n442 B.n441 585
R1077 B.n439 B.n296 585
R1078 B.n437 B.n436 585
R1079 B.n435 B.n297 585
R1080 B.n434 B.n433 585
R1081 B.n431 B.n298 585
R1082 B.n429 B.n428 585
R1083 B.n427 B.n299 585
R1084 B.n426 B.n425 585
R1085 B.n423 B.n300 585
R1086 B.n421 B.n420 585
R1087 B.n419 B.n301 585
R1088 B.n418 B.n417 585
R1089 B.n415 B.n305 585
R1090 B.n413 B.n412 585
R1091 B.n411 B.n306 585
R1092 B.n410 B.n409 585
R1093 B.n407 B.n307 585
R1094 B.n405 B.n404 585
R1095 B.n402 B.n308 585
R1096 B.n401 B.n400 585
R1097 B.n398 B.n311 585
R1098 B.n396 B.n395 585
R1099 B.n394 B.n312 585
R1100 B.n393 B.n392 585
R1101 B.n390 B.n313 585
R1102 B.n388 B.n387 585
R1103 B.n386 B.n314 585
R1104 B.n385 B.n384 585
R1105 B.n382 B.n315 585
R1106 B.n380 B.n379 585
R1107 B.n378 B.n316 585
R1108 B.n377 B.n376 585
R1109 B.n374 B.n317 585
R1110 B.n372 B.n371 585
R1111 B.n370 B.n318 585
R1112 B.n369 B.n368 585
R1113 B.n366 B.n319 585
R1114 B.n364 B.n363 585
R1115 B.n362 B.n320 585
R1116 B.n361 B.n360 585
R1117 B.n358 B.n321 585
R1118 B.n356 B.n355 585
R1119 B.n354 B.n322 585
R1120 B.n353 B.n352 585
R1121 B.n350 B.n323 585
R1122 B.n348 B.n347 585
R1123 B.n346 B.n324 585
R1124 B.n345 B.n344 585
R1125 B.n342 B.n325 585
R1126 B.n340 B.n339 585
R1127 B.n338 B.n326 585
R1128 B.n337 B.n336 585
R1129 B.n334 B.n327 585
R1130 B.n332 B.n331 585
R1131 B.n330 B.n329 585
R1132 B.n279 B.n278 585
R1133 B.n498 B.n497 585
R1134 B.n499 B.n498 585
R1135 B.n275 B.n274 585
R1136 B.n276 B.n275 585
R1137 B.n507 B.n506 585
R1138 B.n506 B.n505 585
R1139 B.n508 B.n273 585
R1140 B.n273 B.n272 585
R1141 B.n510 B.n509 585
R1142 B.n511 B.n510 585
R1143 B.n267 B.n266 585
R1144 B.n268 B.n267 585
R1145 B.n520 B.n519 585
R1146 B.n519 B.n518 585
R1147 B.n521 B.n265 585
R1148 B.n517 B.n265 585
R1149 B.n523 B.n522 585
R1150 B.n524 B.n523 585
R1151 B.n260 B.n259 585
R1152 B.n261 B.n260 585
R1153 B.n532 B.n531 585
R1154 B.n531 B.n530 585
R1155 B.n533 B.n258 585
R1156 B.n258 B.n257 585
R1157 B.n535 B.n534 585
R1158 B.n536 B.n535 585
R1159 B.n252 B.n251 585
R1160 B.n253 B.n252 585
R1161 B.n544 B.n543 585
R1162 B.n543 B.n542 585
R1163 B.n545 B.n250 585
R1164 B.n250 B.n249 585
R1165 B.n547 B.n546 585
R1166 B.n548 B.n547 585
R1167 B.n244 B.n243 585
R1168 B.n245 B.n244 585
R1169 B.n557 B.n556 585
R1170 B.n556 B.n555 585
R1171 B.n558 B.n242 585
R1172 B.n554 B.n242 585
R1173 B.n560 B.n559 585
R1174 B.n561 B.n560 585
R1175 B.n237 B.n236 585
R1176 B.n238 B.n237 585
R1177 B.n569 B.n568 585
R1178 B.n568 B.n567 585
R1179 B.n570 B.n235 585
R1180 B.n235 B.n234 585
R1181 B.n572 B.n571 585
R1182 B.n573 B.n572 585
R1183 B.n229 B.n228 585
R1184 B.n230 B.n229 585
R1185 B.n581 B.n580 585
R1186 B.n580 B.n579 585
R1187 B.n582 B.n227 585
R1188 B.n227 B.n226 585
R1189 B.n584 B.n583 585
R1190 B.n585 B.n584 585
R1191 B.n221 B.n220 585
R1192 B.n222 B.n221 585
R1193 B.n593 B.n592 585
R1194 B.n592 B.n591 585
R1195 B.n594 B.n219 585
R1196 B.n219 B.n218 585
R1197 B.n596 B.n595 585
R1198 B.n597 B.n596 585
R1199 B.n213 B.n212 585
R1200 B.n214 B.n213 585
R1201 B.n605 B.n604 585
R1202 B.n604 B.n603 585
R1203 B.n606 B.n211 585
R1204 B.n211 B.n209 585
R1205 B.n608 B.n607 585
R1206 B.n609 B.n608 585
R1207 B.n205 B.n204 585
R1208 B.n210 B.n205 585
R1209 B.n617 B.n616 585
R1210 B.n616 B.n615 585
R1211 B.n618 B.n203 585
R1212 B.n203 B.n202 585
R1213 B.n620 B.n619 585
R1214 B.n621 B.n620 585
R1215 B.n197 B.n196 585
R1216 B.n198 B.n197 585
R1217 B.n629 B.n628 585
R1218 B.n628 B.n627 585
R1219 B.n630 B.n195 585
R1220 B.n195 B.n194 585
R1221 B.n632 B.n631 585
R1222 B.n633 B.n632 585
R1223 B.n189 B.n188 585
R1224 B.n190 B.n189 585
R1225 B.n641 B.n640 585
R1226 B.n640 B.n639 585
R1227 B.n642 B.n187 585
R1228 B.n187 B.n186 585
R1229 B.n644 B.n643 585
R1230 B.n645 B.n644 585
R1231 B.n181 B.n180 585
R1232 B.n182 B.n181 585
R1233 B.n653 B.n652 585
R1234 B.n652 B.n651 585
R1235 B.n654 B.n179 585
R1236 B.n179 B.n178 585
R1237 B.n656 B.n655 585
R1238 B.n657 B.n656 585
R1239 B.n173 B.n172 585
R1240 B.n174 B.n173 585
R1241 B.n666 B.n665 585
R1242 B.n665 B.n664 585
R1243 B.n667 B.n171 585
R1244 B.n663 B.n171 585
R1245 B.n669 B.n668 585
R1246 B.n670 B.n669 585
R1247 B.n166 B.n165 585
R1248 B.n167 B.n166 585
R1249 B.n679 B.n678 585
R1250 B.n678 B.n677 585
R1251 B.n680 B.n164 585
R1252 B.n164 B.n163 585
R1253 B.n682 B.n681 585
R1254 B.n683 B.n682 585
R1255 B.n2 B.n0 585
R1256 B.n4 B.n2 585
R1257 B.n3 B.n1 585
R1258 B.n1059 B.n3 585
R1259 B.n1057 B.n1056 585
R1260 B.n1058 B.n1057 585
R1261 B.n1055 B.n9 585
R1262 B.n9 B.n8 585
R1263 B.n1054 B.n1053 585
R1264 B.n1053 B.n1052 585
R1265 B.n11 B.n10 585
R1266 B.n1051 B.n11 585
R1267 B.n1049 B.n1048 585
R1268 B.n1050 B.n1049 585
R1269 B.n1047 B.n15 585
R1270 B.n18 B.n15 585
R1271 B.n1046 B.n1045 585
R1272 B.n1045 B.n1044 585
R1273 B.n17 B.n16 585
R1274 B.n1043 B.n17 585
R1275 B.n1041 B.n1040 585
R1276 B.n1042 B.n1041 585
R1277 B.n1039 B.n23 585
R1278 B.n23 B.n22 585
R1279 B.n1038 B.n1037 585
R1280 B.n1037 B.n1036 585
R1281 B.n25 B.n24 585
R1282 B.n1035 B.n25 585
R1283 B.n1033 B.n1032 585
R1284 B.n1034 B.n1033 585
R1285 B.n1031 B.n30 585
R1286 B.n30 B.n29 585
R1287 B.n1030 B.n1029 585
R1288 B.n1029 B.n1028 585
R1289 B.n32 B.n31 585
R1290 B.n1027 B.n32 585
R1291 B.n1025 B.n1024 585
R1292 B.n1026 B.n1025 585
R1293 B.n1023 B.n37 585
R1294 B.n37 B.n36 585
R1295 B.n1022 B.n1021 585
R1296 B.n1021 B.n1020 585
R1297 B.n39 B.n38 585
R1298 B.n1019 B.n39 585
R1299 B.n1017 B.n1016 585
R1300 B.n1018 B.n1017 585
R1301 B.n1015 B.n44 585
R1302 B.n44 B.n43 585
R1303 B.n1014 B.n1013 585
R1304 B.n1013 B.n1012 585
R1305 B.n46 B.n45 585
R1306 B.n1011 B.n46 585
R1307 B.n1009 B.n1008 585
R1308 B.n1010 B.n1009 585
R1309 B.n1007 B.n51 585
R1310 B.n51 B.n50 585
R1311 B.n1006 B.n1005 585
R1312 B.n1005 B.n1004 585
R1313 B.n53 B.n52 585
R1314 B.n1003 B.n53 585
R1315 B.n1001 B.n1000 585
R1316 B.n1002 B.n1001 585
R1317 B.n999 B.n58 585
R1318 B.n58 B.n57 585
R1319 B.n998 B.n997 585
R1320 B.n997 B.n996 585
R1321 B.n60 B.n59 585
R1322 B.n995 B.n60 585
R1323 B.n993 B.n992 585
R1324 B.n994 B.n993 585
R1325 B.n991 B.n65 585
R1326 B.n65 B.n64 585
R1327 B.n990 B.n989 585
R1328 B.n989 B.n988 585
R1329 B.n67 B.n66 585
R1330 B.n987 B.n67 585
R1331 B.n985 B.n984 585
R1332 B.n986 B.n985 585
R1333 B.n983 B.n72 585
R1334 B.n72 B.n71 585
R1335 B.n982 B.n981 585
R1336 B.n981 B.n980 585
R1337 B.n74 B.n73 585
R1338 B.n979 B.n74 585
R1339 B.n977 B.n976 585
R1340 B.n978 B.n977 585
R1341 B.n975 B.n78 585
R1342 B.n81 B.n78 585
R1343 B.n974 B.n973 585
R1344 B.n973 B.n972 585
R1345 B.n80 B.n79 585
R1346 B.n971 B.n80 585
R1347 B.n969 B.n968 585
R1348 B.n970 B.n969 585
R1349 B.n967 B.n86 585
R1350 B.n86 B.n85 585
R1351 B.n966 B.n965 585
R1352 B.n965 B.n964 585
R1353 B.n88 B.n87 585
R1354 B.n963 B.n88 585
R1355 B.n961 B.n960 585
R1356 B.n962 B.n961 585
R1357 B.n959 B.n93 585
R1358 B.n93 B.n92 585
R1359 B.n958 B.n957 585
R1360 B.n957 B.n956 585
R1361 B.n95 B.n94 585
R1362 B.n955 B.n95 585
R1363 B.n953 B.n952 585
R1364 B.n954 B.n953 585
R1365 B.n951 B.n99 585
R1366 B.n102 B.n99 585
R1367 B.n950 B.n949 585
R1368 B.n949 B.n948 585
R1369 B.n101 B.n100 585
R1370 B.n947 B.n101 585
R1371 B.n945 B.n944 585
R1372 B.n946 B.n945 585
R1373 B.n943 B.n107 585
R1374 B.n107 B.n106 585
R1375 B.n942 B.n941 585
R1376 B.n941 B.n940 585
R1377 B.n109 B.n108 585
R1378 B.n939 B.n109 585
R1379 B.n937 B.n936 585
R1380 B.n938 B.n937 585
R1381 B.n1062 B.n1061 585
R1382 B.n1061 B.n1060 585
R1383 B.n498 B.n281 559.769
R1384 B.n937 B.n114 559.769
R1385 B.n500 B.n279 559.769
R1386 B.n766 B.n112 559.769
R1387 B.n309 B.t16 319.286
R1388 B.n141 B.t18 319.286
R1389 B.n302 B.t22 319.286
R1390 B.n133 B.t11 319.286
R1391 B.n309 B.t13 302.363
R1392 B.n302 B.t20 302.363
R1393 B.n133 B.t9 302.363
R1394 B.n141 B.t17 302.363
R1395 B.n310 B.t15 259.748
R1396 B.n142 B.t19 259.748
R1397 B.n303 B.t21 259.748
R1398 B.n134 B.t12 259.748
R1399 B.n767 B.n113 256.663
R1400 B.n773 B.n113 256.663
R1401 B.n775 B.n113 256.663
R1402 B.n781 B.n113 256.663
R1403 B.n783 B.n113 256.663
R1404 B.n789 B.n113 256.663
R1405 B.n791 B.n113 256.663
R1406 B.n797 B.n113 256.663
R1407 B.n799 B.n113 256.663
R1408 B.n805 B.n113 256.663
R1409 B.n807 B.n113 256.663
R1410 B.n813 B.n113 256.663
R1411 B.n815 B.n113 256.663
R1412 B.n821 B.n113 256.663
R1413 B.n823 B.n113 256.663
R1414 B.n829 B.n113 256.663
R1415 B.n831 B.n113 256.663
R1416 B.n837 B.n113 256.663
R1417 B.n839 B.n113 256.663
R1418 B.n846 B.n113 256.663
R1419 B.n848 B.n113 256.663
R1420 B.n854 B.n113 256.663
R1421 B.n136 B.n113 256.663
R1422 B.n860 B.n113 256.663
R1423 B.n866 B.n113 256.663
R1424 B.n868 B.n113 256.663
R1425 B.n874 B.n113 256.663
R1426 B.n876 B.n113 256.663
R1427 B.n882 B.n113 256.663
R1428 B.n884 B.n113 256.663
R1429 B.n890 B.n113 256.663
R1430 B.n892 B.n113 256.663
R1431 B.n898 B.n113 256.663
R1432 B.n900 B.n113 256.663
R1433 B.n906 B.n113 256.663
R1434 B.n908 B.n113 256.663
R1435 B.n914 B.n113 256.663
R1436 B.n916 B.n113 256.663
R1437 B.n922 B.n113 256.663
R1438 B.n924 B.n113 256.663
R1439 B.n930 B.n113 256.663
R1440 B.n932 B.n113 256.663
R1441 B.n493 B.n280 256.663
R1442 B.n283 B.n280 256.663
R1443 B.n486 B.n280 256.663
R1444 B.n480 B.n280 256.663
R1445 B.n478 B.n280 256.663
R1446 B.n472 B.n280 256.663
R1447 B.n470 B.n280 256.663
R1448 B.n464 B.n280 256.663
R1449 B.n462 B.n280 256.663
R1450 B.n456 B.n280 256.663
R1451 B.n454 B.n280 256.663
R1452 B.n448 B.n280 256.663
R1453 B.n446 B.n280 256.663
R1454 B.n440 B.n280 256.663
R1455 B.n438 B.n280 256.663
R1456 B.n432 B.n280 256.663
R1457 B.n430 B.n280 256.663
R1458 B.n424 B.n280 256.663
R1459 B.n422 B.n280 256.663
R1460 B.n416 B.n280 256.663
R1461 B.n414 B.n280 256.663
R1462 B.n408 B.n280 256.663
R1463 B.n406 B.n280 256.663
R1464 B.n399 B.n280 256.663
R1465 B.n397 B.n280 256.663
R1466 B.n391 B.n280 256.663
R1467 B.n389 B.n280 256.663
R1468 B.n383 B.n280 256.663
R1469 B.n381 B.n280 256.663
R1470 B.n375 B.n280 256.663
R1471 B.n373 B.n280 256.663
R1472 B.n367 B.n280 256.663
R1473 B.n365 B.n280 256.663
R1474 B.n359 B.n280 256.663
R1475 B.n357 B.n280 256.663
R1476 B.n351 B.n280 256.663
R1477 B.n349 B.n280 256.663
R1478 B.n343 B.n280 256.663
R1479 B.n341 B.n280 256.663
R1480 B.n335 B.n280 256.663
R1481 B.n333 B.n280 256.663
R1482 B.n328 B.n280 256.663
R1483 B.n498 B.n275 163.367
R1484 B.n506 B.n275 163.367
R1485 B.n506 B.n273 163.367
R1486 B.n510 B.n273 163.367
R1487 B.n510 B.n267 163.367
R1488 B.n519 B.n267 163.367
R1489 B.n519 B.n265 163.367
R1490 B.n523 B.n265 163.367
R1491 B.n523 B.n260 163.367
R1492 B.n531 B.n260 163.367
R1493 B.n531 B.n258 163.367
R1494 B.n535 B.n258 163.367
R1495 B.n535 B.n252 163.367
R1496 B.n543 B.n252 163.367
R1497 B.n543 B.n250 163.367
R1498 B.n547 B.n250 163.367
R1499 B.n547 B.n244 163.367
R1500 B.n556 B.n244 163.367
R1501 B.n556 B.n242 163.367
R1502 B.n560 B.n242 163.367
R1503 B.n560 B.n237 163.367
R1504 B.n568 B.n237 163.367
R1505 B.n568 B.n235 163.367
R1506 B.n572 B.n235 163.367
R1507 B.n572 B.n229 163.367
R1508 B.n580 B.n229 163.367
R1509 B.n580 B.n227 163.367
R1510 B.n584 B.n227 163.367
R1511 B.n584 B.n221 163.367
R1512 B.n592 B.n221 163.367
R1513 B.n592 B.n219 163.367
R1514 B.n596 B.n219 163.367
R1515 B.n596 B.n213 163.367
R1516 B.n604 B.n213 163.367
R1517 B.n604 B.n211 163.367
R1518 B.n608 B.n211 163.367
R1519 B.n608 B.n205 163.367
R1520 B.n616 B.n205 163.367
R1521 B.n616 B.n203 163.367
R1522 B.n620 B.n203 163.367
R1523 B.n620 B.n197 163.367
R1524 B.n628 B.n197 163.367
R1525 B.n628 B.n195 163.367
R1526 B.n632 B.n195 163.367
R1527 B.n632 B.n189 163.367
R1528 B.n640 B.n189 163.367
R1529 B.n640 B.n187 163.367
R1530 B.n644 B.n187 163.367
R1531 B.n644 B.n181 163.367
R1532 B.n652 B.n181 163.367
R1533 B.n652 B.n179 163.367
R1534 B.n656 B.n179 163.367
R1535 B.n656 B.n173 163.367
R1536 B.n665 B.n173 163.367
R1537 B.n665 B.n171 163.367
R1538 B.n669 B.n171 163.367
R1539 B.n669 B.n166 163.367
R1540 B.n678 B.n166 163.367
R1541 B.n678 B.n164 163.367
R1542 B.n682 B.n164 163.367
R1543 B.n682 B.n2 163.367
R1544 B.n1061 B.n2 163.367
R1545 B.n1061 B.n3 163.367
R1546 B.n1057 B.n3 163.367
R1547 B.n1057 B.n9 163.367
R1548 B.n1053 B.n9 163.367
R1549 B.n1053 B.n11 163.367
R1550 B.n1049 B.n11 163.367
R1551 B.n1049 B.n15 163.367
R1552 B.n1045 B.n15 163.367
R1553 B.n1045 B.n17 163.367
R1554 B.n1041 B.n17 163.367
R1555 B.n1041 B.n23 163.367
R1556 B.n1037 B.n23 163.367
R1557 B.n1037 B.n25 163.367
R1558 B.n1033 B.n25 163.367
R1559 B.n1033 B.n30 163.367
R1560 B.n1029 B.n30 163.367
R1561 B.n1029 B.n32 163.367
R1562 B.n1025 B.n32 163.367
R1563 B.n1025 B.n37 163.367
R1564 B.n1021 B.n37 163.367
R1565 B.n1021 B.n39 163.367
R1566 B.n1017 B.n39 163.367
R1567 B.n1017 B.n44 163.367
R1568 B.n1013 B.n44 163.367
R1569 B.n1013 B.n46 163.367
R1570 B.n1009 B.n46 163.367
R1571 B.n1009 B.n51 163.367
R1572 B.n1005 B.n51 163.367
R1573 B.n1005 B.n53 163.367
R1574 B.n1001 B.n53 163.367
R1575 B.n1001 B.n58 163.367
R1576 B.n997 B.n58 163.367
R1577 B.n997 B.n60 163.367
R1578 B.n993 B.n60 163.367
R1579 B.n993 B.n65 163.367
R1580 B.n989 B.n65 163.367
R1581 B.n989 B.n67 163.367
R1582 B.n985 B.n67 163.367
R1583 B.n985 B.n72 163.367
R1584 B.n981 B.n72 163.367
R1585 B.n981 B.n74 163.367
R1586 B.n977 B.n74 163.367
R1587 B.n977 B.n78 163.367
R1588 B.n973 B.n78 163.367
R1589 B.n973 B.n80 163.367
R1590 B.n969 B.n80 163.367
R1591 B.n969 B.n86 163.367
R1592 B.n965 B.n86 163.367
R1593 B.n965 B.n88 163.367
R1594 B.n961 B.n88 163.367
R1595 B.n961 B.n93 163.367
R1596 B.n957 B.n93 163.367
R1597 B.n957 B.n95 163.367
R1598 B.n953 B.n95 163.367
R1599 B.n953 B.n99 163.367
R1600 B.n949 B.n99 163.367
R1601 B.n949 B.n101 163.367
R1602 B.n945 B.n101 163.367
R1603 B.n945 B.n107 163.367
R1604 B.n941 B.n107 163.367
R1605 B.n941 B.n109 163.367
R1606 B.n937 B.n109 163.367
R1607 B.n494 B.n492 163.367
R1608 B.n492 B.n491 163.367
R1609 B.n488 B.n487 163.367
R1610 B.n485 B.n285 163.367
R1611 B.n481 B.n479 163.367
R1612 B.n477 B.n287 163.367
R1613 B.n473 B.n471 163.367
R1614 B.n469 B.n289 163.367
R1615 B.n465 B.n463 163.367
R1616 B.n461 B.n291 163.367
R1617 B.n457 B.n455 163.367
R1618 B.n453 B.n293 163.367
R1619 B.n449 B.n447 163.367
R1620 B.n445 B.n295 163.367
R1621 B.n441 B.n439 163.367
R1622 B.n437 B.n297 163.367
R1623 B.n433 B.n431 163.367
R1624 B.n429 B.n299 163.367
R1625 B.n425 B.n423 163.367
R1626 B.n421 B.n301 163.367
R1627 B.n417 B.n415 163.367
R1628 B.n413 B.n306 163.367
R1629 B.n409 B.n407 163.367
R1630 B.n405 B.n308 163.367
R1631 B.n400 B.n398 163.367
R1632 B.n396 B.n312 163.367
R1633 B.n392 B.n390 163.367
R1634 B.n388 B.n314 163.367
R1635 B.n384 B.n382 163.367
R1636 B.n380 B.n316 163.367
R1637 B.n376 B.n374 163.367
R1638 B.n372 B.n318 163.367
R1639 B.n368 B.n366 163.367
R1640 B.n364 B.n320 163.367
R1641 B.n360 B.n358 163.367
R1642 B.n356 B.n322 163.367
R1643 B.n352 B.n350 163.367
R1644 B.n348 B.n324 163.367
R1645 B.n344 B.n342 163.367
R1646 B.n340 B.n326 163.367
R1647 B.n336 B.n334 163.367
R1648 B.n332 B.n329 163.367
R1649 B.n500 B.n277 163.367
R1650 B.n504 B.n277 163.367
R1651 B.n504 B.n271 163.367
R1652 B.n512 B.n271 163.367
R1653 B.n512 B.n269 163.367
R1654 B.n516 B.n269 163.367
R1655 B.n516 B.n264 163.367
R1656 B.n525 B.n264 163.367
R1657 B.n525 B.n262 163.367
R1658 B.n529 B.n262 163.367
R1659 B.n529 B.n256 163.367
R1660 B.n537 B.n256 163.367
R1661 B.n537 B.n254 163.367
R1662 B.n541 B.n254 163.367
R1663 B.n541 B.n248 163.367
R1664 B.n549 B.n248 163.367
R1665 B.n549 B.n246 163.367
R1666 B.n553 B.n246 163.367
R1667 B.n553 B.n241 163.367
R1668 B.n562 B.n241 163.367
R1669 B.n562 B.n239 163.367
R1670 B.n566 B.n239 163.367
R1671 B.n566 B.n233 163.367
R1672 B.n574 B.n233 163.367
R1673 B.n574 B.n231 163.367
R1674 B.n578 B.n231 163.367
R1675 B.n578 B.n225 163.367
R1676 B.n586 B.n225 163.367
R1677 B.n586 B.n223 163.367
R1678 B.n590 B.n223 163.367
R1679 B.n590 B.n217 163.367
R1680 B.n598 B.n217 163.367
R1681 B.n598 B.n215 163.367
R1682 B.n602 B.n215 163.367
R1683 B.n602 B.n208 163.367
R1684 B.n610 B.n208 163.367
R1685 B.n610 B.n206 163.367
R1686 B.n614 B.n206 163.367
R1687 B.n614 B.n201 163.367
R1688 B.n622 B.n201 163.367
R1689 B.n622 B.n199 163.367
R1690 B.n626 B.n199 163.367
R1691 B.n626 B.n193 163.367
R1692 B.n634 B.n193 163.367
R1693 B.n634 B.n191 163.367
R1694 B.n638 B.n191 163.367
R1695 B.n638 B.n185 163.367
R1696 B.n646 B.n185 163.367
R1697 B.n646 B.n183 163.367
R1698 B.n650 B.n183 163.367
R1699 B.n650 B.n177 163.367
R1700 B.n658 B.n177 163.367
R1701 B.n658 B.n175 163.367
R1702 B.n662 B.n175 163.367
R1703 B.n662 B.n170 163.367
R1704 B.n671 B.n170 163.367
R1705 B.n671 B.n168 163.367
R1706 B.n676 B.n168 163.367
R1707 B.n676 B.n162 163.367
R1708 B.n684 B.n162 163.367
R1709 B.n685 B.n684 163.367
R1710 B.n685 B.n5 163.367
R1711 B.n6 B.n5 163.367
R1712 B.n7 B.n6 163.367
R1713 B.n690 B.n7 163.367
R1714 B.n690 B.n12 163.367
R1715 B.n13 B.n12 163.367
R1716 B.n14 B.n13 163.367
R1717 B.n695 B.n14 163.367
R1718 B.n695 B.n19 163.367
R1719 B.n20 B.n19 163.367
R1720 B.n21 B.n20 163.367
R1721 B.n700 B.n21 163.367
R1722 B.n700 B.n26 163.367
R1723 B.n27 B.n26 163.367
R1724 B.n28 B.n27 163.367
R1725 B.n705 B.n28 163.367
R1726 B.n705 B.n33 163.367
R1727 B.n34 B.n33 163.367
R1728 B.n35 B.n34 163.367
R1729 B.n710 B.n35 163.367
R1730 B.n710 B.n40 163.367
R1731 B.n41 B.n40 163.367
R1732 B.n42 B.n41 163.367
R1733 B.n715 B.n42 163.367
R1734 B.n715 B.n47 163.367
R1735 B.n48 B.n47 163.367
R1736 B.n49 B.n48 163.367
R1737 B.n720 B.n49 163.367
R1738 B.n720 B.n54 163.367
R1739 B.n55 B.n54 163.367
R1740 B.n56 B.n55 163.367
R1741 B.n725 B.n56 163.367
R1742 B.n725 B.n61 163.367
R1743 B.n62 B.n61 163.367
R1744 B.n63 B.n62 163.367
R1745 B.n730 B.n63 163.367
R1746 B.n730 B.n68 163.367
R1747 B.n69 B.n68 163.367
R1748 B.n70 B.n69 163.367
R1749 B.n735 B.n70 163.367
R1750 B.n735 B.n75 163.367
R1751 B.n76 B.n75 163.367
R1752 B.n77 B.n76 163.367
R1753 B.n740 B.n77 163.367
R1754 B.n740 B.n82 163.367
R1755 B.n83 B.n82 163.367
R1756 B.n84 B.n83 163.367
R1757 B.n745 B.n84 163.367
R1758 B.n745 B.n89 163.367
R1759 B.n90 B.n89 163.367
R1760 B.n91 B.n90 163.367
R1761 B.n750 B.n91 163.367
R1762 B.n750 B.n96 163.367
R1763 B.n97 B.n96 163.367
R1764 B.n98 B.n97 163.367
R1765 B.n755 B.n98 163.367
R1766 B.n755 B.n103 163.367
R1767 B.n104 B.n103 163.367
R1768 B.n105 B.n104 163.367
R1769 B.n760 B.n105 163.367
R1770 B.n760 B.n110 163.367
R1771 B.n111 B.n110 163.367
R1772 B.n112 B.n111 163.367
R1773 B.n933 B.n931 163.367
R1774 B.n929 B.n116 163.367
R1775 B.n925 B.n923 163.367
R1776 B.n921 B.n118 163.367
R1777 B.n917 B.n915 163.367
R1778 B.n913 B.n120 163.367
R1779 B.n909 B.n907 163.367
R1780 B.n905 B.n122 163.367
R1781 B.n901 B.n899 163.367
R1782 B.n897 B.n124 163.367
R1783 B.n893 B.n891 163.367
R1784 B.n889 B.n126 163.367
R1785 B.n885 B.n883 163.367
R1786 B.n881 B.n128 163.367
R1787 B.n877 B.n875 163.367
R1788 B.n873 B.n130 163.367
R1789 B.n869 B.n867 163.367
R1790 B.n865 B.n132 163.367
R1791 B.n861 B.n859 163.367
R1792 B.n856 B.n855 163.367
R1793 B.n853 B.n138 163.367
R1794 B.n849 B.n847 163.367
R1795 B.n845 B.n140 163.367
R1796 B.n840 B.n838 163.367
R1797 B.n836 B.n144 163.367
R1798 B.n832 B.n830 163.367
R1799 B.n828 B.n146 163.367
R1800 B.n824 B.n822 163.367
R1801 B.n820 B.n148 163.367
R1802 B.n816 B.n814 163.367
R1803 B.n812 B.n150 163.367
R1804 B.n808 B.n806 163.367
R1805 B.n804 B.n152 163.367
R1806 B.n800 B.n798 163.367
R1807 B.n796 B.n154 163.367
R1808 B.n792 B.n790 163.367
R1809 B.n788 B.n156 163.367
R1810 B.n784 B.n782 163.367
R1811 B.n780 B.n158 163.367
R1812 B.n776 B.n774 163.367
R1813 B.n772 B.n160 163.367
R1814 B.n768 B.n766 163.367
R1815 B.n499 B.n280 98.4669
R1816 B.n938 B.n113 98.4669
R1817 B.n493 B.n281 71.676
R1818 B.n491 B.n283 71.676
R1819 B.n487 B.n486 71.676
R1820 B.n480 B.n285 71.676
R1821 B.n479 B.n478 71.676
R1822 B.n472 B.n287 71.676
R1823 B.n471 B.n470 71.676
R1824 B.n464 B.n289 71.676
R1825 B.n463 B.n462 71.676
R1826 B.n456 B.n291 71.676
R1827 B.n455 B.n454 71.676
R1828 B.n448 B.n293 71.676
R1829 B.n447 B.n446 71.676
R1830 B.n440 B.n295 71.676
R1831 B.n439 B.n438 71.676
R1832 B.n432 B.n297 71.676
R1833 B.n431 B.n430 71.676
R1834 B.n424 B.n299 71.676
R1835 B.n423 B.n422 71.676
R1836 B.n416 B.n301 71.676
R1837 B.n415 B.n414 71.676
R1838 B.n408 B.n306 71.676
R1839 B.n407 B.n406 71.676
R1840 B.n399 B.n308 71.676
R1841 B.n398 B.n397 71.676
R1842 B.n391 B.n312 71.676
R1843 B.n390 B.n389 71.676
R1844 B.n383 B.n314 71.676
R1845 B.n382 B.n381 71.676
R1846 B.n375 B.n316 71.676
R1847 B.n374 B.n373 71.676
R1848 B.n367 B.n318 71.676
R1849 B.n366 B.n365 71.676
R1850 B.n359 B.n320 71.676
R1851 B.n358 B.n357 71.676
R1852 B.n351 B.n322 71.676
R1853 B.n350 B.n349 71.676
R1854 B.n343 B.n324 71.676
R1855 B.n342 B.n341 71.676
R1856 B.n335 B.n326 71.676
R1857 B.n334 B.n333 71.676
R1858 B.n329 B.n328 71.676
R1859 B.n932 B.n114 71.676
R1860 B.n931 B.n930 71.676
R1861 B.n924 B.n116 71.676
R1862 B.n923 B.n922 71.676
R1863 B.n916 B.n118 71.676
R1864 B.n915 B.n914 71.676
R1865 B.n908 B.n120 71.676
R1866 B.n907 B.n906 71.676
R1867 B.n900 B.n122 71.676
R1868 B.n899 B.n898 71.676
R1869 B.n892 B.n124 71.676
R1870 B.n891 B.n890 71.676
R1871 B.n884 B.n126 71.676
R1872 B.n883 B.n882 71.676
R1873 B.n876 B.n128 71.676
R1874 B.n875 B.n874 71.676
R1875 B.n868 B.n130 71.676
R1876 B.n867 B.n866 71.676
R1877 B.n860 B.n132 71.676
R1878 B.n859 B.n136 71.676
R1879 B.n855 B.n854 71.676
R1880 B.n848 B.n138 71.676
R1881 B.n847 B.n846 71.676
R1882 B.n839 B.n140 71.676
R1883 B.n838 B.n837 71.676
R1884 B.n831 B.n144 71.676
R1885 B.n830 B.n829 71.676
R1886 B.n823 B.n146 71.676
R1887 B.n822 B.n821 71.676
R1888 B.n815 B.n148 71.676
R1889 B.n814 B.n813 71.676
R1890 B.n807 B.n150 71.676
R1891 B.n806 B.n805 71.676
R1892 B.n799 B.n152 71.676
R1893 B.n798 B.n797 71.676
R1894 B.n791 B.n154 71.676
R1895 B.n790 B.n789 71.676
R1896 B.n783 B.n156 71.676
R1897 B.n782 B.n781 71.676
R1898 B.n775 B.n158 71.676
R1899 B.n774 B.n773 71.676
R1900 B.n767 B.n160 71.676
R1901 B.n768 B.n767 71.676
R1902 B.n773 B.n772 71.676
R1903 B.n776 B.n775 71.676
R1904 B.n781 B.n780 71.676
R1905 B.n784 B.n783 71.676
R1906 B.n789 B.n788 71.676
R1907 B.n792 B.n791 71.676
R1908 B.n797 B.n796 71.676
R1909 B.n800 B.n799 71.676
R1910 B.n805 B.n804 71.676
R1911 B.n808 B.n807 71.676
R1912 B.n813 B.n812 71.676
R1913 B.n816 B.n815 71.676
R1914 B.n821 B.n820 71.676
R1915 B.n824 B.n823 71.676
R1916 B.n829 B.n828 71.676
R1917 B.n832 B.n831 71.676
R1918 B.n837 B.n836 71.676
R1919 B.n840 B.n839 71.676
R1920 B.n846 B.n845 71.676
R1921 B.n849 B.n848 71.676
R1922 B.n854 B.n853 71.676
R1923 B.n856 B.n136 71.676
R1924 B.n861 B.n860 71.676
R1925 B.n866 B.n865 71.676
R1926 B.n869 B.n868 71.676
R1927 B.n874 B.n873 71.676
R1928 B.n877 B.n876 71.676
R1929 B.n882 B.n881 71.676
R1930 B.n885 B.n884 71.676
R1931 B.n890 B.n889 71.676
R1932 B.n893 B.n892 71.676
R1933 B.n898 B.n897 71.676
R1934 B.n901 B.n900 71.676
R1935 B.n906 B.n905 71.676
R1936 B.n909 B.n908 71.676
R1937 B.n914 B.n913 71.676
R1938 B.n917 B.n916 71.676
R1939 B.n922 B.n921 71.676
R1940 B.n925 B.n924 71.676
R1941 B.n930 B.n929 71.676
R1942 B.n933 B.n932 71.676
R1943 B.n494 B.n493 71.676
R1944 B.n488 B.n283 71.676
R1945 B.n486 B.n485 71.676
R1946 B.n481 B.n480 71.676
R1947 B.n478 B.n477 71.676
R1948 B.n473 B.n472 71.676
R1949 B.n470 B.n469 71.676
R1950 B.n465 B.n464 71.676
R1951 B.n462 B.n461 71.676
R1952 B.n457 B.n456 71.676
R1953 B.n454 B.n453 71.676
R1954 B.n449 B.n448 71.676
R1955 B.n446 B.n445 71.676
R1956 B.n441 B.n440 71.676
R1957 B.n438 B.n437 71.676
R1958 B.n433 B.n432 71.676
R1959 B.n430 B.n429 71.676
R1960 B.n425 B.n424 71.676
R1961 B.n422 B.n421 71.676
R1962 B.n417 B.n416 71.676
R1963 B.n414 B.n413 71.676
R1964 B.n409 B.n408 71.676
R1965 B.n406 B.n405 71.676
R1966 B.n400 B.n399 71.676
R1967 B.n397 B.n396 71.676
R1968 B.n392 B.n391 71.676
R1969 B.n389 B.n388 71.676
R1970 B.n384 B.n383 71.676
R1971 B.n381 B.n380 71.676
R1972 B.n376 B.n375 71.676
R1973 B.n373 B.n372 71.676
R1974 B.n368 B.n367 71.676
R1975 B.n365 B.n364 71.676
R1976 B.n360 B.n359 71.676
R1977 B.n357 B.n356 71.676
R1978 B.n352 B.n351 71.676
R1979 B.n349 B.n348 71.676
R1980 B.n344 B.n343 71.676
R1981 B.n341 B.n340 71.676
R1982 B.n336 B.n335 71.676
R1983 B.n333 B.n332 71.676
R1984 B.n328 B.n279 71.676
R1985 B.n403 B.n310 59.5399
R1986 B.n310 B.n309 59.5399
R1987 B.n304 B.n303 59.5399
R1988 B.n303 B.n302 59.5399
R1989 B.n134 B.n133 59.5399
R1990 B.n135 B.n134 59.5399
R1991 B.n142 B.n141 59.5399
R1992 B.n842 B.n142 59.5399
R1993 B.n499 B.n276 46.8237
R1994 B.n505 B.n276 46.8237
R1995 B.n505 B.n272 46.8237
R1996 B.n511 B.n272 46.8237
R1997 B.n511 B.n268 46.8237
R1998 B.n518 B.n268 46.8237
R1999 B.n518 B.n517 46.8237
R2000 B.n524 B.n261 46.8237
R2001 B.n530 B.n261 46.8237
R2002 B.n530 B.n257 46.8237
R2003 B.n536 B.n257 46.8237
R2004 B.n536 B.n253 46.8237
R2005 B.n542 B.n253 46.8237
R2006 B.n542 B.n249 46.8237
R2007 B.n548 B.n249 46.8237
R2008 B.n548 B.n245 46.8237
R2009 B.n555 B.n245 46.8237
R2010 B.n555 B.n554 46.8237
R2011 B.n561 B.n238 46.8237
R2012 B.n567 B.n238 46.8237
R2013 B.n567 B.n234 46.8237
R2014 B.n573 B.n234 46.8237
R2015 B.n573 B.n230 46.8237
R2016 B.n579 B.n230 46.8237
R2017 B.n579 B.n226 46.8237
R2018 B.n585 B.n226 46.8237
R2019 B.n591 B.n222 46.8237
R2020 B.n591 B.n218 46.8237
R2021 B.n597 B.n218 46.8237
R2022 B.n597 B.n214 46.8237
R2023 B.n603 B.n214 46.8237
R2024 B.n603 B.n209 46.8237
R2025 B.n609 B.n209 46.8237
R2026 B.n609 B.n210 46.8237
R2027 B.n615 B.n202 46.8237
R2028 B.n621 B.n202 46.8237
R2029 B.n621 B.n198 46.8237
R2030 B.n627 B.n198 46.8237
R2031 B.n627 B.n194 46.8237
R2032 B.n633 B.n194 46.8237
R2033 B.n633 B.n190 46.8237
R2034 B.n639 B.n190 46.8237
R2035 B.n645 B.n186 46.8237
R2036 B.n645 B.n182 46.8237
R2037 B.n651 B.n182 46.8237
R2038 B.n651 B.n178 46.8237
R2039 B.n657 B.n178 46.8237
R2040 B.n657 B.n174 46.8237
R2041 B.n664 B.n174 46.8237
R2042 B.n664 B.n663 46.8237
R2043 B.n670 B.n167 46.8237
R2044 B.n677 B.n167 46.8237
R2045 B.n677 B.n163 46.8237
R2046 B.n683 B.n163 46.8237
R2047 B.n683 B.n4 46.8237
R2048 B.n1060 B.n4 46.8237
R2049 B.n1060 B.n1059 46.8237
R2050 B.n1059 B.n1058 46.8237
R2051 B.n1058 B.n8 46.8237
R2052 B.n1052 B.n8 46.8237
R2053 B.n1052 B.n1051 46.8237
R2054 B.n1051 B.n1050 46.8237
R2055 B.n1044 B.n18 46.8237
R2056 B.n1044 B.n1043 46.8237
R2057 B.n1043 B.n1042 46.8237
R2058 B.n1042 B.n22 46.8237
R2059 B.n1036 B.n22 46.8237
R2060 B.n1036 B.n1035 46.8237
R2061 B.n1035 B.n1034 46.8237
R2062 B.n1034 B.n29 46.8237
R2063 B.n1028 B.n1027 46.8237
R2064 B.n1027 B.n1026 46.8237
R2065 B.n1026 B.n36 46.8237
R2066 B.n1020 B.n36 46.8237
R2067 B.n1020 B.n1019 46.8237
R2068 B.n1019 B.n1018 46.8237
R2069 B.n1018 B.n43 46.8237
R2070 B.n1012 B.n43 46.8237
R2071 B.n1011 B.n1010 46.8237
R2072 B.n1010 B.n50 46.8237
R2073 B.n1004 B.n50 46.8237
R2074 B.n1004 B.n1003 46.8237
R2075 B.n1003 B.n1002 46.8237
R2076 B.n1002 B.n57 46.8237
R2077 B.n996 B.n57 46.8237
R2078 B.n996 B.n995 46.8237
R2079 B.n994 B.n64 46.8237
R2080 B.n988 B.n64 46.8237
R2081 B.n988 B.n987 46.8237
R2082 B.n987 B.n986 46.8237
R2083 B.n986 B.n71 46.8237
R2084 B.n980 B.n71 46.8237
R2085 B.n980 B.n979 46.8237
R2086 B.n979 B.n978 46.8237
R2087 B.n972 B.n81 46.8237
R2088 B.n972 B.n971 46.8237
R2089 B.n971 B.n970 46.8237
R2090 B.n970 B.n85 46.8237
R2091 B.n964 B.n85 46.8237
R2092 B.n964 B.n963 46.8237
R2093 B.n963 B.n962 46.8237
R2094 B.n962 B.n92 46.8237
R2095 B.n956 B.n92 46.8237
R2096 B.n956 B.n955 46.8237
R2097 B.n955 B.n954 46.8237
R2098 B.n948 B.n102 46.8237
R2099 B.n948 B.n947 46.8237
R2100 B.n947 B.n946 46.8237
R2101 B.n946 B.n106 46.8237
R2102 B.n940 B.n106 46.8237
R2103 B.n940 B.n939 46.8237
R2104 B.n939 B.n938 46.8237
R2105 B.n663 B.t8 41.3151
R2106 B.n18 B.t4 41.3151
R2107 B.n639 B.t23 39.9379
R2108 B.n1028 B.t1 39.9379
R2109 B.n210 B.t7 38.5607
R2110 B.t2 B.n1011 38.5607
R2111 B.n585 B.t3 37.1836
R2112 B.t5 B.n994 37.1836
R2113 B.n765 B.n764 36.3712
R2114 B.n936 B.n935 36.3712
R2115 B.n501 B.n278 36.3712
R2116 B.n497 B.n496 36.3712
R2117 B.n554 B.t6 35.8064
R2118 B.n81 B.t0 35.8064
R2119 B.n517 B.t14 24.7892
R2120 B.n102 B.t10 24.7892
R2121 B.n524 B.t14 22.0349
R2122 B.n954 B.t10 22.0349
R2123 B B.n1062 18.0485
R2124 B.n561 B.t6 11.0177
R2125 B.n978 B.t0 11.0177
R2126 B.n935 B.n934 10.6151
R2127 B.n934 B.n115 10.6151
R2128 B.n928 B.n115 10.6151
R2129 B.n928 B.n927 10.6151
R2130 B.n927 B.n926 10.6151
R2131 B.n926 B.n117 10.6151
R2132 B.n920 B.n117 10.6151
R2133 B.n920 B.n919 10.6151
R2134 B.n919 B.n918 10.6151
R2135 B.n918 B.n119 10.6151
R2136 B.n912 B.n119 10.6151
R2137 B.n912 B.n911 10.6151
R2138 B.n911 B.n910 10.6151
R2139 B.n910 B.n121 10.6151
R2140 B.n904 B.n121 10.6151
R2141 B.n904 B.n903 10.6151
R2142 B.n903 B.n902 10.6151
R2143 B.n902 B.n123 10.6151
R2144 B.n896 B.n123 10.6151
R2145 B.n896 B.n895 10.6151
R2146 B.n895 B.n894 10.6151
R2147 B.n894 B.n125 10.6151
R2148 B.n888 B.n125 10.6151
R2149 B.n888 B.n887 10.6151
R2150 B.n887 B.n886 10.6151
R2151 B.n886 B.n127 10.6151
R2152 B.n880 B.n127 10.6151
R2153 B.n880 B.n879 10.6151
R2154 B.n879 B.n878 10.6151
R2155 B.n878 B.n129 10.6151
R2156 B.n872 B.n129 10.6151
R2157 B.n872 B.n871 10.6151
R2158 B.n871 B.n870 10.6151
R2159 B.n870 B.n131 10.6151
R2160 B.n864 B.n131 10.6151
R2161 B.n864 B.n863 10.6151
R2162 B.n863 B.n862 10.6151
R2163 B.n858 B.n857 10.6151
R2164 B.n857 B.n137 10.6151
R2165 B.n852 B.n137 10.6151
R2166 B.n852 B.n851 10.6151
R2167 B.n851 B.n850 10.6151
R2168 B.n850 B.n139 10.6151
R2169 B.n844 B.n139 10.6151
R2170 B.n844 B.n843 10.6151
R2171 B.n841 B.n143 10.6151
R2172 B.n835 B.n143 10.6151
R2173 B.n835 B.n834 10.6151
R2174 B.n834 B.n833 10.6151
R2175 B.n833 B.n145 10.6151
R2176 B.n827 B.n145 10.6151
R2177 B.n827 B.n826 10.6151
R2178 B.n826 B.n825 10.6151
R2179 B.n825 B.n147 10.6151
R2180 B.n819 B.n147 10.6151
R2181 B.n819 B.n818 10.6151
R2182 B.n818 B.n817 10.6151
R2183 B.n817 B.n149 10.6151
R2184 B.n811 B.n149 10.6151
R2185 B.n811 B.n810 10.6151
R2186 B.n810 B.n809 10.6151
R2187 B.n809 B.n151 10.6151
R2188 B.n803 B.n151 10.6151
R2189 B.n803 B.n802 10.6151
R2190 B.n802 B.n801 10.6151
R2191 B.n801 B.n153 10.6151
R2192 B.n795 B.n153 10.6151
R2193 B.n795 B.n794 10.6151
R2194 B.n794 B.n793 10.6151
R2195 B.n793 B.n155 10.6151
R2196 B.n787 B.n155 10.6151
R2197 B.n787 B.n786 10.6151
R2198 B.n786 B.n785 10.6151
R2199 B.n785 B.n157 10.6151
R2200 B.n779 B.n157 10.6151
R2201 B.n779 B.n778 10.6151
R2202 B.n778 B.n777 10.6151
R2203 B.n777 B.n159 10.6151
R2204 B.n771 B.n159 10.6151
R2205 B.n771 B.n770 10.6151
R2206 B.n770 B.n769 10.6151
R2207 B.n769 B.n765 10.6151
R2208 B.n502 B.n501 10.6151
R2209 B.n503 B.n502 10.6151
R2210 B.n503 B.n270 10.6151
R2211 B.n513 B.n270 10.6151
R2212 B.n514 B.n513 10.6151
R2213 B.n515 B.n514 10.6151
R2214 B.n515 B.n263 10.6151
R2215 B.n526 B.n263 10.6151
R2216 B.n527 B.n526 10.6151
R2217 B.n528 B.n527 10.6151
R2218 B.n528 B.n255 10.6151
R2219 B.n538 B.n255 10.6151
R2220 B.n539 B.n538 10.6151
R2221 B.n540 B.n539 10.6151
R2222 B.n540 B.n247 10.6151
R2223 B.n550 B.n247 10.6151
R2224 B.n551 B.n550 10.6151
R2225 B.n552 B.n551 10.6151
R2226 B.n552 B.n240 10.6151
R2227 B.n563 B.n240 10.6151
R2228 B.n564 B.n563 10.6151
R2229 B.n565 B.n564 10.6151
R2230 B.n565 B.n232 10.6151
R2231 B.n575 B.n232 10.6151
R2232 B.n576 B.n575 10.6151
R2233 B.n577 B.n576 10.6151
R2234 B.n577 B.n224 10.6151
R2235 B.n587 B.n224 10.6151
R2236 B.n588 B.n587 10.6151
R2237 B.n589 B.n588 10.6151
R2238 B.n589 B.n216 10.6151
R2239 B.n599 B.n216 10.6151
R2240 B.n600 B.n599 10.6151
R2241 B.n601 B.n600 10.6151
R2242 B.n601 B.n207 10.6151
R2243 B.n611 B.n207 10.6151
R2244 B.n612 B.n611 10.6151
R2245 B.n613 B.n612 10.6151
R2246 B.n613 B.n200 10.6151
R2247 B.n623 B.n200 10.6151
R2248 B.n624 B.n623 10.6151
R2249 B.n625 B.n624 10.6151
R2250 B.n625 B.n192 10.6151
R2251 B.n635 B.n192 10.6151
R2252 B.n636 B.n635 10.6151
R2253 B.n637 B.n636 10.6151
R2254 B.n637 B.n184 10.6151
R2255 B.n647 B.n184 10.6151
R2256 B.n648 B.n647 10.6151
R2257 B.n649 B.n648 10.6151
R2258 B.n649 B.n176 10.6151
R2259 B.n659 B.n176 10.6151
R2260 B.n660 B.n659 10.6151
R2261 B.n661 B.n660 10.6151
R2262 B.n661 B.n169 10.6151
R2263 B.n672 B.n169 10.6151
R2264 B.n673 B.n672 10.6151
R2265 B.n675 B.n673 10.6151
R2266 B.n675 B.n674 10.6151
R2267 B.n674 B.n161 10.6151
R2268 B.n686 B.n161 10.6151
R2269 B.n687 B.n686 10.6151
R2270 B.n688 B.n687 10.6151
R2271 B.n689 B.n688 10.6151
R2272 B.n691 B.n689 10.6151
R2273 B.n692 B.n691 10.6151
R2274 B.n693 B.n692 10.6151
R2275 B.n694 B.n693 10.6151
R2276 B.n696 B.n694 10.6151
R2277 B.n697 B.n696 10.6151
R2278 B.n698 B.n697 10.6151
R2279 B.n699 B.n698 10.6151
R2280 B.n701 B.n699 10.6151
R2281 B.n702 B.n701 10.6151
R2282 B.n703 B.n702 10.6151
R2283 B.n704 B.n703 10.6151
R2284 B.n706 B.n704 10.6151
R2285 B.n707 B.n706 10.6151
R2286 B.n708 B.n707 10.6151
R2287 B.n709 B.n708 10.6151
R2288 B.n711 B.n709 10.6151
R2289 B.n712 B.n711 10.6151
R2290 B.n713 B.n712 10.6151
R2291 B.n714 B.n713 10.6151
R2292 B.n716 B.n714 10.6151
R2293 B.n717 B.n716 10.6151
R2294 B.n718 B.n717 10.6151
R2295 B.n719 B.n718 10.6151
R2296 B.n721 B.n719 10.6151
R2297 B.n722 B.n721 10.6151
R2298 B.n723 B.n722 10.6151
R2299 B.n724 B.n723 10.6151
R2300 B.n726 B.n724 10.6151
R2301 B.n727 B.n726 10.6151
R2302 B.n728 B.n727 10.6151
R2303 B.n729 B.n728 10.6151
R2304 B.n731 B.n729 10.6151
R2305 B.n732 B.n731 10.6151
R2306 B.n733 B.n732 10.6151
R2307 B.n734 B.n733 10.6151
R2308 B.n736 B.n734 10.6151
R2309 B.n737 B.n736 10.6151
R2310 B.n738 B.n737 10.6151
R2311 B.n739 B.n738 10.6151
R2312 B.n741 B.n739 10.6151
R2313 B.n742 B.n741 10.6151
R2314 B.n743 B.n742 10.6151
R2315 B.n744 B.n743 10.6151
R2316 B.n746 B.n744 10.6151
R2317 B.n747 B.n746 10.6151
R2318 B.n748 B.n747 10.6151
R2319 B.n749 B.n748 10.6151
R2320 B.n751 B.n749 10.6151
R2321 B.n752 B.n751 10.6151
R2322 B.n753 B.n752 10.6151
R2323 B.n754 B.n753 10.6151
R2324 B.n756 B.n754 10.6151
R2325 B.n757 B.n756 10.6151
R2326 B.n758 B.n757 10.6151
R2327 B.n759 B.n758 10.6151
R2328 B.n761 B.n759 10.6151
R2329 B.n762 B.n761 10.6151
R2330 B.n763 B.n762 10.6151
R2331 B.n764 B.n763 10.6151
R2332 B.n496 B.n495 10.6151
R2333 B.n495 B.n282 10.6151
R2334 B.n490 B.n282 10.6151
R2335 B.n490 B.n489 10.6151
R2336 B.n489 B.n284 10.6151
R2337 B.n484 B.n284 10.6151
R2338 B.n484 B.n483 10.6151
R2339 B.n483 B.n482 10.6151
R2340 B.n482 B.n286 10.6151
R2341 B.n476 B.n286 10.6151
R2342 B.n476 B.n475 10.6151
R2343 B.n475 B.n474 10.6151
R2344 B.n474 B.n288 10.6151
R2345 B.n468 B.n288 10.6151
R2346 B.n468 B.n467 10.6151
R2347 B.n467 B.n466 10.6151
R2348 B.n466 B.n290 10.6151
R2349 B.n460 B.n290 10.6151
R2350 B.n460 B.n459 10.6151
R2351 B.n459 B.n458 10.6151
R2352 B.n458 B.n292 10.6151
R2353 B.n452 B.n292 10.6151
R2354 B.n452 B.n451 10.6151
R2355 B.n451 B.n450 10.6151
R2356 B.n450 B.n294 10.6151
R2357 B.n444 B.n294 10.6151
R2358 B.n444 B.n443 10.6151
R2359 B.n443 B.n442 10.6151
R2360 B.n442 B.n296 10.6151
R2361 B.n436 B.n296 10.6151
R2362 B.n436 B.n435 10.6151
R2363 B.n435 B.n434 10.6151
R2364 B.n434 B.n298 10.6151
R2365 B.n428 B.n298 10.6151
R2366 B.n428 B.n427 10.6151
R2367 B.n427 B.n426 10.6151
R2368 B.n426 B.n300 10.6151
R2369 B.n420 B.n419 10.6151
R2370 B.n419 B.n418 10.6151
R2371 B.n418 B.n305 10.6151
R2372 B.n412 B.n305 10.6151
R2373 B.n412 B.n411 10.6151
R2374 B.n411 B.n410 10.6151
R2375 B.n410 B.n307 10.6151
R2376 B.n404 B.n307 10.6151
R2377 B.n402 B.n401 10.6151
R2378 B.n401 B.n311 10.6151
R2379 B.n395 B.n311 10.6151
R2380 B.n395 B.n394 10.6151
R2381 B.n394 B.n393 10.6151
R2382 B.n393 B.n313 10.6151
R2383 B.n387 B.n313 10.6151
R2384 B.n387 B.n386 10.6151
R2385 B.n386 B.n385 10.6151
R2386 B.n385 B.n315 10.6151
R2387 B.n379 B.n315 10.6151
R2388 B.n379 B.n378 10.6151
R2389 B.n378 B.n377 10.6151
R2390 B.n377 B.n317 10.6151
R2391 B.n371 B.n317 10.6151
R2392 B.n371 B.n370 10.6151
R2393 B.n370 B.n369 10.6151
R2394 B.n369 B.n319 10.6151
R2395 B.n363 B.n319 10.6151
R2396 B.n363 B.n362 10.6151
R2397 B.n362 B.n361 10.6151
R2398 B.n361 B.n321 10.6151
R2399 B.n355 B.n321 10.6151
R2400 B.n355 B.n354 10.6151
R2401 B.n354 B.n353 10.6151
R2402 B.n353 B.n323 10.6151
R2403 B.n347 B.n323 10.6151
R2404 B.n347 B.n346 10.6151
R2405 B.n346 B.n345 10.6151
R2406 B.n345 B.n325 10.6151
R2407 B.n339 B.n325 10.6151
R2408 B.n339 B.n338 10.6151
R2409 B.n338 B.n337 10.6151
R2410 B.n337 B.n327 10.6151
R2411 B.n331 B.n327 10.6151
R2412 B.n331 B.n330 10.6151
R2413 B.n330 B.n278 10.6151
R2414 B.n497 B.n274 10.6151
R2415 B.n507 B.n274 10.6151
R2416 B.n508 B.n507 10.6151
R2417 B.n509 B.n508 10.6151
R2418 B.n509 B.n266 10.6151
R2419 B.n520 B.n266 10.6151
R2420 B.n521 B.n520 10.6151
R2421 B.n522 B.n521 10.6151
R2422 B.n522 B.n259 10.6151
R2423 B.n532 B.n259 10.6151
R2424 B.n533 B.n532 10.6151
R2425 B.n534 B.n533 10.6151
R2426 B.n534 B.n251 10.6151
R2427 B.n544 B.n251 10.6151
R2428 B.n545 B.n544 10.6151
R2429 B.n546 B.n545 10.6151
R2430 B.n546 B.n243 10.6151
R2431 B.n557 B.n243 10.6151
R2432 B.n558 B.n557 10.6151
R2433 B.n559 B.n558 10.6151
R2434 B.n559 B.n236 10.6151
R2435 B.n569 B.n236 10.6151
R2436 B.n570 B.n569 10.6151
R2437 B.n571 B.n570 10.6151
R2438 B.n571 B.n228 10.6151
R2439 B.n581 B.n228 10.6151
R2440 B.n582 B.n581 10.6151
R2441 B.n583 B.n582 10.6151
R2442 B.n583 B.n220 10.6151
R2443 B.n593 B.n220 10.6151
R2444 B.n594 B.n593 10.6151
R2445 B.n595 B.n594 10.6151
R2446 B.n595 B.n212 10.6151
R2447 B.n605 B.n212 10.6151
R2448 B.n606 B.n605 10.6151
R2449 B.n607 B.n606 10.6151
R2450 B.n607 B.n204 10.6151
R2451 B.n617 B.n204 10.6151
R2452 B.n618 B.n617 10.6151
R2453 B.n619 B.n618 10.6151
R2454 B.n619 B.n196 10.6151
R2455 B.n629 B.n196 10.6151
R2456 B.n630 B.n629 10.6151
R2457 B.n631 B.n630 10.6151
R2458 B.n631 B.n188 10.6151
R2459 B.n641 B.n188 10.6151
R2460 B.n642 B.n641 10.6151
R2461 B.n643 B.n642 10.6151
R2462 B.n643 B.n180 10.6151
R2463 B.n653 B.n180 10.6151
R2464 B.n654 B.n653 10.6151
R2465 B.n655 B.n654 10.6151
R2466 B.n655 B.n172 10.6151
R2467 B.n666 B.n172 10.6151
R2468 B.n667 B.n666 10.6151
R2469 B.n668 B.n667 10.6151
R2470 B.n668 B.n165 10.6151
R2471 B.n679 B.n165 10.6151
R2472 B.n680 B.n679 10.6151
R2473 B.n681 B.n680 10.6151
R2474 B.n681 B.n0 10.6151
R2475 B.n1056 B.n1 10.6151
R2476 B.n1056 B.n1055 10.6151
R2477 B.n1055 B.n1054 10.6151
R2478 B.n1054 B.n10 10.6151
R2479 B.n1048 B.n10 10.6151
R2480 B.n1048 B.n1047 10.6151
R2481 B.n1047 B.n1046 10.6151
R2482 B.n1046 B.n16 10.6151
R2483 B.n1040 B.n16 10.6151
R2484 B.n1040 B.n1039 10.6151
R2485 B.n1039 B.n1038 10.6151
R2486 B.n1038 B.n24 10.6151
R2487 B.n1032 B.n24 10.6151
R2488 B.n1032 B.n1031 10.6151
R2489 B.n1031 B.n1030 10.6151
R2490 B.n1030 B.n31 10.6151
R2491 B.n1024 B.n31 10.6151
R2492 B.n1024 B.n1023 10.6151
R2493 B.n1023 B.n1022 10.6151
R2494 B.n1022 B.n38 10.6151
R2495 B.n1016 B.n38 10.6151
R2496 B.n1016 B.n1015 10.6151
R2497 B.n1015 B.n1014 10.6151
R2498 B.n1014 B.n45 10.6151
R2499 B.n1008 B.n45 10.6151
R2500 B.n1008 B.n1007 10.6151
R2501 B.n1007 B.n1006 10.6151
R2502 B.n1006 B.n52 10.6151
R2503 B.n1000 B.n52 10.6151
R2504 B.n1000 B.n999 10.6151
R2505 B.n999 B.n998 10.6151
R2506 B.n998 B.n59 10.6151
R2507 B.n992 B.n59 10.6151
R2508 B.n992 B.n991 10.6151
R2509 B.n991 B.n990 10.6151
R2510 B.n990 B.n66 10.6151
R2511 B.n984 B.n66 10.6151
R2512 B.n984 B.n983 10.6151
R2513 B.n983 B.n982 10.6151
R2514 B.n982 B.n73 10.6151
R2515 B.n976 B.n73 10.6151
R2516 B.n976 B.n975 10.6151
R2517 B.n975 B.n974 10.6151
R2518 B.n974 B.n79 10.6151
R2519 B.n968 B.n79 10.6151
R2520 B.n968 B.n967 10.6151
R2521 B.n967 B.n966 10.6151
R2522 B.n966 B.n87 10.6151
R2523 B.n960 B.n87 10.6151
R2524 B.n960 B.n959 10.6151
R2525 B.n959 B.n958 10.6151
R2526 B.n958 B.n94 10.6151
R2527 B.n952 B.n94 10.6151
R2528 B.n952 B.n951 10.6151
R2529 B.n951 B.n950 10.6151
R2530 B.n950 B.n100 10.6151
R2531 B.n944 B.n100 10.6151
R2532 B.n944 B.n943 10.6151
R2533 B.n943 B.n942 10.6151
R2534 B.n942 B.n108 10.6151
R2535 B.n936 B.n108 10.6151
R2536 B.t3 B.n222 9.64056
R2537 B.n995 B.t5 9.64056
R2538 B.n615 B.t7 8.26341
R2539 B.n1012 B.t2 8.26341
R2540 B.t23 B.n186 6.88626
R2541 B.t1 B.n29 6.88626
R2542 B.n858 B.n135 6.5566
R2543 B.n843 B.n842 6.5566
R2544 B.n420 B.n304 6.5566
R2545 B.n404 B.n403 6.5566
R2546 B.n670 B.t8 5.50911
R2547 B.n1050 B.t4 5.50911
R2548 B.n862 B.n135 4.05904
R2549 B.n842 B.n841 4.05904
R2550 B.n304 B.n300 4.05904
R2551 B.n403 B.n402 4.05904
R2552 B.n1062 B.n0 2.81026
R2553 B.n1062 B.n1 2.81026
R2554 VP.n27 VP.n26 161.3
R2555 VP.n28 VP.n23 161.3
R2556 VP.n30 VP.n29 161.3
R2557 VP.n31 VP.n22 161.3
R2558 VP.n33 VP.n32 161.3
R2559 VP.n34 VP.n21 161.3
R2560 VP.n36 VP.n35 161.3
R2561 VP.n37 VP.n20 161.3
R2562 VP.n39 VP.n38 161.3
R2563 VP.n40 VP.n19 161.3
R2564 VP.n42 VP.n41 161.3
R2565 VP.n43 VP.n18 161.3
R2566 VP.n45 VP.n44 161.3
R2567 VP.n47 VP.n46 161.3
R2568 VP.n48 VP.n16 161.3
R2569 VP.n50 VP.n49 161.3
R2570 VP.n51 VP.n15 161.3
R2571 VP.n53 VP.n52 161.3
R2572 VP.n54 VP.n14 161.3
R2573 VP.n96 VP.n0 161.3
R2574 VP.n95 VP.n94 161.3
R2575 VP.n93 VP.n1 161.3
R2576 VP.n92 VP.n91 161.3
R2577 VP.n90 VP.n2 161.3
R2578 VP.n89 VP.n88 161.3
R2579 VP.n87 VP.n86 161.3
R2580 VP.n85 VP.n4 161.3
R2581 VP.n84 VP.n83 161.3
R2582 VP.n82 VP.n5 161.3
R2583 VP.n81 VP.n80 161.3
R2584 VP.n79 VP.n6 161.3
R2585 VP.n78 VP.n77 161.3
R2586 VP.n76 VP.n7 161.3
R2587 VP.n75 VP.n74 161.3
R2588 VP.n73 VP.n8 161.3
R2589 VP.n72 VP.n71 161.3
R2590 VP.n70 VP.n9 161.3
R2591 VP.n69 VP.n68 161.3
R2592 VP.n66 VP.n10 161.3
R2593 VP.n65 VP.n64 161.3
R2594 VP.n63 VP.n11 161.3
R2595 VP.n62 VP.n61 161.3
R2596 VP.n60 VP.n12 161.3
R2597 VP.n59 VP.n58 161.3
R2598 VP.n24 VP.t4 126.767
R2599 VP.n57 VP.n13 104.022
R2600 VP.n98 VP.n97 104.022
R2601 VP.n56 VP.n55 104.022
R2602 VP.n78 VP.t8 94.1136
R2603 VP.n13 VP.t6 94.1136
R2604 VP.n67 VP.t9 94.1136
R2605 VP.n3 VP.t3 94.1136
R2606 VP.n97 VP.t2 94.1136
R2607 VP.n36 VP.t7 94.1136
R2608 VP.n55 VP.t5 94.1136
R2609 VP.n17 VP.t1 94.1136
R2610 VP.n25 VP.t0 94.1136
R2611 VP.n25 VP.n24 69.6937
R2612 VP.n57 VP.n56 52.8974
R2613 VP.n61 VP.n11 50.7491
R2614 VP.n91 VP.n1 50.7491
R2615 VP.n49 VP.n15 50.7491
R2616 VP.n73 VP.n72 43.9677
R2617 VP.n84 VP.n5 43.9677
R2618 VP.n42 VP.n19 43.9677
R2619 VP.n31 VP.n30 43.9677
R2620 VP.n74 VP.n73 37.1863
R2621 VP.n80 VP.n5 37.1863
R2622 VP.n38 VP.n19 37.1863
R2623 VP.n32 VP.n31 37.1863
R2624 VP.n65 VP.n11 30.405
R2625 VP.n91 VP.n90 30.405
R2626 VP.n49 VP.n48 30.405
R2627 VP.n60 VP.n59 24.5923
R2628 VP.n61 VP.n60 24.5923
R2629 VP.n66 VP.n65 24.5923
R2630 VP.n68 VP.n9 24.5923
R2631 VP.n72 VP.n9 24.5923
R2632 VP.n74 VP.n7 24.5923
R2633 VP.n78 VP.n7 24.5923
R2634 VP.n79 VP.n78 24.5923
R2635 VP.n80 VP.n79 24.5923
R2636 VP.n85 VP.n84 24.5923
R2637 VP.n86 VP.n85 24.5923
R2638 VP.n90 VP.n89 24.5923
R2639 VP.n95 VP.n1 24.5923
R2640 VP.n96 VP.n95 24.5923
R2641 VP.n53 VP.n15 24.5923
R2642 VP.n54 VP.n53 24.5923
R2643 VP.n43 VP.n42 24.5923
R2644 VP.n44 VP.n43 24.5923
R2645 VP.n48 VP.n47 24.5923
R2646 VP.n32 VP.n21 24.5923
R2647 VP.n36 VP.n21 24.5923
R2648 VP.n37 VP.n36 24.5923
R2649 VP.n38 VP.n37 24.5923
R2650 VP.n26 VP.n23 24.5923
R2651 VP.n30 VP.n23 24.5923
R2652 VP.n67 VP.n66 21.1495
R2653 VP.n89 VP.n3 21.1495
R2654 VP.n47 VP.n17 21.1495
R2655 VP.n27 VP.n24 7.0306
R2656 VP.n59 VP.n13 6.88621
R2657 VP.n97 VP.n96 6.88621
R2658 VP.n55 VP.n54 6.88621
R2659 VP.n68 VP.n67 3.44336
R2660 VP.n86 VP.n3 3.44336
R2661 VP.n44 VP.n17 3.44336
R2662 VP.n26 VP.n25 3.44336
R2663 VP.n56 VP.n14 0.278335
R2664 VP.n58 VP.n57 0.278335
R2665 VP.n98 VP.n0 0.278335
R2666 VP.n28 VP.n27 0.189894
R2667 VP.n29 VP.n28 0.189894
R2668 VP.n29 VP.n22 0.189894
R2669 VP.n33 VP.n22 0.189894
R2670 VP.n34 VP.n33 0.189894
R2671 VP.n35 VP.n34 0.189894
R2672 VP.n35 VP.n20 0.189894
R2673 VP.n39 VP.n20 0.189894
R2674 VP.n40 VP.n39 0.189894
R2675 VP.n41 VP.n40 0.189894
R2676 VP.n41 VP.n18 0.189894
R2677 VP.n45 VP.n18 0.189894
R2678 VP.n46 VP.n45 0.189894
R2679 VP.n46 VP.n16 0.189894
R2680 VP.n50 VP.n16 0.189894
R2681 VP.n51 VP.n50 0.189894
R2682 VP.n52 VP.n51 0.189894
R2683 VP.n52 VP.n14 0.189894
R2684 VP.n58 VP.n12 0.189894
R2685 VP.n62 VP.n12 0.189894
R2686 VP.n63 VP.n62 0.189894
R2687 VP.n64 VP.n63 0.189894
R2688 VP.n64 VP.n10 0.189894
R2689 VP.n69 VP.n10 0.189894
R2690 VP.n70 VP.n69 0.189894
R2691 VP.n71 VP.n70 0.189894
R2692 VP.n71 VP.n8 0.189894
R2693 VP.n75 VP.n8 0.189894
R2694 VP.n76 VP.n75 0.189894
R2695 VP.n77 VP.n76 0.189894
R2696 VP.n77 VP.n6 0.189894
R2697 VP.n81 VP.n6 0.189894
R2698 VP.n82 VP.n81 0.189894
R2699 VP.n83 VP.n82 0.189894
R2700 VP.n83 VP.n4 0.189894
R2701 VP.n87 VP.n4 0.189894
R2702 VP.n88 VP.n87 0.189894
R2703 VP.n88 VP.n2 0.189894
R2704 VP.n92 VP.n2 0.189894
R2705 VP.n93 VP.n92 0.189894
R2706 VP.n94 VP.n93 0.189894
R2707 VP.n94 VP.n0 0.189894
R2708 VP VP.n98 0.153485
R2709 VDD1.n52 VDD1.n0 289.615
R2710 VDD1.n111 VDD1.n59 289.615
R2711 VDD1.n53 VDD1.n52 185
R2712 VDD1.n51 VDD1.n50 185
R2713 VDD1.n4 VDD1.n3 185
R2714 VDD1.n45 VDD1.n44 185
R2715 VDD1.n43 VDD1.n42 185
R2716 VDD1.n41 VDD1.n7 185
R2717 VDD1.n11 VDD1.n8 185
R2718 VDD1.n36 VDD1.n35 185
R2719 VDD1.n34 VDD1.n33 185
R2720 VDD1.n13 VDD1.n12 185
R2721 VDD1.n28 VDD1.n27 185
R2722 VDD1.n26 VDD1.n25 185
R2723 VDD1.n17 VDD1.n16 185
R2724 VDD1.n20 VDD1.n19 185
R2725 VDD1.n78 VDD1.n77 185
R2726 VDD1.n75 VDD1.n74 185
R2727 VDD1.n84 VDD1.n83 185
R2728 VDD1.n86 VDD1.n85 185
R2729 VDD1.n71 VDD1.n70 185
R2730 VDD1.n92 VDD1.n91 185
R2731 VDD1.n95 VDD1.n94 185
R2732 VDD1.n93 VDD1.n67 185
R2733 VDD1.n100 VDD1.n66 185
R2734 VDD1.n102 VDD1.n101 185
R2735 VDD1.n104 VDD1.n103 185
R2736 VDD1.n63 VDD1.n62 185
R2737 VDD1.n110 VDD1.n109 185
R2738 VDD1.n112 VDD1.n111 185
R2739 VDD1.t5 VDD1.n18 149.524
R2740 VDD1.t3 VDD1.n76 149.524
R2741 VDD1.n52 VDD1.n51 104.615
R2742 VDD1.n51 VDD1.n3 104.615
R2743 VDD1.n44 VDD1.n3 104.615
R2744 VDD1.n44 VDD1.n43 104.615
R2745 VDD1.n43 VDD1.n7 104.615
R2746 VDD1.n11 VDD1.n7 104.615
R2747 VDD1.n35 VDD1.n11 104.615
R2748 VDD1.n35 VDD1.n34 104.615
R2749 VDD1.n34 VDD1.n12 104.615
R2750 VDD1.n27 VDD1.n12 104.615
R2751 VDD1.n27 VDD1.n26 104.615
R2752 VDD1.n26 VDD1.n16 104.615
R2753 VDD1.n19 VDD1.n16 104.615
R2754 VDD1.n77 VDD1.n74 104.615
R2755 VDD1.n84 VDD1.n74 104.615
R2756 VDD1.n85 VDD1.n84 104.615
R2757 VDD1.n85 VDD1.n70 104.615
R2758 VDD1.n92 VDD1.n70 104.615
R2759 VDD1.n94 VDD1.n92 104.615
R2760 VDD1.n94 VDD1.n93 104.615
R2761 VDD1.n93 VDD1.n66 104.615
R2762 VDD1.n102 VDD1.n66 104.615
R2763 VDD1.n103 VDD1.n102 104.615
R2764 VDD1.n103 VDD1.n62 104.615
R2765 VDD1.n110 VDD1.n62 104.615
R2766 VDD1.n111 VDD1.n110 104.615
R2767 VDD1.n119 VDD1.n118 64.6576
R2768 VDD1.n58 VDD1.n57 62.7282
R2769 VDD1.n121 VDD1.n120 62.728
R2770 VDD1.n117 VDD1.n116 62.728
R2771 VDD1.n19 VDD1.t5 52.3082
R2772 VDD1.n77 VDD1.t3 52.3082
R2773 VDD1.n58 VDD1.n56 51.8986
R2774 VDD1.n117 VDD1.n115 51.8986
R2775 VDD1.n121 VDD1.n119 47.4168
R2776 VDD1.n42 VDD1.n41 13.1884
R2777 VDD1.n101 VDD1.n100 13.1884
R2778 VDD1.n45 VDD1.n6 12.8005
R2779 VDD1.n40 VDD1.n8 12.8005
R2780 VDD1.n99 VDD1.n67 12.8005
R2781 VDD1.n104 VDD1.n65 12.8005
R2782 VDD1.n46 VDD1.n4 12.0247
R2783 VDD1.n37 VDD1.n36 12.0247
R2784 VDD1.n96 VDD1.n95 12.0247
R2785 VDD1.n105 VDD1.n63 12.0247
R2786 VDD1.n50 VDD1.n49 11.249
R2787 VDD1.n33 VDD1.n10 11.249
R2788 VDD1.n91 VDD1.n69 11.249
R2789 VDD1.n109 VDD1.n108 11.249
R2790 VDD1.n53 VDD1.n2 10.4732
R2791 VDD1.n32 VDD1.n13 10.4732
R2792 VDD1.n90 VDD1.n71 10.4732
R2793 VDD1.n112 VDD1.n61 10.4732
R2794 VDD1.n20 VDD1.n18 10.2747
R2795 VDD1.n78 VDD1.n76 10.2747
R2796 VDD1.n54 VDD1.n0 9.69747
R2797 VDD1.n29 VDD1.n28 9.69747
R2798 VDD1.n87 VDD1.n86 9.69747
R2799 VDD1.n113 VDD1.n59 9.69747
R2800 VDD1.n56 VDD1.n55 9.45567
R2801 VDD1.n115 VDD1.n114 9.45567
R2802 VDD1.n22 VDD1.n21 9.3005
R2803 VDD1.n24 VDD1.n23 9.3005
R2804 VDD1.n15 VDD1.n14 9.3005
R2805 VDD1.n30 VDD1.n29 9.3005
R2806 VDD1.n32 VDD1.n31 9.3005
R2807 VDD1.n10 VDD1.n9 9.3005
R2808 VDD1.n38 VDD1.n37 9.3005
R2809 VDD1.n40 VDD1.n39 9.3005
R2810 VDD1.n55 VDD1.n54 9.3005
R2811 VDD1.n2 VDD1.n1 9.3005
R2812 VDD1.n49 VDD1.n48 9.3005
R2813 VDD1.n47 VDD1.n46 9.3005
R2814 VDD1.n6 VDD1.n5 9.3005
R2815 VDD1.n114 VDD1.n113 9.3005
R2816 VDD1.n61 VDD1.n60 9.3005
R2817 VDD1.n108 VDD1.n107 9.3005
R2818 VDD1.n106 VDD1.n105 9.3005
R2819 VDD1.n65 VDD1.n64 9.3005
R2820 VDD1.n80 VDD1.n79 9.3005
R2821 VDD1.n82 VDD1.n81 9.3005
R2822 VDD1.n73 VDD1.n72 9.3005
R2823 VDD1.n88 VDD1.n87 9.3005
R2824 VDD1.n90 VDD1.n89 9.3005
R2825 VDD1.n69 VDD1.n68 9.3005
R2826 VDD1.n97 VDD1.n96 9.3005
R2827 VDD1.n99 VDD1.n98 9.3005
R2828 VDD1.n25 VDD1.n15 8.92171
R2829 VDD1.n83 VDD1.n73 8.92171
R2830 VDD1.n24 VDD1.n17 8.14595
R2831 VDD1.n82 VDD1.n75 8.14595
R2832 VDD1.n21 VDD1.n20 7.3702
R2833 VDD1.n79 VDD1.n78 7.3702
R2834 VDD1.n21 VDD1.n17 5.81868
R2835 VDD1.n79 VDD1.n75 5.81868
R2836 VDD1.n25 VDD1.n24 5.04292
R2837 VDD1.n83 VDD1.n82 5.04292
R2838 VDD1.n56 VDD1.n0 4.26717
R2839 VDD1.n28 VDD1.n15 4.26717
R2840 VDD1.n86 VDD1.n73 4.26717
R2841 VDD1.n115 VDD1.n59 4.26717
R2842 VDD1.n54 VDD1.n53 3.49141
R2843 VDD1.n29 VDD1.n13 3.49141
R2844 VDD1.n87 VDD1.n71 3.49141
R2845 VDD1.n113 VDD1.n112 3.49141
R2846 VDD1.n22 VDD1.n18 2.84303
R2847 VDD1.n80 VDD1.n76 2.84303
R2848 VDD1.n50 VDD1.n2 2.71565
R2849 VDD1.n33 VDD1.n32 2.71565
R2850 VDD1.n91 VDD1.n90 2.71565
R2851 VDD1.n109 VDD1.n61 2.71565
R2852 VDD1.n49 VDD1.n4 1.93989
R2853 VDD1.n36 VDD1.n10 1.93989
R2854 VDD1.n95 VDD1.n69 1.93989
R2855 VDD1.n108 VDD1.n63 1.93989
R2856 VDD1 VDD1.n121 1.92722
R2857 VDD1.n120 VDD1.t8 1.85097
R2858 VDD1.n120 VDD1.t4 1.85097
R2859 VDD1.n57 VDD1.t9 1.85097
R2860 VDD1.n57 VDD1.t2 1.85097
R2861 VDD1.n118 VDD1.t6 1.85097
R2862 VDD1.n118 VDD1.t7 1.85097
R2863 VDD1.n116 VDD1.t0 1.85097
R2864 VDD1.n116 VDD1.t1 1.85097
R2865 VDD1.n46 VDD1.n45 1.16414
R2866 VDD1.n37 VDD1.n8 1.16414
R2867 VDD1.n96 VDD1.n67 1.16414
R2868 VDD1.n105 VDD1.n104 1.16414
R2869 VDD1 VDD1.n58 0.720328
R2870 VDD1.n119 VDD1.n117 0.606792
R2871 VDD1.n42 VDD1.n6 0.388379
R2872 VDD1.n41 VDD1.n40 0.388379
R2873 VDD1.n100 VDD1.n99 0.388379
R2874 VDD1.n101 VDD1.n65 0.388379
R2875 VDD1.n55 VDD1.n1 0.155672
R2876 VDD1.n48 VDD1.n1 0.155672
R2877 VDD1.n48 VDD1.n47 0.155672
R2878 VDD1.n47 VDD1.n5 0.155672
R2879 VDD1.n39 VDD1.n5 0.155672
R2880 VDD1.n39 VDD1.n38 0.155672
R2881 VDD1.n38 VDD1.n9 0.155672
R2882 VDD1.n31 VDD1.n9 0.155672
R2883 VDD1.n31 VDD1.n30 0.155672
R2884 VDD1.n30 VDD1.n14 0.155672
R2885 VDD1.n23 VDD1.n14 0.155672
R2886 VDD1.n23 VDD1.n22 0.155672
R2887 VDD1.n81 VDD1.n80 0.155672
R2888 VDD1.n81 VDD1.n72 0.155672
R2889 VDD1.n88 VDD1.n72 0.155672
R2890 VDD1.n89 VDD1.n88 0.155672
R2891 VDD1.n89 VDD1.n68 0.155672
R2892 VDD1.n97 VDD1.n68 0.155672
R2893 VDD1.n98 VDD1.n97 0.155672
R2894 VDD1.n98 VDD1.n64 0.155672
R2895 VDD1.n106 VDD1.n64 0.155672
R2896 VDD1.n107 VDD1.n106 0.155672
R2897 VDD1.n107 VDD1.n60 0.155672
R2898 VDD1.n114 VDD1.n60 0.155672
C0 VP VTAIL 10.443f
C1 VP VDD2 0.601479f
C2 VP VDD1 10.1144f
C3 VTAIL VDD2 9.89599f
C4 VTAIL VDD1 9.84367f
C5 VDD1 VDD2 2.26406f
C6 VP VN 8.35572f
C7 VN VTAIL 10.4287f
C8 VN VDD2 9.67039f
C9 VN VDD1 0.153821f
C10 VDD2 B 7.161858f
C11 VDD1 B 7.116049f
C12 VTAIL B 7.789729f
C13 VN B 18.68991f
C14 VP B 17.244623f
C15 VDD1.n0 B 0.034048f
C16 VDD1.n1 B 0.024942f
C17 VDD1.n2 B 0.013403f
C18 VDD1.n3 B 0.031679f
C19 VDD1.n4 B 0.014191f
C20 VDD1.n5 B 0.024942f
C21 VDD1.n6 B 0.013403f
C22 VDD1.n7 B 0.031679f
C23 VDD1.n8 B 0.014191f
C24 VDD1.n9 B 0.024942f
C25 VDD1.n10 B 0.013403f
C26 VDD1.n11 B 0.031679f
C27 VDD1.n12 B 0.031679f
C28 VDD1.n13 B 0.014191f
C29 VDD1.n14 B 0.024942f
C30 VDD1.n15 B 0.013403f
C31 VDD1.n16 B 0.031679f
C32 VDD1.n17 B 0.014191f
C33 VDD1.n18 B 0.167381f
C34 VDD1.t5 B 0.05333f
C35 VDD1.n19 B 0.023759f
C36 VDD1.n20 B 0.022395f
C37 VDD1.n21 B 0.013403f
C38 VDD1.n22 B 1.11405f
C39 VDD1.n23 B 0.024942f
C40 VDD1.n24 B 0.013403f
C41 VDD1.n25 B 0.014191f
C42 VDD1.n26 B 0.031679f
C43 VDD1.n27 B 0.031679f
C44 VDD1.n28 B 0.014191f
C45 VDD1.n29 B 0.013403f
C46 VDD1.n30 B 0.024942f
C47 VDD1.n31 B 0.024942f
C48 VDD1.n32 B 0.013403f
C49 VDD1.n33 B 0.014191f
C50 VDD1.n34 B 0.031679f
C51 VDD1.n35 B 0.031679f
C52 VDD1.n36 B 0.014191f
C53 VDD1.n37 B 0.013403f
C54 VDD1.n38 B 0.024942f
C55 VDD1.n39 B 0.024942f
C56 VDD1.n40 B 0.013403f
C57 VDD1.n41 B 0.013797f
C58 VDD1.n42 B 0.013797f
C59 VDD1.n43 B 0.031679f
C60 VDD1.n44 B 0.031679f
C61 VDD1.n45 B 0.014191f
C62 VDD1.n46 B 0.013403f
C63 VDD1.n47 B 0.024942f
C64 VDD1.n48 B 0.024942f
C65 VDD1.n49 B 0.013403f
C66 VDD1.n50 B 0.014191f
C67 VDD1.n51 B 0.031679f
C68 VDD1.n52 B 0.066794f
C69 VDD1.n53 B 0.014191f
C70 VDD1.n54 B 0.013403f
C71 VDD1.n55 B 0.058333f
C72 VDD1.n56 B 0.067743f
C73 VDD1.t9 B 0.210895f
C74 VDD1.t2 B 0.210895f
C75 VDD1.n57 B 1.86589f
C76 VDD1.n58 B 0.722618f
C77 VDD1.n59 B 0.034048f
C78 VDD1.n60 B 0.024942f
C79 VDD1.n61 B 0.013403f
C80 VDD1.n62 B 0.031679f
C81 VDD1.n63 B 0.014191f
C82 VDD1.n64 B 0.024942f
C83 VDD1.n65 B 0.013403f
C84 VDD1.n66 B 0.031679f
C85 VDD1.n67 B 0.014191f
C86 VDD1.n68 B 0.024942f
C87 VDD1.n69 B 0.013403f
C88 VDD1.n70 B 0.031679f
C89 VDD1.n71 B 0.014191f
C90 VDD1.n72 B 0.024942f
C91 VDD1.n73 B 0.013403f
C92 VDD1.n74 B 0.031679f
C93 VDD1.n75 B 0.014191f
C94 VDD1.n76 B 0.167381f
C95 VDD1.t3 B 0.05333f
C96 VDD1.n77 B 0.023759f
C97 VDD1.n78 B 0.022395f
C98 VDD1.n79 B 0.013403f
C99 VDD1.n80 B 1.11405f
C100 VDD1.n81 B 0.024942f
C101 VDD1.n82 B 0.013403f
C102 VDD1.n83 B 0.014191f
C103 VDD1.n84 B 0.031679f
C104 VDD1.n85 B 0.031679f
C105 VDD1.n86 B 0.014191f
C106 VDD1.n87 B 0.013403f
C107 VDD1.n88 B 0.024942f
C108 VDD1.n89 B 0.024942f
C109 VDD1.n90 B 0.013403f
C110 VDD1.n91 B 0.014191f
C111 VDD1.n92 B 0.031679f
C112 VDD1.n93 B 0.031679f
C113 VDD1.n94 B 0.031679f
C114 VDD1.n95 B 0.014191f
C115 VDD1.n96 B 0.013403f
C116 VDD1.n97 B 0.024942f
C117 VDD1.n98 B 0.024942f
C118 VDD1.n99 B 0.013403f
C119 VDD1.n100 B 0.013797f
C120 VDD1.n101 B 0.013797f
C121 VDD1.n102 B 0.031679f
C122 VDD1.n103 B 0.031679f
C123 VDD1.n104 B 0.014191f
C124 VDD1.n105 B 0.013403f
C125 VDD1.n106 B 0.024942f
C126 VDD1.n107 B 0.024942f
C127 VDD1.n108 B 0.013403f
C128 VDD1.n109 B 0.014191f
C129 VDD1.n110 B 0.031679f
C130 VDD1.n111 B 0.066794f
C131 VDD1.n112 B 0.014191f
C132 VDD1.n113 B 0.013403f
C133 VDD1.n114 B 0.058333f
C134 VDD1.n115 B 0.067743f
C135 VDD1.t0 B 0.210895f
C136 VDD1.t1 B 0.210895f
C137 VDD1.n116 B 1.86589f
C138 VDD1.n117 B 0.714455f
C139 VDD1.t6 B 0.210895f
C140 VDD1.t7 B 0.210895f
C141 VDD1.n118 B 1.88327f
C142 VDD1.n119 B 3.01809f
C143 VDD1.t8 B 0.210895f
C144 VDD1.t4 B 0.210895f
C145 VDD1.n120 B 1.86589f
C146 VDD1.n121 B 3.1235f
C147 VP.n0 B 0.028228f
C148 VP.t2 B 1.70445f
C149 VP.n1 B 0.038898f
C150 VP.n2 B 0.021412f
C151 VP.t3 B 1.70445f
C152 VP.n3 B 0.60602f
C153 VP.n4 B 0.021412f
C154 VP.n5 B 0.01763f
C155 VP.n6 B 0.021412f
C156 VP.t8 B 1.70445f
C157 VP.n7 B 0.039706f
C158 VP.n8 B 0.021412f
C159 VP.n9 B 0.039706f
C160 VP.n10 B 0.021412f
C161 VP.t9 B 1.70445f
C162 VP.n11 B 0.020505f
C163 VP.n12 B 0.021412f
C164 VP.t6 B 1.70445f
C165 VP.n13 B 0.67768f
C166 VP.n14 B 0.028228f
C167 VP.t5 B 1.70445f
C168 VP.n15 B 0.038898f
C169 VP.n16 B 0.021412f
C170 VP.t1 B 1.70445f
C171 VP.n17 B 0.60602f
C172 VP.n18 B 0.021412f
C173 VP.n19 B 0.01763f
C174 VP.n20 B 0.021412f
C175 VP.t7 B 1.70445f
C176 VP.n21 B 0.039706f
C177 VP.n22 B 0.021412f
C178 VP.n23 B 0.039706f
C179 VP.t4 B 1.89545f
C180 VP.n24 B 0.645903f
C181 VP.t0 B 1.70445f
C182 VP.n25 B 0.663225f
C183 VP.n26 B 0.022849f
C184 VP.n27 B 0.21001f
C185 VP.n28 B 0.021412f
C186 VP.n29 B 0.021412f
C187 VP.n30 B 0.041434f
C188 VP.n31 B 0.01763f
C189 VP.n32 B 0.042893f
C190 VP.n33 B 0.021412f
C191 VP.n34 B 0.021412f
C192 VP.n35 B 0.021412f
C193 VP.n36 B 0.626124f
C194 VP.n37 B 0.039706f
C195 VP.n38 B 0.042893f
C196 VP.n39 B 0.021412f
C197 VP.n40 B 0.021412f
C198 VP.n41 B 0.021412f
C199 VP.n42 B 0.041434f
C200 VP.n43 B 0.039706f
C201 VP.n44 B 0.022849f
C202 VP.n45 B 0.021412f
C203 VP.n46 B 0.021412f
C204 VP.n47 B 0.036962f
C205 VP.n48 B 0.042554f
C206 VP.n49 B 0.020505f
C207 VP.n50 B 0.021412f
C208 VP.n51 B 0.021412f
C209 VP.n52 B 0.021412f
C210 VP.n53 B 0.039706f
C211 VP.n54 B 0.025593f
C212 VP.n55 B 0.67768f
C213 VP.n56 B 1.29562f
C214 VP.n57 B 1.31021f
C215 VP.n58 B 0.028228f
C216 VP.n59 B 0.025593f
C217 VP.n60 B 0.039706f
C218 VP.n61 B 0.038898f
C219 VP.n62 B 0.021412f
C220 VP.n63 B 0.021412f
C221 VP.n64 B 0.021412f
C222 VP.n65 B 0.042554f
C223 VP.n66 B 0.036962f
C224 VP.n67 B 0.60602f
C225 VP.n68 B 0.022849f
C226 VP.n69 B 0.021412f
C227 VP.n70 B 0.021412f
C228 VP.n71 B 0.021412f
C229 VP.n72 B 0.041434f
C230 VP.n73 B 0.01763f
C231 VP.n74 B 0.042893f
C232 VP.n75 B 0.021412f
C233 VP.n76 B 0.021412f
C234 VP.n77 B 0.021412f
C235 VP.n78 B 0.626124f
C236 VP.n79 B 0.039706f
C237 VP.n80 B 0.042893f
C238 VP.n81 B 0.021412f
C239 VP.n82 B 0.021412f
C240 VP.n83 B 0.021412f
C241 VP.n84 B 0.041434f
C242 VP.n85 B 0.039706f
C243 VP.n86 B 0.022849f
C244 VP.n87 B 0.021412f
C245 VP.n88 B 0.021412f
C246 VP.n89 B 0.036962f
C247 VP.n90 B 0.042554f
C248 VP.n91 B 0.020505f
C249 VP.n92 B 0.021412f
C250 VP.n93 B 0.021412f
C251 VP.n94 B 0.021412f
C252 VP.n95 B 0.039706f
C253 VP.n96 B 0.025593f
C254 VP.n97 B 0.67768f
C255 VP.n98 B 0.037499f
C256 VDD2.n0 B 0.033728f
C257 VDD2.n1 B 0.024707f
C258 VDD2.n2 B 0.013277f
C259 VDD2.n3 B 0.031381f
C260 VDD2.n4 B 0.014058f
C261 VDD2.n5 B 0.024707f
C262 VDD2.n6 B 0.013277f
C263 VDD2.n7 B 0.031381f
C264 VDD2.n8 B 0.014058f
C265 VDD2.n9 B 0.024707f
C266 VDD2.n10 B 0.013277f
C267 VDD2.n11 B 0.031381f
C268 VDD2.n12 B 0.014058f
C269 VDD2.n13 B 0.024707f
C270 VDD2.n14 B 0.013277f
C271 VDD2.n15 B 0.031381f
C272 VDD2.n16 B 0.014058f
C273 VDD2.n17 B 0.165807f
C274 VDD2.t2 B 0.052828f
C275 VDD2.n18 B 0.023536f
C276 VDD2.n19 B 0.022184f
C277 VDD2.n20 B 0.013277f
C278 VDD2.n21 B 1.10358f
C279 VDD2.n22 B 0.024707f
C280 VDD2.n23 B 0.013277f
C281 VDD2.n24 B 0.014058f
C282 VDD2.n25 B 0.031381f
C283 VDD2.n26 B 0.031381f
C284 VDD2.n27 B 0.014058f
C285 VDD2.n28 B 0.013277f
C286 VDD2.n29 B 0.024707f
C287 VDD2.n30 B 0.024707f
C288 VDD2.n31 B 0.013277f
C289 VDD2.n32 B 0.014058f
C290 VDD2.n33 B 0.031381f
C291 VDD2.n34 B 0.031381f
C292 VDD2.n35 B 0.031381f
C293 VDD2.n36 B 0.014058f
C294 VDD2.n37 B 0.013277f
C295 VDD2.n38 B 0.024707f
C296 VDD2.n39 B 0.024707f
C297 VDD2.n40 B 0.013277f
C298 VDD2.n41 B 0.013667f
C299 VDD2.n42 B 0.013667f
C300 VDD2.n43 B 0.031381f
C301 VDD2.n44 B 0.031381f
C302 VDD2.n45 B 0.014058f
C303 VDD2.n46 B 0.013277f
C304 VDD2.n47 B 0.024707f
C305 VDD2.n48 B 0.024707f
C306 VDD2.n49 B 0.013277f
C307 VDD2.n50 B 0.014058f
C308 VDD2.n51 B 0.031381f
C309 VDD2.n52 B 0.066166f
C310 VDD2.n53 B 0.014058f
C311 VDD2.n54 B 0.013277f
C312 VDD2.n55 B 0.057785f
C313 VDD2.n56 B 0.067106f
C314 VDD2.t1 B 0.208912f
C315 VDD2.t0 B 0.208912f
C316 VDD2.n57 B 1.84834f
C317 VDD2.n58 B 0.707737f
C318 VDD2.t5 B 0.208912f
C319 VDD2.t6 B 0.208912f
C320 VDD2.n59 B 1.86556f
C321 VDD2.n60 B 2.86331f
C322 VDD2.n61 B 0.033728f
C323 VDD2.n62 B 0.024707f
C324 VDD2.n63 B 0.013277f
C325 VDD2.n64 B 0.031381f
C326 VDD2.n65 B 0.014058f
C327 VDD2.n66 B 0.024707f
C328 VDD2.n67 B 0.013277f
C329 VDD2.n68 B 0.031381f
C330 VDD2.n69 B 0.014058f
C331 VDD2.n70 B 0.024707f
C332 VDD2.n71 B 0.013277f
C333 VDD2.n72 B 0.031381f
C334 VDD2.n73 B 0.031381f
C335 VDD2.n74 B 0.014058f
C336 VDD2.n75 B 0.024707f
C337 VDD2.n76 B 0.013277f
C338 VDD2.n77 B 0.031381f
C339 VDD2.n78 B 0.014058f
C340 VDD2.n79 B 0.165807f
C341 VDD2.t8 B 0.052828f
C342 VDD2.n80 B 0.023536f
C343 VDD2.n81 B 0.022184f
C344 VDD2.n82 B 0.013277f
C345 VDD2.n83 B 1.10358f
C346 VDD2.n84 B 0.024707f
C347 VDD2.n85 B 0.013277f
C348 VDD2.n86 B 0.014058f
C349 VDD2.n87 B 0.031381f
C350 VDD2.n88 B 0.031381f
C351 VDD2.n89 B 0.014058f
C352 VDD2.n90 B 0.013277f
C353 VDD2.n91 B 0.024707f
C354 VDD2.n92 B 0.024707f
C355 VDD2.n93 B 0.013277f
C356 VDD2.n94 B 0.014058f
C357 VDD2.n95 B 0.031381f
C358 VDD2.n96 B 0.031381f
C359 VDD2.n97 B 0.014058f
C360 VDD2.n98 B 0.013277f
C361 VDD2.n99 B 0.024707f
C362 VDD2.n100 B 0.024707f
C363 VDD2.n101 B 0.013277f
C364 VDD2.n102 B 0.013667f
C365 VDD2.n103 B 0.013667f
C366 VDD2.n104 B 0.031381f
C367 VDD2.n105 B 0.031381f
C368 VDD2.n106 B 0.014058f
C369 VDD2.n107 B 0.013277f
C370 VDD2.n108 B 0.024707f
C371 VDD2.n109 B 0.024707f
C372 VDD2.n110 B 0.013277f
C373 VDD2.n111 B 0.014058f
C374 VDD2.n112 B 0.031381f
C375 VDD2.n113 B 0.066166f
C376 VDD2.n114 B 0.014058f
C377 VDD2.n115 B 0.013277f
C378 VDD2.n116 B 0.057785f
C379 VDD2.n117 B 0.053916f
C380 VDD2.n118 B 2.81154f
C381 VDD2.t3 B 0.208912f
C382 VDD2.t9 B 0.208912f
C383 VDD2.n119 B 1.84835f
C384 VDD2.n120 B 0.470353f
C385 VDD2.t7 B 0.208912f
C386 VDD2.t4 B 0.208912f
C387 VDD2.n121 B 1.86552f
C388 VTAIL.t10 B 0.215218f
C389 VTAIL.t13 B 0.215218f
C390 VTAIL.n0 B 1.83039f
C391 VTAIL.n1 B 0.562247f
C392 VTAIL.n2 B 0.034746f
C393 VTAIL.n3 B 0.025453f
C394 VTAIL.n4 B 0.013677f
C395 VTAIL.n5 B 0.032328f
C396 VTAIL.n6 B 0.014482f
C397 VTAIL.n7 B 0.025453f
C398 VTAIL.n8 B 0.013677f
C399 VTAIL.n9 B 0.032328f
C400 VTAIL.n10 B 0.014482f
C401 VTAIL.n11 B 0.025453f
C402 VTAIL.n12 B 0.013677f
C403 VTAIL.n13 B 0.032328f
C404 VTAIL.n14 B 0.014482f
C405 VTAIL.n15 B 0.025453f
C406 VTAIL.n16 B 0.013677f
C407 VTAIL.n17 B 0.032328f
C408 VTAIL.n18 B 0.014482f
C409 VTAIL.n19 B 0.170812f
C410 VTAIL.t8 B 0.054423f
C411 VTAIL.n20 B 0.024246f
C412 VTAIL.n21 B 0.022854f
C413 VTAIL.n22 B 0.013677f
C414 VTAIL.n23 B 1.13689f
C415 VTAIL.n24 B 0.025453f
C416 VTAIL.n25 B 0.013677f
C417 VTAIL.n26 B 0.014482f
C418 VTAIL.n27 B 0.032328f
C419 VTAIL.n28 B 0.032328f
C420 VTAIL.n29 B 0.014482f
C421 VTAIL.n30 B 0.013677f
C422 VTAIL.n31 B 0.025453f
C423 VTAIL.n32 B 0.025453f
C424 VTAIL.n33 B 0.013677f
C425 VTAIL.n34 B 0.014482f
C426 VTAIL.n35 B 0.032328f
C427 VTAIL.n36 B 0.032328f
C428 VTAIL.n37 B 0.032328f
C429 VTAIL.n38 B 0.014482f
C430 VTAIL.n39 B 0.013677f
C431 VTAIL.n40 B 0.025453f
C432 VTAIL.n41 B 0.025453f
C433 VTAIL.n42 B 0.013677f
C434 VTAIL.n43 B 0.01408f
C435 VTAIL.n44 B 0.01408f
C436 VTAIL.n45 B 0.032328f
C437 VTAIL.n46 B 0.032328f
C438 VTAIL.n47 B 0.014482f
C439 VTAIL.n48 B 0.013677f
C440 VTAIL.n49 B 0.025453f
C441 VTAIL.n50 B 0.025453f
C442 VTAIL.n51 B 0.013677f
C443 VTAIL.n52 B 0.014482f
C444 VTAIL.n53 B 0.032328f
C445 VTAIL.n54 B 0.068163f
C446 VTAIL.n55 B 0.014482f
C447 VTAIL.n56 B 0.013677f
C448 VTAIL.n57 B 0.059529f
C449 VTAIL.n58 B 0.037974f
C450 VTAIL.n59 B 0.386253f
C451 VTAIL.t7 B 0.215218f
C452 VTAIL.t19 B 0.215218f
C453 VTAIL.n60 B 1.83039f
C454 VTAIL.n61 B 0.681735f
C455 VTAIL.t6 B 0.215218f
C456 VTAIL.t3 B 0.215218f
C457 VTAIL.n62 B 1.83039f
C458 VTAIL.n63 B 2.00107f
C459 VTAIL.t12 B 0.215218f
C460 VTAIL.t11 B 0.215218f
C461 VTAIL.n64 B 1.8304f
C462 VTAIL.n65 B 2.00106f
C463 VTAIL.t17 B 0.215218f
C464 VTAIL.t18 B 0.215218f
C465 VTAIL.n66 B 1.8304f
C466 VTAIL.n67 B 0.681724f
C467 VTAIL.n68 B 0.034746f
C468 VTAIL.n69 B 0.025453f
C469 VTAIL.n70 B 0.013677f
C470 VTAIL.n71 B 0.032328f
C471 VTAIL.n72 B 0.014482f
C472 VTAIL.n73 B 0.025453f
C473 VTAIL.n74 B 0.013677f
C474 VTAIL.n75 B 0.032328f
C475 VTAIL.n76 B 0.014482f
C476 VTAIL.n77 B 0.025453f
C477 VTAIL.n78 B 0.013677f
C478 VTAIL.n79 B 0.032328f
C479 VTAIL.n80 B 0.032328f
C480 VTAIL.n81 B 0.014482f
C481 VTAIL.n82 B 0.025453f
C482 VTAIL.n83 B 0.013677f
C483 VTAIL.n84 B 0.032328f
C484 VTAIL.n85 B 0.014482f
C485 VTAIL.n86 B 0.170812f
C486 VTAIL.t16 B 0.054423f
C487 VTAIL.n87 B 0.024246f
C488 VTAIL.n88 B 0.022854f
C489 VTAIL.n89 B 0.013677f
C490 VTAIL.n90 B 1.13689f
C491 VTAIL.n91 B 0.025453f
C492 VTAIL.n92 B 0.013677f
C493 VTAIL.n93 B 0.014482f
C494 VTAIL.n94 B 0.032328f
C495 VTAIL.n95 B 0.032328f
C496 VTAIL.n96 B 0.014482f
C497 VTAIL.n97 B 0.013677f
C498 VTAIL.n98 B 0.025453f
C499 VTAIL.n99 B 0.025453f
C500 VTAIL.n100 B 0.013677f
C501 VTAIL.n101 B 0.014482f
C502 VTAIL.n102 B 0.032328f
C503 VTAIL.n103 B 0.032328f
C504 VTAIL.n104 B 0.014482f
C505 VTAIL.n105 B 0.013677f
C506 VTAIL.n106 B 0.025453f
C507 VTAIL.n107 B 0.025453f
C508 VTAIL.n108 B 0.013677f
C509 VTAIL.n109 B 0.01408f
C510 VTAIL.n110 B 0.01408f
C511 VTAIL.n111 B 0.032328f
C512 VTAIL.n112 B 0.032328f
C513 VTAIL.n113 B 0.014482f
C514 VTAIL.n114 B 0.013677f
C515 VTAIL.n115 B 0.025453f
C516 VTAIL.n116 B 0.025453f
C517 VTAIL.n117 B 0.013677f
C518 VTAIL.n118 B 0.014482f
C519 VTAIL.n119 B 0.032328f
C520 VTAIL.n120 B 0.068163f
C521 VTAIL.n121 B 0.014482f
C522 VTAIL.n122 B 0.013677f
C523 VTAIL.n123 B 0.059529f
C524 VTAIL.n124 B 0.037974f
C525 VTAIL.n125 B 0.386253f
C526 VTAIL.t4 B 0.215218f
C527 VTAIL.t1 B 0.215218f
C528 VTAIL.n126 B 1.8304f
C529 VTAIL.n127 B 0.611728f
C530 VTAIL.t2 B 0.215218f
C531 VTAIL.t5 B 0.215218f
C532 VTAIL.n128 B 1.8304f
C533 VTAIL.n129 B 0.681724f
C534 VTAIL.n130 B 0.034746f
C535 VTAIL.n131 B 0.025453f
C536 VTAIL.n132 B 0.013677f
C537 VTAIL.n133 B 0.032328f
C538 VTAIL.n134 B 0.014482f
C539 VTAIL.n135 B 0.025453f
C540 VTAIL.n136 B 0.013677f
C541 VTAIL.n137 B 0.032328f
C542 VTAIL.n138 B 0.014482f
C543 VTAIL.n139 B 0.025453f
C544 VTAIL.n140 B 0.013677f
C545 VTAIL.n141 B 0.032328f
C546 VTAIL.n142 B 0.032328f
C547 VTAIL.n143 B 0.014482f
C548 VTAIL.n144 B 0.025453f
C549 VTAIL.n145 B 0.013677f
C550 VTAIL.n146 B 0.032328f
C551 VTAIL.n147 B 0.014482f
C552 VTAIL.n148 B 0.170812f
C553 VTAIL.t0 B 0.054423f
C554 VTAIL.n149 B 0.024246f
C555 VTAIL.n150 B 0.022854f
C556 VTAIL.n151 B 0.013677f
C557 VTAIL.n152 B 1.13689f
C558 VTAIL.n153 B 0.025453f
C559 VTAIL.n154 B 0.013677f
C560 VTAIL.n155 B 0.014482f
C561 VTAIL.n156 B 0.032328f
C562 VTAIL.n157 B 0.032328f
C563 VTAIL.n158 B 0.014482f
C564 VTAIL.n159 B 0.013677f
C565 VTAIL.n160 B 0.025453f
C566 VTAIL.n161 B 0.025453f
C567 VTAIL.n162 B 0.013677f
C568 VTAIL.n163 B 0.014482f
C569 VTAIL.n164 B 0.032328f
C570 VTAIL.n165 B 0.032328f
C571 VTAIL.n166 B 0.014482f
C572 VTAIL.n167 B 0.013677f
C573 VTAIL.n168 B 0.025453f
C574 VTAIL.n169 B 0.025453f
C575 VTAIL.n170 B 0.013677f
C576 VTAIL.n171 B 0.01408f
C577 VTAIL.n172 B 0.01408f
C578 VTAIL.n173 B 0.032328f
C579 VTAIL.n174 B 0.032328f
C580 VTAIL.n175 B 0.014482f
C581 VTAIL.n176 B 0.013677f
C582 VTAIL.n177 B 0.025453f
C583 VTAIL.n178 B 0.025453f
C584 VTAIL.n179 B 0.013677f
C585 VTAIL.n180 B 0.014482f
C586 VTAIL.n181 B 0.032328f
C587 VTAIL.n182 B 0.068163f
C588 VTAIL.n183 B 0.014482f
C589 VTAIL.n184 B 0.013677f
C590 VTAIL.n185 B 0.059529f
C591 VTAIL.n186 B 0.037974f
C592 VTAIL.n187 B 1.55852f
C593 VTAIL.n188 B 0.034746f
C594 VTAIL.n189 B 0.025453f
C595 VTAIL.n190 B 0.013677f
C596 VTAIL.n191 B 0.032328f
C597 VTAIL.n192 B 0.014482f
C598 VTAIL.n193 B 0.025453f
C599 VTAIL.n194 B 0.013677f
C600 VTAIL.n195 B 0.032328f
C601 VTAIL.n196 B 0.014482f
C602 VTAIL.n197 B 0.025453f
C603 VTAIL.n198 B 0.013677f
C604 VTAIL.n199 B 0.032328f
C605 VTAIL.n200 B 0.014482f
C606 VTAIL.n201 B 0.025453f
C607 VTAIL.n202 B 0.013677f
C608 VTAIL.n203 B 0.032328f
C609 VTAIL.n204 B 0.014482f
C610 VTAIL.n205 B 0.170812f
C611 VTAIL.t14 B 0.054423f
C612 VTAIL.n206 B 0.024246f
C613 VTAIL.n207 B 0.022854f
C614 VTAIL.n208 B 0.013677f
C615 VTAIL.n209 B 1.13689f
C616 VTAIL.n210 B 0.025453f
C617 VTAIL.n211 B 0.013677f
C618 VTAIL.n212 B 0.014482f
C619 VTAIL.n213 B 0.032328f
C620 VTAIL.n214 B 0.032328f
C621 VTAIL.n215 B 0.014482f
C622 VTAIL.n216 B 0.013677f
C623 VTAIL.n217 B 0.025453f
C624 VTAIL.n218 B 0.025453f
C625 VTAIL.n219 B 0.013677f
C626 VTAIL.n220 B 0.014482f
C627 VTAIL.n221 B 0.032328f
C628 VTAIL.n222 B 0.032328f
C629 VTAIL.n223 B 0.032328f
C630 VTAIL.n224 B 0.014482f
C631 VTAIL.n225 B 0.013677f
C632 VTAIL.n226 B 0.025453f
C633 VTAIL.n227 B 0.025453f
C634 VTAIL.n228 B 0.013677f
C635 VTAIL.n229 B 0.01408f
C636 VTAIL.n230 B 0.01408f
C637 VTAIL.n231 B 0.032328f
C638 VTAIL.n232 B 0.032328f
C639 VTAIL.n233 B 0.014482f
C640 VTAIL.n234 B 0.013677f
C641 VTAIL.n235 B 0.025453f
C642 VTAIL.n236 B 0.025453f
C643 VTAIL.n237 B 0.013677f
C644 VTAIL.n238 B 0.014482f
C645 VTAIL.n239 B 0.032328f
C646 VTAIL.n240 B 0.068163f
C647 VTAIL.n241 B 0.014482f
C648 VTAIL.n242 B 0.013677f
C649 VTAIL.n243 B 0.059529f
C650 VTAIL.n244 B 0.037974f
C651 VTAIL.n245 B 1.55852f
C652 VTAIL.t15 B 0.215218f
C653 VTAIL.t9 B 0.215218f
C654 VTAIL.n246 B 1.83039f
C655 VTAIL.n247 B 0.514168f
C656 VN.n0 B 0.027808f
C657 VN.t3 B 1.67911f
C658 VN.n1 B 0.03832f
C659 VN.n2 B 0.021093f
C660 VN.t4 B 1.67911f
C661 VN.n3 B 0.59701f
C662 VN.n4 B 0.021093f
C663 VN.n5 B 0.017368f
C664 VN.n6 B 0.021093f
C665 VN.t9 B 1.67911f
C666 VN.n7 B 0.039116f
C667 VN.n8 B 0.021093f
C668 VN.n9 B 0.039116f
C669 VN.t7 B 1.86727f
C670 VN.n10 B 0.636301f
C671 VN.t8 B 1.67911f
C672 VN.n11 B 0.653365f
C673 VN.n12 B 0.022509f
C674 VN.n13 B 0.206888f
C675 VN.n14 B 0.021093f
C676 VN.n15 B 0.021093f
C677 VN.n16 B 0.040818f
C678 VN.n17 B 0.017368f
C679 VN.n18 B 0.042255f
C680 VN.n19 B 0.021093f
C681 VN.n20 B 0.021093f
C682 VN.n21 B 0.021093f
C683 VN.n22 B 0.616816f
C684 VN.n23 B 0.039116f
C685 VN.n24 B 0.042255f
C686 VN.n25 B 0.021093f
C687 VN.n26 B 0.021093f
C688 VN.n27 B 0.021093f
C689 VN.n28 B 0.040818f
C690 VN.n29 B 0.039116f
C691 VN.n30 B 0.022509f
C692 VN.n31 B 0.021093f
C693 VN.n32 B 0.021093f
C694 VN.n33 B 0.036412f
C695 VN.n34 B 0.041922f
C696 VN.n35 B 0.0202f
C697 VN.n36 B 0.021093f
C698 VN.n37 B 0.021093f
C699 VN.n38 B 0.021093f
C700 VN.n39 B 0.039116f
C701 VN.n40 B 0.025212f
C702 VN.n41 B 0.667605f
C703 VN.n42 B 0.036942f
C704 VN.n43 B 0.027808f
C705 VN.t1 B 1.67911f
C706 VN.n44 B 0.03832f
C707 VN.n45 B 0.021093f
C708 VN.t6 B 1.67911f
C709 VN.n46 B 0.59701f
C710 VN.n47 B 0.021093f
C711 VN.n48 B 0.017368f
C712 VN.n49 B 0.021093f
C713 VN.t0 B 1.67911f
C714 VN.n50 B 0.039116f
C715 VN.n51 B 0.021093f
C716 VN.n52 B 0.039116f
C717 VN.t5 B 1.86727f
C718 VN.n53 B 0.636301f
C719 VN.t2 B 1.67911f
C720 VN.n54 B 0.653365f
C721 VN.n55 B 0.022509f
C722 VN.n56 B 0.206888f
C723 VN.n57 B 0.021093f
C724 VN.n58 B 0.021093f
C725 VN.n59 B 0.040818f
C726 VN.n60 B 0.017368f
C727 VN.n61 B 0.042255f
C728 VN.n62 B 0.021093f
C729 VN.n63 B 0.021093f
C730 VN.n64 B 0.021093f
C731 VN.n65 B 0.616816f
C732 VN.n66 B 0.039116f
C733 VN.n67 B 0.042255f
C734 VN.n68 B 0.021093f
C735 VN.n69 B 0.021093f
C736 VN.n70 B 0.021093f
C737 VN.n71 B 0.040818f
C738 VN.n72 B 0.039116f
C739 VN.n73 B 0.022509f
C740 VN.n74 B 0.021093f
C741 VN.n75 B 0.021093f
C742 VN.n76 B 0.036412f
C743 VN.n77 B 0.041922f
C744 VN.n78 B 0.0202f
C745 VN.n79 B 0.021093f
C746 VN.n80 B 0.021093f
C747 VN.n81 B 0.021093f
C748 VN.n82 B 0.039116f
C749 VN.n83 B 0.025212f
C750 VN.n84 B 0.667605f
C751 VN.n85 B 1.28759f
.ends

