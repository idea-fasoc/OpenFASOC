* NGSPICE file created from diff_pair_sample_0920.ext - technology: sky130A

.subckt diff_pair_sample_0920 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X1 VTAIL.t14 VP.t1 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=1.82
X2 VDD2.t7 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X3 VDD1.t6 VP.t2 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=1.82
X4 VDD1.t5 VP.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X5 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=1.82
X6 VTAIL.t1 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X7 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=1.82
X8 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=1.82
X9 VDD1.t7 VP.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X10 VDD1.t0 VP.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=1.82
X11 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=1.82
X12 VTAIL.t9 VP.t6 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=1.82
X13 VTAIL.t8 VP.t7 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X14 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=1.0179 ps=6 w=2.61 l=1.82
X15 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=1.82
X16 VTAIL.t6 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
X17 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0.43065 ps=2.94 w=2.61 l=1.82
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0179 pd=6 as=0 ps=0 w=2.61 l=1.82
X19 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.43065 pd=2.94 as=0.43065 ps=2.94 w=2.61 l=1.82
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n20 VP.n19 161.3
R5 VP.n21 VP.n7 161.3
R6 VP.n23 VP.n22 161.3
R7 VP.n24 VP.n6 161.3
R8 VP.n48 VP.n0 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n1 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n41 VP.n2 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n3 161.3
R15 VP.n37 VP.n36 161.3
R16 VP.n34 VP.n4 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n31 VP.n5 161.3
R19 VP.n30 VP.n29 161.3
R20 VP.n28 VP.n27 87.5128
R21 VP.n50 VP.n49 87.5128
R22 VP.n26 VP.n25 87.5128
R23 VP.n10 VP.t1 65.9947
R24 VP.n40 VP.n3 56.5193
R25 VP.n16 VP.n9 56.5193
R26 VP.n11 VP.n10 53.8955
R27 VP.n33 VP.n5 50.2061
R28 VP.n47 VP.n1 50.2061
R29 VP.n23 VP.n7 50.2061
R30 VP.n27 VP.n26 40.1663
R31 VP.n28 VP.t6 34.5615
R32 VP.n35 VP.t4 34.5615
R33 VP.n42 VP.t7 34.5615
R34 VP.n49 VP.t5 34.5615
R35 VP.n25 VP.t2 34.5615
R36 VP.n18 VP.t0 34.5615
R37 VP.n11 VP.t3 34.5615
R38 VP.n29 VP.n5 30.7807
R39 VP.n48 VP.n47 30.7807
R40 VP.n24 VP.n23 30.7807
R41 VP.n34 VP.n33 24.4675
R42 VP.n36 VP.n3 24.4675
R43 VP.n41 VP.n40 24.4675
R44 VP.n43 VP.n1 24.4675
R45 VP.n17 VP.n16 24.4675
R46 VP.n19 VP.n7 24.4675
R47 VP.n12 VP.n9 24.4675
R48 VP.n29 VP.n28 23.2442
R49 VP.n49 VP.n48 23.2442
R50 VP.n25 VP.n24 23.2442
R51 VP.n36 VP.n35 15.9041
R52 VP.n42 VP.n41 15.9041
R53 VP.n18 VP.n17 15.9041
R54 VP.n12 VP.n11 15.9041
R55 VP.n13 VP.n10 12.7761
R56 VP.n35 VP.n34 8.56395
R57 VP.n43 VP.n42 8.56395
R58 VP.n19 VP.n18 8.56395
R59 VP.n26 VP.n6 0.278367
R60 VP.n30 VP.n27 0.278367
R61 VP.n50 VP.n0 0.278367
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153454
R81 VDD1 VDD1.n0 90.0169
R82 VDD1.n3 VDD1.n2 89.9033
R83 VDD1.n3 VDD1.n1 89.9033
R84 VDD1.n5 VDD1.n4 89.0319
R85 VDD1.n5 VDD1.n3 34.8888
R86 VDD1.n4 VDD1.t4 7.58671
R87 VDD1.n4 VDD1.t6 7.58671
R88 VDD1.n0 VDD1.t1 7.58671
R89 VDD1.n0 VDD1.t5 7.58671
R90 VDD1.n2 VDD1.t3 7.58671
R91 VDD1.n2 VDD1.t0 7.58671
R92 VDD1.n1 VDD1.t2 7.58671
R93 VDD1.n1 VDD1.t7 7.58671
R94 VDD1 VDD1.n5 0.869035
R95 VTAIL.n98 VTAIL.n92 289.615
R96 VTAIL.n8 VTAIL.n2 289.615
R97 VTAIL.n20 VTAIL.n14 289.615
R98 VTAIL.n34 VTAIL.n28 289.615
R99 VTAIL.n86 VTAIL.n80 289.615
R100 VTAIL.n72 VTAIL.n66 289.615
R101 VTAIL.n60 VTAIL.n54 289.615
R102 VTAIL.n46 VTAIL.n40 289.615
R103 VTAIL.n97 VTAIL.n96 185
R104 VTAIL.n99 VTAIL.n98 185
R105 VTAIL.n7 VTAIL.n6 185
R106 VTAIL.n9 VTAIL.n8 185
R107 VTAIL.n19 VTAIL.n18 185
R108 VTAIL.n21 VTAIL.n20 185
R109 VTAIL.n33 VTAIL.n32 185
R110 VTAIL.n35 VTAIL.n34 185
R111 VTAIL.n87 VTAIL.n86 185
R112 VTAIL.n85 VTAIL.n84 185
R113 VTAIL.n73 VTAIL.n72 185
R114 VTAIL.n71 VTAIL.n70 185
R115 VTAIL.n61 VTAIL.n60 185
R116 VTAIL.n59 VTAIL.n58 185
R117 VTAIL.n47 VTAIL.n46 185
R118 VTAIL.n45 VTAIL.n44 185
R119 VTAIL.n95 VTAIL.t3 151.613
R120 VTAIL.n5 VTAIL.t2 151.613
R121 VTAIL.n17 VTAIL.t10 151.613
R122 VTAIL.n31 VTAIL.t9 151.613
R123 VTAIL.n83 VTAIL.t13 151.613
R124 VTAIL.n69 VTAIL.t14 151.613
R125 VTAIL.n57 VTAIL.t5 151.613
R126 VTAIL.n43 VTAIL.t0 151.613
R127 VTAIL.n98 VTAIL.n97 104.615
R128 VTAIL.n8 VTAIL.n7 104.615
R129 VTAIL.n20 VTAIL.n19 104.615
R130 VTAIL.n34 VTAIL.n33 104.615
R131 VTAIL.n86 VTAIL.n85 104.615
R132 VTAIL.n72 VTAIL.n71 104.615
R133 VTAIL.n60 VTAIL.n59 104.615
R134 VTAIL.n46 VTAIL.n45 104.615
R135 VTAIL.n79 VTAIL.n78 72.3532
R136 VTAIL.n53 VTAIL.n52 72.3532
R137 VTAIL.n1 VTAIL.n0 72.3531
R138 VTAIL.n27 VTAIL.n26 72.3531
R139 VTAIL.n97 VTAIL.t3 52.3082
R140 VTAIL.n7 VTAIL.t2 52.3082
R141 VTAIL.n19 VTAIL.t10 52.3082
R142 VTAIL.n33 VTAIL.t9 52.3082
R143 VTAIL.n85 VTAIL.t13 52.3082
R144 VTAIL.n71 VTAIL.t14 52.3082
R145 VTAIL.n59 VTAIL.t5 52.3082
R146 VTAIL.n45 VTAIL.t0 52.3082
R147 VTAIL.n103 VTAIL.n102 36.2581
R148 VTAIL.n13 VTAIL.n12 36.2581
R149 VTAIL.n25 VTAIL.n24 36.2581
R150 VTAIL.n39 VTAIL.n38 36.2581
R151 VTAIL.n91 VTAIL.n90 36.2581
R152 VTAIL.n77 VTAIL.n76 36.2581
R153 VTAIL.n65 VTAIL.n64 36.2581
R154 VTAIL.n51 VTAIL.n50 36.2581
R155 VTAIL.n103 VTAIL.n91 16.4703
R156 VTAIL.n51 VTAIL.n39 16.4703
R157 VTAIL.n96 VTAIL.n95 15.3979
R158 VTAIL.n6 VTAIL.n5 15.3979
R159 VTAIL.n18 VTAIL.n17 15.3979
R160 VTAIL.n32 VTAIL.n31 15.3979
R161 VTAIL.n84 VTAIL.n83 15.3979
R162 VTAIL.n70 VTAIL.n69 15.3979
R163 VTAIL.n58 VTAIL.n57 15.3979
R164 VTAIL.n44 VTAIL.n43 15.3979
R165 VTAIL.n99 VTAIL.n94 12.8005
R166 VTAIL.n9 VTAIL.n4 12.8005
R167 VTAIL.n21 VTAIL.n16 12.8005
R168 VTAIL.n35 VTAIL.n30 12.8005
R169 VTAIL.n87 VTAIL.n82 12.8005
R170 VTAIL.n73 VTAIL.n68 12.8005
R171 VTAIL.n61 VTAIL.n56 12.8005
R172 VTAIL.n47 VTAIL.n42 12.8005
R173 VTAIL.n100 VTAIL.n92 12.0247
R174 VTAIL.n10 VTAIL.n2 12.0247
R175 VTAIL.n22 VTAIL.n14 12.0247
R176 VTAIL.n36 VTAIL.n28 12.0247
R177 VTAIL.n88 VTAIL.n80 12.0247
R178 VTAIL.n74 VTAIL.n66 12.0247
R179 VTAIL.n62 VTAIL.n54 12.0247
R180 VTAIL.n48 VTAIL.n40 12.0247
R181 VTAIL.n102 VTAIL.n101 9.45567
R182 VTAIL.n12 VTAIL.n11 9.45567
R183 VTAIL.n24 VTAIL.n23 9.45567
R184 VTAIL.n38 VTAIL.n37 9.45567
R185 VTAIL.n90 VTAIL.n89 9.45567
R186 VTAIL.n76 VTAIL.n75 9.45567
R187 VTAIL.n64 VTAIL.n63 9.45567
R188 VTAIL.n50 VTAIL.n49 9.45567
R189 VTAIL.n101 VTAIL.n100 9.3005
R190 VTAIL.n94 VTAIL.n93 9.3005
R191 VTAIL.n11 VTAIL.n10 9.3005
R192 VTAIL.n4 VTAIL.n3 9.3005
R193 VTAIL.n23 VTAIL.n22 9.3005
R194 VTAIL.n16 VTAIL.n15 9.3005
R195 VTAIL.n37 VTAIL.n36 9.3005
R196 VTAIL.n30 VTAIL.n29 9.3005
R197 VTAIL.n89 VTAIL.n88 9.3005
R198 VTAIL.n82 VTAIL.n81 9.3005
R199 VTAIL.n75 VTAIL.n74 9.3005
R200 VTAIL.n68 VTAIL.n67 9.3005
R201 VTAIL.n63 VTAIL.n62 9.3005
R202 VTAIL.n56 VTAIL.n55 9.3005
R203 VTAIL.n49 VTAIL.n48 9.3005
R204 VTAIL.n42 VTAIL.n41 9.3005
R205 VTAIL.n0 VTAIL.t4 7.58671
R206 VTAIL.n0 VTAIL.t1 7.58671
R207 VTAIL.n26 VTAIL.t11 7.58671
R208 VTAIL.n26 VTAIL.t8 7.58671
R209 VTAIL.n78 VTAIL.t12 7.58671
R210 VTAIL.n78 VTAIL.t15 7.58671
R211 VTAIL.n52 VTAIL.t7 7.58671
R212 VTAIL.n52 VTAIL.t6 7.58671
R213 VTAIL.n95 VTAIL.n93 4.69785
R214 VTAIL.n5 VTAIL.n3 4.69785
R215 VTAIL.n17 VTAIL.n15 4.69785
R216 VTAIL.n31 VTAIL.n29 4.69785
R217 VTAIL.n83 VTAIL.n81 4.69785
R218 VTAIL.n69 VTAIL.n67 4.69785
R219 VTAIL.n57 VTAIL.n55 4.69785
R220 VTAIL.n43 VTAIL.n41 4.69785
R221 VTAIL.n102 VTAIL.n92 1.93989
R222 VTAIL.n12 VTAIL.n2 1.93989
R223 VTAIL.n24 VTAIL.n14 1.93989
R224 VTAIL.n38 VTAIL.n28 1.93989
R225 VTAIL.n90 VTAIL.n80 1.93989
R226 VTAIL.n76 VTAIL.n66 1.93989
R227 VTAIL.n64 VTAIL.n54 1.93989
R228 VTAIL.n50 VTAIL.n40 1.93989
R229 VTAIL.n53 VTAIL.n51 1.85395
R230 VTAIL.n65 VTAIL.n53 1.85395
R231 VTAIL.n79 VTAIL.n77 1.85395
R232 VTAIL.n91 VTAIL.n79 1.85395
R233 VTAIL.n39 VTAIL.n27 1.85395
R234 VTAIL.n27 VTAIL.n25 1.85395
R235 VTAIL.n13 VTAIL.n1 1.85395
R236 VTAIL VTAIL.n103 1.79576
R237 VTAIL.n100 VTAIL.n99 1.16414
R238 VTAIL.n10 VTAIL.n9 1.16414
R239 VTAIL.n22 VTAIL.n21 1.16414
R240 VTAIL.n36 VTAIL.n35 1.16414
R241 VTAIL.n88 VTAIL.n87 1.16414
R242 VTAIL.n74 VTAIL.n73 1.16414
R243 VTAIL.n62 VTAIL.n61 1.16414
R244 VTAIL.n48 VTAIL.n47 1.16414
R245 VTAIL.n77 VTAIL.n65 0.470328
R246 VTAIL.n25 VTAIL.n13 0.470328
R247 VTAIL.n96 VTAIL.n94 0.388379
R248 VTAIL.n6 VTAIL.n4 0.388379
R249 VTAIL.n18 VTAIL.n16 0.388379
R250 VTAIL.n32 VTAIL.n30 0.388379
R251 VTAIL.n84 VTAIL.n82 0.388379
R252 VTAIL.n70 VTAIL.n68 0.388379
R253 VTAIL.n58 VTAIL.n56 0.388379
R254 VTAIL.n44 VTAIL.n42 0.388379
R255 VTAIL.n101 VTAIL.n93 0.155672
R256 VTAIL.n11 VTAIL.n3 0.155672
R257 VTAIL.n23 VTAIL.n15 0.155672
R258 VTAIL.n37 VTAIL.n29 0.155672
R259 VTAIL.n89 VTAIL.n81 0.155672
R260 VTAIL.n75 VTAIL.n67 0.155672
R261 VTAIL.n63 VTAIL.n55 0.155672
R262 VTAIL.n49 VTAIL.n41 0.155672
R263 VTAIL VTAIL.n1 0.0586897
R264 B.n515 B.n514 585
R265 B.n169 B.n93 585
R266 B.n168 B.n167 585
R267 B.n166 B.n165 585
R268 B.n164 B.n163 585
R269 B.n162 B.n161 585
R270 B.n160 B.n159 585
R271 B.n158 B.n157 585
R272 B.n156 B.n155 585
R273 B.n154 B.n153 585
R274 B.n152 B.n151 585
R275 B.n150 B.n149 585
R276 B.n148 B.n147 585
R277 B.n146 B.n145 585
R278 B.n144 B.n143 585
R279 B.n142 B.n141 585
R280 B.n140 B.n139 585
R281 B.n138 B.n137 585
R282 B.n136 B.n135 585
R283 B.n134 B.n133 585
R284 B.n132 B.n131 585
R285 B.n130 B.n129 585
R286 B.n128 B.n127 585
R287 B.n126 B.n125 585
R288 B.n124 B.n123 585
R289 B.n122 B.n121 585
R290 B.n120 B.n119 585
R291 B.n118 B.n117 585
R292 B.n116 B.n115 585
R293 B.n114 B.n113 585
R294 B.n112 B.n111 585
R295 B.n110 B.n109 585
R296 B.n108 B.n107 585
R297 B.n106 B.n105 585
R298 B.n104 B.n103 585
R299 B.n102 B.n101 585
R300 B.n75 B.n74 585
R301 B.n520 B.n519 585
R302 B.n513 B.n94 585
R303 B.n94 B.n72 585
R304 B.n512 B.n71 585
R305 B.n524 B.n71 585
R306 B.n511 B.n70 585
R307 B.n525 B.n70 585
R308 B.n510 B.n69 585
R309 B.n526 B.n69 585
R310 B.n509 B.n508 585
R311 B.n508 B.n65 585
R312 B.n507 B.n64 585
R313 B.n532 B.n64 585
R314 B.n506 B.n63 585
R315 B.n533 B.n63 585
R316 B.n505 B.n62 585
R317 B.n534 B.n62 585
R318 B.n504 B.n503 585
R319 B.n503 B.n58 585
R320 B.n502 B.n57 585
R321 B.n540 B.n57 585
R322 B.n501 B.n56 585
R323 B.n541 B.n56 585
R324 B.n500 B.n55 585
R325 B.n542 B.n55 585
R326 B.n499 B.n498 585
R327 B.n498 B.n51 585
R328 B.n497 B.n50 585
R329 B.n548 B.n50 585
R330 B.n496 B.n49 585
R331 B.n549 B.n49 585
R332 B.n495 B.n48 585
R333 B.n550 B.n48 585
R334 B.n494 B.n493 585
R335 B.n493 B.n44 585
R336 B.n492 B.n43 585
R337 B.n556 B.n43 585
R338 B.n491 B.n42 585
R339 B.n557 B.n42 585
R340 B.n490 B.n41 585
R341 B.n558 B.n41 585
R342 B.n489 B.n488 585
R343 B.n488 B.n37 585
R344 B.n487 B.n36 585
R345 B.n564 B.n36 585
R346 B.n486 B.n35 585
R347 B.n565 B.n35 585
R348 B.n485 B.n34 585
R349 B.n566 B.n34 585
R350 B.n484 B.n483 585
R351 B.n483 B.n30 585
R352 B.n482 B.n29 585
R353 B.n572 B.n29 585
R354 B.n481 B.n28 585
R355 B.n573 B.n28 585
R356 B.n480 B.n27 585
R357 B.n574 B.n27 585
R358 B.n479 B.n478 585
R359 B.n478 B.n26 585
R360 B.n477 B.n22 585
R361 B.n580 B.n22 585
R362 B.n476 B.n21 585
R363 B.n581 B.n21 585
R364 B.n475 B.n20 585
R365 B.n582 B.n20 585
R366 B.n474 B.n473 585
R367 B.n473 B.n16 585
R368 B.n472 B.n15 585
R369 B.n588 B.n15 585
R370 B.n471 B.n14 585
R371 B.n589 B.n14 585
R372 B.n470 B.n13 585
R373 B.n590 B.n13 585
R374 B.n469 B.n468 585
R375 B.n468 B.n12 585
R376 B.n467 B.n466 585
R377 B.n467 B.n8 585
R378 B.n465 B.n7 585
R379 B.n597 B.n7 585
R380 B.n464 B.n6 585
R381 B.n598 B.n6 585
R382 B.n463 B.n5 585
R383 B.n599 B.n5 585
R384 B.n462 B.n461 585
R385 B.n461 B.n4 585
R386 B.n460 B.n170 585
R387 B.n460 B.n459 585
R388 B.n450 B.n171 585
R389 B.n172 B.n171 585
R390 B.n452 B.n451 585
R391 B.n453 B.n452 585
R392 B.n449 B.n176 585
R393 B.n180 B.n176 585
R394 B.n448 B.n447 585
R395 B.n447 B.n446 585
R396 B.n178 B.n177 585
R397 B.n179 B.n178 585
R398 B.n439 B.n438 585
R399 B.n440 B.n439 585
R400 B.n437 B.n185 585
R401 B.n185 B.n184 585
R402 B.n436 B.n435 585
R403 B.n435 B.n434 585
R404 B.n187 B.n186 585
R405 B.n427 B.n187 585
R406 B.n426 B.n425 585
R407 B.n428 B.n426 585
R408 B.n424 B.n192 585
R409 B.n192 B.n191 585
R410 B.n423 B.n422 585
R411 B.n422 B.n421 585
R412 B.n194 B.n193 585
R413 B.n195 B.n194 585
R414 B.n414 B.n413 585
R415 B.n415 B.n414 585
R416 B.n412 B.n199 585
R417 B.n203 B.n199 585
R418 B.n411 B.n410 585
R419 B.n410 B.n409 585
R420 B.n201 B.n200 585
R421 B.n202 B.n201 585
R422 B.n402 B.n401 585
R423 B.n403 B.n402 585
R424 B.n400 B.n208 585
R425 B.n208 B.n207 585
R426 B.n399 B.n398 585
R427 B.n398 B.n397 585
R428 B.n210 B.n209 585
R429 B.n211 B.n210 585
R430 B.n390 B.n389 585
R431 B.n391 B.n390 585
R432 B.n388 B.n216 585
R433 B.n216 B.n215 585
R434 B.n387 B.n386 585
R435 B.n386 B.n385 585
R436 B.n218 B.n217 585
R437 B.n219 B.n218 585
R438 B.n378 B.n377 585
R439 B.n379 B.n378 585
R440 B.n376 B.n224 585
R441 B.n224 B.n223 585
R442 B.n375 B.n374 585
R443 B.n374 B.n373 585
R444 B.n226 B.n225 585
R445 B.n227 B.n226 585
R446 B.n366 B.n365 585
R447 B.n367 B.n366 585
R448 B.n364 B.n231 585
R449 B.n235 B.n231 585
R450 B.n363 B.n362 585
R451 B.n362 B.n361 585
R452 B.n233 B.n232 585
R453 B.n234 B.n233 585
R454 B.n354 B.n353 585
R455 B.n355 B.n354 585
R456 B.n352 B.n240 585
R457 B.n240 B.n239 585
R458 B.n351 B.n350 585
R459 B.n350 B.n349 585
R460 B.n242 B.n241 585
R461 B.n243 B.n242 585
R462 B.n345 B.n344 585
R463 B.n246 B.n245 585
R464 B.n341 B.n340 585
R465 B.n342 B.n341 585
R466 B.n339 B.n265 585
R467 B.n338 B.n337 585
R468 B.n336 B.n335 585
R469 B.n334 B.n333 585
R470 B.n332 B.n331 585
R471 B.n330 B.n329 585
R472 B.n328 B.n327 585
R473 B.n326 B.n325 585
R474 B.n324 B.n323 585
R475 B.n322 B.n321 585
R476 B.n320 B.n319 585
R477 B.n317 B.n316 585
R478 B.n315 B.n314 585
R479 B.n313 B.n312 585
R480 B.n311 B.n310 585
R481 B.n309 B.n308 585
R482 B.n307 B.n306 585
R483 B.n305 B.n304 585
R484 B.n303 B.n302 585
R485 B.n301 B.n300 585
R486 B.n299 B.n298 585
R487 B.n296 B.n295 585
R488 B.n294 B.n293 585
R489 B.n292 B.n291 585
R490 B.n290 B.n289 585
R491 B.n288 B.n287 585
R492 B.n286 B.n285 585
R493 B.n284 B.n283 585
R494 B.n282 B.n281 585
R495 B.n280 B.n279 585
R496 B.n278 B.n277 585
R497 B.n276 B.n275 585
R498 B.n274 B.n273 585
R499 B.n272 B.n271 585
R500 B.n270 B.n264 585
R501 B.n342 B.n264 585
R502 B.n346 B.n244 585
R503 B.n244 B.n243 585
R504 B.n348 B.n347 585
R505 B.n349 B.n348 585
R506 B.n238 B.n237 585
R507 B.n239 B.n238 585
R508 B.n357 B.n356 585
R509 B.n356 B.n355 585
R510 B.n358 B.n236 585
R511 B.n236 B.n234 585
R512 B.n360 B.n359 585
R513 B.n361 B.n360 585
R514 B.n230 B.n229 585
R515 B.n235 B.n230 585
R516 B.n369 B.n368 585
R517 B.n368 B.n367 585
R518 B.n370 B.n228 585
R519 B.n228 B.n227 585
R520 B.n372 B.n371 585
R521 B.n373 B.n372 585
R522 B.n222 B.n221 585
R523 B.n223 B.n222 585
R524 B.n381 B.n380 585
R525 B.n380 B.n379 585
R526 B.n382 B.n220 585
R527 B.n220 B.n219 585
R528 B.n384 B.n383 585
R529 B.n385 B.n384 585
R530 B.n214 B.n213 585
R531 B.n215 B.n214 585
R532 B.n393 B.n392 585
R533 B.n392 B.n391 585
R534 B.n394 B.n212 585
R535 B.n212 B.n211 585
R536 B.n396 B.n395 585
R537 B.n397 B.n396 585
R538 B.n206 B.n205 585
R539 B.n207 B.n206 585
R540 B.n405 B.n404 585
R541 B.n404 B.n403 585
R542 B.n406 B.n204 585
R543 B.n204 B.n202 585
R544 B.n408 B.n407 585
R545 B.n409 B.n408 585
R546 B.n198 B.n197 585
R547 B.n203 B.n198 585
R548 B.n417 B.n416 585
R549 B.n416 B.n415 585
R550 B.n418 B.n196 585
R551 B.n196 B.n195 585
R552 B.n420 B.n419 585
R553 B.n421 B.n420 585
R554 B.n190 B.n189 585
R555 B.n191 B.n190 585
R556 B.n430 B.n429 585
R557 B.n429 B.n428 585
R558 B.n431 B.n188 585
R559 B.n427 B.n188 585
R560 B.n433 B.n432 585
R561 B.n434 B.n433 585
R562 B.n183 B.n182 585
R563 B.n184 B.n183 585
R564 B.n442 B.n441 585
R565 B.n441 B.n440 585
R566 B.n443 B.n181 585
R567 B.n181 B.n179 585
R568 B.n445 B.n444 585
R569 B.n446 B.n445 585
R570 B.n175 B.n174 585
R571 B.n180 B.n175 585
R572 B.n455 B.n454 585
R573 B.n454 B.n453 585
R574 B.n456 B.n173 585
R575 B.n173 B.n172 585
R576 B.n458 B.n457 585
R577 B.n459 B.n458 585
R578 B.n3 B.n0 585
R579 B.n4 B.n3 585
R580 B.n596 B.n1 585
R581 B.n597 B.n596 585
R582 B.n595 B.n594 585
R583 B.n595 B.n8 585
R584 B.n593 B.n9 585
R585 B.n12 B.n9 585
R586 B.n592 B.n591 585
R587 B.n591 B.n590 585
R588 B.n11 B.n10 585
R589 B.n589 B.n11 585
R590 B.n587 B.n586 585
R591 B.n588 B.n587 585
R592 B.n585 B.n17 585
R593 B.n17 B.n16 585
R594 B.n584 B.n583 585
R595 B.n583 B.n582 585
R596 B.n19 B.n18 585
R597 B.n581 B.n19 585
R598 B.n579 B.n578 585
R599 B.n580 B.n579 585
R600 B.n577 B.n23 585
R601 B.n26 B.n23 585
R602 B.n576 B.n575 585
R603 B.n575 B.n574 585
R604 B.n25 B.n24 585
R605 B.n573 B.n25 585
R606 B.n571 B.n570 585
R607 B.n572 B.n571 585
R608 B.n569 B.n31 585
R609 B.n31 B.n30 585
R610 B.n568 B.n567 585
R611 B.n567 B.n566 585
R612 B.n33 B.n32 585
R613 B.n565 B.n33 585
R614 B.n563 B.n562 585
R615 B.n564 B.n563 585
R616 B.n561 B.n38 585
R617 B.n38 B.n37 585
R618 B.n560 B.n559 585
R619 B.n559 B.n558 585
R620 B.n40 B.n39 585
R621 B.n557 B.n40 585
R622 B.n555 B.n554 585
R623 B.n556 B.n555 585
R624 B.n553 B.n45 585
R625 B.n45 B.n44 585
R626 B.n552 B.n551 585
R627 B.n551 B.n550 585
R628 B.n47 B.n46 585
R629 B.n549 B.n47 585
R630 B.n547 B.n546 585
R631 B.n548 B.n547 585
R632 B.n545 B.n52 585
R633 B.n52 B.n51 585
R634 B.n544 B.n543 585
R635 B.n543 B.n542 585
R636 B.n54 B.n53 585
R637 B.n541 B.n54 585
R638 B.n539 B.n538 585
R639 B.n540 B.n539 585
R640 B.n537 B.n59 585
R641 B.n59 B.n58 585
R642 B.n536 B.n535 585
R643 B.n535 B.n534 585
R644 B.n61 B.n60 585
R645 B.n533 B.n61 585
R646 B.n531 B.n530 585
R647 B.n532 B.n531 585
R648 B.n529 B.n66 585
R649 B.n66 B.n65 585
R650 B.n528 B.n527 585
R651 B.n527 B.n526 585
R652 B.n68 B.n67 585
R653 B.n525 B.n68 585
R654 B.n523 B.n522 585
R655 B.n524 B.n523 585
R656 B.n521 B.n73 585
R657 B.n73 B.n72 585
R658 B.n600 B.n599 585
R659 B.n598 B.n2 585
R660 B.n519 B.n73 502.111
R661 B.n515 B.n94 502.111
R662 B.n264 B.n242 502.111
R663 B.n344 B.n244 502.111
R664 B.n517 B.n516 256.663
R665 B.n517 B.n92 256.663
R666 B.n517 B.n91 256.663
R667 B.n517 B.n90 256.663
R668 B.n517 B.n89 256.663
R669 B.n517 B.n88 256.663
R670 B.n517 B.n87 256.663
R671 B.n517 B.n86 256.663
R672 B.n517 B.n85 256.663
R673 B.n517 B.n84 256.663
R674 B.n517 B.n83 256.663
R675 B.n517 B.n82 256.663
R676 B.n517 B.n81 256.663
R677 B.n517 B.n80 256.663
R678 B.n517 B.n79 256.663
R679 B.n517 B.n78 256.663
R680 B.n517 B.n77 256.663
R681 B.n517 B.n76 256.663
R682 B.n518 B.n517 256.663
R683 B.n343 B.n342 256.663
R684 B.n342 B.n247 256.663
R685 B.n342 B.n248 256.663
R686 B.n342 B.n249 256.663
R687 B.n342 B.n250 256.663
R688 B.n342 B.n251 256.663
R689 B.n342 B.n252 256.663
R690 B.n342 B.n253 256.663
R691 B.n342 B.n254 256.663
R692 B.n342 B.n255 256.663
R693 B.n342 B.n256 256.663
R694 B.n342 B.n257 256.663
R695 B.n342 B.n258 256.663
R696 B.n342 B.n259 256.663
R697 B.n342 B.n260 256.663
R698 B.n342 B.n261 256.663
R699 B.n342 B.n262 256.663
R700 B.n342 B.n263 256.663
R701 B.n602 B.n601 256.663
R702 B.n98 B.t12 241.023
R703 B.n95 B.t8 241.023
R704 B.n268 B.t15 241.023
R705 B.n266 B.t19 241.023
R706 B.n342 B.n243 193.912
R707 B.n517 B.n72 193.912
R708 B.n95 B.t10 166.53
R709 B.n268 B.t18 166.53
R710 B.n98 B.t13 166.53
R711 B.n266 B.t21 166.53
R712 B.n101 B.n75 163.367
R713 B.n105 B.n104 163.367
R714 B.n109 B.n108 163.367
R715 B.n113 B.n112 163.367
R716 B.n117 B.n116 163.367
R717 B.n121 B.n120 163.367
R718 B.n125 B.n124 163.367
R719 B.n129 B.n128 163.367
R720 B.n133 B.n132 163.367
R721 B.n137 B.n136 163.367
R722 B.n141 B.n140 163.367
R723 B.n145 B.n144 163.367
R724 B.n149 B.n148 163.367
R725 B.n153 B.n152 163.367
R726 B.n157 B.n156 163.367
R727 B.n161 B.n160 163.367
R728 B.n165 B.n164 163.367
R729 B.n167 B.n93 163.367
R730 B.n350 B.n242 163.367
R731 B.n350 B.n240 163.367
R732 B.n354 B.n240 163.367
R733 B.n354 B.n233 163.367
R734 B.n362 B.n233 163.367
R735 B.n362 B.n231 163.367
R736 B.n366 B.n231 163.367
R737 B.n366 B.n226 163.367
R738 B.n374 B.n226 163.367
R739 B.n374 B.n224 163.367
R740 B.n378 B.n224 163.367
R741 B.n378 B.n218 163.367
R742 B.n386 B.n218 163.367
R743 B.n386 B.n216 163.367
R744 B.n390 B.n216 163.367
R745 B.n390 B.n210 163.367
R746 B.n398 B.n210 163.367
R747 B.n398 B.n208 163.367
R748 B.n402 B.n208 163.367
R749 B.n402 B.n201 163.367
R750 B.n410 B.n201 163.367
R751 B.n410 B.n199 163.367
R752 B.n414 B.n199 163.367
R753 B.n414 B.n194 163.367
R754 B.n422 B.n194 163.367
R755 B.n422 B.n192 163.367
R756 B.n426 B.n192 163.367
R757 B.n426 B.n187 163.367
R758 B.n435 B.n187 163.367
R759 B.n435 B.n185 163.367
R760 B.n439 B.n185 163.367
R761 B.n439 B.n178 163.367
R762 B.n447 B.n178 163.367
R763 B.n447 B.n176 163.367
R764 B.n452 B.n176 163.367
R765 B.n452 B.n171 163.367
R766 B.n460 B.n171 163.367
R767 B.n461 B.n460 163.367
R768 B.n461 B.n5 163.367
R769 B.n6 B.n5 163.367
R770 B.n7 B.n6 163.367
R771 B.n467 B.n7 163.367
R772 B.n468 B.n467 163.367
R773 B.n468 B.n13 163.367
R774 B.n14 B.n13 163.367
R775 B.n15 B.n14 163.367
R776 B.n473 B.n15 163.367
R777 B.n473 B.n20 163.367
R778 B.n21 B.n20 163.367
R779 B.n22 B.n21 163.367
R780 B.n478 B.n22 163.367
R781 B.n478 B.n27 163.367
R782 B.n28 B.n27 163.367
R783 B.n29 B.n28 163.367
R784 B.n483 B.n29 163.367
R785 B.n483 B.n34 163.367
R786 B.n35 B.n34 163.367
R787 B.n36 B.n35 163.367
R788 B.n488 B.n36 163.367
R789 B.n488 B.n41 163.367
R790 B.n42 B.n41 163.367
R791 B.n43 B.n42 163.367
R792 B.n493 B.n43 163.367
R793 B.n493 B.n48 163.367
R794 B.n49 B.n48 163.367
R795 B.n50 B.n49 163.367
R796 B.n498 B.n50 163.367
R797 B.n498 B.n55 163.367
R798 B.n56 B.n55 163.367
R799 B.n57 B.n56 163.367
R800 B.n503 B.n57 163.367
R801 B.n503 B.n62 163.367
R802 B.n63 B.n62 163.367
R803 B.n64 B.n63 163.367
R804 B.n508 B.n64 163.367
R805 B.n508 B.n69 163.367
R806 B.n70 B.n69 163.367
R807 B.n71 B.n70 163.367
R808 B.n94 B.n71 163.367
R809 B.n341 B.n246 163.367
R810 B.n341 B.n265 163.367
R811 B.n337 B.n336 163.367
R812 B.n333 B.n332 163.367
R813 B.n329 B.n328 163.367
R814 B.n325 B.n324 163.367
R815 B.n321 B.n320 163.367
R816 B.n316 B.n315 163.367
R817 B.n312 B.n311 163.367
R818 B.n308 B.n307 163.367
R819 B.n304 B.n303 163.367
R820 B.n300 B.n299 163.367
R821 B.n295 B.n294 163.367
R822 B.n291 B.n290 163.367
R823 B.n287 B.n286 163.367
R824 B.n283 B.n282 163.367
R825 B.n279 B.n278 163.367
R826 B.n275 B.n274 163.367
R827 B.n271 B.n264 163.367
R828 B.n348 B.n244 163.367
R829 B.n348 B.n238 163.367
R830 B.n356 B.n238 163.367
R831 B.n356 B.n236 163.367
R832 B.n360 B.n236 163.367
R833 B.n360 B.n230 163.367
R834 B.n368 B.n230 163.367
R835 B.n368 B.n228 163.367
R836 B.n372 B.n228 163.367
R837 B.n372 B.n222 163.367
R838 B.n380 B.n222 163.367
R839 B.n380 B.n220 163.367
R840 B.n384 B.n220 163.367
R841 B.n384 B.n214 163.367
R842 B.n392 B.n214 163.367
R843 B.n392 B.n212 163.367
R844 B.n396 B.n212 163.367
R845 B.n396 B.n206 163.367
R846 B.n404 B.n206 163.367
R847 B.n404 B.n204 163.367
R848 B.n408 B.n204 163.367
R849 B.n408 B.n198 163.367
R850 B.n416 B.n198 163.367
R851 B.n416 B.n196 163.367
R852 B.n420 B.n196 163.367
R853 B.n420 B.n190 163.367
R854 B.n429 B.n190 163.367
R855 B.n429 B.n188 163.367
R856 B.n433 B.n188 163.367
R857 B.n433 B.n183 163.367
R858 B.n441 B.n183 163.367
R859 B.n441 B.n181 163.367
R860 B.n445 B.n181 163.367
R861 B.n445 B.n175 163.367
R862 B.n454 B.n175 163.367
R863 B.n454 B.n173 163.367
R864 B.n458 B.n173 163.367
R865 B.n458 B.n3 163.367
R866 B.n600 B.n3 163.367
R867 B.n596 B.n2 163.367
R868 B.n596 B.n595 163.367
R869 B.n595 B.n9 163.367
R870 B.n591 B.n9 163.367
R871 B.n591 B.n11 163.367
R872 B.n587 B.n11 163.367
R873 B.n587 B.n17 163.367
R874 B.n583 B.n17 163.367
R875 B.n583 B.n19 163.367
R876 B.n579 B.n19 163.367
R877 B.n579 B.n23 163.367
R878 B.n575 B.n23 163.367
R879 B.n575 B.n25 163.367
R880 B.n571 B.n25 163.367
R881 B.n571 B.n31 163.367
R882 B.n567 B.n31 163.367
R883 B.n567 B.n33 163.367
R884 B.n563 B.n33 163.367
R885 B.n563 B.n38 163.367
R886 B.n559 B.n38 163.367
R887 B.n559 B.n40 163.367
R888 B.n555 B.n40 163.367
R889 B.n555 B.n45 163.367
R890 B.n551 B.n45 163.367
R891 B.n551 B.n47 163.367
R892 B.n547 B.n47 163.367
R893 B.n547 B.n52 163.367
R894 B.n543 B.n52 163.367
R895 B.n543 B.n54 163.367
R896 B.n539 B.n54 163.367
R897 B.n539 B.n59 163.367
R898 B.n535 B.n59 163.367
R899 B.n535 B.n61 163.367
R900 B.n531 B.n61 163.367
R901 B.n531 B.n66 163.367
R902 B.n527 B.n66 163.367
R903 B.n527 B.n68 163.367
R904 B.n523 B.n68 163.367
R905 B.n523 B.n73 163.367
R906 B.n96 B.t11 124.832
R907 B.n269 B.t17 124.832
R908 B.n99 B.t14 124.832
R909 B.n267 B.t20 124.832
R910 B.n349 B.n243 94.8642
R911 B.n349 B.n239 94.8642
R912 B.n355 B.n239 94.8642
R913 B.n355 B.n234 94.8642
R914 B.n361 B.n234 94.8642
R915 B.n361 B.n235 94.8642
R916 B.n367 B.n227 94.8642
R917 B.n373 B.n227 94.8642
R918 B.n373 B.n223 94.8642
R919 B.n379 B.n223 94.8642
R920 B.n379 B.n219 94.8642
R921 B.n385 B.n219 94.8642
R922 B.n385 B.n215 94.8642
R923 B.n391 B.n215 94.8642
R924 B.n397 B.n211 94.8642
R925 B.n397 B.n207 94.8642
R926 B.n403 B.n207 94.8642
R927 B.n403 B.n202 94.8642
R928 B.n409 B.n202 94.8642
R929 B.n409 B.n203 94.8642
R930 B.n415 B.n195 94.8642
R931 B.n421 B.n195 94.8642
R932 B.n421 B.n191 94.8642
R933 B.n428 B.n191 94.8642
R934 B.n428 B.n427 94.8642
R935 B.n434 B.n184 94.8642
R936 B.n440 B.n184 94.8642
R937 B.n440 B.n179 94.8642
R938 B.n446 B.n179 94.8642
R939 B.n446 B.n180 94.8642
R940 B.n453 B.n172 94.8642
R941 B.n459 B.n172 94.8642
R942 B.n459 B.n4 94.8642
R943 B.n599 B.n4 94.8642
R944 B.n599 B.n598 94.8642
R945 B.n598 B.n597 94.8642
R946 B.n597 B.n8 94.8642
R947 B.n12 B.n8 94.8642
R948 B.n590 B.n12 94.8642
R949 B.n589 B.n588 94.8642
R950 B.n588 B.n16 94.8642
R951 B.n582 B.n16 94.8642
R952 B.n582 B.n581 94.8642
R953 B.n581 B.n580 94.8642
R954 B.n574 B.n26 94.8642
R955 B.n574 B.n573 94.8642
R956 B.n573 B.n572 94.8642
R957 B.n572 B.n30 94.8642
R958 B.n566 B.n30 94.8642
R959 B.n565 B.n564 94.8642
R960 B.n564 B.n37 94.8642
R961 B.n558 B.n37 94.8642
R962 B.n558 B.n557 94.8642
R963 B.n557 B.n556 94.8642
R964 B.n556 B.n44 94.8642
R965 B.n550 B.n549 94.8642
R966 B.n549 B.n548 94.8642
R967 B.n548 B.n51 94.8642
R968 B.n542 B.n51 94.8642
R969 B.n542 B.n541 94.8642
R970 B.n541 B.n540 94.8642
R971 B.n540 B.n58 94.8642
R972 B.n534 B.n58 94.8642
R973 B.n533 B.n532 94.8642
R974 B.n532 B.n65 94.8642
R975 B.n526 B.n65 94.8642
R976 B.n526 B.n525 94.8642
R977 B.n525 B.n524 94.8642
R978 B.n524 B.n72 94.8642
R979 B.n415 B.t7 86.4938
R980 B.n566 B.t1 86.4938
R981 B.n367 B.t16 72.5433
R982 B.n391 B.t0 72.5433
R983 B.n550 B.t3 72.5433
R984 B.n534 B.t9 72.5433
R985 B.n519 B.n518 71.676
R986 B.n101 B.n76 71.676
R987 B.n105 B.n77 71.676
R988 B.n109 B.n78 71.676
R989 B.n113 B.n79 71.676
R990 B.n117 B.n80 71.676
R991 B.n121 B.n81 71.676
R992 B.n125 B.n82 71.676
R993 B.n129 B.n83 71.676
R994 B.n133 B.n84 71.676
R995 B.n137 B.n85 71.676
R996 B.n141 B.n86 71.676
R997 B.n145 B.n87 71.676
R998 B.n149 B.n88 71.676
R999 B.n153 B.n89 71.676
R1000 B.n157 B.n90 71.676
R1001 B.n161 B.n91 71.676
R1002 B.n165 B.n92 71.676
R1003 B.n516 B.n93 71.676
R1004 B.n516 B.n515 71.676
R1005 B.n167 B.n92 71.676
R1006 B.n164 B.n91 71.676
R1007 B.n160 B.n90 71.676
R1008 B.n156 B.n89 71.676
R1009 B.n152 B.n88 71.676
R1010 B.n148 B.n87 71.676
R1011 B.n144 B.n86 71.676
R1012 B.n140 B.n85 71.676
R1013 B.n136 B.n84 71.676
R1014 B.n132 B.n83 71.676
R1015 B.n128 B.n82 71.676
R1016 B.n124 B.n81 71.676
R1017 B.n120 B.n80 71.676
R1018 B.n116 B.n79 71.676
R1019 B.n112 B.n78 71.676
R1020 B.n108 B.n77 71.676
R1021 B.n104 B.n76 71.676
R1022 B.n518 B.n75 71.676
R1023 B.n344 B.n343 71.676
R1024 B.n265 B.n247 71.676
R1025 B.n336 B.n248 71.676
R1026 B.n332 B.n249 71.676
R1027 B.n328 B.n250 71.676
R1028 B.n324 B.n251 71.676
R1029 B.n320 B.n252 71.676
R1030 B.n315 B.n253 71.676
R1031 B.n311 B.n254 71.676
R1032 B.n307 B.n255 71.676
R1033 B.n303 B.n256 71.676
R1034 B.n299 B.n257 71.676
R1035 B.n294 B.n258 71.676
R1036 B.n290 B.n259 71.676
R1037 B.n286 B.n260 71.676
R1038 B.n282 B.n261 71.676
R1039 B.n278 B.n262 71.676
R1040 B.n274 B.n263 71.676
R1041 B.n343 B.n246 71.676
R1042 B.n337 B.n247 71.676
R1043 B.n333 B.n248 71.676
R1044 B.n329 B.n249 71.676
R1045 B.n325 B.n250 71.676
R1046 B.n321 B.n251 71.676
R1047 B.n316 B.n252 71.676
R1048 B.n312 B.n253 71.676
R1049 B.n308 B.n254 71.676
R1050 B.n304 B.n255 71.676
R1051 B.n300 B.n256 71.676
R1052 B.n295 B.n257 71.676
R1053 B.n291 B.n258 71.676
R1054 B.n287 B.n259 71.676
R1055 B.n283 B.n260 71.676
R1056 B.n279 B.n261 71.676
R1057 B.n275 B.n262 71.676
R1058 B.n271 B.n263 71.676
R1059 B.n601 B.n600 71.676
R1060 B.n601 B.n2 71.676
R1061 B.n180 B.t5 69.7532
R1062 B.t2 B.n589 69.7532
R1063 B.n100 B.n99 59.5399
R1064 B.n97 B.n96 59.5399
R1065 B.n297 B.n269 59.5399
R1066 B.n318 B.n267 59.5399
R1067 B.n434 B.t6 55.8027
R1068 B.n580 B.t4 55.8027
R1069 B.n99 B.n98 41.6975
R1070 B.n96 B.n95 41.6975
R1071 B.n269 B.n268 41.6975
R1072 B.n267 B.n266 41.6975
R1073 B.n427 B.t6 39.062
R1074 B.n26 B.t4 39.062
R1075 B.n346 B.n345 32.6249
R1076 B.n270 B.n241 32.6249
R1077 B.n514 B.n513 32.6249
R1078 B.n521 B.n520 32.6249
R1079 B.n453 B.t5 25.1115
R1080 B.n590 B.t2 25.1115
R1081 B.n235 B.t16 22.3214
R1082 B.t0 B.n211 22.3214
R1083 B.t3 B.n44 22.3214
R1084 B.t9 B.n533 22.3214
R1085 B B.n602 18.0485
R1086 B.n347 B.n346 10.6151
R1087 B.n347 B.n237 10.6151
R1088 B.n357 B.n237 10.6151
R1089 B.n358 B.n357 10.6151
R1090 B.n359 B.n358 10.6151
R1091 B.n359 B.n229 10.6151
R1092 B.n369 B.n229 10.6151
R1093 B.n370 B.n369 10.6151
R1094 B.n371 B.n370 10.6151
R1095 B.n371 B.n221 10.6151
R1096 B.n381 B.n221 10.6151
R1097 B.n382 B.n381 10.6151
R1098 B.n383 B.n382 10.6151
R1099 B.n383 B.n213 10.6151
R1100 B.n393 B.n213 10.6151
R1101 B.n394 B.n393 10.6151
R1102 B.n395 B.n394 10.6151
R1103 B.n395 B.n205 10.6151
R1104 B.n405 B.n205 10.6151
R1105 B.n406 B.n405 10.6151
R1106 B.n407 B.n406 10.6151
R1107 B.n407 B.n197 10.6151
R1108 B.n417 B.n197 10.6151
R1109 B.n418 B.n417 10.6151
R1110 B.n419 B.n418 10.6151
R1111 B.n419 B.n189 10.6151
R1112 B.n430 B.n189 10.6151
R1113 B.n431 B.n430 10.6151
R1114 B.n432 B.n431 10.6151
R1115 B.n432 B.n182 10.6151
R1116 B.n442 B.n182 10.6151
R1117 B.n443 B.n442 10.6151
R1118 B.n444 B.n443 10.6151
R1119 B.n444 B.n174 10.6151
R1120 B.n455 B.n174 10.6151
R1121 B.n456 B.n455 10.6151
R1122 B.n457 B.n456 10.6151
R1123 B.n457 B.n0 10.6151
R1124 B.n345 B.n245 10.6151
R1125 B.n340 B.n245 10.6151
R1126 B.n340 B.n339 10.6151
R1127 B.n339 B.n338 10.6151
R1128 B.n338 B.n335 10.6151
R1129 B.n335 B.n334 10.6151
R1130 B.n334 B.n331 10.6151
R1131 B.n331 B.n330 10.6151
R1132 B.n330 B.n327 10.6151
R1133 B.n327 B.n326 10.6151
R1134 B.n326 B.n323 10.6151
R1135 B.n323 B.n322 10.6151
R1136 B.n322 B.n319 10.6151
R1137 B.n317 B.n314 10.6151
R1138 B.n314 B.n313 10.6151
R1139 B.n313 B.n310 10.6151
R1140 B.n310 B.n309 10.6151
R1141 B.n309 B.n306 10.6151
R1142 B.n306 B.n305 10.6151
R1143 B.n305 B.n302 10.6151
R1144 B.n302 B.n301 10.6151
R1145 B.n301 B.n298 10.6151
R1146 B.n296 B.n293 10.6151
R1147 B.n293 B.n292 10.6151
R1148 B.n292 B.n289 10.6151
R1149 B.n289 B.n288 10.6151
R1150 B.n288 B.n285 10.6151
R1151 B.n285 B.n284 10.6151
R1152 B.n284 B.n281 10.6151
R1153 B.n281 B.n280 10.6151
R1154 B.n280 B.n277 10.6151
R1155 B.n277 B.n276 10.6151
R1156 B.n276 B.n273 10.6151
R1157 B.n273 B.n272 10.6151
R1158 B.n272 B.n270 10.6151
R1159 B.n351 B.n241 10.6151
R1160 B.n352 B.n351 10.6151
R1161 B.n353 B.n352 10.6151
R1162 B.n353 B.n232 10.6151
R1163 B.n363 B.n232 10.6151
R1164 B.n364 B.n363 10.6151
R1165 B.n365 B.n364 10.6151
R1166 B.n365 B.n225 10.6151
R1167 B.n375 B.n225 10.6151
R1168 B.n376 B.n375 10.6151
R1169 B.n377 B.n376 10.6151
R1170 B.n377 B.n217 10.6151
R1171 B.n387 B.n217 10.6151
R1172 B.n388 B.n387 10.6151
R1173 B.n389 B.n388 10.6151
R1174 B.n389 B.n209 10.6151
R1175 B.n399 B.n209 10.6151
R1176 B.n400 B.n399 10.6151
R1177 B.n401 B.n400 10.6151
R1178 B.n401 B.n200 10.6151
R1179 B.n411 B.n200 10.6151
R1180 B.n412 B.n411 10.6151
R1181 B.n413 B.n412 10.6151
R1182 B.n413 B.n193 10.6151
R1183 B.n423 B.n193 10.6151
R1184 B.n424 B.n423 10.6151
R1185 B.n425 B.n424 10.6151
R1186 B.n425 B.n186 10.6151
R1187 B.n436 B.n186 10.6151
R1188 B.n437 B.n436 10.6151
R1189 B.n438 B.n437 10.6151
R1190 B.n438 B.n177 10.6151
R1191 B.n448 B.n177 10.6151
R1192 B.n449 B.n448 10.6151
R1193 B.n451 B.n449 10.6151
R1194 B.n451 B.n450 10.6151
R1195 B.n450 B.n170 10.6151
R1196 B.n462 B.n170 10.6151
R1197 B.n463 B.n462 10.6151
R1198 B.n464 B.n463 10.6151
R1199 B.n465 B.n464 10.6151
R1200 B.n466 B.n465 10.6151
R1201 B.n469 B.n466 10.6151
R1202 B.n470 B.n469 10.6151
R1203 B.n471 B.n470 10.6151
R1204 B.n472 B.n471 10.6151
R1205 B.n474 B.n472 10.6151
R1206 B.n475 B.n474 10.6151
R1207 B.n476 B.n475 10.6151
R1208 B.n477 B.n476 10.6151
R1209 B.n479 B.n477 10.6151
R1210 B.n480 B.n479 10.6151
R1211 B.n481 B.n480 10.6151
R1212 B.n482 B.n481 10.6151
R1213 B.n484 B.n482 10.6151
R1214 B.n485 B.n484 10.6151
R1215 B.n486 B.n485 10.6151
R1216 B.n487 B.n486 10.6151
R1217 B.n489 B.n487 10.6151
R1218 B.n490 B.n489 10.6151
R1219 B.n491 B.n490 10.6151
R1220 B.n492 B.n491 10.6151
R1221 B.n494 B.n492 10.6151
R1222 B.n495 B.n494 10.6151
R1223 B.n496 B.n495 10.6151
R1224 B.n497 B.n496 10.6151
R1225 B.n499 B.n497 10.6151
R1226 B.n500 B.n499 10.6151
R1227 B.n501 B.n500 10.6151
R1228 B.n502 B.n501 10.6151
R1229 B.n504 B.n502 10.6151
R1230 B.n505 B.n504 10.6151
R1231 B.n506 B.n505 10.6151
R1232 B.n507 B.n506 10.6151
R1233 B.n509 B.n507 10.6151
R1234 B.n510 B.n509 10.6151
R1235 B.n511 B.n510 10.6151
R1236 B.n512 B.n511 10.6151
R1237 B.n513 B.n512 10.6151
R1238 B.n594 B.n1 10.6151
R1239 B.n594 B.n593 10.6151
R1240 B.n593 B.n592 10.6151
R1241 B.n592 B.n10 10.6151
R1242 B.n586 B.n10 10.6151
R1243 B.n586 B.n585 10.6151
R1244 B.n585 B.n584 10.6151
R1245 B.n584 B.n18 10.6151
R1246 B.n578 B.n18 10.6151
R1247 B.n578 B.n577 10.6151
R1248 B.n577 B.n576 10.6151
R1249 B.n576 B.n24 10.6151
R1250 B.n570 B.n24 10.6151
R1251 B.n570 B.n569 10.6151
R1252 B.n569 B.n568 10.6151
R1253 B.n568 B.n32 10.6151
R1254 B.n562 B.n32 10.6151
R1255 B.n562 B.n561 10.6151
R1256 B.n561 B.n560 10.6151
R1257 B.n560 B.n39 10.6151
R1258 B.n554 B.n39 10.6151
R1259 B.n554 B.n553 10.6151
R1260 B.n553 B.n552 10.6151
R1261 B.n552 B.n46 10.6151
R1262 B.n546 B.n46 10.6151
R1263 B.n546 B.n545 10.6151
R1264 B.n545 B.n544 10.6151
R1265 B.n544 B.n53 10.6151
R1266 B.n538 B.n53 10.6151
R1267 B.n538 B.n537 10.6151
R1268 B.n537 B.n536 10.6151
R1269 B.n536 B.n60 10.6151
R1270 B.n530 B.n60 10.6151
R1271 B.n530 B.n529 10.6151
R1272 B.n529 B.n528 10.6151
R1273 B.n528 B.n67 10.6151
R1274 B.n522 B.n67 10.6151
R1275 B.n522 B.n521 10.6151
R1276 B.n520 B.n74 10.6151
R1277 B.n102 B.n74 10.6151
R1278 B.n103 B.n102 10.6151
R1279 B.n106 B.n103 10.6151
R1280 B.n107 B.n106 10.6151
R1281 B.n110 B.n107 10.6151
R1282 B.n111 B.n110 10.6151
R1283 B.n114 B.n111 10.6151
R1284 B.n115 B.n114 10.6151
R1285 B.n118 B.n115 10.6151
R1286 B.n119 B.n118 10.6151
R1287 B.n122 B.n119 10.6151
R1288 B.n123 B.n122 10.6151
R1289 B.n127 B.n126 10.6151
R1290 B.n130 B.n127 10.6151
R1291 B.n131 B.n130 10.6151
R1292 B.n134 B.n131 10.6151
R1293 B.n135 B.n134 10.6151
R1294 B.n138 B.n135 10.6151
R1295 B.n139 B.n138 10.6151
R1296 B.n142 B.n139 10.6151
R1297 B.n143 B.n142 10.6151
R1298 B.n147 B.n146 10.6151
R1299 B.n150 B.n147 10.6151
R1300 B.n151 B.n150 10.6151
R1301 B.n154 B.n151 10.6151
R1302 B.n155 B.n154 10.6151
R1303 B.n158 B.n155 10.6151
R1304 B.n159 B.n158 10.6151
R1305 B.n162 B.n159 10.6151
R1306 B.n163 B.n162 10.6151
R1307 B.n166 B.n163 10.6151
R1308 B.n168 B.n166 10.6151
R1309 B.n169 B.n168 10.6151
R1310 B.n514 B.n169 10.6151
R1311 B.n319 B.n318 9.36635
R1312 B.n297 B.n296 9.36635
R1313 B.n123 B.n100 9.36635
R1314 B.n146 B.n97 9.36635
R1315 B.n203 B.t7 8.37082
R1316 B.t1 B.n565 8.37082
R1317 B.n602 B.n0 8.11757
R1318 B.n602 B.n1 8.11757
R1319 B.n318 B.n317 1.24928
R1320 B.n298 B.n297 1.24928
R1321 B.n126 B.n100 1.24928
R1322 B.n143 B.n97 1.24928
R1323 VN.n39 VN.n21 161.3
R1324 VN.n38 VN.n37 161.3
R1325 VN.n36 VN.n22 161.3
R1326 VN.n35 VN.n34 161.3
R1327 VN.n32 VN.n23 161.3
R1328 VN.n31 VN.n30 161.3
R1329 VN.n29 VN.n24 161.3
R1330 VN.n28 VN.n27 161.3
R1331 VN.n18 VN.n0 161.3
R1332 VN.n17 VN.n16 161.3
R1333 VN.n15 VN.n1 161.3
R1334 VN.n14 VN.n13 161.3
R1335 VN.n11 VN.n2 161.3
R1336 VN.n10 VN.n9 161.3
R1337 VN.n8 VN.n3 161.3
R1338 VN.n7 VN.n6 161.3
R1339 VN.n20 VN.n19 87.5128
R1340 VN.n41 VN.n40 87.5128
R1341 VN.n4 VN.t6 65.9947
R1342 VN.n25 VN.t4 65.9947
R1343 VN.n10 VN.n3 56.5193
R1344 VN.n31 VN.n24 56.5193
R1345 VN.n5 VN.n4 53.8955
R1346 VN.n26 VN.n25 53.8955
R1347 VN.n17 VN.n1 50.2061
R1348 VN.n38 VN.n22 50.2061
R1349 VN VN.n41 40.4451
R1350 VN.n5 VN.t7 34.5615
R1351 VN.n12 VN.t2 34.5615
R1352 VN.n19 VN.t3 34.5615
R1353 VN.n26 VN.t5 34.5615
R1354 VN.n33 VN.t0 34.5615
R1355 VN.n40 VN.t1 34.5615
R1356 VN.n18 VN.n17 30.7807
R1357 VN.n39 VN.n38 30.7807
R1358 VN.n6 VN.n3 24.4675
R1359 VN.n11 VN.n10 24.4675
R1360 VN.n13 VN.n1 24.4675
R1361 VN.n27 VN.n24 24.4675
R1362 VN.n34 VN.n22 24.4675
R1363 VN.n32 VN.n31 24.4675
R1364 VN.n19 VN.n18 23.2442
R1365 VN.n40 VN.n39 23.2442
R1366 VN.n6 VN.n5 15.9041
R1367 VN.n12 VN.n11 15.9041
R1368 VN.n27 VN.n26 15.9041
R1369 VN.n33 VN.n32 15.9041
R1370 VN.n28 VN.n25 12.7761
R1371 VN.n7 VN.n4 12.7761
R1372 VN.n13 VN.n12 8.56395
R1373 VN.n34 VN.n33 8.56395
R1374 VN.n41 VN.n21 0.278367
R1375 VN.n20 VN.n0 0.278367
R1376 VN.n37 VN.n21 0.189894
R1377 VN.n37 VN.n36 0.189894
R1378 VN.n36 VN.n35 0.189894
R1379 VN.n35 VN.n23 0.189894
R1380 VN.n30 VN.n23 0.189894
R1381 VN.n30 VN.n29 0.189894
R1382 VN.n29 VN.n28 0.189894
R1383 VN.n8 VN.n7 0.189894
R1384 VN.n9 VN.n8 0.189894
R1385 VN.n9 VN.n2 0.189894
R1386 VN.n14 VN.n2 0.189894
R1387 VN.n15 VN.n14 0.189894
R1388 VN.n16 VN.n15 0.189894
R1389 VN.n16 VN.n0 0.189894
R1390 VN VN.n20 0.153454
R1391 VDD2.n2 VDD2.n1 89.9033
R1392 VDD2.n2 VDD2.n0 89.9033
R1393 VDD2 VDD2.n5 89.9004
R1394 VDD2.n4 VDD2.n3 89.032
R1395 VDD2.n4 VDD2.n2 34.3058
R1396 VDD2.n5 VDD2.t2 7.58671
R1397 VDD2.n5 VDD2.t3 7.58671
R1398 VDD2.n3 VDD2.t6 7.58671
R1399 VDD2.n3 VDD2.t7 7.58671
R1400 VDD2.n1 VDD2.t5 7.58671
R1401 VDD2.n1 VDD2.t4 7.58671
R1402 VDD2.n0 VDD2.t1 7.58671
R1403 VDD2.n0 VDD2.t0 7.58671
R1404 VDD2 VDD2.n4 0.985414
C0 VN VTAIL 2.80139f
C1 VN VP 4.97887f
C2 VDD2 VTAIL 4.36573f
C3 VDD1 VTAIL 4.31654f
C4 VDD2 VP 0.442562f
C5 VDD1 VP 2.36704f
C6 VDD2 VN 2.08185f
C7 VDD1 VN 0.155405f
C8 VDD2 VDD1 1.3704f
C9 VP VTAIL 2.8155f
C10 VDD2 B 3.8428f
C11 VDD1 B 4.200875f
C12 VTAIL B 4.056247f
C13 VN B 11.67113f
C14 VP B 10.206487f
C15 VDD2.t1 B 0.050759f
C16 VDD2.t0 B 0.050759f
C17 VDD2.n0 B 0.365568f
C18 VDD2.t5 B 0.050759f
C19 VDD2.t4 B 0.050759f
C20 VDD2.n1 B 0.365568f
C21 VDD2.n2 B 2.19063f
C22 VDD2.t6 B 0.050759f
C23 VDD2.t7 B 0.050759f
C24 VDD2.n3 B 0.361589f
C25 VDD2.n4 B 1.89221f
C26 VDD2.t2 B 0.050759f
C27 VDD2.t3 B 0.050759f
C28 VDD2.n5 B 0.365547f
C29 VN.n0 B 0.044442f
C30 VN.t3 B 0.391431f
C31 VN.n1 B 0.061868f
C32 VN.n2 B 0.033709f
C33 VN.t2 B 0.391431f
C34 VN.n3 B 0.049209f
C35 VN.t6 B 0.552646f
C36 VN.n4 B 0.249108f
C37 VN.t7 B 0.391431f
C38 VN.n5 B 0.260766f
C39 VN.n6 B 0.051967f
C40 VN.n7 B 0.246957f
C41 VN.n8 B 0.033709f
C42 VN.n9 B 0.033709f
C43 VN.n10 B 0.049209f
C44 VN.n11 B 0.051967f
C45 VN.n12 B 0.180595f
C46 VN.n13 B 0.042662f
C47 VN.n14 B 0.033709f
C48 VN.n15 B 0.033709f
C49 VN.n16 B 0.033709f
C50 VN.n17 B 0.031844f
C51 VN.n18 B 0.065978f
C52 VN.n19 B 0.281613f
C53 VN.n20 B 0.036646f
C54 VN.n21 B 0.044442f
C55 VN.t1 B 0.391431f
C56 VN.n22 B 0.061868f
C57 VN.n23 B 0.033709f
C58 VN.t0 B 0.391431f
C59 VN.n24 B 0.049209f
C60 VN.t4 B 0.552646f
C61 VN.n25 B 0.249108f
C62 VN.t5 B 0.391431f
C63 VN.n26 B 0.260766f
C64 VN.n27 B 0.051967f
C65 VN.n28 B 0.246957f
C66 VN.n29 B 0.033709f
C67 VN.n30 B 0.033709f
C68 VN.n31 B 0.049209f
C69 VN.n32 B 0.051967f
C70 VN.n33 B 0.180595f
C71 VN.n34 B 0.042662f
C72 VN.n35 B 0.033709f
C73 VN.n36 B 0.033709f
C74 VN.n37 B 0.033709f
C75 VN.n38 B 0.031844f
C76 VN.n39 B 0.065978f
C77 VN.n40 B 0.281613f
C78 VN.n41 B 1.33266f
C79 VTAIL.t4 B 0.056712f
C80 VTAIL.t1 B 0.056712f
C81 VTAIL.n0 B 0.357804f
C82 VTAIL.n1 B 0.383788f
C83 VTAIL.n2 B 0.038835f
C84 VTAIL.n3 B 0.21693f
C85 VTAIL.n4 B 0.014776f
C86 VTAIL.t2 B 0.061639f
C87 VTAIL.n5 B 0.100246f
C88 VTAIL.n6 B 0.01977f
C89 VTAIL.n7 B 0.026193f
C90 VTAIL.n8 B 0.075933f
C91 VTAIL.n9 B 0.015645f
C92 VTAIL.n10 B 0.014776f
C93 VTAIL.n11 B 0.071446f
C94 VTAIL.n12 B 0.042751f
C95 VTAIL.n13 B 0.233793f
C96 VTAIL.n14 B 0.038835f
C97 VTAIL.n15 B 0.21693f
C98 VTAIL.n16 B 0.014776f
C99 VTAIL.t10 B 0.061639f
C100 VTAIL.n17 B 0.100246f
C101 VTAIL.n18 B 0.01977f
C102 VTAIL.n19 B 0.026193f
C103 VTAIL.n20 B 0.075933f
C104 VTAIL.n21 B 0.015645f
C105 VTAIL.n22 B 0.014776f
C106 VTAIL.n23 B 0.071446f
C107 VTAIL.n24 B 0.042751f
C108 VTAIL.n25 B 0.233793f
C109 VTAIL.t11 B 0.056712f
C110 VTAIL.t8 B 0.056712f
C111 VTAIL.n26 B 0.357804f
C112 VTAIL.n27 B 0.54285f
C113 VTAIL.n28 B 0.038835f
C114 VTAIL.n29 B 0.21693f
C115 VTAIL.n30 B 0.014776f
C116 VTAIL.t9 B 0.061639f
C117 VTAIL.n31 B 0.100246f
C118 VTAIL.n32 B 0.01977f
C119 VTAIL.n33 B 0.026193f
C120 VTAIL.n34 B 0.075933f
C121 VTAIL.n35 B 0.015645f
C122 VTAIL.n36 B 0.014776f
C123 VTAIL.n37 B 0.071446f
C124 VTAIL.n38 B 0.042751f
C125 VTAIL.n39 B 0.929248f
C126 VTAIL.n40 B 0.038835f
C127 VTAIL.n41 B 0.21693f
C128 VTAIL.n42 B 0.014776f
C129 VTAIL.t0 B 0.061639f
C130 VTAIL.n43 B 0.100246f
C131 VTAIL.n44 B 0.01977f
C132 VTAIL.n45 B 0.026193f
C133 VTAIL.n46 B 0.075933f
C134 VTAIL.n47 B 0.015645f
C135 VTAIL.n48 B 0.014776f
C136 VTAIL.n49 B 0.071446f
C137 VTAIL.n50 B 0.042751f
C138 VTAIL.n51 B 0.929248f
C139 VTAIL.t7 B 0.056712f
C140 VTAIL.t6 B 0.056712f
C141 VTAIL.n52 B 0.357806f
C142 VTAIL.n53 B 0.542848f
C143 VTAIL.n54 B 0.038835f
C144 VTAIL.n55 B 0.21693f
C145 VTAIL.n56 B 0.014776f
C146 VTAIL.t5 B 0.061639f
C147 VTAIL.n57 B 0.100246f
C148 VTAIL.n58 B 0.01977f
C149 VTAIL.n59 B 0.026193f
C150 VTAIL.n60 B 0.075933f
C151 VTAIL.n61 B 0.015645f
C152 VTAIL.n62 B 0.014776f
C153 VTAIL.n63 B 0.071446f
C154 VTAIL.n64 B 0.042751f
C155 VTAIL.n65 B 0.233793f
C156 VTAIL.n66 B 0.038835f
C157 VTAIL.n67 B 0.21693f
C158 VTAIL.n68 B 0.014776f
C159 VTAIL.t14 B 0.061639f
C160 VTAIL.n69 B 0.100246f
C161 VTAIL.n70 B 0.01977f
C162 VTAIL.n71 B 0.026193f
C163 VTAIL.n72 B 0.075933f
C164 VTAIL.n73 B 0.015645f
C165 VTAIL.n74 B 0.014776f
C166 VTAIL.n75 B 0.071446f
C167 VTAIL.n76 B 0.042751f
C168 VTAIL.n77 B 0.233793f
C169 VTAIL.t12 B 0.056712f
C170 VTAIL.t15 B 0.056712f
C171 VTAIL.n78 B 0.357806f
C172 VTAIL.n79 B 0.542848f
C173 VTAIL.n80 B 0.038835f
C174 VTAIL.n81 B 0.21693f
C175 VTAIL.n82 B 0.014776f
C176 VTAIL.t13 B 0.061639f
C177 VTAIL.n83 B 0.100246f
C178 VTAIL.n84 B 0.01977f
C179 VTAIL.n85 B 0.026193f
C180 VTAIL.n86 B 0.075933f
C181 VTAIL.n87 B 0.015645f
C182 VTAIL.n88 B 0.014776f
C183 VTAIL.n89 B 0.071446f
C184 VTAIL.n90 B 0.042751f
C185 VTAIL.n91 B 0.929248f
C186 VTAIL.n92 B 0.038835f
C187 VTAIL.n93 B 0.21693f
C188 VTAIL.n94 B 0.014776f
C189 VTAIL.t3 B 0.061639f
C190 VTAIL.n95 B 0.100246f
C191 VTAIL.n96 B 0.01977f
C192 VTAIL.n97 B 0.026193f
C193 VTAIL.n98 B 0.075933f
C194 VTAIL.n99 B 0.015645f
C195 VTAIL.n100 B 0.014776f
C196 VTAIL.n101 B 0.071446f
C197 VTAIL.n102 B 0.042751f
C198 VTAIL.n103 B 0.924092f
C199 VDD1.t1 B 0.0516f
C200 VDD1.t5 B 0.0516f
C201 VDD1.n0 B 0.372235f
C202 VDD1.t2 B 0.0516f
C203 VDD1.t7 B 0.0516f
C204 VDD1.n1 B 0.371619f
C205 VDD1.t3 B 0.0516f
C206 VDD1.t0 B 0.0516f
C207 VDD1.n2 B 0.371619f
C208 VDD1.n3 B 2.2797f
C209 VDD1.t4 B 0.0516f
C210 VDD1.t6 B 0.0516f
C211 VDD1.n4 B 0.367573f
C212 VDD1.n5 B 1.95375f
C213 VP.n0 B 0.046009f
C214 VP.t5 B 0.405233f
C215 VP.n1 B 0.064049f
C216 VP.n2 B 0.034897f
C217 VP.t7 B 0.405233f
C218 VP.n3 B 0.050944f
C219 VP.n4 B 0.034897f
C220 VP.t4 B 0.405233f
C221 VP.n5 B 0.032967f
C222 VP.n6 B 0.046009f
C223 VP.t2 B 0.405233f
C224 VP.n7 B 0.064049f
C225 VP.n8 B 0.034897f
C226 VP.t0 B 0.405233f
C227 VP.n9 B 0.050944f
C228 VP.t1 B 0.572132f
C229 VP.n10 B 0.257891f
C230 VP.t3 B 0.405233f
C231 VP.n11 B 0.26996f
C232 VP.n12 B 0.0538f
C233 VP.n13 B 0.255665f
C234 VP.n14 B 0.034897f
C235 VP.n15 B 0.034897f
C236 VP.n16 B 0.050944f
C237 VP.n17 B 0.0538f
C238 VP.n18 B 0.186962f
C239 VP.n19 B 0.044166f
C240 VP.n20 B 0.034897f
C241 VP.n21 B 0.034897f
C242 VP.n22 B 0.034897f
C243 VP.n23 B 0.032967f
C244 VP.n24 B 0.068304f
C245 VP.n25 B 0.291542f
C246 VP.n26 B 1.36017f
C247 VP.n27 B 1.3914f
C248 VP.t6 B 0.405233f
C249 VP.n28 B 0.291542f
C250 VP.n29 B 0.068304f
C251 VP.n30 B 0.046009f
C252 VP.n31 B 0.034897f
C253 VP.n32 B 0.034897f
C254 VP.n33 B 0.064049f
C255 VP.n34 B 0.044166f
C256 VP.n35 B 0.186962f
C257 VP.n36 B 0.0538f
C258 VP.n37 B 0.034897f
C259 VP.n38 B 0.034897f
C260 VP.n39 B 0.034897f
C261 VP.n40 B 0.050944f
C262 VP.n41 B 0.0538f
C263 VP.n42 B 0.186962f
C264 VP.n43 B 0.044166f
C265 VP.n44 B 0.034897f
C266 VP.n45 B 0.034897f
C267 VP.n46 B 0.034897f
C268 VP.n47 B 0.032967f
C269 VP.n48 B 0.068304f
C270 VP.n49 B 0.291542f
C271 VP.n50 B 0.037938f
.ends

