* NGSPICE file created from diff_pair_sample_0679.ext - technology: sky130A

.subckt diff_pair_sample_0679 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=0 ps=0 w=10.24 l=2.78
X1 VDD1.t9 VP.t0 VTAIL.t10 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X2 B.t8 B.t6 B.t7 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=0 ps=0 w=10.24 l=2.78
X3 VDD2.t9 VN.t0 VTAIL.t7 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X4 B.t5 B.t3 B.t4 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=0 ps=0 w=10.24 l=2.78
X5 VDD2.t8 VN.t1 VTAIL.t9 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=1.6896 ps=10.57 w=10.24 l=2.78
X6 VTAIL.t3 VN.t2 VDD2.t7 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X7 VDD2.t6 VN.t3 VTAIL.t0 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=3.9936 ps=21.26 w=10.24 l=2.78
X8 VDD1.t8 VP.t1 VTAIL.t11 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=3.9936 ps=21.26 w=10.24 l=2.78
X9 VDD1.t7 VP.t2 VTAIL.t12 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=3.9936 ps=21.26 w=10.24 l=2.78
X10 VTAIL.t6 VN.t4 VDD2.t5 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X11 VDD1.t6 VP.t3 VTAIL.t13 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=1.6896 ps=10.57 w=10.24 l=2.78
X12 VDD2.t4 VN.t5 VTAIL.t2 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X13 VDD2.t3 VN.t6 VTAIL.t8 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=3.9936 ps=21.26 w=10.24 l=2.78
X14 VTAIL.t14 VP.t4 VDD1.t5 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X15 VTAIL.t15 VP.t5 VDD1.t4 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X16 VTAIL.t4 VN.t7 VDD2.t2 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X17 VDD2.t1 VN.t8 VTAIL.t1 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=1.6896 ps=10.57 w=10.24 l=2.78
X18 VDD1.t3 VP.t6 VTAIL.t16 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=1.6896 ps=10.57 w=10.24 l=2.78
X19 VTAIL.t17 VP.t7 VDD1.t2 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X20 VDD1.t1 VP.t8 VTAIL.t18 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X21 VTAIL.t19 VP.t9 VDD1.t0 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
X22 B.t2 B.t0 B.t1 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=3.9936 pd=21.26 as=0 ps=0 w=10.24 l=2.78
X23 VTAIL.t5 VN.t9 VDD2.t0 w_n4702_n3016# sky130_fd_pr__pfet_01v8 ad=1.6896 pd=10.57 as=1.6896 ps=10.57 w=10.24 l=2.78
R0 B.n628 B.n79 585
R1 B.n630 B.n629 585
R2 B.n631 B.n78 585
R3 B.n633 B.n632 585
R4 B.n634 B.n77 585
R5 B.n636 B.n635 585
R6 B.n637 B.n76 585
R7 B.n639 B.n638 585
R8 B.n640 B.n75 585
R9 B.n642 B.n641 585
R10 B.n643 B.n74 585
R11 B.n645 B.n644 585
R12 B.n646 B.n73 585
R13 B.n648 B.n647 585
R14 B.n649 B.n72 585
R15 B.n651 B.n650 585
R16 B.n652 B.n71 585
R17 B.n654 B.n653 585
R18 B.n655 B.n70 585
R19 B.n657 B.n656 585
R20 B.n658 B.n69 585
R21 B.n660 B.n659 585
R22 B.n661 B.n68 585
R23 B.n663 B.n662 585
R24 B.n664 B.n67 585
R25 B.n666 B.n665 585
R26 B.n667 B.n66 585
R27 B.n669 B.n668 585
R28 B.n670 B.n65 585
R29 B.n672 B.n671 585
R30 B.n673 B.n64 585
R31 B.n675 B.n674 585
R32 B.n676 B.n63 585
R33 B.n678 B.n677 585
R34 B.n679 B.n59 585
R35 B.n681 B.n680 585
R36 B.n682 B.n58 585
R37 B.n684 B.n683 585
R38 B.n685 B.n57 585
R39 B.n687 B.n686 585
R40 B.n688 B.n56 585
R41 B.n690 B.n689 585
R42 B.n691 B.n55 585
R43 B.n693 B.n692 585
R44 B.n694 B.n54 585
R45 B.n696 B.n695 585
R46 B.n698 B.n51 585
R47 B.n700 B.n699 585
R48 B.n701 B.n50 585
R49 B.n703 B.n702 585
R50 B.n704 B.n49 585
R51 B.n706 B.n705 585
R52 B.n707 B.n48 585
R53 B.n709 B.n708 585
R54 B.n710 B.n47 585
R55 B.n712 B.n711 585
R56 B.n713 B.n46 585
R57 B.n715 B.n714 585
R58 B.n716 B.n45 585
R59 B.n718 B.n717 585
R60 B.n719 B.n44 585
R61 B.n721 B.n720 585
R62 B.n722 B.n43 585
R63 B.n724 B.n723 585
R64 B.n725 B.n42 585
R65 B.n727 B.n726 585
R66 B.n728 B.n41 585
R67 B.n730 B.n729 585
R68 B.n731 B.n40 585
R69 B.n733 B.n732 585
R70 B.n734 B.n39 585
R71 B.n736 B.n735 585
R72 B.n737 B.n38 585
R73 B.n739 B.n738 585
R74 B.n740 B.n37 585
R75 B.n742 B.n741 585
R76 B.n743 B.n36 585
R77 B.n745 B.n744 585
R78 B.n746 B.n35 585
R79 B.n748 B.n747 585
R80 B.n749 B.n34 585
R81 B.n751 B.n750 585
R82 B.n627 B.n626 585
R83 B.n625 B.n80 585
R84 B.n624 B.n623 585
R85 B.n622 B.n81 585
R86 B.n621 B.n620 585
R87 B.n619 B.n82 585
R88 B.n618 B.n617 585
R89 B.n616 B.n83 585
R90 B.n615 B.n614 585
R91 B.n613 B.n84 585
R92 B.n612 B.n611 585
R93 B.n610 B.n85 585
R94 B.n609 B.n608 585
R95 B.n607 B.n86 585
R96 B.n606 B.n605 585
R97 B.n604 B.n87 585
R98 B.n603 B.n602 585
R99 B.n601 B.n88 585
R100 B.n600 B.n599 585
R101 B.n598 B.n89 585
R102 B.n597 B.n596 585
R103 B.n595 B.n90 585
R104 B.n594 B.n593 585
R105 B.n592 B.n91 585
R106 B.n591 B.n590 585
R107 B.n589 B.n92 585
R108 B.n588 B.n587 585
R109 B.n586 B.n93 585
R110 B.n585 B.n584 585
R111 B.n583 B.n94 585
R112 B.n582 B.n581 585
R113 B.n580 B.n95 585
R114 B.n579 B.n578 585
R115 B.n577 B.n96 585
R116 B.n576 B.n575 585
R117 B.n574 B.n97 585
R118 B.n573 B.n572 585
R119 B.n571 B.n98 585
R120 B.n570 B.n569 585
R121 B.n568 B.n99 585
R122 B.n567 B.n566 585
R123 B.n565 B.n100 585
R124 B.n564 B.n563 585
R125 B.n562 B.n101 585
R126 B.n561 B.n560 585
R127 B.n559 B.n102 585
R128 B.n558 B.n557 585
R129 B.n556 B.n103 585
R130 B.n555 B.n554 585
R131 B.n553 B.n104 585
R132 B.n552 B.n551 585
R133 B.n550 B.n105 585
R134 B.n549 B.n548 585
R135 B.n547 B.n106 585
R136 B.n546 B.n545 585
R137 B.n544 B.n107 585
R138 B.n543 B.n542 585
R139 B.n541 B.n108 585
R140 B.n540 B.n539 585
R141 B.n538 B.n109 585
R142 B.n537 B.n536 585
R143 B.n535 B.n110 585
R144 B.n534 B.n533 585
R145 B.n532 B.n111 585
R146 B.n531 B.n530 585
R147 B.n529 B.n112 585
R148 B.n528 B.n527 585
R149 B.n526 B.n113 585
R150 B.n525 B.n524 585
R151 B.n523 B.n114 585
R152 B.n522 B.n521 585
R153 B.n520 B.n115 585
R154 B.n519 B.n518 585
R155 B.n517 B.n116 585
R156 B.n516 B.n515 585
R157 B.n514 B.n117 585
R158 B.n513 B.n512 585
R159 B.n511 B.n118 585
R160 B.n510 B.n509 585
R161 B.n508 B.n119 585
R162 B.n507 B.n506 585
R163 B.n505 B.n120 585
R164 B.n504 B.n503 585
R165 B.n502 B.n121 585
R166 B.n501 B.n500 585
R167 B.n499 B.n122 585
R168 B.n498 B.n497 585
R169 B.n496 B.n123 585
R170 B.n495 B.n494 585
R171 B.n493 B.n124 585
R172 B.n492 B.n491 585
R173 B.n490 B.n125 585
R174 B.n489 B.n488 585
R175 B.n487 B.n126 585
R176 B.n486 B.n485 585
R177 B.n484 B.n127 585
R178 B.n483 B.n482 585
R179 B.n481 B.n128 585
R180 B.n480 B.n479 585
R181 B.n478 B.n129 585
R182 B.n477 B.n476 585
R183 B.n475 B.n130 585
R184 B.n474 B.n473 585
R185 B.n472 B.n131 585
R186 B.n471 B.n470 585
R187 B.n469 B.n132 585
R188 B.n468 B.n467 585
R189 B.n466 B.n133 585
R190 B.n465 B.n464 585
R191 B.n463 B.n134 585
R192 B.n462 B.n461 585
R193 B.n460 B.n135 585
R194 B.n459 B.n458 585
R195 B.n457 B.n136 585
R196 B.n456 B.n455 585
R197 B.n454 B.n137 585
R198 B.n453 B.n452 585
R199 B.n451 B.n138 585
R200 B.n450 B.n449 585
R201 B.n448 B.n139 585
R202 B.n447 B.n446 585
R203 B.n445 B.n140 585
R204 B.n444 B.n443 585
R205 B.n442 B.n141 585
R206 B.n441 B.n440 585
R207 B.n439 B.n142 585
R208 B.n438 B.n437 585
R209 B.n313 B.n188 585
R210 B.n315 B.n314 585
R211 B.n316 B.n187 585
R212 B.n318 B.n317 585
R213 B.n319 B.n186 585
R214 B.n321 B.n320 585
R215 B.n322 B.n185 585
R216 B.n324 B.n323 585
R217 B.n325 B.n184 585
R218 B.n327 B.n326 585
R219 B.n328 B.n183 585
R220 B.n330 B.n329 585
R221 B.n331 B.n182 585
R222 B.n333 B.n332 585
R223 B.n334 B.n181 585
R224 B.n336 B.n335 585
R225 B.n337 B.n180 585
R226 B.n339 B.n338 585
R227 B.n340 B.n179 585
R228 B.n342 B.n341 585
R229 B.n343 B.n178 585
R230 B.n345 B.n344 585
R231 B.n346 B.n177 585
R232 B.n348 B.n347 585
R233 B.n349 B.n176 585
R234 B.n351 B.n350 585
R235 B.n352 B.n175 585
R236 B.n354 B.n353 585
R237 B.n355 B.n174 585
R238 B.n357 B.n356 585
R239 B.n358 B.n173 585
R240 B.n360 B.n359 585
R241 B.n361 B.n172 585
R242 B.n363 B.n362 585
R243 B.n364 B.n171 585
R244 B.n366 B.n365 585
R245 B.n368 B.n168 585
R246 B.n370 B.n369 585
R247 B.n371 B.n167 585
R248 B.n373 B.n372 585
R249 B.n374 B.n166 585
R250 B.n376 B.n375 585
R251 B.n377 B.n165 585
R252 B.n379 B.n378 585
R253 B.n380 B.n164 585
R254 B.n382 B.n381 585
R255 B.n384 B.n383 585
R256 B.n385 B.n160 585
R257 B.n387 B.n386 585
R258 B.n388 B.n159 585
R259 B.n390 B.n389 585
R260 B.n391 B.n158 585
R261 B.n393 B.n392 585
R262 B.n394 B.n157 585
R263 B.n396 B.n395 585
R264 B.n397 B.n156 585
R265 B.n399 B.n398 585
R266 B.n400 B.n155 585
R267 B.n402 B.n401 585
R268 B.n403 B.n154 585
R269 B.n405 B.n404 585
R270 B.n406 B.n153 585
R271 B.n408 B.n407 585
R272 B.n409 B.n152 585
R273 B.n411 B.n410 585
R274 B.n412 B.n151 585
R275 B.n414 B.n413 585
R276 B.n415 B.n150 585
R277 B.n417 B.n416 585
R278 B.n418 B.n149 585
R279 B.n420 B.n419 585
R280 B.n421 B.n148 585
R281 B.n423 B.n422 585
R282 B.n424 B.n147 585
R283 B.n426 B.n425 585
R284 B.n427 B.n146 585
R285 B.n429 B.n428 585
R286 B.n430 B.n145 585
R287 B.n432 B.n431 585
R288 B.n433 B.n144 585
R289 B.n435 B.n434 585
R290 B.n436 B.n143 585
R291 B.n312 B.n311 585
R292 B.n310 B.n189 585
R293 B.n309 B.n308 585
R294 B.n307 B.n190 585
R295 B.n306 B.n305 585
R296 B.n304 B.n191 585
R297 B.n303 B.n302 585
R298 B.n301 B.n192 585
R299 B.n300 B.n299 585
R300 B.n298 B.n193 585
R301 B.n297 B.n296 585
R302 B.n295 B.n194 585
R303 B.n294 B.n293 585
R304 B.n292 B.n195 585
R305 B.n291 B.n290 585
R306 B.n289 B.n196 585
R307 B.n288 B.n287 585
R308 B.n286 B.n197 585
R309 B.n285 B.n284 585
R310 B.n283 B.n198 585
R311 B.n282 B.n281 585
R312 B.n280 B.n199 585
R313 B.n279 B.n278 585
R314 B.n277 B.n200 585
R315 B.n276 B.n275 585
R316 B.n274 B.n201 585
R317 B.n273 B.n272 585
R318 B.n271 B.n202 585
R319 B.n270 B.n269 585
R320 B.n268 B.n203 585
R321 B.n267 B.n266 585
R322 B.n265 B.n204 585
R323 B.n264 B.n263 585
R324 B.n262 B.n205 585
R325 B.n261 B.n260 585
R326 B.n259 B.n206 585
R327 B.n258 B.n257 585
R328 B.n256 B.n207 585
R329 B.n255 B.n254 585
R330 B.n253 B.n208 585
R331 B.n252 B.n251 585
R332 B.n250 B.n209 585
R333 B.n249 B.n248 585
R334 B.n247 B.n210 585
R335 B.n246 B.n245 585
R336 B.n244 B.n211 585
R337 B.n243 B.n242 585
R338 B.n241 B.n212 585
R339 B.n240 B.n239 585
R340 B.n238 B.n213 585
R341 B.n237 B.n236 585
R342 B.n235 B.n214 585
R343 B.n234 B.n233 585
R344 B.n232 B.n215 585
R345 B.n231 B.n230 585
R346 B.n229 B.n216 585
R347 B.n228 B.n227 585
R348 B.n226 B.n217 585
R349 B.n225 B.n224 585
R350 B.n223 B.n218 585
R351 B.n222 B.n221 585
R352 B.n220 B.n219 585
R353 B.n2 B.n0 585
R354 B.n845 B.n1 585
R355 B.n844 B.n843 585
R356 B.n842 B.n3 585
R357 B.n841 B.n840 585
R358 B.n839 B.n4 585
R359 B.n838 B.n837 585
R360 B.n836 B.n5 585
R361 B.n835 B.n834 585
R362 B.n833 B.n6 585
R363 B.n832 B.n831 585
R364 B.n830 B.n7 585
R365 B.n829 B.n828 585
R366 B.n827 B.n8 585
R367 B.n826 B.n825 585
R368 B.n824 B.n9 585
R369 B.n823 B.n822 585
R370 B.n821 B.n10 585
R371 B.n820 B.n819 585
R372 B.n818 B.n11 585
R373 B.n817 B.n816 585
R374 B.n815 B.n12 585
R375 B.n814 B.n813 585
R376 B.n812 B.n13 585
R377 B.n811 B.n810 585
R378 B.n809 B.n14 585
R379 B.n808 B.n807 585
R380 B.n806 B.n15 585
R381 B.n805 B.n804 585
R382 B.n803 B.n16 585
R383 B.n802 B.n801 585
R384 B.n800 B.n17 585
R385 B.n799 B.n798 585
R386 B.n797 B.n18 585
R387 B.n796 B.n795 585
R388 B.n794 B.n19 585
R389 B.n793 B.n792 585
R390 B.n791 B.n20 585
R391 B.n790 B.n789 585
R392 B.n788 B.n21 585
R393 B.n787 B.n786 585
R394 B.n785 B.n22 585
R395 B.n784 B.n783 585
R396 B.n782 B.n23 585
R397 B.n781 B.n780 585
R398 B.n779 B.n24 585
R399 B.n778 B.n777 585
R400 B.n776 B.n25 585
R401 B.n775 B.n774 585
R402 B.n773 B.n26 585
R403 B.n772 B.n771 585
R404 B.n770 B.n27 585
R405 B.n769 B.n768 585
R406 B.n767 B.n28 585
R407 B.n766 B.n765 585
R408 B.n764 B.n29 585
R409 B.n763 B.n762 585
R410 B.n761 B.n30 585
R411 B.n760 B.n759 585
R412 B.n758 B.n31 585
R413 B.n757 B.n756 585
R414 B.n755 B.n32 585
R415 B.n754 B.n753 585
R416 B.n752 B.n33 585
R417 B.n847 B.n846 585
R418 B.n311 B.n188 535.745
R419 B.n750 B.n33 535.745
R420 B.n437 B.n436 535.745
R421 B.n628 B.n627 535.745
R422 B.n161 B.t0 297.075
R423 B.n169 B.t9 297.075
R424 B.n52 B.t6 297.075
R425 B.n60 B.t3 297.075
R426 B.n161 B.t2 168.681
R427 B.n60 B.t4 168.681
R428 B.n169 B.t11 168.669
R429 B.n52 B.t7 168.669
R430 B.n311 B.n310 163.367
R431 B.n310 B.n309 163.367
R432 B.n309 B.n190 163.367
R433 B.n305 B.n190 163.367
R434 B.n305 B.n304 163.367
R435 B.n304 B.n303 163.367
R436 B.n303 B.n192 163.367
R437 B.n299 B.n192 163.367
R438 B.n299 B.n298 163.367
R439 B.n298 B.n297 163.367
R440 B.n297 B.n194 163.367
R441 B.n293 B.n194 163.367
R442 B.n293 B.n292 163.367
R443 B.n292 B.n291 163.367
R444 B.n291 B.n196 163.367
R445 B.n287 B.n196 163.367
R446 B.n287 B.n286 163.367
R447 B.n286 B.n285 163.367
R448 B.n285 B.n198 163.367
R449 B.n281 B.n198 163.367
R450 B.n281 B.n280 163.367
R451 B.n280 B.n279 163.367
R452 B.n279 B.n200 163.367
R453 B.n275 B.n200 163.367
R454 B.n275 B.n274 163.367
R455 B.n274 B.n273 163.367
R456 B.n273 B.n202 163.367
R457 B.n269 B.n202 163.367
R458 B.n269 B.n268 163.367
R459 B.n268 B.n267 163.367
R460 B.n267 B.n204 163.367
R461 B.n263 B.n204 163.367
R462 B.n263 B.n262 163.367
R463 B.n262 B.n261 163.367
R464 B.n261 B.n206 163.367
R465 B.n257 B.n206 163.367
R466 B.n257 B.n256 163.367
R467 B.n256 B.n255 163.367
R468 B.n255 B.n208 163.367
R469 B.n251 B.n208 163.367
R470 B.n251 B.n250 163.367
R471 B.n250 B.n249 163.367
R472 B.n249 B.n210 163.367
R473 B.n245 B.n210 163.367
R474 B.n245 B.n244 163.367
R475 B.n244 B.n243 163.367
R476 B.n243 B.n212 163.367
R477 B.n239 B.n212 163.367
R478 B.n239 B.n238 163.367
R479 B.n238 B.n237 163.367
R480 B.n237 B.n214 163.367
R481 B.n233 B.n214 163.367
R482 B.n233 B.n232 163.367
R483 B.n232 B.n231 163.367
R484 B.n231 B.n216 163.367
R485 B.n227 B.n216 163.367
R486 B.n227 B.n226 163.367
R487 B.n226 B.n225 163.367
R488 B.n225 B.n218 163.367
R489 B.n221 B.n218 163.367
R490 B.n221 B.n220 163.367
R491 B.n220 B.n2 163.367
R492 B.n846 B.n2 163.367
R493 B.n846 B.n845 163.367
R494 B.n845 B.n844 163.367
R495 B.n844 B.n3 163.367
R496 B.n840 B.n3 163.367
R497 B.n840 B.n839 163.367
R498 B.n839 B.n838 163.367
R499 B.n838 B.n5 163.367
R500 B.n834 B.n5 163.367
R501 B.n834 B.n833 163.367
R502 B.n833 B.n832 163.367
R503 B.n832 B.n7 163.367
R504 B.n828 B.n7 163.367
R505 B.n828 B.n827 163.367
R506 B.n827 B.n826 163.367
R507 B.n826 B.n9 163.367
R508 B.n822 B.n9 163.367
R509 B.n822 B.n821 163.367
R510 B.n821 B.n820 163.367
R511 B.n820 B.n11 163.367
R512 B.n816 B.n11 163.367
R513 B.n816 B.n815 163.367
R514 B.n815 B.n814 163.367
R515 B.n814 B.n13 163.367
R516 B.n810 B.n13 163.367
R517 B.n810 B.n809 163.367
R518 B.n809 B.n808 163.367
R519 B.n808 B.n15 163.367
R520 B.n804 B.n15 163.367
R521 B.n804 B.n803 163.367
R522 B.n803 B.n802 163.367
R523 B.n802 B.n17 163.367
R524 B.n798 B.n17 163.367
R525 B.n798 B.n797 163.367
R526 B.n797 B.n796 163.367
R527 B.n796 B.n19 163.367
R528 B.n792 B.n19 163.367
R529 B.n792 B.n791 163.367
R530 B.n791 B.n790 163.367
R531 B.n790 B.n21 163.367
R532 B.n786 B.n21 163.367
R533 B.n786 B.n785 163.367
R534 B.n785 B.n784 163.367
R535 B.n784 B.n23 163.367
R536 B.n780 B.n23 163.367
R537 B.n780 B.n779 163.367
R538 B.n779 B.n778 163.367
R539 B.n778 B.n25 163.367
R540 B.n774 B.n25 163.367
R541 B.n774 B.n773 163.367
R542 B.n773 B.n772 163.367
R543 B.n772 B.n27 163.367
R544 B.n768 B.n27 163.367
R545 B.n768 B.n767 163.367
R546 B.n767 B.n766 163.367
R547 B.n766 B.n29 163.367
R548 B.n762 B.n29 163.367
R549 B.n762 B.n761 163.367
R550 B.n761 B.n760 163.367
R551 B.n760 B.n31 163.367
R552 B.n756 B.n31 163.367
R553 B.n756 B.n755 163.367
R554 B.n755 B.n754 163.367
R555 B.n754 B.n33 163.367
R556 B.n315 B.n188 163.367
R557 B.n316 B.n315 163.367
R558 B.n317 B.n316 163.367
R559 B.n317 B.n186 163.367
R560 B.n321 B.n186 163.367
R561 B.n322 B.n321 163.367
R562 B.n323 B.n322 163.367
R563 B.n323 B.n184 163.367
R564 B.n327 B.n184 163.367
R565 B.n328 B.n327 163.367
R566 B.n329 B.n328 163.367
R567 B.n329 B.n182 163.367
R568 B.n333 B.n182 163.367
R569 B.n334 B.n333 163.367
R570 B.n335 B.n334 163.367
R571 B.n335 B.n180 163.367
R572 B.n339 B.n180 163.367
R573 B.n340 B.n339 163.367
R574 B.n341 B.n340 163.367
R575 B.n341 B.n178 163.367
R576 B.n345 B.n178 163.367
R577 B.n346 B.n345 163.367
R578 B.n347 B.n346 163.367
R579 B.n347 B.n176 163.367
R580 B.n351 B.n176 163.367
R581 B.n352 B.n351 163.367
R582 B.n353 B.n352 163.367
R583 B.n353 B.n174 163.367
R584 B.n357 B.n174 163.367
R585 B.n358 B.n357 163.367
R586 B.n359 B.n358 163.367
R587 B.n359 B.n172 163.367
R588 B.n363 B.n172 163.367
R589 B.n364 B.n363 163.367
R590 B.n365 B.n364 163.367
R591 B.n365 B.n168 163.367
R592 B.n370 B.n168 163.367
R593 B.n371 B.n370 163.367
R594 B.n372 B.n371 163.367
R595 B.n372 B.n166 163.367
R596 B.n376 B.n166 163.367
R597 B.n377 B.n376 163.367
R598 B.n378 B.n377 163.367
R599 B.n378 B.n164 163.367
R600 B.n382 B.n164 163.367
R601 B.n383 B.n382 163.367
R602 B.n383 B.n160 163.367
R603 B.n387 B.n160 163.367
R604 B.n388 B.n387 163.367
R605 B.n389 B.n388 163.367
R606 B.n389 B.n158 163.367
R607 B.n393 B.n158 163.367
R608 B.n394 B.n393 163.367
R609 B.n395 B.n394 163.367
R610 B.n395 B.n156 163.367
R611 B.n399 B.n156 163.367
R612 B.n400 B.n399 163.367
R613 B.n401 B.n400 163.367
R614 B.n401 B.n154 163.367
R615 B.n405 B.n154 163.367
R616 B.n406 B.n405 163.367
R617 B.n407 B.n406 163.367
R618 B.n407 B.n152 163.367
R619 B.n411 B.n152 163.367
R620 B.n412 B.n411 163.367
R621 B.n413 B.n412 163.367
R622 B.n413 B.n150 163.367
R623 B.n417 B.n150 163.367
R624 B.n418 B.n417 163.367
R625 B.n419 B.n418 163.367
R626 B.n419 B.n148 163.367
R627 B.n423 B.n148 163.367
R628 B.n424 B.n423 163.367
R629 B.n425 B.n424 163.367
R630 B.n425 B.n146 163.367
R631 B.n429 B.n146 163.367
R632 B.n430 B.n429 163.367
R633 B.n431 B.n430 163.367
R634 B.n431 B.n144 163.367
R635 B.n435 B.n144 163.367
R636 B.n436 B.n435 163.367
R637 B.n437 B.n142 163.367
R638 B.n441 B.n142 163.367
R639 B.n442 B.n441 163.367
R640 B.n443 B.n442 163.367
R641 B.n443 B.n140 163.367
R642 B.n447 B.n140 163.367
R643 B.n448 B.n447 163.367
R644 B.n449 B.n448 163.367
R645 B.n449 B.n138 163.367
R646 B.n453 B.n138 163.367
R647 B.n454 B.n453 163.367
R648 B.n455 B.n454 163.367
R649 B.n455 B.n136 163.367
R650 B.n459 B.n136 163.367
R651 B.n460 B.n459 163.367
R652 B.n461 B.n460 163.367
R653 B.n461 B.n134 163.367
R654 B.n465 B.n134 163.367
R655 B.n466 B.n465 163.367
R656 B.n467 B.n466 163.367
R657 B.n467 B.n132 163.367
R658 B.n471 B.n132 163.367
R659 B.n472 B.n471 163.367
R660 B.n473 B.n472 163.367
R661 B.n473 B.n130 163.367
R662 B.n477 B.n130 163.367
R663 B.n478 B.n477 163.367
R664 B.n479 B.n478 163.367
R665 B.n479 B.n128 163.367
R666 B.n483 B.n128 163.367
R667 B.n484 B.n483 163.367
R668 B.n485 B.n484 163.367
R669 B.n485 B.n126 163.367
R670 B.n489 B.n126 163.367
R671 B.n490 B.n489 163.367
R672 B.n491 B.n490 163.367
R673 B.n491 B.n124 163.367
R674 B.n495 B.n124 163.367
R675 B.n496 B.n495 163.367
R676 B.n497 B.n496 163.367
R677 B.n497 B.n122 163.367
R678 B.n501 B.n122 163.367
R679 B.n502 B.n501 163.367
R680 B.n503 B.n502 163.367
R681 B.n503 B.n120 163.367
R682 B.n507 B.n120 163.367
R683 B.n508 B.n507 163.367
R684 B.n509 B.n508 163.367
R685 B.n509 B.n118 163.367
R686 B.n513 B.n118 163.367
R687 B.n514 B.n513 163.367
R688 B.n515 B.n514 163.367
R689 B.n515 B.n116 163.367
R690 B.n519 B.n116 163.367
R691 B.n520 B.n519 163.367
R692 B.n521 B.n520 163.367
R693 B.n521 B.n114 163.367
R694 B.n525 B.n114 163.367
R695 B.n526 B.n525 163.367
R696 B.n527 B.n526 163.367
R697 B.n527 B.n112 163.367
R698 B.n531 B.n112 163.367
R699 B.n532 B.n531 163.367
R700 B.n533 B.n532 163.367
R701 B.n533 B.n110 163.367
R702 B.n537 B.n110 163.367
R703 B.n538 B.n537 163.367
R704 B.n539 B.n538 163.367
R705 B.n539 B.n108 163.367
R706 B.n543 B.n108 163.367
R707 B.n544 B.n543 163.367
R708 B.n545 B.n544 163.367
R709 B.n545 B.n106 163.367
R710 B.n549 B.n106 163.367
R711 B.n550 B.n549 163.367
R712 B.n551 B.n550 163.367
R713 B.n551 B.n104 163.367
R714 B.n555 B.n104 163.367
R715 B.n556 B.n555 163.367
R716 B.n557 B.n556 163.367
R717 B.n557 B.n102 163.367
R718 B.n561 B.n102 163.367
R719 B.n562 B.n561 163.367
R720 B.n563 B.n562 163.367
R721 B.n563 B.n100 163.367
R722 B.n567 B.n100 163.367
R723 B.n568 B.n567 163.367
R724 B.n569 B.n568 163.367
R725 B.n569 B.n98 163.367
R726 B.n573 B.n98 163.367
R727 B.n574 B.n573 163.367
R728 B.n575 B.n574 163.367
R729 B.n575 B.n96 163.367
R730 B.n579 B.n96 163.367
R731 B.n580 B.n579 163.367
R732 B.n581 B.n580 163.367
R733 B.n581 B.n94 163.367
R734 B.n585 B.n94 163.367
R735 B.n586 B.n585 163.367
R736 B.n587 B.n586 163.367
R737 B.n587 B.n92 163.367
R738 B.n591 B.n92 163.367
R739 B.n592 B.n591 163.367
R740 B.n593 B.n592 163.367
R741 B.n593 B.n90 163.367
R742 B.n597 B.n90 163.367
R743 B.n598 B.n597 163.367
R744 B.n599 B.n598 163.367
R745 B.n599 B.n88 163.367
R746 B.n603 B.n88 163.367
R747 B.n604 B.n603 163.367
R748 B.n605 B.n604 163.367
R749 B.n605 B.n86 163.367
R750 B.n609 B.n86 163.367
R751 B.n610 B.n609 163.367
R752 B.n611 B.n610 163.367
R753 B.n611 B.n84 163.367
R754 B.n615 B.n84 163.367
R755 B.n616 B.n615 163.367
R756 B.n617 B.n616 163.367
R757 B.n617 B.n82 163.367
R758 B.n621 B.n82 163.367
R759 B.n622 B.n621 163.367
R760 B.n623 B.n622 163.367
R761 B.n623 B.n80 163.367
R762 B.n627 B.n80 163.367
R763 B.n750 B.n749 163.367
R764 B.n749 B.n748 163.367
R765 B.n748 B.n35 163.367
R766 B.n744 B.n35 163.367
R767 B.n744 B.n743 163.367
R768 B.n743 B.n742 163.367
R769 B.n742 B.n37 163.367
R770 B.n738 B.n37 163.367
R771 B.n738 B.n737 163.367
R772 B.n737 B.n736 163.367
R773 B.n736 B.n39 163.367
R774 B.n732 B.n39 163.367
R775 B.n732 B.n731 163.367
R776 B.n731 B.n730 163.367
R777 B.n730 B.n41 163.367
R778 B.n726 B.n41 163.367
R779 B.n726 B.n725 163.367
R780 B.n725 B.n724 163.367
R781 B.n724 B.n43 163.367
R782 B.n720 B.n43 163.367
R783 B.n720 B.n719 163.367
R784 B.n719 B.n718 163.367
R785 B.n718 B.n45 163.367
R786 B.n714 B.n45 163.367
R787 B.n714 B.n713 163.367
R788 B.n713 B.n712 163.367
R789 B.n712 B.n47 163.367
R790 B.n708 B.n47 163.367
R791 B.n708 B.n707 163.367
R792 B.n707 B.n706 163.367
R793 B.n706 B.n49 163.367
R794 B.n702 B.n49 163.367
R795 B.n702 B.n701 163.367
R796 B.n701 B.n700 163.367
R797 B.n700 B.n51 163.367
R798 B.n695 B.n51 163.367
R799 B.n695 B.n694 163.367
R800 B.n694 B.n693 163.367
R801 B.n693 B.n55 163.367
R802 B.n689 B.n55 163.367
R803 B.n689 B.n688 163.367
R804 B.n688 B.n687 163.367
R805 B.n687 B.n57 163.367
R806 B.n683 B.n57 163.367
R807 B.n683 B.n682 163.367
R808 B.n682 B.n681 163.367
R809 B.n681 B.n59 163.367
R810 B.n677 B.n59 163.367
R811 B.n677 B.n676 163.367
R812 B.n676 B.n675 163.367
R813 B.n675 B.n64 163.367
R814 B.n671 B.n64 163.367
R815 B.n671 B.n670 163.367
R816 B.n670 B.n669 163.367
R817 B.n669 B.n66 163.367
R818 B.n665 B.n66 163.367
R819 B.n665 B.n664 163.367
R820 B.n664 B.n663 163.367
R821 B.n663 B.n68 163.367
R822 B.n659 B.n68 163.367
R823 B.n659 B.n658 163.367
R824 B.n658 B.n657 163.367
R825 B.n657 B.n70 163.367
R826 B.n653 B.n70 163.367
R827 B.n653 B.n652 163.367
R828 B.n652 B.n651 163.367
R829 B.n651 B.n72 163.367
R830 B.n647 B.n72 163.367
R831 B.n647 B.n646 163.367
R832 B.n646 B.n645 163.367
R833 B.n645 B.n74 163.367
R834 B.n641 B.n74 163.367
R835 B.n641 B.n640 163.367
R836 B.n640 B.n639 163.367
R837 B.n639 B.n76 163.367
R838 B.n635 B.n76 163.367
R839 B.n635 B.n634 163.367
R840 B.n634 B.n633 163.367
R841 B.n633 B.n78 163.367
R842 B.n629 B.n78 163.367
R843 B.n629 B.n628 163.367
R844 B.n162 B.t1 108.367
R845 B.n61 B.t5 108.367
R846 B.n170 B.t10 108.355
R847 B.n53 B.t8 108.355
R848 B.n162 B.n161 60.3157
R849 B.n170 B.n169 60.3157
R850 B.n53 B.n52 60.3157
R851 B.n61 B.n60 60.3157
R852 B.n163 B.n162 59.5399
R853 B.n367 B.n170 59.5399
R854 B.n697 B.n53 59.5399
R855 B.n62 B.n61 59.5399
R856 B.n752 B.n751 34.8103
R857 B.n626 B.n79 34.8103
R858 B.n438 B.n143 34.8103
R859 B.n313 B.n312 34.8103
R860 B B.n847 18.0485
R861 B.n751 B.n34 10.6151
R862 B.n747 B.n34 10.6151
R863 B.n747 B.n746 10.6151
R864 B.n746 B.n745 10.6151
R865 B.n745 B.n36 10.6151
R866 B.n741 B.n36 10.6151
R867 B.n741 B.n740 10.6151
R868 B.n740 B.n739 10.6151
R869 B.n739 B.n38 10.6151
R870 B.n735 B.n38 10.6151
R871 B.n735 B.n734 10.6151
R872 B.n734 B.n733 10.6151
R873 B.n733 B.n40 10.6151
R874 B.n729 B.n40 10.6151
R875 B.n729 B.n728 10.6151
R876 B.n728 B.n727 10.6151
R877 B.n727 B.n42 10.6151
R878 B.n723 B.n42 10.6151
R879 B.n723 B.n722 10.6151
R880 B.n722 B.n721 10.6151
R881 B.n721 B.n44 10.6151
R882 B.n717 B.n44 10.6151
R883 B.n717 B.n716 10.6151
R884 B.n716 B.n715 10.6151
R885 B.n715 B.n46 10.6151
R886 B.n711 B.n46 10.6151
R887 B.n711 B.n710 10.6151
R888 B.n710 B.n709 10.6151
R889 B.n709 B.n48 10.6151
R890 B.n705 B.n48 10.6151
R891 B.n705 B.n704 10.6151
R892 B.n704 B.n703 10.6151
R893 B.n703 B.n50 10.6151
R894 B.n699 B.n50 10.6151
R895 B.n699 B.n698 10.6151
R896 B.n696 B.n54 10.6151
R897 B.n692 B.n54 10.6151
R898 B.n692 B.n691 10.6151
R899 B.n691 B.n690 10.6151
R900 B.n690 B.n56 10.6151
R901 B.n686 B.n56 10.6151
R902 B.n686 B.n685 10.6151
R903 B.n685 B.n684 10.6151
R904 B.n684 B.n58 10.6151
R905 B.n680 B.n679 10.6151
R906 B.n679 B.n678 10.6151
R907 B.n678 B.n63 10.6151
R908 B.n674 B.n63 10.6151
R909 B.n674 B.n673 10.6151
R910 B.n673 B.n672 10.6151
R911 B.n672 B.n65 10.6151
R912 B.n668 B.n65 10.6151
R913 B.n668 B.n667 10.6151
R914 B.n667 B.n666 10.6151
R915 B.n666 B.n67 10.6151
R916 B.n662 B.n67 10.6151
R917 B.n662 B.n661 10.6151
R918 B.n661 B.n660 10.6151
R919 B.n660 B.n69 10.6151
R920 B.n656 B.n69 10.6151
R921 B.n656 B.n655 10.6151
R922 B.n655 B.n654 10.6151
R923 B.n654 B.n71 10.6151
R924 B.n650 B.n71 10.6151
R925 B.n650 B.n649 10.6151
R926 B.n649 B.n648 10.6151
R927 B.n648 B.n73 10.6151
R928 B.n644 B.n73 10.6151
R929 B.n644 B.n643 10.6151
R930 B.n643 B.n642 10.6151
R931 B.n642 B.n75 10.6151
R932 B.n638 B.n75 10.6151
R933 B.n638 B.n637 10.6151
R934 B.n637 B.n636 10.6151
R935 B.n636 B.n77 10.6151
R936 B.n632 B.n77 10.6151
R937 B.n632 B.n631 10.6151
R938 B.n631 B.n630 10.6151
R939 B.n630 B.n79 10.6151
R940 B.n439 B.n438 10.6151
R941 B.n440 B.n439 10.6151
R942 B.n440 B.n141 10.6151
R943 B.n444 B.n141 10.6151
R944 B.n445 B.n444 10.6151
R945 B.n446 B.n445 10.6151
R946 B.n446 B.n139 10.6151
R947 B.n450 B.n139 10.6151
R948 B.n451 B.n450 10.6151
R949 B.n452 B.n451 10.6151
R950 B.n452 B.n137 10.6151
R951 B.n456 B.n137 10.6151
R952 B.n457 B.n456 10.6151
R953 B.n458 B.n457 10.6151
R954 B.n458 B.n135 10.6151
R955 B.n462 B.n135 10.6151
R956 B.n463 B.n462 10.6151
R957 B.n464 B.n463 10.6151
R958 B.n464 B.n133 10.6151
R959 B.n468 B.n133 10.6151
R960 B.n469 B.n468 10.6151
R961 B.n470 B.n469 10.6151
R962 B.n470 B.n131 10.6151
R963 B.n474 B.n131 10.6151
R964 B.n475 B.n474 10.6151
R965 B.n476 B.n475 10.6151
R966 B.n476 B.n129 10.6151
R967 B.n480 B.n129 10.6151
R968 B.n481 B.n480 10.6151
R969 B.n482 B.n481 10.6151
R970 B.n482 B.n127 10.6151
R971 B.n486 B.n127 10.6151
R972 B.n487 B.n486 10.6151
R973 B.n488 B.n487 10.6151
R974 B.n488 B.n125 10.6151
R975 B.n492 B.n125 10.6151
R976 B.n493 B.n492 10.6151
R977 B.n494 B.n493 10.6151
R978 B.n494 B.n123 10.6151
R979 B.n498 B.n123 10.6151
R980 B.n499 B.n498 10.6151
R981 B.n500 B.n499 10.6151
R982 B.n500 B.n121 10.6151
R983 B.n504 B.n121 10.6151
R984 B.n505 B.n504 10.6151
R985 B.n506 B.n505 10.6151
R986 B.n506 B.n119 10.6151
R987 B.n510 B.n119 10.6151
R988 B.n511 B.n510 10.6151
R989 B.n512 B.n511 10.6151
R990 B.n512 B.n117 10.6151
R991 B.n516 B.n117 10.6151
R992 B.n517 B.n516 10.6151
R993 B.n518 B.n517 10.6151
R994 B.n518 B.n115 10.6151
R995 B.n522 B.n115 10.6151
R996 B.n523 B.n522 10.6151
R997 B.n524 B.n523 10.6151
R998 B.n524 B.n113 10.6151
R999 B.n528 B.n113 10.6151
R1000 B.n529 B.n528 10.6151
R1001 B.n530 B.n529 10.6151
R1002 B.n530 B.n111 10.6151
R1003 B.n534 B.n111 10.6151
R1004 B.n535 B.n534 10.6151
R1005 B.n536 B.n535 10.6151
R1006 B.n536 B.n109 10.6151
R1007 B.n540 B.n109 10.6151
R1008 B.n541 B.n540 10.6151
R1009 B.n542 B.n541 10.6151
R1010 B.n542 B.n107 10.6151
R1011 B.n546 B.n107 10.6151
R1012 B.n547 B.n546 10.6151
R1013 B.n548 B.n547 10.6151
R1014 B.n548 B.n105 10.6151
R1015 B.n552 B.n105 10.6151
R1016 B.n553 B.n552 10.6151
R1017 B.n554 B.n553 10.6151
R1018 B.n554 B.n103 10.6151
R1019 B.n558 B.n103 10.6151
R1020 B.n559 B.n558 10.6151
R1021 B.n560 B.n559 10.6151
R1022 B.n560 B.n101 10.6151
R1023 B.n564 B.n101 10.6151
R1024 B.n565 B.n564 10.6151
R1025 B.n566 B.n565 10.6151
R1026 B.n566 B.n99 10.6151
R1027 B.n570 B.n99 10.6151
R1028 B.n571 B.n570 10.6151
R1029 B.n572 B.n571 10.6151
R1030 B.n572 B.n97 10.6151
R1031 B.n576 B.n97 10.6151
R1032 B.n577 B.n576 10.6151
R1033 B.n578 B.n577 10.6151
R1034 B.n578 B.n95 10.6151
R1035 B.n582 B.n95 10.6151
R1036 B.n583 B.n582 10.6151
R1037 B.n584 B.n583 10.6151
R1038 B.n584 B.n93 10.6151
R1039 B.n588 B.n93 10.6151
R1040 B.n589 B.n588 10.6151
R1041 B.n590 B.n589 10.6151
R1042 B.n590 B.n91 10.6151
R1043 B.n594 B.n91 10.6151
R1044 B.n595 B.n594 10.6151
R1045 B.n596 B.n595 10.6151
R1046 B.n596 B.n89 10.6151
R1047 B.n600 B.n89 10.6151
R1048 B.n601 B.n600 10.6151
R1049 B.n602 B.n601 10.6151
R1050 B.n602 B.n87 10.6151
R1051 B.n606 B.n87 10.6151
R1052 B.n607 B.n606 10.6151
R1053 B.n608 B.n607 10.6151
R1054 B.n608 B.n85 10.6151
R1055 B.n612 B.n85 10.6151
R1056 B.n613 B.n612 10.6151
R1057 B.n614 B.n613 10.6151
R1058 B.n614 B.n83 10.6151
R1059 B.n618 B.n83 10.6151
R1060 B.n619 B.n618 10.6151
R1061 B.n620 B.n619 10.6151
R1062 B.n620 B.n81 10.6151
R1063 B.n624 B.n81 10.6151
R1064 B.n625 B.n624 10.6151
R1065 B.n626 B.n625 10.6151
R1066 B.n314 B.n313 10.6151
R1067 B.n314 B.n187 10.6151
R1068 B.n318 B.n187 10.6151
R1069 B.n319 B.n318 10.6151
R1070 B.n320 B.n319 10.6151
R1071 B.n320 B.n185 10.6151
R1072 B.n324 B.n185 10.6151
R1073 B.n325 B.n324 10.6151
R1074 B.n326 B.n325 10.6151
R1075 B.n326 B.n183 10.6151
R1076 B.n330 B.n183 10.6151
R1077 B.n331 B.n330 10.6151
R1078 B.n332 B.n331 10.6151
R1079 B.n332 B.n181 10.6151
R1080 B.n336 B.n181 10.6151
R1081 B.n337 B.n336 10.6151
R1082 B.n338 B.n337 10.6151
R1083 B.n338 B.n179 10.6151
R1084 B.n342 B.n179 10.6151
R1085 B.n343 B.n342 10.6151
R1086 B.n344 B.n343 10.6151
R1087 B.n344 B.n177 10.6151
R1088 B.n348 B.n177 10.6151
R1089 B.n349 B.n348 10.6151
R1090 B.n350 B.n349 10.6151
R1091 B.n350 B.n175 10.6151
R1092 B.n354 B.n175 10.6151
R1093 B.n355 B.n354 10.6151
R1094 B.n356 B.n355 10.6151
R1095 B.n356 B.n173 10.6151
R1096 B.n360 B.n173 10.6151
R1097 B.n361 B.n360 10.6151
R1098 B.n362 B.n361 10.6151
R1099 B.n362 B.n171 10.6151
R1100 B.n366 B.n171 10.6151
R1101 B.n369 B.n368 10.6151
R1102 B.n369 B.n167 10.6151
R1103 B.n373 B.n167 10.6151
R1104 B.n374 B.n373 10.6151
R1105 B.n375 B.n374 10.6151
R1106 B.n375 B.n165 10.6151
R1107 B.n379 B.n165 10.6151
R1108 B.n380 B.n379 10.6151
R1109 B.n381 B.n380 10.6151
R1110 B.n385 B.n384 10.6151
R1111 B.n386 B.n385 10.6151
R1112 B.n386 B.n159 10.6151
R1113 B.n390 B.n159 10.6151
R1114 B.n391 B.n390 10.6151
R1115 B.n392 B.n391 10.6151
R1116 B.n392 B.n157 10.6151
R1117 B.n396 B.n157 10.6151
R1118 B.n397 B.n396 10.6151
R1119 B.n398 B.n397 10.6151
R1120 B.n398 B.n155 10.6151
R1121 B.n402 B.n155 10.6151
R1122 B.n403 B.n402 10.6151
R1123 B.n404 B.n403 10.6151
R1124 B.n404 B.n153 10.6151
R1125 B.n408 B.n153 10.6151
R1126 B.n409 B.n408 10.6151
R1127 B.n410 B.n409 10.6151
R1128 B.n410 B.n151 10.6151
R1129 B.n414 B.n151 10.6151
R1130 B.n415 B.n414 10.6151
R1131 B.n416 B.n415 10.6151
R1132 B.n416 B.n149 10.6151
R1133 B.n420 B.n149 10.6151
R1134 B.n421 B.n420 10.6151
R1135 B.n422 B.n421 10.6151
R1136 B.n422 B.n147 10.6151
R1137 B.n426 B.n147 10.6151
R1138 B.n427 B.n426 10.6151
R1139 B.n428 B.n427 10.6151
R1140 B.n428 B.n145 10.6151
R1141 B.n432 B.n145 10.6151
R1142 B.n433 B.n432 10.6151
R1143 B.n434 B.n433 10.6151
R1144 B.n434 B.n143 10.6151
R1145 B.n312 B.n189 10.6151
R1146 B.n308 B.n189 10.6151
R1147 B.n308 B.n307 10.6151
R1148 B.n307 B.n306 10.6151
R1149 B.n306 B.n191 10.6151
R1150 B.n302 B.n191 10.6151
R1151 B.n302 B.n301 10.6151
R1152 B.n301 B.n300 10.6151
R1153 B.n300 B.n193 10.6151
R1154 B.n296 B.n193 10.6151
R1155 B.n296 B.n295 10.6151
R1156 B.n295 B.n294 10.6151
R1157 B.n294 B.n195 10.6151
R1158 B.n290 B.n195 10.6151
R1159 B.n290 B.n289 10.6151
R1160 B.n289 B.n288 10.6151
R1161 B.n288 B.n197 10.6151
R1162 B.n284 B.n197 10.6151
R1163 B.n284 B.n283 10.6151
R1164 B.n283 B.n282 10.6151
R1165 B.n282 B.n199 10.6151
R1166 B.n278 B.n199 10.6151
R1167 B.n278 B.n277 10.6151
R1168 B.n277 B.n276 10.6151
R1169 B.n276 B.n201 10.6151
R1170 B.n272 B.n201 10.6151
R1171 B.n272 B.n271 10.6151
R1172 B.n271 B.n270 10.6151
R1173 B.n270 B.n203 10.6151
R1174 B.n266 B.n203 10.6151
R1175 B.n266 B.n265 10.6151
R1176 B.n265 B.n264 10.6151
R1177 B.n264 B.n205 10.6151
R1178 B.n260 B.n205 10.6151
R1179 B.n260 B.n259 10.6151
R1180 B.n259 B.n258 10.6151
R1181 B.n258 B.n207 10.6151
R1182 B.n254 B.n207 10.6151
R1183 B.n254 B.n253 10.6151
R1184 B.n253 B.n252 10.6151
R1185 B.n252 B.n209 10.6151
R1186 B.n248 B.n209 10.6151
R1187 B.n248 B.n247 10.6151
R1188 B.n247 B.n246 10.6151
R1189 B.n246 B.n211 10.6151
R1190 B.n242 B.n211 10.6151
R1191 B.n242 B.n241 10.6151
R1192 B.n241 B.n240 10.6151
R1193 B.n240 B.n213 10.6151
R1194 B.n236 B.n213 10.6151
R1195 B.n236 B.n235 10.6151
R1196 B.n235 B.n234 10.6151
R1197 B.n234 B.n215 10.6151
R1198 B.n230 B.n215 10.6151
R1199 B.n230 B.n229 10.6151
R1200 B.n229 B.n228 10.6151
R1201 B.n228 B.n217 10.6151
R1202 B.n224 B.n217 10.6151
R1203 B.n224 B.n223 10.6151
R1204 B.n223 B.n222 10.6151
R1205 B.n222 B.n219 10.6151
R1206 B.n219 B.n0 10.6151
R1207 B.n843 B.n1 10.6151
R1208 B.n843 B.n842 10.6151
R1209 B.n842 B.n841 10.6151
R1210 B.n841 B.n4 10.6151
R1211 B.n837 B.n4 10.6151
R1212 B.n837 B.n836 10.6151
R1213 B.n836 B.n835 10.6151
R1214 B.n835 B.n6 10.6151
R1215 B.n831 B.n6 10.6151
R1216 B.n831 B.n830 10.6151
R1217 B.n830 B.n829 10.6151
R1218 B.n829 B.n8 10.6151
R1219 B.n825 B.n8 10.6151
R1220 B.n825 B.n824 10.6151
R1221 B.n824 B.n823 10.6151
R1222 B.n823 B.n10 10.6151
R1223 B.n819 B.n10 10.6151
R1224 B.n819 B.n818 10.6151
R1225 B.n818 B.n817 10.6151
R1226 B.n817 B.n12 10.6151
R1227 B.n813 B.n12 10.6151
R1228 B.n813 B.n812 10.6151
R1229 B.n812 B.n811 10.6151
R1230 B.n811 B.n14 10.6151
R1231 B.n807 B.n14 10.6151
R1232 B.n807 B.n806 10.6151
R1233 B.n806 B.n805 10.6151
R1234 B.n805 B.n16 10.6151
R1235 B.n801 B.n16 10.6151
R1236 B.n801 B.n800 10.6151
R1237 B.n800 B.n799 10.6151
R1238 B.n799 B.n18 10.6151
R1239 B.n795 B.n18 10.6151
R1240 B.n795 B.n794 10.6151
R1241 B.n794 B.n793 10.6151
R1242 B.n793 B.n20 10.6151
R1243 B.n789 B.n20 10.6151
R1244 B.n789 B.n788 10.6151
R1245 B.n788 B.n787 10.6151
R1246 B.n787 B.n22 10.6151
R1247 B.n783 B.n22 10.6151
R1248 B.n783 B.n782 10.6151
R1249 B.n782 B.n781 10.6151
R1250 B.n781 B.n24 10.6151
R1251 B.n777 B.n24 10.6151
R1252 B.n777 B.n776 10.6151
R1253 B.n776 B.n775 10.6151
R1254 B.n775 B.n26 10.6151
R1255 B.n771 B.n26 10.6151
R1256 B.n771 B.n770 10.6151
R1257 B.n770 B.n769 10.6151
R1258 B.n769 B.n28 10.6151
R1259 B.n765 B.n28 10.6151
R1260 B.n765 B.n764 10.6151
R1261 B.n764 B.n763 10.6151
R1262 B.n763 B.n30 10.6151
R1263 B.n759 B.n30 10.6151
R1264 B.n759 B.n758 10.6151
R1265 B.n758 B.n757 10.6151
R1266 B.n757 B.n32 10.6151
R1267 B.n753 B.n32 10.6151
R1268 B.n753 B.n752 10.6151
R1269 B.n698 B.n697 9.36635
R1270 B.n680 B.n62 9.36635
R1271 B.n367 B.n366 9.36635
R1272 B.n384 B.n163 9.36635
R1273 B.n847 B.n0 2.81026
R1274 B.n847 B.n1 2.81026
R1275 B.n697 B.n696 1.24928
R1276 B.n62 B.n58 1.24928
R1277 B.n368 B.n367 1.24928
R1278 B.n381 B.n163 1.24928
R1279 VP.n25 VP.n22 161.3
R1280 VP.n27 VP.n26 161.3
R1281 VP.n28 VP.n21 161.3
R1282 VP.n30 VP.n29 161.3
R1283 VP.n31 VP.n20 161.3
R1284 VP.n34 VP.n33 161.3
R1285 VP.n35 VP.n19 161.3
R1286 VP.n37 VP.n36 161.3
R1287 VP.n38 VP.n18 161.3
R1288 VP.n40 VP.n39 161.3
R1289 VP.n41 VP.n17 161.3
R1290 VP.n43 VP.n42 161.3
R1291 VP.n45 VP.n16 161.3
R1292 VP.n47 VP.n46 161.3
R1293 VP.n48 VP.n15 161.3
R1294 VP.n50 VP.n49 161.3
R1295 VP.n51 VP.n14 161.3
R1296 VP.n53 VP.n52 161.3
R1297 VP.n95 VP.n94 161.3
R1298 VP.n93 VP.n1 161.3
R1299 VP.n92 VP.n91 161.3
R1300 VP.n90 VP.n2 161.3
R1301 VP.n89 VP.n88 161.3
R1302 VP.n87 VP.n3 161.3
R1303 VP.n85 VP.n84 161.3
R1304 VP.n83 VP.n4 161.3
R1305 VP.n82 VP.n81 161.3
R1306 VP.n80 VP.n5 161.3
R1307 VP.n79 VP.n78 161.3
R1308 VP.n77 VP.n6 161.3
R1309 VP.n76 VP.n75 161.3
R1310 VP.n73 VP.n7 161.3
R1311 VP.n72 VP.n71 161.3
R1312 VP.n70 VP.n8 161.3
R1313 VP.n69 VP.n68 161.3
R1314 VP.n67 VP.n9 161.3
R1315 VP.n65 VP.n64 161.3
R1316 VP.n63 VP.n10 161.3
R1317 VP.n62 VP.n61 161.3
R1318 VP.n60 VP.n11 161.3
R1319 VP.n59 VP.n58 161.3
R1320 VP.n57 VP.n12 161.3
R1321 VP.n23 VP.t3 120.678
R1322 VP.n55 VP.t6 88.7717
R1323 VP.n66 VP.t4 88.7717
R1324 VP.n74 VP.t0 88.7717
R1325 VP.n86 VP.t7 88.7717
R1326 VP.n0 VP.t2 88.7717
R1327 VP.n13 VP.t1 88.7717
R1328 VP.n44 VP.t5 88.7717
R1329 VP.n32 VP.t8 88.7717
R1330 VP.n24 VP.t9 88.7717
R1331 VP.n56 VP.n55 67.0082
R1332 VP.n96 VP.n0 67.0082
R1333 VP.n54 VP.n13 67.0082
R1334 VP.n72 VP.n8 56.4773
R1335 VP.n81 VP.n80 56.4773
R1336 VP.n39 VP.n38 56.4773
R1337 VP.n30 VP.n21 56.4773
R1338 VP.n24 VP.n23 55.8592
R1339 VP.n56 VP.n54 52.8741
R1340 VP.n61 VP.n60 48.6874
R1341 VP.n92 VP.n2 48.6874
R1342 VP.n50 VP.n15 48.6874
R1343 VP.n60 VP.n59 32.1338
R1344 VP.n93 VP.n92 32.1338
R1345 VP.n51 VP.n50 32.1338
R1346 VP.n59 VP.n12 24.3439
R1347 VP.n61 VP.n10 24.3439
R1348 VP.n65 VP.n10 24.3439
R1349 VP.n68 VP.n67 24.3439
R1350 VP.n68 VP.n8 24.3439
R1351 VP.n73 VP.n72 24.3439
R1352 VP.n75 VP.n73 24.3439
R1353 VP.n79 VP.n6 24.3439
R1354 VP.n80 VP.n79 24.3439
R1355 VP.n81 VP.n4 24.3439
R1356 VP.n85 VP.n4 24.3439
R1357 VP.n88 VP.n87 24.3439
R1358 VP.n88 VP.n2 24.3439
R1359 VP.n94 VP.n93 24.3439
R1360 VP.n52 VP.n51 24.3439
R1361 VP.n39 VP.n17 24.3439
R1362 VP.n43 VP.n17 24.3439
R1363 VP.n46 VP.n45 24.3439
R1364 VP.n46 VP.n15 24.3439
R1365 VP.n31 VP.n30 24.3439
R1366 VP.n33 VP.n31 24.3439
R1367 VP.n37 VP.n19 24.3439
R1368 VP.n38 VP.n37 24.3439
R1369 VP.n26 VP.n25 24.3439
R1370 VP.n26 VP.n21 24.3439
R1371 VP.n55 VP.n12 22.8833
R1372 VP.n94 VP.n0 22.8833
R1373 VP.n52 VP.n13 22.8833
R1374 VP.n67 VP.n66 17.5278
R1375 VP.n86 VP.n85 17.5278
R1376 VP.n44 VP.n43 17.5278
R1377 VP.n25 VP.n24 17.5278
R1378 VP.n75 VP.n74 12.1722
R1379 VP.n74 VP.n6 12.1722
R1380 VP.n33 VP.n32 12.1722
R1381 VP.n32 VP.n19 12.1722
R1382 VP.n66 VP.n65 6.81666
R1383 VP.n87 VP.n86 6.81666
R1384 VP.n45 VP.n44 6.81666
R1385 VP.n23 VP.n22 5.32595
R1386 VP.n54 VP.n53 0.355081
R1387 VP.n57 VP.n56 0.355081
R1388 VP.n96 VP.n95 0.355081
R1389 VP VP.n96 0.26685
R1390 VP.n27 VP.n22 0.189894
R1391 VP.n28 VP.n27 0.189894
R1392 VP.n29 VP.n28 0.189894
R1393 VP.n29 VP.n20 0.189894
R1394 VP.n34 VP.n20 0.189894
R1395 VP.n35 VP.n34 0.189894
R1396 VP.n36 VP.n35 0.189894
R1397 VP.n36 VP.n18 0.189894
R1398 VP.n40 VP.n18 0.189894
R1399 VP.n41 VP.n40 0.189894
R1400 VP.n42 VP.n41 0.189894
R1401 VP.n42 VP.n16 0.189894
R1402 VP.n47 VP.n16 0.189894
R1403 VP.n48 VP.n47 0.189894
R1404 VP.n49 VP.n48 0.189894
R1405 VP.n49 VP.n14 0.189894
R1406 VP.n53 VP.n14 0.189894
R1407 VP.n58 VP.n57 0.189894
R1408 VP.n58 VP.n11 0.189894
R1409 VP.n62 VP.n11 0.189894
R1410 VP.n63 VP.n62 0.189894
R1411 VP.n64 VP.n63 0.189894
R1412 VP.n64 VP.n9 0.189894
R1413 VP.n69 VP.n9 0.189894
R1414 VP.n70 VP.n69 0.189894
R1415 VP.n71 VP.n70 0.189894
R1416 VP.n71 VP.n7 0.189894
R1417 VP.n76 VP.n7 0.189894
R1418 VP.n77 VP.n76 0.189894
R1419 VP.n78 VP.n77 0.189894
R1420 VP.n78 VP.n5 0.189894
R1421 VP.n82 VP.n5 0.189894
R1422 VP.n83 VP.n82 0.189894
R1423 VP.n84 VP.n83 0.189894
R1424 VP.n84 VP.n3 0.189894
R1425 VP.n89 VP.n3 0.189894
R1426 VP.n90 VP.n89 0.189894
R1427 VP.n91 VP.n90 0.189894
R1428 VP.n91 VP.n1 0.189894
R1429 VP.n95 VP.n1 0.189894
R1430 VTAIL.n11 VTAIL.t0 61.4127
R1431 VTAIL.n16 VTAIL.t11 61.4125
R1432 VTAIL.n17 VTAIL.t8 61.4125
R1433 VTAIL.n2 VTAIL.t12 61.4125
R1434 VTAIL.n15 VTAIL.n14 58.2384
R1435 VTAIL.n13 VTAIL.n12 58.2384
R1436 VTAIL.n10 VTAIL.n9 58.2384
R1437 VTAIL.n8 VTAIL.n7 58.2384
R1438 VTAIL.n19 VTAIL.n18 58.2381
R1439 VTAIL.n1 VTAIL.n0 58.2381
R1440 VTAIL.n4 VTAIL.n3 58.2381
R1441 VTAIL.n6 VTAIL.n5 58.2381
R1442 VTAIL.n8 VTAIL.n6 26.5565
R1443 VTAIL.n17 VTAIL.n16 23.8755
R1444 VTAIL.n18 VTAIL.t7 3.17482
R1445 VTAIL.n18 VTAIL.t3 3.17482
R1446 VTAIL.n0 VTAIL.t9 3.17482
R1447 VTAIL.n0 VTAIL.t5 3.17482
R1448 VTAIL.n3 VTAIL.t10 3.17482
R1449 VTAIL.n3 VTAIL.t17 3.17482
R1450 VTAIL.n5 VTAIL.t16 3.17482
R1451 VTAIL.n5 VTAIL.t14 3.17482
R1452 VTAIL.n14 VTAIL.t18 3.17482
R1453 VTAIL.n14 VTAIL.t15 3.17482
R1454 VTAIL.n12 VTAIL.t13 3.17482
R1455 VTAIL.n12 VTAIL.t19 3.17482
R1456 VTAIL.n9 VTAIL.t2 3.17482
R1457 VTAIL.n9 VTAIL.t6 3.17482
R1458 VTAIL.n7 VTAIL.t1 3.17482
R1459 VTAIL.n7 VTAIL.t4 3.17482
R1460 VTAIL.n10 VTAIL.n8 2.68153
R1461 VTAIL.n11 VTAIL.n10 2.68153
R1462 VTAIL.n15 VTAIL.n13 2.68153
R1463 VTAIL.n16 VTAIL.n15 2.68153
R1464 VTAIL.n6 VTAIL.n4 2.68153
R1465 VTAIL.n4 VTAIL.n2 2.68153
R1466 VTAIL.n19 VTAIL.n17 2.68153
R1467 VTAIL VTAIL.n1 2.06947
R1468 VTAIL.n13 VTAIL.n11 1.81084
R1469 VTAIL.n2 VTAIL.n1 1.81084
R1470 VTAIL VTAIL.n19 0.612569
R1471 VDD1.n1 VDD1.t6 80.7725
R1472 VDD1.n3 VDD1.t3 80.7723
R1473 VDD1.n5 VDD1.n4 76.8724
R1474 VDD1.n1 VDD1.n0 74.9172
R1475 VDD1.n7 VDD1.n6 74.917
R1476 VDD1.n3 VDD1.n2 74.9169
R1477 VDD1.n7 VDD1.n5 47.2013
R1478 VDD1.n6 VDD1.t4 3.17482
R1479 VDD1.n6 VDD1.t8 3.17482
R1480 VDD1.n0 VDD1.t0 3.17482
R1481 VDD1.n0 VDD1.t1 3.17482
R1482 VDD1.n4 VDD1.t2 3.17482
R1483 VDD1.n4 VDD1.t7 3.17482
R1484 VDD1.n2 VDD1.t5 3.17482
R1485 VDD1.n2 VDD1.t9 3.17482
R1486 VDD1 VDD1.n7 1.95309
R1487 VDD1 VDD1.n1 0.728948
R1488 VDD1.n5 VDD1.n3 0.615413
R1489 VN.n82 VN.n81 161.3
R1490 VN.n80 VN.n43 161.3
R1491 VN.n79 VN.n78 161.3
R1492 VN.n77 VN.n44 161.3
R1493 VN.n76 VN.n75 161.3
R1494 VN.n74 VN.n45 161.3
R1495 VN.n72 VN.n71 161.3
R1496 VN.n70 VN.n46 161.3
R1497 VN.n69 VN.n68 161.3
R1498 VN.n67 VN.n47 161.3
R1499 VN.n66 VN.n65 161.3
R1500 VN.n64 VN.n48 161.3
R1501 VN.n63 VN.n62 161.3
R1502 VN.n61 VN.n49 161.3
R1503 VN.n60 VN.n59 161.3
R1504 VN.n58 VN.n51 161.3
R1505 VN.n57 VN.n56 161.3
R1506 VN.n55 VN.n52 161.3
R1507 VN.n40 VN.n39 161.3
R1508 VN.n38 VN.n1 161.3
R1509 VN.n37 VN.n36 161.3
R1510 VN.n35 VN.n2 161.3
R1511 VN.n34 VN.n33 161.3
R1512 VN.n32 VN.n3 161.3
R1513 VN.n30 VN.n29 161.3
R1514 VN.n28 VN.n4 161.3
R1515 VN.n27 VN.n26 161.3
R1516 VN.n25 VN.n5 161.3
R1517 VN.n24 VN.n23 161.3
R1518 VN.n22 VN.n6 161.3
R1519 VN.n21 VN.n20 161.3
R1520 VN.n18 VN.n7 161.3
R1521 VN.n17 VN.n16 161.3
R1522 VN.n15 VN.n8 161.3
R1523 VN.n14 VN.n13 161.3
R1524 VN.n12 VN.n9 161.3
R1525 VN.n53 VN.t3 120.678
R1526 VN.n10 VN.t1 120.678
R1527 VN.n11 VN.t9 88.7717
R1528 VN.n19 VN.t0 88.7717
R1529 VN.n31 VN.t2 88.7717
R1530 VN.n0 VN.t6 88.7717
R1531 VN.n54 VN.t4 88.7717
R1532 VN.n50 VN.t5 88.7717
R1533 VN.n73 VN.t7 88.7717
R1534 VN.n42 VN.t8 88.7717
R1535 VN.n41 VN.n0 67.0082
R1536 VN.n83 VN.n42 67.0082
R1537 VN.n17 VN.n8 56.4773
R1538 VN.n26 VN.n25 56.4773
R1539 VN.n60 VN.n51 56.4773
R1540 VN.n68 VN.n67 56.4773
R1541 VN.n11 VN.n10 55.8591
R1542 VN.n54 VN.n53 55.8591
R1543 VN VN.n83 53.0396
R1544 VN.n37 VN.n2 48.6874
R1545 VN.n79 VN.n44 48.6874
R1546 VN.n38 VN.n37 32.1338
R1547 VN.n80 VN.n79 32.1338
R1548 VN.n13 VN.n12 24.3439
R1549 VN.n13 VN.n8 24.3439
R1550 VN.n18 VN.n17 24.3439
R1551 VN.n20 VN.n18 24.3439
R1552 VN.n24 VN.n6 24.3439
R1553 VN.n25 VN.n24 24.3439
R1554 VN.n26 VN.n4 24.3439
R1555 VN.n30 VN.n4 24.3439
R1556 VN.n33 VN.n32 24.3439
R1557 VN.n33 VN.n2 24.3439
R1558 VN.n39 VN.n38 24.3439
R1559 VN.n56 VN.n51 24.3439
R1560 VN.n56 VN.n55 24.3439
R1561 VN.n67 VN.n66 24.3439
R1562 VN.n66 VN.n48 24.3439
R1563 VN.n62 VN.n61 24.3439
R1564 VN.n61 VN.n60 24.3439
R1565 VN.n75 VN.n44 24.3439
R1566 VN.n75 VN.n74 24.3439
R1567 VN.n72 VN.n46 24.3439
R1568 VN.n68 VN.n46 24.3439
R1569 VN.n81 VN.n80 24.3439
R1570 VN.n39 VN.n0 22.8833
R1571 VN.n81 VN.n42 22.8833
R1572 VN.n12 VN.n11 17.5278
R1573 VN.n31 VN.n30 17.5278
R1574 VN.n55 VN.n54 17.5278
R1575 VN.n73 VN.n72 17.5278
R1576 VN.n20 VN.n19 12.1722
R1577 VN.n19 VN.n6 12.1722
R1578 VN.n50 VN.n48 12.1722
R1579 VN.n62 VN.n50 12.1722
R1580 VN.n32 VN.n31 6.81666
R1581 VN.n74 VN.n73 6.81666
R1582 VN.n53 VN.n52 5.32599
R1583 VN.n10 VN.n9 5.32599
R1584 VN.n83 VN.n82 0.355081
R1585 VN.n41 VN.n40 0.355081
R1586 VN VN.n41 0.26685
R1587 VN.n82 VN.n43 0.189894
R1588 VN.n78 VN.n43 0.189894
R1589 VN.n78 VN.n77 0.189894
R1590 VN.n77 VN.n76 0.189894
R1591 VN.n76 VN.n45 0.189894
R1592 VN.n71 VN.n45 0.189894
R1593 VN.n71 VN.n70 0.189894
R1594 VN.n70 VN.n69 0.189894
R1595 VN.n69 VN.n47 0.189894
R1596 VN.n65 VN.n47 0.189894
R1597 VN.n65 VN.n64 0.189894
R1598 VN.n64 VN.n63 0.189894
R1599 VN.n63 VN.n49 0.189894
R1600 VN.n59 VN.n49 0.189894
R1601 VN.n59 VN.n58 0.189894
R1602 VN.n58 VN.n57 0.189894
R1603 VN.n57 VN.n52 0.189894
R1604 VN.n14 VN.n9 0.189894
R1605 VN.n15 VN.n14 0.189894
R1606 VN.n16 VN.n15 0.189894
R1607 VN.n16 VN.n7 0.189894
R1608 VN.n21 VN.n7 0.189894
R1609 VN.n22 VN.n21 0.189894
R1610 VN.n23 VN.n22 0.189894
R1611 VN.n23 VN.n5 0.189894
R1612 VN.n27 VN.n5 0.189894
R1613 VN.n28 VN.n27 0.189894
R1614 VN.n29 VN.n28 0.189894
R1615 VN.n29 VN.n3 0.189894
R1616 VN.n34 VN.n3 0.189894
R1617 VN.n35 VN.n34 0.189894
R1618 VN.n36 VN.n35 0.189894
R1619 VN.n36 VN.n1 0.189894
R1620 VN.n40 VN.n1 0.189894
R1621 VDD2.n1 VDD2.t8 80.7723
R1622 VDD2.n4 VDD2.t1 78.0915
R1623 VDD2.n3 VDD2.n2 76.8724
R1624 VDD2 VDD2.n7 76.8696
R1625 VDD2.n6 VDD2.n5 74.9172
R1626 VDD2.n1 VDD2.n0 74.9169
R1627 VDD2.n4 VDD2.n3 45.2778
R1628 VDD2.n7 VDD2.t5 3.17482
R1629 VDD2.n7 VDD2.t6 3.17482
R1630 VDD2.n5 VDD2.t2 3.17482
R1631 VDD2.n5 VDD2.t4 3.17482
R1632 VDD2.n2 VDD2.t7 3.17482
R1633 VDD2.n2 VDD2.t3 3.17482
R1634 VDD2.n0 VDD2.t0 3.17482
R1635 VDD2.n0 VDD2.t9 3.17482
R1636 VDD2.n6 VDD2.n4 2.68153
R1637 VDD2 VDD2.n6 0.728948
R1638 VDD2.n3 VDD2.n1 0.615413
C0 VTAIL w_n4702_n3016# 2.99299f
C1 VDD1 w_n4702_n3016# 2.73611f
C2 VN VDD2 9.29645f
C3 B w_n4702_n3016# 10.3563f
C4 VN w_n4702_n3016# 10.0994f
C5 VDD2 w_n4702_n3016# 2.88902f
C6 VTAIL VP 10.108f
C7 VP VDD1 9.74552f
C8 VTAIL VDD1 9.65458f
C9 VP B 2.33584f
C10 VTAIL B 3.40551f
C11 B VDD1 2.41119f
C12 VP VN 8.34888f
C13 VTAIL VN 10.0937f
C14 VDD1 VN 0.153451f
C15 VP VDD2 0.606086f
C16 B VN 1.3045f
C17 VTAIL VDD2 9.7073f
C18 VDD1 VDD2 2.29149f
C19 VP w_n4702_n3016# 10.7122f
C20 B VDD2 2.53612f
C21 VDD2 VSUBS 2.215161f
C22 VDD1 VSUBS 1.989924f
C23 VTAIL VSUBS 1.284797f
C24 VN VSUBS 7.94382f
C25 VP VSUBS 4.417873f
C26 B VSUBS 5.442975f
C27 w_n4702_n3016# VSUBS 0.175084p
C28 VDD2.t8 VSUBS 2.5198f
C29 VDD2.t0 VSUBS 0.251126f
C30 VDD2.t9 VSUBS 0.251126f
C31 VDD2.n0 VSUBS 1.89832f
C32 VDD2.n1 VSUBS 1.81508f
C33 VDD2.t7 VSUBS 0.251126f
C34 VDD2.t3 VSUBS 0.251126f
C35 VDD2.n2 VSUBS 1.92494f
C36 VDD2.n3 VSUBS 3.89871f
C37 VDD2.t1 VSUBS 2.48842f
C38 VDD2.n4 VSUBS 4.12387f
C39 VDD2.t2 VSUBS 0.251126f
C40 VDD2.t4 VSUBS 0.251126f
C41 VDD2.n5 VSUBS 1.89832f
C42 VDD2.n6 VSUBS 0.911093f
C43 VDD2.t5 VSUBS 0.251126f
C44 VDD2.t6 VSUBS 0.251126f
C45 VDD2.n7 VSUBS 1.92488f
C46 VN.t6 VSUBS 2.2063f
C47 VN.n0 VSUBS 0.898737f
C48 VN.n1 VSUBS 0.028586f
C49 VN.n2 VSUBS 0.053544f
C50 VN.n3 VSUBS 0.028586f
C51 VN.t2 VSUBS 2.2063f
C52 VN.n4 VSUBS 0.053544f
C53 VN.n5 VSUBS 0.028586f
C54 VN.n6 VSUBS 0.040326f
C55 VN.n7 VSUBS 0.028586f
C56 VN.n8 VSUBS 0.0375f
C57 VN.n9 VSUBS 0.300345f
C58 VN.t9 VSUBS 2.2063f
C59 VN.t1 VSUBS 2.4639f
C60 VN.n10 VSUBS 0.849312f
C61 VN.n11 VSUBS 0.880507f
C62 VN.n12 VSUBS 0.046142f
C63 VN.n13 VSUBS 0.053544f
C64 VN.n14 VSUBS 0.028586f
C65 VN.n15 VSUBS 0.028586f
C66 VN.n16 VSUBS 0.028586f
C67 VN.n17 VSUBS 0.046324f
C68 VN.n18 VSUBS 0.053544f
C69 VN.t0 VSUBS 2.2063f
C70 VN.n19 VSUBS 0.786616f
C71 VN.n20 VSUBS 0.040326f
C72 VN.n21 VSUBS 0.028586f
C73 VN.n22 VSUBS 0.028586f
C74 VN.n23 VSUBS 0.028586f
C75 VN.n24 VSUBS 0.053544f
C76 VN.n25 VSUBS 0.046324f
C77 VN.n26 VSUBS 0.0375f
C78 VN.n27 VSUBS 0.028586f
C79 VN.n28 VSUBS 0.028586f
C80 VN.n29 VSUBS 0.028586f
C81 VN.n30 VSUBS 0.046142f
C82 VN.n31 VSUBS 0.786616f
C83 VN.n32 VSUBS 0.03451f
C84 VN.n33 VSUBS 0.053544f
C85 VN.n34 VSUBS 0.028586f
C86 VN.n35 VSUBS 0.028586f
C87 VN.n36 VSUBS 0.028586f
C88 VN.n37 VSUBS 0.025922f
C89 VN.n38 VSUBS 0.057902f
C90 VN.n39 VSUBS 0.051958f
C91 VN.n40 VSUBS 0.046144f
C92 VN.n41 VSUBS 0.053631f
C93 VN.t8 VSUBS 2.2063f
C94 VN.n42 VSUBS 0.898737f
C95 VN.n43 VSUBS 0.028586f
C96 VN.n44 VSUBS 0.053544f
C97 VN.n45 VSUBS 0.028586f
C98 VN.t7 VSUBS 2.2063f
C99 VN.n46 VSUBS 0.053544f
C100 VN.n47 VSUBS 0.028586f
C101 VN.n48 VSUBS 0.040326f
C102 VN.n49 VSUBS 0.028586f
C103 VN.t5 VSUBS 2.2063f
C104 VN.n50 VSUBS 0.786616f
C105 VN.n51 VSUBS 0.0375f
C106 VN.n52 VSUBS 0.300345f
C107 VN.t4 VSUBS 2.2063f
C108 VN.t3 VSUBS 2.4639f
C109 VN.n53 VSUBS 0.849312f
C110 VN.n54 VSUBS 0.880507f
C111 VN.n55 VSUBS 0.046142f
C112 VN.n56 VSUBS 0.053544f
C113 VN.n57 VSUBS 0.028586f
C114 VN.n58 VSUBS 0.028586f
C115 VN.n59 VSUBS 0.028586f
C116 VN.n60 VSUBS 0.046324f
C117 VN.n61 VSUBS 0.053544f
C118 VN.n62 VSUBS 0.040326f
C119 VN.n63 VSUBS 0.028586f
C120 VN.n64 VSUBS 0.028586f
C121 VN.n65 VSUBS 0.028586f
C122 VN.n66 VSUBS 0.053544f
C123 VN.n67 VSUBS 0.046324f
C124 VN.n68 VSUBS 0.0375f
C125 VN.n69 VSUBS 0.028586f
C126 VN.n70 VSUBS 0.028586f
C127 VN.n71 VSUBS 0.028586f
C128 VN.n72 VSUBS 0.046142f
C129 VN.n73 VSUBS 0.786616f
C130 VN.n74 VSUBS 0.03451f
C131 VN.n75 VSUBS 0.053544f
C132 VN.n76 VSUBS 0.028586f
C133 VN.n77 VSUBS 0.028586f
C134 VN.n78 VSUBS 0.028586f
C135 VN.n79 VSUBS 0.025922f
C136 VN.n80 VSUBS 0.057902f
C137 VN.n81 VSUBS 0.051958f
C138 VN.n82 VSUBS 0.046144f
C139 VN.n83 VSUBS 1.75481f
C140 VDD1.t6 VSUBS 2.51843f
C141 VDD1.t0 VSUBS 0.250989f
C142 VDD1.t1 VSUBS 0.250989f
C143 VDD1.n0 VSUBS 1.89729f
C144 VDD1.n1 VSUBS 1.82426f
C145 VDD1.t3 VSUBS 2.51842f
C146 VDD1.t5 VSUBS 0.250989f
C147 VDD1.t9 VSUBS 0.250989f
C148 VDD1.n2 VSUBS 1.89728f
C149 VDD1.n3 VSUBS 1.81409f
C150 VDD1.t2 VSUBS 0.250989f
C151 VDD1.t7 VSUBS 0.250989f
C152 VDD1.n4 VSUBS 1.92389f
C153 VDD1.n5 VSUBS 4.05616f
C154 VDD1.t4 VSUBS 0.250989f
C155 VDD1.t8 VSUBS 0.250989f
C156 VDD1.n6 VSUBS 1.89728f
C157 VDD1.n7 VSUBS 4.17702f
C158 VTAIL.t9 VSUBS 0.242112f
C159 VTAIL.t5 VSUBS 0.242112f
C160 VTAIL.n0 VSUBS 1.67438f
C161 VTAIL.n1 VSUBS 1.03882f
C162 VTAIL.t12 VSUBS 2.22653f
C163 VTAIL.n2 VSUBS 1.20599f
C164 VTAIL.t10 VSUBS 0.242112f
C165 VTAIL.t17 VSUBS 0.242112f
C166 VTAIL.n3 VSUBS 1.67438f
C167 VTAIL.n4 VSUBS 1.18177f
C168 VTAIL.t16 VSUBS 0.242112f
C169 VTAIL.t14 VSUBS 0.242112f
C170 VTAIL.n5 VSUBS 1.67438f
C171 VTAIL.n6 VSUBS 2.69774f
C172 VTAIL.t1 VSUBS 0.242112f
C173 VTAIL.t4 VSUBS 0.242112f
C174 VTAIL.n7 VSUBS 1.67439f
C175 VTAIL.n8 VSUBS 2.69773f
C176 VTAIL.t2 VSUBS 0.242112f
C177 VTAIL.t6 VSUBS 0.242112f
C178 VTAIL.n9 VSUBS 1.67439f
C179 VTAIL.n10 VSUBS 1.18176f
C180 VTAIL.t0 VSUBS 2.22653f
C181 VTAIL.n11 VSUBS 1.20598f
C182 VTAIL.t13 VSUBS 0.242112f
C183 VTAIL.t19 VSUBS 0.242112f
C184 VTAIL.n12 VSUBS 1.67439f
C185 VTAIL.n13 VSUBS 1.09782f
C186 VTAIL.t18 VSUBS 0.242112f
C187 VTAIL.t15 VSUBS 0.242112f
C188 VTAIL.n14 VSUBS 1.67439f
C189 VTAIL.n15 VSUBS 1.18176f
C190 VTAIL.t11 VSUBS 2.22653f
C191 VTAIL.n16 VSUBS 2.54742f
C192 VTAIL.t8 VSUBS 2.22653f
C193 VTAIL.n17 VSUBS 2.54742f
C194 VTAIL.t7 VSUBS 0.242112f
C195 VTAIL.t3 VSUBS 0.242112f
C196 VTAIL.n18 VSUBS 1.67438f
C197 VTAIL.n19 VSUBS 0.982303f
C198 VP.t2 VSUBS 2.40147f
C199 VP.n0 VSUBS 0.978238f
C200 VP.n1 VSUBS 0.031115f
C201 VP.n2 VSUBS 0.05828f
C202 VP.n3 VSUBS 0.031115f
C203 VP.t7 VSUBS 2.40147f
C204 VP.n4 VSUBS 0.05828f
C205 VP.n5 VSUBS 0.031115f
C206 VP.n6 VSUBS 0.043893f
C207 VP.n7 VSUBS 0.031115f
C208 VP.n8 VSUBS 0.040817f
C209 VP.n9 VSUBS 0.031115f
C210 VP.t4 VSUBS 2.40147f
C211 VP.n10 VSUBS 0.05828f
C212 VP.n11 VSUBS 0.031115f
C213 VP.n12 VSUBS 0.056554f
C214 VP.t1 VSUBS 2.40147f
C215 VP.n13 VSUBS 0.978238f
C216 VP.n14 VSUBS 0.031115f
C217 VP.n15 VSUBS 0.05828f
C218 VP.n16 VSUBS 0.031115f
C219 VP.t5 VSUBS 2.40147f
C220 VP.n17 VSUBS 0.05828f
C221 VP.n18 VSUBS 0.031115f
C222 VP.n19 VSUBS 0.043893f
C223 VP.n20 VSUBS 0.031115f
C224 VP.n21 VSUBS 0.040817f
C225 VP.n22 VSUBS 0.326914f
C226 VP.t9 VSUBS 2.40147f
C227 VP.t3 VSUBS 2.68185f
C228 VP.n23 VSUBS 0.924442f
C229 VP.n24 VSUBS 0.958396f
C230 VP.n25 VSUBS 0.050223f
C231 VP.n26 VSUBS 0.05828f
C232 VP.n27 VSUBS 0.031115f
C233 VP.n28 VSUBS 0.031115f
C234 VP.n29 VSUBS 0.031115f
C235 VP.n30 VSUBS 0.050422f
C236 VP.n31 VSUBS 0.05828f
C237 VP.t8 VSUBS 2.40147f
C238 VP.n32 VSUBS 0.856199f
C239 VP.n33 VSUBS 0.043893f
C240 VP.n34 VSUBS 0.031115f
C241 VP.n35 VSUBS 0.031115f
C242 VP.n36 VSUBS 0.031115f
C243 VP.n37 VSUBS 0.05828f
C244 VP.n38 VSUBS 0.050422f
C245 VP.n39 VSUBS 0.040817f
C246 VP.n40 VSUBS 0.031115f
C247 VP.n41 VSUBS 0.031115f
C248 VP.n42 VSUBS 0.031115f
C249 VP.n43 VSUBS 0.050223f
C250 VP.n44 VSUBS 0.856199f
C251 VP.n45 VSUBS 0.037562f
C252 VP.n46 VSUBS 0.05828f
C253 VP.n47 VSUBS 0.031115f
C254 VP.n48 VSUBS 0.031115f
C255 VP.n49 VSUBS 0.031115f
C256 VP.n50 VSUBS 0.028215f
C257 VP.n51 VSUBS 0.063024f
C258 VP.n52 VSUBS 0.056554f
C259 VP.n53 VSUBS 0.050226f
C260 VP.n54 VSUBS 1.89753f
C261 VP.t6 VSUBS 2.40147f
C262 VP.n55 VSUBS 0.978238f
C263 VP.n56 VSUBS 1.91862f
C264 VP.n57 VSUBS 0.050226f
C265 VP.n58 VSUBS 0.031115f
C266 VP.n59 VSUBS 0.063024f
C267 VP.n60 VSUBS 0.028215f
C268 VP.n61 VSUBS 0.05828f
C269 VP.n62 VSUBS 0.031115f
C270 VP.n63 VSUBS 0.031115f
C271 VP.n64 VSUBS 0.031115f
C272 VP.n65 VSUBS 0.037562f
C273 VP.n66 VSUBS 0.856199f
C274 VP.n67 VSUBS 0.050223f
C275 VP.n68 VSUBS 0.05828f
C276 VP.n69 VSUBS 0.031115f
C277 VP.n70 VSUBS 0.031115f
C278 VP.n71 VSUBS 0.031115f
C279 VP.n72 VSUBS 0.050422f
C280 VP.n73 VSUBS 0.05828f
C281 VP.t0 VSUBS 2.40147f
C282 VP.n74 VSUBS 0.856199f
C283 VP.n75 VSUBS 0.043893f
C284 VP.n76 VSUBS 0.031115f
C285 VP.n77 VSUBS 0.031115f
C286 VP.n78 VSUBS 0.031115f
C287 VP.n79 VSUBS 0.05828f
C288 VP.n80 VSUBS 0.050422f
C289 VP.n81 VSUBS 0.040817f
C290 VP.n82 VSUBS 0.031115f
C291 VP.n83 VSUBS 0.031115f
C292 VP.n84 VSUBS 0.031115f
C293 VP.n85 VSUBS 0.050223f
C294 VP.n86 VSUBS 0.856199f
C295 VP.n87 VSUBS 0.037562f
C296 VP.n88 VSUBS 0.05828f
C297 VP.n89 VSUBS 0.031115f
C298 VP.n90 VSUBS 0.031115f
C299 VP.n91 VSUBS 0.031115f
C300 VP.n92 VSUBS 0.028215f
C301 VP.n93 VSUBS 0.063024f
C302 VP.n94 VSUBS 0.056554f
C303 VP.n95 VSUBS 0.050226f
C304 VP.n96 VSUBS 0.058375f
C305 B.n0 VSUBS 0.006164f
C306 B.n1 VSUBS 0.006164f
C307 B.n2 VSUBS 0.009748f
C308 B.n3 VSUBS 0.009748f
C309 B.n4 VSUBS 0.009748f
C310 B.n5 VSUBS 0.009748f
C311 B.n6 VSUBS 0.009748f
C312 B.n7 VSUBS 0.009748f
C313 B.n8 VSUBS 0.009748f
C314 B.n9 VSUBS 0.009748f
C315 B.n10 VSUBS 0.009748f
C316 B.n11 VSUBS 0.009748f
C317 B.n12 VSUBS 0.009748f
C318 B.n13 VSUBS 0.009748f
C319 B.n14 VSUBS 0.009748f
C320 B.n15 VSUBS 0.009748f
C321 B.n16 VSUBS 0.009748f
C322 B.n17 VSUBS 0.009748f
C323 B.n18 VSUBS 0.009748f
C324 B.n19 VSUBS 0.009748f
C325 B.n20 VSUBS 0.009748f
C326 B.n21 VSUBS 0.009748f
C327 B.n22 VSUBS 0.009748f
C328 B.n23 VSUBS 0.009748f
C329 B.n24 VSUBS 0.009748f
C330 B.n25 VSUBS 0.009748f
C331 B.n26 VSUBS 0.009748f
C332 B.n27 VSUBS 0.009748f
C333 B.n28 VSUBS 0.009748f
C334 B.n29 VSUBS 0.009748f
C335 B.n30 VSUBS 0.009748f
C336 B.n31 VSUBS 0.009748f
C337 B.n32 VSUBS 0.009748f
C338 B.n33 VSUBS 0.023494f
C339 B.n34 VSUBS 0.009748f
C340 B.n35 VSUBS 0.009748f
C341 B.n36 VSUBS 0.009748f
C342 B.n37 VSUBS 0.009748f
C343 B.n38 VSUBS 0.009748f
C344 B.n39 VSUBS 0.009748f
C345 B.n40 VSUBS 0.009748f
C346 B.n41 VSUBS 0.009748f
C347 B.n42 VSUBS 0.009748f
C348 B.n43 VSUBS 0.009748f
C349 B.n44 VSUBS 0.009748f
C350 B.n45 VSUBS 0.009748f
C351 B.n46 VSUBS 0.009748f
C352 B.n47 VSUBS 0.009748f
C353 B.n48 VSUBS 0.009748f
C354 B.n49 VSUBS 0.009748f
C355 B.n50 VSUBS 0.009748f
C356 B.n51 VSUBS 0.009748f
C357 B.t8 VSUBS 0.456179f
C358 B.t7 VSUBS 0.487262f
C359 B.t6 VSUBS 1.83074f
C360 B.n52 VSUBS 0.259322f
C361 B.n53 VSUBS 0.100826f
C362 B.n54 VSUBS 0.009748f
C363 B.n55 VSUBS 0.009748f
C364 B.n56 VSUBS 0.009748f
C365 B.n57 VSUBS 0.009748f
C366 B.n58 VSUBS 0.005448f
C367 B.n59 VSUBS 0.009748f
C368 B.t5 VSUBS 0.456173f
C369 B.t4 VSUBS 0.487256f
C370 B.t3 VSUBS 1.83074f
C371 B.n60 VSUBS 0.259329f
C372 B.n61 VSUBS 0.100833f
C373 B.n62 VSUBS 0.022586f
C374 B.n63 VSUBS 0.009748f
C375 B.n64 VSUBS 0.009748f
C376 B.n65 VSUBS 0.009748f
C377 B.n66 VSUBS 0.009748f
C378 B.n67 VSUBS 0.009748f
C379 B.n68 VSUBS 0.009748f
C380 B.n69 VSUBS 0.009748f
C381 B.n70 VSUBS 0.009748f
C382 B.n71 VSUBS 0.009748f
C383 B.n72 VSUBS 0.009748f
C384 B.n73 VSUBS 0.009748f
C385 B.n74 VSUBS 0.009748f
C386 B.n75 VSUBS 0.009748f
C387 B.n76 VSUBS 0.009748f
C388 B.n77 VSUBS 0.009748f
C389 B.n78 VSUBS 0.009748f
C390 B.n79 VSUBS 0.02302f
C391 B.n80 VSUBS 0.009748f
C392 B.n81 VSUBS 0.009748f
C393 B.n82 VSUBS 0.009748f
C394 B.n83 VSUBS 0.009748f
C395 B.n84 VSUBS 0.009748f
C396 B.n85 VSUBS 0.009748f
C397 B.n86 VSUBS 0.009748f
C398 B.n87 VSUBS 0.009748f
C399 B.n88 VSUBS 0.009748f
C400 B.n89 VSUBS 0.009748f
C401 B.n90 VSUBS 0.009748f
C402 B.n91 VSUBS 0.009748f
C403 B.n92 VSUBS 0.009748f
C404 B.n93 VSUBS 0.009748f
C405 B.n94 VSUBS 0.009748f
C406 B.n95 VSUBS 0.009748f
C407 B.n96 VSUBS 0.009748f
C408 B.n97 VSUBS 0.009748f
C409 B.n98 VSUBS 0.009748f
C410 B.n99 VSUBS 0.009748f
C411 B.n100 VSUBS 0.009748f
C412 B.n101 VSUBS 0.009748f
C413 B.n102 VSUBS 0.009748f
C414 B.n103 VSUBS 0.009748f
C415 B.n104 VSUBS 0.009748f
C416 B.n105 VSUBS 0.009748f
C417 B.n106 VSUBS 0.009748f
C418 B.n107 VSUBS 0.009748f
C419 B.n108 VSUBS 0.009748f
C420 B.n109 VSUBS 0.009748f
C421 B.n110 VSUBS 0.009748f
C422 B.n111 VSUBS 0.009748f
C423 B.n112 VSUBS 0.009748f
C424 B.n113 VSUBS 0.009748f
C425 B.n114 VSUBS 0.009748f
C426 B.n115 VSUBS 0.009748f
C427 B.n116 VSUBS 0.009748f
C428 B.n117 VSUBS 0.009748f
C429 B.n118 VSUBS 0.009748f
C430 B.n119 VSUBS 0.009748f
C431 B.n120 VSUBS 0.009748f
C432 B.n121 VSUBS 0.009748f
C433 B.n122 VSUBS 0.009748f
C434 B.n123 VSUBS 0.009748f
C435 B.n124 VSUBS 0.009748f
C436 B.n125 VSUBS 0.009748f
C437 B.n126 VSUBS 0.009748f
C438 B.n127 VSUBS 0.009748f
C439 B.n128 VSUBS 0.009748f
C440 B.n129 VSUBS 0.009748f
C441 B.n130 VSUBS 0.009748f
C442 B.n131 VSUBS 0.009748f
C443 B.n132 VSUBS 0.009748f
C444 B.n133 VSUBS 0.009748f
C445 B.n134 VSUBS 0.009748f
C446 B.n135 VSUBS 0.009748f
C447 B.n136 VSUBS 0.009748f
C448 B.n137 VSUBS 0.009748f
C449 B.n138 VSUBS 0.009748f
C450 B.n139 VSUBS 0.009748f
C451 B.n140 VSUBS 0.009748f
C452 B.n141 VSUBS 0.009748f
C453 B.n142 VSUBS 0.009748f
C454 B.n143 VSUBS 0.0241f
C455 B.n144 VSUBS 0.009748f
C456 B.n145 VSUBS 0.009748f
C457 B.n146 VSUBS 0.009748f
C458 B.n147 VSUBS 0.009748f
C459 B.n148 VSUBS 0.009748f
C460 B.n149 VSUBS 0.009748f
C461 B.n150 VSUBS 0.009748f
C462 B.n151 VSUBS 0.009748f
C463 B.n152 VSUBS 0.009748f
C464 B.n153 VSUBS 0.009748f
C465 B.n154 VSUBS 0.009748f
C466 B.n155 VSUBS 0.009748f
C467 B.n156 VSUBS 0.009748f
C468 B.n157 VSUBS 0.009748f
C469 B.n158 VSUBS 0.009748f
C470 B.n159 VSUBS 0.009748f
C471 B.n160 VSUBS 0.009748f
C472 B.t1 VSUBS 0.456173f
C473 B.t2 VSUBS 0.487256f
C474 B.t0 VSUBS 1.83074f
C475 B.n161 VSUBS 0.259329f
C476 B.n162 VSUBS 0.100833f
C477 B.n163 VSUBS 0.022586f
C478 B.n164 VSUBS 0.009748f
C479 B.n165 VSUBS 0.009748f
C480 B.n166 VSUBS 0.009748f
C481 B.n167 VSUBS 0.009748f
C482 B.n168 VSUBS 0.009748f
C483 B.t10 VSUBS 0.456179f
C484 B.t11 VSUBS 0.487262f
C485 B.t9 VSUBS 1.83074f
C486 B.n169 VSUBS 0.259322f
C487 B.n170 VSUBS 0.100826f
C488 B.n171 VSUBS 0.009748f
C489 B.n172 VSUBS 0.009748f
C490 B.n173 VSUBS 0.009748f
C491 B.n174 VSUBS 0.009748f
C492 B.n175 VSUBS 0.009748f
C493 B.n176 VSUBS 0.009748f
C494 B.n177 VSUBS 0.009748f
C495 B.n178 VSUBS 0.009748f
C496 B.n179 VSUBS 0.009748f
C497 B.n180 VSUBS 0.009748f
C498 B.n181 VSUBS 0.009748f
C499 B.n182 VSUBS 0.009748f
C500 B.n183 VSUBS 0.009748f
C501 B.n184 VSUBS 0.009748f
C502 B.n185 VSUBS 0.009748f
C503 B.n186 VSUBS 0.009748f
C504 B.n187 VSUBS 0.009748f
C505 B.n188 VSUBS 0.0241f
C506 B.n189 VSUBS 0.009748f
C507 B.n190 VSUBS 0.009748f
C508 B.n191 VSUBS 0.009748f
C509 B.n192 VSUBS 0.009748f
C510 B.n193 VSUBS 0.009748f
C511 B.n194 VSUBS 0.009748f
C512 B.n195 VSUBS 0.009748f
C513 B.n196 VSUBS 0.009748f
C514 B.n197 VSUBS 0.009748f
C515 B.n198 VSUBS 0.009748f
C516 B.n199 VSUBS 0.009748f
C517 B.n200 VSUBS 0.009748f
C518 B.n201 VSUBS 0.009748f
C519 B.n202 VSUBS 0.009748f
C520 B.n203 VSUBS 0.009748f
C521 B.n204 VSUBS 0.009748f
C522 B.n205 VSUBS 0.009748f
C523 B.n206 VSUBS 0.009748f
C524 B.n207 VSUBS 0.009748f
C525 B.n208 VSUBS 0.009748f
C526 B.n209 VSUBS 0.009748f
C527 B.n210 VSUBS 0.009748f
C528 B.n211 VSUBS 0.009748f
C529 B.n212 VSUBS 0.009748f
C530 B.n213 VSUBS 0.009748f
C531 B.n214 VSUBS 0.009748f
C532 B.n215 VSUBS 0.009748f
C533 B.n216 VSUBS 0.009748f
C534 B.n217 VSUBS 0.009748f
C535 B.n218 VSUBS 0.009748f
C536 B.n219 VSUBS 0.009748f
C537 B.n220 VSUBS 0.009748f
C538 B.n221 VSUBS 0.009748f
C539 B.n222 VSUBS 0.009748f
C540 B.n223 VSUBS 0.009748f
C541 B.n224 VSUBS 0.009748f
C542 B.n225 VSUBS 0.009748f
C543 B.n226 VSUBS 0.009748f
C544 B.n227 VSUBS 0.009748f
C545 B.n228 VSUBS 0.009748f
C546 B.n229 VSUBS 0.009748f
C547 B.n230 VSUBS 0.009748f
C548 B.n231 VSUBS 0.009748f
C549 B.n232 VSUBS 0.009748f
C550 B.n233 VSUBS 0.009748f
C551 B.n234 VSUBS 0.009748f
C552 B.n235 VSUBS 0.009748f
C553 B.n236 VSUBS 0.009748f
C554 B.n237 VSUBS 0.009748f
C555 B.n238 VSUBS 0.009748f
C556 B.n239 VSUBS 0.009748f
C557 B.n240 VSUBS 0.009748f
C558 B.n241 VSUBS 0.009748f
C559 B.n242 VSUBS 0.009748f
C560 B.n243 VSUBS 0.009748f
C561 B.n244 VSUBS 0.009748f
C562 B.n245 VSUBS 0.009748f
C563 B.n246 VSUBS 0.009748f
C564 B.n247 VSUBS 0.009748f
C565 B.n248 VSUBS 0.009748f
C566 B.n249 VSUBS 0.009748f
C567 B.n250 VSUBS 0.009748f
C568 B.n251 VSUBS 0.009748f
C569 B.n252 VSUBS 0.009748f
C570 B.n253 VSUBS 0.009748f
C571 B.n254 VSUBS 0.009748f
C572 B.n255 VSUBS 0.009748f
C573 B.n256 VSUBS 0.009748f
C574 B.n257 VSUBS 0.009748f
C575 B.n258 VSUBS 0.009748f
C576 B.n259 VSUBS 0.009748f
C577 B.n260 VSUBS 0.009748f
C578 B.n261 VSUBS 0.009748f
C579 B.n262 VSUBS 0.009748f
C580 B.n263 VSUBS 0.009748f
C581 B.n264 VSUBS 0.009748f
C582 B.n265 VSUBS 0.009748f
C583 B.n266 VSUBS 0.009748f
C584 B.n267 VSUBS 0.009748f
C585 B.n268 VSUBS 0.009748f
C586 B.n269 VSUBS 0.009748f
C587 B.n270 VSUBS 0.009748f
C588 B.n271 VSUBS 0.009748f
C589 B.n272 VSUBS 0.009748f
C590 B.n273 VSUBS 0.009748f
C591 B.n274 VSUBS 0.009748f
C592 B.n275 VSUBS 0.009748f
C593 B.n276 VSUBS 0.009748f
C594 B.n277 VSUBS 0.009748f
C595 B.n278 VSUBS 0.009748f
C596 B.n279 VSUBS 0.009748f
C597 B.n280 VSUBS 0.009748f
C598 B.n281 VSUBS 0.009748f
C599 B.n282 VSUBS 0.009748f
C600 B.n283 VSUBS 0.009748f
C601 B.n284 VSUBS 0.009748f
C602 B.n285 VSUBS 0.009748f
C603 B.n286 VSUBS 0.009748f
C604 B.n287 VSUBS 0.009748f
C605 B.n288 VSUBS 0.009748f
C606 B.n289 VSUBS 0.009748f
C607 B.n290 VSUBS 0.009748f
C608 B.n291 VSUBS 0.009748f
C609 B.n292 VSUBS 0.009748f
C610 B.n293 VSUBS 0.009748f
C611 B.n294 VSUBS 0.009748f
C612 B.n295 VSUBS 0.009748f
C613 B.n296 VSUBS 0.009748f
C614 B.n297 VSUBS 0.009748f
C615 B.n298 VSUBS 0.009748f
C616 B.n299 VSUBS 0.009748f
C617 B.n300 VSUBS 0.009748f
C618 B.n301 VSUBS 0.009748f
C619 B.n302 VSUBS 0.009748f
C620 B.n303 VSUBS 0.009748f
C621 B.n304 VSUBS 0.009748f
C622 B.n305 VSUBS 0.009748f
C623 B.n306 VSUBS 0.009748f
C624 B.n307 VSUBS 0.009748f
C625 B.n308 VSUBS 0.009748f
C626 B.n309 VSUBS 0.009748f
C627 B.n310 VSUBS 0.009748f
C628 B.n311 VSUBS 0.023494f
C629 B.n312 VSUBS 0.023494f
C630 B.n313 VSUBS 0.0241f
C631 B.n314 VSUBS 0.009748f
C632 B.n315 VSUBS 0.009748f
C633 B.n316 VSUBS 0.009748f
C634 B.n317 VSUBS 0.009748f
C635 B.n318 VSUBS 0.009748f
C636 B.n319 VSUBS 0.009748f
C637 B.n320 VSUBS 0.009748f
C638 B.n321 VSUBS 0.009748f
C639 B.n322 VSUBS 0.009748f
C640 B.n323 VSUBS 0.009748f
C641 B.n324 VSUBS 0.009748f
C642 B.n325 VSUBS 0.009748f
C643 B.n326 VSUBS 0.009748f
C644 B.n327 VSUBS 0.009748f
C645 B.n328 VSUBS 0.009748f
C646 B.n329 VSUBS 0.009748f
C647 B.n330 VSUBS 0.009748f
C648 B.n331 VSUBS 0.009748f
C649 B.n332 VSUBS 0.009748f
C650 B.n333 VSUBS 0.009748f
C651 B.n334 VSUBS 0.009748f
C652 B.n335 VSUBS 0.009748f
C653 B.n336 VSUBS 0.009748f
C654 B.n337 VSUBS 0.009748f
C655 B.n338 VSUBS 0.009748f
C656 B.n339 VSUBS 0.009748f
C657 B.n340 VSUBS 0.009748f
C658 B.n341 VSUBS 0.009748f
C659 B.n342 VSUBS 0.009748f
C660 B.n343 VSUBS 0.009748f
C661 B.n344 VSUBS 0.009748f
C662 B.n345 VSUBS 0.009748f
C663 B.n346 VSUBS 0.009748f
C664 B.n347 VSUBS 0.009748f
C665 B.n348 VSUBS 0.009748f
C666 B.n349 VSUBS 0.009748f
C667 B.n350 VSUBS 0.009748f
C668 B.n351 VSUBS 0.009748f
C669 B.n352 VSUBS 0.009748f
C670 B.n353 VSUBS 0.009748f
C671 B.n354 VSUBS 0.009748f
C672 B.n355 VSUBS 0.009748f
C673 B.n356 VSUBS 0.009748f
C674 B.n357 VSUBS 0.009748f
C675 B.n358 VSUBS 0.009748f
C676 B.n359 VSUBS 0.009748f
C677 B.n360 VSUBS 0.009748f
C678 B.n361 VSUBS 0.009748f
C679 B.n362 VSUBS 0.009748f
C680 B.n363 VSUBS 0.009748f
C681 B.n364 VSUBS 0.009748f
C682 B.n365 VSUBS 0.009748f
C683 B.n366 VSUBS 0.009175f
C684 B.n367 VSUBS 0.022586f
C685 B.n368 VSUBS 0.005448f
C686 B.n369 VSUBS 0.009748f
C687 B.n370 VSUBS 0.009748f
C688 B.n371 VSUBS 0.009748f
C689 B.n372 VSUBS 0.009748f
C690 B.n373 VSUBS 0.009748f
C691 B.n374 VSUBS 0.009748f
C692 B.n375 VSUBS 0.009748f
C693 B.n376 VSUBS 0.009748f
C694 B.n377 VSUBS 0.009748f
C695 B.n378 VSUBS 0.009748f
C696 B.n379 VSUBS 0.009748f
C697 B.n380 VSUBS 0.009748f
C698 B.n381 VSUBS 0.005448f
C699 B.n382 VSUBS 0.009748f
C700 B.n383 VSUBS 0.009748f
C701 B.n384 VSUBS 0.009175f
C702 B.n385 VSUBS 0.009748f
C703 B.n386 VSUBS 0.009748f
C704 B.n387 VSUBS 0.009748f
C705 B.n388 VSUBS 0.009748f
C706 B.n389 VSUBS 0.009748f
C707 B.n390 VSUBS 0.009748f
C708 B.n391 VSUBS 0.009748f
C709 B.n392 VSUBS 0.009748f
C710 B.n393 VSUBS 0.009748f
C711 B.n394 VSUBS 0.009748f
C712 B.n395 VSUBS 0.009748f
C713 B.n396 VSUBS 0.009748f
C714 B.n397 VSUBS 0.009748f
C715 B.n398 VSUBS 0.009748f
C716 B.n399 VSUBS 0.009748f
C717 B.n400 VSUBS 0.009748f
C718 B.n401 VSUBS 0.009748f
C719 B.n402 VSUBS 0.009748f
C720 B.n403 VSUBS 0.009748f
C721 B.n404 VSUBS 0.009748f
C722 B.n405 VSUBS 0.009748f
C723 B.n406 VSUBS 0.009748f
C724 B.n407 VSUBS 0.009748f
C725 B.n408 VSUBS 0.009748f
C726 B.n409 VSUBS 0.009748f
C727 B.n410 VSUBS 0.009748f
C728 B.n411 VSUBS 0.009748f
C729 B.n412 VSUBS 0.009748f
C730 B.n413 VSUBS 0.009748f
C731 B.n414 VSUBS 0.009748f
C732 B.n415 VSUBS 0.009748f
C733 B.n416 VSUBS 0.009748f
C734 B.n417 VSUBS 0.009748f
C735 B.n418 VSUBS 0.009748f
C736 B.n419 VSUBS 0.009748f
C737 B.n420 VSUBS 0.009748f
C738 B.n421 VSUBS 0.009748f
C739 B.n422 VSUBS 0.009748f
C740 B.n423 VSUBS 0.009748f
C741 B.n424 VSUBS 0.009748f
C742 B.n425 VSUBS 0.009748f
C743 B.n426 VSUBS 0.009748f
C744 B.n427 VSUBS 0.009748f
C745 B.n428 VSUBS 0.009748f
C746 B.n429 VSUBS 0.009748f
C747 B.n430 VSUBS 0.009748f
C748 B.n431 VSUBS 0.009748f
C749 B.n432 VSUBS 0.009748f
C750 B.n433 VSUBS 0.009748f
C751 B.n434 VSUBS 0.009748f
C752 B.n435 VSUBS 0.009748f
C753 B.n436 VSUBS 0.0241f
C754 B.n437 VSUBS 0.023494f
C755 B.n438 VSUBS 0.023494f
C756 B.n439 VSUBS 0.009748f
C757 B.n440 VSUBS 0.009748f
C758 B.n441 VSUBS 0.009748f
C759 B.n442 VSUBS 0.009748f
C760 B.n443 VSUBS 0.009748f
C761 B.n444 VSUBS 0.009748f
C762 B.n445 VSUBS 0.009748f
C763 B.n446 VSUBS 0.009748f
C764 B.n447 VSUBS 0.009748f
C765 B.n448 VSUBS 0.009748f
C766 B.n449 VSUBS 0.009748f
C767 B.n450 VSUBS 0.009748f
C768 B.n451 VSUBS 0.009748f
C769 B.n452 VSUBS 0.009748f
C770 B.n453 VSUBS 0.009748f
C771 B.n454 VSUBS 0.009748f
C772 B.n455 VSUBS 0.009748f
C773 B.n456 VSUBS 0.009748f
C774 B.n457 VSUBS 0.009748f
C775 B.n458 VSUBS 0.009748f
C776 B.n459 VSUBS 0.009748f
C777 B.n460 VSUBS 0.009748f
C778 B.n461 VSUBS 0.009748f
C779 B.n462 VSUBS 0.009748f
C780 B.n463 VSUBS 0.009748f
C781 B.n464 VSUBS 0.009748f
C782 B.n465 VSUBS 0.009748f
C783 B.n466 VSUBS 0.009748f
C784 B.n467 VSUBS 0.009748f
C785 B.n468 VSUBS 0.009748f
C786 B.n469 VSUBS 0.009748f
C787 B.n470 VSUBS 0.009748f
C788 B.n471 VSUBS 0.009748f
C789 B.n472 VSUBS 0.009748f
C790 B.n473 VSUBS 0.009748f
C791 B.n474 VSUBS 0.009748f
C792 B.n475 VSUBS 0.009748f
C793 B.n476 VSUBS 0.009748f
C794 B.n477 VSUBS 0.009748f
C795 B.n478 VSUBS 0.009748f
C796 B.n479 VSUBS 0.009748f
C797 B.n480 VSUBS 0.009748f
C798 B.n481 VSUBS 0.009748f
C799 B.n482 VSUBS 0.009748f
C800 B.n483 VSUBS 0.009748f
C801 B.n484 VSUBS 0.009748f
C802 B.n485 VSUBS 0.009748f
C803 B.n486 VSUBS 0.009748f
C804 B.n487 VSUBS 0.009748f
C805 B.n488 VSUBS 0.009748f
C806 B.n489 VSUBS 0.009748f
C807 B.n490 VSUBS 0.009748f
C808 B.n491 VSUBS 0.009748f
C809 B.n492 VSUBS 0.009748f
C810 B.n493 VSUBS 0.009748f
C811 B.n494 VSUBS 0.009748f
C812 B.n495 VSUBS 0.009748f
C813 B.n496 VSUBS 0.009748f
C814 B.n497 VSUBS 0.009748f
C815 B.n498 VSUBS 0.009748f
C816 B.n499 VSUBS 0.009748f
C817 B.n500 VSUBS 0.009748f
C818 B.n501 VSUBS 0.009748f
C819 B.n502 VSUBS 0.009748f
C820 B.n503 VSUBS 0.009748f
C821 B.n504 VSUBS 0.009748f
C822 B.n505 VSUBS 0.009748f
C823 B.n506 VSUBS 0.009748f
C824 B.n507 VSUBS 0.009748f
C825 B.n508 VSUBS 0.009748f
C826 B.n509 VSUBS 0.009748f
C827 B.n510 VSUBS 0.009748f
C828 B.n511 VSUBS 0.009748f
C829 B.n512 VSUBS 0.009748f
C830 B.n513 VSUBS 0.009748f
C831 B.n514 VSUBS 0.009748f
C832 B.n515 VSUBS 0.009748f
C833 B.n516 VSUBS 0.009748f
C834 B.n517 VSUBS 0.009748f
C835 B.n518 VSUBS 0.009748f
C836 B.n519 VSUBS 0.009748f
C837 B.n520 VSUBS 0.009748f
C838 B.n521 VSUBS 0.009748f
C839 B.n522 VSUBS 0.009748f
C840 B.n523 VSUBS 0.009748f
C841 B.n524 VSUBS 0.009748f
C842 B.n525 VSUBS 0.009748f
C843 B.n526 VSUBS 0.009748f
C844 B.n527 VSUBS 0.009748f
C845 B.n528 VSUBS 0.009748f
C846 B.n529 VSUBS 0.009748f
C847 B.n530 VSUBS 0.009748f
C848 B.n531 VSUBS 0.009748f
C849 B.n532 VSUBS 0.009748f
C850 B.n533 VSUBS 0.009748f
C851 B.n534 VSUBS 0.009748f
C852 B.n535 VSUBS 0.009748f
C853 B.n536 VSUBS 0.009748f
C854 B.n537 VSUBS 0.009748f
C855 B.n538 VSUBS 0.009748f
C856 B.n539 VSUBS 0.009748f
C857 B.n540 VSUBS 0.009748f
C858 B.n541 VSUBS 0.009748f
C859 B.n542 VSUBS 0.009748f
C860 B.n543 VSUBS 0.009748f
C861 B.n544 VSUBS 0.009748f
C862 B.n545 VSUBS 0.009748f
C863 B.n546 VSUBS 0.009748f
C864 B.n547 VSUBS 0.009748f
C865 B.n548 VSUBS 0.009748f
C866 B.n549 VSUBS 0.009748f
C867 B.n550 VSUBS 0.009748f
C868 B.n551 VSUBS 0.009748f
C869 B.n552 VSUBS 0.009748f
C870 B.n553 VSUBS 0.009748f
C871 B.n554 VSUBS 0.009748f
C872 B.n555 VSUBS 0.009748f
C873 B.n556 VSUBS 0.009748f
C874 B.n557 VSUBS 0.009748f
C875 B.n558 VSUBS 0.009748f
C876 B.n559 VSUBS 0.009748f
C877 B.n560 VSUBS 0.009748f
C878 B.n561 VSUBS 0.009748f
C879 B.n562 VSUBS 0.009748f
C880 B.n563 VSUBS 0.009748f
C881 B.n564 VSUBS 0.009748f
C882 B.n565 VSUBS 0.009748f
C883 B.n566 VSUBS 0.009748f
C884 B.n567 VSUBS 0.009748f
C885 B.n568 VSUBS 0.009748f
C886 B.n569 VSUBS 0.009748f
C887 B.n570 VSUBS 0.009748f
C888 B.n571 VSUBS 0.009748f
C889 B.n572 VSUBS 0.009748f
C890 B.n573 VSUBS 0.009748f
C891 B.n574 VSUBS 0.009748f
C892 B.n575 VSUBS 0.009748f
C893 B.n576 VSUBS 0.009748f
C894 B.n577 VSUBS 0.009748f
C895 B.n578 VSUBS 0.009748f
C896 B.n579 VSUBS 0.009748f
C897 B.n580 VSUBS 0.009748f
C898 B.n581 VSUBS 0.009748f
C899 B.n582 VSUBS 0.009748f
C900 B.n583 VSUBS 0.009748f
C901 B.n584 VSUBS 0.009748f
C902 B.n585 VSUBS 0.009748f
C903 B.n586 VSUBS 0.009748f
C904 B.n587 VSUBS 0.009748f
C905 B.n588 VSUBS 0.009748f
C906 B.n589 VSUBS 0.009748f
C907 B.n590 VSUBS 0.009748f
C908 B.n591 VSUBS 0.009748f
C909 B.n592 VSUBS 0.009748f
C910 B.n593 VSUBS 0.009748f
C911 B.n594 VSUBS 0.009748f
C912 B.n595 VSUBS 0.009748f
C913 B.n596 VSUBS 0.009748f
C914 B.n597 VSUBS 0.009748f
C915 B.n598 VSUBS 0.009748f
C916 B.n599 VSUBS 0.009748f
C917 B.n600 VSUBS 0.009748f
C918 B.n601 VSUBS 0.009748f
C919 B.n602 VSUBS 0.009748f
C920 B.n603 VSUBS 0.009748f
C921 B.n604 VSUBS 0.009748f
C922 B.n605 VSUBS 0.009748f
C923 B.n606 VSUBS 0.009748f
C924 B.n607 VSUBS 0.009748f
C925 B.n608 VSUBS 0.009748f
C926 B.n609 VSUBS 0.009748f
C927 B.n610 VSUBS 0.009748f
C928 B.n611 VSUBS 0.009748f
C929 B.n612 VSUBS 0.009748f
C930 B.n613 VSUBS 0.009748f
C931 B.n614 VSUBS 0.009748f
C932 B.n615 VSUBS 0.009748f
C933 B.n616 VSUBS 0.009748f
C934 B.n617 VSUBS 0.009748f
C935 B.n618 VSUBS 0.009748f
C936 B.n619 VSUBS 0.009748f
C937 B.n620 VSUBS 0.009748f
C938 B.n621 VSUBS 0.009748f
C939 B.n622 VSUBS 0.009748f
C940 B.n623 VSUBS 0.009748f
C941 B.n624 VSUBS 0.009748f
C942 B.n625 VSUBS 0.009748f
C943 B.n626 VSUBS 0.024575f
C944 B.n627 VSUBS 0.023494f
C945 B.n628 VSUBS 0.0241f
C946 B.n629 VSUBS 0.009748f
C947 B.n630 VSUBS 0.009748f
C948 B.n631 VSUBS 0.009748f
C949 B.n632 VSUBS 0.009748f
C950 B.n633 VSUBS 0.009748f
C951 B.n634 VSUBS 0.009748f
C952 B.n635 VSUBS 0.009748f
C953 B.n636 VSUBS 0.009748f
C954 B.n637 VSUBS 0.009748f
C955 B.n638 VSUBS 0.009748f
C956 B.n639 VSUBS 0.009748f
C957 B.n640 VSUBS 0.009748f
C958 B.n641 VSUBS 0.009748f
C959 B.n642 VSUBS 0.009748f
C960 B.n643 VSUBS 0.009748f
C961 B.n644 VSUBS 0.009748f
C962 B.n645 VSUBS 0.009748f
C963 B.n646 VSUBS 0.009748f
C964 B.n647 VSUBS 0.009748f
C965 B.n648 VSUBS 0.009748f
C966 B.n649 VSUBS 0.009748f
C967 B.n650 VSUBS 0.009748f
C968 B.n651 VSUBS 0.009748f
C969 B.n652 VSUBS 0.009748f
C970 B.n653 VSUBS 0.009748f
C971 B.n654 VSUBS 0.009748f
C972 B.n655 VSUBS 0.009748f
C973 B.n656 VSUBS 0.009748f
C974 B.n657 VSUBS 0.009748f
C975 B.n658 VSUBS 0.009748f
C976 B.n659 VSUBS 0.009748f
C977 B.n660 VSUBS 0.009748f
C978 B.n661 VSUBS 0.009748f
C979 B.n662 VSUBS 0.009748f
C980 B.n663 VSUBS 0.009748f
C981 B.n664 VSUBS 0.009748f
C982 B.n665 VSUBS 0.009748f
C983 B.n666 VSUBS 0.009748f
C984 B.n667 VSUBS 0.009748f
C985 B.n668 VSUBS 0.009748f
C986 B.n669 VSUBS 0.009748f
C987 B.n670 VSUBS 0.009748f
C988 B.n671 VSUBS 0.009748f
C989 B.n672 VSUBS 0.009748f
C990 B.n673 VSUBS 0.009748f
C991 B.n674 VSUBS 0.009748f
C992 B.n675 VSUBS 0.009748f
C993 B.n676 VSUBS 0.009748f
C994 B.n677 VSUBS 0.009748f
C995 B.n678 VSUBS 0.009748f
C996 B.n679 VSUBS 0.009748f
C997 B.n680 VSUBS 0.009175f
C998 B.n681 VSUBS 0.009748f
C999 B.n682 VSUBS 0.009748f
C1000 B.n683 VSUBS 0.009748f
C1001 B.n684 VSUBS 0.009748f
C1002 B.n685 VSUBS 0.009748f
C1003 B.n686 VSUBS 0.009748f
C1004 B.n687 VSUBS 0.009748f
C1005 B.n688 VSUBS 0.009748f
C1006 B.n689 VSUBS 0.009748f
C1007 B.n690 VSUBS 0.009748f
C1008 B.n691 VSUBS 0.009748f
C1009 B.n692 VSUBS 0.009748f
C1010 B.n693 VSUBS 0.009748f
C1011 B.n694 VSUBS 0.009748f
C1012 B.n695 VSUBS 0.009748f
C1013 B.n696 VSUBS 0.005448f
C1014 B.n697 VSUBS 0.022586f
C1015 B.n698 VSUBS 0.009175f
C1016 B.n699 VSUBS 0.009748f
C1017 B.n700 VSUBS 0.009748f
C1018 B.n701 VSUBS 0.009748f
C1019 B.n702 VSUBS 0.009748f
C1020 B.n703 VSUBS 0.009748f
C1021 B.n704 VSUBS 0.009748f
C1022 B.n705 VSUBS 0.009748f
C1023 B.n706 VSUBS 0.009748f
C1024 B.n707 VSUBS 0.009748f
C1025 B.n708 VSUBS 0.009748f
C1026 B.n709 VSUBS 0.009748f
C1027 B.n710 VSUBS 0.009748f
C1028 B.n711 VSUBS 0.009748f
C1029 B.n712 VSUBS 0.009748f
C1030 B.n713 VSUBS 0.009748f
C1031 B.n714 VSUBS 0.009748f
C1032 B.n715 VSUBS 0.009748f
C1033 B.n716 VSUBS 0.009748f
C1034 B.n717 VSUBS 0.009748f
C1035 B.n718 VSUBS 0.009748f
C1036 B.n719 VSUBS 0.009748f
C1037 B.n720 VSUBS 0.009748f
C1038 B.n721 VSUBS 0.009748f
C1039 B.n722 VSUBS 0.009748f
C1040 B.n723 VSUBS 0.009748f
C1041 B.n724 VSUBS 0.009748f
C1042 B.n725 VSUBS 0.009748f
C1043 B.n726 VSUBS 0.009748f
C1044 B.n727 VSUBS 0.009748f
C1045 B.n728 VSUBS 0.009748f
C1046 B.n729 VSUBS 0.009748f
C1047 B.n730 VSUBS 0.009748f
C1048 B.n731 VSUBS 0.009748f
C1049 B.n732 VSUBS 0.009748f
C1050 B.n733 VSUBS 0.009748f
C1051 B.n734 VSUBS 0.009748f
C1052 B.n735 VSUBS 0.009748f
C1053 B.n736 VSUBS 0.009748f
C1054 B.n737 VSUBS 0.009748f
C1055 B.n738 VSUBS 0.009748f
C1056 B.n739 VSUBS 0.009748f
C1057 B.n740 VSUBS 0.009748f
C1058 B.n741 VSUBS 0.009748f
C1059 B.n742 VSUBS 0.009748f
C1060 B.n743 VSUBS 0.009748f
C1061 B.n744 VSUBS 0.009748f
C1062 B.n745 VSUBS 0.009748f
C1063 B.n746 VSUBS 0.009748f
C1064 B.n747 VSUBS 0.009748f
C1065 B.n748 VSUBS 0.009748f
C1066 B.n749 VSUBS 0.009748f
C1067 B.n750 VSUBS 0.0241f
C1068 B.n751 VSUBS 0.0241f
C1069 B.n752 VSUBS 0.023494f
C1070 B.n753 VSUBS 0.009748f
C1071 B.n754 VSUBS 0.009748f
C1072 B.n755 VSUBS 0.009748f
C1073 B.n756 VSUBS 0.009748f
C1074 B.n757 VSUBS 0.009748f
C1075 B.n758 VSUBS 0.009748f
C1076 B.n759 VSUBS 0.009748f
C1077 B.n760 VSUBS 0.009748f
C1078 B.n761 VSUBS 0.009748f
C1079 B.n762 VSUBS 0.009748f
C1080 B.n763 VSUBS 0.009748f
C1081 B.n764 VSUBS 0.009748f
C1082 B.n765 VSUBS 0.009748f
C1083 B.n766 VSUBS 0.009748f
C1084 B.n767 VSUBS 0.009748f
C1085 B.n768 VSUBS 0.009748f
C1086 B.n769 VSUBS 0.009748f
C1087 B.n770 VSUBS 0.009748f
C1088 B.n771 VSUBS 0.009748f
C1089 B.n772 VSUBS 0.009748f
C1090 B.n773 VSUBS 0.009748f
C1091 B.n774 VSUBS 0.009748f
C1092 B.n775 VSUBS 0.009748f
C1093 B.n776 VSUBS 0.009748f
C1094 B.n777 VSUBS 0.009748f
C1095 B.n778 VSUBS 0.009748f
C1096 B.n779 VSUBS 0.009748f
C1097 B.n780 VSUBS 0.009748f
C1098 B.n781 VSUBS 0.009748f
C1099 B.n782 VSUBS 0.009748f
C1100 B.n783 VSUBS 0.009748f
C1101 B.n784 VSUBS 0.009748f
C1102 B.n785 VSUBS 0.009748f
C1103 B.n786 VSUBS 0.009748f
C1104 B.n787 VSUBS 0.009748f
C1105 B.n788 VSUBS 0.009748f
C1106 B.n789 VSUBS 0.009748f
C1107 B.n790 VSUBS 0.009748f
C1108 B.n791 VSUBS 0.009748f
C1109 B.n792 VSUBS 0.009748f
C1110 B.n793 VSUBS 0.009748f
C1111 B.n794 VSUBS 0.009748f
C1112 B.n795 VSUBS 0.009748f
C1113 B.n796 VSUBS 0.009748f
C1114 B.n797 VSUBS 0.009748f
C1115 B.n798 VSUBS 0.009748f
C1116 B.n799 VSUBS 0.009748f
C1117 B.n800 VSUBS 0.009748f
C1118 B.n801 VSUBS 0.009748f
C1119 B.n802 VSUBS 0.009748f
C1120 B.n803 VSUBS 0.009748f
C1121 B.n804 VSUBS 0.009748f
C1122 B.n805 VSUBS 0.009748f
C1123 B.n806 VSUBS 0.009748f
C1124 B.n807 VSUBS 0.009748f
C1125 B.n808 VSUBS 0.009748f
C1126 B.n809 VSUBS 0.009748f
C1127 B.n810 VSUBS 0.009748f
C1128 B.n811 VSUBS 0.009748f
C1129 B.n812 VSUBS 0.009748f
C1130 B.n813 VSUBS 0.009748f
C1131 B.n814 VSUBS 0.009748f
C1132 B.n815 VSUBS 0.009748f
C1133 B.n816 VSUBS 0.009748f
C1134 B.n817 VSUBS 0.009748f
C1135 B.n818 VSUBS 0.009748f
C1136 B.n819 VSUBS 0.009748f
C1137 B.n820 VSUBS 0.009748f
C1138 B.n821 VSUBS 0.009748f
C1139 B.n822 VSUBS 0.009748f
C1140 B.n823 VSUBS 0.009748f
C1141 B.n824 VSUBS 0.009748f
C1142 B.n825 VSUBS 0.009748f
C1143 B.n826 VSUBS 0.009748f
C1144 B.n827 VSUBS 0.009748f
C1145 B.n828 VSUBS 0.009748f
C1146 B.n829 VSUBS 0.009748f
C1147 B.n830 VSUBS 0.009748f
C1148 B.n831 VSUBS 0.009748f
C1149 B.n832 VSUBS 0.009748f
C1150 B.n833 VSUBS 0.009748f
C1151 B.n834 VSUBS 0.009748f
C1152 B.n835 VSUBS 0.009748f
C1153 B.n836 VSUBS 0.009748f
C1154 B.n837 VSUBS 0.009748f
C1155 B.n838 VSUBS 0.009748f
C1156 B.n839 VSUBS 0.009748f
C1157 B.n840 VSUBS 0.009748f
C1158 B.n841 VSUBS 0.009748f
C1159 B.n842 VSUBS 0.009748f
C1160 B.n843 VSUBS 0.009748f
C1161 B.n844 VSUBS 0.009748f
C1162 B.n845 VSUBS 0.009748f
C1163 B.n846 VSUBS 0.009748f
C1164 B.n847 VSUBS 0.022073f
.ends

