* NGSPICE file created from diff_pair_sample_1355.ext - technology: sky130A

.subckt diff_pair_sample_1355 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X1 VDD1.t9 VP.t0 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X2 VDD1.t8 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=1.15
X3 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X4 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=1.15
X5 VTAIL.t0 VP.t3 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X6 VDD2.t0 VN.t1 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=1.15
X7 VDD2.t7 VN.t2 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=1.15
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=1.15
X9 VDD2.t4 VN.t3 VTAIL.t15 B.t23 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X10 VDD2.t1 VN.t4 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=1.15
X12 VDD2.t9 VN.t5 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=1.15
X13 VTAIL.t12 VN.t6 VDD2.t5 B.t22 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X14 VTAIL.t8 VP.t4 VDD1.t5 B.t22 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X15 VTAIL.t11 VN.t7 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X16 VDD2.t3 VN.t8 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=1.15
X17 VDD1.t4 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=1.15
X18 VTAIL.t5 VP.t6 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0 ps=0 w=5.64 l=1.15
X20 VTAIL.t9 VN.t9 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X21 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=0.9306 ps=5.97 w=5.64 l=1.15
X22 VDD1.t1 VP.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9306 pd=5.97 as=2.1996 ps=12.06 w=5.64 l=1.15
X23 VDD1.t0 VP.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1996 pd=12.06 as=0.9306 ps=5.97 w=5.64 l=1.15
R0 VN.n4 VN.t2 175.499
R1 VN.n23 VN.t8 175.499
R2 VN.n35 VN.n19 161.3
R3 VN.n34 VN.n33 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n21 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n22 161.3
R8 VN.n26 VN.n25 161.3
R9 VN.n16 VN.n0 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n11 VN.n2 161.3
R13 VN.n10 VN.n9 161.3
R14 VN.n8 VN.n3 161.3
R15 VN.n7 VN.n6 161.3
R16 VN.n17 VN.t5 152.355
R17 VN.n36 VN.t1 152.355
R18 VN.n10 VN.t4 118.195
R19 VN.n5 VN.t6 118.195
R20 VN.n1 VN.t7 118.195
R21 VN.n29 VN.t3 118.195
R22 VN.n24 VN.t0 118.195
R23 VN.n20 VN.t9 118.195
R24 VN.n37 VN.n36 80.6037
R25 VN.n18 VN.n17 80.6037
R26 VN.n12 VN.n11 56.5617
R27 VN.n31 VN.n30 56.5617
R28 VN.n6 VN.n3 56.5617
R29 VN.n25 VN.n22 56.5617
R30 VN.n17 VN.n16 50.9056
R31 VN.n36 VN.n35 50.9056
R32 VN VN.n37 40.9233
R33 VN.n5 VN.n4 33.7965
R34 VN.n24 VN.n23 33.7965
R35 VN.n26 VN.n23 28.0737
R36 VN.n7 VN.n4 28.0737
R37 VN.n10 VN.n3 24.5923
R38 VN.n11 VN.n10 24.5923
R39 VN.n16 VN.n15 24.5923
R40 VN.n30 VN.n29 24.5923
R41 VN.n29 VN.n22 24.5923
R42 VN.n35 VN.n34 24.5923
R43 VN.n6 VN.n5 23.6087
R44 VN.n12 VN.n1 23.6087
R45 VN.n25 VN.n24 23.6087
R46 VN.n31 VN.n20 23.6087
R47 VN.n15 VN.n1 0.984173
R48 VN.n34 VN.n20 0.984173
R49 VN.n37 VN.n19 0.285035
R50 VN.n18 VN.n0 0.285035
R51 VN.n33 VN.n19 0.189894
R52 VN.n33 VN.n32 0.189894
R53 VN.n32 VN.n21 0.189894
R54 VN.n28 VN.n21 0.189894
R55 VN.n28 VN.n27 0.189894
R56 VN.n27 VN.n26 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n9 VN.n8 0.189894
R59 VN.n9 VN.n2 0.189894
R60 VN.n13 VN.n2 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n0 0.189894
R63 VN VN.n18 0.146778
R64 VDD2.n1 VDD2.t7 72.6563
R65 VDD2.n4 VDD2.t0 71.3807
R66 VDD2.n3 VDD2.n2 68.7714
R67 VDD2 VDD2.n7 68.7686
R68 VDD2.n6 VDD2.n5 67.87
R69 VDD2.n1 VDD2.n0 67.8698
R70 VDD2.n4 VDD2.n3 34.6377
R71 VDD2.n7 VDD2.t6 3.51114
R72 VDD2.n7 VDD2.t3 3.51114
R73 VDD2.n5 VDD2.t8 3.51114
R74 VDD2.n5 VDD2.t4 3.51114
R75 VDD2.n2 VDD2.t2 3.51114
R76 VDD2.n2 VDD2.t9 3.51114
R77 VDD2.n0 VDD2.t5 3.51114
R78 VDD2.n0 VDD2.t1 3.51114
R79 VDD2.n6 VDD2.n4 1.27636
R80 VDD2 VDD2.n6 0.377655
R81 VDD2.n3 VDD2.n1 0.26412
R82 VTAIL.n11 VTAIL.t10 54.7019
R83 VTAIL.n17 VTAIL.t13 54.7017
R84 VTAIL.n2 VTAIL.t1 54.7017
R85 VTAIL.n16 VTAIL.t6 54.7017
R86 VTAIL.n15 VTAIL.n14 51.1912
R87 VTAIL.n13 VTAIL.n12 51.1912
R88 VTAIL.n10 VTAIL.n9 51.1912
R89 VTAIL.n8 VTAIL.n7 51.1912
R90 VTAIL.n19 VTAIL.n18 51.191
R91 VTAIL.n1 VTAIL.n0 51.191
R92 VTAIL.n4 VTAIL.n3 51.191
R93 VTAIL.n6 VTAIL.n5 51.191
R94 VTAIL.n8 VTAIL.n6 19.7807
R95 VTAIL.n17 VTAIL.n16 18.5048
R96 VTAIL.n18 VTAIL.t14 3.51114
R97 VTAIL.n18 VTAIL.t11 3.51114
R98 VTAIL.n0 VTAIL.t16 3.51114
R99 VTAIL.n0 VTAIL.t12 3.51114
R100 VTAIL.n3 VTAIL.t19 3.51114
R101 VTAIL.n3 VTAIL.t2 3.51114
R102 VTAIL.n5 VTAIL.t4 3.51114
R103 VTAIL.n5 VTAIL.t5 3.51114
R104 VTAIL.n14 VTAIL.t7 3.51114
R105 VTAIL.n14 VTAIL.t0 3.51114
R106 VTAIL.n12 VTAIL.t3 3.51114
R107 VTAIL.n12 VTAIL.t8 3.51114
R108 VTAIL.n9 VTAIL.t15 3.51114
R109 VTAIL.n9 VTAIL.t18 3.51114
R110 VTAIL.n7 VTAIL.t17 3.51114
R111 VTAIL.n7 VTAIL.t9 3.51114
R112 VTAIL.n10 VTAIL.n8 1.27636
R113 VTAIL.n11 VTAIL.n10 1.27636
R114 VTAIL.n15 VTAIL.n13 1.27636
R115 VTAIL.n16 VTAIL.n15 1.27636
R116 VTAIL.n6 VTAIL.n4 1.27636
R117 VTAIL.n4 VTAIL.n2 1.27636
R118 VTAIL.n19 VTAIL.n17 1.27636
R119 VTAIL.n13 VTAIL.n11 1.10826
R120 VTAIL.n2 VTAIL.n1 1.10826
R121 VTAIL VTAIL.n1 1.01559
R122 VTAIL VTAIL.n19 0.261276
R123 B.n452 B.n451 585
R124 B.n452 B.n64 585
R125 B.n455 B.n454 585
R126 B.n456 B.n96 585
R127 B.n458 B.n457 585
R128 B.n460 B.n95 585
R129 B.n463 B.n462 585
R130 B.n464 B.n94 585
R131 B.n466 B.n465 585
R132 B.n468 B.n93 585
R133 B.n471 B.n470 585
R134 B.n472 B.n92 585
R135 B.n474 B.n473 585
R136 B.n476 B.n91 585
R137 B.n479 B.n478 585
R138 B.n480 B.n90 585
R139 B.n482 B.n481 585
R140 B.n484 B.n89 585
R141 B.n487 B.n486 585
R142 B.n488 B.n88 585
R143 B.n490 B.n489 585
R144 B.n492 B.n87 585
R145 B.n495 B.n494 585
R146 B.n496 B.n84 585
R147 B.n499 B.n498 585
R148 B.n501 B.n83 585
R149 B.n504 B.n503 585
R150 B.n505 B.n82 585
R151 B.n507 B.n506 585
R152 B.n509 B.n81 585
R153 B.n512 B.n511 585
R154 B.n513 B.n77 585
R155 B.n515 B.n514 585
R156 B.n517 B.n76 585
R157 B.n520 B.n519 585
R158 B.n521 B.n75 585
R159 B.n523 B.n522 585
R160 B.n525 B.n74 585
R161 B.n528 B.n527 585
R162 B.n529 B.n73 585
R163 B.n531 B.n530 585
R164 B.n533 B.n72 585
R165 B.n536 B.n535 585
R166 B.n537 B.n71 585
R167 B.n539 B.n538 585
R168 B.n541 B.n70 585
R169 B.n544 B.n543 585
R170 B.n545 B.n69 585
R171 B.n547 B.n546 585
R172 B.n549 B.n68 585
R173 B.n552 B.n551 585
R174 B.n553 B.n67 585
R175 B.n555 B.n554 585
R176 B.n557 B.n66 585
R177 B.n560 B.n559 585
R178 B.n561 B.n65 585
R179 B.n450 B.n63 585
R180 B.n564 B.n63 585
R181 B.n449 B.n62 585
R182 B.n565 B.n62 585
R183 B.n448 B.n61 585
R184 B.n566 B.n61 585
R185 B.n447 B.n446 585
R186 B.n446 B.n57 585
R187 B.n445 B.n56 585
R188 B.n572 B.n56 585
R189 B.n444 B.n55 585
R190 B.n573 B.n55 585
R191 B.n443 B.n54 585
R192 B.n574 B.n54 585
R193 B.n442 B.n441 585
R194 B.n441 B.n50 585
R195 B.n440 B.n49 585
R196 B.n580 B.n49 585
R197 B.n439 B.n48 585
R198 B.n581 B.n48 585
R199 B.n438 B.n47 585
R200 B.n582 B.n47 585
R201 B.n437 B.n436 585
R202 B.n436 B.n43 585
R203 B.n435 B.n42 585
R204 B.n588 B.n42 585
R205 B.n434 B.n41 585
R206 B.n589 B.n41 585
R207 B.n433 B.n40 585
R208 B.n590 B.n40 585
R209 B.n432 B.n431 585
R210 B.n431 B.n36 585
R211 B.n430 B.n35 585
R212 B.n596 B.n35 585
R213 B.n429 B.n34 585
R214 B.n597 B.n34 585
R215 B.n428 B.n33 585
R216 B.n598 B.n33 585
R217 B.n427 B.n426 585
R218 B.n426 B.n29 585
R219 B.n425 B.n28 585
R220 B.n604 B.n28 585
R221 B.n424 B.n27 585
R222 B.n605 B.n27 585
R223 B.n423 B.n26 585
R224 B.n606 B.n26 585
R225 B.n422 B.n421 585
R226 B.n421 B.n22 585
R227 B.n420 B.n21 585
R228 B.n612 B.n21 585
R229 B.n419 B.n20 585
R230 B.n613 B.n20 585
R231 B.n418 B.n19 585
R232 B.n614 B.n19 585
R233 B.n417 B.n416 585
R234 B.n416 B.n15 585
R235 B.n415 B.n14 585
R236 B.n620 B.n14 585
R237 B.n414 B.n13 585
R238 B.n621 B.n13 585
R239 B.n413 B.n12 585
R240 B.n622 B.n12 585
R241 B.n412 B.n411 585
R242 B.n411 B.n8 585
R243 B.n410 B.n7 585
R244 B.n628 B.n7 585
R245 B.n409 B.n6 585
R246 B.n629 B.n6 585
R247 B.n408 B.n5 585
R248 B.n630 B.n5 585
R249 B.n407 B.n406 585
R250 B.n406 B.n4 585
R251 B.n405 B.n97 585
R252 B.n405 B.n404 585
R253 B.n395 B.n98 585
R254 B.n99 B.n98 585
R255 B.n397 B.n396 585
R256 B.n398 B.n397 585
R257 B.n394 B.n104 585
R258 B.n104 B.n103 585
R259 B.n393 B.n392 585
R260 B.n392 B.n391 585
R261 B.n106 B.n105 585
R262 B.n107 B.n106 585
R263 B.n384 B.n383 585
R264 B.n385 B.n384 585
R265 B.n382 B.n111 585
R266 B.n115 B.n111 585
R267 B.n381 B.n380 585
R268 B.n380 B.n379 585
R269 B.n113 B.n112 585
R270 B.n114 B.n113 585
R271 B.n372 B.n371 585
R272 B.n373 B.n372 585
R273 B.n370 B.n119 585
R274 B.n123 B.n119 585
R275 B.n369 B.n368 585
R276 B.n368 B.n367 585
R277 B.n121 B.n120 585
R278 B.n122 B.n121 585
R279 B.n360 B.n359 585
R280 B.n361 B.n360 585
R281 B.n358 B.n127 585
R282 B.n131 B.n127 585
R283 B.n357 B.n356 585
R284 B.n356 B.n355 585
R285 B.n129 B.n128 585
R286 B.n130 B.n129 585
R287 B.n348 B.n347 585
R288 B.n349 B.n348 585
R289 B.n346 B.n136 585
R290 B.n136 B.n135 585
R291 B.n345 B.n344 585
R292 B.n344 B.n343 585
R293 B.n138 B.n137 585
R294 B.n139 B.n138 585
R295 B.n336 B.n335 585
R296 B.n337 B.n336 585
R297 B.n334 B.n144 585
R298 B.n144 B.n143 585
R299 B.n333 B.n332 585
R300 B.n332 B.n331 585
R301 B.n146 B.n145 585
R302 B.n147 B.n146 585
R303 B.n324 B.n323 585
R304 B.n325 B.n324 585
R305 B.n322 B.n151 585
R306 B.n155 B.n151 585
R307 B.n321 B.n320 585
R308 B.n320 B.n319 585
R309 B.n153 B.n152 585
R310 B.n154 B.n153 585
R311 B.n312 B.n311 585
R312 B.n313 B.n312 585
R313 B.n310 B.n160 585
R314 B.n160 B.n159 585
R315 B.n309 B.n308 585
R316 B.n308 B.n307 585
R317 B.n304 B.n164 585
R318 B.n303 B.n302 585
R319 B.n300 B.n165 585
R320 B.n300 B.n163 585
R321 B.n299 B.n298 585
R322 B.n297 B.n296 585
R323 B.n295 B.n167 585
R324 B.n293 B.n292 585
R325 B.n291 B.n168 585
R326 B.n290 B.n289 585
R327 B.n287 B.n169 585
R328 B.n285 B.n284 585
R329 B.n283 B.n170 585
R330 B.n282 B.n281 585
R331 B.n279 B.n171 585
R332 B.n277 B.n276 585
R333 B.n275 B.n172 585
R334 B.n274 B.n273 585
R335 B.n271 B.n173 585
R336 B.n269 B.n268 585
R337 B.n267 B.n174 585
R338 B.n266 B.n265 585
R339 B.n263 B.n175 585
R340 B.n261 B.n260 585
R341 B.n258 B.n176 585
R342 B.n257 B.n256 585
R343 B.n254 B.n179 585
R344 B.n252 B.n251 585
R345 B.n250 B.n180 585
R346 B.n249 B.n248 585
R347 B.n246 B.n181 585
R348 B.n244 B.n243 585
R349 B.n242 B.n182 585
R350 B.n240 B.n239 585
R351 B.n237 B.n185 585
R352 B.n235 B.n234 585
R353 B.n233 B.n186 585
R354 B.n232 B.n231 585
R355 B.n229 B.n187 585
R356 B.n227 B.n226 585
R357 B.n225 B.n188 585
R358 B.n224 B.n223 585
R359 B.n221 B.n189 585
R360 B.n219 B.n218 585
R361 B.n217 B.n190 585
R362 B.n216 B.n215 585
R363 B.n213 B.n191 585
R364 B.n211 B.n210 585
R365 B.n209 B.n192 585
R366 B.n208 B.n207 585
R367 B.n205 B.n193 585
R368 B.n203 B.n202 585
R369 B.n201 B.n194 585
R370 B.n200 B.n199 585
R371 B.n197 B.n195 585
R372 B.n162 B.n161 585
R373 B.n306 B.n305 585
R374 B.n307 B.n306 585
R375 B.n158 B.n157 585
R376 B.n159 B.n158 585
R377 B.n315 B.n314 585
R378 B.n314 B.n313 585
R379 B.n316 B.n156 585
R380 B.n156 B.n154 585
R381 B.n318 B.n317 585
R382 B.n319 B.n318 585
R383 B.n150 B.n149 585
R384 B.n155 B.n150 585
R385 B.n327 B.n326 585
R386 B.n326 B.n325 585
R387 B.n328 B.n148 585
R388 B.n148 B.n147 585
R389 B.n330 B.n329 585
R390 B.n331 B.n330 585
R391 B.n142 B.n141 585
R392 B.n143 B.n142 585
R393 B.n339 B.n338 585
R394 B.n338 B.n337 585
R395 B.n340 B.n140 585
R396 B.n140 B.n139 585
R397 B.n342 B.n341 585
R398 B.n343 B.n342 585
R399 B.n134 B.n133 585
R400 B.n135 B.n134 585
R401 B.n351 B.n350 585
R402 B.n350 B.n349 585
R403 B.n352 B.n132 585
R404 B.n132 B.n130 585
R405 B.n354 B.n353 585
R406 B.n355 B.n354 585
R407 B.n126 B.n125 585
R408 B.n131 B.n126 585
R409 B.n363 B.n362 585
R410 B.n362 B.n361 585
R411 B.n364 B.n124 585
R412 B.n124 B.n122 585
R413 B.n366 B.n365 585
R414 B.n367 B.n366 585
R415 B.n118 B.n117 585
R416 B.n123 B.n118 585
R417 B.n375 B.n374 585
R418 B.n374 B.n373 585
R419 B.n376 B.n116 585
R420 B.n116 B.n114 585
R421 B.n378 B.n377 585
R422 B.n379 B.n378 585
R423 B.n110 B.n109 585
R424 B.n115 B.n110 585
R425 B.n387 B.n386 585
R426 B.n386 B.n385 585
R427 B.n388 B.n108 585
R428 B.n108 B.n107 585
R429 B.n390 B.n389 585
R430 B.n391 B.n390 585
R431 B.n102 B.n101 585
R432 B.n103 B.n102 585
R433 B.n400 B.n399 585
R434 B.n399 B.n398 585
R435 B.n401 B.n100 585
R436 B.n100 B.n99 585
R437 B.n403 B.n402 585
R438 B.n404 B.n403 585
R439 B.n2 B.n0 585
R440 B.n4 B.n2 585
R441 B.n3 B.n1 585
R442 B.n629 B.n3 585
R443 B.n627 B.n626 585
R444 B.n628 B.n627 585
R445 B.n625 B.n9 585
R446 B.n9 B.n8 585
R447 B.n624 B.n623 585
R448 B.n623 B.n622 585
R449 B.n11 B.n10 585
R450 B.n621 B.n11 585
R451 B.n619 B.n618 585
R452 B.n620 B.n619 585
R453 B.n617 B.n16 585
R454 B.n16 B.n15 585
R455 B.n616 B.n615 585
R456 B.n615 B.n614 585
R457 B.n18 B.n17 585
R458 B.n613 B.n18 585
R459 B.n611 B.n610 585
R460 B.n612 B.n611 585
R461 B.n609 B.n23 585
R462 B.n23 B.n22 585
R463 B.n608 B.n607 585
R464 B.n607 B.n606 585
R465 B.n25 B.n24 585
R466 B.n605 B.n25 585
R467 B.n603 B.n602 585
R468 B.n604 B.n603 585
R469 B.n601 B.n30 585
R470 B.n30 B.n29 585
R471 B.n600 B.n599 585
R472 B.n599 B.n598 585
R473 B.n32 B.n31 585
R474 B.n597 B.n32 585
R475 B.n595 B.n594 585
R476 B.n596 B.n595 585
R477 B.n593 B.n37 585
R478 B.n37 B.n36 585
R479 B.n592 B.n591 585
R480 B.n591 B.n590 585
R481 B.n39 B.n38 585
R482 B.n589 B.n39 585
R483 B.n587 B.n586 585
R484 B.n588 B.n587 585
R485 B.n585 B.n44 585
R486 B.n44 B.n43 585
R487 B.n584 B.n583 585
R488 B.n583 B.n582 585
R489 B.n46 B.n45 585
R490 B.n581 B.n46 585
R491 B.n579 B.n578 585
R492 B.n580 B.n579 585
R493 B.n577 B.n51 585
R494 B.n51 B.n50 585
R495 B.n576 B.n575 585
R496 B.n575 B.n574 585
R497 B.n53 B.n52 585
R498 B.n573 B.n53 585
R499 B.n571 B.n570 585
R500 B.n572 B.n571 585
R501 B.n569 B.n58 585
R502 B.n58 B.n57 585
R503 B.n568 B.n567 585
R504 B.n567 B.n566 585
R505 B.n60 B.n59 585
R506 B.n565 B.n60 585
R507 B.n563 B.n562 585
R508 B.n564 B.n563 585
R509 B.n632 B.n631 585
R510 B.n631 B.n630 585
R511 B.n306 B.n164 569.379
R512 B.n563 B.n65 569.379
R513 B.n308 B.n162 569.379
R514 B.n452 B.n63 569.379
R515 B.n183 B.t8 322.043
R516 B.n177 B.t19 322.043
R517 B.n78 B.t16 322.043
R518 B.n85 B.t12 322.043
R519 B.n453 B.n64 256.663
R520 B.n459 B.n64 256.663
R521 B.n461 B.n64 256.663
R522 B.n467 B.n64 256.663
R523 B.n469 B.n64 256.663
R524 B.n475 B.n64 256.663
R525 B.n477 B.n64 256.663
R526 B.n483 B.n64 256.663
R527 B.n485 B.n64 256.663
R528 B.n491 B.n64 256.663
R529 B.n493 B.n64 256.663
R530 B.n500 B.n64 256.663
R531 B.n502 B.n64 256.663
R532 B.n508 B.n64 256.663
R533 B.n510 B.n64 256.663
R534 B.n516 B.n64 256.663
R535 B.n518 B.n64 256.663
R536 B.n524 B.n64 256.663
R537 B.n526 B.n64 256.663
R538 B.n532 B.n64 256.663
R539 B.n534 B.n64 256.663
R540 B.n540 B.n64 256.663
R541 B.n542 B.n64 256.663
R542 B.n548 B.n64 256.663
R543 B.n550 B.n64 256.663
R544 B.n556 B.n64 256.663
R545 B.n558 B.n64 256.663
R546 B.n301 B.n163 256.663
R547 B.n166 B.n163 256.663
R548 B.n294 B.n163 256.663
R549 B.n288 B.n163 256.663
R550 B.n286 B.n163 256.663
R551 B.n280 B.n163 256.663
R552 B.n278 B.n163 256.663
R553 B.n272 B.n163 256.663
R554 B.n270 B.n163 256.663
R555 B.n264 B.n163 256.663
R556 B.n262 B.n163 256.663
R557 B.n255 B.n163 256.663
R558 B.n253 B.n163 256.663
R559 B.n247 B.n163 256.663
R560 B.n245 B.n163 256.663
R561 B.n238 B.n163 256.663
R562 B.n236 B.n163 256.663
R563 B.n230 B.n163 256.663
R564 B.n228 B.n163 256.663
R565 B.n222 B.n163 256.663
R566 B.n220 B.n163 256.663
R567 B.n214 B.n163 256.663
R568 B.n212 B.n163 256.663
R569 B.n206 B.n163 256.663
R570 B.n204 B.n163 256.663
R571 B.n198 B.n163 256.663
R572 B.n196 B.n163 256.663
R573 B.n306 B.n158 163.367
R574 B.n314 B.n158 163.367
R575 B.n314 B.n156 163.367
R576 B.n318 B.n156 163.367
R577 B.n318 B.n150 163.367
R578 B.n326 B.n150 163.367
R579 B.n326 B.n148 163.367
R580 B.n330 B.n148 163.367
R581 B.n330 B.n142 163.367
R582 B.n338 B.n142 163.367
R583 B.n338 B.n140 163.367
R584 B.n342 B.n140 163.367
R585 B.n342 B.n134 163.367
R586 B.n350 B.n134 163.367
R587 B.n350 B.n132 163.367
R588 B.n354 B.n132 163.367
R589 B.n354 B.n126 163.367
R590 B.n362 B.n126 163.367
R591 B.n362 B.n124 163.367
R592 B.n366 B.n124 163.367
R593 B.n366 B.n118 163.367
R594 B.n374 B.n118 163.367
R595 B.n374 B.n116 163.367
R596 B.n378 B.n116 163.367
R597 B.n378 B.n110 163.367
R598 B.n386 B.n110 163.367
R599 B.n386 B.n108 163.367
R600 B.n390 B.n108 163.367
R601 B.n390 B.n102 163.367
R602 B.n399 B.n102 163.367
R603 B.n399 B.n100 163.367
R604 B.n403 B.n100 163.367
R605 B.n403 B.n2 163.367
R606 B.n631 B.n2 163.367
R607 B.n631 B.n3 163.367
R608 B.n627 B.n3 163.367
R609 B.n627 B.n9 163.367
R610 B.n623 B.n9 163.367
R611 B.n623 B.n11 163.367
R612 B.n619 B.n11 163.367
R613 B.n619 B.n16 163.367
R614 B.n615 B.n16 163.367
R615 B.n615 B.n18 163.367
R616 B.n611 B.n18 163.367
R617 B.n611 B.n23 163.367
R618 B.n607 B.n23 163.367
R619 B.n607 B.n25 163.367
R620 B.n603 B.n25 163.367
R621 B.n603 B.n30 163.367
R622 B.n599 B.n30 163.367
R623 B.n599 B.n32 163.367
R624 B.n595 B.n32 163.367
R625 B.n595 B.n37 163.367
R626 B.n591 B.n37 163.367
R627 B.n591 B.n39 163.367
R628 B.n587 B.n39 163.367
R629 B.n587 B.n44 163.367
R630 B.n583 B.n44 163.367
R631 B.n583 B.n46 163.367
R632 B.n579 B.n46 163.367
R633 B.n579 B.n51 163.367
R634 B.n575 B.n51 163.367
R635 B.n575 B.n53 163.367
R636 B.n571 B.n53 163.367
R637 B.n571 B.n58 163.367
R638 B.n567 B.n58 163.367
R639 B.n567 B.n60 163.367
R640 B.n563 B.n60 163.367
R641 B.n302 B.n300 163.367
R642 B.n300 B.n299 163.367
R643 B.n296 B.n295 163.367
R644 B.n293 B.n168 163.367
R645 B.n289 B.n287 163.367
R646 B.n285 B.n170 163.367
R647 B.n281 B.n279 163.367
R648 B.n277 B.n172 163.367
R649 B.n273 B.n271 163.367
R650 B.n269 B.n174 163.367
R651 B.n265 B.n263 163.367
R652 B.n261 B.n176 163.367
R653 B.n256 B.n254 163.367
R654 B.n252 B.n180 163.367
R655 B.n248 B.n246 163.367
R656 B.n244 B.n182 163.367
R657 B.n239 B.n237 163.367
R658 B.n235 B.n186 163.367
R659 B.n231 B.n229 163.367
R660 B.n227 B.n188 163.367
R661 B.n223 B.n221 163.367
R662 B.n219 B.n190 163.367
R663 B.n215 B.n213 163.367
R664 B.n211 B.n192 163.367
R665 B.n207 B.n205 163.367
R666 B.n203 B.n194 163.367
R667 B.n199 B.n197 163.367
R668 B.n308 B.n160 163.367
R669 B.n312 B.n160 163.367
R670 B.n312 B.n153 163.367
R671 B.n320 B.n153 163.367
R672 B.n320 B.n151 163.367
R673 B.n324 B.n151 163.367
R674 B.n324 B.n146 163.367
R675 B.n332 B.n146 163.367
R676 B.n332 B.n144 163.367
R677 B.n336 B.n144 163.367
R678 B.n336 B.n138 163.367
R679 B.n344 B.n138 163.367
R680 B.n344 B.n136 163.367
R681 B.n348 B.n136 163.367
R682 B.n348 B.n129 163.367
R683 B.n356 B.n129 163.367
R684 B.n356 B.n127 163.367
R685 B.n360 B.n127 163.367
R686 B.n360 B.n121 163.367
R687 B.n368 B.n121 163.367
R688 B.n368 B.n119 163.367
R689 B.n372 B.n119 163.367
R690 B.n372 B.n113 163.367
R691 B.n380 B.n113 163.367
R692 B.n380 B.n111 163.367
R693 B.n384 B.n111 163.367
R694 B.n384 B.n106 163.367
R695 B.n392 B.n106 163.367
R696 B.n392 B.n104 163.367
R697 B.n397 B.n104 163.367
R698 B.n397 B.n98 163.367
R699 B.n405 B.n98 163.367
R700 B.n406 B.n405 163.367
R701 B.n406 B.n5 163.367
R702 B.n6 B.n5 163.367
R703 B.n7 B.n6 163.367
R704 B.n411 B.n7 163.367
R705 B.n411 B.n12 163.367
R706 B.n13 B.n12 163.367
R707 B.n14 B.n13 163.367
R708 B.n416 B.n14 163.367
R709 B.n416 B.n19 163.367
R710 B.n20 B.n19 163.367
R711 B.n21 B.n20 163.367
R712 B.n421 B.n21 163.367
R713 B.n421 B.n26 163.367
R714 B.n27 B.n26 163.367
R715 B.n28 B.n27 163.367
R716 B.n426 B.n28 163.367
R717 B.n426 B.n33 163.367
R718 B.n34 B.n33 163.367
R719 B.n35 B.n34 163.367
R720 B.n431 B.n35 163.367
R721 B.n431 B.n40 163.367
R722 B.n41 B.n40 163.367
R723 B.n42 B.n41 163.367
R724 B.n436 B.n42 163.367
R725 B.n436 B.n47 163.367
R726 B.n48 B.n47 163.367
R727 B.n49 B.n48 163.367
R728 B.n441 B.n49 163.367
R729 B.n441 B.n54 163.367
R730 B.n55 B.n54 163.367
R731 B.n56 B.n55 163.367
R732 B.n446 B.n56 163.367
R733 B.n446 B.n61 163.367
R734 B.n62 B.n61 163.367
R735 B.n63 B.n62 163.367
R736 B.n559 B.n557 163.367
R737 B.n555 B.n67 163.367
R738 B.n551 B.n549 163.367
R739 B.n547 B.n69 163.367
R740 B.n543 B.n541 163.367
R741 B.n539 B.n71 163.367
R742 B.n535 B.n533 163.367
R743 B.n531 B.n73 163.367
R744 B.n527 B.n525 163.367
R745 B.n523 B.n75 163.367
R746 B.n519 B.n517 163.367
R747 B.n515 B.n77 163.367
R748 B.n511 B.n509 163.367
R749 B.n507 B.n82 163.367
R750 B.n503 B.n501 163.367
R751 B.n499 B.n84 163.367
R752 B.n494 B.n492 163.367
R753 B.n490 B.n88 163.367
R754 B.n486 B.n484 163.367
R755 B.n482 B.n90 163.367
R756 B.n478 B.n476 163.367
R757 B.n474 B.n92 163.367
R758 B.n470 B.n468 163.367
R759 B.n466 B.n94 163.367
R760 B.n462 B.n460 163.367
R761 B.n458 B.n96 163.367
R762 B.n454 B.n452 163.367
R763 B.n307 B.n163 140.083
R764 B.n564 B.n64 140.083
R765 B.n183 B.t11 102.257
R766 B.n85 B.t14 102.257
R767 B.n177 B.t21 102.251
R768 B.n78 B.t17 102.251
R769 B.n184 B.t10 73.5538
R770 B.n86 B.t15 73.5538
R771 B.n178 B.t20 73.548
R772 B.n79 B.t18 73.548
R773 B.n301 B.n164 71.676
R774 B.n299 B.n166 71.676
R775 B.n295 B.n294 71.676
R776 B.n288 B.n168 71.676
R777 B.n287 B.n286 71.676
R778 B.n280 B.n170 71.676
R779 B.n279 B.n278 71.676
R780 B.n272 B.n172 71.676
R781 B.n271 B.n270 71.676
R782 B.n264 B.n174 71.676
R783 B.n263 B.n262 71.676
R784 B.n255 B.n176 71.676
R785 B.n254 B.n253 71.676
R786 B.n247 B.n180 71.676
R787 B.n246 B.n245 71.676
R788 B.n238 B.n182 71.676
R789 B.n237 B.n236 71.676
R790 B.n230 B.n186 71.676
R791 B.n229 B.n228 71.676
R792 B.n222 B.n188 71.676
R793 B.n221 B.n220 71.676
R794 B.n214 B.n190 71.676
R795 B.n213 B.n212 71.676
R796 B.n206 B.n192 71.676
R797 B.n205 B.n204 71.676
R798 B.n198 B.n194 71.676
R799 B.n197 B.n196 71.676
R800 B.n558 B.n65 71.676
R801 B.n557 B.n556 71.676
R802 B.n550 B.n67 71.676
R803 B.n549 B.n548 71.676
R804 B.n542 B.n69 71.676
R805 B.n541 B.n540 71.676
R806 B.n534 B.n71 71.676
R807 B.n533 B.n532 71.676
R808 B.n526 B.n73 71.676
R809 B.n525 B.n524 71.676
R810 B.n518 B.n75 71.676
R811 B.n517 B.n516 71.676
R812 B.n510 B.n77 71.676
R813 B.n509 B.n508 71.676
R814 B.n502 B.n82 71.676
R815 B.n501 B.n500 71.676
R816 B.n493 B.n84 71.676
R817 B.n492 B.n491 71.676
R818 B.n485 B.n88 71.676
R819 B.n484 B.n483 71.676
R820 B.n477 B.n90 71.676
R821 B.n476 B.n475 71.676
R822 B.n469 B.n92 71.676
R823 B.n468 B.n467 71.676
R824 B.n461 B.n94 71.676
R825 B.n460 B.n459 71.676
R826 B.n453 B.n96 71.676
R827 B.n454 B.n453 71.676
R828 B.n459 B.n458 71.676
R829 B.n462 B.n461 71.676
R830 B.n467 B.n466 71.676
R831 B.n470 B.n469 71.676
R832 B.n475 B.n474 71.676
R833 B.n478 B.n477 71.676
R834 B.n483 B.n482 71.676
R835 B.n486 B.n485 71.676
R836 B.n491 B.n490 71.676
R837 B.n494 B.n493 71.676
R838 B.n500 B.n499 71.676
R839 B.n503 B.n502 71.676
R840 B.n508 B.n507 71.676
R841 B.n511 B.n510 71.676
R842 B.n516 B.n515 71.676
R843 B.n519 B.n518 71.676
R844 B.n524 B.n523 71.676
R845 B.n527 B.n526 71.676
R846 B.n532 B.n531 71.676
R847 B.n535 B.n534 71.676
R848 B.n540 B.n539 71.676
R849 B.n543 B.n542 71.676
R850 B.n548 B.n547 71.676
R851 B.n551 B.n550 71.676
R852 B.n556 B.n555 71.676
R853 B.n559 B.n558 71.676
R854 B.n302 B.n301 71.676
R855 B.n296 B.n166 71.676
R856 B.n294 B.n293 71.676
R857 B.n289 B.n288 71.676
R858 B.n286 B.n285 71.676
R859 B.n281 B.n280 71.676
R860 B.n278 B.n277 71.676
R861 B.n273 B.n272 71.676
R862 B.n270 B.n269 71.676
R863 B.n265 B.n264 71.676
R864 B.n262 B.n261 71.676
R865 B.n256 B.n255 71.676
R866 B.n253 B.n252 71.676
R867 B.n248 B.n247 71.676
R868 B.n245 B.n244 71.676
R869 B.n239 B.n238 71.676
R870 B.n236 B.n235 71.676
R871 B.n231 B.n230 71.676
R872 B.n228 B.n227 71.676
R873 B.n223 B.n222 71.676
R874 B.n220 B.n219 71.676
R875 B.n215 B.n214 71.676
R876 B.n212 B.n211 71.676
R877 B.n207 B.n206 71.676
R878 B.n204 B.n203 71.676
R879 B.n199 B.n198 71.676
R880 B.n196 B.n162 71.676
R881 B.n307 B.n159 68.53
R882 B.n313 B.n159 68.53
R883 B.n313 B.n154 68.53
R884 B.n319 B.n154 68.53
R885 B.n319 B.n155 68.53
R886 B.n325 B.n147 68.53
R887 B.n331 B.n147 68.53
R888 B.n331 B.n143 68.53
R889 B.n337 B.n143 68.53
R890 B.n337 B.n139 68.53
R891 B.n343 B.n139 68.53
R892 B.n349 B.n135 68.53
R893 B.n349 B.n130 68.53
R894 B.n355 B.n130 68.53
R895 B.n355 B.n131 68.53
R896 B.n361 B.n122 68.53
R897 B.n367 B.n122 68.53
R898 B.n367 B.n123 68.53
R899 B.n373 B.n114 68.53
R900 B.n379 B.n114 68.53
R901 B.n379 B.n115 68.53
R902 B.n385 B.n107 68.53
R903 B.n391 B.n107 68.53
R904 B.n391 B.n103 68.53
R905 B.n398 B.n103 68.53
R906 B.n404 B.n99 68.53
R907 B.n404 B.n4 68.53
R908 B.n630 B.n4 68.53
R909 B.n630 B.n629 68.53
R910 B.n629 B.n628 68.53
R911 B.n628 B.n8 68.53
R912 B.n622 B.n621 68.53
R913 B.n621 B.n620 68.53
R914 B.n620 B.n15 68.53
R915 B.n614 B.n15 68.53
R916 B.n613 B.n612 68.53
R917 B.n612 B.n22 68.53
R918 B.n606 B.n22 68.53
R919 B.n605 B.n604 68.53
R920 B.n604 B.n29 68.53
R921 B.n598 B.n29 68.53
R922 B.n597 B.n596 68.53
R923 B.n596 B.n36 68.53
R924 B.n590 B.n36 68.53
R925 B.n590 B.n589 68.53
R926 B.n588 B.n43 68.53
R927 B.n582 B.n43 68.53
R928 B.n582 B.n581 68.53
R929 B.n581 B.n580 68.53
R930 B.n580 B.n50 68.53
R931 B.n574 B.n50 68.53
R932 B.n573 B.n572 68.53
R933 B.n572 B.n57 68.53
R934 B.n566 B.n57 68.53
R935 B.n566 B.n565 68.53
R936 B.n565 B.n564 68.53
R937 B.n241 B.n184 59.5399
R938 B.n259 B.n178 59.5399
R939 B.n80 B.n79 59.5399
R940 B.n497 B.n86 59.5399
R941 B.n115 B.t2 59.46
R942 B.t22 B.n613 59.46
R943 B.n361 B.t5 57.4444
R944 B.n598 B.t0 57.4444
R945 B.n343 B.t4 55.4288
R946 B.t6 B.n588 55.4288
R947 B.t1 B.n99 53.4132
R948 B.t3 B.n8 53.4132
R949 B.n325 B.t9 51.3977
R950 B.n574 B.t13 51.3977
R951 B.n562 B.n561 36.9956
R952 B.n451 B.n450 36.9956
R953 B.n309 B.n161 36.9956
R954 B.n305 B.n304 36.9956
R955 B.n123 B.t23 35.2731
R956 B.t7 B.n605 35.2731
R957 B.n373 B.t23 33.2575
R958 B.n606 B.t7 33.2575
R959 B.n184 B.n183 28.7035
R960 B.n178 B.n177 28.7035
R961 B.n79 B.n78 28.7035
R962 B.n86 B.n85 28.7035
R963 B B.n632 18.0485
R964 B.n155 B.t9 17.1329
R965 B.t13 B.n573 17.1329
R966 B.n398 B.t1 15.1173
R967 B.n622 B.t3 15.1173
R968 B.t4 B.n135 13.1017
R969 B.n589 B.t6 13.1017
R970 B.n131 B.t5 11.0862
R971 B.t0 B.n597 11.0862
R972 B.n561 B.n560 10.6151
R973 B.n560 B.n66 10.6151
R974 B.n554 B.n66 10.6151
R975 B.n554 B.n553 10.6151
R976 B.n553 B.n552 10.6151
R977 B.n552 B.n68 10.6151
R978 B.n546 B.n68 10.6151
R979 B.n546 B.n545 10.6151
R980 B.n545 B.n544 10.6151
R981 B.n544 B.n70 10.6151
R982 B.n538 B.n70 10.6151
R983 B.n538 B.n537 10.6151
R984 B.n537 B.n536 10.6151
R985 B.n536 B.n72 10.6151
R986 B.n530 B.n72 10.6151
R987 B.n530 B.n529 10.6151
R988 B.n529 B.n528 10.6151
R989 B.n528 B.n74 10.6151
R990 B.n522 B.n74 10.6151
R991 B.n522 B.n521 10.6151
R992 B.n521 B.n520 10.6151
R993 B.n520 B.n76 10.6151
R994 B.n514 B.n513 10.6151
R995 B.n513 B.n512 10.6151
R996 B.n512 B.n81 10.6151
R997 B.n506 B.n81 10.6151
R998 B.n506 B.n505 10.6151
R999 B.n505 B.n504 10.6151
R1000 B.n504 B.n83 10.6151
R1001 B.n498 B.n83 10.6151
R1002 B.n496 B.n495 10.6151
R1003 B.n495 B.n87 10.6151
R1004 B.n489 B.n87 10.6151
R1005 B.n489 B.n488 10.6151
R1006 B.n488 B.n487 10.6151
R1007 B.n487 B.n89 10.6151
R1008 B.n481 B.n89 10.6151
R1009 B.n481 B.n480 10.6151
R1010 B.n480 B.n479 10.6151
R1011 B.n479 B.n91 10.6151
R1012 B.n473 B.n91 10.6151
R1013 B.n473 B.n472 10.6151
R1014 B.n472 B.n471 10.6151
R1015 B.n471 B.n93 10.6151
R1016 B.n465 B.n93 10.6151
R1017 B.n465 B.n464 10.6151
R1018 B.n464 B.n463 10.6151
R1019 B.n463 B.n95 10.6151
R1020 B.n457 B.n95 10.6151
R1021 B.n457 B.n456 10.6151
R1022 B.n456 B.n455 10.6151
R1023 B.n455 B.n451 10.6151
R1024 B.n310 B.n309 10.6151
R1025 B.n311 B.n310 10.6151
R1026 B.n311 B.n152 10.6151
R1027 B.n321 B.n152 10.6151
R1028 B.n322 B.n321 10.6151
R1029 B.n323 B.n322 10.6151
R1030 B.n323 B.n145 10.6151
R1031 B.n333 B.n145 10.6151
R1032 B.n334 B.n333 10.6151
R1033 B.n335 B.n334 10.6151
R1034 B.n335 B.n137 10.6151
R1035 B.n345 B.n137 10.6151
R1036 B.n346 B.n345 10.6151
R1037 B.n347 B.n346 10.6151
R1038 B.n347 B.n128 10.6151
R1039 B.n357 B.n128 10.6151
R1040 B.n358 B.n357 10.6151
R1041 B.n359 B.n358 10.6151
R1042 B.n359 B.n120 10.6151
R1043 B.n369 B.n120 10.6151
R1044 B.n370 B.n369 10.6151
R1045 B.n371 B.n370 10.6151
R1046 B.n371 B.n112 10.6151
R1047 B.n381 B.n112 10.6151
R1048 B.n382 B.n381 10.6151
R1049 B.n383 B.n382 10.6151
R1050 B.n383 B.n105 10.6151
R1051 B.n393 B.n105 10.6151
R1052 B.n394 B.n393 10.6151
R1053 B.n396 B.n394 10.6151
R1054 B.n396 B.n395 10.6151
R1055 B.n395 B.n97 10.6151
R1056 B.n407 B.n97 10.6151
R1057 B.n408 B.n407 10.6151
R1058 B.n409 B.n408 10.6151
R1059 B.n410 B.n409 10.6151
R1060 B.n412 B.n410 10.6151
R1061 B.n413 B.n412 10.6151
R1062 B.n414 B.n413 10.6151
R1063 B.n415 B.n414 10.6151
R1064 B.n417 B.n415 10.6151
R1065 B.n418 B.n417 10.6151
R1066 B.n419 B.n418 10.6151
R1067 B.n420 B.n419 10.6151
R1068 B.n422 B.n420 10.6151
R1069 B.n423 B.n422 10.6151
R1070 B.n424 B.n423 10.6151
R1071 B.n425 B.n424 10.6151
R1072 B.n427 B.n425 10.6151
R1073 B.n428 B.n427 10.6151
R1074 B.n429 B.n428 10.6151
R1075 B.n430 B.n429 10.6151
R1076 B.n432 B.n430 10.6151
R1077 B.n433 B.n432 10.6151
R1078 B.n434 B.n433 10.6151
R1079 B.n435 B.n434 10.6151
R1080 B.n437 B.n435 10.6151
R1081 B.n438 B.n437 10.6151
R1082 B.n439 B.n438 10.6151
R1083 B.n440 B.n439 10.6151
R1084 B.n442 B.n440 10.6151
R1085 B.n443 B.n442 10.6151
R1086 B.n444 B.n443 10.6151
R1087 B.n445 B.n444 10.6151
R1088 B.n447 B.n445 10.6151
R1089 B.n448 B.n447 10.6151
R1090 B.n449 B.n448 10.6151
R1091 B.n450 B.n449 10.6151
R1092 B.n304 B.n303 10.6151
R1093 B.n303 B.n165 10.6151
R1094 B.n298 B.n165 10.6151
R1095 B.n298 B.n297 10.6151
R1096 B.n297 B.n167 10.6151
R1097 B.n292 B.n167 10.6151
R1098 B.n292 B.n291 10.6151
R1099 B.n291 B.n290 10.6151
R1100 B.n290 B.n169 10.6151
R1101 B.n284 B.n169 10.6151
R1102 B.n284 B.n283 10.6151
R1103 B.n283 B.n282 10.6151
R1104 B.n282 B.n171 10.6151
R1105 B.n276 B.n171 10.6151
R1106 B.n276 B.n275 10.6151
R1107 B.n275 B.n274 10.6151
R1108 B.n274 B.n173 10.6151
R1109 B.n268 B.n173 10.6151
R1110 B.n268 B.n267 10.6151
R1111 B.n267 B.n266 10.6151
R1112 B.n266 B.n175 10.6151
R1113 B.n260 B.n175 10.6151
R1114 B.n258 B.n257 10.6151
R1115 B.n257 B.n179 10.6151
R1116 B.n251 B.n179 10.6151
R1117 B.n251 B.n250 10.6151
R1118 B.n250 B.n249 10.6151
R1119 B.n249 B.n181 10.6151
R1120 B.n243 B.n181 10.6151
R1121 B.n243 B.n242 10.6151
R1122 B.n240 B.n185 10.6151
R1123 B.n234 B.n185 10.6151
R1124 B.n234 B.n233 10.6151
R1125 B.n233 B.n232 10.6151
R1126 B.n232 B.n187 10.6151
R1127 B.n226 B.n187 10.6151
R1128 B.n226 B.n225 10.6151
R1129 B.n225 B.n224 10.6151
R1130 B.n224 B.n189 10.6151
R1131 B.n218 B.n189 10.6151
R1132 B.n218 B.n217 10.6151
R1133 B.n217 B.n216 10.6151
R1134 B.n216 B.n191 10.6151
R1135 B.n210 B.n191 10.6151
R1136 B.n210 B.n209 10.6151
R1137 B.n209 B.n208 10.6151
R1138 B.n208 B.n193 10.6151
R1139 B.n202 B.n193 10.6151
R1140 B.n202 B.n201 10.6151
R1141 B.n201 B.n200 10.6151
R1142 B.n200 B.n195 10.6151
R1143 B.n195 B.n161 10.6151
R1144 B.n305 B.n157 10.6151
R1145 B.n315 B.n157 10.6151
R1146 B.n316 B.n315 10.6151
R1147 B.n317 B.n316 10.6151
R1148 B.n317 B.n149 10.6151
R1149 B.n327 B.n149 10.6151
R1150 B.n328 B.n327 10.6151
R1151 B.n329 B.n328 10.6151
R1152 B.n329 B.n141 10.6151
R1153 B.n339 B.n141 10.6151
R1154 B.n340 B.n339 10.6151
R1155 B.n341 B.n340 10.6151
R1156 B.n341 B.n133 10.6151
R1157 B.n351 B.n133 10.6151
R1158 B.n352 B.n351 10.6151
R1159 B.n353 B.n352 10.6151
R1160 B.n353 B.n125 10.6151
R1161 B.n363 B.n125 10.6151
R1162 B.n364 B.n363 10.6151
R1163 B.n365 B.n364 10.6151
R1164 B.n365 B.n117 10.6151
R1165 B.n375 B.n117 10.6151
R1166 B.n376 B.n375 10.6151
R1167 B.n377 B.n376 10.6151
R1168 B.n377 B.n109 10.6151
R1169 B.n387 B.n109 10.6151
R1170 B.n388 B.n387 10.6151
R1171 B.n389 B.n388 10.6151
R1172 B.n389 B.n101 10.6151
R1173 B.n400 B.n101 10.6151
R1174 B.n401 B.n400 10.6151
R1175 B.n402 B.n401 10.6151
R1176 B.n402 B.n0 10.6151
R1177 B.n626 B.n1 10.6151
R1178 B.n626 B.n625 10.6151
R1179 B.n625 B.n624 10.6151
R1180 B.n624 B.n10 10.6151
R1181 B.n618 B.n10 10.6151
R1182 B.n618 B.n617 10.6151
R1183 B.n617 B.n616 10.6151
R1184 B.n616 B.n17 10.6151
R1185 B.n610 B.n17 10.6151
R1186 B.n610 B.n609 10.6151
R1187 B.n609 B.n608 10.6151
R1188 B.n608 B.n24 10.6151
R1189 B.n602 B.n24 10.6151
R1190 B.n602 B.n601 10.6151
R1191 B.n601 B.n600 10.6151
R1192 B.n600 B.n31 10.6151
R1193 B.n594 B.n31 10.6151
R1194 B.n594 B.n593 10.6151
R1195 B.n593 B.n592 10.6151
R1196 B.n592 B.n38 10.6151
R1197 B.n586 B.n38 10.6151
R1198 B.n586 B.n585 10.6151
R1199 B.n585 B.n584 10.6151
R1200 B.n584 B.n45 10.6151
R1201 B.n578 B.n45 10.6151
R1202 B.n578 B.n577 10.6151
R1203 B.n577 B.n576 10.6151
R1204 B.n576 B.n52 10.6151
R1205 B.n570 B.n52 10.6151
R1206 B.n570 B.n569 10.6151
R1207 B.n569 B.n568 10.6151
R1208 B.n568 B.n59 10.6151
R1209 B.n562 B.n59 10.6151
R1210 B.n385 B.t2 9.07059
R1211 B.n614 B.t22 9.07059
R1212 B.n514 B.n80 6.5566
R1213 B.n498 B.n497 6.5566
R1214 B.n259 B.n258 6.5566
R1215 B.n242 B.n241 6.5566
R1216 B.n80 B.n76 4.05904
R1217 B.n497 B.n496 4.05904
R1218 B.n260 B.n259 4.05904
R1219 B.n241 B.n240 4.05904
R1220 B.n632 B.n0 2.81026
R1221 B.n632 B.n1 2.81026
R1222 VP.n10 VP.t1 175.499
R1223 VP.n13 VP.n12 161.3
R1224 VP.n14 VP.n9 161.3
R1225 VP.n16 VP.n15 161.3
R1226 VP.n17 VP.n8 161.3
R1227 VP.n19 VP.n18 161.3
R1228 VP.n21 VP.n20 161.3
R1229 VP.n22 VP.n6 161.3
R1230 VP.n40 VP.n0 161.3
R1231 VP.n39 VP.n38 161.3
R1232 VP.n37 VP.n36 161.3
R1233 VP.n35 VP.n2 161.3
R1234 VP.n34 VP.n33 161.3
R1235 VP.n32 VP.n3 161.3
R1236 VP.n31 VP.n30 161.3
R1237 VP.n28 VP.n4 161.3
R1238 VP.n27 VP.n26 161.3
R1239 VP.n5 VP.t9 152.355
R1240 VP.n41 VP.t8 152.355
R1241 VP.n23 VP.t5 152.355
R1242 VP.n34 VP.t0 118.195
R1243 VP.n29 VP.t6 118.195
R1244 VP.n1 VP.t2 118.195
R1245 VP.n16 VP.t7 118.195
R1246 VP.n7 VP.t3 118.195
R1247 VP.n11 VP.t4 118.195
R1248 VP.n24 VP.n23 80.6037
R1249 VP.n42 VP.n41 80.6037
R1250 VP.n25 VP.n5 80.6037
R1251 VP.n36 VP.n35 56.5617
R1252 VP.n12 VP.n9 56.5617
R1253 VP.n30 VP.n3 56.5617
R1254 VP.n18 VP.n17 56.5617
R1255 VP.n27 VP.n5 50.9056
R1256 VP.n41 VP.n40 50.9056
R1257 VP.n23 VP.n22 50.9056
R1258 VP.n25 VP.n24 40.6377
R1259 VP.n11 VP.n10 33.7965
R1260 VP.n13 VP.n10 28.0737
R1261 VP.n28 VP.n27 24.5923
R1262 VP.n34 VP.n3 24.5923
R1263 VP.n35 VP.n34 24.5923
R1264 VP.n40 VP.n39 24.5923
R1265 VP.n22 VP.n21 24.5923
R1266 VP.n16 VP.n9 24.5923
R1267 VP.n17 VP.n16 24.5923
R1268 VP.n30 VP.n29 23.6087
R1269 VP.n36 VP.n1 23.6087
R1270 VP.n18 VP.n7 23.6087
R1271 VP.n12 VP.n11 23.6087
R1272 VP.n29 VP.n28 0.984173
R1273 VP.n39 VP.n1 0.984173
R1274 VP.n21 VP.n7 0.984173
R1275 VP.n24 VP.n6 0.285035
R1276 VP.n26 VP.n25 0.285035
R1277 VP.n42 VP.n0 0.285035
R1278 VP.n14 VP.n13 0.189894
R1279 VP.n15 VP.n14 0.189894
R1280 VP.n15 VP.n8 0.189894
R1281 VP.n19 VP.n8 0.189894
R1282 VP.n20 VP.n19 0.189894
R1283 VP.n20 VP.n6 0.189894
R1284 VP.n26 VP.n4 0.189894
R1285 VP.n31 VP.n4 0.189894
R1286 VP.n32 VP.n31 0.189894
R1287 VP.n33 VP.n32 0.189894
R1288 VP.n33 VP.n2 0.189894
R1289 VP.n37 VP.n2 0.189894
R1290 VP.n38 VP.n37 0.189894
R1291 VP.n38 VP.n0 0.189894
R1292 VP VP.n42 0.146778
R1293 VDD1.n1 VDD1.t8 72.6565
R1294 VDD1.n3 VDD1.t0 72.6563
R1295 VDD1.n5 VDD1.n4 68.7714
R1296 VDD1.n1 VDD1.n0 67.87
R1297 VDD1.n7 VDD1.n6 67.8699
R1298 VDD1.n3 VDD1.n2 67.8698
R1299 VDD1.n7 VDD1.n5 35.8587
R1300 VDD1.n6 VDD1.t6 3.51114
R1301 VDD1.n6 VDD1.t4 3.51114
R1302 VDD1.n0 VDD1.t5 3.51114
R1303 VDD1.n0 VDD1.t2 3.51114
R1304 VDD1.n4 VDD1.t7 3.51114
R1305 VDD1.n4 VDD1.t1 3.51114
R1306 VDD1.n2 VDD1.t3 3.51114
R1307 VDD1.n2 VDD1.t9 3.51114
R1308 VDD1 VDD1.n7 0.899207
R1309 VDD1 VDD1.n1 0.377655
R1310 VDD1.n5 VDD1.n3 0.26412
C0 VTAIL VDD2 7.18145f
C1 VDD1 VP 4.44366f
C2 VN VDD2 4.19816f
C3 VDD1 VDD2 1.24759f
C4 VTAIL VN 4.59061f
C5 VP VDD2 0.398463f
C6 VDD1 VTAIL 7.13998f
C7 VDD1 VN 0.150512f
C8 VTAIL VP 4.60489f
C9 VP VN 5.07559f
C10 VDD2 B 4.371315f
C11 VDD1 B 4.324271f
C12 VTAIL B 4.356688f
C13 VN B 10.686339f
C14 VP B 9.123654f
C15 VDD1.t8 B 1.09718f
C16 VDD1.t5 B 0.103805f
C17 VDD1.t2 B 0.103805f
C18 VDD1.n0 B 0.859106f
C19 VDD1.n1 B 0.649984f
C20 VDD1.t0 B 1.09718f
C21 VDD1.t3 B 0.103805f
C22 VDD1.t9 B 0.103805f
C23 VDD1.n2 B 0.859103f
C24 VDD1.n3 B 0.643518f
C25 VDD1.t7 B 0.103805f
C26 VDD1.t1 B 0.103805f
C27 VDD1.n4 B 0.863839f
C28 VDD1.n5 B 1.71727f
C29 VDD1.t6 B 0.103805f
C30 VDD1.t4 B 0.103805f
C31 VDD1.n6 B 0.859102f
C32 VDD1.n7 B 1.92752f
C33 VP.n0 B 0.049428f
C34 VP.t2 B 0.63351f
C35 VP.n1 B 0.258345f
C36 VP.n2 B 0.037042f
C37 VP.t0 B 0.63351f
C38 VP.n3 B 0.052821f
C39 VP.n4 B 0.037042f
C40 VP.t6 B 0.63351f
C41 VP.t9 B 0.698373f
C42 VP.n5 B 0.325434f
C43 VP.n6 B 0.049428f
C44 VP.t5 B 0.698373f
C45 VP.t3 B 0.63351f
C46 VP.n7 B 0.258345f
C47 VP.n8 B 0.037042f
C48 VP.t7 B 0.63351f
C49 VP.n9 B 0.052821f
C50 VP.t1 B 0.742543f
C51 VP.n10 B 0.307937f
C52 VP.t4 B 0.63351f
C53 VP.n11 B 0.318857f
C54 VP.n12 B 0.053514f
C55 VP.n13 B 0.196357f
C56 VP.n14 B 0.037042f
C57 VP.n15 B 0.037042f
C58 VP.n16 B 0.293125f
C59 VP.n17 B 0.052821f
C60 VP.n18 B 0.053514f
C61 VP.n19 B 0.037042f
C62 VP.n20 B 0.037042f
C63 VP.n21 B 0.036136f
C64 VP.n22 B 0.049178f
C65 VP.n23 B 0.325434f
C66 VP.n24 B 1.45945f
C67 VP.n25 B 1.49231f
C68 VP.n26 B 0.049428f
C69 VP.n27 B 0.049178f
C70 VP.n28 B 0.036136f
C71 VP.n29 B 0.258345f
C72 VP.n30 B 0.053514f
C73 VP.n31 B 0.037042f
C74 VP.n32 B 0.037042f
C75 VP.n33 B 0.037042f
C76 VP.n34 B 0.293125f
C77 VP.n35 B 0.052821f
C78 VP.n36 B 0.053514f
C79 VP.n37 B 0.037042f
C80 VP.n38 B 0.037042f
C81 VP.n39 B 0.036136f
C82 VP.n40 B 0.049178f
C83 VP.t8 B 0.698373f
C84 VP.n41 B 0.325434f
C85 VP.n42 B 0.034691f
C86 VTAIL.t16 B 0.121115f
C87 VTAIL.t12 B 0.121115f
C88 VTAIL.n0 B 0.932617f
C89 VTAIL.n1 B 0.437901f
C90 VTAIL.t1 B 1.18965f
C91 VTAIL.n2 B 0.534015f
C92 VTAIL.t19 B 0.121115f
C93 VTAIL.t2 B 0.121115f
C94 VTAIL.n3 B 0.932617f
C95 VTAIL.n4 B 0.475455f
C96 VTAIL.t4 B 0.121115f
C97 VTAIL.t5 B 0.121115f
C98 VTAIL.n5 B 0.932617f
C99 VTAIL.n6 B 1.38205f
C100 VTAIL.t17 B 0.121115f
C101 VTAIL.t9 B 0.121115f
C102 VTAIL.n7 B 0.932623f
C103 VTAIL.n8 B 1.38204f
C104 VTAIL.t15 B 0.121115f
C105 VTAIL.t18 B 0.121115f
C106 VTAIL.n9 B 0.932623f
C107 VTAIL.n10 B 0.47545f
C108 VTAIL.t10 B 1.18966f
C109 VTAIL.n11 B 0.53401f
C110 VTAIL.t3 B 0.121115f
C111 VTAIL.t8 B 0.121115f
C112 VTAIL.n12 B 0.932623f
C113 VTAIL.n13 B 0.46073f
C114 VTAIL.t7 B 0.121115f
C115 VTAIL.t0 B 0.121115f
C116 VTAIL.n14 B 0.932623f
C117 VTAIL.n15 B 0.47545f
C118 VTAIL.t6 B 1.18965f
C119 VTAIL.n16 B 1.34361f
C120 VTAIL.t13 B 1.18965f
C121 VTAIL.n17 B 1.34361f
C122 VTAIL.t14 B 0.121115f
C123 VTAIL.t11 B 0.121115f
C124 VTAIL.n18 B 0.932617f
C125 VTAIL.n19 B 0.386571f
C126 VDD2.t7 B 1.09584f
C127 VDD2.t5 B 0.103678f
C128 VDD2.t1 B 0.103678f
C129 VDD2.n0 B 0.858051f
C130 VDD2.n1 B 0.64273f
C131 VDD2.t2 B 0.103678f
C132 VDD2.t9 B 0.103678f
C133 VDD2.n2 B 0.862781f
C134 VDD2.n3 B 1.63673f
C135 VDD2.t0 B 1.0898f
C136 VDD2.n4 B 1.90132f
C137 VDD2.t8 B 0.103678f
C138 VDD2.t4 B 0.103678f
C139 VDD2.n5 B 0.858054f
C140 VDD2.n6 B 0.311558f
C141 VDD2.t6 B 0.103678f
C142 VDD2.t3 B 0.103678f
C143 VDD2.n7 B 0.862755f
C144 VN.n0 B 0.048547f
C145 VN.t7 B 0.622226f
C146 VN.n1 B 0.253744f
C147 VN.n2 B 0.036382f
C148 VN.t4 B 0.622226f
C149 VN.n3 B 0.05188f
C150 VN.t2 B 0.729317f
C151 VN.n4 B 0.302452f
C152 VN.t6 B 0.622226f
C153 VN.n5 B 0.313177f
C154 VN.n6 B 0.052561f
C155 VN.n7 B 0.19286f
C156 VN.n8 B 0.036382f
C157 VN.n9 B 0.036382f
C158 VN.n10 B 0.287904f
C159 VN.n11 B 0.05188f
C160 VN.n12 B 0.052561f
C161 VN.n13 B 0.036382f
C162 VN.n14 B 0.036382f
C163 VN.n15 B 0.035493f
C164 VN.n16 B 0.048302f
C165 VN.t5 B 0.685934f
C166 VN.n17 B 0.319638f
C167 VN.n18 B 0.034073f
C168 VN.n19 B 0.048547f
C169 VN.t9 B 0.622226f
C170 VN.n20 B 0.253744f
C171 VN.n21 B 0.036382f
C172 VN.t3 B 0.622226f
C173 VN.n22 B 0.05188f
C174 VN.t8 B 0.729317f
C175 VN.n23 B 0.302452f
C176 VN.t0 B 0.622226f
C177 VN.n24 B 0.313177f
C178 VN.n25 B 0.052561f
C179 VN.n26 B 0.19286f
C180 VN.n27 B 0.036382f
C181 VN.n28 B 0.036382f
C182 VN.n29 B 0.287904f
C183 VN.n30 B 0.05188f
C184 VN.n31 B 0.052561f
C185 VN.n32 B 0.036382f
C186 VN.n33 B 0.036382f
C187 VN.n34 B 0.035493f
C188 VN.n35 B 0.048302f
C189 VN.t1 B 0.685934f
C190 VN.n36 B 0.319638f
C191 VN.n37 B 1.45398f
.ends

