* NGSPICE file created from diff_pair_sample_0269.ext - technology: sky130A

.subckt diff_pair_sample_0269 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.546 ps=3.58 w=1.4 l=2.31
X1 VTAIL.t8 VP.t1 VDD1.t6 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X2 VDD1.t5 VP.t2 VTAIL.t12 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X3 VTAIL.t10 VP.t3 VDD1.t4 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0.231 ps=1.73 w=1.4 l=2.31
X4 B.t11 B.t9 B.t10 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0 ps=0 w=1.4 l=2.31
X5 B.t8 B.t6 B.t7 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0 ps=0 w=1.4 l=2.31
X6 VTAIL.t5 VN.t0 VDD2.t7 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0.231 ps=1.73 w=1.4 l=2.31
X7 VTAIL.t13 VP.t4 VDD1.t3 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0.231 ps=1.73 w=1.4 l=2.31
X8 VDD2.t6 VN.t1 VTAIL.t3 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X9 VDD2.t5 VN.t2 VTAIL.t6 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.546 ps=3.58 w=1.4 l=2.31
X10 B.t5 B.t3 B.t4 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0 ps=0 w=1.4 l=2.31
X11 VDD1.t2 VP.t5 VTAIL.t15 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X12 B.t2 B.t0 B.t1 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0 ps=0 w=1.4 l=2.31
X13 VDD2.t4 VN.t3 VTAIL.t7 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.546 ps=3.58 w=1.4 l=2.31
X14 VDD1.t1 VP.t6 VTAIL.t14 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.546 ps=3.58 w=1.4 l=2.31
X15 VDD2.t3 VN.t4 VTAIL.t4 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X16 VTAIL.t0 VN.t5 VDD2.t2 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X17 VTAIL.t1 VN.t6 VDD2.t1 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X18 VTAIL.t11 VP.t7 VDD1.t0 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.231 pd=1.73 as=0.231 ps=1.73 w=1.4 l=2.31
X19 VTAIL.t2 VN.t7 VDD2.t0 w_n3610_n1248# sky130_fd_pr__pfet_01v8 ad=0.546 pd=3.58 as=0.231 ps=1.73 w=1.4 l=2.31
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n26 VP.n10 161.3
R7 VP.n28 VP.n27 161.3
R8 VP.n29 VP.n9 161.3
R9 VP.n31 VP.n30 161.3
R10 VP.n32 VP.n8 161.3
R11 VP.n62 VP.n0 161.3
R12 VP.n61 VP.n60 161.3
R13 VP.n59 VP.n1 161.3
R14 VP.n58 VP.n57 161.3
R15 VP.n56 VP.n2 161.3
R16 VP.n54 VP.n53 161.3
R17 VP.n52 VP.n3 161.3
R18 VP.n51 VP.n50 161.3
R19 VP.n49 VP.n4 161.3
R20 VP.n48 VP.n47 161.3
R21 VP.n46 VP.n5 161.3
R22 VP.n45 VP.n44 161.3
R23 VP.n42 VP.n6 161.3
R24 VP.n41 VP.n40 161.3
R25 VP.n39 VP.n7 161.3
R26 VP.n38 VP.n37 161.3
R27 VP.n36 VP.n35 100.579
R28 VP.n64 VP.n63 100.579
R29 VP.n34 VP.n33 100.579
R30 VP.n15 VP.n14 68.9827
R31 VP.n50 VP.n49 56.5617
R32 VP.n20 VP.n19 56.5617
R33 VP.n42 VP.n41 51.2335
R34 VP.n57 VP.n1 51.2335
R35 VP.n27 VP.n9 51.2335
R36 VP.n15 VP.t3 45.6612
R37 VP.n35 VP.n34 41.4618
R38 VP.n41 VP.n7 29.9206
R39 VP.n61 VP.n1 29.9206
R40 VP.n31 VP.n9 29.9206
R41 VP.n37 VP.n7 24.5923
R42 VP.n44 VP.n42 24.5923
R43 VP.n48 VP.n5 24.5923
R44 VP.n49 VP.n48 24.5923
R45 VP.n50 VP.n3 24.5923
R46 VP.n54 VP.n3 24.5923
R47 VP.n57 VP.n56 24.5923
R48 VP.n62 VP.n61 24.5923
R49 VP.n32 VP.n31 24.5923
R50 VP.n20 VP.n11 24.5923
R51 VP.n24 VP.n11 24.5923
R52 VP.n27 VP.n26 24.5923
R53 VP.n18 VP.n13 24.5923
R54 VP.n19 VP.n18 24.5923
R55 VP.n44 VP.n43 21.1495
R56 VP.n56 VP.n55 21.1495
R57 VP.n26 VP.n25 21.1495
R58 VP.n36 VP.t4 14.6066
R59 VP.n43 VP.t2 14.6066
R60 VP.n55 VP.t1 14.6066
R61 VP.n63 VP.t6 14.6066
R62 VP.n33 VP.t0 14.6066
R63 VP.n25 VP.t7 14.6066
R64 VP.n14 VP.t5 14.6066
R65 VP.n37 VP.n36 10.3291
R66 VP.n63 VP.n62 10.3291
R67 VP.n33 VP.n32 10.3291
R68 VP.n16 VP.n15 9.96756
R69 VP.n43 VP.n5 3.44336
R70 VP.n55 VP.n54 3.44336
R71 VP.n25 VP.n24 3.44336
R72 VP.n14 VP.n13 3.44336
R73 VP.n34 VP.n8 0.278335
R74 VP.n38 VP.n35 0.278335
R75 VP.n64 VP.n0 0.278335
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153485
R102 VTAIL.n11 VTAIL.t10 255.553
R103 VTAIL.n10 VTAIL.t6 255.553
R104 VTAIL.n7 VTAIL.t2 255.553
R105 VTAIL.n15 VTAIL.t7 255.552
R106 VTAIL.n2 VTAIL.t5 255.552
R107 VTAIL.n3 VTAIL.t14 255.552
R108 VTAIL.n6 VTAIL.t13 255.552
R109 VTAIL.n14 VTAIL.t9 255.552
R110 VTAIL.n13 VTAIL.n12 232.334
R111 VTAIL.n9 VTAIL.n8 232.334
R112 VTAIL.n1 VTAIL.n0 232.334
R113 VTAIL.n5 VTAIL.n4 232.334
R114 VTAIL.n0 VTAIL.t4 23.2184
R115 VTAIL.n0 VTAIL.t1 23.2184
R116 VTAIL.n4 VTAIL.t12 23.2184
R117 VTAIL.n4 VTAIL.t8 23.2184
R118 VTAIL.n12 VTAIL.t15 23.2184
R119 VTAIL.n12 VTAIL.t11 23.2184
R120 VTAIL.n8 VTAIL.t3 23.2184
R121 VTAIL.n8 VTAIL.t0 23.2184
R122 VTAIL.n15 VTAIL.n14 15.8496
R123 VTAIL.n7 VTAIL.n6 15.8496
R124 VTAIL.n9 VTAIL.n7 2.27636
R125 VTAIL.n10 VTAIL.n9 2.27636
R126 VTAIL.n13 VTAIL.n11 2.27636
R127 VTAIL.n14 VTAIL.n13 2.27636
R128 VTAIL.n6 VTAIL.n5 2.27636
R129 VTAIL.n5 VTAIL.n3 2.27636
R130 VTAIL.n2 VTAIL.n1 2.27636
R131 VTAIL VTAIL.n15 2.21817
R132 VTAIL.n11 VTAIL.n10 0.470328
R133 VTAIL.n3 VTAIL.n2 0.470328
R134 VTAIL VTAIL.n1 0.0586897
R135 VDD1 VDD1.n0 250.209
R136 VDD1.n3 VDD1.n2 250.095
R137 VDD1.n3 VDD1.n1 250.095
R138 VDD1.n5 VDD1.n4 249.012
R139 VDD1.n5 VDD1.n3 35.7466
R140 VDD1.n4 VDD1.t0 23.2184
R141 VDD1.n4 VDD1.t7 23.2184
R142 VDD1.n0 VDD1.t4 23.2184
R143 VDD1.n0 VDD1.t2 23.2184
R144 VDD1.n2 VDD1.t6 23.2184
R145 VDD1.n2 VDD1.t1 23.2184
R146 VDD1.n1 VDD1.t3 23.2184
R147 VDD1.n1 VDD1.t5 23.2184
R148 VDD1 VDD1.n5 1.08024
R149 B.n394 B.n45 585
R150 B.n396 B.n395 585
R151 B.n397 B.n44 585
R152 B.n399 B.n398 585
R153 B.n400 B.n43 585
R154 B.n402 B.n401 585
R155 B.n403 B.n42 585
R156 B.n405 B.n404 585
R157 B.n406 B.n41 585
R158 B.n408 B.n407 585
R159 B.n410 B.n38 585
R160 B.n412 B.n411 585
R161 B.n413 B.n37 585
R162 B.n415 B.n414 585
R163 B.n416 B.n36 585
R164 B.n418 B.n417 585
R165 B.n419 B.n35 585
R166 B.n421 B.n420 585
R167 B.n422 B.n31 585
R168 B.n424 B.n423 585
R169 B.n425 B.n30 585
R170 B.n427 B.n426 585
R171 B.n428 B.n29 585
R172 B.n430 B.n429 585
R173 B.n431 B.n28 585
R174 B.n433 B.n432 585
R175 B.n434 B.n27 585
R176 B.n436 B.n435 585
R177 B.n437 B.n26 585
R178 B.n439 B.n438 585
R179 B.n393 B.n392 585
R180 B.n391 B.n46 585
R181 B.n390 B.n389 585
R182 B.n388 B.n47 585
R183 B.n387 B.n386 585
R184 B.n385 B.n48 585
R185 B.n384 B.n383 585
R186 B.n382 B.n49 585
R187 B.n381 B.n380 585
R188 B.n379 B.n50 585
R189 B.n378 B.n377 585
R190 B.n376 B.n51 585
R191 B.n375 B.n374 585
R192 B.n373 B.n52 585
R193 B.n372 B.n371 585
R194 B.n370 B.n53 585
R195 B.n369 B.n368 585
R196 B.n367 B.n54 585
R197 B.n366 B.n365 585
R198 B.n364 B.n55 585
R199 B.n363 B.n362 585
R200 B.n361 B.n56 585
R201 B.n360 B.n359 585
R202 B.n358 B.n57 585
R203 B.n357 B.n356 585
R204 B.n355 B.n58 585
R205 B.n354 B.n353 585
R206 B.n352 B.n59 585
R207 B.n351 B.n350 585
R208 B.n349 B.n60 585
R209 B.n348 B.n347 585
R210 B.n346 B.n61 585
R211 B.n345 B.n344 585
R212 B.n343 B.n62 585
R213 B.n342 B.n341 585
R214 B.n340 B.n63 585
R215 B.n339 B.n338 585
R216 B.n337 B.n64 585
R217 B.n336 B.n335 585
R218 B.n334 B.n65 585
R219 B.n333 B.n332 585
R220 B.n331 B.n66 585
R221 B.n330 B.n329 585
R222 B.n328 B.n67 585
R223 B.n327 B.n326 585
R224 B.n325 B.n68 585
R225 B.n324 B.n323 585
R226 B.n322 B.n69 585
R227 B.n321 B.n320 585
R228 B.n319 B.n70 585
R229 B.n318 B.n317 585
R230 B.n316 B.n71 585
R231 B.n315 B.n314 585
R232 B.n313 B.n72 585
R233 B.n312 B.n311 585
R234 B.n310 B.n73 585
R235 B.n309 B.n308 585
R236 B.n307 B.n74 585
R237 B.n306 B.n305 585
R238 B.n304 B.n75 585
R239 B.n303 B.n302 585
R240 B.n301 B.n76 585
R241 B.n300 B.n299 585
R242 B.n298 B.n77 585
R243 B.n297 B.n296 585
R244 B.n295 B.n78 585
R245 B.n294 B.n293 585
R246 B.n292 B.n79 585
R247 B.n291 B.n290 585
R248 B.n289 B.n80 585
R249 B.n288 B.n287 585
R250 B.n286 B.n81 585
R251 B.n285 B.n284 585
R252 B.n283 B.n82 585
R253 B.n282 B.n281 585
R254 B.n280 B.n83 585
R255 B.n279 B.n278 585
R256 B.n277 B.n84 585
R257 B.n276 B.n275 585
R258 B.n274 B.n85 585
R259 B.n273 B.n272 585
R260 B.n271 B.n86 585
R261 B.n270 B.n269 585
R262 B.n268 B.n87 585
R263 B.n267 B.n266 585
R264 B.n265 B.n88 585
R265 B.n264 B.n263 585
R266 B.n262 B.n89 585
R267 B.n261 B.n260 585
R268 B.n259 B.n90 585
R269 B.n258 B.n257 585
R270 B.n256 B.n91 585
R271 B.n255 B.n254 585
R272 B.n253 B.n92 585
R273 B.n252 B.n251 585
R274 B.n205 B.n112 585
R275 B.n207 B.n206 585
R276 B.n208 B.n111 585
R277 B.n210 B.n209 585
R278 B.n211 B.n110 585
R279 B.n213 B.n212 585
R280 B.n214 B.n109 585
R281 B.n216 B.n215 585
R282 B.n217 B.n108 585
R283 B.n219 B.n218 585
R284 B.n221 B.n220 585
R285 B.n222 B.n104 585
R286 B.n224 B.n223 585
R287 B.n225 B.n103 585
R288 B.n227 B.n226 585
R289 B.n228 B.n102 585
R290 B.n230 B.n229 585
R291 B.n231 B.n101 585
R292 B.n233 B.n232 585
R293 B.n234 B.n98 585
R294 B.n237 B.n236 585
R295 B.n238 B.n97 585
R296 B.n240 B.n239 585
R297 B.n241 B.n96 585
R298 B.n243 B.n242 585
R299 B.n244 B.n95 585
R300 B.n246 B.n245 585
R301 B.n247 B.n94 585
R302 B.n249 B.n248 585
R303 B.n250 B.n93 585
R304 B.n204 B.n203 585
R305 B.n202 B.n113 585
R306 B.n201 B.n200 585
R307 B.n199 B.n114 585
R308 B.n198 B.n197 585
R309 B.n196 B.n115 585
R310 B.n195 B.n194 585
R311 B.n193 B.n116 585
R312 B.n192 B.n191 585
R313 B.n190 B.n117 585
R314 B.n189 B.n188 585
R315 B.n187 B.n118 585
R316 B.n186 B.n185 585
R317 B.n184 B.n119 585
R318 B.n183 B.n182 585
R319 B.n181 B.n120 585
R320 B.n180 B.n179 585
R321 B.n178 B.n121 585
R322 B.n177 B.n176 585
R323 B.n175 B.n122 585
R324 B.n174 B.n173 585
R325 B.n172 B.n123 585
R326 B.n171 B.n170 585
R327 B.n169 B.n124 585
R328 B.n168 B.n167 585
R329 B.n166 B.n125 585
R330 B.n165 B.n164 585
R331 B.n163 B.n126 585
R332 B.n162 B.n161 585
R333 B.n160 B.n127 585
R334 B.n159 B.n158 585
R335 B.n157 B.n128 585
R336 B.n156 B.n155 585
R337 B.n154 B.n129 585
R338 B.n153 B.n152 585
R339 B.n151 B.n130 585
R340 B.n150 B.n149 585
R341 B.n148 B.n131 585
R342 B.n147 B.n146 585
R343 B.n145 B.n132 585
R344 B.n144 B.n143 585
R345 B.n142 B.n133 585
R346 B.n141 B.n140 585
R347 B.n139 B.n134 585
R348 B.n138 B.n137 585
R349 B.n136 B.n135 585
R350 B.n2 B.n0 585
R351 B.n509 B.n1 585
R352 B.n508 B.n507 585
R353 B.n506 B.n3 585
R354 B.n505 B.n504 585
R355 B.n503 B.n4 585
R356 B.n502 B.n501 585
R357 B.n500 B.n5 585
R358 B.n499 B.n498 585
R359 B.n497 B.n6 585
R360 B.n496 B.n495 585
R361 B.n494 B.n7 585
R362 B.n493 B.n492 585
R363 B.n491 B.n8 585
R364 B.n490 B.n489 585
R365 B.n488 B.n9 585
R366 B.n487 B.n486 585
R367 B.n485 B.n10 585
R368 B.n484 B.n483 585
R369 B.n482 B.n11 585
R370 B.n481 B.n480 585
R371 B.n479 B.n12 585
R372 B.n478 B.n477 585
R373 B.n476 B.n13 585
R374 B.n475 B.n474 585
R375 B.n473 B.n14 585
R376 B.n472 B.n471 585
R377 B.n470 B.n15 585
R378 B.n469 B.n468 585
R379 B.n467 B.n16 585
R380 B.n466 B.n465 585
R381 B.n464 B.n17 585
R382 B.n463 B.n462 585
R383 B.n461 B.n18 585
R384 B.n460 B.n459 585
R385 B.n458 B.n19 585
R386 B.n457 B.n456 585
R387 B.n455 B.n20 585
R388 B.n454 B.n453 585
R389 B.n452 B.n21 585
R390 B.n451 B.n450 585
R391 B.n449 B.n22 585
R392 B.n448 B.n447 585
R393 B.n446 B.n23 585
R394 B.n445 B.n444 585
R395 B.n443 B.n24 585
R396 B.n442 B.n441 585
R397 B.n440 B.n25 585
R398 B.n511 B.n510 585
R399 B.n203 B.n112 526.135
R400 B.n438 B.n25 526.135
R401 B.n251 B.n250 526.135
R402 B.n394 B.n393 526.135
R403 B.n99 B.t5 300.257
R404 B.n39 B.t10 300.257
R405 B.n105 B.t2 300.255
R406 B.n32 B.t7 300.255
R407 B.n100 B.t4 249.056
R408 B.n40 B.t11 249.056
R409 B.n106 B.t1 249.055
R410 B.n33 B.t8 249.055
R411 B.n99 B.t3 222.169
R412 B.n105 B.t0 222.169
R413 B.n32 B.t6 222.169
R414 B.n39 B.t9 222.169
R415 B.n203 B.n202 163.367
R416 B.n202 B.n201 163.367
R417 B.n201 B.n114 163.367
R418 B.n197 B.n114 163.367
R419 B.n197 B.n196 163.367
R420 B.n196 B.n195 163.367
R421 B.n195 B.n116 163.367
R422 B.n191 B.n116 163.367
R423 B.n191 B.n190 163.367
R424 B.n190 B.n189 163.367
R425 B.n189 B.n118 163.367
R426 B.n185 B.n118 163.367
R427 B.n185 B.n184 163.367
R428 B.n184 B.n183 163.367
R429 B.n183 B.n120 163.367
R430 B.n179 B.n120 163.367
R431 B.n179 B.n178 163.367
R432 B.n178 B.n177 163.367
R433 B.n177 B.n122 163.367
R434 B.n173 B.n122 163.367
R435 B.n173 B.n172 163.367
R436 B.n172 B.n171 163.367
R437 B.n171 B.n124 163.367
R438 B.n167 B.n124 163.367
R439 B.n167 B.n166 163.367
R440 B.n166 B.n165 163.367
R441 B.n165 B.n126 163.367
R442 B.n161 B.n126 163.367
R443 B.n161 B.n160 163.367
R444 B.n160 B.n159 163.367
R445 B.n159 B.n128 163.367
R446 B.n155 B.n128 163.367
R447 B.n155 B.n154 163.367
R448 B.n154 B.n153 163.367
R449 B.n153 B.n130 163.367
R450 B.n149 B.n130 163.367
R451 B.n149 B.n148 163.367
R452 B.n148 B.n147 163.367
R453 B.n147 B.n132 163.367
R454 B.n143 B.n132 163.367
R455 B.n143 B.n142 163.367
R456 B.n142 B.n141 163.367
R457 B.n141 B.n134 163.367
R458 B.n137 B.n134 163.367
R459 B.n137 B.n136 163.367
R460 B.n136 B.n2 163.367
R461 B.n510 B.n2 163.367
R462 B.n510 B.n509 163.367
R463 B.n509 B.n508 163.367
R464 B.n508 B.n3 163.367
R465 B.n504 B.n3 163.367
R466 B.n504 B.n503 163.367
R467 B.n503 B.n502 163.367
R468 B.n502 B.n5 163.367
R469 B.n498 B.n5 163.367
R470 B.n498 B.n497 163.367
R471 B.n497 B.n496 163.367
R472 B.n496 B.n7 163.367
R473 B.n492 B.n7 163.367
R474 B.n492 B.n491 163.367
R475 B.n491 B.n490 163.367
R476 B.n490 B.n9 163.367
R477 B.n486 B.n9 163.367
R478 B.n486 B.n485 163.367
R479 B.n485 B.n484 163.367
R480 B.n484 B.n11 163.367
R481 B.n480 B.n11 163.367
R482 B.n480 B.n479 163.367
R483 B.n479 B.n478 163.367
R484 B.n478 B.n13 163.367
R485 B.n474 B.n13 163.367
R486 B.n474 B.n473 163.367
R487 B.n473 B.n472 163.367
R488 B.n472 B.n15 163.367
R489 B.n468 B.n15 163.367
R490 B.n468 B.n467 163.367
R491 B.n467 B.n466 163.367
R492 B.n466 B.n17 163.367
R493 B.n462 B.n17 163.367
R494 B.n462 B.n461 163.367
R495 B.n461 B.n460 163.367
R496 B.n460 B.n19 163.367
R497 B.n456 B.n19 163.367
R498 B.n456 B.n455 163.367
R499 B.n455 B.n454 163.367
R500 B.n454 B.n21 163.367
R501 B.n450 B.n21 163.367
R502 B.n450 B.n449 163.367
R503 B.n449 B.n448 163.367
R504 B.n448 B.n23 163.367
R505 B.n444 B.n23 163.367
R506 B.n444 B.n443 163.367
R507 B.n443 B.n442 163.367
R508 B.n442 B.n25 163.367
R509 B.n207 B.n112 163.367
R510 B.n208 B.n207 163.367
R511 B.n209 B.n208 163.367
R512 B.n209 B.n110 163.367
R513 B.n213 B.n110 163.367
R514 B.n214 B.n213 163.367
R515 B.n215 B.n214 163.367
R516 B.n215 B.n108 163.367
R517 B.n219 B.n108 163.367
R518 B.n220 B.n219 163.367
R519 B.n220 B.n104 163.367
R520 B.n224 B.n104 163.367
R521 B.n225 B.n224 163.367
R522 B.n226 B.n225 163.367
R523 B.n226 B.n102 163.367
R524 B.n230 B.n102 163.367
R525 B.n231 B.n230 163.367
R526 B.n232 B.n231 163.367
R527 B.n232 B.n98 163.367
R528 B.n237 B.n98 163.367
R529 B.n238 B.n237 163.367
R530 B.n239 B.n238 163.367
R531 B.n239 B.n96 163.367
R532 B.n243 B.n96 163.367
R533 B.n244 B.n243 163.367
R534 B.n245 B.n244 163.367
R535 B.n245 B.n94 163.367
R536 B.n249 B.n94 163.367
R537 B.n250 B.n249 163.367
R538 B.n251 B.n92 163.367
R539 B.n255 B.n92 163.367
R540 B.n256 B.n255 163.367
R541 B.n257 B.n256 163.367
R542 B.n257 B.n90 163.367
R543 B.n261 B.n90 163.367
R544 B.n262 B.n261 163.367
R545 B.n263 B.n262 163.367
R546 B.n263 B.n88 163.367
R547 B.n267 B.n88 163.367
R548 B.n268 B.n267 163.367
R549 B.n269 B.n268 163.367
R550 B.n269 B.n86 163.367
R551 B.n273 B.n86 163.367
R552 B.n274 B.n273 163.367
R553 B.n275 B.n274 163.367
R554 B.n275 B.n84 163.367
R555 B.n279 B.n84 163.367
R556 B.n280 B.n279 163.367
R557 B.n281 B.n280 163.367
R558 B.n281 B.n82 163.367
R559 B.n285 B.n82 163.367
R560 B.n286 B.n285 163.367
R561 B.n287 B.n286 163.367
R562 B.n287 B.n80 163.367
R563 B.n291 B.n80 163.367
R564 B.n292 B.n291 163.367
R565 B.n293 B.n292 163.367
R566 B.n293 B.n78 163.367
R567 B.n297 B.n78 163.367
R568 B.n298 B.n297 163.367
R569 B.n299 B.n298 163.367
R570 B.n299 B.n76 163.367
R571 B.n303 B.n76 163.367
R572 B.n304 B.n303 163.367
R573 B.n305 B.n304 163.367
R574 B.n305 B.n74 163.367
R575 B.n309 B.n74 163.367
R576 B.n310 B.n309 163.367
R577 B.n311 B.n310 163.367
R578 B.n311 B.n72 163.367
R579 B.n315 B.n72 163.367
R580 B.n316 B.n315 163.367
R581 B.n317 B.n316 163.367
R582 B.n317 B.n70 163.367
R583 B.n321 B.n70 163.367
R584 B.n322 B.n321 163.367
R585 B.n323 B.n322 163.367
R586 B.n323 B.n68 163.367
R587 B.n327 B.n68 163.367
R588 B.n328 B.n327 163.367
R589 B.n329 B.n328 163.367
R590 B.n329 B.n66 163.367
R591 B.n333 B.n66 163.367
R592 B.n334 B.n333 163.367
R593 B.n335 B.n334 163.367
R594 B.n335 B.n64 163.367
R595 B.n339 B.n64 163.367
R596 B.n340 B.n339 163.367
R597 B.n341 B.n340 163.367
R598 B.n341 B.n62 163.367
R599 B.n345 B.n62 163.367
R600 B.n346 B.n345 163.367
R601 B.n347 B.n346 163.367
R602 B.n347 B.n60 163.367
R603 B.n351 B.n60 163.367
R604 B.n352 B.n351 163.367
R605 B.n353 B.n352 163.367
R606 B.n353 B.n58 163.367
R607 B.n357 B.n58 163.367
R608 B.n358 B.n357 163.367
R609 B.n359 B.n358 163.367
R610 B.n359 B.n56 163.367
R611 B.n363 B.n56 163.367
R612 B.n364 B.n363 163.367
R613 B.n365 B.n364 163.367
R614 B.n365 B.n54 163.367
R615 B.n369 B.n54 163.367
R616 B.n370 B.n369 163.367
R617 B.n371 B.n370 163.367
R618 B.n371 B.n52 163.367
R619 B.n375 B.n52 163.367
R620 B.n376 B.n375 163.367
R621 B.n377 B.n376 163.367
R622 B.n377 B.n50 163.367
R623 B.n381 B.n50 163.367
R624 B.n382 B.n381 163.367
R625 B.n383 B.n382 163.367
R626 B.n383 B.n48 163.367
R627 B.n387 B.n48 163.367
R628 B.n388 B.n387 163.367
R629 B.n389 B.n388 163.367
R630 B.n389 B.n46 163.367
R631 B.n393 B.n46 163.367
R632 B.n438 B.n437 163.367
R633 B.n437 B.n436 163.367
R634 B.n436 B.n27 163.367
R635 B.n432 B.n27 163.367
R636 B.n432 B.n431 163.367
R637 B.n431 B.n430 163.367
R638 B.n430 B.n29 163.367
R639 B.n426 B.n29 163.367
R640 B.n426 B.n425 163.367
R641 B.n425 B.n424 163.367
R642 B.n424 B.n31 163.367
R643 B.n420 B.n31 163.367
R644 B.n420 B.n419 163.367
R645 B.n419 B.n418 163.367
R646 B.n418 B.n36 163.367
R647 B.n414 B.n36 163.367
R648 B.n414 B.n413 163.367
R649 B.n413 B.n412 163.367
R650 B.n412 B.n38 163.367
R651 B.n407 B.n38 163.367
R652 B.n407 B.n406 163.367
R653 B.n406 B.n405 163.367
R654 B.n405 B.n42 163.367
R655 B.n401 B.n42 163.367
R656 B.n401 B.n400 163.367
R657 B.n400 B.n399 163.367
R658 B.n399 B.n44 163.367
R659 B.n395 B.n44 163.367
R660 B.n395 B.n394 163.367
R661 B.n235 B.n100 59.5399
R662 B.n107 B.n106 59.5399
R663 B.n34 B.n33 59.5399
R664 B.n409 B.n40 59.5399
R665 B.n100 B.n99 51.2005
R666 B.n106 B.n105 51.2005
R667 B.n33 B.n32 51.2005
R668 B.n40 B.n39 51.2005
R669 B.n440 B.n439 34.1859
R670 B.n392 B.n45 34.1859
R671 B.n252 B.n93 34.1859
R672 B.n205 B.n204 34.1859
R673 B B.n511 18.0485
R674 B.n439 B.n26 10.6151
R675 B.n435 B.n26 10.6151
R676 B.n435 B.n434 10.6151
R677 B.n434 B.n433 10.6151
R678 B.n433 B.n28 10.6151
R679 B.n429 B.n28 10.6151
R680 B.n429 B.n428 10.6151
R681 B.n428 B.n427 10.6151
R682 B.n427 B.n30 10.6151
R683 B.n423 B.n422 10.6151
R684 B.n422 B.n421 10.6151
R685 B.n421 B.n35 10.6151
R686 B.n417 B.n35 10.6151
R687 B.n417 B.n416 10.6151
R688 B.n416 B.n415 10.6151
R689 B.n415 B.n37 10.6151
R690 B.n411 B.n37 10.6151
R691 B.n411 B.n410 10.6151
R692 B.n408 B.n41 10.6151
R693 B.n404 B.n41 10.6151
R694 B.n404 B.n403 10.6151
R695 B.n403 B.n402 10.6151
R696 B.n402 B.n43 10.6151
R697 B.n398 B.n43 10.6151
R698 B.n398 B.n397 10.6151
R699 B.n397 B.n396 10.6151
R700 B.n396 B.n45 10.6151
R701 B.n253 B.n252 10.6151
R702 B.n254 B.n253 10.6151
R703 B.n254 B.n91 10.6151
R704 B.n258 B.n91 10.6151
R705 B.n259 B.n258 10.6151
R706 B.n260 B.n259 10.6151
R707 B.n260 B.n89 10.6151
R708 B.n264 B.n89 10.6151
R709 B.n265 B.n264 10.6151
R710 B.n266 B.n265 10.6151
R711 B.n266 B.n87 10.6151
R712 B.n270 B.n87 10.6151
R713 B.n271 B.n270 10.6151
R714 B.n272 B.n271 10.6151
R715 B.n272 B.n85 10.6151
R716 B.n276 B.n85 10.6151
R717 B.n277 B.n276 10.6151
R718 B.n278 B.n277 10.6151
R719 B.n278 B.n83 10.6151
R720 B.n282 B.n83 10.6151
R721 B.n283 B.n282 10.6151
R722 B.n284 B.n283 10.6151
R723 B.n284 B.n81 10.6151
R724 B.n288 B.n81 10.6151
R725 B.n289 B.n288 10.6151
R726 B.n290 B.n289 10.6151
R727 B.n290 B.n79 10.6151
R728 B.n294 B.n79 10.6151
R729 B.n295 B.n294 10.6151
R730 B.n296 B.n295 10.6151
R731 B.n296 B.n77 10.6151
R732 B.n300 B.n77 10.6151
R733 B.n301 B.n300 10.6151
R734 B.n302 B.n301 10.6151
R735 B.n302 B.n75 10.6151
R736 B.n306 B.n75 10.6151
R737 B.n307 B.n306 10.6151
R738 B.n308 B.n307 10.6151
R739 B.n308 B.n73 10.6151
R740 B.n312 B.n73 10.6151
R741 B.n313 B.n312 10.6151
R742 B.n314 B.n313 10.6151
R743 B.n314 B.n71 10.6151
R744 B.n318 B.n71 10.6151
R745 B.n319 B.n318 10.6151
R746 B.n320 B.n319 10.6151
R747 B.n320 B.n69 10.6151
R748 B.n324 B.n69 10.6151
R749 B.n325 B.n324 10.6151
R750 B.n326 B.n325 10.6151
R751 B.n326 B.n67 10.6151
R752 B.n330 B.n67 10.6151
R753 B.n331 B.n330 10.6151
R754 B.n332 B.n331 10.6151
R755 B.n332 B.n65 10.6151
R756 B.n336 B.n65 10.6151
R757 B.n337 B.n336 10.6151
R758 B.n338 B.n337 10.6151
R759 B.n338 B.n63 10.6151
R760 B.n342 B.n63 10.6151
R761 B.n343 B.n342 10.6151
R762 B.n344 B.n343 10.6151
R763 B.n344 B.n61 10.6151
R764 B.n348 B.n61 10.6151
R765 B.n349 B.n348 10.6151
R766 B.n350 B.n349 10.6151
R767 B.n350 B.n59 10.6151
R768 B.n354 B.n59 10.6151
R769 B.n355 B.n354 10.6151
R770 B.n356 B.n355 10.6151
R771 B.n356 B.n57 10.6151
R772 B.n360 B.n57 10.6151
R773 B.n361 B.n360 10.6151
R774 B.n362 B.n361 10.6151
R775 B.n362 B.n55 10.6151
R776 B.n366 B.n55 10.6151
R777 B.n367 B.n366 10.6151
R778 B.n368 B.n367 10.6151
R779 B.n368 B.n53 10.6151
R780 B.n372 B.n53 10.6151
R781 B.n373 B.n372 10.6151
R782 B.n374 B.n373 10.6151
R783 B.n374 B.n51 10.6151
R784 B.n378 B.n51 10.6151
R785 B.n379 B.n378 10.6151
R786 B.n380 B.n379 10.6151
R787 B.n380 B.n49 10.6151
R788 B.n384 B.n49 10.6151
R789 B.n385 B.n384 10.6151
R790 B.n386 B.n385 10.6151
R791 B.n386 B.n47 10.6151
R792 B.n390 B.n47 10.6151
R793 B.n391 B.n390 10.6151
R794 B.n392 B.n391 10.6151
R795 B.n206 B.n205 10.6151
R796 B.n206 B.n111 10.6151
R797 B.n210 B.n111 10.6151
R798 B.n211 B.n210 10.6151
R799 B.n212 B.n211 10.6151
R800 B.n212 B.n109 10.6151
R801 B.n216 B.n109 10.6151
R802 B.n217 B.n216 10.6151
R803 B.n218 B.n217 10.6151
R804 B.n222 B.n221 10.6151
R805 B.n223 B.n222 10.6151
R806 B.n223 B.n103 10.6151
R807 B.n227 B.n103 10.6151
R808 B.n228 B.n227 10.6151
R809 B.n229 B.n228 10.6151
R810 B.n229 B.n101 10.6151
R811 B.n233 B.n101 10.6151
R812 B.n234 B.n233 10.6151
R813 B.n236 B.n97 10.6151
R814 B.n240 B.n97 10.6151
R815 B.n241 B.n240 10.6151
R816 B.n242 B.n241 10.6151
R817 B.n242 B.n95 10.6151
R818 B.n246 B.n95 10.6151
R819 B.n247 B.n246 10.6151
R820 B.n248 B.n247 10.6151
R821 B.n248 B.n93 10.6151
R822 B.n204 B.n113 10.6151
R823 B.n200 B.n113 10.6151
R824 B.n200 B.n199 10.6151
R825 B.n199 B.n198 10.6151
R826 B.n198 B.n115 10.6151
R827 B.n194 B.n115 10.6151
R828 B.n194 B.n193 10.6151
R829 B.n193 B.n192 10.6151
R830 B.n192 B.n117 10.6151
R831 B.n188 B.n117 10.6151
R832 B.n188 B.n187 10.6151
R833 B.n187 B.n186 10.6151
R834 B.n186 B.n119 10.6151
R835 B.n182 B.n119 10.6151
R836 B.n182 B.n181 10.6151
R837 B.n181 B.n180 10.6151
R838 B.n180 B.n121 10.6151
R839 B.n176 B.n121 10.6151
R840 B.n176 B.n175 10.6151
R841 B.n175 B.n174 10.6151
R842 B.n174 B.n123 10.6151
R843 B.n170 B.n123 10.6151
R844 B.n170 B.n169 10.6151
R845 B.n169 B.n168 10.6151
R846 B.n168 B.n125 10.6151
R847 B.n164 B.n125 10.6151
R848 B.n164 B.n163 10.6151
R849 B.n163 B.n162 10.6151
R850 B.n162 B.n127 10.6151
R851 B.n158 B.n127 10.6151
R852 B.n158 B.n157 10.6151
R853 B.n157 B.n156 10.6151
R854 B.n156 B.n129 10.6151
R855 B.n152 B.n129 10.6151
R856 B.n152 B.n151 10.6151
R857 B.n151 B.n150 10.6151
R858 B.n150 B.n131 10.6151
R859 B.n146 B.n131 10.6151
R860 B.n146 B.n145 10.6151
R861 B.n145 B.n144 10.6151
R862 B.n144 B.n133 10.6151
R863 B.n140 B.n133 10.6151
R864 B.n140 B.n139 10.6151
R865 B.n139 B.n138 10.6151
R866 B.n138 B.n135 10.6151
R867 B.n135 B.n0 10.6151
R868 B.n507 B.n1 10.6151
R869 B.n507 B.n506 10.6151
R870 B.n506 B.n505 10.6151
R871 B.n505 B.n4 10.6151
R872 B.n501 B.n4 10.6151
R873 B.n501 B.n500 10.6151
R874 B.n500 B.n499 10.6151
R875 B.n499 B.n6 10.6151
R876 B.n495 B.n6 10.6151
R877 B.n495 B.n494 10.6151
R878 B.n494 B.n493 10.6151
R879 B.n493 B.n8 10.6151
R880 B.n489 B.n8 10.6151
R881 B.n489 B.n488 10.6151
R882 B.n488 B.n487 10.6151
R883 B.n487 B.n10 10.6151
R884 B.n483 B.n10 10.6151
R885 B.n483 B.n482 10.6151
R886 B.n482 B.n481 10.6151
R887 B.n481 B.n12 10.6151
R888 B.n477 B.n12 10.6151
R889 B.n477 B.n476 10.6151
R890 B.n476 B.n475 10.6151
R891 B.n475 B.n14 10.6151
R892 B.n471 B.n14 10.6151
R893 B.n471 B.n470 10.6151
R894 B.n470 B.n469 10.6151
R895 B.n469 B.n16 10.6151
R896 B.n465 B.n16 10.6151
R897 B.n465 B.n464 10.6151
R898 B.n464 B.n463 10.6151
R899 B.n463 B.n18 10.6151
R900 B.n459 B.n18 10.6151
R901 B.n459 B.n458 10.6151
R902 B.n458 B.n457 10.6151
R903 B.n457 B.n20 10.6151
R904 B.n453 B.n20 10.6151
R905 B.n453 B.n452 10.6151
R906 B.n452 B.n451 10.6151
R907 B.n451 B.n22 10.6151
R908 B.n447 B.n22 10.6151
R909 B.n447 B.n446 10.6151
R910 B.n446 B.n445 10.6151
R911 B.n445 B.n24 10.6151
R912 B.n441 B.n24 10.6151
R913 B.n441 B.n440 10.6151
R914 B.n34 B.n30 9.36635
R915 B.n409 B.n408 9.36635
R916 B.n218 B.n107 9.36635
R917 B.n236 B.n235 9.36635
R918 B.n511 B.n0 2.81026
R919 B.n511 B.n1 2.81026
R920 B.n423 B.n34 1.24928
R921 B.n410 B.n409 1.24928
R922 B.n221 B.n107 1.24928
R923 B.n235 B.n234 1.24928
R924 VN.n51 VN.n27 161.3
R925 VN.n50 VN.n49 161.3
R926 VN.n48 VN.n28 161.3
R927 VN.n47 VN.n46 161.3
R928 VN.n45 VN.n29 161.3
R929 VN.n43 VN.n42 161.3
R930 VN.n41 VN.n30 161.3
R931 VN.n40 VN.n39 161.3
R932 VN.n38 VN.n31 161.3
R933 VN.n37 VN.n36 161.3
R934 VN.n35 VN.n32 161.3
R935 VN.n24 VN.n0 161.3
R936 VN.n23 VN.n22 161.3
R937 VN.n21 VN.n1 161.3
R938 VN.n20 VN.n19 161.3
R939 VN.n18 VN.n2 161.3
R940 VN.n16 VN.n15 161.3
R941 VN.n14 VN.n3 161.3
R942 VN.n13 VN.n12 161.3
R943 VN.n11 VN.n4 161.3
R944 VN.n10 VN.n9 161.3
R945 VN.n8 VN.n5 161.3
R946 VN.n26 VN.n25 100.579
R947 VN.n53 VN.n52 100.579
R948 VN.n7 VN.n6 68.9827
R949 VN.n34 VN.n33 68.9827
R950 VN.n12 VN.n11 56.5617
R951 VN.n39 VN.n38 56.5617
R952 VN.n19 VN.n1 51.2335
R953 VN.n46 VN.n28 51.2335
R954 VN.n7 VN.t0 45.6612
R955 VN.n34 VN.t2 45.6612
R956 VN VN.n53 41.7406
R957 VN.n23 VN.n1 29.9206
R958 VN.n50 VN.n28 29.9206
R959 VN.n10 VN.n5 24.5923
R960 VN.n11 VN.n10 24.5923
R961 VN.n12 VN.n3 24.5923
R962 VN.n16 VN.n3 24.5923
R963 VN.n19 VN.n18 24.5923
R964 VN.n24 VN.n23 24.5923
R965 VN.n38 VN.n37 24.5923
R966 VN.n37 VN.n32 24.5923
R967 VN.n46 VN.n45 24.5923
R968 VN.n43 VN.n30 24.5923
R969 VN.n39 VN.n30 24.5923
R970 VN.n51 VN.n50 24.5923
R971 VN.n18 VN.n17 21.1495
R972 VN.n45 VN.n44 21.1495
R973 VN.n6 VN.t4 14.6066
R974 VN.n17 VN.t6 14.6066
R975 VN.n25 VN.t3 14.6066
R976 VN.n33 VN.t5 14.6066
R977 VN.n44 VN.t1 14.6066
R978 VN.n52 VN.t7 14.6066
R979 VN.n25 VN.n24 10.3291
R980 VN.n52 VN.n51 10.3291
R981 VN.n35 VN.n34 9.96756
R982 VN.n8 VN.n7 9.96756
R983 VN.n6 VN.n5 3.44336
R984 VN.n17 VN.n16 3.44336
R985 VN.n33 VN.n32 3.44336
R986 VN.n44 VN.n43 3.44336
R987 VN.n53 VN.n27 0.278335
R988 VN.n26 VN.n0 0.278335
R989 VN.n49 VN.n27 0.189894
R990 VN.n49 VN.n48 0.189894
R991 VN.n48 VN.n47 0.189894
R992 VN.n47 VN.n29 0.189894
R993 VN.n42 VN.n29 0.189894
R994 VN.n42 VN.n41 0.189894
R995 VN.n41 VN.n40 0.189894
R996 VN.n40 VN.n31 0.189894
R997 VN.n36 VN.n31 0.189894
R998 VN.n36 VN.n35 0.189894
R999 VN.n9 VN.n8 0.189894
R1000 VN.n9 VN.n4 0.189894
R1001 VN.n13 VN.n4 0.189894
R1002 VN.n14 VN.n13 0.189894
R1003 VN.n15 VN.n14 0.189894
R1004 VN.n15 VN.n2 0.189894
R1005 VN.n20 VN.n2 0.189894
R1006 VN.n21 VN.n20 0.189894
R1007 VN.n22 VN.n21 0.189894
R1008 VN.n22 VN.n0 0.189894
R1009 VN VN.n26 0.153485
R1010 VDD2.n2 VDD2.n1 250.095
R1011 VDD2.n2 VDD2.n0 250.095
R1012 VDD2 VDD2.n5 250.093
R1013 VDD2.n4 VDD2.n3 249.013
R1014 VDD2.n4 VDD2.n2 35.1636
R1015 VDD2.n5 VDD2.t2 23.2184
R1016 VDD2.n5 VDD2.t5 23.2184
R1017 VDD2.n3 VDD2.t0 23.2184
R1018 VDD2.n3 VDD2.t6 23.2184
R1019 VDD2.n1 VDD2.t1 23.2184
R1020 VDD2.n1 VDD2.t4 23.2184
R1021 VDD2.n0 VDD2.t7 23.2184
R1022 VDD2.n0 VDD2.t3 23.2184
R1023 VDD2 VDD2.n4 1.19662
C0 w_n3610_n1248# VDD2 1.66944f
C1 B VP 1.80252f
C2 w_n3610_n1248# VP 7.53733f
C3 w_n3610_n1248# B 6.75015f
C4 VN VDD2 1.38939f
C5 VP VN 5.35114f
C6 B VN 1.0209f
C7 w_n3610_n1248# VN 7.076f
C8 VDD1 VDD2 1.62566f
C9 VDD2 VTAIL 4.29652f
C10 VP VDD1 1.72541f
C11 B VDD1 1.27552f
C12 VP VTAIL 2.46849f
C13 B VTAIL 1.30898f
C14 w_n3610_n1248# VDD1 1.56781f
C15 w_n3610_n1248# VTAIL 1.72197f
C16 VDD1 VN 0.15796f
C17 VN VTAIL 2.45438f
C18 VDD1 VTAIL 4.24405f
C19 VP VDD2 0.497054f
C20 B VDD2 1.36287f
C21 VDD2 VSUBS 1.054378f
C22 VDD1 VSUBS 1.621301f
C23 VTAIL VSUBS 0.494052f
C24 VN VSUBS 6.34459f
C25 VP VSUBS 2.668111f
C26 B VSUBS 3.549615f
C27 w_n3610_n1248# VSUBS 57.8322f
C28 VDD2.t7 VSUBS 0.020233f
C29 VDD2.t3 VSUBS 0.020233f
C30 VDD2.n0 VSUBS 0.078427f
C31 VDD2.t1 VSUBS 0.020233f
C32 VDD2.t4 VSUBS 0.020233f
C33 VDD2.n1 VSUBS 0.078427f
C34 VDD2.n2 VSUBS 1.83801f
C35 VDD2.t0 VSUBS 0.020233f
C36 VDD2.t6 VSUBS 0.020233f
C37 VDD2.n3 VSUBS 0.076835f
C38 VDD2.n4 VSUBS 1.48817f
C39 VDD2.t2 VSUBS 0.020233f
C40 VDD2.t5 VSUBS 0.020233f
C41 VDD2.n5 VSUBS 0.078421f
C42 VN.n0 VSUBS 0.07293f
C43 VN.t3 VSUBS 0.382005f
C44 VN.n1 VSUBS 0.053846f
C45 VN.n2 VSUBS 0.055321f
C46 VN.t6 VSUBS 0.382005f
C47 VN.n3 VSUBS 0.102587f
C48 VN.n4 VSUBS 0.055321f
C49 VN.n5 VSUBS 0.059033f
C50 VN.t0 VSUBS 0.732997f
C51 VN.t4 VSUBS 0.382005f
C52 VN.n6 VSUBS 0.348818f
C53 VN.n7 VSUBS 0.349136f
C54 VN.n8 VSUBS 0.47634f
C55 VN.n9 VSUBS 0.055321f
C56 VN.n10 VSUBS 0.102587f
C57 VN.n11 VSUBS 0.080417f
C58 VN.n12 VSUBS 0.080417f
C59 VN.n13 VSUBS 0.055321f
C60 VN.n14 VSUBS 0.055321f
C61 VN.n15 VSUBS 0.055321f
C62 VN.n16 VSUBS 0.059033f
C63 VN.n17 VSUBS 0.217772f
C64 VN.n18 VSUBS 0.095497f
C65 VN.n19 VSUBS 0.099954f
C66 VN.n20 VSUBS 0.055321f
C67 VN.n21 VSUBS 0.055321f
C68 VN.n22 VSUBS 0.055321f
C69 VN.n23 VSUBS 0.109622f
C70 VN.n24 VSUBS 0.073213f
C71 VN.n25 VSUBS 0.381297f
C72 VN.n26 VSUBS 0.084629f
C73 VN.n27 VSUBS 0.07293f
C74 VN.t7 VSUBS 0.382005f
C75 VN.n28 VSUBS 0.053846f
C76 VN.n29 VSUBS 0.055321f
C77 VN.t1 VSUBS 0.382005f
C78 VN.n30 VSUBS 0.102587f
C79 VN.n31 VSUBS 0.055321f
C80 VN.n32 VSUBS 0.059033f
C81 VN.t2 VSUBS 0.732997f
C82 VN.t5 VSUBS 0.382005f
C83 VN.n33 VSUBS 0.348818f
C84 VN.n34 VSUBS 0.349136f
C85 VN.n35 VSUBS 0.47634f
C86 VN.n36 VSUBS 0.055321f
C87 VN.n37 VSUBS 0.102587f
C88 VN.n38 VSUBS 0.080417f
C89 VN.n39 VSUBS 0.080417f
C90 VN.n40 VSUBS 0.055321f
C91 VN.n41 VSUBS 0.055321f
C92 VN.n42 VSUBS 0.055321f
C93 VN.n43 VSUBS 0.059033f
C94 VN.n44 VSUBS 0.217772f
C95 VN.n45 VSUBS 0.095497f
C96 VN.n46 VSUBS 0.099954f
C97 VN.n47 VSUBS 0.055321f
C98 VN.n48 VSUBS 0.055321f
C99 VN.n49 VSUBS 0.055321f
C100 VN.n50 VSUBS 0.109622f
C101 VN.n51 VSUBS 0.073213f
C102 VN.n52 VSUBS 0.381297f
C103 VN.n53 VSUBS 2.32837f
C104 B.n0 VSUBS 0.005939f
C105 B.n1 VSUBS 0.005939f
C106 B.n2 VSUBS 0.009392f
C107 B.n3 VSUBS 0.009392f
C108 B.n4 VSUBS 0.009392f
C109 B.n5 VSUBS 0.009392f
C110 B.n6 VSUBS 0.009392f
C111 B.n7 VSUBS 0.009392f
C112 B.n8 VSUBS 0.009392f
C113 B.n9 VSUBS 0.009392f
C114 B.n10 VSUBS 0.009392f
C115 B.n11 VSUBS 0.009392f
C116 B.n12 VSUBS 0.009392f
C117 B.n13 VSUBS 0.009392f
C118 B.n14 VSUBS 0.009392f
C119 B.n15 VSUBS 0.009392f
C120 B.n16 VSUBS 0.009392f
C121 B.n17 VSUBS 0.009392f
C122 B.n18 VSUBS 0.009392f
C123 B.n19 VSUBS 0.009392f
C124 B.n20 VSUBS 0.009392f
C125 B.n21 VSUBS 0.009392f
C126 B.n22 VSUBS 0.009392f
C127 B.n23 VSUBS 0.009392f
C128 B.n24 VSUBS 0.009392f
C129 B.n25 VSUBS 0.022407f
C130 B.n26 VSUBS 0.009392f
C131 B.n27 VSUBS 0.009392f
C132 B.n28 VSUBS 0.009392f
C133 B.n29 VSUBS 0.009392f
C134 B.n30 VSUBS 0.00884f
C135 B.n31 VSUBS 0.009392f
C136 B.t8 VSUBS 0.037798f
C137 B.t7 VSUBS 0.047009f
C138 B.t6 VSUBS 0.216122f
C139 B.n32 VSUBS 0.083275f
C140 B.n33 VSUBS 0.067418f
C141 B.n34 VSUBS 0.021761f
C142 B.n35 VSUBS 0.009392f
C143 B.n36 VSUBS 0.009392f
C144 B.n37 VSUBS 0.009392f
C145 B.n38 VSUBS 0.009392f
C146 B.t11 VSUBS 0.037798f
C147 B.t10 VSUBS 0.047009f
C148 B.t9 VSUBS 0.216122f
C149 B.n39 VSUBS 0.083275f
C150 B.n40 VSUBS 0.067418f
C151 B.n41 VSUBS 0.009392f
C152 B.n42 VSUBS 0.009392f
C153 B.n43 VSUBS 0.009392f
C154 B.n44 VSUBS 0.009392f
C155 B.n45 VSUBS 0.021838f
C156 B.n46 VSUBS 0.009392f
C157 B.n47 VSUBS 0.009392f
C158 B.n48 VSUBS 0.009392f
C159 B.n49 VSUBS 0.009392f
C160 B.n50 VSUBS 0.009392f
C161 B.n51 VSUBS 0.009392f
C162 B.n52 VSUBS 0.009392f
C163 B.n53 VSUBS 0.009392f
C164 B.n54 VSUBS 0.009392f
C165 B.n55 VSUBS 0.009392f
C166 B.n56 VSUBS 0.009392f
C167 B.n57 VSUBS 0.009392f
C168 B.n58 VSUBS 0.009392f
C169 B.n59 VSUBS 0.009392f
C170 B.n60 VSUBS 0.009392f
C171 B.n61 VSUBS 0.009392f
C172 B.n62 VSUBS 0.009392f
C173 B.n63 VSUBS 0.009392f
C174 B.n64 VSUBS 0.009392f
C175 B.n65 VSUBS 0.009392f
C176 B.n66 VSUBS 0.009392f
C177 B.n67 VSUBS 0.009392f
C178 B.n68 VSUBS 0.009392f
C179 B.n69 VSUBS 0.009392f
C180 B.n70 VSUBS 0.009392f
C181 B.n71 VSUBS 0.009392f
C182 B.n72 VSUBS 0.009392f
C183 B.n73 VSUBS 0.009392f
C184 B.n74 VSUBS 0.009392f
C185 B.n75 VSUBS 0.009392f
C186 B.n76 VSUBS 0.009392f
C187 B.n77 VSUBS 0.009392f
C188 B.n78 VSUBS 0.009392f
C189 B.n79 VSUBS 0.009392f
C190 B.n80 VSUBS 0.009392f
C191 B.n81 VSUBS 0.009392f
C192 B.n82 VSUBS 0.009392f
C193 B.n83 VSUBS 0.009392f
C194 B.n84 VSUBS 0.009392f
C195 B.n85 VSUBS 0.009392f
C196 B.n86 VSUBS 0.009392f
C197 B.n87 VSUBS 0.009392f
C198 B.n88 VSUBS 0.009392f
C199 B.n89 VSUBS 0.009392f
C200 B.n90 VSUBS 0.009392f
C201 B.n91 VSUBS 0.009392f
C202 B.n92 VSUBS 0.009392f
C203 B.n93 VSUBS 0.022898f
C204 B.n94 VSUBS 0.009392f
C205 B.n95 VSUBS 0.009392f
C206 B.n96 VSUBS 0.009392f
C207 B.n97 VSUBS 0.009392f
C208 B.n98 VSUBS 0.009392f
C209 B.t4 VSUBS 0.037798f
C210 B.t5 VSUBS 0.047009f
C211 B.t3 VSUBS 0.216122f
C212 B.n99 VSUBS 0.083275f
C213 B.n100 VSUBS 0.067418f
C214 B.n101 VSUBS 0.009392f
C215 B.n102 VSUBS 0.009392f
C216 B.n103 VSUBS 0.009392f
C217 B.n104 VSUBS 0.009392f
C218 B.t1 VSUBS 0.037798f
C219 B.t2 VSUBS 0.047009f
C220 B.t0 VSUBS 0.216122f
C221 B.n105 VSUBS 0.083275f
C222 B.n106 VSUBS 0.067418f
C223 B.n107 VSUBS 0.021761f
C224 B.n108 VSUBS 0.009392f
C225 B.n109 VSUBS 0.009392f
C226 B.n110 VSUBS 0.009392f
C227 B.n111 VSUBS 0.009392f
C228 B.n112 VSUBS 0.022898f
C229 B.n113 VSUBS 0.009392f
C230 B.n114 VSUBS 0.009392f
C231 B.n115 VSUBS 0.009392f
C232 B.n116 VSUBS 0.009392f
C233 B.n117 VSUBS 0.009392f
C234 B.n118 VSUBS 0.009392f
C235 B.n119 VSUBS 0.009392f
C236 B.n120 VSUBS 0.009392f
C237 B.n121 VSUBS 0.009392f
C238 B.n122 VSUBS 0.009392f
C239 B.n123 VSUBS 0.009392f
C240 B.n124 VSUBS 0.009392f
C241 B.n125 VSUBS 0.009392f
C242 B.n126 VSUBS 0.009392f
C243 B.n127 VSUBS 0.009392f
C244 B.n128 VSUBS 0.009392f
C245 B.n129 VSUBS 0.009392f
C246 B.n130 VSUBS 0.009392f
C247 B.n131 VSUBS 0.009392f
C248 B.n132 VSUBS 0.009392f
C249 B.n133 VSUBS 0.009392f
C250 B.n134 VSUBS 0.009392f
C251 B.n135 VSUBS 0.009392f
C252 B.n136 VSUBS 0.009392f
C253 B.n137 VSUBS 0.009392f
C254 B.n138 VSUBS 0.009392f
C255 B.n139 VSUBS 0.009392f
C256 B.n140 VSUBS 0.009392f
C257 B.n141 VSUBS 0.009392f
C258 B.n142 VSUBS 0.009392f
C259 B.n143 VSUBS 0.009392f
C260 B.n144 VSUBS 0.009392f
C261 B.n145 VSUBS 0.009392f
C262 B.n146 VSUBS 0.009392f
C263 B.n147 VSUBS 0.009392f
C264 B.n148 VSUBS 0.009392f
C265 B.n149 VSUBS 0.009392f
C266 B.n150 VSUBS 0.009392f
C267 B.n151 VSUBS 0.009392f
C268 B.n152 VSUBS 0.009392f
C269 B.n153 VSUBS 0.009392f
C270 B.n154 VSUBS 0.009392f
C271 B.n155 VSUBS 0.009392f
C272 B.n156 VSUBS 0.009392f
C273 B.n157 VSUBS 0.009392f
C274 B.n158 VSUBS 0.009392f
C275 B.n159 VSUBS 0.009392f
C276 B.n160 VSUBS 0.009392f
C277 B.n161 VSUBS 0.009392f
C278 B.n162 VSUBS 0.009392f
C279 B.n163 VSUBS 0.009392f
C280 B.n164 VSUBS 0.009392f
C281 B.n165 VSUBS 0.009392f
C282 B.n166 VSUBS 0.009392f
C283 B.n167 VSUBS 0.009392f
C284 B.n168 VSUBS 0.009392f
C285 B.n169 VSUBS 0.009392f
C286 B.n170 VSUBS 0.009392f
C287 B.n171 VSUBS 0.009392f
C288 B.n172 VSUBS 0.009392f
C289 B.n173 VSUBS 0.009392f
C290 B.n174 VSUBS 0.009392f
C291 B.n175 VSUBS 0.009392f
C292 B.n176 VSUBS 0.009392f
C293 B.n177 VSUBS 0.009392f
C294 B.n178 VSUBS 0.009392f
C295 B.n179 VSUBS 0.009392f
C296 B.n180 VSUBS 0.009392f
C297 B.n181 VSUBS 0.009392f
C298 B.n182 VSUBS 0.009392f
C299 B.n183 VSUBS 0.009392f
C300 B.n184 VSUBS 0.009392f
C301 B.n185 VSUBS 0.009392f
C302 B.n186 VSUBS 0.009392f
C303 B.n187 VSUBS 0.009392f
C304 B.n188 VSUBS 0.009392f
C305 B.n189 VSUBS 0.009392f
C306 B.n190 VSUBS 0.009392f
C307 B.n191 VSUBS 0.009392f
C308 B.n192 VSUBS 0.009392f
C309 B.n193 VSUBS 0.009392f
C310 B.n194 VSUBS 0.009392f
C311 B.n195 VSUBS 0.009392f
C312 B.n196 VSUBS 0.009392f
C313 B.n197 VSUBS 0.009392f
C314 B.n198 VSUBS 0.009392f
C315 B.n199 VSUBS 0.009392f
C316 B.n200 VSUBS 0.009392f
C317 B.n201 VSUBS 0.009392f
C318 B.n202 VSUBS 0.009392f
C319 B.n203 VSUBS 0.022407f
C320 B.n204 VSUBS 0.022407f
C321 B.n205 VSUBS 0.022898f
C322 B.n206 VSUBS 0.009392f
C323 B.n207 VSUBS 0.009392f
C324 B.n208 VSUBS 0.009392f
C325 B.n209 VSUBS 0.009392f
C326 B.n210 VSUBS 0.009392f
C327 B.n211 VSUBS 0.009392f
C328 B.n212 VSUBS 0.009392f
C329 B.n213 VSUBS 0.009392f
C330 B.n214 VSUBS 0.009392f
C331 B.n215 VSUBS 0.009392f
C332 B.n216 VSUBS 0.009392f
C333 B.n217 VSUBS 0.009392f
C334 B.n218 VSUBS 0.00884f
C335 B.n219 VSUBS 0.009392f
C336 B.n220 VSUBS 0.009392f
C337 B.n221 VSUBS 0.005249f
C338 B.n222 VSUBS 0.009392f
C339 B.n223 VSUBS 0.009392f
C340 B.n224 VSUBS 0.009392f
C341 B.n225 VSUBS 0.009392f
C342 B.n226 VSUBS 0.009392f
C343 B.n227 VSUBS 0.009392f
C344 B.n228 VSUBS 0.009392f
C345 B.n229 VSUBS 0.009392f
C346 B.n230 VSUBS 0.009392f
C347 B.n231 VSUBS 0.009392f
C348 B.n232 VSUBS 0.009392f
C349 B.n233 VSUBS 0.009392f
C350 B.n234 VSUBS 0.005249f
C351 B.n235 VSUBS 0.021761f
C352 B.n236 VSUBS 0.00884f
C353 B.n237 VSUBS 0.009392f
C354 B.n238 VSUBS 0.009392f
C355 B.n239 VSUBS 0.009392f
C356 B.n240 VSUBS 0.009392f
C357 B.n241 VSUBS 0.009392f
C358 B.n242 VSUBS 0.009392f
C359 B.n243 VSUBS 0.009392f
C360 B.n244 VSUBS 0.009392f
C361 B.n245 VSUBS 0.009392f
C362 B.n246 VSUBS 0.009392f
C363 B.n247 VSUBS 0.009392f
C364 B.n248 VSUBS 0.009392f
C365 B.n249 VSUBS 0.009392f
C366 B.n250 VSUBS 0.022898f
C367 B.n251 VSUBS 0.022407f
C368 B.n252 VSUBS 0.022407f
C369 B.n253 VSUBS 0.009392f
C370 B.n254 VSUBS 0.009392f
C371 B.n255 VSUBS 0.009392f
C372 B.n256 VSUBS 0.009392f
C373 B.n257 VSUBS 0.009392f
C374 B.n258 VSUBS 0.009392f
C375 B.n259 VSUBS 0.009392f
C376 B.n260 VSUBS 0.009392f
C377 B.n261 VSUBS 0.009392f
C378 B.n262 VSUBS 0.009392f
C379 B.n263 VSUBS 0.009392f
C380 B.n264 VSUBS 0.009392f
C381 B.n265 VSUBS 0.009392f
C382 B.n266 VSUBS 0.009392f
C383 B.n267 VSUBS 0.009392f
C384 B.n268 VSUBS 0.009392f
C385 B.n269 VSUBS 0.009392f
C386 B.n270 VSUBS 0.009392f
C387 B.n271 VSUBS 0.009392f
C388 B.n272 VSUBS 0.009392f
C389 B.n273 VSUBS 0.009392f
C390 B.n274 VSUBS 0.009392f
C391 B.n275 VSUBS 0.009392f
C392 B.n276 VSUBS 0.009392f
C393 B.n277 VSUBS 0.009392f
C394 B.n278 VSUBS 0.009392f
C395 B.n279 VSUBS 0.009392f
C396 B.n280 VSUBS 0.009392f
C397 B.n281 VSUBS 0.009392f
C398 B.n282 VSUBS 0.009392f
C399 B.n283 VSUBS 0.009392f
C400 B.n284 VSUBS 0.009392f
C401 B.n285 VSUBS 0.009392f
C402 B.n286 VSUBS 0.009392f
C403 B.n287 VSUBS 0.009392f
C404 B.n288 VSUBS 0.009392f
C405 B.n289 VSUBS 0.009392f
C406 B.n290 VSUBS 0.009392f
C407 B.n291 VSUBS 0.009392f
C408 B.n292 VSUBS 0.009392f
C409 B.n293 VSUBS 0.009392f
C410 B.n294 VSUBS 0.009392f
C411 B.n295 VSUBS 0.009392f
C412 B.n296 VSUBS 0.009392f
C413 B.n297 VSUBS 0.009392f
C414 B.n298 VSUBS 0.009392f
C415 B.n299 VSUBS 0.009392f
C416 B.n300 VSUBS 0.009392f
C417 B.n301 VSUBS 0.009392f
C418 B.n302 VSUBS 0.009392f
C419 B.n303 VSUBS 0.009392f
C420 B.n304 VSUBS 0.009392f
C421 B.n305 VSUBS 0.009392f
C422 B.n306 VSUBS 0.009392f
C423 B.n307 VSUBS 0.009392f
C424 B.n308 VSUBS 0.009392f
C425 B.n309 VSUBS 0.009392f
C426 B.n310 VSUBS 0.009392f
C427 B.n311 VSUBS 0.009392f
C428 B.n312 VSUBS 0.009392f
C429 B.n313 VSUBS 0.009392f
C430 B.n314 VSUBS 0.009392f
C431 B.n315 VSUBS 0.009392f
C432 B.n316 VSUBS 0.009392f
C433 B.n317 VSUBS 0.009392f
C434 B.n318 VSUBS 0.009392f
C435 B.n319 VSUBS 0.009392f
C436 B.n320 VSUBS 0.009392f
C437 B.n321 VSUBS 0.009392f
C438 B.n322 VSUBS 0.009392f
C439 B.n323 VSUBS 0.009392f
C440 B.n324 VSUBS 0.009392f
C441 B.n325 VSUBS 0.009392f
C442 B.n326 VSUBS 0.009392f
C443 B.n327 VSUBS 0.009392f
C444 B.n328 VSUBS 0.009392f
C445 B.n329 VSUBS 0.009392f
C446 B.n330 VSUBS 0.009392f
C447 B.n331 VSUBS 0.009392f
C448 B.n332 VSUBS 0.009392f
C449 B.n333 VSUBS 0.009392f
C450 B.n334 VSUBS 0.009392f
C451 B.n335 VSUBS 0.009392f
C452 B.n336 VSUBS 0.009392f
C453 B.n337 VSUBS 0.009392f
C454 B.n338 VSUBS 0.009392f
C455 B.n339 VSUBS 0.009392f
C456 B.n340 VSUBS 0.009392f
C457 B.n341 VSUBS 0.009392f
C458 B.n342 VSUBS 0.009392f
C459 B.n343 VSUBS 0.009392f
C460 B.n344 VSUBS 0.009392f
C461 B.n345 VSUBS 0.009392f
C462 B.n346 VSUBS 0.009392f
C463 B.n347 VSUBS 0.009392f
C464 B.n348 VSUBS 0.009392f
C465 B.n349 VSUBS 0.009392f
C466 B.n350 VSUBS 0.009392f
C467 B.n351 VSUBS 0.009392f
C468 B.n352 VSUBS 0.009392f
C469 B.n353 VSUBS 0.009392f
C470 B.n354 VSUBS 0.009392f
C471 B.n355 VSUBS 0.009392f
C472 B.n356 VSUBS 0.009392f
C473 B.n357 VSUBS 0.009392f
C474 B.n358 VSUBS 0.009392f
C475 B.n359 VSUBS 0.009392f
C476 B.n360 VSUBS 0.009392f
C477 B.n361 VSUBS 0.009392f
C478 B.n362 VSUBS 0.009392f
C479 B.n363 VSUBS 0.009392f
C480 B.n364 VSUBS 0.009392f
C481 B.n365 VSUBS 0.009392f
C482 B.n366 VSUBS 0.009392f
C483 B.n367 VSUBS 0.009392f
C484 B.n368 VSUBS 0.009392f
C485 B.n369 VSUBS 0.009392f
C486 B.n370 VSUBS 0.009392f
C487 B.n371 VSUBS 0.009392f
C488 B.n372 VSUBS 0.009392f
C489 B.n373 VSUBS 0.009392f
C490 B.n374 VSUBS 0.009392f
C491 B.n375 VSUBS 0.009392f
C492 B.n376 VSUBS 0.009392f
C493 B.n377 VSUBS 0.009392f
C494 B.n378 VSUBS 0.009392f
C495 B.n379 VSUBS 0.009392f
C496 B.n380 VSUBS 0.009392f
C497 B.n381 VSUBS 0.009392f
C498 B.n382 VSUBS 0.009392f
C499 B.n383 VSUBS 0.009392f
C500 B.n384 VSUBS 0.009392f
C501 B.n385 VSUBS 0.009392f
C502 B.n386 VSUBS 0.009392f
C503 B.n387 VSUBS 0.009392f
C504 B.n388 VSUBS 0.009392f
C505 B.n389 VSUBS 0.009392f
C506 B.n390 VSUBS 0.009392f
C507 B.n391 VSUBS 0.009392f
C508 B.n392 VSUBS 0.023467f
C509 B.n393 VSUBS 0.022407f
C510 B.n394 VSUBS 0.022898f
C511 B.n395 VSUBS 0.009392f
C512 B.n396 VSUBS 0.009392f
C513 B.n397 VSUBS 0.009392f
C514 B.n398 VSUBS 0.009392f
C515 B.n399 VSUBS 0.009392f
C516 B.n400 VSUBS 0.009392f
C517 B.n401 VSUBS 0.009392f
C518 B.n402 VSUBS 0.009392f
C519 B.n403 VSUBS 0.009392f
C520 B.n404 VSUBS 0.009392f
C521 B.n405 VSUBS 0.009392f
C522 B.n406 VSUBS 0.009392f
C523 B.n407 VSUBS 0.009392f
C524 B.n408 VSUBS 0.00884f
C525 B.n409 VSUBS 0.021761f
C526 B.n410 VSUBS 0.005249f
C527 B.n411 VSUBS 0.009392f
C528 B.n412 VSUBS 0.009392f
C529 B.n413 VSUBS 0.009392f
C530 B.n414 VSUBS 0.009392f
C531 B.n415 VSUBS 0.009392f
C532 B.n416 VSUBS 0.009392f
C533 B.n417 VSUBS 0.009392f
C534 B.n418 VSUBS 0.009392f
C535 B.n419 VSUBS 0.009392f
C536 B.n420 VSUBS 0.009392f
C537 B.n421 VSUBS 0.009392f
C538 B.n422 VSUBS 0.009392f
C539 B.n423 VSUBS 0.005249f
C540 B.n424 VSUBS 0.009392f
C541 B.n425 VSUBS 0.009392f
C542 B.n426 VSUBS 0.009392f
C543 B.n427 VSUBS 0.009392f
C544 B.n428 VSUBS 0.009392f
C545 B.n429 VSUBS 0.009392f
C546 B.n430 VSUBS 0.009392f
C547 B.n431 VSUBS 0.009392f
C548 B.n432 VSUBS 0.009392f
C549 B.n433 VSUBS 0.009392f
C550 B.n434 VSUBS 0.009392f
C551 B.n435 VSUBS 0.009392f
C552 B.n436 VSUBS 0.009392f
C553 B.n437 VSUBS 0.009392f
C554 B.n438 VSUBS 0.022898f
C555 B.n439 VSUBS 0.022898f
C556 B.n440 VSUBS 0.022407f
C557 B.n441 VSUBS 0.009392f
C558 B.n442 VSUBS 0.009392f
C559 B.n443 VSUBS 0.009392f
C560 B.n444 VSUBS 0.009392f
C561 B.n445 VSUBS 0.009392f
C562 B.n446 VSUBS 0.009392f
C563 B.n447 VSUBS 0.009392f
C564 B.n448 VSUBS 0.009392f
C565 B.n449 VSUBS 0.009392f
C566 B.n450 VSUBS 0.009392f
C567 B.n451 VSUBS 0.009392f
C568 B.n452 VSUBS 0.009392f
C569 B.n453 VSUBS 0.009392f
C570 B.n454 VSUBS 0.009392f
C571 B.n455 VSUBS 0.009392f
C572 B.n456 VSUBS 0.009392f
C573 B.n457 VSUBS 0.009392f
C574 B.n458 VSUBS 0.009392f
C575 B.n459 VSUBS 0.009392f
C576 B.n460 VSUBS 0.009392f
C577 B.n461 VSUBS 0.009392f
C578 B.n462 VSUBS 0.009392f
C579 B.n463 VSUBS 0.009392f
C580 B.n464 VSUBS 0.009392f
C581 B.n465 VSUBS 0.009392f
C582 B.n466 VSUBS 0.009392f
C583 B.n467 VSUBS 0.009392f
C584 B.n468 VSUBS 0.009392f
C585 B.n469 VSUBS 0.009392f
C586 B.n470 VSUBS 0.009392f
C587 B.n471 VSUBS 0.009392f
C588 B.n472 VSUBS 0.009392f
C589 B.n473 VSUBS 0.009392f
C590 B.n474 VSUBS 0.009392f
C591 B.n475 VSUBS 0.009392f
C592 B.n476 VSUBS 0.009392f
C593 B.n477 VSUBS 0.009392f
C594 B.n478 VSUBS 0.009392f
C595 B.n479 VSUBS 0.009392f
C596 B.n480 VSUBS 0.009392f
C597 B.n481 VSUBS 0.009392f
C598 B.n482 VSUBS 0.009392f
C599 B.n483 VSUBS 0.009392f
C600 B.n484 VSUBS 0.009392f
C601 B.n485 VSUBS 0.009392f
C602 B.n486 VSUBS 0.009392f
C603 B.n487 VSUBS 0.009392f
C604 B.n488 VSUBS 0.009392f
C605 B.n489 VSUBS 0.009392f
C606 B.n490 VSUBS 0.009392f
C607 B.n491 VSUBS 0.009392f
C608 B.n492 VSUBS 0.009392f
C609 B.n493 VSUBS 0.009392f
C610 B.n494 VSUBS 0.009392f
C611 B.n495 VSUBS 0.009392f
C612 B.n496 VSUBS 0.009392f
C613 B.n497 VSUBS 0.009392f
C614 B.n498 VSUBS 0.009392f
C615 B.n499 VSUBS 0.009392f
C616 B.n500 VSUBS 0.009392f
C617 B.n501 VSUBS 0.009392f
C618 B.n502 VSUBS 0.009392f
C619 B.n503 VSUBS 0.009392f
C620 B.n504 VSUBS 0.009392f
C621 B.n505 VSUBS 0.009392f
C622 B.n506 VSUBS 0.009392f
C623 B.n507 VSUBS 0.009392f
C624 B.n508 VSUBS 0.009392f
C625 B.n509 VSUBS 0.009392f
C626 B.n510 VSUBS 0.009392f
C627 B.n511 VSUBS 0.021268f
C628 VDD1.t4 VSUBS 0.019456f
C629 VDD1.t2 VSUBS 0.019456f
C630 VDD1.n0 VSUBS 0.075608f
C631 VDD1.t3 VSUBS 0.019456f
C632 VDD1.t5 VSUBS 0.019456f
C633 VDD1.n1 VSUBS 0.075419f
C634 VDD1.t6 VSUBS 0.019456f
C635 VDD1.t1 VSUBS 0.019456f
C636 VDD1.n2 VSUBS 0.075419f
C637 VDD1.n3 VSUBS 1.80439f
C638 VDD1.t0 VSUBS 0.019456f
C639 VDD1.t7 VSUBS 0.019456f
C640 VDD1.n4 VSUBS 0.073887f
C641 VDD1.n5 VSUBS 1.45255f
C642 VTAIL.t4 VSUBS 0.037701f
C643 VTAIL.t1 VSUBS 0.037701f
C644 VTAIL.n0 VSUBS 0.121942f
C645 VTAIL.n1 VSUBS 0.533484f
C646 VTAIL.t5 VSUBS 0.207769f
C647 VTAIL.n2 VSUBS 0.595681f
C648 VTAIL.t14 VSUBS 0.207769f
C649 VTAIL.n3 VSUBS 0.595681f
C650 VTAIL.t12 VSUBS 0.037701f
C651 VTAIL.t8 VSUBS 0.037701f
C652 VTAIL.n4 VSUBS 0.121942f
C653 VTAIL.n5 VSUBS 0.777002f
C654 VTAIL.t13 VSUBS 0.207769f
C655 VTAIL.n6 VSUBS 1.38944f
C656 VTAIL.t2 VSUBS 0.207769f
C657 VTAIL.n7 VSUBS 1.38944f
C658 VTAIL.t3 VSUBS 0.037701f
C659 VTAIL.t0 VSUBS 0.037701f
C660 VTAIL.n8 VSUBS 0.121942f
C661 VTAIL.n9 VSUBS 0.777001f
C662 VTAIL.t6 VSUBS 0.207769f
C663 VTAIL.n10 VSUBS 0.59568f
C664 VTAIL.t10 VSUBS 0.207769f
C665 VTAIL.n11 VSUBS 0.59568f
C666 VTAIL.t15 VSUBS 0.037701f
C667 VTAIL.t11 VSUBS 0.037701f
C668 VTAIL.n12 VSUBS 0.121942f
C669 VTAIL.n13 VSUBS 0.777001f
C670 VTAIL.t9 VSUBS 0.207769f
C671 VTAIL.n14 VSUBS 1.38944f
C672 VTAIL.t7 VSUBS 0.207769f
C673 VTAIL.n15 VSUBS 1.38305f
C674 VP.n0 VSUBS 0.075266f
C675 VP.t6 VSUBS 0.394236f
C676 VP.n1 VSUBS 0.05557f
C677 VP.n2 VSUBS 0.057092f
C678 VP.t1 VSUBS 0.394236f
C679 VP.n3 VSUBS 0.105872f
C680 VP.n4 VSUBS 0.057092f
C681 VP.n5 VSUBS 0.060923f
C682 VP.n6 VSUBS 0.057092f
C683 VP.n7 VSUBS 0.113132f
C684 VP.n8 VSUBS 0.075266f
C685 VP.t0 VSUBS 0.394236f
C686 VP.n9 VSUBS 0.05557f
C687 VP.n10 VSUBS 0.057092f
C688 VP.t7 VSUBS 0.394236f
C689 VP.n11 VSUBS 0.105872f
C690 VP.n12 VSUBS 0.057092f
C691 VP.n13 VSUBS 0.060923f
C692 VP.t3 VSUBS 0.756465f
C693 VP.t5 VSUBS 0.394236f
C694 VP.n14 VSUBS 0.359986f
C695 VP.n15 VSUBS 0.360314f
C696 VP.n16 VSUBS 0.491591f
C697 VP.n17 VSUBS 0.057092f
C698 VP.n18 VSUBS 0.105872f
C699 VP.n19 VSUBS 0.082992f
C700 VP.n20 VSUBS 0.082992f
C701 VP.n21 VSUBS 0.057092f
C702 VP.n22 VSUBS 0.057092f
C703 VP.n23 VSUBS 0.057092f
C704 VP.n24 VSUBS 0.060923f
C705 VP.n25 VSUBS 0.224744f
C706 VP.n26 VSUBS 0.098554f
C707 VP.n27 VSUBS 0.103154f
C708 VP.n28 VSUBS 0.057092f
C709 VP.n29 VSUBS 0.057092f
C710 VP.n30 VSUBS 0.057092f
C711 VP.n31 VSUBS 0.113132f
C712 VP.n32 VSUBS 0.075557f
C713 VP.n33 VSUBS 0.393505f
C714 VP.n34 VSUBS 2.37123f
C715 VP.n35 VSUBS 2.42088f
C716 VP.t4 VSUBS 0.394236f
C717 VP.n36 VSUBS 0.393505f
C718 VP.n37 VSUBS 0.075557f
C719 VP.n38 VSUBS 0.075266f
C720 VP.n39 VSUBS 0.057092f
C721 VP.n40 VSUBS 0.057092f
C722 VP.n41 VSUBS 0.05557f
C723 VP.n42 VSUBS 0.103154f
C724 VP.t2 VSUBS 0.394236f
C725 VP.n43 VSUBS 0.224744f
C726 VP.n44 VSUBS 0.098554f
C727 VP.n45 VSUBS 0.057092f
C728 VP.n46 VSUBS 0.057092f
C729 VP.n47 VSUBS 0.057092f
C730 VP.n48 VSUBS 0.105872f
C731 VP.n49 VSUBS 0.082992f
C732 VP.n50 VSUBS 0.082992f
C733 VP.n51 VSUBS 0.057092f
C734 VP.n52 VSUBS 0.057092f
C735 VP.n53 VSUBS 0.057092f
C736 VP.n54 VSUBS 0.060923f
C737 VP.n55 VSUBS 0.224744f
C738 VP.n56 VSUBS 0.098554f
C739 VP.n57 VSUBS 0.103154f
C740 VP.n58 VSUBS 0.057092f
C741 VP.n59 VSUBS 0.057092f
C742 VP.n60 VSUBS 0.057092f
C743 VP.n61 VSUBS 0.113132f
C744 VP.n62 VSUBS 0.075557f
C745 VP.n63 VSUBS 0.393505f
C746 VP.n64 VSUBS 0.087339f
.ends

