* NGSPICE file created from diff_pair_sample_1037.ext - technology: sky130A

.subckt diff_pair_sample_1037 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=2.61855 ps=16.2 w=15.87 l=2.56
X1 VDD1.t7 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=6.1893 ps=32.52 w=15.87 l=2.56
X2 VTAIL.t0 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=2.61855 ps=16.2 w=15.87 l=2.56
X3 VDD2.t0 VN.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X4 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=0 ps=0 w=15.87 l=2.56
X5 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=0 ps=0 w=15.87 l=2.56
X6 VTAIL.t13 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X7 VTAIL.t3 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=2.61855 ps=16.2 w=15.87 l=2.56
X8 VDD1.t4 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X9 VDD2.t2 VN.t3 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=6.1893 ps=32.52 w=15.87 l=2.56
X10 VDD2.t5 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X11 VTAIL.t10 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=2.61855 ps=16.2 w=15.87 l=2.56
X12 VTAIL.t2 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X13 VDD2.t7 VN.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=6.1893 ps=32.52 w=15.87 l=2.56
X14 VDD1.t2 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=6.1893 ps=32.52 w=15.87 l=2.56
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=0 ps=0 w=15.87 l=2.56
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1893 pd=32.52 as=0 ps=0 w=15.87 l=2.56
X17 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X18 VDD1.t0 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
X19 VTAIL.t8 VN.t7 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.61855 pd=16.2 as=2.61855 ps=16.2 w=15.87 l=2.56
R0 VN.n7 VN.t0 181.124
R1 VN.n36 VN.t6 181.124
R2 VN.n55 VN.n29 161.3
R3 VN.n54 VN.n53 161.3
R4 VN.n52 VN.n30 161.3
R5 VN.n51 VN.n50 161.3
R6 VN.n49 VN.n31 161.3
R7 VN.n48 VN.n47 161.3
R8 VN.n46 VN.n45 161.3
R9 VN.n44 VN.n33 161.3
R10 VN.n43 VN.n42 161.3
R11 VN.n41 VN.n34 161.3
R12 VN.n40 VN.n39 161.3
R13 VN.n38 VN.n35 161.3
R14 VN.n26 VN.n0 161.3
R15 VN.n25 VN.n24 161.3
R16 VN.n23 VN.n1 161.3
R17 VN.n22 VN.n21 161.3
R18 VN.n20 VN.n2 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n16 161.3
R21 VN.n15 VN.n4 161.3
R22 VN.n14 VN.n13 161.3
R23 VN.n12 VN.n5 161.3
R24 VN.n11 VN.n10 161.3
R25 VN.n9 VN.n6 161.3
R26 VN.n8 VN.t4 149.401
R27 VN.n3 VN.t2 149.401
R28 VN.n27 VN.t3 149.401
R29 VN.n37 VN.t7 149.401
R30 VN.n32 VN.t1 149.401
R31 VN.n56 VN.t5 149.401
R32 VN.n28 VN.n27 106.597
R33 VN.n57 VN.n56 106.597
R34 VN.n8 VN.n7 62.8231
R35 VN.n37 VN.n36 62.8231
R36 VN.n14 VN.n5 56.5193
R37 VN.n43 VN.n34 56.5193
R38 VN.n21 VN.n1 54.0911
R39 VN.n50 VN.n30 54.0911
R40 VN VN.n57 53.8391
R41 VN.n21 VN.n20 26.8957
R42 VN.n50 VN.n49 26.8957
R43 VN.n10 VN.n9 24.4675
R44 VN.n10 VN.n5 24.4675
R45 VN.n15 VN.n14 24.4675
R46 VN.n16 VN.n15 24.4675
R47 VN.n20 VN.n19 24.4675
R48 VN.n25 VN.n1 24.4675
R49 VN.n26 VN.n25 24.4675
R50 VN.n39 VN.n34 24.4675
R51 VN.n39 VN.n38 24.4675
R52 VN.n49 VN.n48 24.4675
R53 VN.n45 VN.n44 24.4675
R54 VN.n44 VN.n43 24.4675
R55 VN.n55 VN.n54 24.4675
R56 VN.n54 VN.n30 24.4675
R57 VN.n19 VN.n3 14.9254
R58 VN.n48 VN.n32 14.9254
R59 VN.n9 VN.n8 9.54263
R60 VN.n16 VN.n3 9.54263
R61 VN.n38 VN.n37 9.54263
R62 VN.n45 VN.n32 9.54263
R63 VN.n36 VN.n35 7.21701
R64 VN.n7 VN.n6 7.21701
R65 VN.n27 VN.n26 4.15989
R66 VN.n56 VN.n55 4.15989
R67 VN.n57 VN.n29 0.278367
R68 VN.n28 VN.n0 0.278367
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153454
R92 VDD2.n2 VDD2.n1 64.9075
R93 VDD2.n2 VDD2.n0 64.9075
R94 VDD2 VDD2.n5 64.9047
R95 VDD2.n4 VDD2.n3 63.7174
R96 VDD2.n4 VDD2.n2 48.6075
R97 VDD2 VDD2.n4 1.30438
R98 VDD2.n5 VDD2.t6 1.24814
R99 VDD2.n5 VDD2.t7 1.24814
R100 VDD2.n3 VDD2.t4 1.24814
R101 VDD2.n3 VDD2.t0 1.24814
R102 VDD2.n1 VDD2.t3 1.24814
R103 VDD2.n1 VDD2.t2 1.24814
R104 VDD2.n0 VDD2.t1 1.24814
R105 VDD2.n0 VDD2.t5 1.24814
R106 VTAIL.n11 VTAIL.t0 48.2862
R107 VTAIL.n10 VTAIL.t9 48.2862
R108 VTAIL.n7 VTAIL.t10 48.2862
R109 VTAIL.n15 VTAIL.t12 48.2861
R110 VTAIL.n2 VTAIL.t15 48.2861
R111 VTAIL.n3 VTAIL.t7 48.2861
R112 VTAIL.n6 VTAIL.t3 48.2861
R113 VTAIL.n14 VTAIL.t4 48.2861
R114 VTAIL.n13 VTAIL.n12 47.0386
R115 VTAIL.n9 VTAIL.n8 47.0386
R116 VTAIL.n1 VTAIL.n0 47.0384
R117 VTAIL.n5 VTAIL.n4 47.0384
R118 VTAIL.n15 VTAIL.n14 28.5393
R119 VTAIL.n7 VTAIL.n6 28.5393
R120 VTAIL.n9 VTAIL.n7 2.49188
R121 VTAIL.n10 VTAIL.n9 2.49188
R122 VTAIL.n13 VTAIL.n11 2.49188
R123 VTAIL.n14 VTAIL.n13 2.49188
R124 VTAIL.n6 VTAIL.n5 2.49188
R125 VTAIL.n5 VTAIL.n3 2.49188
R126 VTAIL.n2 VTAIL.n1 2.49188
R127 VTAIL VTAIL.n15 2.43369
R128 VTAIL.n0 VTAIL.t11 1.24814
R129 VTAIL.n0 VTAIL.t13 1.24814
R130 VTAIL.n4 VTAIL.t6 1.24814
R131 VTAIL.n4 VTAIL.t2 1.24814
R132 VTAIL.n12 VTAIL.t5 1.24814
R133 VTAIL.n12 VTAIL.t1 1.24814
R134 VTAIL.n8 VTAIL.t14 1.24814
R135 VTAIL.n8 VTAIL.t8 1.24814
R136 VTAIL.n11 VTAIL.n10 0.470328
R137 VTAIL.n3 VTAIL.n2 0.470328
R138 VTAIL VTAIL.n1 0.0586897
R139 B.n766 B.n765 585
R140 B.n768 B.n156 585
R141 B.n771 B.n770 585
R142 B.n772 B.n155 585
R143 B.n774 B.n773 585
R144 B.n776 B.n154 585
R145 B.n779 B.n778 585
R146 B.n780 B.n153 585
R147 B.n782 B.n781 585
R148 B.n784 B.n152 585
R149 B.n787 B.n786 585
R150 B.n788 B.n151 585
R151 B.n790 B.n789 585
R152 B.n792 B.n150 585
R153 B.n795 B.n794 585
R154 B.n796 B.n149 585
R155 B.n798 B.n797 585
R156 B.n800 B.n148 585
R157 B.n803 B.n802 585
R158 B.n804 B.n147 585
R159 B.n806 B.n805 585
R160 B.n808 B.n146 585
R161 B.n811 B.n810 585
R162 B.n812 B.n145 585
R163 B.n814 B.n813 585
R164 B.n816 B.n144 585
R165 B.n819 B.n818 585
R166 B.n820 B.n143 585
R167 B.n822 B.n821 585
R168 B.n824 B.n142 585
R169 B.n827 B.n826 585
R170 B.n828 B.n141 585
R171 B.n830 B.n829 585
R172 B.n832 B.n140 585
R173 B.n835 B.n834 585
R174 B.n836 B.n139 585
R175 B.n838 B.n837 585
R176 B.n840 B.n138 585
R177 B.n843 B.n842 585
R178 B.n844 B.n137 585
R179 B.n846 B.n845 585
R180 B.n848 B.n136 585
R181 B.n851 B.n850 585
R182 B.n852 B.n135 585
R183 B.n854 B.n853 585
R184 B.n856 B.n134 585
R185 B.n859 B.n858 585
R186 B.n860 B.n133 585
R187 B.n862 B.n861 585
R188 B.n864 B.n132 585
R189 B.n867 B.n866 585
R190 B.n868 B.n128 585
R191 B.n870 B.n869 585
R192 B.n872 B.n127 585
R193 B.n875 B.n874 585
R194 B.n876 B.n126 585
R195 B.n878 B.n877 585
R196 B.n880 B.n125 585
R197 B.n883 B.n882 585
R198 B.n884 B.n124 585
R199 B.n886 B.n885 585
R200 B.n888 B.n123 585
R201 B.n891 B.n890 585
R202 B.n893 B.n120 585
R203 B.n895 B.n894 585
R204 B.n897 B.n119 585
R205 B.n900 B.n899 585
R206 B.n901 B.n118 585
R207 B.n903 B.n902 585
R208 B.n905 B.n117 585
R209 B.n908 B.n907 585
R210 B.n909 B.n116 585
R211 B.n911 B.n910 585
R212 B.n913 B.n115 585
R213 B.n916 B.n915 585
R214 B.n917 B.n114 585
R215 B.n919 B.n918 585
R216 B.n921 B.n113 585
R217 B.n924 B.n923 585
R218 B.n925 B.n112 585
R219 B.n927 B.n926 585
R220 B.n929 B.n111 585
R221 B.n932 B.n931 585
R222 B.n933 B.n110 585
R223 B.n935 B.n934 585
R224 B.n937 B.n109 585
R225 B.n940 B.n939 585
R226 B.n941 B.n108 585
R227 B.n943 B.n942 585
R228 B.n945 B.n107 585
R229 B.n948 B.n947 585
R230 B.n949 B.n106 585
R231 B.n951 B.n950 585
R232 B.n953 B.n105 585
R233 B.n956 B.n955 585
R234 B.n957 B.n104 585
R235 B.n959 B.n958 585
R236 B.n961 B.n103 585
R237 B.n964 B.n963 585
R238 B.n965 B.n102 585
R239 B.n967 B.n966 585
R240 B.n969 B.n101 585
R241 B.n972 B.n971 585
R242 B.n973 B.n100 585
R243 B.n975 B.n974 585
R244 B.n977 B.n99 585
R245 B.n980 B.n979 585
R246 B.n981 B.n98 585
R247 B.n983 B.n982 585
R248 B.n985 B.n97 585
R249 B.n988 B.n987 585
R250 B.n989 B.n96 585
R251 B.n991 B.n990 585
R252 B.n993 B.n95 585
R253 B.n996 B.n995 585
R254 B.n997 B.n94 585
R255 B.n764 B.n92 585
R256 B.n1000 B.n92 585
R257 B.n763 B.n91 585
R258 B.n1001 B.n91 585
R259 B.n762 B.n90 585
R260 B.n1002 B.n90 585
R261 B.n761 B.n760 585
R262 B.n760 B.n86 585
R263 B.n759 B.n85 585
R264 B.n1008 B.n85 585
R265 B.n758 B.n84 585
R266 B.n1009 B.n84 585
R267 B.n757 B.n83 585
R268 B.n1010 B.n83 585
R269 B.n756 B.n755 585
R270 B.n755 B.n82 585
R271 B.n754 B.n78 585
R272 B.n1016 B.n78 585
R273 B.n753 B.n77 585
R274 B.n1017 B.n77 585
R275 B.n752 B.n76 585
R276 B.n1018 B.n76 585
R277 B.n751 B.n750 585
R278 B.n750 B.n72 585
R279 B.n749 B.n71 585
R280 B.n1024 B.n71 585
R281 B.n748 B.n70 585
R282 B.n1025 B.n70 585
R283 B.n747 B.n69 585
R284 B.n1026 B.n69 585
R285 B.n746 B.n745 585
R286 B.n745 B.n65 585
R287 B.n744 B.n64 585
R288 B.n1032 B.n64 585
R289 B.n743 B.n63 585
R290 B.n1033 B.n63 585
R291 B.n742 B.n62 585
R292 B.n1034 B.n62 585
R293 B.n741 B.n740 585
R294 B.n740 B.n61 585
R295 B.n739 B.n57 585
R296 B.n1040 B.n57 585
R297 B.n738 B.n56 585
R298 B.n1041 B.n56 585
R299 B.n737 B.n55 585
R300 B.n1042 B.n55 585
R301 B.n736 B.n735 585
R302 B.n735 B.n51 585
R303 B.n734 B.n50 585
R304 B.n1048 B.n50 585
R305 B.n733 B.n49 585
R306 B.n1049 B.n49 585
R307 B.n732 B.n48 585
R308 B.n1050 B.n48 585
R309 B.n731 B.n730 585
R310 B.n730 B.n47 585
R311 B.n729 B.n43 585
R312 B.n1056 B.n43 585
R313 B.n728 B.n42 585
R314 B.n1057 B.n42 585
R315 B.n727 B.n41 585
R316 B.n1058 B.n41 585
R317 B.n726 B.n725 585
R318 B.n725 B.n37 585
R319 B.n724 B.n36 585
R320 B.n1064 B.n36 585
R321 B.n723 B.n35 585
R322 B.n1065 B.n35 585
R323 B.n722 B.n34 585
R324 B.n1066 B.n34 585
R325 B.n721 B.n720 585
R326 B.n720 B.n30 585
R327 B.n719 B.n29 585
R328 B.n1072 B.n29 585
R329 B.n718 B.n28 585
R330 B.n1073 B.n28 585
R331 B.n717 B.n27 585
R332 B.n1074 B.n27 585
R333 B.n716 B.n715 585
R334 B.n715 B.n23 585
R335 B.n714 B.n22 585
R336 B.n1080 B.n22 585
R337 B.n713 B.n21 585
R338 B.n1081 B.n21 585
R339 B.n712 B.n20 585
R340 B.n1082 B.n20 585
R341 B.n711 B.n710 585
R342 B.n710 B.n16 585
R343 B.n709 B.n15 585
R344 B.n1088 B.n15 585
R345 B.n708 B.n14 585
R346 B.n1089 B.n14 585
R347 B.n707 B.n13 585
R348 B.n1090 B.n13 585
R349 B.n706 B.n705 585
R350 B.n705 B.n12 585
R351 B.n704 B.n703 585
R352 B.n704 B.n8 585
R353 B.n702 B.n7 585
R354 B.n1097 B.n7 585
R355 B.n701 B.n6 585
R356 B.n1098 B.n6 585
R357 B.n700 B.n5 585
R358 B.n1099 B.n5 585
R359 B.n699 B.n698 585
R360 B.n698 B.n4 585
R361 B.n697 B.n157 585
R362 B.n697 B.n696 585
R363 B.n687 B.n158 585
R364 B.n159 B.n158 585
R365 B.n689 B.n688 585
R366 B.n690 B.n689 585
R367 B.n686 B.n164 585
R368 B.n164 B.n163 585
R369 B.n685 B.n684 585
R370 B.n684 B.n683 585
R371 B.n166 B.n165 585
R372 B.n167 B.n166 585
R373 B.n676 B.n675 585
R374 B.n677 B.n676 585
R375 B.n674 B.n172 585
R376 B.n172 B.n171 585
R377 B.n673 B.n672 585
R378 B.n672 B.n671 585
R379 B.n174 B.n173 585
R380 B.n175 B.n174 585
R381 B.n664 B.n663 585
R382 B.n665 B.n664 585
R383 B.n662 B.n180 585
R384 B.n180 B.n179 585
R385 B.n661 B.n660 585
R386 B.n660 B.n659 585
R387 B.n182 B.n181 585
R388 B.n183 B.n182 585
R389 B.n652 B.n651 585
R390 B.n653 B.n652 585
R391 B.n650 B.n188 585
R392 B.n188 B.n187 585
R393 B.n649 B.n648 585
R394 B.n648 B.n647 585
R395 B.n190 B.n189 585
R396 B.n191 B.n190 585
R397 B.n640 B.n639 585
R398 B.n641 B.n640 585
R399 B.n638 B.n196 585
R400 B.n196 B.n195 585
R401 B.n637 B.n636 585
R402 B.n636 B.n635 585
R403 B.n198 B.n197 585
R404 B.n628 B.n198 585
R405 B.n627 B.n626 585
R406 B.n629 B.n627 585
R407 B.n625 B.n203 585
R408 B.n203 B.n202 585
R409 B.n624 B.n623 585
R410 B.n623 B.n622 585
R411 B.n205 B.n204 585
R412 B.n206 B.n205 585
R413 B.n615 B.n614 585
R414 B.n616 B.n615 585
R415 B.n613 B.n211 585
R416 B.n211 B.n210 585
R417 B.n612 B.n611 585
R418 B.n611 B.n610 585
R419 B.n213 B.n212 585
R420 B.n603 B.n213 585
R421 B.n602 B.n601 585
R422 B.n604 B.n602 585
R423 B.n600 B.n218 585
R424 B.n218 B.n217 585
R425 B.n599 B.n598 585
R426 B.n598 B.n597 585
R427 B.n220 B.n219 585
R428 B.n221 B.n220 585
R429 B.n590 B.n589 585
R430 B.n591 B.n590 585
R431 B.n588 B.n226 585
R432 B.n226 B.n225 585
R433 B.n587 B.n586 585
R434 B.n586 B.n585 585
R435 B.n228 B.n227 585
R436 B.n229 B.n228 585
R437 B.n578 B.n577 585
R438 B.n579 B.n578 585
R439 B.n576 B.n234 585
R440 B.n234 B.n233 585
R441 B.n575 B.n574 585
R442 B.n574 B.n573 585
R443 B.n236 B.n235 585
R444 B.n566 B.n236 585
R445 B.n565 B.n564 585
R446 B.n567 B.n565 585
R447 B.n563 B.n241 585
R448 B.n241 B.n240 585
R449 B.n562 B.n561 585
R450 B.n561 B.n560 585
R451 B.n243 B.n242 585
R452 B.n244 B.n243 585
R453 B.n553 B.n552 585
R454 B.n554 B.n553 585
R455 B.n551 B.n249 585
R456 B.n249 B.n248 585
R457 B.n550 B.n549 585
R458 B.n549 B.n548 585
R459 B.n545 B.n253 585
R460 B.n544 B.n543 585
R461 B.n541 B.n254 585
R462 B.n541 B.n252 585
R463 B.n540 B.n539 585
R464 B.n538 B.n537 585
R465 B.n536 B.n256 585
R466 B.n534 B.n533 585
R467 B.n532 B.n257 585
R468 B.n531 B.n530 585
R469 B.n528 B.n258 585
R470 B.n526 B.n525 585
R471 B.n524 B.n259 585
R472 B.n523 B.n522 585
R473 B.n520 B.n260 585
R474 B.n518 B.n517 585
R475 B.n516 B.n261 585
R476 B.n515 B.n514 585
R477 B.n512 B.n262 585
R478 B.n510 B.n509 585
R479 B.n508 B.n263 585
R480 B.n507 B.n506 585
R481 B.n504 B.n264 585
R482 B.n502 B.n501 585
R483 B.n500 B.n265 585
R484 B.n499 B.n498 585
R485 B.n496 B.n266 585
R486 B.n494 B.n493 585
R487 B.n492 B.n267 585
R488 B.n491 B.n490 585
R489 B.n488 B.n268 585
R490 B.n486 B.n485 585
R491 B.n484 B.n269 585
R492 B.n483 B.n482 585
R493 B.n480 B.n270 585
R494 B.n478 B.n477 585
R495 B.n476 B.n271 585
R496 B.n475 B.n474 585
R497 B.n472 B.n272 585
R498 B.n470 B.n469 585
R499 B.n468 B.n273 585
R500 B.n467 B.n466 585
R501 B.n464 B.n274 585
R502 B.n462 B.n461 585
R503 B.n460 B.n275 585
R504 B.n459 B.n458 585
R505 B.n456 B.n276 585
R506 B.n454 B.n453 585
R507 B.n452 B.n277 585
R508 B.n451 B.n450 585
R509 B.n448 B.n278 585
R510 B.n446 B.n445 585
R511 B.n444 B.n279 585
R512 B.n443 B.n442 585
R513 B.n440 B.n439 585
R514 B.n438 B.n437 585
R515 B.n436 B.n284 585
R516 B.n434 B.n433 585
R517 B.n432 B.n285 585
R518 B.n431 B.n430 585
R519 B.n428 B.n286 585
R520 B.n426 B.n425 585
R521 B.n424 B.n287 585
R522 B.n423 B.n422 585
R523 B.n420 B.n419 585
R524 B.n418 B.n417 585
R525 B.n416 B.n292 585
R526 B.n414 B.n413 585
R527 B.n412 B.n293 585
R528 B.n411 B.n410 585
R529 B.n408 B.n294 585
R530 B.n406 B.n405 585
R531 B.n404 B.n295 585
R532 B.n403 B.n402 585
R533 B.n400 B.n296 585
R534 B.n398 B.n397 585
R535 B.n396 B.n297 585
R536 B.n395 B.n394 585
R537 B.n392 B.n298 585
R538 B.n390 B.n389 585
R539 B.n388 B.n299 585
R540 B.n387 B.n386 585
R541 B.n384 B.n300 585
R542 B.n382 B.n381 585
R543 B.n380 B.n301 585
R544 B.n379 B.n378 585
R545 B.n376 B.n302 585
R546 B.n374 B.n373 585
R547 B.n372 B.n303 585
R548 B.n371 B.n370 585
R549 B.n368 B.n304 585
R550 B.n366 B.n365 585
R551 B.n364 B.n305 585
R552 B.n363 B.n362 585
R553 B.n360 B.n306 585
R554 B.n358 B.n357 585
R555 B.n356 B.n307 585
R556 B.n355 B.n354 585
R557 B.n352 B.n308 585
R558 B.n350 B.n349 585
R559 B.n348 B.n309 585
R560 B.n347 B.n346 585
R561 B.n344 B.n310 585
R562 B.n342 B.n341 585
R563 B.n340 B.n311 585
R564 B.n339 B.n338 585
R565 B.n336 B.n312 585
R566 B.n334 B.n333 585
R567 B.n332 B.n313 585
R568 B.n331 B.n330 585
R569 B.n328 B.n314 585
R570 B.n326 B.n325 585
R571 B.n324 B.n315 585
R572 B.n323 B.n322 585
R573 B.n320 B.n316 585
R574 B.n318 B.n317 585
R575 B.n251 B.n250 585
R576 B.n252 B.n251 585
R577 B.n547 B.n546 585
R578 B.n548 B.n547 585
R579 B.n247 B.n246 585
R580 B.n248 B.n247 585
R581 B.n556 B.n555 585
R582 B.n555 B.n554 585
R583 B.n557 B.n245 585
R584 B.n245 B.n244 585
R585 B.n559 B.n558 585
R586 B.n560 B.n559 585
R587 B.n239 B.n238 585
R588 B.n240 B.n239 585
R589 B.n569 B.n568 585
R590 B.n568 B.n567 585
R591 B.n570 B.n237 585
R592 B.n566 B.n237 585
R593 B.n572 B.n571 585
R594 B.n573 B.n572 585
R595 B.n232 B.n231 585
R596 B.n233 B.n232 585
R597 B.n581 B.n580 585
R598 B.n580 B.n579 585
R599 B.n582 B.n230 585
R600 B.n230 B.n229 585
R601 B.n584 B.n583 585
R602 B.n585 B.n584 585
R603 B.n224 B.n223 585
R604 B.n225 B.n224 585
R605 B.n593 B.n592 585
R606 B.n592 B.n591 585
R607 B.n594 B.n222 585
R608 B.n222 B.n221 585
R609 B.n596 B.n595 585
R610 B.n597 B.n596 585
R611 B.n216 B.n215 585
R612 B.n217 B.n216 585
R613 B.n606 B.n605 585
R614 B.n605 B.n604 585
R615 B.n607 B.n214 585
R616 B.n603 B.n214 585
R617 B.n609 B.n608 585
R618 B.n610 B.n609 585
R619 B.n209 B.n208 585
R620 B.n210 B.n209 585
R621 B.n618 B.n617 585
R622 B.n617 B.n616 585
R623 B.n619 B.n207 585
R624 B.n207 B.n206 585
R625 B.n621 B.n620 585
R626 B.n622 B.n621 585
R627 B.n201 B.n200 585
R628 B.n202 B.n201 585
R629 B.n631 B.n630 585
R630 B.n630 B.n629 585
R631 B.n632 B.n199 585
R632 B.n628 B.n199 585
R633 B.n634 B.n633 585
R634 B.n635 B.n634 585
R635 B.n194 B.n193 585
R636 B.n195 B.n194 585
R637 B.n643 B.n642 585
R638 B.n642 B.n641 585
R639 B.n644 B.n192 585
R640 B.n192 B.n191 585
R641 B.n646 B.n645 585
R642 B.n647 B.n646 585
R643 B.n186 B.n185 585
R644 B.n187 B.n186 585
R645 B.n655 B.n654 585
R646 B.n654 B.n653 585
R647 B.n656 B.n184 585
R648 B.n184 B.n183 585
R649 B.n658 B.n657 585
R650 B.n659 B.n658 585
R651 B.n178 B.n177 585
R652 B.n179 B.n178 585
R653 B.n667 B.n666 585
R654 B.n666 B.n665 585
R655 B.n668 B.n176 585
R656 B.n176 B.n175 585
R657 B.n670 B.n669 585
R658 B.n671 B.n670 585
R659 B.n170 B.n169 585
R660 B.n171 B.n170 585
R661 B.n679 B.n678 585
R662 B.n678 B.n677 585
R663 B.n680 B.n168 585
R664 B.n168 B.n167 585
R665 B.n682 B.n681 585
R666 B.n683 B.n682 585
R667 B.n162 B.n161 585
R668 B.n163 B.n162 585
R669 B.n692 B.n691 585
R670 B.n691 B.n690 585
R671 B.n693 B.n160 585
R672 B.n160 B.n159 585
R673 B.n695 B.n694 585
R674 B.n696 B.n695 585
R675 B.n3 B.n0 585
R676 B.n4 B.n3 585
R677 B.n1096 B.n1 585
R678 B.n1097 B.n1096 585
R679 B.n1095 B.n1094 585
R680 B.n1095 B.n8 585
R681 B.n1093 B.n9 585
R682 B.n12 B.n9 585
R683 B.n1092 B.n1091 585
R684 B.n1091 B.n1090 585
R685 B.n11 B.n10 585
R686 B.n1089 B.n11 585
R687 B.n1087 B.n1086 585
R688 B.n1088 B.n1087 585
R689 B.n1085 B.n17 585
R690 B.n17 B.n16 585
R691 B.n1084 B.n1083 585
R692 B.n1083 B.n1082 585
R693 B.n19 B.n18 585
R694 B.n1081 B.n19 585
R695 B.n1079 B.n1078 585
R696 B.n1080 B.n1079 585
R697 B.n1077 B.n24 585
R698 B.n24 B.n23 585
R699 B.n1076 B.n1075 585
R700 B.n1075 B.n1074 585
R701 B.n26 B.n25 585
R702 B.n1073 B.n26 585
R703 B.n1071 B.n1070 585
R704 B.n1072 B.n1071 585
R705 B.n1069 B.n31 585
R706 B.n31 B.n30 585
R707 B.n1068 B.n1067 585
R708 B.n1067 B.n1066 585
R709 B.n33 B.n32 585
R710 B.n1065 B.n33 585
R711 B.n1063 B.n1062 585
R712 B.n1064 B.n1063 585
R713 B.n1061 B.n38 585
R714 B.n38 B.n37 585
R715 B.n1060 B.n1059 585
R716 B.n1059 B.n1058 585
R717 B.n40 B.n39 585
R718 B.n1057 B.n40 585
R719 B.n1055 B.n1054 585
R720 B.n1056 B.n1055 585
R721 B.n1053 B.n44 585
R722 B.n47 B.n44 585
R723 B.n1052 B.n1051 585
R724 B.n1051 B.n1050 585
R725 B.n46 B.n45 585
R726 B.n1049 B.n46 585
R727 B.n1047 B.n1046 585
R728 B.n1048 B.n1047 585
R729 B.n1045 B.n52 585
R730 B.n52 B.n51 585
R731 B.n1044 B.n1043 585
R732 B.n1043 B.n1042 585
R733 B.n54 B.n53 585
R734 B.n1041 B.n54 585
R735 B.n1039 B.n1038 585
R736 B.n1040 B.n1039 585
R737 B.n1037 B.n58 585
R738 B.n61 B.n58 585
R739 B.n1036 B.n1035 585
R740 B.n1035 B.n1034 585
R741 B.n60 B.n59 585
R742 B.n1033 B.n60 585
R743 B.n1031 B.n1030 585
R744 B.n1032 B.n1031 585
R745 B.n1029 B.n66 585
R746 B.n66 B.n65 585
R747 B.n1028 B.n1027 585
R748 B.n1027 B.n1026 585
R749 B.n68 B.n67 585
R750 B.n1025 B.n68 585
R751 B.n1023 B.n1022 585
R752 B.n1024 B.n1023 585
R753 B.n1021 B.n73 585
R754 B.n73 B.n72 585
R755 B.n1020 B.n1019 585
R756 B.n1019 B.n1018 585
R757 B.n75 B.n74 585
R758 B.n1017 B.n75 585
R759 B.n1015 B.n1014 585
R760 B.n1016 B.n1015 585
R761 B.n1013 B.n79 585
R762 B.n82 B.n79 585
R763 B.n1012 B.n1011 585
R764 B.n1011 B.n1010 585
R765 B.n81 B.n80 585
R766 B.n1009 B.n81 585
R767 B.n1007 B.n1006 585
R768 B.n1008 B.n1007 585
R769 B.n1005 B.n87 585
R770 B.n87 B.n86 585
R771 B.n1004 B.n1003 585
R772 B.n1003 B.n1002 585
R773 B.n89 B.n88 585
R774 B.n1001 B.n89 585
R775 B.n999 B.n998 585
R776 B.n1000 B.n999 585
R777 B.n1100 B.n1099 585
R778 B.n1098 B.n2 585
R779 B.n999 B.n94 482.89
R780 B.n766 B.n92 482.89
R781 B.n549 B.n251 482.89
R782 B.n547 B.n253 482.89
R783 B.n121 B.t16 357.387
R784 B.n129 B.t8 357.387
R785 B.n288 B.t12 357.387
R786 B.n280 B.t19 357.387
R787 B.n767 B.n93 256.663
R788 B.n769 B.n93 256.663
R789 B.n775 B.n93 256.663
R790 B.n777 B.n93 256.663
R791 B.n783 B.n93 256.663
R792 B.n785 B.n93 256.663
R793 B.n791 B.n93 256.663
R794 B.n793 B.n93 256.663
R795 B.n799 B.n93 256.663
R796 B.n801 B.n93 256.663
R797 B.n807 B.n93 256.663
R798 B.n809 B.n93 256.663
R799 B.n815 B.n93 256.663
R800 B.n817 B.n93 256.663
R801 B.n823 B.n93 256.663
R802 B.n825 B.n93 256.663
R803 B.n831 B.n93 256.663
R804 B.n833 B.n93 256.663
R805 B.n839 B.n93 256.663
R806 B.n841 B.n93 256.663
R807 B.n847 B.n93 256.663
R808 B.n849 B.n93 256.663
R809 B.n855 B.n93 256.663
R810 B.n857 B.n93 256.663
R811 B.n863 B.n93 256.663
R812 B.n865 B.n93 256.663
R813 B.n871 B.n93 256.663
R814 B.n873 B.n93 256.663
R815 B.n879 B.n93 256.663
R816 B.n881 B.n93 256.663
R817 B.n887 B.n93 256.663
R818 B.n889 B.n93 256.663
R819 B.n896 B.n93 256.663
R820 B.n898 B.n93 256.663
R821 B.n904 B.n93 256.663
R822 B.n906 B.n93 256.663
R823 B.n912 B.n93 256.663
R824 B.n914 B.n93 256.663
R825 B.n920 B.n93 256.663
R826 B.n922 B.n93 256.663
R827 B.n928 B.n93 256.663
R828 B.n930 B.n93 256.663
R829 B.n936 B.n93 256.663
R830 B.n938 B.n93 256.663
R831 B.n944 B.n93 256.663
R832 B.n946 B.n93 256.663
R833 B.n952 B.n93 256.663
R834 B.n954 B.n93 256.663
R835 B.n960 B.n93 256.663
R836 B.n962 B.n93 256.663
R837 B.n968 B.n93 256.663
R838 B.n970 B.n93 256.663
R839 B.n976 B.n93 256.663
R840 B.n978 B.n93 256.663
R841 B.n984 B.n93 256.663
R842 B.n986 B.n93 256.663
R843 B.n992 B.n93 256.663
R844 B.n994 B.n93 256.663
R845 B.n542 B.n252 256.663
R846 B.n255 B.n252 256.663
R847 B.n535 B.n252 256.663
R848 B.n529 B.n252 256.663
R849 B.n527 B.n252 256.663
R850 B.n521 B.n252 256.663
R851 B.n519 B.n252 256.663
R852 B.n513 B.n252 256.663
R853 B.n511 B.n252 256.663
R854 B.n505 B.n252 256.663
R855 B.n503 B.n252 256.663
R856 B.n497 B.n252 256.663
R857 B.n495 B.n252 256.663
R858 B.n489 B.n252 256.663
R859 B.n487 B.n252 256.663
R860 B.n481 B.n252 256.663
R861 B.n479 B.n252 256.663
R862 B.n473 B.n252 256.663
R863 B.n471 B.n252 256.663
R864 B.n465 B.n252 256.663
R865 B.n463 B.n252 256.663
R866 B.n457 B.n252 256.663
R867 B.n455 B.n252 256.663
R868 B.n449 B.n252 256.663
R869 B.n447 B.n252 256.663
R870 B.n441 B.n252 256.663
R871 B.n283 B.n252 256.663
R872 B.n435 B.n252 256.663
R873 B.n429 B.n252 256.663
R874 B.n427 B.n252 256.663
R875 B.n421 B.n252 256.663
R876 B.n291 B.n252 256.663
R877 B.n415 B.n252 256.663
R878 B.n409 B.n252 256.663
R879 B.n407 B.n252 256.663
R880 B.n401 B.n252 256.663
R881 B.n399 B.n252 256.663
R882 B.n393 B.n252 256.663
R883 B.n391 B.n252 256.663
R884 B.n385 B.n252 256.663
R885 B.n383 B.n252 256.663
R886 B.n377 B.n252 256.663
R887 B.n375 B.n252 256.663
R888 B.n369 B.n252 256.663
R889 B.n367 B.n252 256.663
R890 B.n361 B.n252 256.663
R891 B.n359 B.n252 256.663
R892 B.n353 B.n252 256.663
R893 B.n351 B.n252 256.663
R894 B.n345 B.n252 256.663
R895 B.n343 B.n252 256.663
R896 B.n337 B.n252 256.663
R897 B.n335 B.n252 256.663
R898 B.n329 B.n252 256.663
R899 B.n327 B.n252 256.663
R900 B.n321 B.n252 256.663
R901 B.n319 B.n252 256.663
R902 B.n1102 B.n1101 256.663
R903 B.n995 B.n993 163.367
R904 B.n991 B.n96 163.367
R905 B.n987 B.n985 163.367
R906 B.n983 B.n98 163.367
R907 B.n979 B.n977 163.367
R908 B.n975 B.n100 163.367
R909 B.n971 B.n969 163.367
R910 B.n967 B.n102 163.367
R911 B.n963 B.n961 163.367
R912 B.n959 B.n104 163.367
R913 B.n955 B.n953 163.367
R914 B.n951 B.n106 163.367
R915 B.n947 B.n945 163.367
R916 B.n943 B.n108 163.367
R917 B.n939 B.n937 163.367
R918 B.n935 B.n110 163.367
R919 B.n931 B.n929 163.367
R920 B.n927 B.n112 163.367
R921 B.n923 B.n921 163.367
R922 B.n919 B.n114 163.367
R923 B.n915 B.n913 163.367
R924 B.n911 B.n116 163.367
R925 B.n907 B.n905 163.367
R926 B.n903 B.n118 163.367
R927 B.n899 B.n897 163.367
R928 B.n895 B.n120 163.367
R929 B.n890 B.n888 163.367
R930 B.n886 B.n124 163.367
R931 B.n882 B.n880 163.367
R932 B.n878 B.n126 163.367
R933 B.n874 B.n872 163.367
R934 B.n870 B.n128 163.367
R935 B.n866 B.n864 163.367
R936 B.n862 B.n133 163.367
R937 B.n858 B.n856 163.367
R938 B.n854 B.n135 163.367
R939 B.n850 B.n848 163.367
R940 B.n846 B.n137 163.367
R941 B.n842 B.n840 163.367
R942 B.n838 B.n139 163.367
R943 B.n834 B.n832 163.367
R944 B.n830 B.n141 163.367
R945 B.n826 B.n824 163.367
R946 B.n822 B.n143 163.367
R947 B.n818 B.n816 163.367
R948 B.n814 B.n145 163.367
R949 B.n810 B.n808 163.367
R950 B.n806 B.n147 163.367
R951 B.n802 B.n800 163.367
R952 B.n798 B.n149 163.367
R953 B.n794 B.n792 163.367
R954 B.n790 B.n151 163.367
R955 B.n786 B.n784 163.367
R956 B.n782 B.n153 163.367
R957 B.n778 B.n776 163.367
R958 B.n774 B.n155 163.367
R959 B.n770 B.n768 163.367
R960 B.n549 B.n249 163.367
R961 B.n553 B.n249 163.367
R962 B.n553 B.n243 163.367
R963 B.n561 B.n243 163.367
R964 B.n561 B.n241 163.367
R965 B.n565 B.n241 163.367
R966 B.n565 B.n236 163.367
R967 B.n574 B.n236 163.367
R968 B.n574 B.n234 163.367
R969 B.n578 B.n234 163.367
R970 B.n578 B.n228 163.367
R971 B.n586 B.n228 163.367
R972 B.n586 B.n226 163.367
R973 B.n590 B.n226 163.367
R974 B.n590 B.n220 163.367
R975 B.n598 B.n220 163.367
R976 B.n598 B.n218 163.367
R977 B.n602 B.n218 163.367
R978 B.n602 B.n213 163.367
R979 B.n611 B.n213 163.367
R980 B.n611 B.n211 163.367
R981 B.n615 B.n211 163.367
R982 B.n615 B.n205 163.367
R983 B.n623 B.n205 163.367
R984 B.n623 B.n203 163.367
R985 B.n627 B.n203 163.367
R986 B.n627 B.n198 163.367
R987 B.n636 B.n198 163.367
R988 B.n636 B.n196 163.367
R989 B.n640 B.n196 163.367
R990 B.n640 B.n190 163.367
R991 B.n648 B.n190 163.367
R992 B.n648 B.n188 163.367
R993 B.n652 B.n188 163.367
R994 B.n652 B.n182 163.367
R995 B.n660 B.n182 163.367
R996 B.n660 B.n180 163.367
R997 B.n664 B.n180 163.367
R998 B.n664 B.n174 163.367
R999 B.n672 B.n174 163.367
R1000 B.n672 B.n172 163.367
R1001 B.n676 B.n172 163.367
R1002 B.n676 B.n166 163.367
R1003 B.n684 B.n166 163.367
R1004 B.n684 B.n164 163.367
R1005 B.n689 B.n164 163.367
R1006 B.n689 B.n158 163.367
R1007 B.n697 B.n158 163.367
R1008 B.n698 B.n697 163.367
R1009 B.n698 B.n5 163.367
R1010 B.n6 B.n5 163.367
R1011 B.n7 B.n6 163.367
R1012 B.n704 B.n7 163.367
R1013 B.n705 B.n704 163.367
R1014 B.n705 B.n13 163.367
R1015 B.n14 B.n13 163.367
R1016 B.n15 B.n14 163.367
R1017 B.n710 B.n15 163.367
R1018 B.n710 B.n20 163.367
R1019 B.n21 B.n20 163.367
R1020 B.n22 B.n21 163.367
R1021 B.n715 B.n22 163.367
R1022 B.n715 B.n27 163.367
R1023 B.n28 B.n27 163.367
R1024 B.n29 B.n28 163.367
R1025 B.n720 B.n29 163.367
R1026 B.n720 B.n34 163.367
R1027 B.n35 B.n34 163.367
R1028 B.n36 B.n35 163.367
R1029 B.n725 B.n36 163.367
R1030 B.n725 B.n41 163.367
R1031 B.n42 B.n41 163.367
R1032 B.n43 B.n42 163.367
R1033 B.n730 B.n43 163.367
R1034 B.n730 B.n48 163.367
R1035 B.n49 B.n48 163.367
R1036 B.n50 B.n49 163.367
R1037 B.n735 B.n50 163.367
R1038 B.n735 B.n55 163.367
R1039 B.n56 B.n55 163.367
R1040 B.n57 B.n56 163.367
R1041 B.n740 B.n57 163.367
R1042 B.n740 B.n62 163.367
R1043 B.n63 B.n62 163.367
R1044 B.n64 B.n63 163.367
R1045 B.n745 B.n64 163.367
R1046 B.n745 B.n69 163.367
R1047 B.n70 B.n69 163.367
R1048 B.n71 B.n70 163.367
R1049 B.n750 B.n71 163.367
R1050 B.n750 B.n76 163.367
R1051 B.n77 B.n76 163.367
R1052 B.n78 B.n77 163.367
R1053 B.n755 B.n78 163.367
R1054 B.n755 B.n83 163.367
R1055 B.n84 B.n83 163.367
R1056 B.n85 B.n84 163.367
R1057 B.n760 B.n85 163.367
R1058 B.n760 B.n90 163.367
R1059 B.n91 B.n90 163.367
R1060 B.n92 B.n91 163.367
R1061 B.n543 B.n541 163.367
R1062 B.n541 B.n540 163.367
R1063 B.n537 B.n536 163.367
R1064 B.n534 B.n257 163.367
R1065 B.n530 B.n528 163.367
R1066 B.n526 B.n259 163.367
R1067 B.n522 B.n520 163.367
R1068 B.n518 B.n261 163.367
R1069 B.n514 B.n512 163.367
R1070 B.n510 B.n263 163.367
R1071 B.n506 B.n504 163.367
R1072 B.n502 B.n265 163.367
R1073 B.n498 B.n496 163.367
R1074 B.n494 B.n267 163.367
R1075 B.n490 B.n488 163.367
R1076 B.n486 B.n269 163.367
R1077 B.n482 B.n480 163.367
R1078 B.n478 B.n271 163.367
R1079 B.n474 B.n472 163.367
R1080 B.n470 B.n273 163.367
R1081 B.n466 B.n464 163.367
R1082 B.n462 B.n275 163.367
R1083 B.n458 B.n456 163.367
R1084 B.n454 B.n277 163.367
R1085 B.n450 B.n448 163.367
R1086 B.n446 B.n279 163.367
R1087 B.n442 B.n440 163.367
R1088 B.n437 B.n436 163.367
R1089 B.n434 B.n285 163.367
R1090 B.n430 B.n428 163.367
R1091 B.n426 B.n287 163.367
R1092 B.n422 B.n420 163.367
R1093 B.n417 B.n416 163.367
R1094 B.n414 B.n293 163.367
R1095 B.n410 B.n408 163.367
R1096 B.n406 B.n295 163.367
R1097 B.n402 B.n400 163.367
R1098 B.n398 B.n297 163.367
R1099 B.n394 B.n392 163.367
R1100 B.n390 B.n299 163.367
R1101 B.n386 B.n384 163.367
R1102 B.n382 B.n301 163.367
R1103 B.n378 B.n376 163.367
R1104 B.n374 B.n303 163.367
R1105 B.n370 B.n368 163.367
R1106 B.n366 B.n305 163.367
R1107 B.n362 B.n360 163.367
R1108 B.n358 B.n307 163.367
R1109 B.n354 B.n352 163.367
R1110 B.n350 B.n309 163.367
R1111 B.n346 B.n344 163.367
R1112 B.n342 B.n311 163.367
R1113 B.n338 B.n336 163.367
R1114 B.n334 B.n313 163.367
R1115 B.n330 B.n328 163.367
R1116 B.n326 B.n315 163.367
R1117 B.n322 B.n320 163.367
R1118 B.n318 B.n251 163.367
R1119 B.n547 B.n247 163.367
R1120 B.n555 B.n247 163.367
R1121 B.n555 B.n245 163.367
R1122 B.n559 B.n245 163.367
R1123 B.n559 B.n239 163.367
R1124 B.n568 B.n239 163.367
R1125 B.n568 B.n237 163.367
R1126 B.n572 B.n237 163.367
R1127 B.n572 B.n232 163.367
R1128 B.n580 B.n232 163.367
R1129 B.n580 B.n230 163.367
R1130 B.n584 B.n230 163.367
R1131 B.n584 B.n224 163.367
R1132 B.n592 B.n224 163.367
R1133 B.n592 B.n222 163.367
R1134 B.n596 B.n222 163.367
R1135 B.n596 B.n216 163.367
R1136 B.n605 B.n216 163.367
R1137 B.n605 B.n214 163.367
R1138 B.n609 B.n214 163.367
R1139 B.n609 B.n209 163.367
R1140 B.n617 B.n209 163.367
R1141 B.n617 B.n207 163.367
R1142 B.n621 B.n207 163.367
R1143 B.n621 B.n201 163.367
R1144 B.n630 B.n201 163.367
R1145 B.n630 B.n199 163.367
R1146 B.n634 B.n199 163.367
R1147 B.n634 B.n194 163.367
R1148 B.n642 B.n194 163.367
R1149 B.n642 B.n192 163.367
R1150 B.n646 B.n192 163.367
R1151 B.n646 B.n186 163.367
R1152 B.n654 B.n186 163.367
R1153 B.n654 B.n184 163.367
R1154 B.n658 B.n184 163.367
R1155 B.n658 B.n178 163.367
R1156 B.n666 B.n178 163.367
R1157 B.n666 B.n176 163.367
R1158 B.n670 B.n176 163.367
R1159 B.n670 B.n170 163.367
R1160 B.n678 B.n170 163.367
R1161 B.n678 B.n168 163.367
R1162 B.n682 B.n168 163.367
R1163 B.n682 B.n162 163.367
R1164 B.n691 B.n162 163.367
R1165 B.n691 B.n160 163.367
R1166 B.n695 B.n160 163.367
R1167 B.n695 B.n3 163.367
R1168 B.n1100 B.n3 163.367
R1169 B.n1096 B.n2 163.367
R1170 B.n1096 B.n1095 163.367
R1171 B.n1095 B.n9 163.367
R1172 B.n1091 B.n9 163.367
R1173 B.n1091 B.n11 163.367
R1174 B.n1087 B.n11 163.367
R1175 B.n1087 B.n17 163.367
R1176 B.n1083 B.n17 163.367
R1177 B.n1083 B.n19 163.367
R1178 B.n1079 B.n19 163.367
R1179 B.n1079 B.n24 163.367
R1180 B.n1075 B.n24 163.367
R1181 B.n1075 B.n26 163.367
R1182 B.n1071 B.n26 163.367
R1183 B.n1071 B.n31 163.367
R1184 B.n1067 B.n31 163.367
R1185 B.n1067 B.n33 163.367
R1186 B.n1063 B.n33 163.367
R1187 B.n1063 B.n38 163.367
R1188 B.n1059 B.n38 163.367
R1189 B.n1059 B.n40 163.367
R1190 B.n1055 B.n40 163.367
R1191 B.n1055 B.n44 163.367
R1192 B.n1051 B.n44 163.367
R1193 B.n1051 B.n46 163.367
R1194 B.n1047 B.n46 163.367
R1195 B.n1047 B.n52 163.367
R1196 B.n1043 B.n52 163.367
R1197 B.n1043 B.n54 163.367
R1198 B.n1039 B.n54 163.367
R1199 B.n1039 B.n58 163.367
R1200 B.n1035 B.n58 163.367
R1201 B.n1035 B.n60 163.367
R1202 B.n1031 B.n60 163.367
R1203 B.n1031 B.n66 163.367
R1204 B.n1027 B.n66 163.367
R1205 B.n1027 B.n68 163.367
R1206 B.n1023 B.n68 163.367
R1207 B.n1023 B.n73 163.367
R1208 B.n1019 B.n73 163.367
R1209 B.n1019 B.n75 163.367
R1210 B.n1015 B.n75 163.367
R1211 B.n1015 B.n79 163.367
R1212 B.n1011 B.n79 163.367
R1213 B.n1011 B.n81 163.367
R1214 B.n1007 B.n81 163.367
R1215 B.n1007 B.n87 163.367
R1216 B.n1003 B.n87 163.367
R1217 B.n1003 B.n89 163.367
R1218 B.n999 B.n89 163.367
R1219 B.n129 B.t10 127.903
R1220 B.n288 B.t15 127.903
R1221 B.n121 B.t17 127.882
R1222 B.n280 B.t21 127.882
R1223 B.n130 B.t11 71.8536
R1224 B.n289 B.t14 71.8536
R1225 B.n122 B.t18 71.8329
R1226 B.n281 B.t20 71.8329
R1227 B.n994 B.n94 71.676
R1228 B.n993 B.n992 71.676
R1229 B.n986 B.n96 71.676
R1230 B.n985 B.n984 71.676
R1231 B.n978 B.n98 71.676
R1232 B.n977 B.n976 71.676
R1233 B.n970 B.n100 71.676
R1234 B.n969 B.n968 71.676
R1235 B.n962 B.n102 71.676
R1236 B.n961 B.n960 71.676
R1237 B.n954 B.n104 71.676
R1238 B.n953 B.n952 71.676
R1239 B.n946 B.n106 71.676
R1240 B.n945 B.n944 71.676
R1241 B.n938 B.n108 71.676
R1242 B.n937 B.n936 71.676
R1243 B.n930 B.n110 71.676
R1244 B.n929 B.n928 71.676
R1245 B.n922 B.n112 71.676
R1246 B.n921 B.n920 71.676
R1247 B.n914 B.n114 71.676
R1248 B.n913 B.n912 71.676
R1249 B.n906 B.n116 71.676
R1250 B.n905 B.n904 71.676
R1251 B.n898 B.n118 71.676
R1252 B.n897 B.n896 71.676
R1253 B.n889 B.n120 71.676
R1254 B.n888 B.n887 71.676
R1255 B.n881 B.n124 71.676
R1256 B.n880 B.n879 71.676
R1257 B.n873 B.n126 71.676
R1258 B.n872 B.n871 71.676
R1259 B.n865 B.n128 71.676
R1260 B.n864 B.n863 71.676
R1261 B.n857 B.n133 71.676
R1262 B.n856 B.n855 71.676
R1263 B.n849 B.n135 71.676
R1264 B.n848 B.n847 71.676
R1265 B.n841 B.n137 71.676
R1266 B.n840 B.n839 71.676
R1267 B.n833 B.n139 71.676
R1268 B.n832 B.n831 71.676
R1269 B.n825 B.n141 71.676
R1270 B.n824 B.n823 71.676
R1271 B.n817 B.n143 71.676
R1272 B.n816 B.n815 71.676
R1273 B.n809 B.n145 71.676
R1274 B.n808 B.n807 71.676
R1275 B.n801 B.n147 71.676
R1276 B.n800 B.n799 71.676
R1277 B.n793 B.n149 71.676
R1278 B.n792 B.n791 71.676
R1279 B.n785 B.n151 71.676
R1280 B.n784 B.n783 71.676
R1281 B.n777 B.n153 71.676
R1282 B.n776 B.n775 71.676
R1283 B.n769 B.n155 71.676
R1284 B.n768 B.n767 71.676
R1285 B.n767 B.n766 71.676
R1286 B.n770 B.n769 71.676
R1287 B.n775 B.n774 71.676
R1288 B.n778 B.n777 71.676
R1289 B.n783 B.n782 71.676
R1290 B.n786 B.n785 71.676
R1291 B.n791 B.n790 71.676
R1292 B.n794 B.n793 71.676
R1293 B.n799 B.n798 71.676
R1294 B.n802 B.n801 71.676
R1295 B.n807 B.n806 71.676
R1296 B.n810 B.n809 71.676
R1297 B.n815 B.n814 71.676
R1298 B.n818 B.n817 71.676
R1299 B.n823 B.n822 71.676
R1300 B.n826 B.n825 71.676
R1301 B.n831 B.n830 71.676
R1302 B.n834 B.n833 71.676
R1303 B.n839 B.n838 71.676
R1304 B.n842 B.n841 71.676
R1305 B.n847 B.n846 71.676
R1306 B.n850 B.n849 71.676
R1307 B.n855 B.n854 71.676
R1308 B.n858 B.n857 71.676
R1309 B.n863 B.n862 71.676
R1310 B.n866 B.n865 71.676
R1311 B.n871 B.n870 71.676
R1312 B.n874 B.n873 71.676
R1313 B.n879 B.n878 71.676
R1314 B.n882 B.n881 71.676
R1315 B.n887 B.n886 71.676
R1316 B.n890 B.n889 71.676
R1317 B.n896 B.n895 71.676
R1318 B.n899 B.n898 71.676
R1319 B.n904 B.n903 71.676
R1320 B.n907 B.n906 71.676
R1321 B.n912 B.n911 71.676
R1322 B.n915 B.n914 71.676
R1323 B.n920 B.n919 71.676
R1324 B.n923 B.n922 71.676
R1325 B.n928 B.n927 71.676
R1326 B.n931 B.n930 71.676
R1327 B.n936 B.n935 71.676
R1328 B.n939 B.n938 71.676
R1329 B.n944 B.n943 71.676
R1330 B.n947 B.n946 71.676
R1331 B.n952 B.n951 71.676
R1332 B.n955 B.n954 71.676
R1333 B.n960 B.n959 71.676
R1334 B.n963 B.n962 71.676
R1335 B.n968 B.n967 71.676
R1336 B.n971 B.n970 71.676
R1337 B.n976 B.n975 71.676
R1338 B.n979 B.n978 71.676
R1339 B.n984 B.n983 71.676
R1340 B.n987 B.n986 71.676
R1341 B.n992 B.n991 71.676
R1342 B.n995 B.n994 71.676
R1343 B.n542 B.n253 71.676
R1344 B.n540 B.n255 71.676
R1345 B.n536 B.n535 71.676
R1346 B.n529 B.n257 71.676
R1347 B.n528 B.n527 71.676
R1348 B.n521 B.n259 71.676
R1349 B.n520 B.n519 71.676
R1350 B.n513 B.n261 71.676
R1351 B.n512 B.n511 71.676
R1352 B.n505 B.n263 71.676
R1353 B.n504 B.n503 71.676
R1354 B.n497 B.n265 71.676
R1355 B.n496 B.n495 71.676
R1356 B.n489 B.n267 71.676
R1357 B.n488 B.n487 71.676
R1358 B.n481 B.n269 71.676
R1359 B.n480 B.n479 71.676
R1360 B.n473 B.n271 71.676
R1361 B.n472 B.n471 71.676
R1362 B.n465 B.n273 71.676
R1363 B.n464 B.n463 71.676
R1364 B.n457 B.n275 71.676
R1365 B.n456 B.n455 71.676
R1366 B.n449 B.n277 71.676
R1367 B.n448 B.n447 71.676
R1368 B.n441 B.n279 71.676
R1369 B.n440 B.n283 71.676
R1370 B.n436 B.n435 71.676
R1371 B.n429 B.n285 71.676
R1372 B.n428 B.n427 71.676
R1373 B.n421 B.n287 71.676
R1374 B.n420 B.n291 71.676
R1375 B.n416 B.n415 71.676
R1376 B.n409 B.n293 71.676
R1377 B.n408 B.n407 71.676
R1378 B.n401 B.n295 71.676
R1379 B.n400 B.n399 71.676
R1380 B.n393 B.n297 71.676
R1381 B.n392 B.n391 71.676
R1382 B.n385 B.n299 71.676
R1383 B.n384 B.n383 71.676
R1384 B.n377 B.n301 71.676
R1385 B.n376 B.n375 71.676
R1386 B.n369 B.n303 71.676
R1387 B.n368 B.n367 71.676
R1388 B.n361 B.n305 71.676
R1389 B.n360 B.n359 71.676
R1390 B.n353 B.n307 71.676
R1391 B.n352 B.n351 71.676
R1392 B.n345 B.n309 71.676
R1393 B.n344 B.n343 71.676
R1394 B.n337 B.n311 71.676
R1395 B.n336 B.n335 71.676
R1396 B.n329 B.n313 71.676
R1397 B.n328 B.n327 71.676
R1398 B.n321 B.n315 71.676
R1399 B.n320 B.n319 71.676
R1400 B.n543 B.n542 71.676
R1401 B.n537 B.n255 71.676
R1402 B.n535 B.n534 71.676
R1403 B.n530 B.n529 71.676
R1404 B.n527 B.n526 71.676
R1405 B.n522 B.n521 71.676
R1406 B.n519 B.n518 71.676
R1407 B.n514 B.n513 71.676
R1408 B.n511 B.n510 71.676
R1409 B.n506 B.n505 71.676
R1410 B.n503 B.n502 71.676
R1411 B.n498 B.n497 71.676
R1412 B.n495 B.n494 71.676
R1413 B.n490 B.n489 71.676
R1414 B.n487 B.n486 71.676
R1415 B.n482 B.n481 71.676
R1416 B.n479 B.n478 71.676
R1417 B.n474 B.n473 71.676
R1418 B.n471 B.n470 71.676
R1419 B.n466 B.n465 71.676
R1420 B.n463 B.n462 71.676
R1421 B.n458 B.n457 71.676
R1422 B.n455 B.n454 71.676
R1423 B.n450 B.n449 71.676
R1424 B.n447 B.n446 71.676
R1425 B.n442 B.n441 71.676
R1426 B.n437 B.n283 71.676
R1427 B.n435 B.n434 71.676
R1428 B.n430 B.n429 71.676
R1429 B.n427 B.n426 71.676
R1430 B.n422 B.n421 71.676
R1431 B.n417 B.n291 71.676
R1432 B.n415 B.n414 71.676
R1433 B.n410 B.n409 71.676
R1434 B.n407 B.n406 71.676
R1435 B.n402 B.n401 71.676
R1436 B.n399 B.n398 71.676
R1437 B.n394 B.n393 71.676
R1438 B.n391 B.n390 71.676
R1439 B.n386 B.n385 71.676
R1440 B.n383 B.n382 71.676
R1441 B.n378 B.n377 71.676
R1442 B.n375 B.n374 71.676
R1443 B.n370 B.n369 71.676
R1444 B.n367 B.n366 71.676
R1445 B.n362 B.n361 71.676
R1446 B.n359 B.n358 71.676
R1447 B.n354 B.n353 71.676
R1448 B.n351 B.n350 71.676
R1449 B.n346 B.n345 71.676
R1450 B.n343 B.n342 71.676
R1451 B.n338 B.n337 71.676
R1452 B.n335 B.n334 71.676
R1453 B.n330 B.n329 71.676
R1454 B.n327 B.n326 71.676
R1455 B.n322 B.n321 71.676
R1456 B.n319 B.n318 71.676
R1457 B.n1101 B.n1100 71.676
R1458 B.n1101 B.n2 71.676
R1459 B.n548 B.n252 68.149
R1460 B.n1000 B.n93 68.149
R1461 B.n892 B.n122 59.5399
R1462 B.n131 B.n130 59.5399
R1463 B.n290 B.n289 59.5399
R1464 B.n282 B.n281 59.5399
R1465 B.n122 B.n121 56.049
R1466 B.n130 B.n129 56.049
R1467 B.n289 B.n288 56.049
R1468 B.n281 B.n280 56.049
R1469 B.n548 B.n248 35.3753
R1470 B.n554 B.n248 35.3753
R1471 B.n554 B.n244 35.3753
R1472 B.n560 B.n244 35.3753
R1473 B.n560 B.n240 35.3753
R1474 B.n567 B.n240 35.3753
R1475 B.n567 B.n566 35.3753
R1476 B.n573 B.n233 35.3753
R1477 B.n579 B.n233 35.3753
R1478 B.n579 B.n229 35.3753
R1479 B.n585 B.n229 35.3753
R1480 B.n585 B.n225 35.3753
R1481 B.n591 B.n225 35.3753
R1482 B.n591 B.n221 35.3753
R1483 B.n597 B.n221 35.3753
R1484 B.n597 B.n217 35.3753
R1485 B.n604 B.n217 35.3753
R1486 B.n604 B.n603 35.3753
R1487 B.n610 B.n210 35.3753
R1488 B.n616 B.n210 35.3753
R1489 B.n616 B.n206 35.3753
R1490 B.n622 B.n206 35.3753
R1491 B.n622 B.n202 35.3753
R1492 B.n629 B.n202 35.3753
R1493 B.n629 B.n628 35.3753
R1494 B.n635 B.n195 35.3753
R1495 B.n641 B.n195 35.3753
R1496 B.n641 B.n191 35.3753
R1497 B.n647 B.n191 35.3753
R1498 B.n647 B.n187 35.3753
R1499 B.n653 B.n187 35.3753
R1500 B.n653 B.n183 35.3753
R1501 B.n659 B.n183 35.3753
R1502 B.n665 B.n179 35.3753
R1503 B.n665 B.n175 35.3753
R1504 B.n671 B.n175 35.3753
R1505 B.n671 B.n171 35.3753
R1506 B.n677 B.n171 35.3753
R1507 B.n677 B.n167 35.3753
R1508 B.n683 B.n167 35.3753
R1509 B.n690 B.n163 35.3753
R1510 B.n690 B.n159 35.3753
R1511 B.n696 B.n159 35.3753
R1512 B.n696 B.n4 35.3753
R1513 B.n1099 B.n4 35.3753
R1514 B.n1099 B.n1098 35.3753
R1515 B.n1098 B.n1097 35.3753
R1516 B.n1097 B.n8 35.3753
R1517 B.n12 B.n8 35.3753
R1518 B.n1090 B.n12 35.3753
R1519 B.n1090 B.n1089 35.3753
R1520 B.n1088 B.n16 35.3753
R1521 B.n1082 B.n16 35.3753
R1522 B.n1082 B.n1081 35.3753
R1523 B.n1081 B.n1080 35.3753
R1524 B.n1080 B.n23 35.3753
R1525 B.n1074 B.n23 35.3753
R1526 B.n1074 B.n1073 35.3753
R1527 B.n1072 B.n30 35.3753
R1528 B.n1066 B.n30 35.3753
R1529 B.n1066 B.n1065 35.3753
R1530 B.n1065 B.n1064 35.3753
R1531 B.n1064 B.n37 35.3753
R1532 B.n1058 B.n37 35.3753
R1533 B.n1058 B.n1057 35.3753
R1534 B.n1057 B.n1056 35.3753
R1535 B.n1050 B.n47 35.3753
R1536 B.n1050 B.n1049 35.3753
R1537 B.n1049 B.n1048 35.3753
R1538 B.n1048 B.n51 35.3753
R1539 B.n1042 B.n51 35.3753
R1540 B.n1042 B.n1041 35.3753
R1541 B.n1041 B.n1040 35.3753
R1542 B.n1034 B.n61 35.3753
R1543 B.n1034 B.n1033 35.3753
R1544 B.n1033 B.n1032 35.3753
R1545 B.n1032 B.n65 35.3753
R1546 B.n1026 B.n65 35.3753
R1547 B.n1026 B.n1025 35.3753
R1548 B.n1025 B.n1024 35.3753
R1549 B.n1024 B.n72 35.3753
R1550 B.n1018 B.n72 35.3753
R1551 B.n1018 B.n1017 35.3753
R1552 B.n1017 B.n1016 35.3753
R1553 B.n1010 B.n82 35.3753
R1554 B.n1010 B.n1009 35.3753
R1555 B.n1009 B.n1008 35.3753
R1556 B.n1008 B.n86 35.3753
R1557 B.n1002 B.n86 35.3753
R1558 B.n1002 B.n1001 35.3753
R1559 B.n1001 B.n1000 35.3753
R1560 B.n546 B.n545 31.3761
R1561 B.n550 B.n250 31.3761
R1562 B.n765 B.n764 31.3761
R1563 B.n998 B.n997 31.3761
R1564 B.n610 B.t3 30.1731
R1565 B.t2 B.n179 30.1731
R1566 B.n1073 B.t5 30.1731
R1567 B.n1040 B.t4 30.1731
R1568 B.n628 B.t6 22.8901
R1569 B.n683 B.t7 22.8901
R1570 B.t0 B.n1088 22.8901
R1571 B.n47 B.t1 22.8901
R1572 B.n573 B.t13 19.7688
R1573 B.n1016 B.t9 19.7688
R1574 B B.n1102 18.0485
R1575 B.n566 B.t13 15.607
R1576 B.n82 B.t9 15.607
R1577 B.n635 B.t6 12.4857
R1578 B.t7 B.n163 12.4857
R1579 B.n1089 B.t0 12.4857
R1580 B.n1056 B.t1 12.4857
R1581 B.n546 B.n246 10.6151
R1582 B.n556 B.n246 10.6151
R1583 B.n557 B.n556 10.6151
R1584 B.n558 B.n557 10.6151
R1585 B.n558 B.n238 10.6151
R1586 B.n569 B.n238 10.6151
R1587 B.n570 B.n569 10.6151
R1588 B.n571 B.n570 10.6151
R1589 B.n571 B.n231 10.6151
R1590 B.n581 B.n231 10.6151
R1591 B.n582 B.n581 10.6151
R1592 B.n583 B.n582 10.6151
R1593 B.n583 B.n223 10.6151
R1594 B.n593 B.n223 10.6151
R1595 B.n594 B.n593 10.6151
R1596 B.n595 B.n594 10.6151
R1597 B.n595 B.n215 10.6151
R1598 B.n606 B.n215 10.6151
R1599 B.n607 B.n606 10.6151
R1600 B.n608 B.n607 10.6151
R1601 B.n608 B.n208 10.6151
R1602 B.n618 B.n208 10.6151
R1603 B.n619 B.n618 10.6151
R1604 B.n620 B.n619 10.6151
R1605 B.n620 B.n200 10.6151
R1606 B.n631 B.n200 10.6151
R1607 B.n632 B.n631 10.6151
R1608 B.n633 B.n632 10.6151
R1609 B.n633 B.n193 10.6151
R1610 B.n643 B.n193 10.6151
R1611 B.n644 B.n643 10.6151
R1612 B.n645 B.n644 10.6151
R1613 B.n645 B.n185 10.6151
R1614 B.n655 B.n185 10.6151
R1615 B.n656 B.n655 10.6151
R1616 B.n657 B.n656 10.6151
R1617 B.n657 B.n177 10.6151
R1618 B.n667 B.n177 10.6151
R1619 B.n668 B.n667 10.6151
R1620 B.n669 B.n668 10.6151
R1621 B.n669 B.n169 10.6151
R1622 B.n679 B.n169 10.6151
R1623 B.n680 B.n679 10.6151
R1624 B.n681 B.n680 10.6151
R1625 B.n681 B.n161 10.6151
R1626 B.n692 B.n161 10.6151
R1627 B.n693 B.n692 10.6151
R1628 B.n694 B.n693 10.6151
R1629 B.n694 B.n0 10.6151
R1630 B.n545 B.n544 10.6151
R1631 B.n544 B.n254 10.6151
R1632 B.n539 B.n254 10.6151
R1633 B.n539 B.n538 10.6151
R1634 B.n538 B.n256 10.6151
R1635 B.n533 B.n256 10.6151
R1636 B.n533 B.n532 10.6151
R1637 B.n532 B.n531 10.6151
R1638 B.n531 B.n258 10.6151
R1639 B.n525 B.n258 10.6151
R1640 B.n525 B.n524 10.6151
R1641 B.n524 B.n523 10.6151
R1642 B.n523 B.n260 10.6151
R1643 B.n517 B.n260 10.6151
R1644 B.n517 B.n516 10.6151
R1645 B.n516 B.n515 10.6151
R1646 B.n515 B.n262 10.6151
R1647 B.n509 B.n262 10.6151
R1648 B.n509 B.n508 10.6151
R1649 B.n508 B.n507 10.6151
R1650 B.n507 B.n264 10.6151
R1651 B.n501 B.n264 10.6151
R1652 B.n501 B.n500 10.6151
R1653 B.n500 B.n499 10.6151
R1654 B.n499 B.n266 10.6151
R1655 B.n493 B.n266 10.6151
R1656 B.n493 B.n492 10.6151
R1657 B.n492 B.n491 10.6151
R1658 B.n491 B.n268 10.6151
R1659 B.n485 B.n268 10.6151
R1660 B.n485 B.n484 10.6151
R1661 B.n484 B.n483 10.6151
R1662 B.n483 B.n270 10.6151
R1663 B.n477 B.n270 10.6151
R1664 B.n477 B.n476 10.6151
R1665 B.n476 B.n475 10.6151
R1666 B.n475 B.n272 10.6151
R1667 B.n469 B.n272 10.6151
R1668 B.n469 B.n468 10.6151
R1669 B.n468 B.n467 10.6151
R1670 B.n467 B.n274 10.6151
R1671 B.n461 B.n274 10.6151
R1672 B.n461 B.n460 10.6151
R1673 B.n460 B.n459 10.6151
R1674 B.n459 B.n276 10.6151
R1675 B.n453 B.n276 10.6151
R1676 B.n453 B.n452 10.6151
R1677 B.n452 B.n451 10.6151
R1678 B.n451 B.n278 10.6151
R1679 B.n445 B.n278 10.6151
R1680 B.n445 B.n444 10.6151
R1681 B.n444 B.n443 10.6151
R1682 B.n439 B.n438 10.6151
R1683 B.n438 B.n284 10.6151
R1684 B.n433 B.n284 10.6151
R1685 B.n433 B.n432 10.6151
R1686 B.n432 B.n431 10.6151
R1687 B.n431 B.n286 10.6151
R1688 B.n425 B.n286 10.6151
R1689 B.n425 B.n424 10.6151
R1690 B.n424 B.n423 10.6151
R1691 B.n419 B.n418 10.6151
R1692 B.n418 B.n292 10.6151
R1693 B.n413 B.n292 10.6151
R1694 B.n413 B.n412 10.6151
R1695 B.n412 B.n411 10.6151
R1696 B.n411 B.n294 10.6151
R1697 B.n405 B.n294 10.6151
R1698 B.n405 B.n404 10.6151
R1699 B.n404 B.n403 10.6151
R1700 B.n403 B.n296 10.6151
R1701 B.n397 B.n296 10.6151
R1702 B.n397 B.n396 10.6151
R1703 B.n396 B.n395 10.6151
R1704 B.n395 B.n298 10.6151
R1705 B.n389 B.n298 10.6151
R1706 B.n389 B.n388 10.6151
R1707 B.n388 B.n387 10.6151
R1708 B.n387 B.n300 10.6151
R1709 B.n381 B.n300 10.6151
R1710 B.n381 B.n380 10.6151
R1711 B.n380 B.n379 10.6151
R1712 B.n379 B.n302 10.6151
R1713 B.n373 B.n302 10.6151
R1714 B.n373 B.n372 10.6151
R1715 B.n372 B.n371 10.6151
R1716 B.n371 B.n304 10.6151
R1717 B.n365 B.n304 10.6151
R1718 B.n365 B.n364 10.6151
R1719 B.n364 B.n363 10.6151
R1720 B.n363 B.n306 10.6151
R1721 B.n357 B.n306 10.6151
R1722 B.n357 B.n356 10.6151
R1723 B.n356 B.n355 10.6151
R1724 B.n355 B.n308 10.6151
R1725 B.n349 B.n308 10.6151
R1726 B.n349 B.n348 10.6151
R1727 B.n348 B.n347 10.6151
R1728 B.n347 B.n310 10.6151
R1729 B.n341 B.n310 10.6151
R1730 B.n341 B.n340 10.6151
R1731 B.n340 B.n339 10.6151
R1732 B.n339 B.n312 10.6151
R1733 B.n333 B.n312 10.6151
R1734 B.n333 B.n332 10.6151
R1735 B.n332 B.n331 10.6151
R1736 B.n331 B.n314 10.6151
R1737 B.n325 B.n314 10.6151
R1738 B.n325 B.n324 10.6151
R1739 B.n324 B.n323 10.6151
R1740 B.n323 B.n316 10.6151
R1741 B.n317 B.n316 10.6151
R1742 B.n317 B.n250 10.6151
R1743 B.n551 B.n550 10.6151
R1744 B.n552 B.n551 10.6151
R1745 B.n552 B.n242 10.6151
R1746 B.n562 B.n242 10.6151
R1747 B.n563 B.n562 10.6151
R1748 B.n564 B.n563 10.6151
R1749 B.n564 B.n235 10.6151
R1750 B.n575 B.n235 10.6151
R1751 B.n576 B.n575 10.6151
R1752 B.n577 B.n576 10.6151
R1753 B.n577 B.n227 10.6151
R1754 B.n587 B.n227 10.6151
R1755 B.n588 B.n587 10.6151
R1756 B.n589 B.n588 10.6151
R1757 B.n589 B.n219 10.6151
R1758 B.n599 B.n219 10.6151
R1759 B.n600 B.n599 10.6151
R1760 B.n601 B.n600 10.6151
R1761 B.n601 B.n212 10.6151
R1762 B.n612 B.n212 10.6151
R1763 B.n613 B.n612 10.6151
R1764 B.n614 B.n613 10.6151
R1765 B.n614 B.n204 10.6151
R1766 B.n624 B.n204 10.6151
R1767 B.n625 B.n624 10.6151
R1768 B.n626 B.n625 10.6151
R1769 B.n626 B.n197 10.6151
R1770 B.n637 B.n197 10.6151
R1771 B.n638 B.n637 10.6151
R1772 B.n639 B.n638 10.6151
R1773 B.n639 B.n189 10.6151
R1774 B.n649 B.n189 10.6151
R1775 B.n650 B.n649 10.6151
R1776 B.n651 B.n650 10.6151
R1777 B.n651 B.n181 10.6151
R1778 B.n661 B.n181 10.6151
R1779 B.n662 B.n661 10.6151
R1780 B.n663 B.n662 10.6151
R1781 B.n663 B.n173 10.6151
R1782 B.n673 B.n173 10.6151
R1783 B.n674 B.n673 10.6151
R1784 B.n675 B.n674 10.6151
R1785 B.n675 B.n165 10.6151
R1786 B.n685 B.n165 10.6151
R1787 B.n686 B.n685 10.6151
R1788 B.n688 B.n686 10.6151
R1789 B.n688 B.n687 10.6151
R1790 B.n687 B.n157 10.6151
R1791 B.n699 B.n157 10.6151
R1792 B.n700 B.n699 10.6151
R1793 B.n701 B.n700 10.6151
R1794 B.n702 B.n701 10.6151
R1795 B.n703 B.n702 10.6151
R1796 B.n706 B.n703 10.6151
R1797 B.n707 B.n706 10.6151
R1798 B.n708 B.n707 10.6151
R1799 B.n709 B.n708 10.6151
R1800 B.n711 B.n709 10.6151
R1801 B.n712 B.n711 10.6151
R1802 B.n713 B.n712 10.6151
R1803 B.n714 B.n713 10.6151
R1804 B.n716 B.n714 10.6151
R1805 B.n717 B.n716 10.6151
R1806 B.n718 B.n717 10.6151
R1807 B.n719 B.n718 10.6151
R1808 B.n721 B.n719 10.6151
R1809 B.n722 B.n721 10.6151
R1810 B.n723 B.n722 10.6151
R1811 B.n724 B.n723 10.6151
R1812 B.n726 B.n724 10.6151
R1813 B.n727 B.n726 10.6151
R1814 B.n728 B.n727 10.6151
R1815 B.n729 B.n728 10.6151
R1816 B.n731 B.n729 10.6151
R1817 B.n732 B.n731 10.6151
R1818 B.n733 B.n732 10.6151
R1819 B.n734 B.n733 10.6151
R1820 B.n736 B.n734 10.6151
R1821 B.n737 B.n736 10.6151
R1822 B.n738 B.n737 10.6151
R1823 B.n739 B.n738 10.6151
R1824 B.n741 B.n739 10.6151
R1825 B.n742 B.n741 10.6151
R1826 B.n743 B.n742 10.6151
R1827 B.n744 B.n743 10.6151
R1828 B.n746 B.n744 10.6151
R1829 B.n747 B.n746 10.6151
R1830 B.n748 B.n747 10.6151
R1831 B.n749 B.n748 10.6151
R1832 B.n751 B.n749 10.6151
R1833 B.n752 B.n751 10.6151
R1834 B.n753 B.n752 10.6151
R1835 B.n754 B.n753 10.6151
R1836 B.n756 B.n754 10.6151
R1837 B.n757 B.n756 10.6151
R1838 B.n758 B.n757 10.6151
R1839 B.n759 B.n758 10.6151
R1840 B.n761 B.n759 10.6151
R1841 B.n762 B.n761 10.6151
R1842 B.n763 B.n762 10.6151
R1843 B.n764 B.n763 10.6151
R1844 B.n1094 B.n1 10.6151
R1845 B.n1094 B.n1093 10.6151
R1846 B.n1093 B.n1092 10.6151
R1847 B.n1092 B.n10 10.6151
R1848 B.n1086 B.n10 10.6151
R1849 B.n1086 B.n1085 10.6151
R1850 B.n1085 B.n1084 10.6151
R1851 B.n1084 B.n18 10.6151
R1852 B.n1078 B.n18 10.6151
R1853 B.n1078 B.n1077 10.6151
R1854 B.n1077 B.n1076 10.6151
R1855 B.n1076 B.n25 10.6151
R1856 B.n1070 B.n25 10.6151
R1857 B.n1070 B.n1069 10.6151
R1858 B.n1069 B.n1068 10.6151
R1859 B.n1068 B.n32 10.6151
R1860 B.n1062 B.n32 10.6151
R1861 B.n1062 B.n1061 10.6151
R1862 B.n1061 B.n1060 10.6151
R1863 B.n1060 B.n39 10.6151
R1864 B.n1054 B.n39 10.6151
R1865 B.n1054 B.n1053 10.6151
R1866 B.n1053 B.n1052 10.6151
R1867 B.n1052 B.n45 10.6151
R1868 B.n1046 B.n45 10.6151
R1869 B.n1046 B.n1045 10.6151
R1870 B.n1045 B.n1044 10.6151
R1871 B.n1044 B.n53 10.6151
R1872 B.n1038 B.n53 10.6151
R1873 B.n1038 B.n1037 10.6151
R1874 B.n1037 B.n1036 10.6151
R1875 B.n1036 B.n59 10.6151
R1876 B.n1030 B.n59 10.6151
R1877 B.n1030 B.n1029 10.6151
R1878 B.n1029 B.n1028 10.6151
R1879 B.n1028 B.n67 10.6151
R1880 B.n1022 B.n67 10.6151
R1881 B.n1022 B.n1021 10.6151
R1882 B.n1021 B.n1020 10.6151
R1883 B.n1020 B.n74 10.6151
R1884 B.n1014 B.n74 10.6151
R1885 B.n1014 B.n1013 10.6151
R1886 B.n1013 B.n1012 10.6151
R1887 B.n1012 B.n80 10.6151
R1888 B.n1006 B.n80 10.6151
R1889 B.n1006 B.n1005 10.6151
R1890 B.n1005 B.n1004 10.6151
R1891 B.n1004 B.n88 10.6151
R1892 B.n998 B.n88 10.6151
R1893 B.n997 B.n996 10.6151
R1894 B.n996 B.n95 10.6151
R1895 B.n990 B.n95 10.6151
R1896 B.n990 B.n989 10.6151
R1897 B.n989 B.n988 10.6151
R1898 B.n988 B.n97 10.6151
R1899 B.n982 B.n97 10.6151
R1900 B.n982 B.n981 10.6151
R1901 B.n981 B.n980 10.6151
R1902 B.n980 B.n99 10.6151
R1903 B.n974 B.n99 10.6151
R1904 B.n974 B.n973 10.6151
R1905 B.n973 B.n972 10.6151
R1906 B.n972 B.n101 10.6151
R1907 B.n966 B.n101 10.6151
R1908 B.n966 B.n965 10.6151
R1909 B.n965 B.n964 10.6151
R1910 B.n964 B.n103 10.6151
R1911 B.n958 B.n103 10.6151
R1912 B.n958 B.n957 10.6151
R1913 B.n957 B.n956 10.6151
R1914 B.n956 B.n105 10.6151
R1915 B.n950 B.n105 10.6151
R1916 B.n950 B.n949 10.6151
R1917 B.n949 B.n948 10.6151
R1918 B.n948 B.n107 10.6151
R1919 B.n942 B.n107 10.6151
R1920 B.n942 B.n941 10.6151
R1921 B.n941 B.n940 10.6151
R1922 B.n940 B.n109 10.6151
R1923 B.n934 B.n109 10.6151
R1924 B.n934 B.n933 10.6151
R1925 B.n933 B.n932 10.6151
R1926 B.n932 B.n111 10.6151
R1927 B.n926 B.n111 10.6151
R1928 B.n926 B.n925 10.6151
R1929 B.n925 B.n924 10.6151
R1930 B.n924 B.n113 10.6151
R1931 B.n918 B.n113 10.6151
R1932 B.n918 B.n917 10.6151
R1933 B.n917 B.n916 10.6151
R1934 B.n916 B.n115 10.6151
R1935 B.n910 B.n115 10.6151
R1936 B.n910 B.n909 10.6151
R1937 B.n909 B.n908 10.6151
R1938 B.n908 B.n117 10.6151
R1939 B.n902 B.n117 10.6151
R1940 B.n902 B.n901 10.6151
R1941 B.n901 B.n900 10.6151
R1942 B.n900 B.n119 10.6151
R1943 B.n894 B.n119 10.6151
R1944 B.n894 B.n893 10.6151
R1945 B.n891 B.n123 10.6151
R1946 B.n885 B.n123 10.6151
R1947 B.n885 B.n884 10.6151
R1948 B.n884 B.n883 10.6151
R1949 B.n883 B.n125 10.6151
R1950 B.n877 B.n125 10.6151
R1951 B.n877 B.n876 10.6151
R1952 B.n876 B.n875 10.6151
R1953 B.n875 B.n127 10.6151
R1954 B.n869 B.n868 10.6151
R1955 B.n868 B.n867 10.6151
R1956 B.n867 B.n132 10.6151
R1957 B.n861 B.n132 10.6151
R1958 B.n861 B.n860 10.6151
R1959 B.n860 B.n859 10.6151
R1960 B.n859 B.n134 10.6151
R1961 B.n853 B.n134 10.6151
R1962 B.n853 B.n852 10.6151
R1963 B.n852 B.n851 10.6151
R1964 B.n851 B.n136 10.6151
R1965 B.n845 B.n136 10.6151
R1966 B.n845 B.n844 10.6151
R1967 B.n844 B.n843 10.6151
R1968 B.n843 B.n138 10.6151
R1969 B.n837 B.n138 10.6151
R1970 B.n837 B.n836 10.6151
R1971 B.n836 B.n835 10.6151
R1972 B.n835 B.n140 10.6151
R1973 B.n829 B.n140 10.6151
R1974 B.n829 B.n828 10.6151
R1975 B.n828 B.n827 10.6151
R1976 B.n827 B.n142 10.6151
R1977 B.n821 B.n142 10.6151
R1978 B.n821 B.n820 10.6151
R1979 B.n820 B.n819 10.6151
R1980 B.n819 B.n144 10.6151
R1981 B.n813 B.n144 10.6151
R1982 B.n813 B.n812 10.6151
R1983 B.n812 B.n811 10.6151
R1984 B.n811 B.n146 10.6151
R1985 B.n805 B.n146 10.6151
R1986 B.n805 B.n804 10.6151
R1987 B.n804 B.n803 10.6151
R1988 B.n803 B.n148 10.6151
R1989 B.n797 B.n148 10.6151
R1990 B.n797 B.n796 10.6151
R1991 B.n796 B.n795 10.6151
R1992 B.n795 B.n150 10.6151
R1993 B.n789 B.n150 10.6151
R1994 B.n789 B.n788 10.6151
R1995 B.n788 B.n787 10.6151
R1996 B.n787 B.n152 10.6151
R1997 B.n781 B.n152 10.6151
R1998 B.n781 B.n780 10.6151
R1999 B.n780 B.n779 10.6151
R2000 B.n779 B.n154 10.6151
R2001 B.n773 B.n154 10.6151
R2002 B.n773 B.n772 10.6151
R2003 B.n772 B.n771 10.6151
R2004 B.n771 B.n156 10.6151
R2005 B.n765 B.n156 10.6151
R2006 B.n443 B.n282 9.36635
R2007 B.n419 B.n290 9.36635
R2008 B.n893 B.n892 9.36635
R2009 B.n869 B.n131 9.36635
R2010 B.n1102 B.n0 8.11757
R2011 B.n1102 B.n1 8.11757
R2012 B.n603 B.t3 5.20268
R2013 B.n659 B.t2 5.20268
R2014 B.t5 B.n1072 5.20268
R2015 B.n61 B.t4 5.20268
R2016 B.n439 B.n282 1.24928
R2017 B.n423 B.n290 1.24928
R2018 B.n892 B.n891 1.24928
R2019 B.n131 B.n127 1.24928
R2020 VP.n17 VP.t1 181.124
R2021 VP.n19 VP.n16 161.3
R2022 VP.n21 VP.n20 161.3
R2023 VP.n22 VP.n15 161.3
R2024 VP.n24 VP.n23 161.3
R2025 VP.n25 VP.n14 161.3
R2026 VP.n27 VP.n26 161.3
R2027 VP.n29 VP.n28 161.3
R2028 VP.n30 VP.n12 161.3
R2029 VP.n32 VP.n31 161.3
R2030 VP.n33 VP.n11 161.3
R2031 VP.n35 VP.n34 161.3
R2032 VP.n36 VP.n10 161.3
R2033 VP.n68 VP.n0 161.3
R2034 VP.n67 VP.n66 161.3
R2035 VP.n65 VP.n1 161.3
R2036 VP.n64 VP.n63 161.3
R2037 VP.n62 VP.n2 161.3
R2038 VP.n61 VP.n60 161.3
R2039 VP.n59 VP.n58 161.3
R2040 VP.n57 VP.n4 161.3
R2041 VP.n56 VP.n55 161.3
R2042 VP.n54 VP.n5 161.3
R2043 VP.n53 VP.n52 161.3
R2044 VP.n51 VP.n6 161.3
R2045 VP.n49 VP.n48 161.3
R2046 VP.n47 VP.n7 161.3
R2047 VP.n46 VP.n45 161.3
R2048 VP.n44 VP.n8 161.3
R2049 VP.n43 VP.n42 161.3
R2050 VP.n41 VP.n9 161.3
R2051 VP.n39 VP.t2 149.401
R2052 VP.n50 VP.t7 149.401
R2053 VP.n3 VP.t4 149.401
R2054 VP.n69 VP.t0 149.401
R2055 VP.n37 VP.t5 149.401
R2056 VP.n13 VP.t6 149.401
R2057 VP.n18 VP.t3 149.401
R2058 VP.n40 VP.n39 106.597
R2059 VP.n70 VP.n69 106.597
R2060 VP.n38 VP.n37 106.597
R2061 VP.n18 VP.n17 62.8231
R2062 VP.n56 VP.n5 56.5193
R2063 VP.n24 VP.n15 56.5193
R2064 VP.n45 VP.n44 54.0911
R2065 VP.n63 VP.n1 54.0911
R2066 VP.n31 VP.n11 54.0911
R2067 VP.n40 VP.n38 53.5602
R2068 VP.n45 VP.n7 26.8957
R2069 VP.n63 VP.n62 26.8957
R2070 VP.n31 VP.n30 26.8957
R2071 VP.n43 VP.n9 24.4675
R2072 VP.n44 VP.n43 24.4675
R2073 VP.n49 VP.n7 24.4675
R2074 VP.n52 VP.n51 24.4675
R2075 VP.n52 VP.n5 24.4675
R2076 VP.n57 VP.n56 24.4675
R2077 VP.n58 VP.n57 24.4675
R2078 VP.n62 VP.n61 24.4675
R2079 VP.n67 VP.n1 24.4675
R2080 VP.n68 VP.n67 24.4675
R2081 VP.n35 VP.n11 24.4675
R2082 VP.n36 VP.n35 24.4675
R2083 VP.n25 VP.n24 24.4675
R2084 VP.n26 VP.n25 24.4675
R2085 VP.n30 VP.n29 24.4675
R2086 VP.n20 VP.n19 24.4675
R2087 VP.n20 VP.n15 24.4675
R2088 VP.n50 VP.n49 14.9254
R2089 VP.n61 VP.n3 14.9254
R2090 VP.n29 VP.n13 14.9254
R2091 VP.n51 VP.n50 9.54263
R2092 VP.n58 VP.n3 9.54263
R2093 VP.n26 VP.n13 9.54263
R2094 VP.n19 VP.n18 9.54263
R2095 VP.n17 VP.n16 7.21701
R2096 VP.n39 VP.n9 4.15989
R2097 VP.n69 VP.n68 4.15989
R2098 VP.n37 VP.n36 4.15989
R2099 VP.n38 VP.n10 0.278367
R2100 VP.n41 VP.n40 0.278367
R2101 VP.n70 VP.n0 0.278367
R2102 VP.n21 VP.n16 0.189894
R2103 VP.n22 VP.n21 0.189894
R2104 VP.n23 VP.n22 0.189894
R2105 VP.n23 VP.n14 0.189894
R2106 VP.n27 VP.n14 0.189894
R2107 VP.n28 VP.n27 0.189894
R2108 VP.n28 VP.n12 0.189894
R2109 VP.n32 VP.n12 0.189894
R2110 VP.n33 VP.n32 0.189894
R2111 VP.n34 VP.n33 0.189894
R2112 VP.n34 VP.n10 0.189894
R2113 VP.n42 VP.n41 0.189894
R2114 VP.n42 VP.n8 0.189894
R2115 VP.n46 VP.n8 0.189894
R2116 VP.n47 VP.n46 0.189894
R2117 VP.n48 VP.n47 0.189894
R2118 VP.n48 VP.n6 0.189894
R2119 VP.n53 VP.n6 0.189894
R2120 VP.n54 VP.n53 0.189894
R2121 VP.n55 VP.n54 0.189894
R2122 VP.n55 VP.n4 0.189894
R2123 VP.n59 VP.n4 0.189894
R2124 VP.n60 VP.n59 0.189894
R2125 VP.n60 VP.n2 0.189894
R2126 VP.n64 VP.n2 0.189894
R2127 VP.n65 VP.n64 0.189894
R2128 VP.n66 VP.n65 0.189894
R2129 VP.n66 VP.n0 0.189894
R2130 VP VP.n70 0.153454
R2131 VDD1 VDD1.n0 65.0213
R2132 VDD1.n3 VDD1.n2 64.9075
R2133 VDD1.n3 VDD1.n1 64.9075
R2134 VDD1.n5 VDD1.n4 63.7172
R2135 VDD1.n5 VDD1.n3 49.1905
R2136 VDD1.n4 VDD1.t1 1.24814
R2137 VDD1.n4 VDD1.t2 1.24814
R2138 VDD1.n0 VDD1.t6 1.24814
R2139 VDD1.n0 VDD1.t4 1.24814
R2140 VDD1.n2 VDD1.t3 1.24814
R2141 VDD1.n2 VDD1.t7 1.24814
R2142 VDD1.n1 VDD1.t5 1.24814
R2143 VDD1.n1 VDD1.t0 1.24814
R2144 VDD1 VDD1.n5 1.188
C0 VDD2 VN 11.3162f
C1 VDD1 VP 11.678599f
C2 VP VDD2 0.515413f
C3 VDD1 VTAIL 9.38381f
C4 VTAIL VDD2 9.43796f
C5 VDD1 VDD2 1.75652f
C6 VP VN 8.33372f
C7 VTAIL VN 11.5258f
C8 VTAIL VP 11.539901f
C9 VDD1 VN 0.151654f
C10 VDD2 B 5.601851f
C11 VDD1 B 6.036154f
C12 VTAIL B 12.777831f
C13 VN B 15.676189f
C14 VP B 14.197847f
C15 VDD1.t6 B 0.308766f
C16 VDD1.t4 B 0.308766f
C17 VDD1.n0 B 2.81141f
C18 VDD1.t5 B 0.308766f
C19 VDD1.t0 B 0.308766f
C20 VDD1.n1 B 2.81038f
C21 VDD1.t3 B 0.308766f
C22 VDD1.t7 B 0.308766f
C23 VDD1.n2 B 2.81038f
C24 VDD1.n3 B 3.49044f
C25 VDD1.t1 B 0.308766f
C26 VDD1.t2 B 0.308766f
C27 VDD1.n4 B 2.80117f
C28 VDD1.n5 B 3.20825f
C29 VP.n0 B 0.028903f
C30 VP.t0 B 2.44364f
C31 VP.n1 B 0.038426f
C32 VP.n2 B 0.021923f
C33 VP.t4 B 2.44364f
C34 VP.n3 B 0.852194f
C35 VP.n4 B 0.021923f
C36 VP.n5 B 0.032004f
C37 VP.n6 B 0.021923f
C38 VP.t7 B 2.44364f
C39 VP.n7 B 0.042497f
C40 VP.n8 B 0.021923f
C41 VP.n9 B 0.024115f
C42 VP.n10 B 0.028903f
C43 VP.t5 B 2.44364f
C44 VP.n11 B 0.038426f
C45 VP.n12 B 0.021923f
C46 VP.t6 B 2.44364f
C47 VP.n13 B 0.852194f
C48 VP.n14 B 0.021923f
C49 VP.n15 B 0.032004f
C50 VP.n16 B 0.210582f
C51 VP.t3 B 2.44364f
C52 VP.t1 B 2.61607f
C53 VP.n17 B 0.899371f
C54 VP.n18 B 0.912825f
C55 VP.n19 B 0.028553f
C56 VP.n20 B 0.040859f
C57 VP.n21 B 0.021923f
C58 VP.n22 B 0.021923f
C59 VP.n23 B 0.021923f
C60 VP.n24 B 0.032004f
C61 VP.n25 B 0.040859f
C62 VP.n26 B 0.028553f
C63 VP.n27 B 0.021923f
C64 VP.n28 B 0.021923f
C65 VP.n29 B 0.032991f
C66 VP.n30 B 0.042497f
C67 VP.n31 B 0.023943f
C68 VP.n32 B 0.021923f
C69 VP.n33 B 0.021923f
C70 VP.n34 B 0.021923f
C71 VP.n35 B 0.040859f
C72 VP.n36 B 0.024115f
C73 VP.n37 B 0.917733f
C74 VP.n38 B 1.34915f
C75 VP.t2 B 2.44364f
C76 VP.n39 B 0.917733f
C77 VP.n40 B 1.36386f
C78 VP.n41 B 0.028903f
C79 VP.n42 B 0.021923f
C80 VP.n43 B 0.040859f
C81 VP.n44 B 0.038426f
C82 VP.n45 B 0.023943f
C83 VP.n46 B 0.021923f
C84 VP.n47 B 0.021923f
C85 VP.n48 B 0.021923f
C86 VP.n49 B 0.032991f
C87 VP.n50 B 0.852194f
C88 VP.n51 B 0.028553f
C89 VP.n52 B 0.040859f
C90 VP.n53 B 0.021923f
C91 VP.n54 B 0.021923f
C92 VP.n55 B 0.021923f
C93 VP.n56 B 0.032004f
C94 VP.n57 B 0.040859f
C95 VP.n58 B 0.028553f
C96 VP.n59 B 0.021923f
C97 VP.n60 B 0.021923f
C98 VP.n61 B 0.032991f
C99 VP.n62 B 0.042497f
C100 VP.n63 B 0.023943f
C101 VP.n64 B 0.021923f
C102 VP.n65 B 0.021923f
C103 VP.n66 B 0.021923f
C104 VP.n67 B 0.040859f
C105 VP.n68 B 0.024115f
C106 VP.n69 B 0.917733f
C107 VP.n70 B 0.038255f
C108 VTAIL.t11 B 0.236408f
C109 VTAIL.t13 B 0.236408f
C110 VTAIL.n0 B 2.09187f
C111 VTAIL.n1 B 0.334805f
C112 VTAIL.t15 B 2.67201f
C113 VTAIL.n2 B 0.424418f
C114 VTAIL.t7 B 2.67201f
C115 VTAIL.n3 B 0.424418f
C116 VTAIL.t6 B 0.236408f
C117 VTAIL.t2 B 0.236408f
C118 VTAIL.n4 B 2.09187f
C119 VTAIL.n5 B 0.482601f
C120 VTAIL.t3 B 2.67201f
C121 VTAIL.n6 B 1.63429f
C122 VTAIL.t10 B 2.67202f
C123 VTAIL.n7 B 1.63427f
C124 VTAIL.t14 B 0.236408f
C125 VTAIL.t8 B 0.236408f
C126 VTAIL.n8 B 2.09187f
C127 VTAIL.n9 B 0.482599f
C128 VTAIL.t9 B 2.67202f
C129 VTAIL.n10 B 0.424401f
C130 VTAIL.t0 B 2.67202f
C131 VTAIL.n11 B 0.424401f
C132 VTAIL.t5 B 0.236408f
C133 VTAIL.t1 B 0.236408f
C134 VTAIL.n12 B 2.09187f
C135 VTAIL.n13 B 0.482599f
C136 VTAIL.t4 B 2.67201f
C137 VTAIL.n14 B 1.63429f
C138 VTAIL.t12 B 2.67201f
C139 VTAIL.n15 B 1.63075f
C140 VDD2.t1 B 0.304223f
C141 VDD2.t5 B 0.304223f
C142 VDD2.n0 B 2.76903f
C143 VDD2.t3 B 0.304223f
C144 VDD2.t2 B 0.304223f
C145 VDD2.n1 B 2.76903f
C146 VDD2.n2 B 3.3887f
C147 VDD2.t4 B 0.304223f
C148 VDD2.t0 B 0.304223f
C149 VDD2.n3 B 2.75997f
C150 VDD2.n4 B 3.13094f
C151 VDD2.t6 B 0.304223f
C152 VDD2.t7 B 0.304223f
C153 VDD2.n5 B 2.76899f
C154 VN.n0 B 0.028508f
C155 VN.t3 B 2.41025f
C156 VN.n1 B 0.037902f
C157 VN.n2 B 0.021623f
C158 VN.t2 B 2.41025f
C159 VN.n3 B 0.84055f
C160 VN.n4 B 0.021623f
C161 VN.n5 B 0.031566f
C162 VN.n6 B 0.207705f
C163 VN.t4 B 2.41025f
C164 VN.t0 B 2.58032f
C165 VN.n7 B 0.887082f
C166 VN.n8 B 0.900353f
C167 VN.n9 B 0.028163f
C168 VN.n10 B 0.040301f
C169 VN.n11 B 0.021623f
C170 VN.n12 B 0.021623f
C171 VN.n13 B 0.021623f
C172 VN.n14 B 0.031566f
C173 VN.n15 B 0.040301f
C174 VN.n16 B 0.028163f
C175 VN.n17 B 0.021623f
C176 VN.n18 B 0.021623f
C177 VN.n19 B 0.03254f
C178 VN.n20 B 0.041916f
C179 VN.n21 B 0.023616f
C180 VN.n22 B 0.021623f
C181 VN.n23 B 0.021623f
C182 VN.n24 B 0.021623f
C183 VN.n25 B 0.040301f
C184 VN.n26 B 0.023785f
C185 VN.n27 B 0.905193f
C186 VN.n28 B 0.037732f
C187 VN.n29 B 0.028508f
C188 VN.t5 B 2.41025f
C189 VN.n30 B 0.037902f
C190 VN.n31 B 0.021623f
C191 VN.t1 B 2.41025f
C192 VN.n32 B 0.84055f
C193 VN.n33 B 0.021623f
C194 VN.n34 B 0.031566f
C195 VN.n35 B 0.207705f
C196 VN.t7 B 2.41025f
C197 VN.t6 B 2.58032f
C198 VN.n36 B 0.887082f
C199 VN.n37 B 0.900353f
C200 VN.n38 B 0.028163f
C201 VN.n39 B 0.040301f
C202 VN.n40 B 0.021623f
C203 VN.n41 B 0.021623f
C204 VN.n42 B 0.021623f
C205 VN.n43 B 0.031566f
C206 VN.n44 B 0.040301f
C207 VN.n45 B 0.028163f
C208 VN.n46 B 0.021623f
C209 VN.n47 B 0.021623f
C210 VN.n48 B 0.03254f
C211 VN.n49 B 0.041916f
C212 VN.n50 B 0.023616f
C213 VN.n51 B 0.021623f
C214 VN.n52 B 0.021623f
C215 VN.n53 B 0.021623f
C216 VN.n54 B 0.040301f
C217 VN.n55 B 0.023785f
C218 VN.n56 B 0.905193f
C219 VN.n57 B 1.34221f
.ends

