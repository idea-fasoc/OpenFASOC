* NGSPICE file created from diff_pair_sample_0922.ext - technology: sky130A

.subckt diff_pair_sample_0922 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X1 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=1.5807 ps=9.91 w=9.58 l=2.61
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=0 ps=0 w=9.58 l=2.61
X3 VTAIL.t13 VP.t1 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=1.5807 ps=9.91 w=9.58 l=2.61
X4 VDD1.t7 VP.t2 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=3.7362 ps=19.94 w=9.58 l=2.61
X5 VDD2.t6 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=0 ps=0 w=9.58 l=2.61
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=0 ps=0 w=9.58 l=2.61
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=0 ps=0 w=9.58 l=2.61
X9 VTAIL.t11 VP.t3 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X10 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=3.7362 ps=19.94 w=9.58 l=2.61
X11 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X12 VTAIL.t0 VN.t4 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X13 VTAIL.t10 VP.t4 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=1.5807 ps=9.91 w=9.58 l=2.61
X14 VDD1.t4 VP.t5 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X15 VDD1.t6 VP.t6 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=3.7362 ps=19.94 w=9.58 l=2.61
X16 VDD1.t2 VP.t7 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X17 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=1.5807 ps=9.91 w=9.58 l=2.61
X18 VDD2.t1 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5807 pd=9.91 as=3.7362 ps=19.94 w=9.58 l=2.61
X19 VTAIL.t15 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7362 pd=19.94 as=1.5807 ps=9.91 w=9.58 l=2.61
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n29 VP.n28 161.3
R7 VP.n30 VP.n12 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n33 VP.n11 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n36 VP.n10 161.3
R12 VP.n68 VP.n0 161.3
R13 VP.n67 VP.n66 161.3
R14 VP.n65 VP.n1 161.3
R15 VP.n64 VP.n63 161.3
R16 VP.n62 VP.n2 161.3
R17 VP.n61 VP.n60 161.3
R18 VP.n59 VP.n58 161.3
R19 VP.n57 VP.n4 161.3
R20 VP.n56 VP.n55 161.3
R21 VP.n54 VP.n5 161.3
R22 VP.n53 VP.n52 161.3
R23 VP.n51 VP.n6 161.3
R24 VP.n49 VP.n48 161.3
R25 VP.n47 VP.n7 161.3
R26 VP.n46 VP.n45 161.3
R27 VP.n44 VP.n8 161.3
R28 VP.n43 VP.n42 161.3
R29 VP.n41 VP.n9 161.3
R30 VP.n17 VP.t4 121.51
R31 VP.n40 VP.n39 103.038
R32 VP.n70 VP.n69 103.038
R33 VP.n38 VP.n37 103.038
R34 VP.n39 VP.t1 88.4595
R35 VP.n50 VP.t5 88.4595
R36 VP.n3 VP.t3 88.4595
R37 VP.n69 VP.t2 88.4595
R38 VP.n37 VP.t6 88.4595
R39 VP.n13 VP.t0 88.4595
R40 VP.n18 VP.t7 88.4595
R41 VP.n18 VP.n17 61.7254
R42 VP.n45 VP.n44 56.5617
R43 VP.n56 VP.n5 56.5617
R44 VP.n63 VP.n1 56.5617
R45 VP.n31 VP.n11 56.5617
R46 VP.n24 VP.n15 56.5617
R47 VP.n40 VP.n38 49.0981
R48 VP.n43 VP.n9 24.5923
R49 VP.n44 VP.n43 24.5923
R50 VP.n45 VP.n7 24.5923
R51 VP.n49 VP.n7 24.5923
R52 VP.n52 VP.n51 24.5923
R53 VP.n52 VP.n5 24.5923
R54 VP.n57 VP.n56 24.5923
R55 VP.n58 VP.n57 24.5923
R56 VP.n62 VP.n61 24.5923
R57 VP.n63 VP.n62 24.5923
R58 VP.n67 VP.n1 24.5923
R59 VP.n68 VP.n67 24.5923
R60 VP.n35 VP.n11 24.5923
R61 VP.n36 VP.n35 24.5923
R62 VP.n25 VP.n24 24.5923
R63 VP.n26 VP.n25 24.5923
R64 VP.n30 VP.n29 24.5923
R65 VP.n31 VP.n30 24.5923
R66 VP.n20 VP.n19 24.5923
R67 VP.n20 VP.n15 24.5923
R68 VP.n50 VP.n49 13.7719
R69 VP.n61 VP.n3 13.7719
R70 VP.n29 VP.n13 13.7719
R71 VP.n51 VP.n50 10.8209
R72 VP.n58 VP.n3 10.8209
R73 VP.n26 VP.n13 10.8209
R74 VP.n19 VP.n18 10.8209
R75 VP.n39 VP.n9 7.86989
R76 VP.n69 VP.n68 7.86989
R77 VP.n37 VP.n36 7.86989
R78 VP.n17 VP.n16 6.96699
R79 VP.n38 VP.n10 0.278335
R80 VP.n41 VP.n40 0.278335
R81 VP.n70 VP.n0 0.278335
R82 VP.n21 VP.n16 0.189894
R83 VP.n22 VP.n21 0.189894
R84 VP.n23 VP.n22 0.189894
R85 VP.n23 VP.n14 0.189894
R86 VP.n27 VP.n14 0.189894
R87 VP.n28 VP.n27 0.189894
R88 VP.n28 VP.n12 0.189894
R89 VP.n32 VP.n12 0.189894
R90 VP.n33 VP.n32 0.189894
R91 VP.n34 VP.n33 0.189894
R92 VP.n34 VP.n10 0.189894
R93 VP.n42 VP.n41 0.189894
R94 VP.n42 VP.n8 0.189894
R95 VP.n46 VP.n8 0.189894
R96 VP.n47 VP.n46 0.189894
R97 VP.n48 VP.n47 0.189894
R98 VP.n48 VP.n6 0.189894
R99 VP.n53 VP.n6 0.189894
R100 VP.n54 VP.n53 0.189894
R101 VP.n55 VP.n54 0.189894
R102 VP.n55 VP.n4 0.189894
R103 VP.n59 VP.n4 0.189894
R104 VP.n60 VP.n59 0.189894
R105 VP.n60 VP.n2 0.189894
R106 VP.n64 VP.n2 0.189894
R107 VP.n65 VP.n64 0.189894
R108 VP.n66 VP.n65 0.189894
R109 VP.n66 VP.n0 0.189894
R110 VP VP.n70 0.153485
R111 VDD1 VDD1.n0 63.7497
R112 VDD1.n3 VDD1.n2 63.6359
R113 VDD1.n3 VDD1.n1 63.6359
R114 VDD1.n5 VDD1.n4 62.4241
R115 VDD1.n5 VDD1.n3 43.9621
R116 VDD1.n4 VDD1.t3 2.06731
R117 VDD1.n4 VDD1.t6 2.06731
R118 VDD1.n0 VDD1.t1 2.06731
R119 VDD1.n0 VDD1.t2 2.06731
R120 VDD1.n2 VDD1.t0 2.06731
R121 VDD1.n2 VDD1.t7 2.06731
R122 VDD1.n1 VDD1.t5 2.06731
R123 VDD1.n1 VDD1.t4 2.06731
R124 VDD1 VDD1.n5 1.20955
R125 VTAIL.n11 VTAIL.t10 47.8122
R126 VTAIL.n10 VTAIL.t2 47.8122
R127 VTAIL.n7 VTAIL.t3 47.8122
R128 VTAIL.n15 VTAIL.t5 47.8121
R129 VTAIL.n2 VTAIL.t15 47.8121
R130 VTAIL.n3 VTAIL.t12 47.8121
R131 VTAIL.n6 VTAIL.t13 47.8121
R132 VTAIL.n14 VTAIL.t8 47.8121
R133 VTAIL.n13 VTAIL.n12 45.7454
R134 VTAIL.n9 VTAIL.n8 45.7454
R135 VTAIL.n1 VTAIL.n0 45.7452
R136 VTAIL.n5 VTAIL.n4 45.7452
R137 VTAIL.n15 VTAIL.n14 23.16
R138 VTAIL.n7 VTAIL.n6 23.16
R139 VTAIL.n9 VTAIL.n7 2.53498
R140 VTAIL.n10 VTAIL.n9 2.53498
R141 VTAIL.n13 VTAIL.n11 2.53498
R142 VTAIL.n14 VTAIL.n13 2.53498
R143 VTAIL.n6 VTAIL.n5 2.53498
R144 VTAIL.n5 VTAIL.n3 2.53498
R145 VTAIL.n2 VTAIL.n1 2.53498
R146 VTAIL VTAIL.n15 2.47679
R147 VTAIL.n0 VTAIL.t1 2.06731
R148 VTAIL.n0 VTAIL.t0 2.06731
R149 VTAIL.n4 VTAIL.t9 2.06731
R150 VTAIL.n4 VTAIL.t11 2.06731
R151 VTAIL.n12 VTAIL.t7 2.06731
R152 VTAIL.n12 VTAIL.t14 2.06731
R153 VTAIL.n8 VTAIL.t6 2.06731
R154 VTAIL.n8 VTAIL.t4 2.06731
R155 VTAIL.n11 VTAIL.n10 0.470328
R156 VTAIL.n3 VTAIL.n2 0.470328
R157 VTAIL VTAIL.n1 0.0586897
R158 B.n817 B.n816 585
R159 B.n818 B.n817 585
R160 B.n293 B.n135 585
R161 B.n292 B.n291 585
R162 B.n290 B.n289 585
R163 B.n288 B.n287 585
R164 B.n286 B.n285 585
R165 B.n284 B.n283 585
R166 B.n282 B.n281 585
R167 B.n280 B.n279 585
R168 B.n278 B.n277 585
R169 B.n276 B.n275 585
R170 B.n274 B.n273 585
R171 B.n272 B.n271 585
R172 B.n270 B.n269 585
R173 B.n268 B.n267 585
R174 B.n266 B.n265 585
R175 B.n264 B.n263 585
R176 B.n262 B.n261 585
R177 B.n260 B.n259 585
R178 B.n258 B.n257 585
R179 B.n256 B.n255 585
R180 B.n254 B.n253 585
R181 B.n252 B.n251 585
R182 B.n250 B.n249 585
R183 B.n248 B.n247 585
R184 B.n246 B.n245 585
R185 B.n244 B.n243 585
R186 B.n242 B.n241 585
R187 B.n240 B.n239 585
R188 B.n238 B.n237 585
R189 B.n236 B.n235 585
R190 B.n234 B.n233 585
R191 B.n232 B.n231 585
R192 B.n230 B.n229 585
R193 B.n228 B.n227 585
R194 B.n226 B.n225 585
R195 B.n224 B.n223 585
R196 B.n222 B.n221 585
R197 B.n220 B.n219 585
R198 B.n218 B.n217 585
R199 B.n216 B.n215 585
R200 B.n214 B.n213 585
R201 B.n212 B.n211 585
R202 B.n210 B.n209 585
R203 B.n207 B.n206 585
R204 B.n205 B.n204 585
R205 B.n203 B.n202 585
R206 B.n201 B.n200 585
R207 B.n199 B.n198 585
R208 B.n197 B.n196 585
R209 B.n195 B.n194 585
R210 B.n193 B.n192 585
R211 B.n191 B.n190 585
R212 B.n189 B.n188 585
R213 B.n187 B.n186 585
R214 B.n185 B.n184 585
R215 B.n183 B.n182 585
R216 B.n181 B.n180 585
R217 B.n179 B.n178 585
R218 B.n177 B.n176 585
R219 B.n175 B.n174 585
R220 B.n173 B.n172 585
R221 B.n171 B.n170 585
R222 B.n169 B.n168 585
R223 B.n167 B.n166 585
R224 B.n165 B.n164 585
R225 B.n163 B.n162 585
R226 B.n161 B.n160 585
R227 B.n159 B.n158 585
R228 B.n157 B.n156 585
R229 B.n155 B.n154 585
R230 B.n153 B.n152 585
R231 B.n151 B.n150 585
R232 B.n149 B.n148 585
R233 B.n147 B.n146 585
R234 B.n145 B.n144 585
R235 B.n143 B.n142 585
R236 B.n96 B.n95 585
R237 B.n821 B.n820 585
R238 B.n815 B.n136 585
R239 B.n136 B.n93 585
R240 B.n814 B.n92 585
R241 B.n825 B.n92 585
R242 B.n813 B.n91 585
R243 B.n826 B.n91 585
R244 B.n812 B.n90 585
R245 B.n827 B.n90 585
R246 B.n811 B.n810 585
R247 B.n810 B.n86 585
R248 B.n809 B.n85 585
R249 B.n833 B.n85 585
R250 B.n808 B.n84 585
R251 B.n834 B.n84 585
R252 B.n807 B.n83 585
R253 B.n835 B.n83 585
R254 B.n806 B.n805 585
R255 B.n805 B.n79 585
R256 B.n804 B.n78 585
R257 B.n841 B.n78 585
R258 B.n803 B.n77 585
R259 B.n842 B.n77 585
R260 B.n802 B.n76 585
R261 B.n843 B.n76 585
R262 B.n801 B.n800 585
R263 B.n800 B.n72 585
R264 B.n799 B.n71 585
R265 B.n849 B.n71 585
R266 B.n798 B.n70 585
R267 B.n850 B.n70 585
R268 B.n797 B.n69 585
R269 B.n851 B.n69 585
R270 B.n796 B.n795 585
R271 B.n795 B.n65 585
R272 B.n794 B.n64 585
R273 B.n857 B.n64 585
R274 B.n793 B.n63 585
R275 B.n858 B.n63 585
R276 B.n792 B.n62 585
R277 B.n859 B.n62 585
R278 B.n791 B.n790 585
R279 B.n790 B.n58 585
R280 B.n789 B.n57 585
R281 B.n865 B.n57 585
R282 B.n788 B.n56 585
R283 B.n866 B.n56 585
R284 B.n787 B.n55 585
R285 B.n867 B.n55 585
R286 B.n786 B.n785 585
R287 B.n785 B.n51 585
R288 B.n784 B.n50 585
R289 B.n873 B.n50 585
R290 B.n783 B.n49 585
R291 B.n874 B.n49 585
R292 B.n782 B.n48 585
R293 B.n875 B.n48 585
R294 B.n781 B.n780 585
R295 B.n780 B.n47 585
R296 B.n779 B.n43 585
R297 B.n881 B.n43 585
R298 B.n778 B.n42 585
R299 B.n882 B.n42 585
R300 B.n777 B.n41 585
R301 B.n883 B.n41 585
R302 B.n776 B.n775 585
R303 B.n775 B.n37 585
R304 B.n774 B.n36 585
R305 B.n889 B.n36 585
R306 B.n773 B.n35 585
R307 B.n890 B.n35 585
R308 B.n772 B.n34 585
R309 B.n891 B.n34 585
R310 B.n771 B.n770 585
R311 B.n770 B.n33 585
R312 B.n769 B.n29 585
R313 B.n897 B.n29 585
R314 B.n768 B.n28 585
R315 B.n898 B.n28 585
R316 B.n767 B.n27 585
R317 B.n899 B.n27 585
R318 B.n766 B.n765 585
R319 B.n765 B.n23 585
R320 B.n764 B.n22 585
R321 B.n905 B.n22 585
R322 B.n763 B.n21 585
R323 B.n906 B.n21 585
R324 B.n762 B.n20 585
R325 B.n907 B.n20 585
R326 B.n761 B.n760 585
R327 B.n760 B.n16 585
R328 B.n759 B.n15 585
R329 B.n913 B.n15 585
R330 B.n758 B.n14 585
R331 B.n914 B.n14 585
R332 B.n757 B.n13 585
R333 B.n915 B.n13 585
R334 B.n756 B.n755 585
R335 B.n755 B.n12 585
R336 B.n754 B.n753 585
R337 B.n754 B.n8 585
R338 B.n752 B.n7 585
R339 B.n922 B.n7 585
R340 B.n751 B.n6 585
R341 B.n923 B.n6 585
R342 B.n750 B.n5 585
R343 B.n924 B.n5 585
R344 B.n749 B.n748 585
R345 B.n748 B.n4 585
R346 B.n747 B.n294 585
R347 B.n747 B.n746 585
R348 B.n737 B.n295 585
R349 B.n296 B.n295 585
R350 B.n739 B.n738 585
R351 B.n740 B.n739 585
R352 B.n736 B.n301 585
R353 B.n301 B.n300 585
R354 B.n735 B.n734 585
R355 B.n734 B.n733 585
R356 B.n303 B.n302 585
R357 B.n304 B.n303 585
R358 B.n726 B.n725 585
R359 B.n727 B.n726 585
R360 B.n724 B.n309 585
R361 B.n309 B.n308 585
R362 B.n723 B.n722 585
R363 B.n722 B.n721 585
R364 B.n311 B.n310 585
R365 B.n312 B.n311 585
R366 B.n714 B.n713 585
R367 B.n715 B.n714 585
R368 B.n712 B.n317 585
R369 B.n317 B.n316 585
R370 B.n711 B.n710 585
R371 B.n710 B.n709 585
R372 B.n319 B.n318 585
R373 B.n702 B.n319 585
R374 B.n701 B.n700 585
R375 B.n703 B.n701 585
R376 B.n699 B.n324 585
R377 B.n324 B.n323 585
R378 B.n698 B.n697 585
R379 B.n697 B.n696 585
R380 B.n326 B.n325 585
R381 B.n327 B.n326 585
R382 B.n689 B.n688 585
R383 B.n690 B.n689 585
R384 B.n687 B.n332 585
R385 B.n332 B.n331 585
R386 B.n686 B.n685 585
R387 B.n685 B.n684 585
R388 B.n334 B.n333 585
R389 B.n677 B.n334 585
R390 B.n676 B.n675 585
R391 B.n678 B.n676 585
R392 B.n674 B.n339 585
R393 B.n339 B.n338 585
R394 B.n673 B.n672 585
R395 B.n672 B.n671 585
R396 B.n341 B.n340 585
R397 B.n342 B.n341 585
R398 B.n664 B.n663 585
R399 B.n665 B.n664 585
R400 B.n662 B.n347 585
R401 B.n347 B.n346 585
R402 B.n661 B.n660 585
R403 B.n660 B.n659 585
R404 B.n349 B.n348 585
R405 B.n350 B.n349 585
R406 B.n652 B.n651 585
R407 B.n653 B.n652 585
R408 B.n650 B.n355 585
R409 B.n355 B.n354 585
R410 B.n649 B.n648 585
R411 B.n648 B.n647 585
R412 B.n357 B.n356 585
R413 B.n358 B.n357 585
R414 B.n640 B.n639 585
R415 B.n641 B.n640 585
R416 B.n638 B.n363 585
R417 B.n363 B.n362 585
R418 B.n637 B.n636 585
R419 B.n636 B.n635 585
R420 B.n365 B.n364 585
R421 B.n366 B.n365 585
R422 B.n628 B.n627 585
R423 B.n629 B.n628 585
R424 B.n626 B.n371 585
R425 B.n371 B.n370 585
R426 B.n625 B.n624 585
R427 B.n624 B.n623 585
R428 B.n373 B.n372 585
R429 B.n374 B.n373 585
R430 B.n616 B.n615 585
R431 B.n617 B.n616 585
R432 B.n614 B.n379 585
R433 B.n379 B.n378 585
R434 B.n613 B.n612 585
R435 B.n612 B.n611 585
R436 B.n381 B.n380 585
R437 B.n382 B.n381 585
R438 B.n604 B.n603 585
R439 B.n605 B.n604 585
R440 B.n602 B.n387 585
R441 B.n387 B.n386 585
R442 B.n601 B.n600 585
R443 B.n600 B.n599 585
R444 B.n389 B.n388 585
R445 B.n390 B.n389 585
R446 B.n595 B.n594 585
R447 B.n393 B.n392 585
R448 B.n591 B.n590 585
R449 B.n592 B.n591 585
R450 B.n589 B.n432 585
R451 B.n588 B.n587 585
R452 B.n586 B.n585 585
R453 B.n584 B.n583 585
R454 B.n582 B.n581 585
R455 B.n580 B.n579 585
R456 B.n578 B.n577 585
R457 B.n576 B.n575 585
R458 B.n574 B.n573 585
R459 B.n572 B.n571 585
R460 B.n570 B.n569 585
R461 B.n568 B.n567 585
R462 B.n566 B.n565 585
R463 B.n564 B.n563 585
R464 B.n562 B.n561 585
R465 B.n560 B.n559 585
R466 B.n558 B.n557 585
R467 B.n556 B.n555 585
R468 B.n554 B.n553 585
R469 B.n552 B.n551 585
R470 B.n550 B.n549 585
R471 B.n548 B.n547 585
R472 B.n546 B.n545 585
R473 B.n544 B.n543 585
R474 B.n542 B.n541 585
R475 B.n540 B.n539 585
R476 B.n538 B.n537 585
R477 B.n536 B.n535 585
R478 B.n534 B.n533 585
R479 B.n532 B.n531 585
R480 B.n530 B.n529 585
R481 B.n528 B.n527 585
R482 B.n526 B.n525 585
R483 B.n524 B.n523 585
R484 B.n522 B.n521 585
R485 B.n520 B.n519 585
R486 B.n518 B.n517 585
R487 B.n516 B.n515 585
R488 B.n514 B.n513 585
R489 B.n512 B.n511 585
R490 B.n510 B.n509 585
R491 B.n507 B.n506 585
R492 B.n505 B.n504 585
R493 B.n503 B.n502 585
R494 B.n501 B.n500 585
R495 B.n499 B.n498 585
R496 B.n497 B.n496 585
R497 B.n495 B.n494 585
R498 B.n493 B.n492 585
R499 B.n491 B.n490 585
R500 B.n489 B.n488 585
R501 B.n487 B.n486 585
R502 B.n485 B.n484 585
R503 B.n483 B.n482 585
R504 B.n481 B.n480 585
R505 B.n479 B.n478 585
R506 B.n477 B.n476 585
R507 B.n475 B.n474 585
R508 B.n473 B.n472 585
R509 B.n471 B.n470 585
R510 B.n469 B.n468 585
R511 B.n467 B.n466 585
R512 B.n465 B.n464 585
R513 B.n463 B.n462 585
R514 B.n461 B.n460 585
R515 B.n459 B.n458 585
R516 B.n457 B.n456 585
R517 B.n455 B.n454 585
R518 B.n453 B.n452 585
R519 B.n451 B.n450 585
R520 B.n449 B.n448 585
R521 B.n447 B.n446 585
R522 B.n445 B.n444 585
R523 B.n443 B.n442 585
R524 B.n441 B.n440 585
R525 B.n439 B.n438 585
R526 B.n596 B.n391 585
R527 B.n391 B.n390 585
R528 B.n598 B.n597 585
R529 B.n599 B.n598 585
R530 B.n385 B.n384 585
R531 B.n386 B.n385 585
R532 B.n607 B.n606 585
R533 B.n606 B.n605 585
R534 B.n608 B.n383 585
R535 B.n383 B.n382 585
R536 B.n610 B.n609 585
R537 B.n611 B.n610 585
R538 B.n377 B.n376 585
R539 B.n378 B.n377 585
R540 B.n619 B.n618 585
R541 B.n618 B.n617 585
R542 B.n620 B.n375 585
R543 B.n375 B.n374 585
R544 B.n622 B.n621 585
R545 B.n623 B.n622 585
R546 B.n369 B.n368 585
R547 B.n370 B.n369 585
R548 B.n631 B.n630 585
R549 B.n630 B.n629 585
R550 B.n632 B.n367 585
R551 B.n367 B.n366 585
R552 B.n634 B.n633 585
R553 B.n635 B.n634 585
R554 B.n361 B.n360 585
R555 B.n362 B.n361 585
R556 B.n643 B.n642 585
R557 B.n642 B.n641 585
R558 B.n644 B.n359 585
R559 B.n359 B.n358 585
R560 B.n646 B.n645 585
R561 B.n647 B.n646 585
R562 B.n353 B.n352 585
R563 B.n354 B.n353 585
R564 B.n655 B.n654 585
R565 B.n654 B.n653 585
R566 B.n656 B.n351 585
R567 B.n351 B.n350 585
R568 B.n658 B.n657 585
R569 B.n659 B.n658 585
R570 B.n345 B.n344 585
R571 B.n346 B.n345 585
R572 B.n667 B.n666 585
R573 B.n666 B.n665 585
R574 B.n668 B.n343 585
R575 B.n343 B.n342 585
R576 B.n670 B.n669 585
R577 B.n671 B.n670 585
R578 B.n337 B.n336 585
R579 B.n338 B.n337 585
R580 B.n680 B.n679 585
R581 B.n679 B.n678 585
R582 B.n681 B.n335 585
R583 B.n677 B.n335 585
R584 B.n683 B.n682 585
R585 B.n684 B.n683 585
R586 B.n330 B.n329 585
R587 B.n331 B.n330 585
R588 B.n692 B.n691 585
R589 B.n691 B.n690 585
R590 B.n693 B.n328 585
R591 B.n328 B.n327 585
R592 B.n695 B.n694 585
R593 B.n696 B.n695 585
R594 B.n322 B.n321 585
R595 B.n323 B.n322 585
R596 B.n705 B.n704 585
R597 B.n704 B.n703 585
R598 B.n706 B.n320 585
R599 B.n702 B.n320 585
R600 B.n708 B.n707 585
R601 B.n709 B.n708 585
R602 B.n315 B.n314 585
R603 B.n316 B.n315 585
R604 B.n717 B.n716 585
R605 B.n716 B.n715 585
R606 B.n718 B.n313 585
R607 B.n313 B.n312 585
R608 B.n720 B.n719 585
R609 B.n721 B.n720 585
R610 B.n307 B.n306 585
R611 B.n308 B.n307 585
R612 B.n729 B.n728 585
R613 B.n728 B.n727 585
R614 B.n730 B.n305 585
R615 B.n305 B.n304 585
R616 B.n732 B.n731 585
R617 B.n733 B.n732 585
R618 B.n299 B.n298 585
R619 B.n300 B.n299 585
R620 B.n742 B.n741 585
R621 B.n741 B.n740 585
R622 B.n743 B.n297 585
R623 B.n297 B.n296 585
R624 B.n745 B.n744 585
R625 B.n746 B.n745 585
R626 B.n3 B.n0 585
R627 B.n4 B.n3 585
R628 B.n921 B.n1 585
R629 B.n922 B.n921 585
R630 B.n920 B.n919 585
R631 B.n920 B.n8 585
R632 B.n918 B.n9 585
R633 B.n12 B.n9 585
R634 B.n917 B.n916 585
R635 B.n916 B.n915 585
R636 B.n11 B.n10 585
R637 B.n914 B.n11 585
R638 B.n912 B.n911 585
R639 B.n913 B.n912 585
R640 B.n910 B.n17 585
R641 B.n17 B.n16 585
R642 B.n909 B.n908 585
R643 B.n908 B.n907 585
R644 B.n19 B.n18 585
R645 B.n906 B.n19 585
R646 B.n904 B.n903 585
R647 B.n905 B.n904 585
R648 B.n902 B.n24 585
R649 B.n24 B.n23 585
R650 B.n901 B.n900 585
R651 B.n900 B.n899 585
R652 B.n26 B.n25 585
R653 B.n898 B.n26 585
R654 B.n896 B.n895 585
R655 B.n897 B.n896 585
R656 B.n894 B.n30 585
R657 B.n33 B.n30 585
R658 B.n893 B.n892 585
R659 B.n892 B.n891 585
R660 B.n32 B.n31 585
R661 B.n890 B.n32 585
R662 B.n888 B.n887 585
R663 B.n889 B.n888 585
R664 B.n886 B.n38 585
R665 B.n38 B.n37 585
R666 B.n885 B.n884 585
R667 B.n884 B.n883 585
R668 B.n40 B.n39 585
R669 B.n882 B.n40 585
R670 B.n880 B.n879 585
R671 B.n881 B.n880 585
R672 B.n878 B.n44 585
R673 B.n47 B.n44 585
R674 B.n877 B.n876 585
R675 B.n876 B.n875 585
R676 B.n46 B.n45 585
R677 B.n874 B.n46 585
R678 B.n872 B.n871 585
R679 B.n873 B.n872 585
R680 B.n870 B.n52 585
R681 B.n52 B.n51 585
R682 B.n869 B.n868 585
R683 B.n868 B.n867 585
R684 B.n54 B.n53 585
R685 B.n866 B.n54 585
R686 B.n864 B.n863 585
R687 B.n865 B.n864 585
R688 B.n862 B.n59 585
R689 B.n59 B.n58 585
R690 B.n861 B.n860 585
R691 B.n860 B.n859 585
R692 B.n61 B.n60 585
R693 B.n858 B.n61 585
R694 B.n856 B.n855 585
R695 B.n857 B.n856 585
R696 B.n854 B.n66 585
R697 B.n66 B.n65 585
R698 B.n853 B.n852 585
R699 B.n852 B.n851 585
R700 B.n68 B.n67 585
R701 B.n850 B.n68 585
R702 B.n848 B.n847 585
R703 B.n849 B.n848 585
R704 B.n846 B.n73 585
R705 B.n73 B.n72 585
R706 B.n845 B.n844 585
R707 B.n844 B.n843 585
R708 B.n75 B.n74 585
R709 B.n842 B.n75 585
R710 B.n840 B.n839 585
R711 B.n841 B.n840 585
R712 B.n838 B.n80 585
R713 B.n80 B.n79 585
R714 B.n837 B.n836 585
R715 B.n836 B.n835 585
R716 B.n82 B.n81 585
R717 B.n834 B.n82 585
R718 B.n832 B.n831 585
R719 B.n833 B.n832 585
R720 B.n830 B.n87 585
R721 B.n87 B.n86 585
R722 B.n829 B.n828 585
R723 B.n828 B.n827 585
R724 B.n89 B.n88 585
R725 B.n826 B.n89 585
R726 B.n824 B.n823 585
R727 B.n825 B.n824 585
R728 B.n822 B.n94 585
R729 B.n94 B.n93 585
R730 B.n925 B.n924 585
R731 B.n923 B.n2 585
R732 B.n820 B.n94 439.647
R733 B.n817 B.n136 439.647
R734 B.n438 B.n389 439.647
R735 B.n594 B.n391 439.647
R736 B.n140 B.t15 296.522
R737 B.n137 B.t19 296.522
R738 B.n436 B.t12 296.522
R739 B.n433 B.t8 296.522
R740 B.n818 B.n134 256.663
R741 B.n818 B.n133 256.663
R742 B.n818 B.n132 256.663
R743 B.n818 B.n131 256.663
R744 B.n818 B.n130 256.663
R745 B.n818 B.n129 256.663
R746 B.n818 B.n128 256.663
R747 B.n818 B.n127 256.663
R748 B.n818 B.n126 256.663
R749 B.n818 B.n125 256.663
R750 B.n818 B.n124 256.663
R751 B.n818 B.n123 256.663
R752 B.n818 B.n122 256.663
R753 B.n818 B.n121 256.663
R754 B.n818 B.n120 256.663
R755 B.n818 B.n119 256.663
R756 B.n818 B.n118 256.663
R757 B.n818 B.n117 256.663
R758 B.n818 B.n116 256.663
R759 B.n818 B.n115 256.663
R760 B.n818 B.n114 256.663
R761 B.n818 B.n113 256.663
R762 B.n818 B.n112 256.663
R763 B.n818 B.n111 256.663
R764 B.n818 B.n110 256.663
R765 B.n818 B.n109 256.663
R766 B.n818 B.n108 256.663
R767 B.n818 B.n107 256.663
R768 B.n818 B.n106 256.663
R769 B.n818 B.n105 256.663
R770 B.n818 B.n104 256.663
R771 B.n818 B.n103 256.663
R772 B.n818 B.n102 256.663
R773 B.n818 B.n101 256.663
R774 B.n818 B.n100 256.663
R775 B.n818 B.n99 256.663
R776 B.n818 B.n98 256.663
R777 B.n818 B.n97 256.663
R778 B.n819 B.n818 256.663
R779 B.n593 B.n592 256.663
R780 B.n592 B.n394 256.663
R781 B.n592 B.n395 256.663
R782 B.n592 B.n396 256.663
R783 B.n592 B.n397 256.663
R784 B.n592 B.n398 256.663
R785 B.n592 B.n399 256.663
R786 B.n592 B.n400 256.663
R787 B.n592 B.n401 256.663
R788 B.n592 B.n402 256.663
R789 B.n592 B.n403 256.663
R790 B.n592 B.n404 256.663
R791 B.n592 B.n405 256.663
R792 B.n592 B.n406 256.663
R793 B.n592 B.n407 256.663
R794 B.n592 B.n408 256.663
R795 B.n592 B.n409 256.663
R796 B.n592 B.n410 256.663
R797 B.n592 B.n411 256.663
R798 B.n592 B.n412 256.663
R799 B.n592 B.n413 256.663
R800 B.n592 B.n414 256.663
R801 B.n592 B.n415 256.663
R802 B.n592 B.n416 256.663
R803 B.n592 B.n417 256.663
R804 B.n592 B.n418 256.663
R805 B.n592 B.n419 256.663
R806 B.n592 B.n420 256.663
R807 B.n592 B.n421 256.663
R808 B.n592 B.n422 256.663
R809 B.n592 B.n423 256.663
R810 B.n592 B.n424 256.663
R811 B.n592 B.n425 256.663
R812 B.n592 B.n426 256.663
R813 B.n592 B.n427 256.663
R814 B.n592 B.n428 256.663
R815 B.n592 B.n429 256.663
R816 B.n592 B.n430 256.663
R817 B.n592 B.n431 256.663
R818 B.n927 B.n926 256.663
R819 B.n142 B.n96 163.367
R820 B.n146 B.n145 163.367
R821 B.n150 B.n149 163.367
R822 B.n154 B.n153 163.367
R823 B.n158 B.n157 163.367
R824 B.n162 B.n161 163.367
R825 B.n166 B.n165 163.367
R826 B.n170 B.n169 163.367
R827 B.n174 B.n173 163.367
R828 B.n178 B.n177 163.367
R829 B.n182 B.n181 163.367
R830 B.n186 B.n185 163.367
R831 B.n190 B.n189 163.367
R832 B.n194 B.n193 163.367
R833 B.n198 B.n197 163.367
R834 B.n202 B.n201 163.367
R835 B.n206 B.n205 163.367
R836 B.n211 B.n210 163.367
R837 B.n215 B.n214 163.367
R838 B.n219 B.n218 163.367
R839 B.n223 B.n222 163.367
R840 B.n227 B.n226 163.367
R841 B.n231 B.n230 163.367
R842 B.n235 B.n234 163.367
R843 B.n239 B.n238 163.367
R844 B.n243 B.n242 163.367
R845 B.n247 B.n246 163.367
R846 B.n251 B.n250 163.367
R847 B.n255 B.n254 163.367
R848 B.n259 B.n258 163.367
R849 B.n263 B.n262 163.367
R850 B.n267 B.n266 163.367
R851 B.n271 B.n270 163.367
R852 B.n275 B.n274 163.367
R853 B.n279 B.n278 163.367
R854 B.n283 B.n282 163.367
R855 B.n287 B.n286 163.367
R856 B.n291 B.n290 163.367
R857 B.n817 B.n135 163.367
R858 B.n600 B.n389 163.367
R859 B.n600 B.n387 163.367
R860 B.n604 B.n387 163.367
R861 B.n604 B.n381 163.367
R862 B.n612 B.n381 163.367
R863 B.n612 B.n379 163.367
R864 B.n616 B.n379 163.367
R865 B.n616 B.n373 163.367
R866 B.n624 B.n373 163.367
R867 B.n624 B.n371 163.367
R868 B.n628 B.n371 163.367
R869 B.n628 B.n365 163.367
R870 B.n636 B.n365 163.367
R871 B.n636 B.n363 163.367
R872 B.n640 B.n363 163.367
R873 B.n640 B.n357 163.367
R874 B.n648 B.n357 163.367
R875 B.n648 B.n355 163.367
R876 B.n652 B.n355 163.367
R877 B.n652 B.n349 163.367
R878 B.n660 B.n349 163.367
R879 B.n660 B.n347 163.367
R880 B.n664 B.n347 163.367
R881 B.n664 B.n341 163.367
R882 B.n672 B.n341 163.367
R883 B.n672 B.n339 163.367
R884 B.n676 B.n339 163.367
R885 B.n676 B.n334 163.367
R886 B.n685 B.n334 163.367
R887 B.n685 B.n332 163.367
R888 B.n689 B.n332 163.367
R889 B.n689 B.n326 163.367
R890 B.n697 B.n326 163.367
R891 B.n697 B.n324 163.367
R892 B.n701 B.n324 163.367
R893 B.n701 B.n319 163.367
R894 B.n710 B.n319 163.367
R895 B.n710 B.n317 163.367
R896 B.n714 B.n317 163.367
R897 B.n714 B.n311 163.367
R898 B.n722 B.n311 163.367
R899 B.n722 B.n309 163.367
R900 B.n726 B.n309 163.367
R901 B.n726 B.n303 163.367
R902 B.n734 B.n303 163.367
R903 B.n734 B.n301 163.367
R904 B.n739 B.n301 163.367
R905 B.n739 B.n295 163.367
R906 B.n747 B.n295 163.367
R907 B.n748 B.n747 163.367
R908 B.n748 B.n5 163.367
R909 B.n6 B.n5 163.367
R910 B.n7 B.n6 163.367
R911 B.n754 B.n7 163.367
R912 B.n755 B.n754 163.367
R913 B.n755 B.n13 163.367
R914 B.n14 B.n13 163.367
R915 B.n15 B.n14 163.367
R916 B.n760 B.n15 163.367
R917 B.n760 B.n20 163.367
R918 B.n21 B.n20 163.367
R919 B.n22 B.n21 163.367
R920 B.n765 B.n22 163.367
R921 B.n765 B.n27 163.367
R922 B.n28 B.n27 163.367
R923 B.n29 B.n28 163.367
R924 B.n770 B.n29 163.367
R925 B.n770 B.n34 163.367
R926 B.n35 B.n34 163.367
R927 B.n36 B.n35 163.367
R928 B.n775 B.n36 163.367
R929 B.n775 B.n41 163.367
R930 B.n42 B.n41 163.367
R931 B.n43 B.n42 163.367
R932 B.n780 B.n43 163.367
R933 B.n780 B.n48 163.367
R934 B.n49 B.n48 163.367
R935 B.n50 B.n49 163.367
R936 B.n785 B.n50 163.367
R937 B.n785 B.n55 163.367
R938 B.n56 B.n55 163.367
R939 B.n57 B.n56 163.367
R940 B.n790 B.n57 163.367
R941 B.n790 B.n62 163.367
R942 B.n63 B.n62 163.367
R943 B.n64 B.n63 163.367
R944 B.n795 B.n64 163.367
R945 B.n795 B.n69 163.367
R946 B.n70 B.n69 163.367
R947 B.n71 B.n70 163.367
R948 B.n800 B.n71 163.367
R949 B.n800 B.n76 163.367
R950 B.n77 B.n76 163.367
R951 B.n78 B.n77 163.367
R952 B.n805 B.n78 163.367
R953 B.n805 B.n83 163.367
R954 B.n84 B.n83 163.367
R955 B.n85 B.n84 163.367
R956 B.n810 B.n85 163.367
R957 B.n810 B.n90 163.367
R958 B.n91 B.n90 163.367
R959 B.n92 B.n91 163.367
R960 B.n136 B.n92 163.367
R961 B.n591 B.n393 163.367
R962 B.n591 B.n432 163.367
R963 B.n587 B.n586 163.367
R964 B.n583 B.n582 163.367
R965 B.n579 B.n578 163.367
R966 B.n575 B.n574 163.367
R967 B.n571 B.n570 163.367
R968 B.n567 B.n566 163.367
R969 B.n563 B.n562 163.367
R970 B.n559 B.n558 163.367
R971 B.n555 B.n554 163.367
R972 B.n551 B.n550 163.367
R973 B.n547 B.n546 163.367
R974 B.n543 B.n542 163.367
R975 B.n539 B.n538 163.367
R976 B.n535 B.n534 163.367
R977 B.n531 B.n530 163.367
R978 B.n527 B.n526 163.367
R979 B.n523 B.n522 163.367
R980 B.n519 B.n518 163.367
R981 B.n515 B.n514 163.367
R982 B.n511 B.n510 163.367
R983 B.n506 B.n505 163.367
R984 B.n502 B.n501 163.367
R985 B.n498 B.n497 163.367
R986 B.n494 B.n493 163.367
R987 B.n490 B.n489 163.367
R988 B.n486 B.n485 163.367
R989 B.n482 B.n481 163.367
R990 B.n478 B.n477 163.367
R991 B.n474 B.n473 163.367
R992 B.n470 B.n469 163.367
R993 B.n466 B.n465 163.367
R994 B.n462 B.n461 163.367
R995 B.n458 B.n457 163.367
R996 B.n454 B.n453 163.367
R997 B.n450 B.n449 163.367
R998 B.n446 B.n445 163.367
R999 B.n442 B.n441 163.367
R1000 B.n598 B.n391 163.367
R1001 B.n598 B.n385 163.367
R1002 B.n606 B.n385 163.367
R1003 B.n606 B.n383 163.367
R1004 B.n610 B.n383 163.367
R1005 B.n610 B.n377 163.367
R1006 B.n618 B.n377 163.367
R1007 B.n618 B.n375 163.367
R1008 B.n622 B.n375 163.367
R1009 B.n622 B.n369 163.367
R1010 B.n630 B.n369 163.367
R1011 B.n630 B.n367 163.367
R1012 B.n634 B.n367 163.367
R1013 B.n634 B.n361 163.367
R1014 B.n642 B.n361 163.367
R1015 B.n642 B.n359 163.367
R1016 B.n646 B.n359 163.367
R1017 B.n646 B.n353 163.367
R1018 B.n654 B.n353 163.367
R1019 B.n654 B.n351 163.367
R1020 B.n658 B.n351 163.367
R1021 B.n658 B.n345 163.367
R1022 B.n666 B.n345 163.367
R1023 B.n666 B.n343 163.367
R1024 B.n670 B.n343 163.367
R1025 B.n670 B.n337 163.367
R1026 B.n679 B.n337 163.367
R1027 B.n679 B.n335 163.367
R1028 B.n683 B.n335 163.367
R1029 B.n683 B.n330 163.367
R1030 B.n691 B.n330 163.367
R1031 B.n691 B.n328 163.367
R1032 B.n695 B.n328 163.367
R1033 B.n695 B.n322 163.367
R1034 B.n704 B.n322 163.367
R1035 B.n704 B.n320 163.367
R1036 B.n708 B.n320 163.367
R1037 B.n708 B.n315 163.367
R1038 B.n716 B.n315 163.367
R1039 B.n716 B.n313 163.367
R1040 B.n720 B.n313 163.367
R1041 B.n720 B.n307 163.367
R1042 B.n728 B.n307 163.367
R1043 B.n728 B.n305 163.367
R1044 B.n732 B.n305 163.367
R1045 B.n732 B.n299 163.367
R1046 B.n741 B.n299 163.367
R1047 B.n741 B.n297 163.367
R1048 B.n745 B.n297 163.367
R1049 B.n745 B.n3 163.367
R1050 B.n925 B.n3 163.367
R1051 B.n921 B.n2 163.367
R1052 B.n921 B.n920 163.367
R1053 B.n920 B.n9 163.367
R1054 B.n916 B.n9 163.367
R1055 B.n916 B.n11 163.367
R1056 B.n912 B.n11 163.367
R1057 B.n912 B.n17 163.367
R1058 B.n908 B.n17 163.367
R1059 B.n908 B.n19 163.367
R1060 B.n904 B.n19 163.367
R1061 B.n904 B.n24 163.367
R1062 B.n900 B.n24 163.367
R1063 B.n900 B.n26 163.367
R1064 B.n896 B.n26 163.367
R1065 B.n896 B.n30 163.367
R1066 B.n892 B.n30 163.367
R1067 B.n892 B.n32 163.367
R1068 B.n888 B.n32 163.367
R1069 B.n888 B.n38 163.367
R1070 B.n884 B.n38 163.367
R1071 B.n884 B.n40 163.367
R1072 B.n880 B.n40 163.367
R1073 B.n880 B.n44 163.367
R1074 B.n876 B.n44 163.367
R1075 B.n876 B.n46 163.367
R1076 B.n872 B.n46 163.367
R1077 B.n872 B.n52 163.367
R1078 B.n868 B.n52 163.367
R1079 B.n868 B.n54 163.367
R1080 B.n864 B.n54 163.367
R1081 B.n864 B.n59 163.367
R1082 B.n860 B.n59 163.367
R1083 B.n860 B.n61 163.367
R1084 B.n856 B.n61 163.367
R1085 B.n856 B.n66 163.367
R1086 B.n852 B.n66 163.367
R1087 B.n852 B.n68 163.367
R1088 B.n848 B.n68 163.367
R1089 B.n848 B.n73 163.367
R1090 B.n844 B.n73 163.367
R1091 B.n844 B.n75 163.367
R1092 B.n840 B.n75 163.367
R1093 B.n840 B.n80 163.367
R1094 B.n836 B.n80 163.367
R1095 B.n836 B.n82 163.367
R1096 B.n832 B.n82 163.367
R1097 B.n832 B.n87 163.367
R1098 B.n828 B.n87 163.367
R1099 B.n828 B.n89 163.367
R1100 B.n824 B.n89 163.367
R1101 B.n824 B.n94 163.367
R1102 B.n137 B.t20 126.385
R1103 B.n436 B.t14 126.385
R1104 B.n140 B.t17 126.374
R1105 B.n433 B.t11 126.374
R1106 B.n592 B.n390 83.676
R1107 B.n818 B.n93 83.676
R1108 B.n820 B.n819 71.676
R1109 B.n142 B.n97 71.676
R1110 B.n146 B.n98 71.676
R1111 B.n150 B.n99 71.676
R1112 B.n154 B.n100 71.676
R1113 B.n158 B.n101 71.676
R1114 B.n162 B.n102 71.676
R1115 B.n166 B.n103 71.676
R1116 B.n170 B.n104 71.676
R1117 B.n174 B.n105 71.676
R1118 B.n178 B.n106 71.676
R1119 B.n182 B.n107 71.676
R1120 B.n186 B.n108 71.676
R1121 B.n190 B.n109 71.676
R1122 B.n194 B.n110 71.676
R1123 B.n198 B.n111 71.676
R1124 B.n202 B.n112 71.676
R1125 B.n206 B.n113 71.676
R1126 B.n211 B.n114 71.676
R1127 B.n215 B.n115 71.676
R1128 B.n219 B.n116 71.676
R1129 B.n223 B.n117 71.676
R1130 B.n227 B.n118 71.676
R1131 B.n231 B.n119 71.676
R1132 B.n235 B.n120 71.676
R1133 B.n239 B.n121 71.676
R1134 B.n243 B.n122 71.676
R1135 B.n247 B.n123 71.676
R1136 B.n251 B.n124 71.676
R1137 B.n255 B.n125 71.676
R1138 B.n259 B.n126 71.676
R1139 B.n263 B.n127 71.676
R1140 B.n267 B.n128 71.676
R1141 B.n271 B.n129 71.676
R1142 B.n275 B.n130 71.676
R1143 B.n279 B.n131 71.676
R1144 B.n283 B.n132 71.676
R1145 B.n287 B.n133 71.676
R1146 B.n291 B.n134 71.676
R1147 B.n135 B.n134 71.676
R1148 B.n290 B.n133 71.676
R1149 B.n286 B.n132 71.676
R1150 B.n282 B.n131 71.676
R1151 B.n278 B.n130 71.676
R1152 B.n274 B.n129 71.676
R1153 B.n270 B.n128 71.676
R1154 B.n266 B.n127 71.676
R1155 B.n262 B.n126 71.676
R1156 B.n258 B.n125 71.676
R1157 B.n254 B.n124 71.676
R1158 B.n250 B.n123 71.676
R1159 B.n246 B.n122 71.676
R1160 B.n242 B.n121 71.676
R1161 B.n238 B.n120 71.676
R1162 B.n234 B.n119 71.676
R1163 B.n230 B.n118 71.676
R1164 B.n226 B.n117 71.676
R1165 B.n222 B.n116 71.676
R1166 B.n218 B.n115 71.676
R1167 B.n214 B.n114 71.676
R1168 B.n210 B.n113 71.676
R1169 B.n205 B.n112 71.676
R1170 B.n201 B.n111 71.676
R1171 B.n197 B.n110 71.676
R1172 B.n193 B.n109 71.676
R1173 B.n189 B.n108 71.676
R1174 B.n185 B.n107 71.676
R1175 B.n181 B.n106 71.676
R1176 B.n177 B.n105 71.676
R1177 B.n173 B.n104 71.676
R1178 B.n169 B.n103 71.676
R1179 B.n165 B.n102 71.676
R1180 B.n161 B.n101 71.676
R1181 B.n157 B.n100 71.676
R1182 B.n153 B.n99 71.676
R1183 B.n149 B.n98 71.676
R1184 B.n145 B.n97 71.676
R1185 B.n819 B.n96 71.676
R1186 B.n594 B.n593 71.676
R1187 B.n432 B.n394 71.676
R1188 B.n586 B.n395 71.676
R1189 B.n582 B.n396 71.676
R1190 B.n578 B.n397 71.676
R1191 B.n574 B.n398 71.676
R1192 B.n570 B.n399 71.676
R1193 B.n566 B.n400 71.676
R1194 B.n562 B.n401 71.676
R1195 B.n558 B.n402 71.676
R1196 B.n554 B.n403 71.676
R1197 B.n550 B.n404 71.676
R1198 B.n546 B.n405 71.676
R1199 B.n542 B.n406 71.676
R1200 B.n538 B.n407 71.676
R1201 B.n534 B.n408 71.676
R1202 B.n530 B.n409 71.676
R1203 B.n526 B.n410 71.676
R1204 B.n522 B.n411 71.676
R1205 B.n518 B.n412 71.676
R1206 B.n514 B.n413 71.676
R1207 B.n510 B.n414 71.676
R1208 B.n505 B.n415 71.676
R1209 B.n501 B.n416 71.676
R1210 B.n497 B.n417 71.676
R1211 B.n493 B.n418 71.676
R1212 B.n489 B.n419 71.676
R1213 B.n485 B.n420 71.676
R1214 B.n481 B.n421 71.676
R1215 B.n477 B.n422 71.676
R1216 B.n473 B.n423 71.676
R1217 B.n469 B.n424 71.676
R1218 B.n465 B.n425 71.676
R1219 B.n461 B.n426 71.676
R1220 B.n457 B.n427 71.676
R1221 B.n453 B.n428 71.676
R1222 B.n449 B.n429 71.676
R1223 B.n445 B.n430 71.676
R1224 B.n441 B.n431 71.676
R1225 B.n593 B.n393 71.676
R1226 B.n587 B.n394 71.676
R1227 B.n583 B.n395 71.676
R1228 B.n579 B.n396 71.676
R1229 B.n575 B.n397 71.676
R1230 B.n571 B.n398 71.676
R1231 B.n567 B.n399 71.676
R1232 B.n563 B.n400 71.676
R1233 B.n559 B.n401 71.676
R1234 B.n555 B.n402 71.676
R1235 B.n551 B.n403 71.676
R1236 B.n547 B.n404 71.676
R1237 B.n543 B.n405 71.676
R1238 B.n539 B.n406 71.676
R1239 B.n535 B.n407 71.676
R1240 B.n531 B.n408 71.676
R1241 B.n527 B.n409 71.676
R1242 B.n523 B.n410 71.676
R1243 B.n519 B.n411 71.676
R1244 B.n515 B.n412 71.676
R1245 B.n511 B.n413 71.676
R1246 B.n506 B.n414 71.676
R1247 B.n502 B.n415 71.676
R1248 B.n498 B.n416 71.676
R1249 B.n494 B.n417 71.676
R1250 B.n490 B.n418 71.676
R1251 B.n486 B.n419 71.676
R1252 B.n482 B.n420 71.676
R1253 B.n478 B.n421 71.676
R1254 B.n474 B.n422 71.676
R1255 B.n470 B.n423 71.676
R1256 B.n466 B.n424 71.676
R1257 B.n462 B.n425 71.676
R1258 B.n458 B.n426 71.676
R1259 B.n454 B.n427 71.676
R1260 B.n450 B.n428 71.676
R1261 B.n446 B.n429 71.676
R1262 B.n442 B.n430 71.676
R1263 B.n438 B.n431 71.676
R1264 B.n926 B.n925 71.676
R1265 B.n926 B.n2 71.676
R1266 B.n138 B.t21 69.3669
R1267 B.n437 B.t13 69.3669
R1268 B.n141 B.t18 69.3552
R1269 B.n434 B.t10 69.3552
R1270 B.n208 B.n141 59.5399
R1271 B.n139 B.n138 59.5399
R1272 B.n508 B.n437 59.5399
R1273 B.n435 B.n434 59.5399
R1274 B.n141 B.n140 57.0187
R1275 B.n138 B.n137 57.0187
R1276 B.n437 B.n436 57.0187
R1277 B.n434 B.n433 57.0187
R1278 B.n599 B.n390 50.3539
R1279 B.n599 B.n386 50.3539
R1280 B.n605 B.n386 50.3539
R1281 B.n605 B.n382 50.3539
R1282 B.n611 B.n382 50.3539
R1283 B.n611 B.n378 50.3539
R1284 B.n617 B.n378 50.3539
R1285 B.n623 B.n374 50.3539
R1286 B.n623 B.n370 50.3539
R1287 B.n629 B.n370 50.3539
R1288 B.n629 B.n366 50.3539
R1289 B.n635 B.n366 50.3539
R1290 B.n635 B.n362 50.3539
R1291 B.n641 B.n362 50.3539
R1292 B.n641 B.n358 50.3539
R1293 B.n647 B.n358 50.3539
R1294 B.n647 B.n354 50.3539
R1295 B.n653 B.n354 50.3539
R1296 B.n659 B.n350 50.3539
R1297 B.n659 B.n346 50.3539
R1298 B.n665 B.n346 50.3539
R1299 B.n665 B.n342 50.3539
R1300 B.n671 B.n342 50.3539
R1301 B.n671 B.n338 50.3539
R1302 B.n678 B.n338 50.3539
R1303 B.n678 B.n677 50.3539
R1304 B.n684 B.n331 50.3539
R1305 B.n690 B.n331 50.3539
R1306 B.n690 B.n327 50.3539
R1307 B.n696 B.n327 50.3539
R1308 B.n696 B.n323 50.3539
R1309 B.n703 B.n323 50.3539
R1310 B.n703 B.n702 50.3539
R1311 B.n709 B.n316 50.3539
R1312 B.n715 B.n316 50.3539
R1313 B.n715 B.n312 50.3539
R1314 B.n721 B.n312 50.3539
R1315 B.n721 B.n308 50.3539
R1316 B.n727 B.n308 50.3539
R1317 B.n727 B.n304 50.3539
R1318 B.n733 B.n304 50.3539
R1319 B.n740 B.n300 50.3539
R1320 B.n740 B.n296 50.3539
R1321 B.n746 B.n296 50.3539
R1322 B.n746 B.n4 50.3539
R1323 B.n924 B.n4 50.3539
R1324 B.n924 B.n923 50.3539
R1325 B.n923 B.n922 50.3539
R1326 B.n922 B.n8 50.3539
R1327 B.n12 B.n8 50.3539
R1328 B.n915 B.n12 50.3539
R1329 B.n915 B.n914 50.3539
R1330 B.n913 B.n16 50.3539
R1331 B.n907 B.n16 50.3539
R1332 B.n907 B.n906 50.3539
R1333 B.n906 B.n905 50.3539
R1334 B.n905 B.n23 50.3539
R1335 B.n899 B.n23 50.3539
R1336 B.n899 B.n898 50.3539
R1337 B.n898 B.n897 50.3539
R1338 B.n891 B.n33 50.3539
R1339 B.n891 B.n890 50.3539
R1340 B.n890 B.n889 50.3539
R1341 B.n889 B.n37 50.3539
R1342 B.n883 B.n37 50.3539
R1343 B.n883 B.n882 50.3539
R1344 B.n882 B.n881 50.3539
R1345 B.n875 B.n47 50.3539
R1346 B.n875 B.n874 50.3539
R1347 B.n874 B.n873 50.3539
R1348 B.n873 B.n51 50.3539
R1349 B.n867 B.n51 50.3539
R1350 B.n867 B.n866 50.3539
R1351 B.n866 B.n865 50.3539
R1352 B.n865 B.n58 50.3539
R1353 B.n859 B.n858 50.3539
R1354 B.n858 B.n857 50.3539
R1355 B.n857 B.n65 50.3539
R1356 B.n851 B.n65 50.3539
R1357 B.n851 B.n850 50.3539
R1358 B.n850 B.n849 50.3539
R1359 B.n849 B.n72 50.3539
R1360 B.n843 B.n72 50.3539
R1361 B.n843 B.n842 50.3539
R1362 B.n842 B.n841 50.3539
R1363 B.n841 B.n79 50.3539
R1364 B.n835 B.n834 50.3539
R1365 B.n834 B.n833 50.3539
R1366 B.n833 B.n86 50.3539
R1367 B.n827 B.n86 50.3539
R1368 B.n827 B.n826 50.3539
R1369 B.n826 B.n825 50.3539
R1370 B.n825 B.n93 50.3539
R1371 B.n702 B.t4 46.6515
R1372 B.n33 B.t1 46.6515
R1373 B.n617 B.t9 39.2465
R1374 B.n835 B.t16 39.2465
R1375 B.n684 B.t6 36.2846
R1376 B.n881 B.t0 36.2846
R1377 B.n653 B.t3 31.8416
R1378 B.n859 B.t5 31.8416
R1379 B.n733 B.t2 28.8797
R1380 B.t7 B.n913 28.8797
R1381 B.n816 B.n815 28.5664
R1382 B.n596 B.n595 28.5664
R1383 B.n439 B.n388 28.5664
R1384 B.n822 B.n821 28.5664
R1385 B.t2 B.n300 21.4748
R1386 B.n914 B.t7 21.4748
R1387 B.t3 B.n350 18.5128
R1388 B.t5 B.n58 18.5128
R1389 B B.n927 18.0485
R1390 B.n677 B.t6 14.0698
R1391 B.n47 B.t0 14.0698
R1392 B.t9 B.n374 11.1079
R1393 B.t16 B.n79 11.1079
R1394 B.n597 B.n596 10.6151
R1395 B.n597 B.n384 10.6151
R1396 B.n607 B.n384 10.6151
R1397 B.n608 B.n607 10.6151
R1398 B.n609 B.n608 10.6151
R1399 B.n609 B.n376 10.6151
R1400 B.n619 B.n376 10.6151
R1401 B.n620 B.n619 10.6151
R1402 B.n621 B.n620 10.6151
R1403 B.n621 B.n368 10.6151
R1404 B.n631 B.n368 10.6151
R1405 B.n632 B.n631 10.6151
R1406 B.n633 B.n632 10.6151
R1407 B.n633 B.n360 10.6151
R1408 B.n643 B.n360 10.6151
R1409 B.n644 B.n643 10.6151
R1410 B.n645 B.n644 10.6151
R1411 B.n645 B.n352 10.6151
R1412 B.n655 B.n352 10.6151
R1413 B.n656 B.n655 10.6151
R1414 B.n657 B.n656 10.6151
R1415 B.n657 B.n344 10.6151
R1416 B.n667 B.n344 10.6151
R1417 B.n668 B.n667 10.6151
R1418 B.n669 B.n668 10.6151
R1419 B.n669 B.n336 10.6151
R1420 B.n680 B.n336 10.6151
R1421 B.n681 B.n680 10.6151
R1422 B.n682 B.n681 10.6151
R1423 B.n682 B.n329 10.6151
R1424 B.n692 B.n329 10.6151
R1425 B.n693 B.n692 10.6151
R1426 B.n694 B.n693 10.6151
R1427 B.n694 B.n321 10.6151
R1428 B.n705 B.n321 10.6151
R1429 B.n706 B.n705 10.6151
R1430 B.n707 B.n706 10.6151
R1431 B.n707 B.n314 10.6151
R1432 B.n717 B.n314 10.6151
R1433 B.n718 B.n717 10.6151
R1434 B.n719 B.n718 10.6151
R1435 B.n719 B.n306 10.6151
R1436 B.n729 B.n306 10.6151
R1437 B.n730 B.n729 10.6151
R1438 B.n731 B.n730 10.6151
R1439 B.n731 B.n298 10.6151
R1440 B.n742 B.n298 10.6151
R1441 B.n743 B.n742 10.6151
R1442 B.n744 B.n743 10.6151
R1443 B.n744 B.n0 10.6151
R1444 B.n595 B.n392 10.6151
R1445 B.n590 B.n392 10.6151
R1446 B.n590 B.n589 10.6151
R1447 B.n589 B.n588 10.6151
R1448 B.n588 B.n585 10.6151
R1449 B.n585 B.n584 10.6151
R1450 B.n584 B.n581 10.6151
R1451 B.n581 B.n580 10.6151
R1452 B.n580 B.n577 10.6151
R1453 B.n577 B.n576 10.6151
R1454 B.n576 B.n573 10.6151
R1455 B.n573 B.n572 10.6151
R1456 B.n572 B.n569 10.6151
R1457 B.n569 B.n568 10.6151
R1458 B.n568 B.n565 10.6151
R1459 B.n565 B.n564 10.6151
R1460 B.n564 B.n561 10.6151
R1461 B.n561 B.n560 10.6151
R1462 B.n560 B.n557 10.6151
R1463 B.n557 B.n556 10.6151
R1464 B.n556 B.n553 10.6151
R1465 B.n553 B.n552 10.6151
R1466 B.n552 B.n549 10.6151
R1467 B.n549 B.n548 10.6151
R1468 B.n548 B.n545 10.6151
R1469 B.n545 B.n544 10.6151
R1470 B.n544 B.n541 10.6151
R1471 B.n541 B.n540 10.6151
R1472 B.n540 B.n537 10.6151
R1473 B.n537 B.n536 10.6151
R1474 B.n536 B.n533 10.6151
R1475 B.n533 B.n532 10.6151
R1476 B.n532 B.n529 10.6151
R1477 B.n529 B.n528 10.6151
R1478 B.n525 B.n524 10.6151
R1479 B.n524 B.n521 10.6151
R1480 B.n521 B.n520 10.6151
R1481 B.n520 B.n517 10.6151
R1482 B.n517 B.n516 10.6151
R1483 B.n516 B.n513 10.6151
R1484 B.n513 B.n512 10.6151
R1485 B.n512 B.n509 10.6151
R1486 B.n507 B.n504 10.6151
R1487 B.n504 B.n503 10.6151
R1488 B.n503 B.n500 10.6151
R1489 B.n500 B.n499 10.6151
R1490 B.n499 B.n496 10.6151
R1491 B.n496 B.n495 10.6151
R1492 B.n495 B.n492 10.6151
R1493 B.n492 B.n491 10.6151
R1494 B.n491 B.n488 10.6151
R1495 B.n488 B.n487 10.6151
R1496 B.n487 B.n484 10.6151
R1497 B.n484 B.n483 10.6151
R1498 B.n483 B.n480 10.6151
R1499 B.n480 B.n479 10.6151
R1500 B.n479 B.n476 10.6151
R1501 B.n476 B.n475 10.6151
R1502 B.n475 B.n472 10.6151
R1503 B.n472 B.n471 10.6151
R1504 B.n471 B.n468 10.6151
R1505 B.n468 B.n467 10.6151
R1506 B.n467 B.n464 10.6151
R1507 B.n464 B.n463 10.6151
R1508 B.n463 B.n460 10.6151
R1509 B.n460 B.n459 10.6151
R1510 B.n459 B.n456 10.6151
R1511 B.n456 B.n455 10.6151
R1512 B.n455 B.n452 10.6151
R1513 B.n452 B.n451 10.6151
R1514 B.n451 B.n448 10.6151
R1515 B.n448 B.n447 10.6151
R1516 B.n447 B.n444 10.6151
R1517 B.n444 B.n443 10.6151
R1518 B.n443 B.n440 10.6151
R1519 B.n440 B.n439 10.6151
R1520 B.n601 B.n388 10.6151
R1521 B.n602 B.n601 10.6151
R1522 B.n603 B.n602 10.6151
R1523 B.n603 B.n380 10.6151
R1524 B.n613 B.n380 10.6151
R1525 B.n614 B.n613 10.6151
R1526 B.n615 B.n614 10.6151
R1527 B.n615 B.n372 10.6151
R1528 B.n625 B.n372 10.6151
R1529 B.n626 B.n625 10.6151
R1530 B.n627 B.n626 10.6151
R1531 B.n627 B.n364 10.6151
R1532 B.n637 B.n364 10.6151
R1533 B.n638 B.n637 10.6151
R1534 B.n639 B.n638 10.6151
R1535 B.n639 B.n356 10.6151
R1536 B.n649 B.n356 10.6151
R1537 B.n650 B.n649 10.6151
R1538 B.n651 B.n650 10.6151
R1539 B.n651 B.n348 10.6151
R1540 B.n661 B.n348 10.6151
R1541 B.n662 B.n661 10.6151
R1542 B.n663 B.n662 10.6151
R1543 B.n663 B.n340 10.6151
R1544 B.n673 B.n340 10.6151
R1545 B.n674 B.n673 10.6151
R1546 B.n675 B.n674 10.6151
R1547 B.n675 B.n333 10.6151
R1548 B.n686 B.n333 10.6151
R1549 B.n687 B.n686 10.6151
R1550 B.n688 B.n687 10.6151
R1551 B.n688 B.n325 10.6151
R1552 B.n698 B.n325 10.6151
R1553 B.n699 B.n698 10.6151
R1554 B.n700 B.n699 10.6151
R1555 B.n700 B.n318 10.6151
R1556 B.n711 B.n318 10.6151
R1557 B.n712 B.n711 10.6151
R1558 B.n713 B.n712 10.6151
R1559 B.n713 B.n310 10.6151
R1560 B.n723 B.n310 10.6151
R1561 B.n724 B.n723 10.6151
R1562 B.n725 B.n724 10.6151
R1563 B.n725 B.n302 10.6151
R1564 B.n735 B.n302 10.6151
R1565 B.n736 B.n735 10.6151
R1566 B.n738 B.n736 10.6151
R1567 B.n738 B.n737 10.6151
R1568 B.n737 B.n294 10.6151
R1569 B.n749 B.n294 10.6151
R1570 B.n750 B.n749 10.6151
R1571 B.n751 B.n750 10.6151
R1572 B.n752 B.n751 10.6151
R1573 B.n753 B.n752 10.6151
R1574 B.n756 B.n753 10.6151
R1575 B.n757 B.n756 10.6151
R1576 B.n758 B.n757 10.6151
R1577 B.n759 B.n758 10.6151
R1578 B.n761 B.n759 10.6151
R1579 B.n762 B.n761 10.6151
R1580 B.n763 B.n762 10.6151
R1581 B.n764 B.n763 10.6151
R1582 B.n766 B.n764 10.6151
R1583 B.n767 B.n766 10.6151
R1584 B.n768 B.n767 10.6151
R1585 B.n769 B.n768 10.6151
R1586 B.n771 B.n769 10.6151
R1587 B.n772 B.n771 10.6151
R1588 B.n773 B.n772 10.6151
R1589 B.n774 B.n773 10.6151
R1590 B.n776 B.n774 10.6151
R1591 B.n777 B.n776 10.6151
R1592 B.n778 B.n777 10.6151
R1593 B.n779 B.n778 10.6151
R1594 B.n781 B.n779 10.6151
R1595 B.n782 B.n781 10.6151
R1596 B.n783 B.n782 10.6151
R1597 B.n784 B.n783 10.6151
R1598 B.n786 B.n784 10.6151
R1599 B.n787 B.n786 10.6151
R1600 B.n788 B.n787 10.6151
R1601 B.n789 B.n788 10.6151
R1602 B.n791 B.n789 10.6151
R1603 B.n792 B.n791 10.6151
R1604 B.n793 B.n792 10.6151
R1605 B.n794 B.n793 10.6151
R1606 B.n796 B.n794 10.6151
R1607 B.n797 B.n796 10.6151
R1608 B.n798 B.n797 10.6151
R1609 B.n799 B.n798 10.6151
R1610 B.n801 B.n799 10.6151
R1611 B.n802 B.n801 10.6151
R1612 B.n803 B.n802 10.6151
R1613 B.n804 B.n803 10.6151
R1614 B.n806 B.n804 10.6151
R1615 B.n807 B.n806 10.6151
R1616 B.n808 B.n807 10.6151
R1617 B.n809 B.n808 10.6151
R1618 B.n811 B.n809 10.6151
R1619 B.n812 B.n811 10.6151
R1620 B.n813 B.n812 10.6151
R1621 B.n814 B.n813 10.6151
R1622 B.n815 B.n814 10.6151
R1623 B.n919 B.n1 10.6151
R1624 B.n919 B.n918 10.6151
R1625 B.n918 B.n917 10.6151
R1626 B.n917 B.n10 10.6151
R1627 B.n911 B.n10 10.6151
R1628 B.n911 B.n910 10.6151
R1629 B.n910 B.n909 10.6151
R1630 B.n909 B.n18 10.6151
R1631 B.n903 B.n18 10.6151
R1632 B.n903 B.n902 10.6151
R1633 B.n902 B.n901 10.6151
R1634 B.n901 B.n25 10.6151
R1635 B.n895 B.n25 10.6151
R1636 B.n895 B.n894 10.6151
R1637 B.n894 B.n893 10.6151
R1638 B.n893 B.n31 10.6151
R1639 B.n887 B.n31 10.6151
R1640 B.n887 B.n886 10.6151
R1641 B.n886 B.n885 10.6151
R1642 B.n885 B.n39 10.6151
R1643 B.n879 B.n39 10.6151
R1644 B.n879 B.n878 10.6151
R1645 B.n878 B.n877 10.6151
R1646 B.n877 B.n45 10.6151
R1647 B.n871 B.n45 10.6151
R1648 B.n871 B.n870 10.6151
R1649 B.n870 B.n869 10.6151
R1650 B.n869 B.n53 10.6151
R1651 B.n863 B.n53 10.6151
R1652 B.n863 B.n862 10.6151
R1653 B.n862 B.n861 10.6151
R1654 B.n861 B.n60 10.6151
R1655 B.n855 B.n60 10.6151
R1656 B.n855 B.n854 10.6151
R1657 B.n854 B.n853 10.6151
R1658 B.n853 B.n67 10.6151
R1659 B.n847 B.n67 10.6151
R1660 B.n847 B.n846 10.6151
R1661 B.n846 B.n845 10.6151
R1662 B.n845 B.n74 10.6151
R1663 B.n839 B.n74 10.6151
R1664 B.n839 B.n838 10.6151
R1665 B.n838 B.n837 10.6151
R1666 B.n837 B.n81 10.6151
R1667 B.n831 B.n81 10.6151
R1668 B.n831 B.n830 10.6151
R1669 B.n830 B.n829 10.6151
R1670 B.n829 B.n88 10.6151
R1671 B.n823 B.n88 10.6151
R1672 B.n823 B.n822 10.6151
R1673 B.n821 B.n95 10.6151
R1674 B.n143 B.n95 10.6151
R1675 B.n144 B.n143 10.6151
R1676 B.n147 B.n144 10.6151
R1677 B.n148 B.n147 10.6151
R1678 B.n151 B.n148 10.6151
R1679 B.n152 B.n151 10.6151
R1680 B.n155 B.n152 10.6151
R1681 B.n156 B.n155 10.6151
R1682 B.n159 B.n156 10.6151
R1683 B.n160 B.n159 10.6151
R1684 B.n163 B.n160 10.6151
R1685 B.n164 B.n163 10.6151
R1686 B.n167 B.n164 10.6151
R1687 B.n168 B.n167 10.6151
R1688 B.n171 B.n168 10.6151
R1689 B.n172 B.n171 10.6151
R1690 B.n175 B.n172 10.6151
R1691 B.n176 B.n175 10.6151
R1692 B.n179 B.n176 10.6151
R1693 B.n180 B.n179 10.6151
R1694 B.n183 B.n180 10.6151
R1695 B.n184 B.n183 10.6151
R1696 B.n187 B.n184 10.6151
R1697 B.n188 B.n187 10.6151
R1698 B.n191 B.n188 10.6151
R1699 B.n192 B.n191 10.6151
R1700 B.n195 B.n192 10.6151
R1701 B.n196 B.n195 10.6151
R1702 B.n199 B.n196 10.6151
R1703 B.n200 B.n199 10.6151
R1704 B.n203 B.n200 10.6151
R1705 B.n204 B.n203 10.6151
R1706 B.n207 B.n204 10.6151
R1707 B.n212 B.n209 10.6151
R1708 B.n213 B.n212 10.6151
R1709 B.n216 B.n213 10.6151
R1710 B.n217 B.n216 10.6151
R1711 B.n220 B.n217 10.6151
R1712 B.n221 B.n220 10.6151
R1713 B.n224 B.n221 10.6151
R1714 B.n225 B.n224 10.6151
R1715 B.n229 B.n228 10.6151
R1716 B.n232 B.n229 10.6151
R1717 B.n233 B.n232 10.6151
R1718 B.n236 B.n233 10.6151
R1719 B.n237 B.n236 10.6151
R1720 B.n240 B.n237 10.6151
R1721 B.n241 B.n240 10.6151
R1722 B.n244 B.n241 10.6151
R1723 B.n245 B.n244 10.6151
R1724 B.n248 B.n245 10.6151
R1725 B.n249 B.n248 10.6151
R1726 B.n252 B.n249 10.6151
R1727 B.n253 B.n252 10.6151
R1728 B.n256 B.n253 10.6151
R1729 B.n257 B.n256 10.6151
R1730 B.n260 B.n257 10.6151
R1731 B.n261 B.n260 10.6151
R1732 B.n264 B.n261 10.6151
R1733 B.n265 B.n264 10.6151
R1734 B.n268 B.n265 10.6151
R1735 B.n269 B.n268 10.6151
R1736 B.n272 B.n269 10.6151
R1737 B.n273 B.n272 10.6151
R1738 B.n276 B.n273 10.6151
R1739 B.n277 B.n276 10.6151
R1740 B.n280 B.n277 10.6151
R1741 B.n281 B.n280 10.6151
R1742 B.n284 B.n281 10.6151
R1743 B.n285 B.n284 10.6151
R1744 B.n288 B.n285 10.6151
R1745 B.n289 B.n288 10.6151
R1746 B.n292 B.n289 10.6151
R1747 B.n293 B.n292 10.6151
R1748 B.n816 B.n293 10.6151
R1749 B.n927 B.n0 8.11757
R1750 B.n927 B.n1 8.11757
R1751 B.n525 B.n435 6.5566
R1752 B.n509 B.n508 6.5566
R1753 B.n209 B.n208 6.5566
R1754 B.n225 B.n139 6.5566
R1755 B.n528 B.n435 4.05904
R1756 B.n508 B.n507 4.05904
R1757 B.n208 B.n207 4.05904
R1758 B.n228 B.n139 4.05904
R1759 B.n709 B.t4 3.70296
R1760 B.n897 B.t1 3.70296
R1761 VN.n55 VN.n29 161.3
R1762 VN.n54 VN.n53 161.3
R1763 VN.n52 VN.n30 161.3
R1764 VN.n51 VN.n50 161.3
R1765 VN.n49 VN.n31 161.3
R1766 VN.n48 VN.n47 161.3
R1767 VN.n46 VN.n45 161.3
R1768 VN.n44 VN.n33 161.3
R1769 VN.n43 VN.n42 161.3
R1770 VN.n41 VN.n34 161.3
R1771 VN.n40 VN.n39 161.3
R1772 VN.n38 VN.n35 161.3
R1773 VN.n26 VN.n0 161.3
R1774 VN.n25 VN.n24 161.3
R1775 VN.n23 VN.n1 161.3
R1776 VN.n22 VN.n21 161.3
R1777 VN.n20 VN.n2 161.3
R1778 VN.n19 VN.n18 161.3
R1779 VN.n17 VN.n16 161.3
R1780 VN.n15 VN.n4 161.3
R1781 VN.n14 VN.n13 161.3
R1782 VN.n12 VN.n5 161.3
R1783 VN.n11 VN.n10 161.3
R1784 VN.n9 VN.n6 161.3
R1785 VN.n7 VN.t7 121.51
R1786 VN.n36 VN.t2 121.51
R1787 VN.n28 VN.n27 103.038
R1788 VN.n57 VN.n56 103.038
R1789 VN.n8 VN.t1 88.4595
R1790 VN.n3 VN.t4 88.4595
R1791 VN.n27 VN.t6 88.4595
R1792 VN.n37 VN.t3 88.4595
R1793 VN.n32 VN.t5 88.4595
R1794 VN.n56 VN.t0 88.4595
R1795 VN.n8 VN.n7 61.7254
R1796 VN.n37 VN.n36 61.7254
R1797 VN.n14 VN.n5 56.5617
R1798 VN.n21 VN.n1 56.5617
R1799 VN.n43 VN.n34 56.5617
R1800 VN.n50 VN.n30 56.5617
R1801 VN VN.n57 49.377
R1802 VN.n10 VN.n9 24.5923
R1803 VN.n10 VN.n5 24.5923
R1804 VN.n15 VN.n14 24.5923
R1805 VN.n16 VN.n15 24.5923
R1806 VN.n20 VN.n19 24.5923
R1807 VN.n21 VN.n20 24.5923
R1808 VN.n25 VN.n1 24.5923
R1809 VN.n26 VN.n25 24.5923
R1810 VN.n39 VN.n34 24.5923
R1811 VN.n39 VN.n38 24.5923
R1812 VN.n50 VN.n49 24.5923
R1813 VN.n49 VN.n48 24.5923
R1814 VN.n45 VN.n44 24.5923
R1815 VN.n44 VN.n43 24.5923
R1816 VN.n55 VN.n54 24.5923
R1817 VN.n54 VN.n30 24.5923
R1818 VN.n19 VN.n3 13.7719
R1819 VN.n48 VN.n32 13.7719
R1820 VN.n9 VN.n8 10.8209
R1821 VN.n16 VN.n3 10.8209
R1822 VN.n38 VN.n37 10.8209
R1823 VN.n45 VN.n32 10.8209
R1824 VN.n27 VN.n26 7.86989
R1825 VN.n56 VN.n55 7.86989
R1826 VN.n36 VN.n35 6.96699
R1827 VN.n7 VN.n6 6.96699
R1828 VN.n57 VN.n29 0.278335
R1829 VN.n28 VN.n0 0.278335
R1830 VN.n53 VN.n29 0.189894
R1831 VN.n53 VN.n52 0.189894
R1832 VN.n52 VN.n51 0.189894
R1833 VN.n51 VN.n31 0.189894
R1834 VN.n47 VN.n31 0.189894
R1835 VN.n47 VN.n46 0.189894
R1836 VN.n46 VN.n33 0.189894
R1837 VN.n42 VN.n33 0.189894
R1838 VN.n42 VN.n41 0.189894
R1839 VN.n41 VN.n40 0.189894
R1840 VN.n40 VN.n35 0.189894
R1841 VN.n11 VN.n6 0.189894
R1842 VN.n12 VN.n11 0.189894
R1843 VN.n13 VN.n12 0.189894
R1844 VN.n13 VN.n4 0.189894
R1845 VN.n17 VN.n4 0.189894
R1846 VN.n18 VN.n17 0.189894
R1847 VN.n18 VN.n2 0.189894
R1848 VN.n22 VN.n2 0.189894
R1849 VN.n23 VN.n22 0.189894
R1850 VN.n24 VN.n23 0.189894
R1851 VN.n24 VN.n0 0.189894
R1852 VN VN.n28 0.153485
R1853 VDD2.n2 VDD2.n1 63.6359
R1854 VDD2.n2 VDD2.n0 63.6359
R1855 VDD2 VDD2.n5 63.6331
R1856 VDD2.n4 VDD2.n3 62.4242
R1857 VDD2.n4 VDD2.n2 43.3791
R1858 VDD2.n5 VDD2.t4 2.06731
R1859 VDD2.n5 VDD2.t5 2.06731
R1860 VDD2.n3 VDD2.t7 2.06731
R1861 VDD2.n3 VDD2.t2 2.06731
R1862 VDD2.n1 VDD2.t3 2.06731
R1863 VDD2.n1 VDD2.t1 2.06731
R1864 VDD2.n0 VDD2.t0 2.06731
R1865 VDD2.n0 VDD2.t6 2.06731
R1866 VDD2 VDD2.n4 1.32593
C0 VTAIL VDD2 7.32231f
C1 VTAIL VN 7.53835f
C2 VDD1 VTAIL 7.26783f
C3 VN VDD2 7.03057f
C4 VDD1 VDD2 1.78332f
C5 VTAIL VP 7.55245f
C6 VDD2 VP 0.521174f
C7 VDD1 VN 0.152185f
C8 VN VP 7.22086f
C9 VDD1 VP 7.39816f
C10 VDD2 B 5.165053f
C11 VDD1 B 5.609174f
C12 VTAIL B 9.05217f
C13 VN B 15.331161f
C14 VP B 13.956058f
C15 VDD2.t0 B 0.182976f
C16 VDD2.t6 B 0.182976f
C17 VDD2.n0 B 1.61533f
C18 VDD2.t3 B 0.182976f
C19 VDD2.t1 B 0.182976f
C20 VDD2.n1 B 1.61533f
C21 VDD2.n2 B 3.02472f
C22 VDD2.t7 B 0.182976f
C23 VDD2.t2 B 0.182976f
C24 VDD2.n3 B 1.60583f
C25 VDD2.n4 B 2.67376f
C26 VDD2.t4 B 0.182976f
C27 VDD2.t5 B 0.182976f
C28 VDD2.n5 B 1.61529f
C29 VN.n0 B 0.029872f
C30 VN.t6 B 1.53256f
C31 VN.n1 B 0.036701f
C32 VN.n2 B 0.022659f
C33 VN.t4 B 1.53256f
C34 VN.n3 B 0.550012f
C35 VN.n4 B 0.022659f
C36 VN.n5 B 0.032939f
C37 VN.n6 B 0.219164f
C38 VN.t1 B 1.53256f
C39 VN.t7 B 1.72f
C40 VN.n7 B 0.595518f
C41 VN.n8 B 0.613808f
C42 VN.n9 B 0.030403f
C43 VN.n10 B 0.04202f
C44 VN.n11 B 0.022659f
C45 VN.n12 B 0.022659f
C46 VN.n13 B 0.022659f
C47 VN.n14 B 0.032939f
C48 VN.n15 B 0.04202f
C49 VN.n16 B 0.030403f
C50 VN.n17 B 0.022659f
C51 VN.n18 B 0.022659f
C52 VN.n19 B 0.032893f
C53 VN.n20 B 0.04202f
C54 VN.n21 B 0.029177f
C55 VN.n22 B 0.022659f
C56 VN.n23 B 0.022659f
C57 VN.n24 B 0.022659f
C58 VN.n25 B 0.04202f
C59 VN.n26 B 0.027914f
C60 VN.n27 B 0.623163f
C61 VN.n28 B 0.038135f
C62 VN.n29 B 0.029872f
C63 VN.t0 B 1.53256f
C64 VN.n30 B 0.036701f
C65 VN.n31 B 0.022659f
C66 VN.t5 B 1.53256f
C67 VN.n32 B 0.550012f
C68 VN.n33 B 0.022659f
C69 VN.n34 B 0.032939f
C70 VN.n35 B 0.219164f
C71 VN.t3 B 1.53256f
C72 VN.t2 B 1.72f
C73 VN.n36 B 0.595518f
C74 VN.n37 B 0.613808f
C75 VN.n38 B 0.030403f
C76 VN.n39 B 0.04202f
C77 VN.n40 B 0.022659f
C78 VN.n41 B 0.022659f
C79 VN.n42 B 0.022659f
C80 VN.n43 B 0.032939f
C81 VN.n44 B 0.04202f
C82 VN.n45 B 0.030403f
C83 VN.n46 B 0.022659f
C84 VN.n47 B 0.022659f
C85 VN.n48 B 0.032893f
C86 VN.n49 B 0.04202f
C87 VN.n50 B 0.029177f
C88 VN.n51 B 0.022659f
C89 VN.n52 B 0.022659f
C90 VN.n53 B 0.022659f
C91 VN.n54 B 0.04202f
C92 VN.n55 B 0.027914f
C93 VN.n56 B 0.623163f
C94 VN.n57 B 1.24072f
C95 VTAIL.t1 B 0.156735f
C96 VTAIL.t0 B 0.156735f
C97 VTAIL.n0 B 1.31553f
C98 VTAIL.n1 B 0.373329f
C99 VTAIL.t15 B 1.67441f
C100 VTAIL.n2 B 0.469365f
C101 VTAIL.t12 B 1.67441f
C102 VTAIL.n3 B 0.469365f
C103 VTAIL.t9 B 0.156735f
C104 VTAIL.t11 B 0.156735f
C105 VTAIL.n4 B 1.31553f
C106 VTAIL.n5 B 0.538527f
C107 VTAIL.t13 B 1.67441f
C108 VTAIL.n6 B 1.43928f
C109 VTAIL.t3 B 1.67443f
C110 VTAIL.n7 B 1.43927f
C111 VTAIL.t6 B 0.156735f
C112 VTAIL.t4 B 0.156735f
C113 VTAIL.n8 B 1.31553f
C114 VTAIL.n9 B 0.538523f
C115 VTAIL.t2 B 1.67443f
C116 VTAIL.n10 B 0.469353f
C117 VTAIL.t10 B 1.67443f
C118 VTAIL.n11 B 0.469353f
C119 VTAIL.t7 B 0.156735f
C120 VTAIL.t14 B 0.156735f
C121 VTAIL.n12 B 1.31553f
C122 VTAIL.n13 B 0.538523f
C123 VTAIL.t8 B 1.67441f
C124 VTAIL.n14 B 1.43928f
C125 VTAIL.t5 B 1.67441f
C126 VTAIL.n15 B 1.4354f
C127 VDD1.t1 B 0.186928f
C128 VDD1.t2 B 0.186928f
C129 VDD1.n0 B 1.65128f
C130 VDD1.t5 B 0.186928f
C131 VDD1.t4 B 0.186928f
C132 VDD1.n1 B 1.65021f
C133 VDD1.t0 B 0.186928f
C134 VDD1.t7 B 0.186928f
C135 VDD1.n2 B 1.65021f
C136 VDD1.n3 B 3.14154f
C137 VDD1.t3 B 0.186928f
C138 VDD1.t6 B 0.186928f
C139 VDD1.n4 B 1.6405f
C140 VDD1.n5 B 2.76194f
C141 VP.n0 B 0.030606f
C142 VP.t2 B 1.57017f
C143 VP.n1 B 0.037601f
C144 VP.n2 B 0.023216f
C145 VP.t3 B 1.57017f
C146 VP.n3 B 0.563512f
C147 VP.n4 B 0.023216f
C148 VP.n5 B 0.033748f
C149 VP.n6 B 0.023216f
C150 VP.t5 B 1.57017f
C151 VP.n7 B 0.043051f
C152 VP.n8 B 0.023216f
C153 VP.n9 B 0.028599f
C154 VP.n10 B 0.030606f
C155 VP.t6 B 1.57017f
C156 VP.n11 B 0.037601f
C157 VP.n12 B 0.023216f
C158 VP.t0 B 1.57017f
C159 VP.n13 B 0.563512f
C160 VP.n14 B 0.023216f
C161 VP.n15 B 0.033748f
C162 VP.n16 B 0.224543f
C163 VP.t7 B 1.57017f
C164 VP.t4 B 1.76222f
C165 VP.n17 B 0.610135f
C166 VP.n18 B 0.628874f
C167 VP.n19 B 0.031149f
C168 VP.n20 B 0.043051f
C169 VP.n21 B 0.023216f
C170 VP.n22 B 0.023216f
C171 VP.n23 B 0.023216f
C172 VP.n24 B 0.033748f
C173 VP.n25 B 0.043051f
C174 VP.n26 B 0.031149f
C175 VP.n27 B 0.023216f
C176 VP.n28 B 0.023216f
C177 VP.n29 B 0.0337f
C178 VP.n30 B 0.043051f
C179 VP.n31 B 0.029894f
C180 VP.n32 B 0.023216f
C181 VP.n33 B 0.023216f
C182 VP.n34 B 0.023216f
C183 VP.n35 B 0.043051f
C184 VP.n36 B 0.028599f
C185 VP.n37 B 0.638458f
C186 VP.n38 B 1.25866f
C187 VP.t1 B 1.57017f
C188 VP.n39 B 0.638458f
C189 VP.n40 B 1.27571f
C190 VP.n41 B 0.030606f
C191 VP.n42 B 0.023216f
C192 VP.n43 B 0.043051f
C193 VP.n44 B 0.037601f
C194 VP.n45 B 0.029894f
C195 VP.n46 B 0.023216f
C196 VP.n47 B 0.023216f
C197 VP.n48 B 0.023216f
C198 VP.n49 B 0.0337f
C199 VP.n50 B 0.563512f
C200 VP.n51 B 0.031149f
C201 VP.n52 B 0.043051f
C202 VP.n53 B 0.023216f
C203 VP.n54 B 0.023216f
C204 VP.n55 B 0.023216f
C205 VP.n56 B 0.033748f
C206 VP.n57 B 0.043051f
C207 VP.n58 B 0.031149f
C208 VP.n59 B 0.023216f
C209 VP.n60 B 0.023216f
C210 VP.n61 B 0.0337f
C211 VP.n62 B 0.043051f
C212 VP.n63 B 0.029894f
C213 VP.n64 B 0.023216f
C214 VP.n65 B 0.023216f
C215 VP.n66 B 0.023216f
C216 VP.n67 B 0.043051f
C217 VP.n68 B 0.028599f
C218 VP.n69 B 0.638458f
C219 VP.n70 B 0.039071f
.ends

