* NGSPICE file created from diff_pair_sample_1174.ext - technology: sky130A

.subckt diff_pair_sample_1174 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X1 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0 ps=0 w=4.93 l=1.25
X2 VDD1.t9 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=1.9227 ps=10.64 w=4.93 l=1.25
X3 VTAIL.t16 VN.t1 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X4 VDD1.t8 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X5 VTAIL.t15 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X6 VDD1.t7 VP.t2 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=1.9227 ps=10.64 w=4.93 l=1.25
X7 VDD2.t3 VN.t3 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X8 VDD2.t6 VN.t4 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X9 VTAIL.t6 VP.t3 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X10 VDD1.t5 VP.t4 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0.81345 ps=5.26 w=4.93 l=1.25
X11 VTAIL.t5 VP.t5 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X12 VTAIL.t12 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X13 VDD2.t1 VN.t6 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=1.9227 ps=10.64 w=4.93 l=1.25
X14 VDD2.t4 VN.t7 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0.81345 ps=5.26 w=4.93 l=1.25
X15 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0 ps=0 w=4.93 l=1.25
X16 VDD1.t3 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X17 VDD1.t2 VP.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0.81345 ps=5.26 w=4.93 l=1.25
X18 VDD2.t0 VN.t8 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=1.9227 ps=10.64 w=4.93 l=1.25
X19 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X20 VTAIL.t3 VP.t9 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.81345 pd=5.26 as=0.81345 ps=5.26 w=4.93 l=1.25
X21 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0 ps=0 w=4.93 l=1.25
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0 ps=0 w=4.93 l=1.25
X23 VDD2.t9 VN.t9 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9227 pd=10.64 as=0.81345 ps=5.26 w=4.93 l=1.25
R0 VN.n41 VN.n22 161.3
R1 VN.n40 VN.n39 161.3
R2 VN.n38 VN.n37 161.3
R3 VN.n36 VN.n24 161.3
R4 VN.n35 VN.n34 161.3
R5 VN.n33 VN.n32 161.3
R6 VN.n31 VN.n26 161.3
R7 VN.n30 VN.n29 161.3
R8 VN.n19 VN.n0 161.3
R9 VN.n18 VN.n17 161.3
R10 VN.n16 VN.n15 161.3
R11 VN.n14 VN.n2 161.3
R12 VN.n13 VN.n12 161.3
R13 VN.n11 VN.n10 161.3
R14 VN.n9 VN.n4 161.3
R15 VN.n8 VN.n7 161.3
R16 VN.n6 VN.t9 147.857
R17 VN.n28 VN.t8 147.857
R18 VN.n20 VN.t6 126.671
R19 VN.n42 VN.t7 126.671
R20 VN.n5 VN.t0 95.0509
R21 VN.n3 VN.t4 95.0509
R22 VN.n1 VN.t1 95.0509
R23 VN.n27 VN.t5 95.0509
R24 VN.n25 VN.t3 95.0509
R25 VN.n23 VN.t2 95.0509
R26 VN.n43 VN.n42 80.6037
R27 VN.n21 VN.n20 80.6037
R28 VN.n9 VN.n8 44.3785
R29 VN.n15 VN.n14 44.3785
R30 VN.n31 VN.n30 44.3785
R31 VN.n37 VN.n36 44.3785
R32 VN.n20 VN.n19 41.6278
R33 VN.n42 VN.n41 41.6278
R34 VN VN.n43 40.9157
R35 VN.n6 VN.n5 40.893
R36 VN.n28 VN.n27 40.893
R37 VN.n10 VN.n9 36.6083
R38 VN.n14 VN.n13 36.6083
R39 VN.n32 VN.n31 36.6083
R40 VN.n36 VN.n35 36.6083
R41 VN.n19 VN.n18 28.8382
R42 VN.n41 VN.n40 28.8382
R43 VN.n29 VN.n28 28.8325
R44 VN.n7 VN.n6 28.8325
R45 VN.n8 VN.n5 16.1487
R46 VN.n15 VN.n1 16.1487
R47 VN.n30 VN.n27 16.1487
R48 VN.n37 VN.n23 16.1487
R49 VN.n10 VN.n3 12.234
R50 VN.n13 VN.n3 12.234
R51 VN.n35 VN.n25 12.234
R52 VN.n32 VN.n25 12.234
R53 VN.n18 VN.n1 8.31928
R54 VN.n40 VN.n23 8.31928
R55 VN.n43 VN.n22 0.285035
R56 VN.n21 VN.n0 0.285035
R57 VN.n39 VN.n22 0.189894
R58 VN.n39 VN.n38 0.189894
R59 VN.n38 VN.n24 0.189894
R60 VN.n34 VN.n24 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n26 0.189894
R63 VN.n29 VN.n26 0.189894
R64 VN.n7 VN.n4 0.189894
R65 VN.n11 VN.n4 0.189894
R66 VN.n12 VN.n11 0.189894
R67 VN.n12 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n17 VN.n0 0.189894
R71 VN VN.n21 0.146778
R72 VDD2.n1 VDD2.t9 75.1392
R73 VDD2.n4 VDD2.t4 73.7772
R74 VDD2.n3 VDD2.n2 70.727
R75 VDD2 VDD2.n7 70.7242
R76 VDD2.n6 VDD2.n5 69.761
R77 VDD2.n1 VDD2.n0 69.7608
R78 VDD2.n4 VDD2.n3 34.4351
R79 VDD2.n7 VDD2.t2 4.01673
R80 VDD2.n7 VDD2.t0 4.01673
R81 VDD2.n5 VDD2.t5 4.01673
R82 VDD2.n5 VDD2.t3 4.01673
R83 VDD2.n2 VDD2.t7 4.01673
R84 VDD2.n2 VDD2.t1 4.01673
R85 VDD2.n0 VDD2.t8 4.01673
R86 VDD2.n0 VDD2.t6 4.01673
R87 VDD2.n6 VDD2.n4 1.36257
R88 VDD2 VDD2.n6 0.399207
R89 VDD2.n3 VDD2.n1 0.285671
R90 VTAIL.n11 VTAIL.t9 57.0984
R91 VTAIL.n17 VTAIL.t11 57.0983
R92 VTAIL.n2 VTAIL.t0 57.0983
R93 VTAIL.n16 VTAIL.t18 57.0983
R94 VTAIL.n15 VTAIL.n14 53.0822
R95 VTAIL.n13 VTAIL.n12 53.0822
R96 VTAIL.n10 VTAIL.n9 53.0822
R97 VTAIL.n8 VTAIL.n7 53.0822
R98 VTAIL.n19 VTAIL.n18 53.082
R99 VTAIL.n1 VTAIL.n0 53.082
R100 VTAIL.n4 VTAIL.n3 53.082
R101 VTAIL.n6 VTAIL.n5 53.082
R102 VTAIL.n8 VTAIL.n6 19.341
R103 VTAIL.n17 VTAIL.n16 17.9789
R104 VTAIL.n18 VTAIL.t13 4.01673
R105 VTAIL.n18 VTAIL.t16 4.01673
R106 VTAIL.n0 VTAIL.t8 4.01673
R107 VTAIL.n0 VTAIL.t17 4.01673
R108 VTAIL.n3 VTAIL.t2 4.01673
R109 VTAIL.n3 VTAIL.t1 4.01673
R110 VTAIL.n5 VTAIL.t19 4.01673
R111 VTAIL.n5 VTAIL.t6 4.01673
R112 VTAIL.n14 VTAIL.t7 4.01673
R113 VTAIL.n14 VTAIL.t5 4.01673
R114 VTAIL.n12 VTAIL.t4 4.01673
R115 VTAIL.n12 VTAIL.t3 4.01673
R116 VTAIL.n9 VTAIL.t14 4.01673
R117 VTAIL.n9 VTAIL.t12 4.01673
R118 VTAIL.n7 VTAIL.t10 4.01673
R119 VTAIL.n7 VTAIL.t15 4.01673
R120 VTAIL.n10 VTAIL.n8 1.36257
R121 VTAIL.n11 VTAIL.n10 1.36257
R122 VTAIL.n15 VTAIL.n13 1.36257
R123 VTAIL.n16 VTAIL.n15 1.36257
R124 VTAIL.n6 VTAIL.n4 1.36257
R125 VTAIL.n4 VTAIL.n2 1.36257
R126 VTAIL.n19 VTAIL.n17 1.36257
R127 VTAIL.n13 VTAIL.n11 1.15136
R128 VTAIL.n2 VTAIL.n1 1.15136
R129 VTAIL VTAIL.n1 1.08024
R130 VTAIL VTAIL.n19 0.282828
R131 B.n556 B.n555 585
R132 B.n557 B.n556 585
R133 B.n197 B.n94 585
R134 B.n196 B.n195 585
R135 B.n194 B.n193 585
R136 B.n192 B.n191 585
R137 B.n190 B.n189 585
R138 B.n188 B.n187 585
R139 B.n186 B.n185 585
R140 B.n184 B.n183 585
R141 B.n182 B.n181 585
R142 B.n180 B.n179 585
R143 B.n178 B.n177 585
R144 B.n176 B.n175 585
R145 B.n174 B.n173 585
R146 B.n172 B.n171 585
R147 B.n170 B.n169 585
R148 B.n168 B.n167 585
R149 B.n166 B.n165 585
R150 B.n164 B.n163 585
R151 B.n162 B.n161 585
R152 B.n160 B.n159 585
R153 B.n158 B.n157 585
R154 B.n156 B.n155 585
R155 B.n154 B.n153 585
R156 B.n152 B.n151 585
R157 B.n150 B.n149 585
R158 B.n148 B.n147 585
R159 B.n146 B.n145 585
R160 B.n144 B.n143 585
R161 B.n142 B.n141 585
R162 B.n139 B.n138 585
R163 B.n137 B.n136 585
R164 B.n135 B.n134 585
R165 B.n133 B.n132 585
R166 B.n131 B.n130 585
R167 B.n129 B.n128 585
R168 B.n127 B.n126 585
R169 B.n125 B.n124 585
R170 B.n123 B.n122 585
R171 B.n121 B.n120 585
R172 B.n119 B.n118 585
R173 B.n117 B.n116 585
R174 B.n115 B.n114 585
R175 B.n113 B.n112 585
R176 B.n111 B.n110 585
R177 B.n109 B.n108 585
R178 B.n107 B.n106 585
R179 B.n105 B.n104 585
R180 B.n103 B.n102 585
R181 B.n101 B.n100 585
R182 B.n67 B.n66 585
R183 B.n554 B.n68 585
R184 B.n558 B.n68 585
R185 B.n553 B.n552 585
R186 B.n552 B.n64 585
R187 B.n551 B.n63 585
R188 B.n564 B.n63 585
R189 B.n550 B.n62 585
R190 B.n565 B.n62 585
R191 B.n549 B.n61 585
R192 B.n566 B.n61 585
R193 B.n548 B.n547 585
R194 B.n547 B.n60 585
R195 B.n546 B.n56 585
R196 B.n572 B.n56 585
R197 B.n545 B.n55 585
R198 B.n573 B.n55 585
R199 B.n544 B.n54 585
R200 B.n574 B.n54 585
R201 B.n543 B.n542 585
R202 B.n542 B.n50 585
R203 B.n541 B.n49 585
R204 B.n580 B.n49 585
R205 B.n540 B.n48 585
R206 B.n581 B.n48 585
R207 B.n539 B.n47 585
R208 B.n582 B.n47 585
R209 B.n538 B.n537 585
R210 B.n537 B.n46 585
R211 B.n536 B.n42 585
R212 B.n588 B.n42 585
R213 B.n535 B.n41 585
R214 B.n589 B.n41 585
R215 B.n534 B.n40 585
R216 B.n590 B.n40 585
R217 B.n533 B.n532 585
R218 B.n532 B.n36 585
R219 B.n531 B.n35 585
R220 B.n596 B.n35 585
R221 B.n530 B.n34 585
R222 B.n597 B.n34 585
R223 B.n529 B.n33 585
R224 B.n598 B.n33 585
R225 B.n528 B.n527 585
R226 B.n527 B.n29 585
R227 B.n526 B.n28 585
R228 B.n604 B.n28 585
R229 B.n525 B.n27 585
R230 B.n605 B.n27 585
R231 B.n524 B.n26 585
R232 B.n606 B.n26 585
R233 B.n523 B.n522 585
R234 B.n522 B.n22 585
R235 B.n521 B.n21 585
R236 B.n612 B.n21 585
R237 B.n520 B.n20 585
R238 B.n613 B.n20 585
R239 B.n519 B.n19 585
R240 B.n614 B.n19 585
R241 B.n518 B.n517 585
R242 B.n517 B.n15 585
R243 B.n516 B.n14 585
R244 B.n620 B.n14 585
R245 B.n515 B.n13 585
R246 B.n621 B.n13 585
R247 B.n514 B.n12 585
R248 B.n622 B.n12 585
R249 B.n513 B.n512 585
R250 B.n512 B.n8 585
R251 B.n511 B.n7 585
R252 B.n628 B.n7 585
R253 B.n510 B.n6 585
R254 B.n629 B.n6 585
R255 B.n509 B.n5 585
R256 B.n630 B.n5 585
R257 B.n508 B.n507 585
R258 B.n507 B.n4 585
R259 B.n506 B.n198 585
R260 B.n506 B.n505 585
R261 B.n496 B.n199 585
R262 B.n200 B.n199 585
R263 B.n498 B.n497 585
R264 B.n499 B.n498 585
R265 B.n495 B.n205 585
R266 B.n205 B.n204 585
R267 B.n494 B.n493 585
R268 B.n493 B.n492 585
R269 B.n207 B.n206 585
R270 B.n208 B.n207 585
R271 B.n485 B.n484 585
R272 B.n486 B.n485 585
R273 B.n483 B.n212 585
R274 B.n216 B.n212 585
R275 B.n482 B.n481 585
R276 B.n481 B.n480 585
R277 B.n214 B.n213 585
R278 B.n215 B.n214 585
R279 B.n473 B.n472 585
R280 B.n474 B.n473 585
R281 B.n471 B.n221 585
R282 B.n221 B.n220 585
R283 B.n470 B.n469 585
R284 B.n469 B.n468 585
R285 B.n223 B.n222 585
R286 B.n224 B.n223 585
R287 B.n461 B.n460 585
R288 B.n462 B.n461 585
R289 B.n459 B.n229 585
R290 B.n229 B.n228 585
R291 B.n458 B.n457 585
R292 B.n457 B.n456 585
R293 B.n231 B.n230 585
R294 B.n232 B.n231 585
R295 B.n449 B.n448 585
R296 B.n450 B.n449 585
R297 B.n447 B.n237 585
R298 B.n237 B.n236 585
R299 B.n446 B.n445 585
R300 B.n445 B.n444 585
R301 B.n239 B.n238 585
R302 B.n437 B.n239 585
R303 B.n436 B.n435 585
R304 B.n438 B.n436 585
R305 B.n434 B.n244 585
R306 B.n244 B.n243 585
R307 B.n433 B.n432 585
R308 B.n432 B.n431 585
R309 B.n246 B.n245 585
R310 B.n247 B.n246 585
R311 B.n424 B.n423 585
R312 B.n425 B.n424 585
R313 B.n422 B.n252 585
R314 B.n252 B.n251 585
R315 B.n421 B.n420 585
R316 B.n420 B.n419 585
R317 B.n254 B.n253 585
R318 B.n412 B.n254 585
R319 B.n411 B.n410 585
R320 B.n413 B.n411 585
R321 B.n409 B.n259 585
R322 B.n259 B.n258 585
R323 B.n408 B.n407 585
R324 B.n407 B.n406 585
R325 B.n261 B.n260 585
R326 B.n262 B.n261 585
R327 B.n399 B.n398 585
R328 B.n400 B.n399 585
R329 B.n265 B.n264 585
R330 B.n299 B.n298 585
R331 B.n300 B.n296 585
R332 B.n296 B.n266 585
R333 B.n302 B.n301 585
R334 B.n304 B.n295 585
R335 B.n307 B.n306 585
R336 B.n308 B.n294 585
R337 B.n310 B.n309 585
R338 B.n312 B.n293 585
R339 B.n315 B.n314 585
R340 B.n316 B.n292 585
R341 B.n318 B.n317 585
R342 B.n320 B.n291 585
R343 B.n323 B.n322 585
R344 B.n324 B.n290 585
R345 B.n326 B.n325 585
R346 B.n328 B.n289 585
R347 B.n331 B.n330 585
R348 B.n332 B.n288 585
R349 B.n334 B.n333 585
R350 B.n336 B.n287 585
R351 B.n339 B.n338 585
R352 B.n340 B.n283 585
R353 B.n342 B.n341 585
R354 B.n344 B.n282 585
R355 B.n347 B.n346 585
R356 B.n348 B.n281 585
R357 B.n350 B.n349 585
R358 B.n352 B.n280 585
R359 B.n355 B.n354 585
R360 B.n357 B.n277 585
R361 B.n359 B.n358 585
R362 B.n361 B.n276 585
R363 B.n364 B.n363 585
R364 B.n365 B.n275 585
R365 B.n367 B.n366 585
R366 B.n369 B.n274 585
R367 B.n372 B.n371 585
R368 B.n373 B.n273 585
R369 B.n375 B.n374 585
R370 B.n377 B.n272 585
R371 B.n380 B.n379 585
R372 B.n381 B.n271 585
R373 B.n383 B.n382 585
R374 B.n385 B.n270 585
R375 B.n388 B.n387 585
R376 B.n389 B.n269 585
R377 B.n391 B.n390 585
R378 B.n393 B.n268 585
R379 B.n396 B.n395 585
R380 B.n397 B.n267 585
R381 B.n402 B.n401 585
R382 B.n401 B.n400 585
R383 B.n403 B.n263 585
R384 B.n263 B.n262 585
R385 B.n405 B.n404 585
R386 B.n406 B.n405 585
R387 B.n257 B.n256 585
R388 B.n258 B.n257 585
R389 B.n415 B.n414 585
R390 B.n414 B.n413 585
R391 B.n416 B.n255 585
R392 B.n412 B.n255 585
R393 B.n418 B.n417 585
R394 B.n419 B.n418 585
R395 B.n250 B.n249 585
R396 B.n251 B.n250 585
R397 B.n427 B.n426 585
R398 B.n426 B.n425 585
R399 B.n428 B.n248 585
R400 B.n248 B.n247 585
R401 B.n430 B.n429 585
R402 B.n431 B.n430 585
R403 B.n242 B.n241 585
R404 B.n243 B.n242 585
R405 B.n440 B.n439 585
R406 B.n439 B.n438 585
R407 B.n441 B.n240 585
R408 B.n437 B.n240 585
R409 B.n443 B.n442 585
R410 B.n444 B.n443 585
R411 B.n235 B.n234 585
R412 B.n236 B.n235 585
R413 B.n452 B.n451 585
R414 B.n451 B.n450 585
R415 B.n453 B.n233 585
R416 B.n233 B.n232 585
R417 B.n455 B.n454 585
R418 B.n456 B.n455 585
R419 B.n227 B.n226 585
R420 B.n228 B.n227 585
R421 B.n464 B.n463 585
R422 B.n463 B.n462 585
R423 B.n465 B.n225 585
R424 B.n225 B.n224 585
R425 B.n467 B.n466 585
R426 B.n468 B.n467 585
R427 B.n219 B.n218 585
R428 B.n220 B.n219 585
R429 B.n476 B.n475 585
R430 B.n475 B.n474 585
R431 B.n477 B.n217 585
R432 B.n217 B.n215 585
R433 B.n479 B.n478 585
R434 B.n480 B.n479 585
R435 B.n211 B.n210 585
R436 B.n216 B.n211 585
R437 B.n488 B.n487 585
R438 B.n487 B.n486 585
R439 B.n489 B.n209 585
R440 B.n209 B.n208 585
R441 B.n491 B.n490 585
R442 B.n492 B.n491 585
R443 B.n203 B.n202 585
R444 B.n204 B.n203 585
R445 B.n501 B.n500 585
R446 B.n500 B.n499 585
R447 B.n502 B.n201 585
R448 B.n201 B.n200 585
R449 B.n504 B.n503 585
R450 B.n505 B.n504 585
R451 B.n2 B.n0 585
R452 B.n4 B.n2 585
R453 B.n3 B.n1 585
R454 B.n629 B.n3 585
R455 B.n627 B.n626 585
R456 B.n628 B.n627 585
R457 B.n625 B.n9 585
R458 B.n9 B.n8 585
R459 B.n624 B.n623 585
R460 B.n623 B.n622 585
R461 B.n11 B.n10 585
R462 B.n621 B.n11 585
R463 B.n619 B.n618 585
R464 B.n620 B.n619 585
R465 B.n617 B.n16 585
R466 B.n16 B.n15 585
R467 B.n616 B.n615 585
R468 B.n615 B.n614 585
R469 B.n18 B.n17 585
R470 B.n613 B.n18 585
R471 B.n611 B.n610 585
R472 B.n612 B.n611 585
R473 B.n609 B.n23 585
R474 B.n23 B.n22 585
R475 B.n608 B.n607 585
R476 B.n607 B.n606 585
R477 B.n25 B.n24 585
R478 B.n605 B.n25 585
R479 B.n603 B.n602 585
R480 B.n604 B.n603 585
R481 B.n601 B.n30 585
R482 B.n30 B.n29 585
R483 B.n600 B.n599 585
R484 B.n599 B.n598 585
R485 B.n32 B.n31 585
R486 B.n597 B.n32 585
R487 B.n595 B.n594 585
R488 B.n596 B.n595 585
R489 B.n593 B.n37 585
R490 B.n37 B.n36 585
R491 B.n592 B.n591 585
R492 B.n591 B.n590 585
R493 B.n39 B.n38 585
R494 B.n589 B.n39 585
R495 B.n587 B.n586 585
R496 B.n588 B.n587 585
R497 B.n585 B.n43 585
R498 B.n46 B.n43 585
R499 B.n584 B.n583 585
R500 B.n583 B.n582 585
R501 B.n45 B.n44 585
R502 B.n581 B.n45 585
R503 B.n579 B.n578 585
R504 B.n580 B.n579 585
R505 B.n577 B.n51 585
R506 B.n51 B.n50 585
R507 B.n576 B.n575 585
R508 B.n575 B.n574 585
R509 B.n53 B.n52 585
R510 B.n573 B.n53 585
R511 B.n571 B.n570 585
R512 B.n572 B.n571 585
R513 B.n569 B.n57 585
R514 B.n60 B.n57 585
R515 B.n568 B.n567 585
R516 B.n567 B.n566 585
R517 B.n59 B.n58 585
R518 B.n565 B.n59 585
R519 B.n563 B.n562 585
R520 B.n564 B.n563 585
R521 B.n561 B.n65 585
R522 B.n65 B.n64 585
R523 B.n560 B.n559 585
R524 B.n559 B.n558 585
R525 B.n632 B.n631 585
R526 B.n631 B.n630 585
R527 B.n401 B.n265 516.524
R528 B.n559 B.n67 516.524
R529 B.n399 B.n267 516.524
R530 B.n556 B.n68 516.524
R531 B.n278 B.t14 299.421
R532 B.n284 B.t10 299.421
R533 B.n98 B.t17 299.421
R534 B.n95 B.t21 299.421
R535 B.n557 B.n93 256.663
R536 B.n557 B.n92 256.663
R537 B.n557 B.n91 256.663
R538 B.n557 B.n90 256.663
R539 B.n557 B.n89 256.663
R540 B.n557 B.n88 256.663
R541 B.n557 B.n87 256.663
R542 B.n557 B.n86 256.663
R543 B.n557 B.n85 256.663
R544 B.n557 B.n84 256.663
R545 B.n557 B.n83 256.663
R546 B.n557 B.n82 256.663
R547 B.n557 B.n81 256.663
R548 B.n557 B.n80 256.663
R549 B.n557 B.n79 256.663
R550 B.n557 B.n78 256.663
R551 B.n557 B.n77 256.663
R552 B.n557 B.n76 256.663
R553 B.n557 B.n75 256.663
R554 B.n557 B.n74 256.663
R555 B.n557 B.n73 256.663
R556 B.n557 B.n72 256.663
R557 B.n557 B.n71 256.663
R558 B.n557 B.n70 256.663
R559 B.n557 B.n69 256.663
R560 B.n297 B.n266 256.663
R561 B.n303 B.n266 256.663
R562 B.n305 B.n266 256.663
R563 B.n311 B.n266 256.663
R564 B.n313 B.n266 256.663
R565 B.n319 B.n266 256.663
R566 B.n321 B.n266 256.663
R567 B.n327 B.n266 256.663
R568 B.n329 B.n266 256.663
R569 B.n335 B.n266 256.663
R570 B.n337 B.n266 256.663
R571 B.n343 B.n266 256.663
R572 B.n345 B.n266 256.663
R573 B.n351 B.n266 256.663
R574 B.n353 B.n266 256.663
R575 B.n360 B.n266 256.663
R576 B.n362 B.n266 256.663
R577 B.n368 B.n266 256.663
R578 B.n370 B.n266 256.663
R579 B.n376 B.n266 256.663
R580 B.n378 B.n266 256.663
R581 B.n384 B.n266 256.663
R582 B.n386 B.n266 256.663
R583 B.n392 B.n266 256.663
R584 B.n394 B.n266 256.663
R585 B.n401 B.n263 163.367
R586 B.n405 B.n263 163.367
R587 B.n405 B.n257 163.367
R588 B.n414 B.n257 163.367
R589 B.n414 B.n255 163.367
R590 B.n418 B.n255 163.367
R591 B.n418 B.n250 163.367
R592 B.n426 B.n250 163.367
R593 B.n426 B.n248 163.367
R594 B.n430 B.n248 163.367
R595 B.n430 B.n242 163.367
R596 B.n439 B.n242 163.367
R597 B.n439 B.n240 163.367
R598 B.n443 B.n240 163.367
R599 B.n443 B.n235 163.367
R600 B.n451 B.n235 163.367
R601 B.n451 B.n233 163.367
R602 B.n455 B.n233 163.367
R603 B.n455 B.n227 163.367
R604 B.n463 B.n227 163.367
R605 B.n463 B.n225 163.367
R606 B.n467 B.n225 163.367
R607 B.n467 B.n219 163.367
R608 B.n475 B.n219 163.367
R609 B.n475 B.n217 163.367
R610 B.n479 B.n217 163.367
R611 B.n479 B.n211 163.367
R612 B.n487 B.n211 163.367
R613 B.n487 B.n209 163.367
R614 B.n491 B.n209 163.367
R615 B.n491 B.n203 163.367
R616 B.n500 B.n203 163.367
R617 B.n500 B.n201 163.367
R618 B.n504 B.n201 163.367
R619 B.n504 B.n2 163.367
R620 B.n631 B.n2 163.367
R621 B.n631 B.n3 163.367
R622 B.n627 B.n3 163.367
R623 B.n627 B.n9 163.367
R624 B.n623 B.n9 163.367
R625 B.n623 B.n11 163.367
R626 B.n619 B.n11 163.367
R627 B.n619 B.n16 163.367
R628 B.n615 B.n16 163.367
R629 B.n615 B.n18 163.367
R630 B.n611 B.n18 163.367
R631 B.n611 B.n23 163.367
R632 B.n607 B.n23 163.367
R633 B.n607 B.n25 163.367
R634 B.n603 B.n25 163.367
R635 B.n603 B.n30 163.367
R636 B.n599 B.n30 163.367
R637 B.n599 B.n32 163.367
R638 B.n595 B.n32 163.367
R639 B.n595 B.n37 163.367
R640 B.n591 B.n37 163.367
R641 B.n591 B.n39 163.367
R642 B.n587 B.n39 163.367
R643 B.n587 B.n43 163.367
R644 B.n583 B.n43 163.367
R645 B.n583 B.n45 163.367
R646 B.n579 B.n45 163.367
R647 B.n579 B.n51 163.367
R648 B.n575 B.n51 163.367
R649 B.n575 B.n53 163.367
R650 B.n571 B.n53 163.367
R651 B.n571 B.n57 163.367
R652 B.n567 B.n57 163.367
R653 B.n567 B.n59 163.367
R654 B.n563 B.n59 163.367
R655 B.n563 B.n65 163.367
R656 B.n559 B.n65 163.367
R657 B.n298 B.n296 163.367
R658 B.n302 B.n296 163.367
R659 B.n306 B.n304 163.367
R660 B.n310 B.n294 163.367
R661 B.n314 B.n312 163.367
R662 B.n318 B.n292 163.367
R663 B.n322 B.n320 163.367
R664 B.n326 B.n290 163.367
R665 B.n330 B.n328 163.367
R666 B.n334 B.n288 163.367
R667 B.n338 B.n336 163.367
R668 B.n342 B.n283 163.367
R669 B.n346 B.n344 163.367
R670 B.n350 B.n281 163.367
R671 B.n354 B.n352 163.367
R672 B.n359 B.n277 163.367
R673 B.n363 B.n361 163.367
R674 B.n367 B.n275 163.367
R675 B.n371 B.n369 163.367
R676 B.n375 B.n273 163.367
R677 B.n379 B.n377 163.367
R678 B.n383 B.n271 163.367
R679 B.n387 B.n385 163.367
R680 B.n391 B.n269 163.367
R681 B.n395 B.n393 163.367
R682 B.n399 B.n261 163.367
R683 B.n407 B.n261 163.367
R684 B.n407 B.n259 163.367
R685 B.n411 B.n259 163.367
R686 B.n411 B.n254 163.367
R687 B.n420 B.n254 163.367
R688 B.n420 B.n252 163.367
R689 B.n424 B.n252 163.367
R690 B.n424 B.n246 163.367
R691 B.n432 B.n246 163.367
R692 B.n432 B.n244 163.367
R693 B.n436 B.n244 163.367
R694 B.n436 B.n239 163.367
R695 B.n445 B.n239 163.367
R696 B.n445 B.n237 163.367
R697 B.n449 B.n237 163.367
R698 B.n449 B.n231 163.367
R699 B.n457 B.n231 163.367
R700 B.n457 B.n229 163.367
R701 B.n461 B.n229 163.367
R702 B.n461 B.n223 163.367
R703 B.n469 B.n223 163.367
R704 B.n469 B.n221 163.367
R705 B.n473 B.n221 163.367
R706 B.n473 B.n214 163.367
R707 B.n481 B.n214 163.367
R708 B.n481 B.n212 163.367
R709 B.n485 B.n212 163.367
R710 B.n485 B.n207 163.367
R711 B.n493 B.n207 163.367
R712 B.n493 B.n205 163.367
R713 B.n498 B.n205 163.367
R714 B.n498 B.n199 163.367
R715 B.n506 B.n199 163.367
R716 B.n507 B.n506 163.367
R717 B.n507 B.n5 163.367
R718 B.n6 B.n5 163.367
R719 B.n7 B.n6 163.367
R720 B.n512 B.n7 163.367
R721 B.n512 B.n12 163.367
R722 B.n13 B.n12 163.367
R723 B.n14 B.n13 163.367
R724 B.n517 B.n14 163.367
R725 B.n517 B.n19 163.367
R726 B.n20 B.n19 163.367
R727 B.n21 B.n20 163.367
R728 B.n522 B.n21 163.367
R729 B.n522 B.n26 163.367
R730 B.n27 B.n26 163.367
R731 B.n28 B.n27 163.367
R732 B.n527 B.n28 163.367
R733 B.n527 B.n33 163.367
R734 B.n34 B.n33 163.367
R735 B.n35 B.n34 163.367
R736 B.n532 B.n35 163.367
R737 B.n532 B.n40 163.367
R738 B.n41 B.n40 163.367
R739 B.n42 B.n41 163.367
R740 B.n537 B.n42 163.367
R741 B.n537 B.n47 163.367
R742 B.n48 B.n47 163.367
R743 B.n49 B.n48 163.367
R744 B.n542 B.n49 163.367
R745 B.n542 B.n54 163.367
R746 B.n55 B.n54 163.367
R747 B.n56 B.n55 163.367
R748 B.n547 B.n56 163.367
R749 B.n547 B.n61 163.367
R750 B.n62 B.n61 163.367
R751 B.n63 B.n62 163.367
R752 B.n552 B.n63 163.367
R753 B.n552 B.n68 163.367
R754 B.n102 B.n101 163.367
R755 B.n106 B.n105 163.367
R756 B.n110 B.n109 163.367
R757 B.n114 B.n113 163.367
R758 B.n118 B.n117 163.367
R759 B.n122 B.n121 163.367
R760 B.n126 B.n125 163.367
R761 B.n130 B.n129 163.367
R762 B.n134 B.n133 163.367
R763 B.n138 B.n137 163.367
R764 B.n143 B.n142 163.367
R765 B.n147 B.n146 163.367
R766 B.n151 B.n150 163.367
R767 B.n155 B.n154 163.367
R768 B.n159 B.n158 163.367
R769 B.n163 B.n162 163.367
R770 B.n167 B.n166 163.367
R771 B.n171 B.n170 163.367
R772 B.n175 B.n174 163.367
R773 B.n179 B.n178 163.367
R774 B.n183 B.n182 163.367
R775 B.n187 B.n186 163.367
R776 B.n191 B.n190 163.367
R777 B.n195 B.n194 163.367
R778 B.n556 B.n94 163.367
R779 B.n400 B.n266 132.583
R780 B.n558 B.n557 132.583
R781 B.n278 B.t16 104.183
R782 B.n95 B.t22 104.183
R783 B.n284 B.t13 104.178
R784 B.n98 B.t19 104.178
R785 B.n279 B.t15 73.5411
R786 B.n96 B.t23 73.5411
R787 B.n285 B.t12 73.5363
R788 B.n99 B.t20 73.5363
R789 B.n400 B.n262 73.2979
R790 B.n406 B.n262 73.2979
R791 B.n406 B.n258 73.2979
R792 B.n413 B.n258 73.2979
R793 B.n413 B.n412 73.2979
R794 B.n419 B.n251 73.2979
R795 B.n425 B.n251 73.2979
R796 B.n425 B.n247 73.2979
R797 B.n431 B.n247 73.2979
R798 B.n431 B.n243 73.2979
R799 B.n438 B.n243 73.2979
R800 B.n438 B.n437 73.2979
R801 B.n444 B.n236 73.2979
R802 B.n450 B.n236 73.2979
R803 B.n450 B.n232 73.2979
R804 B.n456 B.n232 73.2979
R805 B.n462 B.n228 73.2979
R806 B.n462 B.n224 73.2979
R807 B.n468 B.n224 73.2979
R808 B.n474 B.n220 73.2979
R809 B.n474 B.n215 73.2979
R810 B.n480 B.n215 73.2979
R811 B.n480 B.n216 73.2979
R812 B.n486 B.n208 73.2979
R813 B.n492 B.n208 73.2979
R814 B.n492 B.n204 73.2979
R815 B.n499 B.n204 73.2979
R816 B.n505 B.n200 73.2979
R817 B.n505 B.n4 73.2979
R818 B.n630 B.n4 73.2979
R819 B.n630 B.n629 73.2979
R820 B.n629 B.n628 73.2979
R821 B.n628 B.n8 73.2979
R822 B.n622 B.n621 73.2979
R823 B.n621 B.n620 73.2979
R824 B.n620 B.n15 73.2979
R825 B.n614 B.n15 73.2979
R826 B.n613 B.n612 73.2979
R827 B.n612 B.n22 73.2979
R828 B.n606 B.n22 73.2979
R829 B.n606 B.n605 73.2979
R830 B.n604 B.n29 73.2979
R831 B.n598 B.n29 73.2979
R832 B.n598 B.n597 73.2979
R833 B.n596 B.n36 73.2979
R834 B.n590 B.n36 73.2979
R835 B.n590 B.n589 73.2979
R836 B.n589 B.n588 73.2979
R837 B.n582 B.n46 73.2979
R838 B.n582 B.n581 73.2979
R839 B.n581 B.n580 73.2979
R840 B.n580 B.n50 73.2979
R841 B.n574 B.n50 73.2979
R842 B.n574 B.n573 73.2979
R843 B.n573 B.n572 73.2979
R844 B.n566 B.n60 73.2979
R845 B.n566 B.n565 73.2979
R846 B.n565 B.n564 73.2979
R847 B.n564 B.n64 73.2979
R848 B.n558 B.n64 73.2979
R849 B.n297 B.n265 71.676
R850 B.n303 B.n302 71.676
R851 B.n306 B.n305 71.676
R852 B.n311 B.n310 71.676
R853 B.n314 B.n313 71.676
R854 B.n319 B.n318 71.676
R855 B.n322 B.n321 71.676
R856 B.n327 B.n326 71.676
R857 B.n330 B.n329 71.676
R858 B.n335 B.n334 71.676
R859 B.n338 B.n337 71.676
R860 B.n343 B.n342 71.676
R861 B.n346 B.n345 71.676
R862 B.n351 B.n350 71.676
R863 B.n354 B.n353 71.676
R864 B.n360 B.n359 71.676
R865 B.n363 B.n362 71.676
R866 B.n368 B.n367 71.676
R867 B.n371 B.n370 71.676
R868 B.n376 B.n375 71.676
R869 B.n379 B.n378 71.676
R870 B.n384 B.n383 71.676
R871 B.n387 B.n386 71.676
R872 B.n392 B.n391 71.676
R873 B.n395 B.n394 71.676
R874 B.n69 B.n67 71.676
R875 B.n102 B.n70 71.676
R876 B.n106 B.n71 71.676
R877 B.n110 B.n72 71.676
R878 B.n114 B.n73 71.676
R879 B.n118 B.n74 71.676
R880 B.n122 B.n75 71.676
R881 B.n126 B.n76 71.676
R882 B.n130 B.n77 71.676
R883 B.n134 B.n78 71.676
R884 B.n138 B.n79 71.676
R885 B.n143 B.n80 71.676
R886 B.n147 B.n81 71.676
R887 B.n151 B.n82 71.676
R888 B.n155 B.n83 71.676
R889 B.n159 B.n84 71.676
R890 B.n163 B.n85 71.676
R891 B.n167 B.n86 71.676
R892 B.n171 B.n87 71.676
R893 B.n175 B.n88 71.676
R894 B.n179 B.n89 71.676
R895 B.n183 B.n90 71.676
R896 B.n187 B.n91 71.676
R897 B.n191 B.n92 71.676
R898 B.n195 B.n93 71.676
R899 B.n94 B.n93 71.676
R900 B.n194 B.n92 71.676
R901 B.n190 B.n91 71.676
R902 B.n186 B.n90 71.676
R903 B.n182 B.n89 71.676
R904 B.n178 B.n88 71.676
R905 B.n174 B.n87 71.676
R906 B.n170 B.n86 71.676
R907 B.n166 B.n85 71.676
R908 B.n162 B.n84 71.676
R909 B.n158 B.n83 71.676
R910 B.n154 B.n82 71.676
R911 B.n150 B.n81 71.676
R912 B.n146 B.n80 71.676
R913 B.n142 B.n79 71.676
R914 B.n137 B.n78 71.676
R915 B.n133 B.n77 71.676
R916 B.n129 B.n76 71.676
R917 B.n125 B.n75 71.676
R918 B.n121 B.n74 71.676
R919 B.n117 B.n73 71.676
R920 B.n113 B.n72 71.676
R921 B.n109 B.n71 71.676
R922 B.n105 B.n70 71.676
R923 B.n101 B.n69 71.676
R924 B.n298 B.n297 71.676
R925 B.n304 B.n303 71.676
R926 B.n305 B.n294 71.676
R927 B.n312 B.n311 71.676
R928 B.n313 B.n292 71.676
R929 B.n320 B.n319 71.676
R930 B.n321 B.n290 71.676
R931 B.n328 B.n327 71.676
R932 B.n329 B.n288 71.676
R933 B.n336 B.n335 71.676
R934 B.n337 B.n283 71.676
R935 B.n344 B.n343 71.676
R936 B.n345 B.n281 71.676
R937 B.n352 B.n351 71.676
R938 B.n353 B.n277 71.676
R939 B.n361 B.n360 71.676
R940 B.n362 B.n275 71.676
R941 B.n369 B.n368 71.676
R942 B.n370 B.n273 71.676
R943 B.n377 B.n376 71.676
R944 B.n378 B.n271 71.676
R945 B.n385 B.n384 71.676
R946 B.n386 B.n269 71.676
R947 B.n393 B.n392 71.676
R948 B.n394 B.n267 71.676
R949 B.t0 B.n200 67.9084
R950 B.t4 B.n8 67.9084
R951 B.t6 B.n228 63.5968
R952 B.n597 B.t5 63.5968
R953 B.n356 B.n279 59.5399
R954 B.n286 B.n285 59.5399
R955 B.n140 B.n99 59.5399
R956 B.n97 B.n96 59.5399
R957 B.n468 B.t2 57.1294
R958 B.t7 B.n604 57.1294
R959 B.n412 B.t11 46.3503
R960 B.n60 B.t18 46.3503
R961 B.n486 B.t1 42.0387
R962 B.n614 B.t3 42.0387
R963 B.n444 B.t8 37.7271
R964 B.n588 B.t9 37.7271
R965 B.n437 B.t8 35.5713
R966 B.n46 B.t9 35.5713
R967 B.n560 B.n66 33.5615
R968 B.n555 B.n554 33.5615
R969 B.n398 B.n397 33.5615
R970 B.n402 B.n264 33.5615
R971 B.n216 B.t1 31.2597
R972 B.t3 B.n613 31.2597
R973 B.n279 B.n278 30.6429
R974 B.n285 B.n284 30.6429
R975 B.n99 B.n98 30.6429
R976 B.n96 B.n95 30.6429
R977 B.n419 B.t11 26.9481
R978 B.n572 B.t18 26.9481
R979 B B.n632 18.0485
R980 B.t2 B.n220 16.169
R981 B.n605 B.t7 16.169
R982 B.n100 B.n66 10.6151
R983 B.n103 B.n100 10.6151
R984 B.n104 B.n103 10.6151
R985 B.n107 B.n104 10.6151
R986 B.n108 B.n107 10.6151
R987 B.n111 B.n108 10.6151
R988 B.n112 B.n111 10.6151
R989 B.n115 B.n112 10.6151
R990 B.n116 B.n115 10.6151
R991 B.n119 B.n116 10.6151
R992 B.n120 B.n119 10.6151
R993 B.n123 B.n120 10.6151
R994 B.n124 B.n123 10.6151
R995 B.n127 B.n124 10.6151
R996 B.n128 B.n127 10.6151
R997 B.n131 B.n128 10.6151
R998 B.n132 B.n131 10.6151
R999 B.n135 B.n132 10.6151
R1000 B.n136 B.n135 10.6151
R1001 B.n139 B.n136 10.6151
R1002 B.n144 B.n141 10.6151
R1003 B.n145 B.n144 10.6151
R1004 B.n148 B.n145 10.6151
R1005 B.n149 B.n148 10.6151
R1006 B.n152 B.n149 10.6151
R1007 B.n153 B.n152 10.6151
R1008 B.n156 B.n153 10.6151
R1009 B.n157 B.n156 10.6151
R1010 B.n161 B.n160 10.6151
R1011 B.n164 B.n161 10.6151
R1012 B.n165 B.n164 10.6151
R1013 B.n168 B.n165 10.6151
R1014 B.n169 B.n168 10.6151
R1015 B.n172 B.n169 10.6151
R1016 B.n173 B.n172 10.6151
R1017 B.n176 B.n173 10.6151
R1018 B.n177 B.n176 10.6151
R1019 B.n180 B.n177 10.6151
R1020 B.n181 B.n180 10.6151
R1021 B.n184 B.n181 10.6151
R1022 B.n185 B.n184 10.6151
R1023 B.n188 B.n185 10.6151
R1024 B.n189 B.n188 10.6151
R1025 B.n192 B.n189 10.6151
R1026 B.n193 B.n192 10.6151
R1027 B.n196 B.n193 10.6151
R1028 B.n197 B.n196 10.6151
R1029 B.n555 B.n197 10.6151
R1030 B.n398 B.n260 10.6151
R1031 B.n408 B.n260 10.6151
R1032 B.n409 B.n408 10.6151
R1033 B.n410 B.n409 10.6151
R1034 B.n410 B.n253 10.6151
R1035 B.n421 B.n253 10.6151
R1036 B.n422 B.n421 10.6151
R1037 B.n423 B.n422 10.6151
R1038 B.n423 B.n245 10.6151
R1039 B.n433 B.n245 10.6151
R1040 B.n434 B.n433 10.6151
R1041 B.n435 B.n434 10.6151
R1042 B.n435 B.n238 10.6151
R1043 B.n446 B.n238 10.6151
R1044 B.n447 B.n446 10.6151
R1045 B.n448 B.n447 10.6151
R1046 B.n448 B.n230 10.6151
R1047 B.n458 B.n230 10.6151
R1048 B.n459 B.n458 10.6151
R1049 B.n460 B.n459 10.6151
R1050 B.n460 B.n222 10.6151
R1051 B.n470 B.n222 10.6151
R1052 B.n471 B.n470 10.6151
R1053 B.n472 B.n471 10.6151
R1054 B.n472 B.n213 10.6151
R1055 B.n482 B.n213 10.6151
R1056 B.n483 B.n482 10.6151
R1057 B.n484 B.n483 10.6151
R1058 B.n484 B.n206 10.6151
R1059 B.n494 B.n206 10.6151
R1060 B.n495 B.n494 10.6151
R1061 B.n497 B.n495 10.6151
R1062 B.n497 B.n496 10.6151
R1063 B.n496 B.n198 10.6151
R1064 B.n508 B.n198 10.6151
R1065 B.n509 B.n508 10.6151
R1066 B.n510 B.n509 10.6151
R1067 B.n511 B.n510 10.6151
R1068 B.n513 B.n511 10.6151
R1069 B.n514 B.n513 10.6151
R1070 B.n515 B.n514 10.6151
R1071 B.n516 B.n515 10.6151
R1072 B.n518 B.n516 10.6151
R1073 B.n519 B.n518 10.6151
R1074 B.n520 B.n519 10.6151
R1075 B.n521 B.n520 10.6151
R1076 B.n523 B.n521 10.6151
R1077 B.n524 B.n523 10.6151
R1078 B.n525 B.n524 10.6151
R1079 B.n526 B.n525 10.6151
R1080 B.n528 B.n526 10.6151
R1081 B.n529 B.n528 10.6151
R1082 B.n530 B.n529 10.6151
R1083 B.n531 B.n530 10.6151
R1084 B.n533 B.n531 10.6151
R1085 B.n534 B.n533 10.6151
R1086 B.n535 B.n534 10.6151
R1087 B.n536 B.n535 10.6151
R1088 B.n538 B.n536 10.6151
R1089 B.n539 B.n538 10.6151
R1090 B.n540 B.n539 10.6151
R1091 B.n541 B.n540 10.6151
R1092 B.n543 B.n541 10.6151
R1093 B.n544 B.n543 10.6151
R1094 B.n545 B.n544 10.6151
R1095 B.n546 B.n545 10.6151
R1096 B.n548 B.n546 10.6151
R1097 B.n549 B.n548 10.6151
R1098 B.n550 B.n549 10.6151
R1099 B.n551 B.n550 10.6151
R1100 B.n553 B.n551 10.6151
R1101 B.n554 B.n553 10.6151
R1102 B.n299 B.n264 10.6151
R1103 B.n300 B.n299 10.6151
R1104 B.n301 B.n300 10.6151
R1105 B.n301 B.n295 10.6151
R1106 B.n307 B.n295 10.6151
R1107 B.n308 B.n307 10.6151
R1108 B.n309 B.n308 10.6151
R1109 B.n309 B.n293 10.6151
R1110 B.n315 B.n293 10.6151
R1111 B.n316 B.n315 10.6151
R1112 B.n317 B.n316 10.6151
R1113 B.n317 B.n291 10.6151
R1114 B.n323 B.n291 10.6151
R1115 B.n324 B.n323 10.6151
R1116 B.n325 B.n324 10.6151
R1117 B.n325 B.n289 10.6151
R1118 B.n331 B.n289 10.6151
R1119 B.n332 B.n331 10.6151
R1120 B.n333 B.n332 10.6151
R1121 B.n333 B.n287 10.6151
R1122 B.n340 B.n339 10.6151
R1123 B.n341 B.n340 10.6151
R1124 B.n341 B.n282 10.6151
R1125 B.n347 B.n282 10.6151
R1126 B.n348 B.n347 10.6151
R1127 B.n349 B.n348 10.6151
R1128 B.n349 B.n280 10.6151
R1129 B.n355 B.n280 10.6151
R1130 B.n358 B.n357 10.6151
R1131 B.n358 B.n276 10.6151
R1132 B.n364 B.n276 10.6151
R1133 B.n365 B.n364 10.6151
R1134 B.n366 B.n365 10.6151
R1135 B.n366 B.n274 10.6151
R1136 B.n372 B.n274 10.6151
R1137 B.n373 B.n372 10.6151
R1138 B.n374 B.n373 10.6151
R1139 B.n374 B.n272 10.6151
R1140 B.n380 B.n272 10.6151
R1141 B.n381 B.n380 10.6151
R1142 B.n382 B.n381 10.6151
R1143 B.n382 B.n270 10.6151
R1144 B.n388 B.n270 10.6151
R1145 B.n389 B.n388 10.6151
R1146 B.n390 B.n389 10.6151
R1147 B.n390 B.n268 10.6151
R1148 B.n396 B.n268 10.6151
R1149 B.n397 B.n396 10.6151
R1150 B.n403 B.n402 10.6151
R1151 B.n404 B.n403 10.6151
R1152 B.n404 B.n256 10.6151
R1153 B.n415 B.n256 10.6151
R1154 B.n416 B.n415 10.6151
R1155 B.n417 B.n416 10.6151
R1156 B.n417 B.n249 10.6151
R1157 B.n427 B.n249 10.6151
R1158 B.n428 B.n427 10.6151
R1159 B.n429 B.n428 10.6151
R1160 B.n429 B.n241 10.6151
R1161 B.n440 B.n241 10.6151
R1162 B.n441 B.n440 10.6151
R1163 B.n442 B.n441 10.6151
R1164 B.n442 B.n234 10.6151
R1165 B.n452 B.n234 10.6151
R1166 B.n453 B.n452 10.6151
R1167 B.n454 B.n453 10.6151
R1168 B.n454 B.n226 10.6151
R1169 B.n464 B.n226 10.6151
R1170 B.n465 B.n464 10.6151
R1171 B.n466 B.n465 10.6151
R1172 B.n466 B.n218 10.6151
R1173 B.n476 B.n218 10.6151
R1174 B.n477 B.n476 10.6151
R1175 B.n478 B.n477 10.6151
R1176 B.n478 B.n210 10.6151
R1177 B.n488 B.n210 10.6151
R1178 B.n489 B.n488 10.6151
R1179 B.n490 B.n489 10.6151
R1180 B.n490 B.n202 10.6151
R1181 B.n501 B.n202 10.6151
R1182 B.n502 B.n501 10.6151
R1183 B.n503 B.n502 10.6151
R1184 B.n503 B.n0 10.6151
R1185 B.n626 B.n1 10.6151
R1186 B.n626 B.n625 10.6151
R1187 B.n625 B.n624 10.6151
R1188 B.n624 B.n10 10.6151
R1189 B.n618 B.n10 10.6151
R1190 B.n618 B.n617 10.6151
R1191 B.n617 B.n616 10.6151
R1192 B.n616 B.n17 10.6151
R1193 B.n610 B.n17 10.6151
R1194 B.n610 B.n609 10.6151
R1195 B.n609 B.n608 10.6151
R1196 B.n608 B.n24 10.6151
R1197 B.n602 B.n24 10.6151
R1198 B.n602 B.n601 10.6151
R1199 B.n601 B.n600 10.6151
R1200 B.n600 B.n31 10.6151
R1201 B.n594 B.n31 10.6151
R1202 B.n594 B.n593 10.6151
R1203 B.n593 B.n592 10.6151
R1204 B.n592 B.n38 10.6151
R1205 B.n586 B.n38 10.6151
R1206 B.n586 B.n585 10.6151
R1207 B.n585 B.n584 10.6151
R1208 B.n584 B.n44 10.6151
R1209 B.n578 B.n44 10.6151
R1210 B.n578 B.n577 10.6151
R1211 B.n577 B.n576 10.6151
R1212 B.n576 B.n52 10.6151
R1213 B.n570 B.n52 10.6151
R1214 B.n570 B.n569 10.6151
R1215 B.n569 B.n568 10.6151
R1216 B.n568 B.n58 10.6151
R1217 B.n562 B.n58 10.6151
R1218 B.n562 B.n561 10.6151
R1219 B.n561 B.n560 10.6151
R1220 B.n456 B.t6 9.70163
R1221 B.t5 B.n596 9.70163
R1222 B.n141 B.n140 6.5566
R1223 B.n157 B.n97 6.5566
R1224 B.n339 B.n286 6.5566
R1225 B.n356 B.n355 6.5566
R1226 B.n499 B.t0 5.39001
R1227 B.n622 B.t4 5.39001
R1228 B.n140 B.n139 4.05904
R1229 B.n160 B.n97 4.05904
R1230 B.n287 B.n286 4.05904
R1231 B.n357 B.n356 4.05904
R1232 B.n632 B.n0 2.81026
R1233 B.n632 B.n1 2.81026
R1234 VP.n15 VP.n14 161.3
R1235 VP.n16 VP.n11 161.3
R1236 VP.n18 VP.n17 161.3
R1237 VP.n20 VP.n19 161.3
R1238 VP.n21 VP.n9 161.3
R1239 VP.n23 VP.n22 161.3
R1240 VP.n25 VP.n24 161.3
R1241 VP.n26 VP.n7 161.3
R1242 VP.n46 VP.n0 161.3
R1243 VP.n45 VP.n44 161.3
R1244 VP.n43 VP.n42 161.3
R1245 VP.n41 VP.n2 161.3
R1246 VP.n40 VP.n39 161.3
R1247 VP.n38 VP.n37 161.3
R1248 VP.n36 VP.n4 161.3
R1249 VP.n35 VP.n34 161.3
R1250 VP.n33 VP.n32 161.3
R1251 VP.n31 VP.n6 161.3
R1252 VP.n13 VP.t7 147.857
R1253 VP.n30 VP.t4 126.671
R1254 VP.n47 VP.t0 126.671
R1255 VP.n27 VP.t2 126.671
R1256 VP.n5 VP.t3 95.0509
R1257 VP.n3 VP.t1 95.0509
R1258 VP.n1 VP.t8 95.0509
R1259 VP.n8 VP.t5 95.0509
R1260 VP.n10 VP.t6 95.0509
R1261 VP.n12 VP.t9 95.0509
R1262 VP.n28 VP.n27 80.6037
R1263 VP.n48 VP.n47 80.6037
R1264 VP.n30 VP.n29 80.6037
R1265 VP.n36 VP.n35 44.3785
R1266 VP.n42 VP.n41 44.3785
R1267 VP.n22 VP.n21 44.3785
R1268 VP.n16 VP.n15 44.3785
R1269 VP.n31 VP.n30 41.6278
R1270 VP.n47 VP.n46 41.6278
R1271 VP.n27 VP.n26 41.6278
R1272 VP.n13 VP.n12 40.893
R1273 VP.n29 VP.n28 40.6302
R1274 VP.n37 VP.n36 36.6083
R1275 VP.n41 VP.n40 36.6083
R1276 VP.n21 VP.n20 36.6083
R1277 VP.n17 VP.n16 36.6083
R1278 VP.n32 VP.n31 28.8382
R1279 VP.n46 VP.n45 28.8382
R1280 VP.n26 VP.n25 28.8382
R1281 VP.n14 VP.n13 28.8325
R1282 VP.n35 VP.n5 16.1487
R1283 VP.n42 VP.n1 16.1487
R1284 VP.n22 VP.n8 16.1487
R1285 VP.n15 VP.n12 16.1487
R1286 VP.n37 VP.n3 12.234
R1287 VP.n40 VP.n3 12.234
R1288 VP.n17 VP.n10 12.234
R1289 VP.n20 VP.n10 12.234
R1290 VP.n32 VP.n5 8.31928
R1291 VP.n45 VP.n1 8.31928
R1292 VP.n25 VP.n8 8.31928
R1293 VP.n28 VP.n7 0.285035
R1294 VP.n29 VP.n6 0.285035
R1295 VP.n48 VP.n0 0.285035
R1296 VP.n14 VP.n11 0.189894
R1297 VP.n18 VP.n11 0.189894
R1298 VP.n19 VP.n18 0.189894
R1299 VP.n19 VP.n9 0.189894
R1300 VP.n23 VP.n9 0.189894
R1301 VP.n24 VP.n23 0.189894
R1302 VP.n24 VP.n7 0.189894
R1303 VP.n33 VP.n6 0.189894
R1304 VP.n34 VP.n33 0.189894
R1305 VP.n34 VP.n4 0.189894
R1306 VP.n38 VP.n4 0.189894
R1307 VP.n39 VP.n38 0.189894
R1308 VP.n39 VP.n2 0.189894
R1309 VP.n43 VP.n2 0.189894
R1310 VP.n44 VP.n43 0.189894
R1311 VP.n44 VP.n0 0.189894
R1312 VP VP.n48 0.146778
R1313 VDD1.n1 VDD1.t2 75.1392
R1314 VDD1.n3 VDD1.t5 75.1392
R1315 VDD1.n5 VDD1.n4 70.727
R1316 VDD1.n1 VDD1.n0 69.761
R1317 VDD1.n7 VDD1.n6 69.7609
R1318 VDD1.n3 VDD1.n2 69.7608
R1319 VDD1.n7 VDD1.n5 35.6992
R1320 VDD1.n6 VDD1.t4 4.01673
R1321 VDD1.n6 VDD1.t7 4.01673
R1322 VDD1.n0 VDD1.t0 4.01673
R1323 VDD1.n0 VDD1.t3 4.01673
R1324 VDD1.n4 VDD1.t1 4.01673
R1325 VDD1.n4 VDD1.t9 4.01673
R1326 VDD1.n2 VDD1.t6 4.01673
R1327 VDD1.n2 VDD1.t8 4.01673
R1328 VDD1 VDD1.n7 0.963862
R1329 VDD1 VDD1.n1 0.399207
R1330 VDD1.n5 VDD1.n3 0.285671
C0 VDD2 VDD1 1.3094f
C1 VTAIL VP 4.34369f
C2 VTAIL VN 4.32944f
C3 VDD1 VP 4.10803f
C4 VDD2 VP 0.414695f
C5 VDD1 VN 0.150092f
C6 VDD2 VN 3.84999f
C7 VDD1 VTAIL 6.57668f
C8 VDD2 VTAIL 6.61924f
C9 VN VP 5.09585f
C10 VDD2 B 4.344955f
C11 VDD1 B 4.312795f
C12 VTAIL B 4.138837f
C13 VN B 11.06816f
C14 VP B 9.54395f
C15 VDD1.t2 B 0.950245f
C16 VDD1.t0 B 0.091487f
C17 VDD1.t3 B 0.091487f
C18 VDD1.n0 B 0.743497f
C19 VDD1.n1 B 0.662048f
C20 VDD1.t5 B 0.950241f
C21 VDD1.t6 B 0.091487f
C22 VDD1.t8 B 0.091487f
C23 VDD1.n2 B 0.743494f
C24 VDD1.n3 B 0.655373f
C25 VDD1.t1 B 0.091487f
C26 VDD1.t9 B 0.091487f
C27 VDD1.n4 B 0.74859f
C28 VDD1.n5 B 1.74116f
C29 VDD1.t4 B 0.091487f
C30 VDD1.t7 B 0.091487f
C31 VDD1.n6 B 0.743493f
C32 VDD1.n7 B 1.9269f
C33 VP.n0 B 0.048225f
C34 VP.t8 B 0.581949f
C35 VP.n1 B 0.241304f
C36 VP.n2 B 0.03614f
C37 VP.t1 B 0.581949f
C38 VP.n3 B 0.241304f
C39 VP.n4 B 0.03614f
C40 VP.t3 B 0.581949f
C41 VP.n5 B 0.241304f
C42 VP.n6 B 0.048225f
C43 VP.n7 B 0.048225f
C44 VP.t2 B 0.651158f
C45 VP.t5 B 0.581949f
C46 VP.n8 B 0.241304f
C47 VP.n9 B 0.03614f
C48 VP.t6 B 0.581949f
C49 VP.n10 B 0.241304f
C50 VP.n11 B 0.03614f
C51 VP.t9 B 0.581949f
C52 VP.n12 B 0.292375f
C53 VP.t7 B 0.697219f
C54 VP.n13 B 0.299684f
C55 VP.n14 B 0.191622f
C56 VP.n15 B 0.058733f
C57 VP.n16 B 0.029966f
C58 VP.n17 B 0.056241f
C59 VP.n18 B 0.03614f
C60 VP.n19 B 0.03614f
C61 VP.n20 B 0.056241f
C62 VP.n21 B 0.029966f
C63 VP.n22 B 0.058733f
C64 VP.n23 B 0.03614f
C65 VP.n24 B 0.03614f
C66 VP.n25 B 0.049539f
C67 VP.n26 B 0.032338f
C68 VP.n27 B 0.313158f
C69 VP.n28 B 1.42352f
C70 VP.n29 B 1.45549f
C71 VP.t4 B 0.651158f
C72 VP.n30 B 0.313158f
C73 VP.n31 B 0.032338f
C74 VP.n32 B 0.049539f
C75 VP.n33 B 0.03614f
C76 VP.n34 B 0.03614f
C77 VP.n35 B 0.058733f
C78 VP.n36 B 0.029966f
C79 VP.n37 B 0.056241f
C80 VP.n38 B 0.03614f
C81 VP.n39 B 0.03614f
C82 VP.n40 B 0.056241f
C83 VP.n41 B 0.029966f
C84 VP.n42 B 0.058733f
C85 VP.n43 B 0.03614f
C86 VP.n44 B 0.03614f
C87 VP.n45 B 0.049539f
C88 VP.n46 B 0.032338f
C89 VP.t0 B 0.651158f
C90 VP.n47 B 0.313158f
C91 VP.n48 B 0.033847f
C92 VTAIL.t8 B 0.108274f
C93 VTAIL.t17 B 0.108274f
C94 VTAIL.n0 B 0.812132f
C95 VTAIL.n1 B 0.450809f
C96 VTAIL.t0 B 1.03714f
C97 VTAIL.n2 B 0.546373f
C98 VTAIL.t2 B 0.108274f
C99 VTAIL.t1 B 0.108274f
C100 VTAIL.n3 B 0.812132f
C101 VTAIL.n4 B 0.495007f
C102 VTAIL.t19 B 0.108274f
C103 VTAIL.t6 B 0.108274f
C104 VTAIL.n5 B 0.812132f
C105 VTAIL.n6 B 1.37511f
C106 VTAIL.t10 B 0.108274f
C107 VTAIL.t15 B 0.108274f
C108 VTAIL.n7 B 0.812136f
C109 VTAIL.n8 B 1.3751f
C110 VTAIL.t14 B 0.108274f
C111 VTAIL.t12 B 0.108274f
C112 VTAIL.n9 B 0.812136f
C113 VTAIL.n10 B 0.495002f
C114 VTAIL.t9 B 1.03715f
C115 VTAIL.n11 B 0.546367f
C116 VTAIL.t4 B 0.108274f
C117 VTAIL.t3 B 0.108274f
C118 VTAIL.n12 B 0.812136f
C119 VTAIL.n13 B 0.476088f
C120 VTAIL.t7 B 0.108274f
C121 VTAIL.t5 B 0.108274f
C122 VTAIL.n14 B 0.812136f
C123 VTAIL.n15 B 0.495002f
C124 VTAIL.t18 B 1.03714f
C125 VTAIL.n16 B 1.32341f
C126 VTAIL.t11 B 1.03714f
C127 VTAIL.n17 B 1.32341f
C128 VTAIL.t13 B 0.108274f
C129 VTAIL.t16 B 0.108274f
C130 VTAIL.n18 B 0.812132f
C131 VTAIL.n19 B 0.398313f
C132 VDD2.t9 B 0.931146f
C133 VDD2.t8 B 0.089648f
C134 VDD2.t6 B 0.089648f
C135 VDD2.n0 B 0.728555f
C136 VDD2.n1 B 0.642203f
C137 VDD2.t7 B 0.089648f
C138 VDD2.t1 B 0.089648f
C139 VDD2.n2 B 0.733547f
C140 VDD2.n3 B 1.62695f
C141 VDD2.t4 B 0.924963f
C142 VDD2.n4 B 1.85907f
C143 VDD2.t5 B 0.089648f
C144 VDD2.t3 B 0.089648f
C145 VDD2.n5 B 0.728557f
C146 VDD2.n6 B 0.313569f
C147 VDD2.t2 B 0.089648f
C148 VDD2.t0 B 0.089648f
C149 VDD2.n7 B 0.733521f
C150 VN.n0 B 0.046976f
C151 VN.t1 B 0.566884f
C152 VN.n1 B 0.235057f
C153 VN.n2 B 0.035205f
C154 VN.t4 B 0.566884f
C155 VN.n3 B 0.235057f
C156 VN.n4 B 0.035205f
C157 VN.t0 B 0.566884f
C158 VN.n5 B 0.284806f
C159 VN.t9 B 0.67917f
C160 VN.n6 B 0.291926f
C161 VN.n7 B 0.186661f
C162 VN.n8 B 0.057212f
C163 VN.n9 B 0.02919f
C164 VN.n10 B 0.054785f
C165 VN.n11 B 0.035205f
C166 VN.n12 B 0.035205f
C167 VN.n13 B 0.054785f
C168 VN.n14 B 0.02919f
C169 VN.n15 B 0.057212f
C170 VN.n16 B 0.035205f
C171 VN.n17 B 0.035205f
C172 VN.n18 B 0.048257f
C173 VN.n19 B 0.031501f
C174 VN.t6 B 0.634301f
C175 VN.n20 B 0.305051f
C176 VN.n21 B 0.032971f
C177 VN.n22 B 0.046976f
C178 VN.t2 B 0.566884f
C179 VN.n23 B 0.235057f
C180 VN.n24 B 0.035205f
C181 VN.t3 B 0.566884f
C182 VN.n25 B 0.235057f
C183 VN.n26 B 0.035205f
C184 VN.t5 B 0.566884f
C185 VN.n27 B 0.284806f
C186 VN.t8 B 0.67917f
C187 VN.n28 B 0.291926f
C188 VN.n29 B 0.186661f
C189 VN.n30 B 0.057212f
C190 VN.n31 B 0.02919f
C191 VN.n32 B 0.054785f
C192 VN.n33 B 0.035205f
C193 VN.n34 B 0.035205f
C194 VN.n35 B 0.054785f
C195 VN.n36 B 0.02919f
C196 VN.n37 B 0.057212f
C197 VN.n38 B 0.035205f
C198 VN.n39 B 0.035205f
C199 VN.n40 B 0.048257f
C200 VN.n41 B 0.031501f
C201 VN.t7 B 0.634301f
C202 VN.n42 B 0.305051f
C203 VN.n43 B 1.40654f
.ends

