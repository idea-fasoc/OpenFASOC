* NGSPICE file created from diff_pair_sample_0572.ext - technology: sky130A

.subckt diff_pair_sample_0572 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=0 ps=0 w=19.77 l=1.26
X1 VDD1.t3 VP.t0 VTAIL.t4 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=3.26205 pd=20.1 as=7.7103 ps=40.32 w=19.77 l=1.26
X2 VDD1.t2 VP.t1 VTAIL.t7 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=3.26205 pd=20.1 as=7.7103 ps=40.32 w=19.77 l=1.26
X3 VTAIL.t2 VN.t0 VDD2.t3 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=3.26205 ps=20.1 w=19.77 l=1.26
X4 VDD2.t2 VN.t1 VTAIL.t1 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=3.26205 pd=20.1 as=7.7103 ps=40.32 w=19.77 l=1.26
X5 B.t8 B.t6 B.t7 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=0 ps=0 w=19.77 l=1.26
X6 B.t5 B.t3 B.t4 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=0 ps=0 w=19.77 l=1.26
X7 VDD2.t1 VN.t2 VTAIL.t3 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=3.26205 pd=20.1 as=7.7103 ps=40.32 w=19.77 l=1.26
X8 VTAIL.t0 VN.t3 VDD2.t0 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=3.26205 ps=20.1 w=19.77 l=1.26
X9 VTAIL.t5 VP.t2 VDD1.t1 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=3.26205 ps=20.1 w=19.77 l=1.26
X10 VTAIL.t6 VP.t3 VDD1.t0 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=3.26205 ps=20.1 w=19.77 l=1.26
X11 B.t2 B.t0 B.t1 w_n1924_n4922# sky130_fd_pr__pfet_01v8 ad=7.7103 pd=40.32 as=0 ps=0 w=19.77 l=1.26
R0 B.n504 B.n503 585
R1 B.n505 B.n86 585
R2 B.n507 B.n506 585
R3 B.n508 B.n85 585
R4 B.n510 B.n509 585
R5 B.n511 B.n84 585
R6 B.n513 B.n512 585
R7 B.n514 B.n83 585
R8 B.n516 B.n515 585
R9 B.n517 B.n82 585
R10 B.n519 B.n518 585
R11 B.n520 B.n81 585
R12 B.n522 B.n521 585
R13 B.n523 B.n80 585
R14 B.n525 B.n524 585
R15 B.n526 B.n79 585
R16 B.n528 B.n527 585
R17 B.n529 B.n78 585
R18 B.n531 B.n530 585
R19 B.n532 B.n77 585
R20 B.n534 B.n533 585
R21 B.n535 B.n76 585
R22 B.n537 B.n536 585
R23 B.n538 B.n75 585
R24 B.n540 B.n539 585
R25 B.n541 B.n74 585
R26 B.n543 B.n542 585
R27 B.n544 B.n73 585
R28 B.n546 B.n545 585
R29 B.n547 B.n72 585
R30 B.n549 B.n548 585
R31 B.n550 B.n71 585
R32 B.n552 B.n551 585
R33 B.n553 B.n70 585
R34 B.n555 B.n554 585
R35 B.n556 B.n69 585
R36 B.n558 B.n557 585
R37 B.n559 B.n68 585
R38 B.n561 B.n560 585
R39 B.n562 B.n67 585
R40 B.n564 B.n563 585
R41 B.n565 B.n66 585
R42 B.n567 B.n566 585
R43 B.n568 B.n65 585
R44 B.n570 B.n569 585
R45 B.n571 B.n64 585
R46 B.n573 B.n572 585
R47 B.n574 B.n63 585
R48 B.n576 B.n575 585
R49 B.n577 B.n62 585
R50 B.n579 B.n578 585
R51 B.n580 B.n61 585
R52 B.n582 B.n581 585
R53 B.n583 B.n60 585
R54 B.n585 B.n584 585
R55 B.n586 B.n59 585
R56 B.n588 B.n587 585
R57 B.n589 B.n58 585
R58 B.n591 B.n590 585
R59 B.n592 B.n57 585
R60 B.n594 B.n593 585
R61 B.n595 B.n56 585
R62 B.n597 B.n596 585
R63 B.n598 B.n55 585
R64 B.n600 B.n599 585
R65 B.n602 B.n601 585
R66 B.n603 B.n51 585
R67 B.n605 B.n604 585
R68 B.n606 B.n50 585
R69 B.n608 B.n607 585
R70 B.n609 B.n49 585
R71 B.n611 B.n610 585
R72 B.n612 B.n48 585
R73 B.n614 B.n613 585
R74 B.n616 B.n45 585
R75 B.n618 B.n617 585
R76 B.n619 B.n44 585
R77 B.n621 B.n620 585
R78 B.n622 B.n43 585
R79 B.n624 B.n623 585
R80 B.n625 B.n42 585
R81 B.n627 B.n626 585
R82 B.n628 B.n41 585
R83 B.n630 B.n629 585
R84 B.n631 B.n40 585
R85 B.n633 B.n632 585
R86 B.n634 B.n39 585
R87 B.n636 B.n635 585
R88 B.n637 B.n38 585
R89 B.n639 B.n638 585
R90 B.n640 B.n37 585
R91 B.n642 B.n641 585
R92 B.n643 B.n36 585
R93 B.n645 B.n644 585
R94 B.n646 B.n35 585
R95 B.n648 B.n647 585
R96 B.n649 B.n34 585
R97 B.n651 B.n650 585
R98 B.n652 B.n33 585
R99 B.n654 B.n653 585
R100 B.n655 B.n32 585
R101 B.n657 B.n656 585
R102 B.n658 B.n31 585
R103 B.n660 B.n659 585
R104 B.n661 B.n30 585
R105 B.n663 B.n662 585
R106 B.n664 B.n29 585
R107 B.n666 B.n665 585
R108 B.n667 B.n28 585
R109 B.n669 B.n668 585
R110 B.n670 B.n27 585
R111 B.n672 B.n671 585
R112 B.n673 B.n26 585
R113 B.n675 B.n674 585
R114 B.n676 B.n25 585
R115 B.n678 B.n677 585
R116 B.n679 B.n24 585
R117 B.n681 B.n680 585
R118 B.n682 B.n23 585
R119 B.n684 B.n683 585
R120 B.n685 B.n22 585
R121 B.n687 B.n686 585
R122 B.n688 B.n21 585
R123 B.n690 B.n689 585
R124 B.n691 B.n20 585
R125 B.n693 B.n692 585
R126 B.n694 B.n19 585
R127 B.n696 B.n695 585
R128 B.n697 B.n18 585
R129 B.n699 B.n698 585
R130 B.n700 B.n17 585
R131 B.n702 B.n701 585
R132 B.n703 B.n16 585
R133 B.n705 B.n704 585
R134 B.n706 B.n15 585
R135 B.n708 B.n707 585
R136 B.n709 B.n14 585
R137 B.n711 B.n710 585
R138 B.n712 B.n13 585
R139 B.n502 B.n87 585
R140 B.n501 B.n500 585
R141 B.n499 B.n88 585
R142 B.n498 B.n497 585
R143 B.n496 B.n89 585
R144 B.n495 B.n494 585
R145 B.n493 B.n90 585
R146 B.n492 B.n491 585
R147 B.n490 B.n91 585
R148 B.n489 B.n488 585
R149 B.n487 B.n92 585
R150 B.n486 B.n485 585
R151 B.n484 B.n93 585
R152 B.n483 B.n482 585
R153 B.n481 B.n94 585
R154 B.n480 B.n479 585
R155 B.n478 B.n95 585
R156 B.n477 B.n476 585
R157 B.n475 B.n96 585
R158 B.n474 B.n473 585
R159 B.n472 B.n97 585
R160 B.n471 B.n470 585
R161 B.n469 B.n98 585
R162 B.n468 B.n467 585
R163 B.n466 B.n99 585
R164 B.n465 B.n464 585
R165 B.n463 B.n100 585
R166 B.n462 B.n461 585
R167 B.n460 B.n101 585
R168 B.n459 B.n458 585
R169 B.n457 B.n102 585
R170 B.n456 B.n455 585
R171 B.n454 B.n103 585
R172 B.n453 B.n452 585
R173 B.n451 B.n104 585
R174 B.n450 B.n449 585
R175 B.n448 B.n105 585
R176 B.n447 B.n446 585
R177 B.n445 B.n106 585
R178 B.n444 B.n443 585
R179 B.n442 B.n107 585
R180 B.n441 B.n440 585
R181 B.n439 B.n108 585
R182 B.n438 B.n437 585
R183 B.n436 B.n109 585
R184 B.n226 B.n183 585
R185 B.n228 B.n227 585
R186 B.n229 B.n182 585
R187 B.n231 B.n230 585
R188 B.n232 B.n181 585
R189 B.n234 B.n233 585
R190 B.n235 B.n180 585
R191 B.n237 B.n236 585
R192 B.n238 B.n179 585
R193 B.n240 B.n239 585
R194 B.n241 B.n178 585
R195 B.n243 B.n242 585
R196 B.n244 B.n177 585
R197 B.n246 B.n245 585
R198 B.n247 B.n176 585
R199 B.n249 B.n248 585
R200 B.n250 B.n175 585
R201 B.n252 B.n251 585
R202 B.n253 B.n174 585
R203 B.n255 B.n254 585
R204 B.n256 B.n173 585
R205 B.n258 B.n257 585
R206 B.n259 B.n172 585
R207 B.n261 B.n260 585
R208 B.n262 B.n171 585
R209 B.n264 B.n263 585
R210 B.n265 B.n170 585
R211 B.n267 B.n266 585
R212 B.n268 B.n169 585
R213 B.n270 B.n269 585
R214 B.n271 B.n168 585
R215 B.n273 B.n272 585
R216 B.n274 B.n167 585
R217 B.n276 B.n275 585
R218 B.n277 B.n166 585
R219 B.n279 B.n278 585
R220 B.n280 B.n165 585
R221 B.n282 B.n281 585
R222 B.n283 B.n164 585
R223 B.n285 B.n284 585
R224 B.n286 B.n163 585
R225 B.n288 B.n287 585
R226 B.n289 B.n162 585
R227 B.n291 B.n290 585
R228 B.n292 B.n161 585
R229 B.n294 B.n293 585
R230 B.n295 B.n160 585
R231 B.n297 B.n296 585
R232 B.n298 B.n159 585
R233 B.n300 B.n299 585
R234 B.n301 B.n158 585
R235 B.n303 B.n302 585
R236 B.n304 B.n157 585
R237 B.n306 B.n305 585
R238 B.n307 B.n156 585
R239 B.n309 B.n308 585
R240 B.n310 B.n155 585
R241 B.n312 B.n311 585
R242 B.n313 B.n154 585
R243 B.n315 B.n314 585
R244 B.n316 B.n153 585
R245 B.n318 B.n317 585
R246 B.n319 B.n152 585
R247 B.n321 B.n320 585
R248 B.n322 B.n149 585
R249 B.n325 B.n324 585
R250 B.n326 B.n148 585
R251 B.n328 B.n327 585
R252 B.n329 B.n147 585
R253 B.n331 B.n330 585
R254 B.n332 B.n146 585
R255 B.n334 B.n333 585
R256 B.n335 B.n145 585
R257 B.n337 B.n336 585
R258 B.n339 B.n338 585
R259 B.n340 B.n141 585
R260 B.n342 B.n341 585
R261 B.n343 B.n140 585
R262 B.n345 B.n344 585
R263 B.n346 B.n139 585
R264 B.n348 B.n347 585
R265 B.n349 B.n138 585
R266 B.n351 B.n350 585
R267 B.n352 B.n137 585
R268 B.n354 B.n353 585
R269 B.n355 B.n136 585
R270 B.n357 B.n356 585
R271 B.n358 B.n135 585
R272 B.n360 B.n359 585
R273 B.n361 B.n134 585
R274 B.n363 B.n362 585
R275 B.n364 B.n133 585
R276 B.n366 B.n365 585
R277 B.n367 B.n132 585
R278 B.n369 B.n368 585
R279 B.n370 B.n131 585
R280 B.n372 B.n371 585
R281 B.n373 B.n130 585
R282 B.n375 B.n374 585
R283 B.n376 B.n129 585
R284 B.n378 B.n377 585
R285 B.n379 B.n128 585
R286 B.n381 B.n380 585
R287 B.n382 B.n127 585
R288 B.n384 B.n383 585
R289 B.n385 B.n126 585
R290 B.n387 B.n386 585
R291 B.n388 B.n125 585
R292 B.n390 B.n389 585
R293 B.n391 B.n124 585
R294 B.n393 B.n392 585
R295 B.n394 B.n123 585
R296 B.n396 B.n395 585
R297 B.n397 B.n122 585
R298 B.n399 B.n398 585
R299 B.n400 B.n121 585
R300 B.n402 B.n401 585
R301 B.n403 B.n120 585
R302 B.n405 B.n404 585
R303 B.n406 B.n119 585
R304 B.n408 B.n407 585
R305 B.n409 B.n118 585
R306 B.n411 B.n410 585
R307 B.n412 B.n117 585
R308 B.n414 B.n413 585
R309 B.n415 B.n116 585
R310 B.n417 B.n416 585
R311 B.n418 B.n115 585
R312 B.n420 B.n419 585
R313 B.n421 B.n114 585
R314 B.n423 B.n422 585
R315 B.n424 B.n113 585
R316 B.n426 B.n425 585
R317 B.n427 B.n112 585
R318 B.n429 B.n428 585
R319 B.n430 B.n111 585
R320 B.n432 B.n431 585
R321 B.n433 B.n110 585
R322 B.n435 B.n434 585
R323 B.n225 B.n224 585
R324 B.n223 B.n184 585
R325 B.n222 B.n221 585
R326 B.n220 B.n185 585
R327 B.n219 B.n218 585
R328 B.n217 B.n186 585
R329 B.n216 B.n215 585
R330 B.n214 B.n187 585
R331 B.n213 B.n212 585
R332 B.n211 B.n188 585
R333 B.n210 B.n209 585
R334 B.n208 B.n189 585
R335 B.n207 B.n206 585
R336 B.n205 B.n190 585
R337 B.n204 B.n203 585
R338 B.n202 B.n191 585
R339 B.n201 B.n200 585
R340 B.n199 B.n192 585
R341 B.n198 B.n197 585
R342 B.n196 B.n193 585
R343 B.n195 B.n194 585
R344 B.n2 B.n0 585
R345 B.n745 B.n1 585
R346 B.n744 B.n743 585
R347 B.n742 B.n3 585
R348 B.n741 B.n740 585
R349 B.n739 B.n4 585
R350 B.n738 B.n737 585
R351 B.n736 B.n5 585
R352 B.n735 B.n734 585
R353 B.n733 B.n6 585
R354 B.n732 B.n731 585
R355 B.n730 B.n7 585
R356 B.n729 B.n728 585
R357 B.n727 B.n8 585
R358 B.n726 B.n725 585
R359 B.n724 B.n9 585
R360 B.n723 B.n722 585
R361 B.n721 B.n10 585
R362 B.n720 B.n719 585
R363 B.n718 B.n11 585
R364 B.n717 B.n716 585
R365 B.n715 B.n12 585
R366 B.n714 B.n713 585
R367 B.n747 B.n746 585
R368 B.n142 B.t0 582.559
R369 B.n150 B.t6 582.559
R370 B.n46 B.t9 582.559
R371 B.n52 B.t3 582.559
R372 B.n224 B.n183 482.89
R373 B.n714 B.n13 482.89
R374 B.n434 B.n109 482.89
R375 B.n504 B.n87 482.89
R376 B.n224 B.n223 163.367
R377 B.n223 B.n222 163.367
R378 B.n222 B.n185 163.367
R379 B.n218 B.n185 163.367
R380 B.n218 B.n217 163.367
R381 B.n217 B.n216 163.367
R382 B.n216 B.n187 163.367
R383 B.n212 B.n187 163.367
R384 B.n212 B.n211 163.367
R385 B.n211 B.n210 163.367
R386 B.n210 B.n189 163.367
R387 B.n206 B.n189 163.367
R388 B.n206 B.n205 163.367
R389 B.n205 B.n204 163.367
R390 B.n204 B.n191 163.367
R391 B.n200 B.n191 163.367
R392 B.n200 B.n199 163.367
R393 B.n199 B.n198 163.367
R394 B.n198 B.n193 163.367
R395 B.n194 B.n193 163.367
R396 B.n194 B.n2 163.367
R397 B.n746 B.n2 163.367
R398 B.n746 B.n745 163.367
R399 B.n745 B.n744 163.367
R400 B.n744 B.n3 163.367
R401 B.n740 B.n3 163.367
R402 B.n740 B.n739 163.367
R403 B.n739 B.n738 163.367
R404 B.n738 B.n5 163.367
R405 B.n734 B.n5 163.367
R406 B.n734 B.n733 163.367
R407 B.n733 B.n732 163.367
R408 B.n732 B.n7 163.367
R409 B.n728 B.n7 163.367
R410 B.n728 B.n727 163.367
R411 B.n727 B.n726 163.367
R412 B.n726 B.n9 163.367
R413 B.n722 B.n9 163.367
R414 B.n722 B.n721 163.367
R415 B.n721 B.n720 163.367
R416 B.n720 B.n11 163.367
R417 B.n716 B.n11 163.367
R418 B.n716 B.n715 163.367
R419 B.n715 B.n714 163.367
R420 B.n228 B.n183 163.367
R421 B.n229 B.n228 163.367
R422 B.n230 B.n229 163.367
R423 B.n230 B.n181 163.367
R424 B.n234 B.n181 163.367
R425 B.n235 B.n234 163.367
R426 B.n236 B.n235 163.367
R427 B.n236 B.n179 163.367
R428 B.n240 B.n179 163.367
R429 B.n241 B.n240 163.367
R430 B.n242 B.n241 163.367
R431 B.n242 B.n177 163.367
R432 B.n246 B.n177 163.367
R433 B.n247 B.n246 163.367
R434 B.n248 B.n247 163.367
R435 B.n248 B.n175 163.367
R436 B.n252 B.n175 163.367
R437 B.n253 B.n252 163.367
R438 B.n254 B.n253 163.367
R439 B.n254 B.n173 163.367
R440 B.n258 B.n173 163.367
R441 B.n259 B.n258 163.367
R442 B.n260 B.n259 163.367
R443 B.n260 B.n171 163.367
R444 B.n264 B.n171 163.367
R445 B.n265 B.n264 163.367
R446 B.n266 B.n265 163.367
R447 B.n266 B.n169 163.367
R448 B.n270 B.n169 163.367
R449 B.n271 B.n270 163.367
R450 B.n272 B.n271 163.367
R451 B.n272 B.n167 163.367
R452 B.n276 B.n167 163.367
R453 B.n277 B.n276 163.367
R454 B.n278 B.n277 163.367
R455 B.n278 B.n165 163.367
R456 B.n282 B.n165 163.367
R457 B.n283 B.n282 163.367
R458 B.n284 B.n283 163.367
R459 B.n284 B.n163 163.367
R460 B.n288 B.n163 163.367
R461 B.n289 B.n288 163.367
R462 B.n290 B.n289 163.367
R463 B.n290 B.n161 163.367
R464 B.n294 B.n161 163.367
R465 B.n295 B.n294 163.367
R466 B.n296 B.n295 163.367
R467 B.n296 B.n159 163.367
R468 B.n300 B.n159 163.367
R469 B.n301 B.n300 163.367
R470 B.n302 B.n301 163.367
R471 B.n302 B.n157 163.367
R472 B.n306 B.n157 163.367
R473 B.n307 B.n306 163.367
R474 B.n308 B.n307 163.367
R475 B.n308 B.n155 163.367
R476 B.n312 B.n155 163.367
R477 B.n313 B.n312 163.367
R478 B.n314 B.n313 163.367
R479 B.n314 B.n153 163.367
R480 B.n318 B.n153 163.367
R481 B.n319 B.n318 163.367
R482 B.n320 B.n319 163.367
R483 B.n320 B.n149 163.367
R484 B.n325 B.n149 163.367
R485 B.n326 B.n325 163.367
R486 B.n327 B.n326 163.367
R487 B.n327 B.n147 163.367
R488 B.n331 B.n147 163.367
R489 B.n332 B.n331 163.367
R490 B.n333 B.n332 163.367
R491 B.n333 B.n145 163.367
R492 B.n337 B.n145 163.367
R493 B.n338 B.n337 163.367
R494 B.n338 B.n141 163.367
R495 B.n342 B.n141 163.367
R496 B.n343 B.n342 163.367
R497 B.n344 B.n343 163.367
R498 B.n344 B.n139 163.367
R499 B.n348 B.n139 163.367
R500 B.n349 B.n348 163.367
R501 B.n350 B.n349 163.367
R502 B.n350 B.n137 163.367
R503 B.n354 B.n137 163.367
R504 B.n355 B.n354 163.367
R505 B.n356 B.n355 163.367
R506 B.n356 B.n135 163.367
R507 B.n360 B.n135 163.367
R508 B.n361 B.n360 163.367
R509 B.n362 B.n361 163.367
R510 B.n362 B.n133 163.367
R511 B.n366 B.n133 163.367
R512 B.n367 B.n366 163.367
R513 B.n368 B.n367 163.367
R514 B.n368 B.n131 163.367
R515 B.n372 B.n131 163.367
R516 B.n373 B.n372 163.367
R517 B.n374 B.n373 163.367
R518 B.n374 B.n129 163.367
R519 B.n378 B.n129 163.367
R520 B.n379 B.n378 163.367
R521 B.n380 B.n379 163.367
R522 B.n380 B.n127 163.367
R523 B.n384 B.n127 163.367
R524 B.n385 B.n384 163.367
R525 B.n386 B.n385 163.367
R526 B.n386 B.n125 163.367
R527 B.n390 B.n125 163.367
R528 B.n391 B.n390 163.367
R529 B.n392 B.n391 163.367
R530 B.n392 B.n123 163.367
R531 B.n396 B.n123 163.367
R532 B.n397 B.n396 163.367
R533 B.n398 B.n397 163.367
R534 B.n398 B.n121 163.367
R535 B.n402 B.n121 163.367
R536 B.n403 B.n402 163.367
R537 B.n404 B.n403 163.367
R538 B.n404 B.n119 163.367
R539 B.n408 B.n119 163.367
R540 B.n409 B.n408 163.367
R541 B.n410 B.n409 163.367
R542 B.n410 B.n117 163.367
R543 B.n414 B.n117 163.367
R544 B.n415 B.n414 163.367
R545 B.n416 B.n415 163.367
R546 B.n416 B.n115 163.367
R547 B.n420 B.n115 163.367
R548 B.n421 B.n420 163.367
R549 B.n422 B.n421 163.367
R550 B.n422 B.n113 163.367
R551 B.n426 B.n113 163.367
R552 B.n427 B.n426 163.367
R553 B.n428 B.n427 163.367
R554 B.n428 B.n111 163.367
R555 B.n432 B.n111 163.367
R556 B.n433 B.n432 163.367
R557 B.n434 B.n433 163.367
R558 B.n438 B.n109 163.367
R559 B.n439 B.n438 163.367
R560 B.n440 B.n439 163.367
R561 B.n440 B.n107 163.367
R562 B.n444 B.n107 163.367
R563 B.n445 B.n444 163.367
R564 B.n446 B.n445 163.367
R565 B.n446 B.n105 163.367
R566 B.n450 B.n105 163.367
R567 B.n451 B.n450 163.367
R568 B.n452 B.n451 163.367
R569 B.n452 B.n103 163.367
R570 B.n456 B.n103 163.367
R571 B.n457 B.n456 163.367
R572 B.n458 B.n457 163.367
R573 B.n458 B.n101 163.367
R574 B.n462 B.n101 163.367
R575 B.n463 B.n462 163.367
R576 B.n464 B.n463 163.367
R577 B.n464 B.n99 163.367
R578 B.n468 B.n99 163.367
R579 B.n469 B.n468 163.367
R580 B.n470 B.n469 163.367
R581 B.n470 B.n97 163.367
R582 B.n474 B.n97 163.367
R583 B.n475 B.n474 163.367
R584 B.n476 B.n475 163.367
R585 B.n476 B.n95 163.367
R586 B.n480 B.n95 163.367
R587 B.n481 B.n480 163.367
R588 B.n482 B.n481 163.367
R589 B.n482 B.n93 163.367
R590 B.n486 B.n93 163.367
R591 B.n487 B.n486 163.367
R592 B.n488 B.n487 163.367
R593 B.n488 B.n91 163.367
R594 B.n492 B.n91 163.367
R595 B.n493 B.n492 163.367
R596 B.n494 B.n493 163.367
R597 B.n494 B.n89 163.367
R598 B.n498 B.n89 163.367
R599 B.n499 B.n498 163.367
R600 B.n500 B.n499 163.367
R601 B.n500 B.n87 163.367
R602 B.n710 B.n13 163.367
R603 B.n710 B.n709 163.367
R604 B.n709 B.n708 163.367
R605 B.n708 B.n15 163.367
R606 B.n704 B.n15 163.367
R607 B.n704 B.n703 163.367
R608 B.n703 B.n702 163.367
R609 B.n702 B.n17 163.367
R610 B.n698 B.n17 163.367
R611 B.n698 B.n697 163.367
R612 B.n697 B.n696 163.367
R613 B.n696 B.n19 163.367
R614 B.n692 B.n19 163.367
R615 B.n692 B.n691 163.367
R616 B.n691 B.n690 163.367
R617 B.n690 B.n21 163.367
R618 B.n686 B.n21 163.367
R619 B.n686 B.n685 163.367
R620 B.n685 B.n684 163.367
R621 B.n684 B.n23 163.367
R622 B.n680 B.n23 163.367
R623 B.n680 B.n679 163.367
R624 B.n679 B.n678 163.367
R625 B.n678 B.n25 163.367
R626 B.n674 B.n25 163.367
R627 B.n674 B.n673 163.367
R628 B.n673 B.n672 163.367
R629 B.n672 B.n27 163.367
R630 B.n668 B.n27 163.367
R631 B.n668 B.n667 163.367
R632 B.n667 B.n666 163.367
R633 B.n666 B.n29 163.367
R634 B.n662 B.n29 163.367
R635 B.n662 B.n661 163.367
R636 B.n661 B.n660 163.367
R637 B.n660 B.n31 163.367
R638 B.n656 B.n31 163.367
R639 B.n656 B.n655 163.367
R640 B.n655 B.n654 163.367
R641 B.n654 B.n33 163.367
R642 B.n650 B.n33 163.367
R643 B.n650 B.n649 163.367
R644 B.n649 B.n648 163.367
R645 B.n648 B.n35 163.367
R646 B.n644 B.n35 163.367
R647 B.n644 B.n643 163.367
R648 B.n643 B.n642 163.367
R649 B.n642 B.n37 163.367
R650 B.n638 B.n37 163.367
R651 B.n638 B.n637 163.367
R652 B.n637 B.n636 163.367
R653 B.n636 B.n39 163.367
R654 B.n632 B.n39 163.367
R655 B.n632 B.n631 163.367
R656 B.n631 B.n630 163.367
R657 B.n630 B.n41 163.367
R658 B.n626 B.n41 163.367
R659 B.n626 B.n625 163.367
R660 B.n625 B.n624 163.367
R661 B.n624 B.n43 163.367
R662 B.n620 B.n43 163.367
R663 B.n620 B.n619 163.367
R664 B.n619 B.n618 163.367
R665 B.n618 B.n45 163.367
R666 B.n613 B.n45 163.367
R667 B.n613 B.n612 163.367
R668 B.n612 B.n611 163.367
R669 B.n611 B.n49 163.367
R670 B.n607 B.n49 163.367
R671 B.n607 B.n606 163.367
R672 B.n606 B.n605 163.367
R673 B.n605 B.n51 163.367
R674 B.n601 B.n51 163.367
R675 B.n601 B.n600 163.367
R676 B.n600 B.n55 163.367
R677 B.n596 B.n55 163.367
R678 B.n596 B.n595 163.367
R679 B.n595 B.n594 163.367
R680 B.n594 B.n57 163.367
R681 B.n590 B.n57 163.367
R682 B.n590 B.n589 163.367
R683 B.n589 B.n588 163.367
R684 B.n588 B.n59 163.367
R685 B.n584 B.n59 163.367
R686 B.n584 B.n583 163.367
R687 B.n583 B.n582 163.367
R688 B.n582 B.n61 163.367
R689 B.n578 B.n61 163.367
R690 B.n578 B.n577 163.367
R691 B.n577 B.n576 163.367
R692 B.n576 B.n63 163.367
R693 B.n572 B.n63 163.367
R694 B.n572 B.n571 163.367
R695 B.n571 B.n570 163.367
R696 B.n570 B.n65 163.367
R697 B.n566 B.n65 163.367
R698 B.n566 B.n565 163.367
R699 B.n565 B.n564 163.367
R700 B.n564 B.n67 163.367
R701 B.n560 B.n67 163.367
R702 B.n560 B.n559 163.367
R703 B.n559 B.n558 163.367
R704 B.n558 B.n69 163.367
R705 B.n554 B.n69 163.367
R706 B.n554 B.n553 163.367
R707 B.n553 B.n552 163.367
R708 B.n552 B.n71 163.367
R709 B.n548 B.n71 163.367
R710 B.n548 B.n547 163.367
R711 B.n547 B.n546 163.367
R712 B.n546 B.n73 163.367
R713 B.n542 B.n73 163.367
R714 B.n542 B.n541 163.367
R715 B.n541 B.n540 163.367
R716 B.n540 B.n75 163.367
R717 B.n536 B.n75 163.367
R718 B.n536 B.n535 163.367
R719 B.n535 B.n534 163.367
R720 B.n534 B.n77 163.367
R721 B.n530 B.n77 163.367
R722 B.n530 B.n529 163.367
R723 B.n529 B.n528 163.367
R724 B.n528 B.n79 163.367
R725 B.n524 B.n79 163.367
R726 B.n524 B.n523 163.367
R727 B.n523 B.n522 163.367
R728 B.n522 B.n81 163.367
R729 B.n518 B.n81 163.367
R730 B.n518 B.n517 163.367
R731 B.n517 B.n516 163.367
R732 B.n516 B.n83 163.367
R733 B.n512 B.n83 163.367
R734 B.n512 B.n511 163.367
R735 B.n511 B.n510 163.367
R736 B.n510 B.n85 163.367
R737 B.n506 B.n85 163.367
R738 B.n506 B.n505 163.367
R739 B.n505 B.n504 163.367
R740 B.n142 B.t2 137.851
R741 B.n52 B.t4 137.851
R742 B.n150 B.t8 137.826
R743 B.n46 B.t10 137.826
R744 B.n143 B.t1 107.014
R745 B.n53 B.t5 107.014
R746 B.n151 B.t7 106.989
R747 B.n47 B.t11 106.989
R748 B.n144 B.n143 59.5399
R749 B.n323 B.n151 59.5399
R750 B.n615 B.n47 59.5399
R751 B.n54 B.n53 59.5399
R752 B.n713 B.n712 31.3761
R753 B.n503 B.n502 31.3761
R754 B.n436 B.n435 31.3761
R755 B.n226 B.n225 31.3761
R756 B.n143 B.n142 30.8369
R757 B.n151 B.n150 30.8369
R758 B.n47 B.n46 30.8369
R759 B.n53 B.n52 30.8369
R760 B B.n747 18.0485
R761 B.n712 B.n711 10.6151
R762 B.n711 B.n14 10.6151
R763 B.n707 B.n14 10.6151
R764 B.n707 B.n706 10.6151
R765 B.n706 B.n705 10.6151
R766 B.n705 B.n16 10.6151
R767 B.n701 B.n16 10.6151
R768 B.n701 B.n700 10.6151
R769 B.n700 B.n699 10.6151
R770 B.n699 B.n18 10.6151
R771 B.n695 B.n18 10.6151
R772 B.n695 B.n694 10.6151
R773 B.n694 B.n693 10.6151
R774 B.n693 B.n20 10.6151
R775 B.n689 B.n20 10.6151
R776 B.n689 B.n688 10.6151
R777 B.n688 B.n687 10.6151
R778 B.n687 B.n22 10.6151
R779 B.n683 B.n22 10.6151
R780 B.n683 B.n682 10.6151
R781 B.n682 B.n681 10.6151
R782 B.n681 B.n24 10.6151
R783 B.n677 B.n24 10.6151
R784 B.n677 B.n676 10.6151
R785 B.n676 B.n675 10.6151
R786 B.n675 B.n26 10.6151
R787 B.n671 B.n26 10.6151
R788 B.n671 B.n670 10.6151
R789 B.n670 B.n669 10.6151
R790 B.n669 B.n28 10.6151
R791 B.n665 B.n28 10.6151
R792 B.n665 B.n664 10.6151
R793 B.n664 B.n663 10.6151
R794 B.n663 B.n30 10.6151
R795 B.n659 B.n30 10.6151
R796 B.n659 B.n658 10.6151
R797 B.n658 B.n657 10.6151
R798 B.n657 B.n32 10.6151
R799 B.n653 B.n32 10.6151
R800 B.n653 B.n652 10.6151
R801 B.n652 B.n651 10.6151
R802 B.n651 B.n34 10.6151
R803 B.n647 B.n34 10.6151
R804 B.n647 B.n646 10.6151
R805 B.n646 B.n645 10.6151
R806 B.n645 B.n36 10.6151
R807 B.n641 B.n36 10.6151
R808 B.n641 B.n640 10.6151
R809 B.n640 B.n639 10.6151
R810 B.n639 B.n38 10.6151
R811 B.n635 B.n38 10.6151
R812 B.n635 B.n634 10.6151
R813 B.n634 B.n633 10.6151
R814 B.n633 B.n40 10.6151
R815 B.n629 B.n40 10.6151
R816 B.n629 B.n628 10.6151
R817 B.n628 B.n627 10.6151
R818 B.n627 B.n42 10.6151
R819 B.n623 B.n42 10.6151
R820 B.n623 B.n622 10.6151
R821 B.n622 B.n621 10.6151
R822 B.n621 B.n44 10.6151
R823 B.n617 B.n44 10.6151
R824 B.n617 B.n616 10.6151
R825 B.n614 B.n48 10.6151
R826 B.n610 B.n48 10.6151
R827 B.n610 B.n609 10.6151
R828 B.n609 B.n608 10.6151
R829 B.n608 B.n50 10.6151
R830 B.n604 B.n50 10.6151
R831 B.n604 B.n603 10.6151
R832 B.n603 B.n602 10.6151
R833 B.n599 B.n598 10.6151
R834 B.n598 B.n597 10.6151
R835 B.n597 B.n56 10.6151
R836 B.n593 B.n56 10.6151
R837 B.n593 B.n592 10.6151
R838 B.n592 B.n591 10.6151
R839 B.n591 B.n58 10.6151
R840 B.n587 B.n58 10.6151
R841 B.n587 B.n586 10.6151
R842 B.n586 B.n585 10.6151
R843 B.n585 B.n60 10.6151
R844 B.n581 B.n60 10.6151
R845 B.n581 B.n580 10.6151
R846 B.n580 B.n579 10.6151
R847 B.n579 B.n62 10.6151
R848 B.n575 B.n62 10.6151
R849 B.n575 B.n574 10.6151
R850 B.n574 B.n573 10.6151
R851 B.n573 B.n64 10.6151
R852 B.n569 B.n64 10.6151
R853 B.n569 B.n568 10.6151
R854 B.n568 B.n567 10.6151
R855 B.n567 B.n66 10.6151
R856 B.n563 B.n66 10.6151
R857 B.n563 B.n562 10.6151
R858 B.n562 B.n561 10.6151
R859 B.n561 B.n68 10.6151
R860 B.n557 B.n68 10.6151
R861 B.n557 B.n556 10.6151
R862 B.n556 B.n555 10.6151
R863 B.n555 B.n70 10.6151
R864 B.n551 B.n70 10.6151
R865 B.n551 B.n550 10.6151
R866 B.n550 B.n549 10.6151
R867 B.n549 B.n72 10.6151
R868 B.n545 B.n72 10.6151
R869 B.n545 B.n544 10.6151
R870 B.n544 B.n543 10.6151
R871 B.n543 B.n74 10.6151
R872 B.n539 B.n74 10.6151
R873 B.n539 B.n538 10.6151
R874 B.n538 B.n537 10.6151
R875 B.n537 B.n76 10.6151
R876 B.n533 B.n76 10.6151
R877 B.n533 B.n532 10.6151
R878 B.n532 B.n531 10.6151
R879 B.n531 B.n78 10.6151
R880 B.n527 B.n78 10.6151
R881 B.n527 B.n526 10.6151
R882 B.n526 B.n525 10.6151
R883 B.n525 B.n80 10.6151
R884 B.n521 B.n80 10.6151
R885 B.n521 B.n520 10.6151
R886 B.n520 B.n519 10.6151
R887 B.n519 B.n82 10.6151
R888 B.n515 B.n82 10.6151
R889 B.n515 B.n514 10.6151
R890 B.n514 B.n513 10.6151
R891 B.n513 B.n84 10.6151
R892 B.n509 B.n84 10.6151
R893 B.n509 B.n508 10.6151
R894 B.n508 B.n507 10.6151
R895 B.n507 B.n86 10.6151
R896 B.n503 B.n86 10.6151
R897 B.n437 B.n436 10.6151
R898 B.n437 B.n108 10.6151
R899 B.n441 B.n108 10.6151
R900 B.n442 B.n441 10.6151
R901 B.n443 B.n442 10.6151
R902 B.n443 B.n106 10.6151
R903 B.n447 B.n106 10.6151
R904 B.n448 B.n447 10.6151
R905 B.n449 B.n448 10.6151
R906 B.n449 B.n104 10.6151
R907 B.n453 B.n104 10.6151
R908 B.n454 B.n453 10.6151
R909 B.n455 B.n454 10.6151
R910 B.n455 B.n102 10.6151
R911 B.n459 B.n102 10.6151
R912 B.n460 B.n459 10.6151
R913 B.n461 B.n460 10.6151
R914 B.n461 B.n100 10.6151
R915 B.n465 B.n100 10.6151
R916 B.n466 B.n465 10.6151
R917 B.n467 B.n466 10.6151
R918 B.n467 B.n98 10.6151
R919 B.n471 B.n98 10.6151
R920 B.n472 B.n471 10.6151
R921 B.n473 B.n472 10.6151
R922 B.n473 B.n96 10.6151
R923 B.n477 B.n96 10.6151
R924 B.n478 B.n477 10.6151
R925 B.n479 B.n478 10.6151
R926 B.n479 B.n94 10.6151
R927 B.n483 B.n94 10.6151
R928 B.n484 B.n483 10.6151
R929 B.n485 B.n484 10.6151
R930 B.n485 B.n92 10.6151
R931 B.n489 B.n92 10.6151
R932 B.n490 B.n489 10.6151
R933 B.n491 B.n490 10.6151
R934 B.n491 B.n90 10.6151
R935 B.n495 B.n90 10.6151
R936 B.n496 B.n495 10.6151
R937 B.n497 B.n496 10.6151
R938 B.n497 B.n88 10.6151
R939 B.n501 B.n88 10.6151
R940 B.n502 B.n501 10.6151
R941 B.n227 B.n226 10.6151
R942 B.n227 B.n182 10.6151
R943 B.n231 B.n182 10.6151
R944 B.n232 B.n231 10.6151
R945 B.n233 B.n232 10.6151
R946 B.n233 B.n180 10.6151
R947 B.n237 B.n180 10.6151
R948 B.n238 B.n237 10.6151
R949 B.n239 B.n238 10.6151
R950 B.n239 B.n178 10.6151
R951 B.n243 B.n178 10.6151
R952 B.n244 B.n243 10.6151
R953 B.n245 B.n244 10.6151
R954 B.n245 B.n176 10.6151
R955 B.n249 B.n176 10.6151
R956 B.n250 B.n249 10.6151
R957 B.n251 B.n250 10.6151
R958 B.n251 B.n174 10.6151
R959 B.n255 B.n174 10.6151
R960 B.n256 B.n255 10.6151
R961 B.n257 B.n256 10.6151
R962 B.n257 B.n172 10.6151
R963 B.n261 B.n172 10.6151
R964 B.n262 B.n261 10.6151
R965 B.n263 B.n262 10.6151
R966 B.n263 B.n170 10.6151
R967 B.n267 B.n170 10.6151
R968 B.n268 B.n267 10.6151
R969 B.n269 B.n268 10.6151
R970 B.n269 B.n168 10.6151
R971 B.n273 B.n168 10.6151
R972 B.n274 B.n273 10.6151
R973 B.n275 B.n274 10.6151
R974 B.n275 B.n166 10.6151
R975 B.n279 B.n166 10.6151
R976 B.n280 B.n279 10.6151
R977 B.n281 B.n280 10.6151
R978 B.n281 B.n164 10.6151
R979 B.n285 B.n164 10.6151
R980 B.n286 B.n285 10.6151
R981 B.n287 B.n286 10.6151
R982 B.n287 B.n162 10.6151
R983 B.n291 B.n162 10.6151
R984 B.n292 B.n291 10.6151
R985 B.n293 B.n292 10.6151
R986 B.n293 B.n160 10.6151
R987 B.n297 B.n160 10.6151
R988 B.n298 B.n297 10.6151
R989 B.n299 B.n298 10.6151
R990 B.n299 B.n158 10.6151
R991 B.n303 B.n158 10.6151
R992 B.n304 B.n303 10.6151
R993 B.n305 B.n304 10.6151
R994 B.n305 B.n156 10.6151
R995 B.n309 B.n156 10.6151
R996 B.n310 B.n309 10.6151
R997 B.n311 B.n310 10.6151
R998 B.n311 B.n154 10.6151
R999 B.n315 B.n154 10.6151
R1000 B.n316 B.n315 10.6151
R1001 B.n317 B.n316 10.6151
R1002 B.n317 B.n152 10.6151
R1003 B.n321 B.n152 10.6151
R1004 B.n322 B.n321 10.6151
R1005 B.n324 B.n148 10.6151
R1006 B.n328 B.n148 10.6151
R1007 B.n329 B.n328 10.6151
R1008 B.n330 B.n329 10.6151
R1009 B.n330 B.n146 10.6151
R1010 B.n334 B.n146 10.6151
R1011 B.n335 B.n334 10.6151
R1012 B.n336 B.n335 10.6151
R1013 B.n340 B.n339 10.6151
R1014 B.n341 B.n340 10.6151
R1015 B.n341 B.n140 10.6151
R1016 B.n345 B.n140 10.6151
R1017 B.n346 B.n345 10.6151
R1018 B.n347 B.n346 10.6151
R1019 B.n347 B.n138 10.6151
R1020 B.n351 B.n138 10.6151
R1021 B.n352 B.n351 10.6151
R1022 B.n353 B.n352 10.6151
R1023 B.n353 B.n136 10.6151
R1024 B.n357 B.n136 10.6151
R1025 B.n358 B.n357 10.6151
R1026 B.n359 B.n358 10.6151
R1027 B.n359 B.n134 10.6151
R1028 B.n363 B.n134 10.6151
R1029 B.n364 B.n363 10.6151
R1030 B.n365 B.n364 10.6151
R1031 B.n365 B.n132 10.6151
R1032 B.n369 B.n132 10.6151
R1033 B.n370 B.n369 10.6151
R1034 B.n371 B.n370 10.6151
R1035 B.n371 B.n130 10.6151
R1036 B.n375 B.n130 10.6151
R1037 B.n376 B.n375 10.6151
R1038 B.n377 B.n376 10.6151
R1039 B.n377 B.n128 10.6151
R1040 B.n381 B.n128 10.6151
R1041 B.n382 B.n381 10.6151
R1042 B.n383 B.n382 10.6151
R1043 B.n383 B.n126 10.6151
R1044 B.n387 B.n126 10.6151
R1045 B.n388 B.n387 10.6151
R1046 B.n389 B.n388 10.6151
R1047 B.n389 B.n124 10.6151
R1048 B.n393 B.n124 10.6151
R1049 B.n394 B.n393 10.6151
R1050 B.n395 B.n394 10.6151
R1051 B.n395 B.n122 10.6151
R1052 B.n399 B.n122 10.6151
R1053 B.n400 B.n399 10.6151
R1054 B.n401 B.n400 10.6151
R1055 B.n401 B.n120 10.6151
R1056 B.n405 B.n120 10.6151
R1057 B.n406 B.n405 10.6151
R1058 B.n407 B.n406 10.6151
R1059 B.n407 B.n118 10.6151
R1060 B.n411 B.n118 10.6151
R1061 B.n412 B.n411 10.6151
R1062 B.n413 B.n412 10.6151
R1063 B.n413 B.n116 10.6151
R1064 B.n417 B.n116 10.6151
R1065 B.n418 B.n417 10.6151
R1066 B.n419 B.n418 10.6151
R1067 B.n419 B.n114 10.6151
R1068 B.n423 B.n114 10.6151
R1069 B.n424 B.n423 10.6151
R1070 B.n425 B.n424 10.6151
R1071 B.n425 B.n112 10.6151
R1072 B.n429 B.n112 10.6151
R1073 B.n430 B.n429 10.6151
R1074 B.n431 B.n430 10.6151
R1075 B.n431 B.n110 10.6151
R1076 B.n435 B.n110 10.6151
R1077 B.n225 B.n184 10.6151
R1078 B.n221 B.n184 10.6151
R1079 B.n221 B.n220 10.6151
R1080 B.n220 B.n219 10.6151
R1081 B.n219 B.n186 10.6151
R1082 B.n215 B.n186 10.6151
R1083 B.n215 B.n214 10.6151
R1084 B.n214 B.n213 10.6151
R1085 B.n213 B.n188 10.6151
R1086 B.n209 B.n188 10.6151
R1087 B.n209 B.n208 10.6151
R1088 B.n208 B.n207 10.6151
R1089 B.n207 B.n190 10.6151
R1090 B.n203 B.n190 10.6151
R1091 B.n203 B.n202 10.6151
R1092 B.n202 B.n201 10.6151
R1093 B.n201 B.n192 10.6151
R1094 B.n197 B.n192 10.6151
R1095 B.n197 B.n196 10.6151
R1096 B.n196 B.n195 10.6151
R1097 B.n195 B.n0 10.6151
R1098 B.n743 B.n1 10.6151
R1099 B.n743 B.n742 10.6151
R1100 B.n742 B.n741 10.6151
R1101 B.n741 B.n4 10.6151
R1102 B.n737 B.n4 10.6151
R1103 B.n737 B.n736 10.6151
R1104 B.n736 B.n735 10.6151
R1105 B.n735 B.n6 10.6151
R1106 B.n731 B.n6 10.6151
R1107 B.n731 B.n730 10.6151
R1108 B.n730 B.n729 10.6151
R1109 B.n729 B.n8 10.6151
R1110 B.n725 B.n8 10.6151
R1111 B.n725 B.n724 10.6151
R1112 B.n724 B.n723 10.6151
R1113 B.n723 B.n10 10.6151
R1114 B.n719 B.n10 10.6151
R1115 B.n719 B.n718 10.6151
R1116 B.n718 B.n717 10.6151
R1117 B.n717 B.n12 10.6151
R1118 B.n713 B.n12 10.6151
R1119 B.n615 B.n614 6.5566
R1120 B.n602 B.n54 6.5566
R1121 B.n324 B.n323 6.5566
R1122 B.n336 B.n144 6.5566
R1123 B.n616 B.n615 4.05904
R1124 B.n599 B.n54 4.05904
R1125 B.n323 B.n322 4.05904
R1126 B.n339 B.n144 4.05904
R1127 B.n747 B.n0 2.81026
R1128 B.n747 B.n1 2.81026
R1129 VP.n2 VP.t2 415.05
R1130 VP.n2 VP.t1 414.827
R1131 VP.n3 VP.t3 378.14
R1132 VP.n9 VP.t0 378.14
R1133 VP.n4 VP.n3 171.332
R1134 VP.n10 VP.n9 171.332
R1135 VP.n8 VP.n0 161.3
R1136 VP.n7 VP.n6 161.3
R1137 VP.n5 VP.n1 161.3
R1138 VP.n4 VP.n2 66.1874
R1139 VP.n7 VP.n1 40.4934
R1140 VP.n8 VP.n7 40.4934
R1141 VP.n3 VP.n1 14.436
R1142 VP.n9 VP.n8 14.436
R1143 VP.n5 VP.n4 0.189894
R1144 VP.n6 VP.n5 0.189894
R1145 VP.n6 VP.n0 0.189894
R1146 VP.n10 VP.n0 0.189894
R1147 VP VP.n10 0.0516364
R1148 VTAIL.n5 VTAIL.t5 54.433
R1149 VTAIL.n4 VTAIL.t1 54.433
R1150 VTAIL.n3 VTAIL.t0 54.433
R1151 VTAIL.n7 VTAIL.t3 54.4328
R1152 VTAIL.n0 VTAIL.t2 54.4328
R1153 VTAIL.n1 VTAIL.t4 54.4328
R1154 VTAIL.n2 VTAIL.t6 54.4328
R1155 VTAIL.n6 VTAIL.t7 54.4328
R1156 VTAIL.n7 VTAIL.n6 30.7807
R1157 VTAIL.n3 VTAIL.n2 30.7807
R1158 VTAIL.n4 VTAIL.n3 1.37119
R1159 VTAIL.n6 VTAIL.n5 1.37119
R1160 VTAIL.n2 VTAIL.n1 1.37119
R1161 VTAIL VTAIL.n0 0.744035
R1162 VTAIL VTAIL.n7 0.627655
R1163 VTAIL.n5 VTAIL.n4 0.470328
R1164 VTAIL.n1 VTAIL.n0 0.470328
R1165 VDD1 VDD1.n1 114.862
R1166 VDD1 VDD1.n0 69.5257
R1167 VDD1.n0 VDD1.t1 1.64466
R1168 VDD1.n0 VDD1.t2 1.64466
R1169 VDD1.n1 VDD1.t0 1.64466
R1170 VDD1.n1 VDD1.t3 1.64466
R1171 VN.n0 VN.t0 415.05
R1172 VN.n1 VN.t1 415.05
R1173 VN.n0 VN.t2 414.827
R1174 VN.n1 VN.t3 414.827
R1175 VN VN.n1 66.568
R1176 VN VN.n0 18.2006
R1177 VDD2.n2 VDD2.n0 114.338
R1178 VDD2.n2 VDD2.n1 69.4675
R1179 VDD2.n1 VDD2.t0 1.64466
R1180 VDD2.n1 VDD2.t2 1.64466
R1181 VDD2.n0 VDD2.t3 1.64466
R1182 VDD2.n0 VDD2.t1 1.64466
R1183 VDD2 VDD2.n2 0.0586897
C0 VN w_n1924_n4922# 3.15994f
C1 VTAIL w_n1924_n4922# 5.9245f
C2 VP VDD1 6.51361f
C3 VDD2 VDD1 0.698925f
C4 VDD2 VP 0.308853f
C5 B VDD1 1.23481f
C6 B VP 1.344f
C7 VDD2 B 1.26512f
C8 VN VDD1 0.147603f
C9 VTAIL VDD1 8.25864f
C10 VN VP 6.66476f
C11 VTAIL VP 5.74698f
C12 VDD2 VN 6.35276f
C13 VDD2 VTAIL 8.303861f
C14 B VN 0.945418f
C15 B VTAIL 6.49774f
C16 VDD1 w_n1924_n4922# 1.39126f
C17 VN VTAIL 5.73288f
C18 VP w_n1924_n4922# 3.40389f
C19 VDD2 w_n1924_n4922# 1.41763f
C20 B w_n1924_n4922# 9.77487f
C21 VDD2 VSUBS 0.937297f
C22 VDD1 VSUBS 6.12363f
C23 VTAIL VSUBS 1.337695f
C24 VN VSUBS 5.78275f
C25 VP VSUBS 1.862512f
C26 B VSUBS 3.767359f
C27 w_n1924_n4922# VSUBS 0.115648p
C28 VDD2.t3 VSUBS 0.42026f
C29 VDD2.t1 VSUBS 0.42026f
C30 VDD2.n0 VSUBS 4.49312f
C31 VDD2.t0 VSUBS 0.42026f
C32 VDD2.t2 VSUBS 0.42026f
C33 VDD2.n1 VSUBS 3.54632f
C34 VDD2.n2 VSUBS 4.85492f
C35 VN.t0 VSUBS 3.1269f
C36 VN.t2 VSUBS 3.12622f
C37 VN.n0 VSUBS 2.25634f
C38 VN.t1 VSUBS 3.1269f
C39 VN.t3 VSUBS 3.12622f
C40 VN.n1 VSUBS 4.05407f
C41 VDD1.t1 VSUBS 0.420278f
C42 VDD1.t2 VSUBS 0.420278f
C43 VDD1.n0 VSUBS 3.54702f
C44 VDD1.t0 VSUBS 0.420278f
C45 VDD1.t3 VSUBS 0.420278f
C46 VDD1.n1 VSUBS 4.52109f
C47 VTAIL.t2 VSUBS 3.53309f
C48 VTAIL.n0 VSUBS 0.703084f
C49 VTAIL.t4 VSUBS 3.53309f
C50 VTAIL.n1 VSUBS 0.746682f
C51 VTAIL.t6 VSUBS 3.53309f
C52 VTAIL.n2 VSUBS 2.28713f
C53 VTAIL.t0 VSUBS 3.53309f
C54 VTAIL.n3 VSUBS 2.28713f
C55 VTAIL.t1 VSUBS 3.53309f
C56 VTAIL.n4 VSUBS 0.746681f
C57 VTAIL.t5 VSUBS 3.53309f
C58 VTAIL.n5 VSUBS 0.746681f
C59 VTAIL.t7 VSUBS 3.53309f
C60 VTAIL.n6 VSUBS 2.28713f
C61 VTAIL.t3 VSUBS 3.53309f
C62 VTAIL.n7 VSUBS 2.23544f
C63 VP.n0 VSUBS 0.044716f
C64 VP.t0 VSUBS 3.06896f
C65 VP.n1 VSUBS 0.072f
C66 VP.t2 VSUBS 3.17847f
C67 VP.t1 VSUBS 3.17779f
C68 VP.n2 VSUBS 4.09585f
C69 VP.t3 VSUBS 3.06896f
C70 VP.n3 VSUBS 1.16439f
C71 VP.n4 VSUBS 3.00738f
C72 VP.n5 VSUBS 0.044716f
C73 VP.n6 VSUBS 0.044716f
C74 VP.n7 VSUBS 0.036148f
C75 VP.n8 VSUBS 0.072f
C76 VP.n9 VSUBS 1.16439f
C77 VP.n10 VSUBS 0.039797f
C78 B.n0 VSUBS 0.004426f
C79 B.n1 VSUBS 0.004426f
C80 B.n2 VSUBS 0.006999f
C81 B.n3 VSUBS 0.006999f
C82 B.n4 VSUBS 0.006999f
C83 B.n5 VSUBS 0.006999f
C84 B.n6 VSUBS 0.006999f
C85 B.n7 VSUBS 0.006999f
C86 B.n8 VSUBS 0.006999f
C87 B.n9 VSUBS 0.006999f
C88 B.n10 VSUBS 0.006999f
C89 B.n11 VSUBS 0.006999f
C90 B.n12 VSUBS 0.006999f
C91 B.n13 VSUBS 0.016636f
C92 B.n14 VSUBS 0.006999f
C93 B.n15 VSUBS 0.006999f
C94 B.n16 VSUBS 0.006999f
C95 B.n17 VSUBS 0.006999f
C96 B.n18 VSUBS 0.006999f
C97 B.n19 VSUBS 0.006999f
C98 B.n20 VSUBS 0.006999f
C99 B.n21 VSUBS 0.006999f
C100 B.n22 VSUBS 0.006999f
C101 B.n23 VSUBS 0.006999f
C102 B.n24 VSUBS 0.006999f
C103 B.n25 VSUBS 0.006999f
C104 B.n26 VSUBS 0.006999f
C105 B.n27 VSUBS 0.006999f
C106 B.n28 VSUBS 0.006999f
C107 B.n29 VSUBS 0.006999f
C108 B.n30 VSUBS 0.006999f
C109 B.n31 VSUBS 0.006999f
C110 B.n32 VSUBS 0.006999f
C111 B.n33 VSUBS 0.006999f
C112 B.n34 VSUBS 0.006999f
C113 B.n35 VSUBS 0.006999f
C114 B.n36 VSUBS 0.006999f
C115 B.n37 VSUBS 0.006999f
C116 B.n38 VSUBS 0.006999f
C117 B.n39 VSUBS 0.006999f
C118 B.n40 VSUBS 0.006999f
C119 B.n41 VSUBS 0.006999f
C120 B.n42 VSUBS 0.006999f
C121 B.n43 VSUBS 0.006999f
C122 B.n44 VSUBS 0.006999f
C123 B.n45 VSUBS 0.006999f
C124 B.t11 VSUBS 0.671465f
C125 B.t10 VSUBS 0.684142f
C126 B.t9 VSUBS 1.03879f
C127 B.n46 VSUBS 0.274496f
C128 B.n47 VSUBS 0.066644f
C129 B.n48 VSUBS 0.006999f
C130 B.n49 VSUBS 0.006999f
C131 B.n50 VSUBS 0.006999f
C132 B.n51 VSUBS 0.006999f
C133 B.t5 VSUBS 0.671436f
C134 B.t4 VSUBS 0.684117f
C135 B.t3 VSUBS 1.03879f
C136 B.n52 VSUBS 0.274521f
C137 B.n53 VSUBS 0.066674f
C138 B.n54 VSUBS 0.016216f
C139 B.n55 VSUBS 0.006999f
C140 B.n56 VSUBS 0.006999f
C141 B.n57 VSUBS 0.006999f
C142 B.n58 VSUBS 0.006999f
C143 B.n59 VSUBS 0.006999f
C144 B.n60 VSUBS 0.006999f
C145 B.n61 VSUBS 0.006999f
C146 B.n62 VSUBS 0.006999f
C147 B.n63 VSUBS 0.006999f
C148 B.n64 VSUBS 0.006999f
C149 B.n65 VSUBS 0.006999f
C150 B.n66 VSUBS 0.006999f
C151 B.n67 VSUBS 0.006999f
C152 B.n68 VSUBS 0.006999f
C153 B.n69 VSUBS 0.006999f
C154 B.n70 VSUBS 0.006999f
C155 B.n71 VSUBS 0.006999f
C156 B.n72 VSUBS 0.006999f
C157 B.n73 VSUBS 0.006999f
C158 B.n74 VSUBS 0.006999f
C159 B.n75 VSUBS 0.006999f
C160 B.n76 VSUBS 0.006999f
C161 B.n77 VSUBS 0.006999f
C162 B.n78 VSUBS 0.006999f
C163 B.n79 VSUBS 0.006999f
C164 B.n80 VSUBS 0.006999f
C165 B.n81 VSUBS 0.006999f
C166 B.n82 VSUBS 0.006999f
C167 B.n83 VSUBS 0.006999f
C168 B.n84 VSUBS 0.006999f
C169 B.n85 VSUBS 0.006999f
C170 B.n86 VSUBS 0.006999f
C171 B.n87 VSUBS 0.015271f
C172 B.n88 VSUBS 0.006999f
C173 B.n89 VSUBS 0.006999f
C174 B.n90 VSUBS 0.006999f
C175 B.n91 VSUBS 0.006999f
C176 B.n92 VSUBS 0.006999f
C177 B.n93 VSUBS 0.006999f
C178 B.n94 VSUBS 0.006999f
C179 B.n95 VSUBS 0.006999f
C180 B.n96 VSUBS 0.006999f
C181 B.n97 VSUBS 0.006999f
C182 B.n98 VSUBS 0.006999f
C183 B.n99 VSUBS 0.006999f
C184 B.n100 VSUBS 0.006999f
C185 B.n101 VSUBS 0.006999f
C186 B.n102 VSUBS 0.006999f
C187 B.n103 VSUBS 0.006999f
C188 B.n104 VSUBS 0.006999f
C189 B.n105 VSUBS 0.006999f
C190 B.n106 VSUBS 0.006999f
C191 B.n107 VSUBS 0.006999f
C192 B.n108 VSUBS 0.006999f
C193 B.n109 VSUBS 0.015271f
C194 B.n110 VSUBS 0.006999f
C195 B.n111 VSUBS 0.006999f
C196 B.n112 VSUBS 0.006999f
C197 B.n113 VSUBS 0.006999f
C198 B.n114 VSUBS 0.006999f
C199 B.n115 VSUBS 0.006999f
C200 B.n116 VSUBS 0.006999f
C201 B.n117 VSUBS 0.006999f
C202 B.n118 VSUBS 0.006999f
C203 B.n119 VSUBS 0.006999f
C204 B.n120 VSUBS 0.006999f
C205 B.n121 VSUBS 0.006999f
C206 B.n122 VSUBS 0.006999f
C207 B.n123 VSUBS 0.006999f
C208 B.n124 VSUBS 0.006999f
C209 B.n125 VSUBS 0.006999f
C210 B.n126 VSUBS 0.006999f
C211 B.n127 VSUBS 0.006999f
C212 B.n128 VSUBS 0.006999f
C213 B.n129 VSUBS 0.006999f
C214 B.n130 VSUBS 0.006999f
C215 B.n131 VSUBS 0.006999f
C216 B.n132 VSUBS 0.006999f
C217 B.n133 VSUBS 0.006999f
C218 B.n134 VSUBS 0.006999f
C219 B.n135 VSUBS 0.006999f
C220 B.n136 VSUBS 0.006999f
C221 B.n137 VSUBS 0.006999f
C222 B.n138 VSUBS 0.006999f
C223 B.n139 VSUBS 0.006999f
C224 B.n140 VSUBS 0.006999f
C225 B.n141 VSUBS 0.006999f
C226 B.t1 VSUBS 0.671436f
C227 B.t2 VSUBS 0.684117f
C228 B.t0 VSUBS 1.03879f
C229 B.n142 VSUBS 0.274521f
C230 B.n143 VSUBS 0.066674f
C231 B.n144 VSUBS 0.016216f
C232 B.n145 VSUBS 0.006999f
C233 B.n146 VSUBS 0.006999f
C234 B.n147 VSUBS 0.006999f
C235 B.n148 VSUBS 0.006999f
C236 B.n149 VSUBS 0.006999f
C237 B.t7 VSUBS 0.671465f
C238 B.t8 VSUBS 0.684142f
C239 B.t6 VSUBS 1.03879f
C240 B.n150 VSUBS 0.274496f
C241 B.n151 VSUBS 0.066644f
C242 B.n152 VSUBS 0.006999f
C243 B.n153 VSUBS 0.006999f
C244 B.n154 VSUBS 0.006999f
C245 B.n155 VSUBS 0.006999f
C246 B.n156 VSUBS 0.006999f
C247 B.n157 VSUBS 0.006999f
C248 B.n158 VSUBS 0.006999f
C249 B.n159 VSUBS 0.006999f
C250 B.n160 VSUBS 0.006999f
C251 B.n161 VSUBS 0.006999f
C252 B.n162 VSUBS 0.006999f
C253 B.n163 VSUBS 0.006999f
C254 B.n164 VSUBS 0.006999f
C255 B.n165 VSUBS 0.006999f
C256 B.n166 VSUBS 0.006999f
C257 B.n167 VSUBS 0.006999f
C258 B.n168 VSUBS 0.006999f
C259 B.n169 VSUBS 0.006999f
C260 B.n170 VSUBS 0.006999f
C261 B.n171 VSUBS 0.006999f
C262 B.n172 VSUBS 0.006999f
C263 B.n173 VSUBS 0.006999f
C264 B.n174 VSUBS 0.006999f
C265 B.n175 VSUBS 0.006999f
C266 B.n176 VSUBS 0.006999f
C267 B.n177 VSUBS 0.006999f
C268 B.n178 VSUBS 0.006999f
C269 B.n179 VSUBS 0.006999f
C270 B.n180 VSUBS 0.006999f
C271 B.n181 VSUBS 0.006999f
C272 B.n182 VSUBS 0.006999f
C273 B.n183 VSUBS 0.016636f
C274 B.n184 VSUBS 0.006999f
C275 B.n185 VSUBS 0.006999f
C276 B.n186 VSUBS 0.006999f
C277 B.n187 VSUBS 0.006999f
C278 B.n188 VSUBS 0.006999f
C279 B.n189 VSUBS 0.006999f
C280 B.n190 VSUBS 0.006999f
C281 B.n191 VSUBS 0.006999f
C282 B.n192 VSUBS 0.006999f
C283 B.n193 VSUBS 0.006999f
C284 B.n194 VSUBS 0.006999f
C285 B.n195 VSUBS 0.006999f
C286 B.n196 VSUBS 0.006999f
C287 B.n197 VSUBS 0.006999f
C288 B.n198 VSUBS 0.006999f
C289 B.n199 VSUBS 0.006999f
C290 B.n200 VSUBS 0.006999f
C291 B.n201 VSUBS 0.006999f
C292 B.n202 VSUBS 0.006999f
C293 B.n203 VSUBS 0.006999f
C294 B.n204 VSUBS 0.006999f
C295 B.n205 VSUBS 0.006999f
C296 B.n206 VSUBS 0.006999f
C297 B.n207 VSUBS 0.006999f
C298 B.n208 VSUBS 0.006999f
C299 B.n209 VSUBS 0.006999f
C300 B.n210 VSUBS 0.006999f
C301 B.n211 VSUBS 0.006999f
C302 B.n212 VSUBS 0.006999f
C303 B.n213 VSUBS 0.006999f
C304 B.n214 VSUBS 0.006999f
C305 B.n215 VSUBS 0.006999f
C306 B.n216 VSUBS 0.006999f
C307 B.n217 VSUBS 0.006999f
C308 B.n218 VSUBS 0.006999f
C309 B.n219 VSUBS 0.006999f
C310 B.n220 VSUBS 0.006999f
C311 B.n221 VSUBS 0.006999f
C312 B.n222 VSUBS 0.006999f
C313 B.n223 VSUBS 0.006999f
C314 B.n224 VSUBS 0.015271f
C315 B.n225 VSUBS 0.015271f
C316 B.n226 VSUBS 0.016636f
C317 B.n227 VSUBS 0.006999f
C318 B.n228 VSUBS 0.006999f
C319 B.n229 VSUBS 0.006999f
C320 B.n230 VSUBS 0.006999f
C321 B.n231 VSUBS 0.006999f
C322 B.n232 VSUBS 0.006999f
C323 B.n233 VSUBS 0.006999f
C324 B.n234 VSUBS 0.006999f
C325 B.n235 VSUBS 0.006999f
C326 B.n236 VSUBS 0.006999f
C327 B.n237 VSUBS 0.006999f
C328 B.n238 VSUBS 0.006999f
C329 B.n239 VSUBS 0.006999f
C330 B.n240 VSUBS 0.006999f
C331 B.n241 VSUBS 0.006999f
C332 B.n242 VSUBS 0.006999f
C333 B.n243 VSUBS 0.006999f
C334 B.n244 VSUBS 0.006999f
C335 B.n245 VSUBS 0.006999f
C336 B.n246 VSUBS 0.006999f
C337 B.n247 VSUBS 0.006999f
C338 B.n248 VSUBS 0.006999f
C339 B.n249 VSUBS 0.006999f
C340 B.n250 VSUBS 0.006999f
C341 B.n251 VSUBS 0.006999f
C342 B.n252 VSUBS 0.006999f
C343 B.n253 VSUBS 0.006999f
C344 B.n254 VSUBS 0.006999f
C345 B.n255 VSUBS 0.006999f
C346 B.n256 VSUBS 0.006999f
C347 B.n257 VSUBS 0.006999f
C348 B.n258 VSUBS 0.006999f
C349 B.n259 VSUBS 0.006999f
C350 B.n260 VSUBS 0.006999f
C351 B.n261 VSUBS 0.006999f
C352 B.n262 VSUBS 0.006999f
C353 B.n263 VSUBS 0.006999f
C354 B.n264 VSUBS 0.006999f
C355 B.n265 VSUBS 0.006999f
C356 B.n266 VSUBS 0.006999f
C357 B.n267 VSUBS 0.006999f
C358 B.n268 VSUBS 0.006999f
C359 B.n269 VSUBS 0.006999f
C360 B.n270 VSUBS 0.006999f
C361 B.n271 VSUBS 0.006999f
C362 B.n272 VSUBS 0.006999f
C363 B.n273 VSUBS 0.006999f
C364 B.n274 VSUBS 0.006999f
C365 B.n275 VSUBS 0.006999f
C366 B.n276 VSUBS 0.006999f
C367 B.n277 VSUBS 0.006999f
C368 B.n278 VSUBS 0.006999f
C369 B.n279 VSUBS 0.006999f
C370 B.n280 VSUBS 0.006999f
C371 B.n281 VSUBS 0.006999f
C372 B.n282 VSUBS 0.006999f
C373 B.n283 VSUBS 0.006999f
C374 B.n284 VSUBS 0.006999f
C375 B.n285 VSUBS 0.006999f
C376 B.n286 VSUBS 0.006999f
C377 B.n287 VSUBS 0.006999f
C378 B.n288 VSUBS 0.006999f
C379 B.n289 VSUBS 0.006999f
C380 B.n290 VSUBS 0.006999f
C381 B.n291 VSUBS 0.006999f
C382 B.n292 VSUBS 0.006999f
C383 B.n293 VSUBS 0.006999f
C384 B.n294 VSUBS 0.006999f
C385 B.n295 VSUBS 0.006999f
C386 B.n296 VSUBS 0.006999f
C387 B.n297 VSUBS 0.006999f
C388 B.n298 VSUBS 0.006999f
C389 B.n299 VSUBS 0.006999f
C390 B.n300 VSUBS 0.006999f
C391 B.n301 VSUBS 0.006999f
C392 B.n302 VSUBS 0.006999f
C393 B.n303 VSUBS 0.006999f
C394 B.n304 VSUBS 0.006999f
C395 B.n305 VSUBS 0.006999f
C396 B.n306 VSUBS 0.006999f
C397 B.n307 VSUBS 0.006999f
C398 B.n308 VSUBS 0.006999f
C399 B.n309 VSUBS 0.006999f
C400 B.n310 VSUBS 0.006999f
C401 B.n311 VSUBS 0.006999f
C402 B.n312 VSUBS 0.006999f
C403 B.n313 VSUBS 0.006999f
C404 B.n314 VSUBS 0.006999f
C405 B.n315 VSUBS 0.006999f
C406 B.n316 VSUBS 0.006999f
C407 B.n317 VSUBS 0.006999f
C408 B.n318 VSUBS 0.006999f
C409 B.n319 VSUBS 0.006999f
C410 B.n320 VSUBS 0.006999f
C411 B.n321 VSUBS 0.006999f
C412 B.n322 VSUBS 0.004837f
C413 B.n323 VSUBS 0.016216f
C414 B.n324 VSUBS 0.005661f
C415 B.n325 VSUBS 0.006999f
C416 B.n326 VSUBS 0.006999f
C417 B.n327 VSUBS 0.006999f
C418 B.n328 VSUBS 0.006999f
C419 B.n329 VSUBS 0.006999f
C420 B.n330 VSUBS 0.006999f
C421 B.n331 VSUBS 0.006999f
C422 B.n332 VSUBS 0.006999f
C423 B.n333 VSUBS 0.006999f
C424 B.n334 VSUBS 0.006999f
C425 B.n335 VSUBS 0.006999f
C426 B.n336 VSUBS 0.005661f
C427 B.n337 VSUBS 0.006999f
C428 B.n338 VSUBS 0.006999f
C429 B.n339 VSUBS 0.004837f
C430 B.n340 VSUBS 0.006999f
C431 B.n341 VSUBS 0.006999f
C432 B.n342 VSUBS 0.006999f
C433 B.n343 VSUBS 0.006999f
C434 B.n344 VSUBS 0.006999f
C435 B.n345 VSUBS 0.006999f
C436 B.n346 VSUBS 0.006999f
C437 B.n347 VSUBS 0.006999f
C438 B.n348 VSUBS 0.006999f
C439 B.n349 VSUBS 0.006999f
C440 B.n350 VSUBS 0.006999f
C441 B.n351 VSUBS 0.006999f
C442 B.n352 VSUBS 0.006999f
C443 B.n353 VSUBS 0.006999f
C444 B.n354 VSUBS 0.006999f
C445 B.n355 VSUBS 0.006999f
C446 B.n356 VSUBS 0.006999f
C447 B.n357 VSUBS 0.006999f
C448 B.n358 VSUBS 0.006999f
C449 B.n359 VSUBS 0.006999f
C450 B.n360 VSUBS 0.006999f
C451 B.n361 VSUBS 0.006999f
C452 B.n362 VSUBS 0.006999f
C453 B.n363 VSUBS 0.006999f
C454 B.n364 VSUBS 0.006999f
C455 B.n365 VSUBS 0.006999f
C456 B.n366 VSUBS 0.006999f
C457 B.n367 VSUBS 0.006999f
C458 B.n368 VSUBS 0.006999f
C459 B.n369 VSUBS 0.006999f
C460 B.n370 VSUBS 0.006999f
C461 B.n371 VSUBS 0.006999f
C462 B.n372 VSUBS 0.006999f
C463 B.n373 VSUBS 0.006999f
C464 B.n374 VSUBS 0.006999f
C465 B.n375 VSUBS 0.006999f
C466 B.n376 VSUBS 0.006999f
C467 B.n377 VSUBS 0.006999f
C468 B.n378 VSUBS 0.006999f
C469 B.n379 VSUBS 0.006999f
C470 B.n380 VSUBS 0.006999f
C471 B.n381 VSUBS 0.006999f
C472 B.n382 VSUBS 0.006999f
C473 B.n383 VSUBS 0.006999f
C474 B.n384 VSUBS 0.006999f
C475 B.n385 VSUBS 0.006999f
C476 B.n386 VSUBS 0.006999f
C477 B.n387 VSUBS 0.006999f
C478 B.n388 VSUBS 0.006999f
C479 B.n389 VSUBS 0.006999f
C480 B.n390 VSUBS 0.006999f
C481 B.n391 VSUBS 0.006999f
C482 B.n392 VSUBS 0.006999f
C483 B.n393 VSUBS 0.006999f
C484 B.n394 VSUBS 0.006999f
C485 B.n395 VSUBS 0.006999f
C486 B.n396 VSUBS 0.006999f
C487 B.n397 VSUBS 0.006999f
C488 B.n398 VSUBS 0.006999f
C489 B.n399 VSUBS 0.006999f
C490 B.n400 VSUBS 0.006999f
C491 B.n401 VSUBS 0.006999f
C492 B.n402 VSUBS 0.006999f
C493 B.n403 VSUBS 0.006999f
C494 B.n404 VSUBS 0.006999f
C495 B.n405 VSUBS 0.006999f
C496 B.n406 VSUBS 0.006999f
C497 B.n407 VSUBS 0.006999f
C498 B.n408 VSUBS 0.006999f
C499 B.n409 VSUBS 0.006999f
C500 B.n410 VSUBS 0.006999f
C501 B.n411 VSUBS 0.006999f
C502 B.n412 VSUBS 0.006999f
C503 B.n413 VSUBS 0.006999f
C504 B.n414 VSUBS 0.006999f
C505 B.n415 VSUBS 0.006999f
C506 B.n416 VSUBS 0.006999f
C507 B.n417 VSUBS 0.006999f
C508 B.n418 VSUBS 0.006999f
C509 B.n419 VSUBS 0.006999f
C510 B.n420 VSUBS 0.006999f
C511 B.n421 VSUBS 0.006999f
C512 B.n422 VSUBS 0.006999f
C513 B.n423 VSUBS 0.006999f
C514 B.n424 VSUBS 0.006999f
C515 B.n425 VSUBS 0.006999f
C516 B.n426 VSUBS 0.006999f
C517 B.n427 VSUBS 0.006999f
C518 B.n428 VSUBS 0.006999f
C519 B.n429 VSUBS 0.006999f
C520 B.n430 VSUBS 0.006999f
C521 B.n431 VSUBS 0.006999f
C522 B.n432 VSUBS 0.006999f
C523 B.n433 VSUBS 0.006999f
C524 B.n434 VSUBS 0.016636f
C525 B.n435 VSUBS 0.016636f
C526 B.n436 VSUBS 0.015271f
C527 B.n437 VSUBS 0.006999f
C528 B.n438 VSUBS 0.006999f
C529 B.n439 VSUBS 0.006999f
C530 B.n440 VSUBS 0.006999f
C531 B.n441 VSUBS 0.006999f
C532 B.n442 VSUBS 0.006999f
C533 B.n443 VSUBS 0.006999f
C534 B.n444 VSUBS 0.006999f
C535 B.n445 VSUBS 0.006999f
C536 B.n446 VSUBS 0.006999f
C537 B.n447 VSUBS 0.006999f
C538 B.n448 VSUBS 0.006999f
C539 B.n449 VSUBS 0.006999f
C540 B.n450 VSUBS 0.006999f
C541 B.n451 VSUBS 0.006999f
C542 B.n452 VSUBS 0.006999f
C543 B.n453 VSUBS 0.006999f
C544 B.n454 VSUBS 0.006999f
C545 B.n455 VSUBS 0.006999f
C546 B.n456 VSUBS 0.006999f
C547 B.n457 VSUBS 0.006999f
C548 B.n458 VSUBS 0.006999f
C549 B.n459 VSUBS 0.006999f
C550 B.n460 VSUBS 0.006999f
C551 B.n461 VSUBS 0.006999f
C552 B.n462 VSUBS 0.006999f
C553 B.n463 VSUBS 0.006999f
C554 B.n464 VSUBS 0.006999f
C555 B.n465 VSUBS 0.006999f
C556 B.n466 VSUBS 0.006999f
C557 B.n467 VSUBS 0.006999f
C558 B.n468 VSUBS 0.006999f
C559 B.n469 VSUBS 0.006999f
C560 B.n470 VSUBS 0.006999f
C561 B.n471 VSUBS 0.006999f
C562 B.n472 VSUBS 0.006999f
C563 B.n473 VSUBS 0.006999f
C564 B.n474 VSUBS 0.006999f
C565 B.n475 VSUBS 0.006999f
C566 B.n476 VSUBS 0.006999f
C567 B.n477 VSUBS 0.006999f
C568 B.n478 VSUBS 0.006999f
C569 B.n479 VSUBS 0.006999f
C570 B.n480 VSUBS 0.006999f
C571 B.n481 VSUBS 0.006999f
C572 B.n482 VSUBS 0.006999f
C573 B.n483 VSUBS 0.006999f
C574 B.n484 VSUBS 0.006999f
C575 B.n485 VSUBS 0.006999f
C576 B.n486 VSUBS 0.006999f
C577 B.n487 VSUBS 0.006999f
C578 B.n488 VSUBS 0.006999f
C579 B.n489 VSUBS 0.006999f
C580 B.n490 VSUBS 0.006999f
C581 B.n491 VSUBS 0.006999f
C582 B.n492 VSUBS 0.006999f
C583 B.n493 VSUBS 0.006999f
C584 B.n494 VSUBS 0.006999f
C585 B.n495 VSUBS 0.006999f
C586 B.n496 VSUBS 0.006999f
C587 B.n497 VSUBS 0.006999f
C588 B.n498 VSUBS 0.006999f
C589 B.n499 VSUBS 0.006999f
C590 B.n500 VSUBS 0.006999f
C591 B.n501 VSUBS 0.006999f
C592 B.n502 VSUBS 0.016132f
C593 B.n503 VSUBS 0.015775f
C594 B.n504 VSUBS 0.016636f
C595 B.n505 VSUBS 0.006999f
C596 B.n506 VSUBS 0.006999f
C597 B.n507 VSUBS 0.006999f
C598 B.n508 VSUBS 0.006999f
C599 B.n509 VSUBS 0.006999f
C600 B.n510 VSUBS 0.006999f
C601 B.n511 VSUBS 0.006999f
C602 B.n512 VSUBS 0.006999f
C603 B.n513 VSUBS 0.006999f
C604 B.n514 VSUBS 0.006999f
C605 B.n515 VSUBS 0.006999f
C606 B.n516 VSUBS 0.006999f
C607 B.n517 VSUBS 0.006999f
C608 B.n518 VSUBS 0.006999f
C609 B.n519 VSUBS 0.006999f
C610 B.n520 VSUBS 0.006999f
C611 B.n521 VSUBS 0.006999f
C612 B.n522 VSUBS 0.006999f
C613 B.n523 VSUBS 0.006999f
C614 B.n524 VSUBS 0.006999f
C615 B.n525 VSUBS 0.006999f
C616 B.n526 VSUBS 0.006999f
C617 B.n527 VSUBS 0.006999f
C618 B.n528 VSUBS 0.006999f
C619 B.n529 VSUBS 0.006999f
C620 B.n530 VSUBS 0.006999f
C621 B.n531 VSUBS 0.006999f
C622 B.n532 VSUBS 0.006999f
C623 B.n533 VSUBS 0.006999f
C624 B.n534 VSUBS 0.006999f
C625 B.n535 VSUBS 0.006999f
C626 B.n536 VSUBS 0.006999f
C627 B.n537 VSUBS 0.006999f
C628 B.n538 VSUBS 0.006999f
C629 B.n539 VSUBS 0.006999f
C630 B.n540 VSUBS 0.006999f
C631 B.n541 VSUBS 0.006999f
C632 B.n542 VSUBS 0.006999f
C633 B.n543 VSUBS 0.006999f
C634 B.n544 VSUBS 0.006999f
C635 B.n545 VSUBS 0.006999f
C636 B.n546 VSUBS 0.006999f
C637 B.n547 VSUBS 0.006999f
C638 B.n548 VSUBS 0.006999f
C639 B.n549 VSUBS 0.006999f
C640 B.n550 VSUBS 0.006999f
C641 B.n551 VSUBS 0.006999f
C642 B.n552 VSUBS 0.006999f
C643 B.n553 VSUBS 0.006999f
C644 B.n554 VSUBS 0.006999f
C645 B.n555 VSUBS 0.006999f
C646 B.n556 VSUBS 0.006999f
C647 B.n557 VSUBS 0.006999f
C648 B.n558 VSUBS 0.006999f
C649 B.n559 VSUBS 0.006999f
C650 B.n560 VSUBS 0.006999f
C651 B.n561 VSUBS 0.006999f
C652 B.n562 VSUBS 0.006999f
C653 B.n563 VSUBS 0.006999f
C654 B.n564 VSUBS 0.006999f
C655 B.n565 VSUBS 0.006999f
C656 B.n566 VSUBS 0.006999f
C657 B.n567 VSUBS 0.006999f
C658 B.n568 VSUBS 0.006999f
C659 B.n569 VSUBS 0.006999f
C660 B.n570 VSUBS 0.006999f
C661 B.n571 VSUBS 0.006999f
C662 B.n572 VSUBS 0.006999f
C663 B.n573 VSUBS 0.006999f
C664 B.n574 VSUBS 0.006999f
C665 B.n575 VSUBS 0.006999f
C666 B.n576 VSUBS 0.006999f
C667 B.n577 VSUBS 0.006999f
C668 B.n578 VSUBS 0.006999f
C669 B.n579 VSUBS 0.006999f
C670 B.n580 VSUBS 0.006999f
C671 B.n581 VSUBS 0.006999f
C672 B.n582 VSUBS 0.006999f
C673 B.n583 VSUBS 0.006999f
C674 B.n584 VSUBS 0.006999f
C675 B.n585 VSUBS 0.006999f
C676 B.n586 VSUBS 0.006999f
C677 B.n587 VSUBS 0.006999f
C678 B.n588 VSUBS 0.006999f
C679 B.n589 VSUBS 0.006999f
C680 B.n590 VSUBS 0.006999f
C681 B.n591 VSUBS 0.006999f
C682 B.n592 VSUBS 0.006999f
C683 B.n593 VSUBS 0.006999f
C684 B.n594 VSUBS 0.006999f
C685 B.n595 VSUBS 0.006999f
C686 B.n596 VSUBS 0.006999f
C687 B.n597 VSUBS 0.006999f
C688 B.n598 VSUBS 0.006999f
C689 B.n599 VSUBS 0.004837f
C690 B.n600 VSUBS 0.006999f
C691 B.n601 VSUBS 0.006999f
C692 B.n602 VSUBS 0.005661f
C693 B.n603 VSUBS 0.006999f
C694 B.n604 VSUBS 0.006999f
C695 B.n605 VSUBS 0.006999f
C696 B.n606 VSUBS 0.006999f
C697 B.n607 VSUBS 0.006999f
C698 B.n608 VSUBS 0.006999f
C699 B.n609 VSUBS 0.006999f
C700 B.n610 VSUBS 0.006999f
C701 B.n611 VSUBS 0.006999f
C702 B.n612 VSUBS 0.006999f
C703 B.n613 VSUBS 0.006999f
C704 B.n614 VSUBS 0.005661f
C705 B.n615 VSUBS 0.016216f
C706 B.n616 VSUBS 0.004837f
C707 B.n617 VSUBS 0.006999f
C708 B.n618 VSUBS 0.006999f
C709 B.n619 VSUBS 0.006999f
C710 B.n620 VSUBS 0.006999f
C711 B.n621 VSUBS 0.006999f
C712 B.n622 VSUBS 0.006999f
C713 B.n623 VSUBS 0.006999f
C714 B.n624 VSUBS 0.006999f
C715 B.n625 VSUBS 0.006999f
C716 B.n626 VSUBS 0.006999f
C717 B.n627 VSUBS 0.006999f
C718 B.n628 VSUBS 0.006999f
C719 B.n629 VSUBS 0.006999f
C720 B.n630 VSUBS 0.006999f
C721 B.n631 VSUBS 0.006999f
C722 B.n632 VSUBS 0.006999f
C723 B.n633 VSUBS 0.006999f
C724 B.n634 VSUBS 0.006999f
C725 B.n635 VSUBS 0.006999f
C726 B.n636 VSUBS 0.006999f
C727 B.n637 VSUBS 0.006999f
C728 B.n638 VSUBS 0.006999f
C729 B.n639 VSUBS 0.006999f
C730 B.n640 VSUBS 0.006999f
C731 B.n641 VSUBS 0.006999f
C732 B.n642 VSUBS 0.006999f
C733 B.n643 VSUBS 0.006999f
C734 B.n644 VSUBS 0.006999f
C735 B.n645 VSUBS 0.006999f
C736 B.n646 VSUBS 0.006999f
C737 B.n647 VSUBS 0.006999f
C738 B.n648 VSUBS 0.006999f
C739 B.n649 VSUBS 0.006999f
C740 B.n650 VSUBS 0.006999f
C741 B.n651 VSUBS 0.006999f
C742 B.n652 VSUBS 0.006999f
C743 B.n653 VSUBS 0.006999f
C744 B.n654 VSUBS 0.006999f
C745 B.n655 VSUBS 0.006999f
C746 B.n656 VSUBS 0.006999f
C747 B.n657 VSUBS 0.006999f
C748 B.n658 VSUBS 0.006999f
C749 B.n659 VSUBS 0.006999f
C750 B.n660 VSUBS 0.006999f
C751 B.n661 VSUBS 0.006999f
C752 B.n662 VSUBS 0.006999f
C753 B.n663 VSUBS 0.006999f
C754 B.n664 VSUBS 0.006999f
C755 B.n665 VSUBS 0.006999f
C756 B.n666 VSUBS 0.006999f
C757 B.n667 VSUBS 0.006999f
C758 B.n668 VSUBS 0.006999f
C759 B.n669 VSUBS 0.006999f
C760 B.n670 VSUBS 0.006999f
C761 B.n671 VSUBS 0.006999f
C762 B.n672 VSUBS 0.006999f
C763 B.n673 VSUBS 0.006999f
C764 B.n674 VSUBS 0.006999f
C765 B.n675 VSUBS 0.006999f
C766 B.n676 VSUBS 0.006999f
C767 B.n677 VSUBS 0.006999f
C768 B.n678 VSUBS 0.006999f
C769 B.n679 VSUBS 0.006999f
C770 B.n680 VSUBS 0.006999f
C771 B.n681 VSUBS 0.006999f
C772 B.n682 VSUBS 0.006999f
C773 B.n683 VSUBS 0.006999f
C774 B.n684 VSUBS 0.006999f
C775 B.n685 VSUBS 0.006999f
C776 B.n686 VSUBS 0.006999f
C777 B.n687 VSUBS 0.006999f
C778 B.n688 VSUBS 0.006999f
C779 B.n689 VSUBS 0.006999f
C780 B.n690 VSUBS 0.006999f
C781 B.n691 VSUBS 0.006999f
C782 B.n692 VSUBS 0.006999f
C783 B.n693 VSUBS 0.006999f
C784 B.n694 VSUBS 0.006999f
C785 B.n695 VSUBS 0.006999f
C786 B.n696 VSUBS 0.006999f
C787 B.n697 VSUBS 0.006999f
C788 B.n698 VSUBS 0.006999f
C789 B.n699 VSUBS 0.006999f
C790 B.n700 VSUBS 0.006999f
C791 B.n701 VSUBS 0.006999f
C792 B.n702 VSUBS 0.006999f
C793 B.n703 VSUBS 0.006999f
C794 B.n704 VSUBS 0.006999f
C795 B.n705 VSUBS 0.006999f
C796 B.n706 VSUBS 0.006999f
C797 B.n707 VSUBS 0.006999f
C798 B.n708 VSUBS 0.006999f
C799 B.n709 VSUBS 0.006999f
C800 B.n710 VSUBS 0.006999f
C801 B.n711 VSUBS 0.006999f
C802 B.n712 VSUBS 0.016636f
C803 B.n713 VSUBS 0.015271f
C804 B.n714 VSUBS 0.015271f
C805 B.n715 VSUBS 0.006999f
C806 B.n716 VSUBS 0.006999f
C807 B.n717 VSUBS 0.006999f
C808 B.n718 VSUBS 0.006999f
C809 B.n719 VSUBS 0.006999f
C810 B.n720 VSUBS 0.006999f
C811 B.n721 VSUBS 0.006999f
C812 B.n722 VSUBS 0.006999f
C813 B.n723 VSUBS 0.006999f
C814 B.n724 VSUBS 0.006999f
C815 B.n725 VSUBS 0.006999f
C816 B.n726 VSUBS 0.006999f
C817 B.n727 VSUBS 0.006999f
C818 B.n728 VSUBS 0.006999f
C819 B.n729 VSUBS 0.006999f
C820 B.n730 VSUBS 0.006999f
C821 B.n731 VSUBS 0.006999f
C822 B.n732 VSUBS 0.006999f
C823 B.n733 VSUBS 0.006999f
C824 B.n734 VSUBS 0.006999f
C825 B.n735 VSUBS 0.006999f
C826 B.n736 VSUBS 0.006999f
C827 B.n737 VSUBS 0.006999f
C828 B.n738 VSUBS 0.006999f
C829 B.n739 VSUBS 0.006999f
C830 B.n740 VSUBS 0.006999f
C831 B.n741 VSUBS 0.006999f
C832 B.n742 VSUBS 0.006999f
C833 B.n743 VSUBS 0.006999f
C834 B.n744 VSUBS 0.006999f
C835 B.n745 VSUBS 0.006999f
C836 B.n746 VSUBS 0.006999f
C837 B.n747 VSUBS 0.015848f
.ends

