* NGSPICE file created from diff_pair_sample_1336.ext - technology: sky130A

.subckt diff_pair_sample_1336 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X1 VTAIL.t17 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X2 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=0 ps=0 w=16.21 l=2.87
X3 VDD1.t7 VP.t2 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=2.67465 ps=16.54 w=16.21 l=2.87
X4 VTAIL.t0 VN.t0 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X5 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=0 ps=0 w=16.21 l=2.87
X6 VTAIL.t15 VP.t3 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X7 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=0 ps=0 w=16.21 l=2.87
X8 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X9 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X10 VDD1.t4 VP.t4 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X11 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X12 VDD1.t3 VP.t5 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=6.3219 ps=33.2 w=16.21 l=2.87
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=0 ps=0 w=16.21 l=2.87
X14 VDD2.t5 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=6.3219 ps=33.2 w=16.21 l=2.87
X15 VTAIL.t12 VP.t6 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X16 VDD1.t1 VP.t7 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=6.3219 ps=33.2 w=16.21 l=2.87
X17 VDD2.t4 VN.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=2.67465 ps=16.54 w=16.21 l=2.87
X18 VDD1.t0 VP.t8 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X19 VTAIL.t19 VN.t6 VDD2.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X20 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=2.67465 ps=16.54 w=16.21 l=2.87
X21 VDD2.t1 VN.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=2.67465 ps=16.54 w=16.21 l=2.87
X22 VDD2.t0 VN.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.67465 pd=16.54 as=6.3219 ps=33.2 w=16.21 l=2.87
X23 VDD1.t9 VP.t9 VTAIL.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.3219 pd=33.2 as=2.67465 ps=16.54 w=16.21 l=2.87
R0 VP.n25 VP.t2 167.798
R1 VP.n27 VP.n26 161.3
R2 VP.n28 VP.n23 161.3
R3 VP.n30 VP.n29 161.3
R4 VP.n31 VP.n22 161.3
R5 VP.n33 VP.n32 161.3
R6 VP.n34 VP.n21 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n20 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n19 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n18 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n47 VP.n17 161.3
R15 VP.n49 VP.n48 161.3
R16 VP.n50 VP.n16 161.3
R17 VP.n52 VP.n51 161.3
R18 VP.n53 VP.n15 161.3
R19 VP.n55 VP.n54 161.3
R20 VP.n97 VP.n96 161.3
R21 VP.n95 VP.n1 161.3
R22 VP.n94 VP.n93 161.3
R23 VP.n92 VP.n2 161.3
R24 VP.n91 VP.n90 161.3
R25 VP.n89 VP.n3 161.3
R26 VP.n87 VP.n86 161.3
R27 VP.n85 VP.n4 161.3
R28 VP.n84 VP.n83 161.3
R29 VP.n82 VP.n5 161.3
R30 VP.n81 VP.n80 161.3
R31 VP.n79 VP.n6 161.3
R32 VP.n78 VP.n77 161.3
R33 VP.n76 VP.n7 161.3
R34 VP.n75 VP.n74 161.3
R35 VP.n73 VP.n8 161.3
R36 VP.n72 VP.n71 161.3
R37 VP.n70 VP.n9 161.3
R38 VP.n69 VP.n68 161.3
R39 VP.n67 VP.n66 161.3
R40 VP.n65 VP.n11 161.3
R41 VP.n64 VP.n63 161.3
R42 VP.n62 VP.n12 161.3
R43 VP.n61 VP.n60 161.3
R44 VP.n59 VP.n13 161.3
R45 VP.n77 VP.t8 136.119
R46 VP.n58 VP.t9 136.119
R47 VP.n10 VP.t1 136.119
R48 VP.n88 VP.t0 136.119
R49 VP.n0 VP.t7 136.119
R50 VP.n35 VP.t4 136.119
R51 VP.n14 VP.t5 136.119
R52 VP.n46 VP.t6 136.119
R53 VP.n24 VP.t3 136.119
R54 VP.n58 VP.n57 70.4938
R55 VP.n98 VP.n0 70.4938
R56 VP.n56 VP.n14 70.4938
R57 VP.n25 VP.n24 63.8389
R58 VP.n57 VP.n56 57.8554
R59 VP.n64 VP.n12 56.5193
R60 VP.n94 VP.n2 56.5193
R61 VP.n52 VP.n16 56.5193
R62 VP.n71 VP.n8 50.2061
R63 VP.n83 VP.n82 50.2061
R64 VP.n41 VP.n40 50.2061
R65 VP.n29 VP.n22 50.2061
R66 VP.n75 VP.n8 30.7807
R67 VP.n82 VP.n81 30.7807
R68 VP.n40 VP.n39 30.7807
R69 VP.n33 VP.n22 30.7807
R70 VP.n60 VP.n59 24.4675
R71 VP.n60 VP.n12 24.4675
R72 VP.n65 VP.n64 24.4675
R73 VP.n66 VP.n65 24.4675
R74 VP.n70 VP.n69 24.4675
R75 VP.n71 VP.n70 24.4675
R76 VP.n76 VP.n75 24.4675
R77 VP.n77 VP.n76 24.4675
R78 VP.n77 VP.n6 24.4675
R79 VP.n81 VP.n6 24.4675
R80 VP.n83 VP.n4 24.4675
R81 VP.n87 VP.n4 24.4675
R82 VP.n90 VP.n89 24.4675
R83 VP.n90 VP.n2 24.4675
R84 VP.n95 VP.n94 24.4675
R85 VP.n96 VP.n95 24.4675
R86 VP.n53 VP.n52 24.4675
R87 VP.n54 VP.n53 24.4675
R88 VP.n41 VP.n18 24.4675
R89 VP.n45 VP.n18 24.4675
R90 VP.n48 VP.n47 24.4675
R91 VP.n48 VP.n16 24.4675
R92 VP.n34 VP.n33 24.4675
R93 VP.n35 VP.n34 24.4675
R94 VP.n35 VP.n20 24.4675
R95 VP.n39 VP.n20 24.4675
R96 VP.n28 VP.n27 24.4675
R97 VP.n29 VP.n28 24.4675
R98 VP.n59 VP.n58 19.5741
R99 VP.n96 VP.n0 19.5741
R100 VP.n54 VP.n14 19.5741
R101 VP.n66 VP.n10 14.6807
R102 VP.n89 VP.n88 14.6807
R103 VP.n47 VP.n46 14.6807
R104 VP.n69 VP.n10 9.7873
R105 VP.n88 VP.n87 9.7873
R106 VP.n46 VP.n45 9.7873
R107 VP.n27 VP.n24 9.7873
R108 VP.n26 VP.n25 5.58426
R109 VP.n56 VP.n55 0.354971
R110 VP.n57 VP.n13 0.354971
R111 VP.n98 VP.n97 0.354971
R112 VP VP.n98 0.26696
R113 VP.n26 VP.n23 0.189894
R114 VP.n30 VP.n23 0.189894
R115 VP.n31 VP.n30 0.189894
R116 VP.n32 VP.n31 0.189894
R117 VP.n32 VP.n21 0.189894
R118 VP.n36 VP.n21 0.189894
R119 VP.n37 VP.n36 0.189894
R120 VP.n38 VP.n37 0.189894
R121 VP.n38 VP.n19 0.189894
R122 VP.n42 VP.n19 0.189894
R123 VP.n43 VP.n42 0.189894
R124 VP.n44 VP.n43 0.189894
R125 VP.n44 VP.n17 0.189894
R126 VP.n49 VP.n17 0.189894
R127 VP.n50 VP.n49 0.189894
R128 VP.n51 VP.n50 0.189894
R129 VP.n51 VP.n15 0.189894
R130 VP.n55 VP.n15 0.189894
R131 VP.n61 VP.n13 0.189894
R132 VP.n62 VP.n61 0.189894
R133 VP.n63 VP.n62 0.189894
R134 VP.n63 VP.n11 0.189894
R135 VP.n67 VP.n11 0.189894
R136 VP.n68 VP.n67 0.189894
R137 VP.n68 VP.n9 0.189894
R138 VP.n72 VP.n9 0.189894
R139 VP.n73 VP.n72 0.189894
R140 VP.n74 VP.n73 0.189894
R141 VP.n74 VP.n7 0.189894
R142 VP.n78 VP.n7 0.189894
R143 VP.n79 VP.n78 0.189894
R144 VP.n80 VP.n79 0.189894
R145 VP.n80 VP.n5 0.189894
R146 VP.n84 VP.n5 0.189894
R147 VP.n85 VP.n84 0.189894
R148 VP.n86 VP.n85 0.189894
R149 VP.n86 VP.n3 0.189894
R150 VP.n91 VP.n3 0.189894
R151 VP.n92 VP.n91 0.189894
R152 VP.n93 VP.n92 0.189894
R153 VP.n93 VP.n1 0.189894
R154 VP.n97 VP.n1 0.189894
R155 VDD1.n84 VDD1.n0 289.615
R156 VDD1.n175 VDD1.n91 289.615
R157 VDD1.n85 VDD1.n84 185
R158 VDD1.n83 VDD1.n82 185
R159 VDD1.n4 VDD1.n3 185
R160 VDD1.n77 VDD1.n76 185
R161 VDD1.n75 VDD1.n6 185
R162 VDD1.n74 VDD1.n73 185
R163 VDD1.n9 VDD1.n7 185
R164 VDD1.n68 VDD1.n67 185
R165 VDD1.n66 VDD1.n65 185
R166 VDD1.n13 VDD1.n12 185
R167 VDD1.n60 VDD1.n59 185
R168 VDD1.n58 VDD1.n57 185
R169 VDD1.n17 VDD1.n16 185
R170 VDD1.n52 VDD1.n51 185
R171 VDD1.n50 VDD1.n49 185
R172 VDD1.n21 VDD1.n20 185
R173 VDD1.n44 VDD1.n43 185
R174 VDD1.n42 VDD1.n41 185
R175 VDD1.n25 VDD1.n24 185
R176 VDD1.n36 VDD1.n35 185
R177 VDD1.n34 VDD1.n33 185
R178 VDD1.n29 VDD1.n28 185
R179 VDD1.n119 VDD1.n118 185
R180 VDD1.n124 VDD1.n123 185
R181 VDD1.n126 VDD1.n125 185
R182 VDD1.n115 VDD1.n114 185
R183 VDD1.n132 VDD1.n131 185
R184 VDD1.n134 VDD1.n133 185
R185 VDD1.n111 VDD1.n110 185
R186 VDD1.n140 VDD1.n139 185
R187 VDD1.n142 VDD1.n141 185
R188 VDD1.n107 VDD1.n106 185
R189 VDD1.n148 VDD1.n147 185
R190 VDD1.n150 VDD1.n149 185
R191 VDD1.n103 VDD1.n102 185
R192 VDD1.n156 VDD1.n155 185
R193 VDD1.n158 VDD1.n157 185
R194 VDD1.n99 VDD1.n98 185
R195 VDD1.n165 VDD1.n164 185
R196 VDD1.n166 VDD1.n97 185
R197 VDD1.n168 VDD1.n167 185
R198 VDD1.n95 VDD1.n94 185
R199 VDD1.n174 VDD1.n173 185
R200 VDD1.n176 VDD1.n175 185
R201 VDD1.n30 VDD1.t7 147.659
R202 VDD1.n120 VDD1.t9 147.659
R203 VDD1.n84 VDD1.n83 104.615
R204 VDD1.n83 VDD1.n3 104.615
R205 VDD1.n76 VDD1.n3 104.615
R206 VDD1.n76 VDD1.n75 104.615
R207 VDD1.n75 VDD1.n74 104.615
R208 VDD1.n74 VDD1.n7 104.615
R209 VDD1.n67 VDD1.n7 104.615
R210 VDD1.n67 VDD1.n66 104.615
R211 VDD1.n66 VDD1.n12 104.615
R212 VDD1.n59 VDD1.n12 104.615
R213 VDD1.n59 VDD1.n58 104.615
R214 VDD1.n58 VDD1.n16 104.615
R215 VDD1.n51 VDD1.n16 104.615
R216 VDD1.n51 VDD1.n50 104.615
R217 VDD1.n50 VDD1.n20 104.615
R218 VDD1.n43 VDD1.n20 104.615
R219 VDD1.n43 VDD1.n42 104.615
R220 VDD1.n42 VDD1.n24 104.615
R221 VDD1.n35 VDD1.n24 104.615
R222 VDD1.n35 VDD1.n34 104.615
R223 VDD1.n34 VDD1.n28 104.615
R224 VDD1.n124 VDD1.n118 104.615
R225 VDD1.n125 VDD1.n124 104.615
R226 VDD1.n125 VDD1.n114 104.615
R227 VDD1.n132 VDD1.n114 104.615
R228 VDD1.n133 VDD1.n132 104.615
R229 VDD1.n133 VDD1.n110 104.615
R230 VDD1.n140 VDD1.n110 104.615
R231 VDD1.n141 VDD1.n140 104.615
R232 VDD1.n141 VDD1.n106 104.615
R233 VDD1.n148 VDD1.n106 104.615
R234 VDD1.n149 VDD1.n148 104.615
R235 VDD1.n149 VDD1.n102 104.615
R236 VDD1.n156 VDD1.n102 104.615
R237 VDD1.n157 VDD1.n156 104.615
R238 VDD1.n157 VDD1.n98 104.615
R239 VDD1.n165 VDD1.n98 104.615
R240 VDD1.n166 VDD1.n165 104.615
R241 VDD1.n167 VDD1.n166 104.615
R242 VDD1.n167 VDD1.n94 104.615
R243 VDD1.n174 VDD1.n94 104.615
R244 VDD1.n175 VDD1.n174 104.615
R245 VDD1.n183 VDD1.n182 65.3124
R246 VDD1.n90 VDD1.n89 63.2989
R247 VDD1.n185 VDD1.n184 63.2988
R248 VDD1.n181 VDD1.n180 63.2988
R249 VDD1.n90 VDD1.n88 54.144
R250 VDD1.n181 VDD1.n179 54.144
R251 VDD1.n185 VDD1.n183 52.7552
R252 VDD1.t7 VDD1.n28 52.3082
R253 VDD1.t9 VDD1.n118 52.3082
R254 VDD1.n30 VDD1.n29 15.6677
R255 VDD1.n120 VDD1.n119 15.6677
R256 VDD1.n77 VDD1.n6 13.1884
R257 VDD1.n168 VDD1.n97 13.1884
R258 VDD1.n78 VDD1.n4 12.8005
R259 VDD1.n73 VDD1.n8 12.8005
R260 VDD1.n33 VDD1.n32 12.8005
R261 VDD1.n123 VDD1.n122 12.8005
R262 VDD1.n164 VDD1.n163 12.8005
R263 VDD1.n169 VDD1.n95 12.8005
R264 VDD1.n82 VDD1.n81 12.0247
R265 VDD1.n72 VDD1.n9 12.0247
R266 VDD1.n36 VDD1.n27 12.0247
R267 VDD1.n126 VDD1.n117 12.0247
R268 VDD1.n162 VDD1.n99 12.0247
R269 VDD1.n173 VDD1.n172 12.0247
R270 VDD1.n85 VDD1.n2 11.249
R271 VDD1.n69 VDD1.n68 11.249
R272 VDD1.n37 VDD1.n25 11.249
R273 VDD1.n127 VDD1.n115 11.249
R274 VDD1.n159 VDD1.n158 11.249
R275 VDD1.n176 VDD1.n93 11.249
R276 VDD1.n86 VDD1.n0 10.4732
R277 VDD1.n65 VDD1.n11 10.4732
R278 VDD1.n41 VDD1.n40 10.4732
R279 VDD1.n131 VDD1.n130 10.4732
R280 VDD1.n155 VDD1.n101 10.4732
R281 VDD1.n177 VDD1.n91 10.4732
R282 VDD1.n64 VDD1.n13 9.69747
R283 VDD1.n44 VDD1.n23 9.69747
R284 VDD1.n134 VDD1.n113 9.69747
R285 VDD1.n154 VDD1.n103 9.69747
R286 VDD1.n88 VDD1.n87 9.45567
R287 VDD1.n179 VDD1.n178 9.45567
R288 VDD1.n56 VDD1.n55 9.3005
R289 VDD1.n15 VDD1.n14 9.3005
R290 VDD1.n62 VDD1.n61 9.3005
R291 VDD1.n64 VDD1.n63 9.3005
R292 VDD1.n11 VDD1.n10 9.3005
R293 VDD1.n70 VDD1.n69 9.3005
R294 VDD1.n72 VDD1.n71 9.3005
R295 VDD1.n8 VDD1.n5 9.3005
R296 VDD1.n87 VDD1.n86 9.3005
R297 VDD1.n2 VDD1.n1 9.3005
R298 VDD1.n81 VDD1.n80 9.3005
R299 VDD1.n79 VDD1.n78 9.3005
R300 VDD1.n54 VDD1.n53 9.3005
R301 VDD1.n19 VDD1.n18 9.3005
R302 VDD1.n48 VDD1.n47 9.3005
R303 VDD1.n46 VDD1.n45 9.3005
R304 VDD1.n23 VDD1.n22 9.3005
R305 VDD1.n40 VDD1.n39 9.3005
R306 VDD1.n38 VDD1.n37 9.3005
R307 VDD1.n27 VDD1.n26 9.3005
R308 VDD1.n32 VDD1.n31 9.3005
R309 VDD1.n178 VDD1.n177 9.3005
R310 VDD1.n93 VDD1.n92 9.3005
R311 VDD1.n172 VDD1.n171 9.3005
R312 VDD1.n170 VDD1.n169 9.3005
R313 VDD1.n109 VDD1.n108 9.3005
R314 VDD1.n138 VDD1.n137 9.3005
R315 VDD1.n136 VDD1.n135 9.3005
R316 VDD1.n113 VDD1.n112 9.3005
R317 VDD1.n130 VDD1.n129 9.3005
R318 VDD1.n128 VDD1.n127 9.3005
R319 VDD1.n117 VDD1.n116 9.3005
R320 VDD1.n122 VDD1.n121 9.3005
R321 VDD1.n144 VDD1.n143 9.3005
R322 VDD1.n146 VDD1.n145 9.3005
R323 VDD1.n105 VDD1.n104 9.3005
R324 VDD1.n152 VDD1.n151 9.3005
R325 VDD1.n154 VDD1.n153 9.3005
R326 VDD1.n101 VDD1.n100 9.3005
R327 VDD1.n160 VDD1.n159 9.3005
R328 VDD1.n162 VDD1.n161 9.3005
R329 VDD1.n163 VDD1.n96 9.3005
R330 VDD1.n61 VDD1.n60 8.92171
R331 VDD1.n45 VDD1.n21 8.92171
R332 VDD1.n135 VDD1.n111 8.92171
R333 VDD1.n151 VDD1.n150 8.92171
R334 VDD1.n57 VDD1.n15 8.14595
R335 VDD1.n49 VDD1.n48 8.14595
R336 VDD1.n139 VDD1.n138 8.14595
R337 VDD1.n147 VDD1.n105 8.14595
R338 VDD1.n56 VDD1.n17 7.3702
R339 VDD1.n52 VDD1.n19 7.3702
R340 VDD1.n142 VDD1.n109 7.3702
R341 VDD1.n146 VDD1.n107 7.3702
R342 VDD1.n53 VDD1.n17 6.59444
R343 VDD1.n53 VDD1.n52 6.59444
R344 VDD1.n143 VDD1.n142 6.59444
R345 VDD1.n143 VDD1.n107 6.59444
R346 VDD1.n57 VDD1.n56 5.81868
R347 VDD1.n49 VDD1.n19 5.81868
R348 VDD1.n139 VDD1.n109 5.81868
R349 VDD1.n147 VDD1.n146 5.81868
R350 VDD1.n60 VDD1.n15 5.04292
R351 VDD1.n48 VDD1.n21 5.04292
R352 VDD1.n138 VDD1.n111 5.04292
R353 VDD1.n150 VDD1.n105 5.04292
R354 VDD1.n31 VDD1.n30 4.38563
R355 VDD1.n121 VDD1.n120 4.38563
R356 VDD1.n61 VDD1.n13 4.26717
R357 VDD1.n45 VDD1.n44 4.26717
R358 VDD1.n135 VDD1.n134 4.26717
R359 VDD1.n151 VDD1.n103 4.26717
R360 VDD1.n88 VDD1.n0 3.49141
R361 VDD1.n65 VDD1.n64 3.49141
R362 VDD1.n41 VDD1.n23 3.49141
R363 VDD1.n131 VDD1.n113 3.49141
R364 VDD1.n155 VDD1.n154 3.49141
R365 VDD1.n179 VDD1.n91 3.49141
R366 VDD1.n86 VDD1.n85 2.71565
R367 VDD1.n68 VDD1.n11 2.71565
R368 VDD1.n40 VDD1.n25 2.71565
R369 VDD1.n130 VDD1.n115 2.71565
R370 VDD1.n158 VDD1.n101 2.71565
R371 VDD1.n177 VDD1.n176 2.71565
R372 VDD1 VDD1.n185 2.01128
R373 VDD1.n82 VDD1.n2 1.93989
R374 VDD1.n69 VDD1.n9 1.93989
R375 VDD1.n37 VDD1.n36 1.93989
R376 VDD1.n127 VDD1.n126 1.93989
R377 VDD1.n159 VDD1.n99 1.93989
R378 VDD1.n173 VDD1.n93 1.93989
R379 VDD1.n184 VDD1.t2 1.22197
R380 VDD1.n184 VDD1.t3 1.22197
R381 VDD1.n89 VDD1.t5 1.22197
R382 VDD1.n89 VDD1.t4 1.22197
R383 VDD1.n182 VDD1.t6 1.22197
R384 VDD1.n182 VDD1.t1 1.22197
R385 VDD1.n180 VDD1.t8 1.22197
R386 VDD1.n180 VDD1.t0 1.22197
R387 VDD1.n81 VDD1.n4 1.16414
R388 VDD1.n73 VDD1.n72 1.16414
R389 VDD1.n33 VDD1.n27 1.16414
R390 VDD1.n123 VDD1.n117 1.16414
R391 VDD1.n164 VDD1.n162 1.16414
R392 VDD1.n172 VDD1.n95 1.16414
R393 VDD1 VDD1.n90 0.748345
R394 VDD1.n183 VDD1.n181 0.634809
R395 VDD1.n78 VDD1.n77 0.388379
R396 VDD1.n8 VDD1.n6 0.388379
R397 VDD1.n32 VDD1.n29 0.388379
R398 VDD1.n122 VDD1.n119 0.388379
R399 VDD1.n163 VDD1.n97 0.388379
R400 VDD1.n169 VDD1.n168 0.388379
R401 VDD1.n87 VDD1.n1 0.155672
R402 VDD1.n80 VDD1.n1 0.155672
R403 VDD1.n80 VDD1.n79 0.155672
R404 VDD1.n79 VDD1.n5 0.155672
R405 VDD1.n71 VDD1.n5 0.155672
R406 VDD1.n71 VDD1.n70 0.155672
R407 VDD1.n70 VDD1.n10 0.155672
R408 VDD1.n63 VDD1.n10 0.155672
R409 VDD1.n63 VDD1.n62 0.155672
R410 VDD1.n62 VDD1.n14 0.155672
R411 VDD1.n55 VDD1.n14 0.155672
R412 VDD1.n55 VDD1.n54 0.155672
R413 VDD1.n54 VDD1.n18 0.155672
R414 VDD1.n47 VDD1.n18 0.155672
R415 VDD1.n47 VDD1.n46 0.155672
R416 VDD1.n46 VDD1.n22 0.155672
R417 VDD1.n39 VDD1.n22 0.155672
R418 VDD1.n39 VDD1.n38 0.155672
R419 VDD1.n38 VDD1.n26 0.155672
R420 VDD1.n31 VDD1.n26 0.155672
R421 VDD1.n121 VDD1.n116 0.155672
R422 VDD1.n128 VDD1.n116 0.155672
R423 VDD1.n129 VDD1.n128 0.155672
R424 VDD1.n129 VDD1.n112 0.155672
R425 VDD1.n136 VDD1.n112 0.155672
R426 VDD1.n137 VDD1.n136 0.155672
R427 VDD1.n137 VDD1.n108 0.155672
R428 VDD1.n144 VDD1.n108 0.155672
R429 VDD1.n145 VDD1.n144 0.155672
R430 VDD1.n145 VDD1.n104 0.155672
R431 VDD1.n152 VDD1.n104 0.155672
R432 VDD1.n153 VDD1.n152 0.155672
R433 VDD1.n153 VDD1.n100 0.155672
R434 VDD1.n160 VDD1.n100 0.155672
R435 VDD1.n161 VDD1.n160 0.155672
R436 VDD1.n161 VDD1.n96 0.155672
R437 VDD1.n170 VDD1.n96 0.155672
R438 VDD1.n171 VDD1.n170 0.155672
R439 VDD1.n171 VDD1.n92 0.155672
R440 VDD1.n178 VDD1.n92 0.155672
R441 VTAIL.n368 VTAIL.n284 289.615
R442 VTAIL.n86 VTAIL.n2 289.615
R443 VTAIL.n278 VTAIL.n194 289.615
R444 VTAIL.n184 VTAIL.n100 289.615
R445 VTAIL.n312 VTAIL.n311 185
R446 VTAIL.n317 VTAIL.n316 185
R447 VTAIL.n319 VTAIL.n318 185
R448 VTAIL.n308 VTAIL.n307 185
R449 VTAIL.n325 VTAIL.n324 185
R450 VTAIL.n327 VTAIL.n326 185
R451 VTAIL.n304 VTAIL.n303 185
R452 VTAIL.n333 VTAIL.n332 185
R453 VTAIL.n335 VTAIL.n334 185
R454 VTAIL.n300 VTAIL.n299 185
R455 VTAIL.n341 VTAIL.n340 185
R456 VTAIL.n343 VTAIL.n342 185
R457 VTAIL.n296 VTAIL.n295 185
R458 VTAIL.n349 VTAIL.n348 185
R459 VTAIL.n351 VTAIL.n350 185
R460 VTAIL.n292 VTAIL.n291 185
R461 VTAIL.n358 VTAIL.n357 185
R462 VTAIL.n359 VTAIL.n290 185
R463 VTAIL.n361 VTAIL.n360 185
R464 VTAIL.n288 VTAIL.n287 185
R465 VTAIL.n367 VTAIL.n366 185
R466 VTAIL.n369 VTAIL.n368 185
R467 VTAIL.n30 VTAIL.n29 185
R468 VTAIL.n35 VTAIL.n34 185
R469 VTAIL.n37 VTAIL.n36 185
R470 VTAIL.n26 VTAIL.n25 185
R471 VTAIL.n43 VTAIL.n42 185
R472 VTAIL.n45 VTAIL.n44 185
R473 VTAIL.n22 VTAIL.n21 185
R474 VTAIL.n51 VTAIL.n50 185
R475 VTAIL.n53 VTAIL.n52 185
R476 VTAIL.n18 VTAIL.n17 185
R477 VTAIL.n59 VTAIL.n58 185
R478 VTAIL.n61 VTAIL.n60 185
R479 VTAIL.n14 VTAIL.n13 185
R480 VTAIL.n67 VTAIL.n66 185
R481 VTAIL.n69 VTAIL.n68 185
R482 VTAIL.n10 VTAIL.n9 185
R483 VTAIL.n76 VTAIL.n75 185
R484 VTAIL.n77 VTAIL.n8 185
R485 VTAIL.n79 VTAIL.n78 185
R486 VTAIL.n6 VTAIL.n5 185
R487 VTAIL.n85 VTAIL.n84 185
R488 VTAIL.n87 VTAIL.n86 185
R489 VTAIL.n279 VTAIL.n278 185
R490 VTAIL.n277 VTAIL.n276 185
R491 VTAIL.n198 VTAIL.n197 185
R492 VTAIL.n271 VTAIL.n270 185
R493 VTAIL.n269 VTAIL.n200 185
R494 VTAIL.n268 VTAIL.n267 185
R495 VTAIL.n203 VTAIL.n201 185
R496 VTAIL.n262 VTAIL.n261 185
R497 VTAIL.n260 VTAIL.n259 185
R498 VTAIL.n207 VTAIL.n206 185
R499 VTAIL.n254 VTAIL.n253 185
R500 VTAIL.n252 VTAIL.n251 185
R501 VTAIL.n211 VTAIL.n210 185
R502 VTAIL.n246 VTAIL.n245 185
R503 VTAIL.n244 VTAIL.n243 185
R504 VTAIL.n215 VTAIL.n214 185
R505 VTAIL.n238 VTAIL.n237 185
R506 VTAIL.n236 VTAIL.n235 185
R507 VTAIL.n219 VTAIL.n218 185
R508 VTAIL.n230 VTAIL.n229 185
R509 VTAIL.n228 VTAIL.n227 185
R510 VTAIL.n223 VTAIL.n222 185
R511 VTAIL.n185 VTAIL.n184 185
R512 VTAIL.n183 VTAIL.n182 185
R513 VTAIL.n104 VTAIL.n103 185
R514 VTAIL.n177 VTAIL.n176 185
R515 VTAIL.n175 VTAIL.n106 185
R516 VTAIL.n174 VTAIL.n173 185
R517 VTAIL.n109 VTAIL.n107 185
R518 VTAIL.n168 VTAIL.n167 185
R519 VTAIL.n166 VTAIL.n165 185
R520 VTAIL.n113 VTAIL.n112 185
R521 VTAIL.n160 VTAIL.n159 185
R522 VTAIL.n158 VTAIL.n157 185
R523 VTAIL.n117 VTAIL.n116 185
R524 VTAIL.n152 VTAIL.n151 185
R525 VTAIL.n150 VTAIL.n149 185
R526 VTAIL.n121 VTAIL.n120 185
R527 VTAIL.n144 VTAIL.n143 185
R528 VTAIL.n142 VTAIL.n141 185
R529 VTAIL.n125 VTAIL.n124 185
R530 VTAIL.n136 VTAIL.n135 185
R531 VTAIL.n134 VTAIL.n133 185
R532 VTAIL.n129 VTAIL.n128 185
R533 VTAIL.n313 VTAIL.t3 147.659
R534 VTAIL.n31 VTAIL.t11 147.659
R535 VTAIL.n224 VTAIL.t13 147.659
R536 VTAIL.n130 VTAIL.t6 147.659
R537 VTAIL.n317 VTAIL.n311 104.615
R538 VTAIL.n318 VTAIL.n317 104.615
R539 VTAIL.n318 VTAIL.n307 104.615
R540 VTAIL.n325 VTAIL.n307 104.615
R541 VTAIL.n326 VTAIL.n325 104.615
R542 VTAIL.n326 VTAIL.n303 104.615
R543 VTAIL.n333 VTAIL.n303 104.615
R544 VTAIL.n334 VTAIL.n333 104.615
R545 VTAIL.n334 VTAIL.n299 104.615
R546 VTAIL.n341 VTAIL.n299 104.615
R547 VTAIL.n342 VTAIL.n341 104.615
R548 VTAIL.n342 VTAIL.n295 104.615
R549 VTAIL.n349 VTAIL.n295 104.615
R550 VTAIL.n350 VTAIL.n349 104.615
R551 VTAIL.n350 VTAIL.n291 104.615
R552 VTAIL.n358 VTAIL.n291 104.615
R553 VTAIL.n359 VTAIL.n358 104.615
R554 VTAIL.n360 VTAIL.n359 104.615
R555 VTAIL.n360 VTAIL.n287 104.615
R556 VTAIL.n367 VTAIL.n287 104.615
R557 VTAIL.n368 VTAIL.n367 104.615
R558 VTAIL.n35 VTAIL.n29 104.615
R559 VTAIL.n36 VTAIL.n35 104.615
R560 VTAIL.n36 VTAIL.n25 104.615
R561 VTAIL.n43 VTAIL.n25 104.615
R562 VTAIL.n44 VTAIL.n43 104.615
R563 VTAIL.n44 VTAIL.n21 104.615
R564 VTAIL.n51 VTAIL.n21 104.615
R565 VTAIL.n52 VTAIL.n51 104.615
R566 VTAIL.n52 VTAIL.n17 104.615
R567 VTAIL.n59 VTAIL.n17 104.615
R568 VTAIL.n60 VTAIL.n59 104.615
R569 VTAIL.n60 VTAIL.n13 104.615
R570 VTAIL.n67 VTAIL.n13 104.615
R571 VTAIL.n68 VTAIL.n67 104.615
R572 VTAIL.n68 VTAIL.n9 104.615
R573 VTAIL.n76 VTAIL.n9 104.615
R574 VTAIL.n77 VTAIL.n76 104.615
R575 VTAIL.n78 VTAIL.n77 104.615
R576 VTAIL.n78 VTAIL.n5 104.615
R577 VTAIL.n85 VTAIL.n5 104.615
R578 VTAIL.n86 VTAIL.n85 104.615
R579 VTAIL.n278 VTAIL.n277 104.615
R580 VTAIL.n277 VTAIL.n197 104.615
R581 VTAIL.n270 VTAIL.n197 104.615
R582 VTAIL.n270 VTAIL.n269 104.615
R583 VTAIL.n269 VTAIL.n268 104.615
R584 VTAIL.n268 VTAIL.n201 104.615
R585 VTAIL.n261 VTAIL.n201 104.615
R586 VTAIL.n261 VTAIL.n260 104.615
R587 VTAIL.n260 VTAIL.n206 104.615
R588 VTAIL.n253 VTAIL.n206 104.615
R589 VTAIL.n253 VTAIL.n252 104.615
R590 VTAIL.n252 VTAIL.n210 104.615
R591 VTAIL.n245 VTAIL.n210 104.615
R592 VTAIL.n245 VTAIL.n244 104.615
R593 VTAIL.n244 VTAIL.n214 104.615
R594 VTAIL.n237 VTAIL.n214 104.615
R595 VTAIL.n237 VTAIL.n236 104.615
R596 VTAIL.n236 VTAIL.n218 104.615
R597 VTAIL.n229 VTAIL.n218 104.615
R598 VTAIL.n229 VTAIL.n228 104.615
R599 VTAIL.n228 VTAIL.n222 104.615
R600 VTAIL.n184 VTAIL.n183 104.615
R601 VTAIL.n183 VTAIL.n103 104.615
R602 VTAIL.n176 VTAIL.n103 104.615
R603 VTAIL.n176 VTAIL.n175 104.615
R604 VTAIL.n175 VTAIL.n174 104.615
R605 VTAIL.n174 VTAIL.n107 104.615
R606 VTAIL.n167 VTAIL.n107 104.615
R607 VTAIL.n167 VTAIL.n166 104.615
R608 VTAIL.n166 VTAIL.n112 104.615
R609 VTAIL.n159 VTAIL.n112 104.615
R610 VTAIL.n159 VTAIL.n158 104.615
R611 VTAIL.n158 VTAIL.n116 104.615
R612 VTAIL.n151 VTAIL.n116 104.615
R613 VTAIL.n151 VTAIL.n150 104.615
R614 VTAIL.n150 VTAIL.n120 104.615
R615 VTAIL.n143 VTAIL.n120 104.615
R616 VTAIL.n143 VTAIL.n142 104.615
R617 VTAIL.n142 VTAIL.n124 104.615
R618 VTAIL.n135 VTAIL.n124 104.615
R619 VTAIL.n135 VTAIL.n134 104.615
R620 VTAIL.n134 VTAIL.n128 104.615
R621 VTAIL.t3 VTAIL.n311 52.3082
R622 VTAIL.t11 VTAIL.n29 52.3082
R623 VTAIL.t13 VTAIL.n222 52.3082
R624 VTAIL.t6 VTAIL.n128 52.3082
R625 VTAIL.n193 VTAIL.n192 46.6202
R626 VTAIL.n191 VTAIL.n190 46.6202
R627 VTAIL.n99 VTAIL.n98 46.6202
R628 VTAIL.n97 VTAIL.n96 46.6202
R629 VTAIL.n375 VTAIL.n374 46.62
R630 VTAIL.n1 VTAIL.n0 46.62
R631 VTAIL.n93 VTAIL.n92 46.62
R632 VTAIL.n95 VTAIL.n94 46.62
R633 VTAIL.n373 VTAIL.n372 34.7066
R634 VTAIL.n91 VTAIL.n90 34.7066
R635 VTAIL.n283 VTAIL.n282 34.7066
R636 VTAIL.n189 VTAIL.n188 34.7066
R637 VTAIL.n97 VTAIL.n95 31.8583
R638 VTAIL.n373 VTAIL.n283 29.0996
R639 VTAIL.n313 VTAIL.n312 15.6677
R640 VTAIL.n31 VTAIL.n30 15.6677
R641 VTAIL.n224 VTAIL.n223 15.6677
R642 VTAIL.n130 VTAIL.n129 15.6677
R643 VTAIL.n361 VTAIL.n290 13.1884
R644 VTAIL.n79 VTAIL.n8 13.1884
R645 VTAIL.n271 VTAIL.n200 13.1884
R646 VTAIL.n177 VTAIL.n106 13.1884
R647 VTAIL.n316 VTAIL.n315 12.8005
R648 VTAIL.n357 VTAIL.n356 12.8005
R649 VTAIL.n362 VTAIL.n288 12.8005
R650 VTAIL.n34 VTAIL.n33 12.8005
R651 VTAIL.n75 VTAIL.n74 12.8005
R652 VTAIL.n80 VTAIL.n6 12.8005
R653 VTAIL.n272 VTAIL.n198 12.8005
R654 VTAIL.n267 VTAIL.n202 12.8005
R655 VTAIL.n227 VTAIL.n226 12.8005
R656 VTAIL.n178 VTAIL.n104 12.8005
R657 VTAIL.n173 VTAIL.n108 12.8005
R658 VTAIL.n133 VTAIL.n132 12.8005
R659 VTAIL.n319 VTAIL.n310 12.0247
R660 VTAIL.n355 VTAIL.n292 12.0247
R661 VTAIL.n366 VTAIL.n365 12.0247
R662 VTAIL.n37 VTAIL.n28 12.0247
R663 VTAIL.n73 VTAIL.n10 12.0247
R664 VTAIL.n84 VTAIL.n83 12.0247
R665 VTAIL.n276 VTAIL.n275 12.0247
R666 VTAIL.n266 VTAIL.n203 12.0247
R667 VTAIL.n230 VTAIL.n221 12.0247
R668 VTAIL.n182 VTAIL.n181 12.0247
R669 VTAIL.n172 VTAIL.n109 12.0247
R670 VTAIL.n136 VTAIL.n127 12.0247
R671 VTAIL.n320 VTAIL.n308 11.249
R672 VTAIL.n352 VTAIL.n351 11.249
R673 VTAIL.n369 VTAIL.n286 11.249
R674 VTAIL.n38 VTAIL.n26 11.249
R675 VTAIL.n70 VTAIL.n69 11.249
R676 VTAIL.n87 VTAIL.n4 11.249
R677 VTAIL.n279 VTAIL.n196 11.249
R678 VTAIL.n263 VTAIL.n262 11.249
R679 VTAIL.n231 VTAIL.n219 11.249
R680 VTAIL.n185 VTAIL.n102 11.249
R681 VTAIL.n169 VTAIL.n168 11.249
R682 VTAIL.n137 VTAIL.n125 11.249
R683 VTAIL.n324 VTAIL.n323 10.4732
R684 VTAIL.n348 VTAIL.n294 10.4732
R685 VTAIL.n370 VTAIL.n284 10.4732
R686 VTAIL.n42 VTAIL.n41 10.4732
R687 VTAIL.n66 VTAIL.n12 10.4732
R688 VTAIL.n88 VTAIL.n2 10.4732
R689 VTAIL.n280 VTAIL.n194 10.4732
R690 VTAIL.n259 VTAIL.n205 10.4732
R691 VTAIL.n235 VTAIL.n234 10.4732
R692 VTAIL.n186 VTAIL.n100 10.4732
R693 VTAIL.n165 VTAIL.n111 10.4732
R694 VTAIL.n141 VTAIL.n140 10.4732
R695 VTAIL.n327 VTAIL.n306 9.69747
R696 VTAIL.n347 VTAIL.n296 9.69747
R697 VTAIL.n45 VTAIL.n24 9.69747
R698 VTAIL.n65 VTAIL.n14 9.69747
R699 VTAIL.n258 VTAIL.n207 9.69747
R700 VTAIL.n238 VTAIL.n217 9.69747
R701 VTAIL.n164 VTAIL.n113 9.69747
R702 VTAIL.n144 VTAIL.n123 9.69747
R703 VTAIL.n372 VTAIL.n371 9.45567
R704 VTAIL.n90 VTAIL.n89 9.45567
R705 VTAIL.n282 VTAIL.n281 9.45567
R706 VTAIL.n188 VTAIL.n187 9.45567
R707 VTAIL.n371 VTAIL.n370 9.3005
R708 VTAIL.n286 VTAIL.n285 9.3005
R709 VTAIL.n365 VTAIL.n364 9.3005
R710 VTAIL.n363 VTAIL.n362 9.3005
R711 VTAIL.n302 VTAIL.n301 9.3005
R712 VTAIL.n331 VTAIL.n330 9.3005
R713 VTAIL.n329 VTAIL.n328 9.3005
R714 VTAIL.n306 VTAIL.n305 9.3005
R715 VTAIL.n323 VTAIL.n322 9.3005
R716 VTAIL.n321 VTAIL.n320 9.3005
R717 VTAIL.n310 VTAIL.n309 9.3005
R718 VTAIL.n315 VTAIL.n314 9.3005
R719 VTAIL.n337 VTAIL.n336 9.3005
R720 VTAIL.n339 VTAIL.n338 9.3005
R721 VTAIL.n298 VTAIL.n297 9.3005
R722 VTAIL.n345 VTAIL.n344 9.3005
R723 VTAIL.n347 VTAIL.n346 9.3005
R724 VTAIL.n294 VTAIL.n293 9.3005
R725 VTAIL.n353 VTAIL.n352 9.3005
R726 VTAIL.n355 VTAIL.n354 9.3005
R727 VTAIL.n356 VTAIL.n289 9.3005
R728 VTAIL.n89 VTAIL.n88 9.3005
R729 VTAIL.n4 VTAIL.n3 9.3005
R730 VTAIL.n83 VTAIL.n82 9.3005
R731 VTAIL.n81 VTAIL.n80 9.3005
R732 VTAIL.n20 VTAIL.n19 9.3005
R733 VTAIL.n49 VTAIL.n48 9.3005
R734 VTAIL.n47 VTAIL.n46 9.3005
R735 VTAIL.n24 VTAIL.n23 9.3005
R736 VTAIL.n41 VTAIL.n40 9.3005
R737 VTAIL.n39 VTAIL.n38 9.3005
R738 VTAIL.n28 VTAIL.n27 9.3005
R739 VTAIL.n33 VTAIL.n32 9.3005
R740 VTAIL.n55 VTAIL.n54 9.3005
R741 VTAIL.n57 VTAIL.n56 9.3005
R742 VTAIL.n16 VTAIL.n15 9.3005
R743 VTAIL.n63 VTAIL.n62 9.3005
R744 VTAIL.n65 VTAIL.n64 9.3005
R745 VTAIL.n12 VTAIL.n11 9.3005
R746 VTAIL.n71 VTAIL.n70 9.3005
R747 VTAIL.n73 VTAIL.n72 9.3005
R748 VTAIL.n74 VTAIL.n7 9.3005
R749 VTAIL.n250 VTAIL.n249 9.3005
R750 VTAIL.n209 VTAIL.n208 9.3005
R751 VTAIL.n256 VTAIL.n255 9.3005
R752 VTAIL.n258 VTAIL.n257 9.3005
R753 VTAIL.n205 VTAIL.n204 9.3005
R754 VTAIL.n264 VTAIL.n263 9.3005
R755 VTAIL.n266 VTAIL.n265 9.3005
R756 VTAIL.n202 VTAIL.n199 9.3005
R757 VTAIL.n281 VTAIL.n280 9.3005
R758 VTAIL.n196 VTAIL.n195 9.3005
R759 VTAIL.n275 VTAIL.n274 9.3005
R760 VTAIL.n273 VTAIL.n272 9.3005
R761 VTAIL.n248 VTAIL.n247 9.3005
R762 VTAIL.n213 VTAIL.n212 9.3005
R763 VTAIL.n242 VTAIL.n241 9.3005
R764 VTAIL.n240 VTAIL.n239 9.3005
R765 VTAIL.n217 VTAIL.n216 9.3005
R766 VTAIL.n234 VTAIL.n233 9.3005
R767 VTAIL.n232 VTAIL.n231 9.3005
R768 VTAIL.n221 VTAIL.n220 9.3005
R769 VTAIL.n226 VTAIL.n225 9.3005
R770 VTAIL.n156 VTAIL.n155 9.3005
R771 VTAIL.n115 VTAIL.n114 9.3005
R772 VTAIL.n162 VTAIL.n161 9.3005
R773 VTAIL.n164 VTAIL.n163 9.3005
R774 VTAIL.n111 VTAIL.n110 9.3005
R775 VTAIL.n170 VTAIL.n169 9.3005
R776 VTAIL.n172 VTAIL.n171 9.3005
R777 VTAIL.n108 VTAIL.n105 9.3005
R778 VTAIL.n187 VTAIL.n186 9.3005
R779 VTAIL.n102 VTAIL.n101 9.3005
R780 VTAIL.n181 VTAIL.n180 9.3005
R781 VTAIL.n179 VTAIL.n178 9.3005
R782 VTAIL.n154 VTAIL.n153 9.3005
R783 VTAIL.n119 VTAIL.n118 9.3005
R784 VTAIL.n148 VTAIL.n147 9.3005
R785 VTAIL.n146 VTAIL.n145 9.3005
R786 VTAIL.n123 VTAIL.n122 9.3005
R787 VTAIL.n140 VTAIL.n139 9.3005
R788 VTAIL.n138 VTAIL.n137 9.3005
R789 VTAIL.n127 VTAIL.n126 9.3005
R790 VTAIL.n132 VTAIL.n131 9.3005
R791 VTAIL.n328 VTAIL.n304 8.92171
R792 VTAIL.n344 VTAIL.n343 8.92171
R793 VTAIL.n46 VTAIL.n22 8.92171
R794 VTAIL.n62 VTAIL.n61 8.92171
R795 VTAIL.n255 VTAIL.n254 8.92171
R796 VTAIL.n239 VTAIL.n215 8.92171
R797 VTAIL.n161 VTAIL.n160 8.92171
R798 VTAIL.n145 VTAIL.n121 8.92171
R799 VTAIL.n332 VTAIL.n331 8.14595
R800 VTAIL.n340 VTAIL.n298 8.14595
R801 VTAIL.n50 VTAIL.n49 8.14595
R802 VTAIL.n58 VTAIL.n16 8.14595
R803 VTAIL.n251 VTAIL.n209 8.14595
R804 VTAIL.n243 VTAIL.n242 8.14595
R805 VTAIL.n157 VTAIL.n115 8.14595
R806 VTAIL.n149 VTAIL.n148 8.14595
R807 VTAIL.n335 VTAIL.n302 7.3702
R808 VTAIL.n339 VTAIL.n300 7.3702
R809 VTAIL.n53 VTAIL.n20 7.3702
R810 VTAIL.n57 VTAIL.n18 7.3702
R811 VTAIL.n250 VTAIL.n211 7.3702
R812 VTAIL.n246 VTAIL.n213 7.3702
R813 VTAIL.n156 VTAIL.n117 7.3702
R814 VTAIL.n152 VTAIL.n119 7.3702
R815 VTAIL.n336 VTAIL.n335 6.59444
R816 VTAIL.n336 VTAIL.n300 6.59444
R817 VTAIL.n54 VTAIL.n53 6.59444
R818 VTAIL.n54 VTAIL.n18 6.59444
R819 VTAIL.n247 VTAIL.n211 6.59444
R820 VTAIL.n247 VTAIL.n246 6.59444
R821 VTAIL.n153 VTAIL.n117 6.59444
R822 VTAIL.n153 VTAIL.n152 6.59444
R823 VTAIL.n332 VTAIL.n302 5.81868
R824 VTAIL.n340 VTAIL.n339 5.81868
R825 VTAIL.n50 VTAIL.n20 5.81868
R826 VTAIL.n58 VTAIL.n57 5.81868
R827 VTAIL.n251 VTAIL.n250 5.81868
R828 VTAIL.n243 VTAIL.n213 5.81868
R829 VTAIL.n157 VTAIL.n156 5.81868
R830 VTAIL.n149 VTAIL.n119 5.81868
R831 VTAIL.n331 VTAIL.n304 5.04292
R832 VTAIL.n343 VTAIL.n298 5.04292
R833 VTAIL.n49 VTAIL.n22 5.04292
R834 VTAIL.n61 VTAIL.n16 5.04292
R835 VTAIL.n254 VTAIL.n209 5.04292
R836 VTAIL.n242 VTAIL.n215 5.04292
R837 VTAIL.n160 VTAIL.n115 5.04292
R838 VTAIL.n148 VTAIL.n121 5.04292
R839 VTAIL.n314 VTAIL.n313 4.38563
R840 VTAIL.n32 VTAIL.n31 4.38563
R841 VTAIL.n225 VTAIL.n224 4.38563
R842 VTAIL.n131 VTAIL.n130 4.38563
R843 VTAIL.n328 VTAIL.n327 4.26717
R844 VTAIL.n344 VTAIL.n296 4.26717
R845 VTAIL.n46 VTAIL.n45 4.26717
R846 VTAIL.n62 VTAIL.n14 4.26717
R847 VTAIL.n255 VTAIL.n207 4.26717
R848 VTAIL.n239 VTAIL.n238 4.26717
R849 VTAIL.n161 VTAIL.n113 4.26717
R850 VTAIL.n145 VTAIL.n144 4.26717
R851 VTAIL.n324 VTAIL.n306 3.49141
R852 VTAIL.n348 VTAIL.n347 3.49141
R853 VTAIL.n372 VTAIL.n284 3.49141
R854 VTAIL.n42 VTAIL.n24 3.49141
R855 VTAIL.n66 VTAIL.n65 3.49141
R856 VTAIL.n90 VTAIL.n2 3.49141
R857 VTAIL.n282 VTAIL.n194 3.49141
R858 VTAIL.n259 VTAIL.n258 3.49141
R859 VTAIL.n235 VTAIL.n217 3.49141
R860 VTAIL.n188 VTAIL.n100 3.49141
R861 VTAIL.n165 VTAIL.n164 3.49141
R862 VTAIL.n141 VTAIL.n123 3.49141
R863 VTAIL.n99 VTAIL.n97 2.75912
R864 VTAIL.n189 VTAIL.n99 2.75912
R865 VTAIL.n193 VTAIL.n191 2.75912
R866 VTAIL.n283 VTAIL.n193 2.75912
R867 VTAIL.n95 VTAIL.n93 2.75912
R868 VTAIL.n93 VTAIL.n91 2.75912
R869 VTAIL.n375 VTAIL.n373 2.75912
R870 VTAIL.n323 VTAIL.n308 2.71565
R871 VTAIL.n351 VTAIL.n294 2.71565
R872 VTAIL.n370 VTAIL.n369 2.71565
R873 VTAIL.n41 VTAIL.n26 2.71565
R874 VTAIL.n69 VTAIL.n12 2.71565
R875 VTAIL.n88 VTAIL.n87 2.71565
R876 VTAIL.n280 VTAIL.n279 2.71565
R877 VTAIL.n262 VTAIL.n205 2.71565
R878 VTAIL.n234 VTAIL.n219 2.71565
R879 VTAIL.n186 VTAIL.n185 2.71565
R880 VTAIL.n168 VTAIL.n111 2.71565
R881 VTAIL.n140 VTAIL.n125 2.71565
R882 VTAIL VTAIL.n1 2.12766
R883 VTAIL.n320 VTAIL.n319 1.93989
R884 VTAIL.n352 VTAIL.n292 1.93989
R885 VTAIL.n366 VTAIL.n286 1.93989
R886 VTAIL.n38 VTAIL.n37 1.93989
R887 VTAIL.n70 VTAIL.n10 1.93989
R888 VTAIL.n84 VTAIL.n4 1.93989
R889 VTAIL.n276 VTAIL.n196 1.93989
R890 VTAIL.n263 VTAIL.n203 1.93989
R891 VTAIL.n231 VTAIL.n230 1.93989
R892 VTAIL.n182 VTAIL.n102 1.93989
R893 VTAIL.n169 VTAIL.n109 1.93989
R894 VTAIL.n137 VTAIL.n136 1.93989
R895 VTAIL.n191 VTAIL.n189 1.84964
R896 VTAIL.n91 VTAIL.n1 1.84964
R897 VTAIL.n374 VTAIL.t5 1.22197
R898 VTAIL.n374 VTAIL.t2 1.22197
R899 VTAIL.n0 VTAIL.t7 1.22197
R900 VTAIL.n0 VTAIL.t4 1.22197
R901 VTAIL.n92 VTAIL.t10 1.22197
R902 VTAIL.n92 VTAIL.t18 1.22197
R903 VTAIL.n94 VTAIL.t9 1.22197
R904 VTAIL.n94 VTAIL.t17 1.22197
R905 VTAIL.n192 VTAIL.t14 1.22197
R906 VTAIL.n192 VTAIL.t12 1.22197
R907 VTAIL.n190 VTAIL.t16 1.22197
R908 VTAIL.n190 VTAIL.t15 1.22197
R909 VTAIL.n98 VTAIL.t1 1.22197
R910 VTAIL.n98 VTAIL.t19 1.22197
R911 VTAIL.n96 VTAIL.t8 1.22197
R912 VTAIL.n96 VTAIL.t0 1.22197
R913 VTAIL.n316 VTAIL.n310 1.16414
R914 VTAIL.n357 VTAIL.n355 1.16414
R915 VTAIL.n365 VTAIL.n288 1.16414
R916 VTAIL.n34 VTAIL.n28 1.16414
R917 VTAIL.n75 VTAIL.n73 1.16414
R918 VTAIL.n83 VTAIL.n6 1.16414
R919 VTAIL.n275 VTAIL.n198 1.16414
R920 VTAIL.n267 VTAIL.n266 1.16414
R921 VTAIL.n227 VTAIL.n221 1.16414
R922 VTAIL.n181 VTAIL.n104 1.16414
R923 VTAIL.n173 VTAIL.n172 1.16414
R924 VTAIL.n133 VTAIL.n127 1.16414
R925 VTAIL VTAIL.n375 0.631965
R926 VTAIL.n315 VTAIL.n312 0.388379
R927 VTAIL.n356 VTAIL.n290 0.388379
R928 VTAIL.n362 VTAIL.n361 0.388379
R929 VTAIL.n33 VTAIL.n30 0.388379
R930 VTAIL.n74 VTAIL.n8 0.388379
R931 VTAIL.n80 VTAIL.n79 0.388379
R932 VTAIL.n272 VTAIL.n271 0.388379
R933 VTAIL.n202 VTAIL.n200 0.388379
R934 VTAIL.n226 VTAIL.n223 0.388379
R935 VTAIL.n178 VTAIL.n177 0.388379
R936 VTAIL.n108 VTAIL.n106 0.388379
R937 VTAIL.n132 VTAIL.n129 0.388379
R938 VTAIL.n314 VTAIL.n309 0.155672
R939 VTAIL.n321 VTAIL.n309 0.155672
R940 VTAIL.n322 VTAIL.n321 0.155672
R941 VTAIL.n322 VTAIL.n305 0.155672
R942 VTAIL.n329 VTAIL.n305 0.155672
R943 VTAIL.n330 VTAIL.n329 0.155672
R944 VTAIL.n330 VTAIL.n301 0.155672
R945 VTAIL.n337 VTAIL.n301 0.155672
R946 VTAIL.n338 VTAIL.n337 0.155672
R947 VTAIL.n338 VTAIL.n297 0.155672
R948 VTAIL.n345 VTAIL.n297 0.155672
R949 VTAIL.n346 VTAIL.n345 0.155672
R950 VTAIL.n346 VTAIL.n293 0.155672
R951 VTAIL.n353 VTAIL.n293 0.155672
R952 VTAIL.n354 VTAIL.n353 0.155672
R953 VTAIL.n354 VTAIL.n289 0.155672
R954 VTAIL.n363 VTAIL.n289 0.155672
R955 VTAIL.n364 VTAIL.n363 0.155672
R956 VTAIL.n364 VTAIL.n285 0.155672
R957 VTAIL.n371 VTAIL.n285 0.155672
R958 VTAIL.n32 VTAIL.n27 0.155672
R959 VTAIL.n39 VTAIL.n27 0.155672
R960 VTAIL.n40 VTAIL.n39 0.155672
R961 VTAIL.n40 VTAIL.n23 0.155672
R962 VTAIL.n47 VTAIL.n23 0.155672
R963 VTAIL.n48 VTAIL.n47 0.155672
R964 VTAIL.n48 VTAIL.n19 0.155672
R965 VTAIL.n55 VTAIL.n19 0.155672
R966 VTAIL.n56 VTAIL.n55 0.155672
R967 VTAIL.n56 VTAIL.n15 0.155672
R968 VTAIL.n63 VTAIL.n15 0.155672
R969 VTAIL.n64 VTAIL.n63 0.155672
R970 VTAIL.n64 VTAIL.n11 0.155672
R971 VTAIL.n71 VTAIL.n11 0.155672
R972 VTAIL.n72 VTAIL.n71 0.155672
R973 VTAIL.n72 VTAIL.n7 0.155672
R974 VTAIL.n81 VTAIL.n7 0.155672
R975 VTAIL.n82 VTAIL.n81 0.155672
R976 VTAIL.n82 VTAIL.n3 0.155672
R977 VTAIL.n89 VTAIL.n3 0.155672
R978 VTAIL.n281 VTAIL.n195 0.155672
R979 VTAIL.n274 VTAIL.n195 0.155672
R980 VTAIL.n274 VTAIL.n273 0.155672
R981 VTAIL.n273 VTAIL.n199 0.155672
R982 VTAIL.n265 VTAIL.n199 0.155672
R983 VTAIL.n265 VTAIL.n264 0.155672
R984 VTAIL.n264 VTAIL.n204 0.155672
R985 VTAIL.n257 VTAIL.n204 0.155672
R986 VTAIL.n257 VTAIL.n256 0.155672
R987 VTAIL.n256 VTAIL.n208 0.155672
R988 VTAIL.n249 VTAIL.n208 0.155672
R989 VTAIL.n249 VTAIL.n248 0.155672
R990 VTAIL.n248 VTAIL.n212 0.155672
R991 VTAIL.n241 VTAIL.n212 0.155672
R992 VTAIL.n241 VTAIL.n240 0.155672
R993 VTAIL.n240 VTAIL.n216 0.155672
R994 VTAIL.n233 VTAIL.n216 0.155672
R995 VTAIL.n233 VTAIL.n232 0.155672
R996 VTAIL.n232 VTAIL.n220 0.155672
R997 VTAIL.n225 VTAIL.n220 0.155672
R998 VTAIL.n187 VTAIL.n101 0.155672
R999 VTAIL.n180 VTAIL.n101 0.155672
R1000 VTAIL.n180 VTAIL.n179 0.155672
R1001 VTAIL.n179 VTAIL.n105 0.155672
R1002 VTAIL.n171 VTAIL.n105 0.155672
R1003 VTAIL.n171 VTAIL.n170 0.155672
R1004 VTAIL.n170 VTAIL.n110 0.155672
R1005 VTAIL.n163 VTAIL.n110 0.155672
R1006 VTAIL.n163 VTAIL.n162 0.155672
R1007 VTAIL.n162 VTAIL.n114 0.155672
R1008 VTAIL.n155 VTAIL.n114 0.155672
R1009 VTAIL.n155 VTAIL.n154 0.155672
R1010 VTAIL.n154 VTAIL.n118 0.155672
R1011 VTAIL.n147 VTAIL.n118 0.155672
R1012 VTAIL.n147 VTAIL.n146 0.155672
R1013 VTAIL.n146 VTAIL.n122 0.155672
R1014 VTAIL.n139 VTAIL.n122 0.155672
R1015 VTAIL.n139 VTAIL.n138 0.155672
R1016 VTAIL.n138 VTAIL.n126 0.155672
R1017 VTAIL.n131 VTAIL.n126 0.155672
R1018 B.n1117 B.n1116 585
R1019 B.n414 B.n177 585
R1020 B.n413 B.n412 585
R1021 B.n411 B.n410 585
R1022 B.n409 B.n408 585
R1023 B.n407 B.n406 585
R1024 B.n405 B.n404 585
R1025 B.n403 B.n402 585
R1026 B.n401 B.n400 585
R1027 B.n399 B.n398 585
R1028 B.n397 B.n396 585
R1029 B.n395 B.n394 585
R1030 B.n393 B.n392 585
R1031 B.n391 B.n390 585
R1032 B.n389 B.n388 585
R1033 B.n387 B.n386 585
R1034 B.n385 B.n384 585
R1035 B.n383 B.n382 585
R1036 B.n381 B.n380 585
R1037 B.n379 B.n378 585
R1038 B.n377 B.n376 585
R1039 B.n375 B.n374 585
R1040 B.n373 B.n372 585
R1041 B.n371 B.n370 585
R1042 B.n369 B.n368 585
R1043 B.n367 B.n366 585
R1044 B.n365 B.n364 585
R1045 B.n363 B.n362 585
R1046 B.n361 B.n360 585
R1047 B.n359 B.n358 585
R1048 B.n357 B.n356 585
R1049 B.n355 B.n354 585
R1050 B.n353 B.n352 585
R1051 B.n351 B.n350 585
R1052 B.n349 B.n348 585
R1053 B.n347 B.n346 585
R1054 B.n345 B.n344 585
R1055 B.n343 B.n342 585
R1056 B.n341 B.n340 585
R1057 B.n339 B.n338 585
R1058 B.n337 B.n336 585
R1059 B.n335 B.n334 585
R1060 B.n333 B.n332 585
R1061 B.n331 B.n330 585
R1062 B.n329 B.n328 585
R1063 B.n327 B.n326 585
R1064 B.n325 B.n324 585
R1065 B.n323 B.n322 585
R1066 B.n321 B.n320 585
R1067 B.n319 B.n318 585
R1068 B.n317 B.n316 585
R1069 B.n315 B.n314 585
R1070 B.n313 B.n312 585
R1071 B.n311 B.n310 585
R1072 B.n309 B.n308 585
R1073 B.n307 B.n306 585
R1074 B.n305 B.n304 585
R1075 B.n303 B.n302 585
R1076 B.n301 B.n300 585
R1077 B.n299 B.n298 585
R1078 B.n297 B.n296 585
R1079 B.n295 B.n294 585
R1080 B.n293 B.n292 585
R1081 B.n291 B.n290 585
R1082 B.n289 B.n288 585
R1083 B.n287 B.n286 585
R1084 B.n285 B.n284 585
R1085 B.n283 B.n282 585
R1086 B.n281 B.n280 585
R1087 B.n279 B.n278 585
R1088 B.n277 B.n276 585
R1089 B.n275 B.n274 585
R1090 B.n273 B.n272 585
R1091 B.n271 B.n270 585
R1092 B.n269 B.n268 585
R1093 B.n267 B.n266 585
R1094 B.n265 B.n264 585
R1095 B.n263 B.n262 585
R1096 B.n261 B.n260 585
R1097 B.n259 B.n258 585
R1098 B.n257 B.n256 585
R1099 B.n255 B.n254 585
R1100 B.n253 B.n252 585
R1101 B.n251 B.n250 585
R1102 B.n249 B.n248 585
R1103 B.n247 B.n246 585
R1104 B.n245 B.n244 585
R1105 B.n243 B.n242 585
R1106 B.n241 B.n240 585
R1107 B.n239 B.n238 585
R1108 B.n237 B.n236 585
R1109 B.n235 B.n234 585
R1110 B.n233 B.n232 585
R1111 B.n231 B.n230 585
R1112 B.n229 B.n228 585
R1113 B.n227 B.n226 585
R1114 B.n225 B.n224 585
R1115 B.n223 B.n222 585
R1116 B.n221 B.n220 585
R1117 B.n219 B.n218 585
R1118 B.n217 B.n216 585
R1119 B.n215 B.n214 585
R1120 B.n213 B.n212 585
R1121 B.n211 B.n210 585
R1122 B.n209 B.n208 585
R1123 B.n207 B.n206 585
R1124 B.n205 B.n204 585
R1125 B.n203 B.n202 585
R1126 B.n201 B.n200 585
R1127 B.n199 B.n198 585
R1128 B.n197 B.n196 585
R1129 B.n195 B.n194 585
R1130 B.n193 B.n192 585
R1131 B.n191 B.n190 585
R1132 B.n189 B.n188 585
R1133 B.n187 B.n186 585
R1134 B.n185 B.n184 585
R1135 B.n117 B.n116 585
R1136 B.n1115 B.n118 585
R1137 B.n1120 B.n118 585
R1138 B.n1114 B.n1113 585
R1139 B.n1113 B.n114 585
R1140 B.n1112 B.n113 585
R1141 B.n1126 B.n113 585
R1142 B.n1111 B.n112 585
R1143 B.n1127 B.n112 585
R1144 B.n1110 B.n111 585
R1145 B.n1128 B.n111 585
R1146 B.n1109 B.n1108 585
R1147 B.n1108 B.n107 585
R1148 B.n1107 B.n106 585
R1149 B.n1134 B.n106 585
R1150 B.n1106 B.n105 585
R1151 B.n1135 B.n105 585
R1152 B.n1105 B.n104 585
R1153 B.n1136 B.n104 585
R1154 B.n1104 B.n1103 585
R1155 B.n1103 B.n100 585
R1156 B.n1102 B.n99 585
R1157 B.n1142 B.n99 585
R1158 B.n1101 B.n98 585
R1159 B.n1143 B.n98 585
R1160 B.n1100 B.n97 585
R1161 B.n1144 B.n97 585
R1162 B.n1099 B.n1098 585
R1163 B.n1098 B.n93 585
R1164 B.n1097 B.n92 585
R1165 B.n1150 B.n92 585
R1166 B.n1096 B.n91 585
R1167 B.n1151 B.n91 585
R1168 B.n1095 B.n90 585
R1169 B.n1152 B.n90 585
R1170 B.n1094 B.n1093 585
R1171 B.n1093 B.n86 585
R1172 B.n1092 B.n85 585
R1173 B.n1158 B.n85 585
R1174 B.n1091 B.n84 585
R1175 B.n1159 B.n84 585
R1176 B.n1090 B.n83 585
R1177 B.n1160 B.n83 585
R1178 B.n1089 B.n1088 585
R1179 B.n1088 B.n79 585
R1180 B.n1087 B.n78 585
R1181 B.n1166 B.n78 585
R1182 B.n1086 B.n77 585
R1183 B.n1167 B.n77 585
R1184 B.n1085 B.n76 585
R1185 B.n1168 B.n76 585
R1186 B.n1084 B.n1083 585
R1187 B.n1083 B.n72 585
R1188 B.n1082 B.n71 585
R1189 B.n1174 B.n71 585
R1190 B.n1081 B.n70 585
R1191 B.n1175 B.n70 585
R1192 B.n1080 B.n69 585
R1193 B.n1176 B.n69 585
R1194 B.n1079 B.n1078 585
R1195 B.n1078 B.n68 585
R1196 B.n1077 B.n64 585
R1197 B.n1182 B.n64 585
R1198 B.n1076 B.n63 585
R1199 B.n1183 B.n63 585
R1200 B.n1075 B.n62 585
R1201 B.n1184 B.n62 585
R1202 B.n1074 B.n1073 585
R1203 B.n1073 B.n58 585
R1204 B.n1072 B.n57 585
R1205 B.n1190 B.n57 585
R1206 B.n1071 B.n56 585
R1207 B.n1191 B.n56 585
R1208 B.n1070 B.n55 585
R1209 B.n1192 B.n55 585
R1210 B.n1069 B.n1068 585
R1211 B.n1068 B.n51 585
R1212 B.n1067 B.n50 585
R1213 B.n1198 B.n50 585
R1214 B.n1066 B.n49 585
R1215 B.n1199 B.n49 585
R1216 B.n1065 B.n48 585
R1217 B.n1200 B.n48 585
R1218 B.n1064 B.n1063 585
R1219 B.n1063 B.n44 585
R1220 B.n1062 B.n43 585
R1221 B.n1206 B.n43 585
R1222 B.n1061 B.n42 585
R1223 B.n1207 B.n42 585
R1224 B.n1060 B.n41 585
R1225 B.n1208 B.n41 585
R1226 B.n1059 B.n1058 585
R1227 B.n1058 B.n37 585
R1228 B.n1057 B.n36 585
R1229 B.n1214 B.n36 585
R1230 B.n1056 B.n35 585
R1231 B.n1215 B.n35 585
R1232 B.n1055 B.n34 585
R1233 B.n1216 B.n34 585
R1234 B.n1054 B.n1053 585
R1235 B.n1053 B.n30 585
R1236 B.n1052 B.n29 585
R1237 B.n1222 B.n29 585
R1238 B.n1051 B.n28 585
R1239 B.n1223 B.n28 585
R1240 B.n1050 B.n27 585
R1241 B.n1224 B.n27 585
R1242 B.n1049 B.n1048 585
R1243 B.n1048 B.n23 585
R1244 B.n1047 B.n22 585
R1245 B.n1230 B.n22 585
R1246 B.n1046 B.n21 585
R1247 B.n1231 B.n21 585
R1248 B.n1045 B.n20 585
R1249 B.n1232 B.n20 585
R1250 B.n1044 B.n1043 585
R1251 B.n1043 B.n16 585
R1252 B.n1042 B.n15 585
R1253 B.n1238 B.n15 585
R1254 B.n1041 B.n14 585
R1255 B.n1239 B.n14 585
R1256 B.n1040 B.n13 585
R1257 B.n1240 B.n13 585
R1258 B.n1039 B.n1038 585
R1259 B.n1038 B.n12 585
R1260 B.n1037 B.n1036 585
R1261 B.n1037 B.n8 585
R1262 B.n1035 B.n7 585
R1263 B.n1247 B.n7 585
R1264 B.n1034 B.n6 585
R1265 B.n1248 B.n6 585
R1266 B.n1033 B.n5 585
R1267 B.n1249 B.n5 585
R1268 B.n1032 B.n1031 585
R1269 B.n1031 B.n4 585
R1270 B.n1030 B.n415 585
R1271 B.n1030 B.n1029 585
R1272 B.n1020 B.n416 585
R1273 B.n417 B.n416 585
R1274 B.n1022 B.n1021 585
R1275 B.n1023 B.n1022 585
R1276 B.n1019 B.n422 585
R1277 B.n422 B.n421 585
R1278 B.n1018 B.n1017 585
R1279 B.n1017 B.n1016 585
R1280 B.n424 B.n423 585
R1281 B.n425 B.n424 585
R1282 B.n1009 B.n1008 585
R1283 B.n1010 B.n1009 585
R1284 B.n1007 B.n430 585
R1285 B.n430 B.n429 585
R1286 B.n1006 B.n1005 585
R1287 B.n1005 B.n1004 585
R1288 B.n432 B.n431 585
R1289 B.n433 B.n432 585
R1290 B.n997 B.n996 585
R1291 B.n998 B.n997 585
R1292 B.n995 B.n438 585
R1293 B.n438 B.n437 585
R1294 B.n994 B.n993 585
R1295 B.n993 B.n992 585
R1296 B.n440 B.n439 585
R1297 B.n441 B.n440 585
R1298 B.n985 B.n984 585
R1299 B.n986 B.n985 585
R1300 B.n983 B.n446 585
R1301 B.n446 B.n445 585
R1302 B.n982 B.n981 585
R1303 B.n981 B.n980 585
R1304 B.n448 B.n447 585
R1305 B.n449 B.n448 585
R1306 B.n973 B.n972 585
R1307 B.n974 B.n973 585
R1308 B.n971 B.n454 585
R1309 B.n454 B.n453 585
R1310 B.n970 B.n969 585
R1311 B.n969 B.n968 585
R1312 B.n456 B.n455 585
R1313 B.n457 B.n456 585
R1314 B.n961 B.n960 585
R1315 B.n962 B.n961 585
R1316 B.n959 B.n461 585
R1317 B.n465 B.n461 585
R1318 B.n958 B.n957 585
R1319 B.n957 B.n956 585
R1320 B.n463 B.n462 585
R1321 B.n464 B.n463 585
R1322 B.n949 B.n948 585
R1323 B.n950 B.n949 585
R1324 B.n947 B.n470 585
R1325 B.n470 B.n469 585
R1326 B.n946 B.n945 585
R1327 B.n945 B.n944 585
R1328 B.n472 B.n471 585
R1329 B.n473 B.n472 585
R1330 B.n937 B.n936 585
R1331 B.n938 B.n937 585
R1332 B.n935 B.n478 585
R1333 B.n478 B.n477 585
R1334 B.n934 B.n933 585
R1335 B.n933 B.n932 585
R1336 B.n480 B.n479 585
R1337 B.n925 B.n480 585
R1338 B.n924 B.n923 585
R1339 B.n926 B.n924 585
R1340 B.n922 B.n485 585
R1341 B.n485 B.n484 585
R1342 B.n921 B.n920 585
R1343 B.n920 B.n919 585
R1344 B.n487 B.n486 585
R1345 B.n488 B.n487 585
R1346 B.n912 B.n911 585
R1347 B.n913 B.n912 585
R1348 B.n910 B.n493 585
R1349 B.n493 B.n492 585
R1350 B.n909 B.n908 585
R1351 B.n908 B.n907 585
R1352 B.n495 B.n494 585
R1353 B.n496 B.n495 585
R1354 B.n900 B.n899 585
R1355 B.n901 B.n900 585
R1356 B.n898 B.n501 585
R1357 B.n501 B.n500 585
R1358 B.n897 B.n896 585
R1359 B.n896 B.n895 585
R1360 B.n503 B.n502 585
R1361 B.n504 B.n503 585
R1362 B.n888 B.n887 585
R1363 B.n889 B.n888 585
R1364 B.n886 B.n509 585
R1365 B.n509 B.n508 585
R1366 B.n885 B.n884 585
R1367 B.n884 B.n883 585
R1368 B.n511 B.n510 585
R1369 B.n512 B.n511 585
R1370 B.n876 B.n875 585
R1371 B.n877 B.n876 585
R1372 B.n874 B.n517 585
R1373 B.n517 B.n516 585
R1374 B.n873 B.n872 585
R1375 B.n872 B.n871 585
R1376 B.n519 B.n518 585
R1377 B.n520 B.n519 585
R1378 B.n864 B.n863 585
R1379 B.n865 B.n864 585
R1380 B.n862 B.n524 585
R1381 B.n528 B.n524 585
R1382 B.n861 B.n860 585
R1383 B.n860 B.n859 585
R1384 B.n526 B.n525 585
R1385 B.n527 B.n526 585
R1386 B.n852 B.n851 585
R1387 B.n853 B.n852 585
R1388 B.n850 B.n533 585
R1389 B.n533 B.n532 585
R1390 B.n849 B.n848 585
R1391 B.n848 B.n847 585
R1392 B.n535 B.n534 585
R1393 B.n536 B.n535 585
R1394 B.n840 B.n839 585
R1395 B.n841 B.n840 585
R1396 B.n539 B.n538 585
R1397 B.n604 B.n602 585
R1398 B.n605 B.n601 585
R1399 B.n605 B.n540 585
R1400 B.n608 B.n607 585
R1401 B.n609 B.n600 585
R1402 B.n611 B.n610 585
R1403 B.n613 B.n599 585
R1404 B.n616 B.n615 585
R1405 B.n617 B.n598 585
R1406 B.n619 B.n618 585
R1407 B.n621 B.n597 585
R1408 B.n624 B.n623 585
R1409 B.n625 B.n596 585
R1410 B.n627 B.n626 585
R1411 B.n629 B.n595 585
R1412 B.n632 B.n631 585
R1413 B.n633 B.n594 585
R1414 B.n635 B.n634 585
R1415 B.n637 B.n593 585
R1416 B.n640 B.n639 585
R1417 B.n641 B.n592 585
R1418 B.n643 B.n642 585
R1419 B.n645 B.n591 585
R1420 B.n648 B.n647 585
R1421 B.n649 B.n590 585
R1422 B.n651 B.n650 585
R1423 B.n653 B.n589 585
R1424 B.n656 B.n655 585
R1425 B.n657 B.n588 585
R1426 B.n659 B.n658 585
R1427 B.n661 B.n587 585
R1428 B.n664 B.n663 585
R1429 B.n665 B.n586 585
R1430 B.n667 B.n666 585
R1431 B.n669 B.n585 585
R1432 B.n672 B.n671 585
R1433 B.n673 B.n584 585
R1434 B.n675 B.n674 585
R1435 B.n677 B.n583 585
R1436 B.n680 B.n679 585
R1437 B.n681 B.n582 585
R1438 B.n683 B.n682 585
R1439 B.n685 B.n581 585
R1440 B.n688 B.n687 585
R1441 B.n689 B.n580 585
R1442 B.n691 B.n690 585
R1443 B.n693 B.n579 585
R1444 B.n696 B.n695 585
R1445 B.n697 B.n578 585
R1446 B.n699 B.n698 585
R1447 B.n701 B.n577 585
R1448 B.n704 B.n703 585
R1449 B.n705 B.n576 585
R1450 B.n710 B.n709 585
R1451 B.n712 B.n575 585
R1452 B.n715 B.n714 585
R1453 B.n716 B.n574 585
R1454 B.n718 B.n717 585
R1455 B.n720 B.n573 585
R1456 B.n723 B.n722 585
R1457 B.n724 B.n572 585
R1458 B.n726 B.n725 585
R1459 B.n728 B.n571 585
R1460 B.n731 B.n730 585
R1461 B.n733 B.n568 585
R1462 B.n735 B.n734 585
R1463 B.n737 B.n567 585
R1464 B.n740 B.n739 585
R1465 B.n741 B.n566 585
R1466 B.n743 B.n742 585
R1467 B.n745 B.n565 585
R1468 B.n748 B.n747 585
R1469 B.n749 B.n564 585
R1470 B.n751 B.n750 585
R1471 B.n753 B.n563 585
R1472 B.n756 B.n755 585
R1473 B.n757 B.n562 585
R1474 B.n759 B.n758 585
R1475 B.n761 B.n561 585
R1476 B.n764 B.n763 585
R1477 B.n765 B.n560 585
R1478 B.n767 B.n766 585
R1479 B.n769 B.n559 585
R1480 B.n772 B.n771 585
R1481 B.n773 B.n558 585
R1482 B.n775 B.n774 585
R1483 B.n777 B.n557 585
R1484 B.n780 B.n779 585
R1485 B.n781 B.n556 585
R1486 B.n783 B.n782 585
R1487 B.n785 B.n555 585
R1488 B.n788 B.n787 585
R1489 B.n789 B.n554 585
R1490 B.n791 B.n790 585
R1491 B.n793 B.n553 585
R1492 B.n796 B.n795 585
R1493 B.n797 B.n552 585
R1494 B.n799 B.n798 585
R1495 B.n801 B.n551 585
R1496 B.n804 B.n803 585
R1497 B.n805 B.n550 585
R1498 B.n807 B.n806 585
R1499 B.n809 B.n549 585
R1500 B.n812 B.n811 585
R1501 B.n813 B.n548 585
R1502 B.n815 B.n814 585
R1503 B.n817 B.n547 585
R1504 B.n820 B.n819 585
R1505 B.n821 B.n546 585
R1506 B.n823 B.n822 585
R1507 B.n825 B.n545 585
R1508 B.n828 B.n827 585
R1509 B.n829 B.n544 585
R1510 B.n831 B.n830 585
R1511 B.n833 B.n543 585
R1512 B.n834 B.n542 585
R1513 B.n837 B.n836 585
R1514 B.n838 B.n541 585
R1515 B.n541 B.n540 585
R1516 B.n843 B.n842 585
R1517 B.n842 B.n841 585
R1518 B.n844 B.n537 585
R1519 B.n537 B.n536 585
R1520 B.n846 B.n845 585
R1521 B.n847 B.n846 585
R1522 B.n531 B.n530 585
R1523 B.n532 B.n531 585
R1524 B.n855 B.n854 585
R1525 B.n854 B.n853 585
R1526 B.n856 B.n529 585
R1527 B.n529 B.n527 585
R1528 B.n858 B.n857 585
R1529 B.n859 B.n858 585
R1530 B.n523 B.n522 585
R1531 B.n528 B.n523 585
R1532 B.n867 B.n866 585
R1533 B.n866 B.n865 585
R1534 B.n868 B.n521 585
R1535 B.n521 B.n520 585
R1536 B.n870 B.n869 585
R1537 B.n871 B.n870 585
R1538 B.n515 B.n514 585
R1539 B.n516 B.n515 585
R1540 B.n879 B.n878 585
R1541 B.n878 B.n877 585
R1542 B.n880 B.n513 585
R1543 B.n513 B.n512 585
R1544 B.n882 B.n881 585
R1545 B.n883 B.n882 585
R1546 B.n507 B.n506 585
R1547 B.n508 B.n507 585
R1548 B.n891 B.n890 585
R1549 B.n890 B.n889 585
R1550 B.n892 B.n505 585
R1551 B.n505 B.n504 585
R1552 B.n894 B.n893 585
R1553 B.n895 B.n894 585
R1554 B.n499 B.n498 585
R1555 B.n500 B.n499 585
R1556 B.n903 B.n902 585
R1557 B.n902 B.n901 585
R1558 B.n904 B.n497 585
R1559 B.n497 B.n496 585
R1560 B.n906 B.n905 585
R1561 B.n907 B.n906 585
R1562 B.n491 B.n490 585
R1563 B.n492 B.n491 585
R1564 B.n915 B.n914 585
R1565 B.n914 B.n913 585
R1566 B.n916 B.n489 585
R1567 B.n489 B.n488 585
R1568 B.n918 B.n917 585
R1569 B.n919 B.n918 585
R1570 B.n483 B.n482 585
R1571 B.n484 B.n483 585
R1572 B.n928 B.n927 585
R1573 B.n927 B.n926 585
R1574 B.n929 B.n481 585
R1575 B.n925 B.n481 585
R1576 B.n931 B.n930 585
R1577 B.n932 B.n931 585
R1578 B.n476 B.n475 585
R1579 B.n477 B.n476 585
R1580 B.n940 B.n939 585
R1581 B.n939 B.n938 585
R1582 B.n941 B.n474 585
R1583 B.n474 B.n473 585
R1584 B.n943 B.n942 585
R1585 B.n944 B.n943 585
R1586 B.n468 B.n467 585
R1587 B.n469 B.n468 585
R1588 B.n952 B.n951 585
R1589 B.n951 B.n950 585
R1590 B.n953 B.n466 585
R1591 B.n466 B.n464 585
R1592 B.n955 B.n954 585
R1593 B.n956 B.n955 585
R1594 B.n460 B.n459 585
R1595 B.n465 B.n460 585
R1596 B.n964 B.n963 585
R1597 B.n963 B.n962 585
R1598 B.n965 B.n458 585
R1599 B.n458 B.n457 585
R1600 B.n967 B.n966 585
R1601 B.n968 B.n967 585
R1602 B.n452 B.n451 585
R1603 B.n453 B.n452 585
R1604 B.n976 B.n975 585
R1605 B.n975 B.n974 585
R1606 B.n977 B.n450 585
R1607 B.n450 B.n449 585
R1608 B.n979 B.n978 585
R1609 B.n980 B.n979 585
R1610 B.n444 B.n443 585
R1611 B.n445 B.n444 585
R1612 B.n988 B.n987 585
R1613 B.n987 B.n986 585
R1614 B.n989 B.n442 585
R1615 B.n442 B.n441 585
R1616 B.n991 B.n990 585
R1617 B.n992 B.n991 585
R1618 B.n436 B.n435 585
R1619 B.n437 B.n436 585
R1620 B.n1000 B.n999 585
R1621 B.n999 B.n998 585
R1622 B.n1001 B.n434 585
R1623 B.n434 B.n433 585
R1624 B.n1003 B.n1002 585
R1625 B.n1004 B.n1003 585
R1626 B.n428 B.n427 585
R1627 B.n429 B.n428 585
R1628 B.n1012 B.n1011 585
R1629 B.n1011 B.n1010 585
R1630 B.n1013 B.n426 585
R1631 B.n426 B.n425 585
R1632 B.n1015 B.n1014 585
R1633 B.n1016 B.n1015 585
R1634 B.n420 B.n419 585
R1635 B.n421 B.n420 585
R1636 B.n1025 B.n1024 585
R1637 B.n1024 B.n1023 585
R1638 B.n1026 B.n418 585
R1639 B.n418 B.n417 585
R1640 B.n1028 B.n1027 585
R1641 B.n1029 B.n1028 585
R1642 B.n3 B.n0 585
R1643 B.n4 B.n3 585
R1644 B.n1246 B.n1 585
R1645 B.n1247 B.n1246 585
R1646 B.n1245 B.n1244 585
R1647 B.n1245 B.n8 585
R1648 B.n1243 B.n9 585
R1649 B.n12 B.n9 585
R1650 B.n1242 B.n1241 585
R1651 B.n1241 B.n1240 585
R1652 B.n11 B.n10 585
R1653 B.n1239 B.n11 585
R1654 B.n1237 B.n1236 585
R1655 B.n1238 B.n1237 585
R1656 B.n1235 B.n17 585
R1657 B.n17 B.n16 585
R1658 B.n1234 B.n1233 585
R1659 B.n1233 B.n1232 585
R1660 B.n19 B.n18 585
R1661 B.n1231 B.n19 585
R1662 B.n1229 B.n1228 585
R1663 B.n1230 B.n1229 585
R1664 B.n1227 B.n24 585
R1665 B.n24 B.n23 585
R1666 B.n1226 B.n1225 585
R1667 B.n1225 B.n1224 585
R1668 B.n26 B.n25 585
R1669 B.n1223 B.n26 585
R1670 B.n1221 B.n1220 585
R1671 B.n1222 B.n1221 585
R1672 B.n1219 B.n31 585
R1673 B.n31 B.n30 585
R1674 B.n1218 B.n1217 585
R1675 B.n1217 B.n1216 585
R1676 B.n33 B.n32 585
R1677 B.n1215 B.n33 585
R1678 B.n1213 B.n1212 585
R1679 B.n1214 B.n1213 585
R1680 B.n1211 B.n38 585
R1681 B.n38 B.n37 585
R1682 B.n1210 B.n1209 585
R1683 B.n1209 B.n1208 585
R1684 B.n40 B.n39 585
R1685 B.n1207 B.n40 585
R1686 B.n1205 B.n1204 585
R1687 B.n1206 B.n1205 585
R1688 B.n1203 B.n45 585
R1689 B.n45 B.n44 585
R1690 B.n1202 B.n1201 585
R1691 B.n1201 B.n1200 585
R1692 B.n47 B.n46 585
R1693 B.n1199 B.n47 585
R1694 B.n1197 B.n1196 585
R1695 B.n1198 B.n1197 585
R1696 B.n1195 B.n52 585
R1697 B.n52 B.n51 585
R1698 B.n1194 B.n1193 585
R1699 B.n1193 B.n1192 585
R1700 B.n54 B.n53 585
R1701 B.n1191 B.n54 585
R1702 B.n1189 B.n1188 585
R1703 B.n1190 B.n1189 585
R1704 B.n1187 B.n59 585
R1705 B.n59 B.n58 585
R1706 B.n1186 B.n1185 585
R1707 B.n1185 B.n1184 585
R1708 B.n61 B.n60 585
R1709 B.n1183 B.n61 585
R1710 B.n1181 B.n1180 585
R1711 B.n1182 B.n1181 585
R1712 B.n1179 B.n65 585
R1713 B.n68 B.n65 585
R1714 B.n1178 B.n1177 585
R1715 B.n1177 B.n1176 585
R1716 B.n67 B.n66 585
R1717 B.n1175 B.n67 585
R1718 B.n1173 B.n1172 585
R1719 B.n1174 B.n1173 585
R1720 B.n1171 B.n73 585
R1721 B.n73 B.n72 585
R1722 B.n1170 B.n1169 585
R1723 B.n1169 B.n1168 585
R1724 B.n75 B.n74 585
R1725 B.n1167 B.n75 585
R1726 B.n1165 B.n1164 585
R1727 B.n1166 B.n1165 585
R1728 B.n1163 B.n80 585
R1729 B.n80 B.n79 585
R1730 B.n1162 B.n1161 585
R1731 B.n1161 B.n1160 585
R1732 B.n82 B.n81 585
R1733 B.n1159 B.n82 585
R1734 B.n1157 B.n1156 585
R1735 B.n1158 B.n1157 585
R1736 B.n1155 B.n87 585
R1737 B.n87 B.n86 585
R1738 B.n1154 B.n1153 585
R1739 B.n1153 B.n1152 585
R1740 B.n89 B.n88 585
R1741 B.n1151 B.n89 585
R1742 B.n1149 B.n1148 585
R1743 B.n1150 B.n1149 585
R1744 B.n1147 B.n94 585
R1745 B.n94 B.n93 585
R1746 B.n1146 B.n1145 585
R1747 B.n1145 B.n1144 585
R1748 B.n96 B.n95 585
R1749 B.n1143 B.n96 585
R1750 B.n1141 B.n1140 585
R1751 B.n1142 B.n1141 585
R1752 B.n1139 B.n101 585
R1753 B.n101 B.n100 585
R1754 B.n1138 B.n1137 585
R1755 B.n1137 B.n1136 585
R1756 B.n103 B.n102 585
R1757 B.n1135 B.n103 585
R1758 B.n1133 B.n1132 585
R1759 B.n1134 B.n1133 585
R1760 B.n1131 B.n108 585
R1761 B.n108 B.n107 585
R1762 B.n1130 B.n1129 585
R1763 B.n1129 B.n1128 585
R1764 B.n110 B.n109 585
R1765 B.n1127 B.n110 585
R1766 B.n1125 B.n1124 585
R1767 B.n1126 B.n1125 585
R1768 B.n1123 B.n115 585
R1769 B.n115 B.n114 585
R1770 B.n1122 B.n1121 585
R1771 B.n1121 B.n1120 585
R1772 B.n1250 B.n1249 585
R1773 B.n1248 B.n2 585
R1774 B.n1121 B.n117 478.086
R1775 B.n1117 B.n118 478.086
R1776 B.n840 B.n541 478.086
R1777 B.n842 B.n539 478.086
R1778 B.n178 B.t12 416.865
R1779 B.n569 B.t20 416.865
R1780 B.n181 B.t15 416.865
R1781 B.n706 B.t23 416.865
R1782 B.n179 B.t13 354.803
R1783 B.n570 B.t19 354.803
R1784 B.n182 B.t16 354.803
R1785 B.n707 B.t22 354.803
R1786 B.n181 B.t14 344.539
R1787 B.n178 B.t10 344.539
R1788 B.n569 B.t17 344.539
R1789 B.n706 B.t21 344.539
R1790 B.n1119 B.n1118 256.663
R1791 B.n1119 B.n176 256.663
R1792 B.n1119 B.n175 256.663
R1793 B.n1119 B.n174 256.663
R1794 B.n1119 B.n173 256.663
R1795 B.n1119 B.n172 256.663
R1796 B.n1119 B.n171 256.663
R1797 B.n1119 B.n170 256.663
R1798 B.n1119 B.n169 256.663
R1799 B.n1119 B.n168 256.663
R1800 B.n1119 B.n167 256.663
R1801 B.n1119 B.n166 256.663
R1802 B.n1119 B.n165 256.663
R1803 B.n1119 B.n164 256.663
R1804 B.n1119 B.n163 256.663
R1805 B.n1119 B.n162 256.663
R1806 B.n1119 B.n161 256.663
R1807 B.n1119 B.n160 256.663
R1808 B.n1119 B.n159 256.663
R1809 B.n1119 B.n158 256.663
R1810 B.n1119 B.n157 256.663
R1811 B.n1119 B.n156 256.663
R1812 B.n1119 B.n155 256.663
R1813 B.n1119 B.n154 256.663
R1814 B.n1119 B.n153 256.663
R1815 B.n1119 B.n152 256.663
R1816 B.n1119 B.n151 256.663
R1817 B.n1119 B.n150 256.663
R1818 B.n1119 B.n149 256.663
R1819 B.n1119 B.n148 256.663
R1820 B.n1119 B.n147 256.663
R1821 B.n1119 B.n146 256.663
R1822 B.n1119 B.n145 256.663
R1823 B.n1119 B.n144 256.663
R1824 B.n1119 B.n143 256.663
R1825 B.n1119 B.n142 256.663
R1826 B.n1119 B.n141 256.663
R1827 B.n1119 B.n140 256.663
R1828 B.n1119 B.n139 256.663
R1829 B.n1119 B.n138 256.663
R1830 B.n1119 B.n137 256.663
R1831 B.n1119 B.n136 256.663
R1832 B.n1119 B.n135 256.663
R1833 B.n1119 B.n134 256.663
R1834 B.n1119 B.n133 256.663
R1835 B.n1119 B.n132 256.663
R1836 B.n1119 B.n131 256.663
R1837 B.n1119 B.n130 256.663
R1838 B.n1119 B.n129 256.663
R1839 B.n1119 B.n128 256.663
R1840 B.n1119 B.n127 256.663
R1841 B.n1119 B.n126 256.663
R1842 B.n1119 B.n125 256.663
R1843 B.n1119 B.n124 256.663
R1844 B.n1119 B.n123 256.663
R1845 B.n1119 B.n122 256.663
R1846 B.n1119 B.n121 256.663
R1847 B.n1119 B.n120 256.663
R1848 B.n1119 B.n119 256.663
R1849 B.n603 B.n540 256.663
R1850 B.n606 B.n540 256.663
R1851 B.n612 B.n540 256.663
R1852 B.n614 B.n540 256.663
R1853 B.n620 B.n540 256.663
R1854 B.n622 B.n540 256.663
R1855 B.n628 B.n540 256.663
R1856 B.n630 B.n540 256.663
R1857 B.n636 B.n540 256.663
R1858 B.n638 B.n540 256.663
R1859 B.n644 B.n540 256.663
R1860 B.n646 B.n540 256.663
R1861 B.n652 B.n540 256.663
R1862 B.n654 B.n540 256.663
R1863 B.n660 B.n540 256.663
R1864 B.n662 B.n540 256.663
R1865 B.n668 B.n540 256.663
R1866 B.n670 B.n540 256.663
R1867 B.n676 B.n540 256.663
R1868 B.n678 B.n540 256.663
R1869 B.n684 B.n540 256.663
R1870 B.n686 B.n540 256.663
R1871 B.n692 B.n540 256.663
R1872 B.n694 B.n540 256.663
R1873 B.n700 B.n540 256.663
R1874 B.n702 B.n540 256.663
R1875 B.n711 B.n540 256.663
R1876 B.n713 B.n540 256.663
R1877 B.n719 B.n540 256.663
R1878 B.n721 B.n540 256.663
R1879 B.n727 B.n540 256.663
R1880 B.n729 B.n540 256.663
R1881 B.n736 B.n540 256.663
R1882 B.n738 B.n540 256.663
R1883 B.n744 B.n540 256.663
R1884 B.n746 B.n540 256.663
R1885 B.n752 B.n540 256.663
R1886 B.n754 B.n540 256.663
R1887 B.n760 B.n540 256.663
R1888 B.n762 B.n540 256.663
R1889 B.n768 B.n540 256.663
R1890 B.n770 B.n540 256.663
R1891 B.n776 B.n540 256.663
R1892 B.n778 B.n540 256.663
R1893 B.n784 B.n540 256.663
R1894 B.n786 B.n540 256.663
R1895 B.n792 B.n540 256.663
R1896 B.n794 B.n540 256.663
R1897 B.n800 B.n540 256.663
R1898 B.n802 B.n540 256.663
R1899 B.n808 B.n540 256.663
R1900 B.n810 B.n540 256.663
R1901 B.n816 B.n540 256.663
R1902 B.n818 B.n540 256.663
R1903 B.n824 B.n540 256.663
R1904 B.n826 B.n540 256.663
R1905 B.n832 B.n540 256.663
R1906 B.n835 B.n540 256.663
R1907 B.n1252 B.n1251 256.663
R1908 B.n186 B.n185 163.367
R1909 B.n190 B.n189 163.367
R1910 B.n194 B.n193 163.367
R1911 B.n198 B.n197 163.367
R1912 B.n202 B.n201 163.367
R1913 B.n206 B.n205 163.367
R1914 B.n210 B.n209 163.367
R1915 B.n214 B.n213 163.367
R1916 B.n218 B.n217 163.367
R1917 B.n222 B.n221 163.367
R1918 B.n226 B.n225 163.367
R1919 B.n230 B.n229 163.367
R1920 B.n234 B.n233 163.367
R1921 B.n238 B.n237 163.367
R1922 B.n242 B.n241 163.367
R1923 B.n246 B.n245 163.367
R1924 B.n250 B.n249 163.367
R1925 B.n254 B.n253 163.367
R1926 B.n258 B.n257 163.367
R1927 B.n262 B.n261 163.367
R1928 B.n266 B.n265 163.367
R1929 B.n270 B.n269 163.367
R1930 B.n274 B.n273 163.367
R1931 B.n278 B.n277 163.367
R1932 B.n282 B.n281 163.367
R1933 B.n286 B.n285 163.367
R1934 B.n290 B.n289 163.367
R1935 B.n294 B.n293 163.367
R1936 B.n298 B.n297 163.367
R1937 B.n302 B.n301 163.367
R1938 B.n306 B.n305 163.367
R1939 B.n310 B.n309 163.367
R1940 B.n314 B.n313 163.367
R1941 B.n318 B.n317 163.367
R1942 B.n322 B.n321 163.367
R1943 B.n326 B.n325 163.367
R1944 B.n330 B.n329 163.367
R1945 B.n334 B.n333 163.367
R1946 B.n338 B.n337 163.367
R1947 B.n342 B.n341 163.367
R1948 B.n346 B.n345 163.367
R1949 B.n350 B.n349 163.367
R1950 B.n354 B.n353 163.367
R1951 B.n358 B.n357 163.367
R1952 B.n362 B.n361 163.367
R1953 B.n366 B.n365 163.367
R1954 B.n370 B.n369 163.367
R1955 B.n374 B.n373 163.367
R1956 B.n378 B.n377 163.367
R1957 B.n382 B.n381 163.367
R1958 B.n386 B.n385 163.367
R1959 B.n390 B.n389 163.367
R1960 B.n394 B.n393 163.367
R1961 B.n398 B.n397 163.367
R1962 B.n402 B.n401 163.367
R1963 B.n406 B.n405 163.367
R1964 B.n410 B.n409 163.367
R1965 B.n412 B.n177 163.367
R1966 B.n840 B.n535 163.367
R1967 B.n848 B.n535 163.367
R1968 B.n848 B.n533 163.367
R1969 B.n852 B.n533 163.367
R1970 B.n852 B.n526 163.367
R1971 B.n860 B.n526 163.367
R1972 B.n860 B.n524 163.367
R1973 B.n864 B.n524 163.367
R1974 B.n864 B.n519 163.367
R1975 B.n872 B.n519 163.367
R1976 B.n872 B.n517 163.367
R1977 B.n876 B.n517 163.367
R1978 B.n876 B.n511 163.367
R1979 B.n884 B.n511 163.367
R1980 B.n884 B.n509 163.367
R1981 B.n888 B.n509 163.367
R1982 B.n888 B.n503 163.367
R1983 B.n896 B.n503 163.367
R1984 B.n896 B.n501 163.367
R1985 B.n900 B.n501 163.367
R1986 B.n900 B.n495 163.367
R1987 B.n908 B.n495 163.367
R1988 B.n908 B.n493 163.367
R1989 B.n912 B.n493 163.367
R1990 B.n912 B.n487 163.367
R1991 B.n920 B.n487 163.367
R1992 B.n920 B.n485 163.367
R1993 B.n924 B.n485 163.367
R1994 B.n924 B.n480 163.367
R1995 B.n933 B.n480 163.367
R1996 B.n933 B.n478 163.367
R1997 B.n937 B.n478 163.367
R1998 B.n937 B.n472 163.367
R1999 B.n945 B.n472 163.367
R2000 B.n945 B.n470 163.367
R2001 B.n949 B.n470 163.367
R2002 B.n949 B.n463 163.367
R2003 B.n957 B.n463 163.367
R2004 B.n957 B.n461 163.367
R2005 B.n961 B.n461 163.367
R2006 B.n961 B.n456 163.367
R2007 B.n969 B.n456 163.367
R2008 B.n969 B.n454 163.367
R2009 B.n973 B.n454 163.367
R2010 B.n973 B.n448 163.367
R2011 B.n981 B.n448 163.367
R2012 B.n981 B.n446 163.367
R2013 B.n985 B.n446 163.367
R2014 B.n985 B.n440 163.367
R2015 B.n993 B.n440 163.367
R2016 B.n993 B.n438 163.367
R2017 B.n997 B.n438 163.367
R2018 B.n997 B.n432 163.367
R2019 B.n1005 B.n432 163.367
R2020 B.n1005 B.n430 163.367
R2021 B.n1009 B.n430 163.367
R2022 B.n1009 B.n424 163.367
R2023 B.n1017 B.n424 163.367
R2024 B.n1017 B.n422 163.367
R2025 B.n1022 B.n422 163.367
R2026 B.n1022 B.n416 163.367
R2027 B.n1030 B.n416 163.367
R2028 B.n1031 B.n1030 163.367
R2029 B.n1031 B.n5 163.367
R2030 B.n6 B.n5 163.367
R2031 B.n7 B.n6 163.367
R2032 B.n1037 B.n7 163.367
R2033 B.n1038 B.n1037 163.367
R2034 B.n1038 B.n13 163.367
R2035 B.n14 B.n13 163.367
R2036 B.n15 B.n14 163.367
R2037 B.n1043 B.n15 163.367
R2038 B.n1043 B.n20 163.367
R2039 B.n21 B.n20 163.367
R2040 B.n22 B.n21 163.367
R2041 B.n1048 B.n22 163.367
R2042 B.n1048 B.n27 163.367
R2043 B.n28 B.n27 163.367
R2044 B.n29 B.n28 163.367
R2045 B.n1053 B.n29 163.367
R2046 B.n1053 B.n34 163.367
R2047 B.n35 B.n34 163.367
R2048 B.n36 B.n35 163.367
R2049 B.n1058 B.n36 163.367
R2050 B.n1058 B.n41 163.367
R2051 B.n42 B.n41 163.367
R2052 B.n43 B.n42 163.367
R2053 B.n1063 B.n43 163.367
R2054 B.n1063 B.n48 163.367
R2055 B.n49 B.n48 163.367
R2056 B.n50 B.n49 163.367
R2057 B.n1068 B.n50 163.367
R2058 B.n1068 B.n55 163.367
R2059 B.n56 B.n55 163.367
R2060 B.n57 B.n56 163.367
R2061 B.n1073 B.n57 163.367
R2062 B.n1073 B.n62 163.367
R2063 B.n63 B.n62 163.367
R2064 B.n64 B.n63 163.367
R2065 B.n1078 B.n64 163.367
R2066 B.n1078 B.n69 163.367
R2067 B.n70 B.n69 163.367
R2068 B.n71 B.n70 163.367
R2069 B.n1083 B.n71 163.367
R2070 B.n1083 B.n76 163.367
R2071 B.n77 B.n76 163.367
R2072 B.n78 B.n77 163.367
R2073 B.n1088 B.n78 163.367
R2074 B.n1088 B.n83 163.367
R2075 B.n84 B.n83 163.367
R2076 B.n85 B.n84 163.367
R2077 B.n1093 B.n85 163.367
R2078 B.n1093 B.n90 163.367
R2079 B.n91 B.n90 163.367
R2080 B.n92 B.n91 163.367
R2081 B.n1098 B.n92 163.367
R2082 B.n1098 B.n97 163.367
R2083 B.n98 B.n97 163.367
R2084 B.n99 B.n98 163.367
R2085 B.n1103 B.n99 163.367
R2086 B.n1103 B.n104 163.367
R2087 B.n105 B.n104 163.367
R2088 B.n106 B.n105 163.367
R2089 B.n1108 B.n106 163.367
R2090 B.n1108 B.n111 163.367
R2091 B.n112 B.n111 163.367
R2092 B.n113 B.n112 163.367
R2093 B.n1113 B.n113 163.367
R2094 B.n1113 B.n118 163.367
R2095 B.n605 B.n604 163.367
R2096 B.n607 B.n605 163.367
R2097 B.n611 B.n600 163.367
R2098 B.n615 B.n613 163.367
R2099 B.n619 B.n598 163.367
R2100 B.n623 B.n621 163.367
R2101 B.n627 B.n596 163.367
R2102 B.n631 B.n629 163.367
R2103 B.n635 B.n594 163.367
R2104 B.n639 B.n637 163.367
R2105 B.n643 B.n592 163.367
R2106 B.n647 B.n645 163.367
R2107 B.n651 B.n590 163.367
R2108 B.n655 B.n653 163.367
R2109 B.n659 B.n588 163.367
R2110 B.n663 B.n661 163.367
R2111 B.n667 B.n586 163.367
R2112 B.n671 B.n669 163.367
R2113 B.n675 B.n584 163.367
R2114 B.n679 B.n677 163.367
R2115 B.n683 B.n582 163.367
R2116 B.n687 B.n685 163.367
R2117 B.n691 B.n580 163.367
R2118 B.n695 B.n693 163.367
R2119 B.n699 B.n578 163.367
R2120 B.n703 B.n701 163.367
R2121 B.n710 B.n576 163.367
R2122 B.n714 B.n712 163.367
R2123 B.n718 B.n574 163.367
R2124 B.n722 B.n720 163.367
R2125 B.n726 B.n572 163.367
R2126 B.n730 B.n728 163.367
R2127 B.n735 B.n568 163.367
R2128 B.n739 B.n737 163.367
R2129 B.n743 B.n566 163.367
R2130 B.n747 B.n745 163.367
R2131 B.n751 B.n564 163.367
R2132 B.n755 B.n753 163.367
R2133 B.n759 B.n562 163.367
R2134 B.n763 B.n761 163.367
R2135 B.n767 B.n560 163.367
R2136 B.n771 B.n769 163.367
R2137 B.n775 B.n558 163.367
R2138 B.n779 B.n777 163.367
R2139 B.n783 B.n556 163.367
R2140 B.n787 B.n785 163.367
R2141 B.n791 B.n554 163.367
R2142 B.n795 B.n793 163.367
R2143 B.n799 B.n552 163.367
R2144 B.n803 B.n801 163.367
R2145 B.n807 B.n550 163.367
R2146 B.n811 B.n809 163.367
R2147 B.n815 B.n548 163.367
R2148 B.n819 B.n817 163.367
R2149 B.n823 B.n546 163.367
R2150 B.n827 B.n825 163.367
R2151 B.n831 B.n544 163.367
R2152 B.n834 B.n833 163.367
R2153 B.n836 B.n541 163.367
R2154 B.n842 B.n537 163.367
R2155 B.n846 B.n537 163.367
R2156 B.n846 B.n531 163.367
R2157 B.n854 B.n531 163.367
R2158 B.n854 B.n529 163.367
R2159 B.n858 B.n529 163.367
R2160 B.n858 B.n523 163.367
R2161 B.n866 B.n523 163.367
R2162 B.n866 B.n521 163.367
R2163 B.n870 B.n521 163.367
R2164 B.n870 B.n515 163.367
R2165 B.n878 B.n515 163.367
R2166 B.n878 B.n513 163.367
R2167 B.n882 B.n513 163.367
R2168 B.n882 B.n507 163.367
R2169 B.n890 B.n507 163.367
R2170 B.n890 B.n505 163.367
R2171 B.n894 B.n505 163.367
R2172 B.n894 B.n499 163.367
R2173 B.n902 B.n499 163.367
R2174 B.n902 B.n497 163.367
R2175 B.n906 B.n497 163.367
R2176 B.n906 B.n491 163.367
R2177 B.n914 B.n491 163.367
R2178 B.n914 B.n489 163.367
R2179 B.n918 B.n489 163.367
R2180 B.n918 B.n483 163.367
R2181 B.n927 B.n483 163.367
R2182 B.n927 B.n481 163.367
R2183 B.n931 B.n481 163.367
R2184 B.n931 B.n476 163.367
R2185 B.n939 B.n476 163.367
R2186 B.n939 B.n474 163.367
R2187 B.n943 B.n474 163.367
R2188 B.n943 B.n468 163.367
R2189 B.n951 B.n468 163.367
R2190 B.n951 B.n466 163.367
R2191 B.n955 B.n466 163.367
R2192 B.n955 B.n460 163.367
R2193 B.n963 B.n460 163.367
R2194 B.n963 B.n458 163.367
R2195 B.n967 B.n458 163.367
R2196 B.n967 B.n452 163.367
R2197 B.n975 B.n452 163.367
R2198 B.n975 B.n450 163.367
R2199 B.n979 B.n450 163.367
R2200 B.n979 B.n444 163.367
R2201 B.n987 B.n444 163.367
R2202 B.n987 B.n442 163.367
R2203 B.n991 B.n442 163.367
R2204 B.n991 B.n436 163.367
R2205 B.n999 B.n436 163.367
R2206 B.n999 B.n434 163.367
R2207 B.n1003 B.n434 163.367
R2208 B.n1003 B.n428 163.367
R2209 B.n1011 B.n428 163.367
R2210 B.n1011 B.n426 163.367
R2211 B.n1015 B.n426 163.367
R2212 B.n1015 B.n420 163.367
R2213 B.n1024 B.n420 163.367
R2214 B.n1024 B.n418 163.367
R2215 B.n1028 B.n418 163.367
R2216 B.n1028 B.n3 163.367
R2217 B.n1250 B.n3 163.367
R2218 B.n1246 B.n2 163.367
R2219 B.n1246 B.n1245 163.367
R2220 B.n1245 B.n9 163.367
R2221 B.n1241 B.n9 163.367
R2222 B.n1241 B.n11 163.367
R2223 B.n1237 B.n11 163.367
R2224 B.n1237 B.n17 163.367
R2225 B.n1233 B.n17 163.367
R2226 B.n1233 B.n19 163.367
R2227 B.n1229 B.n19 163.367
R2228 B.n1229 B.n24 163.367
R2229 B.n1225 B.n24 163.367
R2230 B.n1225 B.n26 163.367
R2231 B.n1221 B.n26 163.367
R2232 B.n1221 B.n31 163.367
R2233 B.n1217 B.n31 163.367
R2234 B.n1217 B.n33 163.367
R2235 B.n1213 B.n33 163.367
R2236 B.n1213 B.n38 163.367
R2237 B.n1209 B.n38 163.367
R2238 B.n1209 B.n40 163.367
R2239 B.n1205 B.n40 163.367
R2240 B.n1205 B.n45 163.367
R2241 B.n1201 B.n45 163.367
R2242 B.n1201 B.n47 163.367
R2243 B.n1197 B.n47 163.367
R2244 B.n1197 B.n52 163.367
R2245 B.n1193 B.n52 163.367
R2246 B.n1193 B.n54 163.367
R2247 B.n1189 B.n54 163.367
R2248 B.n1189 B.n59 163.367
R2249 B.n1185 B.n59 163.367
R2250 B.n1185 B.n61 163.367
R2251 B.n1181 B.n61 163.367
R2252 B.n1181 B.n65 163.367
R2253 B.n1177 B.n65 163.367
R2254 B.n1177 B.n67 163.367
R2255 B.n1173 B.n67 163.367
R2256 B.n1173 B.n73 163.367
R2257 B.n1169 B.n73 163.367
R2258 B.n1169 B.n75 163.367
R2259 B.n1165 B.n75 163.367
R2260 B.n1165 B.n80 163.367
R2261 B.n1161 B.n80 163.367
R2262 B.n1161 B.n82 163.367
R2263 B.n1157 B.n82 163.367
R2264 B.n1157 B.n87 163.367
R2265 B.n1153 B.n87 163.367
R2266 B.n1153 B.n89 163.367
R2267 B.n1149 B.n89 163.367
R2268 B.n1149 B.n94 163.367
R2269 B.n1145 B.n94 163.367
R2270 B.n1145 B.n96 163.367
R2271 B.n1141 B.n96 163.367
R2272 B.n1141 B.n101 163.367
R2273 B.n1137 B.n101 163.367
R2274 B.n1137 B.n103 163.367
R2275 B.n1133 B.n103 163.367
R2276 B.n1133 B.n108 163.367
R2277 B.n1129 B.n108 163.367
R2278 B.n1129 B.n110 163.367
R2279 B.n1125 B.n110 163.367
R2280 B.n1125 B.n115 163.367
R2281 B.n1121 B.n115 163.367
R2282 B.n119 B.n117 71.676
R2283 B.n186 B.n120 71.676
R2284 B.n190 B.n121 71.676
R2285 B.n194 B.n122 71.676
R2286 B.n198 B.n123 71.676
R2287 B.n202 B.n124 71.676
R2288 B.n206 B.n125 71.676
R2289 B.n210 B.n126 71.676
R2290 B.n214 B.n127 71.676
R2291 B.n218 B.n128 71.676
R2292 B.n222 B.n129 71.676
R2293 B.n226 B.n130 71.676
R2294 B.n230 B.n131 71.676
R2295 B.n234 B.n132 71.676
R2296 B.n238 B.n133 71.676
R2297 B.n242 B.n134 71.676
R2298 B.n246 B.n135 71.676
R2299 B.n250 B.n136 71.676
R2300 B.n254 B.n137 71.676
R2301 B.n258 B.n138 71.676
R2302 B.n262 B.n139 71.676
R2303 B.n266 B.n140 71.676
R2304 B.n270 B.n141 71.676
R2305 B.n274 B.n142 71.676
R2306 B.n278 B.n143 71.676
R2307 B.n282 B.n144 71.676
R2308 B.n286 B.n145 71.676
R2309 B.n290 B.n146 71.676
R2310 B.n294 B.n147 71.676
R2311 B.n298 B.n148 71.676
R2312 B.n302 B.n149 71.676
R2313 B.n306 B.n150 71.676
R2314 B.n310 B.n151 71.676
R2315 B.n314 B.n152 71.676
R2316 B.n318 B.n153 71.676
R2317 B.n322 B.n154 71.676
R2318 B.n326 B.n155 71.676
R2319 B.n330 B.n156 71.676
R2320 B.n334 B.n157 71.676
R2321 B.n338 B.n158 71.676
R2322 B.n342 B.n159 71.676
R2323 B.n346 B.n160 71.676
R2324 B.n350 B.n161 71.676
R2325 B.n354 B.n162 71.676
R2326 B.n358 B.n163 71.676
R2327 B.n362 B.n164 71.676
R2328 B.n366 B.n165 71.676
R2329 B.n370 B.n166 71.676
R2330 B.n374 B.n167 71.676
R2331 B.n378 B.n168 71.676
R2332 B.n382 B.n169 71.676
R2333 B.n386 B.n170 71.676
R2334 B.n390 B.n171 71.676
R2335 B.n394 B.n172 71.676
R2336 B.n398 B.n173 71.676
R2337 B.n402 B.n174 71.676
R2338 B.n406 B.n175 71.676
R2339 B.n410 B.n176 71.676
R2340 B.n1118 B.n177 71.676
R2341 B.n1118 B.n1117 71.676
R2342 B.n412 B.n176 71.676
R2343 B.n409 B.n175 71.676
R2344 B.n405 B.n174 71.676
R2345 B.n401 B.n173 71.676
R2346 B.n397 B.n172 71.676
R2347 B.n393 B.n171 71.676
R2348 B.n389 B.n170 71.676
R2349 B.n385 B.n169 71.676
R2350 B.n381 B.n168 71.676
R2351 B.n377 B.n167 71.676
R2352 B.n373 B.n166 71.676
R2353 B.n369 B.n165 71.676
R2354 B.n365 B.n164 71.676
R2355 B.n361 B.n163 71.676
R2356 B.n357 B.n162 71.676
R2357 B.n353 B.n161 71.676
R2358 B.n349 B.n160 71.676
R2359 B.n345 B.n159 71.676
R2360 B.n341 B.n158 71.676
R2361 B.n337 B.n157 71.676
R2362 B.n333 B.n156 71.676
R2363 B.n329 B.n155 71.676
R2364 B.n325 B.n154 71.676
R2365 B.n321 B.n153 71.676
R2366 B.n317 B.n152 71.676
R2367 B.n313 B.n151 71.676
R2368 B.n309 B.n150 71.676
R2369 B.n305 B.n149 71.676
R2370 B.n301 B.n148 71.676
R2371 B.n297 B.n147 71.676
R2372 B.n293 B.n146 71.676
R2373 B.n289 B.n145 71.676
R2374 B.n285 B.n144 71.676
R2375 B.n281 B.n143 71.676
R2376 B.n277 B.n142 71.676
R2377 B.n273 B.n141 71.676
R2378 B.n269 B.n140 71.676
R2379 B.n265 B.n139 71.676
R2380 B.n261 B.n138 71.676
R2381 B.n257 B.n137 71.676
R2382 B.n253 B.n136 71.676
R2383 B.n249 B.n135 71.676
R2384 B.n245 B.n134 71.676
R2385 B.n241 B.n133 71.676
R2386 B.n237 B.n132 71.676
R2387 B.n233 B.n131 71.676
R2388 B.n229 B.n130 71.676
R2389 B.n225 B.n129 71.676
R2390 B.n221 B.n128 71.676
R2391 B.n217 B.n127 71.676
R2392 B.n213 B.n126 71.676
R2393 B.n209 B.n125 71.676
R2394 B.n205 B.n124 71.676
R2395 B.n201 B.n123 71.676
R2396 B.n197 B.n122 71.676
R2397 B.n193 B.n121 71.676
R2398 B.n189 B.n120 71.676
R2399 B.n185 B.n119 71.676
R2400 B.n603 B.n539 71.676
R2401 B.n607 B.n606 71.676
R2402 B.n612 B.n611 71.676
R2403 B.n615 B.n614 71.676
R2404 B.n620 B.n619 71.676
R2405 B.n623 B.n622 71.676
R2406 B.n628 B.n627 71.676
R2407 B.n631 B.n630 71.676
R2408 B.n636 B.n635 71.676
R2409 B.n639 B.n638 71.676
R2410 B.n644 B.n643 71.676
R2411 B.n647 B.n646 71.676
R2412 B.n652 B.n651 71.676
R2413 B.n655 B.n654 71.676
R2414 B.n660 B.n659 71.676
R2415 B.n663 B.n662 71.676
R2416 B.n668 B.n667 71.676
R2417 B.n671 B.n670 71.676
R2418 B.n676 B.n675 71.676
R2419 B.n679 B.n678 71.676
R2420 B.n684 B.n683 71.676
R2421 B.n687 B.n686 71.676
R2422 B.n692 B.n691 71.676
R2423 B.n695 B.n694 71.676
R2424 B.n700 B.n699 71.676
R2425 B.n703 B.n702 71.676
R2426 B.n711 B.n710 71.676
R2427 B.n714 B.n713 71.676
R2428 B.n719 B.n718 71.676
R2429 B.n722 B.n721 71.676
R2430 B.n727 B.n726 71.676
R2431 B.n730 B.n729 71.676
R2432 B.n736 B.n735 71.676
R2433 B.n739 B.n738 71.676
R2434 B.n744 B.n743 71.676
R2435 B.n747 B.n746 71.676
R2436 B.n752 B.n751 71.676
R2437 B.n755 B.n754 71.676
R2438 B.n760 B.n759 71.676
R2439 B.n763 B.n762 71.676
R2440 B.n768 B.n767 71.676
R2441 B.n771 B.n770 71.676
R2442 B.n776 B.n775 71.676
R2443 B.n779 B.n778 71.676
R2444 B.n784 B.n783 71.676
R2445 B.n787 B.n786 71.676
R2446 B.n792 B.n791 71.676
R2447 B.n795 B.n794 71.676
R2448 B.n800 B.n799 71.676
R2449 B.n803 B.n802 71.676
R2450 B.n808 B.n807 71.676
R2451 B.n811 B.n810 71.676
R2452 B.n816 B.n815 71.676
R2453 B.n819 B.n818 71.676
R2454 B.n824 B.n823 71.676
R2455 B.n827 B.n826 71.676
R2456 B.n832 B.n831 71.676
R2457 B.n835 B.n834 71.676
R2458 B.n604 B.n603 71.676
R2459 B.n606 B.n600 71.676
R2460 B.n613 B.n612 71.676
R2461 B.n614 B.n598 71.676
R2462 B.n621 B.n620 71.676
R2463 B.n622 B.n596 71.676
R2464 B.n629 B.n628 71.676
R2465 B.n630 B.n594 71.676
R2466 B.n637 B.n636 71.676
R2467 B.n638 B.n592 71.676
R2468 B.n645 B.n644 71.676
R2469 B.n646 B.n590 71.676
R2470 B.n653 B.n652 71.676
R2471 B.n654 B.n588 71.676
R2472 B.n661 B.n660 71.676
R2473 B.n662 B.n586 71.676
R2474 B.n669 B.n668 71.676
R2475 B.n670 B.n584 71.676
R2476 B.n677 B.n676 71.676
R2477 B.n678 B.n582 71.676
R2478 B.n685 B.n684 71.676
R2479 B.n686 B.n580 71.676
R2480 B.n693 B.n692 71.676
R2481 B.n694 B.n578 71.676
R2482 B.n701 B.n700 71.676
R2483 B.n702 B.n576 71.676
R2484 B.n712 B.n711 71.676
R2485 B.n713 B.n574 71.676
R2486 B.n720 B.n719 71.676
R2487 B.n721 B.n572 71.676
R2488 B.n728 B.n727 71.676
R2489 B.n729 B.n568 71.676
R2490 B.n737 B.n736 71.676
R2491 B.n738 B.n566 71.676
R2492 B.n745 B.n744 71.676
R2493 B.n746 B.n564 71.676
R2494 B.n753 B.n752 71.676
R2495 B.n754 B.n562 71.676
R2496 B.n761 B.n760 71.676
R2497 B.n762 B.n560 71.676
R2498 B.n769 B.n768 71.676
R2499 B.n770 B.n558 71.676
R2500 B.n777 B.n776 71.676
R2501 B.n778 B.n556 71.676
R2502 B.n785 B.n784 71.676
R2503 B.n786 B.n554 71.676
R2504 B.n793 B.n792 71.676
R2505 B.n794 B.n552 71.676
R2506 B.n801 B.n800 71.676
R2507 B.n802 B.n550 71.676
R2508 B.n809 B.n808 71.676
R2509 B.n810 B.n548 71.676
R2510 B.n817 B.n816 71.676
R2511 B.n818 B.n546 71.676
R2512 B.n825 B.n824 71.676
R2513 B.n826 B.n544 71.676
R2514 B.n833 B.n832 71.676
R2515 B.n836 B.n835 71.676
R2516 B.n1251 B.n1250 71.676
R2517 B.n1251 B.n2 71.676
R2518 B.n841 B.n540 66.0466
R2519 B.n1120 B.n1119 66.0466
R2520 B.n182 B.n181 62.0611
R2521 B.n179 B.n178 62.0611
R2522 B.n570 B.n569 62.0611
R2523 B.n707 B.n706 62.0611
R2524 B.n183 B.n182 59.5399
R2525 B.n180 B.n179 59.5399
R2526 B.n732 B.n570 59.5399
R2527 B.n708 B.n707 59.5399
R2528 B.n841 B.n536 34.8155
R2529 B.n847 B.n536 34.8155
R2530 B.n847 B.n532 34.8155
R2531 B.n853 B.n532 34.8155
R2532 B.n853 B.n527 34.8155
R2533 B.n859 B.n527 34.8155
R2534 B.n859 B.n528 34.8155
R2535 B.n865 B.n520 34.8155
R2536 B.n871 B.n520 34.8155
R2537 B.n871 B.n516 34.8155
R2538 B.n877 B.n516 34.8155
R2539 B.n877 B.n512 34.8155
R2540 B.n883 B.n512 34.8155
R2541 B.n883 B.n508 34.8155
R2542 B.n889 B.n508 34.8155
R2543 B.n889 B.n504 34.8155
R2544 B.n895 B.n504 34.8155
R2545 B.n895 B.n500 34.8155
R2546 B.n901 B.n500 34.8155
R2547 B.n907 B.n496 34.8155
R2548 B.n907 B.n492 34.8155
R2549 B.n913 B.n492 34.8155
R2550 B.n913 B.n488 34.8155
R2551 B.n919 B.n488 34.8155
R2552 B.n919 B.n484 34.8155
R2553 B.n926 B.n484 34.8155
R2554 B.n926 B.n925 34.8155
R2555 B.n932 B.n477 34.8155
R2556 B.n938 B.n477 34.8155
R2557 B.n938 B.n473 34.8155
R2558 B.n944 B.n473 34.8155
R2559 B.n944 B.n469 34.8155
R2560 B.n950 B.n469 34.8155
R2561 B.n950 B.n464 34.8155
R2562 B.n956 B.n464 34.8155
R2563 B.n956 B.n465 34.8155
R2564 B.n962 B.n457 34.8155
R2565 B.n968 B.n457 34.8155
R2566 B.n968 B.n453 34.8155
R2567 B.n974 B.n453 34.8155
R2568 B.n974 B.n449 34.8155
R2569 B.n980 B.n449 34.8155
R2570 B.n980 B.n445 34.8155
R2571 B.n986 B.n445 34.8155
R2572 B.n992 B.n441 34.8155
R2573 B.n992 B.n437 34.8155
R2574 B.n998 B.n437 34.8155
R2575 B.n998 B.n433 34.8155
R2576 B.n1004 B.n433 34.8155
R2577 B.n1004 B.n429 34.8155
R2578 B.n1010 B.n429 34.8155
R2579 B.n1010 B.n425 34.8155
R2580 B.n1016 B.n425 34.8155
R2581 B.n1023 B.n421 34.8155
R2582 B.n1023 B.n417 34.8155
R2583 B.n1029 B.n417 34.8155
R2584 B.n1029 B.n4 34.8155
R2585 B.n1249 B.n4 34.8155
R2586 B.n1249 B.n1248 34.8155
R2587 B.n1248 B.n1247 34.8155
R2588 B.n1247 B.n8 34.8155
R2589 B.n12 B.n8 34.8155
R2590 B.n1240 B.n12 34.8155
R2591 B.n1240 B.n1239 34.8155
R2592 B.n1238 B.n16 34.8155
R2593 B.n1232 B.n16 34.8155
R2594 B.n1232 B.n1231 34.8155
R2595 B.n1231 B.n1230 34.8155
R2596 B.n1230 B.n23 34.8155
R2597 B.n1224 B.n23 34.8155
R2598 B.n1224 B.n1223 34.8155
R2599 B.n1223 B.n1222 34.8155
R2600 B.n1222 B.n30 34.8155
R2601 B.n1216 B.n1215 34.8155
R2602 B.n1215 B.n1214 34.8155
R2603 B.n1214 B.n37 34.8155
R2604 B.n1208 B.n37 34.8155
R2605 B.n1208 B.n1207 34.8155
R2606 B.n1207 B.n1206 34.8155
R2607 B.n1206 B.n44 34.8155
R2608 B.n1200 B.n44 34.8155
R2609 B.n1199 B.n1198 34.8155
R2610 B.n1198 B.n51 34.8155
R2611 B.n1192 B.n51 34.8155
R2612 B.n1192 B.n1191 34.8155
R2613 B.n1191 B.n1190 34.8155
R2614 B.n1190 B.n58 34.8155
R2615 B.n1184 B.n58 34.8155
R2616 B.n1184 B.n1183 34.8155
R2617 B.n1183 B.n1182 34.8155
R2618 B.n1176 B.n68 34.8155
R2619 B.n1176 B.n1175 34.8155
R2620 B.n1175 B.n1174 34.8155
R2621 B.n1174 B.n72 34.8155
R2622 B.n1168 B.n72 34.8155
R2623 B.n1168 B.n1167 34.8155
R2624 B.n1167 B.n1166 34.8155
R2625 B.n1166 B.n79 34.8155
R2626 B.n1160 B.n1159 34.8155
R2627 B.n1159 B.n1158 34.8155
R2628 B.n1158 B.n86 34.8155
R2629 B.n1152 B.n86 34.8155
R2630 B.n1152 B.n1151 34.8155
R2631 B.n1151 B.n1150 34.8155
R2632 B.n1150 B.n93 34.8155
R2633 B.n1144 B.n93 34.8155
R2634 B.n1144 B.n1143 34.8155
R2635 B.n1143 B.n1142 34.8155
R2636 B.n1142 B.n100 34.8155
R2637 B.n1136 B.n100 34.8155
R2638 B.n1135 B.n1134 34.8155
R2639 B.n1134 B.n107 34.8155
R2640 B.n1128 B.n107 34.8155
R2641 B.n1128 B.n1127 34.8155
R2642 B.n1127 B.n1126 34.8155
R2643 B.n1126 B.n114 34.8155
R2644 B.n1120 B.n114 34.8155
R2645 B.n925 B.t0 33.2795
R2646 B.n68 B.t2 33.2795
R2647 B.n528 B.t18 32.2556
R2648 B.t11 B.n1135 32.2556
R2649 B.n843 B.n538 31.0639
R2650 B.n839 B.n838 31.0639
R2651 B.n1116 B.n1115 31.0639
R2652 B.n1122 B.n116 31.0639
R2653 B.t6 B.n421 28.1597
R2654 B.n1239 B.t7 28.1597
R2655 B.n986 B.t9 27.1357
R2656 B.n1216 B.t4 27.1357
R2657 B.n962 B.t1 22.0159
R2658 B.n1200 B.t5 22.0159
R2659 B.n901 B.t8 18.9439
R2660 B.n1160 B.t3 18.9439
R2661 B B.n1252 18.0485
R2662 B.t8 B.n496 15.872
R2663 B.t3 B.n79 15.872
R2664 B.n465 B.t1 12.8001
R2665 B.t5 B.n1199 12.8001
R2666 B.n844 B.n843 10.6151
R2667 B.n845 B.n844 10.6151
R2668 B.n845 B.n530 10.6151
R2669 B.n855 B.n530 10.6151
R2670 B.n856 B.n855 10.6151
R2671 B.n857 B.n856 10.6151
R2672 B.n857 B.n522 10.6151
R2673 B.n867 B.n522 10.6151
R2674 B.n868 B.n867 10.6151
R2675 B.n869 B.n868 10.6151
R2676 B.n869 B.n514 10.6151
R2677 B.n879 B.n514 10.6151
R2678 B.n880 B.n879 10.6151
R2679 B.n881 B.n880 10.6151
R2680 B.n881 B.n506 10.6151
R2681 B.n891 B.n506 10.6151
R2682 B.n892 B.n891 10.6151
R2683 B.n893 B.n892 10.6151
R2684 B.n893 B.n498 10.6151
R2685 B.n903 B.n498 10.6151
R2686 B.n904 B.n903 10.6151
R2687 B.n905 B.n904 10.6151
R2688 B.n905 B.n490 10.6151
R2689 B.n915 B.n490 10.6151
R2690 B.n916 B.n915 10.6151
R2691 B.n917 B.n916 10.6151
R2692 B.n917 B.n482 10.6151
R2693 B.n928 B.n482 10.6151
R2694 B.n929 B.n928 10.6151
R2695 B.n930 B.n929 10.6151
R2696 B.n930 B.n475 10.6151
R2697 B.n940 B.n475 10.6151
R2698 B.n941 B.n940 10.6151
R2699 B.n942 B.n941 10.6151
R2700 B.n942 B.n467 10.6151
R2701 B.n952 B.n467 10.6151
R2702 B.n953 B.n952 10.6151
R2703 B.n954 B.n953 10.6151
R2704 B.n954 B.n459 10.6151
R2705 B.n964 B.n459 10.6151
R2706 B.n965 B.n964 10.6151
R2707 B.n966 B.n965 10.6151
R2708 B.n966 B.n451 10.6151
R2709 B.n976 B.n451 10.6151
R2710 B.n977 B.n976 10.6151
R2711 B.n978 B.n977 10.6151
R2712 B.n978 B.n443 10.6151
R2713 B.n988 B.n443 10.6151
R2714 B.n989 B.n988 10.6151
R2715 B.n990 B.n989 10.6151
R2716 B.n990 B.n435 10.6151
R2717 B.n1000 B.n435 10.6151
R2718 B.n1001 B.n1000 10.6151
R2719 B.n1002 B.n1001 10.6151
R2720 B.n1002 B.n427 10.6151
R2721 B.n1012 B.n427 10.6151
R2722 B.n1013 B.n1012 10.6151
R2723 B.n1014 B.n1013 10.6151
R2724 B.n1014 B.n419 10.6151
R2725 B.n1025 B.n419 10.6151
R2726 B.n1026 B.n1025 10.6151
R2727 B.n1027 B.n1026 10.6151
R2728 B.n1027 B.n0 10.6151
R2729 B.n602 B.n538 10.6151
R2730 B.n602 B.n601 10.6151
R2731 B.n608 B.n601 10.6151
R2732 B.n609 B.n608 10.6151
R2733 B.n610 B.n609 10.6151
R2734 B.n610 B.n599 10.6151
R2735 B.n616 B.n599 10.6151
R2736 B.n617 B.n616 10.6151
R2737 B.n618 B.n617 10.6151
R2738 B.n618 B.n597 10.6151
R2739 B.n624 B.n597 10.6151
R2740 B.n625 B.n624 10.6151
R2741 B.n626 B.n625 10.6151
R2742 B.n626 B.n595 10.6151
R2743 B.n632 B.n595 10.6151
R2744 B.n633 B.n632 10.6151
R2745 B.n634 B.n633 10.6151
R2746 B.n634 B.n593 10.6151
R2747 B.n640 B.n593 10.6151
R2748 B.n641 B.n640 10.6151
R2749 B.n642 B.n641 10.6151
R2750 B.n642 B.n591 10.6151
R2751 B.n648 B.n591 10.6151
R2752 B.n649 B.n648 10.6151
R2753 B.n650 B.n649 10.6151
R2754 B.n650 B.n589 10.6151
R2755 B.n656 B.n589 10.6151
R2756 B.n657 B.n656 10.6151
R2757 B.n658 B.n657 10.6151
R2758 B.n658 B.n587 10.6151
R2759 B.n664 B.n587 10.6151
R2760 B.n665 B.n664 10.6151
R2761 B.n666 B.n665 10.6151
R2762 B.n666 B.n585 10.6151
R2763 B.n672 B.n585 10.6151
R2764 B.n673 B.n672 10.6151
R2765 B.n674 B.n673 10.6151
R2766 B.n674 B.n583 10.6151
R2767 B.n680 B.n583 10.6151
R2768 B.n681 B.n680 10.6151
R2769 B.n682 B.n681 10.6151
R2770 B.n682 B.n581 10.6151
R2771 B.n688 B.n581 10.6151
R2772 B.n689 B.n688 10.6151
R2773 B.n690 B.n689 10.6151
R2774 B.n690 B.n579 10.6151
R2775 B.n696 B.n579 10.6151
R2776 B.n697 B.n696 10.6151
R2777 B.n698 B.n697 10.6151
R2778 B.n698 B.n577 10.6151
R2779 B.n704 B.n577 10.6151
R2780 B.n705 B.n704 10.6151
R2781 B.n709 B.n705 10.6151
R2782 B.n715 B.n575 10.6151
R2783 B.n716 B.n715 10.6151
R2784 B.n717 B.n716 10.6151
R2785 B.n717 B.n573 10.6151
R2786 B.n723 B.n573 10.6151
R2787 B.n724 B.n723 10.6151
R2788 B.n725 B.n724 10.6151
R2789 B.n725 B.n571 10.6151
R2790 B.n731 B.n571 10.6151
R2791 B.n734 B.n733 10.6151
R2792 B.n734 B.n567 10.6151
R2793 B.n740 B.n567 10.6151
R2794 B.n741 B.n740 10.6151
R2795 B.n742 B.n741 10.6151
R2796 B.n742 B.n565 10.6151
R2797 B.n748 B.n565 10.6151
R2798 B.n749 B.n748 10.6151
R2799 B.n750 B.n749 10.6151
R2800 B.n750 B.n563 10.6151
R2801 B.n756 B.n563 10.6151
R2802 B.n757 B.n756 10.6151
R2803 B.n758 B.n757 10.6151
R2804 B.n758 B.n561 10.6151
R2805 B.n764 B.n561 10.6151
R2806 B.n765 B.n764 10.6151
R2807 B.n766 B.n765 10.6151
R2808 B.n766 B.n559 10.6151
R2809 B.n772 B.n559 10.6151
R2810 B.n773 B.n772 10.6151
R2811 B.n774 B.n773 10.6151
R2812 B.n774 B.n557 10.6151
R2813 B.n780 B.n557 10.6151
R2814 B.n781 B.n780 10.6151
R2815 B.n782 B.n781 10.6151
R2816 B.n782 B.n555 10.6151
R2817 B.n788 B.n555 10.6151
R2818 B.n789 B.n788 10.6151
R2819 B.n790 B.n789 10.6151
R2820 B.n790 B.n553 10.6151
R2821 B.n796 B.n553 10.6151
R2822 B.n797 B.n796 10.6151
R2823 B.n798 B.n797 10.6151
R2824 B.n798 B.n551 10.6151
R2825 B.n804 B.n551 10.6151
R2826 B.n805 B.n804 10.6151
R2827 B.n806 B.n805 10.6151
R2828 B.n806 B.n549 10.6151
R2829 B.n812 B.n549 10.6151
R2830 B.n813 B.n812 10.6151
R2831 B.n814 B.n813 10.6151
R2832 B.n814 B.n547 10.6151
R2833 B.n820 B.n547 10.6151
R2834 B.n821 B.n820 10.6151
R2835 B.n822 B.n821 10.6151
R2836 B.n822 B.n545 10.6151
R2837 B.n828 B.n545 10.6151
R2838 B.n829 B.n828 10.6151
R2839 B.n830 B.n829 10.6151
R2840 B.n830 B.n543 10.6151
R2841 B.n543 B.n542 10.6151
R2842 B.n837 B.n542 10.6151
R2843 B.n838 B.n837 10.6151
R2844 B.n839 B.n534 10.6151
R2845 B.n849 B.n534 10.6151
R2846 B.n850 B.n849 10.6151
R2847 B.n851 B.n850 10.6151
R2848 B.n851 B.n525 10.6151
R2849 B.n861 B.n525 10.6151
R2850 B.n862 B.n861 10.6151
R2851 B.n863 B.n862 10.6151
R2852 B.n863 B.n518 10.6151
R2853 B.n873 B.n518 10.6151
R2854 B.n874 B.n873 10.6151
R2855 B.n875 B.n874 10.6151
R2856 B.n875 B.n510 10.6151
R2857 B.n885 B.n510 10.6151
R2858 B.n886 B.n885 10.6151
R2859 B.n887 B.n886 10.6151
R2860 B.n887 B.n502 10.6151
R2861 B.n897 B.n502 10.6151
R2862 B.n898 B.n897 10.6151
R2863 B.n899 B.n898 10.6151
R2864 B.n899 B.n494 10.6151
R2865 B.n909 B.n494 10.6151
R2866 B.n910 B.n909 10.6151
R2867 B.n911 B.n910 10.6151
R2868 B.n911 B.n486 10.6151
R2869 B.n921 B.n486 10.6151
R2870 B.n922 B.n921 10.6151
R2871 B.n923 B.n922 10.6151
R2872 B.n923 B.n479 10.6151
R2873 B.n934 B.n479 10.6151
R2874 B.n935 B.n934 10.6151
R2875 B.n936 B.n935 10.6151
R2876 B.n936 B.n471 10.6151
R2877 B.n946 B.n471 10.6151
R2878 B.n947 B.n946 10.6151
R2879 B.n948 B.n947 10.6151
R2880 B.n948 B.n462 10.6151
R2881 B.n958 B.n462 10.6151
R2882 B.n959 B.n958 10.6151
R2883 B.n960 B.n959 10.6151
R2884 B.n960 B.n455 10.6151
R2885 B.n970 B.n455 10.6151
R2886 B.n971 B.n970 10.6151
R2887 B.n972 B.n971 10.6151
R2888 B.n972 B.n447 10.6151
R2889 B.n982 B.n447 10.6151
R2890 B.n983 B.n982 10.6151
R2891 B.n984 B.n983 10.6151
R2892 B.n984 B.n439 10.6151
R2893 B.n994 B.n439 10.6151
R2894 B.n995 B.n994 10.6151
R2895 B.n996 B.n995 10.6151
R2896 B.n996 B.n431 10.6151
R2897 B.n1006 B.n431 10.6151
R2898 B.n1007 B.n1006 10.6151
R2899 B.n1008 B.n1007 10.6151
R2900 B.n1008 B.n423 10.6151
R2901 B.n1018 B.n423 10.6151
R2902 B.n1019 B.n1018 10.6151
R2903 B.n1021 B.n1019 10.6151
R2904 B.n1021 B.n1020 10.6151
R2905 B.n1020 B.n415 10.6151
R2906 B.n1032 B.n415 10.6151
R2907 B.n1033 B.n1032 10.6151
R2908 B.n1034 B.n1033 10.6151
R2909 B.n1035 B.n1034 10.6151
R2910 B.n1036 B.n1035 10.6151
R2911 B.n1039 B.n1036 10.6151
R2912 B.n1040 B.n1039 10.6151
R2913 B.n1041 B.n1040 10.6151
R2914 B.n1042 B.n1041 10.6151
R2915 B.n1044 B.n1042 10.6151
R2916 B.n1045 B.n1044 10.6151
R2917 B.n1046 B.n1045 10.6151
R2918 B.n1047 B.n1046 10.6151
R2919 B.n1049 B.n1047 10.6151
R2920 B.n1050 B.n1049 10.6151
R2921 B.n1051 B.n1050 10.6151
R2922 B.n1052 B.n1051 10.6151
R2923 B.n1054 B.n1052 10.6151
R2924 B.n1055 B.n1054 10.6151
R2925 B.n1056 B.n1055 10.6151
R2926 B.n1057 B.n1056 10.6151
R2927 B.n1059 B.n1057 10.6151
R2928 B.n1060 B.n1059 10.6151
R2929 B.n1061 B.n1060 10.6151
R2930 B.n1062 B.n1061 10.6151
R2931 B.n1064 B.n1062 10.6151
R2932 B.n1065 B.n1064 10.6151
R2933 B.n1066 B.n1065 10.6151
R2934 B.n1067 B.n1066 10.6151
R2935 B.n1069 B.n1067 10.6151
R2936 B.n1070 B.n1069 10.6151
R2937 B.n1071 B.n1070 10.6151
R2938 B.n1072 B.n1071 10.6151
R2939 B.n1074 B.n1072 10.6151
R2940 B.n1075 B.n1074 10.6151
R2941 B.n1076 B.n1075 10.6151
R2942 B.n1077 B.n1076 10.6151
R2943 B.n1079 B.n1077 10.6151
R2944 B.n1080 B.n1079 10.6151
R2945 B.n1081 B.n1080 10.6151
R2946 B.n1082 B.n1081 10.6151
R2947 B.n1084 B.n1082 10.6151
R2948 B.n1085 B.n1084 10.6151
R2949 B.n1086 B.n1085 10.6151
R2950 B.n1087 B.n1086 10.6151
R2951 B.n1089 B.n1087 10.6151
R2952 B.n1090 B.n1089 10.6151
R2953 B.n1091 B.n1090 10.6151
R2954 B.n1092 B.n1091 10.6151
R2955 B.n1094 B.n1092 10.6151
R2956 B.n1095 B.n1094 10.6151
R2957 B.n1096 B.n1095 10.6151
R2958 B.n1097 B.n1096 10.6151
R2959 B.n1099 B.n1097 10.6151
R2960 B.n1100 B.n1099 10.6151
R2961 B.n1101 B.n1100 10.6151
R2962 B.n1102 B.n1101 10.6151
R2963 B.n1104 B.n1102 10.6151
R2964 B.n1105 B.n1104 10.6151
R2965 B.n1106 B.n1105 10.6151
R2966 B.n1107 B.n1106 10.6151
R2967 B.n1109 B.n1107 10.6151
R2968 B.n1110 B.n1109 10.6151
R2969 B.n1111 B.n1110 10.6151
R2970 B.n1112 B.n1111 10.6151
R2971 B.n1114 B.n1112 10.6151
R2972 B.n1115 B.n1114 10.6151
R2973 B.n1244 B.n1 10.6151
R2974 B.n1244 B.n1243 10.6151
R2975 B.n1243 B.n1242 10.6151
R2976 B.n1242 B.n10 10.6151
R2977 B.n1236 B.n10 10.6151
R2978 B.n1236 B.n1235 10.6151
R2979 B.n1235 B.n1234 10.6151
R2980 B.n1234 B.n18 10.6151
R2981 B.n1228 B.n18 10.6151
R2982 B.n1228 B.n1227 10.6151
R2983 B.n1227 B.n1226 10.6151
R2984 B.n1226 B.n25 10.6151
R2985 B.n1220 B.n25 10.6151
R2986 B.n1220 B.n1219 10.6151
R2987 B.n1219 B.n1218 10.6151
R2988 B.n1218 B.n32 10.6151
R2989 B.n1212 B.n32 10.6151
R2990 B.n1212 B.n1211 10.6151
R2991 B.n1211 B.n1210 10.6151
R2992 B.n1210 B.n39 10.6151
R2993 B.n1204 B.n39 10.6151
R2994 B.n1204 B.n1203 10.6151
R2995 B.n1203 B.n1202 10.6151
R2996 B.n1202 B.n46 10.6151
R2997 B.n1196 B.n46 10.6151
R2998 B.n1196 B.n1195 10.6151
R2999 B.n1195 B.n1194 10.6151
R3000 B.n1194 B.n53 10.6151
R3001 B.n1188 B.n53 10.6151
R3002 B.n1188 B.n1187 10.6151
R3003 B.n1187 B.n1186 10.6151
R3004 B.n1186 B.n60 10.6151
R3005 B.n1180 B.n60 10.6151
R3006 B.n1180 B.n1179 10.6151
R3007 B.n1179 B.n1178 10.6151
R3008 B.n1178 B.n66 10.6151
R3009 B.n1172 B.n66 10.6151
R3010 B.n1172 B.n1171 10.6151
R3011 B.n1171 B.n1170 10.6151
R3012 B.n1170 B.n74 10.6151
R3013 B.n1164 B.n74 10.6151
R3014 B.n1164 B.n1163 10.6151
R3015 B.n1163 B.n1162 10.6151
R3016 B.n1162 B.n81 10.6151
R3017 B.n1156 B.n81 10.6151
R3018 B.n1156 B.n1155 10.6151
R3019 B.n1155 B.n1154 10.6151
R3020 B.n1154 B.n88 10.6151
R3021 B.n1148 B.n88 10.6151
R3022 B.n1148 B.n1147 10.6151
R3023 B.n1147 B.n1146 10.6151
R3024 B.n1146 B.n95 10.6151
R3025 B.n1140 B.n95 10.6151
R3026 B.n1140 B.n1139 10.6151
R3027 B.n1139 B.n1138 10.6151
R3028 B.n1138 B.n102 10.6151
R3029 B.n1132 B.n102 10.6151
R3030 B.n1132 B.n1131 10.6151
R3031 B.n1131 B.n1130 10.6151
R3032 B.n1130 B.n109 10.6151
R3033 B.n1124 B.n109 10.6151
R3034 B.n1124 B.n1123 10.6151
R3035 B.n1123 B.n1122 10.6151
R3036 B.n184 B.n116 10.6151
R3037 B.n187 B.n184 10.6151
R3038 B.n188 B.n187 10.6151
R3039 B.n191 B.n188 10.6151
R3040 B.n192 B.n191 10.6151
R3041 B.n195 B.n192 10.6151
R3042 B.n196 B.n195 10.6151
R3043 B.n199 B.n196 10.6151
R3044 B.n200 B.n199 10.6151
R3045 B.n203 B.n200 10.6151
R3046 B.n204 B.n203 10.6151
R3047 B.n207 B.n204 10.6151
R3048 B.n208 B.n207 10.6151
R3049 B.n211 B.n208 10.6151
R3050 B.n212 B.n211 10.6151
R3051 B.n215 B.n212 10.6151
R3052 B.n216 B.n215 10.6151
R3053 B.n219 B.n216 10.6151
R3054 B.n220 B.n219 10.6151
R3055 B.n223 B.n220 10.6151
R3056 B.n224 B.n223 10.6151
R3057 B.n227 B.n224 10.6151
R3058 B.n228 B.n227 10.6151
R3059 B.n231 B.n228 10.6151
R3060 B.n232 B.n231 10.6151
R3061 B.n235 B.n232 10.6151
R3062 B.n236 B.n235 10.6151
R3063 B.n239 B.n236 10.6151
R3064 B.n240 B.n239 10.6151
R3065 B.n243 B.n240 10.6151
R3066 B.n244 B.n243 10.6151
R3067 B.n247 B.n244 10.6151
R3068 B.n248 B.n247 10.6151
R3069 B.n251 B.n248 10.6151
R3070 B.n252 B.n251 10.6151
R3071 B.n255 B.n252 10.6151
R3072 B.n256 B.n255 10.6151
R3073 B.n259 B.n256 10.6151
R3074 B.n260 B.n259 10.6151
R3075 B.n263 B.n260 10.6151
R3076 B.n264 B.n263 10.6151
R3077 B.n267 B.n264 10.6151
R3078 B.n268 B.n267 10.6151
R3079 B.n271 B.n268 10.6151
R3080 B.n272 B.n271 10.6151
R3081 B.n275 B.n272 10.6151
R3082 B.n276 B.n275 10.6151
R3083 B.n279 B.n276 10.6151
R3084 B.n280 B.n279 10.6151
R3085 B.n283 B.n280 10.6151
R3086 B.n284 B.n283 10.6151
R3087 B.n287 B.n284 10.6151
R3088 B.n288 B.n287 10.6151
R3089 B.n292 B.n291 10.6151
R3090 B.n295 B.n292 10.6151
R3091 B.n296 B.n295 10.6151
R3092 B.n299 B.n296 10.6151
R3093 B.n300 B.n299 10.6151
R3094 B.n303 B.n300 10.6151
R3095 B.n304 B.n303 10.6151
R3096 B.n307 B.n304 10.6151
R3097 B.n308 B.n307 10.6151
R3098 B.n312 B.n311 10.6151
R3099 B.n315 B.n312 10.6151
R3100 B.n316 B.n315 10.6151
R3101 B.n319 B.n316 10.6151
R3102 B.n320 B.n319 10.6151
R3103 B.n323 B.n320 10.6151
R3104 B.n324 B.n323 10.6151
R3105 B.n327 B.n324 10.6151
R3106 B.n328 B.n327 10.6151
R3107 B.n331 B.n328 10.6151
R3108 B.n332 B.n331 10.6151
R3109 B.n335 B.n332 10.6151
R3110 B.n336 B.n335 10.6151
R3111 B.n339 B.n336 10.6151
R3112 B.n340 B.n339 10.6151
R3113 B.n343 B.n340 10.6151
R3114 B.n344 B.n343 10.6151
R3115 B.n347 B.n344 10.6151
R3116 B.n348 B.n347 10.6151
R3117 B.n351 B.n348 10.6151
R3118 B.n352 B.n351 10.6151
R3119 B.n355 B.n352 10.6151
R3120 B.n356 B.n355 10.6151
R3121 B.n359 B.n356 10.6151
R3122 B.n360 B.n359 10.6151
R3123 B.n363 B.n360 10.6151
R3124 B.n364 B.n363 10.6151
R3125 B.n367 B.n364 10.6151
R3126 B.n368 B.n367 10.6151
R3127 B.n371 B.n368 10.6151
R3128 B.n372 B.n371 10.6151
R3129 B.n375 B.n372 10.6151
R3130 B.n376 B.n375 10.6151
R3131 B.n379 B.n376 10.6151
R3132 B.n380 B.n379 10.6151
R3133 B.n383 B.n380 10.6151
R3134 B.n384 B.n383 10.6151
R3135 B.n387 B.n384 10.6151
R3136 B.n388 B.n387 10.6151
R3137 B.n391 B.n388 10.6151
R3138 B.n392 B.n391 10.6151
R3139 B.n395 B.n392 10.6151
R3140 B.n396 B.n395 10.6151
R3141 B.n399 B.n396 10.6151
R3142 B.n400 B.n399 10.6151
R3143 B.n403 B.n400 10.6151
R3144 B.n404 B.n403 10.6151
R3145 B.n407 B.n404 10.6151
R3146 B.n408 B.n407 10.6151
R3147 B.n411 B.n408 10.6151
R3148 B.n413 B.n411 10.6151
R3149 B.n414 B.n413 10.6151
R3150 B.n1116 B.n414 10.6151
R3151 B.n709 B.n708 9.36635
R3152 B.n733 B.n732 9.36635
R3153 B.n288 B.n183 9.36635
R3154 B.n311 B.n180 9.36635
R3155 B.n1252 B.n0 8.11757
R3156 B.n1252 B.n1 8.11757
R3157 B.t9 B.n441 7.68028
R3158 B.t4 B.n30 7.68028
R3159 B.n1016 B.t6 6.65631
R3160 B.t7 B.n1238 6.65631
R3161 B.n865 B.t18 2.56043
R3162 B.n1136 B.t11 2.56043
R3163 B.n932 B.t0 1.53646
R3164 B.n1182 B.t2 1.53646
R3165 B.n708 B.n575 1.24928
R3166 B.n732 B.n731 1.24928
R3167 B.n291 B.n183 1.24928
R3168 B.n308 B.n180 1.24928
R3169 VN.n11 VN.t8 167.799
R3170 VN.n54 VN.t4 167.799
R3171 VN.n84 VN.n83 161.3
R3172 VN.n82 VN.n44 161.3
R3173 VN.n81 VN.n80 161.3
R3174 VN.n79 VN.n45 161.3
R3175 VN.n78 VN.n77 161.3
R3176 VN.n76 VN.n46 161.3
R3177 VN.n74 VN.n73 161.3
R3178 VN.n72 VN.n47 161.3
R3179 VN.n71 VN.n70 161.3
R3180 VN.n69 VN.n48 161.3
R3181 VN.n68 VN.n67 161.3
R3182 VN.n66 VN.n49 161.3
R3183 VN.n65 VN.n64 161.3
R3184 VN.n63 VN.n50 161.3
R3185 VN.n62 VN.n61 161.3
R3186 VN.n60 VN.n51 161.3
R3187 VN.n59 VN.n58 161.3
R3188 VN.n57 VN.n52 161.3
R3189 VN.n56 VN.n55 161.3
R3190 VN.n41 VN.n40 161.3
R3191 VN.n39 VN.n1 161.3
R3192 VN.n38 VN.n37 161.3
R3193 VN.n36 VN.n2 161.3
R3194 VN.n35 VN.n34 161.3
R3195 VN.n33 VN.n3 161.3
R3196 VN.n31 VN.n30 161.3
R3197 VN.n29 VN.n4 161.3
R3198 VN.n28 VN.n27 161.3
R3199 VN.n26 VN.n5 161.3
R3200 VN.n25 VN.n24 161.3
R3201 VN.n23 VN.n6 161.3
R3202 VN.n22 VN.n21 161.3
R3203 VN.n20 VN.n7 161.3
R3204 VN.n19 VN.n18 161.3
R3205 VN.n17 VN.n8 161.3
R3206 VN.n16 VN.n15 161.3
R3207 VN.n14 VN.n9 161.3
R3208 VN.n13 VN.n12 161.3
R3209 VN.n21 VN.t7 136.119
R3210 VN.n10 VN.t2 136.119
R3211 VN.n32 VN.t3 136.119
R3212 VN.n0 VN.t9 136.119
R3213 VN.n64 VN.t1 136.119
R3214 VN.n53 VN.t6 136.119
R3215 VN.n75 VN.t0 136.119
R3216 VN.n43 VN.t5 136.119
R3217 VN.n42 VN.n0 70.4938
R3218 VN.n85 VN.n43 70.4938
R3219 VN.n11 VN.n10 63.8388
R3220 VN.n54 VN.n53 63.8388
R3221 VN VN.n85 58.0207
R3222 VN.n38 VN.n2 56.5193
R3223 VN.n81 VN.n45 56.5193
R3224 VN.n15 VN.n8 50.2061
R3225 VN.n27 VN.n26 50.2061
R3226 VN.n58 VN.n51 50.2061
R3227 VN.n70 VN.n69 50.2061
R3228 VN.n19 VN.n8 30.7807
R3229 VN.n26 VN.n25 30.7807
R3230 VN.n62 VN.n51 30.7807
R3231 VN.n69 VN.n68 30.7807
R3232 VN.n14 VN.n13 24.4675
R3233 VN.n15 VN.n14 24.4675
R3234 VN.n20 VN.n19 24.4675
R3235 VN.n21 VN.n20 24.4675
R3236 VN.n21 VN.n6 24.4675
R3237 VN.n25 VN.n6 24.4675
R3238 VN.n27 VN.n4 24.4675
R3239 VN.n31 VN.n4 24.4675
R3240 VN.n34 VN.n33 24.4675
R3241 VN.n34 VN.n2 24.4675
R3242 VN.n39 VN.n38 24.4675
R3243 VN.n40 VN.n39 24.4675
R3244 VN.n58 VN.n57 24.4675
R3245 VN.n57 VN.n56 24.4675
R3246 VN.n68 VN.n49 24.4675
R3247 VN.n64 VN.n49 24.4675
R3248 VN.n64 VN.n63 24.4675
R3249 VN.n63 VN.n62 24.4675
R3250 VN.n77 VN.n45 24.4675
R3251 VN.n77 VN.n76 24.4675
R3252 VN.n74 VN.n47 24.4675
R3253 VN.n70 VN.n47 24.4675
R3254 VN.n83 VN.n82 24.4675
R3255 VN.n82 VN.n81 24.4675
R3256 VN.n40 VN.n0 19.5741
R3257 VN.n83 VN.n43 19.5741
R3258 VN.n33 VN.n32 14.6807
R3259 VN.n76 VN.n75 14.6807
R3260 VN.n13 VN.n10 9.7873
R3261 VN.n32 VN.n31 9.7873
R3262 VN.n56 VN.n53 9.7873
R3263 VN.n75 VN.n74 9.7873
R3264 VN.n55 VN.n54 5.5843
R3265 VN.n12 VN.n11 5.5843
R3266 VN.n85 VN.n84 0.354971
R3267 VN.n42 VN.n41 0.354971
R3268 VN VN.n42 0.26696
R3269 VN.n84 VN.n44 0.189894
R3270 VN.n80 VN.n44 0.189894
R3271 VN.n80 VN.n79 0.189894
R3272 VN.n79 VN.n78 0.189894
R3273 VN.n78 VN.n46 0.189894
R3274 VN.n73 VN.n46 0.189894
R3275 VN.n73 VN.n72 0.189894
R3276 VN.n72 VN.n71 0.189894
R3277 VN.n71 VN.n48 0.189894
R3278 VN.n67 VN.n48 0.189894
R3279 VN.n67 VN.n66 0.189894
R3280 VN.n66 VN.n65 0.189894
R3281 VN.n65 VN.n50 0.189894
R3282 VN.n61 VN.n50 0.189894
R3283 VN.n61 VN.n60 0.189894
R3284 VN.n60 VN.n59 0.189894
R3285 VN.n59 VN.n52 0.189894
R3286 VN.n55 VN.n52 0.189894
R3287 VN.n12 VN.n9 0.189894
R3288 VN.n16 VN.n9 0.189894
R3289 VN.n17 VN.n16 0.189894
R3290 VN.n18 VN.n17 0.189894
R3291 VN.n18 VN.n7 0.189894
R3292 VN.n22 VN.n7 0.189894
R3293 VN.n23 VN.n22 0.189894
R3294 VN.n24 VN.n23 0.189894
R3295 VN.n24 VN.n5 0.189894
R3296 VN.n28 VN.n5 0.189894
R3297 VN.n29 VN.n28 0.189894
R3298 VN.n30 VN.n29 0.189894
R3299 VN.n30 VN.n3 0.189894
R3300 VN.n35 VN.n3 0.189894
R3301 VN.n36 VN.n35 0.189894
R3302 VN.n37 VN.n36 0.189894
R3303 VN.n37 VN.n1 0.189894
R3304 VN.n41 VN.n1 0.189894
R3305 VDD2.n177 VDD2.n93 289.615
R3306 VDD2.n84 VDD2.n0 289.615
R3307 VDD2.n178 VDD2.n177 185
R3308 VDD2.n176 VDD2.n175 185
R3309 VDD2.n97 VDD2.n96 185
R3310 VDD2.n170 VDD2.n169 185
R3311 VDD2.n168 VDD2.n99 185
R3312 VDD2.n167 VDD2.n166 185
R3313 VDD2.n102 VDD2.n100 185
R3314 VDD2.n161 VDD2.n160 185
R3315 VDD2.n159 VDD2.n158 185
R3316 VDD2.n106 VDD2.n105 185
R3317 VDD2.n153 VDD2.n152 185
R3318 VDD2.n151 VDD2.n150 185
R3319 VDD2.n110 VDD2.n109 185
R3320 VDD2.n145 VDD2.n144 185
R3321 VDD2.n143 VDD2.n142 185
R3322 VDD2.n114 VDD2.n113 185
R3323 VDD2.n137 VDD2.n136 185
R3324 VDD2.n135 VDD2.n134 185
R3325 VDD2.n118 VDD2.n117 185
R3326 VDD2.n129 VDD2.n128 185
R3327 VDD2.n127 VDD2.n126 185
R3328 VDD2.n122 VDD2.n121 185
R3329 VDD2.n28 VDD2.n27 185
R3330 VDD2.n33 VDD2.n32 185
R3331 VDD2.n35 VDD2.n34 185
R3332 VDD2.n24 VDD2.n23 185
R3333 VDD2.n41 VDD2.n40 185
R3334 VDD2.n43 VDD2.n42 185
R3335 VDD2.n20 VDD2.n19 185
R3336 VDD2.n49 VDD2.n48 185
R3337 VDD2.n51 VDD2.n50 185
R3338 VDD2.n16 VDD2.n15 185
R3339 VDD2.n57 VDD2.n56 185
R3340 VDD2.n59 VDD2.n58 185
R3341 VDD2.n12 VDD2.n11 185
R3342 VDD2.n65 VDD2.n64 185
R3343 VDD2.n67 VDD2.n66 185
R3344 VDD2.n8 VDD2.n7 185
R3345 VDD2.n74 VDD2.n73 185
R3346 VDD2.n75 VDD2.n6 185
R3347 VDD2.n77 VDD2.n76 185
R3348 VDD2.n4 VDD2.n3 185
R3349 VDD2.n83 VDD2.n82 185
R3350 VDD2.n85 VDD2.n84 185
R3351 VDD2.n123 VDD2.t4 147.659
R3352 VDD2.n29 VDD2.t1 147.659
R3353 VDD2.n177 VDD2.n176 104.615
R3354 VDD2.n176 VDD2.n96 104.615
R3355 VDD2.n169 VDD2.n96 104.615
R3356 VDD2.n169 VDD2.n168 104.615
R3357 VDD2.n168 VDD2.n167 104.615
R3358 VDD2.n167 VDD2.n100 104.615
R3359 VDD2.n160 VDD2.n100 104.615
R3360 VDD2.n160 VDD2.n159 104.615
R3361 VDD2.n159 VDD2.n105 104.615
R3362 VDD2.n152 VDD2.n105 104.615
R3363 VDD2.n152 VDD2.n151 104.615
R3364 VDD2.n151 VDD2.n109 104.615
R3365 VDD2.n144 VDD2.n109 104.615
R3366 VDD2.n144 VDD2.n143 104.615
R3367 VDD2.n143 VDD2.n113 104.615
R3368 VDD2.n136 VDD2.n113 104.615
R3369 VDD2.n136 VDD2.n135 104.615
R3370 VDD2.n135 VDD2.n117 104.615
R3371 VDD2.n128 VDD2.n117 104.615
R3372 VDD2.n128 VDD2.n127 104.615
R3373 VDD2.n127 VDD2.n121 104.615
R3374 VDD2.n33 VDD2.n27 104.615
R3375 VDD2.n34 VDD2.n33 104.615
R3376 VDD2.n34 VDD2.n23 104.615
R3377 VDD2.n41 VDD2.n23 104.615
R3378 VDD2.n42 VDD2.n41 104.615
R3379 VDD2.n42 VDD2.n19 104.615
R3380 VDD2.n49 VDD2.n19 104.615
R3381 VDD2.n50 VDD2.n49 104.615
R3382 VDD2.n50 VDD2.n15 104.615
R3383 VDD2.n57 VDD2.n15 104.615
R3384 VDD2.n58 VDD2.n57 104.615
R3385 VDD2.n58 VDD2.n11 104.615
R3386 VDD2.n65 VDD2.n11 104.615
R3387 VDD2.n66 VDD2.n65 104.615
R3388 VDD2.n66 VDD2.n7 104.615
R3389 VDD2.n74 VDD2.n7 104.615
R3390 VDD2.n75 VDD2.n74 104.615
R3391 VDD2.n76 VDD2.n75 104.615
R3392 VDD2.n76 VDD2.n3 104.615
R3393 VDD2.n83 VDD2.n3 104.615
R3394 VDD2.n84 VDD2.n83 104.615
R3395 VDD2.n92 VDD2.n91 65.3124
R3396 VDD2 VDD2.n185 65.3095
R3397 VDD2.n184 VDD2.n183 63.2989
R3398 VDD2.n90 VDD2.n89 63.2988
R3399 VDD2.n90 VDD2.n88 54.144
R3400 VDD2.t4 VDD2.n121 52.3082
R3401 VDD2.t1 VDD2.n27 52.3082
R3402 VDD2.n182 VDD2.n181 51.3853
R3403 VDD2.n182 VDD2.n92 50.7929
R3404 VDD2.n123 VDD2.n122 15.6677
R3405 VDD2.n29 VDD2.n28 15.6677
R3406 VDD2.n170 VDD2.n99 13.1884
R3407 VDD2.n77 VDD2.n6 13.1884
R3408 VDD2.n171 VDD2.n97 12.8005
R3409 VDD2.n166 VDD2.n101 12.8005
R3410 VDD2.n126 VDD2.n125 12.8005
R3411 VDD2.n32 VDD2.n31 12.8005
R3412 VDD2.n73 VDD2.n72 12.8005
R3413 VDD2.n78 VDD2.n4 12.8005
R3414 VDD2.n175 VDD2.n174 12.0247
R3415 VDD2.n165 VDD2.n102 12.0247
R3416 VDD2.n129 VDD2.n120 12.0247
R3417 VDD2.n35 VDD2.n26 12.0247
R3418 VDD2.n71 VDD2.n8 12.0247
R3419 VDD2.n82 VDD2.n81 12.0247
R3420 VDD2.n178 VDD2.n95 11.249
R3421 VDD2.n162 VDD2.n161 11.249
R3422 VDD2.n130 VDD2.n118 11.249
R3423 VDD2.n36 VDD2.n24 11.249
R3424 VDD2.n68 VDD2.n67 11.249
R3425 VDD2.n85 VDD2.n2 11.249
R3426 VDD2.n179 VDD2.n93 10.4732
R3427 VDD2.n158 VDD2.n104 10.4732
R3428 VDD2.n134 VDD2.n133 10.4732
R3429 VDD2.n40 VDD2.n39 10.4732
R3430 VDD2.n64 VDD2.n10 10.4732
R3431 VDD2.n86 VDD2.n0 10.4732
R3432 VDD2.n157 VDD2.n106 9.69747
R3433 VDD2.n137 VDD2.n116 9.69747
R3434 VDD2.n43 VDD2.n22 9.69747
R3435 VDD2.n63 VDD2.n12 9.69747
R3436 VDD2.n181 VDD2.n180 9.45567
R3437 VDD2.n88 VDD2.n87 9.45567
R3438 VDD2.n149 VDD2.n148 9.3005
R3439 VDD2.n108 VDD2.n107 9.3005
R3440 VDD2.n155 VDD2.n154 9.3005
R3441 VDD2.n157 VDD2.n156 9.3005
R3442 VDD2.n104 VDD2.n103 9.3005
R3443 VDD2.n163 VDD2.n162 9.3005
R3444 VDD2.n165 VDD2.n164 9.3005
R3445 VDD2.n101 VDD2.n98 9.3005
R3446 VDD2.n180 VDD2.n179 9.3005
R3447 VDD2.n95 VDD2.n94 9.3005
R3448 VDD2.n174 VDD2.n173 9.3005
R3449 VDD2.n172 VDD2.n171 9.3005
R3450 VDD2.n147 VDD2.n146 9.3005
R3451 VDD2.n112 VDD2.n111 9.3005
R3452 VDD2.n141 VDD2.n140 9.3005
R3453 VDD2.n139 VDD2.n138 9.3005
R3454 VDD2.n116 VDD2.n115 9.3005
R3455 VDD2.n133 VDD2.n132 9.3005
R3456 VDD2.n131 VDD2.n130 9.3005
R3457 VDD2.n120 VDD2.n119 9.3005
R3458 VDD2.n125 VDD2.n124 9.3005
R3459 VDD2.n87 VDD2.n86 9.3005
R3460 VDD2.n2 VDD2.n1 9.3005
R3461 VDD2.n81 VDD2.n80 9.3005
R3462 VDD2.n79 VDD2.n78 9.3005
R3463 VDD2.n18 VDD2.n17 9.3005
R3464 VDD2.n47 VDD2.n46 9.3005
R3465 VDD2.n45 VDD2.n44 9.3005
R3466 VDD2.n22 VDD2.n21 9.3005
R3467 VDD2.n39 VDD2.n38 9.3005
R3468 VDD2.n37 VDD2.n36 9.3005
R3469 VDD2.n26 VDD2.n25 9.3005
R3470 VDD2.n31 VDD2.n30 9.3005
R3471 VDD2.n53 VDD2.n52 9.3005
R3472 VDD2.n55 VDD2.n54 9.3005
R3473 VDD2.n14 VDD2.n13 9.3005
R3474 VDD2.n61 VDD2.n60 9.3005
R3475 VDD2.n63 VDD2.n62 9.3005
R3476 VDD2.n10 VDD2.n9 9.3005
R3477 VDD2.n69 VDD2.n68 9.3005
R3478 VDD2.n71 VDD2.n70 9.3005
R3479 VDD2.n72 VDD2.n5 9.3005
R3480 VDD2.n154 VDD2.n153 8.92171
R3481 VDD2.n138 VDD2.n114 8.92171
R3482 VDD2.n44 VDD2.n20 8.92171
R3483 VDD2.n60 VDD2.n59 8.92171
R3484 VDD2.n150 VDD2.n108 8.14595
R3485 VDD2.n142 VDD2.n141 8.14595
R3486 VDD2.n48 VDD2.n47 8.14595
R3487 VDD2.n56 VDD2.n14 8.14595
R3488 VDD2.n149 VDD2.n110 7.3702
R3489 VDD2.n145 VDD2.n112 7.3702
R3490 VDD2.n51 VDD2.n18 7.3702
R3491 VDD2.n55 VDD2.n16 7.3702
R3492 VDD2.n146 VDD2.n110 6.59444
R3493 VDD2.n146 VDD2.n145 6.59444
R3494 VDD2.n52 VDD2.n51 6.59444
R3495 VDD2.n52 VDD2.n16 6.59444
R3496 VDD2.n150 VDD2.n149 5.81868
R3497 VDD2.n142 VDD2.n112 5.81868
R3498 VDD2.n48 VDD2.n18 5.81868
R3499 VDD2.n56 VDD2.n55 5.81868
R3500 VDD2.n153 VDD2.n108 5.04292
R3501 VDD2.n141 VDD2.n114 5.04292
R3502 VDD2.n47 VDD2.n20 5.04292
R3503 VDD2.n59 VDD2.n14 5.04292
R3504 VDD2.n124 VDD2.n123 4.38563
R3505 VDD2.n30 VDD2.n29 4.38563
R3506 VDD2.n154 VDD2.n106 4.26717
R3507 VDD2.n138 VDD2.n137 4.26717
R3508 VDD2.n44 VDD2.n43 4.26717
R3509 VDD2.n60 VDD2.n12 4.26717
R3510 VDD2.n181 VDD2.n93 3.49141
R3511 VDD2.n158 VDD2.n157 3.49141
R3512 VDD2.n134 VDD2.n116 3.49141
R3513 VDD2.n40 VDD2.n22 3.49141
R3514 VDD2.n64 VDD2.n63 3.49141
R3515 VDD2.n88 VDD2.n0 3.49141
R3516 VDD2.n184 VDD2.n182 2.75912
R3517 VDD2.n179 VDD2.n178 2.71565
R3518 VDD2.n161 VDD2.n104 2.71565
R3519 VDD2.n133 VDD2.n118 2.71565
R3520 VDD2.n39 VDD2.n24 2.71565
R3521 VDD2.n67 VDD2.n10 2.71565
R3522 VDD2.n86 VDD2.n85 2.71565
R3523 VDD2.n175 VDD2.n95 1.93989
R3524 VDD2.n162 VDD2.n102 1.93989
R3525 VDD2.n130 VDD2.n129 1.93989
R3526 VDD2.n36 VDD2.n35 1.93989
R3527 VDD2.n68 VDD2.n8 1.93989
R3528 VDD2.n82 VDD2.n2 1.93989
R3529 VDD2.n185 VDD2.t3 1.22197
R3530 VDD2.n185 VDD2.t5 1.22197
R3531 VDD2.n183 VDD2.t9 1.22197
R3532 VDD2.n183 VDD2.t8 1.22197
R3533 VDD2.n91 VDD2.t6 1.22197
R3534 VDD2.n91 VDD2.t0 1.22197
R3535 VDD2.n89 VDD2.t7 1.22197
R3536 VDD2.n89 VDD2.t2 1.22197
R3537 VDD2.n174 VDD2.n97 1.16414
R3538 VDD2.n166 VDD2.n165 1.16414
R3539 VDD2.n126 VDD2.n120 1.16414
R3540 VDD2.n32 VDD2.n26 1.16414
R3541 VDD2.n73 VDD2.n71 1.16414
R3542 VDD2.n81 VDD2.n4 1.16414
R3543 VDD2 VDD2.n184 0.748345
R3544 VDD2.n92 VDD2.n90 0.634809
R3545 VDD2.n171 VDD2.n170 0.388379
R3546 VDD2.n101 VDD2.n99 0.388379
R3547 VDD2.n125 VDD2.n122 0.388379
R3548 VDD2.n31 VDD2.n28 0.388379
R3549 VDD2.n72 VDD2.n6 0.388379
R3550 VDD2.n78 VDD2.n77 0.388379
R3551 VDD2.n180 VDD2.n94 0.155672
R3552 VDD2.n173 VDD2.n94 0.155672
R3553 VDD2.n173 VDD2.n172 0.155672
R3554 VDD2.n172 VDD2.n98 0.155672
R3555 VDD2.n164 VDD2.n98 0.155672
R3556 VDD2.n164 VDD2.n163 0.155672
R3557 VDD2.n163 VDD2.n103 0.155672
R3558 VDD2.n156 VDD2.n103 0.155672
R3559 VDD2.n156 VDD2.n155 0.155672
R3560 VDD2.n155 VDD2.n107 0.155672
R3561 VDD2.n148 VDD2.n107 0.155672
R3562 VDD2.n148 VDD2.n147 0.155672
R3563 VDD2.n147 VDD2.n111 0.155672
R3564 VDD2.n140 VDD2.n111 0.155672
R3565 VDD2.n140 VDD2.n139 0.155672
R3566 VDD2.n139 VDD2.n115 0.155672
R3567 VDD2.n132 VDD2.n115 0.155672
R3568 VDD2.n132 VDD2.n131 0.155672
R3569 VDD2.n131 VDD2.n119 0.155672
R3570 VDD2.n124 VDD2.n119 0.155672
R3571 VDD2.n30 VDD2.n25 0.155672
R3572 VDD2.n37 VDD2.n25 0.155672
R3573 VDD2.n38 VDD2.n37 0.155672
R3574 VDD2.n38 VDD2.n21 0.155672
R3575 VDD2.n45 VDD2.n21 0.155672
R3576 VDD2.n46 VDD2.n45 0.155672
R3577 VDD2.n46 VDD2.n17 0.155672
R3578 VDD2.n53 VDD2.n17 0.155672
R3579 VDD2.n54 VDD2.n53 0.155672
R3580 VDD2.n54 VDD2.n13 0.155672
R3581 VDD2.n61 VDD2.n13 0.155672
R3582 VDD2.n62 VDD2.n61 0.155672
R3583 VDD2.n62 VDD2.n9 0.155672
R3584 VDD2.n69 VDD2.n9 0.155672
R3585 VDD2.n70 VDD2.n69 0.155672
R3586 VDD2.n70 VDD2.n5 0.155672
R3587 VDD2.n79 VDD2.n5 0.155672
R3588 VDD2.n80 VDD2.n79 0.155672
R3589 VDD2.n80 VDD2.n1 0.155672
R3590 VDD2.n87 VDD2.n1 0.155672
C0 VTAIL VN 15.0698f
C1 VDD1 VP 14.960401f
C2 VDD2 VN 14.500599f
C3 VDD1 VN 0.154017f
C4 VP VN 9.580719f
C5 VTAIL VDD2 12.373199f
C6 VTAIL VDD1 12.321099f
C7 VDD1 VDD2 2.35094f
C8 VTAIL VP 15.0841f
C9 VDD2 VP 0.618373f
C10 VDD2 B 8.261911f
C11 VDD1 B 8.240893f
C12 VTAIL B 10.113239f
C13 VN B 19.783161f
C14 VP B 18.274967f
C15 VDD2.n0 B 0.033611f
C16 VDD2.n1 B 0.023798f
C17 VDD2.n2 B 0.012788f
C18 VDD2.n3 B 0.030226f
C19 VDD2.n4 B 0.01354f
C20 VDD2.n5 B 0.023798f
C21 VDD2.n6 B 0.013164f
C22 VDD2.n7 B 0.030226f
C23 VDD2.n8 B 0.01354f
C24 VDD2.n9 B 0.023798f
C25 VDD2.n10 B 0.012788f
C26 VDD2.n11 B 0.030226f
C27 VDD2.n12 B 0.01354f
C28 VDD2.n13 B 0.023798f
C29 VDD2.n14 B 0.012788f
C30 VDD2.n15 B 0.030226f
C31 VDD2.n16 B 0.01354f
C32 VDD2.n17 B 0.023798f
C33 VDD2.n18 B 0.012788f
C34 VDD2.n19 B 0.030226f
C35 VDD2.n20 B 0.01354f
C36 VDD2.n21 B 0.023798f
C37 VDD2.n22 B 0.012788f
C38 VDD2.n23 B 0.030226f
C39 VDD2.n24 B 0.01354f
C40 VDD2.n25 B 0.023798f
C41 VDD2.n26 B 0.012788f
C42 VDD2.n27 B 0.02267f
C43 VDD2.n28 B 0.017855f
C44 VDD2.t1 B 0.049938f
C45 VDD2.n29 B 0.162435f
C46 VDD2.n30 B 1.6803f
C47 VDD2.n31 B 0.012788f
C48 VDD2.n32 B 0.01354f
C49 VDD2.n33 B 0.030226f
C50 VDD2.n34 B 0.030226f
C51 VDD2.n35 B 0.01354f
C52 VDD2.n36 B 0.012788f
C53 VDD2.n37 B 0.023798f
C54 VDD2.n38 B 0.023798f
C55 VDD2.n39 B 0.012788f
C56 VDD2.n40 B 0.01354f
C57 VDD2.n41 B 0.030226f
C58 VDD2.n42 B 0.030226f
C59 VDD2.n43 B 0.01354f
C60 VDD2.n44 B 0.012788f
C61 VDD2.n45 B 0.023798f
C62 VDD2.n46 B 0.023798f
C63 VDD2.n47 B 0.012788f
C64 VDD2.n48 B 0.01354f
C65 VDD2.n49 B 0.030226f
C66 VDD2.n50 B 0.030226f
C67 VDD2.n51 B 0.01354f
C68 VDD2.n52 B 0.012788f
C69 VDD2.n53 B 0.023798f
C70 VDD2.n54 B 0.023798f
C71 VDD2.n55 B 0.012788f
C72 VDD2.n56 B 0.01354f
C73 VDD2.n57 B 0.030226f
C74 VDD2.n58 B 0.030226f
C75 VDD2.n59 B 0.01354f
C76 VDD2.n60 B 0.012788f
C77 VDD2.n61 B 0.023798f
C78 VDD2.n62 B 0.023798f
C79 VDD2.n63 B 0.012788f
C80 VDD2.n64 B 0.01354f
C81 VDD2.n65 B 0.030226f
C82 VDD2.n66 B 0.030226f
C83 VDD2.n67 B 0.01354f
C84 VDD2.n68 B 0.012788f
C85 VDD2.n69 B 0.023798f
C86 VDD2.n70 B 0.023798f
C87 VDD2.n71 B 0.012788f
C88 VDD2.n72 B 0.012788f
C89 VDD2.n73 B 0.01354f
C90 VDD2.n74 B 0.030226f
C91 VDD2.n75 B 0.030226f
C92 VDD2.n76 B 0.030226f
C93 VDD2.n77 B 0.013164f
C94 VDD2.n78 B 0.012788f
C95 VDD2.n79 B 0.023798f
C96 VDD2.n80 B 0.023798f
C97 VDD2.n81 B 0.012788f
C98 VDD2.n82 B 0.01354f
C99 VDD2.n83 B 0.030226f
C100 VDD2.n84 B 0.065719f
C101 VDD2.n85 B 0.01354f
C102 VDD2.n86 B 0.012788f
C103 VDD2.n87 B 0.059234f
C104 VDD2.n88 B 0.066564f
C105 VDD2.t7 B 0.304843f
C106 VDD2.t2 B 0.304843f
C107 VDD2.n89 B 2.7677f
C108 VDD2.n90 B 0.701076f
C109 VDD2.t6 B 0.304843f
C110 VDD2.t0 B 0.304843f
C111 VDD2.n91 B 2.78526f
C112 VDD2.n92 B 3.14823f
C113 VDD2.n93 B 0.033611f
C114 VDD2.n94 B 0.023798f
C115 VDD2.n95 B 0.012788f
C116 VDD2.n96 B 0.030226f
C117 VDD2.n97 B 0.01354f
C118 VDD2.n98 B 0.023798f
C119 VDD2.n99 B 0.013164f
C120 VDD2.n100 B 0.030226f
C121 VDD2.n101 B 0.012788f
C122 VDD2.n102 B 0.01354f
C123 VDD2.n103 B 0.023798f
C124 VDD2.n104 B 0.012788f
C125 VDD2.n105 B 0.030226f
C126 VDD2.n106 B 0.01354f
C127 VDD2.n107 B 0.023798f
C128 VDD2.n108 B 0.012788f
C129 VDD2.n109 B 0.030226f
C130 VDD2.n110 B 0.01354f
C131 VDD2.n111 B 0.023798f
C132 VDD2.n112 B 0.012788f
C133 VDD2.n113 B 0.030226f
C134 VDD2.n114 B 0.01354f
C135 VDD2.n115 B 0.023798f
C136 VDD2.n116 B 0.012788f
C137 VDD2.n117 B 0.030226f
C138 VDD2.n118 B 0.01354f
C139 VDD2.n119 B 0.023798f
C140 VDD2.n120 B 0.012788f
C141 VDD2.n121 B 0.02267f
C142 VDD2.n122 B 0.017855f
C143 VDD2.t4 B 0.049938f
C144 VDD2.n123 B 0.162435f
C145 VDD2.n124 B 1.6803f
C146 VDD2.n125 B 0.012788f
C147 VDD2.n126 B 0.01354f
C148 VDD2.n127 B 0.030226f
C149 VDD2.n128 B 0.030226f
C150 VDD2.n129 B 0.01354f
C151 VDD2.n130 B 0.012788f
C152 VDD2.n131 B 0.023798f
C153 VDD2.n132 B 0.023798f
C154 VDD2.n133 B 0.012788f
C155 VDD2.n134 B 0.01354f
C156 VDD2.n135 B 0.030226f
C157 VDD2.n136 B 0.030226f
C158 VDD2.n137 B 0.01354f
C159 VDD2.n138 B 0.012788f
C160 VDD2.n139 B 0.023798f
C161 VDD2.n140 B 0.023798f
C162 VDD2.n141 B 0.012788f
C163 VDD2.n142 B 0.01354f
C164 VDD2.n143 B 0.030226f
C165 VDD2.n144 B 0.030226f
C166 VDD2.n145 B 0.01354f
C167 VDD2.n146 B 0.012788f
C168 VDD2.n147 B 0.023798f
C169 VDD2.n148 B 0.023798f
C170 VDD2.n149 B 0.012788f
C171 VDD2.n150 B 0.01354f
C172 VDD2.n151 B 0.030226f
C173 VDD2.n152 B 0.030226f
C174 VDD2.n153 B 0.01354f
C175 VDD2.n154 B 0.012788f
C176 VDD2.n155 B 0.023798f
C177 VDD2.n156 B 0.023798f
C178 VDD2.n157 B 0.012788f
C179 VDD2.n158 B 0.01354f
C180 VDD2.n159 B 0.030226f
C181 VDD2.n160 B 0.030226f
C182 VDD2.n161 B 0.01354f
C183 VDD2.n162 B 0.012788f
C184 VDD2.n163 B 0.023798f
C185 VDD2.n164 B 0.023798f
C186 VDD2.n165 B 0.012788f
C187 VDD2.n166 B 0.01354f
C188 VDD2.n167 B 0.030226f
C189 VDD2.n168 B 0.030226f
C190 VDD2.n169 B 0.030226f
C191 VDD2.n170 B 0.013164f
C192 VDD2.n171 B 0.012788f
C193 VDD2.n172 B 0.023798f
C194 VDD2.n173 B 0.023798f
C195 VDD2.n174 B 0.012788f
C196 VDD2.n175 B 0.01354f
C197 VDD2.n176 B 0.030226f
C198 VDD2.n177 B 0.065719f
C199 VDD2.n178 B 0.01354f
C200 VDD2.n179 B 0.012788f
C201 VDD2.n180 B 0.059234f
C202 VDD2.n181 B 0.053328f
C203 VDD2.n182 B 3.15981f
C204 VDD2.t9 B 0.304843f
C205 VDD2.t8 B 0.304843f
C206 VDD2.n183 B 2.76771f
C207 VDD2.n184 B 0.462357f
C208 VDD2.t3 B 0.304843f
C209 VDD2.t5 B 0.304843f
C210 VDD2.n185 B 2.78522f
C211 VN.t9 B 2.48159f
C212 VN.n0 B 0.935725f
C213 VN.n1 B 0.019433f
C214 VN.n2 B 0.031077f
C215 VN.n3 B 0.019433f
C216 VN.t3 B 2.48159f
C217 VN.n4 B 0.036219f
C218 VN.n5 B 0.019433f
C219 VN.n6 B 0.036219f
C220 VN.n7 B 0.019433f
C221 VN.t7 B 2.48159f
C222 VN.n8 B 0.018358f
C223 VN.n9 B 0.019433f
C224 VN.t2 B 2.48159f
C225 VN.n10 B 0.920924f
C226 VN.t8 B 2.66818f
C227 VN.n11 B 0.897724f
C228 VN.n12 B 0.207347f
C229 VN.n13 B 0.02549f
C230 VN.n14 B 0.036219f
C231 VN.n15 B 0.035667f
C232 VN.n16 B 0.019433f
C233 VN.n17 B 0.019433f
C234 VN.n18 B 0.019433f
C235 VN.n19 B 0.038932f
C236 VN.n20 B 0.036219f
C237 VN.n21 B 0.880783f
C238 VN.n22 B 0.019433f
C239 VN.n23 B 0.019433f
C240 VN.n24 B 0.019433f
C241 VN.n25 B 0.038932f
C242 VN.n26 B 0.018358f
C243 VN.n27 B 0.035667f
C244 VN.n28 B 0.019433f
C245 VN.n29 B 0.019433f
C246 VN.n30 B 0.019433f
C247 VN.n31 B 0.02549f
C248 VN.n32 B 0.862446f
C249 VN.n33 B 0.029066f
C250 VN.n34 B 0.036219f
C251 VN.n35 B 0.019433f
C252 VN.n36 B 0.019433f
C253 VN.n37 B 0.019433f
C254 VN.n38 B 0.025662f
C255 VN.n39 B 0.036219f
C256 VN.n40 B 0.032643f
C257 VN.n41 B 0.031365f
C258 VN.n42 B 0.039968f
C259 VN.t5 B 2.48159f
C260 VN.n43 B 0.935725f
C261 VN.n44 B 0.019433f
C262 VN.n45 B 0.031077f
C263 VN.n46 B 0.019433f
C264 VN.t0 B 2.48159f
C265 VN.n47 B 0.036219f
C266 VN.n48 B 0.019433f
C267 VN.n49 B 0.036219f
C268 VN.n50 B 0.019433f
C269 VN.t1 B 2.48159f
C270 VN.n51 B 0.018358f
C271 VN.n52 B 0.019433f
C272 VN.t6 B 2.48159f
C273 VN.n53 B 0.920924f
C274 VN.t4 B 2.66818f
C275 VN.n54 B 0.897724f
C276 VN.n55 B 0.207347f
C277 VN.n56 B 0.02549f
C278 VN.n57 B 0.036219f
C279 VN.n58 B 0.035667f
C280 VN.n59 B 0.019433f
C281 VN.n60 B 0.019433f
C282 VN.n61 B 0.019433f
C283 VN.n62 B 0.038932f
C284 VN.n63 B 0.036219f
C285 VN.n64 B 0.880783f
C286 VN.n65 B 0.019433f
C287 VN.n66 B 0.019433f
C288 VN.n67 B 0.019433f
C289 VN.n68 B 0.038932f
C290 VN.n69 B 0.018358f
C291 VN.n70 B 0.035667f
C292 VN.n71 B 0.019433f
C293 VN.n72 B 0.019433f
C294 VN.n73 B 0.019433f
C295 VN.n74 B 0.02549f
C296 VN.n75 B 0.862446f
C297 VN.n76 B 0.029066f
C298 VN.n77 B 0.036219f
C299 VN.n78 B 0.019433f
C300 VN.n79 B 0.019433f
C301 VN.n80 B 0.019433f
C302 VN.n81 B 0.025662f
C303 VN.n82 B 0.036219f
C304 VN.n83 B 0.032643f
C305 VN.n84 B 0.031365f
C306 VN.n85 B 1.35401f
C307 VTAIL.t7 B 0.309068f
C308 VTAIL.t4 B 0.309068f
C309 VTAIL.n0 B 2.73753f
C310 VTAIL.n1 B 0.541043f
C311 VTAIL.n2 B 0.034077f
C312 VTAIL.n3 B 0.024128f
C313 VTAIL.n4 B 0.012965f
C314 VTAIL.n5 B 0.030645f
C315 VTAIL.n6 B 0.013728f
C316 VTAIL.n7 B 0.024128f
C317 VTAIL.n8 B 0.013347f
C318 VTAIL.n9 B 0.030645f
C319 VTAIL.n10 B 0.013728f
C320 VTAIL.n11 B 0.024128f
C321 VTAIL.n12 B 0.012965f
C322 VTAIL.n13 B 0.030645f
C323 VTAIL.n14 B 0.013728f
C324 VTAIL.n15 B 0.024128f
C325 VTAIL.n16 B 0.012965f
C326 VTAIL.n17 B 0.030645f
C327 VTAIL.n18 B 0.013728f
C328 VTAIL.n19 B 0.024128f
C329 VTAIL.n20 B 0.012965f
C330 VTAIL.n21 B 0.030645f
C331 VTAIL.n22 B 0.013728f
C332 VTAIL.n23 B 0.024128f
C333 VTAIL.n24 B 0.012965f
C334 VTAIL.n25 B 0.030645f
C335 VTAIL.n26 B 0.013728f
C336 VTAIL.n27 B 0.024128f
C337 VTAIL.n28 B 0.012965f
C338 VTAIL.n29 B 0.022984f
C339 VTAIL.n30 B 0.018103f
C340 VTAIL.t11 B 0.05063f
C341 VTAIL.n31 B 0.164687f
C342 VTAIL.n32 B 1.70359f
C343 VTAIL.n33 B 0.012965f
C344 VTAIL.n34 B 0.013728f
C345 VTAIL.n35 B 0.030645f
C346 VTAIL.n36 B 0.030645f
C347 VTAIL.n37 B 0.013728f
C348 VTAIL.n38 B 0.012965f
C349 VTAIL.n39 B 0.024128f
C350 VTAIL.n40 B 0.024128f
C351 VTAIL.n41 B 0.012965f
C352 VTAIL.n42 B 0.013728f
C353 VTAIL.n43 B 0.030645f
C354 VTAIL.n44 B 0.030645f
C355 VTAIL.n45 B 0.013728f
C356 VTAIL.n46 B 0.012965f
C357 VTAIL.n47 B 0.024128f
C358 VTAIL.n48 B 0.024128f
C359 VTAIL.n49 B 0.012965f
C360 VTAIL.n50 B 0.013728f
C361 VTAIL.n51 B 0.030645f
C362 VTAIL.n52 B 0.030645f
C363 VTAIL.n53 B 0.013728f
C364 VTAIL.n54 B 0.012965f
C365 VTAIL.n55 B 0.024128f
C366 VTAIL.n56 B 0.024128f
C367 VTAIL.n57 B 0.012965f
C368 VTAIL.n58 B 0.013728f
C369 VTAIL.n59 B 0.030645f
C370 VTAIL.n60 B 0.030645f
C371 VTAIL.n61 B 0.013728f
C372 VTAIL.n62 B 0.012965f
C373 VTAIL.n63 B 0.024128f
C374 VTAIL.n64 B 0.024128f
C375 VTAIL.n65 B 0.012965f
C376 VTAIL.n66 B 0.013728f
C377 VTAIL.n67 B 0.030645f
C378 VTAIL.n68 B 0.030645f
C379 VTAIL.n69 B 0.013728f
C380 VTAIL.n70 B 0.012965f
C381 VTAIL.n71 B 0.024128f
C382 VTAIL.n72 B 0.024128f
C383 VTAIL.n73 B 0.012965f
C384 VTAIL.n74 B 0.012965f
C385 VTAIL.n75 B 0.013728f
C386 VTAIL.n76 B 0.030645f
C387 VTAIL.n77 B 0.030645f
C388 VTAIL.n78 B 0.030645f
C389 VTAIL.n79 B 0.013347f
C390 VTAIL.n80 B 0.012965f
C391 VTAIL.n81 B 0.024128f
C392 VTAIL.n82 B 0.024128f
C393 VTAIL.n83 B 0.012965f
C394 VTAIL.n84 B 0.013728f
C395 VTAIL.n85 B 0.030645f
C396 VTAIL.n86 B 0.066629f
C397 VTAIL.n87 B 0.013728f
C398 VTAIL.n88 B 0.012965f
C399 VTAIL.n89 B 0.060055f
C400 VTAIL.n90 B 0.037439f
C401 VTAIL.n91 B 0.381261f
C402 VTAIL.t10 B 0.309068f
C403 VTAIL.t18 B 0.309068f
C404 VTAIL.n92 B 2.73753f
C405 VTAIL.n93 B 0.660844f
C406 VTAIL.t9 B 0.309068f
C407 VTAIL.t17 B 0.309068f
C408 VTAIL.n94 B 2.73753f
C409 VTAIL.n95 B 2.28948f
C410 VTAIL.t8 B 0.309068f
C411 VTAIL.t0 B 0.309068f
C412 VTAIL.n96 B 2.73754f
C413 VTAIL.n97 B 2.28947f
C414 VTAIL.t1 B 0.309068f
C415 VTAIL.t19 B 0.309068f
C416 VTAIL.n98 B 2.73754f
C417 VTAIL.n99 B 0.660832f
C418 VTAIL.n100 B 0.034077f
C419 VTAIL.n101 B 0.024128f
C420 VTAIL.n102 B 0.012965f
C421 VTAIL.n103 B 0.030645f
C422 VTAIL.n104 B 0.013728f
C423 VTAIL.n105 B 0.024128f
C424 VTAIL.n106 B 0.013347f
C425 VTAIL.n107 B 0.030645f
C426 VTAIL.n108 B 0.012965f
C427 VTAIL.n109 B 0.013728f
C428 VTAIL.n110 B 0.024128f
C429 VTAIL.n111 B 0.012965f
C430 VTAIL.n112 B 0.030645f
C431 VTAIL.n113 B 0.013728f
C432 VTAIL.n114 B 0.024128f
C433 VTAIL.n115 B 0.012965f
C434 VTAIL.n116 B 0.030645f
C435 VTAIL.n117 B 0.013728f
C436 VTAIL.n118 B 0.024128f
C437 VTAIL.n119 B 0.012965f
C438 VTAIL.n120 B 0.030645f
C439 VTAIL.n121 B 0.013728f
C440 VTAIL.n122 B 0.024128f
C441 VTAIL.n123 B 0.012965f
C442 VTAIL.n124 B 0.030645f
C443 VTAIL.n125 B 0.013728f
C444 VTAIL.n126 B 0.024128f
C445 VTAIL.n127 B 0.012965f
C446 VTAIL.n128 B 0.022984f
C447 VTAIL.n129 B 0.018103f
C448 VTAIL.t6 B 0.05063f
C449 VTAIL.n130 B 0.164687f
C450 VTAIL.n131 B 1.70359f
C451 VTAIL.n132 B 0.012965f
C452 VTAIL.n133 B 0.013728f
C453 VTAIL.n134 B 0.030645f
C454 VTAIL.n135 B 0.030645f
C455 VTAIL.n136 B 0.013728f
C456 VTAIL.n137 B 0.012965f
C457 VTAIL.n138 B 0.024128f
C458 VTAIL.n139 B 0.024128f
C459 VTAIL.n140 B 0.012965f
C460 VTAIL.n141 B 0.013728f
C461 VTAIL.n142 B 0.030645f
C462 VTAIL.n143 B 0.030645f
C463 VTAIL.n144 B 0.013728f
C464 VTAIL.n145 B 0.012965f
C465 VTAIL.n146 B 0.024128f
C466 VTAIL.n147 B 0.024128f
C467 VTAIL.n148 B 0.012965f
C468 VTAIL.n149 B 0.013728f
C469 VTAIL.n150 B 0.030645f
C470 VTAIL.n151 B 0.030645f
C471 VTAIL.n152 B 0.013728f
C472 VTAIL.n153 B 0.012965f
C473 VTAIL.n154 B 0.024128f
C474 VTAIL.n155 B 0.024128f
C475 VTAIL.n156 B 0.012965f
C476 VTAIL.n157 B 0.013728f
C477 VTAIL.n158 B 0.030645f
C478 VTAIL.n159 B 0.030645f
C479 VTAIL.n160 B 0.013728f
C480 VTAIL.n161 B 0.012965f
C481 VTAIL.n162 B 0.024128f
C482 VTAIL.n163 B 0.024128f
C483 VTAIL.n164 B 0.012965f
C484 VTAIL.n165 B 0.013728f
C485 VTAIL.n166 B 0.030645f
C486 VTAIL.n167 B 0.030645f
C487 VTAIL.n168 B 0.013728f
C488 VTAIL.n169 B 0.012965f
C489 VTAIL.n170 B 0.024128f
C490 VTAIL.n171 B 0.024128f
C491 VTAIL.n172 B 0.012965f
C492 VTAIL.n173 B 0.013728f
C493 VTAIL.n174 B 0.030645f
C494 VTAIL.n175 B 0.030645f
C495 VTAIL.n176 B 0.030645f
C496 VTAIL.n177 B 0.013347f
C497 VTAIL.n178 B 0.012965f
C498 VTAIL.n179 B 0.024128f
C499 VTAIL.n180 B 0.024128f
C500 VTAIL.n181 B 0.012965f
C501 VTAIL.n182 B 0.013728f
C502 VTAIL.n183 B 0.030645f
C503 VTAIL.n184 B 0.066629f
C504 VTAIL.n185 B 0.013728f
C505 VTAIL.n186 B 0.012965f
C506 VTAIL.n187 B 0.060055f
C507 VTAIL.n188 B 0.037439f
C508 VTAIL.n189 B 0.381261f
C509 VTAIL.t16 B 0.309068f
C510 VTAIL.t15 B 0.309068f
C511 VTAIL.n190 B 2.73754f
C512 VTAIL.n191 B 0.590124f
C513 VTAIL.t14 B 0.309068f
C514 VTAIL.t12 B 0.309068f
C515 VTAIL.n192 B 2.73754f
C516 VTAIL.n193 B 0.660832f
C517 VTAIL.n194 B 0.034077f
C518 VTAIL.n195 B 0.024128f
C519 VTAIL.n196 B 0.012965f
C520 VTAIL.n197 B 0.030645f
C521 VTAIL.n198 B 0.013728f
C522 VTAIL.n199 B 0.024128f
C523 VTAIL.n200 B 0.013347f
C524 VTAIL.n201 B 0.030645f
C525 VTAIL.n202 B 0.012965f
C526 VTAIL.n203 B 0.013728f
C527 VTAIL.n204 B 0.024128f
C528 VTAIL.n205 B 0.012965f
C529 VTAIL.n206 B 0.030645f
C530 VTAIL.n207 B 0.013728f
C531 VTAIL.n208 B 0.024128f
C532 VTAIL.n209 B 0.012965f
C533 VTAIL.n210 B 0.030645f
C534 VTAIL.n211 B 0.013728f
C535 VTAIL.n212 B 0.024128f
C536 VTAIL.n213 B 0.012965f
C537 VTAIL.n214 B 0.030645f
C538 VTAIL.n215 B 0.013728f
C539 VTAIL.n216 B 0.024128f
C540 VTAIL.n217 B 0.012965f
C541 VTAIL.n218 B 0.030645f
C542 VTAIL.n219 B 0.013728f
C543 VTAIL.n220 B 0.024128f
C544 VTAIL.n221 B 0.012965f
C545 VTAIL.n222 B 0.022984f
C546 VTAIL.n223 B 0.018103f
C547 VTAIL.t13 B 0.05063f
C548 VTAIL.n224 B 0.164687f
C549 VTAIL.n225 B 1.70359f
C550 VTAIL.n226 B 0.012965f
C551 VTAIL.n227 B 0.013728f
C552 VTAIL.n228 B 0.030645f
C553 VTAIL.n229 B 0.030645f
C554 VTAIL.n230 B 0.013728f
C555 VTAIL.n231 B 0.012965f
C556 VTAIL.n232 B 0.024128f
C557 VTAIL.n233 B 0.024128f
C558 VTAIL.n234 B 0.012965f
C559 VTAIL.n235 B 0.013728f
C560 VTAIL.n236 B 0.030645f
C561 VTAIL.n237 B 0.030645f
C562 VTAIL.n238 B 0.013728f
C563 VTAIL.n239 B 0.012965f
C564 VTAIL.n240 B 0.024128f
C565 VTAIL.n241 B 0.024128f
C566 VTAIL.n242 B 0.012965f
C567 VTAIL.n243 B 0.013728f
C568 VTAIL.n244 B 0.030645f
C569 VTAIL.n245 B 0.030645f
C570 VTAIL.n246 B 0.013728f
C571 VTAIL.n247 B 0.012965f
C572 VTAIL.n248 B 0.024128f
C573 VTAIL.n249 B 0.024128f
C574 VTAIL.n250 B 0.012965f
C575 VTAIL.n251 B 0.013728f
C576 VTAIL.n252 B 0.030645f
C577 VTAIL.n253 B 0.030645f
C578 VTAIL.n254 B 0.013728f
C579 VTAIL.n255 B 0.012965f
C580 VTAIL.n256 B 0.024128f
C581 VTAIL.n257 B 0.024128f
C582 VTAIL.n258 B 0.012965f
C583 VTAIL.n259 B 0.013728f
C584 VTAIL.n260 B 0.030645f
C585 VTAIL.n261 B 0.030645f
C586 VTAIL.n262 B 0.013728f
C587 VTAIL.n263 B 0.012965f
C588 VTAIL.n264 B 0.024128f
C589 VTAIL.n265 B 0.024128f
C590 VTAIL.n266 B 0.012965f
C591 VTAIL.n267 B 0.013728f
C592 VTAIL.n268 B 0.030645f
C593 VTAIL.n269 B 0.030645f
C594 VTAIL.n270 B 0.030645f
C595 VTAIL.n271 B 0.013347f
C596 VTAIL.n272 B 0.012965f
C597 VTAIL.n273 B 0.024128f
C598 VTAIL.n274 B 0.024128f
C599 VTAIL.n275 B 0.012965f
C600 VTAIL.n276 B 0.013728f
C601 VTAIL.n277 B 0.030645f
C602 VTAIL.n278 B 0.066629f
C603 VTAIL.n279 B 0.013728f
C604 VTAIL.n280 B 0.012965f
C605 VTAIL.n281 B 0.060055f
C606 VTAIL.n282 B 0.037439f
C607 VTAIL.n283 B 1.86614f
C608 VTAIL.n284 B 0.034077f
C609 VTAIL.n285 B 0.024128f
C610 VTAIL.n286 B 0.012965f
C611 VTAIL.n287 B 0.030645f
C612 VTAIL.n288 B 0.013728f
C613 VTAIL.n289 B 0.024128f
C614 VTAIL.n290 B 0.013347f
C615 VTAIL.n291 B 0.030645f
C616 VTAIL.n292 B 0.013728f
C617 VTAIL.n293 B 0.024128f
C618 VTAIL.n294 B 0.012965f
C619 VTAIL.n295 B 0.030645f
C620 VTAIL.n296 B 0.013728f
C621 VTAIL.n297 B 0.024128f
C622 VTAIL.n298 B 0.012965f
C623 VTAIL.n299 B 0.030645f
C624 VTAIL.n300 B 0.013728f
C625 VTAIL.n301 B 0.024128f
C626 VTAIL.n302 B 0.012965f
C627 VTAIL.n303 B 0.030645f
C628 VTAIL.n304 B 0.013728f
C629 VTAIL.n305 B 0.024128f
C630 VTAIL.n306 B 0.012965f
C631 VTAIL.n307 B 0.030645f
C632 VTAIL.n308 B 0.013728f
C633 VTAIL.n309 B 0.024128f
C634 VTAIL.n310 B 0.012965f
C635 VTAIL.n311 B 0.022984f
C636 VTAIL.n312 B 0.018103f
C637 VTAIL.t3 B 0.05063f
C638 VTAIL.n313 B 0.164687f
C639 VTAIL.n314 B 1.70359f
C640 VTAIL.n315 B 0.012965f
C641 VTAIL.n316 B 0.013728f
C642 VTAIL.n317 B 0.030645f
C643 VTAIL.n318 B 0.030645f
C644 VTAIL.n319 B 0.013728f
C645 VTAIL.n320 B 0.012965f
C646 VTAIL.n321 B 0.024128f
C647 VTAIL.n322 B 0.024128f
C648 VTAIL.n323 B 0.012965f
C649 VTAIL.n324 B 0.013728f
C650 VTAIL.n325 B 0.030645f
C651 VTAIL.n326 B 0.030645f
C652 VTAIL.n327 B 0.013728f
C653 VTAIL.n328 B 0.012965f
C654 VTAIL.n329 B 0.024128f
C655 VTAIL.n330 B 0.024128f
C656 VTAIL.n331 B 0.012965f
C657 VTAIL.n332 B 0.013728f
C658 VTAIL.n333 B 0.030645f
C659 VTAIL.n334 B 0.030645f
C660 VTAIL.n335 B 0.013728f
C661 VTAIL.n336 B 0.012965f
C662 VTAIL.n337 B 0.024128f
C663 VTAIL.n338 B 0.024128f
C664 VTAIL.n339 B 0.012965f
C665 VTAIL.n340 B 0.013728f
C666 VTAIL.n341 B 0.030645f
C667 VTAIL.n342 B 0.030645f
C668 VTAIL.n343 B 0.013728f
C669 VTAIL.n344 B 0.012965f
C670 VTAIL.n345 B 0.024128f
C671 VTAIL.n346 B 0.024128f
C672 VTAIL.n347 B 0.012965f
C673 VTAIL.n348 B 0.013728f
C674 VTAIL.n349 B 0.030645f
C675 VTAIL.n350 B 0.030645f
C676 VTAIL.n351 B 0.013728f
C677 VTAIL.n352 B 0.012965f
C678 VTAIL.n353 B 0.024128f
C679 VTAIL.n354 B 0.024128f
C680 VTAIL.n355 B 0.012965f
C681 VTAIL.n356 B 0.012965f
C682 VTAIL.n357 B 0.013728f
C683 VTAIL.n358 B 0.030645f
C684 VTAIL.n359 B 0.030645f
C685 VTAIL.n360 B 0.030645f
C686 VTAIL.n361 B 0.013347f
C687 VTAIL.n362 B 0.012965f
C688 VTAIL.n363 B 0.024128f
C689 VTAIL.n364 B 0.024128f
C690 VTAIL.n365 B 0.012965f
C691 VTAIL.n366 B 0.013728f
C692 VTAIL.n367 B 0.030645f
C693 VTAIL.n368 B 0.066629f
C694 VTAIL.n369 B 0.013728f
C695 VTAIL.n370 B 0.012965f
C696 VTAIL.n371 B 0.060055f
C697 VTAIL.n372 B 0.037439f
C698 VTAIL.n373 B 1.86614f
C699 VTAIL.t5 B 0.309068f
C700 VTAIL.t2 B 0.309068f
C701 VTAIL.n374 B 2.73753f
C702 VTAIL.n375 B 0.495468f
C703 VDD1.n0 B 0.033968f
C704 VDD1.n1 B 0.024051f
C705 VDD1.n2 B 0.012924f
C706 VDD1.n3 B 0.030547f
C707 VDD1.n4 B 0.013684f
C708 VDD1.n5 B 0.024051f
C709 VDD1.n6 B 0.013304f
C710 VDD1.n7 B 0.030547f
C711 VDD1.n8 B 0.012924f
C712 VDD1.n9 B 0.013684f
C713 VDD1.n10 B 0.024051f
C714 VDD1.n11 B 0.012924f
C715 VDD1.n12 B 0.030547f
C716 VDD1.n13 B 0.013684f
C717 VDD1.n14 B 0.024051f
C718 VDD1.n15 B 0.012924f
C719 VDD1.n16 B 0.030547f
C720 VDD1.n17 B 0.013684f
C721 VDD1.n18 B 0.024051f
C722 VDD1.n19 B 0.012924f
C723 VDD1.n20 B 0.030547f
C724 VDD1.n21 B 0.013684f
C725 VDD1.n22 B 0.024051f
C726 VDD1.n23 B 0.012924f
C727 VDD1.n24 B 0.030547f
C728 VDD1.n25 B 0.013684f
C729 VDD1.n26 B 0.024051f
C730 VDD1.n27 B 0.012924f
C731 VDD1.n28 B 0.02291f
C732 VDD1.n29 B 0.018045f
C733 VDD1.t7 B 0.050469f
C734 VDD1.n30 B 0.16416f
C735 VDD1.n31 B 1.69815f
C736 VDD1.n32 B 0.012924f
C737 VDD1.n33 B 0.013684f
C738 VDD1.n34 B 0.030547f
C739 VDD1.n35 B 0.030547f
C740 VDD1.n36 B 0.013684f
C741 VDD1.n37 B 0.012924f
C742 VDD1.n38 B 0.024051f
C743 VDD1.n39 B 0.024051f
C744 VDD1.n40 B 0.012924f
C745 VDD1.n41 B 0.013684f
C746 VDD1.n42 B 0.030547f
C747 VDD1.n43 B 0.030547f
C748 VDD1.n44 B 0.013684f
C749 VDD1.n45 B 0.012924f
C750 VDD1.n46 B 0.024051f
C751 VDD1.n47 B 0.024051f
C752 VDD1.n48 B 0.012924f
C753 VDD1.n49 B 0.013684f
C754 VDD1.n50 B 0.030547f
C755 VDD1.n51 B 0.030547f
C756 VDD1.n52 B 0.013684f
C757 VDD1.n53 B 0.012924f
C758 VDD1.n54 B 0.024051f
C759 VDD1.n55 B 0.024051f
C760 VDD1.n56 B 0.012924f
C761 VDD1.n57 B 0.013684f
C762 VDD1.n58 B 0.030547f
C763 VDD1.n59 B 0.030547f
C764 VDD1.n60 B 0.013684f
C765 VDD1.n61 B 0.012924f
C766 VDD1.n62 B 0.024051f
C767 VDD1.n63 B 0.024051f
C768 VDD1.n64 B 0.012924f
C769 VDD1.n65 B 0.013684f
C770 VDD1.n66 B 0.030547f
C771 VDD1.n67 B 0.030547f
C772 VDD1.n68 B 0.013684f
C773 VDD1.n69 B 0.012924f
C774 VDD1.n70 B 0.024051f
C775 VDD1.n71 B 0.024051f
C776 VDD1.n72 B 0.012924f
C777 VDD1.n73 B 0.013684f
C778 VDD1.n74 B 0.030547f
C779 VDD1.n75 B 0.030547f
C780 VDD1.n76 B 0.030547f
C781 VDD1.n77 B 0.013304f
C782 VDD1.n78 B 0.012924f
C783 VDD1.n79 B 0.024051f
C784 VDD1.n80 B 0.024051f
C785 VDD1.n81 B 0.012924f
C786 VDD1.n82 B 0.013684f
C787 VDD1.n83 B 0.030547f
C788 VDD1.n84 B 0.066416f
C789 VDD1.n85 B 0.013684f
C790 VDD1.n86 B 0.012924f
C791 VDD1.n87 B 0.059863f
C792 VDD1.n88 B 0.067271f
C793 VDD1.t5 B 0.308081f
C794 VDD1.t4 B 0.308081f
C795 VDD1.n89 B 2.79711f
C796 VDD1.n90 B 0.716432f
C797 VDD1.n91 B 0.033968f
C798 VDD1.n92 B 0.024051f
C799 VDD1.n93 B 0.012924f
C800 VDD1.n94 B 0.030547f
C801 VDD1.n95 B 0.013684f
C802 VDD1.n96 B 0.024051f
C803 VDD1.n97 B 0.013304f
C804 VDD1.n98 B 0.030547f
C805 VDD1.n99 B 0.013684f
C806 VDD1.n100 B 0.024051f
C807 VDD1.n101 B 0.012924f
C808 VDD1.n102 B 0.030547f
C809 VDD1.n103 B 0.013684f
C810 VDD1.n104 B 0.024051f
C811 VDD1.n105 B 0.012924f
C812 VDD1.n106 B 0.030547f
C813 VDD1.n107 B 0.013684f
C814 VDD1.n108 B 0.024051f
C815 VDD1.n109 B 0.012924f
C816 VDD1.n110 B 0.030547f
C817 VDD1.n111 B 0.013684f
C818 VDD1.n112 B 0.024051f
C819 VDD1.n113 B 0.012924f
C820 VDD1.n114 B 0.030547f
C821 VDD1.n115 B 0.013684f
C822 VDD1.n116 B 0.024051f
C823 VDD1.n117 B 0.012924f
C824 VDD1.n118 B 0.02291f
C825 VDD1.n119 B 0.018045f
C826 VDD1.t9 B 0.050469f
C827 VDD1.n120 B 0.16416f
C828 VDD1.n121 B 1.69815f
C829 VDD1.n122 B 0.012924f
C830 VDD1.n123 B 0.013684f
C831 VDD1.n124 B 0.030547f
C832 VDD1.n125 B 0.030547f
C833 VDD1.n126 B 0.013684f
C834 VDD1.n127 B 0.012924f
C835 VDD1.n128 B 0.024051f
C836 VDD1.n129 B 0.024051f
C837 VDD1.n130 B 0.012924f
C838 VDD1.n131 B 0.013684f
C839 VDD1.n132 B 0.030547f
C840 VDD1.n133 B 0.030547f
C841 VDD1.n134 B 0.013684f
C842 VDD1.n135 B 0.012924f
C843 VDD1.n136 B 0.024051f
C844 VDD1.n137 B 0.024051f
C845 VDD1.n138 B 0.012924f
C846 VDD1.n139 B 0.013684f
C847 VDD1.n140 B 0.030547f
C848 VDD1.n141 B 0.030547f
C849 VDD1.n142 B 0.013684f
C850 VDD1.n143 B 0.012924f
C851 VDD1.n144 B 0.024051f
C852 VDD1.n145 B 0.024051f
C853 VDD1.n146 B 0.012924f
C854 VDD1.n147 B 0.013684f
C855 VDD1.n148 B 0.030547f
C856 VDD1.n149 B 0.030547f
C857 VDD1.n150 B 0.013684f
C858 VDD1.n151 B 0.012924f
C859 VDD1.n152 B 0.024051f
C860 VDD1.n153 B 0.024051f
C861 VDD1.n154 B 0.012924f
C862 VDD1.n155 B 0.013684f
C863 VDD1.n156 B 0.030547f
C864 VDD1.n157 B 0.030547f
C865 VDD1.n158 B 0.013684f
C866 VDD1.n159 B 0.012924f
C867 VDD1.n160 B 0.024051f
C868 VDD1.n161 B 0.024051f
C869 VDD1.n162 B 0.012924f
C870 VDD1.n163 B 0.012924f
C871 VDD1.n164 B 0.013684f
C872 VDD1.n165 B 0.030547f
C873 VDD1.n166 B 0.030547f
C874 VDD1.n167 B 0.030547f
C875 VDD1.n168 B 0.013304f
C876 VDD1.n169 B 0.012924f
C877 VDD1.n170 B 0.024051f
C878 VDD1.n171 B 0.024051f
C879 VDD1.n172 B 0.012924f
C880 VDD1.n173 B 0.013684f
C881 VDD1.n174 B 0.030547f
C882 VDD1.n175 B 0.066416f
C883 VDD1.n176 B 0.013684f
C884 VDD1.n177 B 0.012924f
C885 VDD1.n178 B 0.059863f
C886 VDD1.n179 B 0.067271f
C887 VDD1.t8 B 0.308081f
C888 VDD1.t0 B 0.308081f
C889 VDD1.n180 B 2.7971f
C890 VDD1.n181 B 0.708521f
C891 VDD1.t6 B 0.308081f
C892 VDD1.t1 B 0.308081f
C893 VDD1.n182 B 2.81484f
C894 VDD1.n183 B 3.31165f
C895 VDD1.t2 B 0.308081f
C896 VDD1.t3 B 0.308081f
C897 VDD1.n184 B 2.7971f
C898 VDD1.n185 B 3.46451f
C899 VP.t7 B 2.515f
C900 VP.n0 B 0.948322f
C901 VP.n1 B 0.019695f
C902 VP.n2 B 0.031495f
C903 VP.n3 B 0.019695f
C904 VP.t0 B 2.515f
C905 VP.n4 B 0.036706f
C906 VP.n5 B 0.019695f
C907 VP.n6 B 0.036706f
C908 VP.n7 B 0.019695f
C909 VP.t8 B 2.515f
C910 VP.n8 B 0.018605f
C911 VP.n9 B 0.019695f
C912 VP.t1 B 2.515f
C913 VP.n10 B 0.874056f
C914 VP.n11 B 0.019695f
C915 VP.n12 B 0.026007f
C916 VP.n13 B 0.031787f
C917 VP.t9 B 2.515f
C918 VP.t5 B 2.515f
C919 VP.n14 B 0.948322f
C920 VP.n15 B 0.019695f
C921 VP.n16 B 0.031495f
C922 VP.n17 B 0.019695f
C923 VP.t6 B 2.515f
C924 VP.n18 B 0.036706f
C925 VP.n19 B 0.019695f
C926 VP.n20 B 0.036706f
C927 VP.n21 B 0.019695f
C928 VP.t4 B 2.515f
C929 VP.n22 B 0.018605f
C930 VP.n23 B 0.019695f
C931 VP.t3 B 2.515f
C932 VP.n24 B 0.933321f
C933 VP.t2 B 2.70409f
C934 VP.n25 B 0.909809f
C935 VP.n26 B 0.210139f
C936 VP.n27 B 0.025833f
C937 VP.n28 B 0.036706f
C938 VP.n29 B 0.036147f
C939 VP.n30 B 0.019695f
C940 VP.n31 B 0.019695f
C941 VP.n32 B 0.019695f
C942 VP.n33 B 0.039456f
C943 VP.n34 B 0.036706f
C944 VP.n35 B 0.89264f
C945 VP.n36 B 0.019695f
C946 VP.n37 B 0.019695f
C947 VP.n38 B 0.019695f
C948 VP.n39 B 0.039456f
C949 VP.n40 B 0.018605f
C950 VP.n41 B 0.036147f
C951 VP.n42 B 0.019695f
C952 VP.n43 B 0.019695f
C953 VP.n44 B 0.019695f
C954 VP.n45 B 0.025833f
C955 VP.n46 B 0.874056f
C956 VP.n47 B 0.029458f
C957 VP.n48 B 0.036706f
C958 VP.n49 B 0.019695f
C959 VP.n50 B 0.019695f
C960 VP.n51 B 0.019695f
C961 VP.n52 B 0.026007f
C962 VP.n53 B 0.036706f
C963 VP.n54 B 0.033082f
C964 VP.n55 B 0.031787f
C965 VP.n56 B 1.36454f
C966 VP.n57 B 1.37678f
C967 VP.n58 B 0.948322f
C968 VP.n59 B 0.033082f
C969 VP.n60 B 0.036706f
C970 VP.n61 B 0.019695f
C971 VP.n62 B 0.019695f
C972 VP.n63 B 0.019695f
C973 VP.n64 B 0.031495f
C974 VP.n65 B 0.036706f
C975 VP.n66 B 0.029458f
C976 VP.n67 B 0.019695f
C977 VP.n68 B 0.019695f
C978 VP.n69 B 0.025833f
C979 VP.n70 B 0.036706f
C980 VP.n71 B 0.036147f
C981 VP.n72 B 0.019695f
C982 VP.n73 B 0.019695f
C983 VP.n74 B 0.019695f
C984 VP.n75 B 0.039456f
C985 VP.n76 B 0.036706f
C986 VP.n77 B 0.89264f
C987 VP.n78 B 0.019695f
C988 VP.n79 B 0.019695f
C989 VP.n80 B 0.019695f
C990 VP.n81 B 0.039456f
C991 VP.n82 B 0.018605f
C992 VP.n83 B 0.036147f
C993 VP.n84 B 0.019695f
C994 VP.n85 B 0.019695f
C995 VP.n86 B 0.019695f
C996 VP.n87 B 0.025833f
C997 VP.n88 B 0.874056f
C998 VP.n89 B 0.029458f
C999 VP.n90 B 0.036706f
C1000 VP.n91 B 0.019695f
C1001 VP.n92 B 0.019695f
C1002 VP.n93 B 0.019695f
C1003 VP.n94 B 0.026007f
C1004 VP.n95 B 0.036706f
C1005 VP.n96 B 0.033082f
C1006 VP.n97 B 0.031787f
C1007 VP.n98 B 0.040506f
.ends

