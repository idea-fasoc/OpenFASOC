* NGSPICE file created from diff_pair_sample_0330.ext - technology: sky130A

.subckt diff_pair_sample_0330 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=4.5474 ps=24.1 w=11.66 l=3.56
X1 VDD2.t7 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=0 ps=0 w=11.66 l=3.56
X3 VTAIL.t8 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X4 VDD1.t5 VP.t2 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X5 VDD1.t4 VP.t3 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X6 VDD2.t6 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=4.5474 ps=24.1 w=11.66 l=3.56
X7 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X8 VTAIL.t15 VP.t4 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=1.9239 ps=11.99 w=11.66 l=3.56
X9 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X10 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=0 ps=0 w=11.66 l=3.56
X11 VTAIL.t10 VP.t5 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=1.9239 ps=11.99 w=11.66 l=3.56
X12 VTAIL.t2 VN.t4 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=1.9239 ps=11.99 w=11.66 l=3.56
X13 VTAIL.t5 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=1.9239 ps=11.99 w=11.66 l=3.56
X14 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=0 ps=0 w=11.66 l=3.56
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5474 pd=24.1 as=0 ps=0 w=11.66 l=3.56
X16 VDD2.t1 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=4.5474 ps=24.1 w=11.66 l=3.56
X17 VDD1.t1 VP.t6 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=4.5474 ps=24.1 w=11.66 l=3.56
X18 VTAIL.t13 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
X19 VDD2.t0 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9239 pd=11.99 as=1.9239 ps=11.99 w=11.66 l=3.56
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n23 VP.t5 111.246
R41 VP.n51 VP.n50 86.0649
R42 VP.n90 VP.n0 86.0649
R43 VP.n49 VP.n13 86.0649
R44 VP.n50 VP.t4 78.9348
R45 VP.n62 VP.t2 78.9348
R46 VP.n75 VP.t1 78.9348
R47 VP.n0 VP.t6 78.9348
R48 VP.n13 VP.t0 78.9348
R49 VP.n34 VP.t7 78.9348
R50 VP.n22 VP.t3 78.9348
R51 VP.n23 VP.n22 65.1845
R52 VP.n69 VP.n6 56.5617
R53 VP.n28 VP.n19 56.5617
R54 VP.n51 VP.n49 55.1435
R55 VP.n56 VP.n10 54.1398
R56 VP.n82 VP.n2 54.1398
R57 VP.n41 VP.n15 54.1398
R58 VP.n60 VP.n10 27.0143
R59 VP.n82 VP.n81 27.0143
R60 VP.n41 VP.n40 27.0143
R61 VP.n54 VP.n12 24.5923
R62 VP.n55 VP.n54 24.5923
R63 VP.n56 VP.n55 24.5923
R64 VP.n61 VP.n60 24.5923
R65 VP.n63 VP.n61 24.5923
R66 VP.n67 VP.n8 24.5923
R67 VP.n68 VP.n67 24.5923
R68 VP.n69 VP.n68 24.5923
R69 VP.n73 VP.n6 24.5923
R70 VP.n74 VP.n73 24.5923
R71 VP.n76 VP.n74 24.5923
R72 VP.n80 VP.n4 24.5923
R73 VP.n81 VP.n80 24.5923
R74 VP.n86 VP.n2 24.5923
R75 VP.n87 VP.n86 24.5923
R76 VP.n88 VP.n87 24.5923
R77 VP.n45 VP.n15 24.5923
R78 VP.n46 VP.n45 24.5923
R79 VP.n47 VP.n46 24.5923
R80 VP.n32 VP.n19 24.5923
R81 VP.n33 VP.n32 24.5923
R82 VP.n35 VP.n33 24.5923
R83 VP.n39 VP.n17 24.5923
R84 VP.n40 VP.n39 24.5923
R85 VP.n26 VP.n21 24.5923
R86 VP.n27 VP.n26 24.5923
R87 VP.n28 VP.n27 24.5923
R88 VP.n63 VP.n62 15.0015
R89 VP.n75 VP.n4 15.0015
R90 VP.n34 VP.n17 15.0015
R91 VP.n62 VP.n8 9.59132
R92 VP.n76 VP.n75 9.59132
R93 VP.n35 VP.n34 9.59132
R94 VP.n22 VP.n21 9.59132
R95 VP.n50 VP.n12 4.18111
R96 VP.n88 VP.n0 4.18111
R97 VP.n47 VP.n13 4.18111
R98 VP.n24 VP.n23 3.3307
R99 VP.n49 VP.n48 0.354861
R100 VP.n52 VP.n51 0.354861
R101 VP.n90 VP.n89 0.354861
R102 VP VP.n90 0.267071
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VTAIL.n11 VTAIL.t10 45.06
R142 VTAIL.n10 VTAIL.t1 45.06
R143 VTAIL.n7 VTAIL.t2 45.06
R144 VTAIL.n15 VTAIL.t3 45.0597
R145 VTAIL.n2 VTAIL.t5 45.0597
R146 VTAIL.n3 VTAIL.t12 45.0597
R147 VTAIL.n6 VTAIL.t15 45.0597
R148 VTAIL.n14 VTAIL.t14 45.0597
R149 VTAIL.n13 VTAIL.n12 43.3618
R150 VTAIL.n9 VTAIL.n8 43.3618
R151 VTAIL.n1 VTAIL.n0 43.3616
R152 VTAIL.n5 VTAIL.n4 43.3616
R153 VTAIL.n15 VTAIL.n14 25.7721
R154 VTAIL.n7 VTAIL.n6 25.7721
R155 VTAIL.n9 VTAIL.n7 3.35395
R156 VTAIL.n10 VTAIL.n9 3.35395
R157 VTAIL.n13 VTAIL.n11 3.35395
R158 VTAIL.n14 VTAIL.n13 3.35395
R159 VTAIL.n6 VTAIL.n5 3.35395
R160 VTAIL.n5 VTAIL.n3 3.35395
R161 VTAIL.n2 VTAIL.n1 3.35395
R162 VTAIL VTAIL.n15 3.29576
R163 VTAIL.n0 VTAIL.t7 1.69861
R164 VTAIL.n0 VTAIL.t0 1.69861
R165 VTAIL.n4 VTAIL.t11 1.69861
R166 VTAIL.n4 VTAIL.t8 1.69861
R167 VTAIL.n12 VTAIL.t9 1.69861
R168 VTAIL.n12 VTAIL.t13 1.69861
R169 VTAIL.n8 VTAIL.t4 1.69861
R170 VTAIL.n8 VTAIL.t6 1.69861
R171 VTAIL.n11 VTAIL.n10 0.470328
R172 VTAIL.n3 VTAIL.n2 0.470328
R173 VTAIL VTAIL.n1 0.0586897
R174 VDD1 VDD1.n0 61.7755
R175 VDD1.n3 VDD1.n2 61.6618
R176 VDD1.n3 VDD1.n1 61.6618
R177 VDD1.n5 VDD1.n4 60.0405
R178 VDD1.n5 VDD1.n3 49.4406
R179 VDD1.n4 VDD1.t0 1.69861
R180 VDD1.n4 VDD1.t7 1.69861
R181 VDD1.n0 VDD1.t2 1.69861
R182 VDD1.n0 VDD1.t4 1.69861
R183 VDD1.n2 VDD1.t6 1.69861
R184 VDD1.n2 VDD1.t1 1.69861
R185 VDD1.n1 VDD1.t3 1.69861
R186 VDD1.n1 VDD1.t5 1.69861
R187 VDD1 VDD1.n5 1.61903
R188 B.n992 B.n991 585
R189 B.n993 B.n992 585
R190 B.n350 B.n165 585
R191 B.n349 B.n348 585
R192 B.n347 B.n346 585
R193 B.n345 B.n344 585
R194 B.n343 B.n342 585
R195 B.n341 B.n340 585
R196 B.n339 B.n338 585
R197 B.n337 B.n336 585
R198 B.n335 B.n334 585
R199 B.n333 B.n332 585
R200 B.n331 B.n330 585
R201 B.n329 B.n328 585
R202 B.n327 B.n326 585
R203 B.n325 B.n324 585
R204 B.n323 B.n322 585
R205 B.n321 B.n320 585
R206 B.n319 B.n318 585
R207 B.n317 B.n316 585
R208 B.n315 B.n314 585
R209 B.n313 B.n312 585
R210 B.n311 B.n310 585
R211 B.n309 B.n308 585
R212 B.n307 B.n306 585
R213 B.n305 B.n304 585
R214 B.n303 B.n302 585
R215 B.n301 B.n300 585
R216 B.n299 B.n298 585
R217 B.n297 B.n296 585
R218 B.n295 B.n294 585
R219 B.n293 B.n292 585
R220 B.n291 B.n290 585
R221 B.n289 B.n288 585
R222 B.n287 B.n286 585
R223 B.n285 B.n284 585
R224 B.n283 B.n282 585
R225 B.n281 B.n280 585
R226 B.n279 B.n278 585
R227 B.n277 B.n276 585
R228 B.n275 B.n274 585
R229 B.n273 B.n272 585
R230 B.n271 B.n270 585
R231 B.n269 B.n268 585
R232 B.n267 B.n266 585
R233 B.n265 B.n264 585
R234 B.n263 B.n262 585
R235 B.n261 B.n260 585
R236 B.n259 B.n258 585
R237 B.n257 B.n256 585
R238 B.n255 B.n254 585
R239 B.n252 B.n251 585
R240 B.n250 B.n249 585
R241 B.n248 B.n247 585
R242 B.n246 B.n245 585
R243 B.n244 B.n243 585
R244 B.n242 B.n241 585
R245 B.n240 B.n239 585
R246 B.n238 B.n237 585
R247 B.n236 B.n235 585
R248 B.n234 B.n233 585
R249 B.n232 B.n231 585
R250 B.n230 B.n229 585
R251 B.n228 B.n227 585
R252 B.n226 B.n225 585
R253 B.n224 B.n223 585
R254 B.n222 B.n221 585
R255 B.n220 B.n219 585
R256 B.n218 B.n217 585
R257 B.n216 B.n215 585
R258 B.n214 B.n213 585
R259 B.n212 B.n211 585
R260 B.n210 B.n209 585
R261 B.n208 B.n207 585
R262 B.n206 B.n205 585
R263 B.n204 B.n203 585
R264 B.n202 B.n201 585
R265 B.n200 B.n199 585
R266 B.n198 B.n197 585
R267 B.n196 B.n195 585
R268 B.n194 B.n193 585
R269 B.n192 B.n191 585
R270 B.n190 B.n189 585
R271 B.n188 B.n187 585
R272 B.n186 B.n185 585
R273 B.n184 B.n183 585
R274 B.n182 B.n181 585
R275 B.n180 B.n179 585
R276 B.n178 B.n177 585
R277 B.n176 B.n175 585
R278 B.n174 B.n173 585
R279 B.n172 B.n171 585
R280 B.n990 B.n119 585
R281 B.n994 B.n119 585
R282 B.n989 B.n118 585
R283 B.n995 B.n118 585
R284 B.n988 B.n987 585
R285 B.n987 B.n114 585
R286 B.n986 B.n113 585
R287 B.n1001 B.n113 585
R288 B.n985 B.n112 585
R289 B.n1002 B.n112 585
R290 B.n984 B.n111 585
R291 B.n1003 B.n111 585
R292 B.n983 B.n982 585
R293 B.n982 B.n107 585
R294 B.n981 B.n106 585
R295 B.n1009 B.n106 585
R296 B.n980 B.n105 585
R297 B.n1010 B.n105 585
R298 B.n979 B.n104 585
R299 B.n1011 B.n104 585
R300 B.n978 B.n977 585
R301 B.n977 B.n100 585
R302 B.n976 B.n99 585
R303 B.n1017 B.n99 585
R304 B.n975 B.n98 585
R305 B.n1018 B.n98 585
R306 B.n974 B.n97 585
R307 B.n1019 B.n97 585
R308 B.n973 B.n972 585
R309 B.n972 B.n93 585
R310 B.n971 B.n92 585
R311 B.n1025 B.n92 585
R312 B.n970 B.n91 585
R313 B.n1026 B.n91 585
R314 B.n969 B.n90 585
R315 B.n1027 B.n90 585
R316 B.n968 B.n967 585
R317 B.n967 B.n86 585
R318 B.n966 B.n85 585
R319 B.n1033 B.n85 585
R320 B.n965 B.n84 585
R321 B.n1034 B.n84 585
R322 B.n964 B.n83 585
R323 B.n1035 B.n83 585
R324 B.n963 B.n962 585
R325 B.n962 B.n79 585
R326 B.n961 B.n78 585
R327 B.n1041 B.n78 585
R328 B.n960 B.n77 585
R329 B.n1042 B.n77 585
R330 B.n959 B.n76 585
R331 B.n1043 B.n76 585
R332 B.n958 B.n957 585
R333 B.n957 B.n72 585
R334 B.n956 B.n71 585
R335 B.n1049 B.n71 585
R336 B.n955 B.n70 585
R337 B.n1050 B.n70 585
R338 B.n954 B.n69 585
R339 B.n1051 B.n69 585
R340 B.n953 B.n952 585
R341 B.n952 B.n65 585
R342 B.n951 B.n64 585
R343 B.n1057 B.n64 585
R344 B.n950 B.n63 585
R345 B.n1058 B.n63 585
R346 B.n949 B.n62 585
R347 B.n1059 B.n62 585
R348 B.n948 B.n947 585
R349 B.n947 B.n58 585
R350 B.n946 B.n57 585
R351 B.n1065 B.n57 585
R352 B.n945 B.n56 585
R353 B.n1066 B.n56 585
R354 B.n944 B.n55 585
R355 B.n1067 B.n55 585
R356 B.n943 B.n942 585
R357 B.n942 B.n51 585
R358 B.n941 B.n50 585
R359 B.n1073 B.n50 585
R360 B.n940 B.n49 585
R361 B.n1074 B.n49 585
R362 B.n939 B.n48 585
R363 B.n1075 B.n48 585
R364 B.n938 B.n937 585
R365 B.n937 B.n44 585
R366 B.n936 B.n43 585
R367 B.n1081 B.n43 585
R368 B.n935 B.n42 585
R369 B.n1082 B.n42 585
R370 B.n934 B.n41 585
R371 B.n1083 B.n41 585
R372 B.n933 B.n932 585
R373 B.n932 B.n40 585
R374 B.n931 B.n36 585
R375 B.n1089 B.n36 585
R376 B.n930 B.n35 585
R377 B.n1090 B.n35 585
R378 B.n929 B.n34 585
R379 B.n1091 B.n34 585
R380 B.n928 B.n927 585
R381 B.n927 B.n30 585
R382 B.n926 B.n29 585
R383 B.n1097 B.n29 585
R384 B.n925 B.n28 585
R385 B.n1098 B.n28 585
R386 B.n924 B.n27 585
R387 B.n1099 B.n27 585
R388 B.n923 B.n922 585
R389 B.n922 B.n23 585
R390 B.n921 B.n22 585
R391 B.n1105 B.n22 585
R392 B.n920 B.n21 585
R393 B.n1106 B.n21 585
R394 B.n919 B.n20 585
R395 B.n1107 B.n20 585
R396 B.n918 B.n917 585
R397 B.n917 B.n19 585
R398 B.n916 B.n15 585
R399 B.n1113 B.n15 585
R400 B.n915 B.n14 585
R401 B.n1114 B.n14 585
R402 B.n914 B.n13 585
R403 B.n1115 B.n13 585
R404 B.n913 B.n912 585
R405 B.n912 B.n12 585
R406 B.n911 B.n910 585
R407 B.n911 B.n8 585
R408 B.n909 B.n7 585
R409 B.n1122 B.n7 585
R410 B.n908 B.n6 585
R411 B.n1123 B.n6 585
R412 B.n907 B.n5 585
R413 B.n1124 B.n5 585
R414 B.n906 B.n905 585
R415 B.n905 B.n4 585
R416 B.n904 B.n351 585
R417 B.n904 B.n903 585
R418 B.n894 B.n352 585
R419 B.n353 B.n352 585
R420 B.n896 B.n895 585
R421 B.n897 B.n896 585
R422 B.n893 B.n358 585
R423 B.n358 B.n357 585
R424 B.n892 B.n891 585
R425 B.n891 B.n890 585
R426 B.n360 B.n359 585
R427 B.n883 B.n360 585
R428 B.n882 B.n881 585
R429 B.n884 B.n882 585
R430 B.n880 B.n365 585
R431 B.n365 B.n364 585
R432 B.n879 B.n878 585
R433 B.n878 B.n877 585
R434 B.n367 B.n366 585
R435 B.n368 B.n367 585
R436 B.n870 B.n869 585
R437 B.n871 B.n870 585
R438 B.n868 B.n373 585
R439 B.n373 B.n372 585
R440 B.n867 B.n866 585
R441 B.n866 B.n865 585
R442 B.n375 B.n374 585
R443 B.n376 B.n375 585
R444 B.n858 B.n857 585
R445 B.n859 B.n858 585
R446 B.n856 B.n381 585
R447 B.n381 B.n380 585
R448 B.n855 B.n854 585
R449 B.n854 B.n853 585
R450 B.n383 B.n382 585
R451 B.n846 B.n383 585
R452 B.n845 B.n844 585
R453 B.n847 B.n845 585
R454 B.n843 B.n388 585
R455 B.n388 B.n387 585
R456 B.n842 B.n841 585
R457 B.n841 B.n840 585
R458 B.n390 B.n389 585
R459 B.n391 B.n390 585
R460 B.n833 B.n832 585
R461 B.n834 B.n833 585
R462 B.n831 B.n396 585
R463 B.n396 B.n395 585
R464 B.n830 B.n829 585
R465 B.n829 B.n828 585
R466 B.n398 B.n397 585
R467 B.n399 B.n398 585
R468 B.n821 B.n820 585
R469 B.n822 B.n821 585
R470 B.n819 B.n404 585
R471 B.n404 B.n403 585
R472 B.n818 B.n817 585
R473 B.n817 B.n816 585
R474 B.n406 B.n405 585
R475 B.n407 B.n406 585
R476 B.n809 B.n808 585
R477 B.n810 B.n809 585
R478 B.n807 B.n412 585
R479 B.n412 B.n411 585
R480 B.n806 B.n805 585
R481 B.n805 B.n804 585
R482 B.n414 B.n413 585
R483 B.n415 B.n414 585
R484 B.n797 B.n796 585
R485 B.n798 B.n797 585
R486 B.n795 B.n420 585
R487 B.n420 B.n419 585
R488 B.n794 B.n793 585
R489 B.n793 B.n792 585
R490 B.n422 B.n421 585
R491 B.n423 B.n422 585
R492 B.n785 B.n784 585
R493 B.n786 B.n785 585
R494 B.n783 B.n428 585
R495 B.n428 B.n427 585
R496 B.n782 B.n781 585
R497 B.n781 B.n780 585
R498 B.n430 B.n429 585
R499 B.n431 B.n430 585
R500 B.n773 B.n772 585
R501 B.n774 B.n773 585
R502 B.n771 B.n436 585
R503 B.n436 B.n435 585
R504 B.n770 B.n769 585
R505 B.n769 B.n768 585
R506 B.n438 B.n437 585
R507 B.n439 B.n438 585
R508 B.n761 B.n760 585
R509 B.n762 B.n761 585
R510 B.n759 B.n444 585
R511 B.n444 B.n443 585
R512 B.n758 B.n757 585
R513 B.n757 B.n756 585
R514 B.n446 B.n445 585
R515 B.n447 B.n446 585
R516 B.n749 B.n748 585
R517 B.n750 B.n749 585
R518 B.n747 B.n452 585
R519 B.n452 B.n451 585
R520 B.n746 B.n745 585
R521 B.n745 B.n744 585
R522 B.n454 B.n453 585
R523 B.n455 B.n454 585
R524 B.n737 B.n736 585
R525 B.n738 B.n737 585
R526 B.n735 B.n460 585
R527 B.n460 B.n459 585
R528 B.n734 B.n733 585
R529 B.n733 B.n732 585
R530 B.n462 B.n461 585
R531 B.n463 B.n462 585
R532 B.n725 B.n724 585
R533 B.n726 B.n725 585
R534 B.n723 B.n468 585
R535 B.n468 B.n467 585
R536 B.n722 B.n721 585
R537 B.n721 B.n720 585
R538 B.n470 B.n469 585
R539 B.n471 B.n470 585
R540 B.n713 B.n712 585
R541 B.n714 B.n713 585
R542 B.n711 B.n476 585
R543 B.n476 B.n475 585
R544 B.n705 B.n704 585
R545 B.n703 B.n523 585
R546 B.n702 B.n522 585
R547 B.n707 B.n522 585
R548 B.n701 B.n700 585
R549 B.n699 B.n698 585
R550 B.n697 B.n696 585
R551 B.n695 B.n694 585
R552 B.n693 B.n692 585
R553 B.n691 B.n690 585
R554 B.n689 B.n688 585
R555 B.n687 B.n686 585
R556 B.n685 B.n684 585
R557 B.n683 B.n682 585
R558 B.n681 B.n680 585
R559 B.n679 B.n678 585
R560 B.n677 B.n676 585
R561 B.n675 B.n674 585
R562 B.n673 B.n672 585
R563 B.n671 B.n670 585
R564 B.n669 B.n668 585
R565 B.n667 B.n666 585
R566 B.n665 B.n664 585
R567 B.n663 B.n662 585
R568 B.n661 B.n660 585
R569 B.n659 B.n658 585
R570 B.n657 B.n656 585
R571 B.n655 B.n654 585
R572 B.n653 B.n652 585
R573 B.n651 B.n650 585
R574 B.n649 B.n648 585
R575 B.n647 B.n646 585
R576 B.n645 B.n644 585
R577 B.n643 B.n642 585
R578 B.n641 B.n640 585
R579 B.n639 B.n638 585
R580 B.n637 B.n636 585
R581 B.n635 B.n634 585
R582 B.n633 B.n632 585
R583 B.n631 B.n630 585
R584 B.n629 B.n628 585
R585 B.n627 B.n626 585
R586 B.n625 B.n624 585
R587 B.n623 B.n622 585
R588 B.n621 B.n620 585
R589 B.n619 B.n618 585
R590 B.n617 B.n616 585
R591 B.n615 B.n614 585
R592 B.n613 B.n612 585
R593 B.n611 B.n610 585
R594 B.n609 B.n608 585
R595 B.n606 B.n605 585
R596 B.n604 B.n603 585
R597 B.n602 B.n601 585
R598 B.n600 B.n599 585
R599 B.n598 B.n597 585
R600 B.n596 B.n595 585
R601 B.n594 B.n593 585
R602 B.n592 B.n591 585
R603 B.n590 B.n589 585
R604 B.n588 B.n587 585
R605 B.n586 B.n585 585
R606 B.n584 B.n583 585
R607 B.n582 B.n581 585
R608 B.n580 B.n579 585
R609 B.n578 B.n577 585
R610 B.n576 B.n575 585
R611 B.n574 B.n573 585
R612 B.n572 B.n571 585
R613 B.n570 B.n569 585
R614 B.n568 B.n567 585
R615 B.n566 B.n565 585
R616 B.n564 B.n563 585
R617 B.n562 B.n561 585
R618 B.n560 B.n559 585
R619 B.n558 B.n557 585
R620 B.n556 B.n555 585
R621 B.n554 B.n553 585
R622 B.n552 B.n551 585
R623 B.n550 B.n549 585
R624 B.n548 B.n547 585
R625 B.n546 B.n545 585
R626 B.n544 B.n543 585
R627 B.n542 B.n541 585
R628 B.n540 B.n539 585
R629 B.n538 B.n537 585
R630 B.n536 B.n535 585
R631 B.n534 B.n533 585
R632 B.n532 B.n531 585
R633 B.n530 B.n529 585
R634 B.n478 B.n477 585
R635 B.n710 B.n709 585
R636 B.n474 B.n473 585
R637 B.n475 B.n474 585
R638 B.n716 B.n715 585
R639 B.n715 B.n714 585
R640 B.n717 B.n472 585
R641 B.n472 B.n471 585
R642 B.n719 B.n718 585
R643 B.n720 B.n719 585
R644 B.n466 B.n465 585
R645 B.n467 B.n466 585
R646 B.n728 B.n727 585
R647 B.n727 B.n726 585
R648 B.n729 B.n464 585
R649 B.n464 B.n463 585
R650 B.n731 B.n730 585
R651 B.n732 B.n731 585
R652 B.n458 B.n457 585
R653 B.n459 B.n458 585
R654 B.n740 B.n739 585
R655 B.n739 B.n738 585
R656 B.n741 B.n456 585
R657 B.n456 B.n455 585
R658 B.n743 B.n742 585
R659 B.n744 B.n743 585
R660 B.n450 B.n449 585
R661 B.n451 B.n450 585
R662 B.n752 B.n751 585
R663 B.n751 B.n750 585
R664 B.n753 B.n448 585
R665 B.n448 B.n447 585
R666 B.n755 B.n754 585
R667 B.n756 B.n755 585
R668 B.n442 B.n441 585
R669 B.n443 B.n442 585
R670 B.n764 B.n763 585
R671 B.n763 B.n762 585
R672 B.n765 B.n440 585
R673 B.n440 B.n439 585
R674 B.n767 B.n766 585
R675 B.n768 B.n767 585
R676 B.n434 B.n433 585
R677 B.n435 B.n434 585
R678 B.n776 B.n775 585
R679 B.n775 B.n774 585
R680 B.n777 B.n432 585
R681 B.n432 B.n431 585
R682 B.n779 B.n778 585
R683 B.n780 B.n779 585
R684 B.n426 B.n425 585
R685 B.n427 B.n426 585
R686 B.n788 B.n787 585
R687 B.n787 B.n786 585
R688 B.n789 B.n424 585
R689 B.n424 B.n423 585
R690 B.n791 B.n790 585
R691 B.n792 B.n791 585
R692 B.n418 B.n417 585
R693 B.n419 B.n418 585
R694 B.n800 B.n799 585
R695 B.n799 B.n798 585
R696 B.n801 B.n416 585
R697 B.n416 B.n415 585
R698 B.n803 B.n802 585
R699 B.n804 B.n803 585
R700 B.n410 B.n409 585
R701 B.n411 B.n410 585
R702 B.n812 B.n811 585
R703 B.n811 B.n810 585
R704 B.n813 B.n408 585
R705 B.n408 B.n407 585
R706 B.n815 B.n814 585
R707 B.n816 B.n815 585
R708 B.n402 B.n401 585
R709 B.n403 B.n402 585
R710 B.n824 B.n823 585
R711 B.n823 B.n822 585
R712 B.n825 B.n400 585
R713 B.n400 B.n399 585
R714 B.n827 B.n826 585
R715 B.n828 B.n827 585
R716 B.n394 B.n393 585
R717 B.n395 B.n394 585
R718 B.n836 B.n835 585
R719 B.n835 B.n834 585
R720 B.n837 B.n392 585
R721 B.n392 B.n391 585
R722 B.n839 B.n838 585
R723 B.n840 B.n839 585
R724 B.n386 B.n385 585
R725 B.n387 B.n386 585
R726 B.n849 B.n848 585
R727 B.n848 B.n847 585
R728 B.n850 B.n384 585
R729 B.n846 B.n384 585
R730 B.n852 B.n851 585
R731 B.n853 B.n852 585
R732 B.n379 B.n378 585
R733 B.n380 B.n379 585
R734 B.n861 B.n860 585
R735 B.n860 B.n859 585
R736 B.n862 B.n377 585
R737 B.n377 B.n376 585
R738 B.n864 B.n863 585
R739 B.n865 B.n864 585
R740 B.n371 B.n370 585
R741 B.n372 B.n371 585
R742 B.n873 B.n872 585
R743 B.n872 B.n871 585
R744 B.n874 B.n369 585
R745 B.n369 B.n368 585
R746 B.n876 B.n875 585
R747 B.n877 B.n876 585
R748 B.n363 B.n362 585
R749 B.n364 B.n363 585
R750 B.n886 B.n885 585
R751 B.n885 B.n884 585
R752 B.n887 B.n361 585
R753 B.n883 B.n361 585
R754 B.n889 B.n888 585
R755 B.n890 B.n889 585
R756 B.n356 B.n355 585
R757 B.n357 B.n356 585
R758 B.n899 B.n898 585
R759 B.n898 B.n897 585
R760 B.n900 B.n354 585
R761 B.n354 B.n353 585
R762 B.n902 B.n901 585
R763 B.n903 B.n902 585
R764 B.n3 B.n0 585
R765 B.n4 B.n3 585
R766 B.n1121 B.n1 585
R767 B.n1122 B.n1121 585
R768 B.n1120 B.n1119 585
R769 B.n1120 B.n8 585
R770 B.n1118 B.n9 585
R771 B.n12 B.n9 585
R772 B.n1117 B.n1116 585
R773 B.n1116 B.n1115 585
R774 B.n11 B.n10 585
R775 B.n1114 B.n11 585
R776 B.n1112 B.n1111 585
R777 B.n1113 B.n1112 585
R778 B.n1110 B.n16 585
R779 B.n19 B.n16 585
R780 B.n1109 B.n1108 585
R781 B.n1108 B.n1107 585
R782 B.n18 B.n17 585
R783 B.n1106 B.n18 585
R784 B.n1104 B.n1103 585
R785 B.n1105 B.n1104 585
R786 B.n1102 B.n24 585
R787 B.n24 B.n23 585
R788 B.n1101 B.n1100 585
R789 B.n1100 B.n1099 585
R790 B.n26 B.n25 585
R791 B.n1098 B.n26 585
R792 B.n1096 B.n1095 585
R793 B.n1097 B.n1096 585
R794 B.n1094 B.n31 585
R795 B.n31 B.n30 585
R796 B.n1093 B.n1092 585
R797 B.n1092 B.n1091 585
R798 B.n33 B.n32 585
R799 B.n1090 B.n33 585
R800 B.n1088 B.n1087 585
R801 B.n1089 B.n1088 585
R802 B.n1086 B.n37 585
R803 B.n40 B.n37 585
R804 B.n1085 B.n1084 585
R805 B.n1084 B.n1083 585
R806 B.n39 B.n38 585
R807 B.n1082 B.n39 585
R808 B.n1080 B.n1079 585
R809 B.n1081 B.n1080 585
R810 B.n1078 B.n45 585
R811 B.n45 B.n44 585
R812 B.n1077 B.n1076 585
R813 B.n1076 B.n1075 585
R814 B.n47 B.n46 585
R815 B.n1074 B.n47 585
R816 B.n1072 B.n1071 585
R817 B.n1073 B.n1072 585
R818 B.n1070 B.n52 585
R819 B.n52 B.n51 585
R820 B.n1069 B.n1068 585
R821 B.n1068 B.n1067 585
R822 B.n54 B.n53 585
R823 B.n1066 B.n54 585
R824 B.n1064 B.n1063 585
R825 B.n1065 B.n1064 585
R826 B.n1062 B.n59 585
R827 B.n59 B.n58 585
R828 B.n1061 B.n1060 585
R829 B.n1060 B.n1059 585
R830 B.n61 B.n60 585
R831 B.n1058 B.n61 585
R832 B.n1056 B.n1055 585
R833 B.n1057 B.n1056 585
R834 B.n1054 B.n66 585
R835 B.n66 B.n65 585
R836 B.n1053 B.n1052 585
R837 B.n1052 B.n1051 585
R838 B.n68 B.n67 585
R839 B.n1050 B.n68 585
R840 B.n1048 B.n1047 585
R841 B.n1049 B.n1048 585
R842 B.n1046 B.n73 585
R843 B.n73 B.n72 585
R844 B.n1045 B.n1044 585
R845 B.n1044 B.n1043 585
R846 B.n75 B.n74 585
R847 B.n1042 B.n75 585
R848 B.n1040 B.n1039 585
R849 B.n1041 B.n1040 585
R850 B.n1038 B.n80 585
R851 B.n80 B.n79 585
R852 B.n1037 B.n1036 585
R853 B.n1036 B.n1035 585
R854 B.n82 B.n81 585
R855 B.n1034 B.n82 585
R856 B.n1032 B.n1031 585
R857 B.n1033 B.n1032 585
R858 B.n1030 B.n87 585
R859 B.n87 B.n86 585
R860 B.n1029 B.n1028 585
R861 B.n1028 B.n1027 585
R862 B.n89 B.n88 585
R863 B.n1026 B.n89 585
R864 B.n1024 B.n1023 585
R865 B.n1025 B.n1024 585
R866 B.n1022 B.n94 585
R867 B.n94 B.n93 585
R868 B.n1021 B.n1020 585
R869 B.n1020 B.n1019 585
R870 B.n96 B.n95 585
R871 B.n1018 B.n96 585
R872 B.n1016 B.n1015 585
R873 B.n1017 B.n1016 585
R874 B.n1014 B.n101 585
R875 B.n101 B.n100 585
R876 B.n1013 B.n1012 585
R877 B.n1012 B.n1011 585
R878 B.n103 B.n102 585
R879 B.n1010 B.n103 585
R880 B.n1008 B.n1007 585
R881 B.n1009 B.n1008 585
R882 B.n1006 B.n108 585
R883 B.n108 B.n107 585
R884 B.n1005 B.n1004 585
R885 B.n1004 B.n1003 585
R886 B.n110 B.n109 585
R887 B.n1002 B.n110 585
R888 B.n1000 B.n999 585
R889 B.n1001 B.n1000 585
R890 B.n998 B.n115 585
R891 B.n115 B.n114 585
R892 B.n997 B.n996 585
R893 B.n996 B.n995 585
R894 B.n117 B.n116 585
R895 B.n994 B.n117 585
R896 B.n1125 B.n1124 585
R897 B.n1123 B.n2 585
R898 B.n171 B.n117 454.062
R899 B.n992 B.n119 454.062
R900 B.n709 B.n476 454.062
R901 B.n705 B.n474 454.062
R902 B.n169 B.t19 288.082
R903 B.n166 B.t15 288.082
R904 B.n527 B.t12 288.082
R905 B.n524 B.t8 288.082
R906 B.n993 B.n164 256.663
R907 B.n993 B.n163 256.663
R908 B.n993 B.n162 256.663
R909 B.n993 B.n161 256.663
R910 B.n993 B.n160 256.663
R911 B.n993 B.n159 256.663
R912 B.n993 B.n158 256.663
R913 B.n993 B.n157 256.663
R914 B.n993 B.n156 256.663
R915 B.n993 B.n155 256.663
R916 B.n993 B.n154 256.663
R917 B.n993 B.n153 256.663
R918 B.n993 B.n152 256.663
R919 B.n993 B.n151 256.663
R920 B.n993 B.n150 256.663
R921 B.n993 B.n149 256.663
R922 B.n993 B.n148 256.663
R923 B.n993 B.n147 256.663
R924 B.n993 B.n146 256.663
R925 B.n993 B.n145 256.663
R926 B.n993 B.n144 256.663
R927 B.n993 B.n143 256.663
R928 B.n993 B.n142 256.663
R929 B.n993 B.n141 256.663
R930 B.n993 B.n140 256.663
R931 B.n993 B.n139 256.663
R932 B.n993 B.n138 256.663
R933 B.n993 B.n137 256.663
R934 B.n993 B.n136 256.663
R935 B.n993 B.n135 256.663
R936 B.n993 B.n134 256.663
R937 B.n993 B.n133 256.663
R938 B.n993 B.n132 256.663
R939 B.n993 B.n131 256.663
R940 B.n993 B.n130 256.663
R941 B.n993 B.n129 256.663
R942 B.n993 B.n128 256.663
R943 B.n993 B.n127 256.663
R944 B.n993 B.n126 256.663
R945 B.n993 B.n125 256.663
R946 B.n993 B.n124 256.663
R947 B.n993 B.n123 256.663
R948 B.n993 B.n122 256.663
R949 B.n993 B.n121 256.663
R950 B.n993 B.n120 256.663
R951 B.n707 B.n706 256.663
R952 B.n707 B.n479 256.663
R953 B.n707 B.n480 256.663
R954 B.n707 B.n481 256.663
R955 B.n707 B.n482 256.663
R956 B.n707 B.n483 256.663
R957 B.n707 B.n484 256.663
R958 B.n707 B.n485 256.663
R959 B.n707 B.n486 256.663
R960 B.n707 B.n487 256.663
R961 B.n707 B.n488 256.663
R962 B.n707 B.n489 256.663
R963 B.n707 B.n490 256.663
R964 B.n707 B.n491 256.663
R965 B.n707 B.n492 256.663
R966 B.n707 B.n493 256.663
R967 B.n707 B.n494 256.663
R968 B.n707 B.n495 256.663
R969 B.n707 B.n496 256.663
R970 B.n707 B.n497 256.663
R971 B.n707 B.n498 256.663
R972 B.n707 B.n499 256.663
R973 B.n707 B.n500 256.663
R974 B.n707 B.n501 256.663
R975 B.n707 B.n502 256.663
R976 B.n707 B.n503 256.663
R977 B.n707 B.n504 256.663
R978 B.n707 B.n505 256.663
R979 B.n707 B.n506 256.663
R980 B.n707 B.n507 256.663
R981 B.n707 B.n508 256.663
R982 B.n707 B.n509 256.663
R983 B.n707 B.n510 256.663
R984 B.n707 B.n511 256.663
R985 B.n707 B.n512 256.663
R986 B.n707 B.n513 256.663
R987 B.n707 B.n514 256.663
R988 B.n707 B.n515 256.663
R989 B.n707 B.n516 256.663
R990 B.n707 B.n517 256.663
R991 B.n707 B.n518 256.663
R992 B.n707 B.n519 256.663
R993 B.n707 B.n520 256.663
R994 B.n707 B.n521 256.663
R995 B.n708 B.n707 256.663
R996 B.n1127 B.n1126 256.663
R997 B.n175 B.n174 163.367
R998 B.n179 B.n178 163.367
R999 B.n183 B.n182 163.367
R1000 B.n187 B.n186 163.367
R1001 B.n191 B.n190 163.367
R1002 B.n195 B.n194 163.367
R1003 B.n199 B.n198 163.367
R1004 B.n203 B.n202 163.367
R1005 B.n207 B.n206 163.367
R1006 B.n211 B.n210 163.367
R1007 B.n215 B.n214 163.367
R1008 B.n219 B.n218 163.367
R1009 B.n223 B.n222 163.367
R1010 B.n227 B.n226 163.367
R1011 B.n231 B.n230 163.367
R1012 B.n235 B.n234 163.367
R1013 B.n239 B.n238 163.367
R1014 B.n243 B.n242 163.367
R1015 B.n247 B.n246 163.367
R1016 B.n251 B.n250 163.367
R1017 B.n256 B.n255 163.367
R1018 B.n260 B.n259 163.367
R1019 B.n264 B.n263 163.367
R1020 B.n268 B.n267 163.367
R1021 B.n272 B.n271 163.367
R1022 B.n276 B.n275 163.367
R1023 B.n280 B.n279 163.367
R1024 B.n284 B.n283 163.367
R1025 B.n288 B.n287 163.367
R1026 B.n292 B.n291 163.367
R1027 B.n296 B.n295 163.367
R1028 B.n300 B.n299 163.367
R1029 B.n304 B.n303 163.367
R1030 B.n308 B.n307 163.367
R1031 B.n312 B.n311 163.367
R1032 B.n316 B.n315 163.367
R1033 B.n320 B.n319 163.367
R1034 B.n324 B.n323 163.367
R1035 B.n328 B.n327 163.367
R1036 B.n332 B.n331 163.367
R1037 B.n336 B.n335 163.367
R1038 B.n340 B.n339 163.367
R1039 B.n344 B.n343 163.367
R1040 B.n348 B.n347 163.367
R1041 B.n992 B.n165 163.367
R1042 B.n713 B.n476 163.367
R1043 B.n713 B.n470 163.367
R1044 B.n721 B.n470 163.367
R1045 B.n721 B.n468 163.367
R1046 B.n725 B.n468 163.367
R1047 B.n725 B.n462 163.367
R1048 B.n733 B.n462 163.367
R1049 B.n733 B.n460 163.367
R1050 B.n737 B.n460 163.367
R1051 B.n737 B.n454 163.367
R1052 B.n745 B.n454 163.367
R1053 B.n745 B.n452 163.367
R1054 B.n749 B.n452 163.367
R1055 B.n749 B.n446 163.367
R1056 B.n757 B.n446 163.367
R1057 B.n757 B.n444 163.367
R1058 B.n761 B.n444 163.367
R1059 B.n761 B.n438 163.367
R1060 B.n769 B.n438 163.367
R1061 B.n769 B.n436 163.367
R1062 B.n773 B.n436 163.367
R1063 B.n773 B.n430 163.367
R1064 B.n781 B.n430 163.367
R1065 B.n781 B.n428 163.367
R1066 B.n785 B.n428 163.367
R1067 B.n785 B.n422 163.367
R1068 B.n793 B.n422 163.367
R1069 B.n793 B.n420 163.367
R1070 B.n797 B.n420 163.367
R1071 B.n797 B.n414 163.367
R1072 B.n805 B.n414 163.367
R1073 B.n805 B.n412 163.367
R1074 B.n809 B.n412 163.367
R1075 B.n809 B.n406 163.367
R1076 B.n817 B.n406 163.367
R1077 B.n817 B.n404 163.367
R1078 B.n821 B.n404 163.367
R1079 B.n821 B.n398 163.367
R1080 B.n829 B.n398 163.367
R1081 B.n829 B.n396 163.367
R1082 B.n833 B.n396 163.367
R1083 B.n833 B.n390 163.367
R1084 B.n841 B.n390 163.367
R1085 B.n841 B.n388 163.367
R1086 B.n845 B.n388 163.367
R1087 B.n845 B.n383 163.367
R1088 B.n854 B.n383 163.367
R1089 B.n854 B.n381 163.367
R1090 B.n858 B.n381 163.367
R1091 B.n858 B.n375 163.367
R1092 B.n866 B.n375 163.367
R1093 B.n866 B.n373 163.367
R1094 B.n870 B.n373 163.367
R1095 B.n870 B.n367 163.367
R1096 B.n878 B.n367 163.367
R1097 B.n878 B.n365 163.367
R1098 B.n882 B.n365 163.367
R1099 B.n882 B.n360 163.367
R1100 B.n891 B.n360 163.367
R1101 B.n891 B.n358 163.367
R1102 B.n896 B.n358 163.367
R1103 B.n896 B.n352 163.367
R1104 B.n904 B.n352 163.367
R1105 B.n905 B.n904 163.367
R1106 B.n905 B.n5 163.367
R1107 B.n6 B.n5 163.367
R1108 B.n7 B.n6 163.367
R1109 B.n911 B.n7 163.367
R1110 B.n912 B.n911 163.367
R1111 B.n912 B.n13 163.367
R1112 B.n14 B.n13 163.367
R1113 B.n15 B.n14 163.367
R1114 B.n917 B.n15 163.367
R1115 B.n917 B.n20 163.367
R1116 B.n21 B.n20 163.367
R1117 B.n22 B.n21 163.367
R1118 B.n922 B.n22 163.367
R1119 B.n922 B.n27 163.367
R1120 B.n28 B.n27 163.367
R1121 B.n29 B.n28 163.367
R1122 B.n927 B.n29 163.367
R1123 B.n927 B.n34 163.367
R1124 B.n35 B.n34 163.367
R1125 B.n36 B.n35 163.367
R1126 B.n932 B.n36 163.367
R1127 B.n932 B.n41 163.367
R1128 B.n42 B.n41 163.367
R1129 B.n43 B.n42 163.367
R1130 B.n937 B.n43 163.367
R1131 B.n937 B.n48 163.367
R1132 B.n49 B.n48 163.367
R1133 B.n50 B.n49 163.367
R1134 B.n942 B.n50 163.367
R1135 B.n942 B.n55 163.367
R1136 B.n56 B.n55 163.367
R1137 B.n57 B.n56 163.367
R1138 B.n947 B.n57 163.367
R1139 B.n947 B.n62 163.367
R1140 B.n63 B.n62 163.367
R1141 B.n64 B.n63 163.367
R1142 B.n952 B.n64 163.367
R1143 B.n952 B.n69 163.367
R1144 B.n70 B.n69 163.367
R1145 B.n71 B.n70 163.367
R1146 B.n957 B.n71 163.367
R1147 B.n957 B.n76 163.367
R1148 B.n77 B.n76 163.367
R1149 B.n78 B.n77 163.367
R1150 B.n962 B.n78 163.367
R1151 B.n962 B.n83 163.367
R1152 B.n84 B.n83 163.367
R1153 B.n85 B.n84 163.367
R1154 B.n967 B.n85 163.367
R1155 B.n967 B.n90 163.367
R1156 B.n91 B.n90 163.367
R1157 B.n92 B.n91 163.367
R1158 B.n972 B.n92 163.367
R1159 B.n972 B.n97 163.367
R1160 B.n98 B.n97 163.367
R1161 B.n99 B.n98 163.367
R1162 B.n977 B.n99 163.367
R1163 B.n977 B.n104 163.367
R1164 B.n105 B.n104 163.367
R1165 B.n106 B.n105 163.367
R1166 B.n982 B.n106 163.367
R1167 B.n982 B.n111 163.367
R1168 B.n112 B.n111 163.367
R1169 B.n113 B.n112 163.367
R1170 B.n987 B.n113 163.367
R1171 B.n987 B.n118 163.367
R1172 B.n119 B.n118 163.367
R1173 B.n523 B.n522 163.367
R1174 B.n700 B.n522 163.367
R1175 B.n698 B.n697 163.367
R1176 B.n694 B.n693 163.367
R1177 B.n690 B.n689 163.367
R1178 B.n686 B.n685 163.367
R1179 B.n682 B.n681 163.367
R1180 B.n678 B.n677 163.367
R1181 B.n674 B.n673 163.367
R1182 B.n670 B.n669 163.367
R1183 B.n666 B.n665 163.367
R1184 B.n662 B.n661 163.367
R1185 B.n658 B.n657 163.367
R1186 B.n654 B.n653 163.367
R1187 B.n650 B.n649 163.367
R1188 B.n646 B.n645 163.367
R1189 B.n642 B.n641 163.367
R1190 B.n638 B.n637 163.367
R1191 B.n634 B.n633 163.367
R1192 B.n630 B.n629 163.367
R1193 B.n626 B.n625 163.367
R1194 B.n622 B.n621 163.367
R1195 B.n618 B.n617 163.367
R1196 B.n614 B.n613 163.367
R1197 B.n610 B.n609 163.367
R1198 B.n605 B.n604 163.367
R1199 B.n601 B.n600 163.367
R1200 B.n597 B.n596 163.367
R1201 B.n593 B.n592 163.367
R1202 B.n589 B.n588 163.367
R1203 B.n585 B.n584 163.367
R1204 B.n581 B.n580 163.367
R1205 B.n577 B.n576 163.367
R1206 B.n573 B.n572 163.367
R1207 B.n569 B.n568 163.367
R1208 B.n565 B.n564 163.367
R1209 B.n561 B.n560 163.367
R1210 B.n557 B.n556 163.367
R1211 B.n553 B.n552 163.367
R1212 B.n549 B.n548 163.367
R1213 B.n545 B.n544 163.367
R1214 B.n541 B.n540 163.367
R1215 B.n537 B.n536 163.367
R1216 B.n533 B.n532 163.367
R1217 B.n529 B.n478 163.367
R1218 B.n715 B.n474 163.367
R1219 B.n715 B.n472 163.367
R1220 B.n719 B.n472 163.367
R1221 B.n719 B.n466 163.367
R1222 B.n727 B.n466 163.367
R1223 B.n727 B.n464 163.367
R1224 B.n731 B.n464 163.367
R1225 B.n731 B.n458 163.367
R1226 B.n739 B.n458 163.367
R1227 B.n739 B.n456 163.367
R1228 B.n743 B.n456 163.367
R1229 B.n743 B.n450 163.367
R1230 B.n751 B.n450 163.367
R1231 B.n751 B.n448 163.367
R1232 B.n755 B.n448 163.367
R1233 B.n755 B.n442 163.367
R1234 B.n763 B.n442 163.367
R1235 B.n763 B.n440 163.367
R1236 B.n767 B.n440 163.367
R1237 B.n767 B.n434 163.367
R1238 B.n775 B.n434 163.367
R1239 B.n775 B.n432 163.367
R1240 B.n779 B.n432 163.367
R1241 B.n779 B.n426 163.367
R1242 B.n787 B.n426 163.367
R1243 B.n787 B.n424 163.367
R1244 B.n791 B.n424 163.367
R1245 B.n791 B.n418 163.367
R1246 B.n799 B.n418 163.367
R1247 B.n799 B.n416 163.367
R1248 B.n803 B.n416 163.367
R1249 B.n803 B.n410 163.367
R1250 B.n811 B.n410 163.367
R1251 B.n811 B.n408 163.367
R1252 B.n815 B.n408 163.367
R1253 B.n815 B.n402 163.367
R1254 B.n823 B.n402 163.367
R1255 B.n823 B.n400 163.367
R1256 B.n827 B.n400 163.367
R1257 B.n827 B.n394 163.367
R1258 B.n835 B.n394 163.367
R1259 B.n835 B.n392 163.367
R1260 B.n839 B.n392 163.367
R1261 B.n839 B.n386 163.367
R1262 B.n848 B.n386 163.367
R1263 B.n848 B.n384 163.367
R1264 B.n852 B.n384 163.367
R1265 B.n852 B.n379 163.367
R1266 B.n860 B.n379 163.367
R1267 B.n860 B.n377 163.367
R1268 B.n864 B.n377 163.367
R1269 B.n864 B.n371 163.367
R1270 B.n872 B.n371 163.367
R1271 B.n872 B.n369 163.367
R1272 B.n876 B.n369 163.367
R1273 B.n876 B.n363 163.367
R1274 B.n885 B.n363 163.367
R1275 B.n885 B.n361 163.367
R1276 B.n889 B.n361 163.367
R1277 B.n889 B.n356 163.367
R1278 B.n898 B.n356 163.367
R1279 B.n898 B.n354 163.367
R1280 B.n902 B.n354 163.367
R1281 B.n902 B.n3 163.367
R1282 B.n1125 B.n3 163.367
R1283 B.n1121 B.n2 163.367
R1284 B.n1121 B.n1120 163.367
R1285 B.n1120 B.n9 163.367
R1286 B.n1116 B.n9 163.367
R1287 B.n1116 B.n11 163.367
R1288 B.n1112 B.n11 163.367
R1289 B.n1112 B.n16 163.367
R1290 B.n1108 B.n16 163.367
R1291 B.n1108 B.n18 163.367
R1292 B.n1104 B.n18 163.367
R1293 B.n1104 B.n24 163.367
R1294 B.n1100 B.n24 163.367
R1295 B.n1100 B.n26 163.367
R1296 B.n1096 B.n26 163.367
R1297 B.n1096 B.n31 163.367
R1298 B.n1092 B.n31 163.367
R1299 B.n1092 B.n33 163.367
R1300 B.n1088 B.n33 163.367
R1301 B.n1088 B.n37 163.367
R1302 B.n1084 B.n37 163.367
R1303 B.n1084 B.n39 163.367
R1304 B.n1080 B.n39 163.367
R1305 B.n1080 B.n45 163.367
R1306 B.n1076 B.n45 163.367
R1307 B.n1076 B.n47 163.367
R1308 B.n1072 B.n47 163.367
R1309 B.n1072 B.n52 163.367
R1310 B.n1068 B.n52 163.367
R1311 B.n1068 B.n54 163.367
R1312 B.n1064 B.n54 163.367
R1313 B.n1064 B.n59 163.367
R1314 B.n1060 B.n59 163.367
R1315 B.n1060 B.n61 163.367
R1316 B.n1056 B.n61 163.367
R1317 B.n1056 B.n66 163.367
R1318 B.n1052 B.n66 163.367
R1319 B.n1052 B.n68 163.367
R1320 B.n1048 B.n68 163.367
R1321 B.n1048 B.n73 163.367
R1322 B.n1044 B.n73 163.367
R1323 B.n1044 B.n75 163.367
R1324 B.n1040 B.n75 163.367
R1325 B.n1040 B.n80 163.367
R1326 B.n1036 B.n80 163.367
R1327 B.n1036 B.n82 163.367
R1328 B.n1032 B.n82 163.367
R1329 B.n1032 B.n87 163.367
R1330 B.n1028 B.n87 163.367
R1331 B.n1028 B.n89 163.367
R1332 B.n1024 B.n89 163.367
R1333 B.n1024 B.n94 163.367
R1334 B.n1020 B.n94 163.367
R1335 B.n1020 B.n96 163.367
R1336 B.n1016 B.n96 163.367
R1337 B.n1016 B.n101 163.367
R1338 B.n1012 B.n101 163.367
R1339 B.n1012 B.n103 163.367
R1340 B.n1008 B.n103 163.367
R1341 B.n1008 B.n108 163.367
R1342 B.n1004 B.n108 163.367
R1343 B.n1004 B.n110 163.367
R1344 B.n1000 B.n110 163.367
R1345 B.n1000 B.n115 163.367
R1346 B.n996 B.n115 163.367
R1347 B.n996 B.n117 163.367
R1348 B.n166 B.t17 145.22
R1349 B.n527 B.t14 145.22
R1350 B.n169 B.t20 145.204
R1351 B.n524 B.t11 145.204
R1352 B.n170 B.n169 75.4429
R1353 B.n167 B.n166 75.4429
R1354 B.n528 B.n527 75.4429
R1355 B.n525 B.n524 75.4429
R1356 B.n707 B.n475 72.0997
R1357 B.n994 B.n993 72.0997
R1358 B.n171 B.n120 71.676
R1359 B.n175 B.n121 71.676
R1360 B.n179 B.n122 71.676
R1361 B.n183 B.n123 71.676
R1362 B.n187 B.n124 71.676
R1363 B.n191 B.n125 71.676
R1364 B.n195 B.n126 71.676
R1365 B.n199 B.n127 71.676
R1366 B.n203 B.n128 71.676
R1367 B.n207 B.n129 71.676
R1368 B.n211 B.n130 71.676
R1369 B.n215 B.n131 71.676
R1370 B.n219 B.n132 71.676
R1371 B.n223 B.n133 71.676
R1372 B.n227 B.n134 71.676
R1373 B.n231 B.n135 71.676
R1374 B.n235 B.n136 71.676
R1375 B.n239 B.n137 71.676
R1376 B.n243 B.n138 71.676
R1377 B.n247 B.n139 71.676
R1378 B.n251 B.n140 71.676
R1379 B.n256 B.n141 71.676
R1380 B.n260 B.n142 71.676
R1381 B.n264 B.n143 71.676
R1382 B.n268 B.n144 71.676
R1383 B.n272 B.n145 71.676
R1384 B.n276 B.n146 71.676
R1385 B.n280 B.n147 71.676
R1386 B.n284 B.n148 71.676
R1387 B.n288 B.n149 71.676
R1388 B.n292 B.n150 71.676
R1389 B.n296 B.n151 71.676
R1390 B.n300 B.n152 71.676
R1391 B.n304 B.n153 71.676
R1392 B.n308 B.n154 71.676
R1393 B.n312 B.n155 71.676
R1394 B.n316 B.n156 71.676
R1395 B.n320 B.n157 71.676
R1396 B.n324 B.n158 71.676
R1397 B.n328 B.n159 71.676
R1398 B.n332 B.n160 71.676
R1399 B.n336 B.n161 71.676
R1400 B.n340 B.n162 71.676
R1401 B.n344 B.n163 71.676
R1402 B.n348 B.n164 71.676
R1403 B.n165 B.n164 71.676
R1404 B.n347 B.n163 71.676
R1405 B.n343 B.n162 71.676
R1406 B.n339 B.n161 71.676
R1407 B.n335 B.n160 71.676
R1408 B.n331 B.n159 71.676
R1409 B.n327 B.n158 71.676
R1410 B.n323 B.n157 71.676
R1411 B.n319 B.n156 71.676
R1412 B.n315 B.n155 71.676
R1413 B.n311 B.n154 71.676
R1414 B.n307 B.n153 71.676
R1415 B.n303 B.n152 71.676
R1416 B.n299 B.n151 71.676
R1417 B.n295 B.n150 71.676
R1418 B.n291 B.n149 71.676
R1419 B.n287 B.n148 71.676
R1420 B.n283 B.n147 71.676
R1421 B.n279 B.n146 71.676
R1422 B.n275 B.n145 71.676
R1423 B.n271 B.n144 71.676
R1424 B.n267 B.n143 71.676
R1425 B.n263 B.n142 71.676
R1426 B.n259 B.n141 71.676
R1427 B.n255 B.n140 71.676
R1428 B.n250 B.n139 71.676
R1429 B.n246 B.n138 71.676
R1430 B.n242 B.n137 71.676
R1431 B.n238 B.n136 71.676
R1432 B.n234 B.n135 71.676
R1433 B.n230 B.n134 71.676
R1434 B.n226 B.n133 71.676
R1435 B.n222 B.n132 71.676
R1436 B.n218 B.n131 71.676
R1437 B.n214 B.n130 71.676
R1438 B.n210 B.n129 71.676
R1439 B.n206 B.n128 71.676
R1440 B.n202 B.n127 71.676
R1441 B.n198 B.n126 71.676
R1442 B.n194 B.n125 71.676
R1443 B.n190 B.n124 71.676
R1444 B.n186 B.n123 71.676
R1445 B.n182 B.n122 71.676
R1446 B.n178 B.n121 71.676
R1447 B.n174 B.n120 71.676
R1448 B.n706 B.n705 71.676
R1449 B.n700 B.n479 71.676
R1450 B.n697 B.n480 71.676
R1451 B.n693 B.n481 71.676
R1452 B.n689 B.n482 71.676
R1453 B.n685 B.n483 71.676
R1454 B.n681 B.n484 71.676
R1455 B.n677 B.n485 71.676
R1456 B.n673 B.n486 71.676
R1457 B.n669 B.n487 71.676
R1458 B.n665 B.n488 71.676
R1459 B.n661 B.n489 71.676
R1460 B.n657 B.n490 71.676
R1461 B.n653 B.n491 71.676
R1462 B.n649 B.n492 71.676
R1463 B.n645 B.n493 71.676
R1464 B.n641 B.n494 71.676
R1465 B.n637 B.n495 71.676
R1466 B.n633 B.n496 71.676
R1467 B.n629 B.n497 71.676
R1468 B.n625 B.n498 71.676
R1469 B.n621 B.n499 71.676
R1470 B.n617 B.n500 71.676
R1471 B.n613 B.n501 71.676
R1472 B.n609 B.n502 71.676
R1473 B.n604 B.n503 71.676
R1474 B.n600 B.n504 71.676
R1475 B.n596 B.n505 71.676
R1476 B.n592 B.n506 71.676
R1477 B.n588 B.n507 71.676
R1478 B.n584 B.n508 71.676
R1479 B.n580 B.n509 71.676
R1480 B.n576 B.n510 71.676
R1481 B.n572 B.n511 71.676
R1482 B.n568 B.n512 71.676
R1483 B.n564 B.n513 71.676
R1484 B.n560 B.n514 71.676
R1485 B.n556 B.n515 71.676
R1486 B.n552 B.n516 71.676
R1487 B.n548 B.n517 71.676
R1488 B.n544 B.n518 71.676
R1489 B.n540 B.n519 71.676
R1490 B.n536 B.n520 71.676
R1491 B.n532 B.n521 71.676
R1492 B.n708 B.n478 71.676
R1493 B.n706 B.n523 71.676
R1494 B.n698 B.n479 71.676
R1495 B.n694 B.n480 71.676
R1496 B.n690 B.n481 71.676
R1497 B.n686 B.n482 71.676
R1498 B.n682 B.n483 71.676
R1499 B.n678 B.n484 71.676
R1500 B.n674 B.n485 71.676
R1501 B.n670 B.n486 71.676
R1502 B.n666 B.n487 71.676
R1503 B.n662 B.n488 71.676
R1504 B.n658 B.n489 71.676
R1505 B.n654 B.n490 71.676
R1506 B.n650 B.n491 71.676
R1507 B.n646 B.n492 71.676
R1508 B.n642 B.n493 71.676
R1509 B.n638 B.n494 71.676
R1510 B.n634 B.n495 71.676
R1511 B.n630 B.n496 71.676
R1512 B.n626 B.n497 71.676
R1513 B.n622 B.n498 71.676
R1514 B.n618 B.n499 71.676
R1515 B.n614 B.n500 71.676
R1516 B.n610 B.n501 71.676
R1517 B.n605 B.n502 71.676
R1518 B.n601 B.n503 71.676
R1519 B.n597 B.n504 71.676
R1520 B.n593 B.n505 71.676
R1521 B.n589 B.n506 71.676
R1522 B.n585 B.n507 71.676
R1523 B.n581 B.n508 71.676
R1524 B.n577 B.n509 71.676
R1525 B.n573 B.n510 71.676
R1526 B.n569 B.n511 71.676
R1527 B.n565 B.n512 71.676
R1528 B.n561 B.n513 71.676
R1529 B.n557 B.n514 71.676
R1530 B.n553 B.n515 71.676
R1531 B.n549 B.n516 71.676
R1532 B.n545 B.n517 71.676
R1533 B.n541 B.n518 71.676
R1534 B.n537 B.n519 71.676
R1535 B.n533 B.n520 71.676
R1536 B.n529 B.n521 71.676
R1537 B.n709 B.n708 71.676
R1538 B.n1126 B.n1125 71.676
R1539 B.n1126 B.n2 71.676
R1540 B.n167 B.t18 69.7769
R1541 B.n528 B.t13 69.7769
R1542 B.n170 B.t21 69.7622
R1543 B.n525 B.t10 69.7622
R1544 B.n253 B.n170 59.5399
R1545 B.n168 B.n167 59.5399
R1546 B.n607 B.n528 59.5399
R1547 B.n526 B.n525 59.5399
R1548 B.n714 B.n475 44.1694
R1549 B.n714 B.n471 44.1694
R1550 B.n720 B.n471 44.1694
R1551 B.n720 B.n467 44.1694
R1552 B.n726 B.n467 44.1694
R1553 B.n726 B.n463 44.1694
R1554 B.n732 B.n463 44.1694
R1555 B.n732 B.n459 44.1694
R1556 B.n738 B.n459 44.1694
R1557 B.n744 B.n455 44.1694
R1558 B.n744 B.n451 44.1694
R1559 B.n750 B.n451 44.1694
R1560 B.n750 B.n447 44.1694
R1561 B.n756 B.n447 44.1694
R1562 B.n756 B.n443 44.1694
R1563 B.n762 B.n443 44.1694
R1564 B.n762 B.n439 44.1694
R1565 B.n768 B.n439 44.1694
R1566 B.n768 B.n435 44.1694
R1567 B.n774 B.n435 44.1694
R1568 B.n774 B.n431 44.1694
R1569 B.n780 B.n431 44.1694
R1570 B.n786 B.n427 44.1694
R1571 B.n786 B.n423 44.1694
R1572 B.n792 B.n423 44.1694
R1573 B.n792 B.n419 44.1694
R1574 B.n798 B.n419 44.1694
R1575 B.n798 B.n415 44.1694
R1576 B.n804 B.n415 44.1694
R1577 B.n804 B.n411 44.1694
R1578 B.n810 B.n411 44.1694
R1579 B.n810 B.n407 44.1694
R1580 B.n816 B.n407 44.1694
R1581 B.n822 B.n403 44.1694
R1582 B.n822 B.n399 44.1694
R1583 B.n828 B.n399 44.1694
R1584 B.n828 B.n395 44.1694
R1585 B.n834 B.n395 44.1694
R1586 B.n834 B.n391 44.1694
R1587 B.n840 B.n391 44.1694
R1588 B.n840 B.n387 44.1694
R1589 B.n847 B.n387 44.1694
R1590 B.n847 B.n846 44.1694
R1591 B.n853 B.n380 44.1694
R1592 B.n859 B.n380 44.1694
R1593 B.n859 B.n376 44.1694
R1594 B.n865 B.n376 44.1694
R1595 B.n865 B.n372 44.1694
R1596 B.n871 B.n372 44.1694
R1597 B.n871 B.n368 44.1694
R1598 B.n877 B.n368 44.1694
R1599 B.n877 B.n364 44.1694
R1600 B.n884 B.n364 44.1694
R1601 B.n884 B.n883 44.1694
R1602 B.n890 B.n357 44.1694
R1603 B.n897 B.n357 44.1694
R1604 B.n897 B.n353 44.1694
R1605 B.n903 B.n353 44.1694
R1606 B.n903 B.n4 44.1694
R1607 B.n1124 B.n4 44.1694
R1608 B.n1124 B.n1123 44.1694
R1609 B.n1123 B.n1122 44.1694
R1610 B.n1122 B.n8 44.1694
R1611 B.n12 B.n8 44.1694
R1612 B.n1115 B.n12 44.1694
R1613 B.n1115 B.n1114 44.1694
R1614 B.n1114 B.n1113 44.1694
R1615 B.n1107 B.n19 44.1694
R1616 B.n1107 B.n1106 44.1694
R1617 B.n1106 B.n1105 44.1694
R1618 B.n1105 B.n23 44.1694
R1619 B.n1099 B.n23 44.1694
R1620 B.n1099 B.n1098 44.1694
R1621 B.n1098 B.n1097 44.1694
R1622 B.n1097 B.n30 44.1694
R1623 B.n1091 B.n30 44.1694
R1624 B.n1091 B.n1090 44.1694
R1625 B.n1090 B.n1089 44.1694
R1626 B.n1083 B.n40 44.1694
R1627 B.n1083 B.n1082 44.1694
R1628 B.n1082 B.n1081 44.1694
R1629 B.n1081 B.n44 44.1694
R1630 B.n1075 B.n44 44.1694
R1631 B.n1075 B.n1074 44.1694
R1632 B.n1074 B.n1073 44.1694
R1633 B.n1073 B.n51 44.1694
R1634 B.n1067 B.n51 44.1694
R1635 B.n1067 B.n1066 44.1694
R1636 B.n1065 B.n58 44.1694
R1637 B.n1059 B.n58 44.1694
R1638 B.n1059 B.n1058 44.1694
R1639 B.n1058 B.n1057 44.1694
R1640 B.n1057 B.n65 44.1694
R1641 B.n1051 B.n65 44.1694
R1642 B.n1051 B.n1050 44.1694
R1643 B.n1050 B.n1049 44.1694
R1644 B.n1049 B.n72 44.1694
R1645 B.n1043 B.n72 44.1694
R1646 B.n1043 B.n1042 44.1694
R1647 B.n1041 B.n79 44.1694
R1648 B.n1035 B.n79 44.1694
R1649 B.n1035 B.n1034 44.1694
R1650 B.n1034 B.n1033 44.1694
R1651 B.n1033 B.n86 44.1694
R1652 B.n1027 B.n86 44.1694
R1653 B.n1027 B.n1026 44.1694
R1654 B.n1026 B.n1025 44.1694
R1655 B.n1025 B.n93 44.1694
R1656 B.n1019 B.n93 44.1694
R1657 B.n1019 B.n1018 44.1694
R1658 B.n1018 B.n1017 44.1694
R1659 B.n1017 B.n100 44.1694
R1660 B.n1011 B.n1010 44.1694
R1661 B.n1010 B.n1009 44.1694
R1662 B.n1009 B.n107 44.1694
R1663 B.n1003 B.n107 44.1694
R1664 B.n1003 B.n1002 44.1694
R1665 B.n1002 B.n1001 44.1694
R1666 B.n1001 B.n114 44.1694
R1667 B.n995 B.n114 44.1694
R1668 B.n995 B.n994 44.1694
R1669 B.n780 B.t2 37.674
R1670 B.t3 B.n1041 37.674
R1671 B.n890 B.t1 36.3749
R1672 B.n1113 B.t5 36.3749
R1673 B.t9 B.n455 35.0758
R1674 B.t16 B.n100 35.0758
R1675 B.n846 B.t6 32.4776
R1676 B.n40 B.t7 32.4776
R1677 B.t4 B.n403 31.1785
R1678 B.n1066 B.t0 31.1785
R1679 B.n704 B.n473 29.5029
R1680 B.n711 B.n710 29.5029
R1681 B.n172 B.n116 29.5029
R1682 B.n991 B.n990 29.5029
R1683 B B.n1127 18.0485
R1684 B.n816 B.t4 12.9913
R1685 B.t0 B.n1065 12.9913
R1686 B.n853 B.t6 11.6923
R1687 B.n1089 B.t7 11.6923
R1688 B.n716 B.n473 10.6151
R1689 B.n717 B.n716 10.6151
R1690 B.n718 B.n717 10.6151
R1691 B.n718 B.n465 10.6151
R1692 B.n728 B.n465 10.6151
R1693 B.n729 B.n728 10.6151
R1694 B.n730 B.n729 10.6151
R1695 B.n730 B.n457 10.6151
R1696 B.n740 B.n457 10.6151
R1697 B.n741 B.n740 10.6151
R1698 B.n742 B.n741 10.6151
R1699 B.n742 B.n449 10.6151
R1700 B.n752 B.n449 10.6151
R1701 B.n753 B.n752 10.6151
R1702 B.n754 B.n753 10.6151
R1703 B.n754 B.n441 10.6151
R1704 B.n764 B.n441 10.6151
R1705 B.n765 B.n764 10.6151
R1706 B.n766 B.n765 10.6151
R1707 B.n766 B.n433 10.6151
R1708 B.n776 B.n433 10.6151
R1709 B.n777 B.n776 10.6151
R1710 B.n778 B.n777 10.6151
R1711 B.n778 B.n425 10.6151
R1712 B.n788 B.n425 10.6151
R1713 B.n789 B.n788 10.6151
R1714 B.n790 B.n789 10.6151
R1715 B.n790 B.n417 10.6151
R1716 B.n800 B.n417 10.6151
R1717 B.n801 B.n800 10.6151
R1718 B.n802 B.n801 10.6151
R1719 B.n802 B.n409 10.6151
R1720 B.n812 B.n409 10.6151
R1721 B.n813 B.n812 10.6151
R1722 B.n814 B.n813 10.6151
R1723 B.n814 B.n401 10.6151
R1724 B.n824 B.n401 10.6151
R1725 B.n825 B.n824 10.6151
R1726 B.n826 B.n825 10.6151
R1727 B.n826 B.n393 10.6151
R1728 B.n836 B.n393 10.6151
R1729 B.n837 B.n836 10.6151
R1730 B.n838 B.n837 10.6151
R1731 B.n838 B.n385 10.6151
R1732 B.n849 B.n385 10.6151
R1733 B.n850 B.n849 10.6151
R1734 B.n851 B.n850 10.6151
R1735 B.n851 B.n378 10.6151
R1736 B.n861 B.n378 10.6151
R1737 B.n862 B.n861 10.6151
R1738 B.n863 B.n862 10.6151
R1739 B.n863 B.n370 10.6151
R1740 B.n873 B.n370 10.6151
R1741 B.n874 B.n873 10.6151
R1742 B.n875 B.n874 10.6151
R1743 B.n875 B.n362 10.6151
R1744 B.n886 B.n362 10.6151
R1745 B.n887 B.n886 10.6151
R1746 B.n888 B.n887 10.6151
R1747 B.n888 B.n355 10.6151
R1748 B.n899 B.n355 10.6151
R1749 B.n900 B.n899 10.6151
R1750 B.n901 B.n900 10.6151
R1751 B.n901 B.n0 10.6151
R1752 B.n704 B.n703 10.6151
R1753 B.n703 B.n702 10.6151
R1754 B.n702 B.n701 10.6151
R1755 B.n701 B.n699 10.6151
R1756 B.n699 B.n696 10.6151
R1757 B.n696 B.n695 10.6151
R1758 B.n695 B.n692 10.6151
R1759 B.n692 B.n691 10.6151
R1760 B.n691 B.n688 10.6151
R1761 B.n688 B.n687 10.6151
R1762 B.n687 B.n684 10.6151
R1763 B.n684 B.n683 10.6151
R1764 B.n683 B.n680 10.6151
R1765 B.n680 B.n679 10.6151
R1766 B.n679 B.n676 10.6151
R1767 B.n676 B.n675 10.6151
R1768 B.n675 B.n672 10.6151
R1769 B.n672 B.n671 10.6151
R1770 B.n671 B.n668 10.6151
R1771 B.n668 B.n667 10.6151
R1772 B.n667 B.n664 10.6151
R1773 B.n664 B.n663 10.6151
R1774 B.n663 B.n660 10.6151
R1775 B.n660 B.n659 10.6151
R1776 B.n659 B.n656 10.6151
R1777 B.n656 B.n655 10.6151
R1778 B.n655 B.n652 10.6151
R1779 B.n652 B.n651 10.6151
R1780 B.n651 B.n648 10.6151
R1781 B.n648 B.n647 10.6151
R1782 B.n647 B.n644 10.6151
R1783 B.n644 B.n643 10.6151
R1784 B.n643 B.n640 10.6151
R1785 B.n640 B.n639 10.6151
R1786 B.n639 B.n636 10.6151
R1787 B.n636 B.n635 10.6151
R1788 B.n635 B.n632 10.6151
R1789 B.n632 B.n631 10.6151
R1790 B.n631 B.n628 10.6151
R1791 B.n628 B.n627 10.6151
R1792 B.n624 B.n623 10.6151
R1793 B.n623 B.n620 10.6151
R1794 B.n620 B.n619 10.6151
R1795 B.n619 B.n616 10.6151
R1796 B.n616 B.n615 10.6151
R1797 B.n615 B.n612 10.6151
R1798 B.n612 B.n611 10.6151
R1799 B.n611 B.n608 10.6151
R1800 B.n606 B.n603 10.6151
R1801 B.n603 B.n602 10.6151
R1802 B.n602 B.n599 10.6151
R1803 B.n599 B.n598 10.6151
R1804 B.n598 B.n595 10.6151
R1805 B.n595 B.n594 10.6151
R1806 B.n594 B.n591 10.6151
R1807 B.n591 B.n590 10.6151
R1808 B.n590 B.n587 10.6151
R1809 B.n587 B.n586 10.6151
R1810 B.n586 B.n583 10.6151
R1811 B.n583 B.n582 10.6151
R1812 B.n582 B.n579 10.6151
R1813 B.n579 B.n578 10.6151
R1814 B.n578 B.n575 10.6151
R1815 B.n575 B.n574 10.6151
R1816 B.n574 B.n571 10.6151
R1817 B.n571 B.n570 10.6151
R1818 B.n570 B.n567 10.6151
R1819 B.n567 B.n566 10.6151
R1820 B.n566 B.n563 10.6151
R1821 B.n563 B.n562 10.6151
R1822 B.n562 B.n559 10.6151
R1823 B.n559 B.n558 10.6151
R1824 B.n558 B.n555 10.6151
R1825 B.n555 B.n554 10.6151
R1826 B.n554 B.n551 10.6151
R1827 B.n551 B.n550 10.6151
R1828 B.n550 B.n547 10.6151
R1829 B.n547 B.n546 10.6151
R1830 B.n546 B.n543 10.6151
R1831 B.n543 B.n542 10.6151
R1832 B.n542 B.n539 10.6151
R1833 B.n539 B.n538 10.6151
R1834 B.n538 B.n535 10.6151
R1835 B.n535 B.n534 10.6151
R1836 B.n534 B.n531 10.6151
R1837 B.n531 B.n530 10.6151
R1838 B.n530 B.n477 10.6151
R1839 B.n710 B.n477 10.6151
R1840 B.n712 B.n711 10.6151
R1841 B.n712 B.n469 10.6151
R1842 B.n722 B.n469 10.6151
R1843 B.n723 B.n722 10.6151
R1844 B.n724 B.n723 10.6151
R1845 B.n724 B.n461 10.6151
R1846 B.n734 B.n461 10.6151
R1847 B.n735 B.n734 10.6151
R1848 B.n736 B.n735 10.6151
R1849 B.n736 B.n453 10.6151
R1850 B.n746 B.n453 10.6151
R1851 B.n747 B.n746 10.6151
R1852 B.n748 B.n747 10.6151
R1853 B.n748 B.n445 10.6151
R1854 B.n758 B.n445 10.6151
R1855 B.n759 B.n758 10.6151
R1856 B.n760 B.n759 10.6151
R1857 B.n760 B.n437 10.6151
R1858 B.n770 B.n437 10.6151
R1859 B.n771 B.n770 10.6151
R1860 B.n772 B.n771 10.6151
R1861 B.n772 B.n429 10.6151
R1862 B.n782 B.n429 10.6151
R1863 B.n783 B.n782 10.6151
R1864 B.n784 B.n783 10.6151
R1865 B.n784 B.n421 10.6151
R1866 B.n794 B.n421 10.6151
R1867 B.n795 B.n794 10.6151
R1868 B.n796 B.n795 10.6151
R1869 B.n796 B.n413 10.6151
R1870 B.n806 B.n413 10.6151
R1871 B.n807 B.n806 10.6151
R1872 B.n808 B.n807 10.6151
R1873 B.n808 B.n405 10.6151
R1874 B.n818 B.n405 10.6151
R1875 B.n819 B.n818 10.6151
R1876 B.n820 B.n819 10.6151
R1877 B.n820 B.n397 10.6151
R1878 B.n830 B.n397 10.6151
R1879 B.n831 B.n830 10.6151
R1880 B.n832 B.n831 10.6151
R1881 B.n832 B.n389 10.6151
R1882 B.n842 B.n389 10.6151
R1883 B.n843 B.n842 10.6151
R1884 B.n844 B.n843 10.6151
R1885 B.n844 B.n382 10.6151
R1886 B.n855 B.n382 10.6151
R1887 B.n856 B.n855 10.6151
R1888 B.n857 B.n856 10.6151
R1889 B.n857 B.n374 10.6151
R1890 B.n867 B.n374 10.6151
R1891 B.n868 B.n867 10.6151
R1892 B.n869 B.n868 10.6151
R1893 B.n869 B.n366 10.6151
R1894 B.n879 B.n366 10.6151
R1895 B.n880 B.n879 10.6151
R1896 B.n881 B.n880 10.6151
R1897 B.n881 B.n359 10.6151
R1898 B.n892 B.n359 10.6151
R1899 B.n893 B.n892 10.6151
R1900 B.n895 B.n893 10.6151
R1901 B.n895 B.n894 10.6151
R1902 B.n894 B.n351 10.6151
R1903 B.n906 B.n351 10.6151
R1904 B.n907 B.n906 10.6151
R1905 B.n908 B.n907 10.6151
R1906 B.n909 B.n908 10.6151
R1907 B.n910 B.n909 10.6151
R1908 B.n913 B.n910 10.6151
R1909 B.n914 B.n913 10.6151
R1910 B.n915 B.n914 10.6151
R1911 B.n916 B.n915 10.6151
R1912 B.n918 B.n916 10.6151
R1913 B.n919 B.n918 10.6151
R1914 B.n920 B.n919 10.6151
R1915 B.n921 B.n920 10.6151
R1916 B.n923 B.n921 10.6151
R1917 B.n924 B.n923 10.6151
R1918 B.n925 B.n924 10.6151
R1919 B.n926 B.n925 10.6151
R1920 B.n928 B.n926 10.6151
R1921 B.n929 B.n928 10.6151
R1922 B.n930 B.n929 10.6151
R1923 B.n931 B.n930 10.6151
R1924 B.n933 B.n931 10.6151
R1925 B.n934 B.n933 10.6151
R1926 B.n935 B.n934 10.6151
R1927 B.n936 B.n935 10.6151
R1928 B.n938 B.n936 10.6151
R1929 B.n939 B.n938 10.6151
R1930 B.n940 B.n939 10.6151
R1931 B.n941 B.n940 10.6151
R1932 B.n943 B.n941 10.6151
R1933 B.n944 B.n943 10.6151
R1934 B.n945 B.n944 10.6151
R1935 B.n946 B.n945 10.6151
R1936 B.n948 B.n946 10.6151
R1937 B.n949 B.n948 10.6151
R1938 B.n950 B.n949 10.6151
R1939 B.n951 B.n950 10.6151
R1940 B.n953 B.n951 10.6151
R1941 B.n954 B.n953 10.6151
R1942 B.n955 B.n954 10.6151
R1943 B.n956 B.n955 10.6151
R1944 B.n958 B.n956 10.6151
R1945 B.n959 B.n958 10.6151
R1946 B.n960 B.n959 10.6151
R1947 B.n961 B.n960 10.6151
R1948 B.n963 B.n961 10.6151
R1949 B.n964 B.n963 10.6151
R1950 B.n965 B.n964 10.6151
R1951 B.n966 B.n965 10.6151
R1952 B.n968 B.n966 10.6151
R1953 B.n969 B.n968 10.6151
R1954 B.n970 B.n969 10.6151
R1955 B.n971 B.n970 10.6151
R1956 B.n973 B.n971 10.6151
R1957 B.n974 B.n973 10.6151
R1958 B.n975 B.n974 10.6151
R1959 B.n976 B.n975 10.6151
R1960 B.n978 B.n976 10.6151
R1961 B.n979 B.n978 10.6151
R1962 B.n980 B.n979 10.6151
R1963 B.n981 B.n980 10.6151
R1964 B.n983 B.n981 10.6151
R1965 B.n984 B.n983 10.6151
R1966 B.n985 B.n984 10.6151
R1967 B.n986 B.n985 10.6151
R1968 B.n988 B.n986 10.6151
R1969 B.n989 B.n988 10.6151
R1970 B.n990 B.n989 10.6151
R1971 B.n1119 B.n1 10.6151
R1972 B.n1119 B.n1118 10.6151
R1973 B.n1118 B.n1117 10.6151
R1974 B.n1117 B.n10 10.6151
R1975 B.n1111 B.n10 10.6151
R1976 B.n1111 B.n1110 10.6151
R1977 B.n1110 B.n1109 10.6151
R1978 B.n1109 B.n17 10.6151
R1979 B.n1103 B.n17 10.6151
R1980 B.n1103 B.n1102 10.6151
R1981 B.n1102 B.n1101 10.6151
R1982 B.n1101 B.n25 10.6151
R1983 B.n1095 B.n25 10.6151
R1984 B.n1095 B.n1094 10.6151
R1985 B.n1094 B.n1093 10.6151
R1986 B.n1093 B.n32 10.6151
R1987 B.n1087 B.n32 10.6151
R1988 B.n1087 B.n1086 10.6151
R1989 B.n1086 B.n1085 10.6151
R1990 B.n1085 B.n38 10.6151
R1991 B.n1079 B.n38 10.6151
R1992 B.n1079 B.n1078 10.6151
R1993 B.n1078 B.n1077 10.6151
R1994 B.n1077 B.n46 10.6151
R1995 B.n1071 B.n46 10.6151
R1996 B.n1071 B.n1070 10.6151
R1997 B.n1070 B.n1069 10.6151
R1998 B.n1069 B.n53 10.6151
R1999 B.n1063 B.n53 10.6151
R2000 B.n1063 B.n1062 10.6151
R2001 B.n1062 B.n1061 10.6151
R2002 B.n1061 B.n60 10.6151
R2003 B.n1055 B.n60 10.6151
R2004 B.n1055 B.n1054 10.6151
R2005 B.n1054 B.n1053 10.6151
R2006 B.n1053 B.n67 10.6151
R2007 B.n1047 B.n67 10.6151
R2008 B.n1047 B.n1046 10.6151
R2009 B.n1046 B.n1045 10.6151
R2010 B.n1045 B.n74 10.6151
R2011 B.n1039 B.n74 10.6151
R2012 B.n1039 B.n1038 10.6151
R2013 B.n1038 B.n1037 10.6151
R2014 B.n1037 B.n81 10.6151
R2015 B.n1031 B.n81 10.6151
R2016 B.n1031 B.n1030 10.6151
R2017 B.n1030 B.n1029 10.6151
R2018 B.n1029 B.n88 10.6151
R2019 B.n1023 B.n88 10.6151
R2020 B.n1023 B.n1022 10.6151
R2021 B.n1022 B.n1021 10.6151
R2022 B.n1021 B.n95 10.6151
R2023 B.n1015 B.n95 10.6151
R2024 B.n1015 B.n1014 10.6151
R2025 B.n1014 B.n1013 10.6151
R2026 B.n1013 B.n102 10.6151
R2027 B.n1007 B.n102 10.6151
R2028 B.n1007 B.n1006 10.6151
R2029 B.n1006 B.n1005 10.6151
R2030 B.n1005 B.n109 10.6151
R2031 B.n999 B.n109 10.6151
R2032 B.n999 B.n998 10.6151
R2033 B.n998 B.n997 10.6151
R2034 B.n997 B.n116 10.6151
R2035 B.n173 B.n172 10.6151
R2036 B.n176 B.n173 10.6151
R2037 B.n177 B.n176 10.6151
R2038 B.n180 B.n177 10.6151
R2039 B.n181 B.n180 10.6151
R2040 B.n184 B.n181 10.6151
R2041 B.n185 B.n184 10.6151
R2042 B.n188 B.n185 10.6151
R2043 B.n189 B.n188 10.6151
R2044 B.n192 B.n189 10.6151
R2045 B.n193 B.n192 10.6151
R2046 B.n196 B.n193 10.6151
R2047 B.n197 B.n196 10.6151
R2048 B.n200 B.n197 10.6151
R2049 B.n201 B.n200 10.6151
R2050 B.n204 B.n201 10.6151
R2051 B.n205 B.n204 10.6151
R2052 B.n208 B.n205 10.6151
R2053 B.n209 B.n208 10.6151
R2054 B.n212 B.n209 10.6151
R2055 B.n213 B.n212 10.6151
R2056 B.n216 B.n213 10.6151
R2057 B.n217 B.n216 10.6151
R2058 B.n220 B.n217 10.6151
R2059 B.n221 B.n220 10.6151
R2060 B.n224 B.n221 10.6151
R2061 B.n225 B.n224 10.6151
R2062 B.n228 B.n225 10.6151
R2063 B.n229 B.n228 10.6151
R2064 B.n232 B.n229 10.6151
R2065 B.n233 B.n232 10.6151
R2066 B.n236 B.n233 10.6151
R2067 B.n237 B.n236 10.6151
R2068 B.n240 B.n237 10.6151
R2069 B.n241 B.n240 10.6151
R2070 B.n244 B.n241 10.6151
R2071 B.n245 B.n244 10.6151
R2072 B.n248 B.n245 10.6151
R2073 B.n249 B.n248 10.6151
R2074 B.n252 B.n249 10.6151
R2075 B.n257 B.n254 10.6151
R2076 B.n258 B.n257 10.6151
R2077 B.n261 B.n258 10.6151
R2078 B.n262 B.n261 10.6151
R2079 B.n265 B.n262 10.6151
R2080 B.n266 B.n265 10.6151
R2081 B.n269 B.n266 10.6151
R2082 B.n270 B.n269 10.6151
R2083 B.n274 B.n273 10.6151
R2084 B.n277 B.n274 10.6151
R2085 B.n278 B.n277 10.6151
R2086 B.n281 B.n278 10.6151
R2087 B.n282 B.n281 10.6151
R2088 B.n285 B.n282 10.6151
R2089 B.n286 B.n285 10.6151
R2090 B.n289 B.n286 10.6151
R2091 B.n290 B.n289 10.6151
R2092 B.n293 B.n290 10.6151
R2093 B.n294 B.n293 10.6151
R2094 B.n297 B.n294 10.6151
R2095 B.n298 B.n297 10.6151
R2096 B.n301 B.n298 10.6151
R2097 B.n302 B.n301 10.6151
R2098 B.n305 B.n302 10.6151
R2099 B.n306 B.n305 10.6151
R2100 B.n309 B.n306 10.6151
R2101 B.n310 B.n309 10.6151
R2102 B.n313 B.n310 10.6151
R2103 B.n314 B.n313 10.6151
R2104 B.n317 B.n314 10.6151
R2105 B.n318 B.n317 10.6151
R2106 B.n321 B.n318 10.6151
R2107 B.n322 B.n321 10.6151
R2108 B.n325 B.n322 10.6151
R2109 B.n326 B.n325 10.6151
R2110 B.n329 B.n326 10.6151
R2111 B.n330 B.n329 10.6151
R2112 B.n333 B.n330 10.6151
R2113 B.n334 B.n333 10.6151
R2114 B.n337 B.n334 10.6151
R2115 B.n338 B.n337 10.6151
R2116 B.n341 B.n338 10.6151
R2117 B.n342 B.n341 10.6151
R2118 B.n345 B.n342 10.6151
R2119 B.n346 B.n345 10.6151
R2120 B.n349 B.n346 10.6151
R2121 B.n350 B.n349 10.6151
R2122 B.n991 B.n350 10.6151
R2123 B.n738 B.t9 9.09409
R2124 B.n1011 B.t16 9.09409
R2125 B.n1127 B.n0 8.11757
R2126 B.n1127 B.n1 8.11757
R2127 B.n883 B.t1 7.79501
R2128 B.n19 B.t5 7.79501
R2129 B.n624 B.n526 6.5566
R2130 B.n608 B.n607 6.5566
R2131 B.n254 B.n253 6.5566
R2132 B.n270 B.n168 6.5566
R2133 B.t2 B.n427 6.49592
R2134 B.n1042 B.t3 6.49592
R2135 B.n627 B.n526 4.05904
R2136 B.n607 B.n606 4.05904
R2137 B.n253 B.n252 4.05904
R2138 B.n273 B.n168 4.05904
R2139 VN.n72 VN.n71 161.3
R2140 VN.n70 VN.n38 161.3
R2141 VN.n69 VN.n68 161.3
R2142 VN.n67 VN.n39 161.3
R2143 VN.n66 VN.n65 161.3
R2144 VN.n64 VN.n40 161.3
R2145 VN.n63 VN.n62 161.3
R2146 VN.n61 VN.n41 161.3
R2147 VN.n60 VN.n59 161.3
R2148 VN.n58 VN.n42 161.3
R2149 VN.n57 VN.n56 161.3
R2150 VN.n55 VN.n44 161.3
R2151 VN.n54 VN.n53 161.3
R2152 VN.n52 VN.n45 161.3
R2153 VN.n51 VN.n50 161.3
R2154 VN.n49 VN.n46 161.3
R2155 VN.n35 VN.n34 161.3
R2156 VN.n33 VN.n1 161.3
R2157 VN.n32 VN.n31 161.3
R2158 VN.n30 VN.n2 161.3
R2159 VN.n29 VN.n28 161.3
R2160 VN.n27 VN.n3 161.3
R2161 VN.n26 VN.n25 161.3
R2162 VN.n24 VN.n4 161.3
R2163 VN.n23 VN.n22 161.3
R2164 VN.n20 VN.n5 161.3
R2165 VN.n19 VN.n18 161.3
R2166 VN.n17 VN.n6 161.3
R2167 VN.n16 VN.n15 161.3
R2168 VN.n14 VN.n7 161.3
R2169 VN.n13 VN.n12 161.3
R2170 VN.n11 VN.n8 161.3
R2171 VN.n48 VN.t6 111.246
R2172 VN.n10 VN.t5 111.246
R2173 VN.n36 VN.n0 86.0649
R2174 VN.n73 VN.n37 86.0649
R2175 VN.n9 VN.t7 78.9348
R2176 VN.n21 VN.t2 78.9348
R2177 VN.n0 VN.t1 78.9348
R2178 VN.n47 VN.t3 78.9348
R2179 VN.n43 VN.t0 78.9348
R2180 VN.n37 VN.t4 78.9348
R2181 VN.n10 VN.n9 65.1845
R2182 VN.n48 VN.n47 65.1845
R2183 VN.n15 VN.n6 56.5617
R2184 VN.n53 VN.n44 56.5617
R2185 VN VN.n73 55.3087
R2186 VN.n28 VN.n2 54.1398
R2187 VN.n65 VN.n39 54.1398
R2188 VN.n28 VN.n27 27.0143
R2189 VN.n65 VN.n64 27.0143
R2190 VN.n13 VN.n8 24.5923
R2191 VN.n14 VN.n13 24.5923
R2192 VN.n15 VN.n14 24.5923
R2193 VN.n19 VN.n6 24.5923
R2194 VN.n20 VN.n19 24.5923
R2195 VN.n22 VN.n20 24.5923
R2196 VN.n26 VN.n4 24.5923
R2197 VN.n27 VN.n26 24.5923
R2198 VN.n32 VN.n2 24.5923
R2199 VN.n33 VN.n32 24.5923
R2200 VN.n34 VN.n33 24.5923
R2201 VN.n53 VN.n52 24.5923
R2202 VN.n52 VN.n51 24.5923
R2203 VN.n51 VN.n46 24.5923
R2204 VN.n64 VN.n63 24.5923
R2205 VN.n63 VN.n41 24.5923
R2206 VN.n59 VN.n58 24.5923
R2207 VN.n58 VN.n57 24.5923
R2208 VN.n57 VN.n44 24.5923
R2209 VN.n71 VN.n70 24.5923
R2210 VN.n70 VN.n69 24.5923
R2211 VN.n69 VN.n39 24.5923
R2212 VN.n21 VN.n4 15.0015
R2213 VN.n43 VN.n41 15.0015
R2214 VN.n9 VN.n8 9.59132
R2215 VN.n22 VN.n21 9.59132
R2216 VN.n47 VN.n46 9.59132
R2217 VN.n59 VN.n43 9.59132
R2218 VN.n34 VN.n0 4.18111
R2219 VN.n71 VN.n37 4.18111
R2220 VN.n49 VN.n48 3.33072
R2221 VN.n11 VN.n10 3.33072
R2222 VN.n73 VN.n72 0.354861
R2223 VN.n36 VN.n35 0.354861
R2224 VN VN.n36 0.267071
R2225 VN.n72 VN.n38 0.189894
R2226 VN.n68 VN.n38 0.189894
R2227 VN.n68 VN.n67 0.189894
R2228 VN.n67 VN.n66 0.189894
R2229 VN.n66 VN.n40 0.189894
R2230 VN.n62 VN.n40 0.189894
R2231 VN.n62 VN.n61 0.189894
R2232 VN.n61 VN.n60 0.189894
R2233 VN.n60 VN.n42 0.189894
R2234 VN.n56 VN.n42 0.189894
R2235 VN.n56 VN.n55 0.189894
R2236 VN.n55 VN.n54 0.189894
R2237 VN.n54 VN.n45 0.189894
R2238 VN.n50 VN.n45 0.189894
R2239 VN.n50 VN.n49 0.189894
R2240 VN.n12 VN.n11 0.189894
R2241 VN.n12 VN.n7 0.189894
R2242 VN.n16 VN.n7 0.189894
R2243 VN.n17 VN.n16 0.189894
R2244 VN.n18 VN.n17 0.189894
R2245 VN.n18 VN.n5 0.189894
R2246 VN.n23 VN.n5 0.189894
R2247 VN.n24 VN.n23 0.189894
R2248 VN.n25 VN.n24 0.189894
R2249 VN.n25 VN.n3 0.189894
R2250 VN.n29 VN.n3 0.189894
R2251 VN.n30 VN.n29 0.189894
R2252 VN.n31 VN.n30 0.189894
R2253 VN.n31 VN.n1 0.189894
R2254 VN.n35 VN.n1 0.189894
R2255 VDD2.n2 VDD2.n1 61.6618
R2256 VDD2.n2 VDD2.n0 61.6618
R2257 VDD2 VDD2.n5 61.659
R2258 VDD2.n4 VDD2.n3 60.0406
R2259 VDD2.n4 VDD2.n2 48.8575
R2260 VDD2 VDD2.n4 1.73541
R2261 VDD2.n5 VDD2.t4 1.69861
R2262 VDD2.n5 VDD2.t1 1.69861
R2263 VDD2.n3 VDD2.t3 1.69861
R2264 VDD2.n3 VDD2.t7 1.69861
R2265 VDD2.n1 VDD2.t5 1.69861
R2266 VDD2.n1 VDD2.t6 1.69861
R2267 VDD2.n0 VDD2.t2 1.69861
R2268 VDD2.n0 VDD2.t0 1.69861
C0 VDD2 VP 0.622191f
C1 VN VP 8.77037f
C2 VDD2 VDD1 2.27529f
C3 VDD1 VN 0.15383f
C4 VTAIL VP 9.670549f
C5 VDD1 VTAIL 8.36542f
C6 VDD2 VN 8.923389f
C7 VDD1 VP 9.38987f
C8 VDD2 VTAIL 8.42627f
C9 VTAIL VN 9.656441f
C10 VDD2 B 6.346554f
C11 VDD1 B 6.89369f
C12 VTAIL B 10.93149f
C13 VN B 19.18117f
C14 VP B 17.836304f
C15 VDD2.t2 B 0.250435f
C16 VDD2.t0 B 0.250435f
C17 VDD2.n0 B 2.24282f
C18 VDD2.t5 B 0.250435f
C19 VDD2.t6 B 0.250435f
C20 VDD2.n1 B 2.24282f
C21 VDD2.n2 B 4.1488f
C22 VDD2.t3 B 0.250435f
C23 VDD2.t7 B 0.250435f
C24 VDD2.n3 B 2.2251f
C25 VDD2.n4 B 3.54484f
C26 VDD2.t4 B 0.250435f
C27 VDD2.t1 B 0.250435f
C28 VDD2.n5 B 2.24276f
C29 VN.t1 B 2.0548f
C30 VN.n0 B 0.786634f
C31 VN.n1 B 0.018183f
C32 VN.n2 B 0.031721f
C33 VN.n3 B 0.018183f
C34 VN.n4 B 0.027227f
C35 VN.n5 B 0.018183f
C36 VN.n6 B 0.026433f
C37 VN.n7 B 0.018183f
C38 VN.n8 B 0.023565f
C39 VN.t7 B 2.0548f
C40 VN.n9 B 0.782463f
C41 VN.t5 B 2.30361f
C42 VN.n10 B 0.746515f
C43 VN.n11 B 0.227319f
C44 VN.n12 B 0.018183f
C45 VN.n13 B 0.03372f
C46 VN.n14 B 0.03372f
C47 VN.n15 B 0.026433f
C48 VN.n16 B 0.018183f
C49 VN.n17 B 0.018183f
C50 VN.n18 B 0.018183f
C51 VN.n19 B 0.03372f
C52 VN.n20 B 0.03372f
C53 VN.t2 B 2.0548f
C54 VN.n21 B 0.721736f
C55 VN.n22 B 0.023565f
C56 VN.n23 B 0.018183f
C57 VN.n24 B 0.018183f
C58 VN.n25 B 0.018183f
C59 VN.n26 B 0.03372f
C60 VN.n27 B 0.035063f
C61 VN.n28 B 0.019801f
C62 VN.n29 B 0.018183f
C63 VN.n30 B 0.018183f
C64 VN.n31 B 0.018183f
C65 VN.n32 B 0.03372f
C66 VN.n33 B 0.03372f
C67 VN.n34 B 0.019903f
C68 VN.n35 B 0.029343f
C69 VN.n36 B 0.052715f
C70 VN.t4 B 2.0548f
C71 VN.n37 B 0.786634f
C72 VN.n38 B 0.018183f
C73 VN.n39 B 0.031721f
C74 VN.n40 B 0.018183f
C75 VN.n41 B 0.027227f
C76 VN.n42 B 0.018183f
C77 VN.t0 B 2.0548f
C78 VN.n43 B 0.721736f
C79 VN.n44 B 0.026433f
C80 VN.n45 B 0.018183f
C81 VN.n46 B 0.023565f
C82 VN.t6 B 2.30361f
C83 VN.t3 B 2.0548f
C84 VN.n47 B 0.782463f
C85 VN.n48 B 0.746515f
C86 VN.n49 B 0.227319f
C87 VN.n50 B 0.018183f
C88 VN.n51 B 0.03372f
C89 VN.n52 B 0.03372f
C90 VN.n53 B 0.026433f
C91 VN.n54 B 0.018183f
C92 VN.n55 B 0.018183f
C93 VN.n56 B 0.018183f
C94 VN.n57 B 0.03372f
C95 VN.n58 B 0.03372f
C96 VN.n59 B 0.023565f
C97 VN.n60 B 0.018183f
C98 VN.n61 B 0.018183f
C99 VN.n62 B 0.018183f
C100 VN.n63 B 0.03372f
C101 VN.n64 B 0.035063f
C102 VN.n65 B 0.019801f
C103 VN.n66 B 0.018183f
C104 VN.n67 B 0.018183f
C105 VN.n68 B 0.018183f
C106 VN.n69 B 0.03372f
C107 VN.n70 B 0.03372f
C108 VN.n71 B 0.019903f
C109 VN.n72 B 0.029343f
C110 VN.n73 B 1.20214f
C111 VDD1.t2 B 0.255515f
C112 VDD1.t4 B 0.255515f
C113 VDD1.n0 B 2.28982f
C114 VDD1.t3 B 0.255515f
C115 VDD1.t5 B 0.255515f
C116 VDD1.n1 B 2.28831f
C117 VDD1.t6 B 0.255515f
C118 VDD1.t1 B 0.255515f
C119 VDD1.n2 B 2.28831f
C120 VDD1.n3 B 4.29017f
C121 VDD1.t0 B 0.255515f
C122 VDD1.t7 B 0.255515f
C123 VDD1.n4 B 2.27022f
C124 VDD1.n5 B 3.65156f
C125 VTAIL.t7 B 0.190915f
C126 VTAIL.t0 B 0.190915f
C127 VTAIL.n0 B 1.63122f
C128 VTAIL.n1 B 0.437698f
C129 VTAIL.t5 B 2.078f
C130 VTAIL.n2 B 0.539083f
C131 VTAIL.t12 B 2.078f
C132 VTAIL.n3 B 0.539083f
C133 VTAIL.t11 B 0.190915f
C134 VTAIL.t8 B 0.190915f
C135 VTAIL.n4 B 1.63122f
C136 VTAIL.n5 B 0.657703f
C137 VTAIL.t15 B 2.078f
C138 VTAIL.n6 B 1.68416f
C139 VTAIL.t2 B 2.07801f
C140 VTAIL.n7 B 1.68415f
C141 VTAIL.t4 B 0.190915f
C142 VTAIL.t6 B 0.190915f
C143 VTAIL.n8 B 1.63123f
C144 VTAIL.n9 B 0.657698f
C145 VTAIL.t1 B 2.07801f
C146 VTAIL.n10 B 0.539077f
C147 VTAIL.t10 B 2.07801f
C148 VTAIL.n11 B 0.539077f
C149 VTAIL.t9 B 0.190915f
C150 VTAIL.t13 B 0.190915f
C151 VTAIL.n12 B 1.63123f
C152 VTAIL.n13 B 0.657698f
C153 VTAIL.t14 B 2.078f
C154 VTAIL.n14 B 1.68416f
C155 VTAIL.t3 B 2.078f
C156 VTAIL.n15 B 1.68027f
C157 VP.t6 B 2.09425f
C158 VP.n0 B 0.801737f
C159 VP.n1 B 0.018533f
C160 VP.n2 B 0.03233f
C161 VP.n3 B 0.018533f
C162 VP.n4 B 0.02775f
C163 VP.n5 B 0.018533f
C164 VP.n6 B 0.02694f
C165 VP.n7 B 0.018533f
C166 VP.n8 B 0.024018f
C167 VP.n9 B 0.018533f
C168 VP.n10 B 0.020181f
C169 VP.n11 B 0.018533f
C170 VP.n12 B 0.020285f
C171 VP.t0 B 2.09425f
C172 VP.n13 B 0.801737f
C173 VP.n14 B 0.018533f
C174 VP.n15 B 0.03233f
C175 VP.n16 B 0.018533f
C176 VP.n17 B 0.02775f
C177 VP.n18 B 0.018533f
C178 VP.n19 B 0.02694f
C179 VP.n20 B 0.018533f
C180 VP.n21 B 0.024018f
C181 VP.t5 B 2.34784f
C182 VP.t3 B 2.09425f
C183 VP.n22 B 0.797485f
C184 VP.n23 B 0.760848f
C185 VP.n24 B 0.231684f
C186 VP.n25 B 0.018533f
C187 VP.n26 B 0.034367f
C188 VP.n27 B 0.034367f
C189 VP.n28 B 0.02694f
C190 VP.n29 B 0.018533f
C191 VP.n30 B 0.018533f
C192 VP.n31 B 0.018533f
C193 VP.n32 B 0.034367f
C194 VP.n33 B 0.034367f
C195 VP.t7 B 2.09425f
C196 VP.n34 B 0.735593f
C197 VP.n35 B 0.024018f
C198 VP.n36 B 0.018533f
C199 VP.n37 B 0.018533f
C200 VP.n38 B 0.018533f
C201 VP.n39 B 0.034367f
C202 VP.n40 B 0.035736f
C203 VP.n41 B 0.020181f
C204 VP.n42 B 0.018533f
C205 VP.n43 B 0.018533f
C206 VP.n44 B 0.018533f
C207 VP.n45 B 0.034367f
C208 VP.n46 B 0.034367f
C209 VP.n47 B 0.020285f
C210 VP.n48 B 0.029906f
C211 VP.n49 B 1.21788f
C212 VP.t4 B 2.09425f
C213 VP.n50 B 0.801737f
C214 VP.n51 B 1.23f
C215 VP.n52 B 0.029906f
C216 VP.n53 B 0.018533f
C217 VP.n54 B 0.034367f
C218 VP.n55 B 0.034367f
C219 VP.n56 B 0.03233f
C220 VP.n57 B 0.018533f
C221 VP.n58 B 0.018533f
C222 VP.n59 B 0.018533f
C223 VP.n60 B 0.035736f
C224 VP.n61 B 0.034367f
C225 VP.t2 B 2.09425f
C226 VP.n62 B 0.735593f
C227 VP.n63 B 0.02775f
C228 VP.n64 B 0.018533f
C229 VP.n65 B 0.018533f
C230 VP.n66 B 0.018533f
C231 VP.n67 B 0.034367f
C232 VP.n68 B 0.034367f
C233 VP.n69 B 0.02694f
C234 VP.n70 B 0.018533f
C235 VP.n71 B 0.018533f
C236 VP.n72 B 0.018533f
C237 VP.n73 B 0.034367f
C238 VP.n74 B 0.034367f
C239 VP.t1 B 2.09425f
C240 VP.n75 B 0.735593f
C241 VP.n76 B 0.024018f
C242 VP.n77 B 0.018533f
C243 VP.n78 B 0.018533f
C244 VP.n79 B 0.018533f
C245 VP.n80 B 0.034367f
C246 VP.n81 B 0.035736f
C247 VP.n82 B 0.020181f
C248 VP.n83 B 0.018533f
C249 VP.n84 B 0.018533f
C250 VP.n85 B 0.018533f
C251 VP.n86 B 0.034367f
C252 VP.n87 B 0.034367f
C253 VP.n88 B 0.020285f
C254 VP.n89 B 0.029906f
C255 VP.n90 B 0.053727f
.ends

