* NGSPICE file created from diff_pair_sample_1700.ext - technology: sky130A

.subckt diff_pair_sample_1700 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=0 ps=0 w=14.39 l=1.24
X1 VDD1.t9 VP.t0 VTAIL.t13 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=5.6121 ps=29.56 w=14.39 l=1.24
X2 VDD1.t8 VP.t1 VTAIL.t18 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=2.37435 ps=14.72 w=14.39 l=1.24
X3 B.t8 B.t6 B.t7 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=0 ps=0 w=14.39 l=1.24
X4 VTAIL.t7 VN.t0 VDD2.t9 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X5 VTAIL.t2 VN.t1 VDD2.t8 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X6 B.t5 B.t3 B.t4 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=0 ps=0 w=14.39 l=1.24
X7 VDD1.t7 VP.t2 VTAIL.t14 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X8 VTAIL.t12 VP.t3 VDD1.t6 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X9 VDD2.t7 VN.t2 VTAIL.t6 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=5.6121 ps=29.56 w=14.39 l=1.24
X10 VDD1.t5 VP.t4 VTAIL.t15 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X11 VDD1.t4 VP.t5 VTAIL.t16 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=5.6121 ps=29.56 w=14.39 l=1.24
X12 VDD2.t6 VN.t3 VTAIL.t1 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X13 VDD2.t5 VN.t4 VTAIL.t0 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X14 VTAIL.t4 VN.t5 VDD2.t4 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X15 VTAIL.t17 VP.t6 VDD1.t3 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X16 VDD2.t3 VN.t6 VTAIL.t8 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=2.37435 ps=14.72 w=14.39 l=1.24
X17 VDD2.t2 VN.t7 VTAIL.t3 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=5.6121 ps=29.56 w=14.39 l=1.24
X18 VDD1.t2 VP.t7 VTAIL.t10 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=2.37435 ps=14.72 w=14.39 l=1.24
X19 VDD2.t1 VN.t8 VTAIL.t9 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=2.37435 ps=14.72 w=14.39 l=1.24
X20 VTAIL.t19 VP.t8 VDD1.t1 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X21 VTAIL.t11 VP.t9 VDD1.t0 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
X22 B.t2 B.t0 B.t1 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=5.6121 pd=29.56 as=0 ps=0 w=14.39 l=1.24
X23 VTAIL.t5 VN.t9 VDD2.t0 w_n2854_n3846# sky130_fd_pr__pfet_01v8 ad=2.37435 pd=14.72 as=2.37435 ps=14.72 w=14.39 l=1.24
R0 B.n515 B.n78 585
R1 B.n517 B.n516 585
R2 B.n518 B.n77 585
R3 B.n520 B.n519 585
R4 B.n521 B.n76 585
R5 B.n523 B.n522 585
R6 B.n524 B.n75 585
R7 B.n526 B.n525 585
R8 B.n527 B.n74 585
R9 B.n529 B.n528 585
R10 B.n530 B.n73 585
R11 B.n532 B.n531 585
R12 B.n533 B.n72 585
R13 B.n535 B.n534 585
R14 B.n536 B.n71 585
R15 B.n538 B.n537 585
R16 B.n539 B.n70 585
R17 B.n541 B.n540 585
R18 B.n542 B.n69 585
R19 B.n544 B.n543 585
R20 B.n545 B.n68 585
R21 B.n547 B.n546 585
R22 B.n548 B.n67 585
R23 B.n550 B.n549 585
R24 B.n551 B.n66 585
R25 B.n553 B.n552 585
R26 B.n554 B.n65 585
R27 B.n556 B.n555 585
R28 B.n557 B.n64 585
R29 B.n559 B.n558 585
R30 B.n560 B.n63 585
R31 B.n562 B.n561 585
R32 B.n563 B.n62 585
R33 B.n565 B.n564 585
R34 B.n566 B.n61 585
R35 B.n568 B.n567 585
R36 B.n569 B.n60 585
R37 B.n571 B.n570 585
R38 B.n572 B.n59 585
R39 B.n574 B.n573 585
R40 B.n575 B.n58 585
R41 B.n577 B.n576 585
R42 B.n578 B.n57 585
R43 B.n580 B.n579 585
R44 B.n581 B.n56 585
R45 B.n583 B.n582 585
R46 B.n584 B.n55 585
R47 B.n586 B.n585 585
R48 B.n587 B.n52 585
R49 B.n590 B.n589 585
R50 B.n591 B.n51 585
R51 B.n593 B.n592 585
R52 B.n594 B.n50 585
R53 B.n596 B.n595 585
R54 B.n597 B.n49 585
R55 B.n599 B.n598 585
R56 B.n600 B.n45 585
R57 B.n602 B.n601 585
R58 B.n603 B.n44 585
R59 B.n605 B.n604 585
R60 B.n606 B.n43 585
R61 B.n608 B.n607 585
R62 B.n609 B.n42 585
R63 B.n611 B.n610 585
R64 B.n612 B.n41 585
R65 B.n614 B.n613 585
R66 B.n615 B.n40 585
R67 B.n617 B.n616 585
R68 B.n618 B.n39 585
R69 B.n620 B.n619 585
R70 B.n621 B.n38 585
R71 B.n623 B.n622 585
R72 B.n624 B.n37 585
R73 B.n626 B.n625 585
R74 B.n627 B.n36 585
R75 B.n629 B.n628 585
R76 B.n630 B.n35 585
R77 B.n632 B.n631 585
R78 B.n633 B.n34 585
R79 B.n635 B.n634 585
R80 B.n636 B.n33 585
R81 B.n638 B.n637 585
R82 B.n639 B.n32 585
R83 B.n641 B.n640 585
R84 B.n642 B.n31 585
R85 B.n644 B.n643 585
R86 B.n645 B.n30 585
R87 B.n647 B.n646 585
R88 B.n648 B.n29 585
R89 B.n650 B.n649 585
R90 B.n651 B.n28 585
R91 B.n653 B.n652 585
R92 B.n654 B.n27 585
R93 B.n656 B.n655 585
R94 B.n657 B.n26 585
R95 B.n659 B.n658 585
R96 B.n660 B.n25 585
R97 B.n662 B.n661 585
R98 B.n663 B.n24 585
R99 B.n665 B.n664 585
R100 B.n666 B.n23 585
R101 B.n668 B.n667 585
R102 B.n669 B.n22 585
R103 B.n671 B.n670 585
R104 B.n672 B.n21 585
R105 B.n674 B.n673 585
R106 B.n675 B.n20 585
R107 B.n514 B.n513 585
R108 B.n512 B.n79 585
R109 B.n511 B.n510 585
R110 B.n509 B.n80 585
R111 B.n508 B.n507 585
R112 B.n506 B.n81 585
R113 B.n505 B.n504 585
R114 B.n503 B.n82 585
R115 B.n502 B.n501 585
R116 B.n500 B.n83 585
R117 B.n499 B.n498 585
R118 B.n497 B.n84 585
R119 B.n496 B.n495 585
R120 B.n494 B.n85 585
R121 B.n493 B.n492 585
R122 B.n491 B.n86 585
R123 B.n490 B.n489 585
R124 B.n488 B.n87 585
R125 B.n487 B.n486 585
R126 B.n485 B.n88 585
R127 B.n484 B.n483 585
R128 B.n482 B.n89 585
R129 B.n481 B.n480 585
R130 B.n479 B.n90 585
R131 B.n478 B.n477 585
R132 B.n476 B.n91 585
R133 B.n475 B.n474 585
R134 B.n473 B.n92 585
R135 B.n472 B.n471 585
R136 B.n470 B.n93 585
R137 B.n469 B.n468 585
R138 B.n467 B.n94 585
R139 B.n466 B.n465 585
R140 B.n464 B.n95 585
R141 B.n463 B.n462 585
R142 B.n461 B.n96 585
R143 B.n460 B.n459 585
R144 B.n458 B.n97 585
R145 B.n457 B.n456 585
R146 B.n455 B.n98 585
R147 B.n454 B.n453 585
R148 B.n452 B.n99 585
R149 B.n451 B.n450 585
R150 B.n449 B.n100 585
R151 B.n448 B.n447 585
R152 B.n446 B.n101 585
R153 B.n445 B.n444 585
R154 B.n443 B.n102 585
R155 B.n442 B.n441 585
R156 B.n440 B.n103 585
R157 B.n439 B.n438 585
R158 B.n437 B.n104 585
R159 B.n436 B.n435 585
R160 B.n434 B.n105 585
R161 B.n433 B.n432 585
R162 B.n431 B.n106 585
R163 B.n430 B.n429 585
R164 B.n428 B.n107 585
R165 B.n427 B.n426 585
R166 B.n425 B.n108 585
R167 B.n424 B.n423 585
R168 B.n422 B.n109 585
R169 B.n421 B.n420 585
R170 B.n419 B.n110 585
R171 B.n418 B.n417 585
R172 B.n416 B.n111 585
R173 B.n415 B.n414 585
R174 B.n413 B.n112 585
R175 B.n412 B.n411 585
R176 B.n410 B.n113 585
R177 B.n409 B.n408 585
R178 B.n407 B.n114 585
R179 B.n406 B.n405 585
R180 B.n241 B.n170 585
R181 B.n243 B.n242 585
R182 B.n244 B.n169 585
R183 B.n246 B.n245 585
R184 B.n247 B.n168 585
R185 B.n249 B.n248 585
R186 B.n250 B.n167 585
R187 B.n252 B.n251 585
R188 B.n253 B.n166 585
R189 B.n255 B.n254 585
R190 B.n256 B.n165 585
R191 B.n258 B.n257 585
R192 B.n259 B.n164 585
R193 B.n261 B.n260 585
R194 B.n262 B.n163 585
R195 B.n264 B.n263 585
R196 B.n265 B.n162 585
R197 B.n267 B.n266 585
R198 B.n268 B.n161 585
R199 B.n270 B.n269 585
R200 B.n271 B.n160 585
R201 B.n273 B.n272 585
R202 B.n274 B.n159 585
R203 B.n276 B.n275 585
R204 B.n277 B.n158 585
R205 B.n279 B.n278 585
R206 B.n280 B.n157 585
R207 B.n282 B.n281 585
R208 B.n283 B.n156 585
R209 B.n285 B.n284 585
R210 B.n286 B.n155 585
R211 B.n288 B.n287 585
R212 B.n289 B.n154 585
R213 B.n291 B.n290 585
R214 B.n292 B.n153 585
R215 B.n294 B.n293 585
R216 B.n295 B.n152 585
R217 B.n297 B.n296 585
R218 B.n298 B.n151 585
R219 B.n300 B.n299 585
R220 B.n301 B.n150 585
R221 B.n303 B.n302 585
R222 B.n304 B.n149 585
R223 B.n306 B.n305 585
R224 B.n307 B.n148 585
R225 B.n309 B.n308 585
R226 B.n310 B.n147 585
R227 B.n312 B.n311 585
R228 B.n313 B.n144 585
R229 B.n316 B.n315 585
R230 B.n317 B.n143 585
R231 B.n319 B.n318 585
R232 B.n320 B.n142 585
R233 B.n322 B.n321 585
R234 B.n323 B.n141 585
R235 B.n325 B.n324 585
R236 B.n326 B.n140 585
R237 B.n331 B.n330 585
R238 B.n332 B.n139 585
R239 B.n334 B.n333 585
R240 B.n335 B.n138 585
R241 B.n337 B.n336 585
R242 B.n338 B.n137 585
R243 B.n340 B.n339 585
R244 B.n341 B.n136 585
R245 B.n343 B.n342 585
R246 B.n344 B.n135 585
R247 B.n346 B.n345 585
R248 B.n347 B.n134 585
R249 B.n349 B.n348 585
R250 B.n350 B.n133 585
R251 B.n352 B.n351 585
R252 B.n353 B.n132 585
R253 B.n355 B.n354 585
R254 B.n356 B.n131 585
R255 B.n358 B.n357 585
R256 B.n359 B.n130 585
R257 B.n361 B.n360 585
R258 B.n362 B.n129 585
R259 B.n364 B.n363 585
R260 B.n365 B.n128 585
R261 B.n367 B.n366 585
R262 B.n368 B.n127 585
R263 B.n370 B.n369 585
R264 B.n371 B.n126 585
R265 B.n373 B.n372 585
R266 B.n374 B.n125 585
R267 B.n376 B.n375 585
R268 B.n377 B.n124 585
R269 B.n379 B.n378 585
R270 B.n380 B.n123 585
R271 B.n382 B.n381 585
R272 B.n383 B.n122 585
R273 B.n385 B.n384 585
R274 B.n386 B.n121 585
R275 B.n388 B.n387 585
R276 B.n389 B.n120 585
R277 B.n391 B.n390 585
R278 B.n392 B.n119 585
R279 B.n394 B.n393 585
R280 B.n395 B.n118 585
R281 B.n397 B.n396 585
R282 B.n398 B.n117 585
R283 B.n400 B.n399 585
R284 B.n401 B.n116 585
R285 B.n403 B.n402 585
R286 B.n404 B.n115 585
R287 B.n240 B.n239 585
R288 B.n238 B.n171 585
R289 B.n237 B.n236 585
R290 B.n235 B.n172 585
R291 B.n234 B.n233 585
R292 B.n232 B.n173 585
R293 B.n231 B.n230 585
R294 B.n229 B.n174 585
R295 B.n228 B.n227 585
R296 B.n226 B.n175 585
R297 B.n225 B.n224 585
R298 B.n223 B.n176 585
R299 B.n222 B.n221 585
R300 B.n220 B.n177 585
R301 B.n219 B.n218 585
R302 B.n217 B.n178 585
R303 B.n216 B.n215 585
R304 B.n214 B.n179 585
R305 B.n213 B.n212 585
R306 B.n211 B.n180 585
R307 B.n210 B.n209 585
R308 B.n208 B.n181 585
R309 B.n207 B.n206 585
R310 B.n205 B.n182 585
R311 B.n204 B.n203 585
R312 B.n202 B.n183 585
R313 B.n201 B.n200 585
R314 B.n199 B.n184 585
R315 B.n198 B.n197 585
R316 B.n196 B.n185 585
R317 B.n195 B.n194 585
R318 B.n193 B.n186 585
R319 B.n192 B.n191 585
R320 B.n190 B.n187 585
R321 B.n189 B.n188 585
R322 B.n2 B.n0 585
R323 B.n729 B.n1 585
R324 B.n728 B.n727 585
R325 B.n726 B.n3 585
R326 B.n725 B.n724 585
R327 B.n723 B.n4 585
R328 B.n722 B.n721 585
R329 B.n720 B.n5 585
R330 B.n719 B.n718 585
R331 B.n717 B.n6 585
R332 B.n716 B.n715 585
R333 B.n714 B.n7 585
R334 B.n713 B.n712 585
R335 B.n711 B.n8 585
R336 B.n710 B.n709 585
R337 B.n708 B.n9 585
R338 B.n707 B.n706 585
R339 B.n705 B.n10 585
R340 B.n704 B.n703 585
R341 B.n702 B.n11 585
R342 B.n701 B.n700 585
R343 B.n699 B.n12 585
R344 B.n698 B.n697 585
R345 B.n696 B.n13 585
R346 B.n695 B.n694 585
R347 B.n693 B.n14 585
R348 B.n692 B.n691 585
R349 B.n690 B.n15 585
R350 B.n689 B.n688 585
R351 B.n687 B.n16 585
R352 B.n686 B.n685 585
R353 B.n684 B.n17 585
R354 B.n683 B.n682 585
R355 B.n681 B.n18 585
R356 B.n680 B.n679 585
R357 B.n678 B.n19 585
R358 B.n677 B.n676 585
R359 B.n731 B.n730 585
R360 B.n327 B.t6 483.998
R361 B.n145 B.t9 483.998
R362 B.n46 B.t3 483.998
R363 B.n53 B.t0 483.998
R364 B.n239 B.n170 458.866
R365 B.n676 B.n675 458.866
R366 B.n405 B.n404 458.866
R367 B.n513 B.n78 458.866
R368 B.n239 B.n238 163.367
R369 B.n238 B.n237 163.367
R370 B.n237 B.n172 163.367
R371 B.n233 B.n172 163.367
R372 B.n233 B.n232 163.367
R373 B.n232 B.n231 163.367
R374 B.n231 B.n174 163.367
R375 B.n227 B.n174 163.367
R376 B.n227 B.n226 163.367
R377 B.n226 B.n225 163.367
R378 B.n225 B.n176 163.367
R379 B.n221 B.n176 163.367
R380 B.n221 B.n220 163.367
R381 B.n220 B.n219 163.367
R382 B.n219 B.n178 163.367
R383 B.n215 B.n178 163.367
R384 B.n215 B.n214 163.367
R385 B.n214 B.n213 163.367
R386 B.n213 B.n180 163.367
R387 B.n209 B.n180 163.367
R388 B.n209 B.n208 163.367
R389 B.n208 B.n207 163.367
R390 B.n207 B.n182 163.367
R391 B.n203 B.n182 163.367
R392 B.n203 B.n202 163.367
R393 B.n202 B.n201 163.367
R394 B.n201 B.n184 163.367
R395 B.n197 B.n184 163.367
R396 B.n197 B.n196 163.367
R397 B.n196 B.n195 163.367
R398 B.n195 B.n186 163.367
R399 B.n191 B.n186 163.367
R400 B.n191 B.n190 163.367
R401 B.n190 B.n189 163.367
R402 B.n189 B.n2 163.367
R403 B.n730 B.n2 163.367
R404 B.n730 B.n729 163.367
R405 B.n729 B.n728 163.367
R406 B.n728 B.n3 163.367
R407 B.n724 B.n3 163.367
R408 B.n724 B.n723 163.367
R409 B.n723 B.n722 163.367
R410 B.n722 B.n5 163.367
R411 B.n718 B.n5 163.367
R412 B.n718 B.n717 163.367
R413 B.n717 B.n716 163.367
R414 B.n716 B.n7 163.367
R415 B.n712 B.n7 163.367
R416 B.n712 B.n711 163.367
R417 B.n711 B.n710 163.367
R418 B.n710 B.n9 163.367
R419 B.n706 B.n9 163.367
R420 B.n706 B.n705 163.367
R421 B.n705 B.n704 163.367
R422 B.n704 B.n11 163.367
R423 B.n700 B.n11 163.367
R424 B.n700 B.n699 163.367
R425 B.n699 B.n698 163.367
R426 B.n698 B.n13 163.367
R427 B.n694 B.n13 163.367
R428 B.n694 B.n693 163.367
R429 B.n693 B.n692 163.367
R430 B.n692 B.n15 163.367
R431 B.n688 B.n15 163.367
R432 B.n688 B.n687 163.367
R433 B.n687 B.n686 163.367
R434 B.n686 B.n17 163.367
R435 B.n682 B.n17 163.367
R436 B.n682 B.n681 163.367
R437 B.n681 B.n680 163.367
R438 B.n680 B.n19 163.367
R439 B.n676 B.n19 163.367
R440 B.n243 B.n170 163.367
R441 B.n244 B.n243 163.367
R442 B.n245 B.n244 163.367
R443 B.n245 B.n168 163.367
R444 B.n249 B.n168 163.367
R445 B.n250 B.n249 163.367
R446 B.n251 B.n250 163.367
R447 B.n251 B.n166 163.367
R448 B.n255 B.n166 163.367
R449 B.n256 B.n255 163.367
R450 B.n257 B.n256 163.367
R451 B.n257 B.n164 163.367
R452 B.n261 B.n164 163.367
R453 B.n262 B.n261 163.367
R454 B.n263 B.n262 163.367
R455 B.n263 B.n162 163.367
R456 B.n267 B.n162 163.367
R457 B.n268 B.n267 163.367
R458 B.n269 B.n268 163.367
R459 B.n269 B.n160 163.367
R460 B.n273 B.n160 163.367
R461 B.n274 B.n273 163.367
R462 B.n275 B.n274 163.367
R463 B.n275 B.n158 163.367
R464 B.n279 B.n158 163.367
R465 B.n280 B.n279 163.367
R466 B.n281 B.n280 163.367
R467 B.n281 B.n156 163.367
R468 B.n285 B.n156 163.367
R469 B.n286 B.n285 163.367
R470 B.n287 B.n286 163.367
R471 B.n287 B.n154 163.367
R472 B.n291 B.n154 163.367
R473 B.n292 B.n291 163.367
R474 B.n293 B.n292 163.367
R475 B.n293 B.n152 163.367
R476 B.n297 B.n152 163.367
R477 B.n298 B.n297 163.367
R478 B.n299 B.n298 163.367
R479 B.n299 B.n150 163.367
R480 B.n303 B.n150 163.367
R481 B.n304 B.n303 163.367
R482 B.n305 B.n304 163.367
R483 B.n305 B.n148 163.367
R484 B.n309 B.n148 163.367
R485 B.n310 B.n309 163.367
R486 B.n311 B.n310 163.367
R487 B.n311 B.n144 163.367
R488 B.n316 B.n144 163.367
R489 B.n317 B.n316 163.367
R490 B.n318 B.n317 163.367
R491 B.n318 B.n142 163.367
R492 B.n322 B.n142 163.367
R493 B.n323 B.n322 163.367
R494 B.n324 B.n323 163.367
R495 B.n324 B.n140 163.367
R496 B.n331 B.n140 163.367
R497 B.n332 B.n331 163.367
R498 B.n333 B.n332 163.367
R499 B.n333 B.n138 163.367
R500 B.n337 B.n138 163.367
R501 B.n338 B.n337 163.367
R502 B.n339 B.n338 163.367
R503 B.n339 B.n136 163.367
R504 B.n343 B.n136 163.367
R505 B.n344 B.n343 163.367
R506 B.n345 B.n344 163.367
R507 B.n345 B.n134 163.367
R508 B.n349 B.n134 163.367
R509 B.n350 B.n349 163.367
R510 B.n351 B.n350 163.367
R511 B.n351 B.n132 163.367
R512 B.n355 B.n132 163.367
R513 B.n356 B.n355 163.367
R514 B.n357 B.n356 163.367
R515 B.n357 B.n130 163.367
R516 B.n361 B.n130 163.367
R517 B.n362 B.n361 163.367
R518 B.n363 B.n362 163.367
R519 B.n363 B.n128 163.367
R520 B.n367 B.n128 163.367
R521 B.n368 B.n367 163.367
R522 B.n369 B.n368 163.367
R523 B.n369 B.n126 163.367
R524 B.n373 B.n126 163.367
R525 B.n374 B.n373 163.367
R526 B.n375 B.n374 163.367
R527 B.n375 B.n124 163.367
R528 B.n379 B.n124 163.367
R529 B.n380 B.n379 163.367
R530 B.n381 B.n380 163.367
R531 B.n381 B.n122 163.367
R532 B.n385 B.n122 163.367
R533 B.n386 B.n385 163.367
R534 B.n387 B.n386 163.367
R535 B.n387 B.n120 163.367
R536 B.n391 B.n120 163.367
R537 B.n392 B.n391 163.367
R538 B.n393 B.n392 163.367
R539 B.n393 B.n118 163.367
R540 B.n397 B.n118 163.367
R541 B.n398 B.n397 163.367
R542 B.n399 B.n398 163.367
R543 B.n399 B.n116 163.367
R544 B.n403 B.n116 163.367
R545 B.n404 B.n403 163.367
R546 B.n405 B.n114 163.367
R547 B.n409 B.n114 163.367
R548 B.n410 B.n409 163.367
R549 B.n411 B.n410 163.367
R550 B.n411 B.n112 163.367
R551 B.n415 B.n112 163.367
R552 B.n416 B.n415 163.367
R553 B.n417 B.n416 163.367
R554 B.n417 B.n110 163.367
R555 B.n421 B.n110 163.367
R556 B.n422 B.n421 163.367
R557 B.n423 B.n422 163.367
R558 B.n423 B.n108 163.367
R559 B.n427 B.n108 163.367
R560 B.n428 B.n427 163.367
R561 B.n429 B.n428 163.367
R562 B.n429 B.n106 163.367
R563 B.n433 B.n106 163.367
R564 B.n434 B.n433 163.367
R565 B.n435 B.n434 163.367
R566 B.n435 B.n104 163.367
R567 B.n439 B.n104 163.367
R568 B.n440 B.n439 163.367
R569 B.n441 B.n440 163.367
R570 B.n441 B.n102 163.367
R571 B.n445 B.n102 163.367
R572 B.n446 B.n445 163.367
R573 B.n447 B.n446 163.367
R574 B.n447 B.n100 163.367
R575 B.n451 B.n100 163.367
R576 B.n452 B.n451 163.367
R577 B.n453 B.n452 163.367
R578 B.n453 B.n98 163.367
R579 B.n457 B.n98 163.367
R580 B.n458 B.n457 163.367
R581 B.n459 B.n458 163.367
R582 B.n459 B.n96 163.367
R583 B.n463 B.n96 163.367
R584 B.n464 B.n463 163.367
R585 B.n465 B.n464 163.367
R586 B.n465 B.n94 163.367
R587 B.n469 B.n94 163.367
R588 B.n470 B.n469 163.367
R589 B.n471 B.n470 163.367
R590 B.n471 B.n92 163.367
R591 B.n475 B.n92 163.367
R592 B.n476 B.n475 163.367
R593 B.n477 B.n476 163.367
R594 B.n477 B.n90 163.367
R595 B.n481 B.n90 163.367
R596 B.n482 B.n481 163.367
R597 B.n483 B.n482 163.367
R598 B.n483 B.n88 163.367
R599 B.n487 B.n88 163.367
R600 B.n488 B.n487 163.367
R601 B.n489 B.n488 163.367
R602 B.n489 B.n86 163.367
R603 B.n493 B.n86 163.367
R604 B.n494 B.n493 163.367
R605 B.n495 B.n494 163.367
R606 B.n495 B.n84 163.367
R607 B.n499 B.n84 163.367
R608 B.n500 B.n499 163.367
R609 B.n501 B.n500 163.367
R610 B.n501 B.n82 163.367
R611 B.n505 B.n82 163.367
R612 B.n506 B.n505 163.367
R613 B.n507 B.n506 163.367
R614 B.n507 B.n80 163.367
R615 B.n511 B.n80 163.367
R616 B.n512 B.n511 163.367
R617 B.n513 B.n512 163.367
R618 B.n675 B.n674 163.367
R619 B.n674 B.n21 163.367
R620 B.n670 B.n21 163.367
R621 B.n670 B.n669 163.367
R622 B.n669 B.n668 163.367
R623 B.n668 B.n23 163.367
R624 B.n664 B.n23 163.367
R625 B.n664 B.n663 163.367
R626 B.n663 B.n662 163.367
R627 B.n662 B.n25 163.367
R628 B.n658 B.n25 163.367
R629 B.n658 B.n657 163.367
R630 B.n657 B.n656 163.367
R631 B.n656 B.n27 163.367
R632 B.n652 B.n27 163.367
R633 B.n652 B.n651 163.367
R634 B.n651 B.n650 163.367
R635 B.n650 B.n29 163.367
R636 B.n646 B.n29 163.367
R637 B.n646 B.n645 163.367
R638 B.n645 B.n644 163.367
R639 B.n644 B.n31 163.367
R640 B.n640 B.n31 163.367
R641 B.n640 B.n639 163.367
R642 B.n639 B.n638 163.367
R643 B.n638 B.n33 163.367
R644 B.n634 B.n33 163.367
R645 B.n634 B.n633 163.367
R646 B.n633 B.n632 163.367
R647 B.n632 B.n35 163.367
R648 B.n628 B.n35 163.367
R649 B.n628 B.n627 163.367
R650 B.n627 B.n626 163.367
R651 B.n626 B.n37 163.367
R652 B.n622 B.n37 163.367
R653 B.n622 B.n621 163.367
R654 B.n621 B.n620 163.367
R655 B.n620 B.n39 163.367
R656 B.n616 B.n39 163.367
R657 B.n616 B.n615 163.367
R658 B.n615 B.n614 163.367
R659 B.n614 B.n41 163.367
R660 B.n610 B.n41 163.367
R661 B.n610 B.n609 163.367
R662 B.n609 B.n608 163.367
R663 B.n608 B.n43 163.367
R664 B.n604 B.n43 163.367
R665 B.n604 B.n603 163.367
R666 B.n603 B.n602 163.367
R667 B.n602 B.n45 163.367
R668 B.n598 B.n45 163.367
R669 B.n598 B.n597 163.367
R670 B.n597 B.n596 163.367
R671 B.n596 B.n50 163.367
R672 B.n592 B.n50 163.367
R673 B.n592 B.n591 163.367
R674 B.n591 B.n590 163.367
R675 B.n590 B.n52 163.367
R676 B.n585 B.n52 163.367
R677 B.n585 B.n584 163.367
R678 B.n584 B.n583 163.367
R679 B.n583 B.n56 163.367
R680 B.n579 B.n56 163.367
R681 B.n579 B.n578 163.367
R682 B.n578 B.n577 163.367
R683 B.n577 B.n58 163.367
R684 B.n573 B.n58 163.367
R685 B.n573 B.n572 163.367
R686 B.n572 B.n571 163.367
R687 B.n571 B.n60 163.367
R688 B.n567 B.n60 163.367
R689 B.n567 B.n566 163.367
R690 B.n566 B.n565 163.367
R691 B.n565 B.n62 163.367
R692 B.n561 B.n62 163.367
R693 B.n561 B.n560 163.367
R694 B.n560 B.n559 163.367
R695 B.n559 B.n64 163.367
R696 B.n555 B.n64 163.367
R697 B.n555 B.n554 163.367
R698 B.n554 B.n553 163.367
R699 B.n553 B.n66 163.367
R700 B.n549 B.n66 163.367
R701 B.n549 B.n548 163.367
R702 B.n548 B.n547 163.367
R703 B.n547 B.n68 163.367
R704 B.n543 B.n68 163.367
R705 B.n543 B.n542 163.367
R706 B.n542 B.n541 163.367
R707 B.n541 B.n70 163.367
R708 B.n537 B.n70 163.367
R709 B.n537 B.n536 163.367
R710 B.n536 B.n535 163.367
R711 B.n535 B.n72 163.367
R712 B.n531 B.n72 163.367
R713 B.n531 B.n530 163.367
R714 B.n530 B.n529 163.367
R715 B.n529 B.n74 163.367
R716 B.n525 B.n74 163.367
R717 B.n525 B.n524 163.367
R718 B.n524 B.n523 163.367
R719 B.n523 B.n76 163.367
R720 B.n519 B.n76 163.367
R721 B.n519 B.n518 163.367
R722 B.n518 B.n517 163.367
R723 B.n517 B.n78 163.367
R724 B.n327 B.t8 139.234
R725 B.n53 B.t1 139.234
R726 B.n145 B.t11 139.216
R727 B.n46 B.t4 139.216
R728 B.n328 B.t7 108.785
R729 B.n54 B.t2 108.785
R730 B.n146 B.t10 108.767
R731 B.n47 B.t5 108.767
R732 B.n329 B.n328 59.5399
R733 B.n314 B.n146 59.5399
R734 B.n48 B.n47 59.5399
R735 B.n588 B.n54 59.5399
R736 B.n328 B.n327 30.449
R737 B.n146 B.n145 30.449
R738 B.n47 B.n46 30.449
R739 B.n54 B.n53 30.449
R740 B.n677 B.n20 29.8151
R741 B.n406 B.n115 29.8151
R742 B.n241 B.n240 29.8151
R743 B.n515 B.n514 29.8151
R744 B B.n731 18.0485
R745 B.n673 B.n20 10.6151
R746 B.n673 B.n672 10.6151
R747 B.n672 B.n671 10.6151
R748 B.n671 B.n22 10.6151
R749 B.n667 B.n22 10.6151
R750 B.n667 B.n666 10.6151
R751 B.n666 B.n665 10.6151
R752 B.n665 B.n24 10.6151
R753 B.n661 B.n24 10.6151
R754 B.n661 B.n660 10.6151
R755 B.n660 B.n659 10.6151
R756 B.n659 B.n26 10.6151
R757 B.n655 B.n26 10.6151
R758 B.n655 B.n654 10.6151
R759 B.n654 B.n653 10.6151
R760 B.n653 B.n28 10.6151
R761 B.n649 B.n28 10.6151
R762 B.n649 B.n648 10.6151
R763 B.n648 B.n647 10.6151
R764 B.n647 B.n30 10.6151
R765 B.n643 B.n30 10.6151
R766 B.n643 B.n642 10.6151
R767 B.n642 B.n641 10.6151
R768 B.n641 B.n32 10.6151
R769 B.n637 B.n32 10.6151
R770 B.n637 B.n636 10.6151
R771 B.n636 B.n635 10.6151
R772 B.n635 B.n34 10.6151
R773 B.n631 B.n34 10.6151
R774 B.n631 B.n630 10.6151
R775 B.n630 B.n629 10.6151
R776 B.n629 B.n36 10.6151
R777 B.n625 B.n36 10.6151
R778 B.n625 B.n624 10.6151
R779 B.n624 B.n623 10.6151
R780 B.n623 B.n38 10.6151
R781 B.n619 B.n38 10.6151
R782 B.n619 B.n618 10.6151
R783 B.n618 B.n617 10.6151
R784 B.n617 B.n40 10.6151
R785 B.n613 B.n40 10.6151
R786 B.n613 B.n612 10.6151
R787 B.n612 B.n611 10.6151
R788 B.n611 B.n42 10.6151
R789 B.n607 B.n42 10.6151
R790 B.n607 B.n606 10.6151
R791 B.n606 B.n605 10.6151
R792 B.n605 B.n44 10.6151
R793 B.n601 B.n600 10.6151
R794 B.n600 B.n599 10.6151
R795 B.n599 B.n49 10.6151
R796 B.n595 B.n49 10.6151
R797 B.n595 B.n594 10.6151
R798 B.n594 B.n593 10.6151
R799 B.n593 B.n51 10.6151
R800 B.n589 B.n51 10.6151
R801 B.n587 B.n586 10.6151
R802 B.n586 B.n55 10.6151
R803 B.n582 B.n55 10.6151
R804 B.n582 B.n581 10.6151
R805 B.n581 B.n580 10.6151
R806 B.n580 B.n57 10.6151
R807 B.n576 B.n57 10.6151
R808 B.n576 B.n575 10.6151
R809 B.n575 B.n574 10.6151
R810 B.n574 B.n59 10.6151
R811 B.n570 B.n59 10.6151
R812 B.n570 B.n569 10.6151
R813 B.n569 B.n568 10.6151
R814 B.n568 B.n61 10.6151
R815 B.n564 B.n61 10.6151
R816 B.n564 B.n563 10.6151
R817 B.n563 B.n562 10.6151
R818 B.n562 B.n63 10.6151
R819 B.n558 B.n63 10.6151
R820 B.n558 B.n557 10.6151
R821 B.n557 B.n556 10.6151
R822 B.n556 B.n65 10.6151
R823 B.n552 B.n65 10.6151
R824 B.n552 B.n551 10.6151
R825 B.n551 B.n550 10.6151
R826 B.n550 B.n67 10.6151
R827 B.n546 B.n67 10.6151
R828 B.n546 B.n545 10.6151
R829 B.n545 B.n544 10.6151
R830 B.n544 B.n69 10.6151
R831 B.n540 B.n69 10.6151
R832 B.n540 B.n539 10.6151
R833 B.n539 B.n538 10.6151
R834 B.n538 B.n71 10.6151
R835 B.n534 B.n71 10.6151
R836 B.n534 B.n533 10.6151
R837 B.n533 B.n532 10.6151
R838 B.n532 B.n73 10.6151
R839 B.n528 B.n73 10.6151
R840 B.n528 B.n527 10.6151
R841 B.n527 B.n526 10.6151
R842 B.n526 B.n75 10.6151
R843 B.n522 B.n75 10.6151
R844 B.n522 B.n521 10.6151
R845 B.n521 B.n520 10.6151
R846 B.n520 B.n77 10.6151
R847 B.n516 B.n77 10.6151
R848 B.n516 B.n515 10.6151
R849 B.n407 B.n406 10.6151
R850 B.n408 B.n407 10.6151
R851 B.n408 B.n113 10.6151
R852 B.n412 B.n113 10.6151
R853 B.n413 B.n412 10.6151
R854 B.n414 B.n413 10.6151
R855 B.n414 B.n111 10.6151
R856 B.n418 B.n111 10.6151
R857 B.n419 B.n418 10.6151
R858 B.n420 B.n419 10.6151
R859 B.n420 B.n109 10.6151
R860 B.n424 B.n109 10.6151
R861 B.n425 B.n424 10.6151
R862 B.n426 B.n425 10.6151
R863 B.n426 B.n107 10.6151
R864 B.n430 B.n107 10.6151
R865 B.n431 B.n430 10.6151
R866 B.n432 B.n431 10.6151
R867 B.n432 B.n105 10.6151
R868 B.n436 B.n105 10.6151
R869 B.n437 B.n436 10.6151
R870 B.n438 B.n437 10.6151
R871 B.n438 B.n103 10.6151
R872 B.n442 B.n103 10.6151
R873 B.n443 B.n442 10.6151
R874 B.n444 B.n443 10.6151
R875 B.n444 B.n101 10.6151
R876 B.n448 B.n101 10.6151
R877 B.n449 B.n448 10.6151
R878 B.n450 B.n449 10.6151
R879 B.n450 B.n99 10.6151
R880 B.n454 B.n99 10.6151
R881 B.n455 B.n454 10.6151
R882 B.n456 B.n455 10.6151
R883 B.n456 B.n97 10.6151
R884 B.n460 B.n97 10.6151
R885 B.n461 B.n460 10.6151
R886 B.n462 B.n461 10.6151
R887 B.n462 B.n95 10.6151
R888 B.n466 B.n95 10.6151
R889 B.n467 B.n466 10.6151
R890 B.n468 B.n467 10.6151
R891 B.n468 B.n93 10.6151
R892 B.n472 B.n93 10.6151
R893 B.n473 B.n472 10.6151
R894 B.n474 B.n473 10.6151
R895 B.n474 B.n91 10.6151
R896 B.n478 B.n91 10.6151
R897 B.n479 B.n478 10.6151
R898 B.n480 B.n479 10.6151
R899 B.n480 B.n89 10.6151
R900 B.n484 B.n89 10.6151
R901 B.n485 B.n484 10.6151
R902 B.n486 B.n485 10.6151
R903 B.n486 B.n87 10.6151
R904 B.n490 B.n87 10.6151
R905 B.n491 B.n490 10.6151
R906 B.n492 B.n491 10.6151
R907 B.n492 B.n85 10.6151
R908 B.n496 B.n85 10.6151
R909 B.n497 B.n496 10.6151
R910 B.n498 B.n497 10.6151
R911 B.n498 B.n83 10.6151
R912 B.n502 B.n83 10.6151
R913 B.n503 B.n502 10.6151
R914 B.n504 B.n503 10.6151
R915 B.n504 B.n81 10.6151
R916 B.n508 B.n81 10.6151
R917 B.n509 B.n508 10.6151
R918 B.n510 B.n509 10.6151
R919 B.n510 B.n79 10.6151
R920 B.n514 B.n79 10.6151
R921 B.n242 B.n241 10.6151
R922 B.n242 B.n169 10.6151
R923 B.n246 B.n169 10.6151
R924 B.n247 B.n246 10.6151
R925 B.n248 B.n247 10.6151
R926 B.n248 B.n167 10.6151
R927 B.n252 B.n167 10.6151
R928 B.n253 B.n252 10.6151
R929 B.n254 B.n253 10.6151
R930 B.n254 B.n165 10.6151
R931 B.n258 B.n165 10.6151
R932 B.n259 B.n258 10.6151
R933 B.n260 B.n259 10.6151
R934 B.n260 B.n163 10.6151
R935 B.n264 B.n163 10.6151
R936 B.n265 B.n264 10.6151
R937 B.n266 B.n265 10.6151
R938 B.n266 B.n161 10.6151
R939 B.n270 B.n161 10.6151
R940 B.n271 B.n270 10.6151
R941 B.n272 B.n271 10.6151
R942 B.n272 B.n159 10.6151
R943 B.n276 B.n159 10.6151
R944 B.n277 B.n276 10.6151
R945 B.n278 B.n277 10.6151
R946 B.n278 B.n157 10.6151
R947 B.n282 B.n157 10.6151
R948 B.n283 B.n282 10.6151
R949 B.n284 B.n283 10.6151
R950 B.n284 B.n155 10.6151
R951 B.n288 B.n155 10.6151
R952 B.n289 B.n288 10.6151
R953 B.n290 B.n289 10.6151
R954 B.n290 B.n153 10.6151
R955 B.n294 B.n153 10.6151
R956 B.n295 B.n294 10.6151
R957 B.n296 B.n295 10.6151
R958 B.n296 B.n151 10.6151
R959 B.n300 B.n151 10.6151
R960 B.n301 B.n300 10.6151
R961 B.n302 B.n301 10.6151
R962 B.n302 B.n149 10.6151
R963 B.n306 B.n149 10.6151
R964 B.n307 B.n306 10.6151
R965 B.n308 B.n307 10.6151
R966 B.n308 B.n147 10.6151
R967 B.n312 B.n147 10.6151
R968 B.n313 B.n312 10.6151
R969 B.n315 B.n143 10.6151
R970 B.n319 B.n143 10.6151
R971 B.n320 B.n319 10.6151
R972 B.n321 B.n320 10.6151
R973 B.n321 B.n141 10.6151
R974 B.n325 B.n141 10.6151
R975 B.n326 B.n325 10.6151
R976 B.n330 B.n326 10.6151
R977 B.n334 B.n139 10.6151
R978 B.n335 B.n334 10.6151
R979 B.n336 B.n335 10.6151
R980 B.n336 B.n137 10.6151
R981 B.n340 B.n137 10.6151
R982 B.n341 B.n340 10.6151
R983 B.n342 B.n341 10.6151
R984 B.n342 B.n135 10.6151
R985 B.n346 B.n135 10.6151
R986 B.n347 B.n346 10.6151
R987 B.n348 B.n347 10.6151
R988 B.n348 B.n133 10.6151
R989 B.n352 B.n133 10.6151
R990 B.n353 B.n352 10.6151
R991 B.n354 B.n353 10.6151
R992 B.n354 B.n131 10.6151
R993 B.n358 B.n131 10.6151
R994 B.n359 B.n358 10.6151
R995 B.n360 B.n359 10.6151
R996 B.n360 B.n129 10.6151
R997 B.n364 B.n129 10.6151
R998 B.n365 B.n364 10.6151
R999 B.n366 B.n365 10.6151
R1000 B.n366 B.n127 10.6151
R1001 B.n370 B.n127 10.6151
R1002 B.n371 B.n370 10.6151
R1003 B.n372 B.n371 10.6151
R1004 B.n372 B.n125 10.6151
R1005 B.n376 B.n125 10.6151
R1006 B.n377 B.n376 10.6151
R1007 B.n378 B.n377 10.6151
R1008 B.n378 B.n123 10.6151
R1009 B.n382 B.n123 10.6151
R1010 B.n383 B.n382 10.6151
R1011 B.n384 B.n383 10.6151
R1012 B.n384 B.n121 10.6151
R1013 B.n388 B.n121 10.6151
R1014 B.n389 B.n388 10.6151
R1015 B.n390 B.n389 10.6151
R1016 B.n390 B.n119 10.6151
R1017 B.n394 B.n119 10.6151
R1018 B.n395 B.n394 10.6151
R1019 B.n396 B.n395 10.6151
R1020 B.n396 B.n117 10.6151
R1021 B.n400 B.n117 10.6151
R1022 B.n401 B.n400 10.6151
R1023 B.n402 B.n401 10.6151
R1024 B.n402 B.n115 10.6151
R1025 B.n240 B.n171 10.6151
R1026 B.n236 B.n171 10.6151
R1027 B.n236 B.n235 10.6151
R1028 B.n235 B.n234 10.6151
R1029 B.n234 B.n173 10.6151
R1030 B.n230 B.n173 10.6151
R1031 B.n230 B.n229 10.6151
R1032 B.n229 B.n228 10.6151
R1033 B.n228 B.n175 10.6151
R1034 B.n224 B.n175 10.6151
R1035 B.n224 B.n223 10.6151
R1036 B.n223 B.n222 10.6151
R1037 B.n222 B.n177 10.6151
R1038 B.n218 B.n177 10.6151
R1039 B.n218 B.n217 10.6151
R1040 B.n217 B.n216 10.6151
R1041 B.n216 B.n179 10.6151
R1042 B.n212 B.n179 10.6151
R1043 B.n212 B.n211 10.6151
R1044 B.n211 B.n210 10.6151
R1045 B.n210 B.n181 10.6151
R1046 B.n206 B.n181 10.6151
R1047 B.n206 B.n205 10.6151
R1048 B.n205 B.n204 10.6151
R1049 B.n204 B.n183 10.6151
R1050 B.n200 B.n183 10.6151
R1051 B.n200 B.n199 10.6151
R1052 B.n199 B.n198 10.6151
R1053 B.n198 B.n185 10.6151
R1054 B.n194 B.n185 10.6151
R1055 B.n194 B.n193 10.6151
R1056 B.n193 B.n192 10.6151
R1057 B.n192 B.n187 10.6151
R1058 B.n188 B.n187 10.6151
R1059 B.n188 B.n0 10.6151
R1060 B.n727 B.n1 10.6151
R1061 B.n727 B.n726 10.6151
R1062 B.n726 B.n725 10.6151
R1063 B.n725 B.n4 10.6151
R1064 B.n721 B.n4 10.6151
R1065 B.n721 B.n720 10.6151
R1066 B.n720 B.n719 10.6151
R1067 B.n719 B.n6 10.6151
R1068 B.n715 B.n6 10.6151
R1069 B.n715 B.n714 10.6151
R1070 B.n714 B.n713 10.6151
R1071 B.n713 B.n8 10.6151
R1072 B.n709 B.n8 10.6151
R1073 B.n709 B.n708 10.6151
R1074 B.n708 B.n707 10.6151
R1075 B.n707 B.n10 10.6151
R1076 B.n703 B.n10 10.6151
R1077 B.n703 B.n702 10.6151
R1078 B.n702 B.n701 10.6151
R1079 B.n701 B.n12 10.6151
R1080 B.n697 B.n12 10.6151
R1081 B.n697 B.n696 10.6151
R1082 B.n696 B.n695 10.6151
R1083 B.n695 B.n14 10.6151
R1084 B.n691 B.n14 10.6151
R1085 B.n691 B.n690 10.6151
R1086 B.n690 B.n689 10.6151
R1087 B.n689 B.n16 10.6151
R1088 B.n685 B.n16 10.6151
R1089 B.n685 B.n684 10.6151
R1090 B.n684 B.n683 10.6151
R1091 B.n683 B.n18 10.6151
R1092 B.n679 B.n18 10.6151
R1093 B.n679 B.n678 10.6151
R1094 B.n678 B.n677 10.6151
R1095 B.n601 B.n48 6.5566
R1096 B.n589 B.n588 6.5566
R1097 B.n315 B.n314 6.5566
R1098 B.n330 B.n329 6.5566
R1099 B.n48 B.n44 4.05904
R1100 B.n588 B.n587 4.05904
R1101 B.n314 B.n313 4.05904
R1102 B.n329 B.n139 4.05904
R1103 B.n731 B.n0 2.81026
R1104 B.n731 B.n1 2.81026
R1105 VP.n13 VP.t1 332.315
R1106 VP.n30 VP.t7 311.551
R1107 VP.n47 VP.t0 311.551
R1108 VP.n27 VP.t5 311.551
R1109 VP.n5 VP.t6 279.678
R1110 VP.n3 VP.t4 279.678
R1111 VP.n1 VP.t3 279.678
R1112 VP.n8 VP.t8 279.678
R1113 VP.n10 VP.t2 279.678
R1114 VP.n12 VP.t9 279.678
R1115 VP.n15 VP.n14 161.3
R1116 VP.n16 VP.n11 161.3
R1117 VP.n18 VP.n17 161.3
R1118 VP.n20 VP.n19 161.3
R1119 VP.n21 VP.n9 161.3
R1120 VP.n23 VP.n22 161.3
R1121 VP.n25 VP.n24 161.3
R1122 VP.n26 VP.n7 161.3
R1123 VP.n46 VP.n0 161.3
R1124 VP.n45 VP.n44 161.3
R1125 VP.n43 VP.n42 161.3
R1126 VP.n41 VP.n2 161.3
R1127 VP.n40 VP.n39 161.3
R1128 VP.n38 VP.n37 161.3
R1129 VP.n36 VP.n4 161.3
R1130 VP.n35 VP.n34 161.3
R1131 VP.n33 VP.n32 161.3
R1132 VP.n31 VP.n6 161.3
R1133 VP.n28 VP.n27 80.6037
R1134 VP.n48 VP.n47 80.6037
R1135 VP.n30 VP.n29 80.6037
R1136 VP.n29 VP.n28 47.7249
R1137 VP.n36 VP.n35 43.8928
R1138 VP.n42 VP.n41 43.8928
R1139 VP.n22 VP.n21 43.8928
R1140 VP.n16 VP.n15 43.8928
R1141 VP.n13 VP.n12 41.5283
R1142 VP.n31 VP.n30 39.4369
R1143 VP.n47 VP.n46 39.4369
R1144 VP.n27 VP.n26 39.4369
R1145 VP.n37 VP.n36 37.094
R1146 VP.n41 VP.n40 37.094
R1147 VP.n21 VP.n20 37.094
R1148 VP.n17 VP.n16 37.094
R1149 VP.n32 VP.n31 30.2951
R1150 VP.n46 VP.n45 30.2951
R1151 VP.n26 VP.n25 30.2951
R1152 VP.n14 VP.n13 28.9721
R1153 VP.n35 VP.n5 15.6594
R1154 VP.n42 VP.n1 15.6594
R1155 VP.n22 VP.n8 15.6594
R1156 VP.n15 VP.n12 15.6594
R1157 VP.n37 VP.n3 12.234
R1158 VP.n40 VP.n3 12.234
R1159 VP.n17 VP.n10 12.234
R1160 VP.n20 VP.n10 12.234
R1161 VP.n32 VP.n5 8.80862
R1162 VP.n45 VP.n1 8.80862
R1163 VP.n25 VP.n8 8.80862
R1164 VP.n28 VP.n7 0.285035
R1165 VP.n29 VP.n6 0.285035
R1166 VP.n48 VP.n0 0.285035
R1167 VP.n14 VP.n11 0.189894
R1168 VP.n18 VP.n11 0.189894
R1169 VP.n19 VP.n18 0.189894
R1170 VP.n19 VP.n9 0.189894
R1171 VP.n23 VP.n9 0.189894
R1172 VP.n24 VP.n23 0.189894
R1173 VP.n24 VP.n7 0.189894
R1174 VP.n33 VP.n6 0.189894
R1175 VP.n34 VP.n33 0.189894
R1176 VP.n34 VP.n4 0.189894
R1177 VP.n38 VP.n4 0.189894
R1178 VP.n39 VP.n38 0.189894
R1179 VP.n39 VP.n2 0.189894
R1180 VP.n43 VP.n2 0.189894
R1181 VP.n44 VP.n43 0.189894
R1182 VP.n44 VP.n0 0.189894
R1183 VP VP.n48 0.146778
R1184 VTAIL.n11 VTAIL.t6 58.7559
R1185 VTAIL.n17 VTAIL.t3 58.7558
R1186 VTAIL.n2 VTAIL.t13 58.7558
R1187 VTAIL.n16 VTAIL.t16 58.7558
R1188 VTAIL.n15 VTAIL.n14 56.4971
R1189 VTAIL.n13 VTAIL.n12 56.4971
R1190 VTAIL.n10 VTAIL.n9 56.4971
R1191 VTAIL.n8 VTAIL.n7 56.4971
R1192 VTAIL.n19 VTAIL.n18 56.4969
R1193 VTAIL.n1 VTAIL.n0 56.4969
R1194 VTAIL.n4 VTAIL.n3 56.4969
R1195 VTAIL.n6 VTAIL.n5 56.4969
R1196 VTAIL.n8 VTAIL.n6 27.4789
R1197 VTAIL.n17 VTAIL.n16 26.1255
R1198 VTAIL.n18 VTAIL.t1 2.25936
R1199 VTAIL.n18 VTAIL.t4 2.25936
R1200 VTAIL.n0 VTAIL.t9 2.25936
R1201 VTAIL.n0 VTAIL.t2 2.25936
R1202 VTAIL.n3 VTAIL.t15 2.25936
R1203 VTAIL.n3 VTAIL.t12 2.25936
R1204 VTAIL.n5 VTAIL.t10 2.25936
R1205 VTAIL.n5 VTAIL.t17 2.25936
R1206 VTAIL.n14 VTAIL.t14 2.25936
R1207 VTAIL.n14 VTAIL.t19 2.25936
R1208 VTAIL.n12 VTAIL.t18 2.25936
R1209 VTAIL.n12 VTAIL.t11 2.25936
R1210 VTAIL.n9 VTAIL.t0 2.25936
R1211 VTAIL.n9 VTAIL.t5 2.25936
R1212 VTAIL.n7 VTAIL.t8 2.25936
R1213 VTAIL.n7 VTAIL.t7 2.25936
R1214 VTAIL.n10 VTAIL.n8 1.35395
R1215 VTAIL.n11 VTAIL.n10 1.35395
R1216 VTAIL.n15 VTAIL.n13 1.35395
R1217 VTAIL.n16 VTAIL.n15 1.35395
R1218 VTAIL.n6 VTAIL.n4 1.35395
R1219 VTAIL.n4 VTAIL.n2 1.35395
R1220 VTAIL.n19 VTAIL.n17 1.35395
R1221 VTAIL.n13 VTAIL.n11 1.14705
R1222 VTAIL.n2 VTAIL.n1 1.14705
R1223 VTAIL VTAIL.n1 1.07378
R1224 VTAIL VTAIL.n19 0.280672
R1225 VDD1.n1 VDD1.t8 76.7882
R1226 VDD1.n3 VDD1.t2 76.788
R1227 VDD1.n5 VDD1.n4 74.1354
R1228 VDD1.n1 VDD1.n0 73.1759
R1229 VDD1.n7 VDD1.n6 73.1757
R1230 VDD1.n3 VDD1.n2 73.1757
R1231 VDD1.n7 VDD1.n5 43.8091
R1232 VDD1.n6 VDD1.t1 2.25936
R1233 VDD1.n6 VDD1.t4 2.25936
R1234 VDD1.n0 VDD1.t0 2.25936
R1235 VDD1.n0 VDD1.t7 2.25936
R1236 VDD1.n4 VDD1.t6 2.25936
R1237 VDD1.n4 VDD1.t9 2.25936
R1238 VDD1.n2 VDD1.t3 2.25936
R1239 VDD1.n2 VDD1.t5 2.25936
R1240 VDD1 VDD1.n7 0.957397
R1241 VDD1 VDD1.n1 0.397052
R1242 VDD1.n5 VDD1.n3 0.283516
R1243 VN.n6 VN.t8 332.315
R1244 VN.n28 VN.t2 332.315
R1245 VN.n20 VN.t7 311.551
R1246 VN.n42 VN.t6 311.551
R1247 VN.n5 VN.t1 279.678
R1248 VN.n3 VN.t3 279.678
R1249 VN.n1 VN.t5 279.678
R1250 VN.n27 VN.t9 279.678
R1251 VN.n25 VN.t4 279.678
R1252 VN.n23 VN.t0 279.678
R1253 VN.n41 VN.n22 161.3
R1254 VN.n40 VN.n39 161.3
R1255 VN.n38 VN.n37 161.3
R1256 VN.n36 VN.n24 161.3
R1257 VN.n35 VN.n34 161.3
R1258 VN.n33 VN.n32 161.3
R1259 VN.n31 VN.n26 161.3
R1260 VN.n30 VN.n29 161.3
R1261 VN.n19 VN.n0 161.3
R1262 VN.n18 VN.n17 161.3
R1263 VN.n16 VN.n15 161.3
R1264 VN.n14 VN.n2 161.3
R1265 VN.n13 VN.n12 161.3
R1266 VN.n11 VN.n10 161.3
R1267 VN.n9 VN.n4 161.3
R1268 VN.n8 VN.n7 161.3
R1269 VN.n43 VN.n42 80.6037
R1270 VN.n21 VN.n20 80.6037
R1271 VN VN.n43 48.0104
R1272 VN.n9 VN.n8 43.8928
R1273 VN.n15 VN.n14 43.8928
R1274 VN.n31 VN.n30 43.8928
R1275 VN.n37 VN.n36 43.8928
R1276 VN.n6 VN.n5 41.5283
R1277 VN.n28 VN.n27 41.5283
R1278 VN.n20 VN.n19 39.4369
R1279 VN.n42 VN.n41 39.4369
R1280 VN.n10 VN.n9 37.094
R1281 VN.n14 VN.n13 37.094
R1282 VN.n32 VN.n31 37.094
R1283 VN.n36 VN.n35 37.094
R1284 VN.n19 VN.n18 30.2951
R1285 VN.n41 VN.n40 30.2951
R1286 VN.n29 VN.n28 28.9721
R1287 VN.n7 VN.n6 28.9721
R1288 VN.n8 VN.n5 15.6594
R1289 VN.n15 VN.n1 15.6594
R1290 VN.n30 VN.n27 15.6594
R1291 VN.n37 VN.n23 15.6594
R1292 VN.n10 VN.n3 12.234
R1293 VN.n13 VN.n3 12.234
R1294 VN.n35 VN.n25 12.234
R1295 VN.n32 VN.n25 12.234
R1296 VN.n18 VN.n1 8.80862
R1297 VN.n40 VN.n23 8.80862
R1298 VN.n43 VN.n22 0.285035
R1299 VN.n21 VN.n0 0.285035
R1300 VN.n39 VN.n22 0.189894
R1301 VN.n39 VN.n38 0.189894
R1302 VN.n38 VN.n24 0.189894
R1303 VN.n34 VN.n24 0.189894
R1304 VN.n34 VN.n33 0.189894
R1305 VN.n33 VN.n26 0.189894
R1306 VN.n29 VN.n26 0.189894
R1307 VN.n7 VN.n4 0.189894
R1308 VN.n11 VN.n4 0.189894
R1309 VN.n12 VN.n11 0.189894
R1310 VN.n12 VN.n2 0.189894
R1311 VN.n16 VN.n2 0.189894
R1312 VN.n17 VN.n16 0.189894
R1313 VN.n17 VN.n0 0.189894
R1314 VN VN.n21 0.146778
R1315 VDD2.n1 VDD2.t1 76.788
R1316 VDD2.n4 VDD2.t3 75.4347
R1317 VDD2.n3 VDD2.n2 74.1354
R1318 VDD2 VDD2.n7 74.1326
R1319 VDD2.n6 VDD2.n5 73.1759
R1320 VDD2.n1 VDD2.n0 73.1757
R1321 VDD2.n4 VDD2.n3 42.5493
R1322 VDD2.n7 VDD2.t0 2.25936
R1323 VDD2.n7 VDD2.t7 2.25936
R1324 VDD2.n5 VDD2.t9 2.25936
R1325 VDD2.n5 VDD2.t5 2.25936
R1326 VDD2.n2 VDD2.t4 2.25936
R1327 VDD2.n2 VDD2.t2 2.25936
R1328 VDD2.n0 VDD2.t8 2.25936
R1329 VDD2.n0 VDD2.t6 2.25936
R1330 VDD2.n6 VDD2.n4 1.35395
R1331 VDD2 VDD2.n6 0.397052
R1332 VDD2.n3 VDD2.n1 0.283516
C0 VP w_n2854_n3846# 6.10093f
C1 w_n2854_n3846# VDD2 2.5081f
C2 VDD1 B 2.11363f
C3 VP VDD2 0.410343f
C4 VN VTAIL 10.2815f
C5 w_n2854_n3846# VTAIL 3.40218f
C6 VN B 0.965178f
C7 w_n2854_n3846# B 8.929621f
C8 VDD1 VN 0.150034f
C9 VP VTAIL 10.296f
C10 VDD1 w_n2854_n3846# 2.43521f
C11 VDD2 VTAIL 13.165999f
C12 VP B 1.57545f
C13 B VDD2 2.17862f
C14 VP VDD1 10.5564f
C15 VDD1 VDD2 1.30471f
C16 w_n2854_n3846# VN 5.73355f
C17 B VTAIL 3.53656f
C18 VP VN 6.83379f
C19 VN VDD2 10.301f
C20 VDD1 VTAIL 13.1274f
C21 VDD2 VSUBS 1.716866f
C22 VDD1 VSUBS 1.457181f
C23 VTAIL VSUBS 1.032807f
C24 VN VSUBS 5.73825f
C25 VP VSUBS 2.608884f
C26 B VSUBS 3.882902f
C27 w_n2854_n3846# VSUBS 0.134697p
C28 VDD2.t1 VSUBS 3.28604f
C29 VDD2.t8 VSUBS 0.310931f
C30 VDD2.t6 VSUBS 0.310931f
C31 VDD2.n0 VSUBS 2.51657f
C32 VDD2.n1 VSUBS 1.37833f
C33 VDD2.t4 VSUBS 0.310931f
C34 VDD2.t2 VSUBS 0.310931f
C35 VDD2.n2 VSUBS 2.52598f
C36 VDD2.n3 VSUBS 2.84049f
C37 VDD2.t3 VSUBS 3.27313f
C38 VDD2.n4 VSUBS 3.34773f
C39 VDD2.t9 VSUBS 0.310931f
C40 VDD2.t5 VSUBS 0.310931f
C41 VDD2.n5 VSUBS 2.51657f
C42 VDD2.n6 VSUBS 0.665744f
C43 VDD2.t0 VSUBS 0.310931f
C44 VDD2.t7 VSUBS 0.310931f
C45 VDD2.n7 VSUBS 2.52594f
C46 VN.n0 VSUBS 0.052947f
C47 VN.t5 VSUBS 1.93824f
C48 VN.n1 VSUBS 0.697912f
C49 VN.n2 VSUBS 0.039679f
C50 VN.t3 VSUBS 1.93824f
C51 VN.n3 VSUBS 0.697912f
C52 VN.n4 VSUBS 0.039679f
C53 VN.t1 VSUBS 1.93824f
C54 VN.n5 VSUBS 0.75304f
C55 VN.t8 VSUBS 2.06265f
C56 VN.n6 VSUBS 0.76216f
C57 VN.n7 VSUBS 0.209189f
C58 VN.n8 VSUBS 0.06404f
C59 VN.n9 VSUBS 0.032707f
C60 VN.n10 VSUBS 0.061662f
C61 VN.n11 VSUBS 0.039679f
C62 VN.n12 VSUBS 0.039679f
C63 VN.n13 VSUBS 0.061662f
C64 VN.n14 VSUBS 0.032707f
C65 VN.n15 VSUBS 0.06404f
C66 VN.n16 VSUBS 0.039679f
C67 VN.n17 VSUBS 0.039679f
C68 VN.n18 VSUBS 0.055923f
C69 VN.n19 VSUBS 0.032882f
C70 VN.t7 VSUBS 2.01362f
C71 VN.n20 VSUBS 0.775582f
C72 VN.n21 VSUBS 0.037161f
C73 VN.n22 VSUBS 0.052947f
C74 VN.t0 VSUBS 1.93824f
C75 VN.n23 VSUBS 0.697912f
C76 VN.n24 VSUBS 0.039679f
C77 VN.t4 VSUBS 1.93824f
C78 VN.n25 VSUBS 0.697912f
C79 VN.n26 VSUBS 0.039679f
C80 VN.t9 VSUBS 1.93824f
C81 VN.n27 VSUBS 0.75304f
C82 VN.t2 VSUBS 2.06265f
C83 VN.n28 VSUBS 0.76216f
C84 VN.n29 VSUBS 0.209189f
C85 VN.n30 VSUBS 0.06404f
C86 VN.n31 VSUBS 0.032707f
C87 VN.n32 VSUBS 0.061662f
C88 VN.n33 VSUBS 0.039679f
C89 VN.n34 VSUBS 0.039679f
C90 VN.n35 VSUBS 0.061662f
C91 VN.n36 VSUBS 0.032707f
C92 VN.n37 VSUBS 0.06404f
C93 VN.n38 VSUBS 0.039679f
C94 VN.n39 VSUBS 0.039679f
C95 VN.n40 VSUBS 0.055923f
C96 VN.n41 VSUBS 0.032882f
C97 VN.t6 VSUBS 2.01362f
C98 VN.n42 VSUBS 0.775582f
C99 VN.n43 VSUBS 2.04553f
C100 VDD1.t8 VSUBS 3.27433f
C101 VDD1.t0 VSUBS 0.309821f
C102 VDD1.t7 VSUBS 0.309821f
C103 VDD1.n0 VSUBS 2.50759f
C104 VDD1.n1 VSUBS 1.38113f
C105 VDD1.t2 VSUBS 3.27431f
C106 VDD1.t3 VSUBS 0.309821f
C107 VDD1.t5 VSUBS 0.309821f
C108 VDD1.n2 VSUBS 2.50759f
C109 VDD1.n3 VSUBS 1.37341f
C110 VDD1.t6 VSUBS 0.309821f
C111 VDD1.t9 VSUBS 0.309821f
C112 VDD1.n4 VSUBS 2.51697f
C113 VDD1.n5 VSUBS 2.92951f
C114 VDD1.t1 VSUBS 0.309821f
C115 VDD1.t4 VSUBS 0.309821f
C116 VDD1.n6 VSUBS 2.50758f
C117 VDD1.n7 VSUBS 3.33018f
C118 VTAIL.t9 VSUBS 0.314772f
C119 VTAIL.t2 VSUBS 0.314772f
C120 VTAIL.n0 VSUBS 2.39632f
C121 VTAIL.n1 VSUBS 0.829585f
C122 VTAIL.t13 VSUBS 3.14175f
C123 VTAIL.n2 VSUBS 0.967614f
C124 VTAIL.t15 VSUBS 0.314772f
C125 VTAIL.t12 VSUBS 0.314772f
C126 VTAIL.n3 VSUBS 2.39632f
C127 VTAIL.n4 VSUBS 0.873028f
C128 VTAIL.t10 VSUBS 0.314772f
C129 VTAIL.t17 VSUBS 0.314772f
C130 VTAIL.n5 VSUBS 2.39632f
C131 VTAIL.n6 VSUBS 2.47623f
C132 VTAIL.t8 VSUBS 0.314772f
C133 VTAIL.t7 VSUBS 0.314772f
C134 VTAIL.n7 VSUBS 2.39633f
C135 VTAIL.n8 VSUBS 2.47623f
C136 VTAIL.t0 VSUBS 0.314772f
C137 VTAIL.t5 VSUBS 0.314772f
C138 VTAIL.n9 VSUBS 2.39633f
C139 VTAIL.n10 VSUBS 0.873024f
C140 VTAIL.t6 VSUBS 3.14178f
C141 VTAIL.n11 VSUBS 0.96759f
C142 VTAIL.t18 VSUBS 0.314772f
C143 VTAIL.t11 VSUBS 0.314772f
C144 VTAIL.n12 VSUBS 2.39633f
C145 VTAIL.n13 VSUBS 0.85457f
C146 VTAIL.t14 VSUBS 0.314772f
C147 VTAIL.t19 VSUBS 0.314772f
C148 VTAIL.n14 VSUBS 2.39633f
C149 VTAIL.n15 VSUBS 0.873024f
C150 VTAIL.t16 VSUBS 3.14175f
C151 VTAIL.n16 VSUBS 2.46855f
C152 VTAIL.t3 VSUBS 3.14175f
C153 VTAIL.n17 VSUBS 2.46855f
C154 VTAIL.t1 VSUBS 0.314772f
C155 VTAIL.t4 VSUBS 0.314772f
C156 VTAIL.n18 VSUBS 2.39632f
C157 VTAIL.n19 VSUBS 0.777298f
C158 VP.n0 VSUBS 0.054158f
C159 VP.t3 VSUBS 1.98257f
C160 VP.n1 VSUBS 0.713874f
C161 VP.n2 VSUBS 0.040587f
C162 VP.t4 VSUBS 1.98257f
C163 VP.n3 VSUBS 0.713874f
C164 VP.n4 VSUBS 0.040587f
C165 VP.t6 VSUBS 1.98257f
C166 VP.n5 VSUBS 0.713874f
C167 VP.n6 VSUBS 0.054158f
C168 VP.n7 VSUBS 0.054158f
C169 VP.t5 VSUBS 2.05967f
C170 VP.t8 VSUBS 1.98257f
C171 VP.n8 VSUBS 0.713874f
C172 VP.n9 VSUBS 0.040587f
C173 VP.t2 VSUBS 1.98257f
C174 VP.n10 VSUBS 0.713874f
C175 VP.n11 VSUBS 0.040587f
C176 VP.t9 VSUBS 1.98257f
C177 VP.n12 VSUBS 0.770263f
C178 VP.t1 VSUBS 2.10982f
C179 VP.n13 VSUBS 0.779591f
C180 VP.n14 VSUBS 0.213974f
C181 VP.n15 VSUBS 0.065505f
C182 VP.n16 VSUBS 0.033455f
C183 VP.n17 VSUBS 0.063073f
C184 VP.n18 VSUBS 0.040587f
C185 VP.n19 VSUBS 0.040587f
C186 VP.n20 VSUBS 0.063073f
C187 VP.n21 VSUBS 0.033455f
C188 VP.n22 VSUBS 0.065505f
C189 VP.n23 VSUBS 0.040587f
C190 VP.n24 VSUBS 0.040587f
C191 VP.n25 VSUBS 0.057202f
C192 VP.n26 VSUBS 0.033634f
C193 VP.n27 VSUBS 0.793321f
C194 VP.n28 VSUBS 2.07002f
C195 VP.n29 VSUBS 2.10059f
C196 VP.t7 VSUBS 2.05967f
C197 VP.n30 VSUBS 0.793321f
C198 VP.n31 VSUBS 0.033634f
C199 VP.n32 VSUBS 0.057202f
C200 VP.n33 VSUBS 0.040587f
C201 VP.n34 VSUBS 0.040587f
C202 VP.n35 VSUBS 0.065505f
C203 VP.n36 VSUBS 0.033455f
C204 VP.n37 VSUBS 0.063073f
C205 VP.n38 VSUBS 0.040587f
C206 VP.n39 VSUBS 0.040587f
C207 VP.n40 VSUBS 0.063073f
C208 VP.n41 VSUBS 0.033455f
C209 VP.n42 VSUBS 0.065505f
C210 VP.n43 VSUBS 0.040587f
C211 VP.n44 VSUBS 0.040587f
C212 VP.n45 VSUBS 0.057202f
C213 VP.n46 VSUBS 0.033634f
C214 VP.t0 VSUBS 2.05967f
C215 VP.n47 VSUBS 0.793321f
C216 VP.n48 VSUBS 0.038011f
C217 B.n0 VSUBS 0.005598f
C218 B.n1 VSUBS 0.005598f
C219 B.n2 VSUBS 0.008852f
C220 B.n3 VSUBS 0.008852f
C221 B.n4 VSUBS 0.008852f
C222 B.n5 VSUBS 0.008852f
C223 B.n6 VSUBS 0.008852f
C224 B.n7 VSUBS 0.008852f
C225 B.n8 VSUBS 0.008852f
C226 B.n9 VSUBS 0.008852f
C227 B.n10 VSUBS 0.008852f
C228 B.n11 VSUBS 0.008852f
C229 B.n12 VSUBS 0.008852f
C230 B.n13 VSUBS 0.008852f
C231 B.n14 VSUBS 0.008852f
C232 B.n15 VSUBS 0.008852f
C233 B.n16 VSUBS 0.008852f
C234 B.n17 VSUBS 0.008852f
C235 B.n18 VSUBS 0.008852f
C236 B.n19 VSUBS 0.008852f
C237 B.n20 VSUBS 0.01996f
C238 B.n21 VSUBS 0.008852f
C239 B.n22 VSUBS 0.008852f
C240 B.n23 VSUBS 0.008852f
C241 B.n24 VSUBS 0.008852f
C242 B.n25 VSUBS 0.008852f
C243 B.n26 VSUBS 0.008852f
C244 B.n27 VSUBS 0.008852f
C245 B.n28 VSUBS 0.008852f
C246 B.n29 VSUBS 0.008852f
C247 B.n30 VSUBS 0.008852f
C248 B.n31 VSUBS 0.008852f
C249 B.n32 VSUBS 0.008852f
C250 B.n33 VSUBS 0.008852f
C251 B.n34 VSUBS 0.008852f
C252 B.n35 VSUBS 0.008852f
C253 B.n36 VSUBS 0.008852f
C254 B.n37 VSUBS 0.008852f
C255 B.n38 VSUBS 0.008852f
C256 B.n39 VSUBS 0.008852f
C257 B.n40 VSUBS 0.008852f
C258 B.n41 VSUBS 0.008852f
C259 B.n42 VSUBS 0.008852f
C260 B.n43 VSUBS 0.008852f
C261 B.n44 VSUBS 0.006119f
C262 B.n45 VSUBS 0.008852f
C263 B.t5 VSUBS 0.603622f
C264 B.t4 VSUBS 0.619203f
C265 B.t3 VSUBS 0.960104f
C266 B.n46 VSUBS 0.25204f
C267 B.n47 VSUBS 0.083866f
C268 B.n48 VSUBS 0.02051f
C269 B.n49 VSUBS 0.008852f
C270 B.n50 VSUBS 0.008852f
C271 B.n51 VSUBS 0.008852f
C272 B.n52 VSUBS 0.008852f
C273 B.t2 VSUBS 0.603606f
C274 B.t1 VSUBS 0.619188f
C275 B.t0 VSUBS 0.960104f
C276 B.n53 VSUBS 0.252054f
C277 B.n54 VSUBS 0.083882f
C278 B.n55 VSUBS 0.008852f
C279 B.n56 VSUBS 0.008852f
C280 B.n57 VSUBS 0.008852f
C281 B.n58 VSUBS 0.008852f
C282 B.n59 VSUBS 0.008852f
C283 B.n60 VSUBS 0.008852f
C284 B.n61 VSUBS 0.008852f
C285 B.n62 VSUBS 0.008852f
C286 B.n63 VSUBS 0.008852f
C287 B.n64 VSUBS 0.008852f
C288 B.n65 VSUBS 0.008852f
C289 B.n66 VSUBS 0.008852f
C290 B.n67 VSUBS 0.008852f
C291 B.n68 VSUBS 0.008852f
C292 B.n69 VSUBS 0.008852f
C293 B.n70 VSUBS 0.008852f
C294 B.n71 VSUBS 0.008852f
C295 B.n72 VSUBS 0.008852f
C296 B.n73 VSUBS 0.008852f
C297 B.n74 VSUBS 0.008852f
C298 B.n75 VSUBS 0.008852f
C299 B.n76 VSUBS 0.008852f
C300 B.n77 VSUBS 0.008852f
C301 B.n78 VSUBS 0.01996f
C302 B.n79 VSUBS 0.008852f
C303 B.n80 VSUBS 0.008852f
C304 B.n81 VSUBS 0.008852f
C305 B.n82 VSUBS 0.008852f
C306 B.n83 VSUBS 0.008852f
C307 B.n84 VSUBS 0.008852f
C308 B.n85 VSUBS 0.008852f
C309 B.n86 VSUBS 0.008852f
C310 B.n87 VSUBS 0.008852f
C311 B.n88 VSUBS 0.008852f
C312 B.n89 VSUBS 0.008852f
C313 B.n90 VSUBS 0.008852f
C314 B.n91 VSUBS 0.008852f
C315 B.n92 VSUBS 0.008852f
C316 B.n93 VSUBS 0.008852f
C317 B.n94 VSUBS 0.008852f
C318 B.n95 VSUBS 0.008852f
C319 B.n96 VSUBS 0.008852f
C320 B.n97 VSUBS 0.008852f
C321 B.n98 VSUBS 0.008852f
C322 B.n99 VSUBS 0.008852f
C323 B.n100 VSUBS 0.008852f
C324 B.n101 VSUBS 0.008852f
C325 B.n102 VSUBS 0.008852f
C326 B.n103 VSUBS 0.008852f
C327 B.n104 VSUBS 0.008852f
C328 B.n105 VSUBS 0.008852f
C329 B.n106 VSUBS 0.008852f
C330 B.n107 VSUBS 0.008852f
C331 B.n108 VSUBS 0.008852f
C332 B.n109 VSUBS 0.008852f
C333 B.n110 VSUBS 0.008852f
C334 B.n111 VSUBS 0.008852f
C335 B.n112 VSUBS 0.008852f
C336 B.n113 VSUBS 0.008852f
C337 B.n114 VSUBS 0.008852f
C338 B.n115 VSUBS 0.01996f
C339 B.n116 VSUBS 0.008852f
C340 B.n117 VSUBS 0.008852f
C341 B.n118 VSUBS 0.008852f
C342 B.n119 VSUBS 0.008852f
C343 B.n120 VSUBS 0.008852f
C344 B.n121 VSUBS 0.008852f
C345 B.n122 VSUBS 0.008852f
C346 B.n123 VSUBS 0.008852f
C347 B.n124 VSUBS 0.008852f
C348 B.n125 VSUBS 0.008852f
C349 B.n126 VSUBS 0.008852f
C350 B.n127 VSUBS 0.008852f
C351 B.n128 VSUBS 0.008852f
C352 B.n129 VSUBS 0.008852f
C353 B.n130 VSUBS 0.008852f
C354 B.n131 VSUBS 0.008852f
C355 B.n132 VSUBS 0.008852f
C356 B.n133 VSUBS 0.008852f
C357 B.n134 VSUBS 0.008852f
C358 B.n135 VSUBS 0.008852f
C359 B.n136 VSUBS 0.008852f
C360 B.n137 VSUBS 0.008852f
C361 B.n138 VSUBS 0.008852f
C362 B.n139 VSUBS 0.006119f
C363 B.n140 VSUBS 0.008852f
C364 B.n141 VSUBS 0.008852f
C365 B.n142 VSUBS 0.008852f
C366 B.n143 VSUBS 0.008852f
C367 B.n144 VSUBS 0.008852f
C368 B.t10 VSUBS 0.603622f
C369 B.t11 VSUBS 0.619203f
C370 B.t9 VSUBS 0.960104f
C371 B.n145 VSUBS 0.25204f
C372 B.n146 VSUBS 0.083866f
C373 B.n147 VSUBS 0.008852f
C374 B.n148 VSUBS 0.008852f
C375 B.n149 VSUBS 0.008852f
C376 B.n150 VSUBS 0.008852f
C377 B.n151 VSUBS 0.008852f
C378 B.n152 VSUBS 0.008852f
C379 B.n153 VSUBS 0.008852f
C380 B.n154 VSUBS 0.008852f
C381 B.n155 VSUBS 0.008852f
C382 B.n156 VSUBS 0.008852f
C383 B.n157 VSUBS 0.008852f
C384 B.n158 VSUBS 0.008852f
C385 B.n159 VSUBS 0.008852f
C386 B.n160 VSUBS 0.008852f
C387 B.n161 VSUBS 0.008852f
C388 B.n162 VSUBS 0.008852f
C389 B.n163 VSUBS 0.008852f
C390 B.n164 VSUBS 0.008852f
C391 B.n165 VSUBS 0.008852f
C392 B.n166 VSUBS 0.008852f
C393 B.n167 VSUBS 0.008852f
C394 B.n168 VSUBS 0.008852f
C395 B.n169 VSUBS 0.008852f
C396 B.n170 VSUBS 0.01996f
C397 B.n171 VSUBS 0.008852f
C398 B.n172 VSUBS 0.008852f
C399 B.n173 VSUBS 0.008852f
C400 B.n174 VSUBS 0.008852f
C401 B.n175 VSUBS 0.008852f
C402 B.n176 VSUBS 0.008852f
C403 B.n177 VSUBS 0.008852f
C404 B.n178 VSUBS 0.008852f
C405 B.n179 VSUBS 0.008852f
C406 B.n180 VSUBS 0.008852f
C407 B.n181 VSUBS 0.008852f
C408 B.n182 VSUBS 0.008852f
C409 B.n183 VSUBS 0.008852f
C410 B.n184 VSUBS 0.008852f
C411 B.n185 VSUBS 0.008852f
C412 B.n186 VSUBS 0.008852f
C413 B.n187 VSUBS 0.008852f
C414 B.n188 VSUBS 0.008852f
C415 B.n189 VSUBS 0.008852f
C416 B.n190 VSUBS 0.008852f
C417 B.n191 VSUBS 0.008852f
C418 B.n192 VSUBS 0.008852f
C419 B.n193 VSUBS 0.008852f
C420 B.n194 VSUBS 0.008852f
C421 B.n195 VSUBS 0.008852f
C422 B.n196 VSUBS 0.008852f
C423 B.n197 VSUBS 0.008852f
C424 B.n198 VSUBS 0.008852f
C425 B.n199 VSUBS 0.008852f
C426 B.n200 VSUBS 0.008852f
C427 B.n201 VSUBS 0.008852f
C428 B.n202 VSUBS 0.008852f
C429 B.n203 VSUBS 0.008852f
C430 B.n204 VSUBS 0.008852f
C431 B.n205 VSUBS 0.008852f
C432 B.n206 VSUBS 0.008852f
C433 B.n207 VSUBS 0.008852f
C434 B.n208 VSUBS 0.008852f
C435 B.n209 VSUBS 0.008852f
C436 B.n210 VSUBS 0.008852f
C437 B.n211 VSUBS 0.008852f
C438 B.n212 VSUBS 0.008852f
C439 B.n213 VSUBS 0.008852f
C440 B.n214 VSUBS 0.008852f
C441 B.n215 VSUBS 0.008852f
C442 B.n216 VSUBS 0.008852f
C443 B.n217 VSUBS 0.008852f
C444 B.n218 VSUBS 0.008852f
C445 B.n219 VSUBS 0.008852f
C446 B.n220 VSUBS 0.008852f
C447 B.n221 VSUBS 0.008852f
C448 B.n222 VSUBS 0.008852f
C449 B.n223 VSUBS 0.008852f
C450 B.n224 VSUBS 0.008852f
C451 B.n225 VSUBS 0.008852f
C452 B.n226 VSUBS 0.008852f
C453 B.n227 VSUBS 0.008852f
C454 B.n228 VSUBS 0.008852f
C455 B.n229 VSUBS 0.008852f
C456 B.n230 VSUBS 0.008852f
C457 B.n231 VSUBS 0.008852f
C458 B.n232 VSUBS 0.008852f
C459 B.n233 VSUBS 0.008852f
C460 B.n234 VSUBS 0.008852f
C461 B.n235 VSUBS 0.008852f
C462 B.n236 VSUBS 0.008852f
C463 B.n237 VSUBS 0.008852f
C464 B.n238 VSUBS 0.008852f
C465 B.n239 VSUBS 0.019094f
C466 B.n240 VSUBS 0.019094f
C467 B.n241 VSUBS 0.01996f
C468 B.n242 VSUBS 0.008852f
C469 B.n243 VSUBS 0.008852f
C470 B.n244 VSUBS 0.008852f
C471 B.n245 VSUBS 0.008852f
C472 B.n246 VSUBS 0.008852f
C473 B.n247 VSUBS 0.008852f
C474 B.n248 VSUBS 0.008852f
C475 B.n249 VSUBS 0.008852f
C476 B.n250 VSUBS 0.008852f
C477 B.n251 VSUBS 0.008852f
C478 B.n252 VSUBS 0.008852f
C479 B.n253 VSUBS 0.008852f
C480 B.n254 VSUBS 0.008852f
C481 B.n255 VSUBS 0.008852f
C482 B.n256 VSUBS 0.008852f
C483 B.n257 VSUBS 0.008852f
C484 B.n258 VSUBS 0.008852f
C485 B.n259 VSUBS 0.008852f
C486 B.n260 VSUBS 0.008852f
C487 B.n261 VSUBS 0.008852f
C488 B.n262 VSUBS 0.008852f
C489 B.n263 VSUBS 0.008852f
C490 B.n264 VSUBS 0.008852f
C491 B.n265 VSUBS 0.008852f
C492 B.n266 VSUBS 0.008852f
C493 B.n267 VSUBS 0.008852f
C494 B.n268 VSUBS 0.008852f
C495 B.n269 VSUBS 0.008852f
C496 B.n270 VSUBS 0.008852f
C497 B.n271 VSUBS 0.008852f
C498 B.n272 VSUBS 0.008852f
C499 B.n273 VSUBS 0.008852f
C500 B.n274 VSUBS 0.008852f
C501 B.n275 VSUBS 0.008852f
C502 B.n276 VSUBS 0.008852f
C503 B.n277 VSUBS 0.008852f
C504 B.n278 VSUBS 0.008852f
C505 B.n279 VSUBS 0.008852f
C506 B.n280 VSUBS 0.008852f
C507 B.n281 VSUBS 0.008852f
C508 B.n282 VSUBS 0.008852f
C509 B.n283 VSUBS 0.008852f
C510 B.n284 VSUBS 0.008852f
C511 B.n285 VSUBS 0.008852f
C512 B.n286 VSUBS 0.008852f
C513 B.n287 VSUBS 0.008852f
C514 B.n288 VSUBS 0.008852f
C515 B.n289 VSUBS 0.008852f
C516 B.n290 VSUBS 0.008852f
C517 B.n291 VSUBS 0.008852f
C518 B.n292 VSUBS 0.008852f
C519 B.n293 VSUBS 0.008852f
C520 B.n294 VSUBS 0.008852f
C521 B.n295 VSUBS 0.008852f
C522 B.n296 VSUBS 0.008852f
C523 B.n297 VSUBS 0.008852f
C524 B.n298 VSUBS 0.008852f
C525 B.n299 VSUBS 0.008852f
C526 B.n300 VSUBS 0.008852f
C527 B.n301 VSUBS 0.008852f
C528 B.n302 VSUBS 0.008852f
C529 B.n303 VSUBS 0.008852f
C530 B.n304 VSUBS 0.008852f
C531 B.n305 VSUBS 0.008852f
C532 B.n306 VSUBS 0.008852f
C533 B.n307 VSUBS 0.008852f
C534 B.n308 VSUBS 0.008852f
C535 B.n309 VSUBS 0.008852f
C536 B.n310 VSUBS 0.008852f
C537 B.n311 VSUBS 0.008852f
C538 B.n312 VSUBS 0.008852f
C539 B.n313 VSUBS 0.006119f
C540 B.n314 VSUBS 0.02051f
C541 B.n315 VSUBS 0.00716f
C542 B.n316 VSUBS 0.008852f
C543 B.n317 VSUBS 0.008852f
C544 B.n318 VSUBS 0.008852f
C545 B.n319 VSUBS 0.008852f
C546 B.n320 VSUBS 0.008852f
C547 B.n321 VSUBS 0.008852f
C548 B.n322 VSUBS 0.008852f
C549 B.n323 VSUBS 0.008852f
C550 B.n324 VSUBS 0.008852f
C551 B.n325 VSUBS 0.008852f
C552 B.n326 VSUBS 0.008852f
C553 B.t7 VSUBS 0.603606f
C554 B.t8 VSUBS 0.619188f
C555 B.t6 VSUBS 0.960104f
C556 B.n327 VSUBS 0.252054f
C557 B.n328 VSUBS 0.083882f
C558 B.n329 VSUBS 0.02051f
C559 B.n330 VSUBS 0.00716f
C560 B.n331 VSUBS 0.008852f
C561 B.n332 VSUBS 0.008852f
C562 B.n333 VSUBS 0.008852f
C563 B.n334 VSUBS 0.008852f
C564 B.n335 VSUBS 0.008852f
C565 B.n336 VSUBS 0.008852f
C566 B.n337 VSUBS 0.008852f
C567 B.n338 VSUBS 0.008852f
C568 B.n339 VSUBS 0.008852f
C569 B.n340 VSUBS 0.008852f
C570 B.n341 VSUBS 0.008852f
C571 B.n342 VSUBS 0.008852f
C572 B.n343 VSUBS 0.008852f
C573 B.n344 VSUBS 0.008852f
C574 B.n345 VSUBS 0.008852f
C575 B.n346 VSUBS 0.008852f
C576 B.n347 VSUBS 0.008852f
C577 B.n348 VSUBS 0.008852f
C578 B.n349 VSUBS 0.008852f
C579 B.n350 VSUBS 0.008852f
C580 B.n351 VSUBS 0.008852f
C581 B.n352 VSUBS 0.008852f
C582 B.n353 VSUBS 0.008852f
C583 B.n354 VSUBS 0.008852f
C584 B.n355 VSUBS 0.008852f
C585 B.n356 VSUBS 0.008852f
C586 B.n357 VSUBS 0.008852f
C587 B.n358 VSUBS 0.008852f
C588 B.n359 VSUBS 0.008852f
C589 B.n360 VSUBS 0.008852f
C590 B.n361 VSUBS 0.008852f
C591 B.n362 VSUBS 0.008852f
C592 B.n363 VSUBS 0.008852f
C593 B.n364 VSUBS 0.008852f
C594 B.n365 VSUBS 0.008852f
C595 B.n366 VSUBS 0.008852f
C596 B.n367 VSUBS 0.008852f
C597 B.n368 VSUBS 0.008852f
C598 B.n369 VSUBS 0.008852f
C599 B.n370 VSUBS 0.008852f
C600 B.n371 VSUBS 0.008852f
C601 B.n372 VSUBS 0.008852f
C602 B.n373 VSUBS 0.008852f
C603 B.n374 VSUBS 0.008852f
C604 B.n375 VSUBS 0.008852f
C605 B.n376 VSUBS 0.008852f
C606 B.n377 VSUBS 0.008852f
C607 B.n378 VSUBS 0.008852f
C608 B.n379 VSUBS 0.008852f
C609 B.n380 VSUBS 0.008852f
C610 B.n381 VSUBS 0.008852f
C611 B.n382 VSUBS 0.008852f
C612 B.n383 VSUBS 0.008852f
C613 B.n384 VSUBS 0.008852f
C614 B.n385 VSUBS 0.008852f
C615 B.n386 VSUBS 0.008852f
C616 B.n387 VSUBS 0.008852f
C617 B.n388 VSUBS 0.008852f
C618 B.n389 VSUBS 0.008852f
C619 B.n390 VSUBS 0.008852f
C620 B.n391 VSUBS 0.008852f
C621 B.n392 VSUBS 0.008852f
C622 B.n393 VSUBS 0.008852f
C623 B.n394 VSUBS 0.008852f
C624 B.n395 VSUBS 0.008852f
C625 B.n396 VSUBS 0.008852f
C626 B.n397 VSUBS 0.008852f
C627 B.n398 VSUBS 0.008852f
C628 B.n399 VSUBS 0.008852f
C629 B.n400 VSUBS 0.008852f
C630 B.n401 VSUBS 0.008852f
C631 B.n402 VSUBS 0.008852f
C632 B.n403 VSUBS 0.008852f
C633 B.n404 VSUBS 0.01996f
C634 B.n405 VSUBS 0.019094f
C635 B.n406 VSUBS 0.019094f
C636 B.n407 VSUBS 0.008852f
C637 B.n408 VSUBS 0.008852f
C638 B.n409 VSUBS 0.008852f
C639 B.n410 VSUBS 0.008852f
C640 B.n411 VSUBS 0.008852f
C641 B.n412 VSUBS 0.008852f
C642 B.n413 VSUBS 0.008852f
C643 B.n414 VSUBS 0.008852f
C644 B.n415 VSUBS 0.008852f
C645 B.n416 VSUBS 0.008852f
C646 B.n417 VSUBS 0.008852f
C647 B.n418 VSUBS 0.008852f
C648 B.n419 VSUBS 0.008852f
C649 B.n420 VSUBS 0.008852f
C650 B.n421 VSUBS 0.008852f
C651 B.n422 VSUBS 0.008852f
C652 B.n423 VSUBS 0.008852f
C653 B.n424 VSUBS 0.008852f
C654 B.n425 VSUBS 0.008852f
C655 B.n426 VSUBS 0.008852f
C656 B.n427 VSUBS 0.008852f
C657 B.n428 VSUBS 0.008852f
C658 B.n429 VSUBS 0.008852f
C659 B.n430 VSUBS 0.008852f
C660 B.n431 VSUBS 0.008852f
C661 B.n432 VSUBS 0.008852f
C662 B.n433 VSUBS 0.008852f
C663 B.n434 VSUBS 0.008852f
C664 B.n435 VSUBS 0.008852f
C665 B.n436 VSUBS 0.008852f
C666 B.n437 VSUBS 0.008852f
C667 B.n438 VSUBS 0.008852f
C668 B.n439 VSUBS 0.008852f
C669 B.n440 VSUBS 0.008852f
C670 B.n441 VSUBS 0.008852f
C671 B.n442 VSUBS 0.008852f
C672 B.n443 VSUBS 0.008852f
C673 B.n444 VSUBS 0.008852f
C674 B.n445 VSUBS 0.008852f
C675 B.n446 VSUBS 0.008852f
C676 B.n447 VSUBS 0.008852f
C677 B.n448 VSUBS 0.008852f
C678 B.n449 VSUBS 0.008852f
C679 B.n450 VSUBS 0.008852f
C680 B.n451 VSUBS 0.008852f
C681 B.n452 VSUBS 0.008852f
C682 B.n453 VSUBS 0.008852f
C683 B.n454 VSUBS 0.008852f
C684 B.n455 VSUBS 0.008852f
C685 B.n456 VSUBS 0.008852f
C686 B.n457 VSUBS 0.008852f
C687 B.n458 VSUBS 0.008852f
C688 B.n459 VSUBS 0.008852f
C689 B.n460 VSUBS 0.008852f
C690 B.n461 VSUBS 0.008852f
C691 B.n462 VSUBS 0.008852f
C692 B.n463 VSUBS 0.008852f
C693 B.n464 VSUBS 0.008852f
C694 B.n465 VSUBS 0.008852f
C695 B.n466 VSUBS 0.008852f
C696 B.n467 VSUBS 0.008852f
C697 B.n468 VSUBS 0.008852f
C698 B.n469 VSUBS 0.008852f
C699 B.n470 VSUBS 0.008852f
C700 B.n471 VSUBS 0.008852f
C701 B.n472 VSUBS 0.008852f
C702 B.n473 VSUBS 0.008852f
C703 B.n474 VSUBS 0.008852f
C704 B.n475 VSUBS 0.008852f
C705 B.n476 VSUBS 0.008852f
C706 B.n477 VSUBS 0.008852f
C707 B.n478 VSUBS 0.008852f
C708 B.n479 VSUBS 0.008852f
C709 B.n480 VSUBS 0.008852f
C710 B.n481 VSUBS 0.008852f
C711 B.n482 VSUBS 0.008852f
C712 B.n483 VSUBS 0.008852f
C713 B.n484 VSUBS 0.008852f
C714 B.n485 VSUBS 0.008852f
C715 B.n486 VSUBS 0.008852f
C716 B.n487 VSUBS 0.008852f
C717 B.n488 VSUBS 0.008852f
C718 B.n489 VSUBS 0.008852f
C719 B.n490 VSUBS 0.008852f
C720 B.n491 VSUBS 0.008852f
C721 B.n492 VSUBS 0.008852f
C722 B.n493 VSUBS 0.008852f
C723 B.n494 VSUBS 0.008852f
C724 B.n495 VSUBS 0.008852f
C725 B.n496 VSUBS 0.008852f
C726 B.n497 VSUBS 0.008852f
C727 B.n498 VSUBS 0.008852f
C728 B.n499 VSUBS 0.008852f
C729 B.n500 VSUBS 0.008852f
C730 B.n501 VSUBS 0.008852f
C731 B.n502 VSUBS 0.008852f
C732 B.n503 VSUBS 0.008852f
C733 B.n504 VSUBS 0.008852f
C734 B.n505 VSUBS 0.008852f
C735 B.n506 VSUBS 0.008852f
C736 B.n507 VSUBS 0.008852f
C737 B.n508 VSUBS 0.008852f
C738 B.n509 VSUBS 0.008852f
C739 B.n510 VSUBS 0.008852f
C740 B.n511 VSUBS 0.008852f
C741 B.n512 VSUBS 0.008852f
C742 B.n513 VSUBS 0.019094f
C743 B.n514 VSUBS 0.02024f
C744 B.n515 VSUBS 0.018815f
C745 B.n516 VSUBS 0.008852f
C746 B.n517 VSUBS 0.008852f
C747 B.n518 VSUBS 0.008852f
C748 B.n519 VSUBS 0.008852f
C749 B.n520 VSUBS 0.008852f
C750 B.n521 VSUBS 0.008852f
C751 B.n522 VSUBS 0.008852f
C752 B.n523 VSUBS 0.008852f
C753 B.n524 VSUBS 0.008852f
C754 B.n525 VSUBS 0.008852f
C755 B.n526 VSUBS 0.008852f
C756 B.n527 VSUBS 0.008852f
C757 B.n528 VSUBS 0.008852f
C758 B.n529 VSUBS 0.008852f
C759 B.n530 VSUBS 0.008852f
C760 B.n531 VSUBS 0.008852f
C761 B.n532 VSUBS 0.008852f
C762 B.n533 VSUBS 0.008852f
C763 B.n534 VSUBS 0.008852f
C764 B.n535 VSUBS 0.008852f
C765 B.n536 VSUBS 0.008852f
C766 B.n537 VSUBS 0.008852f
C767 B.n538 VSUBS 0.008852f
C768 B.n539 VSUBS 0.008852f
C769 B.n540 VSUBS 0.008852f
C770 B.n541 VSUBS 0.008852f
C771 B.n542 VSUBS 0.008852f
C772 B.n543 VSUBS 0.008852f
C773 B.n544 VSUBS 0.008852f
C774 B.n545 VSUBS 0.008852f
C775 B.n546 VSUBS 0.008852f
C776 B.n547 VSUBS 0.008852f
C777 B.n548 VSUBS 0.008852f
C778 B.n549 VSUBS 0.008852f
C779 B.n550 VSUBS 0.008852f
C780 B.n551 VSUBS 0.008852f
C781 B.n552 VSUBS 0.008852f
C782 B.n553 VSUBS 0.008852f
C783 B.n554 VSUBS 0.008852f
C784 B.n555 VSUBS 0.008852f
C785 B.n556 VSUBS 0.008852f
C786 B.n557 VSUBS 0.008852f
C787 B.n558 VSUBS 0.008852f
C788 B.n559 VSUBS 0.008852f
C789 B.n560 VSUBS 0.008852f
C790 B.n561 VSUBS 0.008852f
C791 B.n562 VSUBS 0.008852f
C792 B.n563 VSUBS 0.008852f
C793 B.n564 VSUBS 0.008852f
C794 B.n565 VSUBS 0.008852f
C795 B.n566 VSUBS 0.008852f
C796 B.n567 VSUBS 0.008852f
C797 B.n568 VSUBS 0.008852f
C798 B.n569 VSUBS 0.008852f
C799 B.n570 VSUBS 0.008852f
C800 B.n571 VSUBS 0.008852f
C801 B.n572 VSUBS 0.008852f
C802 B.n573 VSUBS 0.008852f
C803 B.n574 VSUBS 0.008852f
C804 B.n575 VSUBS 0.008852f
C805 B.n576 VSUBS 0.008852f
C806 B.n577 VSUBS 0.008852f
C807 B.n578 VSUBS 0.008852f
C808 B.n579 VSUBS 0.008852f
C809 B.n580 VSUBS 0.008852f
C810 B.n581 VSUBS 0.008852f
C811 B.n582 VSUBS 0.008852f
C812 B.n583 VSUBS 0.008852f
C813 B.n584 VSUBS 0.008852f
C814 B.n585 VSUBS 0.008852f
C815 B.n586 VSUBS 0.008852f
C816 B.n587 VSUBS 0.006119f
C817 B.n588 VSUBS 0.02051f
C818 B.n589 VSUBS 0.00716f
C819 B.n590 VSUBS 0.008852f
C820 B.n591 VSUBS 0.008852f
C821 B.n592 VSUBS 0.008852f
C822 B.n593 VSUBS 0.008852f
C823 B.n594 VSUBS 0.008852f
C824 B.n595 VSUBS 0.008852f
C825 B.n596 VSUBS 0.008852f
C826 B.n597 VSUBS 0.008852f
C827 B.n598 VSUBS 0.008852f
C828 B.n599 VSUBS 0.008852f
C829 B.n600 VSUBS 0.008852f
C830 B.n601 VSUBS 0.00716f
C831 B.n602 VSUBS 0.008852f
C832 B.n603 VSUBS 0.008852f
C833 B.n604 VSUBS 0.008852f
C834 B.n605 VSUBS 0.008852f
C835 B.n606 VSUBS 0.008852f
C836 B.n607 VSUBS 0.008852f
C837 B.n608 VSUBS 0.008852f
C838 B.n609 VSUBS 0.008852f
C839 B.n610 VSUBS 0.008852f
C840 B.n611 VSUBS 0.008852f
C841 B.n612 VSUBS 0.008852f
C842 B.n613 VSUBS 0.008852f
C843 B.n614 VSUBS 0.008852f
C844 B.n615 VSUBS 0.008852f
C845 B.n616 VSUBS 0.008852f
C846 B.n617 VSUBS 0.008852f
C847 B.n618 VSUBS 0.008852f
C848 B.n619 VSUBS 0.008852f
C849 B.n620 VSUBS 0.008852f
C850 B.n621 VSUBS 0.008852f
C851 B.n622 VSUBS 0.008852f
C852 B.n623 VSUBS 0.008852f
C853 B.n624 VSUBS 0.008852f
C854 B.n625 VSUBS 0.008852f
C855 B.n626 VSUBS 0.008852f
C856 B.n627 VSUBS 0.008852f
C857 B.n628 VSUBS 0.008852f
C858 B.n629 VSUBS 0.008852f
C859 B.n630 VSUBS 0.008852f
C860 B.n631 VSUBS 0.008852f
C861 B.n632 VSUBS 0.008852f
C862 B.n633 VSUBS 0.008852f
C863 B.n634 VSUBS 0.008852f
C864 B.n635 VSUBS 0.008852f
C865 B.n636 VSUBS 0.008852f
C866 B.n637 VSUBS 0.008852f
C867 B.n638 VSUBS 0.008852f
C868 B.n639 VSUBS 0.008852f
C869 B.n640 VSUBS 0.008852f
C870 B.n641 VSUBS 0.008852f
C871 B.n642 VSUBS 0.008852f
C872 B.n643 VSUBS 0.008852f
C873 B.n644 VSUBS 0.008852f
C874 B.n645 VSUBS 0.008852f
C875 B.n646 VSUBS 0.008852f
C876 B.n647 VSUBS 0.008852f
C877 B.n648 VSUBS 0.008852f
C878 B.n649 VSUBS 0.008852f
C879 B.n650 VSUBS 0.008852f
C880 B.n651 VSUBS 0.008852f
C881 B.n652 VSUBS 0.008852f
C882 B.n653 VSUBS 0.008852f
C883 B.n654 VSUBS 0.008852f
C884 B.n655 VSUBS 0.008852f
C885 B.n656 VSUBS 0.008852f
C886 B.n657 VSUBS 0.008852f
C887 B.n658 VSUBS 0.008852f
C888 B.n659 VSUBS 0.008852f
C889 B.n660 VSUBS 0.008852f
C890 B.n661 VSUBS 0.008852f
C891 B.n662 VSUBS 0.008852f
C892 B.n663 VSUBS 0.008852f
C893 B.n664 VSUBS 0.008852f
C894 B.n665 VSUBS 0.008852f
C895 B.n666 VSUBS 0.008852f
C896 B.n667 VSUBS 0.008852f
C897 B.n668 VSUBS 0.008852f
C898 B.n669 VSUBS 0.008852f
C899 B.n670 VSUBS 0.008852f
C900 B.n671 VSUBS 0.008852f
C901 B.n672 VSUBS 0.008852f
C902 B.n673 VSUBS 0.008852f
C903 B.n674 VSUBS 0.008852f
C904 B.n675 VSUBS 0.01996f
C905 B.n676 VSUBS 0.019094f
C906 B.n677 VSUBS 0.019094f
C907 B.n678 VSUBS 0.008852f
C908 B.n679 VSUBS 0.008852f
C909 B.n680 VSUBS 0.008852f
C910 B.n681 VSUBS 0.008852f
C911 B.n682 VSUBS 0.008852f
C912 B.n683 VSUBS 0.008852f
C913 B.n684 VSUBS 0.008852f
C914 B.n685 VSUBS 0.008852f
C915 B.n686 VSUBS 0.008852f
C916 B.n687 VSUBS 0.008852f
C917 B.n688 VSUBS 0.008852f
C918 B.n689 VSUBS 0.008852f
C919 B.n690 VSUBS 0.008852f
C920 B.n691 VSUBS 0.008852f
C921 B.n692 VSUBS 0.008852f
C922 B.n693 VSUBS 0.008852f
C923 B.n694 VSUBS 0.008852f
C924 B.n695 VSUBS 0.008852f
C925 B.n696 VSUBS 0.008852f
C926 B.n697 VSUBS 0.008852f
C927 B.n698 VSUBS 0.008852f
C928 B.n699 VSUBS 0.008852f
C929 B.n700 VSUBS 0.008852f
C930 B.n701 VSUBS 0.008852f
C931 B.n702 VSUBS 0.008852f
C932 B.n703 VSUBS 0.008852f
C933 B.n704 VSUBS 0.008852f
C934 B.n705 VSUBS 0.008852f
C935 B.n706 VSUBS 0.008852f
C936 B.n707 VSUBS 0.008852f
C937 B.n708 VSUBS 0.008852f
C938 B.n709 VSUBS 0.008852f
C939 B.n710 VSUBS 0.008852f
C940 B.n711 VSUBS 0.008852f
C941 B.n712 VSUBS 0.008852f
C942 B.n713 VSUBS 0.008852f
C943 B.n714 VSUBS 0.008852f
C944 B.n715 VSUBS 0.008852f
C945 B.n716 VSUBS 0.008852f
C946 B.n717 VSUBS 0.008852f
C947 B.n718 VSUBS 0.008852f
C948 B.n719 VSUBS 0.008852f
C949 B.n720 VSUBS 0.008852f
C950 B.n721 VSUBS 0.008852f
C951 B.n722 VSUBS 0.008852f
C952 B.n723 VSUBS 0.008852f
C953 B.n724 VSUBS 0.008852f
C954 B.n725 VSUBS 0.008852f
C955 B.n726 VSUBS 0.008852f
C956 B.n727 VSUBS 0.008852f
C957 B.n728 VSUBS 0.008852f
C958 B.n729 VSUBS 0.008852f
C959 B.n730 VSUBS 0.008852f
C960 B.n731 VSUBS 0.020045f
.ends

