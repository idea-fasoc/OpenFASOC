* NGSPICE file created from diff_pair_sample_1640.ext - technology: sky130A

.subckt diff_pair_sample_1640 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t1 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X1 VTAIL.t2 VN.t0 VDD2.t9 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X2 B.t11 B.t9 B.t10 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=0 ps=0 w=10.8 l=3.93
X3 VDD2.t8 VN.t1 VTAIL.t6 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X4 VTAIL.t16 VP.t1 VDD1.t0 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X5 VTAIL.t1 VN.t2 VDD2.t7 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X6 VDD2.t6 VN.t3 VTAIL.t3 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=1.782 ps=11.13 w=10.8 l=3.93
X7 B.t8 B.t6 B.t7 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=0 ps=0 w=10.8 l=3.93
X8 VDD1.t3 VP.t2 VTAIL.t15 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=1.782 ps=11.13 w=10.8 l=3.93
X9 VDD2.t5 VN.t4 VTAIL.t0 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=4.212 ps=22.38 w=10.8 l=3.93
X10 B.t5 B.t3 B.t4 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=0 ps=0 w=10.8 l=3.93
X11 VDD1.t2 VP.t3 VTAIL.t14 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=1.782 ps=11.13 w=10.8 l=3.93
X12 VDD1.t5 VP.t4 VTAIL.t13 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=4.212 ps=22.38 w=10.8 l=3.93
X13 VTAIL.t5 VN.t5 VDD2.t4 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X14 VDD1.t4 VP.t5 VTAIL.t12 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X15 VDD2.t3 VN.t6 VTAIL.t18 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X16 VDD2.t2 VN.t7 VTAIL.t4 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=4.212 ps=22.38 w=10.8 l=3.93
X17 VDD1.t9 VP.t6 VTAIL.t11 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X18 VDD2.t1 VN.t8 VTAIL.t19 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=1.782 ps=11.13 w=10.8 l=3.93
X19 VDD1.t8 VP.t7 VTAIL.t10 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=4.212 ps=22.38 w=10.8 l=3.93
X20 VTAIL.t9 VP.t8 VDD1.t7 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X21 VTAIL.t7 VN.t9 VDD2.t0 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X22 VTAIL.t8 VP.t9 VDD1.t6 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=1.782 pd=11.13 as=1.782 ps=11.13 w=10.8 l=3.93
X23 B.t2 B.t0 B.t1 w_n6082_n3128# sky130_fd_pr__pfet_01v8 ad=4.212 pd=22.38 as=0 ps=0 w=10.8 l=3.93
R0 VP.n35 VP.n32 161.3
R1 VP.n37 VP.n36 161.3
R2 VP.n38 VP.n31 161.3
R3 VP.n40 VP.n39 161.3
R4 VP.n41 VP.n30 161.3
R5 VP.n43 VP.n42 161.3
R6 VP.n44 VP.n29 161.3
R7 VP.n46 VP.n45 161.3
R8 VP.n47 VP.n28 161.3
R9 VP.n49 VP.n48 161.3
R10 VP.n50 VP.n27 161.3
R11 VP.n52 VP.n51 161.3
R12 VP.n53 VP.n26 161.3
R13 VP.n55 VP.n54 161.3
R14 VP.n56 VP.n25 161.3
R15 VP.n58 VP.n57 161.3
R16 VP.n59 VP.n24 161.3
R17 VP.n62 VP.n61 161.3
R18 VP.n63 VP.n23 161.3
R19 VP.n65 VP.n64 161.3
R20 VP.n66 VP.n22 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n69 VP.n21 161.3
R23 VP.n71 VP.n70 161.3
R24 VP.n72 VP.n20 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n131 VP.n130 161.3
R27 VP.n129 VP.n1 161.3
R28 VP.n128 VP.n127 161.3
R29 VP.n126 VP.n2 161.3
R30 VP.n125 VP.n124 161.3
R31 VP.n123 VP.n3 161.3
R32 VP.n122 VP.n121 161.3
R33 VP.n120 VP.n4 161.3
R34 VP.n119 VP.n118 161.3
R35 VP.n116 VP.n5 161.3
R36 VP.n115 VP.n114 161.3
R37 VP.n113 VP.n6 161.3
R38 VP.n112 VP.n111 161.3
R39 VP.n110 VP.n7 161.3
R40 VP.n109 VP.n108 161.3
R41 VP.n107 VP.n8 161.3
R42 VP.n106 VP.n105 161.3
R43 VP.n104 VP.n9 161.3
R44 VP.n103 VP.n102 161.3
R45 VP.n101 VP.n10 161.3
R46 VP.n100 VP.n99 161.3
R47 VP.n98 VP.n11 161.3
R48 VP.n97 VP.n96 161.3
R49 VP.n95 VP.n12 161.3
R50 VP.n94 VP.n93 161.3
R51 VP.n92 VP.n13 161.3
R52 VP.n90 VP.n89 161.3
R53 VP.n88 VP.n14 161.3
R54 VP.n87 VP.n86 161.3
R55 VP.n85 VP.n15 161.3
R56 VP.n84 VP.n83 161.3
R57 VP.n82 VP.n16 161.3
R58 VP.n81 VP.n80 161.3
R59 VP.n79 VP.n17 161.3
R60 VP.n78 VP.n77 161.3
R61 VP.n33 VP.t3 98.442
R62 VP.n76 VP.n18 88.9173
R63 VP.n132 VP.n0 88.9173
R64 VP.n75 VP.n19 88.9173
R65 VP.n104 VP.t5 66.2295
R66 VP.n18 VP.t2 66.2295
R67 VP.n91 VP.t8 66.2295
R68 VP.n117 VP.t9 66.2295
R69 VP.n0 VP.t4 66.2295
R70 VP.n47 VP.t6 66.2295
R71 VP.n19 VP.t7 66.2295
R72 VP.n60 VP.t1 66.2295
R73 VP.n34 VP.t0 66.2295
R74 VP.n34 VP.n33 62.2666
R75 VP.n76 VP.n75 59.4915
R76 VP.n98 VP.n97 53.0692
R77 VP.n111 VP.n110 53.0692
R78 VP.n54 VP.n53 53.0692
R79 VP.n41 VP.n40 53.0692
R80 VP.n85 VP.n84 51.1217
R81 VP.n124 VP.n123 51.1217
R82 VP.n67 VP.n66 51.1217
R83 VP.n84 VP.n16 29.6995
R84 VP.n124 VP.n2 29.6995
R85 VP.n67 VP.n21 29.6995
R86 VP.n99 VP.n98 27.752
R87 VP.n110 VP.n109 27.752
R88 VP.n53 VP.n52 27.752
R89 VP.n42 VP.n41 27.752
R90 VP.n79 VP.n78 24.3439
R91 VP.n80 VP.n79 24.3439
R92 VP.n80 VP.n16 24.3439
R93 VP.n86 VP.n85 24.3439
R94 VP.n86 VP.n14 24.3439
R95 VP.n90 VP.n14 24.3439
R96 VP.n93 VP.n92 24.3439
R97 VP.n93 VP.n12 24.3439
R98 VP.n97 VP.n12 24.3439
R99 VP.n99 VP.n10 24.3439
R100 VP.n103 VP.n10 24.3439
R101 VP.n104 VP.n103 24.3439
R102 VP.n105 VP.n104 24.3439
R103 VP.n105 VP.n8 24.3439
R104 VP.n109 VP.n8 24.3439
R105 VP.n111 VP.n6 24.3439
R106 VP.n115 VP.n6 24.3439
R107 VP.n116 VP.n115 24.3439
R108 VP.n118 VP.n4 24.3439
R109 VP.n122 VP.n4 24.3439
R110 VP.n123 VP.n122 24.3439
R111 VP.n128 VP.n2 24.3439
R112 VP.n129 VP.n128 24.3439
R113 VP.n130 VP.n129 24.3439
R114 VP.n71 VP.n21 24.3439
R115 VP.n72 VP.n71 24.3439
R116 VP.n73 VP.n72 24.3439
R117 VP.n54 VP.n25 24.3439
R118 VP.n58 VP.n25 24.3439
R119 VP.n59 VP.n58 24.3439
R120 VP.n61 VP.n23 24.3439
R121 VP.n65 VP.n23 24.3439
R122 VP.n66 VP.n65 24.3439
R123 VP.n42 VP.n29 24.3439
R124 VP.n46 VP.n29 24.3439
R125 VP.n47 VP.n46 24.3439
R126 VP.n48 VP.n47 24.3439
R127 VP.n48 VP.n27 24.3439
R128 VP.n52 VP.n27 24.3439
R129 VP.n36 VP.n35 24.3439
R130 VP.n36 VP.n31 24.3439
R131 VP.n40 VP.n31 24.3439
R132 VP.n92 VP.n91 12.6591
R133 VP.n117 VP.n116 12.6591
R134 VP.n60 VP.n59 12.6591
R135 VP.n35 VP.n34 12.6591
R136 VP.n91 VP.n90 11.6853
R137 VP.n118 VP.n117 11.6853
R138 VP.n61 VP.n60 11.6853
R139 VP.n33 VP.n32 2.52182
R140 VP.n78 VP.n18 0.974237
R141 VP.n130 VP.n0 0.974237
R142 VP.n73 VP.n19 0.974237
R143 VP.n75 VP.n74 0.355081
R144 VP.n77 VP.n76 0.355081
R145 VP.n132 VP.n131 0.355081
R146 VP VP.n132 0.26685
R147 VP.n37 VP.n32 0.189894
R148 VP.n38 VP.n37 0.189894
R149 VP.n39 VP.n38 0.189894
R150 VP.n39 VP.n30 0.189894
R151 VP.n43 VP.n30 0.189894
R152 VP.n44 VP.n43 0.189894
R153 VP.n45 VP.n44 0.189894
R154 VP.n45 VP.n28 0.189894
R155 VP.n49 VP.n28 0.189894
R156 VP.n50 VP.n49 0.189894
R157 VP.n51 VP.n50 0.189894
R158 VP.n51 VP.n26 0.189894
R159 VP.n55 VP.n26 0.189894
R160 VP.n56 VP.n55 0.189894
R161 VP.n57 VP.n56 0.189894
R162 VP.n57 VP.n24 0.189894
R163 VP.n62 VP.n24 0.189894
R164 VP.n63 VP.n62 0.189894
R165 VP.n64 VP.n63 0.189894
R166 VP.n64 VP.n22 0.189894
R167 VP.n68 VP.n22 0.189894
R168 VP.n69 VP.n68 0.189894
R169 VP.n70 VP.n69 0.189894
R170 VP.n70 VP.n20 0.189894
R171 VP.n74 VP.n20 0.189894
R172 VP.n77 VP.n17 0.189894
R173 VP.n81 VP.n17 0.189894
R174 VP.n82 VP.n81 0.189894
R175 VP.n83 VP.n82 0.189894
R176 VP.n83 VP.n15 0.189894
R177 VP.n87 VP.n15 0.189894
R178 VP.n88 VP.n87 0.189894
R179 VP.n89 VP.n88 0.189894
R180 VP.n89 VP.n13 0.189894
R181 VP.n94 VP.n13 0.189894
R182 VP.n95 VP.n94 0.189894
R183 VP.n96 VP.n95 0.189894
R184 VP.n96 VP.n11 0.189894
R185 VP.n100 VP.n11 0.189894
R186 VP.n101 VP.n100 0.189894
R187 VP.n102 VP.n101 0.189894
R188 VP.n102 VP.n9 0.189894
R189 VP.n106 VP.n9 0.189894
R190 VP.n107 VP.n106 0.189894
R191 VP.n108 VP.n107 0.189894
R192 VP.n108 VP.n7 0.189894
R193 VP.n112 VP.n7 0.189894
R194 VP.n113 VP.n112 0.189894
R195 VP.n114 VP.n113 0.189894
R196 VP.n114 VP.n5 0.189894
R197 VP.n119 VP.n5 0.189894
R198 VP.n120 VP.n119 0.189894
R199 VP.n121 VP.n120 0.189894
R200 VP.n121 VP.n3 0.189894
R201 VP.n125 VP.n3 0.189894
R202 VP.n126 VP.n125 0.189894
R203 VP.n127 VP.n126 0.189894
R204 VP.n127 VP.n1 0.189894
R205 VP.n131 VP.n1 0.189894
R206 VDD1.n52 VDD1.n0 756.745
R207 VDD1.n111 VDD1.n59 756.745
R208 VDD1.n53 VDD1.n52 585
R209 VDD1.n51 VDD1.n50 585
R210 VDD1.n4 VDD1.n3 585
R211 VDD1.n45 VDD1.n44 585
R212 VDD1.n43 VDD1.n42 585
R213 VDD1.n41 VDD1.n7 585
R214 VDD1.n11 VDD1.n8 585
R215 VDD1.n36 VDD1.n35 585
R216 VDD1.n34 VDD1.n33 585
R217 VDD1.n13 VDD1.n12 585
R218 VDD1.n28 VDD1.n27 585
R219 VDD1.n26 VDD1.n25 585
R220 VDD1.n17 VDD1.n16 585
R221 VDD1.n20 VDD1.n19 585
R222 VDD1.n78 VDD1.n77 585
R223 VDD1.n75 VDD1.n74 585
R224 VDD1.n84 VDD1.n83 585
R225 VDD1.n86 VDD1.n85 585
R226 VDD1.n71 VDD1.n70 585
R227 VDD1.n92 VDD1.n91 585
R228 VDD1.n95 VDD1.n94 585
R229 VDD1.n93 VDD1.n67 585
R230 VDD1.n100 VDD1.n66 585
R231 VDD1.n102 VDD1.n101 585
R232 VDD1.n104 VDD1.n103 585
R233 VDD1.n63 VDD1.n62 585
R234 VDD1.n110 VDD1.n109 585
R235 VDD1.n112 VDD1.n111 585
R236 VDD1.t2 VDD1.n18 329.038
R237 VDD1.t3 VDD1.n76 329.038
R238 VDD1.n52 VDD1.n51 171.744
R239 VDD1.n51 VDD1.n3 171.744
R240 VDD1.n44 VDD1.n3 171.744
R241 VDD1.n44 VDD1.n43 171.744
R242 VDD1.n43 VDD1.n7 171.744
R243 VDD1.n11 VDD1.n7 171.744
R244 VDD1.n35 VDD1.n11 171.744
R245 VDD1.n35 VDD1.n34 171.744
R246 VDD1.n34 VDD1.n12 171.744
R247 VDD1.n27 VDD1.n12 171.744
R248 VDD1.n27 VDD1.n26 171.744
R249 VDD1.n26 VDD1.n16 171.744
R250 VDD1.n19 VDD1.n16 171.744
R251 VDD1.n77 VDD1.n74 171.744
R252 VDD1.n84 VDD1.n74 171.744
R253 VDD1.n85 VDD1.n84 171.744
R254 VDD1.n85 VDD1.n70 171.744
R255 VDD1.n92 VDD1.n70 171.744
R256 VDD1.n94 VDD1.n92 171.744
R257 VDD1.n94 VDD1.n93 171.744
R258 VDD1.n93 VDD1.n66 171.744
R259 VDD1.n102 VDD1.n66 171.744
R260 VDD1.n103 VDD1.n102 171.744
R261 VDD1.n103 VDD1.n62 171.744
R262 VDD1.n110 VDD1.n62 171.744
R263 VDD1.n111 VDD1.n110 171.744
R264 VDD1.n19 VDD1.t2 85.8723
R265 VDD1.n77 VDD1.t3 85.8723
R266 VDD1.n119 VDD1.n118 80.8922
R267 VDD1.n58 VDD1.n57 78.1934
R268 VDD1.n121 VDD1.n120 78.1932
R269 VDD1.n117 VDD1.n116 78.1932
R270 VDD1.n58 VDD1.n56 54.8638
R271 VDD1.n117 VDD1.n115 54.8638
R272 VDD1.n121 VDD1.n119 52.8888
R273 VDD1.n42 VDD1.n41 13.1884
R274 VDD1.n101 VDD1.n100 13.1884
R275 VDD1.n45 VDD1.n6 12.8005
R276 VDD1.n40 VDD1.n8 12.8005
R277 VDD1.n99 VDD1.n67 12.8005
R278 VDD1.n104 VDD1.n65 12.8005
R279 VDD1.n46 VDD1.n4 12.0247
R280 VDD1.n37 VDD1.n36 12.0247
R281 VDD1.n96 VDD1.n95 12.0247
R282 VDD1.n105 VDD1.n63 12.0247
R283 VDD1.n50 VDD1.n49 11.249
R284 VDD1.n33 VDD1.n10 11.249
R285 VDD1.n91 VDD1.n69 11.249
R286 VDD1.n109 VDD1.n108 11.249
R287 VDD1.n20 VDD1.n18 10.7239
R288 VDD1.n78 VDD1.n76 10.7239
R289 VDD1.n53 VDD1.n2 10.4732
R290 VDD1.n32 VDD1.n13 10.4732
R291 VDD1.n90 VDD1.n71 10.4732
R292 VDD1.n112 VDD1.n61 10.4732
R293 VDD1.n54 VDD1.n0 9.69747
R294 VDD1.n29 VDD1.n28 9.69747
R295 VDD1.n87 VDD1.n86 9.69747
R296 VDD1.n113 VDD1.n59 9.69747
R297 VDD1.n56 VDD1.n55 9.45567
R298 VDD1.n115 VDD1.n114 9.45567
R299 VDD1.n22 VDD1.n21 9.3005
R300 VDD1.n24 VDD1.n23 9.3005
R301 VDD1.n15 VDD1.n14 9.3005
R302 VDD1.n30 VDD1.n29 9.3005
R303 VDD1.n32 VDD1.n31 9.3005
R304 VDD1.n10 VDD1.n9 9.3005
R305 VDD1.n38 VDD1.n37 9.3005
R306 VDD1.n40 VDD1.n39 9.3005
R307 VDD1.n55 VDD1.n54 9.3005
R308 VDD1.n2 VDD1.n1 9.3005
R309 VDD1.n49 VDD1.n48 9.3005
R310 VDD1.n47 VDD1.n46 9.3005
R311 VDD1.n6 VDD1.n5 9.3005
R312 VDD1.n114 VDD1.n113 9.3005
R313 VDD1.n61 VDD1.n60 9.3005
R314 VDD1.n108 VDD1.n107 9.3005
R315 VDD1.n106 VDD1.n105 9.3005
R316 VDD1.n65 VDD1.n64 9.3005
R317 VDD1.n80 VDD1.n79 9.3005
R318 VDD1.n82 VDD1.n81 9.3005
R319 VDD1.n73 VDD1.n72 9.3005
R320 VDD1.n88 VDD1.n87 9.3005
R321 VDD1.n90 VDD1.n89 9.3005
R322 VDD1.n69 VDD1.n68 9.3005
R323 VDD1.n97 VDD1.n96 9.3005
R324 VDD1.n99 VDD1.n98 9.3005
R325 VDD1.n25 VDD1.n15 8.92171
R326 VDD1.n83 VDD1.n73 8.92171
R327 VDD1.n24 VDD1.n17 8.14595
R328 VDD1.n82 VDD1.n75 8.14595
R329 VDD1.n21 VDD1.n20 7.3702
R330 VDD1.n79 VDD1.n78 7.3702
R331 VDD1.n21 VDD1.n17 5.81868
R332 VDD1.n79 VDD1.n75 5.81868
R333 VDD1.n25 VDD1.n24 5.04292
R334 VDD1.n83 VDD1.n82 5.04292
R335 VDD1.n56 VDD1.n0 4.26717
R336 VDD1.n28 VDD1.n15 4.26717
R337 VDD1.n86 VDD1.n73 4.26717
R338 VDD1.n115 VDD1.n59 4.26717
R339 VDD1.n54 VDD1.n53 3.49141
R340 VDD1.n29 VDD1.n13 3.49141
R341 VDD1.n87 VDD1.n71 3.49141
R342 VDD1.n113 VDD1.n112 3.49141
R343 VDD1.n120 VDD1.t0 3.01022
R344 VDD1.n120 VDD1.t8 3.01022
R345 VDD1.n57 VDD1.t1 3.01022
R346 VDD1.n57 VDD1.t9 3.01022
R347 VDD1.n118 VDD1.t6 3.01022
R348 VDD1.n118 VDD1.t5 3.01022
R349 VDD1.n116 VDD1.t7 3.01022
R350 VDD1.n116 VDD1.t4 3.01022
R351 VDD1.n50 VDD1.n2 2.71565
R352 VDD1.n33 VDD1.n32 2.71565
R353 VDD1.n91 VDD1.n90 2.71565
R354 VDD1.n109 VDD1.n61 2.71565
R355 VDD1 VDD1.n121 2.69662
R356 VDD1.n22 VDD1.n18 2.41282
R357 VDD1.n80 VDD1.n76 2.41282
R358 VDD1.n49 VDD1.n4 1.93989
R359 VDD1.n36 VDD1.n10 1.93989
R360 VDD1.n95 VDD1.n69 1.93989
R361 VDD1.n108 VDD1.n63 1.93989
R362 VDD1.n46 VDD1.n45 1.16414
R363 VDD1.n37 VDD1.n8 1.16414
R364 VDD1.n96 VDD1.n67 1.16414
R365 VDD1.n105 VDD1.n104 1.16414
R366 VDD1 VDD1.n58 0.976793
R367 VDD1.n119 VDD1.n117 0.863257
R368 VDD1.n42 VDD1.n6 0.388379
R369 VDD1.n41 VDD1.n40 0.388379
R370 VDD1.n100 VDD1.n99 0.388379
R371 VDD1.n101 VDD1.n65 0.388379
R372 VDD1.n55 VDD1.n1 0.155672
R373 VDD1.n48 VDD1.n1 0.155672
R374 VDD1.n48 VDD1.n47 0.155672
R375 VDD1.n47 VDD1.n5 0.155672
R376 VDD1.n39 VDD1.n5 0.155672
R377 VDD1.n39 VDD1.n38 0.155672
R378 VDD1.n38 VDD1.n9 0.155672
R379 VDD1.n31 VDD1.n9 0.155672
R380 VDD1.n31 VDD1.n30 0.155672
R381 VDD1.n30 VDD1.n14 0.155672
R382 VDD1.n23 VDD1.n14 0.155672
R383 VDD1.n23 VDD1.n22 0.155672
R384 VDD1.n81 VDD1.n80 0.155672
R385 VDD1.n81 VDD1.n72 0.155672
R386 VDD1.n88 VDD1.n72 0.155672
R387 VDD1.n89 VDD1.n88 0.155672
R388 VDD1.n89 VDD1.n68 0.155672
R389 VDD1.n97 VDD1.n68 0.155672
R390 VDD1.n98 VDD1.n97 0.155672
R391 VDD1.n98 VDD1.n64 0.155672
R392 VDD1.n106 VDD1.n64 0.155672
R393 VDD1.n107 VDD1.n106 0.155672
R394 VDD1.n107 VDD1.n60 0.155672
R395 VDD1.n114 VDD1.n60 0.155672
R396 VTAIL.n240 VTAIL.n188 756.745
R397 VTAIL.n54 VTAIL.n2 756.745
R398 VTAIL.n182 VTAIL.n130 756.745
R399 VTAIL.n120 VTAIL.n68 756.745
R400 VTAIL.n207 VTAIL.n206 585
R401 VTAIL.n204 VTAIL.n203 585
R402 VTAIL.n213 VTAIL.n212 585
R403 VTAIL.n215 VTAIL.n214 585
R404 VTAIL.n200 VTAIL.n199 585
R405 VTAIL.n221 VTAIL.n220 585
R406 VTAIL.n224 VTAIL.n223 585
R407 VTAIL.n222 VTAIL.n196 585
R408 VTAIL.n229 VTAIL.n195 585
R409 VTAIL.n231 VTAIL.n230 585
R410 VTAIL.n233 VTAIL.n232 585
R411 VTAIL.n192 VTAIL.n191 585
R412 VTAIL.n239 VTAIL.n238 585
R413 VTAIL.n241 VTAIL.n240 585
R414 VTAIL.n21 VTAIL.n20 585
R415 VTAIL.n18 VTAIL.n17 585
R416 VTAIL.n27 VTAIL.n26 585
R417 VTAIL.n29 VTAIL.n28 585
R418 VTAIL.n14 VTAIL.n13 585
R419 VTAIL.n35 VTAIL.n34 585
R420 VTAIL.n38 VTAIL.n37 585
R421 VTAIL.n36 VTAIL.n10 585
R422 VTAIL.n43 VTAIL.n9 585
R423 VTAIL.n45 VTAIL.n44 585
R424 VTAIL.n47 VTAIL.n46 585
R425 VTAIL.n6 VTAIL.n5 585
R426 VTAIL.n53 VTAIL.n52 585
R427 VTAIL.n55 VTAIL.n54 585
R428 VTAIL.n183 VTAIL.n182 585
R429 VTAIL.n181 VTAIL.n180 585
R430 VTAIL.n134 VTAIL.n133 585
R431 VTAIL.n175 VTAIL.n174 585
R432 VTAIL.n173 VTAIL.n172 585
R433 VTAIL.n171 VTAIL.n137 585
R434 VTAIL.n141 VTAIL.n138 585
R435 VTAIL.n166 VTAIL.n165 585
R436 VTAIL.n164 VTAIL.n163 585
R437 VTAIL.n143 VTAIL.n142 585
R438 VTAIL.n158 VTAIL.n157 585
R439 VTAIL.n156 VTAIL.n155 585
R440 VTAIL.n147 VTAIL.n146 585
R441 VTAIL.n150 VTAIL.n149 585
R442 VTAIL.n121 VTAIL.n120 585
R443 VTAIL.n119 VTAIL.n118 585
R444 VTAIL.n72 VTAIL.n71 585
R445 VTAIL.n113 VTAIL.n112 585
R446 VTAIL.n111 VTAIL.n110 585
R447 VTAIL.n109 VTAIL.n75 585
R448 VTAIL.n79 VTAIL.n76 585
R449 VTAIL.n104 VTAIL.n103 585
R450 VTAIL.n102 VTAIL.n101 585
R451 VTAIL.n81 VTAIL.n80 585
R452 VTAIL.n96 VTAIL.n95 585
R453 VTAIL.n94 VTAIL.n93 585
R454 VTAIL.n85 VTAIL.n84 585
R455 VTAIL.n88 VTAIL.n87 585
R456 VTAIL.t10 VTAIL.n148 329.038
R457 VTAIL.t0 VTAIL.n86 329.038
R458 VTAIL.t4 VTAIL.n205 329.038
R459 VTAIL.t13 VTAIL.n19 329.038
R460 VTAIL.n206 VTAIL.n203 171.744
R461 VTAIL.n213 VTAIL.n203 171.744
R462 VTAIL.n214 VTAIL.n213 171.744
R463 VTAIL.n214 VTAIL.n199 171.744
R464 VTAIL.n221 VTAIL.n199 171.744
R465 VTAIL.n223 VTAIL.n221 171.744
R466 VTAIL.n223 VTAIL.n222 171.744
R467 VTAIL.n222 VTAIL.n195 171.744
R468 VTAIL.n231 VTAIL.n195 171.744
R469 VTAIL.n232 VTAIL.n231 171.744
R470 VTAIL.n232 VTAIL.n191 171.744
R471 VTAIL.n239 VTAIL.n191 171.744
R472 VTAIL.n240 VTAIL.n239 171.744
R473 VTAIL.n20 VTAIL.n17 171.744
R474 VTAIL.n27 VTAIL.n17 171.744
R475 VTAIL.n28 VTAIL.n27 171.744
R476 VTAIL.n28 VTAIL.n13 171.744
R477 VTAIL.n35 VTAIL.n13 171.744
R478 VTAIL.n37 VTAIL.n35 171.744
R479 VTAIL.n37 VTAIL.n36 171.744
R480 VTAIL.n36 VTAIL.n9 171.744
R481 VTAIL.n45 VTAIL.n9 171.744
R482 VTAIL.n46 VTAIL.n45 171.744
R483 VTAIL.n46 VTAIL.n5 171.744
R484 VTAIL.n53 VTAIL.n5 171.744
R485 VTAIL.n54 VTAIL.n53 171.744
R486 VTAIL.n182 VTAIL.n181 171.744
R487 VTAIL.n181 VTAIL.n133 171.744
R488 VTAIL.n174 VTAIL.n133 171.744
R489 VTAIL.n174 VTAIL.n173 171.744
R490 VTAIL.n173 VTAIL.n137 171.744
R491 VTAIL.n141 VTAIL.n137 171.744
R492 VTAIL.n165 VTAIL.n141 171.744
R493 VTAIL.n165 VTAIL.n164 171.744
R494 VTAIL.n164 VTAIL.n142 171.744
R495 VTAIL.n157 VTAIL.n142 171.744
R496 VTAIL.n157 VTAIL.n156 171.744
R497 VTAIL.n156 VTAIL.n146 171.744
R498 VTAIL.n149 VTAIL.n146 171.744
R499 VTAIL.n120 VTAIL.n119 171.744
R500 VTAIL.n119 VTAIL.n71 171.744
R501 VTAIL.n112 VTAIL.n71 171.744
R502 VTAIL.n112 VTAIL.n111 171.744
R503 VTAIL.n111 VTAIL.n75 171.744
R504 VTAIL.n79 VTAIL.n75 171.744
R505 VTAIL.n103 VTAIL.n79 171.744
R506 VTAIL.n103 VTAIL.n102 171.744
R507 VTAIL.n102 VTAIL.n80 171.744
R508 VTAIL.n95 VTAIL.n80 171.744
R509 VTAIL.n95 VTAIL.n94 171.744
R510 VTAIL.n94 VTAIL.n84 171.744
R511 VTAIL.n87 VTAIL.n84 171.744
R512 VTAIL.n206 VTAIL.t4 85.8723
R513 VTAIL.n20 VTAIL.t13 85.8723
R514 VTAIL.n149 VTAIL.t10 85.8723
R515 VTAIL.n87 VTAIL.t0 85.8723
R516 VTAIL.n129 VTAIL.n128 61.5146
R517 VTAIL.n127 VTAIL.n126 61.5146
R518 VTAIL.n67 VTAIL.n66 61.5146
R519 VTAIL.n65 VTAIL.n64 61.5146
R520 VTAIL.n247 VTAIL.n246 61.5145
R521 VTAIL.n1 VTAIL.n0 61.5145
R522 VTAIL.n61 VTAIL.n60 61.5145
R523 VTAIL.n63 VTAIL.n62 61.5145
R524 VTAIL.n245 VTAIL.n244 34.5126
R525 VTAIL.n59 VTAIL.n58 34.5126
R526 VTAIL.n187 VTAIL.n186 34.5126
R527 VTAIL.n125 VTAIL.n124 34.5126
R528 VTAIL.n65 VTAIL.n63 29.0221
R529 VTAIL.n245 VTAIL.n187 25.3496
R530 VTAIL.n230 VTAIL.n229 13.1884
R531 VTAIL.n44 VTAIL.n43 13.1884
R532 VTAIL.n172 VTAIL.n171 13.1884
R533 VTAIL.n110 VTAIL.n109 13.1884
R534 VTAIL.n228 VTAIL.n196 12.8005
R535 VTAIL.n233 VTAIL.n194 12.8005
R536 VTAIL.n42 VTAIL.n10 12.8005
R537 VTAIL.n47 VTAIL.n8 12.8005
R538 VTAIL.n175 VTAIL.n136 12.8005
R539 VTAIL.n170 VTAIL.n138 12.8005
R540 VTAIL.n113 VTAIL.n74 12.8005
R541 VTAIL.n108 VTAIL.n76 12.8005
R542 VTAIL.n225 VTAIL.n224 12.0247
R543 VTAIL.n234 VTAIL.n192 12.0247
R544 VTAIL.n39 VTAIL.n38 12.0247
R545 VTAIL.n48 VTAIL.n6 12.0247
R546 VTAIL.n176 VTAIL.n134 12.0247
R547 VTAIL.n167 VTAIL.n166 12.0247
R548 VTAIL.n114 VTAIL.n72 12.0247
R549 VTAIL.n105 VTAIL.n104 12.0247
R550 VTAIL.n220 VTAIL.n198 11.249
R551 VTAIL.n238 VTAIL.n237 11.249
R552 VTAIL.n34 VTAIL.n12 11.249
R553 VTAIL.n52 VTAIL.n51 11.249
R554 VTAIL.n180 VTAIL.n179 11.249
R555 VTAIL.n163 VTAIL.n140 11.249
R556 VTAIL.n118 VTAIL.n117 11.249
R557 VTAIL.n101 VTAIL.n78 11.249
R558 VTAIL.n207 VTAIL.n205 10.7239
R559 VTAIL.n21 VTAIL.n19 10.7239
R560 VTAIL.n150 VTAIL.n148 10.7239
R561 VTAIL.n88 VTAIL.n86 10.7239
R562 VTAIL.n219 VTAIL.n200 10.4732
R563 VTAIL.n241 VTAIL.n190 10.4732
R564 VTAIL.n33 VTAIL.n14 10.4732
R565 VTAIL.n55 VTAIL.n4 10.4732
R566 VTAIL.n183 VTAIL.n132 10.4732
R567 VTAIL.n162 VTAIL.n143 10.4732
R568 VTAIL.n121 VTAIL.n70 10.4732
R569 VTAIL.n100 VTAIL.n81 10.4732
R570 VTAIL.n216 VTAIL.n215 9.69747
R571 VTAIL.n242 VTAIL.n188 9.69747
R572 VTAIL.n30 VTAIL.n29 9.69747
R573 VTAIL.n56 VTAIL.n2 9.69747
R574 VTAIL.n184 VTAIL.n130 9.69747
R575 VTAIL.n159 VTAIL.n158 9.69747
R576 VTAIL.n122 VTAIL.n68 9.69747
R577 VTAIL.n97 VTAIL.n96 9.69747
R578 VTAIL.n244 VTAIL.n243 9.45567
R579 VTAIL.n58 VTAIL.n57 9.45567
R580 VTAIL.n186 VTAIL.n185 9.45567
R581 VTAIL.n124 VTAIL.n123 9.45567
R582 VTAIL.n243 VTAIL.n242 9.3005
R583 VTAIL.n190 VTAIL.n189 9.3005
R584 VTAIL.n237 VTAIL.n236 9.3005
R585 VTAIL.n235 VTAIL.n234 9.3005
R586 VTAIL.n194 VTAIL.n193 9.3005
R587 VTAIL.n209 VTAIL.n208 9.3005
R588 VTAIL.n211 VTAIL.n210 9.3005
R589 VTAIL.n202 VTAIL.n201 9.3005
R590 VTAIL.n217 VTAIL.n216 9.3005
R591 VTAIL.n219 VTAIL.n218 9.3005
R592 VTAIL.n198 VTAIL.n197 9.3005
R593 VTAIL.n226 VTAIL.n225 9.3005
R594 VTAIL.n228 VTAIL.n227 9.3005
R595 VTAIL.n57 VTAIL.n56 9.3005
R596 VTAIL.n4 VTAIL.n3 9.3005
R597 VTAIL.n51 VTAIL.n50 9.3005
R598 VTAIL.n49 VTAIL.n48 9.3005
R599 VTAIL.n8 VTAIL.n7 9.3005
R600 VTAIL.n23 VTAIL.n22 9.3005
R601 VTAIL.n25 VTAIL.n24 9.3005
R602 VTAIL.n16 VTAIL.n15 9.3005
R603 VTAIL.n31 VTAIL.n30 9.3005
R604 VTAIL.n33 VTAIL.n32 9.3005
R605 VTAIL.n12 VTAIL.n11 9.3005
R606 VTAIL.n40 VTAIL.n39 9.3005
R607 VTAIL.n42 VTAIL.n41 9.3005
R608 VTAIL.n152 VTAIL.n151 9.3005
R609 VTAIL.n154 VTAIL.n153 9.3005
R610 VTAIL.n145 VTAIL.n144 9.3005
R611 VTAIL.n160 VTAIL.n159 9.3005
R612 VTAIL.n162 VTAIL.n161 9.3005
R613 VTAIL.n140 VTAIL.n139 9.3005
R614 VTAIL.n168 VTAIL.n167 9.3005
R615 VTAIL.n170 VTAIL.n169 9.3005
R616 VTAIL.n185 VTAIL.n184 9.3005
R617 VTAIL.n132 VTAIL.n131 9.3005
R618 VTAIL.n179 VTAIL.n178 9.3005
R619 VTAIL.n177 VTAIL.n176 9.3005
R620 VTAIL.n136 VTAIL.n135 9.3005
R621 VTAIL.n90 VTAIL.n89 9.3005
R622 VTAIL.n92 VTAIL.n91 9.3005
R623 VTAIL.n83 VTAIL.n82 9.3005
R624 VTAIL.n98 VTAIL.n97 9.3005
R625 VTAIL.n100 VTAIL.n99 9.3005
R626 VTAIL.n78 VTAIL.n77 9.3005
R627 VTAIL.n106 VTAIL.n105 9.3005
R628 VTAIL.n108 VTAIL.n107 9.3005
R629 VTAIL.n123 VTAIL.n122 9.3005
R630 VTAIL.n70 VTAIL.n69 9.3005
R631 VTAIL.n117 VTAIL.n116 9.3005
R632 VTAIL.n115 VTAIL.n114 9.3005
R633 VTAIL.n74 VTAIL.n73 9.3005
R634 VTAIL.n212 VTAIL.n202 8.92171
R635 VTAIL.n26 VTAIL.n16 8.92171
R636 VTAIL.n155 VTAIL.n145 8.92171
R637 VTAIL.n93 VTAIL.n83 8.92171
R638 VTAIL.n211 VTAIL.n204 8.14595
R639 VTAIL.n25 VTAIL.n18 8.14595
R640 VTAIL.n154 VTAIL.n147 8.14595
R641 VTAIL.n92 VTAIL.n85 8.14595
R642 VTAIL.n208 VTAIL.n207 7.3702
R643 VTAIL.n22 VTAIL.n21 7.3702
R644 VTAIL.n151 VTAIL.n150 7.3702
R645 VTAIL.n89 VTAIL.n88 7.3702
R646 VTAIL.n208 VTAIL.n204 5.81868
R647 VTAIL.n22 VTAIL.n18 5.81868
R648 VTAIL.n151 VTAIL.n147 5.81868
R649 VTAIL.n89 VTAIL.n85 5.81868
R650 VTAIL.n212 VTAIL.n211 5.04292
R651 VTAIL.n26 VTAIL.n25 5.04292
R652 VTAIL.n155 VTAIL.n154 5.04292
R653 VTAIL.n93 VTAIL.n92 5.04292
R654 VTAIL.n215 VTAIL.n202 4.26717
R655 VTAIL.n244 VTAIL.n188 4.26717
R656 VTAIL.n29 VTAIL.n16 4.26717
R657 VTAIL.n58 VTAIL.n2 4.26717
R658 VTAIL.n186 VTAIL.n130 4.26717
R659 VTAIL.n158 VTAIL.n145 4.26717
R660 VTAIL.n124 VTAIL.n68 4.26717
R661 VTAIL.n96 VTAIL.n83 4.26717
R662 VTAIL.n67 VTAIL.n65 3.67291
R663 VTAIL.n125 VTAIL.n67 3.67291
R664 VTAIL.n129 VTAIL.n127 3.67291
R665 VTAIL.n187 VTAIL.n129 3.67291
R666 VTAIL.n63 VTAIL.n61 3.67291
R667 VTAIL.n61 VTAIL.n59 3.67291
R668 VTAIL.n247 VTAIL.n245 3.67291
R669 VTAIL.n216 VTAIL.n200 3.49141
R670 VTAIL.n242 VTAIL.n241 3.49141
R671 VTAIL.n30 VTAIL.n14 3.49141
R672 VTAIL.n56 VTAIL.n55 3.49141
R673 VTAIL.n184 VTAIL.n183 3.49141
R674 VTAIL.n159 VTAIL.n143 3.49141
R675 VTAIL.n122 VTAIL.n121 3.49141
R676 VTAIL.n97 VTAIL.n81 3.49141
R677 VTAIL.n246 VTAIL.t18 3.01022
R678 VTAIL.n246 VTAIL.t7 3.01022
R679 VTAIL.n0 VTAIL.t19 3.01022
R680 VTAIL.n0 VTAIL.t1 3.01022
R681 VTAIL.n60 VTAIL.t12 3.01022
R682 VTAIL.n60 VTAIL.t8 3.01022
R683 VTAIL.n62 VTAIL.t15 3.01022
R684 VTAIL.n62 VTAIL.t9 3.01022
R685 VTAIL.n128 VTAIL.t11 3.01022
R686 VTAIL.n128 VTAIL.t16 3.01022
R687 VTAIL.n126 VTAIL.t14 3.01022
R688 VTAIL.n126 VTAIL.t17 3.01022
R689 VTAIL.n66 VTAIL.t6 3.01022
R690 VTAIL.n66 VTAIL.t2 3.01022
R691 VTAIL.n64 VTAIL.t3 3.01022
R692 VTAIL.n64 VTAIL.t5 3.01022
R693 VTAIL VTAIL.n1 2.813
R694 VTAIL.n220 VTAIL.n219 2.71565
R695 VTAIL.n238 VTAIL.n190 2.71565
R696 VTAIL.n34 VTAIL.n33 2.71565
R697 VTAIL.n52 VTAIL.n4 2.71565
R698 VTAIL.n180 VTAIL.n132 2.71565
R699 VTAIL.n163 VTAIL.n162 2.71565
R700 VTAIL.n118 VTAIL.n70 2.71565
R701 VTAIL.n101 VTAIL.n100 2.71565
R702 VTAIL.n209 VTAIL.n205 2.41282
R703 VTAIL.n23 VTAIL.n19 2.41282
R704 VTAIL.n152 VTAIL.n148 2.41282
R705 VTAIL.n90 VTAIL.n86 2.41282
R706 VTAIL.n127 VTAIL.n125 2.30653
R707 VTAIL.n59 VTAIL.n1 2.30653
R708 VTAIL.n224 VTAIL.n198 1.93989
R709 VTAIL.n237 VTAIL.n192 1.93989
R710 VTAIL.n38 VTAIL.n12 1.93989
R711 VTAIL.n51 VTAIL.n6 1.93989
R712 VTAIL.n179 VTAIL.n134 1.93989
R713 VTAIL.n166 VTAIL.n140 1.93989
R714 VTAIL.n117 VTAIL.n72 1.93989
R715 VTAIL.n104 VTAIL.n78 1.93989
R716 VTAIL.n225 VTAIL.n196 1.16414
R717 VTAIL.n234 VTAIL.n233 1.16414
R718 VTAIL.n39 VTAIL.n10 1.16414
R719 VTAIL.n48 VTAIL.n47 1.16414
R720 VTAIL.n176 VTAIL.n175 1.16414
R721 VTAIL.n167 VTAIL.n138 1.16414
R722 VTAIL.n114 VTAIL.n113 1.16414
R723 VTAIL.n105 VTAIL.n76 1.16414
R724 VTAIL VTAIL.n247 0.860414
R725 VTAIL.n229 VTAIL.n228 0.388379
R726 VTAIL.n230 VTAIL.n194 0.388379
R727 VTAIL.n43 VTAIL.n42 0.388379
R728 VTAIL.n44 VTAIL.n8 0.388379
R729 VTAIL.n172 VTAIL.n136 0.388379
R730 VTAIL.n171 VTAIL.n170 0.388379
R731 VTAIL.n110 VTAIL.n74 0.388379
R732 VTAIL.n109 VTAIL.n108 0.388379
R733 VTAIL.n210 VTAIL.n209 0.155672
R734 VTAIL.n210 VTAIL.n201 0.155672
R735 VTAIL.n217 VTAIL.n201 0.155672
R736 VTAIL.n218 VTAIL.n217 0.155672
R737 VTAIL.n218 VTAIL.n197 0.155672
R738 VTAIL.n226 VTAIL.n197 0.155672
R739 VTAIL.n227 VTAIL.n226 0.155672
R740 VTAIL.n227 VTAIL.n193 0.155672
R741 VTAIL.n235 VTAIL.n193 0.155672
R742 VTAIL.n236 VTAIL.n235 0.155672
R743 VTAIL.n236 VTAIL.n189 0.155672
R744 VTAIL.n243 VTAIL.n189 0.155672
R745 VTAIL.n24 VTAIL.n23 0.155672
R746 VTAIL.n24 VTAIL.n15 0.155672
R747 VTAIL.n31 VTAIL.n15 0.155672
R748 VTAIL.n32 VTAIL.n31 0.155672
R749 VTAIL.n32 VTAIL.n11 0.155672
R750 VTAIL.n40 VTAIL.n11 0.155672
R751 VTAIL.n41 VTAIL.n40 0.155672
R752 VTAIL.n41 VTAIL.n7 0.155672
R753 VTAIL.n49 VTAIL.n7 0.155672
R754 VTAIL.n50 VTAIL.n49 0.155672
R755 VTAIL.n50 VTAIL.n3 0.155672
R756 VTAIL.n57 VTAIL.n3 0.155672
R757 VTAIL.n185 VTAIL.n131 0.155672
R758 VTAIL.n178 VTAIL.n131 0.155672
R759 VTAIL.n178 VTAIL.n177 0.155672
R760 VTAIL.n177 VTAIL.n135 0.155672
R761 VTAIL.n169 VTAIL.n135 0.155672
R762 VTAIL.n169 VTAIL.n168 0.155672
R763 VTAIL.n168 VTAIL.n139 0.155672
R764 VTAIL.n161 VTAIL.n139 0.155672
R765 VTAIL.n161 VTAIL.n160 0.155672
R766 VTAIL.n160 VTAIL.n144 0.155672
R767 VTAIL.n153 VTAIL.n144 0.155672
R768 VTAIL.n153 VTAIL.n152 0.155672
R769 VTAIL.n123 VTAIL.n69 0.155672
R770 VTAIL.n116 VTAIL.n69 0.155672
R771 VTAIL.n116 VTAIL.n115 0.155672
R772 VTAIL.n115 VTAIL.n73 0.155672
R773 VTAIL.n107 VTAIL.n73 0.155672
R774 VTAIL.n107 VTAIL.n106 0.155672
R775 VTAIL.n106 VTAIL.n77 0.155672
R776 VTAIL.n99 VTAIL.n77 0.155672
R777 VTAIL.n99 VTAIL.n98 0.155672
R778 VTAIL.n98 VTAIL.n82 0.155672
R779 VTAIL.n91 VTAIL.n82 0.155672
R780 VTAIL.n91 VTAIL.n90 0.155672
R781 VN.n112 VN.n111 161.3
R782 VN.n110 VN.n58 161.3
R783 VN.n109 VN.n108 161.3
R784 VN.n107 VN.n59 161.3
R785 VN.n106 VN.n105 161.3
R786 VN.n104 VN.n60 161.3
R787 VN.n103 VN.n102 161.3
R788 VN.n101 VN.n61 161.3
R789 VN.n100 VN.n99 161.3
R790 VN.n97 VN.n62 161.3
R791 VN.n96 VN.n95 161.3
R792 VN.n94 VN.n63 161.3
R793 VN.n93 VN.n92 161.3
R794 VN.n91 VN.n64 161.3
R795 VN.n90 VN.n89 161.3
R796 VN.n88 VN.n65 161.3
R797 VN.n87 VN.n86 161.3
R798 VN.n85 VN.n66 161.3
R799 VN.n84 VN.n83 161.3
R800 VN.n82 VN.n67 161.3
R801 VN.n81 VN.n80 161.3
R802 VN.n79 VN.n68 161.3
R803 VN.n78 VN.n77 161.3
R804 VN.n76 VN.n69 161.3
R805 VN.n75 VN.n74 161.3
R806 VN.n73 VN.n70 161.3
R807 VN.n55 VN.n54 161.3
R808 VN.n53 VN.n1 161.3
R809 VN.n52 VN.n51 161.3
R810 VN.n50 VN.n2 161.3
R811 VN.n49 VN.n48 161.3
R812 VN.n47 VN.n3 161.3
R813 VN.n46 VN.n45 161.3
R814 VN.n44 VN.n4 161.3
R815 VN.n43 VN.n42 161.3
R816 VN.n40 VN.n5 161.3
R817 VN.n39 VN.n38 161.3
R818 VN.n37 VN.n6 161.3
R819 VN.n36 VN.n35 161.3
R820 VN.n34 VN.n7 161.3
R821 VN.n33 VN.n32 161.3
R822 VN.n31 VN.n8 161.3
R823 VN.n30 VN.n29 161.3
R824 VN.n28 VN.n9 161.3
R825 VN.n27 VN.n26 161.3
R826 VN.n25 VN.n10 161.3
R827 VN.n24 VN.n23 161.3
R828 VN.n22 VN.n11 161.3
R829 VN.n21 VN.n20 161.3
R830 VN.n19 VN.n12 161.3
R831 VN.n18 VN.n17 161.3
R832 VN.n16 VN.n13 161.3
R833 VN.n71 VN.t4 98.4421
R834 VN.n14 VN.t8 98.4421
R835 VN.n56 VN.n0 88.9173
R836 VN.n113 VN.n57 88.9173
R837 VN.n28 VN.t6 66.2295
R838 VN.n15 VN.t2 66.2295
R839 VN.n41 VN.t9 66.2295
R840 VN.n0 VN.t7 66.2295
R841 VN.n85 VN.t1 66.2295
R842 VN.n72 VN.t0 66.2295
R843 VN.n98 VN.t5 66.2295
R844 VN.n57 VN.t3 66.2295
R845 VN.n15 VN.n14 62.2666
R846 VN.n72 VN.n71 62.2666
R847 VN VN.n113 59.657
R848 VN.n22 VN.n21 53.0692
R849 VN.n35 VN.n34 53.0692
R850 VN.n79 VN.n78 53.0692
R851 VN.n92 VN.n91 53.0692
R852 VN.n48 VN.n47 51.1217
R853 VN.n105 VN.n104 51.1217
R854 VN.n48 VN.n2 29.6995
R855 VN.n105 VN.n59 29.6995
R856 VN.n23 VN.n22 27.752
R857 VN.n34 VN.n33 27.752
R858 VN.n80 VN.n79 27.752
R859 VN.n91 VN.n90 27.752
R860 VN.n17 VN.n16 24.3439
R861 VN.n17 VN.n12 24.3439
R862 VN.n21 VN.n12 24.3439
R863 VN.n23 VN.n10 24.3439
R864 VN.n27 VN.n10 24.3439
R865 VN.n28 VN.n27 24.3439
R866 VN.n29 VN.n28 24.3439
R867 VN.n29 VN.n8 24.3439
R868 VN.n33 VN.n8 24.3439
R869 VN.n35 VN.n6 24.3439
R870 VN.n39 VN.n6 24.3439
R871 VN.n40 VN.n39 24.3439
R872 VN.n42 VN.n4 24.3439
R873 VN.n46 VN.n4 24.3439
R874 VN.n47 VN.n46 24.3439
R875 VN.n52 VN.n2 24.3439
R876 VN.n53 VN.n52 24.3439
R877 VN.n54 VN.n53 24.3439
R878 VN.n78 VN.n69 24.3439
R879 VN.n74 VN.n69 24.3439
R880 VN.n74 VN.n73 24.3439
R881 VN.n90 VN.n65 24.3439
R882 VN.n86 VN.n65 24.3439
R883 VN.n86 VN.n85 24.3439
R884 VN.n85 VN.n84 24.3439
R885 VN.n84 VN.n67 24.3439
R886 VN.n80 VN.n67 24.3439
R887 VN.n104 VN.n103 24.3439
R888 VN.n103 VN.n61 24.3439
R889 VN.n99 VN.n61 24.3439
R890 VN.n97 VN.n96 24.3439
R891 VN.n96 VN.n63 24.3439
R892 VN.n92 VN.n63 24.3439
R893 VN.n111 VN.n110 24.3439
R894 VN.n110 VN.n109 24.3439
R895 VN.n109 VN.n59 24.3439
R896 VN.n16 VN.n15 12.6591
R897 VN.n41 VN.n40 12.6591
R898 VN.n73 VN.n72 12.6591
R899 VN.n98 VN.n97 12.6591
R900 VN.n42 VN.n41 11.6853
R901 VN.n99 VN.n98 11.6853
R902 VN.n71 VN.n70 2.52182
R903 VN.n14 VN.n13 2.52182
R904 VN.n54 VN.n0 0.974237
R905 VN.n111 VN.n57 0.974237
R906 VN.n113 VN.n112 0.355081
R907 VN.n56 VN.n55 0.355081
R908 VN VN.n56 0.26685
R909 VN.n112 VN.n58 0.189894
R910 VN.n108 VN.n58 0.189894
R911 VN.n108 VN.n107 0.189894
R912 VN.n107 VN.n106 0.189894
R913 VN.n106 VN.n60 0.189894
R914 VN.n102 VN.n60 0.189894
R915 VN.n102 VN.n101 0.189894
R916 VN.n101 VN.n100 0.189894
R917 VN.n100 VN.n62 0.189894
R918 VN.n95 VN.n62 0.189894
R919 VN.n95 VN.n94 0.189894
R920 VN.n94 VN.n93 0.189894
R921 VN.n93 VN.n64 0.189894
R922 VN.n89 VN.n64 0.189894
R923 VN.n89 VN.n88 0.189894
R924 VN.n88 VN.n87 0.189894
R925 VN.n87 VN.n66 0.189894
R926 VN.n83 VN.n66 0.189894
R927 VN.n83 VN.n82 0.189894
R928 VN.n82 VN.n81 0.189894
R929 VN.n81 VN.n68 0.189894
R930 VN.n77 VN.n68 0.189894
R931 VN.n77 VN.n76 0.189894
R932 VN.n76 VN.n75 0.189894
R933 VN.n75 VN.n70 0.189894
R934 VN.n18 VN.n13 0.189894
R935 VN.n19 VN.n18 0.189894
R936 VN.n20 VN.n19 0.189894
R937 VN.n20 VN.n11 0.189894
R938 VN.n24 VN.n11 0.189894
R939 VN.n25 VN.n24 0.189894
R940 VN.n26 VN.n25 0.189894
R941 VN.n26 VN.n9 0.189894
R942 VN.n30 VN.n9 0.189894
R943 VN.n31 VN.n30 0.189894
R944 VN.n32 VN.n31 0.189894
R945 VN.n32 VN.n7 0.189894
R946 VN.n36 VN.n7 0.189894
R947 VN.n37 VN.n36 0.189894
R948 VN.n38 VN.n37 0.189894
R949 VN.n38 VN.n5 0.189894
R950 VN.n43 VN.n5 0.189894
R951 VN.n44 VN.n43 0.189894
R952 VN.n45 VN.n44 0.189894
R953 VN.n45 VN.n3 0.189894
R954 VN.n49 VN.n3 0.189894
R955 VN.n50 VN.n49 0.189894
R956 VN.n51 VN.n50 0.189894
R957 VN.n51 VN.n1 0.189894
R958 VN.n55 VN.n1 0.189894
R959 VDD2.n113 VDD2.n61 756.745
R960 VDD2.n52 VDD2.n0 756.745
R961 VDD2.n114 VDD2.n113 585
R962 VDD2.n112 VDD2.n111 585
R963 VDD2.n65 VDD2.n64 585
R964 VDD2.n106 VDD2.n105 585
R965 VDD2.n104 VDD2.n103 585
R966 VDD2.n102 VDD2.n68 585
R967 VDD2.n72 VDD2.n69 585
R968 VDD2.n97 VDD2.n96 585
R969 VDD2.n95 VDD2.n94 585
R970 VDD2.n74 VDD2.n73 585
R971 VDD2.n89 VDD2.n88 585
R972 VDD2.n87 VDD2.n86 585
R973 VDD2.n78 VDD2.n77 585
R974 VDD2.n81 VDD2.n80 585
R975 VDD2.n19 VDD2.n18 585
R976 VDD2.n16 VDD2.n15 585
R977 VDD2.n25 VDD2.n24 585
R978 VDD2.n27 VDD2.n26 585
R979 VDD2.n12 VDD2.n11 585
R980 VDD2.n33 VDD2.n32 585
R981 VDD2.n36 VDD2.n35 585
R982 VDD2.n34 VDD2.n8 585
R983 VDD2.n41 VDD2.n7 585
R984 VDD2.n43 VDD2.n42 585
R985 VDD2.n45 VDD2.n44 585
R986 VDD2.n4 VDD2.n3 585
R987 VDD2.n51 VDD2.n50 585
R988 VDD2.n53 VDD2.n52 585
R989 VDD2.t6 VDD2.n79 329.038
R990 VDD2.t1 VDD2.n17 329.038
R991 VDD2.n113 VDD2.n112 171.744
R992 VDD2.n112 VDD2.n64 171.744
R993 VDD2.n105 VDD2.n64 171.744
R994 VDD2.n105 VDD2.n104 171.744
R995 VDD2.n104 VDD2.n68 171.744
R996 VDD2.n72 VDD2.n68 171.744
R997 VDD2.n96 VDD2.n72 171.744
R998 VDD2.n96 VDD2.n95 171.744
R999 VDD2.n95 VDD2.n73 171.744
R1000 VDD2.n88 VDD2.n73 171.744
R1001 VDD2.n88 VDD2.n87 171.744
R1002 VDD2.n87 VDD2.n77 171.744
R1003 VDD2.n80 VDD2.n77 171.744
R1004 VDD2.n18 VDD2.n15 171.744
R1005 VDD2.n25 VDD2.n15 171.744
R1006 VDD2.n26 VDD2.n25 171.744
R1007 VDD2.n26 VDD2.n11 171.744
R1008 VDD2.n33 VDD2.n11 171.744
R1009 VDD2.n35 VDD2.n33 171.744
R1010 VDD2.n35 VDD2.n34 171.744
R1011 VDD2.n34 VDD2.n7 171.744
R1012 VDD2.n43 VDD2.n7 171.744
R1013 VDD2.n44 VDD2.n43 171.744
R1014 VDD2.n44 VDD2.n3 171.744
R1015 VDD2.n51 VDD2.n3 171.744
R1016 VDD2.n52 VDD2.n51 171.744
R1017 VDD2.n80 VDD2.t6 85.8723
R1018 VDD2.n18 VDD2.t1 85.8723
R1019 VDD2.n60 VDD2.n59 80.8922
R1020 VDD2 VDD2.n121 80.8894
R1021 VDD2.n120 VDD2.n119 78.1934
R1022 VDD2.n58 VDD2.n57 78.1932
R1023 VDD2.n58 VDD2.n56 54.8638
R1024 VDD2.n118 VDD2.n117 51.1914
R1025 VDD2.n118 VDD2.n60 50.4696
R1026 VDD2.n103 VDD2.n102 13.1884
R1027 VDD2.n42 VDD2.n41 13.1884
R1028 VDD2.n106 VDD2.n67 12.8005
R1029 VDD2.n101 VDD2.n69 12.8005
R1030 VDD2.n40 VDD2.n8 12.8005
R1031 VDD2.n45 VDD2.n6 12.8005
R1032 VDD2.n107 VDD2.n65 12.0247
R1033 VDD2.n98 VDD2.n97 12.0247
R1034 VDD2.n37 VDD2.n36 12.0247
R1035 VDD2.n46 VDD2.n4 12.0247
R1036 VDD2.n111 VDD2.n110 11.249
R1037 VDD2.n94 VDD2.n71 11.249
R1038 VDD2.n32 VDD2.n10 11.249
R1039 VDD2.n50 VDD2.n49 11.249
R1040 VDD2.n81 VDD2.n79 10.7239
R1041 VDD2.n19 VDD2.n17 10.7239
R1042 VDD2.n114 VDD2.n63 10.4732
R1043 VDD2.n93 VDD2.n74 10.4732
R1044 VDD2.n31 VDD2.n12 10.4732
R1045 VDD2.n53 VDD2.n2 10.4732
R1046 VDD2.n115 VDD2.n61 9.69747
R1047 VDD2.n90 VDD2.n89 9.69747
R1048 VDD2.n28 VDD2.n27 9.69747
R1049 VDD2.n54 VDD2.n0 9.69747
R1050 VDD2.n117 VDD2.n116 9.45567
R1051 VDD2.n56 VDD2.n55 9.45567
R1052 VDD2.n83 VDD2.n82 9.3005
R1053 VDD2.n85 VDD2.n84 9.3005
R1054 VDD2.n76 VDD2.n75 9.3005
R1055 VDD2.n91 VDD2.n90 9.3005
R1056 VDD2.n93 VDD2.n92 9.3005
R1057 VDD2.n71 VDD2.n70 9.3005
R1058 VDD2.n99 VDD2.n98 9.3005
R1059 VDD2.n101 VDD2.n100 9.3005
R1060 VDD2.n116 VDD2.n115 9.3005
R1061 VDD2.n63 VDD2.n62 9.3005
R1062 VDD2.n110 VDD2.n109 9.3005
R1063 VDD2.n108 VDD2.n107 9.3005
R1064 VDD2.n67 VDD2.n66 9.3005
R1065 VDD2.n55 VDD2.n54 9.3005
R1066 VDD2.n2 VDD2.n1 9.3005
R1067 VDD2.n49 VDD2.n48 9.3005
R1068 VDD2.n47 VDD2.n46 9.3005
R1069 VDD2.n6 VDD2.n5 9.3005
R1070 VDD2.n21 VDD2.n20 9.3005
R1071 VDD2.n23 VDD2.n22 9.3005
R1072 VDD2.n14 VDD2.n13 9.3005
R1073 VDD2.n29 VDD2.n28 9.3005
R1074 VDD2.n31 VDD2.n30 9.3005
R1075 VDD2.n10 VDD2.n9 9.3005
R1076 VDD2.n38 VDD2.n37 9.3005
R1077 VDD2.n40 VDD2.n39 9.3005
R1078 VDD2.n86 VDD2.n76 8.92171
R1079 VDD2.n24 VDD2.n14 8.92171
R1080 VDD2.n85 VDD2.n78 8.14595
R1081 VDD2.n23 VDD2.n16 8.14595
R1082 VDD2.n82 VDD2.n81 7.3702
R1083 VDD2.n20 VDD2.n19 7.3702
R1084 VDD2.n82 VDD2.n78 5.81868
R1085 VDD2.n20 VDD2.n16 5.81868
R1086 VDD2.n86 VDD2.n85 5.04292
R1087 VDD2.n24 VDD2.n23 5.04292
R1088 VDD2.n117 VDD2.n61 4.26717
R1089 VDD2.n89 VDD2.n76 4.26717
R1090 VDD2.n27 VDD2.n14 4.26717
R1091 VDD2.n56 VDD2.n0 4.26717
R1092 VDD2.n120 VDD2.n118 3.67291
R1093 VDD2.n115 VDD2.n114 3.49141
R1094 VDD2.n90 VDD2.n74 3.49141
R1095 VDD2.n28 VDD2.n12 3.49141
R1096 VDD2.n54 VDD2.n53 3.49141
R1097 VDD2.n121 VDD2.t9 3.01022
R1098 VDD2.n121 VDD2.t5 3.01022
R1099 VDD2.n119 VDD2.t4 3.01022
R1100 VDD2.n119 VDD2.t8 3.01022
R1101 VDD2.n59 VDD2.t0 3.01022
R1102 VDD2.n59 VDD2.t2 3.01022
R1103 VDD2.n57 VDD2.t7 3.01022
R1104 VDD2.n57 VDD2.t3 3.01022
R1105 VDD2.n111 VDD2.n63 2.71565
R1106 VDD2.n94 VDD2.n93 2.71565
R1107 VDD2.n32 VDD2.n31 2.71565
R1108 VDD2.n50 VDD2.n2 2.71565
R1109 VDD2.n83 VDD2.n79 2.41282
R1110 VDD2.n21 VDD2.n17 2.41282
R1111 VDD2.n110 VDD2.n65 1.93989
R1112 VDD2.n97 VDD2.n71 1.93989
R1113 VDD2.n36 VDD2.n10 1.93989
R1114 VDD2.n49 VDD2.n4 1.93989
R1115 VDD2.n107 VDD2.n106 1.16414
R1116 VDD2.n98 VDD2.n69 1.16414
R1117 VDD2.n37 VDD2.n8 1.16414
R1118 VDD2.n46 VDD2.n45 1.16414
R1119 VDD2 VDD2.n120 0.976793
R1120 VDD2.n60 VDD2.n58 0.863257
R1121 VDD2.n103 VDD2.n67 0.388379
R1122 VDD2.n102 VDD2.n101 0.388379
R1123 VDD2.n41 VDD2.n40 0.388379
R1124 VDD2.n42 VDD2.n6 0.388379
R1125 VDD2.n116 VDD2.n62 0.155672
R1126 VDD2.n109 VDD2.n62 0.155672
R1127 VDD2.n109 VDD2.n108 0.155672
R1128 VDD2.n108 VDD2.n66 0.155672
R1129 VDD2.n100 VDD2.n66 0.155672
R1130 VDD2.n100 VDD2.n99 0.155672
R1131 VDD2.n99 VDD2.n70 0.155672
R1132 VDD2.n92 VDD2.n70 0.155672
R1133 VDD2.n92 VDD2.n91 0.155672
R1134 VDD2.n91 VDD2.n75 0.155672
R1135 VDD2.n84 VDD2.n75 0.155672
R1136 VDD2.n84 VDD2.n83 0.155672
R1137 VDD2.n22 VDD2.n21 0.155672
R1138 VDD2.n22 VDD2.n13 0.155672
R1139 VDD2.n29 VDD2.n13 0.155672
R1140 VDD2.n30 VDD2.n29 0.155672
R1141 VDD2.n30 VDD2.n9 0.155672
R1142 VDD2.n38 VDD2.n9 0.155672
R1143 VDD2.n39 VDD2.n38 0.155672
R1144 VDD2.n39 VDD2.n5 0.155672
R1145 VDD2.n47 VDD2.n5 0.155672
R1146 VDD2.n48 VDD2.n47 0.155672
R1147 VDD2.n48 VDD2.n1 0.155672
R1148 VDD2.n55 VDD2.n1 0.155672
R1149 B.n517 B.n516 585
R1150 B.n515 B.n176 585
R1151 B.n514 B.n513 585
R1152 B.n512 B.n177 585
R1153 B.n511 B.n510 585
R1154 B.n509 B.n178 585
R1155 B.n508 B.n507 585
R1156 B.n506 B.n179 585
R1157 B.n505 B.n504 585
R1158 B.n503 B.n180 585
R1159 B.n502 B.n501 585
R1160 B.n500 B.n181 585
R1161 B.n499 B.n498 585
R1162 B.n497 B.n182 585
R1163 B.n496 B.n495 585
R1164 B.n494 B.n183 585
R1165 B.n493 B.n492 585
R1166 B.n491 B.n184 585
R1167 B.n490 B.n489 585
R1168 B.n488 B.n185 585
R1169 B.n487 B.n486 585
R1170 B.n485 B.n186 585
R1171 B.n484 B.n483 585
R1172 B.n482 B.n187 585
R1173 B.n481 B.n480 585
R1174 B.n479 B.n188 585
R1175 B.n478 B.n477 585
R1176 B.n476 B.n189 585
R1177 B.n475 B.n474 585
R1178 B.n473 B.n190 585
R1179 B.n472 B.n471 585
R1180 B.n470 B.n191 585
R1181 B.n469 B.n468 585
R1182 B.n467 B.n192 585
R1183 B.n466 B.n465 585
R1184 B.n464 B.n193 585
R1185 B.n463 B.n462 585
R1186 B.n461 B.n194 585
R1187 B.n459 B.n458 585
R1188 B.n457 B.n197 585
R1189 B.n456 B.n455 585
R1190 B.n454 B.n198 585
R1191 B.n453 B.n452 585
R1192 B.n451 B.n199 585
R1193 B.n450 B.n449 585
R1194 B.n448 B.n200 585
R1195 B.n447 B.n446 585
R1196 B.n445 B.n201 585
R1197 B.n444 B.n443 585
R1198 B.n439 B.n202 585
R1199 B.n438 B.n437 585
R1200 B.n436 B.n203 585
R1201 B.n435 B.n434 585
R1202 B.n433 B.n204 585
R1203 B.n432 B.n431 585
R1204 B.n430 B.n205 585
R1205 B.n429 B.n428 585
R1206 B.n427 B.n206 585
R1207 B.n426 B.n425 585
R1208 B.n424 B.n207 585
R1209 B.n423 B.n422 585
R1210 B.n421 B.n208 585
R1211 B.n420 B.n419 585
R1212 B.n418 B.n209 585
R1213 B.n417 B.n416 585
R1214 B.n415 B.n210 585
R1215 B.n414 B.n413 585
R1216 B.n412 B.n211 585
R1217 B.n411 B.n410 585
R1218 B.n409 B.n212 585
R1219 B.n408 B.n407 585
R1220 B.n406 B.n213 585
R1221 B.n405 B.n404 585
R1222 B.n403 B.n214 585
R1223 B.n402 B.n401 585
R1224 B.n400 B.n215 585
R1225 B.n399 B.n398 585
R1226 B.n397 B.n216 585
R1227 B.n396 B.n395 585
R1228 B.n394 B.n217 585
R1229 B.n393 B.n392 585
R1230 B.n391 B.n218 585
R1231 B.n390 B.n389 585
R1232 B.n388 B.n219 585
R1233 B.n387 B.n386 585
R1234 B.n385 B.n220 585
R1235 B.n518 B.n175 585
R1236 B.n520 B.n519 585
R1237 B.n521 B.n174 585
R1238 B.n523 B.n522 585
R1239 B.n524 B.n173 585
R1240 B.n526 B.n525 585
R1241 B.n527 B.n172 585
R1242 B.n529 B.n528 585
R1243 B.n530 B.n171 585
R1244 B.n532 B.n531 585
R1245 B.n533 B.n170 585
R1246 B.n535 B.n534 585
R1247 B.n536 B.n169 585
R1248 B.n538 B.n537 585
R1249 B.n539 B.n168 585
R1250 B.n541 B.n540 585
R1251 B.n542 B.n167 585
R1252 B.n544 B.n543 585
R1253 B.n545 B.n166 585
R1254 B.n547 B.n546 585
R1255 B.n548 B.n165 585
R1256 B.n550 B.n549 585
R1257 B.n551 B.n164 585
R1258 B.n553 B.n552 585
R1259 B.n554 B.n163 585
R1260 B.n556 B.n555 585
R1261 B.n557 B.n162 585
R1262 B.n559 B.n558 585
R1263 B.n560 B.n161 585
R1264 B.n562 B.n561 585
R1265 B.n563 B.n160 585
R1266 B.n565 B.n564 585
R1267 B.n566 B.n159 585
R1268 B.n568 B.n567 585
R1269 B.n569 B.n158 585
R1270 B.n571 B.n570 585
R1271 B.n572 B.n157 585
R1272 B.n574 B.n573 585
R1273 B.n575 B.n156 585
R1274 B.n577 B.n576 585
R1275 B.n578 B.n155 585
R1276 B.n580 B.n579 585
R1277 B.n581 B.n154 585
R1278 B.n583 B.n582 585
R1279 B.n584 B.n153 585
R1280 B.n586 B.n585 585
R1281 B.n587 B.n152 585
R1282 B.n589 B.n588 585
R1283 B.n590 B.n151 585
R1284 B.n592 B.n591 585
R1285 B.n593 B.n150 585
R1286 B.n595 B.n594 585
R1287 B.n596 B.n149 585
R1288 B.n598 B.n597 585
R1289 B.n599 B.n148 585
R1290 B.n601 B.n600 585
R1291 B.n602 B.n147 585
R1292 B.n604 B.n603 585
R1293 B.n605 B.n146 585
R1294 B.n607 B.n606 585
R1295 B.n608 B.n145 585
R1296 B.n610 B.n609 585
R1297 B.n611 B.n144 585
R1298 B.n613 B.n612 585
R1299 B.n614 B.n143 585
R1300 B.n616 B.n615 585
R1301 B.n617 B.n142 585
R1302 B.n619 B.n618 585
R1303 B.n620 B.n141 585
R1304 B.n622 B.n621 585
R1305 B.n623 B.n140 585
R1306 B.n625 B.n624 585
R1307 B.n626 B.n139 585
R1308 B.n628 B.n627 585
R1309 B.n629 B.n138 585
R1310 B.n631 B.n630 585
R1311 B.n632 B.n137 585
R1312 B.n634 B.n633 585
R1313 B.n635 B.n136 585
R1314 B.n637 B.n636 585
R1315 B.n638 B.n135 585
R1316 B.n640 B.n639 585
R1317 B.n641 B.n134 585
R1318 B.n643 B.n642 585
R1319 B.n644 B.n133 585
R1320 B.n646 B.n645 585
R1321 B.n647 B.n132 585
R1322 B.n649 B.n648 585
R1323 B.n650 B.n131 585
R1324 B.n652 B.n651 585
R1325 B.n653 B.n130 585
R1326 B.n655 B.n654 585
R1327 B.n656 B.n129 585
R1328 B.n658 B.n657 585
R1329 B.n659 B.n128 585
R1330 B.n661 B.n660 585
R1331 B.n662 B.n127 585
R1332 B.n664 B.n663 585
R1333 B.n665 B.n126 585
R1334 B.n667 B.n666 585
R1335 B.n668 B.n125 585
R1336 B.n670 B.n669 585
R1337 B.n671 B.n124 585
R1338 B.n673 B.n672 585
R1339 B.n674 B.n123 585
R1340 B.n676 B.n675 585
R1341 B.n677 B.n122 585
R1342 B.n679 B.n678 585
R1343 B.n680 B.n121 585
R1344 B.n682 B.n681 585
R1345 B.n683 B.n120 585
R1346 B.n685 B.n684 585
R1347 B.n686 B.n119 585
R1348 B.n688 B.n687 585
R1349 B.n689 B.n118 585
R1350 B.n691 B.n690 585
R1351 B.n692 B.n117 585
R1352 B.n694 B.n693 585
R1353 B.n695 B.n116 585
R1354 B.n697 B.n696 585
R1355 B.n698 B.n115 585
R1356 B.n700 B.n699 585
R1357 B.n701 B.n114 585
R1358 B.n703 B.n702 585
R1359 B.n704 B.n113 585
R1360 B.n706 B.n705 585
R1361 B.n707 B.n112 585
R1362 B.n709 B.n708 585
R1363 B.n710 B.n111 585
R1364 B.n712 B.n711 585
R1365 B.n713 B.n110 585
R1366 B.n715 B.n714 585
R1367 B.n716 B.n109 585
R1368 B.n718 B.n717 585
R1369 B.n719 B.n108 585
R1370 B.n721 B.n720 585
R1371 B.n722 B.n107 585
R1372 B.n724 B.n723 585
R1373 B.n725 B.n106 585
R1374 B.n727 B.n726 585
R1375 B.n728 B.n105 585
R1376 B.n730 B.n729 585
R1377 B.n731 B.n104 585
R1378 B.n733 B.n732 585
R1379 B.n734 B.n103 585
R1380 B.n736 B.n735 585
R1381 B.n737 B.n102 585
R1382 B.n739 B.n738 585
R1383 B.n740 B.n101 585
R1384 B.n742 B.n741 585
R1385 B.n743 B.n100 585
R1386 B.n745 B.n744 585
R1387 B.n746 B.n99 585
R1388 B.n748 B.n747 585
R1389 B.n749 B.n98 585
R1390 B.n751 B.n750 585
R1391 B.n752 B.n97 585
R1392 B.n754 B.n753 585
R1393 B.n755 B.n96 585
R1394 B.n757 B.n756 585
R1395 B.n758 B.n95 585
R1396 B.n760 B.n759 585
R1397 B.n761 B.n94 585
R1398 B.n763 B.n762 585
R1399 B.n764 B.n93 585
R1400 B.n766 B.n765 585
R1401 B.n767 B.n92 585
R1402 B.n769 B.n768 585
R1403 B.n899 B.n898 585
R1404 B.n897 B.n44 585
R1405 B.n896 B.n895 585
R1406 B.n894 B.n45 585
R1407 B.n893 B.n892 585
R1408 B.n891 B.n46 585
R1409 B.n890 B.n889 585
R1410 B.n888 B.n47 585
R1411 B.n887 B.n886 585
R1412 B.n885 B.n48 585
R1413 B.n884 B.n883 585
R1414 B.n882 B.n49 585
R1415 B.n881 B.n880 585
R1416 B.n879 B.n50 585
R1417 B.n878 B.n877 585
R1418 B.n876 B.n51 585
R1419 B.n875 B.n874 585
R1420 B.n873 B.n52 585
R1421 B.n872 B.n871 585
R1422 B.n870 B.n53 585
R1423 B.n869 B.n868 585
R1424 B.n867 B.n54 585
R1425 B.n866 B.n865 585
R1426 B.n864 B.n55 585
R1427 B.n863 B.n862 585
R1428 B.n861 B.n56 585
R1429 B.n860 B.n859 585
R1430 B.n858 B.n57 585
R1431 B.n857 B.n856 585
R1432 B.n855 B.n58 585
R1433 B.n854 B.n853 585
R1434 B.n852 B.n59 585
R1435 B.n851 B.n850 585
R1436 B.n849 B.n60 585
R1437 B.n848 B.n847 585
R1438 B.n846 B.n61 585
R1439 B.n845 B.n844 585
R1440 B.n843 B.n62 585
R1441 B.n842 B.n841 585
R1442 B.n840 B.n63 585
R1443 B.n839 B.n838 585
R1444 B.n837 B.n67 585
R1445 B.n836 B.n835 585
R1446 B.n834 B.n68 585
R1447 B.n833 B.n832 585
R1448 B.n831 B.n69 585
R1449 B.n830 B.n829 585
R1450 B.n828 B.n70 585
R1451 B.n826 B.n825 585
R1452 B.n824 B.n73 585
R1453 B.n823 B.n822 585
R1454 B.n821 B.n74 585
R1455 B.n820 B.n819 585
R1456 B.n818 B.n75 585
R1457 B.n817 B.n816 585
R1458 B.n815 B.n76 585
R1459 B.n814 B.n813 585
R1460 B.n812 B.n77 585
R1461 B.n811 B.n810 585
R1462 B.n809 B.n78 585
R1463 B.n808 B.n807 585
R1464 B.n806 B.n79 585
R1465 B.n805 B.n804 585
R1466 B.n803 B.n80 585
R1467 B.n802 B.n801 585
R1468 B.n800 B.n81 585
R1469 B.n799 B.n798 585
R1470 B.n797 B.n82 585
R1471 B.n796 B.n795 585
R1472 B.n794 B.n83 585
R1473 B.n793 B.n792 585
R1474 B.n791 B.n84 585
R1475 B.n790 B.n789 585
R1476 B.n788 B.n85 585
R1477 B.n787 B.n786 585
R1478 B.n785 B.n86 585
R1479 B.n784 B.n783 585
R1480 B.n782 B.n87 585
R1481 B.n781 B.n780 585
R1482 B.n779 B.n88 585
R1483 B.n778 B.n777 585
R1484 B.n776 B.n89 585
R1485 B.n775 B.n774 585
R1486 B.n773 B.n90 585
R1487 B.n772 B.n771 585
R1488 B.n770 B.n91 585
R1489 B.n900 B.n43 585
R1490 B.n902 B.n901 585
R1491 B.n903 B.n42 585
R1492 B.n905 B.n904 585
R1493 B.n906 B.n41 585
R1494 B.n908 B.n907 585
R1495 B.n909 B.n40 585
R1496 B.n911 B.n910 585
R1497 B.n912 B.n39 585
R1498 B.n914 B.n913 585
R1499 B.n915 B.n38 585
R1500 B.n917 B.n916 585
R1501 B.n918 B.n37 585
R1502 B.n920 B.n919 585
R1503 B.n921 B.n36 585
R1504 B.n923 B.n922 585
R1505 B.n924 B.n35 585
R1506 B.n926 B.n925 585
R1507 B.n927 B.n34 585
R1508 B.n929 B.n928 585
R1509 B.n930 B.n33 585
R1510 B.n932 B.n931 585
R1511 B.n933 B.n32 585
R1512 B.n935 B.n934 585
R1513 B.n936 B.n31 585
R1514 B.n938 B.n937 585
R1515 B.n939 B.n30 585
R1516 B.n941 B.n940 585
R1517 B.n942 B.n29 585
R1518 B.n944 B.n943 585
R1519 B.n945 B.n28 585
R1520 B.n947 B.n946 585
R1521 B.n948 B.n27 585
R1522 B.n950 B.n949 585
R1523 B.n951 B.n26 585
R1524 B.n953 B.n952 585
R1525 B.n954 B.n25 585
R1526 B.n956 B.n955 585
R1527 B.n957 B.n24 585
R1528 B.n959 B.n958 585
R1529 B.n960 B.n23 585
R1530 B.n962 B.n961 585
R1531 B.n963 B.n22 585
R1532 B.n965 B.n964 585
R1533 B.n966 B.n21 585
R1534 B.n968 B.n967 585
R1535 B.n969 B.n20 585
R1536 B.n971 B.n970 585
R1537 B.n972 B.n19 585
R1538 B.n974 B.n973 585
R1539 B.n975 B.n18 585
R1540 B.n977 B.n976 585
R1541 B.n978 B.n17 585
R1542 B.n980 B.n979 585
R1543 B.n981 B.n16 585
R1544 B.n983 B.n982 585
R1545 B.n984 B.n15 585
R1546 B.n986 B.n985 585
R1547 B.n987 B.n14 585
R1548 B.n989 B.n988 585
R1549 B.n990 B.n13 585
R1550 B.n992 B.n991 585
R1551 B.n993 B.n12 585
R1552 B.n995 B.n994 585
R1553 B.n996 B.n11 585
R1554 B.n998 B.n997 585
R1555 B.n999 B.n10 585
R1556 B.n1001 B.n1000 585
R1557 B.n1002 B.n9 585
R1558 B.n1004 B.n1003 585
R1559 B.n1005 B.n8 585
R1560 B.n1007 B.n1006 585
R1561 B.n1008 B.n7 585
R1562 B.n1010 B.n1009 585
R1563 B.n1011 B.n6 585
R1564 B.n1013 B.n1012 585
R1565 B.n1014 B.n5 585
R1566 B.n1016 B.n1015 585
R1567 B.n1017 B.n4 585
R1568 B.n1019 B.n1018 585
R1569 B.n1020 B.n3 585
R1570 B.n1022 B.n1021 585
R1571 B.n1023 B.n0 585
R1572 B.n2 B.n1 585
R1573 B.n262 B.n261 585
R1574 B.n264 B.n263 585
R1575 B.n265 B.n260 585
R1576 B.n267 B.n266 585
R1577 B.n268 B.n259 585
R1578 B.n270 B.n269 585
R1579 B.n271 B.n258 585
R1580 B.n273 B.n272 585
R1581 B.n274 B.n257 585
R1582 B.n276 B.n275 585
R1583 B.n277 B.n256 585
R1584 B.n279 B.n278 585
R1585 B.n280 B.n255 585
R1586 B.n282 B.n281 585
R1587 B.n283 B.n254 585
R1588 B.n285 B.n284 585
R1589 B.n286 B.n253 585
R1590 B.n288 B.n287 585
R1591 B.n289 B.n252 585
R1592 B.n291 B.n290 585
R1593 B.n292 B.n251 585
R1594 B.n294 B.n293 585
R1595 B.n295 B.n250 585
R1596 B.n297 B.n296 585
R1597 B.n298 B.n249 585
R1598 B.n300 B.n299 585
R1599 B.n301 B.n248 585
R1600 B.n303 B.n302 585
R1601 B.n304 B.n247 585
R1602 B.n306 B.n305 585
R1603 B.n307 B.n246 585
R1604 B.n309 B.n308 585
R1605 B.n310 B.n245 585
R1606 B.n312 B.n311 585
R1607 B.n313 B.n244 585
R1608 B.n315 B.n314 585
R1609 B.n316 B.n243 585
R1610 B.n318 B.n317 585
R1611 B.n319 B.n242 585
R1612 B.n321 B.n320 585
R1613 B.n322 B.n241 585
R1614 B.n324 B.n323 585
R1615 B.n325 B.n240 585
R1616 B.n327 B.n326 585
R1617 B.n328 B.n239 585
R1618 B.n330 B.n329 585
R1619 B.n331 B.n238 585
R1620 B.n333 B.n332 585
R1621 B.n334 B.n237 585
R1622 B.n336 B.n335 585
R1623 B.n337 B.n236 585
R1624 B.n339 B.n338 585
R1625 B.n340 B.n235 585
R1626 B.n342 B.n341 585
R1627 B.n343 B.n234 585
R1628 B.n345 B.n344 585
R1629 B.n346 B.n233 585
R1630 B.n348 B.n347 585
R1631 B.n349 B.n232 585
R1632 B.n351 B.n350 585
R1633 B.n352 B.n231 585
R1634 B.n354 B.n353 585
R1635 B.n355 B.n230 585
R1636 B.n357 B.n356 585
R1637 B.n358 B.n229 585
R1638 B.n360 B.n359 585
R1639 B.n361 B.n228 585
R1640 B.n363 B.n362 585
R1641 B.n364 B.n227 585
R1642 B.n366 B.n365 585
R1643 B.n367 B.n226 585
R1644 B.n369 B.n368 585
R1645 B.n370 B.n225 585
R1646 B.n372 B.n371 585
R1647 B.n373 B.n224 585
R1648 B.n375 B.n374 585
R1649 B.n376 B.n223 585
R1650 B.n378 B.n377 585
R1651 B.n379 B.n222 585
R1652 B.n381 B.n380 585
R1653 B.n382 B.n221 585
R1654 B.n384 B.n383 585
R1655 B.n383 B.n220 444.452
R1656 B.n518 B.n517 444.452
R1657 B.n770 B.n769 444.452
R1658 B.n898 B.n43 444.452
R1659 B.n195 B.t7 436.762
R1660 B.n71 B.t2 436.762
R1661 B.n440 B.t10 436.762
R1662 B.n64 B.t5 436.762
R1663 B.n196 B.t8 354.144
R1664 B.n72 B.t1 354.144
R1665 B.n441 B.t11 354.144
R1666 B.n65 B.t4 354.144
R1667 B.n440 B.t9 275.671
R1668 B.n195 B.t6 275.671
R1669 B.n71 B.t0 275.671
R1670 B.n64 B.t3 275.671
R1671 B.n1025 B.n1024 256.663
R1672 B.n1024 B.n1023 235.042
R1673 B.n1024 B.n2 235.042
R1674 B.n387 B.n220 163.367
R1675 B.n388 B.n387 163.367
R1676 B.n389 B.n388 163.367
R1677 B.n389 B.n218 163.367
R1678 B.n393 B.n218 163.367
R1679 B.n394 B.n393 163.367
R1680 B.n395 B.n394 163.367
R1681 B.n395 B.n216 163.367
R1682 B.n399 B.n216 163.367
R1683 B.n400 B.n399 163.367
R1684 B.n401 B.n400 163.367
R1685 B.n401 B.n214 163.367
R1686 B.n405 B.n214 163.367
R1687 B.n406 B.n405 163.367
R1688 B.n407 B.n406 163.367
R1689 B.n407 B.n212 163.367
R1690 B.n411 B.n212 163.367
R1691 B.n412 B.n411 163.367
R1692 B.n413 B.n412 163.367
R1693 B.n413 B.n210 163.367
R1694 B.n417 B.n210 163.367
R1695 B.n418 B.n417 163.367
R1696 B.n419 B.n418 163.367
R1697 B.n419 B.n208 163.367
R1698 B.n423 B.n208 163.367
R1699 B.n424 B.n423 163.367
R1700 B.n425 B.n424 163.367
R1701 B.n425 B.n206 163.367
R1702 B.n429 B.n206 163.367
R1703 B.n430 B.n429 163.367
R1704 B.n431 B.n430 163.367
R1705 B.n431 B.n204 163.367
R1706 B.n435 B.n204 163.367
R1707 B.n436 B.n435 163.367
R1708 B.n437 B.n436 163.367
R1709 B.n437 B.n202 163.367
R1710 B.n444 B.n202 163.367
R1711 B.n445 B.n444 163.367
R1712 B.n446 B.n445 163.367
R1713 B.n446 B.n200 163.367
R1714 B.n450 B.n200 163.367
R1715 B.n451 B.n450 163.367
R1716 B.n452 B.n451 163.367
R1717 B.n452 B.n198 163.367
R1718 B.n456 B.n198 163.367
R1719 B.n457 B.n456 163.367
R1720 B.n458 B.n457 163.367
R1721 B.n458 B.n194 163.367
R1722 B.n463 B.n194 163.367
R1723 B.n464 B.n463 163.367
R1724 B.n465 B.n464 163.367
R1725 B.n465 B.n192 163.367
R1726 B.n469 B.n192 163.367
R1727 B.n470 B.n469 163.367
R1728 B.n471 B.n470 163.367
R1729 B.n471 B.n190 163.367
R1730 B.n475 B.n190 163.367
R1731 B.n476 B.n475 163.367
R1732 B.n477 B.n476 163.367
R1733 B.n477 B.n188 163.367
R1734 B.n481 B.n188 163.367
R1735 B.n482 B.n481 163.367
R1736 B.n483 B.n482 163.367
R1737 B.n483 B.n186 163.367
R1738 B.n487 B.n186 163.367
R1739 B.n488 B.n487 163.367
R1740 B.n489 B.n488 163.367
R1741 B.n489 B.n184 163.367
R1742 B.n493 B.n184 163.367
R1743 B.n494 B.n493 163.367
R1744 B.n495 B.n494 163.367
R1745 B.n495 B.n182 163.367
R1746 B.n499 B.n182 163.367
R1747 B.n500 B.n499 163.367
R1748 B.n501 B.n500 163.367
R1749 B.n501 B.n180 163.367
R1750 B.n505 B.n180 163.367
R1751 B.n506 B.n505 163.367
R1752 B.n507 B.n506 163.367
R1753 B.n507 B.n178 163.367
R1754 B.n511 B.n178 163.367
R1755 B.n512 B.n511 163.367
R1756 B.n513 B.n512 163.367
R1757 B.n513 B.n176 163.367
R1758 B.n517 B.n176 163.367
R1759 B.n769 B.n92 163.367
R1760 B.n765 B.n92 163.367
R1761 B.n765 B.n764 163.367
R1762 B.n764 B.n763 163.367
R1763 B.n763 B.n94 163.367
R1764 B.n759 B.n94 163.367
R1765 B.n759 B.n758 163.367
R1766 B.n758 B.n757 163.367
R1767 B.n757 B.n96 163.367
R1768 B.n753 B.n96 163.367
R1769 B.n753 B.n752 163.367
R1770 B.n752 B.n751 163.367
R1771 B.n751 B.n98 163.367
R1772 B.n747 B.n98 163.367
R1773 B.n747 B.n746 163.367
R1774 B.n746 B.n745 163.367
R1775 B.n745 B.n100 163.367
R1776 B.n741 B.n100 163.367
R1777 B.n741 B.n740 163.367
R1778 B.n740 B.n739 163.367
R1779 B.n739 B.n102 163.367
R1780 B.n735 B.n102 163.367
R1781 B.n735 B.n734 163.367
R1782 B.n734 B.n733 163.367
R1783 B.n733 B.n104 163.367
R1784 B.n729 B.n104 163.367
R1785 B.n729 B.n728 163.367
R1786 B.n728 B.n727 163.367
R1787 B.n727 B.n106 163.367
R1788 B.n723 B.n106 163.367
R1789 B.n723 B.n722 163.367
R1790 B.n722 B.n721 163.367
R1791 B.n721 B.n108 163.367
R1792 B.n717 B.n108 163.367
R1793 B.n717 B.n716 163.367
R1794 B.n716 B.n715 163.367
R1795 B.n715 B.n110 163.367
R1796 B.n711 B.n110 163.367
R1797 B.n711 B.n710 163.367
R1798 B.n710 B.n709 163.367
R1799 B.n709 B.n112 163.367
R1800 B.n705 B.n112 163.367
R1801 B.n705 B.n704 163.367
R1802 B.n704 B.n703 163.367
R1803 B.n703 B.n114 163.367
R1804 B.n699 B.n114 163.367
R1805 B.n699 B.n698 163.367
R1806 B.n698 B.n697 163.367
R1807 B.n697 B.n116 163.367
R1808 B.n693 B.n116 163.367
R1809 B.n693 B.n692 163.367
R1810 B.n692 B.n691 163.367
R1811 B.n691 B.n118 163.367
R1812 B.n687 B.n118 163.367
R1813 B.n687 B.n686 163.367
R1814 B.n686 B.n685 163.367
R1815 B.n685 B.n120 163.367
R1816 B.n681 B.n120 163.367
R1817 B.n681 B.n680 163.367
R1818 B.n680 B.n679 163.367
R1819 B.n679 B.n122 163.367
R1820 B.n675 B.n122 163.367
R1821 B.n675 B.n674 163.367
R1822 B.n674 B.n673 163.367
R1823 B.n673 B.n124 163.367
R1824 B.n669 B.n124 163.367
R1825 B.n669 B.n668 163.367
R1826 B.n668 B.n667 163.367
R1827 B.n667 B.n126 163.367
R1828 B.n663 B.n126 163.367
R1829 B.n663 B.n662 163.367
R1830 B.n662 B.n661 163.367
R1831 B.n661 B.n128 163.367
R1832 B.n657 B.n128 163.367
R1833 B.n657 B.n656 163.367
R1834 B.n656 B.n655 163.367
R1835 B.n655 B.n130 163.367
R1836 B.n651 B.n130 163.367
R1837 B.n651 B.n650 163.367
R1838 B.n650 B.n649 163.367
R1839 B.n649 B.n132 163.367
R1840 B.n645 B.n132 163.367
R1841 B.n645 B.n644 163.367
R1842 B.n644 B.n643 163.367
R1843 B.n643 B.n134 163.367
R1844 B.n639 B.n134 163.367
R1845 B.n639 B.n638 163.367
R1846 B.n638 B.n637 163.367
R1847 B.n637 B.n136 163.367
R1848 B.n633 B.n136 163.367
R1849 B.n633 B.n632 163.367
R1850 B.n632 B.n631 163.367
R1851 B.n631 B.n138 163.367
R1852 B.n627 B.n138 163.367
R1853 B.n627 B.n626 163.367
R1854 B.n626 B.n625 163.367
R1855 B.n625 B.n140 163.367
R1856 B.n621 B.n140 163.367
R1857 B.n621 B.n620 163.367
R1858 B.n620 B.n619 163.367
R1859 B.n619 B.n142 163.367
R1860 B.n615 B.n142 163.367
R1861 B.n615 B.n614 163.367
R1862 B.n614 B.n613 163.367
R1863 B.n613 B.n144 163.367
R1864 B.n609 B.n144 163.367
R1865 B.n609 B.n608 163.367
R1866 B.n608 B.n607 163.367
R1867 B.n607 B.n146 163.367
R1868 B.n603 B.n146 163.367
R1869 B.n603 B.n602 163.367
R1870 B.n602 B.n601 163.367
R1871 B.n601 B.n148 163.367
R1872 B.n597 B.n148 163.367
R1873 B.n597 B.n596 163.367
R1874 B.n596 B.n595 163.367
R1875 B.n595 B.n150 163.367
R1876 B.n591 B.n150 163.367
R1877 B.n591 B.n590 163.367
R1878 B.n590 B.n589 163.367
R1879 B.n589 B.n152 163.367
R1880 B.n585 B.n152 163.367
R1881 B.n585 B.n584 163.367
R1882 B.n584 B.n583 163.367
R1883 B.n583 B.n154 163.367
R1884 B.n579 B.n154 163.367
R1885 B.n579 B.n578 163.367
R1886 B.n578 B.n577 163.367
R1887 B.n577 B.n156 163.367
R1888 B.n573 B.n156 163.367
R1889 B.n573 B.n572 163.367
R1890 B.n572 B.n571 163.367
R1891 B.n571 B.n158 163.367
R1892 B.n567 B.n158 163.367
R1893 B.n567 B.n566 163.367
R1894 B.n566 B.n565 163.367
R1895 B.n565 B.n160 163.367
R1896 B.n561 B.n160 163.367
R1897 B.n561 B.n560 163.367
R1898 B.n560 B.n559 163.367
R1899 B.n559 B.n162 163.367
R1900 B.n555 B.n162 163.367
R1901 B.n555 B.n554 163.367
R1902 B.n554 B.n553 163.367
R1903 B.n553 B.n164 163.367
R1904 B.n549 B.n164 163.367
R1905 B.n549 B.n548 163.367
R1906 B.n548 B.n547 163.367
R1907 B.n547 B.n166 163.367
R1908 B.n543 B.n166 163.367
R1909 B.n543 B.n542 163.367
R1910 B.n542 B.n541 163.367
R1911 B.n541 B.n168 163.367
R1912 B.n537 B.n168 163.367
R1913 B.n537 B.n536 163.367
R1914 B.n536 B.n535 163.367
R1915 B.n535 B.n170 163.367
R1916 B.n531 B.n170 163.367
R1917 B.n531 B.n530 163.367
R1918 B.n530 B.n529 163.367
R1919 B.n529 B.n172 163.367
R1920 B.n525 B.n172 163.367
R1921 B.n525 B.n524 163.367
R1922 B.n524 B.n523 163.367
R1923 B.n523 B.n174 163.367
R1924 B.n519 B.n174 163.367
R1925 B.n519 B.n518 163.367
R1926 B.n898 B.n897 163.367
R1927 B.n897 B.n896 163.367
R1928 B.n896 B.n45 163.367
R1929 B.n892 B.n45 163.367
R1930 B.n892 B.n891 163.367
R1931 B.n891 B.n890 163.367
R1932 B.n890 B.n47 163.367
R1933 B.n886 B.n47 163.367
R1934 B.n886 B.n885 163.367
R1935 B.n885 B.n884 163.367
R1936 B.n884 B.n49 163.367
R1937 B.n880 B.n49 163.367
R1938 B.n880 B.n879 163.367
R1939 B.n879 B.n878 163.367
R1940 B.n878 B.n51 163.367
R1941 B.n874 B.n51 163.367
R1942 B.n874 B.n873 163.367
R1943 B.n873 B.n872 163.367
R1944 B.n872 B.n53 163.367
R1945 B.n868 B.n53 163.367
R1946 B.n868 B.n867 163.367
R1947 B.n867 B.n866 163.367
R1948 B.n866 B.n55 163.367
R1949 B.n862 B.n55 163.367
R1950 B.n862 B.n861 163.367
R1951 B.n861 B.n860 163.367
R1952 B.n860 B.n57 163.367
R1953 B.n856 B.n57 163.367
R1954 B.n856 B.n855 163.367
R1955 B.n855 B.n854 163.367
R1956 B.n854 B.n59 163.367
R1957 B.n850 B.n59 163.367
R1958 B.n850 B.n849 163.367
R1959 B.n849 B.n848 163.367
R1960 B.n848 B.n61 163.367
R1961 B.n844 B.n61 163.367
R1962 B.n844 B.n843 163.367
R1963 B.n843 B.n842 163.367
R1964 B.n842 B.n63 163.367
R1965 B.n838 B.n63 163.367
R1966 B.n838 B.n837 163.367
R1967 B.n837 B.n836 163.367
R1968 B.n836 B.n68 163.367
R1969 B.n832 B.n68 163.367
R1970 B.n832 B.n831 163.367
R1971 B.n831 B.n830 163.367
R1972 B.n830 B.n70 163.367
R1973 B.n825 B.n70 163.367
R1974 B.n825 B.n824 163.367
R1975 B.n824 B.n823 163.367
R1976 B.n823 B.n74 163.367
R1977 B.n819 B.n74 163.367
R1978 B.n819 B.n818 163.367
R1979 B.n818 B.n817 163.367
R1980 B.n817 B.n76 163.367
R1981 B.n813 B.n76 163.367
R1982 B.n813 B.n812 163.367
R1983 B.n812 B.n811 163.367
R1984 B.n811 B.n78 163.367
R1985 B.n807 B.n78 163.367
R1986 B.n807 B.n806 163.367
R1987 B.n806 B.n805 163.367
R1988 B.n805 B.n80 163.367
R1989 B.n801 B.n80 163.367
R1990 B.n801 B.n800 163.367
R1991 B.n800 B.n799 163.367
R1992 B.n799 B.n82 163.367
R1993 B.n795 B.n82 163.367
R1994 B.n795 B.n794 163.367
R1995 B.n794 B.n793 163.367
R1996 B.n793 B.n84 163.367
R1997 B.n789 B.n84 163.367
R1998 B.n789 B.n788 163.367
R1999 B.n788 B.n787 163.367
R2000 B.n787 B.n86 163.367
R2001 B.n783 B.n86 163.367
R2002 B.n783 B.n782 163.367
R2003 B.n782 B.n781 163.367
R2004 B.n781 B.n88 163.367
R2005 B.n777 B.n88 163.367
R2006 B.n777 B.n776 163.367
R2007 B.n776 B.n775 163.367
R2008 B.n775 B.n90 163.367
R2009 B.n771 B.n90 163.367
R2010 B.n771 B.n770 163.367
R2011 B.n902 B.n43 163.367
R2012 B.n903 B.n902 163.367
R2013 B.n904 B.n903 163.367
R2014 B.n904 B.n41 163.367
R2015 B.n908 B.n41 163.367
R2016 B.n909 B.n908 163.367
R2017 B.n910 B.n909 163.367
R2018 B.n910 B.n39 163.367
R2019 B.n914 B.n39 163.367
R2020 B.n915 B.n914 163.367
R2021 B.n916 B.n915 163.367
R2022 B.n916 B.n37 163.367
R2023 B.n920 B.n37 163.367
R2024 B.n921 B.n920 163.367
R2025 B.n922 B.n921 163.367
R2026 B.n922 B.n35 163.367
R2027 B.n926 B.n35 163.367
R2028 B.n927 B.n926 163.367
R2029 B.n928 B.n927 163.367
R2030 B.n928 B.n33 163.367
R2031 B.n932 B.n33 163.367
R2032 B.n933 B.n932 163.367
R2033 B.n934 B.n933 163.367
R2034 B.n934 B.n31 163.367
R2035 B.n938 B.n31 163.367
R2036 B.n939 B.n938 163.367
R2037 B.n940 B.n939 163.367
R2038 B.n940 B.n29 163.367
R2039 B.n944 B.n29 163.367
R2040 B.n945 B.n944 163.367
R2041 B.n946 B.n945 163.367
R2042 B.n946 B.n27 163.367
R2043 B.n950 B.n27 163.367
R2044 B.n951 B.n950 163.367
R2045 B.n952 B.n951 163.367
R2046 B.n952 B.n25 163.367
R2047 B.n956 B.n25 163.367
R2048 B.n957 B.n956 163.367
R2049 B.n958 B.n957 163.367
R2050 B.n958 B.n23 163.367
R2051 B.n962 B.n23 163.367
R2052 B.n963 B.n962 163.367
R2053 B.n964 B.n963 163.367
R2054 B.n964 B.n21 163.367
R2055 B.n968 B.n21 163.367
R2056 B.n969 B.n968 163.367
R2057 B.n970 B.n969 163.367
R2058 B.n970 B.n19 163.367
R2059 B.n974 B.n19 163.367
R2060 B.n975 B.n974 163.367
R2061 B.n976 B.n975 163.367
R2062 B.n976 B.n17 163.367
R2063 B.n980 B.n17 163.367
R2064 B.n981 B.n980 163.367
R2065 B.n982 B.n981 163.367
R2066 B.n982 B.n15 163.367
R2067 B.n986 B.n15 163.367
R2068 B.n987 B.n986 163.367
R2069 B.n988 B.n987 163.367
R2070 B.n988 B.n13 163.367
R2071 B.n992 B.n13 163.367
R2072 B.n993 B.n992 163.367
R2073 B.n994 B.n993 163.367
R2074 B.n994 B.n11 163.367
R2075 B.n998 B.n11 163.367
R2076 B.n999 B.n998 163.367
R2077 B.n1000 B.n999 163.367
R2078 B.n1000 B.n9 163.367
R2079 B.n1004 B.n9 163.367
R2080 B.n1005 B.n1004 163.367
R2081 B.n1006 B.n1005 163.367
R2082 B.n1006 B.n7 163.367
R2083 B.n1010 B.n7 163.367
R2084 B.n1011 B.n1010 163.367
R2085 B.n1012 B.n1011 163.367
R2086 B.n1012 B.n5 163.367
R2087 B.n1016 B.n5 163.367
R2088 B.n1017 B.n1016 163.367
R2089 B.n1018 B.n1017 163.367
R2090 B.n1018 B.n3 163.367
R2091 B.n1022 B.n3 163.367
R2092 B.n1023 B.n1022 163.367
R2093 B.n262 B.n2 163.367
R2094 B.n263 B.n262 163.367
R2095 B.n263 B.n260 163.367
R2096 B.n267 B.n260 163.367
R2097 B.n268 B.n267 163.367
R2098 B.n269 B.n268 163.367
R2099 B.n269 B.n258 163.367
R2100 B.n273 B.n258 163.367
R2101 B.n274 B.n273 163.367
R2102 B.n275 B.n274 163.367
R2103 B.n275 B.n256 163.367
R2104 B.n279 B.n256 163.367
R2105 B.n280 B.n279 163.367
R2106 B.n281 B.n280 163.367
R2107 B.n281 B.n254 163.367
R2108 B.n285 B.n254 163.367
R2109 B.n286 B.n285 163.367
R2110 B.n287 B.n286 163.367
R2111 B.n287 B.n252 163.367
R2112 B.n291 B.n252 163.367
R2113 B.n292 B.n291 163.367
R2114 B.n293 B.n292 163.367
R2115 B.n293 B.n250 163.367
R2116 B.n297 B.n250 163.367
R2117 B.n298 B.n297 163.367
R2118 B.n299 B.n298 163.367
R2119 B.n299 B.n248 163.367
R2120 B.n303 B.n248 163.367
R2121 B.n304 B.n303 163.367
R2122 B.n305 B.n304 163.367
R2123 B.n305 B.n246 163.367
R2124 B.n309 B.n246 163.367
R2125 B.n310 B.n309 163.367
R2126 B.n311 B.n310 163.367
R2127 B.n311 B.n244 163.367
R2128 B.n315 B.n244 163.367
R2129 B.n316 B.n315 163.367
R2130 B.n317 B.n316 163.367
R2131 B.n317 B.n242 163.367
R2132 B.n321 B.n242 163.367
R2133 B.n322 B.n321 163.367
R2134 B.n323 B.n322 163.367
R2135 B.n323 B.n240 163.367
R2136 B.n327 B.n240 163.367
R2137 B.n328 B.n327 163.367
R2138 B.n329 B.n328 163.367
R2139 B.n329 B.n238 163.367
R2140 B.n333 B.n238 163.367
R2141 B.n334 B.n333 163.367
R2142 B.n335 B.n334 163.367
R2143 B.n335 B.n236 163.367
R2144 B.n339 B.n236 163.367
R2145 B.n340 B.n339 163.367
R2146 B.n341 B.n340 163.367
R2147 B.n341 B.n234 163.367
R2148 B.n345 B.n234 163.367
R2149 B.n346 B.n345 163.367
R2150 B.n347 B.n346 163.367
R2151 B.n347 B.n232 163.367
R2152 B.n351 B.n232 163.367
R2153 B.n352 B.n351 163.367
R2154 B.n353 B.n352 163.367
R2155 B.n353 B.n230 163.367
R2156 B.n357 B.n230 163.367
R2157 B.n358 B.n357 163.367
R2158 B.n359 B.n358 163.367
R2159 B.n359 B.n228 163.367
R2160 B.n363 B.n228 163.367
R2161 B.n364 B.n363 163.367
R2162 B.n365 B.n364 163.367
R2163 B.n365 B.n226 163.367
R2164 B.n369 B.n226 163.367
R2165 B.n370 B.n369 163.367
R2166 B.n371 B.n370 163.367
R2167 B.n371 B.n224 163.367
R2168 B.n375 B.n224 163.367
R2169 B.n376 B.n375 163.367
R2170 B.n377 B.n376 163.367
R2171 B.n377 B.n222 163.367
R2172 B.n381 B.n222 163.367
R2173 B.n382 B.n381 163.367
R2174 B.n383 B.n382 163.367
R2175 B.n441 B.n440 82.6187
R2176 B.n196 B.n195 82.6187
R2177 B.n72 B.n71 82.6187
R2178 B.n65 B.n64 82.6187
R2179 B.n442 B.n441 59.5399
R2180 B.n460 B.n196 59.5399
R2181 B.n827 B.n72 59.5399
R2182 B.n66 B.n65 59.5399
R2183 B.n900 B.n899 28.8785
R2184 B.n768 B.n91 28.8785
R2185 B.n385 B.n384 28.8785
R2186 B.n516 B.n175 28.8785
R2187 B B.n1025 18.0485
R2188 B.n901 B.n900 10.6151
R2189 B.n901 B.n42 10.6151
R2190 B.n905 B.n42 10.6151
R2191 B.n906 B.n905 10.6151
R2192 B.n907 B.n906 10.6151
R2193 B.n907 B.n40 10.6151
R2194 B.n911 B.n40 10.6151
R2195 B.n912 B.n911 10.6151
R2196 B.n913 B.n912 10.6151
R2197 B.n913 B.n38 10.6151
R2198 B.n917 B.n38 10.6151
R2199 B.n918 B.n917 10.6151
R2200 B.n919 B.n918 10.6151
R2201 B.n919 B.n36 10.6151
R2202 B.n923 B.n36 10.6151
R2203 B.n924 B.n923 10.6151
R2204 B.n925 B.n924 10.6151
R2205 B.n925 B.n34 10.6151
R2206 B.n929 B.n34 10.6151
R2207 B.n930 B.n929 10.6151
R2208 B.n931 B.n930 10.6151
R2209 B.n931 B.n32 10.6151
R2210 B.n935 B.n32 10.6151
R2211 B.n936 B.n935 10.6151
R2212 B.n937 B.n936 10.6151
R2213 B.n937 B.n30 10.6151
R2214 B.n941 B.n30 10.6151
R2215 B.n942 B.n941 10.6151
R2216 B.n943 B.n942 10.6151
R2217 B.n943 B.n28 10.6151
R2218 B.n947 B.n28 10.6151
R2219 B.n948 B.n947 10.6151
R2220 B.n949 B.n948 10.6151
R2221 B.n949 B.n26 10.6151
R2222 B.n953 B.n26 10.6151
R2223 B.n954 B.n953 10.6151
R2224 B.n955 B.n954 10.6151
R2225 B.n955 B.n24 10.6151
R2226 B.n959 B.n24 10.6151
R2227 B.n960 B.n959 10.6151
R2228 B.n961 B.n960 10.6151
R2229 B.n961 B.n22 10.6151
R2230 B.n965 B.n22 10.6151
R2231 B.n966 B.n965 10.6151
R2232 B.n967 B.n966 10.6151
R2233 B.n967 B.n20 10.6151
R2234 B.n971 B.n20 10.6151
R2235 B.n972 B.n971 10.6151
R2236 B.n973 B.n972 10.6151
R2237 B.n973 B.n18 10.6151
R2238 B.n977 B.n18 10.6151
R2239 B.n978 B.n977 10.6151
R2240 B.n979 B.n978 10.6151
R2241 B.n979 B.n16 10.6151
R2242 B.n983 B.n16 10.6151
R2243 B.n984 B.n983 10.6151
R2244 B.n985 B.n984 10.6151
R2245 B.n985 B.n14 10.6151
R2246 B.n989 B.n14 10.6151
R2247 B.n990 B.n989 10.6151
R2248 B.n991 B.n990 10.6151
R2249 B.n991 B.n12 10.6151
R2250 B.n995 B.n12 10.6151
R2251 B.n996 B.n995 10.6151
R2252 B.n997 B.n996 10.6151
R2253 B.n997 B.n10 10.6151
R2254 B.n1001 B.n10 10.6151
R2255 B.n1002 B.n1001 10.6151
R2256 B.n1003 B.n1002 10.6151
R2257 B.n1003 B.n8 10.6151
R2258 B.n1007 B.n8 10.6151
R2259 B.n1008 B.n1007 10.6151
R2260 B.n1009 B.n1008 10.6151
R2261 B.n1009 B.n6 10.6151
R2262 B.n1013 B.n6 10.6151
R2263 B.n1014 B.n1013 10.6151
R2264 B.n1015 B.n1014 10.6151
R2265 B.n1015 B.n4 10.6151
R2266 B.n1019 B.n4 10.6151
R2267 B.n1020 B.n1019 10.6151
R2268 B.n1021 B.n1020 10.6151
R2269 B.n1021 B.n0 10.6151
R2270 B.n899 B.n44 10.6151
R2271 B.n895 B.n44 10.6151
R2272 B.n895 B.n894 10.6151
R2273 B.n894 B.n893 10.6151
R2274 B.n893 B.n46 10.6151
R2275 B.n889 B.n46 10.6151
R2276 B.n889 B.n888 10.6151
R2277 B.n888 B.n887 10.6151
R2278 B.n887 B.n48 10.6151
R2279 B.n883 B.n48 10.6151
R2280 B.n883 B.n882 10.6151
R2281 B.n882 B.n881 10.6151
R2282 B.n881 B.n50 10.6151
R2283 B.n877 B.n50 10.6151
R2284 B.n877 B.n876 10.6151
R2285 B.n876 B.n875 10.6151
R2286 B.n875 B.n52 10.6151
R2287 B.n871 B.n52 10.6151
R2288 B.n871 B.n870 10.6151
R2289 B.n870 B.n869 10.6151
R2290 B.n869 B.n54 10.6151
R2291 B.n865 B.n54 10.6151
R2292 B.n865 B.n864 10.6151
R2293 B.n864 B.n863 10.6151
R2294 B.n863 B.n56 10.6151
R2295 B.n859 B.n56 10.6151
R2296 B.n859 B.n858 10.6151
R2297 B.n858 B.n857 10.6151
R2298 B.n857 B.n58 10.6151
R2299 B.n853 B.n58 10.6151
R2300 B.n853 B.n852 10.6151
R2301 B.n852 B.n851 10.6151
R2302 B.n851 B.n60 10.6151
R2303 B.n847 B.n60 10.6151
R2304 B.n847 B.n846 10.6151
R2305 B.n846 B.n845 10.6151
R2306 B.n845 B.n62 10.6151
R2307 B.n841 B.n840 10.6151
R2308 B.n840 B.n839 10.6151
R2309 B.n839 B.n67 10.6151
R2310 B.n835 B.n67 10.6151
R2311 B.n835 B.n834 10.6151
R2312 B.n834 B.n833 10.6151
R2313 B.n833 B.n69 10.6151
R2314 B.n829 B.n69 10.6151
R2315 B.n829 B.n828 10.6151
R2316 B.n826 B.n73 10.6151
R2317 B.n822 B.n73 10.6151
R2318 B.n822 B.n821 10.6151
R2319 B.n821 B.n820 10.6151
R2320 B.n820 B.n75 10.6151
R2321 B.n816 B.n75 10.6151
R2322 B.n816 B.n815 10.6151
R2323 B.n815 B.n814 10.6151
R2324 B.n814 B.n77 10.6151
R2325 B.n810 B.n77 10.6151
R2326 B.n810 B.n809 10.6151
R2327 B.n809 B.n808 10.6151
R2328 B.n808 B.n79 10.6151
R2329 B.n804 B.n79 10.6151
R2330 B.n804 B.n803 10.6151
R2331 B.n803 B.n802 10.6151
R2332 B.n802 B.n81 10.6151
R2333 B.n798 B.n81 10.6151
R2334 B.n798 B.n797 10.6151
R2335 B.n797 B.n796 10.6151
R2336 B.n796 B.n83 10.6151
R2337 B.n792 B.n83 10.6151
R2338 B.n792 B.n791 10.6151
R2339 B.n791 B.n790 10.6151
R2340 B.n790 B.n85 10.6151
R2341 B.n786 B.n85 10.6151
R2342 B.n786 B.n785 10.6151
R2343 B.n785 B.n784 10.6151
R2344 B.n784 B.n87 10.6151
R2345 B.n780 B.n87 10.6151
R2346 B.n780 B.n779 10.6151
R2347 B.n779 B.n778 10.6151
R2348 B.n778 B.n89 10.6151
R2349 B.n774 B.n89 10.6151
R2350 B.n774 B.n773 10.6151
R2351 B.n773 B.n772 10.6151
R2352 B.n772 B.n91 10.6151
R2353 B.n768 B.n767 10.6151
R2354 B.n767 B.n766 10.6151
R2355 B.n766 B.n93 10.6151
R2356 B.n762 B.n93 10.6151
R2357 B.n762 B.n761 10.6151
R2358 B.n761 B.n760 10.6151
R2359 B.n760 B.n95 10.6151
R2360 B.n756 B.n95 10.6151
R2361 B.n756 B.n755 10.6151
R2362 B.n755 B.n754 10.6151
R2363 B.n754 B.n97 10.6151
R2364 B.n750 B.n97 10.6151
R2365 B.n750 B.n749 10.6151
R2366 B.n749 B.n748 10.6151
R2367 B.n748 B.n99 10.6151
R2368 B.n744 B.n99 10.6151
R2369 B.n744 B.n743 10.6151
R2370 B.n743 B.n742 10.6151
R2371 B.n742 B.n101 10.6151
R2372 B.n738 B.n101 10.6151
R2373 B.n738 B.n737 10.6151
R2374 B.n737 B.n736 10.6151
R2375 B.n736 B.n103 10.6151
R2376 B.n732 B.n103 10.6151
R2377 B.n732 B.n731 10.6151
R2378 B.n731 B.n730 10.6151
R2379 B.n730 B.n105 10.6151
R2380 B.n726 B.n105 10.6151
R2381 B.n726 B.n725 10.6151
R2382 B.n725 B.n724 10.6151
R2383 B.n724 B.n107 10.6151
R2384 B.n720 B.n107 10.6151
R2385 B.n720 B.n719 10.6151
R2386 B.n719 B.n718 10.6151
R2387 B.n718 B.n109 10.6151
R2388 B.n714 B.n109 10.6151
R2389 B.n714 B.n713 10.6151
R2390 B.n713 B.n712 10.6151
R2391 B.n712 B.n111 10.6151
R2392 B.n708 B.n111 10.6151
R2393 B.n708 B.n707 10.6151
R2394 B.n707 B.n706 10.6151
R2395 B.n706 B.n113 10.6151
R2396 B.n702 B.n113 10.6151
R2397 B.n702 B.n701 10.6151
R2398 B.n701 B.n700 10.6151
R2399 B.n700 B.n115 10.6151
R2400 B.n696 B.n115 10.6151
R2401 B.n696 B.n695 10.6151
R2402 B.n695 B.n694 10.6151
R2403 B.n694 B.n117 10.6151
R2404 B.n690 B.n117 10.6151
R2405 B.n690 B.n689 10.6151
R2406 B.n689 B.n688 10.6151
R2407 B.n688 B.n119 10.6151
R2408 B.n684 B.n119 10.6151
R2409 B.n684 B.n683 10.6151
R2410 B.n683 B.n682 10.6151
R2411 B.n682 B.n121 10.6151
R2412 B.n678 B.n121 10.6151
R2413 B.n678 B.n677 10.6151
R2414 B.n677 B.n676 10.6151
R2415 B.n676 B.n123 10.6151
R2416 B.n672 B.n123 10.6151
R2417 B.n672 B.n671 10.6151
R2418 B.n671 B.n670 10.6151
R2419 B.n670 B.n125 10.6151
R2420 B.n666 B.n125 10.6151
R2421 B.n666 B.n665 10.6151
R2422 B.n665 B.n664 10.6151
R2423 B.n664 B.n127 10.6151
R2424 B.n660 B.n127 10.6151
R2425 B.n660 B.n659 10.6151
R2426 B.n659 B.n658 10.6151
R2427 B.n658 B.n129 10.6151
R2428 B.n654 B.n129 10.6151
R2429 B.n654 B.n653 10.6151
R2430 B.n653 B.n652 10.6151
R2431 B.n652 B.n131 10.6151
R2432 B.n648 B.n131 10.6151
R2433 B.n648 B.n647 10.6151
R2434 B.n647 B.n646 10.6151
R2435 B.n646 B.n133 10.6151
R2436 B.n642 B.n133 10.6151
R2437 B.n642 B.n641 10.6151
R2438 B.n641 B.n640 10.6151
R2439 B.n640 B.n135 10.6151
R2440 B.n636 B.n135 10.6151
R2441 B.n636 B.n635 10.6151
R2442 B.n635 B.n634 10.6151
R2443 B.n634 B.n137 10.6151
R2444 B.n630 B.n137 10.6151
R2445 B.n630 B.n629 10.6151
R2446 B.n629 B.n628 10.6151
R2447 B.n628 B.n139 10.6151
R2448 B.n624 B.n139 10.6151
R2449 B.n624 B.n623 10.6151
R2450 B.n623 B.n622 10.6151
R2451 B.n622 B.n141 10.6151
R2452 B.n618 B.n141 10.6151
R2453 B.n618 B.n617 10.6151
R2454 B.n617 B.n616 10.6151
R2455 B.n616 B.n143 10.6151
R2456 B.n612 B.n143 10.6151
R2457 B.n612 B.n611 10.6151
R2458 B.n611 B.n610 10.6151
R2459 B.n610 B.n145 10.6151
R2460 B.n606 B.n145 10.6151
R2461 B.n606 B.n605 10.6151
R2462 B.n605 B.n604 10.6151
R2463 B.n604 B.n147 10.6151
R2464 B.n600 B.n147 10.6151
R2465 B.n600 B.n599 10.6151
R2466 B.n599 B.n598 10.6151
R2467 B.n598 B.n149 10.6151
R2468 B.n594 B.n149 10.6151
R2469 B.n594 B.n593 10.6151
R2470 B.n593 B.n592 10.6151
R2471 B.n592 B.n151 10.6151
R2472 B.n588 B.n151 10.6151
R2473 B.n588 B.n587 10.6151
R2474 B.n587 B.n586 10.6151
R2475 B.n586 B.n153 10.6151
R2476 B.n582 B.n153 10.6151
R2477 B.n582 B.n581 10.6151
R2478 B.n581 B.n580 10.6151
R2479 B.n580 B.n155 10.6151
R2480 B.n576 B.n155 10.6151
R2481 B.n576 B.n575 10.6151
R2482 B.n575 B.n574 10.6151
R2483 B.n574 B.n157 10.6151
R2484 B.n570 B.n157 10.6151
R2485 B.n570 B.n569 10.6151
R2486 B.n569 B.n568 10.6151
R2487 B.n568 B.n159 10.6151
R2488 B.n564 B.n159 10.6151
R2489 B.n564 B.n563 10.6151
R2490 B.n563 B.n562 10.6151
R2491 B.n562 B.n161 10.6151
R2492 B.n558 B.n161 10.6151
R2493 B.n558 B.n557 10.6151
R2494 B.n557 B.n556 10.6151
R2495 B.n556 B.n163 10.6151
R2496 B.n552 B.n163 10.6151
R2497 B.n552 B.n551 10.6151
R2498 B.n551 B.n550 10.6151
R2499 B.n550 B.n165 10.6151
R2500 B.n546 B.n165 10.6151
R2501 B.n546 B.n545 10.6151
R2502 B.n545 B.n544 10.6151
R2503 B.n544 B.n167 10.6151
R2504 B.n540 B.n167 10.6151
R2505 B.n540 B.n539 10.6151
R2506 B.n539 B.n538 10.6151
R2507 B.n538 B.n169 10.6151
R2508 B.n534 B.n169 10.6151
R2509 B.n534 B.n533 10.6151
R2510 B.n533 B.n532 10.6151
R2511 B.n532 B.n171 10.6151
R2512 B.n528 B.n171 10.6151
R2513 B.n528 B.n527 10.6151
R2514 B.n527 B.n526 10.6151
R2515 B.n526 B.n173 10.6151
R2516 B.n522 B.n173 10.6151
R2517 B.n522 B.n521 10.6151
R2518 B.n521 B.n520 10.6151
R2519 B.n520 B.n175 10.6151
R2520 B.n261 B.n1 10.6151
R2521 B.n264 B.n261 10.6151
R2522 B.n265 B.n264 10.6151
R2523 B.n266 B.n265 10.6151
R2524 B.n266 B.n259 10.6151
R2525 B.n270 B.n259 10.6151
R2526 B.n271 B.n270 10.6151
R2527 B.n272 B.n271 10.6151
R2528 B.n272 B.n257 10.6151
R2529 B.n276 B.n257 10.6151
R2530 B.n277 B.n276 10.6151
R2531 B.n278 B.n277 10.6151
R2532 B.n278 B.n255 10.6151
R2533 B.n282 B.n255 10.6151
R2534 B.n283 B.n282 10.6151
R2535 B.n284 B.n283 10.6151
R2536 B.n284 B.n253 10.6151
R2537 B.n288 B.n253 10.6151
R2538 B.n289 B.n288 10.6151
R2539 B.n290 B.n289 10.6151
R2540 B.n290 B.n251 10.6151
R2541 B.n294 B.n251 10.6151
R2542 B.n295 B.n294 10.6151
R2543 B.n296 B.n295 10.6151
R2544 B.n296 B.n249 10.6151
R2545 B.n300 B.n249 10.6151
R2546 B.n301 B.n300 10.6151
R2547 B.n302 B.n301 10.6151
R2548 B.n302 B.n247 10.6151
R2549 B.n306 B.n247 10.6151
R2550 B.n307 B.n306 10.6151
R2551 B.n308 B.n307 10.6151
R2552 B.n308 B.n245 10.6151
R2553 B.n312 B.n245 10.6151
R2554 B.n313 B.n312 10.6151
R2555 B.n314 B.n313 10.6151
R2556 B.n314 B.n243 10.6151
R2557 B.n318 B.n243 10.6151
R2558 B.n319 B.n318 10.6151
R2559 B.n320 B.n319 10.6151
R2560 B.n320 B.n241 10.6151
R2561 B.n324 B.n241 10.6151
R2562 B.n325 B.n324 10.6151
R2563 B.n326 B.n325 10.6151
R2564 B.n326 B.n239 10.6151
R2565 B.n330 B.n239 10.6151
R2566 B.n331 B.n330 10.6151
R2567 B.n332 B.n331 10.6151
R2568 B.n332 B.n237 10.6151
R2569 B.n336 B.n237 10.6151
R2570 B.n337 B.n336 10.6151
R2571 B.n338 B.n337 10.6151
R2572 B.n338 B.n235 10.6151
R2573 B.n342 B.n235 10.6151
R2574 B.n343 B.n342 10.6151
R2575 B.n344 B.n343 10.6151
R2576 B.n344 B.n233 10.6151
R2577 B.n348 B.n233 10.6151
R2578 B.n349 B.n348 10.6151
R2579 B.n350 B.n349 10.6151
R2580 B.n350 B.n231 10.6151
R2581 B.n354 B.n231 10.6151
R2582 B.n355 B.n354 10.6151
R2583 B.n356 B.n355 10.6151
R2584 B.n356 B.n229 10.6151
R2585 B.n360 B.n229 10.6151
R2586 B.n361 B.n360 10.6151
R2587 B.n362 B.n361 10.6151
R2588 B.n362 B.n227 10.6151
R2589 B.n366 B.n227 10.6151
R2590 B.n367 B.n366 10.6151
R2591 B.n368 B.n367 10.6151
R2592 B.n368 B.n225 10.6151
R2593 B.n372 B.n225 10.6151
R2594 B.n373 B.n372 10.6151
R2595 B.n374 B.n373 10.6151
R2596 B.n374 B.n223 10.6151
R2597 B.n378 B.n223 10.6151
R2598 B.n379 B.n378 10.6151
R2599 B.n380 B.n379 10.6151
R2600 B.n380 B.n221 10.6151
R2601 B.n384 B.n221 10.6151
R2602 B.n386 B.n385 10.6151
R2603 B.n386 B.n219 10.6151
R2604 B.n390 B.n219 10.6151
R2605 B.n391 B.n390 10.6151
R2606 B.n392 B.n391 10.6151
R2607 B.n392 B.n217 10.6151
R2608 B.n396 B.n217 10.6151
R2609 B.n397 B.n396 10.6151
R2610 B.n398 B.n397 10.6151
R2611 B.n398 B.n215 10.6151
R2612 B.n402 B.n215 10.6151
R2613 B.n403 B.n402 10.6151
R2614 B.n404 B.n403 10.6151
R2615 B.n404 B.n213 10.6151
R2616 B.n408 B.n213 10.6151
R2617 B.n409 B.n408 10.6151
R2618 B.n410 B.n409 10.6151
R2619 B.n410 B.n211 10.6151
R2620 B.n414 B.n211 10.6151
R2621 B.n415 B.n414 10.6151
R2622 B.n416 B.n415 10.6151
R2623 B.n416 B.n209 10.6151
R2624 B.n420 B.n209 10.6151
R2625 B.n421 B.n420 10.6151
R2626 B.n422 B.n421 10.6151
R2627 B.n422 B.n207 10.6151
R2628 B.n426 B.n207 10.6151
R2629 B.n427 B.n426 10.6151
R2630 B.n428 B.n427 10.6151
R2631 B.n428 B.n205 10.6151
R2632 B.n432 B.n205 10.6151
R2633 B.n433 B.n432 10.6151
R2634 B.n434 B.n433 10.6151
R2635 B.n434 B.n203 10.6151
R2636 B.n438 B.n203 10.6151
R2637 B.n439 B.n438 10.6151
R2638 B.n443 B.n439 10.6151
R2639 B.n447 B.n201 10.6151
R2640 B.n448 B.n447 10.6151
R2641 B.n449 B.n448 10.6151
R2642 B.n449 B.n199 10.6151
R2643 B.n453 B.n199 10.6151
R2644 B.n454 B.n453 10.6151
R2645 B.n455 B.n454 10.6151
R2646 B.n455 B.n197 10.6151
R2647 B.n459 B.n197 10.6151
R2648 B.n462 B.n461 10.6151
R2649 B.n462 B.n193 10.6151
R2650 B.n466 B.n193 10.6151
R2651 B.n467 B.n466 10.6151
R2652 B.n468 B.n467 10.6151
R2653 B.n468 B.n191 10.6151
R2654 B.n472 B.n191 10.6151
R2655 B.n473 B.n472 10.6151
R2656 B.n474 B.n473 10.6151
R2657 B.n474 B.n189 10.6151
R2658 B.n478 B.n189 10.6151
R2659 B.n479 B.n478 10.6151
R2660 B.n480 B.n479 10.6151
R2661 B.n480 B.n187 10.6151
R2662 B.n484 B.n187 10.6151
R2663 B.n485 B.n484 10.6151
R2664 B.n486 B.n485 10.6151
R2665 B.n486 B.n185 10.6151
R2666 B.n490 B.n185 10.6151
R2667 B.n491 B.n490 10.6151
R2668 B.n492 B.n491 10.6151
R2669 B.n492 B.n183 10.6151
R2670 B.n496 B.n183 10.6151
R2671 B.n497 B.n496 10.6151
R2672 B.n498 B.n497 10.6151
R2673 B.n498 B.n181 10.6151
R2674 B.n502 B.n181 10.6151
R2675 B.n503 B.n502 10.6151
R2676 B.n504 B.n503 10.6151
R2677 B.n504 B.n179 10.6151
R2678 B.n508 B.n179 10.6151
R2679 B.n509 B.n508 10.6151
R2680 B.n510 B.n509 10.6151
R2681 B.n510 B.n177 10.6151
R2682 B.n514 B.n177 10.6151
R2683 B.n515 B.n514 10.6151
R2684 B.n516 B.n515 10.6151
R2685 B.n66 B.n62 9.36635
R2686 B.n827 B.n826 9.36635
R2687 B.n443 B.n442 9.36635
R2688 B.n461 B.n460 9.36635
R2689 B.n1025 B.n0 8.11757
R2690 B.n1025 B.n1 8.11757
R2691 B.n841 B.n66 1.24928
R2692 B.n828 B.n827 1.24928
R2693 B.n442 B.n201 1.24928
R2694 B.n460 B.n459 1.24928
C0 VN w_n6082_n3128# 13.406099f
C1 w_n6082_n3128# B 12.4462f
C2 VDD2 VDD1 3.04095f
C3 VP VDD2 0.752304f
C4 VP VDD1 10.9307f
C5 VDD2 VTAIL 10.712501f
C6 VTAIL VDD1 10.651401f
C7 VN VDD2 10.3378f
C8 VN VDD1 0.156074f
C9 VP VTAIL 11.6227f
C10 VDD2 B 3.06853f
C11 B VDD1 2.89882f
C12 VP VN 10.1467f
C13 VN VTAIL 11.607901f
C14 VP B 2.94845f
C15 B VTAIL 3.93781f
C16 VN B 1.60268f
C17 VDD2 w_n6082_n3128# 3.42108f
C18 w_n6082_n3128# VDD1 3.20841f
C19 VP w_n6082_n3128# 14.2021f
C20 w_n6082_n3128# VTAIL 3.24112f
C21 VDD2 VSUBS 2.65856f
C22 VDD1 VSUBS 2.5031f
C23 VTAIL VSUBS 1.585821f
C24 VN VSUBS 9.912081f
C25 VP VSUBS 5.885824f
C26 B VSUBS 6.913374f
C27 w_n6082_n3128# VSUBS 0.234644p
C28 B.n0 VSUBS 0.008042f
C29 B.n1 VSUBS 0.008042f
C30 B.n2 VSUBS 0.011894f
C31 B.n3 VSUBS 0.009114f
C32 B.n4 VSUBS 0.009114f
C33 B.n5 VSUBS 0.009114f
C34 B.n6 VSUBS 0.009114f
C35 B.n7 VSUBS 0.009114f
C36 B.n8 VSUBS 0.009114f
C37 B.n9 VSUBS 0.009114f
C38 B.n10 VSUBS 0.009114f
C39 B.n11 VSUBS 0.009114f
C40 B.n12 VSUBS 0.009114f
C41 B.n13 VSUBS 0.009114f
C42 B.n14 VSUBS 0.009114f
C43 B.n15 VSUBS 0.009114f
C44 B.n16 VSUBS 0.009114f
C45 B.n17 VSUBS 0.009114f
C46 B.n18 VSUBS 0.009114f
C47 B.n19 VSUBS 0.009114f
C48 B.n20 VSUBS 0.009114f
C49 B.n21 VSUBS 0.009114f
C50 B.n22 VSUBS 0.009114f
C51 B.n23 VSUBS 0.009114f
C52 B.n24 VSUBS 0.009114f
C53 B.n25 VSUBS 0.009114f
C54 B.n26 VSUBS 0.009114f
C55 B.n27 VSUBS 0.009114f
C56 B.n28 VSUBS 0.009114f
C57 B.n29 VSUBS 0.009114f
C58 B.n30 VSUBS 0.009114f
C59 B.n31 VSUBS 0.009114f
C60 B.n32 VSUBS 0.009114f
C61 B.n33 VSUBS 0.009114f
C62 B.n34 VSUBS 0.009114f
C63 B.n35 VSUBS 0.009114f
C64 B.n36 VSUBS 0.009114f
C65 B.n37 VSUBS 0.009114f
C66 B.n38 VSUBS 0.009114f
C67 B.n39 VSUBS 0.009114f
C68 B.n40 VSUBS 0.009114f
C69 B.n41 VSUBS 0.009114f
C70 B.n42 VSUBS 0.009114f
C71 B.n43 VSUBS 0.019213f
C72 B.n44 VSUBS 0.009114f
C73 B.n45 VSUBS 0.009114f
C74 B.n46 VSUBS 0.009114f
C75 B.n47 VSUBS 0.009114f
C76 B.n48 VSUBS 0.009114f
C77 B.n49 VSUBS 0.009114f
C78 B.n50 VSUBS 0.009114f
C79 B.n51 VSUBS 0.009114f
C80 B.n52 VSUBS 0.009114f
C81 B.n53 VSUBS 0.009114f
C82 B.n54 VSUBS 0.009114f
C83 B.n55 VSUBS 0.009114f
C84 B.n56 VSUBS 0.009114f
C85 B.n57 VSUBS 0.009114f
C86 B.n58 VSUBS 0.009114f
C87 B.n59 VSUBS 0.009114f
C88 B.n60 VSUBS 0.009114f
C89 B.n61 VSUBS 0.009114f
C90 B.n62 VSUBS 0.008578f
C91 B.n63 VSUBS 0.009114f
C92 B.t4 VSUBS 0.240639f
C93 B.t5 VSUBS 0.297334f
C94 B.t3 VSUBS 2.59599f
C95 B.n64 VSUBS 0.475247f
C96 B.n65 VSUBS 0.312716f
C97 B.n66 VSUBS 0.021117f
C98 B.n67 VSUBS 0.009114f
C99 B.n68 VSUBS 0.009114f
C100 B.n69 VSUBS 0.009114f
C101 B.n70 VSUBS 0.009114f
C102 B.t1 VSUBS 0.240643f
C103 B.t2 VSUBS 0.297337f
C104 B.t0 VSUBS 2.59599f
C105 B.n71 VSUBS 0.475244f
C106 B.n72 VSUBS 0.312712f
C107 B.n73 VSUBS 0.009114f
C108 B.n74 VSUBS 0.009114f
C109 B.n75 VSUBS 0.009114f
C110 B.n76 VSUBS 0.009114f
C111 B.n77 VSUBS 0.009114f
C112 B.n78 VSUBS 0.009114f
C113 B.n79 VSUBS 0.009114f
C114 B.n80 VSUBS 0.009114f
C115 B.n81 VSUBS 0.009114f
C116 B.n82 VSUBS 0.009114f
C117 B.n83 VSUBS 0.009114f
C118 B.n84 VSUBS 0.009114f
C119 B.n85 VSUBS 0.009114f
C120 B.n86 VSUBS 0.009114f
C121 B.n87 VSUBS 0.009114f
C122 B.n88 VSUBS 0.009114f
C123 B.n89 VSUBS 0.009114f
C124 B.n90 VSUBS 0.009114f
C125 B.n91 VSUBS 0.020194f
C126 B.n92 VSUBS 0.009114f
C127 B.n93 VSUBS 0.009114f
C128 B.n94 VSUBS 0.009114f
C129 B.n95 VSUBS 0.009114f
C130 B.n96 VSUBS 0.009114f
C131 B.n97 VSUBS 0.009114f
C132 B.n98 VSUBS 0.009114f
C133 B.n99 VSUBS 0.009114f
C134 B.n100 VSUBS 0.009114f
C135 B.n101 VSUBS 0.009114f
C136 B.n102 VSUBS 0.009114f
C137 B.n103 VSUBS 0.009114f
C138 B.n104 VSUBS 0.009114f
C139 B.n105 VSUBS 0.009114f
C140 B.n106 VSUBS 0.009114f
C141 B.n107 VSUBS 0.009114f
C142 B.n108 VSUBS 0.009114f
C143 B.n109 VSUBS 0.009114f
C144 B.n110 VSUBS 0.009114f
C145 B.n111 VSUBS 0.009114f
C146 B.n112 VSUBS 0.009114f
C147 B.n113 VSUBS 0.009114f
C148 B.n114 VSUBS 0.009114f
C149 B.n115 VSUBS 0.009114f
C150 B.n116 VSUBS 0.009114f
C151 B.n117 VSUBS 0.009114f
C152 B.n118 VSUBS 0.009114f
C153 B.n119 VSUBS 0.009114f
C154 B.n120 VSUBS 0.009114f
C155 B.n121 VSUBS 0.009114f
C156 B.n122 VSUBS 0.009114f
C157 B.n123 VSUBS 0.009114f
C158 B.n124 VSUBS 0.009114f
C159 B.n125 VSUBS 0.009114f
C160 B.n126 VSUBS 0.009114f
C161 B.n127 VSUBS 0.009114f
C162 B.n128 VSUBS 0.009114f
C163 B.n129 VSUBS 0.009114f
C164 B.n130 VSUBS 0.009114f
C165 B.n131 VSUBS 0.009114f
C166 B.n132 VSUBS 0.009114f
C167 B.n133 VSUBS 0.009114f
C168 B.n134 VSUBS 0.009114f
C169 B.n135 VSUBS 0.009114f
C170 B.n136 VSUBS 0.009114f
C171 B.n137 VSUBS 0.009114f
C172 B.n138 VSUBS 0.009114f
C173 B.n139 VSUBS 0.009114f
C174 B.n140 VSUBS 0.009114f
C175 B.n141 VSUBS 0.009114f
C176 B.n142 VSUBS 0.009114f
C177 B.n143 VSUBS 0.009114f
C178 B.n144 VSUBS 0.009114f
C179 B.n145 VSUBS 0.009114f
C180 B.n146 VSUBS 0.009114f
C181 B.n147 VSUBS 0.009114f
C182 B.n148 VSUBS 0.009114f
C183 B.n149 VSUBS 0.009114f
C184 B.n150 VSUBS 0.009114f
C185 B.n151 VSUBS 0.009114f
C186 B.n152 VSUBS 0.009114f
C187 B.n153 VSUBS 0.009114f
C188 B.n154 VSUBS 0.009114f
C189 B.n155 VSUBS 0.009114f
C190 B.n156 VSUBS 0.009114f
C191 B.n157 VSUBS 0.009114f
C192 B.n158 VSUBS 0.009114f
C193 B.n159 VSUBS 0.009114f
C194 B.n160 VSUBS 0.009114f
C195 B.n161 VSUBS 0.009114f
C196 B.n162 VSUBS 0.009114f
C197 B.n163 VSUBS 0.009114f
C198 B.n164 VSUBS 0.009114f
C199 B.n165 VSUBS 0.009114f
C200 B.n166 VSUBS 0.009114f
C201 B.n167 VSUBS 0.009114f
C202 B.n168 VSUBS 0.009114f
C203 B.n169 VSUBS 0.009114f
C204 B.n170 VSUBS 0.009114f
C205 B.n171 VSUBS 0.009114f
C206 B.n172 VSUBS 0.009114f
C207 B.n173 VSUBS 0.009114f
C208 B.n174 VSUBS 0.009114f
C209 B.n175 VSUBS 0.020431f
C210 B.n176 VSUBS 0.009114f
C211 B.n177 VSUBS 0.009114f
C212 B.n178 VSUBS 0.009114f
C213 B.n179 VSUBS 0.009114f
C214 B.n180 VSUBS 0.009114f
C215 B.n181 VSUBS 0.009114f
C216 B.n182 VSUBS 0.009114f
C217 B.n183 VSUBS 0.009114f
C218 B.n184 VSUBS 0.009114f
C219 B.n185 VSUBS 0.009114f
C220 B.n186 VSUBS 0.009114f
C221 B.n187 VSUBS 0.009114f
C222 B.n188 VSUBS 0.009114f
C223 B.n189 VSUBS 0.009114f
C224 B.n190 VSUBS 0.009114f
C225 B.n191 VSUBS 0.009114f
C226 B.n192 VSUBS 0.009114f
C227 B.n193 VSUBS 0.009114f
C228 B.n194 VSUBS 0.009114f
C229 B.t8 VSUBS 0.240643f
C230 B.t7 VSUBS 0.297337f
C231 B.t6 VSUBS 2.59599f
C232 B.n195 VSUBS 0.475244f
C233 B.n196 VSUBS 0.312712f
C234 B.n197 VSUBS 0.009114f
C235 B.n198 VSUBS 0.009114f
C236 B.n199 VSUBS 0.009114f
C237 B.n200 VSUBS 0.009114f
C238 B.n201 VSUBS 0.005093f
C239 B.n202 VSUBS 0.009114f
C240 B.n203 VSUBS 0.009114f
C241 B.n204 VSUBS 0.009114f
C242 B.n205 VSUBS 0.009114f
C243 B.n206 VSUBS 0.009114f
C244 B.n207 VSUBS 0.009114f
C245 B.n208 VSUBS 0.009114f
C246 B.n209 VSUBS 0.009114f
C247 B.n210 VSUBS 0.009114f
C248 B.n211 VSUBS 0.009114f
C249 B.n212 VSUBS 0.009114f
C250 B.n213 VSUBS 0.009114f
C251 B.n214 VSUBS 0.009114f
C252 B.n215 VSUBS 0.009114f
C253 B.n216 VSUBS 0.009114f
C254 B.n217 VSUBS 0.009114f
C255 B.n218 VSUBS 0.009114f
C256 B.n219 VSUBS 0.009114f
C257 B.n220 VSUBS 0.020194f
C258 B.n221 VSUBS 0.009114f
C259 B.n222 VSUBS 0.009114f
C260 B.n223 VSUBS 0.009114f
C261 B.n224 VSUBS 0.009114f
C262 B.n225 VSUBS 0.009114f
C263 B.n226 VSUBS 0.009114f
C264 B.n227 VSUBS 0.009114f
C265 B.n228 VSUBS 0.009114f
C266 B.n229 VSUBS 0.009114f
C267 B.n230 VSUBS 0.009114f
C268 B.n231 VSUBS 0.009114f
C269 B.n232 VSUBS 0.009114f
C270 B.n233 VSUBS 0.009114f
C271 B.n234 VSUBS 0.009114f
C272 B.n235 VSUBS 0.009114f
C273 B.n236 VSUBS 0.009114f
C274 B.n237 VSUBS 0.009114f
C275 B.n238 VSUBS 0.009114f
C276 B.n239 VSUBS 0.009114f
C277 B.n240 VSUBS 0.009114f
C278 B.n241 VSUBS 0.009114f
C279 B.n242 VSUBS 0.009114f
C280 B.n243 VSUBS 0.009114f
C281 B.n244 VSUBS 0.009114f
C282 B.n245 VSUBS 0.009114f
C283 B.n246 VSUBS 0.009114f
C284 B.n247 VSUBS 0.009114f
C285 B.n248 VSUBS 0.009114f
C286 B.n249 VSUBS 0.009114f
C287 B.n250 VSUBS 0.009114f
C288 B.n251 VSUBS 0.009114f
C289 B.n252 VSUBS 0.009114f
C290 B.n253 VSUBS 0.009114f
C291 B.n254 VSUBS 0.009114f
C292 B.n255 VSUBS 0.009114f
C293 B.n256 VSUBS 0.009114f
C294 B.n257 VSUBS 0.009114f
C295 B.n258 VSUBS 0.009114f
C296 B.n259 VSUBS 0.009114f
C297 B.n260 VSUBS 0.009114f
C298 B.n261 VSUBS 0.009114f
C299 B.n262 VSUBS 0.009114f
C300 B.n263 VSUBS 0.009114f
C301 B.n264 VSUBS 0.009114f
C302 B.n265 VSUBS 0.009114f
C303 B.n266 VSUBS 0.009114f
C304 B.n267 VSUBS 0.009114f
C305 B.n268 VSUBS 0.009114f
C306 B.n269 VSUBS 0.009114f
C307 B.n270 VSUBS 0.009114f
C308 B.n271 VSUBS 0.009114f
C309 B.n272 VSUBS 0.009114f
C310 B.n273 VSUBS 0.009114f
C311 B.n274 VSUBS 0.009114f
C312 B.n275 VSUBS 0.009114f
C313 B.n276 VSUBS 0.009114f
C314 B.n277 VSUBS 0.009114f
C315 B.n278 VSUBS 0.009114f
C316 B.n279 VSUBS 0.009114f
C317 B.n280 VSUBS 0.009114f
C318 B.n281 VSUBS 0.009114f
C319 B.n282 VSUBS 0.009114f
C320 B.n283 VSUBS 0.009114f
C321 B.n284 VSUBS 0.009114f
C322 B.n285 VSUBS 0.009114f
C323 B.n286 VSUBS 0.009114f
C324 B.n287 VSUBS 0.009114f
C325 B.n288 VSUBS 0.009114f
C326 B.n289 VSUBS 0.009114f
C327 B.n290 VSUBS 0.009114f
C328 B.n291 VSUBS 0.009114f
C329 B.n292 VSUBS 0.009114f
C330 B.n293 VSUBS 0.009114f
C331 B.n294 VSUBS 0.009114f
C332 B.n295 VSUBS 0.009114f
C333 B.n296 VSUBS 0.009114f
C334 B.n297 VSUBS 0.009114f
C335 B.n298 VSUBS 0.009114f
C336 B.n299 VSUBS 0.009114f
C337 B.n300 VSUBS 0.009114f
C338 B.n301 VSUBS 0.009114f
C339 B.n302 VSUBS 0.009114f
C340 B.n303 VSUBS 0.009114f
C341 B.n304 VSUBS 0.009114f
C342 B.n305 VSUBS 0.009114f
C343 B.n306 VSUBS 0.009114f
C344 B.n307 VSUBS 0.009114f
C345 B.n308 VSUBS 0.009114f
C346 B.n309 VSUBS 0.009114f
C347 B.n310 VSUBS 0.009114f
C348 B.n311 VSUBS 0.009114f
C349 B.n312 VSUBS 0.009114f
C350 B.n313 VSUBS 0.009114f
C351 B.n314 VSUBS 0.009114f
C352 B.n315 VSUBS 0.009114f
C353 B.n316 VSUBS 0.009114f
C354 B.n317 VSUBS 0.009114f
C355 B.n318 VSUBS 0.009114f
C356 B.n319 VSUBS 0.009114f
C357 B.n320 VSUBS 0.009114f
C358 B.n321 VSUBS 0.009114f
C359 B.n322 VSUBS 0.009114f
C360 B.n323 VSUBS 0.009114f
C361 B.n324 VSUBS 0.009114f
C362 B.n325 VSUBS 0.009114f
C363 B.n326 VSUBS 0.009114f
C364 B.n327 VSUBS 0.009114f
C365 B.n328 VSUBS 0.009114f
C366 B.n329 VSUBS 0.009114f
C367 B.n330 VSUBS 0.009114f
C368 B.n331 VSUBS 0.009114f
C369 B.n332 VSUBS 0.009114f
C370 B.n333 VSUBS 0.009114f
C371 B.n334 VSUBS 0.009114f
C372 B.n335 VSUBS 0.009114f
C373 B.n336 VSUBS 0.009114f
C374 B.n337 VSUBS 0.009114f
C375 B.n338 VSUBS 0.009114f
C376 B.n339 VSUBS 0.009114f
C377 B.n340 VSUBS 0.009114f
C378 B.n341 VSUBS 0.009114f
C379 B.n342 VSUBS 0.009114f
C380 B.n343 VSUBS 0.009114f
C381 B.n344 VSUBS 0.009114f
C382 B.n345 VSUBS 0.009114f
C383 B.n346 VSUBS 0.009114f
C384 B.n347 VSUBS 0.009114f
C385 B.n348 VSUBS 0.009114f
C386 B.n349 VSUBS 0.009114f
C387 B.n350 VSUBS 0.009114f
C388 B.n351 VSUBS 0.009114f
C389 B.n352 VSUBS 0.009114f
C390 B.n353 VSUBS 0.009114f
C391 B.n354 VSUBS 0.009114f
C392 B.n355 VSUBS 0.009114f
C393 B.n356 VSUBS 0.009114f
C394 B.n357 VSUBS 0.009114f
C395 B.n358 VSUBS 0.009114f
C396 B.n359 VSUBS 0.009114f
C397 B.n360 VSUBS 0.009114f
C398 B.n361 VSUBS 0.009114f
C399 B.n362 VSUBS 0.009114f
C400 B.n363 VSUBS 0.009114f
C401 B.n364 VSUBS 0.009114f
C402 B.n365 VSUBS 0.009114f
C403 B.n366 VSUBS 0.009114f
C404 B.n367 VSUBS 0.009114f
C405 B.n368 VSUBS 0.009114f
C406 B.n369 VSUBS 0.009114f
C407 B.n370 VSUBS 0.009114f
C408 B.n371 VSUBS 0.009114f
C409 B.n372 VSUBS 0.009114f
C410 B.n373 VSUBS 0.009114f
C411 B.n374 VSUBS 0.009114f
C412 B.n375 VSUBS 0.009114f
C413 B.n376 VSUBS 0.009114f
C414 B.n377 VSUBS 0.009114f
C415 B.n378 VSUBS 0.009114f
C416 B.n379 VSUBS 0.009114f
C417 B.n380 VSUBS 0.009114f
C418 B.n381 VSUBS 0.009114f
C419 B.n382 VSUBS 0.009114f
C420 B.n383 VSUBS 0.019213f
C421 B.n384 VSUBS 0.019213f
C422 B.n385 VSUBS 0.020194f
C423 B.n386 VSUBS 0.009114f
C424 B.n387 VSUBS 0.009114f
C425 B.n388 VSUBS 0.009114f
C426 B.n389 VSUBS 0.009114f
C427 B.n390 VSUBS 0.009114f
C428 B.n391 VSUBS 0.009114f
C429 B.n392 VSUBS 0.009114f
C430 B.n393 VSUBS 0.009114f
C431 B.n394 VSUBS 0.009114f
C432 B.n395 VSUBS 0.009114f
C433 B.n396 VSUBS 0.009114f
C434 B.n397 VSUBS 0.009114f
C435 B.n398 VSUBS 0.009114f
C436 B.n399 VSUBS 0.009114f
C437 B.n400 VSUBS 0.009114f
C438 B.n401 VSUBS 0.009114f
C439 B.n402 VSUBS 0.009114f
C440 B.n403 VSUBS 0.009114f
C441 B.n404 VSUBS 0.009114f
C442 B.n405 VSUBS 0.009114f
C443 B.n406 VSUBS 0.009114f
C444 B.n407 VSUBS 0.009114f
C445 B.n408 VSUBS 0.009114f
C446 B.n409 VSUBS 0.009114f
C447 B.n410 VSUBS 0.009114f
C448 B.n411 VSUBS 0.009114f
C449 B.n412 VSUBS 0.009114f
C450 B.n413 VSUBS 0.009114f
C451 B.n414 VSUBS 0.009114f
C452 B.n415 VSUBS 0.009114f
C453 B.n416 VSUBS 0.009114f
C454 B.n417 VSUBS 0.009114f
C455 B.n418 VSUBS 0.009114f
C456 B.n419 VSUBS 0.009114f
C457 B.n420 VSUBS 0.009114f
C458 B.n421 VSUBS 0.009114f
C459 B.n422 VSUBS 0.009114f
C460 B.n423 VSUBS 0.009114f
C461 B.n424 VSUBS 0.009114f
C462 B.n425 VSUBS 0.009114f
C463 B.n426 VSUBS 0.009114f
C464 B.n427 VSUBS 0.009114f
C465 B.n428 VSUBS 0.009114f
C466 B.n429 VSUBS 0.009114f
C467 B.n430 VSUBS 0.009114f
C468 B.n431 VSUBS 0.009114f
C469 B.n432 VSUBS 0.009114f
C470 B.n433 VSUBS 0.009114f
C471 B.n434 VSUBS 0.009114f
C472 B.n435 VSUBS 0.009114f
C473 B.n436 VSUBS 0.009114f
C474 B.n437 VSUBS 0.009114f
C475 B.n438 VSUBS 0.009114f
C476 B.n439 VSUBS 0.009114f
C477 B.t11 VSUBS 0.240639f
C478 B.t10 VSUBS 0.297334f
C479 B.t9 VSUBS 2.59599f
C480 B.n440 VSUBS 0.475247f
C481 B.n441 VSUBS 0.312716f
C482 B.n442 VSUBS 0.021117f
C483 B.n443 VSUBS 0.008578f
C484 B.n444 VSUBS 0.009114f
C485 B.n445 VSUBS 0.009114f
C486 B.n446 VSUBS 0.009114f
C487 B.n447 VSUBS 0.009114f
C488 B.n448 VSUBS 0.009114f
C489 B.n449 VSUBS 0.009114f
C490 B.n450 VSUBS 0.009114f
C491 B.n451 VSUBS 0.009114f
C492 B.n452 VSUBS 0.009114f
C493 B.n453 VSUBS 0.009114f
C494 B.n454 VSUBS 0.009114f
C495 B.n455 VSUBS 0.009114f
C496 B.n456 VSUBS 0.009114f
C497 B.n457 VSUBS 0.009114f
C498 B.n458 VSUBS 0.009114f
C499 B.n459 VSUBS 0.005093f
C500 B.n460 VSUBS 0.021117f
C501 B.n461 VSUBS 0.008578f
C502 B.n462 VSUBS 0.009114f
C503 B.n463 VSUBS 0.009114f
C504 B.n464 VSUBS 0.009114f
C505 B.n465 VSUBS 0.009114f
C506 B.n466 VSUBS 0.009114f
C507 B.n467 VSUBS 0.009114f
C508 B.n468 VSUBS 0.009114f
C509 B.n469 VSUBS 0.009114f
C510 B.n470 VSUBS 0.009114f
C511 B.n471 VSUBS 0.009114f
C512 B.n472 VSUBS 0.009114f
C513 B.n473 VSUBS 0.009114f
C514 B.n474 VSUBS 0.009114f
C515 B.n475 VSUBS 0.009114f
C516 B.n476 VSUBS 0.009114f
C517 B.n477 VSUBS 0.009114f
C518 B.n478 VSUBS 0.009114f
C519 B.n479 VSUBS 0.009114f
C520 B.n480 VSUBS 0.009114f
C521 B.n481 VSUBS 0.009114f
C522 B.n482 VSUBS 0.009114f
C523 B.n483 VSUBS 0.009114f
C524 B.n484 VSUBS 0.009114f
C525 B.n485 VSUBS 0.009114f
C526 B.n486 VSUBS 0.009114f
C527 B.n487 VSUBS 0.009114f
C528 B.n488 VSUBS 0.009114f
C529 B.n489 VSUBS 0.009114f
C530 B.n490 VSUBS 0.009114f
C531 B.n491 VSUBS 0.009114f
C532 B.n492 VSUBS 0.009114f
C533 B.n493 VSUBS 0.009114f
C534 B.n494 VSUBS 0.009114f
C535 B.n495 VSUBS 0.009114f
C536 B.n496 VSUBS 0.009114f
C537 B.n497 VSUBS 0.009114f
C538 B.n498 VSUBS 0.009114f
C539 B.n499 VSUBS 0.009114f
C540 B.n500 VSUBS 0.009114f
C541 B.n501 VSUBS 0.009114f
C542 B.n502 VSUBS 0.009114f
C543 B.n503 VSUBS 0.009114f
C544 B.n504 VSUBS 0.009114f
C545 B.n505 VSUBS 0.009114f
C546 B.n506 VSUBS 0.009114f
C547 B.n507 VSUBS 0.009114f
C548 B.n508 VSUBS 0.009114f
C549 B.n509 VSUBS 0.009114f
C550 B.n510 VSUBS 0.009114f
C551 B.n511 VSUBS 0.009114f
C552 B.n512 VSUBS 0.009114f
C553 B.n513 VSUBS 0.009114f
C554 B.n514 VSUBS 0.009114f
C555 B.n515 VSUBS 0.009114f
C556 B.n516 VSUBS 0.018976f
C557 B.n517 VSUBS 0.020194f
C558 B.n518 VSUBS 0.019213f
C559 B.n519 VSUBS 0.009114f
C560 B.n520 VSUBS 0.009114f
C561 B.n521 VSUBS 0.009114f
C562 B.n522 VSUBS 0.009114f
C563 B.n523 VSUBS 0.009114f
C564 B.n524 VSUBS 0.009114f
C565 B.n525 VSUBS 0.009114f
C566 B.n526 VSUBS 0.009114f
C567 B.n527 VSUBS 0.009114f
C568 B.n528 VSUBS 0.009114f
C569 B.n529 VSUBS 0.009114f
C570 B.n530 VSUBS 0.009114f
C571 B.n531 VSUBS 0.009114f
C572 B.n532 VSUBS 0.009114f
C573 B.n533 VSUBS 0.009114f
C574 B.n534 VSUBS 0.009114f
C575 B.n535 VSUBS 0.009114f
C576 B.n536 VSUBS 0.009114f
C577 B.n537 VSUBS 0.009114f
C578 B.n538 VSUBS 0.009114f
C579 B.n539 VSUBS 0.009114f
C580 B.n540 VSUBS 0.009114f
C581 B.n541 VSUBS 0.009114f
C582 B.n542 VSUBS 0.009114f
C583 B.n543 VSUBS 0.009114f
C584 B.n544 VSUBS 0.009114f
C585 B.n545 VSUBS 0.009114f
C586 B.n546 VSUBS 0.009114f
C587 B.n547 VSUBS 0.009114f
C588 B.n548 VSUBS 0.009114f
C589 B.n549 VSUBS 0.009114f
C590 B.n550 VSUBS 0.009114f
C591 B.n551 VSUBS 0.009114f
C592 B.n552 VSUBS 0.009114f
C593 B.n553 VSUBS 0.009114f
C594 B.n554 VSUBS 0.009114f
C595 B.n555 VSUBS 0.009114f
C596 B.n556 VSUBS 0.009114f
C597 B.n557 VSUBS 0.009114f
C598 B.n558 VSUBS 0.009114f
C599 B.n559 VSUBS 0.009114f
C600 B.n560 VSUBS 0.009114f
C601 B.n561 VSUBS 0.009114f
C602 B.n562 VSUBS 0.009114f
C603 B.n563 VSUBS 0.009114f
C604 B.n564 VSUBS 0.009114f
C605 B.n565 VSUBS 0.009114f
C606 B.n566 VSUBS 0.009114f
C607 B.n567 VSUBS 0.009114f
C608 B.n568 VSUBS 0.009114f
C609 B.n569 VSUBS 0.009114f
C610 B.n570 VSUBS 0.009114f
C611 B.n571 VSUBS 0.009114f
C612 B.n572 VSUBS 0.009114f
C613 B.n573 VSUBS 0.009114f
C614 B.n574 VSUBS 0.009114f
C615 B.n575 VSUBS 0.009114f
C616 B.n576 VSUBS 0.009114f
C617 B.n577 VSUBS 0.009114f
C618 B.n578 VSUBS 0.009114f
C619 B.n579 VSUBS 0.009114f
C620 B.n580 VSUBS 0.009114f
C621 B.n581 VSUBS 0.009114f
C622 B.n582 VSUBS 0.009114f
C623 B.n583 VSUBS 0.009114f
C624 B.n584 VSUBS 0.009114f
C625 B.n585 VSUBS 0.009114f
C626 B.n586 VSUBS 0.009114f
C627 B.n587 VSUBS 0.009114f
C628 B.n588 VSUBS 0.009114f
C629 B.n589 VSUBS 0.009114f
C630 B.n590 VSUBS 0.009114f
C631 B.n591 VSUBS 0.009114f
C632 B.n592 VSUBS 0.009114f
C633 B.n593 VSUBS 0.009114f
C634 B.n594 VSUBS 0.009114f
C635 B.n595 VSUBS 0.009114f
C636 B.n596 VSUBS 0.009114f
C637 B.n597 VSUBS 0.009114f
C638 B.n598 VSUBS 0.009114f
C639 B.n599 VSUBS 0.009114f
C640 B.n600 VSUBS 0.009114f
C641 B.n601 VSUBS 0.009114f
C642 B.n602 VSUBS 0.009114f
C643 B.n603 VSUBS 0.009114f
C644 B.n604 VSUBS 0.009114f
C645 B.n605 VSUBS 0.009114f
C646 B.n606 VSUBS 0.009114f
C647 B.n607 VSUBS 0.009114f
C648 B.n608 VSUBS 0.009114f
C649 B.n609 VSUBS 0.009114f
C650 B.n610 VSUBS 0.009114f
C651 B.n611 VSUBS 0.009114f
C652 B.n612 VSUBS 0.009114f
C653 B.n613 VSUBS 0.009114f
C654 B.n614 VSUBS 0.009114f
C655 B.n615 VSUBS 0.009114f
C656 B.n616 VSUBS 0.009114f
C657 B.n617 VSUBS 0.009114f
C658 B.n618 VSUBS 0.009114f
C659 B.n619 VSUBS 0.009114f
C660 B.n620 VSUBS 0.009114f
C661 B.n621 VSUBS 0.009114f
C662 B.n622 VSUBS 0.009114f
C663 B.n623 VSUBS 0.009114f
C664 B.n624 VSUBS 0.009114f
C665 B.n625 VSUBS 0.009114f
C666 B.n626 VSUBS 0.009114f
C667 B.n627 VSUBS 0.009114f
C668 B.n628 VSUBS 0.009114f
C669 B.n629 VSUBS 0.009114f
C670 B.n630 VSUBS 0.009114f
C671 B.n631 VSUBS 0.009114f
C672 B.n632 VSUBS 0.009114f
C673 B.n633 VSUBS 0.009114f
C674 B.n634 VSUBS 0.009114f
C675 B.n635 VSUBS 0.009114f
C676 B.n636 VSUBS 0.009114f
C677 B.n637 VSUBS 0.009114f
C678 B.n638 VSUBS 0.009114f
C679 B.n639 VSUBS 0.009114f
C680 B.n640 VSUBS 0.009114f
C681 B.n641 VSUBS 0.009114f
C682 B.n642 VSUBS 0.009114f
C683 B.n643 VSUBS 0.009114f
C684 B.n644 VSUBS 0.009114f
C685 B.n645 VSUBS 0.009114f
C686 B.n646 VSUBS 0.009114f
C687 B.n647 VSUBS 0.009114f
C688 B.n648 VSUBS 0.009114f
C689 B.n649 VSUBS 0.009114f
C690 B.n650 VSUBS 0.009114f
C691 B.n651 VSUBS 0.009114f
C692 B.n652 VSUBS 0.009114f
C693 B.n653 VSUBS 0.009114f
C694 B.n654 VSUBS 0.009114f
C695 B.n655 VSUBS 0.009114f
C696 B.n656 VSUBS 0.009114f
C697 B.n657 VSUBS 0.009114f
C698 B.n658 VSUBS 0.009114f
C699 B.n659 VSUBS 0.009114f
C700 B.n660 VSUBS 0.009114f
C701 B.n661 VSUBS 0.009114f
C702 B.n662 VSUBS 0.009114f
C703 B.n663 VSUBS 0.009114f
C704 B.n664 VSUBS 0.009114f
C705 B.n665 VSUBS 0.009114f
C706 B.n666 VSUBS 0.009114f
C707 B.n667 VSUBS 0.009114f
C708 B.n668 VSUBS 0.009114f
C709 B.n669 VSUBS 0.009114f
C710 B.n670 VSUBS 0.009114f
C711 B.n671 VSUBS 0.009114f
C712 B.n672 VSUBS 0.009114f
C713 B.n673 VSUBS 0.009114f
C714 B.n674 VSUBS 0.009114f
C715 B.n675 VSUBS 0.009114f
C716 B.n676 VSUBS 0.009114f
C717 B.n677 VSUBS 0.009114f
C718 B.n678 VSUBS 0.009114f
C719 B.n679 VSUBS 0.009114f
C720 B.n680 VSUBS 0.009114f
C721 B.n681 VSUBS 0.009114f
C722 B.n682 VSUBS 0.009114f
C723 B.n683 VSUBS 0.009114f
C724 B.n684 VSUBS 0.009114f
C725 B.n685 VSUBS 0.009114f
C726 B.n686 VSUBS 0.009114f
C727 B.n687 VSUBS 0.009114f
C728 B.n688 VSUBS 0.009114f
C729 B.n689 VSUBS 0.009114f
C730 B.n690 VSUBS 0.009114f
C731 B.n691 VSUBS 0.009114f
C732 B.n692 VSUBS 0.009114f
C733 B.n693 VSUBS 0.009114f
C734 B.n694 VSUBS 0.009114f
C735 B.n695 VSUBS 0.009114f
C736 B.n696 VSUBS 0.009114f
C737 B.n697 VSUBS 0.009114f
C738 B.n698 VSUBS 0.009114f
C739 B.n699 VSUBS 0.009114f
C740 B.n700 VSUBS 0.009114f
C741 B.n701 VSUBS 0.009114f
C742 B.n702 VSUBS 0.009114f
C743 B.n703 VSUBS 0.009114f
C744 B.n704 VSUBS 0.009114f
C745 B.n705 VSUBS 0.009114f
C746 B.n706 VSUBS 0.009114f
C747 B.n707 VSUBS 0.009114f
C748 B.n708 VSUBS 0.009114f
C749 B.n709 VSUBS 0.009114f
C750 B.n710 VSUBS 0.009114f
C751 B.n711 VSUBS 0.009114f
C752 B.n712 VSUBS 0.009114f
C753 B.n713 VSUBS 0.009114f
C754 B.n714 VSUBS 0.009114f
C755 B.n715 VSUBS 0.009114f
C756 B.n716 VSUBS 0.009114f
C757 B.n717 VSUBS 0.009114f
C758 B.n718 VSUBS 0.009114f
C759 B.n719 VSUBS 0.009114f
C760 B.n720 VSUBS 0.009114f
C761 B.n721 VSUBS 0.009114f
C762 B.n722 VSUBS 0.009114f
C763 B.n723 VSUBS 0.009114f
C764 B.n724 VSUBS 0.009114f
C765 B.n725 VSUBS 0.009114f
C766 B.n726 VSUBS 0.009114f
C767 B.n727 VSUBS 0.009114f
C768 B.n728 VSUBS 0.009114f
C769 B.n729 VSUBS 0.009114f
C770 B.n730 VSUBS 0.009114f
C771 B.n731 VSUBS 0.009114f
C772 B.n732 VSUBS 0.009114f
C773 B.n733 VSUBS 0.009114f
C774 B.n734 VSUBS 0.009114f
C775 B.n735 VSUBS 0.009114f
C776 B.n736 VSUBS 0.009114f
C777 B.n737 VSUBS 0.009114f
C778 B.n738 VSUBS 0.009114f
C779 B.n739 VSUBS 0.009114f
C780 B.n740 VSUBS 0.009114f
C781 B.n741 VSUBS 0.009114f
C782 B.n742 VSUBS 0.009114f
C783 B.n743 VSUBS 0.009114f
C784 B.n744 VSUBS 0.009114f
C785 B.n745 VSUBS 0.009114f
C786 B.n746 VSUBS 0.009114f
C787 B.n747 VSUBS 0.009114f
C788 B.n748 VSUBS 0.009114f
C789 B.n749 VSUBS 0.009114f
C790 B.n750 VSUBS 0.009114f
C791 B.n751 VSUBS 0.009114f
C792 B.n752 VSUBS 0.009114f
C793 B.n753 VSUBS 0.009114f
C794 B.n754 VSUBS 0.009114f
C795 B.n755 VSUBS 0.009114f
C796 B.n756 VSUBS 0.009114f
C797 B.n757 VSUBS 0.009114f
C798 B.n758 VSUBS 0.009114f
C799 B.n759 VSUBS 0.009114f
C800 B.n760 VSUBS 0.009114f
C801 B.n761 VSUBS 0.009114f
C802 B.n762 VSUBS 0.009114f
C803 B.n763 VSUBS 0.009114f
C804 B.n764 VSUBS 0.009114f
C805 B.n765 VSUBS 0.009114f
C806 B.n766 VSUBS 0.009114f
C807 B.n767 VSUBS 0.009114f
C808 B.n768 VSUBS 0.019213f
C809 B.n769 VSUBS 0.019213f
C810 B.n770 VSUBS 0.020194f
C811 B.n771 VSUBS 0.009114f
C812 B.n772 VSUBS 0.009114f
C813 B.n773 VSUBS 0.009114f
C814 B.n774 VSUBS 0.009114f
C815 B.n775 VSUBS 0.009114f
C816 B.n776 VSUBS 0.009114f
C817 B.n777 VSUBS 0.009114f
C818 B.n778 VSUBS 0.009114f
C819 B.n779 VSUBS 0.009114f
C820 B.n780 VSUBS 0.009114f
C821 B.n781 VSUBS 0.009114f
C822 B.n782 VSUBS 0.009114f
C823 B.n783 VSUBS 0.009114f
C824 B.n784 VSUBS 0.009114f
C825 B.n785 VSUBS 0.009114f
C826 B.n786 VSUBS 0.009114f
C827 B.n787 VSUBS 0.009114f
C828 B.n788 VSUBS 0.009114f
C829 B.n789 VSUBS 0.009114f
C830 B.n790 VSUBS 0.009114f
C831 B.n791 VSUBS 0.009114f
C832 B.n792 VSUBS 0.009114f
C833 B.n793 VSUBS 0.009114f
C834 B.n794 VSUBS 0.009114f
C835 B.n795 VSUBS 0.009114f
C836 B.n796 VSUBS 0.009114f
C837 B.n797 VSUBS 0.009114f
C838 B.n798 VSUBS 0.009114f
C839 B.n799 VSUBS 0.009114f
C840 B.n800 VSUBS 0.009114f
C841 B.n801 VSUBS 0.009114f
C842 B.n802 VSUBS 0.009114f
C843 B.n803 VSUBS 0.009114f
C844 B.n804 VSUBS 0.009114f
C845 B.n805 VSUBS 0.009114f
C846 B.n806 VSUBS 0.009114f
C847 B.n807 VSUBS 0.009114f
C848 B.n808 VSUBS 0.009114f
C849 B.n809 VSUBS 0.009114f
C850 B.n810 VSUBS 0.009114f
C851 B.n811 VSUBS 0.009114f
C852 B.n812 VSUBS 0.009114f
C853 B.n813 VSUBS 0.009114f
C854 B.n814 VSUBS 0.009114f
C855 B.n815 VSUBS 0.009114f
C856 B.n816 VSUBS 0.009114f
C857 B.n817 VSUBS 0.009114f
C858 B.n818 VSUBS 0.009114f
C859 B.n819 VSUBS 0.009114f
C860 B.n820 VSUBS 0.009114f
C861 B.n821 VSUBS 0.009114f
C862 B.n822 VSUBS 0.009114f
C863 B.n823 VSUBS 0.009114f
C864 B.n824 VSUBS 0.009114f
C865 B.n825 VSUBS 0.009114f
C866 B.n826 VSUBS 0.008578f
C867 B.n827 VSUBS 0.021117f
C868 B.n828 VSUBS 0.005093f
C869 B.n829 VSUBS 0.009114f
C870 B.n830 VSUBS 0.009114f
C871 B.n831 VSUBS 0.009114f
C872 B.n832 VSUBS 0.009114f
C873 B.n833 VSUBS 0.009114f
C874 B.n834 VSUBS 0.009114f
C875 B.n835 VSUBS 0.009114f
C876 B.n836 VSUBS 0.009114f
C877 B.n837 VSUBS 0.009114f
C878 B.n838 VSUBS 0.009114f
C879 B.n839 VSUBS 0.009114f
C880 B.n840 VSUBS 0.009114f
C881 B.n841 VSUBS 0.005093f
C882 B.n842 VSUBS 0.009114f
C883 B.n843 VSUBS 0.009114f
C884 B.n844 VSUBS 0.009114f
C885 B.n845 VSUBS 0.009114f
C886 B.n846 VSUBS 0.009114f
C887 B.n847 VSUBS 0.009114f
C888 B.n848 VSUBS 0.009114f
C889 B.n849 VSUBS 0.009114f
C890 B.n850 VSUBS 0.009114f
C891 B.n851 VSUBS 0.009114f
C892 B.n852 VSUBS 0.009114f
C893 B.n853 VSUBS 0.009114f
C894 B.n854 VSUBS 0.009114f
C895 B.n855 VSUBS 0.009114f
C896 B.n856 VSUBS 0.009114f
C897 B.n857 VSUBS 0.009114f
C898 B.n858 VSUBS 0.009114f
C899 B.n859 VSUBS 0.009114f
C900 B.n860 VSUBS 0.009114f
C901 B.n861 VSUBS 0.009114f
C902 B.n862 VSUBS 0.009114f
C903 B.n863 VSUBS 0.009114f
C904 B.n864 VSUBS 0.009114f
C905 B.n865 VSUBS 0.009114f
C906 B.n866 VSUBS 0.009114f
C907 B.n867 VSUBS 0.009114f
C908 B.n868 VSUBS 0.009114f
C909 B.n869 VSUBS 0.009114f
C910 B.n870 VSUBS 0.009114f
C911 B.n871 VSUBS 0.009114f
C912 B.n872 VSUBS 0.009114f
C913 B.n873 VSUBS 0.009114f
C914 B.n874 VSUBS 0.009114f
C915 B.n875 VSUBS 0.009114f
C916 B.n876 VSUBS 0.009114f
C917 B.n877 VSUBS 0.009114f
C918 B.n878 VSUBS 0.009114f
C919 B.n879 VSUBS 0.009114f
C920 B.n880 VSUBS 0.009114f
C921 B.n881 VSUBS 0.009114f
C922 B.n882 VSUBS 0.009114f
C923 B.n883 VSUBS 0.009114f
C924 B.n884 VSUBS 0.009114f
C925 B.n885 VSUBS 0.009114f
C926 B.n886 VSUBS 0.009114f
C927 B.n887 VSUBS 0.009114f
C928 B.n888 VSUBS 0.009114f
C929 B.n889 VSUBS 0.009114f
C930 B.n890 VSUBS 0.009114f
C931 B.n891 VSUBS 0.009114f
C932 B.n892 VSUBS 0.009114f
C933 B.n893 VSUBS 0.009114f
C934 B.n894 VSUBS 0.009114f
C935 B.n895 VSUBS 0.009114f
C936 B.n896 VSUBS 0.009114f
C937 B.n897 VSUBS 0.009114f
C938 B.n898 VSUBS 0.020194f
C939 B.n899 VSUBS 0.020194f
C940 B.n900 VSUBS 0.019213f
C941 B.n901 VSUBS 0.009114f
C942 B.n902 VSUBS 0.009114f
C943 B.n903 VSUBS 0.009114f
C944 B.n904 VSUBS 0.009114f
C945 B.n905 VSUBS 0.009114f
C946 B.n906 VSUBS 0.009114f
C947 B.n907 VSUBS 0.009114f
C948 B.n908 VSUBS 0.009114f
C949 B.n909 VSUBS 0.009114f
C950 B.n910 VSUBS 0.009114f
C951 B.n911 VSUBS 0.009114f
C952 B.n912 VSUBS 0.009114f
C953 B.n913 VSUBS 0.009114f
C954 B.n914 VSUBS 0.009114f
C955 B.n915 VSUBS 0.009114f
C956 B.n916 VSUBS 0.009114f
C957 B.n917 VSUBS 0.009114f
C958 B.n918 VSUBS 0.009114f
C959 B.n919 VSUBS 0.009114f
C960 B.n920 VSUBS 0.009114f
C961 B.n921 VSUBS 0.009114f
C962 B.n922 VSUBS 0.009114f
C963 B.n923 VSUBS 0.009114f
C964 B.n924 VSUBS 0.009114f
C965 B.n925 VSUBS 0.009114f
C966 B.n926 VSUBS 0.009114f
C967 B.n927 VSUBS 0.009114f
C968 B.n928 VSUBS 0.009114f
C969 B.n929 VSUBS 0.009114f
C970 B.n930 VSUBS 0.009114f
C971 B.n931 VSUBS 0.009114f
C972 B.n932 VSUBS 0.009114f
C973 B.n933 VSUBS 0.009114f
C974 B.n934 VSUBS 0.009114f
C975 B.n935 VSUBS 0.009114f
C976 B.n936 VSUBS 0.009114f
C977 B.n937 VSUBS 0.009114f
C978 B.n938 VSUBS 0.009114f
C979 B.n939 VSUBS 0.009114f
C980 B.n940 VSUBS 0.009114f
C981 B.n941 VSUBS 0.009114f
C982 B.n942 VSUBS 0.009114f
C983 B.n943 VSUBS 0.009114f
C984 B.n944 VSUBS 0.009114f
C985 B.n945 VSUBS 0.009114f
C986 B.n946 VSUBS 0.009114f
C987 B.n947 VSUBS 0.009114f
C988 B.n948 VSUBS 0.009114f
C989 B.n949 VSUBS 0.009114f
C990 B.n950 VSUBS 0.009114f
C991 B.n951 VSUBS 0.009114f
C992 B.n952 VSUBS 0.009114f
C993 B.n953 VSUBS 0.009114f
C994 B.n954 VSUBS 0.009114f
C995 B.n955 VSUBS 0.009114f
C996 B.n956 VSUBS 0.009114f
C997 B.n957 VSUBS 0.009114f
C998 B.n958 VSUBS 0.009114f
C999 B.n959 VSUBS 0.009114f
C1000 B.n960 VSUBS 0.009114f
C1001 B.n961 VSUBS 0.009114f
C1002 B.n962 VSUBS 0.009114f
C1003 B.n963 VSUBS 0.009114f
C1004 B.n964 VSUBS 0.009114f
C1005 B.n965 VSUBS 0.009114f
C1006 B.n966 VSUBS 0.009114f
C1007 B.n967 VSUBS 0.009114f
C1008 B.n968 VSUBS 0.009114f
C1009 B.n969 VSUBS 0.009114f
C1010 B.n970 VSUBS 0.009114f
C1011 B.n971 VSUBS 0.009114f
C1012 B.n972 VSUBS 0.009114f
C1013 B.n973 VSUBS 0.009114f
C1014 B.n974 VSUBS 0.009114f
C1015 B.n975 VSUBS 0.009114f
C1016 B.n976 VSUBS 0.009114f
C1017 B.n977 VSUBS 0.009114f
C1018 B.n978 VSUBS 0.009114f
C1019 B.n979 VSUBS 0.009114f
C1020 B.n980 VSUBS 0.009114f
C1021 B.n981 VSUBS 0.009114f
C1022 B.n982 VSUBS 0.009114f
C1023 B.n983 VSUBS 0.009114f
C1024 B.n984 VSUBS 0.009114f
C1025 B.n985 VSUBS 0.009114f
C1026 B.n986 VSUBS 0.009114f
C1027 B.n987 VSUBS 0.009114f
C1028 B.n988 VSUBS 0.009114f
C1029 B.n989 VSUBS 0.009114f
C1030 B.n990 VSUBS 0.009114f
C1031 B.n991 VSUBS 0.009114f
C1032 B.n992 VSUBS 0.009114f
C1033 B.n993 VSUBS 0.009114f
C1034 B.n994 VSUBS 0.009114f
C1035 B.n995 VSUBS 0.009114f
C1036 B.n996 VSUBS 0.009114f
C1037 B.n997 VSUBS 0.009114f
C1038 B.n998 VSUBS 0.009114f
C1039 B.n999 VSUBS 0.009114f
C1040 B.n1000 VSUBS 0.009114f
C1041 B.n1001 VSUBS 0.009114f
C1042 B.n1002 VSUBS 0.009114f
C1043 B.n1003 VSUBS 0.009114f
C1044 B.n1004 VSUBS 0.009114f
C1045 B.n1005 VSUBS 0.009114f
C1046 B.n1006 VSUBS 0.009114f
C1047 B.n1007 VSUBS 0.009114f
C1048 B.n1008 VSUBS 0.009114f
C1049 B.n1009 VSUBS 0.009114f
C1050 B.n1010 VSUBS 0.009114f
C1051 B.n1011 VSUBS 0.009114f
C1052 B.n1012 VSUBS 0.009114f
C1053 B.n1013 VSUBS 0.009114f
C1054 B.n1014 VSUBS 0.009114f
C1055 B.n1015 VSUBS 0.009114f
C1056 B.n1016 VSUBS 0.009114f
C1057 B.n1017 VSUBS 0.009114f
C1058 B.n1018 VSUBS 0.009114f
C1059 B.n1019 VSUBS 0.009114f
C1060 B.n1020 VSUBS 0.009114f
C1061 B.n1021 VSUBS 0.009114f
C1062 B.n1022 VSUBS 0.009114f
C1063 B.n1023 VSUBS 0.011894f
C1064 B.n1024 VSUBS 0.01267f
C1065 B.n1025 VSUBS 0.025195f
C1066 VDD2.n0 VSUBS 0.035427f
C1067 VDD2.n1 VSUBS 0.031872f
C1068 VDD2.n2 VSUBS 0.017126f
C1069 VDD2.n3 VSUBS 0.040481f
C1070 VDD2.n4 VSUBS 0.018134f
C1071 VDD2.n5 VSUBS 0.031872f
C1072 VDD2.n6 VSUBS 0.017126f
C1073 VDD2.n7 VSUBS 0.040481f
C1074 VDD2.n8 VSUBS 0.018134f
C1075 VDD2.n9 VSUBS 0.031872f
C1076 VDD2.n10 VSUBS 0.017126f
C1077 VDD2.n11 VSUBS 0.040481f
C1078 VDD2.n12 VSUBS 0.018134f
C1079 VDD2.n13 VSUBS 0.031872f
C1080 VDD2.n14 VSUBS 0.017126f
C1081 VDD2.n15 VSUBS 0.040481f
C1082 VDD2.n16 VSUBS 0.018134f
C1083 VDD2.n17 VSUBS 0.233728f
C1084 VDD2.t1 VSUBS 0.087118f
C1085 VDD2.n18 VSUBS 0.03036f
C1086 VDD2.n19 VSUBS 0.030452f
C1087 VDD2.n20 VSUBS 0.017126f
C1088 VDD2.n21 VSUBS 1.39834f
C1089 VDD2.n22 VSUBS 0.031872f
C1090 VDD2.n23 VSUBS 0.017126f
C1091 VDD2.n24 VSUBS 0.018134f
C1092 VDD2.n25 VSUBS 0.040481f
C1093 VDD2.n26 VSUBS 0.040481f
C1094 VDD2.n27 VSUBS 0.018134f
C1095 VDD2.n28 VSUBS 0.017126f
C1096 VDD2.n29 VSUBS 0.031872f
C1097 VDD2.n30 VSUBS 0.031872f
C1098 VDD2.n31 VSUBS 0.017126f
C1099 VDD2.n32 VSUBS 0.018134f
C1100 VDD2.n33 VSUBS 0.040481f
C1101 VDD2.n34 VSUBS 0.040481f
C1102 VDD2.n35 VSUBS 0.040481f
C1103 VDD2.n36 VSUBS 0.018134f
C1104 VDD2.n37 VSUBS 0.017126f
C1105 VDD2.n38 VSUBS 0.031872f
C1106 VDD2.n39 VSUBS 0.031872f
C1107 VDD2.n40 VSUBS 0.017126f
C1108 VDD2.n41 VSUBS 0.01763f
C1109 VDD2.n42 VSUBS 0.01763f
C1110 VDD2.n43 VSUBS 0.040481f
C1111 VDD2.n44 VSUBS 0.040481f
C1112 VDD2.n45 VSUBS 0.018134f
C1113 VDD2.n46 VSUBS 0.017126f
C1114 VDD2.n47 VSUBS 0.031872f
C1115 VDD2.n48 VSUBS 0.031872f
C1116 VDD2.n49 VSUBS 0.017126f
C1117 VDD2.n50 VSUBS 0.018134f
C1118 VDD2.n51 VSUBS 0.040481f
C1119 VDD2.n52 VSUBS 0.099386f
C1120 VDD2.n53 VSUBS 0.018134f
C1121 VDD2.n54 VSUBS 0.017126f
C1122 VDD2.n55 VSUBS 0.078894f
C1123 VDD2.n56 VSUBS 0.101719f
C1124 VDD2.t7 VSUBS 0.272007f
C1125 VDD2.t3 VSUBS 0.272007f
C1126 VDD2.n57 VSUBS 2.09236f
C1127 VDD2.n58 VSUBS 1.45549f
C1128 VDD2.t0 VSUBS 0.272007f
C1129 VDD2.t2 VSUBS 0.272007f
C1130 VDD2.n59 VSUBS 2.13388f
C1131 VDD2.n60 VSUBS 4.80119f
C1132 VDD2.n61 VSUBS 0.035427f
C1133 VDD2.n62 VSUBS 0.031872f
C1134 VDD2.n63 VSUBS 0.017126f
C1135 VDD2.n64 VSUBS 0.040481f
C1136 VDD2.n65 VSUBS 0.018134f
C1137 VDD2.n66 VSUBS 0.031872f
C1138 VDD2.n67 VSUBS 0.017126f
C1139 VDD2.n68 VSUBS 0.040481f
C1140 VDD2.n69 VSUBS 0.018134f
C1141 VDD2.n70 VSUBS 0.031872f
C1142 VDD2.n71 VSUBS 0.017126f
C1143 VDD2.n72 VSUBS 0.040481f
C1144 VDD2.n73 VSUBS 0.040481f
C1145 VDD2.n74 VSUBS 0.018134f
C1146 VDD2.n75 VSUBS 0.031872f
C1147 VDD2.n76 VSUBS 0.017126f
C1148 VDD2.n77 VSUBS 0.040481f
C1149 VDD2.n78 VSUBS 0.018134f
C1150 VDD2.n79 VSUBS 0.233728f
C1151 VDD2.t6 VSUBS 0.087118f
C1152 VDD2.n80 VSUBS 0.03036f
C1153 VDD2.n81 VSUBS 0.030452f
C1154 VDD2.n82 VSUBS 0.017126f
C1155 VDD2.n83 VSUBS 1.39834f
C1156 VDD2.n84 VSUBS 0.031872f
C1157 VDD2.n85 VSUBS 0.017126f
C1158 VDD2.n86 VSUBS 0.018134f
C1159 VDD2.n87 VSUBS 0.040481f
C1160 VDD2.n88 VSUBS 0.040481f
C1161 VDD2.n89 VSUBS 0.018134f
C1162 VDD2.n90 VSUBS 0.017126f
C1163 VDD2.n91 VSUBS 0.031872f
C1164 VDD2.n92 VSUBS 0.031872f
C1165 VDD2.n93 VSUBS 0.017126f
C1166 VDD2.n94 VSUBS 0.018134f
C1167 VDD2.n95 VSUBS 0.040481f
C1168 VDD2.n96 VSUBS 0.040481f
C1169 VDD2.n97 VSUBS 0.018134f
C1170 VDD2.n98 VSUBS 0.017126f
C1171 VDD2.n99 VSUBS 0.031872f
C1172 VDD2.n100 VSUBS 0.031872f
C1173 VDD2.n101 VSUBS 0.017126f
C1174 VDD2.n102 VSUBS 0.01763f
C1175 VDD2.n103 VSUBS 0.01763f
C1176 VDD2.n104 VSUBS 0.040481f
C1177 VDD2.n105 VSUBS 0.040481f
C1178 VDD2.n106 VSUBS 0.018134f
C1179 VDD2.n107 VSUBS 0.017126f
C1180 VDD2.n108 VSUBS 0.031872f
C1181 VDD2.n109 VSUBS 0.031872f
C1182 VDD2.n110 VSUBS 0.017126f
C1183 VDD2.n111 VSUBS 0.018134f
C1184 VDD2.n112 VSUBS 0.040481f
C1185 VDD2.n113 VSUBS 0.099386f
C1186 VDD2.n114 VSUBS 0.018134f
C1187 VDD2.n115 VSUBS 0.017126f
C1188 VDD2.n116 VSUBS 0.078894f
C1189 VDD2.n117 VSUBS 0.072166f
C1190 VDD2.n118 VSUBS 4.23226f
C1191 VDD2.t4 VSUBS 0.272007f
C1192 VDD2.t8 VSUBS 0.272007f
C1193 VDD2.n119 VSUBS 2.09237f
C1194 VDD2.n120 VSUBS 1.05433f
C1195 VDD2.t9 VSUBS 0.272007f
C1196 VDD2.t5 VSUBS 0.272007f
C1197 VDD2.n121 VSUBS 2.13382f
C1198 VN.t7 VSUBS 2.72474f
C1199 VN.n0 VSUBS 1.04886f
C1200 VN.n1 VSUBS 0.023636f
C1201 VN.n2 VSUBS 0.047348f
C1202 VN.n3 VSUBS 0.023636f
C1203 VN.n4 VSUBS 0.044273f
C1204 VN.n5 VSUBS 0.023636f
C1205 VN.t9 VSUBS 2.72474f
C1206 VN.n6 VSUBS 0.044273f
C1207 VN.n7 VSUBS 0.023636f
C1208 VN.n8 VSUBS 0.044273f
C1209 VN.n9 VSUBS 0.023636f
C1210 VN.t6 VSUBS 2.72474f
C1211 VN.n10 VSUBS 0.044273f
C1212 VN.n11 VSUBS 0.023636f
C1213 VN.n12 VSUBS 0.044273f
C1214 VN.n13 VSUBS 0.309051f
C1215 VN.t2 VSUBS 2.72474f
C1216 VN.t8 VSUBS 3.10156f
C1217 VN.n14 VSUBS 0.999688f
C1218 VN.n15 VSUBS 1.046f
C1219 VN.n16 VSUBS 0.033781f
C1220 VN.n17 VSUBS 0.044273f
C1221 VN.n18 VSUBS 0.023636f
C1222 VN.n19 VSUBS 0.023636f
C1223 VN.n20 VSUBS 0.023636f
C1224 VN.n21 VSUBS 0.042144f
C1225 VN.n22 VSUBS 0.024858f
C1226 VN.n23 VSUBS 0.046582f
C1227 VN.n24 VSUBS 0.023636f
C1228 VN.n25 VSUBS 0.023636f
C1229 VN.n26 VSUBS 0.023636f
C1230 VN.n27 VSUBS 0.044273f
C1231 VN.n28 VSUBS 0.981446f
C1232 VN.n29 VSUBS 0.044273f
C1233 VN.n30 VSUBS 0.023636f
C1234 VN.n31 VSUBS 0.023636f
C1235 VN.n32 VSUBS 0.023636f
C1236 VN.n33 VSUBS 0.046582f
C1237 VN.n34 VSUBS 0.024858f
C1238 VN.n35 VSUBS 0.042144f
C1239 VN.n36 VSUBS 0.023636f
C1240 VN.n37 VSUBS 0.023636f
C1241 VN.n38 VSUBS 0.023636f
C1242 VN.n39 VSUBS 0.044273f
C1243 VN.n40 VSUBS 0.033781f
C1244 VN.n41 VSUBS 0.959032f
C1245 VN.n42 VSUBS 0.032907f
C1246 VN.n43 VSUBS 0.023636f
C1247 VN.n44 VSUBS 0.023636f
C1248 VN.n45 VSUBS 0.023636f
C1249 VN.n46 VSUBS 0.044273f
C1250 VN.n47 VSUBS 0.043128f
C1251 VN.n48 VSUBS 0.023107f
C1252 VN.n49 VSUBS 0.023636f
C1253 VN.n50 VSUBS 0.023636f
C1254 VN.n51 VSUBS 0.023636f
C1255 VN.n52 VSUBS 0.044273f
C1256 VN.n53 VSUBS 0.044273f
C1257 VN.n54 VSUBS 0.023288f
C1258 VN.n55 VSUBS 0.038155f
C1259 VN.n56 VSUBS 0.075781f
C1260 VN.t3 VSUBS 2.72474f
C1261 VN.n57 VSUBS 1.04886f
C1262 VN.n58 VSUBS 0.023636f
C1263 VN.n59 VSUBS 0.047348f
C1264 VN.n60 VSUBS 0.023636f
C1265 VN.n61 VSUBS 0.044273f
C1266 VN.n62 VSUBS 0.023636f
C1267 VN.t5 VSUBS 2.72474f
C1268 VN.n63 VSUBS 0.044273f
C1269 VN.n64 VSUBS 0.023636f
C1270 VN.n65 VSUBS 0.044273f
C1271 VN.n66 VSUBS 0.023636f
C1272 VN.t1 VSUBS 2.72474f
C1273 VN.n67 VSUBS 0.044273f
C1274 VN.n68 VSUBS 0.023636f
C1275 VN.n69 VSUBS 0.044273f
C1276 VN.n70 VSUBS 0.309051f
C1277 VN.t0 VSUBS 2.72474f
C1278 VN.t4 VSUBS 3.10156f
C1279 VN.n71 VSUBS 0.999688f
C1280 VN.n72 VSUBS 1.046f
C1281 VN.n73 VSUBS 0.033781f
C1282 VN.n74 VSUBS 0.044273f
C1283 VN.n75 VSUBS 0.023636f
C1284 VN.n76 VSUBS 0.023636f
C1285 VN.n77 VSUBS 0.023636f
C1286 VN.n78 VSUBS 0.042144f
C1287 VN.n79 VSUBS 0.024858f
C1288 VN.n80 VSUBS 0.046582f
C1289 VN.n81 VSUBS 0.023636f
C1290 VN.n82 VSUBS 0.023636f
C1291 VN.n83 VSUBS 0.023636f
C1292 VN.n84 VSUBS 0.044273f
C1293 VN.n85 VSUBS 0.981446f
C1294 VN.n86 VSUBS 0.044273f
C1295 VN.n87 VSUBS 0.023636f
C1296 VN.n88 VSUBS 0.023636f
C1297 VN.n89 VSUBS 0.023636f
C1298 VN.n90 VSUBS 0.046582f
C1299 VN.n91 VSUBS 0.024858f
C1300 VN.n92 VSUBS 0.042144f
C1301 VN.n93 VSUBS 0.023636f
C1302 VN.n94 VSUBS 0.023636f
C1303 VN.n95 VSUBS 0.023636f
C1304 VN.n96 VSUBS 0.044273f
C1305 VN.n97 VSUBS 0.033781f
C1306 VN.n98 VSUBS 0.959032f
C1307 VN.n99 VSUBS 0.032907f
C1308 VN.n100 VSUBS 0.023636f
C1309 VN.n101 VSUBS 0.023636f
C1310 VN.n102 VSUBS 0.023636f
C1311 VN.n103 VSUBS 0.044273f
C1312 VN.n104 VSUBS 0.043128f
C1313 VN.n105 VSUBS 0.023107f
C1314 VN.n106 VSUBS 0.023636f
C1315 VN.n107 VSUBS 0.023636f
C1316 VN.n108 VSUBS 0.023636f
C1317 VN.n109 VSUBS 0.044273f
C1318 VN.n110 VSUBS 0.044273f
C1319 VN.n111 VSUBS 0.023288f
C1320 VN.n112 VSUBS 0.038155f
C1321 VN.n113 VSUBS 1.73958f
C1322 VTAIL.t19 VSUBS 0.262209f
C1323 VTAIL.t1 VSUBS 0.262209f
C1324 VTAIL.n0 VSUBS 1.86778f
C1325 VTAIL.n1 VSUBS 1.17032f
C1326 VTAIL.n2 VSUBS 0.034151f
C1327 VTAIL.n3 VSUBS 0.030723f
C1328 VTAIL.n4 VSUBS 0.01651f
C1329 VTAIL.n5 VSUBS 0.039022f
C1330 VTAIL.n6 VSUBS 0.017481f
C1331 VTAIL.n7 VSUBS 0.030723f
C1332 VTAIL.n8 VSUBS 0.01651f
C1333 VTAIL.n9 VSUBS 0.039022f
C1334 VTAIL.n10 VSUBS 0.017481f
C1335 VTAIL.n11 VSUBS 0.030723f
C1336 VTAIL.n12 VSUBS 0.01651f
C1337 VTAIL.n13 VSUBS 0.039022f
C1338 VTAIL.n14 VSUBS 0.017481f
C1339 VTAIL.n15 VSUBS 0.030723f
C1340 VTAIL.n16 VSUBS 0.01651f
C1341 VTAIL.n17 VSUBS 0.039022f
C1342 VTAIL.n18 VSUBS 0.017481f
C1343 VTAIL.n19 VSUBS 0.225308f
C1344 VTAIL.t13 VSUBS 0.083979f
C1345 VTAIL.n20 VSUBS 0.029267f
C1346 VTAIL.n21 VSUBS 0.029355f
C1347 VTAIL.n22 VSUBS 0.01651f
C1348 VTAIL.n23 VSUBS 1.34797f
C1349 VTAIL.n24 VSUBS 0.030723f
C1350 VTAIL.n25 VSUBS 0.01651f
C1351 VTAIL.n26 VSUBS 0.017481f
C1352 VTAIL.n27 VSUBS 0.039022f
C1353 VTAIL.n28 VSUBS 0.039022f
C1354 VTAIL.n29 VSUBS 0.017481f
C1355 VTAIL.n30 VSUBS 0.01651f
C1356 VTAIL.n31 VSUBS 0.030723f
C1357 VTAIL.n32 VSUBS 0.030723f
C1358 VTAIL.n33 VSUBS 0.01651f
C1359 VTAIL.n34 VSUBS 0.017481f
C1360 VTAIL.n35 VSUBS 0.039022f
C1361 VTAIL.n36 VSUBS 0.039022f
C1362 VTAIL.n37 VSUBS 0.039022f
C1363 VTAIL.n38 VSUBS 0.017481f
C1364 VTAIL.n39 VSUBS 0.01651f
C1365 VTAIL.n40 VSUBS 0.030723f
C1366 VTAIL.n41 VSUBS 0.030723f
C1367 VTAIL.n42 VSUBS 0.01651f
C1368 VTAIL.n43 VSUBS 0.016995f
C1369 VTAIL.n44 VSUBS 0.016995f
C1370 VTAIL.n45 VSUBS 0.039022f
C1371 VTAIL.n46 VSUBS 0.039022f
C1372 VTAIL.n47 VSUBS 0.017481f
C1373 VTAIL.n48 VSUBS 0.01651f
C1374 VTAIL.n49 VSUBS 0.030723f
C1375 VTAIL.n50 VSUBS 0.030723f
C1376 VTAIL.n51 VSUBS 0.01651f
C1377 VTAIL.n52 VSUBS 0.017481f
C1378 VTAIL.n53 VSUBS 0.039022f
C1379 VTAIL.n54 VSUBS 0.095806f
C1380 VTAIL.n55 VSUBS 0.017481f
C1381 VTAIL.n56 VSUBS 0.01651f
C1382 VTAIL.n57 VSUBS 0.076052f
C1383 VTAIL.n58 VSUBS 0.048389f
C1384 VTAIL.n59 VSUBS 0.620941f
C1385 VTAIL.t12 VSUBS 0.262209f
C1386 VTAIL.t8 VSUBS 0.262209f
C1387 VTAIL.n60 VSUBS 1.86778f
C1388 VTAIL.n61 VSUBS 1.39072f
C1389 VTAIL.t15 VSUBS 0.262209f
C1390 VTAIL.t9 VSUBS 0.262209f
C1391 VTAIL.n62 VSUBS 1.86778f
C1392 VTAIL.n63 VSUBS 3.09332f
C1393 VTAIL.t3 VSUBS 0.262209f
C1394 VTAIL.t5 VSUBS 0.262209f
C1395 VTAIL.n64 VSUBS 1.86779f
C1396 VTAIL.n65 VSUBS 3.09331f
C1397 VTAIL.t6 VSUBS 0.262209f
C1398 VTAIL.t2 VSUBS 0.262209f
C1399 VTAIL.n66 VSUBS 1.86779f
C1400 VTAIL.n67 VSUBS 1.39071f
C1401 VTAIL.n68 VSUBS 0.034151f
C1402 VTAIL.n69 VSUBS 0.030723f
C1403 VTAIL.n70 VSUBS 0.01651f
C1404 VTAIL.n71 VSUBS 0.039022f
C1405 VTAIL.n72 VSUBS 0.017481f
C1406 VTAIL.n73 VSUBS 0.030723f
C1407 VTAIL.n74 VSUBS 0.01651f
C1408 VTAIL.n75 VSUBS 0.039022f
C1409 VTAIL.n76 VSUBS 0.017481f
C1410 VTAIL.n77 VSUBS 0.030723f
C1411 VTAIL.n78 VSUBS 0.01651f
C1412 VTAIL.n79 VSUBS 0.039022f
C1413 VTAIL.n80 VSUBS 0.039022f
C1414 VTAIL.n81 VSUBS 0.017481f
C1415 VTAIL.n82 VSUBS 0.030723f
C1416 VTAIL.n83 VSUBS 0.01651f
C1417 VTAIL.n84 VSUBS 0.039022f
C1418 VTAIL.n85 VSUBS 0.017481f
C1419 VTAIL.n86 VSUBS 0.225308f
C1420 VTAIL.t0 VSUBS 0.083979f
C1421 VTAIL.n87 VSUBS 0.029267f
C1422 VTAIL.n88 VSUBS 0.029355f
C1423 VTAIL.n89 VSUBS 0.01651f
C1424 VTAIL.n90 VSUBS 1.34797f
C1425 VTAIL.n91 VSUBS 0.030723f
C1426 VTAIL.n92 VSUBS 0.01651f
C1427 VTAIL.n93 VSUBS 0.017481f
C1428 VTAIL.n94 VSUBS 0.039022f
C1429 VTAIL.n95 VSUBS 0.039022f
C1430 VTAIL.n96 VSUBS 0.017481f
C1431 VTAIL.n97 VSUBS 0.01651f
C1432 VTAIL.n98 VSUBS 0.030723f
C1433 VTAIL.n99 VSUBS 0.030723f
C1434 VTAIL.n100 VSUBS 0.01651f
C1435 VTAIL.n101 VSUBS 0.017481f
C1436 VTAIL.n102 VSUBS 0.039022f
C1437 VTAIL.n103 VSUBS 0.039022f
C1438 VTAIL.n104 VSUBS 0.017481f
C1439 VTAIL.n105 VSUBS 0.01651f
C1440 VTAIL.n106 VSUBS 0.030723f
C1441 VTAIL.n107 VSUBS 0.030723f
C1442 VTAIL.n108 VSUBS 0.01651f
C1443 VTAIL.n109 VSUBS 0.016995f
C1444 VTAIL.n110 VSUBS 0.016995f
C1445 VTAIL.n111 VSUBS 0.039022f
C1446 VTAIL.n112 VSUBS 0.039022f
C1447 VTAIL.n113 VSUBS 0.017481f
C1448 VTAIL.n114 VSUBS 0.01651f
C1449 VTAIL.n115 VSUBS 0.030723f
C1450 VTAIL.n116 VSUBS 0.030723f
C1451 VTAIL.n117 VSUBS 0.01651f
C1452 VTAIL.n118 VSUBS 0.017481f
C1453 VTAIL.n119 VSUBS 0.039022f
C1454 VTAIL.n120 VSUBS 0.095806f
C1455 VTAIL.n121 VSUBS 0.017481f
C1456 VTAIL.n122 VSUBS 0.01651f
C1457 VTAIL.n123 VSUBS 0.076052f
C1458 VTAIL.n124 VSUBS 0.048389f
C1459 VTAIL.n125 VSUBS 0.620941f
C1460 VTAIL.t14 VSUBS 0.262209f
C1461 VTAIL.t17 VSUBS 0.262209f
C1462 VTAIL.n126 VSUBS 1.86779f
C1463 VTAIL.n127 VSUBS 1.25544f
C1464 VTAIL.t11 VSUBS 0.262209f
C1465 VTAIL.t16 VSUBS 0.262209f
C1466 VTAIL.n128 VSUBS 1.86779f
C1467 VTAIL.n129 VSUBS 1.39071f
C1468 VTAIL.n130 VSUBS 0.034151f
C1469 VTAIL.n131 VSUBS 0.030723f
C1470 VTAIL.n132 VSUBS 0.01651f
C1471 VTAIL.n133 VSUBS 0.039022f
C1472 VTAIL.n134 VSUBS 0.017481f
C1473 VTAIL.n135 VSUBS 0.030723f
C1474 VTAIL.n136 VSUBS 0.01651f
C1475 VTAIL.n137 VSUBS 0.039022f
C1476 VTAIL.n138 VSUBS 0.017481f
C1477 VTAIL.n139 VSUBS 0.030723f
C1478 VTAIL.n140 VSUBS 0.01651f
C1479 VTAIL.n141 VSUBS 0.039022f
C1480 VTAIL.n142 VSUBS 0.039022f
C1481 VTAIL.n143 VSUBS 0.017481f
C1482 VTAIL.n144 VSUBS 0.030723f
C1483 VTAIL.n145 VSUBS 0.01651f
C1484 VTAIL.n146 VSUBS 0.039022f
C1485 VTAIL.n147 VSUBS 0.017481f
C1486 VTAIL.n148 VSUBS 0.225308f
C1487 VTAIL.t10 VSUBS 0.083979f
C1488 VTAIL.n149 VSUBS 0.029267f
C1489 VTAIL.n150 VSUBS 0.029355f
C1490 VTAIL.n151 VSUBS 0.01651f
C1491 VTAIL.n152 VSUBS 1.34797f
C1492 VTAIL.n153 VSUBS 0.030723f
C1493 VTAIL.n154 VSUBS 0.01651f
C1494 VTAIL.n155 VSUBS 0.017481f
C1495 VTAIL.n156 VSUBS 0.039022f
C1496 VTAIL.n157 VSUBS 0.039022f
C1497 VTAIL.n158 VSUBS 0.017481f
C1498 VTAIL.n159 VSUBS 0.01651f
C1499 VTAIL.n160 VSUBS 0.030723f
C1500 VTAIL.n161 VSUBS 0.030723f
C1501 VTAIL.n162 VSUBS 0.01651f
C1502 VTAIL.n163 VSUBS 0.017481f
C1503 VTAIL.n164 VSUBS 0.039022f
C1504 VTAIL.n165 VSUBS 0.039022f
C1505 VTAIL.n166 VSUBS 0.017481f
C1506 VTAIL.n167 VSUBS 0.01651f
C1507 VTAIL.n168 VSUBS 0.030723f
C1508 VTAIL.n169 VSUBS 0.030723f
C1509 VTAIL.n170 VSUBS 0.01651f
C1510 VTAIL.n171 VSUBS 0.016995f
C1511 VTAIL.n172 VSUBS 0.016995f
C1512 VTAIL.n173 VSUBS 0.039022f
C1513 VTAIL.n174 VSUBS 0.039022f
C1514 VTAIL.n175 VSUBS 0.017481f
C1515 VTAIL.n176 VSUBS 0.01651f
C1516 VTAIL.n177 VSUBS 0.030723f
C1517 VTAIL.n178 VSUBS 0.030723f
C1518 VTAIL.n179 VSUBS 0.01651f
C1519 VTAIL.n180 VSUBS 0.017481f
C1520 VTAIL.n181 VSUBS 0.039022f
C1521 VTAIL.n182 VSUBS 0.095806f
C1522 VTAIL.n183 VSUBS 0.017481f
C1523 VTAIL.n184 VSUBS 0.01651f
C1524 VTAIL.n185 VSUBS 0.076052f
C1525 VTAIL.n186 VSUBS 0.048389f
C1526 VTAIL.n187 VSUBS 2.09526f
C1527 VTAIL.n188 VSUBS 0.034151f
C1528 VTAIL.n189 VSUBS 0.030723f
C1529 VTAIL.n190 VSUBS 0.01651f
C1530 VTAIL.n191 VSUBS 0.039022f
C1531 VTAIL.n192 VSUBS 0.017481f
C1532 VTAIL.n193 VSUBS 0.030723f
C1533 VTAIL.n194 VSUBS 0.01651f
C1534 VTAIL.n195 VSUBS 0.039022f
C1535 VTAIL.n196 VSUBS 0.017481f
C1536 VTAIL.n197 VSUBS 0.030723f
C1537 VTAIL.n198 VSUBS 0.01651f
C1538 VTAIL.n199 VSUBS 0.039022f
C1539 VTAIL.n200 VSUBS 0.017481f
C1540 VTAIL.n201 VSUBS 0.030723f
C1541 VTAIL.n202 VSUBS 0.01651f
C1542 VTAIL.n203 VSUBS 0.039022f
C1543 VTAIL.n204 VSUBS 0.017481f
C1544 VTAIL.n205 VSUBS 0.225308f
C1545 VTAIL.t4 VSUBS 0.083979f
C1546 VTAIL.n206 VSUBS 0.029267f
C1547 VTAIL.n207 VSUBS 0.029355f
C1548 VTAIL.n208 VSUBS 0.01651f
C1549 VTAIL.n209 VSUBS 1.34797f
C1550 VTAIL.n210 VSUBS 0.030723f
C1551 VTAIL.n211 VSUBS 0.01651f
C1552 VTAIL.n212 VSUBS 0.017481f
C1553 VTAIL.n213 VSUBS 0.039022f
C1554 VTAIL.n214 VSUBS 0.039022f
C1555 VTAIL.n215 VSUBS 0.017481f
C1556 VTAIL.n216 VSUBS 0.01651f
C1557 VTAIL.n217 VSUBS 0.030723f
C1558 VTAIL.n218 VSUBS 0.030723f
C1559 VTAIL.n219 VSUBS 0.01651f
C1560 VTAIL.n220 VSUBS 0.017481f
C1561 VTAIL.n221 VSUBS 0.039022f
C1562 VTAIL.n222 VSUBS 0.039022f
C1563 VTAIL.n223 VSUBS 0.039022f
C1564 VTAIL.n224 VSUBS 0.017481f
C1565 VTAIL.n225 VSUBS 0.01651f
C1566 VTAIL.n226 VSUBS 0.030723f
C1567 VTAIL.n227 VSUBS 0.030723f
C1568 VTAIL.n228 VSUBS 0.01651f
C1569 VTAIL.n229 VSUBS 0.016995f
C1570 VTAIL.n230 VSUBS 0.016995f
C1571 VTAIL.n231 VSUBS 0.039022f
C1572 VTAIL.n232 VSUBS 0.039022f
C1573 VTAIL.n233 VSUBS 0.017481f
C1574 VTAIL.n234 VSUBS 0.01651f
C1575 VTAIL.n235 VSUBS 0.030723f
C1576 VTAIL.n236 VSUBS 0.030723f
C1577 VTAIL.n237 VSUBS 0.01651f
C1578 VTAIL.n238 VSUBS 0.017481f
C1579 VTAIL.n239 VSUBS 0.039022f
C1580 VTAIL.n240 VSUBS 0.095806f
C1581 VTAIL.n241 VSUBS 0.017481f
C1582 VTAIL.n242 VSUBS 0.01651f
C1583 VTAIL.n243 VSUBS 0.076052f
C1584 VTAIL.n244 VSUBS 0.048389f
C1585 VTAIL.n245 VSUBS 2.09526f
C1586 VTAIL.t18 VSUBS 0.262209f
C1587 VTAIL.t7 VSUBS 0.262209f
C1588 VTAIL.n246 VSUBS 1.86778f
C1589 VTAIL.n247 VSUBS 1.11229f
C1590 VDD1.n0 VSUBS 0.035522f
C1591 VDD1.n1 VSUBS 0.031957f
C1592 VDD1.n2 VSUBS 0.017172f
C1593 VDD1.n3 VSUBS 0.040589f
C1594 VDD1.n4 VSUBS 0.018183f
C1595 VDD1.n5 VSUBS 0.031957f
C1596 VDD1.n6 VSUBS 0.017172f
C1597 VDD1.n7 VSUBS 0.040589f
C1598 VDD1.n8 VSUBS 0.018183f
C1599 VDD1.n9 VSUBS 0.031957f
C1600 VDD1.n10 VSUBS 0.017172f
C1601 VDD1.n11 VSUBS 0.040589f
C1602 VDD1.n12 VSUBS 0.040589f
C1603 VDD1.n13 VSUBS 0.018183f
C1604 VDD1.n14 VSUBS 0.031957f
C1605 VDD1.n15 VSUBS 0.017172f
C1606 VDD1.n16 VSUBS 0.040589f
C1607 VDD1.n17 VSUBS 0.018183f
C1608 VDD1.n18 VSUBS 0.234356f
C1609 VDD1.t2 VSUBS 0.087352f
C1610 VDD1.n19 VSUBS 0.030442f
C1611 VDD1.n20 VSUBS 0.030534f
C1612 VDD1.n21 VSUBS 0.017172f
C1613 VDD1.n22 VSUBS 1.4021f
C1614 VDD1.n23 VSUBS 0.031957f
C1615 VDD1.n24 VSUBS 0.017172f
C1616 VDD1.n25 VSUBS 0.018183f
C1617 VDD1.n26 VSUBS 0.040589f
C1618 VDD1.n27 VSUBS 0.040589f
C1619 VDD1.n28 VSUBS 0.018183f
C1620 VDD1.n29 VSUBS 0.017172f
C1621 VDD1.n30 VSUBS 0.031957f
C1622 VDD1.n31 VSUBS 0.031957f
C1623 VDD1.n32 VSUBS 0.017172f
C1624 VDD1.n33 VSUBS 0.018183f
C1625 VDD1.n34 VSUBS 0.040589f
C1626 VDD1.n35 VSUBS 0.040589f
C1627 VDD1.n36 VSUBS 0.018183f
C1628 VDD1.n37 VSUBS 0.017172f
C1629 VDD1.n38 VSUBS 0.031957f
C1630 VDD1.n39 VSUBS 0.031957f
C1631 VDD1.n40 VSUBS 0.017172f
C1632 VDD1.n41 VSUBS 0.017677f
C1633 VDD1.n42 VSUBS 0.017677f
C1634 VDD1.n43 VSUBS 0.040589f
C1635 VDD1.n44 VSUBS 0.040589f
C1636 VDD1.n45 VSUBS 0.018183f
C1637 VDD1.n46 VSUBS 0.017172f
C1638 VDD1.n47 VSUBS 0.031957f
C1639 VDD1.n48 VSUBS 0.031957f
C1640 VDD1.n49 VSUBS 0.017172f
C1641 VDD1.n50 VSUBS 0.018183f
C1642 VDD1.n51 VSUBS 0.040589f
C1643 VDD1.n52 VSUBS 0.099653f
C1644 VDD1.n53 VSUBS 0.018183f
C1645 VDD1.n54 VSUBS 0.017172f
C1646 VDD1.n55 VSUBS 0.079106f
C1647 VDD1.n56 VSUBS 0.101993f
C1648 VDD1.t1 VSUBS 0.272738f
C1649 VDD1.t9 VSUBS 0.272738f
C1650 VDD1.n57 VSUBS 2.09799f
C1651 VDD1.n58 VSUBS 1.47023f
C1652 VDD1.n59 VSUBS 0.035522f
C1653 VDD1.n60 VSUBS 0.031957f
C1654 VDD1.n61 VSUBS 0.017172f
C1655 VDD1.n62 VSUBS 0.040589f
C1656 VDD1.n63 VSUBS 0.018183f
C1657 VDD1.n64 VSUBS 0.031957f
C1658 VDD1.n65 VSUBS 0.017172f
C1659 VDD1.n66 VSUBS 0.040589f
C1660 VDD1.n67 VSUBS 0.018183f
C1661 VDD1.n68 VSUBS 0.031957f
C1662 VDD1.n69 VSUBS 0.017172f
C1663 VDD1.n70 VSUBS 0.040589f
C1664 VDD1.n71 VSUBS 0.018183f
C1665 VDD1.n72 VSUBS 0.031957f
C1666 VDD1.n73 VSUBS 0.017172f
C1667 VDD1.n74 VSUBS 0.040589f
C1668 VDD1.n75 VSUBS 0.018183f
C1669 VDD1.n76 VSUBS 0.234356f
C1670 VDD1.t3 VSUBS 0.087352f
C1671 VDD1.n77 VSUBS 0.030442f
C1672 VDD1.n78 VSUBS 0.030534f
C1673 VDD1.n79 VSUBS 0.017172f
C1674 VDD1.n80 VSUBS 1.4021f
C1675 VDD1.n81 VSUBS 0.031957f
C1676 VDD1.n82 VSUBS 0.017172f
C1677 VDD1.n83 VSUBS 0.018183f
C1678 VDD1.n84 VSUBS 0.040589f
C1679 VDD1.n85 VSUBS 0.040589f
C1680 VDD1.n86 VSUBS 0.018183f
C1681 VDD1.n87 VSUBS 0.017172f
C1682 VDD1.n88 VSUBS 0.031957f
C1683 VDD1.n89 VSUBS 0.031957f
C1684 VDD1.n90 VSUBS 0.017172f
C1685 VDD1.n91 VSUBS 0.018183f
C1686 VDD1.n92 VSUBS 0.040589f
C1687 VDD1.n93 VSUBS 0.040589f
C1688 VDD1.n94 VSUBS 0.040589f
C1689 VDD1.n95 VSUBS 0.018183f
C1690 VDD1.n96 VSUBS 0.017172f
C1691 VDD1.n97 VSUBS 0.031957f
C1692 VDD1.n98 VSUBS 0.031957f
C1693 VDD1.n99 VSUBS 0.017172f
C1694 VDD1.n100 VSUBS 0.017677f
C1695 VDD1.n101 VSUBS 0.017677f
C1696 VDD1.n102 VSUBS 0.040589f
C1697 VDD1.n103 VSUBS 0.040589f
C1698 VDD1.n104 VSUBS 0.018183f
C1699 VDD1.n105 VSUBS 0.017172f
C1700 VDD1.n106 VSUBS 0.031957f
C1701 VDD1.n107 VSUBS 0.031957f
C1702 VDD1.n108 VSUBS 0.017172f
C1703 VDD1.n109 VSUBS 0.018183f
C1704 VDD1.n110 VSUBS 0.040589f
C1705 VDD1.n111 VSUBS 0.099653f
C1706 VDD1.n112 VSUBS 0.018183f
C1707 VDD1.n113 VSUBS 0.017172f
C1708 VDD1.n114 VSUBS 0.079106f
C1709 VDD1.n115 VSUBS 0.101993f
C1710 VDD1.t7 VSUBS 0.272738f
C1711 VDD1.t4 VSUBS 0.272738f
C1712 VDD1.n116 VSUBS 2.09798f
C1713 VDD1.n117 VSUBS 1.4594f
C1714 VDD1.t6 VSUBS 0.272738f
C1715 VDD1.t5 VSUBS 0.272738f
C1716 VDD1.n118 VSUBS 2.13961f
C1717 VDD1.n119 VSUBS 5.019741f
C1718 VDD1.t0 VSUBS 0.272738f
C1719 VDD1.t8 VSUBS 0.272738f
C1720 VDD1.n120 VSUBS 2.09798f
C1721 VDD1.n121 VSUBS 4.96046f
C1722 VP.t4 VSUBS 2.985f
C1723 VP.n0 VSUBS 1.14904f
C1724 VP.n1 VSUBS 0.025894f
C1725 VP.n2 VSUBS 0.05187f
C1726 VP.n3 VSUBS 0.025894f
C1727 VP.n4 VSUBS 0.048502f
C1728 VP.n5 VSUBS 0.025894f
C1729 VP.t9 VSUBS 2.985f
C1730 VP.n6 VSUBS 0.048502f
C1731 VP.n7 VSUBS 0.025894f
C1732 VP.n8 VSUBS 0.048502f
C1733 VP.n9 VSUBS 0.025894f
C1734 VP.t5 VSUBS 2.985f
C1735 VP.n10 VSUBS 0.048502f
C1736 VP.n11 VSUBS 0.025894f
C1737 VP.n12 VSUBS 0.048502f
C1738 VP.n13 VSUBS 0.025894f
C1739 VP.t8 VSUBS 2.985f
C1740 VP.n14 VSUBS 0.048502f
C1741 VP.n15 VSUBS 0.025894f
C1742 VP.n16 VSUBS 0.05187f
C1743 VP.n17 VSUBS 0.025894f
C1744 VP.t2 VSUBS 2.985f
C1745 VP.n18 VSUBS 1.14904f
C1746 VP.t7 VSUBS 2.985f
C1747 VP.n19 VSUBS 1.14904f
C1748 VP.n20 VSUBS 0.025894f
C1749 VP.n21 VSUBS 0.05187f
C1750 VP.n22 VSUBS 0.025894f
C1751 VP.n23 VSUBS 0.048502f
C1752 VP.n24 VSUBS 0.025894f
C1753 VP.t1 VSUBS 2.985f
C1754 VP.n25 VSUBS 0.048502f
C1755 VP.n26 VSUBS 0.025894f
C1756 VP.n27 VSUBS 0.048502f
C1757 VP.n28 VSUBS 0.025894f
C1758 VP.t6 VSUBS 2.985f
C1759 VP.n29 VSUBS 0.048502f
C1760 VP.n30 VSUBS 0.025894f
C1761 VP.n31 VSUBS 0.048502f
C1762 VP.n32 VSUBS 0.33857f
C1763 VP.t0 VSUBS 2.985f
C1764 VP.t3 VSUBS 3.3978f
C1765 VP.n33 VSUBS 1.09517f
C1766 VP.n34 VSUBS 1.14591f
C1767 VP.n35 VSUBS 0.037007f
C1768 VP.n36 VSUBS 0.048502f
C1769 VP.n37 VSUBS 0.025894f
C1770 VP.n38 VSUBS 0.025894f
C1771 VP.n39 VSUBS 0.025894f
C1772 VP.n40 VSUBS 0.046169f
C1773 VP.n41 VSUBS 0.027233f
C1774 VP.n42 VSUBS 0.051031f
C1775 VP.n43 VSUBS 0.025894f
C1776 VP.n44 VSUBS 0.025894f
C1777 VP.n45 VSUBS 0.025894f
C1778 VP.n46 VSUBS 0.048502f
C1779 VP.n47 VSUBS 1.07519f
C1780 VP.n48 VSUBS 0.048502f
C1781 VP.n49 VSUBS 0.025894f
C1782 VP.n50 VSUBS 0.025894f
C1783 VP.n51 VSUBS 0.025894f
C1784 VP.n52 VSUBS 0.051031f
C1785 VP.n53 VSUBS 0.027233f
C1786 VP.n54 VSUBS 0.046169f
C1787 VP.n55 VSUBS 0.025894f
C1788 VP.n56 VSUBS 0.025894f
C1789 VP.n57 VSUBS 0.025894f
C1790 VP.n58 VSUBS 0.048502f
C1791 VP.n59 VSUBS 0.037007f
C1792 VP.n60 VSUBS 1.05063f
C1793 VP.n61 VSUBS 0.03605f
C1794 VP.n62 VSUBS 0.025894f
C1795 VP.n63 VSUBS 0.025894f
C1796 VP.n64 VSUBS 0.025894f
C1797 VP.n65 VSUBS 0.048502f
C1798 VP.n66 VSUBS 0.047248f
C1799 VP.n67 VSUBS 0.025315f
C1800 VP.n68 VSUBS 0.025894f
C1801 VP.n69 VSUBS 0.025894f
C1802 VP.n70 VSUBS 0.025894f
C1803 VP.n71 VSUBS 0.048502f
C1804 VP.n72 VSUBS 0.048502f
C1805 VP.n73 VSUBS 0.025513f
C1806 VP.n74 VSUBS 0.041799f
C1807 VP.n75 VSUBS 1.89573f
C1808 VP.n76 VSUBS 1.91133f
C1809 VP.n77 VSUBS 0.041799f
C1810 VP.n78 VSUBS 0.025513f
C1811 VP.n79 VSUBS 0.048502f
C1812 VP.n80 VSUBS 0.048502f
C1813 VP.n81 VSUBS 0.025894f
C1814 VP.n82 VSUBS 0.025894f
C1815 VP.n83 VSUBS 0.025894f
C1816 VP.n84 VSUBS 0.025315f
C1817 VP.n85 VSUBS 0.047248f
C1818 VP.n86 VSUBS 0.048502f
C1819 VP.n87 VSUBS 0.025894f
C1820 VP.n88 VSUBS 0.025894f
C1821 VP.n89 VSUBS 0.025894f
C1822 VP.n90 VSUBS 0.03605f
C1823 VP.n91 VSUBS 1.05063f
C1824 VP.n92 VSUBS 0.037007f
C1825 VP.n93 VSUBS 0.048502f
C1826 VP.n94 VSUBS 0.025894f
C1827 VP.n95 VSUBS 0.025894f
C1828 VP.n96 VSUBS 0.025894f
C1829 VP.n97 VSUBS 0.046169f
C1830 VP.n98 VSUBS 0.027233f
C1831 VP.n99 VSUBS 0.051031f
C1832 VP.n100 VSUBS 0.025894f
C1833 VP.n101 VSUBS 0.025894f
C1834 VP.n102 VSUBS 0.025894f
C1835 VP.n103 VSUBS 0.048502f
C1836 VP.n104 VSUBS 1.07519f
C1837 VP.n105 VSUBS 0.048502f
C1838 VP.n106 VSUBS 0.025894f
C1839 VP.n107 VSUBS 0.025894f
C1840 VP.n108 VSUBS 0.025894f
C1841 VP.n109 VSUBS 0.051031f
C1842 VP.n110 VSUBS 0.027233f
C1843 VP.n111 VSUBS 0.046169f
C1844 VP.n112 VSUBS 0.025894f
C1845 VP.n113 VSUBS 0.025894f
C1846 VP.n114 VSUBS 0.025894f
C1847 VP.n115 VSUBS 0.048502f
C1848 VP.n116 VSUBS 0.037007f
C1849 VP.n117 VSUBS 1.05063f
C1850 VP.n118 VSUBS 0.03605f
C1851 VP.n119 VSUBS 0.025894f
C1852 VP.n120 VSUBS 0.025894f
C1853 VP.n121 VSUBS 0.025894f
C1854 VP.n122 VSUBS 0.048502f
C1855 VP.n123 VSUBS 0.047248f
C1856 VP.n124 VSUBS 0.025315f
C1857 VP.n125 VSUBS 0.025894f
C1858 VP.n126 VSUBS 0.025894f
C1859 VP.n127 VSUBS 0.025894f
C1860 VP.n128 VSUBS 0.048502f
C1861 VP.n129 VSUBS 0.048502f
C1862 VP.n130 VSUBS 0.025513f
C1863 VP.n131 VSUBS 0.041799f
C1864 VP.n132 VSUBS 0.083019f
.ends

