*
* 4k spice models for n-channel thin oxide mosfets (std VTH). 
*
*
* this scaled model was extracted by coolcad electroncis llc,
* akin akturk, akin.akturk@coolcadelectronics.com
*
* measurements used in model extraction correspond to the 
* following W (um)/L (um) devices:    
*'nshort; w=1.68; l=0.15; m=1';
*'nshort; w=7.0; l=8.0; m=1';
*'nshort; w=7.0; l=0.15; m=1';
*'nshort; w=0.42; l=8.0; m=1';
*'nshort; w=0.42; l=0.15; m=1';
*
* to use the models, please set the circuit temperature
* to -269 in celcius. for standard spice, this can be done 
* by adding the following line to netlist: .options temp=-269
*
* 
*
*
.MODEL nshort NMOS 
+ LEVEL = 54 
+ VERSION = 4.6.5 
+ BINUNIT = 2 
+ PARAMCHK = 1 
+ MOBMOD = 1 
+ MTRLMOD = 0 
+ RDSMOD = 0 
+ IGCMOD = 0 
+ IGBMOD = 0 
+ CVCHARGEMOD = 0 
+ CAPMOD = 2 
+ RGATEMOD = 0 
+ RBODYMOD = 0 
+ TRNQSMOD = 0 
+ ACNQSMOD = 0 
+ FNOIMOD = 1 
+ TNOIMOD = 0 
+ DIOMOD = 1 
+ TEMPMOD = 0 
+ PERMOD = 1 
+ GEOMOD = 0 
+ WPEMOD = 0 
+ EPSROX = 3.9 
+ TOXE = 4.0840E-009 
+ EOT = 4.0840E-009 
+ TOXP = 4.0840E-009 
+ TOXM = 4.0840E-009 
+ DTOX = 0 
+ XJ = 1.5E-007 
+ NDEP = 1.7E+017 
+ NGATE = 1E+022 
+ NSD = 1E+020 
+ XT = 1.55E-007 
+ RSH = 0 
+ RSHG = 0.1 
+ VTH0 = 0.665 
+ WVTH0 = -0.02E-7 
+ LVTH0 = 0.22E-7
+ PVTH0 = 0.08E-14
+ VDDEOT = 1.5 
+ LEFFEOT = 1 
+ WEFFEOT = 10 
+ TEMPEOT = 300.1 
+ PHIN = 0 
+ EASUB = 4.05 
+ EPSRSUB = 11.7 
+ NI0SUB = 1.45E+010 
+ BG0SUB = 1.16 
+ TBGASUB = 0.000702 
+ TBGBSUB = 1108 
+ ADOS = 1 
+ BDOS = 1 
+ VFB = -1 
+ K1 = 0.4
+ K2 = 0.01
+ LK2 = 0.01E-6 
+ PK2 = 0.008E-13
+ K3 = 15 
+ K3B = 0 
+ WK1 = -0.0225E-6
+ LK1 = -0.045E-6
+ PK1 = -0.5E-15 
+ W0 = 9.222E-007 
+ LPE0 = 1.899E-008 
+ LPEB = 6.702E-008 
+ VBM = -3 
+ DVT0 = 0.001
+ DVT1 = 0.1135 
+ DVT2 = -2.864 
+ DVTP0 = 5.919E-009 
+ DVTP1 = 2.966 
+ DVT0W = -10.37 
+ DVT1W = 5.3E+006 
+ DVT2W = -0.032 
+ U0 = 0.25
+ LU0 = -0.036E-6
+ WU0 = -0.02E-6
+ PU0 = 0.01E-12 
+ UA = -1.986E-009 
+ LUA = -5E-0117
+ UB = 0.47E-017 
+ WUB = -2E-025 
+ LUB = -5E-025
+ PUB = 12E-032
+ UC = -0.07076 
+ UD = 3.228 
+ UCS = 1.67 
+ UP = 0.3928 
+ LP = 1.39E-005
+ EU = 1.6 
+ VSAT = 1.8e+004 
+ WVSAT = -1.8E-3
+ LVSAT = 20E-3
+ PVSAT = 1.5e-9
+ A0 = 2.2
+ AGS = 1.4
+ B0 = 0 
+ B1 = 0 
+ KETA = -0.02134 
+ A1 = 0 
+ A2 = 0.8779 
+ WINT = -3.6E-008 
+ LINT = -2.4E-008 
+ DWG = 6.974E-009 
+ LDWG = -5E-015
+ DWB = 0 
+ VOFF = -0.1 
+ VOFFL = 15E-009 
+ MINV = -7
+ LMINV = -15e-7
+ NFACTOR = 2 
+ ETA0 = 2.686 
+ ETAB = -1.412 
+ DSUB = 0.6654 
+ CIT = 0 
+ CDSC = 4.441E-016 
+ CDSCB = -6.337E-006 
+ CDSCD = 0 
+ PCLM = 0.5
+ LPCLM = 0.7E-6
+ WPCLM = -0.1E-6
+ PDIBLC1 = 0.001E-10 
+ PDIBLC2 = 1E-006 
+ PDIBLCB = 0 
+ DROUT = 0.56 
+ PSCBE1 = 1.5E+008 
+ PSCBE2 = 0.15E-006 
+ PVAG = 5 
+ DELTA = 0.01 
+ FPROUT = 0 
+ PDITS = 0.01 
+ PDITSL = 1.392E+006 
+ PDITSD = 1 
+ LAMBDA = 0 
+ VTL = 2E+005 
+ LC = 0 
+ XN = 4 
+ PHIG = 4.05 
+ EPSRGATE = 11.7 
+ RDSW = 0.0 
+ RDSWMIN = 5.0 
+ RDW = 100 
+ RDWMIN = 0 
+ RSW = 100 
+ RSWMIN = 0 
+ PRWG = 0.4 
+ PRWB = -0.1169 
+ WR = 8.882E-016 
+ ALPHA0 = 1E-005 
+ ALPHA1 = 0 
+ BETA0 = 15 
+ AGIDL = 1E-015 
+ BGIDL = 2.3E+009 
+ CGIDL = 0.5 
+ EGIDL = 0.8 
+ AGISL = 0 
+ BGISL = 2.3E+009 
+ CGISL = 0.5 
+ EGISL = 0.8 
+ AIGBACC = 0.43 
+ BIGBACC = 0.054 
+ CIGBACC = 0.075 
+ NIGBACC = 1 
+ AIGBINV = 0.35 
+ BIGBINV = 0.03 
+ CIGBINV = 0.006 
+ EIGBINV = 1.1 
+ NIGBINV = 3 
+ AIGC = 0.54 
+ BIGC = 0.054 
+ CIGC = 0.075 
+ AIGSD = 0.43 
+ BIGSD = 0.054 
+ CIGSD = 0.075 
+ DLCIG = 1.051E-008 
+ AIGS = 0.0136 
+ BIGS = 0.00171 
+ CIGS = 0.075 
+ AIGD = 0.0136 
+ BIGD = 0.00171 
+ CIGD = 0.075 
+ DLCIGD = 0 
+ NIGC = 1 
+ POXEDGE = 1 
+ PIGCD = 1 
+ NTOX = 1 
+ TOXREF = 4.0840E-009 
+ VFBSDOFF = 0 
+ XPART = 0 
+ CGSO = 3E-011 
+ CGDO = 3E-011 
+ CGBO = 0 
+ CGSL = 1.343E-010 
+ CGDL = 1.343E-010 
+ CKAPPAS = 0.6 
+ CKAPPAD = 0.6 
+ CF = 2.977E-010 
+ CLC = 1E-007 
+ CLE = 0.6 
+ DLC = 1.051E-008 
+ DWC = 0 
+ VFBCV = -1 
+ NOFF = 2 
+ VOFFCV = 0.051 
+ VOFFCVL = 0 
+ MINVCV = 0 
+ ACDE = 1 
+ MOIN = 15 
+ XRCRG1 = 12 
+ XRCRG2 = 1 
+ RBPB = 50 
+ RBPD = 50 
+ RBPS = 15 
+ RBDB = 50 
+ RBSB = 50 
+ GBMIN = 1E-012 
+ RBPS0 = 50 
+ RBPSL = 0 
+ RBPSW = 0 
+ RBPSNF = 0 
+ RBPD0 = 50 
+ RBPDL = 0 
+ RBPDW = 0 
+ RBPDNF = 0 
+ RBPBX0 = 100 
+ RBPBXL = 0 
+ RBPBXW = 0 
+ RBPBXNF = 0 
+ RBPBY0 = 100 
+ RBPBYL = 0 
+ RBPBYW = 0 
+ RBPBYNF = 0 
+ RBSBX0 = 100 
+ RBSBY0 = 100 
+ RBDBX0 = 100 
+ RBDBY0 = 100 
+ RBSDBXL = 0 
+ RBSDBXW = 0 
+ RBSDBXNF = 0 
+ RBSDBYL = 0 
+ RBSDBYW = 0 
+ RBSDBYNF = 0 
+ NOIA = 6.25E+041 
+ NOIB = 3.125E+026 
+ NOIC = 8.75 
+ EM = 4.1E+007 
+ AF = 1 
+ EF = 1 
+ KF = 0 
+ LINTNOI = 0 
+ NTNOI = 1 
+ TNOIA = 1.5 
+ TNOIB = 3.5 
+ RNOIA = 0.577 
+ RNOIB = 0.5164 
+ DMCG = 0 
+ DMCI = 0 
+ DMDG = 0 
+ DMCGT = 0 
+ DWJ = 0 
+ XGW = 0 
+ XGL = 0 
+ XL = 0 
+ XW = 5E-8 
+ NGCON = 1 
+ IJTHSREV = 0.0044 
+ IJTHSFWD = 0.0044 
+ XJBVS = 1 
+ BVS = 10 
+ JSS = 1.487E-8 
+ JSWS = 1E-18 
+ JSWGS = 0 
+ JTSS = 0 
+ JTSSWS = 0 
+ JTSSWGS = 0 
+ JTWEFF = 0 
+ NJS = 15 
+ NJTS = 20 
+ NJTSSW = 20 
+ NJTSSWG = 20 
+ XTSS = 0.02 
+ XTSSWS = 0.02 
+ XTSSWGS = 0.02 
+ VTSS = 10 
+ VTSSWS = 10 
+ VTSSWGS = 10 
+ TNJTS = 0 
+ TNJTSSW = 0 
+ TNJTSSWG = 0 
+ CJS = 0.001283 
+ MJS = 0.3296 
+ MJSWS = 0.33 
+ CJSWS = 3.5E-011 
+ CJSWGS = 3.5E-011 
+ MJSWGS = 0.33 
+ PBS = 0.9641 
+ PBSWS = 1 
+ PBSWGS = 1 
+ IJTHDREV = 0.0044 
+ IJTHDFWD = 0.0044 
+ XJBVD = 1 
+ BVD = 10 
+ JSD = 1.487E-8 
+ JSWD = 1E-18 
+ JSWGD = 0 
+ JTSD = 0 
+ JTSSWD = 0 
+ JTSSWGD = 0 
+ NJD = 15 
+ NJTSD = 20 
+ NJTSSWD = 20 
+ NJTSSWGD = 20 
+ XTSD = 0.02 
+ XTSSWD = 0.02 
+ XTSSWGD = 0.02 
+ VTSD = 10 
+ VTSSWD = 10 
+ VTSSWGD = 10 
+ TNJTSD = 0 
+ TNJTSSWD = 0 
+ TNJTSSWGD = 0 
+ CJD = 0.001283 
+ MJD = 0.3296 
+ MJSWD = 0.33 
+ CJSWD = 3.5E-011 
+ CJSWGD = 3.5E-011 
+ MJSWGD = 0.33 
+ PBD = 0.9641 
+ PBSWD = 1 
+ PBSWGD = 1 
+ TNOM = -253 
+ UTE = 0 
+ UCSTE = -0.004775 
+ KT1 = 0 
+ KT1L = 0 
+ KT2 = 0 
+ UA1 = 0 
+ UB1 = 0 
+ UC1 = 0 
+ UD1 = 0 
+ AT = 0 
+ PRT = 0 
+ XTIS = 3 
+ XTID = 3 
+ TPB = 0 
+ TPBSW = 0 
+ TPBSWG = 0 
+ TCJ = 0 
+ TCJSW = 0 
+ TCJSWG = 0 
+ TVOFF = 0 
+ TVFBSDOFF = 0 
+ SAREF = 0 
+ SBREF = 0 
+ WLOD = 2E-006 
+ KU0 = 4E-006 
+ KVSAT = 0.0 
+ TKU0 = 0 
+ LKU0 = 1E-006 
+ WKU0 = 1E-006 
+ PKU0 = 0 
+ LLODKU0 = 1.1 
+ WLODKU0 = 1.1 
+ KVTH0 = -2E-008 
+ LKVTH0 = 1.1E-006 
+ WKVTH0 = 1.1E-006 
+ PKVTH0 = 0 
+ LLODVTH = 1 
+ WLODVTH = 1 
+ STK2 = 0 
+ LODK2 = 1 
+ STETA0 = 0 
+ LODETA0 = 1 
+ WEB = 0 
+ WEC = 0 
+ KVTH0WE = 0 
+ K2WE = 0 
+ KU0WE = 0 
+ SCREF = 1E-006 
+ WL = 1E-014 
+ WLN = 1.056 
+ WW = 10.807E-015 
+ WWN = 1.03 
+ WWL = -1.419E-021 
+ LL = -1.609E-015 
+ LLN = 0.9 
+ LW = -7.92E-015 
+ LWN = 1.012 
+ LWL = 6.569E-021 
+ LLC = 0 
+ LWC = 0 
+ LWLC = 0 
+ WLC = 0 
+ WWC = 0 
+ WWLC = 0 
*
*
