* NGSPICE file created from diff_pair_sample_1014.ext - technology: sky130A

.subckt diff_pair_sample_1014 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=2.28195 ps=14.16 w=13.83 l=3.2
X1 VTAIL.t7 VP.t0 VDD1.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X2 VDD1.t8 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=5.3937 ps=28.44 w=13.83 l=3.2
X3 VDD1.t7 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=5.3937 ps=28.44 w=13.83 l=3.2
X4 VTAIL.t4 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X5 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=0 ps=0 w=13.83 l=3.2
X6 VDD1.t5 VP.t4 VTAIL.t18 B.t22 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X7 VDD2.t8 VN.t1 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=2.28195 ps=14.16 w=13.83 l=3.2
X8 VTAIL.t16 VN.t2 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X9 VTAIL.t8 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X10 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=0 ps=0 w=13.83 l=3.2
X11 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=0 ps=0 w=13.83 l=3.2
X12 VTAIL.t13 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X13 VTAIL.t3 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X14 VTAIL.t9 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X15 VDD2.t3 VN.t6 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=5.3937 ps=28.44 w=13.83 l=3.2
X16 VDD2.t2 VN.t7 VTAIL.t10 B.t23 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X17 VDD1.t3 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=2.28195 ps=14.16 w=13.83 l=3.2
X18 VDD1.t2 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=2.28195 ps=14.16 w=13.83 l=3.2
X19 VDD2.t1 VN.t8 VTAIL.t17 B.t22 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X20 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
X21 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3937 pd=28.44 as=0 ps=0 w=13.83 l=3.2
X22 VDD2.t0 VN.t9 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=5.3937 ps=28.44 w=13.83 l=3.2
X23 VDD1.t0 VP.t9 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=2.28195 pd=14.16 as=2.28195 ps=14.16 w=13.83 l=3.2
R0 VN.n94 VN.n93 161.3
R1 VN.n92 VN.n49 161.3
R2 VN.n91 VN.n90 161.3
R3 VN.n89 VN.n50 161.3
R4 VN.n88 VN.n87 161.3
R5 VN.n86 VN.n51 161.3
R6 VN.n85 VN.n84 161.3
R7 VN.n83 VN.n82 161.3
R8 VN.n81 VN.n53 161.3
R9 VN.n80 VN.n79 161.3
R10 VN.n78 VN.n54 161.3
R11 VN.n77 VN.n76 161.3
R12 VN.n75 VN.n55 161.3
R13 VN.n74 VN.n73 161.3
R14 VN.n72 VN.n71 161.3
R15 VN.n70 VN.n57 161.3
R16 VN.n69 VN.n68 161.3
R17 VN.n67 VN.n58 161.3
R18 VN.n66 VN.n65 161.3
R19 VN.n64 VN.n59 161.3
R20 VN.n63 VN.n62 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n1 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n2 161.3
R25 VN.n40 VN.n39 161.3
R26 VN.n38 VN.n3 161.3
R27 VN.n37 VN.n36 161.3
R28 VN.n35 VN.n34 161.3
R29 VN.n33 VN.n5 161.3
R30 VN.n32 VN.n31 161.3
R31 VN.n30 VN.n6 161.3
R32 VN.n29 VN.n28 161.3
R33 VN.n27 VN.n7 161.3
R34 VN.n26 VN.n25 161.3
R35 VN.n24 VN.n23 161.3
R36 VN.n22 VN.n9 161.3
R37 VN.n21 VN.n20 161.3
R38 VN.n19 VN.n10 161.3
R39 VN.n18 VN.n17 161.3
R40 VN.n16 VN.n11 161.3
R41 VN.n15 VN.n14 161.3
R42 VN.n61 VN.t6 137.179
R43 VN.n13 VN.t0 137.179
R44 VN.n12 VN.t4 104.157
R45 VN.n8 VN.t8 104.157
R46 VN.n4 VN.t3 104.157
R47 VN.n0 VN.t9 104.157
R48 VN.n60 VN.t5 104.157
R49 VN.n56 VN.t7 104.157
R50 VN.n52 VN.t2 104.157
R51 VN.n48 VN.t1 104.157
R52 VN.n47 VN.n0 74.8979
R53 VN.n95 VN.n48 74.8979
R54 VN.n13 VN.n12 60.5137
R55 VN.n61 VN.n60 60.5137
R56 VN VN.n95 58.0245
R57 VN.n43 VN.n2 44.8641
R58 VN.n91 VN.n50 44.8641
R59 VN.n17 VN.n10 41.9503
R60 VN.n32 VN.n6 41.9503
R61 VN.n65 VN.n58 41.9503
R62 VN.n80 VN.n54 41.9503
R63 VN.n21 VN.n10 39.0365
R64 VN.n28 VN.n6 39.0365
R65 VN.n69 VN.n58 39.0365
R66 VN.n76 VN.n54 39.0365
R67 VN.n39 VN.n2 36.1227
R68 VN.n87 VN.n50 36.1227
R69 VN.n16 VN.n15 24.4675
R70 VN.n17 VN.n16 24.4675
R71 VN.n22 VN.n21 24.4675
R72 VN.n23 VN.n22 24.4675
R73 VN.n27 VN.n26 24.4675
R74 VN.n28 VN.n27 24.4675
R75 VN.n33 VN.n32 24.4675
R76 VN.n34 VN.n33 24.4675
R77 VN.n38 VN.n37 24.4675
R78 VN.n39 VN.n38 24.4675
R79 VN.n44 VN.n43 24.4675
R80 VN.n45 VN.n44 24.4675
R81 VN.n65 VN.n64 24.4675
R82 VN.n64 VN.n63 24.4675
R83 VN.n76 VN.n75 24.4675
R84 VN.n75 VN.n74 24.4675
R85 VN.n71 VN.n70 24.4675
R86 VN.n70 VN.n69 24.4675
R87 VN.n87 VN.n86 24.4675
R88 VN.n86 VN.n85 24.4675
R89 VN.n82 VN.n81 24.4675
R90 VN.n81 VN.n80 24.4675
R91 VN.n93 VN.n92 24.4675
R92 VN.n92 VN.n91 24.4675
R93 VN.n45 VN.n0 15.17
R94 VN.n93 VN.n48 15.17
R95 VN.n15 VN.n12 13.702
R96 VN.n34 VN.n4 13.702
R97 VN.n63 VN.n60 13.702
R98 VN.n82 VN.n52 13.702
R99 VN.n23 VN.n8 12.234
R100 VN.n26 VN.n8 12.234
R101 VN.n74 VN.n56 12.234
R102 VN.n71 VN.n56 12.234
R103 VN.n37 VN.n4 10.766
R104 VN.n85 VN.n52 10.766
R105 VN.n62 VN.n61 4.13481
R106 VN.n14 VN.n13 4.13481
R107 VN.n95 VN.n94 0.354971
R108 VN.n47 VN.n46 0.354971
R109 VN VN.n47 0.26696
R110 VN.n94 VN.n49 0.189894
R111 VN.n90 VN.n49 0.189894
R112 VN.n90 VN.n89 0.189894
R113 VN.n89 VN.n88 0.189894
R114 VN.n88 VN.n51 0.189894
R115 VN.n84 VN.n51 0.189894
R116 VN.n84 VN.n83 0.189894
R117 VN.n83 VN.n53 0.189894
R118 VN.n79 VN.n53 0.189894
R119 VN.n79 VN.n78 0.189894
R120 VN.n78 VN.n77 0.189894
R121 VN.n77 VN.n55 0.189894
R122 VN.n73 VN.n55 0.189894
R123 VN.n73 VN.n72 0.189894
R124 VN.n72 VN.n57 0.189894
R125 VN.n68 VN.n57 0.189894
R126 VN.n68 VN.n67 0.189894
R127 VN.n67 VN.n66 0.189894
R128 VN.n66 VN.n59 0.189894
R129 VN.n62 VN.n59 0.189894
R130 VN.n14 VN.n11 0.189894
R131 VN.n18 VN.n11 0.189894
R132 VN.n19 VN.n18 0.189894
R133 VN.n20 VN.n19 0.189894
R134 VN.n20 VN.n9 0.189894
R135 VN.n24 VN.n9 0.189894
R136 VN.n25 VN.n24 0.189894
R137 VN.n25 VN.n7 0.189894
R138 VN.n29 VN.n7 0.189894
R139 VN.n30 VN.n29 0.189894
R140 VN.n31 VN.n30 0.189894
R141 VN.n31 VN.n5 0.189894
R142 VN.n35 VN.n5 0.189894
R143 VN.n36 VN.n35 0.189894
R144 VN.n36 VN.n3 0.189894
R145 VN.n40 VN.n3 0.189894
R146 VN.n41 VN.n40 0.189894
R147 VN.n42 VN.n41 0.189894
R148 VN.n42 VN.n1 0.189894
R149 VN.n46 VN.n1 0.189894
R150 VTAIL.n16 VTAIL.t6 44.4957
R151 VTAIL.n11 VTAIL.t14 44.4957
R152 VTAIL.n17 VTAIL.t15 44.4956
R153 VTAIL.n2 VTAIL.t5 44.4956
R154 VTAIL.n15 VTAIL.n14 43.0641
R155 VTAIL.n13 VTAIL.n12 43.0641
R156 VTAIL.n10 VTAIL.n9 43.0641
R157 VTAIL.n8 VTAIL.n7 43.0641
R158 VTAIL.n19 VTAIL.n18 43.064
R159 VTAIL.n1 VTAIL.n0 43.064
R160 VTAIL.n4 VTAIL.n3 43.064
R161 VTAIL.n6 VTAIL.n5 43.064
R162 VTAIL.n8 VTAIL.n6 30.3755
R163 VTAIL.n17 VTAIL.n16 27.3324
R164 VTAIL.n10 VTAIL.n8 3.0436
R165 VTAIL.n11 VTAIL.n10 3.0436
R166 VTAIL.n15 VTAIL.n13 3.0436
R167 VTAIL.n16 VTAIL.n15 3.0436
R168 VTAIL.n6 VTAIL.n4 3.0436
R169 VTAIL.n4 VTAIL.n2 3.0436
R170 VTAIL.n19 VTAIL.n17 3.0436
R171 VTAIL VTAIL.n1 2.34102
R172 VTAIL.n13 VTAIL.n11 1.99188
R173 VTAIL.n2 VTAIL.n1 1.99188
R174 VTAIL.n18 VTAIL.t17 1.43217
R175 VTAIL.n18 VTAIL.t8 1.43217
R176 VTAIL.n0 VTAIL.t11 1.43217
R177 VTAIL.n0 VTAIL.t13 1.43217
R178 VTAIL.n3 VTAIL.t19 1.43217
R179 VTAIL.n3 VTAIL.t1 1.43217
R180 VTAIL.n5 VTAIL.t2 1.43217
R181 VTAIL.n5 VTAIL.t7 1.43217
R182 VTAIL.n14 VTAIL.t18 1.43217
R183 VTAIL.n14 VTAIL.t4 1.43217
R184 VTAIL.n12 VTAIL.t0 1.43217
R185 VTAIL.n12 VTAIL.t3 1.43217
R186 VTAIL.n9 VTAIL.t10 1.43217
R187 VTAIL.n9 VTAIL.t9 1.43217
R188 VTAIL.n7 VTAIL.t12 1.43217
R189 VTAIL.n7 VTAIL.t16 1.43217
R190 VTAIL VTAIL.n19 0.703086
R191 VDD2.n1 VDD2.t9 64.2174
R192 VDD2.n3 VDD2.n2 61.9698
R193 VDD2 VDD2.n7 61.967
R194 VDD2.n4 VDD2.t8 61.1745
R195 VDD2.n6 VDD2.n5 59.7429
R196 VDD2.n1 VDD2.n0 59.7428
R197 VDD2.n4 VDD2.n3 50.0924
R198 VDD2.n6 VDD2.n4 3.0436
R199 VDD2.n7 VDD2.t4 1.43217
R200 VDD2.n7 VDD2.t3 1.43217
R201 VDD2.n5 VDD2.t7 1.43217
R202 VDD2.n5 VDD2.t2 1.43217
R203 VDD2.n2 VDD2.t6 1.43217
R204 VDD2.n2 VDD2.t0 1.43217
R205 VDD2.n0 VDD2.t5 1.43217
R206 VDD2.n0 VDD2.t1 1.43217
R207 VDD2 VDD2.n6 0.819465
R208 VDD2.n3 VDD2.n1 0.70593
R209 B.n890 B.n889 585
R210 B.n892 B.n185 585
R211 B.n895 B.n894 585
R212 B.n896 B.n184 585
R213 B.n898 B.n897 585
R214 B.n900 B.n183 585
R215 B.n903 B.n902 585
R216 B.n904 B.n182 585
R217 B.n906 B.n905 585
R218 B.n908 B.n181 585
R219 B.n911 B.n910 585
R220 B.n912 B.n180 585
R221 B.n914 B.n913 585
R222 B.n916 B.n179 585
R223 B.n919 B.n918 585
R224 B.n920 B.n178 585
R225 B.n922 B.n921 585
R226 B.n924 B.n177 585
R227 B.n927 B.n926 585
R228 B.n928 B.n176 585
R229 B.n930 B.n929 585
R230 B.n932 B.n175 585
R231 B.n935 B.n934 585
R232 B.n936 B.n174 585
R233 B.n938 B.n937 585
R234 B.n940 B.n173 585
R235 B.n943 B.n942 585
R236 B.n944 B.n172 585
R237 B.n946 B.n945 585
R238 B.n948 B.n171 585
R239 B.n951 B.n950 585
R240 B.n952 B.n170 585
R241 B.n954 B.n953 585
R242 B.n956 B.n169 585
R243 B.n959 B.n958 585
R244 B.n960 B.n168 585
R245 B.n962 B.n961 585
R246 B.n964 B.n167 585
R247 B.n967 B.n966 585
R248 B.n968 B.n166 585
R249 B.n970 B.n969 585
R250 B.n972 B.n165 585
R251 B.n975 B.n974 585
R252 B.n976 B.n164 585
R253 B.n978 B.n977 585
R254 B.n980 B.n163 585
R255 B.n983 B.n982 585
R256 B.n985 B.n160 585
R257 B.n987 B.n986 585
R258 B.n989 B.n159 585
R259 B.n992 B.n991 585
R260 B.n993 B.n158 585
R261 B.n995 B.n994 585
R262 B.n997 B.n157 585
R263 B.n1000 B.n999 585
R264 B.n1001 B.n153 585
R265 B.n1003 B.n1002 585
R266 B.n1005 B.n152 585
R267 B.n1008 B.n1007 585
R268 B.n1009 B.n151 585
R269 B.n1011 B.n1010 585
R270 B.n1013 B.n150 585
R271 B.n1016 B.n1015 585
R272 B.n1017 B.n149 585
R273 B.n1019 B.n1018 585
R274 B.n1021 B.n148 585
R275 B.n1024 B.n1023 585
R276 B.n1025 B.n147 585
R277 B.n1027 B.n1026 585
R278 B.n1029 B.n146 585
R279 B.n1032 B.n1031 585
R280 B.n1033 B.n145 585
R281 B.n1035 B.n1034 585
R282 B.n1037 B.n144 585
R283 B.n1040 B.n1039 585
R284 B.n1041 B.n143 585
R285 B.n1043 B.n1042 585
R286 B.n1045 B.n142 585
R287 B.n1048 B.n1047 585
R288 B.n1049 B.n141 585
R289 B.n1051 B.n1050 585
R290 B.n1053 B.n140 585
R291 B.n1056 B.n1055 585
R292 B.n1057 B.n139 585
R293 B.n1059 B.n1058 585
R294 B.n1061 B.n138 585
R295 B.n1064 B.n1063 585
R296 B.n1065 B.n137 585
R297 B.n1067 B.n1066 585
R298 B.n1069 B.n136 585
R299 B.n1072 B.n1071 585
R300 B.n1073 B.n135 585
R301 B.n1075 B.n1074 585
R302 B.n1077 B.n134 585
R303 B.n1080 B.n1079 585
R304 B.n1081 B.n133 585
R305 B.n1083 B.n1082 585
R306 B.n1085 B.n132 585
R307 B.n1088 B.n1087 585
R308 B.n1089 B.n131 585
R309 B.n1091 B.n1090 585
R310 B.n1093 B.n130 585
R311 B.n1096 B.n1095 585
R312 B.n1097 B.n129 585
R313 B.n888 B.n127 585
R314 B.n1100 B.n127 585
R315 B.n887 B.n126 585
R316 B.n1101 B.n126 585
R317 B.n886 B.n125 585
R318 B.n1102 B.n125 585
R319 B.n885 B.n884 585
R320 B.n884 B.n121 585
R321 B.n883 B.n120 585
R322 B.n1108 B.n120 585
R323 B.n882 B.n119 585
R324 B.n1109 B.n119 585
R325 B.n881 B.n118 585
R326 B.n1110 B.n118 585
R327 B.n880 B.n879 585
R328 B.n879 B.n114 585
R329 B.n878 B.n113 585
R330 B.n1116 B.n113 585
R331 B.n877 B.n112 585
R332 B.n1117 B.n112 585
R333 B.n876 B.n111 585
R334 B.n1118 B.n111 585
R335 B.n875 B.n874 585
R336 B.n874 B.n107 585
R337 B.n873 B.n106 585
R338 B.n1124 B.n106 585
R339 B.n872 B.n105 585
R340 B.n1125 B.n105 585
R341 B.n871 B.n104 585
R342 B.n1126 B.n104 585
R343 B.n870 B.n869 585
R344 B.n869 B.n100 585
R345 B.n868 B.n99 585
R346 B.n1132 B.n99 585
R347 B.n867 B.n98 585
R348 B.n1133 B.n98 585
R349 B.n866 B.n97 585
R350 B.n1134 B.n97 585
R351 B.n865 B.n864 585
R352 B.n864 B.n93 585
R353 B.n863 B.n92 585
R354 B.n1140 B.n92 585
R355 B.n862 B.n91 585
R356 B.n1141 B.n91 585
R357 B.n861 B.n90 585
R358 B.n1142 B.n90 585
R359 B.n860 B.n859 585
R360 B.n859 B.n86 585
R361 B.n858 B.n85 585
R362 B.n1148 B.n85 585
R363 B.n857 B.n84 585
R364 B.n1149 B.n84 585
R365 B.n856 B.n83 585
R366 B.n1150 B.n83 585
R367 B.n855 B.n854 585
R368 B.n854 B.n79 585
R369 B.n853 B.n78 585
R370 B.n1156 B.n78 585
R371 B.n852 B.n77 585
R372 B.n1157 B.n77 585
R373 B.n851 B.n76 585
R374 B.n1158 B.n76 585
R375 B.n850 B.n849 585
R376 B.n849 B.n72 585
R377 B.n848 B.n71 585
R378 B.n1164 B.n71 585
R379 B.n847 B.n70 585
R380 B.n1165 B.n70 585
R381 B.n846 B.n69 585
R382 B.n1166 B.n69 585
R383 B.n845 B.n844 585
R384 B.n844 B.n65 585
R385 B.n843 B.n64 585
R386 B.n1172 B.n64 585
R387 B.n842 B.n63 585
R388 B.n1173 B.n63 585
R389 B.n841 B.n62 585
R390 B.n1174 B.n62 585
R391 B.n840 B.n839 585
R392 B.n839 B.n58 585
R393 B.n838 B.n57 585
R394 B.n1180 B.n57 585
R395 B.n837 B.n56 585
R396 B.n1181 B.n56 585
R397 B.n836 B.n55 585
R398 B.n1182 B.n55 585
R399 B.n835 B.n834 585
R400 B.n834 B.n51 585
R401 B.n833 B.n50 585
R402 B.n1188 B.n50 585
R403 B.n832 B.n49 585
R404 B.n1189 B.n49 585
R405 B.n831 B.n48 585
R406 B.n1190 B.n48 585
R407 B.n830 B.n829 585
R408 B.n829 B.n44 585
R409 B.n828 B.n43 585
R410 B.n1196 B.n43 585
R411 B.n827 B.n42 585
R412 B.n1197 B.n42 585
R413 B.n826 B.n41 585
R414 B.n1198 B.n41 585
R415 B.n825 B.n824 585
R416 B.n824 B.n37 585
R417 B.n823 B.n36 585
R418 B.n1204 B.n36 585
R419 B.n822 B.n35 585
R420 B.n1205 B.n35 585
R421 B.n821 B.n34 585
R422 B.n1206 B.n34 585
R423 B.n820 B.n819 585
R424 B.n819 B.n30 585
R425 B.n818 B.n29 585
R426 B.n1212 B.n29 585
R427 B.n817 B.n28 585
R428 B.n1213 B.n28 585
R429 B.n816 B.n27 585
R430 B.n1214 B.n27 585
R431 B.n815 B.n814 585
R432 B.n814 B.n23 585
R433 B.n813 B.n22 585
R434 B.n1220 B.n22 585
R435 B.n812 B.n21 585
R436 B.n1221 B.n21 585
R437 B.n811 B.n20 585
R438 B.n1222 B.n20 585
R439 B.n810 B.n809 585
R440 B.n809 B.n19 585
R441 B.n808 B.n15 585
R442 B.n1228 B.n15 585
R443 B.n807 B.n14 585
R444 B.n1229 B.n14 585
R445 B.n806 B.n13 585
R446 B.n1230 B.n13 585
R447 B.n805 B.n804 585
R448 B.n804 B.n12 585
R449 B.n803 B.n802 585
R450 B.n803 B.n8 585
R451 B.n801 B.n7 585
R452 B.n1237 B.n7 585
R453 B.n800 B.n6 585
R454 B.n1238 B.n6 585
R455 B.n799 B.n5 585
R456 B.n1239 B.n5 585
R457 B.n798 B.n797 585
R458 B.n797 B.n4 585
R459 B.n796 B.n186 585
R460 B.n796 B.n795 585
R461 B.n786 B.n187 585
R462 B.n188 B.n187 585
R463 B.n788 B.n787 585
R464 B.n789 B.n788 585
R465 B.n785 B.n193 585
R466 B.n193 B.n192 585
R467 B.n784 B.n783 585
R468 B.n783 B.n782 585
R469 B.n195 B.n194 585
R470 B.n775 B.n195 585
R471 B.n774 B.n773 585
R472 B.n776 B.n774 585
R473 B.n772 B.n200 585
R474 B.n200 B.n199 585
R475 B.n771 B.n770 585
R476 B.n770 B.n769 585
R477 B.n202 B.n201 585
R478 B.n203 B.n202 585
R479 B.n762 B.n761 585
R480 B.n763 B.n762 585
R481 B.n760 B.n208 585
R482 B.n208 B.n207 585
R483 B.n759 B.n758 585
R484 B.n758 B.n757 585
R485 B.n210 B.n209 585
R486 B.n211 B.n210 585
R487 B.n750 B.n749 585
R488 B.n751 B.n750 585
R489 B.n748 B.n215 585
R490 B.n219 B.n215 585
R491 B.n747 B.n746 585
R492 B.n746 B.n745 585
R493 B.n217 B.n216 585
R494 B.n218 B.n217 585
R495 B.n738 B.n737 585
R496 B.n739 B.n738 585
R497 B.n736 B.n224 585
R498 B.n224 B.n223 585
R499 B.n735 B.n734 585
R500 B.n734 B.n733 585
R501 B.n226 B.n225 585
R502 B.n227 B.n226 585
R503 B.n726 B.n725 585
R504 B.n727 B.n726 585
R505 B.n724 B.n232 585
R506 B.n232 B.n231 585
R507 B.n723 B.n722 585
R508 B.n722 B.n721 585
R509 B.n234 B.n233 585
R510 B.n235 B.n234 585
R511 B.n714 B.n713 585
R512 B.n715 B.n714 585
R513 B.n712 B.n240 585
R514 B.n240 B.n239 585
R515 B.n711 B.n710 585
R516 B.n710 B.n709 585
R517 B.n242 B.n241 585
R518 B.n243 B.n242 585
R519 B.n702 B.n701 585
R520 B.n703 B.n702 585
R521 B.n700 B.n248 585
R522 B.n248 B.n247 585
R523 B.n699 B.n698 585
R524 B.n698 B.n697 585
R525 B.n250 B.n249 585
R526 B.n251 B.n250 585
R527 B.n690 B.n689 585
R528 B.n691 B.n690 585
R529 B.n688 B.n256 585
R530 B.n256 B.n255 585
R531 B.n687 B.n686 585
R532 B.n686 B.n685 585
R533 B.n258 B.n257 585
R534 B.n259 B.n258 585
R535 B.n678 B.n677 585
R536 B.n679 B.n678 585
R537 B.n676 B.n264 585
R538 B.n264 B.n263 585
R539 B.n675 B.n674 585
R540 B.n674 B.n673 585
R541 B.n266 B.n265 585
R542 B.n267 B.n266 585
R543 B.n666 B.n665 585
R544 B.n667 B.n666 585
R545 B.n664 B.n272 585
R546 B.n272 B.n271 585
R547 B.n663 B.n662 585
R548 B.n662 B.n661 585
R549 B.n274 B.n273 585
R550 B.n275 B.n274 585
R551 B.n654 B.n653 585
R552 B.n655 B.n654 585
R553 B.n652 B.n280 585
R554 B.n280 B.n279 585
R555 B.n651 B.n650 585
R556 B.n650 B.n649 585
R557 B.n282 B.n281 585
R558 B.n283 B.n282 585
R559 B.n642 B.n641 585
R560 B.n643 B.n642 585
R561 B.n640 B.n288 585
R562 B.n288 B.n287 585
R563 B.n639 B.n638 585
R564 B.n638 B.n637 585
R565 B.n290 B.n289 585
R566 B.n291 B.n290 585
R567 B.n630 B.n629 585
R568 B.n631 B.n630 585
R569 B.n628 B.n296 585
R570 B.n296 B.n295 585
R571 B.n627 B.n626 585
R572 B.n626 B.n625 585
R573 B.n298 B.n297 585
R574 B.n299 B.n298 585
R575 B.n618 B.n617 585
R576 B.n619 B.n618 585
R577 B.n616 B.n304 585
R578 B.n304 B.n303 585
R579 B.n615 B.n614 585
R580 B.n614 B.n613 585
R581 B.n306 B.n305 585
R582 B.n307 B.n306 585
R583 B.n606 B.n605 585
R584 B.n607 B.n606 585
R585 B.n604 B.n312 585
R586 B.n312 B.n311 585
R587 B.n603 B.n602 585
R588 B.n602 B.n601 585
R589 B.n314 B.n313 585
R590 B.n315 B.n314 585
R591 B.n594 B.n593 585
R592 B.n595 B.n594 585
R593 B.n592 B.n320 585
R594 B.n320 B.n319 585
R595 B.n591 B.n590 585
R596 B.n590 B.n589 585
R597 B.n586 B.n324 585
R598 B.n585 B.n584 585
R599 B.n582 B.n325 585
R600 B.n582 B.n323 585
R601 B.n581 B.n580 585
R602 B.n579 B.n578 585
R603 B.n577 B.n327 585
R604 B.n575 B.n574 585
R605 B.n573 B.n328 585
R606 B.n572 B.n571 585
R607 B.n569 B.n329 585
R608 B.n567 B.n566 585
R609 B.n565 B.n330 585
R610 B.n564 B.n563 585
R611 B.n561 B.n331 585
R612 B.n559 B.n558 585
R613 B.n557 B.n332 585
R614 B.n556 B.n555 585
R615 B.n553 B.n333 585
R616 B.n551 B.n550 585
R617 B.n549 B.n334 585
R618 B.n548 B.n547 585
R619 B.n545 B.n335 585
R620 B.n543 B.n542 585
R621 B.n541 B.n336 585
R622 B.n540 B.n539 585
R623 B.n537 B.n337 585
R624 B.n535 B.n534 585
R625 B.n533 B.n338 585
R626 B.n532 B.n531 585
R627 B.n529 B.n339 585
R628 B.n527 B.n526 585
R629 B.n525 B.n340 585
R630 B.n524 B.n523 585
R631 B.n521 B.n341 585
R632 B.n519 B.n518 585
R633 B.n517 B.n342 585
R634 B.n516 B.n515 585
R635 B.n513 B.n343 585
R636 B.n511 B.n510 585
R637 B.n509 B.n344 585
R638 B.n508 B.n507 585
R639 B.n505 B.n345 585
R640 B.n503 B.n502 585
R641 B.n501 B.n346 585
R642 B.n500 B.n499 585
R643 B.n497 B.n347 585
R644 B.n495 B.n494 585
R645 B.n492 B.n348 585
R646 B.n491 B.n490 585
R647 B.n488 B.n351 585
R648 B.n486 B.n485 585
R649 B.n484 B.n352 585
R650 B.n483 B.n482 585
R651 B.n480 B.n353 585
R652 B.n478 B.n477 585
R653 B.n476 B.n354 585
R654 B.n475 B.n474 585
R655 B.n472 B.n471 585
R656 B.n470 B.n469 585
R657 B.n468 B.n359 585
R658 B.n466 B.n465 585
R659 B.n464 B.n360 585
R660 B.n463 B.n462 585
R661 B.n460 B.n361 585
R662 B.n458 B.n457 585
R663 B.n456 B.n362 585
R664 B.n455 B.n454 585
R665 B.n452 B.n363 585
R666 B.n450 B.n449 585
R667 B.n448 B.n364 585
R668 B.n447 B.n446 585
R669 B.n444 B.n365 585
R670 B.n442 B.n441 585
R671 B.n440 B.n366 585
R672 B.n439 B.n438 585
R673 B.n436 B.n367 585
R674 B.n434 B.n433 585
R675 B.n432 B.n368 585
R676 B.n431 B.n430 585
R677 B.n428 B.n369 585
R678 B.n426 B.n425 585
R679 B.n424 B.n370 585
R680 B.n423 B.n422 585
R681 B.n420 B.n371 585
R682 B.n418 B.n417 585
R683 B.n416 B.n372 585
R684 B.n415 B.n414 585
R685 B.n412 B.n373 585
R686 B.n410 B.n409 585
R687 B.n408 B.n374 585
R688 B.n407 B.n406 585
R689 B.n404 B.n375 585
R690 B.n402 B.n401 585
R691 B.n400 B.n376 585
R692 B.n399 B.n398 585
R693 B.n396 B.n377 585
R694 B.n394 B.n393 585
R695 B.n392 B.n378 585
R696 B.n391 B.n390 585
R697 B.n388 B.n379 585
R698 B.n386 B.n385 585
R699 B.n384 B.n380 585
R700 B.n383 B.n382 585
R701 B.n322 B.n321 585
R702 B.n323 B.n322 585
R703 B.n588 B.n587 585
R704 B.n589 B.n588 585
R705 B.n318 B.n317 585
R706 B.n319 B.n318 585
R707 B.n597 B.n596 585
R708 B.n596 B.n595 585
R709 B.n598 B.n316 585
R710 B.n316 B.n315 585
R711 B.n600 B.n599 585
R712 B.n601 B.n600 585
R713 B.n310 B.n309 585
R714 B.n311 B.n310 585
R715 B.n609 B.n608 585
R716 B.n608 B.n607 585
R717 B.n610 B.n308 585
R718 B.n308 B.n307 585
R719 B.n612 B.n611 585
R720 B.n613 B.n612 585
R721 B.n302 B.n301 585
R722 B.n303 B.n302 585
R723 B.n621 B.n620 585
R724 B.n620 B.n619 585
R725 B.n622 B.n300 585
R726 B.n300 B.n299 585
R727 B.n624 B.n623 585
R728 B.n625 B.n624 585
R729 B.n294 B.n293 585
R730 B.n295 B.n294 585
R731 B.n633 B.n632 585
R732 B.n632 B.n631 585
R733 B.n634 B.n292 585
R734 B.n292 B.n291 585
R735 B.n636 B.n635 585
R736 B.n637 B.n636 585
R737 B.n286 B.n285 585
R738 B.n287 B.n286 585
R739 B.n645 B.n644 585
R740 B.n644 B.n643 585
R741 B.n646 B.n284 585
R742 B.n284 B.n283 585
R743 B.n648 B.n647 585
R744 B.n649 B.n648 585
R745 B.n278 B.n277 585
R746 B.n279 B.n278 585
R747 B.n657 B.n656 585
R748 B.n656 B.n655 585
R749 B.n658 B.n276 585
R750 B.n276 B.n275 585
R751 B.n660 B.n659 585
R752 B.n661 B.n660 585
R753 B.n270 B.n269 585
R754 B.n271 B.n270 585
R755 B.n669 B.n668 585
R756 B.n668 B.n667 585
R757 B.n670 B.n268 585
R758 B.n268 B.n267 585
R759 B.n672 B.n671 585
R760 B.n673 B.n672 585
R761 B.n262 B.n261 585
R762 B.n263 B.n262 585
R763 B.n681 B.n680 585
R764 B.n680 B.n679 585
R765 B.n682 B.n260 585
R766 B.n260 B.n259 585
R767 B.n684 B.n683 585
R768 B.n685 B.n684 585
R769 B.n254 B.n253 585
R770 B.n255 B.n254 585
R771 B.n693 B.n692 585
R772 B.n692 B.n691 585
R773 B.n694 B.n252 585
R774 B.n252 B.n251 585
R775 B.n696 B.n695 585
R776 B.n697 B.n696 585
R777 B.n246 B.n245 585
R778 B.n247 B.n246 585
R779 B.n705 B.n704 585
R780 B.n704 B.n703 585
R781 B.n706 B.n244 585
R782 B.n244 B.n243 585
R783 B.n708 B.n707 585
R784 B.n709 B.n708 585
R785 B.n238 B.n237 585
R786 B.n239 B.n238 585
R787 B.n717 B.n716 585
R788 B.n716 B.n715 585
R789 B.n718 B.n236 585
R790 B.n236 B.n235 585
R791 B.n720 B.n719 585
R792 B.n721 B.n720 585
R793 B.n230 B.n229 585
R794 B.n231 B.n230 585
R795 B.n729 B.n728 585
R796 B.n728 B.n727 585
R797 B.n730 B.n228 585
R798 B.n228 B.n227 585
R799 B.n732 B.n731 585
R800 B.n733 B.n732 585
R801 B.n222 B.n221 585
R802 B.n223 B.n222 585
R803 B.n741 B.n740 585
R804 B.n740 B.n739 585
R805 B.n742 B.n220 585
R806 B.n220 B.n218 585
R807 B.n744 B.n743 585
R808 B.n745 B.n744 585
R809 B.n214 B.n213 585
R810 B.n219 B.n214 585
R811 B.n753 B.n752 585
R812 B.n752 B.n751 585
R813 B.n754 B.n212 585
R814 B.n212 B.n211 585
R815 B.n756 B.n755 585
R816 B.n757 B.n756 585
R817 B.n206 B.n205 585
R818 B.n207 B.n206 585
R819 B.n765 B.n764 585
R820 B.n764 B.n763 585
R821 B.n766 B.n204 585
R822 B.n204 B.n203 585
R823 B.n768 B.n767 585
R824 B.n769 B.n768 585
R825 B.n198 B.n197 585
R826 B.n199 B.n198 585
R827 B.n778 B.n777 585
R828 B.n777 B.n776 585
R829 B.n779 B.n196 585
R830 B.n775 B.n196 585
R831 B.n781 B.n780 585
R832 B.n782 B.n781 585
R833 B.n191 B.n190 585
R834 B.n192 B.n191 585
R835 B.n791 B.n790 585
R836 B.n790 B.n789 585
R837 B.n792 B.n189 585
R838 B.n189 B.n188 585
R839 B.n794 B.n793 585
R840 B.n795 B.n794 585
R841 B.n3 B.n0 585
R842 B.n4 B.n3 585
R843 B.n1236 B.n1 585
R844 B.n1237 B.n1236 585
R845 B.n1235 B.n1234 585
R846 B.n1235 B.n8 585
R847 B.n1233 B.n9 585
R848 B.n12 B.n9 585
R849 B.n1232 B.n1231 585
R850 B.n1231 B.n1230 585
R851 B.n11 B.n10 585
R852 B.n1229 B.n11 585
R853 B.n1227 B.n1226 585
R854 B.n1228 B.n1227 585
R855 B.n1225 B.n16 585
R856 B.n19 B.n16 585
R857 B.n1224 B.n1223 585
R858 B.n1223 B.n1222 585
R859 B.n18 B.n17 585
R860 B.n1221 B.n18 585
R861 B.n1219 B.n1218 585
R862 B.n1220 B.n1219 585
R863 B.n1217 B.n24 585
R864 B.n24 B.n23 585
R865 B.n1216 B.n1215 585
R866 B.n1215 B.n1214 585
R867 B.n26 B.n25 585
R868 B.n1213 B.n26 585
R869 B.n1211 B.n1210 585
R870 B.n1212 B.n1211 585
R871 B.n1209 B.n31 585
R872 B.n31 B.n30 585
R873 B.n1208 B.n1207 585
R874 B.n1207 B.n1206 585
R875 B.n33 B.n32 585
R876 B.n1205 B.n33 585
R877 B.n1203 B.n1202 585
R878 B.n1204 B.n1203 585
R879 B.n1201 B.n38 585
R880 B.n38 B.n37 585
R881 B.n1200 B.n1199 585
R882 B.n1199 B.n1198 585
R883 B.n40 B.n39 585
R884 B.n1197 B.n40 585
R885 B.n1195 B.n1194 585
R886 B.n1196 B.n1195 585
R887 B.n1193 B.n45 585
R888 B.n45 B.n44 585
R889 B.n1192 B.n1191 585
R890 B.n1191 B.n1190 585
R891 B.n47 B.n46 585
R892 B.n1189 B.n47 585
R893 B.n1187 B.n1186 585
R894 B.n1188 B.n1187 585
R895 B.n1185 B.n52 585
R896 B.n52 B.n51 585
R897 B.n1184 B.n1183 585
R898 B.n1183 B.n1182 585
R899 B.n54 B.n53 585
R900 B.n1181 B.n54 585
R901 B.n1179 B.n1178 585
R902 B.n1180 B.n1179 585
R903 B.n1177 B.n59 585
R904 B.n59 B.n58 585
R905 B.n1176 B.n1175 585
R906 B.n1175 B.n1174 585
R907 B.n61 B.n60 585
R908 B.n1173 B.n61 585
R909 B.n1171 B.n1170 585
R910 B.n1172 B.n1171 585
R911 B.n1169 B.n66 585
R912 B.n66 B.n65 585
R913 B.n1168 B.n1167 585
R914 B.n1167 B.n1166 585
R915 B.n68 B.n67 585
R916 B.n1165 B.n68 585
R917 B.n1163 B.n1162 585
R918 B.n1164 B.n1163 585
R919 B.n1161 B.n73 585
R920 B.n73 B.n72 585
R921 B.n1160 B.n1159 585
R922 B.n1159 B.n1158 585
R923 B.n75 B.n74 585
R924 B.n1157 B.n75 585
R925 B.n1155 B.n1154 585
R926 B.n1156 B.n1155 585
R927 B.n1153 B.n80 585
R928 B.n80 B.n79 585
R929 B.n1152 B.n1151 585
R930 B.n1151 B.n1150 585
R931 B.n82 B.n81 585
R932 B.n1149 B.n82 585
R933 B.n1147 B.n1146 585
R934 B.n1148 B.n1147 585
R935 B.n1145 B.n87 585
R936 B.n87 B.n86 585
R937 B.n1144 B.n1143 585
R938 B.n1143 B.n1142 585
R939 B.n89 B.n88 585
R940 B.n1141 B.n89 585
R941 B.n1139 B.n1138 585
R942 B.n1140 B.n1139 585
R943 B.n1137 B.n94 585
R944 B.n94 B.n93 585
R945 B.n1136 B.n1135 585
R946 B.n1135 B.n1134 585
R947 B.n96 B.n95 585
R948 B.n1133 B.n96 585
R949 B.n1131 B.n1130 585
R950 B.n1132 B.n1131 585
R951 B.n1129 B.n101 585
R952 B.n101 B.n100 585
R953 B.n1128 B.n1127 585
R954 B.n1127 B.n1126 585
R955 B.n103 B.n102 585
R956 B.n1125 B.n103 585
R957 B.n1123 B.n1122 585
R958 B.n1124 B.n1123 585
R959 B.n1121 B.n108 585
R960 B.n108 B.n107 585
R961 B.n1120 B.n1119 585
R962 B.n1119 B.n1118 585
R963 B.n110 B.n109 585
R964 B.n1117 B.n110 585
R965 B.n1115 B.n1114 585
R966 B.n1116 B.n1115 585
R967 B.n1113 B.n115 585
R968 B.n115 B.n114 585
R969 B.n1112 B.n1111 585
R970 B.n1111 B.n1110 585
R971 B.n117 B.n116 585
R972 B.n1109 B.n117 585
R973 B.n1107 B.n1106 585
R974 B.n1108 B.n1107 585
R975 B.n1105 B.n122 585
R976 B.n122 B.n121 585
R977 B.n1104 B.n1103 585
R978 B.n1103 B.n1102 585
R979 B.n124 B.n123 585
R980 B.n1101 B.n124 585
R981 B.n1099 B.n1098 585
R982 B.n1100 B.n1099 585
R983 B.n1240 B.n1239 585
R984 B.n1238 B.n2 585
R985 B.n1099 B.n129 449.257
R986 B.n890 B.n127 449.257
R987 B.n590 B.n322 449.257
R988 B.n588 B.n324 449.257
R989 B.n154 B.t15 312.959
R990 B.n161 B.t19 312.959
R991 B.n355 B.t8 312.959
R992 B.n349 B.t12 312.959
R993 B.n891 B.n128 256.663
R994 B.n893 B.n128 256.663
R995 B.n899 B.n128 256.663
R996 B.n901 B.n128 256.663
R997 B.n907 B.n128 256.663
R998 B.n909 B.n128 256.663
R999 B.n915 B.n128 256.663
R1000 B.n917 B.n128 256.663
R1001 B.n923 B.n128 256.663
R1002 B.n925 B.n128 256.663
R1003 B.n931 B.n128 256.663
R1004 B.n933 B.n128 256.663
R1005 B.n939 B.n128 256.663
R1006 B.n941 B.n128 256.663
R1007 B.n947 B.n128 256.663
R1008 B.n949 B.n128 256.663
R1009 B.n955 B.n128 256.663
R1010 B.n957 B.n128 256.663
R1011 B.n963 B.n128 256.663
R1012 B.n965 B.n128 256.663
R1013 B.n971 B.n128 256.663
R1014 B.n973 B.n128 256.663
R1015 B.n979 B.n128 256.663
R1016 B.n981 B.n128 256.663
R1017 B.n988 B.n128 256.663
R1018 B.n990 B.n128 256.663
R1019 B.n996 B.n128 256.663
R1020 B.n998 B.n128 256.663
R1021 B.n1004 B.n128 256.663
R1022 B.n1006 B.n128 256.663
R1023 B.n1012 B.n128 256.663
R1024 B.n1014 B.n128 256.663
R1025 B.n1020 B.n128 256.663
R1026 B.n1022 B.n128 256.663
R1027 B.n1028 B.n128 256.663
R1028 B.n1030 B.n128 256.663
R1029 B.n1036 B.n128 256.663
R1030 B.n1038 B.n128 256.663
R1031 B.n1044 B.n128 256.663
R1032 B.n1046 B.n128 256.663
R1033 B.n1052 B.n128 256.663
R1034 B.n1054 B.n128 256.663
R1035 B.n1060 B.n128 256.663
R1036 B.n1062 B.n128 256.663
R1037 B.n1068 B.n128 256.663
R1038 B.n1070 B.n128 256.663
R1039 B.n1076 B.n128 256.663
R1040 B.n1078 B.n128 256.663
R1041 B.n1084 B.n128 256.663
R1042 B.n1086 B.n128 256.663
R1043 B.n1092 B.n128 256.663
R1044 B.n1094 B.n128 256.663
R1045 B.n583 B.n323 256.663
R1046 B.n326 B.n323 256.663
R1047 B.n576 B.n323 256.663
R1048 B.n570 B.n323 256.663
R1049 B.n568 B.n323 256.663
R1050 B.n562 B.n323 256.663
R1051 B.n560 B.n323 256.663
R1052 B.n554 B.n323 256.663
R1053 B.n552 B.n323 256.663
R1054 B.n546 B.n323 256.663
R1055 B.n544 B.n323 256.663
R1056 B.n538 B.n323 256.663
R1057 B.n536 B.n323 256.663
R1058 B.n530 B.n323 256.663
R1059 B.n528 B.n323 256.663
R1060 B.n522 B.n323 256.663
R1061 B.n520 B.n323 256.663
R1062 B.n514 B.n323 256.663
R1063 B.n512 B.n323 256.663
R1064 B.n506 B.n323 256.663
R1065 B.n504 B.n323 256.663
R1066 B.n498 B.n323 256.663
R1067 B.n496 B.n323 256.663
R1068 B.n489 B.n323 256.663
R1069 B.n487 B.n323 256.663
R1070 B.n481 B.n323 256.663
R1071 B.n479 B.n323 256.663
R1072 B.n473 B.n323 256.663
R1073 B.n358 B.n323 256.663
R1074 B.n467 B.n323 256.663
R1075 B.n461 B.n323 256.663
R1076 B.n459 B.n323 256.663
R1077 B.n453 B.n323 256.663
R1078 B.n451 B.n323 256.663
R1079 B.n445 B.n323 256.663
R1080 B.n443 B.n323 256.663
R1081 B.n437 B.n323 256.663
R1082 B.n435 B.n323 256.663
R1083 B.n429 B.n323 256.663
R1084 B.n427 B.n323 256.663
R1085 B.n421 B.n323 256.663
R1086 B.n419 B.n323 256.663
R1087 B.n413 B.n323 256.663
R1088 B.n411 B.n323 256.663
R1089 B.n405 B.n323 256.663
R1090 B.n403 B.n323 256.663
R1091 B.n397 B.n323 256.663
R1092 B.n395 B.n323 256.663
R1093 B.n389 B.n323 256.663
R1094 B.n387 B.n323 256.663
R1095 B.n381 B.n323 256.663
R1096 B.n1242 B.n1241 256.663
R1097 B.n1095 B.n1093 163.367
R1098 B.n1091 B.n131 163.367
R1099 B.n1087 B.n1085 163.367
R1100 B.n1083 B.n133 163.367
R1101 B.n1079 B.n1077 163.367
R1102 B.n1075 B.n135 163.367
R1103 B.n1071 B.n1069 163.367
R1104 B.n1067 B.n137 163.367
R1105 B.n1063 B.n1061 163.367
R1106 B.n1059 B.n139 163.367
R1107 B.n1055 B.n1053 163.367
R1108 B.n1051 B.n141 163.367
R1109 B.n1047 B.n1045 163.367
R1110 B.n1043 B.n143 163.367
R1111 B.n1039 B.n1037 163.367
R1112 B.n1035 B.n145 163.367
R1113 B.n1031 B.n1029 163.367
R1114 B.n1027 B.n147 163.367
R1115 B.n1023 B.n1021 163.367
R1116 B.n1019 B.n149 163.367
R1117 B.n1015 B.n1013 163.367
R1118 B.n1011 B.n151 163.367
R1119 B.n1007 B.n1005 163.367
R1120 B.n1003 B.n153 163.367
R1121 B.n999 B.n997 163.367
R1122 B.n995 B.n158 163.367
R1123 B.n991 B.n989 163.367
R1124 B.n987 B.n160 163.367
R1125 B.n982 B.n980 163.367
R1126 B.n978 B.n164 163.367
R1127 B.n974 B.n972 163.367
R1128 B.n970 B.n166 163.367
R1129 B.n966 B.n964 163.367
R1130 B.n962 B.n168 163.367
R1131 B.n958 B.n956 163.367
R1132 B.n954 B.n170 163.367
R1133 B.n950 B.n948 163.367
R1134 B.n946 B.n172 163.367
R1135 B.n942 B.n940 163.367
R1136 B.n938 B.n174 163.367
R1137 B.n934 B.n932 163.367
R1138 B.n930 B.n176 163.367
R1139 B.n926 B.n924 163.367
R1140 B.n922 B.n178 163.367
R1141 B.n918 B.n916 163.367
R1142 B.n914 B.n180 163.367
R1143 B.n910 B.n908 163.367
R1144 B.n906 B.n182 163.367
R1145 B.n902 B.n900 163.367
R1146 B.n898 B.n184 163.367
R1147 B.n894 B.n892 163.367
R1148 B.n590 B.n320 163.367
R1149 B.n594 B.n320 163.367
R1150 B.n594 B.n314 163.367
R1151 B.n602 B.n314 163.367
R1152 B.n602 B.n312 163.367
R1153 B.n606 B.n312 163.367
R1154 B.n606 B.n306 163.367
R1155 B.n614 B.n306 163.367
R1156 B.n614 B.n304 163.367
R1157 B.n618 B.n304 163.367
R1158 B.n618 B.n298 163.367
R1159 B.n626 B.n298 163.367
R1160 B.n626 B.n296 163.367
R1161 B.n630 B.n296 163.367
R1162 B.n630 B.n290 163.367
R1163 B.n638 B.n290 163.367
R1164 B.n638 B.n288 163.367
R1165 B.n642 B.n288 163.367
R1166 B.n642 B.n282 163.367
R1167 B.n650 B.n282 163.367
R1168 B.n650 B.n280 163.367
R1169 B.n654 B.n280 163.367
R1170 B.n654 B.n274 163.367
R1171 B.n662 B.n274 163.367
R1172 B.n662 B.n272 163.367
R1173 B.n666 B.n272 163.367
R1174 B.n666 B.n266 163.367
R1175 B.n674 B.n266 163.367
R1176 B.n674 B.n264 163.367
R1177 B.n678 B.n264 163.367
R1178 B.n678 B.n258 163.367
R1179 B.n686 B.n258 163.367
R1180 B.n686 B.n256 163.367
R1181 B.n690 B.n256 163.367
R1182 B.n690 B.n250 163.367
R1183 B.n698 B.n250 163.367
R1184 B.n698 B.n248 163.367
R1185 B.n702 B.n248 163.367
R1186 B.n702 B.n242 163.367
R1187 B.n710 B.n242 163.367
R1188 B.n710 B.n240 163.367
R1189 B.n714 B.n240 163.367
R1190 B.n714 B.n234 163.367
R1191 B.n722 B.n234 163.367
R1192 B.n722 B.n232 163.367
R1193 B.n726 B.n232 163.367
R1194 B.n726 B.n226 163.367
R1195 B.n734 B.n226 163.367
R1196 B.n734 B.n224 163.367
R1197 B.n738 B.n224 163.367
R1198 B.n738 B.n217 163.367
R1199 B.n746 B.n217 163.367
R1200 B.n746 B.n215 163.367
R1201 B.n750 B.n215 163.367
R1202 B.n750 B.n210 163.367
R1203 B.n758 B.n210 163.367
R1204 B.n758 B.n208 163.367
R1205 B.n762 B.n208 163.367
R1206 B.n762 B.n202 163.367
R1207 B.n770 B.n202 163.367
R1208 B.n770 B.n200 163.367
R1209 B.n774 B.n200 163.367
R1210 B.n774 B.n195 163.367
R1211 B.n783 B.n195 163.367
R1212 B.n783 B.n193 163.367
R1213 B.n788 B.n193 163.367
R1214 B.n788 B.n187 163.367
R1215 B.n796 B.n187 163.367
R1216 B.n797 B.n796 163.367
R1217 B.n797 B.n5 163.367
R1218 B.n6 B.n5 163.367
R1219 B.n7 B.n6 163.367
R1220 B.n803 B.n7 163.367
R1221 B.n804 B.n803 163.367
R1222 B.n804 B.n13 163.367
R1223 B.n14 B.n13 163.367
R1224 B.n15 B.n14 163.367
R1225 B.n809 B.n15 163.367
R1226 B.n809 B.n20 163.367
R1227 B.n21 B.n20 163.367
R1228 B.n22 B.n21 163.367
R1229 B.n814 B.n22 163.367
R1230 B.n814 B.n27 163.367
R1231 B.n28 B.n27 163.367
R1232 B.n29 B.n28 163.367
R1233 B.n819 B.n29 163.367
R1234 B.n819 B.n34 163.367
R1235 B.n35 B.n34 163.367
R1236 B.n36 B.n35 163.367
R1237 B.n824 B.n36 163.367
R1238 B.n824 B.n41 163.367
R1239 B.n42 B.n41 163.367
R1240 B.n43 B.n42 163.367
R1241 B.n829 B.n43 163.367
R1242 B.n829 B.n48 163.367
R1243 B.n49 B.n48 163.367
R1244 B.n50 B.n49 163.367
R1245 B.n834 B.n50 163.367
R1246 B.n834 B.n55 163.367
R1247 B.n56 B.n55 163.367
R1248 B.n57 B.n56 163.367
R1249 B.n839 B.n57 163.367
R1250 B.n839 B.n62 163.367
R1251 B.n63 B.n62 163.367
R1252 B.n64 B.n63 163.367
R1253 B.n844 B.n64 163.367
R1254 B.n844 B.n69 163.367
R1255 B.n70 B.n69 163.367
R1256 B.n71 B.n70 163.367
R1257 B.n849 B.n71 163.367
R1258 B.n849 B.n76 163.367
R1259 B.n77 B.n76 163.367
R1260 B.n78 B.n77 163.367
R1261 B.n854 B.n78 163.367
R1262 B.n854 B.n83 163.367
R1263 B.n84 B.n83 163.367
R1264 B.n85 B.n84 163.367
R1265 B.n859 B.n85 163.367
R1266 B.n859 B.n90 163.367
R1267 B.n91 B.n90 163.367
R1268 B.n92 B.n91 163.367
R1269 B.n864 B.n92 163.367
R1270 B.n864 B.n97 163.367
R1271 B.n98 B.n97 163.367
R1272 B.n99 B.n98 163.367
R1273 B.n869 B.n99 163.367
R1274 B.n869 B.n104 163.367
R1275 B.n105 B.n104 163.367
R1276 B.n106 B.n105 163.367
R1277 B.n874 B.n106 163.367
R1278 B.n874 B.n111 163.367
R1279 B.n112 B.n111 163.367
R1280 B.n113 B.n112 163.367
R1281 B.n879 B.n113 163.367
R1282 B.n879 B.n118 163.367
R1283 B.n119 B.n118 163.367
R1284 B.n120 B.n119 163.367
R1285 B.n884 B.n120 163.367
R1286 B.n884 B.n125 163.367
R1287 B.n126 B.n125 163.367
R1288 B.n127 B.n126 163.367
R1289 B.n584 B.n582 163.367
R1290 B.n582 B.n581 163.367
R1291 B.n578 B.n577 163.367
R1292 B.n575 B.n328 163.367
R1293 B.n571 B.n569 163.367
R1294 B.n567 B.n330 163.367
R1295 B.n563 B.n561 163.367
R1296 B.n559 B.n332 163.367
R1297 B.n555 B.n553 163.367
R1298 B.n551 B.n334 163.367
R1299 B.n547 B.n545 163.367
R1300 B.n543 B.n336 163.367
R1301 B.n539 B.n537 163.367
R1302 B.n535 B.n338 163.367
R1303 B.n531 B.n529 163.367
R1304 B.n527 B.n340 163.367
R1305 B.n523 B.n521 163.367
R1306 B.n519 B.n342 163.367
R1307 B.n515 B.n513 163.367
R1308 B.n511 B.n344 163.367
R1309 B.n507 B.n505 163.367
R1310 B.n503 B.n346 163.367
R1311 B.n499 B.n497 163.367
R1312 B.n495 B.n348 163.367
R1313 B.n490 B.n488 163.367
R1314 B.n486 B.n352 163.367
R1315 B.n482 B.n480 163.367
R1316 B.n478 B.n354 163.367
R1317 B.n474 B.n472 163.367
R1318 B.n469 B.n468 163.367
R1319 B.n466 B.n360 163.367
R1320 B.n462 B.n460 163.367
R1321 B.n458 B.n362 163.367
R1322 B.n454 B.n452 163.367
R1323 B.n450 B.n364 163.367
R1324 B.n446 B.n444 163.367
R1325 B.n442 B.n366 163.367
R1326 B.n438 B.n436 163.367
R1327 B.n434 B.n368 163.367
R1328 B.n430 B.n428 163.367
R1329 B.n426 B.n370 163.367
R1330 B.n422 B.n420 163.367
R1331 B.n418 B.n372 163.367
R1332 B.n414 B.n412 163.367
R1333 B.n410 B.n374 163.367
R1334 B.n406 B.n404 163.367
R1335 B.n402 B.n376 163.367
R1336 B.n398 B.n396 163.367
R1337 B.n394 B.n378 163.367
R1338 B.n390 B.n388 163.367
R1339 B.n386 B.n380 163.367
R1340 B.n382 B.n322 163.367
R1341 B.n588 B.n318 163.367
R1342 B.n596 B.n318 163.367
R1343 B.n596 B.n316 163.367
R1344 B.n600 B.n316 163.367
R1345 B.n600 B.n310 163.367
R1346 B.n608 B.n310 163.367
R1347 B.n608 B.n308 163.367
R1348 B.n612 B.n308 163.367
R1349 B.n612 B.n302 163.367
R1350 B.n620 B.n302 163.367
R1351 B.n620 B.n300 163.367
R1352 B.n624 B.n300 163.367
R1353 B.n624 B.n294 163.367
R1354 B.n632 B.n294 163.367
R1355 B.n632 B.n292 163.367
R1356 B.n636 B.n292 163.367
R1357 B.n636 B.n286 163.367
R1358 B.n644 B.n286 163.367
R1359 B.n644 B.n284 163.367
R1360 B.n648 B.n284 163.367
R1361 B.n648 B.n278 163.367
R1362 B.n656 B.n278 163.367
R1363 B.n656 B.n276 163.367
R1364 B.n660 B.n276 163.367
R1365 B.n660 B.n270 163.367
R1366 B.n668 B.n270 163.367
R1367 B.n668 B.n268 163.367
R1368 B.n672 B.n268 163.367
R1369 B.n672 B.n262 163.367
R1370 B.n680 B.n262 163.367
R1371 B.n680 B.n260 163.367
R1372 B.n684 B.n260 163.367
R1373 B.n684 B.n254 163.367
R1374 B.n692 B.n254 163.367
R1375 B.n692 B.n252 163.367
R1376 B.n696 B.n252 163.367
R1377 B.n696 B.n246 163.367
R1378 B.n704 B.n246 163.367
R1379 B.n704 B.n244 163.367
R1380 B.n708 B.n244 163.367
R1381 B.n708 B.n238 163.367
R1382 B.n716 B.n238 163.367
R1383 B.n716 B.n236 163.367
R1384 B.n720 B.n236 163.367
R1385 B.n720 B.n230 163.367
R1386 B.n728 B.n230 163.367
R1387 B.n728 B.n228 163.367
R1388 B.n732 B.n228 163.367
R1389 B.n732 B.n222 163.367
R1390 B.n740 B.n222 163.367
R1391 B.n740 B.n220 163.367
R1392 B.n744 B.n220 163.367
R1393 B.n744 B.n214 163.367
R1394 B.n752 B.n214 163.367
R1395 B.n752 B.n212 163.367
R1396 B.n756 B.n212 163.367
R1397 B.n756 B.n206 163.367
R1398 B.n764 B.n206 163.367
R1399 B.n764 B.n204 163.367
R1400 B.n768 B.n204 163.367
R1401 B.n768 B.n198 163.367
R1402 B.n777 B.n198 163.367
R1403 B.n777 B.n196 163.367
R1404 B.n781 B.n196 163.367
R1405 B.n781 B.n191 163.367
R1406 B.n790 B.n191 163.367
R1407 B.n790 B.n189 163.367
R1408 B.n794 B.n189 163.367
R1409 B.n794 B.n3 163.367
R1410 B.n1240 B.n3 163.367
R1411 B.n1236 B.n2 163.367
R1412 B.n1236 B.n1235 163.367
R1413 B.n1235 B.n9 163.367
R1414 B.n1231 B.n9 163.367
R1415 B.n1231 B.n11 163.367
R1416 B.n1227 B.n11 163.367
R1417 B.n1227 B.n16 163.367
R1418 B.n1223 B.n16 163.367
R1419 B.n1223 B.n18 163.367
R1420 B.n1219 B.n18 163.367
R1421 B.n1219 B.n24 163.367
R1422 B.n1215 B.n24 163.367
R1423 B.n1215 B.n26 163.367
R1424 B.n1211 B.n26 163.367
R1425 B.n1211 B.n31 163.367
R1426 B.n1207 B.n31 163.367
R1427 B.n1207 B.n33 163.367
R1428 B.n1203 B.n33 163.367
R1429 B.n1203 B.n38 163.367
R1430 B.n1199 B.n38 163.367
R1431 B.n1199 B.n40 163.367
R1432 B.n1195 B.n40 163.367
R1433 B.n1195 B.n45 163.367
R1434 B.n1191 B.n45 163.367
R1435 B.n1191 B.n47 163.367
R1436 B.n1187 B.n47 163.367
R1437 B.n1187 B.n52 163.367
R1438 B.n1183 B.n52 163.367
R1439 B.n1183 B.n54 163.367
R1440 B.n1179 B.n54 163.367
R1441 B.n1179 B.n59 163.367
R1442 B.n1175 B.n59 163.367
R1443 B.n1175 B.n61 163.367
R1444 B.n1171 B.n61 163.367
R1445 B.n1171 B.n66 163.367
R1446 B.n1167 B.n66 163.367
R1447 B.n1167 B.n68 163.367
R1448 B.n1163 B.n68 163.367
R1449 B.n1163 B.n73 163.367
R1450 B.n1159 B.n73 163.367
R1451 B.n1159 B.n75 163.367
R1452 B.n1155 B.n75 163.367
R1453 B.n1155 B.n80 163.367
R1454 B.n1151 B.n80 163.367
R1455 B.n1151 B.n82 163.367
R1456 B.n1147 B.n82 163.367
R1457 B.n1147 B.n87 163.367
R1458 B.n1143 B.n87 163.367
R1459 B.n1143 B.n89 163.367
R1460 B.n1139 B.n89 163.367
R1461 B.n1139 B.n94 163.367
R1462 B.n1135 B.n94 163.367
R1463 B.n1135 B.n96 163.367
R1464 B.n1131 B.n96 163.367
R1465 B.n1131 B.n101 163.367
R1466 B.n1127 B.n101 163.367
R1467 B.n1127 B.n103 163.367
R1468 B.n1123 B.n103 163.367
R1469 B.n1123 B.n108 163.367
R1470 B.n1119 B.n108 163.367
R1471 B.n1119 B.n110 163.367
R1472 B.n1115 B.n110 163.367
R1473 B.n1115 B.n115 163.367
R1474 B.n1111 B.n115 163.367
R1475 B.n1111 B.n117 163.367
R1476 B.n1107 B.n117 163.367
R1477 B.n1107 B.n122 163.367
R1478 B.n1103 B.n122 163.367
R1479 B.n1103 B.n124 163.367
R1480 B.n1099 B.n124 163.367
R1481 B.n161 B.t20 140.495
R1482 B.n355 B.t11 140.495
R1483 B.n154 B.t17 140.477
R1484 B.n349 B.t14 140.477
R1485 B.n162 B.t21 72.0347
R1486 B.n356 B.t10 72.0347
R1487 B.n155 B.t18 72.0169
R1488 B.n350 B.t13 72.0169
R1489 B.n1094 B.n129 71.676
R1490 B.n1093 B.n1092 71.676
R1491 B.n1086 B.n131 71.676
R1492 B.n1085 B.n1084 71.676
R1493 B.n1078 B.n133 71.676
R1494 B.n1077 B.n1076 71.676
R1495 B.n1070 B.n135 71.676
R1496 B.n1069 B.n1068 71.676
R1497 B.n1062 B.n137 71.676
R1498 B.n1061 B.n1060 71.676
R1499 B.n1054 B.n139 71.676
R1500 B.n1053 B.n1052 71.676
R1501 B.n1046 B.n141 71.676
R1502 B.n1045 B.n1044 71.676
R1503 B.n1038 B.n143 71.676
R1504 B.n1037 B.n1036 71.676
R1505 B.n1030 B.n145 71.676
R1506 B.n1029 B.n1028 71.676
R1507 B.n1022 B.n147 71.676
R1508 B.n1021 B.n1020 71.676
R1509 B.n1014 B.n149 71.676
R1510 B.n1013 B.n1012 71.676
R1511 B.n1006 B.n151 71.676
R1512 B.n1005 B.n1004 71.676
R1513 B.n998 B.n153 71.676
R1514 B.n997 B.n996 71.676
R1515 B.n990 B.n158 71.676
R1516 B.n989 B.n988 71.676
R1517 B.n981 B.n160 71.676
R1518 B.n980 B.n979 71.676
R1519 B.n973 B.n164 71.676
R1520 B.n972 B.n971 71.676
R1521 B.n965 B.n166 71.676
R1522 B.n964 B.n963 71.676
R1523 B.n957 B.n168 71.676
R1524 B.n956 B.n955 71.676
R1525 B.n949 B.n170 71.676
R1526 B.n948 B.n947 71.676
R1527 B.n941 B.n172 71.676
R1528 B.n940 B.n939 71.676
R1529 B.n933 B.n174 71.676
R1530 B.n932 B.n931 71.676
R1531 B.n925 B.n176 71.676
R1532 B.n924 B.n923 71.676
R1533 B.n917 B.n178 71.676
R1534 B.n916 B.n915 71.676
R1535 B.n909 B.n180 71.676
R1536 B.n908 B.n907 71.676
R1537 B.n901 B.n182 71.676
R1538 B.n900 B.n899 71.676
R1539 B.n893 B.n184 71.676
R1540 B.n892 B.n891 71.676
R1541 B.n891 B.n890 71.676
R1542 B.n894 B.n893 71.676
R1543 B.n899 B.n898 71.676
R1544 B.n902 B.n901 71.676
R1545 B.n907 B.n906 71.676
R1546 B.n910 B.n909 71.676
R1547 B.n915 B.n914 71.676
R1548 B.n918 B.n917 71.676
R1549 B.n923 B.n922 71.676
R1550 B.n926 B.n925 71.676
R1551 B.n931 B.n930 71.676
R1552 B.n934 B.n933 71.676
R1553 B.n939 B.n938 71.676
R1554 B.n942 B.n941 71.676
R1555 B.n947 B.n946 71.676
R1556 B.n950 B.n949 71.676
R1557 B.n955 B.n954 71.676
R1558 B.n958 B.n957 71.676
R1559 B.n963 B.n962 71.676
R1560 B.n966 B.n965 71.676
R1561 B.n971 B.n970 71.676
R1562 B.n974 B.n973 71.676
R1563 B.n979 B.n978 71.676
R1564 B.n982 B.n981 71.676
R1565 B.n988 B.n987 71.676
R1566 B.n991 B.n990 71.676
R1567 B.n996 B.n995 71.676
R1568 B.n999 B.n998 71.676
R1569 B.n1004 B.n1003 71.676
R1570 B.n1007 B.n1006 71.676
R1571 B.n1012 B.n1011 71.676
R1572 B.n1015 B.n1014 71.676
R1573 B.n1020 B.n1019 71.676
R1574 B.n1023 B.n1022 71.676
R1575 B.n1028 B.n1027 71.676
R1576 B.n1031 B.n1030 71.676
R1577 B.n1036 B.n1035 71.676
R1578 B.n1039 B.n1038 71.676
R1579 B.n1044 B.n1043 71.676
R1580 B.n1047 B.n1046 71.676
R1581 B.n1052 B.n1051 71.676
R1582 B.n1055 B.n1054 71.676
R1583 B.n1060 B.n1059 71.676
R1584 B.n1063 B.n1062 71.676
R1585 B.n1068 B.n1067 71.676
R1586 B.n1071 B.n1070 71.676
R1587 B.n1076 B.n1075 71.676
R1588 B.n1079 B.n1078 71.676
R1589 B.n1084 B.n1083 71.676
R1590 B.n1087 B.n1086 71.676
R1591 B.n1092 B.n1091 71.676
R1592 B.n1095 B.n1094 71.676
R1593 B.n583 B.n324 71.676
R1594 B.n581 B.n326 71.676
R1595 B.n577 B.n576 71.676
R1596 B.n570 B.n328 71.676
R1597 B.n569 B.n568 71.676
R1598 B.n562 B.n330 71.676
R1599 B.n561 B.n560 71.676
R1600 B.n554 B.n332 71.676
R1601 B.n553 B.n552 71.676
R1602 B.n546 B.n334 71.676
R1603 B.n545 B.n544 71.676
R1604 B.n538 B.n336 71.676
R1605 B.n537 B.n536 71.676
R1606 B.n530 B.n338 71.676
R1607 B.n529 B.n528 71.676
R1608 B.n522 B.n340 71.676
R1609 B.n521 B.n520 71.676
R1610 B.n514 B.n342 71.676
R1611 B.n513 B.n512 71.676
R1612 B.n506 B.n344 71.676
R1613 B.n505 B.n504 71.676
R1614 B.n498 B.n346 71.676
R1615 B.n497 B.n496 71.676
R1616 B.n489 B.n348 71.676
R1617 B.n488 B.n487 71.676
R1618 B.n481 B.n352 71.676
R1619 B.n480 B.n479 71.676
R1620 B.n473 B.n354 71.676
R1621 B.n472 B.n358 71.676
R1622 B.n468 B.n467 71.676
R1623 B.n461 B.n360 71.676
R1624 B.n460 B.n459 71.676
R1625 B.n453 B.n362 71.676
R1626 B.n452 B.n451 71.676
R1627 B.n445 B.n364 71.676
R1628 B.n444 B.n443 71.676
R1629 B.n437 B.n366 71.676
R1630 B.n436 B.n435 71.676
R1631 B.n429 B.n368 71.676
R1632 B.n428 B.n427 71.676
R1633 B.n421 B.n370 71.676
R1634 B.n420 B.n419 71.676
R1635 B.n413 B.n372 71.676
R1636 B.n412 B.n411 71.676
R1637 B.n405 B.n374 71.676
R1638 B.n404 B.n403 71.676
R1639 B.n397 B.n376 71.676
R1640 B.n396 B.n395 71.676
R1641 B.n389 B.n378 71.676
R1642 B.n388 B.n387 71.676
R1643 B.n381 B.n380 71.676
R1644 B.n584 B.n583 71.676
R1645 B.n578 B.n326 71.676
R1646 B.n576 B.n575 71.676
R1647 B.n571 B.n570 71.676
R1648 B.n568 B.n567 71.676
R1649 B.n563 B.n562 71.676
R1650 B.n560 B.n559 71.676
R1651 B.n555 B.n554 71.676
R1652 B.n552 B.n551 71.676
R1653 B.n547 B.n546 71.676
R1654 B.n544 B.n543 71.676
R1655 B.n539 B.n538 71.676
R1656 B.n536 B.n535 71.676
R1657 B.n531 B.n530 71.676
R1658 B.n528 B.n527 71.676
R1659 B.n523 B.n522 71.676
R1660 B.n520 B.n519 71.676
R1661 B.n515 B.n514 71.676
R1662 B.n512 B.n511 71.676
R1663 B.n507 B.n506 71.676
R1664 B.n504 B.n503 71.676
R1665 B.n499 B.n498 71.676
R1666 B.n496 B.n495 71.676
R1667 B.n490 B.n489 71.676
R1668 B.n487 B.n486 71.676
R1669 B.n482 B.n481 71.676
R1670 B.n479 B.n478 71.676
R1671 B.n474 B.n473 71.676
R1672 B.n469 B.n358 71.676
R1673 B.n467 B.n466 71.676
R1674 B.n462 B.n461 71.676
R1675 B.n459 B.n458 71.676
R1676 B.n454 B.n453 71.676
R1677 B.n451 B.n450 71.676
R1678 B.n446 B.n445 71.676
R1679 B.n443 B.n442 71.676
R1680 B.n438 B.n437 71.676
R1681 B.n435 B.n434 71.676
R1682 B.n430 B.n429 71.676
R1683 B.n427 B.n426 71.676
R1684 B.n422 B.n421 71.676
R1685 B.n419 B.n418 71.676
R1686 B.n414 B.n413 71.676
R1687 B.n411 B.n410 71.676
R1688 B.n406 B.n405 71.676
R1689 B.n403 B.n402 71.676
R1690 B.n398 B.n397 71.676
R1691 B.n395 B.n394 71.676
R1692 B.n390 B.n389 71.676
R1693 B.n387 B.n386 71.676
R1694 B.n382 B.n381 71.676
R1695 B.n1241 B.n1240 71.676
R1696 B.n1241 B.n2 71.676
R1697 B.n155 B.n154 68.4611
R1698 B.n162 B.n161 68.4611
R1699 B.n356 B.n355 68.4611
R1700 B.n350 B.n349 68.4611
R1701 B.n589 B.n323 67.3651
R1702 B.n1100 B.n128 67.3651
R1703 B.n156 B.n155 59.5399
R1704 B.n984 B.n162 59.5399
R1705 B.n357 B.n356 59.5399
R1706 B.n493 B.n350 59.5399
R1707 B.n589 B.n319 39.1526
R1708 B.n595 B.n319 39.1526
R1709 B.n595 B.n315 39.1526
R1710 B.n601 B.n315 39.1526
R1711 B.n601 B.n311 39.1526
R1712 B.n607 B.n311 39.1526
R1713 B.n607 B.n307 39.1526
R1714 B.n613 B.n307 39.1526
R1715 B.n619 B.n303 39.1526
R1716 B.n619 B.n299 39.1526
R1717 B.n625 B.n299 39.1526
R1718 B.n625 B.n295 39.1526
R1719 B.n631 B.n295 39.1526
R1720 B.n631 B.n291 39.1526
R1721 B.n637 B.n291 39.1526
R1722 B.n637 B.n287 39.1526
R1723 B.n643 B.n287 39.1526
R1724 B.n643 B.n283 39.1526
R1725 B.n649 B.n283 39.1526
R1726 B.n649 B.n279 39.1526
R1727 B.n655 B.n279 39.1526
R1728 B.n661 B.n275 39.1526
R1729 B.n661 B.n271 39.1526
R1730 B.n667 B.n271 39.1526
R1731 B.n667 B.n267 39.1526
R1732 B.n673 B.n267 39.1526
R1733 B.n673 B.n263 39.1526
R1734 B.n679 B.n263 39.1526
R1735 B.n679 B.n259 39.1526
R1736 B.n685 B.n259 39.1526
R1737 B.n691 B.n255 39.1526
R1738 B.n691 B.n251 39.1526
R1739 B.n697 B.n251 39.1526
R1740 B.n697 B.n247 39.1526
R1741 B.n703 B.n247 39.1526
R1742 B.n703 B.n243 39.1526
R1743 B.n709 B.n243 39.1526
R1744 B.n709 B.n239 39.1526
R1745 B.n715 B.n239 39.1526
R1746 B.n721 B.n235 39.1526
R1747 B.n721 B.n231 39.1526
R1748 B.n727 B.n231 39.1526
R1749 B.n727 B.n227 39.1526
R1750 B.n733 B.n227 39.1526
R1751 B.n733 B.n223 39.1526
R1752 B.n739 B.n223 39.1526
R1753 B.n739 B.n218 39.1526
R1754 B.n745 B.n218 39.1526
R1755 B.n745 B.n219 39.1526
R1756 B.n751 B.n211 39.1526
R1757 B.n757 B.n211 39.1526
R1758 B.n757 B.n207 39.1526
R1759 B.n763 B.n207 39.1526
R1760 B.n763 B.n203 39.1526
R1761 B.n769 B.n203 39.1526
R1762 B.n769 B.n199 39.1526
R1763 B.n776 B.n199 39.1526
R1764 B.n776 B.n775 39.1526
R1765 B.n782 B.n192 39.1526
R1766 B.n789 B.n192 39.1526
R1767 B.n789 B.n188 39.1526
R1768 B.n795 B.n188 39.1526
R1769 B.n795 B.n4 39.1526
R1770 B.n1239 B.n4 39.1526
R1771 B.n1239 B.n1238 39.1526
R1772 B.n1238 B.n1237 39.1526
R1773 B.n1237 B.n8 39.1526
R1774 B.n12 B.n8 39.1526
R1775 B.n1230 B.n12 39.1526
R1776 B.n1230 B.n1229 39.1526
R1777 B.n1229 B.n1228 39.1526
R1778 B.n1222 B.n19 39.1526
R1779 B.n1222 B.n1221 39.1526
R1780 B.n1221 B.n1220 39.1526
R1781 B.n1220 B.n23 39.1526
R1782 B.n1214 B.n23 39.1526
R1783 B.n1214 B.n1213 39.1526
R1784 B.n1213 B.n1212 39.1526
R1785 B.n1212 B.n30 39.1526
R1786 B.n1206 B.n30 39.1526
R1787 B.n1205 B.n1204 39.1526
R1788 B.n1204 B.n37 39.1526
R1789 B.n1198 B.n37 39.1526
R1790 B.n1198 B.n1197 39.1526
R1791 B.n1197 B.n1196 39.1526
R1792 B.n1196 B.n44 39.1526
R1793 B.n1190 B.n44 39.1526
R1794 B.n1190 B.n1189 39.1526
R1795 B.n1189 B.n1188 39.1526
R1796 B.n1188 B.n51 39.1526
R1797 B.n1182 B.n1181 39.1526
R1798 B.n1181 B.n1180 39.1526
R1799 B.n1180 B.n58 39.1526
R1800 B.n1174 B.n58 39.1526
R1801 B.n1174 B.n1173 39.1526
R1802 B.n1173 B.n1172 39.1526
R1803 B.n1172 B.n65 39.1526
R1804 B.n1166 B.n65 39.1526
R1805 B.n1166 B.n1165 39.1526
R1806 B.n1164 B.n72 39.1526
R1807 B.n1158 B.n72 39.1526
R1808 B.n1158 B.n1157 39.1526
R1809 B.n1157 B.n1156 39.1526
R1810 B.n1156 B.n79 39.1526
R1811 B.n1150 B.n79 39.1526
R1812 B.n1150 B.n1149 39.1526
R1813 B.n1149 B.n1148 39.1526
R1814 B.n1148 B.n86 39.1526
R1815 B.n1142 B.n1141 39.1526
R1816 B.n1141 B.n1140 39.1526
R1817 B.n1140 B.n93 39.1526
R1818 B.n1134 B.n93 39.1526
R1819 B.n1134 B.n1133 39.1526
R1820 B.n1133 B.n1132 39.1526
R1821 B.n1132 B.n100 39.1526
R1822 B.n1126 B.n100 39.1526
R1823 B.n1126 B.n1125 39.1526
R1824 B.n1125 B.n1124 39.1526
R1825 B.n1124 B.n107 39.1526
R1826 B.n1118 B.n107 39.1526
R1827 B.n1118 B.n1117 39.1526
R1828 B.n1116 B.n114 39.1526
R1829 B.n1110 B.n114 39.1526
R1830 B.n1110 B.n1109 39.1526
R1831 B.n1109 B.n1108 39.1526
R1832 B.n1108 B.n121 39.1526
R1833 B.n1102 B.n121 39.1526
R1834 B.n1102 B.n1101 39.1526
R1835 B.n1101 B.n1100 39.1526
R1836 B.n715 B.t23 36.8495
R1837 B.n1182 B.t22 36.8495
R1838 B.t2 B.n275 32.2434
R1839 B.t6 B.n86 32.2434
R1840 B.n889 B.n888 29.1907
R1841 B.n587 B.n586 29.1907
R1842 B.n591 B.n321 29.1907
R1843 B.n1098 B.n1097 29.1907
R1844 B.n775 B.t5 27.6372
R1845 B.n19 B.t0 27.6372
R1846 B.n751 B.t1 26.4857
R1847 B.n1206 B.t3 26.4857
R1848 B.n613 B.t9 23.0311
R1849 B.t16 B.n1116 23.0311
R1850 B.n685 B.t7 21.8796
R1851 B.t4 B.n1164 21.8796
R1852 B B.n1242 18.0485
R1853 B.t7 B.n255 17.2735
R1854 B.n1165 B.t4 17.2735
R1855 B.t9 B.n303 16.1219
R1856 B.n1117 B.t16 16.1219
R1857 B.n219 B.t1 12.6673
R1858 B.t3 B.n1205 12.6673
R1859 B.n782 B.t5 11.5158
R1860 B.n1228 B.t0 11.5158
R1861 B.n587 B.n317 10.6151
R1862 B.n597 B.n317 10.6151
R1863 B.n598 B.n597 10.6151
R1864 B.n599 B.n598 10.6151
R1865 B.n599 B.n309 10.6151
R1866 B.n609 B.n309 10.6151
R1867 B.n610 B.n609 10.6151
R1868 B.n611 B.n610 10.6151
R1869 B.n611 B.n301 10.6151
R1870 B.n621 B.n301 10.6151
R1871 B.n622 B.n621 10.6151
R1872 B.n623 B.n622 10.6151
R1873 B.n623 B.n293 10.6151
R1874 B.n633 B.n293 10.6151
R1875 B.n634 B.n633 10.6151
R1876 B.n635 B.n634 10.6151
R1877 B.n635 B.n285 10.6151
R1878 B.n645 B.n285 10.6151
R1879 B.n646 B.n645 10.6151
R1880 B.n647 B.n646 10.6151
R1881 B.n647 B.n277 10.6151
R1882 B.n657 B.n277 10.6151
R1883 B.n658 B.n657 10.6151
R1884 B.n659 B.n658 10.6151
R1885 B.n659 B.n269 10.6151
R1886 B.n669 B.n269 10.6151
R1887 B.n670 B.n669 10.6151
R1888 B.n671 B.n670 10.6151
R1889 B.n671 B.n261 10.6151
R1890 B.n681 B.n261 10.6151
R1891 B.n682 B.n681 10.6151
R1892 B.n683 B.n682 10.6151
R1893 B.n683 B.n253 10.6151
R1894 B.n693 B.n253 10.6151
R1895 B.n694 B.n693 10.6151
R1896 B.n695 B.n694 10.6151
R1897 B.n695 B.n245 10.6151
R1898 B.n705 B.n245 10.6151
R1899 B.n706 B.n705 10.6151
R1900 B.n707 B.n706 10.6151
R1901 B.n707 B.n237 10.6151
R1902 B.n717 B.n237 10.6151
R1903 B.n718 B.n717 10.6151
R1904 B.n719 B.n718 10.6151
R1905 B.n719 B.n229 10.6151
R1906 B.n729 B.n229 10.6151
R1907 B.n730 B.n729 10.6151
R1908 B.n731 B.n730 10.6151
R1909 B.n731 B.n221 10.6151
R1910 B.n741 B.n221 10.6151
R1911 B.n742 B.n741 10.6151
R1912 B.n743 B.n742 10.6151
R1913 B.n743 B.n213 10.6151
R1914 B.n753 B.n213 10.6151
R1915 B.n754 B.n753 10.6151
R1916 B.n755 B.n754 10.6151
R1917 B.n755 B.n205 10.6151
R1918 B.n765 B.n205 10.6151
R1919 B.n766 B.n765 10.6151
R1920 B.n767 B.n766 10.6151
R1921 B.n767 B.n197 10.6151
R1922 B.n778 B.n197 10.6151
R1923 B.n779 B.n778 10.6151
R1924 B.n780 B.n779 10.6151
R1925 B.n780 B.n190 10.6151
R1926 B.n791 B.n190 10.6151
R1927 B.n792 B.n791 10.6151
R1928 B.n793 B.n792 10.6151
R1929 B.n793 B.n0 10.6151
R1930 B.n586 B.n585 10.6151
R1931 B.n585 B.n325 10.6151
R1932 B.n580 B.n325 10.6151
R1933 B.n580 B.n579 10.6151
R1934 B.n579 B.n327 10.6151
R1935 B.n574 B.n327 10.6151
R1936 B.n574 B.n573 10.6151
R1937 B.n573 B.n572 10.6151
R1938 B.n572 B.n329 10.6151
R1939 B.n566 B.n329 10.6151
R1940 B.n566 B.n565 10.6151
R1941 B.n565 B.n564 10.6151
R1942 B.n564 B.n331 10.6151
R1943 B.n558 B.n331 10.6151
R1944 B.n558 B.n557 10.6151
R1945 B.n557 B.n556 10.6151
R1946 B.n556 B.n333 10.6151
R1947 B.n550 B.n333 10.6151
R1948 B.n550 B.n549 10.6151
R1949 B.n549 B.n548 10.6151
R1950 B.n548 B.n335 10.6151
R1951 B.n542 B.n335 10.6151
R1952 B.n542 B.n541 10.6151
R1953 B.n541 B.n540 10.6151
R1954 B.n540 B.n337 10.6151
R1955 B.n534 B.n337 10.6151
R1956 B.n534 B.n533 10.6151
R1957 B.n533 B.n532 10.6151
R1958 B.n532 B.n339 10.6151
R1959 B.n526 B.n339 10.6151
R1960 B.n526 B.n525 10.6151
R1961 B.n525 B.n524 10.6151
R1962 B.n524 B.n341 10.6151
R1963 B.n518 B.n341 10.6151
R1964 B.n518 B.n517 10.6151
R1965 B.n517 B.n516 10.6151
R1966 B.n516 B.n343 10.6151
R1967 B.n510 B.n343 10.6151
R1968 B.n510 B.n509 10.6151
R1969 B.n509 B.n508 10.6151
R1970 B.n508 B.n345 10.6151
R1971 B.n502 B.n345 10.6151
R1972 B.n502 B.n501 10.6151
R1973 B.n501 B.n500 10.6151
R1974 B.n500 B.n347 10.6151
R1975 B.n494 B.n347 10.6151
R1976 B.n492 B.n491 10.6151
R1977 B.n491 B.n351 10.6151
R1978 B.n485 B.n351 10.6151
R1979 B.n485 B.n484 10.6151
R1980 B.n484 B.n483 10.6151
R1981 B.n483 B.n353 10.6151
R1982 B.n477 B.n353 10.6151
R1983 B.n477 B.n476 10.6151
R1984 B.n476 B.n475 10.6151
R1985 B.n471 B.n470 10.6151
R1986 B.n470 B.n359 10.6151
R1987 B.n465 B.n359 10.6151
R1988 B.n465 B.n464 10.6151
R1989 B.n464 B.n463 10.6151
R1990 B.n463 B.n361 10.6151
R1991 B.n457 B.n361 10.6151
R1992 B.n457 B.n456 10.6151
R1993 B.n456 B.n455 10.6151
R1994 B.n455 B.n363 10.6151
R1995 B.n449 B.n363 10.6151
R1996 B.n449 B.n448 10.6151
R1997 B.n448 B.n447 10.6151
R1998 B.n447 B.n365 10.6151
R1999 B.n441 B.n365 10.6151
R2000 B.n441 B.n440 10.6151
R2001 B.n440 B.n439 10.6151
R2002 B.n439 B.n367 10.6151
R2003 B.n433 B.n367 10.6151
R2004 B.n433 B.n432 10.6151
R2005 B.n432 B.n431 10.6151
R2006 B.n431 B.n369 10.6151
R2007 B.n425 B.n369 10.6151
R2008 B.n425 B.n424 10.6151
R2009 B.n424 B.n423 10.6151
R2010 B.n423 B.n371 10.6151
R2011 B.n417 B.n371 10.6151
R2012 B.n417 B.n416 10.6151
R2013 B.n416 B.n415 10.6151
R2014 B.n415 B.n373 10.6151
R2015 B.n409 B.n373 10.6151
R2016 B.n409 B.n408 10.6151
R2017 B.n408 B.n407 10.6151
R2018 B.n407 B.n375 10.6151
R2019 B.n401 B.n375 10.6151
R2020 B.n401 B.n400 10.6151
R2021 B.n400 B.n399 10.6151
R2022 B.n399 B.n377 10.6151
R2023 B.n393 B.n377 10.6151
R2024 B.n393 B.n392 10.6151
R2025 B.n392 B.n391 10.6151
R2026 B.n391 B.n379 10.6151
R2027 B.n385 B.n379 10.6151
R2028 B.n385 B.n384 10.6151
R2029 B.n384 B.n383 10.6151
R2030 B.n383 B.n321 10.6151
R2031 B.n592 B.n591 10.6151
R2032 B.n593 B.n592 10.6151
R2033 B.n593 B.n313 10.6151
R2034 B.n603 B.n313 10.6151
R2035 B.n604 B.n603 10.6151
R2036 B.n605 B.n604 10.6151
R2037 B.n605 B.n305 10.6151
R2038 B.n615 B.n305 10.6151
R2039 B.n616 B.n615 10.6151
R2040 B.n617 B.n616 10.6151
R2041 B.n617 B.n297 10.6151
R2042 B.n627 B.n297 10.6151
R2043 B.n628 B.n627 10.6151
R2044 B.n629 B.n628 10.6151
R2045 B.n629 B.n289 10.6151
R2046 B.n639 B.n289 10.6151
R2047 B.n640 B.n639 10.6151
R2048 B.n641 B.n640 10.6151
R2049 B.n641 B.n281 10.6151
R2050 B.n651 B.n281 10.6151
R2051 B.n652 B.n651 10.6151
R2052 B.n653 B.n652 10.6151
R2053 B.n653 B.n273 10.6151
R2054 B.n663 B.n273 10.6151
R2055 B.n664 B.n663 10.6151
R2056 B.n665 B.n664 10.6151
R2057 B.n665 B.n265 10.6151
R2058 B.n675 B.n265 10.6151
R2059 B.n676 B.n675 10.6151
R2060 B.n677 B.n676 10.6151
R2061 B.n677 B.n257 10.6151
R2062 B.n687 B.n257 10.6151
R2063 B.n688 B.n687 10.6151
R2064 B.n689 B.n688 10.6151
R2065 B.n689 B.n249 10.6151
R2066 B.n699 B.n249 10.6151
R2067 B.n700 B.n699 10.6151
R2068 B.n701 B.n700 10.6151
R2069 B.n701 B.n241 10.6151
R2070 B.n711 B.n241 10.6151
R2071 B.n712 B.n711 10.6151
R2072 B.n713 B.n712 10.6151
R2073 B.n713 B.n233 10.6151
R2074 B.n723 B.n233 10.6151
R2075 B.n724 B.n723 10.6151
R2076 B.n725 B.n724 10.6151
R2077 B.n725 B.n225 10.6151
R2078 B.n735 B.n225 10.6151
R2079 B.n736 B.n735 10.6151
R2080 B.n737 B.n736 10.6151
R2081 B.n737 B.n216 10.6151
R2082 B.n747 B.n216 10.6151
R2083 B.n748 B.n747 10.6151
R2084 B.n749 B.n748 10.6151
R2085 B.n749 B.n209 10.6151
R2086 B.n759 B.n209 10.6151
R2087 B.n760 B.n759 10.6151
R2088 B.n761 B.n760 10.6151
R2089 B.n761 B.n201 10.6151
R2090 B.n771 B.n201 10.6151
R2091 B.n772 B.n771 10.6151
R2092 B.n773 B.n772 10.6151
R2093 B.n773 B.n194 10.6151
R2094 B.n784 B.n194 10.6151
R2095 B.n785 B.n784 10.6151
R2096 B.n787 B.n785 10.6151
R2097 B.n787 B.n786 10.6151
R2098 B.n786 B.n186 10.6151
R2099 B.n798 B.n186 10.6151
R2100 B.n799 B.n798 10.6151
R2101 B.n800 B.n799 10.6151
R2102 B.n801 B.n800 10.6151
R2103 B.n802 B.n801 10.6151
R2104 B.n805 B.n802 10.6151
R2105 B.n806 B.n805 10.6151
R2106 B.n807 B.n806 10.6151
R2107 B.n808 B.n807 10.6151
R2108 B.n810 B.n808 10.6151
R2109 B.n811 B.n810 10.6151
R2110 B.n812 B.n811 10.6151
R2111 B.n813 B.n812 10.6151
R2112 B.n815 B.n813 10.6151
R2113 B.n816 B.n815 10.6151
R2114 B.n817 B.n816 10.6151
R2115 B.n818 B.n817 10.6151
R2116 B.n820 B.n818 10.6151
R2117 B.n821 B.n820 10.6151
R2118 B.n822 B.n821 10.6151
R2119 B.n823 B.n822 10.6151
R2120 B.n825 B.n823 10.6151
R2121 B.n826 B.n825 10.6151
R2122 B.n827 B.n826 10.6151
R2123 B.n828 B.n827 10.6151
R2124 B.n830 B.n828 10.6151
R2125 B.n831 B.n830 10.6151
R2126 B.n832 B.n831 10.6151
R2127 B.n833 B.n832 10.6151
R2128 B.n835 B.n833 10.6151
R2129 B.n836 B.n835 10.6151
R2130 B.n837 B.n836 10.6151
R2131 B.n838 B.n837 10.6151
R2132 B.n840 B.n838 10.6151
R2133 B.n841 B.n840 10.6151
R2134 B.n842 B.n841 10.6151
R2135 B.n843 B.n842 10.6151
R2136 B.n845 B.n843 10.6151
R2137 B.n846 B.n845 10.6151
R2138 B.n847 B.n846 10.6151
R2139 B.n848 B.n847 10.6151
R2140 B.n850 B.n848 10.6151
R2141 B.n851 B.n850 10.6151
R2142 B.n852 B.n851 10.6151
R2143 B.n853 B.n852 10.6151
R2144 B.n855 B.n853 10.6151
R2145 B.n856 B.n855 10.6151
R2146 B.n857 B.n856 10.6151
R2147 B.n858 B.n857 10.6151
R2148 B.n860 B.n858 10.6151
R2149 B.n861 B.n860 10.6151
R2150 B.n862 B.n861 10.6151
R2151 B.n863 B.n862 10.6151
R2152 B.n865 B.n863 10.6151
R2153 B.n866 B.n865 10.6151
R2154 B.n867 B.n866 10.6151
R2155 B.n868 B.n867 10.6151
R2156 B.n870 B.n868 10.6151
R2157 B.n871 B.n870 10.6151
R2158 B.n872 B.n871 10.6151
R2159 B.n873 B.n872 10.6151
R2160 B.n875 B.n873 10.6151
R2161 B.n876 B.n875 10.6151
R2162 B.n877 B.n876 10.6151
R2163 B.n878 B.n877 10.6151
R2164 B.n880 B.n878 10.6151
R2165 B.n881 B.n880 10.6151
R2166 B.n882 B.n881 10.6151
R2167 B.n883 B.n882 10.6151
R2168 B.n885 B.n883 10.6151
R2169 B.n886 B.n885 10.6151
R2170 B.n887 B.n886 10.6151
R2171 B.n888 B.n887 10.6151
R2172 B.n1234 B.n1 10.6151
R2173 B.n1234 B.n1233 10.6151
R2174 B.n1233 B.n1232 10.6151
R2175 B.n1232 B.n10 10.6151
R2176 B.n1226 B.n10 10.6151
R2177 B.n1226 B.n1225 10.6151
R2178 B.n1225 B.n1224 10.6151
R2179 B.n1224 B.n17 10.6151
R2180 B.n1218 B.n17 10.6151
R2181 B.n1218 B.n1217 10.6151
R2182 B.n1217 B.n1216 10.6151
R2183 B.n1216 B.n25 10.6151
R2184 B.n1210 B.n25 10.6151
R2185 B.n1210 B.n1209 10.6151
R2186 B.n1209 B.n1208 10.6151
R2187 B.n1208 B.n32 10.6151
R2188 B.n1202 B.n32 10.6151
R2189 B.n1202 B.n1201 10.6151
R2190 B.n1201 B.n1200 10.6151
R2191 B.n1200 B.n39 10.6151
R2192 B.n1194 B.n39 10.6151
R2193 B.n1194 B.n1193 10.6151
R2194 B.n1193 B.n1192 10.6151
R2195 B.n1192 B.n46 10.6151
R2196 B.n1186 B.n46 10.6151
R2197 B.n1186 B.n1185 10.6151
R2198 B.n1185 B.n1184 10.6151
R2199 B.n1184 B.n53 10.6151
R2200 B.n1178 B.n53 10.6151
R2201 B.n1178 B.n1177 10.6151
R2202 B.n1177 B.n1176 10.6151
R2203 B.n1176 B.n60 10.6151
R2204 B.n1170 B.n60 10.6151
R2205 B.n1170 B.n1169 10.6151
R2206 B.n1169 B.n1168 10.6151
R2207 B.n1168 B.n67 10.6151
R2208 B.n1162 B.n67 10.6151
R2209 B.n1162 B.n1161 10.6151
R2210 B.n1161 B.n1160 10.6151
R2211 B.n1160 B.n74 10.6151
R2212 B.n1154 B.n74 10.6151
R2213 B.n1154 B.n1153 10.6151
R2214 B.n1153 B.n1152 10.6151
R2215 B.n1152 B.n81 10.6151
R2216 B.n1146 B.n81 10.6151
R2217 B.n1146 B.n1145 10.6151
R2218 B.n1145 B.n1144 10.6151
R2219 B.n1144 B.n88 10.6151
R2220 B.n1138 B.n88 10.6151
R2221 B.n1138 B.n1137 10.6151
R2222 B.n1137 B.n1136 10.6151
R2223 B.n1136 B.n95 10.6151
R2224 B.n1130 B.n95 10.6151
R2225 B.n1130 B.n1129 10.6151
R2226 B.n1129 B.n1128 10.6151
R2227 B.n1128 B.n102 10.6151
R2228 B.n1122 B.n102 10.6151
R2229 B.n1122 B.n1121 10.6151
R2230 B.n1121 B.n1120 10.6151
R2231 B.n1120 B.n109 10.6151
R2232 B.n1114 B.n109 10.6151
R2233 B.n1114 B.n1113 10.6151
R2234 B.n1113 B.n1112 10.6151
R2235 B.n1112 B.n116 10.6151
R2236 B.n1106 B.n116 10.6151
R2237 B.n1106 B.n1105 10.6151
R2238 B.n1105 B.n1104 10.6151
R2239 B.n1104 B.n123 10.6151
R2240 B.n1098 B.n123 10.6151
R2241 B.n1097 B.n1096 10.6151
R2242 B.n1096 B.n130 10.6151
R2243 B.n1090 B.n130 10.6151
R2244 B.n1090 B.n1089 10.6151
R2245 B.n1089 B.n1088 10.6151
R2246 B.n1088 B.n132 10.6151
R2247 B.n1082 B.n132 10.6151
R2248 B.n1082 B.n1081 10.6151
R2249 B.n1081 B.n1080 10.6151
R2250 B.n1080 B.n134 10.6151
R2251 B.n1074 B.n134 10.6151
R2252 B.n1074 B.n1073 10.6151
R2253 B.n1073 B.n1072 10.6151
R2254 B.n1072 B.n136 10.6151
R2255 B.n1066 B.n136 10.6151
R2256 B.n1066 B.n1065 10.6151
R2257 B.n1065 B.n1064 10.6151
R2258 B.n1064 B.n138 10.6151
R2259 B.n1058 B.n138 10.6151
R2260 B.n1058 B.n1057 10.6151
R2261 B.n1057 B.n1056 10.6151
R2262 B.n1056 B.n140 10.6151
R2263 B.n1050 B.n140 10.6151
R2264 B.n1050 B.n1049 10.6151
R2265 B.n1049 B.n1048 10.6151
R2266 B.n1048 B.n142 10.6151
R2267 B.n1042 B.n142 10.6151
R2268 B.n1042 B.n1041 10.6151
R2269 B.n1041 B.n1040 10.6151
R2270 B.n1040 B.n144 10.6151
R2271 B.n1034 B.n144 10.6151
R2272 B.n1034 B.n1033 10.6151
R2273 B.n1033 B.n1032 10.6151
R2274 B.n1032 B.n146 10.6151
R2275 B.n1026 B.n146 10.6151
R2276 B.n1026 B.n1025 10.6151
R2277 B.n1025 B.n1024 10.6151
R2278 B.n1024 B.n148 10.6151
R2279 B.n1018 B.n148 10.6151
R2280 B.n1018 B.n1017 10.6151
R2281 B.n1017 B.n1016 10.6151
R2282 B.n1016 B.n150 10.6151
R2283 B.n1010 B.n150 10.6151
R2284 B.n1010 B.n1009 10.6151
R2285 B.n1009 B.n1008 10.6151
R2286 B.n1008 B.n152 10.6151
R2287 B.n1002 B.n1001 10.6151
R2288 B.n1001 B.n1000 10.6151
R2289 B.n1000 B.n157 10.6151
R2290 B.n994 B.n157 10.6151
R2291 B.n994 B.n993 10.6151
R2292 B.n993 B.n992 10.6151
R2293 B.n992 B.n159 10.6151
R2294 B.n986 B.n159 10.6151
R2295 B.n986 B.n985 10.6151
R2296 B.n983 B.n163 10.6151
R2297 B.n977 B.n163 10.6151
R2298 B.n977 B.n976 10.6151
R2299 B.n976 B.n975 10.6151
R2300 B.n975 B.n165 10.6151
R2301 B.n969 B.n165 10.6151
R2302 B.n969 B.n968 10.6151
R2303 B.n968 B.n967 10.6151
R2304 B.n967 B.n167 10.6151
R2305 B.n961 B.n167 10.6151
R2306 B.n961 B.n960 10.6151
R2307 B.n960 B.n959 10.6151
R2308 B.n959 B.n169 10.6151
R2309 B.n953 B.n169 10.6151
R2310 B.n953 B.n952 10.6151
R2311 B.n952 B.n951 10.6151
R2312 B.n951 B.n171 10.6151
R2313 B.n945 B.n171 10.6151
R2314 B.n945 B.n944 10.6151
R2315 B.n944 B.n943 10.6151
R2316 B.n943 B.n173 10.6151
R2317 B.n937 B.n173 10.6151
R2318 B.n937 B.n936 10.6151
R2319 B.n936 B.n935 10.6151
R2320 B.n935 B.n175 10.6151
R2321 B.n929 B.n175 10.6151
R2322 B.n929 B.n928 10.6151
R2323 B.n928 B.n927 10.6151
R2324 B.n927 B.n177 10.6151
R2325 B.n921 B.n177 10.6151
R2326 B.n921 B.n920 10.6151
R2327 B.n920 B.n919 10.6151
R2328 B.n919 B.n179 10.6151
R2329 B.n913 B.n179 10.6151
R2330 B.n913 B.n912 10.6151
R2331 B.n912 B.n911 10.6151
R2332 B.n911 B.n181 10.6151
R2333 B.n905 B.n181 10.6151
R2334 B.n905 B.n904 10.6151
R2335 B.n904 B.n903 10.6151
R2336 B.n903 B.n183 10.6151
R2337 B.n897 B.n183 10.6151
R2338 B.n897 B.n896 10.6151
R2339 B.n896 B.n895 10.6151
R2340 B.n895 B.n185 10.6151
R2341 B.n889 B.n185 10.6151
R2342 B.n494 B.n493 9.36635
R2343 B.n471 B.n357 9.36635
R2344 B.n156 B.n152 9.36635
R2345 B.n984 B.n983 9.36635
R2346 B.n1242 B.n0 8.11757
R2347 B.n1242 B.n1 8.11757
R2348 B.n655 B.t2 6.90969
R2349 B.n1142 B.t6 6.90969
R2350 B.t23 B.n235 2.30356
R2351 B.t22 B.n51 2.30356
R2352 B.n493 B.n492 1.24928
R2353 B.n475 B.n357 1.24928
R2354 B.n1002 B.n156 1.24928
R2355 B.n985 B.n984 1.24928
R2356 VP.n32 VP.n31 161.3
R2357 VP.n33 VP.n28 161.3
R2358 VP.n35 VP.n34 161.3
R2359 VP.n36 VP.n27 161.3
R2360 VP.n38 VP.n37 161.3
R2361 VP.n39 VP.n26 161.3
R2362 VP.n41 VP.n40 161.3
R2363 VP.n43 VP.n42 161.3
R2364 VP.n44 VP.n24 161.3
R2365 VP.n46 VP.n45 161.3
R2366 VP.n47 VP.n23 161.3
R2367 VP.n49 VP.n48 161.3
R2368 VP.n50 VP.n22 161.3
R2369 VP.n52 VP.n51 161.3
R2370 VP.n54 VP.n53 161.3
R2371 VP.n55 VP.n20 161.3
R2372 VP.n57 VP.n56 161.3
R2373 VP.n58 VP.n19 161.3
R2374 VP.n60 VP.n59 161.3
R2375 VP.n61 VP.n18 161.3
R2376 VP.n63 VP.n62 161.3
R2377 VP.n109 VP.n108 161.3
R2378 VP.n107 VP.n1 161.3
R2379 VP.n106 VP.n105 161.3
R2380 VP.n104 VP.n2 161.3
R2381 VP.n103 VP.n102 161.3
R2382 VP.n101 VP.n3 161.3
R2383 VP.n100 VP.n99 161.3
R2384 VP.n98 VP.n97 161.3
R2385 VP.n96 VP.n5 161.3
R2386 VP.n95 VP.n94 161.3
R2387 VP.n93 VP.n6 161.3
R2388 VP.n92 VP.n91 161.3
R2389 VP.n90 VP.n7 161.3
R2390 VP.n89 VP.n88 161.3
R2391 VP.n87 VP.n86 161.3
R2392 VP.n85 VP.n9 161.3
R2393 VP.n84 VP.n83 161.3
R2394 VP.n82 VP.n10 161.3
R2395 VP.n81 VP.n80 161.3
R2396 VP.n79 VP.n11 161.3
R2397 VP.n78 VP.n77 161.3
R2398 VP.n76 VP.n75 161.3
R2399 VP.n74 VP.n13 161.3
R2400 VP.n73 VP.n72 161.3
R2401 VP.n71 VP.n14 161.3
R2402 VP.n70 VP.n69 161.3
R2403 VP.n68 VP.n15 161.3
R2404 VP.n67 VP.n66 161.3
R2405 VP.n30 VP.t6 137.179
R2406 VP.n16 VP.t7 104.157
R2407 VP.n12 VP.t0 104.157
R2408 VP.n8 VP.t9 104.157
R2409 VP.n4 VP.t8 104.157
R2410 VP.n0 VP.t2 104.157
R2411 VP.n17 VP.t1 104.157
R2412 VP.n21 VP.t3 104.157
R2413 VP.n25 VP.t4 104.157
R2414 VP.n29 VP.t5 104.157
R2415 VP.n65 VP.n16 74.8979
R2416 VP.n110 VP.n0 74.8979
R2417 VP.n64 VP.n17 74.8979
R2418 VP.n30 VP.n29 60.5138
R2419 VP.n65 VP.n64 57.8592
R2420 VP.n69 VP.n14 44.8641
R2421 VP.n106 VP.n2 44.8641
R2422 VP.n60 VP.n19 44.8641
R2423 VP.n80 VP.n10 41.9503
R2424 VP.n95 VP.n6 41.9503
R2425 VP.n49 VP.n23 41.9503
R2426 VP.n34 VP.n27 41.9503
R2427 VP.n84 VP.n10 39.0365
R2428 VP.n91 VP.n6 39.0365
R2429 VP.n45 VP.n23 39.0365
R2430 VP.n38 VP.n27 39.0365
R2431 VP.n73 VP.n14 36.1227
R2432 VP.n102 VP.n2 36.1227
R2433 VP.n56 VP.n19 36.1227
R2434 VP.n68 VP.n67 24.4675
R2435 VP.n69 VP.n68 24.4675
R2436 VP.n74 VP.n73 24.4675
R2437 VP.n75 VP.n74 24.4675
R2438 VP.n79 VP.n78 24.4675
R2439 VP.n80 VP.n79 24.4675
R2440 VP.n85 VP.n84 24.4675
R2441 VP.n86 VP.n85 24.4675
R2442 VP.n90 VP.n89 24.4675
R2443 VP.n91 VP.n90 24.4675
R2444 VP.n96 VP.n95 24.4675
R2445 VP.n97 VP.n96 24.4675
R2446 VP.n101 VP.n100 24.4675
R2447 VP.n102 VP.n101 24.4675
R2448 VP.n107 VP.n106 24.4675
R2449 VP.n108 VP.n107 24.4675
R2450 VP.n61 VP.n60 24.4675
R2451 VP.n62 VP.n61 24.4675
R2452 VP.n50 VP.n49 24.4675
R2453 VP.n51 VP.n50 24.4675
R2454 VP.n55 VP.n54 24.4675
R2455 VP.n56 VP.n55 24.4675
R2456 VP.n39 VP.n38 24.4675
R2457 VP.n40 VP.n39 24.4675
R2458 VP.n44 VP.n43 24.4675
R2459 VP.n45 VP.n44 24.4675
R2460 VP.n33 VP.n32 24.4675
R2461 VP.n34 VP.n33 24.4675
R2462 VP.n67 VP.n16 15.17
R2463 VP.n108 VP.n0 15.17
R2464 VP.n62 VP.n17 15.17
R2465 VP.n78 VP.n12 13.702
R2466 VP.n97 VP.n4 13.702
R2467 VP.n51 VP.n21 13.702
R2468 VP.n32 VP.n29 13.702
R2469 VP.n86 VP.n8 12.234
R2470 VP.n89 VP.n8 12.234
R2471 VP.n40 VP.n25 12.234
R2472 VP.n43 VP.n25 12.234
R2473 VP.n75 VP.n12 10.766
R2474 VP.n100 VP.n4 10.766
R2475 VP.n54 VP.n21 10.766
R2476 VP.n31 VP.n30 4.13478
R2477 VP.n64 VP.n63 0.354971
R2478 VP.n66 VP.n65 0.354971
R2479 VP.n110 VP.n109 0.354971
R2480 VP VP.n110 0.26696
R2481 VP.n31 VP.n28 0.189894
R2482 VP.n35 VP.n28 0.189894
R2483 VP.n36 VP.n35 0.189894
R2484 VP.n37 VP.n36 0.189894
R2485 VP.n37 VP.n26 0.189894
R2486 VP.n41 VP.n26 0.189894
R2487 VP.n42 VP.n41 0.189894
R2488 VP.n42 VP.n24 0.189894
R2489 VP.n46 VP.n24 0.189894
R2490 VP.n47 VP.n46 0.189894
R2491 VP.n48 VP.n47 0.189894
R2492 VP.n48 VP.n22 0.189894
R2493 VP.n52 VP.n22 0.189894
R2494 VP.n53 VP.n52 0.189894
R2495 VP.n53 VP.n20 0.189894
R2496 VP.n57 VP.n20 0.189894
R2497 VP.n58 VP.n57 0.189894
R2498 VP.n59 VP.n58 0.189894
R2499 VP.n59 VP.n18 0.189894
R2500 VP.n63 VP.n18 0.189894
R2501 VP.n66 VP.n15 0.189894
R2502 VP.n70 VP.n15 0.189894
R2503 VP.n71 VP.n70 0.189894
R2504 VP.n72 VP.n71 0.189894
R2505 VP.n72 VP.n13 0.189894
R2506 VP.n76 VP.n13 0.189894
R2507 VP.n77 VP.n76 0.189894
R2508 VP.n77 VP.n11 0.189894
R2509 VP.n81 VP.n11 0.189894
R2510 VP.n82 VP.n81 0.189894
R2511 VP.n83 VP.n82 0.189894
R2512 VP.n83 VP.n9 0.189894
R2513 VP.n87 VP.n9 0.189894
R2514 VP.n88 VP.n87 0.189894
R2515 VP.n88 VP.n7 0.189894
R2516 VP.n92 VP.n7 0.189894
R2517 VP.n93 VP.n92 0.189894
R2518 VP.n94 VP.n93 0.189894
R2519 VP.n94 VP.n5 0.189894
R2520 VP.n98 VP.n5 0.189894
R2521 VP.n99 VP.n98 0.189894
R2522 VP.n99 VP.n3 0.189894
R2523 VP.n103 VP.n3 0.189894
R2524 VP.n104 VP.n103 0.189894
R2525 VP.n105 VP.n104 0.189894
R2526 VP.n105 VP.n1 0.189894
R2527 VP.n109 VP.n1 0.189894
R2528 VDD1.n1 VDD1.t3 64.2176
R2529 VDD1.n3 VDD1.t2 64.2174
R2530 VDD1.n5 VDD1.n4 61.9698
R2531 VDD1.n7 VDD1.n6 59.7429
R2532 VDD1.n1 VDD1.n0 59.7429
R2533 VDD1.n3 VDD1.n2 59.7428
R2534 VDD1.n7 VDD1.n5 52.197
R2535 VDD1 VDD1.n7 2.22464
R2536 VDD1.n6 VDD1.t6 1.43217
R2537 VDD1.n6 VDD1.t8 1.43217
R2538 VDD1.n0 VDD1.t4 1.43217
R2539 VDD1.n0 VDD1.t5 1.43217
R2540 VDD1.n4 VDD1.t1 1.43217
R2541 VDD1.n4 VDD1.t7 1.43217
R2542 VDD1.n2 VDD1.t9 1.43217
R2543 VDD1.n2 VDD1.t0 1.43217
R2544 VDD1 VDD1.n1 0.819465
R2545 VDD1.n5 VDD1.n3 0.70593
C0 VTAIL VDD2 11.4427f
C1 VDD1 VDD2 2.56308f
C2 VP VDD2 0.659926f
C3 VN VDD2 12.6946f
C4 VTAIL VDD1 11.3876f
C5 VTAIL VP 13.5241f
C6 VDD1 VP 13.196f
C7 VTAIL VN 13.5099f
C8 VDD1 VN 0.154406f
C9 VP VN 9.624259f
C10 VDD2 B 8.227177f
C11 VDD1 B 8.198031f
C12 VTAIL B 9.39802f
C13 VN B 21.15284f
C14 VP B 19.704346f
C15 VDD1.t3 B 3.10007f
C16 VDD1.t4 B 0.268565f
C17 VDD1.t5 B 0.268565f
C18 VDD1.n0 B 2.40993f
C19 VDD1.n1 B 1.01506f
C20 VDD1.t2 B 3.10005f
C21 VDD1.t9 B 0.268565f
C22 VDD1.t0 B 0.268565f
C23 VDD1.n2 B 2.40994f
C24 VDD1.n3 B 1.00689f
C25 VDD1.t1 B 0.268565f
C26 VDD1.t7 B 0.268565f
C27 VDD1.n4 B 2.43277f
C28 VDD1.n5 B 3.42024f
C29 VDD1.t6 B 0.268565f
C30 VDD1.t8 B 0.268565f
C31 VDD1.n6 B 2.40993f
C32 VDD1.n7 B 3.50563f
C33 VP.t2 B 2.25726f
C34 VP.n0 B 0.860106f
C35 VP.n1 B 0.018649f
C36 VP.n2 B 0.015568f
C37 VP.n3 B 0.018649f
C38 VP.t8 B 2.25726f
C39 VP.n4 B 0.788163f
C40 VP.n5 B 0.018649f
C41 VP.n6 B 0.015131f
C42 VP.n7 B 0.018649f
C43 VP.t9 B 2.25726f
C44 VP.n8 B 0.788163f
C45 VP.n9 B 0.018649f
C46 VP.n10 B 0.015131f
C47 VP.n11 B 0.018649f
C48 VP.t0 B 2.25726f
C49 VP.n12 B 0.788163f
C50 VP.n13 B 0.018649f
C51 VP.n14 B 0.015568f
C52 VP.n15 B 0.018649f
C53 VP.t7 B 2.25726f
C54 VP.n16 B 0.860106f
C55 VP.t1 B 2.25726f
C56 VP.n17 B 0.860106f
C57 VP.n18 B 0.018649f
C58 VP.n19 B 0.015568f
C59 VP.n20 B 0.018649f
C60 VP.t3 B 2.25726f
C61 VP.n21 B 0.788163f
C62 VP.n22 B 0.018649f
C63 VP.n23 B 0.015131f
C64 VP.n24 B 0.018649f
C65 VP.t4 B 2.25726f
C66 VP.n25 B 0.788163f
C67 VP.n26 B 0.018649f
C68 VP.n27 B 0.015131f
C69 VP.n28 B 0.018649f
C70 VP.t5 B 2.25726f
C71 VP.n29 B 0.850499f
C72 VP.t6 B 2.47861f
C73 VP.n30 B 0.813305f
C74 VP.n31 B 0.21672f
C75 VP.n32 B 0.027207f
C76 VP.n33 B 0.034758f
C77 VP.n34 B 0.03676f
C78 VP.n35 B 0.018649f
C79 VP.n36 B 0.018649f
C80 VP.n37 B 0.018649f
C81 VP.n38 B 0.037319f
C82 VP.n39 B 0.034758f
C83 VP.n40 B 0.026178f
C84 VP.n41 B 0.018649f
C85 VP.n42 B 0.018649f
C86 VP.n43 B 0.026178f
C87 VP.n44 B 0.034758f
C88 VP.n45 B 0.037319f
C89 VP.n46 B 0.018649f
C90 VP.n47 B 0.018649f
C91 VP.n48 B 0.018649f
C92 VP.n49 B 0.03676f
C93 VP.n50 B 0.034758f
C94 VP.n51 B 0.027207f
C95 VP.n52 B 0.018649f
C96 VP.n53 B 0.018649f
C97 VP.n54 B 0.025148f
C98 VP.n55 B 0.034758f
C99 VP.n56 B 0.037637f
C100 VP.n57 B 0.018649f
C101 VP.n58 B 0.018649f
C102 VP.n59 B 0.018649f
C103 VP.n60 B 0.036006f
C104 VP.n61 B 0.034758f
C105 VP.n62 B 0.028237f
C106 VP.n63 B 0.0301f
C107 VP.n64 B 1.29883f
C108 VP.n65 B 1.31042f
C109 VP.n66 B 0.0301f
C110 VP.n67 B 0.028237f
C111 VP.n68 B 0.034758f
C112 VP.n69 B 0.036006f
C113 VP.n70 B 0.018649f
C114 VP.n71 B 0.018649f
C115 VP.n72 B 0.018649f
C116 VP.n73 B 0.037637f
C117 VP.n74 B 0.034758f
C118 VP.n75 B 0.025148f
C119 VP.n76 B 0.018649f
C120 VP.n77 B 0.018649f
C121 VP.n78 B 0.027207f
C122 VP.n79 B 0.034758f
C123 VP.n80 B 0.03676f
C124 VP.n81 B 0.018649f
C125 VP.n82 B 0.018649f
C126 VP.n83 B 0.018649f
C127 VP.n84 B 0.037319f
C128 VP.n85 B 0.034758f
C129 VP.n86 B 0.026178f
C130 VP.n87 B 0.018649f
C131 VP.n88 B 0.018649f
C132 VP.n89 B 0.026178f
C133 VP.n90 B 0.034758f
C134 VP.n91 B 0.037319f
C135 VP.n92 B 0.018649f
C136 VP.n93 B 0.018649f
C137 VP.n94 B 0.018649f
C138 VP.n95 B 0.03676f
C139 VP.n96 B 0.034758f
C140 VP.n97 B 0.027207f
C141 VP.n98 B 0.018649f
C142 VP.n99 B 0.018649f
C143 VP.n100 B 0.025148f
C144 VP.n101 B 0.034758f
C145 VP.n102 B 0.037637f
C146 VP.n103 B 0.018649f
C147 VP.n104 B 0.018649f
C148 VP.n105 B 0.018649f
C149 VP.n106 B 0.036006f
C150 VP.n107 B 0.034758f
C151 VP.n108 B 0.028237f
C152 VP.n109 B 0.0301f
C153 VP.n110 B 0.044004f
C154 VDD2.t9 B 3.05326f
C155 VDD2.t5 B 0.264511f
C156 VDD2.t1 B 0.264511f
C157 VDD2.n0 B 2.37356f
C158 VDD2.n1 B 0.991687f
C159 VDD2.t6 B 0.264511f
C160 VDD2.t0 B 0.264511f
C161 VDD2.n2 B 2.39605f
C162 VDD2.n3 B 3.23042f
C163 VDD2.t8 B 3.02871f
C164 VDD2.n4 B 3.39429f
C165 VDD2.t7 B 0.264511f
C166 VDD2.t2 B 0.264511f
C167 VDD2.n5 B 2.37355f
C168 VDD2.n6 B 0.506087f
C169 VDD2.t4 B 0.264511f
C170 VDD2.t3 B 0.264511f
C171 VDD2.n7 B 2.396f
C172 VTAIL.t11 B 0.271372f
C173 VTAIL.t13 B 0.271372f
C174 VTAIL.n0 B 2.35554f
C175 VTAIL.n1 B 0.602638f
C176 VTAIL.t5 B 3.00475f
C177 VTAIL.n2 B 0.74974f
C178 VTAIL.t19 B 0.271372f
C179 VTAIL.t1 B 0.271372f
C180 VTAIL.n3 B 2.35554f
C181 VTAIL.n4 B 0.743f
C182 VTAIL.t2 B 0.271372f
C183 VTAIL.t7 B 0.271372f
C184 VTAIL.n5 B 2.35554f
C185 VTAIL.n6 B 2.27769f
C186 VTAIL.t12 B 0.271372f
C187 VTAIL.t16 B 0.271372f
C188 VTAIL.n7 B 2.35553f
C189 VTAIL.n8 B 2.27769f
C190 VTAIL.t10 B 0.271372f
C191 VTAIL.t9 B 0.271372f
C192 VTAIL.n9 B 2.35553f
C193 VTAIL.n10 B 0.743002f
C194 VTAIL.t14 B 3.00477f
C195 VTAIL.n11 B 0.749721f
C196 VTAIL.t0 B 0.271372f
C197 VTAIL.t3 B 0.271372f
C198 VTAIL.n12 B 2.35553f
C199 VTAIL.n13 B 0.658853f
C200 VTAIL.t18 B 0.271372f
C201 VTAIL.t4 B 0.271372f
C202 VTAIL.n14 B 2.35553f
C203 VTAIL.n15 B 0.743002f
C204 VTAIL.t6 B 3.00477f
C205 VTAIL.n16 B 2.12508f
C206 VTAIL.t15 B 3.00475f
C207 VTAIL.n17 B 2.1251f
C208 VTAIL.t17 B 0.271372f
C209 VTAIL.t8 B 0.271372f
C210 VTAIL.n18 B 2.35554f
C211 VTAIL.n19 B 0.555735f
C212 VN.t9 B 2.22456f
C213 VN.n0 B 0.847647f
C214 VN.n1 B 0.018379f
C215 VN.n2 B 0.015342f
C216 VN.n3 B 0.018379f
C217 VN.t3 B 2.22456f
C218 VN.n4 B 0.776745f
C219 VN.n5 B 0.018379f
C220 VN.n6 B 0.014912f
C221 VN.n7 B 0.018379f
C222 VN.t8 B 2.22456f
C223 VN.n8 B 0.776745f
C224 VN.n9 B 0.018379f
C225 VN.n10 B 0.014912f
C226 VN.n11 B 0.018379f
C227 VN.t4 B 2.22456f
C228 VN.n12 B 0.838179f
C229 VN.t0 B 2.44271f
C230 VN.n13 B 0.801523f
C231 VN.n14 B 0.21358f
C232 VN.n15 B 0.026813f
C233 VN.n16 B 0.034254f
C234 VN.n17 B 0.036228f
C235 VN.n18 B 0.018379f
C236 VN.n19 B 0.018379f
C237 VN.n20 B 0.018379f
C238 VN.n21 B 0.036779f
C239 VN.n22 B 0.034254f
C240 VN.n23 B 0.025798f
C241 VN.n24 B 0.018379f
C242 VN.n25 B 0.018379f
C243 VN.n26 B 0.025798f
C244 VN.n27 B 0.034254f
C245 VN.n28 B 0.036779f
C246 VN.n29 B 0.018379f
C247 VN.n30 B 0.018379f
C248 VN.n31 B 0.018379f
C249 VN.n32 B 0.036228f
C250 VN.n33 B 0.034254f
C251 VN.n34 B 0.026813f
C252 VN.n35 B 0.018379f
C253 VN.n36 B 0.018379f
C254 VN.n37 B 0.024784f
C255 VN.n38 B 0.034254f
C256 VN.n39 B 0.037092f
C257 VN.n40 B 0.018379f
C258 VN.n41 B 0.018379f
C259 VN.n42 B 0.018379f
C260 VN.n43 B 0.035484f
C261 VN.n44 B 0.034254f
C262 VN.n45 B 0.027828f
C263 VN.n46 B 0.029664f
C264 VN.n47 B 0.043366f
C265 VN.t1 B 2.22456f
C266 VN.n48 B 0.847647f
C267 VN.n49 B 0.018379f
C268 VN.n50 B 0.015342f
C269 VN.n51 B 0.018379f
C270 VN.t2 B 2.22456f
C271 VN.n52 B 0.776745f
C272 VN.n53 B 0.018379f
C273 VN.n54 B 0.014912f
C274 VN.n55 B 0.018379f
C275 VN.t7 B 2.22456f
C276 VN.n56 B 0.776745f
C277 VN.n57 B 0.018379f
C278 VN.n58 B 0.014912f
C279 VN.n59 B 0.018379f
C280 VN.t5 B 2.22456f
C281 VN.n60 B 0.838179f
C282 VN.t6 B 2.44271f
C283 VN.n61 B 0.801523f
C284 VN.n62 B 0.21358f
C285 VN.n63 B 0.026813f
C286 VN.n64 B 0.034254f
C287 VN.n65 B 0.036228f
C288 VN.n66 B 0.018379f
C289 VN.n67 B 0.018379f
C290 VN.n68 B 0.018379f
C291 VN.n69 B 0.036779f
C292 VN.n70 B 0.034254f
C293 VN.n71 B 0.025798f
C294 VN.n72 B 0.018379f
C295 VN.n73 B 0.018379f
C296 VN.n74 B 0.025798f
C297 VN.n75 B 0.034254f
C298 VN.n76 B 0.036779f
C299 VN.n77 B 0.018379f
C300 VN.n78 B 0.018379f
C301 VN.n79 B 0.018379f
C302 VN.n80 B 0.036228f
C303 VN.n81 B 0.034254f
C304 VN.n82 B 0.026813f
C305 VN.n83 B 0.018379f
C306 VN.n84 B 0.018379f
C307 VN.n85 B 0.024784f
C308 VN.n86 B 0.034254f
C309 VN.n87 B 0.037092f
C310 VN.n88 B 0.018379f
C311 VN.n89 B 0.018379f
C312 VN.n90 B 0.018379f
C313 VN.n91 B 0.035484f
C314 VN.n92 B 0.034254f
C315 VN.n93 B 0.027828f
C316 VN.n94 B 0.029664f
C317 VN.n95 B 1.28719f
.ends

