* NGSPICE file created from diff_pair_sample_1210.ext - technology: sky130A

.subckt diff_pair_sample_1210 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=2.42
X1 VDD1.t4 VP.t1 VTAIL.t5 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=2.42
X2 B.t11 B.t9 B.t10 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=2.42
X3 VTAIL.t9 VP.t2 VDD1.t3 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=1.83975 ps=11.48 w=11.15 l=2.42
X4 VDD2.t5 VN.t0 VTAIL.t0 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=2.42
X5 VDD2.t4 VN.t1 VTAIL.t4 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=2.42
X6 VDD2.t3 VN.t2 VTAIL.t3 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=2.42
X7 B.t8 B.t6 B.t7 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=2.42
X8 VDD2.t2 VN.t3 VTAIL.t11 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=2.42
X9 B.t5 B.t3 B.t4 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=2.42
X10 VTAIL.t10 VP.t3 VDD1.t2 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=1.83975 ps=11.48 w=11.15 l=2.42
X11 VTAIL.t1 VN.t4 VDD2.t1 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=1.83975 ps=11.48 w=11.15 l=2.42
X12 VTAIL.t2 VN.t5 VDD2.t0 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=1.83975 ps=11.48 w=11.15 l=2.42
X13 VDD1.t1 VP.t4 VTAIL.t6 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=1.83975 pd=11.48 as=4.3485 ps=23.08 w=11.15 l=2.42
X14 VDD1.t0 VP.t5 VTAIL.t7 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=1.83975 ps=11.48 w=11.15 l=2.42
X15 B.t2 B.t0 B.t1 w_n3170_n3198# sky130_fd_pr__pfet_01v8 ad=4.3485 pd=23.08 as=0 ps=0 w=11.15 l=2.42
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n37 VP.n0 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n34 VP.n1 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n31 VP.n2 161.3
R10 VP.n30 VP.n29 161.3
R11 VP.n28 VP.n3 161.3
R12 VP.n27 VP.n26 161.3
R13 VP.n25 VP.n4 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n5 161.3
R16 VP.n9 VP.t0 145.423
R17 VP.n30 VP.t3 111.04
R18 VP.n20 VP.t5 111.04
R19 VP.n38 VP.t1 111.04
R20 VP.n10 VP.t2 111.04
R21 VP.n18 VP.t4 111.04
R22 VP.n21 VP.n20 98.5229
R23 VP.n39 VP.n38 98.5229
R24 VP.n19 VP.n18 98.5229
R25 VP.n26 VP.n25 52.6342
R26 VP.n32 VP.n1 52.6342
R27 VP.n12 VP.n7 52.6342
R28 VP.n10 VP.n9 48.0049
R29 VP.n21 VP.n19 47.3367
R30 VP.n25 VP.n24 28.3526
R31 VP.n36 VP.n1 28.3526
R32 VP.n16 VP.n7 28.3526
R33 VP.n24 VP.n5 24.4675
R34 VP.n26 VP.n3 24.4675
R35 VP.n30 VP.n3 24.4675
R36 VP.n31 VP.n30 24.4675
R37 VP.n32 VP.n31 24.4675
R38 VP.n37 VP.n36 24.4675
R39 VP.n17 VP.n16 24.4675
R40 VP.n11 VP.n10 24.4675
R41 VP.n12 VP.n11 24.4675
R42 VP.n20 VP.n5 12.234
R43 VP.n38 VP.n37 12.234
R44 VP.n18 VP.n17 12.234
R45 VP.n9 VP.n8 6.69041
R46 VP.n19 VP.n6 0.278367
R47 VP.n22 VP.n21 0.278367
R48 VP.n39 VP.n0 0.278367
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153454
R64 VTAIL.n7 VTAIL.t11 63.6748
R65 VTAIL.n11 VTAIL.t4 63.6747
R66 VTAIL.n2 VTAIL.t5 63.6747
R67 VTAIL.n10 VTAIL.t6 63.6747
R68 VTAIL.n9 VTAIL.n8 60.7596
R69 VTAIL.n6 VTAIL.n5 60.7596
R70 VTAIL.n1 VTAIL.n0 60.7593
R71 VTAIL.n4 VTAIL.n3 60.7593
R72 VTAIL.n6 VTAIL.n4 26.7203
R73 VTAIL.n11 VTAIL.n10 24.3496
R74 VTAIL.n0 VTAIL.t3 2.91575
R75 VTAIL.n0 VTAIL.t1 2.91575
R76 VTAIL.n3 VTAIL.t7 2.91575
R77 VTAIL.n3 VTAIL.t10 2.91575
R78 VTAIL.n8 VTAIL.t8 2.91575
R79 VTAIL.n8 VTAIL.t9 2.91575
R80 VTAIL.n5 VTAIL.t0 2.91575
R81 VTAIL.n5 VTAIL.t2 2.91575
R82 VTAIL.n7 VTAIL.n6 2.37119
R83 VTAIL.n10 VTAIL.n9 2.37119
R84 VTAIL.n4 VTAIL.n2 2.37119
R85 VTAIL VTAIL.n11 1.72033
R86 VTAIL.n9 VTAIL.n7 1.65567
R87 VTAIL.n2 VTAIL.n1 1.65567
R88 VTAIL VTAIL.n1 0.651362
R89 VDD1 VDD1.t5 82.1898
R90 VDD1.n1 VDD1.t0 82.0761
R91 VDD1.n1 VDD1.n0 77.9755
R92 VDD1.n3 VDD1.n2 77.4382
R93 VDD1.n3 VDD1.n1 42.8005
R94 VDD1.n2 VDD1.t3 2.91575
R95 VDD1.n2 VDD1.t1 2.91575
R96 VDD1.n0 VDD1.t2 2.91575
R97 VDD1.n0 VDD1.t4 2.91575
R98 VDD1 VDD1.n3 0.534983
R99 B.n371 B.n112 585
R100 B.n370 B.n369 585
R101 B.n368 B.n113 585
R102 B.n367 B.n366 585
R103 B.n365 B.n114 585
R104 B.n364 B.n363 585
R105 B.n362 B.n115 585
R106 B.n361 B.n360 585
R107 B.n359 B.n116 585
R108 B.n358 B.n357 585
R109 B.n356 B.n117 585
R110 B.n355 B.n354 585
R111 B.n353 B.n118 585
R112 B.n352 B.n351 585
R113 B.n350 B.n119 585
R114 B.n349 B.n348 585
R115 B.n347 B.n120 585
R116 B.n346 B.n345 585
R117 B.n344 B.n121 585
R118 B.n343 B.n342 585
R119 B.n341 B.n122 585
R120 B.n340 B.n339 585
R121 B.n338 B.n123 585
R122 B.n337 B.n336 585
R123 B.n335 B.n124 585
R124 B.n334 B.n333 585
R125 B.n332 B.n125 585
R126 B.n331 B.n330 585
R127 B.n329 B.n126 585
R128 B.n328 B.n327 585
R129 B.n326 B.n127 585
R130 B.n325 B.n324 585
R131 B.n323 B.n128 585
R132 B.n322 B.n321 585
R133 B.n320 B.n129 585
R134 B.n319 B.n318 585
R135 B.n317 B.n130 585
R136 B.n316 B.n315 585
R137 B.n314 B.n131 585
R138 B.n313 B.n312 585
R139 B.n308 B.n132 585
R140 B.n307 B.n306 585
R141 B.n305 B.n133 585
R142 B.n304 B.n303 585
R143 B.n302 B.n134 585
R144 B.n301 B.n300 585
R145 B.n299 B.n135 585
R146 B.n298 B.n297 585
R147 B.n296 B.n136 585
R148 B.n294 B.n293 585
R149 B.n292 B.n139 585
R150 B.n291 B.n290 585
R151 B.n289 B.n140 585
R152 B.n288 B.n287 585
R153 B.n286 B.n141 585
R154 B.n285 B.n284 585
R155 B.n283 B.n142 585
R156 B.n282 B.n281 585
R157 B.n280 B.n143 585
R158 B.n279 B.n278 585
R159 B.n277 B.n144 585
R160 B.n276 B.n275 585
R161 B.n274 B.n145 585
R162 B.n273 B.n272 585
R163 B.n271 B.n146 585
R164 B.n270 B.n269 585
R165 B.n268 B.n147 585
R166 B.n267 B.n266 585
R167 B.n265 B.n148 585
R168 B.n264 B.n263 585
R169 B.n262 B.n149 585
R170 B.n261 B.n260 585
R171 B.n259 B.n150 585
R172 B.n258 B.n257 585
R173 B.n256 B.n151 585
R174 B.n255 B.n254 585
R175 B.n253 B.n152 585
R176 B.n252 B.n251 585
R177 B.n250 B.n153 585
R178 B.n249 B.n248 585
R179 B.n247 B.n154 585
R180 B.n246 B.n245 585
R181 B.n244 B.n155 585
R182 B.n243 B.n242 585
R183 B.n241 B.n156 585
R184 B.n240 B.n239 585
R185 B.n238 B.n157 585
R186 B.n237 B.n236 585
R187 B.n373 B.n372 585
R188 B.n374 B.n111 585
R189 B.n376 B.n375 585
R190 B.n377 B.n110 585
R191 B.n379 B.n378 585
R192 B.n380 B.n109 585
R193 B.n382 B.n381 585
R194 B.n383 B.n108 585
R195 B.n385 B.n384 585
R196 B.n386 B.n107 585
R197 B.n388 B.n387 585
R198 B.n389 B.n106 585
R199 B.n391 B.n390 585
R200 B.n392 B.n105 585
R201 B.n394 B.n393 585
R202 B.n395 B.n104 585
R203 B.n397 B.n396 585
R204 B.n398 B.n103 585
R205 B.n400 B.n399 585
R206 B.n401 B.n102 585
R207 B.n403 B.n402 585
R208 B.n404 B.n101 585
R209 B.n406 B.n405 585
R210 B.n407 B.n100 585
R211 B.n409 B.n408 585
R212 B.n410 B.n99 585
R213 B.n412 B.n411 585
R214 B.n413 B.n98 585
R215 B.n415 B.n414 585
R216 B.n416 B.n97 585
R217 B.n418 B.n417 585
R218 B.n419 B.n96 585
R219 B.n421 B.n420 585
R220 B.n422 B.n95 585
R221 B.n424 B.n423 585
R222 B.n425 B.n94 585
R223 B.n427 B.n426 585
R224 B.n428 B.n93 585
R225 B.n430 B.n429 585
R226 B.n431 B.n92 585
R227 B.n433 B.n432 585
R228 B.n434 B.n91 585
R229 B.n436 B.n435 585
R230 B.n437 B.n90 585
R231 B.n439 B.n438 585
R232 B.n440 B.n89 585
R233 B.n442 B.n441 585
R234 B.n443 B.n88 585
R235 B.n445 B.n444 585
R236 B.n446 B.n87 585
R237 B.n448 B.n447 585
R238 B.n449 B.n86 585
R239 B.n451 B.n450 585
R240 B.n452 B.n85 585
R241 B.n454 B.n453 585
R242 B.n455 B.n84 585
R243 B.n457 B.n456 585
R244 B.n458 B.n83 585
R245 B.n460 B.n459 585
R246 B.n461 B.n82 585
R247 B.n463 B.n462 585
R248 B.n464 B.n81 585
R249 B.n466 B.n465 585
R250 B.n467 B.n80 585
R251 B.n469 B.n468 585
R252 B.n470 B.n79 585
R253 B.n472 B.n471 585
R254 B.n473 B.n78 585
R255 B.n475 B.n474 585
R256 B.n476 B.n77 585
R257 B.n478 B.n477 585
R258 B.n479 B.n76 585
R259 B.n481 B.n480 585
R260 B.n482 B.n75 585
R261 B.n484 B.n483 585
R262 B.n485 B.n74 585
R263 B.n487 B.n486 585
R264 B.n488 B.n73 585
R265 B.n490 B.n489 585
R266 B.n491 B.n72 585
R267 B.n493 B.n492 585
R268 B.n494 B.n71 585
R269 B.n627 B.n22 585
R270 B.n626 B.n625 585
R271 B.n624 B.n23 585
R272 B.n623 B.n622 585
R273 B.n621 B.n24 585
R274 B.n620 B.n619 585
R275 B.n618 B.n25 585
R276 B.n617 B.n616 585
R277 B.n615 B.n26 585
R278 B.n614 B.n613 585
R279 B.n612 B.n27 585
R280 B.n611 B.n610 585
R281 B.n609 B.n28 585
R282 B.n608 B.n607 585
R283 B.n606 B.n29 585
R284 B.n605 B.n604 585
R285 B.n603 B.n30 585
R286 B.n602 B.n601 585
R287 B.n600 B.n31 585
R288 B.n599 B.n598 585
R289 B.n597 B.n32 585
R290 B.n596 B.n595 585
R291 B.n594 B.n33 585
R292 B.n593 B.n592 585
R293 B.n591 B.n34 585
R294 B.n590 B.n589 585
R295 B.n588 B.n35 585
R296 B.n587 B.n586 585
R297 B.n585 B.n36 585
R298 B.n584 B.n583 585
R299 B.n582 B.n37 585
R300 B.n581 B.n580 585
R301 B.n579 B.n38 585
R302 B.n578 B.n577 585
R303 B.n576 B.n39 585
R304 B.n575 B.n574 585
R305 B.n573 B.n40 585
R306 B.n572 B.n571 585
R307 B.n570 B.n41 585
R308 B.n568 B.n567 585
R309 B.n566 B.n44 585
R310 B.n565 B.n564 585
R311 B.n563 B.n45 585
R312 B.n562 B.n561 585
R313 B.n560 B.n46 585
R314 B.n559 B.n558 585
R315 B.n557 B.n47 585
R316 B.n556 B.n555 585
R317 B.n554 B.n48 585
R318 B.n553 B.n552 585
R319 B.n551 B.n49 585
R320 B.n550 B.n549 585
R321 B.n548 B.n53 585
R322 B.n547 B.n546 585
R323 B.n545 B.n54 585
R324 B.n544 B.n543 585
R325 B.n542 B.n55 585
R326 B.n541 B.n540 585
R327 B.n539 B.n56 585
R328 B.n538 B.n537 585
R329 B.n536 B.n57 585
R330 B.n535 B.n534 585
R331 B.n533 B.n58 585
R332 B.n532 B.n531 585
R333 B.n530 B.n59 585
R334 B.n529 B.n528 585
R335 B.n527 B.n60 585
R336 B.n526 B.n525 585
R337 B.n524 B.n61 585
R338 B.n523 B.n522 585
R339 B.n521 B.n62 585
R340 B.n520 B.n519 585
R341 B.n518 B.n63 585
R342 B.n517 B.n516 585
R343 B.n515 B.n64 585
R344 B.n514 B.n513 585
R345 B.n512 B.n65 585
R346 B.n511 B.n510 585
R347 B.n509 B.n66 585
R348 B.n508 B.n507 585
R349 B.n506 B.n67 585
R350 B.n505 B.n504 585
R351 B.n503 B.n68 585
R352 B.n502 B.n501 585
R353 B.n500 B.n69 585
R354 B.n499 B.n498 585
R355 B.n497 B.n70 585
R356 B.n496 B.n495 585
R357 B.n629 B.n628 585
R358 B.n630 B.n21 585
R359 B.n632 B.n631 585
R360 B.n633 B.n20 585
R361 B.n635 B.n634 585
R362 B.n636 B.n19 585
R363 B.n638 B.n637 585
R364 B.n639 B.n18 585
R365 B.n641 B.n640 585
R366 B.n642 B.n17 585
R367 B.n644 B.n643 585
R368 B.n645 B.n16 585
R369 B.n647 B.n646 585
R370 B.n648 B.n15 585
R371 B.n650 B.n649 585
R372 B.n651 B.n14 585
R373 B.n653 B.n652 585
R374 B.n654 B.n13 585
R375 B.n656 B.n655 585
R376 B.n657 B.n12 585
R377 B.n659 B.n658 585
R378 B.n660 B.n11 585
R379 B.n662 B.n661 585
R380 B.n663 B.n10 585
R381 B.n665 B.n664 585
R382 B.n666 B.n9 585
R383 B.n668 B.n667 585
R384 B.n669 B.n8 585
R385 B.n671 B.n670 585
R386 B.n672 B.n7 585
R387 B.n674 B.n673 585
R388 B.n675 B.n6 585
R389 B.n677 B.n676 585
R390 B.n678 B.n5 585
R391 B.n680 B.n679 585
R392 B.n681 B.n4 585
R393 B.n683 B.n682 585
R394 B.n684 B.n3 585
R395 B.n686 B.n685 585
R396 B.n687 B.n0 585
R397 B.n2 B.n1 585
R398 B.n178 B.n177 585
R399 B.n180 B.n179 585
R400 B.n181 B.n176 585
R401 B.n183 B.n182 585
R402 B.n184 B.n175 585
R403 B.n186 B.n185 585
R404 B.n187 B.n174 585
R405 B.n189 B.n188 585
R406 B.n190 B.n173 585
R407 B.n192 B.n191 585
R408 B.n193 B.n172 585
R409 B.n195 B.n194 585
R410 B.n196 B.n171 585
R411 B.n198 B.n197 585
R412 B.n199 B.n170 585
R413 B.n201 B.n200 585
R414 B.n202 B.n169 585
R415 B.n204 B.n203 585
R416 B.n205 B.n168 585
R417 B.n207 B.n206 585
R418 B.n208 B.n167 585
R419 B.n210 B.n209 585
R420 B.n211 B.n166 585
R421 B.n213 B.n212 585
R422 B.n214 B.n165 585
R423 B.n216 B.n215 585
R424 B.n217 B.n164 585
R425 B.n219 B.n218 585
R426 B.n220 B.n163 585
R427 B.n222 B.n221 585
R428 B.n223 B.n162 585
R429 B.n225 B.n224 585
R430 B.n226 B.n161 585
R431 B.n228 B.n227 585
R432 B.n229 B.n160 585
R433 B.n231 B.n230 585
R434 B.n232 B.n159 585
R435 B.n234 B.n233 585
R436 B.n235 B.n158 585
R437 B.n237 B.n158 478.086
R438 B.n373 B.n112 478.086
R439 B.n495 B.n494 478.086
R440 B.n628 B.n627 478.086
R441 B.n137 B.t9 318.798
R442 B.n309 B.t6 318.798
R443 B.n50 B.t3 318.798
R444 B.n42 B.t0 318.798
R445 B.n689 B.n688 256.663
R446 B.n688 B.n687 235.042
R447 B.n688 B.n2 235.042
R448 B.n309 B.t7 165.889
R449 B.n50 B.t5 165.889
R450 B.n137 B.t10 165.875
R451 B.n42 B.t2 165.875
R452 B.n238 B.n237 163.367
R453 B.n239 B.n238 163.367
R454 B.n239 B.n156 163.367
R455 B.n243 B.n156 163.367
R456 B.n244 B.n243 163.367
R457 B.n245 B.n244 163.367
R458 B.n245 B.n154 163.367
R459 B.n249 B.n154 163.367
R460 B.n250 B.n249 163.367
R461 B.n251 B.n250 163.367
R462 B.n251 B.n152 163.367
R463 B.n255 B.n152 163.367
R464 B.n256 B.n255 163.367
R465 B.n257 B.n256 163.367
R466 B.n257 B.n150 163.367
R467 B.n261 B.n150 163.367
R468 B.n262 B.n261 163.367
R469 B.n263 B.n262 163.367
R470 B.n263 B.n148 163.367
R471 B.n267 B.n148 163.367
R472 B.n268 B.n267 163.367
R473 B.n269 B.n268 163.367
R474 B.n269 B.n146 163.367
R475 B.n273 B.n146 163.367
R476 B.n274 B.n273 163.367
R477 B.n275 B.n274 163.367
R478 B.n275 B.n144 163.367
R479 B.n279 B.n144 163.367
R480 B.n280 B.n279 163.367
R481 B.n281 B.n280 163.367
R482 B.n281 B.n142 163.367
R483 B.n285 B.n142 163.367
R484 B.n286 B.n285 163.367
R485 B.n287 B.n286 163.367
R486 B.n287 B.n140 163.367
R487 B.n291 B.n140 163.367
R488 B.n292 B.n291 163.367
R489 B.n293 B.n292 163.367
R490 B.n293 B.n136 163.367
R491 B.n298 B.n136 163.367
R492 B.n299 B.n298 163.367
R493 B.n300 B.n299 163.367
R494 B.n300 B.n134 163.367
R495 B.n304 B.n134 163.367
R496 B.n305 B.n304 163.367
R497 B.n306 B.n305 163.367
R498 B.n306 B.n132 163.367
R499 B.n313 B.n132 163.367
R500 B.n314 B.n313 163.367
R501 B.n315 B.n314 163.367
R502 B.n315 B.n130 163.367
R503 B.n319 B.n130 163.367
R504 B.n320 B.n319 163.367
R505 B.n321 B.n320 163.367
R506 B.n321 B.n128 163.367
R507 B.n325 B.n128 163.367
R508 B.n326 B.n325 163.367
R509 B.n327 B.n326 163.367
R510 B.n327 B.n126 163.367
R511 B.n331 B.n126 163.367
R512 B.n332 B.n331 163.367
R513 B.n333 B.n332 163.367
R514 B.n333 B.n124 163.367
R515 B.n337 B.n124 163.367
R516 B.n338 B.n337 163.367
R517 B.n339 B.n338 163.367
R518 B.n339 B.n122 163.367
R519 B.n343 B.n122 163.367
R520 B.n344 B.n343 163.367
R521 B.n345 B.n344 163.367
R522 B.n345 B.n120 163.367
R523 B.n349 B.n120 163.367
R524 B.n350 B.n349 163.367
R525 B.n351 B.n350 163.367
R526 B.n351 B.n118 163.367
R527 B.n355 B.n118 163.367
R528 B.n356 B.n355 163.367
R529 B.n357 B.n356 163.367
R530 B.n357 B.n116 163.367
R531 B.n361 B.n116 163.367
R532 B.n362 B.n361 163.367
R533 B.n363 B.n362 163.367
R534 B.n363 B.n114 163.367
R535 B.n367 B.n114 163.367
R536 B.n368 B.n367 163.367
R537 B.n369 B.n368 163.367
R538 B.n369 B.n112 163.367
R539 B.n494 B.n493 163.367
R540 B.n493 B.n72 163.367
R541 B.n489 B.n72 163.367
R542 B.n489 B.n488 163.367
R543 B.n488 B.n487 163.367
R544 B.n487 B.n74 163.367
R545 B.n483 B.n74 163.367
R546 B.n483 B.n482 163.367
R547 B.n482 B.n481 163.367
R548 B.n481 B.n76 163.367
R549 B.n477 B.n76 163.367
R550 B.n477 B.n476 163.367
R551 B.n476 B.n475 163.367
R552 B.n475 B.n78 163.367
R553 B.n471 B.n78 163.367
R554 B.n471 B.n470 163.367
R555 B.n470 B.n469 163.367
R556 B.n469 B.n80 163.367
R557 B.n465 B.n80 163.367
R558 B.n465 B.n464 163.367
R559 B.n464 B.n463 163.367
R560 B.n463 B.n82 163.367
R561 B.n459 B.n82 163.367
R562 B.n459 B.n458 163.367
R563 B.n458 B.n457 163.367
R564 B.n457 B.n84 163.367
R565 B.n453 B.n84 163.367
R566 B.n453 B.n452 163.367
R567 B.n452 B.n451 163.367
R568 B.n451 B.n86 163.367
R569 B.n447 B.n86 163.367
R570 B.n447 B.n446 163.367
R571 B.n446 B.n445 163.367
R572 B.n445 B.n88 163.367
R573 B.n441 B.n88 163.367
R574 B.n441 B.n440 163.367
R575 B.n440 B.n439 163.367
R576 B.n439 B.n90 163.367
R577 B.n435 B.n90 163.367
R578 B.n435 B.n434 163.367
R579 B.n434 B.n433 163.367
R580 B.n433 B.n92 163.367
R581 B.n429 B.n92 163.367
R582 B.n429 B.n428 163.367
R583 B.n428 B.n427 163.367
R584 B.n427 B.n94 163.367
R585 B.n423 B.n94 163.367
R586 B.n423 B.n422 163.367
R587 B.n422 B.n421 163.367
R588 B.n421 B.n96 163.367
R589 B.n417 B.n96 163.367
R590 B.n417 B.n416 163.367
R591 B.n416 B.n415 163.367
R592 B.n415 B.n98 163.367
R593 B.n411 B.n98 163.367
R594 B.n411 B.n410 163.367
R595 B.n410 B.n409 163.367
R596 B.n409 B.n100 163.367
R597 B.n405 B.n100 163.367
R598 B.n405 B.n404 163.367
R599 B.n404 B.n403 163.367
R600 B.n403 B.n102 163.367
R601 B.n399 B.n102 163.367
R602 B.n399 B.n398 163.367
R603 B.n398 B.n397 163.367
R604 B.n397 B.n104 163.367
R605 B.n393 B.n104 163.367
R606 B.n393 B.n392 163.367
R607 B.n392 B.n391 163.367
R608 B.n391 B.n106 163.367
R609 B.n387 B.n106 163.367
R610 B.n387 B.n386 163.367
R611 B.n386 B.n385 163.367
R612 B.n385 B.n108 163.367
R613 B.n381 B.n108 163.367
R614 B.n381 B.n380 163.367
R615 B.n380 B.n379 163.367
R616 B.n379 B.n110 163.367
R617 B.n375 B.n110 163.367
R618 B.n375 B.n374 163.367
R619 B.n374 B.n373 163.367
R620 B.n627 B.n626 163.367
R621 B.n626 B.n23 163.367
R622 B.n622 B.n23 163.367
R623 B.n622 B.n621 163.367
R624 B.n621 B.n620 163.367
R625 B.n620 B.n25 163.367
R626 B.n616 B.n25 163.367
R627 B.n616 B.n615 163.367
R628 B.n615 B.n614 163.367
R629 B.n614 B.n27 163.367
R630 B.n610 B.n27 163.367
R631 B.n610 B.n609 163.367
R632 B.n609 B.n608 163.367
R633 B.n608 B.n29 163.367
R634 B.n604 B.n29 163.367
R635 B.n604 B.n603 163.367
R636 B.n603 B.n602 163.367
R637 B.n602 B.n31 163.367
R638 B.n598 B.n31 163.367
R639 B.n598 B.n597 163.367
R640 B.n597 B.n596 163.367
R641 B.n596 B.n33 163.367
R642 B.n592 B.n33 163.367
R643 B.n592 B.n591 163.367
R644 B.n591 B.n590 163.367
R645 B.n590 B.n35 163.367
R646 B.n586 B.n35 163.367
R647 B.n586 B.n585 163.367
R648 B.n585 B.n584 163.367
R649 B.n584 B.n37 163.367
R650 B.n580 B.n37 163.367
R651 B.n580 B.n579 163.367
R652 B.n579 B.n578 163.367
R653 B.n578 B.n39 163.367
R654 B.n574 B.n39 163.367
R655 B.n574 B.n573 163.367
R656 B.n573 B.n572 163.367
R657 B.n572 B.n41 163.367
R658 B.n567 B.n41 163.367
R659 B.n567 B.n566 163.367
R660 B.n566 B.n565 163.367
R661 B.n565 B.n45 163.367
R662 B.n561 B.n45 163.367
R663 B.n561 B.n560 163.367
R664 B.n560 B.n559 163.367
R665 B.n559 B.n47 163.367
R666 B.n555 B.n47 163.367
R667 B.n555 B.n554 163.367
R668 B.n554 B.n553 163.367
R669 B.n553 B.n49 163.367
R670 B.n549 B.n49 163.367
R671 B.n549 B.n548 163.367
R672 B.n548 B.n547 163.367
R673 B.n547 B.n54 163.367
R674 B.n543 B.n54 163.367
R675 B.n543 B.n542 163.367
R676 B.n542 B.n541 163.367
R677 B.n541 B.n56 163.367
R678 B.n537 B.n56 163.367
R679 B.n537 B.n536 163.367
R680 B.n536 B.n535 163.367
R681 B.n535 B.n58 163.367
R682 B.n531 B.n58 163.367
R683 B.n531 B.n530 163.367
R684 B.n530 B.n529 163.367
R685 B.n529 B.n60 163.367
R686 B.n525 B.n60 163.367
R687 B.n525 B.n524 163.367
R688 B.n524 B.n523 163.367
R689 B.n523 B.n62 163.367
R690 B.n519 B.n62 163.367
R691 B.n519 B.n518 163.367
R692 B.n518 B.n517 163.367
R693 B.n517 B.n64 163.367
R694 B.n513 B.n64 163.367
R695 B.n513 B.n512 163.367
R696 B.n512 B.n511 163.367
R697 B.n511 B.n66 163.367
R698 B.n507 B.n66 163.367
R699 B.n507 B.n506 163.367
R700 B.n506 B.n505 163.367
R701 B.n505 B.n68 163.367
R702 B.n501 B.n68 163.367
R703 B.n501 B.n500 163.367
R704 B.n500 B.n499 163.367
R705 B.n499 B.n70 163.367
R706 B.n495 B.n70 163.367
R707 B.n628 B.n21 163.367
R708 B.n632 B.n21 163.367
R709 B.n633 B.n632 163.367
R710 B.n634 B.n633 163.367
R711 B.n634 B.n19 163.367
R712 B.n638 B.n19 163.367
R713 B.n639 B.n638 163.367
R714 B.n640 B.n639 163.367
R715 B.n640 B.n17 163.367
R716 B.n644 B.n17 163.367
R717 B.n645 B.n644 163.367
R718 B.n646 B.n645 163.367
R719 B.n646 B.n15 163.367
R720 B.n650 B.n15 163.367
R721 B.n651 B.n650 163.367
R722 B.n652 B.n651 163.367
R723 B.n652 B.n13 163.367
R724 B.n656 B.n13 163.367
R725 B.n657 B.n656 163.367
R726 B.n658 B.n657 163.367
R727 B.n658 B.n11 163.367
R728 B.n662 B.n11 163.367
R729 B.n663 B.n662 163.367
R730 B.n664 B.n663 163.367
R731 B.n664 B.n9 163.367
R732 B.n668 B.n9 163.367
R733 B.n669 B.n668 163.367
R734 B.n670 B.n669 163.367
R735 B.n670 B.n7 163.367
R736 B.n674 B.n7 163.367
R737 B.n675 B.n674 163.367
R738 B.n676 B.n675 163.367
R739 B.n676 B.n5 163.367
R740 B.n680 B.n5 163.367
R741 B.n681 B.n680 163.367
R742 B.n682 B.n681 163.367
R743 B.n682 B.n3 163.367
R744 B.n686 B.n3 163.367
R745 B.n687 B.n686 163.367
R746 B.n178 B.n2 163.367
R747 B.n179 B.n178 163.367
R748 B.n179 B.n176 163.367
R749 B.n183 B.n176 163.367
R750 B.n184 B.n183 163.367
R751 B.n185 B.n184 163.367
R752 B.n185 B.n174 163.367
R753 B.n189 B.n174 163.367
R754 B.n190 B.n189 163.367
R755 B.n191 B.n190 163.367
R756 B.n191 B.n172 163.367
R757 B.n195 B.n172 163.367
R758 B.n196 B.n195 163.367
R759 B.n197 B.n196 163.367
R760 B.n197 B.n170 163.367
R761 B.n201 B.n170 163.367
R762 B.n202 B.n201 163.367
R763 B.n203 B.n202 163.367
R764 B.n203 B.n168 163.367
R765 B.n207 B.n168 163.367
R766 B.n208 B.n207 163.367
R767 B.n209 B.n208 163.367
R768 B.n209 B.n166 163.367
R769 B.n213 B.n166 163.367
R770 B.n214 B.n213 163.367
R771 B.n215 B.n214 163.367
R772 B.n215 B.n164 163.367
R773 B.n219 B.n164 163.367
R774 B.n220 B.n219 163.367
R775 B.n221 B.n220 163.367
R776 B.n221 B.n162 163.367
R777 B.n225 B.n162 163.367
R778 B.n226 B.n225 163.367
R779 B.n227 B.n226 163.367
R780 B.n227 B.n160 163.367
R781 B.n231 B.n160 163.367
R782 B.n232 B.n231 163.367
R783 B.n233 B.n232 163.367
R784 B.n233 B.n158 163.367
R785 B.n310 B.t8 112.555
R786 B.n51 B.t4 112.555
R787 B.n138 B.t11 112.543
R788 B.n43 B.t1 112.543
R789 B.n295 B.n138 59.5399
R790 B.n311 B.n310 59.5399
R791 B.n52 B.n51 59.5399
R792 B.n569 B.n43 59.5399
R793 B.n138 B.n137 53.3338
R794 B.n310 B.n309 53.3338
R795 B.n51 B.n50 53.3338
R796 B.n43 B.n42 53.3338
R797 B.n629 B.n22 31.0639
R798 B.n496 B.n71 31.0639
R799 B.n372 B.n371 31.0639
R800 B.n236 B.n235 31.0639
R801 B B.n689 18.0485
R802 B.n630 B.n629 10.6151
R803 B.n631 B.n630 10.6151
R804 B.n631 B.n20 10.6151
R805 B.n635 B.n20 10.6151
R806 B.n636 B.n635 10.6151
R807 B.n637 B.n636 10.6151
R808 B.n637 B.n18 10.6151
R809 B.n641 B.n18 10.6151
R810 B.n642 B.n641 10.6151
R811 B.n643 B.n642 10.6151
R812 B.n643 B.n16 10.6151
R813 B.n647 B.n16 10.6151
R814 B.n648 B.n647 10.6151
R815 B.n649 B.n648 10.6151
R816 B.n649 B.n14 10.6151
R817 B.n653 B.n14 10.6151
R818 B.n654 B.n653 10.6151
R819 B.n655 B.n654 10.6151
R820 B.n655 B.n12 10.6151
R821 B.n659 B.n12 10.6151
R822 B.n660 B.n659 10.6151
R823 B.n661 B.n660 10.6151
R824 B.n661 B.n10 10.6151
R825 B.n665 B.n10 10.6151
R826 B.n666 B.n665 10.6151
R827 B.n667 B.n666 10.6151
R828 B.n667 B.n8 10.6151
R829 B.n671 B.n8 10.6151
R830 B.n672 B.n671 10.6151
R831 B.n673 B.n672 10.6151
R832 B.n673 B.n6 10.6151
R833 B.n677 B.n6 10.6151
R834 B.n678 B.n677 10.6151
R835 B.n679 B.n678 10.6151
R836 B.n679 B.n4 10.6151
R837 B.n683 B.n4 10.6151
R838 B.n684 B.n683 10.6151
R839 B.n685 B.n684 10.6151
R840 B.n685 B.n0 10.6151
R841 B.n625 B.n22 10.6151
R842 B.n625 B.n624 10.6151
R843 B.n624 B.n623 10.6151
R844 B.n623 B.n24 10.6151
R845 B.n619 B.n24 10.6151
R846 B.n619 B.n618 10.6151
R847 B.n618 B.n617 10.6151
R848 B.n617 B.n26 10.6151
R849 B.n613 B.n26 10.6151
R850 B.n613 B.n612 10.6151
R851 B.n612 B.n611 10.6151
R852 B.n611 B.n28 10.6151
R853 B.n607 B.n28 10.6151
R854 B.n607 B.n606 10.6151
R855 B.n606 B.n605 10.6151
R856 B.n605 B.n30 10.6151
R857 B.n601 B.n30 10.6151
R858 B.n601 B.n600 10.6151
R859 B.n600 B.n599 10.6151
R860 B.n599 B.n32 10.6151
R861 B.n595 B.n32 10.6151
R862 B.n595 B.n594 10.6151
R863 B.n594 B.n593 10.6151
R864 B.n593 B.n34 10.6151
R865 B.n589 B.n34 10.6151
R866 B.n589 B.n588 10.6151
R867 B.n588 B.n587 10.6151
R868 B.n587 B.n36 10.6151
R869 B.n583 B.n36 10.6151
R870 B.n583 B.n582 10.6151
R871 B.n582 B.n581 10.6151
R872 B.n581 B.n38 10.6151
R873 B.n577 B.n38 10.6151
R874 B.n577 B.n576 10.6151
R875 B.n576 B.n575 10.6151
R876 B.n575 B.n40 10.6151
R877 B.n571 B.n40 10.6151
R878 B.n571 B.n570 10.6151
R879 B.n568 B.n44 10.6151
R880 B.n564 B.n44 10.6151
R881 B.n564 B.n563 10.6151
R882 B.n563 B.n562 10.6151
R883 B.n562 B.n46 10.6151
R884 B.n558 B.n46 10.6151
R885 B.n558 B.n557 10.6151
R886 B.n557 B.n556 10.6151
R887 B.n556 B.n48 10.6151
R888 B.n552 B.n551 10.6151
R889 B.n551 B.n550 10.6151
R890 B.n550 B.n53 10.6151
R891 B.n546 B.n53 10.6151
R892 B.n546 B.n545 10.6151
R893 B.n545 B.n544 10.6151
R894 B.n544 B.n55 10.6151
R895 B.n540 B.n55 10.6151
R896 B.n540 B.n539 10.6151
R897 B.n539 B.n538 10.6151
R898 B.n538 B.n57 10.6151
R899 B.n534 B.n57 10.6151
R900 B.n534 B.n533 10.6151
R901 B.n533 B.n532 10.6151
R902 B.n532 B.n59 10.6151
R903 B.n528 B.n59 10.6151
R904 B.n528 B.n527 10.6151
R905 B.n527 B.n526 10.6151
R906 B.n526 B.n61 10.6151
R907 B.n522 B.n61 10.6151
R908 B.n522 B.n521 10.6151
R909 B.n521 B.n520 10.6151
R910 B.n520 B.n63 10.6151
R911 B.n516 B.n63 10.6151
R912 B.n516 B.n515 10.6151
R913 B.n515 B.n514 10.6151
R914 B.n514 B.n65 10.6151
R915 B.n510 B.n65 10.6151
R916 B.n510 B.n509 10.6151
R917 B.n509 B.n508 10.6151
R918 B.n508 B.n67 10.6151
R919 B.n504 B.n67 10.6151
R920 B.n504 B.n503 10.6151
R921 B.n503 B.n502 10.6151
R922 B.n502 B.n69 10.6151
R923 B.n498 B.n69 10.6151
R924 B.n498 B.n497 10.6151
R925 B.n497 B.n496 10.6151
R926 B.n492 B.n71 10.6151
R927 B.n492 B.n491 10.6151
R928 B.n491 B.n490 10.6151
R929 B.n490 B.n73 10.6151
R930 B.n486 B.n73 10.6151
R931 B.n486 B.n485 10.6151
R932 B.n485 B.n484 10.6151
R933 B.n484 B.n75 10.6151
R934 B.n480 B.n75 10.6151
R935 B.n480 B.n479 10.6151
R936 B.n479 B.n478 10.6151
R937 B.n478 B.n77 10.6151
R938 B.n474 B.n77 10.6151
R939 B.n474 B.n473 10.6151
R940 B.n473 B.n472 10.6151
R941 B.n472 B.n79 10.6151
R942 B.n468 B.n79 10.6151
R943 B.n468 B.n467 10.6151
R944 B.n467 B.n466 10.6151
R945 B.n466 B.n81 10.6151
R946 B.n462 B.n81 10.6151
R947 B.n462 B.n461 10.6151
R948 B.n461 B.n460 10.6151
R949 B.n460 B.n83 10.6151
R950 B.n456 B.n83 10.6151
R951 B.n456 B.n455 10.6151
R952 B.n455 B.n454 10.6151
R953 B.n454 B.n85 10.6151
R954 B.n450 B.n85 10.6151
R955 B.n450 B.n449 10.6151
R956 B.n449 B.n448 10.6151
R957 B.n448 B.n87 10.6151
R958 B.n444 B.n87 10.6151
R959 B.n444 B.n443 10.6151
R960 B.n443 B.n442 10.6151
R961 B.n442 B.n89 10.6151
R962 B.n438 B.n89 10.6151
R963 B.n438 B.n437 10.6151
R964 B.n437 B.n436 10.6151
R965 B.n436 B.n91 10.6151
R966 B.n432 B.n91 10.6151
R967 B.n432 B.n431 10.6151
R968 B.n431 B.n430 10.6151
R969 B.n430 B.n93 10.6151
R970 B.n426 B.n93 10.6151
R971 B.n426 B.n425 10.6151
R972 B.n425 B.n424 10.6151
R973 B.n424 B.n95 10.6151
R974 B.n420 B.n95 10.6151
R975 B.n420 B.n419 10.6151
R976 B.n419 B.n418 10.6151
R977 B.n418 B.n97 10.6151
R978 B.n414 B.n97 10.6151
R979 B.n414 B.n413 10.6151
R980 B.n413 B.n412 10.6151
R981 B.n412 B.n99 10.6151
R982 B.n408 B.n99 10.6151
R983 B.n408 B.n407 10.6151
R984 B.n407 B.n406 10.6151
R985 B.n406 B.n101 10.6151
R986 B.n402 B.n101 10.6151
R987 B.n402 B.n401 10.6151
R988 B.n401 B.n400 10.6151
R989 B.n400 B.n103 10.6151
R990 B.n396 B.n103 10.6151
R991 B.n396 B.n395 10.6151
R992 B.n395 B.n394 10.6151
R993 B.n394 B.n105 10.6151
R994 B.n390 B.n105 10.6151
R995 B.n390 B.n389 10.6151
R996 B.n389 B.n388 10.6151
R997 B.n388 B.n107 10.6151
R998 B.n384 B.n107 10.6151
R999 B.n384 B.n383 10.6151
R1000 B.n383 B.n382 10.6151
R1001 B.n382 B.n109 10.6151
R1002 B.n378 B.n109 10.6151
R1003 B.n378 B.n377 10.6151
R1004 B.n377 B.n376 10.6151
R1005 B.n376 B.n111 10.6151
R1006 B.n372 B.n111 10.6151
R1007 B.n177 B.n1 10.6151
R1008 B.n180 B.n177 10.6151
R1009 B.n181 B.n180 10.6151
R1010 B.n182 B.n181 10.6151
R1011 B.n182 B.n175 10.6151
R1012 B.n186 B.n175 10.6151
R1013 B.n187 B.n186 10.6151
R1014 B.n188 B.n187 10.6151
R1015 B.n188 B.n173 10.6151
R1016 B.n192 B.n173 10.6151
R1017 B.n193 B.n192 10.6151
R1018 B.n194 B.n193 10.6151
R1019 B.n194 B.n171 10.6151
R1020 B.n198 B.n171 10.6151
R1021 B.n199 B.n198 10.6151
R1022 B.n200 B.n199 10.6151
R1023 B.n200 B.n169 10.6151
R1024 B.n204 B.n169 10.6151
R1025 B.n205 B.n204 10.6151
R1026 B.n206 B.n205 10.6151
R1027 B.n206 B.n167 10.6151
R1028 B.n210 B.n167 10.6151
R1029 B.n211 B.n210 10.6151
R1030 B.n212 B.n211 10.6151
R1031 B.n212 B.n165 10.6151
R1032 B.n216 B.n165 10.6151
R1033 B.n217 B.n216 10.6151
R1034 B.n218 B.n217 10.6151
R1035 B.n218 B.n163 10.6151
R1036 B.n222 B.n163 10.6151
R1037 B.n223 B.n222 10.6151
R1038 B.n224 B.n223 10.6151
R1039 B.n224 B.n161 10.6151
R1040 B.n228 B.n161 10.6151
R1041 B.n229 B.n228 10.6151
R1042 B.n230 B.n229 10.6151
R1043 B.n230 B.n159 10.6151
R1044 B.n234 B.n159 10.6151
R1045 B.n235 B.n234 10.6151
R1046 B.n236 B.n157 10.6151
R1047 B.n240 B.n157 10.6151
R1048 B.n241 B.n240 10.6151
R1049 B.n242 B.n241 10.6151
R1050 B.n242 B.n155 10.6151
R1051 B.n246 B.n155 10.6151
R1052 B.n247 B.n246 10.6151
R1053 B.n248 B.n247 10.6151
R1054 B.n248 B.n153 10.6151
R1055 B.n252 B.n153 10.6151
R1056 B.n253 B.n252 10.6151
R1057 B.n254 B.n253 10.6151
R1058 B.n254 B.n151 10.6151
R1059 B.n258 B.n151 10.6151
R1060 B.n259 B.n258 10.6151
R1061 B.n260 B.n259 10.6151
R1062 B.n260 B.n149 10.6151
R1063 B.n264 B.n149 10.6151
R1064 B.n265 B.n264 10.6151
R1065 B.n266 B.n265 10.6151
R1066 B.n266 B.n147 10.6151
R1067 B.n270 B.n147 10.6151
R1068 B.n271 B.n270 10.6151
R1069 B.n272 B.n271 10.6151
R1070 B.n272 B.n145 10.6151
R1071 B.n276 B.n145 10.6151
R1072 B.n277 B.n276 10.6151
R1073 B.n278 B.n277 10.6151
R1074 B.n278 B.n143 10.6151
R1075 B.n282 B.n143 10.6151
R1076 B.n283 B.n282 10.6151
R1077 B.n284 B.n283 10.6151
R1078 B.n284 B.n141 10.6151
R1079 B.n288 B.n141 10.6151
R1080 B.n289 B.n288 10.6151
R1081 B.n290 B.n289 10.6151
R1082 B.n290 B.n139 10.6151
R1083 B.n294 B.n139 10.6151
R1084 B.n297 B.n296 10.6151
R1085 B.n297 B.n135 10.6151
R1086 B.n301 B.n135 10.6151
R1087 B.n302 B.n301 10.6151
R1088 B.n303 B.n302 10.6151
R1089 B.n303 B.n133 10.6151
R1090 B.n307 B.n133 10.6151
R1091 B.n308 B.n307 10.6151
R1092 B.n312 B.n308 10.6151
R1093 B.n316 B.n131 10.6151
R1094 B.n317 B.n316 10.6151
R1095 B.n318 B.n317 10.6151
R1096 B.n318 B.n129 10.6151
R1097 B.n322 B.n129 10.6151
R1098 B.n323 B.n322 10.6151
R1099 B.n324 B.n323 10.6151
R1100 B.n324 B.n127 10.6151
R1101 B.n328 B.n127 10.6151
R1102 B.n329 B.n328 10.6151
R1103 B.n330 B.n329 10.6151
R1104 B.n330 B.n125 10.6151
R1105 B.n334 B.n125 10.6151
R1106 B.n335 B.n334 10.6151
R1107 B.n336 B.n335 10.6151
R1108 B.n336 B.n123 10.6151
R1109 B.n340 B.n123 10.6151
R1110 B.n341 B.n340 10.6151
R1111 B.n342 B.n341 10.6151
R1112 B.n342 B.n121 10.6151
R1113 B.n346 B.n121 10.6151
R1114 B.n347 B.n346 10.6151
R1115 B.n348 B.n347 10.6151
R1116 B.n348 B.n119 10.6151
R1117 B.n352 B.n119 10.6151
R1118 B.n353 B.n352 10.6151
R1119 B.n354 B.n353 10.6151
R1120 B.n354 B.n117 10.6151
R1121 B.n358 B.n117 10.6151
R1122 B.n359 B.n358 10.6151
R1123 B.n360 B.n359 10.6151
R1124 B.n360 B.n115 10.6151
R1125 B.n364 B.n115 10.6151
R1126 B.n365 B.n364 10.6151
R1127 B.n366 B.n365 10.6151
R1128 B.n366 B.n113 10.6151
R1129 B.n370 B.n113 10.6151
R1130 B.n371 B.n370 10.6151
R1131 B.n570 B.n569 9.36635
R1132 B.n552 B.n52 9.36635
R1133 B.n295 B.n294 9.36635
R1134 B.n311 B.n131 9.36635
R1135 B.n689 B.n0 8.11757
R1136 B.n689 B.n1 8.11757
R1137 B.n569 B.n568 1.24928
R1138 B.n52 B.n48 1.24928
R1139 B.n296 B.n295 1.24928
R1140 B.n312 B.n311 1.24928
R1141 VN.n25 VN.n14 161.3
R1142 VN.n24 VN.n23 161.3
R1143 VN.n22 VN.n15 161.3
R1144 VN.n21 VN.n20 161.3
R1145 VN.n19 VN.n16 161.3
R1146 VN.n11 VN.n0 161.3
R1147 VN.n10 VN.n9 161.3
R1148 VN.n8 VN.n1 161.3
R1149 VN.n7 VN.n6 161.3
R1150 VN.n5 VN.n2 161.3
R1151 VN.n3 VN.t2 145.423
R1152 VN.n17 VN.t3 145.423
R1153 VN.n4 VN.t4 111.04
R1154 VN.n12 VN.t1 111.04
R1155 VN.n18 VN.t5 111.04
R1156 VN.n26 VN.t0 111.04
R1157 VN.n13 VN.n12 98.5229
R1158 VN.n27 VN.n26 98.5229
R1159 VN.n6 VN.n1 52.6342
R1160 VN.n20 VN.n15 52.6342
R1161 VN.n4 VN.n3 48.0049
R1162 VN.n18 VN.n17 48.0049
R1163 VN VN.n27 47.6156
R1164 VN.n10 VN.n1 28.3526
R1165 VN.n24 VN.n15 28.3526
R1166 VN.n5 VN.n4 24.4675
R1167 VN.n6 VN.n5 24.4675
R1168 VN.n11 VN.n10 24.4675
R1169 VN.n20 VN.n19 24.4675
R1170 VN.n19 VN.n18 24.4675
R1171 VN.n25 VN.n24 24.4675
R1172 VN.n12 VN.n11 12.234
R1173 VN.n26 VN.n25 12.234
R1174 VN.n17 VN.n16 6.69041
R1175 VN.n3 VN.n2 6.69041
R1176 VN.n27 VN.n14 0.278367
R1177 VN.n13 VN.n0 0.278367
R1178 VN.n23 VN.n14 0.189894
R1179 VN.n23 VN.n22 0.189894
R1180 VN.n22 VN.n21 0.189894
R1181 VN.n21 VN.n16 0.189894
R1182 VN.n7 VN.n2 0.189894
R1183 VN.n8 VN.n7 0.189894
R1184 VN.n9 VN.n8 0.189894
R1185 VN.n9 VN.n0 0.189894
R1186 VN VN.n13 0.153454
R1187 VDD2.n1 VDD2.t3 82.0761
R1188 VDD2.n2 VDD2.t5 80.3536
R1189 VDD2.n1 VDD2.n0 77.9755
R1190 VDD2 VDD2.n3 77.9727
R1191 VDD2.n2 VDD2.n1 41.0321
R1192 VDD2.n3 VDD2.t0 2.91575
R1193 VDD2.n3 VDD2.t2 2.91575
R1194 VDD2.n0 VDD2.t1 2.91575
R1195 VDD2.n0 VDD2.t4 2.91575
R1196 VDD2 VDD2.n2 1.83671
C0 VDD1 VDD2 1.33679f
C1 VDD2 VP 0.442995f
C2 B VTAIL 3.4315f
C3 VTAIL w_n3170_n3198# 2.84202f
C4 B VDD1 1.97939f
C5 VDD1 w_n3170_n3198# 2.18873f
C6 B VP 1.8017f
C7 w_n3170_n3198# VP 6.35469f
C8 VN VTAIL 6.33844f
C9 B VDD2 2.04917f
C10 VDD2 w_n3170_n3198# 2.26808f
C11 VN VDD1 0.150492f
C12 VN VP 6.59454f
C13 VN VDD2 6.18628f
C14 B w_n3170_n3198# 9.189111f
C15 VDD1 VTAIL 7.38994f
C16 VTAIL VP 6.35273f
C17 VDD2 VTAIL 7.43958f
C18 B VN 1.11918f
C19 VN w_n3170_n3198# 5.94535f
C20 VDD1 VP 6.4757f
C21 VDD2 VSUBS 1.835434f
C22 VDD1 VSUBS 2.191307f
C23 VTAIL VSUBS 1.123398f
C24 VN VSUBS 5.618f
C25 VP VSUBS 2.764218f
C26 B VSUBS 4.38511f
C27 w_n3170_n3198# VSUBS 0.124961p
C28 VDD2.t3 VSUBS 2.52849f
C29 VDD2.t1 VSUBS 0.248317f
C30 VDD2.t4 VSUBS 0.248317f
C31 VDD2.n0 VSUBS 1.92584f
C32 VDD2.n1 VSUBS 3.70081f
C33 VDD2.t5 VSUBS 2.51239f
C34 VDD2.n2 VSUBS 3.31426f
C35 VDD2.t0 VSUBS 0.248317f
C36 VDD2.t2 VSUBS 0.248317f
C37 VDD2.n3 VSUBS 1.92579f
C38 VN.n0 VSUBS 0.042408f
C39 VN.t1 VSUBS 2.35968f
C40 VN.n1 VSUBS 0.033098f
C41 VN.n2 VSUBS 0.305109f
C42 VN.t4 VSUBS 2.35968f
C43 VN.t2 VSUBS 2.60375f
C44 VN.n3 VSUBS 0.901983f
C45 VN.n4 VSUBS 0.946757f
C46 VN.n5 VSUBS 0.05995f
C47 VN.n6 VSUBS 0.057416f
C48 VN.n7 VSUBS 0.032166f
C49 VN.n8 VSUBS 0.032166f
C50 VN.n9 VSUBS 0.032166f
C51 VN.n10 VSUBS 0.063357f
C52 VN.n11 VSUBS 0.045152f
C53 VN.n12 VSUBS 0.944442f
C54 VN.n13 VSUBS 0.048744f
C55 VN.n14 VSUBS 0.042408f
C56 VN.t0 VSUBS 2.35968f
C57 VN.n15 VSUBS 0.033098f
C58 VN.n16 VSUBS 0.305109f
C59 VN.t5 VSUBS 2.35968f
C60 VN.t3 VSUBS 2.60375f
C61 VN.n17 VSUBS 0.901983f
C62 VN.n18 VSUBS 0.946757f
C63 VN.n19 VSUBS 0.05995f
C64 VN.n20 VSUBS 0.057416f
C65 VN.n21 VSUBS 0.032166f
C66 VN.n22 VSUBS 0.032166f
C67 VN.n23 VSUBS 0.032166f
C68 VN.n24 VSUBS 0.063357f
C69 VN.n25 VSUBS 0.045152f
C70 VN.n26 VSUBS 0.944442f
C71 VN.n27 VSUBS 1.66332f
C72 B.n0 VSUBS 0.006483f
C73 B.n1 VSUBS 0.006483f
C74 B.n2 VSUBS 0.009588f
C75 B.n3 VSUBS 0.007348f
C76 B.n4 VSUBS 0.007348f
C77 B.n5 VSUBS 0.007348f
C78 B.n6 VSUBS 0.007348f
C79 B.n7 VSUBS 0.007348f
C80 B.n8 VSUBS 0.007348f
C81 B.n9 VSUBS 0.007348f
C82 B.n10 VSUBS 0.007348f
C83 B.n11 VSUBS 0.007348f
C84 B.n12 VSUBS 0.007348f
C85 B.n13 VSUBS 0.007348f
C86 B.n14 VSUBS 0.007348f
C87 B.n15 VSUBS 0.007348f
C88 B.n16 VSUBS 0.007348f
C89 B.n17 VSUBS 0.007348f
C90 B.n18 VSUBS 0.007348f
C91 B.n19 VSUBS 0.007348f
C92 B.n20 VSUBS 0.007348f
C93 B.n21 VSUBS 0.007348f
C94 B.n22 VSUBS 0.017119f
C95 B.n23 VSUBS 0.007348f
C96 B.n24 VSUBS 0.007348f
C97 B.n25 VSUBS 0.007348f
C98 B.n26 VSUBS 0.007348f
C99 B.n27 VSUBS 0.007348f
C100 B.n28 VSUBS 0.007348f
C101 B.n29 VSUBS 0.007348f
C102 B.n30 VSUBS 0.007348f
C103 B.n31 VSUBS 0.007348f
C104 B.n32 VSUBS 0.007348f
C105 B.n33 VSUBS 0.007348f
C106 B.n34 VSUBS 0.007348f
C107 B.n35 VSUBS 0.007348f
C108 B.n36 VSUBS 0.007348f
C109 B.n37 VSUBS 0.007348f
C110 B.n38 VSUBS 0.007348f
C111 B.n39 VSUBS 0.007348f
C112 B.n40 VSUBS 0.007348f
C113 B.n41 VSUBS 0.007348f
C114 B.t1 VSUBS 0.378297f
C115 B.t2 VSUBS 0.398886f
C116 B.t0 VSUBS 1.28967f
C117 B.n42 VSUBS 0.2057f
C118 B.n43 VSUBS 0.074515f
C119 B.n44 VSUBS 0.007348f
C120 B.n45 VSUBS 0.007348f
C121 B.n46 VSUBS 0.007348f
C122 B.n47 VSUBS 0.007348f
C123 B.n48 VSUBS 0.004106f
C124 B.n49 VSUBS 0.007348f
C125 B.t4 VSUBS 0.378291f
C126 B.t5 VSUBS 0.39888f
C127 B.t3 VSUBS 1.28967f
C128 B.n50 VSUBS 0.205706f
C129 B.n51 VSUBS 0.074521f
C130 B.n52 VSUBS 0.017024f
C131 B.n53 VSUBS 0.007348f
C132 B.n54 VSUBS 0.007348f
C133 B.n55 VSUBS 0.007348f
C134 B.n56 VSUBS 0.007348f
C135 B.n57 VSUBS 0.007348f
C136 B.n58 VSUBS 0.007348f
C137 B.n59 VSUBS 0.007348f
C138 B.n60 VSUBS 0.007348f
C139 B.n61 VSUBS 0.007348f
C140 B.n62 VSUBS 0.007348f
C141 B.n63 VSUBS 0.007348f
C142 B.n64 VSUBS 0.007348f
C143 B.n65 VSUBS 0.007348f
C144 B.n66 VSUBS 0.007348f
C145 B.n67 VSUBS 0.007348f
C146 B.n68 VSUBS 0.007348f
C147 B.n69 VSUBS 0.007348f
C148 B.n70 VSUBS 0.007348f
C149 B.n71 VSUBS 0.016162f
C150 B.n72 VSUBS 0.007348f
C151 B.n73 VSUBS 0.007348f
C152 B.n74 VSUBS 0.007348f
C153 B.n75 VSUBS 0.007348f
C154 B.n76 VSUBS 0.007348f
C155 B.n77 VSUBS 0.007348f
C156 B.n78 VSUBS 0.007348f
C157 B.n79 VSUBS 0.007348f
C158 B.n80 VSUBS 0.007348f
C159 B.n81 VSUBS 0.007348f
C160 B.n82 VSUBS 0.007348f
C161 B.n83 VSUBS 0.007348f
C162 B.n84 VSUBS 0.007348f
C163 B.n85 VSUBS 0.007348f
C164 B.n86 VSUBS 0.007348f
C165 B.n87 VSUBS 0.007348f
C166 B.n88 VSUBS 0.007348f
C167 B.n89 VSUBS 0.007348f
C168 B.n90 VSUBS 0.007348f
C169 B.n91 VSUBS 0.007348f
C170 B.n92 VSUBS 0.007348f
C171 B.n93 VSUBS 0.007348f
C172 B.n94 VSUBS 0.007348f
C173 B.n95 VSUBS 0.007348f
C174 B.n96 VSUBS 0.007348f
C175 B.n97 VSUBS 0.007348f
C176 B.n98 VSUBS 0.007348f
C177 B.n99 VSUBS 0.007348f
C178 B.n100 VSUBS 0.007348f
C179 B.n101 VSUBS 0.007348f
C180 B.n102 VSUBS 0.007348f
C181 B.n103 VSUBS 0.007348f
C182 B.n104 VSUBS 0.007348f
C183 B.n105 VSUBS 0.007348f
C184 B.n106 VSUBS 0.007348f
C185 B.n107 VSUBS 0.007348f
C186 B.n108 VSUBS 0.007348f
C187 B.n109 VSUBS 0.007348f
C188 B.n110 VSUBS 0.007348f
C189 B.n111 VSUBS 0.007348f
C190 B.n112 VSUBS 0.017119f
C191 B.n113 VSUBS 0.007348f
C192 B.n114 VSUBS 0.007348f
C193 B.n115 VSUBS 0.007348f
C194 B.n116 VSUBS 0.007348f
C195 B.n117 VSUBS 0.007348f
C196 B.n118 VSUBS 0.007348f
C197 B.n119 VSUBS 0.007348f
C198 B.n120 VSUBS 0.007348f
C199 B.n121 VSUBS 0.007348f
C200 B.n122 VSUBS 0.007348f
C201 B.n123 VSUBS 0.007348f
C202 B.n124 VSUBS 0.007348f
C203 B.n125 VSUBS 0.007348f
C204 B.n126 VSUBS 0.007348f
C205 B.n127 VSUBS 0.007348f
C206 B.n128 VSUBS 0.007348f
C207 B.n129 VSUBS 0.007348f
C208 B.n130 VSUBS 0.007348f
C209 B.n131 VSUBS 0.006916f
C210 B.n132 VSUBS 0.007348f
C211 B.n133 VSUBS 0.007348f
C212 B.n134 VSUBS 0.007348f
C213 B.n135 VSUBS 0.007348f
C214 B.n136 VSUBS 0.007348f
C215 B.t11 VSUBS 0.378297f
C216 B.t10 VSUBS 0.398886f
C217 B.t9 VSUBS 1.28967f
C218 B.n137 VSUBS 0.2057f
C219 B.n138 VSUBS 0.074515f
C220 B.n139 VSUBS 0.007348f
C221 B.n140 VSUBS 0.007348f
C222 B.n141 VSUBS 0.007348f
C223 B.n142 VSUBS 0.007348f
C224 B.n143 VSUBS 0.007348f
C225 B.n144 VSUBS 0.007348f
C226 B.n145 VSUBS 0.007348f
C227 B.n146 VSUBS 0.007348f
C228 B.n147 VSUBS 0.007348f
C229 B.n148 VSUBS 0.007348f
C230 B.n149 VSUBS 0.007348f
C231 B.n150 VSUBS 0.007348f
C232 B.n151 VSUBS 0.007348f
C233 B.n152 VSUBS 0.007348f
C234 B.n153 VSUBS 0.007348f
C235 B.n154 VSUBS 0.007348f
C236 B.n155 VSUBS 0.007348f
C237 B.n156 VSUBS 0.007348f
C238 B.n157 VSUBS 0.007348f
C239 B.n158 VSUBS 0.016162f
C240 B.n159 VSUBS 0.007348f
C241 B.n160 VSUBS 0.007348f
C242 B.n161 VSUBS 0.007348f
C243 B.n162 VSUBS 0.007348f
C244 B.n163 VSUBS 0.007348f
C245 B.n164 VSUBS 0.007348f
C246 B.n165 VSUBS 0.007348f
C247 B.n166 VSUBS 0.007348f
C248 B.n167 VSUBS 0.007348f
C249 B.n168 VSUBS 0.007348f
C250 B.n169 VSUBS 0.007348f
C251 B.n170 VSUBS 0.007348f
C252 B.n171 VSUBS 0.007348f
C253 B.n172 VSUBS 0.007348f
C254 B.n173 VSUBS 0.007348f
C255 B.n174 VSUBS 0.007348f
C256 B.n175 VSUBS 0.007348f
C257 B.n176 VSUBS 0.007348f
C258 B.n177 VSUBS 0.007348f
C259 B.n178 VSUBS 0.007348f
C260 B.n179 VSUBS 0.007348f
C261 B.n180 VSUBS 0.007348f
C262 B.n181 VSUBS 0.007348f
C263 B.n182 VSUBS 0.007348f
C264 B.n183 VSUBS 0.007348f
C265 B.n184 VSUBS 0.007348f
C266 B.n185 VSUBS 0.007348f
C267 B.n186 VSUBS 0.007348f
C268 B.n187 VSUBS 0.007348f
C269 B.n188 VSUBS 0.007348f
C270 B.n189 VSUBS 0.007348f
C271 B.n190 VSUBS 0.007348f
C272 B.n191 VSUBS 0.007348f
C273 B.n192 VSUBS 0.007348f
C274 B.n193 VSUBS 0.007348f
C275 B.n194 VSUBS 0.007348f
C276 B.n195 VSUBS 0.007348f
C277 B.n196 VSUBS 0.007348f
C278 B.n197 VSUBS 0.007348f
C279 B.n198 VSUBS 0.007348f
C280 B.n199 VSUBS 0.007348f
C281 B.n200 VSUBS 0.007348f
C282 B.n201 VSUBS 0.007348f
C283 B.n202 VSUBS 0.007348f
C284 B.n203 VSUBS 0.007348f
C285 B.n204 VSUBS 0.007348f
C286 B.n205 VSUBS 0.007348f
C287 B.n206 VSUBS 0.007348f
C288 B.n207 VSUBS 0.007348f
C289 B.n208 VSUBS 0.007348f
C290 B.n209 VSUBS 0.007348f
C291 B.n210 VSUBS 0.007348f
C292 B.n211 VSUBS 0.007348f
C293 B.n212 VSUBS 0.007348f
C294 B.n213 VSUBS 0.007348f
C295 B.n214 VSUBS 0.007348f
C296 B.n215 VSUBS 0.007348f
C297 B.n216 VSUBS 0.007348f
C298 B.n217 VSUBS 0.007348f
C299 B.n218 VSUBS 0.007348f
C300 B.n219 VSUBS 0.007348f
C301 B.n220 VSUBS 0.007348f
C302 B.n221 VSUBS 0.007348f
C303 B.n222 VSUBS 0.007348f
C304 B.n223 VSUBS 0.007348f
C305 B.n224 VSUBS 0.007348f
C306 B.n225 VSUBS 0.007348f
C307 B.n226 VSUBS 0.007348f
C308 B.n227 VSUBS 0.007348f
C309 B.n228 VSUBS 0.007348f
C310 B.n229 VSUBS 0.007348f
C311 B.n230 VSUBS 0.007348f
C312 B.n231 VSUBS 0.007348f
C313 B.n232 VSUBS 0.007348f
C314 B.n233 VSUBS 0.007348f
C315 B.n234 VSUBS 0.007348f
C316 B.n235 VSUBS 0.016162f
C317 B.n236 VSUBS 0.017119f
C318 B.n237 VSUBS 0.017119f
C319 B.n238 VSUBS 0.007348f
C320 B.n239 VSUBS 0.007348f
C321 B.n240 VSUBS 0.007348f
C322 B.n241 VSUBS 0.007348f
C323 B.n242 VSUBS 0.007348f
C324 B.n243 VSUBS 0.007348f
C325 B.n244 VSUBS 0.007348f
C326 B.n245 VSUBS 0.007348f
C327 B.n246 VSUBS 0.007348f
C328 B.n247 VSUBS 0.007348f
C329 B.n248 VSUBS 0.007348f
C330 B.n249 VSUBS 0.007348f
C331 B.n250 VSUBS 0.007348f
C332 B.n251 VSUBS 0.007348f
C333 B.n252 VSUBS 0.007348f
C334 B.n253 VSUBS 0.007348f
C335 B.n254 VSUBS 0.007348f
C336 B.n255 VSUBS 0.007348f
C337 B.n256 VSUBS 0.007348f
C338 B.n257 VSUBS 0.007348f
C339 B.n258 VSUBS 0.007348f
C340 B.n259 VSUBS 0.007348f
C341 B.n260 VSUBS 0.007348f
C342 B.n261 VSUBS 0.007348f
C343 B.n262 VSUBS 0.007348f
C344 B.n263 VSUBS 0.007348f
C345 B.n264 VSUBS 0.007348f
C346 B.n265 VSUBS 0.007348f
C347 B.n266 VSUBS 0.007348f
C348 B.n267 VSUBS 0.007348f
C349 B.n268 VSUBS 0.007348f
C350 B.n269 VSUBS 0.007348f
C351 B.n270 VSUBS 0.007348f
C352 B.n271 VSUBS 0.007348f
C353 B.n272 VSUBS 0.007348f
C354 B.n273 VSUBS 0.007348f
C355 B.n274 VSUBS 0.007348f
C356 B.n275 VSUBS 0.007348f
C357 B.n276 VSUBS 0.007348f
C358 B.n277 VSUBS 0.007348f
C359 B.n278 VSUBS 0.007348f
C360 B.n279 VSUBS 0.007348f
C361 B.n280 VSUBS 0.007348f
C362 B.n281 VSUBS 0.007348f
C363 B.n282 VSUBS 0.007348f
C364 B.n283 VSUBS 0.007348f
C365 B.n284 VSUBS 0.007348f
C366 B.n285 VSUBS 0.007348f
C367 B.n286 VSUBS 0.007348f
C368 B.n287 VSUBS 0.007348f
C369 B.n288 VSUBS 0.007348f
C370 B.n289 VSUBS 0.007348f
C371 B.n290 VSUBS 0.007348f
C372 B.n291 VSUBS 0.007348f
C373 B.n292 VSUBS 0.007348f
C374 B.n293 VSUBS 0.007348f
C375 B.n294 VSUBS 0.006916f
C376 B.n295 VSUBS 0.017024f
C377 B.n296 VSUBS 0.004106f
C378 B.n297 VSUBS 0.007348f
C379 B.n298 VSUBS 0.007348f
C380 B.n299 VSUBS 0.007348f
C381 B.n300 VSUBS 0.007348f
C382 B.n301 VSUBS 0.007348f
C383 B.n302 VSUBS 0.007348f
C384 B.n303 VSUBS 0.007348f
C385 B.n304 VSUBS 0.007348f
C386 B.n305 VSUBS 0.007348f
C387 B.n306 VSUBS 0.007348f
C388 B.n307 VSUBS 0.007348f
C389 B.n308 VSUBS 0.007348f
C390 B.t8 VSUBS 0.378291f
C391 B.t7 VSUBS 0.39888f
C392 B.t6 VSUBS 1.28967f
C393 B.n309 VSUBS 0.205706f
C394 B.n310 VSUBS 0.074521f
C395 B.n311 VSUBS 0.017024f
C396 B.n312 VSUBS 0.004106f
C397 B.n313 VSUBS 0.007348f
C398 B.n314 VSUBS 0.007348f
C399 B.n315 VSUBS 0.007348f
C400 B.n316 VSUBS 0.007348f
C401 B.n317 VSUBS 0.007348f
C402 B.n318 VSUBS 0.007348f
C403 B.n319 VSUBS 0.007348f
C404 B.n320 VSUBS 0.007348f
C405 B.n321 VSUBS 0.007348f
C406 B.n322 VSUBS 0.007348f
C407 B.n323 VSUBS 0.007348f
C408 B.n324 VSUBS 0.007348f
C409 B.n325 VSUBS 0.007348f
C410 B.n326 VSUBS 0.007348f
C411 B.n327 VSUBS 0.007348f
C412 B.n328 VSUBS 0.007348f
C413 B.n329 VSUBS 0.007348f
C414 B.n330 VSUBS 0.007348f
C415 B.n331 VSUBS 0.007348f
C416 B.n332 VSUBS 0.007348f
C417 B.n333 VSUBS 0.007348f
C418 B.n334 VSUBS 0.007348f
C419 B.n335 VSUBS 0.007348f
C420 B.n336 VSUBS 0.007348f
C421 B.n337 VSUBS 0.007348f
C422 B.n338 VSUBS 0.007348f
C423 B.n339 VSUBS 0.007348f
C424 B.n340 VSUBS 0.007348f
C425 B.n341 VSUBS 0.007348f
C426 B.n342 VSUBS 0.007348f
C427 B.n343 VSUBS 0.007348f
C428 B.n344 VSUBS 0.007348f
C429 B.n345 VSUBS 0.007348f
C430 B.n346 VSUBS 0.007348f
C431 B.n347 VSUBS 0.007348f
C432 B.n348 VSUBS 0.007348f
C433 B.n349 VSUBS 0.007348f
C434 B.n350 VSUBS 0.007348f
C435 B.n351 VSUBS 0.007348f
C436 B.n352 VSUBS 0.007348f
C437 B.n353 VSUBS 0.007348f
C438 B.n354 VSUBS 0.007348f
C439 B.n355 VSUBS 0.007348f
C440 B.n356 VSUBS 0.007348f
C441 B.n357 VSUBS 0.007348f
C442 B.n358 VSUBS 0.007348f
C443 B.n359 VSUBS 0.007348f
C444 B.n360 VSUBS 0.007348f
C445 B.n361 VSUBS 0.007348f
C446 B.n362 VSUBS 0.007348f
C447 B.n363 VSUBS 0.007348f
C448 B.n364 VSUBS 0.007348f
C449 B.n365 VSUBS 0.007348f
C450 B.n366 VSUBS 0.007348f
C451 B.n367 VSUBS 0.007348f
C452 B.n368 VSUBS 0.007348f
C453 B.n369 VSUBS 0.007348f
C454 B.n370 VSUBS 0.007348f
C455 B.n371 VSUBS 0.016206f
C456 B.n372 VSUBS 0.017075f
C457 B.n373 VSUBS 0.016162f
C458 B.n374 VSUBS 0.007348f
C459 B.n375 VSUBS 0.007348f
C460 B.n376 VSUBS 0.007348f
C461 B.n377 VSUBS 0.007348f
C462 B.n378 VSUBS 0.007348f
C463 B.n379 VSUBS 0.007348f
C464 B.n380 VSUBS 0.007348f
C465 B.n381 VSUBS 0.007348f
C466 B.n382 VSUBS 0.007348f
C467 B.n383 VSUBS 0.007348f
C468 B.n384 VSUBS 0.007348f
C469 B.n385 VSUBS 0.007348f
C470 B.n386 VSUBS 0.007348f
C471 B.n387 VSUBS 0.007348f
C472 B.n388 VSUBS 0.007348f
C473 B.n389 VSUBS 0.007348f
C474 B.n390 VSUBS 0.007348f
C475 B.n391 VSUBS 0.007348f
C476 B.n392 VSUBS 0.007348f
C477 B.n393 VSUBS 0.007348f
C478 B.n394 VSUBS 0.007348f
C479 B.n395 VSUBS 0.007348f
C480 B.n396 VSUBS 0.007348f
C481 B.n397 VSUBS 0.007348f
C482 B.n398 VSUBS 0.007348f
C483 B.n399 VSUBS 0.007348f
C484 B.n400 VSUBS 0.007348f
C485 B.n401 VSUBS 0.007348f
C486 B.n402 VSUBS 0.007348f
C487 B.n403 VSUBS 0.007348f
C488 B.n404 VSUBS 0.007348f
C489 B.n405 VSUBS 0.007348f
C490 B.n406 VSUBS 0.007348f
C491 B.n407 VSUBS 0.007348f
C492 B.n408 VSUBS 0.007348f
C493 B.n409 VSUBS 0.007348f
C494 B.n410 VSUBS 0.007348f
C495 B.n411 VSUBS 0.007348f
C496 B.n412 VSUBS 0.007348f
C497 B.n413 VSUBS 0.007348f
C498 B.n414 VSUBS 0.007348f
C499 B.n415 VSUBS 0.007348f
C500 B.n416 VSUBS 0.007348f
C501 B.n417 VSUBS 0.007348f
C502 B.n418 VSUBS 0.007348f
C503 B.n419 VSUBS 0.007348f
C504 B.n420 VSUBS 0.007348f
C505 B.n421 VSUBS 0.007348f
C506 B.n422 VSUBS 0.007348f
C507 B.n423 VSUBS 0.007348f
C508 B.n424 VSUBS 0.007348f
C509 B.n425 VSUBS 0.007348f
C510 B.n426 VSUBS 0.007348f
C511 B.n427 VSUBS 0.007348f
C512 B.n428 VSUBS 0.007348f
C513 B.n429 VSUBS 0.007348f
C514 B.n430 VSUBS 0.007348f
C515 B.n431 VSUBS 0.007348f
C516 B.n432 VSUBS 0.007348f
C517 B.n433 VSUBS 0.007348f
C518 B.n434 VSUBS 0.007348f
C519 B.n435 VSUBS 0.007348f
C520 B.n436 VSUBS 0.007348f
C521 B.n437 VSUBS 0.007348f
C522 B.n438 VSUBS 0.007348f
C523 B.n439 VSUBS 0.007348f
C524 B.n440 VSUBS 0.007348f
C525 B.n441 VSUBS 0.007348f
C526 B.n442 VSUBS 0.007348f
C527 B.n443 VSUBS 0.007348f
C528 B.n444 VSUBS 0.007348f
C529 B.n445 VSUBS 0.007348f
C530 B.n446 VSUBS 0.007348f
C531 B.n447 VSUBS 0.007348f
C532 B.n448 VSUBS 0.007348f
C533 B.n449 VSUBS 0.007348f
C534 B.n450 VSUBS 0.007348f
C535 B.n451 VSUBS 0.007348f
C536 B.n452 VSUBS 0.007348f
C537 B.n453 VSUBS 0.007348f
C538 B.n454 VSUBS 0.007348f
C539 B.n455 VSUBS 0.007348f
C540 B.n456 VSUBS 0.007348f
C541 B.n457 VSUBS 0.007348f
C542 B.n458 VSUBS 0.007348f
C543 B.n459 VSUBS 0.007348f
C544 B.n460 VSUBS 0.007348f
C545 B.n461 VSUBS 0.007348f
C546 B.n462 VSUBS 0.007348f
C547 B.n463 VSUBS 0.007348f
C548 B.n464 VSUBS 0.007348f
C549 B.n465 VSUBS 0.007348f
C550 B.n466 VSUBS 0.007348f
C551 B.n467 VSUBS 0.007348f
C552 B.n468 VSUBS 0.007348f
C553 B.n469 VSUBS 0.007348f
C554 B.n470 VSUBS 0.007348f
C555 B.n471 VSUBS 0.007348f
C556 B.n472 VSUBS 0.007348f
C557 B.n473 VSUBS 0.007348f
C558 B.n474 VSUBS 0.007348f
C559 B.n475 VSUBS 0.007348f
C560 B.n476 VSUBS 0.007348f
C561 B.n477 VSUBS 0.007348f
C562 B.n478 VSUBS 0.007348f
C563 B.n479 VSUBS 0.007348f
C564 B.n480 VSUBS 0.007348f
C565 B.n481 VSUBS 0.007348f
C566 B.n482 VSUBS 0.007348f
C567 B.n483 VSUBS 0.007348f
C568 B.n484 VSUBS 0.007348f
C569 B.n485 VSUBS 0.007348f
C570 B.n486 VSUBS 0.007348f
C571 B.n487 VSUBS 0.007348f
C572 B.n488 VSUBS 0.007348f
C573 B.n489 VSUBS 0.007348f
C574 B.n490 VSUBS 0.007348f
C575 B.n491 VSUBS 0.007348f
C576 B.n492 VSUBS 0.007348f
C577 B.n493 VSUBS 0.007348f
C578 B.n494 VSUBS 0.016162f
C579 B.n495 VSUBS 0.017119f
C580 B.n496 VSUBS 0.017119f
C581 B.n497 VSUBS 0.007348f
C582 B.n498 VSUBS 0.007348f
C583 B.n499 VSUBS 0.007348f
C584 B.n500 VSUBS 0.007348f
C585 B.n501 VSUBS 0.007348f
C586 B.n502 VSUBS 0.007348f
C587 B.n503 VSUBS 0.007348f
C588 B.n504 VSUBS 0.007348f
C589 B.n505 VSUBS 0.007348f
C590 B.n506 VSUBS 0.007348f
C591 B.n507 VSUBS 0.007348f
C592 B.n508 VSUBS 0.007348f
C593 B.n509 VSUBS 0.007348f
C594 B.n510 VSUBS 0.007348f
C595 B.n511 VSUBS 0.007348f
C596 B.n512 VSUBS 0.007348f
C597 B.n513 VSUBS 0.007348f
C598 B.n514 VSUBS 0.007348f
C599 B.n515 VSUBS 0.007348f
C600 B.n516 VSUBS 0.007348f
C601 B.n517 VSUBS 0.007348f
C602 B.n518 VSUBS 0.007348f
C603 B.n519 VSUBS 0.007348f
C604 B.n520 VSUBS 0.007348f
C605 B.n521 VSUBS 0.007348f
C606 B.n522 VSUBS 0.007348f
C607 B.n523 VSUBS 0.007348f
C608 B.n524 VSUBS 0.007348f
C609 B.n525 VSUBS 0.007348f
C610 B.n526 VSUBS 0.007348f
C611 B.n527 VSUBS 0.007348f
C612 B.n528 VSUBS 0.007348f
C613 B.n529 VSUBS 0.007348f
C614 B.n530 VSUBS 0.007348f
C615 B.n531 VSUBS 0.007348f
C616 B.n532 VSUBS 0.007348f
C617 B.n533 VSUBS 0.007348f
C618 B.n534 VSUBS 0.007348f
C619 B.n535 VSUBS 0.007348f
C620 B.n536 VSUBS 0.007348f
C621 B.n537 VSUBS 0.007348f
C622 B.n538 VSUBS 0.007348f
C623 B.n539 VSUBS 0.007348f
C624 B.n540 VSUBS 0.007348f
C625 B.n541 VSUBS 0.007348f
C626 B.n542 VSUBS 0.007348f
C627 B.n543 VSUBS 0.007348f
C628 B.n544 VSUBS 0.007348f
C629 B.n545 VSUBS 0.007348f
C630 B.n546 VSUBS 0.007348f
C631 B.n547 VSUBS 0.007348f
C632 B.n548 VSUBS 0.007348f
C633 B.n549 VSUBS 0.007348f
C634 B.n550 VSUBS 0.007348f
C635 B.n551 VSUBS 0.007348f
C636 B.n552 VSUBS 0.006916f
C637 B.n553 VSUBS 0.007348f
C638 B.n554 VSUBS 0.007348f
C639 B.n555 VSUBS 0.007348f
C640 B.n556 VSUBS 0.007348f
C641 B.n557 VSUBS 0.007348f
C642 B.n558 VSUBS 0.007348f
C643 B.n559 VSUBS 0.007348f
C644 B.n560 VSUBS 0.007348f
C645 B.n561 VSUBS 0.007348f
C646 B.n562 VSUBS 0.007348f
C647 B.n563 VSUBS 0.007348f
C648 B.n564 VSUBS 0.007348f
C649 B.n565 VSUBS 0.007348f
C650 B.n566 VSUBS 0.007348f
C651 B.n567 VSUBS 0.007348f
C652 B.n568 VSUBS 0.004106f
C653 B.n569 VSUBS 0.017024f
C654 B.n570 VSUBS 0.006916f
C655 B.n571 VSUBS 0.007348f
C656 B.n572 VSUBS 0.007348f
C657 B.n573 VSUBS 0.007348f
C658 B.n574 VSUBS 0.007348f
C659 B.n575 VSUBS 0.007348f
C660 B.n576 VSUBS 0.007348f
C661 B.n577 VSUBS 0.007348f
C662 B.n578 VSUBS 0.007348f
C663 B.n579 VSUBS 0.007348f
C664 B.n580 VSUBS 0.007348f
C665 B.n581 VSUBS 0.007348f
C666 B.n582 VSUBS 0.007348f
C667 B.n583 VSUBS 0.007348f
C668 B.n584 VSUBS 0.007348f
C669 B.n585 VSUBS 0.007348f
C670 B.n586 VSUBS 0.007348f
C671 B.n587 VSUBS 0.007348f
C672 B.n588 VSUBS 0.007348f
C673 B.n589 VSUBS 0.007348f
C674 B.n590 VSUBS 0.007348f
C675 B.n591 VSUBS 0.007348f
C676 B.n592 VSUBS 0.007348f
C677 B.n593 VSUBS 0.007348f
C678 B.n594 VSUBS 0.007348f
C679 B.n595 VSUBS 0.007348f
C680 B.n596 VSUBS 0.007348f
C681 B.n597 VSUBS 0.007348f
C682 B.n598 VSUBS 0.007348f
C683 B.n599 VSUBS 0.007348f
C684 B.n600 VSUBS 0.007348f
C685 B.n601 VSUBS 0.007348f
C686 B.n602 VSUBS 0.007348f
C687 B.n603 VSUBS 0.007348f
C688 B.n604 VSUBS 0.007348f
C689 B.n605 VSUBS 0.007348f
C690 B.n606 VSUBS 0.007348f
C691 B.n607 VSUBS 0.007348f
C692 B.n608 VSUBS 0.007348f
C693 B.n609 VSUBS 0.007348f
C694 B.n610 VSUBS 0.007348f
C695 B.n611 VSUBS 0.007348f
C696 B.n612 VSUBS 0.007348f
C697 B.n613 VSUBS 0.007348f
C698 B.n614 VSUBS 0.007348f
C699 B.n615 VSUBS 0.007348f
C700 B.n616 VSUBS 0.007348f
C701 B.n617 VSUBS 0.007348f
C702 B.n618 VSUBS 0.007348f
C703 B.n619 VSUBS 0.007348f
C704 B.n620 VSUBS 0.007348f
C705 B.n621 VSUBS 0.007348f
C706 B.n622 VSUBS 0.007348f
C707 B.n623 VSUBS 0.007348f
C708 B.n624 VSUBS 0.007348f
C709 B.n625 VSUBS 0.007348f
C710 B.n626 VSUBS 0.007348f
C711 B.n627 VSUBS 0.017119f
C712 B.n628 VSUBS 0.016162f
C713 B.n629 VSUBS 0.016162f
C714 B.n630 VSUBS 0.007348f
C715 B.n631 VSUBS 0.007348f
C716 B.n632 VSUBS 0.007348f
C717 B.n633 VSUBS 0.007348f
C718 B.n634 VSUBS 0.007348f
C719 B.n635 VSUBS 0.007348f
C720 B.n636 VSUBS 0.007348f
C721 B.n637 VSUBS 0.007348f
C722 B.n638 VSUBS 0.007348f
C723 B.n639 VSUBS 0.007348f
C724 B.n640 VSUBS 0.007348f
C725 B.n641 VSUBS 0.007348f
C726 B.n642 VSUBS 0.007348f
C727 B.n643 VSUBS 0.007348f
C728 B.n644 VSUBS 0.007348f
C729 B.n645 VSUBS 0.007348f
C730 B.n646 VSUBS 0.007348f
C731 B.n647 VSUBS 0.007348f
C732 B.n648 VSUBS 0.007348f
C733 B.n649 VSUBS 0.007348f
C734 B.n650 VSUBS 0.007348f
C735 B.n651 VSUBS 0.007348f
C736 B.n652 VSUBS 0.007348f
C737 B.n653 VSUBS 0.007348f
C738 B.n654 VSUBS 0.007348f
C739 B.n655 VSUBS 0.007348f
C740 B.n656 VSUBS 0.007348f
C741 B.n657 VSUBS 0.007348f
C742 B.n658 VSUBS 0.007348f
C743 B.n659 VSUBS 0.007348f
C744 B.n660 VSUBS 0.007348f
C745 B.n661 VSUBS 0.007348f
C746 B.n662 VSUBS 0.007348f
C747 B.n663 VSUBS 0.007348f
C748 B.n664 VSUBS 0.007348f
C749 B.n665 VSUBS 0.007348f
C750 B.n666 VSUBS 0.007348f
C751 B.n667 VSUBS 0.007348f
C752 B.n668 VSUBS 0.007348f
C753 B.n669 VSUBS 0.007348f
C754 B.n670 VSUBS 0.007348f
C755 B.n671 VSUBS 0.007348f
C756 B.n672 VSUBS 0.007348f
C757 B.n673 VSUBS 0.007348f
C758 B.n674 VSUBS 0.007348f
C759 B.n675 VSUBS 0.007348f
C760 B.n676 VSUBS 0.007348f
C761 B.n677 VSUBS 0.007348f
C762 B.n678 VSUBS 0.007348f
C763 B.n679 VSUBS 0.007348f
C764 B.n680 VSUBS 0.007348f
C765 B.n681 VSUBS 0.007348f
C766 B.n682 VSUBS 0.007348f
C767 B.n683 VSUBS 0.007348f
C768 B.n684 VSUBS 0.007348f
C769 B.n685 VSUBS 0.007348f
C770 B.n686 VSUBS 0.007348f
C771 B.n687 VSUBS 0.009588f
C772 B.n688 VSUBS 0.010214f
C773 B.n689 VSUBS 0.020312f
C774 VDD1.t5 VSUBS 2.26222f
C775 VDD1.t0 VSUBS 2.26108f
C776 VDD1.t2 VSUBS 0.222056f
C777 VDD1.t4 VSUBS 0.222056f
C778 VDD1.n0 VSUBS 1.72216f
C779 VDD1.n1 VSUBS 3.42918f
C780 VDD1.t3 VSUBS 0.222056f
C781 VDD1.t1 VSUBS 0.222056f
C782 VDD1.n2 VSUBS 1.71729f
C783 VDD1.n3 VSUBS 2.94767f
C784 VTAIL.t3 VSUBS 0.257463f
C785 VTAIL.t1 VSUBS 0.257463f
C786 VTAIL.n0 VSUBS 1.84632f
C787 VTAIL.n1 VSUBS 0.855238f
C788 VTAIL.t5 VSUBS 2.4436f
C789 VTAIL.n2 VSUBS 1.12207f
C790 VTAIL.t7 VSUBS 0.257463f
C791 VTAIL.t10 VSUBS 0.257463f
C792 VTAIL.n3 VSUBS 1.84632f
C793 VTAIL.n4 VSUBS 2.6097f
C794 VTAIL.t0 VSUBS 0.257463f
C795 VTAIL.t2 VSUBS 0.257463f
C796 VTAIL.n5 VSUBS 1.84633f
C797 VTAIL.n6 VSUBS 2.60969f
C798 VTAIL.t11 VSUBS 2.44361f
C799 VTAIL.n7 VSUBS 1.12205f
C800 VTAIL.t8 VSUBS 0.257463f
C801 VTAIL.t9 VSUBS 0.257463f
C802 VTAIL.n8 VSUBS 1.84633f
C803 VTAIL.n9 VSUBS 1.01716f
C804 VTAIL.t6 VSUBS 2.4436f
C805 VTAIL.n10 VSUBS 2.49138f
C806 VTAIL.t4 VSUBS 2.4436f
C807 VTAIL.n11 VSUBS 2.4301f
C808 VP.n0 VSUBS 0.044015f
C809 VP.t1 VSUBS 2.44906f
C810 VP.n1 VSUBS 0.034352f
C811 VP.n2 VSUBS 0.033385f
C812 VP.t3 VSUBS 2.44906f
C813 VP.n3 VSUBS 0.062221f
C814 VP.n4 VSUBS 0.033385f
C815 VP.n5 VSUBS 0.046862f
C816 VP.n6 VSUBS 0.044015f
C817 VP.t4 VSUBS 2.44906f
C818 VP.n7 VSUBS 0.034352f
C819 VP.n8 VSUBS 0.316666f
C820 VP.t2 VSUBS 2.44906f
C821 VP.t0 VSUBS 2.70237f
C822 VP.n9 VSUBS 0.936148f
C823 VP.n10 VSUBS 0.982618f
C824 VP.n11 VSUBS 0.062221f
C825 VP.n12 VSUBS 0.059591f
C826 VP.n13 VSUBS 0.033385f
C827 VP.n14 VSUBS 0.033385f
C828 VP.n15 VSUBS 0.033385f
C829 VP.n16 VSUBS 0.065757f
C830 VP.n17 VSUBS 0.046862f
C831 VP.n18 VSUBS 0.980215f
C832 VP.n19 VSUBS 1.70823f
C833 VP.t5 VSUBS 2.44906f
C834 VP.n20 VSUBS 0.980215f
C835 VP.n21 VSUBS 1.73358f
C836 VP.n22 VSUBS 0.044015f
C837 VP.n23 VSUBS 0.033385f
C838 VP.n24 VSUBS 0.065757f
C839 VP.n25 VSUBS 0.034352f
C840 VP.n26 VSUBS 0.059591f
C841 VP.n27 VSUBS 0.033385f
C842 VP.n28 VSUBS 0.033385f
C843 VP.n29 VSUBS 0.033385f
C844 VP.n30 VSUBS 0.903733f
C845 VP.n31 VSUBS 0.062221f
C846 VP.n32 VSUBS 0.059591f
C847 VP.n33 VSUBS 0.033385f
C848 VP.n34 VSUBS 0.033385f
C849 VP.n35 VSUBS 0.033385f
C850 VP.n36 VSUBS 0.065757f
C851 VP.n37 VSUBS 0.046862f
C852 VP.n38 VSUBS 0.980215f
C853 VP.n39 VSUBS 0.05059f
.ends

