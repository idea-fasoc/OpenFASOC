* NGSPICE file created from diff_pair_sample_1408.ext - technology: sky130A

.subckt diff_pair_sample_1408 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=1.04
X1 B.t8 B.t6 B.t7 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=1.04
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=1.04
X3 VDD1.t1 VP.t0 VTAIL.t3 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=1.04
X4 B.t5 B.t3 B.t4 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=1.04
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=1.04
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0.39 ps=2.78 w=1 l=1.04
X7 B.t2 B.t0 B.t1 w_n1518_n1172# sky130_fd_pr__pfet_01v8 ad=0.39 pd=2.78 as=0 ps=0 w=1 l=1.04
R0 B.n51 B.t8 673.167
R1 B.n57 B.t2 673.167
R2 B.n16 B.t4 673.167
R3 B.n23 B.t10 673.167
R4 B.n52 B.t7 646.596
R5 B.n58 B.t1 646.596
R6 B.n17 B.t5 646.596
R7 B.n24 B.t11 646.596
R8 B.n188 B.n187 585
R9 B.n189 B.n28 585
R10 B.n191 B.n190 585
R11 B.n192 B.n27 585
R12 B.n194 B.n193 585
R13 B.n195 B.n26 585
R14 B.n197 B.n196 585
R15 B.n198 B.n25 585
R16 B.n200 B.n199 585
R17 B.n202 B.n22 585
R18 B.n204 B.n203 585
R19 B.n205 B.n21 585
R20 B.n207 B.n206 585
R21 B.n208 B.n20 585
R22 B.n210 B.n209 585
R23 B.n211 B.n19 585
R24 B.n213 B.n212 585
R25 B.n214 B.n15 585
R26 B.n216 B.n215 585
R27 B.n217 B.n14 585
R28 B.n219 B.n218 585
R29 B.n220 B.n13 585
R30 B.n222 B.n221 585
R31 B.n223 B.n12 585
R32 B.n225 B.n224 585
R33 B.n226 B.n11 585
R34 B.n228 B.n227 585
R35 B.n229 B.n10 585
R36 B.n186 B.n29 585
R37 B.n185 B.n184 585
R38 B.n183 B.n30 585
R39 B.n182 B.n181 585
R40 B.n180 B.n31 585
R41 B.n179 B.n178 585
R42 B.n177 B.n32 585
R43 B.n176 B.n175 585
R44 B.n174 B.n33 585
R45 B.n173 B.n172 585
R46 B.n171 B.n34 585
R47 B.n170 B.n169 585
R48 B.n168 B.n35 585
R49 B.n167 B.n166 585
R50 B.n165 B.n36 585
R51 B.n164 B.n163 585
R52 B.n162 B.n37 585
R53 B.n161 B.n160 585
R54 B.n159 B.n38 585
R55 B.n158 B.n157 585
R56 B.n156 B.n39 585
R57 B.n155 B.n154 585
R58 B.n153 B.n40 585
R59 B.n152 B.n151 585
R60 B.n150 B.n41 585
R61 B.n149 B.n148 585
R62 B.n147 B.n42 585
R63 B.n146 B.n145 585
R64 B.n144 B.n43 585
R65 B.n143 B.n142 585
R66 B.n141 B.n44 585
R67 B.n140 B.n139 585
R68 B.n138 B.n45 585
R69 B.n95 B.n94 585
R70 B.n96 B.n63 585
R71 B.n98 B.n97 585
R72 B.n99 B.n62 585
R73 B.n101 B.n100 585
R74 B.n102 B.n61 585
R75 B.n104 B.n103 585
R76 B.n105 B.n60 585
R77 B.n107 B.n106 585
R78 B.n109 B.n108 585
R79 B.n110 B.n56 585
R80 B.n112 B.n111 585
R81 B.n113 B.n55 585
R82 B.n115 B.n114 585
R83 B.n116 B.n54 585
R84 B.n118 B.n117 585
R85 B.n119 B.n53 585
R86 B.n121 B.n120 585
R87 B.n122 B.n50 585
R88 B.n125 B.n124 585
R89 B.n126 B.n49 585
R90 B.n128 B.n127 585
R91 B.n129 B.n48 585
R92 B.n131 B.n130 585
R93 B.n132 B.n47 585
R94 B.n134 B.n133 585
R95 B.n135 B.n46 585
R96 B.n137 B.n136 585
R97 B.n93 B.n64 585
R98 B.n92 B.n91 585
R99 B.n90 B.n65 585
R100 B.n89 B.n88 585
R101 B.n87 B.n66 585
R102 B.n86 B.n85 585
R103 B.n84 B.n67 585
R104 B.n83 B.n82 585
R105 B.n81 B.n68 585
R106 B.n80 B.n79 585
R107 B.n78 B.n69 585
R108 B.n77 B.n76 585
R109 B.n75 B.n70 585
R110 B.n74 B.n73 585
R111 B.n72 B.n71 585
R112 B.n2 B.n0 585
R113 B.n253 B.n1 585
R114 B.n252 B.n251 585
R115 B.n250 B.n3 585
R116 B.n249 B.n248 585
R117 B.n247 B.n4 585
R118 B.n246 B.n245 585
R119 B.n244 B.n5 585
R120 B.n243 B.n242 585
R121 B.n241 B.n6 585
R122 B.n240 B.n239 585
R123 B.n238 B.n7 585
R124 B.n237 B.n236 585
R125 B.n235 B.n8 585
R126 B.n234 B.n233 585
R127 B.n232 B.n9 585
R128 B.n231 B.n230 585
R129 B.n255 B.n254 585
R130 B.n95 B.n64 545.355
R131 B.n230 B.n229 545.355
R132 B.n138 B.n137 545.355
R133 B.n187 B.n186 545.355
R134 B.n51 B.t6 226.363
R135 B.n57 B.t0 226.363
R136 B.n16 B.t3 226.363
R137 B.n23 B.t9 226.363
R138 B.n91 B.n64 163.367
R139 B.n91 B.n90 163.367
R140 B.n90 B.n89 163.367
R141 B.n89 B.n66 163.367
R142 B.n85 B.n66 163.367
R143 B.n85 B.n84 163.367
R144 B.n84 B.n83 163.367
R145 B.n83 B.n68 163.367
R146 B.n79 B.n68 163.367
R147 B.n79 B.n78 163.367
R148 B.n78 B.n77 163.367
R149 B.n77 B.n70 163.367
R150 B.n73 B.n70 163.367
R151 B.n73 B.n72 163.367
R152 B.n72 B.n2 163.367
R153 B.n254 B.n2 163.367
R154 B.n254 B.n253 163.367
R155 B.n253 B.n252 163.367
R156 B.n252 B.n3 163.367
R157 B.n248 B.n3 163.367
R158 B.n248 B.n247 163.367
R159 B.n247 B.n246 163.367
R160 B.n246 B.n5 163.367
R161 B.n242 B.n5 163.367
R162 B.n242 B.n241 163.367
R163 B.n241 B.n240 163.367
R164 B.n240 B.n7 163.367
R165 B.n236 B.n7 163.367
R166 B.n236 B.n235 163.367
R167 B.n235 B.n234 163.367
R168 B.n234 B.n9 163.367
R169 B.n230 B.n9 163.367
R170 B.n96 B.n95 163.367
R171 B.n97 B.n96 163.367
R172 B.n97 B.n62 163.367
R173 B.n101 B.n62 163.367
R174 B.n102 B.n101 163.367
R175 B.n103 B.n102 163.367
R176 B.n103 B.n60 163.367
R177 B.n107 B.n60 163.367
R178 B.n108 B.n107 163.367
R179 B.n108 B.n56 163.367
R180 B.n112 B.n56 163.367
R181 B.n113 B.n112 163.367
R182 B.n114 B.n113 163.367
R183 B.n114 B.n54 163.367
R184 B.n118 B.n54 163.367
R185 B.n119 B.n118 163.367
R186 B.n120 B.n119 163.367
R187 B.n120 B.n50 163.367
R188 B.n125 B.n50 163.367
R189 B.n126 B.n125 163.367
R190 B.n127 B.n126 163.367
R191 B.n127 B.n48 163.367
R192 B.n131 B.n48 163.367
R193 B.n132 B.n131 163.367
R194 B.n133 B.n132 163.367
R195 B.n133 B.n46 163.367
R196 B.n137 B.n46 163.367
R197 B.n139 B.n138 163.367
R198 B.n139 B.n44 163.367
R199 B.n143 B.n44 163.367
R200 B.n144 B.n143 163.367
R201 B.n145 B.n144 163.367
R202 B.n145 B.n42 163.367
R203 B.n149 B.n42 163.367
R204 B.n150 B.n149 163.367
R205 B.n151 B.n150 163.367
R206 B.n151 B.n40 163.367
R207 B.n155 B.n40 163.367
R208 B.n156 B.n155 163.367
R209 B.n157 B.n156 163.367
R210 B.n157 B.n38 163.367
R211 B.n161 B.n38 163.367
R212 B.n162 B.n161 163.367
R213 B.n163 B.n162 163.367
R214 B.n163 B.n36 163.367
R215 B.n167 B.n36 163.367
R216 B.n168 B.n167 163.367
R217 B.n169 B.n168 163.367
R218 B.n169 B.n34 163.367
R219 B.n173 B.n34 163.367
R220 B.n174 B.n173 163.367
R221 B.n175 B.n174 163.367
R222 B.n175 B.n32 163.367
R223 B.n179 B.n32 163.367
R224 B.n180 B.n179 163.367
R225 B.n181 B.n180 163.367
R226 B.n181 B.n30 163.367
R227 B.n185 B.n30 163.367
R228 B.n186 B.n185 163.367
R229 B.n229 B.n228 163.367
R230 B.n228 B.n11 163.367
R231 B.n224 B.n11 163.367
R232 B.n224 B.n223 163.367
R233 B.n223 B.n222 163.367
R234 B.n222 B.n13 163.367
R235 B.n218 B.n13 163.367
R236 B.n218 B.n217 163.367
R237 B.n217 B.n216 163.367
R238 B.n216 B.n15 163.367
R239 B.n212 B.n15 163.367
R240 B.n212 B.n211 163.367
R241 B.n211 B.n210 163.367
R242 B.n210 B.n20 163.367
R243 B.n206 B.n20 163.367
R244 B.n206 B.n205 163.367
R245 B.n205 B.n204 163.367
R246 B.n204 B.n22 163.367
R247 B.n199 B.n22 163.367
R248 B.n199 B.n198 163.367
R249 B.n198 B.n197 163.367
R250 B.n197 B.n26 163.367
R251 B.n193 B.n26 163.367
R252 B.n193 B.n192 163.367
R253 B.n192 B.n191 163.367
R254 B.n191 B.n28 163.367
R255 B.n187 B.n28 163.367
R256 B.n123 B.n52 59.5399
R257 B.n59 B.n58 59.5399
R258 B.n18 B.n17 59.5399
R259 B.n201 B.n24 59.5399
R260 B.n188 B.n29 35.4346
R261 B.n231 B.n10 35.4346
R262 B.n136 B.n45 35.4346
R263 B.n94 B.n93 35.4346
R264 B.n52 B.n51 26.5702
R265 B.n58 B.n57 26.5702
R266 B.n17 B.n16 26.5702
R267 B.n24 B.n23 26.5702
R268 B B.n255 18.0485
R269 B.n227 B.n10 10.6151
R270 B.n227 B.n226 10.6151
R271 B.n226 B.n225 10.6151
R272 B.n225 B.n12 10.6151
R273 B.n221 B.n12 10.6151
R274 B.n221 B.n220 10.6151
R275 B.n220 B.n219 10.6151
R276 B.n219 B.n14 10.6151
R277 B.n215 B.n214 10.6151
R278 B.n214 B.n213 10.6151
R279 B.n213 B.n19 10.6151
R280 B.n209 B.n19 10.6151
R281 B.n209 B.n208 10.6151
R282 B.n208 B.n207 10.6151
R283 B.n207 B.n21 10.6151
R284 B.n203 B.n21 10.6151
R285 B.n203 B.n202 10.6151
R286 B.n200 B.n25 10.6151
R287 B.n196 B.n25 10.6151
R288 B.n196 B.n195 10.6151
R289 B.n195 B.n194 10.6151
R290 B.n194 B.n27 10.6151
R291 B.n190 B.n27 10.6151
R292 B.n190 B.n189 10.6151
R293 B.n189 B.n188 10.6151
R294 B.n140 B.n45 10.6151
R295 B.n141 B.n140 10.6151
R296 B.n142 B.n141 10.6151
R297 B.n142 B.n43 10.6151
R298 B.n146 B.n43 10.6151
R299 B.n147 B.n146 10.6151
R300 B.n148 B.n147 10.6151
R301 B.n148 B.n41 10.6151
R302 B.n152 B.n41 10.6151
R303 B.n153 B.n152 10.6151
R304 B.n154 B.n153 10.6151
R305 B.n154 B.n39 10.6151
R306 B.n158 B.n39 10.6151
R307 B.n159 B.n158 10.6151
R308 B.n160 B.n159 10.6151
R309 B.n160 B.n37 10.6151
R310 B.n164 B.n37 10.6151
R311 B.n165 B.n164 10.6151
R312 B.n166 B.n165 10.6151
R313 B.n166 B.n35 10.6151
R314 B.n170 B.n35 10.6151
R315 B.n171 B.n170 10.6151
R316 B.n172 B.n171 10.6151
R317 B.n172 B.n33 10.6151
R318 B.n176 B.n33 10.6151
R319 B.n177 B.n176 10.6151
R320 B.n178 B.n177 10.6151
R321 B.n178 B.n31 10.6151
R322 B.n182 B.n31 10.6151
R323 B.n183 B.n182 10.6151
R324 B.n184 B.n183 10.6151
R325 B.n184 B.n29 10.6151
R326 B.n94 B.n63 10.6151
R327 B.n98 B.n63 10.6151
R328 B.n99 B.n98 10.6151
R329 B.n100 B.n99 10.6151
R330 B.n100 B.n61 10.6151
R331 B.n104 B.n61 10.6151
R332 B.n105 B.n104 10.6151
R333 B.n106 B.n105 10.6151
R334 B.n110 B.n109 10.6151
R335 B.n111 B.n110 10.6151
R336 B.n111 B.n55 10.6151
R337 B.n115 B.n55 10.6151
R338 B.n116 B.n115 10.6151
R339 B.n117 B.n116 10.6151
R340 B.n117 B.n53 10.6151
R341 B.n121 B.n53 10.6151
R342 B.n122 B.n121 10.6151
R343 B.n124 B.n49 10.6151
R344 B.n128 B.n49 10.6151
R345 B.n129 B.n128 10.6151
R346 B.n130 B.n129 10.6151
R347 B.n130 B.n47 10.6151
R348 B.n134 B.n47 10.6151
R349 B.n135 B.n134 10.6151
R350 B.n136 B.n135 10.6151
R351 B.n93 B.n92 10.6151
R352 B.n92 B.n65 10.6151
R353 B.n88 B.n65 10.6151
R354 B.n88 B.n87 10.6151
R355 B.n87 B.n86 10.6151
R356 B.n86 B.n67 10.6151
R357 B.n82 B.n67 10.6151
R358 B.n82 B.n81 10.6151
R359 B.n81 B.n80 10.6151
R360 B.n80 B.n69 10.6151
R361 B.n76 B.n69 10.6151
R362 B.n76 B.n75 10.6151
R363 B.n75 B.n74 10.6151
R364 B.n74 B.n71 10.6151
R365 B.n71 B.n0 10.6151
R366 B.n251 B.n1 10.6151
R367 B.n251 B.n250 10.6151
R368 B.n250 B.n249 10.6151
R369 B.n249 B.n4 10.6151
R370 B.n245 B.n4 10.6151
R371 B.n245 B.n244 10.6151
R372 B.n244 B.n243 10.6151
R373 B.n243 B.n6 10.6151
R374 B.n239 B.n6 10.6151
R375 B.n239 B.n238 10.6151
R376 B.n238 B.n237 10.6151
R377 B.n237 B.n8 10.6151
R378 B.n233 B.n8 10.6151
R379 B.n233 B.n232 10.6151
R380 B.n232 B.n231 10.6151
R381 B.n18 B.n14 8.74196
R382 B.n201 B.n200 8.74196
R383 B.n106 B.n59 8.74196
R384 B.n124 B.n123 8.74196
R385 B.n255 B.n0 2.81026
R386 B.n255 B.n1 2.81026
R387 B.n215 B.n18 1.87367
R388 B.n202 B.n201 1.87367
R389 B.n109 B.n59 1.87367
R390 B.n123 B.n122 1.87367
R391 VN VN.t1 254.827
R392 VN VN.t0 222.297
R393 VTAIL.n2 VTAIL.t3 655.96
R394 VTAIL.n1 VTAIL.t2 655.96
R395 VTAIL.n3 VTAIL.t1 655.958
R396 VTAIL.n0 VTAIL.t0 655.958
R397 VTAIL.n1 VTAIL.n0 15.6083
R398 VTAIL.n3 VTAIL.n2 14.4272
R399 VTAIL.n2 VTAIL.n1 1.06084
R400 VTAIL VTAIL.n0 0.823776
R401 VTAIL VTAIL.n3 0.237569
R402 VDD2.n0 VDD2.t1 699.538
R403 VDD2.n0 VDD2.t0 672.638
R404 VDD2 VDD2.n0 0.353948
R405 VP.n0 VP.t0 254.446
R406 VP.n0 VP.t1 222.245
R407 VP VP.n0 0.0516364
R408 VDD1 VDD1.t0 700.357
R409 VDD1 VDD1.t1 672.991
C0 VTAIL VDD2 1.71371f
C1 VTAIL VN 0.583329f
C2 VP VDD2 0.276756f
C3 VP VN 2.68488f
C4 VTAIL w_n1518_n1172# 1.03103f
C5 VDD2 B 0.671029f
C6 VP w_n1518_n1172# 1.86841f
C7 VN B 0.619164f
C8 VDD1 VDD2 0.493777f
C9 VDD1 VN 0.156804f
C10 w_n1518_n1172# B 4.03577f
C11 VDD1 w_n1518_n1172# 0.799368f
C12 VTAIL VP 0.59747f
C13 VDD2 VN 0.412416f
C14 VTAIL B 0.732673f
C15 VTAIL VDD1 1.67132f
C16 VP B 0.924027f
C17 VDD2 w_n1518_n1172# 0.806356f
C18 VN w_n1518_n1172# 1.68616f
C19 VDD1 VP 0.530806f
C20 VDD1 B 0.653739f
C21 VDD2 VSUBS 0.336008f
C22 VDD1 VSUBS 0.502982f
C23 VTAIL VSUBS 0.194008f
C24 VN VSUBS 3.38328f
C25 VP VSUBS 0.708415f
C26 B VSUBS 1.72982f
C27 w_n1518_n1172# VSUBS 22.933899f
C28 VP.t0 VSUBS 0.378465f
C29 VP.t1 VSUBS 0.241074f
C30 VP.n0 VSUBS 2.05752f
C31 VN.t0 VSUBS 0.23604f
C32 VN.t1 VSUBS 0.375364f
C33 B.n0 VSUBS 0.006702f
C34 B.n1 VSUBS 0.006702f
C35 B.n2 VSUBS 0.010598f
C36 B.n3 VSUBS 0.010598f
C37 B.n4 VSUBS 0.010598f
C38 B.n5 VSUBS 0.010598f
C39 B.n6 VSUBS 0.010598f
C40 B.n7 VSUBS 0.010598f
C41 B.n8 VSUBS 0.010598f
C42 B.n9 VSUBS 0.010598f
C43 B.n10 VSUBS 0.02679f
C44 B.n11 VSUBS 0.010598f
C45 B.n12 VSUBS 0.010598f
C46 B.n13 VSUBS 0.010598f
C47 B.n14 VSUBS 0.009663f
C48 B.n15 VSUBS 0.010598f
C49 B.t5 VSUBS 0.029464f
C50 B.t4 VSUBS 0.031211f
C51 B.t3 VSUBS 0.080361f
C52 B.n16 VSUBS 0.066709f
C53 B.n17 VSUBS 0.059399f
C54 B.n18 VSUBS 0.024555f
C55 B.n19 VSUBS 0.010598f
C56 B.n20 VSUBS 0.010598f
C57 B.n21 VSUBS 0.010598f
C58 B.n22 VSUBS 0.010598f
C59 B.t11 VSUBS 0.029464f
C60 B.t10 VSUBS 0.031211f
C61 B.t9 VSUBS 0.080361f
C62 B.n23 VSUBS 0.066709f
C63 B.n24 VSUBS 0.059399f
C64 B.n25 VSUBS 0.010598f
C65 B.n26 VSUBS 0.010598f
C66 B.n27 VSUBS 0.010598f
C67 B.n28 VSUBS 0.010598f
C68 B.n29 VSUBS 0.026733f
C69 B.n30 VSUBS 0.010598f
C70 B.n31 VSUBS 0.010598f
C71 B.n32 VSUBS 0.010598f
C72 B.n33 VSUBS 0.010598f
C73 B.n34 VSUBS 0.010598f
C74 B.n35 VSUBS 0.010598f
C75 B.n36 VSUBS 0.010598f
C76 B.n37 VSUBS 0.010598f
C77 B.n38 VSUBS 0.010598f
C78 B.n39 VSUBS 0.010598f
C79 B.n40 VSUBS 0.010598f
C80 B.n41 VSUBS 0.010598f
C81 B.n42 VSUBS 0.010598f
C82 B.n43 VSUBS 0.010598f
C83 B.n44 VSUBS 0.010598f
C84 B.n45 VSUBS 0.025579f
C85 B.n46 VSUBS 0.010598f
C86 B.n47 VSUBS 0.010598f
C87 B.n48 VSUBS 0.010598f
C88 B.n49 VSUBS 0.010598f
C89 B.n50 VSUBS 0.010598f
C90 B.t7 VSUBS 0.029464f
C91 B.t8 VSUBS 0.031211f
C92 B.t6 VSUBS 0.080361f
C93 B.n51 VSUBS 0.066709f
C94 B.n52 VSUBS 0.059399f
C95 B.n53 VSUBS 0.010598f
C96 B.n54 VSUBS 0.010598f
C97 B.n55 VSUBS 0.010598f
C98 B.n56 VSUBS 0.010598f
C99 B.t1 VSUBS 0.029464f
C100 B.t2 VSUBS 0.031211f
C101 B.t0 VSUBS 0.080361f
C102 B.n57 VSUBS 0.066709f
C103 B.n58 VSUBS 0.059399f
C104 B.n59 VSUBS 0.024555f
C105 B.n60 VSUBS 0.010598f
C106 B.n61 VSUBS 0.010598f
C107 B.n62 VSUBS 0.010598f
C108 B.n63 VSUBS 0.010598f
C109 B.n64 VSUBS 0.025579f
C110 B.n65 VSUBS 0.010598f
C111 B.n66 VSUBS 0.010598f
C112 B.n67 VSUBS 0.010598f
C113 B.n68 VSUBS 0.010598f
C114 B.n69 VSUBS 0.010598f
C115 B.n70 VSUBS 0.010598f
C116 B.n71 VSUBS 0.010598f
C117 B.n72 VSUBS 0.010598f
C118 B.n73 VSUBS 0.010598f
C119 B.n74 VSUBS 0.010598f
C120 B.n75 VSUBS 0.010598f
C121 B.n76 VSUBS 0.010598f
C122 B.n77 VSUBS 0.010598f
C123 B.n78 VSUBS 0.010598f
C124 B.n79 VSUBS 0.010598f
C125 B.n80 VSUBS 0.010598f
C126 B.n81 VSUBS 0.010598f
C127 B.n82 VSUBS 0.010598f
C128 B.n83 VSUBS 0.010598f
C129 B.n84 VSUBS 0.010598f
C130 B.n85 VSUBS 0.010598f
C131 B.n86 VSUBS 0.010598f
C132 B.n87 VSUBS 0.010598f
C133 B.n88 VSUBS 0.010598f
C134 B.n89 VSUBS 0.010598f
C135 B.n90 VSUBS 0.010598f
C136 B.n91 VSUBS 0.010598f
C137 B.n92 VSUBS 0.010598f
C138 B.n93 VSUBS 0.025579f
C139 B.n94 VSUBS 0.02679f
C140 B.n95 VSUBS 0.02679f
C141 B.n96 VSUBS 0.010598f
C142 B.n97 VSUBS 0.010598f
C143 B.n98 VSUBS 0.010598f
C144 B.n99 VSUBS 0.010598f
C145 B.n100 VSUBS 0.010598f
C146 B.n101 VSUBS 0.010598f
C147 B.n102 VSUBS 0.010598f
C148 B.n103 VSUBS 0.010598f
C149 B.n104 VSUBS 0.010598f
C150 B.n105 VSUBS 0.010598f
C151 B.n106 VSUBS 0.009663f
C152 B.n107 VSUBS 0.010598f
C153 B.n108 VSUBS 0.010598f
C154 B.n109 VSUBS 0.006234f
C155 B.n110 VSUBS 0.010598f
C156 B.n111 VSUBS 0.010598f
C157 B.n112 VSUBS 0.010598f
C158 B.n113 VSUBS 0.010598f
C159 B.n114 VSUBS 0.010598f
C160 B.n115 VSUBS 0.010598f
C161 B.n116 VSUBS 0.010598f
C162 B.n117 VSUBS 0.010598f
C163 B.n118 VSUBS 0.010598f
C164 B.n119 VSUBS 0.010598f
C165 B.n120 VSUBS 0.010598f
C166 B.n121 VSUBS 0.010598f
C167 B.n122 VSUBS 0.006234f
C168 B.n123 VSUBS 0.024555f
C169 B.n124 VSUBS 0.009663f
C170 B.n125 VSUBS 0.010598f
C171 B.n126 VSUBS 0.010598f
C172 B.n127 VSUBS 0.010598f
C173 B.n128 VSUBS 0.010598f
C174 B.n129 VSUBS 0.010598f
C175 B.n130 VSUBS 0.010598f
C176 B.n131 VSUBS 0.010598f
C177 B.n132 VSUBS 0.010598f
C178 B.n133 VSUBS 0.010598f
C179 B.n134 VSUBS 0.010598f
C180 B.n135 VSUBS 0.010598f
C181 B.n136 VSUBS 0.02679f
C182 B.n137 VSUBS 0.02679f
C183 B.n138 VSUBS 0.025579f
C184 B.n139 VSUBS 0.010598f
C185 B.n140 VSUBS 0.010598f
C186 B.n141 VSUBS 0.010598f
C187 B.n142 VSUBS 0.010598f
C188 B.n143 VSUBS 0.010598f
C189 B.n144 VSUBS 0.010598f
C190 B.n145 VSUBS 0.010598f
C191 B.n146 VSUBS 0.010598f
C192 B.n147 VSUBS 0.010598f
C193 B.n148 VSUBS 0.010598f
C194 B.n149 VSUBS 0.010598f
C195 B.n150 VSUBS 0.010598f
C196 B.n151 VSUBS 0.010598f
C197 B.n152 VSUBS 0.010598f
C198 B.n153 VSUBS 0.010598f
C199 B.n154 VSUBS 0.010598f
C200 B.n155 VSUBS 0.010598f
C201 B.n156 VSUBS 0.010598f
C202 B.n157 VSUBS 0.010598f
C203 B.n158 VSUBS 0.010598f
C204 B.n159 VSUBS 0.010598f
C205 B.n160 VSUBS 0.010598f
C206 B.n161 VSUBS 0.010598f
C207 B.n162 VSUBS 0.010598f
C208 B.n163 VSUBS 0.010598f
C209 B.n164 VSUBS 0.010598f
C210 B.n165 VSUBS 0.010598f
C211 B.n166 VSUBS 0.010598f
C212 B.n167 VSUBS 0.010598f
C213 B.n168 VSUBS 0.010598f
C214 B.n169 VSUBS 0.010598f
C215 B.n170 VSUBS 0.010598f
C216 B.n171 VSUBS 0.010598f
C217 B.n172 VSUBS 0.010598f
C218 B.n173 VSUBS 0.010598f
C219 B.n174 VSUBS 0.010598f
C220 B.n175 VSUBS 0.010598f
C221 B.n176 VSUBS 0.010598f
C222 B.n177 VSUBS 0.010598f
C223 B.n178 VSUBS 0.010598f
C224 B.n179 VSUBS 0.010598f
C225 B.n180 VSUBS 0.010598f
C226 B.n181 VSUBS 0.010598f
C227 B.n182 VSUBS 0.010598f
C228 B.n183 VSUBS 0.010598f
C229 B.n184 VSUBS 0.010598f
C230 B.n185 VSUBS 0.010598f
C231 B.n186 VSUBS 0.025579f
C232 B.n187 VSUBS 0.02679f
C233 B.n188 VSUBS 0.025635f
C234 B.n189 VSUBS 0.010598f
C235 B.n190 VSUBS 0.010598f
C236 B.n191 VSUBS 0.010598f
C237 B.n192 VSUBS 0.010598f
C238 B.n193 VSUBS 0.010598f
C239 B.n194 VSUBS 0.010598f
C240 B.n195 VSUBS 0.010598f
C241 B.n196 VSUBS 0.010598f
C242 B.n197 VSUBS 0.010598f
C243 B.n198 VSUBS 0.010598f
C244 B.n199 VSUBS 0.010598f
C245 B.n200 VSUBS 0.009663f
C246 B.n201 VSUBS 0.024555f
C247 B.n202 VSUBS 0.006234f
C248 B.n203 VSUBS 0.010598f
C249 B.n204 VSUBS 0.010598f
C250 B.n205 VSUBS 0.010598f
C251 B.n206 VSUBS 0.010598f
C252 B.n207 VSUBS 0.010598f
C253 B.n208 VSUBS 0.010598f
C254 B.n209 VSUBS 0.010598f
C255 B.n210 VSUBS 0.010598f
C256 B.n211 VSUBS 0.010598f
C257 B.n212 VSUBS 0.010598f
C258 B.n213 VSUBS 0.010598f
C259 B.n214 VSUBS 0.010598f
C260 B.n215 VSUBS 0.006234f
C261 B.n216 VSUBS 0.010598f
C262 B.n217 VSUBS 0.010598f
C263 B.n218 VSUBS 0.010598f
C264 B.n219 VSUBS 0.010598f
C265 B.n220 VSUBS 0.010598f
C266 B.n221 VSUBS 0.010598f
C267 B.n222 VSUBS 0.010598f
C268 B.n223 VSUBS 0.010598f
C269 B.n224 VSUBS 0.010598f
C270 B.n225 VSUBS 0.010598f
C271 B.n226 VSUBS 0.010598f
C272 B.n227 VSUBS 0.010598f
C273 B.n228 VSUBS 0.010598f
C274 B.n229 VSUBS 0.02679f
C275 B.n230 VSUBS 0.025579f
C276 B.n231 VSUBS 0.025579f
C277 B.n232 VSUBS 0.010598f
C278 B.n233 VSUBS 0.010598f
C279 B.n234 VSUBS 0.010598f
C280 B.n235 VSUBS 0.010598f
C281 B.n236 VSUBS 0.010598f
C282 B.n237 VSUBS 0.010598f
C283 B.n238 VSUBS 0.010598f
C284 B.n239 VSUBS 0.010598f
C285 B.n240 VSUBS 0.010598f
C286 B.n241 VSUBS 0.010598f
C287 B.n242 VSUBS 0.010598f
C288 B.n243 VSUBS 0.010598f
C289 B.n244 VSUBS 0.010598f
C290 B.n245 VSUBS 0.010598f
C291 B.n246 VSUBS 0.010598f
C292 B.n247 VSUBS 0.010598f
C293 B.n248 VSUBS 0.010598f
C294 B.n249 VSUBS 0.010598f
C295 B.n250 VSUBS 0.010598f
C296 B.n251 VSUBS 0.010598f
C297 B.n252 VSUBS 0.010598f
C298 B.n253 VSUBS 0.010598f
C299 B.n254 VSUBS 0.010598f
C300 B.n255 VSUBS 0.023999f
.ends

