* NGSPICE file created from diff_pair_sample_0497.ext - technology: sky130A

.subckt diff_pair_sample_0497 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=0.19
X1 VTAIL.t5 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X2 VDD1.t4 VP.t1 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=0.19
X3 VTAIL.t13 VP.t2 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=0.19
X4 VTAIL.t6 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=0.19
X5 VDD1.t0 VP.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X6 VDD1.t3 VP.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=0.19
X7 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X8 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X9 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=0.19
X10 VDD1.t2 VP.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X11 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=0.19
X12 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=0.19
X13 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=0.19
X14 VDD2.t2 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X15 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=2.94525 ps=18.18 w=17.85 l=0.19
X16 VTAIL.t9 VP.t6 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.9615 pd=36.48 as=0 ps=0 w=17.85 l=0.19
X18 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=6.9615 ps=36.48 w=17.85 l=0.19
X19 VTAIL.t8 VP.t7 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.94525 pd=18.18 as=2.94525 ps=18.18 w=17.85 l=0.19
R0 VP.n13 VP.t1 2471.19
R1 VP.n9 VP.t0 2471.19
R2 VP.n2 VP.t2 2471.19
R3 VP.n6 VP.t4 2471.19
R4 VP.n12 VP.t6 2430.29
R5 VP.n10 VP.t3 2430.29
R6 VP.n3 VP.t5 2430.29
R7 VP.n5 VP.t7 2430.29
R8 VP.n2 VP.n1 161.489
R9 VP.n14 VP.n13 161.3
R10 VP.n4 VP.n1 161.3
R11 VP.n7 VP.n6 161.3
R12 VP.n11 VP.n0 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n8 VP.n7 44.0914
R15 VP.n11 VP.n10 37.9763
R16 VP.n12 VP.n11 37.9763
R17 VP.n4 VP.n3 37.9763
R18 VP.n5 VP.n4 37.9763
R19 VP.n10 VP.n9 35.055
R20 VP.n13 VP.n12 35.055
R21 VP.n3 VP.n2 35.055
R22 VP.n6 VP.n5 35.055
R23 VP.n7 VP.n1 0.189894
R24 VP.n8 VP.n0 0.189894
R25 VP.n14 VP.n0 0.189894
R26 VP VP.n14 0.0516364
R27 VDD1 VDD1.n0 60.3645
R28 VDD1.n3 VDD1.n2 60.2507
R29 VDD1.n3 VDD1.n1 60.2507
R30 VDD1.n5 VDD1.n4 60.082
R31 VDD1.n5 VDD1.n3 41.7035
R32 VDD1.n4 VDD1.t6 1.10974
R33 VDD1.n4 VDD1.t3 1.10974
R34 VDD1.n0 VDD1.t1 1.10974
R35 VDD1.n0 VDD1.t2 1.10974
R36 VDD1.n2 VDD1.t7 1.10974
R37 VDD1.n2 VDD1.t4 1.10974
R38 VDD1.n1 VDD1.t5 1.10974
R39 VDD1.n1 VDD1.t0 1.10974
R40 VDD1 VDD1.n5 0.166448
R41 VTAIL.n11 VTAIL.t13 44.5126
R42 VTAIL.n10 VTAIL.t0 44.5126
R43 VTAIL.n7 VTAIL.t2 44.5126
R44 VTAIL.n15 VTAIL.t4 44.5124
R45 VTAIL.n2 VTAIL.t6 44.5124
R46 VTAIL.n3 VTAIL.t14 44.5124
R47 VTAIL.n6 VTAIL.t15 44.5124
R48 VTAIL.n14 VTAIL.t11 44.5124
R49 VTAIL.n13 VTAIL.n12 43.4034
R50 VTAIL.n9 VTAIL.n8 43.4034
R51 VTAIL.n1 VTAIL.n0 43.4032
R52 VTAIL.n5 VTAIL.n4 43.4032
R53 VTAIL.n15 VTAIL.n14 28.2031
R54 VTAIL.n7 VTAIL.n6 28.2031
R55 VTAIL.n0 VTAIL.t3 1.10974
R56 VTAIL.n0 VTAIL.t1 1.10974
R57 VTAIL.n4 VTAIL.t12 1.10974
R58 VTAIL.n4 VTAIL.t9 1.10974
R59 VTAIL.n12 VTAIL.t10 1.10974
R60 VTAIL.n12 VTAIL.t8 1.10974
R61 VTAIL.n8 VTAIL.t7 1.10974
R62 VTAIL.n8 VTAIL.t5 1.10974
R63 VTAIL.n11 VTAIL.n10 0.470328
R64 VTAIL.n3 VTAIL.n2 0.470328
R65 VTAIL.n9 VTAIL.n7 0.448776
R66 VTAIL.n10 VTAIL.n9 0.448776
R67 VTAIL.n13 VTAIL.n11 0.448776
R68 VTAIL.n14 VTAIL.n13 0.448776
R69 VTAIL.n6 VTAIL.n5 0.448776
R70 VTAIL.n5 VTAIL.n3 0.448776
R71 VTAIL.n2 VTAIL.n1 0.448776
R72 VTAIL VTAIL.n15 0.390586
R73 VTAIL VTAIL.n1 0.0586897
R74 B.n101 B.t19 2503.65
R75 B.n98 B.t8 2503.65
R76 B.n450 B.t16 2503.65
R77 B.n447 B.t12 2503.65
R78 B.n772 B.n771 585
R79 B.n773 B.n772 585
R80 B.n354 B.n97 585
R81 B.n353 B.n352 585
R82 B.n351 B.n350 585
R83 B.n349 B.n348 585
R84 B.n347 B.n346 585
R85 B.n345 B.n344 585
R86 B.n343 B.n342 585
R87 B.n341 B.n340 585
R88 B.n339 B.n338 585
R89 B.n337 B.n336 585
R90 B.n335 B.n334 585
R91 B.n333 B.n332 585
R92 B.n331 B.n330 585
R93 B.n329 B.n328 585
R94 B.n327 B.n326 585
R95 B.n325 B.n324 585
R96 B.n323 B.n322 585
R97 B.n321 B.n320 585
R98 B.n319 B.n318 585
R99 B.n317 B.n316 585
R100 B.n315 B.n314 585
R101 B.n313 B.n312 585
R102 B.n311 B.n310 585
R103 B.n309 B.n308 585
R104 B.n307 B.n306 585
R105 B.n305 B.n304 585
R106 B.n303 B.n302 585
R107 B.n301 B.n300 585
R108 B.n299 B.n298 585
R109 B.n297 B.n296 585
R110 B.n295 B.n294 585
R111 B.n293 B.n292 585
R112 B.n291 B.n290 585
R113 B.n289 B.n288 585
R114 B.n287 B.n286 585
R115 B.n285 B.n284 585
R116 B.n283 B.n282 585
R117 B.n281 B.n280 585
R118 B.n279 B.n278 585
R119 B.n277 B.n276 585
R120 B.n275 B.n274 585
R121 B.n273 B.n272 585
R122 B.n271 B.n270 585
R123 B.n269 B.n268 585
R124 B.n267 B.n266 585
R125 B.n265 B.n264 585
R126 B.n263 B.n262 585
R127 B.n261 B.n260 585
R128 B.n259 B.n258 585
R129 B.n257 B.n256 585
R130 B.n255 B.n254 585
R131 B.n253 B.n252 585
R132 B.n251 B.n250 585
R133 B.n249 B.n248 585
R134 B.n247 B.n246 585
R135 B.n245 B.n244 585
R136 B.n243 B.n242 585
R137 B.n241 B.n240 585
R138 B.n239 B.n238 585
R139 B.n237 B.n236 585
R140 B.n235 B.n234 585
R141 B.n233 B.n232 585
R142 B.n231 B.n230 585
R143 B.n229 B.n228 585
R144 B.n227 B.n226 585
R145 B.n225 B.n224 585
R146 B.n223 B.n222 585
R147 B.n220 B.n219 585
R148 B.n218 B.n217 585
R149 B.n216 B.n215 585
R150 B.n214 B.n213 585
R151 B.n212 B.n211 585
R152 B.n210 B.n209 585
R153 B.n208 B.n207 585
R154 B.n206 B.n205 585
R155 B.n204 B.n203 585
R156 B.n202 B.n201 585
R157 B.n200 B.n199 585
R158 B.n198 B.n197 585
R159 B.n196 B.n195 585
R160 B.n194 B.n193 585
R161 B.n192 B.n191 585
R162 B.n190 B.n189 585
R163 B.n188 B.n187 585
R164 B.n186 B.n185 585
R165 B.n184 B.n183 585
R166 B.n182 B.n181 585
R167 B.n180 B.n179 585
R168 B.n178 B.n177 585
R169 B.n176 B.n175 585
R170 B.n174 B.n173 585
R171 B.n172 B.n171 585
R172 B.n170 B.n169 585
R173 B.n168 B.n167 585
R174 B.n166 B.n165 585
R175 B.n164 B.n163 585
R176 B.n162 B.n161 585
R177 B.n160 B.n159 585
R178 B.n158 B.n157 585
R179 B.n156 B.n155 585
R180 B.n154 B.n153 585
R181 B.n152 B.n151 585
R182 B.n150 B.n149 585
R183 B.n148 B.n147 585
R184 B.n146 B.n145 585
R185 B.n144 B.n143 585
R186 B.n142 B.n141 585
R187 B.n140 B.n139 585
R188 B.n138 B.n137 585
R189 B.n136 B.n135 585
R190 B.n134 B.n133 585
R191 B.n132 B.n131 585
R192 B.n130 B.n129 585
R193 B.n128 B.n127 585
R194 B.n126 B.n125 585
R195 B.n124 B.n123 585
R196 B.n122 B.n121 585
R197 B.n120 B.n119 585
R198 B.n118 B.n117 585
R199 B.n116 B.n115 585
R200 B.n114 B.n113 585
R201 B.n112 B.n111 585
R202 B.n110 B.n109 585
R203 B.n108 B.n107 585
R204 B.n106 B.n105 585
R205 B.n104 B.n103 585
R206 B.n770 B.n33 585
R207 B.n774 B.n33 585
R208 B.n769 B.n32 585
R209 B.n775 B.n32 585
R210 B.n768 B.n767 585
R211 B.n767 B.n28 585
R212 B.n766 B.n27 585
R213 B.n781 B.n27 585
R214 B.n765 B.n26 585
R215 B.n782 B.n26 585
R216 B.n764 B.n25 585
R217 B.n783 B.n25 585
R218 B.n763 B.n762 585
R219 B.n762 B.n21 585
R220 B.n761 B.n20 585
R221 B.n789 B.n20 585
R222 B.n760 B.n19 585
R223 B.n790 B.n19 585
R224 B.n759 B.n18 585
R225 B.n791 B.n18 585
R226 B.n758 B.n757 585
R227 B.n757 B.n17 585
R228 B.n756 B.n12 585
R229 B.n797 B.n12 585
R230 B.n755 B.n11 585
R231 B.n798 B.n11 585
R232 B.n754 B.n10 585
R233 B.n799 B.n10 585
R234 B.n753 B.n7 585
R235 B.n802 B.n7 585
R236 B.n752 B.n6 585
R237 B.n803 B.n6 585
R238 B.n751 B.n5 585
R239 B.n804 B.n5 585
R240 B.n750 B.n749 585
R241 B.n749 B.n4 585
R242 B.n748 B.n355 585
R243 B.n748 B.n747 585
R244 B.n738 B.n356 585
R245 B.n357 B.n356 585
R246 B.n740 B.n739 585
R247 B.n741 B.n740 585
R248 B.n737 B.n361 585
R249 B.n364 B.n361 585
R250 B.n736 B.n735 585
R251 B.n735 B.n734 585
R252 B.n363 B.n362 585
R253 B.n727 B.n363 585
R254 B.n726 B.n725 585
R255 B.n728 B.n726 585
R256 B.n724 B.n369 585
R257 B.n369 B.n368 585
R258 B.n723 B.n722 585
R259 B.n722 B.n721 585
R260 B.n371 B.n370 585
R261 B.n372 B.n371 585
R262 B.n714 B.n713 585
R263 B.n715 B.n714 585
R264 B.n712 B.n377 585
R265 B.n377 B.n376 585
R266 B.n711 B.n710 585
R267 B.n710 B.n709 585
R268 B.n379 B.n378 585
R269 B.n380 B.n379 585
R270 B.n705 B.n704 585
R271 B.n383 B.n382 585
R272 B.n701 B.n700 585
R273 B.n702 B.n701 585
R274 B.n699 B.n446 585
R275 B.n698 B.n697 585
R276 B.n696 B.n695 585
R277 B.n694 B.n693 585
R278 B.n692 B.n691 585
R279 B.n690 B.n689 585
R280 B.n688 B.n687 585
R281 B.n686 B.n685 585
R282 B.n684 B.n683 585
R283 B.n682 B.n681 585
R284 B.n680 B.n679 585
R285 B.n678 B.n677 585
R286 B.n676 B.n675 585
R287 B.n674 B.n673 585
R288 B.n672 B.n671 585
R289 B.n670 B.n669 585
R290 B.n668 B.n667 585
R291 B.n666 B.n665 585
R292 B.n664 B.n663 585
R293 B.n662 B.n661 585
R294 B.n660 B.n659 585
R295 B.n658 B.n657 585
R296 B.n656 B.n655 585
R297 B.n654 B.n653 585
R298 B.n652 B.n651 585
R299 B.n650 B.n649 585
R300 B.n648 B.n647 585
R301 B.n646 B.n645 585
R302 B.n644 B.n643 585
R303 B.n642 B.n641 585
R304 B.n640 B.n639 585
R305 B.n638 B.n637 585
R306 B.n636 B.n635 585
R307 B.n634 B.n633 585
R308 B.n632 B.n631 585
R309 B.n630 B.n629 585
R310 B.n628 B.n627 585
R311 B.n626 B.n625 585
R312 B.n624 B.n623 585
R313 B.n622 B.n621 585
R314 B.n620 B.n619 585
R315 B.n618 B.n617 585
R316 B.n616 B.n615 585
R317 B.n614 B.n613 585
R318 B.n612 B.n611 585
R319 B.n610 B.n609 585
R320 B.n608 B.n607 585
R321 B.n606 B.n605 585
R322 B.n604 B.n603 585
R323 B.n602 B.n601 585
R324 B.n600 B.n599 585
R325 B.n598 B.n597 585
R326 B.n596 B.n595 585
R327 B.n594 B.n593 585
R328 B.n592 B.n591 585
R329 B.n590 B.n589 585
R330 B.n588 B.n587 585
R331 B.n586 B.n585 585
R332 B.n584 B.n583 585
R333 B.n582 B.n581 585
R334 B.n580 B.n579 585
R335 B.n578 B.n577 585
R336 B.n576 B.n575 585
R337 B.n574 B.n573 585
R338 B.n572 B.n571 585
R339 B.n569 B.n568 585
R340 B.n567 B.n566 585
R341 B.n565 B.n564 585
R342 B.n563 B.n562 585
R343 B.n561 B.n560 585
R344 B.n559 B.n558 585
R345 B.n557 B.n556 585
R346 B.n555 B.n554 585
R347 B.n553 B.n552 585
R348 B.n551 B.n550 585
R349 B.n549 B.n548 585
R350 B.n547 B.n546 585
R351 B.n545 B.n544 585
R352 B.n543 B.n542 585
R353 B.n541 B.n540 585
R354 B.n539 B.n538 585
R355 B.n537 B.n536 585
R356 B.n535 B.n534 585
R357 B.n533 B.n532 585
R358 B.n531 B.n530 585
R359 B.n529 B.n528 585
R360 B.n527 B.n526 585
R361 B.n525 B.n524 585
R362 B.n523 B.n522 585
R363 B.n521 B.n520 585
R364 B.n519 B.n518 585
R365 B.n517 B.n516 585
R366 B.n515 B.n514 585
R367 B.n513 B.n512 585
R368 B.n511 B.n510 585
R369 B.n509 B.n508 585
R370 B.n507 B.n506 585
R371 B.n505 B.n504 585
R372 B.n503 B.n502 585
R373 B.n501 B.n500 585
R374 B.n499 B.n498 585
R375 B.n497 B.n496 585
R376 B.n495 B.n494 585
R377 B.n493 B.n492 585
R378 B.n491 B.n490 585
R379 B.n489 B.n488 585
R380 B.n487 B.n486 585
R381 B.n485 B.n484 585
R382 B.n483 B.n482 585
R383 B.n481 B.n480 585
R384 B.n479 B.n478 585
R385 B.n477 B.n476 585
R386 B.n475 B.n474 585
R387 B.n473 B.n472 585
R388 B.n471 B.n470 585
R389 B.n469 B.n468 585
R390 B.n467 B.n466 585
R391 B.n465 B.n464 585
R392 B.n463 B.n462 585
R393 B.n461 B.n460 585
R394 B.n459 B.n458 585
R395 B.n457 B.n456 585
R396 B.n455 B.n454 585
R397 B.n453 B.n452 585
R398 B.n706 B.n381 585
R399 B.n381 B.n380 585
R400 B.n708 B.n707 585
R401 B.n709 B.n708 585
R402 B.n375 B.n374 585
R403 B.n376 B.n375 585
R404 B.n717 B.n716 585
R405 B.n716 B.n715 585
R406 B.n718 B.n373 585
R407 B.n373 B.n372 585
R408 B.n720 B.n719 585
R409 B.n721 B.n720 585
R410 B.n367 B.n366 585
R411 B.n368 B.n367 585
R412 B.n730 B.n729 585
R413 B.n729 B.n728 585
R414 B.n731 B.n365 585
R415 B.n727 B.n365 585
R416 B.n733 B.n732 585
R417 B.n734 B.n733 585
R418 B.n360 B.n359 585
R419 B.n364 B.n360 585
R420 B.n743 B.n742 585
R421 B.n742 B.n741 585
R422 B.n744 B.n358 585
R423 B.n358 B.n357 585
R424 B.n746 B.n745 585
R425 B.n747 B.n746 585
R426 B.n3 B.n0 585
R427 B.n4 B.n3 585
R428 B.n801 B.n1 585
R429 B.n802 B.n801 585
R430 B.n800 B.n9 585
R431 B.n800 B.n799 585
R432 B.n14 B.n8 585
R433 B.n798 B.n8 585
R434 B.n796 B.n795 585
R435 B.n797 B.n796 585
R436 B.n794 B.n13 585
R437 B.n17 B.n13 585
R438 B.n793 B.n792 585
R439 B.n792 B.n791 585
R440 B.n16 B.n15 585
R441 B.n790 B.n16 585
R442 B.n788 B.n787 585
R443 B.n789 B.n788 585
R444 B.n786 B.n22 585
R445 B.n22 B.n21 585
R446 B.n785 B.n784 585
R447 B.n784 B.n783 585
R448 B.n24 B.n23 585
R449 B.n782 B.n24 585
R450 B.n780 B.n779 585
R451 B.n781 B.n780 585
R452 B.n778 B.n29 585
R453 B.n29 B.n28 585
R454 B.n777 B.n776 585
R455 B.n776 B.n775 585
R456 B.n31 B.n30 585
R457 B.n774 B.n31 585
R458 B.n805 B.n804 585
R459 B.n803 B.n2 585
R460 B.n103 B.n31 559.769
R461 B.n772 B.n33 559.769
R462 B.n452 B.n379 559.769
R463 B.n704 B.n381 559.769
R464 B.n773 B.n96 256.663
R465 B.n773 B.n95 256.663
R466 B.n773 B.n94 256.663
R467 B.n773 B.n93 256.663
R468 B.n773 B.n92 256.663
R469 B.n773 B.n91 256.663
R470 B.n773 B.n90 256.663
R471 B.n773 B.n89 256.663
R472 B.n773 B.n88 256.663
R473 B.n773 B.n87 256.663
R474 B.n773 B.n86 256.663
R475 B.n773 B.n85 256.663
R476 B.n773 B.n84 256.663
R477 B.n773 B.n83 256.663
R478 B.n773 B.n82 256.663
R479 B.n773 B.n81 256.663
R480 B.n773 B.n80 256.663
R481 B.n773 B.n79 256.663
R482 B.n773 B.n78 256.663
R483 B.n773 B.n77 256.663
R484 B.n773 B.n76 256.663
R485 B.n773 B.n75 256.663
R486 B.n773 B.n74 256.663
R487 B.n773 B.n73 256.663
R488 B.n773 B.n72 256.663
R489 B.n773 B.n71 256.663
R490 B.n773 B.n70 256.663
R491 B.n773 B.n69 256.663
R492 B.n773 B.n68 256.663
R493 B.n773 B.n67 256.663
R494 B.n773 B.n66 256.663
R495 B.n773 B.n65 256.663
R496 B.n773 B.n64 256.663
R497 B.n773 B.n63 256.663
R498 B.n773 B.n62 256.663
R499 B.n773 B.n61 256.663
R500 B.n773 B.n60 256.663
R501 B.n773 B.n59 256.663
R502 B.n773 B.n58 256.663
R503 B.n773 B.n57 256.663
R504 B.n773 B.n56 256.663
R505 B.n773 B.n55 256.663
R506 B.n773 B.n54 256.663
R507 B.n773 B.n53 256.663
R508 B.n773 B.n52 256.663
R509 B.n773 B.n51 256.663
R510 B.n773 B.n50 256.663
R511 B.n773 B.n49 256.663
R512 B.n773 B.n48 256.663
R513 B.n773 B.n47 256.663
R514 B.n773 B.n46 256.663
R515 B.n773 B.n45 256.663
R516 B.n773 B.n44 256.663
R517 B.n773 B.n43 256.663
R518 B.n773 B.n42 256.663
R519 B.n773 B.n41 256.663
R520 B.n773 B.n40 256.663
R521 B.n773 B.n39 256.663
R522 B.n773 B.n38 256.663
R523 B.n773 B.n37 256.663
R524 B.n773 B.n36 256.663
R525 B.n773 B.n35 256.663
R526 B.n773 B.n34 256.663
R527 B.n703 B.n702 256.663
R528 B.n702 B.n384 256.663
R529 B.n702 B.n385 256.663
R530 B.n702 B.n386 256.663
R531 B.n702 B.n387 256.663
R532 B.n702 B.n388 256.663
R533 B.n702 B.n389 256.663
R534 B.n702 B.n390 256.663
R535 B.n702 B.n391 256.663
R536 B.n702 B.n392 256.663
R537 B.n702 B.n393 256.663
R538 B.n702 B.n394 256.663
R539 B.n702 B.n395 256.663
R540 B.n702 B.n396 256.663
R541 B.n702 B.n397 256.663
R542 B.n702 B.n398 256.663
R543 B.n702 B.n399 256.663
R544 B.n702 B.n400 256.663
R545 B.n702 B.n401 256.663
R546 B.n702 B.n402 256.663
R547 B.n702 B.n403 256.663
R548 B.n702 B.n404 256.663
R549 B.n702 B.n405 256.663
R550 B.n702 B.n406 256.663
R551 B.n702 B.n407 256.663
R552 B.n702 B.n408 256.663
R553 B.n702 B.n409 256.663
R554 B.n702 B.n410 256.663
R555 B.n702 B.n411 256.663
R556 B.n702 B.n412 256.663
R557 B.n702 B.n413 256.663
R558 B.n702 B.n414 256.663
R559 B.n702 B.n415 256.663
R560 B.n702 B.n416 256.663
R561 B.n702 B.n417 256.663
R562 B.n702 B.n418 256.663
R563 B.n702 B.n419 256.663
R564 B.n702 B.n420 256.663
R565 B.n702 B.n421 256.663
R566 B.n702 B.n422 256.663
R567 B.n702 B.n423 256.663
R568 B.n702 B.n424 256.663
R569 B.n702 B.n425 256.663
R570 B.n702 B.n426 256.663
R571 B.n702 B.n427 256.663
R572 B.n702 B.n428 256.663
R573 B.n702 B.n429 256.663
R574 B.n702 B.n430 256.663
R575 B.n702 B.n431 256.663
R576 B.n702 B.n432 256.663
R577 B.n702 B.n433 256.663
R578 B.n702 B.n434 256.663
R579 B.n702 B.n435 256.663
R580 B.n702 B.n436 256.663
R581 B.n702 B.n437 256.663
R582 B.n702 B.n438 256.663
R583 B.n702 B.n439 256.663
R584 B.n702 B.n440 256.663
R585 B.n702 B.n441 256.663
R586 B.n702 B.n442 256.663
R587 B.n702 B.n443 256.663
R588 B.n702 B.n444 256.663
R589 B.n702 B.n445 256.663
R590 B.n807 B.n806 256.663
R591 B.n107 B.n106 163.367
R592 B.n111 B.n110 163.367
R593 B.n115 B.n114 163.367
R594 B.n119 B.n118 163.367
R595 B.n123 B.n122 163.367
R596 B.n127 B.n126 163.367
R597 B.n131 B.n130 163.367
R598 B.n135 B.n134 163.367
R599 B.n139 B.n138 163.367
R600 B.n143 B.n142 163.367
R601 B.n147 B.n146 163.367
R602 B.n151 B.n150 163.367
R603 B.n155 B.n154 163.367
R604 B.n159 B.n158 163.367
R605 B.n163 B.n162 163.367
R606 B.n167 B.n166 163.367
R607 B.n171 B.n170 163.367
R608 B.n175 B.n174 163.367
R609 B.n179 B.n178 163.367
R610 B.n183 B.n182 163.367
R611 B.n187 B.n186 163.367
R612 B.n191 B.n190 163.367
R613 B.n195 B.n194 163.367
R614 B.n199 B.n198 163.367
R615 B.n203 B.n202 163.367
R616 B.n207 B.n206 163.367
R617 B.n211 B.n210 163.367
R618 B.n215 B.n214 163.367
R619 B.n219 B.n218 163.367
R620 B.n224 B.n223 163.367
R621 B.n228 B.n227 163.367
R622 B.n232 B.n231 163.367
R623 B.n236 B.n235 163.367
R624 B.n240 B.n239 163.367
R625 B.n244 B.n243 163.367
R626 B.n248 B.n247 163.367
R627 B.n252 B.n251 163.367
R628 B.n256 B.n255 163.367
R629 B.n260 B.n259 163.367
R630 B.n264 B.n263 163.367
R631 B.n268 B.n267 163.367
R632 B.n272 B.n271 163.367
R633 B.n276 B.n275 163.367
R634 B.n280 B.n279 163.367
R635 B.n284 B.n283 163.367
R636 B.n288 B.n287 163.367
R637 B.n292 B.n291 163.367
R638 B.n296 B.n295 163.367
R639 B.n300 B.n299 163.367
R640 B.n304 B.n303 163.367
R641 B.n308 B.n307 163.367
R642 B.n312 B.n311 163.367
R643 B.n316 B.n315 163.367
R644 B.n320 B.n319 163.367
R645 B.n324 B.n323 163.367
R646 B.n328 B.n327 163.367
R647 B.n332 B.n331 163.367
R648 B.n336 B.n335 163.367
R649 B.n340 B.n339 163.367
R650 B.n344 B.n343 163.367
R651 B.n348 B.n347 163.367
R652 B.n352 B.n351 163.367
R653 B.n772 B.n97 163.367
R654 B.n710 B.n379 163.367
R655 B.n710 B.n377 163.367
R656 B.n714 B.n377 163.367
R657 B.n714 B.n371 163.367
R658 B.n722 B.n371 163.367
R659 B.n722 B.n369 163.367
R660 B.n726 B.n369 163.367
R661 B.n726 B.n363 163.367
R662 B.n735 B.n363 163.367
R663 B.n735 B.n361 163.367
R664 B.n740 B.n361 163.367
R665 B.n740 B.n356 163.367
R666 B.n748 B.n356 163.367
R667 B.n749 B.n748 163.367
R668 B.n749 B.n5 163.367
R669 B.n6 B.n5 163.367
R670 B.n7 B.n6 163.367
R671 B.n10 B.n7 163.367
R672 B.n11 B.n10 163.367
R673 B.n12 B.n11 163.367
R674 B.n757 B.n12 163.367
R675 B.n757 B.n18 163.367
R676 B.n19 B.n18 163.367
R677 B.n20 B.n19 163.367
R678 B.n762 B.n20 163.367
R679 B.n762 B.n25 163.367
R680 B.n26 B.n25 163.367
R681 B.n27 B.n26 163.367
R682 B.n767 B.n27 163.367
R683 B.n767 B.n32 163.367
R684 B.n33 B.n32 163.367
R685 B.n701 B.n383 163.367
R686 B.n701 B.n446 163.367
R687 B.n697 B.n696 163.367
R688 B.n693 B.n692 163.367
R689 B.n689 B.n688 163.367
R690 B.n685 B.n684 163.367
R691 B.n681 B.n680 163.367
R692 B.n677 B.n676 163.367
R693 B.n673 B.n672 163.367
R694 B.n669 B.n668 163.367
R695 B.n665 B.n664 163.367
R696 B.n661 B.n660 163.367
R697 B.n657 B.n656 163.367
R698 B.n653 B.n652 163.367
R699 B.n649 B.n648 163.367
R700 B.n645 B.n644 163.367
R701 B.n641 B.n640 163.367
R702 B.n637 B.n636 163.367
R703 B.n633 B.n632 163.367
R704 B.n629 B.n628 163.367
R705 B.n625 B.n624 163.367
R706 B.n621 B.n620 163.367
R707 B.n617 B.n616 163.367
R708 B.n613 B.n612 163.367
R709 B.n609 B.n608 163.367
R710 B.n605 B.n604 163.367
R711 B.n601 B.n600 163.367
R712 B.n597 B.n596 163.367
R713 B.n593 B.n592 163.367
R714 B.n589 B.n588 163.367
R715 B.n585 B.n584 163.367
R716 B.n581 B.n580 163.367
R717 B.n577 B.n576 163.367
R718 B.n573 B.n572 163.367
R719 B.n568 B.n567 163.367
R720 B.n564 B.n563 163.367
R721 B.n560 B.n559 163.367
R722 B.n556 B.n555 163.367
R723 B.n552 B.n551 163.367
R724 B.n548 B.n547 163.367
R725 B.n544 B.n543 163.367
R726 B.n540 B.n539 163.367
R727 B.n536 B.n535 163.367
R728 B.n532 B.n531 163.367
R729 B.n528 B.n527 163.367
R730 B.n524 B.n523 163.367
R731 B.n520 B.n519 163.367
R732 B.n516 B.n515 163.367
R733 B.n512 B.n511 163.367
R734 B.n508 B.n507 163.367
R735 B.n504 B.n503 163.367
R736 B.n500 B.n499 163.367
R737 B.n496 B.n495 163.367
R738 B.n492 B.n491 163.367
R739 B.n488 B.n487 163.367
R740 B.n484 B.n483 163.367
R741 B.n480 B.n479 163.367
R742 B.n476 B.n475 163.367
R743 B.n472 B.n471 163.367
R744 B.n468 B.n467 163.367
R745 B.n464 B.n463 163.367
R746 B.n460 B.n459 163.367
R747 B.n456 B.n455 163.367
R748 B.n708 B.n381 163.367
R749 B.n708 B.n375 163.367
R750 B.n716 B.n375 163.367
R751 B.n716 B.n373 163.367
R752 B.n720 B.n373 163.367
R753 B.n720 B.n367 163.367
R754 B.n729 B.n367 163.367
R755 B.n729 B.n365 163.367
R756 B.n733 B.n365 163.367
R757 B.n733 B.n360 163.367
R758 B.n742 B.n360 163.367
R759 B.n742 B.n358 163.367
R760 B.n746 B.n358 163.367
R761 B.n746 B.n3 163.367
R762 B.n805 B.n3 163.367
R763 B.n801 B.n2 163.367
R764 B.n801 B.n800 163.367
R765 B.n800 B.n8 163.367
R766 B.n796 B.n8 163.367
R767 B.n796 B.n13 163.367
R768 B.n792 B.n13 163.367
R769 B.n792 B.n16 163.367
R770 B.n788 B.n16 163.367
R771 B.n788 B.n22 163.367
R772 B.n784 B.n22 163.367
R773 B.n784 B.n24 163.367
R774 B.n780 B.n24 163.367
R775 B.n780 B.n29 163.367
R776 B.n776 B.n29 163.367
R777 B.n776 B.n31 163.367
R778 B.n98 B.t10 80.6394
R779 B.n450 B.t18 80.6394
R780 B.n101 B.t20 80.6157
R781 B.n447 B.t15 80.6157
R782 B.n103 B.n34 71.676
R783 B.n107 B.n35 71.676
R784 B.n111 B.n36 71.676
R785 B.n115 B.n37 71.676
R786 B.n119 B.n38 71.676
R787 B.n123 B.n39 71.676
R788 B.n127 B.n40 71.676
R789 B.n131 B.n41 71.676
R790 B.n135 B.n42 71.676
R791 B.n139 B.n43 71.676
R792 B.n143 B.n44 71.676
R793 B.n147 B.n45 71.676
R794 B.n151 B.n46 71.676
R795 B.n155 B.n47 71.676
R796 B.n159 B.n48 71.676
R797 B.n163 B.n49 71.676
R798 B.n167 B.n50 71.676
R799 B.n171 B.n51 71.676
R800 B.n175 B.n52 71.676
R801 B.n179 B.n53 71.676
R802 B.n183 B.n54 71.676
R803 B.n187 B.n55 71.676
R804 B.n191 B.n56 71.676
R805 B.n195 B.n57 71.676
R806 B.n199 B.n58 71.676
R807 B.n203 B.n59 71.676
R808 B.n207 B.n60 71.676
R809 B.n211 B.n61 71.676
R810 B.n215 B.n62 71.676
R811 B.n219 B.n63 71.676
R812 B.n224 B.n64 71.676
R813 B.n228 B.n65 71.676
R814 B.n232 B.n66 71.676
R815 B.n236 B.n67 71.676
R816 B.n240 B.n68 71.676
R817 B.n244 B.n69 71.676
R818 B.n248 B.n70 71.676
R819 B.n252 B.n71 71.676
R820 B.n256 B.n72 71.676
R821 B.n260 B.n73 71.676
R822 B.n264 B.n74 71.676
R823 B.n268 B.n75 71.676
R824 B.n272 B.n76 71.676
R825 B.n276 B.n77 71.676
R826 B.n280 B.n78 71.676
R827 B.n284 B.n79 71.676
R828 B.n288 B.n80 71.676
R829 B.n292 B.n81 71.676
R830 B.n296 B.n82 71.676
R831 B.n300 B.n83 71.676
R832 B.n304 B.n84 71.676
R833 B.n308 B.n85 71.676
R834 B.n312 B.n86 71.676
R835 B.n316 B.n87 71.676
R836 B.n320 B.n88 71.676
R837 B.n324 B.n89 71.676
R838 B.n328 B.n90 71.676
R839 B.n332 B.n91 71.676
R840 B.n336 B.n92 71.676
R841 B.n340 B.n93 71.676
R842 B.n344 B.n94 71.676
R843 B.n348 B.n95 71.676
R844 B.n352 B.n96 71.676
R845 B.n97 B.n96 71.676
R846 B.n351 B.n95 71.676
R847 B.n347 B.n94 71.676
R848 B.n343 B.n93 71.676
R849 B.n339 B.n92 71.676
R850 B.n335 B.n91 71.676
R851 B.n331 B.n90 71.676
R852 B.n327 B.n89 71.676
R853 B.n323 B.n88 71.676
R854 B.n319 B.n87 71.676
R855 B.n315 B.n86 71.676
R856 B.n311 B.n85 71.676
R857 B.n307 B.n84 71.676
R858 B.n303 B.n83 71.676
R859 B.n299 B.n82 71.676
R860 B.n295 B.n81 71.676
R861 B.n291 B.n80 71.676
R862 B.n287 B.n79 71.676
R863 B.n283 B.n78 71.676
R864 B.n279 B.n77 71.676
R865 B.n275 B.n76 71.676
R866 B.n271 B.n75 71.676
R867 B.n267 B.n74 71.676
R868 B.n263 B.n73 71.676
R869 B.n259 B.n72 71.676
R870 B.n255 B.n71 71.676
R871 B.n251 B.n70 71.676
R872 B.n247 B.n69 71.676
R873 B.n243 B.n68 71.676
R874 B.n239 B.n67 71.676
R875 B.n235 B.n66 71.676
R876 B.n231 B.n65 71.676
R877 B.n227 B.n64 71.676
R878 B.n223 B.n63 71.676
R879 B.n218 B.n62 71.676
R880 B.n214 B.n61 71.676
R881 B.n210 B.n60 71.676
R882 B.n206 B.n59 71.676
R883 B.n202 B.n58 71.676
R884 B.n198 B.n57 71.676
R885 B.n194 B.n56 71.676
R886 B.n190 B.n55 71.676
R887 B.n186 B.n54 71.676
R888 B.n182 B.n53 71.676
R889 B.n178 B.n52 71.676
R890 B.n174 B.n51 71.676
R891 B.n170 B.n50 71.676
R892 B.n166 B.n49 71.676
R893 B.n162 B.n48 71.676
R894 B.n158 B.n47 71.676
R895 B.n154 B.n46 71.676
R896 B.n150 B.n45 71.676
R897 B.n146 B.n44 71.676
R898 B.n142 B.n43 71.676
R899 B.n138 B.n42 71.676
R900 B.n134 B.n41 71.676
R901 B.n130 B.n40 71.676
R902 B.n126 B.n39 71.676
R903 B.n122 B.n38 71.676
R904 B.n118 B.n37 71.676
R905 B.n114 B.n36 71.676
R906 B.n110 B.n35 71.676
R907 B.n106 B.n34 71.676
R908 B.n704 B.n703 71.676
R909 B.n446 B.n384 71.676
R910 B.n696 B.n385 71.676
R911 B.n692 B.n386 71.676
R912 B.n688 B.n387 71.676
R913 B.n684 B.n388 71.676
R914 B.n680 B.n389 71.676
R915 B.n676 B.n390 71.676
R916 B.n672 B.n391 71.676
R917 B.n668 B.n392 71.676
R918 B.n664 B.n393 71.676
R919 B.n660 B.n394 71.676
R920 B.n656 B.n395 71.676
R921 B.n652 B.n396 71.676
R922 B.n648 B.n397 71.676
R923 B.n644 B.n398 71.676
R924 B.n640 B.n399 71.676
R925 B.n636 B.n400 71.676
R926 B.n632 B.n401 71.676
R927 B.n628 B.n402 71.676
R928 B.n624 B.n403 71.676
R929 B.n620 B.n404 71.676
R930 B.n616 B.n405 71.676
R931 B.n612 B.n406 71.676
R932 B.n608 B.n407 71.676
R933 B.n604 B.n408 71.676
R934 B.n600 B.n409 71.676
R935 B.n596 B.n410 71.676
R936 B.n592 B.n411 71.676
R937 B.n588 B.n412 71.676
R938 B.n584 B.n413 71.676
R939 B.n580 B.n414 71.676
R940 B.n576 B.n415 71.676
R941 B.n572 B.n416 71.676
R942 B.n567 B.n417 71.676
R943 B.n563 B.n418 71.676
R944 B.n559 B.n419 71.676
R945 B.n555 B.n420 71.676
R946 B.n551 B.n421 71.676
R947 B.n547 B.n422 71.676
R948 B.n543 B.n423 71.676
R949 B.n539 B.n424 71.676
R950 B.n535 B.n425 71.676
R951 B.n531 B.n426 71.676
R952 B.n527 B.n427 71.676
R953 B.n523 B.n428 71.676
R954 B.n519 B.n429 71.676
R955 B.n515 B.n430 71.676
R956 B.n511 B.n431 71.676
R957 B.n507 B.n432 71.676
R958 B.n503 B.n433 71.676
R959 B.n499 B.n434 71.676
R960 B.n495 B.n435 71.676
R961 B.n491 B.n436 71.676
R962 B.n487 B.n437 71.676
R963 B.n483 B.n438 71.676
R964 B.n479 B.n439 71.676
R965 B.n475 B.n440 71.676
R966 B.n471 B.n441 71.676
R967 B.n467 B.n442 71.676
R968 B.n463 B.n443 71.676
R969 B.n459 B.n444 71.676
R970 B.n455 B.n445 71.676
R971 B.n703 B.n383 71.676
R972 B.n697 B.n384 71.676
R973 B.n693 B.n385 71.676
R974 B.n689 B.n386 71.676
R975 B.n685 B.n387 71.676
R976 B.n681 B.n388 71.676
R977 B.n677 B.n389 71.676
R978 B.n673 B.n390 71.676
R979 B.n669 B.n391 71.676
R980 B.n665 B.n392 71.676
R981 B.n661 B.n393 71.676
R982 B.n657 B.n394 71.676
R983 B.n653 B.n395 71.676
R984 B.n649 B.n396 71.676
R985 B.n645 B.n397 71.676
R986 B.n641 B.n398 71.676
R987 B.n637 B.n399 71.676
R988 B.n633 B.n400 71.676
R989 B.n629 B.n401 71.676
R990 B.n625 B.n402 71.676
R991 B.n621 B.n403 71.676
R992 B.n617 B.n404 71.676
R993 B.n613 B.n405 71.676
R994 B.n609 B.n406 71.676
R995 B.n605 B.n407 71.676
R996 B.n601 B.n408 71.676
R997 B.n597 B.n409 71.676
R998 B.n593 B.n410 71.676
R999 B.n589 B.n411 71.676
R1000 B.n585 B.n412 71.676
R1001 B.n581 B.n413 71.676
R1002 B.n577 B.n414 71.676
R1003 B.n573 B.n415 71.676
R1004 B.n568 B.n416 71.676
R1005 B.n564 B.n417 71.676
R1006 B.n560 B.n418 71.676
R1007 B.n556 B.n419 71.676
R1008 B.n552 B.n420 71.676
R1009 B.n548 B.n421 71.676
R1010 B.n544 B.n422 71.676
R1011 B.n540 B.n423 71.676
R1012 B.n536 B.n424 71.676
R1013 B.n532 B.n425 71.676
R1014 B.n528 B.n426 71.676
R1015 B.n524 B.n427 71.676
R1016 B.n520 B.n428 71.676
R1017 B.n516 B.n429 71.676
R1018 B.n512 B.n430 71.676
R1019 B.n508 B.n431 71.676
R1020 B.n504 B.n432 71.676
R1021 B.n500 B.n433 71.676
R1022 B.n496 B.n434 71.676
R1023 B.n492 B.n435 71.676
R1024 B.n488 B.n436 71.676
R1025 B.n484 B.n437 71.676
R1026 B.n480 B.n438 71.676
R1027 B.n476 B.n439 71.676
R1028 B.n472 B.n440 71.676
R1029 B.n468 B.n441 71.676
R1030 B.n464 B.n442 71.676
R1031 B.n460 B.n443 71.676
R1032 B.n456 B.n444 71.676
R1033 B.n452 B.n445 71.676
R1034 B.n806 B.n805 71.676
R1035 B.n806 B.n2 71.676
R1036 B.n99 B.t11 70.5546
R1037 B.n451 B.t17 70.5546
R1038 B.n102 B.t21 70.5309
R1039 B.n448 B.t14 70.5309
R1040 B.n702 B.n380 67.0708
R1041 B.n774 B.n773 67.0708
R1042 B.n221 B.n102 59.5399
R1043 B.n100 B.n99 59.5399
R1044 B.n570 B.n451 59.5399
R1045 B.n449 B.n448 59.5399
R1046 B.n771 B.n770 36.3712
R1047 B.n706 B.n705 36.3712
R1048 B.n453 B.n378 36.3712
R1049 B.n104 B.n30 36.3712
R1050 B.n709 B.n380 32.3464
R1051 B.n709 B.n376 32.3464
R1052 B.n715 B.n376 32.3464
R1053 B.n721 B.n372 32.3464
R1054 B.n721 B.n368 32.3464
R1055 B.n728 B.n368 32.3464
R1056 B.n728 B.n727 32.3464
R1057 B.n734 B.n364 32.3464
R1058 B.n747 B.n357 32.3464
R1059 B.n804 B.n4 32.3464
R1060 B.n804 B.n803 32.3464
R1061 B.n803 B.n802 32.3464
R1062 B.n799 B.n798 32.3464
R1063 B.n791 B.n17 32.3464
R1064 B.n790 B.n789 32.3464
R1065 B.n789 B.n21 32.3464
R1066 B.n783 B.n21 32.3464
R1067 B.n783 B.n782 32.3464
R1068 B.n781 B.n28 32.3464
R1069 B.n775 B.n28 32.3464
R1070 B.n775 B.n774 32.3464
R1071 B.n741 B.t7 29.9681
R1072 B.n797 B.t1 29.9681
R1073 B.t0 B.n4 28.0654
R1074 B.n802 B.t6 28.0654
R1075 B.n715 B.t13 26.1627
R1076 B.t9 B.n781 26.1627
R1077 B.n741 B.t5 19.5032
R1078 B.t3 B.n797 19.5032
R1079 B B.n807 18.0485
R1080 B.n727 B.t2 17.6005
R1081 B.t4 B.n790 17.6005
R1082 B.n734 B.t2 14.7464
R1083 B.n791 B.t4 14.7464
R1084 B.t5 B.n357 12.8437
R1085 B.n798 B.t3 12.8437
R1086 B.n707 B.n706 10.6151
R1087 B.n707 B.n374 10.6151
R1088 B.n717 B.n374 10.6151
R1089 B.n718 B.n717 10.6151
R1090 B.n719 B.n718 10.6151
R1091 B.n719 B.n366 10.6151
R1092 B.n730 B.n366 10.6151
R1093 B.n731 B.n730 10.6151
R1094 B.n732 B.n731 10.6151
R1095 B.n732 B.n359 10.6151
R1096 B.n743 B.n359 10.6151
R1097 B.n744 B.n743 10.6151
R1098 B.n745 B.n744 10.6151
R1099 B.n745 B.n0 10.6151
R1100 B.n705 B.n382 10.6151
R1101 B.n700 B.n382 10.6151
R1102 B.n700 B.n699 10.6151
R1103 B.n699 B.n698 10.6151
R1104 B.n698 B.n695 10.6151
R1105 B.n695 B.n694 10.6151
R1106 B.n694 B.n691 10.6151
R1107 B.n691 B.n690 10.6151
R1108 B.n690 B.n687 10.6151
R1109 B.n687 B.n686 10.6151
R1110 B.n686 B.n683 10.6151
R1111 B.n683 B.n682 10.6151
R1112 B.n682 B.n679 10.6151
R1113 B.n679 B.n678 10.6151
R1114 B.n678 B.n675 10.6151
R1115 B.n675 B.n674 10.6151
R1116 B.n674 B.n671 10.6151
R1117 B.n671 B.n670 10.6151
R1118 B.n670 B.n667 10.6151
R1119 B.n667 B.n666 10.6151
R1120 B.n666 B.n663 10.6151
R1121 B.n663 B.n662 10.6151
R1122 B.n662 B.n659 10.6151
R1123 B.n659 B.n658 10.6151
R1124 B.n658 B.n655 10.6151
R1125 B.n655 B.n654 10.6151
R1126 B.n654 B.n651 10.6151
R1127 B.n651 B.n650 10.6151
R1128 B.n650 B.n647 10.6151
R1129 B.n647 B.n646 10.6151
R1130 B.n646 B.n643 10.6151
R1131 B.n643 B.n642 10.6151
R1132 B.n642 B.n639 10.6151
R1133 B.n639 B.n638 10.6151
R1134 B.n638 B.n635 10.6151
R1135 B.n635 B.n634 10.6151
R1136 B.n634 B.n631 10.6151
R1137 B.n631 B.n630 10.6151
R1138 B.n630 B.n627 10.6151
R1139 B.n627 B.n626 10.6151
R1140 B.n626 B.n623 10.6151
R1141 B.n623 B.n622 10.6151
R1142 B.n622 B.n619 10.6151
R1143 B.n619 B.n618 10.6151
R1144 B.n618 B.n615 10.6151
R1145 B.n615 B.n614 10.6151
R1146 B.n614 B.n611 10.6151
R1147 B.n611 B.n610 10.6151
R1148 B.n610 B.n607 10.6151
R1149 B.n607 B.n606 10.6151
R1150 B.n606 B.n603 10.6151
R1151 B.n603 B.n602 10.6151
R1152 B.n602 B.n599 10.6151
R1153 B.n599 B.n598 10.6151
R1154 B.n598 B.n595 10.6151
R1155 B.n595 B.n594 10.6151
R1156 B.n594 B.n591 10.6151
R1157 B.n591 B.n590 10.6151
R1158 B.n587 B.n586 10.6151
R1159 B.n586 B.n583 10.6151
R1160 B.n583 B.n582 10.6151
R1161 B.n582 B.n579 10.6151
R1162 B.n579 B.n578 10.6151
R1163 B.n578 B.n575 10.6151
R1164 B.n575 B.n574 10.6151
R1165 B.n574 B.n571 10.6151
R1166 B.n569 B.n566 10.6151
R1167 B.n566 B.n565 10.6151
R1168 B.n565 B.n562 10.6151
R1169 B.n562 B.n561 10.6151
R1170 B.n561 B.n558 10.6151
R1171 B.n558 B.n557 10.6151
R1172 B.n557 B.n554 10.6151
R1173 B.n554 B.n553 10.6151
R1174 B.n553 B.n550 10.6151
R1175 B.n550 B.n549 10.6151
R1176 B.n549 B.n546 10.6151
R1177 B.n546 B.n545 10.6151
R1178 B.n545 B.n542 10.6151
R1179 B.n542 B.n541 10.6151
R1180 B.n541 B.n538 10.6151
R1181 B.n538 B.n537 10.6151
R1182 B.n537 B.n534 10.6151
R1183 B.n534 B.n533 10.6151
R1184 B.n533 B.n530 10.6151
R1185 B.n530 B.n529 10.6151
R1186 B.n529 B.n526 10.6151
R1187 B.n526 B.n525 10.6151
R1188 B.n525 B.n522 10.6151
R1189 B.n522 B.n521 10.6151
R1190 B.n521 B.n518 10.6151
R1191 B.n518 B.n517 10.6151
R1192 B.n517 B.n514 10.6151
R1193 B.n514 B.n513 10.6151
R1194 B.n513 B.n510 10.6151
R1195 B.n510 B.n509 10.6151
R1196 B.n509 B.n506 10.6151
R1197 B.n506 B.n505 10.6151
R1198 B.n505 B.n502 10.6151
R1199 B.n502 B.n501 10.6151
R1200 B.n501 B.n498 10.6151
R1201 B.n498 B.n497 10.6151
R1202 B.n497 B.n494 10.6151
R1203 B.n494 B.n493 10.6151
R1204 B.n493 B.n490 10.6151
R1205 B.n490 B.n489 10.6151
R1206 B.n489 B.n486 10.6151
R1207 B.n486 B.n485 10.6151
R1208 B.n485 B.n482 10.6151
R1209 B.n482 B.n481 10.6151
R1210 B.n481 B.n478 10.6151
R1211 B.n478 B.n477 10.6151
R1212 B.n477 B.n474 10.6151
R1213 B.n474 B.n473 10.6151
R1214 B.n473 B.n470 10.6151
R1215 B.n470 B.n469 10.6151
R1216 B.n469 B.n466 10.6151
R1217 B.n466 B.n465 10.6151
R1218 B.n465 B.n462 10.6151
R1219 B.n462 B.n461 10.6151
R1220 B.n461 B.n458 10.6151
R1221 B.n458 B.n457 10.6151
R1222 B.n457 B.n454 10.6151
R1223 B.n454 B.n453 10.6151
R1224 B.n711 B.n378 10.6151
R1225 B.n712 B.n711 10.6151
R1226 B.n713 B.n712 10.6151
R1227 B.n713 B.n370 10.6151
R1228 B.n723 B.n370 10.6151
R1229 B.n724 B.n723 10.6151
R1230 B.n725 B.n724 10.6151
R1231 B.n725 B.n362 10.6151
R1232 B.n736 B.n362 10.6151
R1233 B.n737 B.n736 10.6151
R1234 B.n739 B.n737 10.6151
R1235 B.n739 B.n738 10.6151
R1236 B.n738 B.n355 10.6151
R1237 B.n750 B.n355 10.6151
R1238 B.n751 B.n750 10.6151
R1239 B.n752 B.n751 10.6151
R1240 B.n753 B.n752 10.6151
R1241 B.n754 B.n753 10.6151
R1242 B.n755 B.n754 10.6151
R1243 B.n756 B.n755 10.6151
R1244 B.n758 B.n756 10.6151
R1245 B.n759 B.n758 10.6151
R1246 B.n760 B.n759 10.6151
R1247 B.n761 B.n760 10.6151
R1248 B.n763 B.n761 10.6151
R1249 B.n764 B.n763 10.6151
R1250 B.n765 B.n764 10.6151
R1251 B.n766 B.n765 10.6151
R1252 B.n768 B.n766 10.6151
R1253 B.n769 B.n768 10.6151
R1254 B.n770 B.n769 10.6151
R1255 B.n9 B.n1 10.6151
R1256 B.n14 B.n9 10.6151
R1257 B.n795 B.n14 10.6151
R1258 B.n795 B.n794 10.6151
R1259 B.n794 B.n793 10.6151
R1260 B.n793 B.n15 10.6151
R1261 B.n787 B.n15 10.6151
R1262 B.n787 B.n786 10.6151
R1263 B.n786 B.n785 10.6151
R1264 B.n785 B.n23 10.6151
R1265 B.n779 B.n23 10.6151
R1266 B.n779 B.n778 10.6151
R1267 B.n778 B.n777 10.6151
R1268 B.n777 B.n30 10.6151
R1269 B.n105 B.n104 10.6151
R1270 B.n108 B.n105 10.6151
R1271 B.n109 B.n108 10.6151
R1272 B.n112 B.n109 10.6151
R1273 B.n113 B.n112 10.6151
R1274 B.n116 B.n113 10.6151
R1275 B.n117 B.n116 10.6151
R1276 B.n120 B.n117 10.6151
R1277 B.n121 B.n120 10.6151
R1278 B.n124 B.n121 10.6151
R1279 B.n125 B.n124 10.6151
R1280 B.n128 B.n125 10.6151
R1281 B.n129 B.n128 10.6151
R1282 B.n132 B.n129 10.6151
R1283 B.n133 B.n132 10.6151
R1284 B.n136 B.n133 10.6151
R1285 B.n137 B.n136 10.6151
R1286 B.n140 B.n137 10.6151
R1287 B.n141 B.n140 10.6151
R1288 B.n144 B.n141 10.6151
R1289 B.n145 B.n144 10.6151
R1290 B.n148 B.n145 10.6151
R1291 B.n149 B.n148 10.6151
R1292 B.n152 B.n149 10.6151
R1293 B.n153 B.n152 10.6151
R1294 B.n156 B.n153 10.6151
R1295 B.n157 B.n156 10.6151
R1296 B.n160 B.n157 10.6151
R1297 B.n161 B.n160 10.6151
R1298 B.n164 B.n161 10.6151
R1299 B.n165 B.n164 10.6151
R1300 B.n168 B.n165 10.6151
R1301 B.n169 B.n168 10.6151
R1302 B.n172 B.n169 10.6151
R1303 B.n173 B.n172 10.6151
R1304 B.n176 B.n173 10.6151
R1305 B.n177 B.n176 10.6151
R1306 B.n180 B.n177 10.6151
R1307 B.n181 B.n180 10.6151
R1308 B.n184 B.n181 10.6151
R1309 B.n185 B.n184 10.6151
R1310 B.n188 B.n185 10.6151
R1311 B.n189 B.n188 10.6151
R1312 B.n192 B.n189 10.6151
R1313 B.n193 B.n192 10.6151
R1314 B.n196 B.n193 10.6151
R1315 B.n197 B.n196 10.6151
R1316 B.n200 B.n197 10.6151
R1317 B.n201 B.n200 10.6151
R1318 B.n204 B.n201 10.6151
R1319 B.n205 B.n204 10.6151
R1320 B.n208 B.n205 10.6151
R1321 B.n209 B.n208 10.6151
R1322 B.n212 B.n209 10.6151
R1323 B.n213 B.n212 10.6151
R1324 B.n216 B.n213 10.6151
R1325 B.n217 B.n216 10.6151
R1326 B.n220 B.n217 10.6151
R1327 B.n225 B.n222 10.6151
R1328 B.n226 B.n225 10.6151
R1329 B.n229 B.n226 10.6151
R1330 B.n230 B.n229 10.6151
R1331 B.n233 B.n230 10.6151
R1332 B.n234 B.n233 10.6151
R1333 B.n237 B.n234 10.6151
R1334 B.n238 B.n237 10.6151
R1335 B.n242 B.n241 10.6151
R1336 B.n245 B.n242 10.6151
R1337 B.n246 B.n245 10.6151
R1338 B.n249 B.n246 10.6151
R1339 B.n250 B.n249 10.6151
R1340 B.n253 B.n250 10.6151
R1341 B.n254 B.n253 10.6151
R1342 B.n257 B.n254 10.6151
R1343 B.n258 B.n257 10.6151
R1344 B.n261 B.n258 10.6151
R1345 B.n262 B.n261 10.6151
R1346 B.n265 B.n262 10.6151
R1347 B.n266 B.n265 10.6151
R1348 B.n269 B.n266 10.6151
R1349 B.n270 B.n269 10.6151
R1350 B.n273 B.n270 10.6151
R1351 B.n274 B.n273 10.6151
R1352 B.n277 B.n274 10.6151
R1353 B.n278 B.n277 10.6151
R1354 B.n281 B.n278 10.6151
R1355 B.n282 B.n281 10.6151
R1356 B.n285 B.n282 10.6151
R1357 B.n286 B.n285 10.6151
R1358 B.n289 B.n286 10.6151
R1359 B.n290 B.n289 10.6151
R1360 B.n293 B.n290 10.6151
R1361 B.n294 B.n293 10.6151
R1362 B.n297 B.n294 10.6151
R1363 B.n298 B.n297 10.6151
R1364 B.n301 B.n298 10.6151
R1365 B.n302 B.n301 10.6151
R1366 B.n305 B.n302 10.6151
R1367 B.n306 B.n305 10.6151
R1368 B.n309 B.n306 10.6151
R1369 B.n310 B.n309 10.6151
R1370 B.n313 B.n310 10.6151
R1371 B.n314 B.n313 10.6151
R1372 B.n317 B.n314 10.6151
R1373 B.n318 B.n317 10.6151
R1374 B.n321 B.n318 10.6151
R1375 B.n322 B.n321 10.6151
R1376 B.n325 B.n322 10.6151
R1377 B.n326 B.n325 10.6151
R1378 B.n329 B.n326 10.6151
R1379 B.n330 B.n329 10.6151
R1380 B.n333 B.n330 10.6151
R1381 B.n334 B.n333 10.6151
R1382 B.n337 B.n334 10.6151
R1383 B.n338 B.n337 10.6151
R1384 B.n341 B.n338 10.6151
R1385 B.n342 B.n341 10.6151
R1386 B.n345 B.n342 10.6151
R1387 B.n346 B.n345 10.6151
R1388 B.n349 B.n346 10.6151
R1389 B.n350 B.n349 10.6151
R1390 B.n353 B.n350 10.6151
R1391 B.n354 B.n353 10.6151
R1392 B.n771 B.n354 10.6151
R1393 B.n102 B.n101 10.0853
R1394 B.n99 B.n98 10.0853
R1395 B.n451 B.n450 10.0853
R1396 B.n448 B.n447 10.0853
R1397 B.n807 B.n0 8.11757
R1398 B.n807 B.n1 8.11757
R1399 B.n587 B.n449 6.5566
R1400 B.n571 B.n570 6.5566
R1401 B.n222 B.n221 6.5566
R1402 B.n238 B.n100 6.5566
R1403 B.t13 B.n372 6.18428
R1404 B.n782 B.t9 6.18428
R1405 B.n747 B.t0 4.28158
R1406 B.n799 B.t6 4.28158
R1407 B.n590 B.n449 4.05904
R1408 B.n570 B.n569 4.05904
R1409 B.n221 B.n220 4.05904
R1410 B.n241 B.n100 4.05904
R1411 B.n364 B.t7 2.37888
R1412 B.n17 B.t1 2.37888
R1413 VN.n5 VN.t7 2471.19
R1414 VN.n1 VN.t1 2471.19
R1415 VN.n12 VN.t6 2471.19
R1416 VN.n8 VN.t4 2471.19
R1417 VN.n4 VN.t3 2430.29
R1418 VN.n2 VN.t5 2430.29
R1419 VN.n11 VN.t2 2430.29
R1420 VN.n9 VN.t0 2430.29
R1421 VN.n8 VN.n7 161.489
R1422 VN.n1 VN.n0 161.489
R1423 VN.n6 VN.n5 161.3
R1424 VN.n13 VN.n12 161.3
R1425 VN.n10 VN.n7 161.3
R1426 VN.n3 VN.n0 161.3
R1427 VN VN.n13 44.4721
R1428 VN.n3 VN.n2 37.9763
R1429 VN.n4 VN.n3 37.9763
R1430 VN.n11 VN.n10 37.9763
R1431 VN.n10 VN.n9 37.9763
R1432 VN.n2 VN.n1 35.055
R1433 VN.n5 VN.n4 35.055
R1434 VN.n12 VN.n11 35.055
R1435 VN.n9 VN.n8 35.055
R1436 VN.n13 VN.n7 0.189894
R1437 VN.n6 VN.n0 0.189894
R1438 VN VN.n6 0.0516364
R1439 VDD2.n2 VDD2.n1 60.2507
R1440 VDD2.n2 VDD2.n0 60.2507
R1441 VDD2 VDD2.n5 60.2479
R1442 VDD2.n4 VDD2.n3 60.0822
R1443 VDD2.n4 VDD2.n2 41.1205
R1444 VDD2.n5 VDD2.t7 1.10974
R1445 VDD2.n5 VDD2.t3 1.10974
R1446 VDD2.n3 VDD2.t1 1.10974
R1447 VDD2.n3 VDD2.t5 1.10974
R1448 VDD2.n1 VDD2.t4 1.10974
R1449 VDD2.n1 VDD2.t0 1.10974
R1450 VDD2.n0 VDD2.t6 1.10974
R1451 VDD2.n0 VDD2.t2 1.10974
R1452 VDD2 VDD2.n4 0.282828
C0 VP VN 5.79999f
C1 VDD1 VTAIL 28.774902f
C2 VDD1 VDD2 0.577749f
C3 VTAIL VDD2 28.813099f
C4 VDD1 VN 0.146868f
C5 VDD1 VP 3.71683f
C6 VTAIL VN 2.84048f
C7 VTAIL VP 2.85459f
C8 VDD2 VN 3.60115f
C9 VP VDD2 0.262718f
C10 VDD2 B 3.534835f
C11 VDD1 B 3.703358f
C12 VTAIL B 11.45969f
C13 VN B 7.83287f
C14 VP B 5.03589f
C15 VDD2.t6 B 0.549934f
C16 VDD2.t2 B 0.549934f
C17 VDD2.n0 B 5.00776f
C18 VDD2.t4 B 0.549934f
C19 VDD2.t0 B 0.549934f
C20 VDD2.n1 B 5.00776f
C21 VDD2.n2 B 3.49412f
C22 VDD2.t1 B 0.549934f
C23 VDD2.t5 B 0.549934f
C24 VDD2.n3 B 5.00658f
C25 VDD2.n4 B 4.00322f
C26 VDD2.t7 B 0.549934f
C27 VDD2.t3 B 0.549934f
C28 VDD2.n5 B 5.00771f
C29 VN.n0 B 0.1287f
C30 VN.t3 B 0.571503f
C31 VN.t5 B 0.571503f
C32 VN.t1 B 0.575154f
C33 VN.n1 B 0.237627f
C34 VN.n2 B 0.221734f
C35 VN.n3 B 0.020569f
C36 VN.n4 B 0.221734f
C37 VN.t7 B 0.575154f
C38 VN.n5 B 0.237546f
C39 VN.n6 B 0.04633f
C40 VN.n7 B 0.1287f
C41 VN.t6 B 0.575154f
C42 VN.t2 B 0.571503f
C43 VN.t0 B 0.571503f
C44 VN.t4 B 0.575154f
C45 VN.n8 B 0.237627f
C46 VN.n9 B 0.221734f
C47 VN.n10 B 0.020569f
C48 VN.n11 B 0.221734f
C49 VN.n12 B 0.237546f
C50 VN.n13 B 2.71152f
C51 VTAIL.t3 B 0.382712f
C52 VTAIL.t1 B 0.382712f
C53 VTAIL.n0 B 3.39917f
C54 VTAIL.n1 B 0.318829f
C55 VTAIL.t6 B 4.34175f
C56 VTAIL.n2 B 0.455998f
C57 VTAIL.t14 B 4.34175f
C58 VTAIL.n3 B 0.455998f
C59 VTAIL.t12 B 0.382712f
C60 VTAIL.t9 B 0.382712f
C61 VTAIL.n4 B 3.39917f
C62 VTAIL.n5 B 0.352933f
C63 VTAIL.t15 B 4.34175f
C64 VTAIL.n6 B 2.16796f
C65 VTAIL.t2 B 4.34176f
C66 VTAIL.n7 B 2.16796f
C67 VTAIL.t7 B 0.382712f
C68 VTAIL.t5 B 0.382712f
C69 VTAIL.n8 B 3.39918f
C70 VTAIL.n9 B 0.352928f
C71 VTAIL.t0 B 4.34176f
C72 VTAIL.n10 B 0.455993f
C73 VTAIL.t13 B 4.34176f
C74 VTAIL.n11 B 0.455993f
C75 VTAIL.t10 B 0.382712f
C76 VTAIL.t8 B 0.382712f
C77 VTAIL.n12 B 3.39918f
C78 VTAIL.n13 B 0.352928f
C79 VTAIL.t11 B 4.34175f
C80 VTAIL.n14 B 2.16796f
C81 VTAIL.t4 B 4.34175f
C82 VTAIL.n15 B 2.16287f
C83 VDD1.t1 B 0.549191f
C84 VDD1.t2 B 0.549191f
C85 VDD1.n0 B 5.00183f
C86 VDD1.t5 B 0.549191f
C87 VDD1.t0 B 0.549191f
C88 VDD1.n1 B 5.00099f
C89 VDD1.t7 B 0.549191f
C90 VDD1.t4 B 0.549191f
C91 VDD1.n2 B 5.00099f
C92 VDD1.n3 B 3.57254f
C93 VDD1.t6 B 0.549191f
C94 VDD1.t3 B 0.549191f
C95 VDD1.n4 B 4.99979f
C96 VDD1.n5 B 4.04388f
C97 VP.n0 B 0.061185f
C98 VP.t6 B 0.5849f
C99 VP.t3 B 0.5849f
C100 VP.t0 B 0.588637f
C101 VP.n1 B 0.131717f
C102 VP.t7 B 0.5849f
C103 VP.t5 B 0.5849f
C104 VP.t2 B 0.588637f
C105 VP.n2 B 0.243198f
C106 VP.n3 B 0.226932f
C107 VP.n4 B 0.021051f
C108 VP.n5 B 0.226932f
C109 VP.t4 B 0.588637f
C110 VP.n6 B 0.243115f
C111 VP.n7 B 2.73504f
C112 VP.n8 B 2.78492f
C113 VP.n9 B 0.243115f
C114 VP.n10 B 0.226932f
C115 VP.n11 B 0.021051f
C116 VP.n12 B 0.226932f
C117 VP.t1 B 0.588637f
C118 VP.n13 B 0.243115f
C119 VP.n14 B 0.047416f
.ends

