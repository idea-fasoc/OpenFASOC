* NGSPICE file created from diff_pair_sample_0789.ext - technology: sky130A

.subckt diff_pair_sample_0789 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=0 ps=0 w=7.91 l=1.7
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=3.0849 ps=16.6 w=7.91 l=1.7
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=3.0849 ps=16.6 w=7.91 l=1.7
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=3.0849 ps=16.6 w=7.91 l=1.7
X4 VDD2.t0 VN.t1 VTAIL.t1 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=3.0849 ps=16.6 w=7.91 l=1.7
X5 B.t8 B.t6 B.t7 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=0 ps=0 w=7.91 l=1.7
X6 B.t5 B.t3 B.t4 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=0 ps=0 w=7.91 l=1.7
X7 B.t2 B.t0 B.t1 w_n1782_n2550# sky130_fd_pr__pfet_01v8 ad=3.0849 pd=16.6 as=0 ps=0 w=7.91 l=1.7
R0 B.n315 B.n50 585
R1 B.n317 B.n316 585
R2 B.n318 B.n49 585
R3 B.n320 B.n319 585
R4 B.n321 B.n48 585
R5 B.n323 B.n322 585
R6 B.n324 B.n47 585
R7 B.n326 B.n325 585
R8 B.n327 B.n46 585
R9 B.n329 B.n328 585
R10 B.n330 B.n45 585
R11 B.n332 B.n331 585
R12 B.n333 B.n44 585
R13 B.n335 B.n334 585
R14 B.n336 B.n43 585
R15 B.n338 B.n337 585
R16 B.n339 B.n42 585
R17 B.n341 B.n340 585
R18 B.n342 B.n41 585
R19 B.n344 B.n343 585
R20 B.n345 B.n40 585
R21 B.n347 B.n346 585
R22 B.n348 B.n39 585
R23 B.n350 B.n349 585
R24 B.n351 B.n38 585
R25 B.n353 B.n352 585
R26 B.n354 B.n37 585
R27 B.n356 B.n355 585
R28 B.n357 B.n36 585
R29 B.n359 B.n358 585
R30 B.n361 B.n33 585
R31 B.n363 B.n362 585
R32 B.n364 B.n32 585
R33 B.n366 B.n365 585
R34 B.n367 B.n31 585
R35 B.n369 B.n368 585
R36 B.n370 B.n30 585
R37 B.n372 B.n371 585
R38 B.n373 B.n27 585
R39 B.n376 B.n375 585
R40 B.n377 B.n26 585
R41 B.n379 B.n378 585
R42 B.n380 B.n25 585
R43 B.n382 B.n381 585
R44 B.n383 B.n24 585
R45 B.n385 B.n384 585
R46 B.n386 B.n23 585
R47 B.n388 B.n387 585
R48 B.n389 B.n22 585
R49 B.n391 B.n390 585
R50 B.n392 B.n21 585
R51 B.n394 B.n393 585
R52 B.n395 B.n20 585
R53 B.n397 B.n396 585
R54 B.n398 B.n19 585
R55 B.n400 B.n399 585
R56 B.n401 B.n18 585
R57 B.n403 B.n402 585
R58 B.n404 B.n17 585
R59 B.n406 B.n405 585
R60 B.n407 B.n16 585
R61 B.n409 B.n408 585
R62 B.n410 B.n15 585
R63 B.n412 B.n411 585
R64 B.n413 B.n14 585
R65 B.n415 B.n414 585
R66 B.n416 B.n13 585
R67 B.n418 B.n417 585
R68 B.n419 B.n12 585
R69 B.n314 B.n313 585
R70 B.n312 B.n51 585
R71 B.n311 B.n310 585
R72 B.n309 B.n52 585
R73 B.n308 B.n307 585
R74 B.n306 B.n53 585
R75 B.n305 B.n304 585
R76 B.n303 B.n54 585
R77 B.n302 B.n301 585
R78 B.n300 B.n55 585
R79 B.n299 B.n298 585
R80 B.n297 B.n56 585
R81 B.n296 B.n295 585
R82 B.n294 B.n57 585
R83 B.n293 B.n292 585
R84 B.n291 B.n58 585
R85 B.n290 B.n289 585
R86 B.n288 B.n59 585
R87 B.n287 B.n286 585
R88 B.n285 B.n60 585
R89 B.n284 B.n283 585
R90 B.n282 B.n61 585
R91 B.n281 B.n280 585
R92 B.n279 B.n62 585
R93 B.n278 B.n277 585
R94 B.n276 B.n63 585
R95 B.n275 B.n274 585
R96 B.n273 B.n64 585
R97 B.n272 B.n271 585
R98 B.n270 B.n65 585
R99 B.n269 B.n268 585
R100 B.n267 B.n66 585
R101 B.n266 B.n265 585
R102 B.n264 B.n67 585
R103 B.n263 B.n262 585
R104 B.n261 B.n68 585
R105 B.n260 B.n259 585
R106 B.n258 B.n69 585
R107 B.n257 B.n256 585
R108 B.n255 B.n70 585
R109 B.n254 B.n253 585
R110 B.n149 B.n148 585
R111 B.n150 B.n109 585
R112 B.n152 B.n151 585
R113 B.n153 B.n108 585
R114 B.n155 B.n154 585
R115 B.n156 B.n107 585
R116 B.n158 B.n157 585
R117 B.n159 B.n106 585
R118 B.n161 B.n160 585
R119 B.n162 B.n105 585
R120 B.n164 B.n163 585
R121 B.n165 B.n104 585
R122 B.n167 B.n166 585
R123 B.n168 B.n103 585
R124 B.n170 B.n169 585
R125 B.n171 B.n102 585
R126 B.n173 B.n172 585
R127 B.n174 B.n101 585
R128 B.n176 B.n175 585
R129 B.n177 B.n100 585
R130 B.n179 B.n178 585
R131 B.n180 B.n99 585
R132 B.n182 B.n181 585
R133 B.n183 B.n98 585
R134 B.n185 B.n184 585
R135 B.n186 B.n97 585
R136 B.n188 B.n187 585
R137 B.n189 B.n96 585
R138 B.n191 B.n190 585
R139 B.n192 B.n93 585
R140 B.n195 B.n194 585
R141 B.n196 B.n92 585
R142 B.n198 B.n197 585
R143 B.n199 B.n91 585
R144 B.n201 B.n200 585
R145 B.n202 B.n90 585
R146 B.n204 B.n203 585
R147 B.n205 B.n89 585
R148 B.n207 B.n206 585
R149 B.n209 B.n208 585
R150 B.n210 B.n85 585
R151 B.n212 B.n211 585
R152 B.n213 B.n84 585
R153 B.n215 B.n214 585
R154 B.n216 B.n83 585
R155 B.n218 B.n217 585
R156 B.n219 B.n82 585
R157 B.n221 B.n220 585
R158 B.n222 B.n81 585
R159 B.n224 B.n223 585
R160 B.n225 B.n80 585
R161 B.n227 B.n226 585
R162 B.n228 B.n79 585
R163 B.n230 B.n229 585
R164 B.n231 B.n78 585
R165 B.n233 B.n232 585
R166 B.n234 B.n77 585
R167 B.n236 B.n235 585
R168 B.n237 B.n76 585
R169 B.n239 B.n238 585
R170 B.n240 B.n75 585
R171 B.n242 B.n241 585
R172 B.n243 B.n74 585
R173 B.n245 B.n244 585
R174 B.n246 B.n73 585
R175 B.n248 B.n247 585
R176 B.n249 B.n72 585
R177 B.n251 B.n250 585
R178 B.n252 B.n71 585
R179 B.n147 B.n110 585
R180 B.n146 B.n145 585
R181 B.n144 B.n111 585
R182 B.n143 B.n142 585
R183 B.n141 B.n112 585
R184 B.n140 B.n139 585
R185 B.n138 B.n113 585
R186 B.n137 B.n136 585
R187 B.n135 B.n114 585
R188 B.n134 B.n133 585
R189 B.n132 B.n115 585
R190 B.n131 B.n130 585
R191 B.n129 B.n116 585
R192 B.n128 B.n127 585
R193 B.n126 B.n117 585
R194 B.n125 B.n124 585
R195 B.n123 B.n118 585
R196 B.n122 B.n121 585
R197 B.n120 B.n119 585
R198 B.n2 B.n0 585
R199 B.n449 B.n1 585
R200 B.n448 B.n447 585
R201 B.n446 B.n3 585
R202 B.n445 B.n444 585
R203 B.n443 B.n4 585
R204 B.n442 B.n441 585
R205 B.n440 B.n5 585
R206 B.n439 B.n438 585
R207 B.n437 B.n6 585
R208 B.n436 B.n435 585
R209 B.n434 B.n7 585
R210 B.n433 B.n432 585
R211 B.n431 B.n8 585
R212 B.n430 B.n429 585
R213 B.n428 B.n9 585
R214 B.n427 B.n426 585
R215 B.n425 B.n10 585
R216 B.n424 B.n423 585
R217 B.n422 B.n11 585
R218 B.n421 B.n420 585
R219 B.n451 B.n450 585
R220 B.n148 B.n147 487.695
R221 B.n420 B.n419 487.695
R222 B.n254 B.n71 487.695
R223 B.n315 B.n314 487.695
R224 B.n86 B.t11 341.315
R225 B.n34 B.t7 341.315
R226 B.n94 B.t5 341.315
R227 B.n28 B.t1 341.315
R228 B.n86 B.t9 318.25
R229 B.n94 B.t3 318.25
R230 B.n28 B.t0 318.25
R231 B.n34 B.t6 318.25
R232 B.n87 B.t10 301.945
R233 B.n35 B.t8 301.945
R234 B.n95 B.t4 301.945
R235 B.n29 B.t2 301.945
R236 B.n147 B.n146 163.367
R237 B.n146 B.n111 163.367
R238 B.n142 B.n111 163.367
R239 B.n142 B.n141 163.367
R240 B.n141 B.n140 163.367
R241 B.n140 B.n113 163.367
R242 B.n136 B.n113 163.367
R243 B.n136 B.n135 163.367
R244 B.n135 B.n134 163.367
R245 B.n134 B.n115 163.367
R246 B.n130 B.n115 163.367
R247 B.n130 B.n129 163.367
R248 B.n129 B.n128 163.367
R249 B.n128 B.n117 163.367
R250 B.n124 B.n117 163.367
R251 B.n124 B.n123 163.367
R252 B.n123 B.n122 163.367
R253 B.n122 B.n119 163.367
R254 B.n119 B.n2 163.367
R255 B.n450 B.n2 163.367
R256 B.n450 B.n449 163.367
R257 B.n449 B.n448 163.367
R258 B.n448 B.n3 163.367
R259 B.n444 B.n3 163.367
R260 B.n444 B.n443 163.367
R261 B.n443 B.n442 163.367
R262 B.n442 B.n5 163.367
R263 B.n438 B.n5 163.367
R264 B.n438 B.n437 163.367
R265 B.n437 B.n436 163.367
R266 B.n436 B.n7 163.367
R267 B.n432 B.n7 163.367
R268 B.n432 B.n431 163.367
R269 B.n431 B.n430 163.367
R270 B.n430 B.n9 163.367
R271 B.n426 B.n9 163.367
R272 B.n426 B.n425 163.367
R273 B.n425 B.n424 163.367
R274 B.n424 B.n11 163.367
R275 B.n420 B.n11 163.367
R276 B.n148 B.n109 163.367
R277 B.n152 B.n109 163.367
R278 B.n153 B.n152 163.367
R279 B.n154 B.n153 163.367
R280 B.n154 B.n107 163.367
R281 B.n158 B.n107 163.367
R282 B.n159 B.n158 163.367
R283 B.n160 B.n159 163.367
R284 B.n160 B.n105 163.367
R285 B.n164 B.n105 163.367
R286 B.n165 B.n164 163.367
R287 B.n166 B.n165 163.367
R288 B.n166 B.n103 163.367
R289 B.n170 B.n103 163.367
R290 B.n171 B.n170 163.367
R291 B.n172 B.n171 163.367
R292 B.n172 B.n101 163.367
R293 B.n176 B.n101 163.367
R294 B.n177 B.n176 163.367
R295 B.n178 B.n177 163.367
R296 B.n178 B.n99 163.367
R297 B.n182 B.n99 163.367
R298 B.n183 B.n182 163.367
R299 B.n184 B.n183 163.367
R300 B.n184 B.n97 163.367
R301 B.n188 B.n97 163.367
R302 B.n189 B.n188 163.367
R303 B.n190 B.n189 163.367
R304 B.n190 B.n93 163.367
R305 B.n195 B.n93 163.367
R306 B.n196 B.n195 163.367
R307 B.n197 B.n196 163.367
R308 B.n197 B.n91 163.367
R309 B.n201 B.n91 163.367
R310 B.n202 B.n201 163.367
R311 B.n203 B.n202 163.367
R312 B.n203 B.n89 163.367
R313 B.n207 B.n89 163.367
R314 B.n208 B.n207 163.367
R315 B.n208 B.n85 163.367
R316 B.n212 B.n85 163.367
R317 B.n213 B.n212 163.367
R318 B.n214 B.n213 163.367
R319 B.n214 B.n83 163.367
R320 B.n218 B.n83 163.367
R321 B.n219 B.n218 163.367
R322 B.n220 B.n219 163.367
R323 B.n220 B.n81 163.367
R324 B.n224 B.n81 163.367
R325 B.n225 B.n224 163.367
R326 B.n226 B.n225 163.367
R327 B.n226 B.n79 163.367
R328 B.n230 B.n79 163.367
R329 B.n231 B.n230 163.367
R330 B.n232 B.n231 163.367
R331 B.n232 B.n77 163.367
R332 B.n236 B.n77 163.367
R333 B.n237 B.n236 163.367
R334 B.n238 B.n237 163.367
R335 B.n238 B.n75 163.367
R336 B.n242 B.n75 163.367
R337 B.n243 B.n242 163.367
R338 B.n244 B.n243 163.367
R339 B.n244 B.n73 163.367
R340 B.n248 B.n73 163.367
R341 B.n249 B.n248 163.367
R342 B.n250 B.n249 163.367
R343 B.n250 B.n71 163.367
R344 B.n255 B.n254 163.367
R345 B.n256 B.n255 163.367
R346 B.n256 B.n69 163.367
R347 B.n260 B.n69 163.367
R348 B.n261 B.n260 163.367
R349 B.n262 B.n261 163.367
R350 B.n262 B.n67 163.367
R351 B.n266 B.n67 163.367
R352 B.n267 B.n266 163.367
R353 B.n268 B.n267 163.367
R354 B.n268 B.n65 163.367
R355 B.n272 B.n65 163.367
R356 B.n273 B.n272 163.367
R357 B.n274 B.n273 163.367
R358 B.n274 B.n63 163.367
R359 B.n278 B.n63 163.367
R360 B.n279 B.n278 163.367
R361 B.n280 B.n279 163.367
R362 B.n280 B.n61 163.367
R363 B.n284 B.n61 163.367
R364 B.n285 B.n284 163.367
R365 B.n286 B.n285 163.367
R366 B.n286 B.n59 163.367
R367 B.n290 B.n59 163.367
R368 B.n291 B.n290 163.367
R369 B.n292 B.n291 163.367
R370 B.n292 B.n57 163.367
R371 B.n296 B.n57 163.367
R372 B.n297 B.n296 163.367
R373 B.n298 B.n297 163.367
R374 B.n298 B.n55 163.367
R375 B.n302 B.n55 163.367
R376 B.n303 B.n302 163.367
R377 B.n304 B.n303 163.367
R378 B.n304 B.n53 163.367
R379 B.n308 B.n53 163.367
R380 B.n309 B.n308 163.367
R381 B.n310 B.n309 163.367
R382 B.n310 B.n51 163.367
R383 B.n314 B.n51 163.367
R384 B.n419 B.n418 163.367
R385 B.n418 B.n13 163.367
R386 B.n414 B.n13 163.367
R387 B.n414 B.n413 163.367
R388 B.n413 B.n412 163.367
R389 B.n412 B.n15 163.367
R390 B.n408 B.n15 163.367
R391 B.n408 B.n407 163.367
R392 B.n407 B.n406 163.367
R393 B.n406 B.n17 163.367
R394 B.n402 B.n17 163.367
R395 B.n402 B.n401 163.367
R396 B.n401 B.n400 163.367
R397 B.n400 B.n19 163.367
R398 B.n396 B.n19 163.367
R399 B.n396 B.n395 163.367
R400 B.n395 B.n394 163.367
R401 B.n394 B.n21 163.367
R402 B.n390 B.n21 163.367
R403 B.n390 B.n389 163.367
R404 B.n389 B.n388 163.367
R405 B.n388 B.n23 163.367
R406 B.n384 B.n23 163.367
R407 B.n384 B.n383 163.367
R408 B.n383 B.n382 163.367
R409 B.n382 B.n25 163.367
R410 B.n378 B.n25 163.367
R411 B.n378 B.n377 163.367
R412 B.n377 B.n376 163.367
R413 B.n376 B.n27 163.367
R414 B.n371 B.n27 163.367
R415 B.n371 B.n370 163.367
R416 B.n370 B.n369 163.367
R417 B.n369 B.n31 163.367
R418 B.n365 B.n31 163.367
R419 B.n365 B.n364 163.367
R420 B.n364 B.n363 163.367
R421 B.n363 B.n33 163.367
R422 B.n358 B.n33 163.367
R423 B.n358 B.n357 163.367
R424 B.n357 B.n356 163.367
R425 B.n356 B.n37 163.367
R426 B.n352 B.n37 163.367
R427 B.n352 B.n351 163.367
R428 B.n351 B.n350 163.367
R429 B.n350 B.n39 163.367
R430 B.n346 B.n39 163.367
R431 B.n346 B.n345 163.367
R432 B.n345 B.n344 163.367
R433 B.n344 B.n41 163.367
R434 B.n340 B.n41 163.367
R435 B.n340 B.n339 163.367
R436 B.n339 B.n338 163.367
R437 B.n338 B.n43 163.367
R438 B.n334 B.n43 163.367
R439 B.n334 B.n333 163.367
R440 B.n333 B.n332 163.367
R441 B.n332 B.n45 163.367
R442 B.n328 B.n45 163.367
R443 B.n328 B.n327 163.367
R444 B.n327 B.n326 163.367
R445 B.n326 B.n47 163.367
R446 B.n322 B.n47 163.367
R447 B.n322 B.n321 163.367
R448 B.n321 B.n320 163.367
R449 B.n320 B.n49 163.367
R450 B.n316 B.n49 163.367
R451 B.n316 B.n315 163.367
R452 B.n88 B.n87 59.5399
R453 B.n193 B.n95 59.5399
R454 B.n374 B.n29 59.5399
R455 B.n360 B.n35 59.5399
R456 B.n87 B.n86 39.3702
R457 B.n95 B.n94 39.3702
R458 B.n29 B.n28 39.3702
R459 B.n35 B.n34 39.3702
R460 B.n421 B.n12 31.6883
R461 B.n313 B.n50 31.6883
R462 B.n253 B.n252 31.6883
R463 B.n149 B.n110 31.6883
R464 B B.n451 18.0485
R465 B.n417 B.n12 10.6151
R466 B.n417 B.n416 10.6151
R467 B.n416 B.n415 10.6151
R468 B.n415 B.n14 10.6151
R469 B.n411 B.n14 10.6151
R470 B.n411 B.n410 10.6151
R471 B.n410 B.n409 10.6151
R472 B.n409 B.n16 10.6151
R473 B.n405 B.n16 10.6151
R474 B.n405 B.n404 10.6151
R475 B.n404 B.n403 10.6151
R476 B.n403 B.n18 10.6151
R477 B.n399 B.n18 10.6151
R478 B.n399 B.n398 10.6151
R479 B.n398 B.n397 10.6151
R480 B.n397 B.n20 10.6151
R481 B.n393 B.n20 10.6151
R482 B.n393 B.n392 10.6151
R483 B.n392 B.n391 10.6151
R484 B.n391 B.n22 10.6151
R485 B.n387 B.n22 10.6151
R486 B.n387 B.n386 10.6151
R487 B.n386 B.n385 10.6151
R488 B.n385 B.n24 10.6151
R489 B.n381 B.n24 10.6151
R490 B.n381 B.n380 10.6151
R491 B.n380 B.n379 10.6151
R492 B.n379 B.n26 10.6151
R493 B.n375 B.n26 10.6151
R494 B.n373 B.n372 10.6151
R495 B.n372 B.n30 10.6151
R496 B.n368 B.n30 10.6151
R497 B.n368 B.n367 10.6151
R498 B.n367 B.n366 10.6151
R499 B.n366 B.n32 10.6151
R500 B.n362 B.n32 10.6151
R501 B.n362 B.n361 10.6151
R502 B.n359 B.n36 10.6151
R503 B.n355 B.n36 10.6151
R504 B.n355 B.n354 10.6151
R505 B.n354 B.n353 10.6151
R506 B.n353 B.n38 10.6151
R507 B.n349 B.n38 10.6151
R508 B.n349 B.n348 10.6151
R509 B.n348 B.n347 10.6151
R510 B.n347 B.n40 10.6151
R511 B.n343 B.n40 10.6151
R512 B.n343 B.n342 10.6151
R513 B.n342 B.n341 10.6151
R514 B.n341 B.n42 10.6151
R515 B.n337 B.n42 10.6151
R516 B.n337 B.n336 10.6151
R517 B.n336 B.n335 10.6151
R518 B.n335 B.n44 10.6151
R519 B.n331 B.n44 10.6151
R520 B.n331 B.n330 10.6151
R521 B.n330 B.n329 10.6151
R522 B.n329 B.n46 10.6151
R523 B.n325 B.n46 10.6151
R524 B.n325 B.n324 10.6151
R525 B.n324 B.n323 10.6151
R526 B.n323 B.n48 10.6151
R527 B.n319 B.n48 10.6151
R528 B.n319 B.n318 10.6151
R529 B.n318 B.n317 10.6151
R530 B.n317 B.n50 10.6151
R531 B.n253 B.n70 10.6151
R532 B.n257 B.n70 10.6151
R533 B.n258 B.n257 10.6151
R534 B.n259 B.n258 10.6151
R535 B.n259 B.n68 10.6151
R536 B.n263 B.n68 10.6151
R537 B.n264 B.n263 10.6151
R538 B.n265 B.n264 10.6151
R539 B.n265 B.n66 10.6151
R540 B.n269 B.n66 10.6151
R541 B.n270 B.n269 10.6151
R542 B.n271 B.n270 10.6151
R543 B.n271 B.n64 10.6151
R544 B.n275 B.n64 10.6151
R545 B.n276 B.n275 10.6151
R546 B.n277 B.n276 10.6151
R547 B.n277 B.n62 10.6151
R548 B.n281 B.n62 10.6151
R549 B.n282 B.n281 10.6151
R550 B.n283 B.n282 10.6151
R551 B.n283 B.n60 10.6151
R552 B.n287 B.n60 10.6151
R553 B.n288 B.n287 10.6151
R554 B.n289 B.n288 10.6151
R555 B.n289 B.n58 10.6151
R556 B.n293 B.n58 10.6151
R557 B.n294 B.n293 10.6151
R558 B.n295 B.n294 10.6151
R559 B.n295 B.n56 10.6151
R560 B.n299 B.n56 10.6151
R561 B.n300 B.n299 10.6151
R562 B.n301 B.n300 10.6151
R563 B.n301 B.n54 10.6151
R564 B.n305 B.n54 10.6151
R565 B.n306 B.n305 10.6151
R566 B.n307 B.n306 10.6151
R567 B.n307 B.n52 10.6151
R568 B.n311 B.n52 10.6151
R569 B.n312 B.n311 10.6151
R570 B.n313 B.n312 10.6151
R571 B.n150 B.n149 10.6151
R572 B.n151 B.n150 10.6151
R573 B.n151 B.n108 10.6151
R574 B.n155 B.n108 10.6151
R575 B.n156 B.n155 10.6151
R576 B.n157 B.n156 10.6151
R577 B.n157 B.n106 10.6151
R578 B.n161 B.n106 10.6151
R579 B.n162 B.n161 10.6151
R580 B.n163 B.n162 10.6151
R581 B.n163 B.n104 10.6151
R582 B.n167 B.n104 10.6151
R583 B.n168 B.n167 10.6151
R584 B.n169 B.n168 10.6151
R585 B.n169 B.n102 10.6151
R586 B.n173 B.n102 10.6151
R587 B.n174 B.n173 10.6151
R588 B.n175 B.n174 10.6151
R589 B.n175 B.n100 10.6151
R590 B.n179 B.n100 10.6151
R591 B.n180 B.n179 10.6151
R592 B.n181 B.n180 10.6151
R593 B.n181 B.n98 10.6151
R594 B.n185 B.n98 10.6151
R595 B.n186 B.n185 10.6151
R596 B.n187 B.n186 10.6151
R597 B.n187 B.n96 10.6151
R598 B.n191 B.n96 10.6151
R599 B.n192 B.n191 10.6151
R600 B.n194 B.n92 10.6151
R601 B.n198 B.n92 10.6151
R602 B.n199 B.n198 10.6151
R603 B.n200 B.n199 10.6151
R604 B.n200 B.n90 10.6151
R605 B.n204 B.n90 10.6151
R606 B.n205 B.n204 10.6151
R607 B.n206 B.n205 10.6151
R608 B.n210 B.n209 10.6151
R609 B.n211 B.n210 10.6151
R610 B.n211 B.n84 10.6151
R611 B.n215 B.n84 10.6151
R612 B.n216 B.n215 10.6151
R613 B.n217 B.n216 10.6151
R614 B.n217 B.n82 10.6151
R615 B.n221 B.n82 10.6151
R616 B.n222 B.n221 10.6151
R617 B.n223 B.n222 10.6151
R618 B.n223 B.n80 10.6151
R619 B.n227 B.n80 10.6151
R620 B.n228 B.n227 10.6151
R621 B.n229 B.n228 10.6151
R622 B.n229 B.n78 10.6151
R623 B.n233 B.n78 10.6151
R624 B.n234 B.n233 10.6151
R625 B.n235 B.n234 10.6151
R626 B.n235 B.n76 10.6151
R627 B.n239 B.n76 10.6151
R628 B.n240 B.n239 10.6151
R629 B.n241 B.n240 10.6151
R630 B.n241 B.n74 10.6151
R631 B.n245 B.n74 10.6151
R632 B.n246 B.n245 10.6151
R633 B.n247 B.n246 10.6151
R634 B.n247 B.n72 10.6151
R635 B.n251 B.n72 10.6151
R636 B.n252 B.n251 10.6151
R637 B.n145 B.n110 10.6151
R638 B.n145 B.n144 10.6151
R639 B.n144 B.n143 10.6151
R640 B.n143 B.n112 10.6151
R641 B.n139 B.n112 10.6151
R642 B.n139 B.n138 10.6151
R643 B.n138 B.n137 10.6151
R644 B.n137 B.n114 10.6151
R645 B.n133 B.n114 10.6151
R646 B.n133 B.n132 10.6151
R647 B.n132 B.n131 10.6151
R648 B.n131 B.n116 10.6151
R649 B.n127 B.n116 10.6151
R650 B.n127 B.n126 10.6151
R651 B.n126 B.n125 10.6151
R652 B.n125 B.n118 10.6151
R653 B.n121 B.n118 10.6151
R654 B.n121 B.n120 10.6151
R655 B.n120 B.n0 10.6151
R656 B.n447 B.n1 10.6151
R657 B.n447 B.n446 10.6151
R658 B.n446 B.n445 10.6151
R659 B.n445 B.n4 10.6151
R660 B.n441 B.n4 10.6151
R661 B.n441 B.n440 10.6151
R662 B.n440 B.n439 10.6151
R663 B.n439 B.n6 10.6151
R664 B.n435 B.n6 10.6151
R665 B.n435 B.n434 10.6151
R666 B.n434 B.n433 10.6151
R667 B.n433 B.n8 10.6151
R668 B.n429 B.n8 10.6151
R669 B.n429 B.n428 10.6151
R670 B.n428 B.n427 10.6151
R671 B.n427 B.n10 10.6151
R672 B.n423 B.n10 10.6151
R673 B.n423 B.n422 10.6151
R674 B.n422 B.n421 10.6151
R675 B.n374 B.n373 6.5566
R676 B.n361 B.n360 6.5566
R677 B.n194 B.n193 6.5566
R678 B.n206 B.n88 6.5566
R679 B.n375 B.n374 4.05904
R680 B.n360 B.n359 4.05904
R681 B.n193 B.n192 4.05904
R682 B.n209 B.n88 4.05904
R683 B.n451 B.n0 2.81026
R684 B.n451 B.n1 2.81026
R685 VP.n0 VP.t0 210.168
R686 VP.n0 VP.t1 170.998
R687 VP VP.n0 0.241678
R688 VTAIL.n162 VTAIL.n126 756.745
R689 VTAIL.n36 VTAIL.n0 756.745
R690 VTAIL.n120 VTAIL.n84 756.745
R691 VTAIL.n78 VTAIL.n42 756.745
R692 VTAIL.n138 VTAIL.n137 585
R693 VTAIL.n143 VTAIL.n142 585
R694 VTAIL.n145 VTAIL.n144 585
R695 VTAIL.n134 VTAIL.n133 585
R696 VTAIL.n151 VTAIL.n150 585
R697 VTAIL.n153 VTAIL.n152 585
R698 VTAIL.n130 VTAIL.n129 585
R699 VTAIL.n160 VTAIL.n159 585
R700 VTAIL.n161 VTAIL.n128 585
R701 VTAIL.n163 VTAIL.n162 585
R702 VTAIL.n12 VTAIL.n11 585
R703 VTAIL.n17 VTAIL.n16 585
R704 VTAIL.n19 VTAIL.n18 585
R705 VTAIL.n8 VTAIL.n7 585
R706 VTAIL.n25 VTAIL.n24 585
R707 VTAIL.n27 VTAIL.n26 585
R708 VTAIL.n4 VTAIL.n3 585
R709 VTAIL.n34 VTAIL.n33 585
R710 VTAIL.n35 VTAIL.n2 585
R711 VTAIL.n37 VTAIL.n36 585
R712 VTAIL.n121 VTAIL.n120 585
R713 VTAIL.n119 VTAIL.n86 585
R714 VTAIL.n118 VTAIL.n117 585
R715 VTAIL.n89 VTAIL.n87 585
R716 VTAIL.n112 VTAIL.n111 585
R717 VTAIL.n110 VTAIL.n109 585
R718 VTAIL.n93 VTAIL.n92 585
R719 VTAIL.n104 VTAIL.n103 585
R720 VTAIL.n102 VTAIL.n101 585
R721 VTAIL.n97 VTAIL.n96 585
R722 VTAIL.n79 VTAIL.n78 585
R723 VTAIL.n77 VTAIL.n44 585
R724 VTAIL.n76 VTAIL.n75 585
R725 VTAIL.n47 VTAIL.n45 585
R726 VTAIL.n70 VTAIL.n69 585
R727 VTAIL.n68 VTAIL.n67 585
R728 VTAIL.n51 VTAIL.n50 585
R729 VTAIL.n62 VTAIL.n61 585
R730 VTAIL.n60 VTAIL.n59 585
R731 VTAIL.n55 VTAIL.n54 585
R732 VTAIL.n139 VTAIL.t1 329.043
R733 VTAIL.n13 VTAIL.t2 329.043
R734 VTAIL.n98 VTAIL.t3 329.043
R735 VTAIL.n56 VTAIL.t0 329.043
R736 VTAIL.n143 VTAIL.n137 171.744
R737 VTAIL.n144 VTAIL.n143 171.744
R738 VTAIL.n144 VTAIL.n133 171.744
R739 VTAIL.n151 VTAIL.n133 171.744
R740 VTAIL.n152 VTAIL.n151 171.744
R741 VTAIL.n152 VTAIL.n129 171.744
R742 VTAIL.n160 VTAIL.n129 171.744
R743 VTAIL.n161 VTAIL.n160 171.744
R744 VTAIL.n162 VTAIL.n161 171.744
R745 VTAIL.n17 VTAIL.n11 171.744
R746 VTAIL.n18 VTAIL.n17 171.744
R747 VTAIL.n18 VTAIL.n7 171.744
R748 VTAIL.n25 VTAIL.n7 171.744
R749 VTAIL.n26 VTAIL.n25 171.744
R750 VTAIL.n26 VTAIL.n3 171.744
R751 VTAIL.n34 VTAIL.n3 171.744
R752 VTAIL.n35 VTAIL.n34 171.744
R753 VTAIL.n36 VTAIL.n35 171.744
R754 VTAIL.n120 VTAIL.n119 171.744
R755 VTAIL.n119 VTAIL.n118 171.744
R756 VTAIL.n118 VTAIL.n87 171.744
R757 VTAIL.n111 VTAIL.n87 171.744
R758 VTAIL.n111 VTAIL.n110 171.744
R759 VTAIL.n110 VTAIL.n92 171.744
R760 VTAIL.n103 VTAIL.n92 171.744
R761 VTAIL.n103 VTAIL.n102 171.744
R762 VTAIL.n102 VTAIL.n96 171.744
R763 VTAIL.n78 VTAIL.n77 171.744
R764 VTAIL.n77 VTAIL.n76 171.744
R765 VTAIL.n76 VTAIL.n45 171.744
R766 VTAIL.n69 VTAIL.n45 171.744
R767 VTAIL.n69 VTAIL.n68 171.744
R768 VTAIL.n68 VTAIL.n50 171.744
R769 VTAIL.n61 VTAIL.n50 171.744
R770 VTAIL.n61 VTAIL.n60 171.744
R771 VTAIL.n60 VTAIL.n54 171.744
R772 VTAIL.t1 VTAIL.n137 85.8723
R773 VTAIL.t2 VTAIL.n11 85.8723
R774 VTAIL.t3 VTAIL.n96 85.8723
R775 VTAIL.t0 VTAIL.n54 85.8723
R776 VTAIL.n167 VTAIL.n166 34.3187
R777 VTAIL.n41 VTAIL.n40 34.3187
R778 VTAIL.n125 VTAIL.n124 34.3187
R779 VTAIL.n83 VTAIL.n82 34.3187
R780 VTAIL.n83 VTAIL.n41 22.6858
R781 VTAIL.n167 VTAIL.n125 20.9358
R782 VTAIL.n163 VTAIL.n128 13.1884
R783 VTAIL.n37 VTAIL.n2 13.1884
R784 VTAIL.n121 VTAIL.n86 13.1884
R785 VTAIL.n79 VTAIL.n44 13.1884
R786 VTAIL.n159 VTAIL.n158 12.8005
R787 VTAIL.n164 VTAIL.n126 12.8005
R788 VTAIL.n33 VTAIL.n32 12.8005
R789 VTAIL.n38 VTAIL.n0 12.8005
R790 VTAIL.n122 VTAIL.n84 12.8005
R791 VTAIL.n117 VTAIL.n88 12.8005
R792 VTAIL.n80 VTAIL.n42 12.8005
R793 VTAIL.n75 VTAIL.n46 12.8005
R794 VTAIL.n157 VTAIL.n130 12.0247
R795 VTAIL.n31 VTAIL.n4 12.0247
R796 VTAIL.n116 VTAIL.n89 12.0247
R797 VTAIL.n74 VTAIL.n47 12.0247
R798 VTAIL.n154 VTAIL.n153 11.249
R799 VTAIL.n28 VTAIL.n27 11.249
R800 VTAIL.n113 VTAIL.n112 11.249
R801 VTAIL.n71 VTAIL.n70 11.249
R802 VTAIL.n139 VTAIL.n138 10.7238
R803 VTAIL.n13 VTAIL.n12 10.7238
R804 VTAIL.n98 VTAIL.n97 10.7238
R805 VTAIL.n56 VTAIL.n55 10.7238
R806 VTAIL.n150 VTAIL.n132 10.4732
R807 VTAIL.n24 VTAIL.n6 10.4732
R808 VTAIL.n109 VTAIL.n91 10.4732
R809 VTAIL.n67 VTAIL.n49 10.4732
R810 VTAIL.n149 VTAIL.n134 9.69747
R811 VTAIL.n23 VTAIL.n8 9.69747
R812 VTAIL.n108 VTAIL.n93 9.69747
R813 VTAIL.n66 VTAIL.n51 9.69747
R814 VTAIL.n166 VTAIL.n165 9.45567
R815 VTAIL.n40 VTAIL.n39 9.45567
R816 VTAIL.n124 VTAIL.n123 9.45567
R817 VTAIL.n82 VTAIL.n81 9.45567
R818 VTAIL.n165 VTAIL.n164 9.3005
R819 VTAIL.n141 VTAIL.n140 9.3005
R820 VTAIL.n136 VTAIL.n135 9.3005
R821 VTAIL.n147 VTAIL.n146 9.3005
R822 VTAIL.n149 VTAIL.n148 9.3005
R823 VTAIL.n132 VTAIL.n131 9.3005
R824 VTAIL.n155 VTAIL.n154 9.3005
R825 VTAIL.n157 VTAIL.n156 9.3005
R826 VTAIL.n158 VTAIL.n127 9.3005
R827 VTAIL.n39 VTAIL.n38 9.3005
R828 VTAIL.n15 VTAIL.n14 9.3005
R829 VTAIL.n10 VTAIL.n9 9.3005
R830 VTAIL.n21 VTAIL.n20 9.3005
R831 VTAIL.n23 VTAIL.n22 9.3005
R832 VTAIL.n6 VTAIL.n5 9.3005
R833 VTAIL.n29 VTAIL.n28 9.3005
R834 VTAIL.n31 VTAIL.n30 9.3005
R835 VTAIL.n32 VTAIL.n1 9.3005
R836 VTAIL.n100 VTAIL.n99 9.3005
R837 VTAIL.n95 VTAIL.n94 9.3005
R838 VTAIL.n106 VTAIL.n105 9.3005
R839 VTAIL.n108 VTAIL.n107 9.3005
R840 VTAIL.n91 VTAIL.n90 9.3005
R841 VTAIL.n114 VTAIL.n113 9.3005
R842 VTAIL.n116 VTAIL.n115 9.3005
R843 VTAIL.n88 VTAIL.n85 9.3005
R844 VTAIL.n123 VTAIL.n122 9.3005
R845 VTAIL.n58 VTAIL.n57 9.3005
R846 VTAIL.n53 VTAIL.n52 9.3005
R847 VTAIL.n64 VTAIL.n63 9.3005
R848 VTAIL.n66 VTAIL.n65 9.3005
R849 VTAIL.n49 VTAIL.n48 9.3005
R850 VTAIL.n72 VTAIL.n71 9.3005
R851 VTAIL.n74 VTAIL.n73 9.3005
R852 VTAIL.n46 VTAIL.n43 9.3005
R853 VTAIL.n81 VTAIL.n80 9.3005
R854 VTAIL.n146 VTAIL.n145 8.92171
R855 VTAIL.n20 VTAIL.n19 8.92171
R856 VTAIL.n105 VTAIL.n104 8.92171
R857 VTAIL.n63 VTAIL.n62 8.92171
R858 VTAIL.n142 VTAIL.n136 8.14595
R859 VTAIL.n16 VTAIL.n10 8.14595
R860 VTAIL.n101 VTAIL.n95 8.14595
R861 VTAIL.n59 VTAIL.n53 8.14595
R862 VTAIL.n141 VTAIL.n138 7.3702
R863 VTAIL.n15 VTAIL.n12 7.3702
R864 VTAIL.n100 VTAIL.n97 7.3702
R865 VTAIL.n58 VTAIL.n55 7.3702
R866 VTAIL.n142 VTAIL.n141 5.81868
R867 VTAIL.n16 VTAIL.n15 5.81868
R868 VTAIL.n101 VTAIL.n100 5.81868
R869 VTAIL.n59 VTAIL.n58 5.81868
R870 VTAIL.n145 VTAIL.n136 5.04292
R871 VTAIL.n19 VTAIL.n10 5.04292
R872 VTAIL.n104 VTAIL.n95 5.04292
R873 VTAIL.n62 VTAIL.n53 5.04292
R874 VTAIL.n146 VTAIL.n134 4.26717
R875 VTAIL.n20 VTAIL.n8 4.26717
R876 VTAIL.n105 VTAIL.n93 4.26717
R877 VTAIL.n63 VTAIL.n51 4.26717
R878 VTAIL.n150 VTAIL.n149 3.49141
R879 VTAIL.n24 VTAIL.n23 3.49141
R880 VTAIL.n109 VTAIL.n108 3.49141
R881 VTAIL.n67 VTAIL.n66 3.49141
R882 VTAIL.n153 VTAIL.n132 2.71565
R883 VTAIL.n27 VTAIL.n6 2.71565
R884 VTAIL.n112 VTAIL.n91 2.71565
R885 VTAIL.n70 VTAIL.n49 2.71565
R886 VTAIL.n140 VTAIL.n139 2.4129
R887 VTAIL.n14 VTAIL.n13 2.4129
R888 VTAIL.n99 VTAIL.n98 2.4129
R889 VTAIL.n57 VTAIL.n56 2.4129
R890 VTAIL.n154 VTAIL.n130 1.93989
R891 VTAIL.n28 VTAIL.n4 1.93989
R892 VTAIL.n113 VTAIL.n89 1.93989
R893 VTAIL.n71 VTAIL.n47 1.93989
R894 VTAIL.n125 VTAIL.n83 1.34533
R895 VTAIL.n159 VTAIL.n157 1.16414
R896 VTAIL.n166 VTAIL.n126 1.16414
R897 VTAIL.n33 VTAIL.n31 1.16414
R898 VTAIL.n40 VTAIL.n0 1.16414
R899 VTAIL.n124 VTAIL.n84 1.16414
R900 VTAIL.n117 VTAIL.n116 1.16414
R901 VTAIL.n82 VTAIL.n42 1.16414
R902 VTAIL.n75 VTAIL.n74 1.16414
R903 VTAIL VTAIL.n41 0.966017
R904 VTAIL.n158 VTAIL.n128 0.388379
R905 VTAIL.n164 VTAIL.n163 0.388379
R906 VTAIL.n32 VTAIL.n2 0.388379
R907 VTAIL.n38 VTAIL.n37 0.388379
R908 VTAIL.n122 VTAIL.n121 0.388379
R909 VTAIL.n88 VTAIL.n86 0.388379
R910 VTAIL.n80 VTAIL.n79 0.388379
R911 VTAIL.n46 VTAIL.n44 0.388379
R912 VTAIL VTAIL.n167 0.37981
R913 VTAIL.n140 VTAIL.n135 0.155672
R914 VTAIL.n147 VTAIL.n135 0.155672
R915 VTAIL.n148 VTAIL.n147 0.155672
R916 VTAIL.n148 VTAIL.n131 0.155672
R917 VTAIL.n155 VTAIL.n131 0.155672
R918 VTAIL.n156 VTAIL.n155 0.155672
R919 VTAIL.n156 VTAIL.n127 0.155672
R920 VTAIL.n165 VTAIL.n127 0.155672
R921 VTAIL.n14 VTAIL.n9 0.155672
R922 VTAIL.n21 VTAIL.n9 0.155672
R923 VTAIL.n22 VTAIL.n21 0.155672
R924 VTAIL.n22 VTAIL.n5 0.155672
R925 VTAIL.n29 VTAIL.n5 0.155672
R926 VTAIL.n30 VTAIL.n29 0.155672
R927 VTAIL.n30 VTAIL.n1 0.155672
R928 VTAIL.n39 VTAIL.n1 0.155672
R929 VTAIL.n123 VTAIL.n85 0.155672
R930 VTAIL.n115 VTAIL.n85 0.155672
R931 VTAIL.n115 VTAIL.n114 0.155672
R932 VTAIL.n114 VTAIL.n90 0.155672
R933 VTAIL.n107 VTAIL.n90 0.155672
R934 VTAIL.n107 VTAIL.n106 0.155672
R935 VTAIL.n106 VTAIL.n94 0.155672
R936 VTAIL.n99 VTAIL.n94 0.155672
R937 VTAIL.n81 VTAIL.n43 0.155672
R938 VTAIL.n73 VTAIL.n43 0.155672
R939 VTAIL.n73 VTAIL.n72 0.155672
R940 VTAIL.n72 VTAIL.n48 0.155672
R941 VTAIL.n65 VTAIL.n48 0.155672
R942 VTAIL.n65 VTAIL.n64 0.155672
R943 VTAIL.n64 VTAIL.n52 0.155672
R944 VTAIL.n57 VTAIL.n52 0.155672
R945 VDD1.n36 VDD1.n0 756.745
R946 VDD1.n77 VDD1.n41 756.745
R947 VDD1.n37 VDD1.n36 585
R948 VDD1.n35 VDD1.n2 585
R949 VDD1.n34 VDD1.n33 585
R950 VDD1.n5 VDD1.n3 585
R951 VDD1.n28 VDD1.n27 585
R952 VDD1.n26 VDD1.n25 585
R953 VDD1.n9 VDD1.n8 585
R954 VDD1.n20 VDD1.n19 585
R955 VDD1.n18 VDD1.n17 585
R956 VDD1.n13 VDD1.n12 585
R957 VDD1.n53 VDD1.n52 585
R958 VDD1.n58 VDD1.n57 585
R959 VDD1.n60 VDD1.n59 585
R960 VDD1.n49 VDD1.n48 585
R961 VDD1.n66 VDD1.n65 585
R962 VDD1.n68 VDD1.n67 585
R963 VDD1.n45 VDD1.n44 585
R964 VDD1.n75 VDD1.n74 585
R965 VDD1.n76 VDD1.n43 585
R966 VDD1.n78 VDD1.n77 585
R967 VDD1.n14 VDD1.t1 329.043
R968 VDD1.n54 VDD1.t0 329.043
R969 VDD1.n36 VDD1.n35 171.744
R970 VDD1.n35 VDD1.n34 171.744
R971 VDD1.n34 VDD1.n3 171.744
R972 VDD1.n27 VDD1.n3 171.744
R973 VDD1.n27 VDD1.n26 171.744
R974 VDD1.n26 VDD1.n8 171.744
R975 VDD1.n19 VDD1.n8 171.744
R976 VDD1.n19 VDD1.n18 171.744
R977 VDD1.n18 VDD1.n12 171.744
R978 VDD1.n58 VDD1.n52 171.744
R979 VDD1.n59 VDD1.n58 171.744
R980 VDD1.n59 VDD1.n48 171.744
R981 VDD1.n66 VDD1.n48 171.744
R982 VDD1.n67 VDD1.n66 171.744
R983 VDD1.n67 VDD1.n44 171.744
R984 VDD1.n75 VDD1.n44 171.744
R985 VDD1.n76 VDD1.n75 171.744
R986 VDD1.n77 VDD1.n76 171.744
R987 VDD1 VDD1.n81 85.9382
R988 VDD1.t1 VDD1.n12 85.8723
R989 VDD1.t0 VDD1.n52 85.8723
R990 VDD1 VDD1.n40 51.4932
R991 VDD1.n37 VDD1.n2 13.1884
R992 VDD1.n78 VDD1.n43 13.1884
R993 VDD1.n38 VDD1.n0 12.8005
R994 VDD1.n33 VDD1.n4 12.8005
R995 VDD1.n74 VDD1.n73 12.8005
R996 VDD1.n79 VDD1.n41 12.8005
R997 VDD1.n32 VDD1.n5 12.0247
R998 VDD1.n72 VDD1.n45 12.0247
R999 VDD1.n29 VDD1.n28 11.249
R1000 VDD1.n69 VDD1.n68 11.249
R1001 VDD1.n14 VDD1.n13 10.7238
R1002 VDD1.n54 VDD1.n53 10.7238
R1003 VDD1.n25 VDD1.n7 10.4732
R1004 VDD1.n65 VDD1.n47 10.4732
R1005 VDD1.n24 VDD1.n9 9.69747
R1006 VDD1.n64 VDD1.n49 9.69747
R1007 VDD1.n40 VDD1.n39 9.45567
R1008 VDD1.n81 VDD1.n80 9.45567
R1009 VDD1.n16 VDD1.n15 9.3005
R1010 VDD1.n11 VDD1.n10 9.3005
R1011 VDD1.n22 VDD1.n21 9.3005
R1012 VDD1.n24 VDD1.n23 9.3005
R1013 VDD1.n7 VDD1.n6 9.3005
R1014 VDD1.n30 VDD1.n29 9.3005
R1015 VDD1.n32 VDD1.n31 9.3005
R1016 VDD1.n4 VDD1.n1 9.3005
R1017 VDD1.n39 VDD1.n38 9.3005
R1018 VDD1.n80 VDD1.n79 9.3005
R1019 VDD1.n56 VDD1.n55 9.3005
R1020 VDD1.n51 VDD1.n50 9.3005
R1021 VDD1.n62 VDD1.n61 9.3005
R1022 VDD1.n64 VDD1.n63 9.3005
R1023 VDD1.n47 VDD1.n46 9.3005
R1024 VDD1.n70 VDD1.n69 9.3005
R1025 VDD1.n72 VDD1.n71 9.3005
R1026 VDD1.n73 VDD1.n42 9.3005
R1027 VDD1.n21 VDD1.n20 8.92171
R1028 VDD1.n61 VDD1.n60 8.92171
R1029 VDD1.n17 VDD1.n11 8.14595
R1030 VDD1.n57 VDD1.n51 8.14595
R1031 VDD1.n16 VDD1.n13 7.3702
R1032 VDD1.n56 VDD1.n53 7.3702
R1033 VDD1.n17 VDD1.n16 5.81868
R1034 VDD1.n57 VDD1.n56 5.81868
R1035 VDD1.n20 VDD1.n11 5.04292
R1036 VDD1.n60 VDD1.n51 5.04292
R1037 VDD1.n21 VDD1.n9 4.26717
R1038 VDD1.n61 VDD1.n49 4.26717
R1039 VDD1.n25 VDD1.n24 3.49141
R1040 VDD1.n65 VDD1.n64 3.49141
R1041 VDD1.n28 VDD1.n7 2.71565
R1042 VDD1.n68 VDD1.n47 2.71565
R1043 VDD1.n15 VDD1.n14 2.4129
R1044 VDD1.n55 VDD1.n54 2.4129
R1045 VDD1.n29 VDD1.n5 1.93989
R1046 VDD1.n69 VDD1.n45 1.93989
R1047 VDD1.n40 VDD1.n0 1.16414
R1048 VDD1.n33 VDD1.n32 1.16414
R1049 VDD1.n74 VDD1.n72 1.16414
R1050 VDD1.n81 VDD1.n41 1.16414
R1051 VDD1.n38 VDD1.n37 0.388379
R1052 VDD1.n4 VDD1.n2 0.388379
R1053 VDD1.n73 VDD1.n43 0.388379
R1054 VDD1.n79 VDD1.n78 0.388379
R1055 VDD1.n39 VDD1.n1 0.155672
R1056 VDD1.n31 VDD1.n1 0.155672
R1057 VDD1.n31 VDD1.n30 0.155672
R1058 VDD1.n30 VDD1.n6 0.155672
R1059 VDD1.n23 VDD1.n6 0.155672
R1060 VDD1.n23 VDD1.n22 0.155672
R1061 VDD1.n22 VDD1.n10 0.155672
R1062 VDD1.n15 VDD1.n10 0.155672
R1063 VDD1.n55 VDD1.n50 0.155672
R1064 VDD1.n62 VDD1.n50 0.155672
R1065 VDD1.n63 VDD1.n62 0.155672
R1066 VDD1.n63 VDD1.n46 0.155672
R1067 VDD1.n70 VDD1.n46 0.155672
R1068 VDD1.n71 VDD1.n70 0.155672
R1069 VDD1.n71 VDD1.n42 0.155672
R1070 VDD1.n80 VDD1.n42 0.155672
R1071 VN VN.t0 210.359
R1072 VN VN.t1 171.238
R1073 VDD2.n77 VDD2.n41 756.745
R1074 VDD2.n36 VDD2.n0 756.745
R1075 VDD2.n78 VDD2.n77 585
R1076 VDD2.n76 VDD2.n43 585
R1077 VDD2.n75 VDD2.n74 585
R1078 VDD2.n46 VDD2.n44 585
R1079 VDD2.n69 VDD2.n68 585
R1080 VDD2.n67 VDD2.n66 585
R1081 VDD2.n50 VDD2.n49 585
R1082 VDD2.n61 VDD2.n60 585
R1083 VDD2.n59 VDD2.n58 585
R1084 VDD2.n54 VDD2.n53 585
R1085 VDD2.n12 VDD2.n11 585
R1086 VDD2.n17 VDD2.n16 585
R1087 VDD2.n19 VDD2.n18 585
R1088 VDD2.n8 VDD2.n7 585
R1089 VDD2.n25 VDD2.n24 585
R1090 VDD2.n27 VDD2.n26 585
R1091 VDD2.n4 VDD2.n3 585
R1092 VDD2.n34 VDD2.n33 585
R1093 VDD2.n35 VDD2.n2 585
R1094 VDD2.n37 VDD2.n36 585
R1095 VDD2.n55 VDD2.t1 329.043
R1096 VDD2.n13 VDD2.t0 329.043
R1097 VDD2.n77 VDD2.n76 171.744
R1098 VDD2.n76 VDD2.n75 171.744
R1099 VDD2.n75 VDD2.n44 171.744
R1100 VDD2.n68 VDD2.n44 171.744
R1101 VDD2.n68 VDD2.n67 171.744
R1102 VDD2.n67 VDD2.n49 171.744
R1103 VDD2.n60 VDD2.n49 171.744
R1104 VDD2.n60 VDD2.n59 171.744
R1105 VDD2.n59 VDD2.n53 171.744
R1106 VDD2.n17 VDD2.n11 171.744
R1107 VDD2.n18 VDD2.n17 171.744
R1108 VDD2.n18 VDD2.n7 171.744
R1109 VDD2.n25 VDD2.n7 171.744
R1110 VDD2.n26 VDD2.n25 171.744
R1111 VDD2.n26 VDD2.n3 171.744
R1112 VDD2.n34 VDD2.n3 171.744
R1113 VDD2.n35 VDD2.n34 171.744
R1114 VDD2.n36 VDD2.n35 171.744
R1115 VDD2.t1 VDD2.n53 85.8723
R1116 VDD2.t0 VDD2.n11 85.8723
R1117 VDD2.n82 VDD2.n40 84.9759
R1118 VDD2.n82 VDD2.n81 50.9975
R1119 VDD2.n78 VDD2.n43 13.1884
R1120 VDD2.n37 VDD2.n2 13.1884
R1121 VDD2.n79 VDD2.n41 12.8005
R1122 VDD2.n74 VDD2.n45 12.8005
R1123 VDD2.n33 VDD2.n32 12.8005
R1124 VDD2.n38 VDD2.n0 12.8005
R1125 VDD2.n73 VDD2.n46 12.0247
R1126 VDD2.n31 VDD2.n4 12.0247
R1127 VDD2.n70 VDD2.n69 11.249
R1128 VDD2.n28 VDD2.n27 11.249
R1129 VDD2.n55 VDD2.n54 10.7238
R1130 VDD2.n13 VDD2.n12 10.7238
R1131 VDD2.n66 VDD2.n48 10.4732
R1132 VDD2.n24 VDD2.n6 10.4732
R1133 VDD2.n65 VDD2.n50 9.69747
R1134 VDD2.n23 VDD2.n8 9.69747
R1135 VDD2.n81 VDD2.n80 9.45567
R1136 VDD2.n40 VDD2.n39 9.45567
R1137 VDD2.n57 VDD2.n56 9.3005
R1138 VDD2.n52 VDD2.n51 9.3005
R1139 VDD2.n63 VDD2.n62 9.3005
R1140 VDD2.n65 VDD2.n64 9.3005
R1141 VDD2.n48 VDD2.n47 9.3005
R1142 VDD2.n71 VDD2.n70 9.3005
R1143 VDD2.n73 VDD2.n72 9.3005
R1144 VDD2.n45 VDD2.n42 9.3005
R1145 VDD2.n80 VDD2.n79 9.3005
R1146 VDD2.n39 VDD2.n38 9.3005
R1147 VDD2.n15 VDD2.n14 9.3005
R1148 VDD2.n10 VDD2.n9 9.3005
R1149 VDD2.n21 VDD2.n20 9.3005
R1150 VDD2.n23 VDD2.n22 9.3005
R1151 VDD2.n6 VDD2.n5 9.3005
R1152 VDD2.n29 VDD2.n28 9.3005
R1153 VDD2.n31 VDD2.n30 9.3005
R1154 VDD2.n32 VDD2.n1 9.3005
R1155 VDD2.n62 VDD2.n61 8.92171
R1156 VDD2.n20 VDD2.n19 8.92171
R1157 VDD2.n58 VDD2.n52 8.14595
R1158 VDD2.n16 VDD2.n10 8.14595
R1159 VDD2.n57 VDD2.n54 7.3702
R1160 VDD2.n15 VDD2.n12 7.3702
R1161 VDD2.n58 VDD2.n57 5.81868
R1162 VDD2.n16 VDD2.n15 5.81868
R1163 VDD2.n61 VDD2.n52 5.04292
R1164 VDD2.n19 VDD2.n10 5.04292
R1165 VDD2.n62 VDD2.n50 4.26717
R1166 VDD2.n20 VDD2.n8 4.26717
R1167 VDD2.n66 VDD2.n65 3.49141
R1168 VDD2.n24 VDD2.n23 3.49141
R1169 VDD2.n69 VDD2.n48 2.71565
R1170 VDD2.n27 VDD2.n6 2.71565
R1171 VDD2.n56 VDD2.n55 2.4129
R1172 VDD2.n14 VDD2.n13 2.4129
R1173 VDD2.n70 VDD2.n46 1.93989
R1174 VDD2.n28 VDD2.n4 1.93989
R1175 VDD2.n81 VDD2.n41 1.16414
R1176 VDD2.n74 VDD2.n73 1.16414
R1177 VDD2.n33 VDD2.n31 1.16414
R1178 VDD2.n40 VDD2.n0 1.16414
R1179 VDD2 VDD2.n82 0.49619
R1180 VDD2.n79 VDD2.n78 0.388379
R1181 VDD2.n45 VDD2.n43 0.388379
R1182 VDD2.n32 VDD2.n2 0.388379
R1183 VDD2.n38 VDD2.n37 0.388379
R1184 VDD2.n80 VDD2.n42 0.155672
R1185 VDD2.n72 VDD2.n42 0.155672
R1186 VDD2.n72 VDD2.n71 0.155672
R1187 VDD2.n71 VDD2.n47 0.155672
R1188 VDD2.n64 VDD2.n47 0.155672
R1189 VDD2.n64 VDD2.n63 0.155672
R1190 VDD2.n63 VDD2.n51 0.155672
R1191 VDD2.n56 VDD2.n51 0.155672
R1192 VDD2.n14 VDD2.n9 0.155672
R1193 VDD2.n21 VDD2.n9 0.155672
R1194 VDD2.n22 VDD2.n21 0.155672
R1195 VDD2.n22 VDD2.n5 0.155672
R1196 VDD2.n29 VDD2.n5 0.155672
R1197 VDD2.n30 VDD2.n29 0.155672
R1198 VDD2.n30 VDD2.n1 0.155672
R1199 VDD2.n39 VDD2.n1 0.155672
C0 VDD2 w_n1782_n2550# 1.40562f
C1 B w_n1782_n2550# 6.68967f
C2 VN w_n1782_n2550# 2.31364f
C3 VTAIL w_n1782_n2550# 2.17587f
C4 VP VDD1 1.92188f
C5 VDD2 VDD1 0.568077f
C6 VDD2 VP 0.29492f
C7 B VDD1 1.26439f
C8 B VP 1.21615f
C9 VDD2 B 1.28651f
C10 VN VDD1 0.147709f
C11 VTAIL VDD1 3.85492f
C12 VN VP 4.27847f
C13 VTAIL VP 1.57267f
C14 VDD2 VN 1.77685f
C15 VDD2 VTAIL 3.89959f
C16 B VN 0.849765f
C17 B VTAIL 2.41068f
C18 VDD1 w_n1782_n2550# 1.39054f
C19 VN VTAIL 1.55838f
C20 VP w_n1782_n2550# 2.5387f
C21 VDD2 VSUBS 0.659124f
C22 VDD1 VSUBS 2.271446f
C23 VTAIL VSUBS 0.723651f
C24 VN VSUBS 5.19744f
C25 VP VSUBS 1.252447f
C26 B VSUBS 2.881903f
C27 w_n1782_n2550# VSUBS 56.389603f
C28 VDD2.n0 VSUBS 0.01465f
C29 VDD2.n1 VSUBS 0.014093f
C30 VDD2.n2 VSUBS 0.007796f
C31 VDD2.n3 VSUBS 0.0179f
C32 VDD2.n4 VSUBS 0.008019f
C33 VDD2.n5 VSUBS 0.014093f
C34 VDD2.n6 VSUBS 0.007573f
C35 VDD2.n7 VSUBS 0.0179f
C36 VDD2.n8 VSUBS 0.008019f
C37 VDD2.n9 VSUBS 0.014093f
C38 VDD2.n10 VSUBS 0.007573f
C39 VDD2.n11 VSUBS 0.013425f
C40 VDD2.n12 VSUBS 0.013465f
C41 VDD2.t0 VSUBS 0.038439f
C42 VDD2.n13 VSUBS 0.084981f
C43 VDD2.n14 VSUBS 0.439778f
C44 VDD2.n15 VSUBS 0.007573f
C45 VDD2.n16 VSUBS 0.008019f
C46 VDD2.n17 VSUBS 0.0179f
C47 VDD2.n18 VSUBS 0.0179f
C48 VDD2.n19 VSUBS 0.008019f
C49 VDD2.n20 VSUBS 0.007573f
C50 VDD2.n21 VSUBS 0.014093f
C51 VDD2.n22 VSUBS 0.014093f
C52 VDD2.n23 VSUBS 0.007573f
C53 VDD2.n24 VSUBS 0.008019f
C54 VDD2.n25 VSUBS 0.0179f
C55 VDD2.n26 VSUBS 0.0179f
C56 VDD2.n27 VSUBS 0.008019f
C57 VDD2.n28 VSUBS 0.007573f
C58 VDD2.n29 VSUBS 0.014093f
C59 VDD2.n30 VSUBS 0.014093f
C60 VDD2.n31 VSUBS 0.007573f
C61 VDD2.n32 VSUBS 0.007573f
C62 VDD2.n33 VSUBS 0.008019f
C63 VDD2.n34 VSUBS 0.0179f
C64 VDD2.n35 VSUBS 0.0179f
C65 VDD2.n36 VSUBS 0.040488f
C66 VDD2.n37 VSUBS 0.007796f
C67 VDD2.n38 VSUBS 0.007573f
C68 VDD2.n39 VSUBS 0.034694f
C69 VDD2.n40 VSUBS 0.297621f
C70 VDD2.n41 VSUBS 0.01465f
C71 VDD2.n42 VSUBS 0.014093f
C72 VDD2.n43 VSUBS 0.007796f
C73 VDD2.n44 VSUBS 0.0179f
C74 VDD2.n45 VSUBS 0.007573f
C75 VDD2.n46 VSUBS 0.008019f
C76 VDD2.n47 VSUBS 0.014093f
C77 VDD2.n48 VSUBS 0.007573f
C78 VDD2.n49 VSUBS 0.0179f
C79 VDD2.n50 VSUBS 0.008019f
C80 VDD2.n51 VSUBS 0.014093f
C81 VDD2.n52 VSUBS 0.007573f
C82 VDD2.n53 VSUBS 0.013425f
C83 VDD2.n54 VSUBS 0.013465f
C84 VDD2.t1 VSUBS 0.038439f
C85 VDD2.n55 VSUBS 0.084981f
C86 VDD2.n56 VSUBS 0.439778f
C87 VDD2.n57 VSUBS 0.007573f
C88 VDD2.n58 VSUBS 0.008019f
C89 VDD2.n59 VSUBS 0.0179f
C90 VDD2.n60 VSUBS 0.0179f
C91 VDD2.n61 VSUBS 0.008019f
C92 VDD2.n62 VSUBS 0.007573f
C93 VDD2.n63 VSUBS 0.014093f
C94 VDD2.n64 VSUBS 0.014093f
C95 VDD2.n65 VSUBS 0.007573f
C96 VDD2.n66 VSUBS 0.008019f
C97 VDD2.n67 VSUBS 0.0179f
C98 VDD2.n68 VSUBS 0.0179f
C99 VDD2.n69 VSUBS 0.008019f
C100 VDD2.n70 VSUBS 0.007573f
C101 VDD2.n71 VSUBS 0.014093f
C102 VDD2.n72 VSUBS 0.014093f
C103 VDD2.n73 VSUBS 0.007573f
C104 VDD2.n74 VSUBS 0.008019f
C105 VDD2.n75 VSUBS 0.0179f
C106 VDD2.n76 VSUBS 0.0179f
C107 VDD2.n77 VSUBS 0.040488f
C108 VDD2.n78 VSUBS 0.007796f
C109 VDD2.n79 VSUBS 0.007573f
C110 VDD2.n80 VSUBS 0.034694f
C111 VDD2.n81 VSUBS 0.030014f
C112 VDD2.n82 VSUBS 1.38641f
C113 VN.t1 VSUBS 1.48443f
C114 VN.t0 VSUBS 1.81909f
C115 VDD1.n0 VSUBS 0.014457f
C116 VDD1.n1 VSUBS 0.013908f
C117 VDD1.n2 VSUBS 0.007693f
C118 VDD1.n3 VSUBS 0.017664f
C119 VDD1.n4 VSUBS 0.007473f
C120 VDD1.n5 VSUBS 0.007913f
C121 VDD1.n6 VSUBS 0.013908f
C122 VDD1.n7 VSUBS 0.007473f
C123 VDD1.n8 VSUBS 0.017664f
C124 VDD1.n9 VSUBS 0.007913f
C125 VDD1.n10 VSUBS 0.013908f
C126 VDD1.n11 VSUBS 0.007473f
C127 VDD1.n12 VSUBS 0.013248f
C128 VDD1.n13 VSUBS 0.013288f
C129 VDD1.t1 VSUBS 0.037932f
C130 VDD1.n14 VSUBS 0.083862f
C131 VDD1.n15 VSUBS 0.433986f
C132 VDD1.n16 VSUBS 0.007473f
C133 VDD1.n17 VSUBS 0.007913f
C134 VDD1.n18 VSUBS 0.017664f
C135 VDD1.n19 VSUBS 0.017664f
C136 VDD1.n20 VSUBS 0.007913f
C137 VDD1.n21 VSUBS 0.007473f
C138 VDD1.n22 VSUBS 0.013908f
C139 VDD1.n23 VSUBS 0.013908f
C140 VDD1.n24 VSUBS 0.007473f
C141 VDD1.n25 VSUBS 0.007913f
C142 VDD1.n26 VSUBS 0.017664f
C143 VDD1.n27 VSUBS 0.017664f
C144 VDD1.n28 VSUBS 0.007913f
C145 VDD1.n29 VSUBS 0.007473f
C146 VDD1.n30 VSUBS 0.013908f
C147 VDD1.n31 VSUBS 0.013908f
C148 VDD1.n32 VSUBS 0.007473f
C149 VDD1.n33 VSUBS 0.007913f
C150 VDD1.n34 VSUBS 0.017664f
C151 VDD1.n35 VSUBS 0.017664f
C152 VDD1.n36 VSUBS 0.039955f
C153 VDD1.n37 VSUBS 0.007693f
C154 VDD1.n38 VSUBS 0.007473f
C155 VDD1.n39 VSUBS 0.034237f
C156 VDD1.n40 VSUBS 0.030102f
C157 VDD1.n41 VSUBS 0.014457f
C158 VDD1.n42 VSUBS 0.013908f
C159 VDD1.n43 VSUBS 0.007693f
C160 VDD1.n44 VSUBS 0.017664f
C161 VDD1.n45 VSUBS 0.007913f
C162 VDD1.n46 VSUBS 0.013908f
C163 VDD1.n47 VSUBS 0.007473f
C164 VDD1.n48 VSUBS 0.017664f
C165 VDD1.n49 VSUBS 0.007913f
C166 VDD1.n50 VSUBS 0.013908f
C167 VDD1.n51 VSUBS 0.007473f
C168 VDD1.n52 VSUBS 0.013248f
C169 VDD1.n53 VSUBS 0.013288f
C170 VDD1.t0 VSUBS 0.037932f
C171 VDD1.n54 VSUBS 0.083862f
C172 VDD1.n55 VSUBS 0.433986f
C173 VDD1.n56 VSUBS 0.007473f
C174 VDD1.n57 VSUBS 0.007913f
C175 VDD1.n58 VSUBS 0.017664f
C176 VDD1.n59 VSUBS 0.017664f
C177 VDD1.n60 VSUBS 0.007913f
C178 VDD1.n61 VSUBS 0.007473f
C179 VDD1.n62 VSUBS 0.013908f
C180 VDD1.n63 VSUBS 0.013908f
C181 VDD1.n64 VSUBS 0.007473f
C182 VDD1.n65 VSUBS 0.007913f
C183 VDD1.n66 VSUBS 0.017664f
C184 VDD1.n67 VSUBS 0.017664f
C185 VDD1.n68 VSUBS 0.007913f
C186 VDD1.n69 VSUBS 0.007473f
C187 VDD1.n70 VSUBS 0.013908f
C188 VDD1.n71 VSUBS 0.013908f
C189 VDD1.n72 VSUBS 0.007473f
C190 VDD1.n73 VSUBS 0.007473f
C191 VDD1.n74 VSUBS 0.007913f
C192 VDD1.n75 VSUBS 0.017664f
C193 VDD1.n76 VSUBS 0.017664f
C194 VDD1.n77 VSUBS 0.039955f
C195 VDD1.n78 VSUBS 0.007693f
C196 VDD1.n79 VSUBS 0.007473f
C197 VDD1.n80 VSUBS 0.034237f
C198 VDD1.n81 VSUBS 0.314499f
C199 VTAIL.n0 VSUBS 0.025563f
C200 VTAIL.n1 VSUBS 0.024592f
C201 VTAIL.n2 VSUBS 0.013603f
C202 VTAIL.n3 VSUBS 0.031235f
C203 VTAIL.n4 VSUBS 0.013992f
C204 VTAIL.n5 VSUBS 0.024592f
C205 VTAIL.n6 VSUBS 0.013215f
C206 VTAIL.n7 VSUBS 0.031235f
C207 VTAIL.n8 VSUBS 0.013992f
C208 VTAIL.n9 VSUBS 0.024592f
C209 VTAIL.n10 VSUBS 0.013215f
C210 VTAIL.n11 VSUBS 0.023426f
C211 VTAIL.n12 VSUBS 0.023496f
C212 VTAIL.t2 VSUBS 0.067073f
C213 VTAIL.n13 VSUBS 0.148286f
C214 VTAIL.n14 VSUBS 0.767382f
C215 VTAIL.n15 VSUBS 0.013215f
C216 VTAIL.n16 VSUBS 0.013992f
C217 VTAIL.n17 VSUBS 0.031235f
C218 VTAIL.n18 VSUBS 0.031235f
C219 VTAIL.n19 VSUBS 0.013992f
C220 VTAIL.n20 VSUBS 0.013215f
C221 VTAIL.n21 VSUBS 0.024592f
C222 VTAIL.n22 VSUBS 0.024592f
C223 VTAIL.n23 VSUBS 0.013215f
C224 VTAIL.n24 VSUBS 0.013992f
C225 VTAIL.n25 VSUBS 0.031235f
C226 VTAIL.n26 VSUBS 0.031235f
C227 VTAIL.n27 VSUBS 0.013992f
C228 VTAIL.n28 VSUBS 0.013215f
C229 VTAIL.n29 VSUBS 0.024592f
C230 VTAIL.n30 VSUBS 0.024592f
C231 VTAIL.n31 VSUBS 0.013215f
C232 VTAIL.n32 VSUBS 0.013215f
C233 VTAIL.n33 VSUBS 0.013992f
C234 VTAIL.n34 VSUBS 0.031235f
C235 VTAIL.n35 VSUBS 0.031235f
C236 VTAIL.n36 VSUBS 0.070649f
C237 VTAIL.n37 VSUBS 0.013603f
C238 VTAIL.n38 VSUBS 0.013215f
C239 VTAIL.n39 VSUBS 0.060539f
C240 VTAIL.n40 VSUBS 0.035419f
C241 VTAIL.n41 VSUBS 1.25134f
C242 VTAIL.n42 VSUBS 0.025563f
C243 VTAIL.n43 VSUBS 0.024592f
C244 VTAIL.n44 VSUBS 0.013603f
C245 VTAIL.n45 VSUBS 0.031235f
C246 VTAIL.n46 VSUBS 0.013215f
C247 VTAIL.n47 VSUBS 0.013992f
C248 VTAIL.n48 VSUBS 0.024592f
C249 VTAIL.n49 VSUBS 0.013215f
C250 VTAIL.n50 VSUBS 0.031235f
C251 VTAIL.n51 VSUBS 0.013992f
C252 VTAIL.n52 VSUBS 0.024592f
C253 VTAIL.n53 VSUBS 0.013215f
C254 VTAIL.n54 VSUBS 0.023426f
C255 VTAIL.n55 VSUBS 0.023496f
C256 VTAIL.t0 VSUBS 0.067073f
C257 VTAIL.n56 VSUBS 0.148286f
C258 VTAIL.n57 VSUBS 0.767382f
C259 VTAIL.n58 VSUBS 0.013215f
C260 VTAIL.n59 VSUBS 0.013992f
C261 VTAIL.n60 VSUBS 0.031235f
C262 VTAIL.n61 VSUBS 0.031235f
C263 VTAIL.n62 VSUBS 0.013992f
C264 VTAIL.n63 VSUBS 0.013215f
C265 VTAIL.n64 VSUBS 0.024592f
C266 VTAIL.n65 VSUBS 0.024592f
C267 VTAIL.n66 VSUBS 0.013215f
C268 VTAIL.n67 VSUBS 0.013992f
C269 VTAIL.n68 VSUBS 0.031235f
C270 VTAIL.n69 VSUBS 0.031235f
C271 VTAIL.n70 VSUBS 0.013992f
C272 VTAIL.n71 VSUBS 0.013215f
C273 VTAIL.n72 VSUBS 0.024592f
C274 VTAIL.n73 VSUBS 0.024592f
C275 VTAIL.n74 VSUBS 0.013215f
C276 VTAIL.n75 VSUBS 0.013992f
C277 VTAIL.n76 VSUBS 0.031235f
C278 VTAIL.n77 VSUBS 0.031235f
C279 VTAIL.n78 VSUBS 0.070649f
C280 VTAIL.n79 VSUBS 0.013603f
C281 VTAIL.n80 VSUBS 0.013215f
C282 VTAIL.n81 VSUBS 0.060539f
C283 VTAIL.n82 VSUBS 0.035419f
C284 VTAIL.n83 VSUBS 1.2814f
C285 VTAIL.n84 VSUBS 0.025563f
C286 VTAIL.n85 VSUBS 0.024592f
C287 VTAIL.n86 VSUBS 0.013603f
C288 VTAIL.n87 VSUBS 0.031235f
C289 VTAIL.n88 VSUBS 0.013215f
C290 VTAIL.n89 VSUBS 0.013992f
C291 VTAIL.n90 VSUBS 0.024592f
C292 VTAIL.n91 VSUBS 0.013215f
C293 VTAIL.n92 VSUBS 0.031235f
C294 VTAIL.n93 VSUBS 0.013992f
C295 VTAIL.n94 VSUBS 0.024592f
C296 VTAIL.n95 VSUBS 0.013215f
C297 VTAIL.n96 VSUBS 0.023426f
C298 VTAIL.n97 VSUBS 0.023496f
C299 VTAIL.t3 VSUBS 0.067073f
C300 VTAIL.n98 VSUBS 0.148286f
C301 VTAIL.n99 VSUBS 0.767382f
C302 VTAIL.n100 VSUBS 0.013215f
C303 VTAIL.n101 VSUBS 0.013992f
C304 VTAIL.n102 VSUBS 0.031235f
C305 VTAIL.n103 VSUBS 0.031235f
C306 VTAIL.n104 VSUBS 0.013992f
C307 VTAIL.n105 VSUBS 0.013215f
C308 VTAIL.n106 VSUBS 0.024592f
C309 VTAIL.n107 VSUBS 0.024592f
C310 VTAIL.n108 VSUBS 0.013215f
C311 VTAIL.n109 VSUBS 0.013992f
C312 VTAIL.n110 VSUBS 0.031235f
C313 VTAIL.n111 VSUBS 0.031235f
C314 VTAIL.n112 VSUBS 0.013992f
C315 VTAIL.n113 VSUBS 0.013215f
C316 VTAIL.n114 VSUBS 0.024592f
C317 VTAIL.n115 VSUBS 0.024592f
C318 VTAIL.n116 VSUBS 0.013215f
C319 VTAIL.n117 VSUBS 0.013992f
C320 VTAIL.n118 VSUBS 0.031235f
C321 VTAIL.n119 VSUBS 0.031235f
C322 VTAIL.n120 VSUBS 0.070649f
C323 VTAIL.n121 VSUBS 0.013603f
C324 VTAIL.n122 VSUBS 0.013215f
C325 VTAIL.n123 VSUBS 0.060539f
C326 VTAIL.n124 VSUBS 0.035419f
C327 VTAIL.n125 VSUBS 1.14273f
C328 VTAIL.n126 VSUBS 0.025563f
C329 VTAIL.n127 VSUBS 0.024592f
C330 VTAIL.n128 VSUBS 0.013603f
C331 VTAIL.n129 VSUBS 0.031235f
C332 VTAIL.n130 VSUBS 0.013992f
C333 VTAIL.n131 VSUBS 0.024592f
C334 VTAIL.n132 VSUBS 0.013215f
C335 VTAIL.n133 VSUBS 0.031235f
C336 VTAIL.n134 VSUBS 0.013992f
C337 VTAIL.n135 VSUBS 0.024592f
C338 VTAIL.n136 VSUBS 0.013215f
C339 VTAIL.n137 VSUBS 0.023426f
C340 VTAIL.n138 VSUBS 0.023496f
C341 VTAIL.t1 VSUBS 0.067073f
C342 VTAIL.n139 VSUBS 0.148286f
C343 VTAIL.n140 VSUBS 0.767382f
C344 VTAIL.n141 VSUBS 0.013215f
C345 VTAIL.n142 VSUBS 0.013992f
C346 VTAIL.n143 VSUBS 0.031235f
C347 VTAIL.n144 VSUBS 0.031235f
C348 VTAIL.n145 VSUBS 0.013992f
C349 VTAIL.n146 VSUBS 0.013215f
C350 VTAIL.n147 VSUBS 0.024592f
C351 VTAIL.n148 VSUBS 0.024592f
C352 VTAIL.n149 VSUBS 0.013215f
C353 VTAIL.n150 VSUBS 0.013992f
C354 VTAIL.n151 VSUBS 0.031235f
C355 VTAIL.n152 VSUBS 0.031235f
C356 VTAIL.n153 VSUBS 0.013992f
C357 VTAIL.n154 VSUBS 0.013215f
C358 VTAIL.n155 VSUBS 0.024592f
C359 VTAIL.n156 VSUBS 0.024592f
C360 VTAIL.n157 VSUBS 0.013215f
C361 VTAIL.n158 VSUBS 0.013215f
C362 VTAIL.n159 VSUBS 0.013992f
C363 VTAIL.n160 VSUBS 0.031235f
C364 VTAIL.n161 VSUBS 0.031235f
C365 VTAIL.n162 VSUBS 0.070649f
C366 VTAIL.n163 VSUBS 0.013603f
C367 VTAIL.n164 VSUBS 0.013215f
C368 VTAIL.n165 VSUBS 0.060539f
C369 VTAIL.n166 VSUBS 0.035419f
C370 VTAIL.n167 VSUBS 1.06622f
C371 VP.t0 VSUBS 1.8837f
C372 VP.t1 VSUBS 1.54016f
C373 VP.n0 VSUBS 3.32377f
C374 B.n0 VSUBS 0.004723f
C375 B.n1 VSUBS 0.004723f
C376 B.n2 VSUBS 0.007469f
C377 B.n3 VSUBS 0.007469f
C378 B.n4 VSUBS 0.007469f
C379 B.n5 VSUBS 0.007469f
C380 B.n6 VSUBS 0.007469f
C381 B.n7 VSUBS 0.007469f
C382 B.n8 VSUBS 0.007469f
C383 B.n9 VSUBS 0.007469f
C384 B.n10 VSUBS 0.007469f
C385 B.n11 VSUBS 0.007469f
C386 B.n12 VSUBS 0.0177f
C387 B.n13 VSUBS 0.007469f
C388 B.n14 VSUBS 0.007469f
C389 B.n15 VSUBS 0.007469f
C390 B.n16 VSUBS 0.007469f
C391 B.n17 VSUBS 0.007469f
C392 B.n18 VSUBS 0.007469f
C393 B.n19 VSUBS 0.007469f
C394 B.n20 VSUBS 0.007469f
C395 B.n21 VSUBS 0.007469f
C396 B.n22 VSUBS 0.007469f
C397 B.n23 VSUBS 0.007469f
C398 B.n24 VSUBS 0.007469f
C399 B.n25 VSUBS 0.007469f
C400 B.n26 VSUBS 0.007469f
C401 B.n27 VSUBS 0.007469f
C402 B.t2 VSUBS 0.133078f
C403 B.t1 VSUBS 0.154807f
C404 B.t0 VSUBS 0.651536f
C405 B.n28 VSUBS 0.259378f
C406 B.n29 VSUBS 0.199031f
C407 B.n30 VSUBS 0.007469f
C408 B.n31 VSUBS 0.007469f
C409 B.n32 VSUBS 0.007469f
C410 B.n33 VSUBS 0.007469f
C411 B.t8 VSUBS 0.133081f
C412 B.t7 VSUBS 0.154809f
C413 B.t6 VSUBS 0.651536f
C414 B.n34 VSUBS 0.259376f
C415 B.n35 VSUBS 0.199029f
C416 B.n36 VSUBS 0.007469f
C417 B.n37 VSUBS 0.007469f
C418 B.n38 VSUBS 0.007469f
C419 B.n39 VSUBS 0.007469f
C420 B.n40 VSUBS 0.007469f
C421 B.n41 VSUBS 0.007469f
C422 B.n42 VSUBS 0.007469f
C423 B.n43 VSUBS 0.007469f
C424 B.n44 VSUBS 0.007469f
C425 B.n45 VSUBS 0.007469f
C426 B.n46 VSUBS 0.007469f
C427 B.n47 VSUBS 0.007469f
C428 B.n48 VSUBS 0.007469f
C429 B.n49 VSUBS 0.007469f
C430 B.n50 VSUBS 0.016791f
C431 B.n51 VSUBS 0.007469f
C432 B.n52 VSUBS 0.007469f
C433 B.n53 VSUBS 0.007469f
C434 B.n54 VSUBS 0.007469f
C435 B.n55 VSUBS 0.007469f
C436 B.n56 VSUBS 0.007469f
C437 B.n57 VSUBS 0.007469f
C438 B.n58 VSUBS 0.007469f
C439 B.n59 VSUBS 0.007469f
C440 B.n60 VSUBS 0.007469f
C441 B.n61 VSUBS 0.007469f
C442 B.n62 VSUBS 0.007469f
C443 B.n63 VSUBS 0.007469f
C444 B.n64 VSUBS 0.007469f
C445 B.n65 VSUBS 0.007469f
C446 B.n66 VSUBS 0.007469f
C447 B.n67 VSUBS 0.007469f
C448 B.n68 VSUBS 0.007469f
C449 B.n69 VSUBS 0.007469f
C450 B.n70 VSUBS 0.007469f
C451 B.n71 VSUBS 0.0177f
C452 B.n72 VSUBS 0.007469f
C453 B.n73 VSUBS 0.007469f
C454 B.n74 VSUBS 0.007469f
C455 B.n75 VSUBS 0.007469f
C456 B.n76 VSUBS 0.007469f
C457 B.n77 VSUBS 0.007469f
C458 B.n78 VSUBS 0.007469f
C459 B.n79 VSUBS 0.007469f
C460 B.n80 VSUBS 0.007469f
C461 B.n81 VSUBS 0.007469f
C462 B.n82 VSUBS 0.007469f
C463 B.n83 VSUBS 0.007469f
C464 B.n84 VSUBS 0.007469f
C465 B.n85 VSUBS 0.007469f
C466 B.t10 VSUBS 0.133081f
C467 B.t11 VSUBS 0.154809f
C468 B.t9 VSUBS 0.651536f
C469 B.n86 VSUBS 0.259376f
C470 B.n87 VSUBS 0.199029f
C471 B.n88 VSUBS 0.017305f
C472 B.n89 VSUBS 0.007469f
C473 B.n90 VSUBS 0.007469f
C474 B.n91 VSUBS 0.007469f
C475 B.n92 VSUBS 0.007469f
C476 B.n93 VSUBS 0.007469f
C477 B.t4 VSUBS 0.133078f
C478 B.t5 VSUBS 0.154807f
C479 B.t3 VSUBS 0.651536f
C480 B.n94 VSUBS 0.259378f
C481 B.n95 VSUBS 0.199031f
C482 B.n96 VSUBS 0.007469f
C483 B.n97 VSUBS 0.007469f
C484 B.n98 VSUBS 0.007469f
C485 B.n99 VSUBS 0.007469f
C486 B.n100 VSUBS 0.007469f
C487 B.n101 VSUBS 0.007469f
C488 B.n102 VSUBS 0.007469f
C489 B.n103 VSUBS 0.007469f
C490 B.n104 VSUBS 0.007469f
C491 B.n105 VSUBS 0.007469f
C492 B.n106 VSUBS 0.007469f
C493 B.n107 VSUBS 0.007469f
C494 B.n108 VSUBS 0.007469f
C495 B.n109 VSUBS 0.007469f
C496 B.n110 VSUBS 0.016569f
C497 B.n111 VSUBS 0.007469f
C498 B.n112 VSUBS 0.007469f
C499 B.n113 VSUBS 0.007469f
C500 B.n114 VSUBS 0.007469f
C501 B.n115 VSUBS 0.007469f
C502 B.n116 VSUBS 0.007469f
C503 B.n117 VSUBS 0.007469f
C504 B.n118 VSUBS 0.007469f
C505 B.n119 VSUBS 0.007469f
C506 B.n120 VSUBS 0.007469f
C507 B.n121 VSUBS 0.007469f
C508 B.n122 VSUBS 0.007469f
C509 B.n123 VSUBS 0.007469f
C510 B.n124 VSUBS 0.007469f
C511 B.n125 VSUBS 0.007469f
C512 B.n126 VSUBS 0.007469f
C513 B.n127 VSUBS 0.007469f
C514 B.n128 VSUBS 0.007469f
C515 B.n129 VSUBS 0.007469f
C516 B.n130 VSUBS 0.007469f
C517 B.n131 VSUBS 0.007469f
C518 B.n132 VSUBS 0.007469f
C519 B.n133 VSUBS 0.007469f
C520 B.n134 VSUBS 0.007469f
C521 B.n135 VSUBS 0.007469f
C522 B.n136 VSUBS 0.007469f
C523 B.n137 VSUBS 0.007469f
C524 B.n138 VSUBS 0.007469f
C525 B.n139 VSUBS 0.007469f
C526 B.n140 VSUBS 0.007469f
C527 B.n141 VSUBS 0.007469f
C528 B.n142 VSUBS 0.007469f
C529 B.n143 VSUBS 0.007469f
C530 B.n144 VSUBS 0.007469f
C531 B.n145 VSUBS 0.007469f
C532 B.n146 VSUBS 0.007469f
C533 B.n147 VSUBS 0.016569f
C534 B.n148 VSUBS 0.0177f
C535 B.n149 VSUBS 0.0177f
C536 B.n150 VSUBS 0.007469f
C537 B.n151 VSUBS 0.007469f
C538 B.n152 VSUBS 0.007469f
C539 B.n153 VSUBS 0.007469f
C540 B.n154 VSUBS 0.007469f
C541 B.n155 VSUBS 0.007469f
C542 B.n156 VSUBS 0.007469f
C543 B.n157 VSUBS 0.007469f
C544 B.n158 VSUBS 0.007469f
C545 B.n159 VSUBS 0.007469f
C546 B.n160 VSUBS 0.007469f
C547 B.n161 VSUBS 0.007469f
C548 B.n162 VSUBS 0.007469f
C549 B.n163 VSUBS 0.007469f
C550 B.n164 VSUBS 0.007469f
C551 B.n165 VSUBS 0.007469f
C552 B.n166 VSUBS 0.007469f
C553 B.n167 VSUBS 0.007469f
C554 B.n168 VSUBS 0.007469f
C555 B.n169 VSUBS 0.007469f
C556 B.n170 VSUBS 0.007469f
C557 B.n171 VSUBS 0.007469f
C558 B.n172 VSUBS 0.007469f
C559 B.n173 VSUBS 0.007469f
C560 B.n174 VSUBS 0.007469f
C561 B.n175 VSUBS 0.007469f
C562 B.n176 VSUBS 0.007469f
C563 B.n177 VSUBS 0.007469f
C564 B.n178 VSUBS 0.007469f
C565 B.n179 VSUBS 0.007469f
C566 B.n180 VSUBS 0.007469f
C567 B.n181 VSUBS 0.007469f
C568 B.n182 VSUBS 0.007469f
C569 B.n183 VSUBS 0.007469f
C570 B.n184 VSUBS 0.007469f
C571 B.n185 VSUBS 0.007469f
C572 B.n186 VSUBS 0.007469f
C573 B.n187 VSUBS 0.007469f
C574 B.n188 VSUBS 0.007469f
C575 B.n189 VSUBS 0.007469f
C576 B.n190 VSUBS 0.007469f
C577 B.n191 VSUBS 0.007469f
C578 B.n192 VSUBS 0.005162f
C579 B.n193 VSUBS 0.017305f
C580 B.n194 VSUBS 0.006041f
C581 B.n195 VSUBS 0.007469f
C582 B.n196 VSUBS 0.007469f
C583 B.n197 VSUBS 0.007469f
C584 B.n198 VSUBS 0.007469f
C585 B.n199 VSUBS 0.007469f
C586 B.n200 VSUBS 0.007469f
C587 B.n201 VSUBS 0.007469f
C588 B.n202 VSUBS 0.007469f
C589 B.n203 VSUBS 0.007469f
C590 B.n204 VSUBS 0.007469f
C591 B.n205 VSUBS 0.007469f
C592 B.n206 VSUBS 0.006041f
C593 B.n207 VSUBS 0.007469f
C594 B.n208 VSUBS 0.007469f
C595 B.n209 VSUBS 0.005162f
C596 B.n210 VSUBS 0.007469f
C597 B.n211 VSUBS 0.007469f
C598 B.n212 VSUBS 0.007469f
C599 B.n213 VSUBS 0.007469f
C600 B.n214 VSUBS 0.007469f
C601 B.n215 VSUBS 0.007469f
C602 B.n216 VSUBS 0.007469f
C603 B.n217 VSUBS 0.007469f
C604 B.n218 VSUBS 0.007469f
C605 B.n219 VSUBS 0.007469f
C606 B.n220 VSUBS 0.007469f
C607 B.n221 VSUBS 0.007469f
C608 B.n222 VSUBS 0.007469f
C609 B.n223 VSUBS 0.007469f
C610 B.n224 VSUBS 0.007469f
C611 B.n225 VSUBS 0.007469f
C612 B.n226 VSUBS 0.007469f
C613 B.n227 VSUBS 0.007469f
C614 B.n228 VSUBS 0.007469f
C615 B.n229 VSUBS 0.007469f
C616 B.n230 VSUBS 0.007469f
C617 B.n231 VSUBS 0.007469f
C618 B.n232 VSUBS 0.007469f
C619 B.n233 VSUBS 0.007469f
C620 B.n234 VSUBS 0.007469f
C621 B.n235 VSUBS 0.007469f
C622 B.n236 VSUBS 0.007469f
C623 B.n237 VSUBS 0.007469f
C624 B.n238 VSUBS 0.007469f
C625 B.n239 VSUBS 0.007469f
C626 B.n240 VSUBS 0.007469f
C627 B.n241 VSUBS 0.007469f
C628 B.n242 VSUBS 0.007469f
C629 B.n243 VSUBS 0.007469f
C630 B.n244 VSUBS 0.007469f
C631 B.n245 VSUBS 0.007469f
C632 B.n246 VSUBS 0.007469f
C633 B.n247 VSUBS 0.007469f
C634 B.n248 VSUBS 0.007469f
C635 B.n249 VSUBS 0.007469f
C636 B.n250 VSUBS 0.007469f
C637 B.n251 VSUBS 0.007469f
C638 B.n252 VSUBS 0.0177f
C639 B.n253 VSUBS 0.016569f
C640 B.n254 VSUBS 0.016569f
C641 B.n255 VSUBS 0.007469f
C642 B.n256 VSUBS 0.007469f
C643 B.n257 VSUBS 0.007469f
C644 B.n258 VSUBS 0.007469f
C645 B.n259 VSUBS 0.007469f
C646 B.n260 VSUBS 0.007469f
C647 B.n261 VSUBS 0.007469f
C648 B.n262 VSUBS 0.007469f
C649 B.n263 VSUBS 0.007469f
C650 B.n264 VSUBS 0.007469f
C651 B.n265 VSUBS 0.007469f
C652 B.n266 VSUBS 0.007469f
C653 B.n267 VSUBS 0.007469f
C654 B.n268 VSUBS 0.007469f
C655 B.n269 VSUBS 0.007469f
C656 B.n270 VSUBS 0.007469f
C657 B.n271 VSUBS 0.007469f
C658 B.n272 VSUBS 0.007469f
C659 B.n273 VSUBS 0.007469f
C660 B.n274 VSUBS 0.007469f
C661 B.n275 VSUBS 0.007469f
C662 B.n276 VSUBS 0.007469f
C663 B.n277 VSUBS 0.007469f
C664 B.n278 VSUBS 0.007469f
C665 B.n279 VSUBS 0.007469f
C666 B.n280 VSUBS 0.007469f
C667 B.n281 VSUBS 0.007469f
C668 B.n282 VSUBS 0.007469f
C669 B.n283 VSUBS 0.007469f
C670 B.n284 VSUBS 0.007469f
C671 B.n285 VSUBS 0.007469f
C672 B.n286 VSUBS 0.007469f
C673 B.n287 VSUBS 0.007469f
C674 B.n288 VSUBS 0.007469f
C675 B.n289 VSUBS 0.007469f
C676 B.n290 VSUBS 0.007469f
C677 B.n291 VSUBS 0.007469f
C678 B.n292 VSUBS 0.007469f
C679 B.n293 VSUBS 0.007469f
C680 B.n294 VSUBS 0.007469f
C681 B.n295 VSUBS 0.007469f
C682 B.n296 VSUBS 0.007469f
C683 B.n297 VSUBS 0.007469f
C684 B.n298 VSUBS 0.007469f
C685 B.n299 VSUBS 0.007469f
C686 B.n300 VSUBS 0.007469f
C687 B.n301 VSUBS 0.007469f
C688 B.n302 VSUBS 0.007469f
C689 B.n303 VSUBS 0.007469f
C690 B.n304 VSUBS 0.007469f
C691 B.n305 VSUBS 0.007469f
C692 B.n306 VSUBS 0.007469f
C693 B.n307 VSUBS 0.007469f
C694 B.n308 VSUBS 0.007469f
C695 B.n309 VSUBS 0.007469f
C696 B.n310 VSUBS 0.007469f
C697 B.n311 VSUBS 0.007469f
C698 B.n312 VSUBS 0.007469f
C699 B.n313 VSUBS 0.017479f
C700 B.n314 VSUBS 0.016569f
C701 B.n315 VSUBS 0.0177f
C702 B.n316 VSUBS 0.007469f
C703 B.n317 VSUBS 0.007469f
C704 B.n318 VSUBS 0.007469f
C705 B.n319 VSUBS 0.007469f
C706 B.n320 VSUBS 0.007469f
C707 B.n321 VSUBS 0.007469f
C708 B.n322 VSUBS 0.007469f
C709 B.n323 VSUBS 0.007469f
C710 B.n324 VSUBS 0.007469f
C711 B.n325 VSUBS 0.007469f
C712 B.n326 VSUBS 0.007469f
C713 B.n327 VSUBS 0.007469f
C714 B.n328 VSUBS 0.007469f
C715 B.n329 VSUBS 0.007469f
C716 B.n330 VSUBS 0.007469f
C717 B.n331 VSUBS 0.007469f
C718 B.n332 VSUBS 0.007469f
C719 B.n333 VSUBS 0.007469f
C720 B.n334 VSUBS 0.007469f
C721 B.n335 VSUBS 0.007469f
C722 B.n336 VSUBS 0.007469f
C723 B.n337 VSUBS 0.007469f
C724 B.n338 VSUBS 0.007469f
C725 B.n339 VSUBS 0.007469f
C726 B.n340 VSUBS 0.007469f
C727 B.n341 VSUBS 0.007469f
C728 B.n342 VSUBS 0.007469f
C729 B.n343 VSUBS 0.007469f
C730 B.n344 VSUBS 0.007469f
C731 B.n345 VSUBS 0.007469f
C732 B.n346 VSUBS 0.007469f
C733 B.n347 VSUBS 0.007469f
C734 B.n348 VSUBS 0.007469f
C735 B.n349 VSUBS 0.007469f
C736 B.n350 VSUBS 0.007469f
C737 B.n351 VSUBS 0.007469f
C738 B.n352 VSUBS 0.007469f
C739 B.n353 VSUBS 0.007469f
C740 B.n354 VSUBS 0.007469f
C741 B.n355 VSUBS 0.007469f
C742 B.n356 VSUBS 0.007469f
C743 B.n357 VSUBS 0.007469f
C744 B.n358 VSUBS 0.007469f
C745 B.n359 VSUBS 0.005162f
C746 B.n360 VSUBS 0.017305f
C747 B.n361 VSUBS 0.006041f
C748 B.n362 VSUBS 0.007469f
C749 B.n363 VSUBS 0.007469f
C750 B.n364 VSUBS 0.007469f
C751 B.n365 VSUBS 0.007469f
C752 B.n366 VSUBS 0.007469f
C753 B.n367 VSUBS 0.007469f
C754 B.n368 VSUBS 0.007469f
C755 B.n369 VSUBS 0.007469f
C756 B.n370 VSUBS 0.007469f
C757 B.n371 VSUBS 0.007469f
C758 B.n372 VSUBS 0.007469f
C759 B.n373 VSUBS 0.006041f
C760 B.n374 VSUBS 0.017305f
C761 B.n375 VSUBS 0.005162f
C762 B.n376 VSUBS 0.007469f
C763 B.n377 VSUBS 0.007469f
C764 B.n378 VSUBS 0.007469f
C765 B.n379 VSUBS 0.007469f
C766 B.n380 VSUBS 0.007469f
C767 B.n381 VSUBS 0.007469f
C768 B.n382 VSUBS 0.007469f
C769 B.n383 VSUBS 0.007469f
C770 B.n384 VSUBS 0.007469f
C771 B.n385 VSUBS 0.007469f
C772 B.n386 VSUBS 0.007469f
C773 B.n387 VSUBS 0.007469f
C774 B.n388 VSUBS 0.007469f
C775 B.n389 VSUBS 0.007469f
C776 B.n390 VSUBS 0.007469f
C777 B.n391 VSUBS 0.007469f
C778 B.n392 VSUBS 0.007469f
C779 B.n393 VSUBS 0.007469f
C780 B.n394 VSUBS 0.007469f
C781 B.n395 VSUBS 0.007469f
C782 B.n396 VSUBS 0.007469f
C783 B.n397 VSUBS 0.007469f
C784 B.n398 VSUBS 0.007469f
C785 B.n399 VSUBS 0.007469f
C786 B.n400 VSUBS 0.007469f
C787 B.n401 VSUBS 0.007469f
C788 B.n402 VSUBS 0.007469f
C789 B.n403 VSUBS 0.007469f
C790 B.n404 VSUBS 0.007469f
C791 B.n405 VSUBS 0.007469f
C792 B.n406 VSUBS 0.007469f
C793 B.n407 VSUBS 0.007469f
C794 B.n408 VSUBS 0.007469f
C795 B.n409 VSUBS 0.007469f
C796 B.n410 VSUBS 0.007469f
C797 B.n411 VSUBS 0.007469f
C798 B.n412 VSUBS 0.007469f
C799 B.n413 VSUBS 0.007469f
C800 B.n414 VSUBS 0.007469f
C801 B.n415 VSUBS 0.007469f
C802 B.n416 VSUBS 0.007469f
C803 B.n417 VSUBS 0.007469f
C804 B.n418 VSUBS 0.007469f
C805 B.n419 VSUBS 0.0177f
C806 B.n420 VSUBS 0.016569f
C807 B.n421 VSUBS 0.016569f
C808 B.n422 VSUBS 0.007469f
C809 B.n423 VSUBS 0.007469f
C810 B.n424 VSUBS 0.007469f
C811 B.n425 VSUBS 0.007469f
C812 B.n426 VSUBS 0.007469f
C813 B.n427 VSUBS 0.007469f
C814 B.n428 VSUBS 0.007469f
C815 B.n429 VSUBS 0.007469f
C816 B.n430 VSUBS 0.007469f
C817 B.n431 VSUBS 0.007469f
C818 B.n432 VSUBS 0.007469f
C819 B.n433 VSUBS 0.007469f
C820 B.n434 VSUBS 0.007469f
C821 B.n435 VSUBS 0.007469f
C822 B.n436 VSUBS 0.007469f
C823 B.n437 VSUBS 0.007469f
C824 B.n438 VSUBS 0.007469f
C825 B.n439 VSUBS 0.007469f
C826 B.n440 VSUBS 0.007469f
C827 B.n441 VSUBS 0.007469f
C828 B.n442 VSUBS 0.007469f
C829 B.n443 VSUBS 0.007469f
C830 B.n444 VSUBS 0.007469f
C831 B.n445 VSUBS 0.007469f
C832 B.n446 VSUBS 0.007469f
C833 B.n447 VSUBS 0.007469f
C834 B.n448 VSUBS 0.007469f
C835 B.n449 VSUBS 0.007469f
C836 B.n450 VSUBS 0.007469f
C837 B.n451 VSUBS 0.016912f
.ends

