* NGSPICE file created from diff_pair_sample_1001.ext - technology: sky130A

.subckt diff_pair_sample_1001 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=3.73
X1 VDD1.t7 VP.t0 VTAIL.t9 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=3.73
X2 B.t8 B.t6 B.t7 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=3.73
X3 VDD2.t7 VN.t0 VTAIL.t2 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X4 VTAIL.t12 VN.t1 VDD2.t6 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X5 VTAIL.t4 VP.t1 VDD1.t6 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X6 VTAIL.t3 VP.t2 VDD1.t5 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=3.73
X7 B.t5 B.t3 B.t4 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=3.73
X8 VTAIL.t13 VN.t2 VDD2.t5 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=3.73
X9 VDD2.t4 VN.t3 VTAIL.t14 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=3.73
X10 VDD1.t4 VP.t3 VTAIL.t10 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X11 VTAIL.t15 VN.t4 VDD2.t3 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X12 VTAIL.t7 VP.t4 VDD1.t3 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X13 B.t2 B.t0 B.t1 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=0 ps=0 w=19.44 l=3.73
X14 VTAIL.t1 VN.t5 VDD2.t2 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=3.73
X15 VDD1.t2 VP.t5 VTAIL.t5 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=3.73
X16 VTAIL.t8 VP.t6 VDD1.t1 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=7.5816 pd=39.66 as=3.2076 ps=19.77 w=19.44 l=3.73
X17 VDD2.t1 VN.t6 VTAIL.t11 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=7.5816 ps=39.66 w=19.44 l=3.73
X18 VDD1.t0 VP.t7 VTAIL.t6 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
X19 VDD2.t0 VN.t7 VTAIL.t0 w_n5030_n4856# sky130_fd_pr__pfet_01v8 ad=3.2076 pd=19.77 as=3.2076 ps=19.77 w=19.44 l=3.73
R0 B.n210 B.t5 588.221
R1 B.n76 B.t7 588.221
R2 B.n216 B.t2 588.221
R3 B.n68 B.t10 588.221
R4 B.n798 B.n797 585
R5 B.n799 B.n108 585
R6 B.n801 B.n800 585
R7 B.n802 B.n107 585
R8 B.n804 B.n803 585
R9 B.n805 B.n106 585
R10 B.n807 B.n806 585
R11 B.n808 B.n105 585
R12 B.n810 B.n809 585
R13 B.n811 B.n104 585
R14 B.n813 B.n812 585
R15 B.n814 B.n103 585
R16 B.n816 B.n815 585
R17 B.n817 B.n102 585
R18 B.n819 B.n818 585
R19 B.n820 B.n101 585
R20 B.n822 B.n821 585
R21 B.n823 B.n100 585
R22 B.n825 B.n824 585
R23 B.n826 B.n99 585
R24 B.n828 B.n827 585
R25 B.n829 B.n98 585
R26 B.n831 B.n830 585
R27 B.n832 B.n97 585
R28 B.n834 B.n833 585
R29 B.n835 B.n96 585
R30 B.n837 B.n836 585
R31 B.n838 B.n95 585
R32 B.n840 B.n839 585
R33 B.n841 B.n94 585
R34 B.n843 B.n842 585
R35 B.n844 B.n93 585
R36 B.n846 B.n845 585
R37 B.n847 B.n92 585
R38 B.n849 B.n848 585
R39 B.n850 B.n91 585
R40 B.n852 B.n851 585
R41 B.n853 B.n90 585
R42 B.n855 B.n854 585
R43 B.n856 B.n89 585
R44 B.n858 B.n857 585
R45 B.n859 B.n88 585
R46 B.n861 B.n860 585
R47 B.n862 B.n87 585
R48 B.n864 B.n863 585
R49 B.n865 B.n86 585
R50 B.n867 B.n866 585
R51 B.n868 B.n85 585
R52 B.n870 B.n869 585
R53 B.n871 B.n84 585
R54 B.n873 B.n872 585
R55 B.n874 B.n83 585
R56 B.n876 B.n875 585
R57 B.n877 B.n82 585
R58 B.n879 B.n878 585
R59 B.n880 B.n81 585
R60 B.n882 B.n881 585
R61 B.n883 B.n80 585
R62 B.n885 B.n884 585
R63 B.n886 B.n79 585
R64 B.n888 B.n887 585
R65 B.n889 B.n78 585
R66 B.n891 B.n890 585
R67 B.n892 B.n75 585
R68 B.n895 B.n894 585
R69 B.n896 B.n74 585
R70 B.n898 B.n897 585
R71 B.n899 B.n73 585
R72 B.n901 B.n900 585
R73 B.n902 B.n72 585
R74 B.n904 B.n903 585
R75 B.n905 B.n71 585
R76 B.n907 B.n906 585
R77 B.n909 B.n908 585
R78 B.n910 B.n67 585
R79 B.n912 B.n911 585
R80 B.n913 B.n66 585
R81 B.n915 B.n914 585
R82 B.n916 B.n65 585
R83 B.n918 B.n917 585
R84 B.n919 B.n64 585
R85 B.n921 B.n920 585
R86 B.n922 B.n63 585
R87 B.n924 B.n923 585
R88 B.n925 B.n62 585
R89 B.n927 B.n926 585
R90 B.n928 B.n61 585
R91 B.n930 B.n929 585
R92 B.n931 B.n60 585
R93 B.n933 B.n932 585
R94 B.n934 B.n59 585
R95 B.n936 B.n935 585
R96 B.n937 B.n58 585
R97 B.n939 B.n938 585
R98 B.n940 B.n57 585
R99 B.n942 B.n941 585
R100 B.n943 B.n56 585
R101 B.n945 B.n944 585
R102 B.n946 B.n55 585
R103 B.n948 B.n947 585
R104 B.n949 B.n54 585
R105 B.n951 B.n950 585
R106 B.n952 B.n53 585
R107 B.n954 B.n953 585
R108 B.n955 B.n52 585
R109 B.n957 B.n956 585
R110 B.n958 B.n51 585
R111 B.n960 B.n959 585
R112 B.n961 B.n50 585
R113 B.n963 B.n962 585
R114 B.n964 B.n49 585
R115 B.n966 B.n965 585
R116 B.n967 B.n48 585
R117 B.n969 B.n968 585
R118 B.n970 B.n47 585
R119 B.n972 B.n971 585
R120 B.n973 B.n46 585
R121 B.n975 B.n974 585
R122 B.n976 B.n45 585
R123 B.n978 B.n977 585
R124 B.n979 B.n44 585
R125 B.n981 B.n980 585
R126 B.n982 B.n43 585
R127 B.n984 B.n983 585
R128 B.n985 B.n42 585
R129 B.n987 B.n986 585
R130 B.n988 B.n41 585
R131 B.n990 B.n989 585
R132 B.n991 B.n40 585
R133 B.n993 B.n992 585
R134 B.n994 B.n39 585
R135 B.n996 B.n995 585
R136 B.n997 B.n38 585
R137 B.n999 B.n998 585
R138 B.n1000 B.n37 585
R139 B.n1002 B.n1001 585
R140 B.n1003 B.n36 585
R141 B.n796 B.n109 585
R142 B.n795 B.n794 585
R143 B.n793 B.n110 585
R144 B.n792 B.n791 585
R145 B.n790 B.n111 585
R146 B.n789 B.n788 585
R147 B.n787 B.n112 585
R148 B.n786 B.n785 585
R149 B.n784 B.n113 585
R150 B.n783 B.n782 585
R151 B.n781 B.n114 585
R152 B.n780 B.n779 585
R153 B.n778 B.n115 585
R154 B.n777 B.n776 585
R155 B.n775 B.n116 585
R156 B.n774 B.n773 585
R157 B.n772 B.n117 585
R158 B.n771 B.n770 585
R159 B.n769 B.n118 585
R160 B.n768 B.n767 585
R161 B.n766 B.n119 585
R162 B.n765 B.n764 585
R163 B.n763 B.n120 585
R164 B.n762 B.n761 585
R165 B.n760 B.n121 585
R166 B.n759 B.n758 585
R167 B.n757 B.n122 585
R168 B.n756 B.n755 585
R169 B.n754 B.n123 585
R170 B.n753 B.n752 585
R171 B.n751 B.n124 585
R172 B.n750 B.n749 585
R173 B.n748 B.n125 585
R174 B.n747 B.n746 585
R175 B.n745 B.n126 585
R176 B.n744 B.n743 585
R177 B.n742 B.n127 585
R178 B.n741 B.n740 585
R179 B.n739 B.n128 585
R180 B.n738 B.n737 585
R181 B.n736 B.n129 585
R182 B.n735 B.n734 585
R183 B.n733 B.n130 585
R184 B.n732 B.n731 585
R185 B.n730 B.n131 585
R186 B.n729 B.n728 585
R187 B.n727 B.n132 585
R188 B.n726 B.n725 585
R189 B.n724 B.n133 585
R190 B.n723 B.n722 585
R191 B.n721 B.n134 585
R192 B.n720 B.n719 585
R193 B.n718 B.n135 585
R194 B.n717 B.n716 585
R195 B.n715 B.n136 585
R196 B.n714 B.n713 585
R197 B.n712 B.n137 585
R198 B.n711 B.n710 585
R199 B.n709 B.n138 585
R200 B.n708 B.n707 585
R201 B.n706 B.n139 585
R202 B.n705 B.n704 585
R203 B.n703 B.n140 585
R204 B.n702 B.n701 585
R205 B.n700 B.n141 585
R206 B.n699 B.n698 585
R207 B.n697 B.n142 585
R208 B.n696 B.n695 585
R209 B.n694 B.n143 585
R210 B.n693 B.n692 585
R211 B.n691 B.n144 585
R212 B.n690 B.n689 585
R213 B.n688 B.n145 585
R214 B.n687 B.n686 585
R215 B.n685 B.n146 585
R216 B.n684 B.n683 585
R217 B.n682 B.n147 585
R218 B.n681 B.n680 585
R219 B.n679 B.n148 585
R220 B.n678 B.n677 585
R221 B.n676 B.n149 585
R222 B.n675 B.n674 585
R223 B.n673 B.n150 585
R224 B.n672 B.n671 585
R225 B.n670 B.n151 585
R226 B.n669 B.n668 585
R227 B.n667 B.n152 585
R228 B.n666 B.n665 585
R229 B.n664 B.n153 585
R230 B.n663 B.n662 585
R231 B.n661 B.n154 585
R232 B.n660 B.n659 585
R233 B.n658 B.n155 585
R234 B.n657 B.n656 585
R235 B.n655 B.n156 585
R236 B.n654 B.n653 585
R237 B.n652 B.n157 585
R238 B.n651 B.n650 585
R239 B.n649 B.n158 585
R240 B.n648 B.n647 585
R241 B.n646 B.n159 585
R242 B.n645 B.n644 585
R243 B.n643 B.n160 585
R244 B.n642 B.n641 585
R245 B.n640 B.n161 585
R246 B.n639 B.n638 585
R247 B.n637 B.n162 585
R248 B.n636 B.n635 585
R249 B.n634 B.n163 585
R250 B.n633 B.n632 585
R251 B.n631 B.n164 585
R252 B.n630 B.n629 585
R253 B.n628 B.n165 585
R254 B.n627 B.n626 585
R255 B.n625 B.n166 585
R256 B.n624 B.n623 585
R257 B.n622 B.n167 585
R258 B.n621 B.n620 585
R259 B.n619 B.n168 585
R260 B.n618 B.n617 585
R261 B.n616 B.n169 585
R262 B.n615 B.n614 585
R263 B.n613 B.n170 585
R264 B.n612 B.n611 585
R265 B.n610 B.n171 585
R266 B.n609 B.n608 585
R267 B.n607 B.n172 585
R268 B.n606 B.n605 585
R269 B.n604 B.n173 585
R270 B.n603 B.n602 585
R271 B.n601 B.n174 585
R272 B.n600 B.n599 585
R273 B.n598 B.n175 585
R274 B.n597 B.n596 585
R275 B.n595 B.n176 585
R276 B.n594 B.n593 585
R277 B.n592 B.n177 585
R278 B.n385 B.n250 585
R279 B.n387 B.n386 585
R280 B.n388 B.n249 585
R281 B.n390 B.n389 585
R282 B.n391 B.n248 585
R283 B.n393 B.n392 585
R284 B.n394 B.n247 585
R285 B.n396 B.n395 585
R286 B.n397 B.n246 585
R287 B.n399 B.n398 585
R288 B.n400 B.n245 585
R289 B.n402 B.n401 585
R290 B.n403 B.n244 585
R291 B.n405 B.n404 585
R292 B.n406 B.n243 585
R293 B.n408 B.n407 585
R294 B.n409 B.n242 585
R295 B.n411 B.n410 585
R296 B.n412 B.n241 585
R297 B.n414 B.n413 585
R298 B.n415 B.n240 585
R299 B.n417 B.n416 585
R300 B.n418 B.n239 585
R301 B.n420 B.n419 585
R302 B.n421 B.n238 585
R303 B.n423 B.n422 585
R304 B.n424 B.n237 585
R305 B.n426 B.n425 585
R306 B.n427 B.n236 585
R307 B.n429 B.n428 585
R308 B.n430 B.n235 585
R309 B.n432 B.n431 585
R310 B.n433 B.n234 585
R311 B.n435 B.n434 585
R312 B.n436 B.n233 585
R313 B.n438 B.n437 585
R314 B.n439 B.n232 585
R315 B.n441 B.n440 585
R316 B.n442 B.n231 585
R317 B.n444 B.n443 585
R318 B.n445 B.n230 585
R319 B.n447 B.n446 585
R320 B.n448 B.n229 585
R321 B.n450 B.n449 585
R322 B.n451 B.n228 585
R323 B.n453 B.n452 585
R324 B.n454 B.n227 585
R325 B.n456 B.n455 585
R326 B.n457 B.n226 585
R327 B.n459 B.n458 585
R328 B.n460 B.n225 585
R329 B.n462 B.n461 585
R330 B.n463 B.n224 585
R331 B.n465 B.n464 585
R332 B.n466 B.n223 585
R333 B.n468 B.n467 585
R334 B.n469 B.n222 585
R335 B.n471 B.n470 585
R336 B.n472 B.n221 585
R337 B.n474 B.n473 585
R338 B.n475 B.n220 585
R339 B.n477 B.n476 585
R340 B.n478 B.n219 585
R341 B.n480 B.n479 585
R342 B.n482 B.n481 585
R343 B.n483 B.n215 585
R344 B.n485 B.n484 585
R345 B.n486 B.n214 585
R346 B.n488 B.n487 585
R347 B.n489 B.n213 585
R348 B.n491 B.n490 585
R349 B.n492 B.n212 585
R350 B.n494 B.n493 585
R351 B.n496 B.n209 585
R352 B.n498 B.n497 585
R353 B.n499 B.n208 585
R354 B.n501 B.n500 585
R355 B.n502 B.n207 585
R356 B.n504 B.n503 585
R357 B.n505 B.n206 585
R358 B.n507 B.n506 585
R359 B.n508 B.n205 585
R360 B.n510 B.n509 585
R361 B.n511 B.n204 585
R362 B.n513 B.n512 585
R363 B.n514 B.n203 585
R364 B.n516 B.n515 585
R365 B.n517 B.n202 585
R366 B.n519 B.n518 585
R367 B.n520 B.n201 585
R368 B.n522 B.n521 585
R369 B.n523 B.n200 585
R370 B.n525 B.n524 585
R371 B.n526 B.n199 585
R372 B.n528 B.n527 585
R373 B.n529 B.n198 585
R374 B.n531 B.n530 585
R375 B.n532 B.n197 585
R376 B.n534 B.n533 585
R377 B.n535 B.n196 585
R378 B.n537 B.n536 585
R379 B.n538 B.n195 585
R380 B.n540 B.n539 585
R381 B.n541 B.n194 585
R382 B.n543 B.n542 585
R383 B.n544 B.n193 585
R384 B.n546 B.n545 585
R385 B.n547 B.n192 585
R386 B.n549 B.n548 585
R387 B.n550 B.n191 585
R388 B.n552 B.n551 585
R389 B.n553 B.n190 585
R390 B.n555 B.n554 585
R391 B.n556 B.n189 585
R392 B.n558 B.n557 585
R393 B.n559 B.n188 585
R394 B.n561 B.n560 585
R395 B.n562 B.n187 585
R396 B.n564 B.n563 585
R397 B.n565 B.n186 585
R398 B.n567 B.n566 585
R399 B.n568 B.n185 585
R400 B.n570 B.n569 585
R401 B.n571 B.n184 585
R402 B.n573 B.n572 585
R403 B.n574 B.n183 585
R404 B.n576 B.n575 585
R405 B.n577 B.n182 585
R406 B.n579 B.n578 585
R407 B.n580 B.n181 585
R408 B.n582 B.n581 585
R409 B.n583 B.n180 585
R410 B.n585 B.n584 585
R411 B.n586 B.n179 585
R412 B.n588 B.n587 585
R413 B.n589 B.n178 585
R414 B.n591 B.n590 585
R415 B.n384 B.n383 585
R416 B.n382 B.n251 585
R417 B.n381 B.n380 585
R418 B.n379 B.n252 585
R419 B.n378 B.n377 585
R420 B.n376 B.n253 585
R421 B.n375 B.n374 585
R422 B.n373 B.n254 585
R423 B.n372 B.n371 585
R424 B.n370 B.n255 585
R425 B.n369 B.n368 585
R426 B.n367 B.n256 585
R427 B.n366 B.n365 585
R428 B.n364 B.n257 585
R429 B.n363 B.n362 585
R430 B.n361 B.n258 585
R431 B.n360 B.n359 585
R432 B.n358 B.n259 585
R433 B.n357 B.n356 585
R434 B.n355 B.n260 585
R435 B.n354 B.n353 585
R436 B.n352 B.n261 585
R437 B.n351 B.n350 585
R438 B.n349 B.n262 585
R439 B.n348 B.n347 585
R440 B.n346 B.n263 585
R441 B.n345 B.n344 585
R442 B.n343 B.n264 585
R443 B.n342 B.n341 585
R444 B.n340 B.n265 585
R445 B.n339 B.n338 585
R446 B.n337 B.n266 585
R447 B.n336 B.n335 585
R448 B.n334 B.n267 585
R449 B.n333 B.n332 585
R450 B.n331 B.n268 585
R451 B.n330 B.n329 585
R452 B.n328 B.n269 585
R453 B.n327 B.n326 585
R454 B.n325 B.n270 585
R455 B.n324 B.n323 585
R456 B.n322 B.n271 585
R457 B.n321 B.n320 585
R458 B.n319 B.n272 585
R459 B.n318 B.n317 585
R460 B.n316 B.n273 585
R461 B.n315 B.n314 585
R462 B.n313 B.n274 585
R463 B.n312 B.n311 585
R464 B.n310 B.n275 585
R465 B.n309 B.n308 585
R466 B.n307 B.n276 585
R467 B.n306 B.n305 585
R468 B.n304 B.n277 585
R469 B.n303 B.n302 585
R470 B.n301 B.n278 585
R471 B.n300 B.n299 585
R472 B.n298 B.n279 585
R473 B.n297 B.n296 585
R474 B.n295 B.n280 585
R475 B.n294 B.n293 585
R476 B.n292 B.n281 585
R477 B.n291 B.n290 585
R478 B.n289 B.n282 585
R479 B.n288 B.n287 585
R480 B.n286 B.n283 585
R481 B.n285 B.n284 585
R482 B.n2 B.n0 585
R483 B.n1105 B.n1 585
R484 B.n1104 B.n1103 585
R485 B.n1102 B.n3 585
R486 B.n1101 B.n1100 585
R487 B.n1099 B.n4 585
R488 B.n1098 B.n1097 585
R489 B.n1096 B.n5 585
R490 B.n1095 B.n1094 585
R491 B.n1093 B.n6 585
R492 B.n1092 B.n1091 585
R493 B.n1090 B.n7 585
R494 B.n1089 B.n1088 585
R495 B.n1087 B.n8 585
R496 B.n1086 B.n1085 585
R497 B.n1084 B.n9 585
R498 B.n1083 B.n1082 585
R499 B.n1081 B.n10 585
R500 B.n1080 B.n1079 585
R501 B.n1078 B.n11 585
R502 B.n1077 B.n1076 585
R503 B.n1075 B.n12 585
R504 B.n1074 B.n1073 585
R505 B.n1072 B.n13 585
R506 B.n1071 B.n1070 585
R507 B.n1069 B.n14 585
R508 B.n1068 B.n1067 585
R509 B.n1066 B.n15 585
R510 B.n1065 B.n1064 585
R511 B.n1063 B.n16 585
R512 B.n1062 B.n1061 585
R513 B.n1060 B.n17 585
R514 B.n1059 B.n1058 585
R515 B.n1057 B.n18 585
R516 B.n1056 B.n1055 585
R517 B.n1054 B.n19 585
R518 B.n1053 B.n1052 585
R519 B.n1051 B.n20 585
R520 B.n1050 B.n1049 585
R521 B.n1048 B.n21 585
R522 B.n1047 B.n1046 585
R523 B.n1045 B.n22 585
R524 B.n1044 B.n1043 585
R525 B.n1042 B.n23 585
R526 B.n1041 B.n1040 585
R527 B.n1039 B.n24 585
R528 B.n1038 B.n1037 585
R529 B.n1036 B.n25 585
R530 B.n1035 B.n1034 585
R531 B.n1033 B.n26 585
R532 B.n1032 B.n1031 585
R533 B.n1030 B.n27 585
R534 B.n1029 B.n1028 585
R535 B.n1027 B.n28 585
R536 B.n1026 B.n1025 585
R537 B.n1024 B.n29 585
R538 B.n1023 B.n1022 585
R539 B.n1021 B.n30 585
R540 B.n1020 B.n1019 585
R541 B.n1018 B.n31 585
R542 B.n1017 B.n1016 585
R543 B.n1015 B.n32 585
R544 B.n1014 B.n1013 585
R545 B.n1012 B.n33 585
R546 B.n1011 B.n1010 585
R547 B.n1009 B.n34 585
R548 B.n1008 B.n1007 585
R549 B.n1006 B.n35 585
R550 B.n1005 B.n1004 585
R551 B.n1107 B.n1106 585
R552 B.n211 B.t4 509.483
R553 B.n77 B.t8 509.483
R554 B.n217 B.t1 509.483
R555 B.n69 B.t11 509.483
R556 B.n385 B.n384 434.841
R557 B.n1004 B.n1003 434.841
R558 B.n590 B.n177 434.841
R559 B.n798 B.n109 434.841
R560 B.n210 B.t3 334.894
R561 B.n216 B.t0 334.894
R562 B.n68 B.t9 334.894
R563 B.n76 B.t6 334.894
R564 B.n384 B.n251 163.367
R565 B.n380 B.n251 163.367
R566 B.n380 B.n379 163.367
R567 B.n379 B.n378 163.367
R568 B.n378 B.n253 163.367
R569 B.n374 B.n253 163.367
R570 B.n374 B.n373 163.367
R571 B.n373 B.n372 163.367
R572 B.n372 B.n255 163.367
R573 B.n368 B.n255 163.367
R574 B.n368 B.n367 163.367
R575 B.n367 B.n366 163.367
R576 B.n366 B.n257 163.367
R577 B.n362 B.n257 163.367
R578 B.n362 B.n361 163.367
R579 B.n361 B.n360 163.367
R580 B.n360 B.n259 163.367
R581 B.n356 B.n259 163.367
R582 B.n356 B.n355 163.367
R583 B.n355 B.n354 163.367
R584 B.n354 B.n261 163.367
R585 B.n350 B.n261 163.367
R586 B.n350 B.n349 163.367
R587 B.n349 B.n348 163.367
R588 B.n348 B.n263 163.367
R589 B.n344 B.n263 163.367
R590 B.n344 B.n343 163.367
R591 B.n343 B.n342 163.367
R592 B.n342 B.n265 163.367
R593 B.n338 B.n265 163.367
R594 B.n338 B.n337 163.367
R595 B.n337 B.n336 163.367
R596 B.n336 B.n267 163.367
R597 B.n332 B.n267 163.367
R598 B.n332 B.n331 163.367
R599 B.n331 B.n330 163.367
R600 B.n330 B.n269 163.367
R601 B.n326 B.n269 163.367
R602 B.n326 B.n325 163.367
R603 B.n325 B.n324 163.367
R604 B.n324 B.n271 163.367
R605 B.n320 B.n271 163.367
R606 B.n320 B.n319 163.367
R607 B.n319 B.n318 163.367
R608 B.n318 B.n273 163.367
R609 B.n314 B.n273 163.367
R610 B.n314 B.n313 163.367
R611 B.n313 B.n312 163.367
R612 B.n312 B.n275 163.367
R613 B.n308 B.n275 163.367
R614 B.n308 B.n307 163.367
R615 B.n307 B.n306 163.367
R616 B.n306 B.n277 163.367
R617 B.n302 B.n277 163.367
R618 B.n302 B.n301 163.367
R619 B.n301 B.n300 163.367
R620 B.n300 B.n279 163.367
R621 B.n296 B.n279 163.367
R622 B.n296 B.n295 163.367
R623 B.n295 B.n294 163.367
R624 B.n294 B.n281 163.367
R625 B.n290 B.n281 163.367
R626 B.n290 B.n289 163.367
R627 B.n289 B.n288 163.367
R628 B.n288 B.n283 163.367
R629 B.n284 B.n283 163.367
R630 B.n284 B.n2 163.367
R631 B.n1106 B.n2 163.367
R632 B.n1106 B.n1105 163.367
R633 B.n1105 B.n1104 163.367
R634 B.n1104 B.n3 163.367
R635 B.n1100 B.n3 163.367
R636 B.n1100 B.n1099 163.367
R637 B.n1099 B.n1098 163.367
R638 B.n1098 B.n5 163.367
R639 B.n1094 B.n5 163.367
R640 B.n1094 B.n1093 163.367
R641 B.n1093 B.n1092 163.367
R642 B.n1092 B.n7 163.367
R643 B.n1088 B.n7 163.367
R644 B.n1088 B.n1087 163.367
R645 B.n1087 B.n1086 163.367
R646 B.n1086 B.n9 163.367
R647 B.n1082 B.n9 163.367
R648 B.n1082 B.n1081 163.367
R649 B.n1081 B.n1080 163.367
R650 B.n1080 B.n11 163.367
R651 B.n1076 B.n11 163.367
R652 B.n1076 B.n1075 163.367
R653 B.n1075 B.n1074 163.367
R654 B.n1074 B.n13 163.367
R655 B.n1070 B.n13 163.367
R656 B.n1070 B.n1069 163.367
R657 B.n1069 B.n1068 163.367
R658 B.n1068 B.n15 163.367
R659 B.n1064 B.n15 163.367
R660 B.n1064 B.n1063 163.367
R661 B.n1063 B.n1062 163.367
R662 B.n1062 B.n17 163.367
R663 B.n1058 B.n17 163.367
R664 B.n1058 B.n1057 163.367
R665 B.n1057 B.n1056 163.367
R666 B.n1056 B.n19 163.367
R667 B.n1052 B.n19 163.367
R668 B.n1052 B.n1051 163.367
R669 B.n1051 B.n1050 163.367
R670 B.n1050 B.n21 163.367
R671 B.n1046 B.n21 163.367
R672 B.n1046 B.n1045 163.367
R673 B.n1045 B.n1044 163.367
R674 B.n1044 B.n23 163.367
R675 B.n1040 B.n23 163.367
R676 B.n1040 B.n1039 163.367
R677 B.n1039 B.n1038 163.367
R678 B.n1038 B.n25 163.367
R679 B.n1034 B.n25 163.367
R680 B.n1034 B.n1033 163.367
R681 B.n1033 B.n1032 163.367
R682 B.n1032 B.n27 163.367
R683 B.n1028 B.n27 163.367
R684 B.n1028 B.n1027 163.367
R685 B.n1027 B.n1026 163.367
R686 B.n1026 B.n29 163.367
R687 B.n1022 B.n29 163.367
R688 B.n1022 B.n1021 163.367
R689 B.n1021 B.n1020 163.367
R690 B.n1020 B.n31 163.367
R691 B.n1016 B.n31 163.367
R692 B.n1016 B.n1015 163.367
R693 B.n1015 B.n1014 163.367
R694 B.n1014 B.n33 163.367
R695 B.n1010 B.n33 163.367
R696 B.n1010 B.n1009 163.367
R697 B.n1009 B.n1008 163.367
R698 B.n1008 B.n35 163.367
R699 B.n1004 B.n35 163.367
R700 B.n386 B.n385 163.367
R701 B.n386 B.n249 163.367
R702 B.n390 B.n249 163.367
R703 B.n391 B.n390 163.367
R704 B.n392 B.n391 163.367
R705 B.n392 B.n247 163.367
R706 B.n396 B.n247 163.367
R707 B.n397 B.n396 163.367
R708 B.n398 B.n397 163.367
R709 B.n398 B.n245 163.367
R710 B.n402 B.n245 163.367
R711 B.n403 B.n402 163.367
R712 B.n404 B.n403 163.367
R713 B.n404 B.n243 163.367
R714 B.n408 B.n243 163.367
R715 B.n409 B.n408 163.367
R716 B.n410 B.n409 163.367
R717 B.n410 B.n241 163.367
R718 B.n414 B.n241 163.367
R719 B.n415 B.n414 163.367
R720 B.n416 B.n415 163.367
R721 B.n416 B.n239 163.367
R722 B.n420 B.n239 163.367
R723 B.n421 B.n420 163.367
R724 B.n422 B.n421 163.367
R725 B.n422 B.n237 163.367
R726 B.n426 B.n237 163.367
R727 B.n427 B.n426 163.367
R728 B.n428 B.n427 163.367
R729 B.n428 B.n235 163.367
R730 B.n432 B.n235 163.367
R731 B.n433 B.n432 163.367
R732 B.n434 B.n433 163.367
R733 B.n434 B.n233 163.367
R734 B.n438 B.n233 163.367
R735 B.n439 B.n438 163.367
R736 B.n440 B.n439 163.367
R737 B.n440 B.n231 163.367
R738 B.n444 B.n231 163.367
R739 B.n445 B.n444 163.367
R740 B.n446 B.n445 163.367
R741 B.n446 B.n229 163.367
R742 B.n450 B.n229 163.367
R743 B.n451 B.n450 163.367
R744 B.n452 B.n451 163.367
R745 B.n452 B.n227 163.367
R746 B.n456 B.n227 163.367
R747 B.n457 B.n456 163.367
R748 B.n458 B.n457 163.367
R749 B.n458 B.n225 163.367
R750 B.n462 B.n225 163.367
R751 B.n463 B.n462 163.367
R752 B.n464 B.n463 163.367
R753 B.n464 B.n223 163.367
R754 B.n468 B.n223 163.367
R755 B.n469 B.n468 163.367
R756 B.n470 B.n469 163.367
R757 B.n470 B.n221 163.367
R758 B.n474 B.n221 163.367
R759 B.n475 B.n474 163.367
R760 B.n476 B.n475 163.367
R761 B.n476 B.n219 163.367
R762 B.n480 B.n219 163.367
R763 B.n481 B.n480 163.367
R764 B.n481 B.n215 163.367
R765 B.n485 B.n215 163.367
R766 B.n486 B.n485 163.367
R767 B.n487 B.n486 163.367
R768 B.n487 B.n213 163.367
R769 B.n491 B.n213 163.367
R770 B.n492 B.n491 163.367
R771 B.n493 B.n492 163.367
R772 B.n493 B.n209 163.367
R773 B.n498 B.n209 163.367
R774 B.n499 B.n498 163.367
R775 B.n500 B.n499 163.367
R776 B.n500 B.n207 163.367
R777 B.n504 B.n207 163.367
R778 B.n505 B.n504 163.367
R779 B.n506 B.n505 163.367
R780 B.n506 B.n205 163.367
R781 B.n510 B.n205 163.367
R782 B.n511 B.n510 163.367
R783 B.n512 B.n511 163.367
R784 B.n512 B.n203 163.367
R785 B.n516 B.n203 163.367
R786 B.n517 B.n516 163.367
R787 B.n518 B.n517 163.367
R788 B.n518 B.n201 163.367
R789 B.n522 B.n201 163.367
R790 B.n523 B.n522 163.367
R791 B.n524 B.n523 163.367
R792 B.n524 B.n199 163.367
R793 B.n528 B.n199 163.367
R794 B.n529 B.n528 163.367
R795 B.n530 B.n529 163.367
R796 B.n530 B.n197 163.367
R797 B.n534 B.n197 163.367
R798 B.n535 B.n534 163.367
R799 B.n536 B.n535 163.367
R800 B.n536 B.n195 163.367
R801 B.n540 B.n195 163.367
R802 B.n541 B.n540 163.367
R803 B.n542 B.n541 163.367
R804 B.n542 B.n193 163.367
R805 B.n546 B.n193 163.367
R806 B.n547 B.n546 163.367
R807 B.n548 B.n547 163.367
R808 B.n548 B.n191 163.367
R809 B.n552 B.n191 163.367
R810 B.n553 B.n552 163.367
R811 B.n554 B.n553 163.367
R812 B.n554 B.n189 163.367
R813 B.n558 B.n189 163.367
R814 B.n559 B.n558 163.367
R815 B.n560 B.n559 163.367
R816 B.n560 B.n187 163.367
R817 B.n564 B.n187 163.367
R818 B.n565 B.n564 163.367
R819 B.n566 B.n565 163.367
R820 B.n566 B.n185 163.367
R821 B.n570 B.n185 163.367
R822 B.n571 B.n570 163.367
R823 B.n572 B.n571 163.367
R824 B.n572 B.n183 163.367
R825 B.n576 B.n183 163.367
R826 B.n577 B.n576 163.367
R827 B.n578 B.n577 163.367
R828 B.n578 B.n181 163.367
R829 B.n582 B.n181 163.367
R830 B.n583 B.n582 163.367
R831 B.n584 B.n583 163.367
R832 B.n584 B.n179 163.367
R833 B.n588 B.n179 163.367
R834 B.n589 B.n588 163.367
R835 B.n590 B.n589 163.367
R836 B.n594 B.n177 163.367
R837 B.n595 B.n594 163.367
R838 B.n596 B.n595 163.367
R839 B.n596 B.n175 163.367
R840 B.n600 B.n175 163.367
R841 B.n601 B.n600 163.367
R842 B.n602 B.n601 163.367
R843 B.n602 B.n173 163.367
R844 B.n606 B.n173 163.367
R845 B.n607 B.n606 163.367
R846 B.n608 B.n607 163.367
R847 B.n608 B.n171 163.367
R848 B.n612 B.n171 163.367
R849 B.n613 B.n612 163.367
R850 B.n614 B.n613 163.367
R851 B.n614 B.n169 163.367
R852 B.n618 B.n169 163.367
R853 B.n619 B.n618 163.367
R854 B.n620 B.n619 163.367
R855 B.n620 B.n167 163.367
R856 B.n624 B.n167 163.367
R857 B.n625 B.n624 163.367
R858 B.n626 B.n625 163.367
R859 B.n626 B.n165 163.367
R860 B.n630 B.n165 163.367
R861 B.n631 B.n630 163.367
R862 B.n632 B.n631 163.367
R863 B.n632 B.n163 163.367
R864 B.n636 B.n163 163.367
R865 B.n637 B.n636 163.367
R866 B.n638 B.n637 163.367
R867 B.n638 B.n161 163.367
R868 B.n642 B.n161 163.367
R869 B.n643 B.n642 163.367
R870 B.n644 B.n643 163.367
R871 B.n644 B.n159 163.367
R872 B.n648 B.n159 163.367
R873 B.n649 B.n648 163.367
R874 B.n650 B.n649 163.367
R875 B.n650 B.n157 163.367
R876 B.n654 B.n157 163.367
R877 B.n655 B.n654 163.367
R878 B.n656 B.n655 163.367
R879 B.n656 B.n155 163.367
R880 B.n660 B.n155 163.367
R881 B.n661 B.n660 163.367
R882 B.n662 B.n661 163.367
R883 B.n662 B.n153 163.367
R884 B.n666 B.n153 163.367
R885 B.n667 B.n666 163.367
R886 B.n668 B.n667 163.367
R887 B.n668 B.n151 163.367
R888 B.n672 B.n151 163.367
R889 B.n673 B.n672 163.367
R890 B.n674 B.n673 163.367
R891 B.n674 B.n149 163.367
R892 B.n678 B.n149 163.367
R893 B.n679 B.n678 163.367
R894 B.n680 B.n679 163.367
R895 B.n680 B.n147 163.367
R896 B.n684 B.n147 163.367
R897 B.n685 B.n684 163.367
R898 B.n686 B.n685 163.367
R899 B.n686 B.n145 163.367
R900 B.n690 B.n145 163.367
R901 B.n691 B.n690 163.367
R902 B.n692 B.n691 163.367
R903 B.n692 B.n143 163.367
R904 B.n696 B.n143 163.367
R905 B.n697 B.n696 163.367
R906 B.n698 B.n697 163.367
R907 B.n698 B.n141 163.367
R908 B.n702 B.n141 163.367
R909 B.n703 B.n702 163.367
R910 B.n704 B.n703 163.367
R911 B.n704 B.n139 163.367
R912 B.n708 B.n139 163.367
R913 B.n709 B.n708 163.367
R914 B.n710 B.n709 163.367
R915 B.n710 B.n137 163.367
R916 B.n714 B.n137 163.367
R917 B.n715 B.n714 163.367
R918 B.n716 B.n715 163.367
R919 B.n716 B.n135 163.367
R920 B.n720 B.n135 163.367
R921 B.n721 B.n720 163.367
R922 B.n722 B.n721 163.367
R923 B.n722 B.n133 163.367
R924 B.n726 B.n133 163.367
R925 B.n727 B.n726 163.367
R926 B.n728 B.n727 163.367
R927 B.n728 B.n131 163.367
R928 B.n732 B.n131 163.367
R929 B.n733 B.n732 163.367
R930 B.n734 B.n733 163.367
R931 B.n734 B.n129 163.367
R932 B.n738 B.n129 163.367
R933 B.n739 B.n738 163.367
R934 B.n740 B.n739 163.367
R935 B.n740 B.n127 163.367
R936 B.n744 B.n127 163.367
R937 B.n745 B.n744 163.367
R938 B.n746 B.n745 163.367
R939 B.n746 B.n125 163.367
R940 B.n750 B.n125 163.367
R941 B.n751 B.n750 163.367
R942 B.n752 B.n751 163.367
R943 B.n752 B.n123 163.367
R944 B.n756 B.n123 163.367
R945 B.n757 B.n756 163.367
R946 B.n758 B.n757 163.367
R947 B.n758 B.n121 163.367
R948 B.n762 B.n121 163.367
R949 B.n763 B.n762 163.367
R950 B.n764 B.n763 163.367
R951 B.n764 B.n119 163.367
R952 B.n768 B.n119 163.367
R953 B.n769 B.n768 163.367
R954 B.n770 B.n769 163.367
R955 B.n770 B.n117 163.367
R956 B.n774 B.n117 163.367
R957 B.n775 B.n774 163.367
R958 B.n776 B.n775 163.367
R959 B.n776 B.n115 163.367
R960 B.n780 B.n115 163.367
R961 B.n781 B.n780 163.367
R962 B.n782 B.n781 163.367
R963 B.n782 B.n113 163.367
R964 B.n786 B.n113 163.367
R965 B.n787 B.n786 163.367
R966 B.n788 B.n787 163.367
R967 B.n788 B.n111 163.367
R968 B.n792 B.n111 163.367
R969 B.n793 B.n792 163.367
R970 B.n794 B.n793 163.367
R971 B.n794 B.n109 163.367
R972 B.n1003 B.n1002 163.367
R973 B.n1002 B.n37 163.367
R974 B.n998 B.n37 163.367
R975 B.n998 B.n997 163.367
R976 B.n997 B.n996 163.367
R977 B.n996 B.n39 163.367
R978 B.n992 B.n39 163.367
R979 B.n992 B.n991 163.367
R980 B.n991 B.n990 163.367
R981 B.n990 B.n41 163.367
R982 B.n986 B.n41 163.367
R983 B.n986 B.n985 163.367
R984 B.n985 B.n984 163.367
R985 B.n984 B.n43 163.367
R986 B.n980 B.n43 163.367
R987 B.n980 B.n979 163.367
R988 B.n979 B.n978 163.367
R989 B.n978 B.n45 163.367
R990 B.n974 B.n45 163.367
R991 B.n974 B.n973 163.367
R992 B.n973 B.n972 163.367
R993 B.n972 B.n47 163.367
R994 B.n968 B.n47 163.367
R995 B.n968 B.n967 163.367
R996 B.n967 B.n966 163.367
R997 B.n966 B.n49 163.367
R998 B.n962 B.n49 163.367
R999 B.n962 B.n961 163.367
R1000 B.n961 B.n960 163.367
R1001 B.n960 B.n51 163.367
R1002 B.n956 B.n51 163.367
R1003 B.n956 B.n955 163.367
R1004 B.n955 B.n954 163.367
R1005 B.n954 B.n53 163.367
R1006 B.n950 B.n53 163.367
R1007 B.n950 B.n949 163.367
R1008 B.n949 B.n948 163.367
R1009 B.n948 B.n55 163.367
R1010 B.n944 B.n55 163.367
R1011 B.n944 B.n943 163.367
R1012 B.n943 B.n942 163.367
R1013 B.n942 B.n57 163.367
R1014 B.n938 B.n57 163.367
R1015 B.n938 B.n937 163.367
R1016 B.n937 B.n936 163.367
R1017 B.n936 B.n59 163.367
R1018 B.n932 B.n59 163.367
R1019 B.n932 B.n931 163.367
R1020 B.n931 B.n930 163.367
R1021 B.n930 B.n61 163.367
R1022 B.n926 B.n61 163.367
R1023 B.n926 B.n925 163.367
R1024 B.n925 B.n924 163.367
R1025 B.n924 B.n63 163.367
R1026 B.n920 B.n63 163.367
R1027 B.n920 B.n919 163.367
R1028 B.n919 B.n918 163.367
R1029 B.n918 B.n65 163.367
R1030 B.n914 B.n65 163.367
R1031 B.n914 B.n913 163.367
R1032 B.n913 B.n912 163.367
R1033 B.n912 B.n67 163.367
R1034 B.n908 B.n67 163.367
R1035 B.n908 B.n907 163.367
R1036 B.n907 B.n71 163.367
R1037 B.n903 B.n71 163.367
R1038 B.n903 B.n902 163.367
R1039 B.n902 B.n901 163.367
R1040 B.n901 B.n73 163.367
R1041 B.n897 B.n73 163.367
R1042 B.n897 B.n896 163.367
R1043 B.n896 B.n895 163.367
R1044 B.n895 B.n75 163.367
R1045 B.n890 B.n75 163.367
R1046 B.n890 B.n889 163.367
R1047 B.n889 B.n888 163.367
R1048 B.n888 B.n79 163.367
R1049 B.n884 B.n79 163.367
R1050 B.n884 B.n883 163.367
R1051 B.n883 B.n882 163.367
R1052 B.n882 B.n81 163.367
R1053 B.n878 B.n81 163.367
R1054 B.n878 B.n877 163.367
R1055 B.n877 B.n876 163.367
R1056 B.n876 B.n83 163.367
R1057 B.n872 B.n83 163.367
R1058 B.n872 B.n871 163.367
R1059 B.n871 B.n870 163.367
R1060 B.n870 B.n85 163.367
R1061 B.n866 B.n85 163.367
R1062 B.n866 B.n865 163.367
R1063 B.n865 B.n864 163.367
R1064 B.n864 B.n87 163.367
R1065 B.n860 B.n87 163.367
R1066 B.n860 B.n859 163.367
R1067 B.n859 B.n858 163.367
R1068 B.n858 B.n89 163.367
R1069 B.n854 B.n89 163.367
R1070 B.n854 B.n853 163.367
R1071 B.n853 B.n852 163.367
R1072 B.n852 B.n91 163.367
R1073 B.n848 B.n91 163.367
R1074 B.n848 B.n847 163.367
R1075 B.n847 B.n846 163.367
R1076 B.n846 B.n93 163.367
R1077 B.n842 B.n93 163.367
R1078 B.n842 B.n841 163.367
R1079 B.n841 B.n840 163.367
R1080 B.n840 B.n95 163.367
R1081 B.n836 B.n95 163.367
R1082 B.n836 B.n835 163.367
R1083 B.n835 B.n834 163.367
R1084 B.n834 B.n97 163.367
R1085 B.n830 B.n97 163.367
R1086 B.n830 B.n829 163.367
R1087 B.n829 B.n828 163.367
R1088 B.n828 B.n99 163.367
R1089 B.n824 B.n99 163.367
R1090 B.n824 B.n823 163.367
R1091 B.n823 B.n822 163.367
R1092 B.n822 B.n101 163.367
R1093 B.n818 B.n101 163.367
R1094 B.n818 B.n817 163.367
R1095 B.n817 B.n816 163.367
R1096 B.n816 B.n103 163.367
R1097 B.n812 B.n103 163.367
R1098 B.n812 B.n811 163.367
R1099 B.n811 B.n810 163.367
R1100 B.n810 B.n105 163.367
R1101 B.n806 B.n105 163.367
R1102 B.n806 B.n805 163.367
R1103 B.n805 B.n804 163.367
R1104 B.n804 B.n107 163.367
R1105 B.n800 B.n107 163.367
R1106 B.n800 B.n799 163.367
R1107 B.n799 B.n798 163.367
R1108 B.n211 B.n210 78.7399
R1109 B.n217 B.n216 78.7399
R1110 B.n69 B.n68 78.7399
R1111 B.n77 B.n76 78.7399
R1112 B.n495 B.n211 59.5399
R1113 B.n218 B.n217 59.5399
R1114 B.n70 B.n69 59.5399
R1115 B.n893 B.n77 59.5399
R1116 B.n1005 B.n36 28.2542
R1117 B.n797 B.n796 28.2542
R1118 B.n592 B.n591 28.2542
R1119 B.n383 B.n250 28.2542
R1120 B B.n1107 18.0485
R1121 B.n1001 B.n36 10.6151
R1122 B.n1001 B.n1000 10.6151
R1123 B.n1000 B.n999 10.6151
R1124 B.n999 B.n38 10.6151
R1125 B.n995 B.n38 10.6151
R1126 B.n995 B.n994 10.6151
R1127 B.n994 B.n993 10.6151
R1128 B.n993 B.n40 10.6151
R1129 B.n989 B.n40 10.6151
R1130 B.n989 B.n988 10.6151
R1131 B.n988 B.n987 10.6151
R1132 B.n987 B.n42 10.6151
R1133 B.n983 B.n42 10.6151
R1134 B.n983 B.n982 10.6151
R1135 B.n982 B.n981 10.6151
R1136 B.n981 B.n44 10.6151
R1137 B.n977 B.n44 10.6151
R1138 B.n977 B.n976 10.6151
R1139 B.n976 B.n975 10.6151
R1140 B.n975 B.n46 10.6151
R1141 B.n971 B.n46 10.6151
R1142 B.n971 B.n970 10.6151
R1143 B.n970 B.n969 10.6151
R1144 B.n969 B.n48 10.6151
R1145 B.n965 B.n48 10.6151
R1146 B.n965 B.n964 10.6151
R1147 B.n964 B.n963 10.6151
R1148 B.n963 B.n50 10.6151
R1149 B.n959 B.n50 10.6151
R1150 B.n959 B.n958 10.6151
R1151 B.n958 B.n957 10.6151
R1152 B.n957 B.n52 10.6151
R1153 B.n953 B.n52 10.6151
R1154 B.n953 B.n952 10.6151
R1155 B.n952 B.n951 10.6151
R1156 B.n951 B.n54 10.6151
R1157 B.n947 B.n54 10.6151
R1158 B.n947 B.n946 10.6151
R1159 B.n946 B.n945 10.6151
R1160 B.n945 B.n56 10.6151
R1161 B.n941 B.n56 10.6151
R1162 B.n941 B.n940 10.6151
R1163 B.n940 B.n939 10.6151
R1164 B.n939 B.n58 10.6151
R1165 B.n935 B.n58 10.6151
R1166 B.n935 B.n934 10.6151
R1167 B.n934 B.n933 10.6151
R1168 B.n933 B.n60 10.6151
R1169 B.n929 B.n60 10.6151
R1170 B.n929 B.n928 10.6151
R1171 B.n928 B.n927 10.6151
R1172 B.n927 B.n62 10.6151
R1173 B.n923 B.n62 10.6151
R1174 B.n923 B.n922 10.6151
R1175 B.n922 B.n921 10.6151
R1176 B.n921 B.n64 10.6151
R1177 B.n917 B.n64 10.6151
R1178 B.n917 B.n916 10.6151
R1179 B.n916 B.n915 10.6151
R1180 B.n915 B.n66 10.6151
R1181 B.n911 B.n66 10.6151
R1182 B.n911 B.n910 10.6151
R1183 B.n910 B.n909 10.6151
R1184 B.n906 B.n905 10.6151
R1185 B.n905 B.n904 10.6151
R1186 B.n904 B.n72 10.6151
R1187 B.n900 B.n72 10.6151
R1188 B.n900 B.n899 10.6151
R1189 B.n899 B.n898 10.6151
R1190 B.n898 B.n74 10.6151
R1191 B.n894 B.n74 10.6151
R1192 B.n892 B.n891 10.6151
R1193 B.n891 B.n78 10.6151
R1194 B.n887 B.n78 10.6151
R1195 B.n887 B.n886 10.6151
R1196 B.n886 B.n885 10.6151
R1197 B.n885 B.n80 10.6151
R1198 B.n881 B.n80 10.6151
R1199 B.n881 B.n880 10.6151
R1200 B.n880 B.n879 10.6151
R1201 B.n879 B.n82 10.6151
R1202 B.n875 B.n82 10.6151
R1203 B.n875 B.n874 10.6151
R1204 B.n874 B.n873 10.6151
R1205 B.n873 B.n84 10.6151
R1206 B.n869 B.n84 10.6151
R1207 B.n869 B.n868 10.6151
R1208 B.n868 B.n867 10.6151
R1209 B.n867 B.n86 10.6151
R1210 B.n863 B.n86 10.6151
R1211 B.n863 B.n862 10.6151
R1212 B.n862 B.n861 10.6151
R1213 B.n861 B.n88 10.6151
R1214 B.n857 B.n88 10.6151
R1215 B.n857 B.n856 10.6151
R1216 B.n856 B.n855 10.6151
R1217 B.n855 B.n90 10.6151
R1218 B.n851 B.n90 10.6151
R1219 B.n851 B.n850 10.6151
R1220 B.n850 B.n849 10.6151
R1221 B.n849 B.n92 10.6151
R1222 B.n845 B.n92 10.6151
R1223 B.n845 B.n844 10.6151
R1224 B.n844 B.n843 10.6151
R1225 B.n843 B.n94 10.6151
R1226 B.n839 B.n94 10.6151
R1227 B.n839 B.n838 10.6151
R1228 B.n838 B.n837 10.6151
R1229 B.n837 B.n96 10.6151
R1230 B.n833 B.n96 10.6151
R1231 B.n833 B.n832 10.6151
R1232 B.n832 B.n831 10.6151
R1233 B.n831 B.n98 10.6151
R1234 B.n827 B.n98 10.6151
R1235 B.n827 B.n826 10.6151
R1236 B.n826 B.n825 10.6151
R1237 B.n825 B.n100 10.6151
R1238 B.n821 B.n100 10.6151
R1239 B.n821 B.n820 10.6151
R1240 B.n820 B.n819 10.6151
R1241 B.n819 B.n102 10.6151
R1242 B.n815 B.n102 10.6151
R1243 B.n815 B.n814 10.6151
R1244 B.n814 B.n813 10.6151
R1245 B.n813 B.n104 10.6151
R1246 B.n809 B.n104 10.6151
R1247 B.n809 B.n808 10.6151
R1248 B.n808 B.n807 10.6151
R1249 B.n807 B.n106 10.6151
R1250 B.n803 B.n106 10.6151
R1251 B.n803 B.n802 10.6151
R1252 B.n802 B.n801 10.6151
R1253 B.n801 B.n108 10.6151
R1254 B.n797 B.n108 10.6151
R1255 B.n593 B.n592 10.6151
R1256 B.n593 B.n176 10.6151
R1257 B.n597 B.n176 10.6151
R1258 B.n598 B.n597 10.6151
R1259 B.n599 B.n598 10.6151
R1260 B.n599 B.n174 10.6151
R1261 B.n603 B.n174 10.6151
R1262 B.n604 B.n603 10.6151
R1263 B.n605 B.n604 10.6151
R1264 B.n605 B.n172 10.6151
R1265 B.n609 B.n172 10.6151
R1266 B.n610 B.n609 10.6151
R1267 B.n611 B.n610 10.6151
R1268 B.n611 B.n170 10.6151
R1269 B.n615 B.n170 10.6151
R1270 B.n616 B.n615 10.6151
R1271 B.n617 B.n616 10.6151
R1272 B.n617 B.n168 10.6151
R1273 B.n621 B.n168 10.6151
R1274 B.n622 B.n621 10.6151
R1275 B.n623 B.n622 10.6151
R1276 B.n623 B.n166 10.6151
R1277 B.n627 B.n166 10.6151
R1278 B.n628 B.n627 10.6151
R1279 B.n629 B.n628 10.6151
R1280 B.n629 B.n164 10.6151
R1281 B.n633 B.n164 10.6151
R1282 B.n634 B.n633 10.6151
R1283 B.n635 B.n634 10.6151
R1284 B.n635 B.n162 10.6151
R1285 B.n639 B.n162 10.6151
R1286 B.n640 B.n639 10.6151
R1287 B.n641 B.n640 10.6151
R1288 B.n641 B.n160 10.6151
R1289 B.n645 B.n160 10.6151
R1290 B.n646 B.n645 10.6151
R1291 B.n647 B.n646 10.6151
R1292 B.n647 B.n158 10.6151
R1293 B.n651 B.n158 10.6151
R1294 B.n652 B.n651 10.6151
R1295 B.n653 B.n652 10.6151
R1296 B.n653 B.n156 10.6151
R1297 B.n657 B.n156 10.6151
R1298 B.n658 B.n657 10.6151
R1299 B.n659 B.n658 10.6151
R1300 B.n659 B.n154 10.6151
R1301 B.n663 B.n154 10.6151
R1302 B.n664 B.n663 10.6151
R1303 B.n665 B.n664 10.6151
R1304 B.n665 B.n152 10.6151
R1305 B.n669 B.n152 10.6151
R1306 B.n670 B.n669 10.6151
R1307 B.n671 B.n670 10.6151
R1308 B.n671 B.n150 10.6151
R1309 B.n675 B.n150 10.6151
R1310 B.n676 B.n675 10.6151
R1311 B.n677 B.n676 10.6151
R1312 B.n677 B.n148 10.6151
R1313 B.n681 B.n148 10.6151
R1314 B.n682 B.n681 10.6151
R1315 B.n683 B.n682 10.6151
R1316 B.n683 B.n146 10.6151
R1317 B.n687 B.n146 10.6151
R1318 B.n688 B.n687 10.6151
R1319 B.n689 B.n688 10.6151
R1320 B.n689 B.n144 10.6151
R1321 B.n693 B.n144 10.6151
R1322 B.n694 B.n693 10.6151
R1323 B.n695 B.n694 10.6151
R1324 B.n695 B.n142 10.6151
R1325 B.n699 B.n142 10.6151
R1326 B.n700 B.n699 10.6151
R1327 B.n701 B.n700 10.6151
R1328 B.n701 B.n140 10.6151
R1329 B.n705 B.n140 10.6151
R1330 B.n706 B.n705 10.6151
R1331 B.n707 B.n706 10.6151
R1332 B.n707 B.n138 10.6151
R1333 B.n711 B.n138 10.6151
R1334 B.n712 B.n711 10.6151
R1335 B.n713 B.n712 10.6151
R1336 B.n713 B.n136 10.6151
R1337 B.n717 B.n136 10.6151
R1338 B.n718 B.n717 10.6151
R1339 B.n719 B.n718 10.6151
R1340 B.n719 B.n134 10.6151
R1341 B.n723 B.n134 10.6151
R1342 B.n724 B.n723 10.6151
R1343 B.n725 B.n724 10.6151
R1344 B.n725 B.n132 10.6151
R1345 B.n729 B.n132 10.6151
R1346 B.n730 B.n729 10.6151
R1347 B.n731 B.n730 10.6151
R1348 B.n731 B.n130 10.6151
R1349 B.n735 B.n130 10.6151
R1350 B.n736 B.n735 10.6151
R1351 B.n737 B.n736 10.6151
R1352 B.n737 B.n128 10.6151
R1353 B.n741 B.n128 10.6151
R1354 B.n742 B.n741 10.6151
R1355 B.n743 B.n742 10.6151
R1356 B.n743 B.n126 10.6151
R1357 B.n747 B.n126 10.6151
R1358 B.n748 B.n747 10.6151
R1359 B.n749 B.n748 10.6151
R1360 B.n749 B.n124 10.6151
R1361 B.n753 B.n124 10.6151
R1362 B.n754 B.n753 10.6151
R1363 B.n755 B.n754 10.6151
R1364 B.n755 B.n122 10.6151
R1365 B.n759 B.n122 10.6151
R1366 B.n760 B.n759 10.6151
R1367 B.n761 B.n760 10.6151
R1368 B.n761 B.n120 10.6151
R1369 B.n765 B.n120 10.6151
R1370 B.n766 B.n765 10.6151
R1371 B.n767 B.n766 10.6151
R1372 B.n767 B.n118 10.6151
R1373 B.n771 B.n118 10.6151
R1374 B.n772 B.n771 10.6151
R1375 B.n773 B.n772 10.6151
R1376 B.n773 B.n116 10.6151
R1377 B.n777 B.n116 10.6151
R1378 B.n778 B.n777 10.6151
R1379 B.n779 B.n778 10.6151
R1380 B.n779 B.n114 10.6151
R1381 B.n783 B.n114 10.6151
R1382 B.n784 B.n783 10.6151
R1383 B.n785 B.n784 10.6151
R1384 B.n785 B.n112 10.6151
R1385 B.n789 B.n112 10.6151
R1386 B.n790 B.n789 10.6151
R1387 B.n791 B.n790 10.6151
R1388 B.n791 B.n110 10.6151
R1389 B.n795 B.n110 10.6151
R1390 B.n796 B.n795 10.6151
R1391 B.n387 B.n250 10.6151
R1392 B.n388 B.n387 10.6151
R1393 B.n389 B.n388 10.6151
R1394 B.n389 B.n248 10.6151
R1395 B.n393 B.n248 10.6151
R1396 B.n394 B.n393 10.6151
R1397 B.n395 B.n394 10.6151
R1398 B.n395 B.n246 10.6151
R1399 B.n399 B.n246 10.6151
R1400 B.n400 B.n399 10.6151
R1401 B.n401 B.n400 10.6151
R1402 B.n401 B.n244 10.6151
R1403 B.n405 B.n244 10.6151
R1404 B.n406 B.n405 10.6151
R1405 B.n407 B.n406 10.6151
R1406 B.n407 B.n242 10.6151
R1407 B.n411 B.n242 10.6151
R1408 B.n412 B.n411 10.6151
R1409 B.n413 B.n412 10.6151
R1410 B.n413 B.n240 10.6151
R1411 B.n417 B.n240 10.6151
R1412 B.n418 B.n417 10.6151
R1413 B.n419 B.n418 10.6151
R1414 B.n419 B.n238 10.6151
R1415 B.n423 B.n238 10.6151
R1416 B.n424 B.n423 10.6151
R1417 B.n425 B.n424 10.6151
R1418 B.n425 B.n236 10.6151
R1419 B.n429 B.n236 10.6151
R1420 B.n430 B.n429 10.6151
R1421 B.n431 B.n430 10.6151
R1422 B.n431 B.n234 10.6151
R1423 B.n435 B.n234 10.6151
R1424 B.n436 B.n435 10.6151
R1425 B.n437 B.n436 10.6151
R1426 B.n437 B.n232 10.6151
R1427 B.n441 B.n232 10.6151
R1428 B.n442 B.n441 10.6151
R1429 B.n443 B.n442 10.6151
R1430 B.n443 B.n230 10.6151
R1431 B.n447 B.n230 10.6151
R1432 B.n448 B.n447 10.6151
R1433 B.n449 B.n448 10.6151
R1434 B.n449 B.n228 10.6151
R1435 B.n453 B.n228 10.6151
R1436 B.n454 B.n453 10.6151
R1437 B.n455 B.n454 10.6151
R1438 B.n455 B.n226 10.6151
R1439 B.n459 B.n226 10.6151
R1440 B.n460 B.n459 10.6151
R1441 B.n461 B.n460 10.6151
R1442 B.n461 B.n224 10.6151
R1443 B.n465 B.n224 10.6151
R1444 B.n466 B.n465 10.6151
R1445 B.n467 B.n466 10.6151
R1446 B.n467 B.n222 10.6151
R1447 B.n471 B.n222 10.6151
R1448 B.n472 B.n471 10.6151
R1449 B.n473 B.n472 10.6151
R1450 B.n473 B.n220 10.6151
R1451 B.n477 B.n220 10.6151
R1452 B.n478 B.n477 10.6151
R1453 B.n479 B.n478 10.6151
R1454 B.n483 B.n482 10.6151
R1455 B.n484 B.n483 10.6151
R1456 B.n484 B.n214 10.6151
R1457 B.n488 B.n214 10.6151
R1458 B.n489 B.n488 10.6151
R1459 B.n490 B.n489 10.6151
R1460 B.n490 B.n212 10.6151
R1461 B.n494 B.n212 10.6151
R1462 B.n497 B.n496 10.6151
R1463 B.n497 B.n208 10.6151
R1464 B.n501 B.n208 10.6151
R1465 B.n502 B.n501 10.6151
R1466 B.n503 B.n502 10.6151
R1467 B.n503 B.n206 10.6151
R1468 B.n507 B.n206 10.6151
R1469 B.n508 B.n507 10.6151
R1470 B.n509 B.n508 10.6151
R1471 B.n509 B.n204 10.6151
R1472 B.n513 B.n204 10.6151
R1473 B.n514 B.n513 10.6151
R1474 B.n515 B.n514 10.6151
R1475 B.n515 B.n202 10.6151
R1476 B.n519 B.n202 10.6151
R1477 B.n520 B.n519 10.6151
R1478 B.n521 B.n520 10.6151
R1479 B.n521 B.n200 10.6151
R1480 B.n525 B.n200 10.6151
R1481 B.n526 B.n525 10.6151
R1482 B.n527 B.n526 10.6151
R1483 B.n527 B.n198 10.6151
R1484 B.n531 B.n198 10.6151
R1485 B.n532 B.n531 10.6151
R1486 B.n533 B.n532 10.6151
R1487 B.n533 B.n196 10.6151
R1488 B.n537 B.n196 10.6151
R1489 B.n538 B.n537 10.6151
R1490 B.n539 B.n538 10.6151
R1491 B.n539 B.n194 10.6151
R1492 B.n543 B.n194 10.6151
R1493 B.n544 B.n543 10.6151
R1494 B.n545 B.n544 10.6151
R1495 B.n545 B.n192 10.6151
R1496 B.n549 B.n192 10.6151
R1497 B.n550 B.n549 10.6151
R1498 B.n551 B.n550 10.6151
R1499 B.n551 B.n190 10.6151
R1500 B.n555 B.n190 10.6151
R1501 B.n556 B.n555 10.6151
R1502 B.n557 B.n556 10.6151
R1503 B.n557 B.n188 10.6151
R1504 B.n561 B.n188 10.6151
R1505 B.n562 B.n561 10.6151
R1506 B.n563 B.n562 10.6151
R1507 B.n563 B.n186 10.6151
R1508 B.n567 B.n186 10.6151
R1509 B.n568 B.n567 10.6151
R1510 B.n569 B.n568 10.6151
R1511 B.n569 B.n184 10.6151
R1512 B.n573 B.n184 10.6151
R1513 B.n574 B.n573 10.6151
R1514 B.n575 B.n574 10.6151
R1515 B.n575 B.n182 10.6151
R1516 B.n579 B.n182 10.6151
R1517 B.n580 B.n579 10.6151
R1518 B.n581 B.n580 10.6151
R1519 B.n581 B.n180 10.6151
R1520 B.n585 B.n180 10.6151
R1521 B.n586 B.n585 10.6151
R1522 B.n587 B.n586 10.6151
R1523 B.n587 B.n178 10.6151
R1524 B.n591 B.n178 10.6151
R1525 B.n383 B.n382 10.6151
R1526 B.n382 B.n381 10.6151
R1527 B.n381 B.n252 10.6151
R1528 B.n377 B.n252 10.6151
R1529 B.n377 B.n376 10.6151
R1530 B.n376 B.n375 10.6151
R1531 B.n375 B.n254 10.6151
R1532 B.n371 B.n254 10.6151
R1533 B.n371 B.n370 10.6151
R1534 B.n370 B.n369 10.6151
R1535 B.n369 B.n256 10.6151
R1536 B.n365 B.n256 10.6151
R1537 B.n365 B.n364 10.6151
R1538 B.n364 B.n363 10.6151
R1539 B.n363 B.n258 10.6151
R1540 B.n359 B.n258 10.6151
R1541 B.n359 B.n358 10.6151
R1542 B.n358 B.n357 10.6151
R1543 B.n357 B.n260 10.6151
R1544 B.n353 B.n260 10.6151
R1545 B.n353 B.n352 10.6151
R1546 B.n352 B.n351 10.6151
R1547 B.n351 B.n262 10.6151
R1548 B.n347 B.n262 10.6151
R1549 B.n347 B.n346 10.6151
R1550 B.n346 B.n345 10.6151
R1551 B.n345 B.n264 10.6151
R1552 B.n341 B.n264 10.6151
R1553 B.n341 B.n340 10.6151
R1554 B.n340 B.n339 10.6151
R1555 B.n339 B.n266 10.6151
R1556 B.n335 B.n266 10.6151
R1557 B.n335 B.n334 10.6151
R1558 B.n334 B.n333 10.6151
R1559 B.n333 B.n268 10.6151
R1560 B.n329 B.n268 10.6151
R1561 B.n329 B.n328 10.6151
R1562 B.n328 B.n327 10.6151
R1563 B.n327 B.n270 10.6151
R1564 B.n323 B.n270 10.6151
R1565 B.n323 B.n322 10.6151
R1566 B.n322 B.n321 10.6151
R1567 B.n321 B.n272 10.6151
R1568 B.n317 B.n272 10.6151
R1569 B.n317 B.n316 10.6151
R1570 B.n316 B.n315 10.6151
R1571 B.n315 B.n274 10.6151
R1572 B.n311 B.n274 10.6151
R1573 B.n311 B.n310 10.6151
R1574 B.n310 B.n309 10.6151
R1575 B.n309 B.n276 10.6151
R1576 B.n305 B.n276 10.6151
R1577 B.n305 B.n304 10.6151
R1578 B.n304 B.n303 10.6151
R1579 B.n303 B.n278 10.6151
R1580 B.n299 B.n278 10.6151
R1581 B.n299 B.n298 10.6151
R1582 B.n298 B.n297 10.6151
R1583 B.n297 B.n280 10.6151
R1584 B.n293 B.n280 10.6151
R1585 B.n293 B.n292 10.6151
R1586 B.n292 B.n291 10.6151
R1587 B.n291 B.n282 10.6151
R1588 B.n287 B.n282 10.6151
R1589 B.n287 B.n286 10.6151
R1590 B.n286 B.n285 10.6151
R1591 B.n285 B.n0 10.6151
R1592 B.n1103 B.n1 10.6151
R1593 B.n1103 B.n1102 10.6151
R1594 B.n1102 B.n1101 10.6151
R1595 B.n1101 B.n4 10.6151
R1596 B.n1097 B.n4 10.6151
R1597 B.n1097 B.n1096 10.6151
R1598 B.n1096 B.n1095 10.6151
R1599 B.n1095 B.n6 10.6151
R1600 B.n1091 B.n6 10.6151
R1601 B.n1091 B.n1090 10.6151
R1602 B.n1090 B.n1089 10.6151
R1603 B.n1089 B.n8 10.6151
R1604 B.n1085 B.n8 10.6151
R1605 B.n1085 B.n1084 10.6151
R1606 B.n1084 B.n1083 10.6151
R1607 B.n1083 B.n10 10.6151
R1608 B.n1079 B.n10 10.6151
R1609 B.n1079 B.n1078 10.6151
R1610 B.n1078 B.n1077 10.6151
R1611 B.n1077 B.n12 10.6151
R1612 B.n1073 B.n12 10.6151
R1613 B.n1073 B.n1072 10.6151
R1614 B.n1072 B.n1071 10.6151
R1615 B.n1071 B.n14 10.6151
R1616 B.n1067 B.n14 10.6151
R1617 B.n1067 B.n1066 10.6151
R1618 B.n1066 B.n1065 10.6151
R1619 B.n1065 B.n16 10.6151
R1620 B.n1061 B.n16 10.6151
R1621 B.n1061 B.n1060 10.6151
R1622 B.n1060 B.n1059 10.6151
R1623 B.n1059 B.n18 10.6151
R1624 B.n1055 B.n18 10.6151
R1625 B.n1055 B.n1054 10.6151
R1626 B.n1054 B.n1053 10.6151
R1627 B.n1053 B.n20 10.6151
R1628 B.n1049 B.n20 10.6151
R1629 B.n1049 B.n1048 10.6151
R1630 B.n1048 B.n1047 10.6151
R1631 B.n1047 B.n22 10.6151
R1632 B.n1043 B.n22 10.6151
R1633 B.n1043 B.n1042 10.6151
R1634 B.n1042 B.n1041 10.6151
R1635 B.n1041 B.n24 10.6151
R1636 B.n1037 B.n24 10.6151
R1637 B.n1037 B.n1036 10.6151
R1638 B.n1036 B.n1035 10.6151
R1639 B.n1035 B.n26 10.6151
R1640 B.n1031 B.n26 10.6151
R1641 B.n1031 B.n1030 10.6151
R1642 B.n1030 B.n1029 10.6151
R1643 B.n1029 B.n28 10.6151
R1644 B.n1025 B.n28 10.6151
R1645 B.n1025 B.n1024 10.6151
R1646 B.n1024 B.n1023 10.6151
R1647 B.n1023 B.n30 10.6151
R1648 B.n1019 B.n30 10.6151
R1649 B.n1019 B.n1018 10.6151
R1650 B.n1018 B.n1017 10.6151
R1651 B.n1017 B.n32 10.6151
R1652 B.n1013 B.n32 10.6151
R1653 B.n1013 B.n1012 10.6151
R1654 B.n1012 B.n1011 10.6151
R1655 B.n1011 B.n34 10.6151
R1656 B.n1007 B.n34 10.6151
R1657 B.n1007 B.n1006 10.6151
R1658 B.n1006 B.n1005 10.6151
R1659 B.n906 B.n70 6.5566
R1660 B.n894 B.n893 6.5566
R1661 B.n482 B.n218 6.5566
R1662 B.n495 B.n494 6.5566
R1663 B.n909 B.n70 4.05904
R1664 B.n893 B.n892 4.05904
R1665 B.n479 B.n218 4.05904
R1666 B.n496 B.n495 4.05904
R1667 B.n1107 B.n0 2.81026
R1668 B.n1107 B.n1 2.81026
R1669 VP.n25 VP.n24 161.3
R1670 VP.n26 VP.n21 161.3
R1671 VP.n28 VP.n27 161.3
R1672 VP.n29 VP.n20 161.3
R1673 VP.n31 VP.n30 161.3
R1674 VP.n32 VP.n19 161.3
R1675 VP.n34 VP.n33 161.3
R1676 VP.n35 VP.n18 161.3
R1677 VP.n38 VP.n37 161.3
R1678 VP.n39 VP.n17 161.3
R1679 VP.n41 VP.n40 161.3
R1680 VP.n42 VP.n16 161.3
R1681 VP.n44 VP.n43 161.3
R1682 VP.n45 VP.n15 161.3
R1683 VP.n47 VP.n46 161.3
R1684 VP.n48 VP.n14 161.3
R1685 VP.n50 VP.n49 161.3
R1686 VP.n93 VP.n92 161.3
R1687 VP.n91 VP.n1 161.3
R1688 VP.n90 VP.n89 161.3
R1689 VP.n88 VP.n2 161.3
R1690 VP.n87 VP.n86 161.3
R1691 VP.n85 VP.n3 161.3
R1692 VP.n84 VP.n83 161.3
R1693 VP.n82 VP.n4 161.3
R1694 VP.n81 VP.n80 161.3
R1695 VP.n78 VP.n5 161.3
R1696 VP.n77 VP.n76 161.3
R1697 VP.n75 VP.n6 161.3
R1698 VP.n74 VP.n73 161.3
R1699 VP.n72 VP.n7 161.3
R1700 VP.n71 VP.n70 161.3
R1701 VP.n69 VP.n8 161.3
R1702 VP.n68 VP.n67 161.3
R1703 VP.n65 VP.n9 161.3
R1704 VP.n64 VP.n63 161.3
R1705 VP.n62 VP.n10 161.3
R1706 VP.n61 VP.n60 161.3
R1707 VP.n59 VP.n11 161.3
R1708 VP.n58 VP.n57 161.3
R1709 VP.n56 VP.n12 161.3
R1710 VP.n55 VP.n54 161.3
R1711 VP.n22 VP.t2 157.768
R1712 VP.n53 VP.t6 125.605
R1713 VP.n66 VP.t3 125.605
R1714 VP.n79 VP.t1 125.605
R1715 VP.n0 VP.t5 125.605
R1716 VP.n13 VP.t0 125.605
R1717 VP.n36 VP.t4 125.605
R1718 VP.n23 VP.t7 125.605
R1719 VP.n53 VP.n52 85.5092
R1720 VP.n94 VP.n0 85.5092
R1721 VP.n51 VP.n13 85.5092
R1722 VP.n23 VP.n22 73.2467
R1723 VP.n52 VP.n51 61.8779
R1724 VP.n60 VP.n59 46.253
R1725 VP.n86 VP.n2 46.253
R1726 VP.n43 VP.n15 46.253
R1727 VP.n73 VP.n72 40.4106
R1728 VP.n73 VP.n6 40.4106
R1729 VP.n30 VP.n19 40.4106
R1730 VP.n30 VP.n29 40.4106
R1731 VP.n60 VP.n10 34.5682
R1732 VP.n86 VP.n85 34.5682
R1733 VP.n43 VP.n42 34.5682
R1734 VP.n54 VP.n12 24.3439
R1735 VP.n58 VP.n12 24.3439
R1736 VP.n59 VP.n58 24.3439
R1737 VP.n64 VP.n10 24.3439
R1738 VP.n65 VP.n64 24.3439
R1739 VP.n67 VP.n8 24.3439
R1740 VP.n71 VP.n8 24.3439
R1741 VP.n72 VP.n71 24.3439
R1742 VP.n77 VP.n6 24.3439
R1743 VP.n78 VP.n77 24.3439
R1744 VP.n80 VP.n78 24.3439
R1745 VP.n84 VP.n4 24.3439
R1746 VP.n85 VP.n84 24.3439
R1747 VP.n90 VP.n2 24.3439
R1748 VP.n91 VP.n90 24.3439
R1749 VP.n92 VP.n91 24.3439
R1750 VP.n47 VP.n15 24.3439
R1751 VP.n48 VP.n47 24.3439
R1752 VP.n49 VP.n48 24.3439
R1753 VP.n34 VP.n19 24.3439
R1754 VP.n35 VP.n34 24.3439
R1755 VP.n37 VP.n35 24.3439
R1756 VP.n41 VP.n17 24.3439
R1757 VP.n42 VP.n41 24.3439
R1758 VP.n24 VP.n21 24.3439
R1759 VP.n28 VP.n21 24.3439
R1760 VP.n29 VP.n28 24.3439
R1761 VP.n66 VP.n65 22.8833
R1762 VP.n79 VP.n4 22.8833
R1763 VP.n36 VP.n17 22.8833
R1764 VP.n54 VP.n53 4.38232
R1765 VP.n92 VP.n0 4.38232
R1766 VP.n49 VP.n13 4.38232
R1767 VP.n25 VP.n22 3.34239
R1768 VP.n67 VP.n66 1.46111
R1769 VP.n80 VP.n79 1.46111
R1770 VP.n37 VP.n36 1.46111
R1771 VP.n24 VP.n23 1.46111
R1772 VP.n51 VP.n50 0.355081
R1773 VP.n55 VP.n52 0.355081
R1774 VP.n94 VP.n93 0.355081
R1775 VP VP.n94 0.26685
R1776 VP.n26 VP.n25 0.189894
R1777 VP.n27 VP.n26 0.189894
R1778 VP.n27 VP.n20 0.189894
R1779 VP.n31 VP.n20 0.189894
R1780 VP.n32 VP.n31 0.189894
R1781 VP.n33 VP.n32 0.189894
R1782 VP.n33 VP.n18 0.189894
R1783 VP.n38 VP.n18 0.189894
R1784 VP.n39 VP.n38 0.189894
R1785 VP.n40 VP.n39 0.189894
R1786 VP.n40 VP.n16 0.189894
R1787 VP.n44 VP.n16 0.189894
R1788 VP.n45 VP.n44 0.189894
R1789 VP.n46 VP.n45 0.189894
R1790 VP.n46 VP.n14 0.189894
R1791 VP.n50 VP.n14 0.189894
R1792 VP.n56 VP.n55 0.189894
R1793 VP.n57 VP.n56 0.189894
R1794 VP.n57 VP.n11 0.189894
R1795 VP.n61 VP.n11 0.189894
R1796 VP.n62 VP.n61 0.189894
R1797 VP.n63 VP.n62 0.189894
R1798 VP.n63 VP.n9 0.189894
R1799 VP.n68 VP.n9 0.189894
R1800 VP.n69 VP.n68 0.189894
R1801 VP.n70 VP.n69 0.189894
R1802 VP.n70 VP.n7 0.189894
R1803 VP.n74 VP.n7 0.189894
R1804 VP.n75 VP.n74 0.189894
R1805 VP.n76 VP.n75 0.189894
R1806 VP.n76 VP.n5 0.189894
R1807 VP.n81 VP.n5 0.189894
R1808 VP.n82 VP.n81 0.189894
R1809 VP.n83 VP.n82 0.189894
R1810 VP.n83 VP.n3 0.189894
R1811 VP.n87 VP.n3 0.189894
R1812 VP.n88 VP.n87 0.189894
R1813 VP.n89 VP.n88 0.189894
R1814 VP.n89 VP.n1 0.189894
R1815 VP.n93 VP.n1 0.189894
R1816 VTAIL.n785 VTAIL.n784 585
R1817 VTAIL.n782 VTAIL.n781 585
R1818 VTAIL.n791 VTAIL.n790 585
R1819 VTAIL.n793 VTAIL.n792 585
R1820 VTAIL.n778 VTAIL.n777 585
R1821 VTAIL.n799 VTAIL.n798 585
R1822 VTAIL.n802 VTAIL.n801 585
R1823 VTAIL.n800 VTAIL.n774 585
R1824 VTAIL.n807 VTAIL.n773 585
R1825 VTAIL.n809 VTAIL.n808 585
R1826 VTAIL.n811 VTAIL.n810 585
R1827 VTAIL.n770 VTAIL.n769 585
R1828 VTAIL.n817 VTAIL.n816 585
R1829 VTAIL.n819 VTAIL.n818 585
R1830 VTAIL.n766 VTAIL.n765 585
R1831 VTAIL.n825 VTAIL.n824 585
R1832 VTAIL.n827 VTAIL.n826 585
R1833 VTAIL.n762 VTAIL.n761 585
R1834 VTAIL.n833 VTAIL.n832 585
R1835 VTAIL.n835 VTAIL.n834 585
R1836 VTAIL.n758 VTAIL.n757 585
R1837 VTAIL.n841 VTAIL.n840 585
R1838 VTAIL.n843 VTAIL.n842 585
R1839 VTAIL.n754 VTAIL.n753 585
R1840 VTAIL.n849 VTAIL.n848 585
R1841 VTAIL.n851 VTAIL.n850 585
R1842 VTAIL.n37 VTAIL.n36 585
R1843 VTAIL.n34 VTAIL.n33 585
R1844 VTAIL.n43 VTAIL.n42 585
R1845 VTAIL.n45 VTAIL.n44 585
R1846 VTAIL.n30 VTAIL.n29 585
R1847 VTAIL.n51 VTAIL.n50 585
R1848 VTAIL.n54 VTAIL.n53 585
R1849 VTAIL.n52 VTAIL.n26 585
R1850 VTAIL.n59 VTAIL.n25 585
R1851 VTAIL.n61 VTAIL.n60 585
R1852 VTAIL.n63 VTAIL.n62 585
R1853 VTAIL.n22 VTAIL.n21 585
R1854 VTAIL.n69 VTAIL.n68 585
R1855 VTAIL.n71 VTAIL.n70 585
R1856 VTAIL.n18 VTAIL.n17 585
R1857 VTAIL.n77 VTAIL.n76 585
R1858 VTAIL.n79 VTAIL.n78 585
R1859 VTAIL.n14 VTAIL.n13 585
R1860 VTAIL.n85 VTAIL.n84 585
R1861 VTAIL.n87 VTAIL.n86 585
R1862 VTAIL.n10 VTAIL.n9 585
R1863 VTAIL.n93 VTAIL.n92 585
R1864 VTAIL.n95 VTAIL.n94 585
R1865 VTAIL.n6 VTAIL.n5 585
R1866 VTAIL.n101 VTAIL.n100 585
R1867 VTAIL.n103 VTAIL.n102 585
R1868 VTAIL.n143 VTAIL.n142 585
R1869 VTAIL.n140 VTAIL.n139 585
R1870 VTAIL.n149 VTAIL.n148 585
R1871 VTAIL.n151 VTAIL.n150 585
R1872 VTAIL.n136 VTAIL.n135 585
R1873 VTAIL.n157 VTAIL.n156 585
R1874 VTAIL.n160 VTAIL.n159 585
R1875 VTAIL.n158 VTAIL.n132 585
R1876 VTAIL.n165 VTAIL.n131 585
R1877 VTAIL.n167 VTAIL.n166 585
R1878 VTAIL.n169 VTAIL.n168 585
R1879 VTAIL.n128 VTAIL.n127 585
R1880 VTAIL.n175 VTAIL.n174 585
R1881 VTAIL.n177 VTAIL.n176 585
R1882 VTAIL.n124 VTAIL.n123 585
R1883 VTAIL.n183 VTAIL.n182 585
R1884 VTAIL.n185 VTAIL.n184 585
R1885 VTAIL.n120 VTAIL.n119 585
R1886 VTAIL.n191 VTAIL.n190 585
R1887 VTAIL.n193 VTAIL.n192 585
R1888 VTAIL.n116 VTAIL.n115 585
R1889 VTAIL.n199 VTAIL.n198 585
R1890 VTAIL.n201 VTAIL.n200 585
R1891 VTAIL.n112 VTAIL.n111 585
R1892 VTAIL.n207 VTAIL.n206 585
R1893 VTAIL.n209 VTAIL.n208 585
R1894 VTAIL.n251 VTAIL.n250 585
R1895 VTAIL.n248 VTAIL.n247 585
R1896 VTAIL.n257 VTAIL.n256 585
R1897 VTAIL.n259 VTAIL.n258 585
R1898 VTAIL.n244 VTAIL.n243 585
R1899 VTAIL.n265 VTAIL.n264 585
R1900 VTAIL.n268 VTAIL.n267 585
R1901 VTAIL.n266 VTAIL.n240 585
R1902 VTAIL.n273 VTAIL.n239 585
R1903 VTAIL.n275 VTAIL.n274 585
R1904 VTAIL.n277 VTAIL.n276 585
R1905 VTAIL.n236 VTAIL.n235 585
R1906 VTAIL.n283 VTAIL.n282 585
R1907 VTAIL.n285 VTAIL.n284 585
R1908 VTAIL.n232 VTAIL.n231 585
R1909 VTAIL.n291 VTAIL.n290 585
R1910 VTAIL.n293 VTAIL.n292 585
R1911 VTAIL.n228 VTAIL.n227 585
R1912 VTAIL.n299 VTAIL.n298 585
R1913 VTAIL.n301 VTAIL.n300 585
R1914 VTAIL.n224 VTAIL.n223 585
R1915 VTAIL.n307 VTAIL.n306 585
R1916 VTAIL.n309 VTAIL.n308 585
R1917 VTAIL.n220 VTAIL.n219 585
R1918 VTAIL.n315 VTAIL.n314 585
R1919 VTAIL.n317 VTAIL.n316 585
R1920 VTAIL.n745 VTAIL.n744 585
R1921 VTAIL.n743 VTAIL.n742 585
R1922 VTAIL.n648 VTAIL.n647 585
R1923 VTAIL.n737 VTAIL.n736 585
R1924 VTAIL.n735 VTAIL.n734 585
R1925 VTAIL.n652 VTAIL.n651 585
R1926 VTAIL.n729 VTAIL.n728 585
R1927 VTAIL.n727 VTAIL.n726 585
R1928 VTAIL.n656 VTAIL.n655 585
R1929 VTAIL.n721 VTAIL.n720 585
R1930 VTAIL.n719 VTAIL.n718 585
R1931 VTAIL.n660 VTAIL.n659 585
R1932 VTAIL.n713 VTAIL.n712 585
R1933 VTAIL.n711 VTAIL.n710 585
R1934 VTAIL.n664 VTAIL.n663 585
R1935 VTAIL.n705 VTAIL.n704 585
R1936 VTAIL.n703 VTAIL.n702 585
R1937 VTAIL.n701 VTAIL.n667 585
R1938 VTAIL.n671 VTAIL.n668 585
R1939 VTAIL.n696 VTAIL.n695 585
R1940 VTAIL.n694 VTAIL.n693 585
R1941 VTAIL.n673 VTAIL.n672 585
R1942 VTAIL.n688 VTAIL.n687 585
R1943 VTAIL.n686 VTAIL.n685 585
R1944 VTAIL.n677 VTAIL.n676 585
R1945 VTAIL.n680 VTAIL.n679 585
R1946 VTAIL.n637 VTAIL.n636 585
R1947 VTAIL.n635 VTAIL.n634 585
R1948 VTAIL.n540 VTAIL.n539 585
R1949 VTAIL.n629 VTAIL.n628 585
R1950 VTAIL.n627 VTAIL.n626 585
R1951 VTAIL.n544 VTAIL.n543 585
R1952 VTAIL.n621 VTAIL.n620 585
R1953 VTAIL.n619 VTAIL.n618 585
R1954 VTAIL.n548 VTAIL.n547 585
R1955 VTAIL.n613 VTAIL.n612 585
R1956 VTAIL.n611 VTAIL.n610 585
R1957 VTAIL.n552 VTAIL.n551 585
R1958 VTAIL.n605 VTAIL.n604 585
R1959 VTAIL.n603 VTAIL.n602 585
R1960 VTAIL.n556 VTAIL.n555 585
R1961 VTAIL.n597 VTAIL.n596 585
R1962 VTAIL.n595 VTAIL.n594 585
R1963 VTAIL.n593 VTAIL.n559 585
R1964 VTAIL.n563 VTAIL.n560 585
R1965 VTAIL.n588 VTAIL.n587 585
R1966 VTAIL.n586 VTAIL.n585 585
R1967 VTAIL.n565 VTAIL.n564 585
R1968 VTAIL.n580 VTAIL.n579 585
R1969 VTAIL.n578 VTAIL.n577 585
R1970 VTAIL.n569 VTAIL.n568 585
R1971 VTAIL.n572 VTAIL.n571 585
R1972 VTAIL.n531 VTAIL.n530 585
R1973 VTAIL.n529 VTAIL.n528 585
R1974 VTAIL.n434 VTAIL.n433 585
R1975 VTAIL.n523 VTAIL.n522 585
R1976 VTAIL.n521 VTAIL.n520 585
R1977 VTAIL.n438 VTAIL.n437 585
R1978 VTAIL.n515 VTAIL.n514 585
R1979 VTAIL.n513 VTAIL.n512 585
R1980 VTAIL.n442 VTAIL.n441 585
R1981 VTAIL.n507 VTAIL.n506 585
R1982 VTAIL.n505 VTAIL.n504 585
R1983 VTAIL.n446 VTAIL.n445 585
R1984 VTAIL.n499 VTAIL.n498 585
R1985 VTAIL.n497 VTAIL.n496 585
R1986 VTAIL.n450 VTAIL.n449 585
R1987 VTAIL.n491 VTAIL.n490 585
R1988 VTAIL.n489 VTAIL.n488 585
R1989 VTAIL.n487 VTAIL.n453 585
R1990 VTAIL.n457 VTAIL.n454 585
R1991 VTAIL.n482 VTAIL.n481 585
R1992 VTAIL.n480 VTAIL.n479 585
R1993 VTAIL.n459 VTAIL.n458 585
R1994 VTAIL.n474 VTAIL.n473 585
R1995 VTAIL.n472 VTAIL.n471 585
R1996 VTAIL.n463 VTAIL.n462 585
R1997 VTAIL.n466 VTAIL.n465 585
R1998 VTAIL.n423 VTAIL.n422 585
R1999 VTAIL.n421 VTAIL.n420 585
R2000 VTAIL.n326 VTAIL.n325 585
R2001 VTAIL.n415 VTAIL.n414 585
R2002 VTAIL.n413 VTAIL.n412 585
R2003 VTAIL.n330 VTAIL.n329 585
R2004 VTAIL.n407 VTAIL.n406 585
R2005 VTAIL.n405 VTAIL.n404 585
R2006 VTAIL.n334 VTAIL.n333 585
R2007 VTAIL.n399 VTAIL.n398 585
R2008 VTAIL.n397 VTAIL.n396 585
R2009 VTAIL.n338 VTAIL.n337 585
R2010 VTAIL.n391 VTAIL.n390 585
R2011 VTAIL.n389 VTAIL.n388 585
R2012 VTAIL.n342 VTAIL.n341 585
R2013 VTAIL.n383 VTAIL.n382 585
R2014 VTAIL.n381 VTAIL.n380 585
R2015 VTAIL.n379 VTAIL.n345 585
R2016 VTAIL.n349 VTAIL.n346 585
R2017 VTAIL.n374 VTAIL.n373 585
R2018 VTAIL.n372 VTAIL.n371 585
R2019 VTAIL.n351 VTAIL.n350 585
R2020 VTAIL.n366 VTAIL.n365 585
R2021 VTAIL.n364 VTAIL.n363 585
R2022 VTAIL.n355 VTAIL.n354 585
R2023 VTAIL.n358 VTAIL.n357 585
R2024 VTAIL.n850 VTAIL.n750 498.474
R2025 VTAIL.n102 VTAIL.n2 498.474
R2026 VTAIL.n208 VTAIL.n108 498.474
R2027 VTAIL.n316 VTAIL.n216 498.474
R2028 VTAIL.n744 VTAIL.n644 498.474
R2029 VTAIL.n636 VTAIL.n536 498.474
R2030 VTAIL.n530 VTAIL.n430 498.474
R2031 VTAIL.n422 VTAIL.n322 498.474
R2032 VTAIL.t11 VTAIL.n783 329.036
R2033 VTAIL.t1 VTAIL.n35 329.036
R2034 VTAIL.t5 VTAIL.n141 329.036
R2035 VTAIL.t8 VTAIL.n249 329.036
R2036 VTAIL.t9 VTAIL.n678 329.036
R2037 VTAIL.t3 VTAIL.n570 329.036
R2038 VTAIL.t14 VTAIL.n464 329.036
R2039 VTAIL.t13 VTAIL.n356 329.036
R2040 VTAIL.n784 VTAIL.n781 171.744
R2041 VTAIL.n791 VTAIL.n781 171.744
R2042 VTAIL.n792 VTAIL.n791 171.744
R2043 VTAIL.n792 VTAIL.n777 171.744
R2044 VTAIL.n799 VTAIL.n777 171.744
R2045 VTAIL.n801 VTAIL.n799 171.744
R2046 VTAIL.n801 VTAIL.n800 171.744
R2047 VTAIL.n800 VTAIL.n773 171.744
R2048 VTAIL.n809 VTAIL.n773 171.744
R2049 VTAIL.n810 VTAIL.n809 171.744
R2050 VTAIL.n810 VTAIL.n769 171.744
R2051 VTAIL.n817 VTAIL.n769 171.744
R2052 VTAIL.n818 VTAIL.n817 171.744
R2053 VTAIL.n818 VTAIL.n765 171.744
R2054 VTAIL.n825 VTAIL.n765 171.744
R2055 VTAIL.n826 VTAIL.n825 171.744
R2056 VTAIL.n826 VTAIL.n761 171.744
R2057 VTAIL.n833 VTAIL.n761 171.744
R2058 VTAIL.n834 VTAIL.n833 171.744
R2059 VTAIL.n834 VTAIL.n757 171.744
R2060 VTAIL.n841 VTAIL.n757 171.744
R2061 VTAIL.n842 VTAIL.n841 171.744
R2062 VTAIL.n842 VTAIL.n753 171.744
R2063 VTAIL.n849 VTAIL.n753 171.744
R2064 VTAIL.n850 VTAIL.n849 171.744
R2065 VTAIL.n36 VTAIL.n33 171.744
R2066 VTAIL.n43 VTAIL.n33 171.744
R2067 VTAIL.n44 VTAIL.n43 171.744
R2068 VTAIL.n44 VTAIL.n29 171.744
R2069 VTAIL.n51 VTAIL.n29 171.744
R2070 VTAIL.n53 VTAIL.n51 171.744
R2071 VTAIL.n53 VTAIL.n52 171.744
R2072 VTAIL.n52 VTAIL.n25 171.744
R2073 VTAIL.n61 VTAIL.n25 171.744
R2074 VTAIL.n62 VTAIL.n61 171.744
R2075 VTAIL.n62 VTAIL.n21 171.744
R2076 VTAIL.n69 VTAIL.n21 171.744
R2077 VTAIL.n70 VTAIL.n69 171.744
R2078 VTAIL.n70 VTAIL.n17 171.744
R2079 VTAIL.n77 VTAIL.n17 171.744
R2080 VTAIL.n78 VTAIL.n77 171.744
R2081 VTAIL.n78 VTAIL.n13 171.744
R2082 VTAIL.n85 VTAIL.n13 171.744
R2083 VTAIL.n86 VTAIL.n85 171.744
R2084 VTAIL.n86 VTAIL.n9 171.744
R2085 VTAIL.n93 VTAIL.n9 171.744
R2086 VTAIL.n94 VTAIL.n93 171.744
R2087 VTAIL.n94 VTAIL.n5 171.744
R2088 VTAIL.n101 VTAIL.n5 171.744
R2089 VTAIL.n102 VTAIL.n101 171.744
R2090 VTAIL.n142 VTAIL.n139 171.744
R2091 VTAIL.n149 VTAIL.n139 171.744
R2092 VTAIL.n150 VTAIL.n149 171.744
R2093 VTAIL.n150 VTAIL.n135 171.744
R2094 VTAIL.n157 VTAIL.n135 171.744
R2095 VTAIL.n159 VTAIL.n157 171.744
R2096 VTAIL.n159 VTAIL.n158 171.744
R2097 VTAIL.n158 VTAIL.n131 171.744
R2098 VTAIL.n167 VTAIL.n131 171.744
R2099 VTAIL.n168 VTAIL.n167 171.744
R2100 VTAIL.n168 VTAIL.n127 171.744
R2101 VTAIL.n175 VTAIL.n127 171.744
R2102 VTAIL.n176 VTAIL.n175 171.744
R2103 VTAIL.n176 VTAIL.n123 171.744
R2104 VTAIL.n183 VTAIL.n123 171.744
R2105 VTAIL.n184 VTAIL.n183 171.744
R2106 VTAIL.n184 VTAIL.n119 171.744
R2107 VTAIL.n191 VTAIL.n119 171.744
R2108 VTAIL.n192 VTAIL.n191 171.744
R2109 VTAIL.n192 VTAIL.n115 171.744
R2110 VTAIL.n199 VTAIL.n115 171.744
R2111 VTAIL.n200 VTAIL.n199 171.744
R2112 VTAIL.n200 VTAIL.n111 171.744
R2113 VTAIL.n207 VTAIL.n111 171.744
R2114 VTAIL.n208 VTAIL.n207 171.744
R2115 VTAIL.n250 VTAIL.n247 171.744
R2116 VTAIL.n257 VTAIL.n247 171.744
R2117 VTAIL.n258 VTAIL.n257 171.744
R2118 VTAIL.n258 VTAIL.n243 171.744
R2119 VTAIL.n265 VTAIL.n243 171.744
R2120 VTAIL.n267 VTAIL.n265 171.744
R2121 VTAIL.n267 VTAIL.n266 171.744
R2122 VTAIL.n266 VTAIL.n239 171.744
R2123 VTAIL.n275 VTAIL.n239 171.744
R2124 VTAIL.n276 VTAIL.n275 171.744
R2125 VTAIL.n276 VTAIL.n235 171.744
R2126 VTAIL.n283 VTAIL.n235 171.744
R2127 VTAIL.n284 VTAIL.n283 171.744
R2128 VTAIL.n284 VTAIL.n231 171.744
R2129 VTAIL.n291 VTAIL.n231 171.744
R2130 VTAIL.n292 VTAIL.n291 171.744
R2131 VTAIL.n292 VTAIL.n227 171.744
R2132 VTAIL.n299 VTAIL.n227 171.744
R2133 VTAIL.n300 VTAIL.n299 171.744
R2134 VTAIL.n300 VTAIL.n223 171.744
R2135 VTAIL.n307 VTAIL.n223 171.744
R2136 VTAIL.n308 VTAIL.n307 171.744
R2137 VTAIL.n308 VTAIL.n219 171.744
R2138 VTAIL.n315 VTAIL.n219 171.744
R2139 VTAIL.n316 VTAIL.n315 171.744
R2140 VTAIL.n744 VTAIL.n743 171.744
R2141 VTAIL.n743 VTAIL.n647 171.744
R2142 VTAIL.n736 VTAIL.n647 171.744
R2143 VTAIL.n736 VTAIL.n735 171.744
R2144 VTAIL.n735 VTAIL.n651 171.744
R2145 VTAIL.n728 VTAIL.n651 171.744
R2146 VTAIL.n728 VTAIL.n727 171.744
R2147 VTAIL.n727 VTAIL.n655 171.744
R2148 VTAIL.n720 VTAIL.n655 171.744
R2149 VTAIL.n720 VTAIL.n719 171.744
R2150 VTAIL.n719 VTAIL.n659 171.744
R2151 VTAIL.n712 VTAIL.n659 171.744
R2152 VTAIL.n712 VTAIL.n711 171.744
R2153 VTAIL.n711 VTAIL.n663 171.744
R2154 VTAIL.n704 VTAIL.n663 171.744
R2155 VTAIL.n704 VTAIL.n703 171.744
R2156 VTAIL.n703 VTAIL.n667 171.744
R2157 VTAIL.n671 VTAIL.n667 171.744
R2158 VTAIL.n695 VTAIL.n671 171.744
R2159 VTAIL.n695 VTAIL.n694 171.744
R2160 VTAIL.n694 VTAIL.n672 171.744
R2161 VTAIL.n687 VTAIL.n672 171.744
R2162 VTAIL.n687 VTAIL.n686 171.744
R2163 VTAIL.n686 VTAIL.n676 171.744
R2164 VTAIL.n679 VTAIL.n676 171.744
R2165 VTAIL.n636 VTAIL.n635 171.744
R2166 VTAIL.n635 VTAIL.n539 171.744
R2167 VTAIL.n628 VTAIL.n539 171.744
R2168 VTAIL.n628 VTAIL.n627 171.744
R2169 VTAIL.n627 VTAIL.n543 171.744
R2170 VTAIL.n620 VTAIL.n543 171.744
R2171 VTAIL.n620 VTAIL.n619 171.744
R2172 VTAIL.n619 VTAIL.n547 171.744
R2173 VTAIL.n612 VTAIL.n547 171.744
R2174 VTAIL.n612 VTAIL.n611 171.744
R2175 VTAIL.n611 VTAIL.n551 171.744
R2176 VTAIL.n604 VTAIL.n551 171.744
R2177 VTAIL.n604 VTAIL.n603 171.744
R2178 VTAIL.n603 VTAIL.n555 171.744
R2179 VTAIL.n596 VTAIL.n555 171.744
R2180 VTAIL.n596 VTAIL.n595 171.744
R2181 VTAIL.n595 VTAIL.n559 171.744
R2182 VTAIL.n563 VTAIL.n559 171.744
R2183 VTAIL.n587 VTAIL.n563 171.744
R2184 VTAIL.n587 VTAIL.n586 171.744
R2185 VTAIL.n586 VTAIL.n564 171.744
R2186 VTAIL.n579 VTAIL.n564 171.744
R2187 VTAIL.n579 VTAIL.n578 171.744
R2188 VTAIL.n578 VTAIL.n568 171.744
R2189 VTAIL.n571 VTAIL.n568 171.744
R2190 VTAIL.n530 VTAIL.n529 171.744
R2191 VTAIL.n529 VTAIL.n433 171.744
R2192 VTAIL.n522 VTAIL.n433 171.744
R2193 VTAIL.n522 VTAIL.n521 171.744
R2194 VTAIL.n521 VTAIL.n437 171.744
R2195 VTAIL.n514 VTAIL.n437 171.744
R2196 VTAIL.n514 VTAIL.n513 171.744
R2197 VTAIL.n513 VTAIL.n441 171.744
R2198 VTAIL.n506 VTAIL.n441 171.744
R2199 VTAIL.n506 VTAIL.n505 171.744
R2200 VTAIL.n505 VTAIL.n445 171.744
R2201 VTAIL.n498 VTAIL.n445 171.744
R2202 VTAIL.n498 VTAIL.n497 171.744
R2203 VTAIL.n497 VTAIL.n449 171.744
R2204 VTAIL.n490 VTAIL.n449 171.744
R2205 VTAIL.n490 VTAIL.n489 171.744
R2206 VTAIL.n489 VTAIL.n453 171.744
R2207 VTAIL.n457 VTAIL.n453 171.744
R2208 VTAIL.n481 VTAIL.n457 171.744
R2209 VTAIL.n481 VTAIL.n480 171.744
R2210 VTAIL.n480 VTAIL.n458 171.744
R2211 VTAIL.n473 VTAIL.n458 171.744
R2212 VTAIL.n473 VTAIL.n472 171.744
R2213 VTAIL.n472 VTAIL.n462 171.744
R2214 VTAIL.n465 VTAIL.n462 171.744
R2215 VTAIL.n422 VTAIL.n421 171.744
R2216 VTAIL.n421 VTAIL.n325 171.744
R2217 VTAIL.n414 VTAIL.n325 171.744
R2218 VTAIL.n414 VTAIL.n413 171.744
R2219 VTAIL.n413 VTAIL.n329 171.744
R2220 VTAIL.n406 VTAIL.n329 171.744
R2221 VTAIL.n406 VTAIL.n405 171.744
R2222 VTAIL.n405 VTAIL.n333 171.744
R2223 VTAIL.n398 VTAIL.n333 171.744
R2224 VTAIL.n398 VTAIL.n397 171.744
R2225 VTAIL.n397 VTAIL.n337 171.744
R2226 VTAIL.n390 VTAIL.n337 171.744
R2227 VTAIL.n390 VTAIL.n389 171.744
R2228 VTAIL.n389 VTAIL.n341 171.744
R2229 VTAIL.n382 VTAIL.n341 171.744
R2230 VTAIL.n382 VTAIL.n381 171.744
R2231 VTAIL.n381 VTAIL.n345 171.744
R2232 VTAIL.n349 VTAIL.n345 171.744
R2233 VTAIL.n373 VTAIL.n349 171.744
R2234 VTAIL.n373 VTAIL.n372 171.744
R2235 VTAIL.n372 VTAIL.n350 171.744
R2236 VTAIL.n365 VTAIL.n350 171.744
R2237 VTAIL.n365 VTAIL.n364 171.744
R2238 VTAIL.n364 VTAIL.n354 171.744
R2239 VTAIL.n357 VTAIL.n354 171.744
R2240 VTAIL.n784 VTAIL.t11 85.8723
R2241 VTAIL.n36 VTAIL.t1 85.8723
R2242 VTAIL.n142 VTAIL.t5 85.8723
R2243 VTAIL.n250 VTAIL.t8 85.8723
R2244 VTAIL.n679 VTAIL.t9 85.8723
R2245 VTAIL.n571 VTAIL.t3 85.8723
R2246 VTAIL.n465 VTAIL.t14 85.8723
R2247 VTAIL.n357 VTAIL.t13 85.8723
R2248 VTAIL.n643 VTAIL.n642 53.4917
R2249 VTAIL.n429 VTAIL.n428 53.4917
R2250 VTAIL.n1 VTAIL.n0 53.4916
R2251 VTAIL.n215 VTAIL.n214 53.4916
R2252 VTAIL.n855 VTAIL.n854 34.5126
R2253 VTAIL.n107 VTAIL.n106 34.5126
R2254 VTAIL.n213 VTAIL.n212 34.5126
R2255 VTAIL.n321 VTAIL.n320 34.5126
R2256 VTAIL.n749 VTAIL.n748 34.5126
R2257 VTAIL.n641 VTAIL.n640 34.5126
R2258 VTAIL.n535 VTAIL.n534 34.5126
R2259 VTAIL.n427 VTAIL.n426 34.5126
R2260 VTAIL.n855 VTAIL.n749 32.6255
R2261 VTAIL.n427 VTAIL.n321 32.6255
R2262 VTAIL.n808 VTAIL.n807 13.1884
R2263 VTAIL.n60 VTAIL.n59 13.1884
R2264 VTAIL.n166 VTAIL.n165 13.1884
R2265 VTAIL.n274 VTAIL.n273 13.1884
R2266 VTAIL.n702 VTAIL.n701 13.1884
R2267 VTAIL.n594 VTAIL.n593 13.1884
R2268 VTAIL.n488 VTAIL.n487 13.1884
R2269 VTAIL.n380 VTAIL.n379 13.1884
R2270 VTAIL.n806 VTAIL.n774 12.8005
R2271 VTAIL.n811 VTAIL.n772 12.8005
R2272 VTAIL.n852 VTAIL.n851 12.8005
R2273 VTAIL.n58 VTAIL.n26 12.8005
R2274 VTAIL.n63 VTAIL.n24 12.8005
R2275 VTAIL.n104 VTAIL.n103 12.8005
R2276 VTAIL.n164 VTAIL.n132 12.8005
R2277 VTAIL.n169 VTAIL.n130 12.8005
R2278 VTAIL.n210 VTAIL.n209 12.8005
R2279 VTAIL.n272 VTAIL.n240 12.8005
R2280 VTAIL.n277 VTAIL.n238 12.8005
R2281 VTAIL.n318 VTAIL.n317 12.8005
R2282 VTAIL.n746 VTAIL.n745 12.8005
R2283 VTAIL.n705 VTAIL.n666 12.8005
R2284 VTAIL.n700 VTAIL.n668 12.8005
R2285 VTAIL.n638 VTAIL.n637 12.8005
R2286 VTAIL.n597 VTAIL.n558 12.8005
R2287 VTAIL.n592 VTAIL.n560 12.8005
R2288 VTAIL.n532 VTAIL.n531 12.8005
R2289 VTAIL.n491 VTAIL.n452 12.8005
R2290 VTAIL.n486 VTAIL.n454 12.8005
R2291 VTAIL.n424 VTAIL.n423 12.8005
R2292 VTAIL.n383 VTAIL.n344 12.8005
R2293 VTAIL.n378 VTAIL.n346 12.8005
R2294 VTAIL.n803 VTAIL.n802 12.0247
R2295 VTAIL.n812 VTAIL.n770 12.0247
R2296 VTAIL.n848 VTAIL.n752 12.0247
R2297 VTAIL.n55 VTAIL.n54 12.0247
R2298 VTAIL.n64 VTAIL.n22 12.0247
R2299 VTAIL.n100 VTAIL.n4 12.0247
R2300 VTAIL.n161 VTAIL.n160 12.0247
R2301 VTAIL.n170 VTAIL.n128 12.0247
R2302 VTAIL.n206 VTAIL.n110 12.0247
R2303 VTAIL.n269 VTAIL.n268 12.0247
R2304 VTAIL.n278 VTAIL.n236 12.0247
R2305 VTAIL.n314 VTAIL.n218 12.0247
R2306 VTAIL.n742 VTAIL.n646 12.0247
R2307 VTAIL.n706 VTAIL.n664 12.0247
R2308 VTAIL.n697 VTAIL.n696 12.0247
R2309 VTAIL.n634 VTAIL.n538 12.0247
R2310 VTAIL.n598 VTAIL.n556 12.0247
R2311 VTAIL.n589 VTAIL.n588 12.0247
R2312 VTAIL.n528 VTAIL.n432 12.0247
R2313 VTAIL.n492 VTAIL.n450 12.0247
R2314 VTAIL.n483 VTAIL.n482 12.0247
R2315 VTAIL.n420 VTAIL.n324 12.0247
R2316 VTAIL.n384 VTAIL.n342 12.0247
R2317 VTAIL.n375 VTAIL.n374 12.0247
R2318 VTAIL.n798 VTAIL.n776 11.249
R2319 VTAIL.n816 VTAIL.n815 11.249
R2320 VTAIL.n847 VTAIL.n754 11.249
R2321 VTAIL.n50 VTAIL.n28 11.249
R2322 VTAIL.n68 VTAIL.n67 11.249
R2323 VTAIL.n99 VTAIL.n6 11.249
R2324 VTAIL.n156 VTAIL.n134 11.249
R2325 VTAIL.n174 VTAIL.n173 11.249
R2326 VTAIL.n205 VTAIL.n112 11.249
R2327 VTAIL.n264 VTAIL.n242 11.249
R2328 VTAIL.n282 VTAIL.n281 11.249
R2329 VTAIL.n313 VTAIL.n220 11.249
R2330 VTAIL.n741 VTAIL.n648 11.249
R2331 VTAIL.n710 VTAIL.n709 11.249
R2332 VTAIL.n693 VTAIL.n670 11.249
R2333 VTAIL.n633 VTAIL.n540 11.249
R2334 VTAIL.n602 VTAIL.n601 11.249
R2335 VTAIL.n585 VTAIL.n562 11.249
R2336 VTAIL.n527 VTAIL.n434 11.249
R2337 VTAIL.n496 VTAIL.n495 11.249
R2338 VTAIL.n479 VTAIL.n456 11.249
R2339 VTAIL.n419 VTAIL.n326 11.249
R2340 VTAIL.n388 VTAIL.n387 11.249
R2341 VTAIL.n371 VTAIL.n348 11.249
R2342 VTAIL.n785 VTAIL.n783 10.7239
R2343 VTAIL.n37 VTAIL.n35 10.7239
R2344 VTAIL.n143 VTAIL.n141 10.7239
R2345 VTAIL.n251 VTAIL.n249 10.7239
R2346 VTAIL.n680 VTAIL.n678 10.7239
R2347 VTAIL.n572 VTAIL.n570 10.7239
R2348 VTAIL.n466 VTAIL.n464 10.7239
R2349 VTAIL.n358 VTAIL.n356 10.7239
R2350 VTAIL.n797 VTAIL.n778 10.4732
R2351 VTAIL.n819 VTAIL.n768 10.4732
R2352 VTAIL.n844 VTAIL.n843 10.4732
R2353 VTAIL.n49 VTAIL.n30 10.4732
R2354 VTAIL.n71 VTAIL.n20 10.4732
R2355 VTAIL.n96 VTAIL.n95 10.4732
R2356 VTAIL.n155 VTAIL.n136 10.4732
R2357 VTAIL.n177 VTAIL.n126 10.4732
R2358 VTAIL.n202 VTAIL.n201 10.4732
R2359 VTAIL.n263 VTAIL.n244 10.4732
R2360 VTAIL.n285 VTAIL.n234 10.4732
R2361 VTAIL.n310 VTAIL.n309 10.4732
R2362 VTAIL.n738 VTAIL.n737 10.4732
R2363 VTAIL.n713 VTAIL.n662 10.4732
R2364 VTAIL.n692 VTAIL.n673 10.4732
R2365 VTAIL.n630 VTAIL.n629 10.4732
R2366 VTAIL.n605 VTAIL.n554 10.4732
R2367 VTAIL.n584 VTAIL.n565 10.4732
R2368 VTAIL.n524 VTAIL.n523 10.4732
R2369 VTAIL.n499 VTAIL.n448 10.4732
R2370 VTAIL.n478 VTAIL.n459 10.4732
R2371 VTAIL.n416 VTAIL.n415 10.4732
R2372 VTAIL.n391 VTAIL.n340 10.4732
R2373 VTAIL.n370 VTAIL.n351 10.4732
R2374 VTAIL.n794 VTAIL.n793 9.69747
R2375 VTAIL.n820 VTAIL.n766 9.69747
R2376 VTAIL.n840 VTAIL.n756 9.69747
R2377 VTAIL.n46 VTAIL.n45 9.69747
R2378 VTAIL.n72 VTAIL.n18 9.69747
R2379 VTAIL.n92 VTAIL.n8 9.69747
R2380 VTAIL.n152 VTAIL.n151 9.69747
R2381 VTAIL.n178 VTAIL.n124 9.69747
R2382 VTAIL.n198 VTAIL.n114 9.69747
R2383 VTAIL.n260 VTAIL.n259 9.69747
R2384 VTAIL.n286 VTAIL.n232 9.69747
R2385 VTAIL.n306 VTAIL.n222 9.69747
R2386 VTAIL.n734 VTAIL.n650 9.69747
R2387 VTAIL.n714 VTAIL.n660 9.69747
R2388 VTAIL.n689 VTAIL.n688 9.69747
R2389 VTAIL.n626 VTAIL.n542 9.69747
R2390 VTAIL.n606 VTAIL.n552 9.69747
R2391 VTAIL.n581 VTAIL.n580 9.69747
R2392 VTAIL.n520 VTAIL.n436 9.69747
R2393 VTAIL.n500 VTAIL.n446 9.69747
R2394 VTAIL.n475 VTAIL.n474 9.69747
R2395 VTAIL.n412 VTAIL.n328 9.69747
R2396 VTAIL.n392 VTAIL.n338 9.69747
R2397 VTAIL.n367 VTAIL.n366 9.69747
R2398 VTAIL.n854 VTAIL.n853 9.45567
R2399 VTAIL.n106 VTAIL.n105 9.45567
R2400 VTAIL.n212 VTAIL.n211 9.45567
R2401 VTAIL.n320 VTAIL.n319 9.45567
R2402 VTAIL.n748 VTAIL.n747 9.45567
R2403 VTAIL.n640 VTAIL.n639 9.45567
R2404 VTAIL.n534 VTAIL.n533 9.45567
R2405 VTAIL.n426 VTAIL.n425 9.45567
R2406 VTAIL.n829 VTAIL.n828 9.3005
R2407 VTAIL.n764 VTAIL.n763 9.3005
R2408 VTAIL.n823 VTAIL.n822 9.3005
R2409 VTAIL.n821 VTAIL.n820 9.3005
R2410 VTAIL.n768 VTAIL.n767 9.3005
R2411 VTAIL.n815 VTAIL.n814 9.3005
R2412 VTAIL.n813 VTAIL.n812 9.3005
R2413 VTAIL.n772 VTAIL.n771 9.3005
R2414 VTAIL.n787 VTAIL.n786 9.3005
R2415 VTAIL.n789 VTAIL.n788 9.3005
R2416 VTAIL.n780 VTAIL.n779 9.3005
R2417 VTAIL.n795 VTAIL.n794 9.3005
R2418 VTAIL.n797 VTAIL.n796 9.3005
R2419 VTAIL.n776 VTAIL.n775 9.3005
R2420 VTAIL.n804 VTAIL.n803 9.3005
R2421 VTAIL.n806 VTAIL.n805 9.3005
R2422 VTAIL.n831 VTAIL.n830 9.3005
R2423 VTAIL.n760 VTAIL.n759 9.3005
R2424 VTAIL.n837 VTAIL.n836 9.3005
R2425 VTAIL.n839 VTAIL.n838 9.3005
R2426 VTAIL.n756 VTAIL.n755 9.3005
R2427 VTAIL.n845 VTAIL.n844 9.3005
R2428 VTAIL.n847 VTAIL.n846 9.3005
R2429 VTAIL.n752 VTAIL.n751 9.3005
R2430 VTAIL.n853 VTAIL.n852 9.3005
R2431 VTAIL.n81 VTAIL.n80 9.3005
R2432 VTAIL.n16 VTAIL.n15 9.3005
R2433 VTAIL.n75 VTAIL.n74 9.3005
R2434 VTAIL.n73 VTAIL.n72 9.3005
R2435 VTAIL.n20 VTAIL.n19 9.3005
R2436 VTAIL.n67 VTAIL.n66 9.3005
R2437 VTAIL.n65 VTAIL.n64 9.3005
R2438 VTAIL.n24 VTAIL.n23 9.3005
R2439 VTAIL.n39 VTAIL.n38 9.3005
R2440 VTAIL.n41 VTAIL.n40 9.3005
R2441 VTAIL.n32 VTAIL.n31 9.3005
R2442 VTAIL.n47 VTAIL.n46 9.3005
R2443 VTAIL.n49 VTAIL.n48 9.3005
R2444 VTAIL.n28 VTAIL.n27 9.3005
R2445 VTAIL.n56 VTAIL.n55 9.3005
R2446 VTAIL.n58 VTAIL.n57 9.3005
R2447 VTAIL.n83 VTAIL.n82 9.3005
R2448 VTAIL.n12 VTAIL.n11 9.3005
R2449 VTAIL.n89 VTAIL.n88 9.3005
R2450 VTAIL.n91 VTAIL.n90 9.3005
R2451 VTAIL.n8 VTAIL.n7 9.3005
R2452 VTAIL.n97 VTAIL.n96 9.3005
R2453 VTAIL.n99 VTAIL.n98 9.3005
R2454 VTAIL.n4 VTAIL.n3 9.3005
R2455 VTAIL.n105 VTAIL.n104 9.3005
R2456 VTAIL.n187 VTAIL.n186 9.3005
R2457 VTAIL.n122 VTAIL.n121 9.3005
R2458 VTAIL.n181 VTAIL.n180 9.3005
R2459 VTAIL.n179 VTAIL.n178 9.3005
R2460 VTAIL.n126 VTAIL.n125 9.3005
R2461 VTAIL.n173 VTAIL.n172 9.3005
R2462 VTAIL.n171 VTAIL.n170 9.3005
R2463 VTAIL.n130 VTAIL.n129 9.3005
R2464 VTAIL.n145 VTAIL.n144 9.3005
R2465 VTAIL.n147 VTAIL.n146 9.3005
R2466 VTAIL.n138 VTAIL.n137 9.3005
R2467 VTAIL.n153 VTAIL.n152 9.3005
R2468 VTAIL.n155 VTAIL.n154 9.3005
R2469 VTAIL.n134 VTAIL.n133 9.3005
R2470 VTAIL.n162 VTAIL.n161 9.3005
R2471 VTAIL.n164 VTAIL.n163 9.3005
R2472 VTAIL.n189 VTAIL.n188 9.3005
R2473 VTAIL.n118 VTAIL.n117 9.3005
R2474 VTAIL.n195 VTAIL.n194 9.3005
R2475 VTAIL.n197 VTAIL.n196 9.3005
R2476 VTAIL.n114 VTAIL.n113 9.3005
R2477 VTAIL.n203 VTAIL.n202 9.3005
R2478 VTAIL.n205 VTAIL.n204 9.3005
R2479 VTAIL.n110 VTAIL.n109 9.3005
R2480 VTAIL.n211 VTAIL.n210 9.3005
R2481 VTAIL.n295 VTAIL.n294 9.3005
R2482 VTAIL.n230 VTAIL.n229 9.3005
R2483 VTAIL.n289 VTAIL.n288 9.3005
R2484 VTAIL.n287 VTAIL.n286 9.3005
R2485 VTAIL.n234 VTAIL.n233 9.3005
R2486 VTAIL.n281 VTAIL.n280 9.3005
R2487 VTAIL.n279 VTAIL.n278 9.3005
R2488 VTAIL.n238 VTAIL.n237 9.3005
R2489 VTAIL.n253 VTAIL.n252 9.3005
R2490 VTAIL.n255 VTAIL.n254 9.3005
R2491 VTAIL.n246 VTAIL.n245 9.3005
R2492 VTAIL.n261 VTAIL.n260 9.3005
R2493 VTAIL.n263 VTAIL.n262 9.3005
R2494 VTAIL.n242 VTAIL.n241 9.3005
R2495 VTAIL.n270 VTAIL.n269 9.3005
R2496 VTAIL.n272 VTAIL.n271 9.3005
R2497 VTAIL.n297 VTAIL.n296 9.3005
R2498 VTAIL.n226 VTAIL.n225 9.3005
R2499 VTAIL.n303 VTAIL.n302 9.3005
R2500 VTAIL.n305 VTAIL.n304 9.3005
R2501 VTAIL.n222 VTAIL.n221 9.3005
R2502 VTAIL.n311 VTAIL.n310 9.3005
R2503 VTAIL.n313 VTAIL.n312 9.3005
R2504 VTAIL.n218 VTAIL.n217 9.3005
R2505 VTAIL.n319 VTAIL.n318 9.3005
R2506 VTAIL.n682 VTAIL.n681 9.3005
R2507 VTAIL.n684 VTAIL.n683 9.3005
R2508 VTAIL.n675 VTAIL.n674 9.3005
R2509 VTAIL.n690 VTAIL.n689 9.3005
R2510 VTAIL.n692 VTAIL.n691 9.3005
R2511 VTAIL.n670 VTAIL.n669 9.3005
R2512 VTAIL.n698 VTAIL.n697 9.3005
R2513 VTAIL.n700 VTAIL.n699 9.3005
R2514 VTAIL.n654 VTAIL.n653 9.3005
R2515 VTAIL.n731 VTAIL.n730 9.3005
R2516 VTAIL.n733 VTAIL.n732 9.3005
R2517 VTAIL.n650 VTAIL.n649 9.3005
R2518 VTAIL.n739 VTAIL.n738 9.3005
R2519 VTAIL.n741 VTAIL.n740 9.3005
R2520 VTAIL.n646 VTAIL.n645 9.3005
R2521 VTAIL.n747 VTAIL.n746 9.3005
R2522 VTAIL.n725 VTAIL.n724 9.3005
R2523 VTAIL.n723 VTAIL.n722 9.3005
R2524 VTAIL.n658 VTAIL.n657 9.3005
R2525 VTAIL.n717 VTAIL.n716 9.3005
R2526 VTAIL.n715 VTAIL.n714 9.3005
R2527 VTAIL.n662 VTAIL.n661 9.3005
R2528 VTAIL.n709 VTAIL.n708 9.3005
R2529 VTAIL.n707 VTAIL.n706 9.3005
R2530 VTAIL.n666 VTAIL.n665 9.3005
R2531 VTAIL.n574 VTAIL.n573 9.3005
R2532 VTAIL.n576 VTAIL.n575 9.3005
R2533 VTAIL.n567 VTAIL.n566 9.3005
R2534 VTAIL.n582 VTAIL.n581 9.3005
R2535 VTAIL.n584 VTAIL.n583 9.3005
R2536 VTAIL.n562 VTAIL.n561 9.3005
R2537 VTAIL.n590 VTAIL.n589 9.3005
R2538 VTAIL.n592 VTAIL.n591 9.3005
R2539 VTAIL.n546 VTAIL.n545 9.3005
R2540 VTAIL.n623 VTAIL.n622 9.3005
R2541 VTAIL.n625 VTAIL.n624 9.3005
R2542 VTAIL.n542 VTAIL.n541 9.3005
R2543 VTAIL.n631 VTAIL.n630 9.3005
R2544 VTAIL.n633 VTAIL.n632 9.3005
R2545 VTAIL.n538 VTAIL.n537 9.3005
R2546 VTAIL.n639 VTAIL.n638 9.3005
R2547 VTAIL.n617 VTAIL.n616 9.3005
R2548 VTAIL.n615 VTAIL.n614 9.3005
R2549 VTAIL.n550 VTAIL.n549 9.3005
R2550 VTAIL.n609 VTAIL.n608 9.3005
R2551 VTAIL.n607 VTAIL.n606 9.3005
R2552 VTAIL.n554 VTAIL.n553 9.3005
R2553 VTAIL.n601 VTAIL.n600 9.3005
R2554 VTAIL.n599 VTAIL.n598 9.3005
R2555 VTAIL.n558 VTAIL.n557 9.3005
R2556 VTAIL.n468 VTAIL.n467 9.3005
R2557 VTAIL.n470 VTAIL.n469 9.3005
R2558 VTAIL.n461 VTAIL.n460 9.3005
R2559 VTAIL.n476 VTAIL.n475 9.3005
R2560 VTAIL.n478 VTAIL.n477 9.3005
R2561 VTAIL.n456 VTAIL.n455 9.3005
R2562 VTAIL.n484 VTAIL.n483 9.3005
R2563 VTAIL.n486 VTAIL.n485 9.3005
R2564 VTAIL.n440 VTAIL.n439 9.3005
R2565 VTAIL.n517 VTAIL.n516 9.3005
R2566 VTAIL.n519 VTAIL.n518 9.3005
R2567 VTAIL.n436 VTAIL.n435 9.3005
R2568 VTAIL.n525 VTAIL.n524 9.3005
R2569 VTAIL.n527 VTAIL.n526 9.3005
R2570 VTAIL.n432 VTAIL.n431 9.3005
R2571 VTAIL.n533 VTAIL.n532 9.3005
R2572 VTAIL.n511 VTAIL.n510 9.3005
R2573 VTAIL.n509 VTAIL.n508 9.3005
R2574 VTAIL.n444 VTAIL.n443 9.3005
R2575 VTAIL.n503 VTAIL.n502 9.3005
R2576 VTAIL.n501 VTAIL.n500 9.3005
R2577 VTAIL.n448 VTAIL.n447 9.3005
R2578 VTAIL.n495 VTAIL.n494 9.3005
R2579 VTAIL.n493 VTAIL.n492 9.3005
R2580 VTAIL.n452 VTAIL.n451 9.3005
R2581 VTAIL.n360 VTAIL.n359 9.3005
R2582 VTAIL.n362 VTAIL.n361 9.3005
R2583 VTAIL.n353 VTAIL.n352 9.3005
R2584 VTAIL.n368 VTAIL.n367 9.3005
R2585 VTAIL.n370 VTAIL.n369 9.3005
R2586 VTAIL.n348 VTAIL.n347 9.3005
R2587 VTAIL.n376 VTAIL.n375 9.3005
R2588 VTAIL.n378 VTAIL.n377 9.3005
R2589 VTAIL.n332 VTAIL.n331 9.3005
R2590 VTAIL.n409 VTAIL.n408 9.3005
R2591 VTAIL.n411 VTAIL.n410 9.3005
R2592 VTAIL.n328 VTAIL.n327 9.3005
R2593 VTAIL.n417 VTAIL.n416 9.3005
R2594 VTAIL.n419 VTAIL.n418 9.3005
R2595 VTAIL.n324 VTAIL.n323 9.3005
R2596 VTAIL.n425 VTAIL.n424 9.3005
R2597 VTAIL.n403 VTAIL.n402 9.3005
R2598 VTAIL.n401 VTAIL.n400 9.3005
R2599 VTAIL.n336 VTAIL.n335 9.3005
R2600 VTAIL.n395 VTAIL.n394 9.3005
R2601 VTAIL.n393 VTAIL.n392 9.3005
R2602 VTAIL.n340 VTAIL.n339 9.3005
R2603 VTAIL.n387 VTAIL.n386 9.3005
R2604 VTAIL.n385 VTAIL.n384 9.3005
R2605 VTAIL.n344 VTAIL.n343 9.3005
R2606 VTAIL.n790 VTAIL.n780 8.92171
R2607 VTAIL.n824 VTAIL.n823 8.92171
R2608 VTAIL.n839 VTAIL.n758 8.92171
R2609 VTAIL.n42 VTAIL.n32 8.92171
R2610 VTAIL.n76 VTAIL.n75 8.92171
R2611 VTAIL.n91 VTAIL.n10 8.92171
R2612 VTAIL.n148 VTAIL.n138 8.92171
R2613 VTAIL.n182 VTAIL.n181 8.92171
R2614 VTAIL.n197 VTAIL.n116 8.92171
R2615 VTAIL.n256 VTAIL.n246 8.92171
R2616 VTAIL.n290 VTAIL.n289 8.92171
R2617 VTAIL.n305 VTAIL.n224 8.92171
R2618 VTAIL.n733 VTAIL.n652 8.92171
R2619 VTAIL.n718 VTAIL.n717 8.92171
R2620 VTAIL.n685 VTAIL.n675 8.92171
R2621 VTAIL.n625 VTAIL.n544 8.92171
R2622 VTAIL.n610 VTAIL.n609 8.92171
R2623 VTAIL.n577 VTAIL.n567 8.92171
R2624 VTAIL.n519 VTAIL.n438 8.92171
R2625 VTAIL.n504 VTAIL.n503 8.92171
R2626 VTAIL.n471 VTAIL.n461 8.92171
R2627 VTAIL.n411 VTAIL.n330 8.92171
R2628 VTAIL.n396 VTAIL.n395 8.92171
R2629 VTAIL.n363 VTAIL.n353 8.92171
R2630 VTAIL.n789 VTAIL.n782 8.14595
R2631 VTAIL.n827 VTAIL.n764 8.14595
R2632 VTAIL.n836 VTAIL.n835 8.14595
R2633 VTAIL.n41 VTAIL.n34 8.14595
R2634 VTAIL.n79 VTAIL.n16 8.14595
R2635 VTAIL.n88 VTAIL.n87 8.14595
R2636 VTAIL.n147 VTAIL.n140 8.14595
R2637 VTAIL.n185 VTAIL.n122 8.14595
R2638 VTAIL.n194 VTAIL.n193 8.14595
R2639 VTAIL.n255 VTAIL.n248 8.14595
R2640 VTAIL.n293 VTAIL.n230 8.14595
R2641 VTAIL.n302 VTAIL.n301 8.14595
R2642 VTAIL.n730 VTAIL.n729 8.14595
R2643 VTAIL.n721 VTAIL.n658 8.14595
R2644 VTAIL.n684 VTAIL.n677 8.14595
R2645 VTAIL.n622 VTAIL.n621 8.14595
R2646 VTAIL.n613 VTAIL.n550 8.14595
R2647 VTAIL.n576 VTAIL.n569 8.14595
R2648 VTAIL.n516 VTAIL.n515 8.14595
R2649 VTAIL.n507 VTAIL.n444 8.14595
R2650 VTAIL.n470 VTAIL.n463 8.14595
R2651 VTAIL.n408 VTAIL.n407 8.14595
R2652 VTAIL.n399 VTAIL.n336 8.14595
R2653 VTAIL.n362 VTAIL.n355 8.14595
R2654 VTAIL.n854 VTAIL.n750 7.75445
R2655 VTAIL.n106 VTAIL.n2 7.75445
R2656 VTAIL.n212 VTAIL.n108 7.75445
R2657 VTAIL.n320 VTAIL.n216 7.75445
R2658 VTAIL.n748 VTAIL.n644 7.75445
R2659 VTAIL.n640 VTAIL.n536 7.75445
R2660 VTAIL.n534 VTAIL.n430 7.75445
R2661 VTAIL.n426 VTAIL.n322 7.75445
R2662 VTAIL.n786 VTAIL.n785 7.3702
R2663 VTAIL.n828 VTAIL.n762 7.3702
R2664 VTAIL.n832 VTAIL.n760 7.3702
R2665 VTAIL.n38 VTAIL.n37 7.3702
R2666 VTAIL.n80 VTAIL.n14 7.3702
R2667 VTAIL.n84 VTAIL.n12 7.3702
R2668 VTAIL.n144 VTAIL.n143 7.3702
R2669 VTAIL.n186 VTAIL.n120 7.3702
R2670 VTAIL.n190 VTAIL.n118 7.3702
R2671 VTAIL.n252 VTAIL.n251 7.3702
R2672 VTAIL.n294 VTAIL.n228 7.3702
R2673 VTAIL.n298 VTAIL.n226 7.3702
R2674 VTAIL.n726 VTAIL.n654 7.3702
R2675 VTAIL.n722 VTAIL.n656 7.3702
R2676 VTAIL.n681 VTAIL.n680 7.3702
R2677 VTAIL.n618 VTAIL.n546 7.3702
R2678 VTAIL.n614 VTAIL.n548 7.3702
R2679 VTAIL.n573 VTAIL.n572 7.3702
R2680 VTAIL.n512 VTAIL.n440 7.3702
R2681 VTAIL.n508 VTAIL.n442 7.3702
R2682 VTAIL.n467 VTAIL.n466 7.3702
R2683 VTAIL.n404 VTAIL.n332 7.3702
R2684 VTAIL.n400 VTAIL.n334 7.3702
R2685 VTAIL.n359 VTAIL.n358 7.3702
R2686 VTAIL.n831 VTAIL.n762 6.59444
R2687 VTAIL.n832 VTAIL.n831 6.59444
R2688 VTAIL.n83 VTAIL.n14 6.59444
R2689 VTAIL.n84 VTAIL.n83 6.59444
R2690 VTAIL.n189 VTAIL.n120 6.59444
R2691 VTAIL.n190 VTAIL.n189 6.59444
R2692 VTAIL.n297 VTAIL.n228 6.59444
R2693 VTAIL.n298 VTAIL.n297 6.59444
R2694 VTAIL.n726 VTAIL.n725 6.59444
R2695 VTAIL.n725 VTAIL.n656 6.59444
R2696 VTAIL.n618 VTAIL.n617 6.59444
R2697 VTAIL.n617 VTAIL.n548 6.59444
R2698 VTAIL.n512 VTAIL.n511 6.59444
R2699 VTAIL.n511 VTAIL.n442 6.59444
R2700 VTAIL.n404 VTAIL.n403 6.59444
R2701 VTAIL.n403 VTAIL.n334 6.59444
R2702 VTAIL.n852 VTAIL.n750 6.08283
R2703 VTAIL.n104 VTAIL.n2 6.08283
R2704 VTAIL.n210 VTAIL.n108 6.08283
R2705 VTAIL.n318 VTAIL.n216 6.08283
R2706 VTAIL.n746 VTAIL.n644 6.08283
R2707 VTAIL.n638 VTAIL.n536 6.08283
R2708 VTAIL.n532 VTAIL.n430 6.08283
R2709 VTAIL.n424 VTAIL.n322 6.08283
R2710 VTAIL.n786 VTAIL.n782 5.81868
R2711 VTAIL.n828 VTAIL.n827 5.81868
R2712 VTAIL.n835 VTAIL.n760 5.81868
R2713 VTAIL.n38 VTAIL.n34 5.81868
R2714 VTAIL.n80 VTAIL.n79 5.81868
R2715 VTAIL.n87 VTAIL.n12 5.81868
R2716 VTAIL.n144 VTAIL.n140 5.81868
R2717 VTAIL.n186 VTAIL.n185 5.81868
R2718 VTAIL.n193 VTAIL.n118 5.81868
R2719 VTAIL.n252 VTAIL.n248 5.81868
R2720 VTAIL.n294 VTAIL.n293 5.81868
R2721 VTAIL.n301 VTAIL.n226 5.81868
R2722 VTAIL.n729 VTAIL.n654 5.81868
R2723 VTAIL.n722 VTAIL.n721 5.81868
R2724 VTAIL.n681 VTAIL.n677 5.81868
R2725 VTAIL.n621 VTAIL.n546 5.81868
R2726 VTAIL.n614 VTAIL.n613 5.81868
R2727 VTAIL.n573 VTAIL.n569 5.81868
R2728 VTAIL.n515 VTAIL.n440 5.81868
R2729 VTAIL.n508 VTAIL.n507 5.81868
R2730 VTAIL.n467 VTAIL.n463 5.81868
R2731 VTAIL.n407 VTAIL.n332 5.81868
R2732 VTAIL.n400 VTAIL.n399 5.81868
R2733 VTAIL.n359 VTAIL.n355 5.81868
R2734 VTAIL.n790 VTAIL.n789 5.04292
R2735 VTAIL.n824 VTAIL.n764 5.04292
R2736 VTAIL.n836 VTAIL.n758 5.04292
R2737 VTAIL.n42 VTAIL.n41 5.04292
R2738 VTAIL.n76 VTAIL.n16 5.04292
R2739 VTAIL.n88 VTAIL.n10 5.04292
R2740 VTAIL.n148 VTAIL.n147 5.04292
R2741 VTAIL.n182 VTAIL.n122 5.04292
R2742 VTAIL.n194 VTAIL.n116 5.04292
R2743 VTAIL.n256 VTAIL.n255 5.04292
R2744 VTAIL.n290 VTAIL.n230 5.04292
R2745 VTAIL.n302 VTAIL.n224 5.04292
R2746 VTAIL.n730 VTAIL.n652 5.04292
R2747 VTAIL.n718 VTAIL.n658 5.04292
R2748 VTAIL.n685 VTAIL.n684 5.04292
R2749 VTAIL.n622 VTAIL.n544 5.04292
R2750 VTAIL.n610 VTAIL.n550 5.04292
R2751 VTAIL.n577 VTAIL.n576 5.04292
R2752 VTAIL.n516 VTAIL.n438 5.04292
R2753 VTAIL.n504 VTAIL.n444 5.04292
R2754 VTAIL.n471 VTAIL.n470 5.04292
R2755 VTAIL.n408 VTAIL.n330 5.04292
R2756 VTAIL.n396 VTAIL.n336 5.04292
R2757 VTAIL.n363 VTAIL.n362 5.04292
R2758 VTAIL.n793 VTAIL.n780 4.26717
R2759 VTAIL.n823 VTAIL.n766 4.26717
R2760 VTAIL.n840 VTAIL.n839 4.26717
R2761 VTAIL.n45 VTAIL.n32 4.26717
R2762 VTAIL.n75 VTAIL.n18 4.26717
R2763 VTAIL.n92 VTAIL.n91 4.26717
R2764 VTAIL.n151 VTAIL.n138 4.26717
R2765 VTAIL.n181 VTAIL.n124 4.26717
R2766 VTAIL.n198 VTAIL.n197 4.26717
R2767 VTAIL.n259 VTAIL.n246 4.26717
R2768 VTAIL.n289 VTAIL.n232 4.26717
R2769 VTAIL.n306 VTAIL.n305 4.26717
R2770 VTAIL.n734 VTAIL.n733 4.26717
R2771 VTAIL.n717 VTAIL.n660 4.26717
R2772 VTAIL.n688 VTAIL.n675 4.26717
R2773 VTAIL.n626 VTAIL.n625 4.26717
R2774 VTAIL.n609 VTAIL.n552 4.26717
R2775 VTAIL.n580 VTAIL.n567 4.26717
R2776 VTAIL.n520 VTAIL.n519 4.26717
R2777 VTAIL.n503 VTAIL.n446 4.26717
R2778 VTAIL.n474 VTAIL.n461 4.26717
R2779 VTAIL.n412 VTAIL.n411 4.26717
R2780 VTAIL.n395 VTAIL.n338 4.26717
R2781 VTAIL.n366 VTAIL.n353 4.26717
R2782 VTAIL.n429 VTAIL.n427 3.5005
R2783 VTAIL.n535 VTAIL.n429 3.5005
R2784 VTAIL.n643 VTAIL.n641 3.5005
R2785 VTAIL.n749 VTAIL.n643 3.5005
R2786 VTAIL.n321 VTAIL.n215 3.5005
R2787 VTAIL.n215 VTAIL.n213 3.5005
R2788 VTAIL.n107 VTAIL.n1 3.5005
R2789 VTAIL.n794 VTAIL.n778 3.49141
R2790 VTAIL.n820 VTAIL.n819 3.49141
R2791 VTAIL.n843 VTAIL.n756 3.49141
R2792 VTAIL.n46 VTAIL.n30 3.49141
R2793 VTAIL.n72 VTAIL.n71 3.49141
R2794 VTAIL.n95 VTAIL.n8 3.49141
R2795 VTAIL.n152 VTAIL.n136 3.49141
R2796 VTAIL.n178 VTAIL.n177 3.49141
R2797 VTAIL.n201 VTAIL.n114 3.49141
R2798 VTAIL.n260 VTAIL.n244 3.49141
R2799 VTAIL.n286 VTAIL.n285 3.49141
R2800 VTAIL.n309 VTAIL.n222 3.49141
R2801 VTAIL.n737 VTAIL.n650 3.49141
R2802 VTAIL.n714 VTAIL.n713 3.49141
R2803 VTAIL.n689 VTAIL.n673 3.49141
R2804 VTAIL.n629 VTAIL.n542 3.49141
R2805 VTAIL.n606 VTAIL.n605 3.49141
R2806 VTAIL.n581 VTAIL.n565 3.49141
R2807 VTAIL.n523 VTAIL.n436 3.49141
R2808 VTAIL.n500 VTAIL.n499 3.49141
R2809 VTAIL.n475 VTAIL.n459 3.49141
R2810 VTAIL.n415 VTAIL.n328 3.49141
R2811 VTAIL.n392 VTAIL.n391 3.49141
R2812 VTAIL.n367 VTAIL.n351 3.49141
R2813 VTAIL VTAIL.n855 3.44231
R2814 VTAIL.n798 VTAIL.n797 2.71565
R2815 VTAIL.n816 VTAIL.n768 2.71565
R2816 VTAIL.n844 VTAIL.n754 2.71565
R2817 VTAIL.n50 VTAIL.n49 2.71565
R2818 VTAIL.n68 VTAIL.n20 2.71565
R2819 VTAIL.n96 VTAIL.n6 2.71565
R2820 VTAIL.n156 VTAIL.n155 2.71565
R2821 VTAIL.n174 VTAIL.n126 2.71565
R2822 VTAIL.n202 VTAIL.n112 2.71565
R2823 VTAIL.n264 VTAIL.n263 2.71565
R2824 VTAIL.n282 VTAIL.n234 2.71565
R2825 VTAIL.n310 VTAIL.n220 2.71565
R2826 VTAIL.n738 VTAIL.n648 2.71565
R2827 VTAIL.n710 VTAIL.n662 2.71565
R2828 VTAIL.n693 VTAIL.n692 2.71565
R2829 VTAIL.n630 VTAIL.n540 2.71565
R2830 VTAIL.n602 VTAIL.n554 2.71565
R2831 VTAIL.n585 VTAIL.n584 2.71565
R2832 VTAIL.n524 VTAIL.n434 2.71565
R2833 VTAIL.n496 VTAIL.n448 2.71565
R2834 VTAIL.n479 VTAIL.n478 2.71565
R2835 VTAIL.n416 VTAIL.n326 2.71565
R2836 VTAIL.n388 VTAIL.n340 2.71565
R2837 VTAIL.n371 VTAIL.n370 2.71565
R2838 VTAIL.n682 VTAIL.n678 2.41282
R2839 VTAIL.n574 VTAIL.n570 2.41282
R2840 VTAIL.n468 VTAIL.n464 2.41282
R2841 VTAIL.n360 VTAIL.n356 2.41282
R2842 VTAIL.n787 VTAIL.n783 2.41282
R2843 VTAIL.n39 VTAIL.n35 2.41282
R2844 VTAIL.n145 VTAIL.n141 2.41282
R2845 VTAIL.n253 VTAIL.n249 2.41282
R2846 VTAIL.n802 VTAIL.n776 1.93989
R2847 VTAIL.n815 VTAIL.n770 1.93989
R2848 VTAIL.n848 VTAIL.n847 1.93989
R2849 VTAIL.n54 VTAIL.n28 1.93989
R2850 VTAIL.n67 VTAIL.n22 1.93989
R2851 VTAIL.n100 VTAIL.n99 1.93989
R2852 VTAIL.n160 VTAIL.n134 1.93989
R2853 VTAIL.n173 VTAIL.n128 1.93989
R2854 VTAIL.n206 VTAIL.n205 1.93989
R2855 VTAIL.n268 VTAIL.n242 1.93989
R2856 VTAIL.n281 VTAIL.n236 1.93989
R2857 VTAIL.n314 VTAIL.n313 1.93989
R2858 VTAIL.n742 VTAIL.n741 1.93989
R2859 VTAIL.n709 VTAIL.n664 1.93989
R2860 VTAIL.n696 VTAIL.n670 1.93989
R2861 VTAIL.n634 VTAIL.n633 1.93989
R2862 VTAIL.n601 VTAIL.n556 1.93989
R2863 VTAIL.n588 VTAIL.n562 1.93989
R2864 VTAIL.n528 VTAIL.n527 1.93989
R2865 VTAIL.n495 VTAIL.n450 1.93989
R2866 VTAIL.n482 VTAIL.n456 1.93989
R2867 VTAIL.n420 VTAIL.n419 1.93989
R2868 VTAIL.n387 VTAIL.n342 1.93989
R2869 VTAIL.n374 VTAIL.n348 1.93989
R2870 VTAIL.n0 VTAIL.t2 1.67257
R2871 VTAIL.n0 VTAIL.t15 1.67257
R2872 VTAIL.n214 VTAIL.t10 1.67257
R2873 VTAIL.n214 VTAIL.t4 1.67257
R2874 VTAIL.n642 VTAIL.t6 1.67257
R2875 VTAIL.n642 VTAIL.t7 1.67257
R2876 VTAIL.n428 VTAIL.t0 1.67257
R2877 VTAIL.n428 VTAIL.t12 1.67257
R2878 VTAIL.n803 VTAIL.n774 1.16414
R2879 VTAIL.n812 VTAIL.n811 1.16414
R2880 VTAIL.n851 VTAIL.n752 1.16414
R2881 VTAIL.n55 VTAIL.n26 1.16414
R2882 VTAIL.n64 VTAIL.n63 1.16414
R2883 VTAIL.n103 VTAIL.n4 1.16414
R2884 VTAIL.n161 VTAIL.n132 1.16414
R2885 VTAIL.n170 VTAIL.n169 1.16414
R2886 VTAIL.n209 VTAIL.n110 1.16414
R2887 VTAIL.n269 VTAIL.n240 1.16414
R2888 VTAIL.n278 VTAIL.n277 1.16414
R2889 VTAIL.n317 VTAIL.n218 1.16414
R2890 VTAIL.n745 VTAIL.n646 1.16414
R2891 VTAIL.n706 VTAIL.n705 1.16414
R2892 VTAIL.n697 VTAIL.n668 1.16414
R2893 VTAIL.n637 VTAIL.n538 1.16414
R2894 VTAIL.n598 VTAIL.n597 1.16414
R2895 VTAIL.n589 VTAIL.n560 1.16414
R2896 VTAIL.n531 VTAIL.n432 1.16414
R2897 VTAIL.n492 VTAIL.n491 1.16414
R2898 VTAIL.n483 VTAIL.n454 1.16414
R2899 VTAIL.n423 VTAIL.n324 1.16414
R2900 VTAIL.n384 VTAIL.n383 1.16414
R2901 VTAIL.n375 VTAIL.n346 1.16414
R2902 VTAIL.n641 VTAIL.n535 0.470328
R2903 VTAIL.n213 VTAIL.n107 0.470328
R2904 VTAIL.n807 VTAIL.n806 0.388379
R2905 VTAIL.n808 VTAIL.n772 0.388379
R2906 VTAIL.n59 VTAIL.n58 0.388379
R2907 VTAIL.n60 VTAIL.n24 0.388379
R2908 VTAIL.n165 VTAIL.n164 0.388379
R2909 VTAIL.n166 VTAIL.n130 0.388379
R2910 VTAIL.n273 VTAIL.n272 0.388379
R2911 VTAIL.n274 VTAIL.n238 0.388379
R2912 VTAIL.n702 VTAIL.n666 0.388379
R2913 VTAIL.n701 VTAIL.n700 0.388379
R2914 VTAIL.n594 VTAIL.n558 0.388379
R2915 VTAIL.n593 VTAIL.n592 0.388379
R2916 VTAIL.n488 VTAIL.n452 0.388379
R2917 VTAIL.n487 VTAIL.n486 0.388379
R2918 VTAIL.n380 VTAIL.n344 0.388379
R2919 VTAIL.n379 VTAIL.n378 0.388379
R2920 VTAIL.n788 VTAIL.n787 0.155672
R2921 VTAIL.n788 VTAIL.n779 0.155672
R2922 VTAIL.n795 VTAIL.n779 0.155672
R2923 VTAIL.n796 VTAIL.n795 0.155672
R2924 VTAIL.n796 VTAIL.n775 0.155672
R2925 VTAIL.n804 VTAIL.n775 0.155672
R2926 VTAIL.n805 VTAIL.n804 0.155672
R2927 VTAIL.n805 VTAIL.n771 0.155672
R2928 VTAIL.n813 VTAIL.n771 0.155672
R2929 VTAIL.n814 VTAIL.n813 0.155672
R2930 VTAIL.n814 VTAIL.n767 0.155672
R2931 VTAIL.n821 VTAIL.n767 0.155672
R2932 VTAIL.n822 VTAIL.n821 0.155672
R2933 VTAIL.n822 VTAIL.n763 0.155672
R2934 VTAIL.n829 VTAIL.n763 0.155672
R2935 VTAIL.n830 VTAIL.n829 0.155672
R2936 VTAIL.n830 VTAIL.n759 0.155672
R2937 VTAIL.n837 VTAIL.n759 0.155672
R2938 VTAIL.n838 VTAIL.n837 0.155672
R2939 VTAIL.n838 VTAIL.n755 0.155672
R2940 VTAIL.n845 VTAIL.n755 0.155672
R2941 VTAIL.n846 VTAIL.n845 0.155672
R2942 VTAIL.n846 VTAIL.n751 0.155672
R2943 VTAIL.n853 VTAIL.n751 0.155672
R2944 VTAIL.n40 VTAIL.n39 0.155672
R2945 VTAIL.n40 VTAIL.n31 0.155672
R2946 VTAIL.n47 VTAIL.n31 0.155672
R2947 VTAIL.n48 VTAIL.n47 0.155672
R2948 VTAIL.n48 VTAIL.n27 0.155672
R2949 VTAIL.n56 VTAIL.n27 0.155672
R2950 VTAIL.n57 VTAIL.n56 0.155672
R2951 VTAIL.n57 VTAIL.n23 0.155672
R2952 VTAIL.n65 VTAIL.n23 0.155672
R2953 VTAIL.n66 VTAIL.n65 0.155672
R2954 VTAIL.n66 VTAIL.n19 0.155672
R2955 VTAIL.n73 VTAIL.n19 0.155672
R2956 VTAIL.n74 VTAIL.n73 0.155672
R2957 VTAIL.n74 VTAIL.n15 0.155672
R2958 VTAIL.n81 VTAIL.n15 0.155672
R2959 VTAIL.n82 VTAIL.n81 0.155672
R2960 VTAIL.n82 VTAIL.n11 0.155672
R2961 VTAIL.n89 VTAIL.n11 0.155672
R2962 VTAIL.n90 VTAIL.n89 0.155672
R2963 VTAIL.n90 VTAIL.n7 0.155672
R2964 VTAIL.n97 VTAIL.n7 0.155672
R2965 VTAIL.n98 VTAIL.n97 0.155672
R2966 VTAIL.n98 VTAIL.n3 0.155672
R2967 VTAIL.n105 VTAIL.n3 0.155672
R2968 VTAIL.n146 VTAIL.n145 0.155672
R2969 VTAIL.n146 VTAIL.n137 0.155672
R2970 VTAIL.n153 VTAIL.n137 0.155672
R2971 VTAIL.n154 VTAIL.n153 0.155672
R2972 VTAIL.n154 VTAIL.n133 0.155672
R2973 VTAIL.n162 VTAIL.n133 0.155672
R2974 VTAIL.n163 VTAIL.n162 0.155672
R2975 VTAIL.n163 VTAIL.n129 0.155672
R2976 VTAIL.n171 VTAIL.n129 0.155672
R2977 VTAIL.n172 VTAIL.n171 0.155672
R2978 VTAIL.n172 VTAIL.n125 0.155672
R2979 VTAIL.n179 VTAIL.n125 0.155672
R2980 VTAIL.n180 VTAIL.n179 0.155672
R2981 VTAIL.n180 VTAIL.n121 0.155672
R2982 VTAIL.n187 VTAIL.n121 0.155672
R2983 VTAIL.n188 VTAIL.n187 0.155672
R2984 VTAIL.n188 VTAIL.n117 0.155672
R2985 VTAIL.n195 VTAIL.n117 0.155672
R2986 VTAIL.n196 VTAIL.n195 0.155672
R2987 VTAIL.n196 VTAIL.n113 0.155672
R2988 VTAIL.n203 VTAIL.n113 0.155672
R2989 VTAIL.n204 VTAIL.n203 0.155672
R2990 VTAIL.n204 VTAIL.n109 0.155672
R2991 VTAIL.n211 VTAIL.n109 0.155672
R2992 VTAIL.n254 VTAIL.n253 0.155672
R2993 VTAIL.n254 VTAIL.n245 0.155672
R2994 VTAIL.n261 VTAIL.n245 0.155672
R2995 VTAIL.n262 VTAIL.n261 0.155672
R2996 VTAIL.n262 VTAIL.n241 0.155672
R2997 VTAIL.n270 VTAIL.n241 0.155672
R2998 VTAIL.n271 VTAIL.n270 0.155672
R2999 VTAIL.n271 VTAIL.n237 0.155672
R3000 VTAIL.n279 VTAIL.n237 0.155672
R3001 VTAIL.n280 VTAIL.n279 0.155672
R3002 VTAIL.n280 VTAIL.n233 0.155672
R3003 VTAIL.n287 VTAIL.n233 0.155672
R3004 VTAIL.n288 VTAIL.n287 0.155672
R3005 VTAIL.n288 VTAIL.n229 0.155672
R3006 VTAIL.n295 VTAIL.n229 0.155672
R3007 VTAIL.n296 VTAIL.n295 0.155672
R3008 VTAIL.n296 VTAIL.n225 0.155672
R3009 VTAIL.n303 VTAIL.n225 0.155672
R3010 VTAIL.n304 VTAIL.n303 0.155672
R3011 VTAIL.n304 VTAIL.n221 0.155672
R3012 VTAIL.n311 VTAIL.n221 0.155672
R3013 VTAIL.n312 VTAIL.n311 0.155672
R3014 VTAIL.n312 VTAIL.n217 0.155672
R3015 VTAIL.n319 VTAIL.n217 0.155672
R3016 VTAIL.n747 VTAIL.n645 0.155672
R3017 VTAIL.n740 VTAIL.n645 0.155672
R3018 VTAIL.n740 VTAIL.n739 0.155672
R3019 VTAIL.n739 VTAIL.n649 0.155672
R3020 VTAIL.n732 VTAIL.n649 0.155672
R3021 VTAIL.n732 VTAIL.n731 0.155672
R3022 VTAIL.n731 VTAIL.n653 0.155672
R3023 VTAIL.n724 VTAIL.n653 0.155672
R3024 VTAIL.n724 VTAIL.n723 0.155672
R3025 VTAIL.n723 VTAIL.n657 0.155672
R3026 VTAIL.n716 VTAIL.n657 0.155672
R3027 VTAIL.n716 VTAIL.n715 0.155672
R3028 VTAIL.n715 VTAIL.n661 0.155672
R3029 VTAIL.n708 VTAIL.n661 0.155672
R3030 VTAIL.n708 VTAIL.n707 0.155672
R3031 VTAIL.n707 VTAIL.n665 0.155672
R3032 VTAIL.n699 VTAIL.n665 0.155672
R3033 VTAIL.n699 VTAIL.n698 0.155672
R3034 VTAIL.n698 VTAIL.n669 0.155672
R3035 VTAIL.n691 VTAIL.n669 0.155672
R3036 VTAIL.n691 VTAIL.n690 0.155672
R3037 VTAIL.n690 VTAIL.n674 0.155672
R3038 VTAIL.n683 VTAIL.n674 0.155672
R3039 VTAIL.n683 VTAIL.n682 0.155672
R3040 VTAIL.n639 VTAIL.n537 0.155672
R3041 VTAIL.n632 VTAIL.n537 0.155672
R3042 VTAIL.n632 VTAIL.n631 0.155672
R3043 VTAIL.n631 VTAIL.n541 0.155672
R3044 VTAIL.n624 VTAIL.n541 0.155672
R3045 VTAIL.n624 VTAIL.n623 0.155672
R3046 VTAIL.n623 VTAIL.n545 0.155672
R3047 VTAIL.n616 VTAIL.n545 0.155672
R3048 VTAIL.n616 VTAIL.n615 0.155672
R3049 VTAIL.n615 VTAIL.n549 0.155672
R3050 VTAIL.n608 VTAIL.n549 0.155672
R3051 VTAIL.n608 VTAIL.n607 0.155672
R3052 VTAIL.n607 VTAIL.n553 0.155672
R3053 VTAIL.n600 VTAIL.n553 0.155672
R3054 VTAIL.n600 VTAIL.n599 0.155672
R3055 VTAIL.n599 VTAIL.n557 0.155672
R3056 VTAIL.n591 VTAIL.n557 0.155672
R3057 VTAIL.n591 VTAIL.n590 0.155672
R3058 VTAIL.n590 VTAIL.n561 0.155672
R3059 VTAIL.n583 VTAIL.n561 0.155672
R3060 VTAIL.n583 VTAIL.n582 0.155672
R3061 VTAIL.n582 VTAIL.n566 0.155672
R3062 VTAIL.n575 VTAIL.n566 0.155672
R3063 VTAIL.n575 VTAIL.n574 0.155672
R3064 VTAIL.n533 VTAIL.n431 0.155672
R3065 VTAIL.n526 VTAIL.n431 0.155672
R3066 VTAIL.n526 VTAIL.n525 0.155672
R3067 VTAIL.n525 VTAIL.n435 0.155672
R3068 VTAIL.n518 VTAIL.n435 0.155672
R3069 VTAIL.n518 VTAIL.n517 0.155672
R3070 VTAIL.n517 VTAIL.n439 0.155672
R3071 VTAIL.n510 VTAIL.n439 0.155672
R3072 VTAIL.n510 VTAIL.n509 0.155672
R3073 VTAIL.n509 VTAIL.n443 0.155672
R3074 VTAIL.n502 VTAIL.n443 0.155672
R3075 VTAIL.n502 VTAIL.n501 0.155672
R3076 VTAIL.n501 VTAIL.n447 0.155672
R3077 VTAIL.n494 VTAIL.n447 0.155672
R3078 VTAIL.n494 VTAIL.n493 0.155672
R3079 VTAIL.n493 VTAIL.n451 0.155672
R3080 VTAIL.n485 VTAIL.n451 0.155672
R3081 VTAIL.n485 VTAIL.n484 0.155672
R3082 VTAIL.n484 VTAIL.n455 0.155672
R3083 VTAIL.n477 VTAIL.n455 0.155672
R3084 VTAIL.n477 VTAIL.n476 0.155672
R3085 VTAIL.n476 VTAIL.n460 0.155672
R3086 VTAIL.n469 VTAIL.n460 0.155672
R3087 VTAIL.n469 VTAIL.n468 0.155672
R3088 VTAIL.n425 VTAIL.n323 0.155672
R3089 VTAIL.n418 VTAIL.n323 0.155672
R3090 VTAIL.n418 VTAIL.n417 0.155672
R3091 VTAIL.n417 VTAIL.n327 0.155672
R3092 VTAIL.n410 VTAIL.n327 0.155672
R3093 VTAIL.n410 VTAIL.n409 0.155672
R3094 VTAIL.n409 VTAIL.n331 0.155672
R3095 VTAIL.n402 VTAIL.n331 0.155672
R3096 VTAIL.n402 VTAIL.n401 0.155672
R3097 VTAIL.n401 VTAIL.n335 0.155672
R3098 VTAIL.n394 VTAIL.n335 0.155672
R3099 VTAIL.n394 VTAIL.n393 0.155672
R3100 VTAIL.n393 VTAIL.n339 0.155672
R3101 VTAIL.n386 VTAIL.n339 0.155672
R3102 VTAIL.n386 VTAIL.n385 0.155672
R3103 VTAIL.n385 VTAIL.n343 0.155672
R3104 VTAIL.n377 VTAIL.n343 0.155672
R3105 VTAIL.n377 VTAIL.n376 0.155672
R3106 VTAIL.n376 VTAIL.n347 0.155672
R3107 VTAIL.n369 VTAIL.n347 0.155672
R3108 VTAIL.n369 VTAIL.n368 0.155672
R3109 VTAIL.n368 VTAIL.n352 0.155672
R3110 VTAIL.n361 VTAIL.n352 0.155672
R3111 VTAIL.n361 VTAIL.n360 0.155672
R3112 VTAIL VTAIL.n1 0.0586897
R3113 VDD1 VDD1.n0 71.9787
R3114 VDD1.n3 VDD1.n2 71.865
R3115 VDD1.n3 VDD1.n1 71.865
R3116 VDD1.n5 VDD1.n4 70.1704
R3117 VDD1.n5 VDD1.n3 56.8069
R3118 VDD1 VDD1.n5 1.69231
R3119 VDD1.n4 VDD1.t3 1.67257
R3120 VDD1.n4 VDD1.t7 1.67257
R3121 VDD1.n0 VDD1.t5 1.67257
R3122 VDD1.n0 VDD1.t0 1.67257
R3123 VDD1.n2 VDD1.t6 1.67257
R3124 VDD1.n2 VDD1.t2 1.67257
R3125 VDD1.n1 VDD1.t1 1.67257
R3126 VDD1.n1 VDD1.t4 1.67257
R3127 VN.n76 VN.n75 161.3
R3128 VN.n74 VN.n40 161.3
R3129 VN.n73 VN.n72 161.3
R3130 VN.n71 VN.n41 161.3
R3131 VN.n70 VN.n69 161.3
R3132 VN.n68 VN.n42 161.3
R3133 VN.n67 VN.n66 161.3
R3134 VN.n65 VN.n43 161.3
R3135 VN.n64 VN.n63 161.3
R3136 VN.n62 VN.n44 161.3
R3137 VN.n61 VN.n60 161.3
R3138 VN.n59 VN.n46 161.3
R3139 VN.n58 VN.n57 161.3
R3140 VN.n56 VN.n47 161.3
R3141 VN.n55 VN.n54 161.3
R3142 VN.n53 VN.n48 161.3
R3143 VN.n52 VN.n51 161.3
R3144 VN.n37 VN.n36 161.3
R3145 VN.n35 VN.n1 161.3
R3146 VN.n34 VN.n33 161.3
R3147 VN.n32 VN.n2 161.3
R3148 VN.n31 VN.n30 161.3
R3149 VN.n29 VN.n3 161.3
R3150 VN.n28 VN.n27 161.3
R3151 VN.n26 VN.n4 161.3
R3152 VN.n25 VN.n24 161.3
R3153 VN.n22 VN.n5 161.3
R3154 VN.n21 VN.n20 161.3
R3155 VN.n19 VN.n6 161.3
R3156 VN.n18 VN.n17 161.3
R3157 VN.n16 VN.n7 161.3
R3158 VN.n15 VN.n14 161.3
R3159 VN.n13 VN.n8 161.3
R3160 VN.n12 VN.n11 161.3
R3161 VN.n49 VN.t3 157.768
R3162 VN.n9 VN.t5 157.768
R3163 VN.n10 VN.t0 125.605
R3164 VN.n23 VN.t4 125.605
R3165 VN.n0 VN.t6 125.605
R3166 VN.n50 VN.t1 125.605
R3167 VN.n45 VN.t7 125.605
R3168 VN.n39 VN.t2 125.605
R3169 VN.n38 VN.n0 85.5092
R3170 VN.n77 VN.n39 85.5092
R3171 VN.n50 VN.n49 73.2467
R3172 VN.n10 VN.n9 73.2466
R3173 VN VN.n77 62.0434
R3174 VN.n30 VN.n2 46.253
R3175 VN.n69 VN.n41 46.253
R3176 VN.n17 VN.n16 40.4106
R3177 VN.n17 VN.n6 40.4106
R3178 VN.n57 VN.n56 40.4106
R3179 VN.n57 VN.n46 40.4106
R3180 VN.n30 VN.n29 34.5682
R3181 VN.n69 VN.n68 34.5682
R3182 VN.n11 VN.n8 24.3439
R3183 VN.n15 VN.n8 24.3439
R3184 VN.n16 VN.n15 24.3439
R3185 VN.n21 VN.n6 24.3439
R3186 VN.n22 VN.n21 24.3439
R3187 VN.n24 VN.n22 24.3439
R3188 VN.n28 VN.n4 24.3439
R3189 VN.n29 VN.n28 24.3439
R3190 VN.n34 VN.n2 24.3439
R3191 VN.n35 VN.n34 24.3439
R3192 VN.n36 VN.n35 24.3439
R3193 VN.n56 VN.n55 24.3439
R3194 VN.n55 VN.n48 24.3439
R3195 VN.n51 VN.n48 24.3439
R3196 VN.n68 VN.n67 24.3439
R3197 VN.n67 VN.n43 24.3439
R3198 VN.n63 VN.n62 24.3439
R3199 VN.n62 VN.n61 24.3439
R3200 VN.n61 VN.n46 24.3439
R3201 VN.n75 VN.n74 24.3439
R3202 VN.n74 VN.n73 24.3439
R3203 VN.n73 VN.n41 24.3439
R3204 VN.n23 VN.n4 22.8833
R3205 VN.n45 VN.n43 22.8833
R3206 VN.n36 VN.n0 4.38232
R3207 VN.n75 VN.n39 4.38232
R3208 VN.n52 VN.n49 3.3424
R3209 VN.n12 VN.n9 3.3424
R3210 VN.n11 VN.n10 1.46111
R3211 VN.n24 VN.n23 1.46111
R3212 VN.n51 VN.n50 1.46111
R3213 VN.n63 VN.n45 1.46111
R3214 VN.n77 VN.n76 0.355081
R3215 VN.n38 VN.n37 0.355081
R3216 VN VN.n38 0.26685
R3217 VN.n76 VN.n40 0.189894
R3218 VN.n72 VN.n40 0.189894
R3219 VN.n72 VN.n71 0.189894
R3220 VN.n71 VN.n70 0.189894
R3221 VN.n70 VN.n42 0.189894
R3222 VN.n66 VN.n42 0.189894
R3223 VN.n66 VN.n65 0.189894
R3224 VN.n65 VN.n64 0.189894
R3225 VN.n64 VN.n44 0.189894
R3226 VN.n60 VN.n44 0.189894
R3227 VN.n60 VN.n59 0.189894
R3228 VN.n59 VN.n58 0.189894
R3229 VN.n58 VN.n47 0.189894
R3230 VN.n54 VN.n47 0.189894
R3231 VN.n54 VN.n53 0.189894
R3232 VN.n53 VN.n52 0.189894
R3233 VN.n13 VN.n12 0.189894
R3234 VN.n14 VN.n13 0.189894
R3235 VN.n14 VN.n7 0.189894
R3236 VN.n18 VN.n7 0.189894
R3237 VN.n19 VN.n18 0.189894
R3238 VN.n20 VN.n19 0.189894
R3239 VN.n20 VN.n5 0.189894
R3240 VN.n25 VN.n5 0.189894
R3241 VN.n26 VN.n25 0.189894
R3242 VN.n27 VN.n26 0.189894
R3243 VN.n27 VN.n3 0.189894
R3244 VN.n31 VN.n3 0.189894
R3245 VN.n32 VN.n31 0.189894
R3246 VN.n33 VN.n32 0.189894
R3247 VN.n33 VN.n1 0.189894
R3248 VN.n37 VN.n1 0.189894
R3249 VDD2.n2 VDD2.n1 71.865
R3250 VDD2.n2 VDD2.n0 71.865
R3251 VDD2 VDD2.n5 71.8622
R3252 VDD2.n4 VDD2.n3 70.1705
R3253 VDD2.n4 VDD2.n2 56.2239
R3254 VDD2 VDD2.n4 1.80869
R3255 VDD2.n5 VDD2.t6 1.67257
R3256 VDD2.n5 VDD2.t4 1.67257
R3257 VDD2.n3 VDD2.t5 1.67257
R3258 VDD2.n3 VDD2.t0 1.67257
R3259 VDD2.n1 VDD2.t3 1.67257
R3260 VDD2.n1 VDD2.t1 1.67257
R3261 VDD2.n0 VDD2.t2 1.67257
R3262 VDD2.n0 VDD2.t7 1.67257
C0 B VN 1.57085f
C1 VN VDD1 0.153193f
C2 B VDD1 2.19499f
C3 w_n5030_n4856# VDD2 2.67544f
C4 w_n5030_n4856# VP 11.3665f
C5 w_n5030_n4856# VTAIL 5.91953f
C6 w_n5030_n4856# VN 10.7102f
C7 w_n5030_n4856# B 13.930901f
C8 w_n5030_n4856# VDD1 2.51333f
C9 VDD2 VP 0.639337f
C10 VDD2 VTAIL 10.704901f
C11 VDD2 VN 14.6708f
C12 B VDD2 2.32657f
C13 VDD2 VDD1 2.36204f
C14 VP VTAIL 15.1039f
C15 VP VN 10.431201f
C16 B VP 2.6771f
C17 VN VTAIL 15.089801f
C18 VP VDD1 15.155f
C19 B VTAIL 8.01912f
C20 VTAIL VDD1 10.6429f
C21 VDD2 VSUBS 2.5792f
C22 VDD1 VSUBS 3.41835f
C23 VTAIL VSUBS 1.868108f
C24 VN VSUBS 8.4998f
C25 VP VSUBS 5.010191f
C26 B VSUBS 6.891747f
C27 w_n5030_n4856# VSUBS 0.298359p
C28 VDD2.t2 VSUBS 0.477568f
C29 VDD2.t7 VSUBS 0.477568f
C30 VDD2.n0 VSUBS 4.05248f
C31 VDD2.t3 VSUBS 0.477568f
C32 VDD2.t1 VSUBS 0.477568f
C33 VDD2.n1 VSUBS 4.05248f
C34 VDD2.n2 VSUBS 6.15023f
C35 VDD2.t5 VSUBS 0.477568f
C36 VDD2.t0 VSUBS 0.477568f
C37 VDD2.n3 VSUBS 4.02583f
C38 VDD2.n4 VSUBS 5.192009f
C39 VDD2.t6 VSUBS 0.477568f
C40 VDD2.t4 VSUBS 0.477568f
C41 VDD2.n5 VSUBS 4.05242f
C42 VN.t6 VSUBS 4.12816f
C43 VN.n0 VSUBS 1.49761f
C44 VN.n1 VSUBS 0.020669f
C45 VN.n2 VSUBS 0.039621f
C46 VN.n3 VSUBS 0.020669f
C47 VN.n4 VSUBS 0.037568f
C48 VN.n5 VSUBS 0.020669f
C49 VN.n6 VSUBS 0.041299f
C50 VN.n7 VSUBS 0.020669f
C51 VN.n8 VSUBS 0.038715f
C52 VN.t5 VSUBS 4.44998f
C53 VN.n9 VSUBS 1.42533f
C54 VN.t0 VSUBS 4.12816f
C55 VN.n10 VSUBS 1.48561f
C56 VN.n11 VSUBS 0.020747f
C57 VN.n12 VSUBS 0.26329f
C58 VN.n13 VSUBS 0.020669f
C59 VN.n14 VSUBS 0.020669f
C60 VN.n15 VSUBS 0.038715f
C61 VN.n16 VSUBS 0.041299f
C62 VN.n17 VSUBS 0.016726f
C63 VN.n18 VSUBS 0.020669f
C64 VN.n19 VSUBS 0.020669f
C65 VN.n20 VSUBS 0.020669f
C66 VN.n21 VSUBS 0.038715f
C67 VN.n22 VSUBS 0.038715f
C68 VN.t4 VSUBS 4.12816f
C69 VN.n23 VSUBS 1.41917f
C70 VN.n24 VSUBS 0.020747f
C71 VN.n25 VSUBS 0.020669f
C72 VN.n26 VSUBS 0.020669f
C73 VN.n27 VSUBS 0.020669f
C74 VN.n28 VSUBS 0.038715f
C75 VN.n29 VSUBS 0.041994f
C76 VN.n30 VSUBS 0.017709f
C77 VN.n31 VSUBS 0.020669f
C78 VN.n32 VSUBS 0.020669f
C79 VN.n33 VSUBS 0.020669f
C80 VN.n34 VSUBS 0.038715f
C81 VN.n35 VSUBS 0.038715f
C82 VN.n36 VSUBS 0.023041f
C83 VN.n37 VSUBS 0.033365f
C84 VN.n38 VSUBS 0.061839f
C85 VN.t2 VSUBS 4.12816f
C86 VN.n39 VSUBS 1.49761f
C87 VN.n40 VSUBS 0.020669f
C88 VN.n41 VSUBS 0.039621f
C89 VN.n42 VSUBS 0.020669f
C90 VN.n43 VSUBS 0.037568f
C91 VN.n44 VSUBS 0.020669f
C92 VN.t7 VSUBS 4.12816f
C93 VN.n45 VSUBS 1.41917f
C94 VN.n46 VSUBS 0.041299f
C95 VN.n47 VSUBS 0.020669f
C96 VN.n48 VSUBS 0.038715f
C97 VN.t3 VSUBS 4.44998f
C98 VN.n49 VSUBS 1.42533f
C99 VN.t1 VSUBS 4.12816f
C100 VN.n50 VSUBS 1.48561f
C101 VN.n51 VSUBS 0.020747f
C102 VN.n52 VSUBS 0.26329f
C103 VN.n53 VSUBS 0.020669f
C104 VN.n54 VSUBS 0.020669f
C105 VN.n55 VSUBS 0.038715f
C106 VN.n56 VSUBS 0.041299f
C107 VN.n57 VSUBS 0.016726f
C108 VN.n58 VSUBS 0.020669f
C109 VN.n59 VSUBS 0.020669f
C110 VN.n60 VSUBS 0.020669f
C111 VN.n61 VSUBS 0.038715f
C112 VN.n62 VSUBS 0.038715f
C113 VN.n63 VSUBS 0.020747f
C114 VN.n64 VSUBS 0.020669f
C115 VN.n65 VSUBS 0.020669f
C116 VN.n66 VSUBS 0.020669f
C117 VN.n67 VSUBS 0.038715f
C118 VN.n68 VSUBS 0.041994f
C119 VN.n69 VSUBS 0.017709f
C120 VN.n70 VSUBS 0.020669f
C121 VN.n71 VSUBS 0.020669f
C122 VN.n72 VSUBS 0.020669f
C123 VN.n73 VSUBS 0.038715f
C124 VN.n74 VSUBS 0.038715f
C125 VN.n75 VSUBS 0.023041f
C126 VN.n76 VSUBS 0.033365f
C127 VN.n77 VSUBS 1.59676f
C128 VDD1.t5 VSUBS 0.477353f
C129 VDD1.t0 VSUBS 0.477353f
C130 VDD1.n0 VSUBS 4.05269f
C131 VDD1.t1 VSUBS 0.477353f
C132 VDD1.t4 VSUBS 0.477353f
C133 VDD1.n1 VSUBS 4.05066f
C134 VDD1.t6 VSUBS 0.477353f
C135 VDD1.t2 VSUBS 0.477353f
C136 VDD1.n2 VSUBS 4.05066f
C137 VDD1.n3 VSUBS 6.21113f
C138 VDD1.t3 VSUBS 0.477353f
C139 VDD1.t7 VSUBS 0.477353f
C140 VDD1.n4 VSUBS 4.024f
C141 VDD1.n5 VSUBS 5.22914f
C142 VTAIL.t2 VSUBS 0.368242f
C143 VTAIL.t15 VSUBS 0.368242f
C144 VTAIL.n0 VSUBS 2.96201f
C145 VTAIL.n1 VSUBS 0.845116f
C146 VTAIL.n2 VSUBS 0.025427f
C147 VTAIL.n3 VSUBS 0.023971f
C148 VTAIL.n4 VSUBS 0.012881f
C149 VTAIL.n5 VSUBS 0.030446f
C150 VTAIL.n6 VSUBS 0.013639f
C151 VTAIL.n7 VSUBS 0.023971f
C152 VTAIL.n8 VSUBS 0.012881f
C153 VTAIL.n9 VSUBS 0.030446f
C154 VTAIL.n10 VSUBS 0.013639f
C155 VTAIL.n11 VSUBS 0.023971f
C156 VTAIL.n12 VSUBS 0.012881f
C157 VTAIL.n13 VSUBS 0.030446f
C158 VTAIL.n14 VSUBS 0.013639f
C159 VTAIL.n15 VSUBS 0.023971f
C160 VTAIL.n16 VSUBS 0.012881f
C161 VTAIL.n17 VSUBS 0.030446f
C162 VTAIL.n18 VSUBS 0.013639f
C163 VTAIL.n19 VSUBS 0.023971f
C164 VTAIL.n20 VSUBS 0.012881f
C165 VTAIL.n21 VSUBS 0.030446f
C166 VTAIL.n22 VSUBS 0.013639f
C167 VTAIL.n23 VSUBS 0.023971f
C168 VTAIL.n24 VSUBS 0.012881f
C169 VTAIL.n25 VSUBS 0.030446f
C170 VTAIL.n26 VSUBS 0.013639f
C171 VTAIL.n27 VSUBS 0.023971f
C172 VTAIL.n28 VSUBS 0.012881f
C173 VTAIL.n29 VSUBS 0.030446f
C174 VTAIL.n30 VSUBS 0.013639f
C175 VTAIL.n31 VSUBS 0.023971f
C176 VTAIL.n32 VSUBS 0.012881f
C177 VTAIL.n33 VSUBS 0.030446f
C178 VTAIL.n34 VSUBS 0.013639f
C179 VTAIL.n35 VSUBS 0.269424f
C180 VTAIL.t1 VSUBS 0.06621f
C181 VTAIL.n36 VSUBS 0.022834f
C182 VTAIL.n37 VSUBS 0.022903f
C183 VTAIL.n38 VSUBS 0.012881f
C184 VTAIL.n39 VSUBS 1.9592f
C185 VTAIL.n40 VSUBS 0.023971f
C186 VTAIL.n41 VSUBS 0.012881f
C187 VTAIL.n42 VSUBS 0.013639f
C188 VTAIL.n43 VSUBS 0.030446f
C189 VTAIL.n44 VSUBS 0.030446f
C190 VTAIL.n45 VSUBS 0.013639f
C191 VTAIL.n46 VSUBS 0.012881f
C192 VTAIL.n47 VSUBS 0.023971f
C193 VTAIL.n48 VSUBS 0.023971f
C194 VTAIL.n49 VSUBS 0.012881f
C195 VTAIL.n50 VSUBS 0.013639f
C196 VTAIL.n51 VSUBS 0.030446f
C197 VTAIL.n52 VSUBS 0.030446f
C198 VTAIL.n53 VSUBS 0.030446f
C199 VTAIL.n54 VSUBS 0.013639f
C200 VTAIL.n55 VSUBS 0.012881f
C201 VTAIL.n56 VSUBS 0.023971f
C202 VTAIL.n57 VSUBS 0.023971f
C203 VTAIL.n58 VSUBS 0.012881f
C204 VTAIL.n59 VSUBS 0.01326f
C205 VTAIL.n60 VSUBS 0.01326f
C206 VTAIL.n61 VSUBS 0.030446f
C207 VTAIL.n62 VSUBS 0.030446f
C208 VTAIL.n63 VSUBS 0.013639f
C209 VTAIL.n64 VSUBS 0.012881f
C210 VTAIL.n65 VSUBS 0.023971f
C211 VTAIL.n66 VSUBS 0.023971f
C212 VTAIL.n67 VSUBS 0.012881f
C213 VTAIL.n68 VSUBS 0.013639f
C214 VTAIL.n69 VSUBS 0.030446f
C215 VTAIL.n70 VSUBS 0.030446f
C216 VTAIL.n71 VSUBS 0.013639f
C217 VTAIL.n72 VSUBS 0.012881f
C218 VTAIL.n73 VSUBS 0.023971f
C219 VTAIL.n74 VSUBS 0.023971f
C220 VTAIL.n75 VSUBS 0.012881f
C221 VTAIL.n76 VSUBS 0.013639f
C222 VTAIL.n77 VSUBS 0.030446f
C223 VTAIL.n78 VSUBS 0.030446f
C224 VTAIL.n79 VSUBS 0.013639f
C225 VTAIL.n80 VSUBS 0.012881f
C226 VTAIL.n81 VSUBS 0.023971f
C227 VTAIL.n82 VSUBS 0.023971f
C228 VTAIL.n83 VSUBS 0.012881f
C229 VTAIL.n84 VSUBS 0.013639f
C230 VTAIL.n85 VSUBS 0.030446f
C231 VTAIL.n86 VSUBS 0.030446f
C232 VTAIL.n87 VSUBS 0.013639f
C233 VTAIL.n88 VSUBS 0.012881f
C234 VTAIL.n89 VSUBS 0.023971f
C235 VTAIL.n90 VSUBS 0.023971f
C236 VTAIL.n91 VSUBS 0.012881f
C237 VTAIL.n92 VSUBS 0.013639f
C238 VTAIL.n93 VSUBS 0.030446f
C239 VTAIL.n94 VSUBS 0.030446f
C240 VTAIL.n95 VSUBS 0.013639f
C241 VTAIL.n96 VSUBS 0.012881f
C242 VTAIL.n97 VSUBS 0.023971f
C243 VTAIL.n98 VSUBS 0.023971f
C244 VTAIL.n99 VSUBS 0.012881f
C245 VTAIL.n100 VSUBS 0.013639f
C246 VTAIL.n101 VSUBS 0.030446f
C247 VTAIL.n102 VSUBS 0.074904f
C248 VTAIL.n103 VSUBS 0.013639f
C249 VTAIL.n104 VSUBS 0.025295f
C250 VTAIL.n105 VSUBS 0.059337f
C251 VTAIL.n106 VSUBS 0.056987f
C252 VTAIL.n107 VSUBS 0.329322f
C253 VTAIL.n108 VSUBS 0.025427f
C254 VTAIL.n109 VSUBS 0.023971f
C255 VTAIL.n110 VSUBS 0.012881f
C256 VTAIL.n111 VSUBS 0.030446f
C257 VTAIL.n112 VSUBS 0.013639f
C258 VTAIL.n113 VSUBS 0.023971f
C259 VTAIL.n114 VSUBS 0.012881f
C260 VTAIL.n115 VSUBS 0.030446f
C261 VTAIL.n116 VSUBS 0.013639f
C262 VTAIL.n117 VSUBS 0.023971f
C263 VTAIL.n118 VSUBS 0.012881f
C264 VTAIL.n119 VSUBS 0.030446f
C265 VTAIL.n120 VSUBS 0.013639f
C266 VTAIL.n121 VSUBS 0.023971f
C267 VTAIL.n122 VSUBS 0.012881f
C268 VTAIL.n123 VSUBS 0.030446f
C269 VTAIL.n124 VSUBS 0.013639f
C270 VTAIL.n125 VSUBS 0.023971f
C271 VTAIL.n126 VSUBS 0.012881f
C272 VTAIL.n127 VSUBS 0.030446f
C273 VTAIL.n128 VSUBS 0.013639f
C274 VTAIL.n129 VSUBS 0.023971f
C275 VTAIL.n130 VSUBS 0.012881f
C276 VTAIL.n131 VSUBS 0.030446f
C277 VTAIL.n132 VSUBS 0.013639f
C278 VTAIL.n133 VSUBS 0.023971f
C279 VTAIL.n134 VSUBS 0.012881f
C280 VTAIL.n135 VSUBS 0.030446f
C281 VTAIL.n136 VSUBS 0.013639f
C282 VTAIL.n137 VSUBS 0.023971f
C283 VTAIL.n138 VSUBS 0.012881f
C284 VTAIL.n139 VSUBS 0.030446f
C285 VTAIL.n140 VSUBS 0.013639f
C286 VTAIL.n141 VSUBS 0.269424f
C287 VTAIL.t5 VSUBS 0.06621f
C288 VTAIL.n142 VSUBS 0.022834f
C289 VTAIL.n143 VSUBS 0.022903f
C290 VTAIL.n144 VSUBS 0.012881f
C291 VTAIL.n145 VSUBS 1.9592f
C292 VTAIL.n146 VSUBS 0.023971f
C293 VTAIL.n147 VSUBS 0.012881f
C294 VTAIL.n148 VSUBS 0.013639f
C295 VTAIL.n149 VSUBS 0.030446f
C296 VTAIL.n150 VSUBS 0.030446f
C297 VTAIL.n151 VSUBS 0.013639f
C298 VTAIL.n152 VSUBS 0.012881f
C299 VTAIL.n153 VSUBS 0.023971f
C300 VTAIL.n154 VSUBS 0.023971f
C301 VTAIL.n155 VSUBS 0.012881f
C302 VTAIL.n156 VSUBS 0.013639f
C303 VTAIL.n157 VSUBS 0.030446f
C304 VTAIL.n158 VSUBS 0.030446f
C305 VTAIL.n159 VSUBS 0.030446f
C306 VTAIL.n160 VSUBS 0.013639f
C307 VTAIL.n161 VSUBS 0.012881f
C308 VTAIL.n162 VSUBS 0.023971f
C309 VTAIL.n163 VSUBS 0.023971f
C310 VTAIL.n164 VSUBS 0.012881f
C311 VTAIL.n165 VSUBS 0.01326f
C312 VTAIL.n166 VSUBS 0.01326f
C313 VTAIL.n167 VSUBS 0.030446f
C314 VTAIL.n168 VSUBS 0.030446f
C315 VTAIL.n169 VSUBS 0.013639f
C316 VTAIL.n170 VSUBS 0.012881f
C317 VTAIL.n171 VSUBS 0.023971f
C318 VTAIL.n172 VSUBS 0.023971f
C319 VTAIL.n173 VSUBS 0.012881f
C320 VTAIL.n174 VSUBS 0.013639f
C321 VTAIL.n175 VSUBS 0.030446f
C322 VTAIL.n176 VSUBS 0.030446f
C323 VTAIL.n177 VSUBS 0.013639f
C324 VTAIL.n178 VSUBS 0.012881f
C325 VTAIL.n179 VSUBS 0.023971f
C326 VTAIL.n180 VSUBS 0.023971f
C327 VTAIL.n181 VSUBS 0.012881f
C328 VTAIL.n182 VSUBS 0.013639f
C329 VTAIL.n183 VSUBS 0.030446f
C330 VTAIL.n184 VSUBS 0.030446f
C331 VTAIL.n185 VSUBS 0.013639f
C332 VTAIL.n186 VSUBS 0.012881f
C333 VTAIL.n187 VSUBS 0.023971f
C334 VTAIL.n188 VSUBS 0.023971f
C335 VTAIL.n189 VSUBS 0.012881f
C336 VTAIL.n190 VSUBS 0.013639f
C337 VTAIL.n191 VSUBS 0.030446f
C338 VTAIL.n192 VSUBS 0.030446f
C339 VTAIL.n193 VSUBS 0.013639f
C340 VTAIL.n194 VSUBS 0.012881f
C341 VTAIL.n195 VSUBS 0.023971f
C342 VTAIL.n196 VSUBS 0.023971f
C343 VTAIL.n197 VSUBS 0.012881f
C344 VTAIL.n198 VSUBS 0.013639f
C345 VTAIL.n199 VSUBS 0.030446f
C346 VTAIL.n200 VSUBS 0.030446f
C347 VTAIL.n201 VSUBS 0.013639f
C348 VTAIL.n202 VSUBS 0.012881f
C349 VTAIL.n203 VSUBS 0.023971f
C350 VTAIL.n204 VSUBS 0.023971f
C351 VTAIL.n205 VSUBS 0.012881f
C352 VTAIL.n206 VSUBS 0.013639f
C353 VTAIL.n207 VSUBS 0.030446f
C354 VTAIL.n208 VSUBS 0.074904f
C355 VTAIL.n209 VSUBS 0.013639f
C356 VTAIL.n210 VSUBS 0.025295f
C357 VTAIL.n211 VSUBS 0.059337f
C358 VTAIL.n212 VSUBS 0.056987f
C359 VTAIL.n213 VSUBS 0.329322f
C360 VTAIL.t10 VSUBS 0.368242f
C361 VTAIL.t4 VSUBS 0.368242f
C362 VTAIL.n214 VSUBS 2.96201f
C363 VTAIL.n215 VSUBS 1.11096f
C364 VTAIL.n216 VSUBS 0.025427f
C365 VTAIL.n217 VSUBS 0.023971f
C366 VTAIL.n218 VSUBS 0.012881f
C367 VTAIL.n219 VSUBS 0.030446f
C368 VTAIL.n220 VSUBS 0.013639f
C369 VTAIL.n221 VSUBS 0.023971f
C370 VTAIL.n222 VSUBS 0.012881f
C371 VTAIL.n223 VSUBS 0.030446f
C372 VTAIL.n224 VSUBS 0.013639f
C373 VTAIL.n225 VSUBS 0.023971f
C374 VTAIL.n226 VSUBS 0.012881f
C375 VTAIL.n227 VSUBS 0.030446f
C376 VTAIL.n228 VSUBS 0.013639f
C377 VTAIL.n229 VSUBS 0.023971f
C378 VTAIL.n230 VSUBS 0.012881f
C379 VTAIL.n231 VSUBS 0.030446f
C380 VTAIL.n232 VSUBS 0.013639f
C381 VTAIL.n233 VSUBS 0.023971f
C382 VTAIL.n234 VSUBS 0.012881f
C383 VTAIL.n235 VSUBS 0.030446f
C384 VTAIL.n236 VSUBS 0.013639f
C385 VTAIL.n237 VSUBS 0.023971f
C386 VTAIL.n238 VSUBS 0.012881f
C387 VTAIL.n239 VSUBS 0.030446f
C388 VTAIL.n240 VSUBS 0.013639f
C389 VTAIL.n241 VSUBS 0.023971f
C390 VTAIL.n242 VSUBS 0.012881f
C391 VTAIL.n243 VSUBS 0.030446f
C392 VTAIL.n244 VSUBS 0.013639f
C393 VTAIL.n245 VSUBS 0.023971f
C394 VTAIL.n246 VSUBS 0.012881f
C395 VTAIL.n247 VSUBS 0.030446f
C396 VTAIL.n248 VSUBS 0.013639f
C397 VTAIL.n249 VSUBS 0.269424f
C398 VTAIL.t8 VSUBS 0.06621f
C399 VTAIL.n250 VSUBS 0.022834f
C400 VTAIL.n251 VSUBS 0.022903f
C401 VTAIL.n252 VSUBS 0.012881f
C402 VTAIL.n253 VSUBS 1.9592f
C403 VTAIL.n254 VSUBS 0.023971f
C404 VTAIL.n255 VSUBS 0.012881f
C405 VTAIL.n256 VSUBS 0.013639f
C406 VTAIL.n257 VSUBS 0.030446f
C407 VTAIL.n258 VSUBS 0.030446f
C408 VTAIL.n259 VSUBS 0.013639f
C409 VTAIL.n260 VSUBS 0.012881f
C410 VTAIL.n261 VSUBS 0.023971f
C411 VTAIL.n262 VSUBS 0.023971f
C412 VTAIL.n263 VSUBS 0.012881f
C413 VTAIL.n264 VSUBS 0.013639f
C414 VTAIL.n265 VSUBS 0.030446f
C415 VTAIL.n266 VSUBS 0.030446f
C416 VTAIL.n267 VSUBS 0.030446f
C417 VTAIL.n268 VSUBS 0.013639f
C418 VTAIL.n269 VSUBS 0.012881f
C419 VTAIL.n270 VSUBS 0.023971f
C420 VTAIL.n271 VSUBS 0.023971f
C421 VTAIL.n272 VSUBS 0.012881f
C422 VTAIL.n273 VSUBS 0.01326f
C423 VTAIL.n274 VSUBS 0.01326f
C424 VTAIL.n275 VSUBS 0.030446f
C425 VTAIL.n276 VSUBS 0.030446f
C426 VTAIL.n277 VSUBS 0.013639f
C427 VTAIL.n278 VSUBS 0.012881f
C428 VTAIL.n279 VSUBS 0.023971f
C429 VTAIL.n280 VSUBS 0.023971f
C430 VTAIL.n281 VSUBS 0.012881f
C431 VTAIL.n282 VSUBS 0.013639f
C432 VTAIL.n283 VSUBS 0.030446f
C433 VTAIL.n284 VSUBS 0.030446f
C434 VTAIL.n285 VSUBS 0.013639f
C435 VTAIL.n286 VSUBS 0.012881f
C436 VTAIL.n287 VSUBS 0.023971f
C437 VTAIL.n288 VSUBS 0.023971f
C438 VTAIL.n289 VSUBS 0.012881f
C439 VTAIL.n290 VSUBS 0.013639f
C440 VTAIL.n291 VSUBS 0.030446f
C441 VTAIL.n292 VSUBS 0.030446f
C442 VTAIL.n293 VSUBS 0.013639f
C443 VTAIL.n294 VSUBS 0.012881f
C444 VTAIL.n295 VSUBS 0.023971f
C445 VTAIL.n296 VSUBS 0.023971f
C446 VTAIL.n297 VSUBS 0.012881f
C447 VTAIL.n298 VSUBS 0.013639f
C448 VTAIL.n299 VSUBS 0.030446f
C449 VTAIL.n300 VSUBS 0.030446f
C450 VTAIL.n301 VSUBS 0.013639f
C451 VTAIL.n302 VSUBS 0.012881f
C452 VTAIL.n303 VSUBS 0.023971f
C453 VTAIL.n304 VSUBS 0.023971f
C454 VTAIL.n305 VSUBS 0.012881f
C455 VTAIL.n306 VSUBS 0.013639f
C456 VTAIL.n307 VSUBS 0.030446f
C457 VTAIL.n308 VSUBS 0.030446f
C458 VTAIL.n309 VSUBS 0.013639f
C459 VTAIL.n310 VSUBS 0.012881f
C460 VTAIL.n311 VSUBS 0.023971f
C461 VTAIL.n312 VSUBS 0.023971f
C462 VTAIL.n313 VSUBS 0.012881f
C463 VTAIL.n314 VSUBS 0.013639f
C464 VTAIL.n315 VSUBS 0.030446f
C465 VTAIL.n316 VSUBS 0.074904f
C466 VTAIL.n317 VSUBS 0.013639f
C467 VTAIL.n318 VSUBS 0.025295f
C468 VTAIL.n319 VSUBS 0.059337f
C469 VTAIL.n320 VSUBS 0.056987f
C470 VTAIL.n321 VSUBS 2.18342f
C471 VTAIL.n322 VSUBS 0.025427f
C472 VTAIL.n323 VSUBS 0.023971f
C473 VTAIL.n324 VSUBS 0.012881f
C474 VTAIL.n325 VSUBS 0.030446f
C475 VTAIL.n326 VSUBS 0.013639f
C476 VTAIL.n327 VSUBS 0.023971f
C477 VTAIL.n328 VSUBS 0.012881f
C478 VTAIL.n329 VSUBS 0.030446f
C479 VTAIL.n330 VSUBS 0.013639f
C480 VTAIL.n331 VSUBS 0.023971f
C481 VTAIL.n332 VSUBS 0.012881f
C482 VTAIL.n333 VSUBS 0.030446f
C483 VTAIL.n334 VSUBS 0.013639f
C484 VTAIL.n335 VSUBS 0.023971f
C485 VTAIL.n336 VSUBS 0.012881f
C486 VTAIL.n337 VSUBS 0.030446f
C487 VTAIL.n338 VSUBS 0.013639f
C488 VTAIL.n339 VSUBS 0.023971f
C489 VTAIL.n340 VSUBS 0.012881f
C490 VTAIL.n341 VSUBS 0.030446f
C491 VTAIL.n342 VSUBS 0.013639f
C492 VTAIL.n343 VSUBS 0.023971f
C493 VTAIL.n344 VSUBS 0.012881f
C494 VTAIL.n345 VSUBS 0.030446f
C495 VTAIL.n346 VSUBS 0.013639f
C496 VTAIL.n347 VSUBS 0.023971f
C497 VTAIL.n348 VSUBS 0.012881f
C498 VTAIL.n349 VSUBS 0.030446f
C499 VTAIL.n350 VSUBS 0.030446f
C500 VTAIL.n351 VSUBS 0.013639f
C501 VTAIL.n352 VSUBS 0.023971f
C502 VTAIL.n353 VSUBS 0.012881f
C503 VTAIL.n354 VSUBS 0.030446f
C504 VTAIL.n355 VSUBS 0.013639f
C505 VTAIL.n356 VSUBS 0.269424f
C506 VTAIL.t13 VSUBS 0.06621f
C507 VTAIL.n357 VSUBS 0.022834f
C508 VTAIL.n358 VSUBS 0.022903f
C509 VTAIL.n359 VSUBS 0.012881f
C510 VTAIL.n360 VSUBS 1.9592f
C511 VTAIL.n361 VSUBS 0.023971f
C512 VTAIL.n362 VSUBS 0.012881f
C513 VTAIL.n363 VSUBS 0.013639f
C514 VTAIL.n364 VSUBS 0.030446f
C515 VTAIL.n365 VSUBS 0.030446f
C516 VTAIL.n366 VSUBS 0.013639f
C517 VTAIL.n367 VSUBS 0.012881f
C518 VTAIL.n368 VSUBS 0.023971f
C519 VTAIL.n369 VSUBS 0.023971f
C520 VTAIL.n370 VSUBS 0.012881f
C521 VTAIL.n371 VSUBS 0.013639f
C522 VTAIL.n372 VSUBS 0.030446f
C523 VTAIL.n373 VSUBS 0.030446f
C524 VTAIL.n374 VSUBS 0.013639f
C525 VTAIL.n375 VSUBS 0.012881f
C526 VTAIL.n376 VSUBS 0.023971f
C527 VTAIL.n377 VSUBS 0.023971f
C528 VTAIL.n378 VSUBS 0.012881f
C529 VTAIL.n379 VSUBS 0.01326f
C530 VTAIL.n380 VSUBS 0.01326f
C531 VTAIL.n381 VSUBS 0.030446f
C532 VTAIL.n382 VSUBS 0.030446f
C533 VTAIL.n383 VSUBS 0.013639f
C534 VTAIL.n384 VSUBS 0.012881f
C535 VTAIL.n385 VSUBS 0.023971f
C536 VTAIL.n386 VSUBS 0.023971f
C537 VTAIL.n387 VSUBS 0.012881f
C538 VTAIL.n388 VSUBS 0.013639f
C539 VTAIL.n389 VSUBS 0.030446f
C540 VTAIL.n390 VSUBS 0.030446f
C541 VTAIL.n391 VSUBS 0.013639f
C542 VTAIL.n392 VSUBS 0.012881f
C543 VTAIL.n393 VSUBS 0.023971f
C544 VTAIL.n394 VSUBS 0.023971f
C545 VTAIL.n395 VSUBS 0.012881f
C546 VTAIL.n396 VSUBS 0.013639f
C547 VTAIL.n397 VSUBS 0.030446f
C548 VTAIL.n398 VSUBS 0.030446f
C549 VTAIL.n399 VSUBS 0.013639f
C550 VTAIL.n400 VSUBS 0.012881f
C551 VTAIL.n401 VSUBS 0.023971f
C552 VTAIL.n402 VSUBS 0.023971f
C553 VTAIL.n403 VSUBS 0.012881f
C554 VTAIL.n404 VSUBS 0.013639f
C555 VTAIL.n405 VSUBS 0.030446f
C556 VTAIL.n406 VSUBS 0.030446f
C557 VTAIL.n407 VSUBS 0.013639f
C558 VTAIL.n408 VSUBS 0.012881f
C559 VTAIL.n409 VSUBS 0.023971f
C560 VTAIL.n410 VSUBS 0.023971f
C561 VTAIL.n411 VSUBS 0.012881f
C562 VTAIL.n412 VSUBS 0.013639f
C563 VTAIL.n413 VSUBS 0.030446f
C564 VTAIL.n414 VSUBS 0.030446f
C565 VTAIL.n415 VSUBS 0.013639f
C566 VTAIL.n416 VSUBS 0.012881f
C567 VTAIL.n417 VSUBS 0.023971f
C568 VTAIL.n418 VSUBS 0.023971f
C569 VTAIL.n419 VSUBS 0.012881f
C570 VTAIL.n420 VSUBS 0.013639f
C571 VTAIL.n421 VSUBS 0.030446f
C572 VTAIL.n422 VSUBS 0.074904f
C573 VTAIL.n423 VSUBS 0.013639f
C574 VTAIL.n424 VSUBS 0.025295f
C575 VTAIL.n425 VSUBS 0.059337f
C576 VTAIL.n426 VSUBS 0.056987f
C577 VTAIL.n427 VSUBS 2.18342f
C578 VTAIL.t0 VSUBS 0.368242f
C579 VTAIL.t12 VSUBS 0.368242f
C580 VTAIL.n428 VSUBS 2.96203f
C581 VTAIL.n429 VSUBS 1.11094f
C582 VTAIL.n430 VSUBS 0.025427f
C583 VTAIL.n431 VSUBS 0.023971f
C584 VTAIL.n432 VSUBS 0.012881f
C585 VTAIL.n433 VSUBS 0.030446f
C586 VTAIL.n434 VSUBS 0.013639f
C587 VTAIL.n435 VSUBS 0.023971f
C588 VTAIL.n436 VSUBS 0.012881f
C589 VTAIL.n437 VSUBS 0.030446f
C590 VTAIL.n438 VSUBS 0.013639f
C591 VTAIL.n439 VSUBS 0.023971f
C592 VTAIL.n440 VSUBS 0.012881f
C593 VTAIL.n441 VSUBS 0.030446f
C594 VTAIL.n442 VSUBS 0.013639f
C595 VTAIL.n443 VSUBS 0.023971f
C596 VTAIL.n444 VSUBS 0.012881f
C597 VTAIL.n445 VSUBS 0.030446f
C598 VTAIL.n446 VSUBS 0.013639f
C599 VTAIL.n447 VSUBS 0.023971f
C600 VTAIL.n448 VSUBS 0.012881f
C601 VTAIL.n449 VSUBS 0.030446f
C602 VTAIL.n450 VSUBS 0.013639f
C603 VTAIL.n451 VSUBS 0.023971f
C604 VTAIL.n452 VSUBS 0.012881f
C605 VTAIL.n453 VSUBS 0.030446f
C606 VTAIL.n454 VSUBS 0.013639f
C607 VTAIL.n455 VSUBS 0.023971f
C608 VTAIL.n456 VSUBS 0.012881f
C609 VTAIL.n457 VSUBS 0.030446f
C610 VTAIL.n458 VSUBS 0.030446f
C611 VTAIL.n459 VSUBS 0.013639f
C612 VTAIL.n460 VSUBS 0.023971f
C613 VTAIL.n461 VSUBS 0.012881f
C614 VTAIL.n462 VSUBS 0.030446f
C615 VTAIL.n463 VSUBS 0.013639f
C616 VTAIL.n464 VSUBS 0.269424f
C617 VTAIL.t14 VSUBS 0.06621f
C618 VTAIL.n465 VSUBS 0.022834f
C619 VTAIL.n466 VSUBS 0.022903f
C620 VTAIL.n467 VSUBS 0.012881f
C621 VTAIL.n468 VSUBS 1.9592f
C622 VTAIL.n469 VSUBS 0.023971f
C623 VTAIL.n470 VSUBS 0.012881f
C624 VTAIL.n471 VSUBS 0.013639f
C625 VTAIL.n472 VSUBS 0.030446f
C626 VTAIL.n473 VSUBS 0.030446f
C627 VTAIL.n474 VSUBS 0.013639f
C628 VTAIL.n475 VSUBS 0.012881f
C629 VTAIL.n476 VSUBS 0.023971f
C630 VTAIL.n477 VSUBS 0.023971f
C631 VTAIL.n478 VSUBS 0.012881f
C632 VTAIL.n479 VSUBS 0.013639f
C633 VTAIL.n480 VSUBS 0.030446f
C634 VTAIL.n481 VSUBS 0.030446f
C635 VTAIL.n482 VSUBS 0.013639f
C636 VTAIL.n483 VSUBS 0.012881f
C637 VTAIL.n484 VSUBS 0.023971f
C638 VTAIL.n485 VSUBS 0.023971f
C639 VTAIL.n486 VSUBS 0.012881f
C640 VTAIL.n487 VSUBS 0.01326f
C641 VTAIL.n488 VSUBS 0.01326f
C642 VTAIL.n489 VSUBS 0.030446f
C643 VTAIL.n490 VSUBS 0.030446f
C644 VTAIL.n491 VSUBS 0.013639f
C645 VTAIL.n492 VSUBS 0.012881f
C646 VTAIL.n493 VSUBS 0.023971f
C647 VTAIL.n494 VSUBS 0.023971f
C648 VTAIL.n495 VSUBS 0.012881f
C649 VTAIL.n496 VSUBS 0.013639f
C650 VTAIL.n497 VSUBS 0.030446f
C651 VTAIL.n498 VSUBS 0.030446f
C652 VTAIL.n499 VSUBS 0.013639f
C653 VTAIL.n500 VSUBS 0.012881f
C654 VTAIL.n501 VSUBS 0.023971f
C655 VTAIL.n502 VSUBS 0.023971f
C656 VTAIL.n503 VSUBS 0.012881f
C657 VTAIL.n504 VSUBS 0.013639f
C658 VTAIL.n505 VSUBS 0.030446f
C659 VTAIL.n506 VSUBS 0.030446f
C660 VTAIL.n507 VSUBS 0.013639f
C661 VTAIL.n508 VSUBS 0.012881f
C662 VTAIL.n509 VSUBS 0.023971f
C663 VTAIL.n510 VSUBS 0.023971f
C664 VTAIL.n511 VSUBS 0.012881f
C665 VTAIL.n512 VSUBS 0.013639f
C666 VTAIL.n513 VSUBS 0.030446f
C667 VTAIL.n514 VSUBS 0.030446f
C668 VTAIL.n515 VSUBS 0.013639f
C669 VTAIL.n516 VSUBS 0.012881f
C670 VTAIL.n517 VSUBS 0.023971f
C671 VTAIL.n518 VSUBS 0.023971f
C672 VTAIL.n519 VSUBS 0.012881f
C673 VTAIL.n520 VSUBS 0.013639f
C674 VTAIL.n521 VSUBS 0.030446f
C675 VTAIL.n522 VSUBS 0.030446f
C676 VTAIL.n523 VSUBS 0.013639f
C677 VTAIL.n524 VSUBS 0.012881f
C678 VTAIL.n525 VSUBS 0.023971f
C679 VTAIL.n526 VSUBS 0.023971f
C680 VTAIL.n527 VSUBS 0.012881f
C681 VTAIL.n528 VSUBS 0.013639f
C682 VTAIL.n529 VSUBS 0.030446f
C683 VTAIL.n530 VSUBS 0.074904f
C684 VTAIL.n531 VSUBS 0.013639f
C685 VTAIL.n532 VSUBS 0.025295f
C686 VTAIL.n533 VSUBS 0.059337f
C687 VTAIL.n534 VSUBS 0.056987f
C688 VTAIL.n535 VSUBS 0.329322f
C689 VTAIL.n536 VSUBS 0.025427f
C690 VTAIL.n537 VSUBS 0.023971f
C691 VTAIL.n538 VSUBS 0.012881f
C692 VTAIL.n539 VSUBS 0.030446f
C693 VTAIL.n540 VSUBS 0.013639f
C694 VTAIL.n541 VSUBS 0.023971f
C695 VTAIL.n542 VSUBS 0.012881f
C696 VTAIL.n543 VSUBS 0.030446f
C697 VTAIL.n544 VSUBS 0.013639f
C698 VTAIL.n545 VSUBS 0.023971f
C699 VTAIL.n546 VSUBS 0.012881f
C700 VTAIL.n547 VSUBS 0.030446f
C701 VTAIL.n548 VSUBS 0.013639f
C702 VTAIL.n549 VSUBS 0.023971f
C703 VTAIL.n550 VSUBS 0.012881f
C704 VTAIL.n551 VSUBS 0.030446f
C705 VTAIL.n552 VSUBS 0.013639f
C706 VTAIL.n553 VSUBS 0.023971f
C707 VTAIL.n554 VSUBS 0.012881f
C708 VTAIL.n555 VSUBS 0.030446f
C709 VTAIL.n556 VSUBS 0.013639f
C710 VTAIL.n557 VSUBS 0.023971f
C711 VTAIL.n558 VSUBS 0.012881f
C712 VTAIL.n559 VSUBS 0.030446f
C713 VTAIL.n560 VSUBS 0.013639f
C714 VTAIL.n561 VSUBS 0.023971f
C715 VTAIL.n562 VSUBS 0.012881f
C716 VTAIL.n563 VSUBS 0.030446f
C717 VTAIL.n564 VSUBS 0.030446f
C718 VTAIL.n565 VSUBS 0.013639f
C719 VTAIL.n566 VSUBS 0.023971f
C720 VTAIL.n567 VSUBS 0.012881f
C721 VTAIL.n568 VSUBS 0.030446f
C722 VTAIL.n569 VSUBS 0.013639f
C723 VTAIL.n570 VSUBS 0.269424f
C724 VTAIL.t3 VSUBS 0.06621f
C725 VTAIL.n571 VSUBS 0.022834f
C726 VTAIL.n572 VSUBS 0.022903f
C727 VTAIL.n573 VSUBS 0.012881f
C728 VTAIL.n574 VSUBS 1.9592f
C729 VTAIL.n575 VSUBS 0.023971f
C730 VTAIL.n576 VSUBS 0.012881f
C731 VTAIL.n577 VSUBS 0.013639f
C732 VTAIL.n578 VSUBS 0.030446f
C733 VTAIL.n579 VSUBS 0.030446f
C734 VTAIL.n580 VSUBS 0.013639f
C735 VTAIL.n581 VSUBS 0.012881f
C736 VTAIL.n582 VSUBS 0.023971f
C737 VTAIL.n583 VSUBS 0.023971f
C738 VTAIL.n584 VSUBS 0.012881f
C739 VTAIL.n585 VSUBS 0.013639f
C740 VTAIL.n586 VSUBS 0.030446f
C741 VTAIL.n587 VSUBS 0.030446f
C742 VTAIL.n588 VSUBS 0.013639f
C743 VTAIL.n589 VSUBS 0.012881f
C744 VTAIL.n590 VSUBS 0.023971f
C745 VTAIL.n591 VSUBS 0.023971f
C746 VTAIL.n592 VSUBS 0.012881f
C747 VTAIL.n593 VSUBS 0.01326f
C748 VTAIL.n594 VSUBS 0.01326f
C749 VTAIL.n595 VSUBS 0.030446f
C750 VTAIL.n596 VSUBS 0.030446f
C751 VTAIL.n597 VSUBS 0.013639f
C752 VTAIL.n598 VSUBS 0.012881f
C753 VTAIL.n599 VSUBS 0.023971f
C754 VTAIL.n600 VSUBS 0.023971f
C755 VTAIL.n601 VSUBS 0.012881f
C756 VTAIL.n602 VSUBS 0.013639f
C757 VTAIL.n603 VSUBS 0.030446f
C758 VTAIL.n604 VSUBS 0.030446f
C759 VTAIL.n605 VSUBS 0.013639f
C760 VTAIL.n606 VSUBS 0.012881f
C761 VTAIL.n607 VSUBS 0.023971f
C762 VTAIL.n608 VSUBS 0.023971f
C763 VTAIL.n609 VSUBS 0.012881f
C764 VTAIL.n610 VSUBS 0.013639f
C765 VTAIL.n611 VSUBS 0.030446f
C766 VTAIL.n612 VSUBS 0.030446f
C767 VTAIL.n613 VSUBS 0.013639f
C768 VTAIL.n614 VSUBS 0.012881f
C769 VTAIL.n615 VSUBS 0.023971f
C770 VTAIL.n616 VSUBS 0.023971f
C771 VTAIL.n617 VSUBS 0.012881f
C772 VTAIL.n618 VSUBS 0.013639f
C773 VTAIL.n619 VSUBS 0.030446f
C774 VTAIL.n620 VSUBS 0.030446f
C775 VTAIL.n621 VSUBS 0.013639f
C776 VTAIL.n622 VSUBS 0.012881f
C777 VTAIL.n623 VSUBS 0.023971f
C778 VTAIL.n624 VSUBS 0.023971f
C779 VTAIL.n625 VSUBS 0.012881f
C780 VTAIL.n626 VSUBS 0.013639f
C781 VTAIL.n627 VSUBS 0.030446f
C782 VTAIL.n628 VSUBS 0.030446f
C783 VTAIL.n629 VSUBS 0.013639f
C784 VTAIL.n630 VSUBS 0.012881f
C785 VTAIL.n631 VSUBS 0.023971f
C786 VTAIL.n632 VSUBS 0.023971f
C787 VTAIL.n633 VSUBS 0.012881f
C788 VTAIL.n634 VSUBS 0.013639f
C789 VTAIL.n635 VSUBS 0.030446f
C790 VTAIL.n636 VSUBS 0.074904f
C791 VTAIL.n637 VSUBS 0.013639f
C792 VTAIL.n638 VSUBS 0.025295f
C793 VTAIL.n639 VSUBS 0.059337f
C794 VTAIL.n640 VSUBS 0.056987f
C795 VTAIL.n641 VSUBS 0.329322f
C796 VTAIL.t6 VSUBS 0.368242f
C797 VTAIL.t7 VSUBS 0.368242f
C798 VTAIL.n642 VSUBS 2.96203f
C799 VTAIL.n643 VSUBS 1.11094f
C800 VTAIL.n644 VSUBS 0.025427f
C801 VTAIL.n645 VSUBS 0.023971f
C802 VTAIL.n646 VSUBS 0.012881f
C803 VTAIL.n647 VSUBS 0.030446f
C804 VTAIL.n648 VSUBS 0.013639f
C805 VTAIL.n649 VSUBS 0.023971f
C806 VTAIL.n650 VSUBS 0.012881f
C807 VTAIL.n651 VSUBS 0.030446f
C808 VTAIL.n652 VSUBS 0.013639f
C809 VTAIL.n653 VSUBS 0.023971f
C810 VTAIL.n654 VSUBS 0.012881f
C811 VTAIL.n655 VSUBS 0.030446f
C812 VTAIL.n656 VSUBS 0.013639f
C813 VTAIL.n657 VSUBS 0.023971f
C814 VTAIL.n658 VSUBS 0.012881f
C815 VTAIL.n659 VSUBS 0.030446f
C816 VTAIL.n660 VSUBS 0.013639f
C817 VTAIL.n661 VSUBS 0.023971f
C818 VTAIL.n662 VSUBS 0.012881f
C819 VTAIL.n663 VSUBS 0.030446f
C820 VTAIL.n664 VSUBS 0.013639f
C821 VTAIL.n665 VSUBS 0.023971f
C822 VTAIL.n666 VSUBS 0.012881f
C823 VTAIL.n667 VSUBS 0.030446f
C824 VTAIL.n668 VSUBS 0.013639f
C825 VTAIL.n669 VSUBS 0.023971f
C826 VTAIL.n670 VSUBS 0.012881f
C827 VTAIL.n671 VSUBS 0.030446f
C828 VTAIL.n672 VSUBS 0.030446f
C829 VTAIL.n673 VSUBS 0.013639f
C830 VTAIL.n674 VSUBS 0.023971f
C831 VTAIL.n675 VSUBS 0.012881f
C832 VTAIL.n676 VSUBS 0.030446f
C833 VTAIL.n677 VSUBS 0.013639f
C834 VTAIL.n678 VSUBS 0.269424f
C835 VTAIL.t9 VSUBS 0.06621f
C836 VTAIL.n679 VSUBS 0.022834f
C837 VTAIL.n680 VSUBS 0.022903f
C838 VTAIL.n681 VSUBS 0.012881f
C839 VTAIL.n682 VSUBS 1.9592f
C840 VTAIL.n683 VSUBS 0.023971f
C841 VTAIL.n684 VSUBS 0.012881f
C842 VTAIL.n685 VSUBS 0.013639f
C843 VTAIL.n686 VSUBS 0.030446f
C844 VTAIL.n687 VSUBS 0.030446f
C845 VTAIL.n688 VSUBS 0.013639f
C846 VTAIL.n689 VSUBS 0.012881f
C847 VTAIL.n690 VSUBS 0.023971f
C848 VTAIL.n691 VSUBS 0.023971f
C849 VTAIL.n692 VSUBS 0.012881f
C850 VTAIL.n693 VSUBS 0.013639f
C851 VTAIL.n694 VSUBS 0.030446f
C852 VTAIL.n695 VSUBS 0.030446f
C853 VTAIL.n696 VSUBS 0.013639f
C854 VTAIL.n697 VSUBS 0.012881f
C855 VTAIL.n698 VSUBS 0.023971f
C856 VTAIL.n699 VSUBS 0.023971f
C857 VTAIL.n700 VSUBS 0.012881f
C858 VTAIL.n701 VSUBS 0.01326f
C859 VTAIL.n702 VSUBS 0.01326f
C860 VTAIL.n703 VSUBS 0.030446f
C861 VTAIL.n704 VSUBS 0.030446f
C862 VTAIL.n705 VSUBS 0.013639f
C863 VTAIL.n706 VSUBS 0.012881f
C864 VTAIL.n707 VSUBS 0.023971f
C865 VTAIL.n708 VSUBS 0.023971f
C866 VTAIL.n709 VSUBS 0.012881f
C867 VTAIL.n710 VSUBS 0.013639f
C868 VTAIL.n711 VSUBS 0.030446f
C869 VTAIL.n712 VSUBS 0.030446f
C870 VTAIL.n713 VSUBS 0.013639f
C871 VTAIL.n714 VSUBS 0.012881f
C872 VTAIL.n715 VSUBS 0.023971f
C873 VTAIL.n716 VSUBS 0.023971f
C874 VTAIL.n717 VSUBS 0.012881f
C875 VTAIL.n718 VSUBS 0.013639f
C876 VTAIL.n719 VSUBS 0.030446f
C877 VTAIL.n720 VSUBS 0.030446f
C878 VTAIL.n721 VSUBS 0.013639f
C879 VTAIL.n722 VSUBS 0.012881f
C880 VTAIL.n723 VSUBS 0.023971f
C881 VTAIL.n724 VSUBS 0.023971f
C882 VTAIL.n725 VSUBS 0.012881f
C883 VTAIL.n726 VSUBS 0.013639f
C884 VTAIL.n727 VSUBS 0.030446f
C885 VTAIL.n728 VSUBS 0.030446f
C886 VTAIL.n729 VSUBS 0.013639f
C887 VTAIL.n730 VSUBS 0.012881f
C888 VTAIL.n731 VSUBS 0.023971f
C889 VTAIL.n732 VSUBS 0.023971f
C890 VTAIL.n733 VSUBS 0.012881f
C891 VTAIL.n734 VSUBS 0.013639f
C892 VTAIL.n735 VSUBS 0.030446f
C893 VTAIL.n736 VSUBS 0.030446f
C894 VTAIL.n737 VSUBS 0.013639f
C895 VTAIL.n738 VSUBS 0.012881f
C896 VTAIL.n739 VSUBS 0.023971f
C897 VTAIL.n740 VSUBS 0.023971f
C898 VTAIL.n741 VSUBS 0.012881f
C899 VTAIL.n742 VSUBS 0.013639f
C900 VTAIL.n743 VSUBS 0.030446f
C901 VTAIL.n744 VSUBS 0.074904f
C902 VTAIL.n745 VSUBS 0.013639f
C903 VTAIL.n746 VSUBS 0.025295f
C904 VTAIL.n747 VSUBS 0.059337f
C905 VTAIL.n748 VSUBS 0.056987f
C906 VTAIL.n749 VSUBS 2.18342f
C907 VTAIL.n750 VSUBS 0.025427f
C908 VTAIL.n751 VSUBS 0.023971f
C909 VTAIL.n752 VSUBS 0.012881f
C910 VTAIL.n753 VSUBS 0.030446f
C911 VTAIL.n754 VSUBS 0.013639f
C912 VTAIL.n755 VSUBS 0.023971f
C913 VTAIL.n756 VSUBS 0.012881f
C914 VTAIL.n757 VSUBS 0.030446f
C915 VTAIL.n758 VSUBS 0.013639f
C916 VTAIL.n759 VSUBS 0.023971f
C917 VTAIL.n760 VSUBS 0.012881f
C918 VTAIL.n761 VSUBS 0.030446f
C919 VTAIL.n762 VSUBS 0.013639f
C920 VTAIL.n763 VSUBS 0.023971f
C921 VTAIL.n764 VSUBS 0.012881f
C922 VTAIL.n765 VSUBS 0.030446f
C923 VTAIL.n766 VSUBS 0.013639f
C924 VTAIL.n767 VSUBS 0.023971f
C925 VTAIL.n768 VSUBS 0.012881f
C926 VTAIL.n769 VSUBS 0.030446f
C927 VTAIL.n770 VSUBS 0.013639f
C928 VTAIL.n771 VSUBS 0.023971f
C929 VTAIL.n772 VSUBS 0.012881f
C930 VTAIL.n773 VSUBS 0.030446f
C931 VTAIL.n774 VSUBS 0.013639f
C932 VTAIL.n775 VSUBS 0.023971f
C933 VTAIL.n776 VSUBS 0.012881f
C934 VTAIL.n777 VSUBS 0.030446f
C935 VTAIL.n778 VSUBS 0.013639f
C936 VTAIL.n779 VSUBS 0.023971f
C937 VTAIL.n780 VSUBS 0.012881f
C938 VTAIL.n781 VSUBS 0.030446f
C939 VTAIL.n782 VSUBS 0.013639f
C940 VTAIL.n783 VSUBS 0.269424f
C941 VTAIL.t11 VSUBS 0.06621f
C942 VTAIL.n784 VSUBS 0.022834f
C943 VTAIL.n785 VSUBS 0.022903f
C944 VTAIL.n786 VSUBS 0.012881f
C945 VTAIL.n787 VSUBS 1.9592f
C946 VTAIL.n788 VSUBS 0.023971f
C947 VTAIL.n789 VSUBS 0.012881f
C948 VTAIL.n790 VSUBS 0.013639f
C949 VTAIL.n791 VSUBS 0.030446f
C950 VTAIL.n792 VSUBS 0.030446f
C951 VTAIL.n793 VSUBS 0.013639f
C952 VTAIL.n794 VSUBS 0.012881f
C953 VTAIL.n795 VSUBS 0.023971f
C954 VTAIL.n796 VSUBS 0.023971f
C955 VTAIL.n797 VSUBS 0.012881f
C956 VTAIL.n798 VSUBS 0.013639f
C957 VTAIL.n799 VSUBS 0.030446f
C958 VTAIL.n800 VSUBS 0.030446f
C959 VTAIL.n801 VSUBS 0.030446f
C960 VTAIL.n802 VSUBS 0.013639f
C961 VTAIL.n803 VSUBS 0.012881f
C962 VTAIL.n804 VSUBS 0.023971f
C963 VTAIL.n805 VSUBS 0.023971f
C964 VTAIL.n806 VSUBS 0.012881f
C965 VTAIL.n807 VSUBS 0.01326f
C966 VTAIL.n808 VSUBS 0.01326f
C967 VTAIL.n809 VSUBS 0.030446f
C968 VTAIL.n810 VSUBS 0.030446f
C969 VTAIL.n811 VSUBS 0.013639f
C970 VTAIL.n812 VSUBS 0.012881f
C971 VTAIL.n813 VSUBS 0.023971f
C972 VTAIL.n814 VSUBS 0.023971f
C973 VTAIL.n815 VSUBS 0.012881f
C974 VTAIL.n816 VSUBS 0.013639f
C975 VTAIL.n817 VSUBS 0.030446f
C976 VTAIL.n818 VSUBS 0.030446f
C977 VTAIL.n819 VSUBS 0.013639f
C978 VTAIL.n820 VSUBS 0.012881f
C979 VTAIL.n821 VSUBS 0.023971f
C980 VTAIL.n822 VSUBS 0.023971f
C981 VTAIL.n823 VSUBS 0.012881f
C982 VTAIL.n824 VSUBS 0.013639f
C983 VTAIL.n825 VSUBS 0.030446f
C984 VTAIL.n826 VSUBS 0.030446f
C985 VTAIL.n827 VSUBS 0.013639f
C986 VTAIL.n828 VSUBS 0.012881f
C987 VTAIL.n829 VSUBS 0.023971f
C988 VTAIL.n830 VSUBS 0.023971f
C989 VTAIL.n831 VSUBS 0.012881f
C990 VTAIL.n832 VSUBS 0.013639f
C991 VTAIL.n833 VSUBS 0.030446f
C992 VTAIL.n834 VSUBS 0.030446f
C993 VTAIL.n835 VSUBS 0.013639f
C994 VTAIL.n836 VSUBS 0.012881f
C995 VTAIL.n837 VSUBS 0.023971f
C996 VTAIL.n838 VSUBS 0.023971f
C997 VTAIL.n839 VSUBS 0.012881f
C998 VTAIL.n840 VSUBS 0.013639f
C999 VTAIL.n841 VSUBS 0.030446f
C1000 VTAIL.n842 VSUBS 0.030446f
C1001 VTAIL.n843 VSUBS 0.013639f
C1002 VTAIL.n844 VSUBS 0.012881f
C1003 VTAIL.n845 VSUBS 0.023971f
C1004 VTAIL.n846 VSUBS 0.023971f
C1005 VTAIL.n847 VSUBS 0.012881f
C1006 VTAIL.n848 VSUBS 0.013639f
C1007 VTAIL.n849 VSUBS 0.030446f
C1008 VTAIL.n850 VSUBS 0.074904f
C1009 VTAIL.n851 VSUBS 0.013639f
C1010 VTAIL.n852 VSUBS 0.025295f
C1011 VTAIL.n853 VSUBS 0.059337f
C1012 VTAIL.n854 VSUBS 0.056987f
C1013 VTAIL.n855 VSUBS 2.17892f
C1014 VP.t5 VSUBS 4.447f
C1015 VP.n0 VSUBS 1.61328f
C1016 VP.n1 VSUBS 0.022265f
C1017 VP.n2 VSUBS 0.042681f
C1018 VP.n3 VSUBS 0.022265f
C1019 VP.n4 VSUBS 0.04047f
C1020 VP.n5 VSUBS 0.022265f
C1021 VP.n6 VSUBS 0.044489f
C1022 VP.n7 VSUBS 0.022265f
C1023 VP.n8 VSUBS 0.041705f
C1024 VP.n9 VSUBS 0.022265f
C1025 VP.t3 VSUBS 4.447f
C1026 VP.n10 VSUBS 0.045238f
C1027 VP.n11 VSUBS 0.022265f
C1028 VP.n12 VSUBS 0.041705f
C1029 VP.t0 VSUBS 4.447f
C1030 VP.n13 VSUBS 1.61328f
C1031 VP.n14 VSUBS 0.022265f
C1032 VP.n15 VSUBS 0.042681f
C1033 VP.n16 VSUBS 0.022265f
C1034 VP.n17 VSUBS 0.04047f
C1035 VP.n18 VSUBS 0.022265f
C1036 VP.n19 VSUBS 0.044489f
C1037 VP.n20 VSUBS 0.022265f
C1038 VP.n21 VSUBS 0.041705f
C1039 VP.t2 VSUBS 4.79368f
C1040 VP.n22 VSUBS 1.53541f
C1041 VP.t7 VSUBS 4.447f
C1042 VP.n23 VSUBS 1.60036f
C1043 VP.n24 VSUBS 0.022349f
C1044 VP.n25 VSUBS 0.283626f
C1045 VP.n26 VSUBS 0.022265f
C1046 VP.n27 VSUBS 0.022265f
C1047 VP.n28 VSUBS 0.041705f
C1048 VP.n29 VSUBS 0.044489f
C1049 VP.n30 VSUBS 0.018018f
C1050 VP.n31 VSUBS 0.022265f
C1051 VP.n32 VSUBS 0.022265f
C1052 VP.n33 VSUBS 0.022265f
C1053 VP.n34 VSUBS 0.041705f
C1054 VP.n35 VSUBS 0.041705f
C1055 VP.t4 VSUBS 4.447f
C1056 VP.n36 VSUBS 1.52878f
C1057 VP.n37 VSUBS 0.022349f
C1058 VP.n38 VSUBS 0.022265f
C1059 VP.n39 VSUBS 0.022265f
C1060 VP.n40 VSUBS 0.022265f
C1061 VP.n41 VSUBS 0.041705f
C1062 VP.n42 VSUBS 0.045238f
C1063 VP.n43 VSUBS 0.019077f
C1064 VP.n44 VSUBS 0.022265f
C1065 VP.n45 VSUBS 0.022265f
C1066 VP.n46 VSUBS 0.022265f
C1067 VP.n47 VSUBS 0.041705f
C1068 VP.n48 VSUBS 0.041705f
C1069 VP.n49 VSUBS 0.02482f
C1070 VP.n50 VSUBS 0.035942f
C1071 VP.n51 VSUBS 1.71158f
C1072 VP.n52 VSUBS 1.72448f
C1073 VP.t6 VSUBS 4.447f
C1074 VP.n53 VSUBS 1.61328f
C1075 VP.n54 VSUBS 0.02482f
C1076 VP.n55 VSUBS 0.035942f
C1077 VP.n56 VSUBS 0.022265f
C1078 VP.n57 VSUBS 0.022265f
C1079 VP.n58 VSUBS 0.041705f
C1080 VP.n59 VSUBS 0.042681f
C1081 VP.n60 VSUBS 0.019077f
C1082 VP.n61 VSUBS 0.022265f
C1083 VP.n62 VSUBS 0.022265f
C1084 VP.n63 VSUBS 0.022265f
C1085 VP.n64 VSUBS 0.041705f
C1086 VP.n65 VSUBS 0.04047f
C1087 VP.n66 VSUBS 1.52878f
C1088 VP.n67 VSUBS 0.022349f
C1089 VP.n68 VSUBS 0.022265f
C1090 VP.n69 VSUBS 0.022265f
C1091 VP.n70 VSUBS 0.022265f
C1092 VP.n71 VSUBS 0.041705f
C1093 VP.n72 VSUBS 0.044489f
C1094 VP.n73 VSUBS 0.018018f
C1095 VP.n74 VSUBS 0.022265f
C1096 VP.n75 VSUBS 0.022265f
C1097 VP.n76 VSUBS 0.022265f
C1098 VP.n77 VSUBS 0.041705f
C1099 VP.n78 VSUBS 0.041705f
C1100 VP.t1 VSUBS 4.447f
C1101 VP.n79 VSUBS 1.52878f
C1102 VP.n80 VSUBS 0.022349f
C1103 VP.n81 VSUBS 0.022265f
C1104 VP.n82 VSUBS 0.022265f
C1105 VP.n83 VSUBS 0.022265f
C1106 VP.n84 VSUBS 0.041705f
C1107 VP.n85 VSUBS 0.045238f
C1108 VP.n86 VSUBS 0.019077f
C1109 VP.n87 VSUBS 0.022265f
C1110 VP.n88 VSUBS 0.022265f
C1111 VP.n89 VSUBS 0.022265f
C1112 VP.n90 VSUBS 0.041705f
C1113 VP.n91 VSUBS 0.041705f
C1114 VP.n92 VSUBS 0.02482f
C1115 VP.n93 VSUBS 0.035942f
C1116 VP.n94 VSUBS 0.066615f
C1117 B.n0 VSUBS 0.00453f
C1118 B.n1 VSUBS 0.00453f
C1119 B.n2 VSUBS 0.007164f
C1120 B.n3 VSUBS 0.007164f
C1121 B.n4 VSUBS 0.007164f
C1122 B.n5 VSUBS 0.007164f
C1123 B.n6 VSUBS 0.007164f
C1124 B.n7 VSUBS 0.007164f
C1125 B.n8 VSUBS 0.007164f
C1126 B.n9 VSUBS 0.007164f
C1127 B.n10 VSUBS 0.007164f
C1128 B.n11 VSUBS 0.007164f
C1129 B.n12 VSUBS 0.007164f
C1130 B.n13 VSUBS 0.007164f
C1131 B.n14 VSUBS 0.007164f
C1132 B.n15 VSUBS 0.007164f
C1133 B.n16 VSUBS 0.007164f
C1134 B.n17 VSUBS 0.007164f
C1135 B.n18 VSUBS 0.007164f
C1136 B.n19 VSUBS 0.007164f
C1137 B.n20 VSUBS 0.007164f
C1138 B.n21 VSUBS 0.007164f
C1139 B.n22 VSUBS 0.007164f
C1140 B.n23 VSUBS 0.007164f
C1141 B.n24 VSUBS 0.007164f
C1142 B.n25 VSUBS 0.007164f
C1143 B.n26 VSUBS 0.007164f
C1144 B.n27 VSUBS 0.007164f
C1145 B.n28 VSUBS 0.007164f
C1146 B.n29 VSUBS 0.007164f
C1147 B.n30 VSUBS 0.007164f
C1148 B.n31 VSUBS 0.007164f
C1149 B.n32 VSUBS 0.007164f
C1150 B.n33 VSUBS 0.007164f
C1151 B.n34 VSUBS 0.007164f
C1152 B.n35 VSUBS 0.007164f
C1153 B.n36 VSUBS 0.015764f
C1154 B.n37 VSUBS 0.007164f
C1155 B.n38 VSUBS 0.007164f
C1156 B.n39 VSUBS 0.007164f
C1157 B.n40 VSUBS 0.007164f
C1158 B.n41 VSUBS 0.007164f
C1159 B.n42 VSUBS 0.007164f
C1160 B.n43 VSUBS 0.007164f
C1161 B.n44 VSUBS 0.007164f
C1162 B.n45 VSUBS 0.007164f
C1163 B.n46 VSUBS 0.007164f
C1164 B.n47 VSUBS 0.007164f
C1165 B.n48 VSUBS 0.007164f
C1166 B.n49 VSUBS 0.007164f
C1167 B.n50 VSUBS 0.007164f
C1168 B.n51 VSUBS 0.007164f
C1169 B.n52 VSUBS 0.007164f
C1170 B.n53 VSUBS 0.007164f
C1171 B.n54 VSUBS 0.007164f
C1172 B.n55 VSUBS 0.007164f
C1173 B.n56 VSUBS 0.007164f
C1174 B.n57 VSUBS 0.007164f
C1175 B.n58 VSUBS 0.007164f
C1176 B.n59 VSUBS 0.007164f
C1177 B.n60 VSUBS 0.007164f
C1178 B.n61 VSUBS 0.007164f
C1179 B.n62 VSUBS 0.007164f
C1180 B.n63 VSUBS 0.007164f
C1181 B.n64 VSUBS 0.007164f
C1182 B.n65 VSUBS 0.007164f
C1183 B.n66 VSUBS 0.007164f
C1184 B.n67 VSUBS 0.007164f
C1185 B.t11 VSUBS 0.394974f
C1186 B.t10 VSUBS 0.44163f
C1187 B.t9 VSUBS 3.36082f
C1188 B.n68 VSUBS 0.707321f
C1189 B.n69 VSUBS 0.358767f
C1190 B.n70 VSUBS 0.016597f
C1191 B.n71 VSUBS 0.007164f
C1192 B.n72 VSUBS 0.007164f
C1193 B.n73 VSUBS 0.007164f
C1194 B.n74 VSUBS 0.007164f
C1195 B.n75 VSUBS 0.007164f
C1196 B.t8 VSUBS 0.394977f
C1197 B.t7 VSUBS 0.441633f
C1198 B.t6 VSUBS 3.36082f
C1199 B.n76 VSUBS 0.707317f
C1200 B.n77 VSUBS 0.358763f
C1201 B.n78 VSUBS 0.007164f
C1202 B.n79 VSUBS 0.007164f
C1203 B.n80 VSUBS 0.007164f
C1204 B.n81 VSUBS 0.007164f
C1205 B.n82 VSUBS 0.007164f
C1206 B.n83 VSUBS 0.007164f
C1207 B.n84 VSUBS 0.007164f
C1208 B.n85 VSUBS 0.007164f
C1209 B.n86 VSUBS 0.007164f
C1210 B.n87 VSUBS 0.007164f
C1211 B.n88 VSUBS 0.007164f
C1212 B.n89 VSUBS 0.007164f
C1213 B.n90 VSUBS 0.007164f
C1214 B.n91 VSUBS 0.007164f
C1215 B.n92 VSUBS 0.007164f
C1216 B.n93 VSUBS 0.007164f
C1217 B.n94 VSUBS 0.007164f
C1218 B.n95 VSUBS 0.007164f
C1219 B.n96 VSUBS 0.007164f
C1220 B.n97 VSUBS 0.007164f
C1221 B.n98 VSUBS 0.007164f
C1222 B.n99 VSUBS 0.007164f
C1223 B.n100 VSUBS 0.007164f
C1224 B.n101 VSUBS 0.007164f
C1225 B.n102 VSUBS 0.007164f
C1226 B.n103 VSUBS 0.007164f
C1227 B.n104 VSUBS 0.007164f
C1228 B.n105 VSUBS 0.007164f
C1229 B.n106 VSUBS 0.007164f
C1230 B.n107 VSUBS 0.007164f
C1231 B.n108 VSUBS 0.007164f
C1232 B.n109 VSUBS 0.014786f
C1233 B.n110 VSUBS 0.007164f
C1234 B.n111 VSUBS 0.007164f
C1235 B.n112 VSUBS 0.007164f
C1236 B.n113 VSUBS 0.007164f
C1237 B.n114 VSUBS 0.007164f
C1238 B.n115 VSUBS 0.007164f
C1239 B.n116 VSUBS 0.007164f
C1240 B.n117 VSUBS 0.007164f
C1241 B.n118 VSUBS 0.007164f
C1242 B.n119 VSUBS 0.007164f
C1243 B.n120 VSUBS 0.007164f
C1244 B.n121 VSUBS 0.007164f
C1245 B.n122 VSUBS 0.007164f
C1246 B.n123 VSUBS 0.007164f
C1247 B.n124 VSUBS 0.007164f
C1248 B.n125 VSUBS 0.007164f
C1249 B.n126 VSUBS 0.007164f
C1250 B.n127 VSUBS 0.007164f
C1251 B.n128 VSUBS 0.007164f
C1252 B.n129 VSUBS 0.007164f
C1253 B.n130 VSUBS 0.007164f
C1254 B.n131 VSUBS 0.007164f
C1255 B.n132 VSUBS 0.007164f
C1256 B.n133 VSUBS 0.007164f
C1257 B.n134 VSUBS 0.007164f
C1258 B.n135 VSUBS 0.007164f
C1259 B.n136 VSUBS 0.007164f
C1260 B.n137 VSUBS 0.007164f
C1261 B.n138 VSUBS 0.007164f
C1262 B.n139 VSUBS 0.007164f
C1263 B.n140 VSUBS 0.007164f
C1264 B.n141 VSUBS 0.007164f
C1265 B.n142 VSUBS 0.007164f
C1266 B.n143 VSUBS 0.007164f
C1267 B.n144 VSUBS 0.007164f
C1268 B.n145 VSUBS 0.007164f
C1269 B.n146 VSUBS 0.007164f
C1270 B.n147 VSUBS 0.007164f
C1271 B.n148 VSUBS 0.007164f
C1272 B.n149 VSUBS 0.007164f
C1273 B.n150 VSUBS 0.007164f
C1274 B.n151 VSUBS 0.007164f
C1275 B.n152 VSUBS 0.007164f
C1276 B.n153 VSUBS 0.007164f
C1277 B.n154 VSUBS 0.007164f
C1278 B.n155 VSUBS 0.007164f
C1279 B.n156 VSUBS 0.007164f
C1280 B.n157 VSUBS 0.007164f
C1281 B.n158 VSUBS 0.007164f
C1282 B.n159 VSUBS 0.007164f
C1283 B.n160 VSUBS 0.007164f
C1284 B.n161 VSUBS 0.007164f
C1285 B.n162 VSUBS 0.007164f
C1286 B.n163 VSUBS 0.007164f
C1287 B.n164 VSUBS 0.007164f
C1288 B.n165 VSUBS 0.007164f
C1289 B.n166 VSUBS 0.007164f
C1290 B.n167 VSUBS 0.007164f
C1291 B.n168 VSUBS 0.007164f
C1292 B.n169 VSUBS 0.007164f
C1293 B.n170 VSUBS 0.007164f
C1294 B.n171 VSUBS 0.007164f
C1295 B.n172 VSUBS 0.007164f
C1296 B.n173 VSUBS 0.007164f
C1297 B.n174 VSUBS 0.007164f
C1298 B.n175 VSUBS 0.007164f
C1299 B.n176 VSUBS 0.007164f
C1300 B.n177 VSUBS 0.014786f
C1301 B.n178 VSUBS 0.007164f
C1302 B.n179 VSUBS 0.007164f
C1303 B.n180 VSUBS 0.007164f
C1304 B.n181 VSUBS 0.007164f
C1305 B.n182 VSUBS 0.007164f
C1306 B.n183 VSUBS 0.007164f
C1307 B.n184 VSUBS 0.007164f
C1308 B.n185 VSUBS 0.007164f
C1309 B.n186 VSUBS 0.007164f
C1310 B.n187 VSUBS 0.007164f
C1311 B.n188 VSUBS 0.007164f
C1312 B.n189 VSUBS 0.007164f
C1313 B.n190 VSUBS 0.007164f
C1314 B.n191 VSUBS 0.007164f
C1315 B.n192 VSUBS 0.007164f
C1316 B.n193 VSUBS 0.007164f
C1317 B.n194 VSUBS 0.007164f
C1318 B.n195 VSUBS 0.007164f
C1319 B.n196 VSUBS 0.007164f
C1320 B.n197 VSUBS 0.007164f
C1321 B.n198 VSUBS 0.007164f
C1322 B.n199 VSUBS 0.007164f
C1323 B.n200 VSUBS 0.007164f
C1324 B.n201 VSUBS 0.007164f
C1325 B.n202 VSUBS 0.007164f
C1326 B.n203 VSUBS 0.007164f
C1327 B.n204 VSUBS 0.007164f
C1328 B.n205 VSUBS 0.007164f
C1329 B.n206 VSUBS 0.007164f
C1330 B.n207 VSUBS 0.007164f
C1331 B.n208 VSUBS 0.007164f
C1332 B.n209 VSUBS 0.007164f
C1333 B.t4 VSUBS 0.394977f
C1334 B.t5 VSUBS 0.441633f
C1335 B.t3 VSUBS 3.36082f
C1336 B.n210 VSUBS 0.707317f
C1337 B.n211 VSUBS 0.358763f
C1338 B.n212 VSUBS 0.007164f
C1339 B.n213 VSUBS 0.007164f
C1340 B.n214 VSUBS 0.007164f
C1341 B.n215 VSUBS 0.007164f
C1342 B.t1 VSUBS 0.394974f
C1343 B.t2 VSUBS 0.44163f
C1344 B.t0 VSUBS 3.36082f
C1345 B.n216 VSUBS 0.707321f
C1346 B.n217 VSUBS 0.358767f
C1347 B.n218 VSUBS 0.016597f
C1348 B.n219 VSUBS 0.007164f
C1349 B.n220 VSUBS 0.007164f
C1350 B.n221 VSUBS 0.007164f
C1351 B.n222 VSUBS 0.007164f
C1352 B.n223 VSUBS 0.007164f
C1353 B.n224 VSUBS 0.007164f
C1354 B.n225 VSUBS 0.007164f
C1355 B.n226 VSUBS 0.007164f
C1356 B.n227 VSUBS 0.007164f
C1357 B.n228 VSUBS 0.007164f
C1358 B.n229 VSUBS 0.007164f
C1359 B.n230 VSUBS 0.007164f
C1360 B.n231 VSUBS 0.007164f
C1361 B.n232 VSUBS 0.007164f
C1362 B.n233 VSUBS 0.007164f
C1363 B.n234 VSUBS 0.007164f
C1364 B.n235 VSUBS 0.007164f
C1365 B.n236 VSUBS 0.007164f
C1366 B.n237 VSUBS 0.007164f
C1367 B.n238 VSUBS 0.007164f
C1368 B.n239 VSUBS 0.007164f
C1369 B.n240 VSUBS 0.007164f
C1370 B.n241 VSUBS 0.007164f
C1371 B.n242 VSUBS 0.007164f
C1372 B.n243 VSUBS 0.007164f
C1373 B.n244 VSUBS 0.007164f
C1374 B.n245 VSUBS 0.007164f
C1375 B.n246 VSUBS 0.007164f
C1376 B.n247 VSUBS 0.007164f
C1377 B.n248 VSUBS 0.007164f
C1378 B.n249 VSUBS 0.007164f
C1379 B.n250 VSUBS 0.015764f
C1380 B.n251 VSUBS 0.007164f
C1381 B.n252 VSUBS 0.007164f
C1382 B.n253 VSUBS 0.007164f
C1383 B.n254 VSUBS 0.007164f
C1384 B.n255 VSUBS 0.007164f
C1385 B.n256 VSUBS 0.007164f
C1386 B.n257 VSUBS 0.007164f
C1387 B.n258 VSUBS 0.007164f
C1388 B.n259 VSUBS 0.007164f
C1389 B.n260 VSUBS 0.007164f
C1390 B.n261 VSUBS 0.007164f
C1391 B.n262 VSUBS 0.007164f
C1392 B.n263 VSUBS 0.007164f
C1393 B.n264 VSUBS 0.007164f
C1394 B.n265 VSUBS 0.007164f
C1395 B.n266 VSUBS 0.007164f
C1396 B.n267 VSUBS 0.007164f
C1397 B.n268 VSUBS 0.007164f
C1398 B.n269 VSUBS 0.007164f
C1399 B.n270 VSUBS 0.007164f
C1400 B.n271 VSUBS 0.007164f
C1401 B.n272 VSUBS 0.007164f
C1402 B.n273 VSUBS 0.007164f
C1403 B.n274 VSUBS 0.007164f
C1404 B.n275 VSUBS 0.007164f
C1405 B.n276 VSUBS 0.007164f
C1406 B.n277 VSUBS 0.007164f
C1407 B.n278 VSUBS 0.007164f
C1408 B.n279 VSUBS 0.007164f
C1409 B.n280 VSUBS 0.007164f
C1410 B.n281 VSUBS 0.007164f
C1411 B.n282 VSUBS 0.007164f
C1412 B.n283 VSUBS 0.007164f
C1413 B.n284 VSUBS 0.007164f
C1414 B.n285 VSUBS 0.007164f
C1415 B.n286 VSUBS 0.007164f
C1416 B.n287 VSUBS 0.007164f
C1417 B.n288 VSUBS 0.007164f
C1418 B.n289 VSUBS 0.007164f
C1419 B.n290 VSUBS 0.007164f
C1420 B.n291 VSUBS 0.007164f
C1421 B.n292 VSUBS 0.007164f
C1422 B.n293 VSUBS 0.007164f
C1423 B.n294 VSUBS 0.007164f
C1424 B.n295 VSUBS 0.007164f
C1425 B.n296 VSUBS 0.007164f
C1426 B.n297 VSUBS 0.007164f
C1427 B.n298 VSUBS 0.007164f
C1428 B.n299 VSUBS 0.007164f
C1429 B.n300 VSUBS 0.007164f
C1430 B.n301 VSUBS 0.007164f
C1431 B.n302 VSUBS 0.007164f
C1432 B.n303 VSUBS 0.007164f
C1433 B.n304 VSUBS 0.007164f
C1434 B.n305 VSUBS 0.007164f
C1435 B.n306 VSUBS 0.007164f
C1436 B.n307 VSUBS 0.007164f
C1437 B.n308 VSUBS 0.007164f
C1438 B.n309 VSUBS 0.007164f
C1439 B.n310 VSUBS 0.007164f
C1440 B.n311 VSUBS 0.007164f
C1441 B.n312 VSUBS 0.007164f
C1442 B.n313 VSUBS 0.007164f
C1443 B.n314 VSUBS 0.007164f
C1444 B.n315 VSUBS 0.007164f
C1445 B.n316 VSUBS 0.007164f
C1446 B.n317 VSUBS 0.007164f
C1447 B.n318 VSUBS 0.007164f
C1448 B.n319 VSUBS 0.007164f
C1449 B.n320 VSUBS 0.007164f
C1450 B.n321 VSUBS 0.007164f
C1451 B.n322 VSUBS 0.007164f
C1452 B.n323 VSUBS 0.007164f
C1453 B.n324 VSUBS 0.007164f
C1454 B.n325 VSUBS 0.007164f
C1455 B.n326 VSUBS 0.007164f
C1456 B.n327 VSUBS 0.007164f
C1457 B.n328 VSUBS 0.007164f
C1458 B.n329 VSUBS 0.007164f
C1459 B.n330 VSUBS 0.007164f
C1460 B.n331 VSUBS 0.007164f
C1461 B.n332 VSUBS 0.007164f
C1462 B.n333 VSUBS 0.007164f
C1463 B.n334 VSUBS 0.007164f
C1464 B.n335 VSUBS 0.007164f
C1465 B.n336 VSUBS 0.007164f
C1466 B.n337 VSUBS 0.007164f
C1467 B.n338 VSUBS 0.007164f
C1468 B.n339 VSUBS 0.007164f
C1469 B.n340 VSUBS 0.007164f
C1470 B.n341 VSUBS 0.007164f
C1471 B.n342 VSUBS 0.007164f
C1472 B.n343 VSUBS 0.007164f
C1473 B.n344 VSUBS 0.007164f
C1474 B.n345 VSUBS 0.007164f
C1475 B.n346 VSUBS 0.007164f
C1476 B.n347 VSUBS 0.007164f
C1477 B.n348 VSUBS 0.007164f
C1478 B.n349 VSUBS 0.007164f
C1479 B.n350 VSUBS 0.007164f
C1480 B.n351 VSUBS 0.007164f
C1481 B.n352 VSUBS 0.007164f
C1482 B.n353 VSUBS 0.007164f
C1483 B.n354 VSUBS 0.007164f
C1484 B.n355 VSUBS 0.007164f
C1485 B.n356 VSUBS 0.007164f
C1486 B.n357 VSUBS 0.007164f
C1487 B.n358 VSUBS 0.007164f
C1488 B.n359 VSUBS 0.007164f
C1489 B.n360 VSUBS 0.007164f
C1490 B.n361 VSUBS 0.007164f
C1491 B.n362 VSUBS 0.007164f
C1492 B.n363 VSUBS 0.007164f
C1493 B.n364 VSUBS 0.007164f
C1494 B.n365 VSUBS 0.007164f
C1495 B.n366 VSUBS 0.007164f
C1496 B.n367 VSUBS 0.007164f
C1497 B.n368 VSUBS 0.007164f
C1498 B.n369 VSUBS 0.007164f
C1499 B.n370 VSUBS 0.007164f
C1500 B.n371 VSUBS 0.007164f
C1501 B.n372 VSUBS 0.007164f
C1502 B.n373 VSUBS 0.007164f
C1503 B.n374 VSUBS 0.007164f
C1504 B.n375 VSUBS 0.007164f
C1505 B.n376 VSUBS 0.007164f
C1506 B.n377 VSUBS 0.007164f
C1507 B.n378 VSUBS 0.007164f
C1508 B.n379 VSUBS 0.007164f
C1509 B.n380 VSUBS 0.007164f
C1510 B.n381 VSUBS 0.007164f
C1511 B.n382 VSUBS 0.007164f
C1512 B.n383 VSUBS 0.014786f
C1513 B.n384 VSUBS 0.014786f
C1514 B.n385 VSUBS 0.015764f
C1515 B.n386 VSUBS 0.007164f
C1516 B.n387 VSUBS 0.007164f
C1517 B.n388 VSUBS 0.007164f
C1518 B.n389 VSUBS 0.007164f
C1519 B.n390 VSUBS 0.007164f
C1520 B.n391 VSUBS 0.007164f
C1521 B.n392 VSUBS 0.007164f
C1522 B.n393 VSUBS 0.007164f
C1523 B.n394 VSUBS 0.007164f
C1524 B.n395 VSUBS 0.007164f
C1525 B.n396 VSUBS 0.007164f
C1526 B.n397 VSUBS 0.007164f
C1527 B.n398 VSUBS 0.007164f
C1528 B.n399 VSUBS 0.007164f
C1529 B.n400 VSUBS 0.007164f
C1530 B.n401 VSUBS 0.007164f
C1531 B.n402 VSUBS 0.007164f
C1532 B.n403 VSUBS 0.007164f
C1533 B.n404 VSUBS 0.007164f
C1534 B.n405 VSUBS 0.007164f
C1535 B.n406 VSUBS 0.007164f
C1536 B.n407 VSUBS 0.007164f
C1537 B.n408 VSUBS 0.007164f
C1538 B.n409 VSUBS 0.007164f
C1539 B.n410 VSUBS 0.007164f
C1540 B.n411 VSUBS 0.007164f
C1541 B.n412 VSUBS 0.007164f
C1542 B.n413 VSUBS 0.007164f
C1543 B.n414 VSUBS 0.007164f
C1544 B.n415 VSUBS 0.007164f
C1545 B.n416 VSUBS 0.007164f
C1546 B.n417 VSUBS 0.007164f
C1547 B.n418 VSUBS 0.007164f
C1548 B.n419 VSUBS 0.007164f
C1549 B.n420 VSUBS 0.007164f
C1550 B.n421 VSUBS 0.007164f
C1551 B.n422 VSUBS 0.007164f
C1552 B.n423 VSUBS 0.007164f
C1553 B.n424 VSUBS 0.007164f
C1554 B.n425 VSUBS 0.007164f
C1555 B.n426 VSUBS 0.007164f
C1556 B.n427 VSUBS 0.007164f
C1557 B.n428 VSUBS 0.007164f
C1558 B.n429 VSUBS 0.007164f
C1559 B.n430 VSUBS 0.007164f
C1560 B.n431 VSUBS 0.007164f
C1561 B.n432 VSUBS 0.007164f
C1562 B.n433 VSUBS 0.007164f
C1563 B.n434 VSUBS 0.007164f
C1564 B.n435 VSUBS 0.007164f
C1565 B.n436 VSUBS 0.007164f
C1566 B.n437 VSUBS 0.007164f
C1567 B.n438 VSUBS 0.007164f
C1568 B.n439 VSUBS 0.007164f
C1569 B.n440 VSUBS 0.007164f
C1570 B.n441 VSUBS 0.007164f
C1571 B.n442 VSUBS 0.007164f
C1572 B.n443 VSUBS 0.007164f
C1573 B.n444 VSUBS 0.007164f
C1574 B.n445 VSUBS 0.007164f
C1575 B.n446 VSUBS 0.007164f
C1576 B.n447 VSUBS 0.007164f
C1577 B.n448 VSUBS 0.007164f
C1578 B.n449 VSUBS 0.007164f
C1579 B.n450 VSUBS 0.007164f
C1580 B.n451 VSUBS 0.007164f
C1581 B.n452 VSUBS 0.007164f
C1582 B.n453 VSUBS 0.007164f
C1583 B.n454 VSUBS 0.007164f
C1584 B.n455 VSUBS 0.007164f
C1585 B.n456 VSUBS 0.007164f
C1586 B.n457 VSUBS 0.007164f
C1587 B.n458 VSUBS 0.007164f
C1588 B.n459 VSUBS 0.007164f
C1589 B.n460 VSUBS 0.007164f
C1590 B.n461 VSUBS 0.007164f
C1591 B.n462 VSUBS 0.007164f
C1592 B.n463 VSUBS 0.007164f
C1593 B.n464 VSUBS 0.007164f
C1594 B.n465 VSUBS 0.007164f
C1595 B.n466 VSUBS 0.007164f
C1596 B.n467 VSUBS 0.007164f
C1597 B.n468 VSUBS 0.007164f
C1598 B.n469 VSUBS 0.007164f
C1599 B.n470 VSUBS 0.007164f
C1600 B.n471 VSUBS 0.007164f
C1601 B.n472 VSUBS 0.007164f
C1602 B.n473 VSUBS 0.007164f
C1603 B.n474 VSUBS 0.007164f
C1604 B.n475 VSUBS 0.007164f
C1605 B.n476 VSUBS 0.007164f
C1606 B.n477 VSUBS 0.007164f
C1607 B.n478 VSUBS 0.007164f
C1608 B.n479 VSUBS 0.004951f
C1609 B.n480 VSUBS 0.007164f
C1610 B.n481 VSUBS 0.007164f
C1611 B.n482 VSUBS 0.005794f
C1612 B.n483 VSUBS 0.007164f
C1613 B.n484 VSUBS 0.007164f
C1614 B.n485 VSUBS 0.007164f
C1615 B.n486 VSUBS 0.007164f
C1616 B.n487 VSUBS 0.007164f
C1617 B.n488 VSUBS 0.007164f
C1618 B.n489 VSUBS 0.007164f
C1619 B.n490 VSUBS 0.007164f
C1620 B.n491 VSUBS 0.007164f
C1621 B.n492 VSUBS 0.007164f
C1622 B.n493 VSUBS 0.007164f
C1623 B.n494 VSUBS 0.005794f
C1624 B.n495 VSUBS 0.016597f
C1625 B.n496 VSUBS 0.004951f
C1626 B.n497 VSUBS 0.007164f
C1627 B.n498 VSUBS 0.007164f
C1628 B.n499 VSUBS 0.007164f
C1629 B.n500 VSUBS 0.007164f
C1630 B.n501 VSUBS 0.007164f
C1631 B.n502 VSUBS 0.007164f
C1632 B.n503 VSUBS 0.007164f
C1633 B.n504 VSUBS 0.007164f
C1634 B.n505 VSUBS 0.007164f
C1635 B.n506 VSUBS 0.007164f
C1636 B.n507 VSUBS 0.007164f
C1637 B.n508 VSUBS 0.007164f
C1638 B.n509 VSUBS 0.007164f
C1639 B.n510 VSUBS 0.007164f
C1640 B.n511 VSUBS 0.007164f
C1641 B.n512 VSUBS 0.007164f
C1642 B.n513 VSUBS 0.007164f
C1643 B.n514 VSUBS 0.007164f
C1644 B.n515 VSUBS 0.007164f
C1645 B.n516 VSUBS 0.007164f
C1646 B.n517 VSUBS 0.007164f
C1647 B.n518 VSUBS 0.007164f
C1648 B.n519 VSUBS 0.007164f
C1649 B.n520 VSUBS 0.007164f
C1650 B.n521 VSUBS 0.007164f
C1651 B.n522 VSUBS 0.007164f
C1652 B.n523 VSUBS 0.007164f
C1653 B.n524 VSUBS 0.007164f
C1654 B.n525 VSUBS 0.007164f
C1655 B.n526 VSUBS 0.007164f
C1656 B.n527 VSUBS 0.007164f
C1657 B.n528 VSUBS 0.007164f
C1658 B.n529 VSUBS 0.007164f
C1659 B.n530 VSUBS 0.007164f
C1660 B.n531 VSUBS 0.007164f
C1661 B.n532 VSUBS 0.007164f
C1662 B.n533 VSUBS 0.007164f
C1663 B.n534 VSUBS 0.007164f
C1664 B.n535 VSUBS 0.007164f
C1665 B.n536 VSUBS 0.007164f
C1666 B.n537 VSUBS 0.007164f
C1667 B.n538 VSUBS 0.007164f
C1668 B.n539 VSUBS 0.007164f
C1669 B.n540 VSUBS 0.007164f
C1670 B.n541 VSUBS 0.007164f
C1671 B.n542 VSUBS 0.007164f
C1672 B.n543 VSUBS 0.007164f
C1673 B.n544 VSUBS 0.007164f
C1674 B.n545 VSUBS 0.007164f
C1675 B.n546 VSUBS 0.007164f
C1676 B.n547 VSUBS 0.007164f
C1677 B.n548 VSUBS 0.007164f
C1678 B.n549 VSUBS 0.007164f
C1679 B.n550 VSUBS 0.007164f
C1680 B.n551 VSUBS 0.007164f
C1681 B.n552 VSUBS 0.007164f
C1682 B.n553 VSUBS 0.007164f
C1683 B.n554 VSUBS 0.007164f
C1684 B.n555 VSUBS 0.007164f
C1685 B.n556 VSUBS 0.007164f
C1686 B.n557 VSUBS 0.007164f
C1687 B.n558 VSUBS 0.007164f
C1688 B.n559 VSUBS 0.007164f
C1689 B.n560 VSUBS 0.007164f
C1690 B.n561 VSUBS 0.007164f
C1691 B.n562 VSUBS 0.007164f
C1692 B.n563 VSUBS 0.007164f
C1693 B.n564 VSUBS 0.007164f
C1694 B.n565 VSUBS 0.007164f
C1695 B.n566 VSUBS 0.007164f
C1696 B.n567 VSUBS 0.007164f
C1697 B.n568 VSUBS 0.007164f
C1698 B.n569 VSUBS 0.007164f
C1699 B.n570 VSUBS 0.007164f
C1700 B.n571 VSUBS 0.007164f
C1701 B.n572 VSUBS 0.007164f
C1702 B.n573 VSUBS 0.007164f
C1703 B.n574 VSUBS 0.007164f
C1704 B.n575 VSUBS 0.007164f
C1705 B.n576 VSUBS 0.007164f
C1706 B.n577 VSUBS 0.007164f
C1707 B.n578 VSUBS 0.007164f
C1708 B.n579 VSUBS 0.007164f
C1709 B.n580 VSUBS 0.007164f
C1710 B.n581 VSUBS 0.007164f
C1711 B.n582 VSUBS 0.007164f
C1712 B.n583 VSUBS 0.007164f
C1713 B.n584 VSUBS 0.007164f
C1714 B.n585 VSUBS 0.007164f
C1715 B.n586 VSUBS 0.007164f
C1716 B.n587 VSUBS 0.007164f
C1717 B.n588 VSUBS 0.007164f
C1718 B.n589 VSUBS 0.007164f
C1719 B.n590 VSUBS 0.015764f
C1720 B.n591 VSUBS 0.015764f
C1721 B.n592 VSUBS 0.014786f
C1722 B.n593 VSUBS 0.007164f
C1723 B.n594 VSUBS 0.007164f
C1724 B.n595 VSUBS 0.007164f
C1725 B.n596 VSUBS 0.007164f
C1726 B.n597 VSUBS 0.007164f
C1727 B.n598 VSUBS 0.007164f
C1728 B.n599 VSUBS 0.007164f
C1729 B.n600 VSUBS 0.007164f
C1730 B.n601 VSUBS 0.007164f
C1731 B.n602 VSUBS 0.007164f
C1732 B.n603 VSUBS 0.007164f
C1733 B.n604 VSUBS 0.007164f
C1734 B.n605 VSUBS 0.007164f
C1735 B.n606 VSUBS 0.007164f
C1736 B.n607 VSUBS 0.007164f
C1737 B.n608 VSUBS 0.007164f
C1738 B.n609 VSUBS 0.007164f
C1739 B.n610 VSUBS 0.007164f
C1740 B.n611 VSUBS 0.007164f
C1741 B.n612 VSUBS 0.007164f
C1742 B.n613 VSUBS 0.007164f
C1743 B.n614 VSUBS 0.007164f
C1744 B.n615 VSUBS 0.007164f
C1745 B.n616 VSUBS 0.007164f
C1746 B.n617 VSUBS 0.007164f
C1747 B.n618 VSUBS 0.007164f
C1748 B.n619 VSUBS 0.007164f
C1749 B.n620 VSUBS 0.007164f
C1750 B.n621 VSUBS 0.007164f
C1751 B.n622 VSUBS 0.007164f
C1752 B.n623 VSUBS 0.007164f
C1753 B.n624 VSUBS 0.007164f
C1754 B.n625 VSUBS 0.007164f
C1755 B.n626 VSUBS 0.007164f
C1756 B.n627 VSUBS 0.007164f
C1757 B.n628 VSUBS 0.007164f
C1758 B.n629 VSUBS 0.007164f
C1759 B.n630 VSUBS 0.007164f
C1760 B.n631 VSUBS 0.007164f
C1761 B.n632 VSUBS 0.007164f
C1762 B.n633 VSUBS 0.007164f
C1763 B.n634 VSUBS 0.007164f
C1764 B.n635 VSUBS 0.007164f
C1765 B.n636 VSUBS 0.007164f
C1766 B.n637 VSUBS 0.007164f
C1767 B.n638 VSUBS 0.007164f
C1768 B.n639 VSUBS 0.007164f
C1769 B.n640 VSUBS 0.007164f
C1770 B.n641 VSUBS 0.007164f
C1771 B.n642 VSUBS 0.007164f
C1772 B.n643 VSUBS 0.007164f
C1773 B.n644 VSUBS 0.007164f
C1774 B.n645 VSUBS 0.007164f
C1775 B.n646 VSUBS 0.007164f
C1776 B.n647 VSUBS 0.007164f
C1777 B.n648 VSUBS 0.007164f
C1778 B.n649 VSUBS 0.007164f
C1779 B.n650 VSUBS 0.007164f
C1780 B.n651 VSUBS 0.007164f
C1781 B.n652 VSUBS 0.007164f
C1782 B.n653 VSUBS 0.007164f
C1783 B.n654 VSUBS 0.007164f
C1784 B.n655 VSUBS 0.007164f
C1785 B.n656 VSUBS 0.007164f
C1786 B.n657 VSUBS 0.007164f
C1787 B.n658 VSUBS 0.007164f
C1788 B.n659 VSUBS 0.007164f
C1789 B.n660 VSUBS 0.007164f
C1790 B.n661 VSUBS 0.007164f
C1791 B.n662 VSUBS 0.007164f
C1792 B.n663 VSUBS 0.007164f
C1793 B.n664 VSUBS 0.007164f
C1794 B.n665 VSUBS 0.007164f
C1795 B.n666 VSUBS 0.007164f
C1796 B.n667 VSUBS 0.007164f
C1797 B.n668 VSUBS 0.007164f
C1798 B.n669 VSUBS 0.007164f
C1799 B.n670 VSUBS 0.007164f
C1800 B.n671 VSUBS 0.007164f
C1801 B.n672 VSUBS 0.007164f
C1802 B.n673 VSUBS 0.007164f
C1803 B.n674 VSUBS 0.007164f
C1804 B.n675 VSUBS 0.007164f
C1805 B.n676 VSUBS 0.007164f
C1806 B.n677 VSUBS 0.007164f
C1807 B.n678 VSUBS 0.007164f
C1808 B.n679 VSUBS 0.007164f
C1809 B.n680 VSUBS 0.007164f
C1810 B.n681 VSUBS 0.007164f
C1811 B.n682 VSUBS 0.007164f
C1812 B.n683 VSUBS 0.007164f
C1813 B.n684 VSUBS 0.007164f
C1814 B.n685 VSUBS 0.007164f
C1815 B.n686 VSUBS 0.007164f
C1816 B.n687 VSUBS 0.007164f
C1817 B.n688 VSUBS 0.007164f
C1818 B.n689 VSUBS 0.007164f
C1819 B.n690 VSUBS 0.007164f
C1820 B.n691 VSUBS 0.007164f
C1821 B.n692 VSUBS 0.007164f
C1822 B.n693 VSUBS 0.007164f
C1823 B.n694 VSUBS 0.007164f
C1824 B.n695 VSUBS 0.007164f
C1825 B.n696 VSUBS 0.007164f
C1826 B.n697 VSUBS 0.007164f
C1827 B.n698 VSUBS 0.007164f
C1828 B.n699 VSUBS 0.007164f
C1829 B.n700 VSUBS 0.007164f
C1830 B.n701 VSUBS 0.007164f
C1831 B.n702 VSUBS 0.007164f
C1832 B.n703 VSUBS 0.007164f
C1833 B.n704 VSUBS 0.007164f
C1834 B.n705 VSUBS 0.007164f
C1835 B.n706 VSUBS 0.007164f
C1836 B.n707 VSUBS 0.007164f
C1837 B.n708 VSUBS 0.007164f
C1838 B.n709 VSUBS 0.007164f
C1839 B.n710 VSUBS 0.007164f
C1840 B.n711 VSUBS 0.007164f
C1841 B.n712 VSUBS 0.007164f
C1842 B.n713 VSUBS 0.007164f
C1843 B.n714 VSUBS 0.007164f
C1844 B.n715 VSUBS 0.007164f
C1845 B.n716 VSUBS 0.007164f
C1846 B.n717 VSUBS 0.007164f
C1847 B.n718 VSUBS 0.007164f
C1848 B.n719 VSUBS 0.007164f
C1849 B.n720 VSUBS 0.007164f
C1850 B.n721 VSUBS 0.007164f
C1851 B.n722 VSUBS 0.007164f
C1852 B.n723 VSUBS 0.007164f
C1853 B.n724 VSUBS 0.007164f
C1854 B.n725 VSUBS 0.007164f
C1855 B.n726 VSUBS 0.007164f
C1856 B.n727 VSUBS 0.007164f
C1857 B.n728 VSUBS 0.007164f
C1858 B.n729 VSUBS 0.007164f
C1859 B.n730 VSUBS 0.007164f
C1860 B.n731 VSUBS 0.007164f
C1861 B.n732 VSUBS 0.007164f
C1862 B.n733 VSUBS 0.007164f
C1863 B.n734 VSUBS 0.007164f
C1864 B.n735 VSUBS 0.007164f
C1865 B.n736 VSUBS 0.007164f
C1866 B.n737 VSUBS 0.007164f
C1867 B.n738 VSUBS 0.007164f
C1868 B.n739 VSUBS 0.007164f
C1869 B.n740 VSUBS 0.007164f
C1870 B.n741 VSUBS 0.007164f
C1871 B.n742 VSUBS 0.007164f
C1872 B.n743 VSUBS 0.007164f
C1873 B.n744 VSUBS 0.007164f
C1874 B.n745 VSUBS 0.007164f
C1875 B.n746 VSUBS 0.007164f
C1876 B.n747 VSUBS 0.007164f
C1877 B.n748 VSUBS 0.007164f
C1878 B.n749 VSUBS 0.007164f
C1879 B.n750 VSUBS 0.007164f
C1880 B.n751 VSUBS 0.007164f
C1881 B.n752 VSUBS 0.007164f
C1882 B.n753 VSUBS 0.007164f
C1883 B.n754 VSUBS 0.007164f
C1884 B.n755 VSUBS 0.007164f
C1885 B.n756 VSUBS 0.007164f
C1886 B.n757 VSUBS 0.007164f
C1887 B.n758 VSUBS 0.007164f
C1888 B.n759 VSUBS 0.007164f
C1889 B.n760 VSUBS 0.007164f
C1890 B.n761 VSUBS 0.007164f
C1891 B.n762 VSUBS 0.007164f
C1892 B.n763 VSUBS 0.007164f
C1893 B.n764 VSUBS 0.007164f
C1894 B.n765 VSUBS 0.007164f
C1895 B.n766 VSUBS 0.007164f
C1896 B.n767 VSUBS 0.007164f
C1897 B.n768 VSUBS 0.007164f
C1898 B.n769 VSUBS 0.007164f
C1899 B.n770 VSUBS 0.007164f
C1900 B.n771 VSUBS 0.007164f
C1901 B.n772 VSUBS 0.007164f
C1902 B.n773 VSUBS 0.007164f
C1903 B.n774 VSUBS 0.007164f
C1904 B.n775 VSUBS 0.007164f
C1905 B.n776 VSUBS 0.007164f
C1906 B.n777 VSUBS 0.007164f
C1907 B.n778 VSUBS 0.007164f
C1908 B.n779 VSUBS 0.007164f
C1909 B.n780 VSUBS 0.007164f
C1910 B.n781 VSUBS 0.007164f
C1911 B.n782 VSUBS 0.007164f
C1912 B.n783 VSUBS 0.007164f
C1913 B.n784 VSUBS 0.007164f
C1914 B.n785 VSUBS 0.007164f
C1915 B.n786 VSUBS 0.007164f
C1916 B.n787 VSUBS 0.007164f
C1917 B.n788 VSUBS 0.007164f
C1918 B.n789 VSUBS 0.007164f
C1919 B.n790 VSUBS 0.007164f
C1920 B.n791 VSUBS 0.007164f
C1921 B.n792 VSUBS 0.007164f
C1922 B.n793 VSUBS 0.007164f
C1923 B.n794 VSUBS 0.007164f
C1924 B.n795 VSUBS 0.007164f
C1925 B.n796 VSUBS 0.015764f
C1926 B.n797 VSUBS 0.014786f
C1927 B.n798 VSUBS 0.015764f
C1928 B.n799 VSUBS 0.007164f
C1929 B.n800 VSUBS 0.007164f
C1930 B.n801 VSUBS 0.007164f
C1931 B.n802 VSUBS 0.007164f
C1932 B.n803 VSUBS 0.007164f
C1933 B.n804 VSUBS 0.007164f
C1934 B.n805 VSUBS 0.007164f
C1935 B.n806 VSUBS 0.007164f
C1936 B.n807 VSUBS 0.007164f
C1937 B.n808 VSUBS 0.007164f
C1938 B.n809 VSUBS 0.007164f
C1939 B.n810 VSUBS 0.007164f
C1940 B.n811 VSUBS 0.007164f
C1941 B.n812 VSUBS 0.007164f
C1942 B.n813 VSUBS 0.007164f
C1943 B.n814 VSUBS 0.007164f
C1944 B.n815 VSUBS 0.007164f
C1945 B.n816 VSUBS 0.007164f
C1946 B.n817 VSUBS 0.007164f
C1947 B.n818 VSUBS 0.007164f
C1948 B.n819 VSUBS 0.007164f
C1949 B.n820 VSUBS 0.007164f
C1950 B.n821 VSUBS 0.007164f
C1951 B.n822 VSUBS 0.007164f
C1952 B.n823 VSUBS 0.007164f
C1953 B.n824 VSUBS 0.007164f
C1954 B.n825 VSUBS 0.007164f
C1955 B.n826 VSUBS 0.007164f
C1956 B.n827 VSUBS 0.007164f
C1957 B.n828 VSUBS 0.007164f
C1958 B.n829 VSUBS 0.007164f
C1959 B.n830 VSUBS 0.007164f
C1960 B.n831 VSUBS 0.007164f
C1961 B.n832 VSUBS 0.007164f
C1962 B.n833 VSUBS 0.007164f
C1963 B.n834 VSUBS 0.007164f
C1964 B.n835 VSUBS 0.007164f
C1965 B.n836 VSUBS 0.007164f
C1966 B.n837 VSUBS 0.007164f
C1967 B.n838 VSUBS 0.007164f
C1968 B.n839 VSUBS 0.007164f
C1969 B.n840 VSUBS 0.007164f
C1970 B.n841 VSUBS 0.007164f
C1971 B.n842 VSUBS 0.007164f
C1972 B.n843 VSUBS 0.007164f
C1973 B.n844 VSUBS 0.007164f
C1974 B.n845 VSUBS 0.007164f
C1975 B.n846 VSUBS 0.007164f
C1976 B.n847 VSUBS 0.007164f
C1977 B.n848 VSUBS 0.007164f
C1978 B.n849 VSUBS 0.007164f
C1979 B.n850 VSUBS 0.007164f
C1980 B.n851 VSUBS 0.007164f
C1981 B.n852 VSUBS 0.007164f
C1982 B.n853 VSUBS 0.007164f
C1983 B.n854 VSUBS 0.007164f
C1984 B.n855 VSUBS 0.007164f
C1985 B.n856 VSUBS 0.007164f
C1986 B.n857 VSUBS 0.007164f
C1987 B.n858 VSUBS 0.007164f
C1988 B.n859 VSUBS 0.007164f
C1989 B.n860 VSUBS 0.007164f
C1990 B.n861 VSUBS 0.007164f
C1991 B.n862 VSUBS 0.007164f
C1992 B.n863 VSUBS 0.007164f
C1993 B.n864 VSUBS 0.007164f
C1994 B.n865 VSUBS 0.007164f
C1995 B.n866 VSUBS 0.007164f
C1996 B.n867 VSUBS 0.007164f
C1997 B.n868 VSUBS 0.007164f
C1998 B.n869 VSUBS 0.007164f
C1999 B.n870 VSUBS 0.007164f
C2000 B.n871 VSUBS 0.007164f
C2001 B.n872 VSUBS 0.007164f
C2002 B.n873 VSUBS 0.007164f
C2003 B.n874 VSUBS 0.007164f
C2004 B.n875 VSUBS 0.007164f
C2005 B.n876 VSUBS 0.007164f
C2006 B.n877 VSUBS 0.007164f
C2007 B.n878 VSUBS 0.007164f
C2008 B.n879 VSUBS 0.007164f
C2009 B.n880 VSUBS 0.007164f
C2010 B.n881 VSUBS 0.007164f
C2011 B.n882 VSUBS 0.007164f
C2012 B.n883 VSUBS 0.007164f
C2013 B.n884 VSUBS 0.007164f
C2014 B.n885 VSUBS 0.007164f
C2015 B.n886 VSUBS 0.007164f
C2016 B.n887 VSUBS 0.007164f
C2017 B.n888 VSUBS 0.007164f
C2018 B.n889 VSUBS 0.007164f
C2019 B.n890 VSUBS 0.007164f
C2020 B.n891 VSUBS 0.007164f
C2021 B.n892 VSUBS 0.004951f
C2022 B.n893 VSUBS 0.016597f
C2023 B.n894 VSUBS 0.005794f
C2024 B.n895 VSUBS 0.007164f
C2025 B.n896 VSUBS 0.007164f
C2026 B.n897 VSUBS 0.007164f
C2027 B.n898 VSUBS 0.007164f
C2028 B.n899 VSUBS 0.007164f
C2029 B.n900 VSUBS 0.007164f
C2030 B.n901 VSUBS 0.007164f
C2031 B.n902 VSUBS 0.007164f
C2032 B.n903 VSUBS 0.007164f
C2033 B.n904 VSUBS 0.007164f
C2034 B.n905 VSUBS 0.007164f
C2035 B.n906 VSUBS 0.005794f
C2036 B.n907 VSUBS 0.007164f
C2037 B.n908 VSUBS 0.007164f
C2038 B.n909 VSUBS 0.004951f
C2039 B.n910 VSUBS 0.007164f
C2040 B.n911 VSUBS 0.007164f
C2041 B.n912 VSUBS 0.007164f
C2042 B.n913 VSUBS 0.007164f
C2043 B.n914 VSUBS 0.007164f
C2044 B.n915 VSUBS 0.007164f
C2045 B.n916 VSUBS 0.007164f
C2046 B.n917 VSUBS 0.007164f
C2047 B.n918 VSUBS 0.007164f
C2048 B.n919 VSUBS 0.007164f
C2049 B.n920 VSUBS 0.007164f
C2050 B.n921 VSUBS 0.007164f
C2051 B.n922 VSUBS 0.007164f
C2052 B.n923 VSUBS 0.007164f
C2053 B.n924 VSUBS 0.007164f
C2054 B.n925 VSUBS 0.007164f
C2055 B.n926 VSUBS 0.007164f
C2056 B.n927 VSUBS 0.007164f
C2057 B.n928 VSUBS 0.007164f
C2058 B.n929 VSUBS 0.007164f
C2059 B.n930 VSUBS 0.007164f
C2060 B.n931 VSUBS 0.007164f
C2061 B.n932 VSUBS 0.007164f
C2062 B.n933 VSUBS 0.007164f
C2063 B.n934 VSUBS 0.007164f
C2064 B.n935 VSUBS 0.007164f
C2065 B.n936 VSUBS 0.007164f
C2066 B.n937 VSUBS 0.007164f
C2067 B.n938 VSUBS 0.007164f
C2068 B.n939 VSUBS 0.007164f
C2069 B.n940 VSUBS 0.007164f
C2070 B.n941 VSUBS 0.007164f
C2071 B.n942 VSUBS 0.007164f
C2072 B.n943 VSUBS 0.007164f
C2073 B.n944 VSUBS 0.007164f
C2074 B.n945 VSUBS 0.007164f
C2075 B.n946 VSUBS 0.007164f
C2076 B.n947 VSUBS 0.007164f
C2077 B.n948 VSUBS 0.007164f
C2078 B.n949 VSUBS 0.007164f
C2079 B.n950 VSUBS 0.007164f
C2080 B.n951 VSUBS 0.007164f
C2081 B.n952 VSUBS 0.007164f
C2082 B.n953 VSUBS 0.007164f
C2083 B.n954 VSUBS 0.007164f
C2084 B.n955 VSUBS 0.007164f
C2085 B.n956 VSUBS 0.007164f
C2086 B.n957 VSUBS 0.007164f
C2087 B.n958 VSUBS 0.007164f
C2088 B.n959 VSUBS 0.007164f
C2089 B.n960 VSUBS 0.007164f
C2090 B.n961 VSUBS 0.007164f
C2091 B.n962 VSUBS 0.007164f
C2092 B.n963 VSUBS 0.007164f
C2093 B.n964 VSUBS 0.007164f
C2094 B.n965 VSUBS 0.007164f
C2095 B.n966 VSUBS 0.007164f
C2096 B.n967 VSUBS 0.007164f
C2097 B.n968 VSUBS 0.007164f
C2098 B.n969 VSUBS 0.007164f
C2099 B.n970 VSUBS 0.007164f
C2100 B.n971 VSUBS 0.007164f
C2101 B.n972 VSUBS 0.007164f
C2102 B.n973 VSUBS 0.007164f
C2103 B.n974 VSUBS 0.007164f
C2104 B.n975 VSUBS 0.007164f
C2105 B.n976 VSUBS 0.007164f
C2106 B.n977 VSUBS 0.007164f
C2107 B.n978 VSUBS 0.007164f
C2108 B.n979 VSUBS 0.007164f
C2109 B.n980 VSUBS 0.007164f
C2110 B.n981 VSUBS 0.007164f
C2111 B.n982 VSUBS 0.007164f
C2112 B.n983 VSUBS 0.007164f
C2113 B.n984 VSUBS 0.007164f
C2114 B.n985 VSUBS 0.007164f
C2115 B.n986 VSUBS 0.007164f
C2116 B.n987 VSUBS 0.007164f
C2117 B.n988 VSUBS 0.007164f
C2118 B.n989 VSUBS 0.007164f
C2119 B.n990 VSUBS 0.007164f
C2120 B.n991 VSUBS 0.007164f
C2121 B.n992 VSUBS 0.007164f
C2122 B.n993 VSUBS 0.007164f
C2123 B.n994 VSUBS 0.007164f
C2124 B.n995 VSUBS 0.007164f
C2125 B.n996 VSUBS 0.007164f
C2126 B.n997 VSUBS 0.007164f
C2127 B.n998 VSUBS 0.007164f
C2128 B.n999 VSUBS 0.007164f
C2129 B.n1000 VSUBS 0.007164f
C2130 B.n1001 VSUBS 0.007164f
C2131 B.n1002 VSUBS 0.007164f
C2132 B.n1003 VSUBS 0.015764f
C2133 B.n1004 VSUBS 0.014786f
C2134 B.n1005 VSUBS 0.014786f
C2135 B.n1006 VSUBS 0.007164f
C2136 B.n1007 VSUBS 0.007164f
C2137 B.n1008 VSUBS 0.007164f
C2138 B.n1009 VSUBS 0.007164f
C2139 B.n1010 VSUBS 0.007164f
C2140 B.n1011 VSUBS 0.007164f
C2141 B.n1012 VSUBS 0.007164f
C2142 B.n1013 VSUBS 0.007164f
C2143 B.n1014 VSUBS 0.007164f
C2144 B.n1015 VSUBS 0.007164f
C2145 B.n1016 VSUBS 0.007164f
C2146 B.n1017 VSUBS 0.007164f
C2147 B.n1018 VSUBS 0.007164f
C2148 B.n1019 VSUBS 0.007164f
C2149 B.n1020 VSUBS 0.007164f
C2150 B.n1021 VSUBS 0.007164f
C2151 B.n1022 VSUBS 0.007164f
C2152 B.n1023 VSUBS 0.007164f
C2153 B.n1024 VSUBS 0.007164f
C2154 B.n1025 VSUBS 0.007164f
C2155 B.n1026 VSUBS 0.007164f
C2156 B.n1027 VSUBS 0.007164f
C2157 B.n1028 VSUBS 0.007164f
C2158 B.n1029 VSUBS 0.007164f
C2159 B.n1030 VSUBS 0.007164f
C2160 B.n1031 VSUBS 0.007164f
C2161 B.n1032 VSUBS 0.007164f
C2162 B.n1033 VSUBS 0.007164f
C2163 B.n1034 VSUBS 0.007164f
C2164 B.n1035 VSUBS 0.007164f
C2165 B.n1036 VSUBS 0.007164f
C2166 B.n1037 VSUBS 0.007164f
C2167 B.n1038 VSUBS 0.007164f
C2168 B.n1039 VSUBS 0.007164f
C2169 B.n1040 VSUBS 0.007164f
C2170 B.n1041 VSUBS 0.007164f
C2171 B.n1042 VSUBS 0.007164f
C2172 B.n1043 VSUBS 0.007164f
C2173 B.n1044 VSUBS 0.007164f
C2174 B.n1045 VSUBS 0.007164f
C2175 B.n1046 VSUBS 0.007164f
C2176 B.n1047 VSUBS 0.007164f
C2177 B.n1048 VSUBS 0.007164f
C2178 B.n1049 VSUBS 0.007164f
C2179 B.n1050 VSUBS 0.007164f
C2180 B.n1051 VSUBS 0.007164f
C2181 B.n1052 VSUBS 0.007164f
C2182 B.n1053 VSUBS 0.007164f
C2183 B.n1054 VSUBS 0.007164f
C2184 B.n1055 VSUBS 0.007164f
C2185 B.n1056 VSUBS 0.007164f
C2186 B.n1057 VSUBS 0.007164f
C2187 B.n1058 VSUBS 0.007164f
C2188 B.n1059 VSUBS 0.007164f
C2189 B.n1060 VSUBS 0.007164f
C2190 B.n1061 VSUBS 0.007164f
C2191 B.n1062 VSUBS 0.007164f
C2192 B.n1063 VSUBS 0.007164f
C2193 B.n1064 VSUBS 0.007164f
C2194 B.n1065 VSUBS 0.007164f
C2195 B.n1066 VSUBS 0.007164f
C2196 B.n1067 VSUBS 0.007164f
C2197 B.n1068 VSUBS 0.007164f
C2198 B.n1069 VSUBS 0.007164f
C2199 B.n1070 VSUBS 0.007164f
C2200 B.n1071 VSUBS 0.007164f
C2201 B.n1072 VSUBS 0.007164f
C2202 B.n1073 VSUBS 0.007164f
C2203 B.n1074 VSUBS 0.007164f
C2204 B.n1075 VSUBS 0.007164f
C2205 B.n1076 VSUBS 0.007164f
C2206 B.n1077 VSUBS 0.007164f
C2207 B.n1078 VSUBS 0.007164f
C2208 B.n1079 VSUBS 0.007164f
C2209 B.n1080 VSUBS 0.007164f
C2210 B.n1081 VSUBS 0.007164f
C2211 B.n1082 VSUBS 0.007164f
C2212 B.n1083 VSUBS 0.007164f
C2213 B.n1084 VSUBS 0.007164f
C2214 B.n1085 VSUBS 0.007164f
C2215 B.n1086 VSUBS 0.007164f
C2216 B.n1087 VSUBS 0.007164f
C2217 B.n1088 VSUBS 0.007164f
C2218 B.n1089 VSUBS 0.007164f
C2219 B.n1090 VSUBS 0.007164f
C2220 B.n1091 VSUBS 0.007164f
C2221 B.n1092 VSUBS 0.007164f
C2222 B.n1093 VSUBS 0.007164f
C2223 B.n1094 VSUBS 0.007164f
C2224 B.n1095 VSUBS 0.007164f
C2225 B.n1096 VSUBS 0.007164f
C2226 B.n1097 VSUBS 0.007164f
C2227 B.n1098 VSUBS 0.007164f
C2228 B.n1099 VSUBS 0.007164f
C2229 B.n1100 VSUBS 0.007164f
C2230 B.n1101 VSUBS 0.007164f
C2231 B.n1102 VSUBS 0.007164f
C2232 B.n1103 VSUBS 0.007164f
C2233 B.n1104 VSUBS 0.007164f
C2234 B.n1105 VSUBS 0.007164f
C2235 B.n1106 VSUBS 0.007164f
C2236 B.n1107 VSUBS 0.016221f
.ends

