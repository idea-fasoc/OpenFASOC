* NGSPICE file created from diff_pair_sample_1646.ext - technology: sky130A

.subckt diff_pair_sample_1646 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=2.9055 ps=15.68 w=7.45 l=0.6
X1 B.t11 B.t9 B.t10 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=0 ps=0 w=7.45 l=0.6
X2 VDD1.t1 VP.t0 VTAIL.t0 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=2.9055 ps=15.68 w=7.45 l=0.6
X3 B.t8 B.t6 B.t7 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=0 ps=0 w=7.45 l=0.6
X4 B.t5 B.t3 B.t4 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=0 ps=0 w=7.45 l=0.6
X5 B.t2 B.t0 B.t1 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=0 ps=0 w=7.45 l=0.6
X6 VDD2.t0 VN.t1 VTAIL.t3 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=2.9055 ps=15.68 w=7.45 l=0.6
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1342_n2462# sky130_fd_pr__pfet_01v8 ad=2.9055 pd=15.68 as=2.9055 ps=15.68 w=7.45 l=0.6
R0 VN VN.t1 562.716
R1 VN VN.t0 526.466
R2 VTAIL.n154 VTAIL.n120 756.745
R3 VTAIL.n34 VTAIL.n0 756.745
R4 VTAIL.n114 VTAIL.n80 756.745
R5 VTAIL.n74 VTAIL.n40 756.745
R6 VTAIL.n132 VTAIL.n131 585
R7 VTAIL.n137 VTAIL.n136 585
R8 VTAIL.n139 VTAIL.n138 585
R9 VTAIL.n128 VTAIL.n127 585
R10 VTAIL.n145 VTAIL.n144 585
R11 VTAIL.n147 VTAIL.n146 585
R12 VTAIL.n124 VTAIL.n123 585
R13 VTAIL.n153 VTAIL.n152 585
R14 VTAIL.n155 VTAIL.n154 585
R15 VTAIL.n12 VTAIL.n11 585
R16 VTAIL.n17 VTAIL.n16 585
R17 VTAIL.n19 VTAIL.n18 585
R18 VTAIL.n8 VTAIL.n7 585
R19 VTAIL.n25 VTAIL.n24 585
R20 VTAIL.n27 VTAIL.n26 585
R21 VTAIL.n4 VTAIL.n3 585
R22 VTAIL.n33 VTAIL.n32 585
R23 VTAIL.n35 VTAIL.n34 585
R24 VTAIL.n115 VTAIL.n114 585
R25 VTAIL.n113 VTAIL.n112 585
R26 VTAIL.n84 VTAIL.n83 585
R27 VTAIL.n107 VTAIL.n106 585
R28 VTAIL.n105 VTAIL.n104 585
R29 VTAIL.n88 VTAIL.n87 585
R30 VTAIL.n99 VTAIL.n98 585
R31 VTAIL.n97 VTAIL.n96 585
R32 VTAIL.n92 VTAIL.n91 585
R33 VTAIL.n75 VTAIL.n74 585
R34 VTAIL.n73 VTAIL.n72 585
R35 VTAIL.n44 VTAIL.n43 585
R36 VTAIL.n67 VTAIL.n66 585
R37 VTAIL.n65 VTAIL.n64 585
R38 VTAIL.n48 VTAIL.n47 585
R39 VTAIL.n59 VTAIL.n58 585
R40 VTAIL.n57 VTAIL.n56 585
R41 VTAIL.n52 VTAIL.n51 585
R42 VTAIL.n133 VTAIL.t2 327.483
R43 VTAIL.n13 VTAIL.t0 327.483
R44 VTAIL.n93 VTAIL.t1 327.483
R45 VTAIL.n53 VTAIL.t3 327.483
R46 VTAIL.n137 VTAIL.n131 171.744
R47 VTAIL.n138 VTAIL.n137 171.744
R48 VTAIL.n138 VTAIL.n127 171.744
R49 VTAIL.n145 VTAIL.n127 171.744
R50 VTAIL.n146 VTAIL.n145 171.744
R51 VTAIL.n146 VTAIL.n123 171.744
R52 VTAIL.n153 VTAIL.n123 171.744
R53 VTAIL.n154 VTAIL.n153 171.744
R54 VTAIL.n17 VTAIL.n11 171.744
R55 VTAIL.n18 VTAIL.n17 171.744
R56 VTAIL.n18 VTAIL.n7 171.744
R57 VTAIL.n25 VTAIL.n7 171.744
R58 VTAIL.n26 VTAIL.n25 171.744
R59 VTAIL.n26 VTAIL.n3 171.744
R60 VTAIL.n33 VTAIL.n3 171.744
R61 VTAIL.n34 VTAIL.n33 171.744
R62 VTAIL.n114 VTAIL.n113 171.744
R63 VTAIL.n113 VTAIL.n83 171.744
R64 VTAIL.n106 VTAIL.n83 171.744
R65 VTAIL.n106 VTAIL.n105 171.744
R66 VTAIL.n105 VTAIL.n87 171.744
R67 VTAIL.n98 VTAIL.n87 171.744
R68 VTAIL.n98 VTAIL.n97 171.744
R69 VTAIL.n97 VTAIL.n91 171.744
R70 VTAIL.n74 VTAIL.n73 171.744
R71 VTAIL.n73 VTAIL.n43 171.744
R72 VTAIL.n66 VTAIL.n43 171.744
R73 VTAIL.n66 VTAIL.n65 171.744
R74 VTAIL.n65 VTAIL.n47 171.744
R75 VTAIL.n58 VTAIL.n47 171.744
R76 VTAIL.n58 VTAIL.n57 171.744
R77 VTAIL.n57 VTAIL.n51 171.744
R78 VTAIL.t2 VTAIL.n131 85.8723
R79 VTAIL.t0 VTAIL.n11 85.8723
R80 VTAIL.t1 VTAIL.n91 85.8723
R81 VTAIL.t3 VTAIL.n51 85.8723
R82 VTAIL.n159 VTAIL.n158 32.3793
R83 VTAIL.n39 VTAIL.n38 32.3793
R84 VTAIL.n119 VTAIL.n118 32.3793
R85 VTAIL.n79 VTAIL.n78 32.3793
R86 VTAIL.n79 VTAIL.n39 20.41
R87 VTAIL.n159 VTAIL.n119 19.6083
R88 VTAIL.n133 VTAIL.n132 16.3891
R89 VTAIL.n13 VTAIL.n12 16.3891
R90 VTAIL.n93 VTAIL.n92 16.3891
R91 VTAIL.n53 VTAIL.n52 16.3891
R92 VTAIL.n136 VTAIL.n135 12.8005
R93 VTAIL.n16 VTAIL.n15 12.8005
R94 VTAIL.n96 VTAIL.n95 12.8005
R95 VTAIL.n56 VTAIL.n55 12.8005
R96 VTAIL.n139 VTAIL.n130 12.0247
R97 VTAIL.n19 VTAIL.n10 12.0247
R98 VTAIL.n99 VTAIL.n90 12.0247
R99 VTAIL.n59 VTAIL.n50 12.0247
R100 VTAIL.n140 VTAIL.n128 11.249
R101 VTAIL.n20 VTAIL.n8 11.249
R102 VTAIL.n100 VTAIL.n88 11.249
R103 VTAIL.n60 VTAIL.n48 11.249
R104 VTAIL.n144 VTAIL.n143 10.4732
R105 VTAIL.n24 VTAIL.n23 10.4732
R106 VTAIL.n104 VTAIL.n103 10.4732
R107 VTAIL.n64 VTAIL.n63 10.4732
R108 VTAIL.n147 VTAIL.n126 9.69747
R109 VTAIL.n27 VTAIL.n6 9.69747
R110 VTAIL.n107 VTAIL.n86 9.69747
R111 VTAIL.n67 VTAIL.n46 9.69747
R112 VTAIL.n158 VTAIL.n157 9.45567
R113 VTAIL.n38 VTAIL.n37 9.45567
R114 VTAIL.n118 VTAIL.n117 9.45567
R115 VTAIL.n78 VTAIL.n77 9.45567
R116 VTAIL.n157 VTAIL.n156 9.3005
R117 VTAIL.n151 VTAIL.n150 9.3005
R118 VTAIL.n149 VTAIL.n148 9.3005
R119 VTAIL.n126 VTAIL.n125 9.3005
R120 VTAIL.n143 VTAIL.n142 9.3005
R121 VTAIL.n141 VTAIL.n140 9.3005
R122 VTAIL.n130 VTAIL.n129 9.3005
R123 VTAIL.n135 VTAIL.n134 9.3005
R124 VTAIL.n122 VTAIL.n121 9.3005
R125 VTAIL.n37 VTAIL.n36 9.3005
R126 VTAIL.n31 VTAIL.n30 9.3005
R127 VTAIL.n29 VTAIL.n28 9.3005
R128 VTAIL.n6 VTAIL.n5 9.3005
R129 VTAIL.n23 VTAIL.n22 9.3005
R130 VTAIL.n21 VTAIL.n20 9.3005
R131 VTAIL.n10 VTAIL.n9 9.3005
R132 VTAIL.n15 VTAIL.n14 9.3005
R133 VTAIL.n2 VTAIL.n1 9.3005
R134 VTAIL.n117 VTAIL.n116 9.3005
R135 VTAIL.n82 VTAIL.n81 9.3005
R136 VTAIL.n111 VTAIL.n110 9.3005
R137 VTAIL.n109 VTAIL.n108 9.3005
R138 VTAIL.n86 VTAIL.n85 9.3005
R139 VTAIL.n103 VTAIL.n102 9.3005
R140 VTAIL.n101 VTAIL.n100 9.3005
R141 VTAIL.n90 VTAIL.n89 9.3005
R142 VTAIL.n95 VTAIL.n94 9.3005
R143 VTAIL.n77 VTAIL.n76 9.3005
R144 VTAIL.n42 VTAIL.n41 9.3005
R145 VTAIL.n71 VTAIL.n70 9.3005
R146 VTAIL.n69 VTAIL.n68 9.3005
R147 VTAIL.n46 VTAIL.n45 9.3005
R148 VTAIL.n63 VTAIL.n62 9.3005
R149 VTAIL.n61 VTAIL.n60 9.3005
R150 VTAIL.n50 VTAIL.n49 9.3005
R151 VTAIL.n55 VTAIL.n54 9.3005
R152 VTAIL.n148 VTAIL.n124 8.92171
R153 VTAIL.n28 VTAIL.n4 8.92171
R154 VTAIL.n108 VTAIL.n84 8.92171
R155 VTAIL.n68 VTAIL.n44 8.92171
R156 VTAIL.n152 VTAIL.n151 8.14595
R157 VTAIL.n32 VTAIL.n31 8.14595
R158 VTAIL.n112 VTAIL.n111 8.14595
R159 VTAIL.n72 VTAIL.n71 8.14595
R160 VTAIL.n155 VTAIL.n122 7.3702
R161 VTAIL.n158 VTAIL.n120 7.3702
R162 VTAIL.n35 VTAIL.n2 7.3702
R163 VTAIL.n38 VTAIL.n0 7.3702
R164 VTAIL.n118 VTAIL.n80 7.3702
R165 VTAIL.n115 VTAIL.n82 7.3702
R166 VTAIL.n78 VTAIL.n40 7.3702
R167 VTAIL.n75 VTAIL.n42 7.3702
R168 VTAIL.n156 VTAIL.n155 6.59444
R169 VTAIL.n156 VTAIL.n120 6.59444
R170 VTAIL.n36 VTAIL.n35 6.59444
R171 VTAIL.n36 VTAIL.n0 6.59444
R172 VTAIL.n116 VTAIL.n80 6.59444
R173 VTAIL.n116 VTAIL.n115 6.59444
R174 VTAIL.n76 VTAIL.n40 6.59444
R175 VTAIL.n76 VTAIL.n75 6.59444
R176 VTAIL.n152 VTAIL.n122 5.81868
R177 VTAIL.n32 VTAIL.n2 5.81868
R178 VTAIL.n112 VTAIL.n82 5.81868
R179 VTAIL.n72 VTAIL.n42 5.81868
R180 VTAIL.n151 VTAIL.n124 5.04292
R181 VTAIL.n31 VTAIL.n4 5.04292
R182 VTAIL.n111 VTAIL.n84 5.04292
R183 VTAIL.n71 VTAIL.n44 5.04292
R184 VTAIL.n148 VTAIL.n147 4.26717
R185 VTAIL.n28 VTAIL.n27 4.26717
R186 VTAIL.n108 VTAIL.n107 4.26717
R187 VTAIL.n68 VTAIL.n67 4.26717
R188 VTAIL.n134 VTAIL.n133 3.71019
R189 VTAIL.n14 VTAIL.n13 3.71019
R190 VTAIL.n94 VTAIL.n93 3.71019
R191 VTAIL.n54 VTAIL.n53 3.71019
R192 VTAIL.n144 VTAIL.n126 3.49141
R193 VTAIL.n24 VTAIL.n6 3.49141
R194 VTAIL.n104 VTAIL.n86 3.49141
R195 VTAIL.n64 VTAIL.n46 3.49141
R196 VTAIL.n143 VTAIL.n128 2.71565
R197 VTAIL.n23 VTAIL.n8 2.71565
R198 VTAIL.n103 VTAIL.n88 2.71565
R199 VTAIL.n63 VTAIL.n48 2.71565
R200 VTAIL.n140 VTAIL.n139 1.93989
R201 VTAIL.n20 VTAIL.n19 1.93989
R202 VTAIL.n100 VTAIL.n99 1.93989
R203 VTAIL.n60 VTAIL.n59 1.93989
R204 VTAIL.n136 VTAIL.n130 1.16414
R205 VTAIL.n16 VTAIL.n10 1.16414
R206 VTAIL.n96 VTAIL.n90 1.16414
R207 VTAIL.n56 VTAIL.n50 1.16414
R208 VTAIL.n119 VTAIL.n79 0.87119
R209 VTAIL VTAIL.n39 0.728948
R210 VTAIL.n135 VTAIL.n132 0.388379
R211 VTAIL.n15 VTAIL.n12 0.388379
R212 VTAIL.n95 VTAIL.n92 0.388379
R213 VTAIL.n55 VTAIL.n52 0.388379
R214 VTAIL.n134 VTAIL.n129 0.155672
R215 VTAIL.n141 VTAIL.n129 0.155672
R216 VTAIL.n142 VTAIL.n141 0.155672
R217 VTAIL.n142 VTAIL.n125 0.155672
R218 VTAIL.n149 VTAIL.n125 0.155672
R219 VTAIL.n150 VTAIL.n149 0.155672
R220 VTAIL.n150 VTAIL.n121 0.155672
R221 VTAIL.n157 VTAIL.n121 0.155672
R222 VTAIL.n14 VTAIL.n9 0.155672
R223 VTAIL.n21 VTAIL.n9 0.155672
R224 VTAIL.n22 VTAIL.n21 0.155672
R225 VTAIL.n22 VTAIL.n5 0.155672
R226 VTAIL.n29 VTAIL.n5 0.155672
R227 VTAIL.n30 VTAIL.n29 0.155672
R228 VTAIL.n30 VTAIL.n1 0.155672
R229 VTAIL.n37 VTAIL.n1 0.155672
R230 VTAIL.n117 VTAIL.n81 0.155672
R231 VTAIL.n110 VTAIL.n81 0.155672
R232 VTAIL.n110 VTAIL.n109 0.155672
R233 VTAIL.n109 VTAIL.n85 0.155672
R234 VTAIL.n102 VTAIL.n85 0.155672
R235 VTAIL.n102 VTAIL.n101 0.155672
R236 VTAIL.n101 VTAIL.n89 0.155672
R237 VTAIL.n94 VTAIL.n89 0.155672
R238 VTAIL.n77 VTAIL.n41 0.155672
R239 VTAIL.n70 VTAIL.n41 0.155672
R240 VTAIL.n70 VTAIL.n69 0.155672
R241 VTAIL.n69 VTAIL.n45 0.155672
R242 VTAIL.n62 VTAIL.n45 0.155672
R243 VTAIL.n62 VTAIL.n61 0.155672
R244 VTAIL.n61 VTAIL.n49 0.155672
R245 VTAIL.n54 VTAIL.n49 0.155672
R246 VTAIL VTAIL.n159 0.142741
R247 VDD2.n73 VDD2.n39 756.745
R248 VDD2.n34 VDD2.n0 756.745
R249 VDD2.n74 VDD2.n73 585
R250 VDD2.n72 VDD2.n71 585
R251 VDD2.n43 VDD2.n42 585
R252 VDD2.n66 VDD2.n65 585
R253 VDD2.n64 VDD2.n63 585
R254 VDD2.n47 VDD2.n46 585
R255 VDD2.n58 VDD2.n57 585
R256 VDD2.n56 VDD2.n55 585
R257 VDD2.n51 VDD2.n50 585
R258 VDD2.n12 VDD2.n11 585
R259 VDD2.n17 VDD2.n16 585
R260 VDD2.n19 VDD2.n18 585
R261 VDD2.n8 VDD2.n7 585
R262 VDD2.n25 VDD2.n24 585
R263 VDD2.n27 VDD2.n26 585
R264 VDD2.n4 VDD2.n3 585
R265 VDD2.n33 VDD2.n32 585
R266 VDD2.n35 VDD2.n34 585
R267 VDD2.n52 VDD2.t0 327.483
R268 VDD2.n13 VDD2.t1 327.483
R269 VDD2.n73 VDD2.n72 171.744
R270 VDD2.n72 VDD2.n42 171.744
R271 VDD2.n65 VDD2.n42 171.744
R272 VDD2.n65 VDD2.n64 171.744
R273 VDD2.n64 VDD2.n46 171.744
R274 VDD2.n57 VDD2.n46 171.744
R275 VDD2.n57 VDD2.n56 171.744
R276 VDD2.n56 VDD2.n50 171.744
R277 VDD2.n17 VDD2.n11 171.744
R278 VDD2.n18 VDD2.n17 171.744
R279 VDD2.n18 VDD2.n7 171.744
R280 VDD2.n25 VDD2.n7 171.744
R281 VDD2.n26 VDD2.n25 171.744
R282 VDD2.n26 VDD2.n3 171.744
R283 VDD2.n33 VDD2.n3 171.744
R284 VDD2.n34 VDD2.n33 171.744
R285 VDD2.t0 VDD2.n50 85.8723
R286 VDD2.t1 VDD2.n11 85.8723
R287 VDD2.n78 VDD2.n38 80.7606
R288 VDD2.n78 VDD2.n77 49.0581
R289 VDD2.n52 VDD2.n51 16.3891
R290 VDD2.n13 VDD2.n12 16.3891
R291 VDD2.n55 VDD2.n54 12.8005
R292 VDD2.n16 VDD2.n15 12.8005
R293 VDD2.n58 VDD2.n49 12.0247
R294 VDD2.n19 VDD2.n10 12.0247
R295 VDD2.n59 VDD2.n47 11.249
R296 VDD2.n20 VDD2.n8 11.249
R297 VDD2.n63 VDD2.n62 10.4732
R298 VDD2.n24 VDD2.n23 10.4732
R299 VDD2.n66 VDD2.n45 9.69747
R300 VDD2.n27 VDD2.n6 9.69747
R301 VDD2.n77 VDD2.n76 9.45567
R302 VDD2.n38 VDD2.n37 9.45567
R303 VDD2.n76 VDD2.n75 9.3005
R304 VDD2.n41 VDD2.n40 9.3005
R305 VDD2.n70 VDD2.n69 9.3005
R306 VDD2.n68 VDD2.n67 9.3005
R307 VDD2.n45 VDD2.n44 9.3005
R308 VDD2.n62 VDD2.n61 9.3005
R309 VDD2.n60 VDD2.n59 9.3005
R310 VDD2.n49 VDD2.n48 9.3005
R311 VDD2.n54 VDD2.n53 9.3005
R312 VDD2.n37 VDD2.n36 9.3005
R313 VDD2.n31 VDD2.n30 9.3005
R314 VDD2.n29 VDD2.n28 9.3005
R315 VDD2.n6 VDD2.n5 9.3005
R316 VDD2.n23 VDD2.n22 9.3005
R317 VDD2.n21 VDD2.n20 9.3005
R318 VDD2.n10 VDD2.n9 9.3005
R319 VDD2.n15 VDD2.n14 9.3005
R320 VDD2.n2 VDD2.n1 9.3005
R321 VDD2.n67 VDD2.n43 8.92171
R322 VDD2.n28 VDD2.n4 8.92171
R323 VDD2.n71 VDD2.n70 8.14595
R324 VDD2.n32 VDD2.n31 8.14595
R325 VDD2.n77 VDD2.n39 7.3702
R326 VDD2.n74 VDD2.n41 7.3702
R327 VDD2.n35 VDD2.n2 7.3702
R328 VDD2.n38 VDD2.n0 7.3702
R329 VDD2.n75 VDD2.n39 6.59444
R330 VDD2.n75 VDD2.n74 6.59444
R331 VDD2.n36 VDD2.n35 6.59444
R332 VDD2.n36 VDD2.n0 6.59444
R333 VDD2.n71 VDD2.n41 5.81868
R334 VDD2.n32 VDD2.n2 5.81868
R335 VDD2.n70 VDD2.n43 5.04292
R336 VDD2.n31 VDD2.n4 5.04292
R337 VDD2.n67 VDD2.n66 4.26717
R338 VDD2.n28 VDD2.n27 4.26717
R339 VDD2.n53 VDD2.n52 3.71019
R340 VDD2.n14 VDD2.n13 3.71019
R341 VDD2.n63 VDD2.n45 3.49141
R342 VDD2.n24 VDD2.n6 3.49141
R343 VDD2.n62 VDD2.n47 2.71565
R344 VDD2.n23 VDD2.n8 2.71565
R345 VDD2.n59 VDD2.n58 1.93989
R346 VDD2.n20 VDD2.n19 1.93989
R347 VDD2.n55 VDD2.n49 1.16414
R348 VDD2.n16 VDD2.n10 1.16414
R349 VDD2.n54 VDD2.n51 0.388379
R350 VDD2.n15 VDD2.n12 0.388379
R351 VDD2 VDD2.n78 0.259121
R352 VDD2.n76 VDD2.n40 0.155672
R353 VDD2.n69 VDD2.n40 0.155672
R354 VDD2.n69 VDD2.n68 0.155672
R355 VDD2.n68 VDD2.n44 0.155672
R356 VDD2.n61 VDD2.n44 0.155672
R357 VDD2.n61 VDD2.n60 0.155672
R358 VDD2.n60 VDD2.n48 0.155672
R359 VDD2.n53 VDD2.n48 0.155672
R360 VDD2.n14 VDD2.n9 0.155672
R361 VDD2.n21 VDD2.n9 0.155672
R362 VDD2.n22 VDD2.n21 0.155672
R363 VDD2.n22 VDD2.n5 0.155672
R364 VDD2.n29 VDD2.n5 0.155672
R365 VDD2.n30 VDD2.n29 0.155672
R366 VDD2.n30 VDD2.n1 0.155672
R367 VDD2.n37 VDD2.n1 0.155672
R368 B.n222 B.n221 585
R369 B.n220 B.n61 585
R370 B.n219 B.n218 585
R371 B.n217 B.n62 585
R372 B.n216 B.n215 585
R373 B.n214 B.n63 585
R374 B.n213 B.n212 585
R375 B.n211 B.n64 585
R376 B.n210 B.n209 585
R377 B.n208 B.n65 585
R378 B.n207 B.n206 585
R379 B.n205 B.n66 585
R380 B.n204 B.n203 585
R381 B.n202 B.n67 585
R382 B.n201 B.n200 585
R383 B.n199 B.n68 585
R384 B.n198 B.n197 585
R385 B.n196 B.n69 585
R386 B.n195 B.n194 585
R387 B.n193 B.n70 585
R388 B.n192 B.n191 585
R389 B.n190 B.n71 585
R390 B.n189 B.n188 585
R391 B.n187 B.n72 585
R392 B.n186 B.n185 585
R393 B.n184 B.n73 585
R394 B.n183 B.n182 585
R395 B.n181 B.n74 585
R396 B.n179 B.n178 585
R397 B.n177 B.n77 585
R398 B.n176 B.n175 585
R399 B.n174 B.n78 585
R400 B.n173 B.n172 585
R401 B.n171 B.n79 585
R402 B.n170 B.n169 585
R403 B.n168 B.n80 585
R404 B.n167 B.n166 585
R405 B.n165 B.n81 585
R406 B.n164 B.n163 585
R407 B.n159 B.n82 585
R408 B.n158 B.n157 585
R409 B.n156 B.n83 585
R410 B.n155 B.n154 585
R411 B.n153 B.n84 585
R412 B.n152 B.n151 585
R413 B.n150 B.n85 585
R414 B.n149 B.n148 585
R415 B.n147 B.n86 585
R416 B.n146 B.n145 585
R417 B.n144 B.n87 585
R418 B.n143 B.n142 585
R419 B.n141 B.n88 585
R420 B.n140 B.n139 585
R421 B.n138 B.n89 585
R422 B.n137 B.n136 585
R423 B.n135 B.n90 585
R424 B.n134 B.n133 585
R425 B.n132 B.n91 585
R426 B.n131 B.n130 585
R427 B.n129 B.n92 585
R428 B.n128 B.n127 585
R429 B.n126 B.n93 585
R430 B.n125 B.n124 585
R431 B.n123 B.n94 585
R432 B.n122 B.n121 585
R433 B.n120 B.n95 585
R434 B.n223 B.n60 585
R435 B.n225 B.n224 585
R436 B.n226 B.n59 585
R437 B.n228 B.n227 585
R438 B.n229 B.n58 585
R439 B.n231 B.n230 585
R440 B.n232 B.n57 585
R441 B.n234 B.n233 585
R442 B.n235 B.n56 585
R443 B.n237 B.n236 585
R444 B.n238 B.n55 585
R445 B.n240 B.n239 585
R446 B.n241 B.n54 585
R447 B.n243 B.n242 585
R448 B.n244 B.n53 585
R449 B.n246 B.n245 585
R450 B.n247 B.n52 585
R451 B.n249 B.n248 585
R452 B.n250 B.n51 585
R453 B.n252 B.n251 585
R454 B.n253 B.n50 585
R455 B.n255 B.n254 585
R456 B.n256 B.n49 585
R457 B.n258 B.n257 585
R458 B.n259 B.n48 585
R459 B.n261 B.n260 585
R460 B.n262 B.n47 585
R461 B.n264 B.n263 585
R462 B.n364 B.n363 585
R463 B.n362 B.n9 585
R464 B.n361 B.n360 585
R465 B.n359 B.n10 585
R466 B.n358 B.n357 585
R467 B.n356 B.n11 585
R468 B.n355 B.n354 585
R469 B.n353 B.n12 585
R470 B.n352 B.n351 585
R471 B.n350 B.n13 585
R472 B.n349 B.n348 585
R473 B.n347 B.n14 585
R474 B.n346 B.n345 585
R475 B.n344 B.n15 585
R476 B.n343 B.n342 585
R477 B.n341 B.n16 585
R478 B.n340 B.n339 585
R479 B.n338 B.n17 585
R480 B.n337 B.n336 585
R481 B.n335 B.n18 585
R482 B.n334 B.n333 585
R483 B.n332 B.n19 585
R484 B.n331 B.n330 585
R485 B.n329 B.n20 585
R486 B.n328 B.n327 585
R487 B.n326 B.n21 585
R488 B.n325 B.n324 585
R489 B.n323 B.n22 585
R490 B.n322 B.n321 585
R491 B.n320 B.n23 585
R492 B.n319 B.n318 585
R493 B.n317 B.n27 585
R494 B.n316 B.n315 585
R495 B.n314 B.n28 585
R496 B.n313 B.n312 585
R497 B.n311 B.n29 585
R498 B.n310 B.n309 585
R499 B.n308 B.n30 585
R500 B.n306 B.n305 585
R501 B.n304 B.n33 585
R502 B.n303 B.n302 585
R503 B.n301 B.n34 585
R504 B.n300 B.n299 585
R505 B.n298 B.n35 585
R506 B.n297 B.n296 585
R507 B.n295 B.n36 585
R508 B.n294 B.n293 585
R509 B.n292 B.n37 585
R510 B.n291 B.n290 585
R511 B.n289 B.n38 585
R512 B.n288 B.n287 585
R513 B.n286 B.n39 585
R514 B.n285 B.n284 585
R515 B.n283 B.n40 585
R516 B.n282 B.n281 585
R517 B.n280 B.n41 585
R518 B.n279 B.n278 585
R519 B.n277 B.n42 585
R520 B.n276 B.n275 585
R521 B.n274 B.n43 585
R522 B.n273 B.n272 585
R523 B.n271 B.n44 585
R524 B.n270 B.n269 585
R525 B.n268 B.n45 585
R526 B.n267 B.n266 585
R527 B.n265 B.n46 585
R528 B.n365 B.n8 585
R529 B.n367 B.n366 585
R530 B.n368 B.n7 585
R531 B.n370 B.n369 585
R532 B.n371 B.n6 585
R533 B.n373 B.n372 585
R534 B.n374 B.n5 585
R535 B.n376 B.n375 585
R536 B.n377 B.n4 585
R537 B.n379 B.n378 585
R538 B.n380 B.n3 585
R539 B.n382 B.n381 585
R540 B.n383 B.n0 585
R541 B.n2 B.n1 585
R542 B.n102 B.n101 585
R543 B.n104 B.n103 585
R544 B.n105 B.n100 585
R545 B.n107 B.n106 585
R546 B.n108 B.n99 585
R547 B.n110 B.n109 585
R548 B.n111 B.n98 585
R549 B.n113 B.n112 585
R550 B.n114 B.n97 585
R551 B.n116 B.n115 585
R552 B.n117 B.n96 585
R553 B.n119 B.n118 585
R554 B.n120 B.n119 526.135
R555 B.n221 B.n60 526.135
R556 B.n263 B.n46 526.135
R557 B.n365 B.n364 526.135
R558 B.n160 B.t6 503.642
R559 B.n75 B.t3 503.642
R560 B.n31 B.t0 503.642
R561 B.n24 B.t9 503.642
R562 B.n75 B.t4 312.077
R563 B.n31 B.t2 312.077
R564 B.n160 B.t7 312.077
R565 B.n24 B.t11 312.077
R566 B.n76 B.t5 294.041
R567 B.n32 B.t1 294.041
R568 B.n161 B.t8 294.041
R569 B.n25 B.t10 294.041
R570 B.n385 B.n384 256.663
R571 B.n384 B.n383 235.042
R572 B.n384 B.n2 235.042
R573 B.n121 B.n120 163.367
R574 B.n121 B.n94 163.367
R575 B.n125 B.n94 163.367
R576 B.n126 B.n125 163.367
R577 B.n127 B.n126 163.367
R578 B.n127 B.n92 163.367
R579 B.n131 B.n92 163.367
R580 B.n132 B.n131 163.367
R581 B.n133 B.n132 163.367
R582 B.n133 B.n90 163.367
R583 B.n137 B.n90 163.367
R584 B.n138 B.n137 163.367
R585 B.n139 B.n138 163.367
R586 B.n139 B.n88 163.367
R587 B.n143 B.n88 163.367
R588 B.n144 B.n143 163.367
R589 B.n145 B.n144 163.367
R590 B.n145 B.n86 163.367
R591 B.n149 B.n86 163.367
R592 B.n150 B.n149 163.367
R593 B.n151 B.n150 163.367
R594 B.n151 B.n84 163.367
R595 B.n155 B.n84 163.367
R596 B.n156 B.n155 163.367
R597 B.n157 B.n156 163.367
R598 B.n157 B.n82 163.367
R599 B.n164 B.n82 163.367
R600 B.n165 B.n164 163.367
R601 B.n166 B.n165 163.367
R602 B.n166 B.n80 163.367
R603 B.n170 B.n80 163.367
R604 B.n171 B.n170 163.367
R605 B.n172 B.n171 163.367
R606 B.n172 B.n78 163.367
R607 B.n176 B.n78 163.367
R608 B.n177 B.n176 163.367
R609 B.n178 B.n177 163.367
R610 B.n178 B.n74 163.367
R611 B.n183 B.n74 163.367
R612 B.n184 B.n183 163.367
R613 B.n185 B.n184 163.367
R614 B.n185 B.n72 163.367
R615 B.n189 B.n72 163.367
R616 B.n190 B.n189 163.367
R617 B.n191 B.n190 163.367
R618 B.n191 B.n70 163.367
R619 B.n195 B.n70 163.367
R620 B.n196 B.n195 163.367
R621 B.n197 B.n196 163.367
R622 B.n197 B.n68 163.367
R623 B.n201 B.n68 163.367
R624 B.n202 B.n201 163.367
R625 B.n203 B.n202 163.367
R626 B.n203 B.n66 163.367
R627 B.n207 B.n66 163.367
R628 B.n208 B.n207 163.367
R629 B.n209 B.n208 163.367
R630 B.n209 B.n64 163.367
R631 B.n213 B.n64 163.367
R632 B.n214 B.n213 163.367
R633 B.n215 B.n214 163.367
R634 B.n215 B.n62 163.367
R635 B.n219 B.n62 163.367
R636 B.n220 B.n219 163.367
R637 B.n221 B.n220 163.367
R638 B.n263 B.n262 163.367
R639 B.n262 B.n261 163.367
R640 B.n261 B.n48 163.367
R641 B.n257 B.n48 163.367
R642 B.n257 B.n256 163.367
R643 B.n256 B.n255 163.367
R644 B.n255 B.n50 163.367
R645 B.n251 B.n50 163.367
R646 B.n251 B.n250 163.367
R647 B.n250 B.n249 163.367
R648 B.n249 B.n52 163.367
R649 B.n245 B.n52 163.367
R650 B.n245 B.n244 163.367
R651 B.n244 B.n243 163.367
R652 B.n243 B.n54 163.367
R653 B.n239 B.n54 163.367
R654 B.n239 B.n238 163.367
R655 B.n238 B.n237 163.367
R656 B.n237 B.n56 163.367
R657 B.n233 B.n56 163.367
R658 B.n233 B.n232 163.367
R659 B.n232 B.n231 163.367
R660 B.n231 B.n58 163.367
R661 B.n227 B.n58 163.367
R662 B.n227 B.n226 163.367
R663 B.n226 B.n225 163.367
R664 B.n225 B.n60 163.367
R665 B.n364 B.n9 163.367
R666 B.n360 B.n9 163.367
R667 B.n360 B.n359 163.367
R668 B.n359 B.n358 163.367
R669 B.n358 B.n11 163.367
R670 B.n354 B.n11 163.367
R671 B.n354 B.n353 163.367
R672 B.n353 B.n352 163.367
R673 B.n352 B.n13 163.367
R674 B.n348 B.n13 163.367
R675 B.n348 B.n347 163.367
R676 B.n347 B.n346 163.367
R677 B.n346 B.n15 163.367
R678 B.n342 B.n15 163.367
R679 B.n342 B.n341 163.367
R680 B.n341 B.n340 163.367
R681 B.n340 B.n17 163.367
R682 B.n336 B.n17 163.367
R683 B.n336 B.n335 163.367
R684 B.n335 B.n334 163.367
R685 B.n334 B.n19 163.367
R686 B.n330 B.n19 163.367
R687 B.n330 B.n329 163.367
R688 B.n329 B.n328 163.367
R689 B.n328 B.n21 163.367
R690 B.n324 B.n21 163.367
R691 B.n324 B.n323 163.367
R692 B.n323 B.n322 163.367
R693 B.n322 B.n23 163.367
R694 B.n318 B.n23 163.367
R695 B.n318 B.n317 163.367
R696 B.n317 B.n316 163.367
R697 B.n316 B.n28 163.367
R698 B.n312 B.n28 163.367
R699 B.n312 B.n311 163.367
R700 B.n311 B.n310 163.367
R701 B.n310 B.n30 163.367
R702 B.n305 B.n30 163.367
R703 B.n305 B.n304 163.367
R704 B.n304 B.n303 163.367
R705 B.n303 B.n34 163.367
R706 B.n299 B.n34 163.367
R707 B.n299 B.n298 163.367
R708 B.n298 B.n297 163.367
R709 B.n297 B.n36 163.367
R710 B.n293 B.n36 163.367
R711 B.n293 B.n292 163.367
R712 B.n292 B.n291 163.367
R713 B.n291 B.n38 163.367
R714 B.n287 B.n38 163.367
R715 B.n287 B.n286 163.367
R716 B.n286 B.n285 163.367
R717 B.n285 B.n40 163.367
R718 B.n281 B.n40 163.367
R719 B.n281 B.n280 163.367
R720 B.n280 B.n279 163.367
R721 B.n279 B.n42 163.367
R722 B.n275 B.n42 163.367
R723 B.n275 B.n274 163.367
R724 B.n274 B.n273 163.367
R725 B.n273 B.n44 163.367
R726 B.n269 B.n44 163.367
R727 B.n269 B.n268 163.367
R728 B.n268 B.n267 163.367
R729 B.n267 B.n46 163.367
R730 B.n366 B.n365 163.367
R731 B.n366 B.n7 163.367
R732 B.n370 B.n7 163.367
R733 B.n371 B.n370 163.367
R734 B.n372 B.n371 163.367
R735 B.n372 B.n5 163.367
R736 B.n376 B.n5 163.367
R737 B.n377 B.n376 163.367
R738 B.n378 B.n377 163.367
R739 B.n378 B.n3 163.367
R740 B.n382 B.n3 163.367
R741 B.n383 B.n382 163.367
R742 B.n102 B.n2 163.367
R743 B.n103 B.n102 163.367
R744 B.n103 B.n100 163.367
R745 B.n107 B.n100 163.367
R746 B.n108 B.n107 163.367
R747 B.n109 B.n108 163.367
R748 B.n109 B.n98 163.367
R749 B.n113 B.n98 163.367
R750 B.n114 B.n113 163.367
R751 B.n115 B.n114 163.367
R752 B.n115 B.n96 163.367
R753 B.n119 B.n96 163.367
R754 B.n162 B.n161 59.5399
R755 B.n180 B.n76 59.5399
R756 B.n307 B.n32 59.5399
R757 B.n26 B.n25 59.5399
R758 B.n363 B.n8 34.1859
R759 B.n265 B.n264 34.1859
R760 B.n223 B.n222 34.1859
R761 B.n118 B.n95 34.1859
R762 B B.n385 18.0485
R763 B.n161 B.n160 18.0369
R764 B.n76 B.n75 18.0369
R765 B.n32 B.n31 18.0369
R766 B.n25 B.n24 18.0369
R767 B.n367 B.n8 10.6151
R768 B.n368 B.n367 10.6151
R769 B.n369 B.n368 10.6151
R770 B.n369 B.n6 10.6151
R771 B.n373 B.n6 10.6151
R772 B.n374 B.n373 10.6151
R773 B.n375 B.n374 10.6151
R774 B.n375 B.n4 10.6151
R775 B.n379 B.n4 10.6151
R776 B.n380 B.n379 10.6151
R777 B.n381 B.n380 10.6151
R778 B.n381 B.n0 10.6151
R779 B.n363 B.n362 10.6151
R780 B.n362 B.n361 10.6151
R781 B.n361 B.n10 10.6151
R782 B.n357 B.n10 10.6151
R783 B.n357 B.n356 10.6151
R784 B.n356 B.n355 10.6151
R785 B.n355 B.n12 10.6151
R786 B.n351 B.n12 10.6151
R787 B.n351 B.n350 10.6151
R788 B.n350 B.n349 10.6151
R789 B.n349 B.n14 10.6151
R790 B.n345 B.n14 10.6151
R791 B.n345 B.n344 10.6151
R792 B.n344 B.n343 10.6151
R793 B.n343 B.n16 10.6151
R794 B.n339 B.n16 10.6151
R795 B.n339 B.n338 10.6151
R796 B.n338 B.n337 10.6151
R797 B.n337 B.n18 10.6151
R798 B.n333 B.n18 10.6151
R799 B.n333 B.n332 10.6151
R800 B.n332 B.n331 10.6151
R801 B.n331 B.n20 10.6151
R802 B.n327 B.n20 10.6151
R803 B.n327 B.n326 10.6151
R804 B.n326 B.n325 10.6151
R805 B.n325 B.n22 10.6151
R806 B.n321 B.n320 10.6151
R807 B.n320 B.n319 10.6151
R808 B.n319 B.n27 10.6151
R809 B.n315 B.n27 10.6151
R810 B.n315 B.n314 10.6151
R811 B.n314 B.n313 10.6151
R812 B.n313 B.n29 10.6151
R813 B.n309 B.n29 10.6151
R814 B.n309 B.n308 10.6151
R815 B.n306 B.n33 10.6151
R816 B.n302 B.n33 10.6151
R817 B.n302 B.n301 10.6151
R818 B.n301 B.n300 10.6151
R819 B.n300 B.n35 10.6151
R820 B.n296 B.n35 10.6151
R821 B.n296 B.n295 10.6151
R822 B.n295 B.n294 10.6151
R823 B.n294 B.n37 10.6151
R824 B.n290 B.n37 10.6151
R825 B.n290 B.n289 10.6151
R826 B.n289 B.n288 10.6151
R827 B.n288 B.n39 10.6151
R828 B.n284 B.n39 10.6151
R829 B.n284 B.n283 10.6151
R830 B.n283 B.n282 10.6151
R831 B.n282 B.n41 10.6151
R832 B.n278 B.n41 10.6151
R833 B.n278 B.n277 10.6151
R834 B.n277 B.n276 10.6151
R835 B.n276 B.n43 10.6151
R836 B.n272 B.n43 10.6151
R837 B.n272 B.n271 10.6151
R838 B.n271 B.n270 10.6151
R839 B.n270 B.n45 10.6151
R840 B.n266 B.n45 10.6151
R841 B.n266 B.n265 10.6151
R842 B.n264 B.n47 10.6151
R843 B.n260 B.n47 10.6151
R844 B.n260 B.n259 10.6151
R845 B.n259 B.n258 10.6151
R846 B.n258 B.n49 10.6151
R847 B.n254 B.n49 10.6151
R848 B.n254 B.n253 10.6151
R849 B.n253 B.n252 10.6151
R850 B.n252 B.n51 10.6151
R851 B.n248 B.n51 10.6151
R852 B.n248 B.n247 10.6151
R853 B.n247 B.n246 10.6151
R854 B.n246 B.n53 10.6151
R855 B.n242 B.n53 10.6151
R856 B.n242 B.n241 10.6151
R857 B.n241 B.n240 10.6151
R858 B.n240 B.n55 10.6151
R859 B.n236 B.n55 10.6151
R860 B.n236 B.n235 10.6151
R861 B.n235 B.n234 10.6151
R862 B.n234 B.n57 10.6151
R863 B.n230 B.n57 10.6151
R864 B.n230 B.n229 10.6151
R865 B.n229 B.n228 10.6151
R866 B.n228 B.n59 10.6151
R867 B.n224 B.n59 10.6151
R868 B.n224 B.n223 10.6151
R869 B.n101 B.n1 10.6151
R870 B.n104 B.n101 10.6151
R871 B.n105 B.n104 10.6151
R872 B.n106 B.n105 10.6151
R873 B.n106 B.n99 10.6151
R874 B.n110 B.n99 10.6151
R875 B.n111 B.n110 10.6151
R876 B.n112 B.n111 10.6151
R877 B.n112 B.n97 10.6151
R878 B.n116 B.n97 10.6151
R879 B.n117 B.n116 10.6151
R880 B.n118 B.n117 10.6151
R881 B.n122 B.n95 10.6151
R882 B.n123 B.n122 10.6151
R883 B.n124 B.n123 10.6151
R884 B.n124 B.n93 10.6151
R885 B.n128 B.n93 10.6151
R886 B.n129 B.n128 10.6151
R887 B.n130 B.n129 10.6151
R888 B.n130 B.n91 10.6151
R889 B.n134 B.n91 10.6151
R890 B.n135 B.n134 10.6151
R891 B.n136 B.n135 10.6151
R892 B.n136 B.n89 10.6151
R893 B.n140 B.n89 10.6151
R894 B.n141 B.n140 10.6151
R895 B.n142 B.n141 10.6151
R896 B.n142 B.n87 10.6151
R897 B.n146 B.n87 10.6151
R898 B.n147 B.n146 10.6151
R899 B.n148 B.n147 10.6151
R900 B.n148 B.n85 10.6151
R901 B.n152 B.n85 10.6151
R902 B.n153 B.n152 10.6151
R903 B.n154 B.n153 10.6151
R904 B.n154 B.n83 10.6151
R905 B.n158 B.n83 10.6151
R906 B.n159 B.n158 10.6151
R907 B.n163 B.n159 10.6151
R908 B.n167 B.n81 10.6151
R909 B.n168 B.n167 10.6151
R910 B.n169 B.n168 10.6151
R911 B.n169 B.n79 10.6151
R912 B.n173 B.n79 10.6151
R913 B.n174 B.n173 10.6151
R914 B.n175 B.n174 10.6151
R915 B.n175 B.n77 10.6151
R916 B.n179 B.n77 10.6151
R917 B.n182 B.n181 10.6151
R918 B.n182 B.n73 10.6151
R919 B.n186 B.n73 10.6151
R920 B.n187 B.n186 10.6151
R921 B.n188 B.n187 10.6151
R922 B.n188 B.n71 10.6151
R923 B.n192 B.n71 10.6151
R924 B.n193 B.n192 10.6151
R925 B.n194 B.n193 10.6151
R926 B.n194 B.n69 10.6151
R927 B.n198 B.n69 10.6151
R928 B.n199 B.n198 10.6151
R929 B.n200 B.n199 10.6151
R930 B.n200 B.n67 10.6151
R931 B.n204 B.n67 10.6151
R932 B.n205 B.n204 10.6151
R933 B.n206 B.n205 10.6151
R934 B.n206 B.n65 10.6151
R935 B.n210 B.n65 10.6151
R936 B.n211 B.n210 10.6151
R937 B.n212 B.n211 10.6151
R938 B.n212 B.n63 10.6151
R939 B.n216 B.n63 10.6151
R940 B.n217 B.n216 10.6151
R941 B.n218 B.n217 10.6151
R942 B.n218 B.n61 10.6151
R943 B.n222 B.n61 10.6151
R944 B.n26 B.n22 8.74196
R945 B.n307 B.n306 8.74196
R946 B.n163 B.n162 8.74196
R947 B.n181 B.n180 8.74196
R948 B.n385 B.n0 8.11757
R949 B.n385 B.n1 8.11757
R950 B.n321 B.n26 1.87367
R951 B.n308 B.n307 1.87367
R952 B.n162 B.n81 1.87367
R953 B.n180 B.n179 1.87367
R954 VP.n0 VP.t1 562.336
R955 VP.n0 VP.t0 526.415
R956 VP VP.n0 0.0516364
R957 VDD1.n34 VDD1.n0 756.745
R958 VDD1.n73 VDD1.n39 756.745
R959 VDD1.n35 VDD1.n34 585
R960 VDD1.n33 VDD1.n32 585
R961 VDD1.n4 VDD1.n3 585
R962 VDD1.n27 VDD1.n26 585
R963 VDD1.n25 VDD1.n24 585
R964 VDD1.n8 VDD1.n7 585
R965 VDD1.n19 VDD1.n18 585
R966 VDD1.n17 VDD1.n16 585
R967 VDD1.n12 VDD1.n11 585
R968 VDD1.n51 VDD1.n50 585
R969 VDD1.n56 VDD1.n55 585
R970 VDD1.n58 VDD1.n57 585
R971 VDD1.n47 VDD1.n46 585
R972 VDD1.n64 VDD1.n63 585
R973 VDD1.n66 VDD1.n65 585
R974 VDD1.n43 VDD1.n42 585
R975 VDD1.n72 VDD1.n71 585
R976 VDD1.n74 VDD1.n73 585
R977 VDD1.n13 VDD1.t0 327.483
R978 VDD1.n52 VDD1.t1 327.483
R979 VDD1.n34 VDD1.n33 171.744
R980 VDD1.n33 VDD1.n3 171.744
R981 VDD1.n26 VDD1.n3 171.744
R982 VDD1.n26 VDD1.n25 171.744
R983 VDD1.n25 VDD1.n7 171.744
R984 VDD1.n18 VDD1.n7 171.744
R985 VDD1.n18 VDD1.n17 171.744
R986 VDD1.n17 VDD1.n11 171.744
R987 VDD1.n56 VDD1.n50 171.744
R988 VDD1.n57 VDD1.n56 171.744
R989 VDD1.n57 VDD1.n46 171.744
R990 VDD1.n64 VDD1.n46 171.744
R991 VDD1.n65 VDD1.n64 171.744
R992 VDD1.n65 VDD1.n42 171.744
R993 VDD1.n72 VDD1.n42 171.744
R994 VDD1.n73 VDD1.n72 171.744
R995 VDD1.t0 VDD1.n11 85.8723
R996 VDD1.t1 VDD1.n50 85.8723
R997 VDD1 VDD1.n77 81.4859
R998 VDD1 VDD1.n38 49.3167
R999 VDD1.n13 VDD1.n12 16.3891
R1000 VDD1.n52 VDD1.n51 16.3891
R1001 VDD1.n16 VDD1.n15 12.8005
R1002 VDD1.n55 VDD1.n54 12.8005
R1003 VDD1.n19 VDD1.n10 12.0247
R1004 VDD1.n58 VDD1.n49 12.0247
R1005 VDD1.n20 VDD1.n8 11.249
R1006 VDD1.n59 VDD1.n47 11.249
R1007 VDD1.n24 VDD1.n23 10.4732
R1008 VDD1.n63 VDD1.n62 10.4732
R1009 VDD1.n27 VDD1.n6 9.69747
R1010 VDD1.n66 VDD1.n45 9.69747
R1011 VDD1.n38 VDD1.n37 9.45567
R1012 VDD1.n77 VDD1.n76 9.45567
R1013 VDD1.n37 VDD1.n36 9.3005
R1014 VDD1.n2 VDD1.n1 9.3005
R1015 VDD1.n31 VDD1.n30 9.3005
R1016 VDD1.n29 VDD1.n28 9.3005
R1017 VDD1.n6 VDD1.n5 9.3005
R1018 VDD1.n23 VDD1.n22 9.3005
R1019 VDD1.n21 VDD1.n20 9.3005
R1020 VDD1.n10 VDD1.n9 9.3005
R1021 VDD1.n15 VDD1.n14 9.3005
R1022 VDD1.n76 VDD1.n75 9.3005
R1023 VDD1.n70 VDD1.n69 9.3005
R1024 VDD1.n68 VDD1.n67 9.3005
R1025 VDD1.n45 VDD1.n44 9.3005
R1026 VDD1.n62 VDD1.n61 9.3005
R1027 VDD1.n60 VDD1.n59 9.3005
R1028 VDD1.n49 VDD1.n48 9.3005
R1029 VDD1.n54 VDD1.n53 9.3005
R1030 VDD1.n41 VDD1.n40 9.3005
R1031 VDD1.n28 VDD1.n4 8.92171
R1032 VDD1.n67 VDD1.n43 8.92171
R1033 VDD1.n32 VDD1.n31 8.14595
R1034 VDD1.n71 VDD1.n70 8.14595
R1035 VDD1.n38 VDD1.n0 7.3702
R1036 VDD1.n35 VDD1.n2 7.3702
R1037 VDD1.n74 VDD1.n41 7.3702
R1038 VDD1.n77 VDD1.n39 7.3702
R1039 VDD1.n36 VDD1.n0 6.59444
R1040 VDD1.n36 VDD1.n35 6.59444
R1041 VDD1.n75 VDD1.n74 6.59444
R1042 VDD1.n75 VDD1.n39 6.59444
R1043 VDD1.n32 VDD1.n2 5.81868
R1044 VDD1.n71 VDD1.n41 5.81868
R1045 VDD1.n31 VDD1.n4 5.04292
R1046 VDD1.n70 VDD1.n43 5.04292
R1047 VDD1.n28 VDD1.n27 4.26717
R1048 VDD1.n67 VDD1.n66 4.26717
R1049 VDD1.n14 VDD1.n13 3.71019
R1050 VDD1.n53 VDD1.n52 3.71019
R1051 VDD1.n24 VDD1.n6 3.49141
R1052 VDD1.n63 VDD1.n45 3.49141
R1053 VDD1.n23 VDD1.n8 2.71565
R1054 VDD1.n62 VDD1.n47 2.71565
R1055 VDD1.n20 VDD1.n19 1.93989
R1056 VDD1.n59 VDD1.n58 1.93989
R1057 VDD1.n16 VDD1.n10 1.16414
R1058 VDD1.n55 VDD1.n49 1.16414
R1059 VDD1.n15 VDD1.n12 0.388379
R1060 VDD1.n54 VDD1.n51 0.388379
R1061 VDD1.n37 VDD1.n1 0.155672
R1062 VDD1.n30 VDD1.n1 0.155672
R1063 VDD1.n30 VDD1.n29 0.155672
R1064 VDD1.n29 VDD1.n5 0.155672
R1065 VDD1.n22 VDD1.n5 0.155672
R1066 VDD1.n22 VDD1.n21 0.155672
R1067 VDD1.n21 VDD1.n9 0.155672
R1068 VDD1.n14 VDD1.n9 0.155672
R1069 VDD1.n53 VDD1.n48 0.155672
R1070 VDD1.n60 VDD1.n48 0.155672
R1071 VDD1.n61 VDD1.n60 0.155672
R1072 VDD1.n61 VDD1.n44 0.155672
R1073 VDD1.n68 VDD1.n44 0.155672
R1074 VDD1.n69 VDD1.n68 0.155672
R1075 VDD1.n69 VDD1.n40 0.155672
R1076 VDD1.n76 VDD1.n40 0.155672
C0 B VDD2 1.08255f
C1 VTAIL VN 0.93448f
C2 VP VTAIL 0.948917f
C3 VDD1 B 1.06872f
C4 VTAIL VDD2 4.12031f
C5 VDD1 VTAIL 4.08486f
C6 w_n1342_n2462# VN 1.60184f
C7 VP w_n1342_n2462# 1.76847f
C8 VTAIL B 1.86261f
C9 w_n1342_n2462# VDD2 1.22777f
C10 VP VN 3.67395f
C11 VDD1 w_n1342_n2462# 1.22413f
C12 VDD2 VN 1.25203f
C13 VDD1 VN 0.148543f
C14 VP VDD2 0.250128f
C15 w_n1342_n2462# B 5.376009f
C16 VDD1 VP 1.35074f
C17 VDD1 VDD2 0.451376f
C18 B VN 0.656697f
C19 w_n1342_n2462# VTAIL 2.17554f
C20 VP B 0.922625f
C21 VDD2 VSUBS 0.57873f
C22 VDD1 VSUBS 2.160297f
C23 VTAIL VSUBS 0.577435f
C24 VN VSUBS 3.98307f
C25 VP VSUBS 0.907275f
C26 B VSUBS 2.036955f
C27 w_n1342_n2462# VSUBS 41.0491f
C28 VDD1.n0 VSUBS 0.01819f
C29 VDD1.n1 VSUBS 0.016058f
C30 VDD1.n2 VSUBS 0.008629f
C31 VDD1.n3 VSUBS 0.020396f
C32 VDD1.n4 VSUBS 0.009136f
C33 VDD1.n5 VSUBS 0.016058f
C34 VDD1.n6 VSUBS 0.008629f
C35 VDD1.n7 VSUBS 0.020396f
C36 VDD1.n8 VSUBS 0.009136f
C37 VDD1.n9 VSUBS 0.016058f
C38 VDD1.n10 VSUBS 0.008629f
C39 VDD1.n11 VSUBS 0.015297f
C40 VDD1.n12 VSUBS 0.012974f
C41 VDD1.t0 VSUBS 0.043551f
C42 VDD1.n13 VSUBS 0.077622f
C43 VDD1.n14 VSUBS 0.474576f
C44 VDD1.n15 VSUBS 0.008629f
C45 VDD1.n16 VSUBS 0.009136f
C46 VDD1.n17 VSUBS 0.020396f
C47 VDD1.n18 VSUBS 0.020396f
C48 VDD1.n19 VSUBS 0.009136f
C49 VDD1.n20 VSUBS 0.008629f
C50 VDD1.n21 VSUBS 0.016058f
C51 VDD1.n22 VSUBS 0.016058f
C52 VDD1.n23 VSUBS 0.008629f
C53 VDD1.n24 VSUBS 0.009136f
C54 VDD1.n25 VSUBS 0.020396f
C55 VDD1.n26 VSUBS 0.020396f
C56 VDD1.n27 VSUBS 0.009136f
C57 VDD1.n28 VSUBS 0.008629f
C58 VDD1.n29 VSUBS 0.016058f
C59 VDD1.n30 VSUBS 0.016058f
C60 VDD1.n31 VSUBS 0.008629f
C61 VDD1.n32 VSUBS 0.009136f
C62 VDD1.n33 VSUBS 0.020396f
C63 VDD1.n34 VSUBS 0.051234f
C64 VDD1.n35 VSUBS 0.009136f
C65 VDD1.n36 VSUBS 0.008629f
C66 VDD1.n37 VSUBS 0.037337f
C67 VDD1.n38 VSUBS 0.037173f
C68 VDD1.n39 VSUBS 0.01819f
C69 VDD1.n40 VSUBS 0.016058f
C70 VDD1.n41 VSUBS 0.008629f
C71 VDD1.n42 VSUBS 0.020396f
C72 VDD1.n43 VSUBS 0.009136f
C73 VDD1.n44 VSUBS 0.016058f
C74 VDD1.n45 VSUBS 0.008629f
C75 VDD1.n46 VSUBS 0.020396f
C76 VDD1.n47 VSUBS 0.009136f
C77 VDD1.n48 VSUBS 0.016058f
C78 VDD1.n49 VSUBS 0.008629f
C79 VDD1.n50 VSUBS 0.015297f
C80 VDD1.n51 VSUBS 0.012974f
C81 VDD1.t1 VSUBS 0.043551f
C82 VDD1.n52 VSUBS 0.077622f
C83 VDD1.n53 VSUBS 0.474576f
C84 VDD1.n54 VSUBS 0.008629f
C85 VDD1.n55 VSUBS 0.009136f
C86 VDD1.n56 VSUBS 0.020396f
C87 VDD1.n57 VSUBS 0.020396f
C88 VDD1.n58 VSUBS 0.009136f
C89 VDD1.n59 VSUBS 0.008629f
C90 VDD1.n60 VSUBS 0.016058f
C91 VDD1.n61 VSUBS 0.016058f
C92 VDD1.n62 VSUBS 0.008629f
C93 VDD1.n63 VSUBS 0.009136f
C94 VDD1.n64 VSUBS 0.020396f
C95 VDD1.n65 VSUBS 0.020396f
C96 VDD1.n66 VSUBS 0.009136f
C97 VDD1.n67 VSUBS 0.008629f
C98 VDD1.n68 VSUBS 0.016058f
C99 VDD1.n69 VSUBS 0.016058f
C100 VDD1.n70 VSUBS 0.008629f
C101 VDD1.n71 VSUBS 0.009136f
C102 VDD1.n72 VSUBS 0.020396f
C103 VDD1.n73 VSUBS 0.051234f
C104 VDD1.n74 VSUBS 0.009136f
C105 VDD1.n75 VSUBS 0.008629f
C106 VDD1.n76 VSUBS 0.037337f
C107 VDD1.n77 VSUBS 0.31827f
C108 VP.t1 VSUBS 0.619079f
C109 VP.t0 VSUBS 0.536358f
C110 VP.n0 VSUBS 2.53401f
C111 B.n0 VSUBS 0.005481f
C112 B.n1 VSUBS 0.005481f
C113 B.n2 VSUBS 0.008107f
C114 B.n3 VSUBS 0.006212f
C115 B.n4 VSUBS 0.006212f
C116 B.n5 VSUBS 0.006212f
C117 B.n6 VSUBS 0.006212f
C118 B.n7 VSUBS 0.006212f
C119 B.n8 VSUBS 0.014649f
C120 B.n9 VSUBS 0.006212f
C121 B.n10 VSUBS 0.006212f
C122 B.n11 VSUBS 0.006212f
C123 B.n12 VSUBS 0.006212f
C124 B.n13 VSUBS 0.006212f
C125 B.n14 VSUBS 0.006212f
C126 B.n15 VSUBS 0.006212f
C127 B.n16 VSUBS 0.006212f
C128 B.n17 VSUBS 0.006212f
C129 B.n18 VSUBS 0.006212f
C130 B.n19 VSUBS 0.006212f
C131 B.n20 VSUBS 0.006212f
C132 B.n21 VSUBS 0.006212f
C133 B.n22 VSUBS 0.005664f
C134 B.n23 VSUBS 0.006212f
C135 B.t10 VSUBS 0.103141f
C136 B.t11 VSUBS 0.111546f
C137 B.t9 VSUBS 0.167031f
C138 B.n24 VSUBS 0.180884f
C139 B.n25 VSUBS 0.154287f
C140 B.n26 VSUBS 0.014393f
C141 B.n27 VSUBS 0.006212f
C142 B.n28 VSUBS 0.006212f
C143 B.n29 VSUBS 0.006212f
C144 B.n30 VSUBS 0.006212f
C145 B.t1 VSUBS 0.103143f
C146 B.t2 VSUBS 0.111548f
C147 B.t0 VSUBS 0.167031f
C148 B.n31 VSUBS 0.180882f
C149 B.n32 VSUBS 0.154285f
C150 B.n33 VSUBS 0.006212f
C151 B.n34 VSUBS 0.006212f
C152 B.n35 VSUBS 0.006212f
C153 B.n36 VSUBS 0.006212f
C154 B.n37 VSUBS 0.006212f
C155 B.n38 VSUBS 0.006212f
C156 B.n39 VSUBS 0.006212f
C157 B.n40 VSUBS 0.006212f
C158 B.n41 VSUBS 0.006212f
C159 B.n42 VSUBS 0.006212f
C160 B.n43 VSUBS 0.006212f
C161 B.n44 VSUBS 0.006212f
C162 B.n45 VSUBS 0.006212f
C163 B.n46 VSUBS 0.015316f
C164 B.n47 VSUBS 0.006212f
C165 B.n48 VSUBS 0.006212f
C166 B.n49 VSUBS 0.006212f
C167 B.n50 VSUBS 0.006212f
C168 B.n51 VSUBS 0.006212f
C169 B.n52 VSUBS 0.006212f
C170 B.n53 VSUBS 0.006212f
C171 B.n54 VSUBS 0.006212f
C172 B.n55 VSUBS 0.006212f
C173 B.n56 VSUBS 0.006212f
C174 B.n57 VSUBS 0.006212f
C175 B.n58 VSUBS 0.006212f
C176 B.n59 VSUBS 0.006212f
C177 B.n60 VSUBS 0.014649f
C178 B.n61 VSUBS 0.006212f
C179 B.n62 VSUBS 0.006212f
C180 B.n63 VSUBS 0.006212f
C181 B.n64 VSUBS 0.006212f
C182 B.n65 VSUBS 0.006212f
C183 B.n66 VSUBS 0.006212f
C184 B.n67 VSUBS 0.006212f
C185 B.n68 VSUBS 0.006212f
C186 B.n69 VSUBS 0.006212f
C187 B.n70 VSUBS 0.006212f
C188 B.n71 VSUBS 0.006212f
C189 B.n72 VSUBS 0.006212f
C190 B.n73 VSUBS 0.006212f
C191 B.n74 VSUBS 0.006212f
C192 B.t5 VSUBS 0.103143f
C193 B.t4 VSUBS 0.111548f
C194 B.t3 VSUBS 0.167031f
C195 B.n75 VSUBS 0.180882f
C196 B.n76 VSUBS 0.154285f
C197 B.n77 VSUBS 0.006212f
C198 B.n78 VSUBS 0.006212f
C199 B.n79 VSUBS 0.006212f
C200 B.n80 VSUBS 0.006212f
C201 B.n81 VSUBS 0.003654f
C202 B.n82 VSUBS 0.006212f
C203 B.n83 VSUBS 0.006212f
C204 B.n84 VSUBS 0.006212f
C205 B.n85 VSUBS 0.006212f
C206 B.n86 VSUBS 0.006212f
C207 B.n87 VSUBS 0.006212f
C208 B.n88 VSUBS 0.006212f
C209 B.n89 VSUBS 0.006212f
C210 B.n90 VSUBS 0.006212f
C211 B.n91 VSUBS 0.006212f
C212 B.n92 VSUBS 0.006212f
C213 B.n93 VSUBS 0.006212f
C214 B.n94 VSUBS 0.006212f
C215 B.n95 VSUBS 0.015316f
C216 B.n96 VSUBS 0.006212f
C217 B.n97 VSUBS 0.006212f
C218 B.n98 VSUBS 0.006212f
C219 B.n99 VSUBS 0.006212f
C220 B.n100 VSUBS 0.006212f
C221 B.n101 VSUBS 0.006212f
C222 B.n102 VSUBS 0.006212f
C223 B.n103 VSUBS 0.006212f
C224 B.n104 VSUBS 0.006212f
C225 B.n105 VSUBS 0.006212f
C226 B.n106 VSUBS 0.006212f
C227 B.n107 VSUBS 0.006212f
C228 B.n108 VSUBS 0.006212f
C229 B.n109 VSUBS 0.006212f
C230 B.n110 VSUBS 0.006212f
C231 B.n111 VSUBS 0.006212f
C232 B.n112 VSUBS 0.006212f
C233 B.n113 VSUBS 0.006212f
C234 B.n114 VSUBS 0.006212f
C235 B.n115 VSUBS 0.006212f
C236 B.n116 VSUBS 0.006212f
C237 B.n117 VSUBS 0.006212f
C238 B.n118 VSUBS 0.014649f
C239 B.n119 VSUBS 0.014649f
C240 B.n120 VSUBS 0.015316f
C241 B.n121 VSUBS 0.006212f
C242 B.n122 VSUBS 0.006212f
C243 B.n123 VSUBS 0.006212f
C244 B.n124 VSUBS 0.006212f
C245 B.n125 VSUBS 0.006212f
C246 B.n126 VSUBS 0.006212f
C247 B.n127 VSUBS 0.006212f
C248 B.n128 VSUBS 0.006212f
C249 B.n129 VSUBS 0.006212f
C250 B.n130 VSUBS 0.006212f
C251 B.n131 VSUBS 0.006212f
C252 B.n132 VSUBS 0.006212f
C253 B.n133 VSUBS 0.006212f
C254 B.n134 VSUBS 0.006212f
C255 B.n135 VSUBS 0.006212f
C256 B.n136 VSUBS 0.006212f
C257 B.n137 VSUBS 0.006212f
C258 B.n138 VSUBS 0.006212f
C259 B.n139 VSUBS 0.006212f
C260 B.n140 VSUBS 0.006212f
C261 B.n141 VSUBS 0.006212f
C262 B.n142 VSUBS 0.006212f
C263 B.n143 VSUBS 0.006212f
C264 B.n144 VSUBS 0.006212f
C265 B.n145 VSUBS 0.006212f
C266 B.n146 VSUBS 0.006212f
C267 B.n147 VSUBS 0.006212f
C268 B.n148 VSUBS 0.006212f
C269 B.n149 VSUBS 0.006212f
C270 B.n150 VSUBS 0.006212f
C271 B.n151 VSUBS 0.006212f
C272 B.n152 VSUBS 0.006212f
C273 B.n153 VSUBS 0.006212f
C274 B.n154 VSUBS 0.006212f
C275 B.n155 VSUBS 0.006212f
C276 B.n156 VSUBS 0.006212f
C277 B.n157 VSUBS 0.006212f
C278 B.n158 VSUBS 0.006212f
C279 B.n159 VSUBS 0.006212f
C280 B.t8 VSUBS 0.103141f
C281 B.t7 VSUBS 0.111546f
C282 B.t6 VSUBS 0.167031f
C283 B.n160 VSUBS 0.180884f
C284 B.n161 VSUBS 0.154287f
C285 B.n162 VSUBS 0.014393f
C286 B.n163 VSUBS 0.005664f
C287 B.n164 VSUBS 0.006212f
C288 B.n165 VSUBS 0.006212f
C289 B.n166 VSUBS 0.006212f
C290 B.n167 VSUBS 0.006212f
C291 B.n168 VSUBS 0.006212f
C292 B.n169 VSUBS 0.006212f
C293 B.n170 VSUBS 0.006212f
C294 B.n171 VSUBS 0.006212f
C295 B.n172 VSUBS 0.006212f
C296 B.n173 VSUBS 0.006212f
C297 B.n174 VSUBS 0.006212f
C298 B.n175 VSUBS 0.006212f
C299 B.n176 VSUBS 0.006212f
C300 B.n177 VSUBS 0.006212f
C301 B.n178 VSUBS 0.006212f
C302 B.n179 VSUBS 0.003654f
C303 B.n180 VSUBS 0.014393f
C304 B.n181 VSUBS 0.005664f
C305 B.n182 VSUBS 0.006212f
C306 B.n183 VSUBS 0.006212f
C307 B.n184 VSUBS 0.006212f
C308 B.n185 VSUBS 0.006212f
C309 B.n186 VSUBS 0.006212f
C310 B.n187 VSUBS 0.006212f
C311 B.n188 VSUBS 0.006212f
C312 B.n189 VSUBS 0.006212f
C313 B.n190 VSUBS 0.006212f
C314 B.n191 VSUBS 0.006212f
C315 B.n192 VSUBS 0.006212f
C316 B.n193 VSUBS 0.006212f
C317 B.n194 VSUBS 0.006212f
C318 B.n195 VSUBS 0.006212f
C319 B.n196 VSUBS 0.006212f
C320 B.n197 VSUBS 0.006212f
C321 B.n198 VSUBS 0.006212f
C322 B.n199 VSUBS 0.006212f
C323 B.n200 VSUBS 0.006212f
C324 B.n201 VSUBS 0.006212f
C325 B.n202 VSUBS 0.006212f
C326 B.n203 VSUBS 0.006212f
C327 B.n204 VSUBS 0.006212f
C328 B.n205 VSUBS 0.006212f
C329 B.n206 VSUBS 0.006212f
C330 B.n207 VSUBS 0.006212f
C331 B.n208 VSUBS 0.006212f
C332 B.n209 VSUBS 0.006212f
C333 B.n210 VSUBS 0.006212f
C334 B.n211 VSUBS 0.006212f
C335 B.n212 VSUBS 0.006212f
C336 B.n213 VSUBS 0.006212f
C337 B.n214 VSUBS 0.006212f
C338 B.n215 VSUBS 0.006212f
C339 B.n216 VSUBS 0.006212f
C340 B.n217 VSUBS 0.006212f
C341 B.n218 VSUBS 0.006212f
C342 B.n219 VSUBS 0.006212f
C343 B.n220 VSUBS 0.006212f
C344 B.n221 VSUBS 0.015316f
C345 B.n222 VSUBS 0.014615f
C346 B.n223 VSUBS 0.01535f
C347 B.n224 VSUBS 0.006212f
C348 B.n225 VSUBS 0.006212f
C349 B.n226 VSUBS 0.006212f
C350 B.n227 VSUBS 0.006212f
C351 B.n228 VSUBS 0.006212f
C352 B.n229 VSUBS 0.006212f
C353 B.n230 VSUBS 0.006212f
C354 B.n231 VSUBS 0.006212f
C355 B.n232 VSUBS 0.006212f
C356 B.n233 VSUBS 0.006212f
C357 B.n234 VSUBS 0.006212f
C358 B.n235 VSUBS 0.006212f
C359 B.n236 VSUBS 0.006212f
C360 B.n237 VSUBS 0.006212f
C361 B.n238 VSUBS 0.006212f
C362 B.n239 VSUBS 0.006212f
C363 B.n240 VSUBS 0.006212f
C364 B.n241 VSUBS 0.006212f
C365 B.n242 VSUBS 0.006212f
C366 B.n243 VSUBS 0.006212f
C367 B.n244 VSUBS 0.006212f
C368 B.n245 VSUBS 0.006212f
C369 B.n246 VSUBS 0.006212f
C370 B.n247 VSUBS 0.006212f
C371 B.n248 VSUBS 0.006212f
C372 B.n249 VSUBS 0.006212f
C373 B.n250 VSUBS 0.006212f
C374 B.n251 VSUBS 0.006212f
C375 B.n252 VSUBS 0.006212f
C376 B.n253 VSUBS 0.006212f
C377 B.n254 VSUBS 0.006212f
C378 B.n255 VSUBS 0.006212f
C379 B.n256 VSUBS 0.006212f
C380 B.n257 VSUBS 0.006212f
C381 B.n258 VSUBS 0.006212f
C382 B.n259 VSUBS 0.006212f
C383 B.n260 VSUBS 0.006212f
C384 B.n261 VSUBS 0.006212f
C385 B.n262 VSUBS 0.006212f
C386 B.n263 VSUBS 0.014649f
C387 B.n264 VSUBS 0.014649f
C388 B.n265 VSUBS 0.015316f
C389 B.n266 VSUBS 0.006212f
C390 B.n267 VSUBS 0.006212f
C391 B.n268 VSUBS 0.006212f
C392 B.n269 VSUBS 0.006212f
C393 B.n270 VSUBS 0.006212f
C394 B.n271 VSUBS 0.006212f
C395 B.n272 VSUBS 0.006212f
C396 B.n273 VSUBS 0.006212f
C397 B.n274 VSUBS 0.006212f
C398 B.n275 VSUBS 0.006212f
C399 B.n276 VSUBS 0.006212f
C400 B.n277 VSUBS 0.006212f
C401 B.n278 VSUBS 0.006212f
C402 B.n279 VSUBS 0.006212f
C403 B.n280 VSUBS 0.006212f
C404 B.n281 VSUBS 0.006212f
C405 B.n282 VSUBS 0.006212f
C406 B.n283 VSUBS 0.006212f
C407 B.n284 VSUBS 0.006212f
C408 B.n285 VSUBS 0.006212f
C409 B.n286 VSUBS 0.006212f
C410 B.n287 VSUBS 0.006212f
C411 B.n288 VSUBS 0.006212f
C412 B.n289 VSUBS 0.006212f
C413 B.n290 VSUBS 0.006212f
C414 B.n291 VSUBS 0.006212f
C415 B.n292 VSUBS 0.006212f
C416 B.n293 VSUBS 0.006212f
C417 B.n294 VSUBS 0.006212f
C418 B.n295 VSUBS 0.006212f
C419 B.n296 VSUBS 0.006212f
C420 B.n297 VSUBS 0.006212f
C421 B.n298 VSUBS 0.006212f
C422 B.n299 VSUBS 0.006212f
C423 B.n300 VSUBS 0.006212f
C424 B.n301 VSUBS 0.006212f
C425 B.n302 VSUBS 0.006212f
C426 B.n303 VSUBS 0.006212f
C427 B.n304 VSUBS 0.006212f
C428 B.n305 VSUBS 0.006212f
C429 B.n306 VSUBS 0.005664f
C430 B.n307 VSUBS 0.014393f
C431 B.n308 VSUBS 0.003654f
C432 B.n309 VSUBS 0.006212f
C433 B.n310 VSUBS 0.006212f
C434 B.n311 VSUBS 0.006212f
C435 B.n312 VSUBS 0.006212f
C436 B.n313 VSUBS 0.006212f
C437 B.n314 VSUBS 0.006212f
C438 B.n315 VSUBS 0.006212f
C439 B.n316 VSUBS 0.006212f
C440 B.n317 VSUBS 0.006212f
C441 B.n318 VSUBS 0.006212f
C442 B.n319 VSUBS 0.006212f
C443 B.n320 VSUBS 0.006212f
C444 B.n321 VSUBS 0.003654f
C445 B.n322 VSUBS 0.006212f
C446 B.n323 VSUBS 0.006212f
C447 B.n324 VSUBS 0.006212f
C448 B.n325 VSUBS 0.006212f
C449 B.n326 VSUBS 0.006212f
C450 B.n327 VSUBS 0.006212f
C451 B.n328 VSUBS 0.006212f
C452 B.n329 VSUBS 0.006212f
C453 B.n330 VSUBS 0.006212f
C454 B.n331 VSUBS 0.006212f
C455 B.n332 VSUBS 0.006212f
C456 B.n333 VSUBS 0.006212f
C457 B.n334 VSUBS 0.006212f
C458 B.n335 VSUBS 0.006212f
C459 B.n336 VSUBS 0.006212f
C460 B.n337 VSUBS 0.006212f
C461 B.n338 VSUBS 0.006212f
C462 B.n339 VSUBS 0.006212f
C463 B.n340 VSUBS 0.006212f
C464 B.n341 VSUBS 0.006212f
C465 B.n342 VSUBS 0.006212f
C466 B.n343 VSUBS 0.006212f
C467 B.n344 VSUBS 0.006212f
C468 B.n345 VSUBS 0.006212f
C469 B.n346 VSUBS 0.006212f
C470 B.n347 VSUBS 0.006212f
C471 B.n348 VSUBS 0.006212f
C472 B.n349 VSUBS 0.006212f
C473 B.n350 VSUBS 0.006212f
C474 B.n351 VSUBS 0.006212f
C475 B.n352 VSUBS 0.006212f
C476 B.n353 VSUBS 0.006212f
C477 B.n354 VSUBS 0.006212f
C478 B.n355 VSUBS 0.006212f
C479 B.n356 VSUBS 0.006212f
C480 B.n357 VSUBS 0.006212f
C481 B.n358 VSUBS 0.006212f
C482 B.n359 VSUBS 0.006212f
C483 B.n360 VSUBS 0.006212f
C484 B.n361 VSUBS 0.006212f
C485 B.n362 VSUBS 0.006212f
C486 B.n363 VSUBS 0.015316f
C487 B.n364 VSUBS 0.015316f
C488 B.n365 VSUBS 0.014649f
C489 B.n366 VSUBS 0.006212f
C490 B.n367 VSUBS 0.006212f
C491 B.n368 VSUBS 0.006212f
C492 B.n369 VSUBS 0.006212f
C493 B.n370 VSUBS 0.006212f
C494 B.n371 VSUBS 0.006212f
C495 B.n372 VSUBS 0.006212f
C496 B.n373 VSUBS 0.006212f
C497 B.n374 VSUBS 0.006212f
C498 B.n375 VSUBS 0.006212f
C499 B.n376 VSUBS 0.006212f
C500 B.n377 VSUBS 0.006212f
C501 B.n378 VSUBS 0.006212f
C502 B.n379 VSUBS 0.006212f
C503 B.n380 VSUBS 0.006212f
C504 B.n381 VSUBS 0.006212f
C505 B.n382 VSUBS 0.006212f
C506 B.n383 VSUBS 0.008107f
C507 B.n384 VSUBS 0.008636f
C508 B.n385 VSUBS 0.017173f
C509 VDD2.n0 VSUBS 0.018457f
C510 VDD2.n1 VSUBS 0.016294f
C511 VDD2.n2 VSUBS 0.008756f
C512 VDD2.n3 VSUBS 0.020695f
C513 VDD2.n4 VSUBS 0.009271f
C514 VDD2.n5 VSUBS 0.016294f
C515 VDD2.n6 VSUBS 0.008756f
C516 VDD2.n7 VSUBS 0.020695f
C517 VDD2.n8 VSUBS 0.009271f
C518 VDD2.n9 VSUBS 0.016294f
C519 VDD2.n10 VSUBS 0.008756f
C520 VDD2.n11 VSUBS 0.015521f
C521 VDD2.n12 VSUBS 0.013164f
C522 VDD2.t1 VSUBS 0.04419f
C523 VDD2.n13 VSUBS 0.078761f
C524 VDD2.n14 VSUBS 0.481542f
C525 VDD2.n15 VSUBS 0.008756f
C526 VDD2.n16 VSUBS 0.009271f
C527 VDD2.n17 VSUBS 0.020695f
C528 VDD2.n18 VSUBS 0.020695f
C529 VDD2.n19 VSUBS 0.009271f
C530 VDD2.n20 VSUBS 0.008756f
C531 VDD2.n21 VSUBS 0.016294f
C532 VDD2.n22 VSUBS 0.016294f
C533 VDD2.n23 VSUBS 0.008756f
C534 VDD2.n24 VSUBS 0.009271f
C535 VDD2.n25 VSUBS 0.020695f
C536 VDD2.n26 VSUBS 0.020695f
C537 VDD2.n27 VSUBS 0.009271f
C538 VDD2.n28 VSUBS 0.008756f
C539 VDD2.n29 VSUBS 0.016294f
C540 VDD2.n30 VSUBS 0.016294f
C541 VDD2.n31 VSUBS 0.008756f
C542 VDD2.n32 VSUBS 0.009271f
C543 VDD2.n33 VSUBS 0.020695f
C544 VDD2.n34 VSUBS 0.051986f
C545 VDD2.n35 VSUBS 0.009271f
C546 VDD2.n36 VSUBS 0.008756f
C547 VDD2.n37 VSUBS 0.037885f
C548 VDD2.n38 VSUBS 0.303515f
C549 VDD2.n39 VSUBS 0.018457f
C550 VDD2.n40 VSUBS 0.016294f
C551 VDD2.n41 VSUBS 0.008756f
C552 VDD2.n42 VSUBS 0.020695f
C553 VDD2.n43 VSUBS 0.009271f
C554 VDD2.n44 VSUBS 0.016294f
C555 VDD2.n45 VSUBS 0.008756f
C556 VDD2.n46 VSUBS 0.020695f
C557 VDD2.n47 VSUBS 0.009271f
C558 VDD2.n48 VSUBS 0.016294f
C559 VDD2.n49 VSUBS 0.008756f
C560 VDD2.n50 VSUBS 0.015521f
C561 VDD2.n51 VSUBS 0.013164f
C562 VDD2.t0 VSUBS 0.04419f
C563 VDD2.n52 VSUBS 0.078761f
C564 VDD2.n53 VSUBS 0.481542f
C565 VDD2.n54 VSUBS 0.008756f
C566 VDD2.n55 VSUBS 0.009271f
C567 VDD2.n56 VSUBS 0.020695f
C568 VDD2.n57 VSUBS 0.020695f
C569 VDD2.n58 VSUBS 0.009271f
C570 VDD2.n59 VSUBS 0.008756f
C571 VDD2.n60 VSUBS 0.016294f
C572 VDD2.n61 VSUBS 0.016294f
C573 VDD2.n62 VSUBS 0.008756f
C574 VDD2.n63 VSUBS 0.009271f
C575 VDD2.n64 VSUBS 0.020695f
C576 VDD2.n65 VSUBS 0.020695f
C577 VDD2.n66 VSUBS 0.009271f
C578 VDD2.n67 VSUBS 0.008756f
C579 VDD2.n68 VSUBS 0.016294f
C580 VDD2.n69 VSUBS 0.016294f
C581 VDD2.n70 VSUBS 0.008756f
C582 VDD2.n71 VSUBS 0.009271f
C583 VDD2.n72 VSUBS 0.020695f
C584 VDD2.n73 VSUBS 0.051986f
C585 VDD2.n74 VSUBS 0.009271f
C586 VDD2.n75 VSUBS 0.008756f
C587 VDD2.n76 VSUBS 0.037885f
C588 VDD2.n77 VSUBS 0.037482f
C589 VDD2.n78 VSUBS 1.41714f
C590 VTAIL.n0 VSUBS 0.025773f
C591 VTAIL.n1 VSUBS 0.022752f
C592 VTAIL.n2 VSUBS 0.012226f
C593 VTAIL.n3 VSUBS 0.028898f
C594 VTAIL.n4 VSUBS 0.012945f
C595 VTAIL.n5 VSUBS 0.022752f
C596 VTAIL.n6 VSUBS 0.012226f
C597 VTAIL.n7 VSUBS 0.028898f
C598 VTAIL.n8 VSUBS 0.012945f
C599 VTAIL.n9 VSUBS 0.022752f
C600 VTAIL.n10 VSUBS 0.012226f
C601 VTAIL.n11 VSUBS 0.021674f
C602 VTAIL.n12 VSUBS 0.018382f
C603 VTAIL.t0 VSUBS 0.061707f
C604 VTAIL.n13 VSUBS 0.109981f
C605 VTAIL.n14 VSUBS 0.672419f
C606 VTAIL.n15 VSUBS 0.012226f
C607 VTAIL.n16 VSUBS 0.012945f
C608 VTAIL.n17 VSUBS 0.028898f
C609 VTAIL.n18 VSUBS 0.028898f
C610 VTAIL.n19 VSUBS 0.012945f
C611 VTAIL.n20 VSUBS 0.012226f
C612 VTAIL.n21 VSUBS 0.022752f
C613 VTAIL.n22 VSUBS 0.022752f
C614 VTAIL.n23 VSUBS 0.012226f
C615 VTAIL.n24 VSUBS 0.012945f
C616 VTAIL.n25 VSUBS 0.028898f
C617 VTAIL.n26 VSUBS 0.028898f
C618 VTAIL.n27 VSUBS 0.012945f
C619 VTAIL.n28 VSUBS 0.012226f
C620 VTAIL.n29 VSUBS 0.022752f
C621 VTAIL.n30 VSUBS 0.022752f
C622 VTAIL.n31 VSUBS 0.012226f
C623 VTAIL.n32 VSUBS 0.012945f
C624 VTAIL.n33 VSUBS 0.028898f
C625 VTAIL.n34 VSUBS 0.072592f
C626 VTAIL.n35 VSUBS 0.012945f
C627 VTAIL.n36 VSUBS 0.012226f
C628 VTAIL.n37 VSUBS 0.052902f
C629 VTAIL.n38 VSUBS 0.036632f
C630 VTAIL.n39 VSUBS 0.971745f
C631 VTAIL.n40 VSUBS 0.025773f
C632 VTAIL.n41 VSUBS 0.022752f
C633 VTAIL.n42 VSUBS 0.012226f
C634 VTAIL.n43 VSUBS 0.028898f
C635 VTAIL.n44 VSUBS 0.012945f
C636 VTAIL.n45 VSUBS 0.022752f
C637 VTAIL.n46 VSUBS 0.012226f
C638 VTAIL.n47 VSUBS 0.028898f
C639 VTAIL.n48 VSUBS 0.012945f
C640 VTAIL.n49 VSUBS 0.022752f
C641 VTAIL.n50 VSUBS 0.012226f
C642 VTAIL.n51 VSUBS 0.021674f
C643 VTAIL.n52 VSUBS 0.018382f
C644 VTAIL.t3 VSUBS 0.061707f
C645 VTAIL.n53 VSUBS 0.109981f
C646 VTAIL.n54 VSUBS 0.672419f
C647 VTAIL.n55 VSUBS 0.012226f
C648 VTAIL.n56 VSUBS 0.012945f
C649 VTAIL.n57 VSUBS 0.028898f
C650 VTAIL.n58 VSUBS 0.028898f
C651 VTAIL.n59 VSUBS 0.012945f
C652 VTAIL.n60 VSUBS 0.012226f
C653 VTAIL.n61 VSUBS 0.022752f
C654 VTAIL.n62 VSUBS 0.022752f
C655 VTAIL.n63 VSUBS 0.012226f
C656 VTAIL.n64 VSUBS 0.012945f
C657 VTAIL.n65 VSUBS 0.028898f
C658 VTAIL.n66 VSUBS 0.028898f
C659 VTAIL.n67 VSUBS 0.012945f
C660 VTAIL.n68 VSUBS 0.012226f
C661 VTAIL.n69 VSUBS 0.022752f
C662 VTAIL.n70 VSUBS 0.022752f
C663 VTAIL.n71 VSUBS 0.012226f
C664 VTAIL.n72 VSUBS 0.012945f
C665 VTAIL.n73 VSUBS 0.028898f
C666 VTAIL.n74 VSUBS 0.072592f
C667 VTAIL.n75 VSUBS 0.012945f
C668 VTAIL.n76 VSUBS 0.012226f
C669 VTAIL.n77 VSUBS 0.052902f
C670 VTAIL.n78 VSUBS 0.036632f
C671 VTAIL.n79 VSUBS 0.982173f
C672 VTAIL.n80 VSUBS 0.025773f
C673 VTAIL.n81 VSUBS 0.022752f
C674 VTAIL.n82 VSUBS 0.012226f
C675 VTAIL.n83 VSUBS 0.028898f
C676 VTAIL.n84 VSUBS 0.012945f
C677 VTAIL.n85 VSUBS 0.022752f
C678 VTAIL.n86 VSUBS 0.012226f
C679 VTAIL.n87 VSUBS 0.028898f
C680 VTAIL.n88 VSUBS 0.012945f
C681 VTAIL.n89 VSUBS 0.022752f
C682 VTAIL.n90 VSUBS 0.012226f
C683 VTAIL.n91 VSUBS 0.021674f
C684 VTAIL.n92 VSUBS 0.018382f
C685 VTAIL.t1 VSUBS 0.061707f
C686 VTAIL.n93 VSUBS 0.109981f
C687 VTAIL.n94 VSUBS 0.672419f
C688 VTAIL.n95 VSUBS 0.012226f
C689 VTAIL.n96 VSUBS 0.012945f
C690 VTAIL.n97 VSUBS 0.028898f
C691 VTAIL.n98 VSUBS 0.028898f
C692 VTAIL.n99 VSUBS 0.012945f
C693 VTAIL.n100 VSUBS 0.012226f
C694 VTAIL.n101 VSUBS 0.022752f
C695 VTAIL.n102 VSUBS 0.022752f
C696 VTAIL.n103 VSUBS 0.012226f
C697 VTAIL.n104 VSUBS 0.012945f
C698 VTAIL.n105 VSUBS 0.028898f
C699 VTAIL.n106 VSUBS 0.028898f
C700 VTAIL.n107 VSUBS 0.012945f
C701 VTAIL.n108 VSUBS 0.012226f
C702 VTAIL.n109 VSUBS 0.022752f
C703 VTAIL.n110 VSUBS 0.022752f
C704 VTAIL.n111 VSUBS 0.012226f
C705 VTAIL.n112 VSUBS 0.012945f
C706 VTAIL.n113 VSUBS 0.028898f
C707 VTAIL.n114 VSUBS 0.072592f
C708 VTAIL.n115 VSUBS 0.012945f
C709 VTAIL.n116 VSUBS 0.012226f
C710 VTAIL.n117 VSUBS 0.052902f
C711 VTAIL.n118 VSUBS 0.036632f
C712 VTAIL.n119 VSUBS 0.923396f
C713 VTAIL.n120 VSUBS 0.025773f
C714 VTAIL.n121 VSUBS 0.022752f
C715 VTAIL.n122 VSUBS 0.012226f
C716 VTAIL.n123 VSUBS 0.028898f
C717 VTAIL.n124 VSUBS 0.012945f
C718 VTAIL.n125 VSUBS 0.022752f
C719 VTAIL.n126 VSUBS 0.012226f
C720 VTAIL.n127 VSUBS 0.028898f
C721 VTAIL.n128 VSUBS 0.012945f
C722 VTAIL.n129 VSUBS 0.022752f
C723 VTAIL.n130 VSUBS 0.012226f
C724 VTAIL.n131 VSUBS 0.021674f
C725 VTAIL.n132 VSUBS 0.018382f
C726 VTAIL.t2 VSUBS 0.061707f
C727 VTAIL.n133 VSUBS 0.109981f
C728 VTAIL.n134 VSUBS 0.672419f
C729 VTAIL.n135 VSUBS 0.012226f
C730 VTAIL.n136 VSUBS 0.012945f
C731 VTAIL.n137 VSUBS 0.028898f
C732 VTAIL.n138 VSUBS 0.028898f
C733 VTAIL.n139 VSUBS 0.012945f
C734 VTAIL.n140 VSUBS 0.012226f
C735 VTAIL.n141 VSUBS 0.022752f
C736 VTAIL.n142 VSUBS 0.022752f
C737 VTAIL.n143 VSUBS 0.012226f
C738 VTAIL.n144 VSUBS 0.012945f
C739 VTAIL.n145 VSUBS 0.028898f
C740 VTAIL.n146 VSUBS 0.028898f
C741 VTAIL.n147 VSUBS 0.012945f
C742 VTAIL.n148 VSUBS 0.012226f
C743 VTAIL.n149 VSUBS 0.022752f
C744 VTAIL.n150 VSUBS 0.022752f
C745 VTAIL.n151 VSUBS 0.012226f
C746 VTAIL.n152 VSUBS 0.012945f
C747 VTAIL.n153 VSUBS 0.028898f
C748 VTAIL.n154 VSUBS 0.072592f
C749 VTAIL.n155 VSUBS 0.012945f
C750 VTAIL.n156 VSUBS 0.012226f
C751 VTAIL.n157 VSUBS 0.052902f
C752 VTAIL.n158 VSUBS 0.036632f
C753 VTAIL.n159 VSUBS 0.869991f
C754 VN.t0 VSUBS 0.528975f
C755 VN.t1 VSUBS 0.612902f
.ends

