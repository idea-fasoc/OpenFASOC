* NGSPICE file created from diff_pair_sample_0947.ext - technology: sky130A

.subckt diff_pair_sample_0947 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=1.3806 ps=7.86 w=3.54 l=2.02
X1 VTAIL.t7 VP.t1 VDD1.t4 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=0.5841 ps=3.87 w=3.54 l=2.02
X2 VDD2.t5 VN.t0 VTAIL.t4 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0.5841 ps=3.87 w=3.54 l=2.02
X3 VDD2.t4 VN.t1 VTAIL.t3 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=1.3806 ps=7.86 w=3.54 l=2.02
X4 VDD2.t3 VN.t2 VTAIL.t5 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=1.3806 ps=7.86 w=3.54 l=2.02
X5 B.t11 B.t9 B.t10 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0 ps=0 w=3.54 l=2.02
X6 B.t8 B.t6 B.t7 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0 ps=0 w=3.54 l=2.02
X7 VTAIL.t2 VN.t3 VDD2.t2 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=0.5841 ps=3.87 w=3.54 l=2.02
X8 B.t5 B.t3 B.t4 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0 ps=0 w=3.54 l=2.02
X9 VDD1.t3 VP.t2 VTAIL.t10 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=1.3806 ps=7.86 w=3.54 l=2.02
X10 VDD1.t2 VP.t3 VTAIL.t9 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0.5841 ps=3.87 w=3.54 l=2.02
X11 VTAIL.t1 VN.t4 VDD2.t1 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=0.5841 ps=3.87 w=3.54 l=2.02
X12 VDD2.t0 VN.t5 VTAIL.t0 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0.5841 ps=3.87 w=3.54 l=2.02
X13 VDD1.t1 VP.t4 VTAIL.t6 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0.5841 ps=3.87 w=3.54 l=2.02
X14 B.t2 B.t0 B.t1 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=1.3806 pd=7.86 as=0 ps=0 w=3.54 l=2.02
X15 VTAIL.t11 VP.t5 VDD1.t0 w_n2850_n1676# sky130_fd_pr__pfet_01v8 ad=0.5841 pd=3.87 as=0.5841 ps=3.87 w=3.54 l=2.02
R0 VP.n10 VP.n9 161.3
R1 VP.n11 VP.n6 161.3
R2 VP.n13 VP.n12 161.3
R3 VP.n14 VP.n5 161.3
R4 VP.n31 VP.n0 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n28 VP.n1 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n25 VP.n2 161.3
R9 VP.n24 VP.n23 161.3
R10 VP.n22 VP.n3 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n19 VP.n4 161.3
R13 VP.n18 VP.n17 93.694
R14 VP.n33 VP.n32 93.694
R15 VP.n16 VP.n15 93.694
R16 VP.n7 VP.t4 75.9506
R17 VP.n20 VP.n3 56.5617
R18 VP.n30 VP.n1 56.5617
R19 VP.n13 VP.n6 56.5617
R20 VP.n8 VP.n7 45.9066
R21 VP.n25 VP.t5 42.2352
R22 VP.n18 VP.t3 42.2352
R23 VP.n32 VP.t2 42.2352
R24 VP.n8 VP.t1 42.2352
R25 VP.n15 VP.t0 42.2352
R26 VP.n17 VP.n16 39.9807
R27 VP.n20 VP.n19 24.5923
R28 VP.n24 VP.n3 24.5923
R29 VP.n25 VP.n24 24.5923
R30 VP.n26 VP.n25 24.5923
R31 VP.n26 VP.n1 24.5923
R32 VP.n31 VP.n30 24.5923
R33 VP.n14 VP.n13 24.5923
R34 VP.n9 VP.n8 24.5923
R35 VP.n9 VP.n6 24.5923
R36 VP.n19 VP.n18 17.2148
R37 VP.n32 VP.n31 17.2148
R38 VP.n15 VP.n14 17.2148
R39 VP.n10 VP.n7 9.21706
R40 VP.n16 VP.n5 0.278335
R41 VP.n17 VP.n4 0.278335
R42 VP.n33 VP.n0 0.278335
R43 VP.n11 VP.n10 0.189894
R44 VP.n12 VP.n11 0.189894
R45 VP.n12 VP.n5 0.189894
R46 VP.n21 VP.n4 0.189894
R47 VP.n22 VP.n21 0.189894
R48 VP.n23 VP.n22 0.189894
R49 VP.n23 VP.n2 0.189894
R50 VP.n27 VP.n2 0.189894
R51 VP.n28 VP.n27 0.189894
R52 VP.n29 VP.n28 0.189894
R53 VP.n29 VP.n0 0.189894
R54 VP VP.n33 0.153485
R55 VTAIL.n7 VTAIL.t3 113.576
R56 VTAIL.n11 VTAIL.t5 113.576
R57 VTAIL.n2 VTAIL.t10 113.576
R58 VTAIL.n10 VTAIL.t8 113.576
R59 VTAIL.n9 VTAIL.n8 104.394
R60 VTAIL.n6 VTAIL.n5 104.394
R61 VTAIL.n1 VTAIL.n0 104.392
R62 VTAIL.n4 VTAIL.n3 104.392
R63 VTAIL.n6 VTAIL.n4 19.4703
R64 VTAIL.n11 VTAIL.n10 17.4445
R65 VTAIL.n0 VTAIL.t4 9.1827
R66 VTAIL.n0 VTAIL.t2 9.1827
R67 VTAIL.n3 VTAIL.t9 9.1827
R68 VTAIL.n3 VTAIL.t11 9.1827
R69 VTAIL.n8 VTAIL.t6 9.1827
R70 VTAIL.n8 VTAIL.t7 9.1827
R71 VTAIL.n5 VTAIL.t0 9.1827
R72 VTAIL.n5 VTAIL.t1 9.1827
R73 VTAIL.n7 VTAIL.n6 2.02636
R74 VTAIL.n10 VTAIL.n9 2.02636
R75 VTAIL.n4 VTAIL.n2 2.02636
R76 VTAIL.n9 VTAIL.n7 1.48326
R77 VTAIL.n2 VTAIL.n1 1.48326
R78 VTAIL VTAIL.n11 1.46171
R79 VTAIL VTAIL.n1 0.565155
R80 VDD1 VDD1.t1 131.832
R81 VDD1.n1 VDD1.t2 131.719
R82 VDD1.n1 VDD1.n0 121.522
R83 VDD1.n3 VDD1.n2 121.072
R84 VDD1.n3 VDD1.n1 34.947
R85 VDD1.n2 VDD1.t4 9.1827
R86 VDD1.n2 VDD1.t5 9.1827
R87 VDD1.n0 VDD1.t0 9.1827
R88 VDD1.n0 VDD1.t3 9.1827
R89 VDD1 VDD1.n3 0.448776
R90 VN.n21 VN.n12 161.3
R91 VN.n20 VN.n19 161.3
R92 VN.n18 VN.n13 161.3
R93 VN.n17 VN.n16 161.3
R94 VN.n9 VN.n0 161.3
R95 VN.n8 VN.n7 161.3
R96 VN.n6 VN.n1 161.3
R97 VN.n5 VN.n4 161.3
R98 VN.n11 VN.n10 93.694
R99 VN.n23 VN.n22 93.694
R100 VN.n2 VN.t0 75.9506
R101 VN.n14 VN.t1 75.9506
R102 VN.n8 VN.n1 56.5617
R103 VN.n20 VN.n13 56.5617
R104 VN.n15 VN.n14 45.9066
R105 VN.n3 VN.n2 45.9066
R106 VN.n3 VN.t3 42.2352
R107 VN.n10 VN.t2 42.2352
R108 VN.n15 VN.t4 42.2352
R109 VN.n22 VN.t5 42.2352
R110 VN VN.n23 40.2596
R111 VN.n4 VN.n3 24.5923
R112 VN.n4 VN.n1 24.5923
R113 VN.n9 VN.n8 24.5923
R114 VN.n16 VN.n13 24.5923
R115 VN.n16 VN.n15 24.5923
R116 VN.n21 VN.n20 24.5923
R117 VN.n10 VN.n9 17.2148
R118 VN.n22 VN.n21 17.2148
R119 VN.n17 VN.n14 9.21706
R120 VN.n5 VN.n2 9.21706
R121 VN.n23 VN.n12 0.278335
R122 VN.n11 VN.n0 0.278335
R123 VN.n19 VN.n12 0.189894
R124 VN.n19 VN.n18 0.189894
R125 VN.n18 VN.n17 0.189894
R126 VN.n6 VN.n5 0.189894
R127 VN.n7 VN.n6 0.189894
R128 VN.n7 VN.n0 0.189894
R129 VN VN.n11 0.153485
R130 VDD2.n1 VDD2.t5 131.719
R131 VDD2.n2 VDD2.t0 130.255
R132 VDD2.n1 VDD2.n0 121.522
R133 VDD2 VDD2.n3 121.52
R134 VDD2.n2 VDD2.n1 33.3511
R135 VDD2.n3 VDD2.t1 9.1827
R136 VDD2.n3 VDD2.t4 9.1827
R137 VDD2.n0 VDD2.t2 9.1827
R138 VDD2.n0 VDD2.t3 9.1827
R139 VDD2 VDD2.n2 1.57809
R140 B.n241 B.n240 585
R141 B.n239 B.n82 585
R142 B.n238 B.n237 585
R143 B.n236 B.n83 585
R144 B.n235 B.n234 585
R145 B.n233 B.n84 585
R146 B.n232 B.n231 585
R147 B.n230 B.n85 585
R148 B.n229 B.n228 585
R149 B.n227 B.n86 585
R150 B.n226 B.n225 585
R151 B.n224 B.n87 585
R152 B.n223 B.n222 585
R153 B.n221 B.n88 585
R154 B.n220 B.n219 585
R155 B.n218 B.n89 585
R156 B.n217 B.n216 585
R157 B.n215 B.n214 585
R158 B.n213 B.n93 585
R159 B.n212 B.n211 585
R160 B.n210 B.n94 585
R161 B.n209 B.n208 585
R162 B.n207 B.n95 585
R163 B.n206 B.n205 585
R164 B.n204 B.n96 585
R165 B.n203 B.n202 585
R166 B.n200 B.n97 585
R167 B.n199 B.n198 585
R168 B.n197 B.n100 585
R169 B.n196 B.n195 585
R170 B.n194 B.n101 585
R171 B.n193 B.n192 585
R172 B.n191 B.n102 585
R173 B.n190 B.n189 585
R174 B.n188 B.n103 585
R175 B.n187 B.n186 585
R176 B.n185 B.n104 585
R177 B.n184 B.n183 585
R178 B.n182 B.n105 585
R179 B.n181 B.n180 585
R180 B.n179 B.n106 585
R181 B.n178 B.n177 585
R182 B.n176 B.n107 585
R183 B.n242 B.n81 585
R184 B.n244 B.n243 585
R185 B.n245 B.n80 585
R186 B.n247 B.n246 585
R187 B.n248 B.n79 585
R188 B.n250 B.n249 585
R189 B.n251 B.n78 585
R190 B.n253 B.n252 585
R191 B.n254 B.n77 585
R192 B.n256 B.n255 585
R193 B.n257 B.n76 585
R194 B.n259 B.n258 585
R195 B.n260 B.n75 585
R196 B.n262 B.n261 585
R197 B.n263 B.n74 585
R198 B.n265 B.n264 585
R199 B.n266 B.n73 585
R200 B.n268 B.n267 585
R201 B.n269 B.n72 585
R202 B.n271 B.n270 585
R203 B.n272 B.n71 585
R204 B.n274 B.n273 585
R205 B.n275 B.n70 585
R206 B.n277 B.n276 585
R207 B.n278 B.n69 585
R208 B.n280 B.n279 585
R209 B.n281 B.n68 585
R210 B.n283 B.n282 585
R211 B.n284 B.n67 585
R212 B.n286 B.n285 585
R213 B.n287 B.n66 585
R214 B.n289 B.n288 585
R215 B.n290 B.n65 585
R216 B.n292 B.n291 585
R217 B.n293 B.n64 585
R218 B.n295 B.n294 585
R219 B.n296 B.n63 585
R220 B.n298 B.n297 585
R221 B.n299 B.n62 585
R222 B.n301 B.n300 585
R223 B.n302 B.n61 585
R224 B.n304 B.n303 585
R225 B.n305 B.n60 585
R226 B.n307 B.n306 585
R227 B.n308 B.n59 585
R228 B.n310 B.n309 585
R229 B.n311 B.n58 585
R230 B.n313 B.n312 585
R231 B.n314 B.n57 585
R232 B.n316 B.n315 585
R233 B.n317 B.n56 585
R234 B.n319 B.n318 585
R235 B.n320 B.n55 585
R236 B.n322 B.n321 585
R237 B.n323 B.n54 585
R238 B.n325 B.n324 585
R239 B.n326 B.n53 585
R240 B.n328 B.n327 585
R241 B.n329 B.n52 585
R242 B.n331 B.n330 585
R243 B.n332 B.n51 585
R244 B.n334 B.n333 585
R245 B.n335 B.n50 585
R246 B.n337 B.n336 585
R247 B.n338 B.n49 585
R248 B.n340 B.n339 585
R249 B.n341 B.n48 585
R250 B.n343 B.n342 585
R251 B.n344 B.n47 585
R252 B.n346 B.n345 585
R253 B.n347 B.n46 585
R254 B.n349 B.n348 585
R255 B.n415 B.n414 585
R256 B.n413 B.n20 585
R257 B.n412 B.n411 585
R258 B.n410 B.n21 585
R259 B.n409 B.n408 585
R260 B.n407 B.n22 585
R261 B.n406 B.n405 585
R262 B.n404 B.n23 585
R263 B.n403 B.n402 585
R264 B.n401 B.n24 585
R265 B.n400 B.n399 585
R266 B.n398 B.n25 585
R267 B.n397 B.n396 585
R268 B.n395 B.n26 585
R269 B.n394 B.n393 585
R270 B.n392 B.n27 585
R271 B.n391 B.n390 585
R272 B.n389 B.n388 585
R273 B.n387 B.n31 585
R274 B.n386 B.n385 585
R275 B.n384 B.n32 585
R276 B.n383 B.n382 585
R277 B.n381 B.n33 585
R278 B.n380 B.n379 585
R279 B.n378 B.n34 585
R280 B.n377 B.n376 585
R281 B.n374 B.n35 585
R282 B.n373 B.n372 585
R283 B.n371 B.n38 585
R284 B.n370 B.n369 585
R285 B.n368 B.n39 585
R286 B.n367 B.n366 585
R287 B.n365 B.n40 585
R288 B.n364 B.n363 585
R289 B.n362 B.n41 585
R290 B.n361 B.n360 585
R291 B.n359 B.n42 585
R292 B.n358 B.n357 585
R293 B.n356 B.n43 585
R294 B.n355 B.n354 585
R295 B.n353 B.n44 585
R296 B.n352 B.n351 585
R297 B.n350 B.n45 585
R298 B.n416 B.n19 585
R299 B.n418 B.n417 585
R300 B.n419 B.n18 585
R301 B.n421 B.n420 585
R302 B.n422 B.n17 585
R303 B.n424 B.n423 585
R304 B.n425 B.n16 585
R305 B.n427 B.n426 585
R306 B.n428 B.n15 585
R307 B.n430 B.n429 585
R308 B.n431 B.n14 585
R309 B.n433 B.n432 585
R310 B.n434 B.n13 585
R311 B.n436 B.n435 585
R312 B.n437 B.n12 585
R313 B.n439 B.n438 585
R314 B.n440 B.n11 585
R315 B.n442 B.n441 585
R316 B.n443 B.n10 585
R317 B.n445 B.n444 585
R318 B.n446 B.n9 585
R319 B.n448 B.n447 585
R320 B.n449 B.n8 585
R321 B.n451 B.n450 585
R322 B.n452 B.n7 585
R323 B.n454 B.n453 585
R324 B.n455 B.n6 585
R325 B.n457 B.n456 585
R326 B.n458 B.n5 585
R327 B.n460 B.n459 585
R328 B.n461 B.n4 585
R329 B.n463 B.n462 585
R330 B.n464 B.n3 585
R331 B.n466 B.n465 585
R332 B.n467 B.n0 585
R333 B.n2 B.n1 585
R334 B.n125 B.n124 585
R335 B.n127 B.n126 585
R336 B.n128 B.n123 585
R337 B.n130 B.n129 585
R338 B.n131 B.n122 585
R339 B.n133 B.n132 585
R340 B.n134 B.n121 585
R341 B.n136 B.n135 585
R342 B.n137 B.n120 585
R343 B.n139 B.n138 585
R344 B.n140 B.n119 585
R345 B.n142 B.n141 585
R346 B.n143 B.n118 585
R347 B.n145 B.n144 585
R348 B.n146 B.n117 585
R349 B.n148 B.n147 585
R350 B.n149 B.n116 585
R351 B.n151 B.n150 585
R352 B.n152 B.n115 585
R353 B.n154 B.n153 585
R354 B.n155 B.n114 585
R355 B.n157 B.n156 585
R356 B.n158 B.n113 585
R357 B.n160 B.n159 585
R358 B.n161 B.n112 585
R359 B.n163 B.n162 585
R360 B.n164 B.n111 585
R361 B.n166 B.n165 585
R362 B.n167 B.n110 585
R363 B.n169 B.n168 585
R364 B.n170 B.n109 585
R365 B.n172 B.n171 585
R366 B.n173 B.n108 585
R367 B.n175 B.n174 585
R368 B.n174 B.n107 545.355
R369 B.n240 B.n81 545.355
R370 B.n348 B.n45 545.355
R371 B.n414 B.n19 545.355
R372 B.n469 B.n468 256.663
R373 B.n98 B.t9 249.2
R374 B.n90 B.t3 249.2
R375 B.n36 B.t0 249.2
R376 B.n28 B.t6 249.2
R377 B.n468 B.n467 235.042
R378 B.n468 B.n2 235.042
R379 B.n90 B.t4 174.542
R380 B.n36 B.t2 174.542
R381 B.n98 B.t10 174.54
R382 B.n28 B.t8 174.54
R383 B.n178 B.n107 163.367
R384 B.n179 B.n178 163.367
R385 B.n180 B.n179 163.367
R386 B.n180 B.n105 163.367
R387 B.n184 B.n105 163.367
R388 B.n185 B.n184 163.367
R389 B.n186 B.n185 163.367
R390 B.n186 B.n103 163.367
R391 B.n190 B.n103 163.367
R392 B.n191 B.n190 163.367
R393 B.n192 B.n191 163.367
R394 B.n192 B.n101 163.367
R395 B.n196 B.n101 163.367
R396 B.n197 B.n196 163.367
R397 B.n198 B.n197 163.367
R398 B.n198 B.n97 163.367
R399 B.n203 B.n97 163.367
R400 B.n204 B.n203 163.367
R401 B.n205 B.n204 163.367
R402 B.n205 B.n95 163.367
R403 B.n209 B.n95 163.367
R404 B.n210 B.n209 163.367
R405 B.n211 B.n210 163.367
R406 B.n211 B.n93 163.367
R407 B.n215 B.n93 163.367
R408 B.n216 B.n215 163.367
R409 B.n216 B.n89 163.367
R410 B.n220 B.n89 163.367
R411 B.n221 B.n220 163.367
R412 B.n222 B.n221 163.367
R413 B.n222 B.n87 163.367
R414 B.n226 B.n87 163.367
R415 B.n227 B.n226 163.367
R416 B.n228 B.n227 163.367
R417 B.n228 B.n85 163.367
R418 B.n232 B.n85 163.367
R419 B.n233 B.n232 163.367
R420 B.n234 B.n233 163.367
R421 B.n234 B.n83 163.367
R422 B.n238 B.n83 163.367
R423 B.n239 B.n238 163.367
R424 B.n240 B.n239 163.367
R425 B.n348 B.n347 163.367
R426 B.n347 B.n346 163.367
R427 B.n346 B.n47 163.367
R428 B.n342 B.n47 163.367
R429 B.n342 B.n341 163.367
R430 B.n341 B.n340 163.367
R431 B.n340 B.n49 163.367
R432 B.n336 B.n49 163.367
R433 B.n336 B.n335 163.367
R434 B.n335 B.n334 163.367
R435 B.n334 B.n51 163.367
R436 B.n330 B.n51 163.367
R437 B.n330 B.n329 163.367
R438 B.n329 B.n328 163.367
R439 B.n328 B.n53 163.367
R440 B.n324 B.n53 163.367
R441 B.n324 B.n323 163.367
R442 B.n323 B.n322 163.367
R443 B.n322 B.n55 163.367
R444 B.n318 B.n55 163.367
R445 B.n318 B.n317 163.367
R446 B.n317 B.n316 163.367
R447 B.n316 B.n57 163.367
R448 B.n312 B.n57 163.367
R449 B.n312 B.n311 163.367
R450 B.n311 B.n310 163.367
R451 B.n310 B.n59 163.367
R452 B.n306 B.n59 163.367
R453 B.n306 B.n305 163.367
R454 B.n305 B.n304 163.367
R455 B.n304 B.n61 163.367
R456 B.n300 B.n61 163.367
R457 B.n300 B.n299 163.367
R458 B.n299 B.n298 163.367
R459 B.n298 B.n63 163.367
R460 B.n294 B.n63 163.367
R461 B.n294 B.n293 163.367
R462 B.n293 B.n292 163.367
R463 B.n292 B.n65 163.367
R464 B.n288 B.n65 163.367
R465 B.n288 B.n287 163.367
R466 B.n287 B.n286 163.367
R467 B.n286 B.n67 163.367
R468 B.n282 B.n67 163.367
R469 B.n282 B.n281 163.367
R470 B.n281 B.n280 163.367
R471 B.n280 B.n69 163.367
R472 B.n276 B.n69 163.367
R473 B.n276 B.n275 163.367
R474 B.n275 B.n274 163.367
R475 B.n274 B.n71 163.367
R476 B.n270 B.n71 163.367
R477 B.n270 B.n269 163.367
R478 B.n269 B.n268 163.367
R479 B.n268 B.n73 163.367
R480 B.n264 B.n73 163.367
R481 B.n264 B.n263 163.367
R482 B.n263 B.n262 163.367
R483 B.n262 B.n75 163.367
R484 B.n258 B.n75 163.367
R485 B.n258 B.n257 163.367
R486 B.n257 B.n256 163.367
R487 B.n256 B.n77 163.367
R488 B.n252 B.n77 163.367
R489 B.n252 B.n251 163.367
R490 B.n251 B.n250 163.367
R491 B.n250 B.n79 163.367
R492 B.n246 B.n79 163.367
R493 B.n246 B.n245 163.367
R494 B.n245 B.n244 163.367
R495 B.n244 B.n81 163.367
R496 B.n414 B.n413 163.367
R497 B.n413 B.n412 163.367
R498 B.n412 B.n21 163.367
R499 B.n408 B.n21 163.367
R500 B.n408 B.n407 163.367
R501 B.n407 B.n406 163.367
R502 B.n406 B.n23 163.367
R503 B.n402 B.n23 163.367
R504 B.n402 B.n401 163.367
R505 B.n401 B.n400 163.367
R506 B.n400 B.n25 163.367
R507 B.n396 B.n25 163.367
R508 B.n396 B.n395 163.367
R509 B.n395 B.n394 163.367
R510 B.n394 B.n27 163.367
R511 B.n390 B.n27 163.367
R512 B.n390 B.n389 163.367
R513 B.n389 B.n31 163.367
R514 B.n385 B.n31 163.367
R515 B.n385 B.n384 163.367
R516 B.n384 B.n383 163.367
R517 B.n383 B.n33 163.367
R518 B.n379 B.n33 163.367
R519 B.n379 B.n378 163.367
R520 B.n378 B.n377 163.367
R521 B.n377 B.n35 163.367
R522 B.n372 B.n35 163.367
R523 B.n372 B.n371 163.367
R524 B.n371 B.n370 163.367
R525 B.n370 B.n39 163.367
R526 B.n366 B.n39 163.367
R527 B.n366 B.n365 163.367
R528 B.n365 B.n364 163.367
R529 B.n364 B.n41 163.367
R530 B.n360 B.n41 163.367
R531 B.n360 B.n359 163.367
R532 B.n359 B.n358 163.367
R533 B.n358 B.n43 163.367
R534 B.n354 B.n43 163.367
R535 B.n354 B.n353 163.367
R536 B.n353 B.n352 163.367
R537 B.n352 B.n45 163.367
R538 B.n418 B.n19 163.367
R539 B.n419 B.n418 163.367
R540 B.n420 B.n419 163.367
R541 B.n420 B.n17 163.367
R542 B.n424 B.n17 163.367
R543 B.n425 B.n424 163.367
R544 B.n426 B.n425 163.367
R545 B.n426 B.n15 163.367
R546 B.n430 B.n15 163.367
R547 B.n431 B.n430 163.367
R548 B.n432 B.n431 163.367
R549 B.n432 B.n13 163.367
R550 B.n436 B.n13 163.367
R551 B.n437 B.n436 163.367
R552 B.n438 B.n437 163.367
R553 B.n438 B.n11 163.367
R554 B.n442 B.n11 163.367
R555 B.n443 B.n442 163.367
R556 B.n444 B.n443 163.367
R557 B.n444 B.n9 163.367
R558 B.n448 B.n9 163.367
R559 B.n449 B.n448 163.367
R560 B.n450 B.n449 163.367
R561 B.n450 B.n7 163.367
R562 B.n454 B.n7 163.367
R563 B.n455 B.n454 163.367
R564 B.n456 B.n455 163.367
R565 B.n456 B.n5 163.367
R566 B.n460 B.n5 163.367
R567 B.n461 B.n460 163.367
R568 B.n462 B.n461 163.367
R569 B.n462 B.n3 163.367
R570 B.n466 B.n3 163.367
R571 B.n467 B.n466 163.367
R572 B.n125 B.n2 163.367
R573 B.n126 B.n125 163.367
R574 B.n126 B.n123 163.367
R575 B.n130 B.n123 163.367
R576 B.n131 B.n130 163.367
R577 B.n132 B.n131 163.367
R578 B.n132 B.n121 163.367
R579 B.n136 B.n121 163.367
R580 B.n137 B.n136 163.367
R581 B.n138 B.n137 163.367
R582 B.n138 B.n119 163.367
R583 B.n142 B.n119 163.367
R584 B.n143 B.n142 163.367
R585 B.n144 B.n143 163.367
R586 B.n144 B.n117 163.367
R587 B.n148 B.n117 163.367
R588 B.n149 B.n148 163.367
R589 B.n150 B.n149 163.367
R590 B.n150 B.n115 163.367
R591 B.n154 B.n115 163.367
R592 B.n155 B.n154 163.367
R593 B.n156 B.n155 163.367
R594 B.n156 B.n113 163.367
R595 B.n160 B.n113 163.367
R596 B.n161 B.n160 163.367
R597 B.n162 B.n161 163.367
R598 B.n162 B.n111 163.367
R599 B.n166 B.n111 163.367
R600 B.n167 B.n166 163.367
R601 B.n168 B.n167 163.367
R602 B.n168 B.n109 163.367
R603 B.n172 B.n109 163.367
R604 B.n173 B.n172 163.367
R605 B.n174 B.n173 163.367
R606 B.n91 B.t5 128.965
R607 B.n37 B.t1 128.965
R608 B.n99 B.t11 128.964
R609 B.n29 B.t7 128.964
R610 B.n201 B.n99 59.5399
R611 B.n92 B.n91 59.5399
R612 B.n375 B.n37 59.5399
R613 B.n30 B.n29 59.5399
R614 B.n99 B.n98 45.5763
R615 B.n91 B.n90 45.5763
R616 B.n37 B.n36 45.5763
R617 B.n29 B.n28 45.5763
R618 B.n416 B.n415 35.4346
R619 B.n350 B.n349 35.4346
R620 B.n242 B.n241 35.4346
R621 B.n176 B.n175 35.4346
R622 B B.n469 18.0485
R623 B.n417 B.n416 10.6151
R624 B.n417 B.n18 10.6151
R625 B.n421 B.n18 10.6151
R626 B.n422 B.n421 10.6151
R627 B.n423 B.n422 10.6151
R628 B.n423 B.n16 10.6151
R629 B.n427 B.n16 10.6151
R630 B.n428 B.n427 10.6151
R631 B.n429 B.n428 10.6151
R632 B.n429 B.n14 10.6151
R633 B.n433 B.n14 10.6151
R634 B.n434 B.n433 10.6151
R635 B.n435 B.n434 10.6151
R636 B.n435 B.n12 10.6151
R637 B.n439 B.n12 10.6151
R638 B.n440 B.n439 10.6151
R639 B.n441 B.n440 10.6151
R640 B.n441 B.n10 10.6151
R641 B.n445 B.n10 10.6151
R642 B.n446 B.n445 10.6151
R643 B.n447 B.n446 10.6151
R644 B.n447 B.n8 10.6151
R645 B.n451 B.n8 10.6151
R646 B.n452 B.n451 10.6151
R647 B.n453 B.n452 10.6151
R648 B.n453 B.n6 10.6151
R649 B.n457 B.n6 10.6151
R650 B.n458 B.n457 10.6151
R651 B.n459 B.n458 10.6151
R652 B.n459 B.n4 10.6151
R653 B.n463 B.n4 10.6151
R654 B.n464 B.n463 10.6151
R655 B.n465 B.n464 10.6151
R656 B.n465 B.n0 10.6151
R657 B.n415 B.n20 10.6151
R658 B.n411 B.n20 10.6151
R659 B.n411 B.n410 10.6151
R660 B.n410 B.n409 10.6151
R661 B.n409 B.n22 10.6151
R662 B.n405 B.n22 10.6151
R663 B.n405 B.n404 10.6151
R664 B.n404 B.n403 10.6151
R665 B.n403 B.n24 10.6151
R666 B.n399 B.n24 10.6151
R667 B.n399 B.n398 10.6151
R668 B.n398 B.n397 10.6151
R669 B.n397 B.n26 10.6151
R670 B.n393 B.n26 10.6151
R671 B.n393 B.n392 10.6151
R672 B.n392 B.n391 10.6151
R673 B.n388 B.n387 10.6151
R674 B.n387 B.n386 10.6151
R675 B.n386 B.n32 10.6151
R676 B.n382 B.n32 10.6151
R677 B.n382 B.n381 10.6151
R678 B.n381 B.n380 10.6151
R679 B.n380 B.n34 10.6151
R680 B.n376 B.n34 10.6151
R681 B.n374 B.n373 10.6151
R682 B.n373 B.n38 10.6151
R683 B.n369 B.n38 10.6151
R684 B.n369 B.n368 10.6151
R685 B.n368 B.n367 10.6151
R686 B.n367 B.n40 10.6151
R687 B.n363 B.n40 10.6151
R688 B.n363 B.n362 10.6151
R689 B.n362 B.n361 10.6151
R690 B.n361 B.n42 10.6151
R691 B.n357 B.n42 10.6151
R692 B.n357 B.n356 10.6151
R693 B.n356 B.n355 10.6151
R694 B.n355 B.n44 10.6151
R695 B.n351 B.n44 10.6151
R696 B.n351 B.n350 10.6151
R697 B.n349 B.n46 10.6151
R698 B.n345 B.n46 10.6151
R699 B.n345 B.n344 10.6151
R700 B.n344 B.n343 10.6151
R701 B.n343 B.n48 10.6151
R702 B.n339 B.n48 10.6151
R703 B.n339 B.n338 10.6151
R704 B.n338 B.n337 10.6151
R705 B.n337 B.n50 10.6151
R706 B.n333 B.n50 10.6151
R707 B.n333 B.n332 10.6151
R708 B.n332 B.n331 10.6151
R709 B.n331 B.n52 10.6151
R710 B.n327 B.n52 10.6151
R711 B.n327 B.n326 10.6151
R712 B.n326 B.n325 10.6151
R713 B.n325 B.n54 10.6151
R714 B.n321 B.n54 10.6151
R715 B.n321 B.n320 10.6151
R716 B.n320 B.n319 10.6151
R717 B.n319 B.n56 10.6151
R718 B.n315 B.n56 10.6151
R719 B.n315 B.n314 10.6151
R720 B.n314 B.n313 10.6151
R721 B.n313 B.n58 10.6151
R722 B.n309 B.n58 10.6151
R723 B.n309 B.n308 10.6151
R724 B.n308 B.n307 10.6151
R725 B.n307 B.n60 10.6151
R726 B.n303 B.n60 10.6151
R727 B.n303 B.n302 10.6151
R728 B.n302 B.n301 10.6151
R729 B.n301 B.n62 10.6151
R730 B.n297 B.n62 10.6151
R731 B.n297 B.n296 10.6151
R732 B.n296 B.n295 10.6151
R733 B.n295 B.n64 10.6151
R734 B.n291 B.n64 10.6151
R735 B.n291 B.n290 10.6151
R736 B.n290 B.n289 10.6151
R737 B.n289 B.n66 10.6151
R738 B.n285 B.n66 10.6151
R739 B.n285 B.n284 10.6151
R740 B.n284 B.n283 10.6151
R741 B.n283 B.n68 10.6151
R742 B.n279 B.n68 10.6151
R743 B.n279 B.n278 10.6151
R744 B.n278 B.n277 10.6151
R745 B.n277 B.n70 10.6151
R746 B.n273 B.n70 10.6151
R747 B.n273 B.n272 10.6151
R748 B.n272 B.n271 10.6151
R749 B.n271 B.n72 10.6151
R750 B.n267 B.n72 10.6151
R751 B.n267 B.n266 10.6151
R752 B.n266 B.n265 10.6151
R753 B.n265 B.n74 10.6151
R754 B.n261 B.n74 10.6151
R755 B.n261 B.n260 10.6151
R756 B.n260 B.n259 10.6151
R757 B.n259 B.n76 10.6151
R758 B.n255 B.n76 10.6151
R759 B.n255 B.n254 10.6151
R760 B.n254 B.n253 10.6151
R761 B.n253 B.n78 10.6151
R762 B.n249 B.n78 10.6151
R763 B.n249 B.n248 10.6151
R764 B.n248 B.n247 10.6151
R765 B.n247 B.n80 10.6151
R766 B.n243 B.n80 10.6151
R767 B.n243 B.n242 10.6151
R768 B.n124 B.n1 10.6151
R769 B.n127 B.n124 10.6151
R770 B.n128 B.n127 10.6151
R771 B.n129 B.n128 10.6151
R772 B.n129 B.n122 10.6151
R773 B.n133 B.n122 10.6151
R774 B.n134 B.n133 10.6151
R775 B.n135 B.n134 10.6151
R776 B.n135 B.n120 10.6151
R777 B.n139 B.n120 10.6151
R778 B.n140 B.n139 10.6151
R779 B.n141 B.n140 10.6151
R780 B.n141 B.n118 10.6151
R781 B.n145 B.n118 10.6151
R782 B.n146 B.n145 10.6151
R783 B.n147 B.n146 10.6151
R784 B.n147 B.n116 10.6151
R785 B.n151 B.n116 10.6151
R786 B.n152 B.n151 10.6151
R787 B.n153 B.n152 10.6151
R788 B.n153 B.n114 10.6151
R789 B.n157 B.n114 10.6151
R790 B.n158 B.n157 10.6151
R791 B.n159 B.n158 10.6151
R792 B.n159 B.n112 10.6151
R793 B.n163 B.n112 10.6151
R794 B.n164 B.n163 10.6151
R795 B.n165 B.n164 10.6151
R796 B.n165 B.n110 10.6151
R797 B.n169 B.n110 10.6151
R798 B.n170 B.n169 10.6151
R799 B.n171 B.n170 10.6151
R800 B.n171 B.n108 10.6151
R801 B.n175 B.n108 10.6151
R802 B.n177 B.n176 10.6151
R803 B.n177 B.n106 10.6151
R804 B.n181 B.n106 10.6151
R805 B.n182 B.n181 10.6151
R806 B.n183 B.n182 10.6151
R807 B.n183 B.n104 10.6151
R808 B.n187 B.n104 10.6151
R809 B.n188 B.n187 10.6151
R810 B.n189 B.n188 10.6151
R811 B.n189 B.n102 10.6151
R812 B.n193 B.n102 10.6151
R813 B.n194 B.n193 10.6151
R814 B.n195 B.n194 10.6151
R815 B.n195 B.n100 10.6151
R816 B.n199 B.n100 10.6151
R817 B.n200 B.n199 10.6151
R818 B.n202 B.n96 10.6151
R819 B.n206 B.n96 10.6151
R820 B.n207 B.n206 10.6151
R821 B.n208 B.n207 10.6151
R822 B.n208 B.n94 10.6151
R823 B.n212 B.n94 10.6151
R824 B.n213 B.n212 10.6151
R825 B.n214 B.n213 10.6151
R826 B.n218 B.n217 10.6151
R827 B.n219 B.n218 10.6151
R828 B.n219 B.n88 10.6151
R829 B.n223 B.n88 10.6151
R830 B.n224 B.n223 10.6151
R831 B.n225 B.n224 10.6151
R832 B.n225 B.n86 10.6151
R833 B.n229 B.n86 10.6151
R834 B.n230 B.n229 10.6151
R835 B.n231 B.n230 10.6151
R836 B.n231 B.n84 10.6151
R837 B.n235 B.n84 10.6151
R838 B.n236 B.n235 10.6151
R839 B.n237 B.n236 10.6151
R840 B.n237 B.n82 10.6151
R841 B.n241 B.n82 10.6151
R842 B.n469 B.n0 8.11757
R843 B.n469 B.n1 8.11757
R844 B.n388 B.n30 6.5566
R845 B.n376 B.n375 6.5566
R846 B.n202 B.n201 6.5566
R847 B.n214 B.n92 6.5566
R848 B.n391 B.n30 4.05904
R849 B.n375 B.n374 4.05904
R850 B.n201 B.n200 4.05904
R851 B.n217 B.n92 4.05904
C0 VDD2 VTAIL 4.38042f
C1 B VDD1 1.28023f
C2 VP B 1.56583f
C3 B w_n2850_n1676# 6.51606f
C4 VDD2 VN 2.14246f
C5 VTAIL VN 2.67871f
C6 VDD2 VDD1 1.1893f
C7 VTAIL VDD1 4.33174f
C8 VP VDD2 0.41397f
C9 VP VTAIL 2.69289f
C10 VDD2 w_n2850_n1676# 1.62059f
C11 w_n2850_n1676# VTAIL 1.70444f
C12 VDD1 VN 0.154979f
C13 VP VN 4.80127f
C14 VP VDD1 2.3992f
C15 w_n2850_n1676# VN 5.098721f
C16 w_n2850_n1676# VDD1 1.55443f
C17 VP w_n2850_n1676# 5.46405f
C18 VDD2 B 1.34056f
C19 B VTAIL 1.59482f
C20 B VN 0.956548f
C21 VDD2 VSUBS 1.182884f
C22 VDD1 VSUBS 1.587059f
C23 VTAIL VSUBS 0.506811f
C24 VN VSUBS 5.02248f
C25 VP VSUBS 2.003238f
C26 B VSUBS 3.160277f
C27 w_n2850_n1676# VSUBS 60.294605f
C28 B.n0 VSUBS 0.006495f
C29 B.n1 VSUBS 0.006495f
C30 B.n2 VSUBS 0.009606f
C31 B.n3 VSUBS 0.007361f
C32 B.n4 VSUBS 0.007361f
C33 B.n5 VSUBS 0.007361f
C34 B.n6 VSUBS 0.007361f
C35 B.n7 VSUBS 0.007361f
C36 B.n8 VSUBS 0.007361f
C37 B.n9 VSUBS 0.007361f
C38 B.n10 VSUBS 0.007361f
C39 B.n11 VSUBS 0.007361f
C40 B.n12 VSUBS 0.007361f
C41 B.n13 VSUBS 0.007361f
C42 B.n14 VSUBS 0.007361f
C43 B.n15 VSUBS 0.007361f
C44 B.n16 VSUBS 0.007361f
C45 B.n17 VSUBS 0.007361f
C46 B.n18 VSUBS 0.007361f
C47 B.n19 VSUBS 0.017649f
C48 B.n20 VSUBS 0.007361f
C49 B.n21 VSUBS 0.007361f
C50 B.n22 VSUBS 0.007361f
C51 B.n23 VSUBS 0.007361f
C52 B.n24 VSUBS 0.007361f
C53 B.n25 VSUBS 0.007361f
C54 B.n26 VSUBS 0.007361f
C55 B.n27 VSUBS 0.007361f
C56 B.t7 VSUBS 0.094314f
C57 B.t8 VSUBS 0.109394f
C58 B.t6 VSUBS 0.360214f
C59 B.n28 VSUBS 0.086298f
C60 B.n29 VSUBS 0.06825f
C61 B.n30 VSUBS 0.017055f
C62 B.n31 VSUBS 0.007361f
C63 B.n32 VSUBS 0.007361f
C64 B.n33 VSUBS 0.007361f
C65 B.n34 VSUBS 0.007361f
C66 B.n35 VSUBS 0.007361f
C67 B.t1 VSUBS 0.094314f
C68 B.t2 VSUBS 0.109394f
C69 B.t0 VSUBS 0.360214f
C70 B.n36 VSUBS 0.086298f
C71 B.n37 VSUBS 0.06825f
C72 B.n38 VSUBS 0.007361f
C73 B.n39 VSUBS 0.007361f
C74 B.n40 VSUBS 0.007361f
C75 B.n41 VSUBS 0.007361f
C76 B.n42 VSUBS 0.007361f
C77 B.n43 VSUBS 0.007361f
C78 B.n44 VSUBS 0.007361f
C79 B.n45 VSUBS 0.018725f
C80 B.n46 VSUBS 0.007361f
C81 B.n47 VSUBS 0.007361f
C82 B.n48 VSUBS 0.007361f
C83 B.n49 VSUBS 0.007361f
C84 B.n50 VSUBS 0.007361f
C85 B.n51 VSUBS 0.007361f
C86 B.n52 VSUBS 0.007361f
C87 B.n53 VSUBS 0.007361f
C88 B.n54 VSUBS 0.007361f
C89 B.n55 VSUBS 0.007361f
C90 B.n56 VSUBS 0.007361f
C91 B.n57 VSUBS 0.007361f
C92 B.n58 VSUBS 0.007361f
C93 B.n59 VSUBS 0.007361f
C94 B.n60 VSUBS 0.007361f
C95 B.n61 VSUBS 0.007361f
C96 B.n62 VSUBS 0.007361f
C97 B.n63 VSUBS 0.007361f
C98 B.n64 VSUBS 0.007361f
C99 B.n65 VSUBS 0.007361f
C100 B.n66 VSUBS 0.007361f
C101 B.n67 VSUBS 0.007361f
C102 B.n68 VSUBS 0.007361f
C103 B.n69 VSUBS 0.007361f
C104 B.n70 VSUBS 0.007361f
C105 B.n71 VSUBS 0.007361f
C106 B.n72 VSUBS 0.007361f
C107 B.n73 VSUBS 0.007361f
C108 B.n74 VSUBS 0.007361f
C109 B.n75 VSUBS 0.007361f
C110 B.n76 VSUBS 0.007361f
C111 B.n77 VSUBS 0.007361f
C112 B.n78 VSUBS 0.007361f
C113 B.n79 VSUBS 0.007361f
C114 B.n80 VSUBS 0.007361f
C115 B.n81 VSUBS 0.017649f
C116 B.n82 VSUBS 0.007361f
C117 B.n83 VSUBS 0.007361f
C118 B.n84 VSUBS 0.007361f
C119 B.n85 VSUBS 0.007361f
C120 B.n86 VSUBS 0.007361f
C121 B.n87 VSUBS 0.007361f
C122 B.n88 VSUBS 0.007361f
C123 B.n89 VSUBS 0.007361f
C124 B.t5 VSUBS 0.094314f
C125 B.t4 VSUBS 0.109394f
C126 B.t3 VSUBS 0.360214f
C127 B.n90 VSUBS 0.086298f
C128 B.n91 VSUBS 0.06825f
C129 B.n92 VSUBS 0.017055f
C130 B.n93 VSUBS 0.007361f
C131 B.n94 VSUBS 0.007361f
C132 B.n95 VSUBS 0.007361f
C133 B.n96 VSUBS 0.007361f
C134 B.n97 VSUBS 0.007361f
C135 B.t11 VSUBS 0.094314f
C136 B.t10 VSUBS 0.109394f
C137 B.t9 VSUBS 0.360214f
C138 B.n98 VSUBS 0.086298f
C139 B.n99 VSUBS 0.06825f
C140 B.n100 VSUBS 0.007361f
C141 B.n101 VSUBS 0.007361f
C142 B.n102 VSUBS 0.007361f
C143 B.n103 VSUBS 0.007361f
C144 B.n104 VSUBS 0.007361f
C145 B.n105 VSUBS 0.007361f
C146 B.n106 VSUBS 0.007361f
C147 B.n107 VSUBS 0.018725f
C148 B.n108 VSUBS 0.007361f
C149 B.n109 VSUBS 0.007361f
C150 B.n110 VSUBS 0.007361f
C151 B.n111 VSUBS 0.007361f
C152 B.n112 VSUBS 0.007361f
C153 B.n113 VSUBS 0.007361f
C154 B.n114 VSUBS 0.007361f
C155 B.n115 VSUBS 0.007361f
C156 B.n116 VSUBS 0.007361f
C157 B.n117 VSUBS 0.007361f
C158 B.n118 VSUBS 0.007361f
C159 B.n119 VSUBS 0.007361f
C160 B.n120 VSUBS 0.007361f
C161 B.n121 VSUBS 0.007361f
C162 B.n122 VSUBS 0.007361f
C163 B.n123 VSUBS 0.007361f
C164 B.n124 VSUBS 0.007361f
C165 B.n125 VSUBS 0.007361f
C166 B.n126 VSUBS 0.007361f
C167 B.n127 VSUBS 0.007361f
C168 B.n128 VSUBS 0.007361f
C169 B.n129 VSUBS 0.007361f
C170 B.n130 VSUBS 0.007361f
C171 B.n131 VSUBS 0.007361f
C172 B.n132 VSUBS 0.007361f
C173 B.n133 VSUBS 0.007361f
C174 B.n134 VSUBS 0.007361f
C175 B.n135 VSUBS 0.007361f
C176 B.n136 VSUBS 0.007361f
C177 B.n137 VSUBS 0.007361f
C178 B.n138 VSUBS 0.007361f
C179 B.n139 VSUBS 0.007361f
C180 B.n140 VSUBS 0.007361f
C181 B.n141 VSUBS 0.007361f
C182 B.n142 VSUBS 0.007361f
C183 B.n143 VSUBS 0.007361f
C184 B.n144 VSUBS 0.007361f
C185 B.n145 VSUBS 0.007361f
C186 B.n146 VSUBS 0.007361f
C187 B.n147 VSUBS 0.007361f
C188 B.n148 VSUBS 0.007361f
C189 B.n149 VSUBS 0.007361f
C190 B.n150 VSUBS 0.007361f
C191 B.n151 VSUBS 0.007361f
C192 B.n152 VSUBS 0.007361f
C193 B.n153 VSUBS 0.007361f
C194 B.n154 VSUBS 0.007361f
C195 B.n155 VSUBS 0.007361f
C196 B.n156 VSUBS 0.007361f
C197 B.n157 VSUBS 0.007361f
C198 B.n158 VSUBS 0.007361f
C199 B.n159 VSUBS 0.007361f
C200 B.n160 VSUBS 0.007361f
C201 B.n161 VSUBS 0.007361f
C202 B.n162 VSUBS 0.007361f
C203 B.n163 VSUBS 0.007361f
C204 B.n164 VSUBS 0.007361f
C205 B.n165 VSUBS 0.007361f
C206 B.n166 VSUBS 0.007361f
C207 B.n167 VSUBS 0.007361f
C208 B.n168 VSUBS 0.007361f
C209 B.n169 VSUBS 0.007361f
C210 B.n170 VSUBS 0.007361f
C211 B.n171 VSUBS 0.007361f
C212 B.n172 VSUBS 0.007361f
C213 B.n173 VSUBS 0.007361f
C214 B.n174 VSUBS 0.017649f
C215 B.n175 VSUBS 0.017649f
C216 B.n176 VSUBS 0.018725f
C217 B.n177 VSUBS 0.007361f
C218 B.n178 VSUBS 0.007361f
C219 B.n179 VSUBS 0.007361f
C220 B.n180 VSUBS 0.007361f
C221 B.n181 VSUBS 0.007361f
C222 B.n182 VSUBS 0.007361f
C223 B.n183 VSUBS 0.007361f
C224 B.n184 VSUBS 0.007361f
C225 B.n185 VSUBS 0.007361f
C226 B.n186 VSUBS 0.007361f
C227 B.n187 VSUBS 0.007361f
C228 B.n188 VSUBS 0.007361f
C229 B.n189 VSUBS 0.007361f
C230 B.n190 VSUBS 0.007361f
C231 B.n191 VSUBS 0.007361f
C232 B.n192 VSUBS 0.007361f
C233 B.n193 VSUBS 0.007361f
C234 B.n194 VSUBS 0.007361f
C235 B.n195 VSUBS 0.007361f
C236 B.n196 VSUBS 0.007361f
C237 B.n197 VSUBS 0.007361f
C238 B.n198 VSUBS 0.007361f
C239 B.n199 VSUBS 0.007361f
C240 B.n200 VSUBS 0.005088f
C241 B.n201 VSUBS 0.017055f
C242 B.n202 VSUBS 0.005954f
C243 B.n203 VSUBS 0.007361f
C244 B.n204 VSUBS 0.007361f
C245 B.n205 VSUBS 0.007361f
C246 B.n206 VSUBS 0.007361f
C247 B.n207 VSUBS 0.007361f
C248 B.n208 VSUBS 0.007361f
C249 B.n209 VSUBS 0.007361f
C250 B.n210 VSUBS 0.007361f
C251 B.n211 VSUBS 0.007361f
C252 B.n212 VSUBS 0.007361f
C253 B.n213 VSUBS 0.007361f
C254 B.n214 VSUBS 0.005954f
C255 B.n215 VSUBS 0.007361f
C256 B.n216 VSUBS 0.007361f
C257 B.n217 VSUBS 0.005088f
C258 B.n218 VSUBS 0.007361f
C259 B.n219 VSUBS 0.007361f
C260 B.n220 VSUBS 0.007361f
C261 B.n221 VSUBS 0.007361f
C262 B.n222 VSUBS 0.007361f
C263 B.n223 VSUBS 0.007361f
C264 B.n224 VSUBS 0.007361f
C265 B.n225 VSUBS 0.007361f
C266 B.n226 VSUBS 0.007361f
C267 B.n227 VSUBS 0.007361f
C268 B.n228 VSUBS 0.007361f
C269 B.n229 VSUBS 0.007361f
C270 B.n230 VSUBS 0.007361f
C271 B.n231 VSUBS 0.007361f
C272 B.n232 VSUBS 0.007361f
C273 B.n233 VSUBS 0.007361f
C274 B.n234 VSUBS 0.007361f
C275 B.n235 VSUBS 0.007361f
C276 B.n236 VSUBS 0.007361f
C277 B.n237 VSUBS 0.007361f
C278 B.n238 VSUBS 0.007361f
C279 B.n239 VSUBS 0.007361f
C280 B.n240 VSUBS 0.018725f
C281 B.n241 VSUBS 0.017923f
C282 B.n242 VSUBS 0.018451f
C283 B.n243 VSUBS 0.007361f
C284 B.n244 VSUBS 0.007361f
C285 B.n245 VSUBS 0.007361f
C286 B.n246 VSUBS 0.007361f
C287 B.n247 VSUBS 0.007361f
C288 B.n248 VSUBS 0.007361f
C289 B.n249 VSUBS 0.007361f
C290 B.n250 VSUBS 0.007361f
C291 B.n251 VSUBS 0.007361f
C292 B.n252 VSUBS 0.007361f
C293 B.n253 VSUBS 0.007361f
C294 B.n254 VSUBS 0.007361f
C295 B.n255 VSUBS 0.007361f
C296 B.n256 VSUBS 0.007361f
C297 B.n257 VSUBS 0.007361f
C298 B.n258 VSUBS 0.007361f
C299 B.n259 VSUBS 0.007361f
C300 B.n260 VSUBS 0.007361f
C301 B.n261 VSUBS 0.007361f
C302 B.n262 VSUBS 0.007361f
C303 B.n263 VSUBS 0.007361f
C304 B.n264 VSUBS 0.007361f
C305 B.n265 VSUBS 0.007361f
C306 B.n266 VSUBS 0.007361f
C307 B.n267 VSUBS 0.007361f
C308 B.n268 VSUBS 0.007361f
C309 B.n269 VSUBS 0.007361f
C310 B.n270 VSUBS 0.007361f
C311 B.n271 VSUBS 0.007361f
C312 B.n272 VSUBS 0.007361f
C313 B.n273 VSUBS 0.007361f
C314 B.n274 VSUBS 0.007361f
C315 B.n275 VSUBS 0.007361f
C316 B.n276 VSUBS 0.007361f
C317 B.n277 VSUBS 0.007361f
C318 B.n278 VSUBS 0.007361f
C319 B.n279 VSUBS 0.007361f
C320 B.n280 VSUBS 0.007361f
C321 B.n281 VSUBS 0.007361f
C322 B.n282 VSUBS 0.007361f
C323 B.n283 VSUBS 0.007361f
C324 B.n284 VSUBS 0.007361f
C325 B.n285 VSUBS 0.007361f
C326 B.n286 VSUBS 0.007361f
C327 B.n287 VSUBS 0.007361f
C328 B.n288 VSUBS 0.007361f
C329 B.n289 VSUBS 0.007361f
C330 B.n290 VSUBS 0.007361f
C331 B.n291 VSUBS 0.007361f
C332 B.n292 VSUBS 0.007361f
C333 B.n293 VSUBS 0.007361f
C334 B.n294 VSUBS 0.007361f
C335 B.n295 VSUBS 0.007361f
C336 B.n296 VSUBS 0.007361f
C337 B.n297 VSUBS 0.007361f
C338 B.n298 VSUBS 0.007361f
C339 B.n299 VSUBS 0.007361f
C340 B.n300 VSUBS 0.007361f
C341 B.n301 VSUBS 0.007361f
C342 B.n302 VSUBS 0.007361f
C343 B.n303 VSUBS 0.007361f
C344 B.n304 VSUBS 0.007361f
C345 B.n305 VSUBS 0.007361f
C346 B.n306 VSUBS 0.007361f
C347 B.n307 VSUBS 0.007361f
C348 B.n308 VSUBS 0.007361f
C349 B.n309 VSUBS 0.007361f
C350 B.n310 VSUBS 0.007361f
C351 B.n311 VSUBS 0.007361f
C352 B.n312 VSUBS 0.007361f
C353 B.n313 VSUBS 0.007361f
C354 B.n314 VSUBS 0.007361f
C355 B.n315 VSUBS 0.007361f
C356 B.n316 VSUBS 0.007361f
C357 B.n317 VSUBS 0.007361f
C358 B.n318 VSUBS 0.007361f
C359 B.n319 VSUBS 0.007361f
C360 B.n320 VSUBS 0.007361f
C361 B.n321 VSUBS 0.007361f
C362 B.n322 VSUBS 0.007361f
C363 B.n323 VSUBS 0.007361f
C364 B.n324 VSUBS 0.007361f
C365 B.n325 VSUBS 0.007361f
C366 B.n326 VSUBS 0.007361f
C367 B.n327 VSUBS 0.007361f
C368 B.n328 VSUBS 0.007361f
C369 B.n329 VSUBS 0.007361f
C370 B.n330 VSUBS 0.007361f
C371 B.n331 VSUBS 0.007361f
C372 B.n332 VSUBS 0.007361f
C373 B.n333 VSUBS 0.007361f
C374 B.n334 VSUBS 0.007361f
C375 B.n335 VSUBS 0.007361f
C376 B.n336 VSUBS 0.007361f
C377 B.n337 VSUBS 0.007361f
C378 B.n338 VSUBS 0.007361f
C379 B.n339 VSUBS 0.007361f
C380 B.n340 VSUBS 0.007361f
C381 B.n341 VSUBS 0.007361f
C382 B.n342 VSUBS 0.007361f
C383 B.n343 VSUBS 0.007361f
C384 B.n344 VSUBS 0.007361f
C385 B.n345 VSUBS 0.007361f
C386 B.n346 VSUBS 0.007361f
C387 B.n347 VSUBS 0.007361f
C388 B.n348 VSUBS 0.017649f
C389 B.n349 VSUBS 0.017649f
C390 B.n350 VSUBS 0.018725f
C391 B.n351 VSUBS 0.007361f
C392 B.n352 VSUBS 0.007361f
C393 B.n353 VSUBS 0.007361f
C394 B.n354 VSUBS 0.007361f
C395 B.n355 VSUBS 0.007361f
C396 B.n356 VSUBS 0.007361f
C397 B.n357 VSUBS 0.007361f
C398 B.n358 VSUBS 0.007361f
C399 B.n359 VSUBS 0.007361f
C400 B.n360 VSUBS 0.007361f
C401 B.n361 VSUBS 0.007361f
C402 B.n362 VSUBS 0.007361f
C403 B.n363 VSUBS 0.007361f
C404 B.n364 VSUBS 0.007361f
C405 B.n365 VSUBS 0.007361f
C406 B.n366 VSUBS 0.007361f
C407 B.n367 VSUBS 0.007361f
C408 B.n368 VSUBS 0.007361f
C409 B.n369 VSUBS 0.007361f
C410 B.n370 VSUBS 0.007361f
C411 B.n371 VSUBS 0.007361f
C412 B.n372 VSUBS 0.007361f
C413 B.n373 VSUBS 0.007361f
C414 B.n374 VSUBS 0.005088f
C415 B.n375 VSUBS 0.017055f
C416 B.n376 VSUBS 0.005954f
C417 B.n377 VSUBS 0.007361f
C418 B.n378 VSUBS 0.007361f
C419 B.n379 VSUBS 0.007361f
C420 B.n380 VSUBS 0.007361f
C421 B.n381 VSUBS 0.007361f
C422 B.n382 VSUBS 0.007361f
C423 B.n383 VSUBS 0.007361f
C424 B.n384 VSUBS 0.007361f
C425 B.n385 VSUBS 0.007361f
C426 B.n386 VSUBS 0.007361f
C427 B.n387 VSUBS 0.007361f
C428 B.n388 VSUBS 0.005954f
C429 B.n389 VSUBS 0.007361f
C430 B.n390 VSUBS 0.007361f
C431 B.n391 VSUBS 0.005088f
C432 B.n392 VSUBS 0.007361f
C433 B.n393 VSUBS 0.007361f
C434 B.n394 VSUBS 0.007361f
C435 B.n395 VSUBS 0.007361f
C436 B.n396 VSUBS 0.007361f
C437 B.n397 VSUBS 0.007361f
C438 B.n398 VSUBS 0.007361f
C439 B.n399 VSUBS 0.007361f
C440 B.n400 VSUBS 0.007361f
C441 B.n401 VSUBS 0.007361f
C442 B.n402 VSUBS 0.007361f
C443 B.n403 VSUBS 0.007361f
C444 B.n404 VSUBS 0.007361f
C445 B.n405 VSUBS 0.007361f
C446 B.n406 VSUBS 0.007361f
C447 B.n407 VSUBS 0.007361f
C448 B.n408 VSUBS 0.007361f
C449 B.n409 VSUBS 0.007361f
C450 B.n410 VSUBS 0.007361f
C451 B.n411 VSUBS 0.007361f
C452 B.n412 VSUBS 0.007361f
C453 B.n413 VSUBS 0.007361f
C454 B.n414 VSUBS 0.018725f
C455 B.n415 VSUBS 0.018725f
C456 B.n416 VSUBS 0.017649f
C457 B.n417 VSUBS 0.007361f
C458 B.n418 VSUBS 0.007361f
C459 B.n419 VSUBS 0.007361f
C460 B.n420 VSUBS 0.007361f
C461 B.n421 VSUBS 0.007361f
C462 B.n422 VSUBS 0.007361f
C463 B.n423 VSUBS 0.007361f
C464 B.n424 VSUBS 0.007361f
C465 B.n425 VSUBS 0.007361f
C466 B.n426 VSUBS 0.007361f
C467 B.n427 VSUBS 0.007361f
C468 B.n428 VSUBS 0.007361f
C469 B.n429 VSUBS 0.007361f
C470 B.n430 VSUBS 0.007361f
C471 B.n431 VSUBS 0.007361f
C472 B.n432 VSUBS 0.007361f
C473 B.n433 VSUBS 0.007361f
C474 B.n434 VSUBS 0.007361f
C475 B.n435 VSUBS 0.007361f
C476 B.n436 VSUBS 0.007361f
C477 B.n437 VSUBS 0.007361f
C478 B.n438 VSUBS 0.007361f
C479 B.n439 VSUBS 0.007361f
C480 B.n440 VSUBS 0.007361f
C481 B.n441 VSUBS 0.007361f
C482 B.n442 VSUBS 0.007361f
C483 B.n443 VSUBS 0.007361f
C484 B.n444 VSUBS 0.007361f
C485 B.n445 VSUBS 0.007361f
C486 B.n446 VSUBS 0.007361f
C487 B.n447 VSUBS 0.007361f
C488 B.n448 VSUBS 0.007361f
C489 B.n449 VSUBS 0.007361f
C490 B.n450 VSUBS 0.007361f
C491 B.n451 VSUBS 0.007361f
C492 B.n452 VSUBS 0.007361f
C493 B.n453 VSUBS 0.007361f
C494 B.n454 VSUBS 0.007361f
C495 B.n455 VSUBS 0.007361f
C496 B.n456 VSUBS 0.007361f
C497 B.n457 VSUBS 0.007361f
C498 B.n458 VSUBS 0.007361f
C499 B.n459 VSUBS 0.007361f
C500 B.n460 VSUBS 0.007361f
C501 B.n461 VSUBS 0.007361f
C502 B.n462 VSUBS 0.007361f
C503 B.n463 VSUBS 0.007361f
C504 B.n464 VSUBS 0.007361f
C505 B.n465 VSUBS 0.007361f
C506 B.n466 VSUBS 0.007361f
C507 B.n467 VSUBS 0.009606f
C508 B.n468 VSUBS 0.010233f
C509 B.n469 VSUBS 0.020349f
C510 VDD2.t5 VSUBS 0.489308f
C511 VDD2.t2 VSUBS 0.062008f
C512 VDD2.t3 VSUBS 0.062008f
C513 VDD2.n0 VSUBS 0.349087f
C514 VDD2.n1 VSUBS 2.11877f
C515 VDD2.t0 VSUBS 0.484364f
C516 VDD2.n2 VSUBS 1.83369f
C517 VDD2.t1 VSUBS 0.062008f
C518 VDD2.t4 VSUBS 0.062008f
C519 VDD2.n3 VSUBS 0.34907f
C520 VN.n0 VSUBS 0.065148f
C521 VN.t2 VSUBS 0.897066f
C522 VN.n1 VSUBS 0.061581f
C523 VN.t0 VSUBS 1.17598f
C524 VN.n2 VSUBS 0.473284f
C525 VN.t3 VSUBS 0.897066f
C526 VN.n3 VSUBS 0.51948f
C527 VN.n4 VSUBS 0.09164f
C528 VN.n5 VSUBS 0.412352f
C529 VN.n6 VSUBS 0.049417f
C530 VN.n7 VSUBS 0.049417f
C531 VN.n8 VSUBS 0.08209f
C532 VN.n9 VSUBS 0.078068f
C533 VN.n10 VSUBS 0.519762f
C534 VN.n11 VSUBS 0.063763f
C535 VN.n12 VSUBS 0.065148f
C536 VN.t5 VSUBS 0.897066f
C537 VN.n13 VSUBS 0.061581f
C538 VN.t1 VSUBS 1.17598f
C539 VN.n14 VSUBS 0.473284f
C540 VN.t4 VSUBS 0.897066f
C541 VN.n15 VSUBS 0.51948f
C542 VN.n16 VSUBS 0.09164f
C543 VN.n17 VSUBS 0.412352f
C544 VN.n18 VSUBS 0.049417f
C545 VN.n19 VSUBS 0.049417f
C546 VN.n20 VSUBS 0.08209f
C547 VN.n21 VSUBS 0.078068f
C548 VN.n22 VSUBS 0.519762f
C549 VN.n23 VSUBS 1.94825f
C550 VDD1.t1 VSUBS 0.498573f
C551 VDD1.t2 VSUBS 0.49809f
C552 VDD1.t0 VSUBS 0.063121f
C553 VDD1.t3 VSUBS 0.063121f
C554 VDD1.n0 VSUBS 0.355352f
C555 VDD1.n1 VSUBS 2.24862f
C556 VDD1.t4 VSUBS 0.063121f
C557 VDD1.t5 VSUBS 0.063121f
C558 VDD1.n2 VSUBS 0.353515f
C559 VDD1.n3 VSUBS 1.8907f
C560 VTAIL.t4 VSUBS 0.082261f
C561 VTAIL.t2 VSUBS 0.082261f
C562 VTAIL.n0 VSUBS 0.398207f
C563 VTAIL.n1 VSUBS 0.613378f
C564 VTAIL.t10 VSUBS 0.578875f
C565 VTAIL.n2 VSUBS 0.795514f
C566 VTAIL.t9 VSUBS 0.082261f
C567 VTAIL.t11 VSUBS 0.082261f
C568 VTAIL.n3 VSUBS 0.398207f
C569 VTAIL.n4 VSUBS 1.68386f
C570 VTAIL.t0 VSUBS 0.082261f
C571 VTAIL.t1 VSUBS 0.082261f
C572 VTAIL.n5 VSUBS 0.398209f
C573 VTAIL.n6 VSUBS 1.68386f
C574 VTAIL.t3 VSUBS 0.578878f
C575 VTAIL.n7 VSUBS 0.795511f
C576 VTAIL.t6 VSUBS 0.082261f
C577 VTAIL.t7 VSUBS 0.082261f
C578 VTAIL.n8 VSUBS 0.398209f
C579 VTAIL.n9 VSUBS 0.75183f
C580 VTAIL.t8 VSUBS 0.578875f
C581 VTAIL.n10 VSUBS 1.53558f
C582 VTAIL.t5 VSUBS 0.578875f
C583 VTAIL.n11 VSUBS 1.48208f
C584 VP.n0 VSUBS 0.068574f
C585 VP.t2 VSUBS 0.944246f
C586 VP.n1 VSUBS 0.06482f
C587 VP.n2 VSUBS 0.052016f
C588 VP.t5 VSUBS 0.944246f
C589 VP.n3 VSUBS 0.06482f
C590 VP.n4 VSUBS 0.068574f
C591 VP.t3 VSUBS 0.944246f
C592 VP.n5 VSUBS 0.068574f
C593 VP.t0 VSUBS 0.944246f
C594 VP.n6 VSUBS 0.06482f
C595 VP.t4 VSUBS 1.23783f
C596 VP.n7 VSUBS 0.498175f
C597 VP.t1 VSUBS 0.944246f
C598 VP.n8 VSUBS 0.546801f
C599 VP.n9 VSUBS 0.096459f
C600 VP.n10 VSUBS 0.434039f
C601 VP.n11 VSUBS 0.052016f
C602 VP.n12 VSUBS 0.052016f
C603 VP.n13 VSUBS 0.086407f
C604 VP.n14 VSUBS 0.082173f
C605 VP.n15 VSUBS 0.547098f
C606 VP.n16 VSUBS 2.02165f
C607 VP.n17 VSUBS 2.06856f
C608 VP.n18 VSUBS 0.547098f
C609 VP.n19 VSUBS 0.082173f
C610 VP.n20 VSUBS 0.086407f
C611 VP.n21 VSUBS 0.052016f
C612 VP.n22 VSUBS 0.052016f
C613 VP.n23 VSUBS 0.052016f
C614 VP.n24 VSUBS 0.096459f
C615 VP.n25 VSUBS 0.443926f
C616 VP.n26 VSUBS 0.096459f
C617 VP.n27 VSUBS 0.052016f
C618 VP.n28 VSUBS 0.052016f
C619 VP.n29 VSUBS 0.052016f
C620 VP.n30 VSUBS 0.086407f
C621 VP.n31 VSUBS 0.082173f
C622 VP.n32 VSUBS 0.547098f
C623 VP.n33 VSUBS 0.067117f
.ends

