* NGSPICE file created from diff_pair_sample_0419.ext - technology: sky130A

.subckt diff_pair_sample_0419 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0 ps=0 w=0.64 l=1.31
X1 B.t8 B.t6 B.t7 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0 ps=0 w=0.64 l=1.31
X2 VDD1.t7 VP.t0 VTAIL.t10 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X3 VDD2.t7 VN.t0 VTAIL.t7 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.2496 ps=2.06 w=0.64 l=1.31
X4 VDD2.t6 VN.t1 VTAIL.t0 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.2496 ps=2.06 w=0.64 l=1.31
X5 VTAIL.t4 VN.t2 VDD2.t5 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X6 VDD2.t4 VN.t3 VTAIL.t6 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X7 B.t5 B.t3 B.t4 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0 ps=0 w=0.64 l=1.31
X8 B.t2 B.t0 B.t1 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0 ps=0 w=0.64 l=1.31
X9 VTAIL.t2 VN.t4 VDD2.t3 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X10 VDD1.t6 VP.t1 VTAIL.t8 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.2496 ps=2.06 w=0.64 l=1.31
X11 VTAIL.t9 VP.t2 VDD1.t5 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X12 VTAIL.t15 VP.t3 VDD1.t4 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X13 VTAIL.t3 VN.t5 VDD2.t2 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0.1056 ps=0.97 w=0.64 l=1.31
X14 VDD1.t3 VP.t4 VTAIL.t11 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X15 VTAIL.t14 VP.t5 VDD1.t2 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0.1056 ps=0.97 w=0.64 l=1.31
X16 VDD2.t1 VN.t6 VTAIL.t5 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.1056 ps=0.97 w=0.64 l=1.31
X17 VDD1.t1 VP.t6 VTAIL.t13 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.1056 pd=0.97 as=0.2496 ps=2.06 w=0.64 l=1.31
X18 VTAIL.t1 VN.t7 VDD2.t0 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0.1056 ps=0.97 w=0.64 l=1.31
X19 VTAIL.t12 VP.t7 VDD1.t0 w_n2610_n1096# sky130_fd_pr__pfet_01v8 ad=0.2496 pd=2.06 as=0.1056 ps=0.97 w=0.64 l=1.31
R0 B.n72 B.t11 689.899
R1 B.n80 B.t8 689.899
R2 B.n22 B.t1 689.899
R3 B.n30 B.t4 689.899
R4 B.n73 B.t10 658.092
R5 B.n81 B.t7 658.092
R6 B.n23 B.t2 658.092
R7 B.n31 B.t5 658.092
R8 B.n286 B.n35 585
R9 B.n288 B.n287 585
R10 B.n289 B.n34 585
R11 B.n291 B.n290 585
R12 B.n292 B.n33 585
R13 B.n294 B.n293 585
R14 B.n295 B.n32 585
R15 B.n297 B.n296 585
R16 B.n299 B.n29 585
R17 B.n301 B.n300 585
R18 B.n302 B.n28 585
R19 B.n304 B.n303 585
R20 B.n305 B.n27 585
R21 B.n307 B.n306 585
R22 B.n308 B.n26 585
R23 B.n310 B.n309 585
R24 B.n311 B.n25 585
R25 B.n313 B.n312 585
R26 B.n315 B.n314 585
R27 B.n316 B.n21 585
R28 B.n318 B.n317 585
R29 B.n319 B.n20 585
R30 B.n321 B.n320 585
R31 B.n322 B.n19 585
R32 B.n324 B.n323 585
R33 B.n325 B.n18 585
R34 B.n285 B.n284 585
R35 B.n283 B.n36 585
R36 B.n282 B.n281 585
R37 B.n280 B.n37 585
R38 B.n279 B.n278 585
R39 B.n277 B.n38 585
R40 B.n276 B.n275 585
R41 B.n274 B.n39 585
R42 B.n273 B.n272 585
R43 B.n271 B.n40 585
R44 B.n270 B.n269 585
R45 B.n268 B.n41 585
R46 B.n267 B.n266 585
R47 B.n265 B.n42 585
R48 B.n264 B.n263 585
R49 B.n262 B.n43 585
R50 B.n261 B.n260 585
R51 B.n259 B.n44 585
R52 B.n258 B.n257 585
R53 B.n256 B.n45 585
R54 B.n255 B.n254 585
R55 B.n253 B.n46 585
R56 B.n252 B.n251 585
R57 B.n250 B.n47 585
R58 B.n249 B.n248 585
R59 B.n247 B.n48 585
R60 B.n246 B.n245 585
R61 B.n244 B.n49 585
R62 B.n243 B.n242 585
R63 B.n241 B.n50 585
R64 B.n240 B.n239 585
R65 B.n238 B.n51 585
R66 B.n237 B.n236 585
R67 B.n235 B.n52 585
R68 B.n234 B.n233 585
R69 B.n232 B.n53 585
R70 B.n231 B.n230 585
R71 B.n229 B.n54 585
R72 B.n228 B.n227 585
R73 B.n226 B.n55 585
R74 B.n225 B.n224 585
R75 B.n223 B.n56 585
R76 B.n222 B.n221 585
R77 B.n220 B.n57 585
R78 B.n219 B.n218 585
R79 B.n217 B.n58 585
R80 B.n216 B.n215 585
R81 B.n214 B.n59 585
R82 B.n213 B.n212 585
R83 B.n211 B.n60 585
R84 B.n210 B.n209 585
R85 B.n208 B.n61 585
R86 B.n207 B.n206 585
R87 B.n205 B.n62 585
R88 B.n204 B.n203 585
R89 B.n202 B.n63 585
R90 B.n201 B.n200 585
R91 B.n199 B.n64 585
R92 B.n198 B.n197 585
R93 B.n196 B.n65 585
R94 B.n195 B.n194 585
R95 B.n193 B.n66 585
R96 B.n192 B.n191 585
R97 B.n190 B.n67 585
R98 B.n189 B.n188 585
R99 B.n148 B.n85 585
R100 B.n150 B.n149 585
R101 B.n151 B.n84 585
R102 B.n153 B.n152 585
R103 B.n154 B.n83 585
R104 B.n156 B.n155 585
R105 B.n157 B.n82 585
R106 B.n159 B.n158 585
R107 B.n161 B.n79 585
R108 B.n163 B.n162 585
R109 B.n164 B.n78 585
R110 B.n166 B.n165 585
R111 B.n167 B.n77 585
R112 B.n169 B.n168 585
R113 B.n170 B.n76 585
R114 B.n172 B.n171 585
R115 B.n173 B.n75 585
R116 B.n175 B.n174 585
R117 B.n177 B.n176 585
R118 B.n178 B.n71 585
R119 B.n180 B.n179 585
R120 B.n181 B.n70 585
R121 B.n183 B.n182 585
R122 B.n184 B.n69 585
R123 B.n186 B.n185 585
R124 B.n187 B.n68 585
R125 B.n147 B.n146 585
R126 B.n145 B.n86 585
R127 B.n144 B.n143 585
R128 B.n142 B.n87 585
R129 B.n141 B.n140 585
R130 B.n139 B.n88 585
R131 B.n138 B.n137 585
R132 B.n136 B.n89 585
R133 B.n135 B.n134 585
R134 B.n133 B.n90 585
R135 B.n132 B.n131 585
R136 B.n130 B.n91 585
R137 B.n129 B.n128 585
R138 B.n127 B.n92 585
R139 B.n126 B.n125 585
R140 B.n124 B.n93 585
R141 B.n123 B.n122 585
R142 B.n121 B.n94 585
R143 B.n120 B.n119 585
R144 B.n118 B.n95 585
R145 B.n117 B.n116 585
R146 B.n115 B.n96 585
R147 B.n114 B.n113 585
R148 B.n112 B.n97 585
R149 B.n111 B.n110 585
R150 B.n109 B.n98 585
R151 B.n108 B.n107 585
R152 B.n106 B.n99 585
R153 B.n105 B.n104 585
R154 B.n103 B.n100 585
R155 B.n102 B.n101 585
R156 B.n2 B.n0 585
R157 B.n373 B.n1 585
R158 B.n372 B.n371 585
R159 B.n370 B.n3 585
R160 B.n369 B.n368 585
R161 B.n367 B.n4 585
R162 B.n366 B.n365 585
R163 B.n364 B.n5 585
R164 B.n363 B.n362 585
R165 B.n361 B.n6 585
R166 B.n360 B.n359 585
R167 B.n358 B.n7 585
R168 B.n357 B.n356 585
R169 B.n355 B.n8 585
R170 B.n354 B.n353 585
R171 B.n352 B.n9 585
R172 B.n351 B.n350 585
R173 B.n349 B.n10 585
R174 B.n348 B.n347 585
R175 B.n346 B.n11 585
R176 B.n345 B.n344 585
R177 B.n343 B.n12 585
R178 B.n342 B.n341 585
R179 B.n340 B.n13 585
R180 B.n339 B.n338 585
R181 B.n337 B.n14 585
R182 B.n336 B.n335 585
R183 B.n334 B.n15 585
R184 B.n333 B.n332 585
R185 B.n331 B.n16 585
R186 B.n330 B.n329 585
R187 B.n328 B.n17 585
R188 B.n327 B.n326 585
R189 B.n375 B.n374 585
R190 B.n146 B.n85 535.745
R191 B.n326 B.n325 535.745
R192 B.n188 B.n187 535.745
R193 B.n284 B.n35 535.745
R194 B.n72 B.t9 207.482
R195 B.n30 B.t3 207.482
R196 B.n80 B.t6 207.084
R197 B.n22 B.t0 207.084
R198 B.n146 B.n145 163.367
R199 B.n145 B.n144 163.367
R200 B.n144 B.n87 163.367
R201 B.n140 B.n87 163.367
R202 B.n140 B.n139 163.367
R203 B.n139 B.n138 163.367
R204 B.n138 B.n89 163.367
R205 B.n134 B.n89 163.367
R206 B.n134 B.n133 163.367
R207 B.n133 B.n132 163.367
R208 B.n132 B.n91 163.367
R209 B.n128 B.n91 163.367
R210 B.n128 B.n127 163.367
R211 B.n127 B.n126 163.367
R212 B.n126 B.n93 163.367
R213 B.n122 B.n93 163.367
R214 B.n122 B.n121 163.367
R215 B.n121 B.n120 163.367
R216 B.n120 B.n95 163.367
R217 B.n116 B.n95 163.367
R218 B.n116 B.n115 163.367
R219 B.n115 B.n114 163.367
R220 B.n114 B.n97 163.367
R221 B.n110 B.n97 163.367
R222 B.n110 B.n109 163.367
R223 B.n109 B.n108 163.367
R224 B.n108 B.n99 163.367
R225 B.n104 B.n99 163.367
R226 B.n104 B.n103 163.367
R227 B.n103 B.n102 163.367
R228 B.n102 B.n2 163.367
R229 B.n374 B.n2 163.367
R230 B.n374 B.n373 163.367
R231 B.n373 B.n372 163.367
R232 B.n372 B.n3 163.367
R233 B.n368 B.n3 163.367
R234 B.n368 B.n367 163.367
R235 B.n367 B.n366 163.367
R236 B.n366 B.n5 163.367
R237 B.n362 B.n5 163.367
R238 B.n362 B.n361 163.367
R239 B.n361 B.n360 163.367
R240 B.n360 B.n7 163.367
R241 B.n356 B.n7 163.367
R242 B.n356 B.n355 163.367
R243 B.n355 B.n354 163.367
R244 B.n354 B.n9 163.367
R245 B.n350 B.n9 163.367
R246 B.n350 B.n349 163.367
R247 B.n349 B.n348 163.367
R248 B.n348 B.n11 163.367
R249 B.n344 B.n11 163.367
R250 B.n344 B.n343 163.367
R251 B.n343 B.n342 163.367
R252 B.n342 B.n13 163.367
R253 B.n338 B.n13 163.367
R254 B.n338 B.n337 163.367
R255 B.n337 B.n336 163.367
R256 B.n336 B.n15 163.367
R257 B.n332 B.n15 163.367
R258 B.n332 B.n331 163.367
R259 B.n331 B.n330 163.367
R260 B.n330 B.n17 163.367
R261 B.n326 B.n17 163.367
R262 B.n150 B.n85 163.367
R263 B.n151 B.n150 163.367
R264 B.n152 B.n151 163.367
R265 B.n152 B.n83 163.367
R266 B.n156 B.n83 163.367
R267 B.n157 B.n156 163.367
R268 B.n158 B.n157 163.367
R269 B.n158 B.n79 163.367
R270 B.n163 B.n79 163.367
R271 B.n164 B.n163 163.367
R272 B.n165 B.n164 163.367
R273 B.n165 B.n77 163.367
R274 B.n169 B.n77 163.367
R275 B.n170 B.n169 163.367
R276 B.n171 B.n170 163.367
R277 B.n171 B.n75 163.367
R278 B.n175 B.n75 163.367
R279 B.n176 B.n175 163.367
R280 B.n176 B.n71 163.367
R281 B.n180 B.n71 163.367
R282 B.n181 B.n180 163.367
R283 B.n182 B.n181 163.367
R284 B.n182 B.n69 163.367
R285 B.n186 B.n69 163.367
R286 B.n187 B.n186 163.367
R287 B.n188 B.n67 163.367
R288 B.n192 B.n67 163.367
R289 B.n193 B.n192 163.367
R290 B.n194 B.n193 163.367
R291 B.n194 B.n65 163.367
R292 B.n198 B.n65 163.367
R293 B.n199 B.n198 163.367
R294 B.n200 B.n199 163.367
R295 B.n200 B.n63 163.367
R296 B.n204 B.n63 163.367
R297 B.n205 B.n204 163.367
R298 B.n206 B.n205 163.367
R299 B.n206 B.n61 163.367
R300 B.n210 B.n61 163.367
R301 B.n211 B.n210 163.367
R302 B.n212 B.n211 163.367
R303 B.n212 B.n59 163.367
R304 B.n216 B.n59 163.367
R305 B.n217 B.n216 163.367
R306 B.n218 B.n217 163.367
R307 B.n218 B.n57 163.367
R308 B.n222 B.n57 163.367
R309 B.n223 B.n222 163.367
R310 B.n224 B.n223 163.367
R311 B.n224 B.n55 163.367
R312 B.n228 B.n55 163.367
R313 B.n229 B.n228 163.367
R314 B.n230 B.n229 163.367
R315 B.n230 B.n53 163.367
R316 B.n234 B.n53 163.367
R317 B.n235 B.n234 163.367
R318 B.n236 B.n235 163.367
R319 B.n236 B.n51 163.367
R320 B.n240 B.n51 163.367
R321 B.n241 B.n240 163.367
R322 B.n242 B.n241 163.367
R323 B.n242 B.n49 163.367
R324 B.n246 B.n49 163.367
R325 B.n247 B.n246 163.367
R326 B.n248 B.n247 163.367
R327 B.n248 B.n47 163.367
R328 B.n252 B.n47 163.367
R329 B.n253 B.n252 163.367
R330 B.n254 B.n253 163.367
R331 B.n254 B.n45 163.367
R332 B.n258 B.n45 163.367
R333 B.n259 B.n258 163.367
R334 B.n260 B.n259 163.367
R335 B.n260 B.n43 163.367
R336 B.n264 B.n43 163.367
R337 B.n265 B.n264 163.367
R338 B.n266 B.n265 163.367
R339 B.n266 B.n41 163.367
R340 B.n270 B.n41 163.367
R341 B.n271 B.n270 163.367
R342 B.n272 B.n271 163.367
R343 B.n272 B.n39 163.367
R344 B.n276 B.n39 163.367
R345 B.n277 B.n276 163.367
R346 B.n278 B.n277 163.367
R347 B.n278 B.n37 163.367
R348 B.n282 B.n37 163.367
R349 B.n283 B.n282 163.367
R350 B.n284 B.n283 163.367
R351 B.n325 B.n324 163.367
R352 B.n324 B.n19 163.367
R353 B.n320 B.n19 163.367
R354 B.n320 B.n319 163.367
R355 B.n319 B.n318 163.367
R356 B.n318 B.n21 163.367
R357 B.n314 B.n21 163.367
R358 B.n314 B.n313 163.367
R359 B.n313 B.n25 163.367
R360 B.n309 B.n25 163.367
R361 B.n309 B.n308 163.367
R362 B.n308 B.n307 163.367
R363 B.n307 B.n27 163.367
R364 B.n303 B.n27 163.367
R365 B.n303 B.n302 163.367
R366 B.n302 B.n301 163.367
R367 B.n301 B.n29 163.367
R368 B.n296 B.n29 163.367
R369 B.n296 B.n295 163.367
R370 B.n295 B.n294 163.367
R371 B.n294 B.n33 163.367
R372 B.n290 B.n33 163.367
R373 B.n290 B.n289 163.367
R374 B.n289 B.n288 163.367
R375 B.n288 B.n35 163.367
R376 B.n74 B.n73 59.5399
R377 B.n160 B.n81 59.5399
R378 B.n24 B.n23 59.5399
R379 B.n298 B.n31 59.5399
R380 B.n327 B.n18 34.8103
R381 B.n286 B.n285 34.8103
R382 B.n189 B.n68 34.8103
R383 B.n148 B.n147 34.8103
R384 B.n73 B.n72 31.8066
R385 B.n81 B.n80 31.8066
R386 B.n23 B.n22 31.8066
R387 B.n31 B.n30 31.8066
R388 B B.n375 18.0485
R389 B.n323 B.n18 10.6151
R390 B.n323 B.n322 10.6151
R391 B.n322 B.n321 10.6151
R392 B.n321 B.n20 10.6151
R393 B.n317 B.n20 10.6151
R394 B.n317 B.n316 10.6151
R395 B.n316 B.n315 10.6151
R396 B.n312 B.n311 10.6151
R397 B.n311 B.n310 10.6151
R398 B.n310 B.n26 10.6151
R399 B.n306 B.n26 10.6151
R400 B.n306 B.n305 10.6151
R401 B.n305 B.n304 10.6151
R402 B.n304 B.n28 10.6151
R403 B.n300 B.n28 10.6151
R404 B.n300 B.n299 10.6151
R405 B.n297 B.n32 10.6151
R406 B.n293 B.n32 10.6151
R407 B.n293 B.n292 10.6151
R408 B.n292 B.n291 10.6151
R409 B.n291 B.n34 10.6151
R410 B.n287 B.n34 10.6151
R411 B.n287 B.n286 10.6151
R412 B.n190 B.n189 10.6151
R413 B.n191 B.n190 10.6151
R414 B.n191 B.n66 10.6151
R415 B.n195 B.n66 10.6151
R416 B.n196 B.n195 10.6151
R417 B.n197 B.n196 10.6151
R418 B.n197 B.n64 10.6151
R419 B.n201 B.n64 10.6151
R420 B.n202 B.n201 10.6151
R421 B.n203 B.n202 10.6151
R422 B.n203 B.n62 10.6151
R423 B.n207 B.n62 10.6151
R424 B.n208 B.n207 10.6151
R425 B.n209 B.n208 10.6151
R426 B.n209 B.n60 10.6151
R427 B.n213 B.n60 10.6151
R428 B.n214 B.n213 10.6151
R429 B.n215 B.n214 10.6151
R430 B.n215 B.n58 10.6151
R431 B.n219 B.n58 10.6151
R432 B.n220 B.n219 10.6151
R433 B.n221 B.n220 10.6151
R434 B.n221 B.n56 10.6151
R435 B.n225 B.n56 10.6151
R436 B.n226 B.n225 10.6151
R437 B.n227 B.n226 10.6151
R438 B.n227 B.n54 10.6151
R439 B.n231 B.n54 10.6151
R440 B.n232 B.n231 10.6151
R441 B.n233 B.n232 10.6151
R442 B.n233 B.n52 10.6151
R443 B.n237 B.n52 10.6151
R444 B.n238 B.n237 10.6151
R445 B.n239 B.n238 10.6151
R446 B.n239 B.n50 10.6151
R447 B.n243 B.n50 10.6151
R448 B.n244 B.n243 10.6151
R449 B.n245 B.n244 10.6151
R450 B.n245 B.n48 10.6151
R451 B.n249 B.n48 10.6151
R452 B.n250 B.n249 10.6151
R453 B.n251 B.n250 10.6151
R454 B.n251 B.n46 10.6151
R455 B.n255 B.n46 10.6151
R456 B.n256 B.n255 10.6151
R457 B.n257 B.n256 10.6151
R458 B.n257 B.n44 10.6151
R459 B.n261 B.n44 10.6151
R460 B.n262 B.n261 10.6151
R461 B.n263 B.n262 10.6151
R462 B.n263 B.n42 10.6151
R463 B.n267 B.n42 10.6151
R464 B.n268 B.n267 10.6151
R465 B.n269 B.n268 10.6151
R466 B.n269 B.n40 10.6151
R467 B.n273 B.n40 10.6151
R468 B.n274 B.n273 10.6151
R469 B.n275 B.n274 10.6151
R470 B.n275 B.n38 10.6151
R471 B.n279 B.n38 10.6151
R472 B.n280 B.n279 10.6151
R473 B.n281 B.n280 10.6151
R474 B.n281 B.n36 10.6151
R475 B.n285 B.n36 10.6151
R476 B.n149 B.n148 10.6151
R477 B.n149 B.n84 10.6151
R478 B.n153 B.n84 10.6151
R479 B.n154 B.n153 10.6151
R480 B.n155 B.n154 10.6151
R481 B.n155 B.n82 10.6151
R482 B.n159 B.n82 10.6151
R483 B.n162 B.n161 10.6151
R484 B.n162 B.n78 10.6151
R485 B.n166 B.n78 10.6151
R486 B.n167 B.n166 10.6151
R487 B.n168 B.n167 10.6151
R488 B.n168 B.n76 10.6151
R489 B.n172 B.n76 10.6151
R490 B.n173 B.n172 10.6151
R491 B.n174 B.n173 10.6151
R492 B.n178 B.n177 10.6151
R493 B.n179 B.n178 10.6151
R494 B.n179 B.n70 10.6151
R495 B.n183 B.n70 10.6151
R496 B.n184 B.n183 10.6151
R497 B.n185 B.n184 10.6151
R498 B.n185 B.n68 10.6151
R499 B.n147 B.n86 10.6151
R500 B.n143 B.n86 10.6151
R501 B.n143 B.n142 10.6151
R502 B.n142 B.n141 10.6151
R503 B.n141 B.n88 10.6151
R504 B.n137 B.n88 10.6151
R505 B.n137 B.n136 10.6151
R506 B.n136 B.n135 10.6151
R507 B.n135 B.n90 10.6151
R508 B.n131 B.n90 10.6151
R509 B.n131 B.n130 10.6151
R510 B.n130 B.n129 10.6151
R511 B.n129 B.n92 10.6151
R512 B.n125 B.n92 10.6151
R513 B.n125 B.n124 10.6151
R514 B.n124 B.n123 10.6151
R515 B.n123 B.n94 10.6151
R516 B.n119 B.n94 10.6151
R517 B.n119 B.n118 10.6151
R518 B.n118 B.n117 10.6151
R519 B.n117 B.n96 10.6151
R520 B.n113 B.n96 10.6151
R521 B.n113 B.n112 10.6151
R522 B.n112 B.n111 10.6151
R523 B.n111 B.n98 10.6151
R524 B.n107 B.n98 10.6151
R525 B.n107 B.n106 10.6151
R526 B.n106 B.n105 10.6151
R527 B.n105 B.n100 10.6151
R528 B.n101 B.n100 10.6151
R529 B.n101 B.n0 10.6151
R530 B.n371 B.n1 10.6151
R531 B.n371 B.n370 10.6151
R532 B.n370 B.n369 10.6151
R533 B.n369 B.n4 10.6151
R534 B.n365 B.n4 10.6151
R535 B.n365 B.n364 10.6151
R536 B.n364 B.n363 10.6151
R537 B.n363 B.n6 10.6151
R538 B.n359 B.n6 10.6151
R539 B.n359 B.n358 10.6151
R540 B.n358 B.n357 10.6151
R541 B.n357 B.n8 10.6151
R542 B.n353 B.n8 10.6151
R543 B.n353 B.n352 10.6151
R544 B.n352 B.n351 10.6151
R545 B.n351 B.n10 10.6151
R546 B.n347 B.n10 10.6151
R547 B.n347 B.n346 10.6151
R548 B.n346 B.n345 10.6151
R549 B.n345 B.n12 10.6151
R550 B.n341 B.n12 10.6151
R551 B.n341 B.n340 10.6151
R552 B.n340 B.n339 10.6151
R553 B.n339 B.n14 10.6151
R554 B.n335 B.n14 10.6151
R555 B.n335 B.n334 10.6151
R556 B.n334 B.n333 10.6151
R557 B.n333 B.n16 10.6151
R558 B.n329 B.n16 10.6151
R559 B.n329 B.n328 10.6151
R560 B.n328 B.n327 10.6151
R561 B.n315 B.n24 9.52245
R562 B.n298 B.n297 9.52245
R563 B.n160 B.n159 9.52245
R564 B.n177 B.n74 9.52245
R565 B.n375 B.n0 2.81026
R566 B.n375 B.n1 2.81026
R567 B.n312 B.n24 1.09318
R568 B.n299 B.n298 1.09318
R569 B.n161 B.n160 1.09318
R570 B.n174 B.n74 1.09318
R571 VP.n25 VP.n5 175.419
R572 VP.n44 VP.n43 175.419
R573 VP.n24 VP.n23 175.419
R574 VP.n12 VP.n9 161.3
R575 VP.n14 VP.n13 161.3
R576 VP.n15 VP.n8 161.3
R577 VP.n18 VP.n17 161.3
R578 VP.n19 VP.n7 161.3
R579 VP.n21 VP.n20 161.3
R580 VP.n22 VP.n6 161.3
R581 VP.n42 VP.n0 161.3
R582 VP.n41 VP.n40 161.3
R583 VP.n39 VP.n1 161.3
R584 VP.n38 VP.n37 161.3
R585 VP.n35 VP.n2 161.3
R586 VP.n34 VP.n33 161.3
R587 VP.n32 VP.n3 161.3
R588 VP.n31 VP.n30 161.3
R589 VP.n28 VP.n4 161.3
R590 VP.n27 VP.n26 161.3
R591 VP.n11 VP.n10 61.8956
R592 VP.n35 VP.n34 56.4773
R593 VP.n15 VP.n14 56.4773
R594 VP.n30 VP.n28 51.1217
R595 VP.n41 VP.n1 51.1217
R596 VP.n21 VP.n7 51.1217
R597 VP.n11 VP.t5 39.2192
R598 VP.n25 VP.n24 36.1369
R599 VP.n28 VP.n27 29.6995
R600 VP.n42 VP.n41 29.6995
R601 VP.n22 VP.n21 29.6995
R602 VP.n12 VP.n11 27.6663
R603 VP.n34 VP.n3 24.3439
R604 VP.n37 VP.n35 24.3439
R605 VP.n17 VP.n15 24.3439
R606 VP.n14 VP.n9 24.3439
R607 VP.n30 VP.n29 20.9359
R608 VP.n36 VP.n1 20.9359
R609 VP.n16 VP.n7 20.9359
R610 VP.n5 VP.t7 11.7745
R611 VP.n29 VP.t0 11.7745
R612 VP.n36 VP.t2 11.7745
R613 VP.n43 VP.t6 11.7745
R614 VP.n23 VP.t1 11.7745
R615 VP.n16 VP.t3 11.7745
R616 VP.n10 VP.t4 11.7745
R617 VP.n27 VP.n5 10.2247
R618 VP.n43 VP.n42 10.2247
R619 VP.n23 VP.n22 10.2247
R620 VP.n29 VP.n3 3.40858
R621 VP.n37 VP.n36 3.40858
R622 VP.n17 VP.n16 3.40858
R623 VP.n10 VP.n9 3.40858
R624 VP.n13 VP.n12 0.189894
R625 VP.n13 VP.n8 0.189894
R626 VP.n18 VP.n8 0.189894
R627 VP.n19 VP.n18 0.189894
R628 VP.n20 VP.n19 0.189894
R629 VP.n20 VP.n6 0.189894
R630 VP.n24 VP.n6 0.189894
R631 VP.n26 VP.n25 0.189894
R632 VP.n26 VP.n4 0.189894
R633 VP.n31 VP.n4 0.189894
R634 VP.n32 VP.n31 0.189894
R635 VP.n33 VP.n32 0.189894
R636 VP.n33 VP.n2 0.189894
R637 VP.n38 VP.n2 0.189894
R638 VP.n39 VP.n38 0.189894
R639 VP.n40 VP.n39 0.189894
R640 VP.n40 VP.n0 0.189894
R641 VP.n44 VP.n0 0.189894
R642 VP VP.n44 0.0516364
R643 VTAIL.n15 VTAIL.t7 668.75
R644 VTAIL.n2 VTAIL.t1 668.75
R645 VTAIL.n3 VTAIL.t13 668.75
R646 VTAIL.n6 VTAIL.t12 668.75
R647 VTAIL.n14 VTAIL.t8 668.75
R648 VTAIL.n11 VTAIL.t14 668.75
R649 VTAIL.n10 VTAIL.t0 668.75
R650 VTAIL.n7 VTAIL.t3 668.75
R651 VTAIL.n1 VTAIL.n0 617.962
R652 VTAIL.n5 VTAIL.n4 617.962
R653 VTAIL.n13 VTAIL.n12 617.962
R654 VTAIL.n9 VTAIL.n8 617.962
R655 VTAIL.n0 VTAIL.t5 50.7896
R656 VTAIL.n0 VTAIL.t2 50.7896
R657 VTAIL.n4 VTAIL.t10 50.7896
R658 VTAIL.n4 VTAIL.t9 50.7896
R659 VTAIL.n12 VTAIL.t11 50.7896
R660 VTAIL.n12 VTAIL.t15 50.7896
R661 VTAIL.n8 VTAIL.t6 50.7896
R662 VTAIL.n8 VTAIL.t4 50.7896
R663 VTAIL.n15 VTAIL.n14 14.3324
R664 VTAIL.n7 VTAIL.n6 14.3324
R665 VTAIL.n9 VTAIL.n7 1.41429
R666 VTAIL.n10 VTAIL.n9 1.41429
R667 VTAIL.n13 VTAIL.n11 1.41429
R668 VTAIL.n14 VTAIL.n13 1.41429
R669 VTAIL.n6 VTAIL.n5 1.41429
R670 VTAIL.n5 VTAIL.n3 1.41429
R671 VTAIL.n2 VTAIL.n1 1.41429
R672 VTAIL VTAIL.n15 1.3561
R673 VTAIL.n11 VTAIL.n10 0.470328
R674 VTAIL.n3 VTAIL.n2 0.470328
R675 VTAIL VTAIL.n1 0.0586897
R676 VDD1 VDD1.n0 635.404
R677 VDD1.n3 VDD1.n2 635.292
R678 VDD1.n3 VDD1.n1 635.292
R679 VDD1.n5 VDD1.n4 634.639
R680 VDD1.n4 VDD1.t4 50.7896
R681 VDD1.n4 VDD1.t6 50.7896
R682 VDD1.n0 VDD1.t2 50.7896
R683 VDD1.n0 VDD1.t3 50.7896
R684 VDD1.n2 VDD1.t5 50.7896
R685 VDD1.n2 VDD1.t1 50.7896
R686 VDD1.n1 VDD1.t0 50.7896
R687 VDD1.n1 VDD1.t7 50.7896
R688 VDD1.n5 VDD1.n3 31.2121
R689 VDD1 VDD1.n5 0.649207
R690 VN.n18 VN.n17 175.419
R691 VN.n37 VN.n36 175.419
R692 VN.n35 VN.n19 161.3
R693 VN.n34 VN.n33 161.3
R694 VN.n32 VN.n20 161.3
R695 VN.n31 VN.n30 161.3
R696 VN.n29 VN.n21 161.3
R697 VN.n28 VN.n27 161.3
R698 VN.n26 VN.n23 161.3
R699 VN.n16 VN.n0 161.3
R700 VN.n15 VN.n14 161.3
R701 VN.n13 VN.n1 161.3
R702 VN.n12 VN.n11 161.3
R703 VN.n9 VN.n2 161.3
R704 VN.n8 VN.n7 161.3
R705 VN.n6 VN.n3 161.3
R706 VN.n5 VN.n4 61.8956
R707 VN.n25 VN.n24 61.8956
R708 VN.n9 VN.n8 56.4773
R709 VN.n29 VN.n28 56.4773
R710 VN.n15 VN.n1 51.1217
R711 VN.n34 VN.n20 51.1217
R712 VN.n5 VN.t7 39.2192
R713 VN.n25 VN.t1 39.2192
R714 VN VN.n37 36.5175
R715 VN.n16 VN.n15 29.6995
R716 VN.n35 VN.n34 29.6995
R717 VN.n26 VN.n25 27.6663
R718 VN.n6 VN.n5 27.6663
R719 VN.n8 VN.n3 24.3439
R720 VN.n11 VN.n9 24.3439
R721 VN.n28 VN.n23 24.3439
R722 VN.n30 VN.n29 24.3439
R723 VN.n10 VN.n1 20.9359
R724 VN.n22 VN.n20 20.9359
R725 VN.n4 VN.t6 11.7745
R726 VN.n10 VN.t4 11.7745
R727 VN.n17 VN.t0 11.7745
R728 VN.n24 VN.t2 11.7745
R729 VN.n22 VN.t3 11.7745
R730 VN.n36 VN.t5 11.7745
R731 VN.n17 VN.n16 10.2247
R732 VN.n36 VN.n35 10.2247
R733 VN.n4 VN.n3 3.40858
R734 VN.n11 VN.n10 3.40858
R735 VN.n24 VN.n23 3.40858
R736 VN.n30 VN.n22 3.40858
R737 VN.n37 VN.n19 0.189894
R738 VN.n33 VN.n19 0.189894
R739 VN.n33 VN.n32 0.189894
R740 VN.n32 VN.n31 0.189894
R741 VN.n31 VN.n21 0.189894
R742 VN.n27 VN.n21 0.189894
R743 VN.n27 VN.n26 0.189894
R744 VN.n7 VN.n6 0.189894
R745 VN.n7 VN.n2 0.189894
R746 VN.n12 VN.n2 0.189894
R747 VN.n13 VN.n12 0.189894
R748 VN.n14 VN.n13 0.189894
R749 VN.n14 VN.n0 0.189894
R750 VN.n18 VN.n0 0.189894
R751 VN VN.n18 0.0516364
R752 VDD2.n2 VDD2.n1 635.292
R753 VDD2.n2 VDD2.n0 635.292
R754 VDD2 VDD2.n5 635.288
R755 VDD2.n4 VDD2.n3 634.639
R756 VDD2.n5 VDD2.t5 50.7896
R757 VDD2.n5 VDD2.t6 50.7896
R758 VDD2.n3 VDD2.t2 50.7896
R759 VDD2.n3 VDD2.t4 50.7896
R760 VDD2.n1 VDD2.t3 50.7896
R761 VDD2.n1 VDD2.t7 50.7896
R762 VDD2.n0 VDD2.t0 50.7896
R763 VDD2.n0 VDD2.t1 50.7896
R764 VDD2.n4 VDD2.n2 30.6291
R765 VDD2 VDD2.n4 0.765586
C0 VP VTAIL 1.51447f
C1 VP VN 3.99785f
C2 VTAIL VN 1.50037f
C3 VP VDD2 0.391417f
C4 VP w_n2610_n1096# 5.06157f
C5 VDD2 VTAIL 3.08736f
C6 VTAIL w_n2610_n1096# 1.34919f
C7 VP B 1.30921f
C8 VP VDD1 1.01976f
C9 VTAIL B 0.825735f
C10 VTAIL VDD1 3.04159f
C11 VN w_n2610_n1096# 4.7356f
C12 VDD2 VN 0.787808f
C13 VN B 0.755955f
C14 VDD1 VN 0.156658f
C15 VDD2 w_n2610_n1096# 1.2671f
C16 B w_n2610_n1096# 4.98528f
C17 VDD2 B 1.00544f
C18 VDD1 w_n2610_n1096# 1.20789f
C19 VDD2 VDD1 1.13138f
C20 VDD1 B 0.949385f
C21 VDD2 VSUBS 0.715795f
C22 VDD1 VSUBS 1.111634f
C23 VTAIL VSUBS 0.346701f
C24 VN VSUBS 4.65122f
C25 VP VSUBS 1.6774f
C26 B VSUBS 2.45563f
C27 w_n2610_n1096# VSUBS 37.0516f
C28 VDD2.t0 VSUBS 0.010844f
C29 VDD2.t1 VSUBS 0.010844f
C30 VDD2.n0 VSUBS 0.023976f
C31 VDD2.t3 VSUBS 0.010844f
C32 VDD2.t7 VSUBS 0.010844f
C33 VDD2.n1 VSUBS 0.023976f
C34 VDD2.n2 VSUBS 1.36064f
C35 VDD2.t2 VSUBS 0.010844f
C36 VDD2.t4 VSUBS 0.010844f
C37 VDD2.n3 VSUBS 0.023761f
C38 VDD2.n4 VSUBS 1.25057f
C39 VDD2.t5 VSUBS 0.010844f
C40 VDD2.t6 VSUBS 0.010844f
C41 VDD2.n5 VSUBS 0.023974f
C42 VN.n0 VSUBS 0.060057f
C43 VN.t0 VSUBS 0.066145f
C44 VN.n1 VSUBS 0.101807f
C45 VN.n2 VSUBS 0.060057f
C46 VN.n3 VSUBS 0.064727f
C47 VN.t7 VSUBS 0.271085f
C48 VN.t6 VSUBS 0.066145f
C49 VN.n4 VSUBS 0.183148f
C50 VN.n5 VSUBS 0.174105f
C51 VN.n6 VSUBS 0.315091f
C52 VN.n7 VSUBS 0.060057f
C53 VN.n8 VSUBS 0.088054f
C54 VN.n9 VSUBS 0.088054f
C55 VN.t4 VSUBS 0.066145f
C56 VN.n10 VSUBS 0.102578f
C57 VN.n11 VSUBS 0.064727f
C58 VN.n12 VSUBS 0.060057f
C59 VN.n13 VSUBS 0.060057f
C60 VN.n14 VSUBS 0.060057f
C61 VN.n15 VSUBS 0.058713f
C62 VN.n16 VSUBS 0.088091f
C63 VN.n17 VSUBS 0.20806f
C64 VN.n18 VSUBS 0.055775f
C65 VN.n19 VSUBS 0.060057f
C66 VN.t5 VSUBS 0.066145f
C67 VN.n20 VSUBS 0.101807f
C68 VN.n21 VSUBS 0.060057f
C69 VN.t3 VSUBS 0.066145f
C70 VN.n22 VSUBS 0.102578f
C71 VN.n23 VSUBS 0.064727f
C72 VN.t1 VSUBS 0.271085f
C73 VN.t2 VSUBS 0.066145f
C74 VN.n24 VSUBS 0.183148f
C75 VN.n25 VSUBS 0.174105f
C76 VN.n26 VSUBS 0.315091f
C77 VN.n27 VSUBS 0.060057f
C78 VN.n28 VSUBS 0.088054f
C79 VN.n29 VSUBS 0.088054f
C80 VN.n30 VSUBS 0.064727f
C81 VN.n31 VSUBS 0.060057f
C82 VN.n32 VSUBS 0.060057f
C83 VN.n33 VSUBS 0.060057f
C84 VN.n34 VSUBS 0.058713f
C85 VN.n35 VSUBS 0.088091f
C86 VN.n36 VSUBS 0.20806f
C87 VN.n37 VSUBS 1.95081f
C88 VDD1.t2 VSUBS 0.010233f
C89 VDD1.t3 VSUBS 0.010233f
C90 VDD1.n0 VSUBS 0.022668f
C91 VDD1.t0 VSUBS 0.010233f
C92 VDD1.t7 VSUBS 0.010233f
C93 VDD1.n1 VSUBS 0.022625f
C94 VDD1.t5 VSUBS 0.010233f
C95 VDD1.t1 VSUBS 0.010233f
C96 VDD1.n2 VSUBS 0.022625f
C97 VDD1.n3 VSUBS 1.32689f
C98 VDD1.t4 VSUBS 0.010233f
C99 VDD1.t6 VSUBS 0.010233f
C100 VDD1.n4 VSUBS 0.022422f
C101 VDD1.n5 VSUBS 1.20428f
C102 VTAIL.t5 VSUBS 0.015197f
C103 VTAIL.t2 VSUBS 0.015197f
C104 VTAIL.n0 VSUBS 0.03127f
C105 VTAIL.n1 VSUBS 0.18464f
C106 VTAIL.t1 VSUBS 0.068349f
C107 VTAIL.n2 VSUBS 0.228865f
C108 VTAIL.t13 VSUBS 0.068349f
C109 VTAIL.n3 VSUBS 0.228865f
C110 VTAIL.t10 VSUBS 0.015197f
C111 VTAIL.t9 VSUBS 0.015197f
C112 VTAIL.n4 VSUBS 0.03127f
C113 VTAIL.n5 VSUBS 0.315898f
C114 VTAIL.t12 VSUBS 0.068349f
C115 VTAIL.n6 VSUBS 0.781875f
C116 VTAIL.t3 VSUBS 0.068349f
C117 VTAIL.n7 VSUBS 0.781875f
C118 VTAIL.t6 VSUBS 0.015197f
C119 VTAIL.t4 VSUBS 0.015197f
C120 VTAIL.n8 VSUBS 0.03127f
C121 VTAIL.n9 VSUBS 0.315898f
C122 VTAIL.t0 VSUBS 0.068349f
C123 VTAIL.n10 VSUBS 0.228865f
C124 VTAIL.t14 VSUBS 0.068349f
C125 VTAIL.n11 VSUBS 0.228865f
C126 VTAIL.t11 VSUBS 0.015197f
C127 VTAIL.t15 VSUBS 0.015197f
C128 VTAIL.n12 VSUBS 0.03127f
C129 VTAIL.n13 VSUBS 0.315898f
C130 VTAIL.t8 VSUBS 0.068349f
C131 VTAIL.n14 VSUBS 0.781875f
C132 VTAIL.t7 VSUBS 0.068349f
C133 VTAIL.n15 VSUBS 0.776241f
C134 VP.n0 VSUBS 0.063434f
C135 VP.t6 VSUBS 0.069864f
C136 VP.n1 VSUBS 0.107532f
C137 VP.n2 VSUBS 0.063434f
C138 VP.n3 VSUBS 0.068366f
C139 VP.n4 VSUBS 0.063434f
C140 VP.t7 VSUBS 0.069864f
C141 VP.n5 VSUBS 0.219758f
C142 VP.n6 VSUBS 0.063434f
C143 VP.t1 VSUBS 0.069864f
C144 VP.n7 VSUBS 0.107532f
C145 VP.n8 VSUBS 0.063434f
C146 VP.n9 VSUBS 0.068366f
C147 VP.t5 VSUBS 0.286327f
C148 VP.t4 VSUBS 0.069864f
C149 VP.n10 VSUBS 0.193446f
C150 VP.n11 VSUBS 0.183895f
C151 VP.n12 VSUBS 0.332807f
C152 VP.n13 VSUBS 0.063434f
C153 VP.n14 VSUBS 0.093005f
C154 VP.n15 VSUBS 0.093005f
C155 VP.t3 VSUBS 0.069864f
C156 VP.n16 VSUBS 0.108346f
C157 VP.n17 VSUBS 0.068366f
C158 VP.n18 VSUBS 0.063434f
C159 VP.n19 VSUBS 0.063434f
C160 VP.n20 VSUBS 0.063434f
C161 VP.n21 VSUBS 0.062014f
C162 VP.n22 VSUBS 0.093044f
C163 VP.n23 VSUBS 0.219758f
C164 VP.n24 VSUBS 2.01843f
C165 VP.n25 VSUBS 2.08135f
C166 VP.n26 VSUBS 0.063434f
C167 VP.n27 VSUBS 0.093044f
C168 VP.n28 VSUBS 0.062014f
C169 VP.t0 VSUBS 0.069864f
C170 VP.n29 VSUBS 0.108346f
C171 VP.n30 VSUBS 0.107532f
C172 VP.n31 VSUBS 0.063434f
C173 VP.n32 VSUBS 0.063434f
C174 VP.n33 VSUBS 0.063434f
C175 VP.n34 VSUBS 0.093005f
C176 VP.n35 VSUBS 0.093005f
C177 VP.t2 VSUBS 0.069864f
C178 VP.n36 VSUBS 0.108346f
C179 VP.n37 VSUBS 0.068366f
C180 VP.n38 VSUBS 0.063434f
C181 VP.n39 VSUBS 0.063434f
C182 VP.n40 VSUBS 0.063434f
C183 VP.n41 VSUBS 0.062014f
C184 VP.n42 VSUBS 0.093044f
C185 VP.n43 VSUBS 0.219758f
C186 VP.n44 VSUBS 0.058911f
C187 B.n0 VSUBS 0.006602f
C188 B.n1 VSUBS 0.006602f
C189 B.n2 VSUBS 0.01044f
C190 B.n3 VSUBS 0.01044f
C191 B.n4 VSUBS 0.01044f
C192 B.n5 VSUBS 0.01044f
C193 B.n6 VSUBS 0.01044f
C194 B.n7 VSUBS 0.01044f
C195 B.n8 VSUBS 0.01044f
C196 B.n9 VSUBS 0.01044f
C197 B.n10 VSUBS 0.01044f
C198 B.n11 VSUBS 0.01044f
C199 B.n12 VSUBS 0.01044f
C200 B.n13 VSUBS 0.01044f
C201 B.n14 VSUBS 0.01044f
C202 B.n15 VSUBS 0.01044f
C203 B.n16 VSUBS 0.01044f
C204 B.n17 VSUBS 0.01044f
C205 B.n18 VSUBS 0.026262f
C206 B.n19 VSUBS 0.01044f
C207 B.n20 VSUBS 0.01044f
C208 B.n21 VSUBS 0.01044f
C209 B.t2 VSUBS 0.018064f
C210 B.t1 VSUBS 0.019768f
C211 B.t0 VSUBS 0.066891f
C212 B.n22 VSUBS 0.05957f
C213 B.n23 VSUBS 0.051849f
C214 B.n24 VSUBS 0.024188f
C215 B.n25 VSUBS 0.01044f
C216 B.n26 VSUBS 0.01044f
C217 B.n27 VSUBS 0.01044f
C218 B.n28 VSUBS 0.01044f
C219 B.n29 VSUBS 0.01044f
C220 B.t5 VSUBS 0.018064f
C221 B.t4 VSUBS 0.019768f
C222 B.t3 VSUBS 0.06692f
C223 B.n30 VSUBS 0.059541f
C224 B.n31 VSUBS 0.051849f
C225 B.n32 VSUBS 0.01044f
C226 B.n33 VSUBS 0.01044f
C227 B.n34 VSUBS 0.01044f
C228 B.n35 VSUBS 0.026262f
C229 B.n36 VSUBS 0.01044f
C230 B.n37 VSUBS 0.01044f
C231 B.n38 VSUBS 0.01044f
C232 B.n39 VSUBS 0.01044f
C233 B.n40 VSUBS 0.01044f
C234 B.n41 VSUBS 0.01044f
C235 B.n42 VSUBS 0.01044f
C236 B.n43 VSUBS 0.01044f
C237 B.n44 VSUBS 0.01044f
C238 B.n45 VSUBS 0.01044f
C239 B.n46 VSUBS 0.01044f
C240 B.n47 VSUBS 0.01044f
C241 B.n48 VSUBS 0.01044f
C242 B.n49 VSUBS 0.01044f
C243 B.n50 VSUBS 0.01044f
C244 B.n51 VSUBS 0.01044f
C245 B.n52 VSUBS 0.01044f
C246 B.n53 VSUBS 0.01044f
C247 B.n54 VSUBS 0.01044f
C248 B.n55 VSUBS 0.01044f
C249 B.n56 VSUBS 0.01044f
C250 B.n57 VSUBS 0.01044f
C251 B.n58 VSUBS 0.01044f
C252 B.n59 VSUBS 0.01044f
C253 B.n60 VSUBS 0.01044f
C254 B.n61 VSUBS 0.01044f
C255 B.n62 VSUBS 0.01044f
C256 B.n63 VSUBS 0.01044f
C257 B.n64 VSUBS 0.01044f
C258 B.n65 VSUBS 0.01044f
C259 B.n66 VSUBS 0.01044f
C260 B.n67 VSUBS 0.01044f
C261 B.n68 VSUBS 0.026262f
C262 B.n69 VSUBS 0.01044f
C263 B.n70 VSUBS 0.01044f
C264 B.n71 VSUBS 0.01044f
C265 B.t10 VSUBS 0.018064f
C266 B.t11 VSUBS 0.019768f
C267 B.t9 VSUBS 0.06692f
C268 B.n72 VSUBS 0.059541f
C269 B.n73 VSUBS 0.051849f
C270 B.n74 VSUBS 0.024188f
C271 B.n75 VSUBS 0.01044f
C272 B.n76 VSUBS 0.01044f
C273 B.n77 VSUBS 0.01044f
C274 B.n78 VSUBS 0.01044f
C275 B.n79 VSUBS 0.01044f
C276 B.t7 VSUBS 0.018064f
C277 B.t8 VSUBS 0.019768f
C278 B.t6 VSUBS 0.066891f
C279 B.n80 VSUBS 0.05957f
C280 B.n81 VSUBS 0.051849f
C281 B.n82 VSUBS 0.01044f
C282 B.n83 VSUBS 0.01044f
C283 B.n84 VSUBS 0.01044f
C284 B.n85 VSUBS 0.026262f
C285 B.n86 VSUBS 0.01044f
C286 B.n87 VSUBS 0.01044f
C287 B.n88 VSUBS 0.01044f
C288 B.n89 VSUBS 0.01044f
C289 B.n90 VSUBS 0.01044f
C290 B.n91 VSUBS 0.01044f
C291 B.n92 VSUBS 0.01044f
C292 B.n93 VSUBS 0.01044f
C293 B.n94 VSUBS 0.01044f
C294 B.n95 VSUBS 0.01044f
C295 B.n96 VSUBS 0.01044f
C296 B.n97 VSUBS 0.01044f
C297 B.n98 VSUBS 0.01044f
C298 B.n99 VSUBS 0.01044f
C299 B.n100 VSUBS 0.01044f
C300 B.n101 VSUBS 0.01044f
C301 B.n102 VSUBS 0.01044f
C302 B.n103 VSUBS 0.01044f
C303 B.n104 VSUBS 0.01044f
C304 B.n105 VSUBS 0.01044f
C305 B.n106 VSUBS 0.01044f
C306 B.n107 VSUBS 0.01044f
C307 B.n108 VSUBS 0.01044f
C308 B.n109 VSUBS 0.01044f
C309 B.n110 VSUBS 0.01044f
C310 B.n111 VSUBS 0.01044f
C311 B.n112 VSUBS 0.01044f
C312 B.n113 VSUBS 0.01044f
C313 B.n114 VSUBS 0.01044f
C314 B.n115 VSUBS 0.01044f
C315 B.n116 VSUBS 0.01044f
C316 B.n117 VSUBS 0.01044f
C317 B.n118 VSUBS 0.01044f
C318 B.n119 VSUBS 0.01044f
C319 B.n120 VSUBS 0.01044f
C320 B.n121 VSUBS 0.01044f
C321 B.n122 VSUBS 0.01044f
C322 B.n123 VSUBS 0.01044f
C323 B.n124 VSUBS 0.01044f
C324 B.n125 VSUBS 0.01044f
C325 B.n126 VSUBS 0.01044f
C326 B.n127 VSUBS 0.01044f
C327 B.n128 VSUBS 0.01044f
C328 B.n129 VSUBS 0.01044f
C329 B.n130 VSUBS 0.01044f
C330 B.n131 VSUBS 0.01044f
C331 B.n132 VSUBS 0.01044f
C332 B.n133 VSUBS 0.01044f
C333 B.n134 VSUBS 0.01044f
C334 B.n135 VSUBS 0.01044f
C335 B.n136 VSUBS 0.01044f
C336 B.n137 VSUBS 0.01044f
C337 B.n138 VSUBS 0.01044f
C338 B.n139 VSUBS 0.01044f
C339 B.n140 VSUBS 0.01044f
C340 B.n141 VSUBS 0.01044f
C341 B.n142 VSUBS 0.01044f
C342 B.n143 VSUBS 0.01044f
C343 B.n144 VSUBS 0.01044f
C344 B.n145 VSUBS 0.01044f
C345 B.n146 VSUBS 0.024709f
C346 B.n147 VSUBS 0.024709f
C347 B.n148 VSUBS 0.026262f
C348 B.n149 VSUBS 0.01044f
C349 B.n150 VSUBS 0.01044f
C350 B.n151 VSUBS 0.01044f
C351 B.n152 VSUBS 0.01044f
C352 B.n153 VSUBS 0.01044f
C353 B.n154 VSUBS 0.01044f
C354 B.n155 VSUBS 0.01044f
C355 B.n156 VSUBS 0.01044f
C356 B.n157 VSUBS 0.01044f
C357 B.n158 VSUBS 0.01044f
C358 B.n159 VSUBS 0.009903f
C359 B.n160 VSUBS 0.024188f
C360 B.n161 VSUBS 0.005757f
C361 B.n162 VSUBS 0.01044f
C362 B.n163 VSUBS 0.01044f
C363 B.n164 VSUBS 0.01044f
C364 B.n165 VSUBS 0.01044f
C365 B.n166 VSUBS 0.01044f
C366 B.n167 VSUBS 0.01044f
C367 B.n168 VSUBS 0.01044f
C368 B.n169 VSUBS 0.01044f
C369 B.n170 VSUBS 0.01044f
C370 B.n171 VSUBS 0.01044f
C371 B.n172 VSUBS 0.01044f
C372 B.n173 VSUBS 0.01044f
C373 B.n174 VSUBS 0.005757f
C374 B.n175 VSUBS 0.01044f
C375 B.n176 VSUBS 0.01044f
C376 B.n177 VSUBS 0.009903f
C377 B.n178 VSUBS 0.01044f
C378 B.n179 VSUBS 0.01044f
C379 B.n180 VSUBS 0.01044f
C380 B.n181 VSUBS 0.01044f
C381 B.n182 VSUBS 0.01044f
C382 B.n183 VSUBS 0.01044f
C383 B.n184 VSUBS 0.01044f
C384 B.n185 VSUBS 0.01044f
C385 B.n186 VSUBS 0.01044f
C386 B.n187 VSUBS 0.026262f
C387 B.n188 VSUBS 0.024709f
C388 B.n189 VSUBS 0.024709f
C389 B.n190 VSUBS 0.01044f
C390 B.n191 VSUBS 0.01044f
C391 B.n192 VSUBS 0.01044f
C392 B.n193 VSUBS 0.01044f
C393 B.n194 VSUBS 0.01044f
C394 B.n195 VSUBS 0.01044f
C395 B.n196 VSUBS 0.01044f
C396 B.n197 VSUBS 0.01044f
C397 B.n198 VSUBS 0.01044f
C398 B.n199 VSUBS 0.01044f
C399 B.n200 VSUBS 0.01044f
C400 B.n201 VSUBS 0.01044f
C401 B.n202 VSUBS 0.01044f
C402 B.n203 VSUBS 0.01044f
C403 B.n204 VSUBS 0.01044f
C404 B.n205 VSUBS 0.01044f
C405 B.n206 VSUBS 0.01044f
C406 B.n207 VSUBS 0.01044f
C407 B.n208 VSUBS 0.01044f
C408 B.n209 VSUBS 0.01044f
C409 B.n210 VSUBS 0.01044f
C410 B.n211 VSUBS 0.01044f
C411 B.n212 VSUBS 0.01044f
C412 B.n213 VSUBS 0.01044f
C413 B.n214 VSUBS 0.01044f
C414 B.n215 VSUBS 0.01044f
C415 B.n216 VSUBS 0.01044f
C416 B.n217 VSUBS 0.01044f
C417 B.n218 VSUBS 0.01044f
C418 B.n219 VSUBS 0.01044f
C419 B.n220 VSUBS 0.01044f
C420 B.n221 VSUBS 0.01044f
C421 B.n222 VSUBS 0.01044f
C422 B.n223 VSUBS 0.01044f
C423 B.n224 VSUBS 0.01044f
C424 B.n225 VSUBS 0.01044f
C425 B.n226 VSUBS 0.01044f
C426 B.n227 VSUBS 0.01044f
C427 B.n228 VSUBS 0.01044f
C428 B.n229 VSUBS 0.01044f
C429 B.n230 VSUBS 0.01044f
C430 B.n231 VSUBS 0.01044f
C431 B.n232 VSUBS 0.01044f
C432 B.n233 VSUBS 0.01044f
C433 B.n234 VSUBS 0.01044f
C434 B.n235 VSUBS 0.01044f
C435 B.n236 VSUBS 0.01044f
C436 B.n237 VSUBS 0.01044f
C437 B.n238 VSUBS 0.01044f
C438 B.n239 VSUBS 0.01044f
C439 B.n240 VSUBS 0.01044f
C440 B.n241 VSUBS 0.01044f
C441 B.n242 VSUBS 0.01044f
C442 B.n243 VSUBS 0.01044f
C443 B.n244 VSUBS 0.01044f
C444 B.n245 VSUBS 0.01044f
C445 B.n246 VSUBS 0.01044f
C446 B.n247 VSUBS 0.01044f
C447 B.n248 VSUBS 0.01044f
C448 B.n249 VSUBS 0.01044f
C449 B.n250 VSUBS 0.01044f
C450 B.n251 VSUBS 0.01044f
C451 B.n252 VSUBS 0.01044f
C452 B.n253 VSUBS 0.01044f
C453 B.n254 VSUBS 0.01044f
C454 B.n255 VSUBS 0.01044f
C455 B.n256 VSUBS 0.01044f
C456 B.n257 VSUBS 0.01044f
C457 B.n258 VSUBS 0.01044f
C458 B.n259 VSUBS 0.01044f
C459 B.n260 VSUBS 0.01044f
C460 B.n261 VSUBS 0.01044f
C461 B.n262 VSUBS 0.01044f
C462 B.n263 VSUBS 0.01044f
C463 B.n264 VSUBS 0.01044f
C464 B.n265 VSUBS 0.01044f
C465 B.n266 VSUBS 0.01044f
C466 B.n267 VSUBS 0.01044f
C467 B.n268 VSUBS 0.01044f
C468 B.n269 VSUBS 0.01044f
C469 B.n270 VSUBS 0.01044f
C470 B.n271 VSUBS 0.01044f
C471 B.n272 VSUBS 0.01044f
C472 B.n273 VSUBS 0.01044f
C473 B.n274 VSUBS 0.01044f
C474 B.n275 VSUBS 0.01044f
C475 B.n276 VSUBS 0.01044f
C476 B.n277 VSUBS 0.01044f
C477 B.n278 VSUBS 0.01044f
C478 B.n279 VSUBS 0.01044f
C479 B.n280 VSUBS 0.01044f
C480 B.n281 VSUBS 0.01044f
C481 B.n282 VSUBS 0.01044f
C482 B.n283 VSUBS 0.01044f
C483 B.n284 VSUBS 0.024709f
C484 B.n285 VSUBS 0.025867f
C485 B.n286 VSUBS 0.025105f
C486 B.n287 VSUBS 0.01044f
C487 B.n288 VSUBS 0.01044f
C488 B.n289 VSUBS 0.01044f
C489 B.n290 VSUBS 0.01044f
C490 B.n291 VSUBS 0.01044f
C491 B.n292 VSUBS 0.01044f
C492 B.n293 VSUBS 0.01044f
C493 B.n294 VSUBS 0.01044f
C494 B.n295 VSUBS 0.01044f
C495 B.n296 VSUBS 0.01044f
C496 B.n297 VSUBS 0.009903f
C497 B.n298 VSUBS 0.024188f
C498 B.n299 VSUBS 0.005757f
C499 B.n300 VSUBS 0.01044f
C500 B.n301 VSUBS 0.01044f
C501 B.n302 VSUBS 0.01044f
C502 B.n303 VSUBS 0.01044f
C503 B.n304 VSUBS 0.01044f
C504 B.n305 VSUBS 0.01044f
C505 B.n306 VSUBS 0.01044f
C506 B.n307 VSUBS 0.01044f
C507 B.n308 VSUBS 0.01044f
C508 B.n309 VSUBS 0.01044f
C509 B.n310 VSUBS 0.01044f
C510 B.n311 VSUBS 0.01044f
C511 B.n312 VSUBS 0.005757f
C512 B.n313 VSUBS 0.01044f
C513 B.n314 VSUBS 0.01044f
C514 B.n315 VSUBS 0.009903f
C515 B.n316 VSUBS 0.01044f
C516 B.n317 VSUBS 0.01044f
C517 B.n318 VSUBS 0.01044f
C518 B.n319 VSUBS 0.01044f
C519 B.n320 VSUBS 0.01044f
C520 B.n321 VSUBS 0.01044f
C521 B.n322 VSUBS 0.01044f
C522 B.n323 VSUBS 0.01044f
C523 B.n324 VSUBS 0.01044f
C524 B.n325 VSUBS 0.026262f
C525 B.n326 VSUBS 0.024709f
C526 B.n327 VSUBS 0.024709f
C527 B.n328 VSUBS 0.01044f
C528 B.n329 VSUBS 0.01044f
C529 B.n330 VSUBS 0.01044f
C530 B.n331 VSUBS 0.01044f
C531 B.n332 VSUBS 0.01044f
C532 B.n333 VSUBS 0.01044f
C533 B.n334 VSUBS 0.01044f
C534 B.n335 VSUBS 0.01044f
C535 B.n336 VSUBS 0.01044f
C536 B.n337 VSUBS 0.01044f
C537 B.n338 VSUBS 0.01044f
C538 B.n339 VSUBS 0.01044f
C539 B.n340 VSUBS 0.01044f
C540 B.n341 VSUBS 0.01044f
C541 B.n342 VSUBS 0.01044f
C542 B.n343 VSUBS 0.01044f
C543 B.n344 VSUBS 0.01044f
C544 B.n345 VSUBS 0.01044f
C545 B.n346 VSUBS 0.01044f
C546 B.n347 VSUBS 0.01044f
C547 B.n348 VSUBS 0.01044f
C548 B.n349 VSUBS 0.01044f
C549 B.n350 VSUBS 0.01044f
C550 B.n351 VSUBS 0.01044f
C551 B.n352 VSUBS 0.01044f
C552 B.n353 VSUBS 0.01044f
C553 B.n354 VSUBS 0.01044f
C554 B.n355 VSUBS 0.01044f
C555 B.n356 VSUBS 0.01044f
C556 B.n357 VSUBS 0.01044f
C557 B.n358 VSUBS 0.01044f
C558 B.n359 VSUBS 0.01044f
C559 B.n360 VSUBS 0.01044f
C560 B.n361 VSUBS 0.01044f
C561 B.n362 VSUBS 0.01044f
C562 B.n363 VSUBS 0.01044f
C563 B.n364 VSUBS 0.01044f
C564 B.n365 VSUBS 0.01044f
C565 B.n366 VSUBS 0.01044f
C566 B.n367 VSUBS 0.01044f
C567 B.n368 VSUBS 0.01044f
C568 B.n369 VSUBS 0.01044f
C569 B.n370 VSUBS 0.01044f
C570 B.n371 VSUBS 0.01044f
C571 B.n372 VSUBS 0.01044f
C572 B.n373 VSUBS 0.01044f
C573 B.n374 VSUBS 0.01044f
C574 B.n375 VSUBS 0.02364f
.ends

