* NGSPICE file created from diff_pair_sample_0453.ext - technology: sky130A

.subckt diff_pair_sample_0453 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=0 ps=0 w=3.59 l=1.19
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=0 ps=0 w=3.59 l=1.19
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=1.4001 ps=7.96 w=3.59 l=1.19
X3 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=1.4001 ps=7.96 w=3.59 l=1.19
X4 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=1.4001 ps=7.96 w=3.59 l=1.19
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=1.4001 ps=7.96 w=3.59 l=1.19
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=0 ps=0 w=3.59 l=1.19
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4001 pd=7.96 as=0 ps=0 w=3.59 l=1.19
R0 B.n365 B.n364 585
R1 B.n366 B.n365 585
R2 B.n145 B.n56 585
R3 B.n144 B.n143 585
R4 B.n142 B.n141 585
R5 B.n140 B.n139 585
R6 B.n138 B.n137 585
R7 B.n136 B.n135 585
R8 B.n134 B.n133 585
R9 B.n132 B.n131 585
R10 B.n130 B.n129 585
R11 B.n128 B.n127 585
R12 B.n126 B.n125 585
R13 B.n124 B.n123 585
R14 B.n122 B.n121 585
R15 B.n120 B.n119 585
R16 B.n118 B.n117 585
R17 B.n116 B.n115 585
R18 B.n114 B.n113 585
R19 B.n112 B.n111 585
R20 B.n110 B.n109 585
R21 B.n108 B.n107 585
R22 B.n106 B.n105 585
R23 B.n104 B.n103 585
R24 B.n102 B.n101 585
R25 B.n100 B.n99 585
R26 B.n98 B.n97 585
R27 B.n95 B.n94 585
R28 B.n93 B.n92 585
R29 B.n91 B.n90 585
R30 B.n89 B.n88 585
R31 B.n87 B.n86 585
R32 B.n85 B.n84 585
R33 B.n83 B.n82 585
R34 B.n81 B.n80 585
R35 B.n79 B.n78 585
R36 B.n77 B.n76 585
R37 B.n75 B.n74 585
R38 B.n73 B.n72 585
R39 B.n71 B.n70 585
R40 B.n69 B.n68 585
R41 B.n67 B.n66 585
R42 B.n65 B.n64 585
R43 B.n63 B.n62 585
R44 B.n363 B.n34 585
R45 B.n367 B.n34 585
R46 B.n362 B.n33 585
R47 B.n368 B.n33 585
R48 B.n361 B.n360 585
R49 B.n360 B.n29 585
R50 B.n359 B.n28 585
R51 B.n374 B.n28 585
R52 B.n358 B.n27 585
R53 B.n375 B.n27 585
R54 B.n357 B.n26 585
R55 B.n376 B.n26 585
R56 B.n356 B.n355 585
R57 B.n355 B.n22 585
R58 B.n354 B.n21 585
R59 B.n382 B.n21 585
R60 B.n353 B.n20 585
R61 B.n383 B.n20 585
R62 B.n352 B.n19 585
R63 B.n384 B.n19 585
R64 B.n351 B.n350 585
R65 B.n350 B.n15 585
R66 B.n349 B.n14 585
R67 B.n390 B.n14 585
R68 B.n348 B.n13 585
R69 B.n391 B.n13 585
R70 B.n347 B.n12 585
R71 B.n392 B.n12 585
R72 B.n346 B.n345 585
R73 B.n345 B.n8 585
R74 B.n344 B.n7 585
R75 B.n398 B.n7 585
R76 B.n343 B.n6 585
R77 B.n399 B.n6 585
R78 B.n342 B.n5 585
R79 B.n400 B.n5 585
R80 B.n341 B.n340 585
R81 B.n340 B.n4 585
R82 B.n339 B.n146 585
R83 B.n339 B.n338 585
R84 B.n329 B.n147 585
R85 B.n148 B.n147 585
R86 B.n331 B.n330 585
R87 B.n332 B.n331 585
R88 B.n328 B.n153 585
R89 B.n153 B.n152 585
R90 B.n327 B.n326 585
R91 B.n326 B.n325 585
R92 B.n155 B.n154 585
R93 B.n156 B.n155 585
R94 B.n318 B.n317 585
R95 B.n319 B.n318 585
R96 B.n316 B.n161 585
R97 B.n161 B.n160 585
R98 B.n315 B.n314 585
R99 B.n314 B.n313 585
R100 B.n163 B.n162 585
R101 B.n164 B.n163 585
R102 B.n306 B.n305 585
R103 B.n307 B.n306 585
R104 B.n304 B.n169 585
R105 B.n169 B.n168 585
R106 B.n303 B.n302 585
R107 B.n302 B.n301 585
R108 B.n171 B.n170 585
R109 B.n172 B.n171 585
R110 B.n294 B.n293 585
R111 B.n295 B.n294 585
R112 B.n292 B.n177 585
R113 B.n177 B.n176 585
R114 B.n286 B.n285 585
R115 B.n284 B.n200 585
R116 B.n283 B.n199 585
R117 B.n288 B.n199 585
R118 B.n282 B.n281 585
R119 B.n280 B.n279 585
R120 B.n278 B.n277 585
R121 B.n276 B.n275 585
R122 B.n274 B.n273 585
R123 B.n272 B.n271 585
R124 B.n270 B.n269 585
R125 B.n268 B.n267 585
R126 B.n266 B.n265 585
R127 B.n264 B.n263 585
R128 B.n262 B.n261 585
R129 B.n260 B.n259 585
R130 B.n258 B.n257 585
R131 B.n256 B.n255 585
R132 B.n254 B.n253 585
R133 B.n252 B.n251 585
R134 B.n250 B.n249 585
R135 B.n248 B.n247 585
R136 B.n246 B.n245 585
R137 B.n244 B.n243 585
R138 B.n242 B.n241 585
R139 B.n240 B.n239 585
R140 B.n238 B.n237 585
R141 B.n235 B.n234 585
R142 B.n233 B.n232 585
R143 B.n231 B.n230 585
R144 B.n229 B.n228 585
R145 B.n227 B.n226 585
R146 B.n225 B.n224 585
R147 B.n223 B.n222 585
R148 B.n221 B.n220 585
R149 B.n219 B.n218 585
R150 B.n217 B.n216 585
R151 B.n215 B.n214 585
R152 B.n213 B.n212 585
R153 B.n211 B.n210 585
R154 B.n209 B.n208 585
R155 B.n207 B.n206 585
R156 B.n179 B.n178 585
R157 B.n291 B.n290 585
R158 B.n175 B.n174 585
R159 B.n176 B.n175 585
R160 B.n297 B.n296 585
R161 B.n296 B.n295 585
R162 B.n298 B.n173 585
R163 B.n173 B.n172 585
R164 B.n300 B.n299 585
R165 B.n301 B.n300 585
R166 B.n167 B.n166 585
R167 B.n168 B.n167 585
R168 B.n309 B.n308 585
R169 B.n308 B.n307 585
R170 B.n310 B.n165 585
R171 B.n165 B.n164 585
R172 B.n312 B.n311 585
R173 B.n313 B.n312 585
R174 B.n159 B.n158 585
R175 B.n160 B.n159 585
R176 B.n321 B.n320 585
R177 B.n320 B.n319 585
R178 B.n322 B.n157 585
R179 B.n157 B.n156 585
R180 B.n324 B.n323 585
R181 B.n325 B.n324 585
R182 B.n151 B.n150 585
R183 B.n152 B.n151 585
R184 B.n334 B.n333 585
R185 B.n333 B.n332 585
R186 B.n335 B.n149 585
R187 B.n149 B.n148 585
R188 B.n337 B.n336 585
R189 B.n338 B.n337 585
R190 B.n2 B.n0 585
R191 B.n4 B.n2 585
R192 B.n3 B.n1 585
R193 B.n399 B.n3 585
R194 B.n397 B.n396 585
R195 B.n398 B.n397 585
R196 B.n395 B.n9 585
R197 B.n9 B.n8 585
R198 B.n394 B.n393 585
R199 B.n393 B.n392 585
R200 B.n11 B.n10 585
R201 B.n391 B.n11 585
R202 B.n389 B.n388 585
R203 B.n390 B.n389 585
R204 B.n387 B.n16 585
R205 B.n16 B.n15 585
R206 B.n386 B.n385 585
R207 B.n385 B.n384 585
R208 B.n18 B.n17 585
R209 B.n383 B.n18 585
R210 B.n381 B.n380 585
R211 B.n382 B.n381 585
R212 B.n379 B.n23 585
R213 B.n23 B.n22 585
R214 B.n378 B.n377 585
R215 B.n377 B.n376 585
R216 B.n25 B.n24 585
R217 B.n375 B.n25 585
R218 B.n373 B.n372 585
R219 B.n374 B.n373 585
R220 B.n371 B.n30 585
R221 B.n30 B.n29 585
R222 B.n370 B.n369 585
R223 B.n369 B.n368 585
R224 B.n32 B.n31 585
R225 B.n367 B.n32 585
R226 B.n402 B.n401 585
R227 B.n401 B.n400 585
R228 B.n286 B.n175 535.745
R229 B.n62 B.n32 535.745
R230 B.n290 B.n177 535.745
R231 B.n365 B.n34 535.745
R232 B.n204 B.t2 276.769
R233 B.n201 B.t6 276.769
R234 B.n60 B.t9 276.769
R235 B.n57 B.t13 276.769
R236 B.n366 B.n55 256.663
R237 B.n366 B.n54 256.663
R238 B.n366 B.n53 256.663
R239 B.n366 B.n52 256.663
R240 B.n366 B.n51 256.663
R241 B.n366 B.n50 256.663
R242 B.n366 B.n49 256.663
R243 B.n366 B.n48 256.663
R244 B.n366 B.n47 256.663
R245 B.n366 B.n46 256.663
R246 B.n366 B.n45 256.663
R247 B.n366 B.n44 256.663
R248 B.n366 B.n43 256.663
R249 B.n366 B.n42 256.663
R250 B.n366 B.n41 256.663
R251 B.n366 B.n40 256.663
R252 B.n366 B.n39 256.663
R253 B.n366 B.n38 256.663
R254 B.n366 B.n37 256.663
R255 B.n366 B.n36 256.663
R256 B.n366 B.n35 256.663
R257 B.n288 B.n287 256.663
R258 B.n288 B.n180 256.663
R259 B.n288 B.n181 256.663
R260 B.n288 B.n182 256.663
R261 B.n288 B.n183 256.663
R262 B.n288 B.n184 256.663
R263 B.n288 B.n185 256.663
R264 B.n288 B.n186 256.663
R265 B.n288 B.n187 256.663
R266 B.n288 B.n188 256.663
R267 B.n288 B.n189 256.663
R268 B.n288 B.n190 256.663
R269 B.n288 B.n191 256.663
R270 B.n288 B.n192 256.663
R271 B.n288 B.n193 256.663
R272 B.n288 B.n194 256.663
R273 B.n288 B.n195 256.663
R274 B.n288 B.n196 256.663
R275 B.n288 B.n197 256.663
R276 B.n288 B.n198 256.663
R277 B.n289 B.n288 256.663
R278 B.n296 B.n175 163.367
R279 B.n296 B.n173 163.367
R280 B.n300 B.n173 163.367
R281 B.n300 B.n167 163.367
R282 B.n308 B.n167 163.367
R283 B.n308 B.n165 163.367
R284 B.n312 B.n165 163.367
R285 B.n312 B.n159 163.367
R286 B.n320 B.n159 163.367
R287 B.n320 B.n157 163.367
R288 B.n324 B.n157 163.367
R289 B.n324 B.n151 163.367
R290 B.n333 B.n151 163.367
R291 B.n333 B.n149 163.367
R292 B.n337 B.n149 163.367
R293 B.n337 B.n2 163.367
R294 B.n401 B.n2 163.367
R295 B.n401 B.n3 163.367
R296 B.n397 B.n3 163.367
R297 B.n397 B.n9 163.367
R298 B.n393 B.n9 163.367
R299 B.n393 B.n11 163.367
R300 B.n389 B.n11 163.367
R301 B.n389 B.n16 163.367
R302 B.n385 B.n16 163.367
R303 B.n385 B.n18 163.367
R304 B.n381 B.n18 163.367
R305 B.n381 B.n23 163.367
R306 B.n377 B.n23 163.367
R307 B.n377 B.n25 163.367
R308 B.n373 B.n25 163.367
R309 B.n373 B.n30 163.367
R310 B.n369 B.n30 163.367
R311 B.n369 B.n32 163.367
R312 B.n200 B.n199 163.367
R313 B.n281 B.n199 163.367
R314 B.n279 B.n278 163.367
R315 B.n275 B.n274 163.367
R316 B.n271 B.n270 163.367
R317 B.n267 B.n266 163.367
R318 B.n263 B.n262 163.367
R319 B.n259 B.n258 163.367
R320 B.n255 B.n254 163.367
R321 B.n251 B.n250 163.367
R322 B.n247 B.n246 163.367
R323 B.n243 B.n242 163.367
R324 B.n239 B.n238 163.367
R325 B.n234 B.n233 163.367
R326 B.n230 B.n229 163.367
R327 B.n226 B.n225 163.367
R328 B.n222 B.n221 163.367
R329 B.n218 B.n217 163.367
R330 B.n214 B.n213 163.367
R331 B.n210 B.n209 163.367
R332 B.n206 B.n179 163.367
R333 B.n294 B.n177 163.367
R334 B.n294 B.n171 163.367
R335 B.n302 B.n171 163.367
R336 B.n302 B.n169 163.367
R337 B.n306 B.n169 163.367
R338 B.n306 B.n163 163.367
R339 B.n314 B.n163 163.367
R340 B.n314 B.n161 163.367
R341 B.n318 B.n161 163.367
R342 B.n318 B.n155 163.367
R343 B.n326 B.n155 163.367
R344 B.n326 B.n153 163.367
R345 B.n331 B.n153 163.367
R346 B.n331 B.n147 163.367
R347 B.n339 B.n147 163.367
R348 B.n340 B.n339 163.367
R349 B.n340 B.n5 163.367
R350 B.n6 B.n5 163.367
R351 B.n7 B.n6 163.367
R352 B.n345 B.n7 163.367
R353 B.n345 B.n12 163.367
R354 B.n13 B.n12 163.367
R355 B.n14 B.n13 163.367
R356 B.n350 B.n14 163.367
R357 B.n350 B.n19 163.367
R358 B.n20 B.n19 163.367
R359 B.n21 B.n20 163.367
R360 B.n355 B.n21 163.367
R361 B.n355 B.n26 163.367
R362 B.n27 B.n26 163.367
R363 B.n28 B.n27 163.367
R364 B.n360 B.n28 163.367
R365 B.n360 B.n33 163.367
R366 B.n34 B.n33 163.367
R367 B.n66 B.n65 163.367
R368 B.n70 B.n69 163.367
R369 B.n74 B.n73 163.367
R370 B.n78 B.n77 163.367
R371 B.n82 B.n81 163.367
R372 B.n86 B.n85 163.367
R373 B.n90 B.n89 163.367
R374 B.n94 B.n93 163.367
R375 B.n99 B.n98 163.367
R376 B.n103 B.n102 163.367
R377 B.n107 B.n106 163.367
R378 B.n111 B.n110 163.367
R379 B.n115 B.n114 163.367
R380 B.n119 B.n118 163.367
R381 B.n123 B.n122 163.367
R382 B.n127 B.n126 163.367
R383 B.n131 B.n130 163.367
R384 B.n135 B.n134 163.367
R385 B.n139 B.n138 163.367
R386 B.n143 B.n142 163.367
R387 B.n365 B.n56 163.367
R388 B.n288 B.n176 157.587
R389 B.n367 B.n366 157.587
R390 B.n204 B.t5 105.641
R391 B.n57 B.t14 105.641
R392 B.n201 B.t8 105.638
R393 B.n60 B.t11 105.638
R394 B.n295 B.n176 84.3773
R395 B.n295 B.n172 84.3773
R396 B.n301 B.n172 84.3773
R397 B.n301 B.n168 84.3773
R398 B.n307 B.n168 84.3773
R399 B.n313 B.n164 84.3773
R400 B.n313 B.n160 84.3773
R401 B.n319 B.n160 84.3773
R402 B.n319 B.n156 84.3773
R403 B.n325 B.n156 84.3773
R404 B.n325 B.n152 84.3773
R405 B.n332 B.n152 84.3773
R406 B.n338 B.n148 84.3773
R407 B.n338 B.n4 84.3773
R408 B.n400 B.n4 84.3773
R409 B.n400 B.n399 84.3773
R410 B.n399 B.n398 84.3773
R411 B.n398 B.n8 84.3773
R412 B.n392 B.n391 84.3773
R413 B.n391 B.n390 84.3773
R414 B.n390 B.n15 84.3773
R415 B.n384 B.n15 84.3773
R416 B.n384 B.n383 84.3773
R417 B.n383 B.n382 84.3773
R418 B.n382 B.n22 84.3773
R419 B.n376 B.n375 84.3773
R420 B.n375 B.n374 84.3773
R421 B.n374 B.n29 84.3773
R422 B.n368 B.n29 84.3773
R423 B.n368 B.n367 84.3773
R424 B.n205 B.t4 76.1617
R425 B.n58 B.t15 76.1617
R426 B.n202 B.t7 76.1588
R427 B.n61 B.t12 76.1588
R428 B.n287 B.n286 71.676
R429 B.n281 B.n180 71.676
R430 B.n278 B.n181 71.676
R431 B.n274 B.n182 71.676
R432 B.n270 B.n183 71.676
R433 B.n266 B.n184 71.676
R434 B.n262 B.n185 71.676
R435 B.n258 B.n186 71.676
R436 B.n254 B.n187 71.676
R437 B.n250 B.n188 71.676
R438 B.n246 B.n189 71.676
R439 B.n242 B.n190 71.676
R440 B.n238 B.n191 71.676
R441 B.n233 B.n192 71.676
R442 B.n229 B.n193 71.676
R443 B.n225 B.n194 71.676
R444 B.n221 B.n195 71.676
R445 B.n217 B.n196 71.676
R446 B.n213 B.n197 71.676
R447 B.n209 B.n198 71.676
R448 B.n289 B.n179 71.676
R449 B.n62 B.n35 71.676
R450 B.n66 B.n36 71.676
R451 B.n70 B.n37 71.676
R452 B.n74 B.n38 71.676
R453 B.n78 B.n39 71.676
R454 B.n82 B.n40 71.676
R455 B.n86 B.n41 71.676
R456 B.n90 B.n42 71.676
R457 B.n94 B.n43 71.676
R458 B.n99 B.n44 71.676
R459 B.n103 B.n45 71.676
R460 B.n107 B.n46 71.676
R461 B.n111 B.n47 71.676
R462 B.n115 B.n48 71.676
R463 B.n119 B.n49 71.676
R464 B.n123 B.n50 71.676
R465 B.n127 B.n51 71.676
R466 B.n131 B.n52 71.676
R467 B.n135 B.n53 71.676
R468 B.n139 B.n54 71.676
R469 B.n143 B.n55 71.676
R470 B.n56 B.n55 71.676
R471 B.n142 B.n54 71.676
R472 B.n138 B.n53 71.676
R473 B.n134 B.n52 71.676
R474 B.n130 B.n51 71.676
R475 B.n126 B.n50 71.676
R476 B.n122 B.n49 71.676
R477 B.n118 B.n48 71.676
R478 B.n114 B.n47 71.676
R479 B.n110 B.n46 71.676
R480 B.n106 B.n45 71.676
R481 B.n102 B.n44 71.676
R482 B.n98 B.n43 71.676
R483 B.n93 B.n42 71.676
R484 B.n89 B.n41 71.676
R485 B.n85 B.n40 71.676
R486 B.n81 B.n39 71.676
R487 B.n77 B.n38 71.676
R488 B.n73 B.n37 71.676
R489 B.n69 B.n36 71.676
R490 B.n65 B.n35 71.676
R491 B.n287 B.n200 71.676
R492 B.n279 B.n180 71.676
R493 B.n275 B.n181 71.676
R494 B.n271 B.n182 71.676
R495 B.n267 B.n183 71.676
R496 B.n263 B.n184 71.676
R497 B.n259 B.n185 71.676
R498 B.n255 B.n186 71.676
R499 B.n251 B.n187 71.676
R500 B.n247 B.n188 71.676
R501 B.n243 B.n189 71.676
R502 B.n239 B.n190 71.676
R503 B.n234 B.n191 71.676
R504 B.n230 B.n192 71.676
R505 B.n226 B.n193 71.676
R506 B.n222 B.n194 71.676
R507 B.n218 B.n195 71.676
R508 B.n214 B.n196 71.676
R509 B.n210 B.n197 71.676
R510 B.n206 B.n198 71.676
R511 B.n290 B.n289 71.676
R512 B.t0 B.n148 70.7281
R513 B.t1 B.n8 70.7281
R514 B.n236 B.n205 59.5399
R515 B.n203 B.n202 59.5399
R516 B.n96 B.n61 59.5399
R517 B.n59 B.n58 59.5399
R518 B.t3 B.n164 43.4297
R519 B.t10 B.n22 43.4297
R520 B.n307 B.t3 40.948
R521 B.n376 B.t10 40.948
R522 B.n63 B.n31 34.8103
R523 B.n364 B.n363 34.8103
R524 B.n292 B.n291 34.8103
R525 B.n285 B.n174 34.8103
R526 B.n205 B.n204 29.4793
R527 B.n202 B.n201 29.4793
R528 B.n61 B.n60 29.4793
R529 B.n58 B.n57 29.4793
R530 B B.n402 18.0485
R531 B.n332 B.t0 13.6497
R532 B.n392 B.t1 13.6497
R533 B.n64 B.n63 10.6151
R534 B.n67 B.n64 10.6151
R535 B.n68 B.n67 10.6151
R536 B.n71 B.n68 10.6151
R537 B.n72 B.n71 10.6151
R538 B.n75 B.n72 10.6151
R539 B.n76 B.n75 10.6151
R540 B.n79 B.n76 10.6151
R541 B.n80 B.n79 10.6151
R542 B.n83 B.n80 10.6151
R543 B.n84 B.n83 10.6151
R544 B.n87 B.n84 10.6151
R545 B.n88 B.n87 10.6151
R546 B.n91 B.n88 10.6151
R547 B.n92 B.n91 10.6151
R548 B.n95 B.n92 10.6151
R549 B.n100 B.n97 10.6151
R550 B.n101 B.n100 10.6151
R551 B.n104 B.n101 10.6151
R552 B.n105 B.n104 10.6151
R553 B.n108 B.n105 10.6151
R554 B.n109 B.n108 10.6151
R555 B.n112 B.n109 10.6151
R556 B.n113 B.n112 10.6151
R557 B.n117 B.n116 10.6151
R558 B.n120 B.n117 10.6151
R559 B.n121 B.n120 10.6151
R560 B.n124 B.n121 10.6151
R561 B.n125 B.n124 10.6151
R562 B.n128 B.n125 10.6151
R563 B.n129 B.n128 10.6151
R564 B.n132 B.n129 10.6151
R565 B.n133 B.n132 10.6151
R566 B.n136 B.n133 10.6151
R567 B.n137 B.n136 10.6151
R568 B.n140 B.n137 10.6151
R569 B.n141 B.n140 10.6151
R570 B.n144 B.n141 10.6151
R571 B.n145 B.n144 10.6151
R572 B.n364 B.n145 10.6151
R573 B.n293 B.n292 10.6151
R574 B.n293 B.n170 10.6151
R575 B.n303 B.n170 10.6151
R576 B.n304 B.n303 10.6151
R577 B.n305 B.n304 10.6151
R578 B.n305 B.n162 10.6151
R579 B.n315 B.n162 10.6151
R580 B.n316 B.n315 10.6151
R581 B.n317 B.n316 10.6151
R582 B.n317 B.n154 10.6151
R583 B.n327 B.n154 10.6151
R584 B.n328 B.n327 10.6151
R585 B.n330 B.n328 10.6151
R586 B.n330 B.n329 10.6151
R587 B.n329 B.n146 10.6151
R588 B.n341 B.n146 10.6151
R589 B.n342 B.n341 10.6151
R590 B.n343 B.n342 10.6151
R591 B.n344 B.n343 10.6151
R592 B.n346 B.n344 10.6151
R593 B.n347 B.n346 10.6151
R594 B.n348 B.n347 10.6151
R595 B.n349 B.n348 10.6151
R596 B.n351 B.n349 10.6151
R597 B.n352 B.n351 10.6151
R598 B.n353 B.n352 10.6151
R599 B.n354 B.n353 10.6151
R600 B.n356 B.n354 10.6151
R601 B.n357 B.n356 10.6151
R602 B.n358 B.n357 10.6151
R603 B.n359 B.n358 10.6151
R604 B.n361 B.n359 10.6151
R605 B.n362 B.n361 10.6151
R606 B.n363 B.n362 10.6151
R607 B.n285 B.n284 10.6151
R608 B.n284 B.n283 10.6151
R609 B.n283 B.n282 10.6151
R610 B.n282 B.n280 10.6151
R611 B.n280 B.n277 10.6151
R612 B.n277 B.n276 10.6151
R613 B.n276 B.n273 10.6151
R614 B.n273 B.n272 10.6151
R615 B.n272 B.n269 10.6151
R616 B.n269 B.n268 10.6151
R617 B.n268 B.n265 10.6151
R618 B.n265 B.n264 10.6151
R619 B.n264 B.n261 10.6151
R620 B.n261 B.n260 10.6151
R621 B.n260 B.n257 10.6151
R622 B.n257 B.n256 10.6151
R623 B.n253 B.n252 10.6151
R624 B.n252 B.n249 10.6151
R625 B.n249 B.n248 10.6151
R626 B.n248 B.n245 10.6151
R627 B.n245 B.n244 10.6151
R628 B.n244 B.n241 10.6151
R629 B.n241 B.n240 10.6151
R630 B.n240 B.n237 10.6151
R631 B.n235 B.n232 10.6151
R632 B.n232 B.n231 10.6151
R633 B.n231 B.n228 10.6151
R634 B.n228 B.n227 10.6151
R635 B.n227 B.n224 10.6151
R636 B.n224 B.n223 10.6151
R637 B.n223 B.n220 10.6151
R638 B.n220 B.n219 10.6151
R639 B.n219 B.n216 10.6151
R640 B.n216 B.n215 10.6151
R641 B.n215 B.n212 10.6151
R642 B.n212 B.n211 10.6151
R643 B.n211 B.n208 10.6151
R644 B.n208 B.n207 10.6151
R645 B.n207 B.n178 10.6151
R646 B.n291 B.n178 10.6151
R647 B.n297 B.n174 10.6151
R648 B.n298 B.n297 10.6151
R649 B.n299 B.n298 10.6151
R650 B.n299 B.n166 10.6151
R651 B.n309 B.n166 10.6151
R652 B.n310 B.n309 10.6151
R653 B.n311 B.n310 10.6151
R654 B.n311 B.n158 10.6151
R655 B.n321 B.n158 10.6151
R656 B.n322 B.n321 10.6151
R657 B.n323 B.n322 10.6151
R658 B.n323 B.n150 10.6151
R659 B.n334 B.n150 10.6151
R660 B.n335 B.n334 10.6151
R661 B.n336 B.n335 10.6151
R662 B.n336 B.n0 10.6151
R663 B.n396 B.n1 10.6151
R664 B.n396 B.n395 10.6151
R665 B.n395 B.n394 10.6151
R666 B.n394 B.n10 10.6151
R667 B.n388 B.n10 10.6151
R668 B.n388 B.n387 10.6151
R669 B.n387 B.n386 10.6151
R670 B.n386 B.n17 10.6151
R671 B.n380 B.n17 10.6151
R672 B.n380 B.n379 10.6151
R673 B.n379 B.n378 10.6151
R674 B.n378 B.n24 10.6151
R675 B.n372 B.n24 10.6151
R676 B.n372 B.n371 10.6151
R677 B.n371 B.n370 10.6151
R678 B.n370 B.n31 10.6151
R679 B.n97 B.n96 6.5566
R680 B.n113 B.n59 6.5566
R681 B.n253 B.n203 6.5566
R682 B.n237 B.n236 6.5566
R683 B.n96 B.n95 4.05904
R684 B.n116 B.n59 4.05904
R685 B.n256 B.n203 4.05904
R686 B.n236 B.n235 4.05904
R687 B.n402 B.n0 2.81026
R688 B.n402 B.n1 2.81026
R689 VN VN.t1 221.355
R690 VN VN.t0 186.668
R691 VTAIL.n1 VTAIL.t2 66.3304
R692 VTAIL.n3 VTAIL.t3 66.3304
R693 VTAIL.n0 VTAIL.t0 66.3304
R694 VTAIL.n2 VTAIL.t1 66.3304
R695 VTAIL.n1 VTAIL.n0 18.0824
R696 VTAIL.n3 VTAIL.n2 16.7721
R697 VTAIL.n2 VTAIL.n1 1.1255
R698 VTAIL VTAIL.n0 0.856103
R699 VTAIL VTAIL.n3 0.269897
R700 VDD2.n0 VDD2.t1 112.385
R701 VDD2.n0 VDD2.t0 83.0092
R702 VDD2 VDD2.n0 0.386276
R703 VP.n0 VP.t1 221.069
R704 VP.n0 VP.t0 186.523
R705 VP VP.n0 0.146778
R706 VDD1 VDD1.t1 113.237
R707 VDD1 VDD1.t0 83.3949
C0 VDD2 VP 0.277923f
C1 VDD2 VTAIL 2.56938f
C2 VDD2 VDD1 0.510401f
C3 VN VP 3.24483f
C4 VTAIL VN 0.872988f
C5 VDD1 VN 0.152015f
C6 VTAIL VP 0.887206f
C7 VDD2 VN 0.875061f
C8 VDD1 VP 0.999282f
C9 VDD1 VTAIL 2.52705f
C10 VDD2 B 2.390563f
C11 VDD1 B 3.96387f
C12 VTAIL B 3.197478f
C13 VN B 6.08476f
C14 VP B 3.953375f
C15 VDD1.t0 B 0.418371f
C16 VDD1.t1 B 0.601341f
C17 VP.t1 B 0.669687f
C18 VP.t0 B 0.500486f
C19 VP.n0 B 2.00256f
C20 VDD2.t1 B 0.624594f
C21 VDD2.t0 B 0.444158f
C22 VDD2.n0 B 1.47722f
C23 VTAIL.t0 B 0.467748f
C24 VTAIL.n0 B 0.830079f
C25 VTAIL.t2 B 0.467751f
C26 VTAIL.n1 B 0.846017f
C27 VTAIL.t1 B 0.467748f
C28 VTAIL.n2 B 0.768485f
C29 VTAIL.t3 B 0.467748f
C30 VTAIL.n3 B 0.717857f
C31 VN.t0 B 0.493629f
C32 VN.t1 B 0.664415f
.ends

