* NGSPICE file created from diff_pair_sample_1746.ext - technology: sky130A

.subckt diff_pair_sample_1746 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X1 VTAIL.t19 VN.t0 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X2 VDD1.t7 VP.t1 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X3 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0.9603 ps=6.15 w=5.82 l=3.63
X4 VDD1.t3 VP.t2 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X5 VTAIL.t2 VN.t2 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X6 VTAIL.t15 VP.t3 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X7 VDD2.t6 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X8 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0 ps=0 w=5.82 l=3.63
X9 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X10 VTAIL.t14 VP.t4 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X11 VDD1.t2 VP.t5 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=2.2698 ps=12.42 w=5.82 l=3.63
X12 VDD1.t6 VP.t6 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0.9603 ps=6.15 w=5.82 l=3.63
X13 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0 ps=0 w=5.82 l=3.63
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0 ps=0 w=5.82 l=3.63
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0 ps=0 w=5.82 l=3.63
X16 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=2.2698 ps=12.42 w=5.82 l=3.63
X17 VTAIL.t6 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X18 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0.9603 ps=6.15 w=5.82 l=3.63
X19 VDD2.t1 VN.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=2.2698 ps=12.42 w=5.82 l=3.63
X20 VTAIL.t8 VN.t9 VDD2.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X21 VTAIL.t11 VP.t7 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=0.9603 ps=6.15 w=5.82 l=3.63
X22 VDD1.t8 VP.t8 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9603 pd=6.15 as=2.2698 ps=12.42 w=5.82 l=3.63
X23 VDD1.t0 VP.t9 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2698 pd=12.42 as=0.9603 ps=6.15 w=5.82 l=3.63
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n72 VP.n71 81.8843
R57 VP.n124 VP.n0 81.8843
R58 VP.n70 VP.n17 81.8843
R59 VP.n31 VP.t9 71.8349
R60 VP.n31 VP.n30 64.4539
R61 VP.n77 VP.n14 56.5617
R62 VP.n116 VP.n2 56.5617
R63 VP.n62 VP.n19 56.5617
R64 VP.n90 VP.n10 56.5617
R65 VP.n103 VP.n6 56.5617
R66 VP.n49 VP.n23 56.5617
R67 VP.n36 VP.n27 56.5617
R68 VP.n72 VP.n70 54.1283
R69 VP.n71 VP.t6 38.6402
R70 VP.n83 VP.t7 38.6402
R71 VP.n96 VP.t2 38.6402
R72 VP.n109 VP.t4 38.6402
R73 VP.n0 VP.t5 38.6402
R74 VP.n17 VP.t8 38.6402
R75 VP.n55 VP.t0 38.6402
R76 VP.n42 VP.t1 38.6402
R77 VP.n30 VP.t3 38.6402
R78 VP.n75 VP.n16 24.5923
R79 VP.n76 VP.n75 24.5923
R80 VP.n77 VP.n76 24.5923
R81 VP.n81 VP.n14 24.5923
R82 VP.n82 VP.n81 24.5923
R83 VP.n84 VP.n82 24.5923
R84 VP.n88 VP.n12 24.5923
R85 VP.n89 VP.n88 24.5923
R86 VP.n90 VP.n89 24.5923
R87 VP.n94 VP.n10 24.5923
R88 VP.n95 VP.n94 24.5923
R89 VP.n97 VP.n95 24.5923
R90 VP.n101 VP.n8 24.5923
R91 VP.n102 VP.n101 24.5923
R92 VP.n103 VP.n102 24.5923
R93 VP.n107 VP.n6 24.5923
R94 VP.n108 VP.n107 24.5923
R95 VP.n110 VP.n108 24.5923
R96 VP.n114 VP.n4 24.5923
R97 VP.n115 VP.n114 24.5923
R98 VP.n116 VP.n115 24.5923
R99 VP.n120 VP.n2 24.5923
R100 VP.n121 VP.n120 24.5923
R101 VP.n122 VP.n121 24.5923
R102 VP.n66 VP.n19 24.5923
R103 VP.n67 VP.n66 24.5923
R104 VP.n68 VP.n67 24.5923
R105 VP.n53 VP.n23 24.5923
R106 VP.n54 VP.n53 24.5923
R107 VP.n56 VP.n54 24.5923
R108 VP.n60 VP.n21 24.5923
R109 VP.n61 VP.n60 24.5923
R110 VP.n62 VP.n61 24.5923
R111 VP.n40 VP.n27 24.5923
R112 VP.n41 VP.n40 24.5923
R113 VP.n43 VP.n41 24.5923
R114 VP.n47 VP.n25 24.5923
R115 VP.n48 VP.n47 24.5923
R116 VP.n49 VP.n48 24.5923
R117 VP.n34 VP.n29 24.5923
R118 VP.n35 VP.n34 24.5923
R119 VP.n36 VP.n35 24.5923
R120 VP.n84 VP.n83 14.2638
R121 VP.n109 VP.n4 14.2638
R122 VP.n55 VP.n21 14.2638
R123 VP.n97 VP.n96 12.2964
R124 VP.n96 VP.n8 12.2964
R125 VP.n43 VP.n42 12.2964
R126 VP.n42 VP.n25 12.2964
R127 VP.n83 VP.n12 10.3291
R128 VP.n110 VP.n109 10.3291
R129 VP.n56 VP.n55 10.3291
R130 VP.n30 VP.n29 10.3291
R131 VP.n71 VP.n16 8.36172
R132 VP.n122 VP.n0 8.36172
R133 VP.n68 VP.n17 8.36172
R134 VP.n32 VP.n31 3.19892
R135 VP.n70 VP.n69 0.354861
R136 VP.n73 VP.n72 0.354861
R137 VP.n124 VP.n123 0.354861
R138 VP VP.n124 0.267071
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VDD1.n28 VDD1.n27 289.615
R194 VDD1.n59 VDD1.n58 289.615
R195 VDD1.n27 VDD1.n26 185
R196 VDD1.n2 VDD1.n1 185
R197 VDD1.n21 VDD1.n20 185
R198 VDD1.n19 VDD1.n18 185
R199 VDD1.n6 VDD1.n5 185
R200 VDD1.n13 VDD1.n12 185
R201 VDD1.n11 VDD1.n10 185
R202 VDD1.n42 VDD1.n41 185
R203 VDD1.n44 VDD1.n43 185
R204 VDD1.n37 VDD1.n36 185
R205 VDD1.n50 VDD1.n49 185
R206 VDD1.n52 VDD1.n51 185
R207 VDD1.n33 VDD1.n32 185
R208 VDD1.n58 VDD1.n57 185
R209 VDD1.n9 VDD1.t0 149.528
R210 VDD1.n40 VDD1.t6 149.528
R211 VDD1.n27 VDD1.n1 104.615
R212 VDD1.n20 VDD1.n1 104.615
R213 VDD1.n20 VDD1.n19 104.615
R214 VDD1.n19 VDD1.n5 104.615
R215 VDD1.n12 VDD1.n5 104.615
R216 VDD1.n12 VDD1.n11 104.615
R217 VDD1.n43 VDD1.n42 104.615
R218 VDD1.n43 VDD1.n36 104.615
R219 VDD1.n50 VDD1.n36 104.615
R220 VDD1.n51 VDD1.n50 104.615
R221 VDD1.n51 VDD1.n32 104.615
R222 VDD1.n58 VDD1.n32 104.615
R223 VDD1.n63 VDD1.n62 72.3701
R224 VDD1.n30 VDD1.n29 69.8661
R225 VDD1.n61 VDD1.n60 69.8651
R226 VDD1.n65 VDD1.n64 69.865
R227 VDD1.n30 VDD1.n28 54.6052
R228 VDD1.n61 VDD1.n59 54.6052
R229 VDD1.n11 VDD1.t0 52.3082
R230 VDD1.n42 VDD1.t6 52.3082
R231 VDD1.n65 VDD1.n63 47.238
R232 VDD1.n26 VDD1.n0 12.0247
R233 VDD1.n57 VDD1.n31 12.0247
R234 VDD1.n25 VDD1.n2 11.249
R235 VDD1.n56 VDD1.n33 11.249
R236 VDD1.n22 VDD1.n21 10.4732
R237 VDD1.n53 VDD1.n52 10.4732
R238 VDD1.n10 VDD1.n9 10.2745
R239 VDD1.n41 VDD1.n40 10.2745
R240 VDD1.n18 VDD1.n4 9.69747
R241 VDD1.n49 VDD1.n35 9.69747
R242 VDD1.n24 VDD1.n0 9.45567
R243 VDD1.n55 VDD1.n31 9.45567
R244 VDD1.n15 VDD1.n14 9.3005
R245 VDD1.n17 VDD1.n16 9.3005
R246 VDD1.n4 VDD1.n3 9.3005
R247 VDD1.n23 VDD1.n22 9.3005
R248 VDD1.n25 VDD1.n24 9.3005
R249 VDD1.n8 VDD1.n7 9.3005
R250 VDD1.n39 VDD1.n38 9.3005
R251 VDD1.n46 VDD1.n45 9.3005
R252 VDD1.n48 VDD1.n47 9.3005
R253 VDD1.n35 VDD1.n34 9.3005
R254 VDD1.n54 VDD1.n53 9.3005
R255 VDD1.n56 VDD1.n55 9.3005
R256 VDD1.n17 VDD1.n6 8.92171
R257 VDD1.n48 VDD1.n37 8.92171
R258 VDD1.n14 VDD1.n13 8.14595
R259 VDD1.n45 VDD1.n44 8.14595
R260 VDD1.n10 VDD1.n8 7.3702
R261 VDD1.n41 VDD1.n39 7.3702
R262 VDD1.n13 VDD1.n8 5.81868
R263 VDD1.n44 VDD1.n39 5.81868
R264 VDD1.n14 VDD1.n6 5.04292
R265 VDD1.n45 VDD1.n37 5.04292
R266 VDD1.n18 VDD1.n17 4.26717
R267 VDD1.n49 VDD1.n48 4.26717
R268 VDD1.n21 VDD1.n4 3.49141
R269 VDD1.n52 VDD1.n35 3.49141
R270 VDD1.n64 VDD1.t9 3.40256
R271 VDD1.n64 VDD1.t8 3.40256
R272 VDD1.n29 VDD1.t5 3.40256
R273 VDD1.n29 VDD1.t7 3.40256
R274 VDD1.n62 VDD1.t1 3.40256
R275 VDD1.n62 VDD1.t2 3.40256
R276 VDD1.n60 VDD1.t4 3.40256
R277 VDD1.n60 VDD1.t3 3.40256
R278 VDD1.n9 VDD1.n7 2.84323
R279 VDD1.n40 VDD1.n38 2.84323
R280 VDD1.n22 VDD1.n2 2.71565
R281 VDD1.n53 VDD1.n33 2.71565
R282 VDD1 VDD1.n65 2.50266
R283 VDD1.n26 VDD1.n25 1.93989
R284 VDD1.n57 VDD1.n56 1.93989
R285 VDD1.n28 VDD1.n0 1.16414
R286 VDD1.n59 VDD1.n31 1.16414
R287 VDD1 VDD1.n30 0.912138
R288 VDD1.n63 VDD1.n61 0.798602
R289 VDD1.n24 VDD1.n23 0.155672
R290 VDD1.n23 VDD1.n3 0.155672
R291 VDD1.n16 VDD1.n3 0.155672
R292 VDD1.n16 VDD1.n15 0.155672
R293 VDD1.n15 VDD1.n7 0.155672
R294 VDD1.n46 VDD1.n38 0.155672
R295 VDD1.n47 VDD1.n46 0.155672
R296 VDD1.n47 VDD1.n34 0.155672
R297 VDD1.n54 VDD1.n34 0.155672
R298 VDD1.n55 VDD1.n54 0.155672
R299 VTAIL.n132 VTAIL.n131 289.615
R300 VTAIL.n30 VTAIL.n29 289.615
R301 VTAIL.n102 VTAIL.n101 289.615
R302 VTAIL.n68 VTAIL.n67 289.615
R303 VTAIL.n115 VTAIL.n114 185
R304 VTAIL.n117 VTAIL.n116 185
R305 VTAIL.n110 VTAIL.n109 185
R306 VTAIL.n123 VTAIL.n122 185
R307 VTAIL.n125 VTAIL.n124 185
R308 VTAIL.n106 VTAIL.n105 185
R309 VTAIL.n131 VTAIL.n130 185
R310 VTAIL.n13 VTAIL.n12 185
R311 VTAIL.n15 VTAIL.n14 185
R312 VTAIL.n8 VTAIL.n7 185
R313 VTAIL.n21 VTAIL.n20 185
R314 VTAIL.n23 VTAIL.n22 185
R315 VTAIL.n4 VTAIL.n3 185
R316 VTAIL.n29 VTAIL.n28 185
R317 VTAIL.n101 VTAIL.n100 185
R318 VTAIL.n76 VTAIL.n75 185
R319 VTAIL.n95 VTAIL.n94 185
R320 VTAIL.n93 VTAIL.n92 185
R321 VTAIL.n80 VTAIL.n79 185
R322 VTAIL.n87 VTAIL.n86 185
R323 VTAIL.n85 VTAIL.n84 185
R324 VTAIL.n67 VTAIL.n66 185
R325 VTAIL.n42 VTAIL.n41 185
R326 VTAIL.n61 VTAIL.n60 185
R327 VTAIL.n59 VTAIL.n58 185
R328 VTAIL.n46 VTAIL.n45 185
R329 VTAIL.n53 VTAIL.n52 185
R330 VTAIL.n51 VTAIL.n50 185
R331 VTAIL.n113 VTAIL.t7 149.528
R332 VTAIL.n11 VTAIL.t13 149.528
R333 VTAIL.n83 VTAIL.t10 149.528
R334 VTAIL.n49 VTAIL.t4 149.528
R335 VTAIL.n116 VTAIL.n115 104.615
R336 VTAIL.n116 VTAIL.n109 104.615
R337 VTAIL.n123 VTAIL.n109 104.615
R338 VTAIL.n124 VTAIL.n123 104.615
R339 VTAIL.n124 VTAIL.n105 104.615
R340 VTAIL.n131 VTAIL.n105 104.615
R341 VTAIL.n14 VTAIL.n13 104.615
R342 VTAIL.n14 VTAIL.n7 104.615
R343 VTAIL.n21 VTAIL.n7 104.615
R344 VTAIL.n22 VTAIL.n21 104.615
R345 VTAIL.n22 VTAIL.n3 104.615
R346 VTAIL.n29 VTAIL.n3 104.615
R347 VTAIL.n101 VTAIL.n75 104.615
R348 VTAIL.n94 VTAIL.n75 104.615
R349 VTAIL.n94 VTAIL.n93 104.615
R350 VTAIL.n93 VTAIL.n79 104.615
R351 VTAIL.n86 VTAIL.n79 104.615
R352 VTAIL.n86 VTAIL.n85 104.615
R353 VTAIL.n67 VTAIL.n41 104.615
R354 VTAIL.n60 VTAIL.n41 104.615
R355 VTAIL.n60 VTAIL.n59 104.615
R356 VTAIL.n59 VTAIL.n45 104.615
R357 VTAIL.n52 VTAIL.n45 104.615
R358 VTAIL.n52 VTAIL.n51 104.615
R359 VTAIL.n73 VTAIL.n72 53.1873
R360 VTAIL.n71 VTAIL.n70 53.1873
R361 VTAIL.n39 VTAIL.n38 53.1873
R362 VTAIL.n37 VTAIL.n36 53.1873
R363 VTAIL.n135 VTAIL.n134 53.1863
R364 VTAIL.n1 VTAIL.n0 53.1863
R365 VTAIL.n33 VTAIL.n32 53.1863
R366 VTAIL.n35 VTAIL.n34 53.1863
R367 VTAIL.n115 VTAIL.t7 52.3082
R368 VTAIL.n13 VTAIL.t13 52.3082
R369 VTAIL.n85 VTAIL.t10 52.3082
R370 VTAIL.n51 VTAIL.t4 52.3082
R371 VTAIL.n133 VTAIL.n132 34.5126
R372 VTAIL.n31 VTAIL.n30 34.5126
R373 VTAIL.n103 VTAIL.n102 34.5126
R374 VTAIL.n69 VTAIL.n68 34.5126
R375 VTAIL.n37 VTAIL.n35 24.2117
R376 VTAIL.n133 VTAIL.n103 20.7979
R377 VTAIL.n130 VTAIL.n104 12.0247
R378 VTAIL.n28 VTAIL.n2 12.0247
R379 VTAIL.n100 VTAIL.n74 12.0247
R380 VTAIL.n66 VTAIL.n40 12.0247
R381 VTAIL.n129 VTAIL.n106 11.249
R382 VTAIL.n27 VTAIL.n4 11.249
R383 VTAIL.n99 VTAIL.n76 11.249
R384 VTAIL.n65 VTAIL.n42 11.249
R385 VTAIL.n126 VTAIL.n125 10.4732
R386 VTAIL.n24 VTAIL.n23 10.4732
R387 VTAIL.n96 VTAIL.n95 10.4732
R388 VTAIL.n62 VTAIL.n61 10.4732
R389 VTAIL.n114 VTAIL.n113 10.2745
R390 VTAIL.n12 VTAIL.n11 10.2745
R391 VTAIL.n84 VTAIL.n83 10.2745
R392 VTAIL.n50 VTAIL.n49 10.2745
R393 VTAIL.n122 VTAIL.n108 9.69747
R394 VTAIL.n20 VTAIL.n6 9.69747
R395 VTAIL.n92 VTAIL.n78 9.69747
R396 VTAIL.n58 VTAIL.n44 9.69747
R397 VTAIL.n128 VTAIL.n104 9.45567
R398 VTAIL.n26 VTAIL.n2 9.45567
R399 VTAIL.n98 VTAIL.n74 9.45567
R400 VTAIL.n64 VTAIL.n40 9.45567
R401 VTAIL.n112 VTAIL.n111 9.3005
R402 VTAIL.n119 VTAIL.n118 9.3005
R403 VTAIL.n121 VTAIL.n120 9.3005
R404 VTAIL.n108 VTAIL.n107 9.3005
R405 VTAIL.n127 VTAIL.n126 9.3005
R406 VTAIL.n129 VTAIL.n128 9.3005
R407 VTAIL.n10 VTAIL.n9 9.3005
R408 VTAIL.n17 VTAIL.n16 9.3005
R409 VTAIL.n19 VTAIL.n18 9.3005
R410 VTAIL.n6 VTAIL.n5 9.3005
R411 VTAIL.n25 VTAIL.n24 9.3005
R412 VTAIL.n27 VTAIL.n26 9.3005
R413 VTAIL.n99 VTAIL.n98 9.3005
R414 VTAIL.n97 VTAIL.n96 9.3005
R415 VTAIL.n78 VTAIL.n77 9.3005
R416 VTAIL.n91 VTAIL.n90 9.3005
R417 VTAIL.n89 VTAIL.n88 9.3005
R418 VTAIL.n82 VTAIL.n81 9.3005
R419 VTAIL.n55 VTAIL.n54 9.3005
R420 VTAIL.n57 VTAIL.n56 9.3005
R421 VTAIL.n44 VTAIL.n43 9.3005
R422 VTAIL.n63 VTAIL.n62 9.3005
R423 VTAIL.n65 VTAIL.n64 9.3005
R424 VTAIL.n48 VTAIL.n47 9.3005
R425 VTAIL.n121 VTAIL.n110 8.92171
R426 VTAIL.n19 VTAIL.n8 8.92171
R427 VTAIL.n91 VTAIL.n80 8.92171
R428 VTAIL.n57 VTAIL.n46 8.92171
R429 VTAIL.n118 VTAIL.n117 8.14595
R430 VTAIL.n16 VTAIL.n15 8.14595
R431 VTAIL.n88 VTAIL.n87 8.14595
R432 VTAIL.n54 VTAIL.n53 8.14595
R433 VTAIL.n114 VTAIL.n112 7.3702
R434 VTAIL.n12 VTAIL.n10 7.3702
R435 VTAIL.n84 VTAIL.n82 7.3702
R436 VTAIL.n50 VTAIL.n48 7.3702
R437 VTAIL.n117 VTAIL.n112 5.81868
R438 VTAIL.n15 VTAIL.n10 5.81868
R439 VTAIL.n87 VTAIL.n82 5.81868
R440 VTAIL.n53 VTAIL.n48 5.81868
R441 VTAIL.n118 VTAIL.n110 5.04292
R442 VTAIL.n16 VTAIL.n8 5.04292
R443 VTAIL.n88 VTAIL.n80 5.04292
R444 VTAIL.n54 VTAIL.n46 5.04292
R445 VTAIL.n122 VTAIL.n121 4.26717
R446 VTAIL.n20 VTAIL.n19 4.26717
R447 VTAIL.n92 VTAIL.n91 4.26717
R448 VTAIL.n58 VTAIL.n57 4.26717
R449 VTAIL.n125 VTAIL.n108 3.49141
R450 VTAIL.n23 VTAIL.n6 3.49141
R451 VTAIL.n95 VTAIL.n78 3.49141
R452 VTAIL.n61 VTAIL.n44 3.49141
R453 VTAIL.n39 VTAIL.n37 3.41429
R454 VTAIL.n69 VTAIL.n39 3.41429
R455 VTAIL.n73 VTAIL.n71 3.41429
R456 VTAIL.n103 VTAIL.n73 3.41429
R457 VTAIL.n35 VTAIL.n33 3.41429
R458 VTAIL.n33 VTAIL.n31 3.41429
R459 VTAIL.n135 VTAIL.n133 3.41429
R460 VTAIL.n134 VTAIL.t1 3.40256
R461 VTAIL.n134 VTAIL.t19 3.40256
R462 VTAIL.n0 VTAIL.t5 3.40256
R463 VTAIL.n0 VTAIL.t6 3.40256
R464 VTAIL.n32 VTAIL.t16 3.40256
R465 VTAIL.n32 VTAIL.t14 3.40256
R466 VTAIL.n34 VTAIL.t12 3.40256
R467 VTAIL.n34 VTAIL.t11 3.40256
R468 VTAIL.n72 VTAIL.t17 3.40256
R469 VTAIL.n72 VTAIL.t18 3.40256
R470 VTAIL.n70 VTAIL.t9 3.40256
R471 VTAIL.n70 VTAIL.t15 3.40256
R472 VTAIL.n38 VTAIL.t0 3.40256
R473 VTAIL.n38 VTAIL.t8 3.40256
R474 VTAIL.n36 VTAIL.t3 3.40256
R475 VTAIL.n36 VTAIL.t2 3.40256
R476 VTAIL.n83 VTAIL.n81 2.84323
R477 VTAIL.n49 VTAIL.n47 2.84323
R478 VTAIL.n113 VTAIL.n111 2.84323
R479 VTAIL.n11 VTAIL.n9 2.84323
R480 VTAIL.n126 VTAIL.n106 2.71565
R481 VTAIL.n24 VTAIL.n4 2.71565
R482 VTAIL.n96 VTAIL.n76 2.71565
R483 VTAIL.n62 VTAIL.n42 2.71565
R484 VTAIL VTAIL.n1 2.61903
R485 VTAIL.n71 VTAIL.n69 2.17722
R486 VTAIL.n31 VTAIL.n1 2.17722
R487 VTAIL.n130 VTAIL.n129 1.93989
R488 VTAIL.n28 VTAIL.n27 1.93989
R489 VTAIL.n100 VTAIL.n99 1.93989
R490 VTAIL.n66 VTAIL.n65 1.93989
R491 VTAIL.n132 VTAIL.n104 1.16414
R492 VTAIL.n30 VTAIL.n2 1.16414
R493 VTAIL.n102 VTAIL.n74 1.16414
R494 VTAIL.n68 VTAIL.n40 1.16414
R495 VTAIL VTAIL.n135 0.795759
R496 VTAIL.n119 VTAIL.n111 0.155672
R497 VTAIL.n120 VTAIL.n119 0.155672
R498 VTAIL.n120 VTAIL.n107 0.155672
R499 VTAIL.n127 VTAIL.n107 0.155672
R500 VTAIL.n128 VTAIL.n127 0.155672
R501 VTAIL.n17 VTAIL.n9 0.155672
R502 VTAIL.n18 VTAIL.n17 0.155672
R503 VTAIL.n18 VTAIL.n5 0.155672
R504 VTAIL.n25 VTAIL.n5 0.155672
R505 VTAIL.n26 VTAIL.n25 0.155672
R506 VTAIL.n98 VTAIL.n97 0.155672
R507 VTAIL.n97 VTAIL.n77 0.155672
R508 VTAIL.n90 VTAIL.n77 0.155672
R509 VTAIL.n90 VTAIL.n89 0.155672
R510 VTAIL.n89 VTAIL.n81 0.155672
R511 VTAIL.n64 VTAIL.n63 0.155672
R512 VTAIL.n63 VTAIL.n43 0.155672
R513 VTAIL.n56 VTAIL.n43 0.155672
R514 VTAIL.n56 VTAIL.n55 0.155672
R515 VTAIL.n55 VTAIL.n47 0.155672
R516 B.n807 B.n806 585
R517 B.n809 B.n174 585
R518 B.n812 B.n811 585
R519 B.n813 B.n173 585
R520 B.n815 B.n814 585
R521 B.n817 B.n172 585
R522 B.n820 B.n819 585
R523 B.n821 B.n171 585
R524 B.n823 B.n822 585
R525 B.n825 B.n170 585
R526 B.n828 B.n827 585
R527 B.n829 B.n169 585
R528 B.n831 B.n830 585
R529 B.n833 B.n168 585
R530 B.n836 B.n835 585
R531 B.n837 B.n167 585
R532 B.n839 B.n838 585
R533 B.n841 B.n166 585
R534 B.n844 B.n843 585
R535 B.n845 B.n165 585
R536 B.n847 B.n846 585
R537 B.n849 B.n164 585
R538 B.n852 B.n851 585
R539 B.n854 B.n161 585
R540 B.n856 B.n855 585
R541 B.n858 B.n160 585
R542 B.n861 B.n860 585
R543 B.n862 B.n159 585
R544 B.n864 B.n863 585
R545 B.n866 B.n158 585
R546 B.n869 B.n868 585
R547 B.n870 B.n154 585
R548 B.n872 B.n871 585
R549 B.n874 B.n153 585
R550 B.n877 B.n876 585
R551 B.n878 B.n152 585
R552 B.n880 B.n879 585
R553 B.n882 B.n151 585
R554 B.n885 B.n884 585
R555 B.n886 B.n150 585
R556 B.n888 B.n887 585
R557 B.n890 B.n149 585
R558 B.n893 B.n892 585
R559 B.n894 B.n148 585
R560 B.n896 B.n895 585
R561 B.n898 B.n147 585
R562 B.n901 B.n900 585
R563 B.n902 B.n146 585
R564 B.n904 B.n903 585
R565 B.n906 B.n145 585
R566 B.n909 B.n908 585
R567 B.n910 B.n144 585
R568 B.n912 B.n911 585
R569 B.n914 B.n143 585
R570 B.n917 B.n916 585
R571 B.n918 B.n142 585
R572 B.n805 B.n140 585
R573 B.n921 B.n140 585
R574 B.n804 B.n139 585
R575 B.n922 B.n139 585
R576 B.n803 B.n138 585
R577 B.n923 B.n138 585
R578 B.n802 B.n801 585
R579 B.n801 B.n134 585
R580 B.n800 B.n133 585
R581 B.n929 B.n133 585
R582 B.n799 B.n132 585
R583 B.n930 B.n132 585
R584 B.n798 B.n131 585
R585 B.n931 B.n131 585
R586 B.n797 B.n796 585
R587 B.n796 B.n127 585
R588 B.n795 B.n126 585
R589 B.n937 B.n126 585
R590 B.n794 B.n125 585
R591 B.n938 B.n125 585
R592 B.n793 B.n124 585
R593 B.n939 B.n124 585
R594 B.n792 B.n791 585
R595 B.n791 B.n120 585
R596 B.n790 B.n119 585
R597 B.n945 B.n119 585
R598 B.n789 B.n118 585
R599 B.n946 B.n118 585
R600 B.n788 B.n117 585
R601 B.n947 B.n117 585
R602 B.n787 B.n786 585
R603 B.n786 B.n113 585
R604 B.n785 B.n112 585
R605 B.n953 B.n112 585
R606 B.n784 B.n111 585
R607 B.n954 B.n111 585
R608 B.n783 B.n110 585
R609 B.n955 B.n110 585
R610 B.n782 B.n781 585
R611 B.n781 B.n106 585
R612 B.n780 B.n105 585
R613 B.n961 B.n105 585
R614 B.n779 B.n104 585
R615 B.n962 B.n104 585
R616 B.n778 B.n103 585
R617 B.n963 B.n103 585
R618 B.n777 B.n776 585
R619 B.n776 B.n102 585
R620 B.n775 B.n98 585
R621 B.n969 B.n98 585
R622 B.n774 B.n97 585
R623 B.n970 B.n97 585
R624 B.n773 B.n96 585
R625 B.n971 B.n96 585
R626 B.n772 B.n771 585
R627 B.n771 B.n92 585
R628 B.n770 B.n91 585
R629 B.n977 B.n91 585
R630 B.n769 B.n90 585
R631 B.n978 B.n90 585
R632 B.n768 B.n89 585
R633 B.n979 B.n89 585
R634 B.n767 B.n766 585
R635 B.n766 B.n85 585
R636 B.n765 B.n84 585
R637 B.n985 B.n84 585
R638 B.n764 B.n83 585
R639 B.n986 B.n83 585
R640 B.n763 B.n82 585
R641 B.n987 B.n82 585
R642 B.n762 B.n761 585
R643 B.n761 B.n81 585
R644 B.n760 B.n77 585
R645 B.n993 B.n77 585
R646 B.n759 B.n76 585
R647 B.n994 B.n76 585
R648 B.n758 B.n75 585
R649 B.n995 B.n75 585
R650 B.n757 B.n756 585
R651 B.n756 B.n71 585
R652 B.n755 B.n70 585
R653 B.n1001 B.n70 585
R654 B.n754 B.n69 585
R655 B.n1002 B.n69 585
R656 B.n753 B.n68 585
R657 B.n1003 B.n68 585
R658 B.n752 B.n751 585
R659 B.n751 B.n64 585
R660 B.n750 B.n63 585
R661 B.n1009 B.n63 585
R662 B.n749 B.n62 585
R663 B.n1010 B.n62 585
R664 B.n748 B.n61 585
R665 B.n1011 B.n61 585
R666 B.n747 B.n746 585
R667 B.n746 B.n60 585
R668 B.n745 B.n56 585
R669 B.n1017 B.n56 585
R670 B.n744 B.n55 585
R671 B.n1018 B.n55 585
R672 B.n743 B.n54 585
R673 B.n1019 B.n54 585
R674 B.n742 B.n741 585
R675 B.n741 B.n50 585
R676 B.n740 B.n49 585
R677 B.n1025 B.n49 585
R678 B.n739 B.n48 585
R679 B.n1026 B.n48 585
R680 B.n738 B.n47 585
R681 B.n1027 B.n47 585
R682 B.n737 B.n736 585
R683 B.n736 B.n43 585
R684 B.n735 B.n42 585
R685 B.n1033 B.n42 585
R686 B.n734 B.n41 585
R687 B.n1034 B.n41 585
R688 B.n733 B.n40 585
R689 B.n1035 B.n40 585
R690 B.n732 B.n731 585
R691 B.n731 B.n36 585
R692 B.n730 B.n35 585
R693 B.n1041 B.n35 585
R694 B.n729 B.n34 585
R695 B.n1042 B.n34 585
R696 B.n728 B.n33 585
R697 B.n1043 B.n33 585
R698 B.n727 B.n726 585
R699 B.n726 B.n29 585
R700 B.n725 B.n28 585
R701 B.n1049 B.n28 585
R702 B.n724 B.n27 585
R703 B.n1050 B.n27 585
R704 B.n723 B.n26 585
R705 B.n1051 B.n26 585
R706 B.n722 B.n721 585
R707 B.n721 B.n22 585
R708 B.n720 B.n21 585
R709 B.n1057 B.n21 585
R710 B.n719 B.n20 585
R711 B.n1058 B.n20 585
R712 B.n718 B.n19 585
R713 B.n1059 B.n19 585
R714 B.n717 B.n716 585
R715 B.n716 B.n15 585
R716 B.n715 B.n14 585
R717 B.n1065 B.n14 585
R718 B.n714 B.n13 585
R719 B.n1066 B.n13 585
R720 B.n713 B.n12 585
R721 B.n1067 B.n12 585
R722 B.n712 B.n711 585
R723 B.n711 B.n8 585
R724 B.n710 B.n7 585
R725 B.n1073 B.n7 585
R726 B.n709 B.n6 585
R727 B.n1074 B.n6 585
R728 B.n708 B.n5 585
R729 B.n1075 B.n5 585
R730 B.n707 B.n706 585
R731 B.n706 B.n4 585
R732 B.n705 B.n175 585
R733 B.n705 B.n704 585
R734 B.n695 B.n176 585
R735 B.n177 B.n176 585
R736 B.n697 B.n696 585
R737 B.n698 B.n697 585
R738 B.n694 B.n182 585
R739 B.n182 B.n181 585
R740 B.n693 B.n692 585
R741 B.n692 B.n691 585
R742 B.n184 B.n183 585
R743 B.n185 B.n184 585
R744 B.n684 B.n683 585
R745 B.n685 B.n684 585
R746 B.n682 B.n190 585
R747 B.n190 B.n189 585
R748 B.n681 B.n680 585
R749 B.n680 B.n679 585
R750 B.n192 B.n191 585
R751 B.n193 B.n192 585
R752 B.n672 B.n671 585
R753 B.n673 B.n672 585
R754 B.n670 B.n198 585
R755 B.n198 B.n197 585
R756 B.n669 B.n668 585
R757 B.n668 B.n667 585
R758 B.n200 B.n199 585
R759 B.n201 B.n200 585
R760 B.n660 B.n659 585
R761 B.n661 B.n660 585
R762 B.n658 B.n206 585
R763 B.n206 B.n205 585
R764 B.n657 B.n656 585
R765 B.n656 B.n655 585
R766 B.n208 B.n207 585
R767 B.n209 B.n208 585
R768 B.n648 B.n647 585
R769 B.n649 B.n648 585
R770 B.n646 B.n214 585
R771 B.n214 B.n213 585
R772 B.n645 B.n644 585
R773 B.n644 B.n643 585
R774 B.n216 B.n215 585
R775 B.n217 B.n216 585
R776 B.n636 B.n635 585
R777 B.n637 B.n636 585
R778 B.n634 B.n222 585
R779 B.n222 B.n221 585
R780 B.n633 B.n632 585
R781 B.n632 B.n631 585
R782 B.n224 B.n223 585
R783 B.n225 B.n224 585
R784 B.n624 B.n623 585
R785 B.n625 B.n624 585
R786 B.n622 B.n230 585
R787 B.n230 B.n229 585
R788 B.n621 B.n620 585
R789 B.n620 B.n619 585
R790 B.n232 B.n231 585
R791 B.n612 B.n232 585
R792 B.n611 B.n610 585
R793 B.n613 B.n611 585
R794 B.n609 B.n237 585
R795 B.n237 B.n236 585
R796 B.n608 B.n607 585
R797 B.n607 B.n606 585
R798 B.n239 B.n238 585
R799 B.n240 B.n239 585
R800 B.n599 B.n598 585
R801 B.n600 B.n599 585
R802 B.n597 B.n245 585
R803 B.n245 B.n244 585
R804 B.n596 B.n595 585
R805 B.n595 B.n594 585
R806 B.n247 B.n246 585
R807 B.n248 B.n247 585
R808 B.n587 B.n586 585
R809 B.n588 B.n587 585
R810 B.n585 B.n253 585
R811 B.n253 B.n252 585
R812 B.n584 B.n583 585
R813 B.n583 B.n582 585
R814 B.n255 B.n254 585
R815 B.n575 B.n255 585
R816 B.n574 B.n573 585
R817 B.n576 B.n574 585
R818 B.n572 B.n260 585
R819 B.n260 B.n259 585
R820 B.n571 B.n570 585
R821 B.n570 B.n569 585
R822 B.n262 B.n261 585
R823 B.n263 B.n262 585
R824 B.n562 B.n561 585
R825 B.n563 B.n562 585
R826 B.n560 B.n268 585
R827 B.n268 B.n267 585
R828 B.n559 B.n558 585
R829 B.n558 B.n557 585
R830 B.n270 B.n269 585
R831 B.n271 B.n270 585
R832 B.n550 B.n549 585
R833 B.n551 B.n550 585
R834 B.n548 B.n276 585
R835 B.n276 B.n275 585
R836 B.n547 B.n546 585
R837 B.n546 B.n545 585
R838 B.n278 B.n277 585
R839 B.n538 B.n278 585
R840 B.n537 B.n536 585
R841 B.n539 B.n537 585
R842 B.n535 B.n283 585
R843 B.n283 B.n282 585
R844 B.n534 B.n533 585
R845 B.n533 B.n532 585
R846 B.n285 B.n284 585
R847 B.n286 B.n285 585
R848 B.n525 B.n524 585
R849 B.n526 B.n525 585
R850 B.n523 B.n291 585
R851 B.n291 B.n290 585
R852 B.n522 B.n521 585
R853 B.n521 B.n520 585
R854 B.n293 B.n292 585
R855 B.n294 B.n293 585
R856 B.n513 B.n512 585
R857 B.n514 B.n513 585
R858 B.n511 B.n299 585
R859 B.n299 B.n298 585
R860 B.n510 B.n509 585
R861 B.n509 B.n508 585
R862 B.n301 B.n300 585
R863 B.n302 B.n301 585
R864 B.n501 B.n500 585
R865 B.n502 B.n501 585
R866 B.n499 B.n306 585
R867 B.n310 B.n306 585
R868 B.n498 B.n497 585
R869 B.n497 B.n496 585
R870 B.n308 B.n307 585
R871 B.n309 B.n308 585
R872 B.n489 B.n488 585
R873 B.n490 B.n489 585
R874 B.n487 B.n315 585
R875 B.n315 B.n314 585
R876 B.n486 B.n485 585
R877 B.n485 B.n484 585
R878 B.n317 B.n316 585
R879 B.n318 B.n317 585
R880 B.n477 B.n476 585
R881 B.n478 B.n477 585
R882 B.n475 B.n323 585
R883 B.n323 B.n322 585
R884 B.n474 B.n473 585
R885 B.n473 B.n472 585
R886 B.n469 B.n327 585
R887 B.n468 B.n467 585
R888 B.n465 B.n328 585
R889 B.n465 B.n326 585
R890 B.n464 B.n463 585
R891 B.n462 B.n461 585
R892 B.n460 B.n330 585
R893 B.n458 B.n457 585
R894 B.n456 B.n331 585
R895 B.n455 B.n454 585
R896 B.n452 B.n332 585
R897 B.n450 B.n449 585
R898 B.n448 B.n333 585
R899 B.n447 B.n446 585
R900 B.n444 B.n334 585
R901 B.n442 B.n441 585
R902 B.n440 B.n335 585
R903 B.n439 B.n438 585
R904 B.n436 B.n336 585
R905 B.n434 B.n433 585
R906 B.n432 B.n337 585
R907 B.n431 B.n430 585
R908 B.n428 B.n338 585
R909 B.n426 B.n425 585
R910 B.n423 B.n339 585
R911 B.n422 B.n421 585
R912 B.n419 B.n342 585
R913 B.n417 B.n416 585
R914 B.n415 B.n343 585
R915 B.n414 B.n413 585
R916 B.n411 B.n344 585
R917 B.n409 B.n408 585
R918 B.n407 B.n345 585
R919 B.n406 B.n405 585
R920 B.n403 B.n402 585
R921 B.n401 B.n400 585
R922 B.n399 B.n350 585
R923 B.n397 B.n396 585
R924 B.n395 B.n351 585
R925 B.n394 B.n393 585
R926 B.n391 B.n352 585
R927 B.n389 B.n388 585
R928 B.n387 B.n353 585
R929 B.n386 B.n385 585
R930 B.n383 B.n354 585
R931 B.n381 B.n380 585
R932 B.n379 B.n355 585
R933 B.n378 B.n377 585
R934 B.n375 B.n356 585
R935 B.n373 B.n372 585
R936 B.n371 B.n357 585
R937 B.n370 B.n369 585
R938 B.n367 B.n358 585
R939 B.n365 B.n364 585
R940 B.n363 B.n359 585
R941 B.n362 B.n361 585
R942 B.n325 B.n324 585
R943 B.n326 B.n325 585
R944 B.n471 B.n470 585
R945 B.n472 B.n471 585
R946 B.n321 B.n320 585
R947 B.n322 B.n321 585
R948 B.n480 B.n479 585
R949 B.n479 B.n478 585
R950 B.n481 B.n319 585
R951 B.n319 B.n318 585
R952 B.n483 B.n482 585
R953 B.n484 B.n483 585
R954 B.n313 B.n312 585
R955 B.n314 B.n313 585
R956 B.n492 B.n491 585
R957 B.n491 B.n490 585
R958 B.n493 B.n311 585
R959 B.n311 B.n309 585
R960 B.n495 B.n494 585
R961 B.n496 B.n495 585
R962 B.n305 B.n304 585
R963 B.n310 B.n305 585
R964 B.n504 B.n503 585
R965 B.n503 B.n502 585
R966 B.n505 B.n303 585
R967 B.n303 B.n302 585
R968 B.n507 B.n506 585
R969 B.n508 B.n507 585
R970 B.n297 B.n296 585
R971 B.n298 B.n297 585
R972 B.n516 B.n515 585
R973 B.n515 B.n514 585
R974 B.n517 B.n295 585
R975 B.n295 B.n294 585
R976 B.n519 B.n518 585
R977 B.n520 B.n519 585
R978 B.n289 B.n288 585
R979 B.n290 B.n289 585
R980 B.n528 B.n527 585
R981 B.n527 B.n526 585
R982 B.n529 B.n287 585
R983 B.n287 B.n286 585
R984 B.n531 B.n530 585
R985 B.n532 B.n531 585
R986 B.n281 B.n280 585
R987 B.n282 B.n281 585
R988 B.n541 B.n540 585
R989 B.n540 B.n539 585
R990 B.n542 B.n279 585
R991 B.n538 B.n279 585
R992 B.n544 B.n543 585
R993 B.n545 B.n544 585
R994 B.n274 B.n273 585
R995 B.n275 B.n274 585
R996 B.n553 B.n552 585
R997 B.n552 B.n551 585
R998 B.n554 B.n272 585
R999 B.n272 B.n271 585
R1000 B.n556 B.n555 585
R1001 B.n557 B.n556 585
R1002 B.n266 B.n265 585
R1003 B.n267 B.n266 585
R1004 B.n565 B.n564 585
R1005 B.n564 B.n563 585
R1006 B.n566 B.n264 585
R1007 B.n264 B.n263 585
R1008 B.n568 B.n567 585
R1009 B.n569 B.n568 585
R1010 B.n258 B.n257 585
R1011 B.n259 B.n258 585
R1012 B.n578 B.n577 585
R1013 B.n577 B.n576 585
R1014 B.n579 B.n256 585
R1015 B.n575 B.n256 585
R1016 B.n581 B.n580 585
R1017 B.n582 B.n581 585
R1018 B.n251 B.n250 585
R1019 B.n252 B.n251 585
R1020 B.n590 B.n589 585
R1021 B.n589 B.n588 585
R1022 B.n591 B.n249 585
R1023 B.n249 B.n248 585
R1024 B.n593 B.n592 585
R1025 B.n594 B.n593 585
R1026 B.n243 B.n242 585
R1027 B.n244 B.n243 585
R1028 B.n602 B.n601 585
R1029 B.n601 B.n600 585
R1030 B.n603 B.n241 585
R1031 B.n241 B.n240 585
R1032 B.n605 B.n604 585
R1033 B.n606 B.n605 585
R1034 B.n235 B.n234 585
R1035 B.n236 B.n235 585
R1036 B.n615 B.n614 585
R1037 B.n614 B.n613 585
R1038 B.n616 B.n233 585
R1039 B.n612 B.n233 585
R1040 B.n618 B.n617 585
R1041 B.n619 B.n618 585
R1042 B.n228 B.n227 585
R1043 B.n229 B.n228 585
R1044 B.n627 B.n626 585
R1045 B.n626 B.n625 585
R1046 B.n628 B.n226 585
R1047 B.n226 B.n225 585
R1048 B.n630 B.n629 585
R1049 B.n631 B.n630 585
R1050 B.n220 B.n219 585
R1051 B.n221 B.n220 585
R1052 B.n639 B.n638 585
R1053 B.n638 B.n637 585
R1054 B.n640 B.n218 585
R1055 B.n218 B.n217 585
R1056 B.n642 B.n641 585
R1057 B.n643 B.n642 585
R1058 B.n212 B.n211 585
R1059 B.n213 B.n212 585
R1060 B.n651 B.n650 585
R1061 B.n650 B.n649 585
R1062 B.n652 B.n210 585
R1063 B.n210 B.n209 585
R1064 B.n654 B.n653 585
R1065 B.n655 B.n654 585
R1066 B.n204 B.n203 585
R1067 B.n205 B.n204 585
R1068 B.n663 B.n662 585
R1069 B.n662 B.n661 585
R1070 B.n664 B.n202 585
R1071 B.n202 B.n201 585
R1072 B.n666 B.n665 585
R1073 B.n667 B.n666 585
R1074 B.n196 B.n195 585
R1075 B.n197 B.n196 585
R1076 B.n675 B.n674 585
R1077 B.n674 B.n673 585
R1078 B.n676 B.n194 585
R1079 B.n194 B.n193 585
R1080 B.n678 B.n677 585
R1081 B.n679 B.n678 585
R1082 B.n188 B.n187 585
R1083 B.n189 B.n188 585
R1084 B.n687 B.n686 585
R1085 B.n686 B.n685 585
R1086 B.n688 B.n186 585
R1087 B.n186 B.n185 585
R1088 B.n690 B.n689 585
R1089 B.n691 B.n690 585
R1090 B.n180 B.n179 585
R1091 B.n181 B.n180 585
R1092 B.n700 B.n699 585
R1093 B.n699 B.n698 585
R1094 B.n701 B.n178 585
R1095 B.n178 B.n177 585
R1096 B.n703 B.n702 585
R1097 B.n704 B.n703 585
R1098 B.n2 B.n0 585
R1099 B.n4 B.n2 585
R1100 B.n3 B.n1 585
R1101 B.n1074 B.n3 585
R1102 B.n1072 B.n1071 585
R1103 B.n1073 B.n1072 585
R1104 B.n1070 B.n9 585
R1105 B.n9 B.n8 585
R1106 B.n1069 B.n1068 585
R1107 B.n1068 B.n1067 585
R1108 B.n11 B.n10 585
R1109 B.n1066 B.n11 585
R1110 B.n1064 B.n1063 585
R1111 B.n1065 B.n1064 585
R1112 B.n1062 B.n16 585
R1113 B.n16 B.n15 585
R1114 B.n1061 B.n1060 585
R1115 B.n1060 B.n1059 585
R1116 B.n18 B.n17 585
R1117 B.n1058 B.n18 585
R1118 B.n1056 B.n1055 585
R1119 B.n1057 B.n1056 585
R1120 B.n1054 B.n23 585
R1121 B.n23 B.n22 585
R1122 B.n1053 B.n1052 585
R1123 B.n1052 B.n1051 585
R1124 B.n25 B.n24 585
R1125 B.n1050 B.n25 585
R1126 B.n1048 B.n1047 585
R1127 B.n1049 B.n1048 585
R1128 B.n1046 B.n30 585
R1129 B.n30 B.n29 585
R1130 B.n1045 B.n1044 585
R1131 B.n1044 B.n1043 585
R1132 B.n32 B.n31 585
R1133 B.n1042 B.n32 585
R1134 B.n1040 B.n1039 585
R1135 B.n1041 B.n1040 585
R1136 B.n1038 B.n37 585
R1137 B.n37 B.n36 585
R1138 B.n1037 B.n1036 585
R1139 B.n1036 B.n1035 585
R1140 B.n39 B.n38 585
R1141 B.n1034 B.n39 585
R1142 B.n1032 B.n1031 585
R1143 B.n1033 B.n1032 585
R1144 B.n1030 B.n44 585
R1145 B.n44 B.n43 585
R1146 B.n1029 B.n1028 585
R1147 B.n1028 B.n1027 585
R1148 B.n46 B.n45 585
R1149 B.n1026 B.n46 585
R1150 B.n1024 B.n1023 585
R1151 B.n1025 B.n1024 585
R1152 B.n1022 B.n51 585
R1153 B.n51 B.n50 585
R1154 B.n1021 B.n1020 585
R1155 B.n1020 B.n1019 585
R1156 B.n53 B.n52 585
R1157 B.n1018 B.n53 585
R1158 B.n1016 B.n1015 585
R1159 B.n1017 B.n1016 585
R1160 B.n1014 B.n57 585
R1161 B.n60 B.n57 585
R1162 B.n1013 B.n1012 585
R1163 B.n1012 B.n1011 585
R1164 B.n59 B.n58 585
R1165 B.n1010 B.n59 585
R1166 B.n1008 B.n1007 585
R1167 B.n1009 B.n1008 585
R1168 B.n1006 B.n65 585
R1169 B.n65 B.n64 585
R1170 B.n1005 B.n1004 585
R1171 B.n1004 B.n1003 585
R1172 B.n67 B.n66 585
R1173 B.n1002 B.n67 585
R1174 B.n1000 B.n999 585
R1175 B.n1001 B.n1000 585
R1176 B.n998 B.n72 585
R1177 B.n72 B.n71 585
R1178 B.n997 B.n996 585
R1179 B.n996 B.n995 585
R1180 B.n74 B.n73 585
R1181 B.n994 B.n74 585
R1182 B.n992 B.n991 585
R1183 B.n993 B.n992 585
R1184 B.n990 B.n78 585
R1185 B.n81 B.n78 585
R1186 B.n989 B.n988 585
R1187 B.n988 B.n987 585
R1188 B.n80 B.n79 585
R1189 B.n986 B.n80 585
R1190 B.n984 B.n983 585
R1191 B.n985 B.n984 585
R1192 B.n982 B.n86 585
R1193 B.n86 B.n85 585
R1194 B.n981 B.n980 585
R1195 B.n980 B.n979 585
R1196 B.n88 B.n87 585
R1197 B.n978 B.n88 585
R1198 B.n976 B.n975 585
R1199 B.n977 B.n976 585
R1200 B.n974 B.n93 585
R1201 B.n93 B.n92 585
R1202 B.n973 B.n972 585
R1203 B.n972 B.n971 585
R1204 B.n95 B.n94 585
R1205 B.n970 B.n95 585
R1206 B.n968 B.n967 585
R1207 B.n969 B.n968 585
R1208 B.n966 B.n99 585
R1209 B.n102 B.n99 585
R1210 B.n965 B.n964 585
R1211 B.n964 B.n963 585
R1212 B.n101 B.n100 585
R1213 B.n962 B.n101 585
R1214 B.n960 B.n959 585
R1215 B.n961 B.n960 585
R1216 B.n958 B.n107 585
R1217 B.n107 B.n106 585
R1218 B.n957 B.n956 585
R1219 B.n956 B.n955 585
R1220 B.n109 B.n108 585
R1221 B.n954 B.n109 585
R1222 B.n952 B.n951 585
R1223 B.n953 B.n952 585
R1224 B.n950 B.n114 585
R1225 B.n114 B.n113 585
R1226 B.n949 B.n948 585
R1227 B.n948 B.n947 585
R1228 B.n116 B.n115 585
R1229 B.n946 B.n116 585
R1230 B.n944 B.n943 585
R1231 B.n945 B.n944 585
R1232 B.n942 B.n121 585
R1233 B.n121 B.n120 585
R1234 B.n941 B.n940 585
R1235 B.n940 B.n939 585
R1236 B.n123 B.n122 585
R1237 B.n938 B.n123 585
R1238 B.n936 B.n935 585
R1239 B.n937 B.n936 585
R1240 B.n934 B.n128 585
R1241 B.n128 B.n127 585
R1242 B.n933 B.n932 585
R1243 B.n932 B.n931 585
R1244 B.n130 B.n129 585
R1245 B.n930 B.n130 585
R1246 B.n928 B.n927 585
R1247 B.n929 B.n928 585
R1248 B.n926 B.n135 585
R1249 B.n135 B.n134 585
R1250 B.n925 B.n924 585
R1251 B.n924 B.n923 585
R1252 B.n137 B.n136 585
R1253 B.n922 B.n137 585
R1254 B.n920 B.n919 585
R1255 B.n921 B.n920 585
R1256 B.n1077 B.n1076 585
R1257 B.n1076 B.n1075 585
R1258 B.n471 B.n327 535.745
R1259 B.n920 B.n142 535.745
R1260 B.n473 B.n325 535.745
R1261 B.n807 B.n140 535.745
R1262 B.n808 B.n141 256.663
R1263 B.n810 B.n141 256.663
R1264 B.n816 B.n141 256.663
R1265 B.n818 B.n141 256.663
R1266 B.n824 B.n141 256.663
R1267 B.n826 B.n141 256.663
R1268 B.n832 B.n141 256.663
R1269 B.n834 B.n141 256.663
R1270 B.n840 B.n141 256.663
R1271 B.n842 B.n141 256.663
R1272 B.n848 B.n141 256.663
R1273 B.n850 B.n141 256.663
R1274 B.n857 B.n141 256.663
R1275 B.n859 B.n141 256.663
R1276 B.n865 B.n141 256.663
R1277 B.n867 B.n141 256.663
R1278 B.n873 B.n141 256.663
R1279 B.n875 B.n141 256.663
R1280 B.n881 B.n141 256.663
R1281 B.n883 B.n141 256.663
R1282 B.n889 B.n141 256.663
R1283 B.n891 B.n141 256.663
R1284 B.n897 B.n141 256.663
R1285 B.n899 B.n141 256.663
R1286 B.n905 B.n141 256.663
R1287 B.n907 B.n141 256.663
R1288 B.n913 B.n141 256.663
R1289 B.n915 B.n141 256.663
R1290 B.n466 B.n326 256.663
R1291 B.n329 B.n326 256.663
R1292 B.n459 B.n326 256.663
R1293 B.n453 B.n326 256.663
R1294 B.n451 B.n326 256.663
R1295 B.n445 B.n326 256.663
R1296 B.n443 B.n326 256.663
R1297 B.n437 B.n326 256.663
R1298 B.n435 B.n326 256.663
R1299 B.n429 B.n326 256.663
R1300 B.n427 B.n326 256.663
R1301 B.n420 B.n326 256.663
R1302 B.n418 B.n326 256.663
R1303 B.n412 B.n326 256.663
R1304 B.n410 B.n326 256.663
R1305 B.n404 B.n326 256.663
R1306 B.n349 B.n326 256.663
R1307 B.n398 B.n326 256.663
R1308 B.n392 B.n326 256.663
R1309 B.n390 B.n326 256.663
R1310 B.n384 B.n326 256.663
R1311 B.n382 B.n326 256.663
R1312 B.n376 B.n326 256.663
R1313 B.n374 B.n326 256.663
R1314 B.n368 B.n326 256.663
R1315 B.n366 B.n326 256.663
R1316 B.n360 B.n326 256.663
R1317 B.n346 B.t23 252.296
R1318 B.n162 B.t12 252.296
R1319 B.n340 B.t17 252.296
R1320 B.n155 B.t19 252.296
R1321 B.n346 B.t21 247.846
R1322 B.n340 B.t14 247.846
R1323 B.n155 B.t18 247.846
R1324 B.n162 B.t10 247.846
R1325 B.n347 B.t22 175.495
R1326 B.n163 B.t13 175.495
R1327 B.n341 B.t16 175.495
R1328 B.n156 B.t20 175.495
R1329 B.n471 B.n321 163.367
R1330 B.n479 B.n321 163.367
R1331 B.n479 B.n319 163.367
R1332 B.n483 B.n319 163.367
R1333 B.n483 B.n313 163.367
R1334 B.n491 B.n313 163.367
R1335 B.n491 B.n311 163.367
R1336 B.n495 B.n311 163.367
R1337 B.n495 B.n305 163.367
R1338 B.n503 B.n305 163.367
R1339 B.n503 B.n303 163.367
R1340 B.n507 B.n303 163.367
R1341 B.n507 B.n297 163.367
R1342 B.n515 B.n297 163.367
R1343 B.n515 B.n295 163.367
R1344 B.n519 B.n295 163.367
R1345 B.n519 B.n289 163.367
R1346 B.n527 B.n289 163.367
R1347 B.n527 B.n287 163.367
R1348 B.n531 B.n287 163.367
R1349 B.n531 B.n281 163.367
R1350 B.n540 B.n281 163.367
R1351 B.n540 B.n279 163.367
R1352 B.n544 B.n279 163.367
R1353 B.n544 B.n274 163.367
R1354 B.n552 B.n274 163.367
R1355 B.n552 B.n272 163.367
R1356 B.n556 B.n272 163.367
R1357 B.n556 B.n266 163.367
R1358 B.n564 B.n266 163.367
R1359 B.n564 B.n264 163.367
R1360 B.n568 B.n264 163.367
R1361 B.n568 B.n258 163.367
R1362 B.n577 B.n258 163.367
R1363 B.n577 B.n256 163.367
R1364 B.n581 B.n256 163.367
R1365 B.n581 B.n251 163.367
R1366 B.n589 B.n251 163.367
R1367 B.n589 B.n249 163.367
R1368 B.n593 B.n249 163.367
R1369 B.n593 B.n243 163.367
R1370 B.n601 B.n243 163.367
R1371 B.n601 B.n241 163.367
R1372 B.n605 B.n241 163.367
R1373 B.n605 B.n235 163.367
R1374 B.n614 B.n235 163.367
R1375 B.n614 B.n233 163.367
R1376 B.n618 B.n233 163.367
R1377 B.n618 B.n228 163.367
R1378 B.n626 B.n228 163.367
R1379 B.n626 B.n226 163.367
R1380 B.n630 B.n226 163.367
R1381 B.n630 B.n220 163.367
R1382 B.n638 B.n220 163.367
R1383 B.n638 B.n218 163.367
R1384 B.n642 B.n218 163.367
R1385 B.n642 B.n212 163.367
R1386 B.n650 B.n212 163.367
R1387 B.n650 B.n210 163.367
R1388 B.n654 B.n210 163.367
R1389 B.n654 B.n204 163.367
R1390 B.n662 B.n204 163.367
R1391 B.n662 B.n202 163.367
R1392 B.n666 B.n202 163.367
R1393 B.n666 B.n196 163.367
R1394 B.n674 B.n196 163.367
R1395 B.n674 B.n194 163.367
R1396 B.n678 B.n194 163.367
R1397 B.n678 B.n188 163.367
R1398 B.n686 B.n188 163.367
R1399 B.n686 B.n186 163.367
R1400 B.n690 B.n186 163.367
R1401 B.n690 B.n180 163.367
R1402 B.n699 B.n180 163.367
R1403 B.n699 B.n178 163.367
R1404 B.n703 B.n178 163.367
R1405 B.n703 B.n2 163.367
R1406 B.n1076 B.n2 163.367
R1407 B.n1076 B.n3 163.367
R1408 B.n1072 B.n3 163.367
R1409 B.n1072 B.n9 163.367
R1410 B.n1068 B.n9 163.367
R1411 B.n1068 B.n11 163.367
R1412 B.n1064 B.n11 163.367
R1413 B.n1064 B.n16 163.367
R1414 B.n1060 B.n16 163.367
R1415 B.n1060 B.n18 163.367
R1416 B.n1056 B.n18 163.367
R1417 B.n1056 B.n23 163.367
R1418 B.n1052 B.n23 163.367
R1419 B.n1052 B.n25 163.367
R1420 B.n1048 B.n25 163.367
R1421 B.n1048 B.n30 163.367
R1422 B.n1044 B.n30 163.367
R1423 B.n1044 B.n32 163.367
R1424 B.n1040 B.n32 163.367
R1425 B.n1040 B.n37 163.367
R1426 B.n1036 B.n37 163.367
R1427 B.n1036 B.n39 163.367
R1428 B.n1032 B.n39 163.367
R1429 B.n1032 B.n44 163.367
R1430 B.n1028 B.n44 163.367
R1431 B.n1028 B.n46 163.367
R1432 B.n1024 B.n46 163.367
R1433 B.n1024 B.n51 163.367
R1434 B.n1020 B.n51 163.367
R1435 B.n1020 B.n53 163.367
R1436 B.n1016 B.n53 163.367
R1437 B.n1016 B.n57 163.367
R1438 B.n1012 B.n57 163.367
R1439 B.n1012 B.n59 163.367
R1440 B.n1008 B.n59 163.367
R1441 B.n1008 B.n65 163.367
R1442 B.n1004 B.n65 163.367
R1443 B.n1004 B.n67 163.367
R1444 B.n1000 B.n67 163.367
R1445 B.n1000 B.n72 163.367
R1446 B.n996 B.n72 163.367
R1447 B.n996 B.n74 163.367
R1448 B.n992 B.n74 163.367
R1449 B.n992 B.n78 163.367
R1450 B.n988 B.n78 163.367
R1451 B.n988 B.n80 163.367
R1452 B.n984 B.n80 163.367
R1453 B.n984 B.n86 163.367
R1454 B.n980 B.n86 163.367
R1455 B.n980 B.n88 163.367
R1456 B.n976 B.n88 163.367
R1457 B.n976 B.n93 163.367
R1458 B.n972 B.n93 163.367
R1459 B.n972 B.n95 163.367
R1460 B.n968 B.n95 163.367
R1461 B.n968 B.n99 163.367
R1462 B.n964 B.n99 163.367
R1463 B.n964 B.n101 163.367
R1464 B.n960 B.n101 163.367
R1465 B.n960 B.n107 163.367
R1466 B.n956 B.n107 163.367
R1467 B.n956 B.n109 163.367
R1468 B.n952 B.n109 163.367
R1469 B.n952 B.n114 163.367
R1470 B.n948 B.n114 163.367
R1471 B.n948 B.n116 163.367
R1472 B.n944 B.n116 163.367
R1473 B.n944 B.n121 163.367
R1474 B.n940 B.n121 163.367
R1475 B.n940 B.n123 163.367
R1476 B.n936 B.n123 163.367
R1477 B.n936 B.n128 163.367
R1478 B.n932 B.n128 163.367
R1479 B.n932 B.n130 163.367
R1480 B.n928 B.n130 163.367
R1481 B.n928 B.n135 163.367
R1482 B.n924 B.n135 163.367
R1483 B.n924 B.n137 163.367
R1484 B.n920 B.n137 163.367
R1485 B.n467 B.n465 163.367
R1486 B.n465 B.n464 163.367
R1487 B.n461 B.n460 163.367
R1488 B.n458 B.n331 163.367
R1489 B.n454 B.n452 163.367
R1490 B.n450 B.n333 163.367
R1491 B.n446 B.n444 163.367
R1492 B.n442 B.n335 163.367
R1493 B.n438 B.n436 163.367
R1494 B.n434 B.n337 163.367
R1495 B.n430 B.n428 163.367
R1496 B.n426 B.n339 163.367
R1497 B.n421 B.n419 163.367
R1498 B.n417 B.n343 163.367
R1499 B.n413 B.n411 163.367
R1500 B.n409 B.n345 163.367
R1501 B.n405 B.n403 163.367
R1502 B.n400 B.n399 163.367
R1503 B.n397 B.n351 163.367
R1504 B.n393 B.n391 163.367
R1505 B.n389 B.n353 163.367
R1506 B.n385 B.n383 163.367
R1507 B.n381 B.n355 163.367
R1508 B.n377 B.n375 163.367
R1509 B.n373 B.n357 163.367
R1510 B.n369 B.n367 163.367
R1511 B.n365 B.n359 163.367
R1512 B.n361 B.n325 163.367
R1513 B.n473 B.n323 163.367
R1514 B.n477 B.n323 163.367
R1515 B.n477 B.n317 163.367
R1516 B.n485 B.n317 163.367
R1517 B.n485 B.n315 163.367
R1518 B.n489 B.n315 163.367
R1519 B.n489 B.n308 163.367
R1520 B.n497 B.n308 163.367
R1521 B.n497 B.n306 163.367
R1522 B.n501 B.n306 163.367
R1523 B.n501 B.n301 163.367
R1524 B.n509 B.n301 163.367
R1525 B.n509 B.n299 163.367
R1526 B.n513 B.n299 163.367
R1527 B.n513 B.n293 163.367
R1528 B.n521 B.n293 163.367
R1529 B.n521 B.n291 163.367
R1530 B.n525 B.n291 163.367
R1531 B.n525 B.n285 163.367
R1532 B.n533 B.n285 163.367
R1533 B.n533 B.n283 163.367
R1534 B.n537 B.n283 163.367
R1535 B.n537 B.n278 163.367
R1536 B.n546 B.n278 163.367
R1537 B.n546 B.n276 163.367
R1538 B.n550 B.n276 163.367
R1539 B.n550 B.n270 163.367
R1540 B.n558 B.n270 163.367
R1541 B.n558 B.n268 163.367
R1542 B.n562 B.n268 163.367
R1543 B.n562 B.n262 163.367
R1544 B.n570 B.n262 163.367
R1545 B.n570 B.n260 163.367
R1546 B.n574 B.n260 163.367
R1547 B.n574 B.n255 163.367
R1548 B.n583 B.n255 163.367
R1549 B.n583 B.n253 163.367
R1550 B.n587 B.n253 163.367
R1551 B.n587 B.n247 163.367
R1552 B.n595 B.n247 163.367
R1553 B.n595 B.n245 163.367
R1554 B.n599 B.n245 163.367
R1555 B.n599 B.n239 163.367
R1556 B.n607 B.n239 163.367
R1557 B.n607 B.n237 163.367
R1558 B.n611 B.n237 163.367
R1559 B.n611 B.n232 163.367
R1560 B.n620 B.n232 163.367
R1561 B.n620 B.n230 163.367
R1562 B.n624 B.n230 163.367
R1563 B.n624 B.n224 163.367
R1564 B.n632 B.n224 163.367
R1565 B.n632 B.n222 163.367
R1566 B.n636 B.n222 163.367
R1567 B.n636 B.n216 163.367
R1568 B.n644 B.n216 163.367
R1569 B.n644 B.n214 163.367
R1570 B.n648 B.n214 163.367
R1571 B.n648 B.n208 163.367
R1572 B.n656 B.n208 163.367
R1573 B.n656 B.n206 163.367
R1574 B.n660 B.n206 163.367
R1575 B.n660 B.n200 163.367
R1576 B.n668 B.n200 163.367
R1577 B.n668 B.n198 163.367
R1578 B.n672 B.n198 163.367
R1579 B.n672 B.n192 163.367
R1580 B.n680 B.n192 163.367
R1581 B.n680 B.n190 163.367
R1582 B.n684 B.n190 163.367
R1583 B.n684 B.n184 163.367
R1584 B.n692 B.n184 163.367
R1585 B.n692 B.n182 163.367
R1586 B.n697 B.n182 163.367
R1587 B.n697 B.n176 163.367
R1588 B.n705 B.n176 163.367
R1589 B.n706 B.n705 163.367
R1590 B.n706 B.n5 163.367
R1591 B.n6 B.n5 163.367
R1592 B.n7 B.n6 163.367
R1593 B.n711 B.n7 163.367
R1594 B.n711 B.n12 163.367
R1595 B.n13 B.n12 163.367
R1596 B.n14 B.n13 163.367
R1597 B.n716 B.n14 163.367
R1598 B.n716 B.n19 163.367
R1599 B.n20 B.n19 163.367
R1600 B.n21 B.n20 163.367
R1601 B.n721 B.n21 163.367
R1602 B.n721 B.n26 163.367
R1603 B.n27 B.n26 163.367
R1604 B.n28 B.n27 163.367
R1605 B.n726 B.n28 163.367
R1606 B.n726 B.n33 163.367
R1607 B.n34 B.n33 163.367
R1608 B.n35 B.n34 163.367
R1609 B.n731 B.n35 163.367
R1610 B.n731 B.n40 163.367
R1611 B.n41 B.n40 163.367
R1612 B.n42 B.n41 163.367
R1613 B.n736 B.n42 163.367
R1614 B.n736 B.n47 163.367
R1615 B.n48 B.n47 163.367
R1616 B.n49 B.n48 163.367
R1617 B.n741 B.n49 163.367
R1618 B.n741 B.n54 163.367
R1619 B.n55 B.n54 163.367
R1620 B.n56 B.n55 163.367
R1621 B.n746 B.n56 163.367
R1622 B.n746 B.n61 163.367
R1623 B.n62 B.n61 163.367
R1624 B.n63 B.n62 163.367
R1625 B.n751 B.n63 163.367
R1626 B.n751 B.n68 163.367
R1627 B.n69 B.n68 163.367
R1628 B.n70 B.n69 163.367
R1629 B.n756 B.n70 163.367
R1630 B.n756 B.n75 163.367
R1631 B.n76 B.n75 163.367
R1632 B.n77 B.n76 163.367
R1633 B.n761 B.n77 163.367
R1634 B.n761 B.n82 163.367
R1635 B.n83 B.n82 163.367
R1636 B.n84 B.n83 163.367
R1637 B.n766 B.n84 163.367
R1638 B.n766 B.n89 163.367
R1639 B.n90 B.n89 163.367
R1640 B.n91 B.n90 163.367
R1641 B.n771 B.n91 163.367
R1642 B.n771 B.n96 163.367
R1643 B.n97 B.n96 163.367
R1644 B.n98 B.n97 163.367
R1645 B.n776 B.n98 163.367
R1646 B.n776 B.n103 163.367
R1647 B.n104 B.n103 163.367
R1648 B.n105 B.n104 163.367
R1649 B.n781 B.n105 163.367
R1650 B.n781 B.n110 163.367
R1651 B.n111 B.n110 163.367
R1652 B.n112 B.n111 163.367
R1653 B.n786 B.n112 163.367
R1654 B.n786 B.n117 163.367
R1655 B.n118 B.n117 163.367
R1656 B.n119 B.n118 163.367
R1657 B.n791 B.n119 163.367
R1658 B.n791 B.n124 163.367
R1659 B.n125 B.n124 163.367
R1660 B.n126 B.n125 163.367
R1661 B.n796 B.n126 163.367
R1662 B.n796 B.n131 163.367
R1663 B.n132 B.n131 163.367
R1664 B.n133 B.n132 163.367
R1665 B.n801 B.n133 163.367
R1666 B.n801 B.n138 163.367
R1667 B.n139 B.n138 163.367
R1668 B.n140 B.n139 163.367
R1669 B.n916 B.n914 163.367
R1670 B.n912 B.n144 163.367
R1671 B.n908 B.n906 163.367
R1672 B.n904 B.n146 163.367
R1673 B.n900 B.n898 163.367
R1674 B.n896 B.n148 163.367
R1675 B.n892 B.n890 163.367
R1676 B.n888 B.n150 163.367
R1677 B.n884 B.n882 163.367
R1678 B.n880 B.n152 163.367
R1679 B.n876 B.n874 163.367
R1680 B.n872 B.n154 163.367
R1681 B.n868 B.n866 163.367
R1682 B.n864 B.n159 163.367
R1683 B.n860 B.n858 163.367
R1684 B.n856 B.n161 163.367
R1685 B.n851 B.n849 163.367
R1686 B.n847 B.n165 163.367
R1687 B.n843 B.n841 163.367
R1688 B.n839 B.n167 163.367
R1689 B.n835 B.n833 163.367
R1690 B.n831 B.n169 163.367
R1691 B.n827 B.n825 163.367
R1692 B.n823 B.n171 163.367
R1693 B.n819 B.n817 163.367
R1694 B.n815 B.n173 163.367
R1695 B.n811 B.n809 163.367
R1696 B.n472 B.n326 121.948
R1697 B.n921 B.n141 121.948
R1698 B.n347 B.n346 76.8005
R1699 B.n341 B.n340 76.8005
R1700 B.n156 B.n155 76.8005
R1701 B.n163 B.n162 76.8005
R1702 B.n466 B.n327 71.676
R1703 B.n464 B.n329 71.676
R1704 B.n460 B.n459 71.676
R1705 B.n453 B.n331 71.676
R1706 B.n452 B.n451 71.676
R1707 B.n445 B.n333 71.676
R1708 B.n444 B.n443 71.676
R1709 B.n437 B.n335 71.676
R1710 B.n436 B.n435 71.676
R1711 B.n429 B.n337 71.676
R1712 B.n428 B.n427 71.676
R1713 B.n420 B.n339 71.676
R1714 B.n419 B.n418 71.676
R1715 B.n412 B.n343 71.676
R1716 B.n411 B.n410 71.676
R1717 B.n404 B.n345 71.676
R1718 B.n403 B.n349 71.676
R1719 B.n399 B.n398 71.676
R1720 B.n392 B.n351 71.676
R1721 B.n391 B.n390 71.676
R1722 B.n384 B.n353 71.676
R1723 B.n383 B.n382 71.676
R1724 B.n376 B.n355 71.676
R1725 B.n375 B.n374 71.676
R1726 B.n368 B.n357 71.676
R1727 B.n367 B.n366 71.676
R1728 B.n360 B.n359 71.676
R1729 B.n915 B.n142 71.676
R1730 B.n914 B.n913 71.676
R1731 B.n907 B.n144 71.676
R1732 B.n906 B.n905 71.676
R1733 B.n899 B.n146 71.676
R1734 B.n898 B.n897 71.676
R1735 B.n891 B.n148 71.676
R1736 B.n890 B.n889 71.676
R1737 B.n883 B.n150 71.676
R1738 B.n882 B.n881 71.676
R1739 B.n875 B.n152 71.676
R1740 B.n874 B.n873 71.676
R1741 B.n867 B.n154 71.676
R1742 B.n866 B.n865 71.676
R1743 B.n859 B.n159 71.676
R1744 B.n858 B.n857 71.676
R1745 B.n850 B.n161 71.676
R1746 B.n849 B.n848 71.676
R1747 B.n842 B.n165 71.676
R1748 B.n841 B.n840 71.676
R1749 B.n834 B.n167 71.676
R1750 B.n833 B.n832 71.676
R1751 B.n826 B.n169 71.676
R1752 B.n825 B.n824 71.676
R1753 B.n818 B.n171 71.676
R1754 B.n817 B.n816 71.676
R1755 B.n810 B.n173 71.676
R1756 B.n809 B.n808 71.676
R1757 B.n808 B.n807 71.676
R1758 B.n811 B.n810 71.676
R1759 B.n816 B.n815 71.676
R1760 B.n819 B.n818 71.676
R1761 B.n824 B.n823 71.676
R1762 B.n827 B.n826 71.676
R1763 B.n832 B.n831 71.676
R1764 B.n835 B.n834 71.676
R1765 B.n840 B.n839 71.676
R1766 B.n843 B.n842 71.676
R1767 B.n848 B.n847 71.676
R1768 B.n851 B.n850 71.676
R1769 B.n857 B.n856 71.676
R1770 B.n860 B.n859 71.676
R1771 B.n865 B.n864 71.676
R1772 B.n868 B.n867 71.676
R1773 B.n873 B.n872 71.676
R1774 B.n876 B.n875 71.676
R1775 B.n881 B.n880 71.676
R1776 B.n884 B.n883 71.676
R1777 B.n889 B.n888 71.676
R1778 B.n892 B.n891 71.676
R1779 B.n897 B.n896 71.676
R1780 B.n900 B.n899 71.676
R1781 B.n905 B.n904 71.676
R1782 B.n908 B.n907 71.676
R1783 B.n913 B.n912 71.676
R1784 B.n916 B.n915 71.676
R1785 B.n467 B.n466 71.676
R1786 B.n461 B.n329 71.676
R1787 B.n459 B.n458 71.676
R1788 B.n454 B.n453 71.676
R1789 B.n451 B.n450 71.676
R1790 B.n446 B.n445 71.676
R1791 B.n443 B.n442 71.676
R1792 B.n438 B.n437 71.676
R1793 B.n435 B.n434 71.676
R1794 B.n430 B.n429 71.676
R1795 B.n427 B.n426 71.676
R1796 B.n421 B.n420 71.676
R1797 B.n418 B.n417 71.676
R1798 B.n413 B.n412 71.676
R1799 B.n410 B.n409 71.676
R1800 B.n405 B.n404 71.676
R1801 B.n400 B.n349 71.676
R1802 B.n398 B.n397 71.676
R1803 B.n393 B.n392 71.676
R1804 B.n390 B.n389 71.676
R1805 B.n385 B.n384 71.676
R1806 B.n382 B.n381 71.676
R1807 B.n377 B.n376 71.676
R1808 B.n374 B.n373 71.676
R1809 B.n369 B.n368 71.676
R1810 B.n366 B.n365 71.676
R1811 B.n361 B.n360 71.676
R1812 B.n472 B.n322 67.4183
R1813 B.n478 B.n322 67.4183
R1814 B.n478 B.n318 67.4183
R1815 B.n484 B.n318 67.4183
R1816 B.n484 B.n314 67.4183
R1817 B.n490 B.n314 67.4183
R1818 B.n490 B.n309 67.4183
R1819 B.n496 B.n309 67.4183
R1820 B.n496 B.n310 67.4183
R1821 B.n502 B.n302 67.4183
R1822 B.n508 B.n302 67.4183
R1823 B.n508 B.n298 67.4183
R1824 B.n514 B.n298 67.4183
R1825 B.n514 B.n294 67.4183
R1826 B.n520 B.n294 67.4183
R1827 B.n520 B.n290 67.4183
R1828 B.n526 B.n290 67.4183
R1829 B.n526 B.n286 67.4183
R1830 B.n532 B.n286 67.4183
R1831 B.n532 B.n282 67.4183
R1832 B.n539 B.n282 67.4183
R1833 B.n539 B.n538 67.4183
R1834 B.n545 B.n275 67.4183
R1835 B.n551 B.n275 67.4183
R1836 B.n551 B.n271 67.4183
R1837 B.n557 B.n271 67.4183
R1838 B.n557 B.n267 67.4183
R1839 B.n563 B.n267 67.4183
R1840 B.n563 B.n263 67.4183
R1841 B.n569 B.n263 67.4183
R1842 B.n569 B.n259 67.4183
R1843 B.n576 B.n259 67.4183
R1844 B.n576 B.n575 67.4183
R1845 B.n582 B.n252 67.4183
R1846 B.n588 B.n252 67.4183
R1847 B.n588 B.n248 67.4183
R1848 B.n594 B.n248 67.4183
R1849 B.n594 B.n244 67.4183
R1850 B.n600 B.n244 67.4183
R1851 B.n600 B.n240 67.4183
R1852 B.n606 B.n240 67.4183
R1853 B.n606 B.n236 67.4183
R1854 B.n613 B.n236 67.4183
R1855 B.n613 B.n612 67.4183
R1856 B.n619 B.n229 67.4183
R1857 B.n625 B.n229 67.4183
R1858 B.n625 B.n225 67.4183
R1859 B.n631 B.n225 67.4183
R1860 B.n631 B.n221 67.4183
R1861 B.n637 B.n221 67.4183
R1862 B.n637 B.n217 67.4183
R1863 B.n643 B.n217 67.4183
R1864 B.n643 B.n213 67.4183
R1865 B.n649 B.n213 67.4183
R1866 B.n655 B.n209 67.4183
R1867 B.n655 B.n205 67.4183
R1868 B.n661 B.n205 67.4183
R1869 B.n661 B.n201 67.4183
R1870 B.n667 B.n201 67.4183
R1871 B.n667 B.n197 67.4183
R1872 B.n673 B.n197 67.4183
R1873 B.n673 B.n193 67.4183
R1874 B.n679 B.n193 67.4183
R1875 B.n679 B.n189 67.4183
R1876 B.n685 B.n189 67.4183
R1877 B.n691 B.n185 67.4183
R1878 B.n691 B.n181 67.4183
R1879 B.n698 B.n181 67.4183
R1880 B.n698 B.n177 67.4183
R1881 B.n704 B.n177 67.4183
R1882 B.n704 B.n4 67.4183
R1883 B.n1075 B.n4 67.4183
R1884 B.n1075 B.n1074 67.4183
R1885 B.n1074 B.n1073 67.4183
R1886 B.n1073 B.n8 67.4183
R1887 B.n1067 B.n8 67.4183
R1888 B.n1067 B.n1066 67.4183
R1889 B.n1066 B.n1065 67.4183
R1890 B.n1065 B.n15 67.4183
R1891 B.n1059 B.n1058 67.4183
R1892 B.n1058 B.n1057 67.4183
R1893 B.n1057 B.n22 67.4183
R1894 B.n1051 B.n22 67.4183
R1895 B.n1051 B.n1050 67.4183
R1896 B.n1050 B.n1049 67.4183
R1897 B.n1049 B.n29 67.4183
R1898 B.n1043 B.n29 67.4183
R1899 B.n1043 B.n1042 67.4183
R1900 B.n1042 B.n1041 67.4183
R1901 B.n1041 B.n36 67.4183
R1902 B.n1035 B.n1034 67.4183
R1903 B.n1034 B.n1033 67.4183
R1904 B.n1033 B.n43 67.4183
R1905 B.n1027 B.n43 67.4183
R1906 B.n1027 B.n1026 67.4183
R1907 B.n1026 B.n1025 67.4183
R1908 B.n1025 B.n50 67.4183
R1909 B.n1019 B.n50 67.4183
R1910 B.n1019 B.n1018 67.4183
R1911 B.n1018 B.n1017 67.4183
R1912 B.n1011 B.n60 67.4183
R1913 B.n1011 B.n1010 67.4183
R1914 B.n1010 B.n1009 67.4183
R1915 B.n1009 B.n64 67.4183
R1916 B.n1003 B.n64 67.4183
R1917 B.n1003 B.n1002 67.4183
R1918 B.n1002 B.n1001 67.4183
R1919 B.n1001 B.n71 67.4183
R1920 B.n995 B.n71 67.4183
R1921 B.n995 B.n994 67.4183
R1922 B.n994 B.n993 67.4183
R1923 B.n987 B.n81 67.4183
R1924 B.n987 B.n986 67.4183
R1925 B.n986 B.n985 67.4183
R1926 B.n985 B.n85 67.4183
R1927 B.n979 B.n85 67.4183
R1928 B.n979 B.n978 67.4183
R1929 B.n978 B.n977 67.4183
R1930 B.n977 B.n92 67.4183
R1931 B.n971 B.n92 67.4183
R1932 B.n971 B.n970 67.4183
R1933 B.n970 B.n969 67.4183
R1934 B.n963 B.n102 67.4183
R1935 B.n963 B.n962 67.4183
R1936 B.n962 B.n961 67.4183
R1937 B.n961 B.n106 67.4183
R1938 B.n955 B.n106 67.4183
R1939 B.n955 B.n954 67.4183
R1940 B.n954 B.n953 67.4183
R1941 B.n953 B.n113 67.4183
R1942 B.n947 B.n113 67.4183
R1943 B.n947 B.n946 67.4183
R1944 B.n946 B.n945 67.4183
R1945 B.n945 B.n120 67.4183
R1946 B.n939 B.n120 67.4183
R1947 B.n938 B.n937 67.4183
R1948 B.n937 B.n127 67.4183
R1949 B.n931 B.n127 67.4183
R1950 B.n931 B.n930 67.4183
R1951 B.n930 B.n929 67.4183
R1952 B.n929 B.n134 67.4183
R1953 B.n923 B.n134 67.4183
R1954 B.n923 B.n922 67.4183
R1955 B.n922 B.n921 67.4183
R1956 B.n538 B.t3 66.4268
R1957 B.n102 B.t7 66.4268
R1958 B.n649 B.t8 62.4611
R1959 B.n1035 B.t6 62.4611
R1960 B.n348 B.n347 59.5399
R1961 B.n424 B.n341 59.5399
R1962 B.n157 B.n156 59.5399
R1963 B.n853 B.n163 59.5399
R1964 B.n502 B.t15 58.4953
R1965 B.n939 B.t11 58.4953
R1966 B.n619 B.t0 48.5809
R1967 B.n1017 B.t1 48.5809
R1968 B.n575 B.t2 42.6323
R1969 B.n81 B.t9 42.6323
R1970 B.n685 B.t4 38.6666
R1971 B.n1059 B.t5 38.6666
R1972 B.n919 B.n918 34.8103
R1973 B.n806 B.n805 34.8103
R1974 B.n474 B.n324 34.8103
R1975 B.n470 B.n469 34.8103
R1976 B.t4 B.n185 28.7522
R1977 B.t5 B.n15 28.7522
R1978 B.n582 B.t2 24.7864
R1979 B.n993 B.t9 24.7864
R1980 B.n612 B.t0 18.8378
R1981 B.n60 B.t1 18.8378
R1982 B B.n1077 18.0485
R1983 B.n918 B.n917 10.6151
R1984 B.n917 B.n143 10.6151
R1985 B.n911 B.n143 10.6151
R1986 B.n911 B.n910 10.6151
R1987 B.n910 B.n909 10.6151
R1988 B.n909 B.n145 10.6151
R1989 B.n903 B.n145 10.6151
R1990 B.n903 B.n902 10.6151
R1991 B.n902 B.n901 10.6151
R1992 B.n901 B.n147 10.6151
R1993 B.n895 B.n147 10.6151
R1994 B.n895 B.n894 10.6151
R1995 B.n894 B.n893 10.6151
R1996 B.n893 B.n149 10.6151
R1997 B.n887 B.n149 10.6151
R1998 B.n887 B.n886 10.6151
R1999 B.n886 B.n885 10.6151
R2000 B.n885 B.n151 10.6151
R2001 B.n879 B.n151 10.6151
R2002 B.n879 B.n878 10.6151
R2003 B.n878 B.n877 10.6151
R2004 B.n877 B.n153 10.6151
R2005 B.n871 B.n870 10.6151
R2006 B.n870 B.n869 10.6151
R2007 B.n869 B.n158 10.6151
R2008 B.n863 B.n158 10.6151
R2009 B.n863 B.n862 10.6151
R2010 B.n862 B.n861 10.6151
R2011 B.n861 B.n160 10.6151
R2012 B.n855 B.n160 10.6151
R2013 B.n855 B.n854 10.6151
R2014 B.n852 B.n164 10.6151
R2015 B.n846 B.n164 10.6151
R2016 B.n846 B.n845 10.6151
R2017 B.n845 B.n844 10.6151
R2018 B.n844 B.n166 10.6151
R2019 B.n838 B.n166 10.6151
R2020 B.n838 B.n837 10.6151
R2021 B.n837 B.n836 10.6151
R2022 B.n836 B.n168 10.6151
R2023 B.n830 B.n168 10.6151
R2024 B.n830 B.n829 10.6151
R2025 B.n829 B.n828 10.6151
R2026 B.n828 B.n170 10.6151
R2027 B.n822 B.n170 10.6151
R2028 B.n822 B.n821 10.6151
R2029 B.n821 B.n820 10.6151
R2030 B.n820 B.n172 10.6151
R2031 B.n814 B.n172 10.6151
R2032 B.n814 B.n813 10.6151
R2033 B.n813 B.n812 10.6151
R2034 B.n812 B.n174 10.6151
R2035 B.n806 B.n174 10.6151
R2036 B.n475 B.n474 10.6151
R2037 B.n476 B.n475 10.6151
R2038 B.n476 B.n316 10.6151
R2039 B.n486 B.n316 10.6151
R2040 B.n487 B.n486 10.6151
R2041 B.n488 B.n487 10.6151
R2042 B.n488 B.n307 10.6151
R2043 B.n498 B.n307 10.6151
R2044 B.n499 B.n498 10.6151
R2045 B.n500 B.n499 10.6151
R2046 B.n500 B.n300 10.6151
R2047 B.n510 B.n300 10.6151
R2048 B.n511 B.n510 10.6151
R2049 B.n512 B.n511 10.6151
R2050 B.n512 B.n292 10.6151
R2051 B.n522 B.n292 10.6151
R2052 B.n523 B.n522 10.6151
R2053 B.n524 B.n523 10.6151
R2054 B.n524 B.n284 10.6151
R2055 B.n534 B.n284 10.6151
R2056 B.n535 B.n534 10.6151
R2057 B.n536 B.n535 10.6151
R2058 B.n536 B.n277 10.6151
R2059 B.n547 B.n277 10.6151
R2060 B.n548 B.n547 10.6151
R2061 B.n549 B.n548 10.6151
R2062 B.n549 B.n269 10.6151
R2063 B.n559 B.n269 10.6151
R2064 B.n560 B.n559 10.6151
R2065 B.n561 B.n560 10.6151
R2066 B.n561 B.n261 10.6151
R2067 B.n571 B.n261 10.6151
R2068 B.n572 B.n571 10.6151
R2069 B.n573 B.n572 10.6151
R2070 B.n573 B.n254 10.6151
R2071 B.n584 B.n254 10.6151
R2072 B.n585 B.n584 10.6151
R2073 B.n586 B.n585 10.6151
R2074 B.n586 B.n246 10.6151
R2075 B.n596 B.n246 10.6151
R2076 B.n597 B.n596 10.6151
R2077 B.n598 B.n597 10.6151
R2078 B.n598 B.n238 10.6151
R2079 B.n608 B.n238 10.6151
R2080 B.n609 B.n608 10.6151
R2081 B.n610 B.n609 10.6151
R2082 B.n610 B.n231 10.6151
R2083 B.n621 B.n231 10.6151
R2084 B.n622 B.n621 10.6151
R2085 B.n623 B.n622 10.6151
R2086 B.n623 B.n223 10.6151
R2087 B.n633 B.n223 10.6151
R2088 B.n634 B.n633 10.6151
R2089 B.n635 B.n634 10.6151
R2090 B.n635 B.n215 10.6151
R2091 B.n645 B.n215 10.6151
R2092 B.n646 B.n645 10.6151
R2093 B.n647 B.n646 10.6151
R2094 B.n647 B.n207 10.6151
R2095 B.n657 B.n207 10.6151
R2096 B.n658 B.n657 10.6151
R2097 B.n659 B.n658 10.6151
R2098 B.n659 B.n199 10.6151
R2099 B.n669 B.n199 10.6151
R2100 B.n670 B.n669 10.6151
R2101 B.n671 B.n670 10.6151
R2102 B.n671 B.n191 10.6151
R2103 B.n681 B.n191 10.6151
R2104 B.n682 B.n681 10.6151
R2105 B.n683 B.n682 10.6151
R2106 B.n683 B.n183 10.6151
R2107 B.n693 B.n183 10.6151
R2108 B.n694 B.n693 10.6151
R2109 B.n696 B.n694 10.6151
R2110 B.n696 B.n695 10.6151
R2111 B.n695 B.n175 10.6151
R2112 B.n707 B.n175 10.6151
R2113 B.n708 B.n707 10.6151
R2114 B.n709 B.n708 10.6151
R2115 B.n710 B.n709 10.6151
R2116 B.n712 B.n710 10.6151
R2117 B.n713 B.n712 10.6151
R2118 B.n714 B.n713 10.6151
R2119 B.n715 B.n714 10.6151
R2120 B.n717 B.n715 10.6151
R2121 B.n718 B.n717 10.6151
R2122 B.n719 B.n718 10.6151
R2123 B.n720 B.n719 10.6151
R2124 B.n722 B.n720 10.6151
R2125 B.n723 B.n722 10.6151
R2126 B.n724 B.n723 10.6151
R2127 B.n725 B.n724 10.6151
R2128 B.n727 B.n725 10.6151
R2129 B.n728 B.n727 10.6151
R2130 B.n729 B.n728 10.6151
R2131 B.n730 B.n729 10.6151
R2132 B.n732 B.n730 10.6151
R2133 B.n733 B.n732 10.6151
R2134 B.n734 B.n733 10.6151
R2135 B.n735 B.n734 10.6151
R2136 B.n737 B.n735 10.6151
R2137 B.n738 B.n737 10.6151
R2138 B.n739 B.n738 10.6151
R2139 B.n740 B.n739 10.6151
R2140 B.n742 B.n740 10.6151
R2141 B.n743 B.n742 10.6151
R2142 B.n744 B.n743 10.6151
R2143 B.n745 B.n744 10.6151
R2144 B.n747 B.n745 10.6151
R2145 B.n748 B.n747 10.6151
R2146 B.n749 B.n748 10.6151
R2147 B.n750 B.n749 10.6151
R2148 B.n752 B.n750 10.6151
R2149 B.n753 B.n752 10.6151
R2150 B.n754 B.n753 10.6151
R2151 B.n755 B.n754 10.6151
R2152 B.n757 B.n755 10.6151
R2153 B.n758 B.n757 10.6151
R2154 B.n759 B.n758 10.6151
R2155 B.n760 B.n759 10.6151
R2156 B.n762 B.n760 10.6151
R2157 B.n763 B.n762 10.6151
R2158 B.n764 B.n763 10.6151
R2159 B.n765 B.n764 10.6151
R2160 B.n767 B.n765 10.6151
R2161 B.n768 B.n767 10.6151
R2162 B.n769 B.n768 10.6151
R2163 B.n770 B.n769 10.6151
R2164 B.n772 B.n770 10.6151
R2165 B.n773 B.n772 10.6151
R2166 B.n774 B.n773 10.6151
R2167 B.n775 B.n774 10.6151
R2168 B.n777 B.n775 10.6151
R2169 B.n778 B.n777 10.6151
R2170 B.n779 B.n778 10.6151
R2171 B.n780 B.n779 10.6151
R2172 B.n782 B.n780 10.6151
R2173 B.n783 B.n782 10.6151
R2174 B.n784 B.n783 10.6151
R2175 B.n785 B.n784 10.6151
R2176 B.n787 B.n785 10.6151
R2177 B.n788 B.n787 10.6151
R2178 B.n789 B.n788 10.6151
R2179 B.n790 B.n789 10.6151
R2180 B.n792 B.n790 10.6151
R2181 B.n793 B.n792 10.6151
R2182 B.n794 B.n793 10.6151
R2183 B.n795 B.n794 10.6151
R2184 B.n797 B.n795 10.6151
R2185 B.n798 B.n797 10.6151
R2186 B.n799 B.n798 10.6151
R2187 B.n800 B.n799 10.6151
R2188 B.n802 B.n800 10.6151
R2189 B.n803 B.n802 10.6151
R2190 B.n804 B.n803 10.6151
R2191 B.n805 B.n804 10.6151
R2192 B.n469 B.n468 10.6151
R2193 B.n468 B.n328 10.6151
R2194 B.n463 B.n328 10.6151
R2195 B.n463 B.n462 10.6151
R2196 B.n462 B.n330 10.6151
R2197 B.n457 B.n330 10.6151
R2198 B.n457 B.n456 10.6151
R2199 B.n456 B.n455 10.6151
R2200 B.n455 B.n332 10.6151
R2201 B.n449 B.n332 10.6151
R2202 B.n449 B.n448 10.6151
R2203 B.n448 B.n447 10.6151
R2204 B.n447 B.n334 10.6151
R2205 B.n441 B.n334 10.6151
R2206 B.n441 B.n440 10.6151
R2207 B.n440 B.n439 10.6151
R2208 B.n439 B.n336 10.6151
R2209 B.n433 B.n336 10.6151
R2210 B.n433 B.n432 10.6151
R2211 B.n432 B.n431 10.6151
R2212 B.n431 B.n338 10.6151
R2213 B.n425 B.n338 10.6151
R2214 B.n423 B.n422 10.6151
R2215 B.n422 B.n342 10.6151
R2216 B.n416 B.n342 10.6151
R2217 B.n416 B.n415 10.6151
R2218 B.n415 B.n414 10.6151
R2219 B.n414 B.n344 10.6151
R2220 B.n408 B.n344 10.6151
R2221 B.n408 B.n407 10.6151
R2222 B.n407 B.n406 10.6151
R2223 B.n402 B.n401 10.6151
R2224 B.n401 B.n350 10.6151
R2225 B.n396 B.n350 10.6151
R2226 B.n396 B.n395 10.6151
R2227 B.n395 B.n394 10.6151
R2228 B.n394 B.n352 10.6151
R2229 B.n388 B.n352 10.6151
R2230 B.n388 B.n387 10.6151
R2231 B.n387 B.n386 10.6151
R2232 B.n386 B.n354 10.6151
R2233 B.n380 B.n354 10.6151
R2234 B.n380 B.n379 10.6151
R2235 B.n379 B.n378 10.6151
R2236 B.n378 B.n356 10.6151
R2237 B.n372 B.n356 10.6151
R2238 B.n372 B.n371 10.6151
R2239 B.n371 B.n370 10.6151
R2240 B.n370 B.n358 10.6151
R2241 B.n364 B.n358 10.6151
R2242 B.n364 B.n363 10.6151
R2243 B.n363 B.n362 10.6151
R2244 B.n362 B.n324 10.6151
R2245 B.n470 B.n320 10.6151
R2246 B.n480 B.n320 10.6151
R2247 B.n481 B.n480 10.6151
R2248 B.n482 B.n481 10.6151
R2249 B.n482 B.n312 10.6151
R2250 B.n492 B.n312 10.6151
R2251 B.n493 B.n492 10.6151
R2252 B.n494 B.n493 10.6151
R2253 B.n494 B.n304 10.6151
R2254 B.n504 B.n304 10.6151
R2255 B.n505 B.n504 10.6151
R2256 B.n506 B.n505 10.6151
R2257 B.n506 B.n296 10.6151
R2258 B.n516 B.n296 10.6151
R2259 B.n517 B.n516 10.6151
R2260 B.n518 B.n517 10.6151
R2261 B.n518 B.n288 10.6151
R2262 B.n528 B.n288 10.6151
R2263 B.n529 B.n528 10.6151
R2264 B.n530 B.n529 10.6151
R2265 B.n530 B.n280 10.6151
R2266 B.n541 B.n280 10.6151
R2267 B.n542 B.n541 10.6151
R2268 B.n543 B.n542 10.6151
R2269 B.n543 B.n273 10.6151
R2270 B.n553 B.n273 10.6151
R2271 B.n554 B.n553 10.6151
R2272 B.n555 B.n554 10.6151
R2273 B.n555 B.n265 10.6151
R2274 B.n565 B.n265 10.6151
R2275 B.n566 B.n565 10.6151
R2276 B.n567 B.n566 10.6151
R2277 B.n567 B.n257 10.6151
R2278 B.n578 B.n257 10.6151
R2279 B.n579 B.n578 10.6151
R2280 B.n580 B.n579 10.6151
R2281 B.n580 B.n250 10.6151
R2282 B.n590 B.n250 10.6151
R2283 B.n591 B.n590 10.6151
R2284 B.n592 B.n591 10.6151
R2285 B.n592 B.n242 10.6151
R2286 B.n602 B.n242 10.6151
R2287 B.n603 B.n602 10.6151
R2288 B.n604 B.n603 10.6151
R2289 B.n604 B.n234 10.6151
R2290 B.n615 B.n234 10.6151
R2291 B.n616 B.n615 10.6151
R2292 B.n617 B.n616 10.6151
R2293 B.n617 B.n227 10.6151
R2294 B.n627 B.n227 10.6151
R2295 B.n628 B.n627 10.6151
R2296 B.n629 B.n628 10.6151
R2297 B.n629 B.n219 10.6151
R2298 B.n639 B.n219 10.6151
R2299 B.n640 B.n639 10.6151
R2300 B.n641 B.n640 10.6151
R2301 B.n641 B.n211 10.6151
R2302 B.n651 B.n211 10.6151
R2303 B.n652 B.n651 10.6151
R2304 B.n653 B.n652 10.6151
R2305 B.n653 B.n203 10.6151
R2306 B.n663 B.n203 10.6151
R2307 B.n664 B.n663 10.6151
R2308 B.n665 B.n664 10.6151
R2309 B.n665 B.n195 10.6151
R2310 B.n675 B.n195 10.6151
R2311 B.n676 B.n675 10.6151
R2312 B.n677 B.n676 10.6151
R2313 B.n677 B.n187 10.6151
R2314 B.n687 B.n187 10.6151
R2315 B.n688 B.n687 10.6151
R2316 B.n689 B.n688 10.6151
R2317 B.n689 B.n179 10.6151
R2318 B.n700 B.n179 10.6151
R2319 B.n701 B.n700 10.6151
R2320 B.n702 B.n701 10.6151
R2321 B.n702 B.n0 10.6151
R2322 B.n1071 B.n1 10.6151
R2323 B.n1071 B.n1070 10.6151
R2324 B.n1070 B.n1069 10.6151
R2325 B.n1069 B.n10 10.6151
R2326 B.n1063 B.n10 10.6151
R2327 B.n1063 B.n1062 10.6151
R2328 B.n1062 B.n1061 10.6151
R2329 B.n1061 B.n17 10.6151
R2330 B.n1055 B.n17 10.6151
R2331 B.n1055 B.n1054 10.6151
R2332 B.n1054 B.n1053 10.6151
R2333 B.n1053 B.n24 10.6151
R2334 B.n1047 B.n24 10.6151
R2335 B.n1047 B.n1046 10.6151
R2336 B.n1046 B.n1045 10.6151
R2337 B.n1045 B.n31 10.6151
R2338 B.n1039 B.n31 10.6151
R2339 B.n1039 B.n1038 10.6151
R2340 B.n1038 B.n1037 10.6151
R2341 B.n1037 B.n38 10.6151
R2342 B.n1031 B.n38 10.6151
R2343 B.n1031 B.n1030 10.6151
R2344 B.n1030 B.n1029 10.6151
R2345 B.n1029 B.n45 10.6151
R2346 B.n1023 B.n45 10.6151
R2347 B.n1023 B.n1022 10.6151
R2348 B.n1022 B.n1021 10.6151
R2349 B.n1021 B.n52 10.6151
R2350 B.n1015 B.n52 10.6151
R2351 B.n1015 B.n1014 10.6151
R2352 B.n1014 B.n1013 10.6151
R2353 B.n1013 B.n58 10.6151
R2354 B.n1007 B.n58 10.6151
R2355 B.n1007 B.n1006 10.6151
R2356 B.n1006 B.n1005 10.6151
R2357 B.n1005 B.n66 10.6151
R2358 B.n999 B.n66 10.6151
R2359 B.n999 B.n998 10.6151
R2360 B.n998 B.n997 10.6151
R2361 B.n997 B.n73 10.6151
R2362 B.n991 B.n73 10.6151
R2363 B.n991 B.n990 10.6151
R2364 B.n990 B.n989 10.6151
R2365 B.n989 B.n79 10.6151
R2366 B.n983 B.n79 10.6151
R2367 B.n983 B.n982 10.6151
R2368 B.n982 B.n981 10.6151
R2369 B.n981 B.n87 10.6151
R2370 B.n975 B.n87 10.6151
R2371 B.n975 B.n974 10.6151
R2372 B.n974 B.n973 10.6151
R2373 B.n973 B.n94 10.6151
R2374 B.n967 B.n94 10.6151
R2375 B.n967 B.n966 10.6151
R2376 B.n966 B.n965 10.6151
R2377 B.n965 B.n100 10.6151
R2378 B.n959 B.n100 10.6151
R2379 B.n959 B.n958 10.6151
R2380 B.n958 B.n957 10.6151
R2381 B.n957 B.n108 10.6151
R2382 B.n951 B.n108 10.6151
R2383 B.n951 B.n950 10.6151
R2384 B.n950 B.n949 10.6151
R2385 B.n949 B.n115 10.6151
R2386 B.n943 B.n115 10.6151
R2387 B.n943 B.n942 10.6151
R2388 B.n942 B.n941 10.6151
R2389 B.n941 B.n122 10.6151
R2390 B.n935 B.n122 10.6151
R2391 B.n935 B.n934 10.6151
R2392 B.n934 B.n933 10.6151
R2393 B.n933 B.n129 10.6151
R2394 B.n927 B.n129 10.6151
R2395 B.n927 B.n926 10.6151
R2396 B.n926 B.n925 10.6151
R2397 B.n925 B.n136 10.6151
R2398 B.n919 B.n136 10.6151
R2399 B.n157 B.n153 9.36635
R2400 B.n853 B.n852 9.36635
R2401 B.n425 B.n424 9.36635
R2402 B.n402 B.n348 9.36635
R2403 B.n310 B.t15 8.92344
R2404 B.t11 B.n938 8.92344
R2405 B.t8 B.n209 4.95769
R2406 B.t6 B.n36 4.95769
R2407 B.n1077 B.n0 2.81026
R2408 B.n1077 B.n1 2.81026
R2409 B.n871 B.n157 1.24928
R2410 B.n854 B.n853 1.24928
R2411 B.n424 B.n423 1.24928
R2412 B.n406 B.n348 1.24928
R2413 B.n545 B.t3 0.991938
R2414 B.n969 B.t7 0.991938
R2415 VN.n106 VN.n105 161.3
R2416 VN.n104 VN.n55 161.3
R2417 VN.n103 VN.n102 161.3
R2418 VN.n101 VN.n56 161.3
R2419 VN.n100 VN.n99 161.3
R2420 VN.n98 VN.n57 161.3
R2421 VN.n97 VN.n96 161.3
R2422 VN.n95 VN.n58 161.3
R2423 VN.n94 VN.n93 161.3
R2424 VN.n92 VN.n59 161.3
R2425 VN.n91 VN.n90 161.3
R2426 VN.n89 VN.n61 161.3
R2427 VN.n88 VN.n87 161.3
R2428 VN.n86 VN.n62 161.3
R2429 VN.n85 VN.n84 161.3
R2430 VN.n83 VN.n63 161.3
R2431 VN.n82 VN.n81 161.3
R2432 VN.n80 VN.n64 161.3
R2433 VN.n79 VN.n78 161.3
R2434 VN.n77 VN.n66 161.3
R2435 VN.n76 VN.n75 161.3
R2436 VN.n74 VN.n67 161.3
R2437 VN.n73 VN.n72 161.3
R2438 VN.n71 VN.n68 161.3
R2439 VN.n52 VN.n51 161.3
R2440 VN.n50 VN.n1 161.3
R2441 VN.n49 VN.n48 161.3
R2442 VN.n47 VN.n2 161.3
R2443 VN.n46 VN.n45 161.3
R2444 VN.n44 VN.n3 161.3
R2445 VN.n43 VN.n42 161.3
R2446 VN.n41 VN.n4 161.3
R2447 VN.n40 VN.n39 161.3
R2448 VN.n37 VN.n5 161.3
R2449 VN.n36 VN.n35 161.3
R2450 VN.n34 VN.n6 161.3
R2451 VN.n33 VN.n32 161.3
R2452 VN.n31 VN.n7 161.3
R2453 VN.n30 VN.n29 161.3
R2454 VN.n28 VN.n8 161.3
R2455 VN.n27 VN.n26 161.3
R2456 VN.n24 VN.n9 161.3
R2457 VN.n23 VN.n22 161.3
R2458 VN.n21 VN.n10 161.3
R2459 VN.n20 VN.n19 161.3
R2460 VN.n18 VN.n11 161.3
R2461 VN.n17 VN.n16 161.3
R2462 VN.n15 VN.n12 161.3
R2463 VN.n53 VN.n0 81.8843
R2464 VN.n107 VN.n54 81.8843
R2465 VN.n14 VN.t7 71.835
R2466 VN.n70 VN.t5 71.835
R2467 VN.n14 VN.n13 64.4539
R2468 VN.n70 VN.n69 64.4539
R2469 VN.n45 VN.n2 56.5617
R2470 VN.n99 VN.n56 56.5617
R2471 VN.n19 VN.n10 56.5617
R2472 VN.n32 VN.n6 56.5617
R2473 VN.n75 VN.n66 56.5617
R2474 VN.n87 VN.n61 56.5617
R2475 VN VN.n107 54.2936
R2476 VN.n13 VN.t6 38.6402
R2477 VN.n25 VN.t4 38.6402
R2478 VN.n38 VN.t0 38.6402
R2479 VN.n0 VN.t8 38.6402
R2480 VN.n69 VN.t9 38.6402
R2481 VN.n65 VN.t3 38.6402
R2482 VN.n60 VN.t2 38.6402
R2483 VN.n54 VN.t1 38.6402
R2484 VN.n17 VN.n12 24.5923
R2485 VN.n18 VN.n17 24.5923
R2486 VN.n19 VN.n18 24.5923
R2487 VN.n23 VN.n10 24.5923
R2488 VN.n24 VN.n23 24.5923
R2489 VN.n26 VN.n24 24.5923
R2490 VN.n30 VN.n8 24.5923
R2491 VN.n31 VN.n30 24.5923
R2492 VN.n32 VN.n31 24.5923
R2493 VN.n36 VN.n6 24.5923
R2494 VN.n37 VN.n36 24.5923
R2495 VN.n39 VN.n37 24.5923
R2496 VN.n43 VN.n4 24.5923
R2497 VN.n44 VN.n43 24.5923
R2498 VN.n45 VN.n44 24.5923
R2499 VN.n49 VN.n2 24.5923
R2500 VN.n50 VN.n49 24.5923
R2501 VN.n51 VN.n50 24.5923
R2502 VN.n75 VN.n74 24.5923
R2503 VN.n74 VN.n73 24.5923
R2504 VN.n73 VN.n68 24.5923
R2505 VN.n87 VN.n86 24.5923
R2506 VN.n86 VN.n85 24.5923
R2507 VN.n85 VN.n63 24.5923
R2508 VN.n81 VN.n80 24.5923
R2509 VN.n80 VN.n79 24.5923
R2510 VN.n79 VN.n66 24.5923
R2511 VN.n99 VN.n98 24.5923
R2512 VN.n98 VN.n97 24.5923
R2513 VN.n97 VN.n58 24.5923
R2514 VN.n93 VN.n92 24.5923
R2515 VN.n92 VN.n91 24.5923
R2516 VN.n91 VN.n61 24.5923
R2517 VN.n105 VN.n104 24.5923
R2518 VN.n104 VN.n103 24.5923
R2519 VN.n103 VN.n56 24.5923
R2520 VN.n38 VN.n4 14.2638
R2521 VN.n60 VN.n58 14.2638
R2522 VN.n26 VN.n25 12.2964
R2523 VN.n25 VN.n8 12.2964
R2524 VN.n65 VN.n63 12.2964
R2525 VN.n81 VN.n65 12.2964
R2526 VN.n13 VN.n12 10.3291
R2527 VN.n39 VN.n38 10.3291
R2528 VN.n69 VN.n68 10.3291
R2529 VN.n93 VN.n60 10.3291
R2530 VN.n51 VN.n0 8.36172
R2531 VN.n105 VN.n54 8.36172
R2532 VN.n15 VN.n14 3.19893
R2533 VN.n71 VN.n70 3.19893
R2534 VN.n107 VN.n106 0.354861
R2535 VN.n53 VN.n52 0.354861
R2536 VN VN.n53 0.267071
R2537 VN.n106 VN.n55 0.189894
R2538 VN.n102 VN.n55 0.189894
R2539 VN.n102 VN.n101 0.189894
R2540 VN.n101 VN.n100 0.189894
R2541 VN.n100 VN.n57 0.189894
R2542 VN.n96 VN.n57 0.189894
R2543 VN.n96 VN.n95 0.189894
R2544 VN.n95 VN.n94 0.189894
R2545 VN.n94 VN.n59 0.189894
R2546 VN.n90 VN.n59 0.189894
R2547 VN.n90 VN.n89 0.189894
R2548 VN.n89 VN.n88 0.189894
R2549 VN.n88 VN.n62 0.189894
R2550 VN.n84 VN.n62 0.189894
R2551 VN.n84 VN.n83 0.189894
R2552 VN.n83 VN.n82 0.189894
R2553 VN.n82 VN.n64 0.189894
R2554 VN.n78 VN.n64 0.189894
R2555 VN.n78 VN.n77 0.189894
R2556 VN.n77 VN.n76 0.189894
R2557 VN.n76 VN.n67 0.189894
R2558 VN.n72 VN.n67 0.189894
R2559 VN.n72 VN.n71 0.189894
R2560 VN.n16 VN.n15 0.189894
R2561 VN.n16 VN.n11 0.189894
R2562 VN.n20 VN.n11 0.189894
R2563 VN.n21 VN.n20 0.189894
R2564 VN.n22 VN.n21 0.189894
R2565 VN.n22 VN.n9 0.189894
R2566 VN.n27 VN.n9 0.189894
R2567 VN.n28 VN.n27 0.189894
R2568 VN.n29 VN.n28 0.189894
R2569 VN.n29 VN.n7 0.189894
R2570 VN.n33 VN.n7 0.189894
R2571 VN.n34 VN.n33 0.189894
R2572 VN.n35 VN.n34 0.189894
R2573 VN.n35 VN.n5 0.189894
R2574 VN.n40 VN.n5 0.189894
R2575 VN.n41 VN.n40 0.189894
R2576 VN.n42 VN.n41 0.189894
R2577 VN.n42 VN.n3 0.189894
R2578 VN.n46 VN.n3 0.189894
R2579 VN.n47 VN.n46 0.189894
R2580 VN.n48 VN.n47 0.189894
R2581 VN.n48 VN.n1 0.189894
R2582 VN.n52 VN.n1 0.189894
R2583 VDD2.n61 VDD2.n60 289.615
R2584 VDD2.n28 VDD2.n27 289.615
R2585 VDD2.n60 VDD2.n59 185
R2586 VDD2.n35 VDD2.n34 185
R2587 VDD2.n54 VDD2.n53 185
R2588 VDD2.n52 VDD2.n51 185
R2589 VDD2.n39 VDD2.n38 185
R2590 VDD2.n46 VDD2.n45 185
R2591 VDD2.n44 VDD2.n43 185
R2592 VDD2.n11 VDD2.n10 185
R2593 VDD2.n13 VDD2.n12 185
R2594 VDD2.n6 VDD2.n5 185
R2595 VDD2.n19 VDD2.n18 185
R2596 VDD2.n21 VDD2.n20 185
R2597 VDD2.n2 VDD2.n1 185
R2598 VDD2.n27 VDD2.n26 185
R2599 VDD2.n42 VDD2.t8 149.528
R2600 VDD2.n9 VDD2.t2 149.528
R2601 VDD2.n60 VDD2.n34 104.615
R2602 VDD2.n53 VDD2.n34 104.615
R2603 VDD2.n53 VDD2.n52 104.615
R2604 VDD2.n52 VDD2.n38 104.615
R2605 VDD2.n45 VDD2.n38 104.615
R2606 VDD2.n45 VDD2.n44 104.615
R2607 VDD2.n12 VDD2.n11 104.615
R2608 VDD2.n12 VDD2.n5 104.615
R2609 VDD2.n19 VDD2.n5 104.615
R2610 VDD2.n20 VDD2.n19 104.615
R2611 VDD2.n20 VDD2.n1 104.615
R2612 VDD2.n27 VDD2.n1 104.615
R2613 VDD2.n32 VDD2.n31 72.3701
R2614 VDD2 VDD2.n65 72.3671
R2615 VDD2.n64 VDD2.n63 69.8661
R2616 VDD2.n30 VDD2.n29 69.8651
R2617 VDD2.n30 VDD2.n28 54.6052
R2618 VDD2.n44 VDD2.t8 52.3082
R2619 VDD2.n11 VDD2.t2 52.3082
R2620 VDD2.n62 VDD2.n61 51.1914
R2621 VDD2.n62 VDD2.n32 44.9481
R2622 VDD2.n59 VDD2.n33 12.0247
R2623 VDD2.n26 VDD2.n0 12.0247
R2624 VDD2.n58 VDD2.n35 11.249
R2625 VDD2.n25 VDD2.n2 11.249
R2626 VDD2.n55 VDD2.n54 10.4732
R2627 VDD2.n22 VDD2.n21 10.4732
R2628 VDD2.n43 VDD2.n42 10.2745
R2629 VDD2.n10 VDD2.n9 10.2745
R2630 VDD2.n51 VDD2.n37 9.69747
R2631 VDD2.n18 VDD2.n4 9.69747
R2632 VDD2.n57 VDD2.n33 9.45567
R2633 VDD2.n24 VDD2.n0 9.45567
R2634 VDD2.n48 VDD2.n47 9.3005
R2635 VDD2.n50 VDD2.n49 9.3005
R2636 VDD2.n37 VDD2.n36 9.3005
R2637 VDD2.n56 VDD2.n55 9.3005
R2638 VDD2.n58 VDD2.n57 9.3005
R2639 VDD2.n41 VDD2.n40 9.3005
R2640 VDD2.n8 VDD2.n7 9.3005
R2641 VDD2.n15 VDD2.n14 9.3005
R2642 VDD2.n17 VDD2.n16 9.3005
R2643 VDD2.n4 VDD2.n3 9.3005
R2644 VDD2.n23 VDD2.n22 9.3005
R2645 VDD2.n25 VDD2.n24 9.3005
R2646 VDD2.n50 VDD2.n39 8.92171
R2647 VDD2.n17 VDD2.n6 8.92171
R2648 VDD2.n47 VDD2.n46 8.14595
R2649 VDD2.n14 VDD2.n13 8.14595
R2650 VDD2.n43 VDD2.n41 7.3702
R2651 VDD2.n10 VDD2.n8 7.3702
R2652 VDD2.n46 VDD2.n41 5.81868
R2653 VDD2.n13 VDD2.n8 5.81868
R2654 VDD2.n47 VDD2.n39 5.04292
R2655 VDD2.n14 VDD2.n6 5.04292
R2656 VDD2.n51 VDD2.n50 4.26717
R2657 VDD2.n18 VDD2.n17 4.26717
R2658 VDD2.n54 VDD2.n37 3.49141
R2659 VDD2.n21 VDD2.n4 3.49141
R2660 VDD2.n64 VDD2.n62 3.41429
R2661 VDD2.n65 VDD2.t0 3.40256
R2662 VDD2.n65 VDD2.t4 3.40256
R2663 VDD2.n63 VDD2.t7 3.40256
R2664 VDD2.n63 VDD2.t6 3.40256
R2665 VDD2.n31 VDD2.t9 3.40256
R2666 VDD2.n31 VDD2.t1 3.40256
R2667 VDD2.n29 VDD2.t3 3.40256
R2668 VDD2.n29 VDD2.t5 3.40256
R2669 VDD2.n42 VDD2.n40 2.84323
R2670 VDD2.n9 VDD2.n7 2.84323
R2671 VDD2.n55 VDD2.n35 2.71565
R2672 VDD2.n22 VDD2.n2 2.71565
R2673 VDD2.n59 VDD2.n58 1.93989
R2674 VDD2.n26 VDD2.n25 1.93989
R2675 VDD2.n61 VDD2.n33 1.16414
R2676 VDD2.n28 VDD2.n0 1.16414
R2677 VDD2 VDD2.n64 0.912138
R2678 VDD2.n32 VDD2.n30 0.798602
R2679 VDD2.n57 VDD2.n56 0.155672
R2680 VDD2.n56 VDD2.n36 0.155672
R2681 VDD2.n49 VDD2.n36 0.155672
R2682 VDD2.n49 VDD2.n48 0.155672
R2683 VDD2.n48 VDD2.n40 0.155672
R2684 VDD2.n15 VDD2.n7 0.155672
R2685 VDD2.n16 VDD2.n15 0.155672
R2686 VDD2.n16 VDD2.n3 0.155672
R2687 VDD2.n23 VDD2.n3 0.155672
R2688 VDD2.n24 VDD2.n23 0.155672
C0 VTAIL VDD1 8.44897f
C1 VP VN 8.76389f
C2 VP VDD2 0.715072f
C3 VN VDD2 5.75993f
C4 VP VTAIL 7.42699f
C5 VN VTAIL 7.41275f
C6 VP VDD1 6.31569f
C7 VTAIL VDD2 8.508691f
C8 VN VDD1 0.156225f
C9 VDD1 VDD2 2.84616f
C10 VDD2 B 7.38302f
C11 VDD1 B 7.308465f
C12 VTAIL B 5.896188f
C13 VN B 22.381142f
C14 VP B 20.921171f
C15 VDD2.n0 B 0.01516f
C16 VDD2.n1 B 0.03418f
C17 VDD2.n2 B 0.015311f
C18 VDD2.n3 B 0.026911f
C19 VDD2.n4 B 0.014461f
C20 VDD2.n5 B 0.03418f
C21 VDD2.n6 B 0.015311f
C22 VDD2.n7 B 0.617499f
C23 VDD2.n8 B 0.014461f
C24 VDD2.t2 B 0.056973f
C25 VDD2.n9 B 0.130427f
C26 VDD2.n10 B 0.024161f
C27 VDD2.n11 B 0.025635f
C28 VDD2.n12 B 0.03418f
C29 VDD2.n13 B 0.015311f
C30 VDD2.n14 B 0.014461f
C31 VDD2.n15 B 0.026911f
C32 VDD2.n16 B 0.026911f
C33 VDD2.n17 B 0.014461f
C34 VDD2.n18 B 0.015311f
C35 VDD2.n19 B 0.03418f
C36 VDD2.n20 B 0.03418f
C37 VDD2.n21 B 0.015311f
C38 VDD2.n22 B 0.014461f
C39 VDD2.n23 B 0.026911f
C40 VDD2.n24 B 0.068821f
C41 VDD2.n25 B 0.014461f
C42 VDD2.n26 B 0.015311f
C43 VDD2.n27 B 0.068215f
C44 VDD2.n28 B 0.098019f
C45 VDD2.t3 B 0.123767f
C46 VDD2.t5 B 0.123767f
C47 VDD2.n29 B 1.03988f
C48 VDD2.n30 B 0.900732f
C49 VDD2.t9 B 0.123767f
C50 VDD2.t1 B 0.123767f
C51 VDD2.n31 B 1.06517f
C52 VDD2.n32 B 3.2833f
C53 VDD2.n33 B 0.01516f
C54 VDD2.n34 B 0.03418f
C55 VDD2.n35 B 0.015311f
C56 VDD2.n36 B 0.026911f
C57 VDD2.n37 B 0.014461f
C58 VDD2.n38 B 0.03418f
C59 VDD2.n39 B 0.015311f
C60 VDD2.n40 B 0.617499f
C61 VDD2.n41 B 0.014461f
C62 VDD2.t8 B 0.056973f
C63 VDD2.n42 B 0.130427f
C64 VDD2.n43 B 0.024161f
C65 VDD2.n44 B 0.025635f
C66 VDD2.n45 B 0.03418f
C67 VDD2.n46 B 0.015311f
C68 VDD2.n47 B 0.014461f
C69 VDD2.n48 B 0.026911f
C70 VDD2.n49 B 0.026911f
C71 VDD2.n50 B 0.014461f
C72 VDD2.n51 B 0.015311f
C73 VDD2.n52 B 0.03418f
C74 VDD2.n53 B 0.03418f
C75 VDD2.n54 B 0.015311f
C76 VDD2.n55 B 0.014461f
C77 VDD2.n56 B 0.026911f
C78 VDD2.n57 B 0.068821f
C79 VDD2.n58 B 0.014461f
C80 VDD2.n59 B 0.015311f
C81 VDD2.n60 B 0.068215f
C82 VDD2.n61 B 0.076115f
C83 VDD2.n62 B 3.03131f
C84 VDD2.t7 B 0.123767f
C85 VDD2.t6 B 0.123767f
C86 VDD2.n63 B 1.03988f
C87 VDD2.n64 B 0.581335f
C88 VDD2.t0 B 0.123767f
C89 VDD2.t4 B 0.123767f
C90 VDD2.n65 B 1.06512f
C91 VN.t8 B 1.12557f
C92 VN.n0 B 0.494376f
C93 VN.n1 B 0.020166f
C94 VN.n2 B 0.032662f
C95 VN.n3 B 0.020166f
C96 VN.n4 B 0.029642f
C97 VN.n5 B 0.020166f
C98 VN.n6 B 0.03043f
C99 VN.n7 B 0.020166f
C100 VN.n8 B 0.028165f
C101 VN.n9 B 0.020166f
C102 VN.n10 B 0.028198f
C103 VN.n11 B 0.020166f
C104 VN.n12 B 0.026688f
C105 VN.t6 B 1.12557f
C106 VN.n13 B 0.484791f
C107 VN.t7 B 1.38858f
C108 VN.n14 B 0.466524f
C109 VN.n15 B 0.252734f
C110 VN.n16 B 0.020166f
C111 VN.n17 B 0.037396f
C112 VN.n18 B 0.037396f
C113 VN.n19 B 0.03043f
C114 VN.n20 B 0.020166f
C115 VN.n21 B 0.020166f
C116 VN.n22 B 0.020166f
C117 VN.n23 B 0.037396f
C118 VN.n24 B 0.037396f
C119 VN.t4 B 1.12557f
C120 VN.n25 B 0.416446f
C121 VN.n26 B 0.028165f
C122 VN.n27 B 0.020166f
C123 VN.n28 B 0.020166f
C124 VN.n29 B 0.020166f
C125 VN.n30 B 0.037396f
C126 VN.n31 B 0.037396f
C127 VN.n32 B 0.028198f
C128 VN.n33 B 0.020166f
C129 VN.n34 B 0.020166f
C130 VN.n35 B 0.020166f
C131 VN.n36 B 0.037396f
C132 VN.n37 B 0.037396f
C133 VN.t0 B 1.12557f
C134 VN.n38 B 0.416446f
C135 VN.n39 B 0.026688f
C136 VN.n40 B 0.020166f
C137 VN.n41 B 0.020166f
C138 VN.n42 B 0.020166f
C139 VN.n43 B 0.037396f
C140 VN.n44 B 0.037396f
C141 VN.n45 B 0.025967f
C142 VN.n46 B 0.020166f
C143 VN.n47 B 0.020166f
C144 VN.n48 B 0.020166f
C145 VN.n49 B 0.037396f
C146 VN.n50 B 0.037396f
C147 VN.n51 B 0.025211f
C148 VN.n52 B 0.032542f
C149 VN.n53 B 0.056555f
C150 VN.t1 B 1.12557f
C151 VN.n54 B 0.494376f
C152 VN.n55 B 0.020166f
C153 VN.n56 B 0.032662f
C154 VN.n57 B 0.020166f
C155 VN.n58 B 0.029642f
C156 VN.n59 B 0.020166f
C157 VN.t2 B 1.12557f
C158 VN.n60 B 0.416446f
C159 VN.n61 B 0.03043f
C160 VN.n62 B 0.020166f
C161 VN.n63 B 0.028165f
C162 VN.n64 B 0.020166f
C163 VN.t3 B 1.12557f
C164 VN.n65 B 0.416446f
C165 VN.n66 B 0.028198f
C166 VN.n67 B 0.020166f
C167 VN.n68 B 0.026688f
C168 VN.t5 B 1.38858f
C169 VN.t9 B 1.12557f
C170 VN.n69 B 0.484791f
C171 VN.n70 B 0.466524f
C172 VN.n71 B 0.252734f
C173 VN.n72 B 0.020166f
C174 VN.n73 B 0.037396f
C175 VN.n74 B 0.037396f
C176 VN.n75 B 0.03043f
C177 VN.n76 B 0.020166f
C178 VN.n77 B 0.020166f
C179 VN.n78 B 0.020166f
C180 VN.n79 B 0.037396f
C181 VN.n80 B 0.037396f
C182 VN.n81 B 0.028165f
C183 VN.n82 B 0.020166f
C184 VN.n83 B 0.020166f
C185 VN.n84 B 0.020166f
C186 VN.n85 B 0.037396f
C187 VN.n86 B 0.037396f
C188 VN.n87 B 0.028198f
C189 VN.n88 B 0.020166f
C190 VN.n89 B 0.020166f
C191 VN.n90 B 0.020166f
C192 VN.n91 B 0.037396f
C193 VN.n92 B 0.037396f
C194 VN.n93 B 0.026688f
C195 VN.n94 B 0.020166f
C196 VN.n95 B 0.020166f
C197 VN.n96 B 0.020166f
C198 VN.n97 B 0.037396f
C199 VN.n98 B 0.037396f
C200 VN.n99 B 0.025967f
C201 VN.n100 B 0.020166f
C202 VN.n101 B 0.020166f
C203 VN.n102 B 0.020166f
C204 VN.n103 B 0.037396f
C205 VN.n104 B 0.037396f
C206 VN.n105 B 0.025211f
C207 VN.n106 B 0.032542f
C208 VN.n107 B 1.29957f
C209 VTAIL.t5 B 0.138563f
C210 VTAIL.t6 B 0.138563f
C211 VTAIL.n0 B 1.09357f
C212 VTAIL.n1 B 0.726104f
C213 VTAIL.n2 B 0.016972f
C214 VTAIL.n3 B 0.038266f
C215 VTAIL.n4 B 0.017142f
C216 VTAIL.n5 B 0.030128f
C217 VTAIL.n6 B 0.01619f
C218 VTAIL.n7 B 0.038266f
C219 VTAIL.n8 B 0.017142f
C220 VTAIL.n9 B 0.691315f
C221 VTAIL.n10 B 0.01619f
C222 VTAIL.t13 B 0.063783f
C223 VTAIL.n11 B 0.146018f
C224 VTAIL.n12 B 0.02705f
C225 VTAIL.n13 B 0.028699f
C226 VTAIL.n14 B 0.038266f
C227 VTAIL.n15 B 0.017142f
C228 VTAIL.n16 B 0.01619f
C229 VTAIL.n17 B 0.030128f
C230 VTAIL.n18 B 0.030128f
C231 VTAIL.n19 B 0.01619f
C232 VTAIL.n20 B 0.017142f
C233 VTAIL.n21 B 0.038266f
C234 VTAIL.n22 B 0.038266f
C235 VTAIL.n23 B 0.017142f
C236 VTAIL.n24 B 0.01619f
C237 VTAIL.n25 B 0.030128f
C238 VTAIL.n26 B 0.077048f
C239 VTAIL.n27 B 0.01619f
C240 VTAIL.n28 B 0.017142f
C241 VTAIL.n29 B 0.076369f
C242 VTAIL.n30 B 0.064447f
C243 VTAIL.n31 B 0.571246f
C244 VTAIL.t16 B 0.138563f
C245 VTAIL.t14 B 0.138563f
C246 VTAIL.n32 B 1.09357f
C247 VTAIL.n33 B 0.9234f
C248 VTAIL.t12 B 0.138563f
C249 VTAIL.t11 B 0.138563f
C250 VTAIL.n34 B 1.09357f
C251 VTAIL.n35 B 2.15113f
C252 VTAIL.t3 B 0.138563f
C253 VTAIL.t2 B 0.138563f
C254 VTAIL.n36 B 1.09357f
C255 VTAIL.n37 B 2.15113f
C256 VTAIL.t0 B 0.138563f
C257 VTAIL.t8 B 0.138563f
C258 VTAIL.n38 B 1.09357f
C259 VTAIL.n39 B 0.923401f
C260 VTAIL.n40 B 0.016972f
C261 VTAIL.n41 B 0.038266f
C262 VTAIL.n42 B 0.017142f
C263 VTAIL.n43 B 0.030128f
C264 VTAIL.n44 B 0.01619f
C265 VTAIL.n45 B 0.038266f
C266 VTAIL.n46 B 0.017142f
C267 VTAIL.n47 B 0.691315f
C268 VTAIL.n48 B 0.01619f
C269 VTAIL.t4 B 0.063783f
C270 VTAIL.n49 B 0.146018f
C271 VTAIL.n50 B 0.02705f
C272 VTAIL.n51 B 0.028699f
C273 VTAIL.n52 B 0.038266f
C274 VTAIL.n53 B 0.017142f
C275 VTAIL.n54 B 0.01619f
C276 VTAIL.n55 B 0.030128f
C277 VTAIL.n56 B 0.030128f
C278 VTAIL.n57 B 0.01619f
C279 VTAIL.n58 B 0.017142f
C280 VTAIL.n59 B 0.038266f
C281 VTAIL.n60 B 0.038266f
C282 VTAIL.n61 B 0.017142f
C283 VTAIL.n62 B 0.01619f
C284 VTAIL.n63 B 0.030128f
C285 VTAIL.n64 B 0.077048f
C286 VTAIL.n65 B 0.01619f
C287 VTAIL.n66 B 0.017142f
C288 VTAIL.n67 B 0.076369f
C289 VTAIL.n68 B 0.064447f
C290 VTAIL.n69 B 0.571246f
C291 VTAIL.t9 B 0.138563f
C292 VTAIL.t15 B 0.138563f
C293 VTAIL.n70 B 1.09357f
C294 VTAIL.n71 B 0.803308f
C295 VTAIL.t17 B 0.138563f
C296 VTAIL.t18 B 0.138563f
C297 VTAIL.n72 B 1.09357f
C298 VTAIL.n73 B 0.923401f
C299 VTAIL.n74 B 0.016972f
C300 VTAIL.n75 B 0.038266f
C301 VTAIL.n76 B 0.017142f
C302 VTAIL.n77 B 0.030128f
C303 VTAIL.n78 B 0.01619f
C304 VTAIL.n79 B 0.038266f
C305 VTAIL.n80 B 0.017142f
C306 VTAIL.n81 B 0.691315f
C307 VTAIL.n82 B 0.01619f
C308 VTAIL.t10 B 0.063783f
C309 VTAIL.n83 B 0.146018f
C310 VTAIL.n84 B 0.02705f
C311 VTAIL.n85 B 0.028699f
C312 VTAIL.n86 B 0.038266f
C313 VTAIL.n87 B 0.017142f
C314 VTAIL.n88 B 0.01619f
C315 VTAIL.n89 B 0.030128f
C316 VTAIL.n90 B 0.030128f
C317 VTAIL.n91 B 0.01619f
C318 VTAIL.n92 B 0.017142f
C319 VTAIL.n93 B 0.038266f
C320 VTAIL.n94 B 0.038266f
C321 VTAIL.n95 B 0.017142f
C322 VTAIL.n96 B 0.01619f
C323 VTAIL.n97 B 0.030128f
C324 VTAIL.n98 B 0.077048f
C325 VTAIL.n99 B 0.01619f
C326 VTAIL.n100 B 0.017142f
C327 VTAIL.n101 B 0.076369f
C328 VTAIL.n102 B 0.064447f
C329 VTAIL.n103 B 1.58766f
C330 VTAIL.n104 B 0.016972f
C331 VTAIL.n105 B 0.038266f
C332 VTAIL.n106 B 0.017142f
C333 VTAIL.n107 B 0.030128f
C334 VTAIL.n108 B 0.01619f
C335 VTAIL.n109 B 0.038266f
C336 VTAIL.n110 B 0.017142f
C337 VTAIL.n111 B 0.691315f
C338 VTAIL.n112 B 0.01619f
C339 VTAIL.t7 B 0.063783f
C340 VTAIL.n113 B 0.146018f
C341 VTAIL.n114 B 0.02705f
C342 VTAIL.n115 B 0.028699f
C343 VTAIL.n116 B 0.038266f
C344 VTAIL.n117 B 0.017142f
C345 VTAIL.n118 B 0.01619f
C346 VTAIL.n119 B 0.030128f
C347 VTAIL.n120 B 0.030128f
C348 VTAIL.n121 B 0.01619f
C349 VTAIL.n122 B 0.017142f
C350 VTAIL.n123 B 0.038266f
C351 VTAIL.n124 B 0.038266f
C352 VTAIL.n125 B 0.017142f
C353 VTAIL.n126 B 0.01619f
C354 VTAIL.n127 B 0.030128f
C355 VTAIL.n128 B 0.077048f
C356 VTAIL.n129 B 0.01619f
C357 VTAIL.n130 B 0.017142f
C358 VTAIL.n131 B 0.076369f
C359 VTAIL.n132 B 0.064447f
C360 VTAIL.n133 B 1.58766f
C361 VTAIL.t1 B 0.138563f
C362 VTAIL.t19 B 0.138563f
C363 VTAIL.n134 B 1.09357f
C364 VTAIL.n135 B 0.669195f
C365 VDD1.n0 B 0.015425f
C366 VDD1.n1 B 0.034777f
C367 VDD1.n2 B 0.015579f
C368 VDD1.n3 B 0.027381f
C369 VDD1.n4 B 0.014713f
C370 VDD1.n5 B 0.034777f
C371 VDD1.n6 B 0.015579f
C372 VDD1.n7 B 0.628291f
C373 VDD1.n8 B 0.014713f
C374 VDD1.t0 B 0.057969f
C375 VDD1.n9 B 0.132706f
C376 VDD1.n10 B 0.024584f
C377 VDD1.n11 B 0.026083f
C378 VDD1.n12 B 0.034777f
C379 VDD1.n13 B 0.015579f
C380 VDD1.n14 B 0.014713f
C381 VDD1.n15 B 0.027381f
C382 VDD1.n16 B 0.027381f
C383 VDD1.n17 B 0.014713f
C384 VDD1.n18 B 0.015579f
C385 VDD1.n19 B 0.034777f
C386 VDD1.n20 B 0.034777f
C387 VDD1.n21 B 0.015579f
C388 VDD1.n22 B 0.014713f
C389 VDD1.n23 B 0.027381f
C390 VDD1.n24 B 0.070024f
C391 VDD1.n25 B 0.014713f
C392 VDD1.n26 B 0.015579f
C393 VDD1.n27 B 0.069407f
C394 VDD1.n28 B 0.099732f
C395 VDD1.t5 B 0.12593f
C396 VDD1.t7 B 0.12593f
C397 VDD1.n29 B 1.05805f
C398 VDD1.n30 B 0.925698f
C399 VDD1.n31 B 0.015425f
C400 VDD1.n32 B 0.034777f
C401 VDD1.n33 B 0.015579f
C402 VDD1.n34 B 0.027381f
C403 VDD1.n35 B 0.014713f
C404 VDD1.n36 B 0.034777f
C405 VDD1.n37 B 0.015579f
C406 VDD1.n38 B 0.628291f
C407 VDD1.n39 B 0.014713f
C408 VDD1.t6 B 0.057969f
C409 VDD1.n40 B 0.132706f
C410 VDD1.n41 B 0.024584f
C411 VDD1.n42 B 0.026083f
C412 VDD1.n43 B 0.034777f
C413 VDD1.n44 B 0.015579f
C414 VDD1.n45 B 0.014713f
C415 VDD1.n46 B 0.027381f
C416 VDD1.n47 B 0.027381f
C417 VDD1.n48 B 0.014713f
C418 VDD1.n49 B 0.015579f
C419 VDD1.n50 B 0.034777f
C420 VDD1.n51 B 0.034777f
C421 VDD1.n52 B 0.015579f
C422 VDD1.n53 B 0.014713f
C423 VDD1.n54 B 0.027381f
C424 VDD1.n55 B 0.070024f
C425 VDD1.n56 B 0.014713f
C426 VDD1.n57 B 0.015579f
C427 VDD1.n58 B 0.069407f
C428 VDD1.n59 B 0.099732f
C429 VDD1.t4 B 0.12593f
C430 VDD1.t3 B 0.12593f
C431 VDD1.n60 B 1.05805f
C432 VDD1.n61 B 0.916474f
C433 VDD1.t1 B 0.12593f
C434 VDD1.t2 B 0.12593f
C435 VDD1.n62 B 1.08378f
C436 VDD1.n63 B 3.50246f
C437 VDD1.t9 B 0.12593f
C438 VDD1.t8 B 0.12593f
C439 VDD1.n64 B 1.05805f
C440 VDD1.n65 B 3.41001f
C441 VP.t5 B 1.15264f
C442 VP.n0 B 0.506264f
C443 VP.n1 B 0.020651f
C444 VP.n2 B 0.033447f
C445 VP.n3 B 0.020651f
C446 VP.n4 B 0.030355f
C447 VP.n5 B 0.020651f
C448 VP.n6 B 0.031162f
C449 VP.n7 B 0.020651f
C450 VP.n8 B 0.028842f
C451 VP.n9 B 0.020651f
C452 VP.n10 B 0.028876f
C453 VP.n11 B 0.020651f
C454 VP.n12 B 0.02733f
C455 VP.n13 B 0.020651f
C456 VP.n14 B 0.026591f
C457 VP.n15 B 0.020651f
C458 VP.n16 B 0.025818f
C459 VP.t8 B 1.15264f
C460 VP.n17 B 0.506264f
C461 VP.n18 B 0.020651f
C462 VP.n19 B 0.033447f
C463 VP.n20 B 0.020651f
C464 VP.n21 B 0.030355f
C465 VP.n22 B 0.020651f
C466 VP.n23 B 0.031162f
C467 VP.n24 B 0.020651f
C468 VP.n25 B 0.028842f
C469 VP.n26 B 0.020651f
C470 VP.n27 B 0.028876f
C471 VP.n28 B 0.020651f
C472 VP.n29 B 0.02733f
C473 VP.t9 B 1.42197f
C474 VP.t3 B 1.15264f
C475 VP.n30 B 0.496448f
C476 VP.n31 B 0.477743f
C477 VP.n32 B 0.258811f
C478 VP.n33 B 0.020651f
C479 VP.n34 B 0.038295f
C480 VP.n35 B 0.038295f
C481 VP.n36 B 0.031162f
C482 VP.n37 B 0.020651f
C483 VP.n38 B 0.020651f
C484 VP.n39 B 0.020651f
C485 VP.n40 B 0.038295f
C486 VP.n41 B 0.038295f
C487 VP.t1 B 1.15264f
C488 VP.n42 B 0.42646f
C489 VP.n43 B 0.028842f
C490 VP.n44 B 0.020651f
C491 VP.n45 B 0.020651f
C492 VP.n46 B 0.020651f
C493 VP.n47 B 0.038295f
C494 VP.n48 B 0.038295f
C495 VP.n49 B 0.028876f
C496 VP.n50 B 0.020651f
C497 VP.n51 B 0.020651f
C498 VP.n52 B 0.020651f
C499 VP.n53 B 0.038295f
C500 VP.n54 B 0.038295f
C501 VP.t0 B 1.15264f
C502 VP.n55 B 0.42646f
C503 VP.n56 B 0.02733f
C504 VP.n57 B 0.020651f
C505 VP.n58 B 0.020651f
C506 VP.n59 B 0.020651f
C507 VP.n60 B 0.038295f
C508 VP.n61 B 0.038295f
C509 VP.n62 B 0.026591f
C510 VP.n63 B 0.020651f
C511 VP.n64 B 0.020651f
C512 VP.n65 B 0.020651f
C513 VP.n66 B 0.038295f
C514 VP.n67 B 0.038295f
C515 VP.n68 B 0.025818f
C516 VP.n69 B 0.033325f
C517 VP.n70 B 1.3226f
C518 VP.t6 B 1.15264f
C519 VP.n71 B 0.506264f
C520 VP.n72 B 1.33635f
C521 VP.n73 B 0.033325f
C522 VP.n74 B 0.020651f
C523 VP.n75 B 0.038295f
C524 VP.n76 B 0.038295f
C525 VP.n77 B 0.033447f
C526 VP.n78 B 0.020651f
C527 VP.n79 B 0.020651f
C528 VP.n80 B 0.020651f
C529 VP.n81 B 0.038295f
C530 VP.n82 B 0.038295f
C531 VP.t7 B 1.15264f
C532 VP.n83 B 0.42646f
C533 VP.n84 B 0.030355f
C534 VP.n85 B 0.020651f
C535 VP.n86 B 0.020651f
C536 VP.n87 B 0.020651f
C537 VP.n88 B 0.038295f
C538 VP.n89 B 0.038295f
C539 VP.n90 B 0.031162f
C540 VP.n91 B 0.020651f
C541 VP.n92 B 0.020651f
C542 VP.n93 B 0.020651f
C543 VP.n94 B 0.038295f
C544 VP.n95 B 0.038295f
C545 VP.t2 B 1.15264f
C546 VP.n96 B 0.42646f
C547 VP.n97 B 0.028842f
C548 VP.n98 B 0.020651f
C549 VP.n99 B 0.020651f
C550 VP.n100 B 0.020651f
C551 VP.n101 B 0.038295f
C552 VP.n102 B 0.038295f
C553 VP.n103 B 0.028876f
C554 VP.n104 B 0.020651f
C555 VP.n105 B 0.020651f
C556 VP.n106 B 0.020651f
C557 VP.n107 B 0.038295f
C558 VP.n108 B 0.038295f
C559 VP.t4 B 1.15264f
C560 VP.n109 B 0.42646f
C561 VP.n110 B 0.02733f
C562 VP.n111 B 0.020651f
C563 VP.n112 B 0.020651f
C564 VP.n113 B 0.020651f
C565 VP.n114 B 0.038295f
C566 VP.n115 B 0.038295f
C567 VP.n116 B 0.026591f
C568 VP.n117 B 0.020651f
C569 VP.n118 B 0.020651f
C570 VP.n119 B 0.020651f
C571 VP.n120 B 0.038295f
C572 VP.n121 B 0.038295f
C573 VP.n122 B 0.025818f
C574 VP.n123 B 0.033325f
C575 VP.n124 B 0.057915f
.ends

