* NGSPICE file created from diff_pair_sample_0416.ext - technology: sky130A

.subckt diff_pair_sample_0416 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3629 pd=8.59 as=3.2214 ps=17.3 w=8.26 l=2.06
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=0 ps=0 w=8.26 l=2.06
X2 VDD1.t2 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3629 pd=8.59 as=3.2214 ps=17.3 w=8.26 l=2.06
X3 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=1.3629 ps=8.59 w=8.26 l=2.06
X4 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=1.3629 ps=8.59 w=8.26 l=2.06
X5 VTAIL.t4 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=1.3629 ps=8.59 w=8.26 l=2.06
X6 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=0 ps=0 w=8.26 l=2.06
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=0 ps=0 w=8.26 l=2.06
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3629 pd=8.59 as=3.2214 ps=17.3 w=8.26 l=2.06
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=0 ps=0 w=8.26 l=2.06
X10 VTAIL.t7 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2214 pd=17.3 as=1.3629 ps=8.59 w=8.26 l=2.06
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3629 pd=8.59 as=3.2214 ps=17.3 w=8.26 l=2.06
R0 VP.n10 VP.n0 161.3
R1 VP.n9 VP.n8 161.3
R2 VP.n7 VP.n1 161.3
R3 VP.n6 VP.n5 161.3
R4 VP.n2 VP.t2 132.62
R5 VP.n2 VP.t0 132.078
R6 VP.n4 VP.t3 96.6345
R7 VP.n11 VP.t1 96.6345
R8 VP.n4 VP.n3 89.0215
R9 VP.n12 VP.n11 89.0215
R10 VP.n9 VP.n1 56.5617
R11 VP.n3 VP.n2 48.8659
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 21.8872
R15 VP.n11 VP.n10 21.8872
R16 VP.n6 VP.n3 0.278335
R17 VP.n12 VP.n0 0.278335
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153485
R22 VTAIL.n5 VTAIL.t4 51.3533
R23 VTAIL.n4 VTAIL.t2 51.3533
R24 VTAIL.n3 VTAIL.t3 51.3533
R25 VTAIL.n7 VTAIL.t0 51.3533
R26 VTAIL.n0 VTAIL.t1 51.3533
R27 VTAIL.n1 VTAIL.t6 51.3533
R28 VTAIL.n2 VTAIL.t7 51.3533
R29 VTAIL.n6 VTAIL.t5 51.3533
R30 VTAIL.n7 VTAIL.n6 21.5479
R31 VTAIL.n3 VTAIL.n2 21.5479
R32 VTAIL.n4 VTAIL.n3 2.06084
R33 VTAIL.n6 VTAIL.n5 2.06084
R34 VTAIL.n2 VTAIL.n1 2.06084
R35 VTAIL VTAIL.n0 1.08886
R36 VTAIL VTAIL.n7 0.972483
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 103.177
R40 VDD1 VDD1.n0 65.6931
R41 VDD1.n0 VDD1.t1 2.39759
R42 VDD1.n0 VDD1.t3 2.39759
R43 VDD1.n1 VDD1.t0 2.39759
R44 VDD1.n1 VDD1.t2 2.39759
R45 B.n601 B.n600 585
R46 B.n602 B.n601 585
R47 B.n236 B.n91 585
R48 B.n235 B.n234 585
R49 B.n233 B.n232 585
R50 B.n231 B.n230 585
R51 B.n229 B.n228 585
R52 B.n227 B.n226 585
R53 B.n225 B.n224 585
R54 B.n223 B.n222 585
R55 B.n221 B.n220 585
R56 B.n219 B.n218 585
R57 B.n217 B.n216 585
R58 B.n215 B.n214 585
R59 B.n213 B.n212 585
R60 B.n211 B.n210 585
R61 B.n209 B.n208 585
R62 B.n207 B.n206 585
R63 B.n205 B.n204 585
R64 B.n203 B.n202 585
R65 B.n201 B.n200 585
R66 B.n199 B.n198 585
R67 B.n197 B.n196 585
R68 B.n195 B.n194 585
R69 B.n193 B.n192 585
R70 B.n191 B.n190 585
R71 B.n189 B.n188 585
R72 B.n187 B.n186 585
R73 B.n185 B.n184 585
R74 B.n183 B.n182 585
R75 B.n181 B.n180 585
R76 B.n179 B.n178 585
R77 B.n177 B.n176 585
R78 B.n175 B.n174 585
R79 B.n173 B.n172 585
R80 B.n171 B.n170 585
R81 B.n169 B.n168 585
R82 B.n167 B.n166 585
R83 B.n165 B.n164 585
R84 B.n163 B.n162 585
R85 B.n161 B.n160 585
R86 B.n158 B.n157 585
R87 B.n156 B.n155 585
R88 B.n154 B.n153 585
R89 B.n152 B.n151 585
R90 B.n150 B.n149 585
R91 B.n148 B.n147 585
R92 B.n146 B.n145 585
R93 B.n144 B.n143 585
R94 B.n142 B.n141 585
R95 B.n140 B.n139 585
R96 B.n138 B.n137 585
R97 B.n136 B.n135 585
R98 B.n134 B.n133 585
R99 B.n132 B.n131 585
R100 B.n130 B.n129 585
R101 B.n128 B.n127 585
R102 B.n126 B.n125 585
R103 B.n124 B.n123 585
R104 B.n122 B.n121 585
R105 B.n120 B.n119 585
R106 B.n118 B.n117 585
R107 B.n116 B.n115 585
R108 B.n114 B.n113 585
R109 B.n112 B.n111 585
R110 B.n110 B.n109 585
R111 B.n108 B.n107 585
R112 B.n106 B.n105 585
R113 B.n104 B.n103 585
R114 B.n102 B.n101 585
R115 B.n100 B.n99 585
R116 B.n98 B.n97 585
R117 B.n599 B.n55 585
R118 B.n603 B.n55 585
R119 B.n598 B.n54 585
R120 B.n604 B.n54 585
R121 B.n597 B.n596 585
R122 B.n596 B.n50 585
R123 B.n595 B.n49 585
R124 B.n610 B.n49 585
R125 B.n594 B.n48 585
R126 B.n611 B.n48 585
R127 B.n593 B.n47 585
R128 B.n612 B.n47 585
R129 B.n592 B.n591 585
R130 B.n591 B.n46 585
R131 B.n590 B.n42 585
R132 B.n618 B.n42 585
R133 B.n589 B.n41 585
R134 B.n619 B.n41 585
R135 B.n588 B.n40 585
R136 B.n620 B.n40 585
R137 B.n587 B.n586 585
R138 B.n586 B.n36 585
R139 B.n585 B.n35 585
R140 B.n626 B.n35 585
R141 B.n584 B.n34 585
R142 B.n627 B.n34 585
R143 B.n583 B.n33 585
R144 B.n628 B.n33 585
R145 B.n582 B.n581 585
R146 B.n581 B.n29 585
R147 B.n580 B.n28 585
R148 B.n634 B.n28 585
R149 B.n579 B.n27 585
R150 B.n635 B.n27 585
R151 B.n578 B.n26 585
R152 B.n636 B.n26 585
R153 B.n577 B.n576 585
R154 B.n576 B.n22 585
R155 B.n575 B.n21 585
R156 B.n642 B.n21 585
R157 B.n574 B.n20 585
R158 B.n643 B.n20 585
R159 B.n573 B.n19 585
R160 B.n644 B.n19 585
R161 B.n572 B.n571 585
R162 B.n571 B.n15 585
R163 B.n570 B.n14 585
R164 B.n650 B.n14 585
R165 B.n569 B.n13 585
R166 B.n651 B.n13 585
R167 B.n568 B.n12 585
R168 B.n652 B.n12 585
R169 B.n567 B.n566 585
R170 B.n566 B.n8 585
R171 B.n565 B.n7 585
R172 B.n658 B.n7 585
R173 B.n564 B.n6 585
R174 B.n659 B.n6 585
R175 B.n563 B.n5 585
R176 B.n660 B.n5 585
R177 B.n562 B.n561 585
R178 B.n561 B.n4 585
R179 B.n560 B.n237 585
R180 B.n560 B.n559 585
R181 B.n550 B.n238 585
R182 B.n239 B.n238 585
R183 B.n552 B.n551 585
R184 B.n553 B.n552 585
R185 B.n549 B.n244 585
R186 B.n244 B.n243 585
R187 B.n548 B.n547 585
R188 B.n547 B.n546 585
R189 B.n246 B.n245 585
R190 B.n247 B.n246 585
R191 B.n539 B.n538 585
R192 B.n540 B.n539 585
R193 B.n537 B.n252 585
R194 B.n252 B.n251 585
R195 B.n536 B.n535 585
R196 B.n535 B.n534 585
R197 B.n254 B.n253 585
R198 B.n255 B.n254 585
R199 B.n527 B.n526 585
R200 B.n528 B.n527 585
R201 B.n525 B.n259 585
R202 B.n263 B.n259 585
R203 B.n524 B.n523 585
R204 B.n523 B.n522 585
R205 B.n261 B.n260 585
R206 B.n262 B.n261 585
R207 B.n515 B.n514 585
R208 B.n516 B.n515 585
R209 B.n513 B.n268 585
R210 B.n268 B.n267 585
R211 B.n512 B.n511 585
R212 B.n511 B.n510 585
R213 B.n270 B.n269 585
R214 B.n271 B.n270 585
R215 B.n503 B.n502 585
R216 B.n504 B.n503 585
R217 B.n501 B.n276 585
R218 B.n276 B.n275 585
R219 B.n500 B.n499 585
R220 B.n499 B.n498 585
R221 B.n278 B.n277 585
R222 B.n491 B.n278 585
R223 B.n490 B.n489 585
R224 B.n492 B.n490 585
R225 B.n488 B.n283 585
R226 B.n283 B.n282 585
R227 B.n487 B.n486 585
R228 B.n486 B.n485 585
R229 B.n285 B.n284 585
R230 B.n286 B.n285 585
R231 B.n478 B.n477 585
R232 B.n479 B.n478 585
R233 B.n476 B.n291 585
R234 B.n291 B.n290 585
R235 B.n470 B.n469 585
R236 B.n468 B.n328 585
R237 B.n467 B.n327 585
R238 B.n472 B.n327 585
R239 B.n466 B.n465 585
R240 B.n464 B.n463 585
R241 B.n462 B.n461 585
R242 B.n460 B.n459 585
R243 B.n458 B.n457 585
R244 B.n456 B.n455 585
R245 B.n454 B.n453 585
R246 B.n452 B.n451 585
R247 B.n450 B.n449 585
R248 B.n448 B.n447 585
R249 B.n446 B.n445 585
R250 B.n444 B.n443 585
R251 B.n442 B.n441 585
R252 B.n440 B.n439 585
R253 B.n438 B.n437 585
R254 B.n436 B.n435 585
R255 B.n434 B.n433 585
R256 B.n432 B.n431 585
R257 B.n430 B.n429 585
R258 B.n428 B.n427 585
R259 B.n426 B.n425 585
R260 B.n424 B.n423 585
R261 B.n422 B.n421 585
R262 B.n420 B.n419 585
R263 B.n418 B.n417 585
R264 B.n416 B.n415 585
R265 B.n414 B.n413 585
R266 B.n412 B.n411 585
R267 B.n410 B.n409 585
R268 B.n408 B.n407 585
R269 B.n406 B.n405 585
R270 B.n404 B.n403 585
R271 B.n402 B.n401 585
R272 B.n400 B.n399 585
R273 B.n398 B.n397 585
R274 B.n396 B.n395 585
R275 B.n394 B.n393 585
R276 B.n391 B.n390 585
R277 B.n389 B.n388 585
R278 B.n387 B.n386 585
R279 B.n385 B.n384 585
R280 B.n383 B.n382 585
R281 B.n381 B.n380 585
R282 B.n379 B.n378 585
R283 B.n377 B.n376 585
R284 B.n375 B.n374 585
R285 B.n373 B.n372 585
R286 B.n371 B.n370 585
R287 B.n369 B.n368 585
R288 B.n367 B.n366 585
R289 B.n365 B.n364 585
R290 B.n363 B.n362 585
R291 B.n361 B.n360 585
R292 B.n359 B.n358 585
R293 B.n357 B.n356 585
R294 B.n355 B.n354 585
R295 B.n353 B.n352 585
R296 B.n351 B.n350 585
R297 B.n349 B.n348 585
R298 B.n347 B.n346 585
R299 B.n345 B.n344 585
R300 B.n343 B.n342 585
R301 B.n341 B.n340 585
R302 B.n339 B.n338 585
R303 B.n337 B.n336 585
R304 B.n335 B.n334 585
R305 B.n293 B.n292 585
R306 B.n475 B.n474 585
R307 B.n289 B.n288 585
R308 B.n290 B.n289 585
R309 B.n481 B.n480 585
R310 B.n480 B.n479 585
R311 B.n482 B.n287 585
R312 B.n287 B.n286 585
R313 B.n484 B.n483 585
R314 B.n485 B.n484 585
R315 B.n281 B.n280 585
R316 B.n282 B.n281 585
R317 B.n494 B.n493 585
R318 B.n493 B.n492 585
R319 B.n495 B.n279 585
R320 B.n491 B.n279 585
R321 B.n497 B.n496 585
R322 B.n498 B.n497 585
R323 B.n274 B.n273 585
R324 B.n275 B.n274 585
R325 B.n506 B.n505 585
R326 B.n505 B.n504 585
R327 B.n507 B.n272 585
R328 B.n272 B.n271 585
R329 B.n509 B.n508 585
R330 B.n510 B.n509 585
R331 B.n266 B.n265 585
R332 B.n267 B.n266 585
R333 B.n518 B.n517 585
R334 B.n517 B.n516 585
R335 B.n519 B.n264 585
R336 B.n264 B.n262 585
R337 B.n521 B.n520 585
R338 B.n522 B.n521 585
R339 B.n258 B.n257 585
R340 B.n263 B.n258 585
R341 B.n530 B.n529 585
R342 B.n529 B.n528 585
R343 B.n531 B.n256 585
R344 B.n256 B.n255 585
R345 B.n533 B.n532 585
R346 B.n534 B.n533 585
R347 B.n250 B.n249 585
R348 B.n251 B.n250 585
R349 B.n542 B.n541 585
R350 B.n541 B.n540 585
R351 B.n543 B.n248 585
R352 B.n248 B.n247 585
R353 B.n545 B.n544 585
R354 B.n546 B.n545 585
R355 B.n242 B.n241 585
R356 B.n243 B.n242 585
R357 B.n555 B.n554 585
R358 B.n554 B.n553 585
R359 B.n556 B.n240 585
R360 B.n240 B.n239 585
R361 B.n558 B.n557 585
R362 B.n559 B.n558 585
R363 B.n2 B.n0 585
R364 B.n4 B.n2 585
R365 B.n3 B.n1 585
R366 B.n659 B.n3 585
R367 B.n657 B.n656 585
R368 B.n658 B.n657 585
R369 B.n655 B.n9 585
R370 B.n9 B.n8 585
R371 B.n654 B.n653 585
R372 B.n653 B.n652 585
R373 B.n11 B.n10 585
R374 B.n651 B.n11 585
R375 B.n649 B.n648 585
R376 B.n650 B.n649 585
R377 B.n647 B.n16 585
R378 B.n16 B.n15 585
R379 B.n646 B.n645 585
R380 B.n645 B.n644 585
R381 B.n18 B.n17 585
R382 B.n643 B.n18 585
R383 B.n641 B.n640 585
R384 B.n642 B.n641 585
R385 B.n639 B.n23 585
R386 B.n23 B.n22 585
R387 B.n638 B.n637 585
R388 B.n637 B.n636 585
R389 B.n25 B.n24 585
R390 B.n635 B.n25 585
R391 B.n633 B.n632 585
R392 B.n634 B.n633 585
R393 B.n631 B.n30 585
R394 B.n30 B.n29 585
R395 B.n630 B.n629 585
R396 B.n629 B.n628 585
R397 B.n32 B.n31 585
R398 B.n627 B.n32 585
R399 B.n625 B.n624 585
R400 B.n626 B.n625 585
R401 B.n623 B.n37 585
R402 B.n37 B.n36 585
R403 B.n622 B.n621 585
R404 B.n621 B.n620 585
R405 B.n39 B.n38 585
R406 B.n619 B.n39 585
R407 B.n617 B.n616 585
R408 B.n618 B.n617 585
R409 B.n615 B.n43 585
R410 B.n46 B.n43 585
R411 B.n614 B.n613 585
R412 B.n613 B.n612 585
R413 B.n45 B.n44 585
R414 B.n611 B.n45 585
R415 B.n609 B.n608 585
R416 B.n610 B.n609 585
R417 B.n607 B.n51 585
R418 B.n51 B.n50 585
R419 B.n606 B.n605 585
R420 B.n605 B.n604 585
R421 B.n53 B.n52 585
R422 B.n603 B.n53 585
R423 B.n662 B.n661 585
R424 B.n661 B.n660 585
R425 B.n470 B.n289 516.524
R426 B.n97 B.n53 516.524
R427 B.n474 B.n291 516.524
R428 B.n601 B.n55 516.524
R429 B.n332 B.t12 303.69
R430 B.n329 B.t8 303.69
R431 B.n95 B.t15 303.69
R432 B.n92 B.t4 303.69
R433 B.n602 B.n90 256.663
R434 B.n602 B.n89 256.663
R435 B.n602 B.n88 256.663
R436 B.n602 B.n87 256.663
R437 B.n602 B.n86 256.663
R438 B.n602 B.n85 256.663
R439 B.n602 B.n84 256.663
R440 B.n602 B.n83 256.663
R441 B.n602 B.n82 256.663
R442 B.n602 B.n81 256.663
R443 B.n602 B.n80 256.663
R444 B.n602 B.n79 256.663
R445 B.n602 B.n78 256.663
R446 B.n602 B.n77 256.663
R447 B.n602 B.n76 256.663
R448 B.n602 B.n75 256.663
R449 B.n602 B.n74 256.663
R450 B.n602 B.n73 256.663
R451 B.n602 B.n72 256.663
R452 B.n602 B.n71 256.663
R453 B.n602 B.n70 256.663
R454 B.n602 B.n69 256.663
R455 B.n602 B.n68 256.663
R456 B.n602 B.n67 256.663
R457 B.n602 B.n66 256.663
R458 B.n602 B.n65 256.663
R459 B.n602 B.n64 256.663
R460 B.n602 B.n63 256.663
R461 B.n602 B.n62 256.663
R462 B.n602 B.n61 256.663
R463 B.n602 B.n60 256.663
R464 B.n602 B.n59 256.663
R465 B.n602 B.n58 256.663
R466 B.n602 B.n57 256.663
R467 B.n602 B.n56 256.663
R468 B.n472 B.n471 256.663
R469 B.n472 B.n294 256.663
R470 B.n472 B.n295 256.663
R471 B.n472 B.n296 256.663
R472 B.n472 B.n297 256.663
R473 B.n472 B.n298 256.663
R474 B.n472 B.n299 256.663
R475 B.n472 B.n300 256.663
R476 B.n472 B.n301 256.663
R477 B.n472 B.n302 256.663
R478 B.n472 B.n303 256.663
R479 B.n472 B.n304 256.663
R480 B.n472 B.n305 256.663
R481 B.n472 B.n306 256.663
R482 B.n472 B.n307 256.663
R483 B.n472 B.n308 256.663
R484 B.n472 B.n309 256.663
R485 B.n472 B.n310 256.663
R486 B.n472 B.n311 256.663
R487 B.n472 B.n312 256.663
R488 B.n472 B.n313 256.663
R489 B.n472 B.n314 256.663
R490 B.n472 B.n315 256.663
R491 B.n472 B.n316 256.663
R492 B.n472 B.n317 256.663
R493 B.n472 B.n318 256.663
R494 B.n472 B.n319 256.663
R495 B.n472 B.n320 256.663
R496 B.n472 B.n321 256.663
R497 B.n472 B.n322 256.663
R498 B.n472 B.n323 256.663
R499 B.n472 B.n324 256.663
R500 B.n472 B.n325 256.663
R501 B.n472 B.n326 256.663
R502 B.n473 B.n472 256.663
R503 B.n480 B.n289 163.367
R504 B.n480 B.n287 163.367
R505 B.n484 B.n287 163.367
R506 B.n484 B.n281 163.367
R507 B.n493 B.n281 163.367
R508 B.n493 B.n279 163.367
R509 B.n497 B.n279 163.367
R510 B.n497 B.n274 163.367
R511 B.n505 B.n274 163.367
R512 B.n505 B.n272 163.367
R513 B.n509 B.n272 163.367
R514 B.n509 B.n266 163.367
R515 B.n517 B.n266 163.367
R516 B.n517 B.n264 163.367
R517 B.n521 B.n264 163.367
R518 B.n521 B.n258 163.367
R519 B.n529 B.n258 163.367
R520 B.n529 B.n256 163.367
R521 B.n533 B.n256 163.367
R522 B.n533 B.n250 163.367
R523 B.n541 B.n250 163.367
R524 B.n541 B.n248 163.367
R525 B.n545 B.n248 163.367
R526 B.n545 B.n242 163.367
R527 B.n554 B.n242 163.367
R528 B.n554 B.n240 163.367
R529 B.n558 B.n240 163.367
R530 B.n558 B.n2 163.367
R531 B.n661 B.n2 163.367
R532 B.n661 B.n3 163.367
R533 B.n657 B.n3 163.367
R534 B.n657 B.n9 163.367
R535 B.n653 B.n9 163.367
R536 B.n653 B.n11 163.367
R537 B.n649 B.n11 163.367
R538 B.n649 B.n16 163.367
R539 B.n645 B.n16 163.367
R540 B.n645 B.n18 163.367
R541 B.n641 B.n18 163.367
R542 B.n641 B.n23 163.367
R543 B.n637 B.n23 163.367
R544 B.n637 B.n25 163.367
R545 B.n633 B.n25 163.367
R546 B.n633 B.n30 163.367
R547 B.n629 B.n30 163.367
R548 B.n629 B.n32 163.367
R549 B.n625 B.n32 163.367
R550 B.n625 B.n37 163.367
R551 B.n621 B.n37 163.367
R552 B.n621 B.n39 163.367
R553 B.n617 B.n39 163.367
R554 B.n617 B.n43 163.367
R555 B.n613 B.n43 163.367
R556 B.n613 B.n45 163.367
R557 B.n609 B.n45 163.367
R558 B.n609 B.n51 163.367
R559 B.n605 B.n51 163.367
R560 B.n605 B.n53 163.367
R561 B.n328 B.n327 163.367
R562 B.n465 B.n327 163.367
R563 B.n463 B.n462 163.367
R564 B.n459 B.n458 163.367
R565 B.n455 B.n454 163.367
R566 B.n451 B.n450 163.367
R567 B.n447 B.n446 163.367
R568 B.n443 B.n442 163.367
R569 B.n439 B.n438 163.367
R570 B.n435 B.n434 163.367
R571 B.n431 B.n430 163.367
R572 B.n427 B.n426 163.367
R573 B.n423 B.n422 163.367
R574 B.n419 B.n418 163.367
R575 B.n415 B.n414 163.367
R576 B.n411 B.n410 163.367
R577 B.n407 B.n406 163.367
R578 B.n403 B.n402 163.367
R579 B.n399 B.n398 163.367
R580 B.n395 B.n394 163.367
R581 B.n390 B.n389 163.367
R582 B.n386 B.n385 163.367
R583 B.n382 B.n381 163.367
R584 B.n378 B.n377 163.367
R585 B.n374 B.n373 163.367
R586 B.n370 B.n369 163.367
R587 B.n366 B.n365 163.367
R588 B.n362 B.n361 163.367
R589 B.n358 B.n357 163.367
R590 B.n354 B.n353 163.367
R591 B.n350 B.n349 163.367
R592 B.n346 B.n345 163.367
R593 B.n342 B.n341 163.367
R594 B.n338 B.n337 163.367
R595 B.n334 B.n293 163.367
R596 B.n478 B.n291 163.367
R597 B.n478 B.n285 163.367
R598 B.n486 B.n285 163.367
R599 B.n486 B.n283 163.367
R600 B.n490 B.n283 163.367
R601 B.n490 B.n278 163.367
R602 B.n499 B.n278 163.367
R603 B.n499 B.n276 163.367
R604 B.n503 B.n276 163.367
R605 B.n503 B.n270 163.367
R606 B.n511 B.n270 163.367
R607 B.n511 B.n268 163.367
R608 B.n515 B.n268 163.367
R609 B.n515 B.n261 163.367
R610 B.n523 B.n261 163.367
R611 B.n523 B.n259 163.367
R612 B.n527 B.n259 163.367
R613 B.n527 B.n254 163.367
R614 B.n535 B.n254 163.367
R615 B.n535 B.n252 163.367
R616 B.n539 B.n252 163.367
R617 B.n539 B.n246 163.367
R618 B.n547 B.n246 163.367
R619 B.n547 B.n244 163.367
R620 B.n552 B.n244 163.367
R621 B.n552 B.n238 163.367
R622 B.n560 B.n238 163.367
R623 B.n561 B.n560 163.367
R624 B.n561 B.n5 163.367
R625 B.n6 B.n5 163.367
R626 B.n7 B.n6 163.367
R627 B.n566 B.n7 163.367
R628 B.n566 B.n12 163.367
R629 B.n13 B.n12 163.367
R630 B.n14 B.n13 163.367
R631 B.n571 B.n14 163.367
R632 B.n571 B.n19 163.367
R633 B.n20 B.n19 163.367
R634 B.n21 B.n20 163.367
R635 B.n576 B.n21 163.367
R636 B.n576 B.n26 163.367
R637 B.n27 B.n26 163.367
R638 B.n28 B.n27 163.367
R639 B.n581 B.n28 163.367
R640 B.n581 B.n33 163.367
R641 B.n34 B.n33 163.367
R642 B.n35 B.n34 163.367
R643 B.n586 B.n35 163.367
R644 B.n586 B.n40 163.367
R645 B.n41 B.n40 163.367
R646 B.n42 B.n41 163.367
R647 B.n591 B.n42 163.367
R648 B.n591 B.n47 163.367
R649 B.n48 B.n47 163.367
R650 B.n49 B.n48 163.367
R651 B.n596 B.n49 163.367
R652 B.n596 B.n54 163.367
R653 B.n55 B.n54 163.367
R654 B.n101 B.n100 163.367
R655 B.n105 B.n104 163.367
R656 B.n109 B.n108 163.367
R657 B.n113 B.n112 163.367
R658 B.n117 B.n116 163.367
R659 B.n121 B.n120 163.367
R660 B.n125 B.n124 163.367
R661 B.n129 B.n128 163.367
R662 B.n133 B.n132 163.367
R663 B.n137 B.n136 163.367
R664 B.n141 B.n140 163.367
R665 B.n145 B.n144 163.367
R666 B.n149 B.n148 163.367
R667 B.n153 B.n152 163.367
R668 B.n157 B.n156 163.367
R669 B.n162 B.n161 163.367
R670 B.n166 B.n165 163.367
R671 B.n170 B.n169 163.367
R672 B.n174 B.n173 163.367
R673 B.n178 B.n177 163.367
R674 B.n182 B.n181 163.367
R675 B.n186 B.n185 163.367
R676 B.n190 B.n189 163.367
R677 B.n194 B.n193 163.367
R678 B.n198 B.n197 163.367
R679 B.n202 B.n201 163.367
R680 B.n206 B.n205 163.367
R681 B.n210 B.n209 163.367
R682 B.n214 B.n213 163.367
R683 B.n218 B.n217 163.367
R684 B.n222 B.n221 163.367
R685 B.n226 B.n225 163.367
R686 B.n230 B.n229 163.367
R687 B.n234 B.n233 163.367
R688 B.n601 B.n91 163.367
R689 B.n332 B.t14 116.823
R690 B.n92 B.t6 116.823
R691 B.n329 B.t11 116.814
R692 B.n95 B.t16 116.814
R693 B.n472 B.n290 111.341
R694 B.n603 B.n602 111.341
R695 B.n471 B.n470 71.676
R696 B.n465 B.n294 71.676
R697 B.n462 B.n295 71.676
R698 B.n458 B.n296 71.676
R699 B.n454 B.n297 71.676
R700 B.n450 B.n298 71.676
R701 B.n446 B.n299 71.676
R702 B.n442 B.n300 71.676
R703 B.n438 B.n301 71.676
R704 B.n434 B.n302 71.676
R705 B.n430 B.n303 71.676
R706 B.n426 B.n304 71.676
R707 B.n422 B.n305 71.676
R708 B.n418 B.n306 71.676
R709 B.n414 B.n307 71.676
R710 B.n410 B.n308 71.676
R711 B.n406 B.n309 71.676
R712 B.n402 B.n310 71.676
R713 B.n398 B.n311 71.676
R714 B.n394 B.n312 71.676
R715 B.n389 B.n313 71.676
R716 B.n385 B.n314 71.676
R717 B.n381 B.n315 71.676
R718 B.n377 B.n316 71.676
R719 B.n373 B.n317 71.676
R720 B.n369 B.n318 71.676
R721 B.n365 B.n319 71.676
R722 B.n361 B.n320 71.676
R723 B.n357 B.n321 71.676
R724 B.n353 B.n322 71.676
R725 B.n349 B.n323 71.676
R726 B.n345 B.n324 71.676
R727 B.n341 B.n325 71.676
R728 B.n337 B.n326 71.676
R729 B.n473 B.n293 71.676
R730 B.n97 B.n56 71.676
R731 B.n101 B.n57 71.676
R732 B.n105 B.n58 71.676
R733 B.n109 B.n59 71.676
R734 B.n113 B.n60 71.676
R735 B.n117 B.n61 71.676
R736 B.n121 B.n62 71.676
R737 B.n125 B.n63 71.676
R738 B.n129 B.n64 71.676
R739 B.n133 B.n65 71.676
R740 B.n137 B.n66 71.676
R741 B.n141 B.n67 71.676
R742 B.n145 B.n68 71.676
R743 B.n149 B.n69 71.676
R744 B.n153 B.n70 71.676
R745 B.n157 B.n71 71.676
R746 B.n162 B.n72 71.676
R747 B.n166 B.n73 71.676
R748 B.n170 B.n74 71.676
R749 B.n174 B.n75 71.676
R750 B.n178 B.n76 71.676
R751 B.n182 B.n77 71.676
R752 B.n186 B.n78 71.676
R753 B.n190 B.n79 71.676
R754 B.n194 B.n80 71.676
R755 B.n198 B.n81 71.676
R756 B.n202 B.n82 71.676
R757 B.n206 B.n83 71.676
R758 B.n210 B.n84 71.676
R759 B.n214 B.n85 71.676
R760 B.n218 B.n86 71.676
R761 B.n222 B.n87 71.676
R762 B.n226 B.n88 71.676
R763 B.n230 B.n89 71.676
R764 B.n234 B.n90 71.676
R765 B.n91 B.n90 71.676
R766 B.n233 B.n89 71.676
R767 B.n229 B.n88 71.676
R768 B.n225 B.n87 71.676
R769 B.n221 B.n86 71.676
R770 B.n217 B.n85 71.676
R771 B.n213 B.n84 71.676
R772 B.n209 B.n83 71.676
R773 B.n205 B.n82 71.676
R774 B.n201 B.n81 71.676
R775 B.n197 B.n80 71.676
R776 B.n193 B.n79 71.676
R777 B.n189 B.n78 71.676
R778 B.n185 B.n77 71.676
R779 B.n181 B.n76 71.676
R780 B.n177 B.n75 71.676
R781 B.n173 B.n74 71.676
R782 B.n169 B.n73 71.676
R783 B.n165 B.n72 71.676
R784 B.n161 B.n71 71.676
R785 B.n156 B.n70 71.676
R786 B.n152 B.n69 71.676
R787 B.n148 B.n68 71.676
R788 B.n144 B.n67 71.676
R789 B.n140 B.n66 71.676
R790 B.n136 B.n65 71.676
R791 B.n132 B.n64 71.676
R792 B.n128 B.n63 71.676
R793 B.n124 B.n62 71.676
R794 B.n120 B.n61 71.676
R795 B.n116 B.n60 71.676
R796 B.n112 B.n59 71.676
R797 B.n108 B.n58 71.676
R798 B.n104 B.n57 71.676
R799 B.n100 B.n56 71.676
R800 B.n471 B.n328 71.676
R801 B.n463 B.n294 71.676
R802 B.n459 B.n295 71.676
R803 B.n455 B.n296 71.676
R804 B.n451 B.n297 71.676
R805 B.n447 B.n298 71.676
R806 B.n443 B.n299 71.676
R807 B.n439 B.n300 71.676
R808 B.n435 B.n301 71.676
R809 B.n431 B.n302 71.676
R810 B.n427 B.n303 71.676
R811 B.n423 B.n304 71.676
R812 B.n419 B.n305 71.676
R813 B.n415 B.n306 71.676
R814 B.n411 B.n307 71.676
R815 B.n407 B.n308 71.676
R816 B.n403 B.n309 71.676
R817 B.n399 B.n310 71.676
R818 B.n395 B.n311 71.676
R819 B.n390 B.n312 71.676
R820 B.n386 B.n313 71.676
R821 B.n382 B.n314 71.676
R822 B.n378 B.n315 71.676
R823 B.n374 B.n316 71.676
R824 B.n370 B.n317 71.676
R825 B.n366 B.n318 71.676
R826 B.n362 B.n319 71.676
R827 B.n358 B.n320 71.676
R828 B.n354 B.n321 71.676
R829 B.n350 B.n322 71.676
R830 B.n346 B.n323 71.676
R831 B.n342 B.n324 71.676
R832 B.n338 B.n325 71.676
R833 B.n334 B.n326 71.676
R834 B.n474 B.n473 71.676
R835 B.n333 B.t13 70.4714
R836 B.n93 B.t7 70.4714
R837 B.n330 B.t10 70.4616
R838 B.n96 B.t17 70.4616
R839 B.n392 B.n333 59.5399
R840 B.n331 B.n330 59.5399
R841 B.n159 B.n96 59.5399
R842 B.n94 B.n93 59.5399
R843 B.n479 B.n290 55.2646
R844 B.n479 B.n286 55.2646
R845 B.n485 B.n286 55.2646
R846 B.n485 B.n282 55.2646
R847 B.n492 B.n282 55.2646
R848 B.n492 B.n491 55.2646
R849 B.n498 B.n275 55.2646
R850 B.n504 B.n275 55.2646
R851 B.n504 B.n271 55.2646
R852 B.n510 B.n271 55.2646
R853 B.n510 B.n267 55.2646
R854 B.n516 B.n267 55.2646
R855 B.n516 B.n262 55.2646
R856 B.n522 B.n262 55.2646
R857 B.n522 B.n263 55.2646
R858 B.n528 B.n255 55.2646
R859 B.n534 B.n255 55.2646
R860 B.n534 B.n251 55.2646
R861 B.n540 B.n251 55.2646
R862 B.n540 B.n247 55.2646
R863 B.n546 B.n247 55.2646
R864 B.n553 B.n243 55.2646
R865 B.n553 B.n239 55.2646
R866 B.n559 B.n239 55.2646
R867 B.n559 B.n4 55.2646
R868 B.n660 B.n4 55.2646
R869 B.n660 B.n659 55.2646
R870 B.n659 B.n658 55.2646
R871 B.n658 B.n8 55.2646
R872 B.n652 B.n8 55.2646
R873 B.n652 B.n651 55.2646
R874 B.n650 B.n15 55.2646
R875 B.n644 B.n15 55.2646
R876 B.n644 B.n643 55.2646
R877 B.n643 B.n642 55.2646
R878 B.n642 B.n22 55.2646
R879 B.n636 B.n22 55.2646
R880 B.n635 B.n634 55.2646
R881 B.n634 B.n29 55.2646
R882 B.n628 B.n29 55.2646
R883 B.n628 B.n627 55.2646
R884 B.n627 B.n626 55.2646
R885 B.n626 B.n36 55.2646
R886 B.n620 B.n36 55.2646
R887 B.n620 B.n619 55.2646
R888 B.n619 B.n618 55.2646
R889 B.n612 B.n46 55.2646
R890 B.n612 B.n611 55.2646
R891 B.n611 B.n610 55.2646
R892 B.n610 B.n50 55.2646
R893 B.n604 B.n50 55.2646
R894 B.n604 B.n603 55.2646
R895 B.n546 B.t2 48.763
R896 B.t1 B.n650 48.763
R897 B.n263 B.t3 47.1376
R898 B.t0 B.n635 47.1376
R899 B.n333 B.n332 46.352
R900 B.n330 B.n329 46.352
R901 B.n96 B.n95 46.352
R902 B.n93 B.n92 46.352
R903 B.n491 B.t9 34.1342
R904 B.n46 B.t5 34.1342
R905 B.n98 B.n52 33.5615
R906 B.n600 B.n599 33.5615
R907 B.n476 B.n475 33.5615
R908 B.n469 B.n288 33.5615
R909 B.n498 B.t9 21.1309
R910 B.n618 B.t5 21.1309
R911 B B.n662 18.0485
R912 B.n99 B.n98 10.6151
R913 B.n102 B.n99 10.6151
R914 B.n103 B.n102 10.6151
R915 B.n106 B.n103 10.6151
R916 B.n107 B.n106 10.6151
R917 B.n110 B.n107 10.6151
R918 B.n111 B.n110 10.6151
R919 B.n114 B.n111 10.6151
R920 B.n115 B.n114 10.6151
R921 B.n118 B.n115 10.6151
R922 B.n119 B.n118 10.6151
R923 B.n122 B.n119 10.6151
R924 B.n123 B.n122 10.6151
R925 B.n126 B.n123 10.6151
R926 B.n127 B.n126 10.6151
R927 B.n130 B.n127 10.6151
R928 B.n131 B.n130 10.6151
R929 B.n134 B.n131 10.6151
R930 B.n135 B.n134 10.6151
R931 B.n138 B.n135 10.6151
R932 B.n139 B.n138 10.6151
R933 B.n142 B.n139 10.6151
R934 B.n143 B.n142 10.6151
R935 B.n146 B.n143 10.6151
R936 B.n147 B.n146 10.6151
R937 B.n150 B.n147 10.6151
R938 B.n151 B.n150 10.6151
R939 B.n154 B.n151 10.6151
R940 B.n155 B.n154 10.6151
R941 B.n158 B.n155 10.6151
R942 B.n163 B.n160 10.6151
R943 B.n164 B.n163 10.6151
R944 B.n167 B.n164 10.6151
R945 B.n168 B.n167 10.6151
R946 B.n171 B.n168 10.6151
R947 B.n172 B.n171 10.6151
R948 B.n175 B.n172 10.6151
R949 B.n176 B.n175 10.6151
R950 B.n180 B.n179 10.6151
R951 B.n183 B.n180 10.6151
R952 B.n184 B.n183 10.6151
R953 B.n187 B.n184 10.6151
R954 B.n188 B.n187 10.6151
R955 B.n191 B.n188 10.6151
R956 B.n192 B.n191 10.6151
R957 B.n195 B.n192 10.6151
R958 B.n196 B.n195 10.6151
R959 B.n199 B.n196 10.6151
R960 B.n200 B.n199 10.6151
R961 B.n203 B.n200 10.6151
R962 B.n204 B.n203 10.6151
R963 B.n207 B.n204 10.6151
R964 B.n208 B.n207 10.6151
R965 B.n211 B.n208 10.6151
R966 B.n212 B.n211 10.6151
R967 B.n215 B.n212 10.6151
R968 B.n216 B.n215 10.6151
R969 B.n219 B.n216 10.6151
R970 B.n220 B.n219 10.6151
R971 B.n223 B.n220 10.6151
R972 B.n224 B.n223 10.6151
R973 B.n227 B.n224 10.6151
R974 B.n228 B.n227 10.6151
R975 B.n231 B.n228 10.6151
R976 B.n232 B.n231 10.6151
R977 B.n235 B.n232 10.6151
R978 B.n236 B.n235 10.6151
R979 B.n600 B.n236 10.6151
R980 B.n477 B.n476 10.6151
R981 B.n477 B.n284 10.6151
R982 B.n487 B.n284 10.6151
R983 B.n488 B.n487 10.6151
R984 B.n489 B.n488 10.6151
R985 B.n489 B.n277 10.6151
R986 B.n500 B.n277 10.6151
R987 B.n501 B.n500 10.6151
R988 B.n502 B.n501 10.6151
R989 B.n502 B.n269 10.6151
R990 B.n512 B.n269 10.6151
R991 B.n513 B.n512 10.6151
R992 B.n514 B.n513 10.6151
R993 B.n514 B.n260 10.6151
R994 B.n524 B.n260 10.6151
R995 B.n525 B.n524 10.6151
R996 B.n526 B.n525 10.6151
R997 B.n526 B.n253 10.6151
R998 B.n536 B.n253 10.6151
R999 B.n537 B.n536 10.6151
R1000 B.n538 B.n537 10.6151
R1001 B.n538 B.n245 10.6151
R1002 B.n548 B.n245 10.6151
R1003 B.n549 B.n548 10.6151
R1004 B.n551 B.n549 10.6151
R1005 B.n551 B.n550 10.6151
R1006 B.n550 B.n237 10.6151
R1007 B.n562 B.n237 10.6151
R1008 B.n563 B.n562 10.6151
R1009 B.n564 B.n563 10.6151
R1010 B.n565 B.n564 10.6151
R1011 B.n567 B.n565 10.6151
R1012 B.n568 B.n567 10.6151
R1013 B.n569 B.n568 10.6151
R1014 B.n570 B.n569 10.6151
R1015 B.n572 B.n570 10.6151
R1016 B.n573 B.n572 10.6151
R1017 B.n574 B.n573 10.6151
R1018 B.n575 B.n574 10.6151
R1019 B.n577 B.n575 10.6151
R1020 B.n578 B.n577 10.6151
R1021 B.n579 B.n578 10.6151
R1022 B.n580 B.n579 10.6151
R1023 B.n582 B.n580 10.6151
R1024 B.n583 B.n582 10.6151
R1025 B.n584 B.n583 10.6151
R1026 B.n585 B.n584 10.6151
R1027 B.n587 B.n585 10.6151
R1028 B.n588 B.n587 10.6151
R1029 B.n589 B.n588 10.6151
R1030 B.n590 B.n589 10.6151
R1031 B.n592 B.n590 10.6151
R1032 B.n593 B.n592 10.6151
R1033 B.n594 B.n593 10.6151
R1034 B.n595 B.n594 10.6151
R1035 B.n597 B.n595 10.6151
R1036 B.n598 B.n597 10.6151
R1037 B.n599 B.n598 10.6151
R1038 B.n469 B.n468 10.6151
R1039 B.n468 B.n467 10.6151
R1040 B.n467 B.n466 10.6151
R1041 B.n466 B.n464 10.6151
R1042 B.n464 B.n461 10.6151
R1043 B.n461 B.n460 10.6151
R1044 B.n460 B.n457 10.6151
R1045 B.n457 B.n456 10.6151
R1046 B.n456 B.n453 10.6151
R1047 B.n453 B.n452 10.6151
R1048 B.n452 B.n449 10.6151
R1049 B.n449 B.n448 10.6151
R1050 B.n448 B.n445 10.6151
R1051 B.n445 B.n444 10.6151
R1052 B.n444 B.n441 10.6151
R1053 B.n441 B.n440 10.6151
R1054 B.n440 B.n437 10.6151
R1055 B.n437 B.n436 10.6151
R1056 B.n436 B.n433 10.6151
R1057 B.n433 B.n432 10.6151
R1058 B.n432 B.n429 10.6151
R1059 B.n429 B.n428 10.6151
R1060 B.n428 B.n425 10.6151
R1061 B.n425 B.n424 10.6151
R1062 B.n424 B.n421 10.6151
R1063 B.n421 B.n420 10.6151
R1064 B.n420 B.n417 10.6151
R1065 B.n417 B.n416 10.6151
R1066 B.n416 B.n413 10.6151
R1067 B.n413 B.n412 10.6151
R1068 B.n409 B.n408 10.6151
R1069 B.n408 B.n405 10.6151
R1070 B.n405 B.n404 10.6151
R1071 B.n404 B.n401 10.6151
R1072 B.n401 B.n400 10.6151
R1073 B.n400 B.n397 10.6151
R1074 B.n397 B.n396 10.6151
R1075 B.n396 B.n393 10.6151
R1076 B.n391 B.n388 10.6151
R1077 B.n388 B.n387 10.6151
R1078 B.n387 B.n384 10.6151
R1079 B.n384 B.n383 10.6151
R1080 B.n383 B.n380 10.6151
R1081 B.n380 B.n379 10.6151
R1082 B.n379 B.n376 10.6151
R1083 B.n376 B.n375 10.6151
R1084 B.n375 B.n372 10.6151
R1085 B.n372 B.n371 10.6151
R1086 B.n371 B.n368 10.6151
R1087 B.n368 B.n367 10.6151
R1088 B.n367 B.n364 10.6151
R1089 B.n364 B.n363 10.6151
R1090 B.n363 B.n360 10.6151
R1091 B.n360 B.n359 10.6151
R1092 B.n359 B.n356 10.6151
R1093 B.n356 B.n355 10.6151
R1094 B.n355 B.n352 10.6151
R1095 B.n352 B.n351 10.6151
R1096 B.n351 B.n348 10.6151
R1097 B.n348 B.n347 10.6151
R1098 B.n347 B.n344 10.6151
R1099 B.n344 B.n343 10.6151
R1100 B.n343 B.n340 10.6151
R1101 B.n340 B.n339 10.6151
R1102 B.n339 B.n336 10.6151
R1103 B.n336 B.n335 10.6151
R1104 B.n335 B.n292 10.6151
R1105 B.n475 B.n292 10.6151
R1106 B.n481 B.n288 10.6151
R1107 B.n482 B.n481 10.6151
R1108 B.n483 B.n482 10.6151
R1109 B.n483 B.n280 10.6151
R1110 B.n494 B.n280 10.6151
R1111 B.n495 B.n494 10.6151
R1112 B.n496 B.n495 10.6151
R1113 B.n496 B.n273 10.6151
R1114 B.n506 B.n273 10.6151
R1115 B.n507 B.n506 10.6151
R1116 B.n508 B.n507 10.6151
R1117 B.n508 B.n265 10.6151
R1118 B.n518 B.n265 10.6151
R1119 B.n519 B.n518 10.6151
R1120 B.n520 B.n519 10.6151
R1121 B.n520 B.n257 10.6151
R1122 B.n530 B.n257 10.6151
R1123 B.n531 B.n530 10.6151
R1124 B.n532 B.n531 10.6151
R1125 B.n532 B.n249 10.6151
R1126 B.n542 B.n249 10.6151
R1127 B.n543 B.n542 10.6151
R1128 B.n544 B.n543 10.6151
R1129 B.n544 B.n241 10.6151
R1130 B.n555 B.n241 10.6151
R1131 B.n556 B.n555 10.6151
R1132 B.n557 B.n556 10.6151
R1133 B.n557 B.n0 10.6151
R1134 B.n656 B.n1 10.6151
R1135 B.n656 B.n655 10.6151
R1136 B.n655 B.n654 10.6151
R1137 B.n654 B.n10 10.6151
R1138 B.n648 B.n10 10.6151
R1139 B.n648 B.n647 10.6151
R1140 B.n647 B.n646 10.6151
R1141 B.n646 B.n17 10.6151
R1142 B.n640 B.n17 10.6151
R1143 B.n640 B.n639 10.6151
R1144 B.n639 B.n638 10.6151
R1145 B.n638 B.n24 10.6151
R1146 B.n632 B.n24 10.6151
R1147 B.n632 B.n631 10.6151
R1148 B.n631 B.n630 10.6151
R1149 B.n630 B.n31 10.6151
R1150 B.n624 B.n31 10.6151
R1151 B.n624 B.n623 10.6151
R1152 B.n623 B.n622 10.6151
R1153 B.n622 B.n38 10.6151
R1154 B.n616 B.n38 10.6151
R1155 B.n616 B.n615 10.6151
R1156 B.n615 B.n614 10.6151
R1157 B.n614 B.n44 10.6151
R1158 B.n608 B.n44 10.6151
R1159 B.n608 B.n607 10.6151
R1160 B.n607 B.n606 10.6151
R1161 B.n606 B.n52 10.6151
R1162 B.n528 B.t3 8.12758
R1163 B.n636 B.t0 8.12758
R1164 B.n160 B.n159 6.5566
R1165 B.n176 B.n94 6.5566
R1166 B.n409 B.n331 6.5566
R1167 B.n393 B.n392 6.5566
R1168 B.t2 B.n243 6.50216
R1169 B.n651 B.t1 6.50216
R1170 B.n159 B.n158 4.05904
R1171 B.n179 B.n94 4.05904
R1172 B.n412 B.n331 4.05904
R1173 B.n392 B.n391 4.05904
R1174 B.n662 B.n0 2.81026
R1175 B.n662 B.n1 2.81026
R1176 VN.n0 VN.t1 132.62
R1177 VN.n1 VN.t2 132.62
R1178 VN.n0 VN.t3 132.078
R1179 VN.n1 VN.t0 132.078
R1180 VN VN.n1 49.1447
R1181 VN VN.n0 7.03488
R1182 VDD2.n2 VDD2.n0 102.651
R1183 VDD2.n2 VDD2.n1 65.635
R1184 VDD2.n1 VDD2.t3 2.39759
R1185 VDD2.n1 VDD2.t1 2.39759
R1186 VDD2.n0 VDD2.t2 2.39759
R1187 VDD2.n0 VDD2.t0 2.39759
R1188 VDD2 VDD2.n2 0.0586897
C0 VP VDD1 3.42436f
C1 VTAIL VP 3.22566f
C2 VDD2 VN 3.21353f
C3 VTAIL VDD1 4.39904f
C4 VP VN 5.105f
C5 VN VDD1 0.148972f
C6 VP VDD2 0.360404f
C7 VTAIL VN 3.21155f
C8 VDD2 VDD1 0.898815f
C9 VTAIL VDD2 4.44963f
C10 VDD2 B 3.169241f
C11 VDD1 B 6.72363f
C12 VTAIL B 7.535985f
C13 VN B 9.37871f
C14 VP B 7.538539f
C15 VDD2.t2 B 0.174579f
C16 VDD2.t0 B 0.174579f
C17 VDD2.n0 B 2.01337f
C18 VDD2.t3 B 0.174579f
C19 VDD2.t1 B 0.174579f
C20 VDD2.n1 B 1.51626f
C21 VDD2.n2 B 3.18874f
C22 VN.t1 B 1.58167f
C23 VN.t3 B 1.57892f
C24 VN.n0 B 1.06826f
C25 VN.t2 B 1.58167f
C26 VN.t0 B 1.57892f
C27 VN.n1 B 2.36048f
C28 VDD1.t1 B 0.176874f
C29 VDD1.t3 B 0.176874f
C30 VDD1.n0 B 1.53655f
C31 VDD1.t0 B 0.176874f
C32 VDD1.t2 B 0.176874f
C33 VDD1.n1 B 2.06425f
C34 VTAIL.t1 B 1.18749f
C35 VTAIL.n0 B 0.298961f
C36 VTAIL.t6 B 1.18749f
C37 VTAIL.n1 B 0.353021f
C38 VTAIL.t7 B 1.18749f
C39 VTAIL.n2 B 1.072f
C40 VTAIL.t3 B 1.1875f
C41 VTAIL.n3 B 1.07199f
C42 VTAIL.t2 B 1.1875f
C43 VTAIL.n4 B 0.353013f
C44 VTAIL.t4 B 1.1875f
C45 VTAIL.n5 B 0.353013f
C46 VTAIL.t5 B 1.18749f
C47 VTAIL.n6 B 1.072f
C48 VTAIL.t0 B 1.18749f
C49 VTAIL.n7 B 1.01146f
C50 VP.n0 B 0.041105f
C51 VP.t1 B 1.42684f
C52 VP.n1 B 0.045325f
C53 VP.t0 B 1.61239f
C54 VP.t2 B 1.6152f
C55 VP.n2 B 2.39447f
C56 VP.n3 B 1.55265f
C57 VP.t3 B 1.42684f
C58 VP.n4 B 0.625849f
C59 VP.n5 B 0.054681f
C60 VP.n6 B 0.041105f
C61 VP.n7 B 0.03118f
C62 VP.n8 B 0.03118f
C63 VP.n9 B 0.045325f
C64 VP.n10 B 0.054681f
C65 VP.n11 B 0.625849f
C66 VP.n12 B 0.036211f
.ends

