* NGSPICE file created from diff_pair_sample_0514.ext - technology: sky130A

.subckt diff_pair_sample_0514 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.77
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.77
X2 B.t8 B.t6 B.t7 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.77
X3 B.t5 B.t3 B.t4 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.77
X4 VDD2.t1 VN.t0 VTAIL.t0 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.77
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.77
X6 B.t2 B.t0 B.t1 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.77
X7 VDD1.t0 VP.t1 VTAIL.t2 w_n1810_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.77
R0 B.n289 B.n288 585
R1 B.n287 B.n80 585
R2 B.n286 B.n285 585
R3 B.n284 B.n81 585
R4 B.n283 B.n282 585
R5 B.n281 B.n82 585
R6 B.n280 B.n279 585
R7 B.n278 B.n83 585
R8 B.n277 B.n276 585
R9 B.n275 B.n84 585
R10 B.n274 B.n273 585
R11 B.n272 B.n85 585
R12 B.n271 B.n270 585
R13 B.n269 B.n86 585
R14 B.n268 B.n267 585
R15 B.n266 B.n87 585
R16 B.n265 B.n264 585
R17 B.n263 B.n88 585
R18 B.n262 B.n261 585
R19 B.n260 B.n89 585
R20 B.n259 B.n258 585
R21 B.n257 B.n90 585
R22 B.n256 B.n255 585
R23 B.n254 B.n91 585
R24 B.n253 B.n252 585
R25 B.n251 B.n92 585
R26 B.n250 B.n249 585
R27 B.n248 B.n93 585
R28 B.n247 B.n246 585
R29 B.n245 B.n94 585
R30 B.n244 B.n243 585
R31 B.n242 B.n95 585
R32 B.n241 B.n240 585
R33 B.n239 B.n96 585
R34 B.n238 B.n237 585
R35 B.n236 B.n97 585
R36 B.n235 B.n234 585
R37 B.n232 B.n98 585
R38 B.n231 B.n230 585
R39 B.n229 B.n101 585
R40 B.n228 B.n227 585
R41 B.n226 B.n102 585
R42 B.n225 B.n224 585
R43 B.n223 B.n103 585
R44 B.n222 B.n221 585
R45 B.n220 B.n104 585
R46 B.n218 B.n217 585
R47 B.n216 B.n107 585
R48 B.n215 B.n214 585
R49 B.n213 B.n108 585
R50 B.n212 B.n211 585
R51 B.n210 B.n109 585
R52 B.n209 B.n208 585
R53 B.n207 B.n110 585
R54 B.n206 B.n205 585
R55 B.n204 B.n111 585
R56 B.n203 B.n202 585
R57 B.n201 B.n112 585
R58 B.n200 B.n199 585
R59 B.n198 B.n113 585
R60 B.n197 B.n196 585
R61 B.n195 B.n114 585
R62 B.n194 B.n193 585
R63 B.n192 B.n115 585
R64 B.n191 B.n190 585
R65 B.n189 B.n116 585
R66 B.n188 B.n187 585
R67 B.n186 B.n117 585
R68 B.n185 B.n184 585
R69 B.n183 B.n118 585
R70 B.n182 B.n181 585
R71 B.n180 B.n119 585
R72 B.n179 B.n178 585
R73 B.n177 B.n120 585
R74 B.n176 B.n175 585
R75 B.n174 B.n121 585
R76 B.n173 B.n172 585
R77 B.n171 B.n122 585
R78 B.n170 B.n169 585
R79 B.n168 B.n123 585
R80 B.n167 B.n166 585
R81 B.n165 B.n124 585
R82 B.n164 B.n163 585
R83 B.n290 B.n79 585
R84 B.n292 B.n291 585
R85 B.n293 B.n78 585
R86 B.n295 B.n294 585
R87 B.n296 B.n77 585
R88 B.n298 B.n297 585
R89 B.n299 B.n76 585
R90 B.n301 B.n300 585
R91 B.n302 B.n75 585
R92 B.n304 B.n303 585
R93 B.n305 B.n74 585
R94 B.n307 B.n306 585
R95 B.n308 B.n73 585
R96 B.n310 B.n309 585
R97 B.n311 B.n72 585
R98 B.n313 B.n312 585
R99 B.n314 B.n71 585
R100 B.n316 B.n315 585
R101 B.n317 B.n70 585
R102 B.n319 B.n318 585
R103 B.n320 B.n69 585
R104 B.n322 B.n321 585
R105 B.n323 B.n68 585
R106 B.n325 B.n324 585
R107 B.n326 B.n67 585
R108 B.n328 B.n327 585
R109 B.n329 B.n66 585
R110 B.n331 B.n330 585
R111 B.n332 B.n65 585
R112 B.n334 B.n333 585
R113 B.n335 B.n64 585
R114 B.n337 B.n336 585
R115 B.n338 B.n63 585
R116 B.n340 B.n339 585
R117 B.n341 B.n62 585
R118 B.n343 B.n342 585
R119 B.n344 B.n61 585
R120 B.n346 B.n345 585
R121 B.n347 B.n60 585
R122 B.n349 B.n348 585
R123 B.n350 B.n59 585
R124 B.n352 B.n351 585
R125 B.n477 B.n12 585
R126 B.n476 B.n475 585
R127 B.n474 B.n13 585
R128 B.n473 B.n472 585
R129 B.n471 B.n14 585
R130 B.n470 B.n469 585
R131 B.n468 B.n15 585
R132 B.n467 B.n466 585
R133 B.n465 B.n16 585
R134 B.n464 B.n463 585
R135 B.n462 B.n17 585
R136 B.n461 B.n460 585
R137 B.n459 B.n18 585
R138 B.n458 B.n457 585
R139 B.n456 B.n19 585
R140 B.n455 B.n454 585
R141 B.n453 B.n20 585
R142 B.n452 B.n451 585
R143 B.n450 B.n21 585
R144 B.n449 B.n448 585
R145 B.n447 B.n22 585
R146 B.n446 B.n445 585
R147 B.n444 B.n23 585
R148 B.n443 B.n442 585
R149 B.n441 B.n24 585
R150 B.n440 B.n439 585
R151 B.n438 B.n25 585
R152 B.n437 B.n436 585
R153 B.n435 B.n26 585
R154 B.n434 B.n433 585
R155 B.n432 B.n27 585
R156 B.n431 B.n430 585
R157 B.n429 B.n28 585
R158 B.n428 B.n427 585
R159 B.n426 B.n29 585
R160 B.n425 B.n424 585
R161 B.n423 B.n30 585
R162 B.n422 B.n421 585
R163 B.n420 B.n31 585
R164 B.n419 B.n418 585
R165 B.n417 B.n35 585
R166 B.n416 B.n415 585
R167 B.n414 B.n36 585
R168 B.n413 B.n412 585
R169 B.n411 B.n37 585
R170 B.n410 B.n409 585
R171 B.n407 B.n38 585
R172 B.n406 B.n405 585
R173 B.n404 B.n41 585
R174 B.n403 B.n402 585
R175 B.n401 B.n42 585
R176 B.n400 B.n399 585
R177 B.n398 B.n43 585
R178 B.n397 B.n396 585
R179 B.n395 B.n44 585
R180 B.n394 B.n393 585
R181 B.n392 B.n45 585
R182 B.n391 B.n390 585
R183 B.n389 B.n46 585
R184 B.n388 B.n387 585
R185 B.n386 B.n47 585
R186 B.n385 B.n384 585
R187 B.n383 B.n48 585
R188 B.n382 B.n381 585
R189 B.n380 B.n49 585
R190 B.n379 B.n378 585
R191 B.n377 B.n50 585
R192 B.n376 B.n375 585
R193 B.n374 B.n51 585
R194 B.n373 B.n372 585
R195 B.n371 B.n52 585
R196 B.n370 B.n369 585
R197 B.n368 B.n53 585
R198 B.n367 B.n366 585
R199 B.n365 B.n54 585
R200 B.n364 B.n363 585
R201 B.n362 B.n55 585
R202 B.n361 B.n360 585
R203 B.n359 B.n56 585
R204 B.n358 B.n357 585
R205 B.n356 B.n57 585
R206 B.n355 B.n354 585
R207 B.n353 B.n58 585
R208 B.n479 B.n478 585
R209 B.n480 B.n11 585
R210 B.n482 B.n481 585
R211 B.n483 B.n10 585
R212 B.n485 B.n484 585
R213 B.n486 B.n9 585
R214 B.n488 B.n487 585
R215 B.n489 B.n8 585
R216 B.n491 B.n490 585
R217 B.n492 B.n7 585
R218 B.n494 B.n493 585
R219 B.n495 B.n6 585
R220 B.n497 B.n496 585
R221 B.n498 B.n5 585
R222 B.n500 B.n499 585
R223 B.n501 B.n4 585
R224 B.n503 B.n502 585
R225 B.n504 B.n3 585
R226 B.n506 B.n505 585
R227 B.n507 B.n0 585
R228 B.n2 B.n1 585
R229 B.n135 B.n134 585
R230 B.n137 B.n136 585
R231 B.n138 B.n133 585
R232 B.n140 B.n139 585
R233 B.n141 B.n132 585
R234 B.n143 B.n142 585
R235 B.n144 B.n131 585
R236 B.n146 B.n145 585
R237 B.n147 B.n130 585
R238 B.n149 B.n148 585
R239 B.n150 B.n129 585
R240 B.n152 B.n151 585
R241 B.n153 B.n128 585
R242 B.n155 B.n154 585
R243 B.n156 B.n127 585
R244 B.n158 B.n157 585
R245 B.n159 B.n126 585
R246 B.n161 B.n160 585
R247 B.n162 B.n125 585
R248 B.n163 B.n162 506.916
R249 B.n290 B.n289 506.916
R250 B.n351 B.n58 506.916
R251 B.n478 B.n477 506.916
R252 B.n105 B.t0 347.382
R253 B.n99 B.t9 347.382
R254 B.n39 B.t3 347.382
R255 B.n32 B.t6 347.382
R256 B.n509 B.n508 256.663
R257 B.n508 B.n507 235.042
R258 B.n508 B.n2 235.042
R259 B.n163 B.n124 163.367
R260 B.n167 B.n124 163.367
R261 B.n168 B.n167 163.367
R262 B.n169 B.n168 163.367
R263 B.n169 B.n122 163.367
R264 B.n173 B.n122 163.367
R265 B.n174 B.n173 163.367
R266 B.n175 B.n174 163.367
R267 B.n175 B.n120 163.367
R268 B.n179 B.n120 163.367
R269 B.n180 B.n179 163.367
R270 B.n181 B.n180 163.367
R271 B.n181 B.n118 163.367
R272 B.n185 B.n118 163.367
R273 B.n186 B.n185 163.367
R274 B.n187 B.n186 163.367
R275 B.n187 B.n116 163.367
R276 B.n191 B.n116 163.367
R277 B.n192 B.n191 163.367
R278 B.n193 B.n192 163.367
R279 B.n193 B.n114 163.367
R280 B.n197 B.n114 163.367
R281 B.n198 B.n197 163.367
R282 B.n199 B.n198 163.367
R283 B.n199 B.n112 163.367
R284 B.n203 B.n112 163.367
R285 B.n204 B.n203 163.367
R286 B.n205 B.n204 163.367
R287 B.n205 B.n110 163.367
R288 B.n209 B.n110 163.367
R289 B.n210 B.n209 163.367
R290 B.n211 B.n210 163.367
R291 B.n211 B.n108 163.367
R292 B.n215 B.n108 163.367
R293 B.n216 B.n215 163.367
R294 B.n217 B.n216 163.367
R295 B.n217 B.n104 163.367
R296 B.n222 B.n104 163.367
R297 B.n223 B.n222 163.367
R298 B.n224 B.n223 163.367
R299 B.n224 B.n102 163.367
R300 B.n228 B.n102 163.367
R301 B.n229 B.n228 163.367
R302 B.n230 B.n229 163.367
R303 B.n230 B.n98 163.367
R304 B.n235 B.n98 163.367
R305 B.n236 B.n235 163.367
R306 B.n237 B.n236 163.367
R307 B.n237 B.n96 163.367
R308 B.n241 B.n96 163.367
R309 B.n242 B.n241 163.367
R310 B.n243 B.n242 163.367
R311 B.n243 B.n94 163.367
R312 B.n247 B.n94 163.367
R313 B.n248 B.n247 163.367
R314 B.n249 B.n248 163.367
R315 B.n249 B.n92 163.367
R316 B.n253 B.n92 163.367
R317 B.n254 B.n253 163.367
R318 B.n255 B.n254 163.367
R319 B.n255 B.n90 163.367
R320 B.n259 B.n90 163.367
R321 B.n260 B.n259 163.367
R322 B.n261 B.n260 163.367
R323 B.n261 B.n88 163.367
R324 B.n265 B.n88 163.367
R325 B.n266 B.n265 163.367
R326 B.n267 B.n266 163.367
R327 B.n267 B.n86 163.367
R328 B.n271 B.n86 163.367
R329 B.n272 B.n271 163.367
R330 B.n273 B.n272 163.367
R331 B.n273 B.n84 163.367
R332 B.n277 B.n84 163.367
R333 B.n278 B.n277 163.367
R334 B.n279 B.n278 163.367
R335 B.n279 B.n82 163.367
R336 B.n283 B.n82 163.367
R337 B.n284 B.n283 163.367
R338 B.n285 B.n284 163.367
R339 B.n285 B.n80 163.367
R340 B.n289 B.n80 163.367
R341 B.n351 B.n350 163.367
R342 B.n350 B.n349 163.367
R343 B.n349 B.n60 163.367
R344 B.n345 B.n60 163.367
R345 B.n345 B.n344 163.367
R346 B.n344 B.n343 163.367
R347 B.n343 B.n62 163.367
R348 B.n339 B.n62 163.367
R349 B.n339 B.n338 163.367
R350 B.n338 B.n337 163.367
R351 B.n337 B.n64 163.367
R352 B.n333 B.n64 163.367
R353 B.n333 B.n332 163.367
R354 B.n332 B.n331 163.367
R355 B.n331 B.n66 163.367
R356 B.n327 B.n66 163.367
R357 B.n327 B.n326 163.367
R358 B.n326 B.n325 163.367
R359 B.n325 B.n68 163.367
R360 B.n321 B.n68 163.367
R361 B.n321 B.n320 163.367
R362 B.n320 B.n319 163.367
R363 B.n319 B.n70 163.367
R364 B.n315 B.n70 163.367
R365 B.n315 B.n314 163.367
R366 B.n314 B.n313 163.367
R367 B.n313 B.n72 163.367
R368 B.n309 B.n72 163.367
R369 B.n309 B.n308 163.367
R370 B.n308 B.n307 163.367
R371 B.n307 B.n74 163.367
R372 B.n303 B.n74 163.367
R373 B.n303 B.n302 163.367
R374 B.n302 B.n301 163.367
R375 B.n301 B.n76 163.367
R376 B.n297 B.n76 163.367
R377 B.n297 B.n296 163.367
R378 B.n296 B.n295 163.367
R379 B.n295 B.n78 163.367
R380 B.n291 B.n78 163.367
R381 B.n291 B.n290 163.367
R382 B.n477 B.n476 163.367
R383 B.n476 B.n13 163.367
R384 B.n472 B.n13 163.367
R385 B.n472 B.n471 163.367
R386 B.n471 B.n470 163.367
R387 B.n470 B.n15 163.367
R388 B.n466 B.n15 163.367
R389 B.n466 B.n465 163.367
R390 B.n465 B.n464 163.367
R391 B.n464 B.n17 163.367
R392 B.n460 B.n17 163.367
R393 B.n460 B.n459 163.367
R394 B.n459 B.n458 163.367
R395 B.n458 B.n19 163.367
R396 B.n454 B.n19 163.367
R397 B.n454 B.n453 163.367
R398 B.n453 B.n452 163.367
R399 B.n452 B.n21 163.367
R400 B.n448 B.n21 163.367
R401 B.n448 B.n447 163.367
R402 B.n447 B.n446 163.367
R403 B.n446 B.n23 163.367
R404 B.n442 B.n23 163.367
R405 B.n442 B.n441 163.367
R406 B.n441 B.n440 163.367
R407 B.n440 B.n25 163.367
R408 B.n436 B.n25 163.367
R409 B.n436 B.n435 163.367
R410 B.n435 B.n434 163.367
R411 B.n434 B.n27 163.367
R412 B.n430 B.n27 163.367
R413 B.n430 B.n429 163.367
R414 B.n429 B.n428 163.367
R415 B.n428 B.n29 163.367
R416 B.n424 B.n29 163.367
R417 B.n424 B.n423 163.367
R418 B.n423 B.n422 163.367
R419 B.n422 B.n31 163.367
R420 B.n418 B.n31 163.367
R421 B.n418 B.n417 163.367
R422 B.n417 B.n416 163.367
R423 B.n416 B.n36 163.367
R424 B.n412 B.n36 163.367
R425 B.n412 B.n411 163.367
R426 B.n411 B.n410 163.367
R427 B.n410 B.n38 163.367
R428 B.n405 B.n38 163.367
R429 B.n405 B.n404 163.367
R430 B.n404 B.n403 163.367
R431 B.n403 B.n42 163.367
R432 B.n399 B.n42 163.367
R433 B.n399 B.n398 163.367
R434 B.n398 B.n397 163.367
R435 B.n397 B.n44 163.367
R436 B.n393 B.n44 163.367
R437 B.n393 B.n392 163.367
R438 B.n392 B.n391 163.367
R439 B.n391 B.n46 163.367
R440 B.n387 B.n46 163.367
R441 B.n387 B.n386 163.367
R442 B.n386 B.n385 163.367
R443 B.n385 B.n48 163.367
R444 B.n381 B.n48 163.367
R445 B.n381 B.n380 163.367
R446 B.n380 B.n379 163.367
R447 B.n379 B.n50 163.367
R448 B.n375 B.n50 163.367
R449 B.n375 B.n374 163.367
R450 B.n374 B.n373 163.367
R451 B.n373 B.n52 163.367
R452 B.n369 B.n52 163.367
R453 B.n369 B.n368 163.367
R454 B.n368 B.n367 163.367
R455 B.n367 B.n54 163.367
R456 B.n363 B.n54 163.367
R457 B.n363 B.n362 163.367
R458 B.n362 B.n361 163.367
R459 B.n361 B.n56 163.367
R460 B.n357 B.n56 163.367
R461 B.n357 B.n356 163.367
R462 B.n356 B.n355 163.367
R463 B.n355 B.n58 163.367
R464 B.n478 B.n11 163.367
R465 B.n482 B.n11 163.367
R466 B.n483 B.n482 163.367
R467 B.n484 B.n483 163.367
R468 B.n484 B.n9 163.367
R469 B.n488 B.n9 163.367
R470 B.n489 B.n488 163.367
R471 B.n490 B.n489 163.367
R472 B.n490 B.n7 163.367
R473 B.n494 B.n7 163.367
R474 B.n495 B.n494 163.367
R475 B.n496 B.n495 163.367
R476 B.n496 B.n5 163.367
R477 B.n500 B.n5 163.367
R478 B.n501 B.n500 163.367
R479 B.n502 B.n501 163.367
R480 B.n502 B.n3 163.367
R481 B.n506 B.n3 163.367
R482 B.n507 B.n506 163.367
R483 B.n134 B.n2 163.367
R484 B.n137 B.n134 163.367
R485 B.n138 B.n137 163.367
R486 B.n139 B.n138 163.367
R487 B.n139 B.n132 163.367
R488 B.n143 B.n132 163.367
R489 B.n144 B.n143 163.367
R490 B.n145 B.n144 163.367
R491 B.n145 B.n130 163.367
R492 B.n149 B.n130 163.367
R493 B.n150 B.n149 163.367
R494 B.n151 B.n150 163.367
R495 B.n151 B.n128 163.367
R496 B.n155 B.n128 163.367
R497 B.n156 B.n155 163.367
R498 B.n157 B.n156 163.367
R499 B.n157 B.n126 163.367
R500 B.n161 B.n126 163.367
R501 B.n162 B.n161 163.367
R502 B.n99 B.t10 151.385
R503 B.n39 B.t5 151.385
R504 B.n105 B.t1 151.373
R505 B.n32 B.t8 151.373
R506 B.n100 B.t11 110.656
R507 B.n40 B.t4 110.656
R508 B.n106 B.t2 110.644
R509 B.n33 B.t7 110.644
R510 B.n219 B.n106 59.5399
R511 B.n233 B.n100 59.5399
R512 B.n408 B.n40 59.5399
R513 B.n34 B.n33 59.5399
R514 B.n106 B.n105 40.7278
R515 B.n100 B.n99 40.7278
R516 B.n40 B.n39 40.7278
R517 B.n33 B.n32 40.7278
R518 B.n479 B.n12 32.9371
R519 B.n353 B.n352 32.9371
R520 B.n288 B.n79 32.9371
R521 B.n164 B.n125 32.9371
R522 B B.n509 18.0485
R523 B.n480 B.n479 10.6151
R524 B.n481 B.n480 10.6151
R525 B.n481 B.n10 10.6151
R526 B.n485 B.n10 10.6151
R527 B.n486 B.n485 10.6151
R528 B.n487 B.n486 10.6151
R529 B.n487 B.n8 10.6151
R530 B.n491 B.n8 10.6151
R531 B.n492 B.n491 10.6151
R532 B.n493 B.n492 10.6151
R533 B.n493 B.n6 10.6151
R534 B.n497 B.n6 10.6151
R535 B.n498 B.n497 10.6151
R536 B.n499 B.n498 10.6151
R537 B.n499 B.n4 10.6151
R538 B.n503 B.n4 10.6151
R539 B.n504 B.n503 10.6151
R540 B.n505 B.n504 10.6151
R541 B.n505 B.n0 10.6151
R542 B.n475 B.n12 10.6151
R543 B.n475 B.n474 10.6151
R544 B.n474 B.n473 10.6151
R545 B.n473 B.n14 10.6151
R546 B.n469 B.n14 10.6151
R547 B.n469 B.n468 10.6151
R548 B.n468 B.n467 10.6151
R549 B.n467 B.n16 10.6151
R550 B.n463 B.n16 10.6151
R551 B.n463 B.n462 10.6151
R552 B.n462 B.n461 10.6151
R553 B.n461 B.n18 10.6151
R554 B.n457 B.n18 10.6151
R555 B.n457 B.n456 10.6151
R556 B.n456 B.n455 10.6151
R557 B.n455 B.n20 10.6151
R558 B.n451 B.n20 10.6151
R559 B.n451 B.n450 10.6151
R560 B.n450 B.n449 10.6151
R561 B.n449 B.n22 10.6151
R562 B.n445 B.n22 10.6151
R563 B.n445 B.n444 10.6151
R564 B.n444 B.n443 10.6151
R565 B.n443 B.n24 10.6151
R566 B.n439 B.n24 10.6151
R567 B.n439 B.n438 10.6151
R568 B.n438 B.n437 10.6151
R569 B.n437 B.n26 10.6151
R570 B.n433 B.n26 10.6151
R571 B.n433 B.n432 10.6151
R572 B.n432 B.n431 10.6151
R573 B.n431 B.n28 10.6151
R574 B.n427 B.n28 10.6151
R575 B.n427 B.n426 10.6151
R576 B.n426 B.n425 10.6151
R577 B.n425 B.n30 10.6151
R578 B.n421 B.n420 10.6151
R579 B.n420 B.n419 10.6151
R580 B.n419 B.n35 10.6151
R581 B.n415 B.n35 10.6151
R582 B.n415 B.n414 10.6151
R583 B.n414 B.n413 10.6151
R584 B.n413 B.n37 10.6151
R585 B.n409 B.n37 10.6151
R586 B.n407 B.n406 10.6151
R587 B.n406 B.n41 10.6151
R588 B.n402 B.n41 10.6151
R589 B.n402 B.n401 10.6151
R590 B.n401 B.n400 10.6151
R591 B.n400 B.n43 10.6151
R592 B.n396 B.n43 10.6151
R593 B.n396 B.n395 10.6151
R594 B.n395 B.n394 10.6151
R595 B.n394 B.n45 10.6151
R596 B.n390 B.n45 10.6151
R597 B.n390 B.n389 10.6151
R598 B.n389 B.n388 10.6151
R599 B.n388 B.n47 10.6151
R600 B.n384 B.n47 10.6151
R601 B.n384 B.n383 10.6151
R602 B.n383 B.n382 10.6151
R603 B.n382 B.n49 10.6151
R604 B.n378 B.n49 10.6151
R605 B.n378 B.n377 10.6151
R606 B.n377 B.n376 10.6151
R607 B.n376 B.n51 10.6151
R608 B.n372 B.n51 10.6151
R609 B.n372 B.n371 10.6151
R610 B.n371 B.n370 10.6151
R611 B.n370 B.n53 10.6151
R612 B.n366 B.n53 10.6151
R613 B.n366 B.n365 10.6151
R614 B.n365 B.n364 10.6151
R615 B.n364 B.n55 10.6151
R616 B.n360 B.n55 10.6151
R617 B.n360 B.n359 10.6151
R618 B.n359 B.n358 10.6151
R619 B.n358 B.n57 10.6151
R620 B.n354 B.n57 10.6151
R621 B.n354 B.n353 10.6151
R622 B.n352 B.n59 10.6151
R623 B.n348 B.n59 10.6151
R624 B.n348 B.n347 10.6151
R625 B.n347 B.n346 10.6151
R626 B.n346 B.n61 10.6151
R627 B.n342 B.n61 10.6151
R628 B.n342 B.n341 10.6151
R629 B.n341 B.n340 10.6151
R630 B.n340 B.n63 10.6151
R631 B.n336 B.n63 10.6151
R632 B.n336 B.n335 10.6151
R633 B.n335 B.n334 10.6151
R634 B.n334 B.n65 10.6151
R635 B.n330 B.n65 10.6151
R636 B.n330 B.n329 10.6151
R637 B.n329 B.n328 10.6151
R638 B.n328 B.n67 10.6151
R639 B.n324 B.n67 10.6151
R640 B.n324 B.n323 10.6151
R641 B.n323 B.n322 10.6151
R642 B.n322 B.n69 10.6151
R643 B.n318 B.n69 10.6151
R644 B.n318 B.n317 10.6151
R645 B.n317 B.n316 10.6151
R646 B.n316 B.n71 10.6151
R647 B.n312 B.n71 10.6151
R648 B.n312 B.n311 10.6151
R649 B.n311 B.n310 10.6151
R650 B.n310 B.n73 10.6151
R651 B.n306 B.n73 10.6151
R652 B.n306 B.n305 10.6151
R653 B.n305 B.n304 10.6151
R654 B.n304 B.n75 10.6151
R655 B.n300 B.n75 10.6151
R656 B.n300 B.n299 10.6151
R657 B.n299 B.n298 10.6151
R658 B.n298 B.n77 10.6151
R659 B.n294 B.n77 10.6151
R660 B.n294 B.n293 10.6151
R661 B.n293 B.n292 10.6151
R662 B.n292 B.n79 10.6151
R663 B.n135 B.n1 10.6151
R664 B.n136 B.n135 10.6151
R665 B.n136 B.n133 10.6151
R666 B.n140 B.n133 10.6151
R667 B.n141 B.n140 10.6151
R668 B.n142 B.n141 10.6151
R669 B.n142 B.n131 10.6151
R670 B.n146 B.n131 10.6151
R671 B.n147 B.n146 10.6151
R672 B.n148 B.n147 10.6151
R673 B.n148 B.n129 10.6151
R674 B.n152 B.n129 10.6151
R675 B.n153 B.n152 10.6151
R676 B.n154 B.n153 10.6151
R677 B.n154 B.n127 10.6151
R678 B.n158 B.n127 10.6151
R679 B.n159 B.n158 10.6151
R680 B.n160 B.n159 10.6151
R681 B.n160 B.n125 10.6151
R682 B.n165 B.n164 10.6151
R683 B.n166 B.n165 10.6151
R684 B.n166 B.n123 10.6151
R685 B.n170 B.n123 10.6151
R686 B.n171 B.n170 10.6151
R687 B.n172 B.n171 10.6151
R688 B.n172 B.n121 10.6151
R689 B.n176 B.n121 10.6151
R690 B.n177 B.n176 10.6151
R691 B.n178 B.n177 10.6151
R692 B.n178 B.n119 10.6151
R693 B.n182 B.n119 10.6151
R694 B.n183 B.n182 10.6151
R695 B.n184 B.n183 10.6151
R696 B.n184 B.n117 10.6151
R697 B.n188 B.n117 10.6151
R698 B.n189 B.n188 10.6151
R699 B.n190 B.n189 10.6151
R700 B.n190 B.n115 10.6151
R701 B.n194 B.n115 10.6151
R702 B.n195 B.n194 10.6151
R703 B.n196 B.n195 10.6151
R704 B.n196 B.n113 10.6151
R705 B.n200 B.n113 10.6151
R706 B.n201 B.n200 10.6151
R707 B.n202 B.n201 10.6151
R708 B.n202 B.n111 10.6151
R709 B.n206 B.n111 10.6151
R710 B.n207 B.n206 10.6151
R711 B.n208 B.n207 10.6151
R712 B.n208 B.n109 10.6151
R713 B.n212 B.n109 10.6151
R714 B.n213 B.n212 10.6151
R715 B.n214 B.n213 10.6151
R716 B.n214 B.n107 10.6151
R717 B.n218 B.n107 10.6151
R718 B.n221 B.n220 10.6151
R719 B.n221 B.n103 10.6151
R720 B.n225 B.n103 10.6151
R721 B.n226 B.n225 10.6151
R722 B.n227 B.n226 10.6151
R723 B.n227 B.n101 10.6151
R724 B.n231 B.n101 10.6151
R725 B.n232 B.n231 10.6151
R726 B.n234 B.n97 10.6151
R727 B.n238 B.n97 10.6151
R728 B.n239 B.n238 10.6151
R729 B.n240 B.n239 10.6151
R730 B.n240 B.n95 10.6151
R731 B.n244 B.n95 10.6151
R732 B.n245 B.n244 10.6151
R733 B.n246 B.n245 10.6151
R734 B.n246 B.n93 10.6151
R735 B.n250 B.n93 10.6151
R736 B.n251 B.n250 10.6151
R737 B.n252 B.n251 10.6151
R738 B.n252 B.n91 10.6151
R739 B.n256 B.n91 10.6151
R740 B.n257 B.n256 10.6151
R741 B.n258 B.n257 10.6151
R742 B.n258 B.n89 10.6151
R743 B.n262 B.n89 10.6151
R744 B.n263 B.n262 10.6151
R745 B.n264 B.n263 10.6151
R746 B.n264 B.n87 10.6151
R747 B.n268 B.n87 10.6151
R748 B.n269 B.n268 10.6151
R749 B.n270 B.n269 10.6151
R750 B.n270 B.n85 10.6151
R751 B.n274 B.n85 10.6151
R752 B.n275 B.n274 10.6151
R753 B.n276 B.n275 10.6151
R754 B.n276 B.n83 10.6151
R755 B.n280 B.n83 10.6151
R756 B.n281 B.n280 10.6151
R757 B.n282 B.n281 10.6151
R758 B.n282 B.n81 10.6151
R759 B.n286 B.n81 10.6151
R760 B.n287 B.n286 10.6151
R761 B.n288 B.n287 10.6151
R762 B.n509 B.n0 8.11757
R763 B.n509 B.n1 8.11757
R764 B.n421 B.n34 6.5566
R765 B.n409 B.n408 6.5566
R766 B.n220 B.n219 6.5566
R767 B.n233 B.n232 6.5566
R768 B.n34 B.n30 4.05904
R769 B.n408 B.n407 4.05904
R770 B.n219 B.n218 4.05904
R771 B.n234 B.n233 4.05904
R772 VP.n0 VP.t1 241.16
R773 VP.n0 VP.t0 199.946
R774 VP VP.n0 0.241678
R775 VTAIL.n1 VTAIL.t0 63.7032
R776 VTAIL.n2 VTAIL.t2 63.703
R777 VTAIL.n3 VTAIL.t1 63.703
R778 VTAIL.n0 VTAIL.t3 63.703
R779 VTAIL.n1 VTAIL.n0 24.9186
R780 VTAIL.n3 VTAIL.n2 23.1083
R781 VTAIL.n2 VTAIL.n1 1.3755
R782 VTAIL VTAIL.n0 0.981103
R783 VTAIL VTAIL.n3 0.394897
R784 VDD1 VDD1.t1 117.57
R785 VDD1 VDD1.t0 80.8925
R786 VN VN.t0 241.351
R787 VN VN.t1 200.188
R788 VDD2.n0 VDD2.t0 116.593
R789 VDD2.n0 VDD2.t1 80.3818
R790 VDD2 VDD2.n0 0.511276
C0 w_n1810_n3040# VTAIL 2.53876f
C1 B VP 1.26622f
C2 B VN 0.893441f
C3 B VDD1 1.4628f
C4 VP VDD2 0.298444f
C5 VDD2 VN 2.2715f
C6 VDD2 VDD1 0.576498f
C7 B VDD2 1.48554f
C8 w_n1810_n3040# VP 2.62836f
C9 w_n1810_n3040# VN 2.39959f
C10 w_n1810_n3040# VDD1 1.57237f
C11 w_n1810_n3040# B 7.4524f
C12 w_n1810_n3040# VDD2 1.58827f
C13 VTAIL VP 1.96514f
C14 VTAIL VN 1.9508f
C15 VTAIL VDD1 4.5583f
C16 VTAIL B 2.94972f
C17 VTAIL VDD2 4.60273f
C18 VP VN 4.76128f
C19 VP VDD1 2.41917f
C20 VN VDD1 0.148075f
C21 VDD2 VSUBS 0.771135f
C22 VDD1 VSUBS 4.060982f
C23 VTAIL VSUBS 0.819879f
C24 VN VSUBS 6.48158f
C25 VP VSUBS 1.373274f
C26 B VSUBS 3.139782f
C27 w_n1810_n3040# VSUBS 67.9184f
C28 VDD2.t0 VSUBS 2.12682f
C29 VDD2.t1 VSUBS 1.66398f
C30 VDD2.n0 VSUBS 3.01567f
C31 VN.t1 VSUBS 2.31376f
C32 VN.t0 VSUBS 2.72621f
C33 VDD1.t0 VSUBS 1.67287f
C34 VDD1.t1 VSUBS 2.16207f
C35 VTAIL.t3 VSUBS 1.77162f
C36 VTAIL.n0 VSUBS 1.91665f
C37 VTAIL.t0 VSUBS 1.77163f
C38 VTAIL.n1 VSUBS 1.9462f
C39 VTAIL.t2 VSUBS 1.77162f
C40 VTAIL.n2 VSUBS 1.81055f
C41 VTAIL.t1 VSUBS 1.77162f
C42 VTAIL.n3 VSUBS 1.73707f
C43 VP.t1 VSUBS 2.82441f
C44 VP.t0 VSUBS 2.4004f
C45 VP.n0 VSUBS 4.51159f
C46 B.n0 VSUBS 0.006031f
C47 B.n1 VSUBS 0.006031f
C48 B.n2 VSUBS 0.00892f
C49 B.n3 VSUBS 0.006835f
C50 B.n4 VSUBS 0.006835f
C51 B.n5 VSUBS 0.006835f
C52 B.n6 VSUBS 0.006835f
C53 B.n7 VSUBS 0.006835f
C54 B.n8 VSUBS 0.006835f
C55 B.n9 VSUBS 0.006835f
C56 B.n10 VSUBS 0.006835f
C57 B.n11 VSUBS 0.006835f
C58 B.n12 VSUBS 0.016386f
C59 B.n13 VSUBS 0.006835f
C60 B.n14 VSUBS 0.006835f
C61 B.n15 VSUBS 0.006835f
C62 B.n16 VSUBS 0.006835f
C63 B.n17 VSUBS 0.006835f
C64 B.n18 VSUBS 0.006835f
C65 B.n19 VSUBS 0.006835f
C66 B.n20 VSUBS 0.006835f
C67 B.n21 VSUBS 0.006835f
C68 B.n22 VSUBS 0.006835f
C69 B.n23 VSUBS 0.006835f
C70 B.n24 VSUBS 0.006835f
C71 B.n25 VSUBS 0.006835f
C72 B.n26 VSUBS 0.006835f
C73 B.n27 VSUBS 0.006835f
C74 B.n28 VSUBS 0.006835f
C75 B.n29 VSUBS 0.006835f
C76 B.n30 VSUBS 0.004724f
C77 B.n31 VSUBS 0.006835f
C78 B.t7 VSUBS 0.32409f
C79 B.t8 VSUBS 0.339391f
C80 B.t6 VSUBS 0.801162f
C81 B.n32 VSUBS 0.161864f
C82 B.n33 VSUBS 0.066616f
C83 B.n34 VSUBS 0.015836f
C84 B.n35 VSUBS 0.006835f
C85 B.n36 VSUBS 0.006835f
C86 B.n37 VSUBS 0.006835f
C87 B.n38 VSUBS 0.006835f
C88 B.t4 VSUBS 0.324086f
C89 B.t5 VSUBS 0.339386f
C90 B.t3 VSUBS 0.801162f
C91 B.n39 VSUBS 0.161869f
C92 B.n40 VSUBS 0.066621f
C93 B.n41 VSUBS 0.006835f
C94 B.n42 VSUBS 0.006835f
C95 B.n43 VSUBS 0.006835f
C96 B.n44 VSUBS 0.006835f
C97 B.n45 VSUBS 0.006835f
C98 B.n46 VSUBS 0.006835f
C99 B.n47 VSUBS 0.006835f
C100 B.n48 VSUBS 0.006835f
C101 B.n49 VSUBS 0.006835f
C102 B.n50 VSUBS 0.006835f
C103 B.n51 VSUBS 0.006835f
C104 B.n52 VSUBS 0.006835f
C105 B.n53 VSUBS 0.006835f
C106 B.n54 VSUBS 0.006835f
C107 B.n55 VSUBS 0.006835f
C108 B.n56 VSUBS 0.006835f
C109 B.n57 VSUBS 0.006835f
C110 B.n58 VSUBS 0.016386f
C111 B.n59 VSUBS 0.006835f
C112 B.n60 VSUBS 0.006835f
C113 B.n61 VSUBS 0.006835f
C114 B.n62 VSUBS 0.006835f
C115 B.n63 VSUBS 0.006835f
C116 B.n64 VSUBS 0.006835f
C117 B.n65 VSUBS 0.006835f
C118 B.n66 VSUBS 0.006835f
C119 B.n67 VSUBS 0.006835f
C120 B.n68 VSUBS 0.006835f
C121 B.n69 VSUBS 0.006835f
C122 B.n70 VSUBS 0.006835f
C123 B.n71 VSUBS 0.006835f
C124 B.n72 VSUBS 0.006835f
C125 B.n73 VSUBS 0.006835f
C126 B.n74 VSUBS 0.006835f
C127 B.n75 VSUBS 0.006835f
C128 B.n76 VSUBS 0.006835f
C129 B.n77 VSUBS 0.006835f
C130 B.n78 VSUBS 0.006835f
C131 B.n79 VSUBS 0.016581f
C132 B.n80 VSUBS 0.006835f
C133 B.n81 VSUBS 0.006835f
C134 B.n82 VSUBS 0.006835f
C135 B.n83 VSUBS 0.006835f
C136 B.n84 VSUBS 0.006835f
C137 B.n85 VSUBS 0.006835f
C138 B.n86 VSUBS 0.006835f
C139 B.n87 VSUBS 0.006835f
C140 B.n88 VSUBS 0.006835f
C141 B.n89 VSUBS 0.006835f
C142 B.n90 VSUBS 0.006835f
C143 B.n91 VSUBS 0.006835f
C144 B.n92 VSUBS 0.006835f
C145 B.n93 VSUBS 0.006835f
C146 B.n94 VSUBS 0.006835f
C147 B.n95 VSUBS 0.006835f
C148 B.n96 VSUBS 0.006835f
C149 B.n97 VSUBS 0.006835f
C150 B.n98 VSUBS 0.006835f
C151 B.t11 VSUBS 0.324086f
C152 B.t10 VSUBS 0.339386f
C153 B.t9 VSUBS 0.801162f
C154 B.n99 VSUBS 0.161869f
C155 B.n100 VSUBS 0.066621f
C156 B.n101 VSUBS 0.006835f
C157 B.n102 VSUBS 0.006835f
C158 B.n103 VSUBS 0.006835f
C159 B.n104 VSUBS 0.006835f
C160 B.t2 VSUBS 0.32409f
C161 B.t1 VSUBS 0.339391f
C162 B.t0 VSUBS 0.801162f
C163 B.n105 VSUBS 0.161864f
C164 B.n106 VSUBS 0.066616f
C165 B.n107 VSUBS 0.006835f
C166 B.n108 VSUBS 0.006835f
C167 B.n109 VSUBS 0.006835f
C168 B.n110 VSUBS 0.006835f
C169 B.n111 VSUBS 0.006835f
C170 B.n112 VSUBS 0.006835f
C171 B.n113 VSUBS 0.006835f
C172 B.n114 VSUBS 0.006835f
C173 B.n115 VSUBS 0.006835f
C174 B.n116 VSUBS 0.006835f
C175 B.n117 VSUBS 0.006835f
C176 B.n118 VSUBS 0.006835f
C177 B.n119 VSUBS 0.006835f
C178 B.n120 VSUBS 0.006835f
C179 B.n121 VSUBS 0.006835f
C180 B.n122 VSUBS 0.006835f
C181 B.n123 VSUBS 0.006835f
C182 B.n124 VSUBS 0.006835f
C183 B.n125 VSUBS 0.01578f
C184 B.n126 VSUBS 0.006835f
C185 B.n127 VSUBS 0.006835f
C186 B.n128 VSUBS 0.006835f
C187 B.n129 VSUBS 0.006835f
C188 B.n130 VSUBS 0.006835f
C189 B.n131 VSUBS 0.006835f
C190 B.n132 VSUBS 0.006835f
C191 B.n133 VSUBS 0.006835f
C192 B.n134 VSUBS 0.006835f
C193 B.n135 VSUBS 0.006835f
C194 B.n136 VSUBS 0.006835f
C195 B.n137 VSUBS 0.006835f
C196 B.n138 VSUBS 0.006835f
C197 B.n139 VSUBS 0.006835f
C198 B.n140 VSUBS 0.006835f
C199 B.n141 VSUBS 0.006835f
C200 B.n142 VSUBS 0.006835f
C201 B.n143 VSUBS 0.006835f
C202 B.n144 VSUBS 0.006835f
C203 B.n145 VSUBS 0.006835f
C204 B.n146 VSUBS 0.006835f
C205 B.n147 VSUBS 0.006835f
C206 B.n148 VSUBS 0.006835f
C207 B.n149 VSUBS 0.006835f
C208 B.n150 VSUBS 0.006835f
C209 B.n151 VSUBS 0.006835f
C210 B.n152 VSUBS 0.006835f
C211 B.n153 VSUBS 0.006835f
C212 B.n154 VSUBS 0.006835f
C213 B.n155 VSUBS 0.006835f
C214 B.n156 VSUBS 0.006835f
C215 B.n157 VSUBS 0.006835f
C216 B.n158 VSUBS 0.006835f
C217 B.n159 VSUBS 0.006835f
C218 B.n160 VSUBS 0.006835f
C219 B.n161 VSUBS 0.006835f
C220 B.n162 VSUBS 0.01578f
C221 B.n163 VSUBS 0.016386f
C222 B.n164 VSUBS 0.016386f
C223 B.n165 VSUBS 0.006835f
C224 B.n166 VSUBS 0.006835f
C225 B.n167 VSUBS 0.006835f
C226 B.n168 VSUBS 0.006835f
C227 B.n169 VSUBS 0.006835f
C228 B.n170 VSUBS 0.006835f
C229 B.n171 VSUBS 0.006835f
C230 B.n172 VSUBS 0.006835f
C231 B.n173 VSUBS 0.006835f
C232 B.n174 VSUBS 0.006835f
C233 B.n175 VSUBS 0.006835f
C234 B.n176 VSUBS 0.006835f
C235 B.n177 VSUBS 0.006835f
C236 B.n178 VSUBS 0.006835f
C237 B.n179 VSUBS 0.006835f
C238 B.n180 VSUBS 0.006835f
C239 B.n181 VSUBS 0.006835f
C240 B.n182 VSUBS 0.006835f
C241 B.n183 VSUBS 0.006835f
C242 B.n184 VSUBS 0.006835f
C243 B.n185 VSUBS 0.006835f
C244 B.n186 VSUBS 0.006835f
C245 B.n187 VSUBS 0.006835f
C246 B.n188 VSUBS 0.006835f
C247 B.n189 VSUBS 0.006835f
C248 B.n190 VSUBS 0.006835f
C249 B.n191 VSUBS 0.006835f
C250 B.n192 VSUBS 0.006835f
C251 B.n193 VSUBS 0.006835f
C252 B.n194 VSUBS 0.006835f
C253 B.n195 VSUBS 0.006835f
C254 B.n196 VSUBS 0.006835f
C255 B.n197 VSUBS 0.006835f
C256 B.n198 VSUBS 0.006835f
C257 B.n199 VSUBS 0.006835f
C258 B.n200 VSUBS 0.006835f
C259 B.n201 VSUBS 0.006835f
C260 B.n202 VSUBS 0.006835f
C261 B.n203 VSUBS 0.006835f
C262 B.n204 VSUBS 0.006835f
C263 B.n205 VSUBS 0.006835f
C264 B.n206 VSUBS 0.006835f
C265 B.n207 VSUBS 0.006835f
C266 B.n208 VSUBS 0.006835f
C267 B.n209 VSUBS 0.006835f
C268 B.n210 VSUBS 0.006835f
C269 B.n211 VSUBS 0.006835f
C270 B.n212 VSUBS 0.006835f
C271 B.n213 VSUBS 0.006835f
C272 B.n214 VSUBS 0.006835f
C273 B.n215 VSUBS 0.006835f
C274 B.n216 VSUBS 0.006835f
C275 B.n217 VSUBS 0.006835f
C276 B.n218 VSUBS 0.004724f
C277 B.n219 VSUBS 0.015836f
C278 B.n220 VSUBS 0.005528f
C279 B.n221 VSUBS 0.006835f
C280 B.n222 VSUBS 0.006835f
C281 B.n223 VSUBS 0.006835f
C282 B.n224 VSUBS 0.006835f
C283 B.n225 VSUBS 0.006835f
C284 B.n226 VSUBS 0.006835f
C285 B.n227 VSUBS 0.006835f
C286 B.n228 VSUBS 0.006835f
C287 B.n229 VSUBS 0.006835f
C288 B.n230 VSUBS 0.006835f
C289 B.n231 VSUBS 0.006835f
C290 B.n232 VSUBS 0.005528f
C291 B.n233 VSUBS 0.015836f
C292 B.n234 VSUBS 0.004724f
C293 B.n235 VSUBS 0.006835f
C294 B.n236 VSUBS 0.006835f
C295 B.n237 VSUBS 0.006835f
C296 B.n238 VSUBS 0.006835f
C297 B.n239 VSUBS 0.006835f
C298 B.n240 VSUBS 0.006835f
C299 B.n241 VSUBS 0.006835f
C300 B.n242 VSUBS 0.006835f
C301 B.n243 VSUBS 0.006835f
C302 B.n244 VSUBS 0.006835f
C303 B.n245 VSUBS 0.006835f
C304 B.n246 VSUBS 0.006835f
C305 B.n247 VSUBS 0.006835f
C306 B.n248 VSUBS 0.006835f
C307 B.n249 VSUBS 0.006835f
C308 B.n250 VSUBS 0.006835f
C309 B.n251 VSUBS 0.006835f
C310 B.n252 VSUBS 0.006835f
C311 B.n253 VSUBS 0.006835f
C312 B.n254 VSUBS 0.006835f
C313 B.n255 VSUBS 0.006835f
C314 B.n256 VSUBS 0.006835f
C315 B.n257 VSUBS 0.006835f
C316 B.n258 VSUBS 0.006835f
C317 B.n259 VSUBS 0.006835f
C318 B.n260 VSUBS 0.006835f
C319 B.n261 VSUBS 0.006835f
C320 B.n262 VSUBS 0.006835f
C321 B.n263 VSUBS 0.006835f
C322 B.n264 VSUBS 0.006835f
C323 B.n265 VSUBS 0.006835f
C324 B.n266 VSUBS 0.006835f
C325 B.n267 VSUBS 0.006835f
C326 B.n268 VSUBS 0.006835f
C327 B.n269 VSUBS 0.006835f
C328 B.n270 VSUBS 0.006835f
C329 B.n271 VSUBS 0.006835f
C330 B.n272 VSUBS 0.006835f
C331 B.n273 VSUBS 0.006835f
C332 B.n274 VSUBS 0.006835f
C333 B.n275 VSUBS 0.006835f
C334 B.n276 VSUBS 0.006835f
C335 B.n277 VSUBS 0.006835f
C336 B.n278 VSUBS 0.006835f
C337 B.n279 VSUBS 0.006835f
C338 B.n280 VSUBS 0.006835f
C339 B.n281 VSUBS 0.006835f
C340 B.n282 VSUBS 0.006835f
C341 B.n283 VSUBS 0.006835f
C342 B.n284 VSUBS 0.006835f
C343 B.n285 VSUBS 0.006835f
C344 B.n286 VSUBS 0.006835f
C345 B.n287 VSUBS 0.006835f
C346 B.n288 VSUBS 0.015585f
C347 B.n289 VSUBS 0.016386f
C348 B.n290 VSUBS 0.01578f
C349 B.n291 VSUBS 0.006835f
C350 B.n292 VSUBS 0.006835f
C351 B.n293 VSUBS 0.006835f
C352 B.n294 VSUBS 0.006835f
C353 B.n295 VSUBS 0.006835f
C354 B.n296 VSUBS 0.006835f
C355 B.n297 VSUBS 0.006835f
C356 B.n298 VSUBS 0.006835f
C357 B.n299 VSUBS 0.006835f
C358 B.n300 VSUBS 0.006835f
C359 B.n301 VSUBS 0.006835f
C360 B.n302 VSUBS 0.006835f
C361 B.n303 VSUBS 0.006835f
C362 B.n304 VSUBS 0.006835f
C363 B.n305 VSUBS 0.006835f
C364 B.n306 VSUBS 0.006835f
C365 B.n307 VSUBS 0.006835f
C366 B.n308 VSUBS 0.006835f
C367 B.n309 VSUBS 0.006835f
C368 B.n310 VSUBS 0.006835f
C369 B.n311 VSUBS 0.006835f
C370 B.n312 VSUBS 0.006835f
C371 B.n313 VSUBS 0.006835f
C372 B.n314 VSUBS 0.006835f
C373 B.n315 VSUBS 0.006835f
C374 B.n316 VSUBS 0.006835f
C375 B.n317 VSUBS 0.006835f
C376 B.n318 VSUBS 0.006835f
C377 B.n319 VSUBS 0.006835f
C378 B.n320 VSUBS 0.006835f
C379 B.n321 VSUBS 0.006835f
C380 B.n322 VSUBS 0.006835f
C381 B.n323 VSUBS 0.006835f
C382 B.n324 VSUBS 0.006835f
C383 B.n325 VSUBS 0.006835f
C384 B.n326 VSUBS 0.006835f
C385 B.n327 VSUBS 0.006835f
C386 B.n328 VSUBS 0.006835f
C387 B.n329 VSUBS 0.006835f
C388 B.n330 VSUBS 0.006835f
C389 B.n331 VSUBS 0.006835f
C390 B.n332 VSUBS 0.006835f
C391 B.n333 VSUBS 0.006835f
C392 B.n334 VSUBS 0.006835f
C393 B.n335 VSUBS 0.006835f
C394 B.n336 VSUBS 0.006835f
C395 B.n337 VSUBS 0.006835f
C396 B.n338 VSUBS 0.006835f
C397 B.n339 VSUBS 0.006835f
C398 B.n340 VSUBS 0.006835f
C399 B.n341 VSUBS 0.006835f
C400 B.n342 VSUBS 0.006835f
C401 B.n343 VSUBS 0.006835f
C402 B.n344 VSUBS 0.006835f
C403 B.n345 VSUBS 0.006835f
C404 B.n346 VSUBS 0.006835f
C405 B.n347 VSUBS 0.006835f
C406 B.n348 VSUBS 0.006835f
C407 B.n349 VSUBS 0.006835f
C408 B.n350 VSUBS 0.006835f
C409 B.n351 VSUBS 0.01578f
C410 B.n352 VSUBS 0.01578f
C411 B.n353 VSUBS 0.016386f
C412 B.n354 VSUBS 0.006835f
C413 B.n355 VSUBS 0.006835f
C414 B.n356 VSUBS 0.006835f
C415 B.n357 VSUBS 0.006835f
C416 B.n358 VSUBS 0.006835f
C417 B.n359 VSUBS 0.006835f
C418 B.n360 VSUBS 0.006835f
C419 B.n361 VSUBS 0.006835f
C420 B.n362 VSUBS 0.006835f
C421 B.n363 VSUBS 0.006835f
C422 B.n364 VSUBS 0.006835f
C423 B.n365 VSUBS 0.006835f
C424 B.n366 VSUBS 0.006835f
C425 B.n367 VSUBS 0.006835f
C426 B.n368 VSUBS 0.006835f
C427 B.n369 VSUBS 0.006835f
C428 B.n370 VSUBS 0.006835f
C429 B.n371 VSUBS 0.006835f
C430 B.n372 VSUBS 0.006835f
C431 B.n373 VSUBS 0.006835f
C432 B.n374 VSUBS 0.006835f
C433 B.n375 VSUBS 0.006835f
C434 B.n376 VSUBS 0.006835f
C435 B.n377 VSUBS 0.006835f
C436 B.n378 VSUBS 0.006835f
C437 B.n379 VSUBS 0.006835f
C438 B.n380 VSUBS 0.006835f
C439 B.n381 VSUBS 0.006835f
C440 B.n382 VSUBS 0.006835f
C441 B.n383 VSUBS 0.006835f
C442 B.n384 VSUBS 0.006835f
C443 B.n385 VSUBS 0.006835f
C444 B.n386 VSUBS 0.006835f
C445 B.n387 VSUBS 0.006835f
C446 B.n388 VSUBS 0.006835f
C447 B.n389 VSUBS 0.006835f
C448 B.n390 VSUBS 0.006835f
C449 B.n391 VSUBS 0.006835f
C450 B.n392 VSUBS 0.006835f
C451 B.n393 VSUBS 0.006835f
C452 B.n394 VSUBS 0.006835f
C453 B.n395 VSUBS 0.006835f
C454 B.n396 VSUBS 0.006835f
C455 B.n397 VSUBS 0.006835f
C456 B.n398 VSUBS 0.006835f
C457 B.n399 VSUBS 0.006835f
C458 B.n400 VSUBS 0.006835f
C459 B.n401 VSUBS 0.006835f
C460 B.n402 VSUBS 0.006835f
C461 B.n403 VSUBS 0.006835f
C462 B.n404 VSUBS 0.006835f
C463 B.n405 VSUBS 0.006835f
C464 B.n406 VSUBS 0.006835f
C465 B.n407 VSUBS 0.004724f
C466 B.n408 VSUBS 0.015836f
C467 B.n409 VSUBS 0.005528f
C468 B.n410 VSUBS 0.006835f
C469 B.n411 VSUBS 0.006835f
C470 B.n412 VSUBS 0.006835f
C471 B.n413 VSUBS 0.006835f
C472 B.n414 VSUBS 0.006835f
C473 B.n415 VSUBS 0.006835f
C474 B.n416 VSUBS 0.006835f
C475 B.n417 VSUBS 0.006835f
C476 B.n418 VSUBS 0.006835f
C477 B.n419 VSUBS 0.006835f
C478 B.n420 VSUBS 0.006835f
C479 B.n421 VSUBS 0.005528f
C480 B.n422 VSUBS 0.006835f
C481 B.n423 VSUBS 0.006835f
C482 B.n424 VSUBS 0.006835f
C483 B.n425 VSUBS 0.006835f
C484 B.n426 VSUBS 0.006835f
C485 B.n427 VSUBS 0.006835f
C486 B.n428 VSUBS 0.006835f
C487 B.n429 VSUBS 0.006835f
C488 B.n430 VSUBS 0.006835f
C489 B.n431 VSUBS 0.006835f
C490 B.n432 VSUBS 0.006835f
C491 B.n433 VSUBS 0.006835f
C492 B.n434 VSUBS 0.006835f
C493 B.n435 VSUBS 0.006835f
C494 B.n436 VSUBS 0.006835f
C495 B.n437 VSUBS 0.006835f
C496 B.n438 VSUBS 0.006835f
C497 B.n439 VSUBS 0.006835f
C498 B.n440 VSUBS 0.006835f
C499 B.n441 VSUBS 0.006835f
C500 B.n442 VSUBS 0.006835f
C501 B.n443 VSUBS 0.006835f
C502 B.n444 VSUBS 0.006835f
C503 B.n445 VSUBS 0.006835f
C504 B.n446 VSUBS 0.006835f
C505 B.n447 VSUBS 0.006835f
C506 B.n448 VSUBS 0.006835f
C507 B.n449 VSUBS 0.006835f
C508 B.n450 VSUBS 0.006835f
C509 B.n451 VSUBS 0.006835f
C510 B.n452 VSUBS 0.006835f
C511 B.n453 VSUBS 0.006835f
C512 B.n454 VSUBS 0.006835f
C513 B.n455 VSUBS 0.006835f
C514 B.n456 VSUBS 0.006835f
C515 B.n457 VSUBS 0.006835f
C516 B.n458 VSUBS 0.006835f
C517 B.n459 VSUBS 0.006835f
C518 B.n460 VSUBS 0.006835f
C519 B.n461 VSUBS 0.006835f
C520 B.n462 VSUBS 0.006835f
C521 B.n463 VSUBS 0.006835f
C522 B.n464 VSUBS 0.006835f
C523 B.n465 VSUBS 0.006835f
C524 B.n466 VSUBS 0.006835f
C525 B.n467 VSUBS 0.006835f
C526 B.n468 VSUBS 0.006835f
C527 B.n469 VSUBS 0.006835f
C528 B.n470 VSUBS 0.006835f
C529 B.n471 VSUBS 0.006835f
C530 B.n472 VSUBS 0.006835f
C531 B.n473 VSUBS 0.006835f
C532 B.n474 VSUBS 0.006835f
C533 B.n475 VSUBS 0.006835f
C534 B.n476 VSUBS 0.006835f
C535 B.n477 VSUBS 0.016386f
C536 B.n478 VSUBS 0.01578f
C537 B.n479 VSUBS 0.01578f
C538 B.n480 VSUBS 0.006835f
C539 B.n481 VSUBS 0.006835f
C540 B.n482 VSUBS 0.006835f
C541 B.n483 VSUBS 0.006835f
C542 B.n484 VSUBS 0.006835f
C543 B.n485 VSUBS 0.006835f
C544 B.n486 VSUBS 0.006835f
C545 B.n487 VSUBS 0.006835f
C546 B.n488 VSUBS 0.006835f
C547 B.n489 VSUBS 0.006835f
C548 B.n490 VSUBS 0.006835f
C549 B.n491 VSUBS 0.006835f
C550 B.n492 VSUBS 0.006835f
C551 B.n493 VSUBS 0.006835f
C552 B.n494 VSUBS 0.006835f
C553 B.n495 VSUBS 0.006835f
C554 B.n496 VSUBS 0.006835f
C555 B.n497 VSUBS 0.006835f
C556 B.n498 VSUBS 0.006835f
C557 B.n499 VSUBS 0.006835f
C558 B.n500 VSUBS 0.006835f
C559 B.n501 VSUBS 0.006835f
C560 B.n502 VSUBS 0.006835f
C561 B.n503 VSUBS 0.006835f
C562 B.n504 VSUBS 0.006835f
C563 B.n505 VSUBS 0.006835f
C564 B.n506 VSUBS 0.006835f
C565 B.n507 VSUBS 0.00892f
C566 B.n508 VSUBS 0.009502f
C567 B.n509 VSUBS 0.018895f
.ends

