* NGSPICE file created from diff_pair_sample_1226.ext - technology: sky130A

.subckt diff_pair_sample_1226 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t15 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=0.72
X1 B.t11 B.t9 B.t10 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=0.72
X2 VDD2.t8 VN.t1 VTAIL.t16 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X3 VTAIL.t2 VP.t0 VDD1.t9 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X4 B.t8 B.t6 B.t7 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=0.72
X5 VTAIL.t13 VN.t2 VDD2.t7 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X6 VDD2.t6 VN.t3 VTAIL.t7 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=0.72
X7 VDD1.t8 VP.t1 VTAIL.t18 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X8 VTAIL.t5 VP.t2 VDD1.t7 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X9 VTAIL.t0 VP.t3 VDD1.t6 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X10 VDD2.t5 VN.t4 VTAIL.t14 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=0.72
X11 VDD1.t5 VP.t4 VTAIL.t19 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=0.72
X12 B.t5 B.t3 B.t4 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=0.72
X13 VDD1.t4 VP.t5 VTAIL.t1 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=1.7355 ps=9.68 w=4.45 l=0.72
X14 VTAIL.t8 VN.t5 VDD2.t4 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X15 VDD2.t3 VN.t6 VTAIL.t10 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=0.72
X16 VTAIL.t12 VN.t7 VDD2.t2 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X17 VDD1.t3 VP.t6 VTAIL.t3 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=0.72
X18 B.t2 B.t0 B.t1 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0 ps=0 w=4.45 l=0.72
X19 VDD1.t2 VP.t7 VTAIL.t17 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X20 VDD2.t1 VN.t8 VTAIL.t9 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X21 VTAIL.t6 VP.t8 VDD1.t1 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X22 VTAIL.t11 VN.t9 VDD2.t0 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=0.73425 pd=4.78 as=0.73425 ps=4.78 w=4.45 l=0.72
X23 VDD1.t0 VP.t9 VTAIL.t4 w_n2230_n1858# sky130_fd_pr__pfet_01v8 ad=1.7355 pd=9.68 as=0.73425 ps=4.78 w=4.45 l=0.72
R0 VN.n3 VN.t6 227.692
R1 VN.n17 VN.t4 227.692
R2 VN.n4 VN.t2 203.846
R3 VN.n6 VN.t1 203.846
R4 VN.n10 VN.t7 203.846
R5 VN.n12 VN.t3 203.846
R6 VN.n18 VN.t5 203.846
R7 VN.n20 VN.t8 203.846
R8 VN.n24 VN.t9 203.846
R9 VN.n26 VN.t0 203.846
R10 VN.n13 VN.n12 161.3
R11 VN.n27 VN.n26 161.3
R12 VN.n25 VN.n14 161.3
R13 VN.n24 VN.n23 161.3
R14 VN.n22 VN.n15 161.3
R15 VN.n21 VN.n20 161.3
R16 VN.n19 VN.n16 161.3
R17 VN.n11 VN.n0 161.3
R18 VN.n10 VN.n9 161.3
R19 VN.n8 VN.n1 161.3
R20 VN.n7 VN.n6 161.3
R21 VN.n5 VN.n2 161.3
R22 VN.n17 VN.n16 44.9119
R23 VN.n3 VN.n2 44.9119
R24 VN VN.n27 37.5895
R25 VN.n12 VN.n11 35.055
R26 VN.n26 VN.n25 35.055
R27 VN.n5 VN.n4 27.752
R28 VN.n10 VN.n1 27.752
R29 VN.n19 VN.n18 27.752
R30 VN.n24 VN.n15 27.752
R31 VN.n6 VN.n5 20.449
R32 VN.n6 VN.n1 20.449
R33 VN.n20 VN.n19 20.449
R34 VN.n20 VN.n15 20.449
R35 VN.n4 VN.n3 17.739
R36 VN.n18 VN.n17 17.739
R37 VN.n11 VN.n10 13.146
R38 VN.n25 VN.n24 13.146
R39 VN.n27 VN.n14 0.189894
R40 VN.n23 VN.n14 0.189894
R41 VN.n23 VN.n22 0.189894
R42 VN.n22 VN.n21 0.189894
R43 VN.n21 VN.n16 0.189894
R44 VN.n7 VN.n2 0.189894
R45 VN.n8 VN.n7 0.189894
R46 VN.n9 VN.n8 0.189894
R47 VN.n9 VN.n0 0.189894
R48 VN.n13 VN.n0 0.189894
R49 VN VN.n13 0.0516364
R50 VTAIL.n104 VTAIL.n86 756.745
R51 VTAIL.n20 VTAIL.n2 756.745
R52 VTAIL.n80 VTAIL.n62 756.745
R53 VTAIL.n52 VTAIL.n34 756.745
R54 VTAIL.n95 VTAIL.n94 585
R55 VTAIL.n97 VTAIL.n96 585
R56 VTAIL.n90 VTAIL.n89 585
R57 VTAIL.n103 VTAIL.n102 585
R58 VTAIL.n105 VTAIL.n104 585
R59 VTAIL.n11 VTAIL.n10 585
R60 VTAIL.n13 VTAIL.n12 585
R61 VTAIL.n6 VTAIL.n5 585
R62 VTAIL.n19 VTAIL.n18 585
R63 VTAIL.n21 VTAIL.n20 585
R64 VTAIL.n81 VTAIL.n80 585
R65 VTAIL.n79 VTAIL.n78 585
R66 VTAIL.n66 VTAIL.n65 585
R67 VTAIL.n73 VTAIL.n72 585
R68 VTAIL.n71 VTAIL.n70 585
R69 VTAIL.n53 VTAIL.n52 585
R70 VTAIL.n51 VTAIL.n50 585
R71 VTAIL.n38 VTAIL.n37 585
R72 VTAIL.n45 VTAIL.n44 585
R73 VTAIL.n43 VTAIL.n42 585
R74 VTAIL.n93 VTAIL.t7 328.587
R75 VTAIL.n9 VTAIL.t1 328.587
R76 VTAIL.n69 VTAIL.t19 328.587
R77 VTAIL.n41 VTAIL.t14 328.587
R78 VTAIL.n96 VTAIL.n95 171.744
R79 VTAIL.n96 VTAIL.n89 171.744
R80 VTAIL.n103 VTAIL.n89 171.744
R81 VTAIL.n104 VTAIL.n103 171.744
R82 VTAIL.n12 VTAIL.n11 171.744
R83 VTAIL.n12 VTAIL.n5 171.744
R84 VTAIL.n19 VTAIL.n5 171.744
R85 VTAIL.n20 VTAIL.n19 171.744
R86 VTAIL.n80 VTAIL.n79 171.744
R87 VTAIL.n79 VTAIL.n65 171.744
R88 VTAIL.n72 VTAIL.n65 171.744
R89 VTAIL.n72 VTAIL.n71 171.744
R90 VTAIL.n52 VTAIL.n51 171.744
R91 VTAIL.n51 VTAIL.n37 171.744
R92 VTAIL.n44 VTAIL.n37 171.744
R93 VTAIL.n44 VTAIL.n43 171.744
R94 VTAIL.n95 VTAIL.t7 85.8723
R95 VTAIL.n11 VTAIL.t1 85.8723
R96 VTAIL.n71 VTAIL.t19 85.8723
R97 VTAIL.n43 VTAIL.t14 85.8723
R98 VTAIL.n61 VTAIL.n60 85.2677
R99 VTAIL.n59 VTAIL.n58 85.2677
R100 VTAIL.n33 VTAIL.n32 85.2677
R101 VTAIL.n31 VTAIL.n30 85.2677
R102 VTAIL.n111 VTAIL.n110 85.2675
R103 VTAIL.n1 VTAIL.n0 85.2675
R104 VTAIL.n27 VTAIL.n26 85.2675
R105 VTAIL.n29 VTAIL.n28 85.2675
R106 VTAIL.n109 VTAIL.n108 30.052
R107 VTAIL.n25 VTAIL.n24 30.052
R108 VTAIL.n85 VTAIL.n84 30.052
R109 VTAIL.n57 VTAIL.n56 30.052
R110 VTAIL.n31 VTAIL.n29 18.0134
R111 VTAIL.n109 VTAIL.n85 17.1083
R112 VTAIL.n94 VTAIL.n93 16.3651
R113 VTAIL.n10 VTAIL.n9 16.3651
R114 VTAIL.n70 VTAIL.n69 16.3651
R115 VTAIL.n42 VTAIL.n41 16.3651
R116 VTAIL.n97 VTAIL.n92 12.8005
R117 VTAIL.n13 VTAIL.n8 12.8005
R118 VTAIL.n73 VTAIL.n68 12.8005
R119 VTAIL.n45 VTAIL.n40 12.8005
R120 VTAIL.n98 VTAIL.n90 12.0247
R121 VTAIL.n14 VTAIL.n6 12.0247
R122 VTAIL.n74 VTAIL.n66 12.0247
R123 VTAIL.n46 VTAIL.n38 12.0247
R124 VTAIL.n102 VTAIL.n101 11.249
R125 VTAIL.n18 VTAIL.n17 11.249
R126 VTAIL.n78 VTAIL.n77 11.249
R127 VTAIL.n50 VTAIL.n49 11.249
R128 VTAIL.n105 VTAIL.n88 10.4732
R129 VTAIL.n21 VTAIL.n4 10.4732
R130 VTAIL.n81 VTAIL.n64 10.4732
R131 VTAIL.n53 VTAIL.n36 10.4732
R132 VTAIL.n106 VTAIL.n86 9.69747
R133 VTAIL.n22 VTAIL.n2 9.69747
R134 VTAIL.n82 VTAIL.n62 9.69747
R135 VTAIL.n54 VTAIL.n34 9.69747
R136 VTAIL.n108 VTAIL.n107 9.45567
R137 VTAIL.n24 VTAIL.n23 9.45567
R138 VTAIL.n84 VTAIL.n83 9.45567
R139 VTAIL.n56 VTAIL.n55 9.45567
R140 VTAIL.n107 VTAIL.n106 9.3005
R141 VTAIL.n88 VTAIL.n87 9.3005
R142 VTAIL.n101 VTAIL.n100 9.3005
R143 VTAIL.n99 VTAIL.n98 9.3005
R144 VTAIL.n92 VTAIL.n91 9.3005
R145 VTAIL.n23 VTAIL.n22 9.3005
R146 VTAIL.n4 VTAIL.n3 9.3005
R147 VTAIL.n17 VTAIL.n16 9.3005
R148 VTAIL.n15 VTAIL.n14 9.3005
R149 VTAIL.n8 VTAIL.n7 9.3005
R150 VTAIL.n83 VTAIL.n82 9.3005
R151 VTAIL.n64 VTAIL.n63 9.3005
R152 VTAIL.n77 VTAIL.n76 9.3005
R153 VTAIL.n75 VTAIL.n74 9.3005
R154 VTAIL.n68 VTAIL.n67 9.3005
R155 VTAIL.n55 VTAIL.n54 9.3005
R156 VTAIL.n36 VTAIL.n35 9.3005
R157 VTAIL.n49 VTAIL.n48 9.3005
R158 VTAIL.n47 VTAIL.n46 9.3005
R159 VTAIL.n40 VTAIL.n39 9.3005
R160 VTAIL.n110 VTAIL.t16 7.30499
R161 VTAIL.n110 VTAIL.t12 7.30499
R162 VTAIL.n0 VTAIL.t10 7.30499
R163 VTAIL.n0 VTAIL.t13 7.30499
R164 VTAIL.n26 VTAIL.t17 7.30499
R165 VTAIL.n26 VTAIL.t2 7.30499
R166 VTAIL.n28 VTAIL.t4 7.30499
R167 VTAIL.n28 VTAIL.t5 7.30499
R168 VTAIL.n60 VTAIL.t18 7.30499
R169 VTAIL.n60 VTAIL.t0 7.30499
R170 VTAIL.n58 VTAIL.t3 7.30499
R171 VTAIL.n58 VTAIL.t6 7.30499
R172 VTAIL.n32 VTAIL.t9 7.30499
R173 VTAIL.n32 VTAIL.t8 7.30499
R174 VTAIL.n30 VTAIL.t15 7.30499
R175 VTAIL.n30 VTAIL.t11 7.30499
R176 VTAIL.n108 VTAIL.n86 4.26717
R177 VTAIL.n24 VTAIL.n2 4.26717
R178 VTAIL.n84 VTAIL.n62 4.26717
R179 VTAIL.n56 VTAIL.n34 4.26717
R180 VTAIL.n93 VTAIL.n91 3.73474
R181 VTAIL.n9 VTAIL.n7 3.73474
R182 VTAIL.n69 VTAIL.n67 3.73474
R183 VTAIL.n41 VTAIL.n39 3.73474
R184 VTAIL.n106 VTAIL.n105 3.49141
R185 VTAIL.n22 VTAIL.n21 3.49141
R186 VTAIL.n82 VTAIL.n81 3.49141
R187 VTAIL.n54 VTAIL.n53 3.49141
R188 VTAIL.n102 VTAIL.n88 2.71565
R189 VTAIL.n18 VTAIL.n4 2.71565
R190 VTAIL.n78 VTAIL.n64 2.71565
R191 VTAIL.n50 VTAIL.n36 2.71565
R192 VTAIL.n101 VTAIL.n90 1.93989
R193 VTAIL.n17 VTAIL.n6 1.93989
R194 VTAIL.n77 VTAIL.n66 1.93989
R195 VTAIL.n49 VTAIL.n38 1.93989
R196 VTAIL.n98 VTAIL.n97 1.16414
R197 VTAIL.n14 VTAIL.n13 1.16414
R198 VTAIL.n74 VTAIL.n73 1.16414
R199 VTAIL.n46 VTAIL.n45 1.16414
R200 VTAIL.n59 VTAIL.n57 0.922914
R201 VTAIL.n25 VTAIL.n1 0.922914
R202 VTAIL.n33 VTAIL.n31 0.905672
R203 VTAIL.n57 VTAIL.n33 0.905672
R204 VTAIL.n61 VTAIL.n59 0.905672
R205 VTAIL.n85 VTAIL.n61 0.905672
R206 VTAIL.n29 VTAIL.n27 0.905672
R207 VTAIL.n27 VTAIL.n25 0.905672
R208 VTAIL.n111 VTAIL.n109 0.905672
R209 VTAIL VTAIL.n1 0.737569
R210 VTAIL.n94 VTAIL.n92 0.388379
R211 VTAIL.n10 VTAIL.n8 0.388379
R212 VTAIL.n70 VTAIL.n68 0.388379
R213 VTAIL.n42 VTAIL.n40 0.388379
R214 VTAIL VTAIL.n111 0.168603
R215 VTAIL.n99 VTAIL.n91 0.155672
R216 VTAIL.n100 VTAIL.n99 0.155672
R217 VTAIL.n100 VTAIL.n87 0.155672
R218 VTAIL.n107 VTAIL.n87 0.155672
R219 VTAIL.n15 VTAIL.n7 0.155672
R220 VTAIL.n16 VTAIL.n15 0.155672
R221 VTAIL.n16 VTAIL.n3 0.155672
R222 VTAIL.n23 VTAIL.n3 0.155672
R223 VTAIL.n83 VTAIL.n63 0.155672
R224 VTAIL.n76 VTAIL.n63 0.155672
R225 VTAIL.n76 VTAIL.n75 0.155672
R226 VTAIL.n75 VTAIL.n67 0.155672
R227 VTAIL.n55 VTAIL.n35 0.155672
R228 VTAIL.n48 VTAIL.n35 0.155672
R229 VTAIL.n48 VTAIL.n47 0.155672
R230 VTAIL.n47 VTAIL.n39 0.155672
R231 VDD2.n45 VDD2.n27 756.745
R232 VDD2.n18 VDD2.n0 756.745
R233 VDD2.n46 VDD2.n45 585
R234 VDD2.n44 VDD2.n43 585
R235 VDD2.n31 VDD2.n30 585
R236 VDD2.n38 VDD2.n37 585
R237 VDD2.n36 VDD2.n35 585
R238 VDD2.n9 VDD2.n8 585
R239 VDD2.n11 VDD2.n10 585
R240 VDD2.n4 VDD2.n3 585
R241 VDD2.n17 VDD2.n16 585
R242 VDD2.n19 VDD2.n18 585
R243 VDD2.n34 VDD2.t9 328.587
R244 VDD2.n7 VDD2.t3 328.587
R245 VDD2.n45 VDD2.n44 171.744
R246 VDD2.n44 VDD2.n30 171.744
R247 VDD2.n37 VDD2.n30 171.744
R248 VDD2.n37 VDD2.n36 171.744
R249 VDD2.n10 VDD2.n9 171.744
R250 VDD2.n10 VDD2.n3 171.744
R251 VDD2.n17 VDD2.n3 171.744
R252 VDD2.n18 VDD2.n17 171.744
R253 VDD2.n26 VDD2.n25 102.57
R254 VDD2 VDD2.n53 102.567
R255 VDD2.n52 VDD2.n51 101.947
R256 VDD2.n24 VDD2.n23 101.947
R257 VDD2.n36 VDD2.t9 85.8723
R258 VDD2.n9 VDD2.t3 85.8723
R259 VDD2.n24 VDD2.n22 47.636
R260 VDD2.n50 VDD2.n49 46.7308
R261 VDD2.n50 VDD2.n26 31.8511
R262 VDD2.n35 VDD2.n34 16.3651
R263 VDD2.n8 VDD2.n7 16.3651
R264 VDD2.n38 VDD2.n33 12.8005
R265 VDD2.n11 VDD2.n6 12.8005
R266 VDD2.n39 VDD2.n31 12.0247
R267 VDD2.n12 VDD2.n4 12.0247
R268 VDD2.n43 VDD2.n42 11.249
R269 VDD2.n16 VDD2.n15 11.249
R270 VDD2.n46 VDD2.n29 10.4732
R271 VDD2.n19 VDD2.n2 10.4732
R272 VDD2.n47 VDD2.n27 9.69747
R273 VDD2.n20 VDD2.n0 9.69747
R274 VDD2.n49 VDD2.n48 9.45567
R275 VDD2.n22 VDD2.n21 9.45567
R276 VDD2.n48 VDD2.n47 9.3005
R277 VDD2.n29 VDD2.n28 9.3005
R278 VDD2.n42 VDD2.n41 9.3005
R279 VDD2.n40 VDD2.n39 9.3005
R280 VDD2.n33 VDD2.n32 9.3005
R281 VDD2.n21 VDD2.n20 9.3005
R282 VDD2.n2 VDD2.n1 9.3005
R283 VDD2.n15 VDD2.n14 9.3005
R284 VDD2.n13 VDD2.n12 9.3005
R285 VDD2.n6 VDD2.n5 9.3005
R286 VDD2.n53 VDD2.t4 7.30499
R287 VDD2.n53 VDD2.t5 7.30499
R288 VDD2.n51 VDD2.t0 7.30499
R289 VDD2.n51 VDD2.t1 7.30499
R290 VDD2.n25 VDD2.t2 7.30499
R291 VDD2.n25 VDD2.t6 7.30499
R292 VDD2.n23 VDD2.t7 7.30499
R293 VDD2.n23 VDD2.t8 7.30499
R294 VDD2.n49 VDD2.n27 4.26717
R295 VDD2.n22 VDD2.n0 4.26717
R296 VDD2.n34 VDD2.n32 3.73474
R297 VDD2.n7 VDD2.n5 3.73474
R298 VDD2.n47 VDD2.n46 3.49141
R299 VDD2.n20 VDD2.n19 3.49141
R300 VDD2.n43 VDD2.n29 2.71565
R301 VDD2.n16 VDD2.n2 2.71565
R302 VDD2.n42 VDD2.n31 1.93989
R303 VDD2.n15 VDD2.n4 1.93989
R304 VDD2.n39 VDD2.n38 1.16414
R305 VDD2.n12 VDD2.n11 1.16414
R306 VDD2.n52 VDD2.n50 0.905672
R307 VDD2.n35 VDD2.n33 0.388379
R308 VDD2.n8 VDD2.n6 0.388379
R309 VDD2 VDD2.n52 0.284983
R310 VDD2.n26 VDD2.n24 0.171447
R311 VDD2.n48 VDD2.n28 0.155672
R312 VDD2.n41 VDD2.n28 0.155672
R313 VDD2.n41 VDD2.n40 0.155672
R314 VDD2.n40 VDD2.n32 0.155672
R315 VDD2.n13 VDD2.n5 0.155672
R316 VDD2.n14 VDD2.n13 0.155672
R317 VDD2.n14 VDD2.n1 0.155672
R318 VDD2.n21 VDD2.n1 0.155672
R319 B.n222 B.n71 585
R320 B.n221 B.n220 585
R321 B.n219 B.n72 585
R322 B.n218 B.n217 585
R323 B.n216 B.n73 585
R324 B.n215 B.n214 585
R325 B.n213 B.n74 585
R326 B.n212 B.n211 585
R327 B.n210 B.n75 585
R328 B.n209 B.n208 585
R329 B.n207 B.n76 585
R330 B.n206 B.n205 585
R331 B.n204 B.n77 585
R332 B.n203 B.n202 585
R333 B.n201 B.n78 585
R334 B.n200 B.n199 585
R335 B.n198 B.n79 585
R336 B.n197 B.n196 585
R337 B.n195 B.n80 585
R338 B.n193 B.n192 585
R339 B.n191 B.n83 585
R340 B.n190 B.n189 585
R341 B.n188 B.n84 585
R342 B.n187 B.n186 585
R343 B.n185 B.n85 585
R344 B.n184 B.n183 585
R345 B.n182 B.n86 585
R346 B.n181 B.n180 585
R347 B.n179 B.n87 585
R348 B.n178 B.n177 585
R349 B.n173 B.n88 585
R350 B.n172 B.n171 585
R351 B.n170 B.n89 585
R352 B.n169 B.n168 585
R353 B.n167 B.n90 585
R354 B.n166 B.n165 585
R355 B.n164 B.n91 585
R356 B.n163 B.n162 585
R357 B.n161 B.n92 585
R358 B.n160 B.n159 585
R359 B.n158 B.n93 585
R360 B.n157 B.n156 585
R361 B.n155 B.n94 585
R362 B.n154 B.n153 585
R363 B.n152 B.n95 585
R364 B.n151 B.n150 585
R365 B.n149 B.n96 585
R366 B.n148 B.n147 585
R367 B.n224 B.n223 585
R368 B.n225 B.n70 585
R369 B.n227 B.n226 585
R370 B.n228 B.n69 585
R371 B.n230 B.n229 585
R372 B.n231 B.n68 585
R373 B.n233 B.n232 585
R374 B.n234 B.n67 585
R375 B.n236 B.n235 585
R376 B.n237 B.n66 585
R377 B.n239 B.n238 585
R378 B.n240 B.n65 585
R379 B.n242 B.n241 585
R380 B.n243 B.n64 585
R381 B.n245 B.n244 585
R382 B.n246 B.n63 585
R383 B.n248 B.n247 585
R384 B.n249 B.n62 585
R385 B.n251 B.n250 585
R386 B.n252 B.n61 585
R387 B.n254 B.n253 585
R388 B.n255 B.n60 585
R389 B.n257 B.n256 585
R390 B.n258 B.n59 585
R391 B.n260 B.n259 585
R392 B.n261 B.n58 585
R393 B.n263 B.n262 585
R394 B.n264 B.n57 585
R395 B.n266 B.n265 585
R396 B.n267 B.n56 585
R397 B.n269 B.n268 585
R398 B.n270 B.n55 585
R399 B.n272 B.n271 585
R400 B.n273 B.n54 585
R401 B.n275 B.n274 585
R402 B.n276 B.n53 585
R403 B.n278 B.n277 585
R404 B.n279 B.n52 585
R405 B.n281 B.n280 585
R406 B.n282 B.n51 585
R407 B.n284 B.n283 585
R408 B.n285 B.n50 585
R409 B.n287 B.n286 585
R410 B.n288 B.n49 585
R411 B.n290 B.n289 585
R412 B.n291 B.n48 585
R413 B.n293 B.n292 585
R414 B.n294 B.n47 585
R415 B.n296 B.n295 585
R416 B.n297 B.n46 585
R417 B.n299 B.n298 585
R418 B.n300 B.n45 585
R419 B.n302 B.n301 585
R420 B.n303 B.n44 585
R421 B.n376 B.n15 585
R422 B.n375 B.n374 585
R423 B.n373 B.n16 585
R424 B.n372 B.n371 585
R425 B.n370 B.n17 585
R426 B.n369 B.n368 585
R427 B.n367 B.n18 585
R428 B.n366 B.n365 585
R429 B.n364 B.n19 585
R430 B.n363 B.n362 585
R431 B.n361 B.n20 585
R432 B.n360 B.n359 585
R433 B.n358 B.n21 585
R434 B.n357 B.n356 585
R435 B.n355 B.n22 585
R436 B.n354 B.n353 585
R437 B.n352 B.n23 585
R438 B.n351 B.n350 585
R439 B.n349 B.n24 585
R440 B.n348 B.n347 585
R441 B.n346 B.n25 585
R442 B.n345 B.n344 585
R443 B.n343 B.n29 585
R444 B.n342 B.n341 585
R445 B.n340 B.n30 585
R446 B.n339 B.n338 585
R447 B.n337 B.n31 585
R448 B.n336 B.n335 585
R449 B.n334 B.n32 585
R450 B.n332 B.n331 585
R451 B.n330 B.n35 585
R452 B.n329 B.n328 585
R453 B.n327 B.n36 585
R454 B.n326 B.n325 585
R455 B.n324 B.n37 585
R456 B.n323 B.n322 585
R457 B.n321 B.n38 585
R458 B.n320 B.n319 585
R459 B.n318 B.n39 585
R460 B.n317 B.n316 585
R461 B.n315 B.n40 585
R462 B.n314 B.n313 585
R463 B.n312 B.n41 585
R464 B.n311 B.n310 585
R465 B.n309 B.n42 585
R466 B.n308 B.n307 585
R467 B.n306 B.n43 585
R468 B.n305 B.n304 585
R469 B.n378 B.n377 585
R470 B.n379 B.n14 585
R471 B.n381 B.n380 585
R472 B.n382 B.n13 585
R473 B.n384 B.n383 585
R474 B.n385 B.n12 585
R475 B.n387 B.n386 585
R476 B.n388 B.n11 585
R477 B.n390 B.n389 585
R478 B.n391 B.n10 585
R479 B.n393 B.n392 585
R480 B.n394 B.n9 585
R481 B.n396 B.n395 585
R482 B.n397 B.n8 585
R483 B.n399 B.n398 585
R484 B.n400 B.n7 585
R485 B.n402 B.n401 585
R486 B.n403 B.n6 585
R487 B.n405 B.n404 585
R488 B.n406 B.n5 585
R489 B.n408 B.n407 585
R490 B.n409 B.n4 585
R491 B.n411 B.n410 585
R492 B.n412 B.n3 585
R493 B.n414 B.n413 585
R494 B.n415 B.n0 585
R495 B.n2 B.n1 585
R496 B.n110 B.n109 585
R497 B.n112 B.n111 585
R498 B.n113 B.n108 585
R499 B.n115 B.n114 585
R500 B.n116 B.n107 585
R501 B.n118 B.n117 585
R502 B.n119 B.n106 585
R503 B.n121 B.n120 585
R504 B.n122 B.n105 585
R505 B.n124 B.n123 585
R506 B.n125 B.n104 585
R507 B.n127 B.n126 585
R508 B.n128 B.n103 585
R509 B.n130 B.n129 585
R510 B.n131 B.n102 585
R511 B.n133 B.n132 585
R512 B.n134 B.n101 585
R513 B.n136 B.n135 585
R514 B.n137 B.n100 585
R515 B.n139 B.n138 585
R516 B.n140 B.n99 585
R517 B.n142 B.n141 585
R518 B.n143 B.n98 585
R519 B.n145 B.n144 585
R520 B.n146 B.n97 585
R521 B.n147 B.n146 554.963
R522 B.n223 B.n222 554.963
R523 B.n305 B.n44 554.963
R524 B.n378 B.n15 554.963
R525 B.n174 B.t6 351.678
R526 B.n81 B.t0 351.678
R527 B.n33 B.t3 351.678
R528 B.n26 B.t9 351.678
R529 B.n81 B.t1 261.8
R530 B.n33 B.t5 261.8
R531 B.n174 B.t7 261.8
R532 B.n26 B.t11 261.8
R533 B.n417 B.n416 256.663
R534 B.n82 B.t2 241.435
R535 B.n34 B.t4 241.435
R536 B.n175 B.t8 241.435
R537 B.n27 B.t10 241.435
R538 B.n416 B.n415 235.042
R539 B.n416 B.n2 235.042
R540 B.n147 B.n96 163.367
R541 B.n151 B.n96 163.367
R542 B.n152 B.n151 163.367
R543 B.n153 B.n152 163.367
R544 B.n153 B.n94 163.367
R545 B.n157 B.n94 163.367
R546 B.n158 B.n157 163.367
R547 B.n159 B.n158 163.367
R548 B.n159 B.n92 163.367
R549 B.n163 B.n92 163.367
R550 B.n164 B.n163 163.367
R551 B.n165 B.n164 163.367
R552 B.n165 B.n90 163.367
R553 B.n169 B.n90 163.367
R554 B.n170 B.n169 163.367
R555 B.n171 B.n170 163.367
R556 B.n171 B.n88 163.367
R557 B.n178 B.n88 163.367
R558 B.n179 B.n178 163.367
R559 B.n180 B.n179 163.367
R560 B.n180 B.n86 163.367
R561 B.n184 B.n86 163.367
R562 B.n185 B.n184 163.367
R563 B.n186 B.n185 163.367
R564 B.n186 B.n84 163.367
R565 B.n190 B.n84 163.367
R566 B.n191 B.n190 163.367
R567 B.n192 B.n191 163.367
R568 B.n192 B.n80 163.367
R569 B.n197 B.n80 163.367
R570 B.n198 B.n197 163.367
R571 B.n199 B.n198 163.367
R572 B.n199 B.n78 163.367
R573 B.n203 B.n78 163.367
R574 B.n204 B.n203 163.367
R575 B.n205 B.n204 163.367
R576 B.n205 B.n76 163.367
R577 B.n209 B.n76 163.367
R578 B.n210 B.n209 163.367
R579 B.n211 B.n210 163.367
R580 B.n211 B.n74 163.367
R581 B.n215 B.n74 163.367
R582 B.n216 B.n215 163.367
R583 B.n217 B.n216 163.367
R584 B.n217 B.n72 163.367
R585 B.n221 B.n72 163.367
R586 B.n222 B.n221 163.367
R587 B.n301 B.n44 163.367
R588 B.n301 B.n300 163.367
R589 B.n300 B.n299 163.367
R590 B.n299 B.n46 163.367
R591 B.n295 B.n46 163.367
R592 B.n295 B.n294 163.367
R593 B.n294 B.n293 163.367
R594 B.n293 B.n48 163.367
R595 B.n289 B.n48 163.367
R596 B.n289 B.n288 163.367
R597 B.n288 B.n287 163.367
R598 B.n287 B.n50 163.367
R599 B.n283 B.n50 163.367
R600 B.n283 B.n282 163.367
R601 B.n282 B.n281 163.367
R602 B.n281 B.n52 163.367
R603 B.n277 B.n52 163.367
R604 B.n277 B.n276 163.367
R605 B.n276 B.n275 163.367
R606 B.n275 B.n54 163.367
R607 B.n271 B.n54 163.367
R608 B.n271 B.n270 163.367
R609 B.n270 B.n269 163.367
R610 B.n269 B.n56 163.367
R611 B.n265 B.n56 163.367
R612 B.n265 B.n264 163.367
R613 B.n264 B.n263 163.367
R614 B.n263 B.n58 163.367
R615 B.n259 B.n58 163.367
R616 B.n259 B.n258 163.367
R617 B.n258 B.n257 163.367
R618 B.n257 B.n60 163.367
R619 B.n253 B.n60 163.367
R620 B.n253 B.n252 163.367
R621 B.n252 B.n251 163.367
R622 B.n251 B.n62 163.367
R623 B.n247 B.n62 163.367
R624 B.n247 B.n246 163.367
R625 B.n246 B.n245 163.367
R626 B.n245 B.n64 163.367
R627 B.n241 B.n64 163.367
R628 B.n241 B.n240 163.367
R629 B.n240 B.n239 163.367
R630 B.n239 B.n66 163.367
R631 B.n235 B.n66 163.367
R632 B.n235 B.n234 163.367
R633 B.n234 B.n233 163.367
R634 B.n233 B.n68 163.367
R635 B.n229 B.n68 163.367
R636 B.n229 B.n228 163.367
R637 B.n228 B.n227 163.367
R638 B.n227 B.n70 163.367
R639 B.n223 B.n70 163.367
R640 B.n374 B.n15 163.367
R641 B.n374 B.n373 163.367
R642 B.n373 B.n372 163.367
R643 B.n372 B.n17 163.367
R644 B.n368 B.n17 163.367
R645 B.n368 B.n367 163.367
R646 B.n367 B.n366 163.367
R647 B.n366 B.n19 163.367
R648 B.n362 B.n19 163.367
R649 B.n362 B.n361 163.367
R650 B.n361 B.n360 163.367
R651 B.n360 B.n21 163.367
R652 B.n356 B.n21 163.367
R653 B.n356 B.n355 163.367
R654 B.n355 B.n354 163.367
R655 B.n354 B.n23 163.367
R656 B.n350 B.n23 163.367
R657 B.n350 B.n349 163.367
R658 B.n349 B.n348 163.367
R659 B.n348 B.n25 163.367
R660 B.n344 B.n25 163.367
R661 B.n344 B.n343 163.367
R662 B.n343 B.n342 163.367
R663 B.n342 B.n30 163.367
R664 B.n338 B.n30 163.367
R665 B.n338 B.n337 163.367
R666 B.n337 B.n336 163.367
R667 B.n336 B.n32 163.367
R668 B.n331 B.n32 163.367
R669 B.n331 B.n330 163.367
R670 B.n330 B.n329 163.367
R671 B.n329 B.n36 163.367
R672 B.n325 B.n36 163.367
R673 B.n325 B.n324 163.367
R674 B.n324 B.n323 163.367
R675 B.n323 B.n38 163.367
R676 B.n319 B.n38 163.367
R677 B.n319 B.n318 163.367
R678 B.n318 B.n317 163.367
R679 B.n317 B.n40 163.367
R680 B.n313 B.n40 163.367
R681 B.n313 B.n312 163.367
R682 B.n312 B.n311 163.367
R683 B.n311 B.n42 163.367
R684 B.n307 B.n42 163.367
R685 B.n307 B.n306 163.367
R686 B.n306 B.n305 163.367
R687 B.n379 B.n378 163.367
R688 B.n380 B.n379 163.367
R689 B.n380 B.n13 163.367
R690 B.n384 B.n13 163.367
R691 B.n385 B.n384 163.367
R692 B.n386 B.n385 163.367
R693 B.n386 B.n11 163.367
R694 B.n390 B.n11 163.367
R695 B.n391 B.n390 163.367
R696 B.n392 B.n391 163.367
R697 B.n392 B.n9 163.367
R698 B.n396 B.n9 163.367
R699 B.n397 B.n396 163.367
R700 B.n398 B.n397 163.367
R701 B.n398 B.n7 163.367
R702 B.n402 B.n7 163.367
R703 B.n403 B.n402 163.367
R704 B.n404 B.n403 163.367
R705 B.n404 B.n5 163.367
R706 B.n408 B.n5 163.367
R707 B.n409 B.n408 163.367
R708 B.n410 B.n409 163.367
R709 B.n410 B.n3 163.367
R710 B.n414 B.n3 163.367
R711 B.n415 B.n414 163.367
R712 B.n110 B.n2 163.367
R713 B.n111 B.n110 163.367
R714 B.n111 B.n108 163.367
R715 B.n115 B.n108 163.367
R716 B.n116 B.n115 163.367
R717 B.n117 B.n116 163.367
R718 B.n117 B.n106 163.367
R719 B.n121 B.n106 163.367
R720 B.n122 B.n121 163.367
R721 B.n123 B.n122 163.367
R722 B.n123 B.n104 163.367
R723 B.n127 B.n104 163.367
R724 B.n128 B.n127 163.367
R725 B.n129 B.n128 163.367
R726 B.n129 B.n102 163.367
R727 B.n133 B.n102 163.367
R728 B.n134 B.n133 163.367
R729 B.n135 B.n134 163.367
R730 B.n135 B.n100 163.367
R731 B.n139 B.n100 163.367
R732 B.n140 B.n139 163.367
R733 B.n141 B.n140 163.367
R734 B.n141 B.n98 163.367
R735 B.n145 B.n98 163.367
R736 B.n146 B.n145 163.367
R737 B.n176 B.n175 59.5399
R738 B.n194 B.n82 59.5399
R739 B.n333 B.n34 59.5399
R740 B.n28 B.n27 59.5399
R741 B.n377 B.n376 36.059
R742 B.n304 B.n303 36.059
R743 B.n148 B.n97 36.059
R744 B.n224 B.n71 36.059
R745 B.n175 B.n174 20.3641
R746 B.n82 B.n81 20.3641
R747 B.n34 B.n33 20.3641
R748 B.n27 B.n26 20.3641
R749 B B.n417 18.0485
R750 B.n377 B.n14 10.6151
R751 B.n381 B.n14 10.6151
R752 B.n382 B.n381 10.6151
R753 B.n383 B.n382 10.6151
R754 B.n383 B.n12 10.6151
R755 B.n387 B.n12 10.6151
R756 B.n388 B.n387 10.6151
R757 B.n389 B.n388 10.6151
R758 B.n389 B.n10 10.6151
R759 B.n393 B.n10 10.6151
R760 B.n394 B.n393 10.6151
R761 B.n395 B.n394 10.6151
R762 B.n395 B.n8 10.6151
R763 B.n399 B.n8 10.6151
R764 B.n400 B.n399 10.6151
R765 B.n401 B.n400 10.6151
R766 B.n401 B.n6 10.6151
R767 B.n405 B.n6 10.6151
R768 B.n406 B.n405 10.6151
R769 B.n407 B.n406 10.6151
R770 B.n407 B.n4 10.6151
R771 B.n411 B.n4 10.6151
R772 B.n412 B.n411 10.6151
R773 B.n413 B.n412 10.6151
R774 B.n413 B.n0 10.6151
R775 B.n376 B.n375 10.6151
R776 B.n375 B.n16 10.6151
R777 B.n371 B.n16 10.6151
R778 B.n371 B.n370 10.6151
R779 B.n370 B.n369 10.6151
R780 B.n369 B.n18 10.6151
R781 B.n365 B.n18 10.6151
R782 B.n365 B.n364 10.6151
R783 B.n364 B.n363 10.6151
R784 B.n363 B.n20 10.6151
R785 B.n359 B.n20 10.6151
R786 B.n359 B.n358 10.6151
R787 B.n358 B.n357 10.6151
R788 B.n357 B.n22 10.6151
R789 B.n353 B.n22 10.6151
R790 B.n353 B.n352 10.6151
R791 B.n352 B.n351 10.6151
R792 B.n351 B.n24 10.6151
R793 B.n347 B.n346 10.6151
R794 B.n346 B.n345 10.6151
R795 B.n345 B.n29 10.6151
R796 B.n341 B.n29 10.6151
R797 B.n341 B.n340 10.6151
R798 B.n340 B.n339 10.6151
R799 B.n339 B.n31 10.6151
R800 B.n335 B.n31 10.6151
R801 B.n335 B.n334 10.6151
R802 B.n332 B.n35 10.6151
R803 B.n328 B.n35 10.6151
R804 B.n328 B.n327 10.6151
R805 B.n327 B.n326 10.6151
R806 B.n326 B.n37 10.6151
R807 B.n322 B.n37 10.6151
R808 B.n322 B.n321 10.6151
R809 B.n321 B.n320 10.6151
R810 B.n320 B.n39 10.6151
R811 B.n316 B.n39 10.6151
R812 B.n316 B.n315 10.6151
R813 B.n315 B.n314 10.6151
R814 B.n314 B.n41 10.6151
R815 B.n310 B.n41 10.6151
R816 B.n310 B.n309 10.6151
R817 B.n309 B.n308 10.6151
R818 B.n308 B.n43 10.6151
R819 B.n304 B.n43 10.6151
R820 B.n303 B.n302 10.6151
R821 B.n302 B.n45 10.6151
R822 B.n298 B.n45 10.6151
R823 B.n298 B.n297 10.6151
R824 B.n297 B.n296 10.6151
R825 B.n296 B.n47 10.6151
R826 B.n292 B.n47 10.6151
R827 B.n292 B.n291 10.6151
R828 B.n291 B.n290 10.6151
R829 B.n290 B.n49 10.6151
R830 B.n286 B.n49 10.6151
R831 B.n286 B.n285 10.6151
R832 B.n285 B.n284 10.6151
R833 B.n284 B.n51 10.6151
R834 B.n280 B.n51 10.6151
R835 B.n280 B.n279 10.6151
R836 B.n279 B.n278 10.6151
R837 B.n278 B.n53 10.6151
R838 B.n274 B.n53 10.6151
R839 B.n274 B.n273 10.6151
R840 B.n273 B.n272 10.6151
R841 B.n272 B.n55 10.6151
R842 B.n268 B.n55 10.6151
R843 B.n268 B.n267 10.6151
R844 B.n267 B.n266 10.6151
R845 B.n266 B.n57 10.6151
R846 B.n262 B.n57 10.6151
R847 B.n262 B.n261 10.6151
R848 B.n261 B.n260 10.6151
R849 B.n260 B.n59 10.6151
R850 B.n256 B.n59 10.6151
R851 B.n256 B.n255 10.6151
R852 B.n255 B.n254 10.6151
R853 B.n254 B.n61 10.6151
R854 B.n250 B.n61 10.6151
R855 B.n250 B.n249 10.6151
R856 B.n249 B.n248 10.6151
R857 B.n248 B.n63 10.6151
R858 B.n244 B.n63 10.6151
R859 B.n244 B.n243 10.6151
R860 B.n243 B.n242 10.6151
R861 B.n242 B.n65 10.6151
R862 B.n238 B.n65 10.6151
R863 B.n238 B.n237 10.6151
R864 B.n237 B.n236 10.6151
R865 B.n236 B.n67 10.6151
R866 B.n232 B.n67 10.6151
R867 B.n232 B.n231 10.6151
R868 B.n231 B.n230 10.6151
R869 B.n230 B.n69 10.6151
R870 B.n226 B.n69 10.6151
R871 B.n226 B.n225 10.6151
R872 B.n225 B.n224 10.6151
R873 B.n109 B.n1 10.6151
R874 B.n112 B.n109 10.6151
R875 B.n113 B.n112 10.6151
R876 B.n114 B.n113 10.6151
R877 B.n114 B.n107 10.6151
R878 B.n118 B.n107 10.6151
R879 B.n119 B.n118 10.6151
R880 B.n120 B.n119 10.6151
R881 B.n120 B.n105 10.6151
R882 B.n124 B.n105 10.6151
R883 B.n125 B.n124 10.6151
R884 B.n126 B.n125 10.6151
R885 B.n126 B.n103 10.6151
R886 B.n130 B.n103 10.6151
R887 B.n131 B.n130 10.6151
R888 B.n132 B.n131 10.6151
R889 B.n132 B.n101 10.6151
R890 B.n136 B.n101 10.6151
R891 B.n137 B.n136 10.6151
R892 B.n138 B.n137 10.6151
R893 B.n138 B.n99 10.6151
R894 B.n142 B.n99 10.6151
R895 B.n143 B.n142 10.6151
R896 B.n144 B.n143 10.6151
R897 B.n144 B.n97 10.6151
R898 B.n149 B.n148 10.6151
R899 B.n150 B.n149 10.6151
R900 B.n150 B.n95 10.6151
R901 B.n154 B.n95 10.6151
R902 B.n155 B.n154 10.6151
R903 B.n156 B.n155 10.6151
R904 B.n156 B.n93 10.6151
R905 B.n160 B.n93 10.6151
R906 B.n161 B.n160 10.6151
R907 B.n162 B.n161 10.6151
R908 B.n162 B.n91 10.6151
R909 B.n166 B.n91 10.6151
R910 B.n167 B.n166 10.6151
R911 B.n168 B.n167 10.6151
R912 B.n168 B.n89 10.6151
R913 B.n172 B.n89 10.6151
R914 B.n173 B.n172 10.6151
R915 B.n177 B.n173 10.6151
R916 B.n181 B.n87 10.6151
R917 B.n182 B.n181 10.6151
R918 B.n183 B.n182 10.6151
R919 B.n183 B.n85 10.6151
R920 B.n187 B.n85 10.6151
R921 B.n188 B.n187 10.6151
R922 B.n189 B.n188 10.6151
R923 B.n189 B.n83 10.6151
R924 B.n193 B.n83 10.6151
R925 B.n196 B.n195 10.6151
R926 B.n196 B.n79 10.6151
R927 B.n200 B.n79 10.6151
R928 B.n201 B.n200 10.6151
R929 B.n202 B.n201 10.6151
R930 B.n202 B.n77 10.6151
R931 B.n206 B.n77 10.6151
R932 B.n207 B.n206 10.6151
R933 B.n208 B.n207 10.6151
R934 B.n208 B.n75 10.6151
R935 B.n212 B.n75 10.6151
R936 B.n213 B.n212 10.6151
R937 B.n214 B.n213 10.6151
R938 B.n214 B.n73 10.6151
R939 B.n218 B.n73 10.6151
R940 B.n219 B.n218 10.6151
R941 B.n220 B.n219 10.6151
R942 B.n220 B.n71 10.6151
R943 B.n28 B.n24 9.36635
R944 B.n333 B.n332 9.36635
R945 B.n177 B.n176 9.36635
R946 B.n195 B.n194 9.36635
R947 B.n417 B.n0 8.11757
R948 B.n417 B.n1 8.11757
R949 B.n347 B.n28 1.24928
R950 B.n334 B.n333 1.24928
R951 B.n176 B.n87 1.24928
R952 B.n194 B.n193 1.24928
R953 VP.n7 VP.t6 227.692
R954 VP.n18 VP.t9 203.846
R955 VP.n22 VP.t2 203.846
R956 VP.n24 VP.t7 203.846
R957 VP.n28 VP.t0 203.846
R958 VP.n30 VP.t5 203.846
R959 VP.n16 VP.t4 203.846
R960 VP.n14 VP.t3 203.846
R961 VP.n6 VP.t1 203.846
R962 VP.n8 VP.t8 203.846
R963 VP.n31 VP.n30 161.3
R964 VP.n10 VP.n9 161.3
R965 VP.n11 VP.n6 161.3
R966 VP.n13 VP.n12 161.3
R967 VP.n14 VP.n5 161.3
R968 VP.n15 VP.n4 161.3
R969 VP.n17 VP.n16 161.3
R970 VP.n29 VP.n0 161.3
R971 VP.n28 VP.n27 161.3
R972 VP.n26 VP.n1 161.3
R973 VP.n25 VP.n24 161.3
R974 VP.n23 VP.n2 161.3
R975 VP.n22 VP.n21 161.3
R976 VP.n20 VP.n3 161.3
R977 VP.n19 VP.n18 161.3
R978 VP.n10 VP.n7 44.9119
R979 VP.n19 VP.n17 37.2088
R980 VP.n18 VP.n3 35.055
R981 VP.n30 VP.n29 35.055
R982 VP.n16 VP.n15 35.055
R983 VP.n23 VP.n22 27.752
R984 VP.n28 VP.n1 27.752
R985 VP.n14 VP.n13 27.752
R986 VP.n9 VP.n8 27.752
R987 VP.n24 VP.n23 20.449
R988 VP.n24 VP.n1 20.449
R989 VP.n13 VP.n6 20.449
R990 VP.n9 VP.n6 20.449
R991 VP.n8 VP.n7 17.739
R992 VP.n22 VP.n3 13.146
R993 VP.n29 VP.n28 13.146
R994 VP.n15 VP.n14 13.146
R995 VP.n11 VP.n10 0.189894
R996 VP.n12 VP.n11 0.189894
R997 VP.n12 VP.n5 0.189894
R998 VP.n5 VP.n4 0.189894
R999 VP.n17 VP.n4 0.189894
R1000 VP.n20 VP.n19 0.189894
R1001 VP.n21 VP.n20 0.189894
R1002 VP.n21 VP.n2 0.189894
R1003 VP.n25 VP.n2 0.189894
R1004 VP.n26 VP.n25 0.189894
R1005 VP.n27 VP.n26 0.189894
R1006 VP.n27 VP.n0 0.189894
R1007 VP.n31 VP.n0 0.189894
R1008 VP VP.n31 0.0516364
R1009 VDD1.n18 VDD1.n0 756.745
R1010 VDD1.n43 VDD1.n25 756.745
R1011 VDD1.n19 VDD1.n18 585
R1012 VDD1.n17 VDD1.n16 585
R1013 VDD1.n4 VDD1.n3 585
R1014 VDD1.n11 VDD1.n10 585
R1015 VDD1.n9 VDD1.n8 585
R1016 VDD1.n34 VDD1.n33 585
R1017 VDD1.n36 VDD1.n35 585
R1018 VDD1.n29 VDD1.n28 585
R1019 VDD1.n42 VDD1.n41 585
R1020 VDD1.n44 VDD1.n43 585
R1021 VDD1.n7 VDD1.t3 328.587
R1022 VDD1.n32 VDD1.t0 328.587
R1023 VDD1.n18 VDD1.n17 171.744
R1024 VDD1.n17 VDD1.n3 171.744
R1025 VDD1.n10 VDD1.n3 171.744
R1026 VDD1.n10 VDD1.n9 171.744
R1027 VDD1.n35 VDD1.n34 171.744
R1028 VDD1.n35 VDD1.n28 171.744
R1029 VDD1.n42 VDD1.n28 171.744
R1030 VDD1.n43 VDD1.n42 171.744
R1031 VDD1.n51 VDD1.n50 102.57
R1032 VDD1.n24 VDD1.n23 101.947
R1033 VDD1.n53 VDD1.n52 101.947
R1034 VDD1.n49 VDD1.n48 101.947
R1035 VDD1.n9 VDD1.t3 85.8723
R1036 VDD1.n34 VDD1.t0 85.8723
R1037 VDD1.n24 VDD1.n22 47.636
R1038 VDD1.n49 VDD1.n47 47.636
R1039 VDD1.n53 VDD1.n51 32.8867
R1040 VDD1.n8 VDD1.n7 16.3651
R1041 VDD1.n33 VDD1.n32 16.3651
R1042 VDD1.n11 VDD1.n6 12.8005
R1043 VDD1.n36 VDD1.n31 12.8005
R1044 VDD1.n12 VDD1.n4 12.0247
R1045 VDD1.n37 VDD1.n29 12.0247
R1046 VDD1.n16 VDD1.n15 11.249
R1047 VDD1.n41 VDD1.n40 11.249
R1048 VDD1.n19 VDD1.n2 10.4732
R1049 VDD1.n44 VDD1.n27 10.4732
R1050 VDD1.n20 VDD1.n0 9.69747
R1051 VDD1.n45 VDD1.n25 9.69747
R1052 VDD1.n22 VDD1.n21 9.45567
R1053 VDD1.n47 VDD1.n46 9.45567
R1054 VDD1.n21 VDD1.n20 9.3005
R1055 VDD1.n2 VDD1.n1 9.3005
R1056 VDD1.n15 VDD1.n14 9.3005
R1057 VDD1.n13 VDD1.n12 9.3005
R1058 VDD1.n6 VDD1.n5 9.3005
R1059 VDD1.n46 VDD1.n45 9.3005
R1060 VDD1.n27 VDD1.n26 9.3005
R1061 VDD1.n40 VDD1.n39 9.3005
R1062 VDD1.n38 VDD1.n37 9.3005
R1063 VDD1.n31 VDD1.n30 9.3005
R1064 VDD1.n52 VDD1.t6 7.30499
R1065 VDD1.n52 VDD1.t5 7.30499
R1066 VDD1.n23 VDD1.t1 7.30499
R1067 VDD1.n23 VDD1.t8 7.30499
R1068 VDD1.n50 VDD1.t9 7.30499
R1069 VDD1.n50 VDD1.t4 7.30499
R1070 VDD1.n48 VDD1.t7 7.30499
R1071 VDD1.n48 VDD1.t2 7.30499
R1072 VDD1.n22 VDD1.n0 4.26717
R1073 VDD1.n47 VDD1.n25 4.26717
R1074 VDD1.n7 VDD1.n5 3.73474
R1075 VDD1.n32 VDD1.n30 3.73474
R1076 VDD1.n20 VDD1.n19 3.49141
R1077 VDD1.n45 VDD1.n44 3.49141
R1078 VDD1.n16 VDD1.n2 2.71565
R1079 VDD1.n41 VDD1.n27 2.71565
R1080 VDD1.n15 VDD1.n4 1.93989
R1081 VDD1.n40 VDD1.n29 1.93989
R1082 VDD1.n12 VDD1.n11 1.16414
R1083 VDD1.n37 VDD1.n36 1.16414
R1084 VDD1 VDD1.n53 0.62119
R1085 VDD1.n8 VDD1.n6 0.388379
R1086 VDD1.n33 VDD1.n31 0.388379
R1087 VDD1 VDD1.n24 0.284983
R1088 VDD1.n51 VDD1.n49 0.171447
R1089 VDD1.n21 VDD1.n1 0.155672
R1090 VDD1.n14 VDD1.n1 0.155672
R1091 VDD1.n14 VDD1.n13 0.155672
R1092 VDD1.n13 VDD1.n5 0.155672
R1093 VDD1.n38 VDD1.n30 0.155672
R1094 VDD1.n39 VDD1.n38 0.155672
R1095 VDD1.n39 VDD1.n26 0.155672
R1096 VDD1.n46 VDD1.n26 0.155672
C0 VP VDD2 0.347096f
C1 VDD1 VN 0.152836f
C2 B VN 0.721511f
C3 VDD1 VDD2 0.980841f
C4 B VDD2 1.20675f
C5 VTAIL VN 3.02234f
C6 VDD1 VP 2.98969f
C7 w_n2230_n1858# VN 4.05588f
C8 VP B 1.18948f
C9 VTAIL VDD2 6.84551f
C10 w_n2230_n1858# VDD2 1.53274f
C11 VP VTAIL 3.03663f
C12 VDD1 B 1.16165f
C13 VP w_n2230_n1858# 4.34012f
C14 VDD1 VTAIL 6.80696f
C15 VDD1 w_n2230_n1858# 1.48743f
C16 VTAIL B 1.38234f
C17 VDD2 VN 2.79788f
C18 w_n2230_n1858# B 5.27112f
C19 VP VN 4.23308f
C20 w_n2230_n1858# VTAIL 1.82184f
C21 VDD2 VSUBS 1.060054f
C22 VDD1 VSUBS 0.91824f
C23 VTAIL VSUBS 0.396475f
C24 VN VSUBS 4.4181f
C25 VP VSUBS 1.442347f
C26 B VSUBS 2.291213f
C27 w_n2230_n1858# VSUBS 52.0482f
C28 VDD1.n0 VSUBS 0.025f
C29 VDD1.n1 VSUBS 0.024653f
C30 VDD1.n2 VSUBS 0.013248f
C31 VDD1.n3 VSUBS 0.031313f
C32 VDD1.n4 VSUBS 0.014027f
C33 VDD1.n5 VSUBS 0.39143f
C34 VDD1.n6 VSUBS 0.013248f
C35 VDD1.t3 VSUBS 0.067567f
C36 VDD1.n7 VSUBS 0.097957f
C37 VDD1.n8 VSUBS 0.019837f
C38 VDD1.n9 VSUBS 0.023484f
C39 VDD1.n10 VSUBS 0.031313f
C40 VDD1.n11 VSUBS 0.014027f
C41 VDD1.n12 VSUBS 0.013248f
C42 VDD1.n13 VSUBS 0.024653f
C43 VDD1.n14 VSUBS 0.024653f
C44 VDD1.n15 VSUBS 0.013248f
C45 VDD1.n16 VSUBS 0.014027f
C46 VDD1.n17 VSUBS 0.031313f
C47 VDD1.n18 VSUBS 0.06869f
C48 VDD1.n19 VSUBS 0.014027f
C49 VDD1.n20 VSUBS 0.013248f
C50 VDD1.n21 VSUBS 0.05328f
C51 VDD1.n22 VSUBS 0.053393f
C52 VDD1.t1 VSUBS 0.086694f
C53 VDD1.t8 VSUBS 0.086694f
C54 VDD1.n23 VSUBS 0.523806f
C55 VDD1.n24 VSUBS 0.573367f
C56 VDD1.n25 VSUBS 0.025f
C57 VDD1.n26 VSUBS 0.024653f
C58 VDD1.n27 VSUBS 0.013248f
C59 VDD1.n28 VSUBS 0.031313f
C60 VDD1.n29 VSUBS 0.014027f
C61 VDD1.n30 VSUBS 0.39143f
C62 VDD1.n31 VSUBS 0.013248f
C63 VDD1.t0 VSUBS 0.067567f
C64 VDD1.n32 VSUBS 0.097957f
C65 VDD1.n33 VSUBS 0.019837f
C66 VDD1.n34 VSUBS 0.023484f
C67 VDD1.n35 VSUBS 0.031313f
C68 VDD1.n36 VSUBS 0.014027f
C69 VDD1.n37 VSUBS 0.013248f
C70 VDD1.n38 VSUBS 0.024653f
C71 VDD1.n39 VSUBS 0.024653f
C72 VDD1.n40 VSUBS 0.013248f
C73 VDD1.n41 VSUBS 0.014027f
C74 VDD1.n42 VSUBS 0.031313f
C75 VDD1.n43 VSUBS 0.06869f
C76 VDD1.n44 VSUBS 0.014027f
C77 VDD1.n45 VSUBS 0.013248f
C78 VDD1.n46 VSUBS 0.05328f
C79 VDD1.n47 VSUBS 0.053393f
C80 VDD1.t7 VSUBS 0.086694f
C81 VDD1.t2 VSUBS 0.086694f
C82 VDD1.n48 VSUBS 0.523804f
C83 VDD1.n49 VSUBS 0.567694f
C84 VDD1.t9 VSUBS 0.086694f
C85 VDD1.t4 VSUBS 0.086694f
C86 VDD1.n50 VSUBS 0.52682f
C87 VDD1.n51 VSUBS 1.68167f
C88 VDD1.t6 VSUBS 0.086694f
C89 VDD1.t5 VSUBS 0.086694f
C90 VDD1.n52 VSUBS 0.523804f
C91 VDD1.n53 VSUBS 1.93181f
C92 VP.n0 VSUBS 0.063735f
C93 VP.n1 VSUBS 0.014463f
C94 VP.n2 VSUBS 0.063735f
C95 VP.n3 VSUBS 0.014463f
C96 VP.n4 VSUBS 0.063735f
C97 VP.t4 VSUBS 0.59972f
C98 VP.t3 VSUBS 0.59972f
C99 VP.n5 VSUBS 0.063735f
C100 VP.t1 VSUBS 0.59972f
C101 VP.n6 VSUBS 0.301855f
C102 VP.t6 VSUBS 0.631424f
C103 VP.n7 VSUBS 0.27649f
C104 VP.t8 VSUBS 0.59972f
C105 VP.n8 VSUBS 0.30975f
C106 VP.n9 VSUBS 0.014463f
C107 VP.n10 VSUBS 0.270103f
C108 VP.n11 VSUBS 0.063735f
C109 VP.n12 VSUBS 0.063735f
C110 VP.n13 VSUBS 0.014463f
C111 VP.n14 VSUBS 0.301855f
C112 VP.n15 VSUBS 0.014463f
C113 VP.n16 VSUBS 0.300284f
C114 VP.n17 VSUBS 2.13024f
C115 VP.t9 VSUBS 0.59972f
C116 VP.n18 VSUBS 0.300284f
C117 VP.n19 VSUBS 2.19182f
C118 VP.n20 VSUBS 0.063735f
C119 VP.n21 VSUBS 0.063735f
C120 VP.t2 VSUBS 0.59972f
C121 VP.n22 VSUBS 0.301855f
C122 VP.n23 VSUBS 0.014463f
C123 VP.t7 VSUBS 0.59972f
C124 VP.n24 VSUBS 0.301855f
C125 VP.n25 VSUBS 0.063735f
C126 VP.n26 VSUBS 0.063735f
C127 VP.n27 VSUBS 0.063735f
C128 VP.t0 VSUBS 0.59972f
C129 VP.n28 VSUBS 0.301855f
C130 VP.n29 VSUBS 0.014463f
C131 VP.t5 VSUBS 0.59972f
C132 VP.n30 VSUBS 0.300284f
C133 VP.n31 VSUBS 0.049392f
C134 B.n0 VSUBS 0.00629f
C135 B.n1 VSUBS 0.00629f
C136 B.n2 VSUBS 0.009302f
C137 B.n3 VSUBS 0.007128f
C138 B.n4 VSUBS 0.007128f
C139 B.n5 VSUBS 0.007128f
C140 B.n6 VSUBS 0.007128f
C141 B.n7 VSUBS 0.007128f
C142 B.n8 VSUBS 0.007128f
C143 B.n9 VSUBS 0.007128f
C144 B.n10 VSUBS 0.007128f
C145 B.n11 VSUBS 0.007128f
C146 B.n12 VSUBS 0.007128f
C147 B.n13 VSUBS 0.007128f
C148 B.n14 VSUBS 0.007128f
C149 B.n15 VSUBS 0.018147f
C150 B.n16 VSUBS 0.007128f
C151 B.n17 VSUBS 0.007128f
C152 B.n18 VSUBS 0.007128f
C153 B.n19 VSUBS 0.007128f
C154 B.n20 VSUBS 0.007128f
C155 B.n21 VSUBS 0.007128f
C156 B.n22 VSUBS 0.007128f
C157 B.n23 VSUBS 0.007128f
C158 B.n24 VSUBS 0.006709f
C159 B.n25 VSUBS 0.007128f
C160 B.t10 VSUBS 0.065039f
C161 B.t11 VSUBS 0.073614f
C162 B.t9 VSUBS 0.144876f
C163 B.n26 VSUBS 0.135051f
C164 B.n27 VSUBS 0.120402f
C165 B.n28 VSUBS 0.016516f
C166 B.n29 VSUBS 0.007128f
C167 B.n30 VSUBS 0.007128f
C168 B.n31 VSUBS 0.007128f
C169 B.n32 VSUBS 0.007128f
C170 B.t4 VSUBS 0.06504f
C171 B.t5 VSUBS 0.073615f
C172 B.t3 VSUBS 0.144876f
C173 B.n33 VSUBS 0.13505f
C174 B.n34 VSUBS 0.120401f
C175 B.n35 VSUBS 0.007128f
C176 B.n36 VSUBS 0.007128f
C177 B.n37 VSUBS 0.007128f
C178 B.n38 VSUBS 0.007128f
C179 B.n39 VSUBS 0.007128f
C180 B.n40 VSUBS 0.007128f
C181 B.n41 VSUBS 0.007128f
C182 B.n42 VSUBS 0.007128f
C183 B.n43 VSUBS 0.007128f
C184 B.n44 VSUBS 0.017495f
C185 B.n45 VSUBS 0.007128f
C186 B.n46 VSUBS 0.007128f
C187 B.n47 VSUBS 0.007128f
C188 B.n48 VSUBS 0.007128f
C189 B.n49 VSUBS 0.007128f
C190 B.n50 VSUBS 0.007128f
C191 B.n51 VSUBS 0.007128f
C192 B.n52 VSUBS 0.007128f
C193 B.n53 VSUBS 0.007128f
C194 B.n54 VSUBS 0.007128f
C195 B.n55 VSUBS 0.007128f
C196 B.n56 VSUBS 0.007128f
C197 B.n57 VSUBS 0.007128f
C198 B.n58 VSUBS 0.007128f
C199 B.n59 VSUBS 0.007128f
C200 B.n60 VSUBS 0.007128f
C201 B.n61 VSUBS 0.007128f
C202 B.n62 VSUBS 0.007128f
C203 B.n63 VSUBS 0.007128f
C204 B.n64 VSUBS 0.007128f
C205 B.n65 VSUBS 0.007128f
C206 B.n66 VSUBS 0.007128f
C207 B.n67 VSUBS 0.007128f
C208 B.n68 VSUBS 0.007128f
C209 B.n69 VSUBS 0.007128f
C210 B.n70 VSUBS 0.007128f
C211 B.n71 VSUBS 0.017384f
C212 B.n72 VSUBS 0.007128f
C213 B.n73 VSUBS 0.007128f
C214 B.n74 VSUBS 0.007128f
C215 B.n75 VSUBS 0.007128f
C216 B.n76 VSUBS 0.007128f
C217 B.n77 VSUBS 0.007128f
C218 B.n78 VSUBS 0.007128f
C219 B.n79 VSUBS 0.007128f
C220 B.n80 VSUBS 0.007128f
C221 B.t2 VSUBS 0.06504f
C222 B.t1 VSUBS 0.073615f
C223 B.t0 VSUBS 0.144876f
C224 B.n81 VSUBS 0.13505f
C225 B.n82 VSUBS 0.120401f
C226 B.n83 VSUBS 0.007128f
C227 B.n84 VSUBS 0.007128f
C228 B.n85 VSUBS 0.007128f
C229 B.n86 VSUBS 0.007128f
C230 B.n87 VSUBS 0.003984f
C231 B.n88 VSUBS 0.007128f
C232 B.n89 VSUBS 0.007128f
C233 B.n90 VSUBS 0.007128f
C234 B.n91 VSUBS 0.007128f
C235 B.n92 VSUBS 0.007128f
C236 B.n93 VSUBS 0.007128f
C237 B.n94 VSUBS 0.007128f
C238 B.n95 VSUBS 0.007128f
C239 B.n96 VSUBS 0.007128f
C240 B.n97 VSUBS 0.017495f
C241 B.n98 VSUBS 0.007128f
C242 B.n99 VSUBS 0.007128f
C243 B.n100 VSUBS 0.007128f
C244 B.n101 VSUBS 0.007128f
C245 B.n102 VSUBS 0.007128f
C246 B.n103 VSUBS 0.007128f
C247 B.n104 VSUBS 0.007128f
C248 B.n105 VSUBS 0.007128f
C249 B.n106 VSUBS 0.007128f
C250 B.n107 VSUBS 0.007128f
C251 B.n108 VSUBS 0.007128f
C252 B.n109 VSUBS 0.007128f
C253 B.n110 VSUBS 0.007128f
C254 B.n111 VSUBS 0.007128f
C255 B.n112 VSUBS 0.007128f
C256 B.n113 VSUBS 0.007128f
C257 B.n114 VSUBS 0.007128f
C258 B.n115 VSUBS 0.007128f
C259 B.n116 VSUBS 0.007128f
C260 B.n117 VSUBS 0.007128f
C261 B.n118 VSUBS 0.007128f
C262 B.n119 VSUBS 0.007128f
C263 B.n120 VSUBS 0.007128f
C264 B.n121 VSUBS 0.007128f
C265 B.n122 VSUBS 0.007128f
C266 B.n123 VSUBS 0.007128f
C267 B.n124 VSUBS 0.007128f
C268 B.n125 VSUBS 0.007128f
C269 B.n126 VSUBS 0.007128f
C270 B.n127 VSUBS 0.007128f
C271 B.n128 VSUBS 0.007128f
C272 B.n129 VSUBS 0.007128f
C273 B.n130 VSUBS 0.007128f
C274 B.n131 VSUBS 0.007128f
C275 B.n132 VSUBS 0.007128f
C276 B.n133 VSUBS 0.007128f
C277 B.n134 VSUBS 0.007128f
C278 B.n135 VSUBS 0.007128f
C279 B.n136 VSUBS 0.007128f
C280 B.n137 VSUBS 0.007128f
C281 B.n138 VSUBS 0.007128f
C282 B.n139 VSUBS 0.007128f
C283 B.n140 VSUBS 0.007128f
C284 B.n141 VSUBS 0.007128f
C285 B.n142 VSUBS 0.007128f
C286 B.n143 VSUBS 0.007128f
C287 B.n144 VSUBS 0.007128f
C288 B.n145 VSUBS 0.007128f
C289 B.n146 VSUBS 0.017495f
C290 B.n147 VSUBS 0.018147f
C291 B.n148 VSUBS 0.018147f
C292 B.n149 VSUBS 0.007128f
C293 B.n150 VSUBS 0.007128f
C294 B.n151 VSUBS 0.007128f
C295 B.n152 VSUBS 0.007128f
C296 B.n153 VSUBS 0.007128f
C297 B.n154 VSUBS 0.007128f
C298 B.n155 VSUBS 0.007128f
C299 B.n156 VSUBS 0.007128f
C300 B.n157 VSUBS 0.007128f
C301 B.n158 VSUBS 0.007128f
C302 B.n159 VSUBS 0.007128f
C303 B.n160 VSUBS 0.007128f
C304 B.n161 VSUBS 0.007128f
C305 B.n162 VSUBS 0.007128f
C306 B.n163 VSUBS 0.007128f
C307 B.n164 VSUBS 0.007128f
C308 B.n165 VSUBS 0.007128f
C309 B.n166 VSUBS 0.007128f
C310 B.n167 VSUBS 0.007128f
C311 B.n168 VSUBS 0.007128f
C312 B.n169 VSUBS 0.007128f
C313 B.n170 VSUBS 0.007128f
C314 B.n171 VSUBS 0.007128f
C315 B.n172 VSUBS 0.007128f
C316 B.n173 VSUBS 0.007128f
C317 B.t8 VSUBS 0.065039f
C318 B.t7 VSUBS 0.073614f
C319 B.t6 VSUBS 0.144876f
C320 B.n174 VSUBS 0.135051f
C321 B.n175 VSUBS 0.120402f
C322 B.n176 VSUBS 0.016516f
C323 B.n177 VSUBS 0.006709f
C324 B.n178 VSUBS 0.007128f
C325 B.n179 VSUBS 0.007128f
C326 B.n180 VSUBS 0.007128f
C327 B.n181 VSUBS 0.007128f
C328 B.n182 VSUBS 0.007128f
C329 B.n183 VSUBS 0.007128f
C330 B.n184 VSUBS 0.007128f
C331 B.n185 VSUBS 0.007128f
C332 B.n186 VSUBS 0.007128f
C333 B.n187 VSUBS 0.007128f
C334 B.n188 VSUBS 0.007128f
C335 B.n189 VSUBS 0.007128f
C336 B.n190 VSUBS 0.007128f
C337 B.n191 VSUBS 0.007128f
C338 B.n192 VSUBS 0.007128f
C339 B.n193 VSUBS 0.003984f
C340 B.n194 VSUBS 0.016516f
C341 B.n195 VSUBS 0.006709f
C342 B.n196 VSUBS 0.007128f
C343 B.n197 VSUBS 0.007128f
C344 B.n198 VSUBS 0.007128f
C345 B.n199 VSUBS 0.007128f
C346 B.n200 VSUBS 0.007128f
C347 B.n201 VSUBS 0.007128f
C348 B.n202 VSUBS 0.007128f
C349 B.n203 VSUBS 0.007128f
C350 B.n204 VSUBS 0.007128f
C351 B.n205 VSUBS 0.007128f
C352 B.n206 VSUBS 0.007128f
C353 B.n207 VSUBS 0.007128f
C354 B.n208 VSUBS 0.007128f
C355 B.n209 VSUBS 0.007128f
C356 B.n210 VSUBS 0.007128f
C357 B.n211 VSUBS 0.007128f
C358 B.n212 VSUBS 0.007128f
C359 B.n213 VSUBS 0.007128f
C360 B.n214 VSUBS 0.007128f
C361 B.n215 VSUBS 0.007128f
C362 B.n216 VSUBS 0.007128f
C363 B.n217 VSUBS 0.007128f
C364 B.n218 VSUBS 0.007128f
C365 B.n219 VSUBS 0.007128f
C366 B.n220 VSUBS 0.007128f
C367 B.n221 VSUBS 0.007128f
C368 B.n222 VSUBS 0.018147f
C369 B.n223 VSUBS 0.017495f
C370 B.n224 VSUBS 0.018258f
C371 B.n225 VSUBS 0.007128f
C372 B.n226 VSUBS 0.007128f
C373 B.n227 VSUBS 0.007128f
C374 B.n228 VSUBS 0.007128f
C375 B.n229 VSUBS 0.007128f
C376 B.n230 VSUBS 0.007128f
C377 B.n231 VSUBS 0.007128f
C378 B.n232 VSUBS 0.007128f
C379 B.n233 VSUBS 0.007128f
C380 B.n234 VSUBS 0.007128f
C381 B.n235 VSUBS 0.007128f
C382 B.n236 VSUBS 0.007128f
C383 B.n237 VSUBS 0.007128f
C384 B.n238 VSUBS 0.007128f
C385 B.n239 VSUBS 0.007128f
C386 B.n240 VSUBS 0.007128f
C387 B.n241 VSUBS 0.007128f
C388 B.n242 VSUBS 0.007128f
C389 B.n243 VSUBS 0.007128f
C390 B.n244 VSUBS 0.007128f
C391 B.n245 VSUBS 0.007128f
C392 B.n246 VSUBS 0.007128f
C393 B.n247 VSUBS 0.007128f
C394 B.n248 VSUBS 0.007128f
C395 B.n249 VSUBS 0.007128f
C396 B.n250 VSUBS 0.007128f
C397 B.n251 VSUBS 0.007128f
C398 B.n252 VSUBS 0.007128f
C399 B.n253 VSUBS 0.007128f
C400 B.n254 VSUBS 0.007128f
C401 B.n255 VSUBS 0.007128f
C402 B.n256 VSUBS 0.007128f
C403 B.n257 VSUBS 0.007128f
C404 B.n258 VSUBS 0.007128f
C405 B.n259 VSUBS 0.007128f
C406 B.n260 VSUBS 0.007128f
C407 B.n261 VSUBS 0.007128f
C408 B.n262 VSUBS 0.007128f
C409 B.n263 VSUBS 0.007128f
C410 B.n264 VSUBS 0.007128f
C411 B.n265 VSUBS 0.007128f
C412 B.n266 VSUBS 0.007128f
C413 B.n267 VSUBS 0.007128f
C414 B.n268 VSUBS 0.007128f
C415 B.n269 VSUBS 0.007128f
C416 B.n270 VSUBS 0.007128f
C417 B.n271 VSUBS 0.007128f
C418 B.n272 VSUBS 0.007128f
C419 B.n273 VSUBS 0.007128f
C420 B.n274 VSUBS 0.007128f
C421 B.n275 VSUBS 0.007128f
C422 B.n276 VSUBS 0.007128f
C423 B.n277 VSUBS 0.007128f
C424 B.n278 VSUBS 0.007128f
C425 B.n279 VSUBS 0.007128f
C426 B.n280 VSUBS 0.007128f
C427 B.n281 VSUBS 0.007128f
C428 B.n282 VSUBS 0.007128f
C429 B.n283 VSUBS 0.007128f
C430 B.n284 VSUBS 0.007128f
C431 B.n285 VSUBS 0.007128f
C432 B.n286 VSUBS 0.007128f
C433 B.n287 VSUBS 0.007128f
C434 B.n288 VSUBS 0.007128f
C435 B.n289 VSUBS 0.007128f
C436 B.n290 VSUBS 0.007128f
C437 B.n291 VSUBS 0.007128f
C438 B.n292 VSUBS 0.007128f
C439 B.n293 VSUBS 0.007128f
C440 B.n294 VSUBS 0.007128f
C441 B.n295 VSUBS 0.007128f
C442 B.n296 VSUBS 0.007128f
C443 B.n297 VSUBS 0.007128f
C444 B.n298 VSUBS 0.007128f
C445 B.n299 VSUBS 0.007128f
C446 B.n300 VSUBS 0.007128f
C447 B.n301 VSUBS 0.007128f
C448 B.n302 VSUBS 0.007128f
C449 B.n303 VSUBS 0.017495f
C450 B.n304 VSUBS 0.018147f
C451 B.n305 VSUBS 0.018147f
C452 B.n306 VSUBS 0.007128f
C453 B.n307 VSUBS 0.007128f
C454 B.n308 VSUBS 0.007128f
C455 B.n309 VSUBS 0.007128f
C456 B.n310 VSUBS 0.007128f
C457 B.n311 VSUBS 0.007128f
C458 B.n312 VSUBS 0.007128f
C459 B.n313 VSUBS 0.007128f
C460 B.n314 VSUBS 0.007128f
C461 B.n315 VSUBS 0.007128f
C462 B.n316 VSUBS 0.007128f
C463 B.n317 VSUBS 0.007128f
C464 B.n318 VSUBS 0.007128f
C465 B.n319 VSUBS 0.007128f
C466 B.n320 VSUBS 0.007128f
C467 B.n321 VSUBS 0.007128f
C468 B.n322 VSUBS 0.007128f
C469 B.n323 VSUBS 0.007128f
C470 B.n324 VSUBS 0.007128f
C471 B.n325 VSUBS 0.007128f
C472 B.n326 VSUBS 0.007128f
C473 B.n327 VSUBS 0.007128f
C474 B.n328 VSUBS 0.007128f
C475 B.n329 VSUBS 0.007128f
C476 B.n330 VSUBS 0.007128f
C477 B.n331 VSUBS 0.007128f
C478 B.n332 VSUBS 0.006709f
C479 B.n333 VSUBS 0.016516f
C480 B.n334 VSUBS 0.003984f
C481 B.n335 VSUBS 0.007128f
C482 B.n336 VSUBS 0.007128f
C483 B.n337 VSUBS 0.007128f
C484 B.n338 VSUBS 0.007128f
C485 B.n339 VSUBS 0.007128f
C486 B.n340 VSUBS 0.007128f
C487 B.n341 VSUBS 0.007128f
C488 B.n342 VSUBS 0.007128f
C489 B.n343 VSUBS 0.007128f
C490 B.n344 VSUBS 0.007128f
C491 B.n345 VSUBS 0.007128f
C492 B.n346 VSUBS 0.007128f
C493 B.n347 VSUBS 0.003984f
C494 B.n348 VSUBS 0.007128f
C495 B.n349 VSUBS 0.007128f
C496 B.n350 VSUBS 0.007128f
C497 B.n351 VSUBS 0.007128f
C498 B.n352 VSUBS 0.007128f
C499 B.n353 VSUBS 0.007128f
C500 B.n354 VSUBS 0.007128f
C501 B.n355 VSUBS 0.007128f
C502 B.n356 VSUBS 0.007128f
C503 B.n357 VSUBS 0.007128f
C504 B.n358 VSUBS 0.007128f
C505 B.n359 VSUBS 0.007128f
C506 B.n360 VSUBS 0.007128f
C507 B.n361 VSUBS 0.007128f
C508 B.n362 VSUBS 0.007128f
C509 B.n363 VSUBS 0.007128f
C510 B.n364 VSUBS 0.007128f
C511 B.n365 VSUBS 0.007128f
C512 B.n366 VSUBS 0.007128f
C513 B.n367 VSUBS 0.007128f
C514 B.n368 VSUBS 0.007128f
C515 B.n369 VSUBS 0.007128f
C516 B.n370 VSUBS 0.007128f
C517 B.n371 VSUBS 0.007128f
C518 B.n372 VSUBS 0.007128f
C519 B.n373 VSUBS 0.007128f
C520 B.n374 VSUBS 0.007128f
C521 B.n375 VSUBS 0.007128f
C522 B.n376 VSUBS 0.018147f
C523 B.n377 VSUBS 0.017495f
C524 B.n378 VSUBS 0.017495f
C525 B.n379 VSUBS 0.007128f
C526 B.n380 VSUBS 0.007128f
C527 B.n381 VSUBS 0.007128f
C528 B.n382 VSUBS 0.007128f
C529 B.n383 VSUBS 0.007128f
C530 B.n384 VSUBS 0.007128f
C531 B.n385 VSUBS 0.007128f
C532 B.n386 VSUBS 0.007128f
C533 B.n387 VSUBS 0.007128f
C534 B.n388 VSUBS 0.007128f
C535 B.n389 VSUBS 0.007128f
C536 B.n390 VSUBS 0.007128f
C537 B.n391 VSUBS 0.007128f
C538 B.n392 VSUBS 0.007128f
C539 B.n393 VSUBS 0.007128f
C540 B.n394 VSUBS 0.007128f
C541 B.n395 VSUBS 0.007128f
C542 B.n396 VSUBS 0.007128f
C543 B.n397 VSUBS 0.007128f
C544 B.n398 VSUBS 0.007128f
C545 B.n399 VSUBS 0.007128f
C546 B.n400 VSUBS 0.007128f
C547 B.n401 VSUBS 0.007128f
C548 B.n402 VSUBS 0.007128f
C549 B.n403 VSUBS 0.007128f
C550 B.n404 VSUBS 0.007128f
C551 B.n405 VSUBS 0.007128f
C552 B.n406 VSUBS 0.007128f
C553 B.n407 VSUBS 0.007128f
C554 B.n408 VSUBS 0.007128f
C555 B.n409 VSUBS 0.007128f
C556 B.n410 VSUBS 0.007128f
C557 B.n411 VSUBS 0.007128f
C558 B.n412 VSUBS 0.007128f
C559 B.n413 VSUBS 0.007128f
C560 B.n414 VSUBS 0.007128f
C561 B.n415 VSUBS 0.009302f
C562 B.n416 VSUBS 0.009909f
C563 B.n417 VSUBS 0.019705f
C564 VDD2.n0 VSUBS 0.02472f
C565 VDD2.n1 VSUBS 0.024377f
C566 VDD2.n2 VSUBS 0.013099f
C567 VDD2.n3 VSUBS 0.030961f
C568 VDD2.n4 VSUBS 0.01387f
C569 VDD2.n5 VSUBS 0.387038f
C570 VDD2.n6 VSUBS 0.013099f
C571 VDD2.t3 VSUBS 0.066809f
C572 VDD2.n7 VSUBS 0.096858f
C573 VDD2.n8 VSUBS 0.019614f
C574 VDD2.n9 VSUBS 0.023221f
C575 VDD2.n10 VSUBS 0.030961f
C576 VDD2.n11 VSUBS 0.01387f
C577 VDD2.n12 VSUBS 0.013099f
C578 VDD2.n13 VSUBS 0.024377f
C579 VDD2.n14 VSUBS 0.024377f
C580 VDD2.n15 VSUBS 0.013099f
C581 VDD2.n16 VSUBS 0.01387f
C582 VDD2.n17 VSUBS 0.030961f
C583 VDD2.n18 VSUBS 0.067919f
C584 VDD2.n19 VSUBS 0.01387f
C585 VDD2.n20 VSUBS 0.013099f
C586 VDD2.n21 VSUBS 0.052682f
C587 VDD2.n22 VSUBS 0.052794f
C588 VDD2.t7 VSUBS 0.085721f
C589 VDD2.t8 VSUBS 0.085721f
C590 VDD2.n23 VSUBS 0.517926f
C591 VDD2.n24 VSUBS 0.561323f
C592 VDD2.t2 VSUBS 0.085721f
C593 VDD2.t6 VSUBS 0.085721f
C594 VDD2.n25 VSUBS 0.520908f
C595 VDD2.n26 VSUBS 1.59051f
C596 VDD2.n27 VSUBS 0.02472f
C597 VDD2.n28 VSUBS 0.024377f
C598 VDD2.n29 VSUBS 0.013099f
C599 VDD2.n30 VSUBS 0.030961f
C600 VDD2.n31 VSUBS 0.01387f
C601 VDD2.n32 VSUBS 0.387038f
C602 VDD2.n33 VSUBS 0.013099f
C603 VDD2.t9 VSUBS 0.066809f
C604 VDD2.n34 VSUBS 0.096858f
C605 VDD2.n35 VSUBS 0.019614f
C606 VDD2.n36 VSUBS 0.023221f
C607 VDD2.n37 VSUBS 0.030961f
C608 VDD2.n38 VSUBS 0.01387f
C609 VDD2.n39 VSUBS 0.013099f
C610 VDD2.n40 VSUBS 0.024377f
C611 VDD2.n41 VSUBS 0.024377f
C612 VDD2.n42 VSUBS 0.013099f
C613 VDD2.n43 VSUBS 0.01387f
C614 VDD2.n44 VSUBS 0.030961f
C615 VDD2.n45 VSUBS 0.067919f
C616 VDD2.n46 VSUBS 0.01387f
C617 VDD2.n47 VSUBS 0.013099f
C618 VDD2.n48 VSUBS 0.052682f
C619 VDD2.n49 VSUBS 0.050591f
C620 VDD2.n50 VSUBS 1.51891f
C621 VDD2.t0 VSUBS 0.085721f
C622 VDD2.t1 VSUBS 0.085721f
C623 VDD2.n51 VSUBS 0.517929f
C624 VDD2.n52 VSUBS 0.453194f
C625 VDD2.t4 VSUBS 0.085721f
C626 VDD2.t5 VSUBS 0.085721f
C627 VDD2.n53 VSUBS 0.520888f
C628 VTAIL.t10 VSUBS 0.099859f
C629 VTAIL.t13 VSUBS 0.099859f
C630 VTAIL.n0 VSUBS 0.52243f
C631 VTAIL.n1 VSUBS 0.613254f
C632 VTAIL.n2 VSUBS 0.028797f
C633 VTAIL.n3 VSUBS 0.028397f
C634 VTAIL.n4 VSUBS 0.015259f
C635 VTAIL.n5 VSUBS 0.036068f
C636 VTAIL.n6 VSUBS 0.016157f
C637 VTAIL.n7 VSUBS 0.450873f
C638 VTAIL.n8 VSUBS 0.015259f
C639 VTAIL.t1 VSUBS 0.077828f
C640 VTAIL.n9 VSUBS 0.112833f
C641 VTAIL.n10 VSUBS 0.022849f
C642 VTAIL.n11 VSUBS 0.027051f
C643 VTAIL.n12 VSUBS 0.036068f
C644 VTAIL.n13 VSUBS 0.016157f
C645 VTAIL.n14 VSUBS 0.015259f
C646 VTAIL.n15 VSUBS 0.028397f
C647 VTAIL.n16 VSUBS 0.028397f
C648 VTAIL.n17 VSUBS 0.015259f
C649 VTAIL.n18 VSUBS 0.016157f
C650 VTAIL.n19 VSUBS 0.036068f
C651 VTAIL.n20 VSUBS 0.079121f
C652 VTAIL.n21 VSUBS 0.016157f
C653 VTAIL.n22 VSUBS 0.015259f
C654 VTAIL.n23 VSUBS 0.061372f
C655 VTAIL.n24 VSUBS 0.03929f
C656 VTAIL.n25 VSUBS 0.189077f
C657 VTAIL.t17 VSUBS 0.099859f
C658 VTAIL.t2 VSUBS 0.099859f
C659 VTAIL.n26 VSUBS 0.52243f
C660 VTAIL.n27 VSUBS 0.627058f
C661 VTAIL.t4 VSUBS 0.099859f
C662 VTAIL.t5 VSUBS 0.099859f
C663 VTAIL.n28 VSUBS 0.52243f
C664 VTAIL.n29 VSUBS 1.44665f
C665 VTAIL.t15 VSUBS 0.099859f
C666 VTAIL.t11 VSUBS 0.099859f
C667 VTAIL.n30 VSUBS 0.522434f
C668 VTAIL.n31 VSUBS 1.44664f
C669 VTAIL.t9 VSUBS 0.099859f
C670 VTAIL.t8 VSUBS 0.099859f
C671 VTAIL.n32 VSUBS 0.522434f
C672 VTAIL.n33 VSUBS 0.627055f
C673 VTAIL.n34 VSUBS 0.028797f
C674 VTAIL.n35 VSUBS 0.028397f
C675 VTAIL.n36 VSUBS 0.015259f
C676 VTAIL.n37 VSUBS 0.036068f
C677 VTAIL.n38 VSUBS 0.016157f
C678 VTAIL.n39 VSUBS 0.450873f
C679 VTAIL.n40 VSUBS 0.015259f
C680 VTAIL.t14 VSUBS 0.077828f
C681 VTAIL.n41 VSUBS 0.112833f
C682 VTAIL.n42 VSUBS 0.022849f
C683 VTAIL.n43 VSUBS 0.027051f
C684 VTAIL.n44 VSUBS 0.036068f
C685 VTAIL.n45 VSUBS 0.016157f
C686 VTAIL.n46 VSUBS 0.015259f
C687 VTAIL.n47 VSUBS 0.028397f
C688 VTAIL.n48 VSUBS 0.028397f
C689 VTAIL.n49 VSUBS 0.015259f
C690 VTAIL.n50 VSUBS 0.016157f
C691 VTAIL.n51 VSUBS 0.036068f
C692 VTAIL.n52 VSUBS 0.079121f
C693 VTAIL.n53 VSUBS 0.016157f
C694 VTAIL.n54 VSUBS 0.015259f
C695 VTAIL.n55 VSUBS 0.061372f
C696 VTAIL.n56 VSUBS 0.03929f
C697 VTAIL.n57 VSUBS 0.189077f
C698 VTAIL.t3 VSUBS 0.099859f
C699 VTAIL.t6 VSUBS 0.099859f
C700 VTAIL.n58 VSUBS 0.522434f
C701 VTAIL.n59 VSUBS 0.628632f
C702 VTAIL.t18 VSUBS 0.099859f
C703 VTAIL.t0 VSUBS 0.099859f
C704 VTAIL.n60 VSUBS 0.522434f
C705 VTAIL.n61 VSUBS 0.627055f
C706 VTAIL.n62 VSUBS 0.028797f
C707 VTAIL.n63 VSUBS 0.028397f
C708 VTAIL.n64 VSUBS 0.015259f
C709 VTAIL.n65 VSUBS 0.036068f
C710 VTAIL.n66 VSUBS 0.016157f
C711 VTAIL.n67 VSUBS 0.450873f
C712 VTAIL.n68 VSUBS 0.015259f
C713 VTAIL.t19 VSUBS 0.077828f
C714 VTAIL.n69 VSUBS 0.112833f
C715 VTAIL.n70 VSUBS 0.022849f
C716 VTAIL.n71 VSUBS 0.027051f
C717 VTAIL.n72 VSUBS 0.036068f
C718 VTAIL.n73 VSUBS 0.016157f
C719 VTAIL.n74 VSUBS 0.015259f
C720 VTAIL.n75 VSUBS 0.028397f
C721 VTAIL.n76 VSUBS 0.028397f
C722 VTAIL.n77 VSUBS 0.015259f
C723 VTAIL.n78 VSUBS 0.016157f
C724 VTAIL.n79 VSUBS 0.036068f
C725 VTAIL.n80 VSUBS 0.079121f
C726 VTAIL.n81 VSUBS 0.016157f
C727 VTAIL.n82 VSUBS 0.015259f
C728 VTAIL.n83 VSUBS 0.061372f
C729 VTAIL.n84 VSUBS 0.03929f
C730 VTAIL.n85 VSUBS 0.924263f
C731 VTAIL.n86 VSUBS 0.028797f
C732 VTAIL.n87 VSUBS 0.028397f
C733 VTAIL.n88 VSUBS 0.015259f
C734 VTAIL.n89 VSUBS 0.036068f
C735 VTAIL.n90 VSUBS 0.016157f
C736 VTAIL.n91 VSUBS 0.450873f
C737 VTAIL.n92 VSUBS 0.015259f
C738 VTAIL.t7 VSUBS 0.077828f
C739 VTAIL.n93 VSUBS 0.112833f
C740 VTAIL.n94 VSUBS 0.022849f
C741 VTAIL.n95 VSUBS 0.027051f
C742 VTAIL.n96 VSUBS 0.036068f
C743 VTAIL.n97 VSUBS 0.016157f
C744 VTAIL.n98 VSUBS 0.015259f
C745 VTAIL.n99 VSUBS 0.028397f
C746 VTAIL.n100 VSUBS 0.028397f
C747 VTAIL.n101 VSUBS 0.015259f
C748 VTAIL.n102 VSUBS 0.016157f
C749 VTAIL.n103 VSUBS 0.036068f
C750 VTAIL.n104 VSUBS 0.079121f
C751 VTAIL.n105 VSUBS 0.016157f
C752 VTAIL.n106 VSUBS 0.015259f
C753 VTAIL.n107 VSUBS 0.061372f
C754 VTAIL.n108 VSUBS 0.03929f
C755 VTAIL.n109 VSUBS 0.924263f
C756 VTAIL.t16 VSUBS 0.099859f
C757 VTAIL.t12 VSUBS 0.099859f
C758 VTAIL.n110 VSUBS 0.52243f
C759 VTAIL.n111 VSUBS 0.559615f
C760 VN.n0 VSUBS 0.061596f
C761 VN.n1 VSUBS 0.013977f
C762 VN.n2 VSUBS 0.261039f
C763 VN.t6 VSUBS 0.610234f
C764 VN.n3 VSUBS 0.267211f
C765 VN.t2 VSUBS 0.579595f
C766 VN.n4 VSUBS 0.299356f
C767 VN.n5 VSUBS 0.013977f
C768 VN.t1 VSUBS 0.579595f
C769 VN.n6 VSUBS 0.291726f
C770 VN.n7 VSUBS 0.061596f
C771 VN.n8 VSUBS 0.061596f
C772 VN.n9 VSUBS 0.061596f
C773 VN.t7 VSUBS 0.579595f
C774 VN.n10 VSUBS 0.291726f
C775 VN.n11 VSUBS 0.013977f
C776 VN.t3 VSUBS 0.579595f
C777 VN.n12 VSUBS 0.290207f
C778 VN.n13 VSUBS 0.047735f
C779 VN.n14 VSUBS 0.061596f
C780 VN.n15 VSUBS 0.013977f
C781 VN.t9 VSUBS 0.579595f
C782 VN.n16 VSUBS 0.261039f
C783 VN.t4 VSUBS 0.610234f
C784 VN.n17 VSUBS 0.267211f
C785 VN.t5 VSUBS 0.579595f
C786 VN.n18 VSUBS 0.299356f
C787 VN.n19 VSUBS 0.013977f
C788 VN.t8 VSUBS 0.579595f
C789 VN.n20 VSUBS 0.291726f
C790 VN.n21 VSUBS 0.061596f
C791 VN.n22 VSUBS 0.061596f
C792 VN.n23 VSUBS 0.061596f
C793 VN.n24 VSUBS 0.291726f
C794 VN.n25 VSUBS 0.013977f
C795 VN.t0 VSUBS 0.579595f
C796 VN.n26 VSUBS 0.290207f
C797 VN.n27 VSUBS 2.09952f
.ends

