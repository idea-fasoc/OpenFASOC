* NGSPICE file created from diff_pair_sample_1476.ext - technology: sky130A

.subckt diff_pair_sample_1476 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=3.12345 ps=19.26 w=18.93 l=2.82
X1 B.t11 B.t9 B.t10 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=0 ps=0 w=18.93 l=2.82
X2 B.t8 B.t6 B.t7 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=0 ps=0 w=18.93 l=2.82
X3 VTAIL.t6 VP.t1 VDD1.t0 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=3.12345 ps=19.26 w=18.93 l=2.82
X4 B.t5 B.t3 B.t4 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=0 ps=0 w=18.93 l=2.82
X5 VDD1.t2 VP.t2 VTAIL.t5 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=3.12345 pd=19.26 as=7.3827 ps=38.64 w=18.93 l=2.82
X6 VDD2.t3 VN.t0 VTAIL.t0 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=3.12345 pd=19.26 as=7.3827 ps=38.64 w=18.93 l=2.82
X7 VDD2.t2 VN.t1 VTAIL.t2 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=3.12345 pd=19.26 as=7.3827 ps=38.64 w=18.93 l=2.82
X8 VDD1.t3 VP.t3 VTAIL.t4 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=3.12345 pd=19.26 as=7.3827 ps=38.64 w=18.93 l=2.82
X9 VTAIL.t3 VN.t2 VDD2.t1 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=3.12345 ps=19.26 w=18.93 l=2.82
X10 VTAIL.t1 VN.t3 VDD2.t0 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=3.12345 ps=19.26 w=18.93 l=2.82
X11 B.t2 B.t0 B.t1 w_n2860_n4754# sky130_fd_pr__pfet_01v8 ad=7.3827 pd=38.64 as=0 ps=0 w=18.93 l=2.82
R0 VP.n4 VP.t1 196.916
R1 VP.n4 VP.t3 196.024
R2 VP.n5 VP.t0 161.779
R3 VP.n17 VP.t2 161.779
R4 VP.n16 VP.n0 161.3
R5 VP.n15 VP.n14 161.3
R6 VP.n13 VP.n1 161.3
R7 VP.n12 VP.n11 161.3
R8 VP.n10 VP.n2 161.3
R9 VP.n9 VP.n8 161.3
R10 VP.n7 VP.n3 161.3
R11 VP.n6 VP.n5 107.087
R12 VP.n18 VP.n17 107.087
R13 VP.n6 VP.n4 55.7043
R14 VP.n11 VP.n10 40.4934
R15 VP.n11 VP.n1 40.4934
R16 VP.n9 VP.n3 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n1 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n5 VP.n3 3.67055
R21 VP.n17 VP.n16 3.67055
R22 VP.n7 VP.n6 0.278367
R23 VP.n18 VP.n0 0.278367
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153454
R31 VDD1 VDD1.n1 116.508
R32 VDD1 VDD1.n0 67.8611
R33 VDD1.n0 VDD1.t0 1.71762
R34 VDD1.n0 VDD1.t3 1.71762
R35 VDD1.n1 VDD1.t1 1.71762
R36 VDD1.n1 VDD1.t2 1.71762
R37 VTAIL.n842 VTAIL.n742 756.745
R38 VTAIL.n100 VTAIL.n0 756.745
R39 VTAIL.n206 VTAIL.n106 756.745
R40 VTAIL.n312 VTAIL.n212 756.745
R41 VTAIL.n736 VTAIL.n636 756.745
R42 VTAIL.n630 VTAIL.n530 756.745
R43 VTAIL.n524 VTAIL.n424 756.745
R44 VTAIL.n418 VTAIL.n318 756.745
R45 VTAIL.n777 VTAIL.n776 585
R46 VTAIL.n774 VTAIL.n773 585
R47 VTAIL.n783 VTAIL.n782 585
R48 VTAIL.n785 VTAIL.n784 585
R49 VTAIL.n770 VTAIL.n769 585
R50 VTAIL.n791 VTAIL.n790 585
R51 VTAIL.n793 VTAIL.n792 585
R52 VTAIL.n766 VTAIL.n765 585
R53 VTAIL.n799 VTAIL.n798 585
R54 VTAIL.n801 VTAIL.n800 585
R55 VTAIL.n762 VTAIL.n761 585
R56 VTAIL.n807 VTAIL.n806 585
R57 VTAIL.n809 VTAIL.n808 585
R58 VTAIL.n758 VTAIL.n757 585
R59 VTAIL.n815 VTAIL.n814 585
R60 VTAIL.n818 VTAIL.n817 585
R61 VTAIL.n816 VTAIL.n754 585
R62 VTAIL.n823 VTAIL.n753 585
R63 VTAIL.n825 VTAIL.n824 585
R64 VTAIL.n827 VTAIL.n826 585
R65 VTAIL.n750 VTAIL.n749 585
R66 VTAIL.n833 VTAIL.n832 585
R67 VTAIL.n835 VTAIL.n834 585
R68 VTAIL.n746 VTAIL.n745 585
R69 VTAIL.n841 VTAIL.n840 585
R70 VTAIL.n843 VTAIL.n842 585
R71 VTAIL.n35 VTAIL.n34 585
R72 VTAIL.n32 VTAIL.n31 585
R73 VTAIL.n41 VTAIL.n40 585
R74 VTAIL.n43 VTAIL.n42 585
R75 VTAIL.n28 VTAIL.n27 585
R76 VTAIL.n49 VTAIL.n48 585
R77 VTAIL.n51 VTAIL.n50 585
R78 VTAIL.n24 VTAIL.n23 585
R79 VTAIL.n57 VTAIL.n56 585
R80 VTAIL.n59 VTAIL.n58 585
R81 VTAIL.n20 VTAIL.n19 585
R82 VTAIL.n65 VTAIL.n64 585
R83 VTAIL.n67 VTAIL.n66 585
R84 VTAIL.n16 VTAIL.n15 585
R85 VTAIL.n73 VTAIL.n72 585
R86 VTAIL.n76 VTAIL.n75 585
R87 VTAIL.n74 VTAIL.n12 585
R88 VTAIL.n81 VTAIL.n11 585
R89 VTAIL.n83 VTAIL.n82 585
R90 VTAIL.n85 VTAIL.n84 585
R91 VTAIL.n8 VTAIL.n7 585
R92 VTAIL.n91 VTAIL.n90 585
R93 VTAIL.n93 VTAIL.n92 585
R94 VTAIL.n4 VTAIL.n3 585
R95 VTAIL.n99 VTAIL.n98 585
R96 VTAIL.n101 VTAIL.n100 585
R97 VTAIL.n141 VTAIL.n140 585
R98 VTAIL.n138 VTAIL.n137 585
R99 VTAIL.n147 VTAIL.n146 585
R100 VTAIL.n149 VTAIL.n148 585
R101 VTAIL.n134 VTAIL.n133 585
R102 VTAIL.n155 VTAIL.n154 585
R103 VTAIL.n157 VTAIL.n156 585
R104 VTAIL.n130 VTAIL.n129 585
R105 VTAIL.n163 VTAIL.n162 585
R106 VTAIL.n165 VTAIL.n164 585
R107 VTAIL.n126 VTAIL.n125 585
R108 VTAIL.n171 VTAIL.n170 585
R109 VTAIL.n173 VTAIL.n172 585
R110 VTAIL.n122 VTAIL.n121 585
R111 VTAIL.n179 VTAIL.n178 585
R112 VTAIL.n182 VTAIL.n181 585
R113 VTAIL.n180 VTAIL.n118 585
R114 VTAIL.n187 VTAIL.n117 585
R115 VTAIL.n189 VTAIL.n188 585
R116 VTAIL.n191 VTAIL.n190 585
R117 VTAIL.n114 VTAIL.n113 585
R118 VTAIL.n197 VTAIL.n196 585
R119 VTAIL.n199 VTAIL.n198 585
R120 VTAIL.n110 VTAIL.n109 585
R121 VTAIL.n205 VTAIL.n204 585
R122 VTAIL.n207 VTAIL.n206 585
R123 VTAIL.n247 VTAIL.n246 585
R124 VTAIL.n244 VTAIL.n243 585
R125 VTAIL.n253 VTAIL.n252 585
R126 VTAIL.n255 VTAIL.n254 585
R127 VTAIL.n240 VTAIL.n239 585
R128 VTAIL.n261 VTAIL.n260 585
R129 VTAIL.n263 VTAIL.n262 585
R130 VTAIL.n236 VTAIL.n235 585
R131 VTAIL.n269 VTAIL.n268 585
R132 VTAIL.n271 VTAIL.n270 585
R133 VTAIL.n232 VTAIL.n231 585
R134 VTAIL.n277 VTAIL.n276 585
R135 VTAIL.n279 VTAIL.n278 585
R136 VTAIL.n228 VTAIL.n227 585
R137 VTAIL.n285 VTAIL.n284 585
R138 VTAIL.n288 VTAIL.n287 585
R139 VTAIL.n286 VTAIL.n224 585
R140 VTAIL.n293 VTAIL.n223 585
R141 VTAIL.n295 VTAIL.n294 585
R142 VTAIL.n297 VTAIL.n296 585
R143 VTAIL.n220 VTAIL.n219 585
R144 VTAIL.n303 VTAIL.n302 585
R145 VTAIL.n305 VTAIL.n304 585
R146 VTAIL.n216 VTAIL.n215 585
R147 VTAIL.n311 VTAIL.n310 585
R148 VTAIL.n313 VTAIL.n312 585
R149 VTAIL.n737 VTAIL.n736 585
R150 VTAIL.n735 VTAIL.n734 585
R151 VTAIL.n640 VTAIL.n639 585
R152 VTAIL.n729 VTAIL.n728 585
R153 VTAIL.n727 VTAIL.n726 585
R154 VTAIL.n644 VTAIL.n643 585
R155 VTAIL.n721 VTAIL.n720 585
R156 VTAIL.n719 VTAIL.n718 585
R157 VTAIL.n717 VTAIL.n647 585
R158 VTAIL.n651 VTAIL.n648 585
R159 VTAIL.n712 VTAIL.n711 585
R160 VTAIL.n710 VTAIL.n709 585
R161 VTAIL.n653 VTAIL.n652 585
R162 VTAIL.n704 VTAIL.n703 585
R163 VTAIL.n702 VTAIL.n701 585
R164 VTAIL.n657 VTAIL.n656 585
R165 VTAIL.n696 VTAIL.n695 585
R166 VTAIL.n694 VTAIL.n693 585
R167 VTAIL.n661 VTAIL.n660 585
R168 VTAIL.n688 VTAIL.n687 585
R169 VTAIL.n686 VTAIL.n685 585
R170 VTAIL.n665 VTAIL.n664 585
R171 VTAIL.n680 VTAIL.n679 585
R172 VTAIL.n678 VTAIL.n677 585
R173 VTAIL.n669 VTAIL.n668 585
R174 VTAIL.n672 VTAIL.n671 585
R175 VTAIL.n631 VTAIL.n630 585
R176 VTAIL.n629 VTAIL.n628 585
R177 VTAIL.n534 VTAIL.n533 585
R178 VTAIL.n623 VTAIL.n622 585
R179 VTAIL.n621 VTAIL.n620 585
R180 VTAIL.n538 VTAIL.n537 585
R181 VTAIL.n615 VTAIL.n614 585
R182 VTAIL.n613 VTAIL.n612 585
R183 VTAIL.n611 VTAIL.n541 585
R184 VTAIL.n545 VTAIL.n542 585
R185 VTAIL.n606 VTAIL.n605 585
R186 VTAIL.n604 VTAIL.n603 585
R187 VTAIL.n547 VTAIL.n546 585
R188 VTAIL.n598 VTAIL.n597 585
R189 VTAIL.n596 VTAIL.n595 585
R190 VTAIL.n551 VTAIL.n550 585
R191 VTAIL.n590 VTAIL.n589 585
R192 VTAIL.n588 VTAIL.n587 585
R193 VTAIL.n555 VTAIL.n554 585
R194 VTAIL.n582 VTAIL.n581 585
R195 VTAIL.n580 VTAIL.n579 585
R196 VTAIL.n559 VTAIL.n558 585
R197 VTAIL.n574 VTAIL.n573 585
R198 VTAIL.n572 VTAIL.n571 585
R199 VTAIL.n563 VTAIL.n562 585
R200 VTAIL.n566 VTAIL.n565 585
R201 VTAIL.n525 VTAIL.n524 585
R202 VTAIL.n523 VTAIL.n522 585
R203 VTAIL.n428 VTAIL.n427 585
R204 VTAIL.n517 VTAIL.n516 585
R205 VTAIL.n515 VTAIL.n514 585
R206 VTAIL.n432 VTAIL.n431 585
R207 VTAIL.n509 VTAIL.n508 585
R208 VTAIL.n507 VTAIL.n506 585
R209 VTAIL.n505 VTAIL.n435 585
R210 VTAIL.n439 VTAIL.n436 585
R211 VTAIL.n500 VTAIL.n499 585
R212 VTAIL.n498 VTAIL.n497 585
R213 VTAIL.n441 VTAIL.n440 585
R214 VTAIL.n492 VTAIL.n491 585
R215 VTAIL.n490 VTAIL.n489 585
R216 VTAIL.n445 VTAIL.n444 585
R217 VTAIL.n484 VTAIL.n483 585
R218 VTAIL.n482 VTAIL.n481 585
R219 VTAIL.n449 VTAIL.n448 585
R220 VTAIL.n476 VTAIL.n475 585
R221 VTAIL.n474 VTAIL.n473 585
R222 VTAIL.n453 VTAIL.n452 585
R223 VTAIL.n468 VTAIL.n467 585
R224 VTAIL.n466 VTAIL.n465 585
R225 VTAIL.n457 VTAIL.n456 585
R226 VTAIL.n460 VTAIL.n459 585
R227 VTAIL.n419 VTAIL.n418 585
R228 VTAIL.n417 VTAIL.n416 585
R229 VTAIL.n322 VTAIL.n321 585
R230 VTAIL.n411 VTAIL.n410 585
R231 VTAIL.n409 VTAIL.n408 585
R232 VTAIL.n326 VTAIL.n325 585
R233 VTAIL.n403 VTAIL.n402 585
R234 VTAIL.n401 VTAIL.n400 585
R235 VTAIL.n399 VTAIL.n329 585
R236 VTAIL.n333 VTAIL.n330 585
R237 VTAIL.n394 VTAIL.n393 585
R238 VTAIL.n392 VTAIL.n391 585
R239 VTAIL.n335 VTAIL.n334 585
R240 VTAIL.n386 VTAIL.n385 585
R241 VTAIL.n384 VTAIL.n383 585
R242 VTAIL.n339 VTAIL.n338 585
R243 VTAIL.n378 VTAIL.n377 585
R244 VTAIL.n376 VTAIL.n375 585
R245 VTAIL.n343 VTAIL.n342 585
R246 VTAIL.n370 VTAIL.n369 585
R247 VTAIL.n368 VTAIL.n367 585
R248 VTAIL.n347 VTAIL.n346 585
R249 VTAIL.n362 VTAIL.n361 585
R250 VTAIL.n360 VTAIL.n359 585
R251 VTAIL.n351 VTAIL.n350 585
R252 VTAIL.n354 VTAIL.n353 585
R253 VTAIL.t4 VTAIL.n670 327.466
R254 VTAIL.t6 VTAIL.n564 327.466
R255 VTAIL.t0 VTAIL.n458 327.466
R256 VTAIL.t3 VTAIL.n352 327.466
R257 VTAIL.t2 VTAIL.n775 327.466
R258 VTAIL.t1 VTAIL.n33 327.466
R259 VTAIL.t5 VTAIL.n139 327.466
R260 VTAIL.t7 VTAIL.n245 327.466
R261 VTAIL.n776 VTAIL.n773 171.744
R262 VTAIL.n783 VTAIL.n773 171.744
R263 VTAIL.n784 VTAIL.n783 171.744
R264 VTAIL.n784 VTAIL.n769 171.744
R265 VTAIL.n791 VTAIL.n769 171.744
R266 VTAIL.n792 VTAIL.n791 171.744
R267 VTAIL.n792 VTAIL.n765 171.744
R268 VTAIL.n799 VTAIL.n765 171.744
R269 VTAIL.n800 VTAIL.n799 171.744
R270 VTAIL.n800 VTAIL.n761 171.744
R271 VTAIL.n807 VTAIL.n761 171.744
R272 VTAIL.n808 VTAIL.n807 171.744
R273 VTAIL.n808 VTAIL.n757 171.744
R274 VTAIL.n815 VTAIL.n757 171.744
R275 VTAIL.n817 VTAIL.n815 171.744
R276 VTAIL.n817 VTAIL.n816 171.744
R277 VTAIL.n816 VTAIL.n753 171.744
R278 VTAIL.n825 VTAIL.n753 171.744
R279 VTAIL.n826 VTAIL.n825 171.744
R280 VTAIL.n826 VTAIL.n749 171.744
R281 VTAIL.n833 VTAIL.n749 171.744
R282 VTAIL.n834 VTAIL.n833 171.744
R283 VTAIL.n834 VTAIL.n745 171.744
R284 VTAIL.n841 VTAIL.n745 171.744
R285 VTAIL.n842 VTAIL.n841 171.744
R286 VTAIL.n34 VTAIL.n31 171.744
R287 VTAIL.n41 VTAIL.n31 171.744
R288 VTAIL.n42 VTAIL.n41 171.744
R289 VTAIL.n42 VTAIL.n27 171.744
R290 VTAIL.n49 VTAIL.n27 171.744
R291 VTAIL.n50 VTAIL.n49 171.744
R292 VTAIL.n50 VTAIL.n23 171.744
R293 VTAIL.n57 VTAIL.n23 171.744
R294 VTAIL.n58 VTAIL.n57 171.744
R295 VTAIL.n58 VTAIL.n19 171.744
R296 VTAIL.n65 VTAIL.n19 171.744
R297 VTAIL.n66 VTAIL.n65 171.744
R298 VTAIL.n66 VTAIL.n15 171.744
R299 VTAIL.n73 VTAIL.n15 171.744
R300 VTAIL.n75 VTAIL.n73 171.744
R301 VTAIL.n75 VTAIL.n74 171.744
R302 VTAIL.n74 VTAIL.n11 171.744
R303 VTAIL.n83 VTAIL.n11 171.744
R304 VTAIL.n84 VTAIL.n83 171.744
R305 VTAIL.n84 VTAIL.n7 171.744
R306 VTAIL.n91 VTAIL.n7 171.744
R307 VTAIL.n92 VTAIL.n91 171.744
R308 VTAIL.n92 VTAIL.n3 171.744
R309 VTAIL.n99 VTAIL.n3 171.744
R310 VTAIL.n100 VTAIL.n99 171.744
R311 VTAIL.n140 VTAIL.n137 171.744
R312 VTAIL.n147 VTAIL.n137 171.744
R313 VTAIL.n148 VTAIL.n147 171.744
R314 VTAIL.n148 VTAIL.n133 171.744
R315 VTAIL.n155 VTAIL.n133 171.744
R316 VTAIL.n156 VTAIL.n155 171.744
R317 VTAIL.n156 VTAIL.n129 171.744
R318 VTAIL.n163 VTAIL.n129 171.744
R319 VTAIL.n164 VTAIL.n163 171.744
R320 VTAIL.n164 VTAIL.n125 171.744
R321 VTAIL.n171 VTAIL.n125 171.744
R322 VTAIL.n172 VTAIL.n171 171.744
R323 VTAIL.n172 VTAIL.n121 171.744
R324 VTAIL.n179 VTAIL.n121 171.744
R325 VTAIL.n181 VTAIL.n179 171.744
R326 VTAIL.n181 VTAIL.n180 171.744
R327 VTAIL.n180 VTAIL.n117 171.744
R328 VTAIL.n189 VTAIL.n117 171.744
R329 VTAIL.n190 VTAIL.n189 171.744
R330 VTAIL.n190 VTAIL.n113 171.744
R331 VTAIL.n197 VTAIL.n113 171.744
R332 VTAIL.n198 VTAIL.n197 171.744
R333 VTAIL.n198 VTAIL.n109 171.744
R334 VTAIL.n205 VTAIL.n109 171.744
R335 VTAIL.n206 VTAIL.n205 171.744
R336 VTAIL.n246 VTAIL.n243 171.744
R337 VTAIL.n253 VTAIL.n243 171.744
R338 VTAIL.n254 VTAIL.n253 171.744
R339 VTAIL.n254 VTAIL.n239 171.744
R340 VTAIL.n261 VTAIL.n239 171.744
R341 VTAIL.n262 VTAIL.n261 171.744
R342 VTAIL.n262 VTAIL.n235 171.744
R343 VTAIL.n269 VTAIL.n235 171.744
R344 VTAIL.n270 VTAIL.n269 171.744
R345 VTAIL.n270 VTAIL.n231 171.744
R346 VTAIL.n277 VTAIL.n231 171.744
R347 VTAIL.n278 VTAIL.n277 171.744
R348 VTAIL.n278 VTAIL.n227 171.744
R349 VTAIL.n285 VTAIL.n227 171.744
R350 VTAIL.n287 VTAIL.n285 171.744
R351 VTAIL.n287 VTAIL.n286 171.744
R352 VTAIL.n286 VTAIL.n223 171.744
R353 VTAIL.n295 VTAIL.n223 171.744
R354 VTAIL.n296 VTAIL.n295 171.744
R355 VTAIL.n296 VTAIL.n219 171.744
R356 VTAIL.n303 VTAIL.n219 171.744
R357 VTAIL.n304 VTAIL.n303 171.744
R358 VTAIL.n304 VTAIL.n215 171.744
R359 VTAIL.n311 VTAIL.n215 171.744
R360 VTAIL.n312 VTAIL.n311 171.744
R361 VTAIL.n736 VTAIL.n735 171.744
R362 VTAIL.n735 VTAIL.n639 171.744
R363 VTAIL.n728 VTAIL.n639 171.744
R364 VTAIL.n728 VTAIL.n727 171.744
R365 VTAIL.n727 VTAIL.n643 171.744
R366 VTAIL.n720 VTAIL.n643 171.744
R367 VTAIL.n720 VTAIL.n719 171.744
R368 VTAIL.n719 VTAIL.n647 171.744
R369 VTAIL.n651 VTAIL.n647 171.744
R370 VTAIL.n711 VTAIL.n651 171.744
R371 VTAIL.n711 VTAIL.n710 171.744
R372 VTAIL.n710 VTAIL.n652 171.744
R373 VTAIL.n703 VTAIL.n652 171.744
R374 VTAIL.n703 VTAIL.n702 171.744
R375 VTAIL.n702 VTAIL.n656 171.744
R376 VTAIL.n695 VTAIL.n656 171.744
R377 VTAIL.n695 VTAIL.n694 171.744
R378 VTAIL.n694 VTAIL.n660 171.744
R379 VTAIL.n687 VTAIL.n660 171.744
R380 VTAIL.n687 VTAIL.n686 171.744
R381 VTAIL.n686 VTAIL.n664 171.744
R382 VTAIL.n679 VTAIL.n664 171.744
R383 VTAIL.n679 VTAIL.n678 171.744
R384 VTAIL.n678 VTAIL.n668 171.744
R385 VTAIL.n671 VTAIL.n668 171.744
R386 VTAIL.n630 VTAIL.n629 171.744
R387 VTAIL.n629 VTAIL.n533 171.744
R388 VTAIL.n622 VTAIL.n533 171.744
R389 VTAIL.n622 VTAIL.n621 171.744
R390 VTAIL.n621 VTAIL.n537 171.744
R391 VTAIL.n614 VTAIL.n537 171.744
R392 VTAIL.n614 VTAIL.n613 171.744
R393 VTAIL.n613 VTAIL.n541 171.744
R394 VTAIL.n545 VTAIL.n541 171.744
R395 VTAIL.n605 VTAIL.n545 171.744
R396 VTAIL.n605 VTAIL.n604 171.744
R397 VTAIL.n604 VTAIL.n546 171.744
R398 VTAIL.n597 VTAIL.n546 171.744
R399 VTAIL.n597 VTAIL.n596 171.744
R400 VTAIL.n596 VTAIL.n550 171.744
R401 VTAIL.n589 VTAIL.n550 171.744
R402 VTAIL.n589 VTAIL.n588 171.744
R403 VTAIL.n588 VTAIL.n554 171.744
R404 VTAIL.n581 VTAIL.n554 171.744
R405 VTAIL.n581 VTAIL.n580 171.744
R406 VTAIL.n580 VTAIL.n558 171.744
R407 VTAIL.n573 VTAIL.n558 171.744
R408 VTAIL.n573 VTAIL.n572 171.744
R409 VTAIL.n572 VTAIL.n562 171.744
R410 VTAIL.n565 VTAIL.n562 171.744
R411 VTAIL.n524 VTAIL.n523 171.744
R412 VTAIL.n523 VTAIL.n427 171.744
R413 VTAIL.n516 VTAIL.n427 171.744
R414 VTAIL.n516 VTAIL.n515 171.744
R415 VTAIL.n515 VTAIL.n431 171.744
R416 VTAIL.n508 VTAIL.n431 171.744
R417 VTAIL.n508 VTAIL.n507 171.744
R418 VTAIL.n507 VTAIL.n435 171.744
R419 VTAIL.n439 VTAIL.n435 171.744
R420 VTAIL.n499 VTAIL.n439 171.744
R421 VTAIL.n499 VTAIL.n498 171.744
R422 VTAIL.n498 VTAIL.n440 171.744
R423 VTAIL.n491 VTAIL.n440 171.744
R424 VTAIL.n491 VTAIL.n490 171.744
R425 VTAIL.n490 VTAIL.n444 171.744
R426 VTAIL.n483 VTAIL.n444 171.744
R427 VTAIL.n483 VTAIL.n482 171.744
R428 VTAIL.n482 VTAIL.n448 171.744
R429 VTAIL.n475 VTAIL.n448 171.744
R430 VTAIL.n475 VTAIL.n474 171.744
R431 VTAIL.n474 VTAIL.n452 171.744
R432 VTAIL.n467 VTAIL.n452 171.744
R433 VTAIL.n467 VTAIL.n466 171.744
R434 VTAIL.n466 VTAIL.n456 171.744
R435 VTAIL.n459 VTAIL.n456 171.744
R436 VTAIL.n418 VTAIL.n417 171.744
R437 VTAIL.n417 VTAIL.n321 171.744
R438 VTAIL.n410 VTAIL.n321 171.744
R439 VTAIL.n410 VTAIL.n409 171.744
R440 VTAIL.n409 VTAIL.n325 171.744
R441 VTAIL.n402 VTAIL.n325 171.744
R442 VTAIL.n402 VTAIL.n401 171.744
R443 VTAIL.n401 VTAIL.n329 171.744
R444 VTAIL.n333 VTAIL.n329 171.744
R445 VTAIL.n393 VTAIL.n333 171.744
R446 VTAIL.n393 VTAIL.n392 171.744
R447 VTAIL.n392 VTAIL.n334 171.744
R448 VTAIL.n385 VTAIL.n334 171.744
R449 VTAIL.n385 VTAIL.n384 171.744
R450 VTAIL.n384 VTAIL.n338 171.744
R451 VTAIL.n377 VTAIL.n338 171.744
R452 VTAIL.n377 VTAIL.n376 171.744
R453 VTAIL.n376 VTAIL.n342 171.744
R454 VTAIL.n369 VTAIL.n342 171.744
R455 VTAIL.n369 VTAIL.n368 171.744
R456 VTAIL.n368 VTAIL.n346 171.744
R457 VTAIL.n361 VTAIL.n346 171.744
R458 VTAIL.n361 VTAIL.n360 171.744
R459 VTAIL.n360 VTAIL.n350 171.744
R460 VTAIL.n353 VTAIL.n350 171.744
R461 VTAIL.n776 VTAIL.t2 85.8723
R462 VTAIL.n34 VTAIL.t1 85.8723
R463 VTAIL.n140 VTAIL.t5 85.8723
R464 VTAIL.n246 VTAIL.t7 85.8723
R465 VTAIL.n671 VTAIL.t4 85.8723
R466 VTAIL.n565 VTAIL.t6 85.8723
R467 VTAIL.n459 VTAIL.t0 85.8723
R468 VTAIL.n353 VTAIL.t3 85.8723
R469 VTAIL.n847 VTAIL.n846 31.6035
R470 VTAIL.n105 VTAIL.n104 31.6035
R471 VTAIL.n211 VTAIL.n210 31.6035
R472 VTAIL.n317 VTAIL.n316 31.6035
R473 VTAIL.n741 VTAIL.n740 31.6035
R474 VTAIL.n635 VTAIL.n634 31.6035
R475 VTAIL.n529 VTAIL.n528 31.6035
R476 VTAIL.n423 VTAIL.n422 31.6035
R477 VTAIL.n847 VTAIL.n741 31.4014
R478 VTAIL.n423 VTAIL.n317 31.4014
R479 VTAIL.n777 VTAIL.n775 16.3895
R480 VTAIL.n35 VTAIL.n33 16.3895
R481 VTAIL.n141 VTAIL.n139 16.3895
R482 VTAIL.n247 VTAIL.n245 16.3895
R483 VTAIL.n672 VTAIL.n670 16.3895
R484 VTAIL.n566 VTAIL.n564 16.3895
R485 VTAIL.n460 VTAIL.n458 16.3895
R486 VTAIL.n354 VTAIL.n352 16.3895
R487 VTAIL.n824 VTAIL.n823 13.1884
R488 VTAIL.n82 VTAIL.n81 13.1884
R489 VTAIL.n188 VTAIL.n187 13.1884
R490 VTAIL.n294 VTAIL.n293 13.1884
R491 VTAIL.n718 VTAIL.n717 13.1884
R492 VTAIL.n612 VTAIL.n611 13.1884
R493 VTAIL.n506 VTAIL.n505 13.1884
R494 VTAIL.n400 VTAIL.n399 13.1884
R495 VTAIL.n778 VTAIL.n774 12.8005
R496 VTAIL.n822 VTAIL.n754 12.8005
R497 VTAIL.n827 VTAIL.n752 12.8005
R498 VTAIL.n36 VTAIL.n32 12.8005
R499 VTAIL.n80 VTAIL.n12 12.8005
R500 VTAIL.n85 VTAIL.n10 12.8005
R501 VTAIL.n142 VTAIL.n138 12.8005
R502 VTAIL.n186 VTAIL.n118 12.8005
R503 VTAIL.n191 VTAIL.n116 12.8005
R504 VTAIL.n248 VTAIL.n244 12.8005
R505 VTAIL.n292 VTAIL.n224 12.8005
R506 VTAIL.n297 VTAIL.n222 12.8005
R507 VTAIL.n721 VTAIL.n646 12.8005
R508 VTAIL.n716 VTAIL.n648 12.8005
R509 VTAIL.n673 VTAIL.n669 12.8005
R510 VTAIL.n615 VTAIL.n540 12.8005
R511 VTAIL.n610 VTAIL.n542 12.8005
R512 VTAIL.n567 VTAIL.n563 12.8005
R513 VTAIL.n509 VTAIL.n434 12.8005
R514 VTAIL.n504 VTAIL.n436 12.8005
R515 VTAIL.n461 VTAIL.n457 12.8005
R516 VTAIL.n403 VTAIL.n328 12.8005
R517 VTAIL.n398 VTAIL.n330 12.8005
R518 VTAIL.n355 VTAIL.n351 12.8005
R519 VTAIL.n782 VTAIL.n781 12.0247
R520 VTAIL.n819 VTAIL.n818 12.0247
R521 VTAIL.n828 VTAIL.n750 12.0247
R522 VTAIL.n40 VTAIL.n39 12.0247
R523 VTAIL.n77 VTAIL.n76 12.0247
R524 VTAIL.n86 VTAIL.n8 12.0247
R525 VTAIL.n146 VTAIL.n145 12.0247
R526 VTAIL.n183 VTAIL.n182 12.0247
R527 VTAIL.n192 VTAIL.n114 12.0247
R528 VTAIL.n252 VTAIL.n251 12.0247
R529 VTAIL.n289 VTAIL.n288 12.0247
R530 VTAIL.n298 VTAIL.n220 12.0247
R531 VTAIL.n722 VTAIL.n644 12.0247
R532 VTAIL.n713 VTAIL.n712 12.0247
R533 VTAIL.n677 VTAIL.n676 12.0247
R534 VTAIL.n616 VTAIL.n538 12.0247
R535 VTAIL.n607 VTAIL.n606 12.0247
R536 VTAIL.n571 VTAIL.n570 12.0247
R537 VTAIL.n510 VTAIL.n432 12.0247
R538 VTAIL.n501 VTAIL.n500 12.0247
R539 VTAIL.n465 VTAIL.n464 12.0247
R540 VTAIL.n404 VTAIL.n326 12.0247
R541 VTAIL.n395 VTAIL.n394 12.0247
R542 VTAIL.n359 VTAIL.n358 12.0247
R543 VTAIL.n785 VTAIL.n772 11.249
R544 VTAIL.n814 VTAIL.n756 11.249
R545 VTAIL.n832 VTAIL.n831 11.249
R546 VTAIL.n43 VTAIL.n30 11.249
R547 VTAIL.n72 VTAIL.n14 11.249
R548 VTAIL.n90 VTAIL.n89 11.249
R549 VTAIL.n149 VTAIL.n136 11.249
R550 VTAIL.n178 VTAIL.n120 11.249
R551 VTAIL.n196 VTAIL.n195 11.249
R552 VTAIL.n255 VTAIL.n242 11.249
R553 VTAIL.n284 VTAIL.n226 11.249
R554 VTAIL.n302 VTAIL.n301 11.249
R555 VTAIL.n726 VTAIL.n725 11.249
R556 VTAIL.n709 VTAIL.n650 11.249
R557 VTAIL.n680 VTAIL.n667 11.249
R558 VTAIL.n620 VTAIL.n619 11.249
R559 VTAIL.n603 VTAIL.n544 11.249
R560 VTAIL.n574 VTAIL.n561 11.249
R561 VTAIL.n514 VTAIL.n513 11.249
R562 VTAIL.n497 VTAIL.n438 11.249
R563 VTAIL.n468 VTAIL.n455 11.249
R564 VTAIL.n408 VTAIL.n407 11.249
R565 VTAIL.n391 VTAIL.n332 11.249
R566 VTAIL.n362 VTAIL.n349 11.249
R567 VTAIL.n786 VTAIL.n770 10.4732
R568 VTAIL.n813 VTAIL.n758 10.4732
R569 VTAIL.n835 VTAIL.n748 10.4732
R570 VTAIL.n44 VTAIL.n28 10.4732
R571 VTAIL.n71 VTAIL.n16 10.4732
R572 VTAIL.n93 VTAIL.n6 10.4732
R573 VTAIL.n150 VTAIL.n134 10.4732
R574 VTAIL.n177 VTAIL.n122 10.4732
R575 VTAIL.n199 VTAIL.n112 10.4732
R576 VTAIL.n256 VTAIL.n240 10.4732
R577 VTAIL.n283 VTAIL.n228 10.4732
R578 VTAIL.n305 VTAIL.n218 10.4732
R579 VTAIL.n729 VTAIL.n642 10.4732
R580 VTAIL.n708 VTAIL.n653 10.4732
R581 VTAIL.n681 VTAIL.n665 10.4732
R582 VTAIL.n623 VTAIL.n536 10.4732
R583 VTAIL.n602 VTAIL.n547 10.4732
R584 VTAIL.n575 VTAIL.n559 10.4732
R585 VTAIL.n517 VTAIL.n430 10.4732
R586 VTAIL.n496 VTAIL.n441 10.4732
R587 VTAIL.n469 VTAIL.n453 10.4732
R588 VTAIL.n411 VTAIL.n324 10.4732
R589 VTAIL.n390 VTAIL.n335 10.4732
R590 VTAIL.n363 VTAIL.n347 10.4732
R591 VTAIL.n790 VTAIL.n789 9.69747
R592 VTAIL.n810 VTAIL.n809 9.69747
R593 VTAIL.n836 VTAIL.n746 9.69747
R594 VTAIL.n48 VTAIL.n47 9.69747
R595 VTAIL.n68 VTAIL.n67 9.69747
R596 VTAIL.n94 VTAIL.n4 9.69747
R597 VTAIL.n154 VTAIL.n153 9.69747
R598 VTAIL.n174 VTAIL.n173 9.69747
R599 VTAIL.n200 VTAIL.n110 9.69747
R600 VTAIL.n260 VTAIL.n259 9.69747
R601 VTAIL.n280 VTAIL.n279 9.69747
R602 VTAIL.n306 VTAIL.n216 9.69747
R603 VTAIL.n730 VTAIL.n640 9.69747
R604 VTAIL.n705 VTAIL.n704 9.69747
R605 VTAIL.n685 VTAIL.n684 9.69747
R606 VTAIL.n624 VTAIL.n534 9.69747
R607 VTAIL.n599 VTAIL.n598 9.69747
R608 VTAIL.n579 VTAIL.n578 9.69747
R609 VTAIL.n518 VTAIL.n428 9.69747
R610 VTAIL.n493 VTAIL.n492 9.69747
R611 VTAIL.n473 VTAIL.n472 9.69747
R612 VTAIL.n412 VTAIL.n322 9.69747
R613 VTAIL.n387 VTAIL.n386 9.69747
R614 VTAIL.n367 VTAIL.n366 9.69747
R615 VTAIL.n846 VTAIL.n845 9.45567
R616 VTAIL.n104 VTAIL.n103 9.45567
R617 VTAIL.n210 VTAIL.n209 9.45567
R618 VTAIL.n316 VTAIL.n315 9.45567
R619 VTAIL.n740 VTAIL.n739 9.45567
R620 VTAIL.n634 VTAIL.n633 9.45567
R621 VTAIL.n528 VTAIL.n527 9.45567
R622 VTAIL.n422 VTAIL.n421 9.45567
R623 VTAIL.n744 VTAIL.n743 9.3005
R624 VTAIL.n839 VTAIL.n838 9.3005
R625 VTAIL.n837 VTAIL.n836 9.3005
R626 VTAIL.n748 VTAIL.n747 9.3005
R627 VTAIL.n831 VTAIL.n830 9.3005
R628 VTAIL.n829 VTAIL.n828 9.3005
R629 VTAIL.n752 VTAIL.n751 9.3005
R630 VTAIL.n797 VTAIL.n796 9.3005
R631 VTAIL.n795 VTAIL.n794 9.3005
R632 VTAIL.n768 VTAIL.n767 9.3005
R633 VTAIL.n789 VTAIL.n788 9.3005
R634 VTAIL.n787 VTAIL.n786 9.3005
R635 VTAIL.n772 VTAIL.n771 9.3005
R636 VTAIL.n781 VTAIL.n780 9.3005
R637 VTAIL.n779 VTAIL.n778 9.3005
R638 VTAIL.n764 VTAIL.n763 9.3005
R639 VTAIL.n803 VTAIL.n802 9.3005
R640 VTAIL.n805 VTAIL.n804 9.3005
R641 VTAIL.n760 VTAIL.n759 9.3005
R642 VTAIL.n811 VTAIL.n810 9.3005
R643 VTAIL.n813 VTAIL.n812 9.3005
R644 VTAIL.n756 VTAIL.n755 9.3005
R645 VTAIL.n820 VTAIL.n819 9.3005
R646 VTAIL.n822 VTAIL.n821 9.3005
R647 VTAIL.n845 VTAIL.n844 9.3005
R648 VTAIL.n2 VTAIL.n1 9.3005
R649 VTAIL.n97 VTAIL.n96 9.3005
R650 VTAIL.n95 VTAIL.n94 9.3005
R651 VTAIL.n6 VTAIL.n5 9.3005
R652 VTAIL.n89 VTAIL.n88 9.3005
R653 VTAIL.n87 VTAIL.n86 9.3005
R654 VTAIL.n10 VTAIL.n9 9.3005
R655 VTAIL.n55 VTAIL.n54 9.3005
R656 VTAIL.n53 VTAIL.n52 9.3005
R657 VTAIL.n26 VTAIL.n25 9.3005
R658 VTAIL.n47 VTAIL.n46 9.3005
R659 VTAIL.n45 VTAIL.n44 9.3005
R660 VTAIL.n30 VTAIL.n29 9.3005
R661 VTAIL.n39 VTAIL.n38 9.3005
R662 VTAIL.n37 VTAIL.n36 9.3005
R663 VTAIL.n22 VTAIL.n21 9.3005
R664 VTAIL.n61 VTAIL.n60 9.3005
R665 VTAIL.n63 VTAIL.n62 9.3005
R666 VTAIL.n18 VTAIL.n17 9.3005
R667 VTAIL.n69 VTAIL.n68 9.3005
R668 VTAIL.n71 VTAIL.n70 9.3005
R669 VTAIL.n14 VTAIL.n13 9.3005
R670 VTAIL.n78 VTAIL.n77 9.3005
R671 VTAIL.n80 VTAIL.n79 9.3005
R672 VTAIL.n103 VTAIL.n102 9.3005
R673 VTAIL.n108 VTAIL.n107 9.3005
R674 VTAIL.n203 VTAIL.n202 9.3005
R675 VTAIL.n201 VTAIL.n200 9.3005
R676 VTAIL.n112 VTAIL.n111 9.3005
R677 VTAIL.n195 VTAIL.n194 9.3005
R678 VTAIL.n193 VTAIL.n192 9.3005
R679 VTAIL.n116 VTAIL.n115 9.3005
R680 VTAIL.n161 VTAIL.n160 9.3005
R681 VTAIL.n159 VTAIL.n158 9.3005
R682 VTAIL.n132 VTAIL.n131 9.3005
R683 VTAIL.n153 VTAIL.n152 9.3005
R684 VTAIL.n151 VTAIL.n150 9.3005
R685 VTAIL.n136 VTAIL.n135 9.3005
R686 VTAIL.n145 VTAIL.n144 9.3005
R687 VTAIL.n143 VTAIL.n142 9.3005
R688 VTAIL.n128 VTAIL.n127 9.3005
R689 VTAIL.n167 VTAIL.n166 9.3005
R690 VTAIL.n169 VTAIL.n168 9.3005
R691 VTAIL.n124 VTAIL.n123 9.3005
R692 VTAIL.n175 VTAIL.n174 9.3005
R693 VTAIL.n177 VTAIL.n176 9.3005
R694 VTAIL.n120 VTAIL.n119 9.3005
R695 VTAIL.n184 VTAIL.n183 9.3005
R696 VTAIL.n186 VTAIL.n185 9.3005
R697 VTAIL.n209 VTAIL.n208 9.3005
R698 VTAIL.n214 VTAIL.n213 9.3005
R699 VTAIL.n309 VTAIL.n308 9.3005
R700 VTAIL.n307 VTAIL.n306 9.3005
R701 VTAIL.n218 VTAIL.n217 9.3005
R702 VTAIL.n301 VTAIL.n300 9.3005
R703 VTAIL.n299 VTAIL.n298 9.3005
R704 VTAIL.n222 VTAIL.n221 9.3005
R705 VTAIL.n267 VTAIL.n266 9.3005
R706 VTAIL.n265 VTAIL.n264 9.3005
R707 VTAIL.n238 VTAIL.n237 9.3005
R708 VTAIL.n259 VTAIL.n258 9.3005
R709 VTAIL.n257 VTAIL.n256 9.3005
R710 VTAIL.n242 VTAIL.n241 9.3005
R711 VTAIL.n251 VTAIL.n250 9.3005
R712 VTAIL.n249 VTAIL.n248 9.3005
R713 VTAIL.n234 VTAIL.n233 9.3005
R714 VTAIL.n273 VTAIL.n272 9.3005
R715 VTAIL.n275 VTAIL.n274 9.3005
R716 VTAIL.n230 VTAIL.n229 9.3005
R717 VTAIL.n281 VTAIL.n280 9.3005
R718 VTAIL.n283 VTAIL.n282 9.3005
R719 VTAIL.n226 VTAIL.n225 9.3005
R720 VTAIL.n290 VTAIL.n289 9.3005
R721 VTAIL.n292 VTAIL.n291 9.3005
R722 VTAIL.n315 VTAIL.n314 9.3005
R723 VTAIL.n698 VTAIL.n697 9.3005
R724 VTAIL.n700 VTAIL.n699 9.3005
R725 VTAIL.n655 VTAIL.n654 9.3005
R726 VTAIL.n706 VTAIL.n705 9.3005
R727 VTAIL.n708 VTAIL.n707 9.3005
R728 VTAIL.n650 VTAIL.n649 9.3005
R729 VTAIL.n714 VTAIL.n713 9.3005
R730 VTAIL.n716 VTAIL.n715 9.3005
R731 VTAIL.n739 VTAIL.n738 9.3005
R732 VTAIL.n638 VTAIL.n637 9.3005
R733 VTAIL.n733 VTAIL.n732 9.3005
R734 VTAIL.n731 VTAIL.n730 9.3005
R735 VTAIL.n642 VTAIL.n641 9.3005
R736 VTAIL.n725 VTAIL.n724 9.3005
R737 VTAIL.n723 VTAIL.n722 9.3005
R738 VTAIL.n646 VTAIL.n645 9.3005
R739 VTAIL.n659 VTAIL.n658 9.3005
R740 VTAIL.n692 VTAIL.n691 9.3005
R741 VTAIL.n690 VTAIL.n689 9.3005
R742 VTAIL.n663 VTAIL.n662 9.3005
R743 VTAIL.n684 VTAIL.n683 9.3005
R744 VTAIL.n682 VTAIL.n681 9.3005
R745 VTAIL.n667 VTAIL.n666 9.3005
R746 VTAIL.n676 VTAIL.n675 9.3005
R747 VTAIL.n674 VTAIL.n673 9.3005
R748 VTAIL.n592 VTAIL.n591 9.3005
R749 VTAIL.n594 VTAIL.n593 9.3005
R750 VTAIL.n549 VTAIL.n548 9.3005
R751 VTAIL.n600 VTAIL.n599 9.3005
R752 VTAIL.n602 VTAIL.n601 9.3005
R753 VTAIL.n544 VTAIL.n543 9.3005
R754 VTAIL.n608 VTAIL.n607 9.3005
R755 VTAIL.n610 VTAIL.n609 9.3005
R756 VTAIL.n633 VTAIL.n632 9.3005
R757 VTAIL.n532 VTAIL.n531 9.3005
R758 VTAIL.n627 VTAIL.n626 9.3005
R759 VTAIL.n625 VTAIL.n624 9.3005
R760 VTAIL.n536 VTAIL.n535 9.3005
R761 VTAIL.n619 VTAIL.n618 9.3005
R762 VTAIL.n617 VTAIL.n616 9.3005
R763 VTAIL.n540 VTAIL.n539 9.3005
R764 VTAIL.n553 VTAIL.n552 9.3005
R765 VTAIL.n586 VTAIL.n585 9.3005
R766 VTAIL.n584 VTAIL.n583 9.3005
R767 VTAIL.n557 VTAIL.n556 9.3005
R768 VTAIL.n578 VTAIL.n577 9.3005
R769 VTAIL.n576 VTAIL.n575 9.3005
R770 VTAIL.n561 VTAIL.n560 9.3005
R771 VTAIL.n570 VTAIL.n569 9.3005
R772 VTAIL.n568 VTAIL.n567 9.3005
R773 VTAIL.n486 VTAIL.n485 9.3005
R774 VTAIL.n488 VTAIL.n487 9.3005
R775 VTAIL.n443 VTAIL.n442 9.3005
R776 VTAIL.n494 VTAIL.n493 9.3005
R777 VTAIL.n496 VTAIL.n495 9.3005
R778 VTAIL.n438 VTAIL.n437 9.3005
R779 VTAIL.n502 VTAIL.n501 9.3005
R780 VTAIL.n504 VTAIL.n503 9.3005
R781 VTAIL.n527 VTAIL.n526 9.3005
R782 VTAIL.n426 VTAIL.n425 9.3005
R783 VTAIL.n521 VTAIL.n520 9.3005
R784 VTAIL.n519 VTAIL.n518 9.3005
R785 VTAIL.n430 VTAIL.n429 9.3005
R786 VTAIL.n513 VTAIL.n512 9.3005
R787 VTAIL.n511 VTAIL.n510 9.3005
R788 VTAIL.n434 VTAIL.n433 9.3005
R789 VTAIL.n447 VTAIL.n446 9.3005
R790 VTAIL.n480 VTAIL.n479 9.3005
R791 VTAIL.n478 VTAIL.n477 9.3005
R792 VTAIL.n451 VTAIL.n450 9.3005
R793 VTAIL.n472 VTAIL.n471 9.3005
R794 VTAIL.n470 VTAIL.n469 9.3005
R795 VTAIL.n455 VTAIL.n454 9.3005
R796 VTAIL.n464 VTAIL.n463 9.3005
R797 VTAIL.n462 VTAIL.n461 9.3005
R798 VTAIL.n380 VTAIL.n379 9.3005
R799 VTAIL.n382 VTAIL.n381 9.3005
R800 VTAIL.n337 VTAIL.n336 9.3005
R801 VTAIL.n388 VTAIL.n387 9.3005
R802 VTAIL.n390 VTAIL.n389 9.3005
R803 VTAIL.n332 VTAIL.n331 9.3005
R804 VTAIL.n396 VTAIL.n395 9.3005
R805 VTAIL.n398 VTAIL.n397 9.3005
R806 VTAIL.n421 VTAIL.n420 9.3005
R807 VTAIL.n320 VTAIL.n319 9.3005
R808 VTAIL.n415 VTAIL.n414 9.3005
R809 VTAIL.n413 VTAIL.n412 9.3005
R810 VTAIL.n324 VTAIL.n323 9.3005
R811 VTAIL.n407 VTAIL.n406 9.3005
R812 VTAIL.n405 VTAIL.n404 9.3005
R813 VTAIL.n328 VTAIL.n327 9.3005
R814 VTAIL.n341 VTAIL.n340 9.3005
R815 VTAIL.n374 VTAIL.n373 9.3005
R816 VTAIL.n372 VTAIL.n371 9.3005
R817 VTAIL.n345 VTAIL.n344 9.3005
R818 VTAIL.n366 VTAIL.n365 9.3005
R819 VTAIL.n364 VTAIL.n363 9.3005
R820 VTAIL.n349 VTAIL.n348 9.3005
R821 VTAIL.n358 VTAIL.n357 9.3005
R822 VTAIL.n356 VTAIL.n355 9.3005
R823 VTAIL.n793 VTAIL.n768 8.92171
R824 VTAIL.n806 VTAIL.n760 8.92171
R825 VTAIL.n840 VTAIL.n839 8.92171
R826 VTAIL.n51 VTAIL.n26 8.92171
R827 VTAIL.n64 VTAIL.n18 8.92171
R828 VTAIL.n98 VTAIL.n97 8.92171
R829 VTAIL.n157 VTAIL.n132 8.92171
R830 VTAIL.n170 VTAIL.n124 8.92171
R831 VTAIL.n204 VTAIL.n203 8.92171
R832 VTAIL.n263 VTAIL.n238 8.92171
R833 VTAIL.n276 VTAIL.n230 8.92171
R834 VTAIL.n310 VTAIL.n309 8.92171
R835 VTAIL.n734 VTAIL.n733 8.92171
R836 VTAIL.n701 VTAIL.n655 8.92171
R837 VTAIL.n688 VTAIL.n663 8.92171
R838 VTAIL.n628 VTAIL.n627 8.92171
R839 VTAIL.n595 VTAIL.n549 8.92171
R840 VTAIL.n582 VTAIL.n557 8.92171
R841 VTAIL.n522 VTAIL.n521 8.92171
R842 VTAIL.n489 VTAIL.n443 8.92171
R843 VTAIL.n476 VTAIL.n451 8.92171
R844 VTAIL.n416 VTAIL.n415 8.92171
R845 VTAIL.n383 VTAIL.n337 8.92171
R846 VTAIL.n370 VTAIL.n345 8.92171
R847 VTAIL.n794 VTAIL.n766 8.14595
R848 VTAIL.n805 VTAIL.n762 8.14595
R849 VTAIL.n843 VTAIL.n744 8.14595
R850 VTAIL.n52 VTAIL.n24 8.14595
R851 VTAIL.n63 VTAIL.n20 8.14595
R852 VTAIL.n101 VTAIL.n2 8.14595
R853 VTAIL.n158 VTAIL.n130 8.14595
R854 VTAIL.n169 VTAIL.n126 8.14595
R855 VTAIL.n207 VTAIL.n108 8.14595
R856 VTAIL.n264 VTAIL.n236 8.14595
R857 VTAIL.n275 VTAIL.n232 8.14595
R858 VTAIL.n313 VTAIL.n214 8.14595
R859 VTAIL.n737 VTAIL.n638 8.14595
R860 VTAIL.n700 VTAIL.n657 8.14595
R861 VTAIL.n689 VTAIL.n661 8.14595
R862 VTAIL.n631 VTAIL.n532 8.14595
R863 VTAIL.n594 VTAIL.n551 8.14595
R864 VTAIL.n583 VTAIL.n555 8.14595
R865 VTAIL.n525 VTAIL.n426 8.14595
R866 VTAIL.n488 VTAIL.n445 8.14595
R867 VTAIL.n477 VTAIL.n449 8.14595
R868 VTAIL.n419 VTAIL.n320 8.14595
R869 VTAIL.n382 VTAIL.n339 8.14595
R870 VTAIL.n371 VTAIL.n343 8.14595
R871 VTAIL.n798 VTAIL.n797 7.3702
R872 VTAIL.n802 VTAIL.n801 7.3702
R873 VTAIL.n844 VTAIL.n742 7.3702
R874 VTAIL.n56 VTAIL.n55 7.3702
R875 VTAIL.n60 VTAIL.n59 7.3702
R876 VTAIL.n102 VTAIL.n0 7.3702
R877 VTAIL.n162 VTAIL.n161 7.3702
R878 VTAIL.n166 VTAIL.n165 7.3702
R879 VTAIL.n208 VTAIL.n106 7.3702
R880 VTAIL.n268 VTAIL.n267 7.3702
R881 VTAIL.n272 VTAIL.n271 7.3702
R882 VTAIL.n314 VTAIL.n212 7.3702
R883 VTAIL.n738 VTAIL.n636 7.3702
R884 VTAIL.n697 VTAIL.n696 7.3702
R885 VTAIL.n693 VTAIL.n692 7.3702
R886 VTAIL.n632 VTAIL.n530 7.3702
R887 VTAIL.n591 VTAIL.n590 7.3702
R888 VTAIL.n587 VTAIL.n586 7.3702
R889 VTAIL.n526 VTAIL.n424 7.3702
R890 VTAIL.n485 VTAIL.n484 7.3702
R891 VTAIL.n481 VTAIL.n480 7.3702
R892 VTAIL.n420 VTAIL.n318 7.3702
R893 VTAIL.n379 VTAIL.n378 7.3702
R894 VTAIL.n375 VTAIL.n374 7.3702
R895 VTAIL.n798 VTAIL.n764 6.59444
R896 VTAIL.n801 VTAIL.n764 6.59444
R897 VTAIL.n846 VTAIL.n742 6.59444
R898 VTAIL.n56 VTAIL.n22 6.59444
R899 VTAIL.n59 VTAIL.n22 6.59444
R900 VTAIL.n104 VTAIL.n0 6.59444
R901 VTAIL.n162 VTAIL.n128 6.59444
R902 VTAIL.n165 VTAIL.n128 6.59444
R903 VTAIL.n210 VTAIL.n106 6.59444
R904 VTAIL.n268 VTAIL.n234 6.59444
R905 VTAIL.n271 VTAIL.n234 6.59444
R906 VTAIL.n316 VTAIL.n212 6.59444
R907 VTAIL.n740 VTAIL.n636 6.59444
R908 VTAIL.n696 VTAIL.n659 6.59444
R909 VTAIL.n693 VTAIL.n659 6.59444
R910 VTAIL.n634 VTAIL.n530 6.59444
R911 VTAIL.n590 VTAIL.n553 6.59444
R912 VTAIL.n587 VTAIL.n553 6.59444
R913 VTAIL.n528 VTAIL.n424 6.59444
R914 VTAIL.n484 VTAIL.n447 6.59444
R915 VTAIL.n481 VTAIL.n447 6.59444
R916 VTAIL.n422 VTAIL.n318 6.59444
R917 VTAIL.n378 VTAIL.n341 6.59444
R918 VTAIL.n375 VTAIL.n341 6.59444
R919 VTAIL.n797 VTAIL.n766 5.81868
R920 VTAIL.n802 VTAIL.n762 5.81868
R921 VTAIL.n844 VTAIL.n843 5.81868
R922 VTAIL.n55 VTAIL.n24 5.81868
R923 VTAIL.n60 VTAIL.n20 5.81868
R924 VTAIL.n102 VTAIL.n101 5.81868
R925 VTAIL.n161 VTAIL.n130 5.81868
R926 VTAIL.n166 VTAIL.n126 5.81868
R927 VTAIL.n208 VTAIL.n207 5.81868
R928 VTAIL.n267 VTAIL.n236 5.81868
R929 VTAIL.n272 VTAIL.n232 5.81868
R930 VTAIL.n314 VTAIL.n313 5.81868
R931 VTAIL.n738 VTAIL.n737 5.81868
R932 VTAIL.n697 VTAIL.n657 5.81868
R933 VTAIL.n692 VTAIL.n661 5.81868
R934 VTAIL.n632 VTAIL.n631 5.81868
R935 VTAIL.n591 VTAIL.n551 5.81868
R936 VTAIL.n586 VTAIL.n555 5.81868
R937 VTAIL.n526 VTAIL.n525 5.81868
R938 VTAIL.n485 VTAIL.n445 5.81868
R939 VTAIL.n480 VTAIL.n449 5.81868
R940 VTAIL.n420 VTAIL.n419 5.81868
R941 VTAIL.n379 VTAIL.n339 5.81868
R942 VTAIL.n374 VTAIL.n343 5.81868
R943 VTAIL.n794 VTAIL.n793 5.04292
R944 VTAIL.n806 VTAIL.n805 5.04292
R945 VTAIL.n840 VTAIL.n744 5.04292
R946 VTAIL.n52 VTAIL.n51 5.04292
R947 VTAIL.n64 VTAIL.n63 5.04292
R948 VTAIL.n98 VTAIL.n2 5.04292
R949 VTAIL.n158 VTAIL.n157 5.04292
R950 VTAIL.n170 VTAIL.n169 5.04292
R951 VTAIL.n204 VTAIL.n108 5.04292
R952 VTAIL.n264 VTAIL.n263 5.04292
R953 VTAIL.n276 VTAIL.n275 5.04292
R954 VTAIL.n310 VTAIL.n214 5.04292
R955 VTAIL.n734 VTAIL.n638 5.04292
R956 VTAIL.n701 VTAIL.n700 5.04292
R957 VTAIL.n689 VTAIL.n688 5.04292
R958 VTAIL.n628 VTAIL.n532 5.04292
R959 VTAIL.n595 VTAIL.n594 5.04292
R960 VTAIL.n583 VTAIL.n582 5.04292
R961 VTAIL.n522 VTAIL.n426 5.04292
R962 VTAIL.n489 VTAIL.n488 5.04292
R963 VTAIL.n477 VTAIL.n476 5.04292
R964 VTAIL.n416 VTAIL.n320 5.04292
R965 VTAIL.n383 VTAIL.n382 5.04292
R966 VTAIL.n371 VTAIL.n370 5.04292
R967 VTAIL.n790 VTAIL.n768 4.26717
R968 VTAIL.n809 VTAIL.n760 4.26717
R969 VTAIL.n839 VTAIL.n746 4.26717
R970 VTAIL.n48 VTAIL.n26 4.26717
R971 VTAIL.n67 VTAIL.n18 4.26717
R972 VTAIL.n97 VTAIL.n4 4.26717
R973 VTAIL.n154 VTAIL.n132 4.26717
R974 VTAIL.n173 VTAIL.n124 4.26717
R975 VTAIL.n203 VTAIL.n110 4.26717
R976 VTAIL.n260 VTAIL.n238 4.26717
R977 VTAIL.n279 VTAIL.n230 4.26717
R978 VTAIL.n309 VTAIL.n216 4.26717
R979 VTAIL.n733 VTAIL.n640 4.26717
R980 VTAIL.n704 VTAIL.n655 4.26717
R981 VTAIL.n685 VTAIL.n663 4.26717
R982 VTAIL.n627 VTAIL.n534 4.26717
R983 VTAIL.n598 VTAIL.n549 4.26717
R984 VTAIL.n579 VTAIL.n557 4.26717
R985 VTAIL.n521 VTAIL.n428 4.26717
R986 VTAIL.n492 VTAIL.n443 4.26717
R987 VTAIL.n473 VTAIL.n451 4.26717
R988 VTAIL.n415 VTAIL.n322 4.26717
R989 VTAIL.n386 VTAIL.n337 4.26717
R990 VTAIL.n367 VTAIL.n345 4.26717
R991 VTAIL.n779 VTAIL.n775 3.70982
R992 VTAIL.n37 VTAIL.n33 3.70982
R993 VTAIL.n143 VTAIL.n139 3.70982
R994 VTAIL.n249 VTAIL.n245 3.70982
R995 VTAIL.n674 VTAIL.n670 3.70982
R996 VTAIL.n568 VTAIL.n564 3.70982
R997 VTAIL.n462 VTAIL.n458 3.70982
R998 VTAIL.n356 VTAIL.n352 3.70982
R999 VTAIL.n789 VTAIL.n770 3.49141
R1000 VTAIL.n810 VTAIL.n758 3.49141
R1001 VTAIL.n836 VTAIL.n835 3.49141
R1002 VTAIL.n47 VTAIL.n28 3.49141
R1003 VTAIL.n68 VTAIL.n16 3.49141
R1004 VTAIL.n94 VTAIL.n93 3.49141
R1005 VTAIL.n153 VTAIL.n134 3.49141
R1006 VTAIL.n174 VTAIL.n122 3.49141
R1007 VTAIL.n200 VTAIL.n199 3.49141
R1008 VTAIL.n259 VTAIL.n240 3.49141
R1009 VTAIL.n280 VTAIL.n228 3.49141
R1010 VTAIL.n306 VTAIL.n305 3.49141
R1011 VTAIL.n730 VTAIL.n729 3.49141
R1012 VTAIL.n705 VTAIL.n653 3.49141
R1013 VTAIL.n684 VTAIL.n665 3.49141
R1014 VTAIL.n624 VTAIL.n623 3.49141
R1015 VTAIL.n599 VTAIL.n547 3.49141
R1016 VTAIL.n578 VTAIL.n559 3.49141
R1017 VTAIL.n518 VTAIL.n517 3.49141
R1018 VTAIL.n493 VTAIL.n441 3.49141
R1019 VTAIL.n472 VTAIL.n453 3.49141
R1020 VTAIL.n412 VTAIL.n411 3.49141
R1021 VTAIL.n387 VTAIL.n335 3.49141
R1022 VTAIL.n366 VTAIL.n347 3.49141
R1023 VTAIL.n529 VTAIL.n423 2.71602
R1024 VTAIL.n741 VTAIL.n635 2.71602
R1025 VTAIL.n317 VTAIL.n211 2.71602
R1026 VTAIL.n786 VTAIL.n785 2.71565
R1027 VTAIL.n814 VTAIL.n813 2.71565
R1028 VTAIL.n832 VTAIL.n748 2.71565
R1029 VTAIL.n44 VTAIL.n43 2.71565
R1030 VTAIL.n72 VTAIL.n71 2.71565
R1031 VTAIL.n90 VTAIL.n6 2.71565
R1032 VTAIL.n150 VTAIL.n149 2.71565
R1033 VTAIL.n178 VTAIL.n177 2.71565
R1034 VTAIL.n196 VTAIL.n112 2.71565
R1035 VTAIL.n256 VTAIL.n255 2.71565
R1036 VTAIL.n284 VTAIL.n283 2.71565
R1037 VTAIL.n302 VTAIL.n218 2.71565
R1038 VTAIL.n726 VTAIL.n642 2.71565
R1039 VTAIL.n709 VTAIL.n708 2.71565
R1040 VTAIL.n681 VTAIL.n680 2.71565
R1041 VTAIL.n620 VTAIL.n536 2.71565
R1042 VTAIL.n603 VTAIL.n602 2.71565
R1043 VTAIL.n575 VTAIL.n574 2.71565
R1044 VTAIL.n514 VTAIL.n430 2.71565
R1045 VTAIL.n497 VTAIL.n496 2.71565
R1046 VTAIL.n469 VTAIL.n468 2.71565
R1047 VTAIL.n408 VTAIL.n324 2.71565
R1048 VTAIL.n391 VTAIL.n390 2.71565
R1049 VTAIL.n363 VTAIL.n362 2.71565
R1050 VTAIL.n782 VTAIL.n772 1.93989
R1051 VTAIL.n818 VTAIL.n756 1.93989
R1052 VTAIL.n831 VTAIL.n750 1.93989
R1053 VTAIL.n40 VTAIL.n30 1.93989
R1054 VTAIL.n76 VTAIL.n14 1.93989
R1055 VTAIL.n89 VTAIL.n8 1.93989
R1056 VTAIL.n146 VTAIL.n136 1.93989
R1057 VTAIL.n182 VTAIL.n120 1.93989
R1058 VTAIL.n195 VTAIL.n114 1.93989
R1059 VTAIL.n252 VTAIL.n242 1.93989
R1060 VTAIL.n288 VTAIL.n226 1.93989
R1061 VTAIL.n301 VTAIL.n220 1.93989
R1062 VTAIL.n725 VTAIL.n644 1.93989
R1063 VTAIL.n712 VTAIL.n650 1.93989
R1064 VTAIL.n677 VTAIL.n667 1.93989
R1065 VTAIL.n619 VTAIL.n538 1.93989
R1066 VTAIL.n606 VTAIL.n544 1.93989
R1067 VTAIL.n571 VTAIL.n561 1.93989
R1068 VTAIL.n513 VTAIL.n432 1.93989
R1069 VTAIL.n500 VTAIL.n438 1.93989
R1070 VTAIL.n465 VTAIL.n455 1.93989
R1071 VTAIL.n407 VTAIL.n326 1.93989
R1072 VTAIL.n394 VTAIL.n332 1.93989
R1073 VTAIL.n359 VTAIL.n349 1.93989
R1074 VTAIL VTAIL.n105 1.41645
R1075 VTAIL VTAIL.n847 1.30007
R1076 VTAIL.n781 VTAIL.n774 1.16414
R1077 VTAIL.n819 VTAIL.n754 1.16414
R1078 VTAIL.n828 VTAIL.n827 1.16414
R1079 VTAIL.n39 VTAIL.n32 1.16414
R1080 VTAIL.n77 VTAIL.n12 1.16414
R1081 VTAIL.n86 VTAIL.n85 1.16414
R1082 VTAIL.n145 VTAIL.n138 1.16414
R1083 VTAIL.n183 VTAIL.n118 1.16414
R1084 VTAIL.n192 VTAIL.n191 1.16414
R1085 VTAIL.n251 VTAIL.n244 1.16414
R1086 VTAIL.n289 VTAIL.n224 1.16414
R1087 VTAIL.n298 VTAIL.n297 1.16414
R1088 VTAIL.n722 VTAIL.n721 1.16414
R1089 VTAIL.n713 VTAIL.n648 1.16414
R1090 VTAIL.n676 VTAIL.n669 1.16414
R1091 VTAIL.n616 VTAIL.n615 1.16414
R1092 VTAIL.n607 VTAIL.n542 1.16414
R1093 VTAIL.n570 VTAIL.n563 1.16414
R1094 VTAIL.n510 VTAIL.n509 1.16414
R1095 VTAIL.n501 VTAIL.n436 1.16414
R1096 VTAIL.n464 VTAIL.n457 1.16414
R1097 VTAIL.n404 VTAIL.n403 1.16414
R1098 VTAIL.n395 VTAIL.n330 1.16414
R1099 VTAIL.n358 VTAIL.n351 1.16414
R1100 VTAIL.n635 VTAIL.n529 0.470328
R1101 VTAIL.n211 VTAIL.n105 0.470328
R1102 VTAIL.n778 VTAIL.n777 0.388379
R1103 VTAIL.n823 VTAIL.n822 0.388379
R1104 VTAIL.n824 VTAIL.n752 0.388379
R1105 VTAIL.n36 VTAIL.n35 0.388379
R1106 VTAIL.n81 VTAIL.n80 0.388379
R1107 VTAIL.n82 VTAIL.n10 0.388379
R1108 VTAIL.n142 VTAIL.n141 0.388379
R1109 VTAIL.n187 VTAIL.n186 0.388379
R1110 VTAIL.n188 VTAIL.n116 0.388379
R1111 VTAIL.n248 VTAIL.n247 0.388379
R1112 VTAIL.n293 VTAIL.n292 0.388379
R1113 VTAIL.n294 VTAIL.n222 0.388379
R1114 VTAIL.n718 VTAIL.n646 0.388379
R1115 VTAIL.n717 VTAIL.n716 0.388379
R1116 VTAIL.n673 VTAIL.n672 0.388379
R1117 VTAIL.n612 VTAIL.n540 0.388379
R1118 VTAIL.n611 VTAIL.n610 0.388379
R1119 VTAIL.n567 VTAIL.n566 0.388379
R1120 VTAIL.n506 VTAIL.n434 0.388379
R1121 VTAIL.n505 VTAIL.n504 0.388379
R1122 VTAIL.n461 VTAIL.n460 0.388379
R1123 VTAIL.n400 VTAIL.n328 0.388379
R1124 VTAIL.n399 VTAIL.n398 0.388379
R1125 VTAIL.n355 VTAIL.n354 0.388379
R1126 VTAIL.n780 VTAIL.n779 0.155672
R1127 VTAIL.n780 VTAIL.n771 0.155672
R1128 VTAIL.n787 VTAIL.n771 0.155672
R1129 VTAIL.n788 VTAIL.n787 0.155672
R1130 VTAIL.n788 VTAIL.n767 0.155672
R1131 VTAIL.n795 VTAIL.n767 0.155672
R1132 VTAIL.n796 VTAIL.n795 0.155672
R1133 VTAIL.n796 VTAIL.n763 0.155672
R1134 VTAIL.n803 VTAIL.n763 0.155672
R1135 VTAIL.n804 VTAIL.n803 0.155672
R1136 VTAIL.n804 VTAIL.n759 0.155672
R1137 VTAIL.n811 VTAIL.n759 0.155672
R1138 VTAIL.n812 VTAIL.n811 0.155672
R1139 VTAIL.n812 VTAIL.n755 0.155672
R1140 VTAIL.n820 VTAIL.n755 0.155672
R1141 VTAIL.n821 VTAIL.n820 0.155672
R1142 VTAIL.n821 VTAIL.n751 0.155672
R1143 VTAIL.n829 VTAIL.n751 0.155672
R1144 VTAIL.n830 VTAIL.n829 0.155672
R1145 VTAIL.n830 VTAIL.n747 0.155672
R1146 VTAIL.n837 VTAIL.n747 0.155672
R1147 VTAIL.n838 VTAIL.n837 0.155672
R1148 VTAIL.n838 VTAIL.n743 0.155672
R1149 VTAIL.n845 VTAIL.n743 0.155672
R1150 VTAIL.n38 VTAIL.n37 0.155672
R1151 VTAIL.n38 VTAIL.n29 0.155672
R1152 VTAIL.n45 VTAIL.n29 0.155672
R1153 VTAIL.n46 VTAIL.n45 0.155672
R1154 VTAIL.n46 VTAIL.n25 0.155672
R1155 VTAIL.n53 VTAIL.n25 0.155672
R1156 VTAIL.n54 VTAIL.n53 0.155672
R1157 VTAIL.n54 VTAIL.n21 0.155672
R1158 VTAIL.n61 VTAIL.n21 0.155672
R1159 VTAIL.n62 VTAIL.n61 0.155672
R1160 VTAIL.n62 VTAIL.n17 0.155672
R1161 VTAIL.n69 VTAIL.n17 0.155672
R1162 VTAIL.n70 VTAIL.n69 0.155672
R1163 VTAIL.n70 VTAIL.n13 0.155672
R1164 VTAIL.n78 VTAIL.n13 0.155672
R1165 VTAIL.n79 VTAIL.n78 0.155672
R1166 VTAIL.n79 VTAIL.n9 0.155672
R1167 VTAIL.n87 VTAIL.n9 0.155672
R1168 VTAIL.n88 VTAIL.n87 0.155672
R1169 VTAIL.n88 VTAIL.n5 0.155672
R1170 VTAIL.n95 VTAIL.n5 0.155672
R1171 VTAIL.n96 VTAIL.n95 0.155672
R1172 VTAIL.n96 VTAIL.n1 0.155672
R1173 VTAIL.n103 VTAIL.n1 0.155672
R1174 VTAIL.n144 VTAIL.n143 0.155672
R1175 VTAIL.n144 VTAIL.n135 0.155672
R1176 VTAIL.n151 VTAIL.n135 0.155672
R1177 VTAIL.n152 VTAIL.n151 0.155672
R1178 VTAIL.n152 VTAIL.n131 0.155672
R1179 VTAIL.n159 VTAIL.n131 0.155672
R1180 VTAIL.n160 VTAIL.n159 0.155672
R1181 VTAIL.n160 VTAIL.n127 0.155672
R1182 VTAIL.n167 VTAIL.n127 0.155672
R1183 VTAIL.n168 VTAIL.n167 0.155672
R1184 VTAIL.n168 VTAIL.n123 0.155672
R1185 VTAIL.n175 VTAIL.n123 0.155672
R1186 VTAIL.n176 VTAIL.n175 0.155672
R1187 VTAIL.n176 VTAIL.n119 0.155672
R1188 VTAIL.n184 VTAIL.n119 0.155672
R1189 VTAIL.n185 VTAIL.n184 0.155672
R1190 VTAIL.n185 VTAIL.n115 0.155672
R1191 VTAIL.n193 VTAIL.n115 0.155672
R1192 VTAIL.n194 VTAIL.n193 0.155672
R1193 VTAIL.n194 VTAIL.n111 0.155672
R1194 VTAIL.n201 VTAIL.n111 0.155672
R1195 VTAIL.n202 VTAIL.n201 0.155672
R1196 VTAIL.n202 VTAIL.n107 0.155672
R1197 VTAIL.n209 VTAIL.n107 0.155672
R1198 VTAIL.n250 VTAIL.n249 0.155672
R1199 VTAIL.n250 VTAIL.n241 0.155672
R1200 VTAIL.n257 VTAIL.n241 0.155672
R1201 VTAIL.n258 VTAIL.n257 0.155672
R1202 VTAIL.n258 VTAIL.n237 0.155672
R1203 VTAIL.n265 VTAIL.n237 0.155672
R1204 VTAIL.n266 VTAIL.n265 0.155672
R1205 VTAIL.n266 VTAIL.n233 0.155672
R1206 VTAIL.n273 VTAIL.n233 0.155672
R1207 VTAIL.n274 VTAIL.n273 0.155672
R1208 VTAIL.n274 VTAIL.n229 0.155672
R1209 VTAIL.n281 VTAIL.n229 0.155672
R1210 VTAIL.n282 VTAIL.n281 0.155672
R1211 VTAIL.n282 VTAIL.n225 0.155672
R1212 VTAIL.n290 VTAIL.n225 0.155672
R1213 VTAIL.n291 VTAIL.n290 0.155672
R1214 VTAIL.n291 VTAIL.n221 0.155672
R1215 VTAIL.n299 VTAIL.n221 0.155672
R1216 VTAIL.n300 VTAIL.n299 0.155672
R1217 VTAIL.n300 VTAIL.n217 0.155672
R1218 VTAIL.n307 VTAIL.n217 0.155672
R1219 VTAIL.n308 VTAIL.n307 0.155672
R1220 VTAIL.n308 VTAIL.n213 0.155672
R1221 VTAIL.n315 VTAIL.n213 0.155672
R1222 VTAIL.n739 VTAIL.n637 0.155672
R1223 VTAIL.n732 VTAIL.n637 0.155672
R1224 VTAIL.n732 VTAIL.n731 0.155672
R1225 VTAIL.n731 VTAIL.n641 0.155672
R1226 VTAIL.n724 VTAIL.n641 0.155672
R1227 VTAIL.n724 VTAIL.n723 0.155672
R1228 VTAIL.n723 VTAIL.n645 0.155672
R1229 VTAIL.n715 VTAIL.n645 0.155672
R1230 VTAIL.n715 VTAIL.n714 0.155672
R1231 VTAIL.n714 VTAIL.n649 0.155672
R1232 VTAIL.n707 VTAIL.n649 0.155672
R1233 VTAIL.n707 VTAIL.n706 0.155672
R1234 VTAIL.n706 VTAIL.n654 0.155672
R1235 VTAIL.n699 VTAIL.n654 0.155672
R1236 VTAIL.n699 VTAIL.n698 0.155672
R1237 VTAIL.n698 VTAIL.n658 0.155672
R1238 VTAIL.n691 VTAIL.n658 0.155672
R1239 VTAIL.n691 VTAIL.n690 0.155672
R1240 VTAIL.n690 VTAIL.n662 0.155672
R1241 VTAIL.n683 VTAIL.n662 0.155672
R1242 VTAIL.n683 VTAIL.n682 0.155672
R1243 VTAIL.n682 VTAIL.n666 0.155672
R1244 VTAIL.n675 VTAIL.n666 0.155672
R1245 VTAIL.n675 VTAIL.n674 0.155672
R1246 VTAIL.n633 VTAIL.n531 0.155672
R1247 VTAIL.n626 VTAIL.n531 0.155672
R1248 VTAIL.n626 VTAIL.n625 0.155672
R1249 VTAIL.n625 VTAIL.n535 0.155672
R1250 VTAIL.n618 VTAIL.n535 0.155672
R1251 VTAIL.n618 VTAIL.n617 0.155672
R1252 VTAIL.n617 VTAIL.n539 0.155672
R1253 VTAIL.n609 VTAIL.n539 0.155672
R1254 VTAIL.n609 VTAIL.n608 0.155672
R1255 VTAIL.n608 VTAIL.n543 0.155672
R1256 VTAIL.n601 VTAIL.n543 0.155672
R1257 VTAIL.n601 VTAIL.n600 0.155672
R1258 VTAIL.n600 VTAIL.n548 0.155672
R1259 VTAIL.n593 VTAIL.n548 0.155672
R1260 VTAIL.n593 VTAIL.n592 0.155672
R1261 VTAIL.n592 VTAIL.n552 0.155672
R1262 VTAIL.n585 VTAIL.n552 0.155672
R1263 VTAIL.n585 VTAIL.n584 0.155672
R1264 VTAIL.n584 VTAIL.n556 0.155672
R1265 VTAIL.n577 VTAIL.n556 0.155672
R1266 VTAIL.n577 VTAIL.n576 0.155672
R1267 VTAIL.n576 VTAIL.n560 0.155672
R1268 VTAIL.n569 VTAIL.n560 0.155672
R1269 VTAIL.n569 VTAIL.n568 0.155672
R1270 VTAIL.n527 VTAIL.n425 0.155672
R1271 VTAIL.n520 VTAIL.n425 0.155672
R1272 VTAIL.n520 VTAIL.n519 0.155672
R1273 VTAIL.n519 VTAIL.n429 0.155672
R1274 VTAIL.n512 VTAIL.n429 0.155672
R1275 VTAIL.n512 VTAIL.n511 0.155672
R1276 VTAIL.n511 VTAIL.n433 0.155672
R1277 VTAIL.n503 VTAIL.n433 0.155672
R1278 VTAIL.n503 VTAIL.n502 0.155672
R1279 VTAIL.n502 VTAIL.n437 0.155672
R1280 VTAIL.n495 VTAIL.n437 0.155672
R1281 VTAIL.n495 VTAIL.n494 0.155672
R1282 VTAIL.n494 VTAIL.n442 0.155672
R1283 VTAIL.n487 VTAIL.n442 0.155672
R1284 VTAIL.n487 VTAIL.n486 0.155672
R1285 VTAIL.n486 VTAIL.n446 0.155672
R1286 VTAIL.n479 VTAIL.n446 0.155672
R1287 VTAIL.n479 VTAIL.n478 0.155672
R1288 VTAIL.n478 VTAIL.n450 0.155672
R1289 VTAIL.n471 VTAIL.n450 0.155672
R1290 VTAIL.n471 VTAIL.n470 0.155672
R1291 VTAIL.n470 VTAIL.n454 0.155672
R1292 VTAIL.n463 VTAIL.n454 0.155672
R1293 VTAIL.n463 VTAIL.n462 0.155672
R1294 VTAIL.n421 VTAIL.n319 0.155672
R1295 VTAIL.n414 VTAIL.n319 0.155672
R1296 VTAIL.n414 VTAIL.n413 0.155672
R1297 VTAIL.n413 VTAIL.n323 0.155672
R1298 VTAIL.n406 VTAIL.n323 0.155672
R1299 VTAIL.n406 VTAIL.n405 0.155672
R1300 VTAIL.n405 VTAIL.n327 0.155672
R1301 VTAIL.n397 VTAIL.n327 0.155672
R1302 VTAIL.n397 VTAIL.n396 0.155672
R1303 VTAIL.n396 VTAIL.n331 0.155672
R1304 VTAIL.n389 VTAIL.n331 0.155672
R1305 VTAIL.n389 VTAIL.n388 0.155672
R1306 VTAIL.n388 VTAIL.n336 0.155672
R1307 VTAIL.n381 VTAIL.n336 0.155672
R1308 VTAIL.n381 VTAIL.n380 0.155672
R1309 VTAIL.n380 VTAIL.n340 0.155672
R1310 VTAIL.n373 VTAIL.n340 0.155672
R1311 VTAIL.n373 VTAIL.n372 0.155672
R1312 VTAIL.n372 VTAIL.n344 0.155672
R1313 VTAIL.n365 VTAIL.n344 0.155672
R1314 VTAIL.n365 VTAIL.n364 0.155672
R1315 VTAIL.n364 VTAIL.n348 0.155672
R1316 VTAIL.n357 VTAIL.n348 0.155672
R1317 VTAIL.n357 VTAIL.n356 0.155672
R1318 B.n582 B.n91 585
R1319 B.n584 B.n583 585
R1320 B.n585 B.n90 585
R1321 B.n587 B.n586 585
R1322 B.n588 B.n89 585
R1323 B.n590 B.n589 585
R1324 B.n591 B.n88 585
R1325 B.n593 B.n592 585
R1326 B.n594 B.n87 585
R1327 B.n596 B.n595 585
R1328 B.n597 B.n86 585
R1329 B.n599 B.n598 585
R1330 B.n600 B.n85 585
R1331 B.n602 B.n601 585
R1332 B.n603 B.n84 585
R1333 B.n605 B.n604 585
R1334 B.n606 B.n83 585
R1335 B.n608 B.n607 585
R1336 B.n609 B.n82 585
R1337 B.n611 B.n610 585
R1338 B.n612 B.n81 585
R1339 B.n614 B.n613 585
R1340 B.n615 B.n80 585
R1341 B.n617 B.n616 585
R1342 B.n618 B.n79 585
R1343 B.n620 B.n619 585
R1344 B.n621 B.n78 585
R1345 B.n623 B.n622 585
R1346 B.n624 B.n77 585
R1347 B.n626 B.n625 585
R1348 B.n627 B.n76 585
R1349 B.n629 B.n628 585
R1350 B.n630 B.n75 585
R1351 B.n632 B.n631 585
R1352 B.n633 B.n74 585
R1353 B.n635 B.n634 585
R1354 B.n636 B.n73 585
R1355 B.n638 B.n637 585
R1356 B.n639 B.n72 585
R1357 B.n641 B.n640 585
R1358 B.n642 B.n71 585
R1359 B.n644 B.n643 585
R1360 B.n645 B.n70 585
R1361 B.n647 B.n646 585
R1362 B.n648 B.n69 585
R1363 B.n650 B.n649 585
R1364 B.n651 B.n68 585
R1365 B.n653 B.n652 585
R1366 B.n654 B.n67 585
R1367 B.n656 B.n655 585
R1368 B.n657 B.n66 585
R1369 B.n659 B.n658 585
R1370 B.n660 B.n65 585
R1371 B.n662 B.n661 585
R1372 B.n663 B.n64 585
R1373 B.n665 B.n664 585
R1374 B.n666 B.n63 585
R1375 B.n668 B.n667 585
R1376 B.n669 B.n62 585
R1377 B.n671 B.n670 585
R1378 B.n672 B.n61 585
R1379 B.n674 B.n673 585
R1380 B.n676 B.n675 585
R1381 B.n677 B.n57 585
R1382 B.n679 B.n678 585
R1383 B.n680 B.n56 585
R1384 B.n682 B.n681 585
R1385 B.n683 B.n55 585
R1386 B.n685 B.n684 585
R1387 B.n686 B.n54 585
R1388 B.n688 B.n687 585
R1389 B.n689 B.n51 585
R1390 B.n692 B.n691 585
R1391 B.n693 B.n50 585
R1392 B.n695 B.n694 585
R1393 B.n696 B.n49 585
R1394 B.n698 B.n697 585
R1395 B.n699 B.n48 585
R1396 B.n701 B.n700 585
R1397 B.n702 B.n47 585
R1398 B.n704 B.n703 585
R1399 B.n705 B.n46 585
R1400 B.n707 B.n706 585
R1401 B.n708 B.n45 585
R1402 B.n710 B.n709 585
R1403 B.n711 B.n44 585
R1404 B.n713 B.n712 585
R1405 B.n714 B.n43 585
R1406 B.n716 B.n715 585
R1407 B.n717 B.n42 585
R1408 B.n719 B.n718 585
R1409 B.n720 B.n41 585
R1410 B.n722 B.n721 585
R1411 B.n723 B.n40 585
R1412 B.n725 B.n724 585
R1413 B.n726 B.n39 585
R1414 B.n728 B.n727 585
R1415 B.n729 B.n38 585
R1416 B.n731 B.n730 585
R1417 B.n732 B.n37 585
R1418 B.n734 B.n733 585
R1419 B.n735 B.n36 585
R1420 B.n737 B.n736 585
R1421 B.n738 B.n35 585
R1422 B.n740 B.n739 585
R1423 B.n741 B.n34 585
R1424 B.n743 B.n742 585
R1425 B.n744 B.n33 585
R1426 B.n746 B.n745 585
R1427 B.n747 B.n32 585
R1428 B.n749 B.n748 585
R1429 B.n750 B.n31 585
R1430 B.n752 B.n751 585
R1431 B.n753 B.n30 585
R1432 B.n755 B.n754 585
R1433 B.n756 B.n29 585
R1434 B.n758 B.n757 585
R1435 B.n759 B.n28 585
R1436 B.n761 B.n760 585
R1437 B.n762 B.n27 585
R1438 B.n764 B.n763 585
R1439 B.n765 B.n26 585
R1440 B.n767 B.n766 585
R1441 B.n768 B.n25 585
R1442 B.n770 B.n769 585
R1443 B.n771 B.n24 585
R1444 B.n773 B.n772 585
R1445 B.n774 B.n23 585
R1446 B.n776 B.n775 585
R1447 B.n777 B.n22 585
R1448 B.n779 B.n778 585
R1449 B.n780 B.n21 585
R1450 B.n782 B.n781 585
R1451 B.n783 B.n20 585
R1452 B.n581 B.n580 585
R1453 B.n579 B.n92 585
R1454 B.n578 B.n577 585
R1455 B.n576 B.n93 585
R1456 B.n575 B.n574 585
R1457 B.n573 B.n94 585
R1458 B.n572 B.n571 585
R1459 B.n570 B.n95 585
R1460 B.n569 B.n568 585
R1461 B.n567 B.n96 585
R1462 B.n566 B.n565 585
R1463 B.n564 B.n97 585
R1464 B.n563 B.n562 585
R1465 B.n561 B.n98 585
R1466 B.n560 B.n559 585
R1467 B.n558 B.n99 585
R1468 B.n557 B.n556 585
R1469 B.n555 B.n100 585
R1470 B.n554 B.n553 585
R1471 B.n552 B.n101 585
R1472 B.n551 B.n550 585
R1473 B.n549 B.n102 585
R1474 B.n548 B.n547 585
R1475 B.n546 B.n103 585
R1476 B.n545 B.n544 585
R1477 B.n543 B.n104 585
R1478 B.n542 B.n541 585
R1479 B.n540 B.n105 585
R1480 B.n539 B.n538 585
R1481 B.n537 B.n106 585
R1482 B.n536 B.n535 585
R1483 B.n534 B.n107 585
R1484 B.n533 B.n532 585
R1485 B.n531 B.n108 585
R1486 B.n530 B.n529 585
R1487 B.n528 B.n109 585
R1488 B.n527 B.n526 585
R1489 B.n525 B.n110 585
R1490 B.n524 B.n523 585
R1491 B.n522 B.n111 585
R1492 B.n521 B.n520 585
R1493 B.n519 B.n112 585
R1494 B.n518 B.n517 585
R1495 B.n516 B.n113 585
R1496 B.n515 B.n514 585
R1497 B.n513 B.n114 585
R1498 B.n512 B.n511 585
R1499 B.n510 B.n115 585
R1500 B.n509 B.n508 585
R1501 B.n507 B.n116 585
R1502 B.n506 B.n505 585
R1503 B.n504 B.n117 585
R1504 B.n503 B.n502 585
R1505 B.n501 B.n118 585
R1506 B.n500 B.n499 585
R1507 B.n498 B.n119 585
R1508 B.n497 B.n496 585
R1509 B.n495 B.n120 585
R1510 B.n494 B.n493 585
R1511 B.n492 B.n121 585
R1512 B.n491 B.n490 585
R1513 B.n489 B.n122 585
R1514 B.n488 B.n487 585
R1515 B.n486 B.n123 585
R1516 B.n485 B.n484 585
R1517 B.n483 B.n124 585
R1518 B.n482 B.n481 585
R1519 B.n480 B.n125 585
R1520 B.n479 B.n478 585
R1521 B.n477 B.n126 585
R1522 B.n476 B.n475 585
R1523 B.n474 B.n127 585
R1524 B.n473 B.n472 585
R1525 B.n270 B.n199 585
R1526 B.n272 B.n271 585
R1527 B.n273 B.n198 585
R1528 B.n275 B.n274 585
R1529 B.n276 B.n197 585
R1530 B.n278 B.n277 585
R1531 B.n279 B.n196 585
R1532 B.n281 B.n280 585
R1533 B.n282 B.n195 585
R1534 B.n284 B.n283 585
R1535 B.n285 B.n194 585
R1536 B.n287 B.n286 585
R1537 B.n288 B.n193 585
R1538 B.n290 B.n289 585
R1539 B.n291 B.n192 585
R1540 B.n293 B.n292 585
R1541 B.n294 B.n191 585
R1542 B.n296 B.n295 585
R1543 B.n297 B.n190 585
R1544 B.n299 B.n298 585
R1545 B.n300 B.n189 585
R1546 B.n302 B.n301 585
R1547 B.n303 B.n188 585
R1548 B.n305 B.n304 585
R1549 B.n306 B.n187 585
R1550 B.n308 B.n307 585
R1551 B.n309 B.n186 585
R1552 B.n311 B.n310 585
R1553 B.n312 B.n185 585
R1554 B.n314 B.n313 585
R1555 B.n315 B.n184 585
R1556 B.n317 B.n316 585
R1557 B.n318 B.n183 585
R1558 B.n320 B.n319 585
R1559 B.n321 B.n182 585
R1560 B.n323 B.n322 585
R1561 B.n324 B.n181 585
R1562 B.n326 B.n325 585
R1563 B.n327 B.n180 585
R1564 B.n329 B.n328 585
R1565 B.n330 B.n179 585
R1566 B.n332 B.n331 585
R1567 B.n333 B.n178 585
R1568 B.n335 B.n334 585
R1569 B.n336 B.n177 585
R1570 B.n338 B.n337 585
R1571 B.n339 B.n176 585
R1572 B.n341 B.n340 585
R1573 B.n342 B.n175 585
R1574 B.n344 B.n343 585
R1575 B.n345 B.n174 585
R1576 B.n347 B.n346 585
R1577 B.n348 B.n173 585
R1578 B.n350 B.n349 585
R1579 B.n351 B.n172 585
R1580 B.n353 B.n352 585
R1581 B.n354 B.n171 585
R1582 B.n356 B.n355 585
R1583 B.n357 B.n170 585
R1584 B.n359 B.n358 585
R1585 B.n360 B.n169 585
R1586 B.n362 B.n361 585
R1587 B.n364 B.n363 585
R1588 B.n365 B.n165 585
R1589 B.n367 B.n366 585
R1590 B.n368 B.n164 585
R1591 B.n370 B.n369 585
R1592 B.n371 B.n163 585
R1593 B.n373 B.n372 585
R1594 B.n374 B.n162 585
R1595 B.n376 B.n375 585
R1596 B.n377 B.n159 585
R1597 B.n380 B.n379 585
R1598 B.n381 B.n158 585
R1599 B.n383 B.n382 585
R1600 B.n384 B.n157 585
R1601 B.n386 B.n385 585
R1602 B.n387 B.n156 585
R1603 B.n389 B.n388 585
R1604 B.n390 B.n155 585
R1605 B.n392 B.n391 585
R1606 B.n393 B.n154 585
R1607 B.n395 B.n394 585
R1608 B.n396 B.n153 585
R1609 B.n398 B.n397 585
R1610 B.n399 B.n152 585
R1611 B.n401 B.n400 585
R1612 B.n402 B.n151 585
R1613 B.n404 B.n403 585
R1614 B.n405 B.n150 585
R1615 B.n407 B.n406 585
R1616 B.n408 B.n149 585
R1617 B.n410 B.n409 585
R1618 B.n411 B.n148 585
R1619 B.n413 B.n412 585
R1620 B.n414 B.n147 585
R1621 B.n416 B.n415 585
R1622 B.n417 B.n146 585
R1623 B.n419 B.n418 585
R1624 B.n420 B.n145 585
R1625 B.n422 B.n421 585
R1626 B.n423 B.n144 585
R1627 B.n425 B.n424 585
R1628 B.n426 B.n143 585
R1629 B.n428 B.n427 585
R1630 B.n429 B.n142 585
R1631 B.n431 B.n430 585
R1632 B.n432 B.n141 585
R1633 B.n434 B.n433 585
R1634 B.n435 B.n140 585
R1635 B.n437 B.n436 585
R1636 B.n438 B.n139 585
R1637 B.n440 B.n439 585
R1638 B.n441 B.n138 585
R1639 B.n443 B.n442 585
R1640 B.n444 B.n137 585
R1641 B.n446 B.n445 585
R1642 B.n447 B.n136 585
R1643 B.n449 B.n448 585
R1644 B.n450 B.n135 585
R1645 B.n452 B.n451 585
R1646 B.n453 B.n134 585
R1647 B.n455 B.n454 585
R1648 B.n456 B.n133 585
R1649 B.n458 B.n457 585
R1650 B.n459 B.n132 585
R1651 B.n461 B.n460 585
R1652 B.n462 B.n131 585
R1653 B.n464 B.n463 585
R1654 B.n465 B.n130 585
R1655 B.n467 B.n466 585
R1656 B.n468 B.n129 585
R1657 B.n470 B.n469 585
R1658 B.n471 B.n128 585
R1659 B.n269 B.n268 585
R1660 B.n267 B.n200 585
R1661 B.n266 B.n265 585
R1662 B.n264 B.n201 585
R1663 B.n263 B.n262 585
R1664 B.n261 B.n202 585
R1665 B.n260 B.n259 585
R1666 B.n258 B.n203 585
R1667 B.n257 B.n256 585
R1668 B.n255 B.n204 585
R1669 B.n254 B.n253 585
R1670 B.n252 B.n205 585
R1671 B.n251 B.n250 585
R1672 B.n249 B.n206 585
R1673 B.n248 B.n247 585
R1674 B.n246 B.n207 585
R1675 B.n245 B.n244 585
R1676 B.n243 B.n208 585
R1677 B.n242 B.n241 585
R1678 B.n240 B.n209 585
R1679 B.n239 B.n238 585
R1680 B.n237 B.n210 585
R1681 B.n236 B.n235 585
R1682 B.n234 B.n211 585
R1683 B.n233 B.n232 585
R1684 B.n231 B.n212 585
R1685 B.n230 B.n229 585
R1686 B.n228 B.n213 585
R1687 B.n227 B.n226 585
R1688 B.n225 B.n214 585
R1689 B.n224 B.n223 585
R1690 B.n222 B.n215 585
R1691 B.n221 B.n220 585
R1692 B.n219 B.n216 585
R1693 B.n218 B.n217 585
R1694 B.n2 B.n0 585
R1695 B.n837 B.n1 585
R1696 B.n836 B.n835 585
R1697 B.n834 B.n3 585
R1698 B.n833 B.n832 585
R1699 B.n831 B.n4 585
R1700 B.n830 B.n829 585
R1701 B.n828 B.n5 585
R1702 B.n827 B.n826 585
R1703 B.n825 B.n6 585
R1704 B.n824 B.n823 585
R1705 B.n822 B.n7 585
R1706 B.n821 B.n820 585
R1707 B.n819 B.n8 585
R1708 B.n818 B.n817 585
R1709 B.n816 B.n9 585
R1710 B.n815 B.n814 585
R1711 B.n813 B.n10 585
R1712 B.n812 B.n811 585
R1713 B.n810 B.n11 585
R1714 B.n809 B.n808 585
R1715 B.n807 B.n12 585
R1716 B.n806 B.n805 585
R1717 B.n804 B.n13 585
R1718 B.n803 B.n802 585
R1719 B.n801 B.n14 585
R1720 B.n800 B.n799 585
R1721 B.n798 B.n15 585
R1722 B.n797 B.n796 585
R1723 B.n795 B.n16 585
R1724 B.n794 B.n793 585
R1725 B.n792 B.n17 585
R1726 B.n791 B.n790 585
R1727 B.n789 B.n18 585
R1728 B.n788 B.n787 585
R1729 B.n786 B.n19 585
R1730 B.n785 B.n784 585
R1731 B.n839 B.n838 585
R1732 B.n160 B.t2 561.622
R1733 B.n58 B.t10 561.622
R1734 B.n166 B.t8 561.622
R1735 B.n52 B.t4 561.622
R1736 B.n161 B.t1 500.531
R1737 B.n59 B.t11 500.531
R1738 B.n167 B.t7 500.531
R1739 B.n53 B.t5 500.531
R1740 B.n268 B.n199 449.257
R1741 B.n784 B.n783 449.257
R1742 B.n472 B.n471 449.257
R1743 B.n580 B.n91 449.257
R1744 B.n160 B.t0 370.135
R1745 B.n166 B.t6 370.135
R1746 B.n52 B.t3 370.135
R1747 B.n58 B.t9 370.135
R1748 B.n268 B.n267 163.367
R1749 B.n267 B.n266 163.367
R1750 B.n266 B.n201 163.367
R1751 B.n262 B.n201 163.367
R1752 B.n262 B.n261 163.367
R1753 B.n261 B.n260 163.367
R1754 B.n260 B.n203 163.367
R1755 B.n256 B.n203 163.367
R1756 B.n256 B.n255 163.367
R1757 B.n255 B.n254 163.367
R1758 B.n254 B.n205 163.367
R1759 B.n250 B.n205 163.367
R1760 B.n250 B.n249 163.367
R1761 B.n249 B.n248 163.367
R1762 B.n248 B.n207 163.367
R1763 B.n244 B.n207 163.367
R1764 B.n244 B.n243 163.367
R1765 B.n243 B.n242 163.367
R1766 B.n242 B.n209 163.367
R1767 B.n238 B.n209 163.367
R1768 B.n238 B.n237 163.367
R1769 B.n237 B.n236 163.367
R1770 B.n236 B.n211 163.367
R1771 B.n232 B.n211 163.367
R1772 B.n232 B.n231 163.367
R1773 B.n231 B.n230 163.367
R1774 B.n230 B.n213 163.367
R1775 B.n226 B.n213 163.367
R1776 B.n226 B.n225 163.367
R1777 B.n225 B.n224 163.367
R1778 B.n224 B.n215 163.367
R1779 B.n220 B.n215 163.367
R1780 B.n220 B.n219 163.367
R1781 B.n219 B.n218 163.367
R1782 B.n218 B.n2 163.367
R1783 B.n838 B.n2 163.367
R1784 B.n838 B.n837 163.367
R1785 B.n837 B.n836 163.367
R1786 B.n836 B.n3 163.367
R1787 B.n832 B.n3 163.367
R1788 B.n832 B.n831 163.367
R1789 B.n831 B.n830 163.367
R1790 B.n830 B.n5 163.367
R1791 B.n826 B.n5 163.367
R1792 B.n826 B.n825 163.367
R1793 B.n825 B.n824 163.367
R1794 B.n824 B.n7 163.367
R1795 B.n820 B.n7 163.367
R1796 B.n820 B.n819 163.367
R1797 B.n819 B.n818 163.367
R1798 B.n818 B.n9 163.367
R1799 B.n814 B.n9 163.367
R1800 B.n814 B.n813 163.367
R1801 B.n813 B.n812 163.367
R1802 B.n812 B.n11 163.367
R1803 B.n808 B.n11 163.367
R1804 B.n808 B.n807 163.367
R1805 B.n807 B.n806 163.367
R1806 B.n806 B.n13 163.367
R1807 B.n802 B.n13 163.367
R1808 B.n802 B.n801 163.367
R1809 B.n801 B.n800 163.367
R1810 B.n800 B.n15 163.367
R1811 B.n796 B.n15 163.367
R1812 B.n796 B.n795 163.367
R1813 B.n795 B.n794 163.367
R1814 B.n794 B.n17 163.367
R1815 B.n790 B.n17 163.367
R1816 B.n790 B.n789 163.367
R1817 B.n789 B.n788 163.367
R1818 B.n788 B.n19 163.367
R1819 B.n784 B.n19 163.367
R1820 B.n272 B.n199 163.367
R1821 B.n273 B.n272 163.367
R1822 B.n274 B.n273 163.367
R1823 B.n274 B.n197 163.367
R1824 B.n278 B.n197 163.367
R1825 B.n279 B.n278 163.367
R1826 B.n280 B.n279 163.367
R1827 B.n280 B.n195 163.367
R1828 B.n284 B.n195 163.367
R1829 B.n285 B.n284 163.367
R1830 B.n286 B.n285 163.367
R1831 B.n286 B.n193 163.367
R1832 B.n290 B.n193 163.367
R1833 B.n291 B.n290 163.367
R1834 B.n292 B.n291 163.367
R1835 B.n292 B.n191 163.367
R1836 B.n296 B.n191 163.367
R1837 B.n297 B.n296 163.367
R1838 B.n298 B.n297 163.367
R1839 B.n298 B.n189 163.367
R1840 B.n302 B.n189 163.367
R1841 B.n303 B.n302 163.367
R1842 B.n304 B.n303 163.367
R1843 B.n304 B.n187 163.367
R1844 B.n308 B.n187 163.367
R1845 B.n309 B.n308 163.367
R1846 B.n310 B.n309 163.367
R1847 B.n310 B.n185 163.367
R1848 B.n314 B.n185 163.367
R1849 B.n315 B.n314 163.367
R1850 B.n316 B.n315 163.367
R1851 B.n316 B.n183 163.367
R1852 B.n320 B.n183 163.367
R1853 B.n321 B.n320 163.367
R1854 B.n322 B.n321 163.367
R1855 B.n322 B.n181 163.367
R1856 B.n326 B.n181 163.367
R1857 B.n327 B.n326 163.367
R1858 B.n328 B.n327 163.367
R1859 B.n328 B.n179 163.367
R1860 B.n332 B.n179 163.367
R1861 B.n333 B.n332 163.367
R1862 B.n334 B.n333 163.367
R1863 B.n334 B.n177 163.367
R1864 B.n338 B.n177 163.367
R1865 B.n339 B.n338 163.367
R1866 B.n340 B.n339 163.367
R1867 B.n340 B.n175 163.367
R1868 B.n344 B.n175 163.367
R1869 B.n345 B.n344 163.367
R1870 B.n346 B.n345 163.367
R1871 B.n346 B.n173 163.367
R1872 B.n350 B.n173 163.367
R1873 B.n351 B.n350 163.367
R1874 B.n352 B.n351 163.367
R1875 B.n352 B.n171 163.367
R1876 B.n356 B.n171 163.367
R1877 B.n357 B.n356 163.367
R1878 B.n358 B.n357 163.367
R1879 B.n358 B.n169 163.367
R1880 B.n362 B.n169 163.367
R1881 B.n363 B.n362 163.367
R1882 B.n363 B.n165 163.367
R1883 B.n367 B.n165 163.367
R1884 B.n368 B.n367 163.367
R1885 B.n369 B.n368 163.367
R1886 B.n369 B.n163 163.367
R1887 B.n373 B.n163 163.367
R1888 B.n374 B.n373 163.367
R1889 B.n375 B.n374 163.367
R1890 B.n375 B.n159 163.367
R1891 B.n380 B.n159 163.367
R1892 B.n381 B.n380 163.367
R1893 B.n382 B.n381 163.367
R1894 B.n382 B.n157 163.367
R1895 B.n386 B.n157 163.367
R1896 B.n387 B.n386 163.367
R1897 B.n388 B.n387 163.367
R1898 B.n388 B.n155 163.367
R1899 B.n392 B.n155 163.367
R1900 B.n393 B.n392 163.367
R1901 B.n394 B.n393 163.367
R1902 B.n394 B.n153 163.367
R1903 B.n398 B.n153 163.367
R1904 B.n399 B.n398 163.367
R1905 B.n400 B.n399 163.367
R1906 B.n400 B.n151 163.367
R1907 B.n404 B.n151 163.367
R1908 B.n405 B.n404 163.367
R1909 B.n406 B.n405 163.367
R1910 B.n406 B.n149 163.367
R1911 B.n410 B.n149 163.367
R1912 B.n411 B.n410 163.367
R1913 B.n412 B.n411 163.367
R1914 B.n412 B.n147 163.367
R1915 B.n416 B.n147 163.367
R1916 B.n417 B.n416 163.367
R1917 B.n418 B.n417 163.367
R1918 B.n418 B.n145 163.367
R1919 B.n422 B.n145 163.367
R1920 B.n423 B.n422 163.367
R1921 B.n424 B.n423 163.367
R1922 B.n424 B.n143 163.367
R1923 B.n428 B.n143 163.367
R1924 B.n429 B.n428 163.367
R1925 B.n430 B.n429 163.367
R1926 B.n430 B.n141 163.367
R1927 B.n434 B.n141 163.367
R1928 B.n435 B.n434 163.367
R1929 B.n436 B.n435 163.367
R1930 B.n436 B.n139 163.367
R1931 B.n440 B.n139 163.367
R1932 B.n441 B.n440 163.367
R1933 B.n442 B.n441 163.367
R1934 B.n442 B.n137 163.367
R1935 B.n446 B.n137 163.367
R1936 B.n447 B.n446 163.367
R1937 B.n448 B.n447 163.367
R1938 B.n448 B.n135 163.367
R1939 B.n452 B.n135 163.367
R1940 B.n453 B.n452 163.367
R1941 B.n454 B.n453 163.367
R1942 B.n454 B.n133 163.367
R1943 B.n458 B.n133 163.367
R1944 B.n459 B.n458 163.367
R1945 B.n460 B.n459 163.367
R1946 B.n460 B.n131 163.367
R1947 B.n464 B.n131 163.367
R1948 B.n465 B.n464 163.367
R1949 B.n466 B.n465 163.367
R1950 B.n466 B.n129 163.367
R1951 B.n470 B.n129 163.367
R1952 B.n471 B.n470 163.367
R1953 B.n472 B.n127 163.367
R1954 B.n476 B.n127 163.367
R1955 B.n477 B.n476 163.367
R1956 B.n478 B.n477 163.367
R1957 B.n478 B.n125 163.367
R1958 B.n482 B.n125 163.367
R1959 B.n483 B.n482 163.367
R1960 B.n484 B.n483 163.367
R1961 B.n484 B.n123 163.367
R1962 B.n488 B.n123 163.367
R1963 B.n489 B.n488 163.367
R1964 B.n490 B.n489 163.367
R1965 B.n490 B.n121 163.367
R1966 B.n494 B.n121 163.367
R1967 B.n495 B.n494 163.367
R1968 B.n496 B.n495 163.367
R1969 B.n496 B.n119 163.367
R1970 B.n500 B.n119 163.367
R1971 B.n501 B.n500 163.367
R1972 B.n502 B.n501 163.367
R1973 B.n502 B.n117 163.367
R1974 B.n506 B.n117 163.367
R1975 B.n507 B.n506 163.367
R1976 B.n508 B.n507 163.367
R1977 B.n508 B.n115 163.367
R1978 B.n512 B.n115 163.367
R1979 B.n513 B.n512 163.367
R1980 B.n514 B.n513 163.367
R1981 B.n514 B.n113 163.367
R1982 B.n518 B.n113 163.367
R1983 B.n519 B.n518 163.367
R1984 B.n520 B.n519 163.367
R1985 B.n520 B.n111 163.367
R1986 B.n524 B.n111 163.367
R1987 B.n525 B.n524 163.367
R1988 B.n526 B.n525 163.367
R1989 B.n526 B.n109 163.367
R1990 B.n530 B.n109 163.367
R1991 B.n531 B.n530 163.367
R1992 B.n532 B.n531 163.367
R1993 B.n532 B.n107 163.367
R1994 B.n536 B.n107 163.367
R1995 B.n537 B.n536 163.367
R1996 B.n538 B.n537 163.367
R1997 B.n538 B.n105 163.367
R1998 B.n542 B.n105 163.367
R1999 B.n543 B.n542 163.367
R2000 B.n544 B.n543 163.367
R2001 B.n544 B.n103 163.367
R2002 B.n548 B.n103 163.367
R2003 B.n549 B.n548 163.367
R2004 B.n550 B.n549 163.367
R2005 B.n550 B.n101 163.367
R2006 B.n554 B.n101 163.367
R2007 B.n555 B.n554 163.367
R2008 B.n556 B.n555 163.367
R2009 B.n556 B.n99 163.367
R2010 B.n560 B.n99 163.367
R2011 B.n561 B.n560 163.367
R2012 B.n562 B.n561 163.367
R2013 B.n562 B.n97 163.367
R2014 B.n566 B.n97 163.367
R2015 B.n567 B.n566 163.367
R2016 B.n568 B.n567 163.367
R2017 B.n568 B.n95 163.367
R2018 B.n572 B.n95 163.367
R2019 B.n573 B.n572 163.367
R2020 B.n574 B.n573 163.367
R2021 B.n574 B.n93 163.367
R2022 B.n578 B.n93 163.367
R2023 B.n579 B.n578 163.367
R2024 B.n580 B.n579 163.367
R2025 B.n783 B.n782 163.367
R2026 B.n782 B.n21 163.367
R2027 B.n778 B.n21 163.367
R2028 B.n778 B.n777 163.367
R2029 B.n777 B.n776 163.367
R2030 B.n776 B.n23 163.367
R2031 B.n772 B.n23 163.367
R2032 B.n772 B.n771 163.367
R2033 B.n771 B.n770 163.367
R2034 B.n770 B.n25 163.367
R2035 B.n766 B.n25 163.367
R2036 B.n766 B.n765 163.367
R2037 B.n765 B.n764 163.367
R2038 B.n764 B.n27 163.367
R2039 B.n760 B.n27 163.367
R2040 B.n760 B.n759 163.367
R2041 B.n759 B.n758 163.367
R2042 B.n758 B.n29 163.367
R2043 B.n754 B.n29 163.367
R2044 B.n754 B.n753 163.367
R2045 B.n753 B.n752 163.367
R2046 B.n752 B.n31 163.367
R2047 B.n748 B.n31 163.367
R2048 B.n748 B.n747 163.367
R2049 B.n747 B.n746 163.367
R2050 B.n746 B.n33 163.367
R2051 B.n742 B.n33 163.367
R2052 B.n742 B.n741 163.367
R2053 B.n741 B.n740 163.367
R2054 B.n740 B.n35 163.367
R2055 B.n736 B.n35 163.367
R2056 B.n736 B.n735 163.367
R2057 B.n735 B.n734 163.367
R2058 B.n734 B.n37 163.367
R2059 B.n730 B.n37 163.367
R2060 B.n730 B.n729 163.367
R2061 B.n729 B.n728 163.367
R2062 B.n728 B.n39 163.367
R2063 B.n724 B.n39 163.367
R2064 B.n724 B.n723 163.367
R2065 B.n723 B.n722 163.367
R2066 B.n722 B.n41 163.367
R2067 B.n718 B.n41 163.367
R2068 B.n718 B.n717 163.367
R2069 B.n717 B.n716 163.367
R2070 B.n716 B.n43 163.367
R2071 B.n712 B.n43 163.367
R2072 B.n712 B.n711 163.367
R2073 B.n711 B.n710 163.367
R2074 B.n710 B.n45 163.367
R2075 B.n706 B.n45 163.367
R2076 B.n706 B.n705 163.367
R2077 B.n705 B.n704 163.367
R2078 B.n704 B.n47 163.367
R2079 B.n700 B.n47 163.367
R2080 B.n700 B.n699 163.367
R2081 B.n699 B.n698 163.367
R2082 B.n698 B.n49 163.367
R2083 B.n694 B.n49 163.367
R2084 B.n694 B.n693 163.367
R2085 B.n693 B.n692 163.367
R2086 B.n692 B.n51 163.367
R2087 B.n687 B.n51 163.367
R2088 B.n687 B.n686 163.367
R2089 B.n686 B.n685 163.367
R2090 B.n685 B.n55 163.367
R2091 B.n681 B.n55 163.367
R2092 B.n681 B.n680 163.367
R2093 B.n680 B.n679 163.367
R2094 B.n679 B.n57 163.367
R2095 B.n675 B.n57 163.367
R2096 B.n675 B.n674 163.367
R2097 B.n674 B.n61 163.367
R2098 B.n670 B.n61 163.367
R2099 B.n670 B.n669 163.367
R2100 B.n669 B.n668 163.367
R2101 B.n668 B.n63 163.367
R2102 B.n664 B.n63 163.367
R2103 B.n664 B.n663 163.367
R2104 B.n663 B.n662 163.367
R2105 B.n662 B.n65 163.367
R2106 B.n658 B.n65 163.367
R2107 B.n658 B.n657 163.367
R2108 B.n657 B.n656 163.367
R2109 B.n656 B.n67 163.367
R2110 B.n652 B.n67 163.367
R2111 B.n652 B.n651 163.367
R2112 B.n651 B.n650 163.367
R2113 B.n650 B.n69 163.367
R2114 B.n646 B.n69 163.367
R2115 B.n646 B.n645 163.367
R2116 B.n645 B.n644 163.367
R2117 B.n644 B.n71 163.367
R2118 B.n640 B.n71 163.367
R2119 B.n640 B.n639 163.367
R2120 B.n639 B.n638 163.367
R2121 B.n638 B.n73 163.367
R2122 B.n634 B.n73 163.367
R2123 B.n634 B.n633 163.367
R2124 B.n633 B.n632 163.367
R2125 B.n632 B.n75 163.367
R2126 B.n628 B.n75 163.367
R2127 B.n628 B.n627 163.367
R2128 B.n627 B.n626 163.367
R2129 B.n626 B.n77 163.367
R2130 B.n622 B.n77 163.367
R2131 B.n622 B.n621 163.367
R2132 B.n621 B.n620 163.367
R2133 B.n620 B.n79 163.367
R2134 B.n616 B.n79 163.367
R2135 B.n616 B.n615 163.367
R2136 B.n615 B.n614 163.367
R2137 B.n614 B.n81 163.367
R2138 B.n610 B.n81 163.367
R2139 B.n610 B.n609 163.367
R2140 B.n609 B.n608 163.367
R2141 B.n608 B.n83 163.367
R2142 B.n604 B.n83 163.367
R2143 B.n604 B.n603 163.367
R2144 B.n603 B.n602 163.367
R2145 B.n602 B.n85 163.367
R2146 B.n598 B.n85 163.367
R2147 B.n598 B.n597 163.367
R2148 B.n597 B.n596 163.367
R2149 B.n596 B.n87 163.367
R2150 B.n592 B.n87 163.367
R2151 B.n592 B.n591 163.367
R2152 B.n591 B.n590 163.367
R2153 B.n590 B.n89 163.367
R2154 B.n586 B.n89 163.367
R2155 B.n586 B.n585 163.367
R2156 B.n585 B.n584 163.367
R2157 B.n584 B.n91 163.367
R2158 B.n161 B.n160 61.0914
R2159 B.n167 B.n166 61.0914
R2160 B.n53 B.n52 61.0914
R2161 B.n59 B.n58 61.0914
R2162 B.n378 B.n161 59.5399
R2163 B.n168 B.n167 59.5399
R2164 B.n690 B.n53 59.5399
R2165 B.n60 B.n59 59.5399
R2166 B.n582 B.n581 29.1907
R2167 B.n785 B.n20 29.1907
R2168 B.n473 B.n128 29.1907
R2169 B.n270 B.n269 29.1907
R2170 B B.n839 18.0485
R2171 B.n781 B.n20 10.6151
R2172 B.n781 B.n780 10.6151
R2173 B.n780 B.n779 10.6151
R2174 B.n779 B.n22 10.6151
R2175 B.n775 B.n22 10.6151
R2176 B.n775 B.n774 10.6151
R2177 B.n774 B.n773 10.6151
R2178 B.n773 B.n24 10.6151
R2179 B.n769 B.n24 10.6151
R2180 B.n769 B.n768 10.6151
R2181 B.n768 B.n767 10.6151
R2182 B.n767 B.n26 10.6151
R2183 B.n763 B.n26 10.6151
R2184 B.n763 B.n762 10.6151
R2185 B.n762 B.n761 10.6151
R2186 B.n761 B.n28 10.6151
R2187 B.n757 B.n28 10.6151
R2188 B.n757 B.n756 10.6151
R2189 B.n756 B.n755 10.6151
R2190 B.n755 B.n30 10.6151
R2191 B.n751 B.n30 10.6151
R2192 B.n751 B.n750 10.6151
R2193 B.n750 B.n749 10.6151
R2194 B.n749 B.n32 10.6151
R2195 B.n745 B.n32 10.6151
R2196 B.n745 B.n744 10.6151
R2197 B.n744 B.n743 10.6151
R2198 B.n743 B.n34 10.6151
R2199 B.n739 B.n34 10.6151
R2200 B.n739 B.n738 10.6151
R2201 B.n738 B.n737 10.6151
R2202 B.n737 B.n36 10.6151
R2203 B.n733 B.n36 10.6151
R2204 B.n733 B.n732 10.6151
R2205 B.n732 B.n731 10.6151
R2206 B.n731 B.n38 10.6151
R2207 B.n727 B.n38 10.6151
R2208 B.n727 B.n726 10.6151
R2209 B.n726 B.n725 10.6151
R2210 B.n725 B.n40 10.6151
R2211 B.n721 B.n40 10.6151
R2212 B.n721 B.n720 10.6151
R2213 B.n720 B.n719 10.6151
R2214 B.n719 B.n42 10.6151
R2215 B.n715 B.n42 10.6151
R2216 B.n715 B.n714 10.6151
R2217 B.n714 B.n713 10.6151
R2218 B.n713 B.n44 10.6151
R2219 B.n709 B.n44 10.6151
R2220 B.n709 B.n708 10.6151
R2221 B.n708 B.n707 10.6151
R2222 B.n707 B.n46 10.6151
R2223 B.n703 B.n46 10.6151
R2224 B.n703 B.n702 10.6151
R2225 B.n702 B.n701 10.6151
R2226 B.n701 B.n48 10.6151
R2227 B.n697 B.n48 10.6151
R2228 B.n697 B.n696 10.6151
R2229 B.n696 B.n695 10.6151
R2230 B.n695 B.n50 10.6151
R2231 B.n691 B.n50 10.6151
R2232 B.n689 B.n688 10.6151
R2233 B.n688 B.n54 10.6151
R2234 B.n684 B.n54 10.6151
R2235 B.n684 B.n683 10.6151
R2236 B.n683 B.n682 10.6151
R2237 B.n682 B.n56 10.6151
R2238 B.n678 B.n56 10.6151
R2239 B.n678 B.n677 10.6151
R2240 B.n677 B.n676 10.6151
R2241 B.n673 B.n672 10.6151
R2242 B.n672 B.n671 10.6151
R2243 B.n671 B.n62 10.6151
R2244 B.n667 B.n62 10.6151
R2245 B.n667 B.n666 10.6151
R2246 B.n666 B.n665 10.6151
R2247 B.n665 B.n64 10.6151
R2248 B.n661 B.n64 10.6151
R2249 B.n661 B.n660 10.6151
R2250 B.n660 B.n659 10.6151
R2251 B.n659 B.n66 10.6151
R2252 B.n655 B.n66 10.6151
R2253 B.n655 B.n654 10.6151
R2254 B.n654 B.n653 10.6151
R2255 B.n653 B.n68 10.6151
R2256 B.n649 B.n68 10.6151
R2257 B.n649 B.n648 10.6151
R2258 B.n648 B.n647 10.6151
R2259 B.n647 B.n70 10.6151
R2260 B.n643 B.n70 10.6151
R2261 B.n643 B.n642 10.6151
R2262 B.n642 B.n641 10.6151
R2263 B.n641 B.n72 10.6151
R2264 B.n637 B.n72 10.6151
R2265 B.n637 B.n636 10.6151
R2266 B.n636 B.n635 10.6151
R2267 B.n635 B.n74 10.6151
R2268 B.n631 B.n74 10.6151
R2269 B.n631 B.n630 10.6151
R2270 B.n630 B.n629 10.6151
R2271 B.n629 B.n76 10.6151
R2272 B.n625 B.n76 10.6151
R2273 B.n625 B.n624 10.6151
R2274 B.n624 B.n623 10.6151
R2275 B.n623 B.n78 10.6151
R2276 B.n619 B.n78 10.6151
R2277 B.n619 B.n618 10.6151
R2278 B.n618 B.n617 10.6151
R2279 B.n617 B.n80 10.6151
R2280 B.n613 B.n80 10.6151
R2281 B.n613 B.n612 10.6151
R2282 B.n612 B.n611 10.6151
R2283 B.n611 B.n82 10.6151
R2284 B.n607 B.n82 10.6151
R2285 B.n607 B.n606 10.6151
R2286 B.n606 B.n605 10.6151
R2287 B.n605 B.n84 10.6151
R2288 B.n601 B.n84 10.6151
R2289 B.n601 B.n600 10.6151
R2290 B.n600 B.n599 10.6151
R2291 B.n599 B.n86 10.6151
R2292 B.n595 B.n86 10.6151
R2293 B.n595 B.n594 10.6151
R2294 B.n594 B.n593 10.6151
R2295 B.n593 B.n88 10.6151
R2296 B.n589 B.n88 10.6151
R2297 B.n589 B.n588 10.6151
R2298 B.n588 B.n587 10.6151
R2299 B.n587 B.n90 10.6151
R2300 B.n583 B.n90 10.6151
R2301 B.n583 B.n582 10.6151
R2302 B.n474 B.n473 10.6151
R2303 B.n475 B.n474 10.6151
R2304 B.n475 B.n126 10.6151
R2305 B.n479 B.n126 10.6151
R2306 B.n480 B.n479 10.6151
R2307 B.n481 B.n480 10.6151
R2308 B.n481 B.n124 10.6151
R2309 B.n485 B.n124 10.6151
R2310 B.n486 B.n485 10.6151
R2311 B.n487 B.n486 10.6151
R2312 B.n487 B.n122 10.6151
R2313 B.n491 B.n122 10.6151
R2314 B.n492 B.n491 10.6151
R2315 B.n493 B.n492 10.6151
R2316 B.n493 B.n120 10.6151
R2317 B.n497 B.n120 10.6151
R2318 B.n498 B.n497 10.6151
R2319 B.n499 B.n498 10.6151
R2320 B.n499 B.n118 10.6151
R2321 B.n503 B.n118 10.6151
R2322 B.n504 B.n503 10.6151
R2323 B.n505 B.n504 10.6151
R2324 B.n505 B.n116 10.6151
R2325 B.n509 B.n116 10.6151
R2326 B.n510 B.n509 10.6151
R2327 B.n511 B.n510 10.6151
R2328 B.n511 B.n114 10.6151
R2329 B.n515 B.n114 10.6151
R2330 B.n516 B.n515 10.6151
R2331 B.n517 B.n516 10.6151
R2332 B.n517 B.n112 10.6151
R2333 B.n521 B.n112 10.6151
R2334 B.n522 B.n521 10.6151
R2335 B.n523 B.n522 10.6151
R2336 B.n523 B.n110 10.6151
R2337 B.n527 B.n110 10.6151
R2338 B.n528 B.n527 10.6151
R2339 B.n529 B.n528 10.6151
R2340 B.n529 B.n108 10.6151
R2341 B.n533 B.n108 10.6151
R2342 B.n534 B.n533 10.6151
R2343 B.n535 B.n534 10.6151
R2344 B.n535 B.n106 10.6151
R2345 B.n539 B.n106 10.6151
R2346 B.n540 B.n539 10.6151
R2347 B.n541 B.n540 10.6151
R2348 B.n541 B.n104 10.6151
R2349 B.n545 B.n104 10.6151
R2350 B.n546 B.n545 10.6151
R2351 B.n547 B.n546 10.6151
R2352 B.n547 B.n102 10.6151
R2353 B.n551 B.n102 10.6151
R2354 B.n552 B.n551 10.6151
R2355 B.n553 B.n552 10.6151
R2356 B.n553 B.n100 10.6151
R2357 B.n557 B.n100 10.6151
R2358 B.n558 B.n557 10.6151
R2359 B.n559 B.n558 10.6151
R2360 B.n559 B.n98 10.6151
R2361 B.n563 B.n98 10.6151
R2362 B.n564 B.n563 10.6151
R2363 B.n565 B.n564 10.6151
R2364 B.n565 B.n96 10.6151
R2365 B.n569 B.n96 10.6151
R2366 B.n570 B.n569 10.6151
R2367 B.n571 B.n570 10.6151
R2368 B.n571 B.n94 10.6151
R2369 B.n575 B.n94 10.6151
R2370 B.n576 B.n575 10.6151
R2371 B.n577 B.n576 10.6151
R2372 B.n577 B.n92 10.6151
R2373 B.n581 B.n92 10.6151
R2374 B.n271 B.n270 10.6151
R2375 B.n271 B.n198 10.6151
R2376 B.n275 B.n198 10.6151
R2377 B.n276 B.n275 10.6151
R2378 B.n277 B.n276 10.6151
R2379 B.n277 B.n196 10.6151
R2380 B.n281 B.n196 10.6151
R2381 B.n282 B.n281 10.6151
R2382 B.n283 B.n282 10.6151
R2383 B.n283 B.n194 10.6151
R2384 B.n287 B.n194 10.6151
R2385 B.n288 B.n287 10.6151
R2386 B.n289 B.n288 10.6151
R2387 B.n289 B.n192 10.6151
R2388 B.n293 B.n192 10.6151
R2389 B.n294 B.n293 10.6151
R2390 B.n295 B.n294 10.6151
R2391 B.n295 B.n190 10.6151
R2392 B.n299 B.n190 10.6151
R2393 B.n300 B.n299 10.6151
R2394 B.n301 B.n300 10.6151
R2395 B.n301 B.n188 10.6151
R2396 B.n305 B.n188 10.6151
R2397 B.n306 B.n305 10.6151
R2398 B.n307 B.n306 10.6151
R2399 B.n307 B.n186 10.6151
R2400 B.n311 B.n186 10.6151
R2401 B.n312 B.n311 10.6151
R2402 B.n313 B.n312 10.6151
R2403 B.n313 B.n184 10.6151
R2404 B.n317 B.n184 10.6151
R2405 B.n318 B.n317 10.6151
R2406 B.n319 B.n318 10.6151
R2407 B.n319 B.n182 10.6151
R2408 B.n323 B.n182 10.6151
R2409 B.n324 B.n323 10.6151
R2410 B.n325 B.n324 10.6151
R2411 B.n325 B.n180 10.6151
R2412 B.n329 B.n180 10.6151
R2413 B.n330 B.n329 10.6151
R2414 B.n331 B.n330 10.6151
R2415 B.n331 B.n178 10.6151
R2416 B.n335 B.n178 10.6151
R2417 B.n336 B.n335 10.6151
R2418 B.n337 B.n336 10.6151
R2419 B.n337 B.n176 10.6151
R2420 B.n341 B.n176 10.6151
R2421 B.n342 B.n341 10.6151
R2422 B.n343 B.n342 10.6151
R2423 B.n343 B.n174 10.6151
R2424 B.n347 B.n174 10.6151
R2425 B.n348 B.n347 10.6151
R2426 B.n349 B.n348 10.6151
R2427 B.n349 B.n172 10.6151
R2428 B.n353 B.n172 10.6151
R2429 B.n354 B.n353 10.6151
R2430 B.n355 B.n354 10.6151
R2431 B.n355 B.n170 10.6151
R2432 B.n359 B.n170 10.6151
R2433 B.n360 B.n359 10.6151
R2434 B.n361 B.n360 10.6151
R2435 B.n365 B.n364 10.6151
R2436 B.n366 B.n365 10.6151
R2437 B.n366 B.n164 10.6151
R2438 B.n370 B.n164 10.6151
R2439 B.n371 B.n370 10.6151
R2440 B.n372 B.n371 10.6151
R2441 B.n372 B.n162 10.6151
R2442 B.n376 B.n162 10.6151
R2443 B.n377 B.n376 10.6151
R2444 B.n379 B.n158 10.6151
R2445 B.n383 B.n158 10.6151
R2446 B.n384 B.n383 10.6151
R2447 B.n385 B.n384 10.6151
R2448 B.n385 B.n156 10.6151
R2449 B.n389 B.n156 10.6151
R2450 B.n390 B.n389 10.6151
R2451 B.n391 B.n390 10.6151
R2452 B.n391 B.n154 10.6151
R2453 B.n395 B.n154 10.6151
R2454 B.n396 B.n395 10.6151
R2455 B.n397 B.n396 10.6151
R2456 B.n397 B.n152 10.6151
R2457 B.n401 B.n152 10.6151
R2458 B.n402 B.n401 10.6151
R2459 B.n403 B.n402 10.6151
R2460 B.n403 B.n150 10.6151
R2461 B.n407 B.n150 10.6151
R2462 B.n408 B.n407 10.6151
R2463 B.n409 B.n408 10.6151
R2464 B.n409 B.n148 10.6151
R2465 B.n413 B.n148 10.6151
R2466 B.n414 B.n413 10.6151
R2467 B.n415 B.n414 10.6151
R2468 B.n415 B.n146 10.6151
R2469 B.n419 B.n146 10.6151
R2470 B.n420 B.n419 10.6151
R2471 B.n421 B.n420 10.6151
R2472 B.n421 B.n144 10.6151
R2473 B.n425 B.n144 10.6151
R2474 B.n426 B.n425 10.6151
R2475 B.n427 B.n426 10.6151
R2476 B.n427 B.n142 10.6151
R2477 B.n431 B.n142 10.6151
R2478 B.n432 B.n431 10.6151
R2479 B.n433 B.n432 10.6151
R2480 B.n433 B.n140 10.6151
R2481 B.n437 B.n140 10.6151
R2482 B.n438 B.n437 10.6151
R2483 B.n439 B.n438 10.6151
R2484 B.n439 B.n138 10.6151
R2485 B.n443 B.n138 10.6151
R2486 B.n444 B.n443 10.6151
R2487 B.n445 B.n444 10.6151
R2488 B.n445 B.n136 10.6151
R2489 B.n449 B.n136 10.6151
R2490 B.n450 B.n449 10.6151
R2491 B.n451 B.n450 10.6151
R2492 B.n451 B.n134 10.6151
R2493 B.n455 B.n134 10.6151
R2494 B.n456 B.n455 10.6151
R2495 B.n457 B.n456 10.6151
R2496 B.n457 B.n132 10.6151
R2497 B.n461 B.n132 10.6151
R2498 B.n462 B.n461 10.6151
R2499 B.n463 B.n462 10.6151
R2500 B.n463 B.n130 10.6151
R2501 B.n467 B.n130 10.6151
R2502 B.n468 B.n467 10.6151
R2503 B.n469 B.n468 10.6151
R2504 B.n469 B.n128 10.6151
R2505 B.n269 B.n200 10.6151
R2506 B.n265 B.n200 10.6151
R2507 B.n265 B.n264 10.6151
R2508 B.n264 B.n263 10.6151
R2509 B.n263 B.n202 10.6151
R2510 B.n259 B.n202 10.6151
R2511 B.n259 B.n258 10.6151
R2512 B.n258 B.n257 10.6151
R2513 B.n257 B.n204 10.6151
R2514 B.n253 B.n204 10.6151
R2515 B.n253 B.n252 10.6151
R2516 B.n252 B.n251 10.6151
R2517 B.n251 B.n206 10.6151
R2518 B.n247 B.n206 10.6151
R2519 B.n247 B.n246 10.6151
R2520 B.n246 B.n245 10.6151
R2521 B.n245 B.n208 10.6151
R2522 B.n241 B.n208 10.6151
R2523 B.n241 B.n240 10.6151
R2524 B.n240 B.n239 10.6151
R2525 B.n239 B.n210 10.6151
R2526 B.n235 B.n210 10.6151
R2527 B.n235 B.n234 10.6151
R2528 B.n234 B.n233 10.6151
R2529 B.n233 B.n212 10.6151
R2530 B.n229 B.n212 10.6151
R2531 B.n229 B.n228 10.6151
R2532 B.n228 B.n227 10.6151
R2533 B.n227 B.n214 10.6151
R2534 B.n223 B.n214 10.6151
R2535 B.n223 B.n222 10.6151
R2536 B.n222 B.n221 10.6151
R2537 B.n221 B.n216 10.6151
R2538 B.n217 B.n216 10.6151
R2539 B.n217 B.n0 10.6151
R2540 B.n835 B.n1 10.6151
R2541 B.n835 B.n834 10.6151
R2542 B.n834 B.n833 10.6151
R2543 B.n833 B.n4 10.6151
R2544 B.n829 B.n4 10.6151
R2545 B.n829 B.n828 10.6151
R2546 B.n828 B.n827 10.6151
R2547 B.n827 B.n6 10.6151
R2548 B.n823 B.n6 10.6151
R2549 B.n823 B.n822 10.6151
R2550 B.n822 B.n821 10.6151
R2551 B.n821 B.n8 10.6151
R2552 B.n817 B.n8 10.6151
R2553 B.n817 B.n816 10.6151
R2554 B.n816 B.n815 10.6151
R2555 B.n815 B.n10 10.6151
R2556 B.n811 B.n10 10.6151
R2557 B.n811 B.n810 10.6151
R2558 B.n810 B.n809 10.6151
R2559 B.n809 B.n12 10.6151
R2560 B.n805 B.n12 10.6151
R2561 B.n805 B.n804 10.6151
R2562 B.n804 B.n803 10.6151
R2563 B.n803 B.n14 10.6151
R2564 B.n799 B.n14 10.6151
R2565 B.n799 B.n798 10.6151
R2566 B.n798 B.n797 10.6151
R2567 B.n797 B.n16 10.6151
R2568 B.n793 B.n16 10.6151
R2569 B.n793 B.n792 10.6151
R2570 B.n792 B.n791 10.6151
R2571 B.n791 B.n18 10.6151
R2572 B.n787 B.n18 10.6151
R2573 B.n787 B.n786 10.6151
R2574 B.n786 B.n785 10.6151
R2575 B.n691 B.n690 9.36635
R2576 B.n673 B.n60 9.36635
R2577 B.n361 B.n168 9.36635
R2578 B.n379 B.n378 9.36635
R2579 B.n839 B.n0 2.81026
R2580 B.n839 B.n1 2.81026
R2581 B.n690 B.n689 1.24928
R2582 B.n676 B.n60 1.24928
R2583 B.n364 B.n168 1.24928
R2584 B.n378 B.n377 1.24928
R2585 VN.n0 VN.t3 196.916
R2586 VN.n1 VN.t0 196.916
R2587 VN.n0 VN.t1 196.024
R2588 VN.n1 VN.t2 196.024
R2589 VN VN.n1 55.9831
R2590 VN VN.n0 3.47936
R2591 VDD2.n2 VDD2.n0 115.984
R2592 VDD2.n2 VDD2.n1 67.8029
R2593 VDD2.n1 VDD2.t1 1.71762
R2594 VDD2.n1 VDD2.t3 1.71762
R2595 VDD2.n0 VDD2.t0 1.71762
R2596 VDD2.n0 VDD2.t2 1.71762
R2597 VDD2 VDD2.n2 0.0586897
C0 w_n2860_n4754# VTAIL 5.52599f
C1 B w_n2860_n4754# 11.4595f
C2 w_n2860_n4754# VN 5.01412f
C3 VP w_n2860_n4754# 5.38234f
C4 B VTAIL 7.34586f
C5 VDD1 VDD2 1.07487f
C6 VN VTAIL 7.04791f
C7 VP VTAIL 7.06202f
C8 B VN 1.23184f
C9 B VP 1.84391f
C10 VP VN 7.63225f
C11 VDD1 w_n2860_n4754# 1.67835f
C12 VDD2 w_n2860_n4754# 1.73935f
C13 VDD1 VTAIL 7.0457f
C14 VDD1 B 1.48665f
C15 VDD2 VTAIL 7.10138f
C16 VDD1 VN 0.149037f
C17 VDD1 VP 7.67955f
C18 VDD2 B 1.54245f
C19 VDD2 VN 7.42124f
C20 VDD2 VP 0.408142f
C21 VDD2 VSUBS 1.150336f
C22 VDD1 VSUBS 6.72053f
C23 VTAIL VSUBS 1.566739f
C24 VN VSUBS 5.8137f
C25 VP VSUBS 2.646377f
C26 B VSUBS 5.05171f
C27 w_n2860_n4754# VSUBS 0.166143p
C28 VDD2.t0 VSUBS 0.395688f
C29 VDD2.t2 VSUBS 0.395688f
C30 VDD2.n0 VSUBS 4.31662f
C31 VDD2.t1 VSUBS 0.395688f
C32 VDD2.t3 VSUBS 0.395688f
C33 VDD2.n1 VSUBS 3.30296f
C34 VDD2.n2 VSUBS 5.06052f
C35 VN.t3 VSUBS 4.38346f
C36 VN.t1 VSUBS 4.37635f
C37 VN.n0 VSUBS 2.79037f
C38 VN.t0 VSUBS 4.38346f
C39 VN.t2 VSUBS 4.37635f
C40 VN.n1 VSUBS 4.61007f
C41 B.n0 VSUBS 0.003696f
C42 B.n1 VSUBS 0.003696f
C43 B.n2 VSUBS 0.005845f
C44 B.n3 VSUBS 0.005845f
C45 B.n4 VSUBS 0.005845f
C46 B.n5 VSUBS 0.005845f
C47 B.n6 VSUBS 0.005845f
C48 B.n7 VSUBS 0.005845f
C49 B.n8 VSUBS 0.005845f
C50 B.n9 VSUBS 0.005845f
C51 B.n10 VSUBS 0.005845f
C52 B.n11 VSUBS 0.005845f
C53 B.n12 VSUBS 0.005845f
C54 B.n13 VSUBS 0.005845f
C55 B.n14 VSUBS 0.005845f
C56 B.n15 VSUBS 0.005845f
C57 B.n16 VSUBS 0.005845f
C58 B.n17 VSUBS 0.005845f
C59 B.n18 VSUBS 0.005845f
C60 B.n19 VSUBS 0.005845f
C61 B.n20 VSUBS 0.013165f
C62 B.n21 VSUBS 0.005845f
C63 B.n22 VSUBS 0.005845f
C64 B.n23 VSUBS 0.005845f
C65 B.n24 VSUBS 0.005845f
C66 B.n25 VSUBS 0.005845f
C67 B.n26 VSUBS 0.005845f
C68 B.n27 VSUBS 0.005845f
C69 B.n28 VSUBS 0.005845f
C70 B.n29 VSUBS 0.005845f
C71 B.n30 VSUBS 0.005845f
C72 B.n31 VSUBS 0.005845f
C73 B.n32 VSUBS 0.005845f
C74 B.n33 VSUBS 0.005845f
C75 B.n34 VSUBS 0.005845f
C76 B.n35 VSUBS 0.005845f
C77 B.n36 VSUBS 0.005845f
C78 B.n37 VSUBS 0.005845f
C79 B.n38 VSUBS 0.005845f
C80 B.n39 VSUBS 0.005845f
C81 B.n40 VSUBS 0.005845f
C82 B.n41 VSUBS 0.005845f
C83 B.n42 VSUBS 0.005845f
C84 B.n43 VSUBS 0.005845f
C85 B.n44 VSUBS 0.005845f
C86 B.n45 VSUBS 0.005845f
C87 B.n46 VSUBS 0.005845f
C88 B.n47 VSUBS 0.005845f
C89 B.n48 VSUBS 0.005845f
C90 B.n49 VSUBS 0.005845f
C91 B.n50 VSUBS 0.005845f
C92 B.n51 VSUBS 0.005845f
C93 B.t5 VSUBS 0.312079f
C94 B.t4 VSUBS 0.342107f
C95 B.t3 VSUBS 1.98241f
C96 B.n52 VSUBS 0.528329f
C97 B.n53 VSUBS 0.284392f
C98 B.n54 VSUBS 0.005845f
C99 B.n55 VSUBS 0.005845f
C100 B.n56 VSUBS 0.005845f
C101 B.n57 VSUBS 0.005845f
C102 B.t11 VSUBS 0.312082f
C103 B.t10 VSUBS 0.34211f
C104 B.t9 VSUBS 1.98241f
C105 B.n58 VSUBS 0.528326f
C106 B.n59 VSUBS 0.284389f
C107 B.n60 VSUBS 0.013542f
C108 B.n61 VSUBS 0.005845f
C109 B.n62 VSUBS 0.005845f
C110 B.n63 VSUBS 0.005845f
C111 B.n64 VSUBS 0.005845f
C112 B.n65 VSUBS 0.005845f
C113 B.n66 VSUBS 0.005845f
C114 B.n67 VSUBS 0.005845f
C115 B.n68 VSUBS 0.005845f
C116 B.n69 VSUBS 0.005845f
C117 B.n70 VSUBS 0.005845f
C118 B.n71 VSUBS 0.005845f
C119 B.n72 VSUBS 0.005845f
C120 B.n73 VSUBS 0.005845f
C121 B.n74 VSUBS 0.005845f
C122 B.n75 VSUBS 0.005845f
C123 B.n76 VSUBS 0.005845f
C124 B.n77 VSUBS 0.005845f
C125 B.n78 VSUBS 0.005845f
C126 B.n79 VSUBS 0.005845f
C127 B.n80 VSUBS 0.005845f
C128 B.n81 VSUBS 0.005845f
C129 B.n82 VSUBS 0.005845f
C130 B.n83 VSUBS 0.005845f
C131 B.n84 VSUBS 0.005845f
C132 B.n85 VSUBS 0.005845f
C133 B.n86 VSUBS 0.005845f
C134 B.n87 VSUBS 0.005845f
C135 B.n88 VSUBS 0.005845f
C136 B.n89 VSUBS 0.005845f
C137 B.n90 VSUBS 0.005845f
C138 B.n91 VSUBS 0.013165f
C139 B.n92 VSUBS 0.005845f
C140 B.n93 VSUBS 0.005845f
C141 B.n94 VSUBS 0.005845f
C142 B.n95 VSUBS 0.005845f
C143 B.n96 VSUBS 0.005845f
C144 B.n97 VSUBS 0.005845f
C145 B.n98 VSUBS 0.005845f
C146 B.n99 VSUBS 0.005845f
C147 B.n100 VSUBS 0.005845f
C148 B.n101 VSUBS 0.005845f
C149 B.n102 VSUBS 0.005845f
C150 B.n103 VSUBS 0.005845f
C151 B.n104 VSUBS 0.005845f
C152 B.n105 VSUBS 0.005845f
C153 B.n106 VSUBS 0.005845f
C154 B.n107 VSUBS 0.005845f
C155 B.n108 VSUBS 0.005845f
C156 B.n109 VSUBS 0.005845f
C157 B.n110 VSUBS 0.005845f
C158 B.n111 VSUBS 0.005845f
C159 B.n112 VSUBS 0.005845f
C160 B.n113 VSUBS 0.005845f
C161 B.n114 VSUBS 0.005845f
C162 B.n115 VSUBS 0.005845f
C163 B.n116 VSUBS 0.005845f
C164 B.n117 VSUBS 0.005845f
C165 B.n118 VSUBS 0.005845f
C166 B.n119 VSUBS 0.005845f
C167 B.n120 VSUBS 0.005845f
C168 B.n121 VSUBS 0.005845f
C169 B.n122 VSUBS 0.005845f
C170 B.n123 VSUBS 0.005845f
C171 B.n124 VSUBS 0.005845f
C172 B.n125 VSUBS 0.005845f
C173 B.n126 VSUBS 0.005845f
C174 B.n127 VSUBS 0.005845f
C175 B.n128 VSUBS 0.013165f
C176 B.n129 VSUBS 0.005845f
C177 B.n130 VSUBS 0.005845f
C178 B.n131 VSUBS 0.005845f
C179 B.n132 VSUBS 0.005845f
C180 B.n133 VSUBS 0.005845f
C181 B.n134 VSUBS 0.005845f
C182 B.n135 VSUBS 0.005845f
C183 B.n136 VSUBS 0.005845f
C184 B.n137 VSUBS 0.005845f
C185 B.n138 VSUBS 0.005845f
C186 B.n139 VSUBS 0.005845f
C187 B.n140 VSUBS 0.005845f
C188 B.n141 VSUBS 0.005845f
C189 B.n142 VSUBS 0.005845f
C190 B.n143 VSUBS 0.005845f
C191 B.n144 VSUBS 0.005845f
C192 B.n145 VSUBS 0.005845f
C193 B.n146 VSUBS 0.005845f
C194 B.n147 VSUBS 0.005845f
C195 B.n148 VSUBS 0.005845f
C196 B.n149 VSUBS 0.005845f
C197 B.n150 VSUBS 0.005845f
C198 B.n151 VSUBS 0.005845f
C199 B.n152 VSUBS 0.005845f
C200 B.n153 VSUBS 0.005845f
C201 B.n154 VSUBS 0.005845f
C202 B.n155 VSUBS 0.005845f
C203 B.n156 VSUBS 0.005845f
C204 B.n157 VSUBS 0.005845f
C205 B.n158 VSUBS 0.005845f
C206 B.n159 VSUBS 0.005845f
C207 B.t1 VSUBS 0.312082f
C208 B.t2 VSUBS 0.34211f
C209 B.t0 VSUBS 1.98241f
C210 B.n160 VSUBS 0.528326f
C211 B.n161 VSUBS 0.284389f
C212 B.n162 VSUBS 0.005845f
C213 B.n163 VSUBS 0.005845f
C214 B.n164 VSUBS 0.005845f
C215 B.n165 VSUBS 0.005845f
C216 B.t7 VSUBS 0.312079f
C217 B.t8 VSUBS 0.342107f
C218 B.t6 VSUBS 1.98241f
C219 B.n166 VSUBS 0.528329f
C220 B.n167 VSUBS 0.284392f
C221 B.n168 VSUBS 0.013542f
C222 B.n169 VSUBS 0.005845f
C223 B.n170 VSUBS 0.005845f
C224 B.n171 VSUBS 0.005845f
C225 B.n172 VSUBS 0.005845f
C226 B.n173 VSUBS 0.005845f
C227 B.n174 VSUBS 0.005845f
C228 B.n175 VSUBS 0.005845f
C229 B.n176 VSUBS 0.005845f
C230 B.n177 VSUBS 0.005845f
C231 B.n178 VSUBS 0.005845f
C232 B.n179 VSUBS 0.005845f
C233 B.n180 VSUBS 0.005845f
C234 B.n181 VSUBS 0.005845f
C235 B.n182 VSUBS 0.005845f
C236 B.n183 VSUBS 0.005845f
C237 B.n184 VSUBS 0.005845f
C238 B.n185 VSUBS 0.005845f
C239 B.n186 VSUBS 0.005845f
C240 B.n187 VSUBS 0.005845f
C241 B.n188 VSUBS 0.005845f
C242 B.n189 VSUBS 0.005845f
C243 B.n190 VSUBS 0.005845f
C244 B.n191 VSUBS 0.005845f
C245 B.n192 VSUBS 0.005845f
C246 B.n193 VSUBS 0.005845f
C247 B.n194 VSUBS 0.005845f
C248 B.n195 VSUBS 0.005845f
C249 B.n196 VSUBS 0.005845f
C250 B.n197 VSUBS 0.005845f
C251 B.n198 VSUBS 0.005845f
C252 B.n199 VSUBS 0.013165f
C253 B.n200 VSUBS 0.005845f
C254 B.n201 VSUBS 0.005845f
C255 B.n202 VSUBS 0.005845f
C256 B.n203 VSUBS 0.005845f
C257 B.n204 VSUBS 0.005845f
C258 B.n205 VSUBS 0.005845f
C259 B.n206 VSUBS 0.005845f
C260 B.n207 VSUBS 0.005845f
C261 B.n208 VSUBS 0.005845f
C262 B.n209 VSUBS 0.005845f
C263 B.n210 VSUBS 0.005845f
C264 B.n211 VSUBS 0.005845f
C265 B.n212 VSUBS 0.005845f
C266 B.n213 VSUBS 0.005845f
C267 B.n214 VSUBS 0.005845f
C268 B.n215 VSUBS 0.005845f
C269 B.n216 VSUBS 0.005845f
C270 B.n217 VSUBS 0.005845f
C271 B.n218 VSUBS 0.005845f
C272 B.n219 VSUBS 0.005845f
C273 B.n220 VSUBS 0.005845f
C274 B.n221 VSUBS 0.005845f
C275 B.n222 VSUBS 0.005845f
C276 B.n223 VSUBS 0.005845f
C277 B.n224 VSUBS 0.005845f
C278 B.n225 VSUBS 0.005845f
C279 B.n226 VSUBS 0.005845f
C280 B.n227 VSUBS 0.005845f
C281 B.n228 VSUBS 0.005845f
C282 B.n229 VSUBS 0.005845f
C283 B.n230 VSUBS 0.005845f
C284 B.n231 VSUBS 0.005845f
C285 B.n232 VSUBS 0.005845f
C286 B.n233 VSUBS 0.005845f
C287 B.n234 VSUBS 0.005845f
C288 B.n235 VSUBS 0.005845f
C289 B.n236 VSUBS 0.005845f
C290 B.n237 VSUBS 0.005845f
C291 B.n238 VSUBS 0.005845f
C292 B.n239 VSUBS 0.005845f
C293 B.n240 VSUBS 0.005845f
C294 B.n241 VSUBS 0.005845f
C295 B.n242 VSUBS 0.005845f
C296 B.n243 VSUBS 0.005845f
C297 B.n244 VSUBS 0.005845f
C298 B.n245 VSUBS 0.005845f
C299 B.n246 VSUBS 0.005845f
C300 B.n247 VSUBS 0.005845f
C301 B.n248 VSUBS 0.005845f
C302 B.n249 VSUBS 0.005845f
C303 B.n250 VSUBS 0.005845f
C304 B.n251 VSUBS 0.005845f
C305 B.n252 VSUBS 0.005845f
C306 B.n253 VSUBS 0.005845f
C307 B.n254 VSUBS 0.005845f
C308 B.n255 VSUBS 0.005845f
C309 B.n256 VSUBS 0.005845f
C310 B.n257 VSUBS 0.005845f
C311 B.n258 VSUBS 0.005845f
C312 B.n259 VSUBS 0.005845f
C313 B.n260 VSUBS 0.005845f
C314 B.n261 VSUBS 0.005845f
C315 B.n262 VSUBS 0.005845f
C316 B.n263 VSUBS 0.005845f
C317 B.n264 VSUBS 0.005845f
C318 B.n265 VSUBS 0.005845f
C319 B.n266 VSUBS 0.005845f
C320 B.n267 VSUBS 0.005845f
C321 B.n268 VSUBS 0.012279f
C322 B.n269 VSUBS 0.012279f
C323 B.n270 VSUBS 0.013165f
C324 B.n271 VSUBS 0.005845f
C325 B.n272 VSUBS 0.005845f
C326 B.n273 VSUBS 0.005845f
C327 B.n274 VSUBS 0.005845f
C328 B.n275 VSUBS 0.005845f
C329 B.n276 VSUBS 0.005845f
C330 B.n277 VSUBS 0.005845f
C331 B.n278 VSUBS 0.005845f
C332 B.n279 VSUBS 0.005845f
C333 B.n280 VSUBS 0.005845f
C334 B.n281 VSUBS 0.005845f
C335 B.n282 VSUBS 0.005845f
C336 B.n283 VSUBS 0.005845f
C337 B.n284 VSUBS 0.005845f
C338 B.n285 VSUBS 0.005845f
C339 B.n286 VSUBS 0.005845f
C340 B.n287 VSUBS 0.005845f
C341 B.n288 VSUBS 0.005845f
C342 B.n289 VSUBS 0.005845f
C343 B.n290 VSUBS 0.005845f
C344 B.n291 VSUBS 0.005845f
C345 B.n292 VSUBS 0.005845f
C346 B.n293 VSUBS 0.005845f
C347 B.n294 VSUBS 0.005845f
C348 B.n295 VSUBS 0.005845f
C349 B.n296 VSUBS 0.005845f
C350 B.n297 VSUBS 0.005845f
C351 B.n298 VSUBS 0.005845f
C352 B.n299 VSUBS 0.005845f
C353 B.n300 VSUBS 0.005845f
C354 B.n301 VSUBS 0.005845f
C355 B.n302 VSUBS 0.005845f
C356 B.n303 VSUBS 0.005845f
C357 B.n304 VSUBS 0.005845f
C358 B.n305 VSUBS 0.005845f
C359 B.n306 VSUBS 0.005845f
C360 B.n307 VSUBS 0.005845f
C361 B.n308 VSUBS 0.005845f
C362 B.n309 VSUBS 0.005845f
C363 B.n310 VSUBS 0.005845f
C364 B.n311 VSUBS 0.005845f
C365 B.n312 VSUBS 0.005845f
C366 B.n313 VSUBS 0.005845f
C367 B.n314 VSUBS 0.005845f
C368 B.n315 VSUBS 0.005845f
C369 B.n316 VSUBS 0.005845f
C370 B.n317 VSUBS 0.005845f
C371 B.n318 VSUBS 0.005845f
C372 B.n319 VSUBS 0.005845f
C373 B.n320 VSUBS 0.005845f
C374 B.n321 VSUBS 0.005845f
C375 B.n322 VSUBS 0.005845f
C376 B.n323 VSUBS 0.005845f
C377 B.n324 VSUBS 0.005845f
C378 B.n325 VSUBS 0.005845f
C379 B.n326 VSUBS 0.005845f
C380 B.n327 VSUBS 0.005845f
C381 B.n328 VSUBS 0.005845f
C382 B.n329 VSUBS 0.005845f
C383 B.n330 VSUBS 0.005845f
C384 B.n331 VSUBS 0.005845f
C385 B.n332 VSUBS 0.005845f
C386 B.n333 VSUBS 0.005845f
C387 B.n334 VSUBS 0.005845f
C388 B.n335 VSUBS 0.005845f
C389 B.n336 VSUBS 0.005845f
C390 B.n337 VSUBS 0.005845f
C391 B.n338 VSUBS 0.005845f
C392 B.n339 VSUBS 0.005845f
C393 B.n340 VSUBS 0.005845f
C394 B.n341 VSUBS 0.005845f
C395 B.n342 VSUBS 0.005845f
C396 B.n343 VSUBS 0.005845f
C397 B.n344 VSUBS 0.005845f
C398 B.n345 VSUBS 0.005845f
C399 B.n346 VSUBS 0.005845f
C400 B.n347 VSUBS 0.005845f
C401 B.n348 VSUBS 0.005845f
C402 B.n349 VSUBS 0.005845f
C403 B.n350 VSUBS 0.005845f
C404 B.n351 VSUBS 0.005845f
C405 B.n352 VSUBS 0.005845f
C406 B.n353 VSUBS 0.005845f
C407 B.n354 VSUBS 0.005845f
C408 B.n355 VSUBS 0.005845f
C409 B.n356 VSUBS 0.005845f
C410 B.n357 VSUBS 0.005845f
C411 B.n358 VSUBS 0.005845f
C412 B.n359 VSUBS 0.005845f
C413 B.n360 VSUBS 0.005845f
C414 B.n361 VSUBS 0.005501f
C415 B.n362 VSUBS 0.005845f
C416 B.n363 VSUBS 0.005845f
C417 B.n364 VSUBS 0.003266f
C418 B.n365 VSUBS 0.005845f
C419 B.n366 VSUBS 0.005845f
C420 B.n367 VSUBS 0.005845f
C421 B.n368 VSUBS 0.005845f
C422 B.n369 VSUBS 0.005845f
C423 B.n370 VSUBS 0.005845f
C424 B.n371 VSUBS 0.005845f
C425 B.n372 VSUBS 0.005845f
C426 B.n373 VSUBS 0.005845f
C427 B.n374 VSUBS 0.005845f
C428 B.n375 VSUBS 0.005845f
C429 B.n376 VSUBS 0.005845f
C430 B.n377 VSUBS 0.003266f
C431 B.n378 VSUBS 0.013542f
C432 B.n379 VSUBS 0.005501f
C433 B.n380 VSUBS 0.005845f
C434 B.n381 VSUBS 0.005845f
C435 B.n382 VSUBS 0.005845f
C436 B.n383 VSUBS 0.005845f
C437 B.n384 VSUBS 0.005845f
C438 B.n385 VSUBS 0.005845f
C439 B.n386 VSUBS 0.005845f
C440 B.n387 VSUBS 0.005845f
C441 B.n388 VSUBS 0.005845f
C442 B.n389 VSUBS 0.005845f
C443 B.n390 VSUBS 0.005845f
C444 B.n391 VSUBS 0.005845f
C445 B.n392 VSUBS 0.005845f
C446 B.n393 VSUBS 0.005845f
C447 B.n394 VSUBS 0.005845f
C448 B.n395 VSUBS 0.005845f
C449 B.n396 VSUBS 0.005845f
C450 B.n397 VSUBS 0.005845f
C451 B.n398 VSUBS 0.005845f
C452 B.n399 VSUBS 0.005845f
C453 B.n400 VSUBS 0.005845f
C454 B.n401 VSUBS 0.005845f
C455 B.n402 VSUBS 0.005845f
C456 B.n403 VSUBS 0.005845f
C457 B.n404 VSUBS 0.005845f
C458 B.n405 VSUBS 0.005845f
C459 B.n406 VSUBS 0.005845f
C460 B.n407 VSUBS 0.005845f
C461 B.n408 VSUBS 0.005845f
C462 B.n409 VSUBS 0.005845f
C463 B.n410 VSUBS 0.005845f
C464 B.n411 VSUBS 0.005845f
C465 B.n412 VSUBS 0.005845f
C466 B.n413 VSUBS 0.005845f
C467 B.n414 VSUBS 0.005845f
C468 B.n415 VSUBS 0.005845f
C469 B.n416 VSUBS 0.005845f
C470 B.n417 VSUBS 0.005845f
C471 B.n418 VSUBS 0.005845f
C472 B.n419 VSUBS 0.005845f
C473 B.n420 VSUBS 0.005845f
C474 B.n421 VSUBS 0.005845f
C475 B.n422 VSUBS 0.005845f
C476 B.n423 VSUBS 0.005845f
C477 B.n424 VSUBS 0.005845f
C478 B.n425 VSUBS 0.005845f
C479 B.n426 VSUBS 0.005845f
C480 B.n427 VSUBS 0.005845f
C481 B.n428 VSUBS 0.005845f
C482 B.n429 VSUBS 0.005845f
C483 B.n430 VSUBS 0.005845f
C484 B.n431 VSUBS 0.005845f
C485 B.n432 VSUBS 0.005845f
C486 B.n433 VSUBS 0.005845f
C487 B.n434 VSUBS 0.005845f
C488 B.n435 VSUBS 0.005845f
C489 B.n436 VSUBS 0.005845f
C490 B.n437 VSUBS 0.005845f
C491 B.n438 VSUBS 0.005845f
C492 B.n439 VSUBS 0.005845f
C493 B.n440 VSUBS 0.005845f
C494 B.n441 VSUBS 0.005845f
C495 B.n442 VSUBS 0.005845f
C496 B.n443 VSUBS 0.005845f
C497 B.n444 VSUBS 0.005845f
C498 B.n445 VSUBS 0.005845f
C499 B.n446 VSUBS 0.005845f
C500 B.n447 VSUBS 0.005845f
C501 B.n448 VSUBS 0.005845f
C502 B.n449 VSUBS 0.005845f
C503 B.n450 VSUBS 0.005845f
C504 B.n451 VSUBS 0.005845f
C505 B.n452 VSUBS 0.005845f
C506 B.n453 VSUBS 0.005845f
C507 B.n454 VSUBS 0.005845f
C508 B.n455 VSUBS 0.005845f
C509 B.n456 VSUBS 0.005845f
C510 B.n457 VSUBS 0.005845f
C511 B.n458 VSUBS 0.005845f
C512 B.n459 VSUBS 0.005845f
C513 B.n460 VSUBS 0.005845f
C514 B.n461 VSUBS 0.005845f
C515 B.n462 VSUBS 0.005845f
C516 B.n463 VSUBS 0.005845f
C517 B.n464 VSUBS 0.005845f
C518 B.n465 VSUBS 0.005845f
C519 B.n466 VSUBS 0.005845f
C520 B.n467 VSUBS 0.005845f
C521 B.n468 VSUBS 0.005845f
C522 B.n469 VSUBS 0.005845f
C523 B.n470 VSUBS 0.005845f
C524 B.n471 VSUBS 0.013165f
C525 B.n472 VSUBS 0.012279f
C526 B.n473 VSUBS 0.012279f
C527 B.n474 VSUBS 0.005845f
C528 B.n475 VSUBS 0.005845f
C529 B.n476 VSUBS 0.005845f
C530 B.n477 VSUBS 0.005845f
C531 B.n478 VSUBS 0.005845f
C532 B.n479 VSUBS 0.005845f
C533 B.n480 VSUBS 0.005845f
C534 B.n481 VSUBS 0.005845f
C535 B.n482 VSUBS 0.005845f
C536 B.n483 VSUBS 0.005845f
C537 B.n484 VSUBS 0.005845f
C538 B.n485 VSUBS 0.005845f
C539 B.n486 VSUBS 0.005845f
C540 B.n487 VSUBS 0.005845f
C541 B.n488 VSUBS 0.005845f
C542 B.n489 VSUBS 0.005845f
C543 B.n490 VSUBS 0.005845f
C544 B.n491 VSUBS 0.005845f
C545 B.n492 VSUBS 0.005845f
C546 B.n493 VSUBS 0.005845f
C547 B.n494 VSUBS 0.005845f
C548 B.n495 VSUBS 0.005845f
C549 B.n496 VSUBS 0.005845f
C550 B.n497 VSUBS 0.005845f
C551 B.n498 VSUBS 0.005845f
C552 B.n499 VSUBS 0.005845f
C553 B.n500 VSUBS 0.005845f
C554 B.n501 VSUBS 0.005845f
C555 B.n502 VSUBS 0.005845f
C556 B.n503 VSUBS 0.005845f
C557 B.n504 VSUBS 0.005845f
C558 B.n505 VSUBS 0.005845f
C559 B.n506 VSUBS 0.005845f
C560 B.n507 VSUBS 0.005845f
C561 B.n508 VSUBS 0.005845f
C562 B.n509 VSUBS 0.005845f
C563 B.n510 VSUBS 0.005845f
C564 B.n511 VSUBS 0.005845f
C565 B.n512 VSUBS 0.005845f
C566 B.n513 VSUBS 0.005845f
C567 B.n514 VSUBS 0.005845f
C568 B.n515 VSUBS 0.005845f
C569 B.n516 VSUBS 0.005845f
C570 B.n517 VSUBS 0.005845f
C571 B.n518 VSUBS 0.005845f
C572 B.n519 VSUBS 0.005845f
C573 B.n520 VSUBS 0.005845f
C574 B.n521 VSUBS 0.005845f
C575 B.n522 VSUBS 0.005845f
C576 B.n523 VSUBS 0.005845f
C577 B.n524 VSUBS 0.005845f
C578 B.n525 VSUBS 0.005845f
C579 B.n526 VSUBS 0.005845f
C580 B.n527 VSUBS 0.005845f
C581 B.n528 VSUBS 0.005845f
C582 B.n529 VSUBS 0.005845f
C583 B.n530 VSUBS 0.005845f
C584 B.n531 VSUBS 0.005845f
C585 B.n532 VSUBS 0.005845f
C586 B.n533 VSUBS 0.005845f
C587 B.n534 VSUBS 0.005845f
C588 B.n535 VSUBS 0.005845f
C589 B.n536 VSUBS 0.005845f
C590 B.n537 VSUBS 0.005845f
C591 B.n538 VSUBS 0.005845f
C592 B.n539 VSUBS 0.005845f
C593 B.n540 VSUBS 0.005845f
C594 B.n541 VSUBS 0.005845f
C595 B.n542 VSUBS 0.005845f
C596 B.n543 VSUBS 0.005845f
C597 B.n544 VSUBS 0.005845f
C598 B.n545 VSUBS 0.005845f
C599 B.n546 VSUBS 0.005845f
C600 B.n547 VSUBS 0.005845f
C601 B.n548 VSUBS 0.005845f
C602 B.n549 VSUBS 0.005845f
C603 B.n550 VSUBS 0.005845f
C604 B.n551 VSUBS 0.005845f
C605 B.n552 VSUBS 0.005845f
C606 B.n553 VSUBS 0.005845f
C607 B.n554 VSUBS 0.005845f
C608 B.n555 VSUBS 0.005845f
C609 B.n556 VSUBS 0.005845f
C610 B.n557 VSUBS 0.005845f
C611 B.n558 VSUBS 0.005845f
C612 B.n559 VSUBS 0.005845f
C613 B.n560 VSUBS 0.005845f
C614 B.n561 VSUBS 0.005845f
C615 B.n562 VSUBS 0.005845f
C616 B.n563 VSUBS 0.005845f
C617 B.n564 VSUBS 0.005845f
C618 B.n565 VSUBS 0.005845f
C619 B.n566 VSUBS 0.005845f
C620 B.n567 VSUBS 0.005845f
C621 B.n568 VSUBS 0.005845f
C622 B.n569 VSUBS 0.005845f
C623 B.n570 VSUBS 0.005845f
C624 B.n571 VSUBS 0.005845f
C625 B.n572 VSUBS 0.005845f
C626 B.n573 VSUBS 0.005845f
C627 B.n574 VSUBS 0.005845f
C628 B.n575 VSUBS 0.005845f
C629 B.n576 VSUBS 0.005845f
C630 B.n577 VSUBS 0.005845f
C631 B.n578 VSUBS 0.005845f
C632 B.n579 VSUBS 0.005845f
C633 B.n580 VSUBS 0.012279f
C634 B.n581 VSUBS 0.013052f
C635 B.n582 VSUBS 0.012392f
C636 B.n583 VSUBS 0.005845f
C637 B.n584 VSUBS 0.005845f
C638 B.n585 VSUBS 0.005845f
C639 B.n586 VSUBS 0.005845f
C640 B.n587 VSUBS 0.005845f
C641 B.n588 VSUBS 0.005845f
C642 B.n589 VSUBS 0.005845f
C643 B.n590 VSUBS 0.005845f
C644 B.n591 VSUBS 0.005845f
C645 B.n592 VSUBS 0.005845f
C646 B.n593 VSUBS 0.005845f
C647 B.n594 VSUBS 0.005845f
C648 B.n595 VSUBS 0.005845f
C649 B.n596 VSUBS 0.005845f
C650 B.n597 VSUBS 0.005845f
C651 B.n598 VSUBS 0.005845f
C652 B.n599 VSUBS 0.005845f
C653 B.n600 VSUBS 0.005845f
C654 B.n601 VSUBS 0.005845f
C655 B.n602 VSUBS 0.005845f
C656 B.n603 VSUBS 0.005845f
C657 B.n604 VSUBS 0.005845f
C658 B.n605 VSUBS 0.005845f
C659 B.n606 VSUBS 0.005845f
C660 B.n607 VSUBS 0.005845f
C661 B.n608 VSUBS 0.005845f
C662 B.n609 VSUBS 0.005845f
C663 B.n610 VSUBS 0.005845f
C664 B.n611 VSUBS 0.005845f
C665 B.n612 VSUBS 0.005845f
C666 B.n613 VSUBS 0.005845f
C667 B.n614 VSUBS 0.005845f
C668 B.n615 VSUBS 0.005845f
C669 B.n616 VSUBS 0.005845f
C670 B.n617 VSUBS 0.005845f
C671 B.n618 VSUBS 0.005845f
C672 B.n619 VSUBS 0.005845f
C673 B.n620 VSUBS 0.005845f
C674 B.n621 VSUBS 0.005845f
C675 B.n622 VSUBS 0.005845f
C676 B.n623 VSUBS 0.005845f
C677 B.n624 VSUBS 0.005845f
C678 B.n625 VSUBS 0.005845f
C679 B.n626 VSUBS 0.005845f
C680 B.n627 VSUBS 0.005845f
C681 B.n628 VSUBS 0.005845f
C682 B.n629 VSUBS 0.005845f
C683 B.n630 VSUBS 0.005845f
C684 B.n631 VSUBS 0.005845f
C685 B.n632 VSUBS 0.005845f
C686 B.n633 VSUBS 0.005845f
C687 B.n634 VSUBS 0.005845f
C688 B.n635 VSUBS 0.005845f
C689 B.n636 VSUBS 0.005845f
C690 B.n637 VSUBS 0.005845f
C691 B.n638 VSUBS 0.005845f
C692 B.n639 VSUBS 0.005845f
C693 B.n640 VSUBS 0.005845f
C694 B.n641 VSUBS 0.005845f
C695 B.n642 VSUBS 0.005845f
C696 B.n643 VSUBS 0.005845f
C697 B.n644 VSUBS 0.005845f
C698 B.n645 VSUBS 0.005845f
C699 B.n646 VSUBS 0.005845f
C700 B.n647 VSUBS 0.005845f
C701 B.n648 VSUBS 0.005845f
C702 B.n649 VSUBS 0.005845f
C703 B.n650 VSUBS 0.005845f
C704 B.n651 VSUBS 0.005845f
C705 B.n652 VSUBS 0.005845f
C706 B.n653 VSUBS 0.005845f
C707 B.n654 VSUBS 0.005845f
C708 B.n655 VSUBS 0.005845f
C709 B.n656 VSUBS 0.005845f
C710 B.n657 VSUBS 0.005845f
C711 B.n658 VSUBS 0.005845f
C712 B.n659 VSUBS 0.005845f
C713 B.n660 VSUBS 0.005845f
C714 B.n661 VSUBS 0.005845f
C715 B.n662 VSUBS 0.005845f
C716 B.n663 VSUBS 0.005845f
C717 B.n664 VSUBS 0.005845f
C718 B.n665 VSUBS 0.005845f
C719 B.n666 VSUBS 0.005845f
C720 B.n667 VSUBS 0.005845f
C721 B.n668 VSUBS 0.005845f
C722 B.n669 VSUBS 0.005845f
C723 B.n670 VSUBS 0.005845f
C724 B.n671 VSUBS 0.005845f
C725 B.n672 VSUBS 0.005845f
C726 B.n673 VSUBS 0.005501f
C727 B.n674 VSUBS 0.005845f
C728 B.n675 VSUBS 0.005845f
C729 B.n676 VSUBS 0.003266f
C730 B.n677 VSUBS 0.005845f
C731 B.n678 VSUBS 0.005845f
C732 B.n679 VSUBS 0.005845f
C733 B.n680 VSUBS 0.005845f
C734 B.n681 VSUBS 0.005845f
C735 B.n682 VSUBS 0.005845f
C736 B.n683 VSUBS 0.005845f
C737 B.n684 VSUBS 0.005845f
C738 B.n685 VSUBS 0.005845f
C739 B.n686 VSUBS 0.005845f
C740 B.n687 VSUBS 0.005845f
C741 B.n688 VSUBS 0.005845f
C742 B.n689 VSUBS 0.003266f
C743 B.n690 VSUBS 0.013542f
C744 B.n691 VSUBS 0.005501f
C745 B.n692 VSUBS 0.005845f
C746 B.n693 VSUBS 0.005845f
C747 B.n694 VSUBS 0.005845f
C748 B.n695 VSUBS 0.005845f
C749 B.n696 VSUBS 0.005845f
C750 B.n697 VSUBS 0.005845f
C751 B.n698 VSUBS 0.005845f
C752 B.n699 VSUBS 0.005845f
C753 B.n700 VSUBS 0.005845f
C754 B.n701 VSUBS 0.005845f
C755 B.n702 VSUBS 0.005845f
C756 B.n703 VSUBS 0.005845f
C757 B.n704 VSUBS 0.005845f
C758 B.n705 VSUBS 0.005845f
C759 B.n706 VSUBS 0.005845f
C760 B.n707 VSUBS 0.005845f
C761 B.n708 VSUBS 0.005845f
C762 B.n709 VSUBS 0.005845f
C763 B.n710 VSUBS 0.005845f
C764 B.n711 VSUBS 0.005845f
C765 B.n712 VSUBS 0.005845f
C766 B.n713 VSUBS 0.005845f
C767 B.n714 VSUBS 0.005845f
C768 B.n715 VSUBS 0.005845f
C769 B.n716 VSUBS 0.005845f
C770 B.n717 VSUBS 0.005845f
C771 B.n718 VSUBS 0.005845f
C772 B.n719 VSUBS 0.005845f
C773 B.n720 VSUBS 0.005845f
C774 B.n721 VSUBS 0.005845f
C775 B.n722 VSUBS 0.005845f
C776 B.n723 VSUBS 0.005845f
C777 B.n724 VSUBS 0.005845f
C778 B.n725 VSUBS 0.005845f
C779 B.n726 VSUBS 0.005845f
C780 B.n727 VSUBS 0.005845f
C781 B.n728 VSUBS 0.005845f
C782 B.n729 VSUBS 0.005845f
C783 B.n730 VSUBS 0.005845f
C784 B.n731 VSUBS 0.005845f
C785 B.n732 VSUBS 0.005845f
C786 B.n733 VSUBS 0.005845f
C787 B.n734 VSUBS 0.005845f
C788 B.n735 VSUBS 0.005845f
C789 B.n736 VSUBS 0.005845f
C790 B.n737 VSUBS 0.005845f
C791 B.n738 VSUBS 0.005845f
C792 B.n739 VSUBS 0.005845f
C793 B.n740 VSUBS 0.005845f
C794 B.n741 VSUBS 0.005845f
C795 B.n742 VSUBS 0.005845f
C796 B.n743 VSUBS 0.005845f
C797 B.n744 VSUBS 0.005845f
C798 B.n745 VSUBS 0.005845f
C799 B.n746 VSUBS 0.005845f
C800 B.n747 VSUBS 0.005845f
C801 B.n748 VSUBS 0.005845f
C802 B.n749 VSUBS 0.005845f
C803 B.n750 VSUBS 0.005845f
C804 B.n751 VSUBS 0.005845f
C805 B.n752 VSUBS 0.005845f
C806 B.n753 VSUBS 0.005845f
C807 B.n754 VSUBS 0.005845f
C808 B.n755 VSUBS 0.005845f
C809 B.n756 VSUBS 0.005845f
C810 B.n757 VSUBS 0.005845f
C811 B.n758 VSUBS 0.005845f
C812 B.n759 VSUBS 0.005845f
C813 B.n760 VSUBS 0.005845f
C814 B.n761 VSUBS 0.005845f
C815 B.n762 VSUBS 0.005845f
C816 B.n763 VSUBS 0.005845f
C817 B.n764 VSUBS 0.005845f
C818 B.n765 VSUBS 0.005845f
C819 B.n766 VSUBS 0.005845f
C820 B.n767 VSUBS 0.005845f
C821 B.n768 VSUBS 0.005845f
C822 B.n769 VSUBS 0.005845f
C823 B.n770 VSUBS 0.005845f
C824 B.n771 VSUBS 0.005845f
C825 B.n772 VSUBS 0.005845f
C826 B.n773 VSUBS 0.005845f
C827 B.n774 VSUBS 0.005845f
C828 B.n775 VSUBS 0.005845f
C829 B.n776 VSUBS 0.005845f
C830 B.n777 VSUBS 0.005845f
C831 B.n778 VSUBS 0.005845f
C832 B.n779 VSUBS 0.005845f
C833 B.n780 VSUBS 0.005845f
C834 B.n781 VSUBS 0.005845f
C835 B.n782 VSUBS 0.005845f
C836 B.n783 VSUBS 0.013165f
C837 B.n784 VSUBS 0.012279f
C838 B.n785 VSUBS 0.012279f
C839 B.n786 VSUBS 0.005845f
C840 B.n787 VSUBS 0.005845f
C841 B.n788 VSUBS 0.005845f
C842 B.n789 VSUBS 0.005845f
C843 B.n790 VSUBS 0.005845f
C844 B.n791 VSUBS 0.005845f
C845 B.n792 VSUBS 0.005845f
C846 B.n793 VSUBS 0.005845f
C847 B.n794 VSUBS 0.005845f
C848 B.n795 VSUBS 0.005845f
C849 B.n796 VSUBS 0.005845f
C850 B.n797 VSUBS 0.005845f
C851 B.n798 VSUBS 0.005845f
C852 B.n799 VSUBS 0.005845f
C853 B.n800 VSUBS 0.005845f
C854 B.n801 VSUBS 0.005845f
C855 B.n802 VSUBS 0.005845f
C856 B.n803 VSUBS 0.005845f
C857 B.n804 VSUBS 0.005845f
C858 B.n805 VSUBS 0.005845f
C859 B.n806 VSUBS 0.005845f
C860 B.n807 VSUBS 0.005845f
C861 B.n808 VSUBS 0.005845f
C862 B.n809 VSUBS 0.005845f
C863 B.n810 VSUBS 0.005845f
C864 B.n811 VSUBS 0.005845f
C865 B.n812 VSUBS 0.005845f
C866 B.n813 VSUBS 0.005845f
C867 B.n814 VSUBS 0.005845f
C868 B.n815 VSUBS 0.005845f
C869 B.n816 VSUBS 0.005845f
C870 B.n817 VSUBS 0.005845f
C871 B.n818 VSUBS 0.005845f
C872 B.n819 VSUBS 0.005845f
C873 B.n820 VSUBS 0.005845f
C874 B.n821 VSUBS 0.005845f
C875 B.n822 VSUBS 0.005845f
C876 B.n823 VSUBS 0.005845f
C877 B.n824 VSUBS 0.005845f
C878 B.n825 VSUBS 0.005845f
C879 B.n826 VSUBS 0.005845f
C880 B.n827 VSUBS 0.005845f
C881 B.n828 VSUBS 0.005845f
C882 B.n829 VSUBS 0.005845f
C883 B.n830 VSUBS 0.005845f
C884 B.n831 VSUBS 0.005845f
C885 B.n832 VSUBS 0.005845f
C886 B.n833 VSUBS 0.005845f
C887 B.n834 VSUBS 0.005845f
C888 B.n835 VSUBS 0.005845f
C889 B.n836 VSUBS 0.005845f
C890 B.n837 VSUBS 0.005845f
C891 B.n838 VSUBS 0.005845f
C892 B.n839 VSUBS 0.013235f
C893 VTAIL.n0 VSUBS 0.024349f
C894 VTAIL.n1 VSUBS 0.022159f
C895 VTAIL.n2 VSUBS 0.011907f
C896 VTAIL.n3 VSUBS 0.028144f
C897 VTAIL.n4 VSUBS 0.012607f
C898 VTAIL.n5 VSUBS 0.022159f
C899 VTAIL.n6 VSUBS 0.011907f
C900 VTAIL.n7 VSUBS 0.028144f
C901 VTAIL.n8 VSUBS 0.012607f
C902 VTAIL.n9 VSUBS 0.022159f
C903 VTAIL.n10 VSUBS 0.011907f
C904 VTAIL.n11 VSUBS 0.028144f
C905 VTAIL.n12 VSUBS 0.012607f
C906 VTAIL.n13 VSUBS 0.022159f
C907 VTAIL.n14 VSUBS 0.011907f
C908 VTAIL.n15 VSUBS 0.028144f
C909 VTAIL.n16 VSUBS 0.012607f
C910 VTAIL.n17 VSUBS 0.022159f
C911 VTAIL.n18 VSUBS 0.011907f
C912 VTAIL.n19 VSUBS 0.028144f
C913 VTAIL.n20 VSUBS 0.012607f
C914 VTAIL.n21 VSUBS 0.022159f
C915 VTAIL.n22 VSUBS 0.011907f
C916 VTAIL.n23 VSUBS 0.028144f
C917 VTAIL.n24 VSUBS 0.012607f
C918 VTAIL.n25 VSUBS 0.022159f
C919 VTAIL.n26 VSUBS 0.011907f
C920 VTAIL.n27 VSUBS 0.028144f
C921 VTAIL.n28 VSUBS 0.012607f
C922 VTAIL.n29 VSUBS 0.022159f
C923 VTAIL.n30 VSUBS 0.011907f
C924 VTAIL.n31 VSUBS 0.028144f
C925 VTAIL.n32 VSUBS 0.012607f
C926 VTAIL.n33 VSUBS 0.181886f
C927 VTAIL.t1 VSUBS 0.060467f
C928 VTAIL.n34 VSUBS 0.021108f
C929 VTAIL.n35 VSUBS 0.017904f
C930 VTAIL.n36 VSUBS 0.011907f
C931 VTAIL.n37 VSUBS 1.81021f
C932 VTAIL.n38 VSUBS 0.022159f
C933 VTAIL.n39 VSUBS 0.011907f
C934 VTAIL.n40 VSUBS 0.012607f
C935 VTAIL.n41 VSUBS 0.028144f
C936 VTAIL.n42 VSUBS 0.028144f
C937 VTAIL.n43 VSUBS 0.012607f
C938 VTAIL.n44 VSUBS 0.011907f
C939 VTAIL.n45 VSUBS 0.022159f
C940 VTAIL.n46 VSUBS 0.022159f
C941 VTAIL.n47 VSUBS 0.011907f
C942 VTAIL.n48 VSUBS 0.012607f
C943 VTAIL.n49 VSUBS 0.028144f
C944 VTAIL.n50 VSUBS 0.028144f
C945 VTAIL.n51 VSUBS 0.012607f
C946 VTAIL.n52 VSUBS 0.011907f
C947 VTAIL.n53 VSUBS 0.022159f
C948 VTAIL.n54 VSUBS 0.022159f
C949 VTAIL.n55 VSUBS 0.011907f
C950 VTAIL.n56 VSUBS 0.012607f
C951 VTAIL.n57 VSUBS 0.028144f
C952 VTAIL.n58 VSUBS 0.028144f
C953 VTAIL.n59 VSUBS 0.012607f
C954 VTAIL.n60 VSUBS 0.011907f
C955 VTAIL.n61 VSUBS 0.022159f
C956 VTAIL.n62 VSUBS 0.022159f
C957 VTAIL.n63 VSUBS 0.011907f
C958 VTAIL.n64 VSUBS 0.012607f
C959 VTAIL.n65 VSUBS 0.028144f
C960 VTAIL.n66 VSUBS 0.028144f
C961 VTAIL.n67 VSUBS 0.012607f
C962 VTAIL.n68 VSUBS 0.011907f
C963 VTAIL.n69 VSUBS 0.022159f
C964 VTAIL.n70 VSUBS 0.022159f
C965 VTAIL.n71 VSUBS 0.011907f
C966 VTAIL.n72 VSUBS 0.012607f
C967 VTAIL.n73 VSUBS 0.028144f
C968 VTAIL.n74 VSUBS 0.028144f
C969 VTAIL.n75 VSUBS 0.028144f
C970 VTAIL.n76 VSUBS 0.012607f
C971 VTAIL.n77 VSUBS 0.011907f
C972 VTAIL.n78 VSUBS 0.022159f
C973 VTAIL.n79 VSUBS 0.022159f
C974 VTAIL.n80 VSUBS 0.011907f
C975 VTAIL.n81 VSUBS 0.012257f
C976 VTAIL.n82 VSUBS 0.012257f
C977 VTAIL.n83 VSUBS 0.028144f
C978 VTAIL.n84 VSUBS 0.028144f
C979 VTAIL.n85 VSUBS 0.012607f
C980 VTAIL.n86 VSUBS 0.011907f
C981 VTAIL.n87 VSUBS 0.022159f
C982 VTAIL.n88 VSUBS 0.022159f
C983 VTAIL.n89 VSUBS 0.011907f
C984 VTAIL.n90 VSUBS 0.012607f
C985 VTAIL.n91 VSUBS 0.028144f
C986 VTAIL.n92 VSUBS 0.028144f
C987 VTAIL.n93 VSUBS 0.012607f
C988 VTAIL.n94 VSUBS 0.011907f
C989 VTAIL.n95 VSUBS 0.022159f
C990 VTAIL.n96 VSUBS 0.022159f
C991 VTAIL.n97 VSUBS 0.011907f
C992 VTAIL.n98 VSUBS 0.012607f
C993 VTAIL.n99 VSUBS 0.028144f
C994 VTAIL.n100 VSUBS 0.068138f
C995 VTAIL.n101 VSUBS 0.012607f
C996 VTAIL.n102 VSUBS 0.011907f
C997 VTAIL.n103 VSUBS 0.050311f
C998 VTAIL.n104 VSUBS 0.034238f
C999 VTAIL.n105 VSUBS 0.153058f
C1000 VTAIL.n106 VSUBS 0.024349f
C1001 VTAIL.n107 VSUBS 0.022159f
C1002 VTAIL.n108 VSUBS 0.011907f
C1003 VTAIL.n109 VSUBS 0.028144f
C1004 VTAIL.n110 VSUBS 0.012607f
C1005 VTAIL.n111 VSUBS 0.022159f
C1006 VTAIL.n112 VSUBS 0.011907f
C1007 VTAIL.n113 VSUBS 0.028144f
C1008 VTAIL.n114 VSUBS 0.012607f
C1009 VTAIL.n115 VSUBS 0.022159f
C1010 VTAIL.n116 VSUBS 0.011907f
C1011 VTAIL.n117 VSUBS 0.028144f
C1012 VTAIL.n118 VSUBS 0.012607f
C1013 VTAIL.n119 VSUBS 0.022159f
C1014 VTAIL.n120 VSUBS 0.011907f
C1015 VTAIL.n121 VSUBS 0.028144f
C1016 VTAIL.n122 VSUBS 0.012607f
C1017 VTAIL.n123 VSUBS 0.022159f
C1018 VTAIL.n124 VSUBS 0.011907f
C1019 VTAIL.n125 VSUBS 0.028144f
C1020 VTAIL.n126 VSUBS 0.012607f
C1021 VTAIL.n127 VSUBS 0.022159f
C1022 VTAIL.n128 VSUBS 0.011907f
C1023 VTAIL.n129 VSUBS 0.028144f
C1024 VTAIL.n130 VSUBS 0.012607f
C1025 VTAIL.n131 VSUBS 0.022159f
C1026 VTAIL.n132 VSUBS 0.011907f
C1027 VTAIL.n133 VSUBS 0.028144f
C1028 VTAIL.n134 VSUBS 0.012607f
C1029 VTAIL.n135 VSUBS 0.022159f
C1030 VTAIL.n136 VSUBS 0.011907f
C1031 VTAIL.n137 VSUBS 0.028144f
C1032 VTAIL.n138 VSUBS 0.012607f
C1033 VTAIL.n139 VSUBS 0.181886f
C1034 VTAIL.t5 VSUBS 0.060467f
C1035 VTAIL.n140 VSUBS 0.021108f
C1036 VTAIL.n141 VSUBS 0.017904f
C1037 VTAIL.n142 VSUBS 0.011907f
C1038 VTAIL.n143 VSUBS 1.81021f
C1039 VTAIL.n144 VSUBS 0.022159f
C1040 VTAIL.n145 VSUBS 0.011907f
C1041 VTAIL.n146 VSUBS 0.012607f
C1042 VTAIL.n147 VSUBS 0.028144f
C1043 VTAIL.n148 VSUBS 0.028144f
C1044 VTAIL.n149 VSUBS 0.012607f
C1045 VTAIL.n150 VSUBS 0.011907f
C1046 VTAIL.n151 VSUBS 0.022159f
C1047 VTAIL.n152 VSUBS 0.022159f
C1048 VTAIL.n153 VSUBS 0.011907f
C1049 VTAIL.n154 VSUBS 0.012607f
C1050 VTAIL.n155 VSUBS 0.028144f
C1051 VTAIL.n156 VSUBS 0.028144f
C1052 VTAIL.n157 VSUBS 0.012607f
C1053 VTAIL.n158 VSUBS 0.011907f
C1054 VTAIL.n159 VSUBS 0.022159f
C1055 VTAIL.n160 VSUBS 0.022159f
C1056 VTAIL.n161 VSUBS 0.011907f
C1057 VTAIL.n162 VSUBS 0.012607f
C1058 VTAIL.n163 VSUBS 0.028144f
C1059 VTAIL.n164 VSUBS 0.028144f
C1060 VTAIL.n165 VSUBS 0.012607f
C1061 VTAIL.n166 VSUBS 0.011907f
C1062 VTAIL.n167 VSUBS 0.022159f
C1063 VTAIL.n168 VSUBS 0.022159f
C1064 VTAIL.n169 VSUBS 0.011907f
C1065 VTAIL.n170 VSUBS 0.012607f
C1066 VTAIL.n171 VSUBS 0.028144f
C1067 VTAIL.n172 VSUBS 0.028144f
C1068 VTAIL.n173 VSUBS 0.012607f
C1069 VTAIL.n174 VSUBS 0.011907f
C1070 VTAIL.n175 VSUBS 0.022159f
C1071 VTAIL.n176 VSUBS 0.022159f
C1072 VTAIL.n177 VSUBS 0.011907f
C1073 VTAIL.n178 VSUBS 0.012607f
C1074 VTAIL.n179 VSUBS 0.028144f
C1075 VTAIL.n180 VSUBS 0.028144f
C1076 VTAIL.n181 VSUBS 0.028144f
C1077 VTAIL.n182 VSUBS 0.012607f
C1078 VTAIL.n183 VSUBS 0.011907f
C1079 VTAIL.n184 VSUBS 0.022159f
C1080 VTAIL.n185 VSUBS 0.022159f
C1081 VTAIL.n186 VSUBS 0.011907f
C1082 VTAIL.n187 VSUBS 0.012257f
C1083 VTAIL.n188 VSUBS 0.012257f
C1084 VTAIL.n189 VSUBS 0.028144f
C1085 VTAIL.n190 VSUBS 0.028144f
C1086 VTAIL.n191 VSUBS 0.012607f
C1087 VTAIL.n192 VSUBS 0.011907f
C1088 VTAIL.n193 VSUBS 0.022159f
C1089 VTAIL.n194 VSUBS 0.022159f
C1090 VTAIL.n195 VSUBS 0.011907f
C1091 VTAIL.n196 VSUBS 0.012607f
C1092 VTAIL.n197 VSUBS 0.028144f
C1093 VTAIL.n198 VSUBS 0.028144f
C1094 VTAIL.n199 VSUBS 0.012607f
C1095 VTAIL.n200 VSUBS 0.011907f
C1096 VTAIL.n201 VSUBS 0.022159f
C1097 VTAIL.n202 VSUBS 0.022159f
C1098 VTAIL.n203 VSUBS 0.011907f
C1099 VTAIL.n204 VSUBS 0.012607f
C1100 VTAIL.n205 VSUBS 0.028144f
C1101 VTAIL.n206 VSUBS 0.068138f
C1102 VTAIL.n207 VSUBS 0.012607f
C1103 VTAIL.n208 VSUBS 0.011907f
C1104 VTAIL.n209 VSUBS 0.050311f
C1105 VTAIL.n210 VSUBS 0.034238f
C1106 VTAIL.n211 VSUBS 0.245847f
C1107 VTAIL.n212 VSUBS 0.024349f
C1108 VTAIL.n213 VSUBS 0.022159f
C1109 VTAIL.n214 VSUBS 0.011907f
C1110 VTAIL.n215 VSUBS 0.028144f
C1111 VTAIL.n216 VSUBS 0.012607f
C1112 VTAIL.n217 VSUBS 0.022159f
C1113 VTAIL.n218 VSUBS 0.011907f
C1114 VTAIL.n219 VSUBS 0.028144f
C1115 VTAIL.n220 VSUBS 0.012607f
C1116 VTAIL.n221 VSUBS 0.022159f
C1117 VTAIL.n222 VSUBS 0.011907f
C1118 VTAIL.n223 VSUBS 0.028144f
C1119 VTAIL.n224 VSUBS 0.012607f
C1120 VTAIL.n225 VSUBS 0.022159f
C1121 VTAIL.n226 VSUBS 0.011907f
C1122 VTAIL.n227 VSUBS 0.028144f
C1123 VTAIL.n228 VSUBS 0.012607f
C1124 VTAIL.n229 VSUBS 0.022159f
C1125 VTAIL.n230 VSUBS 0.011907f
C1126 VTAIL.n231 VSUBS 0.028144f
C1127 VTAIL.n232 VSUBS 0.012607f
C1128 VTAIL.n233 VSUBS 0.022159f
C1129 VTAIL.n234 VSUBS 0.011907f
C1130 VTAIL.n235 VSUBS 0.028144f
C1131 VTAIL.n236 VSUBS 0.012607f
C1132 VTAIL.n237 VSUBS 0.022159f
C1133 VTAIL.n238 VSUBS 0.011907f
C1134 VTAIL.n239 VSUBS 0.028144f
C1135 VTAIL.n240 VSUBS 0.012607f
C1136 VTAIL.n241 VSUBS 0.022159f
C1137 VTAIL.n242 VSUBS 0.011907f
C1138 VTAIL.n243 VSUBS 0.028144f
C1139 VTAIL.n244 VSUBS 0.012607f
C1140 VTAIL.n245 VSUBS 0.181886f
C1141 VTAIL.t7 VSUBS 0.060467f
C1142 VTAIL.n246 VSUBS 0.021108f
C1143 VTAIL.n247 VSUBS 0.017904f
C1144 VTAIL.n248 VSUBS 0.011907f
C1145 VTAIL.n249 VSUBS 1.81021f
C1146 VTAIL.n250 VSUBS 0.022159f
C1147 VTAIL.n251 VSUBS 0.011907f
C1148 VTAIL.n252 VSUBS 0.012607f
C1149 VTAIL.n253 VSUBS 0.028144f
C1150 VTAIL.n254 VSUBS 0.028144f
C1151 VTAIL.n255 VSUBS 0.012607f
C1152 VTAIL.n256 VSUBS 0.011907f
C1153 VTAIL.n257 VSUBS 0.022159f
C1154 VTAIL.n258 VSUBS 0.022159f
C1155 VTAIL.n259 VSUBS 0.011907f
C1156 VTAIL.n260 VSUBS 0.012607f
C1157 VTAIL.n261 VSUBS 0.028144f
C1158 VTAIL.n262 VSUBS 0.028144f
C1159 VTAIL.n263 VSUBS 0.012607f
C1160 VTAIL.n264 VSUBS 0.011907f
C1161 VTAIL.n265 VSUBS 0.022159f
C1162 VTAIL.n266 VSUBS 0.022159f
C1163 VTAIL.n267 VSUBS 0.011907f
C1164 VTAIL.n268 VSUBS 0.012607f
C1165 VTAIL.n269 VSUBS 0.028144f
C1166 VTAIL.n270 VSUBS 0.028144f
C1167 VTAIL.n271 VSUBS 0.012607f
C1168 VTAIL.n272 VSUBS 0.011907f
C1169 VTAIL.n273 VSUBS 0.022159f
C1170 VTAIL.n274 VSUBS 0.022159f
C1171 VTAIL.n275 VSUBS 0.011907f
C1172 VTAIL.n276 VSUBS 0.012607f
C1173 VTAIL.n277 VSUBS 0.028144f
C1174 VTAIL.n278 VSUBS 0.028144f
C1175 VTAIL.n279 VSUBS 0.012607f
C1176 VTAIL.n280 VSUBS 0.011907f
C1177 VTAIL.n281 VSUBS 0.022159f
C1178 VTAIL.n282 VSUBS 0.022159f
C1179 VTAIL.n283 VSUBS 0.011907f
C1180 VTAIL.n284 VSUBS 0.012607f
C1181 VTAIL.n285 VSUBS 0.028144f
C1182 VTAIL.n286 VSUBS 0.028144f
C1183 VTAIL.n287 VSUBS 0.028144f
C1184 VTAIL.n288 VSUBS 0.012607f
C1185 VTAIL.n289 VSUBS 0.011907f
C1186 VTAIL.n290 VSUBS 0.022159f
C1187 VTAIL.n291 VSUBS 0.022159f
C1188 VTAIL.n292 VSUBS 0.011907f
C1189 VTAIL.n293 VSUBS 0.012257f
C1190 VTAIL.n294 VSUBS 0.012257f
C1191 VTAIL.n295 VSUBS 0.028144f
C1192 VTAIL.n296 VSUBS 0.028144f
C1193 VTAIL.n297 VSUBS 0.012607f
C1194 VTAIL.n298 VSUBS 0.011907f
C1195 VTAIL.n299 VSUBS 0.022159f
C1196 VTAIL.n300 VSUBS 0.022159f
C1197 VTAIL.n301 VSUBS 0.011907f
C1198 VTAIL.n302 VSUBS 0.012607f
C1199 VTAIL.n303 VSUBS 0.028144f
C1200 VTAIL.n304 VSUBS 0.028144f
C1201 VTAIL.n305 VSUBS 0.012607f
C1202 VTAIL.n306 VSUBS 0.011907f
C1203 VTAIL.n307 VSUBS 0.022159f
C1204 VTAIL.n308 VSUBS 0.022159f
C1205 VTAIL.n309 VSUBS 0.011907f
C1206 VTAIL.n310 VSUBS 0.012607f
C1207 VTAIL.n311 VSUBS 0.028144f
C1208 VTAIL.n312 VSUBS 0.068138f
C1209 VTAIL.n313 VSUBS 0.012607f
C1210 VTAIL.n314 VSUBS 0.011907f
C1211 VTAIL.n315 VSUBS 0.050311f
C1212 VTAIL.n316 VSUBS 0.034238f
C1213 VTAIL.n317 VSUBS 1.87237f
C1214 VTAIL.n318 VSUBS 0.024349f
C1215 VTAIL.n319 VSUBS 0.022159f
C1216 VTAIL.n320 VSUBS 0.011907f
C1217 VTAIL.n321 VSUBS 0.028144f
C1218 VTAIL.n322 VSUBS 0.012607f
C1219 VTAIL.n323 VSUBS 0.022159f
C1220 VTAIL.n324 VSUBS 0.011907f
C1221 VTAIL.n325 VSUBS 0.028144f
C1222 VTAIL.n326 VSUBS 0.012607f
C1223 VTAIL.n327 VSUBS 0.022159f
C1224 VTAIL.n328 VSUBS 0.011907f
C1225 VTAIL.n329 VSUBS 0.028144f
C1226 VTAIL.n330 VSUBS 0.012607f
C1227 VTAIL.n331 VSUBS 0.022159f
C1228 VTAIL.n332 VSUBS 0.011907f
C1229 VTAIL.n333 VSUBS 0.028144f
C1230 VTAIL.n334 VSUBS 0.028144f
C1231 VTAIL.n335 VSUBS 0.012607f
C1232 VTAIL.n336 VSUBS 0.022159f
C1233 VTAIL.n337 VSUBS 0.011907f
C1234 VTAIL.n338 VSUBS 0.028144f
C1235 VTAIL.n339 VSUBS 0.012607f
C1236 VTAIL.n340 VSUBS 0.022159f
C1237 VTAIL.n341 VSUBS 0.011907f
C1238 VTAIL.n342 VSUBS 0.028144f
C1239 VTAIL.n343 VSUBS 0.012607f
C1240 VTAIL.n344 VSUBS 0.022159f
C1241 VTAIL.n345 VSUBS 0.011907f
C1242 VTAIL.n346 VSUBS 0.028144f
C1243 VTAIL.n347 VSUBS 0.012607f
C1244 VTAIL.n348 VSUBS 0.022159f
C1245 VTAIL.n349 VSUBS 0.011907f
C1246 VTAIL.n350 VSUBS 0.028144f
C1247 VTAIL.n351 VSUBS 0.012607f
C1248 VTAIL.n352 VSUBS 0.181886f
C1249 VTAIL.t3 VSUBS 0.060467f
C1250 VTAIL.n353 VSUBS 0.021108f
C1251 VTAIL.n354 VSUBS 0.017904f
C1252 VTAIL.n355 VSUBS 0.011907f
C1253 VTAIL.n356 VSUBS 1.81021f
C1254 VTAIL.n357 VSUBS 0.022159f
C1255 VTAIL.n358 VSUBS 0.011907f
C1256 VTAIL.n359 VSUBS 0.012607f
C1257 VTAIL.n360 VSUBS 0.028144f
C1258 VTAIL.n361 VSUBS 0.028144f
C1259 VTAIL.n362 VSUBS 0.012607f
C1260 VTAIL.n363 VSUBS 0.011907f
C1261 VTAIL.n364 VSUBS 0.022159f
C1262 VTAIL.n365 VSUBS 0.022159f
C1263 VTAIL.n366 VSUBS 0.011907f
C1264 VTAIL.n367 VSUBS 0.012607f
C1265 VTAIL.n368 VSUBS 0.028144f
C1266 VTAIL.n369 VSUBS 0.028144f
C1267 VTAIL.n370 VSUBS 0.012607f
C1268 VTAIL.n371 VSUBS 0.011907f
C1269 VTAIL.n372 VSUBS 0.022159f
C1270 VTAIL.n373 VSUBS 0.022159f
C1271 VTAIL.n374 VSUBS 0.011907f
C1272 VTAIL.n375 VSUBS 0.012607f
C1273 VTAIL.n376 VSUBS 0.028144f
C1274 VTAIL.n377 VSUBS 0.028144f
C1275 VTAIL.n378 VSUBS 0.012607f
C1276 VTAIL.n379 VSUBS 0.011907f
C1277 VTAIL.n380 VSUBS 0.022159f
C1278 VTAIL.n381 VSUBS 0.022159f
C1279 VTAIL.n382 VSUBS 0.011907f
C1280 VTAIL.n383 VSUBS 0.012607f
C1281 VTAIL.n384 VSUBS 0.028144f
C1282 VTAIL.n385 VSUBS 0.028144f
C1283 VTAIL.n386 VSUBS 0.012607f
C1284 VTAIL.n387 VSUBS 0.011907f
C1285 VTAIL.n388 VSUBS 0.022159f
C1286 VTAIL.n389 VSUBS 0.022159f
C1287 VTAIL.n390 VSUBS 0.011907f
C1288 VTAIL.n391 VSUBS 0.012607f
C1289 VTAIL.n392 VSUBS 0.028144f
C1290 VTAIL.n393 VSUBS 0.028144f
C1291 VTAIL.n394 VSUBS 0.012607f
C1292 VTAIL.n395 VSUBS 0.011907f
C1293 VTAIL.n396 VSUBS 0.022159f
C1294 VTAIL.n397 VSUBS 0.022159f
C1295 VTAIL.n398 VSUBS 0.011907f
C1296 VTAIL.n399 VSUBS 0.012257f
C1297 VTAIL.n400 VSUBS 0.012257f
C1298 VTAIL.n401 VSUBS 0.028144f
C1299 VTAIL.n402 VSUBS 0.028144f
C1300 VTAIL.n403 VSUBS 0.012607f
C1301 VTAIL.n404 VSUBS 0.011907f
C1302 VTAIL.n405 VSUBS 0.022159f
C1303 VTAIL.n406 VSUBS 0.022159f
C1304 VTAIL.n407 VSUBS 0.011907f
C1305 VTAIL.n408 VSUBS 0.012607f
C1306 VTAIL.n409 VSUBS 0.028144f
C1307 VTAIL.n410 VSUBS 0.028144f
C1308 VTAIL.n411 VSUBS 0.012607f
C1309 VTAIL.n412 VSUBS 0.011907f
C1310 VTAIL.n413 VSUBS 0.022159f
C1311 VTAIL.n414 VSUBS 0.022159f
C1312 VTAIL.n415 VSUBS 0.011907f
C1313 VTAIL.n416 VSUBS 0.012607f
C1314 VTAIL.n417 VSUBS 0.028144f
C1315 VTAIL.n418 VSUBS 0.068138f
C1316 VTAIL.n419 VSUBS 0.012607f
C1317 VTAIL.n420 VSUBS 0.011907f
C1318 VTAIL.n421 VSUBS 0.050311f
C1319 VTAIL.n422 VSUBS 0.034238f
C1320 VTAIL.n423 VSUBS 1.87237f
C1321 VTAIL.n424 VSUBS 0.024349f
C1322 VTAIL.n425 VSUBS 0.022159f
C1323 VTAIL.n426 VSUBS 0.011907f
C1324 VTAIL.n427 VSUBS 0.028144f
C1325 VTAIL.n428 VSUBS 0.012607f
C1326 VTAIL.n429 VSUBS 0.022159f
C1327 VTAIL.n430 VSUBS 0.011907f
C1328 VTAIL.n431 VSUBS 0.028144f
C1329 VTAIL.n432 VSUBS 0.012607f
C1330 VTAIL.n433 VSUBS 0.022159f
C1331 VTAIL.n434 VSUBS 0.011907f
C1332 VTAIL.n435 VSUBS 0.028144f
C1333 VTAIL.n436 VSUBS 0.012607f
C1334 VTAIL.n437 VSUBS 0.022159f
C1335 VTAIL.n438 VSUBS 0.011907f
C1336 VTAIL.n439 VSUBS 0.028144f
C1337 VTAIL.n440 VSUBS 0.028144f
C1338 VTAIL.n441 VSUBS 0.012607f
C1339 VTAIL.n442 VSUBS 0.022159f
C1340 VTAIL.n443 VSUBS 0.011907f
C1341 VTAIL.n444 VSUBS 0.028144f
C1342 VTAIL.n445 VSUBS 0.012607f
C1343 VTAIL.n446 VSUBS 0.022159f
C1344 VTAIL.n447 VSUBS 0.011907f
C1345 VTAIL.n448 VSUBS 0.028144f
C1346 VTAIL.n449 VSUBS 0.012607f
C1347 VTAIL.n450 VSUBS 0.022159f
C1348 VTAIL.n451 VSUBS 0.011907f
C1349 VTAIL.n452 VSUBS 0.028144f
C1350 VTAIL.n453 VSUBS 0.012607f
C1351 VTAIL.n454 VSUBS 0.022159f
C1352 VTAIL.n455 VSUBS 0.011907f
C1353 VTAIL.n456 VSUBS 0.028144f
C1354 VTAIL.n457 VSUBS 0.012607f
C1355 VTAIL.n458 VSUBS 0.181886f
C1356 VTAIL.t0 VSUBS 0.060467f
C1357 VTAIL.n459 VSUBS 0.021108f
C1358 VTAIL.n460 VSUBS 0.017904f
C1359 VTAIL.n461 VSUBS 0.011907f
C1360 VTAIL.n462 VSUBS 1.81021f
C1361 VTAIL.n463 VSUBS 0.022159f
C1362 VTAIL.n464 VSUBS 0.011907f
C1363 VTAIL.n465 VSUBS 0.012607f
C1364 VTAIL.n466 VSUBS 0.028144f
C1365 VTAIL.n467 VSUBS 0.028144f
C1366 VTAIL.n468 VSUBS 0.012607f
C1367 VTAIL.n469 VSUBS 0.011907f
C1368 VTAIL.n470 VSUBS 0.022159f
C1369 VTAIL.n471 VSUBS 0.022159f
C1370 VTAIL.n472 VSUBS 0.011907f
C1371 VTAIL.n473 VSUBS 0.012607f
C1372 VTAIL.n474 VSUBS 0.028144f
C1373 VTAIL.n475 VSUBS 0.028144f
C1374 VTAIL.n476 VSUBS 0.012607f
C1375 VTAIL.n477 VSUBS 0.011907f
C1376 VTAIL.n478 VSUBS 0.022159f
C1377 VTAIL.n479 VSUBS 0.022159f
C1378 VTAIL.n480 VSUBS 0.011907f
C1379 VTAIL.n481 VSUBS 0.012607f
C1380 VTAIL.n482 VSUBS 0.028144f
C1381 VTAIL.n483 VSUBS 0.028144f
C1382 VTAIL.n484 VSUBS 0.012607f
C1383 VTAIL.n485 VSUBS 0.011907f
C1384 VTAIL.n486 VSUBS 0.022159f
C1385 VTAIL.n487 VSUBS 0.022159f
C1386 VTAIL.n488 VSUBS 0.011907f
C1387 VTAIL.n489 VSUBS 0.012607f
C1388 VTAIL.n490 VSUBS 0.028144f
C1389 VTAIL.n491 VSUBS 0.028144f
C1390 VTAIL.n492 VSUBS 0.012607f
C1391 VTAIL.n493 VSUBS 0.011907f
C1392 VTAIL.n494 VSUBS 0.022159f
C1393 VTAIL.n495 VSUBS 0.022159f
C1394 VTAIL.n496 VSUBS 0.011907f
C1395 VTAIL.n497 VSUBS 0.012607f
C1396 VTAIL.n498 VSUBS 0.028144f
C1397 VTAIL.n499 VSUBS 0.028144f
C1398 VTAIL.n500 VSUBS 0.012607f
C1399 VTAIL.n501 VSUBS 0.011907f
C1400 VTAIL.n502 VSUBS 0.022159f
C1401 VTAIL.n503 VSUBS 0.022159f
C1402 VTAIL.n504 VSUBS 0.011907f
C1403 VTAIL.n505 VSUBS 0.012257f
C1404 VTAIL.n506 VSUBS 0.012257f
C1405 VTAIL.n507 VSUBS 0.028144f
C1406 VTAIL.n508 VSUBS 0.028144f
C1407 VTAIL.n509 VSUBS 0.012607f
C1408 VTAIL.n510 VSUBS 0.011907f
C1409 VTAIL.n511 VSUBS 0.022159f
C1410 VTAIL.n512 VSUBS 0.022159f
C1411 VTAIL.n513 VSUBS 0.011907f
C1412 VTAIL.n514 VSUBS 0.012607f
C1413 VTAIL.n515 VSUBS 0.028144f
C1414 VTAIL.n516 VSUBS 0.028144f
C1415 VTAIL.n517 VSUBS 0.012607f
C1416 VTAIL.n518 VSUBS 0.011907f
C1417 VTAIL.n519 VSUBS 0.022159f
C1418 VTAIL.n520 VSUBS 0.022159f
C1419 VTAIL.n521 VSUBS 0.011907f
C1420 VTAIL.n522 VSUBS 0.012607f
C1421 VTAIL.n523 VSUBS 0.028144f
C1422 VTAIL.n524 VSUBS 0.068138f
C1423 VTAIL.n525 VSUBS 0.012607f
C1424 VTAIL.n526 VSUBS 0.011907f
C1425 VTAIL.n527 VSUBS 0.050311f
C1426 VTAIL.n528 VSUBS 0.034238f
C1427 VTAIL.n529 VSUBS 0.245847f
C1428 VTAIL.n530 VSUBS 0.024349f
C1429 VTAIL.n531 VSUBS 0.022159f
C1430 VTAIL.n532 VSUBS 0.011907f
C1431 VTAIL.n533 VSUBS 0.028144f
C1432 VTAIL.n534 VSUBS 0.012607f
C1433 VTAIL.n535 VSUBS 0.022159f
C1434 VTAIL.n536 VSUBS 0.011907f
C1435 VTAIL.n537 VSUBS 0.028144f
C1436 VTAIL.n538 VSUBS 0.012607f
C1437 VTAIL.n539 VSUBS 0.022159f
C1438 VTAIL.n540 VSUBS 0.011907f
C1439 VTAIL.n541 VSUBS 0.028144f
C1440 VTAIL.n542 VSUBS 0.012607f
C1441 VTAIL.n543 VSUBS 0.022159f
C1442 VTAIL.n544 VSUBS 0.011907f
C1443 VTAIL.n545 VSUBS 0.028144f
C1444 VTAIL.n546 VSUBS 0.028144f
C1445 VTAIL.n547 VSUBS 0.012607f
C1446 VTAIL.n548 VSUBS 0.022159f
C1447 VTAIL.n549 VSUBS 0.011907f
C1448 VTAIL.n550 VSUBS 0.028144f
C1449 VTAIL.n551 VSUBS 0.012607f
C1450 VTAIL.n552 VSUBS 0.022159f
C1451 VTAIL.n553 VSUBS 0.011907f
C1452 VTAIL.n554 VSUBS 0.028144f
C1453 VTAIL.n555 VSUBS 0.012607f
C1454 VTAIL.n556 VSUBS 0.022159f
C1455 VTAIL.n557 VSUBS 0.011907f
C1456 VTAIL.n558 VSUBS 0.028144f
C1457 VTAIL.n559 VSUBS 0.012607f
C1458 VTAIL.n560 VSUBS 0.022159f
C1459 VTAIL.n561 VSUBS 0.011907f
C1460 VTAIL.n562 VSUBS 0.028144f
C1461 VTAIL.n563 VSUBS 0.012607f
C1462 VTAIL.n564 VSUBS 0.181886f
C1463 VTAIL.t6 VSUBS 0.060467f
C1464 VTAIL.n565 VSUBS 0.021108f
C1465 VTAIL.n566 VSUBS 0.017904f
C1466 VTAIL.n567 VSUBS 0.011907f
C1467 VTAIL.n568 VSUBS 1.81021f
C1468 VTAIL.n569 VSUBS 0.022159f
C1469 VTAIL.n570 VSUBS 0.011907f
C1470 VTAIL.n571 VSUBS 0.012607f
C1471 VTAIL.n572 VSUBS 0.028144f
C1472 VTAIL.n573 VSUBS 0.028144f
C1473 VTAIL.n574 VSUBS 0.012607f
C1474 VTAIL.n575 VSUBS 0.011907f
C1475 VTAIL.n576 VSUBS 0.022159f
C1476 VTAIL.n577 VSUBS 0.022159f
C1477 VTAIL.n578 VSUBS 0.011907f
C1478 VTAIL.n579 VSUBS 0.012607f
C1479 VTAIL.n580 VSUBS 0.028144f
C1480 VTAIL.n581 VSUBS 0.028144f
C1481 VTAIL.n582 VSUBS 0.012607f
C1482 VTAIL.n583 VSUBS 0.011907f
C1483 VTAIL.n584 VSUBS 0.022159f
C1484 VTAIL.n585 VSUBS 0.022159f
C1485 VTAIL.n586 VSUBS 0.011907f
C1486 VTAIL.n587 VSUBS 0.012607f
C1487 VTAIL.n588 VSUBS 0.028144f
C1488 VTAIL.n589 VSUBS 0.028144f
C1489 VTAIL.n590 VSUBS 0.012607f
C1490 VTAIL.n591 VSUBS 0.011907f
C1491 VTAIL.n592 VSUBS 0.022159f
C1492 VTAIL.n593 VSUBS 0.022159f
C1493 VTAIL.n594 VSUBS 0.011907f
C1494 VTAIL.n595 VSUBS 0.012607f
C1495 VTAIL.n596 VSUBS 0.028144f
C1496 VTAIL.n597 VSUBS 0.028144f
C1497 VTAIL.n598 VSUBS 0.012607f
C1498 VTAIL.n599 VSUBS 0.011907f
C1499 VTAIL.n600 VSUBS 0.022159f
C1500 VTAIL.n601 VSUBS 0.022159f
C1501 VTAIL.n602 VSUBS 0.011907f
C1502 VTAIL.n603 VSUBS 0.012607f
C1503 VTAIL.n604 VSUBS 0.028144f
C1504 VTAIL.n605 VSUBS 0.028144f
C1505 VTAIL.n606 VSUBS 0.012607f
C1506 VTAIL.n607 VSUBS 0.011907f
C1507 VTAIL.n608 VSUBS 0.022159f
C1508 VTAIL.n609 VSUBS 0.022159f
C1509 VTAIL.n610 VSUBS 0.011907f
C1510 VTAIL.n611 VSUBS 0.012257f
C1511 VTAIL.n612 VSUBS 0.012257f
C1512 VTAIL.n613 VSUBS 0.028144f
C1513 VTAIL.n614 VSUBS 0.028144f
C1514 VTAIL.n615 VSUBS 0.012607f
C1515 VTAIL.n616 VSUBS 0.011907f
C1516 VTAIL.n617 VSUBS 0.022159f
C1517 VTAIL.n618 VSUBS 0.022159f
C1518 VTAIL.n619 VSUBS 0.011907f
C1519 VTAIL.n620 VSUBS 0.012607f
C1520 VTAIL.n621 VSUBS 0.028144f
C1521 VTAIL.n622 VSUBS 0.028144f
C1522 VTAIL.n623 VSUBS 0.012607f
C1523 VTAIL.n624 VSUBS 0.011907f
C1524 VTAIL.n625 VSUBS 0.022159f
C1525 VTAIL.n626 VSUBS 0.022159f
C1526 VTAIL.n627 VSUBS 0.011907f
C1527 VTAIL.n628 VSUBS 0.012607f
C1528 VTAIL.n629 VSUBS 0.028144f
C1529 VTAIL.n630 VSUBS 0.068138f
C1530 VTAIL.n631 VSUBS 0.012607f
C1531 VTAIL.n632 VSUBS 0.011907f
C1532 VTAIL.n633 VSUBS 0.050311f
C1533 VTAIL.n634 VSUBS 0.034238f
C1534 VTAIL.n635 VSUBS 0.245847f
C1535 VTAIL.n636 VSUBS 0.024349f
C1536 VTAIL.n637 VSUBS 0.022159f
C1537 VTAIL.n638 VSUBS 0.011907f
C1538 VTAIL.n639 VSUBS 0.028144f
C1539 VTAIL.n640 VSUBS 0.012607f
C1540 VTAIL.n641 VSUBS 0.022159f
C1541 VTAIL.n642 VSUBS 0.011907f
C1542 VTAIL.n643 VSUBS 0.028144f
C1543 VTAIL.n644 VSUBS 0.012607f
C1544 VTAIL.n645 VSUBS 0.022159f
C1545 VTAIL.n646 VSUBS 0.011907f
C1546 VTAIL.n647 VSUBS 0.028144f
C1547 VTAIL.n648 VSUBS 0.012607f
C1548 VTAIL.n649 VSUBS 0.022159f
C1549 VTAIL.n650 VSUBS 0.011907f
C1550 VTAIL.n651 VSUBS 0.028144f
C1551 VTAIL.n652 VSUBS 0.028144f
C1552 VTAIL.n653 VSUBS 0.012607f
C1553 VTAIL.n654 VSUBS 0.022159f
C1554 VTAIL.n655 VSUBS 0.011907f
C1555 VTAIL.n656 VSUBS 0.028144f
C1556 VTAIL.n657 VSUBS 0.012607f
C1557 VTAIL.n658 VSUBS 0.022159f
C1558 VTAIL.n659 VSUBS 0.011907f
C1559 VTAIL.n660 VSUBS 0.028144f
C1560 VTAIL.n661 VSUBS 0.012607f
C1561 VTAIL.n662 VSUBS 0.022159f
C1562 VTAIL.n663 VSUBS 0.011907f
C1563 VTAIL.n664 VSUBS 0.028144f
C1564 VTAIL.n665 VSUBS 0.012607f
C1565 VTAIL.n666 VSUBS 0.022159f
C1566 VTAIL.n667 VSUBS 0.011907f
C1567 VTAIL.n668 VSUBS 0.028144f
C1568 VTAIL.n669 VSUBS 0.012607f
C1569 VTAIL.n670 VSUBS 0.181886f
C1570 VTAIL.t4 VSUBS 0.060467f
C1571 VTAIL.n671 VSUBS 0.021108f
C1572 VTAIL.n672 VSUBS 0.017904f
C1573 VTAIL.n673 VSUBS 0.011907f
C1574 VTAIL.n674 VSUBS 1.81021f
C1575 VTAIL.n675 VSUBS 0.022159f
C1576 VTAIL.n676 VSUBS 0.011907f
C1577 VTAIL.n677 VSUBS 0.012607f
C1578 VTAIL.n678 VSUBS 0.028144f
C1579 VTAIL.n679 VSUBS 0.028144f
C1580 VTAIL.n680 VSUBS 0.012607f
C1581 VTAIL.n681 VSUBS 0.011907f
C1582 VTAIL.n682 VSUBS 0.022159f
C1583 VTAIL.n683 VSUBS 0.022159f
C1584 VTAIL.n684 VSUBS 0.011907f
C1585 VTAIL.n685 VSUBS 0.012607f
C1586 VTAIL.n686 VSUBS 0.028144f
C1587 VTAIL.n687 VSUBS 0.028144f
C1588 VTAIL.n688 VSUBS 0.012607f
C1589 VTAIL.n689 VSUBS 0.011907f
C1590 VTAIL.n690 VSUBS 0.022159f
C1591 VTAIL.n691 VSUBS 0.022159f
C1592 VTAIL.n692 VSUBS 0.011907f
C1593 VTAIL.n693 VSUBS 0.012607f
C1594 VTAIL.n694 VSUBS 0.028144f
C1595 VTAIL.n695 VSUBS 0.028144f
C1596 VTAIL.n696 VSUBS 0.012607f
C1597 VTAIL.n697 VSUBS 0.011907f
C1598 VTAIL.n698 VSUBS 0.022159f
C1599 VTAIL.n699 VSUBS 0.022159f
C1600 VTAIL.n700 VSUBS 0.011907f
C1601 VTAIL.n701 VSUBS 0.012607f
C1602 VTAIL.n702 VSUBS 0.028144f
C1603 VTAIL.n703 VSUBS 0.028144f
C1604 VTAIL.n704 VSUBS 0.012607f
C1605 VTAIL.n705 VSUBS 0.011907f
C1606 VTAIL.n706 VSUBS 0.022159f
C1607 VTAIL.n707 VSUBS 0.022159f
C1608 VTAIL.n708 VSUBS 0.011907f
C1609 VTAIL.n709 VSUBS 0.012607f
C1610 VTAIL.n710 VSUBS 0.028144f
C1611 VTAIL.n711 VSUBS 0.028144f
C1612 VTAIL.n712 VSUBS 0.012607f
C1613 VTAIL.n713 VSUBS 0.011907f
C1614 VTAIL.n714 VSUBS 0.022159f
C1615 VTAIL.n715 VSUBS 0.022159f
C1616 VTAIL.n716 VSUBS 0.011907f
C1617 VTAIL.n717 VSUBS 0.012257f
C1618 VTAIL.n718 VSUBS 0.012257f
C1619 VTAIL.n719 VSUBS 0.028144f
C1620 VTAIL.n720 VSUBS 0.028144f
C1621 VTAIL.n721 VSUBS 0.012607f
C1622 VTAIL.n722 VSUBS 0.011907f
C1623 VTAIL.n723 VSUBS 0.022159f
C1624 VTAIL.n724 VSUBS 0.022159f
C1625 VTAIL.n725 VSUBS 0.011907f
C1626 VTAIL.n726 VSUBS 0.012607f
C1627 VTAIL.n727 VSUBS 0.028144f
C1628 VTAIL.n728 VSUBS 0.028144f
C1629 VTAIL.n729 VSUBS 0.012607f
C1630 VTAIL.n730 VSUBS 0.011907f
C1631 VTAIL.n731 VSUBS 0.022159f
C1632 VTAIL.n732 VSUBS 0.022159f
C1633 VTAIL.n733 VSUBS 0.011907f
C1634 VTAIL.n734 VSUBS 0.012607f
C1635 VTAIL.n735 VSUBS 0.028144f
C1636 VTAIL.n736 VSUBS 0.068138f
C1637 VTAIL.n737 VSUBS 0.012607f
C1638 VTAIL.n738 VSUBS 0.011907f
C1639 VTAIL.n739 VSUBS 0.050311f
C1640 VTAIL.n740 VSUBS 0.034238f
C1641 VTAIL.n741 VSUBS 1.87237f
C1642 VTAIL.n742 VSUBS 0.024349f
C1643 VTAIL.n743 VSUBS 0.022159f
C1644 VTAIL.n744 VSUBS 0.011907f
C1645 VTAIL.n745 VSUBS 0.028144f
C1646 VTAIL.n746 VSUBS 0.012607f
C1647 VTAIL.n747 VSUBS 0.022159f
C1648 VTAIL.n748 VSUBS 0.011907f
C1649 VTAIL.n749 VSUBS 0.028144f
C1650 VTAIL.n750 VSUBS 0.012607f
C1651 VTAIL.n751 VSUBS 0.022159f
C1652 VTAIL.n752 VSUBS 0.011907f
C1653 VTAIL.n753 VSUBS 0.028144f
C1654 VTAIL.n754 VSUBS 0.012607f
C1655 VTAIL.n755 VSUBS 0.022159f
C1656 VTAIL.n756 VSUBS 0.011907f
C1657 VTAIL.n757 VSUBS 0.028144f
C1658 VTAIL.n758 VSUBS 0.012607f
C1659 VTAIL.n759 VSUBS 0.022159f
C1660 VTAIL.n760 VSUBS 0.011907f
C1661 VTAIL.n761 VSUBS 0.028144f
C1662 VTAIL.n762 VSUBS 0.012607f
C1663 VTAIL.n763 VSUBS 0.022159f
C1664 VTAIL.n764 VSUBS 0.011907f
C1665 VTAIL.n765 VSUBS 0.028144f
C1666 VTAIL.n766 VSUBS 0.012607f
C1667 VTAIL.n767 VSUBS 0.022159f
C1668 VTAIL.n768 VSUBS 0.011907f
C1669 VTAIL.n769 VSUBS 0.028144f
C1670 VTAIL.n770 VSUBS 0.012607f
C1671 VTAIL.n771 VSUBS 0.022159f
C1672 VTAIL.n772 VSUBS 0.011907f
C1673 VTAIL.n773 VSUBS 0.028144f
C1674 VTAIL.n774 VSUBS 0.012607f
C1675 VTAIL.n775 VSUBS 0.181886f
C1676 VTAIL.t2 VSUBS 0.060467f
C1677 VTAIL.n776 VSUBS 0.021108f
C1678 VTAIL.n777 VSUBS 0.017904f
C1679 VTAIL.n778 VSUBS 0.011907f
C1680 VTAIL.n779 VSUBS 1.81021f
C1681 VTAIL.n780 VSUBS 0.022159f
C1682 VTAIL.n781 VSUBS 0.011907f
C1683 VTAIL.n782 VSUBS 0.012607f
C1684 VTAIL.n783 VSUBS 0.028144f
C1685 VTAIL.n784 VSUBS 0.028144f
C1686 VTAIL.n785 VSUBS 0.012607f
C1687 VTAIL.n786 VSUBS 0.011907f
C1688 VTAIL.n787 VSUBS 0.022159f
C1689 VTAIL.n788 VSUBS 0.022159f
C1690 VTAIL.n789 VSUBS 0.011907f
C1691 VTAIL.n790 VSUBS 0.012607f
C1692 VTAIL.n791 VSUBS 0.028144f
C1693 VTAIL.n792 VSUBS 0.028144f
C1694 VTAIL.n793 VSUBS 0.012607f
C1695 VTAIL.n794 VSUBS 0.011907f
C1696 VTAIL.n795 VSUBS 0.022159f
C1697 VTAIL.n796 VSUBS 0.022159f
C1698 VTAIL.n797 VSUBS 0.011907f
C1699 VTAIL.n798 VSUBS 0.012607f
C1700 VTAIL.n799 VSUBS 0.028144f
C1701 VTAIL.n800 VSUBS 0.028144f
C1702 VTAIL.n801 VSUBS 0.012607f
C1703 VTAIL.n802 VSUBS 0.011907f
C1704 VTAIL.n803 VSUBS 0.022159f
C1705 VTAIL.n804 VSUBS 0.022159f
C1706 VTAIL.n805 VSUBS 0.011907f
C1707 VTAIL.n806 VSUBS 0.012607f
C1708 VTAIL.n807 VSUBS 0.028144f
C1709 VTAIL.n808 VSUBS 0.028144f
C1710 VTAIL.n809 VSUBS 0.012607f
C1711 VTAIL.n810 VSUBS 0.011907f
C1712 VTAIL.n811 VSUBS 0.022159f
C1713 VTAIL.n812 VSUBS 0.022159f
C1714 VTAIL.n813 VSUBS 0.011907f
C1715 VTAIL.n814 VSUBS 0.012607f
C1716 VTAIL.n815 VSUBS 0.028144f
C1717 VTAIL.n816 VSUBS 0.028144f
C1718 VTAIL.n817 VSUBS 0.028144f
C1719 VTAIL.n818 VSUBS 0.012607f
C1720 VTAIL.n819 VSUBS 0.011907f
C1721 VTAIL.n820 VSUBS 0.022159f
C1722 VTAIL.n821 VSUBS 0.022159f
C1723 VTAIL.n822 VSUBS 0.011907f
C1724 VTAIL.n823 VSUBS 0.012257f
C1725 VTAIL.n824 VSUBS 0.012257f
C1726 VTAIL.n825 VSUBS 0.028144f
C1727 VTAIL.n826 VSUBS 0.028144f
C1728 VTAIL.n827 VSUBS 0.012607f
C1729 VTAIL.n828 VSUBS 0.011907f
C1730 VTAIL.n829 VSUBS 0.022159f
C1731 VTAIL.n830 VSUBS 0.022159f
C1732 VTAIL.n831 VSUBS 0.011907f
C1733 VTAIL.n832 VSUBS 0.012607f
C1734 VTAIL.n833 VSUBS 0.028144f
C1735 VTAIL.n834 VSUBS 0.028144f
C1736 VTAIL.n835 VSUBS 0.012607f
C1737 VTAIL.n836 VSUBS 0.011907f
C1738 VTAIL.n837 VSUBS 0.022159f
C1739 VTAIL.n838 VSUBS 0.022159f
C1740 VTAIL.n839 VSUBS 0.011907f
C1741 VTAIL.n840 VSUBS 0.012607f
C1742 VTAIL.n841 VSUBS 0.028144f
C1743 VTAIL.n842 VSUBS 0.068138f
C1744 VTAIL.n843 VSUBS 0.012607f
C1745 VTAIL.n844 VSUBS 0.011907f
C1746 VTAIL.n845 VSUBS 0.050311f
C1747 VTAIL.n846 VSUBS 0.034238f
C1748 VTAIL.n847 VSUBS 1.77127f
C1749 VDD1.t0 VSUBS 0.398461f
C1750 VDD1.t3 VSUBS 0.398461f
C1751 VDD1.n0 VSUBS 3.32678f
C1752 VDD1.t1 VSUBS 0.398461f
C1753 VDD1.t2 VSUBS 0.398461f
C1754 VDD1.n1 VSUBS 4.37516f
C1755 VP.n0 VSUBS 0.03789f
C1756 VP.t2 VSUBS 4.22384f
C1757 VP.n1 VSUBS 0.05712f
C1758 VP.n2 VSUBS 0.02874f
C1759 VP.n3 VSUBS 0.031084f
C1760 VP.t3 VSUBS 4.51257f
C1761 VP.t1 VSUBS 4.5199f
C1762 VP.n4 VSUBS 4.73855f
C1763 VP.t0 VSUBS 4.22384f
C1764 VP.n5 VSUBS 1.55446f
C1765 VP.n6 VSUBS 1.8563f
C1766 VP.n7 VSUBS 0.03789f
C1767 VP.n8 VSUBS 0.02874f
C1768 VP.n9 VSUBS 0.053564f
C1769 VP.n10 VSUBS 0.05712f
C1770 VP.n11 VSUBS 0.023233f
C1771 VP.n12 VSUBS 0.02874f
C1772 VP.n13 VSUBS 0.02874f
C1773 VP.n14 VSUBS 0.02874f
C1774 VP.n15 VSUBS 0.053564f
C1775 VP.n16 VSUBS 0.031084f
C1776 VP.n17 VSUBS 1.55446f
C1777 VP.n18 VSUBS 0.053344f
.ends

