* NGSPICE file created from diff_pair_sample_0871.ext - technology: sky130A

.subckt diff_pair_sample_0871 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X1 B.t22 B.t20 B.t21 B.t14 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=0 ps=0 w=12.92 l=1.49
X2 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X3 B.t19 B.t17 B.t18 B.t10 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=0 ps=0 w=12.92 l=1.49
X4 VDD1.t8 VP.t1 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=2.1318 ps=13.25 w=12.92 l=1.49
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=0 ps=0 w=12.92 l=1.49
X6 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X7 VDD1.t7 VP.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=2.1318 ps=13.25 w=12.92 l=1.49
X8 VDD2.t7 VN.t2 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=2.1318 ps=13.25 w=12.92 l=1.49
X9 VDD2.t6 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=2.1318 ps=13.25 w=12.92 l=1.49
X10 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X11 VTAIL.t16 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X12 VDD1.t5 VP.t4 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=5.0388 ps=26.62 w=12.92 l=1.49
X13 VTAIL.t2 VN.t5 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X14 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.0388 pd=26.62 as=0 ps=0 w=12.92 l=1.49
X15 VDD2.t3 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X16 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=5.0388 ps=26.62 w=12.92 l=1.49
X17 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X18 VDD1.t4 VP.t5 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X19 VDD1.t3 VP.t6 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=5.0388 ps=26.62 w=12.92 l=1.49
X20 VTAIL.t13 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X21 VDD2.t0 VN.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=5.0388 ps=26.62 w=12.92 l=1.49
X22 VTAIL.t14 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
X23 VTAIL.t11 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1318 pd=13.25 as=2.1318 ps=13.25 w=12.92 l=1.49
R0 VP.n15 VP.t2 241.106
R1 VP.n48 VP.t5 208.976
R2 VP.n35 VP.t1 208.976
R3 VP.n41 VP.t9 208.976
R4 VP.n54 VP.t8 208.976
R5 VP.n61 VP.t4 208.976
R6 VP.n20 VP.t0 208.976
R7 VP.n33 VP.t6 208.976
R8 VP.n26 VP.t3 208.976
R9 VP.n14 VP.t7 208.976
R10 VP.n36 VP.n35 179.006
R11 VP.n62 VP.n61 179.006
R12 VP.n34 VP.n33 179.006
R13 VP.n16 VP.n13 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n12 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n11 161.3
R18 VP.n24 VP.n23 161.3
R19 VP.n25 VP.n10 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n29 VP.n9 161.3
R22 VP.n31 VP.n30 161.3
R23 VP.n32 VP.n8 161.3
R24 VP.n60 VP.n0 161.3
R25 VP.n59 VP.n58 161.3
R26 VP.n57 VP.n1 161.3
R27 VP.n56 VP.n55 161.3
R28 VP.n53 VP.n2 161.3
R29 VP.n52 VP.n51 161.3
R30 VP.n50 VP.n3 161.3
R31 VP.n49 VP.n48 161.3
R32 VP.n47 VP.n4 161.3
R33 VP.n46 VP.n45 161.3
R34 VP.n44 VP.n5 161.3
R35 VP.n43 VP.n42 161.3
R36 VP.n40 VP.n6 161.3
R37 VP.n39 VP.n38 161.3
R38 VP.n37 VP.n7 161.3
R39 VP.n40 VP.n39 56.5617
R40 VP.n59 VP.n1 56.5617
R41 VP.n31 VP.n9 56.5617
R42 VP.n15 VP.n14 50.5334
R43 VP.n47 VP.n46 49.296
R44 VP.n52 VP.n3 49.296
R45 VP.n24 VP.n11 49.296
R46 VP.n19 VP.n18 49.296
R47 VP.n36 VP.n34 47.652
R48 VP.n46 VP.n5 31.8581
R49 VP.n53 VP.n52 31.8581
R50 VP.n25 VP.n24 31.8581
R51 VP.n18 VP.n13 31.8581
R52 VP.n39 VP.n7 24.5923
R53 VP.n42 VP.n40 24.5923
R54 VP.n48 VP.n47 24.5923
R55 VP.n48 VP.n3 24.5923
R56 VP.n55 VP.n1 24.5923
R57 VP.n60 VP.n59 24.5923
R58 VP.n32 VP.n31 24.5923
R59 VP.n27 VP.n9 24.5923
R60 VP.n20 VP.n19 24.5923
R61 VP.n20 VP.n11 24.5923
R62 VP.n16 VP.n15 18.0715
R63 VP.n41 VP.n5 15.7393
R64 VP.n54 VP.n53 15.7393
R65 VP.n26 VP.n25 15.7393
R66 VP.n14 VP.n13 15.7393
R67 VP.n42 VP.n41 8.85356
R68 VP.n55 VP.n54 8.85356
R69 VP.n27 VP.n26 8.85356
R70 VP.n35 VP.n7 6.88621
R71 VP.n61 VP.n60 6.88621
R72 VP.n33 VP.n32 6.88621
R73 VP.n17 VP.n16 0.189894
R74 VP.n17 VP.n12 0.189894
R75 VP.n21 VP.n12 0.189894
R76 VP.n22 VP.n21 0.189894
R77 VP.n23 VP.n22 0.189894
R78 VP.n23 VP.n10 0.189894
R79 VP.n28 VP.n10 0.189894
R80 VP.n29 VP.n28 0.189894
R81 VP.n30 VP.n29 0.189894
R82 VP.n30 VP.n8 0.189894
R83 VP.n34 VP.n8 0.189894
R84 VP.n37 VP.n36 0.189894
R85 VP.n38 VP.n37 0.189894
R86 VP.n38 VP.n6 0.189894
R87 VP.n43 VP.n6 0.189894
R88 VP.n44 VP.n43 0.189894
R89 VP.n45 VP.n44 0.189894
R90 VP.n45 VP.n4 0.189894
R91 VP.n49 VP.n4 0.189894
R92 VP.n50 VP.n49 0.189894
R93 VP.n51 VP.n50 0.189894
R94 VP.n51 VP.n2 0.189894
R95 VP.n56 VP.n2 0.189894
R96 VP.n57 VP.n56 0.189894
R97 VP.n58 VP.n57 0.189894
R98 VP.n58 VP.n0 0.189894
R99 VP.n62 VP.n0 0.189894
R100 VP VP.n62 0.0516364
R101 VTAIL.n11 VTAIL.t6 47.5822
R102 VTAIL.n17 VTAIL.t4 47.581
R103 VTAIL.n2 VTAIL.t9 47.581
R104 VTAIL.n16 VTAIL.t15 47.581
R105 VTAIL.n15 VTAIL.n14 46.0497
R106 VTAIL.n13 VTAIL.n12 46.0497
R107 VTAIL.n10 VTAIL.n9 46.0497
R108 VTAIL.n8 VTAIL.n7 46.0497
R109 VTAIL.n19 VTAIL.n18 46.0485
R110 VTAIL.n1 VTAIL.n0 46.0485
R111 VTAIL.n4 VTAIL.n3 46.0485
R112 VTAIL.n6 VTAIL.n5 46.0485
R113 VTAIL.n8 VTAIL.n6 26.6427
R114 VTAIL.n17 VTAIL.n16 25.0738
R115 VTAIL.n10 VTAIL.n8 1.56947
R116 VTAIL.n11 VTAIL.n10 1.56947
R117 VTAIL.n15 VTAIL.n13 1.56947
R118 VTAIL.n16 VTAIL.n15 1.56947
R119 VTAIL.n6 VTAIL.n4 1.56947
R120 VTAIL.n4 VTAIL.n2 1.56947
R121 VTAIL.n19 VTAIL.n17 1.56947
R122 VTAIL.n18 VTAIL.t7 1.53301
R123 VTAIL.n18 VTAIL.t1 1.53301
R124 VTAIL.n0 VTAIL.t3 1.53301
R125 VTAIL.n0 VTAIL.t2 1.53301
R126 VTAIL.n3 VTAIL.t12 1.53301
R127 VTAIL.n3 VTAIL.t14 1.53301
R128 VTAIL.n5 VTAIL.t18 1.53301
R129 VTAIL.n5 VTAIL.t11 1.53301
R130 VTAIL.n14 VTAIL.t17 1.53301
R131 VTAIL.n14 VTAIL.t16 1.53301
R132 VTAIL.n12 VTAIL.t10 1.53301
R133 VTAIL.n12 VTAIL.t13 1.53301
R134 VTAIL.n9 VTAIL.t0 1.53301
R135 VTAIL.n9 VTAIL.t8 1.53301
R136 VTAIL.n7 VTAIL.t19 1.53301
R137 VTAIL.n7 VTAIL.t5 1.53301
R138 VTAIL.n13 VTAIL.n11 1.25481
R139 VTAIL.n2 VTAIL.n1 1.25481
R140 VTAIL VTAIL.n1 1.23541
R141 VTAIL VTAIL.n19 0.334552
R142 VDD1.n1 VDD1.t7 65.8299
R143 VDD1.n3 VDD1.t8 65.8288
R144 VDD1.n5 VDD1.n4 63.8487
R145 VDD1.n1 VDD1.n0 62.7285
R146 VDD1.n7 VDD1.n6 62.7273
R147 VDD1.n3 VDD1.n2 62.7273
R148 VDD1.n7 VDD1.n5 43.6733
R149 VDD1.n6 VDD1.t6 1.53301
R150 VDD1.n6 VDD1.t3 1.53301
R151 VDD1.n0 VDD1.t2 1.53301
R152 VDD1.n0 VDD1.t9 1.53301
R153 VDD1.n4 VDD1.t1 1.53301
R154 VDD1.n4 VDD1.t5 1.53301
R155 VDD1.n2 VDD1.t0 1.53301
R156 VDD1.n2 VDD1.t4 1.53301
R157 VDD1 VDD1.n7 1.11903
R158 VDD1 VDD1.n1 0.450931
R159 VDD1.n5 VDD1.n3 0.337395
R160 B.n822 B.n821 585
R161 B.n321 B.n124 585
R162 B.n320 B.n319 585
R163 B.n318 B.n317 585
R164 B.n316 B.n315 585
R165 B.n314 B.n313 585
R166 B.n312 B.n311 585
R167 B.n310 B.n309 585
R168 B.n308 B.n307 585
R169 B.n306 B.n305 585
R170 B.n304 B.n303 585
R171 B.n302 B.n301 585
R172 B.n300 B.n299 585
R173 B.n298 B.n297 585
R174 B.n296 B.n295 585
R175 B.n294 B.n293 585
R176 B.n292 B.n291 585
R177 B.n290 B.n289 585
R178 B.n288 B.n287 585
R179 B.n286 B.n285 585
R180 B.n284 B.n283 585
R181 B.n282 B.n281 585
R182 B.n280 B.n279 585
R183 B.n278 B.n277 585
R184 B.n276 B.n275 585
R185 B.n274 B.n273 585
R186 B.n272 B.n271 585
R187 B.n270 B.n269 585
R188 B.n268 B.n267 585
R189 B.n266 B.n265 585
R190 B.n264 B.n263 585
R191 B.n262 B.n261 585
R192 B.n260 B.n259 585
R193 B.n258 B.n257 585
R194 B.n256 B.n255 585
R195 B.n254 B.n253 585
R196 B.n252 B.n251 585
R197 B.n250 B.n249 585
R198 B.n248 B.n247 585
R199 B.n246 B.n245 585
R200 B.n244 B.n243 585
R201 B.n242 B.n241 585
R202 B.n240 B.n239 585
R203 B.n238 B.n237 585
R204 B.n236 B.n235 585
R205 B.n234 B.n233 585
R206 B.n232 B.n231 585
R207 B.n230 B.n229 585
R208 B.n228 B.n227 585
R209 B.n226 B.n225 585
R210 B.n224 B.n223 585
R211 B.n222 B.n221 585
R212 B.n220 B.n219 585
R213 B.n218 B.n217 585
R214 B.n216 B.n215 585
R215 B.n214 B.n213 585
R216 B.n212 B.n211 585
R217 B.n210 B.n209 585
R218 B.n208 B.n207 585
R219 B.n206 B.n205 585
R220 B.n204 B.n203 585
R221 B.n202 B.n201 585
R222 B.n200 B.n199 585
R223 B.n198 B.n197 585
R224 B.n196 B.n195 585
R225 B.n194 B.n193 585
R226 B.n192 B.n191 585
R227 B.n190 B.n189 585
R228 B.n188 B.n187 585
R229 B.n186 B.n185 585
R230 B.n184 B.n183 585
R231 B.n182 B.n181 585
R232 B.n180 B.n179 585
R233 B.n178 B.n177 585
R234 B.n176 B.n175 585
R235 B.n174 B.n173 585
R236 B.n172 B.n171 585
R237 B.n170 B.n169 585
R238 B.n168 B.n167 585
R239 B.n166 B.n165 585
R240 B.n164 B.n163 585
R241 B.n162 B.n161 585
R242 B.n160 B.n159 585
R243 B.n158 B.n157 585
R244 B.n156 B.n155 585
R245 B.n154 B.n153 585
R246 B.n152 B.n151 585
R247 B.n150 B.n149 585
R248 B.n148 B.n147 585
R249 B.n146 B.n145 585
R250 B.n144 B.n143 585
R251 B.n142 B.n141 585
R252 B.n140 B.n139 585
R253 B.n138 B.n137 585
R254 B.n136 B.n135 585
R255 B.n134 B.n133 585
R256 B.n132 B.n131 585
R257 B.n74 B.n73 585
R258 B.n820 B.n75 585
R259 B.n825 B.n75 585
R260 B.n819 B.n818 585
R261 B.n818 B.n71 585
R262 B.n817 B.n70 585
R263 B.n831 B.n70 585
R264 B.n816 B.n69 585
R265 B.n832 B.n69 585
R266 B.n815 B.n68 585
R267 B.n833 B.n68 585
R268 B.n814 B.n813 585
R269 B.n813 B.n67 585
R270 B.n812 B.n63 585
R271 B.n839 B.n63 585
R272 B.n811 B.n62 585
R273 B.n840 B.n62 585
R274 B.n810 B.n61 585
R275 B.n841 B.n61 585
R276 B.n809 B.n808 585
R277 B.n808 B.n57 585
R278 B.n807 B.n56 585
R279 B.n847 B.n56 585
R280 B.n806 B.n55 585
R281 B.n848 B.n55 585
R282 B.n805 B.n54 585
R283 B.n849 B.n54 585
R284 B.n804 B.n803 585
R285 B.n803 B.n50 585
R286 B.n802 B.n49 585
R287 B.n855 B.n49 585
R288 B.n801 B.n48 585
R289 B.n856 B.n48 585
R290 B.n800 B.n47 585
R291 B.n857 B.n47 585
R292 B.n799 B.n798 585
R293 B.n798 B.n43 585
R294 B.n797 B.n42 585
R295 B.n863 B.n42 585
R296 B.n796 B.n41 585
R297 B.n864 B.n41 585
R298 B.n795 B.n40 585
R299 B.n865 B.n40 585
R300 B.n794 B.n793 585
R301 B.n793 B.n36 585
R302 B.n792 B.n35 585
R303 B.n871 B.n35 585
R304 B.n791 B.n34 585
R305 B.n872 B.n34 585
R306 B.n790 B.n33 585
R307 B.n873 B.n33 585
R308 B.n789 B.n788 585
R309 B.n788 B.n32 585
R310 B.n787 B.n28 585
R311 B.n879 B.n28 585
R312 B.n786 B.n27 585
R313 B.n880 B.n27 585
R314 B.n785 B.n26 585
R315 B.n881 B.n26 585
R316 B.n784 B.n783 585
R317 B.n783 B.n22 585
R318 B.n782 B.n21 585
R319 B.n887 B.n21 585
R320 B.n781 B.n20 585
R321 B.n888 B.n20 585
R322 B.n780 B.n19 585
R323 B.n889 B.n19 585
R324 B.n779 B.n778 585
R325 B.n778 B.n15 585
R326 B.n777 B.n14 585
R327 B.n895 B.n14 585
R328 B.n776 B.n13 585
R329 B.n896 B.n13 585
R330 B.n775 B.n12 585
R331 B.n897 B.n12 585
R332 B.n774 B.n773 585
R333 B.n773 B.n8 585
R334 B.n772 B.n7 585
R335 B.n903 B.n7 585
R336 B.n771 B.n6 585
R337 B.n904 B.n6 585
R338 B.n770 B.n5 585
R339 B.n905 B.n5 585
R340 B.n769 B.n768 585
R341 B.n768 B.n4 585
R342 B.n767 B.n322 585
R343 B.n767 B.n766 585
R344 B.n757 B.n323 585
R345 B.n324 B.n323 585
R346 B.n759 B.n758 585
R347 B.n760 B.n759 585
R348 B.n756 B.n328 585
R349 B.n332 B.n328 585
R350 B.n755 B.n754 585
R351 B.n754 B.n753 585
R352 B.n330 B.n329 585
R353 B.n331 B.n330 585
R354 B.n746 B.n745 585
R355 B.n747 B.n746 585
R356 B.n744 B.n337 585
R357 B.n337 B.n336 585
R358 B.n743 B.n742 585
R359 B.n742 B.n741 585
R360 B.n339 B.n338 585
R361 B.n340 B.n339 585
R362 B.n734 B.n733 585
R363 B.n735 B.n734 585
R364 B.n732 B.n345 585
R365 B.n345 B.n344 585
R366 B.n731 B.n730 585
R367 B.n730 B.n729 585
R368 B.n347 B.n346 585
R369 B.n722 B.n347 585
R370 B.n721 B.n720 585
R371 B.n723 B.n721 585
R372 B.n719 B.n352 585
R373 B.n352 B.n351 585
R374 B.n718 B.n717 585
R375 B.n717 B.n716 585
R376 B.n354 B.n353 585
R377 B.n355 B.n354 585
R378 B.n709 B.n708 585
R379 B.n710 B.n709 585
R380 B.n707 B.n359 585
R381 B.n363 B.n359 585
R382 B.n706 B.n705 585
R383 B.n705 B.n704 585
R384 B.n361 B.n360 585
R385 B.n362 B.n361 585
R386 B.n697 B.n696 585
R387 B.n698 B.n697 585
R388 B.n695 B.n368 585
R389 B.n368 B.n367 585
R390 B.n694 B.n693 585
R391 B.n693 B.n692 585
R392 B.n370 B.n369 585
R393 B.n371 B.n370 585
R394 B.n685 B.n684 585
R395 B.n686 B.n685 585
R396 B.n683 B.n376 585
R397 B.n376 B.n375 585
R398 B.n682 B.n681 585
R399 B.n681 B.n680 585
R400 B.n378 B.n377 585
R401 B.n379 B.n378 585
R402 B.n673 B.n672 585
R403 B.n674 B.n673 585
R404 B.n671 B.n384 585
R405 B.n384 B.n383 585
R406 B.n670 B.n669 585
R407 B.n669 B.n668 585
R408 B.n386 B.n385 585
R409 B.n661 B.n386 585
R410 B.n660 B.n659 585
R411 B.n662 B.n660 585
R412 B.n658 B.n391 585
R413 B.n391 B.n390 585
R414 B.n657 B.n656 585
R415 B.n656 B.n655 585
R416 B.n393 B.n392 585
R417 B.n394 B.n393 585
R418 B.n648 B.n647 585
R419 B.n649 B.n648 585
R420 B.n397 B.n396 585
R421 B.n452 B.n450 585
R422 B.n453 B.n449 585
R423 B.n453 B.n398 585
R424 B.n456 B.n455 585
R425 B.n457 B.n448 585
R426 B.n459 B.n458 585
R427 B.n461 B.n447 585
R428 B.n464 B.n463 585
R429 B.n465 B.n446 585
R430 B.n467 B.n466 585
R431 B.n469 B.n445 585
R432 B.n472 B.n471 585
R433 B.n473 B.n444 585
R434 B.n475 B.n474 585
R435 B.n477 B.n443 585
R436 B.n480 B.n479 585
R437 B.n481 B.n442 585
R438 B.n483 B.n482 585
R439 B.n485 B.n441 585
R440 B.n488 B.n487 585
R441 B.n489 B.n440 585
R442 B.n491 B.n490 585
R443 B.n493 B.n439 585
R444 B.n496 B.n495 585
R445 B.n497 B.n438 585
R446 B.n499 B.n498 585
R447 B.n501 B.n437 585
R448 B.n504 B.n503 585
R449 B.n505 B.n436 585
R450 B.n507 B.n506 585
R451 B.n509 B.n435 585
R452 B.n512 B.n511 585
R453 B.n513 B.n434 585
R454 B.n515 B.n514 585
R455 B.n517 B.n433 585
R456 B.n520 B.n519 585
R457 B.n521 B.n432 585
R458 B.n523 B.n522 585
R459 B.n525 B.n431 585
R460 B.n528 B.n527 585
R461 B.n529 B.n430 585
R462 B.n531 B.n530 585
R463 B.n533 B.n429 585
R464 B.n536 B.n535 585
R465 B.n538 B.n426 585
R466 B.n540 B.n539 585
R467 B.n542 B.n425 585
R468 B.n545 B.n544 585
R469 B.n546 B.n424 585
R470 B.n548 B.n547 585
R471 B.n550 B.n423 585
R472 B.n553 B.n552 585
R473 B.n554 B.n422 585
R474 B.n559 B.n558 585
R475 B.n561 B.n421 585
R476 B.n564 B.n563 585
R477 B.n565 B.n420 585
R478 B.n567 B.n566 585
R479 B.n569 B.n419 585
R480 B.n572 B.n571 585
R481 B.n573 B.n418 585
R482 B.n575 B.n574 585
R483 B.n577 B.n417 585
R484 B.n580 B.n579 585
R485 B.n581 B.n416 585
R486 B.n583 B.n582 585
R487 B.n585 B.n415 585
R488 B.n588 B.n587 585
R489 B.n589 B.n414 585
R490 B.n591 B.n590 585
R491 B.n593 B.n413 585
R492 B.n596 B.n595 585
R493 B.n597 B.n412 585
R494 B.n599 B.n598 585
R495 B.n601 B.n411 585
R496 B.n604 B.n603 585
R497 B.n605 B.n410 585
R498 B.n607 B.n606 585
R499 B.n609 B.n409 585
R500 B.n612 B.n611 585
R501 B.n613 B.n408 585
R502 B.n615 B.n614 585
R503 B.n617 B.n407 585
R504 B.n620 B.n619 585
R505 B.n621 B.n406 585
R506 B.n623 B.n622 585
R507 B.n625 B.n405 585
R508 B.n628 B.n627 585
R509 B.n629 B.n404 585
R510 B.n631 B.n630 585
R511 B.n633 B.n403 585
R512 B.n636 B.n635 585
R513 B.n637 B.n402 585
R514 B.n639 B.n638 585
R515 B.n641 B.n401 585
R516 B.n642 B.n400 585
R517 B.n645 B.n644 585
R518 B.n646 B.n399 585
R519 B.n399 B.n398 585
R520 B.n651 B.n650 585
R521 B.n650 B.n649 585
R522 B.n652 B.n395 585
R523 B.n395 B.n394 585
R524 B.n654 B.n653 585
R525 B.n655 B.n654 585
R526 B.n389 B.n388 585
R527 B.n390 B.n389 585
R528 B.n664 B.n663 585
R529 B.n663 B.n662 585
R530 B.n665 B.n387 585
R531 B.n661 B.n387 585
R532 B.n667 B.n666 585
R533 B.n668 B.n667 585
R534 B.n382 B.n381 585
R535 B.n383 B.n382 585
R536 B.n676 B.n675 585
R537 B.n675 B.n674 585
R538 B.n677 B.n380 585
R539 B.n380 B.n379 585
R540 B.n679 B.n678 585
R541 B.n680 B.n679 585
R542 B.n374 B.n373 585
R543 B.n375 B.n374 585
R544 B.n688 B.n687 585
R545 B.n687 B.n686 585
R546 B.n689 B.n372 585
R547 B.n372 B.n371 585
R548 B.n691 B.n690 585
R549 B.n692 B.n691 585
R550 B.n366 B.n365 585
R551 B.n367 B.n366 585
R552 B.n700 B.n699 585
R553 B.n699 B.n698 585
R554 B.n701 B.n364 585
R555 B.n364 B.n362 585
R556 B.n703 B.n702 585
R557 B.n704 B.n703 585
R558 B.n358 B.n357 585
R559 B.n363 B.n358 585
R560 B.n712 B.n711 585
R561 B.n711 B.n710 585
R562 B.n713 B.n356 585
R563 B.n356 B.n355 585
R564 B.n715 B.n714 585
R565 B.n716 B.n715 585
R566 B.n350 B.n349 585
R567 B.n351 B.n350 585
R568 B.n725 B.n724 585
R569 B.n724 B.n723 585
R570 B.n726 B.n348 585
R571 B.n722 B.n348 585
R572 B.n728 B.n727 585
R573 B.n729 B.n728 585
R574 B.n343 B.n342 585
R575 B.n344 B.n343 585
R576 B.n737 B.n736 585
R577 B.n736 B.n735 585
R578 B.n738 B.n341 585
R579 B.n341 B.n340 585
R580 B.n740 B.n739 585
R581 B.n741 B.n740 585
R582 B.n335 B.n334 585
R583 B.n336 B.n335 585
R584 B.n749 B.n748 585
R585 B.n748 B.n747 585
R586 B.n750 B.n333 585
R587 B.n333 B.n331 585
R588 B.n752 B.n751 585
R589 B.n753 B.n752 585
R590 B.n327 B.n326 585
R591 B.n332 B.n327 585
R592 B.n762 B.n761 585
R593 B.n761 B.n760 585
R594 B.n763 B.n325 585
R595 B.n325 B.n324 585
R596 B.n765 B.n764 585
R597 B.n766 B.n765 585
R598 B.n2 B.n0 585
R599 B.n4 B.n2 585
R600 B.n3 B.n1 585
R601 B.n904 B.n3 585
R602 B.n902 B.n901 585
R603 B.n903 B.n902 585
R604 B.n900 B.n9 585
R605 B.n9 B.n8 585
R606 B.n899 B.n898 585
R607 B.n898 B.n897 585
R608 B.n11 B.n10 585
R609 B.n896 B.n11 585
R610 B.n894 B.n893 585
R611 B.n895 B.n894 585
R612 B.n892 B.n16 585
R613 B.n16 B.n15 585
R614 B.n891 B.n890 585
R615 B.n890 B.n889 585
R616 B.n18 B.n17 585
R617 B.n888 B.n18 585
R618 B.n886 B.n885 585
R619 B.n887 B.n886 585
R620 B.n884 B.n23 585
R621 B.n23 B.n22 585
R622 B.n883 B.n882 585
R623 B.n882 B.n881 585
R624 B.n25 B.n24 585
R625 B.n880 B.n25 585
R626 B.n878 B.n877 585
R627 B.n879 B.n878 585
R628 B.n876 B.n29 585
R629 B.n32 B.n29 585
R630 B.n875 B.n874 585
R631 B.n874 B.n873 585
R632 B.n31 B.n30 585
R633 B.n872 B.n31 585
R634 B.n870 B.n869 585
R635 B.n871 B.n870 585
R636 B.n868 B.n37 585
R637 B.n37 B.n36 585
R638 B.n867 B.n866 585
R639 B.n866 B.n865 585
R640 B.n39 B.n38 585
R641 B.n864 B.n39 585
R642 B.n862 B.n861 585
R643 B.n863 B.n862 585
R644 B.n860 B.n44 585
R645 B.n44 B.n43 585
R646 B.n859 B.n858 585
R647 B.n858 B.n857 585
R648 B.n46 B.n45 585
R649 B.n856 B.n46 585
R650 B.n854 B.n853 585
R651 B.n855 B.n854 585
R652 B.n852 B.n51 585
R653 B.n51 B.n50 585
R654 B.n851 B.n850 585
R655 B.n850 B.n849 585
R656 B.n53 B.n52 585
R657 B.n848 B.n53 585
R658 B.n846 B.n845 585
R659 B.n847 B.n846 585
R660 B.n844 B.n58 585
R661 B.n58 B.n57 585
R662 B.n843 B.n842 585
R663 B.n842 B.n841 585
R664 B.n60 B.n59 585
R665 B.n840 B.n60 585
R666 B.n838 B.n837 585
R667 B.n839 B.n838 585
R668 B.n836 B.n64 585
R669 B.n67 B.n64 585
R670 B.n835 B.n834 585
R671 B.n834 B.n833 585
R672 B.n66 B.n65 585
R673 B.n832 B.n66 585
R674 B.n830 B.n829 585
R675 B.n831 B.n830 585
R676 B.n828 B.n72 585
R677 B.n72 B.n71 585
R678 B.n827 B.n826 585
R679 B.n826 B.n825 585
R680 B.n907 B.n906 585
R681 B.n906 B.n905 585
R682 B.n650 B.n397 554.963
R683 B.n826 B.n74 554.963
R684 B.n648 B.n399 554.963
R685 B.n822 B.n75 554.963
R686 B.n555 B.t20 414.377
R687 B.n427 B.t13 414.377
R688 B.n128 B.t9 414.377
R689 B.n125 B.t17 414.377
R690 B.n824 B.n823 256.663
R691 B.n824 B.n123 256.663
R692 B.n824 B.n122 256.663
R693 B.n824 B.n121 256.663
R694 B.n824 B.n120 256.663
R695 B.n824 B.n119 256.663
R696 B.n824 B.n118 256.663
R697 B.n824 B.n117 256.663
R698 B.n824 B.n116 256.663
R699 B.n824 B.n115 256.663
R700 B.n824 B.n114 256.663
R701 B.n824 B.n113 256.663
R702 B.n824 B.n112 256.663
R703 B.n824 B.n111 256.663
R704 B.n824 B.n110 256.663
R705 B.n824 B.n109 256.663
R706 B.n824 B.n108 256.663
R707 B.n824 B.n107 256.663
R708 B.n824 B.n106 256.663
R709 B.n824 B.n105 256.663
R710 B.n824 B.n104 256.663
R711 B.n824 B.n103 256.663
R712 B.n824 B.n102 256.663
R713 B.n824 B.n101 256.663
R714 B.n824 B.n100 256.663
R715 B.n824 B.n99 256.663
R716 B.n824 B.n98 256.663
R717 B.n824 B.n97 256.663
R718 B.n824 B.n96 256.663
R719 B.n824 B.n95 256.663
R720 B.n824 B.n94 256.663
R721 B.n824 B.n93 256.663
R722 B.n824 B.n92 256.663
R723 B.n824 B.n91 256.663
R724 B.n824 B.n90 256.663
R725 B.n824 B.n89 256.663
R726 B.n824 B.n88 256.663
R727 B.n824 B.n87 256.663
R728 B.n824 B.n86 256.663
R729 B.n824 B.n85 256.663
R730 B.n824 B.n84 256.663
R731 B.n824 B.n83 256.663
R732 B.n824 B.n82 256.663
R733 B.n824 B.n81 256.663
R734 B.n824 B.n80 256.663
R735 B.n824 B.n79 256.663
R736 B.n824 B.n78 256.663
R737 B.n824 B.n77 256.663
R738 B.n824 B.n76 256.663
R739 B.n451 B.n398 256.663
R740 B.n454 B.n398 256.663
R741 B.n460 B.n398 256.663
R742 B.n462 B.n398 256.663
R743 B.n468 B.n398 256.663
R744 B.n470 B.n398 256.663
R745 B.n476 B.n398 256.663
R746 B.n478 B.n398 256.663
R747 B.n484 B.n398 256.663
R748 B.n486 B.n398 256.663
R749 B.n492 B.n398 256.663
R750 B.n494 B.n398 256.663
R751 B.n500 B.n398 256.663
R752 B.n502 B.n398 256.663
R753 B.n508 B.n398 256.663
R754 B.n510 B.n398 256.663
R755 B.n516 B.n398 256.663
R756 B.n518 B.n398 256.663
R757 B.n524 B.n398 256.663
R758 B.n526 B.n398 256.663
R759 B.n532 B.n398 256.663
R760 B.n534 B.n398 256.663
R761 B.n541 B.n398 256.663
R762 B.n543 B.n398 256.663
R763 B.n549 B.n398 256.663
R764 B.n551 B.n398 256.663
R765 B.n560 B.n398 256.663
R766 B.n562 B.n398 256.663
R767 B.n568 B.n398 256.663
R768 B.n570 B.n398 256.663
R769 B.n576 B.n398 256.663
R770 B.n578 B.n398 256.663
R771 B.n584 B.n398 256.663
R772 B.n586 B.n398 256.663
R773 B.n592 B.n398 256.663
R774 B.n594 B.n398 256.663
R775 B.n600 B.n398 256.663
R776 B.n602 B.n398 256.663
R777 B.n608 B.n398 256.663
R778 B.n610 B.n398 256.663
R779 B.n616 B.n398 256.663
R780 B.n618 B.n398 256.663
R781 B.n624 B.n398 256.663
R782 B.n626 B.n398 256.663
R783 B.n632 B.n398 256.663
R784 B.n634 B.n398 256.663
R785 B.n640 B.n398 256.663
R786 B.n643 B.n398 256.663
R787 B.n650 B.n395 163.367
R788 B.n654 B.n395 163.367
R789 B.n654 B.n389 163.367
R790 B.n663 B.n389 163.367
R791 B.n663 B.n387 163.367
R792 B.n667 B.n387 163.367
R793 B.n667 B.n382 163.367
R794 B.n675 B.n382 163.367
R795 B.n675 B.n380 163.367
R796 B.n679 B.n380 163.367
R797 B.n679 B.n374 163.367
R798 B.n687 B.n374 163.367
R799 B.n687 B.n372 163.367
R800 B.n691 B.n372 163.367
R801 B.n691 B.n366 163.367
R802 B.n699 B.n366 163.367
R803 B.n699 B.n364 163.367
R804 B.n703 B.n364 163.367
R805 B.n703 B.n358 163.367
R806 B.n711 B.n358 163.367
R807 B.n711 B.n356 163.367
R808 B.n715 B.n356 163.367
R809 B.n715 B.n350 163.367
R810 B.n724 B.n350 163.367
R811 B.n724 B.n348 163.367
R812 B.n728 B.n348 163.367
R813 B.n728 B.n343 163.367
R814 B.n736 B.n343 163.367
R815 B.n736 B.n341 163.367
R816 B.n740 B.n341 163.367
R817 B.n740 B.n335 163.367
R818 B.n748 B.n335 163.367
R819 B.n748 B.n333 163.367
R820 B.n752 B.n333 163.367
R821 B.n752 B.n327 163.367
R822 B.n761 B.n327 163.367
R823 B.n761 B.n325 163.367
R824 B.n765 B.n325 163.367
R825 B.n765 B.n2 163.367
R826 B.n906 B.n2 163.367
R827 B.n906 B.n3 163.367
R828 B.n902 B.n3 163.367
R829 B.n902 B.n9 163.367
R830 B.n898 B.n9 163.367
R831 B.n898 B.n11 163.367
R832 B.n894 B.n11 163.367
R833 B.n894 B.n16 163.367
R834 B.n890 B.n16 163.367
R835 B.n890 B.n18 163.367
R836 B.n886 B.n18 163.367
R837 B.n886 B.n23 163.367
R838 B.n882 B.n23 163.367
R839 B.n882 B.n25 163.367
R840 B.n878 B.n25 163.367
R841 B.n878 B.n29 163.367
R842 B.n874 B.n29 163.367
R843 B.n874 B.n31 163.367
R844 B.n870 B.n31 163.367
R845 B.n870 B.n37 163.367
R846 B.n866 B.n37 163.367
R847 B.n866 B.n39 163.367
R848 B.n862 B.n39 163.367
R849 B.n862 B.n44 163.367
R850 B.n858 B.n44 163.367
R851 B.n858 B.n46 163.367
R852 B.n854 B.n46 163.367
R853 B.n854 B.n51 163.367
R854 B.n850 B.n51 163.367
R855 B.n850 B.n53 163.367
R856 B.n846 B.n53 163.367
R857 B.n846 B.n58 163.367
R858 B.n842 B.n58 163.367
R859 B.n842 B.n60 163.367
R860 B.n838 B.n60 163.367
R861 B.n838 B.n64 163.367
R862 B.n834 B.n64 163.367
R863 B.n834 B.n66 163.367
R864 B.n830 B.n66 163.367
R865 B.n830 B.n72 163.367
R866 B.n826 B.n72 163.367
R867 B.n453 B.n452 163.367
R868 B.n455 B.n453 163.367
R869 B.n459 B.n448 163.367
R870 B.n463 B.n461 163.367
R871 B.n467 B.n446 163.367
R872 B.n471 B.n469 163.367
R873 B.n475 B.n444 163.367
R874 B.n479 B.n477 163.367
R875 B.n483 B.n442 163.367
R876 B.n487 B.n485 163.367
R877 B.n491 B.n440 163.367
R878 B.n495 B.n493 163.367
R879 B.n499 B.n438 163.367
R880 B.n503 B.n501 163.367
R881 B.n507 B.n436 163.367
R882 B.n511 B.n509 163.367
R883 B.n515 B.n434 163.367
R884 B.n519 B.n517 163.367
R885 B.n523 B.n432 163.367
R886 B.n527 B.n525 163.367
R887 B.n531 B.n430 163.367
R888 B.n535 B.n533 163.367
R889 B.n540 B.n426 163.367
R890 B.n544 B.n542 163.367
R891 B.n548 B.n424 163.367
R892 B.n552 B.n550 163.367
R893 B.n559 B.n422 163.367
R894 B.n563 B.n561 163.367
R895 B.n567 B.n420 163.367
R896 B.n571 B.n569 163.367
R897 B.n575 B.n418 163.367
R898 B.n579 B.n577 163.367
R899 B.n583 B.n416 163.367
R900 B.n587 B.n585 163.367
R901 B.n591 B.n414 163.367
R902 B.n595 B.n593 163.367
R903 B.n599 B.n412 163.367
R904 B.n603 B.n601 163.367
R905 B.n607 B.n410 163.367
R906 B.n611 B.n609 163.367
R907 B.n615 B.n408 163.367
R908 B.n619 B.n617 163.367
R909 B.n623 B.n406 163.367
R910 B.n627 B.n625 163.367
R911 B.n631 B.n404 163.367
R912 B.n635 B.n633 163.367
R913 B.n639 B.n402 163.367
R914 B.n642 B.n641 163.367
R915 B.n644 B.n399 163.367
R916 B.n648 B.n393 163.367
R917 B.n656 B.n393 163.367
R918 B.n656 B.n391 163.367
R919 B.n660 B.n391 163.367
R920 B.n660 B.n386 163.367
R921 B.n669 B.n386 163.367
R922 B.n669 B.n384 163.367
R923 B.n673 B.n384 163.367
R924 B.n673 B.n378 163.367
R925 B.n681 B.n378 163.367
R926 B.n681 B.n376 163.367
R927 B.n685 B.n376 163.367
R928 B.n685 B.n370 163.367
R929 B.n693 B.n370 163.367
R930 B.n693 B.n368 163.367
R931 B.n697 B.n368 163.367
R932 B.n697 B.n361 163.367
R933 B.n705 B.n361 163.367
R934 B.n705 B.n359 163.367
R935 B.n709 B.n359 163.367
R936 B.n709 B.n354 163.367
R937 B.n717 B.n354 163.367
R938 B.n717 B.n352 163.367
R939 B.n721 B.n352 163.367
R940 B.n721 B.n347 163.367
R941 B.n730 B.n347 163.367
R942 B.n730 B.n345 163.367
R943 B.n734 B.n345 163.367
R944 B.n734 B.n339 163.367
R945 B.n742 B.n339 163.367
R946 B.n742 B.n337 163.367
R947 B.n746 B.n337 163.367
R948 B.n746 B.n330 163.367
R949 B.n754 B.n330 163.367
R950 B.n754 B.n328 163.367
R951 B.n759 B.n328 163.367
R952 B.n759 B.n323 163.367
R953 B.n767 B.n323 163.367
R954 B.n768 B.n767 163.367
R955 B.n768 B.n5 163.367
R956 B.n6 B.n5 163.367
R957 B.n7 B.n6 163.367
R958 B.n773 B.n7 163.367
R959 B.n773 B.n12 163.367
R960 B.n13 B.n12 163.367
R961 B.n14 B.n13 163.367
R962 B.n778 B.n14 163.367
R963 B.n778 B.n19 163.367
R964 B.n20 B.n19 163.367
R965 B.n21 B.n20 163.367
R966 B.n783 B.n21 163.367
R967 B.n783 B.n26 163.367
R968 B.n27 B.n26 163.367
R969 B.n28 B.n27 163.367
R970 B.n788 B.n28 163.367
R971 B.n788 B.n33 163.367
R972 B.n34 B.n33 163.367
R973 B.n35 B.n34 163.367
R974 B.n793 B.n35 163.367
R975 B.n793 B.n40 163.367
R976 B.n41 B.n40 163.367
R977 B.n42 B.n41 163.367
R978 B.n798 B.n42 163.367
R979 B.n798 B.n47 163.367
R980 B.n48 B.n47 163.367
R981 B.n49 B.n48 163.367
R982 B.n803 B.n49 163.367
R983 B.n803 B.n54 163.367
R984 B.n55 B.n54 163.367
R985 B.n56 B.n55 163.367
R986 B.n808 B.n56 163.367
R987 B.n808 B.n61 163.367
R988 B.n62 B.n61 163.367
R989 B.n63 B.n62 163.367
R990 B.n813 B.n63 163.367
R991 B.n813 B.n68 163.367
R992 B.n69 B.n68 163.367
R993 B.n70 B.n69 163.367
R994 B.n818 B.n70 163.367
R995 B.n818 B.n75 163.367
R996 B.n133 B.n132 163.367
R997 B.n137 B.n136 163.367
R998 B.n141 B.n140 163.367
R999 B.n145 B.n144 163.367
R1000 B.n149 B.n148 163.367
R1001 B.n153 B.n152 163.367
R1002 B.n157 B.n156 163.367
R1003 B.n161 B.n160 163.367
R1004 B.n165 B.n164 163.367
R1005 B.n169 B.n168 163.367
R1006 B.n173 B.n172 163.367
R1007 B.n177 B.n176 163.367
R1008 B.n181 B.n180 163.367
R1009 B.n185 B.n184 163.367
R1010 B.n189 B.n188 163.367
R1011 B.n193 B.n192 163.367
R1012 B.n197 B.n196 163.367
R1013 B.n201 B.n200 163.367
R1014 B.n205 B.n204 163.367
R1015 B.n209 B.n208 163.367
R1016 B.n213 B.n212 163.367
R1017 B.n217 B.n216 163.367
R1018 B.n221 B.n220 163.367
R1019 B.n225 B.n224 163.367
R1020 B.n229 B.n228 163.367
R1021 B.n233 B.n232 163.367
R1022 B.n237 B.n236 163.367
R1023 B.n241 B.n240 163.367
R1024 B.n245 B.n244 163.367
R1025 B.n249 B.n248 163.367
R1026 B.n253 B.n252 163.367
R1027 B.n257 B.n256 163.367
R1028 B.n261 B.n260 163.367
R1029 B.n265 B.n264 163.367
R1030 B.n269 B.n268 163.367
R1031 B.n273 B.n272 163.367
R1032 B.n277 B.n276 163.367
R1033 B.n281 B.n280 163.367
R1034 B.n285 B.n284 163.367
R1035 B.n289 B.n288 163.367
R1036 B.n293 B.n292 163.367
R1037 B.n297 B.n296 163.367
R1038 B.n301 B.n300 163.367
R1039 B.n305 B.n304 163.367
R1040 B.n309 B.n308 163.367
R1041 B.n313 B.n312 163.367
R1042 B.n317 B.n316 163.367
R1043 B.n319 B.n124 163.367
R1044 B.n555 B.t22 102.971
R1045 B.n125 B.t18 102.971
R1046 B.n427 B.t16 102.954
R1047 B.n128 B.t11 102.954
R1048 B.n649 B.n398 84.0346
R1049 B.n825 B.n824 84.0346
R1050 B.n451 B.n397 71.676
R1051 B.n455 B.n454 71.676
R1052 B.n460 B.n459 71.676
R1053 B.n463 B.n462 71.676
R1054 B.n468 B.n467 71.676
R1055 B.n471 B.n470 71.676
R1056 B.n476 B.n475 71.676
R1057 B.n479 B.n478 71.676
R1058 B.n484 B.n483 71.676
R1059 B.n487 B.n486 71.676
R1060 B.n492 B.n491 71.676
R1061 B.n495 B.n494 71.676
R1062 B.n500 B.n499 71.676
R1063 B.n503 B.n502 71.676
R1064 B.n508 B.n507 71.676
R1065 B.n511 B.n510 71.676
R1066 B.n516 B.n515 71.676
R1067 B.n519 B.n518 71.676
R1068 B.n524 B.n523 71.676
R1069 B.n527 B.n526 71.676
R1070 B.n532 B.n531 71.676
R1071 B.n535 B.n534 71.676
R1072 B.n541 B.n540 71.676
R1073 B.n544 B.n543 71.676
R1074 B.n549 B.n548 71.676
R1075 B.n552 B.n551 71.676
R1076 B.n560 B.n559 71.676
R1077 B.n563 B.n562 71.676
R1078 B.n568 B.n567 71.676
R1079 B.n571 B.n570 71.676
R1080 B.n576 B.n575 71.676
R1081 B.n579 B.n578 71.676
R1082 B.n584 B.n583 71.676
R1083 B.n587 B.n586 71.676
R1084 B.n592 B.n591 71.676
R1085 B.n595 B.n594 71.676
R1086 B.n600 B.n599 71.676
R1087 B.n603 B.n602 71.676
R1088 B.n608 B.n607 71.676
R1089 B.n611 B.n610 71.676
R1090 B.n616 B.n615 71.676
R1091 B.n619 B.n618 71.676
R1092 B.n624 B.n623 71.676
R1093 B.n627 B.n626 71.676
R1094 B.n632 B.n631 71.676
R1095 B.n635 B.n634 71.676
R1096 B.n640 B.n639 71.676
R1097 B.n643 B.n642 71.676
R1098 B.n76 B.n74 71.676
R1099 B.n133 B.n77 71.676
R1100 B.n137 B.n78 71.676
R1101 B.n141 B.n79 71.676
R1102 B.n145 B.n80 71.676
R1103 B.n149 B.n81 71.676
R1104 B.n153 B.n82 71.676
R1105 B.n157 B.n83 71.676
R1106 B.n161 B.n84 71.676
R1107 B.n165 B.n85 71.676
R1108 B.n169 B.n86 71.676
R1109 B.n173 B.n87 71.676
R1110 B.n177 B.n88 71.676
R1111 B.n181 B.n89 71.676
R1112 B.n185 B.n90 71.676
R1113 B.n189 B.n91 71.676
R1114 B.n193 B.n92 71.676
R1115 B.n197 B.n93 71.676
R1116 B.n201 B.n94 71.676
R1117 B.n205 B.n95 71.676
R1118 B.n209 B.n96 71.676
R1119 B.n213 B.n97 71.676
R1120 B.n217 B.n98 71.676
R1121 B.n221 B.n99 71.676
R1122 B.n225 B.n100 71.676
R1123 B.n229 B.n101 71.676
R1124 B.n233 B.n102 71.676
R1125 B.n237 B.n103 71.676
R1126 B.n241 B.n104 71.676
R1127 B.n245 B.n105 71.676
R1128 B.n249 B.n106 71.676
R1129 B.n253 B.n107 71.676
R1130 B.n257 B.n108 71.676
R1131 B.n261 B.n109 71.676
R1132 B.n265 B.n110 71.676
R1133 B.n269 B.n111 71.676
R1134 B.n273 B.n112 71.676
R1135 B.n277 B.n113 71.676
R1136 B.n281 B.n114 71.676
R1137 B.n285 B.n115 71.676
R1138 B.n289 B.n116 71.676
R1139 B.n293 B.n117 71.676
R1140 B.n297 B.n118 71.676
R1141 B.n301 B.n119 71.676
R1142 B.n305 B.n120 71.676
R1143 B.n309 B.n121 71.676
R1144 B.n313 B.n122 71.676
R1145 B.n317 B.n123 71.676
R1146 B.n823 B.n124 71.676
R1147 B.n823 B.n822 71.676
R1148 B.n319 B.n123 71.676
R1149 B.n316 B.n122 71.676
R1150 B.n312 B.n121 71.676
R1151 B.n308 B.n120 71.676
R1152 B.n304 B.n119 71.676
R1153 B.n300 B.n118 71.676
R1154 B.n296 B.n117 71.676
R1155 B.n292 B.n116 71.676
R1156 B.n288 B.n115 71.676
R1157 B.n284 B.n114 71.676
R1158 B.n280 B.n113 71.676
R1159 B.n276 B.n112 71.676
R1160 B.n272 B.n111 71.676
R1161 B.n268 B.n110 71.676
R1162 B.n264 B.n109 71.676
R1163 B.n260 B.n108 71.676
R1164 B.n256 B.n107 71.676
R1165 B.n252 B.n106 71.676
R1166 B.n248 B.n105 71.676
R1167 B.n244 B.n104 71.676
R1168 B.n240 B.n103 71.676
R1169 B.n236 B.n102 71.676
R1170 B.n232 B.n101 71.676
R1171 B.n228 B.n100 71.676
R1172 B.n224 B.n99 71.676
R1173 B.n220 B.n98 71.676
R1174 B.n216 B.n97 71.676
R1175 B.n212 B.n96 71.676
R1176 B.n208 B.n95 71.676
R1177 B.n204 B.n94 71.676
R1178 B.n200 B.n93 71.676
R1179 B.n196 B.n92 71.676
R1180 B.n192 B.n91 71.676
R1181 B.n188 B.n90 71.676
R1182 B.n184 B.n89 71.676
R1183 B.n180 B.n88 71.676
R1184 B.n176 B.n87 71.676
R1185 B.n172 B.n86 71.676
R1186 B.n168 B.n85 71.676
R1187 B.n164 B.n84 71.676
R1188 B.n160 B.n83 71.676
R1189 B.n156 B.n82 71.676
R1190 B.n152 B.n81 71.676
R1191 B.n148 B.n80 71.676
R1192 B.n144 B.n79 71.676
R1193 B.n140 B.n78 71.676
R1194 B.n136 B.n77 71.676
R1195 B.n132 B.n76 71.676
R1196 B.n452 B.n451 71.676
R1197 B.n454 B.n448 71.676
R1198 B.n461 B.n460 71.676
R1199 B.n462 B.n446 71.676
R1200 B.n469 B.n468 71.676
R1201 B.n470 B.n444 71.676
R1202 B.n477 B.n476 71.676
R1203 B.n478 B.n442 71.676
R1204 B.n485 B.n484 71.676
R1205 B.n486 B.n440 71.676
R1206 B.n493 B.n492 71.676
R1207 B.n494 B.n438 71.676
R1208 B.n501 B.n500 71.676
R1209 B.n502 B.n436 71.676
R1210 B.n509 B.n508 71.676
R1211 B.n510 B.n434 71.676
R1212 B.n517 B.n516 71.676
R1213 B.n518 B.n432 71.676
R1214 B.n525 B.n524 71.676
R1215 B.n526 B.n430 71.676
R1216 B.n533 B.n532 71.676
R1217 B.n534 B.n426 71.676
R1218 B.n542 B.n541 71.676
R1219 B.n543 B.n424 71.676
R1220 B.n550 B.n549 71.676
R1221 B.n551 B.n422 71.676
R1222 B.n561 B.n560 71.676
R1223 B.n562 B.n420 71.676
R1224 B.n569 B.n568 71.676
R1225 B.n570 B.n418 71.676
R1226 B.n577 B.n576 71.676
R1227 B.n578 B.n416 71.676
R1228 B.n585 B.n584 71.676
R1229 B.n586 B.n414 71.676
R1230 B.n593 B.n592 71.676
R1231 B.n594 B.n412 71.676
R1232 B.n601 B.n600 71.676
R1233 B.n602 B.n410 71.676
R1234 B.n609 B.n608 71.676
R1235 B.n610 B.n408 71.676
R1236 B.n617 B.n616 71.676
R1237 B.n618 B.n406 71.676
R1238 B.n625 B.n624 71.676
R1239 B.n626 B.n404 71.676
R1240 B.n633 B.n632 71.676
R1241 B.n634 B.n402 71.676
R1242 B.n641 B.n640 71.676
R1243 B.n644 B.n643 71.676
R1244 B.n556 B.t21 67.6739
R1245 B.n126 B.t19 67.6739
R1246 B.n428 B.t15 67.6572
R1247 B.n129 B.t12 67.6572
R1248 B.n557 B.n556 59.5399
R1249 B.n537 B.n428 59.5399
R1250 B.n130 B.n129 59.5399
R1251 B.n127 B.n126 59.5399
R1252 B.n649 B.n394 41.1107
R1253 B.n655 B.n394 41.1107
R1254 B.n655 B.n390 41.1107
R1255 B.n662 B.n390 41.1107
R1256 B.n662 B.n661 41.1107
R1257 B.n668 B.n383 41.1107
R1258 B.n674 B.n383 41.1107
R1259 B.n674 B.n379 41.1107
R1260 B.n680 B.n379 41.1107
R1261 B.n680 B.n375 41.1107
R1262 B.n686 B.n375 41.1107
R1263 B.n686 B.n371 41.1107
R1264 B.n692 B.n371 41.1107
R1265 B.n698 B.n367 41.1107
R1266 B.n698 B.n362 41.1107
R1267 B.n704 B.n362 41.1107
R1268 B.n704 B.n363 41.1107
R1269 B.n710 B.n355 41.1107
R1270 B.n716 B.n355 41.1107
R1271 B.n716 B.n351 41.1107
R1272 B.n723 B.n351 41.1107
R1273 B.n723 B.n722 41.1107
R1274 B.n729 B.n344 41.1107
R1275 B.n735 B.n344 41.1107
R1276 B.n735 B.n340 41.1107
R1277 B.n741 B.n340 41.1107
R1278 B.n747 B.n336 41.1107
R1279 B.n747 B.n331 41.1107
R1280 B.n753 B.n331 41.1107
R1281 B.n753 B.n332 41.1107
R1282 B.n760 B.n324 41.1107
R1283 B.n766 B.n324 41.1107
R1284 B.n766 B.n4 41.1107
R1285 B.n905 B.n4 41.1107
R1286 B.n905 B.n904 41.1107
R1287 B.n904 B.n903 41.1107
R1288 B.n903 B.n8 41.1107
R1289 B.n897 B.n8 41.1107
R1290 B.n896 B.n895 41.1107
R1291 B.n895 B.n15 41.1107
R1292 B.n889 B.n15 41.1107
R1293 B.n889 B.n888 41.1107
R1294 B.n887 B.n22 41.1107
R1295 B.n881 B.n22 41.1107
R1296 B.n881 B.n880 41.1107
R1297 B.n880 B.n879 41.1107
R1298 B.n873 B.n32 41.1107
R1299 B.n873 B.n872 41.1107
R1300 B.n872 B.n871 41.1107
R1301 B.n871 B.n36 41.1107
R1302 B.n865 B.n36 41.1107
R1303 B.n864 B.n863 41.1107
R1304 B.n863 B.n43 41.1107
R1305 B.n857 B.n43 41.1107
R1306 B.n857 B.n856 41.1107
R1307 B.n855 B.n50 41.1107
R1308 B.n849 B.n50 41.1107
R1309 B.n849 B.n848 41.1107
R1310 B.n848 B.n847 41.1107
R1311 B.n847 B.n57 41.1107
R1312 B.n841 B.n57 41.1107
R1313 B.n841 B.n840 41.1107
R1314 B.n840 B.n839 41.1107
R1315 B.n833 B.n67 41.1107
R1316 B.n833 B.n832 41.1107
R1317 B.n832 B.n831 41.1107
R1318 B.n831 B.n71 41.1107
R1319 B.n825 B.n71 41.1107
R1320 B.n729 B.t0 40.5061
R1321 B.n879 B.t7 40.5061
R1322 B.n821 B.n820 36.059
R1323 B.n827 B.n73 36.059
R1324 B.n647 B.n646 36.059
R1325 B.n651 B.n396 36.059
R1326 B.n556 B.n555 35.2975
R1327 B.n428 B.n427 35.2975
R1328 B.n129 B.n128 35.2975
R1329 B.n126 B.n125 35.2975
R1330 B.n661 B.t14 30.8331
R1331 B.n67 B.t10 30.8331
R1332 B.n332 B.t6 29.624
R1333 B.t3 B.n896 29.624
R1334 B.t23 B.n367 28.4149
R1335 B.n856 B.t4 28.4149
R1336 B.n363 B.t5 27.2058
R1337 B.t1 B.n864 27.2058
R1338 B.t8 B.n336 25.9967
R1339 B.n888 B.t2 25.9967
R1340 B B.n907 18.0485
R1341 B.n741 B.t8 15.1145
R1342 B.t2 B.n887 15.1145
R1343 B.n710 B.t5 13.9054
R1344 B.n865 B.t1 13.9054
R1345 B.n692 B.t23 12.6963
R1346 B.t4 B.n855 12.6963
R1347 B.n760 B.t6 11.4872
R1348 B.n897 B.t3 11.4872
R1349 B.n131 B.n73 10.6151
R1350 B.n134 B.n131 10.6151
R1351 B.n135 B.n134 10.6151
R1352 B.n138 B.n135 10.6151
R1353 B.n139 B.n138 10.6151
R1354 B.n142 B.n139 10.6151
R1355 B.n143 B.n142 10.6151
R1356 B.n146 B.n143 10.6151
R1357 B.n147 B.n146 10.6151
R1358 B.n150 B.n147 10.6151
R1359 B.n151 B.n150 10.6151
R1360 B.n154 B.n151 10.6151
R1361 B.n155 B.n154 10.6151
R1362 B.n158 B.n155 10.6151
R1363 B.n159 B.n158 10.6151
R1364 B.n162 B.n159 10.6151
R1365 B.n163 B.n162 10.6151
R1366 B.n166 B.n163 10.6151
R1367 B.n167 B.n166 10.6151
R1368 B.n170 B.n167 10.6151
R1369 B.n171 B.n170 10.6151
R1370 B.n174 B.n171 10.6151
R1371 B.n175 B.n174 10.6151
R1372 B.n178 B.n175 10.6151
R1373 B.n179 B.n178 10.6151
R1374 B.n182 B.n179 10.6151
R1375 B.n183 B.n182 10.6151
R1376 B.n186 B.n183 10.6151
R1377 B.n187 B.n186 10.6151
R1378 B.n190 B.n187 10.6151
R1379 B.n191 B.n190 10.6151
R1380 B.n194 B.n191 10.6151
R1381 B.n195 B.n194 10.6151
R1382 B.n198 B.n195 10.6151
R1383 B.n199 B.n198 10.6151
R1384 B.n202 B.n199 10.6151
R1385 B.n203 B.n202 10.6151
R1386 B.n206 B.n203 10.6151
R1387 B.n207 B.n206 10.6151
R1388 B.n210 B.n207 10.6151
R1389 B.n211 B.n210 10.6151
R1390 B.n214 B.n211 10.6151
R1391 B.n215 B.n214 10.6151
R1392 B.n219 B.n218 10.6151
R1393 B.n222 B.n219 10.6151
R1394 B.n223 B.n222 10.6151
R1395 B.n226 B.n223 10.6151
R1396 B.n227 B.n226 10.6151
R1397 B.n230 B.n227 10.6151
R1398 B.n231 B.n230 10.6151
R1399 B.n234 B.n231 10.6151
R1400 B.n235 B.n234 10.6151
R1401 B.n239 B.n238 10.6151
R1402 B.n242 B.n239 10.6151
R1403 B.n243 B.n242 10.6151
R1404 B.n246 B.n243 10.6151
R1405 B.n247 B.n246 10.6151
R1406 B.n250 B.n247 10.6151
R1407 B.n251 B.n250 10.6151
R1408 B.n254 B.n251 10.6151
R1409 B.n255 B.n254 10.6151
R1410 B.n258 B.n255 10.6151
R1411 B.n259 B.n258 10.6151
R1412 B.n262 B.n259 10.6151
R1413 B.n263 B.n262 10.6151
R1414 B.n266 B.n263 10.6151
R1415 B.n267 B.n266 10.6151
R1416 B.n270 B.n267 10.6151
R1417 B.n271 B.n270 10.6151
R1418 B.n274 B.n271 10.6151
R1419 B.n275 B.n274 10.6151
R1420 B.n278 B.n275 10.6151
R1421 B.n279 B.n278 10.6151
R1422 B.n282 B.n279 10.6151
R1423 B.n283 B.n282 10.6151
R1424 B.n286 B.n283 10.6151
R1425 B.n287 B.n286 10.6151
R1426 B.n290 B.n287 10.6151
R1427 B.n291 B.n290 10.6151
R1428 B.n294 B.n291 10.6151
R1429 B.n295 B.n294 10.6151
R1430 B.n298 B.n295 10.6151
R1431 B.n299 B.n298 10.6151
R1432 B.n302 B.n299 10.6151
R1433 B.n303 B.n302 10.6151
R1434 B.n306 B.n303 10.6151
R1435 B.n307 B.n306 10.6151
R1436 B.n310 B.n307 10.6151
R1437 B.n311 B.n310 10.6151
R1438 B.n314 B.n311 10.6151
R1439 B.n315 B.n314 10.6151
R1440 B.n318 B.n315 10.6151
R1441 B.n320 B.n318 10.6151
R1442 B.n321 B.n320 10.6151
R1443 B.n821 B.n321 10.6151
R1444 B.n647 B.n392 10.6151
R1445 B.n657 B.n392 10.6151
R1446 B.n658 B.n657 10.6151
R1447 B.n659 B.n658 10.6151
R1448 B.n659 B.n385 10.6151
R1449 B.n670 B.n385 10.6151
R1450 B.n671 B.n670 10.6151
R1451 B.n672 B.n671 10.6151
R1452 B.n672 B.n377 10.6151
R1453 B.n682 B.n377 10.6151
R1454 B.n683 B.n682 10.6151
R1455 B.n684 B.n683 10.6151
R1456 B.n684 B.n369 10.6151
R1457 B.n694 B.n369 10.6151
R1458 B.n695 B.n694 10.6151
R1459 B.n696 B.n695 10.6151
R1460 B.n696 B.n360 10.6151
R1461 B.n706 B.n360 10.6151
R1462 B.n707 B.n706 10.6151
R1463 B.n708 B.n707 10.6151
R1464 B.n708 B.n353 10.6151
R1465 B.n718 B.n353 10.6151
R1466 B.n719 B.n718 10.6151
R1467 B.n720 B.n719 10.6151
R1468 B.n720 B.n346 10.6151
R1469 B.n731 B.n346 10.6151
R1470 B.n732 B.n731 10.6151
R1471 B.n733 B.n732 10.6151
R1472 B.n733 B.n338 10.6151
R1473 B.n743 B.n338 10.6151
R1474 B.n744 B.n743 10.6151
R1475 B.n745 B.n744 10.6151
R1476 B.n745 B.n329 10.6151
R1477 B.n755 B.n329 10.6151
R1478 B.n756 B.n755 10.6151
R1479 B.n758 B.n756 10.6151
R1480 B.n758 B.n757 10.6151
R1481 B.n757 B.n322 10.6151
R1482 B.n769 B.n322 10.6151
R1483 B.n770 B.n769 10.6151
R1484 B.n771 B.n770 10.6151
R1485 B.n772 B.n771 10.6151
R1486 B.n774 B.n772 10.6151
R1487 B.n775 B.n774 10.6151
R1488 B.n776 B.n775 10.6151
R1489 B.n777 B.n776 10.6151
R1490 B.n779 B.n777 10.6151
R1491 B.n780 B.n779 10.6151
R1492 B.n781 B.n780 10.6151
R1493 B.n782 B.n781 10.6151
R1494 B.n784 B.n782 10.6151
R1495 B.n785 B.n784 10.6151
R1496 B.n786 B.n785 10.6151
R1497 B.n787 B.n786 10.6151
R1498 B.n789 B.n787 10.6151
R1499 B.n790 B.n789 10.6151
R1500 B.n791 B.n790 10.6151
R1501 B.n792 B.n791 10.6151
R1502 B.n794 B.n792 10.6151
R1503 B.n795 B.n794 10.6151
R1504 B.n796 B.n795 10.6151
R1505 B.n797 B.n796 10.6151
R1506 B.n799 B.n797 10.6151
R1507 B.n800 B.n799 10.6151
R1508 B.n801 B.n800 10.6151
R1509 B.n802 B.n801 10.6151
R1510 B.n804 B.n802 10.6151
R1511 B.n805 B.n804 10.6151
R1512 B.n806 B.n805 10.6151
R1513 B.n807 B.n806 10.6151
R1514 B.n809 B.n807 10.6151
R1515 B.n810 B.n809 10.6151
R1516 B.n811 B.n810 10.6151
R1517 B.n812 B.n811 10.6151
R1518 B.n814 B.n812 10.6151
R1519 B.n815 B.n814 10.6151
R1520 B.n816 B.n815 10.6151
R1521 B.n817 B.n816 10.6151
R1522 B.n819 B.n817 10.6151
R1523 B.n820 B.n819 10.6151
R1524 B.n450 B.n396 10.6151
R1525 B.n450 B.n449 10.6151
R1526 B.n456 B.n449 10.6151
R1527 B.n457 B.n456 10.6151
R1528 B.n458 B.n457 10.6151
R1529 B.n458 B.n447 10.6151
R1530 B.n464 B.n447 10.6151
R1531 B.n465 B.n464 10.6151
R1532 B.n466 B.n465 10.6151
R1533 B.n466 B.n445 10.6151
R1534 B.n472 B.n445 10.6151
R1535 B.n473 B.n472 10.6151
R1536 B.n474 B.n473 10.6151
R1537 B.n474 B.n443 10.6151
R1538 B.n480 B.n443 10.6151
R1539 B.n481 B.n480 10.6151
R1540 B.n482 B.n481 10.6151
R1541 B.n482 B.n441 10.6151
R1542 B.n488 B.n441 10.6151
R1543 B.n489 B.n488 10.6151
R1544 B.n490 B.n489 10.6151
R1545 B.n490 B.n439 10.6151
R1546 B.n496 B.n439 10.6151
R1547 B.n497 B.n496 10.6151
R1548 B.n498 B.n497 10.6151
R1549 B.n498 B.n437 10.6151
R1550 B.n504 B.n437 10.6151
R1551 B.n505 B.n504 10.6151
R1552 B.n506 B.n505 10.6151
R1553 B.n506 B.n435 10.6151
R1554 B.n512 B.n435 10.6151
R1555 B.n513 B.n512 10.6151
R1556 B.n514 B.n513 10.6151
R1557 B.n514 B.n433 10.6151
R1558 B.n520 B.n433 10.6151
R1559 B.n521 B.n520 10.6151
R1560 B.n522 B.n521 10.6151
R1561 B.n522 B.n431 10.6151
R1562 B.n528 B.n431 10.6151
R1563 B.n529 B.n528 10.6151
R1564 B.n530 B.n529 10.6151
R1565 B.n530 B.n429 10.6151
R1566 B.n536 B.n429 10.6151
R1567 B.n539 B.n538 10.6151
R1568 B.n539 B.n425 10.6151
R1569 B.n545 B.n425 10.6151
R1570 B.n546 B.n545 10.6151
R1571 B.n547 B.n546 10.6151
R1572 B.n547 B.n423 10.6151
R1573 B.n553 B.n423 10.6151
R1574 B.n554 B.n553 10.6151
R1575 B.n558 B.n554 10.6151
R1576 B.n564 B.n421 10.6151
R1577 B.n565 B.n564 10.6151
R1578 B.n566 B.n565 10.6151
R1579 B.n566 B.n419 10.6151
R1580 B.n572 B.n419 10.6151
R1581 B.n573 B.n572 10.6151
R1582 B.n574 B.n573 10.6151
R1583 B.n574 B.n417 10.6151
R1584 B.n580 B.n417 10.6151
R1585 B.n581 B.n580 10.6151
R1586 B.n582 B.n581 10.6151
R1587 B.n582 B.n415 10.6151
R1588 B.n588 B.n415 10.6151
R1589 B.n589 B.n588 10.6151
R1590 B.n590 B.n589 10.6151
R1591 B.n590 B.n413 10.6151
R1592 B.n596 B.n413 10.6151
R1593 B.n597 B.n596 10.6151
R1594 B.n598 B.n597 10.6151
R1595 B.n598 B.n411 10.6151
R1596 B.n604 B.n411 10.6151
R1597 B.n605 B.n604 10.6151
R1598 B.n606 B.n605 10.6151
R1599 B.n606 B.n409 10.6151
R1600 B.n612 B.n409 10.6151
R1601 B.n613 B.n612 10.6151
R1602 B.n614 B.n613 10.6151
R1603 B.n614 B.n407 10.6151
R1604 B.n620 B.n407 10.6151
R1605 B.n621 B.n620 10.6151
R1606 B.n622 B.n621 10.6151
R1607 B.n622 B.n405 10.6151
R1608 B.n628 B.n405 10.6151
R1609 B.n629 B.n628 10.6151
R1610 B.n630 B.n629 10.6151
R1611 B.n630 B.n403 10.6151
R1612 B.n636 B.n403 10.6151
R1613 B.n637 B.n636 10.6151
R1614 B.n638 B.n637 10.6151
R1615 B.n638 B.n401 10.6151
R1616 B.n401 B.n400 10.6151
R1617 B.n645 B.n400 10.6151
R1618 B.n646 B.n645 10.6151
R1619 B.n652 B.n651 10.6151
R1620 B.n653 B.n652 10.6151
R1621 B.n653 B.n388 10.6151
R1622 B.n664 B.n388 10.6151
R1623 B.n665 B.n664 10.6151
R1624 B.n666 B.n665 10.6151
R1625 B.n666 B.n381 10.6151
R1626 B.n676 B.n381 10.6151
R1627 B.n677 B.n676 10.6151
R1628 B.n678 B.n677 10.6151
R1629 B.n678 B.n373 10.6151
R1630 B.n688 B.n373 10.6151
R1631 B.n689 B.n688 10.6151
R1632 B.n690 B.n689 10.6151
R1633 B.n690 B.n365 10.6151
R1634 B.n700 B.n365 10.6151
R1635 B.n701 B.n700 10.6151
R1636 B.n702 B.n701 10.6151
R1637 B.n702 B.n357 10.6151
R1638 B.n712 B.n357 10.6151
R1639 B.n713 B.n712 10.6151
R1640 B.n714 B.n713 10.6151
R1641 B.n714 B.n349 10.6151
R1642 B.n725 B.n349 10.6151
R1643 B.n726 B.n725 10.6151
R1644 B.n727 B.n726 10.6151
R1645 B.n727 B.n342 10.6151
R1646 B.n737 B.n342 10.6151
R1647 B.n738 B.n737 10.6151
R1648 B.n739 B.n738 10.6151
R1649 B.n739 B.n334 10.6151
R1650 B.n749 B.n334 10.6151
R1651 B.n750 B.n749 10.6151
R1652 B.n751 B.n750 10.6151
R1653 B.n751 B.n326 10.6151
R1654 B.n762 B.n326 10.6151
R1655 B.n763 B.n762 10.6151
R1656 B.n764 B.n763 10.6151
R1657 B.n764 B.n0 10.6151
R1658 B.n901 B.n1 10.6151
R1659 B.n901 B.n900 10.6151
R1660 B.n900 B.n899 10.6151
R1661 B.n899 B.n10 10.6151
R1662 B.n893 B.n10 10.6151
R1663 B.n893 B.n892 10.6151
R1664 B.n892 B.n891 10.6151
R1665 B.n891 B.n17 10.6151
R1666 B.n885 B.n17 10.6151
R1667 B.n885 B.n884 10.6151
R1668 B.n884 B.n883 10.6151
R1669 B.n883 B.n24 10.6151
R1670 B.n877 B.n24 10.6151
R1671 B.n877 B.n876 10.6151
R1672 B.n876 B.n875 10.6151
R1673 B.n875 B.n30 10.6151
R1674 B.n869 B.n30 10.6151
R1675 B.n869 B.n868 10.6151
R1676 B.n868 B.n867 10.6151
R1677 B.n867 B.n38 10.6151
R1678 B.n861 B.n38 10.6151
R1679 B.n861 B.n860 10.6151
R1680 B.n860 B.n859 10.6151
R1681 B.n859 B.n45 10.6151
R1682 B.n853 B.n45 10.6151
R1683 B.n853 B.n852 10.6151
R1684 B.n852 B.n851 10.6151
R1685 B.n851 B.n52 10.6151
R1686 B.n845 B.n52 10.6151
R1687 B.n845 B.n844 10.6151
R1688 B.n844 B.n843 10.6151
R1689 B.n843 B.n59 10.6151
R1690 B.n837 B.n59 10.6151
R1691 B.n837 B.n836 10.6151
R1692 B.n836 B.n835 10.6151
R1693 B.n835 B.n65 10.6151
R1694 B.n829 B.n65 10.6151
R1695 B.n829 B.n828 10.6151
R1696 B.n828 B.n827 10.6151
R1697 B.n668 B.t14 10.278
R1698 B.n839 B.t10 10.278
R1699 B.n215 B.n130 9.36635
R1700 B.n238 B.n127 9.36635
R1701 B.n537 B.n536 9.36635
R1702 B.n557 B.n421 9.36635
R1703 B.n907 B.n0 2.81026
R1704 B.n907 B.n1 2.81026
R1705 B.n218 B.n130 1.24928
R1706 B.n235 B.n127 1.24928
R1707 B.n538 B.n537 1.24928
R1708 B.n558 B.n557 1.24928
R1709 B.n722 B.t0 0.605062
R1710 B.n32 B.t7 0.605062
R1711 VN.n7 VN.t3 241.106
R1712 VN.n34 VN.t7 241.106
R1713 VN.n12 VN.t6 208.976
R1714 VN.n6 VN.t5 208.976
R1715 VN.n18 VN.t8 208.976
R1716 VN.n25 VN.t9 208.976
R1717 VN.n39 VN.t4 208.976
R1718 VN.n33 VN.t1 208.976
R1719 VN.n45 VN.t0 208.976
R1720 VN.n52 VN.t2 208.976
R1721 VN.n26 VN.n25 179.006
R1722 VN.n53 VN.n52 179.006
R1723 VN.n51 VN.n27 161.3
R1724 VN.n50 VN.n49 161.3
R1725 VN.n48 VN.n28 161.3
R1726 VN.n47 VN.n46 161.3
R1727 VN.n44 VN.n29 161.3
R1728 VN.n43 VN.n42 161.3
R1729 VN.n41 VN.n30 161.3
R1730 VN.n40 VN.n39 161.3
R1731 VN.n38 VN.n31 161.3
R1732 VN.n37 VN.n36 161.3
R1733 VN.n35 VN.n32 161.3
R1734 VN.n24 VN.n0 161.3
R1735 VN.n23 VN.n22 161.3
R1736 VN.n21 VN.n1 161.3
R1737 VN.n20 VN.n19 161.3
R1738 VN.n17 VN.n2 161.3
R1739 VN.n16 VN.n15 161.3
R1740 VN.n14 VN.n3 161.3
R1741 VN.n13 VN.n12 161.3
R1742 VN.n11 VN.n4 161.3
R1743 VN.n10 VN.n9 161.3
R1744 VN.n8 VN.n5 161.3
R1745 VN.n23 VN.n1 56.5617
R1746 VN.n50 VN.n28 56.5617
R1747 VN.n7 VN.n6 50.5334
R1748 VN.n34 VN.n33 50.5334
R1749 VN.n11 VN.n10 49.296
R1750 VN.n16 VN.n3 49.296
R1751 VN.n38 VN.n37 49.296
R1752 VN.n43 VN.n30 49.296
R1753 VN VN.n53 48.0327
R1754 VN.n10 VN.n5 31.8581
R1755 VN.n17 VN.n16 31.8581
R1756 VN.n37 VN.n32 31.8581
R1757 VN.n44 VN.n43 31.8581
R1758 VN.n12 VN.n11 24.5923
R1759 VN.n12 VN.n3 24.5923
R1760 VN.n19 VN.n1 24.5923
R1761 VN.n24 VN.n23 24.5923
R1762 VN.n39 VN.n30 24.5923
R1763 VN.n39 VN.n38 24.5923
R1764 VN.n46 VN.n28 24.5923
R1765 VN.n51 VN.n50 24.5923
R1766 VN.n35 VN.n34 18.0715
R1767 VN.n8 VN.n7 18.0715
R1768 VN.n6 VN.n5 15.7393
R1769 VN.n18 VN.n17 15.7393
R1770 VN.n33 VN.n32 15.7393
R1771 VN.n45 VN.n44 15.7393
R1772 VN.n19 VN.n18 8.85356
R1773 VN.n46 VN.n45 8.85356
R1774 VN.n25 VN.n24 6.88621
R1775 VN.n52 VN.n51 6.88621
R1776 VN.n53 VN.n27 0.189894
R1777 VN.n49 VN.n27 0.189894
R1778 VN.n49 VN.n48 0.189894
R1779 VN.n48 VN.n47 0.189894
R1780 VN.n47 VN.n29 0.189894
R1781 VN.n42 VN.n29 0.189894
R1782 VN.n42 VN.n41 0.189894
R1783 VN.n41 VN.n40 0.189894
R1784 VN.n40 VN.n31 0.189894
R1785 VN.n36 VN.n31 0.189894
R1786 VN.n36 VN.n35 0.189894
R1787 VN.n9 VN.n8 0.189894
R1788 VN.n9 VN.n4 0.189894
R1789 VN.n13 VN.n4 0.189894
R1790 VN.n14 VN.n13 0.189894
R1791 VN.n15 VN.n14 0.189894
R1792 VN.n15 VN.n2 0.189894
R1793 VN.n20 VN.n2 0.189894
R1794 VN.n21 VN.n20 0.189894
R1795 VN.n22 VN.n21 0.189894
R1796 VN.n22 VN.n0 0.189894
R1797 VN.n26 VN.n0 0.189894
R1798 VN VN.n26 0.0516364
R1799 VDD2.n1 VDD2.t6 65.8288
R1800 VDD2.n4 VDD2.t7 64.261
R1801 VDD2.n3 VDD2.n2 63.8487
R1802 VDD2 VDD2.n7 63.8459
R1803 VDD2.n6 VDD2.n5 62.7285
R1804 VDD2.n1 VDD2.n0 62.7273
R1805 VDD2.n4 VDD2.n3 42.3058
R1806 VDD2.n6 VDD2.n4 1.56947
R1807 VDD2.n7 VDD2.t8 1.53301
R1808 VDD2.n7 VDD2.t2 1.53301
R1809 VDD2.n5 VDD2.t9 1.53301
R1810 VDD2.n5 VDD2.t5 1.53301
R1811 VDD2.n2 VDD2.t1 1.53301
R1812 VDD2.n2 VDD2.t0 1.53301
R1813 VDD2.n0 VDD2.t4 1.53301
R1814 VDD2.n0 VDD2.t3 1.53301
R1815 VDD2 VDD2.n6 0.450931
R1816 VDD2.n3 VDD2.n1 0.337395
C0 VTAIL VDD2 11.5538f
C1 VDD1 VP 10.194799f
C2 VDD1 VN 0.151154f
C3 VDD1 VTAIL 11.5124f
C4 VDD1 VDD2 1.45293f
C5 VP VN 6.92956f
C6 VP VTAIL 10.0645f
C7 VP VDD2 0.442531f
C8 VTAIL VN 10.05f
C9 VN VDD2 9.90775f
C10 VDD2 B 6.068429f
C11 VDD1 B 6.042821f
C12 VTAIL B 7.64399f
C13 VN B 13.03858f
C14 VP B 11.364157f
C15 VDD2.t6 B 2.64141f
C16 VDD2.t4 B 0.229911f
C17 VDD2.t3 B 0.229911f
C18 VDD2.n0 B 2.06445f
C19 VDD2.n1 B 0.673799f
C20 VDD2.t1 B 0.229911f
C21 VDD2.t0 B 0.229911f
C22 VDD2.n2 B 2.07122f
C23 VDD2.n3 B 2.13833f
C24 VDD2.t7 B 2.63279f
C25 VDD2.n4 B 2.48438f
C26 VDD2.t9 B 0.229911f
C27 VDD2.t5 B 0.229911f
C28 VDD2.n5 B 2.06446f
C29 VDD2.n6 B 0.327006f
C30 VDD2.t8 B 0.229911f
C31 VDD2.t2 B 0.229911f
C32 VDD2.n7 B 2.07119f
C33 VN.n0 B 0.029903f
C34 VN.t9 B 1.57164f
C35 VN.n1 B 0.041814f
C36 VN.n2 B 0.029903f
C37 VN.t8 B 1.57164f
C38 VN.n3 B 0.055178f
C39 VN.n4 B 0.029903f
C40 VN.t6 B 1.57164f
C41 VN.n5 B 0.049968f
C42 VN.t3 B 1.66207f
C43 VN.t5 B 1.57164f
C44 VN.n6 B 0.623814f
C45 VN.n7 B 0.636134f
C46 VN.n8 B 0.187457f
C47 VN.n9 B 0.029903f
C48 VN.n10 B 0.027389f
C49 VN.n11 B 0.055178f
C50 VN.n12 B 0.593206f
C51 VN.n13 B 0.029903f
C52 VN.n14 B 0.029903f
C53 VN.n15 B 0.029903f
C54 VN.n16 B 0.027389f
C55 VN.n17 B 0.049968f
C56 VN.n18 B 0.565129f
C57 VN.n19 B 0.037932f
C58 VN.n20 B 0.029903f
C59 VN.n21 B 0.029903f
C60 VN.n22 B 0.029903f
C61 VN.n23 B 0.045123f
C62 VN.n24 B 0.035742f
C63 VN.n25 B 0.62151f
C64 VN.n26 B 0.029363f
C65 VN.n27 B 0.029903f
C66 VN.t2 B 1.57164f
C67 VN.n28 B 0.041814f
C68 VN.n29 B 0.029903f
C69 VN.t0 B 1.57164f
C70 VN.n30 B 0.055178f
C71 VN.n31 B 0.029903f
C72 VN.t4 B 1.57164f
C73 VN.n32 B 0.049968f
C74 VN.t7 B 1.66207f
C75 VN.t1 B 1.57164f
C76 VN.n33 B 0.623814f
C77 VN.n34 B 0.636134f
C78 VN.n35 B 0.187457f
C79 VN.n36 B 0.029903f
C80 VN.n37 B 0.027389f
C81 VN.n38 B 0.055178f
C82 VN.n39 B 0.593206f
C83 VN.n40 B 0.029903f
C84 VN.n41 B 0.029903f
C85 VN.n42 B 0.029903f
C86 VN.n43 B 0.027389f
C87 VN.n44 B 0.049968f
C88 VN.n45 B 0.565129f
C89 VN.n46 B 0.037932f
C90 VN.n47 B 0.029903f
C91 VN.n48 B 0.029903f
C92 VN.n49 B 0.029903f
C93 VN.n50 B 0.045123f
C94 VN.n51 B 0.035742f
C95 VN.n52 B 0.62151f
C96 VN.n53 B 1.53657f
C97 VDD1.t7 B 2.65572f
C98 VDD1.t2 B 0.231156f
C99 VDD1.t9 B 0.231156f
C100 VDD1.n0 B 2.07564f
C101 VDD1.n1 B 0.684155f
C102 VDD1.t8 B 2.65571f
C103 VDD1.t0 B 0.231156f
C104 VDD1.t4 B 0.231156f
C105 VDD1.n2 B 2.07563f
C106 VDD1.n3 B 0.677446f
C107 VDD1.t1 B 0.231156f
C108 VDD1.t5 B 0.231156f
C109 VDD1.n4 B 2.08243f
C110 VDD1.n5 B 2.23742f
C111 VDD1.t6 B 0.231156f
C112 VDD1.t3 B 0.231156f
C113 VDD1.n6 B 2.07563f
C114 VDD1.n7 B 2.51652f
C115 VTAIL.t3 B 0.24836f
C116 VTAIL.t2 B 0.24836f
C117 VTAIL.n0 B 2.16117f
C118 VTAIL.n1 B 0.425956f
C119 VTAIL.t9 B 2.75509f
C120 VTAIL.n2 B 0.535568f
C121 VTAIL.t12 B 0.24836f
C122 VTAIL.t14 B 0.24836f
C123 VTAIL.n3 B 2.16117f
C124 VTAIL.n4 B 0.476804f
C125 VTAIL.t18 B 0.24836f
C126 VTAIL.t11 B 0.24836f
C127 VTAIL.n5 B 2.16117f
C128 VTAIL.n6 B 1.80324f
C129 VTAIL.t19 B 0.24836f
C130 VTAIL.t5 B 0.24836f
C131 VTAIL.n7 B 2.16118f
C132 VTAIL.n8 B 1.80323f
C133 VTAIL.t0 B 0.24836f
C134 VTAIL.t8 B 0.24836f
C135 VTAIL.n9 B 2.16118f
C136 VTAIL.n10 B 0.476793f
C137 VTAIL.t6 B 2.75511f
C138 VTAIL.n11 B 0.535551f
C139 VTAIL.t10 B 0.24836f
C140 VTAIL.t13 B 0.24836f
C141 VTAIL.n12 B 2.16118f
C142 VTAIL.n13 B 0.452129f
C143 VTAIL.t17 B 0.24836f
C144 VTAIL.t16 B 0.24836f
C145 VTAIL.n14 B 2.16118f
C146 VTAIL.n15 B 0.476793f
C147 VTAIL.t15 B 2.75509f
C148 VTAIL.n16 B 1.76369f
C149 VTAIL.t4 B 2.75509f
C150 VTAIL.n17 B 1.76369f
C151 VTAIL.t7 B 0.24836f
C152 VTAIL.t1 B 0.24836f
C153 VTAIL.n18 B 2.16117f
C154 VTAIL.n19 B 0.380008f
C155 VP.n0 B 0.030284f
C156 VP.t4 B 1.59165f
C157 VP.n1 B 0.042346f
C158 VP.n2 B 0.030284f
C159 VP.t8 B 1.59165f
C160 VP.n3 B 0.055881f
C161 VP.n4 B 0.030284f
C162 VP.t5 B 1.59165f
C163 VP.n5 B 0.050604f
C164 VP.n6 B 0.030284f
C165 VP.n7 B 0.036197f
C166 VP.n8 B 0.030284f
C167 VP.t6 B 1.59165f
C168 VP.n9 B 0.042346f
C169 VP.n10 B 0.030284f
C170 VP.t3 B 1.59165f
C171 VP.n11 B 0.055881f
C172 VP.n12 B 0.030284f
C173 VP.t0 B 1.59165f
C174 VP.n13 B 0.050604f
C175 VP.t2 B 1.68324f
C176 VP.t7 B 1.59165f
C177 VP.n14 B 0.631758f
C178 VP.n15 B 0.644235f
C179 VP.n16 B 0.189845f
C180 VP.n17 B 0.030284f
C181 VP.n18 B 0.027738f
C182 VP.n19 B 0.055881f
C183 VP.n20 B 0.600761f
C184 VP.n21 B 0.030284f
C185 VP.n22 B 0.030284f
C186 VP.n23 B 0.030284f
C187 VP.n24 B 0.027738f
C188 VP.n25 B 0.050604f
C189 VP.n26 B 0.572326f
C190 VP.n27 B 0.038415f
C191 VP.n28 B 0.030284f
C192 VP.n29 B 0.030284f
C193 VP.n30 B 0.030284f
C194 VP.n31 B 0.045698f
C195 VP.n32 B 0.036197f
C196 VP.n33 B 0.629425f
C197 VP.n34 B 1.5364f
C198 VP.t1 B 1.59165f
C199 VP.n35 B 0.629425f
C200 VP.n36 B 1.55931f
C201 VP.n37 B 0.030284f
C202 VP.n38 B 0.030284f
C203 VP.n39 B 0.045698f
C204 VP.n40 B 0.042346f
C205 VP.t9 B 1.59165f
C206 VP.n41 B 0.572326f
C207 VP.n42 B 0.038415f
C208 VP.n43 B 0.030284f
C209 VP.n44 B 0.030284f
C210 VP.n45 B 0.030284f
C211 VP.n46 B 0.027738f
C212 VP.n47 B 0.055881f
C213 VP.n48 B 0.600761f
C214 VP.n49 B 0.030284f
C215 VP.n50 B 0.030284f
C216 VP.n51 B 0.030284f
C217 VP.n52 B 0.027738f
C218 VP.n53 B 0.050604f
C219 VP.n54 B 0.572326f
C220 VP.n55 B 0.038415f
C221 VP.n56 B 0.030284f
C222 VP.n57 B 0.030284f
C223 VP.n58 B 0.030284f
C224 VP.n59 B 0.045698f
C225 VP.n60 B 0.036197f
C226 VP.n61 B 0.629425f
C227 VP.n62 B 0.029737f
.ends

