* NGSPICE file created from diff_pair_sample_1235.ext - technology: sky130A

.subckt diff_pair_sample_1235 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=7.605 ps=39.78 w=19.5 l=3.03
X1 VTAIL.t3 VN.t0 VDD2.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X2 VTAIL.t19 VP.t1 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X3 VDD1.t7 VP.t2 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X4 VTAIL.t17 VP.t3 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X5 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X6 VDD2.t7 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=3.2175 ps=19.83 w=19.5 l=3.03
X7 VDD2.t6 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=3.2175 ps=19.83 w=19.5 l=3.03
X8 VDD1.t5 VP.t4 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=7.605 ps=39.78 w=19.5 l=3.03
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=0 ps=0 w=19.5 l=3.03
X10 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=7.605 ps=39.78 w=19.5 l=3.03
X11 VDD1.t4 VP.t5 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=3.2175 ps=19.83 w=19.5 l=3.03
X12 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X13 VDD2.t3 VN.t6 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X14 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=0 ps=0 w=19.5 l=3.03
X15 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=7.605 ps=39.78 w=19.5 l=3.03
X16 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X17 VTAIL.t10 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=0 ps=0 w=19.5 l=3.03
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=0 ps=0 w=19.5 l=3.03
X20 VTAIL.t4 VN.t9 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X21 VDD1.t2 VP.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=7.605 pd=39.78 as=3.2175 ps=19.83 w=19.5 l=3.03
X22 VDD1.t1 VP.t8 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
X23 VTAIL.t13 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2175 pd=19.83 as=3.2175 ps=19.83 w=19.5 l=3.03
R0 VP.n26 VP.t7 186.941
R1 VP.n27 VP.n24 161.3
R2 VP.n29 VP.n28 161.3
R3 VP.n30 VP.n23 161.3
R4 VP.n32 VP.n31 161.3
R5 VP.n33 VP.n22 161.3
R6 VP.n35 VP.n34 161.3
R7 VP.n36 VP.n21 161.3
R8 VP.n39 VP.n38 161.3
R9 VP.n40 VP.n20 161.3
R10 VP.n42 VP.n41 161.3
R11 VP.n43 VP.n19 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n18 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n50 VP.n17 161.3
R16 VP.n52 VP.n51 161.3
R17 VP.n53 VP.n16 161.3
R18 VP.n55 VP.n54 161.3
R19 VP.n56 VP.n15 161.3
R20 VP.n58 VP.n57 161.3
R21 VP.n103 VP.n102 161.3
R22 VP.n101 VP.n1 161.3
R23 VP.n100 VP.n99 161.3
R24 VP.n98 VP.n2 161.3
R25 VP.n97 VP.n96 161.3
R26 VP.n95 VP.n3 161.3
R27 VP.n93 VP.n92 161.3
R28 VP.n91 VP.n4 161.3
R29 VP.n90 VP.n89 161.3
R30 VP.n88 VP.n5 161.3
R31 VP.n87 VP.n86 161.3
R32 VP.n85 VP.n6 161.3
R33 VP.n84 VP.n83 161.3
R34 VP.n81 VP.n7 161.3
R35 VP.n80 VP.n79 161.3
R36 VP.n78 VP.n8 161.3
R37 VP.n77 VP.n76 161.3
R38 VP.n75 VP.n9 161.3
R39 VP.n74 VP.n73 161.3
R40 VP.n72 VP.n10 161.3
R41 VP.n71 VP.n70 161.3
R42 VP.n68 VP.n11 161.3
R43 VP.n67 VP.n66 161.3
R44 VP.n65 VP.n12 161.3
R45 VP.n64 VP.n63 161.3
R46 VP.n62 VP.n13 161.3
R47 VP.n61 VP.t5 155.1
R48 VP.n69 VP.t1 155.1
R49 VP.n82 VP.t8 155.1
R50 VP.n94 VP.t9 155.1
R51 VP.n0 VP.t4 155.1
R52 VP.n14 VP.t0 155.1
R53 VP.n49 VP.t3 155.1
R54 VP.n37 VP.t2 155.1
R55 VP.n25 VP.t6 155.1
R56 VP.n26 VP.n25 68.6895
R57 VP.n61 VP.n60 67.1292
R58 VP.n104 VP.n0 67.1292
R59 VP.n59 VP.n14 67.1292
R60 VP.n60 VP.n59 61.3102
R61 VP.n67 VP.n12 56.5617
R62 VP.n100 VP.n2 56.5617
R63 VP.n55 VP.n16 56.5617
R64 VP.n76 VP.n8 47.3584
R65 VP.n88 VP.n87 47.3584
R66 VP.n43 VP.n42 47.3584
R67 VP.n31 VP.n22 47.3584
R68 VP.n76 VP.n75 33.7956
R69 VP.n89 VP.n88 33.7956
R70 VP.n44 VP.n43 33.7956
R71 VP.n31 VP.n30 33.7956
R72 VP.n63 VP.n62 24.5923
R73 VP.n63 VP.n12 24.5923
R74 VP.n68 VP.n67 24.5923
R75 VP.n70 VP.n68 24.5923
R76 VP.n74 VP.n10 24.5923
R77 VP.n75 VP.n74 24.5923
R78 VP.n80 VP.n8 24.5923
R79 VP.n81 VP.n80 24.5923
R80 VP.n83 VP.n6 24.5923
R81 VP.n87 VP.n6 24.5923
R82 VP.n89 VP.n4 24.5923
R83 VP.n93 VP.n4 24.5923
R84 VP.n96 VP.n95 24.5923
R85 VP.n96 VP.n2 24.5923
R86 VP.n101 VP.n100 24.5923
R87 VP.n102 VP.n101 24.5923
R88 VP.n56 VP.n55 24.5923
R89 VP.n57 VP.n56 24.5923
R90 VP.n44 VP.n18 24.5923
R91 VP.n48 VP.n18 24.5923
R92 VP.n51 VP.n50 24.5923
R93 VP.n51 VP.n16 24.5923
R94 VP.n35 VP.n22 24.5923
R95 VP.n36 VP.n35 24.5923
R96 VP.n38 VP.n20 24.5923
R97 VP.n42 VP.n20 24.5923
R98 VP.n29 VP.n24 24.5923
R99 VP.n30 VP.n29 24.5923
R100 VP.n62 VP.n61 23.1168
R101 VP.n102 VP.n0 23.1168
R102 VP.n57 VP.n14 23.1168
R103 VP.n70 VP.n69 19.1821
R104 VP.n95 VP.n94 19.1821
R105 VP.n50 VP.n49 19.1821
R106 VP.n82 VP.n81 12.2964
R107 VP.n83 VP.n82 12.2964
R108 VP.n37 VP.n36 12.2964
R109 VP.n38 VP.n37 12.2964
R110 VP.n69 VP.n10 5.4107
R111 VP.n94 VP.n93 5.4107
R112 VP.n49 VP.n48 5.4107
R113 VP.n25 VP.n24 5.4107
R114 VP.n27 VP.n26 5.32097
R115 VP.n59 VP.n58 0.354861
R116 VP.n60 VP.n13 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VTAIL.n432 VTAIL.n332 214.453
R164 VTAIL.n102 VTAIL.n2 214.453
R165 VTAIL.n326 VTAIL.n226 214.453
R166 VTAIL.n216 VTAIL.n116 214.453
R167 VTAIL.n367 VTAIL.n366 185
R168 VTAIL.n364 VTAIL.n363 185
R169 VTAIL.n373 VTAIL.n372 185
R170 VTAIL.n375 VTAIL.n374 185
R171 VTAIL.n360 VTAIL.n359 185
R172 VTAIL.n381 VTAIL.n380 185
R173 VTAIL.n384 VTAIL.n383 185
R174 VTAIL.n382 VTAIL.n356 185
R175 VTAIL.n389 VTAIL.n355 185
R176 VTAIL.n391 VTAIL.n390 185
R177 VTAIL.n393 VTAIL.n392 185
R178 VTAIL.n352 VTAIL.n351 185
R179 VTAIL.n399 VTAIL.n398 185
R180 VTAIL.n401 VTAIL.n400 185
R181 VTAIL.n348 VTAIL.n347 185
R182 VTAIL.n407 VTAIL.n406 185
R183 VTAIL.n409 VTAIL.n408 185
R184 VTAIL.n344 VTAIL.n343 185
R185 VTAIL.n415 VTAIL.n414 185
R186 VTAIL.n417 VTAIL.n416 185
R187 VTAIL.n340 VTAIL.n339 185
R188 VTAIL.n423 VTAIL.n422 185
R189 VTAIL.n425 VTAIL.n424 185
R190 VTAIL.n336 VTAIL.n335 185
R191 VTAIL.n431 VTAIL.n430 185
R192 VTAIL.n433 VTAIL.n432 185
R193 VTAIL.n37 VTAIL.n36 185
R194 VTAIL.n34 VTAIL.n33 185
R195 VTAIL.n43 VTAIL.n42 185
R196 VTAIL.n45 VTAIL.n44 185
R197 VTAIL.n30 VTAIL.n29 185
R198 VTAIL.n51 VTAIL.n50 185
R199 VTAIL.n54 VTAIL.n53 185
R200 VTAIL.n52 VTAIL.n26 185
R201 VTAIL.n59 VTAIL.n25 185
R202 VTAIL.n61 VTAIL.n60 185
R203 VTAIL.n63 VTAIL.n62 185
R204 VTAIL.n22 VTAIL.n21 185
R205 VTAIL.n69 VTAIL.n68 185
R206 VTAIL.n71 VTAIL.n70 185
R207 VTAIL.n18 VTAIL.n17 185
R208 VTAIL.n77 VTAIL.n76 185
R209 VTAIL.n79 VTAIL.n78 185
R210 VTAIL.n14 VTAIL.n13 185
R211 VTAIL.n85 VTAIL.n84 185
R212 VTAIL.n87 VTAIL.n86 185
R213 VTAIL.n10 VTAIL.n9 185
R214 VTAIL.n93 VTAIL.n92 185
R215 VTAIL.n95 VTAIL.n94 185
R216 VTAIL.n6 VTAIL.n5 185
R217 VTAIL.n101 VTAIL.n100 185
R218 VTAIL.n103 VTAIL.n102 185
R219 VTAIL.n327 VTAIL.n326 185
R220 VTAIL.n325 VTAIL.n324 185
R221 VTAIL.n230 VTAIL.n229 185
R222 VTAIL.n319 VTAIL.n318 185
R223 VTAIL.n317 VTAIL.n316 185
R224 VTAIL.n234 VTAIL.n233 185
R225 VTAIL.n311 VTAIL.n310 185
R226 VTAIL.n309 VTAIL.n308 185
R227 VTAIL.n238 VTAIL.n237 185
R228 VTAIL.n303 VTAIL.n302 185
R229 VTAIL.n301 VTAIL.n300 185
R230 VTAIL.n242 VTAIL.n241 185
R231 VTAIL.n295 VTAIL.n294 185
R232 VTAIL.n293 VTAIL.n292 185
R233 VTAIL.n246 VTAIL.n245 185
R234 VTAIL.n287 VTAIL.n286 185
R235 VTAIL.n285 VTAIL.n284 185
R236 VTAIL.n283 VTAIL.n249 185
R237 VTAIL.n253 VTAIL.n250 185
R238 VTAIL.n278 VTAIL.n277 185
R239 VTAIL.n276 VTAIL.n275 185
R240 VTAIL.n255 VTAIL.n254 185
R241 VTAIL.n270 VTAIL.n269 185
R242 VTAIL.n268 VTAIL.n267 185
R243 VTAIL.n259 VTAIL.n258 185
R244 VTAIL.n262 VTAIL.n261 185
R245 VTAIL.n217 VTAIL.n216 185
R246 VTAIL.n215 VTAIL.n214 185
R247 VTAIL.n120 VTAIL.n119 185
R248 VTAIL.n209 VTAIL.n208 185
R249 VTAIL.n207 VTAIL.n206 185
R250 VTAIL.n124 VTAIL.n123 185
R251 VTAIL.n201 VTAIL.n200 185
R252 VTAIL.n199 VTAIL.n198 185
R253 VTAIL.n128 VTAIL.n127 185
R254 VTAIL.n193 VTAIL.n192 185
R255 VTAIL.n191 VTAIL.n190 185
R256 VTAIL.n132 VTAIL.n131 185
R257 VTAIL.n185 VTAIL.n184 185
R258 VTAIL.n183 VTAIL.n182 185
R259 VTAIL.n136 VTAIL.n135 185
R260 VTAIL.n177 VTAIL.n176 185
R261 VTAIL.n175 VTAIL.n174 185
R262 VTAIL.n173 VTAIL.n139 185
R263 VTAIL.n143 VTAIL.n140 185
R264 VTAIL.n168 VTAIL.n167 185
R265 VTAIL.n166 VTAIL.n165 185
R266 VTAIL.n145 VTAIL.n144 185
R267 VTAIL.n160 VTAIL.n159 185
R268 VTAIL.n158 VTAIL.n157 185
R269 VTAIL.n149 VTAIL.n148 185
R270 VTAIL.n152 VTAIL.n151 185
R271 VTAIL.t1 VTAIL.n365 149.524
R272 VTAIL.t18 VTAIL.n35 149.524
R273 VTAIL.t14 VTAIL.n260 149.524
R274 VTAIL.t5 VTAIL.n150 149.524
R275 VTAIL.n366 VTAIL.n363 104.615
R276 VTAIL.n373 VTAIL.n363 104.615
R277 VTAIL.n374 VTAIL.n373 104.615
R278 VTAIL.n374 VTAIL.n359 104.615
R279 VTAIL.n381 VTAIL.n359 104.615
R280 VTAIL.n383 VTAIL.n381 104.615
R281 VTAIL.n383 VTAIL.n382 104.615
R282 VTAIL.n382 VTAIL.n355 104.615
R283 VTAIL.n391 VTAIL.n355 104.615
R284 VTAIL.n392 VTAIL.n391 104.615
R285 VTAIL.n392 VTAIL.n351 104.615
R286 VTAIL.n399 VTAIL.n351 104.615
R287 VTAIL.n400 VTAIL.n399 104.615
R288 VTAIL.n400 VTAIL.n347 104.615
R289 VTAIL.n407 VTAIL.n347 104.615
R290 VTAIL.n408 VTAIL.n407 104.615
R291 VTAIL.n408 VTAIL.n343 104.615
R292 VTAIL.n415 VTAIL.n343 104.615
R293 VTAIL.n416 VTAIL.n415 104.615
R294 VTAIL.n416 VTAIL.n339 104.615
R295 VTAIL.n423 VTAIL.n339 104.615
R296 VTAIL.n424 VTAIL.n423 104.615
R297 VTAIL.n424 VTAIL.n335 104.615
R298 VTAIL.n431 VTAIL.n335 104.615
R299 VTAIL.n432 VTAIL.n431 104.615
R300 VTAIL.n36 VTAIL.n33 104.615
R301 VTAIL.n43 VTAIL.n33 104.615
R302 VTAIL.n44 VTAIL.n43 104.615
R303 VTAIL.n44 VTAIL.n29 104.615
R304 VTAIL.n51 VTAIL.n29 104.615
R305 VTAIL.n53 VTAIL.n51 104.615
R306 VTAIL.n53 VTAIL.n52 104.615
R307 VTAIL.n52 VTAIL.n25 104.615
R308 VTAIL.n61 VTAIL.n25 104.615
R309 VTAIL.n62 VTAIL.n61 104.615
R310 VTAIL.n62 VTAIL.n21 104.615
R311 VTAIL.n69 VTAIL.n21 104.615
R312 VTAIL.n70 VTAIL.n69 104.615
R313 VTAIL.n70 VTAIL.n17 104.615
R314 VTAIL.n77 VTAIL.n17 104.615
R315 VTAIL.n78 VTAIL.n77 104.615
R316 VTAIL.n78 VTAIL.n13 104.615
R317 VTAIL.n85 VTAIL.n13 104.615
R318 VTAIL.n86 VTAIL.n85 104.615
R319 VTAIL.n86 VTAIL.n9 104.615
R320 VTAIL.n93 VTAIL.n9 104.615
R321 VTAIL.n94 VTAIL.n93 104.615
R322 VTAIL.n94 VTAIL.n5 104.615
R323 VTAIL.n101 VTAIL.n5 104.615
R324 VTAIL.n102 VTAIL.n101 104.615
R325 VTAIL.n326 VTAIL.n325 104.615
R326 VTAIL.n325 VTAIL.n229 104.615
R327 VTAIL.n318 VTAIL.n229 104.615
R328 VTAIL.n318 VTAIL.n317 104.615
R329 VTAIL.n317 VTAIL.n233 104.615
R330 VTAIL.n310 VTAIL.n233 104.615
R331 VTAIL.n310 VTAIL.n309 104.615
R332 VTAIL.n309 VTAIL.n237 104.615
R333 VTAIL.n302 VTAIL.n237 104.615
R334 VTAIL.n302 VTAIL.n301 104.615
R335 VTAIL.n301 VTAIL.n241 104.615
R336 VTAIL.n294 VTAIL.n241 104.615
R337 VTAIL.n294 VTAIL.n293 104.615
R338 VTAIL.n293 VTAIL.n245 104.615
R339 VTAIL.n286 VTAIL.n245 104.615
R340 VTAIL.n286 VTAIL.n285 104.615
R341 VTAIL.n285 VTAIL.n249 104.615
R342 VTAIL.n253 VTAIL.n249 104.615
R343 VTAIL.n277 VTAIL.n253 104.615
R344 VTAIL.n277 VTAIL.n276 104.615
R345 VTAIL.n276 VTAIL.n254 104.615
R346 VTAIL.n269 VTAIL.n254 104.615
R347 VTAIL.n269 VTAIL.n268 104.615
R348 VTAIL.n268 VTAIL.n258 104.615
R349 VTAIL.n261 VTAIL.n258 104.615
R350 VTAIL.n216 VTAIL.n215 104.615
R351 VTAIL.n215 VTAIL.n119 104.615
R352 VTAIL.n208 VTAIL.n119 104.615
R353 VTAIL.n208 VTAIL.n207 104.615
R354 VTAIL.n207 VTAIL.n123 104.615
R355 VTAIL.n200 VTAIL.n123 104.615
R356 VTAIL.n200 VTAIL.n199 104.615
R357 VTAIL.n199 VTAIL.n127 104.615
R358 VTAIL.n192 VTAIL.n127 104.615
R359 VTAIL.n192 VTAIL.n191 104.615
R360 VTAIL.n191 VTAIL.n131 104.615
R361 VTAIL.n184 VTAIL.n131 104.615
R362 VTAIL.n184 VTAIL.n183 104.615
R363 VTAIL.n183 VTAIL.n135 104.615
R364 VTAIL.n176 VTAIL.n135 104.615
R365 VTAIL.n176 VTAIL.n175 104.615
R366 VTAIL.n175 VTAIL.n139 104.615
R367 VTAIL.n143 VTAIL.n139 104.615
R368 VTAIL.n167 VTAIL.n143 104.615
R369 VTAIL.n167 VTAIL.n166 104.615
R370 VTAIL.n166 VTAIL.n144 104.615
R371 VTAIL.n159 VTAIL.n144 104.615
R372 VTAIL.n159 VTAIL.n158 104.615
R373 VTAIL.n158 VTAIL.n148 104.615
R374 VTAIL.n151 VTAIL.n148 104.615
R375 VTAIL.n366 VTAIL.t1 52.3082
R376 VTAIL.n36 VTAIL.t18 52.3082
R377 VTAIL.n261 VTAIL.t14 52.3082
R378 VTAIL.n151 VTAIL.t5 52.3082
R379 VTAIL.n225 VTAIL.n224 47.0139
R380 VTAIL.n223 VTAIL.n222 47.0139
R381 VTAIL.n115 VTAIL.n114 47.0139
R382 VTAIL.n113 VTAIL.n112 47.0139
R383 VTAIL.n439 VTAIL.n438 47.0138
R384 VTAIL.n1 VTAIL.n0 47.0138
R385 VTAIL.n109 VTAIL.n108 47.0138
R386 VTAIL.n111 VTAIL.n110 47.0138
R387 VTAIL.n437 VTAIL.n436 35.6763
R388 VTAIL.n107 VTAIL.n106 35.6763
R389 VTAIL.n331 VTAIL.n330 35.6763
R390 VTAIL.n221 VTAIL.n220 35.6763
R391 VTAIL.n113 VTAIL.n111 34.9703
R392 VTAIL.n437 VTAIL.n331 32.0738
R393 VTAIL.n390 VTAIL.n389 13.1884
R394 VTAIL.n60 VTAIL.n59 13.1884
R395 VTAIL.n284 VTAIL.n283 13.1884
R396 VTAIL.n174 VTAIL.n173 13.1884
R397 VTAIL.n388 VTAIL.n356 12.8005
R398 VTAIL.n393 VTAIL.n354 12.8005
R399 VTAIL.n434 VTAIL.n433 12.8005
R400 VTAIL.n58 VTAIL.n26 12.8005
R401 VTAIL.n63 VTAIL.n24 12.8005
R402 VTAIL.n104 VTAIL.n103 12.8005
R403 VTAIL.n328 VTAIL.n327 12.8005
R404 VTAIL.n287 VTAIL.n248 12.8005
R405 VTAIL.n282 VTAIL.n250 12.8005
R406 VTAIL.n218 VTAIL.n217 12.8005
R407 VTAIL.n177 VTAIL.n138 12.8005
R408 VTAIL.n172 VTAIL.n140 12.8005
R409 VTAIL.n385 VTAIL.n384 12.0247
R410 VTAIL.n394 VTAIL.n352 12.0247
R411 VTAIL.n430 VTAIL.n334 12.0247
R412 VTAIL.n55 VTAIL.n54 12.0247
R413 VTAIL.n64 VTAIL.n22 12.0247
R414 VTAIL.n100 VTAIL.n4 12.0247
R415 VTAIL.n324 VTAIL.n228 12.0247
R416 VTAIL.n288 VTAIL.n246 12.0247
R417 VTAIL.n279 VTAIL.n278 12.0247
R418 VTAIL.n214 VTAIL.n118 12.0247
R419 VTAIL.n178 VTAIL.n136 12.0247
R420 VTAIL.n169 VTAIL.n168 12.0247
R421 VTAIL.n380 VTAIL.n358 11.249
R422 VTAIL.n398 VTAIL.n397 11.249
R423 VTAIL.n429 VTAIL.n336 11.249
R424 VTAIL.n50 VTAIL.n28 11.249
R425 VTAIL.n68 VTAIL.n67 11.249
R426 VTAIL.n99 VTAIL.n6 11.249
R427 VTAIL.n323 VTAIL.n230 11.249
R428 VTAIL.n292 VTAIL.n291 11.249
R429 VTAIL.n275 VTAIL.n252 11.249
R430 VTAIL.n213 VTAIL.n120 11.249
R431 VTAIL.n182 VTAIL.n181 11.249
R432 VTAIL.n165 VTAIL.n142 11.249
R433 VTAIL.n379 VTAIL.n360 10.4732
R434 VTAIL.n401 VTAIL.n350 10.4732
R435 VTAIL.n426 VTAIL.n425 10.4732
R436 VTAIL.n49 VTAIL.n30 10.4732
R437 VTAIL.n71 VTAIL.n20 10.4732
R438 VTAIL.n96 VTAIL.n95 10.4732
R439 VTAIL.n320 VTAIL.n319 10.4732
R440 VTAIL.n295 VTAIL.n244 10.4732
R441 VTAIL.n274 VTAIL.n255 10.4732
R442 VTAIL.n210 VTAIL.n209 10.4732
R443 VTAIL.n185 VTAIL.n134 10.4732
R444 VTAIL.n164 VTAIL.n145 10.4732
R445 VTAIL.n367 VTAIL.n365 10.2747
R446 VTAIL.n37 VTAIL.n35 10.2747
R447 VTAIL.n262 VTAIL.n260 10.2747
R448 VTAIL.n152 VTAIL.n150 10.2747
R449 VTAIL.n376 VTAIL.n375 9.69747
R450 VTAIL.n402 VTAIL.n348 9.69747
R451 VTAIL.n422 VTAIL.n338 9.69747
R452 VTAIL.n46 VTAIL.n45 9.69747
R453 VTAIL.n72 VTAIL.n18 9.69747
R454 VTAIL.n92 VTAIL.n8 9.69747
R455 VTAIL.n316 VTAIL.n232 9.69747
R456 VTAIL.n296 VTAIL.n242 9.69747
R457 VTAIL.n271 VTAIL.n270 9.69747
R458 VTAIL.n206 VTAIL.n122 9.69747
R459 VTAIL.n186 VTAIL.n132 9.69747
R460 VTAIL.n161 VTAIL.n160 9.69747
R461 VTAIL.n436 VTAIL.n435 9.45567
R462 VTAIL.n106 VTAIL.n105 9.45567
R463 VTAIL.n330 VTAIL.n329 9.45567
R464 VTAIL.n220 VTAIL.n219 9.45567
R465 VTAIL.n411 VTAIL.n410 9.3005
R466 VTAIL.n346 VTAIL.n345 9.3005
R467 VTAIL.n405 VTAIL.n404 9.3005
R468 VTAIL.n403 VTAIL.n402 9.3005
R469 VTAIL.n350 VTAIL.n349 9.3005
R470 VTAIL.n397 VTAIL.n396 9.3005
R471 VTAIL.n395 VTAIL.n394 9.3005
R472 VTAIL.n354 VTAIL.n353 9.3005
R473 VTAIL.n369 VTAIL.n368 9.3005
R474 VTAIL.n371 VTAIL.n370 9.3005
R475 VTAIL.n362 VTAIL.n361 9.3005
R476 VTAIL.n377 VTAIL.n376 9.3005
R477 VTAIL.n379 VTAIL.n378 9.3005
R478 VTAIL.n358 VTAIL.n357 9.3005
R479 VTAIL.n386 VTAIL.n385 9.3005
R480 VTAIL.n388 VTAIL.n387 9.3005
R481 VTAIL.n413 VTAIL.n412 9.3005
R482 VTAIL.n342 VTAIL.n341 9.3005
R483 VTAIL.n419 VTAIL.n418 9.3005
R484 VTAIL.n421 VTAIL.n420 9.3005
R485 VTAIL.n338 VTAIL.n337 9.3005
R486 VTAIL.n427 VTAIL.n426 9.3005
R487 VTAIL.n429 VTAIL.n428 9.3005
R488 VTAIL.n334 VTAIL.n333 9.3005
R489 VTAIL.n435 VTAIL.n434 9.3005
R490 VTAIL.n81 VTAIL.n80 9.3005
R491 VTAIL.n16 VTAIL.n15 9.3005
R492 VTAIL.n75 VTAIL.n74 9.3005
R493 VTAIL.n73 VTAIL.n72 9.3005
R494 VTAIL.n20 VTAIL.n19 9.3005
R495 VTAIL.n67 VTAIL.n66 9.3005
R496 VTAIL.n65 VTAIL.n64 9.3005
R497 VTAIL.n24 VTAIL.n23 9.3005
R498 VTAIL.n39 VTAIL.n38 9.3005
R499 VTAIL.n41 VTAIL.n40 9.3005
R500 VTAIL.n32 VTAIL.n31 9.3005
R501 VTAIL.n47 VTAIL.n46 9.3005
R502 VTAIL.n49 VTAIL.n48 9.3005
R503 VTAIL.n28 VTAIL.n27 9.3005
R504 VTAIL.n56 VTAIL.n55 9.3005
R505 VTAIL.n58 VTAIL.n57 9.3005
R506 VTAIL.n83 VTAIL.n82 9.3005
R507 VTAIL.n12 VTAIL.n11 9.3005
R508 VTAIL.n89 VTAIL.n88 9.3005
R509 VTAIL.n91 VTAIL.n90 9.3005
R510 VTAIL.n8 VTAIL.n7 9.3005
R511 VTAIL.n97 VTAIL.n96 9.3005
R512 VTAIL.n99 VTAIL.n98 9.3005
R513 VTAIL.n4 VTAIL.n3 9.3005
R514 VTAIL.n105 VTAIL.n104 9.3005
R515 VTAIL.n264 VTAIL.n263 9.3005
R516 VTAIL.n266 VTAIL.n265 9.3005
R517 VTAIL.n257 VTAIL.n256 9.3005
R518 VTAIL.n272 VTAIL.n271 9.3005
R519 VTAIL.n274 VTAIL.n273 9.3005
R520 VTAIL.n252 VTAIL.n251 9.3005
R521 VTAIL.n280 VTAIL.n279 9.3005
R522 VTAIL.n282 VTAIL.n281 9.3005
R523 VTAIL.n236 VTAIL.n235 9.3005
R524 VTAIL.n313 VTAIL.n312 9.3005
R525 VTAIL.n315 VTAIL.n314 9.3005
R526 VTAIL.n232 VTAIL.n231 9.3005
R527 VTAIL.n321 VTAIL.n320 9.3005
R528 VTAIL.n323 VTAIL.n322 9.3005
R529 VTAIL.n228 VTAIL.n227 9.3005
R530 VTAIL.n329 VTAIL.n328 9.3005
R531 VTAIL.n307 VTAIL.n306 9.3005
R532 VTAIL.n305 VTAIL.n304 9.3005
R533 VTAIL.n240 VTAIL.n239 9.3005
R534 VTAIL.n299 VTAIL.n298 9.3005
R535 VTAIL.n297 VTAIL.n296 9.3005
R536 VTAIL.n244 VTAIL.n243 9.3005
R537 VTAIL.n291 VTAIL.n290 9.3005
R538 VTAIL.n289 VTAIL.n288 9.3005
R539 VTAIL.n248 VTAIL.n247 9.3005
R540 VTAIL.n154 VTAIL.n153 9.3005
R541 VTAIL.n156 VTAIL.n155 9.3005
R542 VTAIL.n147 VTAIL.n146 9.3005
R543 VTAIL.n162 VTAIL.n161 9.3005
R544 VTAIL.n164 VTAIL.n163 9.3005
R545 VTAIL.n142 VTAIL.n141 9.3005
R546 VTAIL.n170 VTAIL.n169 9.3005
R547 VTAIL.n172 VTAIL.n171 9.3005
R548 VTAIL.n126 VTAIL.n125 9.3005
R549 VTAIL.n203 VTAIL.n202 9.3005
R550 VTAIL.n205 VTAIL.n204 9.3005
R551 VTAIL.n122 VTAIL.n121 9.3005
R552 VTAIL.n211 VTAIL.n210 9.3005
R553 VTAIL.n213 VTAIL.n212 9.3005
R554 VTAIL.n118 VTAIL.n117 9.3005
R555 VTAIL.n219 VTAIL.n218 9.3005
R556 VTAIL.n197 VTAIL.n196 9.3005
R557 VTAIL.n195 VTAIL.n194 9.3005
R558 VTAIL.n130 VTAIL.n129 9.3005
R559 VTAIL.n189 VTAIL.n188 9.3005
R560 VTAIL.n187 VTAIL.n186 9.3005
R561 VTAIL.n134 VTAIL.n133 9.3005
R562 VTAIL.n181 VTAIL.n180 9.3005
R563 VTAIL.n179 VTAIL.n178 9.3005
R564 VTAIL.n138 VTAIL.n137 9.3005
R565 VTAIL.n372 VTAIL.n362 8.92171
R566 VTAIL.n406 VTAIL.n405 8.92171
R567 VTAIL.n421 VTAIL.n340 8.92171
R568 VTAIL.n42 VTAIL.n32 8.92171
R569 VTAIL.n76 VTAIL.n75 8.92171
R570 VTAIL.n91 VTAIL.n10 8.92171
R571 VTAIL.n315 VTAIL.n234 8.92171
R572 VTAIL.n300 VTAIL.n299 8.92171
R573 VTAIL.n267 VTAIL.n257 8.92171
R574 VTAIL.n205 VTAIL.n124 8.92171
R575 VTAIL.n190 VTAIL.n189 8.92171
R576 VTAIL.n157 VTAIL.n147 8.92171
R577 VTAIL.n436 VTAIL.n332 8.2187
R578 VTAIL.n106 VTAIL.n2 8.2187
R579 VTAIL.n330 VTAIL.n226 8.2187
R580 VTAIL.n220 VTAIL.n116 8.2187
R581 VTAIL.n371 VTAIL.n364 8.14595
R582 VTAIL.n409 VTAIL.n346 8.14595
R583 VTAIL.n418 VTAIL.n417 8.14595
R584 VTAIL.n41 VTAIL.n34 8.14595
R585 VTAIL.n79 VTAIL.n16 8.14595
R586 VTAIL.n88 VTAIL.n87 8.14595
R587 VTAIL.n312 VTAIL.n311 8.14595
R588 VTAIL.n303 VTAIL.n240 8.14595
R589 VTAIL.n266 VTAIL.n259 8.14595
R590 VTAIL.n202 VTAIL.n201 8.14595
R591 VTAIL.n193 VTAIL.n130 8.14595
R592 VTAIL.n156 VTAIL.n149 8.14595
R593 VTAIL.n368 VTAIL.n367 7.3702
R594 VTAIL.n410 VTAIL.n344 7.3702
R595 VTAIL.n414 VTAIL.n342 7.3702
R596 VTAIL.n38 VTAIL.n37 7.3702
R597 VTAIL.n80 VTAIL.n14 7.3702
R598 VTAIL.n84 VTAIL.n12 7.3702
R599 VTAIL.n308 VTAIL.n236 7.3702
R600 VTAIL.n304 VTAIL.n238 7.3702
R601 VTAIL.n263 VTAIL.n262 7.3702
R602 VTAIL.n198 VTAIL.n126 7.3702
R603 VTAIL.n194 VTAIL.n128 7.3702
R604 VTAIL.n153 VTAIL.n152 7.3702
R605 VTAIL.n413 VTAIL.n344 6.59444
R606 VTAIL.n414 VTAIL.n413 6.59444
R607 VTAIL.n83 VTAIL.n14 6.59444
R608 VTAIL.n84 VTAIL.n83 6.59444
R609 VTAIL.n308 VTAIL.n307 6.59444
R610 VTAIL.n307 VTAIL.n238 6.59444
R611 VTAIL.n198 VTAIL.n197 6.59444
R612 VTAIL.n197 VTAIL.n128 6.59444
R613 VTAIL.n368 VTAIL.n364 5.81868
R614 VTAIL.n410 VTAIL.n409 5.81868
R615 VTAIL.n417 VTAIL.n342 5.81868
R616 VTAIL.n38 VTAIL.n34 5.81868
R617 VTAIL.n80 VTAIL.n79 5.81868
R618 VTAIL.n87 VTAIL.n12 5.81868
R619 VTAIL.n311 VTAIL.n236 5.81868
R620 VTAIL.n304 VTAIL.n303 5.81868
R621 VTAIL.n263 VTAIL.n259 5.81868
R622 VTAIL.n201 VTAIL.n126 5.81868
R623 VTAIL.n194 VTAIL.n193 5.81868
R624 VTAIL.n153 VTAIL.n149 5.81868
R625 VTAIL.n434 VTAIL.n332 5.3904
R626 VTAIL.n104 VTAIL.n2 5.3904
R627 VTAIL.n328 VTAIL.n226 5.3904
R628 VTAIL.n218 VTAIL.n116 5.3904
R629 VTAIL.n372 VTAIL.n371 5.04292
R630 VTAIL.n406 VTAIL.n346 5.04292
R631 VTAIL.n418 VTAIL.n340 5.04292
R632 VTAIL.n42 VTAIL.n41 5.04292
R633 VTAIL.n76 VTAIL.n16 5.04292
R634 VTAIL.n88 VTAIL.n10 5.04292
R635 VTAIL.n312 VTAIL.n234 5.04292
R636 VTAIL.n300 VTAIL.n240 5.04292
R637 VTAIL.n267 VTAIL.n266 5.04292
R638 VTAIL.n202 VTAIL.n124 5.04292
R639 VTAIL.n190 VTAIL.n130 5.04292
R640 VTAIL.n157 VTAIL.n156 5.04292
R641 VTAIL.n375 VTAIL.n362 4.26717
R642 VTAIL.n405 VTAIL.n348 4.26717
R643 VTAIL.n422 VTAIL.n421 4.26717
R644 VTAIL.n45 VTAIL.n32 4.26717
R645 VTAIL.n75 VTAIL.n18 4.26717
R646 VTAIL.n92 VTAIL.n91 4.26717
R647 VTAIL.n316 VTAIL.n315 4.26717
R648 VTAIL.n299 VTAIL.n242 4.26717
R649 VTAIL.n270 VTAIL.n257 4.26717
R650 VTAIL.n206 VTAIL.n205 4.26717
R651 VTAIL.n189 VTAIL.n132 4.26717
R652 VTAIL.n160 VTAIL.n147 4.26717
R653 VTAIL.n376 VTAIL.n360 3.49141
R654 VTAIL.n402 VTAIL.n401 3.49141
R655 VTAIL.n425 VTAIL.n338 3.49141
R656 VTAIL.n46 VTAIL.n30 3.49141
R657 VTAIL.n72 VTAIL.n71 3.49141
R658 VTAIL.n95 VTAIL.n8 3.49141
R659 VTAIL.n319 VTAIL.n232 3.49141
R660 VTAIL.n296 VTAIL.n295 3.49141
R661 VTAIL.n271 VTAIL.n255 3.49141
R662 VTAIL.n209 VTAIL.n122 3.49141
R663 VTAIL.n186 VTAIL.n185 3.49141
R664 VTAIL.n161 VTAIL.n145 3.49141
R665 VTAIL.n115 VTAIL.n113 2.89705
R666 VTAIL.n221 VTAIL.n115 2.89705
R667 VTAIL.n225 VTAIL.n223 2.89705
R668 VTAIL.n331 VTAIL.n225 2.89705
R669 VTAIL.n111 VTAIL.n109 2.89705
R670 VTAIL.n109 VTAIL.n107 2.89705
R671 VTAIL.n439 VTAIL.n437 2.89705
R672 VTAIL.n369 VTAIL.n365 2.84303
R673 VTAIL.n39 VTAIL.n35 2.84303
R674 VTAIL.n264 VTAIL.n260 2.84303
R675 VTAIL.n154 VTAIL.n150 2.84303
R676 VTAIL.n380 VTAIL.n379 2.71565
R677 VTAIL.n398 VTAIL.n350 2.71565
R678 VTAIL.n426 VTAIL.n336 2.71565
R679 VTAIL.n50 VTAIL.n49 2.71565
R680 VTAIL.n68 VTAIL.n20 2.71565
R681 VTAIL.n96 VTAIL.n6 2.71565
R682 VTAIL.n320 VTAIL.n230 2.71565
R683 VTAIL.n292 VTAIL.n244 2.71565
R684 VTAIL.n275 VTAIL.n274 2.71565
R685 VTAIL.n210 VTAIL.n120 2.71565
R686 VTAIL.n182 VTAIL.n134 2.71565
R687 VTAIL.n165 VTAIL.n164 2.71565
R688 VTAIL VTAIL.n1 2.2311
R689 VTAIL.n384 VTAIL.n358 1.93989
R690 VTAIL.n397 VTAIL.n352 1.93989
R691 VTAIL.n430 VTAIL.n429 1.93989
R692 VTAIL.n54 VTAIL.n28 1.93989
R693 VTAIL.n67 VTAIL.n22 1.93989
R694 VTAIL.n100 VTAIL.n99 1.93989
R695 VTAIL.n324 VTAIL.n323 1.93989
R696 VTAIL.n291 VTAIL.n246 1.93989
R697 VTAIL.n278 VTAIL.n252 1.93989
R698 VTAIL.n214 VTAIL.n213 1.93989
R699 VTAIL.n181 VTAIL.n136 1.93989
R700 VTAIL.n168 VTAIL.n142 1.93989
R701 VTAIL.n223 VTAIL.n221 1.9186
R702 VTAIL.n107 VTAIL.n1 1.9186
R703 VTAIL.n385 VTAIL.n356 1.16414
R704 VTAIL.n394 VTAIL.n393 1.16414
R705 VTAIL.n433 VTAIL.n334 1.16414
R706 VTAIL.n55 VTAIL.n26 1.16414
R707 VTAIL.n64 VTAIL.n63 1.16414
R708 VTAIL.n103 VTAIL.n4 1.16414
R709 VTAIL.n327 VTAIL.n228 1.16414
R710 VTAIL.n288 VTAIL.n287 1.16414
R711 VTAIL.n279 VTAIL.n250 1.16414
R712 VTAIL.n217 VTAIL.n118 1.16414
R713 VTAIL.n178 VTAIL.n177 1.16414
R714 VTAIL.n169 VTAIL.n140 1.16414
R715 VTAIL.n438 VTAIL.t9 1.01588
R716 VTAIL.n438 VTAIL.t3 1.01588
R717 VTAIL.n0 VTAIL.t7 1.01588
R718 VTAIL.n0 VTAIL.t4 1.01588
R719 VTAIL.n108 VTAIL.t16 1.01588
R720 VTAIL.n108 VTAIL.t13 1.01588
R721 VTAIL.n110 VTAIL.t15 1.01588
R722 VTAIL.n110 VTAIL.t19 1.01588
R723 VTAIL.n224 VTAIL.t11 1.01588
R724 VTAIL.n224 VTAIL.t17 1.01588
R725 VTAIL.n222 VTAIL.t12 1.01588
R726 VTAIL.n222 VTAIL.t10 1.01588
R727 VTAIL.n114 VTAIL.t6 1.01588
R728 VTAIL.n114 VTAIL.t0 1.01588
R729 VTAIL.n112 VTAIL.t2 1.01588
R730 VTAIL.n112 VTAIL.t8 1.01588
R731 VTAIL VTAIL.n439 0.666448
R732 VTAIL.n389 VTAIL.n388 0.388379
R733 VTAIL.n390 VTAIL.n354 0.388379
R734 VTAIL.n59 VTAIL.n58 0.388379
R735 VTAIL.n60 VTAIL.n24 0.388379
R736 VTAIL.n284 VTAIL.n248 0.388379
R737 VTAIL.n283 VTAIL.n282 0.388379
R738 VTAIL.n174 VTAIL.n138 0.388379
R739 VTAIL.n173 VTAIL.n172 0.388379
R740 VTAIL.n370 VTAIL.n369 0.155672
R741 VTAIL.n370 VTAIL.n361 0.155672
R742 VTAIL.n377 VTAIL.n361 0.155672
R743 VTAIL.n378 VTAIL.n377 0.155672
R744 VTAIL.n378 VTAIL.n357 0.155672
R745 VTAIL.n386 VTAIL.n357 0.155672
R746 VTAIL.n387 VTAIL.n386 0.155672
R747 VTAIL.n387 VTAIL.n353 0.155672
R748 VTAIL.n395 VTAIL.n353 0.155672
R749 VTAIL.n396 VTAIL.n395 0.155672
R750 VTAIL.n396 VTAIL.n349 0.155672
R751 VTAIL.n403 VTAIL.n349 0.155672
R752 VTAIL.n404 VTAIL.n403 0.155672
R753 VTAIL.n404 VTAIL.n345 0.155672
R754 VTAIL.n411 VTAIL.n345 0.155672
R755 VTAIL.n412 VTAIL.n411 0.155672
R756 VTAIL.n412 VTAIL.n341 0.155672
R757 VTAIL.n419 VTAIL.n341 0.155672
R758 VTAIL.n420 VTAIL.n419 0.155672
R759 VTAIL.n420 VTAIL.n337 0.155672
R760 VTAIL.n427 VTAIL.n337 0.155672
R761 VTAIL.n428 VTAIL.n427 0.155672
R762 VTAIL.n428 VTAIL.n333 0.155672
R763 VTAIL.n435 VTAIL.n333 0.155672
R764 VTAIL.n40 VTAIL.n39 0.155672
R765 VTAIL.n40 VTAIL.n31 0.155672
R766 VTAIL.n47 VTAIL.n31 0.155672
R767 VTAIL.n48 VTAIL.n47 0.155672
R768 VTAIL.n48 VTAIL.n27 0.155672
R769 VTAIL.n56 VTAIL.n27 0.155672
R770 VTAIL.n57 VTAIL.n56 0.155672
R771 VTAIL.n57 VTAIL.n23 0.155672
R772 VTAIL.n65 VTAIL.n23 0.155672
R773 VTAIL.n66 VTAIL.n65 0.155672
R774 VTAIL.n66 VTAIL.n19 0.155672
R775 VTAIL.n73 VTAIL.n19 0.155672
R776 VTAIL.n74 VTAIL.n73 0.155672
R777 VTAIL.n74 VTAIL.n15 0.155672
R778 VTAIL.n81 VTAIL.n15 0.155672
R779 VTAIL.n82 VTAIL.n81 0.155672
R780 VTAIL.n82 VTAIL.n11 0.155672
R781 VTAIL.n89 VTAIL.n11 0.155672
R782 VTAIL.n90 VTAIL.n89 0.155672
R783 VTAIL.n90 VTAIL.n7 0.155672
R784 VTAIL.n97 VTAIL.n7 0.155672
R785 VTAIL.n98 VTAIL.n97 0.155672
R786 VTAIL.n98 VTAIL.n3 0.155672
R787 VTAIL.n105 VTAIL.n3 0.155672
R788 VTAIL.n329 VTAIL.n227 0.155672
R789 VTAIL.n322 VTAIL.n227 0.155672
R790 VTAIL.n322 VTAIL.n321 0.155672
R791 VTAIL.n321 VTAIL.n231 0.155672
R792 VTAIL.n314 VTAIL.n231 0.155672
R793 VTAIL.n314 VTAIL.n313 0.155672
R794 VTAIL.n313 VTAIL.n235 0.155672
R795 VTAIL.n306 VTAIL.n235 0.155672
R796 VTAIL.n306 VTAIL.n305 0.155672
R797 VTAIL.n305 VTAIL.n239 0.155672
R798 VTAIL.n298 VTAIL.n239 0.155672
R799 VTAIL.n298 VTAIL.n297 0.155672
R800 VTAIL.n297 VTAIL.n243 0.155672
R801 VTAIL.n290 VTAIL.n243 0.155672
R802 VTAIL.n290 VTAIL.n289 0.155672
R803 VTAIL.n289 VTAIL.n247 0.155672
R804 VTAIL.n281 VTAIL.n247 0.155672
R805 VTAIL.n281 VTAIL.n280 0.155672
R806 VTAIL.n280 VTAIL.n251 0.155672
R807 VTAIL.n273 VTAIL.n251 0.155672
R808 VTAIL.n273 VTAIL.n272 0.155672
R809 VTAIL.n272 VTAIL.n256 0.155672
R810 VTAIL.n265 VTAIL.n256 0.155672
R811 VTAIL.n265 VTAIL.n264 0.155672
R812 VTAIL.n219 VTAIL.n117 0.155672
R813 VTAIL.n212 VTAIL.n117 0.155672
R814 VTAIL.n212 VTAIL.n211 0.155672
R815 VTAIL.n211 VTAIL.n121 0.155672
R816 VTAIL.n204 VTAIL.n121 0.155672
R817 VTAIL.n204 VTAIL.n203 0.155672
R818 VTAIL.n203 VTAIL.n125 0.155672
R819 VTAIL.n196 VTAIL.n125 0.155672
R820 VTAIL.n196 VTAIL.n195 0.155672
R821 VTAIL.n195 VTAIL.n129 0.155672
R822 VTAIL.n188 VTAIL.n129 0.155672
R823 VTAIL.n188 VTAIL.n187 0.155672
R824 VTAIL.n187 VTAIL.n133 0.155672
R825 VTAIL.n180 VTAIL.n133 0.155672
R826 VTAIL.n180 VTAIL.n179 0.155672
R827 VTAIL.n179 VTAIL.n137 0.155672
R828 VTAIL.n171 VTAIL.n137 0.155672
R829 VTAIL.n171 VTAIL.n170 0.155672
R830 VTAIL.n170 VTAIL.n141 0.155672
R831 VTAIL.n163 VTAIL.n141 0.155672
R832 VTAIL.n163 VTAIL.n162 0.155672
R833 VTAIL.n162 VTAIL.n146 0.155672
R834 VTAIL.n155 VTAIL.n146 0.155672
R835 VTAIL.n155 VTAIL.n154 0.155672
R836 VDD1.n100 VDD1.n0 214.453
R837 VDD1.n207 VDD1.n107 214.453
R838 VDD1.n101 VDD1.n100 185
R839 VDD1.n99 VDD1.n98 185
R840 VDD1.n4 VDD1.n3 185
R841 VDD1.n93 VDD1.n92 185
R842 VDD1.n91 VDD1.n90 185
R843 VDD1.n8 VDD1.n7 185
R844 VDD1.n85 VDD1.n84 185
R845 VDD1.n83 VDD1.n82 185
R846 VDD1.n12 VDD1.n11 185
R847 VDD1.n77 VDD1.n76 185
R848 VDD1.n75 VDD1.n74 185
R849 VDD1.n16 VDD1.n15 185
R850 VDD1.n69 VDD1.n68 185
R851 VDD1.n67 VDD1.n66 185
R852 VDD1.n20 VDD1.n19 185
R853 VDD1.n61 VDD1.n60 185
R854 VDD1.n59 VDD1.n58 185
R855 VDD1.n57 VDD1.n23 185
R856 VDD1.n27 VDD1.n24 185
R857 VDD1.n52 VDD1.n51 185
R858 VDD1.n50 VDD1.n49 185
R859 VDD1.n29 VDD1.n28 185
R860 VDD1.n44 VDD1.n43 185
R861 VDD1.n42 VDD1.n41 185
R862 VDD1.n33 VDD1.n32 185
R863 VDD1.n36 VDD1.n35 185
R864 VDD1.n142 VDD1.n141 185
R865 VDD1.n139 VDD1.n138 185
R866 VDD1.n148 VDD1.n147 185
R867 VDD1.n150 VDD1.n149 185
R868 VDD1.n135 VDD1.n134 185
R869 VDD1.n156 VDD1.n155 185
R870 VDD1.n159 VDD1.n158 185
R871 VDD1.n157 VDD1.n131 185
R872 VDD1.n164 VDD1.n130 185
R873 VDD1.n166 VDD1.n165 185
R874 VDD1.n168 VDD1.n167 185
R875 VDD1.n127 VDD1.n126 185
R876 VDD1.n174 VDD1.n173 185
R877 VDD1.n176 VDD1.n175 185
R878 VDD1.n123 VDD1.n122 185
R879 VDD1.n182 VDD1.n181 185
R880 VDD1.n184 VDD1.n183 185
R881 VDD1.n119 VDD1.n118 185
R882 VDD1.n190 VDD1.n189 185
R883 VDD1.n192 VDD1.n191 185
R884 VDD1.n115 VDD1.n114 185
R885 VDD1.n198 VDD1.n197 185
R886 VDD1.n200 VDD1.n199 185
R887 VDD1.n111 VDD1.n110 185
R888 VDD1.n206 VDD1.n205 185
R889 VDD1.n208 VDD1.n207 185
R890 VDD1.t2 VDD1.n34 149.524
R891 VDD1.t4 VDD1.n140 149.524
R892 VDD1.n100 VDD1.n99 104.615
R893 VDD1.n99 VDD1.n3 104.615
R894 VDD1.n92 VDD1.n3 104.615
R895 VDD1.n92 VDD1.n91 104.615
R896 VDD1.n91 VDD1.n7 104.615
R897 VDD1.n84 VDD1.n7 104.615
R898 VDD1.n84 VDD1.n83 104.615
R899 VDD1.n83 VDD1.n11 104.615
R900 VDD1.n76 VDD1.n11 104.615
R901 VDD1.n76 VDD1.n75 104.615
R902 VDD1.n75 VDD1.n15 104.615
R903 VDD1.n68 VDD1.n15 104.615
R904 VDD1.n68 VDD1.n67 104.615
R905 VDD1.n67 VDD1.n19 104.615
R906 VDD1.n60 VDD1.n19 104.615
R907 VDD1.n60 VDD1.n59 104.615
R908 VDD1.n59 VDD1.n23 104.615
R909 VDD1.n27 VDD1.n23 104.615
R910 VDD1.n51 VDD1.n27 104.615
R911 VDD1.n51 VDD1.n50 104.615
R912 VDD1.n50 VDD1.n28 104.615
R913 VDD1.n43 VDD1.n28 104.615
R914 VDD1.n43 VDD1.n42 104.615
R915 VDD1.n42 VDD1.n32 104.615
R916 VDD1.n35 VDD1.n32 104.615
R917 VDD1.n141 VDD1.n138 104.615
R918 VDD1.n148 VDD1.n138 104.615
R919 VDD1.n149 VDD1.n148 104.615
R920 VDD1.n149 VDD1.n134 104.615
R921 VDD1.n156 VDD1.n134 104.615
R922 VDD1.n158 VDD1.n156 104.615
R923 VDD1.n158 VDD1.n157 104.615
R924 VDD1.n157 VDD1.n130 104.615
R925 VDD1.n166 VDD1.n130 104.615
R926 VDD1.n167 VDD1.n166 104.615
R927 VDD1.n167 VDD1.n126 104.615
R928 VDD1.n174 VDD1.n126 104.615
R929 VDD1.n175 VDD1.n174 104.615
R930 VDD1.n175 VDD1.n122 104.615
R931 VDD1.n182 VDD1.n122 104.615
R932 VDD1.n183 VDD1.n182 104.615
R933 VDD1.n183 VDD1.n118 104.615
R934 VDD1.n190 VDD1.n118 104.615
R935 VDD1.n191 VDD1.n190 104.615
R936 VDD1.n191 VDD1.n114 104.615
R937 VDD1.n198 VDD1.n114 104.615
R938 VDD1.n199 VDD1.n198 104.615
R939 VDD1.n199 VDD1.n110 104.615
R940 VDD1.n206 VDD1.n110 104.615
R941 VDD1.n207 VDD1.n206 104.615
R942 VDD1.n215 VDD1.n214 65.8096
R943 VDD1.n106 VDD1.n105 63.6927
R944 VDD1.n217 VDD1.n216 63.6925
R945 VDD1.n213 VDD1.n212 63.6925
R946 VDD1.n217 VDD1.n215 56.3155
R947 VDD1.n106 VDD1.n104 55.2516
R948 VDD1.n213 VDD1.n211 55.2516
R949 VDD1.n35 VDD1.t2 52.3082
R950 VDD1.n141 VDD1.t4 52.3082
R951 VDD1.n58 VDD1.n57 13.1884
R952 VDD1.n165 VDD1.n164 13.1884
R953 VDD1.n102 VDD1.n101 12.8005
R954 VDD1.n61 VDD1.n22 12.8005
R955 VDD1.n56 VDD1.n24 12.8005
R956 VDD1.n163 VDD1.n131 12.8005
R957 VDD1.n168 VDD1.n129 12.8005
R958 VDD1.n209 VDD1.n208 12.8005
R959 VDD1.n98 VDD1.n2 12.0247
R960 VDD1.n62 VDD1.n20 12.0247
R961 VDD1.n53 VDD1.n52 12.0247
R962 VDD1.n160 VDD1.n159 12.0247
R963 VDD1.n169 VDD1.n127 12.0247
R964 VDD1.n205 VDD1.n109 12.0247
R965 VDD1.n97 VDD1.n4 11.249
R966 VDD1.n66 VDD1.n65 11.249
R967 VDD1.n49 VDD1.n26 11.249
R968 VDD1.n155 VDD1.n133 11.249
R969 VDD1.n173 VDD1.n172 11.249
R970 VDD1.n204 VDD1.n111 11.249
R971 VDD1.n94 VDD1.n93 10.4732
R972 VDD1.n69 VDD1.n18 10.4732
R973 VDD1.n48 VDD1.n29 10.4732
R974 VDD1.n154 VDD1.n135 10.4732
R975 VDD1.n176 VDD1.n125 10.4732
R976 VDD1.n201 VDD1.n200 10.4732
R977 VDD1.n36 VDD1.n34 10.2747
R978 VDD1.n142 VDD1.n140 10.2747
R979 VDD1.n90 VDD1.n6 9.69747
R980 VDD1.n70 VDD1.n16 9.69747
R981 VDD1.n45 VDD1.n44 9.69747
R982 VDD1.n151 VDD1.n150 9.69747
R983 VDD1.n177 VDD1.n123 9.69747
R984 VDD1.n197 VDD1.n113 9.69747
R985 VDD1.n104 VDD1.n103 9.45567
R986 VDD1.n211 VDD1.n210 9.45567
R987 VDD1.n38 VDD1.n37 9.3005
R988 VDD1.n40 VDD1.n39 9.3005
R989 VDD1.n31 VDD1.n30 9.3005
R990 VDD1.n46 VDD1.n45 9.3005
R991 VDD1.n48 VDD1.n47 9.3005
R992 VDD1.n26 VDD1.n25 9.3005
R993 VDD1.n54 VDD1.n53 9.3005
R994 VDD1.n56 VDD1.n55 9.3005
R995 VDD1.n10 VDD1.n9 9.3005
R996 VDD1.n87 VDD1.n86 9.3005
R997 VDD1.n89 VDD1.n88 9.3005
R998 VDD1.n6 VDD1.n5 9.3005
R999 VDD1.n95 VDD1.n94 9.3005
R1000 VDD1.n97 VDD1.n96 9.3005
R1001 VDD1.n2 VDD1.n1 9.3005
R1002 VDD1.n103 VDD1.n102 9.3005
R1003 VDD1.n81 VDD1.n80 9.3005
R1004 VDD1.n79 VDD1.n78 9.3005
R1005 VDD1.n14 VDD1.n13 9.3005
R1006 VDD1.n73 VDD1.n72 9.3005
R1007 VDD1.n71 VDD1.n70 9.3005
R1008 VDD1.n18 VDD1.n17 9.3005
R1009 VDD1.n65 VDD1.n64 9.3005
R1010 VDD1.n63 VDD1.n62 9.3005
R1011 VDD1.n22 VDD1.n21 9.3005
R1012 VDD1.n186 VDD1.n185 9.3005
R1013 VDD1.n121 VDD1.n120 9.3005
R1014 VDD1.n180 VDD1.n179 9.3005
R1015 VDD1.n178 VDD1.n177 9.3005
R1016 VDD1.n125 VDD1.n124 9.3005
R1017 VDD1.n172 VDD1.n171 9.3005
R1018 VDD1.n170 VDD1.n169 9.3005
R1019 VDD1.n129 VDD1.n128 9.3005
R1020 VDD1.n144 VDD1.n143 9.3005
R1021 VDD1.n146 VDD1.n145 9.3005
R1022 VDD1.n137 VDD1.n136 9.3005
R1023 VDD1.n152 VDD1.n151 9.3005
R1024 VDD1.n154 VDD1.n153 9.3005
R1025 VDD1.n133 VDD1.n132 9.3005
R1026 VDD1.n161 VDD1.n160 9.3005
R1027 VDD1.n163 VDD1.n162 9.3005
R1028 VDD1.n188 VDD1.n187 9.3005
R1029 VDD1.n117 VDD1.n116 9.3005
R1030 VDD1.n194 VDD1.n193 9.3005
R1031 VDD1.n196 VDD1.n195 9.3005
R1032 VDD1.n113 VDD1.n112 9.3005
R1033 VDD1.n202 VDD1.n201 9.3005
R1034 VDD1.n204 VDD1.n203 9.3005
R1035 VDD1.n109 VDD1.n108 9.3005
R1036 VDD1.n210 VDD1.n209 9.3005
R1037 VDD1.n89 VDD1.n8 8.92171
R1038 VDD1.n74 VDD1.n73 8.92171
R1039 VDD1.n41 VDD1.n31 8.92171
R1040 VDD1.n147 VDD1.n137 8.92171
R1041 VDD1.n181 VDD1.n180 8.92171
R1042 VDD1.n196 VDD1.n115 8.92171
R1043 VDD1.n104 VDD1.n0 8.2187
R1044 VDD1.n211 VDD1.n107 8.2187
R1045 VDD1.n86 VDD1.n85 8.14595
R1046 VDD1.n77 VDD1.n14 8.14595
R1047 VDD1.n40 VDD1.n33 8.14595
R1048 VDD1.n146 VDD1.n139 8.14595
R1049 VDD1.n184 VDD1.n121 8.14595
R1050 VDD1.n193 VDD1.n192 8.14595
R1051 VDD1.n82 VDD1.n10 7.3702
R1052 VDD1.n78 VDD1.n12 7.3702
R1053 VDD1.n37 VDD1.n36 7.3702
R1054 VDD1.n143 VDD1.n142 7.3702
R1055 VDD1.n185 VDD1.n119 7.3702
R1056 VDD1.n189 VDD1.n117 7.3702
R1057 VDD1.n82 VDD1.n81 6.59444
R1058 VDD1.n81 VDD1.n12 6.59444
R1059 VDD1.n188 VDD1.n119 6.59444
R1060 VDD1.n189 VDD1.n188 6.59444
R1061 VDD1.n85 VDD1.n10 5.81868
R1062 VDD1.n78 VDD1.n77 5.81868
R1063 VDD1.n37 VDD1.n33 5.81868
R1064 VDD1.n143 VDD1.n139 5.81868
R1065 VDD1.n185 VDD1.n184 5.81868
R1066 VDD1.n192 VDD1.n117 5.81868
R1067 VDD1.n102 VDD1.n0 5.3904
R1068 VDD1.n209 VDD1.n107 5.3904
R1069 VDD1.n86 VDD1.n8 5.04292
R1070 VDD1.n74 VDD1.n14 5.04292
R1071 VDD1.n41 VDD1.n40 5.04292
R1072 VDD1.n147 VDD1.n146 5.04292
R1073 VDD1.n181 VDD1.n121 5.04292
R1074 VDD1.n193 VDD1.n115 5.04292
R1075 VDD1.n90 VDD1.n89 4.26717
R1076 VDD1.n73 VDD1.n16 4.26717
R1077 VDD1.n44 VDD1.n31 4.26717
R1078 VDD1.n150 VDD1.n137 4.26717
R1079 VDD1.n180 VDD1.n123 4.26717
R1080 VDD1.n197 VDD1.n196 4.26717
R1081 VDD1.n93 VDD1.n6 3.49141
R1082 VDD1.n70 VDD1.n69 3.49141
R1083 VDD1.n45 VDD1.n29 3.49141
R1084 VDD1.n151 VDD1.n135 3.49141
R1085 VDD1.n177 VDD1.n176 3.49141
R1086 VDD1.n200 VDD1.n113 3.49141
R1087 VDD1.n144 VDD1.n140 2.84303
R1088 VDD1.n38 VDD1.n34 2.84303
R1089 VDD1.n94 VDD1.n4 2.71565
R1090 VDD1.n66 VDD1.n18 2.71565
R1091 VDD1.n49 VDD1.n48 2.71565
R1092 VDD1.n155 VDD1.n154 2.71565
R1093 VDD1.n173 VDD1.n125 2.71565
R1094 VDD1.n201 VDD1.n111 2.71565
R1095 VDD1 VDD1.n217 2.11472
R1096 VDD1.n98 VDD1.n97 1.93989
R1097 VDD1.n65 VDD1.n20 1.93989
R1098 VDD1.n52 VDD1.n26 1.93989
R1099 VDD1.n159 VDD1.n133 1.93989
R1100 VDD1.n172 VDD1.n127 1.93989
R1101 VDD1.n205 VDD1.n204 1.93989
R1102 VDD1.n101 VDD1.n2 1.16414
R1103 VDD1.n62 VDD1.n61 1.16414
R1104 VDD1.n53 VDD1.n24 1.16414
R1105 VDD1.n160 VDD1.n131 1.16414
R1106 VDD1.n169 VDD1.n168 1.16414
R1107 VDD1.n208 VDD1.n109 1.16414
R1108 VDD1.n216 VDD1.t6 1.01588
R1109 VDD1.n216 VDD1.t9 1.01588
R1110 VDD1.n105 VDD1.t3 1.01588
R1111 VDD1.n105 VDD1.t7 1.01588
R1112 VDD1.n214 VDD1.t0 1.01588
R1113 VDD1.n214 VDD1.t5 1.01588
R1114 VDD1.n212 VDD1.t8 1.01588
R1115 VDD1.n212 VDD1.t1 1.01588
R1116 VDD1 VDD1.n106 0.782828
R1117 VDD1.n215 VDD1.n213 0.669292
R1118 VDD1.n58 VDD1.n22 0.388379
R1119 VDD1.n57 VDD1.n56 0.388379
R1120 VDD1.n164 VDD1.n163 0.388379
R1121 VDD1.n165 VDD1.n129 0.388379
R1122 VDD1.n103 VDD1.n1 0.155672
R1123 VDD1.n96 VDD1.n1 0.155672
R1124 VDD1.n96 VDD1.n95 0.155672
R1125 VDD1.n95 VDD1.n5 0.155672
R1126 VDD1.n88 VDD1.n5 0.155672
R1127 VDD1.n88 VDD1.n87 0.155672
R1128 VDD1.n87 VDD1.n9 0.155672
R1129 VDD1.n80 VDD1.n9 0.155672
R1130 VDD1.n80 VDD1.n79 0.155672
R1131 VDD1.n79 VDD1.n13 0.155672
R1132 VDD1.n72 VDD1.n13 0.155672
R1133 VDD1.n72 VDD1.n71 0.155672
R1134 VDD1.n71 VDD1.n17 0.155672
R1135 VDD1.n64 VDD1.n17 0.155672
R1136 VDD1.n64 VDD1.n63 0.155672
R1137 VDD1.n63 VDD1.n21 0.155672
R1138 VDD1.n55 VDD1.n21 0.155672
R1139 VDD1.n55 VDD1.n54 0.155672
R1140 VDD1.n54 VDD1.n25 0.155672
R1141 VDD1.n47 VDD1.n25 0.155672
R1142 VDD1.n47 VDD1.n46 0.155672
R1143 VDD1.n46 VDD1.n30 0.155672
R1144 VDD1.n39 VDD1.n30 0.155672
R1145 VDD1.n39 VDD1.n38 0.155672
R1146 VDD1.n145 VDD1.n144 0.155672
R1147 VDD1.n145 VDD1.n136 0.155672
R1148 VDD1.n152 VDD1.n136 0.155672
R1149 VDD1.n153 VDD1.n152 0.155672
R1150 VDD1.n153 VDD1.n132 0.155672
R1151 VDD1.n161 VDD1.n132 0.155672
R1152 VDD1.n162 VDD1.n161 0.155672
R1153 VDD1.n162 VDD1.n128 0.155672
R1154 VDD1.n170 VDD1.n128 0.155672
R1155 VDD1.n171 VDD1.n170 0.155672
R1156 VDD1.n171 VDD1.n124 0.155672
R1157 VDD1.n178 VDD1.n124 0.155672
R1158 VDD1.n179 VDD1.n178 0.155672
R1159 VDD1.n179 VDD1.n120 0.155672
R1160 VDD1.n186 VDD1.n120 0.155672
R1161 VDD1.n187 VDD1.n186 0.155672
R1162 VDD1.n187 VDD1.n116 0.155672
R1163 VDD1.n194 VDD1.n116 0.155672
R1164 VDD1.n195 VDD1.n194 0.155672
R1165 VDD1.n195 VDD1.n112 0.155672
R1166 VDD1.n202 VDD1.n112 0.155672
R1167 VDD1.n203 VDD1.n202 0.155672
R1168 VDD1.n203 VDD1.n108 0.155672
R1169 VDD1.n210 VDD1.n108 0.155672
R1170 B.n1235 B.n1234 585
R1171 B.n1236 B.n1235 585
R1172 B.n466 B.n192 585
R1173 B.n465 B.n464 585
R1174 B.n463 B.n462 585
R1175 B.n461 B.n460 585
R1176 B.n459 B.n458 585
R1177 B.n457 B.n456 585
R1178 B.n455 B.n454 585
R1179 B.n453 B.n452 585
R1180 B.n451 B.n450 585
R1181 B.n449 B.n448 585
R1182 B.n447 B.n446 585
R1183 B.n445 B.n444 585
R1184 B.n443 B.n442 585
R1185 B.n441 B.n440 585
R1186 B.n439 B.n438 585
R1187 B.n437 B.n436 585
R1188 B.n435 B.n434 585
R1189 B.n433 B.n432 585
R1190 B.n431 B.n430 585
R1191 B.n429 B.n428 585
R1192 B.n427 B.n426 585
R1193 B.n425 B.n424 585
R1194 B.n423 B.n422 585
R1195 B.n421 B.n420 585
R1196 B.n419 B.n418 585
R1197 B.n417 B.n416 585
R1198 B.n415 B.n414 585
R1199 B.n413 B.n412 585
R1200 B.n411 B.n410 585
R1201 B.n409 B.n408 585
R1202 B.n407 B.n406 585
R1203 B.n405 B.n404 585
R1204 B.n403 B.n402 585
R1205 B.n401 B.n400 585
R1206 B.n399 B.n398 585
R1207 B.n397 B.n396 585
R1208 B.n395 B.n394 585
R1209 B.n393 B.n392 585
R1210 B.n391 B.n390 585
R1211 B.n389 B.n388 585
R1212 B.n387 B.n386 585
R1213 B.n385 B.n384 585
R1214 B.n383 B.n382 585
R1215 B.n381 B.n380 585
R1216 B.n379 B.n378 585
R1217 B.n377 B.n376 585
R1218 B.n375 B.n374 585
R1219 B.n373 B.n372 585
R1220 B.n371 B.n370 585
R1221 B.n369 B.n368 585
R1222 B.n367 B.n366 585
R1223 B.n365 B.n364 585
R1224 B.n363 B.n362 585
R1225 B.n361 B.n360 585
R1226 B.n359 B.n358 585
R1227 B.n357 B.n356 585
R1228 B.n355 B.n354 585
R1229 B.n353 B.n352 585
R1230 B.n351 B.n350 585
R1231 B.n349 B.n348 585
R1232 B.n347 B.n346 585
R1233 B.n345 B.n344 585
R1234 B.n343 B.n342 585
R1235 B.n340 B.n339 585
R1236 B.n338 B.n337 585
R1237 B.n336 B.n335 585
R1238 B.n334 B.n333 585
R1239 B.n332 B.n331 585
R1240 B.n330 B.n329 585
R1241 B.n328 B.n327 585
R1242 B.n326 B.n325 585
R1243 B.n324 B.n323 585
R1244 B.n322 B.n321 585
R1245 B.n320 B.n319 585
R1246 B.n318 B.n317 585
R1247 B.n316 B.n315 585
R1248 B.n314 B.n313 585
R1249 B.n312 B.n311 585
R1250 B.n310 B.n309 585
R1251 B.n308 B.n307 585
R1252 B.n306 B.n305 585
R1253 B.n304 B.n303 585
R1254 B.n302 B.n301 585
R1255 B.n300 B.n299 585
R1256 B.n298 B.n297 585
R1257 B.n296 B.n295 585
R1258 B.n294 B.n293 585
R1259 B.n292 B.n291 585
R1260 B.n290 B.n289 585
R1261 B.n288 B.n287 585
R1262 B.n286 B.n285 585
R1263 B.n284 B.n283 585
R1264 B.n282 B.n281 585
R1265 B.n280 B.n279 585
R1266 B.n278 B.n277 585
R1267 B.n276 B.n275 585
R1268 B.n274 B.n273 585
R1269 B.n272 B.n271 585
R1270 B.n270 B.n269 585
R1271 B.n268 B.n267 585
R1272 B.n266 B.n265 585
R1273 B.n264 B.n263 585
R1274 B.n262 B.n261 585
R1275 B.n260 B.n259 585
R1276 B.n258 B.n257 585
R1277 B.n256 B.n255 585
R1278 B.n254 B.n253 585
R1279 B.n252 B.n251 585
R1280 B.n250 B.n249 585
R1281 B.n248 B.n247 585
R1282 B.n246 B.n245 585
R1283 B.n244 B.n243 585
R1284 B.n242 B.n241 585
R1285 B.n240 B.n239 585
R1286 B.n238 B.n237 585
R1287 B.n236 B.n235 585
R1288 B.n234 B.n233 585
R1289 B.n232 B.n231 585
R1290 B.n230 B.n229 585
R1291 B.n228 B.n227 585
R1292 B.n226 B.n225 585
R1293 B.n224 B.n223 585
R1294 B.n222 B.n221 585
R1295 B.n220 B.n219 585
R1296 B.n218 B.n217 585
R1297 B.n216 B.n215 585
R1298 B.n214 B.n213 585
R1299 B.n212 B.n211 585
R1300 B.n210 B.n209 585
R1301 B.n208 B.n207 585
R1302 B.n206 B.n205 585
R1303 B.n204 B.n203 585
R1304 B.n202 B.n201 585
R1305 B.n200 B.n199 585
R1306 B.n124 B.n123 585
R1307 B.n1239 B.n1238 585
R1308 B.n1233 B.n193 585
R1309 B.n193 B.n121 585
R1310 B.n1232 B.n120 585
R1311 B.n1243 B.n120 585
R1312 B.n1231 B.n119 585
R1313 B.n1244 B.n119 585
R1314 B.n1230 B.n118 585
R1315 B.n1245 B.n118 585
R1316 B.n1229 B.n1228 585
R1317 B.n1228 B.n114 585
R1318 B.n1227 B.n113 585
R1319 B.n1251 B.n113 585
R1320 B.n1226 B.n112 585
R1321 B.n1252 B.n112 585
R1322 B.n1225 B.n111 585
R1323 B.n1253 B.n111 585
R1324 B.n1224 B.n1223 585
R1325 B.n1223 B.n110 585
R1326 B.n1222 B.n106 585
R1327 B.n1259 B.n106 585
R1328 B.n1221 B.n105 585
R1329 B.n1260 B.n105 585
R1330 B.n1220 B.n104 585
R1331 B.n1261 B.n104 585
R1332 B.n1219 B.n1218 585
R1333 B.n1218 B.n100 585
R1334 B.n1217 B.n99 585
R1335 B.n1267 B.n99 585
R1336 B.n1216 B.n98 585
R1337 B.n1268 B.n98 585
R1338 B.n1215 B.n97 585
R1339 B.n1269 B.n97 585
R1340 B.n1214 B.n1213 585
R1341 B.n1213 B.n93 585
R1342 B.n1212 B.n92 585
R1343 B.n1275 B.n92 585
R1344 B.n1211 B.n91 585
R1345 B.n1276 B.n91 585
R1346 B.n1210 B.n90 585
R1347 B.n1277 B.n90 585
R1348 B.n1209 B.n1208 585
R1349 B.n1208 B.n86 585
R1350 B.n1207 B.n85 585
R1351 B.n1283 B.n85 585
R1352 B.n1206 B.n84 585
R1353 B.n1284 B.n84 585
R1354 B.n1205 B.n83 585
R1355 B.n1285 B.n83 585
R1356 B.n1204 B.n1203 585
R1357 B.n1203 B.n79 585
R1358 B.n1202 B.n78 585
R1359 B.n1291 B.n78 585
R1360 B.n1201 B.n77 585
R1361 B.n1292 B.n77 585
R1362 B.n1200 B.n76 585
R1363 B.n1293 B.n76 585
R1364 B.n1199 B.n1198 585
R1365 B.n1198 B.n72 585
R1366 B.n1197 B.n71 585
R1367 B.n1299 B.n71 585
R1368 B.n1196 B.n70 585
R1369 B.n1300 B.n70 585
R1370 B.n1195 B.n69 585
R1371 B.n1301 B.n69 585
R1372 B.n1194 B.n1193 585
R1373 B.n1193 B.n65 585
R1374 B.n1192 B.n64 585
R1375 B.n1307 B.n64 585
R1376 B.n1191 B.n63 585
R1377 B.n1308 B.n63 585
R1378 B.n1190 B.n62 585
R1379 B.n1309 B.n62 585
R1380 B.n1189 B.n1188 585
R1381 B.n1188 B.n58 585
R1382 B.n1187 B.n57 585
R1383 B.n1315 B.n57 585
R1384 B.n1186 B.n56 585
R1385 B.n1316 B.n56 585
R1386 B.n1185 B.n55 585
R1387 B.n1317 B.n55 585
R1388 B.n1184 B.n1183 585
R1389 B.n1183 B.n51 585
R1390 B.n1182 B.n50 585
R1391 B.n1323 B.n50 585
R1392 B.n1181 B.n49 585
R1393 B.n1324 B.n49 585
R1394 B.n1180 B.n48 585
R1395 B.n1325 B.n48 585
R1396 B.n1179 B.n1178 585
R1397 B.n1178 B.n44 585
R1398 B.n1177 B.n43 585
R1399 B.n1331 B.n43 585
R1400 B.n1176 B.n42 585
R1401 B.n1332 B.n42 585
R1402 B.n1175 B.n41 585
R1403 B.n1333 B.n41 585
R1404 B.n1174 B.n1173 585
R1405 B.n1173 B.n37 585
R1406 B.n1172 B.n36 585
R1407 B.n1339 B.n36 585
R1408 B.n1171 B.n35 585
R1409 B.n1340 B.n35 585
R1410 B.n1170 B.n34 585
R1411 B.n1341 B.n34 585
R1412 B.n1169 B.n1168 585
R1413 B.n1168 B.n30 585
R1414 B.n1167 B.n29 585
R1415 B.n1347 B.n29 585
R1416 B.n1166 B.n28 585
R1417 B.n1348 B.n28 585
R1418 B.n1165 B.n27 585
R1419 B.n1349 B.n27 585
R1420 B.n1164 B.n1163 585
R1421 B.n1163 B.n23 585
R1422 B.n1162 B.n22 585
R1423 B.n1355 B.n22 585
R1424 B.n1161 B.n21 585
R1425 B.n1356 B.n21 585
R1426 B.n1160 B.n20 585
R1427 B.n1357 B.n20 585
R1428 B.n1159 B.n1158 585
R1429 B.n1158 B.n19 585
R1430 B.n1157 B.n15 585
R1431 B.n1363 B.n15 585
R1432 B.n1156 B.n14 585
R1433 B.n1364 B.n14 585
R1434 B.n1155 B.n13 585
R1435 B.n1365 B.n13 585
R1436 B.n1154 B.n1153 585
R1437 B.n1153 B.n12 585
R1438 B.n1152 B.n1151 585
R1439 B.n1152 B.n8 585
R1440 B.n1150 B.n7 585
R1441 B.n1372 B.n7 585
R1442 B.n1149 B.n6 585
R1443 B.n1373 B.n6 585
R1444 B.n1148 B.n5 585
R1445 B.n1374 B.n5 585
R1446 B.n1147 B.n1146 585
R1447 B.n1146 B.n4 585
R1448 B.n1145 B.n467 585
R1449 B.n1145 B.n1144 585
R1450 B.n1135 B.n468 585
R1451 B.n469 B.n468 585
R1452 B.n1137 B.n1136 585
R1453 B.n1138 B.n1137 585
R1454 B.n1134 B.n474 585
R1455 B.n474 B.n473 585
R1456 B.n1133 B.n1132 585
R1457 B.n1132 B.n1131 585
R1458 B.n476 B.n475 585
R1459 B.n1124 B.n476 585
R1460 B.n1123 B.n1122 585
R1461 B.n1125 B.n1123 585
R1462 B.n1121 B.n481 585
R1463 B.n481 B.n480 585
R1464 B.n1120 B.n1119 585
R1465 B.n1119 B.n1118 585
R1466 B.n483 B.n482 585
R1467 B.n484 B.n483 585
R1468 B.n1111 B.n1110 585
R1469 B.n1112 B.n1111 585
R1470 B.n1109 B.n489 585
R1471 B.n489 B.n488 585
R1472 B.n1108 B.n1107 585
R1473 B.n1107 B.n1106 585
R1474 B.n491 B.n490 585
R1475 B.n492 B.n491 585
R1476 B.n1099 B.n1098 585
R1477 B.n1100 B.n1099 585
R1478 B.n1097 B.n497 585
R1479 B.n497 B.n496 585
R1480 B.n1096 B.n1095 585
R1481 B.n1095 B.n1094 585
R1482 B.n499 B.n498 585
R1483 B.n500 B.n499 585
R1484 B.n1087 B.n1086 585
R1485 B.n1088 B.n1087 585
R1486 B.n1085 B.n505 585
R1487 B.n505 B.n504 585
R1488 B.n1084 B.n1083 585
R1489 B.n1083 B.n1082 585
R1490 B.n507 B.n506 585
R1491 B.n508 B.n507 585
R1492 B.n1075 B.n1074 585
R1493 B.n1076 B.n1075 585
R1494 B.n1073 B.n513 585
R1495 B.n513 B.n512 585
R1496 B.n1072 B.n1071 585
R1497 B.n1071 B.n1070 585
R1498 B.n515 B.n514 585
R1499 B.n516 B.n515 585
R1500 B.n1063 B.n1062 585
R1501 B.n1064 B.n1063 585
R1502 B.n1061 B.n521 585
R1503 B.n521 B.n520 585
R1504 B.n1060 B.n1059 585
R1505 B.n1059 B.n1058 585
R1506 B.n523 B.n522 585
R1507 B.n524 B.n523 585
R1508 B.n1051 B.n1050 585
R1509 B.n1052 B.n1051 585
R1510 B.n1049 B.n529 585
R1511 B.n529 B.n528 585
R1512 B.n1048 B.n1047 585
R1513 B.n1047 B.n1046 585
R1514 B.n531 B.n530 585
R1515 B.n532 B.n531 585
R1516 B.n1039 B.n1038 585
R1517 B.n1040 B.n1039 585
R1518 B.n1037 B.n537 585
R1519 B.n537 B.n536 585
R1520 B.n1036 B.n1035 585
R1521 B.n1035 B.n1034 585
R1522 B.n539 B.n538 585
R1523 B.n540 B.n539 585
R1524 B.n1027 B.n1026 585
R1525 B.n1028 B.n1027 585
R1526 B.n1025 B.n545 585
R1527 B.n545 B.n544 585
R1528 B.n1024 B.n1023 585
R1529 B.n1023 B.n1022 585
R1530 B.n547 B.n546 585
R1531 B.n548 B.n547 585
R1532 B.n1015 B.n1014 585
R1533 B.n1016 B.n1015 585
R1534 B.n1013 B.n553 585
R1535 B.n553 B.n552 585
R1536 B.n1012 B.n1011 585
R1537 B.n1011 B.n1010 585
R1538 B.n555 B.n554 585
R1539 B.n556 B.n555 585
R1540 B.n1003 B.n1002 585
R1541 B.n1004 B.n1003 585
R1542 B.n1001 B.n561 585
R1543 B.n561 B.n560 585
R1544 B.n1000 B.n999 585
R1545 B.n999 B.n998 585
R1546 B.n563 B.n562 585
R1547 B.n564 B.n563 585
R1548 B.n991 B.n990 585
R1549 B.n992 B.n991 585
R1550 B.n989 B.n569 585
R1551 B.n569 B.n568 585
R1552 B.n988 B.n987 585
R1553 B.n987 B.n986 585
R1554 B.n571 B.n570 585
R1555 B.n572 B.n571 585
R1556 B.n979 B.n978 585
R1557 B.n980 B.n979 585
R1558 B.n977 B.n577 585
R1559 B.n577 B.n576 585
R1560 B.n976 B.n975 585
R1561 B.n975 B.n974 585
R1562 B.n579 B.n578 585
R1563 B.n967 B.n579 585
R1564 B.n966 B.n965 585
R1565 B.n968 B.n966 585
R1566 B.n964 B.n584 585
R1567 B.n584 B.n583 585
R1568 B.n963 B.n962 585
R1569 B.n962 B.n961 585
R1570 B.n586 B.n585 585
R1571 B.n587 B.n586 585
R1572 B.n954 B.n953 585
R1573 B.n955 B.n954 585
R1574 B.n952 B.n592 585
R1575 B.n592 B.n591 585
R1576 B.n951 B.n950 585
R1577 B.n950 B.n949 585
R1578 B.n594 B.n593 585
R1579 B.n595 B.n594 585
R1580 B.n945 B.n944 585
R1581 B.n598 B.n597 585
R1582 B.n941 B.n940 585
R1583 B.n942 B.n941 585
R1584 B.n939 B.n666 585
R1585 B.n938 B.n937 585
R1586 B.n936 B.n935 585
R1587 B.n934 B.n933 585
R1588 B.n932 B.n931 585
R1589 B.n930 B.n929 585
R1590 B.n928 B.n927 585
R1591 B.n926 B.n925 585
R1592 B.n924 B.n923 585
R1593 B.n922 B.n921 585
R1594 B.n920 B.n919 585
R1595 B.n918 B.n917 585
R1596 B.n916 B.n915 585
R1597 B.n914 B.n913 585
R1598 B.n912 B.n911 585
R1599 B.n910 B.n909 585
R1600 B.n908 B.n907 585
R1601 B.n906 B.n905 585
R1602 B.n904 B.n903 585
R1603 B.n902 B.n901 585
R1604 B.n900 B.n899 585
R1605 B.n898 B.n897 585
R1606 B.n896 B.n895 585
R1607 B.n894 B.n893 585
R1608 B.n892 B.n891 585
R1609 B.n890 B.n889 585
R1610 B.n888 B.n887 585
R1611 B.n886 B.n885 585
R1612 B.n884 B.n883 585
R1613 B.n882 B.n881 585
R1614 B.n880 B.n879 585
R1615 B.n878 B.n877 585
R1616 B.n876 B.n875 585
R1617 B.n874 B.n873 585
R1618 B.n872 B.n871 585
R1619 B.n870 B.n869 585
R1620 B.n868 B.n867 585
R1621 B.n866 B.n865 585
R1622 B.n864 B.n863 585
R1623 B.n862 B.n861 585
R1624 B.n860 B.n859 585
R1625 B.n858 B.n857 585
R1626 B.n856 B.n855 585
R1627 B.n854 B.n853 585
R1628 B.n852 B.n851 585
R1629 B.n850 B.n849 585
R1630 B.n848 B.n847 585
R1631 B.n846 B.n845 585
R1632 B.n844 B.n843 585
R1633 B.n842 B.n841 585
R1634 B.n840 B.n839 585
R1635 B.n838 B.n837 585
R1636 B.n836 B.n835 585
R1637 B.n834 B.n833 585
R1638 B.n832 B.n831 585
R1639 B.n830 B.n829 585
R1640 B.n828 B.n827 585
R1641 B.n826 B.n825 585
R1642 B.n824 B.n823 585
R1643 B.n822 B.n821 585
R1644 B.n820 B.n819 585
R1645 B.n817 B.n816 585
R1646 B.n815 B.n814 585
R1647 B.n813 B.n812 585
R1648 B.n811 B.n810 585
R1649 B.n809 B.n808 585
R1650 B.n807 B.n806 585
R1651 B.n805 B.n804 585
R1652 B.n803 B.n802 585
R1653 B.n801 B.n800 585
R1654 B.n799 B.n798 585
R1655 B.n797 B.n796 585
R1656 B.n795 B.n794 585
R1657 B.n793 B.n792 585
R1658 B.n791 B.n790 585
R1659 B.n789 B.n788 585
R1660 B.n787 B.n786 585
R1661 B.n785 B.n784 585
R1662 B.n783 B.n782 585
R1663 B.n781 B.n780 585
R1664 B.n779 B.n778 585
R1665 B.n777 B.n776 585
R1666 B.n775 B.n774 585
R1667 B.n773 B.n772 585
R1668 B.n771 B.n770 585
R1669 B.n769 B.n768 585
R1670 B.n767 B.n766 585
R1671 B.n765 B.n764 585
R1672 B.n763 B.n762 585
R1673 B.n761 B.n760 585
R1674 B.n759 B.n758 585
R1675 B.n757 B.n756 585
R1676 B.n755 B.n754 585
R1677 B.n753 B.n752 585
R1678 B.n751 B.n750 585
R1679 B.n749 B.n748 585
R1680 B.n747 B.n746 585
R1681 B.n745 B.n744 585
R1682 B.n743 B.n742 585
R1683 B.n741 B.n740 585
R1684 B.n739 B.n738 585
R1685 B.n737 B.n736 585
R1686 B.n735 B.n734 585
R1687 B.n733 B.n732 585
R1688 B.n731 B.n730 585
R1689 B.n729 B.n728 585
R1690 B.n727 B.n726 585
R1691 B.n725 B.n724 585
R1692 B.n723 B.n722 585
R1693 B.n721 B.n720 585
R1694 B.n719 B.n718 585
R1695 B.n717 B.n716 585
R1696 B.n715 B.n714 585
R1697 B.n713 B.n712 585
R1698 B.n711 B.n710 585
R1699 B.n709 B.n708 585
R1700 B.n707 B.n706 585
R1701 B.n705 B.n704 585
R1702 B.n703 B.n702 585
R1703 B.n701 B.n700 585
R1704 B.n699 B.n698 585
R1705 B.n697 B.n696 585
R1706 B.n695 B.n694 585
R1707 B.n693 B.n692 585
R1708 B.n691 B.n690 585
R1709 B.n689 B.n688 585
R1710 B.n687 B.n686 585
R1711 B.n685 B.n684 585
R1712 B.n683 B.n682 585
R1713 B.n681 B.n680 585
R1714 B.n679 B.n678 585
R1715 B.n677 B.n676 585
R1716 B.n675 B.n674 585
R1717 B.n673 B.n672 585
R1718 B.n946 B.n596 585
R1719 B.n596 B.n595 585
R1720 B.n948 B.n947 585
R1721 B.n949 B.n948 585
R1722 B.n590 B.n589 585
R1723 B.n591 B.n590 585
R1724 B.n957 B.n956 585
R1725 B.n956 B.n955 585
R1726 B.n958 B.n588 585
R1727 B.n588 B.n587 585
R1728 B.n960 B.n959 585
R1729 B.n961 B.n960 585
R1730 B.n582 B.n581 585
R1731 B.n583 B.n582 585
R1732 B.n970 B.n969 585
R1733 B.n969 B.n968 585
R1734 B.n971 B.n580 585
R1735 B.n967 B.n580 585
R1736 B.n973 B.n972 585
R1737 B.n974 B.n973 585
R1738 B.n575 B.n574 585
R1739 B.n576 B.n575 585
R1740 B.n982 B.n981 585
R1741 B.n981 B.n980 585
R1742 B.n983 B.n573 585
R1743 B.n573 B.n572 585
R1744 B.n985 B.n984 585
R1745 B.n986 B.n985 585
R1746 B.n567 B.n566 585
R1747 B.n568 B.n567 585
R1748 B.n994 B.n993 585
R1749 B.n993 B.n992 585
R1750 B.n995 B.n565 585
R1751 B.n565 B.n564 585
R1752 B.n997 B.n996 585
R1753 B.n998 B.n997 585
R1754 B.n559 B.n558 585
R1755 B.n560 B.n559 585
R1756 B.n1006 B.n1005 585
R1757 B.n1005 B.n1004 585
R1758 B.n1007 B.n557 585
R1759 B.n557 B.n556 585
R1760 B.n1009 B.n1008 585
R1761 B.n1010 B.n1009 585
R1762 B.n551 B.n550 585
R1763 B.n552 B.n551 585
R1764 B.n1018 B.n1017 585
R1765 B.n1017 B.n1016 585
R1766 B.n1019 B.n549 585
R1767 B.n549 B.n548 585
R1768 B.n1021 B.n1020 585
R1769 B.n1022 B.n1021 585
R1770 B.n543 B.n542 585
R1771 B.n544 B.n543 585
R1772 B.n1030 B.n1029 585
R1773 B.n1029 B.n1028 585
R1774 B.n1031 B.n541 585
R1775 B.n541 B.n540 585
R1776 B.n1033 B.n1032 585
R1777 B.n1034 B.n1033 585
R1778 B.n535 B.n534 585
R1779 B.n536 B.n535 585
R1780 B.n1042 B.n1041 585
R1781 B.n1041 B.n1040 585
R1782 B.n1043 B.n533 585
R1783 B.n533 B.n532 585
R1784 B.n1045 B.n1044 585
R1785 B.n1046 B.n1045 585
R1786 B.n527 B.n526 585
R1787 B.n528 B.n527 585
R1788 B.n1054 B.n1053 585
R1789 B.n1053 B.n1052 585
R1790 B.n1055 B.n525 585
R1791 B.n525 B.n524 585
R1792 B.n1057 B.n1056 585
R1793 B.n1058 B.n1057 585
R1794 B.n519 B.n518 585
R1795 B.n520 B.n519 585
R1796 B.n1066 B.n1065 585
R1797 B.n1065 B.n1064 585
R1798 B.n1067 B.n517 585
R1799 B.n517 B.n516 585
R1800 B.n1069 B.n1068 585
R1801 B.n1070 B.n1069 585
R1802 B.n511 B.n510 585
R1803 B.n512 B.n511 585
R1804 B.n1078 B.n1077 585
R1805 B.n1077 B.n1076 585
R1806 B.n1079 B.n509 585
R1807 B.n509 B.n508 585
R1808 B.n1081 B.n1080 585
R1809 B.n1082 B.n1081 585
R1810 B.n503 B.n502 585
R1811 B.n504 B.n503 585
R1812 B.n1090 B.n1089 585
R1813 B.n1089 B.n1088 585
R1814 B.n1091 B.n501 585
R1815 B.n501 B.n500 585
R1816 B.n1093 B.n1092 585
R1817 B.n1094 B.n1093 585
R1818 B.n495 B.n494 585
R1819 B.n496 B.n495 585
R1820 B.n1102 B.n1101 585
R1821 B.n1101 B.n1100 585
R1822 B.n1103 B.n493 585
R1823 B.n493 B.n492 585
R1824 B.n1105 B.n1104 585
R1825 B.n1106 B.n1105 585
R1826 B.n487 B.n486 585
R1827 B.n488 B.n487 585
R1828 B.n1114 B.n1113 585
R1829 B.n1113 B.n1112 585
R1830 B.n1115 B.n485 585
R1831 B.n485 B.n484 585
R1832 B.n1117 B.n1116 585
R1833 B.n1118 B.n1117 585
R1834 B.n479 B.n478 585
R1835 B.n480 B.n479 585
R1836 B.n1127 B.n1126 585
R1837 B.n1126 B.n1125 585
R1838 B.n1128 B.n477 585
R1839 B.n1124 B.n477 585
R1840 B.n1130 B.n1129 585
R1841 B.n1131 B.n1130 585
R1842 B.n472 B.n471 585
R1843 B.n473 B.n472 585
R1844 B.n1140 B.n1139 585
R1845 B.n1139 B.n1138 585
R1846 B.n1141 B.n470 585
R1847 B.n470 B.n469 585
R1848 B.n1143 B.n1142 585
R1849 B.n1144 B.n1143 585
R1850 B.n3 B.n0 585
R1851 B.n4 B.n3 585
R1852 B.n1371 B.n1 585
R1853 B.n1372 B.n1371 585
R1854 B.n1370 B.n1369 585
R1855 B.n1370 B.n8 585
R1856 B.n1368 B.n9 585
R1857 B.n12 B.n9 585
R1858 B.n1367 B.n1366 585
R1859 B.n1366 B.n1365 585
R1860 B.n11 B.n10 585
R1861 B.n1364 B.n11 585
R1862 B.n1362 B.n1361 585
R1863 B.n1363 B.n1362 585
R1864 B.n1360 B.n16 585
R1865 B.n19 B.n16 585
R1866 B.n1359 B.n1358 585
R1867 B.n1358 B.n1357 585
R1868 B.n18 B.n17 585
R1869 B.n1356 B.n18 585
R1870 B.n1354 B.n1353 585
R1871 B.n1355 B.n1354 585
R1872 B.n1352 B.n24 585
R1873 B.n24 B.n23 585
R1874 B.n1351 B.n1350 585
R1875 B.n1350 B.n1349 585
R1876 B.n26 B.n25 585
R1877 B.n1348 B.n26 585
R1878 B.n1346 B.n1345 585
R1879 B.n1347 B.n1346 585
R1880 B.n1344 B.n31 585
R1881 B.n31 B.n30 585
R1882 B.n1343 B.n1342 585
R1883 B.n1342 B.n1341 585
R1884 B.n33 B.n32 585
R1885 B.n1340 B.n33 585
R1886 B.n1338 B.n1337 585
R1887 B.n1339 B.n1338 585
R1888 B.n1336 B.n38 585
R1889 B.n38 B.n37 585
R1890 B.n1335 B.n1334 585
R1891 B.n1334 B.n1333 585
R1892 B.n40 B.n39 585
R1893 B.n1332 B.n40 585
R1894 B.n1330 B.n1329 585
R1895 B.n1331 B.n1330 585
R1896 B.n1328 B.n45 585
R1897 B.n45 B.n44 585
R1898 B.n1327 B.n1326 585
R1899 B.n1326 B.n1325 585
R1900 B.n47 B.n46 585
R1901 B.n1324 B.n47 585
R1902 B.n1322 B.n1321 585
R1903 B.n1323 B.n1322 585
R1904 B.n1320 B.n52 585
R1905 B.n52 B.n51 585
R1906 B.n1319 B.n1318 585
R1907 B.n1318 B.n1317 585
R1908 B.n54 B.n53 585
R1909 B.n1316 B.n54 585
R1910 B.n1314 B.n1313 585
R1911 B.n1315 B.n1314 585
R1912 B.n1312 B.n59 585
R1913 B.n59 B.n58 585
R1914 B.n1311 B.n1310 585
R1915 B.n1310 B.n1309 585
R1916 B.n61 B.n60 585
R1917 B.n1308 B.n61 585
R1918 B.n1306 B.n1305 585
R1919 B.n1307 B.n1306 585
R1920 B.n1304 B.n66 585
R1921 B.n66 B.n65 585
R1922 B.n1303 B.n1302 585
R1923 B.n1302 B.n1301 585
R1924 B.n68 B.n67 585
R1925 B.n1300 B.n68 585
R1926 B.n1298 B.n1297 585
R1927 B.n1299 B.n1298 585
R1928 B.n1296 B.n73 585
R1929 B.n73 B.n72 585
R1930 B.n1295 B.n1294 585
R1931 B.n1294 B.n1293 585
R1932 B.n75 B.n74 585
R1933 B.n1292 B.n75 585
R1934 B.n1290 B.n1289 585
R1935 B.n1291 B.n1290 585
R1936 B.n1288 B.n80 585
R1937 B.n80 B.n79 585
R1938 B.n1287 B.n1286 585
R1939 B.n1286 B.n1285 585
R1940 B.n82 B.n81 585
R1941 B.n1284 B.n82 585
R1942 B.n1282 B.n1281 585
R1943 B.n1283 B.n1282 585
R1944 B.n1280 B.n87 585
R1945 B.n87 B.n86 585
R1946 B.n1279 B.n1278 585
R1947 B.n1278 B.n1277 585
R1948 B.n89 B.n88 585
R1949 B.n1276 B.n89 585
R1950 B.n1274 B.n1273 585
R1951 B.n1275 B.n1274 585
R1952 B.n1272 B.n94 585
R1953 B.n94 B.n93 585
R1954 B.n1271 B.n1270 585
R1955 B.n1270 B.n1269 585
R1956 B.n96 B.n95 585
R1957 B.n1268 B.n96 585
R1958 B.n1266 B.n1265 585
R1959 B.n1267 B.n1266 585
R1960 B.n1264 B.n101 585
R1961 B.n101 B.n100 585
R1962 B.n1263 B.n1262 585
R1963 B.n1262 B.n1261 585
R1964 B.n103 B.n102 585
R1965 B.n1260 B.n103 585
R1966 B.n1258 B.n1257 585
R1967 B.n1259 B.n1258 585
R1968 B.n1256 B.n107 585
R1969 B.n110 B.n107 585
R1970 B.n1255 B.n1254 585
R1971 B.n1254 B.n1253 585
R1972 B.n109 B.n108 585
R1973 B.n1252 B.n109 585
R1974 B.n1250 B.n1249 585
R1975 B.n1251 B.n1250 585
R1976 B.n1248 B.n115 585
R1977 B.n115 B.n114 585
R1978 B.n1247 B.n1246 585
R1979 B.n1246 B.n1245 585
R1980 B.n117 B.n116 585
R1981 B.n1244 B.n117 585
R1982 B.n1242 B.n1241 585
R1983 B.n1243 B.n1242 585
R1984 B.n1240 B.n122 585
R1985 B.n122 B.n121 585
R1986 B.n1375 B.n1374 585
R1987 B.n1373 B.n2 585
R1988 B.n1238 B.n122 478.086
R1989 B.n1235 B.n193 478.086
R1990 B.n672 B.n594 478.086
R1991 B.n944 B.n596 478.086
R1992 B.n194 B.t16 476.397
R1993 B.n669 B.t13 476.397
R1994 B.n196 B.t22 476.397
R1995 B.n667 B.t20 476.397
R1996 B.n195 B.t17 411.233
R1997 B.n670 B.t12 411.233
R1998 B.n197 B.t23 411.233
R1999 B.n668 B.t19 411.233
R2000 B.n196 B.t21 363.714
R2001 B.n194 B.t14 363.714
R2002 B.n669 B.t10 363.714
R2003 B.n667 B.t18 363.714
R2004 B.n1236 B.n191 256.663
R2005 B.n1236 B.n190 256.663
R2006 B.n1236 B.n189 256.663
R2007 B.n1236 B.n188 256.663
R2008 B.n1236 B.n187 256.663
R2009 B.n1236 B.n186 256.663
R2010 B.n1236 B.n185 256.663
R2011 B.n1236 B.n184 256.663
R2012 B.n1236 B.n183 256.663
R2013 B.n1236 B.n182 256.663
R2014 B.n1236 B.n181 256.663
R2015 B.n1236 B.n180 256.663
R2016 B.n1236 B.n179 256.663
R2017 B.n1236 B.n178 256.663
R2018 B.n1236 B.n177 256.663
R2019 B.n1236 B.n176 256.663
R2020 B.n1236 B.n175 256.663
R2021 B.n1236 B.n174 256.663
R2022 B.n1236 B.n173 256.663
R2023 B.n1236 B.n172 256.663
R2024 B.n1236 B.n171 256.663
R2025 B.n1236 B.n170 256.663
R2026 B.n1236 B.n169 256.663
R2027 B.n1236 B.n168 256.663
R2028 B.n1236 B.n167 256.663
R2029 B.n1236 B.n166 256.663
R2030 B.n1236 B.n165 256.663
R2031 B.n1236 B.n164 256.663
R2032 B.n1236 B.n163 256.663
R2033 B.n1236 B.n162 256.663
R2034 B.n1236 B.n161 256.663
R2035 B.n1236 B.n160 256.663
R2036 B.n1236 B.n159 256.663
R2037 B.n1236 B.n158 256.663
R2038 B.n1236 B.n157 256.663
R2039 B.n1236 B.n156 256.663
R2040 B.n1236 B.n155 256.663
R2041 B.n1236 B.n154 256.663
R2042 B.n1236 B.n153 256.663
R2043 B.n1236 B.n152 256.663
R2044 B.n1236 B.n151 256.663
R2045 B.n1236 B.n150 256.663
R2046 B.n1236 B.n149 256.663
R2047 B.n1236 B.n148 256.663
R2048 B.n1236 B.n147 256.663
R2049 B.n1236 B.n146 256.663
R2050 B.n1236 B.n145 256.663
R2051 B.n1236 B.n144 256.663
R2052 B.n1236 B.n143 256.663
R2053 B.n1236 B.n142 256.663
R2054 B.n1236 B.n141 256.663
R2055 B.n1236 B.n140 256.663
R2056 B.n1236 B.n139 256.663
R2057 B.n1236 B.n138 256.663
R2058 B.n1236 B.n137 256.663
R2059 B.n1236 B.n136 256.663
R2060 B.n1236 B.n135 256.663
R2061 B.n1236 B.n134 256.663
R2062 B.n1236 B.n133 256.663
R2063 B.n1236 B.n132 256.663
R2064 B.n1236 B.n131 256.663
R2065 B.n1236 B.n130 256.663
R2066 B.n1236 B.n129 256.663
R2067 B.n1236 B.n128 256.663
R2068 B.n1236 B.n127 256.663
R2069 B.n1236 B.n126 256.663
R2070 B.n1236 B.n125 256.663
R2071 B.n1237 B.n1236 256.663
R2072 B.n943 B.n942 256.663
R2073 B.n942 B.n599 256.663
R2074 B.n942 B.n600 256.663
R2075 B.n942 B.n601 256.663
R2076 B.n942 B.n602 256.663
R2077 B.n942 B.n603 256.663
R2078 B.n942 B.n604 256.663
R2079 B.n942 B.n605 256.663
R2080 B.n942 B.n606 256.663
R2081 B.n942 B.n607 256.663
R2082 B.n942 B.n608 256.663
R2083 B.n942 B.n609 256.663
R2084 B.n942 B.n610 256.663
R2085 B.n942 B.n611 256.663
R2086 B.n942 B.n612 256.663
R2087 B.n942 B.n613 256.663
R2088 B.n942 B.n614 256.663
R2089 B.n942 B.n615 256.663
R2090 B.n942 B.n616 256.663
R2091 B.n942 B.n617 256.663
R2092 B.n942 B.n618 256.663
R2093 B.n942 B.n619 256.663
R2094 B.n942 B.n620 256.663
R2095 B.n942 B.n621 256.663
R2096 B.n942 B.n622 256.663
R2097 B.n942 B.n623 256.663
R2098 B.n942 B.n624 256.663
R2099 B.n942 B.n625 256.663
R2100 B.n942 B.n626 256.663
R2101 B.n942 B.n627 256.663
R2102 B.n942 B.n628 256.663
R2103 B.n942 B.n629 256.663
R2104 B.n942 B.n630 256.663
R2105 B.n942 B.n631 256.663
R2106 B.n942 B.n632 256.663
R2107 B.n942 B.n633 256.663
R2108 B.n942 B.n634 256.663
R2109 B.n942 B.n635 256.663
R2110 B.n942 B.n636 256.663
R2111 B.n942 B.n637 256.663
R2112 B.n942 B.n638 256.663
R2113 B.n942 B.n639 256.663
R2114 B.n942 B.n640 256.663
R2115 B.n942 B.n641 256.663
R2116 B.n942 B.n642 256.663
R2117 B.n942 B.n643 256.663
R2118 B.n942 B.n644 256.663
R2119 B.n942 B.n645 256.663
R2120 B.n942 B.n646 256.663
R2121 B.n942 B.n647 256.663
R2122 B.n942 B.n648 256.663
R2123 B.n942 B.n649 256.663
R2124 B.n942 B.n650 256.663
R2125 B.n942 B.n651 256.663
R2126 B.n942 B.n652 256.663
R2127 B.n942 B.n653 256.663
R2128 B.n942 B.n654 256.663
R2129 B.n942 B.n655 256.663
R2130 B.n942 B.n656 256.663
R2131 B.n942 B.n657 256.663
R2132 B.n942 B.n658 256.663
R2133 B.n942 B.n659 256.663
R2134 B.n942 B.n660 256.663
R2135 B.n942 B.n661 256.663
R2136 B.n942 B.n662 256.663
R2137 B.n942 B.n663 256.663
R2138 B.n942 B.n664 256.663
R2139 B.n942 B.n665 256.663
R2140 B.n1377 B.n1376 256.663
R2141 B.n199 B.n124 163.367
R2142 B.n203 B.n202 163.367
R2143 B.n207 B.n206 163.367
R2144 B.n211 B.n210 163.367
R2145 B.n215 B.n214 163.367
R2146 B.n219 B.n218 163.367
R2147 B.n223 B.n222 163.367
R2148 B.n227 B.n226 163.367
R2149 B.n231 B.n230 163.367
R2150 B.n235 B.n234 163.367
R2151 B.n239 B.n238 163.367
R2152 B.n243 B.n242 163.367
R2153 B.n247 B.n246 163.367
R2154 B.n251 B.n250 163.367
R2155 B.n255 B.n254 163.367
R2156 B.n259 B.n258 163.367
R2157 B.n263 B.n262 163.367
R2158 B.n267 B.n266 163.367
R2159 B.n271 B.n270 163.367
R2160 B.n275 B.n274 163.367
R2161 B.n279 B.n278 163.367
R2162 B.n283 B.n282 163.367
R2163 B.n287 B.n286 163.367
R2164 B.n291 B.n290 163.367
R2165 B.n295 B.n294 163.367
R2166 B.n299 B.n298 163.367
R2167 B.n303 B.n302 163.367
R2168 B.n307 B.n306 163.367
R2169 B.n311 B.n310 163.367
R2170 B.n315 B.n314 163.367
R2171 B.n319 B.n318 163.367
R2172 B.n323 B.n322 163.367
R2173 B.n327 B.n326 163.367
R2174 B.n331 B.n330 163.367
R2175 B.n335 B.n334 163.367
R2176 B.n339 B.n338 163.367
R2177 B.n344 B.n343 163.367
R2178 B.n348 B.n347 163.367
R2179 B.n352 B.n351 163.367
R2180 B.n356 B.n355 163.367
R2181 B.n360 B.n359 163.367
R2182 B.n364 B.n363 163.367
R2183 B.n368 B.n367 163.367
R2184 B.n372 B.n371 163.367
R2185 B.n376 B.n375 163.367
R2186 B.n380 B.n379 163.367
R2187 B.n384 B.n383 163.367
R2188 B.n388 B.n387 163.367
R2189 B.n392 B.n391 163.367
R2190 B.n396 B.n395 163.367
R2191 B.n400 B.n399 163.367
R2192 B.n404 B.n403 163.367
R2193 B.n408 B.n407 163.367
R2194 B.n412 B.n411 163.367
R2195 B.n416 B.n415 163.367
R2196 B.n420 B.n419 163.367
R2197 B.n424 B.n423 163.367
R2198 B.n428 B.n427 163.367
R2199 B.n432 B.n431 163.367
R2200 B.n436 B.n435 163.367
R2201 B.n440 B.n439 163.367
R2202 B.n444 B.n443 163.367
R2203 B.n448 B.n447 163.367
R2204 B.n452 B.n451 163.367
R2205 B.n456 B.n455 163.367
R2206 B.n460 B.n459 163.367
R2207 B.n464 B.n463 163.367
R2208 B.n1235 B.n192 163.367
R2209 B.n950 B.n594 163.367
R2210 B.n950 B.n592 163.367
R2211 B.n954 B.n592 163.367
R2212 B.n954 B.n586 163.367
R2213 B.n962 B.n586 163.367
R2214 B.n962 B.n584 163.367
R2215 B.n966 B.n584 163.367
R2216 B.n966 B.n579 163.367
R2217 B.n975 B.n579 163.367
R2218 B.n975 B.n577 163.367
R2219 B.n979 B.n577 163.367
R2220 B.n979 B.n571 163.367
R2221 B.n987 B.n571 163.367
R2222 B.n987 B.n569 163.367
R2223 B.n991 B.n569 163.367
R2224 B.n991 B.n563 163.367
R2225 B.n999 B.n563 163.367
R2226 B.n999 B.n561 163.367
R2227 B.n1003 B.n561 163.367
R2228 B.n1003 B.n555 163.367
R2229 B.n1011 B.n555 163.367
R2230 B.n1011 B.n553 163.367
R2231 B.n1015 B.n553 163.367
R2232 B.n1015 B.n547 163.367
R2233 B.n1023 B.n547 163.367
R2234 B.n1023 B.n545 163.367
R2235 B.n1027 B.n545 163.367
R2236 B.n1027 B.n539 163.367
R2237 B.n1035 B.n539 163.367
R2238 B.n1035 B.n537 163.367
R2239 B.n1039 B.n537 163.367
R2240 B.n1039 B.n531 163.367
R2241 B.n1047 B.n531 163.367
R2242 B.n1047 B.n529 163.367
R2243 B.n1051 B.n529 163.367
R2244 B.n1051 B.n523 163.367
R2245 B.n1059 B.n523 163.367
R2246 B.n1059 B.n521 163.367
R2247 B.n1063 B.n521 163.367
R2248 B.n1063 B.n515 163.367
R2249 B.n1071 B.n515 163.367
R2250 B.n1071 B.n513 163.367
R2251 B.n1075 B.n513 163.367
R2252 B.n1075 B.n507 163.367
R2253 B.n1083 B.n507 163.367
R2254 B.n1083 B.n505 163.367
R2255 B.n1087 B.n505 163.367
R2256 B.n1087 B.n499 163.367
R2257 B.n1095 B.n499 163.367
R2258 B.n1095 B.n497 163.367
R2259 B.n1099 B.n497 163.367
R2260 B.n1099 B.n491 163.367
R2261 B.n1107 B.n491 163.367
R2262 B.n1107 B.n489 163.367
R2263 B.n1111 B.n489 163.367
R2264 B.n1111 B.n483 163.367
R2265 B.n1119 B.n483 163.367
R2266 B.n1119 B.n481 163.367
R2267 B.n1123 B.n481 163.367
R2268 B.n1123 B.n476 163.367
R2269 B.n1132 B.n476 163.367
R2270 B.n1132 B.n474 163.367
R2271 B.n1137 B.n474 163.367
R2272 B.n1137 B.n468 163.367
R2273 B.n1145 B.n468 163.367
R2274 B.n1146 B.n1145 163.367
R2275 B.n1146 B.n5 163.367
R2276 B.n6 B.n5 163.367
R2277 B.n7 B.n6 163.367
R2278 B.n1152 B.n7 163.367
R2279 B.n1153 B.n1152 163.367
R2280 B.n1153 B.n13 163.367
R2281 B.n14 B.n13 163.367
R2282 B.n15 B.n14 163.367
R2283 B.n1158 B.n15 163.367
R2284 B.n1158 B.n20 163.367
R2285 B.n21 B.n20 163.367
R2286 B.n22 B.n21 163.367
R2287 B.n1163 B.n22 163.367
R2288 B.n1163 B.n27 163.367
R2289 B.n28 B.n27 163.367
R2290 B.n29 B.n28 163.367
R2291 B.n1168 B.n29 163.367
R2292 B.n1168 B.n34 163.367
R2293 B.n35 B.n34 163.367
R2294 B.n36 B.n35 163.367
R2295 B.n1173 B.n36 163.367
R2296 B.n1173 B.n41 163.367
R2297 B.n42 B.n41 163.367
R2298 B.n43 B.n42 163.367
R2299 B.n1178 B.n43 163.367
R2300 B.n1178 B.n48 163.367
R2301 B.n49 B.n48 163.367
R2302 B.n50 B.n49 163.367
R2303 B.n1183 B.n50 163.367
R2304 B.n1183 B.n55 163.367
R2305 B.n56 B.n55 163.367
R2306 B.n57 B.n56 163.367
R2307 B.n1188 B.n57 163.367
R2308 B.n1188 B.n62 163.367
R2309 B.n63 B.n62 163.367
R2310 B.n64 B.n63 163.367
R2311 B.n1193 B.n64 163.367
R2312 B.n1193 B.n69 163.367
R2313 B.n70 B.n69 163.367
R2314 B.n71 B.n70 163.367
R2315 B.n1198 B.n71 163.367
R2316 B.n1198 B.n76 163.367
R2317 B.n77 B.n76 163.367
R2318 B.n78 B.n77 163.367
R2319 B.n1203 B.n78 163.367
R2320 B.n1203 B.n83 163.367
R2321 B.n84 B.n83 163.367
R2322 B.n85 B.n84 163.367
R2323 B.n1208 B.n85 163.367
R2324 B.n1208 B.n90 163.367
R2325 B.n91 B.n90 163.367
R2326 B.n92 B.n91 163.367
R2327 B.n1213 B.n92 163.367
R2328 B.n1213 B.n97 163.367
R2329 B.n98 B.n97 163.367
R2330 B.n99 B.n98 163.367
R2331 B.n1218 B.n99 163.367
R2332 B.n1218 B.n104 163.367
R2333 B.n105 B.n104 163.367
R2334 B.n106 B.n105 163.367
R2335 B.n1223 B.n106 163.367
R2336 B.n1223 B.n111 163.367
R2337 B.n112 B.n111 163.367
R2338 B.n113 B.n112 163.367
R2339 B.n1228 B.n113 163.367
R2340 B.n1228 B.n118 163.367
R2341 B.n119 B.n118 163.367
R2342 B.n120 B.n119 163.367
R2343 B.n193 B.n120 163.367
R2344 B.n941 B.n598 163.367
R2345 B.n941 B.n666 163.367
R2346 B.n937 B.n936 163.367
R2347 B.n933 B.n932 163.367
R2348 B.n929 B.n928 163.367
R2349 B.n925 B.n924 163.367
R2350 B.n921 B.n920 163.367
R2351 B.n917 B.n916 163.367
R2352 B.n913 B.n912 163.367
R2353 B.n909 B.n908 163.367
R2354 B.n905 B.n904 163.367
R2355 B.n901 B.n900 163.367
R2356 B.n897 B.n896 163.367
R2357 B.n893 B.n892 163.367
R2358 B.n889 B.n888 163.367
R2359 B.n885 B.n884 163.367
R2360 B.n881 B.n880 163.367
R2361 B.n877 B.n876 163.367
R2362 B.n873 B.n872 163.367
R2363 B.n869 B.n868 163.367
R2364 B.n865 B.n864 163.367
R2365 B.n861 B.n860 163.367
R2366 B.n857 B.n856 163.367
R2367 B.n853 B.n852 163.367
R2368 B.n849 B.n848 163.367
R2369 B.n845 B.n844 163.367
R2370 B.n841 B.n840 163.367
R2371 B.n837 B.n836 163.367
R2372 B.n833 B.n832 163.367
R2373 B.n829 B.n828 163.367
R2374 B.n825 B.n824 163.367
R2375 B.n821 B.n820 163.367
R2376 B.n816 B.n815 163.367
R2377 B.n812 B.n811 163.367
R2378 B.n808 B.n807 163.367
R2379 B.n804 B.n803 163.367
R2380 B.n800 B.n799 163.367
R2381 B.n796 B.n795 163.367
R2382 B.n792 B.n791 163.367
R2383 B.n788 B.n787 163.367
R2384 B.n784 B.n783 163.367
R2385 B.n780 B.n779 163.367
R2386 B.n776 B.n775 163.367
R2387 B.n772 B.n771 163.367
R2388 B.n768 B.n767 163.367
R2389 B.n764 B.n763 163.367
R2390 B.n760 B.n759 163.367
R2391 B.n756 B.n755 163.367
R2392 B.n752 B.n751 163.367
R2393 B.n748 B.n747 163.367
R2394 B.n744 B.n743 163.367
R2395 B.n740 B.n739 163.367
R2396 B.n736 B.n735 163.367
R2397 B.n732 B.n731 163.367
R2398 B.n728 B.n727 163.367
R2399 B.n724 B.n723 163.367
R2400 B.n720 B.n719 163.367
R2401 B.n716 B.n715 163.367
R2402 B.n712 B.n711 163.367
R2403 B.n708 B.n707 163.367
R2404 B.n704 B.n703 163.367
R2405 B.n700 B.n699 163.367
R2406 B.n696 B.n695 163.367
R2407 B.n692 B.n691 163.367
R2408 B.n688 B.n687 163.367
R2409 B.n684 B.n683 163.367
R2410 B.n680 B.n679 163.367
R2411 B.n676 B.n675 163.367
R2412 B.n948 B.n596 163.367
R2413 B.n948 B.n590 163.367
R2414 B.n956 B.n590 163.367
R2415 B.n956 B.n588 163.367
R2416 B.n960 B.n588 163.367
R2417 B.n960 B.n582 163.367
R2418 B.n969 B.n582 163.367
R2419 B.n969 B.n580 163.367
R2420 B.n973 B.n580 163.367
R2421 B.n973 B.n575 163.367
R2422 B.n981 B.n575 163.367
R2423 B.n981 B.n573 163.367
R2424 B.n985 B.n573 163.367
R2425 B.n985 B.n567 163.367
R2426 B.n993 B.n567 163.367
R2427 B.n993 B.n565 163.367
R2428 B.n997 B.n565 163.367
R2429 B.n997 B.n559 163.367
R2430 B.n1005 B.n559 163.367
R2431 B.n1005 B.n557 163.367
R2432 B.n1009 B.n557 163.367
R2433 B.n1009 B.n551 163.367
R2434 B.n1017 B.n551 163.367
R2435 B.n1017 B.n549 163.367
R2436 B.n1021 B.n549 163.367
R2437 B.n1021 B.n543 163.367
R2438 B.n1029 B.n543 163.367
R2439 B.n1029 B.n541 163.367
R2440 B.n1033 B.n541 163.367
R2441 B.n1033 B.n535 163.367
R2442 B.n1041 B.n535 163.367
R2443 B.n1041 B.n533 163.367
R2444 B.n1045 B.n533 163.367
R2445 B.n1045 B.n527 163.367
R2446 B.n1053 B.n527 163.367
R2447 B.n1053 B.n525 163.367
R2448 B.n1057 B.n525 163.367
R2449 B.n1057 B.n519 163.367
R2450 B.n1065 B.n519 163.367
R2451 B.n1065 B.n517 163.367
R2452 B.n1069 B.n517 163.367
R2453 B.n1069 B.n511 163.367
R2454 B.n1077 B.n511 163.367
R2455 B.n1077 B.n509 163.367
R2456 B.n1081 B.n509 163.367
R2457 B.n1081 B.n503 163.367
R2458 B.n1089 B.n503 163.367
R2459 B.n1089 B.n501 163.367
R2460 B.n1093 B.n501 163.367
R2461 B.n1093 B.n495 163.367
R2462 B.n1101 B.n495 163.367
R2463 B.n1101 B.n493 163.367
R2464 B.n1105 B.n493 163.367
R2465 B.n1105 B.n487 163.367
R2466 B.n1113 B.n487 163.367
R2467 B.n1113 B.n485 163.367
R2468 B.n1117 B.n485 163.367
R2469 B.n1117 B.n479 163.367
R2470 B.n1126 B.n479 163.367
R2471 B.n1126 B.n477 163.367
R2472 B.n1130 B.n477 163.367
R2473 B.n1130 B.n472 163.367
R2474 B.n1139 B.n472 163.367
R2475 B.n1139 B.n470 163.367
R2476 B.n1143 B.n470 163.367
R2477 B.n1143 B.n3 163.367
R2478 B.n1375 B.n3 163.367
R2479 B.n1371 B.n2 163.367
R2480 B.n1371 B.n1370 163.367
R2481 B.n1370 B.n9 163.367
R2482 B.n1366 B.n9 163.367
R2483 B.n1366 B.n11 163.367
R2484 B.n1362 B.n11 163.367
R2485 B.n1362 B.n16 163.367
R2486 B.n1358 B.n16 163.367
R2487 B.n1358 B.n18 163.367
R2488 B.n1354 B.n18 163.367
R2489 B.n1354 B.n24 163.367
R2490 B.n1350 B.n24 163.367
R2491 B.n1350 B.n26 163.367
R2492 B.n1346 B.n26 163.367
R2493 B.n1346 B.n31 163.367
R2494 B.n1342 B.n31 163.367
R2495 B.n1342 B.n33 163.367
R2496 B.n1338 B.n33 163.367
R2497 B.n1338 B.n38 163.367
R2498 B.n1334 B.n38 163.367
R2499 B.n1334 B.n40 163.367
R2500 B.n1330 B.n40 163.367
R2501 B.n1330 B.n45 163.367
R2502 B.n1326 B.n45 163.367
R2503 B.n1326 B.n47 163.367
R2504 B.n1322 B.n47 163.367
R2505 B.n1322 B.n52 163.367
R2506 B.n1318 B.n52 163.367
R2507 B.n1318 B.n54 163.367
R2508 B.n1314 B.n54 163.367
R2509 B.n1314 B.n59 163.367
R2510 B.n1310 B.n59 163.367
R2511 B.n1310 B.n61 163.367
R2512 B.n1306 B.n61 163.367
R2513 B.n1306 B.n66 163.367
R2514 B.n1302 B.n66 163.367
R2515 B.n1302 B.n68 163.367
R2516 B.n1298 B.n68 163.367
R2517 B.n1298 B.n73 163.367
R2518 B.n1294 B.n73 163.367
R2519 B.n1294 B.n75 163.367
R2520 B.n1290 B.n75 163.367
R2521 B.n1290 B.n80 163.367
R2522 B.n1286 B.n80 163.367
R2523 B.n1286 B.n82 163.367
R2524 B.n1282 B.n82 163.367
R2525 B.n1282 B.n87 163.367
R2526 B.n1278 B.n87 163.367
R2527 B.n1278 B.n89 163.367
R2528 B.n1274 B.n89 163.367
R2529 B.n1274 B.n94 163.367
R2530 B.n1270 B.n94 163.367
R2531 B.n1270 B.n96 163.367
R2532 B.n1266 B.n96 163.367
R2533 B.n1266 B.n101 163.367
R2534 B.n1262 B.n101 163.367
R2535 B.n1262 B.n103 163.367
R2536 B.n1258 B.n103 163.367
R2537 B.n1258 B.n107 163.367
R2538 B.n1254 B.n107 163.367
R2539 B.n1254 B.n109 163.367
R2540 B.n1250 B.n109 163.367
R2541 B.n1250 B.n115 163.367
R2542 B.n1246 B.n115 163.367
R2543 B.n1246 B.n117 163.367
R2544 B.n1242 B.n117 163.367
R2545 B.n1242 B.n122 163.367
R2546 B.n1238 B.n1237 71.676
R2547 B.n199 B.n125 71.676
R2548 B.n203 B.n126 71.676
R2549 B.n207 B.n127 71.676
R2550 B.n211 B.n128 71.676
R2551 B.n215 B.n129 71.676
R2552 B.n219 B.n130 71.676
R2553 B.n223 B.n131 71.676
R2554 B.n227 B.n132 71.676
R2555 B.n231 B.n133 71.676
R2556 B.n235 B.n134 71.676
R2557 B.n239 B.n135 71.676
R2558 B.n243 B.n136 71.676
R2559 B.n247 B.n137 71.676
R2560 B.n251 B.n138 71.676
R2561 B.n255 B.n139 71.676
R2562 B.n259 B.n140 71.676
R2563 B.n263 B.n141 71.676
R2564 B.n267 B.n142 71.676
R2565 B.n271 B.n143 71.676
R2566 B.n275 B.n144 71.676
R2567 B.n279 B.n145 71.676
R2568 B.n283 B.n146 71.676
R2569 B.n287 B.n147 71.676
R2570 B.n291 B.n148 71.676
R2571 B.n295 B.n149 71.676
R2572 B.n299 B.n150 71.676
R2573 B.n303 B.n151 71.676
R2574 B.n307 B.n152 71.676
R2575 B.n311 B.n153 71.676
R2576 B.n315 B.n154 71.676
R2577 B.n319 B.n155 71.676
R2578 B.n323 B.n156 71.676
R2579 B.n327 B.n157 71.676
R2580 B.n331 B.n158 71.676
R2581 B.n335 B.n159 71.676
R2582 B.n339 B.n160 71.676
R2583 B.n344 B.n161 71.676
R2584 B.n348 B.n162 71.676
R2585 B.n352 B.n163 71.676
R2586 B.n356 B.n164 71.676
R2587 B.n360 B.n165 71.676
R2588 B.n364 B.n166 71.676
R2589 B.n368 B.n167 71.676
R2590 B.n372 B.n168 71.676
R2591 B.n376 B.n169 71.676
R2592 B.n380 B.n170 71.676
R2593 B.n384 B.n171 71.676
R2594 B.n388 B.n172 71.676
R2595 B.n392 B.n173 71.676
R2596 B.n396 B.n174 71.676
R2597 B.n400 B.n175 71.676
R2598 B.n404 B.n176 71.676
R2599 B.n408 B.n177 71.676
R2600 B.n412 B.n178 71.676
R2601 B.n416 B.n179 71.676
R2602 B.n420 B.n180 71.676
R2603 B.n424 B.n181 71.676
R2604 B.n428 B.n182 71.676
R2605 B.n432 B.n183 71.676
R2606 B.n436 B.n184 71.676
R2607 B.n440 B.n185 71.676
R2608 B.n444 B.n186 71.676
R2609 B.n448 B.n187 71.676
R2610 B.n452 B.n188 71.676
R2611 B.n456 B.n189 71.676
R2612 B.n460 B.n190 71.676
R2613 B.n464 B.n191 71.676
R2614 B.n192 B.n191 71.676
R2615 B.n463 B.n190 71.676
R2616 B.n459 B.n189 71.676
R2617 B.n455 B.n188 71.676
R2618 B.n451 B.n187 71.676
R2619 B.n447 B.n186 71.676
R2620 B.n443 B.n185 71.676
R2621 B.n439 B.n184 71.676
R2622 B.n435 B.n183 71.676
R2623 B.n431 B.n182 71.676
R2624 B.n427 B.n181 71.676
R2625 B.n423 B.n180 71.676
R2626 B.n419 B.n179 71.676
R2627 B.n415 B.n178 71.676
R2628 B.n411 B.n177 71.676
R2629 B.n407 B.n176 71.676
R2630 B.n403 B.n175 71.676
R2631 B.n399 B.n174 71.676
R2632 B.n395 B.n173 71.676
R2633 B.n391 B.n172 71.676
R2634 B.n387 B.n171 71.676
R2635 B.n383 B.n170 71.676
R2636 B.n379 B.n169 71.676
R2637 B.n375 B.n168 71.676
R2638 B.n371 B.n167 71.676
R2639 B.n367 B.n166 71.676
R2640 B.n363 B.n165 71.676
R2641 B.n359 B.n164 71.676
R2642 B.n355 B.n163 71.676
R2643 B.n351 B.n162 71.676
R2644 B.n347 B.n161 71.676
R2645 B.n343 B.n160 71.676
R2646 B.n338 B.n159 71.676
R2647 B.n334 B.n158 71.676
R2648 B.n330 B.n157 71.676
R2649 B.n326 B.n156 71.676
R2650 B.n322 B.n155 71.676
R2651 B.n318 B.n154 71.676
R2652 B.n314 B.n153 71.676
R2653 B.n310 B.n152 71.676
R2654 B.n306 B.n151 71.676
R2655 B.n302 B.n150 71.676
R2656 B.n298 B.n149 71.676
R2657 B.n294 B.n148 71.676
R2658 B.n290 B.n147 71.676
R2659 B.n286 B.n146 71.676
R2660 B.n282 B.n145 71.676
R2661 B.n278 B.n144 71.676
R2662 B.n274 B.n143 71.676
R2663 B.n270 B.n142 71.676
R2664 B.n266 B.n141 71.676
R2665 B.n262 B.n140 71.676
R2666 B.n258 B.n139 71.676
R2667 B.n254 B.n138 71.676
R2668 B.n250 B.n137 71.676
R2669 B.n246 B.n136 71.676
R2670 B.n242 B.n135 71.676
R2671 B.n238 B.n134 71.676
R2672 B.n234 B.n133 71.676
R2673 B.n230 B.n132 71.676
R2674 B.n226 B.n131 71.676
R2675 B.n222 B.n130 71.676
R2676 B.n218 B.n129 71.676
R2677 B.n214 B.n128 71.676
R2678 B.n210 B.n127 71.676
R2679 B.n206 B.n126 71.676
R2680 B.n202 B.n125 71.676
R2681 B.n1237 B.n124 71.676
R2682 B.n944 B.n943 71.676
R2683 B.n666 B.n599 71.676
R2684 B.n936 B.n600 71.676
R2685 B.n932 B.n601 71.676
R2686 B.n928 B.n602 71.676
R2687 B.n924 B.n603 71.676
R2688 B.n920 B.n604 71.676
R2689 B.n916 B.n605 71.676
R2690 B.n912 B.n606 71.676
R2691 B.n908 B.n607 71.676
R2692 B.n904 B.n608 71.676
R2693 B.n900 B.n609 71.676
R2694 B.n896 B.n610 71.676
R2695 B.n892 B.n611 71.676
R2696 B.n888 B.n612 71.676
R2697 B.n884 B.n613 71.676
R2698 B.n880 B.n614 71.676
R2699 B.n876 B.n615 71.676
R2700 B.n872 B.n616 71.676
R2701 B.n868 B.n617 71.676
R2702 B.n864 B.n618 71.676
R2703 B.n860 B.n619 71.676
R2704 B.n856 B.n620 71.676
R2705 B.n852 B.n621 71.676
R2706 B.n848 B.n622 71.676
R2707 B.n844 B.n623 71.676
R2708 B.n840 B.n624 71.676
R2709 B.n836 B.n625 71.676
R2710 B.n832 B.n626 71.676
R2711 B.n828 B.n627 71.676
R2712 B.n824 B.n628 71.676
R2713 B.n820 B.n629 71.676
R2714 B.n815 B.n630 71.676
R2715 B.n811 B.n631 71.676
R2716 B.n807 B.n632 71.676
R2717 B.n803 B.n633 71.676
R2718 B.n799 B.n634 71.676
R2719 B.n795 B.n635 71.676
R2720 B.n791 B.n636 71.676
R2721 B.n787 B.n637 71.676
R2722 B.n783 B.n638 71.676
R2723 B.n779 B.n639 71.676
R2724 B.n775 B.n640 71.676
R2725 B.n771 B.n641 71.676
R2726 B.n767 B.n642 71.676
R2727 B.n763 B.n643 71.676
R2728 B.n759 B.n644 71.676
R2729 B.n755 B.n645 71.676
R2730 B.n751 B.n646 71.676
R2731 B.n747 B.n647 71.676
R2732 B.n743 B.n648 71.676
R2733 B.n739 B.n649 71.676
R2734 B.n735 B.n650 71.676
R2735 B.n731 B.n651 71.676
R2736 B.n727 B.n652 71.676
R2737 B.n723 B.n653 71.676
R2738 B.n719 B.n654 71.676
R2739 B.n715 B.n655 71.676
R2740 B.n711 B.n656 71.676
R2741 B.n707 B.n657 71.676
R2742 B.n703 B.n658 71.676
R2743 B.n699 B.n659 71.676
R2744 B.n695 B.n660 71.676
R2745 B.n691 B.n661 71.676
R2746 B.n687 B.n662 71.676
R2747 B.n683 B.n663 71.676
R2748 B.n679 B.n664 71.676
R2749 B.n675 B.n665 71.676
R2750 B.n943 B.n598 71.676
R2751 B.n937 B.n599 71.676
R2752 B.n933 B.n600 71.676
R2753 B.n929 B.n601 71.676
R2754 B.n925 B.n602 71.676
R2755 B.n921 B.n603 71.676
R2756 B.n917 B.n604 71.676
R2757 B.n913 B.n605 71.676
R2758 B.n909 B.n606 71.676
R2759 B.n905 B.n607 71.676
R2760 B.n901 B.n608 71.676
R2761 B.n897 B.n609 71.676
R2762 B.n893 B.n610 71.676
R2763 B.n889 B.n611 71.676
R2764 B.n885 B.n612 71.676
R2765 B.n881 B.n613 71.676
R2766 B.n877 B.n614 71.676
R2767 B.n873 B.n615 71.676
R2768 B.n869 B.n616 71.676
R2769 B.n865 B.n617 71.676
R2770 B.n861 B.n618 71.676
R2771 B.n857 B.n619 71.676
R2772 B.n853 B.n620 71.676
R2773 B.n849 B.n621 71.676
R2774 B.n845 B.n622 71.676
R2775 B.n841 B.n623 71.676
R2776 B.n837 B.n624 71.676
R2777 B.n833 B.n625 71.676
R2778 B.n829 B.n626 71.676
R2779 B.n825 B.n627 71.676
R2780 B.n821 B.n628 71.676
R2781 B.n816 B.n629 71.676
R2782 B.n812 B.n630 71.676
R2783 B.n808 B.n631 71.676
R2784 B.n804 B.n632 71.676
R2785 B.n800 B.n633 71.676
R2786 B.n796 B.n634 71.676
R2787 B.n792 B.n635 71.676
R2788 B.n788 B.n636 71.676
R2789 B.n784 B.n637 71.676
R2790 B.n780 B.n638 71.676
R2791 B.n776 B.n639 71.676
R2792 B.n772 B.n640 71.676
R2793 B.n768 B.n641 71.676
R2794 B.n764 B.n642 71.676
R2795 B.n760 B.n643 71.676
R2796 B.n756 B.n644 71.676
R2797 B.n752 B.n645 71.676
R2798 B.n748 B.n646 71.676
R2799 B.n744 B.n647 71.676
R2800 B.n740 B.n648 71.676
R2801 B.n736 B.n649 71.676
R2802 B.n732 B.n650 71.676
R2803 B.n728 B.n651 71.676
R2804 B.n724 B.n652 71.676
R2805 B.n720 B.n653 71.676
R2806 B.n716 B.n654 71.676
R2807 B.n712 B.n655 71.676
R2808 B.n708 B.n656 71.676
R2809 B.n704 B.n657 71.676
R2810 B.n700 B.n658 71.676
R2811 B.n696 B.n659 71.676
R2812 B.n692 B.n660 71.676
R2813 B.n688 B.n661 71.676
R2814 B.n684 B.n662 71.676
R2815 B.n680 B.n663 71.676
R2816 B.n676 B.n664 71.676
R2817 B.n672 B.n665 71.676
R2818 B.n1376 B.n1375 71.676
R2819 B.n1376 B.n2 71.676
R2820 B.n197 B.n196 65.1641
R2821 B.n195 B.n194 65.1641
R2822 B.n670 B.n669 65.1641
R2823 B.n668 B.n667 65.1641
R2824 B.n198 B.n197 59.5399
R2825 B.n341 B.n195 59.5399
R2826 B.n671 B.n670 59.5399
R2827 B.n818 B.n668 59.5399
R2828 B.n942 B.n595 51.948
R2829 B.n1236 B.n121 51.948
R2830 B.n946 B.n945 31.0639
R2831 B.n673 B.n593 31.0639
R2832 B.n1234 B.n1233 31.0639
R2833 B.n1240 B.n1239 31.0639
R2834 B.n949 B.n595 30.1922
R2835 B.n949 B.n591 30.1922
R2836 B.n955 B.n591 30.1922
R2837 B.n955 B.n587 30.1922
R2838 B.n961 B.n587 30.1922
R2839 B.n961 B.n583 30.1922
R2840 B.n968 B.n583 30.1922
R2841 B.n968 B.n967 30.1922
R2842 B.n974 B.n576 30.1922
R2843 B.n980 B.n576 30.1922
R2844 B.n980 B.n572 30.1922
R2845 B.n986 B.n572 30.1922
R2846 B.n986 B.n568 30.1922
R2847 B.n992 B.n568 30.1922
R2848 B.n992 B.n564 30.1922
R2849 B.n998 B.n564 30.1922
R2850 B.n998 B.n560 30.1922
R2851 B.n1004 B.n560 30.1922
R2852 B.n1004 B.n556 30.1922
R2853 B.n1010 B.n556 30.1922
R2854 B.n1016 B.n552 30.1922
R2855 B.n1016 B.n548 30.1922
R2856 B.n1022 B.n548 30.1922
R2857 B.n1022 B.n544 30.1922
R2858 B.n1028 B.n544 30.1922
R2859 B.n1028 B.n540 30.1922
R2860 B.n1034 B.n540 30.1922
R2861 B.n1034 B.n536 30.1922
R2862 B.n1040 B.n536 30.1922
R2863 B.n1046 B.n532 30.1922
R2864 B.n1046 B.n528 30.1922
R2865 B.n1052 B.n528 30.1922
R2866 B.n1052 B.n524 30.1922
R2867 B.n1058 B.n524 30.1922
R2868 B.n1058 B.n520 30.1922
R2869 B.n1064 B.n520 30.1922
R2870 B.n1064 B.n516 30.1922
R2871 B.n1070 B.n516 30.1922
R2872 B.n1076 B.n512 30.1922
R2873 B.n1076 B.n508 30.1922
R2874 B.n1082 B.n508 30.1922
R2875 B.n1082 B.n504 30.1922
R2876 B.n1088 B.n504 30.1922
R2877 B.n1088 B.n500 30.1922
R2878 B.n1094 B.n500 30.1922
R2879 B.n1094 B.n496 30.1922
R2880 B.n1100 B.n496 30.1922
R2881 B.n1106 B.n492 30.1922
R2882 B.n1106 B.n488 30.1922
R2883 B.n1112 B.n488 30.1922
R2884 B.n1112 B.n484 30.1922
R2885 B.n1118 B.n484 30.1922
R2886 B.n1118 B.n480 30.1922
R2887 B.n1125 B.n480 30.1922
R2888 B.n1125 B.n1124 30.1922
R2889 B.n1131 B.n473 30.1922
R2890 B.n1138 B.n473 30.1922
R2891 B.n1138 B.n469 30.1922
R2892 B.n1144 B.n469 30.1922
R2893 B.n1144 B.n4 30.1922
R2894 B.n1374 B.n4 30.1922
R2895 B.n1374 B.n1373 30.1922
R2896 B.n1373 B.n1372 30.1922
R2897 B.n1372 B.n8 30.1922
R2898 B.n12 B.n8 30.1922
R2899 B.n1365 B.n12 30.1922
R2900 B.n1365 B.n1364 30.1922
R2901 B.n1364 B.n1363 30.1922
R2902 B.n1357 B.n19 30.1922
R2903 B.n1357 B.n1356 30.1922
R2904 B.n1356 B.n1355 30.1922
R2905 B.n1355 B.n23 30.1922
R2906 B.n1349 B.n23 30.1922
R2907 B.n1349 B.n1348 30.1922
R2908 B.n1348 B.n1347 30.1922
R2909 B.n1347 B.n30 30.1922
R2910 B.n1341 B.n1340 30.1922
R2911 B.n1340 B.n1339 30.1922
R2912 B.n1339 B.n37 30.1922
R2913 B.n1333 B.n37 30.1922
R2914 B.n1333 B.n1332 30.1922
R2915 B.n1332 B.n1331 30.1922
R2916 B.n1331 B.n44 30.1922
R2917 B.n1325 B.n44 30.1922
R2918 B.n1325 B.n1324 30.1922
R2919 B.n1323 B.n51 30.1922
R2920 B.n1317 B.n51 30.1922
R2921 B.n1317 B.n1316 30.1922
R2922 B.n1316 B.n1315 30.1922
R2923 B.n1315 B.n58 30.1922
R2924 B.n1309 B.n58 30.1922
R2925 B.n1309 B.n1308 30.1922
R2926 B.n1308 B.n1307 30.1922
R2927 B.n1307 B.n65 30.1922
R2928 B.n1301 B.n1300 30.1922
R2929 B.n1300 B.n1299 30.1922
R2930 B.n1299 B.n72 30.1922
R2931 B.n1293 B.n72 30.1922
R2932 B.n1293 B.n1292 30.1922
R2933 B.n1292 B.n1291 30.1922
R2934 B.n1291 B.n79 30.1922
R2935 B.n1285 B.n79 30.1922
R2936 B.n1285 B.n1284 30.1922
R2937 B.n1283 B.n86 30.1922
R2938 B.n1277 B.n86 30.1922
R2939 B.n1277 B.n1276 30.1922
R2940 B.n1276 B.n1275 30.1922
R2941 B.n1275 B.n93 30.1922
R2942 B.n1269 B.n93 30.1922
R2943 B.n1269 B.n1268 30.1922
R2944 B.n1268 B.n1267 30.1922
R2945 B.n1267 B.n100 30.1922
R2946 B.n1261 B.n100 30.1922
R2947 B.n1261 B.n1260 30.1922
R2948 B.n1260 B.n1259 30.1922
R2949 B.n1253 B.n110 30.1922
R2950 B.n1253 B.n1252 30.1922
R2951 B.n1252 B.n1251 30.1922
R2952 B.n1251 B.n114 30.1922
R2953 B.n1245 B.n114 30.1922
R2954 B.n1245 B.n1244 30.1922
R2955 B.n1244 B.n1243 30.1922
R2956 B.n1243 B.n121 30.1922
R2957 B.n1124 B.t5 28.8602
R2958 B.n19 B.t7 28.8602
R2959 B.t0 B.n492 27.9722
R2960 B.t4 B.n30 27.9722
R2961 B.t6 B.n512 24.4203
R2962 B.n1324 B.t9 24.4203
R2963 B.t8 B.n532 20.8683
R2964 B.t3 B.n65 20.8683
R2965 B.n974 B.t11 19.9803
R2966 B.n1259 B.t15 19.9803
R2967 B B.n1377 18.0485
R2968 B.t2 B.n552 17.3163
R2969 B.n1284 B.t1 17.3163
R2970 B.n1010 B.t2 12.8764
R2971 B.t1 B.n1283 12.8764
R2972 B.n947 B.n946 10.6151
R2973 B.n947 B.n589 10.6151
R2974 B.n957 B.n589 10.6151
R2975 B.n958 B.n957 10.6151
R2976 B.n959 B.n958 10.6151
R2977 B.n959 B.n581 10.6151
R2978 B.n970 B.n581 10.6151
R2979 B.n971 B.n970 10.6151
R2980 B.n972 B.n971 10.6151
R2981 B.n972 B.n574 10.6151
R2982 B.n982 B.n574 10.6151
R2983 B.n983 B.n982 10.6151
R2984 B.n984 B.n983 10.6151
R2985 B.n984 B.n566 10.6151
R2986 B.n994 B.n566 10.6151
R2987 B.n995 B.n994 10.6151
R2988 B.n996 B.n995 10.6151
R2989 B.n996 B.n558 10.6151
R2990 B.n1006 B.n558 10.6151
R2991 B.n1007 B.n1006 10.6151
R2992 B.n1008 B.n1007 10.6151
R2993 B.n1008 B.n550 10.6151
R2994 B.n1018 B.n550 10.6151
R2995 B.n1019 B.n1018 10.6151
R2996 B.n1020 B.n1019 10.6151
R2997 B.n1020 B.n542 10.6151
R2998 B.n1030 B.n542 10.6151
R2999 B.n1031 B.n1030 10.6151
R3000 B.n1032 B.n1031 10.6151
R3001 B.n1032 B.n534 10.6151
R3002 B.n1042 B.n534 10.6151
R3003 B.n1043 B.n1042 10.6151
R3004 B.n1044 B.n1043 10.6151
R3005 B.n1044 B.n526 10.6151
R3006 B.n1054 B.n526 10.6151
R3007 B.n1055 B.n1054 10.6151
R3008 B.n1056 B.n1055 10.6151
R3009 B.n1056 B.n518 10.6151
R3010 B.n1066 B.n518 10.6151
R3011 B.n1067 B.n1066 10.6151
R3012 B.n1068 B.n1067 10.6151
R3013 B.n1068 B.n510 10.6151
R3014 B.n1078 B.n510 10.6151
R3015 B.n1079 B.n1078 10.6151
R3016 B.n1080 B.n1079 10.6151
R3017 B.n1080 B.n502 10.6151
R3018 B.n1090 B.n502 10.6151
R3019 B.n1091 B.n1090 10.6151
R3020 B.n1092 B.n1091 10.6151
R3021 B.n1092 B.n494 10.6151
R3022 B.n1102 B.n494 10.6151
R3023 B.n1103 B.n1102 10.6151
R3024 B.n1104 B.n1103 10.6151
R3025 B.n1104 B.n486 10.6151
R3026 B.n1114 B.n486 10.6151
R3027 B.n1115 B.n1114 10.6151
R3028 B.n1116 B.n1115 10.6151
R3029 B.n1116 B.n478 10.6151
R3030 B.n1127 B.n478 10.6151
R3031 B.n1128 B.n1127 10.6151
R3032 B.n1129 B.n1128 10.6151
R3033 B.n1129 B.n471 10.6151
R3034 B.n1140 B.n471 10.6151
R3035 B.n1141 B.n1140 10.6151
R3036 B.n1142 B.n1141 10.6151
R3037 B.n1142 B.n0 10.6151
R3038 B.n945 B.n597 10.6151
R3039 B.n940 B.n597 10.6151
R3040 B.n940 B.n939 10.6151
R3041 B.n939 B.n938 10.6151
R3042 B.n938 B.n935 10.6151
R3043 B.n935 B.n934 10.6151
R3044 B.n934 B.n931 10.6151
R3045 B.n931 B.n930 10.6151
R3046 B.n930 B.n927 10.6151
R3047 B.n927 B.n926 10.6151
R3048 B.n926 B.n923 10.6151
R3049 B.n923 B.n922 10.6151
R3050 B.n922 B.n919 10.6151
R3051 B.n919 B.n918 10.6151
R3052 B.n918 B.n915 10.6151
R3053 B.n915 B.n914 10.6151
R3054 B.n914 B.n911 10.6151
R3055 B.n911 B.n910 10.6151
R3056 B.n910 B.n907 10.6151
R3057 B.n907 B.n906 10.6151
R3058 B.n906 B.n903 10.6151
R3059 B.n903 B.n902 10.6151
R3060 B.n902 B.n899 10.6151
R3061 B.n899 B.n898 10.6151
R3062 B.n898 B.n895 10.6151
R3063 B.n895 B.n894 10.6151
R3064 B.n894 B.n891 10.6151
R3065 B.n891 B.n890 10.6151
R3066 B.n890 B.n887 10.6151
R3067 B.n887 B.n886 10.6151
R3068 B.n886 B.n883 10.6151
R3069 B.n883 B.n882 10.6151
R3070 B.n882 B.n879 10.6151
R3071 B.n879 B.n878 10.6151
R3072 B.n878 B.n875 10.6151
R3073 B.n875 B.n874 10.6151
R3074 B.n874 B.n871 10.6151
R3075 B.n871 B.n870 10.6151
R3076 B.n870 B.n867 10.6151
R3077 B.n867 B.n866 10.6151
R3078 B.n866 B.n863 10.6151
R3079 B.n863 B.n862 10.6151
R3080 B.n862 B.n859 10.6151
R3081 B.n859 B.n858 10.6151
R3082 B.n858 B.n855 10.6151
R3083 B.n855 B.n854 10.6151
R3084 B.n854 B.n851 10.6151
R3085 B.n851 B.n850 10.6151
R3086 B.n850 B.n847 10.6151
R3087 B.n847 B.n846 10.6151
R3088 B.n846 B.n843 10.6151
R3089 B.n843 B.n842 10.6151
R3090 B.n842 B.n839 10.6151
R3091 B.n839 B.n838 10.6151
R3092 B.n838 B.n835 10.6151
R3093 B.n835 B.n834 10.6151
R3094 B.n834 B.n831 10.6151
R3095 B.n831 B.n830 10.6151
R3096 B.n830 B.n827 10.6151
R3097 B.n827 B.n826 10.6151
R3098 B.n826 B.n823 10.6151
R3099 B.n823 B.n822 10.6151
R3100 B.n822 B.n819 10.6151
R3101 B.n817 B.n814 10.6151
R3102 B.n814 B.n813 10.6151
R3103 B.n813 B.n810 10.6151
R3104 B.n810 B.n809 10.6151
R3105 B.n809 B.n806 10.6151
R3106 B.n806 B.n805 10.6151
R3107 B.n805 B.n802 10.6151
R3108 B.n802 B.n801 10.6151
R3109 B.n798 B.n797 10.6151
R3110 B.n797 B.n794 10.6151
R3111 B.n794 B.n793 10.6151
R3112 B.n793 B.n790 10.6151
R3113 B.n790 B.n789 10.6151
R3114 B.n789 B.n786 10.6151
R3115 B.n786 B.n785 10.6151
R3116 B.n785 B.n782 10.6151
R3117 B.n782 B.n781 10.6151
R3118 B.n781 B.n778 10.6151
R3119 B.n778 B.n777 10.6151
R3120 B.n777 B.n774 10.6151
R3121 B.n774 B.n773 10.6151
R3122 B.n773 B.n770 10.6151
R3123 B.n770 B.n769 10.6151
R3124 B.n769 B.n766 10.6151
R3125 B.n766 B.n765 10.6151
R3126 B.n765 B.n762 10.6151
R3127 B.n762 B.n761 10.6151
R3128 B.n761 B.n758 10.6151
R3129 B.n758 B.n757 10.6151
R3130 B.n757 B.n754 10.6151
R3131 B.n754 B.n753 10.6151
R3132 B.n753 B.n750 10.6151
R3133 B.n750 B.n749 10.6151
R3134 B.n749 B.n746 10.6151
R3135 B.n746 B.n745 10.6151
R3136 B.n745 B.n742 10.6151
R3137 B.n742 B.n741 10.6151
R3138 B.n741 B.n738 10.6151
R3139 B.n738 B.n737 10.6151
R3140 B.n737 B.n734 10.6151
R3141 B.n734 B.n733 10.6151
R3142 B.n733 B.n730 10.6151
R3143 B.n730 B.n729 10.6151
R3144 B.n729 B.n726 10.6151
R3145 B.n726 B.n725 10.6151
R3146 B.n725 B.n722 10.6151
R3147 B.n722 B.n721 10.6151
R3148 B.n721 B.n718 10.6151
R3149 B.n718 B.n717 10.6151
R3150 B.n717 B.n714 10.6151
R3151 B.n714 B.n713 10.6151
R3152 B.n713 B.n710 10.6151
R3153 B.n710 B.n709 10.6151
R3154 B.n709 B.n706 10.6151
R3155 B.n706 B.n705 10.6151
R3156 B.n705 B.n702 10.6151
R3157 B.n702 B.n701 10.6151
R3158 B.n701 B.n698 10.6151
R3159 B.n698 B.n697 10.6151
R3160 B.n697 B.n694 10.6151
R3161 B.n694 B.n693 10.6151
R3162 B.n693 B.n690 10.6151
R3163 B.n690 B.n689 10.6151
R3164 B.n689 B.n686 10.6151
R3165 B.n686 B.n685 10.6151
R3166 B.n685 B.n682 10.6151
R3167 B.n682 B.n681 10.6151
R3168 B.n681 B.n678 10.6151
R3169 B.n678 B.n677 10.6151
R3170 B.n677 B.n674 10.6151
R3171 B.n674 B.n673 10.6151
R3172 B.n951 B.n593 10.6151
R3173 B.n952 B.n951 10.6151
R3174 B.n953 B.n952 10.6151
R3175 B.n953 B.n585 10.6151
R3176 B.n963 B.n585 10.6151
R3177 B.n964 B.n963 10.6151
R3178 B.n965 B.n964 10.6151
R3179 B.n965 B.n578 10.6151
R3180 B.n976 B.n578 10.6151
R3181 B.n977 B.n976 10.6151
R3182 B.n978 B.n977 10.6151
R3183 B.n978 B.n570 10.6151
R3184 B.n988 B.n570 10.6151
R3185 B.n989 B.n988 10.6151
R3186 B.n990 B.n989 10.6151
R3187 B.n990 B.n562 10.6151
R3188 B.n1000 B.n562 10.6151
R3189 B.n1001 B.n1000 10.6151
R3190 B.n1002 B.n1001 10.6151
R3191 B.n1002 B.n554 10.6151
R3192 B.n1012 B.n554 10.6151
R3193 B.n1013 B.n1012 10.6151
R3194 B.n1014 B.n1013 10.6151
R3195 B.n1014 B.n546 10.6151
R3196 B.n1024 B.n546 10.6151
R3197 B.n1025 B.n1024 10.6151
R3198 B.n1026 B.n1025 10.6151
R3199 B.n1026 B.n538 10.6151
R3200 B.n1036 B.n538 10.6151
R3201 B.n1037 B.n1036 10.6151
R3202 B.n1038 B.n1037 10.6151
R3203 B.n1038 B.n530 10.6151
R3204 B.n1048 B.n530 10.6151
R3205 B.n1049 B.n1048 10.6151
R3206 B.n1050 B.n1049 10.6151
R3207 B.n1050 B.n522 10.6151
R3208 B.n1060 B.n522 10.6151
R3209 B.n1061 B.n1060 10.6151
R3210 B.n1062 B.n1061 10.6151
R3211 B.n1062 B.n514 10.6151
R3212 B.n1072 B.n514 10.6151
R3213 B.n1073 B.n1072 10.6151
R3214 B.n1074 B.n1073 10.6151
R3215 B.n1074 B.n506 10.6151
R3216 B.n1084 B.n506 10.6151
R3217 B.n1085 B.n1084 10.6151
R3218 B.n1086 B.n1085 10.6151
R3219 B.n1086 B.n498 10.6151
R3220 B.n1096 B.n498 10.6151
R3221 B.n1097 B.n1096 10.6151
R3222 B.n1098 B.n1097 10.6151
R3223 B.n1098 B.n490 10.6151
R3224 B.n1108 B.n490 10.6151
R3225 B.n1109 B.n1108 10.6151
R3226 B.n1110 B.n1109 10.6151
R3227 B.n1110 B.n482 10.6151
R3228 B.n1120 B.n482 10.6151
R3229 B.n1121 B.n1120 10.6151
R3230 B.n1122 B.n1121 10.6151
R3231 B.n1122 B.n475 10.6151
R3232 B.n1133 B.n475 10.6151
R3233 B.n1134 B.n1133 10.6151
R3234 B.n1136 B.n1134 10.6151
R3235 B.n1136 B.n1135 10.6151
R3236 B.n1135 B.n467 10.6151
R3237 B.n1147 B.n467 10.6151
R3238 B.n1148 B.n1147 10.6151
R3239 B.n1149 B.n1148 10.6151
R3240 B.n1150 B.n1149 10.6151
R3241 B.n1151 B.n1150 10.6151
R3242 B.n1154 B.n1151 10.6151
R3243 B.n1155 B.n1154 10.6151
R3244 B.n1156 B.n1155 10.6151
R3245 B.n1157 B.n1156 10.6151
R3246 B.n1159 B.n1157 10.6151
R3247 B.n1160 B.n1159 10.6151
R3248 B.n1161 B.n1160 10.6151
R3249 B.n1162 B.n1161 10.6151
R3250 B.n1164 B.n1162 10.6151
R3251 B.n1165 B.n1164 10.6151
R3252 B.n1166 B.n1165 10.6151
R3253 B.n1167 B.n1166 10.6151
R3254 B.n1169 B.n1167 10.6151
R3255 B.n1170 B.n1169 10.6151
R3256 B.n1171 B.n1170 10.6151
R3257 B.n1172 B.n1171 10.6151
R3258 B.n1174 B.n1172 10.6151
R3259 B.n1175 B.n1174 10.6151
R3260 B.n1176 B.n1175 10.6151
R3261 B.n1177 B.n1176 10.6151
R3262 B.n1179 B.n1177 10.6151
R3263 B.n1180 B.n1179 10.6151
R3264 B.n1181 B.n1180 10.6151
R3265 B.n1182 B.n1181 10.6151
R3266 B.n1184 B.n1182 10.6151
R3267 B.n1185 B.n1184 10.6151
R3268 B.n1186 B.n1185 10.6151
R3269 B.n1187 B.n1186 10.6151
R3270 B.n1189 B.n1187 10.6151
R3271 B.n1190 B.n1189 10.6151
R3272 B.n1191 B.n1190 10.6151
R3273 B.n1192 B.n1191 10.6151
R3274 B.n1194 B.n1192 10.6151
R3275 B.n1195 B.n1194 10.6151
R3276 B.n1196 B.n1195 10.6151
R3277 B.n1197 B.n1196 10.6151
R3278 B.n1199 B.n1197 10.6151
R3279 B.n1200 B.n1199 10.6151
R3280 B.n1201 B.n1200 10.6151
R3281 B.n1202 B.n1201 10.6151
R3282 B.n1204 B.n1202 10.6151
R3283 B.n1205 B.n1204 10.6151
R3284 B.n1206 B.n1205 10.6151
R3285 B.n1207 B.n1206 10.6151
R3286 B.n1209 B.n1207 10.6151
R3287 B.n1210 B.n1209 10.6151
R3288 B.n1211 B.n1210 10.6151
R3289 B.n1212 B.n1211 10.6151
R3290 B.n1214 B.n1212 10.6151
R3291 B.n1215 B.n1214 10.6151
R3292 B.n1216 B.n1215 10.6151
R3293 B.n1217 B.n1216 10.6151
R3294 B.n1219 B.n1217 10.6151
R3295 B.n1220 B.n1219 10.6151
R3296 B.n1221 B.n1220 10.6151
R3297 B.n1222 B.n1221 10.6151
R3298 B.n1224 B.n1222 10.6151
R3299 B.n1225 B.n1224 10.6151
R3300 B.n1226 B.n1225 10.6151
R3301 B.n1227 B.n1226 10.6151
R3302 B.n1229 B.n1227 10.6151
R3303 B.n1230 B.n1229 10.6151
R3304 B.n1231 B.n1230 10.6151
R3305 B.n1232 B.n1231 10.6151
R3306 B.n1233 B.n1232 10.6151
R3307 B.n1369 B.n1 10.6151
R3308 B.n1369 B.n1368 10.6151
R3309 B.n1368 B.n1367 10.6151
R3310 B.n1367 B.n10 10.6151
R3311 B.n1361 B.n10 10.6151
R3312 B.n1361 B.n1360 10.6151
R3313 B.n1360 B.n1359 10.6151
R3314 B.n1359 B.n17 10.6151
R3315 B.n1353 B.n17 10.6151
R3316 B.n1353 B.n1352 10.6151
R3317 B.n1352 B.n1351 10.6151
R3318 B.n1351 B.n25 10.6151
R3319 B.n1345 B.n25 10.6151
R3320 B.n1345 B.n1344 10.6151
R3321 B.n1344 B.n1343 10.6151
R3322 B.n1343 B.n32 10.6151
R3323 B.n1337 B.n32 10.6151
R3324 B.n1337 B.n1336 10.6151
R3325 B.n1336 B.n1335 10.6151
R3326 B.n1335 B.n39 10.6151
R3327 B.n1329 B.n39 10.6151
R3328 B.n1329 B.n1328 10.6151
R3329 B.n1328 B.n1327 10.6151
R3330 B.n1327 B.n46 10.6151
R3331 B.n1321 B.n46 10.6151
R3332 B.n1321 B.n1320 10.6151
R3333 B.n1320 B.n1319 10.6151
R3334 B.n1319 B.n53 10.6151
R3335 B.n1313 B.n53 10.6151
R3336 B.n1313 B.n1312 10.6151
R3337 B.n1312 B.n1311 10.6151
R3338 B.n1311 B.n60 10.6151
R3339 B.n1305 B.n60 10.6151
R3340 B.n1305 B.n1304 10.6151
R3341 B.n1304 B.n1303 10.6151
R3342 B.n1303 B.n67 10.6151
R3343 B.n1297 B.n67 10.6151
R3344 B.n1297 B.n1296 10.6151
R3345 B.n1296 B.n1295 10.6151
R3346 B.n1295 B.n74 10.6151
R3347 B.n1289 B.n74 10.6151
R3348 B.n1289 B.n1288 10.6151
R3349 B.n1288 B.n1287 10.6151
R3350 B.n1287 B.n81 10.6151
R3351 B.n1281 B.n81 10.6151
R3352 B.n1281 B.n1280 10.6151
R3353 B.n1280 B.n1279 10.6151
R3354 B.n1279 B.n88 10.6151
R3355 B.n1273 B.n88 10.6151
R3356 B.n1273 B.n1272 10.6151
R3357 B.n1272 B.n1271 10.6151
R3358 B.n1271 B.n95 10.6151
R3359 B.n1265 B.n95 10.6151
R3360 B.n1265 B.n1264 10.6151
R3361 B.n1264 B.n1263 10.6151
R3362 B.n1263 B.n102 10.6151
R3363 B.n1257 B.n102 10.6151
R3364 B.n1257 B.n1256 10.6151
R3365 B.n1256 B.n1255 10.6151
R3366 B.n1255 B.n108 10.6151
R3367 B.n1249 B.n108 10.6151
R3368 B.n1249 B.n1248 10.6151
R3369 B.n1248 B.n1247 10.6151
R3370 B.n1247 B.n116 10.6151
R3371 B.n1241 B.n116 10.6151
R3372 B.n1241 B.n1240 10.6151
R3373 B.n1239 B.n123 10.6151
R3374 B.n200 B.n123 10.6151
R3375 B.n201 B.n200 10.6151
R3376 B.n204 B.n201 10.6151
R3377 B.n205 B.n204 10.6151
R3378 B.n208 B.n205 10.6151
R3379 B.n209 B.n208 10.6151
R3380 B.n212 B.n209 10.6151
R3381 B.n213 B.n212 10.6151
R3382 B.n216 B.n213 10.6151
R3383 B.n217 B.n216 10.6151
R3384 B.n220 B.n217 10.6151
R3385 B.n221 B.n220 10.6151
R3386 B.n224 B.n221 10.6151
R3387 B.n225 B.n224 10.6151
R3388 B.n228 B.n225 10.6151
R3389 B.n229 B.n228 10.6151
R3390 B.n232 B.n229 10.6151
R3391 B.n233 B.n232 10.6151
R3392 B.n236 B.n233 10.6151
R3393 B.n237 B.n236 10.6151
R3394 B.n240 B.n237 10.6151
R3395 B.n241 B.n240 10.6151
R3396 B.n244 B.n241 10.6151
R3397 B.n245 B.n244 10.6151
R3398 B.n248 B.n245 10.6151
R3399 B.n249 B.n248 10.6151
R3400 B.n252 B.n249 10.6151
R3401 B.n253 B.n252 10.6151
R3402 B.n256 B.n253 10.6151
R3403 B.n257 B.n256 10.6151
R3404 B.n260 B.n257 10.6151
R3405 B.n261 B.n260 10.6151
R3406 B.n264 B.n261 10.6151
R3407 B.n265 B.n264 10.6151
R3408 B.n268 B.n265 10.6151
R3409 B.n269 B.n268 10.6151
R3410 B.n272 B.n269 10.6151
R3411 B.n273 B.n272 10.6151
R3412 B.n276 B.n273 10.6151
R3413 B.n277 B.n276 10.6151
R3414 B.n280 B.n277 10.6151
R3415 B.n281 B.n280 10.6151
R3416 B.n284 B.n281 10.6151
R3417 B.n285 B.n284 10.6151
R3418 B.n288 B.n285 10.6151
R3419 B.n289 B.n288 10.6151
R3420 B.n292 B.n289 10.6151
R3421 B.n293 B.n292 10.6151
R3422 B.n296 B.n293 10.6151
R3423 B.n297 B.n296 10.6151
R3424 B.n300 B.n297 10.6151
R3425 B.n301 B.n300 10.6151
R3426 B.n304 B.n301 10.6151
R3427 B.n305 B.n304 10.6151
R3428 B.n308 B.n305 10.6151
R3429 B.n309 B.n308 10.6151
R3430 B.n312 B.n309 10.6151
R3431 B.n313 B.n312 10.6151
R3432 B.n316 B.n313 10.6151
R3433 B.n317 B.n316 10.6151
R3434 B.n320 B.n317 10.6151
R3435 B.n321 B.n320 10.6151
R3436 B.n325 B.n324 10.6151
R3437 B.n328 B.n325 10.6151
R3438 B.n329 B.n328 10.6151
R3439 B.n332 B.n329 10.6151
R3440 B.n333 B.n332 10.6151
R3441 B.n336 B.n333 10.6151
R3442 B.n337 B.n336 10.6151
R3443 B.n340 B.n337 10.6151
R3444 B.n345 B.n342 10.6151
R3445 B.n346 B.n345 10.6151
R3446 B.n349 B.n346 10.6151
R3447 B.n350 B.n349 10.6151
R3448 B.n353 B.n350 10.6151
R3449 B.n354 B.n353 10.6151
R3450 B.n357 B.n354 10.6151
R3451 B.n358 B.n357 10.6151
R3452 B.n361 B.n358 10.6151
R3453 B.n362 B.n361 10.6151
R3454 B.n365 B.n362 10.6151
R3455 B.n366 B.n365 10.6151
R3456 B.n369 B.n366 10.6151
R3457 B.n370 B.n369 10.6151
R3458 B.n373 B.n370 10.6151
R3459 B.n374 B.n373 10.6151
R3460 B.n377 B.n374 10.6151
R3461 B.n378 B.n377 10.6151
R3462 B.n381 B.n378 10.6151
R3463 B.n382 B.n381 10.6151
R3464 B.n385 B.n382 10.6151
R3465 B.n386 B.n385 10.6151
R3466 B.n389 B.n386 10.6151
R3467 B.n390 B.n389 10.6151
R3468 B.n393 B.n390 10.6151
R3469 B.n394 B.n393 10.6151
R3470 B.n397 B.n394 10.6151
R3471 B.n398 B.n397 10.6151
R3472 B.n401 B.n398 10.6151
R3473 B.n402 B.n401 10.6151
R3474 B.n405 B.n402 10.6151
R3475 B.n406 B.n405 10.6151
R3476 B.n409 B.n406 10.6151
R3477 B.n410 B.n409 10.6151
R3478 B.n413 B.n410 10.6151
R3479 B.n414 B.n413 10.6151
R3480 B.n417 B.n414 10.6151
R3481 B.n418 B.n417 10.6151
R3482 B.n421 B.n418 10.6151
R3483 B.n422 B.n421 10.6151
R3484 B.n425 B.n422 10.6151
R3485 B.n426 B.n425 10.6151
R3486 B.n429 B.n426 10.6151
R3487 B.n430 B.n429 10.6151
R3488 B.n433 B.n430 10.6151
R3489 B.n434 B.n433 10.6151
R3490 B.n437 B.n434 10.6151
R3491 B.n438 B.n437 10.6151
R3492 B.n441 B.n438 10.6151
R3493 B.n442 B.n441 10.6151
R3494 B.n445 B.n442 10.6151
R3495 B.n446 B.n445 10.6151
R3496 B.n449 B.n446 10.6151
R3497 B.n450 B.n449 10.6151
R3498 B.n453 B.n450 10.6151
R3499 B.n454 B.n453 10.6151
R3500 B.n457 B.n454 10.6151
R3501 B.n458 B.n457 10.6151
R3502 B.n461 B.n458 10.6151
R3503 B.n462 B.n461 10.6151
R3504 B.n465 B.n462 10.6151
R3505 B.n466 B.n465 10.6151
R3506 B.n1234 B.n466 10.6151
R3507 B.n967 B.t11 10.2124
R3508 B.n110 B.t15 10.2124
R3509 B.n1040 B.t8 9.32442
R3510 B.n1301 B.t3 9.32442
R3511 B.n1377 B.n0 8.11757
R3512 B.n1377 B.n1 8.11757
R3513 B.n818 B.n817 6.5566
R3514 B.n801 B.n671 6.5566
R3515 B.n324 B.n198 6.5566
R3516 B.n341 B.n340 6.5566
R3517 B.n1070 B.t6 5.77245
R3518 B.t9 B.n1323 5.77245
R3519 B.n819 B.n818 4.05904
R3520 B.n798 B.n671 4.05904
R3521 B.n321 B.n198 4.05904
R3522 B.n342 B.n341 4.05904
R3523 B.n1100 B.t0 2.22048
R3524 B.n1341 B.t4 2.22048
R3525 B.n1131 B.t5 1.33249
R3526 B.n1363 B.t7 1.33249
R3527 VN.n58 VN.t7 186.941
R3528 VN.n12 VN.t3 186.941
R3529 VN.n90 VN.n89 161.3
R3530 VN.n88 VN.n47 161.3
R3531 VN.n87 VN.n86 161.3
R3532 VN.n85 VN.n48 161.3
R3533 VN.n84 VN.n83 161.3
R3534 VN.n82 VN.n49 161.3
R3535 VN.n80 VN.n79 161.3
R3536 VN.n78 VN.n50 161.3
R3537 VN.n77 VN.n76 161.3
R3538 VN.n75 VN.n51 161.3
R3539 VN.n74 VN.n73 161.3
R3540 VN.n72 VN.n52 161.3
R3541 VN.n71 VN.n70 161.3
R3542 VN.n68 VN.n53 161.3
R3543 VN.n67 VN.n66 161.3
R3544 VN.n65 VN.n54 161.3
R3545 VN.n64 VN.n63 161.3
R3546 VN.n62 VN.n55 161.3
R3547 VN.n61 VN.n60 161.3
R3548 VN.n59 VN.n56 161.3
R3549 VN.n44 VN.n43 161.3
R3550 VN.n42 VN.n1 161.3
R3551 VN.n41 VN.n40 161.3
R3552 VN.n39 VN.n2 161.3
R3553 VN.n38 VN.n37 161.3
R3554 VN.n36 VN.n3 161.3
R3555 VN.n34 VN.n33 161.3
R3556 VN.n32 VN.n4 161.3
R3557 VN.n31 VN.n30 161.3
R3558 VN.n29 VN.n5 161.3
R3559 VN.n28 VN.n27 161.3
R3560 VN.n26 VN.n6 161.3
R3561 VN.n25 VN.n24 161.3
R3562 VN.n22 VN.n7 161.3
R3563 VN.n21 VN.n20 161.3
R3564 VN.n19 VN.n8 161.3
R3565 VN.n18 VN.n17 161.3
R3566 VN.n16 VN.n9 161.3
R3567 VN.n15 VN.n14 161.3
R3568 VN.n13 VN.n10 161.3
R3569 VN.n11 VN.t9 155.1
R3570 VN.n23 VN.t6 155.1
R3571 VN.n35 VN.t0 155.1
R3572 VN.n0 VN.t4 155.1
R3573 VN.n57 VN.t8 155.1
R3574 VN.n69 VN.t5 155.1
R3575 VN.n81 VN.t1 155.1
R3576 VN.n46 VN.t2 155.1
R3577 VN.n12 VN.n11 68.6894
R3578 VN.n58 VN.n57 68.6894
R3579 VN.n45 VN.n0 67.1292
R3580 VN.n91 VN.n46 67.1292
R3581 VN VN.n91 61.4754
R3582 VN.n41 VN.n2 56.5617
R3583 VN.n87 VN.n48 56.5617
R3584 VN.n17 VN.n8 47.3584
R3585 VN.n29 VN.n28 47.3584
R3586 VN.n63 VN.n54 47.3584
R3587 VN.n75 VN.n74 47.3584
R3588 VN.n17 VN.n16 33.7956
R3589 VN.n30 VN.n29 33.7956
R3590 VN.n63 VN.n62 33.7956
R3591 VN.n76 VN.n75 33.7956
R3592 VN.n15 VN.n10 24.5923
R3593 VN.n16 VN.n15 24.5923
R3594 VN.n21 VN.n8 24.5923
R3595 VN.n22 VN.n21 24.5923
R3596 VN.n24 VN.n6 24.5923
R3597 VN.n28 VN.n6 24.5923
R3598 VN.n30 VN.n4 24.5923
R3599 VN.n34 VN.n4 24.5923
R3600 VN.n37 VN.n36 24.5923
R3601 VN.n37 VN.n2 24.5923
R3602 VN.n42 VN.n41 24.5923
R3603 VN.n43 VN.n42 24.5923
R3604 VN.n62 VN.n61 24.5923
R3605 VN.n61 VN.n56 24.5923
R3606 VN.n74 VN.n52 24.5923
R3607 VN.n70 VN.n52 24.5923
R3608 VN.n68 VN.n67 24.5923
R3609 VN.n67 VN.n54 24.5923
R3610 VN.n83 VN.n48 24.5923
R3611 VN.n83 VN.n82 24.5923
R3612 VN.n80 VN.n50 24.5923
R3613 VN.n76 VN.n50 24.5923
R3614 VN.n89 VN.n88 24.5923
R3615 VN.n88 VN.n87 24.5923
R3616 VN.n43 VN.n0 23.1168
R3617 VN.n89 VN.n46 23.1168
R3618 VN.n36 VN.n35 19.1821
R3619 VN.n82 VN.n81 19.1821
R3620 VN.n23 VN.n22 12.2964
R3621 VN.n24 VN.n23 12.2964
R3622 VN.n70 VN.n69 12.2964
R3623 VN.n69 VN.n68 12.2964
R3624 VN.n11 VN.n10 5.4107
R3625 VN.n35 VN.n34 5.4107
R3626 VN.n57 VN.n56 5.4107
R3627 VN.n81 VN.n80 5.4107
R3628 VN.n59 VN.n58 5.32101
R3629 VN.n13 VN.n12 5.32101
R3630 VN.n91 VN.n90 0.354861
R3631 VN.n45 VN.n44 0.354861
R3632 VN VN.n45 0.267071
R3633 VN.n90 VN.n47 0.189894
R3634 VN.n86 VN.n47 0.189894
R3635 VN.n86 VN.n85 0.189894
R3636 VN.n85 VN.n84 0.189894
R3637 VN.n84 VN.n49 0.189894
R3638 VN.n79 VN.n49 0.189894
R3639 VN.n79 VN.n78 0.189894
R3640 VN.n78 VN.n77 0.189894
R3641 VN.n77 VN.n51 0.189894
R3642 VN.n73 VN.n51 0.189894
R3643 VN.n73 VN.n72 0.189894
R3644 VN.n72 VN.n71 0.189894
R3645 VN.n71 VN.n53 0.189894
R3646 VN.n66 VN.n53 0.189894
R3647 VN.n66 VN.n65 0.189894
R3648 VN.n65 VN.n64 0.189894
R3649 VN.n64 VN.n55 0.189894
R3650 VN.n60 VN.n55 0.189894
R3651 VN.n60 VN.n59 0.189894
R3652 VN.n14 VN.n13 0.189894
R3653 VN.n14 VN.n9 0.189894
R3654 VN.n18 VN.n9 0.189894
R3655 VN.n19 VN.n18 0.189894
R3656 VN.n20 VN.n19 0.189894
R3657 VN.n20 VN.n7 0.189894
R3658 VN.n25 VN.n7 0.189894
R3659 VN.n26 VN.n25 0.189894
R3660 VN.n27 VN.n26 0.189894
R3661 VN.n27 VN.n5 0.189894
R3662 VN.n31 VN.n5 0.189894
R3663 VN.n32 VN.n31 0.189894
R3664 VN.n33 VN.n32 0.189894
R3665 VN.n33 VN.n3 0.189894
R3666 VN.n38 VN.n3 0.189894
R3667 VN.n39 VN.n38 0.189894
R3668 VN.n40 VN.n39 0.189894
R3669 VN.n40 VN.n1 0.189894
R3670 VN.n44 VN.n1 0.189894
R3671 VDD2.n209 VDD2.n109 214.453
R3672 VDD2.n100 VDD2.n0 214.453
R3673 VDD2.n210 VDD2.n209 185
R3674 VDD2.n208 VDD2.n207 185
R3675 VDD2.n113 VDD2.n112 185
R3676 VDD2.n202 VDD2.n201 185
R3677 VDD2.n200 VDD2.n199 185
R3678 VDD2.n117 VDD2.n116 185
R3679 VDD2.n194 VDD2.n193 185
R3680 VDD2.n192 VDD2.n191 185
R3681 VDD2.n121 VDD2.n120 185
R3682 VDD2.n186 VDD2.n185 185
R3683 VDD2.n184 VDD2.n183 185
R3684 VDD2.n125 VDD2.n124 185
R3685 VDD2.n178 VDD2.n177 185
R3686 VDD2.n176 VDD2.n175 185
R3687 VDD2.n129 VDD2.n128 185
R3688 VDD2.n170 VDD2.n169 185
R3689 VDD2.n168 VDD2.n167 185
R3690 VDD2.n166 VDD2.n132 185
R3691 VDD2.n136 VDD2.n133 185
R3692 VDD2.n161 VDD2.n160 185
R3693 VDD2.n159 VDD2.n158 185
R3694 VDD2.n138 VDD2.n137 185
R3695 VDD2.n153 VDD2.n152 185
R3696 VDD2.n151 VDD2.n150 185
R3697 VDD2.n142 VDD2.n141 185
R3698 VDD2.n145 VDD2.n144 185
R3699 VDD2.n35 VDD2.n34 185
R3700 VDD2.n32 VDD2.n31 185
R3701 VDD2.n41 VDD2.n40 185
R3702 VDD2.n43 VDD2.n42 185
R3703 VDD2.n28 VDD2.n27 185
R3704 VDD2.n49 VDD2.n48 185
R3705 VDD2.n52 VDD2.n51 185
R3706 VDD2.n50 VDD2.n24 185
R3707 VDD2.n57 VDD2.n23 185
R3708 VDD2.n59 VDD2.n58 185
R3709 VDD2.n61 VDD2.n60 185
R3710 VDD2.n20 VDD2.n19 185
R3711 VDD2.n67 VDD2.n66 185
R3712 VDD2.n69 VDD2.n68 185
R3713 VDD2.n16 VDD2.n15 185
R3714 VDD2.n75 VDD2.n74 185
R3715 VDD2.n77 VDD2.n76 185
R3716 VDD2.n12 VDD2.n11 185
R3717 VDD2.n83 VDD2.n82 185
R3718 VDD2.n85 VDD2.n84 185
R3719 VDD2.n8 VDD2.n7 185
R3720 VDD2.n91 VDD2.n90 185
R3721 VDD2.n93 VDD2.n92 185
R3722 VDD2.n4 VDD2.n3 185
R3723 VDD2.n99 VDD2.n98 185
R3724 VDD2.n101 VDD2.n100 185
R3725 VDD2.t7 VDD2.n143 149.524
R3726 VDD2.t6 VDD2.n33 149.524
R3727 VDD2.n209 VDD2.n208 104.615
R3728 VDD2.n208 VDD2.n112 104.615
R3729 VDD2.n201 VDD2.n112 104.615
R3730 VDD2.n201 VDD2.n200 104.615
R3731 VDD2.n200 VDD2.n116 104.615
R3732 VDD2.n193 VDD2.n116 104.615
R3733 VDD2.n193 VDD2.n192 104.615
R3734 VDD2.n192 VDD2.n120 104.615
R3735 VDD2.n185 VDD2.n120 104.615
R3736 VDD2.n185 VDD2.n184 104.615
R3737 VDD2.n184 VDD2.n124 104.615
R3738 VDD2.n177 VDD2.n124 104.615
R3739 VDD2.n177 VDD2.n176 104.615
R3740 VDD2.n176 VDD2.n128 104.615
R3741 VDD2.n169 VDD2.n128 104.615
R3742 VDD2.n169 VDD2.n168 104.615
R3743 VDD2.n168 VDD2.n132 104.615
R3744 VDD2.n136 VDD2.n132 104.615
R3745 VDD2.n160 VDD2.n136 104.615
R3746 VDD2.n160 VDD2.n159 104.615
R3747 VDD2.n159 VDD2.n137 104.615
R3748 VDD2.n152 VDD2.n137 104.615
R3749 VDD2.n152 VDD2.n151 104.615
R3750 VDD2.n151 VDD2.n141 104.615
R3751 VDD2.n144 VDD2.n141 104.615
R3752 VDD2.n34 VDD2.n31 104.615
R3753 VDD2.n41 VDD2.n31 104.615
R3754 VDD2.n42 VDD2.n41 104.615
R3755 VDD2.n42 VDD2.n27 104.615
R3756 VDD2.n49 VDD2.n27 104.615
R3757 VDD2.n51 VDD2.n49 104.615
R3758 VDD2.n51 VDD2.n50 104.615
R3759 VDD2.n50 VDD2.n23 104.615
R3760 VDD2.n59 VDD2.n23 104.615
R3761 VDD2.n60 VDD2.n59 104.615
R3762 VDD2.n60 VDD2.n19 104.615
R3763 VDD2.n67 VDD2.n19 104.615
R3764 VDD2.n68 VDD2.n67 104.615
R3765 VDD2.n68 VDD2.n15 104.615
R3766 VDD2.n75 VDD2.n15 104.615
R3767 VDD2.n76 VDD2.n75 104.615
R3768 VDD2.n76 VDD2.n11 104.615
R3769 VDD2.n83 VDD2.n11 104.615
R3770 VDD2.n84 VDD2.n83 104.615
R3771 VDD2.n84 VDD2.n7 104.615
R3772 VDD2.n91 VDD2.n7 104.615
R3773 VDD2.n92 VDD2.n91 104.615
R3774 VDD2.n92 VDD2.n3 104.615
R3775 VDD2.n99 VDD2.n3 104.615
R3776 VDD2.n100 VDD2.n99 104.615
R3777 VDD2.n108 VDD2.n107 65.8096
R3778 VDD2 VDD2.n217 65.8068
R3779 VDD2.n216 VDD2.n215 63.6927
R3780 VDD2.n106 VDD2.n105 63.6925
R3781 VDD2.n106 VDD2.n104 55.2516
R3782 VDD2.n214 VDD2.n108 54.2843
R3783 VDD2.n214 VDD2.n213 52.355
R3784 VDD2.n144 VDD2.t7 52.3082
R3785 VDD2.n34 VDD2.t6 52.3082
R3786 VDD2.n167 VDD2.n166 13.1884
R3787 VDD2.n58 VDD2.n57 13.1884
R3788 VDD2.n211 VDD2.n210 12.8005
R3789 VDD2.n170 VDD2.n131 12.8005
R3790 VDD2.n165 VDD2.n133 12.8005
R3791 VDD2.n56 VDD2.n24 12.8005
R3792 VDD2.n61 VDD2.n22 12.8005
R3793 VDD2.n102 VDD2.n101 12.8005
R3794 VDD2.n207 VDD2.n111 12.0247
R3795 VDD2.n171 VDD2.n129 12.0247
R3796 VDD2.n162 VDD2.n161 12.0247
R3797 VDD2.n53 VDD2.n52 12.0247
R3798 VDD2.n62 VDD2.n20 12.0247
R3799 VDD2.n98 VDD2.n2 12.0247
R3800 VDD2.n206 VDD2.n113 11.249
R3801 VDD2.n175 VDD2.n174 11.249
R3802 VDD2.n158 VDD2.n135 11.249
R3803 VDD2.n48 VDD2.n26 11.249
R3804 VDD2.n66 VDD2.n65 11.249
R3805 VDD2.n97 VDD2.n4 11.249
R3806 VDD2.n203 VDD2.n202 10.4732
R3807 VDD2.n178 VDD2.n127 10.4732
R3808 VDD2.n157 VDD2.n138 10.4732
R3809 VDD2.n47 VDD2.n28 10.4732
R3810 VDD2.n69 VDD2.n18 10.4732
R3811 VDD2.n94 VDD2.n93 10.4732
R3812 VDD2.n145 VDD2.n143 10.2747
R3813 VDD2.n35 VDD2.n33 10.2747
R3814 VDD2.n199 VDD2.n115 9.69747
R3815 VDD2.n179 VDD2.n125 9.69747
R3816 VDD2.n154 VDD2.n153 9.69747
R3817 VDD2.n44 VDD2.n43 9.69747
R3818 VDD2.n70 VDD2.n16 9.69747
R3819 VDD2.n90 VDD2.n6 9.69747
R3820 VDD2.n213 VDD2.n212 9.45567
R3821 VDD2.n104 VDD2.n103 9.45567
R3822 VDD2.n147 VDD2.n146 9.3005
R3823 VDD2.n149 VDD2.n148 9.3005
R3824 VDD2.n140 VDD2.n139 9.3005
R3825 VDD2.n155 VDD2.n154 9.3005
R3826 VDD2.n157 VDD2.n156 9.3005
R3827 VDD2.n135 VDD2.n134 9.3005
R3828 VDD2.n163 VDD2.n162 9.3005
R3829 VDD2.n165 VDD2.n164 9.3005
R3830 VDD2.n119 VDD2.n118 9.3005
R3831 VDD2.n196 VDD2.n195 9.3005
R3832 VDD2.n198 VDD2.n197 9.3005
R3833 VDD2.n115 VDD2.n114 9.3005
R3834 VDD2.n204 VDD2.n203 9.3005
R3835 VDD2.n206 VDD2.n205 9.3005
R3836 VDD2.n111 VDD2.n110 9.3005
R3837 VDD2.n212 VDD2.n211 9.3005
R3838 VDD2.n190 VDD2.n189 9.3005
R3839 VDD2.n188 VDD2.n187 9.3005
R3840 VDD2.n123 VDD2.n122 9.3005
R3841 VDD2.n182 VDD2.n181 9.3005
R3842 VDD2.n180 VDD2.n179 9.3005
R3843 VDD2.n127 VDD2.n126 9.3005
R3844 VDD2.n174 VDD2.n173 9.3005
R3845 VDD2.n172 VDD2.n171 9.3005
R3846 VDD2.n131 VDD2.n130 9.3005
R3847 VDD2.n79 VDD2.n78 9.3005
R3848 VDD2.n14 VDD2.n13 9.3005
R3849 VDD2.n73 VDD2.n72 9.3005
R3850 VDD2.n71 VDD2.n70 9.3005
R3851 VDD2.n18 VDD2.n17 9.3005
R3852 VDD2.n65 VDD2.n64 9.3005
R3853 VDD2.n63 VDD2.n62 9.3005
R3854 VDD2.n22 VDD2.n21 9.3005
R3855 VDD2.n37 VDD2.n36 9.3005
R3856 VDD2.n39 VDD2.n38 9.3005
R3857 VDD2.n30 VDD2.n29 9.3005
R3858 VDD2.n45 VDD2.n44 9.3005
R3859 VDD2.n47 VDD2.n46 9.3005
R3860 VDD2.n26 VDD2.n25 9.3005
R3861 VDD2.n54 VDD2.n53 9.3005
R3862 VDD2.n56 VDD2.n55 9.3005
R3863 VDD2.n81 VDD2.n80 9.3005
R3864 VDD2.n10 VDD2.n9 9.3005
R3865 VDD2.n87 VDD2.n86 9.3005
R3866 VDD2.n89 VDD2.n88 9.3005
R3867 VDD2.n6 VDD2.n5 9.3005
R3868 VDD2.n95 VDD2.n94 9.3005
R3869 VDD2.n97 VDD2.n96 9.3005
R3870 VDD2.n2 VDD2.n1 9.3005
R3871 VDD2.n103 VDD2.n102 9.3005
R3872 VDD2.n198 VDD2.n117 8.92171
R3873 VDD2.n183 VDD2.n182 8.92171
R3874 VDD2.n150 VDD2.n140 8.92171
R3875 VDD2.n40 VDD2.n30 8.92171
R3876 VDD2.n74 VDD2.n73 8.92171
R3877 VDD2.n89 VDD2.n8 8.92171
R3878 VDD2.n213 VDD2.n109 8.2187
R3879 VDD2.n104 VDD2.n0 8.2187
R3880 VDD2.n195 VDD2.n194 8.14595
R3881 VDD2.n186 VDD2.n123 8.14595
R3882 VDD2.n149 VDD2.n142 8.14595
R3883 VDD2.n39 VDD2.n32 8.14595
R3884 VDD2.n77 VDD2.n14 8.14595
R3885 VDD2.n86 VDD2.n85 8.14595
R3886 VDD2.n191 VDD2.n119 7.3702
R3887 VDD2.n187 VDD2.n121 7.3702
R3888 VDD2.n146 VDD2.n145 7.3702
R3889 VDD2.n36 VDD2.n35 7.3702
R3890 VDD2.n78 VDD2.n12 7.3702
R3891 VDD2.n82 VDD2.n10 7.3702
R3892 VDD2.n191 VDD2.n190 6.59444
R3893 VDD2.n190 VDD2.n121 6.59444
R3894 VDD2.n81 VDD2.n12 6.59444
R3895 VDD2.n82 VDD2.n81 6.59444
R3896 VDD2.n194 VDD2.n119 5.81868
R3897 VDD2.n187 VDD2.n186 5.81868
R3898 VDD2.n146 VDD2.n142 5.81868
R3899 VDD2.n36 VDD2.n32 5.81868
R3900 VDD2.n78 VDD2.n77 5.81868
R3901 VDD2.n85 VDD2.n10 5.81868
R3902 VDD2.n211 VDD2.n109 5.3904
R3903 VDD2.n102 VDD2.n0 5.3904
R3904 VDD2.n195 VDD2.n117 5.04292
R3905 VDD2.n183 VDD2.n123 5.04292
R3906 VDD2.n150 VDD2.n149 5.04292
R3907 VDD2.n40 VDD2.n39 5.04292
R3908 VDD2.n74 VDD2.n14 5.04292
R3909 VDD2.n86 VDD2.n8 5.04292
R3910 VDD2.n199 VDD2.n198 4.26717
R3911 VDD2.n182 VDD2.n125 4.26717
R3912 VDD2.n153 VDD2.n140 4.26717
R3913 VDD2.n43 VDD2.n30 4.26717
R3914 VDD2.n73 VDD2.n16 4.26717
R3915 VDD2.n90 VDD2.n89 4.26717
R3916 VDD2.n202 VDD2.n115 3.49141
R3917 VDD2.n179 VDD2.n178 3.49141
R3918 VDD2.n154 VDD2.n138 3.49141
R3919 VDD2.n44 VDD2.n28 3.49141
R3920 VDD2.n70 VDD2.n69 3.49141
R3921 VDD2.n93 VDD2.n6 3.49141
R3922 VDD2.n216 VDD2.n214 2.89705
R3923 VDD2.n37 VDD2.n33 2.84303
R3924 VDD2.n147 VDD2.n143 2.84303
R3925 VDD2.n203 VDD2.n113 2.71565
R3926 VDD2.n175 VDD2.n127 2.71565
R3927 VDD2.n158 VDD2.n157 2.71565
R3928 VDD2.n48 VDD2.n47 2.71565
R3929 VDD2.n66 VDD2.n18 2.71565
R3930 VDD2.n94 VDD2.n4 2.71565
R3931 VDD2.n207 VDD2.n206 1.93989
R3932 VDD2.n174 VDD2.n129 1.93989
R3933 VDD2.n161 VDD2.n135 1.93989
R3934 VDD2.n52 VDD2.n26 1.93989
R3935 VDD2.n65 VDD2.n20 1.93989
R3936 VDD2.n98 VDD2.n97 1.93989
R3937 VDD2.n210 VDD2.n111 1.16414
R3938 VDD2.n171 VDD2.n170 1.16414
R3939 VDD2.n162 VDD2.n133 1.16414
R3940 VDD2.n53 VDD2.n24 1.16414
R3941 VDD2.n62 VDD2.n61 1.16414
R3942 VDD2.n101 VDD2.n2 1.16414
R3943 VDD2.n217 VDD2.t1 1.01588
R3944 VDD2.n217 VDD2.t2 1.01588
R3945 VDD2.n215 VDD2.t8 1.01588
R3946 VDD2.n215 VDD2.t4 1.01588
R3947 VDD2.n107 VDD2.t9 1.01588
R3948 VDD2.n107 VDD2.t5 1.01588
R3949 VDD2.n105 VDD2.t0 1.01588
R3950 VDD2.n105 VDD2.t3 1.01588
R3951 VDD2 VDD2.n216 0.782828
R3952 VDD2.n108 VDD2.n106 0.669292
R3953 VDD2.n167 VDD2.n131 0.388379
R3954 VDD2.n166 VDD2.n165 0.388379
R3955 VDD2.n57 VDD2.n56 0.388379
R3956 VDD2.n58 VDD2.n22 0.388379
R3957 VDD2.n212 VDD2.n110 0.155672
R3958 VDD2.n205 VDD2.n110 0.155672
R3959 VDD2.n205 VDD2.n204 0.155672
R3960 VDD2.n204 VDD2.n114 0.155672
R3961 VDD2.n197 VDD2.n114 0.155672
R3962 VDD2.n197 VDD2.n196 0.155672
R3963 VDD2.n196 VDD2.n118 0.155672
R3964 VDD2.n189 VDD2.n118 0.155672
R3965 VDD2.n189 VDD2.n188 0.155672
R3966 VDD2.n188 VDD2.n122 0.155672
R3967 VDD2.n181 VDD2.n122 0.155672
R3968 VDD2.n181 VDD2.n180 0.155672
R3969 VDD2.n180 VDD2.n126 0.155672
R3970 VDD2.n173 VDD2.n126 0.155672
R3971 VDD2.n173 VDD2.n172 0.155672
R3972 VDD2.n172 VDD2.n130 0.155672
R3973 VDD2.n164 VDD2.n130 0.155672
R3974 VDD2.n164 VDD2.n163 0.155672
R3975 VDD2.n163 VDD2.n134 0.155672
R3976 VDD2.n156 VDD2.n134 0.155672
R3977 VDD2.n156 VDD2.n155 0.155672
R3978 VDD2.n155 VDD2.n139 0.155672
R3979 VDD2.n148 VDD2.n139 0.155672
R3980 VDD2.n148 VDD2.n147 0.155672
R3981 VDD2.n38 VDD2.n37 0.155672
R3982 VDD2.n38 VDD2.n29 0.155672
R3983 VDD2.n45 VDD2.n29 0.155672
R3984 VDD2.n46 VDD2.n45 0.155672
R3985 VDD2.n46 VDD2.n25 0.155672
R3986 VDD2.n54 VDD2.n25 0.155672
R3987 VDD2.n55 VDD2.n54 0.155672
R3988 VDD2.n55 VDD2.n21 0.155672
R3989 VDD2.n63 VDD2.n21 0.155672
R3990 VDD2.n64 VDD2.n63 0.155672
R3991 VDD2.n64 VDD2.n17 0.155672
R3992 VDD2.n71 VDD2.n17 0.155672
R3993 VDD2.n72 VDD2.n71 0.155672
R3994 VDD2.n72 VDD2.n13 0.155672
R3995 VDD2.n79 VDD2.n13 0.155672
R3996 VDD2.n80 VDD2.n79 0.155672
R3997 VDD2.n80 VDD2.n9 0.155672
R3998 VDD2.n87 VDD2.n9 0.155672
R3999 VDD2.n88 VDD2.n87 0.155672
R4000 VDD2.n88 VDD2.n5 0.155672
R4001 VDD2.n95 VDD2.n5 0.155672
R4002 VDD2.n96 VDD2.n95 0.155672
R4003 VDD2.n96 VDD2.n1 0.155672
R4004 VDD2.n103 VDD2.n1 0.155672
C0 VDD2 VN 17.5086f
C1 VN VTAIL 17.9947f
C2 VDD2 VTAIL 13.8031f
C3 VN VP 10.413401f
C4 VDD2 VP 0.639288f
C5 VN VDD1 0.154666f
C6 VDD2 VDD1 2.45511f
C7 VTAIL VP 18.008999f
C8 VTAIL VDD1 13.7504f
C9 VDD1 VP 17.9882f
C10 VDD2 B 9.011057f
C11 VDD1 B 9.005048f
C12 VTAIL B 11.565416f
C13 VN B 20.78899f
C14 VP B 19.248999f
C15 VDD2.n0 B 0.032482f
C16 VDD2.n1 B 0.023447f
C17 VDD2.n2 B 0.012599f
C18 VDD2.n3 B 0.02978f
C19 VDD2.n4 B 0.013341f
C20 VDD2.n5 B 0.023447f
C21 VDD2.n6 B 0.012599f
C22 VDD2.n7 B 0.02978f
C23 VDD2.n8 B 0.013341f
C24 VDD2.n9 B 0.023447f
C25 VDD2.n10 B 0.012599f
C26 VDD2.n11 B 0.02978f
C27 VDD2.n12 B 0.013341f
C28 VDD2.n13 B 0.023447f
C29 VDD2.n14 B 0.012599f
C30 VDD2.n15 B 0.02978f
C31 VDD2.n16 B 0.013341f
C32 VDD2.n17 B 0.023447f
C33 VDD2.n18 B 0.012599f
C34 VDD2.n19 B 0.02978f
C35 VDD2.n20 B 0.013341f
C36 VDD2.n21 B 0.023447f
C37 VDD2.n22 B 0.012599f
C38 VDD2.n23 B 0.02978f
C39 VDD2.n24 B 0.013341f
C40 VDD2.n25 B 0.023447f
C41 VDD2.n26 B 0.012599f
C42 VDD2.n27 B 0.02978f
C43 VDD2.n28 B 0.013341f
C44 VDD2.n29 B 0.023447f
C45 VDD2.n30 B 0.012599f
C46 VDD2.n31 B 0.02978f
C47 VDD2.n32 B 0.013341f
C48 VDD2.n33 B 0.236563f
C49 VDD2.t6 B 0.051244f
C50 VDD2.n34 B 0.022335f
C51 VDD2.n35 B 0.021052f
C52 VDD2.n36 B 0.012599f
C53 VDD2.n37 B 1.96503f
C54 VDD2.n38 B 0.023447f
C55 VDD2.n39 B 0.012599f
C56 VDD2.n40 B 0.013341f
C57 VDD2.n41 B 0.02978f
C58 VDD2.n42 B 0.02978f
C59 VDD2.n43 B 0.013341f
C60 VDD2.n44 B 0.012599f
C61 VDD2.n45 B 0.023447f
C62 VDD2.n46 B 0.023447f
C63 VDD2.n47 B 0.012599f
C64 VDD2.n48 B 0.013341f
C65 VDD2.n49 B 0.02978f
C66 VDD2.n50 B 0.02978f
C67 VDD2.n51 B 0.02978f
C68 VDD2.n52 B 0.013341f
C69 VDD2.n53 B 0.012599f
C70 VDD2.n54 B 0.023447f
C71 VDD2.n55 B 0.023447f
C72 VDD2.n56 B 0.012599f
C73 VDD2.n57 B 0.01297f
C74 VDD2.n58 B 0.01297f
C75 VDD2.n59 B 0.02978f
C76 VDD2.n60 B 0.02978f
C77 VDD2.n61 B 0.013341f
C78 VDD2.n62 B 0.012599f
C79 VDD2.n63 B 0.023447f
C80 VDD2.n64 B 0.023447f
C81 VDD2.n65 B 0.012599f
C82 VDD2.n66 B 0.013341f
C83 VDD2.n67 B 0.02978f
C84 VDD2.n68 B 0.02978f
C85 VDD2.n69 B 0.013341f
C86 VDD2.n70 B 0.012599f
C87 VDD2.n71 B 0.023447f
C88 VDD2.n72 B 0.023447f
C89 VDD2.n73 B 0.012599f
C90 VDD2.n74 B 0.013341f
C91 VDD2.n75 B 0.02978f
C92 VDD2.n76 B 0.02978f
C93 VDD2.n77 B 0.013341f
C94 VDD2.n78 B 0.012599f
C95 VDD2.n79 B 0.023447f
C96 VDD2.n80 B 0.023447f
C97 VDD2.n81 B 0.012599f
C98 VDD2.n82 B 0.013341f
C99 VDD2.n83 B 0.02978f
C100 VDD2.n84 B 0.02978f
C101 VDD2.n85 B 0.013341f
C102 VDD2.n86 B 0.012599f
C103 VDD2.n87 B 0.023447f
C104 VDD2.n88 B 0.023447f
C105 VDD2.n89 B 0.012599f
C106 VDD2.n90 B 0.013341f
C107 VDD2.n91 B 0.02978f
C108 VDD2.n92 B 0.02978f
C109 VDD2.n93 B 0.013341f
C110 VDD2.n94 B 0.012599f
C111 VDD2.n95 B 0.023447f
C112 VDD2.n96 B 0.023447f
C113 VDD2.n97 B 0.012599f
C114 VDD2.n98 B 0.013341f
C115 VDD2.n99 B 0.02978f
C116 VDD2.n100 B 0.061367f
C117 VDD2.n101 B 0.013341f
C118 VDD2.n102 B 0.024636f
C119 VDD2.n103 B 0.059962f
C120 VDD2.n104 B 0.094093f
C121 VDD2.t0 B 0.361306f
C122 VDD2.t3 B 0.361306f
C123 VDD2.n105 B 3.30993f
C124 VDD2.n106 B 0.711073f
C125 VDD2.t9 B 0.361306f
C126 VDD2.t5 B 0.361306f
C127 VDD2.n107 B 3.32846f
C128 VDD2.n108 B 3.37307f
C129 VDD2.n109 B 0.032482f
C130 VDD2.n110 B 0.023447f
C131 VDD2.n111 B 0.012599f
C132 VDD2.n112 B 0.02978f
C133 VDD2.n113 B 0.013341f
C134 VDD2.n114 B 0.023447f
C135 VDD2.n115 B 0.012599f
C136 VDD2.n116 B 0.02978f
C137 VDD2.n117 B 0.013341f
C138 VDD2.n118 B 0.023447f
C139 VDD2.n119 B 0.012599f
C140 VDD2.n120 B 0.02978f
C141 VDD2.n121 B 0.013341f
C142 VDD2.n122 B 0.023447f
C143 VDD2.n123 B 0.012599f
C144 VDD2.n124 B 0.02978f
C145 VDD2.n125 B 0.013341f
C146 VDD2.n126 B 0.023447f
C147 VDD2.n127 B 0.012599f
C148 VDD2.n128 B 0.02978f
C149 VDD2.n129 B 0.013341f
C150 VDD2.n130 B 0.023447f
C151 VDD2.n131 B 0.012599f
C152 VDD2.n132 B 0.02978f
C153 VDD2.n133 B 0.013341f
C154 VDD2.n134 B 0.023447f
C155 VDD2.n135 B 0.012599f
C156 VDD2.n136 B 0.02978f
C157 VDD2.n137 B 0.02978f
C158 VDD2.n138 B 0.013341f
C159 VDD2.n139 B 0.023447f
C160 VDD2.n140 B 0.012599f
C161 VDD2.n141 B 0.02978f
C162 VDD2.n142 B 0.013341f
C163 VDD2.n143 B 0.236563f
C164 VDD2.t7 B 0.051244f
C165 VDD2.n144 B 0.022335f
C166 VDD2.n145 B 0.021052f
C167 VDD2.n146 B 0.012599f
C168 VDD2.n147 B 1.96503f
C169 VDD2.n148 B 0.023447f
C170 VDD2.n149 B 0.012599f
C171 VDD2.n150 B 0.013341f
C172 VDD2.n151 B 0.02978f
C173 VDD2.n152 B 0.02978f
C174 VDD2.n153 B 0.013341f
C175 VDD2.n154 B 0.012599f
C176 VDD2.n155 B 0.023447f
C177 VDD2.n156 B 0.023447f
C178 VDD2.n157 B 0.012599f
C179 VDD2.n158 B 0.013341f
C180 VDD2.n159 B 0.02978f
C181 VDD2.n160 B 0.02978f
C182 VDD2.n161 B 0.013341f
C183 VDD2.n162 B 0.012599f
C184 VDD2.n163 B 0.023447f
C185 VDD2.n164 B 0.023447f
C186 VDD2.n165 B 0.012599f
C187 VDD2.n166 B 0.01297f
C188 VDD2.n167 B 0.01297f
C189 VDD2.n168 B 0.02978f
C190 VDD2.n169 B 0.02978f
C191 VDD2.n170 B 0.013341f
C192 VDD2.n171 B 0.012599f
C193 VDD2.n172 B 0.023447f
C194 VDD2.n173 B 0.023447f
C195 VDD2.n174 B 0.012599f
C196 VDD2.n175 B 0.013341f
C197 VDD2.n176 B 0.02978f
C198 VDD2.n177 B 0.02978f
C199 VDD2.n178 B 0.013341f
C200 VDD2.n179 B 0.012599f
C201 VDD2.n180 B 0.023447f
C202 VDD2.n181 B 0.023447f
C203 VDD2.n182 B 0.012599f
C204 VDD2.n183 B 0.013341f
C205 VDD2.n184 B 0.02978f
C206 VDD2.n185 B 0.02978f
C207 VDD2.n186 B 0.013341f
C208 VDD2.n187 B 0.012599f
C209 VDD2.n188 B 0.023447f
C210 VDD2.n189 B 0.023447f
C211 VDD2.n190 B 0.012599f
C212 VDD2.n191 B 0.013341f
C213 VDD2.n192 B 0.02978f
C214 VDD2.n193 B 0.02978f
C215 VDD2.n194 B 0.013341f
C216 VDD2.n195 B 0.012599f
C217 VDD2.n196 B 0.023447f
C218 VDD2.n197 B 0.023447f
C219 VDD2.n198 B 0.012599f
C220 VDD2.n199 B 0.013341f
C221 VDD2.n200 B 0.02978f
C222 VDD2.n201 B 0.02978f
C223 VDD2.n202 B 0.013341f
C224 VDD2.n203 B 0.012599f
C225 VDD2.n204 B 0.023447f
C226 VDD2.n205 B 0.023447f
C227 VDD2.n206 B 0.012599f
C228 VDD2.n207 B 0.013341f
C229 VDD2.n208 B 0.02978f
C230 VDD2.n209 B 0.061367f
C231 VDD2.n210 B 0.013341f
C232 VDD2.n211 B 0.024636f
C233 VDD2.n212 B 0.059962f
C234 VDD2.n213 B 0.08008f
C235 VDD2.n214 B 3.40528f
C236 VDD2.t8 B 0.361306f
C237 VDD2.t4 B 0.361306f
C238 VDD2.n215 B 3.30994f
C239 VDD2.n216 B 0.465551f
C240 VDD2.t1 B 0.361306f
C241 VDD2.t2 B 0.361306f
C242 VDD2.n217 B 3.32842f
C243 VN.t4 B 2.98332f
C244 VN.n0 B 1.10508f
C245 VN.n1 B 0.01833f
C246 VN.n2 B 0.028675f
C247 VN.n3 B 0.01833f
C248 VN.t0 B 2.98332f
C249 VN.n4 B 0.033992f
C250 VN.n5 B 0.01833f
C251 VN.n6 B 0.033992f
C252 VN.n7 B 0.01833f
C253 VN.t6 B 2.98332f
C254 VN.n8 B 0.034476f
C255 VN.n9 B 0.01833f
C256 VN.n10 B 0.020903f
C257 VN.t9 B 2.98332f
C258 VN.n11 B 1.08237f
C259 VN.t3 B 3.17985f
C260 VN.n12 B 1.05557f
C261 VN.n13 B 0.19772f
C262 VN.n14 B 0.01833f
C263 VN.n15 B 0.033992f
C264 VN.n16 B 0.036825f
C265 VN.n17 B 0.015983f
C266 VN.n18 B 0.01833f
C267 VN.n19 B 0.01833f
C268 VN.n20 B 0.01833f
C269 VN.n21 B 0.033992f
C270 VN.n22 B 0.025601f
C271 VN.n23 B 1.02852f
C272 VN.n24 B 0.025601f
C273 VN.n25 B 0.01833f
C274 VN.n26 B 0.01833f
C275 VN.n27 B 0.01833f
C276 VN.n28 B 0.034476f
C277 VN.n29 B 0.015983f
C278 VN.n30 B 0.036825f
C279 VN.n31 B 0.01833f
C280 VN.n32 B 0.01833f
C281 VN.n33 B 0.01833f
C282 VN.n34 B 0.020903f
C283 VN.n35 B 1.02852f
C284 VN.n36 B 0.0303f
C285 VN.n37 B 0.033992f
C286 VN.n38 B 0.01833f
C287 VN.n39 B 0.01833f
C288 VN.n40 B 0.01833f
C289 VN.n41 B 0.024617f
C290 VN.n42 B 0.033992f
C291 VN.n43 B 0.032985f
C292 VN.n44 B 0.02958f
C293 VN.n45 B 0.035616f
C294 VN.t2 B 2.98332f
C295 VN.n46 B 1.10508f
C296 VN.n47 B 0.01833f
C297 VN.n48 B 0.028675f
C298 VN.n49 B 0.01833f
C299 VN.t1 B 2.98332f
C300 VN.n50 B 0.033992f
C301 VN.n51 B 0.01833f
C302 VN.n52 B 0.033992f
C303 VN.n53 B 0.01833f
C304 VN.t5 B 2.98332f
C305 VN.n54 B 0.034476f
C306 VN.n55 B 0.01833f
C307 VN.n56 B 0.020903f
C308 VN.t7 B 3.17985f
C309 VN.t8 B 2.98332f
C310 VN.n57 B 1.08237f
C311 VN.n58 B 1.05557f
C312 VN.n59 B 0.19772f
C313 VN.n60 B 0.01833f
C314 VN.n61 B 0.033992f
C315 VN.n62 B 0.036825f
C316 VN.n63 B 0.015983f
C317 VN.n64 B 0.01833f
C318 VN.n65 B 0.01833f
C319 VN.n66 B 0.01833f
C320 VN.n67 B 0.033992f
C321 VN.n68 B 0.025601f
C322 VN.n69 B 1.02852f
C323 VN.n70 B 0.025601f
C324 VN.n71 B 0.01833f
C325 VN.n72 B 0.01833f
C326 VN.n73 B 0.01833f
C327 VN.n74 B 0.034476f
C328 VN.n75 B 0.015983f
C329 VN.n76 B 0.036825f
C330 VN.n77 B 0.01833f
C331 VN.n78 B 0.01833f
C332 VN.n79 B 0.01833f
C333 VN.n80 B 0.020903f
C334 VN.n81 B 1.02852f
C335 VN.n82 B 0.0303f
C336 VN.n83 B 0.033992f
C337 VN.n84 B 0.01833f
C338 VN.n85 B 0.01833f
C339 VN.n86 B 0.01833f
C340 VN.n87 B 0.024617f
C341 VN.n88 B 0.033992f
C342 VN.n89 B 0.032985f
C343 VN.n90 B 0.02958f
C344 VN.n91 B 1.3802f
C345 VDD1.n0 B 0.032878f
C346 VDD1.n1 B 0.023733f
C347 VDD1.n2 B 0.012753f
C348 VDD1.n3 B 0.030144f
C349 VDD1.n4 B 0.013503f
C350 VDD1.n5 B 0.023733f
C351 VDD1.n6 B 0.012753f
C352 VDD1.n7 B 0.030144f
C353 VDD1.n8 B 0.013503f
C354 VDD1.n9 B 0.023733f
C355 VDD1.n10 B 0.012753f
C356 VDD1.n11 B 0.030144f
C357 VDD1.n12 B 0.013503f
C358 VDD1.n13 B 0.023733f
C359 VDD1.n14 B 0.012753f
C360 VDD1.n15 B 0.030144f
C361 VDD1.n16 B 0.013503f
C362 VDD1.n17 B 0.023733f
C363 VDD1.n18 B 0.012753f
C364 VDD1.n19 B 0.030144f
C365 VDD1.n20 B 0.013503f
C366 VDD1.n21 B 0.023733f
C367 VDD1.n22 B 0.012753f
C368 VDD1.n23 B 0.030144f
C369 VDD1.n24 B 0.013503f
C370 VDD1.n25 B 0.023733f
C371 VDD1.n26 B 0.012753f
C372 VDD1.n27 B 0.030144f
C373 VDD1.n28 B 0.030144f
C374 VDD1.n29 B 0.013503f
C375 VDD1.n30 B 0.023733f
C376 VDD1.n31 B 0.012753f
C377 VDD1.n32 B 0.030144f
C378 VDD1.n33 B 0.013503f
C379 VDD1.n34 B 0.239449f
C380 VDD1.t2 B 0.051869f
C381 VDD1.n35 B 0.022608f
C382 VDD1.n36 B 0.021309f
C383 VDD1.n37 B 0.012753f
C384 VDD1.n38 B 1.989f
C385 VDD1.n39 B 0.023733f
C386 VDD1.n40 B 0.012753f
C387 VDD1.n41 B 0.013503f
C388 VDD1.n42 B 0.030144f
C389 VDD1.n43 B 0.030144f
C390 VDD1.n44 B 0.013503f
C391 VDD1.n45 B 0.012753f
C392 VDD1.n46 B 0.023733f
C393 VDD1.n47 B 0.023733f
C394 VDD1.n48 B 0.012753f
C395 VDD1.n49 B 0.013503f
C396 VDD1.n50 B 0.030144f
C397 VDD1.n51 B 0.030144f
C398 VDD1.n52 B 0.013503f
C399 VDD1.n53 B 0.012753f
C400 VDD1.n54 B 0.023733f
C401 VDD1.n55 B 0.023733f
C402 VDD1.n56 B 0.012753f
C403 VDD1.n57 B 0.013128f
C404 VDD1.n58 B 0.013128f
C405 VDD1.n59 B 0.030144f
C406 VDD1.n60 B 0.030144f
C407 VDD1.n61 B 0.013503f
C408 VDD1.n62 B 0.012753f
C409 VDD1.n63 B 0.023733f
C410 VDD1.n64 B 0.023733f
C411 VDD1.n65 B 0.012753f
C412 VDD1.n66 B 0.013503f
C413 VDD1.n67 B 0.030144f
C414 VDD1.n68 B 0.030144f
C415 VDD1.n69 B 0.013503f
C416 VDD1.n70 B 0.012753f
C417 VDD1.n71 B 0.023733f
C418 VDD1.n72 B 0.023733f
C419 VDD1.n73 B 0.012753f
C420 VDD1.n74 B 0.013503f
C421 VDD1.n75 B 0.030144f
C422 VDD1.n76 B 0.030144f
C423 VDD1.n77 B 0.013503f
C424 VDD1.n78 B 0.012753f
C425 VDD1.n79 B 0.023733f
C426 VDD1.n80 B 0.023733f
C427 VDD1.n81 B 0.012753f
C428 VDD1.n82 B 0.013503f
C429 VDD1.n83 B 0.030144f
C430 VDD1.n84 B 0.030144f
C431 VDD1.n85 B 0.013503f
C432 VDD1.n86 B 0.012753f
C433 VDD1.n87 B 0.023733f
C434 VDD1.n88 B 0.023733f
C435 VDD1.n89 B 0.012753f
C436 VDD1.n90 B 0.013503f
C437 VDD1.n91 B 0.030144f
C438 VDD1.n92 B 0.030144f
C439 VDD1.n93 B 0.013503f
C440 VDD1.n94 B 0.012753f
C441 VDD1.n95 B 0.023733f
C442 VDD1.n96 B 0.023733f
C443 VDD1.n97 B 0.012753f
C444 VDD1.n98 B 0.013503f
C445 VDD1.n99 B 0.030144f
C446 VDD1.n100 B 0.062116f
C447 VDD1.n101 B 0.013503f
C448 VDD1.n102 B 0.024937f
C449 VDD1.n103 B 0.060694f
C450 VDD1.n104 B 0.095241f
C451 VDD1.t3 B 0.365714f
C452 VDD1.t7 B 0.365714f
C453 VDD1.n105 B 3.35032f
C454 VDD1.n106 B 0.727598f
C455 VDD1.n107 B 0.032878f
C456 VDD1.n108 B 0.023733f
C457 VDD1.n109 B 0.012753f
C458 VDD1.n110 B 0.030144f
C459 VDD1.n111 B 0.013503f
C460 VDD1.n112 B 0.023733f
C461 VDD1.n113 B 0.012753f
C462 VDD1.n114 B 0.030144f
C463 VDD1.n115 B 0.013503f
C464 VDD1.n116 B 0.023733f
C465 VDD1.n117 B 0.012753f
C466 VDD1.n118 B 0.030144f
C467 VDD1.n119 B 0.013503f
C468 VDD1.n120 B 0.023733f
C469 VDD1.n121 B 0.012753f
C470 VDD1.n122 B 0.030144f
C471 VDD1.n123 B 0.013503f
C472 VDD1.n124 B 0.023733f
C473 VDD1.n125 B 0.012753f
C474 VDD1.n126 B 0.030144f
C475 VDD1.n127 B 0.013503f
C476 VDD1.n128 B 0.023733f
C477 VDD1.n129 B 0.012753f
C478 VDD1.n130 B 0.030144f
C479 VDD1.n131 B 0.013503f
C480 VDD1.n132 B 0.023733f
C481 VDD1.n133 B 0.012753f
C482 VDD1.n134 B 0.030144f
C483 VDD1.n135 B 0.013503f
C484 VDD1.n136 B 0.023733f
C485 VDD1.n137 B 0.012753f
C486 VDD1.n138 B 0.030144f
C487 VDD1.n139 B 0.013503f
C488 VDD1.n140 B 0.239449f
C489 VDD1.t4 B 0.051869f
C490 VDD1.n141 B 0.022608f
C491 VDD1.n142 B 0.021309f
C492 VDD1.n143 B 0.012753f
C493 VDD1.n144 B 1.989f
C494 VDD1.n145 B 0.023733f
C495 VDD1.n146 B 0.012753f
C496 VDD1.n147 B 0.013503f
C497 VDD1.n148 B 0.030144f
C498 VDD1.n149 B 0.030144f
C499 VDD1.n150 B 0.013503f
C500 VDD1.n151 B 0.012753f
C501 VDD1.n152 B 0.023733f
C502 VDD1.n153 B 0.023733f
C503 VDD1.n154 B 0.012753f
C504 VDD1.n155 B 0.013503f
C505 VDD1.n156 B 0.030144f
C506 VDD1.n157 B 0.030144f
C507 VDD1.n158 B 0.030144f
C508 VDD1.n159 B 0.013503f
C509 VDD1.n160 B 0.012753f
C510 VDD1.n161 B 0.023733f
C511 VDD1.n162 B 0.023733f
C512 VDD1.n163 B 0.012753f
C513 VDD1.n164 B 0.013128f
C514 VDD1.n165 B 0.013128f
C515 VDD1.n166 B 0.030144f
C516 VDD1.n167 B 0.030144f
C517 VDD1.n168 B 0.013503f
C518 VDD1.n169 B 0.012753f
C519 VDD1.n170 B 0.023733f
C520 VDD1.n171 B 0.023733f
C521 VDD1.n172 B 0.012753f
C522 VDD1.n173 B 0.013503f
C523 VDD1.n174 B 0.030144f
C524 VDD1.n175 B 0.030144f
C525 VDD1.n176 B 0.013503f
C526 VDD1.n177 B 0.012753f
C527 VDD1.n178 B 0.023733f
C528 VDD1.n179 B 0.023733f
C529 VDD1.n180 B 0.012753f
C530 VDD1.n181 B 0.013503f
C531 VDD1.n182 B 0.030144f
C532 VDD1.n183 B 0.030144f
C533 VDD1.n184 B 0.013503f
C534 VDD1.n185 B 0.012753f
C535 VDD1.n186 B 0.023733f
C536 VDD1.n187 B 0.023733f
C537 VDD1.n188 B 0.012753f
C538 VDD1.n189 B 0.013503f
C539 VDD1.n190 B 0.030144f
C540 VDD1.n191 B 0.030144f
C541 VDD1.n192 B 0.013503f
C542 VDD1.n193 B 0.012753f
C543 VDD1.n194 B 0.023733f
C544 VDD1.n195 B 0.023733f
C545 VDD1.n196 B 0.012753f
C546 VDD1.n197 B 0.013503f
C547 VDD1.n198 B 0.030144f
C548 VDD1.n199 B 0.030144f
C549 VDD1.n200 B 0.013503f
C550 VDD1.n201 B 0.012753f
C551 VDD1.n202 B 0.023733f
C552 VDD1.n203 B 0.023733f
C553 VDD1.n204 B 0.012753f
C554 VDD1.n205 B 0.013503f
C555 VDD1.n206 B 0.030144f
C556 VDD1.n207 B 0.062116f
C557 VDD1.n208 B 0.013503f
C558 VDD1.n209 B 0.024937f
C559 VDD1.n210 B 0.060694f
C560 VDD1.n211 B 0.095241f
C561 VDD1.t8 B 0.365714f
C562 VDD1.t1 B 0.365714f
C563 VDD1.n212 B 3.35031f
C564 VDD1.n213 B 0.719748f
C565 VDD1.t0 B 0.365714f
C566 VDD1.t5 B 0.365714f
C567 VDD1.n214 B 3.36907f
C568 VDD1.n215 B 3.54845f
C569 VDD1.t6 B 0.365714f
C570 VDD1.t9 B 0.365714f
C571 VDD1.n216 B 3.35031f
C572 VDD1.n217 B 3.71235f
C573 VTAIL.t7 B 0.364407f
C574 VTAIL.t4 B 0.364407f
C575 VTAIL.n0 B 3.2728f
C576 VTAIL.n1 B 0.538749f
C577 VTAIL.n2 B 0.032761f
C578 VTAIL.n3 B 0.023648f
C579 VTAIL.n4 B 0.012707f
C580 VTAIL.n5 B 0.030036f
C581 VTAIL.n6 B 0.013455f
C582 VTAIL.n7 B 0.023648f
C583 VTAIL.n8 B 0.012707f
C584 VTAIL.n9 B 0.030036f
C585 VTAIL.n10 B 0.013455f
C586 VTAIL.n11 B 0.023648f
C587 VTAIL.n12 B 0.012707f
C588 VTAIL.n13 B 0.030036f
C589 VTAIL.n14 B 0.013455f
C590 VTAIL.n15 B 0.023648f
C591 VTAIL.n16 B 0.012707f
C592 VTAIL.n17 B 0.030036f
C593 VTAIL.n18 B 0.013455f
C594 VTAIL.n19 B 0.023648f
C595 VTAIL.n20 B 0.012707f
C596 VTAIL.n21 B 0.030036f
C597 VTAIL.n22 B 0.013455f
C598 VTAIL.n23 B 0.023648f
C599 VTAIL.n24 B 0.012707f
C600 VTAIL.n25 B 0.030036f
C601 VTAIL.n26 B 0.013455f
C602 VTAIL.n27 B 0.023648f
C603 VTAIL.n28 B 0.012707f
C604 VTAIL.n29 B 0.030036f
C605 VTAIL.n30 B 0.013455f
C606 VTAIL.n31 B 0.023648f
C607 VTAIL.n32 B 0.012707f
C608 VTAIL.n33 B 0.030036f
C609 VTAIL.n34 B 0.013455f
C610 VTAIL.n35 B 0.238593f
C611 VTAIL.t18 B 0.051684f
C612 VTAIL.n36 B 0.022527f
C613 VTAIL.n37 B 0.021233f
C614 VTAIL.n38 B 0.012707f
C615 VTAIL.n39 B 1.98189f
C616 VTAIL.n40 B 0.023648f
C617 VTAIL.n41 B 0.012707f
C618 VTAIL.n42 B 0.013455f
C619 VTAIL.n43 B 0.030036f
C620 VTAIL.n44 B 0.030036f
C621 VTAIL.n45 B 0.013455f
C622 VTAIL.n46 B 0.012707f
C623 VTAIL.n47 B 0.023648f
C624 VTAIL.n48 B 0.023648f
C625 VTAIL.n49 B 0.012707f
C626 VTAIL.n50 B 0.013455f
C627 VTAIL.n51 B 0.030036f
C628 VTAIL.n52 B 0.030036f
C629 VTAIL.n53 B 0.030036f
C630 VTAIL.n54 B 0.013455f
C631 VTAIL.n55 B 0.012707f
C632 VTAIL.n56 B 0.023648f
C633 VTAIL.n57 B 0.023648f
C634 VTAIL.n58 B 0.012707f
C635 VTAIL.n59 B 0.013081f
C636 VTAIL.n60 B 0.013081f
C637 VTAIL.n61 B 0.030036f
C638 VTAIL.n62 B 0.030036f
C639 VTAIL.n63 B 0.013455f
C640 VTAIL.n64 B 0.012707f
C641 VTAIL.n65 B 0.023648f
C642 VTAIL.n66 B 0.023648f
C643 VTAIL.n67 B 0.012707f
C644 VTAIL.n68 B 0.013455f
C645 VTAIL.n69 B 0.030036f
C646 VTAIL.n70 B 0.030036f
C647 VTAIL.n71 B 0.013455f
C648 VTAIL.n72 B 0.012707f
C649 VTAIL.n73 B 0.023648f
C650 VTAIL.n74 B 0.023648f
C651 VTAIL.n75 B 0.012707f
C652 VTAIL.n76 B 0.013455f
C653 VTAIL.n77 B 0.030036f
C654 VTAIL.n78 B 0.030036f
C655 VTAIL.n79 B 0.013455f
C656 VTAIL.n80 B 0.012707f
C657 VTAIL.n81 B 0.023648f
C658 VTAIL.n82 B 0.023648f
C659 VTAIL.n83 B 0.012707f
C660 VTAIL.n84 B 0.013455f
C661 VTAIL.n85 B 0.030036f
C662 VTAIL.n86 B 0.030036f
C663 VTAIL.n87 B 0.013455f
C664 VTAIL.n88 B 0.012707f
C665 VTAIL.n89 B 0.023648f
C666 VTAIL.n90 B 0.023648f
C667 VTAIL.n91 B 0.012707f
C668 VTAIL.n92 B 0.013455f
C669 VTAIL.n93 B 0.030036f
C670 VTAIL.n94 B 0.030036f
C671 VTAIL.n95 B 0.013455f
C672 VTAIL.n96 B 0.012707f
C673 VTAIL.n97 B 0.023648f
C674 VTAIL.n98 B 0.023648f
C675 VTAIL.n99 B 0.012707f
C676 VTAIL.n100 B 0.013455f
C677 VTAIL.n101 B 0.030036f
C678 VTAIL.n102 B 0.061894f
C679 VTAIL.n103 B 0.013455f
C680 VTAIL.n104 B 0.024847f
C681 VTAIL.n105 B 0.060477f
C682 VTAIL.n106 B 0.064479f
C683 VTAIL.n107 B 0.390363f
C684 VTAIL.t16 B 0.364407f
C685 VTAIL.t13 B 0.364407f
C686 VTAIL.n108 B 3.2728f
C687 VTAIL.n109 B 0.664052f
C688 VTAIL.t15 B 0.364407f
C689 VTAIL.t19 B 0.364407f
C690 VTAIL.n110 B 3.2728f
C691 VTAIL.n111 B 2.48695f
C692 VTAIL.t2 B 0.364407f
C693 VTAIL.t8 B 0.364407f
C694 VTAIL.n112 B 3.27281f
C695 VTAIL.n113 B 2.48693f
C696 VTAIL.t6 B 0.364407f
C697 VTAIL.t0 B 0.364407f
C698 VTAIL.n114 B 3.27281f
C699 VTAIL.n115 B 0.664038f
C700 VTAIL.n116 B 0.032761f
C701 VTAIL.n117 B 0.023648f
C702 VTAIL.n118 B 0.012707f
C703 VTAIL.n119 B 0.030036f
C704 VTAIL.n120 B 0.013455f
C705 VTAIL.n121 B 0.023648f
C706 VTAIL.n122 B 0.012707f
C707 VTAIL.n123 B 0.030036f
C708 VTAIL.n124 B 0.013455f
C709 VTAIL.n125 B 0.023648f
C710 VTAIL.n126 B 0.012707f
C711 VTAIL.n127 B 0.030036f
C712 VTAIL.n128 B 0.013455f
C713 VTAIL.n129 B 0.023648f
C714 VTAIL.n130 B 0.012707f
C715 VTAIL.n131 B 0.030036f
C716 VTAIL.n132 B 0.013455f
C717 VTAIL.n133 B 0.023648f
C718 VTAIL.n134 B 0.012707f
C719 VTAIL.n135 B 0.030036f
C720 VTAIL.n136 B 0.013455f
C721 VTAIL.n137 B 0.023648f
C722 VTAIL.n138 B 0.012707f
C723 VTAIL.n139 B 0.030036f
C724 VTAIL.n140 B 0.013455f
C725 VTAIL.n141 B 0.023648f
C726 VTAIL.n142 B 0.012707f
C727 VTAIL.n143 B 0.030036f
C728 VTAIL.n144 B 0.030036f
C729 VTAIL.n145 B 0.013455f
C730 VTAIL.n146 B 0.023648f
C731 VTAIL.n147 B 0.012707f
C732 VTAIL.n148 B 0.030036f
C733 VTAIL.n149 B 0.013455f
C734 VTAIL.n150 B 0.238593f
C735 VTAIL.t5 B 0.051684f
C736 VTAIL.n151 B 0.022527f
C737 VTAIL.n152 B 0.021233f
C738 VTAIL.n153 B 0.012707f
C739 VTAIL.n154 B 1.98189f
C740 VTAIL.n155 B 0.023648f
C741 VTAIL.n156 B 0.012707f
C742 VTAIL.n157 B 0.013455f
C743 VTAIL.n158 B 0.030036f
C744 VTAIL.n159 B 0.030036f
C745 VTAIL.n160 B 0.013455f
C746 VTAIL.n161 B 0.012707f
C747 VTAIL.n162 B 0.023648f
C748 VTAIL.n163 B 0.023648f
C749 VTAIL.n164 B 0.012707f
C750 VTAIL.n165 B 0.013455f
C751 VTAIL.n166 B 0.030036f
C752 VTAIL.n167 B 0.030036f
C753 VTAIL.n168 B 0.013455f
C754 VTAIL.n169 B 0.012707f
C755 VTAIL.n170 B 0.023648f
C756 VTAIL.n171 B 0.023648f
C757 VTAIL.n172 B 0.012707f
C758 VTAIL.n173 B 0.013081f
C759 VTAIL.n174 B 0.013081f
C760 VTAIL.n175 B 0.030036f
C761 VTAIL.n176 B 0.030036f
C762 VTAIL.n177 B 0.013455f
C763 VTAIL.n178 B 0.012707f
C764 VTAIL.n179 B 0.023648f
C765 VTAIL.n180 B 0.023648f
C766 VTAIL.n181 B 0.012707f
C767 VTAIL.n182 B 0.013455f
C768 VTAIL.n183 B 0.030036f
C769 VTAIL.n184 B 0.030036f
C770 VTAIL.n185 B 0.013455f
C771 VTAIL.n186 B 0.012707f
C772 VTAIL.n187 B 0.023648f
C773 VTAIL.n188 B 0.023648f
C774 VTAIL.n189 B 0.012707f
C775 VTAIL.n190 B 0.013455f
C776 VTAIL.n191 B 0.030036f
C777 VTAIL.n192 B 0.030036f
C778 VTAIL.n193 B 0.013455f
C779 VTAIL.n194 B 0.012707f
C780 VTAIL.n195 B 0.023648f
C781 VTAIL.n196 B 0.023648f
C782 VTAIL.n197 B 0.012707f
C783 VTAIL.n198 B 0.013455f
C784 VTAIL.n199 B 0.030036f
C785 VTAIL.n200 B 0.030036f
C786 VTAIL.n201 B 0.013455f
C787 VTAIL.n202 B 0.012707f
C788 VTAIL.n203 B 0.023648f
C789 VTAIL.n204 B 0.023648f
C790 VTAIL.n205 B 0.012707f
C791 VTAIL.n206 B 0.013455f
C792 VTAIL.n207 B 0.030036f
C793 VTAIL.n208 B 0.030036f
C794 VTAIL.n209 B 0.013455f
C795 VTAIL.n210 B 0.012707f
C796 VTAIL.n211 B 0.023648f
C797 VTAIL.n212 B 0.023648f
C798 VTAIL.n213 B 0.012707f
C799 VTAIL.n214 B 0.013455f
C800 VTAIL.n215 B 0.030036f
C801 VTAIL.n216 B 0.061894f
C802 VTAIL.n217 B 0.013455f
C803 VTAIL.n218 B 0.024847f
C804 VTAIL.n219 B 0.060477f
C805 VTAIL.n220 B 0.064479f
C806 VTAIL.n221 B 0.390363f
C807 VTAIL.t12 B 0.364407f
C808 VTAIL.t10 B 0.364407f
C809 VTAIL.n222 B 3.27281f
C810 VTAIL.n223 B 0.589481f
C811 VTAIL.t11 B 0.364407f
C812 VTAIL.t17 B 0.364407f
C813 VTAIL.n224 B 3.27281f
C814 VTAIL.n225 B 0.664038f
C815 VTAIL.n226 B 0.032761f
C816 VTAIL.n227 B 0.023648f
C817 VTAIL.n228 B 0.012707f
C818 VTAIL.n229 B 0.030036f
C819 VTAIL.n230 B 0.013455f
C820 VTAIL.n231 B 0.023648f
C821 VTAIL.n232 B 0.012707f
C822 VTAIL.n233 B 0.030036f
C823 VTAIL.n234 B 0.013455f
C824 VTAIL.n235 B 0.023648f
C825 VTAIL.n236 B 0.012707f
C826 VTAIL.n237 B 0.030036f
C827 VTAIL.n238 B 0.013455f
C828 VTAIL.n239 B 0.023648f
C829 VTAIL.n240 B 0.012707f
C830 VTAIL.n241 B 0.030036f
C831 VTAIL.n242 B 0.013455f
C832 VTAIL.n243 B 0.023648f
C833 VTAIL.n244 B 0.012707f
C834 VTAIL.n245 B 0.030036f
C835 VTAIL.n246 B 0.013455f
C836 VTAIL.n247 B 0.023648f
C837 VTAIL.n248 B 0.012707f
C838 VTAIL.n249 B 0.030036f
C839 VTAIL.n250 B 0.013455f
C840 VTAIL.n251 B 0.023648f
C841 VTAIL.n252 B 0.012707f
C842 VTAIL.n253 B 0.030036f
C843 VTAIL.n254 B 0.030036f
C844 VTAIL.n255 B 0.013455f
C845 VTAIL.n256 B 0.023648f
C846 VTAIL.n257 B 0.012707f
C847 VTAIL.n258 B 0.030036f
C848 VTAIL.n259 B 0.013455f
C849 VTAIL.n260 B 0.238593f
C850 VTAIL.t14 B 0.051684f
C851 VTAIL.n261 B 0.022527f
C852 VTAIL.n262 B 0.021233f
C853 VTAIL.n263 B 0.012707f
C854 VTAIL.n264 B 1.98189f
C855 VTAIL.n265 B 0.023648f
C856 VTAIL.n266 B 0.012707f
C857 VTAIL.n267 B 0.013455f
C858 VTAIL.n268 B 0.030036f
C859 VTAIL.n269 B 0.030036f
C860 VTAIL.n270 B 0.013455f
C861 VTAIL.n271 B 0.012707f
C862 VTAIL.n272 B 0.023648f
C863 VTAIL.n273 B 0.023648f
C864 VTAIL.n274 B 0.012707f
C865 VTAIL.n275 B 0.013455f
C866 VTAIL.n276 B 0.030036f
C867 VTAIL.n277 B 0.030036f
C868 VTAIL.n278 B 0.013455f
C869 VTAIL.n279 B 0.012707f
C870 VTAIL.n280 B 0.023648f
C871 VTAIL.n281 B 0.023648f
C872 VTAIL.n282 B 0.012707f
C873 VTAIL.n283 B 0.013081f
C874 VTAIL.n284 B 0.013081f
C875 VTAIL.n285 B 0.030036f
C876 VTAIL.n286 B 0.030036f
C877 VTAIL.n287 B 0.013455f
C878 VTAIL.n288 B 0.012707f
C879 VTAIL.n289 B 0.023648f
C880 VTAIL.n290 B 0.023648f
C881 VTAIL.n291 B 0.012707f
C882 VTAIL.n292 B 0.013455f
C883 VTAIL.n293 B 0.030036f
C884 VTAIL.n294 B 0.030036f
C885 VTAIL.n295 B 0.013455f
C886 VTAIL.n296 B 0.012707f
C887 VTAIL.n297 B 0.023648f
C888 VTAIL.n298 B 0.023648f
C889 VTAIL.n299 B 0.012707f
C890 VTAIL.n300 B 0.013455f
C891 VTAIL.n301 B 0.030036f
C892 VTAIL.n302 B 0.030036f
C893 VTAIL.n303 B 0.013455f
C894 VTAIL.n304 B 0.012707f
C895 VTAIL.n305 B 0.023648f
C896 VTAIL.n306 B 0.023648f
C897 VTAIL.n307 B 0.012707f
C898 VTAIL.n308 B 0.013455f
C899 VTAIL.n309 B 0.030036f
C900 VTAIL.n310 B 0.030036f
C901 VTAIL.n311 B 0.013455f
C902 VTAIL.n312 B 0.012707f
C903 VTAIL.n313 B 0.023648f
C904 VTAIL.n314 B 0.023648f
C905 VTAIL.n315 B 0.012707f
C906 VTAIL.n316 B 0.013455f
C907 VTAIL.n317 B 0.030036f
C908 VTAIL.n318 B 0.030036f
C909 VTAIL.n319 B 0.013455f
C910 VTAIL.n320 B 0.012707f
C911 VTAIL.n321 B 0.023648f
C912 VTAIL.n322 B 0.023648f
C913 VTAIL.n323 B 0.012707f
C914 VTAIL.n324 B 0.013455f
C915 VTAIL.n325 B 0.030036f
C916 VTAIL.n326 B 0.061894f
C917 VTAIL.n327 B 0.013455f
C918 VTAIL.n328 B 0.024847f
C919 VTAIL.n329 B 0.060477f
C920 VTAIL.n330 B 0.064479f
C921 VTAIL.n331 B 2.0671f
C922 VTAIL.n332 B 0.032761f
C923 VTAIL.n333 B 0.023648f
C924 VTAIL.n334 B 0.012707f
C925 VTAIL.n335 B 0.030036f
C926 VTAIL.n336 B 0.013455f
C927 VTAIL.n337 B 0.023648f
C928 VTAIL.n338 B 0.012707f
C929 VTAIL.n339 B 0.030036f
C930 VTAIL.n340 B 0.013455f
C931 VTAIL.n341 B 0.023648f
C932 VTAIL.n342 B 0.012707f
C933 VTAIL.n343 B 0.030036f
C934 VTAIL.n344 B 0.013455f
C935 VTAIL.n345 B 0.023648f
C936 VTAIL.n346 B 0.012707f
C937 VTAIL.n347 B 0.030036f
C938 VTAIL.n348 B 0.013455f
C939 VTAIL.n349 B 0.023648f
C940 VTAIL.n350 B 0.012707f
C941 VTAIL.n351 B 0.030036f
C942 VTAIL.n352 B 0.013455f
C943 VTAIL.n353 B 0.023648f
C944 VTAIL.n354 B 0.012707f
C945 VTAIL.n355 B 0.030036f
C946 VTAIL.n356 B 0.013455f
C947 VTAIL.n357 B 0.023648f
C948 VTAIL.n358 B 0.012707f
C949 VTAIL.n359 B 0.030036f
C950 VTAIL.n360 B 0.013455f
C951 VTAIL.n361 B 0.023648f
C952 VTAIL.n362 B 0.012707f
C953 VTAIL.n363 B 0.030036f
C954 VTAIL.n364 B 0.013455f
C955 VTAIL.n365 B 0.238593f
C956 VTAIL.t1 B 0.051684f
C957 VTAIL.n366 B 0.022527f
C958 VTAIL.n367 B 0.021233f
C959 VTAIL.n368 B 0.012707f
C960 VTAIL.n369 B 1.98189f
C961 VTAIL.n370 B 0.023648f
C962 VTAIL.n371 B 0.012707f
C963 VTAIL.n372 B 0.013455f
C964 VTAIL.n373 B 0.030036f
C965 VTAIL.n374 B 0.030036f
C966 VTAIL.n375 B 0.013455f
C967 VTAIL.n376 B 0.012707f
C968 VTAIL.n377 B 0.023648f
C969 VTAIL.n378 B 0.023648f
C970 VTAIL.n379 B 0.012707f
C971 VTAIL.n380 B 0.013455f
C972 VTAIL.n381 B 0.030036f
C973 VTAIL.n382 B 0.030036f
C974 VTAIL.n383 B 0.030036f
C975 VTAIL.n384 B 0.013455f
C976 VTAIL.n385 B 0.012707f
C977 VTAIL.n386 B 0.023648f
C978 VTAIL.n387 B 0.023648f
C979 VTAIL.n388 B 0.012707f
C980 VTAIL.n389 B 0.013081f
C981 VTAIL.n390 B 0.013081f
C982 VTAIL.n391 B 0.030036f
C983 VTAIL.n392 B 0.030036f
C984 VTAIL.n393 B 0.013455f
C985 VTAIL.n394 B 0.012707f
C986 VTAIL.n395 B 0.023648f
C987 VTAIL.n396 B 0.023648f
C988 VTAIL.n397 B 0.012707f
C989 VTAIL.n398 B 0.013455f
C990 VTAIL.n399 B 0.030036f
C991 VTAIL.n400 B 0.030036f
C992 VTAIL.n401 B 0.013455f
C993 VTAIL.n402 B 0.012707f
C994 VTAIL.n403 B 0.023648f
C995 VTAIL.n404 B 0.023648f
C996 VTAIL.n405 B 0.012707f
C997 VTAIL.n406 B 0.013455f
C998 VTAIL.n407 B 0.030036f
C999 VTAIL.n408 B 0.030036f
C1000 VTAIL.n409 B 0.013455f
C1001 VTAIL.n410 B 0.012707f
C1002 VTAIL.n411 B 0.023648f
C1003 VTAIL.n412 B 0.023648f
C1004 VTAIL.n413 B 0.012707f
C1005 VTAIL.n414 B 0.013455f
C1006 VTAIL.n415 B 0.030036f
C1007 VTAIL.n416 B 0.030036f
C1008 VTAIL.n417 B 0.013455f
C1009 VTAIL.n418 B 0.012707f
C1010 VTAIL.n419 B 0.023648f
C1011 VTAIL.n420 B 0.023648f
C1012 VTAIL.n421 B 0.012707f
C1013 VTAIL.n422 B 0.013455f
C1014 VTAIL.n423 B 0.030036f
C1015 VTAIL.n424 B 0.030036f
C1016 VTAIL.n425 B 0.013455f
C1017 VTAIL.n426 B 0.012707f
C1018 VTAIL.n427 B 0.023648f
C1019 VTAIL.n428 B 0.023648f
C1020 VTAIL.n429 B 0.012707f
C1021 VTAIL.n430 B 0.013455f
C1022 VTAIL.n431 B 0.030036f
C1023 VTAIL.n432 B 0.061894f
C1024 VTAIL.n433 B 0.013455f
C1025 VTAIL.n434 B 0.024847f
C1026 VTAIL.n435 B 0.060477f
C1027 VTAIL.n436 B 0.064479f
C1028 VTAIL.n437 B 2.0671f
C1029 VTAIL.t9 B 0.364407f
C1030 VTAIL.t3 B 0.364407f
C1031 VTAIL.n438 B 3.2728f
C1032 VTAIL.n439 B 0.494081f
C1033 VP.t4 B 3.01752f
C1034 VP.n0 B 1.11774f
C1035 VP.n1 B 0.01854f
C1036 VP.n2 B 0.029003f
C1037 VP.n3 B 0.01854f
C1038 VP.t9 B 3.01752f
C1039 VP.n4 B 0.034382f
C1040 VP.n5 B 0.01854f
C1041 VP.n6 B 0.034382f
C1042 VP.n7 B 0.01854f
C1043 VP.t8 B 3.01752f
C1044 VP.n8 B 0.034871f
C1045 VP.n9 B 0.01854f
C1046 VP.n10 B 0.021142f
C1047 VP.n11 B 0.01854f
C1048 VP.n12 B 0.024899f
C1049 VP.n13 B 0.029919f
C1050 VP.t5 B 3.01752f
C1051 VP.t0 B 3.01752f
C1052 VP.n14 B 1.11774f
C1053 VP.n15 B 0.01854f
C1054 VP.n16 B 0.029003f
C1055 VP.n17 B 0.01854f
C1056 VP.t3 B 3.01752f
C1057 VP.n18 B 0.034382f
C1058 VP.n19 B 0.01854f
C1059 VP.n20 B 0.034382f
C1060 VP.n21 B 0.01854f
C1061 VP.t2 B 3.01752f
C1062 VP.n22 B 0.034871f
C1063 VP.n23 B 0.01854f
C1064 VP.n24 B 0.021142f
C1065 VP.t7 B 3.21629f
C1066 VP.t6 B 3.01752f
C1067 VP.n25 B 1.09477f
C1068 VP.n26 B 1.06767f
C1069 VP.n27 B 0.199987f
C1070 VP.n28 B 0.01854f
C1071 VP.n29 B 0.034382f
C1072 VP.n30 B 0.037247f
C1073 VP.n31 B 0.016166f
C1074 VP.n32 B 0.01854f
C1075 VP.n33 B 0.01854f
C1076 VP.n34 B 0.01854f
C1077 VP.n35 B 0.034382f
C1078 VP.n36 B 0.025895f
C1079 VP.n37 B 1.0403f
C1080 VP.n38 B 0.025895f
C1081 VP.n39 B 0.01854f
C1082 VP.n40 B 0.01854f
C1083 VP.n41 B 0.01854f
C1084 VP.n42 B 0.034871f
C1085 VP.n43 B 0.016166f
C1086 VP.n44 B 0.037247f
C1087 VP.n45 B 0.01854f
C1088 VP.n46 B 0.01854f
C1089 VP.n47 B 0.01854f
C1090 VP.n48 B 0.021142f
C1091 VP.n49 B 1.0403f
C1092 VP.n50 B 0.030647f
C1093 VP.n51 B 0.034382f
C1094 VP.n52 B 0.01854f
C1095 VP.n53 B 0.01854f
C1096 VP.n54 B 0.01854f
C1097 VP.n55 B 0.024899f
C1098 VP.n56 B 0.034382f
C1099 VP.n57 B 0.033363f
C1100 VP.n58 B 0.029919f
C1101 VP.n59 B 1.38892f
C1102 VP.n60 B 1.39982f
C1103 VP.n61 B 1.11774f
C1104 VP.n62 B 0.033363f
C1105 VP.n63 B 0.034382f
C1106 VP.n64 B 0.01854f
C1107 VP.n65 B 0.01854f
C1108 VP.n66 B 0.01854f
C1109 VP.n67 B 0.029003f
C1110 VP.n68 B 0.034382f
C1111 VP.t1 B 3.01752f
C1112 VP.n69 B 1.0403f
C1113 VP.n70 B 0.030647f
C1114 VP.n71 B 0.01854f
C1115 VP.n72 B 0.01854f
C1116 VP.n73 B 0.01854f
C1117 VP.n74 B 0.034382f
C1118 VP.n75 B 0.037247f
C1119 VP.n76 B 0.016166f
C1120 VP.n77 B 0.01854f
C1121 VP.n78 B 0.01854f
C1122 VP.n79 B 0.01854f
C1123 VP.n80 B 0.034382f
C1124 VP.n81 B 0.025895f
C1125 VP.n82 B 1.0403f
C1126 VP.n83 B 0.025895f
C1127 VP.n84 B 0.01854f
C1128 VP.n85 B 0.01854f
C1129 VP.n86 B 0.01854f
C1130 VP.n87 B 0.034871f
C1131 VP.n88 B 0.016166f
C1132 VP.n89 B 0.037247f
C1133 VP.n90 B 0.01854f
C1134 VP.n91 B 0.01854f
C1135 VP.n92 B 0.01854f
C1136 VP.n93 B 0.021142f
C1137 VP.n94 B 1.0403f
C1138 VP.n95 B 0.030647f
C1139 VP.n96 B 0.034382f
C1140 VP.n97 B 0.01854f
C1141 VP.n98 B 0.01854f
C1142 VP.n99 B 0.01854f
C1143 VP.n100 B 0.024899f
C1144 VP.n101 B 0.034382f
C1145 VP.n102 B 0.033363f
C1146 VP.n103 B 0.029919f
C1147 VP.n104 B 0.036024f
.ends

