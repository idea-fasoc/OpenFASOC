* NGSPICE file created from diff_pair_sample_1013.ext - technology: sky130A

.subckt diff_pair_sample_1013 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=6.318 ps=33.18 w=16.2 l=1.72
X1 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X2 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X3 VTAIL.t10 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=2.673 ps=16.53 w=16.2 l=1.72
X4 VDD2.t5 VN.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=6.318 ps=33.18 w=16.2 l=1.72
X5 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=2.673 ps=16.53 w=16.2 l=1.72
X6 VTAIL.t12 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X7 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=0 ps=0 w=16.2 l=1.72
X8 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=0 ps=0 w=16.2 l=1.72
X9 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=0 ps=0 w=16.2 l=1.72
X10 VTAIL.t14 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X11 VDD2.t3 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=6.318 ps=33.18 w=16.2 l=1.72
X12 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X13 VDD1.t3 VP.t4 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X14 VTAIL.t3 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=2.673 ps=16.53 w=16.2 l=1.72
X15 VDD1.t2 VP.t5 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X16 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=2.673 ps=16.53 w=16.2 l=1.72
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=0 ps=0 w=16.2 l=1.72
X18 VDD1.t1 VP.t6 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.673 pd=16.53 as=6.318 ps=33.18 w=16.2 l=1.72
X19 VTAIL.t13 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=6.318 pd=33.18 as=2.673 ps=16.53 w=16.2 l=1.72
R0 VP.n12 VP.t1 256.594
R1 VP.n31 VP.t7 226.988
R2 VP.n38 VP.t4 226.988
R3 VP.n46 VP.t2 226.988
R4 VP.n53 VP.t6 226.988
R5 VP.n28 VP.t0 226.988
R6 VP.n21 VP.t3 226.988
R7 VP.n13 VP.t5 226.988
R8 VP.n31 VP.n30 182.203
R9 VP.n54 VP.n53 182.203
R10 VP.n29 VP.n28 182.203
R11 VP.n14 VP.n11 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n10 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n20 VP.n9 161.3
R16 VP.n23 VP.n22 161.3
R17 VP.n24 VP.n8 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n27 VP.n7 161.3
R20 VP.n52 VP.n0 161.3
R21 VP.n51 VP.n50 161.3
R22 VP.n49 VP.n1 161.3
R23 VP.n48 VP.n47 161.3
R24 VP.n45 VP.n2 161.3
R25 VP.n44 VP.n43 161.3
R26 VP.n42 VP.n3 161.3
R27 VP.n41 VP.n40 161.3
R28 VP.n39 VP.n4 161.3
R29 VP.n37 VP.n36 161.3
R30 VP.n35 VP.n5 161.3
R31 VP.n34 VP.n33 161.3
R32 VP.n32 VP.n6 161.3
R33 VP.n13 VP.n12 67.3815
R34 VP.n30 VP.n29 49.8414
R35 VP.n33 VP.n5 45.4209
R36 VP.n51 VP.n1 45.4209
R37 VP.n26 VP.n8 45.4209
R38 VP.n40 VP.n3 40.577
R39 VP.n44 VP.n3 40.577
R40 VP.n19 VP.n10 40.577
R41 VP.n15 VP.n10 40.577
R42 VP.n37 VP.n5 35.7332
R43 VP.n47 VP.n1 35.7332
R44 VP.n22 VP.n8 35.7332
R45 VP.n33 VP.n32 24.5923
R46 VP.n40 VP.n39 24.5923
R47 VP.n45 VP.n44 24.5923
R48 VP.n52 VP.n51 24.5923
R49 VP.n27 VP.n26 24.5923
R50 VP.n20 VP.n19 24.5923
R51 VP.n15 VP.n14 24.5923
R52 VP.n38 VP.n37 23.3627
R53 VP.n47 VP.n46 23.3627
R54 VP.n22 VP.n21 23.3627
R55 VP.n12 VP.n11 18.5926
R56 VP.n32 VP.n31 3.68928
R57 VP.n53 VP.n52 3.68928
R58 VP.n28 VP.n27 3.68928
R59 VP.n39 VP.n38 1.23009
R60 VP.n46 VP.n45 1.23009
R61 VP.n21 VP.n20 1.23009
R62 VP.n14 VP.n13 1.23009
R63 VP.n16 VP.n11 0.189894
R64 VP.n17 VP.n16 0.189894
R65 VP.n18 VP.n17 0.189894
R66 VP.n18 VP.n9 0.189894
R67 VP.n23 VP.n9 0.189894
R68 VP.n24 VP.n23 0.189894
R69 VP.n25 VP.n24 0.189894
R70 VP.n25 VP.n7 0.189894
R71 VP.n29 VP.n7 0.189894
R72 VP.n30 VP.n6 0.189894
R73 VP.n34 VP.n6 0.189894
R74 VP.n35 VP.n34 0.189894
R75 VP.n36 VP.n35 0.189894
R76 VP.n36 VP.n4 0.189894
R77 VP.n41 VP.n4 0.189894
R78 VP.n42 VP.n41 0.189894
R79 VP.n43 VP.n42 0.189894
R80 VP.n43 VP.n2 0.189894
R81 VP.n48 VP.n2 0.189894
R82 VP.n49 VP.n48 0.189894
R83 VP.n50 VP.n49 0.189894
R84 VP.n50 VP.n0 0.189894
R85 VP.n54 VP.n0 0.189894
R86 VP VP.n54 0.0516364
R87 VTAIL.n722 VTAIL.n638 289.615
R88 VTAIL.n86 VTAIL.n2 289.615
R89 VTAIL.n176 VTAIL.n92 289.615
R90 VTAIL.n268 VTAIL.n184 289.615
R91 VTAIL.n632 VTAIL.n548 289.615
R92 VTAIL.n540 VTAIL.n456 289.615
R93 VTAIL.n450 VTAIL.n366 289.615
R94 VTAIL.n358 VTAIL.n274 289.615
R95 VTAIL.n666 VTAIL.n665 185
R96 VTAIL.n671 VTAIL.n670 185
R97 VTAIL.n673 VTAIL.n672 185
R98 VTAIL.n662 VTAIL.n661 185
R99 VTAIL.n679 VTAIL.n678 185
R100 VTAIL.n681 VTAIL.n680 185
R101 VTAIL.n658 VTAIL.n657 185
R102 VTAIL.n687 VTAIL.n686 185
R103 VTAIL.n689 VTAIL.n688 185
R104 VTAIL.n654 VTAIL.n653 185
R105 VTAIL.n695 VTAIL.n694 185
R106 VTAIL.n697 VTAIL.n696 185
R107 VTAIL.n650 VTAIL.n649 185
R108 VTAIL.n703 VTAIL.n702 185
R109 VTAIL.n705 VTAIL.n704 185
R110 VTAIL.n646 VTAIL.n645 185
R111 VTAIL.n712 VTAIL.n711 185
R112 VTAIL.n713 VTAIL.n644 185
R113 VTAIL.n715 VTAIL.n714 185
R114 VTAIL.n642 VTAIL.n641 185
R115 VTAIL.n721 VTAIL.n720 185
R116 VTAIL.n723 VTAIL.n722 185
R117 VTAIL.n30 VTAIL.n29 185
R118 VTAIL.n35 VTAIL.n34 185
R119 VTAIL.n37 VTAIL.n36 185
R120 VTAIL.n26 VTAIL.n25 185
R121 VTAIL.n43 VTAIL.n42 185
R122 VTAIL.n45 VTAIL.n44 185
R123 VTAIL.n22 VTAIL.n21 185
R124 VTAIL.n51 VTAIL.n50 185
R125 VTAIL.n53 VTAIL.n52 185
R126 VTAIL.n18 VTAIL.n17 185
R127 VTAIL.n59 VTAIL.n58 185
R128 VTAIL.n61 VTAIL.n60 185
R129 VTAIL.n14 VTAIL.n13 185
R130 VTAIL.n67 VTAIL.n66 185
R131 VTAIL.n69 VTAIL.n68 185
R132 VTAIL.n10 VTAIL.n9 185
R133 VTAIL.n76 VTAIL.n75 185
R134 VTAIL.n77 VTAIL.n8 185
R135 VTAIL.n79 VTAIL.n78 185
R136 VTAIL.n6 VTAIL.n5 185
R137 VTAIL.n85 VTAIL.n84 185
R138 VTAIL.n87 VTAIL.n86 185
R139 VTAIL.n120 VTAIL.n119 185
R140 VTAIL.n125 VTAIL.n124 185
R141 VTAIL.n127 VTAIL.n126 185
R142 VTAIL.n116 VTAIL.n115 185
R143 VTAIL.n133 VTAIL.n132 185
R144 VTAIL.n135 VTAIL.n134 185
R145 VTAIL.n112 VTAIL.n111 185
R146 VTAIL.n141 VTAIL.n140 185
R147 VTAIL.n143 VTAIL.n142 185
R148 VTAIL.n108 VTAIL.n107 185
R149 VTAIL.n149 VTAIL.n148 185
R150 VTAIL.n151 VTAIL.n150 185
R151 VTAIL.n104 VTAIL.n103 185
R152 VTAIL.n157 VTAIL.n156 185
R153 VTAIL.n159 VTAIL.n158 185
R154 VTAIL.n100 VTAIL.n99 185
R155 VTAIL.n166 VTAIL.n165 185
R156 VTAIL.n167 VTAIL.n98 185
R157 VTAIL.n169 VTAIL.n168 185
R158 VTAIL.n96 VTAIL.n95 185
R159 VTAIL.n175 VTAIL.n174 185
R160 VTAIL.n177 VTAIL.n176 185
R161 VTAIL.n212 VTAIL.n211 185
R162 VTAIL.n217 VTAIL.n216 185
R163 VTAIL.n219 VTAIL.n218 185
R164 VTAIL.n208 VTAIL.n207 185
R165 VTAIL.n225 VTAIL.n224 185
R166 VTAIL.n227 VTAIL.n226 185
R167 VTAIL.n204 VTAIL.n203 185
R168 VTAIL.n233 VTAIL.n232 185
R169 VTAIL.n235 VTAIL.n234 185
R170 VTAIL.n200 VTAIL.n199 185
R171 VTAIL.n241 VTAIL.n240 185
R172 VTAIL.n243 VTAIL.n242 185
R173 VTAIL.n196 VTAIL.n195 185
R174 VTAIL.n249 VTAIL.n248 185
R175 VTAIL.n251 VTAIL.n250 185
R176 VTAIL.n192 VTAIL.n191 185
R177 VTAIL.n258 VTAIL.n257 185
R178 VTAIL.n259 VTAIL.n190 185
R179 VTAIL.n261 VTAIL.n260 185
R180 VTAIL.n188 VTAIL.n187 185
R181 VTAIL.n267 VTAIL.n266 185
R182 VTAIL.n269 VTAIL.n268 185
R183 VTAIL.n633 VTAIL.n632 185
R184 VTAIL.n631 VTAIL.n630 185
R185 VTAIL.n552 VTAIL.n551 185
R186 VTAIL.n625 VTAIL.n624 185
R187 VTAIL.n623 VTAIL.n554 185
R188 VTAIL.n622 VTAIL.n621 185
R189 VTAIL.n557 VTAIL.n555 185
R190 VTAIL.n616 VTAIL.n615 185
R191 VTAIL.n614 VTAIL.n613 185
R192 VTAIL.n561 VTAIL.n560 185
R193 VTAIL.n608 VTAIL.n607 185
R194 VTAIL.n606 VTAIL.n605 185
R195 VTAIL.n565 VTAIL.n564 185
R196 VTAIL.n600 VTAIL.n599 185
R197 VTAIL.n598 VTAIL.n597 185
R198 VTAIL.n569 VTAIL.n568 185
R199 VTAIL.n592 VTAIL.n591 185
R200 VTAIL.n590 VTAIL.n589 185
R201 VTAIL.n573 VTAIL.n572 185
R202 VTAIL.n584 VTAIL.n583 185
R203 VTAIL.n582 VTAIL.n581 185
R204 VTAIL.n577 VTAIL.n576 185
R205 VTAIL.n541 VTAIL.n540 185
R206 VTAIL.n539 VTAIL.n538 185
R207 VTAIL.n460 VTAIL.n459 185
R208 VTAIL.n533 VTAIL.n532 185
R209 VTAIL.n531 VTAIL.n462 185
R210 VTAIL.n530 VTAIL.n529 185
R211 VTAIL.n465 VTAIL.n463 185
R212 VTAIL.n524 VTAIL.n523 185
R213 VTAIL.n522 VTAIL.n521 185
R214 VTAIL.n469 VTAIL.n468 185
R215 VTAIL.n516 VTAIL.n515 185
R216 VTAIL.n514 VTAIL.n513 185
R217 VTAIL.n473 VTAIL.n472 185
R218 VTAIL.n508 VTAIL.n507 185
R219 VTAIL.n506 VTAIL.n505 185
R220 VTAIL.n477 VTAIL.n476 185
R221 VTAIL.n500 VTAIL.n499 185
R222 VTAIL.n498 VTAIL.n497 185
R223 VTAIL.n481 VTAIL.n480 185
R224 VTAIL.n492 VTAIL.n491 185
R225 VTAIL.n490 VTAIL.n489 185
R226 VTAIL.n485 VTAIL.n484 185
R227 VTAIL.n451 VTAIL.n450 185
R228 VTAIL.n449 VTAIL.n448 185
R229 VTAIL.n370 VTAIL.n369 185
R230 VTAIL.n443 VTAIL.n442 185
R231 VTAIL.n441 VTAIL.n372 185
R232 VTAIL.n440 VTAIL.n439 185
R233 VTAIL.n375 VTAIL.n373 185
R234 VTAIL.n434 VTAIL.n433 185
R235 VTAIL.n432 VTAIL.n431 185
R236 VTAIL.n379 VTAIL.n378 185
R237 VTAIL.n426 VTAIL.n425 185
R238 VTAIL.n424 VTAIL.n423 185
R239 VTAIL.n383 VTAIL.n382 185
R240 VTAIL.n418 VTAIL.n417 185
R241 VTAIL.n416 VTAIL.n415 185
R242 VTAIL.n387 VTAIL.n386 185
R243 VTAIL.n410 VTAIL.n409 185
R244 VTAIL.n408 VTAIL.n407 185
R245 VTAIL.n391 VTAIL.n390 185
R246 VTAIL.n402 VTAIL.n401 185
R247 VTAIL.n400 VTAIL.n399 185
R248 VTAIL.n395 VTAIL.n394 185
R249 VTAIL.n359 VTAIL.n358 185
R250 VTAIL.n357 VTAIL.n356 185
R251 VTAIL.n278 VTAIL.n277 185
R252 VTAIL.n351 VTAIL.n350 185
R253 VTAIL.n349 VTAIL.n280 185
R254 VTAIL.n348 VTAIL.n347 185
R255 VTAIL.n283 VTAIL.n281 185
R256 VTAIL.n342 VTAIL.n341 185
R257 VTAIL.n340 VTAIL.n339 185
R258 VTAIL.n287 VTAIL.n286 185
R259 VTAIL.n334 VTAIL.n333 185
R260 VTAIL.n332 VTAIL.n331 185
R261 VTAIL.n291 VTAIL.n290 185
R262 VTAIL.n326 VTAIL.n325 185
R263 VTAIL.n324 VTAIL.n323 185
R264 VTAIL.n295 VTAIL.n294 185
R265 VTAIL.n318 VTAIL.n317 185
R266 VTAIL.n316 VTAIL.n315 185
R267 VTAIL.n299 VTAIL.n298 185
R268 VTAIL.n310 VTAIL.n309 185
R269 VTAIL.n308 VTAIL.n307 185
R270 VTAIL.n303 VTAIL.n302 185
R271 VTAIL.n667 VTAIL.t5 147.659
R272 VTAIL.n31 VTAIL.t3 147.659
R273 VTAIL.n121 VTAIL.t8 147.659
R274 VTAIL.n213 VTAIL.t13 147.659
R275 VTAIL.n578 VTAIL.t15 147.659
R276 VTAIL.n486 VTAIL.t10 147.659
R277 VTAIL.n396 VTAIL.t7 147.659
R278 VTAIL.n304 VTAIL.t6 147.659
R279 VTAIL.n671 VTAIL.n665 104.615
R280 VTAIL.n672 VTAIL.n671 104.615
R281 VTAIL.n672 VTAIL.n661 104.615
R282 VTAIL.n679 VTAIL.n661 104.615
R283 VTAIL.n680 VTAIL.n679 104.615
R284 VTAIL.n680 VTAIL.n657 104.615
R285 VTAIL.n687 VTAIL.n657 104.615
R286 VTAIL.n688 VTAIL.n687 104.615
R287 VTAIL.n688 VTAIL.n653 104.615
R288 VTAIL.n695 VTAIL.n653 104.615
R289 VTAIL.n696 VTAIL.n695 104.615
R290 VTAIL.n696 VTAIL.n649 104.615
R291 VTAIL.n703 VTAIL.n649 104.615
R292 VTAIL.n704 VTAIL.n703 104.615
R293 VTAIL.n704 VTAIL.n645 104.615
R294 VTAIL.n712 VTAIL.n645 104.615
R295 VTAIL.n713 VTAIL.n712 104.615
R296 VTAIL.n714 VTAIL.n713 104.615
R297 VTAIL.n714 VTAIL.n641 104.615
R298 VTAIL.n721 VTAIL.n641 104.615
R299 VTAIL.n722 VTAIL.n721 104.615
R300 VTAIL.n35 VTAIL.n29 104.615
R301 VTAIL.n36 VTAIL.n35 104.615
R302 VTAIL.n36 VTAIL.n25 104.615
R303 VTAIL.n43 VTAIL.n25 104.615
R304 VTAIL.n44 VTAIL.n43 104.615
R305 VTAIL.n44 VTAIL.n21 104.615
R306 VTAIL.n51 VTAIL.n21 104.615
R307 VTAIL.n52 VTAIL.n51 104.615
R308 VTAIL.n52 VTAIL.n17 104.615
R309 VTAIL.n59 VTAIL.n17 104.615
R310 VTAIL.n60 VTAIL.n59 104.615
R311 VTAIL.n60 VTAIL.n13 104.615
R312 VTAIL.n67 VTAIL.n13 104.615
R313 VTAIL.n68 VTAIL.n67 104.615
R314 VTAIL.n68 VTAIL.n9 104.615
R315 VTAIL.n76 VTAIL.n9 104.615
R316 VTAIL.n77 VTAIL.n76 104.615
R317 VTAIL.n78 VTAIL.n77 104.615
R318 VTAIL.n78 VTAIL.n5 104.615
R319 VTAIL.n85 VTAIL.n5 104.615
R320 VTAIL.n86 VTAIL.n85 104.615
R321 VTAIL.n125 VTAIL.n119 104.615
R322 VTAIL.n126 VTAIL.n125 104.615
R323 VTAIL.n126 VTAIL.n115 104.615
R324 VTAIL.n133 VTAIL.n115 104.615
R325 VTAIL.n134 VTAIL.n133 104.615
R326 VTAIL.n134 VTAIL.n111 104.615
R327 VTAIL.n141 VTAIL.n111 104.615
R328 VTAIL.n142 VTAIL.n141 104.615
R329 VTAIL.n142 VTAIL.n107 104.615
R330 VTAIL.n149 VTAIL.n107 104.615
R331 VTAIL.n150 VTAIL.n149 104.615
R332 VTAIL.n150 VTAIL.n103 104.615
R333 VTAIL.n157 VTAIL.n103 104.615
R334 VTAIL.n158 VTAIL.n157 104.615
R335 VTAIL.n158 VTAIL.n99 104.615
R336 VTAIL.n166 VTAIL.n99 104.615
R337 VTAIL.n167 VTAIL.n166 104.615
R338 VTAIL.n168 VTAIL.n167 104.615
R339 VTAIL.n168 VTAIL.n95 104.615
R340 VTAIL.n175 VTAIL.n95 104.615
R341 VTAIL.n176 VTAIL.n175 104.615
R342 VTAIL.n217 VTAIL.n211 104.615
R343 VTAIL.n218 VTAIL.n217 104.615
R344 VTAIL.n218 VTAIL.n207 104.615
R345 VTAIL.n225 VTAIL.n207 104.615
R346 VTAIL.n226 VTAIL.n225 104.615
R347 VTAIL.n226 VTAIL.n203 104.615
R348 VTAIL.n233 VTAIL.n203 104.615
R349 VTAIL.n234 VTAIL.n233 104.615
R350 VTAIL.n234 VTAIL.n199 104.615
R351 VTAIL.n241 VTAIL.n199 104.615
R352 VTAIL.n242 VTAIL.n241 104.615
R353 VTAIL.n242 VTAIL.n195 104.615
R354 VTAIL.n249 VTAIL.n195 104.615
R355 VTAIL.n250 VTAIL.n249 104.615
R356 VTAIL.n250 VTAIL.n191 104.615
R357 VTAIL.n258 VTAIL.n191 104.615
R358 VTAIL.n259 VTAIL.n258 104.615
R359 VTAIL.n260 VTAIL.n259 104.615
R360 VTAIL.n260 VTAIL.n187 104.615
R361 VTAIL.n267 VTAIL.n187 104.615
R362 VTAIL.n268 VTAIL.n267 104.615
R363 VTAIL.n632 VTAIL.n631 104.615
R364 VTAIL.n631 VTAIL.n551 104.615
R365 VTAIL.n624 VTAIL.n551 104.615
R366 VTAIL.n624 VTAIL.n623 104.615
R367 VTAIL.n623 VTAIL.n622 104.615
R368 VTAIL.n622 VTAIL.n555 104.615
R369 VTAIL.n615 VTAIL.n555 104.615
R370 VTAIL.n615 VTAIL.n614 104.615
R371 VTAIL.n614 VTAIL.n560 104.615
R372 VTAIL.n607 VTAIL.n560 104.615
R373 VTAIL.n607 VTAIL.n606 104.615
R374 VTAIL.n606 VTAIL.n564 104.615
R375 VTAIL.n599 VTAIL.n564 104.615
R376 VTAIL.n599 VTAIL.n598 104.615
R377 VTAIL.n598 VTAIL.n568 104.615
R378 VTAIL.n591 VTAIL.n568 104.615
R379 VTAIL.n591 VTAIL.n590 104.615
R380 VTAIL.n590 VTAIL.n572 104.615
R381 VTAIL.n583 VTAIL.n572 104.615
R382 VTAIL.n583 VTAIL.n582 104.615
R383 VTAIL.n582 VTAIL.n576 104.615
R384 VTAIL.n540 VTAIL.n539 104.615
R385 VTAIL.n539 VTAIL.n459 104.615
R386 VTAIL.n532 VTAIL.n459 104.615
R387 VTAIL.n532 VTAIL.n531 104.615
R388 VTAIL.n531 VTAIL.n530 104.615
R389 VTAIL.n530 VTAIL.n463 104.615
R390 VTAIL.n523 VTAIL.n463 104.615
R391 VTAIL.n523 VTAIL.n522 104.615
R392 VTAIL.n522 VTAIL.n468 104.615
R393 VTAIL.n515 VTAIL.n468 104.615
R394 VTAIL.n515 VTAIL.n514 104.615
R395 VTAIL.n514 VTAIL.n472 104.615
R396 VTAIL.n507 VTAIL.n472 104.615
R397 VTAIL.n507 VTAIL.n506 104.615
R398 VTAIL.n506 VTAIL.n476 104.615
R399 VTAIL.n499 VTAIL.n476 104.615
R400 VTAIL.n499 VTAIL.n498 104.615
R401 VTAIL.n498 VTAIL.n480 104.615
R402 VTAIL.n491 VTAIL.n480 104.615
R403 VTAIL.n491 VTAIL.n490 104.615
R404 VTAIL.n490 VTAIL.n484 104.615
R405 VTAIL.n450 VTAIL.n449 104.615
R406 VTAIL.n449 VTAIL.n369 104.615
R407 VTAIL.n442 VTAIL.n369 104.615
R408 VTAIL.n442 VTAIL.n441 104.615
R409 VTAIL.n441 VTAIL.n440 104.615
R410 VTAIL.n440 VTAIL.n373 104.615
R411 VTAIL.n433 VTAIL.n373 104.615
R412 VTAIL.n433 VTAIL.n432 104.615
R413 VTAIL.n432 VTAIL.n378 104.615
R414 VTAIL.n425 VTAIL.n378 104.615
R415 VTAIL.n425 VTAIL.n424 104.615
R416 VTAIL.n424 VTAIL.n382 104.615
R417 VTAIL.n417 VTAIL.n382 104.615
R418 VTAIL.n417 VTAIL.n416 104.615
R419 VTAIL.n416 VTAIL.n386 104.615
R420 VTAIL.n409 VTAIL.n386 104.615
R421 VTAIL.n409 VTAIL.n408 104.615
R422 VTAIL.n408 VTAIL.n390 104.615
R423 VTAIL.n401 VTAIL.n390 104.615
R424 VTAIL.n401 VTAIL.n400 104.615
R425 VTAIL.n400 VTAIL.n394 104.615
R426 VTAIL.n358 VTAIL.n357 104.615
R427 VTAIL.n357 VTAIL.n277 104.615
R428 VTAIL.n350 VTAIL.n277 104.615
R429 VTAIL.n350 VTAIL.n349 104.615
R430 VTAIL.n349 VTAIL.n348 104.615
R431 VTAIL.n348 VTAIL.n281 104.615
R432 VTAIL.n341 VTAIL.n281 104.615
R433 VTAIL.n341 VTAIL.n340 104.615
R434 VTAIL.n340 VTAIL.n286 104.615
R435 VTAIL.n333 VTAIL.n286 104.615
R436 VTAIL.n333 VTAIL.n332 104.615
R437 VTAIL.n332 VTAIL.n290 104.615
R438 VTAIL.n325 VTAIL.n290 104.615
R439 VTAIL.n325 VTAIL.n324 104.615
R440 VTAIL.n324 VTAIL.n294 104.615
R441 VTAIL.n317 VTAIL.n294 104.615
R442 VTAIL.n317 VTAIL.n316 104.615
R443 VTAIL.n316 VTAIL.n298 104.615
R444 VTAIL.n309 VTAIL.n298 104.615
R445 VTAIL.n309 VTAIL.n308 104.615
R446 VTAIL.n308 VTAIL.n302 104.615
R447 VTAIL.t5 VTAIL.n665 52.3082
R448 VTAIL.t3 VTAIL.n29 52.3082
R449 VTAIL.t8 VTAIL.n119 52.3082
R450 VTAIL.t13 VTAIL.n211 52.3082
R451 VTAIL.t15 VTAIL.n576 52.3082
R452 VTAIL.t10 VTAIL.n484 52.3082
R453 VTAIL.t7 VTAIL.n394 52.3082
R454 VTAIL.t6 VTAIL.n302 52.3082
R455 VTAIL.n547 VTAIL.n546 46.4262
R456 VTAIL.n365 VTAIL.n364 46.4262
R457 VTAIL.n1 VTAIL.n0 46.426
R458 VTAIL.n183 VTAIL.n182 46.426
R459 VTAIL.n727 VTAIL.n726 34.5126
R460 VTAIL.n91 VTAIL.n90 34.5126
R461 VTAIL.n181 VTAIL.n180 34.5126
R462 VTAIL.n273 VTAIL.n272 34.5126
R463 VTAIL.n637 VTAIL.n636 34.5126
R464 VTAIL.n545 VTAIL.n544 34.5126
R465 VTAIL.n455 VTAIL.n454 34.5126
R466 VTAIL.n363 VTAIL.n362 34.5126
R467 VTAIL.n727 VTAIL.n637 28.0996
R468 VTAIL.n363 VTAIL.n273 28.0996
R469 VTAIL.n667 VTAIL.n666 15.6677
R470 VTAIL.n31 VTAIL.n30 15.6677
R471 VTAIL.n121 VTAIL.n120 15.6677
R472 VTAIL.n213 VTAIL.n212 15.6677
R473 VTAIL.n578 VTAIL.n577 15.6677
R474 VTAIL.n486 VTAIL.n485 15.6677
R475 VTAIL.n396 VTAIL.n395 15.6677
R476 VTAIL.n304 VTAIL.n303 15.6677
R477 VTAIL.n715 VTAIL.n644 13.1884
R478 VTAIL.n79 VTAIL.n8 13.1884
R479 VTAIL.n169 VTAIL.n98 13.1884
R480 VTAIL.n261 VTAIL.n190 13.1884
R481 VTAIL.n625 VTAIL.n554 13.1884
R482 VTAIL.n533 VTAIL.n462 13.1884
R483 VTAIL.n443 VTAIL.n372 13.1884
R484 VTAIL.n351 VTAIL.n280 13.1884
R485 VTAIL.n670 VTAIL.n669 12.8005
R486 VTAIL.n711 VTAIL.n710 12.8005
R487 VTAIL.n716 VTAIL.n642 12.8005
R488 VTAIL.n34 VTAIL.n33 12.8005
R489 VTAIL.n75 VTAIL.n74 12.8005
R490 VTAIL.n80 VTAIL.n6 12.8005
R491 VTAIL.n124 VTAIL.n123 12.8005
R492 VTAIL.n165 VTAIL.n164 12.8005
R493 VTAIL.n170 VTAIL.n96 12.8005
R494 VTAIL.n216 VTAIL.n215 12.8005
R495 VTAIL.n257 VTAIL.n256 12.8005
R496 VTAIL.n262 VTAIL.n188 12.8005
R497 VTAIL.n626 VTAIL.n552 12.8005
R498 VTAIL.n621 VTAIL.n556 12.8005
R499 VTAIL.n581 VTAIL.n580 12.8005
R500 VTAIL.n534 VTAIL.n460 12.8005
R501 VTAIL.n529 VTAIL.n464 12.8005
R502 VTAIL.n489 VTAIL.n488 12.8005
R503 VTAIL.n444 VTAIL.n370 12.8005
R504 VTAIL.n439 VTAIL.n374 12.8005
R505 VTAIL.n399 VTAIL.n398 12.8005
R506 VTAIL.n352 VTAIL.n278 12.8005
R507 VTAIL.n347 VTAIL.n282 12.8005
R508 VTAIL.n307 VTAIL.n306 12.8005
R509 VTAIL.n673 VTAIL.n664 12.0247
R510 VTAIL.n709 VTAIL.n646 12.0247
R511 VTAIL.n720 VTAIL.n719 12.0247
R512 VTAIL.n37 VTAIL.n28 12.0247
R513 VTAIL.n73 VTAIL.n10 12.0247
R514 VTAIL.n84 VTAIL.n83 12.0247
R515 VTAIL.n127 VTAIL.n118 12.0247
R516 VTAIL.n163 VTAIL.n100 12.0247
R517 VTAIL.n174 VTAIL.n173 12.0247
R518 VTAIL.n219 VTAIL.n210 12.0247
R519 VTAIL.n255 VTAIL.n192 12.0247
R520 VTAIL.n266 VTAIL.n265 12.0247
R521 VTAIL.n630 VTAIL.n629 12.0247
R522 VTAIL.n620 VTAIL.n557 12.0247
R523 VTAIL.n584 VTAIL.n575 12.0247
R524 VTAIL.n538 VTAIL.n537 12.0247
R525 VTAIL.n528 VTAIL.n465 12.0247
R526 VTAIL.n492 VTAIL.n483 12.0247
R527 VTAIL.n448 VTAIL.n447 12.0247
R528 VTAIL.n438 VTAIL.n375 12.0247
R529 VTAIL.n402 VTAIL.n393 12.0247
R530 VTAIL.n356 VTAIL.n355 12.0247
R531 VTAIL.n346 VTAIL.n283 12.0247
R532 VTAIL.n310 VTAIL.n301 12.0247
R533 VTAIL.n674 VTAIL.n662 11.249
R534 VTAIL.n706 VTAIL.n705 11.249
R535 VTAIL.n723 VTAIL.n640 11.249
R536 VTAIL.n38 VTAIL.n26 11.249
R537 VTAIL.n70 VTAIL.n69 11.249
R538 VTAIL.n87 VTAIL.n4 11.249
R539 VTAIL.n128 VTAIL.n116 11.249
R540 VTAIL.n160 VTAIL.n159 11.249
R541 VTAIL.n177 VTAIL.n94 11.249
R542 VTAIL.n220 VTAIL.n208 11.249
R543 VTAIL.n252 VTAIL.n251 11.249
R544 VTAIL.n269 VTAIL.n186 11.249
R545 VTAIL.n633 VTAIL.n550 11.249
R546 VTAIL.n617 VTAIL.n616 11.249
R547 VTAIL.n585 VTAIL.n573 11.249
R548 VTAIL.n541 VTAIL.n458 11.249
R549 VTAIL.n525 VTAIL.n524 11.249
R550 VTAIL.n493 VTAIL.n481 11.249
R551 VTAIL.n451 VTAIL.n368 11.249
R552 VTAIL.n435 VTAIL.n434 11.249
R553 VTAIL.n403 VTAIL.n391 11.249
R554 VTAIL.n359 VTAIL.n276 11.249
R555 VTAIL.n343 VTAIL.n342 11.249
R556 VTAIL.n311 VTAIL.n299 11.249
R557 VTAIL.n678 VTAIL.n677 10.4732
R558 VTAIL.n702 VTAIL.n648 10.4732
R559 VTAIL.n724 VTAIL.n638 10.4732
R560 VTAIL.n42 VTAIL.n41 10.4732
R561 VTAIL.n66 VTAIL.n12 10.4732
R562 VTAIL.n88 VTAIL.n2 10.4732
R563 VTAIL.n132 VTAIL.n131 10.4732
R564 VTAIL.n156 VTAIL.n102 10.4732
R565 VTAIL.n178 VTAIL.n92 10.4732
R566 VTAIL.n224 VTAIL.n223 10.4732
R567 VTAIL.n248 VTAIL.n194 10.4732
R568 VTAIL.n270 VTAIL.n184 10.4732
R569 VTAIL.n634 VTAIL.n548 10.4732
R570 VTAIL.n613 VTAIL.n559 10.4732
R571 VTAIL.n589 VTAIL.n588 10.4732
R572 VTAIL.n542 VTAIL.n456 10.4732
R573 VTAIL.n521 VTAIL.n467 10.4732
R574 VTAIL.n497 VTAIL.n496 10.4732
R575 VTAIL.n452 VTAIL.n366 10.4732
R576 VTAIL.n431 VTAIL.n377 10.4732
R577 VTAIL.n407 VTAIL.n406 10.4732
R578 VTAIL.n360 VTAIL.n274 10.4732
R579 VTAIL.n339 VTAIL.n285 10.4732
R580 VTAIL.n315 VTAIL.n314 10.4732
R581 VTAIL.n681 VTAIL.n660 9.69747
R582 VTAIL.n701 VTAIL.n650 9.69747
R583 VTAIL.n45 VTAIL.n24 9.69747
R584 VTAIL.n65 VTAIL.n14 9.69747
R585 VTAIL.n135 VTAIL.n114 9.69747
R586 VTAIL.n155 VTAIL.n104 9.69747
R587 VTAIL.n227 VTAIL.n206 9.69747
R588 VTAIL.n247 VTAIL.n196 9.69747
R589 VTAIL.n612 VTAIL.n561 9.69747
R590 VTAIL.n592 VTAIL.n571 9.69747
R591 VTAIL.n520 VTAIL.n469 9.69747
R592 VTAIL.n500 VTAIL.n479 9.69747
R593 VTAIL.n430 VTAIL.n379 9.69747
R594 VTAIL.n410 VTAIL.n389 9.69747
R595 VTAIL.n338 VTAIL.n287 9.69747
R596 VTAIL.n318 VTAIL.n297 9.69747
R597 VTAIL.n726 VTAIL.n725 9.45567
R598 VTAIL.n90 VTAIL.n89 9.45567
R599 VTAIL.n180 VTAIL.n179 9.45567
R600 VTAIL.n272 VTAIL.n271 9.45567
R601 VTAIL.n636 VTAIL.n635 9.45567
R602 VTAIL.n544 VTAIL.n543 9.45567
R603 VTAIL.n454 VTAIL.n453 9.45567
R604 VTAIL.n362 VTAIL.n361 9.45567
R605 VTAIL.n725 VTAIL.n724 9.3005
R606 VTAIL.n640 VTAIL.n639 9.3005
R607 VTAIL.n719 VTAIL.n718 9.3005
R608 VTAIL.n717 VTAIL.n716 9.3005
R609 VTAIL.n656 VTAIL.n655 9.3005
R610 VTAIL.n685 VTAIL.n684 9.3005
R611 VTAIL.n683 VTAIL.n682 9.3005
R612 VTAIL.n660 VTAIL.n659 9.3005
R613 VTAIL.n677 VTAIL.n676 9.3005
R614 VTAIL.n675 VTAIL.n674 9.3005
R615 VTAIL.n664 VTAIL.n663 9.3005
R616 VTAIL.n669 VTAIL.n668 9.3005
R617 VTAIL.n691 VTAIL.n690 9.3005
R618 VTAIL.n693 VTAIL.n692 9.3005
R619 VTAIL.n652 VTAIL.n651 9.3005
R620 VTAIL.n699 VTAIL.n698 9.3005
R621 VTAIL.n701 VTAIL.n700 9.3005
R622 VTAIL.n648 VTAIL.n647 9.3005
R623 VTAIL.n707 VTAIL.n706 9.3005
R624 VTAIL.n709 VTAIL.n708 9.3005
R625 VTAIL.n710 VTAIL.n643 9.3005
R626 VTAIL.n89 VTAIL.n88 9.3005
R627 VTAIL.n4 VTAIL.n3 9.3005
R628 VTAIL.n83 VTAIL.n82 9.3005
R629 VTAIL.n81 VTAIL.n80 9.3005
R630 VTAIL.n20 VTAIL.n19 9.3005
R631 VTAIL.n49 VTAIL.n48 9.3005
R632 VTAIL.n47 VTAIL.n46 9.3005
R633 VTAIL.n24 VTAIL.n23 9.3005
R634 VTAIL.n41 VTAIL.n40 9.3005
R635 VTAIL.n39 VTAIL.n38 9.3005
R636 VTAIL.n28 VTAIL.n27 9.3005
R637 VTAIL.n33 VTAIL.n32 9.3005
R638 VTAIL.n55 VTAIL.n54 9.3005
R639 VTAIL.n57 VTAIL.n56 9.3005
R640 VTAIL.n16 VTAIL.n15 9.3005
R641 VTAIL.n63 VTAIL.n62 9.3005
R642 VTAIL.n65 VTAIL.n64 9.3005
R643 VTAIL.n12 VTAIL.n11 9.3005
R644 VTAIL.n71 VTAIL.n70 9.3005
R645 VTAIL.n73 VTAIL.n72 9.3005
R646 VTAIL.n74 VTAIL.n7 9.3005
R647 VTAIL.n179 VTAIL.n178 9.3005
R648 VTAIL.n94 VTAIL.n93 9.3005
R649 VTAIL.n173 VTAIL.n172 9.3005
R650 VTAIL.n171 VTAIL.n170 9.3005
R651 VTAIL.n110 VTAIL.n109 9.3005
R652 VTAIL.n139 VTAIL.n138 9.3005
R653 VTAIL.n137 VTAIL.n136 9.3005
R654 VTAIL.n114 VTAIL.n113 9.3005
R655 VTAIL.n131 VTAIL.n130 9.3005
R656 VTAIL.n129 VTAIL.n128 9.3005
R657 VTAIL.n118 VTAIL.n117 9.3005
R658 VTAIL.n123 VTAIL.n122 9.3005
R659 VTAIL.n145 VTAIL.n144 9.3005
R660 VTAIL.n147 VTAIL.n146 9.3005
R661 VTAIL.n106 VTAIL.n105 9.3005
R662 VTAIL.n153 VTAIL.n152 9.3005
R663 VTAIL.n155 VTAIL.n154 9.3005
R664 VTAIL.n102 VTAIL.n101 9.3005
R665 VTAIL.n161 VTAIL.n160 9.3005
R666 VTAIL.n163 VTAIL.n162 9.3005
R667 VTAIL.n164 VTAIL.n97 9.3005
R668 VTAIL.n271 VTAIL.n270 9.3005
R669 VTAIL.n186 VTAIL.n185 9.3005
R670 VTAIL.n265 VTAIL.n264 9.3005
R671 VTAIL.n263 VTAIL.n262 9.3005
R672 VTAIL.n202 VTAIL.n201 9.3005
R673 VTAIL.n231 VTAIL.n230 9.3005
R674 VTAIL.n229 VTAIL.n228 9.3005
R675 VTAIL.n206 VTAIL.n205 9.3005
R676 VTAIL.n223 VTAIL.n222 9.3005
R677 VTAIL.n221 VTAIL.n220 9.3005
R678 VTAIL.n210 VTAIL.n209 9.3005
R679 VTAIL.n215 VTAIL.n214 9.3005
R680 VTAIL.n237 VTAIL.n236 9.3005
R681 VTAIL.n239 VTAIL.n238 9.3005
R682 VTAIL.n198 VTAIL.n197 9.3005
R683 VTAIL.n245 VTAIL.n244 9.3005
R684 VTAIL.n247 VTAIL.n246 9.3005
R685 VTAIL.n194 VTAIL.n193 9.3005
R686 VTAIL.n253 VTAIL.n252 9.3005
R687 VTAIL.n255 VTAIL.n254 9.3005
R688 VTAIL.n256 VTAIL.n189 9.3005
R689 VTAIL.n604 VTAIL.n603 9.3005
R690 VTAIL.n563 VTAIL.n562 9.3005
R691 VTAIL.n610 VTAIL.n609 9.3005
R692 VTAIL.n612 VTAIL.n611 9.3005
R693 VTAIL.n559 VTAIL.n558 9.3005
R694 VTAIL.n618 VTAIL.n617 9.3005
R695 VTAIL.n620 VTAIL.n619 9.3005
R696 VTAIL.n556 VTAIL.n553 9.3005
R697 VTAIL.n635 VTAIL.n634 9.3005
R698 VTAIL.n550 VTAIL.n549 9.3005
R699 VTAIL.n629 VTAIL.n628 9.3005
R700 VTAIL.n627 VTAIL.n626 9.3005
R701 VTAIL.n602 VTAIL.n601 9.3005
R702 VTAIL.n567 VTAIL.n566 9.3005
R703 VTAIL.n596 VTAIL.n595 9.3005
R704 VTAIL.n594 VTAIL.n593 9.3005
R705 VTAIL.n571 VTAIL.n570 9.3005
R706 VTAIL.n588 VTAIL.n587 9.3005
R707 VTAIL.n586 VTAIL.n585 9.3005
R708 VTAIL.n575 VTAIL.n574 9.3005
R709 VTAIL.n580 VTAIL.n579 9.3005
R710 VTAIL.n512 VTAIL.n511 9.3005
R711 VTAIL.n471 VTAIL.n470 9.3005
R712 VTAIL.n518 VTAIL.n517 9.3005
R713 VTAIL.n520 VTAIL.n519 9.3005
R714 VTAIL.n467 VTAIL.n466 9.3005
R715 VTAIL.n526 VTAIL.n525 9.3005
R716 VTAIL.n528 VTAIL.n527 9.3005
R717 VTAIL.n464 VTAIL.n461 9.3005
R718 VTAIL.n543 VTAIL.n542 9.3005
R719 VTAIL.n458 VTAIL.n457 9.3005
R720 VTAIL.n537 VTAIL.n536 9.3005
R721 VTAIL.n535 VTAIL.n534 9.3005
R722 VTAIL.n510 VTAIL.n509 9.3005
R723 VTAIL.n475 VTAIL.n474 9.3005
R724 VTAIL.n504 VTAIL.n503 9.3005
R725 VTAIL.n502 VTAIL.n501 9.3005
R726 VTAIL.n479 VTAIL.n478 9.3005
R727 VTAIL.n496 VTAIL.n495 9.3005
R728 VTAIL.n494 VTAIL.n493 9.3005
R729 VTAIL.n483 VTAIL.n482 9.3005
R730 VTAIL.n488 VTAIL.n487 9.3005
R731 VTAIL.n422 VTAIL.n421 9.3005
R732 VTAIL.n381 VTAIL.n380 9.3005
R733 VTAIL.n428 VTAIL.n427 9.3005
R734 VTAIL.n430 VTAIL.n429 9.3005
R735 VTAIL.n377 VTAIL.n376 9.3005
R736 VTAIL.n436 VTAIL.n435 9.3005
R737 VTAIL.n438 VTAIL.n437 9.3005
R738 VTAIL.n374 VTAIL.n371 9.3005
R739 VTAIL.n453 VTAIL.n452 9.3005
R740 VTAIL.n368 VTAIL.n367 9.3005
R741 VTAIL.n447 VTAIL.n446 9.3005
R742 VTAIL.n445 VTAIL.n444 9.3005
R743 VTAIL.n420 VTAIL.n419 9.3005
R744 VTAIL.n385 VTAIL.n384 9.3005
R745 VTAIL.n414 VTAIL.n413 9.3005
R746 VTAIL.n412 VTAIL.n411 9.3005
R747 VTAIL.n389 VTAIL.n388 9.3005
R748 VTAIL.n406 VTAIL.n405 9.3005
R749 VTAIL.n404 VTAIL.n403 9.3005
R750 VTAIL.n393 VTAIL.n392 9.3005
R751 VTAIL.n398 VTAIL.n397 9.3005
R752 VTAIL.n330 VTAIL.n329 9.3005
R753 VTAIL.n289 VTAIL.n288 9.3005
R754 VTAIL.n336 VTAIL.n335 9.3005
R755 VTAIL.n338 VTAIL.n337 9.3005
R756 VTAIL.n285 VTAIL.n284 9.3005
R757 VTAIL.n344 VTAIL.n343 9.3005
R758 VTAIL.n346 VTAIL.n345 9.3005
R759 VTAIL.n282 VTAIL.n279 9.3005
R760 VTAIL.n361 VTAIL.n360 9.3005
R761 VTAIL.n276 VTAIL.n275 9.3005
R762 VTAIL.n355 VTAIL.n354 9.3005
R763 VTAIL.n353 VTAIL.n352 9.3005
R764 VTAIL.n328 VTAIL.n327 9.3005
R765 VTAIL.n293 VTAIL.n292 9.3005
R766 VTAIL.n322 VTAIL.n321 9.3005
R767 VTAIL.n320 VTAIL.n319 9.3005
R768 VTAIL.n297 VTAIL.n296 9.3005
R769 VTAIL.n314 VTAIL.n313 9.3005
R770 VTAIL.n312 VTAIL.n311 9.3005
R771 VTAIL.n301 VTAIL.n300 9.3005
R772 VTAIL.n306 VTAIL.n305 9.3005
R773 VTAIL.n682 VTAIL.n658 8.92171
R774 VTAIL.n698 VTAIL.n697 8.92171
R775 VTAIL.n46 VTAIL.n22 8.92171
R776 VTAIL.n62 VTAIL.n61 8.92171
R777 VTAIL.n136 VTAIL.n112 8.92171
R778 VTAIL.n152 VTAIL.n151 8.92171
R779 VTAIL.n228 VTAIL.n204 8.92171
R780 VTAIL.n244 VTAIL.n243 8.92171
R781 VTAIL.n609 VTAIL.n608 8.92171
R782 VTAIL.n593 VTAIL.n569 8.92171
R783 VTAIL.n517 VTAIL.n516 8.92171
R784 VTAIL.n501 VTAIL.n477 8.92171
R785 VTAIL.n427 VTAIL.n426 8.92171
R786 VTAIL.n411 VTAIL.n387 8.92171
R787 VTAIL.n335 VTAIL.n334 8.92171
R788 VTAIL.n319 VTAIL.n295 8.92171
R789 VTAIL.n686 VTAIL.n685 8.14595
R790 VTAIL.n694 VTAIL.n652 8.14595
R791 VTAIL.n50 VTAIL.n49 8.14595
R792 VTAIL.n58 VTAIL.n16 8.14595
R793 VTAIL.n140 VTAIL.n139 8.14595
R794 VTAIL.n148 VTAIL.n106 8.14595
R795 VTAIL.n232 VTAIL.n231 8.14595
R796 VTAIL.n240 VTAIL.n198 8.14595
R797 VTAIL.n605 VTAIL.n563 8.14595
R798 VTAIL.n597 VTAIL.n596 8.14595
R799 VTAIL.n513 VTAIL.n471 8.14595
R800 VTAIL.n505 VTAIL.n504 8.14595
R801 VTAIL.n423 VTAIL.n381 8.14595
R802 VTAIL.n415 VTAIL.n414 8.14595
R803 VTAIL.n331 VTAIL.n289 8.14595
R804 VTAIL.n323 VTAIL.n322 8.14595
R805 VTAIL.n689 VTAIL.n656 7.3702
R806 VTAIL.n693 VTAIL.n654 7.3702
R807 VTAIL.n53 VTAIL.n20 7.3702
R808 VTAIL.n57 VTAIL.n18 7.3702
R809 VTAIL.n143 VTAIL.n110 7.3702
R810 VTAIL.n147 VTAIL.n108 7.3702
R811 VTAIL.n235 VTAIL.n202 7.3702
R812 VTAIL.n239 VTAIL.n200 7.3702
R813 VTAIL.n604 VTAIL.n565 7.3702
R814 VTAIL.n600 VTAIL.n567 7.3702
R815 VTAIL.n512 VTAIL.n473 7.3702
R816 VTAIL.n508 VTAIL.n475 7.3702
R817 VTAIL.n422 VTAIL.n383 7.3702
R818 VTAIL.n418 VTAIL.n385 7.3702
R819 VTAIL.n330 VTAIL.n291 7.3702
R820 VTAIL.n326 VTAIL.n293 7.3702
R821 VTAIL.n690 VTAIL.n689 6.59444
R822 VTAIL.n690 VTAIL.n654 6.59444
R823 VTAIL.n54 VTAIL.n53 6.59444
R824 VTAIL.n54 VTAIL.n18 6.59444
R825 VTAIL.n144 VTAIL.n143 6.59444
R826 VTAIL.n144 VTAIL.n108 6.59444
R827 VTAIL.n236 VTAIL.n235 6.59444
R828 VTAIL.n236 VTAIL.n200 6.59444
R829 VTAIL.n601 VTAIL.n565 6.59444
R830 VTAIL.n601 VTAIL.n600 6.59444
R831 VTAIL.n509 VTAIL.n473 6.59444
R832 VTAIL.n509 VTAIL.n508 6.59444
R833 VTAIL.n419 VTAIL.n383 6.59444
R834 VTAIL.n419 VTAIL.n418 6.59444
R835 VTAIL.n327 VTAIL.n291 6.59444
R836 VTAIL.n327 VTAIL.n326 6.59444
R837 VTAIL.n686 VTAIL.n656 5.81868
R838 VTAIL.n694 VTAIL.n693 5.81868
R839 VTAIL.n50 VTAIL.n20 5.81868
R840 VTAIL.n58 VTAIL.n57 5.81868
R841 VTAIL.n140 VTAIL.n110 5.81868
R842 VTAIL.n148 VTAIL.n147 5.81868
R843 VTAIL.n232 VTAIL.n202 5.81868
R844 VTAIL.n240 VTAIL.n239 5.81868
R845 VTAIL.n605 VTAIL.n604 5.81868
R846 VTAIL.n597 VTAIL.n567 5.81868
R847 VTAIL.n513 VTAIL.n512 5.81868
R848 VTAIL.n505 VTAIL.n475 5.81868
R849 VTAIL.n423 VTAIL.n422 5.81868
R850 VTAIL.n415 VTAIL.n385 5.81868
R851 VTAIL.n331 VTAIL.n330 5.81868
R852 VTAIL.n323 VTAIL.n293 5.81868
R853 VTAIL.n685 VTAIL.n658 5.04292
R854 VTAIL.n697 VTAIL.n652 5.04292
R855 VTAIL.n49 VTAIL.n22 5.04292
R856 VTAIL.n61 VTAIL.n16 5.04292
R857 VTAIL.n139 VTAIL.n112 5.04292
R858 VTAIL.n151 VTAIL.n106 5.04292
R859 VTAIL.n231 VTAIL.n204 5.04292
R860 VTAIL.n243 VTAIL.n198 5.04292
R861 VTAIL.n608 VTAIL.n563 5.04292
R862 VTAIL.n596 VTAIL.n569 5.04292
R863 VTAIL.n516 VTAIL.n471 5.04292
R864 VTAIL.n504 VTAIL.n477 5.04292
R865 VTAIL.n426 VTAIL.n381 5.04292
R866 VTAIL.n414 VTAIL.n387 5.04292
R867 VTAIL.n334 VTAIL.n289 5.04292
R868 VTAIL.n322 VTAIL.n295 5.04292
R869 VTAIL.n668 VTAIL.n667 4.38563
R870 VTAIL.n32 VTAIL.n31 4.38563
R871 VTAIL.n122 VTAIL.n121 4.38563
R872 VTAIL.n214 VTAIL.n213 4.38563
R873 VTAIL.n579 VTAIL.n578 4.38563
R874 VTAIL.n487 VTAIL.n486 4.38563
R875 VTAIL.n397 VTAIL.n396 4.38563
R876 VTAIL.n305 VTAIL.n304 4.38563
R877 VTAIL.n682 VTAIL.n681 4.26717
R878 VTAIL.n698 VTAIL.n650 4.26717
R879 VTAIL.n46 VTAIL.n45 4.26717
R880 VTAIL.n62 VTAIL.n14 4.26717
R881 VTAIL.n136 VTAIL.n135 4.26717
R882 VTAIL.n152 VTAIL.n104 4.26717
R883 VTAIL.n228 VTAIL.n227 4.26717
R884 VTAIL.n244 VTAIL.n196 4.26717
R885 VTAIL.n609 VTAIL.n561 4.26717
R886 VTAIL.n593 VTAIL.n592 4.26717
R887 VTAIL.n517 VTAIL.n469 4.26717
R888 VTAIL.n501 VTAIL.n500 4.26717
R889 VTAIL.n427 VTAIL.n379 4.26717
R890 VTAIL.n411 VTAIL.n410 4.26717
R891 VTAIL.n335 VTAIL.n287 4.26717
R892 VTAIL.n319 VTAIL.n318 4.26717
R893 VTAIL.n678 VTAIL.n660 3.49141
R894 VTAIL.n702 VTAIL.n701 3.49141
R895 VTAIL.n726 VTAIL.n638 3.49141
R896 VTAIL.n42 VTAIL.n24 3.49141
R897 VTAIL.n66 VTAIL.n65 3.49141
R898 VTAIL.n90 VTAIL.n2 3.49141
R899 VTAIL.n132 VTAIL.n114 3.49141
R900 VTAIL.n156 VTAIL.n155 3.49141
R901 VTAIL.n180 VTAIL.n92 3.49141
R902 VTAIL.n224 VTAIL.n206 3.49141
R903 VTAIL.n248 VTAIL.n247 3.49141
R904 VTAIL.n272 VTAIL.n184 3.49141
R905 VTAIL.n636 VTAIL.n548 3.49141
R906 VTAIL.n613 VTAIL.n612 3.49141
R907 VTAIL.n589 VTAIL.n571 3.49141
R908 VTAIL.n544 VTAIL.n456 3.49141
R909 VTAIL.n521 VTAIL.n520 3.49141
R910 VTAIL.n497 VTAIL.n479 3.49141
R911 VTAIL.n454 VTAIL.n366 3.49141
R912 VTAIL.n431 VTAIL.n430 3.49141
R913 VTAIL.n407 VTAIL.n389 3.49141
R914 VTAIL.n362 VTAIL.n274 3.49141
R915 VTAIL.n339 VTAIL.n338 3.49141
R916 VTAIL.n315 VTAIL.n297 3.49141
R917 VTAIL.n677 VTAIL.n662 2.71565
R918 VTAIL.n705 VTAIL.n648 2.71565
R919 VTAIL.n724 VTAIL.n723 2.71565
R920 VTAIL.n41 VTAIL.n26 2.71565
R921 VTAIL.n69 VTAIL.n12 2.71565
R922 VTAIL.n88 VTAIL.n87 2.71565
R923 VTAIL.n131 VTAIL.n116 2.71565
R924 VTAIL.n159 VTAIL.n102 2.71565
R925 VTAIL.n178 VTAIL.n177 2.71565
R926 VTAIL.n223 VTAIL.n208 2.71565
R927 VTAIL.n251 VTAIL.n194 2.71565
R928 VTAIL.n270 VTAIL.n269 2.71565
R929 VTAIL.n634 VTAIL.n633 2.71565
R930 VTAIL.n616 VTAIL.n559 2.71565
R931 VTAIL.n588 VTAIL.n573 2.71565
R932 VTAIL.n542 VTAIL.n541 2.71565
R933 VTAIL.n524 VTAIL.n467 2.71565
R934 VTAIL.n496 VTAIL.n481 2.71565
R935 VTAIL.n452 VTAIL.n451 2.71565
R936 VTAIL.n434 VTAIL.n377 2.71565
R937 VTAIL.n406 VTAIL.n391 2.71565
R938 VTAIL.n360 VTAIL.n359 2.71565
R939 VTAIL.n342 VTAIL.n285 2.71565
R940 VTAIL.n314 VTAIL.n299 2.71565
R941 VTAIL.n674 VTAIL.n673 1.93989
R942 VTAIL.n706 VTAIL.n646 1.93989
R943 VTAIL.n720 VTAIL.n640 1.93989
R944 VTAIL.n38 VTAIL.n37 1.93989
R945 VTAIL.n70 VTAIL.n10 1.93989
R946 VTAIL.n84 VTAIL.n4 1.93989
R947 VTAIL.n128 VTAIL.n127 1.93989
R948 VTAIL.n160 VTAIL.n100 1.93989
R949 VTAIL.n174 VTAIL.n94 1.93989
R950 VTAIL.n220 VTAIL.n219 1.93989
R951 VTAIL.n252 VTAIL.n192 1.93989
R952 VTAIL.n266 VTAIL.n186 1.93989
R953 VTAIL.n630 VTAIL.n550 1.93989
R954 VTAIL.n617 VTAIL.n557 1.93989
R955 VTAIL.n585 VTAIL.n584 1.93989
R956 VTAIL.n538 VTAIL.n458 1.93989
R957 VTAIL.n525 VTAIL.n465 1.93989
R958 VTAIL.n493 VTAIL.n492 1.93989
R959 VTAIL.n448 VTAIL.n368 1.93989
R960 VTAIL.n435 VTAIL.n375 1.93989
R961 VTAIL.n403 VTAIL.n402 1.93989
R962 VTAIL.n356 VTAIL.n276 1.93989
R963 VTAIL.n343 VTAIL.n283 1.93989
R964 VTAIL.n311 VTAIL.n310 1.93989
R965 VTAIL.n365 VTAIL.n363 1.76774
R966 VTAIL.n455 VTAIL.n365 1.76774
R967 VTAIL.n547 VTAIL.n545 1.76774
R968 VTAIL.n637 VTAIL.n547 1.76774
R969 VTAIL.n273 VTAIL.n183 1.76774
R970 VTAIL.n183 VTAIL.n181 1.76774
R971 VTAIL.n91 VTAIL.n1 1.76774
R972 VTAIL VTAIL.n727 1.70955
R973 VTAIL.n0 VTAIL.t2 1.22272
R974 VTAIL.n0 VTAIL.t4 1.22272
R975 VTAIL.n182 VTAIL.t9 1.22272
R976 VTAIL.n182 VTAIL.t12 1.22272
R977 VTAIL.n546 VTAIL.t11 1.22272
R978 VTAIL.n546 VTAIL.t14 1.22272
R979 VTAIL.n364 VTAIL.t0 1.22272
R980 VTAIL.n364 VTAIL.t1 1.22272
R981 VTAIL.n670 VTAIL.n664 1.16414
R982 VTAIL.n711 VTAIL.n709 1.16414
R983 VTAIL.n719 VTAIL.n642 1.16414
R984 VTAIL.n34 VTAIL.n28 1.16414
R985 VTAIL.n75 VTAIL.n73 1.16414
R986 VTAIL.n83 VTAIL.n6 1.16414
R987 VTAIL.n124 VTAIL.n118 1.16414
R988 VTAIL.n165 VTAIL.n163 1.16414
R989 VTAIL.n173 VTAIL.n96 1.16414
R990 VTAIL.n216 VTAIL.n210 1.16414
R991 VTAIL.n257 VTAIL.n255 1.16414
R992 VTAIL.n265 VTAIL.n188 1.16414
R993 VTAIL.n629 VTAIL.n552 1.16414
R994 VTAIL.n621 VTAIL.n620 1.16414
R995 VTAIL.n581 VTAIL.n575 1.16414
R996 VTAIL.n537 VTAIL.n460 1.16414
R997 VTAIL.n529 VTAIL.n528 1.16414
R998 VTAIL.n489 VTAIL.n483 1.16414
R999 VTAIL.n447 VTAIL.n370 1.16414
R1000 VTAIL.n439 VTAIL.n438 1.16414
R1001 VTAIL.n399 VTAIL.n393 1.16414
R1002 VTAIL.n355 VTAIL.n278 1.16414
R1003 VTAIL.n347 VTAIL.n346 1.16414
R1004 VTAIL.n307 VTAIL.n301 1.16414
R1005 VTAIL.n545 VTAIL.n455 0.470328
R1006 VTAIL.n181 VTAIL.n91 0.470328
R1007 VTAIL.n669 VTAIL.n666 0.388379
R1008 VTAIL.n710 VTAIL.n644 0.388379
R1009 VTAIL.n716 VTAIL.n715 0.388379
R1010 VTAIL.n33 VTAIL.n30 0.388379
R1011 VTAIL.n74 VTAIL.n8 0.388379
R1012 VTAIL.n80 VTAIL.n79 0.388379
R1013 VTAIL.n123 VTAIL.n120 0.388379
R1014 VTAIL.n164 VTAIL.n98 0.388379
R1015 VTAIL.n170 VTAIL.n169 0.388379
R1016 VTAIL.n215 VTAIL.n212 0.388379
R1017 VTAIL.n256 VTAIL.n190 0.388379
R1018 VTAIL.n262 VTAIL.n261 0.388379
R1019 VTAIL.n626 VTAIL.n625 0.388379
R1020 VTAIL.n556 VTAIL.n554 0.388379
R1021 VTAIL.n580 VTAIL.n577 0.388379
R1022 VTAIL.n534 VTAIL.n533 0.388379
R1023 VTAIL.n464 VTAIL.n462 0.388379
R1024 VTAIL.n488 VTAIL.n485 0.388379
R1025 VTAIL.n444 VTAIL.n443 0.388379
R1026 VTAIL.n374 VTAIL.n372 0.388379
R1027 VTAIL.n398 VTAIL.n395 0.388379
R1028 VTAIL.n352 VTAIL.n351 0.388379
R1029 VTAIL.n282 VTAIL.n280 0.388379
R1030 VTAIL.n306 VTAIL.n303 0.388379
R1031 VTAIL.n668 VTAIL.n663 0.155672
R1032 VTAIL.n675 VTAIL.n663 0.155672
R1033 VTAIL.n676 VTAIL.n675 0.155672
R1034 VTAIL.n676 VTAIL.n659 0.155672
R1035 VTAIL.n683 VTAIL.n659 0.155672
R1036 VTAIL.n684 VTAIL.n683 0.155672
R1037 VTAIL.n684 VTAIL.n655 0.155672
R1038 VTAIL.n691 VTAIL.n655 0.155672
R1039 VTAIL.n692 VTAIL.n691 0.155672
R1040 VTAIL.n692 VTAIL.n651 0.155672
R1041 VTAIL.n699 VTAIL.n651 0.155672
R1042 VTAIL.n700 VTAIL.n699 0.155672
R1043 VTAIL.n700 VTAIL.n647 0.155672
R1044 VTAIL.n707 VTAIL.n647 0.155672
R1045 VTAIL.n708 VTAIL.n707 0.155672
R1046 VTAIL.n708 VTAIL.n643 0.155672
R1047 VTAIL.n717 VTAIL.n643 0.155672
R1048 VTAIL.n718 VTAIL.n717 0.155672
R1049 VTAIL.n718 VTAIL.n639 0.155672
R1050 VTAIL.n725 VTAIL.n639 0.155672
R1051 VTAIL.n32 VTAIL.n27 0.155672
R1052 VTAIL.n39 VTAIL.n27 0.155672
R1053 VTAIL.n40 VTAIL.n39 0.155672
R1054 VTAIL.n40 VTAIL.n23 0.155672
R1055 VTAIL.n47 VTAIL.n23 0.155672
R1056 VTAIL.n48 VTAIL.n47 0.155672
R1057 VTAIL.n48 VTAIL.n19 0.155672
R1058 VTAIL.n55 VTAIL.n19 0.155672
R1059 VTAIL.n56 VTAIL.n55 0.155672
R1060 VTAIL.n56 VTAIL.n15 0.155672
R1061 VTAIL.n63 VTAIL.n15 0.155672
R1062 VTAIL.n64 VTAIL.n63 0.155672
R1063 VTAIL.n64 VTAIL.n11 0.155672
R1064 VTAIL.n71 VTAIL.n11 0.155672
R1065 VTAIL.n72 VTAIL.n71 0.155672
R1066 VTAIL.n72 VTAIL.n7 0.155672
R1067 VTAIL.n81 VTAIL.n7 0.155672
R1068 VTAIL.n82 VTAIL.n81 0.155672
R1069 VTAIL.n82 VTAIL.n3 0.155672
R1070 VTAIL.n89 VTAIL.n3 0.155672
R1071 VTAIL.n122 VTAIL.n117 0.155672
R1072 VTAIL.n129 VTAIL.n117 0.155672
R1073 VTAIL.n130 VTAIL.n129 0.155672
R1074 VTAIL.n130 VTAIL.n113 0.155672
R1075 VTAIL.n137 VTAIL.n113 0.155672
R1076 VTAIL.n138 VTAIL.n137 0.155672
R1077 VTAIL.n138 VTAIL.n109 0.155672
R1078 VTAIL.n145 VTAIL.n109 0.155672
R1079 VTAIL.n146 VTAIL.n145 0.155672
R1080 VTAIL.n146 VTAIL.n105 0.155672
R1081 VTAIL.n153 VTAIL.n105 0.155672
R1082 VTAIL.n154 VTAIL.n153 0.155672
R1083 VTAIL.n154 VTAIL.n101 0.155672
R1084 VTAIL.n161 VTAIL.n101 0.155672
R1085 VTAIL.n162 VTAIL.n161 0.155672
R1086 VTAIL.n162 VTAIL.n97 0.155672
R1087 VTAIL.n171 VTAIL.n97 0.155672
R1088 VTAIL.n172 VTAIL.n171 0.155672
R1089 VTAIL.n172 VTAIL.n93 0.155672
R1090 VTAIL.n179 VTAIL.n93 0.155672
R1091 VTAIL.n214 VTAIL.n209 0.155672
R1092 VTAIL.n221 VTAIL.n209 0.155672
R1093 VTAIL.n222 VTAIL.n221 0.155672
R1094 VTAIL.n222 VTAIL.n205 0.155672
R1095 VTAIL.n229 VTAIL.n205 0.155672
R1096 VTAIL.n230 VTAIL.n229 0.155672
R1097 VTAIL.n230 VTAIL.n201 0.155672
R1098 VTAIL.n237 VTAIL.n201 0.155672
R1099 VTAIL.n238 VTAIL.n237 0.155672
R1100 VTAIL.n238 VTAIL.n197 0.155672
R1101 VTAIL.n245 VTAIL.n197 0.155672
R1102 VTAIL.n246 VTAIL.n245 0.155672
R1103 VTAIL.n246 VTAIL.n193 0.155672
R1104 VTAIL.n253 VTAIL.n193 0.155672
R1105 VTAIL.n254 VTAIL.n253 0.155672
R1106 VTAIL.n254 VTAIL.n189 0.155672
R1107 VTAIL.n263 VTAIL.n189 0.155672
R1108 VTAIL.n264 VTAIL.n263 0.155672
R1109 VTAIL.n264 VTAIL.n185 0.155672
R1110 VTAIL.n271 VTAIL.n185 0.155672
R1111 VTAIL.n635 VTAIL.n549 0.155672
R1112 VTAIL.n628 VTAIL.n549 0.155672
R1113 VTAIL.n628 VTAIL.n627 0.155672
R1114 VTAIL.n627 VTAIL.n553 0.155672
R1115 VTAIL.n619 VTAIL.n553 0.155672
R1116 VTAIL.n619 VTAIL.n618 0.155672
R1117 VTAIL.n618 VTAIL.n558 0.155672
R1118 VTAIL.n611 VTAIL.n558 0.155672
R1119 VTAIL.n611 VTAIL.n610 0.155672
R1120 VTAIL.n610 VTAIL.n562 0.155672
R1121 VTAIL.n603 VTAIL.n562 0.155672
R1122 VTAIL.n603 VTAIL.n602 0.155672
R1123 VTAIL.n602 VTAIL.n566 0.155672
R1124 VTAIL.n595 VTAIL.n566 0.155672
R1125 VTAIL.n595 VTAIL.n594 0.155672
R1126 VTAIL.n594 VTAIL.n570 0.155672
R1127 VTAIL.n587 VTAIL.n570 0.155672
R1128 VTAIL.n587 VTAIL.n586 0.155672
R1129 VTAIL.n586 VTAIL.n574 0.155672
R1130 VTAIL.n579 VTAIL.n574 0.155672
R1131 VTAIL.n543 VTAIL.n457 0.155672
R1132 VTAIL.n536 VTAIL.n457 0.155672
R1133 VTAIL.n536 VTAIL.n535 0.155672
R1134 VTAIL.n535 VTAIL.n461 0.155672
R1135 VTAIL.n527 VTAIL.n461 0.155672
R1136 VTAIL.n527 VTAIL.n526 0.155672
R1137 VTAIL.n526 VTAIL.n466 0.155672
R1138 VTAIL.n519 VTAIL.n466 0.155672
R1139 VTAIL.n519 VTAIL.n518 0.155672
R1140 VTAIL.n518 VTAIL.n470 0.155672
R1141 VTAIL.n511 VTAIL.n470 0.155672
R1142 VTAIL.n511 VTAIL.n510 0.155672
R1143 VTAIL.n510 VTAIL.n474 0.155672
R1144 VTAIL.n503 VTAIL.n474 0.155672
R1145 VTAIL.n503 VTAIL.n502 0.155672
R1146 VTAIL.n502 VTAIL.n478 0.155672
R1147 VTAIL.n495 VTAIL.n478 0.155672
R1148 VTAIL.n495 VTAIL.n494 0.155672
R1149 VTAIL.n494 VTAIL.n482 0.155672
R1150 VTAIL.n487 VTAIL.n482 0.155672
R1151 VTAIL.n453 VTAIL.n367 0.155672
R1152 VTAIL.n446 VTAIL.n367 0.155672
R1153 VTAIL.n446 VTAIL.n445 0.155672
R1154 VTAIL.n445 VTAIL.n371 0.155672
R1155 VTAIL.n437 VTAIL.n371 0.155672
R1156 VTAIL.n437 VTAIL.n436 0.155672
R1157 VTAIL.n436 VTAIL.n376 0.155672
R1158 VTAIL.n429 VTAIL.n376 0.155672
R1159 VTAIL.n429 VTAIL.n428 0.155672
R1160 VTAIL.n428 VTAIL.n380 0.155672
R1161 VTAIL.n421 VTAIL.n380 0.155672
R1162 VTAIL.n421 VTAIL.n420 0.155672
R1163 VTAIL.n420 VTAIL.n384 0.155672
R1164 VTAIL.n413 VTAIL.n384 0.155672
R1165 VTAIL.n413 VTAIL.n412 0.155672
R1166 VTAIL.n412 VTAIL.n388 0.155672
R1167 VTAIL.n405 VTAIL.n388 0.155672
R1168 VTAIL.n405 VTAIL.n404 0.155672
R1169 VTAIL.n404 VTAIL.n392 0.155672
R1170 VTAIL.n397 VTAIL.n392 0.155672
R1171 VTAIL.n361 VTAIL.n275 0.155672
R1172 VTAIL.n354 VTAIL.n275 0.155672
R1173 VTAIL.n354 VTAIL.n353 0.155672
R1174 VTAIL.n353 VTAIL.n279 0.155672
R1175 VTAIL.n345 VTAIL.n279 0.155672
R1176 VTAIL.n345 VTAIL.n344 0.155672
R1177 VTAIL.n344 VTAIL.n284 0.155672
R1178 VTAIL.n337 VTAIL.n284 0.155672
R1179 VTAIL.n337 VTAIL.n336 0.155672
R1180 VTAIL.n336 VTAIL.n288 0.155672
R1181 VTAIL.n329 VTAIL.n288 0.155672
R1182 VTAIL.n329 VTAIL.n328 0.155672
R1183 VTAIL.n328 VTAIL.n292 0.155672
R1184 VTAIL.n321 VTAIL.n292 0.155672
R1185 VTAIL.n321 VTAIL.n320 0.155672
R1186 VTAIL.n320 VTAIL.n296 0.155672
R1187 VTAIL.n313 VTAIL.n296 0.155672
R1188 VTAIL.n313 VTAIL.n312 0.155672
R1189 VTAIL.n312 VTAIL.n300 0.155672
R1190 VTAIL.n305 VTAIL.n300 0.155672
R1191 VTAIL VTAIL.n1 0.0586897
R1192 VDD1 VDD1.n0 64.0468
R1193 VDD1.n3 VDD1.n2 63.9331
R1194 VDD1.n3 VDD1.n1 63.9331
R1195 VDD1.n5 VDD1.n4 63.1048
R1196 VDD1.n5 VDD1.n3 46.2164
R1197 VDD1.n4 VDD1.t4 1.22272
R1198 VDD1.n4 VDD1.t7 1.22272
R1199 VDD1.n0 VDD1.t6 1.22272
R1200 VDD1.n0 VDD1.t2 1.22272
R1201 VDD1.n2 VDD1.t5 1.22272
R1202 VDD1.n2 VDD1.t1 1.22272
R1203 VDD1.n1 VDD1.t0 1.22272
R1204 VDD1.n1 VDD1.t3 1.22272
R1205 VDD1 VDD1.n5 0.825931
R1206 B.n675 B.n674 585
R1207 B.n676 B.n136 585
R1208 B.n678 B.n677 585
R1209 B.n680 B.n135 585
R1210 B.n683 B.n682 585
R1211 B.n684 B.n134 585
R1212 B.n686 B.n685 585
R1213 B.n688 B.n133 585
R1214 B.n691 B.n690 585
R1215 B.n692 B.n132 585
R1216 B.n694 B.n693 585
R1217 B.n696 B.n131 585
R1218 B.n699 B.n698 585
R1219 B.n700 B.n130 585
R1220 B.n702 B.n701 585
R1221 B.n704 B.n129 585
R1222 B.n707 B.n706 585
R1223 B.n708 B.n128 585
R1224 B.n710 B.n709 585
R1225 B.n712 B.n127 585
R1226 B.n715 B.n714 585
R1227 B.n716 B.n126 585
R1228 B.n718 B.n717 585
R1229 B.n720 B.n125 585
R1230 B.n723 B.n722 585
R1231 B.n724 B.n124 585
R1232 B.n726 B.n725 585
R1233 B.n728 B.n123 585
R1234 B.n731 B.n730 585
R1235 B.n732 B.n122 585
R1236 B.n734 B.n733 585
R1237 B.n736 B.n121 585
R1238 B.n739 B.n738 585
R1239 B.n740 B.n120 585
R1240 B.n742 B.n741 585
R1241 B.n744 B.n119 585
R1242 B.n747 B.n746 585
R1243 B.n748 B.n118 585
R1244 B.n750 B.n749 585
R1245 B.n752 B.n117 585
R1246 B.n755 B.n754 585
R1247 B.n756 B.n116 585
R1248 B.n758 B.n757 585
R1249 B.n760 B.n115 585
R1250 B.n763 B.n762 585
R1251 B.n764 B.n114 585
R1252 B.n766 B.n765 585
R1253 B.n768 B.n113 585
R1254 B.n771 B.n770 585
R1255 B.n772 B.n112 585
R1256 B.n774 B.n773 585
R1257 B.n776 B.n111 585
R1258 B.n778 B.n777 585
R1259 B.n780 B.n779 585
R1260 B.n783 B.n782 585
R1261 B.n784 B.n106 585
R1262 B.n786 B.n785 585
R1263 B.n788 B.n105 585
R1264 B.n791 B.n790 585
R1265 B.n792 B.n104 585
R1266 B.n794 B.n793 585
R1267 B.n796 B.n103 585
R1268 B.n798 B.n797 585
R1269 B.n800 B.n799 585
R1270 B.n803 B.n802 585
R1271 B.n804 B.n98 585
R1272 B.n806 B.n805 585
R1273 B.n808 B.n97 585
R1274 B.n811 B.n810 585
R1275 B.n812 B.n96 585
R1276 B.n814 B.n813 585
R1277 B.n816 B.n95 585
R1278 B.n819 B.n818 585
R1279 B.n820 B.n94 585
R1280 B.n822 B.n821 585
R1281 B.n824 B.n93 585
R1282 B.n827 B.n826 585
R1283 B.n828 B.n92 585
R1284 B.n830 B.n829 585
R1285 B.n832 B.n91 585
R1286 B.n835 B.n834 585
R1287 B.n836 B.n90 585
R1288 B.n838 B.n837 585
R1289 B.n840 B.n89 585
R1290 B.n843 B.n842 585
R1291 B.n844 B.n88 585
R1292 B.n846 B.n845 585
R1293 B.n848 B.n87 585
R1294 B.n851 B.n850 585
R1295 B.n852 B.n86 585
R1296 B.n854 B.n853 585
R1297 B.n856 B.n85 585
R1298 B.n859 B.n858 585
R1299 B.n860 B.n84 585
R1300 B.n862 B.n861 585
R1301 B.n864 B.n83 585
R1302 B.n867 B.n866 585
R1303 B.n868 B.n82 585
R1304 B.n870 B.n869 585
R1305 B.n872 B.n81 585
R1306 B.n875 B.n874 585
R1307 B.n876 B.n80 585
R1308 B.n878 B.n877 585
R1309 B.n880 B.n79 585
R1310 B.n883 B.n882 585
R1311 B.n884 B.n78 585
R1312 B.n886 B.n885 585
R1313 B.n888 B.n77 585
R1314 B.n891 B.n890 585
R1315 B.n892 B.n76 585
R1316 B.n894 B.n893 585
R1317 B.n896 B.n75 585
R1318 B.n899 B.n898 585
R1319 B.n900 B.n74 585
R1320 B.n902 B.n901 585
R1321 B.n904 B.n73 585
R1322 B.n907 B.n906 585
R1323 B.n908 B.n72 585
R1324 B.n672 B.n70 585
R1325 B.n911 B.n70 585
R1326 B.n671 B.n69 585
R1327 B.n912 B.n69 585
R1328 B.n670 B.n68 585
R1329 B.n913 B.n68 585
R1330 B.n669 B.n668 585
R1331 B.n668 B.n64 585
R1332 B.n667 B.n63 585
R1333 B.n919 B.n63 585
R1334 B.n666 B.n62 585
R1335 B.n920 B.n62 585
R1336 B.n665 B.n61 585
R1337 B.n921 B.n61 585
R1338 B.n664 B.n663 585
R1339 B.n663 B.n57 585
R1340 B.n662 B.n56 585
R1341 B.n927 B.n56 585
R1342 B.n661 B.n55 585
R1343 B.n928 B.n55 585
R1344 B.n660 B.n54 585
R1345 B.n929 B.n54 585
R1346 B.n659 B.n658 585
R1347 B.n658 B.n50 585
R1348 B.n657 B.n49 585
R1349 B.n935 B.n49 585
R1350 B.n656 B.n48 585
R1351 B.n936 B.n48 585
R1352 B.n655 B.n47 585
R1353 B.n937 B.n47 585
R1354 B.n654 B.n653 585
R1355 B.n653 B.n46 585
R1356 B.n652 B.n42 585
R1357 B.n943 B.n42 585
R1358 B.n651 B.n41 585
R1359 B.n944 B.n41 585
R1360 B.n650 B.n40 585
R1361 B.n945 B.n40 585
R1362 B.n649 B.n648 585
R1363 B.n648 B.n36 585
R1364 B.n647 B.n35 585
R1365 B.n951 B.n35 585
R1366 B.n646 B.n34 585
R1367 B.n952 B.n34 585
R1368 B.n645 B.n33 585
R1369 B.n953 B.n33 585
R1370 B.n644 B.n643 585
R1371 B.n643 B.n29 585
R1372 B.n642 B.n28 585
R1373 B.n959 B.n28 585
R1374 B.n641 B.n27 585
R1375 B.n960 B.n27 585
R1376 B.n640 B.n26 585
R1377 B.n961 B.n26 585
R1378 B.n639 B.n638 585
R1379 B.n638 B.n25 585
R1380 B.n637 B.n21 585
R1381 B.n967 B.n21 585
R1382 B.n636 B.n20 585
R1383 B.n968 B.n20 585
R1384 B.n635 B.n19 585
R1385 B.n969 B.n19 585
R1386 B.n634 B.n633 585
R1387 B.n633 B.n15 585
R1388 B.n632 B.n14 585
R1389 B.n975 B.n14 585
R1390 B.n631 B.n13 585
R1391 B.n976 B.n13 585
R1392 B.n630 B.n12 585
R1393 B.n977 B.n12 585
R1394 B.n629 B.n628 585
R1395 B.n628 B.n8 585
R1396 B.n627 B.n7 585
R1397 B.n983 B.n7 585
R1398 B.n626 B.n6 585
R1399 B.n984 B.n6 585
R1400 B.n625 B.n5 585
R1401 B.n985 B.n5 585
R1402 B.n624 B.n623 585
R1403 B.n623 B.n4 585
R1404 B.n622 B.n137 585
R1405 B.n622 B.n621 585
R1406 B.n612 B.n138 585
R1407 B.n139 B.n138 585
R1408 B.n614 B.n613 585
R1409 B.n615 B.n614 585
R1410 B.n611 B.n143 585
R1411 B.n147 B.n143 585
R1412 B.n610 B.n609 585
R1413 B.n609 B.n608 585
R1414 B.n145 B.n144 585
R1415 B.n146 B.n145 585
R1416 B.n601 B.n600 585
R1417 B.n602 B.n601 585
R1418 B.n599 B.n152 585
R1419 B.n152 B.n151 585
R1420 B.n598 B.n597 585
R1421 B.n597 B.n596 585
R1422 B.n154 B.n153 585
R1423 B.n589 B.n154 585
R1424 B.n588 B.n587 585
R1425 B.n590 B.n588 585
R1426 B.n586 B.n159 585
R1427 B.n159 B.n158 585
R1428 B.n585 B.n584 585
R1429 B.n584 B.n583 585
R1430 B.n161 B.n160 585
R1431 B.n162 B.n161 585
R1432 B.n576 B.n575 585
R1433 B.n577 B.n576 585
R1434 B.n574 B.n166 585
R1435 B.n170 B.n166 585
R1436 B.n573 B.n572 585
R1437 B.n572 B.n571 585
R1438 B.n168 B.n167 585
R1439 B.n169 B.n168 585
R1440 B.n564 B.n563 585
R1441 B.n565 B.n564 585
R1442 B.n562 B.n175 585
R1443 B.n175 B.n174 585
R1444 B.n561 B.n560 585
R1445 B.n560 B.n559 585
R1446 B.n177 B.n176 585
R1447 B.n552 B.n177 585
R1448 B.n551 B.n550 585
R1449 B.n553 B.n551 585
R1450 B.n549 B.n182 585
R1451 B.n182 B.n181 585
R1452 B.n548 B.n547 585
R1453 B.n547 B.n546 585
R1454 B.n184 B.n183 585
R1455 B.n185 B.n184 585
R1456 B.n539 B.n538 585
R1457 B.n540 B.n539 585
R1458 B.n537 B.n190 585
R1459 B.n190 B.n189 585
R1460 B.n536 B.n535 585
R1461 B.n535 B.n534 585
R1462 B.n192 B.n191 585
R1463 B.n193 B.n192 585
R1464 B.n527 B.n526 585
R1465 B.n528 B.n527 585
R1466 B.n525 B.n198 585
R1467 B.n198 B.n197 585
R1468 B.n524 B.n523 585
R1469 B.n523 B.n522 585
R1470 B.n200 B.n199 585
R1471 B.n201 B.n200 585
R1472 B.n515 B.n514 585
R1473 B.n516 B.n515 585
R1474 B.n513 B.n206 585
R1475 B.n206 B.n205 585
R1476 B.n512 B.n511 585
R1477 B.n511 B.n510 585
R1478 B.n507 B.n210 585
R1479 B.n506 B.n505 585
R1480 B.n503 B.n211 585
R1481 B.n503 B.n209 585
R1482 B.n502 B.n501 585
R1483 B.n500 B.n499 585
R1484 B.n498 B.n213 585
R1485 B.n496 B.n495 585
R1486 B.n494 B.n214 585
R1487 B.n493 B.n492 585
R1488 B.n490 B.n215 585
R1489 B.n488 B.n487 585
R1490 B.n486 B.n216 585
R1491 B.n485 B.n484 585
R1492 B.n482 B.n217 585
R1493 B.n480 B.n479 585
R1494 B.n478 B.n218 585
R1495 B.n477 B.n476 585
R1496 B.n474 B.n219 585
R1497 B.n472 B.n471 585
R1498 B.n470 B.n220 585
R1499 B.n469 B.n468 585
R1500 B.n466 B.n221 585
R1501 B.n464 B.n463 585
R1502 B.n462 B.n222 585
R1503 B.n461 B.n460 585
R1504 B.n458 B.n223 585
R1505 B.n456 B.n455 585
R1506 B.n454 B.n224 585
R1507 B.n453 B.n452 585
R1508 B.n450 B.n225 585
R1509 B.n448 B.n447 585
R1510 B.n446 B.n226 585
R1511 B.n445 B.n444 585
R1512 B.n442 B.n227 585
R1513 B.n440 B.n439 585
R1514 B.n438 B.n228 585
R1515 B.n437 B.n436 585
R1516 B.n434 B.n229 585
R1517 B.n432 B.n431 585
R1518 B.n430 B.n230 585
R1519 B.n429 B.n428 585
R1520 B.n426 B.n231 585
R1521 B.n424 B.n423 585
R1522 B.n422 B.n232 585
R1523 B.n421 B.n420 585
R1524 B.n418 B.n233 585
R1525 B.n416 B.n415 585
R1526 B.n414 B.n234 585
R1527 B.n413 B.n412 585
R1528 B.n410 B.n235 585
R1529 B.n408 B.n407 585
R1530 B.n406 B.n236 585
R1531 B.n405 B.n404 585
R1532 B.n402 B.n237 585
R1533 B.n400 B.n399 585
R1534 B.n398 B.n238 585
R1535 B.n397 B.n396 585
R1536 B.n394 B.n242 585
R1537 B.n392 B.n391 585
R1538 B.n390 B.n243 585
R1539 B.n389 B.n388 585
R1540 B.n386 B.n244 585
R1541 B.n384 B.n383 585
R1542 B.n382 B.n245 585
R1543 B.n380 B.n379 585
R1544 B.n377 B.n248 585
R1545 B.n375 B.n374 585
R1546 B.n373 B.n249 585
R1547 B.n372 B.n371 585
R1548 B.n369 B.n250 585
R1549 B.n367 B.n366 585
R1550 B.n365 B.n251 585
R1551 B.n364 B.n363 585
R1552 B.n361 B.n252 585
R1553 B.n359 B.n358 585
R1554 B.n357 B.n253 585
R1555 B.n356 B.n355 585
R1556 B.n353 B.n254 585
R1557 B.n351 B.n350 585
R1558 B.n349 B.n255 585
R1559 B.n348 B.n347 585
R1560 B.n345 B.n256 585
R1561 B.n343 B.n342 585
R1562 B.n341 B.n257 585
R1563 B.n340 B.n339 585
R1564 B.n337 B.n258 585
R1565 B.n335 B.n334 585
R1566 B.n333 B.n259 585
R1567 B.n332 B.n331 585
R1568 B.n329 B.n260 585
R1569 B.n327 B.n326 585
R1570 B.n325 B.n261 585
R1571 B.n324 B.n323 585
R1572 B.n321 B.n262 585
R1573 B.n319 B.n318 585
R1574 B.n317 B.n263 585
R1575 B.n316 B.n315 585
R1576 B.n313 B.n264 585
R1577 B.n311 B.n310 585
R1578 B.n309 B.n265 585
R1579 B.n308 B.n307 585
R1580 B.n305 B.n266 585
R1581 B.n303 B.n302 585
R1582 B.n301 B.n267 585
R1583 B.n300 B.n299 585
R1584 B.n297 B.n268 585
R1585 B.n295 B.n294 585
R1586 B.n293 B.n269 585
R1587 B.n292 B.n291 585
R1588 B.n289 B.n270 585
R1589 B.n287 B.n286 585
R1590 B.n285 B.n271 585
R1591 B.n284 B.n283 585
R1592 B.n281 B.n272 585
R1593 B.n279 B.n278 585
R1594 B.n277 B.n273 585
R1595 B.n276 B.n275 585
R1596 B.n208 B.n207 585
R1597 B.n209 B.n208 585
R1598 B.n509 B.n508 585
R1599 B.n510 B.n509 585
R1600 B.n204 B.n203 585
R1601 B.n205 B.n204 585
R1602 B.n518 B.n517 585
R1603 B.n517 B.n516 585
R1604 B.n519 B.n202 585
R1605 B.n202 B.n201 585
R1606 B.n521 B.n520 585
R1607 B.n522 B.n521 585
R1608 B.n196 B.n195 585
R1609 B.n197 B.n196 585
R1610 B.n530 B.n529 585
R1611 B.n529 B.n528 585
R1612 B.n531 B.n194 585
R1613 B.n194 B.n193 585
R1614 B.n533 B.n532 585
R1615 B.n534 B.n533 585
R1616 B.n188 B.n187 585
R1617 B.n189 B.n188 585
R1618 B.n542 B.n541 585
R1619 B.n541 B.n540 585
R1620 B.n543 B.n186 585
R1621 B.n186 B.n185 585
R1622 B.n545 B.n544 585
R1623 B.n546 B.n545 585
R1624 B.n180 B.n179 585
R1625 B.n181 B.n180 585
R1626 B.n555 B.n554 585
R1627 B.n554 B.n553 585
R1628 B.n556 B.n178 585
R1629 B.n552 B.n178 585
R1630 B.n558 B.n557 585
R1631 B.n559 B.n558 585
R1632 B.n173 B.n172 585
R1633 B.n174 B.n173 585
R1634 B.n567 B.n566 585
R1635 B.n566 B.n565 585
R1636 B.n568 B.n171 585
R1637 B.n171 B.n169 585
R1638 B.n570 B.n569 585
R1639 B.n571 B.n570 585
R1640 B.n165 B.n164 585
R1641 B.n170 B.n165 585
R1642 B.n579 B.n578 585
R1643 B.n578 B.n577 585
R1644 B.n580 B.n163 585
R1645 B.n163 B.n162 585
R1646 B.n582 B.n581 585
R1647 B.n583 B.n582 585
R1648 B.n157 B.n156 585
R1649 B.n158 B.n157 585
R1650 B.n592 B.n591 585
R1651 B.n591 B.n590 585
R1652 B.n593 B.n155 585
R1653 B.n589 B.n155 585
R1654 B.n595 B.n594 585
R1655 B.n596 B.n595 585
R1656 B.n150 B.n149 585
R1657 B.n151 B.n150 585
R1658 B.n604 B.n603 585
R1659 B.n603 B.n602 585
R1660 B.n605 B.n148 585
R1661 B.n148 B.n146 585
R1662 B.n607 B.n606 585
R1663 B.n608 B.n607 585
R1664 B.n142 B.n141 585
R1665 B.n147 B.n142 585
R1666 B.n617 B.n616 585
R1667 B.n616 B.n615 585
R1668 B.n618 B.n140 585
R1669 B.n140 B.n139 585
R1670 B.n620 B.n619 585
R1671 B.n621 B.n620 585
R1672 B.n2 B.n0 585
R1673 B.n4 B.n2 585
R1674 B.n3 B.n1 585
R1675 B.n984 B.n3 585
R1676 B.n982 B.n981 585
R1677 B.n983 B.n982 585
R1678 B.n980 B.n9 585
R1679 B.n9 B.n8 585
R1680 B.n979 B.n978 585
R1681 B.n978 B.n977 585
R1682 B.n11 B.n10 585
R1683 B.n976 B.n11 585
R1684 B.n974 B.n973 585
R1685 B.n975 B.n974 585
R1686 B.n972 B.n16 585
R1687 B.n16 B.n15 585
R1688 B.n971 B.n970 585
R1689 B.n970 B.n969 585
R1690 B.n18 B.n17 585
R1691 B.n968 B.n18 585
R1692 B.n966 B.n965 585
R1693 B.n967 B.n966 585
R1694 B.n964 B.n22 585
R1695 B.n25 B.n22 585
R1696 B.n963 B.n962 585
R1697 B.n962 B.n961 585
R1698 B.n24 B.n23 585
R1699 B.n960 B.n24 585
R1700 B.n958 B.n957 585
R1701 B.n959 B.n958 585
R1702 B.n956 B.n30 585
R1703 B.n30 B.n29 585
R1704 B.n955 B.n954 585
R1705 B.n954 B.n953 585
R1706 B.n32 B.n31 585
R1707 B.n952 B.n32 585
R1708 B.n950 B.n949 585
R1709 B.n951 B.n950 585
R1710 B.n948 B.n37 585
R1711 B.n37 B.n36 585
R1712 B.n947 B.n946 585
R1713 B.n946 B.n945 585
R1714 B.n39 B.n38 585
R1715 B.n944 B.n39 585
R1716 B.n942 B.n941 585
R1717 B.n943 B.n942 585
R1718 B.n940 B.n43 585
R1719 B.n46 B.n43 585
R1720 B.n939 B.n938 585
R1721 B.n938 B.n937 585
R1722 B.n45 B.n44 585
R1723 B.n936 B.n45 585
R1724 B.n934 B.n933 585
R1725 B.n935 B.n934 585
R1726 B.n932 B.n51 585
R1727 B.n51 B.n50 585
R1728 B.n931 B.n930 585
R1729 B.n930 B.n929 585
R1730 B.n53 B.n52 585
R1731 B.n928 B.n53 585
R1732 B.n926 B.n925 585
R1733 B.n927 B.n926 585
R1734 B.n924 B.n58 585
R1735 B.n58 B.n57 585
R1736 B.n923 B.n922 585
R1737 B.n922 B.n921 585
R1738 B.n60 B.n59 585
R1739 B.n920 B.n60 585
R1740 B.n918 B.n917 585
R1741 B.n919 B.n918 585
R1742 B.n916 B.n65 585
R1743 B.n65 B.n64 585
R1744 B.n915 B.n914 585
R1745 B.n914 B.n913 585
R1746 B.n67 B.n66 585
R1747 B.n912 B.n67 585
R1748 B.n910 B.n909 585
R1749 B.n911 B.n910 585
R1750 B.n987 B.n986 585
R1751 B.n986 B.n985 585
R1752 B.n509 B.n210 502.111
R1753 B.n910 B.n72 502.111
R1754 B.n511 B.n208 502.111
R1755 B.n674 B.n70 502.111
R1756 B.n246 B.t15 433.163
R1757 B.n239 B.t19 433.163
R1758 B.n99 B.t8 433.163
R1759 B.n107 B.t12 433.163
R1760 B.n246 B.t18 394.368
R1761 B.n239 B.t21 394.368
R1762 B.n99 B.t10 394.368
R1763 B.n107 B.t13 394.368
R1764 B.n247 B.t17 354.61
R1765 B.n108 B.t14 354.61
R1766 B.n240 B.t20 354.61
R1767 B.n100 B.t11 354.61
R1768 B.n673 B.n71 256.663
R1769 B.n679 B.n71 256.663
R1770 B.n681 B.n71 256.663
R1771 B.n687 B.n71 256.663
R1772 B.n689 B.n71 256.663
R1773 B.n695 B.n71 256.663
R1774 B.n697 B.n71 256.663
R1775 B.n703 B.n71 256.663
R1776 B.n705 B.n71 256.663
R1777 B.n711 B.n71 256.663
R1778 B.n713 B.n71 256.663
R1779 B.n719 B.n71 256.663
R1780 B.n721 B.n71 256.663
R1781 B.n727 B.n71 256.663
R1782 B.n729 B.n71 256.663
R1783 B.n735 B.n71 256.663
R1784 B.n737 B.n71 256.663
R1785 B.n743 B.n71 256.663
R1786 B.n745 B.n71 256.663
R1787 B.n751 B.n71 256.663
R1788 B.n753 B.n71 256.663
R1789 B.n759 B.n71 256.663
R1790 B.n761 B.n71 256.663
R1791 B.n767 B.n71 256.663
R1792 B.n769 B.n71 256.663
R1793 B.n775 B.n71 256.663
R1794 B.n110 B.n71 256.663
R1795 B.n781 B.n71 256.663
R1796 B.n787 B.n71 256.663
R1797 B.n789 B.n71 256.663
R1798 B.n795 B.n71 256.663
R1799 B.n102 B.n71 256.663
R1800 B.n801 B.n71 256.663
R1801 B.n807 B.n71 256.663
R1802 B.n809 B.n71 256.663
R1803 B.n815 B.n71 256.663
R1804 B.n817 B.n71 256.663
R1805 B.n823 B.n71 256.663
R1806 B.n825 B.n71 256.663
R1807 B.n831 B.n71 256.663
R1808 B.n833 B.n71 256.663
R1809 B.n839 B.n71 256.663
R1810 B.n841 B.n71 256.663
R1811 B.n847 B.n71 256.663
R1812 B.n849 B.n71 256.663
R1813 B.n855 B.n71 256.663
R1814 B.n857 B.n71 256.663
R1815 B.n863 B.n71 256.663
R1816 B.n865 B.n71 256.663
R1817 B.n871 B.n71 256.663
R1818 B.n873 B.n71 256.663
R1819 B.n879 B.n71 256.663
R1820 B.n881 B.n71 256.663
R1821 B.n887 B.n71 256.663
R1822 B.n889 B.n71 256.663
R1823 B.n895 B.n71 256.663
R1824 B.n897 B.n71 256.663
R1825 B.n903 B.n71 256.663
R1826 B.n905 B.n71 256.663
R1827 B.n504 B.n209 256.663
R1828 B.n212 B.n209 256.663
R1829 B.n497 B.n209 256.663
R1830 B.n491 B.n209 256.663
R1831 B.n489 B.n209 256.663
R1832 B.n483 B.n209 256.663
R1833 B.n481 B.n209 256.663
R1834 B.n475 B.n209 256.663
R1835 B.n473 B.n209 256.663
R1836 B.n467 B.n209 256.663
R1837 B.n465 B.n209 256.663
R1838 B.n459 B.n209 256.663
R1839 B.n457 B.n209 256.663
R1840 B.n451 B.n209 256.663
R1841 B.n449 B.n209 256.663
R1842 B.n443 B.n209 256.663
R1843 B.n441 B.n209 256.663
R1844 B.n435 B.n209 256.663
R1845 B.n433 B.n209 256.663
R1846 B.n427 B.n209 256.663
R1847 B.n425 B.n209 256.663
R1848 B.n419 B.n209 256.663
R1849 B.n417 B.n209 256.663
R1850 B.n411 B.n209 256.663
R1851 B.n409 B.n209 256.663
R1852 B.n403 B.n209 256.663
R1853 B.n401 B.n209 256.663
R1854 B.n395 B.n209 256.663
R1855 B.n393 B.n209 256.663
R1856 B.n387 B.n209 256.663
R1857 B.n385 B.n209 256.663
R1858 B.n378 B.n209 256.663
R1859 B.n376 B.n209 256.663
R1860 B.n370 B.n209 256.663
R1861 B.n368 B.n209 256.663
R1862 B.n362 B.n209 256.663
R1863 B.n360 B.n209 256.663
R1864 B.n354 B.n209 256.663
R1865 B.n352 B.n209 256.663
R1866 B.n346 B.n209 256.663
R1867 B.n344 B.n209 256.663
R1868 B.n338 B.n209 256.663
R1869 B.n336 B.n209 256.663
R1870 B.n330 B.n209 256.663
R1871 B.n328 B.n209 256.663
R1872 B.n322 B.n209 256.663
R1873 B.n320 B.n209 256.663
R1874 B.n314 B.n209 256.663
R1875 B.n312 B.n209 256.663
R1876 B.n306 B.n209 256.663
R1877 B.n304 B.n209 256.663
R1878 B.n298 B.n209 256.663
R1879 B.n296 B.n209 256.663
R1880 B.n290 B.n209 256.663
R1881 B.n288 B.n209 256.663
R1882 B.n282 B.n209 256.663
R1883 B.n280 B.n209 256.663
R1884 B.n274 B.n209 256.663
R1885 B.n509 B.n204 163.367
R1886 B.n517 B.n204 163.367
R1887 B.n517 B.n202 163.367
R1888 B.n521 B.n202 163.367
R1889 B.n521 B.n196 163.367
R1890 B.n529 B.n196 163.367
R1891 B.n529 B.n194 163.367
R1892 B.n533 B.n194 163.367
R1893 B.n533 B.n188 163.367
R1894 B.n541 B.n188 163.367
R1895 B.n541 B.n186 163.367
R1896 B.n545 B.n186 163.367
R1897 B.n545 B.n180 163.367
R1898 B.n554 B.n180 163.367
R1899 B.n554 B.n178 163.367
R1900 B.n558 B.n178 163.367
R1901 B.n558 B.n173 163.367
R1902 B.n566 B.n173 163.367
R1903 B.n566 B.n171 163.367
R1904 B.n570 B.n171 163.367
R1905 B.n570 B.n165 163.367
R1906 B.n578 B.n165 163.367
R1907 B.n578 B.n163 163.367
R1908 B.n582 B.n163 163.367
R1909 B.n582 B.n157 163.367
R1910 B.n591 B.n157 163.367
R1911 B.n591 B.n155 163.367
R1912 B.n595 B.n155 163.367
R1913 B.n595 B.n150 163.367
R1914 B.n603 B.n150 163.367
R1915 B.n603 B.n148 163.367
R1916 B.n607 B.n148 163.367
R1917 B.n607 B.n142 163.367
R1918 B.n616 B.n142 163.367
R1919 B.n616 B.n140 163.367
R1920 B.n620 B.n140 163.367
R1921 B.n620 B.n2 163.367
R1922 B.n986 B.n2 163.367
R1923 B.n986 B.n3 163.367
R1924 B.n982 B.n3 163.367
R1925 B.n982 B.n9 163.367
R1926 B.n978 B.n9 163.367
R1927 B.n978 B.n11 163.367
R1928 B.n974 B.n11 163.367
R1929 B.n974 B.n16 163.367
R1930 B.n970 B.n16 163.367
R1931 B.n970 B.n18 163.367
R1932 B.n966 B.n18 163.367
R1933 B.n966 B.n22 163.367
R1934 B.n962 B.n22 163.367
R1935 B.n962 B.n24 163.367
R1936 B.n958 B.n24 163.367
R1937 B.n958 B.n30 163.367
R1938 B.n954 B.n30 163.367
R1939 B.n954 B.n32 163.367
R1940 B.n950 B.n32 163.367
R1941 B.n950 B.n37 163.367
R1942 B.n946 B.n37 163.367
R1943 B.n946 B.n39 163.367
R1944 B.n942 B.n39 163.367
R1945 B.n942 B.n43 163.367
R1946 B.n938 B.n43 163.367
R1947 B.n938 B.n45 163.367
R1948 B.n934 B.n45 163.367
R1949 B.n934 B.n51 163.367
R1950 B.n930 B.n51 163.367
R1951 B.n930 B.n53 163.367
R1952 B.n926 B.n53 163.367
R1953 B.n926 B.n58 163.367
R1954 B.n922 B.n58 163.367
R1955 B.n922 B.n60 163.367
R1956 B.n918 B.n60 163.367
R1957 B.n918 B.n65 163.367
R1958 B.n914 B.n65 163.367
R1959 B.n914 B.n67 163.367
R1960 B.n910 B.n67 163.367
R1961 B.n505 B.n503 163.367
R1962 B.n503 B.n502 163.367
R1963 B.n499 B.n498 163.367
R1964 B.n496 B.n214 163.367
R1965 B.n492 B.n490 163.367
R1966 B.n488 B.n216 163.367
R1967 B.n484 B.n482 163.367
R1968 B.n480 B.n218 163.367
R1969 B.n476 B.n474 163.367
R1970 B.n472 B.n220 163.367
R1971 B.n468 B.n466 163.367
R1972 B.n464 B.n222 163.367
R1973 B.n460 B.n458 163.367
R1974 B.n456 B.n224 163.367
R1975 B.n452 B.n450 163.367
R1976 B.n448 B.n226 163.367
R1977 B.n444 B.n442 163.367
R1978 B.n440 B.n228 163.367
R1979 B.n436 B.n434 163.367
R1980 B.n432 B.n230 163.367
R1981 B.n428 B.n426 163.367
R1982 B.n424 B.n232 163.367
R1983 B.n420 B.n418 163.367
R1984 B.n416 B.n234 163.367
R1985 B.n412 B.n410 163.367
R1986 B.n408 B.n236 163.367
R1987 B.n404 B.n402 163.367
R1988 B.n400 B.n238 163.367
R1989 B.n396 B.n394 163.367
R1990 B.n392 B.n243 163.367
R1991 B.n388 B.n386 163.367
R1992 B.n384 B.n245 163.367
R1993 B.n379 B.n377 163.367
R1994 B.n375 B.n249 163.367
R1995 B.n371 B.n369 163.367
R1996 B.n367 B.n251 163.367
R1997 B.n363 B.n361 163.367
R1998 B.n359 B.n253 163.367
R1999 B.n355 B.n353 163.367
R2000 B.n351 B.n255 163.367
R2001 B.n347 B.n345 163.367
R2002 B.n343 B.n257 163.367
R2003 B.n339 B.n337 163.367
R2004 B.n335 B.n259 163.367
R2005 B.n331 B.n329 163.367
R2006 B.n327 B.n261 163.367
R2007 B.n323 B.n321 163.367
R2008 B.n319 B.n263 163.367
R2009 B.n315 B.n313 163.367
R2010 B.n311 B.n265 163.367
R2011 B.n307 B.n305 163.367
R2012 B.n303 B.n267 163.367
R2013 B.n299 B.n297 163.367
R2014 B.n295 B.n269 163.367
R2015 B.n291 B.n289 163.367
R2016 B.n287 B.n271 163.367
R2017 B.n283 B.n281 163.367
R2018 B.n279 B.n273 163.367
R2019 B.n275 B.n208 163.367
R2020 B.n511 B.n206 163.367
R2021 B.n515 B.n206 163.367
R2022 B.n515 B.n200 163.367
R2023 B.n523 B.n200 163.367
R2024 B.n523 B.n198 163.367
R2025 B.n527 B.n198 163.367
R2026 B.n527 B.n192 163.367
R2027 B.n535 B.n192 163.367
R2028 B.n535 B.n190 163.367
R2029 B.n539 B.n190 163.367
R2030 B.n539 B.n184 163.367
R2031 B.n547 B.n184 163.367
R2032 B.n547 B.n182 163.367
R2033 B.n551 B.n182 163.367
R2034 B.n551 B.n177 163.367
R2035 B.n560 B.n177 163.367
R2036 B.n560 B.n175 163.367
R2037 B.n564 B.n175 163.367
R2038 B.n564 B.n168 163.367
R2039 B.n572 B.n168 163.367
R2040 B.n572 B.n166 163.367
R2041 B.n576 B.n166 163.367
R2042 B.n576 B.n161 163.367
R2043 B.n584 B.n161 163.367
R2044 B.n584 B.n159 163.367
R2045 B.n588 B.n159 163.367
R2046 B.n588 B.n154 163.367
R2047 B.n597 B.n154 163.367
R2048 B.n597 B.n152 163.367
R2049 B.n601 B.n152 163.367
R2050 B.n601 B.n145 163.367
R2051 B.n609 B.n145 163.367
R2052 B.n609 B.n143 163.367
R2053 B.n614 B.n143 163.367
R2054 B.n614 B.n138 163.367
R2055 B.n622 B.n138 163.367
R2056 B.n623 B.n622 163.367
R2057 B.n623 B.n5 163.367
R2058 B.n6 B.n5 163.367
R2059 B.n7 B.n6 163.367
R2060 B.n628 B.n7 163.367
R2061 B.n628 B.n12 163.367
R2062 B.n13 B.n12 163.367
R2063 B.n14 B.n13 163.367
R2064 B.n633 B.n14 163.367
R2065 B.n633 B.n19 163.367
R2066 B.n20 B.n19 163.367
R2067 B.n21 B.n20 163.367
R2068 B.n638 B.n21 163.367
R2069 B.n638 B.n26 163.367
R2070 B.n27 B.n26 163.367
R2071 B.n28 B.n27 163.367
R2072 B.n643 B.n28 163.367
R2073 B.n643 B.n33 163.367
R2074 B.n34 B.n33 163.367
R2075 B.n35 B.n34 163.367
R2076 B.n648 B.n35 163.367
R2077 B.n648 B.n40 163.367
R2078 B.n41 B.n40 163.367
R2079 B.n42 B.n41 163.367
R2080 B.n653 B.n42 163.367
R2081 B.n653 B.n47 163.367
R2082 B.n48 B.n47 163.367
R2083 B.n49 B.n48 163.367
R2084 B.n658 B.n49 163.367
R2085 B.n658 B.n54 163.367
R2086 B.n55 B.n54 163.367
R2087 B.n56 B.n55 163.367
R2088 B.n663 B.n56 163.367
R2089 B.n663 B.n61 163.367
R2090 B.n62 B.n61 163.367
R2091 B.n63 B.n62 163.367
R2092 B.n668 B.n63 163.367
R2093 B.n668 B.n68 163.367
R2094 B.n69 B.n68 163.367
R2095 B.n70 B.n69 163.367
R2096 B.n906 B.n904 163.367
R2097 B.n902 B.n74 163.367
R2098 B.n898 B.n896 163.367
R2099 B.n894 B.n76 163.367
R2100 B.n890 B.n888 163.367
R2101 B.n886 B.n78 163.367
R2102 B.n882 B.n880 163.367
R2103 B.n878 B.n80 163.367
R2104 B.n874 B.n872 163.367
R2105 B.n870 B.n82 163.367
R2106 B.n866 B.n864 163.367
R2107 B.n862 B.n84 163.367
R2108 B.n858 B.n856 163.367
R2109 B.n854 B.n86 163.367
R2110 B.n850 B.n848 163.367
R2111 B.n846 B.n88 163.367
R2112 B.n842 B.n840 163.367
R2113 B.n838 B.n90 163.367
R2114 B.n834 B.n832 163.367
R2115 B.n830 B.n92 163.367
R2116 B.n826 B.n824 163.367
R2117 B.n822 B.n94 163.367
R2118 B.n818 B.n816 163.367
R2119 B.n814 B.n96 163.367
R2120 B.n810 B.n808 163.367
R2121 B.n806 B.n98 163.367
R2122 B.n802 B.n800 163.367
R2123 B.n797 B.n796 163.367
R2124 B.n794 B.n104 163.367
R2125 B.n790 B.n788 163.367
R2126 B.n786 B.n106 163.367
R2127 B.n782 B.n780 163.367
R2128 B.n777 B.n776 163.367
R2129 B.n774 B.n112 163.367
R2130 B.n770 B.n768 163.367
R2131 B.n766 B.n114 163.367
R2132 B.n762 B.n760 163.367
R2133 B.n758 B.n116 163.367
R2134 B.n754 B.n752 163.367
R2135 B.n750 B.n118 163.367
R2136 B.n746 B.n744 163.367
R2137 B.n742 B.n120 163.367
R2138 B.n738 B.n736 163.367
R2139 B.n734 B.n122 163.367
R2140 B.n730 B.n728 163.367
R2141 B.n726 B.n124 163.367
R2142 B.n722 B.n720 163.367
R2143 B.n718 B.n126 163.367
R2144 B.n714 B.n712 163.367
R2145 B.n710 B.n128 163.367
R2146 B.n706 B.n704 163.367
R2147 B.n702 B.n130 163.367
R2148 B.n698 B.n696 163.367
R2149 B.n694 B.n132 163.367
R2150 B.n690 B.n688 163.367
R2151 B.n686 B.n134 163.367
R2152 B.n682 B.n680 163.367
R2153 B.n678 B.n136 163.367
R2154 B.n510 B.n209 72.224
R2155 B.n911 B.n71 72.224
R2156 B.n504 B.n210 71.676
R2157 B.n502 B.n212 71.676
R2158 B.n498 B.n497 71.676
R2159 B.n491 B.n214 71.676
R2160 B.n490 B.n489 71.676
R2161 B.n483 B.n216 71.676
R2162 B.n482 B.n481 71.676
R2163 B.n475 B.n218 71.676
R2164 B.n474 B.n473 71.676
R2165 B.n467 B.n220 71.676
R2166 B.n466 B.n465 71.676
R2167 B.n459 B.n222 71.676
R2168 B.n458 B.n457 71.676
R2169 B.n451 B.n224 71.676
R2170 B.n450 B.n449 71.676
R2171 B.n443 B.n226 71.676
R2172 B.n442 B.n441 71.676
R2173 B.n435 B.n228 71.676
R2174 B.n434 B.n433 71.676
R2175 B.n427 B.n230 71.676
R2176 B.n426 B.n425 71.676
R2177 B.n419 B.n232 71.676
R2178 B.n418 B.n417 71.676
R2179 B.n411 B.n234 71.676
R2180 B.n410 B.n409 71.676
R2181 B.n403 B.n236 71.676
R2182 B.n402 B.n401 71.676
R2183 B.n395 B.n238 71.676
R2184 B.n394 B.n393 71.676
R2185 B.n387 B.n243 71.676
R2186 B.n386 B.n385 71.676
R2187 B.n378 B.n245 71.676
R2188 B.n377 B.n376 71.676
R2189 B.n370 B.n249 71.676
R2190 B.n369 B.n368 71.676
R2191 B.n362 B.n251 71.676
R2192 B.n361 B.n360 71.676
R2193 B.n354 B.n253 71.676
R2194 B.n353 B.n352 71.676
R2195 B.n346 B.n255 71.676
R2196 B.n345 B.n344 71.676
R2197 B.n338 B.n257 71.676
R2198 B.n337 B.n336 71.676
R2199 B.n330 B.n259 71.676
R2200 B.n329 B.n328 71.676
R2201 B.n322 B.n261 71.676
R2202 B.n321 B.n320 71.676
R2203 B.n314 B.n263 71.676
R2204 B.n313 B.n312 71.676
R2205 B.n306 B.n265 71.676
R2206 B.n305 B.n304 71.676
R2207 B.n298 B.n267 71.676
R2208 B.n297 B.n296 71.676
R2209 B.n290 B.n269 71.676
R2210 B.n289 B.n288 71.676
R2211 B.n282 B.n271 71.676
R2212 B.n281 B.n280 71.676
R2213 B.n274 B.n273 71.676
R2214 B.n905 B.n72 71.676
R2215 B.n904 B.n903 71.676
R2216 B.n897 B.n74 71.676
R2217 B.n896 B.n895 71.676
R2218 B.n889 B.n76 71.676
R2219 B.n888 B.n887 71.676
R2220 B.n881 B.n78 71.676
R2221 B.n880 B.n879 71.676
R2222 B.n873 B.n80 71.676
R2223 B.n872 B.n871 71.676
R2224 B.n865 B.n82 71.676
R2225 B.n864 B.n863 71.676
R2226 B.n857 B.n84 71.676
R2227 B.n856 B.n855 71.676
R2228 B.n849 B.n86 71.676
R2229 B.n848 B.n847 71.676
R2230 B.n841 B.n88 71.676
R2231 B.n840 B.n839 71.676
R2232 B.n833 B.n90 71.676
R2233 B.n832 B.n831 71.676
R2234 B.n825 B.n92 71.676
R2235 B.n824 B.n823 71.676
R2236 B.n817 B.n94 71.676
R2237 B.n816 B.n815 71.676
R2238 B.n809 B.n96 71.676
R2239 B.n808 B.n807 71.676
R2240 B.n801 B.n98 71.676
R2241 B.n800 B.n102 71.676
R2242 B.n796 B.n795 71.676
R2243 B.n789 B.n104 71.676
R2244 B.n788 B.n787 71.676
R2245 B.n781 B.n106 71.676
R2246 B.n780 B.n110 71.676
R2247 B.n776 B.n775 71.676
R2248 B.n769 B.n112 71.676
R2249 B.n768 B.n767 71.676
R2250 B.n761 B.n114 71.676
R2251 B.n760 B.n759 71.676
R2252 B.n753 B.n116 71.676
R2253 B.n752 B.n751 71.676
R2254 B.n745 B.n118 71.676
R2255 B.n744 B.n743 71.676
R2256 B.n737 B.n120 71.676
R2257 B.n736 B.n735 71.676
R2258 B.n729 B.n122 71.676
R2259 B.n728 B.n727 71.676
R2260 B.n721 B.n124 71.676
R2261 B.n720 B.n719 71.676
R2262 B.n713 B.n126 71.676
R2263 B.n712 B.n711 71.676
R2264 B.n705 B.n128 71.676
R2265 B.n704 B.n703 71.676
R2266 B.n697 B.n130 71.676
R2267 B.n696 B.n695 71.676
R2268 B.n689 B.n132 71.676
R2269 B.n688 B.n687 71.676
R2270 B.n681 B.n134 71.676
R2271 B.n680 B.n679 71.676
R2272 B.n673 B.n136 71.676
R2273 B.n674 B.n673 71.676
R2274 B.n679 B.n678 71.676
R2275 B.n682 B.n681 71.676
R2276 B.n687 B.n686 71.676
R2277 B.n690 B.n689 71.676
R2278 B.n695 B.n694 71.676
R2279 B.n698 B.n697 71.676
R2280 B.n703 B.n702 71.676
R2281 B.n706 B.n705 71.676
R2282 B.n711 B.n710 71.676
R2283 B.n714 B.n713 71.676
R2284 B.n719 B.n718 71.676
R2285 B.n722 B.n721 71.676
R2286 B.n727 B.n726 71.676
R2287 B.n730 B.n729 71.676
R2288 B.n735 B.n734 71.676
R2289 B.n738 B.n737 71.676
R2290 B.n743 B.n742 71.676
R2291 B.n746 B.n745 71.676
R2292 B.n751 B.n750 71.676
R2293 B.n754 B.n753 71.676
R2294 B.n759 B.n758 71.676
R2295 B.n762 B.n761 71.676
R2296 B.n767 B.n766 71.676
R2297 B.n770 B.n769 71.676
R2298 B.n775 B.n774 71.676
R2299 B.n777 B.n110 71.676
R2300 B.n782 B.n781 71.676
R2301 B.n787 B.n786 71.676
R2302 B.n790 B.n789 71.676
R2303 B.n795 B.n794 71.676
R2304 B.n797 B.n102 71.676
R2305 B.n802 B.n801 71.676
R2306 B.n807 B.n806 71.676
R2307 B.n810 B.n809 71.676
R2308 B.n815 B.n814 71.676
R2309 B.n818 B.n817 71.676
R2310 B.n823 B.n822 71.676
R2311 B.n826 B.n825 71.676
R2312 B.n831 B.n830 71.676
R2313 B.n834 B.n833 71.676
R2314 B.n839 B.n838 71.676
R2315 B.n842 B.n841 71.676
R2316 B.n847 B.n846 71.676
R2317 B.n850 B.n849 71.676
R2318 B.n855 B.n854 71.676
R2319 B.n858 B.n857 71.676
R2320 B.n863 B.n862 71.676
R2321 B.n866 B.n865 71.676
R2322 B.n871 B.n870 71.676
R2323 B.n874 B.n873 71.676
R2324 B.n879 B.n878 71.676
R2325 B.n882 B.n881 71.676
R2326 B.n887 B.n886 71.676
R2327 B.n890 B.n889 71.676
R2328 B.n895 B.n894 71.676
R2329 B.n898 B.n897 71.676
R2330 B.n903 B.n902 71.676
R2331 B.n906 B.n905 71.676
R2332 B.n505 B.n504 71.676
R2333 B.n499 B.n212 71.676
R2334 B.n497 B.n496 71.676
R2335 B.n492 B.n491 71.676
R2336 B.n489 B.n488 71.676
R2337 B.n484 B.n483 71.676
R2338 B.n481 B.n480 71.676
R2339 B.n476 B.n475 71.676
R2340 B.n473 B.n472 71.676
R2341 B.n468 B.n467 71.676
R2342 B.n465 B.n464 71.676
R2343 B.n460 B.n459 71.676
R2344 B.n457 B.n456 71.676
R2345 B.n452 B.n451 71.676
R2346 B.n449 B.n448 71.676
R2347 B.n444 B.n443 71.676
R2348 B.n441 B.n440 71.676
R2349 B.n436 B.n435 71.676
R2350 B.n433 B.n432 71.676
R2351 B.n428 B.n427 71.676
R2352 B.n425 B.n424 71.676
R2353 B.n420 B.n419 71.676
R2354 B.n417 B.n416 71.676
R2355 B.n412 B.n411 71.676
R2356 B.n409 B.n408 71.676
R2357 B.n404 B.n403 71.676
R2358 B.n401 B.n400 71.676
R2359 B.n396 B.n395 71.676
R2360 B.n393 B.n392 71.676
R2361 B.n388 B.n387 71.676
R2362 B.n385 B.n384 71.676
R2363 B.n379 B.n378 71.676
R2364 B.n376 B.n375 71.676
R2365 B.n371 B.n370 71.676
R2366 B.n368 B.n367 71.676
R2367 B.n363 B.n362 71.676
R2368 B.n360 B.n359 71.676
R2369 B.n355 B.n354 71.676
R2370 B.n352 B.n351 71.676
R2371 B.n347 B.n346 71.676
R2372 B.n344 B.n343 71.676
R2373 B.n339 B.n338 71.676
R2374 B.n336 B.n335 71.676
R2375 B.n331 B.n330 71.676
R2376 B.n328 B.n327 71.676
R2377 B.n323 B.n322 71.676
R2378 B.n320 B.n319 71.676
R2379 B.n315 B.n314 71.676
R2380 B.n312 B.n311 71.676
R2381 B.n307 B.n306 71.676
R2382 B.n304 B.n303 71.676
R2383 B.n299 B.n298 71.676
R2384 B.n296 B.n295 71.676
R2385 B.n291 B.n290 71.676
R2386 B.n288 B.n287 71.676
R2387 B.n283 B.n282 71.676
R2388 B.n280 B.n279 71.676
R2389 B.n275 B.n274 71.676
R2390 B.n381 B.n247 59.5399
R2391 B.n241 B.n240 59.5399
R2392 B.n101 B.n100 59.5399
R2393 B.n109 B.n108 59.5399
R2394 B.n247 B.n246 39.7581
R2395 B.n240 B.n239 39.7581
R2396 B.n100 B.n99 39.7581
R2397 B.n108 B.n107 39.7581
R2398 B.n510 B.n205 34.8317
R2399 B.n516 B.n205 34.8317
R2400 B.n516 B.n201 34.8317
R2401 B.n522 B.n201 34.8317
R2402 B.n522 B.n197 34.8317
R2403 B.n528 B.n197 34.8317
R2404 B.n534 B.n193 34.8317
R2405 B.n534 B.n189 34.8317
R2406 B.n540 B.n189 34.8317
R2407 B.n540 B.n185 34.8317
R2408 B.n546 B.n185 34.8317
R2409 B.n546 B.n181 34.8317
R2410 B.n553 B.n181 34.8317
R2411 B.n553 B.n552 34.8317
R2412 B.n559 B.n174 34.8317
R2413 B.n565 B.n174 34.8317
R2414 B.n565 B.n169 34.8317
R2415 B.n571 B.n169 34.8317
R2416 B.n571 B.n170 34.8317
R2417 B.n577 B.n162 34.8317
R2418 B.n583 B.n162 34.8317
R2419 B.n583 B.n158 34.8317
R2420 B.n590 B.n158 34.8317
R2421 B.n590 B.n589 34.8317
R2422 B.n596 B.n151 34.8317
R2423 B.n602 B.n151 34.8317
R2424 B.n602 B.n146 34.8317
R2425 B.n608 B.n146 34.8317
R2426 B.n608 B.n147 34.8317
R2427 B.n615 B.n139 34.8317
R2428 B.n621 B.n139 34.8317
R2429 B.n621 B.n4 34.8317
R2430 B.n985 B.n4 34.8317
R2431 B.n985 B.n984 34.8317
R2432 B.n984 B.n983 34.8317
R2433 B.n983 B.n8 34.8317
R2434 B.n977 B.n8 34.8317
R2435 B.n976 B.n975 34.8317
R2436 B.n975 B.n15 34.8317
R2437 B.n969 B.n15 34.8317
R2438 B.n969 B.n968 34.8317
R2439 B.n968 B.n967 34.8317
R2440 B.n961 B.n25 34.8317
R2441 B.n961 B.n960 34.8317
R2442 B.n960 B.n959 34.8317
R2443 B.n959 B.n29 34.8317
R2444 B.n953 B.n29 34.8317
R2445 B.n952 B.n951 34.8317
R2446 B.n951 B.n36 34.8317
R2447 B.n945 B.n36 34.8317
R2448 B.n945 B.n944 34.8317
R2449 B.n944 B.n943 34.8317
R2450 B.n937 B.n46 34.8317
R2451 B.n937 B.n936 34.8317
R2452 B.n936 B.n935 34.8317
R2453 B.n935 B.n50 34.8317
R2454 B.n929 B.n50 34.8317
R2455 B.n929 B.n928 34.8317
R2456 B.n928 B.n927 34.8317
R2457 B.n927 B.n57 34.8317
R2458 B.n921 B.n920 34.8317
R2459 B.n920 B.n919 34.8317
R2460 B.n919 B.n64 34.8317
R2461 B.n913 B.n64 34.8317
R2462 B.n913 B.n912 34.8317
R2463 B.n912 B.n911 34.8317
R2464 B.t16 B.n193 32.7828
R2465 B.t9 B.n57 32.7828
R2466 B.n909 B.n908 32.6249
R2467 B.n675 B.n672 32.6249
R2468 B.n512 B.n207 32.6249
R2469 B.n508 B.n507 32.6249
R2470 B.n559 B.t6 24.5872
R2471 B.n943 B.t5 24.5872
R2472 B.n577 B.t0 23.5628
R2473 B.n953 B.t4 23.5628
R2474 B.n596 B.t1 22.5383
R2475 B.n967 B.t2 22.5383
R2476 B.n615 B.t7 21.5139
R2477 B.n977 B.t3 21.5139
R2478 B B.n987 18.0485
R2479 B.n147 B.t7 13.3183
R2480 B.t3 B.n976 13.3183
R2481 B.n589 B.t1 12.2939
R2482 B.n25 B.t2 12.2939
R2483 B.n170 B.t0 11.2694
R2484 B.t4 B.n952 11.2694
R2485 B.n908 B.n907 10.6151
R2486 B.n907 B.n73 10.6151
R2487 B.n901 B.n73 10.6151
R2488 B.n901 B.n900 10.6151
R2489 B.n900 B.n899 10.6151
R2490 B.n899 B.n75 10.6151
R2491 B.n893 B.n75 10.6151
R2492 B.n893 B.n892 10.6151
R2493 B.n892 B.n891 10.6151
R2494 B.n891 B.n77 10.6151
R2495 B.n885 B.n77 10.6151
R2496 B.n885 B.n884 10.6151
R2497 B.n884 B.n883 10.6151
R2498 B.n883 B.n79 10.6151
R2499 B.n877 B.n79 10.6151
R2500 B.n877 B.n876 10.6151
R2501 B.n876 B.n875 10.6151
R2502 B.n875 B.n81 10.6151
R2503 B.n869 B.n81 10.6151
R2504 B.n869 B.n868 10.6151
R2505 B.n868 B.n867 10.6151
R2506 B.n867 B.n83 10.6151
R2507 B.n861 B.n83 10.6151
R2508 B.n861 B.n860 10.6151
R2509 B.n860 B.n859 10.6151
R2510 B.n859 B.n85 10.6151
R2511 B.n853 B.n85 10.6151
R2512 B.n853 B.n852 10.6151
R2513 B.n852 B.n851 10.6151
R2514 B.n851 B.n87 10.6151
R2515 B.n845 B.n87 10.6151
R2516 B.n845 B.n844 10.6151
R2517 B.n844 B.n843 10.6151
R2518 B.n843 B.n89 10.6151
R2519 B.n837 B.n89 10.6151
R2520 B.n837 B.n836 10.6151
R2521 B.n836 B.n835 10.6151
R2522 B.n835 B.n91 10.6151
R2523 B.n829 B.n91 10.6151
R2524 B.n829 B.n828 10.6151
R2525 B.n828 B.n827 10.6151
R2526 B.n827 B.n93 10.6151
R2527 B.n821 B.n93 10.6151
R2528 B.n821 B.n820 10.6151
R2529 B.n820 B.n819 10.6151
R2530 B.n819 B.n95 10.6151
R2531 B.n813 B.n95 10.6151
R2532 B.n813 B.n812 10.6151
R2533 B.n812 B.n811 10.6151
R2534 B.n811 B.n97 10.6151
R2535 B.n805 B.n97 10.6151
R2536 B.n805 B.n804 10.6151
R2537 B.n804 B.n803 10.6151
R2538 B.n799 B.n798 10.6151
R2539 B.n798 B.n103 10.6151
R2540 B.n793 B.n103 10.6151
R2541 B.n793 B.n792 10.6151
R2542 B.n792 B.n791 10.6151
R2543 B.n791 B.n105 10.6151
R2544 B.n785 B.n105 10.6151
R2545 B.n785 B.n784 10.6151
R2546 B.n784 B.n783 10.6151
R2547 B.n779 B.n778 10.6151
R2548 B.n778 B.n111 10.6151
R2549 B.n773 B.n111 10.6151
R2550 B.n773 B.n772 10.6151
R2551 B.n772 B.n771 10.6151
R2552 B.n771 B.n113 10.6151
R2553 B.n765 B.n113 10.6151
R2554 B.n765 B.n764 10.6151
R2555 B.n764 B.n763 10.6151
R2556 B.n763 B.n115 10.6151
R2557 B.n757 B.n115 10.6151
R2558 B.n757 B.n756 10.6151
R2559 B.n756 B.n755 10.6151
R2560 B.n755 B.n117 10.6151
R2561 B.n749 B.n117 10.6151
R2562 B.n749 B.n748 10.6151
R2563 B.n748 B.n747 10.6151
R2564 B.n747 B.n119 10.6151
R2565 B.n741 B.n119 10.6151
R2566 B.n741 B.n740 10.6151
R2567 B.n740 B.n739 10.6151
R2568 B.n739 B.n121 10.6151
R2569 B.n733 B.n121 10.6151
R2570 B.n733 B.n732 10.6151
R2571 B.n732 B.n731 10.6151
R2572 B.n731 B.n123 10.6151
R2573 B.n725 B.n123 10.6151
R2574 B.n725 B.n724 10.6151
R2575 B.n724 B.n723 10.6151
R2576 B.n723 B.n125 10.6151
R2577 B.n717 B.n125 10.6151
R2578 B.n717 B.n716 10.6151
R2579 B.n716 B.n715 10.6151
R2580 B.n715 B.n127 10.6151
R2581 B.n709 B.n127 10.6151
R2582 B.n709 B.n708 10.6151
R2583 B.n708 B.n707 10.6151
R2584 B.n707 B.n129 10.6151
R2585 B.n701 B.n129 10.6151
R2586 B.n701 B.n700 10.6151
R2587 B.n700 B.n699 10.6151
R2588 B.n699 B.n131 10.6151
R2589 B.n693 B.n131 10.6151
R2590 B.n693 B.n692 10.6151
R2591 B.n692 B.n691 10.6151
R2592 B.n691 B.n133 10.6151
R2593 B.n685 B.n133 10.6151
R2594 B.n685 B.n684 10.6151
R2595 B.n684 B.n683 10.6151
R2596 B.n683 B.n135 10.6151
R2597 B.n677 B.n135 10.6151
R2598 B.n677 B.n676 10.6151
R2599 B.n676 B.n675 10.6151
R2600 B.n513 B.n512 10.6151
R2601 B.n514 B.n513 10.6151
R2602 B.n514 B.n199 10.6151
R2603 B.n524 B.n199 10.6151
R2604 B.n525 B.n524 10.6151
R2605 B.n526 B.n525 10.6151
R2606 B.n526 B.n191 10.6151
R2607 B.n536 B.n191 10.6151
R2608 B.n537 B.n536 10.6151
R2609 B.n538 B.n537 10.6151
R2610 B.n538 B.n183 10.6151
R2611 B.n548 B.n183 10.6151
R2612 B.n549 B.n548 10.6151
R2613 B.n550 B.n549 10.6151
R2614 B.n550 B.n176 10.6151
R2615 B.n561 B.n176 10.6151
R2616 B.n562 B.n561 10.6151
R2617 B.n563 B.n562 10.6151
R2618 B.n563 B.n167 10.6151
R2619 B.n573 B.n167 10.6151
R2620 B.n574 B.n573 10.6151
R2621 B.n575 B.n574 10.6151
R2622 B.n575 B.n160 10.6151
R2623 B.n585 B.n160 10.6151
R2624 B.n586 B.n585 10.6151
R2625 B.n587 B.n586 10.6151
R2626 B.n587 B.n153 10.6151
R2627 B.n598 B.n153 10.6151
R2628 B.n599 B.n598 10.6151
R2629 B.n600 B.n599 10.6151
R2630 B.n600 B.n144 10.6151
R2631 B.n610 B.n144 10.6151
R2632 B.n611 B.n610 10.6151
R2633 B.n613 B.n611 10.6151
R2634 B.n613 B.n612 10.6151
R2635 B.n612 B.n137 10.6151
R2636 B.n624 B.n137 10.6151
R2637 B.n625 B.n624 10.6151
R2638 B.n626 B.n625 10.6151
R2639 B.n627 B.n626 10.6151
R2640 B.n629 B.n627 10.6151
R2641 B.n630 B.n629 10.6151
R2642 B.n631 B.n630 10.6151
R2643 B.n632 B.n631 10.6151
R2644 B.n634 B.n632 10.6151
R2645 B.n635 B.n634 10.6151
R2646 B.n636 B.n635 10.6151
R2647 B.n637 B.n636 10.6151
R2648 B.n639 B.n637 10.6151
R2649 B.n640 B.n639 10.6151
R2650 B.n641 B.n640 10.6151
R2651 B.n642 B.n641 10.6151
R2652 B.n644 B.n642 10.6151
R2653 B.n645 B.n644 10.6151
R2654 B.n646 B.n645 10.6151
R2655 B.n647 B.n646 10.6151
R2656 B.n649 B.n647 10.6151
R2657 B.n650 B.n649 10.6151
R2658 B.n651 B.n650 10.6151
R2659 B.n652 B.n651 10.6151
R2660 B.n654 B.n652 10.6151
R2661 B.n655 B.n654 10.6151
R2662 B.n656 B.n655 10.6151
R2663 B.n657 B.n656 10.6151
R2664 B.n659 B.n657 10.6151
R2665 B.n660 B.n659 10.6151
R2666 B.n661 B.n660 10.6151
R2667 B.n662 B.n661 10.6151
R2668 B.n664 B.n662 10.6151
R2669 B.n665 B.n664 10.6151
R2670 B.n666 B.n665 10.6151
R2671 B.n667 B.n666 10.6151
R2672 B.n669 B.n667 10.6151
R2673 B.n670 B.n669 10.6151
R2674 B.n671 B.n670 10.6151
R2675 B.n672 B.n671 10.6151
R2676 B.n507 B.n506 10.6151
R2677 B.n506 B.n211 10.6151
R2678 B.n501 B.n211 10.6151
R2679 B.n501 B.n500 10.6151
R2680 B.n500 B.n213 10.6151
R2681 B.n495 B.n213 10.6151
R2682 B.n495 B.n494 10.6151
R2683 B.n494 B.n493 10.6151
R2684 B.n493 B.n215 10.6151
R2685 B.n487 B.n215 10.6151
R2686 B.n487 B.n486 10.6151
R2687 B.n486 B.n485 10.6151
R2688 B.n485 B.n217 10.6151
R2689 B.n479 B.n217 10.6151
R2690 B.n479 B.n478 10.6151
R2691 B.n478 B.n477 10.6151
R2692 B.n477 B.n219 10.6151
R2693 B.n471 B.n219 10.6151
R2694 B.n471 B.n470 10.6151
R2695 B.n470 B.n469 10.6151
R2696 B.n469 B.n221 10.6151
R2697 B.n463 B.n221 10.6151
R2698 B.n463 B.n462 10.6151
R2699 B.n462 B.n461 10.6151
R2700 B.n461 B.n223 10.6151
R2701 B.n455 B.n223 10.6151
R2702 B.n455 B.n454 10.6151
R2703 B.n454 B.n453 10.6151
R2704 B.n453 B.n225 10.6151
R2705 B.n447 B.n225 10.6151
R2706 B.n447 B.n446 10.6151
R2707 B.n446 B.n445 10.6151
R2708 B.n445 B.n227 10.6151
R2709 B.n439 B.n227 10.6151
R2710 B.n439 B.n438 10.6151
R2711 B.n438 B.n437 10.6151
R2712 B.n437 B.n229 10.6151
R2713 B.n431 B.n229 10.6151
R2714 B.n431 B.n430 10.6151
R2715 B.n430 B.n429 10.6151
R2716 B.n429 B.n231 10.6151
R2717 B.n423 B.n231 10.6151
R2718 B.n423 B.n422 10.6151
R2719 B.n422 B.n421 10.6151
R2720 B.n421 B.n233 10.6151
R2721 B.n415 B.n233 10.6151
R2722 B.n415 B.n414 10.6151
R2723 B.n414 B.n413 10.6151
R2724 B.n413 B.n235 10.6151
R2725 B.n407 B.n235 10.6151
R2726 B.n407 B.n406 10.6151
R2727 B.n406 B.n405 10.6151
R2728 B.n405 B.n237 10.6151
R2729 B.n399 B.n398 10.6151
R2730 B.n398 B.n397 10.6151
R2731 B.n397 B.n242 10.6151
R2732 B.n391 B.n242 10.6151
R2733 B.n391 B.n390 10.6151
R2734 B.n390 B.n389 10.6151
R2735 B.n389 B.n244 10.6151
R2736 B.n383 B.n244 10.6151
R2737 B.n383 B.n382 10.6151
R2738 B.n380 B.n248 10.6151
R2739 B.n374 B.n248 10.6151
R2740 B.n374 B.n373 10.6151
R2741 B.n373 B.n372 10.6151
R2742 B.n372 B.n250 10.6151
R2743 B.n366 B.n250 10.6151
R2744 B.n366 B.n365 10.6151
R2745 B.n365 B.n364 10.6151
R2746 B.n364 B.n252 10.6151
R2747 B.n358 B.n252 10.6151
R2748 B.n358 B.n357 10.6151
R2749 B.n357 B.n356 10.6151
R2750 B.n356 B.n254 10.6151
R2751 B.n350 B.n254 10.6151
R2752 B.n350 B.n349 10.6151
R2753 B.n349 B.n348 10.6151
R2754 B.n348 B.n256 10.6151
R2755 B.n342 B.n256 10.6151
R2756 B.n342 B.n341 10.6151
R2757 B.n341 B.n340 10.6151
R2758 B.n340 B.n258 10.6151
R2759 B.n334 B.n258 10.6151
R2760 B.n334 B.n333 10.6151
R2761 B.n333 B.n332 10.6151
R2762 B.n332 B.n260 10.6151
R2763 B.n326 B.n260 10.6151
R2764 B.n326 B.n325 10.6151
R2765 B.n325 B.n324 10.6151
R2766 B.n324 B.n262 10.6151
R2767 B.n318 B.n262 10.6151
R2768 B.n318 B.n317 10.6151
R2769 B.n317 B.n316 10.6151
R2770 B.n316 B.n264 10.6151
R2771 B.n310 B.n264 10.6151
R2772 B.n310 B.n309 10.6151
R2773 B.n309 B.n308 10.6151
R2774 B.n308 B.n266 10.6151
R2775 B.n302 B.n266 10.6151
R2776 B.n302 B.n301 10.6151
R2777 B.n301 B.n300 10.6151
R2778 B.n300 B.n268 10.6151
R2779 B.n294 B.n268 10.6151
R2780 B.n294 B.n293 10.6151
R2781 B.n293 B.n292 10.6151
R2782 B.n292 B.n270 10.6151
R2783 B.n286 B.n270 10.6151
R2784 B.n286 B.n285 10.6151
R2785 B.n285 B.n284 10.6151
R2786 B.n284 B.n272 10.6151
R2787 B.n278 B.n272 10.6151
R2788 B.n278 B.n277 10.6151
R2789 B.n277 B.n276 10.6151
R2790 B.n276 B.n207 10.6151
R2791 B.n508 B.n203 10.6151
R2792 B.n518 B.n203 10.6151
R2793 B.n519 B.n518 10.6151
R2794 B.n520 B.n519 10.6151
R2795 B.n520 B.n195 10.6151
R2796 B.n530 B.n195 10.6151
R2797 B.n531 B.n530 10.6151
R2798 B.n532 B.n531 10.6151
R2799 B.n532 B.n187 10.6151
R2800 B.n542 B.n187 10.6151
R2801 B.n543 B.n542 10.6151
R2802 B.n544 B.n543 10.6151
R2803 B.n544 B.n179 10.6151
R2804 B.n555 B.n179 10.6151
R2805 B.n556 B.n555 10.6151
R2806 B.n557 B.n556 10.6151
R2807 B.n557 B.n172 10.6151
R2808 B.n567 B.n172 10.6151
R2809 B.n568 B.n567 10.6151
R2810 B.n569 B.n568 10.6151
R2811 B.n569 B.n164 10.6151
R2812 B.n579 B.n164 10.6151
R2813 B.n580 B.n579 10.6151
R2814 B.n581 B.n580 10.6151
R2815 B.n581 B.n156 10.6151
R2816 B.n592 B.n156 10.6151
R2817 B.n593 B.n592 10.6151
R2818 B.n594 B.n593 10.6151
R2819 B.n594 B.n149 10.6151
R2820 B.n604 B.n149 10.6151
R2821 B.n605 B.n604 10.6151
R2822 B.n606 B.n605 10.6151
R2823 B.n606 B.n141 10.6151
R2824 B.n617 B.n141 10.6151
R2825 B.n618 B.n617 10.6151
R2826 B.n619 B.n618 10.6151
R2827 B.n619 B.n0 10.6151
R2828 B.n981 B.n1 10.6151
R2829 B.n981 B.n980 10.6151
R2830 B.n980 B.n979 10.6151
R2831 B.n979 B.n10 10.6151
R2832 B.n973 B.n10 10.6151
R2833 B.n973 B.n972 10.6151
R2834 B.n972 B.n971 10.6151
R2835 B.n971 B.n17 10.6151
R2836 B.n965 B.n17 10.6151
R2837 B.n965 B.n964 10.6151
R2838 B.n964 B.n963 10.6151
R2839 B.n963 B.n23 10.6151
R2840 B.n957 B.n23 10.6151
R2841 B.n957 B.n956 10.6151
R2842 B.n956 B.n955 10.6151
R2843 B.n955 B.n31 10.6151
R2844 B.n949 B.n31 10.6151
R2845 B.n949 B.n948 10.6151
R2846 B.n948 B.n947 10.6151
R2847 B.n947 B.n38 10.6151
R2848 B.n941 B.n38 10.6151
R2849 B.n941 B.n940 10.6151
R2850 B.n940 B.n939 10.6151
R2851 B.n939 B.n44 10.6151
R2852 B.n933 B.n44 10.6151
R2853 B.n933 B.n932 10.6151
R2854 B.n932 B.n931 10.6151
R2855 B.n931 B.n52 10.6151
R2856 B.n925 B.n52 10.6151
R2857 B.n925 B.n924 10.6151
R2858 B.n924 B.n923 10.6151
R2859 B.n923 B.n59 10.6151
R2860 B.n917 B.n59 10.6151
R2861 B.n917 B.n916 10.6151
R2862 B.n916 B.n915 10.6151
R2863 B.n915 B.n66 10.6151
R2864 B.n909 B.n66 10.6151
R2865 B.n552 B.t6 10.245
R2866 B.n46 B.t5 10.245
R2867 B.n803 B.n101 9.36635
R2868 B.n779 B.n109 9.36635
R2869 B.n241 B.n237 9.36635
R2870 B.n381 B.n380 9.36635
R2871 B.n987 B.n0 2.81026
R2872 B.n987 B.n1 2.81026
R2873 B.n528 B.t16 2.04939
R2874 B.n921 B.t9 2.04939
R2875 B.n799 B.n101 1.24928
R2876 B.n783 B.n109 1.24928
R2877 B.n399 B.n241 1.24928
R2878 B.n382 B.n381 1.24928
R2879 VN.n5 VN.t6 256.594
R2880 VN.n28 VN.t4 256.594
R2881 VN.n6 VN.t1 226.988
R2882 VN.n14 VN.t7 226.988
R2883 VN.n21 VN.t2 226.988
R2884 VN.n29 VN.t0 226.988
R2885 VN.n37 VN.t5 226.988
R2886 VN.n44 VN.t3 226.988
R2887 VN.n22 VN.n21 182.203
R2888 VN.n45 VN.n44 182.203
R2889 VN.n43 VN.n23 161.3
R2890 VN.n42 VN.n41 161.3
R2891 VN.n40 VN.n24 161.3
R2892 VN.n39 VN.n38 161.3
R2893 VN.n36 VN.n25 161.3
R2894 VN.n35 VN.n34 161.3
R2895 VN.n33 VN.n26 161.3
R2896 VN.n32 VN.n31 161.3
R2897 VN.n30 VN.n27 161.3
R2898 VN.n20 VN.n0 161.3
R2899 VN.n19 VN.n18 161.3
R2900 VN.n17 VN.n1 161.3
R2901 VN.n16 VN.n15 161.3
R2902 VN.n13 VN.n2 161.3
R2903 VN.n12 VN.n11 161.3
R2904 VN.n10 VN.n3 161.3
R2905 VN.n9 VN.n8 161.3
R2906 VN.n7 VN.n4 161.3
R2907 VN.n6 VN.n5 67.3815
R2908 VN.n29 VN.n28 67.3815
R2909 VN VN.n45 50.2221
R2910 VN.n19 VN.n1 45.4209
R2911 VN.n42 VN.n24 45.4209
R2912 VN.n8 VN.n3 40.577
R2913 VN.n12 VN.n3 40.577
R2914 VN.n31 VN.n26 40.577
R2915 VN.n35 VN.n26 40.577
R2916 VN.n15 VN.n1 35.7332
R2917 VN.n38 VN.n24 35.7332
R2918 VN.n8 VN.n7 24.5923
R2919 VN.n13 VN.n12 24.5923
R2920 VN.n20 VN.n19 24.5923
R2921 VN.n31 VN.n30 24.5923
R2922 VN.n36 VN.n35 24.5923
R2923 VN.n43 VN.n42 24.5923
R2924 VN.n15 VN.n14 23.3627
R2925 VN.n38 VN.n37 23.3627
R2926 VN.n28 VN.n27 18.5926
R2927 VN.n5 VN.n4 18.5926
R2928 VN.n21 VN.n20 3.68928
R2929 VN.n44 VN.n43 3.68928
R2930 VN.n7 VN.n6 1.23009
R2931 VN.n14 VN.n13 1.23009
R2932 VN.n30 VN.n29 1.23009
R2933 VN.n37 VN.n36 1.23009
R2934 VN.n45 VN.n23 0.189894
R2935 VN.n41 VN.n23 0.189894
R2936 VN.n41 VN.n40 0.189894
R2937 VN.n40 VN.n39 0.189894
R2938 VN.n39 VN.n25 0.189894
R2939 VN.n34 VN.n25 0.189894
R2940 VN.n34 VN.n33 0.189894
R2941 VN.n33 VN.n32 0.189894
R2942 VN.n32 VN.n27 0.189894
R2943 VN.n9 VN.n4 0.189894
R2944 VN.n10 VN.n9 0.189894
R2945 VN.n11 VN.n10 0.189894
R2946 VN.n11 VN.n2 0.189894
R2947 VN.n16 VN.n2 0.189894
R2948 VN.n17 VN.n16 0.189894
R2949 VN.n18 VN.n17 0.189894
R2950 VN.n18 VN.n0 0.189894
R2951 VN.n22 VN.n0 0.189894
R2952 VN VN.n22 0.0516364
R2953 VDD2.n2 VDD2.n1 63.9331
R2954 VDD2.n2 VDD2.n0 63.9331
R2955 VDD2 VDD2.n5 63.9303
R2956 VDD2.n4 VDD2.n3 63.105
R2957 VDD2.n4 VDD2.n2 45.6334
R2958 VDD2.n5 VDD2.t7 1.22272
R2959 VDD2.n5 VDD2.t3 1.22272
R2960 VDD2.n3 VDD2.t4 1.22272
R2961 VDD2.n3 VDD2.t2 1.22272
R2962 VDD2.n1 VDD2.t0 1.22272
R2963 VDD2.n1 VDD2.t5 1.22272
R2964 VDD2.n0 VDD2.t1 1.22272
R2965 VDD2.n0 VDD2.t6 1.22272
R2966 VDD2 VDD2.n4 0.94231
C0 VTAIL VDD2 10.091f
C1 VN VDD1 0.150122f
C2 VN VP 7.36002f
C3 VTAIL VDD1 10.0425f
C4 VTAIL VP 10.4463f
C5 VDD1 VDD2 1.31716f
C6 VDD2 VP 0.426015f
C7 VDD1 VP 10.7722f
C8 VN VTAIL 10.4322f
C9 VN VDD2 10.497201f
C10 VDD2 B 4.822366f
C11 VDD1 B 5.163188f
C12 VTAIL B 12.278193f
C13 VN B 12.578011f
C14 VP B 10.90972f
C15 VDD2.t1 B 0.317797f
C16 VDD2.t6 B 0.317797f
C17 VDD2.n0 B 2.89048f
C18 VDD2.t0 B 0.317797f
C19 VDD2.t5 B 0.317797f
C20 VDD2.n1 B 2.89048f
C21 VDD2.n2 B 3.00388f
C22 VDD2.t4 B 0.317797f
C23 VDD2.t2 B 0.317797f
C24 VDD2.n3 B 2.88504f
C25 VDD2.n4 B 2.94195f
C26 VDD2.t7 B 0.317797f
C27 VDD2.t3 B 0.317797f
C28 VDD2.n5 B 2.89045f
C29 VN.n0 B 0.027953f
C30 VN.t2 B 2.13788f
C31 VN.n1 B 0.02348f
C32 VN.n2 B 0.027953f
C33 VN.t7 B 2.13788f
C34 VN.n3 B 0.022577f
C35 VN.n4 B 0.178863f
C36 VN.t1 B 2.13788f
C37 VN.t6 B 2.23845f
C38 VN.n5 B 0.828494f
C39 VN.n6 B 0.80138f
C40 VN.n7 B 0.027525f
C41 VN.n8 B 0.055264f
C42 VN.n9 B 0.027953f
C43 VN.n10 B 0.027953f
C44 VN.n11 B 0.027953f
C45 VN.n12 B 0.055264f
C46 VN.n13 B 0.027525f
C47 VN.n14 B 0.753187f
C48 VN.n15 B 0.054865f
C49 VN.n16 B 0.027953f
C50 VN.n17 B 0.027953f
C51 VN.n18 B 0.027953f
C52 VN.n19 B 0.053479f
C53 VN.n20 B 0.030085f
C54 VN.n21 B 0.812442f
C55 VN.n22 B 0.029341f
C56 VN.n23 B 0.027953f
C57 VN.t3 B 2.13788f
C58 VN.n24 B 0.02348f
C59 VN.n25 B 0.027953f
C60 VN.t5 B 2.13788f
C61 VN.n26 B 0.022577f
C62 VN.n27 B 0.178863f
C63 VN.t0 B 2.13788f
C64 VN.t4 B 2.23845f
C65 VN.n28 B 0.828494f
C66 VN.n29 B 0.80138f
C67 VN.n30 B 0.027525f
C68 VN.n31 B 0.055264f
C69 VN.n32 B 0.027953f
C70 VN.n33 B 0.027953f
C71 VN.n34 B 0.027953f
C72 VN.n35 B 0.055264f
C73 VN.n36 B 0.027525f
C74 VN.n37 B 0.753187f
C75 VN.n38 B 0.054865f
C76 VN.n39 B 0.027953f
C77 VN.n40 B 0.027953f
C78 VN.n41 B 0.027953f
C79 VN.n42 B 0.053479f
C80 VN.n43 B 0.030085f
C81 VN.n44 B 0.812442f
C82 VN.n45 B 1.53829f
C83 VDD1.t6 B 0.319461f
C84 VDD1.t2 B 0.319461f
C85 VDD1.n0 B 2.90648f
C86 VDD1.t0 B 0.319461f
C87 VDD1.t3 B 0.319461f
C88 VDD1.n1 B 2.90561f
C89 VDD1.t5 B 0.319461f
C90 VDD1.t1 B 0.319461f
C91 VDD1.n2 B 2.90561f
C92 VDD1.n3 B 3.07191f
C93 VDD1.t4 B 0.319461f
C94 VDD1.t7 B 0.319461f
C95 VDD1.n4 B 2.90013f
C96 VDD1.n5 B 2.98786f
C97 VTAIL.t2 B 0.23671f
C98 VTAIL.t4 B 0.23671f
C99 VTAIL.n0 B 2.09611f
C100 VTAIL.n1 B 0.286898f
C101 VTAIL.n2 B 0.02599f
C102 VTAIL.n3 B 0.01849f
C103 VTAIL.n4 B 0.009936f
C104 VTAIL.n5 B 0.023485f
C105 VTAIL.n6 B 0.01052f
C106 VTAIL.n7 B 0.01849f
C107 VTAIL.n8 B 0.010228f
C108 VTAIL.n9 B 0.023485f
C109 VTAIL.n10 B 0.01052f
C110 VTAIL.n11 B 0.01849f
C111 VTAIL.n12 B 0.009936f
C112 VTAIL.n13 B 0.023485f
C113 VTAIL.n14 B 0.01052f
C114 VTAIL.n15 B 0.01849f
C115 VTAIL.n16 B 0.009936f
C116 VTAIL.n17 B 0.023485f
C117 VTAIL.n18 B 0.01052f
C118 VTAIL.n19 B 0.01849f
C119 VTAIL.n20 B 0.009936f
C120 VTAIL.n21 B 0.023485f
C121 VTAIL.n22 B 0.01052f
C122 VTAIL.n23 B 0.01849f
C123 VTAIL.n24 B 0.009936f
C124 VTAIL.n25 B 0.023485f
C125 VTAIL.n26 B 0.01052f
C126 VTAIL.n27 B 0.01849f
C127 VTAIL.n28 B 0.009936f
C128 VTAIL.n29 B 0.017614f
C129 VTAIL.n30 B 0.013873f
C130 VTAIL.t3 B 0.0388f
C131 VTAIL.n31 B 0.126162f
C132 VTAIL.n32 B 1.30471f
C133 VTAIL.n33 B 0.009936f
C134 VTAIL.n34 B 0.01052f
C135 VTAIL.n35 B 0.023485f
C136 VTAIL.n36 B 0.023485f
C137 VTAIL.n37 B 0.01052f
C138 VTAIL.n38 B 0.009936f
C139 VTAIL.n39 B 0.01849f
C140 VTAIL.n40 B 0.01849f
C141 VTAIL.n41 B 0.009936f
C142 VTAIL.n42 B 0.01052f
C143 VTAIL.n43 B 0.023485f
C144 VTAIL.n44 B 0.023485f
C145 VTAIL.n45 B 0.01052f
C146 VTAIL.n46 B 0.009936f
C147 VTAIL.n47 B 0.01849f
C148 VTAIL.n48 B 0.01849f
C149 VTAIL.n49 B 0.009936f
C150 VTAIL.n50 B 0.01052f
C151 VTAIL.n51 B 0.023485f
C152 VTAIL.n52 B 0.023485f
C153 VTAIL.n53 B 0.01052f
C154 VTAIL.n54 B 0.009936f
C155 VTAIL.n55 B 0.01849f
C156 VTAIL.n56 B 0.01849f
C157 VTAIL.n57 B 0.009936f
C158 VTAIL.n58 B 0.01052f
C159 VTAIL.n59 B 0.023485f
C160 VTAIL.n60 B 0.023485f
C161 VTAIL.n61 B 0.01052f
C162 VTAIL.n62 B 0.009936f
C163 VTAIL.n63 B 0.01849f
C164 VTAIL.n64 B 0.01849f
C165 VTAIL.n65 B 0.009936f
C166 VTAIL.n66 B 0.01052f
C167 VTAIL.n67 B 0.023485f
C168 VTAIL.n68 B 0.023485f
C169 VTAIL.n69 B 0.01052f
C170 VTAIL.n70 B 0.009936f
C171 VTAIL.n71 B 0.01849f
C172 VTAIL.n72 B 0.01849f
C173 VTAIL.n73 B 0.009936f
C174 VTAIL.n74 B 0.009936f
C175 VTAIL.n75 B 0.01052f
C176 VTAIL.n76 B 0.023485f
C177 VTAIL.n77 B 0.023485f
C178 VTAIL.n78 B 0.023485f
C179 VTAIL.n79 B 0.010228f
C180 VTAIL.n80 B 0.009936f
C181 VTAIL.n81 B 0.01849f
C182 VTAIL.n82 B 0.01849f
C183 VTAIL.n83 B 0.009936f
C184 VTAIL.n84 B 0.01052f
C185 VTAIL.n85 B 0.023485f
C186 VTAIL.n86 B 0.050841f
C187 VTAIL.n87 B 0.01052f
C188 VTAIL.n88 B 0.009936f
C189 VTAIL.n89 B 0.045771f
C190 VTAIL.n90 B 0.028538f
C191 VTAIL.n91 B 0.150791f
C192 VTAIL.n92 B 0.02599f
C193 VTAIL.n93 B 0.01849f
C194 VTAIL.n94 B 0.009936f
C195 VTAIL.n95 B 0.023485f
C196 VTAIL.n96 B 0.01052f
C197 VTAIL.n97 B 0.01849f
C198 VTAIL.n98 B 0.010228f
C199 VTAIL.n99 B 0.023485f
C200 VTAIL.n100 B 0.01052f
C201 VTAIL.n101 B 0.01849f
C202 VTAIL.n102 B 0.009936f
C203 VTAIL.n103 B 0.023485f
C204 VTAIL.n104 B 0.01052f
C205 VTAIL.n105 B 0.01849f
C206 VTAIL.n106 B 0.009936f
C207 VTAIL.n107 B 0.023485f
C208 VTAIL.n108 B 0.01052f
C209 VTAIL.n109 B 0.01849f
C210 VTAIL.n110 B 0.009936f
C211 VTAIL.n111 B 0.023485f
C212 VTAIL.n112 B 0.01052f
C213 VTAIL.n113 B 0.01849f
C214 VTAIL.n114 B 0.009936f
C215 VTAIL.n115 B 0.023485f
C216 VTAIL.n116 B 0.01052f
C217 VTAIL.n117 B 0.01849f
C218 VTAIL.n118 B 0.009936f
C219 VTAIL.n119 B 0.017614f
C220 VTAIL.n120 B 0.013873f
C221 VTAIL.t8 B 0.0388f
C222 VTAIL.n121 B 0.126162f
C223 VTAIL.n122 B 1.30471f
C224 VTAIL.n123 B 0.009936f
C225 VTAIL.n124 B 0.01052f
C226 VTAIL.n125 B 0.023485f
C227 VTAIL.n126 B 0.023485f
C228 VTAIL.n127 B 0.01052f
C229 VTAIL.n128 B 0.009936f
C230 VTAIL.n129 B 0.01849f
C231 VTAIL.n130 B 0.01849f
C232 VTAIL.n131 B 0.009936f
C233 VTAIL.n132 B 0.01052f
C234 VTAIL.n133 B 0.023485f
C235 VTAIL.n134 B 0.023485f
C236 VTAIL.n135 B 0.01052f
C237 VTAIL.n136 B 0.009936f
C238 VTAIL.n137 B 0.01849f
C239 VTAIL.n138 B 0.01849f
C240 VTAIL.n139 B 0.009936f
C241 VTAIL.n140 B 0.01052f
C242 VTAIL.n141 B 0.023485f
C243 VTAIL.n142 B 0.023485f
C244 VTAIL.n143 B 0.01052f
C245 VTAIL.n144 B 0.009936f
C246 VTAIL.n145 B 0.01849f
C247 VTAIL.n146 B 0.01849f
C248 VTAIL.n147 B 0.009936f
C249 VTAIL.n148 B 0.01052f
C250 VTAIL.n149 B 0.023485f
C251 VTAIL.n150 B 0.023485f
C252 VTAIL.n151 B 0.01052f
C253 VTAIL.n152 B 0.009936f
C254 VTAIL.n153 B 0.01849f
C255 VTAIL.n154 B 0.01849f
C256 VTAIL.n155 B 0.009936f
C257 VTAIL.n156 B 0.01052f
C258 VTAIL.n157 B 0.023485f
C259 VTAIL.n158 B 0.023485f
C260 VTAIL.n159 B 0.01052f
C261 VTAIL.n160 B 0.009936f
C262 VTAIL.n161 B 0.01849f
C263 VTAIL.n162 B 0.01849f
C264 VTAIL.n163 B 0.009936f
C265 VTAIL.n164 B 0.009936f
C266 VTAIL.n165 B 0.01052f
C267 VTAIL.n166 B 0.023485f
C268 VTAIL.n167 B 0.023485f
C269 VTAIL.n168 B 0.023485f
C270 VTAIL.n169 B 0.010228f
C271 VTAIL.n170 B 0.009936f
C272 VTAIL.n171 B 0.01849f
C273 VTAIL.n172 B 0.01849f
C274 VTAIL.n173 B 0.009936f
C275 VTAIL.n174 B 0.01052f
C276 VTAIL.n175 B 0.023485f
C277 VTAIL.n176 B 0.050841f
C278 VTAIL.n177 B 0.01052f
C279 VTAIL.n178 B 0.009936f
C280 VTAIL.n179 B 0.045771f
C281 VTAIL.n180 B 0.028538f
C282 VTAIL.n181 B 0.150791f
C283 VTAIL.t9 B 0.23671f
C284 VTAIL.t12 B 0.23671f
C285 VTAIL.n182 B 2.09611f
C286 VTAIL.n183 B 0.388724f
C287 VTAIL.n184 B 0.02599f
C288 VTAIL.n185 B 0.01849f
C289 VTAIL.n186 B 0.009936f
C290 VTAIL.n187 B 0.023485f
C291 VTAIL.n188 B 0.01052f
C292 VTAIL.n189 B 0.01849f
C293 VTAIL.n190 B 0.010228f
C294 VTAIL.n191 B 0.023485f
C295 VTAIL.n192 B 0.01052f
C296 VTAIL.n193 B 0.01849f
C297 VTAIL.n194 B 0.009936f
C298 VTAIL.n195 B 0.023485f
C299 VTAIL.n196 B 0.01052f
C300 VTAIL.n197 B 0.01849f
C301 VTAIL.n198 B 0.009936f
C302 VTAIL.n199 B 0.023485f
C303 VTAIL.n200 B 0.01052f
C304 VTAIL.n201 B 0.01849f
C305 VTAIL.n202 B 0.009936f
C306 VTAIL.n203 B 0.023485f
C307 VTAIL.n204 B 0.01052f
C308 VTAIL.n205 B 0.01849f
C309 VTAIL.n206 B 0.009936f
C310 VTAIL.n207 B 0.023485f
C311 VTAIL.n208 B 0.01052f
C312 VTAIL.n209 B 0.01849f
C313 VTAIL.n210 B 0.009936f
C314 VTAIL.n211 B 0.017614f
C315 VTAIL.n212 B 0.013873f
C316 VTAIL.t13 B 0.0388f
C317 VTAIL.n213 B 0.126162f
C318 VTAIL.n214 B 1.30471f
C319 VTAIL.n215 B 0.009936f
C320 VTAIL.n216 B 0.01052f
C321 VTAIL.n217 B 0.023485f
C322 VTAIL.n218 B 0.023485f
C323 VTAIL.n219 B 0.01052f
C324 VTAIL.n220 B 0.009936f
C325 VTAIL.n221 B 0.01849f
C326 VTAIL.n222 B 0.01849f
C327 VTAIL.n223 B 0.009936f
C328 VTAIL.n224 B 0.01052f
C329 VTAIL.n225 B 0.023485f
C330 VTAIL.n226 B 0.023485f
C331 VTAIL.n227 B 0.01052f
C332 VTAIL.n228 B 0.009936f
C333 VTAIL.n229 B 0.01849f
C334 VTAIL.n230 B 0.01849f
C335 VTAIL.n231 B 0.009936f
C336 VTAIL.n232 B 0.01052f
C337 VTAIL.n233 B 0.023485f
C338 VTAIL.n234 B 0.023485f
C339 VTAIL.n235 B 0.01052f
C340 VTAIL.n236 B 0.009936f
C341 VTAIL.n237 B 0.01849f
C342 VTAIL.n238 B 0.01849f
C343 VTAIL.n239 B 0.009936f
C344 VTAIL.n240 B 0.01052f
C345 VTAIL.n241 B 0.023485f
C346 VTAIL.n242 B 0.023485f
C347 VTAIL.n243 B 0.01052f
C348 VTAIL.n244 B 0.009936f
C349 VTAIL.n245 B 0.01849f
C350 VTAIL.n246 B 0.01849f
C351 VTAIL.n247 B 0.009936f
C352 VTAIL.n248 B 0.01052f
C353 VTAIL.n249 B 0.023485f
C354 VTAIL.n250 B 0.023485f
C355 VTAIL.n251 B 0.01052f
C356 VTAIL.n252 B 0.009936f
C357 VTAIL.n253 B 0.01849f
C358 VTAIL.n254 B 0.01849f
C359 VTAIL.n255 B 0.009936f
C360 VTAIL.n256 B 0.009936f
C361 VTAIL.n257 B 0.01052f
C362 VTAIL.n258 B 0.023485f
C363 VTAIL.n259 B 0.023485f
C364 VTAIL.n260 B 0.023485f
C365 VTAIL.n261 B 0.010228f
C366 VTAIL.n262 B 0.009936f
C367 VTAIL.n263 B 0.01849f
C368 VTAIL.n264 B 0.01849f
C369 VTAIL.n265 B 0.009936f
C370 VTAIL.n266 B 0.01052f
C371 VTAIL.n267 B 0.023485f
C372 VTAIL.n268 B 0.050841f
C373 VTAIL.n269 B 0.01052f
C374 VTAIL.n270 B 0.009936f
C375 VTAIL.n271 B 0.045771f
C376 VTAIL.n272 B 0.028538f
C377 VTAIL.n273 B 1.31133f
C378 VTAIL.n274 B 0.02599f
C379 VTAIL.n275 B 0.01849f
C380 VTAIL.n276 B 0.009936f
C381 VTAIL.n277 B 0.023485f
C382 VTAIL.n278 B 0.01052f
C383 VTAIL.n279 B 0.01849f
C384 VTAIL.n280 B 0.010228f
C385 VTAIL.n281 B 0.023485f
C386 VTAIL.n282 B 0.009936f
C387 VTAIL.n283 B 0.01052f
C388 VTAIL.n284 B 0.01849f
C389 VTAIL.n285 B 0.009936f
C390 VTAIL.n286 B 0.023485f
C391 VTAIL.n287 B 0.01052f
C392 VTAIL.n288 B 0.01849f
C393 VTAIL.n289 B 0.009936f
C394 VTAIL.n290 B 0.023485f
C395 VTAIL.n291 B 0.01052f
C396 VTAIL.n292 B 0.01849f
C397 VTAIL.n293 B 0.009936f
C398 VTAIL.n294 B 0.023485f
C399 VTAIL.n295 B 0.01052f
C400 VTAIL.n296 B 0.01849f
C401 VTAIL.n297 B 0.009936f
C402 VTAIL.n298 B 0.023485f
C403 VTAIL.n299 B 0.01052f
C404 VTAIL.n300 B 0.01849f
C405 VTAIL.n301 B 0.009936f
C406 VTAIL.n302 B 0.017614f
C407 VTAIL.n303 B 0.013873f
C408 VTAIL.t6 B 0.0388f
C409 VTAIL.n304 B 0.126162f
C410 VTAIL.n305 B 1.30471f
C411 VTAIL.n306 B 0.009936f
C412 VTAIL.n307 B 0.01052f
C413 VTAIL.n308 B 0.023485f
C414 VTAIL.n309 B 0.023485f
C415 VTAIL.n310 B 0.01052f
C416 VTAIL.n311 B 0.009936f
C417 VTAIL.n312 B 0.01849f
C418 VTAIL.n313 B 0.01849f
C419 VTAIL.n314 B 0.009936f
C420 VTAIL.n315 B 0.01052f
C421 VTAIL.n316 B 0.023485f
C422 VTAIL.n317 B 0.023485f
C423 VTAIL.n318 B 0.01052f
C424 VTAIL.n319 B 0.009936f
C425 VTAIL.n320 B 0.01849f
C426 VTAIL.n321 B 0.01849f
C427 VTAIL.n322 B 0.009936f
C428 VTAIL.n323 B 0.01052f
C429 VTAIL.n324 B 0.023485f
C430 VTAIL.n325 B 0.023485f
C431 VTAIL.n326 B 0.01052f
C432 VTAIL.n327 B 0.009936f
C433 VTAIL.n328 B 0.01849f
C434 VTAIL.n329 B 0.01849f
C435 VTAIL.n330 B 0.009936f
C436 VTAIL.n331 B 0.01052f
C437 VTAIL.n332 B 0.023485f
C438 VTAIL.n333 B 0.023485f
C439 VTAIL.n334 B 0.01052f
C440 VTAIL.n335 B 0.009936f
C441 VTAIL.n336 B 0.01849f
C442 VTAIL.n337 B 0.01849f
C443 VTAIL.n338 B 0.009936f
C444 VTAIL.n339 B 0.01052f
C445 VTAIL.n340 B 0.023485f
C446 VTAIL.n341 B 0.023485f
C447 VTAIL.n342 B 0.01052f
C448 VTAIL.n343 B 0.009936f
C449 VTAIL.n344 B 0.01849f
C450 VTAIL.n345 B 0.01849f
C451 VTAIL.n346 B 0.009936f
C452 VTAIL.n347 B 0.01052f
C453 VTAIL.n348 B 0.023485f
C454 VTAIL.n349 B 0.023485f
C455 VTAIL.n350 B 0.023485f
C456 VTAIL.n351 B 0.010228f
C457 VTAIL.n352 B 0.009936f
C458 VTAIL.n353 B 0.01849f
C459 VTAIL.n354 B 0.01849f
C460 VTAIL.n355 B 0.009936f
C461 VTAIL.n356 B 0.01052f
C462 VTAIL.n357 B 0.023485f
C463 VTAIL.n358 B 0.050841f
C464 VTAIL.n359 B 0.01052f
C465 VTAIL.n360 B 0.009936f
C466 VTAIL.n361 B 0.045771f
C467 VTAIL.n362 B 0.028538f
C468 VTAIL.n363 B 1.31133f
C469 VTAIL.t0 B 0.23671f
C470 VTAIL.t1 B 0.23671f
C471 VTAIL.n364 B 2.09612f
C472 VTAIL.n365 B 0.388715f
C473 VTAIL.n366 B 0.02599f
C474 VTAIL.n367 B 0.01849f
C475 VTAIL.n368 B 0.009936f
C476 VTAIL.n369 B 0.023485f
C477 VTAIL.n370 B 0.01052f
C478 VTAIL.n371 B 0.01849f
C479 VTAIL.n372 B 0.010228f
C480 VTAIL.n373 B 0.023485f
C481 VTAIL.n374 B 0.009936f
C482 VTAIL.n375 B 0.01052f
C483 VTAIL.n376 B 0.01849f
C484 VTAIL.n377 B 0.009936f
C485 VTAIL.n378 B 0.023485f
C486 VTAIL.n379 B 0.01052f
C487 VTAIL.n380 B 0.01849f
C488 VTAIL.n381 B 0.009936f
C489 VTAIL.n382 B 0.023485f
C490 VTAIL.n383 B 0.01052f
C491 VTAIL.n384 B 0.01849f
C492 VTAIL.n385 B 0.009936f
C493 VTAIL.n386 B 0.023485f
C494 VTAIL.n387 B 0.01052f
C495 VTAIL.n388 B 0.01849f
C496 VTAIL.n389 B 0.009936f
C497 VTAIL.n390 B 0.023485f
C498 VTAIL.n391 B 0.01052f
C499 VTAIL.n392 B 0.01849f
C500 VTAIL.n393 B 0.009936f
C501 VTAIL.n394 B 0.017614f
C502 VTAIL.n395 B 0.013873f
C503 VTAIL.t7 B 0.0388f
C504 VTAIL.n396 B 0.126162f
C505 VTAIL.n397 B 1.30471f
C506 VTAIL.n398 B 0.009936f
C507 VTAIL.n399 B 0.01052f
C508 VTAIL.n400 B 0.023485f
C509 VTAIL.n401 B 0.023485f
C510 VTAIL.n402 B 0.01052f
C511 VTAIL.n403 B 0.009936f
C512 VTAIL.n404 B 0.01849f
C513 VTAIL.n405 B 0.01849f
C514 VTAIL.n406 B 0.009936f
C515 VTAIL.n407 B 0.01052f
C516 VTAIL.n408 B 0.023485f
C517 VTAIL.n409 B 0.023485f
C518 VTAIL.n410 B 0.01052f
C519 VTAIL.n411 B 0.009936f
C520 VTAIL.n412 B 0.01849f
C521 VTAIL.n413 B 0.01849f
C522 VTAIL.n414 B 0.009936f
C523 VTAIL.n415 B 0.01052f
C524 VTAIL.n416 B 0.023485f
C525 VTAIL.n417 B 0.023485f
C526 VTAIL.n418 B 0.01052f
C527 VTAIL.n419 B 0.009936f
C528 VTAIL.n420 B 0.01849f
C529 VTAIL.n421 B 0.01849f
C530 VTAIL.n422 B 0.009936f
C531 VTAIL.n423 B 0.01052f
C532 VTAIL.n424 B 0.023485f
C533 VTAIL.n425 B 0.023485f
C534 VTAIL.n426 B 0.01052f
C535 VTAIL.n427 B 0.009936f
C536 VTAIL.n428 B 0.01849f
C537 VTAIL.n429 B 0.01849f
C538 VTAIL.n430 B 0.009936f
C539 VTAIL.n431 B 0.01052f
C540 VTAIL.n432 B 0.023485f
C541 VTAIL.n433 B 0.023485f
C542 VTAIL.n434 B 0.01052f
C543 VTAIL.n435 B 0.009936f
C544 VTAIL.n436 B 0.01849f
C545 VTAIL.n437 B 0.01849f
C546 VTAIL.n438 B 0.009936f
C547 VTAIL.n439 B 0.01052f
C548 VTAIL.n440 B 0.023485f
C549 VTAIL.n441 B 0.023485f
C550 VTAIL.n442 B 0.023485f
C551 VTAIL.n443 B 0.010228f
C552 VTAIL.n444 B 0.009936f
C553 VTAIL.n445 B 0.01849f
C554 VTAIL.n446 B 0.01849f
C555 VTAIL.n447 B 0.009936f
C556 VTAIL.n448 B 0.01052f
C557 VTAIL.n449 B 0.023485f
C558 VTAIL.n450 B 0.050841f
C559 VTAIL.n451 B 0.01052f
C560 VTAIL.n452 B 0.009936f
C561 VTAIL.n453 B 0.045771f
C562 VTAIL.n454 B 0.028538f
C563 VTAIL.n455 B 0.150791f
C564 VTAIL.n456 B 0.02599f
C565 VTAIL.n457 B 0.01849f
C566 VTAIL.n458 B 0.009936f
C567 VTAIL.n459 B 0.023485f
C568 VTAIL.n460 B 0.01052f
C569 VTAIL.n461 B 0.01849f
C570 VTAIL.n462 B 0.010228f
C571 VTAIL.n463 B 0.023485f
C572 VTAIL.n464 B 0.009936f
C573 VTAIL.n465 B 0.01052f
C574 VTAIL.n466 B 0.01849f
C575 VTAIL.n467 B 0.009936f
C576 VTAIL.n468 B 0.023485f
C577 VTAIL.n469 B 0.01052f
C578 VTAIL.n470 B 0.01849f
C579 VTAIL.n471 B 0.009936f
C580 VTAIL.n472 B 0.023485f
C581 VTAIL.n473 B 0.01052f
C582 VTAIL.n474 B 0.01849f
C583 VTAIL.n475 B 0.009936f
C584 VTAIL.n476 B 0.023485f
C585 VTAIL.n477 B 0.01052f
C586 VTAIL.n478 B 0.01849f
C587 VTAIL.n479 B 0.009936f
C588 VTAIL.n480 B 0.023485f
C589 VTAIL.n481 B 0.01052f
C590 VTAIL.n482 B 0.01849f
C591 VTAIL.n483 B 0.009936f
C592 VTAIL.n484 B 0.017614f
C593 VTAIL.n485 B 0.013873f
C594 VTAIL.t10 B 0.0388f
C595 VTAIL.n486 B 0.126162f
C596 VTAIL.n487 B 1.30471f
C597 VTAIL.n488 B 0.009936f
C598 VTAIL.n489 B 0.01052f
C599 VTAIL.n490 B 0.023485f
C600 VTAIL.n491 B 0.023485f
C601 VTAIL.n492 B 0.01052f
C602 VTAIL.n493 B 0.009936f
C603 VTAIL.n494 B 0.01849f
C604 VTAIL.n495 B 0.01849f
C605 VTAIL.n496 B 0.009936f
C606 VTAIL.n497 B 0.01052f
C607 VTAIL.n498 B 0.023485f
C608 VTAIL.n499 B 0.023485f
C609 VTAIL.n500 B 0.01052f
C610 VTAIL.n501 B 0.009936f
C611 VTAIL.n502 B 0.01849f
C612 VTAIL.n503 B 0.01849f
C613 VTAIL.n504 B 0.009936f
C614 VTAIL.n505 B 0.01052f
C615 VTAIL.n506 B 0.023485f
C616 VTAIL.n507 B 0.023485f
C617 VTAIL.n508 B 0.01052f
C618 VTAIL.n509 B 0.009936f
C619 VTAIL.n510 B 0.01849f
C620 VTAIL.n511 B 0.01849f
C621 VTAIL.n512 B 0.009936f
C622 VTAIL.n513 B 0.01052f
C623 VTAIL.n514 B 0.023485f
C624 VTAIL.n515 B 0.023485f
C625 VTAIL.n516 B 0.01052f
C626 VTAIL.n517 B 0.009936f
C627 VTAIL.n518 B 0.01849f
C628 VTAIL.n519 B 0.01849f
C629 VTAIL.n520 B 0.009936f
C630 VTAIL.n521 B 0.01052f
C631 VTAIL.n522 B 0.023485f
C632 VTAIL.n523 B 0.023485f
C633 VTAIL.n524 B 0.01052f
C634 VTAIL.n525 B 0.009936f
C635 VTAIL.n526 B 0.01849f
C636 VTAIL.n527 B 0.01849f
C637 VTAIL.n528 B 0.009936f
C638 VTAIL.n529 B 0.01052f
C639 VTAIL.n530 B 0.023485f
C640 VTAIL.n531 B 0.023485f
C641 VTAIL.n532 B 0.023485f
C642 VTAIL.n533 B 0.010228f
C643 VTAIL.n534 B 0.009936f
C644 VTAIL.n535 B 0.01849f
C645 VTAIL.n536 B 0.01849f
C646 VTAIL.n537 B 0.009936f
C647 VTAIL.n538 B 0.01052f
C648 VTAIL.n539 B 0.023485f
C649 VTAIL.n540 B 0.050841f
C650 VTAIL.n541 B 0.01052f
C651 VTAIL.n542 B 0.009936f
C652 VTAIL.n543 B 0.045771f
C653 VTAIL.n544 B 0.028538f
C654 VTAIL.n545 B 0.150791f
C655 VTAIL.t11 B 0.23671f
C656 VTAIL.t14 B 0.23671f
C657 VTAIL.n546 B 2.09612f
C658 VTAIL.n547 B 0.388715f
C659 VTAIL.n548 B 0.02599f
C660 VTAIL.n549 B 0.01849f
C661 VTAIL.n550 B 0.009936f
C662 VTAIL.n551 B 0.023485f
C663 VTAIL.n552 B 0.01052f
C664 VTAIL.n553 B 0.01849f
C665 VTAIL.n554 B 0.010228f
C666 VTAIL.n555 B 0.023485f
C667 VTAIL.n556 B 0.009936f
C668 VTAIL.n557 B 0.01052f
C669 VTAIL.n558 B 0.01849f
C670 VTAIL.n559 B 0.009936f
C671 VTAIL.n560 B 0.023485f
C672 VTAIL.n561 B 0.01052f
C673 VTAIL.n562 B 0.01849f
C674 VTAIL.n563 B 0.009936f
C675 VTAIL.n564 B 0.023485f
C676 VTAIL.n565 B 0.01052f
C677 VTAIL.n566 B 0.01849f
C678 VTAIL.n567 B 0.009936f
C679 VTAIL.n568 B 0.023485f
C680 VTAIL.n569 B 0.01052f
C681 VTAIL.n570 B 0.01849f
C682 VTAIL.n571 B 0.009936f
C683 VTAIL.n572 B 0.023485f
C684 VTAIL.n573 B 0.01052f
C685 VTAIL.n574 B 0.01849f
C686 VTAIL.n575 B 0.009936f
C687 VTAIL.n576 B 0.017614f
C688 VTAIL.n577 B 0.013873f
C689 VTAIL.t15 B 0.0388f
C690 VTAIL.n578 B 0.126162f
C691 VTAIL.n579 B 1.30471f
C692 VTAIL.n580 B 0.009936f
C693 VTAIL.n581 B 0.01052f
C694 VTAIL.n582 B 0.023485f
C695 VTAIL.n583 B 0.023485f
C696 VTAIL.n584 B 0.01052f
C697 VTAIL.n585 B 0.009936f
C698 VTAIL.n586 B 0.01849f
C699 VTAIL.n587 B 0.01849f
C700 VTAIL.n588 B 0.009936f
C701 VTAIL.n589 B 0.01052f
C702 VTAIL.n590 B 0.023485f
C703 VTAIL.n591 B 0.023485f
C704 VTAIL.n592 B 0.01052f
C705 VTAIL.n593 B 0.009936f
C706 VTAIL.n594 B 0.01849f
C707 VTAIL.n595 B 0.01849f
C708 VTAIL.n596 B 0.009936f
C709 VTAIL.n597 B 0.01052f
C710 VTAIL.n598 B 0.023485f
C711 VTAIL.n599 B 0.023485f
C712 VTAIL.n600 B 0.01052f
C713 VTAIL.n601 B 0.009936f
C714 VTAIL.n602 B 0.01849f
C715 VTAIL.n603 B 0.01849f
C716 VTAIL.n604 B 0.009936f
C717 VTAIL.n605 B 0.01052f
C718 VTAIL.n606 B 0.023485f
C719 VTAIL.n607 B 0.023485f
C720 VTAIL.n608 B 0.01052f
C721 VTAIL.n609 B 0.009936f
C722 VTAIL.n610 B 0.01849f
C723 VTAIL.n611 B 0.01849f
C724 VTAIL.n612 B 0.009936f
C725 VTAIL.n613 B 0.01052f
C726 VTAIL.n614 B 0.023485f
C727 VTAIL.n615 B 0.023485f
C728 VTAIL.n616 B 0.01052f
C729 VTAIL.n617 B 0.009936f
C730 VTAIL.n618 B 0.01849f
C731 VTAIL.n619 B 0.01849f
C732 VTAIL.n620 B 0.009936f
C733 VTAIL.n621 B 0.01052f
C734 VTAIL.n622 B 0.023485f
C735 VTAIL.n623 B 0.023485f
C736 VTAIL.n624 B 0.023485f
C737 VTAIL.n625 B 0.010228f
C738 VTAIL.n626 B 0.009936f
C739 VTAIL.n627 B 0.01849f
C740 VTAIL.n628 B 0.01849f
C741 VTAIL.n629 B 0.009936f
C742 VTAIL.n630 B 0.01052f
C743 VTAIL.n631 B 0.023485f
C744 VTAIL.n632 B 0.050841f
C745 VTAIL.n633 B 0.01052f
C746 VTAIL.n634 B 0.009936f
C747 VTAIL.n635 B 0.045771f
C748 VTAIL.n636 B 0.028538f
C749 VTAIL.n637 B 1.31133f
C750 VTAIL.n638 B 0.02599f
C751 VTAIL.n639 B 0.01849f
C752 VTAIL.n640 B 0.009936f
C753 VTAIL.n641 B 0.023485f
C754 VTAIL.n642 B 0.01052f
C755 VTAIL.n643 B 0.01849f
C756 VTAIL.n644 B 0.010228f
C757 VTAIL.n645 B 0.023485f
C758 VTAIL.n646 B 0.01052f
C759 VTAIL.n647 B 0.01849f
C760 VTAIL.n648 B 0.009936f
C761 VTAIL.n649 B 0.023485f
C762 VTAIL.n650 B 0.01052f
C763 VTAIL.n651 B 0.01849f
C764 VTAIL.n652 B 0.009936f
C765 VTAIL.n653 B 0.023485f
C766 VTAIL.n654 B 0.01052f
C767 VTAIL.n655 B 0.01849f
C768 VTAIL.n656 B 0.009936f
C769 VTAIL.n657 B 0.023485f
C770 VTAIL.n658 B 0.01052f
C771 VTAIL.n659 B 0.01849f
C772 VTAIL.n660 B 0.009936f
C773 VTAIL.n661 B 0.023485f
C774 VTAIL.n662 B 0.01052f
C775 VTAIL.n663 B 0.01849f
C776 VTAIL.n664 B 0.009936f
C777 VTAIL.n665 B 0.017614f
C778 VTAIL.n666 B 0.013873f
C779 VTAIL.t5 B 0.0388f
C780 VTAIL.n667 B 0.126162f
C781 VTAIL.n668 B 1.30471f
C782 VTAIL.n669 B 0.009936f
C783 VTAIL.n670 B 0.01052f
C784 VTAIL.n671 B 0.023485f
C785 VTAIL.n672 B 0.023485f
C786 VTAIL.n673 B 0.01052f
C787 VTAIL.n674 B 0.009936f
C788 VTAIL.n675 B 0.01849f
C789 VTAIL.n676 B 0.01849f
C790 VTAIL.n677 B 0.009936f
C791 VTAIL.n678 B 0.01052f
C792 VTAIL.n679 B 0.023485f
C793 VTAIL.n680 B 0.023485f
C794 VTAIL.n681 B 0.01052f
C795 VTAIL.n682 B 0.009936f
C796 VTAIL.n683 B 0.01849f
C797 VTAIL.n684 B 0.01849f
C798 VTAIL.n685 B 0.009936f
C799 VTAIL.n686 B 0.01052f
C800 VTAIL.n687 B 0.023485f
C801 VTAIL.n688 B 0.023485f
C802 VTAIL.n689 B 0.01052f
C803 VTAIL.n690 B 0.009936f
C804 VTAIL.n691 B 0.01849f
C805 VTAIL.n692 B 0.01849f
C806 VTAIL.n693 B 0.009936f
C807 VTAIL.n694 B 0.01052f
C808 VTAIL.n695 B 0.023485f
C809 VTAIL.n696 B 0.023485f
C810 VTAIL.n697 B 0.01052f
C811 VTAIL.n698 B 0.009936f
C812 VTAIL.n699 B 0.01849f
C813 VTAIL.n700 B 0.01849f
C814 VTAIL.n701 B 0.009936f
C815 VTAIL.n702 B 0.01052f
C816 VTAIL.n703 B 0.023485f
C817 VTAIL.n704 B 0.023485f
C818 VTAIL.n705 B 0.01052f
C819 VTAIL.n706 B 0.009936f
C820 VTAIL.n707 B 0.01849f
C821 VTAIL.n708 B 0.01849f
C822 VTAIL.n709 B 0.009936f
C823 VTAIL.n710 B 0.009936f
C824 VTAIL.n711 B 0.01052f
C825 VTAIL.n712 B 0.023485f
C826 VTAIL.n713 B 0.023485f
C827 VTAIL.n714 B 0.023485f
C828 VTAIL.n715 B 0.010228f
C829 VTAIL.n716 B 0.009936f
C830 VTAIL.n717 B 0.01849f
C831 VTAIL.n718 B 0.01849f
C832 VTAIL.n719 B 0.009936f
C833 VTAIL.n720 B 0.01052f
C834 VTAIL.n721 B 0.023485f
C835 VTAIL.n722 B 0.050841f
C836 VTAIL.n723 B 0.01052f
C837 VTAIL.n724 B 0.009936f
C838 VTAIL.n725 B 0.045771f
C839 VTAIL.n726 B 0.028538f
C840 VTAIL.n727 B 1.30787f
C841 VP.n0 B 0.028288f
C842 VP.t6 B 2.16354f
C843 VP.n1 B 0.023762f
C844 VP.n2 B 0.028288f
C845 VP.t2 B 2.16354f
C846 VP.n3 B 0.022848f
C847 VP.n4 B 0.028288f
C848 VP.t4 B 2.16354f
C849 VP.n5 B 0.023762f
C850 VP.n6 B 0.028288f
C851 VP.t7 B 2.16354f
C852 VP.n7 B 0.028288f
C853 VP.t0 B 2.16354f
C854 VP.n8 B 0.023762f
C855 VP.n9 B 0.028288f
C856 VP.t3 B 2.16354f
C857 VP.n10 B 0.022848f
C858 VP.n11 B 0.18101f
C859 VP.t5 B 2.16354f
C860 VP.t1 B 2.26532f
C861 VP.n12 B 0.83844f
C862 VP.n13 B 0.811001f
C863 VP.n14 B 0.027856f
C864 VP.n15 B 0.055927f
C865 VP.n16 B 0.028288f
C866 VP.n17 B 0.028288f
C867 VP.n18 B 0.028288f
C868 VP.n19 B 0.055927f
C869 VP.n20 B 0.027856f
C870 VP.n21 B 0.762229f
C871 VP.n22 B 0.055524f
C872 VP.n23 B 0.028288f
C873 VP.n24 B 0.028288f
C874 VP.n25 B 0.028288f
C875 VP.n26 B 0.054121f
C876 VP.n27 B 0.030446f
C877 VP.n28 B 0.822196f
C878 VP.n29 B 1.53836f
C879 VP.n30 B 1.55882f
C880 VP.n31 B 0.822196f
C881 VP.n32 B 0.030446f
C882 VP.n33 B 0.054121f
C883 VP.n34 B 0.028288f
C884 VP.n35 B 0.028288f
C885 VP.n36 B 0.028288f
C886 VP.n37 B 0.055524f
C887 VP.n38 B 0.762229f
C888 VP.n39 B 0.027856f
C889 VP.n40 B 0.055927f
C890 VP.n41 B 0.028288f
C891 VP.n42 B 0.028288f
C892 VP.n43 B 0.028288f
C893 VP.n44 B 0.055927f
C894 VP.n45 B 0.027856f
C895 VP.n46 B 0.762229f
C896 VP.n47 B 0.055524f
C897 VP.n48 B 0.028288f
C898 VP.n49 B 0.028288f
C899 VP.n50 B 0.028288f
C900 VP.n51 B 0.054121f
C901 VP.n52 B 0.030446f
C902 VP.n53 B 0.822196f
C903 VP.n54 B 0.029694f
.ends

