* NGSPICE file created from diff_pair_sample_1140.ext - technology: sky130A

.subckt diff_pair_sample_1140 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=3.03
X1 B.t8 B.t6 B.t7 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=3.03
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=1.5483 ps=8.72 w=3.97 l=3.03
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=1.5483 ps=8.72 w=3.97 l=3.03
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=1.5483 ps=8.72 w=3.97 l=3.03
X5 VDD1.t0 VP.t1 VTAIL.t1 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=1.5483 ps=8.72 w=3.97 l=3.03
X6 B.t5 B.t3 B.t4 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=3.03
X7 B.t2 B.t0 B.t1 w_n2314_n1762# sky130_fd_pr__pfet_01v8 ad=1.5483 pd=8.72 as=0 ps=0 w=3.97 l=3.03
R0 B.n310 B.n43 585
R1 B.n312 B.n311 585
R2 B.n313 B.n42 585
R3 B.n315 B.n314 585
R4 B.n316 B.n41 585
R5 B.n318 B.n317 585
R6 B.n319 B.n40 585
R7 B.n321 B.n320 585
R8 B.n322 B.n39 585
R9 B.n324 B.n323 585
R10 B.n325 B.n38 585
R11 B.n327 B.n326 585
R12 B.n328 B.n37 585
R13 B.n330 B.n329 585
R14 B.n331 B.n36 585
R15 B.n333 B.n332 585
R16 B.n334 B.n35 585
R17 B.n336 B.n335 585
R18 B.n338 B.n337 585
R19 B.n339 B.n31 585
R20 B.n341 B.n340 585
R21 B.n342 B.n30 585
R22 B.n344 B.n343 585
R23 B.n345 B.n29 585
R24 B.n347 B.n346 585
R25 B.n348 B.n28 585
R26 B.n350 B.n349 585
R27 B.n351 B.n25 585
R28 B.n354 B.n353 585
R29 B.n355 B.n24 585
R30 B.n357 B.n356 585
R31 B.n358 B.n23 585
R32 B.n360 B.n359 585
R33 B.n361 B.n22 585
R34 B.n363 B.n362 585
R35 B.n364 B.n21 585
R36 B.n366 B.n365 585
R37 B.n367 B.n20 585
R38 B.n369 B.n368 585
R39 B.n370 B.n19 585
R40 B.n372 B.n371 585
R41 B.n373 B.n18 585
R42 B.n375 B.n374 585
R43 B.n376 B.n17 585
R44 B.n378 B.n377 585
R45 B.n379 B.n16 585
R46 B.n309 B.n308 585
R47 B.n307 B.n44 585
R48 B.n306 B.n305 585
R49 B.n304 B.n45 585
R50 B.n303 B.n302 585
R51 B.n301 B.n46 585
R52 B.n300 B.n299 585
R53 B.n298 B.n47 585
R54 B.n297 B.n296 585
R55 B.n295 B.n48 585
R56 B.n294 B.n293 585
R57 B.n292 B.n49 585
R58 B.n291 B.n290 585
R59 B.n289 B.n50 585
R60 B.n288 B.n287 585
R61 B.n286 B.n51 585
R62 B.n285 B.n284 585
R63 B.n283 B.n52 585
R64 B.n282 B.n281 585
R65 B.n280 B.n53 585
R66 B.n279 B.n278 585
R67 B.n277 B.n54 585
R68 B.n276 B.n275 585
R69 B.n274 B.n55 585
R70 B.n273 B.n272 585
R71 B.n271 B.n56 585
R72 B.n270 B.n269 585
R73 B.n268 B.n57 585
R74 B.n267 B.n266 585
R75 B.n265 B.n58 585
R76 B.n264 B.n263 585
R77 B.n262 B.n59 585
R78 B.n261 B.n260 585
R79 B.n259 B.n60 585
R80 B.n258 B.n257 585
R81 B.n256 B.n61 585
R82 B.n255 B.n254 585
R83 B.n253 B.n62 585
R84 B.n252 B.n251 585
R85 B.n250 B.n63 585
R86 B.n249 B.n248 585
R87 B.n247 B.n64 585
R88 B.n246 B.n245 585
R89 B.n244 B.n65 585
R90 B.n243 B.n242 585
R91 B.n241 B.n66 585
R92 B.n240 B.n239 585
R93 B.n238 B.n67 585
R94 B.n237 B.n236 585
R95 B.n235 B.n68 585
R96 B.n234 B.n233 585
R97 B.n232 B.n69 585
R98 B.n231 B.n230 585
R99 B.n229 B.n70 585
R100 B.n228 B.n227 585
R101 B.n226 B.n71 585
R102 B.n225 B.n224 585
R103 B.n154 B.n99 585
R104 B.n156 B.n155 585
R105 B.n157 B.n98 585
R106 B.n159 B.n158 585
R107 B.n160 B.n97 585
R108 B.n162 B.n161 585
R109 B.n163 B.n96 585
R110 B.n165 B.n164 585
R111 B.n166 B.n95 585
R112 B.n168 B.n167 585
R113 B.n169 B.n94 585
R114 B.n171 B.n170 585
R115 B.n172 B.n93 585
R116 B.n174 B.n173 585
R117 B.n175 B.n92 585
R118 B.n177 B.n176 585
R119 B.n178 B.n91 585
R120 B.n180 B.n179 585
R121 B.n182 B.n181 585
R122 B.n183 B.n87 585
R123 B.n185 B.n184 585
R124 B.n186 B.n86 585
R125 B.n188 B.n187 585
R126 B.n189 B.n85 585
R127 B.n191 B.n190 585
R128 B.n192 B.n84 585
R129 B.n194 B.n193 585
R130 B.n195 B.n81 585
R131 B.n198 B.n197 585
R132 B.n199 B.n80 585
R133 B.n201 B.n200 585
R134 B.n202 B.n79 585
R135 B.n204 B.n203 585
R136 B.n205 B.n78 585
R137 B.n207 B.n206 585
R138 B.n208 B.n77 585
R139 B.n210 B.n209 585
R140 B.n211 B.n76 585
R141 B.n213 B.n212 585
R142 B.n214 B.n75 585
R143 B.n216 B.n215 585
R144 B.n217 B.n74 585
R145 B.n219 B.n218 585
R146 B.n220 B.n73 585
R147 B.n222 B.n221 585
R148 B.n223 B.n72 585
R149 B.n153 B.n152 585
R150 B.n151 B.n100 585
R151 B.n150 B.n149 585
R152 B.n148 B.n101 585
R153 B.n147 B.n146 585
R154 B.n145 B.n102 585
R155 B.n144 B.n143 585
R156 B.n142 B.n103 585
R157 B.n141 B.n140 585
R158 B.n139 B.n104 585
R159 B.n138 B.n137 585
R160 B.n136 B.n105 585
R161 B.n135 B.n134 585
R162 B.n133 B.n106 585
R163 B.n132 B.n131 585
R164 B.n130 B.n107 585
R165 B.n129 B.n128 585
R166 B.n127 B.n108 585
R167 B.n126 B.n125 585
R168 B.n124 B.n109 585
R169 B.n123 B.n122 585
R170 B.n121 B.n110 585
R171 B.n120 B.n119 585
R172 B.n118 B.n111 585
R173 B.n117 B.n116 585
R174 B.n115 B.n112 585
R175 B.n114 B.n113 585
R176 B.n2 B.n0 585
R177 B.n421 B.n1 585
R178 B.n420 B.n419 585
R179 B.n418 B.n3 585
R180 B.n417 B.n416 585
R181 B.n415 B.n4 585
R182 B.n414 B.n413 585
R183 B.n412 B.n5 585
R184 B.n411 B.n410 585
R185 B.n409 B.n6 585
R186 B.n408 B.n407 585
R187 B.n406 B.n7 585
R188 B.n405 B.n404 585
R189 B.n403 B.n8 585
R190 B.n402 B.n401 585
R191 B.n400 B.n9 585
R192 B.n399 B.n398 585
R193 B.n397 B.n10 585
R194 B.n396 B.n395 585
R195 B.n394 B.n11 585
R196 B.n393 B.n392 585
R197 B.n391 B.n12 585
R198 B.n390 B.n389 585
R199 B.n388 B.n13 585
R200 B.n387 B.n386 585
R201 B.n385 B.n14 585
R202 B.n384 B.n383 585
R203 B.n382 B.n15 585
R204 B.n381 B.n380 585
R205 B.n423 B.n422 585
R206 B.n152 B.n99 444.452
R207 B.n380 B.n379 444.452
R208 B.n224 B.n223 444.452
R209 B.n308 B.n43 444.452
R210 B.n82 B.t5 300.406
R211 B.n32 B.t1 300.406
R212 B.n88 B.t8 300.406
R213 B.n26 B.t10 300.406
R214 B.n82 B.t3 240.859
R215 B.n32 B.t0 240.859
R216 B.n88 B.t6 240.567
R217 B.n26 B.t9 240.567
R218 B.n83 B.t4 235.242
R219 B.n33 B.t2 235.242
R220 B.n89 B.t7 235.242
R221 B.n27 B.t11 235.242
R222 B.n152 B.n151 163.367
R223 B.n151 B.n150 163.367
R224 B.n150 B.n101 163.367
R225 B.n146 B.n101 163.367
R226 B.n146 B.n145 163.367
R227 B.n145 B.n144 163.367
R228 B.n144 B.n103 163.367
R229 B.n140 B.n103 163.367
R230 B.n140 B.n139 163.367
R231 B.n139 B.n138 163.367
R232 B.n138 B.n105 163.367
R233 B.n134 B.n105 163.367
R234 B.n134 B.n133 163.367
R235 B.n133 B.n132 163.367
R236 B.n132 B.n107 163.367
R237 B.n128 B.n107 163.367
R238 B.n128 B.n127 163.367
R239 B.n127 B.n126 163.367
R240 B.n126 B.n109 163.367
R241 B.n122 B.n109 163.367
R242 B.n122 B.n121 163.367
R243 B.n121 B.n120 163.367
R244 B.n120 B.n111 163.367
R245 B.n116 B.n111 163.367
R246 B.n116 B.n115 163.367
R247 B.n115 B.n114 163.367
R248 B.n114 B.n2 163.367
R249 B.n422 B.n2 163.367
R250 B.n422 B.n421 163.367
R251 B.n421 B.n420 163.367
R252 B.n420 B.n3 163.367
R253 B.n416 B.n3 163.367
R254 B.n416 B.n415 163.367
R255 B.n415 B.n414 163.367
R256 B.n414 B.n5 163.367
R257 B.n410 B.n5 163.367
R258 B.n410 B.n409 163.367
R259 B.n409 B.n408 163.367
R260 B.n408 B.n7 163.367
R261 B.n404 B.n7 163.367
R262 B.n404 B.n403 163.367
R263 B.n403 B.n402 163.367
R264 B.n402 B.n9 163.367
R265 B.n398 B.n9 163.367
R266 B.n398 B.n397 163.367
R267 B.n397 B.n396 163.367
R268 B.n396 B.n11 163.367
R269 B.n392 B.n11 163.367
R270 B.n392 B.n391 163.367
R271 B.n391 B.n390 163.367
R272 B.n390 B.n13 163.367
R273 B.n386 B.n13 163.367
R274 B.n386 B.n385 163.367
R275 B.n385 B.n384 163.367
R276 B.n384 B.n15 163.367
R277 B.n380 B.n15 163.367
R278 B.n156 B.n99 163.367
R279 B.n157 B.n156 163.367
R280 B.n158 B.n157 163.367
R281 B.n158 B.n97 163.367
R282 B.n162 B.n97 163.367
R283 B.n163 B.n162 163.367
R284 B.n164 B.n163 163.367
R285 B.n164 B.n95 163.367
R286 B.n168 B.n95 163.367
R287 B.n169 B.n168 163.367
R288 B.n170 B.n169 163.367
R289 B.n170 B.n93 163.367
R290 B.n174 B.n93 163.367
R291 B.n175 B.n174 163.367
R292 B.n176 B.n175 163.367
R293 B.n176 B.n91 163.367
R294 B.n180 B.n91 163.367
R295 B.n181 B.n180 163.367
R296 B.n181 B.n87 163.367
R297 B.n185 B.n87 163.367
R298 B.n186 B.n185 163.367
R299 B.n187 B.n186 163.367
R300 B.n187 B.n85 163.367
R301 B.n191 B.n85 163.367
R302 B.n192 B.n191 163.367
R303 B.n193 B.n192 163.367
R304 B.n193 B.n81 163.367
R305 B.n198 B.n81 163.367
R306 B.n199 B.n198 163.367
R307 B.n200 B.n199 163.367
R308 B.n200 B.n79 163.367
R309 B.n204 B.n79 163.367
R310 B.n205 B.n204 163.367
R311 B.n206 B.n205 163.367
R312 B.n206 B.n77 163.367
R313 B.n210 B.n77 163.367
R314 B.n211 B.n210 163.367
R315 B.n212 B.n211 163.367
R316 B.n212 B.n75 163.367
R317 B.n216 B.n75 163.367
R318 B.n217 B.n216 163.367
R319 B.n218 B.n217 163.367
R320 B.n218 B.n73 163.367
R321 B.n222 B.n73 163.367
R322 B.n223 B.n222 163.367
R323 B.n224 B.n71 163.367
R324 B.n228 B.n71 163.367
R325 B.n229 B.n228 163.367
R326 B.n230 B.n229 163.367
R327 B.n230 B.n69 163.367
R328 B.n234 B.n69 163.367
R329 B.n235 B.n234 163.367
R330 B.n236 B.n235 163.367
R331 B.n236 B.n67 163.367
R332 B.n240 B.n67 163.367
R333 B.n241 B.n240 163.367
R334 B.n242 B.n241 163.367
R335 B.n242 B.n65 163.367
R336 B.n246 B.n65 163.367
R337 B.n247 B.n246 163.367
R338 B.n248 B.n247 163.367
R339 B.n248 B.n63 163.367
R340 B.n252 B.n63 163.367
R341 B.n253 B.n252 163.367
R342 B.n254 B.n253 163.367
R343 B.n254 B.n61 163.367
R344 B.n258 B.n61 163.367
R345 B.n259 B.n258 163.367
R346 B.n260 B.n259 163.367
R347 B.n260 B.n59 163.367
R348 B.n264 B.n59 163.367
R349 B.n265 B.n264 163.367
R350 B.n266 B.n265 163.367
R351 B.n266 B.n57 163.367
R352 B.n270 B.n57 163.367
R353 B.n271 B.n270 163.367
R354 B.n272 B.n271 163.367
R355 B.n272 B.n55 163.367
R356 B.n276 B.n55 163.367
R357 B.n277 B.n276 163.367
R358 B.n278 B.n277 163.367
R359 B.n278 B.n53 163.367
R360 B.n282 B.n53 163.367
R361 B.n283 B.n282 163.367
R362 B.n284 B.n283 163.367
R363 B.n284 B.n51 163.367
R364 B.n288 B.n51 163.367
R365 B.n289 B.n288 163.367
R366 B.n290 B.n289 163.367
R367 B.n290 B.n49 163.367
R368 B.n294 B.n49 163.367
R369 B.n295 B.n294 163.367
R370 B.n296 B.n295 163.367
R371 B.n296 B.n47 163.367
R372 B.n300 B.n47 163.367
R373 B.n301 B.n300 163.367
R374 B.n302 B.n301 163.367
R375 B.n302 B.n45 163.367
R376 B.n306 B.n45 163.367
R377 B.n307 B.n306 163.367
R378 B.n308 B.n307 163.367
R379 B.n379 B.n378 163.367
R380 B.n378 B.n17 163.367
R381 B.n374 B.n17 163.367
R382 B.n374 B.n373 163.367
R383 B.n373 B.n372 163.367
R384 B.n372 B.n19 163.367
R385 B.n368 B.n19 163.367
R386 B.n368 B.n367 163.367
R387 B.n367 B.n366 163.367
R388 B.n366 B.n21 163.367
R389 B.n362 B.n21 163.367
R390 B.n362 B.n361 163.367
R391 B.n361 B.n360 163.367
R392 B.n360 B.n23 163.367
R393 B.n356 B.n23 163.367
R394 B.n356 B.n355 163.367
R395 B.n355 B.n354 163.367
R396 B.n354 B.n25 163.367
R397 B.n349 B.n25 163.367
R398 B.n349 B.n348 163.367
R399 B.n348 B.n347 163.367
R400 B.n347 B.n29 163.367
R401 B.n343 B.n29 163.367
R402 B.n343 B.n342 163.367
R403 B.n342 B.n341 163.367
R404 B.n341 B.n31 163.367
R405 B.n337 B.n31 163.367
R406 B.n337 B.n336 163.367
R407 B.n336 B.n35 163.367
R408 B.n332 B.n35 163.367
R409 B.n332 B.n331 163.367
R410 B.n331 B.n330 163.367
R411 B.n330 B.n37 163.367
R412 B.n326 B.n37 163.367
R413 B.n326 B.n325 163.367
R414 B.n325 B.n324 163.367
R415 B.n324 B.n39 163.367
R416 B.n320 B.n39 163.367
R417 B.n320 B.n319 163.367
R418 B.n319 B.n318 163.367
R419 B.n318 B.n41 163.367
R420 B.n314 B.n41 163.367
R421 B.n314 B.n313 163.367
R422 B.n313 B.n312 163.367
R423 B.n312 B.n43 163.367
R424 B.n83 B.n82 65.1641
R425 B.n89 B.n88 65.1641
R426 B.n27 B.n26 65.1641
R427 B.n33 B.n32 65.1641
R428 B.n196 B.n83 59.5399
R429 B.n90 B.n89 59.5399
R430 B.n352 B.n27 59.5399
R431 B.n34 B.n33 59.5399
R432 B.n310 B.n309 28.8785
R433 B.n381 B.n16 28.8785
R434 B.n225 B.n72 28.8785
R435 B.n154 B.n153 28.8785
R436 B B.n423 18.0485
R437 B.n377 B.n16 10.6151
R438 B.n377 B.n376 10.6151
R439 B.n376 B.n375 10.6151
R440 B.n375 B.n18 10.6151
R441 B.n371 B.n18 10.6151
R442 B.n371 B.n370 10.6151
R443 B.n370 B.n369 10.6151
R444 B.n369 B.n20 10.6151
R445 B.n365 B.n20 10.6151
R446 B.n365 B.n364 10.6151
R447 B.n364 B.n363 10.6151
R448 B.n363 B.n22 10.6151
R449 B.n359 B.n22 10.6151
R450 B.n359 B.n358 10.6151
R451 B.n358 B.n357 10.6151
R452 B.n357 B.n24 10.6151
R453 B.n353 B.n24 10.6151
R454 B.n351 B.n350 10.6151
R455 B.n350 B.n28 10.6151
R456 B.n346 B.n28 10.6151
R457 B.n346 B.n345 10.6151
R458 B.n345 B.n344 10.6151
R459 B.n344 B.n30 10.6151
R460 B.n340 B.n30 10.6151
R461 B.n340 B.n339 10.6151
R462 B.n339 B.n338 10.6151
R463 B.n335 B.n334 10.6151
R464 B.n334 B.n333 10.6151
R465 B.n333 B.n36 10.6151
R466 B.n329 B.n36 10.6151
R467 B.n329 B.n328 10.6151
R468 B.n328 B.n327 10.6151
R469 B.n327 B.n38 10.6151
R470 B.n323 B.n38 10.6151
R471 B.n323 B.n322 10.6151
R472 B.n322 B.n321 10.6151
R473 B.n321 B.n40 10.6151
R474 B.n317 B.n40 10.6151
R475 B.n317 B.n316 10.6151
R476 B.n316 B.n315 10.6151
R477 B.n315 B.n42 10.6151
R478 B.n311 B.n42 10.6151
R479 B.n311 B.n310 10.6151
R480 B.n226 B.n225 10.6151
R481 B.n227 B.n226 10.6151
R482 B.n227 B.n70 10.6151
R483 B.n231 B.n70 10.6151
R484 B.n232 B.n231 10.6151
R485 B.n233 B.n232 10.6151
R486 B.n233 B.n68 10.6151
R487 B.n237 B.n68 10.6151
R488 B.n238 B.n237 10.6151
R489 B.n239 B.n238 10.6151
R490 B.n239 B.n66 10.6151
R491 B.n243 B.n66 10.6151
R492 B.n244 B.n243 10.6151
R493 B.n245 B.n244 10.6151
R494 B.n245 B.n64 10.6151
R495 B.n249 B.n64 10.6151
R496 B.n250 B.n249 10.6151
R497 B.n251 B.n250 10.6151
R498 B.n251 B.n62 10.6151
R499 B.n255 B.n62 10.6151
R500 B.n256 B.n255 10.6151
R501 B.n257 B.n256 10.6151
R502 B.n257 B.n60 10.6151
R503 B.n261 B.n60 10.6151
R504 B.n262 B.n261 10.6151
R505 B.n263 B.n262 10.6151
R506 B.n263 B.n58 10.6151
R507 B.n267 B.n58 10.6151
R508 B.n268 B.n267 10.6151
R509 B.n269 B.n268 10.6151
R510 B.n269 B.n56 10.6151
R511 B.n273 B.n56 10.6151
R512 B.n274 B.n273 10.6151
R513 B.n275 B.n274 10.6151
R514 B.n275 B.n54 10.6151
R515 B.n279 B.n54 10.6151
R516 B.n280 B.n279 10.6151
R517 B.n281 B.n280 10.6151
R518 B.n281 B.n52 10.6151
R519 B.n285 B.n52 10.6151
R520 B.n286 B.n285 10.6151
R521 B.n287 B.n286 10.6151
R522 B.n287 B.n50 10.6151
R523 B.n291 B.n50 10.6151
R524 B.n292 B.n291 10.6151
R525 B.n293 B.n292 10.6151
R526 B.n293 B.n48 10.6151
R527 B.n297 B.n48 10.6151
R528 B.n298 B.n297 10.6151
R529 B.n299 B.n298 10.6151
R530 B.n299 B.n46 10.6151
R531 B.n303 B.n46 10.6151
R532 B.n304 B.n303 10.6151
R533 B.n305 B.n304 10.6151
R534 B.n305 B.n44 10.6151
R535 B.n309 B.n44 10.6151
R536 B.n155 B.n154 10.6151
R537 B.n155 B.n98 10.6151
R538 B.n159 B.n98 10.6151
R539 B.n160 B.n159 10.6151
R540 B.n161 B.n160 10.6151
R541 B.n161 B.n96 10.6151
R542 B.n165 B.n96 10.6151
R543 B.n166 B.n165 10.6151
R544 B.n167 B.n166 10.6151
R545 B.n167 B.n94 10.6151
R546 B.n171 B.n94 10.6151
R547 B.n172 B.n171 10.6151
R548 B.n173 B.n172 10.6151
R549 B.n173 B.n92 10.6151
R550 B.n177 B.n92 10.6151
R551 B.n178 B.n177 10.6151
R552 B.n179 B.n178 10.6151
R553 B.n183 B.n182 10.6151
R554 B.n184 B.n183 10.6151
R555 B.n184 B.n86 10.6151
R556 B.n188 B.n86 10.6151
R557 B.n189 B.n188 10.6151
R558 B.n190 B.n189 10.6151
R559 B.n190 B.n84 10.6151
R560 B.n194 B.n84 10.6151
R561 B.n195 B.n194 10.6151
R562 B.n197 B.n80 10.6151
R563 B.n201 B.n80 10.6151
R564 B.n202 B.n201 10.6151
R565 B.n203 B.n202 10.6151
R566 B.n203 B.n78 10.6151
R567 B.n207 B.n78 10.6151
R568 B.n208 B.n207 10.6151
R569 B.n209 B.n208 10.6151
R570 B.n209 B.n76 10.6151
R571 B.n213 B.n76 10.6151
R572 B.n214 B.n213 10.6151
R573 B.n215 B.n214 10.6151
R574 B.n215 B.n74 10.6151
R575 B.n219 B.n74 10.6151
R576 B.n220 B.n219 10.6151
R577 B.n221 B.n220 10.6151
R578 B.n221 B.n72 10.6151
R579 B.n153 B.n100 10.6151
R580 B.n149 B.n100 10.6151
R581 B.n149 B.n148 10.6151
R582 B.n148 B.n147 10.6151
R583 B.n147 B.n102 10.6151
R584 B.n143 B.n102 10.6151
R585 B.n143 B.n142 10.6151
R586 B.n142 B.n141 10.6151
R587 B.n141 B.n104 10.6151
R588 B.n137 B.n104 10.6151
R589 B.n137 B.n136 10.6151
R590 B.n136 B.n135 10.6151
R591 B.n135 B.n106 10.6151
R592 B.n131 B.n106 10.6151
R593 B.n131 B.n130 10.6151
R594 B.n130 B.n129 10.6151
R595 B.n129 B.n108 10.6151
R596 B.n125 B.n108 10.6151
R597 B.n125 B.n124 10.6151
R598 B.n124 B.n123 10.6151
R599 B.n123 B.n110 10.6151
R600 B.n119 B.n110 10.6151
R601 B.n119 B.n118 10.6151
R602 B.n118 B.n117 10.6151
R603 B.n117 B.n112 10.6151
R604 B.n113 B.n112 10.6151
R605 B.n113 B.n0 10.6151
R606 B.n419 B.n1 10.6151
R607 B.n419 B.n418 10.6151
R608 B.n418 B.n417 10.6151
R609 B.n417 B.n4 10.6151
R610 B.n413 B.n4 10.6151
R611 B.n413 B.n412 10.6151
R612 B.n412 B.n411 10.6151
R613 B.n411 B.n6 10.6151
R614 B.n407 B.n6 10.6151
R615 B.n407 B.n406 10.6151
R616 B.n406 B.n405 10.6151
R617 B.n405 B.n8 10.6151
R618 B.n401 B.n8 10.6151
R619 B.n401 B.n400 10.6151
R620 B.n400 B.n399 10.6151
R621 B.n399 B.n10 10.6151
R622 B.n395 B.n10 10.6151
R623 B.n395 B.n394 10.6151
R624 B.n394 B.n393 10.6151
R625 B.n393 B.n12 10.6151
R626 B.n389 B.n12 10.6151
R627 B.n389 B.n388 10.6151
R628 B.n388 B.n387 10.6151
R629 B.n387 B.n14 10.6151
R630 B.n383 B.n14 10.6151
R631 B.n383 B.n382 10.6151
R632 B.n382 B.n381 10.6151
R633 B.n353 B.n352 9.52245
R634 B.n335 B.n34 9.52245
R635 B.n179 B.n90 9.52245
R636 B.n197 B.n196 9.52245
R637 B.n423 B.n0 2.81026
R638 B.n423 B.n1 2.81026
R639 B.n352 B.n351 1.09318
R640 B.n338 B.n34 1.09318
R641 B.n182 B.n90 1.09318
R642 B.n196 B.n195 1.09318
R643 VN VN.t0 112.388
R644 VN VN.t1 73.1041
R645 VTAIL.n74 VTAIL.n60 756.745
R646 VTAIL.n14 VTAIL.n0 756.745
R647 VTAIL.n54 VTAIL.n40 756.745
R648 VTAIL.n34 VTAIL.n20 756.745
R649 VTAIL.n67 VTAIL.n66 585
R650 VTAIL.n64 VTAIL.n63 585
R651 VTAIL.n73 VTAIL.n72 585
R652 VTAIL.n75 VTAIL.n74 585
R653 VTAIL.n7 VTAIL.n6 585
R654 VTAIL.n4 VTAIL.n3 585
R655 VTAIL.n13 VTAIL.n12 585
R656 VTAIL.n15 VTAIL.n14 585
R657 VTAIL.n55 VTAIL.n54 585
R658 VTAIL.n53 VTAIL.n52 585
R659 VTAIL.n44 VTAIL.n43 585
R660 VTAIL.n47 VTAIL.n46 585
R661 VTAIL.n35 VTAIL.n34 585
R662 VTAIL.n33 VTAIL.n32 585
R663 VTAIL.n24 VTAIL.n23 585
R664 VTAIL.n27 VTAIL.n26 585
R665 VTAIL.t2 VTAIL.n65 330.707
R666 VTAIL.t0 VTAIL.n5 330.707
R667 VTAIL.t1 VTAIL.n45 330.707
R668 VTAIL.t3 VTAIL.n25 330.707
R669 VTAIL.n66 VTAIL.n63 171.744
R670 VTAIL.n73 VTAIL.n63 171.744
R671 VTAIL.n74 VTAIL.n73 171.744
R672 VTAIL.n6 VTAIL.n3 171.744
R673 VTAIL.n13 VTAIL.n3 171.744
R674 VTAIL.n14 VTAIL.n13 171.744
R675 VTAIL.n54 VTAIL.n53 171.744
R676 VTAIL.n53 VTAIL.n43 171.744
R677 VTAIL.n46 VTAIL.n43 171.744
R678 VTAIL.n34 VTAIL.n33 171.744
R679 VTAIL.n33 VTAIL.n23 171.744
R680 VTAIL.n26 VTAIL.n23 171.744
R681 VTAIL.n66 VTAIL.t2 85.8723
R682 VTAIL.n6 VTAIL.t0 85.8723
R683 VTAIL.n46 VTAIL.t1 85.8723
R684 VTAIL.n26 VTAIL.t3 85.8723
R685 VTAIL.n79 VTAIL.n78 34.7066
R686 VTAIL.n19 VTAIL.n18 34.7066
R687 VTAIL.n59 VTAIL.n58 34.7066
R688 VTAIL.n39 VTAIL.n38 34.7066
R689 VTAIL.n39 VTAIL.n19 21.5824
R690 VTAIL.n79 VTAIL.n59 18.6858
R691 VTAIL.n67 VTAIL.n65 16.3201
R692 VTAIL.n7 VTAIL.n5 16.3201
R693 VTAIL.n47 VTAIL.n45 16.3201
R694 VTAIL.n27 VTAIL.n25 16.3201
R695 VTAIL.n68 VTAIL.n64 12.8005
R696 VTAIL.n8 VTAIL.n4 12.8005
R697 VTAIL.n48 VTAIL.n44 12.8005
R698 VTAIL.n28 VTAIL.n24 12.8005
R699 VTAIL.n72 VTAIL.n71 12.0247
R700 VTAIL.n12 VTAIL.n11 12.0247
R701 VTAIL.n52 VTAIL.n51 12.0247
R702 VTAIL.n32 VTAIL.n31 12.0247
R703 VTAIL.n75 VTAIL.n62 11.249
R704 VTAIL.n15 VTAIL.n2 11.249
R705 VTAIL.n55 VTAIL.n42 11.249
R706 VTAIL.n35 VTAIL.n22 11.249
R707 VTAIL.n76 VTAIL.n60 10.4732
R708 VTAIL.n16 VTAIL.n0 10.4732
R709 VTAIL.n56 VTAIL.n40 10.4732
R710 VTAIL.n36 VTAIL.n20 10.4732
R711 VTAIL.n78 VTAIL.n77 9.45567
R712 VTAIL.n18 VTAIL.n17 9.45567
R713 VTAIL.n58 VTAIL.n57 9.45567
R714 VTAIL.n38 VTAIL.n37 9.45567
R715 VTAIL.n77 VTAIL.n76 9.3005
R716 VTAIL.n62 VTAIL.n61 9.3005
R717 VTAIL.n71 VTAIL.n70 9.3005
R718 VTAIL.n69 VTAIL.n68 9.3005
R719 VTAIL.n17 VTAIL.n16 9.3005
R720 VTAIL.n2 VTAIL.n1 9.3005
R721 VTAIL.n11 VTAIL.n10 9.3005
R722 VTAIL.n9 VTAIL.n8 9.3005
R723 VTAIL.n57 VTAIL.n56 9.3005
R724 VTAIL.n42 VTAIL.n41 9.3005
R725 VTAIL.n51 VTAIL.n50 9.3005
R726 VTAIL.n49 VTAIL.n48 9.3005
R727 VTAIL.n37 VTAIL.n36 9.3005
R728 VTAIL.n22 VTAIL.n21 9.3005
R729 VTAIL.n31 VTAIL.n30 9.3005
R730 VTAIL.n29 VTAIL.n28 9.3005
R731 VTAIL.n69 VTAIL.n65 3.78097
R732 VTAIL.n9 VTAIL.n5 3.78097
R733 VTAIL.n49 VTAIL.n45 3.78097
R734 VTAIL.n29 VTAIL.n25 3.78097
R735 VTAIL.n78 VTAIL.n60 3.49141
R736 VTAIL.n18 VTAIL.n0 3.49141
R737 VTAIL.n58 VTAIL.n40 3.49141
R738 VTAIL.n38 VTAIL.n20 3.49141
R739 VTAIL.n76 VTAIL.n75 2.71565
R740 VTAIL.n16 VTAIL.n15 2.71565
R741 VTAIL.n56 VTAIL.n55 2.71565
R742 VTAIL.n36 VTAIL.n35 2.71565
R743 VTAIL.n72 VTAIL.n62 1.93989
R744 VTAIL.n12 VTAIL.n2 1.93989
R745 VTAIL.n52 VTAIL.n42 1.93989
R746 VTAIL.n32 VTAIL.n22 1.93989
R747 VTAIL.n59 VTAIL.n39 1.9186
R748 VTAIL VTAIL.n19 1.25266
R749 VTAIL.n71 VTAIL.n64 1.16414
R750 VTAIL.n11 VTAIL.n4 1.16414
R751 VTAIL.n51 VTAIL.n44 1.16414
R752 VTAIL.n31 VTAIL.n24 1.16414
R753 VTAIL VTAIL.n79 0.666448
R754 VTAIL.n68 VTAIL.n67 0.388379
R755 VTAIL.n8 VTAIL.n7 0.388379
R756 VTAIL.n48 VTAIL.n47 0.388379
R757 VTAIL.n28 VTAIL.n27 0.388379
R758 VTAIL.n70 VTAIL.n69 0.155672
R759 VTAIL.n70 VTAIL.n61 0.155672
R760 VTAIL.n77 VTAIL.n61 0.155672
R761 VTAIL.n10 VTAIL.n9 0.155672
R762 VTAIL.n10 VTAIL.n1 0.155672
R763 VTAIL.n17 VTAIL.n1 0.155672
R764 VTAIL.n57 VTAIL.n41 0.155672
R765 VTAIL.n50 VTAIL.n41 0.155672
R766 VTAIL.n50 VTAIL.n49 0.155672
R767 VTAIL.n37 VTAIL.n21 0.155672
R768 VTAIL.n30 VTAIL.n21 0.155672
R769 VTAIL.n30 VTAIL.n29 0.155672
R770 VDD2.n33 VDD2.n19 756.745
R771 VDD2.n14 VDD2.n0 756.745
R772 VDD2.n34 VDD2.n33 585
R773 VDD2.n32 VDD2.n31 585
R774 VDD2.n23 VDD2.n22 585
R775 VDD2.n26 VDD2.n25 585
R776 VDD2.n7 VDD2.n6 585
R777 VDD2.n4 VDD2.n3 585
R778 VDD2.n13 VDD2.n12 585
R779 VDD2.n15 VDD2.n14 585
R780 VDD2.t1 VDD2.n24 330.707
R781 VDD2.t0 VDD2.n5 330.707
R782 VDD2.n33 VDD2.n32 171.744
R783 VDD2.n32 VDD2.n22 171.744
R784 VDD2.n25 VDD2.n22 171.744
R785 VDD2.n6 VDD2.n3 171.744
R786 VDD2.n13 VDD2.n3 171.744
R787 VDD2.n14 VDD2.n13 171.744
R788 VDD2.n25 VDD2.t1 85.8723
R789 VDD2.n6 VDD2.t0 85.8723
R790 VDD2.n38 VDD2.n18 84.2603
R791 VDD2.n38 VDD2.n37 51.3853
R792 VDD2.n26 VDD2.n24 16.3201
R793 VDD2.n7 VDD2.n5 16.3201
R794 VDD2.n27 VDD2.n23 12.8005
R795 VDD2.n8 VDD2.n4 12.8005
R796 VDD2.n31 VDD2.n30 12.0247
R797 VDD2.n12 VDD2.n11 12.0247
R798 VDD2.n34 VDD2.n21 11.249
R799 VDD2.n15 VDD2.n2 11.249
R800 VDD2.n35 VDD2.n19 10.4732
R801 VDD2.n16 VDD2.n0 10.4732
R802 VDD2.n37 VDD2.n36 9.45567
R803 VDD2.n18 VDD2.n17 9.45567
R804 VDD2.n36 VDD2.n35 9.3005
R805 VDD2.n21 VDD2.n20 9.3005
R806 VDD2.n30 VDD2.n29 9.3005
R807 VDD2.n28 VDD2.n27 9.3005
R808 VDD2.n17 VDD2.n16 9.3005
R809 VDD2.n2 VDD2.n1 9.3005
R810 VDD2.n11 VDD2.n10 9.3005
R811 VDD2.n9 VDD2.n8 9.3005
R812 VDD2.n28 VDD2.n24 3.78097
R813 VDD2.n9 VDD2.n5 3.78097
R814 VDD2.n37 VDD2.n19 3.49141
R815 VDD2.n18 VDD2.n0 3.49141
R816 VDD2.n35 VDD2.n34 2.71565
R817 VDD2.n16 VDD2.n15 2.71565
R818 VDD2.n31 VDD2.n21 1.93989
R819 VDD2.n12 VDD2.n2 1.93989
R820 VDD2.n30 VDD2.n23 1.16414
R821 VDD2.n11 VDD2.n4 1.16414
R822 VDD2 VDD2.n38 0.782828
R823 VDD2.n27 VDD2.n26 0.388379
R824 VDD2.n8 VDD2.n7 0.388379
R825 VDD2.n36 VDD2.n20 0.155672
R826 VDD2.n29 VDD2.n20 0.155672
R827 VDD2.n29 VDD2.n28 0.155672
R828 VDD2.n10 VDD2.n9 0.155672
R829 VDD2.n10 VDD2.n1 0.155672
R830 VDD2.n17 VDD2.n1 0.155672
R831 VP.n0 VP.t1 112.386
R832 VP.n0 VP.t0 72.6728
R833 VP VP.n0 0.431811
R834 VDD1.n14 VDD1.n0 756.745
R835 VDD1.n33 VDD1.n19 756.745
R836 VDD1.n15 VDD1.n14 585
R837 VDD1.n13 VDD1.n12 585
R838 VDD1.n4 VDD1.n3 585
R839 VDD1.n7 VDD1.n6 585
R840 VDD1.n26 VDD1.n25 585
R841 VDD1.n23 VDD1.n22 585
R842 VDD1.n32 VDD1.n31 585
R843 VDD1.n34 VDD1.n33 585
R844 VDD1.t0 VDD1.n5 330.707
R845 VDD1.t1 VDD1.n24 330.707
R846 VDD1.n14 VDD1.n13 171.744
R847 VDD1.n13 VDD1.n3 171.744
R848 VDD1.n6 VDD1.n3 171.744
R849 VDD1.n25 VDD1.n22 171.744
R850 VDD1.n32 VDD1.n22 171.744
R851 VDD1.n33 VDD1.n32 171.744
R852 VDD1.n6 VDD1.t0 85.8723
R853 VDD1.n25 VDD1.t1 85.8723
R854 VDD1 VDD1.n37 85.5093
R855 VDD1 VDD1.n18 52.1677
R856 VDD1.n7 VDD1.n5 16.3201
R857 VDD1.n26 VDD1.n24 16.3201
R858 VDD1.n8 VDD1.n4 12.8005
R859 VDD1.n27 VDD1.n23 12.8005
R860 VDD1.n12 VDD1.n11 12.0247
R861 VDD1.n31 VDD1.n30 12.0247
R862 VDD1.n15 VDD1.n2 11.249
R863 VDD1.n34 VDD1.n21 11.249
R864 VDD1.n16 VDD1.n0 10.4732
R865 VDD1.n35 VDD1.n19 10.4732
R866 VDD1.n18 VDD1.n17 9.45567
R867 VDD1.n37 VDD1.n36 9.45567
R868 VDD1.n17 VDD1.n16 9.3005
R869 VDD1.n2 VDD1.n1 9.3005
R870 VDD1.n11 VDD1.n10 9.3005
R871 VDD1.n9 VDD1.n8 9.3005
R872 VDD1.n36 VDD1.n35 9.3005
R873 VDD1.n21 VDD1.n20 9.3005
R874 VDD1.n30 VDD1.n29 9.3005
R875 VDD1.n28 VDD1.n27 9.3005
R876 VDD1.n9 VDD1.n5 3.78097
R877 VDD1.n28 VDD1.n24 3.78097
R878 VDD1.n18 VDD1.n0 3.49141
R879 VDD1.n37 VDD1.n19 3.49141
R880 VDD1.n16 VDD1.n15 2.71565
R881 VDD1.n35 VDD1.n34 2.71565
R882 VDD1.n12 VDD1.n2 1.93989
R883 VDD1.n31 VDD1.n21 1.93989
R884 VDD1.n11 VDD1.n4 1.16414
R885 VDD1.n30 VDD1.n23 1.16414
R886 VDD1.n8 VDD1.n7 0.388379
R887 VDD1.n27 VDD1.n26 0.388379
R888 VDD1.n17 VDD1.n1 0.155672
R889 VDD1.n10 VDD1.n1 0.155672
R890 VDD1.n10 VDD1.n9 0.155672
R891 VDD1.n29 VDD1.n28 0.155672
R892 VDD1.n29 VDD1.n20 0.155672
R893 VDD1.n36 VDD1.n20 0.155672
C0 VTAIL VP 1.31834f
C1 VTAIL w_n2314_n1762# 1.6221f
C2 B VDD2 1.15672f
C3 VP VN 4.1741f
C4 VTAIL B 1.93548f
C5 w_n2314_n1762# VN 3.07945f
C6 VDD1 VDD2 0.726006f
C7 w_n2314_n1762# VP 3.37421f
C8 VDD1 VTAIL 3.07103f
C9 B VN 1.02345f
C10 B VP 1.5111f
C11 B w_n2314_n1762# 7.05573f
C12 VDD1 VN 0.152593f
C13 VDD1 VP 1.31436f
C14 VDD1 w_n2314_n1762# 1.27356f
C15 VTAIL VDD2 3.12654f
C16 VDD1 B 1.12264f
C17 VDD2 VN 1.11325f
C18 VDD2 VP 0.355225f
C19 VTAIL VN 1.30418f
C20 VDD2 w_n2314_n1762# 1.30437f
C21 VDD2 VSUBS 0.633964f
C22 VDD1 VSUBS 2.377773f
C23 VTAIL VSUBS 0.448204f
C24 VN VSUBS 5.53934f
C25 VP VSUBS 1.377228f
C26 B VSUBS 3.36481f
C27 w_n2314_n1762# VSUBS 51.343f
C28 VDD1.n0 VSUBS 0.017125f
C29 VDD1.n1 VSUBS 0.015584f
C30 VDD1.n2 VSUBS 0.008374f
C31 VDD1.n3 VSUBS 0.019794f
C32 VDD1.n4 VSUBS 0.008867f
C33 VDD1.n5 VSUBS 0.060616f
C34 VDD1.t0 VSUBS 0.043879f
C35 VDD1.n6 VSUBS 0.014845f
C36 VDD1.n7 VSUBS 0.01245f
C37 VDD1.n8 VSUBS 0.008374f
C38 VDD1.n9 VSUBS 0.211478f
C39 VDD1.n10 VSUBS 0.015584f
C40 VDD1.n11 VSUBS 0.008374f
C41 VDD1.n12 VSUBS 0.008867f
C42 VDD1.n13 VSUBS 0.019794f
C43 VDD1.n14 VSUBS 0.047921f
C44 VDD1.n15 VSUBS 0.008867f
C45 VDD1.n16 VSUBS 0.008374f
C46 VDD1.n17 VSUBS 0.03879f
C47 VDD1.n18 VSUBS 0.035985f
C48 VDD1.n19 VSUBS 0.017125f
C49 VDD1.n20 VSUBS 0.015584f
C50 VDD1.n21 VSUBS 0.008374f
C51 VDD1.n22 VSUBS 0.019794f
C52 VDD1.n23 VSUBS 0.008867f
C53 VDD1.n24 VSUBS 0.060616f
C54 VDD1.t1 VSUBS 0.043879f
C55 VDD1.n25 VSUBS 0.014845f
C56 VDD1.n26 VSUBS 0.01245f
C57 VDD1.n27 VSUBS 0.008374f
C58 VDD1.n28 VSUBS 0.211478f
C59 VDD1.n29 VSUBS 0.015584f
C60 VDD1.n30 VSUBS 0.008374f
C61 VDD1.n31 VSUBS 0.008867f
C62 VDD1.n32 VSUBS 0.019794f
C63 VDD1.n33 VSUBS 0.047921f
C64 VDD1.n34 VSUBS 0.008867f
C65 VDD1.n35 VSUBS 0.008374f
C66 VDD1.n36 VSUBS 0.03879f
C67 VDD1.n37 VSUBS 0.330106f
C68 VP.t0 VSUBS 1.69246f
C69 VP.t1 VSUBS 2.43077f
C70 VP.n0 VSUBS 3.35546f
C71 VDD2.n0 VSUBS 0.017448f
C72 VDD2.n1 VSUBS 0.015879f
C73 VDD2.n2 VSUBS 0.008533f
C74 VDD2.n3 VSUBS 0.020168f
C75 VDD2.n4 VSUBS 0.009035f
C76 VDD2.n5 VSUBS 0.061763f
C77 VDD2.t0 VSUBS 0.044709f
C78 VDD2.n6 VSUBS 0.015126f
C79 VDD2.n7 VSUBS 0.012685f
C80 VDD2.n8 VSUBS 0.008533f
C81 VDD2.n9 VSUBS 0.215479f
C82 VDD2.n10 VSUBS 0.015879f
C83 VDD2.n11 VSUBS 0.008533f
C84 VDD2.n12 VSUBS 0.009035f
C85 VDD2.n13 VSUBS 0.020168f
C86 VDD2.n14 VSUBS 0.048828f
C87 VDD2.n15 VSUBS 0.009035f
C88 VDD2.n16 VSUBS 0.008533f
C89 VDD2.n17 VSUBS 0.039523f
C90 VDD2.n18 VSUBS 0.308687f
C91 VDD2.n19 VSUBS 0.017448f
C92 VDD2.n20 VSUBS 0.015879f
C93 VDD2.n21 VSUBS 0.008533f
C94 VDD2.n22 VSUBS 0.020168f
C95 VDD2.n23 VSUBS 0.009035f
C96 VDD2.n24 VSUBS 0.061763f
C97 VDD2.t1 VSUBS 0.044709f
C98 VDD2.n25 VSUBS 0.015126f
C99 VDD2.n26 VSUBS 0.012685f
C100 VDD2.n27 VSUBS 0.008533f
C101 VDD2.n28 VSUBS 0.215479f
C102 VDD2.n29 VSUBS 0.015879f
C103 VDD2.n30 VSUBS 0.008533f
C104 VDD2.n31 VSUBS 0.009035f
C105 VDD2.n32 VSUBS 0.020168f
C106 VDD2.n33 VSUBS 0.048828f
C107 VDD2.n34 VSUBS 0.009035f
C108 VDD2.n35 VSUBS 0.008533f
C109 VDD2.n36 VSUBS 0.039523f
C110 VDD2.n37 VSUBS 0.035583f
C111 VDD2.n38 VSUBS 1.46338f
C112 VTAIL.n0 VSUBS 0.020184f
C113 VTAIL.n1 VSUBS 0.018368f
C114 VTAIL.n2 VSUBS 0.00987f
C115 VTAIL.n3 VSUBS 0.02333f
C116 VTAIL.n4 VSUBS 0.010451f
C117 VTAIL.n5 VSUBS 0.071446f
C118 VTAIL.t0 VSUBS 0.051718f
C119 VTAIL.n6 VSUBS 0.017497f
C120 VTAIL.n7 VSUBS 0.014674f
C121 VTAIL.n8 VSUBS 0.00987f
C122 VTAIL.n9 VSUBS 0.249259f
C123 VTAIL.n10 VSUBS 0.018368f
C124 VTAIL.n11 VSUBS 0.00987f
C125 VTAIL.n12 VSUBS 0.010451f
C126 VTAIL.n13 VSUBS 0.02333f
C127 VTAIL.n14 VSUBS 0.056483f
C128 VTAIL.n15 VSUBS 0.010451f
C129 VTAIL.n16 VSUBS 0.00987f
C130 VTAIL.n17 VSUBS 0.04572f
C131 VTAIL.n18 VSUBS 0.028502f
C132 VTAIL.n19 VSUBS 0.886591f
C133 VTAIL.n20 VSUBS 0.020184f
C134 VTAIL.n21 VSUBS 0.018368f
C135 VTAIL.n22 VSUBS 0.00987f
C136 VTAIL.n23 VSUBS 0.02333f
C137 VTAIL.n24 VSUBS 0.010451f
C138 VTAIL.n25 VSUBS 0.071446f
C139 VTAIL.t3 VSUBS 0.051718f
C140 VTAIL.n26 VSUBS 0.017497f
C141 VTAIL.n27 VSUBS 0.014674f
C142 VTAIL.n28 VSUBS 0.00987f
C143 VTAIL.n29 VSUBS 0.249259f
C144 VTAIL.n30 VSUBS 0.018368f
C145 VTAIL.n31 VSUBS 0.00987f
C146 VTAIL.n32 VSUBS 0.010451f
C147 VTAIL.n33 VSUBS 0.02333f
C148 VTAIL.n34 VSUBS 0.056483f
C149 VTAIL.n35 VSUBS 0.010451f
C150 VTAIL.n36 VSUBS 0.00987f
C151 VTAIL.n37 VSUBS 0.04572f
C152 VTAIL.n38 VSUBS 0.028502f
C153 VTAIL.n39 VSUBS 0.926006f
C154 VTAIL.n40 VSUBS 0.020184f
C155 VTAIL.n41 VSUBS 0.018368f
C156 VTAIL.n42 VSUBS 0.00987f
C157 VTAIL.n43 VSUBS 0.02333f
C158 VTAIL.n44 VSUBS 0.010451f
C159 VTAIL.n45 VSUBS 0.071446f
C160 VTAIL.t1 VSUBS 0.051718f
C161 VTAIL.n46 VSUBS 0.017497f
C162 VTAIL.n47 VSUBS 0.014674f
C163 VTAIL.n48 VSUBS 0.00987f
C164 VTAIL.n49 VSUBS 0.249259f
C165 VTAIL.n50 VSUBS 0.018368f
C166 VTAIL.n51 VSUBS 0.00987f
C167 VTAIL.n52 VSUBS 0.010451f
C168 VTAIL.n53 VSUBS 0.02333f
C169 VTAIL.n54 VSUBS 0.056483f
C170 VTAIL.n55 VSUBS 0.010451f
C171 VTAIL.n56 VSUBS 0.00987f
C172 VTAIL.n57 VSUBS 0.04572f
C173 VTAIL.n58 VSUBS 0.028502f
C174 VTAIL.n59 VSUBS 0.754569f
C175 VTAIL.n60 VSUBS 0.020184f
C176 VTAIL.n61 VSUBS 0.018368f
C177 VTAIL.n62 VSUBS 0.00987f
C178 VTAIL.n63 VSUBS 0.02333f
C179 VTAIL.n64 VSUBS 0.010451f
C180 VTAIL.n65 VSUBS 0.071446f
C181 VTAIL.t2 VSUBS 0.051718f
C182 VTAIL.n66 VSUBS 0.017497f
C183 VTAIL.n67 VSUBS 0.014674f
C184 VTAIL.n68 VSUBS 0.00987f
C185 VTAIL.n69 VSUBS 0.249259f
C186 VTAIL.n70 VSUBS 0.018368f
C187 VTAIL.n71 VSUBS 0.00987f
C188 VTAIL.n72 VSUBS 0.010451f
C189 VTAIL.n73 VSUBS 0.02333f
C190 VTAIL.n74 VSUBS 0.056483f
C191 VTAIL.n75 VSUBS 0.010451f
C192 VTAIL.n76 VSUBS 0.00987f
C193 VTAIL.n77 VSUBS 0.04572f
C194 VTAIL.n78 VSUBS 0.028502f
C195 VTAIL.n79 VSUBS 0.680458f
C196 VN.t1 VSUBS 1.61679f
C197 VN.t0 VSUBS 2.32134f
C198 B.n0 VSUBS 0.004501f
C199 B.n1 VSUBS 0.004501f
C200 B.n2 VSUBS 0.007118f
C201 B.n3 VSUBS 0.007118f
C202 B.n4 VSUBS 0.007118f
C203 B.n5 VSUBS 0.007118f
C204 B.n6 VSUBS 0.007118f
C205 B.n7 VSUBS 0.007118f
C206 B.n8 VSUBS 0.007118f
C207 B.n9 VSUBS 0.007118f
C208 B.n10 VSUBS 0.007118f
C209 B.n11 VSUBS 0.007118f
C210 B.n12 VSUBS 0.007118f
C211 B.n13 VSUBS 0.007118f
C212 B.n14 VSUBS 0.007118f
C213 B.n15 VSUBS 0.007118f
C214 B.n16 VSUBS 0.01591f
C215 B.n17 VSUBS 0.007118f
C216 B.n18 VSUBS 0.007118f
C217 B.n19 VSUBS 0.007118f
C218 B.n20 VSUBS 0.007118f
C219 B.n21 VSUBS 0.007118f
C220 B.n22 VSUBS 0.007118f
C221 B.n23 VSUBS 0.007118f
C222 B.n24 VSUBS 0.007118f
C223 B.n25 VSUBS 0.007118f
C224 B.t11 VSUBS 0.058608f
C225 B.t10 VSUBS 0.082161f
C226 B.t9 VSUBS 0.591742f
C227 B.n26 VSUBS 0.141388f
C228 B.n27 VSUBS 0.118733f
C229 B.n28 VSUBS 0.007118f
C230 B.n29 VSUBS 0.007118f
C231 B.n30 VSUBS 0.007118f
C232 B.n31 VSUBS 0.007118f
C233 B.t2 VSUBS 0.058609f
C234 B.t1 VSUBS 0.082162f
C235 B.t0 VSUBS 0.591782f
C236 B.n32 VSUBS 0.141347f
C237 B.n33 VSUBS 0.118732f
C238 B.n34 VSUBS 0.016492f
C239 B.n35 VSUBS 0.007118f
C240 B.n36 VSUBS 0.007118f
C241 B.n37 VSUBS 0.007118f
C242 B.n38 VSUBS 0.007118f
C243 B.n39 VSUBS 0.007118f
C244 B.n40 VSUBS 0.007118f
C245 B.n41 VSUBS 0.007118f
C246 B.n42 VSUBS 0.007118f
C247 B.n43 VSUBS 0.01591f
C248 B.n44 VSUBS 0.007118f
C249 B.n45 VSUBS 0.007118f
C250 B.n46 VSUBS 0.007118f
C251 B.n47 VSUBS 0.007118f
C252 B.n48 VSUBS 0.007118f
C253 B.n49 VSUBS 0.007118f
C254 B.n50 VSUBS 0.007118f
C255 B.n51 VSUBS 0.007118f
C256 B.n52 VSUBS 0.007118f
C257 B.n53 VSUBS 0.007118f
C258 B.n54 VSUBS 0.007118f
C259 B.n55 VSUBS 0.007118f
C260 B.n56 VSUBS 0.007118f
C261 B.n57 VSUBS 0.007118f
C262 B.n58 VSUBS 0.007118f
C263 B.n59 VSUBS 0.007118f
C264 B.n60 VSUBS 0.007118f
C265 B.n61 VSUBS 0.007118f
C266 B.n62 VSUBS 0.007118f
C267 B.n63 VSUBS 0.007118f
C268 B.n64 VSUBS 0.007118f
C269 B.n65 VSUBS 0.007118f
C270 B.n66 VSUBS 0.007118f
C271 B.n67 VSUBS 0.007118f
C272 B.n68 VSUBS 0.007118f
C273 B.n69 VSUBS 0.007118f
C274 B.n70 VSUBS 0.007118f
C275 B.n71 VSUBS 0.007118f
C276 B.n72 VSUBS 0.01591f
C277 B.n73 VSUBS 0.007118f
C278 B.n74 VSUBS 0.007118f
C279 B.n75 VSUBS 0.007118f
C280 B.n76 VSUBS 0.007118f
C281 B.n77 VSUBS 0.007118f
C282 B.n78 VSUBS 0.007118f
C283 B.n79 VSUBS 0.007118f
C284 B.n80 VSUBS 0.007118f
C285 B.n81 VSUBS 0.007118f
C286 B.t4 VSUBS 0.058609f
C287 B.t5 VSUBS 0.082162f
C288 B.t3 VSUBS 0.591782f
C289 B.n82 VSUBS 0.141347f
C290 B.n83 VSUBS 0.118732f
C291 B.n84 VSUBS 0.007118f
C292 B.n85 VSUBS 0.007118f
C293 B.n86 VSUBS 0.007118f
C294 B.n87 VSUBS 0.007118f
C295 B.t7 VSUBS 0.058608f
C296 B.t8 VSUBS 0.082161f
C297 B.t6 VSUBS 0.591742f
C298 B.n88 VSUBS 0.141388f
C299 B.n89 VSUBS 0.118733f
C300 B.n90 VSUBS 0.016492f
C301 B.n91 VSUBS 0.007118f
C302 B.n92 VSUBS 0.007118f
C303 B.n93 VSUBS 0.007118f
C304 B.n94 VSUBS 0.007118f
C305 B.n95 VSUBS 0.007118f
C306 B.n96 VSUBS 0.007118f
C307 B.n97 VSUBS 0.007118f
C308 B.n98 VSUBS 0.007118f
C309 B.n99 VSUBS 0.01591f
C310 B.n100 VSUBS 0.007118f
C311 B.n101 VSUBS 0.007118f
C312 B.n102 VSUBS 0.007118f
C313 B.n103 VSUBS 0.007118f
C314 B.n104 VSUBS 0.007118f
C315 B.n105 VSUBS 0.007118f
C316 B.n106 VSUBS 0.007118f
C317 B.n107 VSUBS 0.007118f
C318 B.n108 VSUBS 0.007118f
C319 B.n109 VSUBS 0.007118f
C320 B.n110 VSUBS 0.007118f
C321 B.n111 VSUBS 0.007118f
C322 B.n112 VSUBS 0.007118f
C323 B.n113 VSUBS 0.007118f
C324 B.n114 VSUBS 0.007118f
C325 B.n115 VSUBS 0.007118f
C326 B.n116 VSUBS 0.007118f
C327 B.n117 VSUBS 0.007118f
C328 B.n118 VSUBS 0.007118f
C329 B.n119 VSUBS 0.007118f
C330 B.n120 VSUBS 0.007118f
C331 B.n121 VSUBS 0.007118f
C332 B.n122 VSUBS 0.007118f
C333 B.n123 VSUBS 0.007118f
C334 B.n124 VSUBS 0.007118f
C335 B.n125 VSUBS 0.007118f
C336 B.n126 VSUBS 0.007118f
C337 B.n127 VSUBS 0.007118f
C338 B.n128 VSUBS 0.007118f
C339 B.n129 VSUBS 0.007118f
C340 B.n130 VSUBS 0.007118f
C341 B.n131 VSUBS 0.007118f
C342 B.n132 VSUBS 0.007118f
C343 B.n133 VSUBS 0.007118f
C344 B.n134 VSUBS 0.007118f
C345 B.n135 VSUBS 0.007118f
C346 B.n136 VSUBS 0.007118f
C347 B.n137 VSUBS 0.007118f
C348 B.n138 VSUBS 0.007118f
C349 B.n139 VSUBS 0.007118f
C350 B.n140 VSUBS 0.007118f
C351 B.n141 VSUBS 0.007118f
C352 B.n142 VSUBS 0.007118f
C353 B.n143 VSUBS 0.007118f
C354 B.n144 VSUBS 0.007118f
C355 B.n145 VSUBS 0.007118f
C356 B.n146 VSUBS 0.007118f
C357 B.n147 VSUBS 0.007118f
C358 B.n148 VSUBS 0.007118f
C359 B.n149 VSUBS 0.007118f
C360 B.n150 VSUBS 0.007118f
C361 B.n151 VSUBS 0.007118f
C362 B.n152 VSUBS 0.014866f
C363 B.n153 VSUBS 0.014866f
C364 B.n154 VSUBS 0.01591f
C365 B.n155 VSUBS 0.007118f
C366 B.n156 VSUBS 0.007118f
C367 B.n157 VSUBS 0.007118f
C368 B.n158 VSUBS 0.007118f
C369 B.n159 VSUBS 0.007118f
C370 B.n160 VSUBS 0.007118f
C371 B.n161 VSUBS 0.007118f
C372 B.n162 VSUBS 0.007118f
C373 B.n163 VSUBS 0.007118f
C374 B.n164 VSUBS 0.007118f
C375 B.n165 VSUBS 0.007118f
C376 B.n166 VSUBS 0.007118f
C377 B.n167 VSUBS 0.007118f
C378 B.n168 VSUBS 0.007118f
C379 B.n169 VSUBS 0.007118f
C380 B.n170 VSUBS 0.007118f
C381 B.n171 VSUBS 0.007118f
C382 B.n172 VSUBS 0.007118f
C383 B.n173 VSUBS 0.007118f
C384 B.n174 VSUBS 0.007118f
C385 B.n175 VSUBS 0.007118f
C386 B.n176 VSUBS 0.007118f
C387 B.n177 VSUBS 0.007118f
C388 B.n178 VSUBS 0.007118f
C389 B.n179 VSUBS 0.006752f
C390 B.n180 VSUBS 0.007118f
C391 B.n181 VSUBS 0.007118f
C392 B.n182 VSUBS 0.003925f
C393 B.n183 VSUBS 0.007118f
C394 B.n184 VSUBS 0.007118f
C395 B.n185 VSUBS 0.007118f
C396 B.n186 VSUBS 0.007118f
C397 B.n187 VSUBS 0.007118f
C398 B.n188 VSUBS 0.007118f
C399 B.n189 VSUBS 0.007118f
C400 B.n190 VSUBS 0.007118f
C401 B.n191 VSUBS 0.007118f
C402 B.n192 VSUBS 0.007118f
C403 B.n193 VSUBS 0.007118f
C404 B.n194 VSUBS 0.007118f
C405 B.n195 VSUBS 0.003925f
C406 B.n196 VSUBS 0.016492f
C407 B.n197 VSUBS 0.006752f
C408 B.n198 VSUBS 0.007118f
C409 B.n199 VSUBS 0.007118f
C410 B.n200 VSUBS 0.007118f
C411 B.n201 VSUBS 0.007118f
C412 B.n202 VSUBS 0.007118f
C413 B.n203 VSUBS 0.007118f
C414 B.n204 VSUBS 0.007118f
C415 B.n205 VSUBS 0.007118f
C416 B.n206 VSUBS 0.007118f
C417 B.n207 VSUBS 0.007118f
C418 B.n208 VSUBS 0.007118f
C419 B.n209 VSUBS 0.007118f
C420 B.n210 VSUBS 0.007118f
C421 B.n211 VSUBS 0.007118f
C422 B.n212 VSUBS 0.007118f
C423 B.n213 VSUBS 0.007118f
C424 B.n214 VSUBS 0.007118f
C425 B.n215 VSUBS 0.007118f
C426 B.n216 VSUBS 0.007118f
C427 B.n217 VSUBS 0.007118f
C428 B.n218 VSUBS 0.007118f
C429 B.n219 VSUBS 0.007118f
C430 B.n220 VSUBS 0.007118f
C431 B.n221 VSUBS 0.007118f
C432 B.n222 VSUBS 0.007118f
C433 B.n223 VSUBS 0.01591f
C434 B.n224 VSUBS 0.014866f
C435 B.n225 VSUBS 0.014866f
C436 B.n226 VSUBS 0.007118f
C437 B.n227 VSUBS 0.007118f
C438 B.n228 VSUBS 0.007118f
C439 B.n229 VSUBS 0.007118f
C440 B.n230 VSUBS 0.007118f
C441 B.n231 VSUBS 0.007118f
C442 B.n232 VSUBS 0.007118f
C443 B.n233 VSUBS 0.007118f
C444 B.n234 VSUBS 0.007118f
C445 B.n235 VSUBS 0.007118f
C446 B.n236 VSUBS 0.007118f
C447 B.n237 VSUBS 0.007118f
C448 B.n238 VSUBS 0.007118f
C449 B.n239 VSUBS 0.007118f
C450 B.n240 VSUBS 0.007118f
C451 B.n241 VSUBS 0.007118f
C452 B.n242 VSUBS 0.007118f
C453 B.n243 VSUBS 0.007118f
C454 B.n244 VSUBS 0.007118f
C455 B.n245 VSUBS 0.007118f
C456 B.n246 VSUBS 0.007118f
C457 B.n247 VSUBS 0.007118f
C458 B.n248 VSUBS 0.007118f
C459 B.n249 VSUBS 0.007118f
C460 B.n250 VSUBS 0.007118f
C461 B.n251 VSUBS 0.007118f
C462 B.n252 VSUBS 0.007118f
C463 B.n253 VSUBS 0.007118f
C464 B.n254 VSUBS 0.007118f
C465 B.n255 VSUBS 0.007118f
C466 B.n256 VSUBS 0.007118f
C467 B.n257 VSUBS 0.007118f
C468 B.n258 VSUBS 0.007118f
C469 B.n259 VSUBS 0.007118f
C470 B.n260 VSUBS 0.007118f
C471 B.n261 VSUBS 0.007118f
C472 B.n262 VSUBS 0.007118f
C473 B.n263 VSUBS 0.007118f
C474 B.n264 VSUBS 0.007118f
C475 B.n265 VSUBS 0.007118f
C476 B.n266 VSUBS 0.007118f
C477 B.n267 VSUBS 0.007118f
C478 B.n268 VSUBS 0.007118f
C479 B.n269 VSUBS 0.007118f
C480 B.n270 VSUBS 0.007118f
C481 B.n271 VSUBS 0.007118f
C482 B.n272 VSUBS 0.007118f
C483 B.n273 VSUBS 0.007118f
C484 B.n274 VSUBS 0.007118f
C485 B.n275 VSUBS 0.007118f
C486 B.n276 VSUBS 0.007118f
C487 B.n277 VSUBS 0.007118f
C488 B.n278 VSUBS 0.007118f
C489 B.n279 VSUBS 0.007118f
C490 B.n280 VSUBS 0.007118f
C491 B.n281 VSUBS 0.007118f
C492 B.n282 VSUBS 0.007118f
C493 B.n283 VSUBS 0.007118f
C494 B.n284 VSUBS 0.007118f
C495 B.n285 VSUBS 0.007118f
C496 B.n286 VSUBS 0.007118f
C497 B.n287 VSUBS 0.007118f
C498 B.n288 VSUBS 0.007118f
C499 B.n289 VSUBS 0.007118f
C500 B.n290 VSUBS 0.007118f
C501 B.n291 VSUBS 0.007118f
C502 B.n292 VSUBS 0.007118f
C503 B.n293 VSUBS 0.007118f
C504 B.n294 VSUBS 0.007118f
C505 B.n295 VSUBS 0.007118f
C506 B.n296 VSUBS 0.007118f
C507 B.n297 VSUBS 0.007118f
C508 B.n298 VSUBS 0.007118f
C509 B.n299 VSUBS 0.007118f
C510 B.n300 VSUBS 0.007118f
C511 B.n301 VSUBS 0.007118f
C512 B.n302 VSUBS 0.007118f
C513 B.n303 VSUBS 0.007118f
C514 B.n304 VSUBS 0.007118f
C515 B.n305 VSUBS 0.007118f
C516 B.n306 VSUBS 0.007118f
C517 B.n307 VSUBS 0.007118f
C518 B.n308 VSUBS 0.014866f
C519 B.n309 VSUBS 0.015817f
C520 B.n310 VSUBS 0.014958f
C521 B.n311 VSUBS 0.007118f
C522 B.n312 VSUBS 0.007118f
C523 B.n313 VSUBS 0.007118f
C524 B.n314 VSUBS 0.007118f
C525 B.n315 VSUBS 0.007118f
C526 B.n316 VSUBS 0.007118f
C527 B.n317 VSUBS 0.007118f
C528 B.n318 VSUBS 0.007118f
C529 B.n319 VSUBS 0.007118f
C530 B.n320 VSUBS 0.007118f
C531 B.n321 VSUBS 0.007118f
C532 B.n322 VSUBS 0.007118f
C533 B.n323 VSUBS 0.007118f
C534 B.n324 VSUBS 0.007118f
C535 B.n325 VSUBS 0.007118f
C536 B.n326 VSUBS 0.007118f
C537 B.n327 VSUBS 0.007118f
C538 B.n328 VSUBS 0.007118f
C539 B.n329 VSUBS 0.007118f
C540 B.n330 VSUBS 0.007118f
C541 B.n331 VSUBS 0.007118f
C542 B.n332 VSUBS 0.007118f
C543 B.n333 VSUBS 0.007118f
C544 B.n334 VSUBS 0.007118f
C545 B.n335 VSUBS 0.006752f
C546 B.n336 VSUBS 0.007118f
C547 B.n337 VSUBS 0.007118f
C548 B.n338 VSUBS 0.003925f
C549 B.n339 VSUBS 0.007118f
C550 B.n340 VSUBS 0.007118f
C551 B.n341 VSUBS 0.007118f
C552 B.n342 VSUBS 0.007118f
C553 B.n343 VSUBS 0.007118f
C554 B.n344 VSUBS 0.007118f
C555 B.n345 VSUBS 0.007118f
C556 B.n346 VSUBS 0.007118f
C557 B.n347 VSUBS 0.007118f
C558 B.n348 VSUBS 0.007118f
C559 B.n349 VSUBS 0.007118f
C560 B.n350 VSUBS 0.007118f
C561 B.n351 VSUBS 0.003925f
C562 B.n352 VSUBS 0.016492f
C563 B.n353 VSUBS 0.006752f
C564 B.n354 VSUBS 0.007118f
C565 B.n355 VSUBS 0.007118f
C566 B.n356 VSUBS 0.007118f
C567 B.n357 VSUBS 0.007118f
C568 B.n358 VSUBS 0.007118f
C569 B.n359 VSUBS 0.007118f
C570 B.n360 VSUBS 0.007118f
C571 B.n361 VSUBS 0.007118f
C572 B.n362 VSUBS 0.007118f
C573 B.n363 VSUBS 0.007118f
C574 B.n364 VSUBS 0.007118f
C575 B.n365 VSUBS 0.007118f
C576 B.n366 VSUBS 0.007118f
C577 B.n367 VSUBS 0.007118f
C578 B.n368 VSUBS 0.007118f
C579 B.n369 VSUBS 0.007118f
C580 B.n370 VSUBS 0.007118f
C581 B.n371 VSUBS 0.007118f
C582 B.n372 VSUBS 0.007118f
C583 B.n373 VSUBS 0.007118f
C584 B.n374 VSUBS 0.007118f
C585 B.n375 VSUBS 0.007118f
C586 B.n376 VSUBS 0.007118f
C587 B.n377 VSUBS 0.007118f
C588 B.n378 VSUBS 0.007118f
C589 B.n379 VSUBS 0.01591f
C590 B.n380 VSUBS 0.014866f
C591 B.n381 VSUBS 0.014866f
C592 B.n382 VSUBS 0.007118f
C593 B.n383 VSUBS 0.007118f
C594 B.n384 VSUBS 0.007118f
C595 B.n385 VSUBS 0.007118f
C596 B.n386 VSUBS 0.007118f
C597 B.n387 VSUBS 0.007118f
C598 B.n388 VSUBS 0.007118f
C599 B.n389 VSUBS 0.007118f
C600 B.n390 VSUBS 0.007118f
C601 B.n391 VSUBS 0.007118f
C602 B.n392 VSUBS 0.007118f
C603 B.n393 VSUBS 0.007118f
C604 B.n394 VSUBS 0.007118f
C605 B.n395 VSUBS 0.007118f
C606 B.n396 VSUBS 0.007118f
C607 B.n397 VSUBS 0.007118f
C608 B.n398 VSUBS 0.007118f
C609 B.n399 VSUBS 0.007118f
C610 B.n400 VSUBS 0.007118f
C611 B.n401 VSUBS 0.007118f
C612 B.n402 VSUBS 0.007118f
C613 B.n403 VSUBS 0.007118f
C614 B.n404 VSUBS 0.007118f
C615 B.n405 VSUBS 0.007118f
C616 B.n406 VSUBS 0.007118f
C617 B.n407 VSUBS 0.007118f
C618 B.n408 VSUBS 0.007118f
C619 B.n409 VSUBS 0.007118f
C620 B.n410 VSUBS 0.007118f
C621 B.n411 VSUBS 0.007118f
C622 B.n412 VSUBS 0.007118f
C623 B.n413 VSUBS 0.007118f
C624 B.n414 VSUBS 0.007118f
C625 B.n415 VSUBS 0.007118f
C626 B.n416 VSUBS 0.007118f
C627 B.n417 VSUBS 0.007118f
C628 B.n418 VSUBS 0.007118f
C629 B.n419 VSUBS 0.007118f
C630 B.n420 VSUBS 0.007118f
C631 B.n421 VSUBS 0.007118f
C632 B.n422 VSUBS 0.007118f
C633 B.n423 VSUBS 0.016118f
.ends

