* NGSPICE file created from diff_pair_sample_1083.ext - technology: sky130A

.subckt diff_pair_sample_1083 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.34155 pd=2.4 as=0.8073 ps=4.92 w=2.07 l=1.98
X1 VDD1.t2 VP.t1 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.34155 pd=2.4 as=0.8073 ps=4.92 w=2.07 l=1.98
X2 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0.34155 ps=2.4 w=2.07 l=1.98
X3 VTAIL.t5 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0.34155 ps=2.4 w=2.07 l=1.98
X4 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0 ps=0 w=2.07 l=1.98
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0 ps=0 w=2.07 l=1.98
X6 VTAIL.t6 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0.34155 ps=2.4 w=2.07 l=1.98
X7 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.34155 pd=2.4 as=0.8073 ps=4.92 w=2.07 l=1.98
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0 ps=0 w=2.07 l=1.98
X9 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.34155 pd=2.4 as=0.8073 ps=4.92 w=2.07 l=1.98
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0 ps=0 w=2.07 l=1.98
X11 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8073 pd=4.92 as=0.34155 ps=2.4 w=2.07 l=1.98
R0 VP.n10 VP.n0 161.3
R1 VP.n9 VP.n8 161.3
R2 VP.n7 VP.n1 161.3
R3 VP.n6 VP.n5 161.3
R4 VP.n4 VP.n3 90.9382
R5 VP.n12 VP.n11 90.9382
R6 VP.n2 VP.t3 60.6711
R7 VP.n2 VP.t1 60.1424
R8 VP.n9 VP.n1 56.5193
R9 VP.n3 VP.n2 44.192
R10 VP.n4 VP.t2 25.196
R11 VP.n11 VP.t0 25.196
R12 VP.n5 VP.n1 24.4675
R13 VP.n10 VP.n9 24.4675
R14 VP.n5 VP.n4 19.8188
R15 VP.n11 VP.n10 19.8188
R16 VP.n6 VP.n3 0.278367
R17 VP.n12 VP.n0 0.278367
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153454
R22 VTAIL.n7 VTAIL.t1 84.2207
R23 VTAIL.n0 VTAIL.t2 84.2207
R24 VTAIL.n1 VTAIL.t7 84.2207
R25 VTAIL.n2 VTAIL.t5 84.2207
R26 VTAIL.n6 VTAIL.t4 84.2207
R27 VTAIL.n5 VTAIL.t6 84.2206
R28 VTAIL.n4 VTAIL.t0 84.2206
R29 VTAIL.n3 VTAIL.t3 84.2206
R30 VTAIL.n7 VTAIL.n6 16.1427
R31 VTAIL.n3 VTAIL.n2 16.1427
R32 VTAIL.n4 VTAIL.n3 1.99188
R33 VTAIL.n6 VTAIL.n5 1.99188
R34 VTAIL.n2 VTAIL.n1 1.99188
R35 VTAIL VTAIL.n0 1.05438
R36 VTAIL VTAIL.n7 0.938
R37 VTAIL.n5 VTAIL.n4 0.470328
R38 VTAIL.n1 VTAIL.n0 0.470328
R39 VDD1 VDD1.n1 123.332
R40 VDD1 VDD1.n0 91.3925
R41 VDD1.n0 VDD1.t0 9.56572
R42 VDD1.n0 VDD1.t2 9.56572
R43 VDD1.n1 VDD1.t1 9.56572
R44 VDD1.n1 VDD1.t3 9.56572
R45 B.n409 B.n408 585
R46 B.n141 B.n72 585
R47 B.n140 B.n139 585
R48 B.n138 B.n137 585
R49 B.n136 B.n135 585
R50 B.n134 B.n133 585
R51 B.n132 B.n131 585
R52 B.n130 B.n129 585
R53 B.n128 B.n127 585
R54 B.n126 B.n125 585
R55 B.n124 B.n123 585
R56 B.n122 B.n121 585
R57 B.n120 B.n119 585
R58 B.n118 B.n117 585
R59 B.n116 B.n115 585
R60 B.n114 B.n113 585
R61 B.n112 B.n111 585
R62 B.n110 B.n109 585
R63 B.n108 B.n107 585
R64 B.n106 B.n105 585
R65 B.n104 B.n103 585
R66 B.n102 B.n101 585
R67 B.n100 B.n99 585
R68 B.n98 B.n97 585
R69 B.n96 B.n95 585
R70 B.n94 B.n93 585
R71 B.n92 B.n91 585
R72 B.n90 B.n89 585
R73 B.n88 B.n87 585
R74 B.n86 B.n85 585
R75 B.n84 B.n83 585
R76 B.n82 B.n81 585
R77 B.n80 B.n79 585
R78 B.n54 B.n53 585
R79 B.n407 B.n55 585
R80 B.n412 B.n55 585
R81 B.n406 B.n405 585
R82 B.n405 B.n51 585
R83 B.n404 B.n50 585
R84 B.n418 B.n50 585
R85 B.n403 B.n49 585
R86 B.n419 B.n49 585
R87 B.n402 B.n48 585
R88 B.n420 B.n48 585
R89 B.n401 B.n400 585
R90 B.n400 B.n44 585
R91 B.n399 B.n43 585
R92 B.n426 B.n43 585
R93 B.n398 B.n42 585
R94 B.n427 B.n42 585
R95 B.n397 B.n41 585
R96 B.n428 B.n41 585
R97 B.n396 B.n395 585
R98 B.n395 B.n37 585
R99 B.n394 B.n36 585
R100 B.n434 B.n36 585
R101 B.n393 B.n35 585
R102 B.n435 B.n35 585
R103 B.n392 B.n34 585
R104 B.n436 B.n34 585
R105 B.n391 B.n390 585
R106 B.n390 B.n30 585
R107 B.n389 B.n29 585
R108 B.n442 B.n29 585
R109 B.n388 B.n28 585
R110 B.n443 B.n28 585
R111 B.n387 B.n27 585
R112 B.n444 B.n27 585
R113 B.n386 B.n385 585
R114 B.n385 B.n23 585
R115 B.n384 B.n22 585
R116 B.n450 B.n22 585
R117 B.n383 B.n21 585
R118 B.n451 B.n21 585
R119 B.n382 B.n20 585
R120 B.n452 B.n20 585
R121 B.n381 B.n380 585
R122 B.n380 B.n16 585
R123 B.n379 B.n15 585
R124 B.n458 B.n15 585
R125 B.n378 B.n14 585
R126 B.n459 B.n14 585
R127 B.n377 B.n13 585
R128 B.n460 B.n13 585
R129 B.n376 B.n375 585
R130 B.n375 B.n12 585
R131 B.n374 B.n373 585
R132 B.n374 B.n8 585
R133 B.n372 B.n7 585
R134 B.n467 B.n7 585
R135 B.n371 B.n6 585
R136 B.n468 B.n6 585
R137 B.n370 B.n5 585
R138 B.n469 B.n5 585
R139 B.n369 B.n368 585
R140 B.n368 B.n4 585
R141 B.n367 B.n142 585
R142 B.n367 B.n366 585
R143 B.n357 B.n143 585
R144 B.n144 B.n143 585
R145 B.n359 B.n358 585
R146 B.n360 B.n359 585
R147 B.n356 B.n148 585
R148 B.n152 B.n148 585
R149 B.n355 B.n354 585
R150 B.n354 B.n353 585
R151 B.n150 B.n149 585
R152 B.n151 B.n150 585
R153 B.n346 B.n345 585
R154 B.n347 B.n346 585
R155 B.n344 B.n157 585
R156 B.n157 B.n156 585
R157 B.n343 B.n342 585
R158 B.n342 B.n341 585
R159 B.n159 B.n158 585
R160 B.n160 B.n159 585
R161 B.n334 B.n333 585
R162 B.n335 B.n334 585
R163 B.n332 B.n165 585
R164 B.n165 B.n164 585
R165 B.n331 B.n330 585
R166 B.n330 B.n329 585
R167 B.n167 B.n166 585
R168 B.n168 B.n167 585
R169 B.n322 B.n321 585
R170 B.n323 B.n322 585
R171 B.n320 B.n173 585
R172 B.n173 B.n172 585
R173 B.n319 B.n318 585
R174 B.n318 B.n317 585
R175 B.n175 B.n174 585
R176 B.n176 B.n175 585
R177 B.n310 B.n309 585
R178 B.n311 B.n310 585
R179 B.n308 B.n181 585
R180 B.n181 B.n180 585
R181 B.n307 B.n306 585
R182 B.n306 B.n305 585
R183 B.n183 B.n182 585
R184 B.n184 B.n183 585
R185 B.n298 B.n297 585
R186 B.n299 B.n298 585
R187 B.n296 B.n189 585
R188 B.n189 B.n188 585
R189 B.n295 B.n294 585
R190 B.n294 B.n293 585
R191 B.n191 B.n190 585
R192 B.n192 B.n191 585
R193 B.n286 B.n285 585
R194 B.n287 B.n286 585
R195 B.n195 B.n194 585
R196 B.n218 B.n216 585
R197 B.n219 B.n215 585
R198 B.n219 B.n196 585
R199 B.n222 B.n221 585
R200 B.n223 B.n214 585
R201 B.n225 B.n224 585
R202 B.n227 B.n213 585
R203 B.n230 B.n229 585
R204 B.n231 B.n212 585
R205 B.n233 B.n232 585
R206 B.n235 B.n211 585
R207 B.n238 B.n237 585
R208 B.n240 B.n208 585
R209 B.n242 B.n241 585
R210 B.n244 B.n207 585
R211 B.n247 B.n246 585
R212 B.n248 B.n206 585
R213 B.n250 B.n249 585
R214 B.n252 B.n205 585
R215 B.n255 B.n254 585
R216 B.n256 B.n204 585
R217 B.n261 B.n260 585
R218 B.n263 B.n203 585
R219 B.n266 B.n265 585
R220 B.n267 B.n202 585
R221 B.n269 B.n268 585
R222 B.n271 B.n201 585
R223 B.n274 B.n273 585
R224 B.n275 B.n200 585
R225 B.n277 B.n276 585
R226 B.n279 B.n199 585
R227 B.n280 B.n198 585
R228 B.n283 B.n282 585
R229 B.n284 B.n197 585
R230 B.n197 B.n196 585
R231 B.n289 B.n288 585
R232 B.n288 B.n287 585
R233 B.n290 B.n193 585
R234 B.n193 B.n192 585
R235 B.n292 B.n291 585
R236 B.n293 B.n292 585
R237 B.n187 B.n186 585
R238 B.n188 B.n187 585
R239 B.n301 B.n300 585
R240 B.n300 B.n299 585
R241 B.n302 B.n185 585
R242 B.n185 B.n184 585
R243 B.n304 B.n303 585
R244 B.n305 B.n304 585
R245 B.n179 B.n178 585
R246 B.n180 B.n179 585
R247 B.n313 B.n312 585
R248 B.n312 B.n311 585
R249 B.n314 B.n177 585
R250 B.n177 B.n176 585
R251 B.n316 B.n315 585
R252 B.n317 B.n316 585
R253 B.n171 B.n170 585
R254 B.n172 B.n171 585
R255 B.n325 B.n324 585
R256 B.n324 B.n323 585
R257 B.n326 B.n169 585
R258 B.n169 B.n168 585
R259 B.n328 B.n327 585
R260 B.n329 B.n328 585
R261 B.n163 B.n162 585
R262 B.n164 B.n163 585
R263 B.n337 B.n336 585
R264 B.n336 B.n335 585
R265 B.n338 B.n161 585
R266 B.n161 B.n160 585
R267 B.n340 B.n339 585
R268 B.n341 B.n340 585
R269 B.n155 B.n154 585
R270 B.n156 B.n155 585
R271 B.n349 B.n348 585
R272 B.n348 B.n347 585
R273 B.n350 B.n153 585
R274 B.n153 B.n151 585
R275 B.n352 B.n351 585
R276 B.n353 B.n352 585
R277 B.n147 B.n146 585
R278 B.n152 B.n147 585
R279 B.n362 B.n361 585
R280 B.n361 B.n360 585
R281 B.n363 B.n145 585
R282 B.n145 B.n144 585
R283 B.n365 B.n364 585
R284 B.n366 B.n365 585
R285 B.n3 B.n0 585
R286 B.n4 B.n3 585
R287 B.n466 B.n1 585
R288 B.n467 B.n466 585
R289 B.n465 B.n464 585
R290 B.n465 B.n8 585
R291 B.n463 B.n9 585
R292 B.n12 B.n9 585
R293 B.n462 B.n461 585
R294 B.n461 B.n460 585
R295 B.n11 B.n10 585
R296 B.n459 B.n11 585
R297 B.n457 B.n456 585
R298 B.n458 B.n457 585
R299 B.n455 B.n17 585
R300 B.n17 B.n16 585
R301 B.n454 B.n453 585
R302 B.n453 B.n452 585
R303 B.n19 B.n18 585
R304 B.n451 B.n19 585
R305 B.n449 B.n448 585
R306 B.n450 B.n449 585
R307 B.n447 B.n24 585
R308 B.n24 B.n23 585
R309 B.n446 B.n445 585
R310 B.n445 B.n444 585
R311 B.n26 B.n25 585
R312 B.n443 B.n26 585
R313 B.n441 B.n440 585
R314 B.n442 B.n441 585
R315 B.n439 B.n31 585
R316 B.n31 B.n30 585
R317 B.n438 B.n437 585
R318 B.n437 B.n436 585
R319 B.n33 B.n32 585
R320 B.n435 B.n33 585
R321 B.n433 B.n432 585
R322 B.n434 B.n433 585
R323 B.n431 B.n38 585
R324 B.n38 B.n37 585
R325 B.n430 B.n429 585
R326 B.n429 B.n428 585
R327 B.n40 B.n39 585
R328 B.n427 B.n40 585
R329 B.n425 B.n424 585
R330 B.n426 B.n425 585
R331 B.n423 B.n45 585
R332 B.n45 B.n44 585
R333 B.n422 B.n421 585
R334 B.n421 B.n420 585
R335 B.n47 B.n46 585
R336 B.n419 B.n47 585
R337 B.n417 B.n416 585
R338 B.n418 B.n417 585
R339 B.n415 B.n52 585
R340 B.n52 B.n51 585
R341 B.n414 B.n413 585
R342 B.n413 B.n412 585
R343 B.n470 B.n469 585
R344 B.n468 B.n2 585
R345 B.n413 B.n54 530.939
R346 B.n409 B.n55 530.939
R347 B.n286 B.n197 530.939
R348 B.n288 B.n195 530.939
R349 B.n411 B.n410 256.663
R350 B.n411 B.n71 256.663
R351 B.n411 B.n70 256.663
R352 B.n411 B.n69 256.663
R353 B.n411 B.n68 256.663
R354 B.n411 B.n67 256.663
R355 B.n411 B.n66 256.663
R356 B.n411 B.n65 256.663
R357 B.n411 B.n64 256.663
R358 B.n411 B.n63 256.663
R359 B.n411 B.n62 256.663
R360 B.n411 B.n61 256.663
R361 B.n411 B.n60 256.663
R362 B.n411 B.n59 256.663
R363 B.n411 B.n58 256.663
R364 B.n411 B.n57 256.663
R365 B.n411 B.n56 256.663
R366 B.n217 B.n196 256.663
R367 B.n220 B.n196 256.663
R368 B.n226 B.n196 256.663
R369 B.n228 B.n196 256.663
R370 B.n234 B.n196 256.663
R371 B.n236 B.n196 256.663
R372 B.n243 B.n196 256.663
R373 B.n245 B.n196 256.663
R374 B.n251 B.n196 256.663
R375 B.n253 B.n196 256.663
R376 B.n262 B.n196 256.663
R377 B.n264 B.n196 256.663
R378 B.n270 B.n196 256.663
R379 B.n272 B.n196 256.663
R380 B.n278 B.n196 256.663
R381 B.n281 B.n196 256.663
R382 B.n472 B.n471 256.663
R383 B.n76 B.t15 232.065
R384 B.n73 B.t8 232.065
R385 B.n257 B.t12 232.065
R386 B.n209 B.t4 232.065
R387 B.n287 B.n196 184.208
R388 B.n412 B.n411 184.208
R389 B.n81 B.n80 163.367
R390 B.n85 B.n84 163.367
R391 B.n89 B.n88 163.367
R392 B.n93 B.n92 163.367
R393 B.n97 B.n96 163.367
R394 B.n101 B.n100 163.367
R395 B.n105 B.n104 163.367
R396 B.n109 B.n108 163.367
R397 B.n113 B.n112 163.367
R398 B.n117 B.n116 163.367
R399 B.n121 B.n120 163.367
R400 B.n125 B.n124 163.367
R401 B.n129 B.n128 163.367
R402 B.n133 B.n132 163.367
R403 B.n137 B.n136 163.367
R404 B.n139 B.n72 163.367
R405 B.n286 B.n191 163.367
R406 B.n294 B.n191 163.367
R407 B.n294 B.n189 163.367
R408 B.n298 B.n189 163.367
R409 B.n298 B.n183 163.367
R410 B.n306 B.n183 163.367
R411 B.n306 B.n181 163.367
R412 B.n310 B.n181 163.367
R413 B.n310 B.n175 163.367
R414 B.n318 B.n175 163.367
R415 B.n318 B.n173 163.367
R416 B.n322 B.n173 163.367
R417 B.n322 B.n167 163.367
R418 B.n330 B.n167 163.367
R419 B.n330 B.n165 163.367
R420 B.n334 B.n165 163.367
R421 B.n334 B.n159 163.367
R422 B.n342 B.n159 163.367
R423 B.n342 B.n157 163.367
R424 B.n346 B.n157 163.367
R425 B.n346 B.n150 163.367
R426 B.n354 B.n150 163.367
R427 B.n354 B.n148 163.367
R428 B.n359 B.n148 163.367
R429 B.n359 B.n143 163.367
R430 B.n367 B.n143 163.367
R431 B.n368 B.n367 163.367
R432 B.n368 B.n5 163.367
R433 B.n6 B.n5 163.367
R434 B.n7 B.n6 163.367
R435 B.n374 B.n7 163.367
R436 B.n375 B.n374 163.367
R437 B.n375 B.n13 163.367
R438 B.n14 B.n13 163.367
R439 B.n15 B.n14 163.367
R440 B.n380 B.n15 163.367
R441 B.n380 B.n20 163.367
R442 B.n21 B.n20 163.367
R443 B.n22 B.n21 163.367
R444 B.n385 B.n22 163.367
R445 B.n385 B.n27 163.367
R446 B.n28 B.n27 163.367
R447 B.n29 B.n28 163.367
R448 B.n390 B.n29 163.367
R449 B.n390 B.n34 163.367
R450 B.n35 B.n34 163.367
R451 B.n36 B.n35 163.367
R452 B.n395 B.n36 163.367
R453 B.n395 B.n41 163.367
R454 B.n42 B.n41 163.367
R455 B.n43 B.n42 163.367
R456 B.n400 B.n43 163.367
R457 B.n400 B.n48 163.367
R458 B.n49 B.n48 163.367
R459 B.n50 B.n49 163.367
R460 B.n405 B.n50 163.367
R461 B.n405 B.n55 163.367
R462 B.n219 B.n218 163.367
R463 B.n221 B.n219 163.367
R464 B.n225 B.n214 163.367
R465 B.n229 B.n227 163.367
R466 B.n233 B.n212 163.367
R467 B.n237 B.n235 163.367
R468 B.n242 B.n208 163.367
R469 B.n246 B.n244 163.367
R470 B.n250 B.n206 163.367
R471 B.n254 B.n252 163.367
R472 B.n261 B.n204 163.367
R473 B.n265 B.n263 163.367
R474 B.n269 B.n202 163.367
R475 B.n273 B.n271 163.367
R476 B.n277 B.n200 163.367
R477 B.n280 B.n279 163.367
R478 B.n282 B.n197 163.367
R479 B.n288 B.n193 163.367
R480 B.n292 B.n193 163.367
R481 B.n292 B.n187 163.367
R482 B.n300 B.n187 163.367
R483 B.n300 B.n185 163.367
R484 B.n304 B.n185 163.367
R485 B.n304 B.n179 163.367
R486 B.n312 B.n179 163.367
R487 B.n312 B.n177 163.367
R488 B.n316 B.n177 163.367
R489 B.n316 B.n171 163.367
R490 B.n324 B.n171 163.367
R491 B.n324 B.n169 163.367
R492 B.n328 B.n169 163.367
R493 B.n328 B.n163 163.367
R494 B.n336 B.n163 163.367
R495 B.n336 B.n161 163.367
R496 B.n340 B.n161 163.367
R497 B.n340 B.n155 163.367
R498 B.n348 B.n155 163.367
R499 B.n348 B.n153 163.367
R500 B.n352 B.n153 163.367
R501 B.n352 B.n147 163.367
R502 B.n361 B.n147 163.367
R503 B.n361 B.n145 163.367
R504 B.n365 B.n145 163.367
R505 B.n365 B.n3 163.367
R506 B.n470 B.n3 163.367
R507 B.n466 B.n2 163.367
R508 B.n466 B.n465 163.367
R509 B.n465 B.n9 163.367
R510 B.n461 B.n9 163.367
R511 B.n461 B.n11 163.367
R512 B.n457 B.n11 163.367
R513 B.n457 B.n17 163.367
R514 B.n453 B.n17 163.367
R515 B.n453 B.n19 163.367
R516 B.n449 B.n19 163.367
R517 B.n449 B.n24 163.367
R518 B.n445 B.n24 163.367
R519 B.n445 B.n26 163.367
R520 B.n441 B.n26 163.367
R521 B.n441 B.n31 163.367
R522 B.n437 B.n31 163.367
R523 B.n437 B.n33 163.367
R524 B.n433 B.n33 163.367
R525 B.n433 B.n38 163.367
R526 B.n429 B.n38 163.367
R527 B.n429 B.n40 163.367
R528 B.n425 B.n40 163.367
R529 B.n425 B.n45 163.367
R530 B.n421 B.n45 163.367
R531 B.n421 B.n47 163.367
R532 B.n417 B.n47 163.367
R533 B.n417 B.n52 163.367
R534 B.n413 B.n52 163.367
R535 B.n73 B.t10 128.552
R536 B.n257 B.t14 128.552
R537 B.n76 B.t16 128.552
R538 B.n209 B.t7 128.552
R539 B.n287 B.n192 101.838
R540 B.n293 B.n192 101.838
R541 B.n293 B.n188 101.838
R542 B.n299 B.n188 101.838
R543 B.n299 B.n184 101.838
R544 B.n305 B.n184 101.838
R545 B.n311 B.n180 101.838
R546 B.n311 B.n176 101.838
R547 B.n317 B.n176 101.838
R548 B.n317 B.n172 101.838
R549 B.n323 B.n172 101.838
R550 B.n323 B.n168 101.838
R551 B.n329 B.n168 101.838
R552 B.n329 B.n164 101.838
R553 B.n335 B.n164 101.838
R554 B.n341 B.n160 101.838
R555 B.n341 B.n156 101.838
R556 B.n347 B.n156 101.838
R557 B.n347 B.n151 101.838
R558 B.n353 B.n151 101.838
R559 B.n353 B.n152 101.838
R560 B.n360 B.n144 101.838
R561 B.n366 B.n144 101.838
R562 B.n366 B.n4 101.838
R563 B.n469 B.n4 101.838
R564 B.n469 B.n468 101.838
R565 B.n468 B.n467 101.838
R566 B.n467 B.n8 101.838
R567 B.n12 B.n8 101.838
R568 B.n460 B.n12 101.838
R569 B.n459 B.n458 101.838
R570 B.n458 B.n16 101.838
R571 B.n452 B.n16 101.838
R572 B.n452 B.n451 101.838
R573 B.n451 B.n450 101.838
R574 B.n450 B.n23 101.838
R575 B.n444 B.n443 101.838
R576 B.n443 B.n442 101.838
R577 B.n442 B.n30 101.838
R578 B.n436 B.n30 101.838
R579 B.n436 B.n435 101.838
R580 B.n435 B.n434 101.838
R581 B.n434 B.n37 101.838
R582 B.n428 B.n37 101.838
R583 B.n428 B.n427 101.838
R584 B.n426 B.n44 101.838
R585 B.n420 B.n44 101.838
R586 B.n420 B.n419 101.838
R587 B.n419 B.n418 101.838
R588 B.n418 B.n51 101.838
R589 B.n412 B.n51 101.838
R590 B.n74 B.t11 83.7518
R591 B.n258 B.t13 83.7518
R592 B.n77 B.t17 83.7515
R593 B.n210 B.t6 83.7515
R594 B.n305 B.t5 71.8861
R595 B.n335 B.t3 71.8861
R596 B.n444 B.t1 71.8861
R597 B.t9 B.n426 71.8861
R598 B.n56 B.n54 71.676
R599 B.n81 B.n57 71.676
R600 B.n85 B.n58 71.676
R601 B.n89 B.n59 71.676
R602 B.n93 B.n60 71.676
R603 B.n97 B.n61 71.676
R604 B.n101 B.n62 71.676
R605 B.n105 B.n63 71.676
R606 B.n109 B.n64 71.676
R607 B.n113 B.n65 71.676
R608 B.n117 B.n66 71.676
R609 B.n121 B.n67 71.676
R610 B.n125 B.n68 71.676
R611 B.n129 B.n69 71.676
R612 B.n133 B.n70 71.676
R613 B.n137 B.n71 71.676
R614 B.n410 B.n72 71.676
R615 B.n410 B.n409 71.676
R616 B.n139 B.n71 71.676
R617 B.n136 B.n70 71.676
R618 B.n132 B.n69 71.676
R619 B.n128 B.n68 71.676
R620 B.n124 B.n67 71.676
R621 B.n120 B.n66 71.676
R622 B.n116 B.n65 71.676
R623 B.n112 B.n64 71.676
R624 B.n108 B.n63 71.676
R625 B.n104 B.n62 71.676
R626 B.n100 B.n61 71.676
R627 B.n96 B.n60 71.676
R628 B.n92 B.n59 71.676
R629 B.n88 B.n58 71.676
R630 B.n84 B.n57 71.676
R631 B.n80 B.n56 71.676
R632 B.n217 B.n195 71.676
R633 B.n221 B.n220 71.676
R634 B.n226 B.n225 71.676
R635 B.n229 B.n228 71.676
R636 B.n234 B.n233 71.676
R637 B.n237 B.n236 71.676
R638 B.n243 B.n242 71.676
R639 B.n246 B.n245 71.676
R640 B.n251 B.n250 71.676
R641 B.n254 B.n253 71.676
R642 B.n262 B.n261 71.676
R643 B.n265 B.n264 71.676
R644 B.n270 B.n269 71.676
R645 B.n273 B.n272 71.676
R646 B.n278 B.n277 71.676
R647 B.n281 B.n280 71.676
R648 B.n218 B.n217 71.676
R649 B.n220 B.n214 71.676
R650 B.n227 B.n226 71.676
R651 B.n228 B.n212 71.676
R652 B.n235 B.n234 71.676
R653 B.n236 B.n208 71.676
R654 B.n244 B.n243 71.676
R655 B.n245 B.n206 71.676
R656 B.n252 B.n251 71.676
R657 B.n253 B.n204 71.676
R658 B.n263 B.n262 71.676
R659 B.n264 B.n202 71.676
R660 B.n271 B.n270 71.676
R661 B.n272 B.n200 71.676
R662 B.n279 B.n278 71.676
R663 B.n282 B.n281 71.676
R664 B.n471 B.n470 71.676
R665 B.n471 B.n2 71.676
R666 B.n78 B.n77 59.5399
R667 B.n75 B.n74 59.5399
R668 B.n259 B.n258 59.5399
R669 B.n239 B.n210 59.5399
R670 B.n152 B.t0 50.9195
R671 B.n360 B.t0 50.9195
R672 B.n460 B.t2 50.9195
R673 B.t2 B.n459 50.9195
R674 B.n77 B.n76 44.8005
R675 B.n74 B.n73 44.8005
R676 B.n258 B.n257 44.8005
R677 B.n210 B.n209 44.8005
R678 B.n289 B.n194 34.4981
R679 B.n285 B.n284 34.4981
R680 B.n408 B.n407 34.4981
R681 B.n414 B.n53 34.4981
R682 B.t5 B.n180 29.9528
R683 B.t3 B.n160 29.9528
R684 B.t1 B.n23 29.9528
R685 B.n427 B.t9 29.9528
R686 B B.n472 18.0485
R687 B.n290 B.n289 10.6151
R688 B.n291 B.n290 10.6151
R689 B.n291 B.n186 10.6151
R690 B.n301 B.n186 10.6151
R691 B.n302 B.n301 10.6151
R692 B.n303 B.n302 10.6151
R693 B.n303 B.n178 10.6151
R694 B.n313 B.n178 10.6151
R695 B.n314 B.n313 10.6151
R696 B.n315 B.n314 10.6151
R697 B.n315 B.n170 10.6151
R698 B.n325 B.n170 10.6151
R699 B.n326 B.n325 10.6151
R700 B.n327 B.n326 10.6151
R701 B.n327 B.n162 10.6151
R702 B.n337 B.n162 10.6151
R703 B.n338 B.n337 10.6151
R704 B.n339 B.n338 10.6151
R705 B.n339 B.n154 10.6151
R706 B.n349 B.n154 10.6151
R707 B.n350 B.n349 10.6151
R708 B.n351 B.n350 10.6151
R709 B.n351 B.n146 10.6151
R710 B.n362 B.n146 10.6151
R711 B.n363 B.n362 10.6151
R712 B.n364 B.n363 10.6151
R713 B.n364 B.n0 10.6151
R714 B.n216 B.n194 10.6151
R715 B.n216 B.n215 10.6151
R716 B.n222 B.n215 10.6151
R717 B.n223 B.n222 10.6151
R718 B.n224 B.n223 10.6151
R719 B.n224 B.n213 10.6151
R720 B.n230 B.n213 10.6151
R721 B.n231 B.n230 10.6151
R722 B.n232 B.n231 10.6151
R723 B.n232 B.n211 10.6151
R724 B.n238 B.n211 10.6151
R725 B.n241 B.n240 10.6151
R726 B.n241 B.n207 10.6151
R727 B.n247 B.n207 10.6151
R728 B.n248 B.n247 10.6151
R729 B.n249 B.n248 10.6151
R730 B.n249 B.n205 10.6151
R731 B.n255 B.n205 10.6151
R732 B.n256 B.n255 10.6151
R733 B.n260 B.n256 10.6151
R734 B.n266 B.n203 10.6151
R735 B.n267 B.n266 10.6151
R736 B.n268 B.n267 10.6151
R737 B.n268 B.n201 10.6151
R738 B.n274 B.n201 10.6151
R739 B.n275 B.n274 10.6151
R740 B.n276 B.n275 10.6151
R741 B.n276 B.n199 10.6151
R742 B.n199 B.n198 10.6151
R743 B.n283 B.n198 10.6151
R744 B.n284 B.n283 10.6151
R745 B.n285 B.n190 10.6151
R746 B.n295 B.n190 10.6151
R747 B.n296 B.n295 10.6151
R748 B.n297 B.n296 10.6151
R749 B.n297 B.n182 10.6151
R750 B.n307 B.n182 10.6151
R751 B.n308 B.n307 10.6151
R752 B.n309 B.n308 10.6151
R753 B.n309 B.n174 10.6151
R754 B.n319 B.n174 10.6151
R755 B.n320 B.n319 10.6151
R756 B.n321 B.n320 10.6151
R757 B.n321 B.n166 10.6151
R758 B.n331 B.n166 10.6151
R759 B.n332 B.n331 10.6151
R760 B.n333 B.n332 10.6151
R761 B.n333 B.n158 10.6151
R762 B.n343 B.n158 10.6151
R763 B.n344 B.n343 10.6151
R764 B.n345 B.n344 10.6151
R765 B.n345 B.n149 10.6151
R766 B.n355 B.n149 10.6151
R767 B.n356 B.n355 10.6151
R768 B.n358 B.n356 10.6151
R769 B.n358 B.n357 10.6151
R770 B.n357 B.n142 10.6151
R771 B.n369 B.n142 10.6151
R772 B.n370 B.n369 10.6151
R773 B.n371 B.n370 10.6151
R774 B.n372 B.n371 10.6151
R775 B.n373 B.n372 10.6151
R776 B.n376 B.n373 10.6151
R777 B.n377 B.n376 10.6151
R778 B.n378 B.n377 10.6151
R779 B.n379 B.n378 10.6151
R780 B.n381 B.n379 10.6151
R781 B.n382 B.n381 10.6151
R782 B.n383 B.n382 10.6151
R783 B.n384 B.n383 10.6151
R784 B.n386 B.n384 10.6151
R785 B.n387 B.n386 10.6151
R786 B.n388 B.n387 10.6151
R787 B.n389 B.n388 10.6151
R788 B.n391 B.n389 10.6151
R789 B.n392 B.n391 10.6151
R790 B.n393 B.n392 10.6151
R791 B.n394 B.n393 10.6151
R792 B.n396 B.n394 10.6151
R793 B.n397 B.n396 10.6151
R794 B.n398 B.n397 10.6151
R795 B.n399 B.n398 10.6151
R796 B.n401 B.n399 10.6151
R797 B.n402 B.n401 10.6151
R798 B.n403 B.n402 10.6151
R799 B.n404 B.n403 10.6151
R800 B.n406 B.n404 10.6151
R801 B.n407 B.n406 10.6151
R802 B.n464 B.n1 10.6151
R803 B.n464 B.n463 10.6151
R804 B.n463 B.n462 10.6151
R805 B.n462 B.n10 10.6151
R806 B.n456 B.n10 10.6151
R807 B.n456 B.n455 10.6151
R808 B.n455 B.n454 10.6151
R809 B.n454 B.n18 10.6151
R810 B.n448 B.n18 10.6151
R811 B.n448 B.n447 10.6151
R812 B.n447 B.n446 10.6151
R813 B.n446 B.n25 10.6151
R814 B.n440 B.n25 10.6151
R815 B.n440 B.n439 10.6151
R816 B.n439 B.n438 10.6151
R817 B.n438 B.n32 10.6151
R818 B.n432 B.n32 10.6151
R819 B.n432 B.n431 10.6151
R820 B.n431 B.n430 10.6151
R821 B.n430 B.n39 10.6151
R822 B.n424 B.n39 10.6151
R823 B.n424 B.n423 10.6151
R824 B.n423 B.n422 10.6151
R825 B.n422 B.n46 10.6151
R826 B.n416 B.n46 10.6151
R827 B.n416 B.n415 10.6151
R828 B.n415 B.n414 10.6151
R829 B.n79 B.n53 10.6151
R830 B.n82 B.n79 10.6151
R831 B.n83 B.n82 10.6151
R832 B.n86 B.n83 10.6151
R833 B.n87 B.n86 10.6151
R834 B.n90 B.n87 10.6151
R835 B.n91 B.n90 10.6151
R836 B.n94 B.n91 10.6151
R837 B.n95 B.n94 10.6151
R838 B.n98 B.n95 10.6151
R839 B.n99 B.n98 10.6151
R840 B.n103 B.n102 10.6151
R841 B.n106 B.n103 10.6151
R842 B.n107 B.n106 10.6151
R843 B.n110 B.n107 10.6151
R844 B.n111 B.n110 10.6151
R845 B.n114 B.n111 10.6151
R846 B.n115 B.n114 10.6151
R847 B.n118 B.n115 10.6151
R848 B.n119 B.n118 10.6151
R849 B.n123 B.n122 10.6151
R850 B.n126 B.n123 10.6151
R851 B.n127 B.n126 10.6151
R852 B.n130 B.n127 10.6151
R853 B.n131 B.n130 10.6151
R854 B.n134 B.n131 10.6151
R855 B.n135 B.n134 10.6151
R856 B.n138 B.n135 10.6151
R857 B.n140 B.n138 10.6151
R858 B.n141 B.n140 10.6151
R859 B.n408 B.n141 10.6151
R860 B.n239 B.n238 9.36635
R861 B.n259 B.n203 9.36635
R862 B.n99 B.n78 9.36635
R863 B.n122 B.n75 9.36635
R864 B.n472 B.n0 8.11757
R865 B.n472 B.n1 8.11757
R866 B.n240 B.n239 1.24928
R867 B.n260 B.n259 1.24928
R868 B.n102 B.n78 1.24928
R869 B.n119 B.n75 1.24928
R870 VN.n0 VN.t3 60.6711
R871 VN.n1 VN.t1 60.6711
R872 VN.n0 VN.t2 60.1424
R873 VN.n1 VN.t0 60.1424
R874 VN VN.n1 44.4709
R875 VN VN.n0 7.35345
R876 VDD2.n2 VDD2.n0 122.808
R877 VDD2.n2 VDD2.n1 91.3343
R878 VDD2.n1 VDD2.t3 9.56572
R879 VDD2.n1 VDD2.t2 9.56572
R880 VDD2.n0 VDD2.t0 9.56572
R881 VDD2.n0 VDD2.t1 9.56572
R882 VDD2 VDD2.n2 0.0586897
C0 VP VN 3.91458f
C1 VDD2 VDD1 0.879017f
C2 VDD2 VTAIL 2.79419f
C3 VDD1 VN 0.15425f
C4 VDD1 VP 1.23926f
C5 VTAIL VN 1.44743f
C6 VTAIL VP 1.46154f
C7 VTAIL VDD1 2.74414f
C8 VDD2 VN 1.03353f
C9 VDD2 VP 0.361477f
C10 VDD2 B 2.591888f
C11 VDD1 B 4.65311f
C12 VTAIL B 3.476648f
C13 VN B 8.02207f
C14 VP B 6.748226f
C15 VDD2.t0 B 0.033677f
C16 VDD2.t1 B 0.033677f
C17 VDD2.n0 B 0.416762f
C18 VDD2.t3 B 0.033677f
C19 VDD2.t2 B 0.033677f
C20 VDD2.n1 B 0.228076f
C21 VDD2.n2 B 1.88391f
C22 VN.t3 B 0.362572f
C23 VN.t2 B 0.360568f
C24 VN.n0 B 0.25054f
C25 VN.t1 B 0.362572f
C26 VN.t0 B 0.360568f
C27 VN.n1 B 1.05596f
C28 VDD1.t0 B 0.031616f
C29 VDD1.t2 B 0.031616f
C30 VDD1.n0 B 0.214288f
C31 VDD1.t1 B 0.031616f
C32 VDD1.t3 B 0.031616f
C33 VDD1.n1 B 0.403669f
C34 VTAIL.t2 B 0.210041f
C35 VTAIL.n0 B 0.225201f
C36 VTAIL.t7 B 0.210041f
C37 VTAIL.n1 B 0.275536f
C38 VTAIL.t5 B 0.210041f
C39 VTAIL.n2 B 0.679381f
C40 VTAIL.t3 B 0.210043f
C41 VTAIL.n3 B 0.67938f
C42 VTAIL.t0 B 0.210043f
C43 VTAIL.n4 B 0.275535f
C44 VTAIL.t6 B 0.210043f
C45 VTAIL.n5 B 0.275535f
C46 VTAIL.t4 B 0.210041f
C47 VTAIL.n6 B 0.679381f
C48 VTAIL.t1 B 0.210041f
C49 VTAIL.n7 B 0.622798f
C50 VP.n0 B 0.031162f
C51 VP.t0 B 0.227772f
C52 VP.n1 B 0.034505f
C53 VP.t1 B 0.36364f
C54 VP.t3 B 0.365661f
C55 VP.n2 B 1.05273f
C56 VP.n3 B 0.98065f
C57 VP.t2 B 0.227772f
C58 VP.n4 B 0.184014f
C59 VP.n5 B 0.039919f
C60 VP.n6 B 0.031162f
C61 VP.n7 B 0.023636f
C62 VP.n8 B 0.023636f
C63 VP.n9 B 0.034505f
C64 VP.n10 B 0.039919f
C65 VP.n11 B 0.184014f
C66 VP.n12 B 0.028596f
.ends

