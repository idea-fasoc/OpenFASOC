* NGSPICE file created from diff_pair_sample_1610.ext - technology: sky130A

.subckt diff_pair_sample_1610 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=0 ps=0 w=15.13 l=2.35
X1 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=0 ps=0 w=15.13 l=2.35
X2 VTAIL.t18 VP.t0 VDD1.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X3 VTAIL.t8 VN.t0 VDD2.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X4 VDD2.t8 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=2.49645 ps=15.46 w=15.13 l=2.35
X5 VTAIL.t7 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=0 ps=0 w=15.13 l=2.35
X7 VDD1.t1 VP.t1 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=2.49645 ps=15.46 w=15.13 l=2.35
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=0 ps=0 w=15.13 l=2.35
X9 VTAIL.t16 VP.t2 VDD1.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X10 VDD1.t6 VP.t3 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X11 VTAIL.t6 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X12 VTAIL.t5 VN.t4 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X13 VDD1.t5 VP.t4 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X14 VTAIL.t13 VP.t5 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X15 VDD2.t4 VN.t5 VTAIL.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X16 VDD1.t9 VP.t6 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=5.9007 ps=31.04 w=15.13 l=2.35
X17 VTAIL.t11 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
X18 VDD2.t3 VN.t6 VTAIL.t19 B.t2 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=5.9007 ps=31.04 w=15.13 l=2.35
X19 VDD1.t2 VP.t8 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=2.49645 ps=15.46 w=15.13 l=2.35
X20 VDD1.t7 VP.t9 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=5.9007 ps=31.04 w=15.13 l=2.35
X21 VDD2.t2 VN.t7 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9007 pd=31.04 as=2.49645 ps=15.46 w=15.13 l=2.35
X22 VDD2.t1 VN.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=5.9007 ps=31.04 w=15.13 l=2.35
X23 VDD2.t0 VN.t9 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.49645 pd=15.46 as=2.49645 ps=15.46 w=15.13 l=2.35
R0 B.n1009 B.n1008 585
R1 B.n1010 B.n1009 585
R2 B.n380 B.n158 585
R3 B.n379 B.n378 585
R4 B.n377 B.n376 585
R5 B.n375 B.n374 585
R6 B.n373 B.n372 585
R7 B.n371 B.n370 585
R8 B.n369 B.n368 585
R9 B.n367 B.n366 585
R10 B.n365 B.n364 585
R11 B.n363 B.n362 585
R12 B.n361 B.n360 585
R13 B.n359 B.n358 585
R14 B.n357 B.n356 585
R15 B.n355 B.n354 585
R16 B.n353 B.n352 585
R17 B.n351 B.n350 585
R18 B.n349 B.n348 585
R19 B.n347 B.n346 585
R20 B.n345 B.n344 585
R21 B.n343 B.n342 585
R22 B.n341 B.n340 585
R23 B.n339 B.n338 585
R24 B.n337 B.n336 585
R25 B.n335 B.n334 585
R26 B.n333 B.n332 585
R27 B.n331 B.n330 585
R28 B.n329 B.n328 585
R29 B.n327 B.n326 585
R30 B.n325 B.n324 585
R31 B.n323 B.n322 585
R32 B.n321 B.n320 585
R33 B.n319 B.n318 585
R34 B.n317 B.n316 585
R35 B.n315 B.n314 585
R36 B.n313 B.n312 585
R37 B.n311 B.n310 585
R38 B.n309 B.n308 585
R39 B.n307 B.n306 585
R40 B.n305 B.n304 585
R41 B.n303 B.n302 585
R42 B.n301 B.n300 585
R43 B.n299 B.n298 585
R44 B.n297 B.n296 585
R45 B.n295 B.n294 585
R46 B.n293 B.n292 585
R47 B.n291 B.n290 585
R48 B.n289 B.n288 585
R49 B.n287 B.n286 585
R50 B.n285 B.n284 585
R51 B.n283 B.n282 585
R52 B.n281 B.n280 585
R53 B.n279 B.n278 585
R54 B.n277 B.n276 585
R55 B.n275 B.n274 585
R56 B.n273 B.n272 585
R57 B.n271 B.n270 585
R58 B.n269 B.n268 585
R59 B.n267 B.n266 585
R60 B.n265 B.n264 585
R61 B.n262 B.n261 585
R62 B.n260 B.n259 585
R63 B.n258 B.n257 585
R64 B.n256 B.n255 585
R65 B.n254 B.n253 585
R66 B.n252 B.n251 585
R67 B.n250 B.n249 585
R68 B.n248 B.n247 585
R69 B.n246 B.n245 585
R70 B.n244 B.n243 585
R71 B.n242 B.n241 585
R72 B.n240 B.n239 585
R73 B.n238 B.n237 585
R74 B.n236 B.n235 585
R75 B.n234 B.n233 585
R76 B.n232 B.n231 585
R77 B.n230 B.n229 585
R78 B.n228 B.n227 585
R79 B.n226 B.n225 585
R80 B.n224 B.n223 585
R81 B.n222 B.n221 585
R82 B.n220 B.n219 585
R83 B.n218 B.n217 585
R84 B.n216 B.n215 585
R85 B.n214 B.n213 585
R86 B.n212 B.n211 585
R87 B.n210 B.n209 585
R88 B.n208 B.n207 585
R89 B.n206 B.n205 585
R90 B.n204 B.n203 585
R91 B.n202 B.n201 585
R92 B.n200 B.n199 585
R93 B.n198 B.n197 585
R94 B.n196 B.n195 585
R95 B.n194 B.n193 585
R96 B.n192 B.n191 585
R97 B.n190 B.n189 585
R98 B.n188 B.n187 585
R99 B.n186 B.n185 585
R100 B.n184 B.n183 585
R101 B.n182 B.n181 585
R102 B.n180 B.n179 585
R103 B.n178 B.n177 585
R104 B.n176 B.n175 585
R105 B.n174 B.n173 585
R106 B.n172 B.n171 585
R107 B.n170 B.n169 585
R108 B.n168 B.n167 585
R109 B.n166 B.n165 585
R110 B.n103 B.n102 585
R111 B.n1013 B.n1012 585
R112 B.n1007 B.n159 585
R113 B.n159 B.n100 585
R114 B.n1006 B.n99 585
R115 B.n1017 B.n99 585
R116 B.n1005 B.n98 585
R117 B.n1018 B.n98 585
R118 B.n1004 B.n97 585
R119 B.n1019 B.n97 585
R120 B.n1003 B.n1002 585
R121 B.n1002 B.n93 585
R122 B.n1001 B.n92 585
R123 B.n1025 B.n92 585
R124 B.n1000 B.n91 585
R125 B.n1026 B.n91 585
R126 B.n999 B.n90 585
R127 B.n1027 B.n90 585
R128 B.n998 B.n997 585
R129 B.n997 B.n86 585
R130 B.n996 B.n85 585
R131 B.n1033 B.n85 585
R132 B.n995 B.n84 585
R133 B.n1034 B.n84 585
R134 B.n994 B.n83 585
R135 B.n1035 B.n83 585
R136 B.n993 B.n992 585
R137 B.n992 B.n79 585
R138 B.n991 B.n78 585
R139 B.n1041 B.n78 585
R140 B.n990 B.n77 585
R141 B.n1042 B.n77 585
R142 B.n989 B.n76 585
R143 B.n1043 B.n76 585
R144 B.n988 B.n987 585
R145 B.n987 B.n72 585
R146 B.n986 B.n71 585
R147 B.n1049 B.n71 585
R148 B.n985 B.n70 585
R149 B.n1050 B.n70 585
R150 B.n984 B.n69 585
R151 B.n1051 B.n69 585
R152 B.n983 B.n982 585
R153 B.n982 B.n65 585
R154 B.n981 B.n64 585
R155 B.n1057 B.n64 585
R156 B.n980 B.n63 585
R157 B.n1058 B.n63 585
R158 B.n979 B.n62 585
R159 B.n1059 B.n62 585
R160 B.n978 B.n977 585
R161 B.n977 B.n58 585
R162 B.n976 B.n57 585
R163 B.n1065 B.n57 585
R164 B.n975 B.n56 585
R165 B.n1066 B.n56 585
R166 B.n974 B.n55 585
R167 B.n1067 B.n55 585
R168 B.n973 B.n972 585
R169 B.n972 B.n51 585
R170 B.n971 B.n50 585
R171 B.n1073 B.n50 585
R172 B.n970 B.n49 585
R173 B.n1074 B.n49 585
R174 B.n969 B.n48 585
R175 B.n1075 B.n48 585
R176 B.n968 B.n967 585
R177 B.n967 B.n44 585
R178 B.n966 B.n43 585
R179 B.n1081 B.n43 585
R180 B.n965 B.n42 585
R181 B.n1082 B.n42 585
R182 B.n964 B.n41 585
R183 B.n1083 B.n41 585
R184 B.n963 B.n962 585
R185 B.n962 B.n37 585
R186 B.n961 B.n36 585
R187 B.n1089 B.n36 585
R188 B.n960 B.n35 585
R189 B.n1090 B.n35 585
R190 B.n959 B.n34 585
R191 B.n1091 B.n34 585
R192 B.n958 B.n957 585
R193 B.n957 B.n30 585
R194 B.n956 B.n29 585
R195 B.n1097 B.n29 585
R196 B.n955 B.n28 585
R197 B.n1098 B.n28 585
R198 B.n954 B.n27 585
R199 B.n1099 B.n27 585
R200 B.n953 B.n952 585
R201 B.n952 B.n23 585
R202 B.n951 B.n22 585
R203 B.n1105 B.n22 585
R204 B.n950 B.n21 585
R205 B.n1106 B.n21 585
R206 B.n949 B.n20 585
R207 B.n1107 B.n20 585
R208 B.n948 B.n947 585
R209 B.n947 B.n16 585
R210 B.n946 B.n15 585
R211 B.n1113 B.n15 585
R212 B.n945 B.n14 585
R213 B.n1114 B.n14 585
R214 B.n944 B.n13 585
R215 B.n1115 B.n13 585
R216 B.n943 B.n942 585
R217 B.n942 B.n12 585
R218 B.n941 B.n940 585
R219 B.n941 B.n8 585
R220 B.n939 B.n7 585
R221 B.n1122 B.n7 585
R222 B.n938 B.n6 585
R223 B.n1123 B.n6 585
R224 B.n937 B.n5 585
R225 B.n1124 B.n5 585
R226 B.n936 B.n935 585
R227 B.n935 B.n4 585
R228 B.n934 B.n381 585
R229 B.n934 B.n933 585
R230 B.n924 B.n382 585
R231 B.n383 B.n382 585
R232 B.n926 B.n925 585
R233 B.n927 B.n926 585
R234 B.n923 B.n388 585
R235 B.n388 B.n387 585
R236 B.n922 B.n921 585
R237 B.n921 B.n920 585
R238 B.n390 B.n389 585
R239 B.n391 B.n390 585
R240 B.n913 B.n912 585
R241 B.n914 B.n913 585
R242 B.n911 B.n396 585
R243 B.n396 B.n395 585
R244 B.n910 B.n909 585
R245 B.n909 B.n908 585
R246 B.n398 B.n397 585
R247 B.n399 B.n398 585
R248 B.n901 B.n900 585
R249 B.n902 B.n901 585
R250 B.n899 B.n403 585
R251 B.n407 B.n403 585
R252 B.n898 B.n897 585
R253 B.n897 B.n896 585
R254 B.n405 B.n404 585
R255 B.n406 B.n405 585
R256 B.n889 B.n888 585
R257 B.n890 B.n889 585
R258 B.n887 B.n412 585
R259 B.n412 B.n411 585
R260 B.n886 B.n885 585
R261 B.n885 B.n884 585
R262 B.n414 B.n413 585
R263 B.n415 B.n414 585
R264 B.n877 B.n876 585
R265 B.n878 B.n877 585
R266 B.n875 B.n419 585
R267 B.n423 B.n419 585
R268 B.n874 B.n873 585
R269 B.n873 B.n872 585
R270 B.n421 B.n420 585
R271 B.n422 B.n421 585
R272 B.n865 B.n864 585
R273 B.n866 B.n865 585
R274 B.n863 B.n428 585
R275 B.n428 B.n427 585
R276 B.n862 B.n861 585
R277 B.n861 B.n860 585
R278 B.n430 B.n429 585
R279 B.n431 B.n430 585
R280 B.n853 B.n852 585
R281 B.n854 B.n853 585
R282 B.n851 B.n435 585
R283 B.n439 B.n435 585
R284 B.n850 B.n849 585
R285 B.n849 B.n848 585
R286 B.n437 B.n436 585
R287 B.n438 B.n437 585
R288 B.n841 B.n840 585
R289 B.n842 B.n841 585
R290 B.n839 B.n444 585
R291 B.n444 B.n443 585
R292 B.n838 B.n837 585
R293 B.n837 B.n836 585
R294 B.n446 B.n445 585
R295 B.n447 B.n446 585
R296 B.n829 B.n828 585
R297 B.n830 B.n829 585
R298 B.n827 B.n451 585
R299 B.n455 B.n451 585
R300 B.n826 B.n825 585
R301 B.n825 B.n824 585
R302 B.n453 B.n452 585
R303 B.n454 B.n453 585
R304 B.n817 B.n816 585
R305 B.n818 B.n817 585
R306 B.n815 B.n460 585
R307 B.n460 B.n459 585
R308 B.n814 B.n813 585
R309 B.n813 B.n812 585
R310 B.n462 B.n461 585
R311 B.n463 B.n462 585
R312 B.n805 B.n804 585
R313 B.n806 B.n805 585
R314 B.n803 B.n468 585
R315 B.n468 B.n467 585
R316 B.n802 B.n801 585
R317 B.n801 B.n800 585
R318 B.n470 B.n469 585
R319 B.n471 B.n470 585
R320 B.n793 B.n792 585
R321 B.n794 B.n793 585
R322 B.n791 B.n476 585
R323 B.n476 B.n475 585
R324 B.n790 B.n789 585
R325 B.n789 B.n788 585
R326 B.n478 B.n477 585
R327 B.n479 B.n478 585
R328 B.n781 B.n780 585
R329 B.n782 B.n781 585
R330 B.n779 B.n484 585
R331 B.n484 B.n483 585
R332 B.n778 B.n777 585
R333 B.n777 B.n776 585
R334 B.n486 B.n485 585
R335 B.n487 B.n486 585
R336 B.n772 B.n771 585
R337 B.n490 B.n489 585
R338 B.n768 B.n767 585
R339 B.n769 B.n768 585
R340 B.n766 B.n545 585
R341 B.n765 B.n764 585
R342 B.n763 B.n762 585
R343 B.n761 B.n760 585
R344 B.n759 B.n758 585
R345 B.n757 B.n756 585
R346 B.n755 B.n754 585
R347 B.n753 B.n752 585
R348 B.n751 B.n750 585
R349 B.n749 B.n748 585
R350 B.n747 B.n746 585
R351 B.n745 B.n744 585
R352 B.n743 B.n742 585
R353 B.n741 B.n740 585
R354 B.n739 B.n738 585
R355 B.n737 B.n736 585
R356 B.n735 B.n734 585
R357 B.n733 B.n732 585
R358 B.n731 B.n730 585
R359 B.n729 B.n728 585
R360 B.n727 B.n726 585
R361 B.n725 B.n724 585
R362 B.n723 B.n722 585
R363 B.n721 B.n720 585
R364 B.n719 B.n718 585
R365 B.n717 B.n716 585
R366 B.n715 B.n714 585
R367 B.n713 B.n712 585
R368 B.n711 B.n710 585
R369 B.n709 B.n708 585
R370 B.n707 B.n706 585
R371 B.n705 B.n704 585
R372 B.n703 B.n702 585
R373 B.n701 B.n700 585
R374 B.n699 B.n698 585
R375 B.n697 B.n696 585
R376 B.n695 B.n694 585
R377 B.n693 B.n692 585
R378 B.n691 B.n690 585
R379 B.n689 B.n688 585
R380 B.n687 B.n686 585
R381 B.n685 B.n684 585
R382 B.n683 B.n682 585
R383 B.n681 B.n680 585
R384 B.n679 B.n678 585
R385 B.n677 B.n676 585
R386 B.n675 B.n674 585
R387 B.n673 B.n672 585
R388 B.n671 B.n670 585
R389 B.n669 B.n668 585
R390 B.n667 B.n666 585
R391 B.n665 B.n664 585
R392 B.n663 B.n662 585
R393 B.n661 B.n660 585
R394 B.n659 B.n658 585
R395 B.n657 B.n656 585
R396 B.n655 B.n654 585
R397 B.n652 B.n651 585
R398 B.n650 B.n649 585
R399 B.n648 B.n647 585
R400 B.n646 B.n645 585
R401 B.n644 B.n643 585
R402 B.n642 B.n641 585
R403 B.n640 B.n639 585
R404 B.n638 B.n637 585
R405 B.n636 B.n635 585
R406 B.n634 B.n633 585
R407 B.n632 B.n631 585
R408 B.n630 B.n629 585
R409 B.n628 B.n627 585
R410 B.n626 B.n625 585
R411 B.n624 B.n623 585
R412 B.n622 B.n621 585
R413 B.n620 B.n619 585
R414 B.n618 B.n617 585
R415 B.n616 B.n615 585
R416 B.n614 B.n613 585
R417 B.n612 B.n611 585
R418 B.n610 B.n609 585
R419 B.n608 B.n607 585
R420 B.n606 B.n605 585
R421 B.n604 B.n603 585
R422 B.n602 B.n601 585
R423 B.n600 B.n599 585
R424 B.n598 B.n597 585
R425 B.n596 B.n595 585
R426 B.n594 B.n593 585
R427 B.n592 B.n591 585
R428 B.n590 B.n589 585
R429 B.n588 B.n587 585
R430 B.n586 B.n585 585
R431 B.n584 B.n583 585
R432 B.n582 B.n581 585
R433 B.n580 B.n579 585
R434 B.n578 B.n577 585
R435 B.n576 B.n575 585
R436 B.n574 B.n573 585
R437 B.n572 B.n571 585
R438 B.n570 B.n569 585
R439 B.n568 B.n567 585
R440 B.n566 B.n565 585
R441 B.n564 B.n563 585
R442 B.n562 B.n561 585
R443 B.n560 B.n559 585
R444 B.n558 B.n557 585
R445 B.n556 B.n555 585
R446 B.n554 B.n553 585
R447 B.n552 B.n551 585
R448 B.n773 B.n488 585
R449 B.n488 B.n487 585
R450 B.n775 B.n774 585
R451 B.n776 B.n775 585
R452 B.n482 B.n481 585
R453 B.n483 B.n482 585
R454 B.n784 B.n783 585
R455 B.n783 B.n782 585
R456 B.n785 B.n480 585
R457 B.n480 B.n479 585
R458 B.n787 B.n786 585
R459 B.n788 B.n787 585
R460 B.n474 B.n473 585
R461 B.n475 B.n474 585
R462 B.n796 B.n795 585
R463 B.n795 B.n794 585
R464 B.n797 B.n472 585
R465 B.n472 B.n471 585
R466 B.n799 B.n798 585
R467 B.n800 B.n799 585
R468 B.n466 B.n465 585
R469 B.n467 B.n466 585
R470 B.n808 B.n807 585
R471 B.n807 B.n806 585
R472 B.n809 B.n464 585
R473 B.n464 B.n463 585
R474 B.n811 B.n810 585
R475 B.n812 B.n811 585
R476 B.n458 B.n457 585
R477 B.n459 B.n458 585
R478 B.n820 B.n819 585
R479 B.n819 B.n818 585
R480 B.n821 B.n456 585
R481 B.n456 B.n454 585
R482 B.n823 B.n822 585
R483 B.n824 B.n823 585
R484 B.n450 B.n449 585
R485 B.n455 B.n450 585
R486 B.n832 B.n831 585
R487 B.n831 B.n830 585
R488 B.n833 B.n448 585
R489 B.n448 B.n447 585
R490 B.n835 B.n834 585
R491 B.n836 B.n835 585
R492 B.n442 B.n441 585
R493 B.n443 B.n442 585
R494 B.n844 B.n843 585
R495 B.n843 B.n842 585
R496 B.n845 B.n440 585
R497 B.n440 B.n438 585
R498 B.n847 B.n846 585
R499 B.n848 B.n847 585
R500 B.n434 B.n433 585
R501 B.n439 B.n434 585
R502 B.n856 B.n855 585
R503 B.n855 B.n854 585
R504 B.n857 B.n432 585
R505 B.n432 B.n431 585
R506 B.n859 B.n858 585
R507 B.n860 B.n859 585
R508 B.n426 B.n425 585
R509 B.n427 B.n426 585
R510 B.n868 B.n867 585
R511 B.n867 B.n866 585
R512 B.n869 B.n424 585
R513 B.n424 B.n422 585
R514 B.n871 B.n870 585
R515 B.n872 B.n871 585
R516 B.n418 B.n417 585
R517 B.n423 B.n418 585
R518 B.n880 B.n879 585
R519 B.n879 B.n878 585
R520 B.n881 B.n416 585
R521 B.n416 B.n415 585
R522 B.n883 B.n882 585
R523 B.n884 B.n883 585
R524 B.n410 B.n409 585
R525 B.n411 B.n410 585
R526 B.n892 B.n891 585
R527 B.n891 B.n890 585
R528 B.n893 B.n408 585
R529 B.n408 B.n406 585
R530 B.n895 B.n894 585
R531 B.n896 B.n895 585
R532 B.n402 B.n401 585
R533 B.n407 B.n402 585
R534 B.n904 B.n903 585
R535 B.n903 B.n902 585
R536 B.n905 B.n400 585
R537 B.n400 B.n399 585
R538 B.n907 B.n906 585
R539 B.n908 B.n907 585
R540 B.n394 B.n393 585
R541 B.n395 B.n394 585
R542 B.n916 B.n915 585
R543 B.n915 B.n914 585
R544 B.n917 B.n392 585
R545 B.n392 B.n391 585
R546 B.n919 B.n918 585
R547 B.n920 B.n919 585
R548 B.n386 B.n385 585
R549 B.n387 B.n386 585
R550 B.n929 B.n928 585
R551 B.n928 B.n927 585
R552 B.n930 B.n384 585
R553 B.n384 B.n383 585
R554 B.n932 B.n931 585
R555 B.n933 B.n932 585
R556 B.n3 B.n0 585
R557 B.n4 B.n3 585
R558 B.n1121 B.n1 585
R559 B.n1122 B.n1121 585
R560 B.n1120 B.n1119 585
R561 B.n1120 B.n8 585
R562 B.n1118 B.n9 585
R563 B.n12 B.n9 585
R564 B.n1117 B.n1116 585
R565 B.n1116 B.n1115 585
R566 B.n11 B.n10 585
R567 B.n1114 B.n11 585
R568 B.n1112 B.n1111 585
R569 B.n1113 B.n1112 585
R570 B.n1110 B.n17 585
R571 B.n17 B.n16 585
R572 B.n1109 B.n1108 585
R573 B.n1108 B.n1107 585
R574 B.n19 B.n18 585
R575 B.n1106 B.n19 585
R576 B.n1104 B.n1103 585
R577 B.n1105 B.n1104 585
R578 B.n1102 B.n24 585
R579 B.n24 B.n23 585
R580 B.n1101 B.n1100 585
R581 B.n1100 B.n1099 585
R582 B.n26 B.n25 585
R583 B.n1098 B.n26 585
R584 B.n1096 B.n1095 585
R585 B.n1097 B.n1096 585
R586 B.n1094 B.n31 585
R587 B.n31 B.n30 585
R588 B.n1093 B.n1092 585
R589 B.n1092 B.n1091 585
R590 B.n33 B.n32 585
R591 B.n1090 B.n33 585
R592 B.n1088 B.n1087 585
R593 B.n1089 B.n1088 585
R594 B.n1086 B.n38 585
R595 B.n38 B.n37 585
R596 B.n1085 B.n1084 585
R597 B.n1084 B.n1083 585
R598 B.n40 B.n39 585
R599 B.n1082 B.n40 585
R600 B.n1080 B.n1079 585
R601 B.n1081 B.n1080 585
R602 B.n1078 B.n45 585
R603 B.n45 B.n44 585
R604 B.n1077 B.n1076 585
R605 B.n1076 B.n1075 585
R606 B.n47 B.n46 585
R607 B.n1074 B.n47 585
R608 B.n1072 B.n1071 585
R609 B.n1073 B.n1072 585
R610 B.n1070 B.n52 585
R611 B.n52 B.n51 585
R612 B.n1069 B.n1068 585
R613 B.n1068 B.n1067 585
R614 B.n54 B.n53 585
R615 B.n1066 B.n54 585
R616 B.n1064 B.n1063 585
R617 B.n1065 B.n1064 585
R618 B.n1062 B.n59 585
R619 B.n59 B.n58 585
R620 B.n1061 B.n1060 585
R621 B.n1060 B.n1059 585
R622 B.n61 B.n60 585
R623 B.n1058 B.n61 585
R624 B.n1056 B.n1055 585
R625 B.n1057 B.n1056 585
R626 B.n1054 B.n66 585
R627 B.n66 B.n65 585
R628 B.n1053 B.n1052 585
R629 B.n1052 B.n1051 585
R630 B.n68 B.n67 585
R631 B.n1050 B.n68 585
R632 B.n1048 B.n1047 585
R633 B.n1049 B.n1048 585
R634 B.n1046 B.n73 585
R635 B.n73 B.n72 585
R636 B.n1045 B.n1044 585
R637 B.n1044 B.n1043 585
R638 B.n75 B.n74 585
R639 B.n1042 B.n75 585
R640 B.n1040 B.n1039 585
R641 B.n1041 B.n1040 585
R642 B.n1038 B.n80 585
R643 B.n80 B.n79 585
R644 B.n1037 B.n1036 585
R645 B.n1036 B.n1035 585
R646 B.n82 B.n81 585
R647 B.n1034 B.n82 585
R648 B.n1032 B.n1031 585
R649 B.n1033 B.n1032 585
R650 B.n1030 B.n87 585
R651 B.n87 B.n86 585
R652 B.n1029 B.n1028 585
R653 B.n1028 B.n1027 585
R654 B.n89 B.n88 585
R655 B.n1026 B.n89 585
R656 B.n1024 B.n1023 585
R657 B.n1025 B.n1024 585
R658 B.n1022 B.n94 585
R659 B.n94 B.n93 585
R660 B.n1021 B.n1020 585
R661 B.n1020 B.n1019 585
R662 B.n96 B.n95 585
R663 B.n1018 B.n96 585
R664 B.n1016 B.n1015 585
R665 B.n1017 B.n1016 585
R666 B.n1014 B.n101 585
R667 B.n101 B.n100 585
R668 B.n1125 B.n1124 585
R669 B.n1123 B.n2 585
R670 B.n1012 B.n101 502.111
R671 B.n1009 B.n159 502.111
R672 B.n551 B.n486 502.111
R673 B.n771 B.n488 502.111
R674 B.n163 B.t10 362.798
R675 B.n160 B.t21 362.798
R676 B.n549 B.t18 362.798
R677 B.n546 B.t14 362.798
R678 B.n1010 B.n157 256.663
R679 B.n1010 B.n156 256.663
R680 B.n1010 B.n155 256.663
R681 B.n1010 B.n154 256.663
R682 B.n1010 B.n153 256.663
R683 B.n1010 B.n152 256.663
R684 B.n1010 B.n151 256.663
R685 B.n1010 B.n150 256.663
R686 B.n1010 B.n149 256.663
R687 B.n1010 B.n148 256.663
R688 B.n1010 B.n147 256.663
R689 B.n1010 B.n146 256.663
R690 B.n1010 B.n145 256.663
R691 B.n1010 B.n144 256.663
R692 B.n1010 B.n143 256.663
R693 B.n1010 B.n142 256.663
R694 B.n1010 B.n141 256.663
R695 B.n1010 B.n140 256.663
R696 B.n1010 B.n139 256.663
R697 B.n1010 B.n138 256.663
R698 B.n1010 B.n137 256.663
R699 B.n1010 B.n136 256.663
R700 B.n1010 B.n135 256.663
R701 B.n1010 B.n134 256.663
R702 B.n1010 B.n133 256.663
R703 B.n1010 B.n132 256.663
R704 B.n1010 B.n131 256.663
R705 B.n1010 B.n130 256.663
R706 B.n1010 B.n129 256.663
R707 B.n1010 B.n128 256.663
R708 B.n1010 B.n127 256.663
R709 B.n1010 B.n126 256.663
R710 B.n1010 B.n125 256.663
R711 B.n1010 B.n124 256.663
R712 B.n1010 B.n123 256.663
R713 B.n1010 B.n122 256.663
R714 B.n1010 B.n121 256.663
R715 B.n1010 B.n120 256.663
R716 B.n1010 B.n119 256.663
R717 B.n1010 B.n118 256.663
R718 B.n1010 B.n117 256.663
R719 B.n1010 B.n116 256.663
R720 B.n1010 B.n115 256.663
R721 B.n1010 B.n114 256.663
R722 B.n1010 B.n113 256.663
R723 B.n1010 B.n112 256.663
R724 B.n1010 B.n111 256.663
R725 B.n1010 B.n110 256.663
R726 B.n1010 B.n109 256.663
R727 B.n1010 B.n108 256.663
R728 B.n1010 B.n107 256.663
R729 B.n1010 B.n106 256.663
R730 B.n1010 B.n105 256.663
R731 B.n1010 B.n104 256.663
R732 B.n1011 B.n1010 256.663
R733 B.n770 B.n769 256.663
R734 B.n769 B.n491 256.663
R735 B.n769 B.n492 256.663
R736 B.n769 B.n493 256.663
R737 B.n769 B.n494 256.663
R738 B.n769 B.n495 256.663
R739 B.n769 B.n496 256.663
R740 B.n769 B.n497 256.663
R741 B.n769 B.n498 256.663
R742 B.n769 B.n499 256.663
R743 B.n769 B.n500 256.663
R744 B.n769 B.n501 256.663
R745 B.n769 B.n502 256.663
R746 B.n769 B.n503 256.663
R747 B.n769 B.n504 256.663
R748 B.n769 B.n505 256.663
R749 B.n769 B.n506 256.663
R750 B.n769 B.n507 256.663
R751 B.n769 B.n508 256.663
R752 B.n769 B.n509 256.663
R753 B.n769 B.n510 256.663
R754 B.n769 B.n511 256.663
R755 B.n769 B.n512 256.663
R756 B.n769 B.n513 256.663
R757 B.n769 B.n514 256.663
R758 B.n769 B.n515 256.663
R759 B.n769 B.n516 256.663
R760 B.n769 B.n517 256.663
R761 B.n769 B.n518 256.663
R762 B.n769 B.n519 256.663
R763 B.n769 B.n520 256.663
R764 B.n769 B.n521 256.663
R765 B.n769 B.n522 256.663
R766 B.n769 B.n523 256.663
R767 B.n769 B.n524 256.663
R768 B.n769 B.n525 256.663
R769 B.n769 B.n526 256.663
R770 B.n769 B.n527 256.663
R771 B.n769 B.n528 256.663
R772 B.n769 B.n529 256.663
R773 B.n769 B.n530 256.663
R774 B.n769 B.n531 256.663
R775 B.n769 B.n532 256.663
R776 B.n769 B.n533 256.663
R777 B.n769 B.n534 256.663
R778 B.n769 B.n535 256.663
R779 B.n769 B.n536 256.663
R780 B.n769 B.n537 256.663
R781 B.n769 B.n538 256.663
R782 B.n769 B.n539 256.663
R783 B.n769 B.n540 256.663
R784 B.n769 B.n541 256.663
R785 B.n769 B.n542 256.663
R786 B.n769 B.n543 256.663
R787 B.n769 B.n544 256.663
R788 B.n1127 B.n1126 256.663
R789 B.n165 B.n103 163.367
R790 B.n169 B.n168 163.367
R791 B.n173 B.n172 163.367
R792 B.n177 B.n176 163.367
R793 B.n181 B.n180 163.367
R794 B.n185 B.n184 163.367
R795 B.n189 B.n188 163.367
R796 B.n193 B.n192 163.367
R797 B.n197 B.n196 163.367
R798 B.n201 B.n200 163.367
R799 B.n205 B.n204 163.367
R800 B.n209 B.n208 163.367
R801 B.n213 B.n212 163.367
R802 B.n217 B.n216 163.367
R803 B.n221 B.n220 163.367
R804 B.n225 B.n224 163.367
R805 B.n229 B.n228 163.367
R806 B.n233 B.n232 163.367
R807 B.n237 B.n236 163.367
R808 B.n241 B.n240 163.367
R809 B.n245 B.n244 163.367
R810 B.n249 B.n248 163.367
R811 B.n253 B.n252 163.367
R812 B.n257 B.n256 163.367
R813 B.n261 B.n260 163.367
R814 B.n266 B.n265 163.367
R815 B.n270 B.n269 163.367
R816 B.n274 B.n273 163.367
R817 B.n278 B.n277 163.367
R818 B.n282 B.n281 163.367
R819 B.n286 B.n285 163.367
R820 B.n290 B.n289 163.367
R821 B.n294 B.n293 163.367
R822 B.n298 B.n297 163.367
R823 B.n302 B.n301 163.367
R824 B.n306 B.n305 163.367
R825 B.n310 B.n309 163.367
R826 B.n314 B.n313 163.367
R827 B.n318 B.n317 163.367
R828 B.n322 B.n321 163.367
R829 B.n326 B.n325 163.367
R830 B.n330 B.n329 163.367
R831 B.n334 B.n333 163.367
R832 B.n338 B.n337 163.367
R833 B.n342 B.n341 163.367
R834 B.n346 B.n345 163.367
R835 B.n350 B.n349 163.367
R836 B.n354 B.n353 163.367
R837 B.n358 B.n357 163.367
R838 B.n362 B.n361 163.367
R839 B.n366 B.n365 163.367
R840 B.n370 B.n369 163.367
R841 B.n374 B.n373 163.367
R842 B.n378 B.n377 163.367
R843 B.n1009 B.n158 163.367
R844 B.n777 B.n486 163.367
R845 B.n777 B.n484 163.367
R846 B.n781 B.n484 163.367
R847 B.n781 B.n478 163.367
R848 B.n789 B.n478 163.367
R849 B.n789 B.n476 163.367
R850 B.n793 B.n476 163.367
R851 B.n793 B.n470 163.367
R852 B.n801 B.n470 163.367
R853 B.n801 B.n468 163.367
R854 B.n805 B.n468 163.367
R855 B.n805 B.n462 163.367
R856 B.n813 B.n462 163.367
R857 B.n813 B.n460 163.367
R858 B.n817 B.n460 163.367
R859 B.n817 B.n453 163.367
R860 B.n825 B.n453 163.367
R861 B.n825 B.n451 163.367
R862 B.n829 B.n451 163.367
R863 B.n829 B.n446 163.367
R864 B.n837 B.n446 163.367
R865 B.n837 B.n444 163.367
R866 B.n841 B.n444 163.367
R867 B.n841 B.n437 163.367
R868 B.n849 B.n437 163.367
R869 B.n849 B.n435 163.367
R870 B.n853 B.n435 163.367
R871 B.n853 B.n430 163.367
R872 B.n861 B.n430 163.367
R873 B.n861 B.n428 163.367
R874 B.n865 B.n428 163.367
R875 B.n865 B.n421 163.367
R876 B.n873 B.n421 163.367
R877 B.n873 B.n419 163.367
R878 B.n877 B.n419 163.367
R879 B.n877 B.n414 163.367
R880 B.n885 B.n414 163.367
R881 B.n885 B.n412 163.367
R882 B.n889 B.n412 163.367
R883 B.n889 B.n405 163.367
R884 B.n897 B.n405 163.367
R885 B.n897 B.n403 163.367
R886 B.n901 B.n403 163.367
R887 B.n901 B.n398 163.367
R888 B.n909 B.n398 163.367
R889 B.n909 B.n396 163.367
R890 B.n913 B.n396 163.367
R891 B.n913 B.n390 163.367
R892 B.n921 B.n390 163.367
R893 B.n921 B.n388 163.367
R894 B.n926 B.n388 163.367
R895 B.n926 B.n382 163.367
R896 B.n934 B.n382 163.367
R897 B.n935 B.n934 163.367
R898 B.n935 B.n5 163.367
R899 B.n6 B.n5 163.367
R900 B.n7 B.n6 163.367
R901 B.n941 B.n7 163.367
R902 B.n942 B.n941 163.367
R903 B.n942 B.n13 163.367
R904 B.n14 B.n13 163.367
R905 B.n15 B.n14 163.367
R906 B.n947 B.n15 163.367
R907 B.n947 B.n20 163.367
R908 B.n21 B.n20 163.367
R909 B.n22 B.n21 163.367
R910 B.n952 B.n22 163.367
R911 B.n952 B.n27 163.367
R912 B.n28 B.n27 163.367
R913 B.n29 B.n28 163.367
R914 B.n957 B.n29 163.367
R915 B.n957 B.n34 163.367
R916 B.n35 B.n34 163.367
R917 B.n36 B.n35 163.367
R918 B.n962 B.n36 163.367
R919 B.n962 B.n41 163.367
R920 B.n42 B.n41 163.367
R921 B.n43 B.n42 163.367
R922 B.n967 B.n43 163.367
R923 B.n967 B.n48 163.367
R924 B.n49 B.n48 163.367
R925 B.n50 B.n49 163.367
R926 B.n972 B.n50 163.367
R927 B.n972 B.n55 163.367
R928 B.n56 B.n55 163.367
R929 B.n57 B.n56 163.367
R930 B.n977 B.n57 163.367
R931 B.n977 B.n62 163.367
R932 B.n63 B.n62 163.367
R933 B.n64 B.n63 163.367
R934 B.n982 B.n64 163.367
R935 B.n982 B.n69 163.367
R936 B.n70 B.n69 163.367
R937 B.n71 B.n70 163.367
R938 B.n987 B.n71 163.367
R939 B.n987 B.n76 163.367
R940 B.n77 B.n76 163.367
R941 B.n78 B.n77 163.367
R942 B.n992 B.n78 163.367
R943 B.n992 B.n83 163.367
R944 B.n84 B.n83 163.367
R945 B.n85 B.n84 163.367
R946 B.n997 B.n85 163.367
R947 B.n997 B.n90 163.367
R948 B.n91 B.n90 163.367
R949 B.n92 B.n91 163.367
R950 B.n1002 B.n92 163.367
R951 B.n1002 B.n97 163.367
R952 B.n98 B.n97 163.367
R953 B.n99 B.n98 163.367
R954 B.n159 B.n99 163.367
R955 B.n768 B.n490 163.367
R956 B.n768 B.n545 163.367
R957 B.n764 B.n763 163.367
R958 B.n760 B.n759 163.367
R959 B.n756 B.n755 163.367
R960 B.n752 B.n751 163.367
R961 B.n748 B.n747 163.367
R962 B.n744 B.n743 163.367
R963 B.n740 B.n739 163.367
R964 B.n736 B.n735 163.367
R965 B.n732 B.n731 163.367
R966 B.n728 B.n727 163.367
R967 B.n724 B.n723 163.367
R968 B.n720 B.n719 163.367
R969 B.n716 B.n715 163.367
R970 B.n712 B.n711 163.367
R971 B.n708 B.n707 163.367
R972 B.n704 B.n703 163.367
R973 B.n700 B.n699 163.367
R974 B.n696 B.n695 163.367
R975 B.n692 B.n691 163.367
R976 B.n688 B.n687 163.367
R977 B.n684 B.n683 163.367
R978 B.n680 B.n679 163.367
R979 B.n676 B.n675 163.367
R980 B.n672 B.n671 163.367
R981 B.n668 B.n667 163.367
R982 B.n664 B.n663 163.367
R983 B.n660 B.n659 163.367
R984 B.n656 B.n655 163.367
R985 B.n651 B.n650 163.367
R986 B.n647 B.n646 163.367
R987 B.n643 B.n642 163.367
R988 B.n639 B.n638 163.367
R989 B.n635 B.n634 163.367
R990 B.n631 B.n630 163.367
R991 B.n627 B.n626 163.367
R992 B.n623 B.n622 163.367
R993 B.n619 B.n618 163.367
R994 B.n615 B.n614 163.367
R995 B.n611 B.n610 163.367
R996 B.n607 B.n606 163.367
R997 B.n603 B.n602 163.367
R998 B.n599 B.n598 163.367
R999 B.n595 B.n594 163.367
R1000 B.n591 B.n590 163.367
R1001 B.n587 B.n586 163.367
R1002 B.n583 B.n582 163.367
R1003 B.n579 B.n578 163.367
R1004 B.n575 B.n574 163.367
R1005 B.n571 B.n570 163.367
R1006 B.n567 B.n566 163.367
R1007 B.n563 B.n562 163.367
R1008 B.n559 B.n558 163.367
R1009 B.n555 B.n554 163.367
R1010 B.n775 B.n488 163.367
R1011 B.n775 B.n482 163.367
R1012 B.n783 B.n482 163.367
R1013 B.n783 B.n480 163.367
R1014 B.n787 B.n480 163.367
R1015 B.n787 B.n474 163.367
R1016 B.n795 B.n474 163.367
R1017 B.n795 B.n472 163.367
R1018 B.n799 B.n472 163.367
R1019 B.n799 B.n466 163.367
R1020 B.n807 B.n466 163.367
R1021 B.n807 B.n464 163.367
R1022 B.n811 B.n464 163.367
R1023 B.n811 B.n458 163.367
R1024 B.n819 B.n458 163.367
R1025 B.n819 B.n456 163.367
R1026 B.n823 B.n456 163.367
R1027 B.n823 B.n450 163.367
R1028 B.n831 B.n450 163.367
R1029 B.n831 B.n448 163.367
R1030 B.n835 B.n448 163.367
R1031 B.n835 B.n442 163.367
R1032 B.n843 B.n442 163.367
R1033 B.n843 B.n440 163.367
R1034 B.n847 B.n440 163.367
R1035 B.n847 B.n434 163.367
R1036 B.n855 B.n434 163.367
R1037 B.n855 B.n432 163.367
R1038 B.n859 B.n432 163.367
R1039 B.n859 B.n426 163.367
R1040 B.n867 B.n426 163.367
R1041 B.n867 B.n424 163.367
R1042 B.n871 B.n424 163.367
R1043 B.n871 B.n418 163.367
R1044 B.n879 B.n418 163.367
R1045 B.n879 B.n416 163.367
R1046 B.n883 B.n416 163.367
R1047 B.n883 B.n410 163.367
R1048 B.n891 B.n410 163.367
R1049 B.n891 B.n408 163.367
R1050 B.n895 B.n408 163.367
R1051 B.n895 B.n402 163.367
R1052 B.n903 B.n402 163.367
R1053 B.n903 B.n400 163.367
R1054 B.n907 B.n400 163.367
R1055 B.n907 B.n394 163.367
R1056 B.n915 B.n394 163.367
R1057 B.n915 B.n392 163.367
R1058 B.n919 B.n392 163.367
R1059 B.n919 B.n386 163.367
R1060 B.n928 B.n386 163.367
R1061 B.n928 B.n384 163.367
R1062 B.n932 B.n384 163.367
R1063 B.n932 B.n3 163.367
R1064 B.n1125 B.n3 163.367
R1065 B.n1121 B.n2 163.367
R1066 B.n1121 B.n1120 163.367
R1067 B.n1120 B.n9 163.367
R1068 B.n1116 B.n9 163.367
R1069 B.n1116 B.n11 163.367
R1070 B.n1112 B.n11 163.367
R1071 B.n1112 B.n17 163.367
R1072 B.n1108 B.n17 163.367
R1073 B.n1108 B.n19 163.367
R1074 B.n1104 B.n19 163.367
R1075 B.n1104 B.n24 163.367
R1076 B.n1100 B.n24 163.367
R1077 B.n1100 B.n26 163.367
R1078 B.n1096 B.n26 163.367
R1079 B.n1096 B.n31 163.367
R1080 B.n1092 B.n31 163.367
R1081 B.n1092 B.n33 163.367
R1082 B.n1088 B.n33 163.367
R1083 B.n1088 B.n38 163.367
R1084 B.n1084 B.n38 163.367
R1085 B.n1084 B.n40 163.367
R1086 B.n1080 B.n40 163.367
R1087 B.n1080 B.n45 163.367
R1088 B.n1076 B.n45 163.367
R1089 B.n1076 B.n47 163.367
R1090 B.n1072 B.n47 163.367
R1091 B.n1072 B.n52 163.367
R1092 B.n1068 B.n52 163.367
R1093 B.n1068 B.n54 163.367
R1094 B.n1064 B.n54 163.367
R1095 B.n1064 B.n59 163.367
R1096 B.n1060 B.n59 163.367
R1097 B.n1060 B.n61 163.367
R1098 B.n1056 B.n61 163.367
R1099 B.n1056 B.n66 163.367
R1100 B.n1052 B.n66 163.367
R1101 B.n1052 B.n68 163.367
R1102 B.n1048 B.n68 163.367
R1103 B.n1048 B.n73 163.367
R1104 B.n1044 B.n73 163.367
R1105 B.n1044 B.n75 163.367
R1106 B.n1040 B.n75 163.367
R1107 B.n1040 B.n80 163.367
R1108 B.n1036 B.n80 163.367
R1109 B.n1036 B.n82 163.367
R1110 B.n1032 B.n82 163.367
R1111 B.n1032 B.n87 163.367
R1112 B.n1028 B.n87 163.367
R1113 B.n1028 B.n89 163.367
R1114 B.n1024 B.n89 163.367
R1115 B.n1024 B.n94 163.367
R1116 B.n1020 B.n94 163.367
R1117 B.n1020 B.n96 163.367
R1118 B.n1016 B.n96 163.367
R1119 B.n1016 B.n101 163.367
R1120 B.n160 B.t22 122.725
R1121 B.n549 B.t20 122.725
R1122 B.n163 B.t12 122.707
R1123 B.n546 B.t17 122.707
R1124 B.n1012 B.n1011 71.676
R1125 B.n165 B.n104 71.676
R1126 B.n169 B.n105 71.676
R1127 B.n173 B.n106 71.676
R1128 B.n177 B.n107 71.676
R1129 B.n181 B.n108 71.676
R1130 B.n185 B.n109 71.676
R1131 B.n189 B.n110 71.676
R1132 B.n193 B.n111 71.676
R1133 B.n197 B.n112 71.676
R1134 B.n201 B.n113 71.676
R1135 B.n205 B.n114 71.676
R1136 B.n209 B.n115 71.676
R1137 B.n213 B.n116 71.676
R1138 B.n217 B.n117 71.676
R1139 B.n221 B.n118 71.676
R1140 B.n225 B.n119 71.676
R1141 B.n229 B.n120 71.676
R1142 B.n233 B.n121 71.676
R1143 B.n237 B.n122 71.676
R1144 B.n241 B.n123 71.676
R1145 B.n245 B.n124 71.676
R1146 B.n249 B.n125 71.676
R1147 B.n253 B.n126 71.676
R1148 B.n257 B.n127 71.676
R1149 B.n261 B.n128 71.676
R1150 B.n266 B.n129 71.676
R1151 B.n270 B.n130 71.676
R1152 B.n274 B.n131 71.676
R1153 B.n278 B.n132 71.676
R1154 B.n282 B.n133 71.676
R1155 B.n286 B.n134 71.676
R1156 B.n290 B.n135 71.676
R1157 B.n294 B.n136 71.676
R1158 B.n298 B.n137 71.676
R1159 B.n302 B.n138 71.676
R1160 B.n306 B.n139 71.676
R1161 B.n310 B.n140 71.676
R1162 B.n314 B.n141 71.676
R1163 B.n318 B.n142 71.676
R1164 B.n322 B.n143 71.676
R1165 B.n326 B.n144 71.676
R1166 B.n330 B.n145 71.676
R1167 B.n334 B.n146 71.676
R1168 B.n338 B.n147 71.676
R1169 B.n342 B.n148 71.676
R1170 B.n346 B.n149 71.676
R1171 B.n350 B.n150 71.676
R1172 B.n354 B.n151 71.676
R1173 B.n358 B.n152 71.676
R1174 B.n362 B.n153 71.676
R1175 B.n366 B.n154 71.676
R1176 B.n370 B.n155 71.676
R1177 B.n374 B.n156 71.676
R1178 B.n378 B.n157 71.676
R1179 B.n158 B.n157 71.676
R1180 B.n377 B.n156 71.676
R1181 B.n373 B.n155 71.676
R1182 B.n369 B.n154 71.676
R1183 B.n365 B.n153 71.676
R1184 B.n361 B.n152 71.676
R1185 B.n357 B.n151 71.676
R1186 B.n353 B.n150 71.676
R1187 B.n349 B.n149 71.676
R1188 B.n345 B.n148 71.676
R1189 B.n341 B.n147 71.676
R1190 B.n337 B.n146 71.676
R1191 B.n333 B.n145 71.676
R1192 B.n329 B.n144 71.676
R1193 B.n325 B.n143 71.676
R1194 B.n321 B.n142 71.676
R1195 B.n317 B.n141 71.676
R1196 B.n313 B.n140 71.676
R1197 B.n309 B.n139 71.676
R1198 B.n305 B.n138 71.676
R1199 B.n301 B.n137 71.676
R1200 B.n297 B.n136 71.676
R1201 B.n293 B.n135 71.676
R1202 B.n289 B.n134 71.676
R1203 B.n285 B.n133 71.676
R1204 B.n281 B.n132 71.676
R1205 B.n277 B.n131 71.676
R1206 B.n273 B.n130 71.676
R1207 B.n269 B.n129 71.676
R1208 B.n265 B.n128 71.676
R1209 B.n260 B.n127 71.676
R1210 B.n256 B.n126 71.676
R1211 B.n252 B.n125 71.676
R1212 B.n248 B.n124 71.676
R1213 B.n244 B.n123 71.676
R1214 B.n240 B.n122 71.676
R1215 B.n236 B.n121 71.676
R1216 B.n232 B.n120 71.676
R1217 B.n228 B.n119 71.676
R1218 B.n224 B.n118 71.676
R1219 B.n220 B.n117 71.676
R1220 B.n216 B.n116 71.676
R1221 B.n212 B.n115 71.676
R1222 B.n208 B.n114 71.676
R1223 B.n204 B.n113 71.676
R1224 B.n200 B.n112 71.676
R1225 B.n196 B.n111 71.676
R1226 B.n192 B.n110 71.676
R1227 B.n188 B.n109 71.676
R1228 B.n184 B.n108 71.676
R1229 B.n180 B.n107 71.676
R1230 B.n176 B.n106 71.676
R1231 B.n172 B.n105 71.676
R1232 B.n168 B.n104 71.676
R1233 B.n1011 B.n103 71.676
R1234 B.n771 B.n770 71.676
R1235 B.n545 B.n491 71.676
R1236 B.n763 B.n492 71.676
R1237 B.n759 B.n493 71.676
R1238 B.n755 B.n494 71.676
R1239 B.n751 B.n495 71.676
R1240 B.n747 B.n496 71.676
R1241 B.n743 B.n497 71.676
R1242 B.n739 B.n498 71.676
R1243 B.n735 B.n499 71.676
R1244 B.n731 B.n500 71.676
R1245 B.n727 B.n501 71.676
R1246 B.n723 B.n502 71.676
R1247 B.n719 B.n503 71.676
R1248 B.n715 B.n504 71.676
R1249 B.n711 B.n505 71.676
R1250 B.n707 B.n506 71.676
R1251 B.n703 B.n507 71.676
R1252 B.n699 B.n508 71.676
R1253 B.n695 B.n509 71.676
R1254 B.n691 B.n510 71.676
R1255 B.n687 B.n511 71.676
R1256 B.n683 B.n512 71.676
R1257 B.n679 B.n513 71.676
R1258 B.n675 B.n514 71.676
R1259 B.n671 B.n515 71.676
R1260 B.n667 B.n516 71.676
R1261 B.n663 B.n517 71.676
R1262 B.n659 B.n518 71.676
R1263 B.n655 B.n519 71.676
R1264 B.n650 B.n520 71.676
R1265 B.n646 B.n521 71.676
R1266 B.n642 B.n522 71.676
R1267 B.n638 B.n523 71.676
R1268 B.n634 B.n524 71.676
R1269 B.n630 B.n525 71.676
R1270 B.n626 B.n526 71.676
R1271 B.n622 B.n527 71.676
R1272 B.n618 B.n528 71.676
R1273 B.n614 B.n529 71.676
R1274 B.n610 B.n530 71.676
R1275 B.n606 B.n531 71.676
R1276 B.n602 B.n532 71.676
R1277 B.n598 B.n533 71.676
R1278 B.n594 B.n534 71.676
R1279 B.n590 B.n535 71.676
R1280 B.n586 B.n536 71.676
R1281 B.n582 B.n537 71.676
R1282 B.n578 B.n538 71.676
R1283 B.n574 B.n539 71.676
R1284 B.n570 B.n540 71.676
R1285 B.n566 B.n541 71.676
R1286 B.n562 B.n542 71.676
R1287 B.n558 B.n543 71.676
R1288 B.n554 B.n544 71.676
R1289 B.n770 B.n490 71.676
R1290 B.n764 B.n491 71.676
R1291 B.n760 B.n492 71.676
R1292 B.n756 B.n493 71.676
R1293 B.n752 B.n494 71.676
R1294 B.n748 B.n495 71.676
R1295 B.n744 B.n496 71.676
R1296 B.n740 B.n497 71.676
R1297 B.n736 B.n498 71.676
R1298 B.n732 B.n499 71.676
R1299 B.n728 B.n500 71.676
R1300 B.n724 B.n501 71.676
R1301 B.n720 B.n502 71.676
R1302 B.n716 B.n503 71.676
R1303 B.n712 B.n504 71.676
R1304 B.n708 B.n505 71.676
R1305 B.n704 B.n506 71.676
R1306 B.n700 B.n507 71.676
R1307 B.n696 B.n508 71.676
R1308 B.n692 B.n509 71.676
R1309 B.n688 B.n510 71.676
R1310 B.n684 B.n511 71.676
R1311 B.n680 B.n512 71.676
R1312 B.n676 B.n513 71.676
R1313 B.n672 B.n514 71.676
R1314 B.n668 B.n515 71.676
R1315 B.n664 B.n516 71.676
R1316 B.n660 B.n517 71.676
R1317 B.n656 B.n518 71.676
R1318 B.n651 B.n519 71.676
R1319 B.n647 B.n520 71.676
R1320 B.n643 B.n521 71.676
R1321 B.n639 B.n522 71.676
R1322 B.n635 B.n523 71.676
R1323 B.n631 B.n524 71.676
R1324 B.n627 B.n525 71.676
R1325 B.n623 B.n526 71.676
R1326 B.n619 B.n527 71.676
R1327 B.n615 B.n528 71.676
R1328 B.n611 B.n529 71.676
R1329 B.n607 B.n530 71.676
R1330 B.n603 B.n531 71.676
R1331 B.n599 B.n532 71.676
R1332 B.n595 B.n533 71.676
R1333 B.n591 B.n534 71.676
R1334 B.n587 B.n535 71.676
R1335 B.n583 B.n536 71.676
R1336 B.n579 B.n537 71.676
R1337 B.n575 B.n538 71.676
R1338 B.n571 B.n539 71.676
R1339 B.n567 B.n540 71.676
R1340 B.n563 B.n541 71.676
R1341 B.n559 B.n542 71.676
R1342 B.n555 B.n543 71.676
R1343 B.n551 B.n544 71.676
R1344 B.n1126 B.n1125 71.676
R1345 B.n1126 B.n2 71.676
R1346 B.n161 B.t23 70.75
R1347 B.n550 B.t19 70.75
R1348 B.n164 B.t13 70.7303
R1349 B.n547 B.t16 70.7303
R1350 B.n769 B.n487 63.0733
R1351 B.n1010 B.n100 63.0733
R1352 B.n263 B.n164 59.5399
R1353 B.n162 B.n161 59.5399
R1354 B.n653 B.n550 59.5399
R1355 B.n548 B.n547 59.5399
R1356 B.n164 B.n163 51.9763
R1357 B.n161 B.n160 51.9763
R1358 B.n550 B.n549 51.9763
R1359 B.n547 B.n546 51.9763
R1360 B.n776 B.n487 36.6582
R1361 B.n776 B.n483 36.6582
R1362 B.n782 B.n483 36.6582
R1363 B.n782 B.n479 36.6582
R1364 B.n788 B.n479 36.6582
R1365 B.n788 B.n475 36.6582
R1366 B.n794 B.n475 36.6582
R1367 B.n800 B.n471 36.6582
R1368 B.n800 B.n467 36.6582
R1369 B.n806 B.n467 36.6582
R1370 B.n806 B.n463 36.6582
R1371 B.n812 B.n463 36.6582
R1372 B.n812 B.n459 36.6582
R1373 B.n818 B.n459 36.6582
R1374 B.n818 B.n454 36.6582
R1375 B.n824 B.n454 36.6582
R1376 B.n824 B.n455 36.6582
R1377 B.n830 B.n447 36.6582
R1378 B.n836 B.n447 36.6582
R1379 B.n836 B.n443 36.6582
R1380 B.n842 B.n443 36.6582
R1381 B.n842 B.n438 36.6582
R1382 B.n848 B.n438 36.6582
R1383 B.n848 B.n439 36.6582
R1384 B.n854 B.n431 36.6582
R1385 B.n860 B.n431 36.6582
R1386 B.n860 B.n427 36.6582
R1387 B.n866 B.n427 36.6582
R1388 B.n866 B.n422 36.6582
R1389 B.n872 B.n422 36.6582
R1390 B.n872 B.n423 36.6582
R1391 B.n878 B.n415 36.6582
R1392 B.n884 B.n415 36.6582
R1393 B.n884 B.n411 36.6582
R1394 B.n890 B.n411 36.6582
R1395 B.n890 B.n406 36.6582
R1396 B.n896 B.n406 36.6582
R1397 B.n896 B.n407 36.6582
R1398 B.n902 B.n399 36.6582
R1399 B.n908 B.n399 36.6582
R1400 B.n908 B.n395 36.6582
R1401 B.n914 B.n395 36.6582
R1402 B.n914 B.n391 36.6582
R1403 B.n920 B.n391 36.6582
R1404 B.n927 B.n387 36.6582
R1405 B.n927 B.n383 36.6582
R1406 B.n933 B.n383 36.6582
R1407 B.n933 B.n4 36.6582
R1408 B.n1124 B.n4 36.6582
R1409 B.n1124 B.n1123 36.6582
R1410 B.n1123 B.n1122 36.6582
R1411 B.n1122 B.n8 36.6582
R1412 B.n12 B.n8 36.6582
R1413 B.n1115 B.n12 36.6582
R1414 B.n1115 B.n1114 36.6582
R1415 B.n1113 B.n16 36.6582
R1416 B.n1107 B.n16 36.6582
R1417 B.n1107 B.n1106 36.6582
R1418 B.n1106 B.n1105 36.6582
R1419 B.n1105 B.n23 36.6582
R1420 B.n1099 B.n23 36.6582
R1421 B.n1098 B.n1097 36.6582
R1422 B.n1097 B.n30 36.6582
R1423 B.n1091 B.n30 36.6582
R1424 B.n1091 B.n1090 36.6582
R1425 B.n1090 B.n1089 36.6582
R1426 B.n1089 B.n37 36.6582
R1427 B.n1083 B.n37 36.6582
R1428 B.n1082 B.n1081 36.6582
R1429 B.n1081 B.n44 36.6582
R1430 B.n1075 B.n44 36.6582
R1431 B.n1075 B.n1074 36.6582
R1432 B.n1074 B.n1073 36.6582
R1433 B.n1073 B.n51 36.6582
R1434 B.n1067 B.n51 36.6582
R1435 B.n1066 B.n1065 36.6582
R1436 B.n1065 B.n58 36.6582
R1437 B.n1059 B.n58 36.6582
R1438 B.n1059 B.n1058 36.6582
R1439 B.n1058 B.n1057 36.6582
R1440 B.n1057 B.n65 36.6582
R1441 B.n1051 B.n65 36.6582
R1442 B.n1050 B.n1049 36.6582
R1443 B.n1049 B.n72 36.6582
R1444 B.n1043 B.n72 36.6582
R1445 B.n1043 B.n1042 36.6582
R1446 B.n1042 B.n1041 36.6582
R1447 B.n1041 B.n79 36.6582
R1448 B.n1035 B.n79 36.6582
R1449 B.n1035 B.n1034 36.6582
R1450 B.n1034 B.n1033 36.6582
R1451 B.n1033 B.n86 36.6582
R1452 B.n1027 B.n1026 36.6582
R1453 B.n1026 B.n1025 36.6582
R1454 B.n1025 B.n93 36.6582
R1455 B.n1019 B.n93 36.6582
R1456 B.n1019 B.n1018 36.6582
R1457 B.n1018 B.n1017 36.6582
R1458 B.n1017 B.n100 36.6582
R1459 B.n920 B.t2 35.0409
R1460 B.t1 B.n1113 35.0409
R1461 B.n902 B.t3 33.9628
R1462 B.n1099 B.t6 33.9628
R1463 B.n773 B.n772 32.6249
R1464 B.n552 B.n485 32.6249
R1465 B.n1008 B.n1007 32.6249
R1466 B.n1014 B.n1013 32.6249
R1467 B.n878 B.t8 29.6501
R1468 B.n1083 B.t4 29.6501
R1469 B.n854 B.t7 25.3374
R1470 B.n1067 B.t9 25.3374
R1471 B.t15 B.n471 24.2593
R1472 B.t11 B.n86 24.2593
R1473 B.n830 B.t5 21.0248
R1474 B.n1051 B.t0 21.0248
R1475 B B.n1127 18.0485
R1476 B.n455 B.t5 15.6339
R1477 B.t0 B.n1050 15.6339
R1478 B.n794 B.t15 12.3994
R1479 B.n1027 B.t11 12.3994
R1480 B.n439 B.t7 11.3213
R1481 B.t9 B.n1066 11.3213
R1482 B.n774 B.n773 10.6151
R1483 B.n774 B.n481 10.6151
R1484 B.n784 B.n481 10.6151
R1485 B.n785 B.n784 10.6151
R1486 B.n786 B.n785 10.6151
R1487 B.n786 B.n473 10.6151
R1488 B.n796 B.n473 10.6151
R1489 B.n797 B.n796 10.6151
R1490 B.n798 B.n797 10.6151
R1491 B.n798 B.n465 10.6151
R1492 B.n808 B.n465 10.6151
R1493 B.n809 B.n808 10.6151
R1494 B.n810 B.n809 10.6151
R1495 B.n810 B.n457 10.6151
R1496 B.n820 B.n457 10.6151
R1497 B.n821 B.n820 10.6151
R1498 B.n822 B.n821 10.6151
R1499 B.n822 B.n449 10.6151
R1500 B.n832 B.n449 10.6151
R1501 B.n833 B.n832 10.6151
R1502 B.n834 B.n833 10.6151
R1503 B.n834 B.n441 10.6151
R1504 B.n844 B.n441 10.6151
R1505 B.n845 B.n844 10.6151
R1506 B.n846 B.n845 10.6151
R1507 B.n846 B.n433 10.6151
R1508 B.n856 B.n433 10.6151
R1509 B.n857 B.n856 10.6151
R1510 B.n858 B.n857 10.6151
R1511 B.n858 B.n425 10.6151
R1512 B.n868 B.n425 10.6151
R1513 B.n869 B.n868 10.6151
R1514 B.n870 B.n869 10.6151
R1515 B.n870 B.n417 10.6151
R1516 B.n880 B.n417 10.6151
R1517 B.n881 B.n880 10.6151
R1518 B.n882 B.n881 10.6151
R1519 B.n882 B.n409 10.6151
R1520 B.n892 B.n409 10.6151
R1521 B.n893 B.n892 10.6151
R1522 B.n894 B.n893 10.6151
R1523 B.n894 B.n401 10.6151
R1524 B.n904 B.n401 10.6151
R1525 B.n905 B.n904 10.6151
R1526 B.n906 B.n905 10.6151
R1527 B.n906 B.n393 10.6151
R1528 B.n916 B.n393 10.6151
R1529 B.n917 B.n916 10.6151
R1530 B.n918 B.n917 10.6151
R1531 B.n918 B.n385 10.6151
R1532 B.n929 B.n385 10.6151
R1533 B.n930 B.n929 10.6151
R1534 B.n931 B.n930 10.6151
R1535 B.n931 B.n0 10.6151
R1536 B.n772 B.n489 10.6151
R1537 B.n767 B.n489 10.6151
R1538 B.n767 B.n766 10.6151
R1539 B.n766 B.n765 10.6151
R1540 B.n765 B.n762 10.6151
R1541 B.n762 B.n761 10.6151
R1542 B.n761 B.n758 10.6151
R1543 B.n758 B.n757 10.6151
R1544 B.n757 B.n754 10.6151
R1545 B.n754 B.n753 10.6151
R1546 B.n753 B.n750 10.6151
R1547 B.n750 B.n749 10.6151
R1548 B.n749 B.n746 10.6151
R1549 B.n746 B.n745 10.6151
R1550 B.n745 B.n742 10.6151
R1551 B.n742 B.n741 10.6151
R1552 B.n741 B.n738 10.6151
R1553 B.n738 B.n737 10.6151
R1554 B.n737 B.n734 10.6151
R1555 B.n734 B.n733 10.6151
R1556 B.n733 B.n730 10.6151
R1557 B.n730 B.n729 10.6151
R1558 B.n729 B.n726 10.6151
R1559 B.n726 B.n725 10.6151
R1560 B.n725 B.n722 10.6151
R1561 B.n722 B.n721 10.6151
R1562 B.n721 B.n718 10.6151
R1563 B.n718 B.n717 10.6151
R1564 B.n717 B.n714 10.6151
R1565 B.n714 B.n713 10.6151
R1566 B.n713 B.n710 10.6151
R1567 B.n710 B.n709 10.6151
R1568 B.n709 B.n706 10.6151
R1569 B.n706 B.n705 10.6151
R1570 B.n705 B.n702 10.6151
R1571 B.n702 B.n701 10.6151
R1572 B.n701 B.n698 10.6151
R1573 B.n698 B.n697 10.6151
R1574 B.n697 B.n694 10.6151
R1575 B.n694 B.n693 10.6151
R1576 B.n693 B.n690 10.6151
R1577 B.n690 B.n689 10.6151
R1578 B.n689 B.n686 10.6151
R1579 B.n686 B.n685 10.6151
R1580 B.n685 B.n682 10.6151
R1581 B.n682 B.n681 10.6151
R1582 B.n681 B.n678 10.6151
R1583 B.n678 B.n677 10.6151
R1584 B.n677 B.n674 10.6151
R1585 B.n674 B.n673 10.6151
R1586 B.n670 B.n669 10.6151
R1587 B.n669 B.n666 10.6151
R1588 B.n666 B.n665 10.6151
R1589 B.n665 B.n662 10.6151
R1590 B.n662 B.n661 10.6151
R1591 B.n661 B.n658 10.6151
R1592 B.n658 B.n657 10.6151
R1593 B.n657 B.n654 10.6151
R1594 B.n652 B.n649 10.6151
R1595 B.n649 B.n648 10.6151
R1596 B.n648 B.n645 10.6151
R1597 B.n645 B.n644 10.6151
R1598 B.n644 B.n641 10.6151
R1599 B.n641 B.n640 10.6151
R1600 B.n640 B.n637 10.6151
R1601 B.n637 B.n636 10.6151
R1602 B.n636 B.n633 10.6151
R1603 B.n633 B.n632 10.6151
R1604 B.n632 B.n629 10.6151
R1605 B.n629 B.n628 10.6151
R1606 B.n628 B.n625 10.6151
R1607 B.n625 B.n624 10.6151
R1608 B.n624 B.n621 10.6151
R1609 B.n621 B.n620 10.6151
R1610 B.n620 B.n617 10.6151
R1611 B.n617 B.n616 10.6151
R1612 B.n616 B.n613 10.6151
R1613 B.n613 B.n612 10.6151
R1614 B.n612 B.n609 10.6151
R1615 B.n609 B.n608 10.6151
R1616 B.n608 B.n605 10.6151
R1617 B.n605 B.n604 10.6151
R1618 B.n604 B.n601 10.6151
R1619 B.n601 B.n600 10.6151
R1620 B.n600 B.n597 10.6151
R1621 B.n597 B.n596 10.6151
R1622 B.n596 B.n593 10.6151
R1623 B.n593 B.n592 10.6151
R1624 B.n592 B.n589 10.6151
R1625 B.n589 B.n588 10.6151
R1626 B.n588 B.n585 10.6151
R1627 B.n585 B.n584 10.6151
R1628 B.n584 B.n581 10.6151
R1629 B.n581 B.n580 10.6151
R1630 B.n580 B.n577 10.6151
R1631 B.n577 B.n576 10.6151
R1632 B.n576 B.n573 10.6151
R1633 B.n573 B.n572 10.6151
R1634 B.n572 B.n569 10.6151
R1635 B.n569 B.n568 10.6151
R1636 B.n568 B.n565 10.6151
R1637 B.n565 B.n564 10.6151
R1638 B.n564 B.n561 10.6151
R1639 B.n561 B.n560 10.6151
R1640 B.n560 B.n557 10.6151
R1641 B.n557 B.n556 10.6151
R1642 B.n556 B.n553 10.6151
R1643 B.n553 B.n552 10.6151
R1644 B.n778 B.n485 10.6151
R1645 B.n779 B.n778 10.6151
R1646 B.n780 B.n779 10.6151
R1647 B.n780 B.n477 10.6151
R1648 B.n790 B.n477 10.6151
R1649 B.n791 B.n790 10.6151
R1650 B.n792 B.n791 10.6151
R1651 B.n792 B.n469 10.6151
R1652 B.n802 B.n469 10.6151
R1653 B.n803 B.n802 10.6151
R1654 B.n804 B.n803 10.6151
R1655 B.n804 B.n461 10.6151
R1656 B.n814 B.n461 10.6151
R1657 B.n815 B.n814 10.6151
R1658 B.n816 B.n815 10.6151
R1659 B.n816 B.n452 10.6151
R1660 B.n826 B.n452 10.6151
R1661 B.n827 B.n826 10.6151
R1662 B.n828 B.n827 10.6151
R1663 B.n828 B.n445 10.6151
R1664 B.n838 B.n445 10.6151
R1665 B.n839 B.n838 10.6151
R1666 B.n840 B.n839 10.6151
R1667 B.n840 B.n436 10.6151
R1668 B.n850 B.n436 10.6151
R1669 B.n851 B.n850 10.6151
R1670 B.n852 B.n851 10.6151
R1671 B.n852 B.n429 10.6151
R1672 B.n862 B.n429 10.6151
R1673 B.n863 B.n862 10.6151
R1674 B.n864 B.n863 10.6151
R1675 B.n864 B.n420 10.6151
R1676 B.n874 B.n420 10.6151
R1677 B.n875 B.n874 10.6151
R1678 B.n876 B.n875 10.6151
R1679 B.n876 B.n413 10.6151
R1680 B.n886 B.n413 10.6151
R1681 B.n887 B.n886 10.6151
R1682 B.n888 B.n887 10.6151
R1683 B.n888 B.n404 10.6151
R1684 B.n898 B.n404 10.6151
R1685 B.n899 B.n898 10.6151
R1686 B.n900 B.n899 10.6151
R1687 B.n900 B.n397 10.6151
R1688 B.n910 B.n397 10.6151
R1689 B.n911 B.n910 10.6151
R1690 B.n912 B.n911 10.6151
R1691 B.n912 B.n389 10.6151
R1692 B.n922 B.n389 10.6151
R1693 B.n923 B.n922 10.6151
R1694 B.n925 B.n923 10.6151
R1695 B.n925 B.n924 10.6151
R1696 B.n924 B.n381 10.6151
R1697 B.n936 B.n381 10.6151
R1698 B.n937 B.n936 10.6151
R1699 B.n938 B.n937 10.6151
R1700 B.n939 B.n938 10.6151
R1701 B.n940 B.n939 10.6151
R1702 B.n943 B.n940 10.6151
R1703 B.n944 B.n943 10.6151
R1704 B.n945 B.n944 10.6151
R1705 B.n946 B.n945 10.6151
R1706 B.n948 B.n946 10.6151
R1707 B.n949 B.n948 10.6151
R1708 B.n950 B.n949 10.6151
R1709 B.n951 B.n950 10.6151
R1710 B.n953 B.n951 10.6151
R1711 B.n954 B.n953 10.6151
R1712 B.n955 B.n954 10.6151
R1713 B.n956 B.n955 10.6151
R1714 B.n958 B.n956 10.6151
R1715 B.n959 B.n958 10.6151
R1716 B.n960 B.n959 10.6151
R1717 B.n961 B.n960 10.6151
R1718 B.n963 B.n961 10.6151
R1719 B.n964 B.n963 10.6151
R1720 B.n965 B.n964 10.6151
R1721 B.n966 B.n965 10.6151
R1722 B.n968 B.n966 10.6151
R1723 B.n969 B.n968 10.6151
R1724 B.n970 B.n969 10.6151
R1725 B.n971 B.n970 10.6151
R1726 B.n973 B.n971 10.6151
R1727 B.n974 B.n973 10.6151
R1728 B.n975 B.n974 10.6151
R1729 B.n976 B.n975 10.6151
R1730 B.n978 B.n976 10.6151
R1731 B.n979 B.n978 10.6151
R1732 B.n980 B.n979 10.6151
R1733 B.n981 B.n980 10.6151
R1734 B.n983 B.n981 10.6151
R1735 B.n984 B.n983 10.6151
R1736 B.n985 B.n984 10.6151
R1737 B.n986 B.n985 10.6151
R1738 B.n988 B.n986 10.6151
R1739 B.n989 B.n988 10.6151
R1740 B.n990 B.n989 10.6151
R1741 B.n991 B.n990 10.6151
R1742 B.n993 B.n991 10.6151
R1743 B.n994 B.n993 10.6151
R1744 B.n995 B.n994 10.6151
R1745 B.n996 B.n995 10.6151
R1746 B.n998 B.n996 10.6151
R1747 B.n999 B.n998 10.6151
R1748 B.n1000 B.n999 10.6151
R1749 B.n1001 B.n1000 10.6151
R1750 B.n1003 B.n1001 10.6151
R1751 B.n1004 B.n1003 10.6151
R1752 B.n1005 B.n1004 10.6151
R1753 B.n1006 B.n1005 10.6151
R1754 B.n1007 B.n1006 10.6151
R1755 B.n1119 B.n1 10.6151
R1756 B.n1119 B.n1118 10.6151
R1757 B.n1118 B.n1117 10.6151
R1758 B.n1117 B.n10 10.6151
R1759 B.n1111 B.n10 10.6151
R1760 B.n1111 B.n1110 10.6151
R1761 B.n1110 B.n1109 10.6151
R1762 B.n1109 B.n18 10.6151
R1763 B.n1103 B.n18 10.6151
R1764 B.n1103 B.n1102 10.6151
R1765 B.n1102 B.n1101 10.6151
R1766 B.n1101 B.n25 10.6151
R1767 B.n1095 B.n25 10.6151
R1768 B.n1095 B.n1094 10.6151
R1769 B.n1094 B.n1093 10.6151
R1770 B.n1093 B.n32 10.6151
R1771 B.n1087 B.n32 10.6151
R1772 B.n1087 B.n1086 10.6151
R1773 B.n1086 B.n1085 10.6151
R1774 B.n1085 B.n39 10.6151
R1775 B.n1079 B.n39 10.6151
R1776 B.n1079 B.n1078 10.6151
R1777 B.n1078 B.n1077 10.6151
R1778 B.n1077 B.n46 10.6151
R1779 B.n1071 B.n46 10.6151
R1780 B.n1071 B.n1070 10.6151
R1781 B.n1070 B.n1069 10.6151
R1782 B.n1069 B.n53 10.6151
R1783 B.n1063 B.n53 10.6151
R1784 B.n1063 B.n1062 10.6151
R1785 B.n1062 B.n1061 10.6151
R1786 B.n1061 B.n60 10.6151
R1787 B.n1055 B.n60 10.6151
R1788 B.n1055 B.n1054 10.6151
R1789 B.n1054 B.n1053 10.6151
R1790 B.n1053 B.n67 10.6151
R1791 B.n1047 B.n67 10.6151
R1792 B.n1047 B.n1046 10.6151
R1793 B.n1046 B.n1045 10.6151
R1794 B.n1045 B.n74 10.6151
R1795 B.n1039 B.n74 10.6151
R1796 B.n1039 B.n1038 10.6151
R1797 B.n1038 B.n1037 10.6151
R1798 B.n1037 B.n81 10.6151
R1799 B.n1031 B.n81 10.6151
R1800 B.n1031 B.n1030 10.6151
R1801 B.n1030 B.n1029 10.6151
R1802 B.n1029 B.n88 10.6151
R1803 B.n1023 B.n88 10.6151
R1804 B.n1023 B.n1022 10.6151
R1805 B.n1022 B.n1021 10.6151
R1806 B.n1021 B.n95 10.6151
R1807 B.n1015 B.n95 10.6151
R1808 B.n1015 B.n1014 10.6151
R1809 B.n1013 B.n102 10.6151
R1810 B.n166 B.n102 10.6151
R1811 B.n167 B.n166 10.6151
R1812 B.n170 B.n167 10.6151
R1813 B.n171 B.n170 10.6151
R1814 B.n174 B.n171 10.6151
R1815 B.n175 B.n174 10.6151
R1816 B.n178 B.n175 10.6151
R1817 B.n179 B.n178 10.6151
R1818 B.n182 B.n179 10.6151
R1819 B.n183 B.n182 10.6151
R1820 B.n186 B.n183 10.6151
R1821 B.n187 B.n186 10.6151
R1822 B.n190 B.n187 10.6151
R1823 B.n191 B.n190 10.6151
R1824 B.n194 B.n191 10.6151
R1825 B.n195 B.n194 10.6151
R1826 B.n198 B.n195 10.6151
R1827 B.n199 B.n198 10.6151
R1828 B.n202 B.n199 10.6151
R1829 B.n203 B.n202 10.6151
R1830 B.n206 B.n203 10.6151
R1831 B.n207 B.n206 10.6151
R1832 B.n210 B.n207 10.6151
R1833 B.n211 B.n210 10.6151
R1834 B.n214 B.n211 10.6151
R1835 B.n215 B.n214 10.6151
R1836 B.n218 B.n215 10.6151
R1837 B.n219 B.n218 10.6151
R1838 B.n222 B.n219 10.6151
R1839 B.n223 B.n222 10.6151
R1840 B.n226 B.n223 10.6151
R1841 B.n227 B.n226 10.6151
R1842 B.n230 B.n227 10.6151
R1843 B.n231 B.n230 10.6151
R1844 B.n234 B.n231 10.6151
R1845 B.n235 B.n234 10.6151
R1846 B.n238 B.n235 10.6151
R1847 B.n239 B.n238 10.6151
R1848 B.n242 B.n239 10.6151
R1849 B.n243 B.n242 10.6151
R1850 B.n246 B.n243 10.6151
R1851 B.n247 B.n246 10.6151
R1852 B.n250 B.n247 10.6151
R1853 B.n251 B.n250 10.6151
R1854 B.n254 B.n251 10.6151
R1855 B.n255 B.n254 10.6151
R1856 B.n258 B.n255 10.6151
R1857 B.n259 B.n258 10.6151
R1858 B.n262 B.n259 10.6151
R1859 B.n267 B.n264 10.6151
R1860 B.n268 B.n267 10.6151
R1861 B.n271 B.n268 10.6151
R1862 B.n272 B.n271 10.6151
R1863 B.n275 B.n272 10.6151
R1864 B.n276 B.n275 10.6151
R1865 B.n279 B.n276 10.6151
R1866 B.n280 B.n279 10.6151
R1867 B.n284 B.n283 10.6151
R1868 B.n287 B.n284 10.6151
R1869 B.n288 B.n287 10.6151
R1870 B.n291 B.n288 10.6151
R1871 B.n292 B.n291 10.6151
R1872 B.n295 B.n292 10.6151
R1873 B.n296 B.n295 10.6151
R1874 B.n299 B.n296 10.6151
R1875 B.n300 B.n299 10.6151
R1876 B.n303 B.n300 10.6151
R1877 B.n304 B.n303 10.6151
R1878 B.n307 B.n304 10.6151
R1879 B.n308 B.n307 10.6151
R1880 B.n311 B.n308 10.6151
R1881 B.n312 B.n311 10.6151
R1882 B.n315 B.n312 10.6151
R1883 B.n316 B.n315 10.6151
R1884 B.n319 B.n316 10.6151
R1885 B.n320 B.n319 10.6151
R1886 B.n323 B.n320 10.6151
R1887 B.n324 B.n323 10.6151
R1888 B.n327 B.n324 10.6151
R1889 B.n328 B.n327 10.6151
R1890 B.n331 B.n328 10.6151
R1891 B.n332 B.n331 10.6151
R1892 B.n335 B.n332 10.6151
R1893 B.n336 B.n335 10.6151
R1894 B.n339 B.n336 10.6151
R1895 B.n340 B.n339 10.6151
R1896 B.n343 B.n340 10.6151
R1897 B.n344 B.n343 10.6151
R1898 B.n347 B.n344 10.6151
R1899 B.n348 B.n347 10.6151
R1900 B.n351 B.n348 10.6151
R1901 B.n352 B.n351 10.6151
R1902 B.n355 B.n352 10.6151
R1903 B.n356 B.n355 10.6151
R1904 B.n359 B.n356 10.6151
R1905 B.n360 B.n359 10.6151
R1906 B.n363 B.n360 10.6151
R1907 B.n364 B.n363 10.6151
R1908 B.n367 B.n364 10.6151
R1909 B.n368 B.n367 10.6151
R1910 B.n371 B.n368 10.6151
R1911 B.n372 B.n371 10.6151
R1912 B.n375 B.n372 10.6151
R1913 B.n376 B.n375 10.6151
R1914 B.n379 B.n376 10.6151
R1915 B.n380 B.n379 10.6151
R1916 B.n1008 B.n380 10.6151
R1917 B.n1127 B.n0 8.11757
R1918 B.n1127 B.n1 8.11757
R1919 B.n423 B.t8 7.00859
R1920 B.t4 B.n1082 7.00859
R1921 B.n670 B.n548 6.5566
R1922 B.n654 B.n653 6.5566
R1923 B.n264 B.n263 6.5566
R1924 B.n280 B.n162 6.5566
R1925 B.n673 B.n548 4.05904
R1926 B.n653 B.n652 4.05904
R1927 B.n263 B.n262 4.05904
R1928 B.n283 B.n162 4.05904
R1929 B.n407 B.t3 2.69592
R1930 B.t6 B.n1098 2.69592
R1931 B.t2 B.n387 1.61775
R1932 B.n1114 B.t1 1.61775
R1933 VP.n19 VP.t8 188.483
R1934 VP.n22 VP.n21 161.3
R1935 VP.n23 VP.n18 161.3
R1936 VP.n25 VP.n24 161.3
R1937 VP.n26 VP.n17 161.3
R1938 VP.n28 VP.n27 161.3
R1939 VP.n29 VP.n16 161.3
R1940 VP.n31 VP.n30 161.3
R1941 VP.n32 VP.n15 161.3
R1942 VP.n34 VP.n33 161.3
R1943 VP.n35 VP.n14 161.3
R1944 VP.n37 VP.n36 161.3
R1945 VP.n39 VP.n13 161.3
R1946 VP.n41 VP.n40 161.3
R1947 VP.n42 VP.n12 161.3
R1948 VP.n44 VP.n43 161.3
R1949 VP.n45 VP.n11 161.3
R1950 VP.n82 VP.n0 161.3
R1951 VP.n81 VP.n80 161.3
R1952 VP.n79 VP.n1 161.3
R1953 VP.n78 VP.n77 161.3
R1954 VP.n76 VP.n2 161.3
R1955 VP.n74 VP.n73 161.3
R1956 VP.n72 VP.n3 161.3
R1957 VP.n71 VP.n70 161.3
R1958 VP.n69 VP.n4 161.3
R1959 VP.n68 VP.n67 161.3
R1960 VP.n66 VP.n5 161.3
R1961 VP.n65 VP.n64 161.3
R1962 VP.n63 VP.n6 161.3
R1963 VP.n62 VP.n61 161.3
R1964 VP.n60 VP.n7 161.3
R1965 VP.n59 VP.n58 161.3
R1966 VP.n56 VP.n8 161.3
R1967 VP.n55 VP.n54 161.3
R1968 VP.n53 VP.n9 161.3
R1969 VP.n52 VP.n51 161.3
R1970 VP.n50 VP.n10 161.3
R1971 VP.n5 VP.t4 155.163
R1972 VP.n49 VP.t1 155.163
R1973 VP.n57 VP.t2 155.163
R1974 VP.n75 VP.t7 155.163
R1975 VP.n83 VP.t6 155.163
R1976 VP.n16 VP.t3 155.163
R1977 VP.n46 VP.t9 155.163
R1978 VP.n38 VP.t0 155.163
R1979 VP.n20 VP.t5 155.163
R1980 VP.n49 VP.n48 93.1402
R1981 VP.n84 VP.n83 93.1402
R1982 VP.n47 VP.n46 93.1402
R1983 VP.n20 VP.n19 63.0043
R1984 VP.n63 VP.n62 56.0336
R1985 VP.n70 VP.n69 56.0336
R1986 VP.n33 VP.n32 56.0336
R1987 VP.n26 VP.n25 56.0336
R1988 VP.n48 VP.n47 54.2041
R1989 VP.n51 VP.n9 42.4359
R1990 VP.n81 VP.n1 42.4359
R1991 VP.n44 VP.n12 42.4359
R1992 VP.n55 VP.n9 38.5509
R1993 VP.n77 VP.n1 38.5509
R1994 VP.n40 VP.n12 38.5509
R1995 VP.n62 VP.n7 24.9531
R1996 VP.n70 VP.n3 24.9531
R1997 VP.n33 VP.n14 24.9531
R1998 VP.n25 VP.n18 24.9531
R1999 VP.n51 VP.n50 24.4675
R2000 VP.n56 VP.n55 24.4675
R2001 VP.n58 VP.n7 24.4675
R2002 VP.n64 VP.n63 24.4675
R2003 VP.n64 VP.n5 24.4675
R2004 VP.n68 VP.n5 24.4675
R2005 VP.n69 VP.n68 24.4675
R2006 VP.n74 VP.n3 24.4675
R2007 VP.n77 VP.n76 24.4675
R2008 VP.n82 VP.n81 24.4675
R2009 VP.n45 VP.n44 24.4675
R2010 VP.n37 VP.n14 24.4675
R2011 VP.n40 VP.n39 24.4675
R2012 VP.n27 VP.n26 24.4675
R2013 VP.n27 VP.n16 24.4675
R2014 VP.n31 VP.n16 24.4675
R2015 VP.n32 VP.n31 24.4675
R2016 VP.n21 VP.n18 24.4675
R2017 VP.n50 VP.n49 17.6167
R2018 VP.n83 VP.n82 17.6167
R2019 VP.n46 VP.n45 17.6167
R2020 VP.n57 VP.n56 15.6594
R2021 VP.n76 VP.n75 15.6594
R2022 VP.n39 VP.n38 15.6594
R2023 VP.n22 VP.n19 9.21387
R2024 VP.n58 VP.n57 8.80862
R2025 VP.n75 VP.n74 8.80862
R2026 VP.n38 VP.n37 8.80862
R2027 VP.n21 VP.n20 8.80862
R2028 VP.n47 VP.n11 0.278367
R2029 VP.n48 VP.n10 0.278367
R2030 VP.n84 VP.n0 0.278367
R2031 VP.n23 VP.n22 0.189894
R2032 VP.n24 VP.n23 0.189894
R2033 VP.n24 VP.n17 0.189894
R2034 VP.n28 VP.n17 0.189894
R2035 VP.n29 VP.n28 0.189894
R2036 VP.n30 VP.n29 0.189894
R2037 VP.n30 VP.n15 0.189894
R2038 VP.n34 VP.n15 0.189894
R2039 VP.n35 VP.n34 0.189894
R2040 VP.n36 VP.n35 0.189894
R2041 VP.n36 VP.n13 0.189894
R2042 VP.n41 VP.n13 0.189894
R2043 VP.n42 VP.n41 0.189894
R2044 VP.n43 VP.n42 0.189894
R2045 VP.n43 VP.n11 0.189894
R2046 VP.n52 VP.n10 0.189894
R2047 VP.n53 VP.n52 0.189894
R2048 VP.n54 VP.n53 0.189894
R2049 VP.n54 VP.n8 0.189894
R2050 VP.n59 VP.n8 0.189894
R2051 VP.n60 VP.n59 0.189894
R2052 VP.n61 VP.n60 0.189894
R2053 VP.n61 VP.n6 0.189894
R2054 VP.n65 VP.n6 0.189894
R2055 VP.n66 VP.n65 0.189894
R2056 VP.n67 VP.n66 0.189894
R2057 VP.n67 VP.n4 0.189894
R2058 VP.n71 VP.n4 0.189894
R2059 VP.n72 VP.n71 0.189894
R2060 VP.n73 VP.n72 0.189894
R2061 VP.n73 VP.n2 0.189894
R2062 VP.n78 VP.n2 0.189894
R2063 VP.n79 VP.n78 0.189894
R2064 VP.n80 VP.n79 0.189894
R2065 VP.n80 VP.n0 0.189894
R2066 VP VP.n84 0.153454
R2067 VDD1.n1 VDD1.t2 67.02
R2068 VDD1.n3 VDD1.t1 67.0198
R2069 VDD1.n5 VDD1.n4 65.0782
R2070 VDD1.n1 VDD1.n0 63.401
R2071 VDD1.n7 VDD1.n6 63.4008
R2072 VDD1.n3 VDD1.n2 63.4008
R2073 VDD1.n7 VDD1.n5 49.4707
R2074 VDD1 VDD1.n7 1.67507
R2075 VDD1.n6 VDD1.t3 1.30916
R2076 VDD1.n6 VDD1.t7 1.30916
R2077 VDD1.n0 VDD1.t4 1.30916
R2078 VDD1.n0 VDD1.t6 1.30916
R2079 VDD1.n4 VDD1.t0 1.30916
R2080 VDD1.n4 VDD1.t9 1.30916
R2081 VDD1.n2 VDD1.t8 1.30916
R2082 VDD1.n2 VDD1.t5 1.30916
R2083 VDD1 VDD1.n1 0.636276
R2084 VDD1.n5 VDD1.n3 0.52274
R2085 VTAIL.n11 VTAIL.t19 48.0309
R2086 VTAIL.n17 VTAIL.t0 48.0306
R2087 VTAIL.n2 VTAIL.t12 48.0306
R2088 VTAIL.n16 VTAIL.t9 48.0306
R2089 VTAIL.n15 VTAIL.n14 46.7222
R2090 VTAIL.n13 VTAIL.n12 46.7222
R2091 VTAIL.n10 VTAIL.n9 46.7222
R2092 VTAIL.n8 VTAIL.n7 46.7222
R2093 VTAIL.n19 VTAIL.n18 46.722
R2094 VTAIL.n1 VTAIL.n0 46.722
R2095 VTAIL.n4 VTAIL.n3 46.722
R2096 VTAIL.n6 VTAIL.n5 46.722
R2097 VTAIL.n8 VTAIL.n6 30.0307
R2098 VTAIL.n17 VTAIL.n16 27.7203
R2099 VTAIL.n10 VTAIL.n8 2.31084
R2100 VTAIL.n11 VTAIL.n10 2.31084
R2101 VTAIL.n15 VTAIL.n13 2.31084
R2102 VTAIL.n16 VTAIL.n15 2.31084
R2103 VTAIL.n6 VTAIL.n4 2.31084
R2104 VTAIL.n4 VTAIL.n2 2.31084
R2105 VTAIL.n19 VTAIL.n17 2.31084
R2106 VTAIL VTAIL.n1 1.79145
R2107 VTAIL.n13 VTAIL.n11 1.6255
R2108 VTAIL.n2 VTAIL.n1 1.6255
R2109 VTAIL.n18 VTAIL.t2 1.30916
R2110 VTAIL.n18 VTAIL.t7 1.30916
R2111 VTAIL.n0 VTAIL.t1 1.30916
R2112 VTAIL.n0 VTAIL.t8 1.30916
R2113 VTAIL.n3 VTAIL.t14 1.30916
R2114 VTAIL.n3 VTAIL.t11 1.30916
R2115 VTAIL.n5 VTAIL.t17 1.30916
R2116 VTAIL.n5 VTAIL.t16 1.30916
R2117 VTAIL.n14 VTAIL.t15 1.30916
R2118 VTAIL.n14 VTAIL.t18 1.30916
R2119 VTAIL.n12 VTAIL.t10 1.30916
R2120 VTAIL.n12 VTAIL.t13 1.30916
R2121 VTAIL.n9 VTAIL.t4 1.30916
R2122 VTAIL.n9 VTAIL.t5 1.30916
R2123 VTAIL.n7 VTAIL.t3 1.30916
R2124 VTAIL.n7 VTAIL.t6 1.30916
R2125 VTAIL VTAIL.n19 0.519897
R2126 VN.n8 VN.t1 188.483
R2127 VN.n45 VN.t6 188.483
R2128 VN.n71 VN.n37 161.3
R2129 VN.n70 VN.n69 161.3
R2130 VN.n68 VN.n38 161.3
R2131 VN.n67 VN.n66 161.3
R2132 VN.n65 VN.n39 161.3
R2133 VN.n63 VN.n62 161.3
R2134 VN.n61 VN.n40 161.3
R2135 VN.n60 VN.n59 161.3
R2136 VN.n58 VN.n41 161.3
R2137 VN.n57 VN.n56 161.3
R2138 VN.n55 VN.n42 161.3
R2139 VN.n54 VN.n53 161.3
R2140 VN.n52 VN.n43 161.3
R2141 VN.n51 VN.n50 161.3
R2142 VN.n49 VN.n44 161.3
R2143 VN.n48 VN.n47 161.3
R2144 VN.n34 VN.n0 161.3
R2145 VN.n33 VN.n32 161.3
R2146 VN.n31 VN.n1 161.3
R2147 VN.n30 VN.n29 161.3
R2148 VN.n28 VN.n2 161.3
R2149 VN.n26 VN.n25 161.3
R2150 VN.n24 VN.n3 161.3
R2151 VN.n23 VN.n22 161.3
R2152 VN.n21 VN.n4 161.3
R2153 VN.n20 VN.n19 161.3
R2154 VN.n18 VN.n5 161.3
R2155 VN.n17 VN.n16 161.3
R2156 VN.n15 VN.n6 161.3
R2157 VN.n14 VN.n13 161.3
R2158 VN.n12 VN.n7 161.3
R2159 VN.n11 VN.n10 161.3
R2160 VN.n5 VN.t9 155.163
R2161 VN.n9 VN.t0 155.163
R2162 VN.n27 VN.t2 155.163
R2163 VN.n35 VN.t8 155.163
R2164 VN.n42 VN.t5 155.163
R2165 VN.n46 VN.t4 155.163
R2166 VN.n64 VN.t3 155.163
R2167 VN.n72 VN.t7 155.163
R2168 VN.n36 VN.n35 93.1402
R2169 VN.n73 VN.n72 93.1402
R2170 VN.n9 VN.n8 63.0043
R2171 VN.n46 VN.n45 63.0043
R2172 VN.n15 VN.n14 56.0336
R2173 VN.n22 VN.n21 56.0336
R2174 VN.n52 VN.n51 56.0336
R2175 VN.n59 VN.n58 56.0336
R2176 VN VN.n73 54.483
R2177 VN.n33 VN.n1 42.4359
R2178 VN.n70 VN.n38 42.4359
R2179 VN.n29 VN.n1 38.5509
R2180 VN.n66 VN.n38 38.5509
R2181 VN.n14 VN.n7 24.9531
R2182 VN.n22 VN.n3 24.9531
R2183 VN.n51 VN.n44 24.9531
R2184 VN.n59 VN.n40 24.9531
R2185 VN.n10 VN.n7 24.4675
R2186 VN.n16 VN.n15 24.4675
R2187 VN.n16 VN.n5 24.4675
R2188 VN.n20 VN.n5 24.4675
R2189 VN.n21 VN.n20 24.4675
R2190 VN.n26 VN.n3 24.4675
R2191 VN.n29 VN.n28 24.4675
R2192 VN.n34 VN.n33 24.4675
R2193 VN.n47 VN.n44 24.4675
R2194 VN.n58 VN.n57 24.4675
R2195 VN.n57 VN.n42 24.4675
R2196 VN.n53 VN.n42 24.4675
R2197 VN.n53 VN.n52 24.4675
R2198 VN.n66 VN.n65 24.4675
R2199 VN.n63 VN.n40 24.4675
R2200 VN.n71 VN.n70 24.4675
R2201 VN.n35 VN.n34 17.6167
R2202 VN.n72 VN.n71 17.6167
R2203 VN.n28 VN.n27 15.6594
R2204 VN.n65 VN.n64 15.6594
R2205 VN.n48 VN.n45 9.21387
R2206 VN.n11 VN.n8 9.21387
R2207 VN.n10 VN.n9 8.80862
R2208 VN.n27 VN.n26 8.80862
R2209 VN.n47 VN.n46 8.80862
R2210 VN.n64 VN.n63 8.80862
R2211 VN.n73 VN.n37 0.278367
R2212 VN.n36 VN.n0 0.278367
R2213 VN.n69 VN.n37 0.189894
R2214 VN.n69 VN.n68 0.189894
R2215 VN.n68 VN.n67 0.189894
R2216 VN.n67 VN.n39 0.189894
R2217 VN.n62 VN.n39 0.189894
R2218 VN.n62 VN.n61 0.189894
R2219 VN.n61 VN.n60 0.189894
R2220 VN.n60 VN.n41 0.189894
R2221 VN.n56 VN.n41 0.189894
R2222 VN.n56 VN.n55 0.189894
R2223 VN.n55 VN.n54 0.189894
R2224 VN.n54 VN.n43 0.189894
R2225 VN.n50 VN.n43 0.189894
R2226 VN.n50 VN.n49 0.189894
R2227 VN.n49 VN.n48 0.189894
R2228 VN.n12 VN.n11 0.189894
R2229 VN.n13 VN.n12 0.189894
R2230 VN.n13 VN.n6 0.189894
R2231 VN.n17 VN.n6 0.189894
R2232 VN.n18 VN.n17 0.189894
R2233 VN.n19 VN.n18 0.189894
R2234 VN.n19 VN.n4 0.189894
R2235 VN.n23 VN.n4 0.189894
R2236 VN.n24 VN.n23 0.189894
R2237 VN.n25 VN.n24 0.189894
R2238 VN.n25 VN.n2 0.189894
R2239 VN.n30 VN.n2 0.189894
R2240 VN.n31 VN.n30 0.189894
R2241 VN.n32 VN.n31 0.189894
R2242 VN.n32 VN.n0 0.189894
R2243 VN VN.n36 0.153454
R2244 VDD2.n1 VDD2.t8 67.0198
R2245 VDD2.n3 VDD2.n2 65.0782
R2246 VDD2 VDD2.n7 65.0754
R2247 VDD2.n4 VDD2.t2 64.7097
R2248 VDD2.n6 VDD2.n5 63.401
R2249 VDD2.n1 VDD2.n0 63.4008
R2250 VDD2.n4 VDD2.n3 47.7325
R2251 VDD2.n6 VDD2.n4 2.31084
R2252 VDD2.n7 VDD2.t5 1.30916
R2253 VDD2.n7 VDD2.t3 1.30916
R2254 VDD2.n5 VDD2.t6 1.30916
R2255 VDD2.n5 VDD2.t4 1.30916
R2256 VDD2.n2 VDD2.t7 1.30916
R2257 VDD2.n2 VDD2.t1 1.30916
R2258 VDD2.n0 VDD2.t9 1.30916
R2259 VDD2.n0 VDD2.t0 1.30916
R2260 VDD2 VDD2.n6 0.636276
R2261 VDD2.n3 VDD2.n1 0.52274
C0 VN VTAIL 13.4388f
C1 VDD2 VP 0.551837f
C2 VP VTAIL 13.453199f
C3 VN VP 8.607151f
C4 VDD1 VDD2 2.01123f
C5 VDD1 VTAIL 11.8878f
C6 VDD1 VN 0.15266f
C7 VDD2 VTAIL 11.936001f
C8 VN VDD2 13.0389f
C9 VDD1 VP 13.433701f
C10 VDD2 B 7.471934f
C11 VDD1 B 7.443674f
C12 VTAIL B 9.245653f
C13 VN B 17.21998f
C14 VP B 15.6724f
C15 VDD2.t8 B 3.28587f
C16 VDD2.t9 B 0.282912f
C17 VDD2.t0 B 0.282912f
C18 VDD2.n0 B 2.56085f
C19 VDD2.n1 B 0.831894f
C20 VDD2.t7 B 0.282912f
C21 VDD2.t1 B 0.282912f
C22 VDD2.n2 B 2.57387f
C23 VDD2.n3 B 2.80723f
C24 VDD2.t2 B 3.27075f
C25 VDD2.n4 B 3.08776f
C26 VDD2.t6 B 0.282912f
C27 VDD2.t4 B 0.282912f
C28 VDD2.n5 B 2.56085f
C29 VDD2.n6 B 0.415945f
C30 VDD2.t5 B 0.282912f
C31 VDD2.t3 B 0.282912f
C32 VDD2.n7 B 2.57383f
C33 VN.n0 B 0.029389f
C34 VN.t8 B 2.17223f
C35 VN.n1 B 0.018135f
C36 VN.n2 B 0.022291f
C37 VN.t2 B 2.17223f
C38 VN.n3 B 0.041935f
C39 VN.n4 B 0.022291f
C40 VN.t9 B 2.17223f
C41 VN.n5 B 0.781933f
C42 VN.n6 B 0.022291f
C43 VN.n7 B 0.041935f
C44 VN.t1 B 2.32944f
C45 VN.n8 B 0.807865f
C46 VN.t0 B 2.17223f
C47 VN.n9 B 0.818238f
C48 VN.n10 B 0.028418f
C49 VN.n11 B 0.192942f
C50 VN.n12 B 0.022291f
C51 VN.n13 B 0.022291f
C52 VN.n14 B 0.026615f
C53 VN.n15 B 0.038077f
C54 VN.n16 B 0.041545f
C55 VN.n17 B 0.022291f
C56 VN.n18 B 0.022291f
C57 VN.n19 B 0.022291f
C58 VN.n20 B 0.041545f
C59 VN.n21 B 0.038077f
C60 VN.n22 B 0.026615f
C61 VN.n23 B 0.022291f
C62 VN.n24 B 0.022291f
C63 VN.n25 B 0.022291f
C64 VN.n26 B 0.028418f
C65 VN.n27 B 0.760899f
C66 VN.n28 B 0.034161f
C67 VN.n29 B 0.044691f
C68 VN.n30 B 0.022291f
C69 VN.n31 B 0.022291f
C70 VN.n32 B 0.022291f
C71 VN.n33 B 0.043802f
C72 VN.n34 B 0.035802f
C73 VN.n35 B 0.837936f
C74 VN.n36 B 0.029944f
C75 VN.n37 B 0.029389f
C76 VN.t7 B 2.17223f
C77 VN.n38 B 0.018135f
C78 VN.n39 B 0.022291f
C79 VN.t3 B 2.17223f
C80 VN.n40 B 0.041935f
C81 VN.n41 B 0.022291f
C82 VN.t5 B 2.17223f
C83 VN.n42 B 0.781933f
C84 VN.n43 B 0.022291f
C85 VN.n44 B 0.041935f
C86 VN.t6 B 2.32944f
C87 VN.n45 B 0.807865f
C88 VN.t4 B 2.17223f
C89 VN.n46 B 0.818238f
C90 VN.n47 B 0.028418f
C91 VN.n48 B 0.192942f
C92 VN.n49 B 0.022291f
C93 VN.n50 B 0.022291f
C94 VN.n51 B 0.026615f
C95 VN.n52 B 0.038077f
C96 VN.n53 B 0.041545f
C97 VN.n54 B 0.022291f
C98 VN.n55 B 0.022291f
C99 VN.n56 B 0.022291f
C100 VN.n57 B 0.041545f
C101 VN.n58 B 0.038077f
C102 VN.n59 B 0.026615f
C103 VN.n60 B 0.022291f
C104 VN.n61 B 0.022291f
C105 VN.n62 B 0.022291f
C106 VN.n63 B 0.028418f
C107 VN.n64 B 0.760899f
C108 VN.n65 B 0.034161f
C109 VN.n66 B 0.044691f
C110 VN.n67 B 0.022291f
C111 VN.n68 B 0.022291f
C112 VN.n69 B 0.022291f
C113 VN.n70 B 0.043802f
C114 VN.n71 B 0.035802f
C115 VN.n72 B 0.837936f
C116 VN.n73 B 1.39936f
C117 VTAIL.t1 B 0.28752f
C118 VTAIL.t8 B 0.28752f
C119 VTAIL.n0 B 2.53478f
C120 VTAIL.n1 B 0.494216f
C121 VTAIL.t12 B 3.23632f
C122 VTAIL.n2 B 0.617058f
C123 VTAIL.t14 B 0.28752f
C124 VTAIL.t11 B 0.28752f
C125 VTAIL.n3 B 2.53478f
C126 VTAIL.n4 B 0.587568f
C127 VTAIL.t17 B 0.28752f
C128 VTAIL.t16 B 0.28752f
C129 VTAIL.n5 B 2.53478f
C130 VTAIL.n6 B 2.10393f
C131 VTAIL.t3 B 0.28752f
C132 VTAIL.t6 B 0.28752f
C133 VTAIL.n7 B 2.53478f
C134 VTAIL.n8 B 2.10392f
C135 VTAIL.t4 B 0.28752f
C136 VTAIL.t5 B 0.28752f
C137 VTAIL.n9 B 2.53478f
C138 VTAIL.n10 B 0.587565f
C139 VTAIL.t19 B 3.23633f
C140 VTAIL.n11 B 0.617055f
C141 VTAIL.t10 B 0.28752f
C142 VTAIL.t13 B 0.28752f
C143 VTAIL.n12 B 2.53478f
C144 VTAIL.n13 B 0.53446f
C145 VTAIL.t15 B 0.28752f
C146 VTAIL.t18 B 0.28752f
C147 VTAIL.n14 B 2.53478f
C148 VTAIL.n15 B 0.587565f
C149 VTAIL.t9 B 3.23633f
C150 VTAIL.n16 B 2.0075f
C151 VTAIL.t0 B 3.23632f
C152 VTAIL.n17 B 2.0075f
C153 VTAIL.t2 B 0.28752f
C154 VTAIL.t7 B 0.28752f
C155 VTAIL.n18 B 2.53478f
C156 VTAIL.n19 B 0.448793f
C157 VDD1.t2 B 3.32394f
C158 VDD1.t4 B 0.286189f
C159 VDD1.t6 B 0.286189f
C160 VDD1.n0 B 2.59051f
C161 VDD1.n1 B 0.84922f
C162 VDD1.t1 B 3.32394f
C163 VDD1.t8 B 0.286189f
C164 VDD1.t5 B 0.286189f
C165 VDD1.n2 B 2.59051f
C166 VDD1.n3 B 0.84153f
C167 VDD1.t0 B 0.286189f
C168 VDD1.t9 B 0.286189f
C169 VDD1.n4 B 2.60368f
C170 VDD1.n5 B 2.95492f
C171 VDD1.t3 B 0.286189f
C172 VDD1.t7 B 0.286189f
C173 VDD1.n6 B 2.5905f
C174 VDD1.n7 B 3.16354f
C175 VP.n0 B 0.029835f
C176 VP.t6 B 2.20524f
C177 VP.n1 B 0.018411f
C178 VP.n2 B 0.02263f
C179 VP.t7 B 2.20524f
C180 VP.n3 B 0.042572f
C181 VP.n4 B 0.02263f
C182 VP.t4 B 2.20524f
C183 VP.n5 B 0.793814f
C184 VP.n6 B 0.02263f
C185 VP.n7 B 0.042572f
C186 VP.n8 B 0.02263f
C187 VP.t2 B 2.20524f
C188 VP.n9 B 0.018411f
C189 VP.n10 B 0.029835f
C190 VP.t1 B 2.20524f
C191 VP.n11 B 0.029835f
C192 VP.t9 B 2.20524f
C193 VP.n12 B 0.018411f
C194 VP.n13 B 0.02263f
C195 VP.t0 B 2.20524f
C196 VP.n14 B 0.042572f
C197 VP.n15 B 0.02263f
C198 VP.t3 B 2.20524f
C199 VP.n16 B 0.793814f
C200 VP.n17 B 0.02263f
C201 VP.n18 B 0.042572f
C202 VP.t8 B 2.36484f
C203 VP.n19 B 0.82014f
C204 VP.t5 B 2.20524f
C205 VP.n20 B 0.830671f
C206 VP.n21 B 0.02885f
C207 VP.n22 B 0.195874f
C208 VP.n23 B 0.02263f
C209 VP.n24 B 0.02263f
C210 VP.n25 B 0.02702f
C211 VP.n26 B 0.038655f
C212 VP.n27 B 0.042176f
C213 VP.n28 B 0.02263f
C214 VP.n29 B 0.02263f
C215 VP.n30 B 0.02263f
C216 VP.n31 B 0.042176f
C217 VP.n32 B 0.038655f
C218 VP.n33 B 0.02702f
C219 VP.n34 B 0.02263f
C220 VP.n35 B 0.02263f
C221 VP.n36 B 0.02263f
C222 VP.n37 B 0.02885f
C223 VP.n38 B 0.772461f
C224 VP.n39 B 0.03468f
C225 VP.n40 B 0.04537f
C226 VP.n41 B 0.02263f
C227 VP.n42 B 0.02263f
C228 VP.n43 B 0.02263f
C229 VP.n44 B 0.044467f
C230 VP.n45 B 0.036346f
C231 VP.n46 B 0.850668f
C232 VP.n47 B 1.40861f
C233 VP.n48 B 1.42362f
C234 VP.n49 B 0.850668f
C235 VP.n50 B 0.036346f
C236 VP.n51 B 0.044467f
C237 VP.n52 B 0.02263f
C238 VP.n53 B 0.02263f
C239 VP.n54 B 0.02263f
C240 VP.n55 B 0.04537f
C241 VP.n56 B 0.03468f
C242 VP.n57 B 0.772461f
C243 VP.n58 B 0.02885f
C244 VP.n59 B 0.02263f
C245 VP.n60 B 0.02263f
C246 VP.n61 B 0.02263f
C247 VP.n62 B 0.02702f
C248 VP.n63 B 0.038655f
C249 VP.n64 B 0.042176f
C250 VP.n65 B 0.02263f
C251 VP.n66 B 0.02263f
C252 VP.n67 B 0.02263f
C253 VP.n68 B 0.042176f
C254 VP.n69 B 0.038655f
C255 VP.n70 B 0.02702f
C256 VP.n71 B 0.02263f
C257 VP.n72 B 0.02263f
C258 VP.n73 B 0.02263f
C259 VP.n74 B 0.02885f
C260 VP.n75 B 0.772461f
C261 VP.n76 B 0.03468f
C262 VP.n77 B 0.04537f
C263 VP.n78 B 0.02263f
C264 VP.n79 B 0.02263f
C265 VP.n80 B 0.02263f
C266 VP.n81 B 0.044467f
C267 VP.n82 B 0.036346f
C268 VP.n83 B 0.850668f
C269 VP.n84 B 0.030399f
.ends

