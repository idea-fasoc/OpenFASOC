* NGSPICE file created from diff_pair_sample_0724.ext - technology: sky130A

.subckt diff_pair_sample_0724 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0 ps=0 w=2.58 l=2.11
X1 VDD1.t7 VP.t0 VTAIL.t15 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X2 VDD2.t7 VN.t0 VTAIL.t7 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=1.0062 ps=5.94 w=2.58 l=2.11
X3 VDD1.t6 VP.t1 VTAIL.t10 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=1.0062 ps=5.94 w=2.58 l=2.11
X4 B.t8 B.t6 B.t7 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0 ps=0 w=2.58 l=2.11
X5 VTAIL.t6 VN.t1 VDD2.t6 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X6 VDD1.t5 VP.t2 VTAIL.t8 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X7 VTAIL.t1 VN.t2 VDD2.t5 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0.4257 ps=2.91 w=2.58 l=2.11
X8 VDD2.t4 VN.t3 VTAIL.t2 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X9 VDD2.t3 VN.t4 VTAIL.t3 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=1.0062 ps=5.94 w=2.58 l=2.11
X10 B.t5 B.t3 B.t4 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0 ps=0 w=2.58 l=2.11
X11 VTAIL.t12 VP.t3 VDD1.t4 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0.4257 ps=2.91 w=2.58 l=2.11
X12 VTAIL.t13 VP.t4 VDD1.t3 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X13 VTAIL.t4 VN.t5 VDD2.t2 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0.4257 ps=2.91 w=2.58 l=2.11
X14 VTAIL.t11 VP.t5 VDD1.t2 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X15 B.t2 B.t0 B.t1 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0 ps=0 w=2.58 l=2.11
X16 VTAIL.t5 VN.t6 VDD2.t1 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X17 VDD1.t1 VP.t6 VTAIL.t9 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=1.0062 ps=5.94 w=2.58 l=2.11
X18 VDD2.t0 VN.t7 VTAIL.t0 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=0.4257 pd=2.91 as=0.4257 ps=2.91 w=2.58 l=2.11
X19 VTAIL.t14 VP.t7 VDD1.t0 w_n3410_n1484# sky130_fd_pr__pfet_01v8 ad=1.0062 pd=5.94 as=0.4257 ps=2.91 w=2.58 l=2.11
R0 B.n391 B.n46 585
R1 B.n393 B.n392 585
R2 B.n394 B.n45 585
R3 B.n396 B.n395 585
R4 B.n397 B.n44 585
R5 B.n399 B.n398 585
R6 B.n400 B.n43 585
R7 B.n402 B.n401 585
R8 B.n403 B.n42 585
R9 B.n405 B.n404 585
R10 B.n406 B.n41 585
R11 B.n408 B.n407 585
R12 B.n409 B.n40 585
R13 B.n411 B.n410 585
R14 B.n413 B.n37 585
R15 B.n415 B.n414 585
R16 B.n416 B.n36 585
R17 B.n418 B.n417 585
R18 B.n419 B.n35 585
R19 B.n421 B.n420 585
R20 B.n422 B.n34 585
R21 B.n424 B.n423 585
R22 B.n425 B.n31 585
R23 B.n428 B.n427 585
R24 B.n429 B.n30 585
R25 B.n431 B.n430 585
R26 B.n432 B.n29 585
R27 B.n434 B.n433 585
R28 B.n435 B.n28 585
R29 B.n437 B.n436 585
R30 B.n438 B.n27 585
R31 B.n440 B.n439 585
R32 B.n441 B.n26 585
R33 B.n443 B.n442 585
R34 B.n444 B.n25 585
R35 B.n446 B.n445 585
R36 B.n447 B.n24 585
R37 B.n390 B.n389 585
R38 B.n388 B.n47 585
R39 B.n387 B.n386 585
R40 B.n385 B.n48 585
R41 B.n384 B.n383 585
R42 B.n382 B.n49 585
R43 B.n381 B.n380 585
R44 B.n379 B.n50 585
R45 B.n378 B.n377 585
R46 B.n376 B.n51 585
R47 B.n375 B.n374 585
R48 B.n373 B.n52 585
R49 B.n372 B.n371 585
R50 B.n370 B.n53 585
R51 B.n369 B.n368 585
R52 B.n367 B.n54 585
R53 B.n366 B.n365 585
R54 B.n364 B.n55 585
R55 B.n363 B.n362 585
R56 B.n361 B.n56 585
R57 B.n360 B.n359 585
R58 B.n358 B.n57 585
R59 B.n357 B.n356 585
R60 B.n355 B.n58 585
R61 B.n354 B.n353 585
R62 B.n352 B.n59 585
R63 B.n351 B.n350 585
R64 B.n349 B.n60 585
R65 B.n348 B.n347 585
R66 B.n346 B.n61 585
R67 B.n345 B.n344 585
R68 B.n343 B.n62 585
R69 B.n342 B.n341 585
R70 B.n340 B.n63 585
R71 B.n339 B.n338 585
R72 B.n337 B.n64 585
R73 B.n336 B.n335 585
R74 B.n334 B.n65 585
R75 B.n333 B.n332 585
R76 B.n331 B.n66 585
R77 B.n330 B.n329 585
R78 B.n328 B.n67 585
R79 B.n327 B.n326 585
R80 B.n325 B.n68 585
R81 B.n324 B.n323 585
R82 B.n322 B.n69 585
R83 B.n321 B.n320 585
R84 B.n319 B.n70 585
R85 B.n318 B.n317 585
R86 B.n316 B.n71 585
R87 B.n315 B.n314 585
R88 B.n313 B.n72 585
R89 B.n312 B.n311 585
R90 B.n310 B.n73 585
R91 B.n309 B.n308 585
R92 B.n307 B.n74 585
R93 B.n306 B.n305 585
R94 B.n304 B.n75 585
R95 B.n303 B.n302 585
R96 B.n301 B.n76 585
R97 B.n300 B.n299 585
R98 B.n298 B.n77 585
R99 B.n297 B.n296 585
R100 B.n295 B.n78 585
R101 B.n294 B.n293 585
R102 B.n292 B.n79 585
R103 B.n291 B.n290 585
R104 B.n289 B.n80 585
R105 B.n288 B.n287 585
R106 B.n286 B.n81 585
R107 B.n285 B.n284 585
R108 B.n283 B.n82 585
R109 B.n282 B.n281 585
R110 B.n280 B.n83 585
R111 B.n279 B.n278 585
R112 B.n277 B.n84 585
R113 B.n276 B.n275 585
R114 B.n274 B.n85 585
R115 B.n273 B.n272 585
R116 B.n271 B.n86 585
R117 B.n270 B.n269 585
R118 B.n268 B.n87 585
R119 B.n267 B.n266 585
R120 B.n265 B.n88 585
R121 B.n264 B.n263 585
R122 B.n262 B.n89 585
R123 B.n261 B.n260 585
R124 B.n259 B.n90 585
R125 B.n258 B.n257 585
R126 B.n201 B.n200 585
R127 B.n202 B.n113 585
R128 B.n204 B.n203 585
R129 B.n205 B.n112 585
R130 B.n207 B.n206 585
R131 B.n208 B.n111 585
R132 B.n210 B.n209 585
R133 B.n211 B.n110 585
R134 B.n213 B.n212 585
R135 B.n214 B.n109 585
R136 B.n216 B.n215 585
R137 B.n217 B.n108 585
R138 B.n219 B.n218 585
R139 B.n220 B.n105 585
R140 B.n223 B.n222 585
R141 B.n224 B.n104 585
R142 B.n226 B.n225 585
R143 B.n227 B.n103 585
R144 B.n229 B.n228 585
R145 B.n230 B.n102 585
R146 B.n232 B.n231 585
R147 B.n233 B.n101 585
R148 B.n235 B.n234 585
R149 B.n237 B.n236 585
R150 B.n238 B.n97 585
R151 B.n240 B.n239 585
R152 B.n241 B.n96 585
R153 B.n243 B.n242 585
R154 B.n244 B.n95 585
R155 B.n246 B.n245 585
R156 B.n247 B.n94 585
R157 B.n249 B.n248 585
R158 B.n250 B.n93 585
R159 B.n252 B.n251 585
R160 B.n253 B.n92 585
R161 B.n255 B.n254 585
R162 B.n256 B.n91 585
R163 B.n199 B.n114 585
R164 B.n198 B.n197 585
R165 B.n196 B.n115 585
R166 B.n195 B.n194 585
R167 B.n193 B.n116 585
R168 B.n192 B.n191 585
R169 B.n190 B.n117 585
R170 B.n189 B.n188 585
R171 B.n187 B.n118 585
R172 B.n186 B.n185 585
R173 B.n184 B.n119 585
R174 B.n183 B.n182 585
R175 B.n181 B.n120 585
R176 B.n180 B.n179 585
R177 B.n178 B.n121 585
R178 B.n177 B.n176 585
R179 B.n175 B.n122 585
R180 B.n174 B.n173 585
R181 B.n172 B.n123 585
R182 B.n171 B.n170 585
R183 B.n169 B.n124 585
R184 B.n168 B.n167 585
R185 B.n166 B.n125 585
R186 B.n165 B.n164 585
R187 B.n163 B.n126 585
R188 B.n162 B.n161 585
R189 B.n160 B.n127 585
R190 B.n159 B.n158 585
R191 B.n157 B.n128 585
R192 B.n156 B.n155 585
R193 B.n154 B.n129 585
R194 B.n153 B.n152 585
R195 B.n151 B.n130 585
R196 B.n150 B.n149 585
R197 B.n148 B.n131 585
R198 B.n147 B.n146 585
R199 B.n145 B.n132 585
R200 B.n144 B.n143 585
R201 B.n142 B.n133 585
R202 B.n141 B.n140 585
R203 B.n139 B.n134 585
R204 B.n138 B.n137 585
R205 B.n136 B.n135 585
R206 B.n2 B.n0 585
R207 B.n513 B.n1 585
R208 B.n512 B.n511 585
R209 B.n510 B.n3 585
R210 B.n509 B.n508 585
R211 B.n507 B.n4 585
R212 B.n506 B.n505 585
R213 B.n504 B.n5 585
R214 B.n503 B.n502 585
R215 B.n501 B.n6 585
R216 B.n500 B.n499 585
R217 B.n498 B.n7 585
R218 B.n497 B.n496 585
R219 B.n495 B.n8 585
R220 B.n494 B.n493 585
R221 B.n492 B.n9 585
R222 B.n491 B.n490 585
R223 B.n489 B.n10 585
R224 B.n488 B.n487 585
R225 B.n486 B.n11 585
R226 B.n485 B.n484 585
R227 B.n483 B.n12 585
R228 B.n482 B.n481 585
R229 B.n480 B.n13 585
R230 B.n479 B.n478 585
R231 B.n477 B.n14 585
R232 B.n476 B.n475 585
R233 B.n474 B.n15 585
R234 B.n473 B.n472 585
R235 B.n471 B.n16 585
R236 B.n470 B.n469 585
R237 B.n468 B.n17 585
R238 B.n467 B.n466 585
R239 B.n465 B.n18 585
R240 B.n464 B.n463 585
R241 B.n462 B.n19 585
R242 B.n461 B.n460 585
R243 B.n459 B.n20 585
R244 B.n458 B.n457 585
R245 B.n456 B.n21 585
R246 B.n455 B.n454 585
R247 B.n453 B.n22 585
R248 B.n452 B.n451 585
R249 B.n450 B.n23 585
R250 B.n449 B.n448 585
R251 B.n515 B.n514 585
R252 B.n200 B.n199 530.939
R253 B.n448 B.n447 530.939
R254 B.n258 B.n91 530.939
R255 B.n391 B.n390 530.939
R256 B.n98 B.t11 273.125
R257 B.n38 B.t7 273.125
R258 B.n106 B.t5 273.123
R259 B.n32 B.t1 273.123
R260 B.n98 B.t9 236.633
R261 B.n106 B.t3 236.633
R262 B.n32 B.t0 236.633
R263 B.n38 B.t6 236.633
R264 B.n99 B.t10 225.803
R265 B.n39 B.t8 225.803
R266 B.n107 B.t4 225.803
R267 B.n33 B.t2 225.803
R268 B.n199 B.n198 163.367
R269 B.n198 B.n115 163.367
R270 B.n194 B.n115 163.367
R271 B.n194 B.n193 163.367
R272 B.n193 B.n192 163.367
R273 B.n192 B.n117 163.367
R274 B.n188 B.n117 163.367
R275 B.n188 B.n187 163.367
R276 B.n187 B.n186 163.367
R277 B.n186 B.n119 163.367
R278 B.n182 B.n119 163.367
R279 B.n182 B.n181 163.367
R280 B.n181 B.n180 163.367
R281 B.n180 B.n121 163.367
R282 B.n176 B.n121 163.367
R283 B.n176 B.n175 163.367
R284 B.n175 B.n174 163.367
R285 B.n174 B.n123 163.367
R286 B.n170 B.n123 163.367
R287 B.n170 B.n169 163.367
R288 B.n169 B.n168 163.367
R289 B.n168 B.n125 163.367
R290 B.n164 B.n125 163.367
R291 B.n164 B.n163 163.367
R292 B.n163 B.n162 163.367
R293 B.n162 B.n127 163.367
R294 B.n158 B.n127 163.367
R295 B.n158 B.n157 163.367
R296 B.n157 B.n156 163.367
R297 B.n156 B.n129 163.367
R298 B.n152 B.n129 163.367
R299 B.n152 B.n151 163.367
R300 B.n151 B.n150 163.367
R301 B.n150 B.n131 163.367
R302 B.n146 B.n131 163.367
R303 B.n146 B.n145 163.367
R304 B.n145 B.n144 163.367
R305 B.n144 B.n133 163.367
R306 B.n140 B.n133 163.367
R307 B.n140 B.n139 163.367
R308 B.n139 B.n138 163.367
R309 B.n138 B.n135 163.367
R310 B.n135 B.n2 163.367
R311 B.n514 B.n2 163.367
R312 B.n514 B.n513 163.367
R313 B.n513 B.n512 163.367
R314 B.n512 B.n3 163.367
R315 B.n508 B.n3 163.367
R316 B.n508 B.n507 163.367
R317 B.n507 B.n506 163.367
R318 B.n506 B.n5 163.367
R319 B.n502 B.n5 163.367
R320 B.n502 B.n501 163.367
R321 B.n501 B.n500 163.367
R322 B.n500 B.n7 163.367
R323 B.n496 B.n7 163.367
R324 B.n496 B.n495 163.367
R325 B.n495 B.n494 163.367
R326 B.n494 B.n9 163.367
R327 B.n490 B.n9 163.367
R328 B.n490 B.n489 163.367
R329 B.n489 B.n488 163.367
R330 B.n488 B.n11 163.367
R331 B.n484 B.n11 163.367
R332 B.n484 B.n483 163.367
R333 B.n483 B.n482 163.367
R334 B.n482 B.n13 163.367
R335 B.n478 B.n13 163.367
R336 B.n478 B.n477 163.367
R337 B.n477 B.n476 163.367
R338 B.n476 B.n15 163.367
R339 B.n472 B.n15 163.367
R340 B.n472 B.n471 163.367
R341 B.n471 B.n470 163.367
R342 B.n470 B.n17 163.367
R343 B.n466 B.n17 163.367
R344 B.n466 B.n465 163.367
R345 B.n465 B.n464 163.367
R346 B.n464 B.n19 163.367
R347 B.n460 B.n19 163.367
R348 B.n460 B.n459 163.367
R349 B.n459 B.n458 163.367
R350 B.n458 B.n21 163.367
R351 B.n454 B.n21 163.367
R352 B.n454 B.n453 163.367
R353 B.n453 B.n452 163.367
R354 B.n452 B.n23 163.367
R355 B.n448 B.n23 163.367
R356 B.n200 B.n113 163.367
R357 B.n204 B.n113 163.367
R358 B.n205 B.n204 163.367
R359 B.n206 B.n205 163.367
R360 B.n206 B.n111 163.367
R361 B.n210 B.n111 163.367
R362 B.n211 B.n210 163.367
R363 B.n212 B.n211 163.367
R364 B.n212 B.n109 163.367
R365 B.n216 B.n109 163.367
R366 B.n217 B.n216 163.367
R367 B.n218 B.n217 163.367
R368 B.n218 B.n105 163.367
R369 B.n223 B.n105 163.367
R370 B.n224 B.n223 163.367
R371 B.n225 B.n224 163.367
R372 B.n225 B.n103 163.367
R373 B.n229 B.n103 163.367
R374 B.n230 B.n229 163.367
R375 B.n231 B.n230 163.367
R376 B.n231 B.n101 163.367
R377 B.n235 B.n101 163.367
R378 B.n236 B.n235 163.367
R379 B.n236 B.n97 163.367
R380 B.n240 B.n97 163.367
R381 B.n241 B.n240 163.367
R382 B.n242 B.n241 163.367
R383 B.n242 B.n95 163.367
R384 B.n246 B.n95 163.367
R385 B.n247 B.n246 163.367
R386 B.n248 B.n247 163.367
R387 B.n248 B.n93 163.367
R388 B.n252 B.n93 163.367
R389 B.n253 B.n252 163.367
R390 B.n254 B.n253 163.367
R391 B.n254 B.n91 163.367
R392 B.n259 B.n258 163.367
R393 B.n260 B.n259 163.367
R394 B.n260 B.n89 163.367
R395 B.n264 B.n89 163.367
R396 B.n265 B.n264 163.367
R397 B.n266 B.n265 163.367
R398 B.n266 B.n87 163.367
R399 B.n270 B.n87 163.367
R400 B.n271 B.n270 163.367
R401 B.n272 B.n271 163.367
R402 B.n272 B.n85 163.367
R403 B.n276 B.n85 163.367
R404 B.n277 B.n276 163.367
R405 B.n278 B.n277 163.367
R406 B.n278 B.n83 163.367
R407 B.n282 B.n83 163.367
R408 B.n283 B.n282 163.367
R409 B.n284 B.n283 163.367
R410 B.n284 B.n81 163.367
R411 B.n288 B.n81 163.367
R412 B.n289 B.n288 163.367
R413 B.n290 B.n289 163.367
R414 B.n290 B.n79 163.367
R415 B.n294 B.n79 163.367
R416 B.n295 B.n294 163.367
R417 B.n296 B.n295 163.367
R418 B.n296 B.n77 163.367
R419 B.n300 B.n77 163.367
R420 B.n301 B.n300 163.367
R421 B.n302 B.n301 163.367
R422 B.n302 B.n75 163.367
R423 B.n306 B.n75 163.367
R424 B.n307 B.n306 163.367
R425 B.n308 B.n307 163.367
R426 B.n308 B.n73 163.367
R427 B.n312 B.n73 163.367
R428 B.n313 B.n312 163.367
R429 B.n314 B.n313 163.367
R430 B.n314 B.n71 163.367
R431 B.n318 B.n71 163.367
R432 B.n319 B.n318 163.367
R433 B.n320 B.n319 163.367
R434 B.n320 B.n69 163.367
R435 B.n324 B.n69 163.367
R436 B.n325 B.n324 163.367
R437 B.n326 B.n325 163.367
R438 B.n326 B.n67 163.367
R439 B.n330 B.n67 163.367
R440 B.n331 B.n330 163.367
R441 B.n332 B.n331 163.367
R442 B.n332 B.n65 163.367
R443 B.n336 B.n65 163.367
R444 B.n337 B.n336 163.367
R445 B.n338 B.n337 163.367
R446 B.n338 B.n63 163.367
R447 B.n342 B.n63 163.367
R448 B.n343 B.n342 163.367
R449 B.n344 B.n343 163.367
R450 B.n344 B.n61 163.367
R451 B.n348 B.n61 163.367
R452 B.n349 B.n348 163.367
R453 B.n350 B.n349 163.367
R454 B.n350 B.n59 163.367
R455 B.n354 B.n59 163.367
R456 B.n355 B.n354 163.367
R457 B.n356 B.n355 163.367
R458 B.n356 B.n57 163.367
R459 B.n360 B.n57 163.367
R460 B.n361 B.n360 163.367
R461 B.n362 B.n361 163.367
R462 B.n362 B.n55 163.367
R463 B.n366 B.n55 163.367
R464 B.n367 B.n366 163.367
R465 B.n368 B.n367 163.367
R466 B.n368 B.n53 163.367
R467 B.n372 B.n53 163.367
R468 B.n373 B.n372 163.367
R469 B.n374 B.n373 163.367
R470 B.n374 B.n51 163.367
R471 B.n378 B.n51 163.367
R472 B.n379 B.n378 163.367
R473 B.n380 B.n379 163.367
R474 B.n380 B.n49 163.367
R475 B.n384 B.n49 163.367
R476 B.n385 B.n384 163.367
R477 B.n386 B.n385 163.367
R478 B.n386 B.n47 163.367
R479 B.n390 B.n47 163.367
R480 B.n447 B.n446 163.367
R481 B.n446 B.n25 163.367
R482 B.n442 B.n25 163.367
R483 B.n442 B.n441 163.367
R484 B.n441 B.n440 163.367
R485 B.n440 B.n27 163.367
R486 B.n436 B.n27 163.367
R487 B.n436 B.n435 163.367
R488 B.n435 B.n434 163.367
R489 B.n434 B.n29 163.367
R490 B.n430 B.n29 163.367
R491 B.n430 B.n429 163.367
R492 B.n429 B.n428 163.367
R493 B.n428 B.n31 163.367
R494 B.n423 B.n31 163.367
R495 B.n423 B.n422 163.367
R496 B.n422 B.n421 163.367
R497 B.n421 B.n35 163.367
R498 B.n417 B.n35 163.367
R499 B.n417 B.n416 163.367
R500 B.n416 B.n415 163.367
R501 B.n415 B.n37 163.367
R502 B.n410 B.n37 163.367
R503 B.n410 B.n409 163.367
R504 B.n409 B.n408 163.367
R505 B.n408 B.n41 163.367
R506 B.n404 B.n41 163.367
R507 B.n404 B.n403 163.367
R508 B.n403 B.n402 163.367
R509 B.n402 B.n43 163.367
R510 B.n398 B.n43 163.367
R511 B.n398 B.n397 163.367
R512 B.n397 B.n396 163.367
R513 B.n396 B.n45 163.367
R514 B.n392 B.n45 163.367
R515 B.n392 B.n391 163.367
R516 B.n100 B.n99 59.5399
R517 B.n221 B.n107 59.5399
R518 B.n426 B.n33 59.5399
R519 B.n412 B.n39 59.5399
R520 B.n99 B.n98 47.3217
R521 B.n107 B.n106 47.3217
R522 B.n33 B.n32 47.3217
R523 B.n39 B.n38 47.3217
R524 B.n449 B.n24 34.4981
R525 B.n389 B.n46 34.4981
R526 B.n257 B.n256 34.4981
R527 B.n201 B.n114 34.4981
R528 B B.n515 18.0485
R529 B.n445 B.n24 10.6151
R530 B.n445 B.n444 10.6151
R531 B.n444 B.n443 10.6151
R532 B.n443 B.n26 10.6151
R533 B.n439 B.n26 10.6151
R534 B.n439 B.n438 10.6151
R535 B.n438 B.n437 10.6151
R536 B.n437 B.n28 10.6151
R537 B.n433 B.n28 10.6151
R538 B.n433 B.n432 10.6151
R539 B.n432 B.n431 10.6151
R540 B.n431 B.n30 10.6151
R541 B.n427 B.n30 10.6151
R542 B.n425 B.n424 10.6151
R543 B.n424 B.n34 10.6151
R544 B.n420 B.n34 10.6151
R545 B.n420 B.n419 10.6151
R546 B.n419 B.n418 10.6151
R547 B.n418 B.n36 10.6151
R548 B.n414 B.n36 10.6151
R549 B.n414 B.n413 10.6151
R550 B.n411 B.n40 10.6151
R551 B.n407 B.n40 10.6151
R552 B.n407 B.n406 10.6151
R553 B.n406 B.n405 10.6151
R554 B.n405 B.n42 10.6151
R555 B.n401 B.n42 10.6151
R556 B.n401 B.n400 10.6151
R557 B.n400 B.n399 10.6151
R558 B.n399 B.n44 10.6151
R559 B.n395 B.n44 10.6151
R560 B.n395 B.n394 10.6151
R561 B.n394 B.n393 10.6151
R562 B.n393 B.n46 10.6151
R563 B.n257 B.n90 10.6151
R564 B.n261 B.n90 10.6151
R565 B.n262 B.n261 10.6151
R566 B.n263 B.n262 10.6151
R567 B.n263 B.n88 10.6151
R568 B.n267 B.n88 10.6151
R569 B.n268 B.n267 10.6151
R570 B.n269 B.n268 10.6151
R571 B.n269 B.n86 10.6151
R572 B.n273 B.n86 10.6151
R573 B.n274 B.n273 10.6151
R574 B.n275 B.n274 10.6151
R575 B.n275 B.n84 10.6151
R576 B.n279 B.n84 10.6151
R577 B.n280 B.n279 10.6151
R578 B.n281 B.n280 10.6151
R579 B.n281 B.n82 10.6151
R580 B.n285 B.n82 10.6151
R581 B.n286 B.n285 10.6151
R582 B.n287 B.n286 10.6151
R583 B.n287 B.n80 10.6151
R584 B.n291 B.n80 10.6151
R585 B.n292 B.n291 10.6151
R586 B.n293 B.n292 10.6151
R587 B.n293 B.n78 10.6151
R588 B.n297 B.n78 10.6151
R589 B.n298 B.n297 10.6151
R590 B.n299 B.n298 10.6151
R591 B.n299 B.n76 10.6151
R592 B.n303 B.n76 10.6151
R593 B.n304 B.n303 10.6151
R594 B.n305 B.n304 10.6151
R595 B.n305 B.n74 10.6151
R596 B.n309 B.n74 10.6151
R597 B.n310 B.n309 10.6151
R598 B.n311 B.n310 10.6151
R599 B.n311 B.n72 10.6151
R600 B.n315 B.n72 10.6151
R601 B.n316 B.n315 10.6151
R602 B.n317 B.n316 10.6151
R603 B.n317 B.n70 10.6151
R604 B.n321 B.n70 10.6151
R605 B.n322 B.n321 10.6151
R606 B.n323 B.n322 10.6151
R607 B.n323 B.n68 10.6151
R608 B.n327 B.n68 10.6151
R609 B.n328 B.n327 10.6151
R610 B.n329 B.n328 10.6151
R611 B.n329 B.n66 10.6151
R612 B.n333 B.n66 10.6151
R613 B.n334 B.n333 10.6151
R614 B.n335 B.n334 10.6151
R615 B.n335 B.n64 10.6151
R616 B.n339 B.n64 10.6151
R617 B.n340 B.n339 10.6151
R618 B.n341 B.n340 10.6151
R619 B.n341 B.n62 10.6151
R620 B.n345 B.n62 10.6151
R621 B.n346 B.n345 10.6151
R622 B.n347 B.n346 10.6151
R623 B.n347 B.n60 10.6151
R624 B.n351 B.n60 10.6151
R625 B.n352 B.n351 10.6151
R626 B.n353 B.n352 10.6151
R627 B.n353 B.n58 10.6151
R628 B.n357 B.n58 10.6151
R629 B.n358 B.n357 10.6151
R630 B.n359 B.n358 10.6151
R631 B.n359 B.n56 10.6151
R632 B.n363 B.n56 10.6151
R633 B.n364 B.n363 10.6151
R634 B.n365 B.n364 10.6151
R635 B.n365 B.n54 10.6151
R636 B.n369 B.n54 10.6151
R637 B.n370 B.n369 10.6151
R638 B.n371 B.n370 10.6151
R639 B.n371 B.n52 10.6151
R640 B.n375 B.n52 10.6151
R641 B.n376 B.n375 10.6151
R642 B.n377 B.n376 10.6151
R643 B.n377 B.n50 10.6151
R644 B.n381 B.n50 10.6151
R645 B.n382 B.n381 10.6151
R646 B.n383 B.n382 10.6151
R647 B.n383 B.n48 10.6151
R648 B.n387 B.n48 10.6151
R649 B.n388 B.n387 10.6151
R650 B.n389 B.n388 10.6151
R651 B.n202 B.n201 10.6151
R652 B.n203 B.n202 10.6151
R653 B.n203 B.n112 10.6151
R654 B.n207 B.n112 10.6151
R655 B.n208 B.n207 10.6151
R656 B.n209 B.n208 10.6151
R657 B.n209 B.n110 10.6151
R658 B.n213 B.n110 10.6151
R659 B.n214 B.n213 10.6151
R660 B.n215 B.n214 10.6151
R661 B.n215 B.n108 10.6151
R662 B.n219 B.n108 10.6151
R663 B.n220 B.n219 10.6151
R664 B.n222 B.n104 10.6151
R665 B.n226 B.n104 10.6151
R666 B.n227 B.n226 10.6151
R667 B.n228 B.n227 10.6151
R668 B.n228 B.n102 10.6151
R669 B.n232 B.n102 10.6151
R670 B.n233 B.n232 10.6151
R671 B.n234 B.n233 10.6151
R672 B.n238 B.n237 10.6151
R673 B.n239 B.n238 10.6151
R674 B.n239 B.n96 10.6151
R675 B.n243 B.n96 10.6151
R676 B.n244 B.n243 10.6151
R677 B.n245 B.n244 10.6151
R678 B.n245 B.n94 10.6151
R679 B.n249 B.n94 10.6151
R680 B.n250 B.n249 10.6151
R681 B.n251 B.n250 10.6151
R682 B.n251 B.n92 10.6151
R683 B.n255 B.n92 10.6151
R684 B.n256 B.n255 10.6151
R685 B.n197 B.n114 10.6151
R686 B.n197 B.n196 10.6151
R687 B.n196 B.n195 10.6151
R688 B.n195 B.n116 10.6151
R689 B.n191 B.n116 10.6151
R690 B.n191 B.n190 10.6151
R691 B.n190 B.n189 10.6151
R692 B.n189 B.n118 10.6151
R693 B.n185 B.n118 10.6151
R694 B.n185 B.n184 10.6151
R695 B.n184 B.n183 10.6151
R696 B.n183 B.n120 10.6151
R697 B.n179 B.n120 10.6151
R698 B.n179 B.n178 10.6151
R699 B.n178 B.n177 10.6151
R700 B.n177 B.n122 10.6151
R701 B.n173 B.n122 10.6151
R702 B.n173 B.n172 10.6151
R703 B.n172 B.n171 10.6151
R704 B.n171 B.n124 10.6151
R705 B.n167 B.n124 10.6151
R706 B.n167 B.n166 10.6151
R707 B.n166 B.n165 10.6151
R708 B.n165 B.n126 10.6151
R709 B.n161 B.n126 10.6151
R710 B.n161 B.n160 10.6151
R711 B.n160 B.n159 10.6151
R712 B.n159 B.n128 10.6151
R713 B.n155 B.n128 10.6151
R714 B.n155 B.n154 10.6151
R715 B.n154 B.n153 10.6151
R716 B.n153 B.n130 10.6151
R717 B.n149 B.n130 10.6151
R718 B.n149 B.n148 10.6151
R719 B.n148 B.n147 10.6151
R720 B.n147 B.n132 10.6151
R721 B.n143 B.n132 10.6151
R722 B.n143 B.n142 10.6151
R723 B.n142 B.n141 10.6151
R724 B.n141 B.n134 10.6151
R725 B.n137 B.n134 10.6151
R726 B.n137 B.n136 10.6151
R727 B.n136 B.n0 10.6151
R728 B.n511 B.n1 10.6151
R729 B.n511 B.n510 10.6151
R730 B.n510 B.n509 10.6151
R731 B.n509 B.n4 10.6151
R732 B.n505 B.n4 10.6151
R733 B.n505 B.n504 10.6151
R734 B.n504 B.n503 10.6151
R735 B.n503 B.n6 10.6151
R736 B.n499 B.n6 10.6151
R737 B.n499 B.n498 10.6151
R738 B.n498 B.n497 10.6151
R739 B.n497 B.n8 10.6151
R740 B.n493 B.n8 10.6151
R741 B.n493 B.n492 10.6151
R742 B.n492 B.n491 10.6151
R743 B.n491 B.n10 10.6151
R744 B.n487 B.n10 10.6151
R745 B.n487 B.n486 10.6151
R746 B.n486 B.n485 10.6151
R747 B.n485 B.n12 10.6151
R748 B.n481 B.n12 10.6151
R749 B.n481 B.n480 10.6151
R750 B.n480 B.n479 10.6151
R751 B.n479 B.n14 10.6151
R752 B.n475 B.n14 10.6151
R753 B.n475 B.n474 10.6151
R754 B.n474 B.n473 10.6151
R755 B.n473 B.n16 10.6151
R756 B.n469 B.n16 10.6151
R757 B.n469 B.n468 10.6151
R758 B.n468 B.n467 10.6151
R759 B.n467 B.n18 10.6151
R760 B.n463 B.n18 10.6151
R761 B.n463 B.n462 10.6151
R762 B.n462 B.n461 10.6151
R763 B.n461 B.n20 10.6151
R764 B.n457 B.n20 10.6151
R765 B.n457 B.n456 10.6151
R766 B.n456 B.n455 10.6151
R767 B.n455 B.n22 10.6151
R768 B.n451 B.n22 10.6151
R769 B.n451 B.n450 10.6151
R770 B.n450 B.n449 10.6151
R771 B.n426 B.n425 6.5566
R772 B.n413 B.n412 6.5566
R773 B.n222 B.n221 6.5566
R774 B.n234 B.n100 6.5566
R775 B.n427 B.n426 4.05904
R776 B.n412 B.n411 4.05904
R777 B.n221 B.n220 4.05904
R778 B.n237 B.n100 4.05904
R779 B.n515 B.n0 2.81026
R780 B.n515 B.n1 2.81026
R781 VP.n15 VP.n12 161.3
R782 VP.n17 VP.n16 161.3
R783 VP.n18 VP.n11 161.3
R784 VP.n20 VP.n19 161.3
R785 VP.n22 VP.n10 161.3
R786 VP.n24 VP.n23 161.3
R787 VP.n25 VP.n9 161.3
R788 VP.n27 VP.n26 161.3
R789 VP.n28 VP.n8 161.3
R790 VP.n54 VP.n0 161.3
R791 VP.n53 VP.n52 161.3
R792 VP.n51 VP.n1 161.3
R793 VP.n50 VP.n49 161.3
R794 VP.n48 VP.n2 161.3
R795 VP.n46 VP.n45 161.3
R796 VP.n44 VP.n3 161.3
R797 VP.n43 VP.n42 161.3
R798 VP.n41 VP.n4 161.3
R799 VP.n39 VP.n38 161.3
R800 VP.n37 VP.n5 161.3
R801 VP.n36 VP.n35 161.3
R802 VP.n34 VP.n6 161.3
R803 VP.n33 VP.n32 161.3
R804 VP.n31 VP.n7 90.7429
R805 VP.n56 VP.n55 90.7429
R806 VP.n30 VP.n29 90.7429
R807 VP.n13 VP.t7 63.7136
R808 VP.n35 VP.n34 56.5617
R809 VP.n42 VP.n3 56.5617
R810 VP.n53 VP.n1 56.5617
R811 VP.n27 VP.n9 56.5617
R812 VP.n16 VP.n11 56.5617
R813 VP.n14 VP.n13 47.6568
R814 VP.n31 VP.n30 41.5224
R815 VP.n7 VP.t3 29.4687
R816 VP.n40 VP.t0 29.4687
R817 VP.n47 VP.t5 29.4687
R818 VP.n55 VP.t1 29.4687
R819 VP.n29 VP.t6 29.4687
R820 VP.n21 VP.t4 29.4687
R821 VP.n14 VP.t2 29.4687
R822 VP.n34 VP.n33 24.5923
R823 VP.n35 VP.n5 24.5923
R824 VP.n39 VP.n5 24.5923
R825 VP.n42 VP.n41 24.5923
R826 VP.n46 VP.n3 24.5923
R827 VP.n49 VP.n48 24.5923
R828 VP.n49 VP.n1 24.5923
R829 VP.n54 VP.n53 24.5923
R830 VP.n28 VP.n27 24.5923
R831 VP.n20 VP.n11 24.5923
R832 VP.n23 VP.n22 24.5923
R833 VP.n23 VP.n9 24.5923
R834 VP.n16 VP.n15 24.5923
R835 VP.n41 VP.n40 23.1168
R836 VP.n47 VP.n46 23.1168
R837 VP.n21 VP.n20 23.1168
R838 VP.n15 VP.n14 23.1168
R839 VP.n33 VP.n7 20.1658
R840 VP.n55 VP.n54 20.1658
R841 VP.n29 VP.n28 20.1658
R842 VP.n13 VP.n12 8.94243
R843 VP.n40 VP.n39 1.47601
R844 VP.n48 VP.n47 1.47601
R845 VP.n22 VP.n21 1.47601
R846 VP.n30 VP.n8 0.278335
R847 VP.n32 VP.n31 0.278335
R848 VP.n56 VP.n0 0.278335
R849 VP.n17 VP.n12 0.189894
R850 VP.n18 VP.n17 0.189894
R851 VP.n19 VP.n18 0.189894
R852 VP.n19 VP.n10 0.189894
R853 VP.n24 VP.n10 0.189894
R854 VP.n25 VP.n24 0.189894
R855 VP.n26 VP.n25 0.189894
R856 VP.n26 VP.n8 0.189894
R857 VP.n32 VP.n6 0.189894
R858 VP.n36 VP.n6 0.189894
R859 VP.n37 VP.n36 0.189894
R860 VP.n38 VP.n37 0.189894
R861 VP.n38 VP.n4 0.189894
R862 VP.n43 VP.n4 0.189894
R863 VP.n44 VP.n43 0.189894
R864 VP.n45 VP.n44 0.189894
R865 VP.n45 VP.n2 0.189894
R866 VP.n50 VP.n2 0.189894
R867 VP.n51 VP.n50 0.189894
R868 VP.n52 VP.n51 0.189894
R869 VP.n52 VP.n0 0.189894
R870 VP VP.n56 0.153485
R871 VTAIL.n98 VTAIL.n92 756.745
R872 VTAIL.n8 VTAIL.n2 756.745
R873 VTAIL.n20 VTAIL.n14 756.745
R874 VTAIL.n34 VTAIL.n28 756.745
R875 VTAIL.n86 VTAIL.n80 756.745
R876 VTAIL.n72 VTAIL.n66 756.745
R877 VTAIL.n60 VTAIL.n54 756.745
R878 VTAIL.n46 VTAIL.n40 756.745
R879 VTAIL.n97 VTAIL.n96 585
R880 VTAIL.n99 VTAIL.n98 585
R881 VTAIL.n7 VTAIL.n6 585
R882 VTAIL.n9 VTAIL.n8 585
R883 VTAIL.n19 VTAIL.n18 585
R884 VTAIL.n21 VTAIL.n20 585
R885 VTAIL.n33 VTAIL.n32 585
R886 VTAIL.n35 VTAIL.n34 585
R887 VTAIL.n87 VTAIL.n86 585
R888 VTAIL.n85 VTAIL.n84 585
R889 VTAIL.n73 VTAIL.n72 585
R890 VTAIL.n71 VTAIL.n70 585
R891 VTAIL.n61 VTAIL.n60 585
R892 VTAIL.n59 VTAIL.n58 585
R893 VTAIL.n47 VTAIL.n46 585
R894 VTAIL.n45 VTAIL.n44 585
R895 VTAIL.n95 VTAIL.t7 355.474
R896 VTAIL.n5 VTAIL.t1 355.474
R897 VTAIL.n17 VTAIL.t10 355.474
R898 VTAIL.n31 VTAIL.t12 355.474
R899 VTAIL.n83 VTAIL.t9 355.474
R900 VTAIL.n69 VTAIL.t14 355.474
R901 VTAIL.n57 VTAIL.t3 355.474
R902 VTAIL.n43 VTAIL.t4 355.474
R903 VTAIL.n98 VTAIL.n97 171.744
R904 VTAIL.n8 VTAIL.n7 171.744
R905 VTAIL.n20 VTAIL.n19 171.744
R906 VTAIL.n34 VTAIL.n33 171.744
R907 VTAIL.n86 VTAIL.n85 171.744
R908 VTAIL.n72 VTAIL.n71 171.744
R909 VTAIL.n60 VTAIL.n59 171.744
R910 VTAIL.n46 VTAIL.n45 171.744
R911 VTAIL.n79 VTAIL.n78 138.532
R912 VTAIL.n53 VTAIL.n52 138.532
R913 VTAIL.n1 VTAIL.n0 138.532
R914 VTAIL.n27 VTAIL.n26 138.532
R915 VTAIL.n97 VTAIL.t7 85.8723
R916 VTAIL.n7 VTAIL.t1 85.8723
R917 VTAIL.n19 VTAIL.t10 85.8723
R918 VTAIL.n33 VTAIL.t12 85.8723
R919 VTAIL.n85 VTAIL.t9 85.8723
R920 VTAIL.n71 VTAIL.t14 85.8723
R921 VTAIL.n59 VTAIL.t3 85.8723
R922 VTAIL.n45 VTAIL.t4 85.8723
R923 VTAIL.n103 VTAIL.n102 35.6763
R924 VTAIL.n13 VTAIL.n12 35.6763
R925 VTAIL.n25 VTAIL.n24 35.6763
R926 VTAIL.n39 VTAIL.n38 35.6763
R927 VTAIL.n91 VTAIL.n90 35.6763
R928 VTAIL.n77 VTAIL.n76 35.6763
R929 VTAIL.n65 VTAIL.n64 35.6763
R930 VTAIL.n51 VTAIL.n50 35.6763
R931 VTAIL.n103 VTAIL.n91 16.6945
R932 VTAIL.n51 VTAIL.n39 16.6945
R933 VTAIL.n96 VTAIL.n95 15.8418
R934 VTAIL.n6 VTAIL.n5 15.8418
R935 VTAIL.n18 VTAIL.n17 15.8418
R936 VTAIL.n32 VTAIL.n31 15.8418
R937 VTAIL.n84 VTAIL.n83 15.8418
R938 VTAIL.n70 VTAIL.n69 15.8418
R939 VTAIL.n58 VTAIL.n57 15.8418
R940 VTAIL.n44 VTAIL.n43 15.8418
R941 VTAIL.n99 VTAIL.n94 12.8005
R942 VTAIL.n9 VTAIL.n4 12.8005
R943 VTAIL.n21 VTAIL.n16 12.8005
R944 VTAIL.n35 VTAIL.n30 12.8005
R945 VTAIL.n87 VTAIL.n82 12.8005
R946 VTAIL.n73 VTAIL.n68 12.8005
R947 VTAIL.n61 VTAIL.n56 12.8005
R948 VTAIL.n47 VTAIL.n42 12.8005
R949 VTAIL.n0 VTAIL.t0 12.5993
R950 VTAIL.n0 VTAIL.t6 12.5993
R951 VTAIL.n26 VTAIL.t15 12.5993
R952 VTAIL.n26 VTAIL.t11 12.5993
R953 VTAIL.n78 VTAIL.t8 12.5993
R954 VTAIL.n78 VTAIL.t13 12.5993
R955 VTAIL.n52 VTAIL.t2 12.5993
R956 VTAIL.n52 VTAIL.t5 12.5993
R957 VTAIL.n100 VTAIL.n92 12.0247
R958 VTAIL.n10 VTAIL.n2 12.0247
R959 VTAIL.n22 VTAIL.n14 12.0247
R960 VTAIL.n36 VTAIL.n28 12.0247
R961 VTAIL.n88 VTAIL.n80 12.0247
R962 VTAIL.n74 VTAIL.n66 12.0247
R963 VTAIL.n62 VTAIL.n54 12.0247
R964 VTAIL.n48 VTAIL.n40 12.0247
R965 VTAIL.n102 VTAIL.n101 9.45567
R966 VTAIL.n12 VTAIL.n11 9.45567
R967 VTAIL.n24 VTAIL.n23 9.45567
R968 VTAIL.n38 VTAIL.n37 9.45567
R969 VTAIL.n90 VTAIL.n89 9.45567
R970 VTAIL.n76 VTAIL.n75 9.45567
R971 VTAIL.n64 VTAIL.n63 9.45567
R972 VTAIL.n50 VTAIL.n49 9.45567
R973 VTAIL.n101 VTAIL.n100 9.3005
R974 VTAIL.n94 VTAIL.n93 9.3005
R975 VTAIL.n11 VTAIL.n10 9.3005
R976 VTAIL.n4 VTAIL.n3 9.3005
R977 VTAIL.n23 VTAIL.n22 9.3005
R978 VTAIL.n16 VTAIL.n15 9.3005
R979 VTAIL.n37 VTAIL.n36 9.3005
R980 VTAIL.n30 VTAIL.n29 9.3005
R981 VTAIL.n89 VTAIL.n88 9.3005
R982 VTAIL.n82 VTAIL.n81 9.3005
R983 VTAIL.n75 VTAIL.n74 9.3005
R984 VTAIL.n68 VTAIL.n67 9.3005
R985 VTAIL.n63 VTAIL.n62 9.3005
R986 VTAIL.n56 VTAIL.n55 9.3005
R987 VTAIL.n49 VTAIL.n48 9.3005
R988 VTAIL.n42 VTAIL.n41 9.3005
R989 VTAIL.n83 VTAIL.n81 4.29255
R990 VTAIL.n69 VTAIL.n67 4.29255
R991 VTAIL.n57 VTAIL.n55 4.29255
R992 VTAIL.n43 VTAIL.n41 4.29255
R993 VTAIL.n95 VTAIL.n93 4.29255
R994 VTAIL.n5 VTAIL.n3 4.29255
R995 VTAIL.n17 VTAIL.n15 4.29255
R996 VTAIL.n31 VTAIL.n29 4.29255
R997 VTAIL.n53 VTAIL.n51 2.10395
R998 VTAIL.n65 VTAIL.n53 2.10395
R999 VTAIL.n79 VTAIL.n77 2.10395
R1000 VTAIL.n91 VTAIL.n79 2.10395
R1001 VTAIL.n39 VTAIL.n27 2.10395
R1002 VTAIL.n27 VTAIL.n25 2.10395
R1003 VTAIL.n13 VTAIL.n1 2.10395
R1004 VTAIL VTAIL.n103 2.04576
R1005 VTAIL.n102 VTAIL.n92 1.93989
R1006 VTAIL.n12 VTAIL.n2 1.93989
R1007 VTAIL.n24 VTAIL.n14 1.93989
R1008 VTAIL.n38 VTAIL.n28 1.93989
R1009 VTAIL.n90 VTAIL.n80 1.93989
R1010 VTAIL.n76 VTAIL.n66 1.93989
R1011 VTAIL.n64 VTAIL.n54 1.93989
R1012 VTAIL.n50 VTAIL.n40 1.93989
R1013 VTAIL.n100 VTAIL.n99 1.16414
R1014 VTAIL.n10 VTAIL.n9 1.16414
R1015 VTAIL.n22 VTAIL.n21 1.16414
R1016 VTAIL.n36 VTAIL.n35 1.16414
R1017 VTAIL.n88 VTAIL.n87 1.16414
R1018 VTAIL.n74 VTAIL.n73 1.16414
R1019 VTAIL.n62 VTAIL.n61 1.16414
R1020 VTAIL.n48 VTAIL.n47 1.16414
R1021 VTAIL.n77 VTAIL.n65 0.470328
R1022 VTAIL.n25 VTAIL.n13 0.470328
R1023 VTAIL.n96 VTAIL.n94 0.388379
R1024 VTAIL.n6 VTAIL.n4 0.388379
R1025 VTAIL.n18 VTAIL.n16 0.388379
R1026 VTAIL.n32 VTAIL.n30 0.388379
R1027 VTAIL.n84 VTAIL.n82 0.388379
R1028 VTAIL.n70 VTAIL.n68 0.388379
R1029 VTAIL.n58 VTAIL.n56 0.388379
R1030 VTAIL.n44 VTAIL.n42 0.388379
R1031 VTAIL.n101 VTAIL.n93 0.155672
R1032 VTAIL.n11 VTAIL.n3 0.155672
R1033 VTAIL.n23 VTAIL.n15 0.155672
R1034 VTAIL.n37 VTAIL.n29 0.155672
R1035 VTAIL.n89 VTAIL.n81 0.155672
R1036 VTAIL.n75 VTAIL.n67 0.155672
R1037 VTAIL.n63 VTAIL.n55 0.155672
R1038 VTAIL.n49 VTAIL.n41 0.155672
R1039 VTAIL VTAIL.n1 0.0586897
R1040 VDD1 VDD1.n0 156.321
R1041 VDD1.n3 VDD1.n2 156.208
R1042 VDD1.n3 VDD1.n1 156.208
R1043 VDD1.n5 VDD1.n4 155.212
R1044 VDD1.n5 VDD1.n3 35.988
R1045 VDD1.n4 VDD1.t3 12.5993
R1046 VDD1.n4 VDD1.t1 12.5993
R1047 VDD1.n0 VDD1.t0 12.5993
R1048 VDD1.n0 VDD1.t5 12.5993
R1049 VDD1.n2 VDD1.t2 12.5993
R1050 VDD1.n2 VDD1.t6 12.5993
R1051 VDD1.n1 VDD1.t4 12.5993
R1052 VDD1.n1 VDD1.t7 12.5993
R1053 VDD1 VDD1.n5 0.994035
R1054 VN.n43 VN.n23 161.3
R1055 VN.n42 VN.n41 161.3
R1056 VN.n40 VN.n24 161.3
R1057 VN.n39 VN.n38 161.3
R1058 VN.n37 VN.n25 161.3
R1059 VN.n35 VN.n34 161.3
R1060 VN.n33 VN.n26 161.3
R1061 VN.n32 VN.n31 161.3
R1062 VN.n30 VN.n27 161.3
R1063 VN.n20 VN.n0 161.3
R1064 VN.n19 VN.n18 161.3
R1065 VN.n17 VN.n1 161.3
R1066 VN.n16 VN.n15 161.3
R1067 VN.n14 VN.n2 161.3
R1068 VN.n12 VN.n11 161.3
R1069 VN.n10 VN.n3 161.3
R1070 VN.n9 VN.n8 161.3
R1071 VN.n7 VN.n4 161.3
R1072 VN.n22 VN.n21 90.7429
R1073 VN.n45 VN.n44 90.7429
R1074 VN.n5 VN.t2 63.7136
R1075 VN.n28 VN.t4 63.7136
R1076 VN.n8 VN.n3 56.5617
R1077 VN.n19 VN.n1 56.5617
R1078 VN.n31 VN.n26 56.5617
R1079 VN.n42 VN.n24 56.5617
R1080 VN.n6 VN.n5 47.6568
R1081 VN.n29 VN.n28 47.6568
R1082 VN VN.n45 41.8012
R1083 VN.n6 VN.t7 29.4687
R1084 VN.n13 VN.t1 29.4687
R1085 VN.n21 VN.t0 29.4687
R1086 VN.n29 VN.t6 29.4687
R1087 VN.n36 VN.t3 29.4687
R1088 VN.n44 VN.t5 29.4687
R1089 VN.n8 VN.n7 24.5923
R1090 VN.n12 VN.n3 24.5923
R1091 VN.n15 VN.n14 24.5923
R1092 VN.n15 VN.n1 24.5923
R1093 VN.n20 VN.n19 24.5923
R1094 VN.n31 VN.n30 24.5923
R1095 VN.n38 VN.n24 24.5923
R1096 VN.n38 VN.n37 24.5923
R1097 VN.n35 VN.n26 24.5923
R1098 VN.n43 VN.n42 24.5923
R1099 VN.n7 VN.n6 23.1168
R1100 VN.n13 VN.n12 23.1168
R1101 VN.n30 VN.n29 23.1168
R1102 VN.n36 VN.n35 23.1168
R1103 VN.n21 VN.n20 20.1658
R1104 VN.n44 VN.n43 20.1658
R1105 VN.n28 VN.n27 8.94243
R1106 VN.n5 VN.n4 8.94243
R1107 VN.n14 VN.n13 1.47601
R1108 VN.n37 VN.n36 1.47601
R1109 VN.n45 VN.n23 0.278335
R1110 VN.n22 VN.n0 0.278335
R1111 VN.n41 VN.n23 0.189894
R1112 VN.n41 VN.n40 0.189894
R1113 VN.n40 VN.n39 0.189894
R1114 VN.n39 VN.n25 0.189894
R1115 VN.n34 VN.n25 0.189894
R1116 VN.n34 VN.n33 0.189894
R1117 VN.n33 VN.n32 0.189894
R1118 VN.n32 VN.n27 0.189894
R1119 VN.n9 VN.n4 0.189894
R1120 VN.n10 VN.n9 0.189894
R1121 VN.n11 VN.n10 0.189894
R1122 VN.n11 VN.n2 0.189894
R1123 VN.n16 VN.n2 0.189894
R1124 VN.n17 VN.n16 0.189894
R1125 VN.n18 VN.n17 0.189894
R1126 VN.n18 VN.n0 0.189894
R1127 VN VN.n22 0.153485
R1128 VDD2.n2 VDD2.n1 156.208
R1129 VDD2.n2 VDD2.n0 156.208
R1130 VDD2 VDD2.n5 156.204
R1131 VDD2.n4 VDD2.n3 155.212
R1132 VDD2.n4 VDD2.n2 35.4049
R1133 VDD2.n5 VDD2.t1 12.5993
R1134 VDD2.n5 VDD2.t3 12.5993
R1135 VDD2.n3 VDD2.t2 12.5993
R1136 VDD2.n3 VDD2.t4 12.5993
R1137 VDD2.n1 VDD2.t6 12.5993
R1138 VDD2.n1 VDD2.t7 12.5993
R1139 VDD2.n0 VDD2.t5 12.5993
R1140 VDD2.n0 VDD2.t0 12.5993
R1141 VDD2 VDD2.n4 1.11041
C0 VP VTAIL 2.99827f
C1 VDD1 B 1.24633f
C2 B VN 1.0106f
C3 VDD1 VTAIL 4.51287f
C4 B VDD2 1.32716f
C5 w_n3410_n1484# B 6.74973f
C6 VTAIL VN 2.98417f
C7 VDD2 VTAIL 4.564f
C8 w_n3410_n1484# VTAIL 1.98879f
C9 VDD1 VP 2.44485f
C10 VP VN 5.32038f
C11 VP VDD2 0.474105f
C12 B VTAIL 1.69008f
C13 VP w_n3410_n1484# 7.05466f
C14 VDD1 VN 0.156549f
C15 VDD1 VDD2 1.52302f
C16 VDD1 w_n3410_n1484# 1.54085f
C17 VDD2 VN 2.1295f
C18 w_n3410_n1484# VN 6.61649f
C19 w_n3410_n1484# VDD2 1.63439f
C20 VP B 1.74711f
C21 VDD2 VSUBS 1.266149f
C22 VDD1 VSUBS 1.830763f
C23 VTAIL VSUBS 0.505627f
C24 VN VSUBS 5.98125f
C25 VP VSUBS 2.535439f
C26 B VSUBS 3.441663f
C27 w_n3410_n1484# VSUBS 64.2853f
C28 VDD2.t5 VSUBS 0.049539f
C29 VDD2.t0 VSUBS 0.049539f
C30 VDD2.n0 VSUBS 0.247172f
C31 VDD2.t6 VSUBS 0.049539f
C32 VDD2.t7 VSUBS 0.049539f
C33 VDD2.n1 VSUBS 0.247172f
C34 VDD2.n2 VSUBS 2.54134f
C35 VDD2.t2 VSUBS 0.049539f
C36 VDD2.t4 VSUBS 0.049539f
C37 VDD2.n3 VSUBS 0.243713f
C38 VDD2.n4 VSUBS 2.07415f
C39 VDD2.t1 VSUBS 0.049539f
C40 VDD2.t3 VSUBS 0.049539f
C41 VDD2.n5 VSUBS 0.247158f
C42 VN.n0 VSUBS 0.068081f
C43 VN.t0 VSUBS 0.686064f
C44 VN.n1 VSUBS 0.066497f
C45 VN.n2 VSUBS 0.051642f
C46 VN.t1 VSUBS 0.686064f
C47 VN.n3 VSUBS 0.07507f
C48 VN.n4 VSUBS 0.43507f
C49 VN.t7 VSUBS 0.686064f
C50 VN.t2 VSUBS 1.00228f
C51 VN.n5 VSUBS 0.412482f
C52 VN.n6 VSUBS 0.46075f
C53 VN.n7 VSUBS 0.092929f
C54 VN.n8 VSUBS 0.07507f
C55 VN.n9 VSUBS 0.051642f
C56 VN.n10 VSUBS 0.051642f
C57 VN.n11 VSUBS 0.051642f
C58 VN.n12 VSUBS 0.092929f
C59 VN.n13 VSUBS 0.309895f
C60 VN.n14 VSUBS 0.051325f
C61 VN.n15 VSUBS 0.095765f
C62 VN.n16 VSUBS 0.051642f
C63 VN.n17 VSUBS 0.051642f
C64 VN.n18 VSUBS 0.051642f
C65 VN.n19 VSUBS 0.083642f
C66 VN.n20 VSUBS 0.087255f
C67 VN.n21 VSUBS 0.476714f
C68 VN.n22 VSUBS 0.063168f
C69 VN.n23 VSUBS 0.068081f
C70 VN.t5 VSUBS 0.686064f
C71 VN.n24 VSUBS 0.066497f
C72 VN.n25 VSUBS 0.051642f
C73 VN.t3 VSUBS 0.686064f
C74 VN.n26 VSUBS 0.07507f
C75 VN.n27 VSUBS 0.43507f
C76 VN.t6 VSUBS 0.686064f
C77 VN.t4 VSUBS 1.00228f
C78 VN.n28 VSUBS 0.412482f
C79 VN.n29 VSUBS 0.46075f
C80 VN.n30 VSUBS 0.092929f
C81 VN.n31 VSUBS 0.07507f
C82 VN.n32 VSUBS 0.051642f
C83 VN.n33 VSUBS 0.051642f
C84 VN.n34 VSUBS 0.051642f
C85 VN.n35 VSUBS 0.092929f
C86 VN.n36 VSUBS 0.309895f
C87 VN.n37 VSUBS 0.051325f
C88 VN.n38 VSUBS 0.095765f
C89 VN.n39 VSUBS 0.051642f
C90 VN.n40 VSUBS 0.051642f
C91 VN.n41 VSUBS 0.051642f
C92 VN.n42 VSUBS 0.083642f
C93 VN.n43 VSUBS 0.087255f
C94 VN.n44 VSUBS 0.476714f
C95 VN.n45 VSUBS 2.16449f
C96 VDD1.t0 VSUBS 0.050343f
C97 VDD1.t5 VSUBS 0.050343f
C98 VDD1.n0 VSUBS 0.251645f
C99 VDD1.t4 VSUBS 0.050343f
C100 VDD1.t7 VSUBS 0.050343f
C101 VDD1.n1 VSUBS 0.251186f
C102 VDD1.t2 VSUBS 0.050343f
C103 VDD1.t6 VSUBS 0.050343f
C104 VDD1.n2 VSUBS 0.251186f
C105 VDD1.n3 VSUBS 2.63454f
C106 VDD1.t3 VSUBS 0.050343f
C107 VDD1.t1 VSUBS 0.050343f
C108 VDD1.n4 VSUBS 0.247669f
C109 VDD1.n5 VSUBS 2.13784f
C110 VTAIL.t0 VSUBS 0.057822f
C111 VTAIL.t6 VSUBS 0.057822f
C112 VTAIL.n0 VSUBS 0.244433f
C113 VTAIL.n1 VSUBS 0.536911f
C114 VTAIL.n2 VSUBS 0.030803f
C115 VTAIL.n3 VSUBS 0.207222f
C116 VTAIL.n4 VSUBS 0.01524f
C117 VTAIL.t1 VSUBS 0.081954f
C118 VTAIL.n5 VSUBS 0.096579f
C119 VTAIL.n6 VSUBS 0.021239f
C120 VTAIL.n7 VSUBS 0.027016f
C121 VTAIL.n8 VSUBS 0.085981f
C122 VTAIL.n9 VSUBS 0.016136f
C123 VTAIL.n10 VSUBS 0.01524f
C124 VTAIL.n11 VSUBS 0.072529f
C125 VTAIL.n12 VSUBS 0.04339f
C126 VTAIL.n13 VSUBS 0.263327f
C127 VTAIL.n14 VSUBS 0.030803f
C128 VTAIL.n15 VSUBS 0.207222f
C129 VTAIL.n16 VSUBS 0.01524f
C130 VTAIL.t10 VSUBS 0.081954f
C131 VTAIL.n17 VSUBS 0.096579f
C132 VTAIL.n18 VSUBS 0.021239f
C133 VTAIL.n19 VSUBS 0.027016f
C134 VTAIL.n20 VSUBS 0.085981f
C135 VTAIL.n21 VSUBS 0.016136f
C136 VTAIL.n22 VSUBS 0.01524f
C137 VTAIL.n23 VSUBS 0.072529f
C138 VTAIL.n24 VSUBS 0.04339f
C139 VTAIL.n25 VSUBS 0.263327f
C140 VTAIL.t15 VSUBS 0.057822f
C141 VTAIL.t11 VSUBS 0.057822f
C142 VTAIL.n26 VSUBS 0.244433f
C143 VTAIL.n27 VSUBS 0.723817f
C144 VTAIL.n28 VSUBS 0.030803f
C145 VTAIL.n29 VSUBS 0.207222f
C146 VTAIL.n30 VSUBS 0.01524f
C147 VTAIL.t12 VSUBS 0.081954f
C148 VTAIL.n31 VSUBS 0.096579f
C149 VTAIL.n32 VSUBS 0.021239f
C150 VTAIL.n33 VSUBS 0.027016f
C151 VTAIL.n34 VSUBS 0.085981f
C152 VTAIL.n35 VSUBS 0.016136f
C153 VTAIL.n36 VSUBS 0.01524f
C154 VTAIL.n37 VSUBS 0.072529f
C155 VTAIL.n38 VSUBS 0.04339f
C156 VTAIL.n39 VSUBS 1.00112f
C157 VTAIL.n40 VSUBS 0.030803f
C158 VTAIL.n41 VSUBS 0.207222f
C159 VTAIL.n42 VSUBS 0.01524f
C160 VTAIL.t4 VSUBS 0.081954f
C161 VTAIL.n43 VSUBS 0.096579f
C162 VTAIL.n44 VSUBS 0.021239f
C163 VTAIL.n45 VSUBS 0.027016f
C164 VTAIL.n46 VSUBS 0.085981f
C165 VTAIL.n47 VSUBS 0.016136f
C166 VTAIL.n48 VSUBS 0.01524f
C167 VTAIL.n49 VSUBS 0.072529f
C168 VTAIL.n50 VSUBS 0.04339f
C169 VTAIL.n51 VSUBS 1.00112f
C170 VTAIL.t2 VSUBS 0.057822f
C171 VTAIL.t5 VSUBS 0.057822f
C172 VTAIL.n52 VSUBS 0.244435f
C173 VTAIL.n53 VSUBS 0.723815f
C174 VTAIL.n54 VSUBS 0.030803f
C175 VTAIL.n55 VSUBS 0.207222f
C176 VTAIL.n56 VSUBS 0.01524f
C177 VTAIL.t3 VSUBS 0.081954f
C178 VTAIL.n57 VSUBS 0.096579f
C179 VTAIL.n58 VSUBS 0.021239f
C180 VTAIL.n59 VSUBS 0.027016f
C181 VTAIL.n60 VSUBS 0.085981f
C182 VTAIL.n61 VSUBS 0.016136f
C183 VTAIL.n62 VSUBS 0.01524f
C184 VTAIL.n63 VSUBS 0.072529f
C185 VTAIL.n64 VSUBS 0.04339f
C186 VTAIL.n65 VSUBS 0.263327f
C187 VTAIL.n66 VSUBS 0.030803f
C188 VTAIL.n67 VSUBS 0.207222f
C189 VTAIL.n68 VSUBS 0.01524f
C190 VTAIL.t14 VSUBS 0.081954f
C191 VTAIL.n69 VSUBS 0.096579f
C192 VTAIL.n70 VSUBS 0.021239f
C193 VTAIL.n71 VSUBS 0.027016f
C194 VTAIL.n72 VSUBS 0.085981f
C195 VTAIL.n73 VSUBS 0.016136f
C196 VTAIL.n74 VSUBS 0.01524f
C197 VTAIL.n75 VSUBS 0.072529f
C198 VTAIL.n76 VSUBS 0.04339f
C199 VTAIL.n77 VSUBS 0.263327f
C200 VTAIL.t8 VSUBS 0.057822f
C201 VTAIL.t13 VSUBS 0.057822f
C202 VTAIL.n78 VSUBS 0.244435f
C203 VTAIL.n79 VSUBS 0.723815f
C204 VTAIL.n80 VSUBS 0.030803f
C205 VTAIL.n81 VSUBS 0.207222f
C206 VTAIL.n82 VSUBS 0.01524f
C207 VTAIL.t9 VSUBS 0.081954f
C208 VTAIL.n83 VSUBS 0.096579f
C209 VTAIL.n84 VSUBS 0.021239f
C210 VTAIL.n85 VSUBS 0.027016f
C211 VTAIL.n86 VSUBS 0.085981f
C212 VTAIL.n87 VSUBS 0.016136f
C213 VTAIL.n88 VSUBS 0.01524f
C214 VTAIL.n89 VSUBS 0.072529f
C215 VTAIL.n90 VSUBS 0.04339f
C216 VTAIL.n91 VSUBS 1.00112f
C217 VTAIL.n92 VSUBS 0.030803f
C218 VTAIL.n93 VSUBS 0.207222f
C219 VTAIL.n94 VSUBS 0.01524f
C220 VTAIL.t7 VSUBS 0.081954f
C221 VTAIL.n95 VSUBS 0.096579f
C222 VTAIL.n96 VSUBS 0.021239f
C223 VTAIL.n97 VSUBS 0.027016f
C224 VTAIL.n98 VSUBS 0.085981f
C225 VTAIL.n99 VSUBS 0.016136f
C226 VTAIL.n100 VSUBS 0.01524f
C227 VTAIL.n101 VSUBS 0.072529f
C228 VTAIL.n102 VSUBS 0.04339f
C229 VTAIL.n103 VSUBS 0.9958f
C230 VP.n0 VSUBS 0.07159f
C231 VP.t1 VSUBS 0.72143f
C232 VP.n1 VSUBS 0.069925f
C233 VP.n2 VSUBS 0.054304f
C234 VP.t5 VSUBS 0.72143f
C235 VP.n3 VSUBS 0.078939f
C236 VP.n4 VSUBS 0.054304f
C237 VP.t0 VSUBS 0.72143f
C238 VP.n5 VSUBS 0.100702f
C239 VP.n6 VSUBS 0.054304f
C240 VP.t3 VSUBS 0.72143f
C241 VP.n7 VSUBS 0.501288f
C242 VP.n8 VSUBS 0.07159f
C243 VP.t6 VSUBS 0.72143f
C244 VP.n9 VSUBS 0.069925f
C245 VP.n10 VSUBS 0.054304f
C246 VP.t4 VSUBS 0.72143f
C247 VP.n11 VSUBS 0.078939f
C248 VP.n12 VSUBS 0.457498f
C249 VP.t2 VSUBS 0.72143f
C250 VP.t7 VSUBS 1.05395f
C251 VP.n13 VSUBS 0.433745f
C252 VP.n14 VSUBS 0.484501f
C253 VP.n15 VSUBS 0.097719f
C254 VP.n16 VSUBS 0.078939f
C255 VP.n17 VSUBS 0.054304f
C256 VP.n18 VSUBS 0.054304f
C257 VP.n19 VSUBS 0.054304f
C258 VP.n20 VSUBS 0.097719f
C259 VP.n21 VSUBS 0.32587f
C260 VP.n22 VSUBS 0.053971f
C261 VP.n23 VSUBS 0.100702f
C262 VP.n24 VSUBS 0.054304f
C263 VP.n25 VSUBS 0.054304f
C264 VP.n26 VSUBS 0.054304f
C265 VP.n27 VSUBS 0.087954f
C266 VP.n28 VSUBS 0.091753f
C267 VP.n29 VSUBS 0.501288f
C268 VP.n30 VSUBS 2.24594f
C269 VP.n31 VSUBS 2.29309f
C270 VP.n32 VSUBS 0.07159f
C271 VP.n33 VSUBS 0.091753f
C272 VP.n34 VSUBS 0.087954f
C273 VP.n35 VSUBS 0.069925f
C274 VP.n36 VSUBS 0.054304f
C275 VP.n37 VSUBS 0.054304f
C276 VP.n38 VSUBS 0.054304f
C277 VP.n39 VSUBS 0.053971f
C278 VP.n40 VSUBS 0.32587f
C279 VP.n41 VSUBS 0.097719f
C280 VP.n42 VSUBS 0.078939f
C281 VP.n43 VSUBS 0.054304f
C282 VP.n44 VSUBS 0.054304f
C283 VP.n45 VSUBS 0.054304f
C284 VP.n46 VSUBS 0.097719f
C285 VP.n47 VSUBS 0.32587f
C286 VP.n48 VSUBS 0.053971f
C287 VP.n49 VSUBS 0.100702f
C288 VP.n50 VSUBS 0.054304f
C289 VP.n51 VSUBS 0.054304f
C290 VP.n52 VSUBS 0.054304f
C291 VP.n53 VSUBS 0.087954f
C292 VP.n54 VSUBS 0.091753f
C293 VP.n55 VSUBS 0.501288f
C294 VP.n56 VSUBS 0.066424f
C295 B.n0 VSUBS 0.005053f
C296 B.n1 VSUBS 0.005053f
C297 B.n2 VSUBS 0.007991f
C298 B.n3 VSUBS 0.007991f
C299 B.n4 VSUBS 0.007991f
C300 B.n5 VSUBS 0.007991f
C301 B.n6 VSUBS 0.007991f
C302 B.n7 VSUBS 0.007991f
C303 B.n8 VSUBS 0.007991f
C304 B.n9 VSUBS 0.007991f
C305 B.n10 VSUBS 0.007991f
C306 B.n11 VSUBS 0.007991f
C307 B.n12 VSUBS 0.007991f
C308 B.n13 VSUBS 0.007991f
C309 B.n14 VSUBS 0.007991f
C310 B.n15 VSUBS 0.007991f
C311 B.n16 VSUBS 0.007991f
C312 B.n17 VSUBS 0.007991f
C313 B.n18 VSUBS 0.007991f
C314 B.n19 VSUBS 0.007991f
C315 B.n20 VSUBS 0.007991f
C316 B.n21 VSUBS 0.007991f
C317 B.n22 VSUBS 0.007991f
C318 B.n23 VSUBS 0.007991f
C319 B.n24 VSUBS 0.019661f
C320 B.n25 VSUBS 0.007991f
C321 B.n26 VSUBS 0.007991f
C322 B.n27 VSUBS 0.007991f
C323 B.n28 VSUBS 0.007991f
C324 B.n29 VSUBS 0.007991f
C325 B.n30 VSUBS 0.007991f
C326 B.n31 VSUBS 0.007991f
C327 B.t2 VSUBS 0.045769f
C328 B.t1 VSUBS 0.059647f
C329 B.t0 VSUBS 0.302104f
C330 B.n32 VSUBS 0.105481f
C331 B.n33 VSUBS 0.091496f
C332 B.n34 VSUBS 0.007991f
C333 B.n35 VSUBS 0.007991f
C334 B.n36 VSUBS 0.007991f
C335 B.n37 VSUBS 0.007991f
C336 B.t8 VSUBS 0.04577f
C337 B.t7 VSUBS 0.059647f
C338 B.t6 VSUBS 0.302104f
C339 B.n38 VSUBS 0.105481f
C340 B.n39 VSUBS 0.091496f
C341 B.n40 VSUBS 0.007991f
C342 B.n41 VSUBS 0.007991f
C343 B.n42 VSUBS 0.007991f
C344 B.n43 VSUBS 0.007991f
C345 B.n44 VSUBS 0.007991f
C346 B.n45 VSUBS 0.007991f
C347 B.n46 VSUBS 0.018768f
C348 B.n47 VSUBS 0.007991f
C349 B.n48 VSUBS 0.007991f
C350 B.n49 VSUBS 0.007991f
C351 B.n50 VSUBS 0.007991f
C352 B.n51 VSUBS 0.007991f
C353 B.n52 VSUBS 0.007991f
C354 B.n53 VSUBS 0.007991f
C355 B.n54 VSUBS 0.007991f
C356 B.n55 VSUBS 0.007991f
C357 B.n56 VSUBS 0.007991f
C358 B.n57 VSUBS 0.007991f
C359 B.n58 VSUBS 0.007991f
C360 B.n59 VSUBS 0.007991f
C361 B.n60 VSUBS 0.007991f
C362 B.n61 VSUBS 0.007991f
C363 B.n62 VSUBS 0.007991f
C364 B.n63 VSUBS 0.007991f
C365 B.n64 VSUBS 0.007991f
C366 B.n65 VSUBS 0.007991f
C367 B.n66 VSUBS 0.007991f
C368 B.n67 VSUBS 0.007991f
C369 B.n68 VSUBS 0.007991f
C370 B.n69 VSUBS 0.007991f
C371 B.n70 VSUBS 0.007991f
C372 B.n71 VSUBS 0.007991f
C373 B.n72 VSUBS 0.007991f
C374 B.n73 VSUBS 0.007991f
C375 B.n74 VSUBS 0.007991f
C376 B.n75 VSUBS 0.007991f
C377 B.n76 VSUBS 0.007991f
C378 B.n77 VSUBS 0.007991f
C379 B.n78 VSUBS 0.007991f
C380 B.n79 VSUBS 0.007991f
C381 B.n80 VSUBS 0.007991f
C382 B.n81 VSUBS 0.007991f
C383 B.n82 VSUBS 0.007991f
C384 B.n83 VSUBS 0.007991f
C385 B.n84 VSUBS 0.007991f
C386 B.n85 VSUBS 0.007991f
C387 B.n86 VSUBS 0.007991f
C388 B.n87 VSUBS 0.007991f
C389 B.n88 VSUBS 0.007991f
C390 B.n89 VSUBS 0.007991f
C391 B.n90 VSUBS 0.007991f
C392 B.n91 VSUBS 0.019661f
C393 B.n92 VSUBS 0.007991f
C394 B.n93 VSUBS 0.007991f
C395 B.n94 VSUBS 0.007991f
C396 B.n95 VSUBS 0.007991f
C397 B.n96 VSUBS 0.007991f
C398 B.n97 VSUBS 0.007991f
C399 B.t10 VSUBS 0.04577f
C400 B.t11 VSUBS 0.059647f
C401 B.t9 VSUBS 0.302104f
C402 B.n98 VSUBS 0.105481f
C403 B.n99 VSUBS 0.091496f
C404 B.n100 VSUBS 0.018513f
C405 B.n101 VSUBS 0.007991f
C406 B.n102 VSUBS 0.007991f
C407 B.n103 VSUBS 0.007991f
C408 B.n104 VSUBS 0.007991f
C409 B.n105 VSUBS 0.007991f
C410 B.t4 VSUBS 0.045769f
C411 B.t5 VSUBS 0.059647f
C412 B.t3 VSUBS 0.302104f
C413 B.n106 VSUBS 0.105481f
C414 B.n107 VSUBS 0.091496f
C415 B.n108 VSUBS 0.007991f
C416 B.n109 VSUBS 0.007991f
C417 B.n110 VSUBS 0.007991f
C418 B.n111 VSUBS 0.007991f
C419 B.n112 VSUBS 0.007991f
C420 B.n113 VSUBS 0.007991f
C421 B.n114 VSUBS 0.019116f
C422 B.n115 VSUBS 0.007991f
C423 B.n116 VSUBS 0.007991f
C424 B.n117 VSUBS 0.007991f
C425 B.n118 VSUBS 0.007991f
C426 B.n119 VSUBS 0.007991f
C427 B.n120 VSUBS 0.007991f
C428 B.n121 VSUBS 0.007991f
C429 B.n122 VSUBS 0.007991f
C430 B.n123 VSUBS 0.007991f
C431 B.n124 VSUBS 0.007991f
C432 B.n125 VSUBS 0.007991f
C433 B.n126 VSUBS 0.007991f
C434 B.n127 VSUBS 0.007991f
C435 B.n128 VSUBS 0.007991f
C436 B.n129 VSUBS 0.007991f
C437 B.n130 VSUBS 0.007991f
C438 B.n131 VSUBS 0.007991f
C439 B.n132 VSUBS 0.007991f
C440 B.n133 VSUBS 0.007991f
C441 B.n134 VSUBS 0.007991f
C442 B.n135 VSUBS 0.007991f
C443 B.n136 VSUBS 0.007991f
C444 B.n137 VSUBS 0.007991f
C445 B.n138 VSUBS 0.007991f
C446 B.n139 VSUBS 0.007991f
C447 B.n140 VSUBS 0.007991f
C448 B.n141 VSUBS 0.007991f
C449 B.n142 VSUBS 0.007991f
C450 B.n143 VSUBS 0.007991f
C451 B.n144 VSUBS 0.007991f
C452 B.n145 VSUBS 0.007991f
C453 B.n146 VSUBS 0.007991f
C454 B.n147 VSUBS 0.007991f
C455 B.n148 VSUBS 0.007991f
C456 B.n149 VSUBS 0.007991f
C457 B.n150 VSUBS 0.007991f
C458 B.n151 VSUBS 0.007991f
C459 B.n152 VSUBS 0.007991f
C460 B.n153 VSUBS 0.007991f
C461 B.n154 VSUBS 0.007991f
C462 B.n155 VSUBS 0.007991f
C463 B.n156 VSUBS 0.007991f
C464 B.n157 VSUBS 0.007991f
C465 B.n158 VSUBS 0.007991f
C466 B.n159 VSUBS 0.007991f
C467 B.n160 VSUBS 0.007991f
C468 B.n161 VSUBS 0.007991f
C469 B.n162 VSUBS 0.007991f
C470 B.n163 VSUBS 0.007991f
C471 B.n164 VSUBS 0.007991f
C472 B.n165 VSUBS 0.007991f
C473 B.n166 VSUBS 0.007991f
C474 B.n167 VSUBS 0.007991f
C475 B.n168 VSUBS 0.007991f
C476 B.n169 VSUBS 0.007991f
C477 B.n170 VSUBS 0.007991f
C478 B.n171 VSUBS 0.007991f
C479 B.n172 VSUBS 0.007991f
C480 B.n173 VSUBS 0.007991f
C481 B.n174 VSUBS 0.007991f
C482 B.n175 VSUBS 0.007991f
C483 B.n176 VSUBS 0.007991f
C484 B.n177 VSUBS 0.007991f
C485 B.n178 VSUBS 0.007991f
C486 B.n179 VSUBS 0.007991f
C487 B.n180 VSUBS 0.007991f
C488 B.n181 VSUBS 0.007991f
C489 B.n182 VSUBS 0.007991f
C490 B.n183 VSUBS 0.007991f
C491 B.n184 VSUBS 0.007991f
C492 B.n185 VSUBS 0.007991f
C493 B.n186 VSUBS 0.007991f
C494 B.n187 VSUBS 0.007991f
C495 B.n188 VSUBS 0.007991f
C496 B.n189 VSUBS 0.007991f
C497 B.n190 VSUBS 0.007991f
C498 B.n191 VSUBS 0.007991f
C499 B.n192 VSUBS 0.007991f
C500 B.n193 VSUBS 0.007991f
C501 B.n194 VSUBS 0.007991f
C502 B.n195 VSUBS 0.007991f
C503 B.n196 VSUBS 0.007991f
C504 B.n197 VSUBS 0.007991f
C505 B.n198 VSUBS 0.007991f
C506 B.n199 VSUBS 0.019116f
C507 B.n200 VSUBS 0.019661f
C508 B.n201 VSUBS 0.019661f
C509 B.n202 VSUBS 0.007991f
C510 B.n203 VSUBS 0.007991f
C511 B.n204 VSUBS 0.007991f
C512 B.n205 VSUBS 0.007991f
C513 B.n206 VSUBS 0.007991f
C514 B.n207 VSUBS 0.007991f
C515 B.n208 VSUBS 0.007991f
C516 B.n209 VSUBS 0.007991f
C517 B.n210 VSUBS 0.007991f
C518 B.n211 VSUBS 0.007991f
C519 B.n212 VSUBS 0.007991f
C520 B.n213 VSUBS 0.007991f
C521 B.n214 VSUBS 0.007991f
C522 B.n215 VSUBS 0.007991f
C523 B.n216 VSUBS 0.007991f
C524 B.n217 VSUBS 0.007991f
C525 B.n218 VSUBS 0.007991f
C526 B.n219 VSUBS 0.007991f
C527 B.n220 VSUBS 0.005523f
C528 B.n221 VSUBS 0.018513f
C529 B.n222 VSUBS 0.006463f
C530 B.n223 VSUBS 0.007991f
C531 B.n224 VSUBS 0.007991f
C532 B.n225 VSUBS 0.007991f
C533 B.n226 VSUBS 0.007991f
C534 B.n227 VSUBS 0.007991f
C535 B.n228 VSUBS 0.007991f
C536 B.n229 VSUBS 0.007991f
C537 B.n230 VSUBS 0.007991f
C538 B.n231 VSUBS 0.007991f
C539 B.n232 VSUBS 0.007991f
C540 B.n233 VSUBS 0.007991f
C541 B.n234 VSUBS 0.006463f
C542 B.n235 VSUBS 0.007991f
C543 B.n236 VSUBS 0.007991f
C544 B.n237 VSUBS 0.005523f
C545 B.n238 VSUBS 0.007991f
C546 B.n239 VSUBS 0.007991f
C547 B.n240 VSUBS 0.007991f
C548 B.n241 VSUBS 0.007991f
C549 B.n242 VSUBS 0.007991f
C550 B.n243 VSUBS 0.007991f
C551 B.n244 VSUBS 0.007991f
C552 B.n245 VSUBS 0.007991f
C553 B.n246 VSUBS 0.007991f
C554 B.n247 VSUBS 0.007991f
C555 B.n248 VSUBS 0.007991f
C556 B.n249 VSUBS 0.007991f
C557 B.n250 VSUBS 0.007991f
C558 B.n251 VSUBS 0.007991f
C559 B.n252 VSUBS 0.007991f
C560 B.n253 VSUBS 0.007991f
C561 B.n254 VSUBS 0.007991f
C562 B.n255 VSUBS 0.007991f
C563 B.n256 VSUBS 0.019661f
C564 B.n257 VSUBS 0.019116f
C565 B.n258 VSUBS 0.019116f
C566 B.n259 VSUBS 0.007991f
C567 B.n260 VSUBS 0.007991f
C568 B.n261 VSUBS 0.007991f
C569 B.n262 VSUBS 0.007991f
C570 B.n263 VSUBS 0.007991f
C571 B.n264 VSUBS 0.007991f
C572 B.n265 VSUBS 0.007991f
C573 B.n266 VSUBS 0.007991f
C574 B.n267 VSUBS 0.007991f
C575 B.n268 VSUBS 0.007991f
C576 B.n269 VSUBS 0.007991f
C577 B.n270 VSUBS 0.007991f
C578 B.n271 VSUBS 0.007991f
C579 B.n272 VSUBS 0.007991f
C580 B.n273 VSUBS 0.007991f
C581 B.n274 VSUBS 0.007991f
C582 B.n275 VSUBS 0.007991f
C583 B.n276 VSUBS 0.007991f
C584 B.n277 VSUBS 0.007991f
C585 B.n278 VSUBS 0.007991f
C586 B.n279 VSUBS 0.007991f
C587 B.n280 VSUBS 0.007991f
C588 B.n281 VSUBS 0.007991f
C589 B.n282 VSUBS 0.007991f
C590 B.n283 VSUBS 0.007991f
C591 B.n284 VSUBS 0.007991f
C592 B.n285 VSUBS 0.007991f
C593 B.n286 VSUBS 0.007991f
C594 B.n287 VSUBS 0.007991f
C595 B.n288 VSUBS 0.007991f
C596 B.n289 VSUBS 0.007991f
C597 B.n290 VSUBS 0.007991f
C598 B.n291 VSUBS 0.007991f
C599 B.n292 VSUBS 0.007991f
C600 B.n293 VSUBS 0.007991f
C601 B.n294 VSUBS 0.007991f
C602 B.n295 VSUBS 0.007991f
C603 B.n296 VSUBS 0.007991f
C604 B.n297 VSUBS 0.007991f
C605 B.n298 VSUBS 0.007991f
C606 B.n299 VSUBS 0.007991f
C607 B.n300 VSUBS 0.007991f
C608 B.n301 VSUBS 0.007991f
C609 B.n302 VSUBS 0.007991f
C610 B.n303 VSUBS 0.007991f
C611 B.n304 VSUBS 0.007991f
C612 B.n305 VSUBS 0.007991f
C613 B.n306 VSUBS 0.007991f
C614 B.n307 VSUBS 0.007991f
C615 B.n308 VSUBS 0.007991f
C616 B.n309 VSUBS 0.007991f
C617 B.n310 VSUBS 0.007991f
C618 B.n311 VSUBS 0.007991f
C619 B.n312 VSUBS 0.007991f
C620 B.n313 VSUBS 0.007991f
C621 B.n314 VSUBS 0.007991f
C622 B.n315 VSUBS 0.007991f
C623 B.n316 VSUBS 0.007991f
C624 B.n317 VSUBS 0.007991f
C625 B.n318 VSUBS 0.007991f
C626 B.n319 VSUBS 0.007991f
C627 B.n320 VSUBS 0.007991f
C628 B.n321 VSUBS 0.007991f
C629 B.n322 VSUBS 0.007991f
C630 B.n323 VSUBS 0.007991f
C631 B.n324 VSUBS 0.007991f
C632 B.n325 VSUBS 0.007991f
C633 B.n326 VSUBS 0.007991f
C634 B.n327 VSUBS 0.007991f
C635 B.n328 VSUBS 0.007991f
C636 B.n329 VSUBS 0.007991f
C637 B.n330 VSUBS 0.007991f
C638 B.n331 VSUBS 0.007991f
C639 B.n332 VSUBS 0.007991f
C640 B.n333 VSUBS 0.007991f
C641 B.n334 VSUBS 0.007991f
C642 B.n335 VSUBS 0.007991f
C643 B.n336 VSUBS 0.007991f
C644 B.n337 VSUBS 0.007991f
C645 B.n338 VSUBS 0.007991f
C646 B.n339 VSUBS 0.007991f
C647 B.n340 VSUBS 0.007991f
C648 B.n341 VSUBS 0.007991f
C649 B.n342 VSUBS 0.007991f
C650 B.n343 VSUBS 0.007991f
C651 B.n344 VSUBS 0.007991f
C652 B.n345 VSUBS 0.007991f
C653 B.n346 VSUBS 0.007991f
C654 B.n347 VSUBS 0.007991f
C655 B.n348 VSUBS 0.007991f
C656 B.n349 VSUBS 0.007991f
C657 B.n350 VSUBS 0.007991f
C658 B.n351 VSUBS 0.007991f
C659 B.n352 VSUBS 0.007991f
C660 B.n353 VSUBS 0.007991f
C661 B.n354 VSUBS 0.007991f
C662 B.n355 VSUBS 0.007991f
C663 B.n356 VSUBS 0.007991f
C664 B.n357 VSUBS 0.007991f
C665 B.n358 VSUBS 0.007991f
C666 B.n359 VSUBS 0.007991f
C667 B.n360 VSUBS 0.007991f
C668 B.n361 VSUBS 0.007991f
C669 B.n362 VSUBS 0.007991f
C670 B.n363 VSUBS 0.007991f
C671 B.n364 VSUBS 0.007991f
C672 B.n365 VSUBS 0.007991f
C673 B.n366 VSUBS 0.007991f
C674 B.n367 VSUBS 0.007991f
C675 B.n368 VSUBS 0.007991f
C676 B.n369 VSUBS 0.007991f
C677 B.n370 VSUBS 0.007991f
C678 B.n371 VSUBS 0.007991f
C679 B.n372 VSUBS 0.007991f
C680 B.n373 VSUBS 0.007991f
C681 B.n374 VSUBS 0.007991f
C682 B.n375 VSUBS 0.007991f
C683 B.n376 VSUBS 0.007991f
C684 B.n377 VSUBS 0.007991f
C685 B.n378 VSUBS 0.007991f
C686 B.n379 VSUBS 0.007991f
C687 B.n380 VSUBS 0.007991f
C688 B.n381 VSUBS 0.007991f
C689 B.n382 VSUBS 0.007991f
C690 B.n383 VSUBS 0.007991f
C691 B.n384 VSUBS 0.007991f
C692 B.n385 VSUBS 0.007991f
C693 B.n386 VSUBS 0.007991f
C694 B.n387 VSUBS 0.007991f
C695 B.n388 VSUBS 0.007991f
C696 B.n389 VSUBS 0.02001f
C697 B.n390 VSUBS 0.019116f
C698 B.n391 VSUBS 0.019661f
C699 B.n392 VSUBS 0.007991f
C700 B.n393 VSUBS 0.007991f
C701 B.n394 VSUBS 0.007991f
C702 B.n395 VSUBS 0.007991f
C703 B.n396 VSUBS 0.007991f
C704 B.n397 VSUBS 0.007991f
C705 B.n398 VSUBS 0.007991f
C706 B.n399 VSUBS 0.007991f
C707 B.n400 VSUBS 0.007991f
C708 B.n401 VSUBS 0.007991f
C709 B.n402 VSUBS 0.007991f
C710 B.n403 VSUBS 0.007991f
C711 B.n404 VSUBS 0.007991f
C712 B.n405 VSUBS 0.007991f
C713 B.n406 VSUBS 0.007991f
C714 B.n407 VSUBS 0.007991f
C715 B.n408 VSUBS 0.007991f
C716 B.n409 VSUBS 0.007991f
C717 B.n410 VSUBS 0.007991f
C718 B.n411 VSUBS 0.005523f
C719 B.n412 VSUBS 0.018513f
C720 B.n413 VSUBS 0.006463f
C721 B.n414 VSUBS 0.007991f
C722 B.n415 VSUBS 0.007991f
C723 B.n416 VSUBS 0.007991f
C724 B.n417 VSUBS 0.007991f
C725 B.n418 VSUBS 0.007991f
C726 B.n419 VSUBS 0.007991f
C727 B.n420 VSUBS 0.007991f
C728 B.n421 VSUBS 0.007991f
C729 B.n422 VSUBS 0.007991f
C730 B.n423 VSUBS 0.007991f
C731 B.n424 VSUBS 0.007991f
C732 B.n425 VSUBS 0.006463f
C733 B.n426 VSUBS 0.018513f
C734 B.n427 VSUBS 0.005523f
C735 B.n428 VSUBS 0.007991f
C736 B.n429 VSUBS 0.007991f
C737 B.n430 VSUBS 0.007991f
C738 B.n431 VSUBS 0.007991f
C739 B.n432 VSUBS 0.007991f
C740 B.n433 VSUBS 0.007991f
C741 B.n434 VSUBS 0.007991f
C742 B.n435 VSUBS 0.007991f
C743 B.n436 VSUBS 0.007991f
C744 B.n437 VSUBS 0.007991f
C745 B.n438 VSUBS 0.007991f
C746 B.n439 VSUBS 0.007991f
C747 B.n440 VSUBS 0.007991f
C748 B.n441 VSUBS 0.007991f
C749 B.n442 VSUBS 0.007991f
C750 B.n443 VSUBS 0.007991f
C751 B.n444 VSUBS 0.007991f
C752 B.n445 VSUBS 0.007991f
C753 B.n446 VSUBS 0.007991f
C754 B.n447 VSUBS 0.019661f
C755 B.n448 VSUBS 0.019116f
C756 B.n449 VSUBS 0.019116f
C757 B.n450 VSUBS 0.007991f
C758 B.n451 VSUBS 0.007991f
C759 B.n452 VSUBS 0.007991f
C760 B.n453 VSUBS 0.007991f
C761 B.n454 VSUBS 0.007991f
C762 B.n455 VSUBS 0.007991f
C763 B.n456 VSUBS 0.007991f
C764 B.n457 VSUBS 0.007991f
C765 B.n458 VSUBS 0.007991f
C766 B.n459 VSUBS 0.007991f
C767 B.n460 VSUBS 0.007991f
C768 B.n461 VSUBS 0.007991f
C769 B.n462 VSUBS 0.007991f
C770 B.n463 VSUBS 0.007991f
C771 B.n464 VSUBS 0.007991f
C772 B.n465 VSUBS 0.007991f
C773 B.n466 VSUBS 0.007991f
C774 B.n467 VSUBS 0.007991f
C775 B.n468 VSUBS 0.007991f
C776 B.n469 VSUBS 0.007991f
C777 B.n470 VSUBS 0.007991f
C778 B.n471 VSUBS 0.007991f
C779 B.n472 VSUBS 0.007991f
C780 B.n473 VSUBS 0.007991f
C781 B.n474 VSUBS 0.007991f
C782 B.n475 VSUBS 0.007991f
C783 B.n476 VSUBS 0.007991f
C784 B.n477 VSUBS 0.007991f
C785 B.n478 VSUBS 0.007991f
C786 B.n479 VSUBS 0.007991f
C787 B.n480 VSUBS 0.007991f
C788 B.n481 VSUBS 0.007991f
C789 B.n482 VSUBS 0.007991f
C790 B.n483 VSUBS 0.007991f
C791 B.n484 VSUBS 0.007991f
C792 B.n485 VSUBS 0.007991f
C793 B.n486 VSUBS 0.007991f
C794 B.n487 VSUBS 0.007991f
C795 B.n488 VSUBS 0.007991f
C796 B.n489 VSUBS 0.007991f
C797 B.n490 VSUBS 0.007991f
C798 B.n491 VSUBS 0.007991f
C799 B.n492 VSUBS 0.007991f
C800 B.n493 VSUBS 0.007991f
C801 B.n494 VSUBS 0.007991f
C802 B.n495 VSUBS 0.007991f
C803 B.n496 VSUBS 0.007991f
C804 B.n497 VSUBS 0.007991f
C805 B.n498 VSUBS 0.007991f
C806 B.n499 VSUBS 0.007991f
C807 B.n500 VSUBS 0.007991f
C808 B.n501 VSUBS 0.007991f
C809 B.n502 VSUBS 0.007991f
C810 B.n503 VSUBS 0.007991f
C811 B.n504 VSUBS 0.007991f
C812 B.n505 VSUBS 0.007991f
C813 B.n506 VSUBS 0.007991f
C814 B.n507 VSUBS 0.007991f
C815 B.n508 VSUBS 0.007991f
C816 B.n509 VSUBS 0.007991f
C817 B.n510 VSUBS 0.007991f
C818 B.n511 VSUBS 0.007991f
C819 B.n512 VSUBS 0.007991f
C820 B.n513 VSUBS 0.007991f
C821 B.n514 VSUBS 0.007991f
C822 B.n515 VSUBS 0.018093f
.ends

