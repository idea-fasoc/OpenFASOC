* NGSPICE file created from diff_pair_sample_0629.ext - technology: sky130A

.subckt diff_pair_sample_0629 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=3.2955 ps=17.68 w=8.45 l=1.62
X1 VDD1.t9 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X2 VTAIL.t2 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X3 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=0 ps=0 w=8.45 l=1.62
X4 VTAIL.t11 VN.t1 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X5 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=0 ps=0 w=8.45 l=1.62
X6 VDD1.t7 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=3.2955 ps=17.68 w=8.45 l=1.62
X7 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=0 ps=0 w=8.45 l=1.62
X8 VDD2.t7 VN.t2 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X9 VTAIL.t18 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X10 VDD2.t5 VN.t4 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=3.2955 ps=17.68 w=8.45 l=1.62
X11 VDD2.t4 VN.t5 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=1.39425 ps=8.78 w=8.45 l=1.62
X12 VDD1.t6 VP.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=1.39425 ps=8.78 w=8.45 l=1.62
X13 VTAIL.t10 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X14 VDD1.t5 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=3.2955 ps=17.68 w=8.45 l=1.62
X15 VDD2.t2 VN.t7 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X16 VTAIL.t7 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X17 VDD1.t3 VP.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=1.39425 ps=8.78 w=8.45 l=1.62
X18 VDD1.t2 VP.t7 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=0 ps=0 w=8.45 l=1.62
X20 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X21 VTAIL.t12 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X22 VTAIL.t0 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.39425 pd=8.78 as=1.39425 ps=8.78 w=8.45 l=1.62
X23 VDD2.t0 VN.t9 VTAIL.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=3.2955 pd=17.68 as=1.39425 ps=8.78 w=8.45 l=1.62
R0 VN.n29 VN.n28 178.428
R1 VN.n59 VN.n58 178.428
R2 VN.n57 VN.n30 161.3
R3 VN.n56 VN.n55 161.3
R4 VN.n54 VN.n31 161.3
R5 VN.n53 VN.n52 161.3
R6 VN.n50 VN.n32 161.3
R7 VN.n49 VN.n48 161.3
R8 VN.n47 VN.n33 161.3
R9 VN.n46 VN.n45 161.3
R10 VN.n43 VN.n34 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n35 161.3
R13 VN.n39 VN.n38 161.3
R14 VN.n27 VN.n0 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n1 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n20 VN.n2 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n3 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n13 VN.n4 161.3
R23 VN.n12 VN.n11 161.3
R24 VN.n10 VN.n5 161.3
R25 VN.n9 VN.n8 161.3
R26 VN.n6 VN.t5 158.025
R27 VN.n36 VN.t4 158.025
R28 VN.n7 VN.t3 125.707
R29 VN.n14 VN.t2 125.707
R30 VN.n21 VN.t1 125.707
R31 VN.n28 VN.t0 125.707
R32 VN.n37 VN.t6 125.707
R33 VN.n44 VN.t7 125.707
R34 VN.n51 VN.t8 125.707
R35 VN.n58 VN.t9 125.707
R36 VN.n12 VN.n5 56.5193
R37 VN.n19 VN.n3 56.5193
R38 VN.n26 VN.n1 56.5193
R39 VN.n42 VN.n35 56.5193
R40 VN.n49 VN.n33 56.5193
R41 VN.n56 VN.n31 56.5193
R42 VN.n7 VN.n6 56.3226
R43 VN.n37 VN.n36 56.3226
R44 VN VN.n59 45.3925
R45 VN.n8 VN.n5 24.4675
R46 VN.n13 VN.n12 24.4675
R47 VN.n15 VN.n3 24.4675
R48 VN.n20 VN.n19 24.4675
R49 VN.n22 VN.n1 24.4675
R50 VN.n27 VN.n26 24.4675
R51 VN.n38 VN.n35 24.4675
R52 VN.n45 VN.n33 24.4675
R53 VN.n43 VN.n42 24.4675
R54 VN.n52 VN.n31 24.4675
R55 VN.n50 VN.n49 24.4675
R56 VN.n57 VN.n56 24.4675
R57 VN.n39 VN.n36 18.0474
R58 VN.n9 VN.n6 18.0474
R59 VN.n22 VN.n21 14.6807
R60 VN.n52 VN.n51 14.6807
R61 VN.n14 VN.n13 12.234
R62 VN.n15 VN.n14 12.234
R63 VN.n45 VN.n44 12.234
R64 VN.n44 VN.n43 12.234
R65 VN.n8 VN.n7 9.7873
R66 VN.n21 VN.n20 9.7873
R67 VN.n38 VN.n37 9.7873
R68 VN.n51 VN.n50 9.7873
R69 VN.n28 VN.n27 7.3406
R70 VN.n58 VN.n57 7.3406
R71 VN.n59 VN.n30 0.189894
R72 VN.n55 VN.n30 0.189894
R73 VN.n55 VN.n54 0.189894
R74 VN.n54 VN.n53 0.189894
R75 VN.n53 VN.n32 0.189894
R76 VN.n48 VN.n32 0.189894
R77 VN.n48 VN.n47 0.189894
R78 VN.n47 VN.n46 0.189894
R79 VN.n46 VN.n34 0.189894
R80 VN.n41 VN.n34 0.189894
R81 VN.n41 VN.n40 0.189894
R82 VN.n40 VN.n39 0.189894
R83 VN.n10 VN.n9 0.189894
R84 VN.n11 VN.n10 0.189894
R85 VN.n11 VN.n4 0.189894
R86 VN.n16 VN.n4 0.189894
R87 VN.n17 VN.n16 0.189894
R88 VN.n18 VN.n17 0.189894
R89 VN.n18 VN.n2 0.189894
R90 VN.n23 VN.n2 0.189894
R91 VN.n24 VN.n23 0.189894
R92 VN.n25 VN.n24 0.189894
R93 VN.n25 VN.n0 0.189894
R94 VN.n29 VN.n0 0.189894
R95 VN VN.n29 0.0516364
R96 VTAIL.n11 VTAIL.t17 48.5129
R97 VTAIL.n16 VTAIL.t3 48.5129
R98 VTAIL.n17 VTAIL.t16 48.5127
R99 VTAIL.n2 VTAIL.t4 48.5127
R100 VTAIL.n15 VTAIL.n14 46.1697
R101 VTAIL.n13 VTAIL.n12 46.1697
R102 VTAIL.n10 VTAIL.n9 46.1697
R103 VTAIL.n8 VTAIL.n7 46.1697
R104 VTAIL.n19 VTAIL.n18 46.1697
R105 VTAIL.n1 VTAIL.n0 46.1697
R106 VTAIL.n4 VTAIL.n3 46.1697
R107 VTAIL.n6 VTAIL.n5 46.1697
R108 VTAIL.n8 VTAIL.n6 23.0134
R109 VTAIL.n17 VTAIL.n16 21.3324
R110 VTAIL.n18 VTAIL.t15 2.3437
R111 VTAIL.n18 VTAIL.t11 2.3437
R112 VTAIL.n0 VTAIL.t13 2.3437
R113 VTAIL.n0 VTAIL.t18 2.3437
R114 VTAIL.n3 VTAIL.t6 2.3437
R115 VTAIL.n3 VTAIL.t2 2.3437
R116 VTAIL.n5 VTAIL.t8 2.3437
R117 VTAIL.n5 VTAIL.t7 2.3437
R118 VTAIL.n14 VTAIL.t19 2.3437
R119 VTAIL.n14 VTAIL.t0 2.3437
R120 VTAIL.n12 VTAIL.t5 2.3437
R121 VTAIL.n12 VTAIL.t1 2.3437
R122 VTAIL.n9 VTAIL.t14 2.3437
R123 VTAIL.n9 VTAIL.t10 2.3437
R124 VTAIL.n7 VTAIL.t9 2.3437
R125 VTAIL.n7 VTAIL.t12 2.3437
R126 VTAIL.n10 VTAIL.n8 1.68153
R127 VTAIL.n11 VTAIL.n10 1.68153
R128 VTAIL.n15 VTAIL.n13 1.68153
R129 VTAIL.n16 VTAIL.n15 1.68153
R130 VTAIL.n6 VTAIL.n4 1.68153
R131 VTAIL.n4 VTAIL.n2 1.68153
R132 VTAIL.n19 VTAIL.n17 1.68153
R133 VTAIL VTAIL.n1 1.31947
R134 VTAIL.n13 VTAIL.n11 1.31084
R135 VTAIL.n2 VTAIL.n1 1.31084
R136 VTAIL VTAIL.n19 0.362569
R137 VDD2.n1 VDD2.t4 66.8725
R138 VDD2.n4 VDD2.t0 65.1917
R139 VDD2.n3 VDD2.n2 64.0539
R140 VDD2 VDD2.n7 64.0511
R141 VDD2.n6 VDD2.n5 62.8485
R142 VDD2.n1 VDD2.n0 62.8485
R143 VDD2.n4 VDD2.n3 38.9847
R144 VDD2.n7 VDD2.t3 2.3437
R145 VDD2.n7 VDD2.t5 2.3437
R146 VDD2.n5 VDD2.t1 2.3437
R147 VDD2.n5 VDD2.t2 2.3437
R148 VDD2.n2 VDD2.t8 2.3437
R149 VDD2.n2 VDD2.t9 2.3437
R150 VDD2.n0 VDD2.t6 2.3437
R151 VDD2.n0 VDD2.t7 2.3437
R152 VDD2.n6 VDD2.n4 1.68153
R153 VDD2 VDD2.n6 0.478948
R154 VDD2.n3 VDD2.n1 0.365413
R155 B.n570 B.n569 585
R156 B.n572 B.n119 585
R157 B.n575 B.n574 585
R158 B.n576 B.n118 585
R159 B.n578 B.n577 585
R160 B.n580 B.n117 585
R161 B.n583 B.n582 585
R162 B.n584 B.n116 585
R163 B.n586 B.n585 585
R164 B.n588 B.n115 585
R165 B.n591 B.n590 585
R166 B.n592 B.n114 585
R167 B.n594 B.n593 585
R168 B.n596 B.n113 585
R169 B.n599 B.n598 585
R170 B.n600 B.n112 585
R171 B.n602 B.n601 585
R172 B.n604 B.n111 585
R173 B.n607 B.n606 585
R174 B.n608 B.n110 585
R175 B.n610 B.n609 585
R176 B.n612 B.n109 585
R177 B.n615 B.n614 585
R178 B.n616 B.n108 585
R179 B.n618 B.n617 585
R180 B.n620 B.n107 585
R181 B.n623 B.n622 585
R182 B.n624 B.n106 585
R183 B.n626 B.n625 585
R184 B.n628 B.n105 585
R185 B.n631 B.n630 585
R186 B.n633 B.n102 585
R187 B.n635 B.n634 585
R188 B.n637 B.n101 585
R189 B.n640 B.n639 585
R190 B.n641 B.n100 585
R191 B.n643 B.n642 585
R192 B.n645 B.n99 585
R193 B.n648 B.n647 585
R194 B.n649 B.n95 585
R195 B.n651 B.n650 585
R196 B.n653 B.n94 585
R197 B.n656 B.n655 585
R198 B.n657 B.n93 585
R199 B.n659 B.n658 585
R200 B.n661 B.n92 585
R201 B.n664 B.n663 585
R202 B.n665 B.n91 585
R203 B.n667 B.n666 585
R204 B.n669 B.n90 585
R205 B.n672 B.n671 585
R206 B.n673 B.n89 585
R207 B.n675 B.n674 585
R208 B.n677 B.n88 585
R209 B.n680 B.n679 585
R210 B.n681 B.n87 585
R211 B.n683 B.n682 585
R212 B.n685 B.n86 585
R213 B.n688 B.n687 585
R214 B.n689 B.n85 585
R215 B.n691 B.n690 585
R216 B.n693 B.n84 585
R217 B.n696 B.n695 585
R218 B.n697 B.n83 585
R219 B.n699 B.n698 585
R220 B.n701 B.n82 585
R221 B.n704 B.n703 585
R222 B.n705 B.n81 585
R223 B.n707 B.n706 585
R224 B.n709 B.n80 585
R225 B.n712 B.n711 585
R226 B.n713 B.n79 585
R227 B.n568 B.n77 585
R228 B.n716 B.n77 585
R229 B.n567 B.n76 585
R230 B.n717 B.n76 585
R231 B.n566 B.n75 585
R232 B.n718 B.n75 585
R233 B.n565 B.n564 585
R234 B.n564 B.n71 585
R235 B.n563 B.n70 585
R236 B.n724 B.n70 585
R237 B.n562 B.n69 585
R238 B.n725 B.n69 585
R239 B.n561 B.n68 585
R240 B.n726 B.n68 585
R241 B.n560 B.n559 585
R242 B.n559 B.n64 585
R243 B.n558 B.n63 585
R244 B.n732 B.n63 585
R245 B.n557 B.n62 585
R246 B.n733 B.n62 585
R247 B.n556 B.n61 585
R248 B.n734 B.n61 585
R249 B.n555 B.n554 585
R250 B.n554 B.n57 585
R251 B.n553 B.n56 585
R252 B.n740 B.n56 585
R253 B.n552 B.n55 585
R254 B.n741 B.n55 585
R255 B.n551 B.n54 585
R256 B.n742 B.n54 585
R257 B.n550 B.n549 585
R258 B.n549 B.n53 585
R259 B.n548 B.n49 585
R260 B.n748 B.n49 585
R261 B.n547 B.n48 585
R262 B.n749 B.n48 585
R263 B.n546 B.n47 585
R264 B.n750 B.n47 585
R265 B.n545 B.n544 585
R266 B.n544 B.n43 585
R267 B.n543 B.n42 585
R268 B.n756 B.n42 585
R269 B.n542 B.n41 585
R270 B.n757 B.n41 585
R271 B.n541 B.n40 585
R272 B.n758 B.n40 585
R273 B.n540 B.n539 585
R274 B.n539 B.n36 585
R275 B.n538 B.n35 585
R276 B.n764 B.n35 585
R277 B.n537 B.n34 585
R278 B.n765 B.n34 585
R279 B.n536 B.n33 585
R280 B.n766 B.n33 585
R281 B.n535 B.n534 585
R282 B.n534 B.n29 585
R283 B.n533 B.n28 585
R284 B.n772 B.n28 585
R285 B.n532 B.n27 585
R286 B.n773 B.n27 585
R287 B.n531 B.n26 585
R288 B.n774 B.n26 585
R289 B.n530 B.n529 585
R290 B.n529 B.n22 585
R291 B.n528 B.n21 585
R292 B.n780 B.n21 585
R293 B.n527 B.n20 585
R294 B.n781 B.n20 585
R295 B.n526 B.n19 585
R296 B.n782 B.n19 585
R297 B.n525 B.n524 585
R298 B.n524 B.n15 585
R299 B.n523 B.n14 585
R300 B.n788 B.n14 585
R301 B.n522 B.n13 585
R302 B.n789 B.n13 585
R303 B.n521 B.n12 585
R304 B.n790 B.n12 585
R305 B.n520 B.n519 585
R306 B.n519 B.n518 585
R307 B.n517 B.n516 585
R308 B.n517 B.n8 585
R309 B.n515 B.n7 585
R310 B.n797 B.n7 585
R311 B.n514 B.n6 585
R312 B.n798 B.n6 585
R313 B.n513 B.n5 585
R314 B.n799 B.n5 585
R315 B.n512 B.n511 585
R316 B.n511 B.n4 585
R317 B.n510 B.n120 585
R318 B.n510 B.n509 585
R319 B.n500 B.n121 585
R320 B.n122 B.n121 585
R321 B.n502 B.n501 585
R322 B.n503 B.n502 585
R323 B.n499 B.n127 585
R324 B.n127 B.n126 585
R325 B.n498 B.n497 585
R326 B.n497 B.n496 585
R327 B.n129 B.n128 585
R328 B.n130 B.n129 585
R329 B.n489 B.n488 585
R330 B.n490 B.n489 585
R331 B.n487 B.n135 585
R332 B.n135 B.n134 585
R333 B.n486 B.n485 585
R334 B.n485 B.n484 585
R335 B.n137 B.n136 585
R336 B.n138 B.n137 585
R337 B.n477 B.n476 585
R338 B.n478 B.n477 585
R339 B.n475 B.n143 585
R340 B.n143 B.n142 585
R341 B.n474 B.n473 585
R342 B.n473 B.n472 585
R343 B.n145 B.n144 585
R344 B.n146 B.n145 585
R345 B.n465 B.n464 585
R346 B.n466 B.n465 585
R347 B.n463 B.n151 585
R348 B.n151 B.n150 585
R349 B.n462 B.n461 585
R350 B.n461 B.n460 585
R351 B.n153 B.n152 585
R352 B.n154 B.n153 585
R353 B.n453 B.n452 585
R354 B.n454 B.n453 585
R355 B.n451 B.n159 585
R356 B.n159 B.n158 585
R357 B.n450 B.n449 585
R358 B.n449 B.n448 585
R359 B.n161 B.n160 585
R360 B.n162 B.n161 585
R361 B.n441 B.n440 585
R362 B.n442 B.n441 585
R363 B.n439 B.n167 585
R364 B.n167 B.n166 585
R365 B.n438 B.n437 585
R366 B.n437 B.n436 585
R367 B.n169 B.n168 585
R368 B.n429 B.n169 585
R369 B.n428 B.n427 585
R370 B.n430 B.n428 585
R371 B.n426 B.n174 585
R372 B.n174 B.n173 585
R373 B.n425 B.n424 585
R374 B.n424 B.n423 585
R375 B.n176 B.n175 585
R376 B.n177 B.n176 585
R377 B.n416 B.n415 585
R378 B.n417 B.n416 585
R379 B.n414 B.n182 585
R380 B.n182 B.n181 585
R381 B.n413 B.n412 585
R382 B.n412 B.n411 585
R383 B.n184 B.n183 585
R384 B.n185 B.n184 585
R385 B.n404 B.n403 585
R386 B.n405 B.n404 585
R387 B.n402 B.n190 585
R388 B.n190 B.n189 585
R389 B.n401 B.n400 585
R390 B.n400 B.n399 585
R391 B.n192 B.n191 585
R392 B.n193 B.n192 585
R393 B.n392 B.n391 585
R394 B.n393 B.n392 585
R395 B.n390 B.n198 585
R396 B.n198 B.n197 585
R397 B.n389 B.n388 585
R398 B.n388 B.n387 585
R399 B.n384 B.n202 585
R400 B.n383 B.n382 585
R401 B.n380 B.n203 585
R402 B.n380 B.n201 585
R403 B.n379 B.n378 585
R404 B.n377 B.n376 585
R405 B.n375 B.n205 585
R406 B.n373 B.n372 585
R407 B.n371 B.n206 585
R408 B.n370 B.n369 585
R409 B.n367 B.n207 585
R410 B.n365 B.n364 585
R411 B.n363 B.n208 585
R412 B.n362 B.n361 585
R413 B.n359 B.n209 585
R414 B.n357 B.n356 585
R415 B.n355 B.n210 585
R416 B.n354 B.n353 585
R417 B.n351 B.n211 585
R418 B.n349 B.n348 585
R419 B.n347 B.n212 585
R420 B.n346 B.n345 585
R421 B.n343 B.n213 585
R422 B.n341 B.n340 585
R423 B.n339 B.n214 585
R424 B.n338 B.n337 585
R425 B.n335 B.n215 585
R426 B.n333 B.n332 585
R427 B.n331 B.n216 585
R428 B.n330 B.n329 585
R429 B.n327 B.n217 585
R430 B.n325 B.n324 585
R431 B.n322 B.n218 585
R432 B.n321 B.n320 585
R433 B.n318 B.n221 585
R434 B.n316 B.n315 585
R435 B.n314 B.n222 585
R436 B.n313 B.n312 585
R437 B.n310 B.n223 585
R438 B.n308 B.n307 585
R439 B.n306 B.n224 585
R440 B.n305 B.n304 585
R441 B.n302 B.n301 585
R442 B.n300 B.n299 585
R443 B.n298 B.n229 585
R444 B.n296 B.n295 585
R445 B.n294 B.n230 585
R446 B.n293 B.n292 585
R447 B.n290 B.n231 585
R448 B.n288 B.n287 585
R449 B.n286 B.n232 585
R450 B.n285 B.n284 585
R451 B.n282 B.n233 585
R452 B.n280 B.n279 585
R453 B.n278 B.n234 585
R454 B.n277 B.n276 585
R455 B.n274 B.n235 585
R456 B.n272 B.n271 585
R457 B.n270 B.n236 585
R458 B.n269 B.n268 585
R459 B.n266 B.n237 585
R460 B.n264 B.n263 585
R461 B.n262 B.n238 585
R462 B.n261 B.n260 585
R463 B.n258 B.n239 585
R464 B.n256 B.n255 585
R465 B.n254 B.n240 585
R466 B.n253 B.n252 585
R467 B.n250 B.n241 585
R468 B.n248 B.n247 585
R469 B.n246 B.n242 585
R470 B.n245 B.n244 585
R471 B.n200 B.n199 585
R472 B.n201 B.n200 585
R473 B.n386 B.n385 585
R474 B.n387 B.n386 585
R475 B.n196 B.n195 585
R476 B.n197 B.n196 585
R477 B.n395 B.n394 585
R478 B.n394 B.n393 585
R479 B.n396 B.n194 585
R480 B.n194 B.n193 585
R481 B.n398 B.n397 585
R482 B.n399 B.n398 585
R483 B.n188 B.n187 585
R484 B.n189 B.n188 585
R485 B.n407 B.n406 585
R486 B.n406 B.n405 585
R487 B.n408 B.n186 585
R488 B.n186 B.n185 585
R489 B.n410 B.n409 585
R490 B.n411 B.n410 585
R491 B.n180 B.n179 585
R492 B.n181 B.n180 585
R493 B.n419 B.n418 585
R494 B.n418 B.n417 585
R495 B.n420 B.n178 585
R496 B.n178 B.n177 585
R497 B.n422 B.n421 585
R498 B.n423 B.n422 585
R499 B.n172 B.n171 585
R500 B.n173 B.n172 585
R501 B.n432 B.n431 585
R502 B.n431 B.n430 585
R503 B.n433 B.n170 585
R504 B.n429 B.n170 585
R505 B.n435 B.n434 585
R506 B.n436 B.n435 585
R507 B.n165 B.n164 585
R508 B.n166 B.n165 585
R509 B.n444 B.n443 585
R510 B.n443 B.n442 585
R511 B.n445 B.n163 585
R512 B.n163 B.n162 585
R513 B.n447 B.n446 585
R514 B.n448 B.n447 585
R515 B.n157 B.n156 585
R516 B.n158 B.n157 585
R517 B.n456 B.n455 585
R518 B.n455 B.n454 585
R519 B.n457 B.n155 585
R520 B.n155 B.n154 585
R521 B.n459 B.n458 585
R522 B.n460 B.n459 585
R523 B.n149 B.n148 585
R524 B.n150 B.n149 585
R525 B.n468 B.n467 585
R526 B.n467 B.n466 585
R527 B.n469 B.n147 585
R528 B.n147 B.n146 585
R529 B.n471 B.n470 585
R530 B.n472 B.n471 585
R531 B.n141 B.n140 585
R532 B.n142 B.n141 585
R533 B.n480 B.n479 585
R534 B.n479 B.n478 585
R535 B.n481 B.n139 585
R536 B.n139 B.n138 585
R537 B.n483 B.n482 585
R538 B.n484 B.n483 585
R539 B.n133 B.n132 585
R540 B.n134 B.n133 585
R541 B.n492 B.n491 585
R542 B.n491 B.n490 585
R543 B.n493 B.n131 585
R544 B.n131 B.n130 585
R545 B.n495 B.n494 585
R546 B.n496 B.n495 585
R547 B.n125 B.n124 585
R548 B.n126 B.n125 585
R549 B.n505 B.n504 585
R550 B.n504 B.n503 585
R551 B.n506 B.n123 585
R552 B.n123 B.n122 585
R553 B.n508 B.n507 585
R554 B.n509 B.n508 585
R555 B.n3 B.n0 585
R556 B.n4 B.n3 585
R557 B.n796 B.n1 585
R558 B.n797 B.n796 585
R559 B.n795 B.n794 585
R560 B.n795 B.n8 585
R561 B.n793 B.n9 585
R562 B.n518 B.n9 585
R563 B.n792 B.n791 585
R564 B.n791 B.n790 585
R565 B.n11 B.n10 585
R566 B.n789 B.n11 585
R567 B.n787 B.n786 585
R568 B.n788 B.n787 585
R569 B.n785 B.n16 585
R570 B.n16 B.n15 585
R571 B.n784 B.n783 585
R572 B.n783 B.n782 585
R573 B.n18 B.n17 585
R574 B.n781 B.n18 585
R575 B.n779 B.n778 585
R576 B.n780 B.n779 585
R577 B.n777 B.n23 585
R578 B.n23 B.n22 585
R579 B.n776 B.n775 585
R580 B.n775 B.n774 585
R581 B.n25 B.n24 585
R582 B.n773 B.n25 585
R583 B.n771 B.n770 585
R584 B.n772 B.n771 585
R585 B.n769 B.n30 585
R586 B.n30 B.n29 585
R587 B.n768 B.n767 585
R588 B.n767 B.n766 585
R589 B.n32 B.n31 585
R590 B.n765 B.n32 585
R591 B.n763 B.n762 585
R592 B.n764 B.n763 585
R593 B.n761 B.n37 585
R594 B.n37 B.n36 585
R595 B.n760 B.n759 585
R596 B.n759 B.n758 585
R597 B.n39 B.n38 585
R598 B.n757 B.n39 585
R599 B.n755 B.n754 585
R600 B.n756 B.n755 585
R601 B.n753 B.n44 585
R602 B.n44 B.n43 585
R603 B.n752 B.n751 585
R604 B.n751 B.n750 585
R605 B.n46 B.n45 585
R606 B.n749 B.n46 585
R607 B.n747 B.n746 585
R608 B.n748 B.n747 585
R609 B.n745 B.n50 585
R610 B.n53 B.n50 585
R611 B.n744 B.n743 585
R612 B.n743 B.n742 585
R613 B.n52 B.n51 585
R614 B.n741 B.n52 585
R615 B.n739 B.n738 585
R616 B.n740 B.n739 585
R617 B.n737 B.n58 585
R618 B.n58 B.n57 585
R619 B.n736 B.n735 585
R620 B.n735 B.n734 585
R621 B.n60 B.n59 585
R622 B.n733 B.n60 585
R623 B.n731 B.n730 585
R624 B.n732 B.n731 585
R625 B.n729 B.n65 585
R626 B.n65 B.n64 585
R627 B.n728 B.n727 585
R628 B.n727 B.n726 585
R629 B.n67 B.n66 585
R630 B.n725 B.n67 585
R631 B.n723 B.n722 585
R632 B.n724 B.n723 585
R633 B.n721 B.n72 585
R634 B.n72 B.n71 585
R635 B.n720 B.n719 585
R636 B.n719 B.n718 585
R637 B.n74 B.n73 585
R638 B.n717 B.n74 585
R639 B.n715 B.n714 585
R640 B.n716 B.n715 585
R641 B.n800 B.n799 585
R642 B.n798 B.n2 585
R643 B.n715 B.n79 497.305
R644 B.n570 B.n77 497.305
R645 B.n388 B.n200 497.305
R646 B.n386 B.n202 497.305
R647 B.n96 B.t18 331.567
R648 B.n103 B.t10 331.567
R649 B.n225 B.t14 331.567
R650 B.n219 B.t21 331.567
R651 B.n571 B.n78 256.663
R652 B.n573 B.n78 256.663
R653 B.n579 B.n78 256.663
R654 B.n581 B.n78 256.663
R655 B.n587 B.n78 256.663
R656 B.n589 B.n78 256.663
R657 B.n595 B.n78 256.663
R658 B.n597 B.n78 256.663
R659 B.n603 B.n78 256.663
R660 B.n605 B.n78 256.663
R661 B.n611 B.n78 256.663
R662 B.n613 B.n78 256.663
R663 B.n619 B.n78 256.663
R664 B.n621 B.n78 256.663
R665 B.n627 B.n78 256.663
R666 B.n629 B.n78 256.663
R667 B.n636 B.n78 256.663
R668 B.n638 B.n78 256.663
R669 B.n644 B.n78 256.663
R670 B.n646 B.n78 256.663
R671 B.n652 B.n78 256.663
R672 B.n654 B.n78 256.663
R673 B.n660 B.n78 256.663
R674 B.n662 B.n78 256.663
R675 B.n668 B.n78 256.663
R676 B.n670 B.n78 256.663
R677 B.n676 B.n78 256.663
R678 B.n678 B.n78 256.663
R679 B.n684 B.n78 256.663
R680 B.n686 B.n78 256.663
R681 B.n692 B.n78 256.663
R682 B.n694 B.n78 256.663
R683 B.n700 B.n78 256.663
R684 B.n702 B.n78 256.663
R685 B.n708 B.n78 256.663
R686 B.n710 B.n78 256.663
R687 B.n381 B.n201 256.663
R688 B.n204 B.n201 256.663
R689 B.n374 B.n201 256.663
R690 B.n368 B.n201 256.663
R691 B.n366 B.n201 256.663
R692 B.n360 B.n201 256.663
R693 B.n358 B.n201 256.663
R694 B.n352 B.n201 256.663
R695 B.n350 B.n201 256.663
R696 B.n344 B.n201 256.663
R697 B.n342 B.n201 256.663
R698 B.n336 B.n201 256.663
R699 B.n334 B.n201 256.663
R700 B.n328 B.n201 256.663
R701 B.n326 B.n201 256.663
R702 B.n319 B.n201 256.663
R703 B.n317 B.n201 256.663
R704 B.n311 B.n201 256.663
R705 B.n309 B.n201 256.663
R706 B.n303 B.n201 256.663
R707 B.n228 B.n201 256.663
R708 B.n297 B.n201 256.663
R709 B.n291 B.n201 256.663
R710 B.n289 B.n201 256.663
R711 B.n283 B.n201 256.663
R712 B.n281 B.n201 256.663
R713 B.n275 B.n201 256.663
R714 B.n273 B.n201 256.663
R715 B.n267 B.n201 256.663
R716 B.n265 B.n201 256.663
R717 B.n259 B.n201 256.663
R718 B.n257 B.n201 256.663
R719 B.n251 B.n201 256.663
R720 B.n249 B.n201 256.663
R721 B.n243 B.n201 256.663
R722 B.n802 B.n801 256.663
R723 B.n711 B.n709 163.367
R724 B.n707 B.n81 163.367
R725 B.n703 B.n701 163.367
R726 B.n699 B.n83 163.367
R727 B.n695 B.n693 163.367
R728 B.n691 B.n85 163.367
R729 B.n687 B.n685 163.367
R730 B.n683 B.n87 163.367
R731 B.n679 B.n677 163.367
R732 B.n675 B.n89 163.367
R733 B.n671 B.n669 163.367
R734 B.n667 B.n91 163.367
R735 B.n663 B.n661 163.367
R736 B.n659 B.n93 163.367
R737 B.n655 B.n653 163.367
R738 B.n651 B.n95 163.367
R739 B.n647 B.n645 163.367
R740 B.n643 B.n100 163.367
R741 B.n639 B.n637 163.367
R742 B.n635 B.n102 163.367
R743 B.n630 B.n628 163.367
R744 B.n626 B.n106 163.367
R745 B.n622 B.n620 163.367
R746 B.n618 B.n108 163.367
R747 B.n614 B.n612 163.367
R748 B.n610 B.n110 163.367
R749 B.n606 B.n604 163.367
R750 B.n602 B.n112 163.367
R751 B.n598 B.n596 163.367
R752 B.n594 B.n114 163.367
R753 B.n590 B.n588 163.367
R754 B.n586 B.n116 163.367
R755 B.n582 B.n580 163.367
R756 B.n578 B.n118 163.367
R757 B.n574 B.n572 163.367
R758 B.n388 B.n198 163.367
R759 B.n392 B.n198 163.367
R760 B.n392 B.n192 163.367
R761 B.n400 B.n192 163.367
R762 B.n400 B.n190 163.367
R763 B.n404 B.n190 163.367
R764 B.n404 B.n184 163.367
R765 B.n412 B.n184 163.367
R766 B.n412 B.n182 163.367
R767 B.n416 B.n182 163.367
R768 B.n416 B.n176 163.367
R769 B.n424 B.n176 163.367
R770 B.n424 B.n174 163.367
R771 B.n428 B.n174 163.367
R772 B.n428 B.n169 163.367
R773 B.n437 B.n169 163.367
R774 B.n437 B.n167 163.367
R775 B.n441 B.n167 163.367
R776 B.n441 B.n161 163.367
R777 B.n449 B.n161 163.367
R778 B.n449 B.n159 163.367
R779 B.n453 B.n159 163.367
R780 B.n453 B.n153 163.367
R781 B.n461 B.n153 163.367
R782 B.n461 B.n151 163.367
R783 B.n465 B.n151 163.367
R784 B.n465 B.n145 163.367
R785 B.n473 B.n145 163.367
R786 B.n473 B.n143 163.367
R787 B.n477 B.n143 163.367
R788 B.n477 B.n137 163.367
R789 B.n485 B.n137 163.367
R790 B.n485 B.n135 163.367
R791 B.n489 B.n135 163.367
R792 B.n489 B.n129 163.367
R793 B.n497 B.n129 163.367
R794 B.n497 B.n127 163.367
R795 B.n502 B.n127 163.367
R796 B.n502 B.n121 163.367
R797 B.n510 B.n121 163.367
R798 B.n511 B.n510 163.367
R799 B.n511 B.n5 163.367
R800 B.n6 B.n5 163.367
R801 B.n7 B.n6 163.367
R802 B.n517 B.n7 163.367
R803 B.n519 B.n517 163.367
R804 B.n519 B.n12 163.367
R805 B.n13 B.n12 163.367
R806 B.n14 B.n13 163.367
R807 B.n524 B.n14 163.367
R808 B.n524 B.n19 163.367
R809 B.n20 B.n19 163.367
R810 B.n21 B.n20 163.367
R811 B.n529 B.n21 163.367
R812 B.n529 B.n26 163.367
R813 B.n27 B.n26 163.367
R814 B.n28 B.n27 163.367
R815 B.n534 B.n28 163.367
R816 B.n534 B.n33 163.367
R817 B.n34 B.n33 163.367
R818 B.n35 B.n34 163.367
R819 B.n539 B.n35 163.367
R820 B.n539 B.n40 163.367
R821 B.n41 B.n40 163.367
R822 B.n42 B.n41 163.367
R823 B.n544 B.n42 163.367
R824 B.n544 B.n47 163.367
R825 B.n48 B.n47 163.367
R826 B.n49 B.n48 163.367
R827 B.n549 B.n49 163.367
R828 B.n549 B.n54 163.367
R829 B.n55 B.n54 163.367
R830 B.n56 B.n55 163.367
R831 B.n554 B.n56 163.367
R832 B.n554 B.n61 163.367
R833 B.n62 B.n61 163.367
R834 B.n63 B.n62 163.367
R835 B.n559 B.n63 163.367
R836 B.n559 B.n68 163.367
R837 B.n69 B.n68 163.367
R838 B.n70 B.n69 163.367
R839 B.n564 B.n70 163.367
R840 B.n564 B.n75 163.367
R841 B.n76 B.n75 163.367
R842 B.n77 B.n76 163.367
R843 B.n382 B.n380 163.367
R844 B.n380 B.n379 163.367
R845 B.n376 B.n375 163.367
R846 B.n373 B.n206 163.367
R847 B.n369 B.n367 163.367
R848 B.n365 B.n208 163.367
R849 B.n361 B.n359 163.367
R850 B.n357 B.n210 163.367
R851 B.n353 B.n351 163.367
R852 B.n349 B.n212 163.367
R853 B.n345 B.n343 163.367
R854 B.n341 B.n214 163.367
R855 B.n337 B.n335 163.367
R856 B.n333 B.n216 163.367
R857 B.n329 B.n327 163.367
R858 B.n325 B.n218 163.367
R859 B.n320 B.n318 163.367
R860 B.n316 B.n222 163.367
R861 B.n312 B.n310 163.367
R862 B.n308 B.n224 163.367
R863 B.n304 B.n302 163.367
R864 B.n299 B.n298 163.367
R865 B.n296 B.n230 163.367
R866 B.n292 B.n290 163.367
R867 B.n288 B.n232 163.367
R868 B.n284 B.n282 163.367
R869 B.n280 B.n234 163.367
R870 B.n276 B.n274 163.367
R871 B.n272 B.n236 163.367
R872 B.n268 B.n266 163.367
R873 B.n264 B.n238 163.367
R874 B.n260 B.n258 163.367
R875 B.n256 B.n240 163.367
R876 B.n252 B.n250 163.367
R877 B.n248 B.n242 163.367
R878 B.n244 B.n200 163.367
R879 B.n386 B.n196 163.367
R880 B.n394 B.n196 163.367
R881 B.n394 B.n194 163.367
R882 B.n398 B.n194 163.367
R883 B.n398 B.n188 163.367
R884 B.n406 B.n188 163.367
R885 B.n406 B.n186 163.367
R886 B.n410 B.n186 163.367
R887 B.n410 B.n180 163.367
R888 B.n418 B.n180 163.367
R889 B.n418 B.n178 163.367
R890 B.n422 B.n178 163.367
R891 B.n422 B.n172 163.367
R892 B.n431 B.n172 163.367
R893 B.n431 B.n170 163.367
R894 B.n435 B.n170 163.367
R895 B.n435 B.n165 163.367
R896 B.n443 B.n165 163.367
R897 B.n443 B.n163 163.367
R898 B.n447 B.n163 163.367
R899 B.n447 B.n157 163.367
R900 B.n455 B.n157 163.367
R901 B.n455 B.n155 163.367
R902 B.n459 B.n155 163.367
R903 B.n459 B.n149 163.367
R904 B.n467 B.n149 163.367
R905 B.n467 B.n147 163.367
R906 B.n471 B.n147 163.367
R907 B.n471 B.n141 163.367
R908 B.n479 B.n141 163.367
R909 B.n479 B.n139 163.367
R910 B.n483 B.n139 163.367
R911 B.n483 B.n133 163.367
R912 B.n491 B.n133 163.367
R913 B.n491 B.n131 163.367
R914 B.n495 B.n131 163.367
R915 B.n495 B.n125 163.367
R916 B.n504 B.n125 163.367
R917 B.n504 B.n123 163.367
R918 B.n508 B.n123 163.367
R919 B.n508 B.n3 163.367
R920 B.n800 B.n3 163.367
R921 B.n796 B.n2 163.367
R922 B.n796 B.n795 163.367
R923 B.n795 B.n9 163.367
R924 B.n791 B.n9 163.367
R925 B.n791 B.n11 163.367
R926 B.n787 B.n11 163.367
R927 B.n787 B.n16 163.367
R928 B.n783 B.n16 163.367
R929 B.n783 B.n18 163.367
R930 B.n779 B.n18 163.367
R931 B.n779 B.n23 163.367
R932 B.n775 B.n23 163.367
R933 B.n775 B.n25 163.367
R934 B.n771 B.n25 163.367
R935 B.n771 B.n30 163.367
R936 B.n767 B.n30 163.367
R937 B.n767 B.n32 163.367
R938 B.n763 B.n32 163.367
R939 B.n763 B.n37 163.367
R940 B.n759 B.n37 163.367
R941 B.n759 B.n39 163.367
R942 B.n755 B.n39 163.367
R943 B.n755 B.n44 163.367
R944 B.n751 B.n44 163.367
R945 B.n751 B.n46 163.367
R946 B.n747 B.n46 163.367
R947 B.n747 B.n50 163.367
R948 B.n743 B.n50 163.367
R949 B.n743 B.n52 163.367
R950 B.n739 B.n52 163.367
R951 B.n739 B.n58 163.367
R952 B.n735 B.n58 163.367
R953 B.n735 B.n60 163.367
R954 B.n731 B.n60 163.367
R955 B.n731 B.n65 163.367
R956 B.n727 B.n65 163.367
R957 B.n727 B.n67 163.367
R958 B.n723 B.n67 163.367
R959 B.n723 B.n72 163.367
R960 B.n719 B.n72 163.367
R961 B.n719 B.n74 163.367
R962 B.n715 B.n74 163.367
R963 B.n103 B.t12 111.921
R964 B.n225 B.t17 111.921
R965 B.n96 B.t19 111.91
R966 B.n219 B.t23 111.91
R967 B.n387 B.n201 100.183
R968 B.n716 B.n78 100.183
R969 B.n104 B.t13 74.1023
R970 B.n226 B.t16 74.1023
R971 B.n97 B.t20 74.0926
R972 B.n220 B.t22 74.0926
R973 B.n710 B.n79 71.676
R974 B.n709 B.n708 71.676
R975 B.n702 B.n81 71.676
R976 B.n701 B.n700 71.676
R977 B.n694 B.n83 71.676
R978 B.n693 B.n692 71.676
R979 B.n686 B.n85 71.676
R980 B.n685 B.n684 71.676
R981 B.n678 B.n87 71.676
R982 B.n677 B.n676 71.676
R983 B.n670 B.n89 71.676
R984 B.n669 B.n668 71.676
R985 B.n662 B.n91 71.676
R986 B.n661 B.n660 71.676
R987 B.n654 B.n93 71.676
R988 B.n653 B.n652 71.676
R989 B.n646 B.n95 71.676
R990 B.n645 B.n644 71.676
R991 B.n638 B.n100 71.676
R992 B.n637 B.n636 71.676
R993 B.n629 B.n102 71.676
R994 B.n628 B.n627 71.676
R995 B.n621 B.n106 71.676
R996 B.n620 B.n619 71.676
R997 B.n613 B.n108 71.676
R998 B.n612 B.n611 71.676
R999 B.n605 B.n110 71.676
R1000 B.n604 B.n603 71.676
R1001 B.n597 B.n112 71.676
R1002 B.n596 B.n595 71.676
R1003 B.n589 B.n114 71.676
R1004 B.n588 B.n587 71.676
R1005 B.n581 B.n116 71.676
R1006 B.n580 B.n579 71.676
R1007 B.n573 B.n118 71.676
R1008 B.n572 B.n571 71.676
R1009 B.n571 B.n570 71.676
R1010 B.n574 B.n573 71.676
R1011 B.n579 B.n578 71.676
R1012 B.n582 B.n581 71.676
R1013 B.n587 B.n586 71.676
R1014 B.n590 B.n589 71.676
R1015 B.n595 B.n594 71.676
R1016 B.n598 B.n597 71.676
R1017 B.n603 B.n602 71.676
R1018 B.n606 B.n605 71.676
R1019 B.n611 B.n610 71.676
R1020 B.n614 B.n613 71.676
R1021 B.n619 B.n618 71.676
R1022 B.n622 B.n621 71.676
R1023 B.n627 B.n626 71.676
R1024 B.n630 B.n629 71.676
R1025 B.n636 B.n635 71.676
R1026 B.n639 B.n638 71.676
R1027 B.n644 B.n643 71.676
R1028 B.n647 B.n646 71.676
R1029 B.n652 B.n651 71.676
R1030 B.n655 B.n654 71.676
R1031 B.n660 B.n659 71.676
R1032 B.n663 B.n662 71.676
R1033 B.n668 B.n667 71.676
R1034 B.n671 B.n670 71.676
R1035 B.n676 B.n675 71.676
R1036 B.n679 B.n678 71.676
R1037 B.n684 B.n683 71.676
R1038 B.n687 B.n686 71.676
R1039 B.n692 B.n691 71.676
R1040 B.n695 B.n694 71.676
R1041 B.n700 B.n699 71.676
R1042 B.n703 B.n702 71.676
R1043 B.n708 B.n707 71.676
R1044 B.n711 B.n710 71.676
R1045 B.n381 B.n202 71.676
R1046 B.n379 B.n204 71.676
R1047 B.n375 B.n374 71.676
R1048 B.n368 B.n206 71.676
R1049 B.n367 B.n366 71.676
R1050 B.n360 B.n208 71.676
R1051 B.n359 B.n358 71.676
R1052 B.n352 B.n210 71.676
R1053 B.n351 B.n350 71.676
R1054 B.n344 B.n212 71.676
R1055 B.n343 B.n342 71.676
R1056 B.n336 B.n214 71.676
R1057 B.n335 B.n334 71.676
R1058 B.n328 B.n216 71.676
R1059 B.n327 B.n326 71.676
R1060 B.n319 B.n218 71.676
R1061 B.n318 B.n317 71.676
R1062 B.n311 B.n222 71.676
R1063 B.n310 B.n309 71.676
R1064 B.n303 B.n224 71.676
R1065 B.n302 B.n228 71.676
R1066 B.n298 B.n297 71.676
R1067 B.n291 B.n230 71.676
R1068 B.n290 B.n289 71.676
R1069 B.n283 B.n232 71.676
R1070 B.n282 B.n281 71.676
R1071 B.n275 B.n234 71.676
R1072 B.n274 B.n273 71.676
R1073 B.n267 B.n236 71.676
R1074 B.n266 B.n265 71.676
R1075 B.n259 B.n238 71.676
R1076 B.n258 B.n257 71.676
R1077 B.n251 B.n240 71.676
R1078 B.n250 B.n249 71.676
R1079 B.n243 B.n242 71.676
R1080 B.n382 B.n381 71.676
R1081 B.n376 B.n204 71.676
R1082 B.n374 B.n373 71.676
R1083 B.n369 B.n368 71.676
R1084 B.n366 B.n365 71.676
R1085 B.n361 B.n360 71.676
R1086 B.n358 B.n357 71.676
R1087 B.n353 B.n352 71.676
R1088 B.n350 B.n349 71.676
R1089 B.n345 B.n344 71.676
R1090 B.n342 B.n341 71.676
R1091 B.n337 B.n336 71.676
R1092 B.n334 B.n333 71.676
R1093 B.n329 B.n328 71.676
R1094 B.n326 B.n325 71.676
R1095 B.n320 B.n319 71.676
R1096 B.n317 B.n316 71.676
R1097 B.n312 B.n311 71.676
R1098 B.n309 B.n308 71.676
R1099 B.n304 B.n303 71.676
R1100 B.n299 B.n228 71.676
R1101 B.n297 B.n296 71.676
R1102 B.n292 B.n291 71.676
R1103 B.n289 B.n288 71.676
R1104 B.n284 B.n283 71.676
R1105 B.n281 B.n280 71.676
R1106 B.n276 B.n275 71.676
R1107 B.n273 B.n272 71.676
R1108 B.n268 B.n267 71.676
R1109 B.n265 B.n264 71.676
R1110 B.n260 B.n259 71.676
R1111 B.n257 B.n256 71.676
R1112 B.n252 B.n251 71.676
R1113 B.n249 B.n248 71.676
R1114 B.n244 B.n243 71.676
R1115 B.n801 B.n800 71.676
R1116 B.n801 B.n2 71.676
R1117 B.n98 B.n97 59.5399
R1118 B.n632 B.n104 59.5399
R1119 B.n227 B.n226 59.5399
R1120 B.n323 B.n220 59.5399
R1121 B.n387 B.n197 54.4996
R1122 B.n393 B.n197 54.4996
R1123 B.n393 B.n193 54.4996
R1124 B.n399 B.n193 54.4996
R1125 B.n399 B.n189 54.4996
R1126 B.n405 B.n189 54.4996
R1127 B.n411 B.n185 54.4996
R1128 B.n411 B.n181 54.4996
R1129 B.n417 B.n181 54.4996
R1130 B.n417 B.n177 54.4996
R1131 B.n423 B.n177 54.4996
R1132 B.n423 B.n173 54.4996
R1133 B.n430 B.n173 54.4996
R1134 B.n430 B.n429 54.4996
R1135 B.n436 B.n166 54.4996
R1136 B.n442 B.n166 54.4996
R1137 B.n442 B.n162 54.4996
R1138 B.n448 B.n162 54.4996
R1139 B.n454 B.n158 54.4996
R1140 B.n454 B.n154 54.4996
R1141 B.n460 B.n154 54.4996
R1142 B.n460 B.n150 54.4996
R1143 B.n466 B.n150 54.4996
R1144 B.n472 B.n146 54.4996
R1145 B.n472 B.n142 54.4996
R1146 B.n478 B.n142 54.4996
R1147 B.n478 B.n138 54.4996
R1148 B.n484 B.n138 54.4996
R1149 B.n490 B.n134 54.4996
R1150 B.n490 B.n130 54.4996
R1151 B.n496 B.n130 54.4996
R1152 B.n496 B.n126 54.4996
R1153 B.n503 B.n126 54.4996
R1154 B.n509 B.n122 54.4996
R1155 B.n509 B.n4 54.4996
R1156 B.n799 B.n4 54.4996
R1157 B.n799 B.n798 54.4996
R1158 B.n798 B.n797 54.4996
R1159 B.n797 B.n8 54.4996
R1160 B.n518 B.n8 54.4996
R1161 B.n790 B.n789 54.4996
R1162 B.n789 B.n788 54.4996
R1163 B.n788 B.n15 54.4996
R1164 B.n782 B.n15 54.4996
R1165 B.n782 B.n781 54.4996
R1166 B.n780 B.n22 54.4996
R1167 B.n774 B.n22 54.4996
R1168 B.n774 B.n773 54.4996
R1169 B.n773 B.n772 54.4996
R1170 B.n772 B.n29 54.4996
R1171 B.n766 B.n765 54.4996
R1172 B.n765 B.n764 54.4996
R1173 B.n764 B.n36 54.4996
R1174 B.n758 B.n36 54.4996
R1175 B.n758 B.n757 54.4996
R1176 B.n756 B.n43 54.4996
R1177 B.n750 B.n43 54.4996
R1178 B.n750 B.n749 54.4996
R1179 B.n749 B.n748 54.4996
R1180 B.n742 B.n53 54.4996
R1181 B.n742 B.n741 54.4996
R1182 B.n741 B.n740 54.4996
R1183 B.n740 B.n57 54.4996
R1184 B.n734 B.n57 54.4996
R1185 B.n734 B.n733 54.4996
R1186 B.n733 B.n732 54.4996
R1187 B.n732 B.n64 54.4996
R1188 B.n726 B.n725 54.4996
R1189 B.n725 B.n724 54.4996
R1190 B.n724 B.n71 54.4996
R1191 B.n718 B.n71 54.4996
R1192 B.n718 B.n717 54.4996
R1193 B.n717 B.n716 54.4996
R1194 B.t4 B.n122 52.8967
R1195 B.n518 B.t5 52.8967
R1196 B.n436 B.t8 49.6908
R1197 B.n748 B.t3 49.6908
R1198 B.t15 B.n185 46.485
R1199 B.t11 B.n64 46.485
R1200 B.n448 B.t7 44.8821
R1201 B.t0 B.n756 44.8821
R1202 B.t2 B.n134 38.4704
R1203 B.n781 B.t1 38.4704
R1204 B.n97 B.n96 37.8187
R1205 B.n104 B.n103 37.8187
R1206 B.n226 B.n225 37.8187
R1207 B.n220 B.n219 37.8187
R1208 B.n385 B.n384 32.3127
R1209 B.n389 B.n199 32.3127
R1210 B.n569 B.n568 32.3127
R1211 B.n714 B.n713 32.3127
R1212 B.n466 B.t6 30.4559
R1213 B.n766 B.t9 30.4559
R1214 B.t6 B.n146 24.0442
R1215 B.t9 B.n29 24.0442
R1216 B B.n802 18.0485
R1217 B.n484 B.t2 16.0296
R1218 B.t1 B.n780 16.0296
R1219 B.n385 B.n195 10.6151
R1220 B.n395 B.n195 10.6151
R1221 B.n396 B.n395 10.6151
R1222 B.n397 B.n396 10.6151
R1223 B.n397 B.n187 10.6151
R1224 B.n407 B.n187 10.6151
R1225 B.n408 B.n407 10.6151
R1226 B.n409 B.n408 10.6151
R1227 B.n409 B.n179 10.6151
R1228 B.n419 B.n179 10.6151
R1229 B.n420 B.n419 10.6151
R1230 B.n421 B.n420 10.6151
R1231 B.n421 B.n171 10.6151
R1232 B.n432 B.n171 10.6151
R1233 B.n433 B.n432 10.6151
R1234 B.n434 B.n433 10.6151
R1235 B.n434 B.n164 10.6151
R1236 B.n444 B.n164 10.6151
R1237 B.n445 B.n444 10.6151
R1238 B.n446 B.n445 10.6151
R1239 B.n446 B.n156 10.6151
R1240 B.n456 B.n156 10.6151
R1241 B.n457 B.n456 10.6151
R1242 B.n458 B.n457 10.6151
R1243 B.n458 B.n148 10.6151
R1244 B.n468 B.n148 10.6151
R1245 B.n469 B.n468 10.6151
R1246 B.n470 B.n469 10.6151
R1247 B.n470 B.n140 10.6151
R1248 B.n480 B.n140 10.6151
R1249 B.n481 B.n480 10.6151
R1250 B.n482 B.n481 10.6151
R1251 B.n482 B.n132 10.6151
R1252 B.n492 B.n132 10.6151
R1253 B.n493 B.n492 10.6151
R1254 B.n494 B.n493 10.6151
R1255 B.n494 B.n124 10.6151
R1256 B.n505 B.n124 10.6151
R1257 B.n506 B.n505 10.6151
R1258 B.n507 B.n506 10.6151
R1259 B.n507 B.n0 10.6151
R1260 B.n384 B.n383 10.6151
R1261 B.n383 B.n203 10.6151
R1262 B.n378 B.n203 10.6151
R1263 B.n378 B.n377 10.6151
R1264 B.n377 B.n205 10.6151
R1265 B.n372 B.n205 10.6151
R1266 B.n372 B.n371 10.6151
R1267 B.n371 B.n370 10.6151
R1268 B.n370 B.n207 10.6151
R1269 B.n364 B.n207 10.6151
R1270 B.n364 B.n363 10.6151
R1271 B.n363 B.n362 10.6151
R1272 B.n362 B.n209 10.6151
R1273 B.n356 B.n209 10.6151
R1274 B.n356 B.n355 10.6151
R1275 B.n355 B.n354 10.6151
R1276 B.n354 B.n211 10.6151
R1277 B.n348 B.n211 10.6151
R1278 B.n348 B.n347 10.6151
R1279 B.n347 B.n346 10.6151
R1280 B.n346 B.n213 10.6151
R1281 B.n340 B.n213 10.6151
R1282 B.n340 B.n339 10.6151
R1283 B.n339 B.n338 10.6151
R1284 B.n338 B.n215 10.6151
R1285 B.n332 B.n215 10.6151
R1286 B.n332 B.n331 10.6151
R1287 B.n331 B.n330 10.6151
R1288 B.n330 B.n217 10.6151
R1289 B.n324 B.n217 10.6151
R1290 B.n322 B.n321 10.6151
R1291 B.n321 B.n221 10.6151
R1292 B.n315 B.n221 10.6151
R1293 B.n315 B.n314 10.6151
R1294 B.n314 B.n313 10.6151
R1295 B.n313 B.n223 10.6151
R1296 B.n307 B.n223 10.6151
R1297 B.n307 B.n306 10.6151
R1298 B.n306 B.n305 10.6151
R1299 B.n301 B.n300 10.6151
R1300 B.n300 B.n229 10.6151
R1301 B.n295 B.n229 10.6151
R1302 B.n295 B.n294 10.6151
R1303 B.n294 B.n293 10.6151
R1304 B.n293 B.n231 10.6151
R1305 B.n287 B.n231 10.6151
R1306 B.n287 B.n286 10.6151
R1307 B.n286 B.n285 10.6151
R1308 B.n285 B.n233 10.6151
R1309 B.n279 B.n233 10.6151
R1310 B.n279 B.n278 10.6151
R1311 B.n278 B.n277 10.6151
R1312 B.n277 B.n235 10.6151
R1313 B.n271 B.n235 10.6151
R1314 B.n271 B.n270 10.6151
R1315 B.n270 B.n269 10.6151
R1316 B.n269 B.n237 10.6151
R1317 B.n263 B.n237 10.6151
R1318 B.n263 B.n262 10.6151
R1319 B.n262 B.n261 10.6151
R1320 B.n261 B.n239 10.6151
R1321 B.n255 B.n239 10.6151
R1322 B.n255 B.n254 10.6151
R1323 B.n254 B.n253 10.6151
R1324 B.n253 B.n241 10.6151
R1325 B.n247 B.n241 10.6151
R1326 B.n247 B.n246 10.6151
R1327 B.n246 B.n245 10.6151
R1328 B.n245 B.n199 10.6151
R1329 B.n390 B.n389 10.6151
R1330 B.n391 B.n390 10.6151
R1331 B.n391 B.n191 10.6151
R1332 B.n401 B.n191 10.6151
R1333 B.n402 B.n401 10.6151
R1334 B.n403 B.n402 10.6151
R1335 B.n403 B.n183 10.6151
R1336 B.n413 B.n183 10.6151
R1337 B.n414 B.n413 10.6151
R1338 B.n415 B.n414 10.6151
R1339 B.n415 B.n175 10.6151
R1340 B.n425 B.n175 10.6151
R1341 B.n426 B.n425 10.6151
R1342 B.n427 B.n426 10.6151
R1343 B.n427 B.n168 10.6151
R1344 B.n438 B.n168 10.6151
R1345 B.n439 B.n438 10.6151
R1346 B.n440 B.n439 10.6151
R1347 B.n440 B.n160 10.6151
R1348 B.n450 B.n160 10.6151
R1349 B.n451 B.n450 10.6151
R1350 B.n452 B.n451 10.6151
R1351 B.n452 B.n152 10.6151
R1352 B.n462 B.n152 10.6151
R1353 B.n463 B.n462 10.6151
R1354 B.n464 B.n463 10.6151
R1355 B.n464 B.n144 10.6151
R1356 B.n474 B.n144 10.6151
R1357 B.n475 B.n474 10.6151
R1358 B.n476 B.n475 10.6151
R1359 B.n476 B.n136 10.6151
R1360 B.n486 B.n136 10.6151
R1361 B.n487 B.n486 10.6151
R1362 B.n488 B.n487 10.6151
R1363 B.n488 B.n128 10.6151
R1364 B.n498 B.n128 10.6151
R1365 B.n499 B.n498 10.6151
R1366 B.n501 B.n499 10.6151
R1367 B.n501 B.n500 10.6151
R1368 B.n500 B.n120 10.6151
R1369 B.n512 B.n120 10.6151
R1370 B.n513 B.n512 10.6151
R1371 B.n514 B.n513 10.6151
R1372 B.n515 B.n514 10.6151
R1373 B.n516 B.n515 10.6151
R1374 B.n520 B.n516 10.6151
R1375 B.n521 B.n520 10.6151
R1376 B.n522 B.n521 10.6151
R1377 B.n523 B.n522 10.6151
R1378 B.n525 B.n523 10.6151
R1379 B.n526 B.n525 10.6151
R1380 B.n527 B.n526 10.6151
R1381 B.n528 B.n527 10.6151
R1382 B.n530 B.n528 10.6151
R1383 B.n531 B.n530 10.6151
R1384 B.n532 B.n531 10.6151
R1385 B.n533 B.n532 10.6151
R1386 B.n535 B.n533 10.6151
R1387 B.n536 B.n535 10.6151
R1388 B.n537 B.n536 10.6151
R1389 B.n538 B.n537 10.6151
R1390 B.n540 B.n538 10.6151
R1391 B.n541 B.n540 10.6151
R1392 B.n542 B.n541 10.6151
R1393 B.n543 B.n542 10.6151
R1394 B.n545 B.n543 10.6151
R1395 B.n546 B.n545 10.6151
R1396 B.n547 B.n546 10.6151
R1397 B.n548 B.n547 10.6151
R1398 B.n550 B.n548 10.6151
R1399 B.n551 B.n550 10.6151
R1400 B.n552 B.n551 10.6151
R1401 B.n553 B.n552 10.6151
R1402 B.n555 B.n553 10.6151
R1403 B.n556 B.n555 10.6151
R1404 B.n557 B.n556 10.6151
R1405 B.n558 B.n557 10.6151
R1406 B.n560 B.n558 10.6151
R1407 B.n561 B.n560 10.6151
R1408 B.n562 B.n561 10.6151
R1409 B.n563 B.n562 10.6151
R1410 B.n565 B.n563 10.6151
R1411 B.n566 B.n565 10.6151
R1412 B.n567 B.n566 10.6151
R1413 B.n568 B.n567 10.6151
R1414 B.n794 B.n1 10.6151
R1415 B.n794 B.n793 10.6151
R1416 B.n793 B.n792 10.6151
R1417 B.n792 B.n10 10.6151
R1418 B.n786 B.n10 10.6151
R1419 B.n786 B.n785 10.6151
R1420 B.n785 B.n784 10.6151
R1421 B.n784 B.n17 10.6151
R1422 B.n778 B.n17 10.6151
R1423 B.n778 B.n777 10.6151
R1424 B.n777 B.n776 10.6151
R1425 B.n776 B.n24 10.6151
R1426 B.n770 B.n24 10.6151
R1427 B.n770 B.n769 10.6151
R1428 B.n769 B.n768 10.6151
R1429 B.n768 B.n31 10.6151
R1430 B.n762 B.n31 10.6151
R1431 B.n762 B.n761 10.6151
R1432 B.n761 B.n760 10.6151
R1433 B.n760 B.n38 10.6151
R1434 B.n754 B.n38 10.6151
R1435 B.n754 B.n753 10.6151
R1436 B.n753 B.n752 10.6151
R1437 B.n752 B.n45 10.6151
R1438 B.n746 B.n45 10.6151
R1439 B.n746 B.n745 10.6151
R1440 B.n745 B.n744 10.6151
R1441 B.n744 B.n51 10.6151
R1442 B.n738 B.n51 10.6151
R1443 B.n738 B.n737 10.6151
R1444 B.n737 B.n736 10.6151
R1445 B.n736 B.n59 10.6151
R1446 B.n730 B.n59 10.6151
R1447 B.n730 B.n729 10.6151
R1448 B.n729 B.n728 10.6151
R1449 B.n728 B.n66 10.6151
R1450 B.n722 B.n66 10.6151
R1451 B.n722 B.n721 10.6151
R1452 B.n721 B.n720 10.6151
R1453 B.n720 B.n73 10.6151
R1454 B.n714 B.n73 10.6151
R1455 B.n713 B.n712 10.6151
R1456 B.n712 B.n80 10.6151
R1457 B.n706 B.n80 10.6151
R1458 B.n706 B.n705 10.6151
R1459 B.n705 B.n704 10.6151
R1460 B.n704 B.n82 10.6151
R1461 B.n698 B.n82 10.6151
R1462 B.n698 B.n697 10.6151
R1463 B.n697 B.n696 10.6151
R1464 B.n696 B.n84 10.6151
R1465 B.n690 B.n84 10.6151
R1466 B.n690 B.n689 10.6151
R1467 B.n689 B.n688 10.6151
R1468 B.n688 B.n86 10.6151
R1469 B.n682 B.n86 10.6151
R1470 B.n682 B.n681 10.6151
R1471 B.n681 B.n680 10.6151
R1472 B.n680 B.n88 10.6151
R1473 B.n674 B.n88 10.6151
R1474 B.n674 B.n673 10.6151
R1475 B.n673 B.n672 10.6151
R1476 B.n672 B.n90 10.6151
R1477 B.n666 B.n90 10.6151
R1478 B.n666 B.n665 10.6151
R1479 B.n665 B.n664 10.6151
R1480 B.n664 B.n92 10.6151
R1481 B.n658 B.n92 10.6151
R1482 B.n658 B.n657 10.6151
R1483 B.n657 B.n656 10.6151
R1484 B.n656 B.n94 10.6151
R1485 B.n650 B.n649 10.6151
R1486 B.n649 B.n648 10.6151
R1487 B.n648 B.n99 10.6151
R1488 B.n642 B.n99 10.6151
R1489 B.n642 B.n641 10.6151
R1490 B.n641 B.n640 10.6151
R1491 B.n640 B.n101 10.6151
R1492 B.n634 B.n101 10.6151
R1493 B.n634 B.n633 10.6151
R1494 B.n631 B.n105 10.6151
R1495 B.n625 B.n105 10.6151
R1496 B.n625 B.n624 10.6151
R1497 B.n624 B.n623 10.6151
R1498 B.n623 B.n107 10.6151
R1499 B.n617 B.n107 10.6151
R1500 B.n617 B.n616 10.6151
R1501 B.n616 B.n615 10.6151
R1502 B.n615 B.n109 10.6151
R1503 B.n609 B.n109 10.6151
R1504 B.n609 B.n608 10.6151
R1505 B.n608 B.n607 10.6151
R1506 B.n607 B.n111 10.6151
R1507 B.n601 B.n111 10.6151
R1508 B.n601 B.n600 10.6151
R1509 B.n600 B.n599 10.6151
R1510 B.n599 B.n113 10.6151
R1511 B.n593 B.n113 10.6151
R1512 B.n593 B.n592 10.6151
R1513 B.n592 B.n591 10.6151
R1514 B.n591 B.n115 10.6151
R1515 B.n585 B.n115 10.6151
R1516 B.n585 B.n584 10.6151
R1517 B.n584 B.n583 10.6151
R1518 B.n583 B.n117 10.6151
R1519 B.n577 B.n117 10.6151
R1520 B.n577 B.n576 10.6151
R1521 B.n576 B.n575 10.6151
R1522 B.n575 B.n119 10.6151
R1523 B.n569 B.n119 10.6151
R1524 B.t7 B.n158 9.61799
R1525 B.n757 B.t0 9.61799
R1526 B.n324 B.n323 9.36635
R1527 B.n301 B.n227 9.36635
R1528 B.n98 B.n94 9.36635
R1529 B.n632 B.n631 9.36635
R1530 B.n802 B.n0 8.11757
R1531 B.n802 B.n1 8.11757
R1532 B.n405 B.t15 8.01507
R1533 B.n726 B.t11 8.01507
R1534 B.n429 B.t8 4.80924
R1535 B.n53 B.t3 4.80924
R1536 B.n503 B.t4 1.60341
R1537 B.n790 B.t5 1.60341
R1538 B.n323 B.n322 1.24928
R1539 B.n305 B.n227 1.24928
R1540 B.n650 B.n98 1.24928
R1541 B.n633 B.n632 1.24928
R1542 VP.n39 VP.n38 178.428
R1543 VP.n68 VP.n67 178.428
R1544 VP.n37 VP.n36 178.428
R1545 VP.n17 VP.n16 161.3
R1546 VP.n18 VP.n13 161.3
R1547 VP.n20 VP.n19 161.3
R1548 VP.n21 VP.n12 161.3
R1549 VP.n24 VP.n23 161.3
R1550 VP.n25 VP.n11 161.3
R1551 VP.n27 VP.n26 161.3
R1552 VP.n28 VP.n10 161.3
R1553 VP.n31 VP.n30 161.3
R1554 VP.n32 VP.n9 161.3
R1555 VP.n34 VP.n33 161.3
R1556 VP.n35 VP.n8 161.3
R1557 VP.n66 VP.n0 161.3
R1558 VP.n65 VP.n64 161.3
R1559 VP.n63 VP.n1 161.3
R1560 VP.n62 VP.n61 161.3
R1561 VP.n59 VP.n2 161.3
R1562 VP.n58 VP.n57 161.3
R1563 VP.n56 VP.n3 161.3
R1564 VP.n55 VP.n54 161.3
R1565 VP.n52 VP.n4 161.3
R1566 VP.n51 VP.n50 161.3
R1567 VP.n49 VP.n5 161.3
R1568 VP.n48 VP.n47 161.3
R1569 VP.n45 VP.n6 161.3
R1570 VP.n44 VP.n43 161.3
R1571 VP.n42 VP.n7 161.3
R1572 VP.n41 VP.n40 161.3
R1573 VP.n14 VP.t6 158.025
R1574 VP.n39 VP.t3 125.707
R1575 VP.n46 VP.t5 125.707
R1576 VP.n53 VP.t0 125.707
R1577 VP.n60 VP.t1 125.707
R1578 VP.n67 VP.t2 125.707
R1579 VP.n36 VP.t4 125.707
R1580 VP.n29 VP.t9 125.707
R1581 VP.n22 VP.t7 125.707
R1582 VP.n15 VP.t8 125.707
R1583 VP.n44 VP.n7 56.5193
R1584 VP.n51 VP.n5 56.5193
R1585 VP.n58 VP.n3 56.5193
R1586 VP.n65 VP.n1 56.5193
R1587 VP.n34 VP.n9 56.5193
R1588 VP.n27 VP.n11 56.5193
R1589 VP.n20 VP.n13 56.5193
R1590 VP.n15 VP.n14 56.3226
R1591 VP.n38 VP.n37 45.0119
R1592 VP.n40 VP.n7 24.4675
R1593 VP.n45 VP.n44 24.4675
R1594 VP.n47 VP.n5 24.4675
R1595 VP.n52 VP.n51 24.4675
R1596 VP.n54 VP.n3 24.4675
R1597 VP.n59 VP.n58 24.4675
R1598 VP.n61 VP.n1 24.4675
R1599 VP.n66 VP.n65 24.4675
R1600 VP.n35 VP.n34 24.4675
R1601 VP.n28 VP.n27 24.4675
R1602 VP.n30 VP.n9 24.4675
R1603 VP.n21 VP.n20 24.4675
R1604 VP.n23 VP.n11 24.4675
R1605 VP.n16 VP.n13 24.4675
R1606 VP.n17 VP.n14 18.0474
R1607 VP.n46 VP.n45 14.6807
R1608 VP.n61 VP.n60 14.6807
R1609 VP.n30 VP.n29 14.6807
R1610 VP.n53 VP.n52 12.234
R1611 VP.n54 VP.n53 12.234
R1612 VP.n22 VP.n21 12.234
R1613 VP.n23 VP.n22 12.234
R1614 VP.n47 VP.n46 9.7873
R1615 VP.n60 VP.n59 9.7873
R1616 VP.n29 VP.n28 9.7873
R1617 VP.n16 VP.n15 9.7873
R1618 VP.n40 VP.n39 7.3406
R1619 VP.n67 VP.n66 7.3406
R1620 VP.n36 VP.n35 7.3406
R1621 VP.n18 VP.n17 0.189894
R1622 VP.n19 VP.n18 0.189894
R1623 VP.n19 VP.n12 0.189894
R1624 VP.n24 VP.n12 0.189894
R1625 VP.n25 VP.n24 0.189894
R1626 VP.n26 VP.n25 0.189894
R1627 VP.n26 VP.n10 0.189894
R1628 VP.n31 VP.n10 0.189894
R1629 VP.n32 VP.n31 0.189894
R1630 VP.n33 VP.n32 0.189894
R1631 VP.n33 VP.n8 0.189894
R1632 VP.n37 VP.n8 0.189894
R1633 VP.n41 VP.n38 0.189894
R1634 VP.n42 VP.n41 0.189894
R1635 VP.n43 VP.n42 0.189894
R1636 VP.n43 VP.n6 0.189894
R1637 VP.n48 VP.n6 0.189894
R1638 VP.n49 VP.n48 0.189894
R1639 VP.n50 VP.n49 0.189894
R1640 VP.n50 VP.n4 0.189894
R1641 VP.n55 VP.n4 0.189894
R1642 VP.n56 VP.n55 0.189894
R1643 VP.n57 VP.n56 0.189894
R1644 VP.n57 VP.n2 0.189894
R1645 VP.n62 VP.n2 0.189894
R1646 VP.n63 VP.n62 0.189894
R1647 VP.n64 VP.n63 0.189894
R1648 VP.n64 VP.n0 0.189894
R1649 VP.n68 VP.n0 0.189894
R1650 VP VP.n68 0.0516364
R1651 VDD1.n1 VDD1.t3 66.8727
R1652 VDD1.n3 VDD1.t6 66.8725
R1653 VDD1.n5 VDD1.n4 64.0539
R1654 VDD1.n7 VDD1.n6 62.8485
R1655 VDD1.n1 VDD1.n0 62.8485
R1656 VDD1.n3 VDD1.n2 62.8485
R1657 VDD1.n7 VDD1.n5 40.4082
R1658 VDD1.n6 VDD1.t0 2.3437
R1659 VDD1.n6 VDD1.t5 2.3437
R1660 VDD1.n0 VDD1.t1 2.3437
R1661 VDD1.n0 VDD1.t2 2.3437
R1662 VDD1.n4 VDD1.t8 2.3437
R1663 VDD1.n4 VDD1.t7 2.3437
R1664 VDD1.n2 VDD1.t4 2.3437
R1665 VDD1.n2 VDD1.t9 2.3437
R1666 VDD1 VDD1.n7 1.20309
R1667 VDD1 VDD1.n1 0.478948
R1668 VDD1.n5 VDD1.n3 0.365413
C0 VN VTAIL 7.19139f
C1 VP VDD1 7.11794f
C2 VTAIL VDD2 8.69339f
C3 VN VDD2 6.81396f
C4 VTAIL VP 7.2057f
C5 VN VP 6.29593f
C6 VP VDD2 0.458411f
C7 VTAIL VDD1 8.64921f
C8 VN VDD1 0.151262f
C9 VDD2 VDD1 1.53752f
C10 VDD2 B 5.434114f
C11 VDD1 B 5.402916f
C12 VTAIL B 6.045504f
C13 VN B 13.2139f
C14 VP B 11.686296f
C15 VDD1.t3 B 1.67615f
C16 VDD1.t1 B 0.151612f
C17 VDD1.t2 B 0.151612f
C18 VDD1.n0 B 1.30961f
C19 VDD1.n1 B 0.718631f
C20 VDD1.t6 B 1.67614f
C21 VDD1.t4 B 0.151612f
C22 VDD1.t9 B 0.151612f
C23 VDD1.n2 B 1.30961f
C24 VDD1.n3 B 0.711774f
C25 VDD1.t8 B 0.151612f
C26 VDD1.t7 B 0.151612f
C27 VDD1.n4 B 1.31735f
C28 VDD1.n5 B 2.06824f
C29 VDD1.t0 B 0.151612f
C30 VDD1.t5 B 0.151612f
C31 VDD1.n6 B 1.30961f
C32 VDD1.n7 B 2.267f
C33 VP.n0 B 0.029949f
C34 VP.t2 B 1.10362f
C35 VP.n1 B 0.037464f
C36 VP.n2 B 0.029949f
C37 VP.t1 B 1.10362f
C38 VP.n3 B 0.041637f
C39 VP.n4 B 0.029949f
C40 VP.t0 B 1.10362f
C41 VP.n5 B 0.04581f
C42 VP.n6 B 0.029949f
C43 VP.t5 B 1.10362f
C44 VP.n7 B 0.049982f
C45 VP.n8 B 0.029949f
C46 VP.t4 B 1.10362f
C47 VP.n9 B 0.037464f
C48 VP.n10 B 0.029949f
C49 VP.t9 B 1.10362f
C50 VP.n11 B 0.041637f
C51 VP.n12 B 0.029949f
C52 VP.t7 B 1.10362f
C53 VP.n13 B 0.04581f
C54 VP.t6 B 1.21277f
C55 VP.n14 B 0.481016f
C56 VP.t8 B 1.10362f
C57 VP.n15 B 0.466812f
C58 VP.n16 B 0.039283f
C59 VP.n17 B 0.191018f
C60 VP.n18 B 0.029949f
C61 VP.n19 B 0.029949f
C62 VP.n20 B 0.041637f
C63 VP.n21 B 0.042039f
C64 VP.n22 B 0.410538f
C65 VP.n23 B 0.042039f
C66 VP.n24 B 0.029949f
C67 VP.n25 B 0.029949f
C68 VP.n26 B 0.029949f
C69 VP.n27 B 0.04581f
C70 VP.n28 B 0.039283f
C71 VP.n29 B 0.410538f
C72 VP.n30 B 0.044795f
C73 VP.n31 B 0.029949f
C74 VP.n32 B 0.029949f
C75 VP.n33 B 0.029949f
C76 VP.n34 B 0.049982f
C77 VP.n35 B 0.036528f
C78 VP.n36 B 0.474451f
C79 VP.n37 B 1.39068f
C80 VP.n38 B 1.41459f
C81 VP.t3 B 1.10362f
C82 VP.n39 B 0.474451f
C83 VP.n40 B 0.036528f
C84 VP.n41 B 0.029949f
C85 VP.n42 B 0.029949f
C86 VP.n43 B 0.029949f
C87 VP.n44 B 0.037464f
C88 VP.n45 B 0.044795f
C89 VP.n46 B 0.410538f
C90 VP.n47 B 0.039283f
C91 VP.n48 B 0.029949f
C92 VP.n49 B 0.029949f
C93 VP.n50 B 0.029949f
C94 VP.n51 B 0.041637f
C95 VP.n52 B 0.042039f
C96 VP.n53 B 0.410538f
C97 VP.n54 B 0.042039f
C98 VP.n55 B 0.029949f
C99 VP.n56 B 0.029949f
C100 VP.n57 B 0.029949f
C101 VP.n58 B 0.04581f
C102 VP.n59 B 0.039283f
C103 VP.n60 B 0.410538f
C104 VP.n61 B 0.044795f
C105 VP.n62 B 0.029949f
C106 VP.n63 B 0.029949f
C107 VP.n64 B 0.029949f
C108 VP.n65 B 0.049982f
C109 VP.n66 B 0.036528f
C110 VP.n67 B 0.474451f
C111 VP.n68 B 0.029996f
C112 VDD2.t4 B 1.66368f
C113 VDD2.t6 B 0.150485f
C114 VDD2.t7 B 0.150485f
C115 VDD2.n0 B 1.29987f
C116 VDD2.n1 B 0.70648f
C117 VDD2.t8 B 0.150485f
C118 VDD2.t9 B 0.150485f
C119 VDD2.n2 B 1.30755f
C120 VDD2.n3 B 1.96511f
C121 VDD2.t0 B 1.65422f
C122 VDD2.n4 B 2.22339f
C123 VDD2.t1 B 0.150485f
C124 VDD2.t2 B 0.150485f
C125 VDD2.n5 B 1.29987f
C126 VDD2.n6 B 0.346177f
C127 VDD2.t3 B 0.150485f
C128 VDD2.t5 B 0.150485f
C129 VDD2.n7 B 1.30753f
C130 VTAIL.t13 B 0.170619f
C131 VTAIL.t18 B 0.170619f
C132 VTAIL.n0 B 1.39798f
C133 VTAIL.n1 B 0.472253f
C134 VTAIL.t4 B 1.78154f
C135 VTAIL.n2 B 0.583826f
C136 VTAIL.t6 B 0.170619f
C137 VTAIL.t2 B 0.170619f
C138 VTAIL.n3 B 1.39798f
C139 VTAIL.n4 B 0.532583f
C140 VTAIL.t8 B 0.170619f
C141 VTAIL.t7 B 0.170619f
C142 VTAIL.n5 B 1.39798f
C143 VTAIL.n6 B 1.61783f
C144 VTAIL.t9 B 0.170619f
C145 VTAIL.t12 B 0.170619f
C146 VTAIL.n7 B 1.39798f
C147 VTAIL.n8 B 1.61782f
C148 VTAIL.t14 B 0.170619f
C149 VTAIL.t10 B 0.170619f
C150 VTAIL.n9 B 1.39798f
C151 VTAIL.n10 B 0.53258f
C152 VTAIL.t17 B 1.78155f
C153 VTAIL.n11 B 0.583818f
C154 VTAIL.t5 B 0.170619f
C155 VTAIL.t1 B 0.170619f
C156 VTAIL.n12 B 1.39798f
C157 VTAIL.n13 B 0.50206f
C158 VTAIL.t19 B 0.170619f
C159 VTAIL.t0 B 0.170619f
C160 VTAIL.n14 B 1.39798f
C161 VTAIL.n15 B 0.53258f
C162 VTAIL.t3 B 1.78155f
C163 VTAIL.n16 B 1.56117f
C164 VTAIL.t16 B 1.78154f
C165 VTAIL.n17 B 1.56118f
C166 VTAIL.t15 B 0.170619f
C167 VTAIL.t11 B 0.170619f
C168 VTAIL.n18 B 1.39798f
C169 VTAIL.n19 B 0.423989f
C170 VN.n0 B 0.029453f
C171 VN.t0 B 1.08533f
C172 VN.n1 B 0.036843f
C173 VN.n2 B 0.029453f
C174 VN.t1 B 1.08533f
C175 VN.n3 B 0.040947f
C176 VN.n4 B 0.029453f
C177 VN.t2 B 1.08533f
C178 VN.n5 B 0.04505f
C179 VN.t5 B 1.19267f
C180 VN.n6 B 0.473045f
C181 VN.t3 B 1.08533f
C182 VN.n7 B 0.459075f
C183 VN.n8 B 0.038632f
C184 VN.n9 B 0.187852f
C185 VN.n10 B 0.029453f
C186 VN.n11 B 0.029453f
C187 VN.n12 B 0.040947f
C188 VN.n13 B 0.041342f
C189 VN.n14 B 0.403734f
C190 VN.n15 B 0.041342f
C191 VN.n16 B 0.029453f
C192 VN.n17 B 0.029453f
C193 VN.n18 B 0.029453f
C194 VN.n19 B 0.04505f
C195 VN.n20 B 0.038632f
C196 VN.n21 B 0.403734f
C197 VN.n22 B 0.044052f
C198 VN.n23 B 0.029453f
C199 VN.n24 B 0.029453f
C200 VN.n25 B 0.029453f
C201 VN.n26 B 0.049154f
C202 VN.n27 B 0.035922f
C203 VN.n28 B 0.466588f
C204 VN.n29 B 0.029499f
C205 VN.n30 B 0.029453f
C206 VN.t9 B 1.08533f
C207 VN.n31 B 0.036843f
C208 VN.n32 B 0.029453f
C209 VN.t8 B 1.08533f
C210 VN.n33 B 0.040947f
C211 VN.n34 B 0.029453f
C212 VN.t7 B 1.08533f
C213 VN.n35 B 0.04505f
C214 VN.t4 B 1.19267f
C215 VN.n36 B 0.473045f
C216 VN.t6 B 1.08533f
C217 VN.n37 B 0.459075f
C218 VN.n38 B 0.038632f
C219 VN.n39 B 0.187852f
C220 VN.n40 B 0.029453f
C221 VN.n41 B 0.029453f
C222 VN.n42 B 0.040947f
C223 VN.n43 B 0.041342f
C224 VN.n44 B 0.403734f
C225 VN.n45 B 0.041342f
C226 VN.n46 B 0.029453f
C227 VN.n47 B 0.029453f
C228 VN.n48 B 0.029453f
C229 VN.n49 B 0.04505f
C230 VN.n50 B 0.038632f
C231 VN.n51 B 0.403734f
C232 VN.n52 B 0.044052f
C233 VN.n53 B 0.029453f
C234 VN.n54 B 0.029453f
C235 VN.n55 B 0.029453f
C236 VN.n56 B 0.049154f
C237 VN.n57 B 0.035922f
C238 VN.n58 B 0.466588f
C239 VN.n59 B 1.38688f
.ends

