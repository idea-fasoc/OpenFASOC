* NGSPICE file created from diff_pair_sample_1120.ext - technology: sky130A

.subckt diff_pair_sample_1120 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X1 VDD2.t7 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X2 VTAIL.t15 VN.t1 VDD2.t6 B.t21 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=1.8843 ps=11.75 w=11.42 l=0.54
X3 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=0 ps=0 w=11.42 l=0.54
X4 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X5 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X6 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=4.4538 ps=23.62 w=11.42 l=0.54
X7 VDD1.t7 VP.t1 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=4.4538 ps=23.62 w=11.42 l=0.54
X8 VDD1.t0 VP.t2 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X9 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=0 ps=0 w=11.42 l=0.54
X10 VTAIL.t4 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X11 VDD1.t4 VP.t3 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X12 VTAIL.t10 VP.t4 VDD1.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=1.8843 ps=11.75 w=11.42 l=0.54
X13 VDD2.t1 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=4.4538 ps=23.62 w=11.42 l=0.54
X14 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=0 ps=0 w=11.42 l=0.54
X15 VTAIL.t9 VP.t5 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=1.8843 ps=11.75 w=11.42 l=0.54
X16 VTAIL.t8 VP.t6 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=1.8843 ps=11.75 w=11.42 l=0.54
X17 VDD1.t1 VP.t7 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8843 pd=11.75 as=4.4538 ps=23.62 w=11.42 l=0.54
X18 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=1.8843 ps=11.75 w=11.42 l=0.54
X19 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.4538 pd=23.62 as=0 ps=0 w=11.42 l=0.54
R0 VP.n4 VP.t4 607.811
R1 VP.n11 VP.t6 582.418
R2 VP.n1 VP.t3 582.418
R3 VP.n16 VP.t5 582.418
R4 VP.n18 VP.t1 582.418
R5 VP.n8 VP.t7 582.418
R6 VP.n6 VP.t0 582.418
R7 VP.n5 VP.t2 582.418
R8 VP.n19 VP.n18 161.3
R9 VP.n6 VP.n3 161.3
R10 VP.n7 VP.n2 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n17 VP.n0 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n14 VP.n1 161.3
R15 VP.n13 VP.n12 161.3
R16 VP.n11 VP.n10 161.3
R17 VP.n16 VP.n1 48.2005
R18 VP.n6 VP.n5 48.2005
R19 VP.n4 VP.n3 45.0031
R20 VP.n12 VP.n11 41.6278
R21 VP.n18 VP.n17 41.6278
R22 VP.n8 VP.n7 41.6278
R23 VP.n10 VP.n9 40.7732
R24 VP.n5 VP.n4 15.6319
R25 VP.n12 VP.n1 6.57323
R26 VP.n17 VP.n16 6.57323
R27 VP.n7 VP.n6 6.57323
R28 VP.n3 VP.n2 0.189894
R29 VP.n9 VP.n2 0.189894
R30 VP.n13 VP.n10 0.189894
R31 VP.n14 VP.n13 0.189894
R32 VP.n15 VP.n14 0.189894
R33 VP.n15 VP.n0 0.189894
R34 VP.n19 VP.n0 0.189894
R35 VP VP.n19 0.0516364
R36 VDD1 VDD1.n0 62.911
R37 VDD1.n3 VDD1.n2 62.7973
R38 VDD1.n3 VDD1.n1 62.7973
R39 VDD1.n5 VDD1.n4 62.4776
R40 VDD1.n5 VDD1.n3 37.5181
R41 VDD1.n4 VDD1.t6 1.7343
R42 VDD1.n4 VDD1.t1 1.7343
R43 VDD1.n0 VDD1.t5 1.7343
R44 VDD1.n0 VDD1.t0 1.7343
R45 VDD1.n2 VDD1.t3 1.7343
R46 VDD1.n2 VDD1.t7 1.7343
R47 VDD1.n1 VDD1.t2 1.7343
R48 VDD1.n1 VDD1.t4 1.7343
R49 VDD1 VDD1.n5 0.31731
R50 VTAIL.n498 VTAIL.n442 289.615
R51 VTAIL.n58 VTAIL.n2 289.615
R52 VTAIL.n120 VTAIL.n64 289.615
R53 VTAIL.n184 VTAIL.n128 289.615
R54 VTAIL.n436 VTAIL.n380 289.615
R55 VTAIL.n372 VTAIL.n316 289.615
R56 VTAIL.n310 VTAIL.n254 289.615
R57 VTAIL.n246 VTAIL.n190 289.615
R58 VTAIL.n463 VTAIL.n462 185
R59 VTAIL.n465 VTAIL.n464 185
R60 VTAIL.n458 VTAIL.n457 185
R61 VTAIL.n471 VTAIL.n470 185
R62 VTAIL.n473 VTAIL.n472 185
R63 VTAIL.n454 VTAIL.n453 185
R64 VTAIL.n480 VTAIL.n479 185
R65 VTAIL.n481 VTAIL.n452 185
R66 VTAIL.n483 VTAIL.n482 185
R67 VTAIL.n450 VTAIL.n449 185
R68 VTAIL.n489 VTAIL.n488 185
R69 VTAIL.n491 VTAIL.n490 185
R70 VTAIL.n446 VTAIL.n445 185
R71 VTAIL.n497 VTAIL.n496 185
R72 VTAIL.n499 VTAIL.n498 185
R73 VTAIL.n23 VTAIL.n22 185
R74 VTAIL.n25 VTAIL.n24 185
R75 VTAIL.n18 VTAIL.n17 185
R76 VTAIL.n31 VTAIL.n30 185
R77 VTAIL.n33 VTAIL.n32 185
R78 VTAIL.n14 VTAIL.n13 185
R79 VTAIL.n40 VTAIL.n39 185
R80 VTAIL.n41 VTAIL.n12 185
R81 VTAIL.n43 VTAIL.n42 185
R82 VTAIL.n10 VTAIL.n9 185
R83 VTAIL.n49 VTAIL.n48 185
R84 VTAIL.n51 VTAIL.n50 185
R85 VTAIL.n6 VTAIL.n5 185
R86 VTAIL.n57 VTAIL.n56 185
R87 VTAIL.n59 VTAIL.n58 185
R88 VTAIL.n85 VTAIL.n84 185
R89 VTAIL.n87 VTAIL.n86 185
R90 VTAIL.n80 VTAIL.n79 185
R91 VTAIL.n93 VTAIL.n92 185
R92 VTAIL.n95 VTAIL.n94 185
R93 VTAIL.n76 VTAIL.n75 185
R94 VTAIL.n102 VTAIL.n101 185
R95 VTAIL.n103 VTAIL.n74 185
R96 VTAIL.n105 VTAIL.n104 185
R97 VTAIL.n72 VTAIL.n71 185
R98 VTAIL.n111 VTAIL.n110 185
R99 VTAIL.n113 VTAIL.n112 185
R100 VTAIL.n68 VTAIL.n67 185
R101 VTAIL.n119 VTAIL.n118 185
R102 VTAIL.n121 VTAIL.n120 185
R103 VTAIL.n149 VTAIL.n148 185
R104 VTAIL.n151 VTAIL.n150 185
R105 VTAIL.n144 VTAIL.n143 185
R106 VTAIL.n157 VTAIL.n156 185
R107 VTAIL.n159 VTAIL.n158 185
R108 VTAIL.n140 VTAIL.n139 185
R109 VTAIL.n166 VTAIL.n165 185
R110 VTAIL.n167 VTAIL.n138 185
R111 VTAIL.n169 VTAIL.n168 185
R112 VTAIL.n136 VTAIL.n135 185
R113 VTAIL.n175 VTAIL.n174 185
R114 VTAIL.n177 VTAIL.n176 185
R115 VTAIL.n132 VTAIL.n131 185
R116 VTAIL.n183 VTAIL.n182 185
R117 VTAIL.n185 VTAIL.n184 185
R118 VTAIL.n437 VTAIL.n436 185
R119 VTAIL.n435 VTAIL.n434 185
R120 VTAIL.n384 VTAIL.n383 185
R121 VTAIL.n429 VTAIL.n428 185
R122 VTAIL.n427 VTAIL.n426 185
R123 VTAIL.n388 VTAIL.n387 185
R124 VTAIL.n392 VTAIL.n390 185
R125 VTAIL.n421 VTAIL.n420 185
R126 VTAIL.n419 VTAIL.n418 185
R127 VTAIL.n394 VTAIL.n393 185
R128 VTAIL.n413 VTAIL.n412 185
R129 VTAIL.n411 VTAIL.n410 185
R130 VTAIL.n398 VTAIL.n397 185
R131 VTAIL.n405 VTAIL.n404 185
R132 VTAIL.n403 VTAIL.n402 185
R133 VTAIL.n373 VTAIL.n372 185
R134 VTAIL.n371 VTAIL.n370 185
R135 VTAIL.n320 VTAIL.n319 185
R136 VTAIL.n365 VTAIL.n364 185
R137 VTAIL.n363 VTAIL.n362 185
R138 VTAIL.n324 VTAIL.n323 185
R139 VTAIL.n328 VTAIL.n326 185
R140 VTAIL.n357 VTAIL.n356 185
R141 VTAIL.n355 VTAIL.n354 185
R142 VTAIL.n330 VTAIL.n329 185
R143 VTAIL.n349 VTAIL.n348 185
R144 VTAIL.n347 VTAIL.n346 185
R145 VTAIL.n334 VTAIL.n333 185
R146 VTAIL.n341 VTAIL.n340 185
R147 VTAIL.n339 VTAIL.n338 185
R148 VTAIL.n311 VTAIL.n310 185
R149 VTAIL.n309 VTAIL.n308 185
R150 VTAIL.n258 VTAIL.n257 185
R151 VTAIL.n303 VTAIL.n302 185
R152 VTAIL.n301 VTAIL.n300 185
R153 VTAIL.n262 VTAIL.n261 185
R154 VTAIL.n266 VTAIL.n264 185
R155 VTAIL.n295 VTAIL.n294 185
R156 VTAIL.n293 VTAIL.n292 185
R157 VTAIL.n268 VTAIL.n267 185
R158 VTAIL.n287 VTAIL.n286 185
R159 VTAIL.n285 VTAIL.n284 185
R160 VTAIL.n272 VTAIL.n271 185
R161 VTAIL.n279 VTAIL.n278 185
R162 VTAIL.n277 VTAIL.n276 185
R163 VTAIL.n247 VTAIL.n246 185
R164 VTAIL.n245 VTAIL.n244 185
R165 VTAIL.n194 VTAIL.n193 185
R166 VTAIL.n239 VTAIL.n238 185
R167 VTAIL.n237 VTAIL.n236 185
R168 VTAIL.n198 VTAIL.n197 185
R169 VTAIL.n202 VTAIL.n200 185
R170 VTAIL.n231 VTAIL.n230 185
R171 VTAIL.n229 VTAIL.n228 185
R172 VTAIL.n204 VTAIL.n203 185
R173 VTAIL.n223 VTAIL.n222 185
R174 VTAIL.n221 VTAIL.n220 185
R175 VTAIL.n208 VTAIL.n207 185
R176 VTAIL.n215 VTAIL.n214 185
R177 VTAIL.n213 VTAIL.n212 185
R178 VTAIL.n461 VTAIL.t5 149.524
R179 VTAIL.n21 VTAIL.t15 149.524
R180 VTAIL.n83 VTAIL.t13 149.524
R181 VTAIL.n147 VTAIL.t8 149.524
R182 VTAIL.n401 VTAIL.t7 149.524
R183 VTAIL.n337 VTAIL.t10 149.524
R184 VTAIL.n275 VTAIL.t1 149.524
R185 VTAIL.n211 VTAIL.t3 149.524
R186 VTAIL.n464 VTAIL.n463 104.615
R187 VTAIL.n464 VTAIL.n457 104.615
R188 VTAIL.n471 VTAIL.n457 104.615
R189 VTAIL.n472 VTAIL.n471 104.615
R190 VTAIL.n472 VTAIL.n453 104.615
R191 VTAIL.n480 VTAIL.n453 104.615
R192 VTAIL.n481 VTAIL.n480 104.615
R193 VTAIL.n482 VTAIL.n481 104.615
R194 VTAIL.n482 VTAIL.n449 104.615
R195 VTAIL.n489 VTAIL.n449 104.615
R196 VTAIL.n490 VTAIL.n489 104.615
R197 VTAIL.n490 VTAIL.n445 104.615
R198 VTAIL.n497 VTAIL.n445 104.615
R199 VTAIL.n498 VTAIL.n497 104.615
R200 VTAIL.n24 VTAIL.n23 104.615
R201 VTAIL.n24 VTAIL.n17 104.615
R202 VTAIL.n31 VTAIL.n17 104.615
R203 VTAIL.n32 VTAIL.n31 104.615
R204 VTAIL.n32 VTAIL.n13 104.615
R205 VTAIL.n40 VTAIL.n13 104.615
R206 VTAIL.n41 VTAIL.n40 104.615
R207 VTAIL.n42 VTAIL.n41 104.615
R208 VTAIL.n42 VTAIL.n9 104.615
R209 VTAIL.n49 VTAIL.n9 104.615
R210 VTAIL.n50 VTAIL.n49 104.615
R211 VTAIL.n50 VTAIL.n5 104.615
R212 VTAIL.n57 VTAIL.n5 104.615
R213 VTAIL.n58 VTAIL.n57 104.615
R214 VTAIL.n86 VTAIL.n85 104.615
R215 VTAIL.n86 VTAIL.n79 104.615
R216 VTAIL.n93 VTAIL.n79 104.615
R217 VTAIL.n94 VTAIL.n93 104.615
R218 VTAIL.n94 VTAIL.n75 104.615
R219 VTAIL.n102 VTAIL.n75 104.615
R220 VTAIL.n103 VTAIL.n102 104.615
R221 VTAIL.n104 VTAIL.n103 104.615
R222 VTAIL.n104 VTAIL.n71 104.615
R223 VTAIL.n111 VTAIL.n71 104.615
R224 VTAIL.n112 VTAIL.n111 104.615
R225 VTAIL.n112 VTAIL.n67 104.615
R226 VTAIL.n119 VTAIL.n67 104.615
R227 VTAIL.n120 VTAIL.n119 104.615
R228 VTAIL.n150 VTAIL.n149 104.615
R229 VTAIL.n150 VTAIL.n143 104.615
R230 VTAIL.n157 VTAIL.n143 104.615
R231 VTAIL.n158 VTAIL.n157 104.615
R232 VTAIL.n158 VTAIL.n139 104.615
R233 VTAIL.n166 VTAIL.n139 104.615
R234 VTAIL.n167 VTAIL.n166 104.615
R235 VTAIL.n168 VTAIL.n167 104.615
R236 VTAIL.n168 VTAIL.n135 104.615
R237 VTAIL.n175 VTAIL.n135 104.615
R238 VTAIL.n176 VTAIL.n175 104.615
R239 VTAIL.n176 VTAIL.n131 104.615
R240 VTAIL.n183 VTAIL.n131 104.615
R241 VTAIL.n184 VTAIL.n183 104.615
R242 VTAIL.n436 VTAIL.n435 104.615
R243 VTAIL.n435 VTAIL.n383 104.615
R244 VTAIL.n428 VTAIL.n383 104.615
R245 VTAIL.n428 VTAIL.n427 104.615
R246 VTAIL.n427 VTAIL.n387 104.615
R247 VTAIL.n392 VTAIL.n387 104.615
R248 VTAIL.n420 VTAIL.n392 104.615
R249 VTAIL.n420 VTAIL.n419 104.615
R250 VTAIL.n419 VTAIL.n393 104.615
R251 VTAIL.n412 VTAIL.n393 104.615
R252 VTAIL.n412 VTAIL.n411 104.615
R253 VTAIL.n411 VTAIL.n397 104.615
R254 VTAIL.n404 VTAIL.n397 104.615
R255 VTAIL.n404 VTAIL.n403 104.615
R256 VTAIL.n372 VTAIL.n371 104.615
R257 VTAIL.n371 VTAIL.n319 104.615
R258 VTAIL.n364 VTAIL.n319 104.615
R259 VTAIL.n364 VTAIL.n363 104.615
R260 VTAIL.n363 VTAIL.n323 104.615
R261 VTAIL.n328 VTAIL.n323 104.615
R262 VTAIL.n356 VTAIL.n328 104.615
R263 VTAIL.n356 VTAIL.n355 104.615
R264 VTAIL.n355 VTAIL.n329 104.615
R265 VTAIL.n348 VTAIL.n329 104.615
R266 VTAIL.n348 VTAIL.n347 104.615
R267 VTAIL.n347 VTAIL.n333 104.615
R268 VTAIL.n340 VTAIL.n333 104.615
R269 VTAIL.n340 VTAIL.n339 104.615
R270 VTAIL.n310 VTAIL.n309 104.615
R271 VTAIL.n309 VTAIL.n257 104.615
R272 VTAIL.n302 VTAIL.n257 104.615
R273 VTAIL.n302 VTAIL.n301 104.615
R274 VTAIL.n301 VTAIL.n261 104.615
R275 VTAIL.n266 VTAIL.n261 104.615
R276 VTAIL.n294 VTAIL.n266 104.615
R277 VTAIL.n294 VTAIL.n293 104.615
R278 VTAIL.n293 VTAIL.n267 104.615
R279 VTAIL.n286 VTAIL.n267 104.615
R280 VTAIL.n286 VTAIL.n285 104.615
R281 VTAIL.n285 VTAIL.n271 104.615
R282 VTAIL.n278 VTAIL.n271 104.615
R283 VTAIL.n278 VTAIL.n277 104.615
R284 VTAIL.n246 VTAIL.n245 104.615
R285 VTAIL.n245 VTAIL.n193 104.615
R286 VTAIL.n238 VTAIL.n193 104.615
R287 VTAIL.n238 VTAIL.n237 104.615
R288 VTAIL.n237 VTAIL.n197 104.615
R289 VTAIL.n202 VTAIL.n197 104.615
R290 VTAIL.n230 VTAIL.n202 104.615
R291 VTAIL.n230 VTAIL.n229 104.615
R292 VTAIL.n229 VTAIL.n203 104.615
R293 VTAIL.n222 VTAIL.n203 104.615
R294 VTAIL.n222 VTAIL.n221 104.615
R295 VTAIL.n221 VTAIL.n207 104.615
R296 VTAIL.n214 VTAIL.n207 104.615
R297 VTAIL.n214 VTAIL.n213 104.615
R298 VTAIL.n463 VTAIL.t5 52.3082
R299 VTAIL.n23 VTAIL.t15 52.3082
R300 VTAIL.n85 VTAIL.t13 52.3082
R301 VTAIL.n149 VTAIL.t8 52.3082
R302 VTAIL.n403 VTAIL.t7 52.3082
R303 VTAIL.n339 VTAIL.t10 52.3082
R304 VTAIL.n277 VTAIL.t1 52.3082
R305 VTAIL.n213 VTAIL.t3 52.3082
R306 VTAIL.n379 VTAIL.n378 45.799
R307 VTAIL.n253 VTAIL.n252 45.799
R308 VTAIL.n1 VTAIL.n0 45.7988
R309 VTAIL.n127 VTAIL.n126 45.7988
R310 VTAIL.n503 VTAIL.n502 32.5732
R311 VTAIL.n63 VTAIL.n62 32.5732
R312 VTAIL.n125 VTAIL.n124 32.5732
R313 VTAIL.n189 VTAIL.n188 32.5732
R314 VTAIL.n441 VTAIL.n440 32.5732
R315 VTAIL.n377 VTAIL.n376 32.5732
R316 VTAIL.n315 VTAIL.n314 32.5732
R317 VTAIL.n251 VTAIL.n250 32.5732
R318 VTAIL.n503 VTAIL.n441 22.9617
R319 VTAIL.n251 VTAIL.n189 22.9617
R320 VTAIL.n483 VTAIL.n450 13.1884
R321 VTAIL.n43 VTAIL.n10 13.1884
R322 VTAIL.n105 VTAIL.n72 13.1884
R323 VTAIL.n169 VTAIL.n136 13.1884
R324 VTAIL.n390 VTAIL.n388 13.1884
R325 VTAIL.n326 VTAIL.n324 13.1884
R326 VTAIL.n264 VTAIL.n262 13.1884
R327 VTAIL.n200 VTAIL.n198 13.1884
R328 VTAIL.n484 VTAIL.n452 12.8005
R329 VTAIL.n488 VTAIL.n487 12.8005
R330 VTAIL.n44 VTAIL.n12 12.8005
R331 VTAIL.n48 VTAIL.n47 12.8005
R332 VTAIL.n106 VTAIL.n74 12.8005
R333 VTAIL.n110 VTAIL.n109 12.8005
R334 VTAIL.n170 VTAIL.n138 12.8005
R335 VTAIL.n174 VTAIL.n173 12.8005
R336 VTAIL.n426 VTAIL.n425 12.8005
R337 VTAIL.n422 VTAIL.n421 12.8005
R338 VTAIL.n362 VTAIL.n361 12.8005
R339 VTAIL.n358 VTAIL.n357 12.8005
R340 VTAIL.n300 VTAIL.n299 12.8005
R341 VTAIL.n296 VTAIL.n295 12.8005
R342 VTAIL.n236 VTAIL.n235 12.8005
R343 VTAIL.n232 VTAIL.n231 12.8005
R344 VTAIL.n479 VTAIL.n478 12.0247
R345 VTAIL.n491 VTAIL.n448 12.0247
R346 VTAIL.n39 VTAIL.n38 12.0247
R347 VTAIL.n51 VTAIL.n8 12.0247
R348 VTAIL.n101 VTAIL.n100 12.0247
R349 VTAIL.n113 VTAIL.n70 12.0247
R350 VTAIL.n165 VTAIL.n164 12.0247
R351 VTAIL.n177 VTAIL.n134 12.0247
R352 VTAIL.n429 VTAIL.n386 12.0247
R353 VTAIL.n418 VTAIL.n391 12.0247
R354 VTAIL.n365 VTAIL.n322 12.0247
R355 VTAIL.n354 VTAIL.n327 12.0247
R356 VTAIL.n303 VTAIL.n260 12.0247
R357 VTAIL.n292 VTAIL.n265 12.0247
R358 VTAIL.n239 VTAIL.n196 12.0247
R359 VTAIL.n228 VTAIL.n201 12.0247
R360 VTAIL.n477 VTAIL.n454 11.249
R361 VTAIL.n492 VTAIL.n446 11.249
R362 VTAIL.n37 VTAIL.n14 11.249
R363 VTAIL.n52 VTAIL.n6 11.249
R364 VTAIL.n99 VTAIL.n76 11.249
R365 VTAIL.n114 VTAIL.n68 11.249
R366 VTAIL.n163 VTAIL.n140 11.249
R367 VTAIL.n178 VTAIL.n132 11.249
R368 VTAIL.n430 VTAIL.n384 11.249
R369 VTAIL.n417 VTAIL.n394 11.249
R370 VTAIL.n366 VTAIL.n320 11.249
R371 VTAIL.n353 VTAIL.n330 11.249
R372 VTAIL.n304 VTAIL.n258 11.249
R373 VTAIL.n291 VTAIL.n268 11.249
R374 VTAIL.n240 VTAIL.n194 11.249
R375 VTAIL.n227 VTAIL.n204 11.249
R376 VTAIL.n474 VTAIL.n473 10.4732
R377 VTAIL.n496 VTAIL.n495 10.4732
R378 VTAIL.n34 VTAIL.n33 10.4732
R379 VTAIL.n56 VTAIL.n55 10.4732
R380 VTAIL.n96 VTAIL.n95 10.4732
R381 VTAIL.n118 VTAIL.n117 10.4732
R382 VTAIL.n160 VTAIL.n159 10.4732
R383 VTAIL.n182 VTAIL.n181 10.4732
R384 VTAIL.n434 VTAIL.n433 10.4732
R385 VTAIL.n414 VTAIL.n413 10.4732
R386 VTAIL.n370 VTAIL.n369 10.4732
R387 VTAIL.n350 VTAIL.n349 10.4732
R388 VTAIL.n308 VTAIL.n307 10.4732
R389 VTAIL.n288 VTAIL.n287 10.4732
R390 VTAIL.n244 VTAIL.n243 10.4732
R391 VTAIL.n224 VTAIL.n223 10.4732
R392 VTAIL.n462 VTAIL.n461 10.2747
R393 VTAIL.n22 VTAIL.n21 10.2747
R394 VTAIL.n84 VTAIL.n83 10.2747
R395 VTAIL.n148 VTAIL.n147 10.2747
R396 VTAIL.n402 VTAIL.n401 10.2747
R397 VTAIL.n338 VTAIL.n337 10.2747
R398 VTAIL.n276 VTAIL.n275 10.2747
R399 VTAIL.n212 VTAIL.n211 10.2747
R400 VTAIL.n470 VTAIL.n456 9.69747
R401 VTAIL.n499 VTAIL.n444 9.69747
R402 VTAIL.n30 VTAIL.n16 9.69747
R403 VTAIL.n59 VTAIL.n4 9.69747
R404 VTAIL.n92 VTAIL.n78 9.69747
R405 VTAIL.n121 VTAIL.n66 9.69747
R406 VTAIL.n156 VTAIL.n142 9.69747
R407 VTAIL.n185 VTAIL.n130 9.69747
R408 VTAIL.n437 VTAIL.n382 9.69747
R409 VTAIL.n410 VTAIL.n396 9.69747
R410 VTAIL.n373 VTAIL.n318 9.69747
R411 VTAIL.n346 VTAIL.n332 9.69747
R412 VTAIL.n311 VTAIL.n256 9.69747
R413 VTAIL.n284 VTAIL.n270 9.69747
R414 VTAIL.n247 VTAIL.n192 9.69747
R415 VTAIL.n220 VTAIL.n206 9.69747
R416 VTAIL.n502 VTAIL.n501 9.45567
R417 VTAIL.n62 VTAIL.n61 9.45567
R418 VTAIL.n124 VTAIL.n123 9.45567
R419 VTAIL.n188 VTAIL.n187 9.45567
R420 VTAIL.n440 VTAIL.n439 9.45567
R421 VTAIL.n376 VTAIL.n375 9.45567
R422 VTAIL.n314 VTAIL.n313 9.45567
R423 VTAIL.n250 VTAIL.n249 9.45567
R424 VTAIL.n501 VTAIL.n500 9.3005
R425 VTAIL.n444 VTAIL.n443 9.3005
R426 VTAIL.n495 VTAIL.n494 9.3005
R427 VTAIL.n493 VTAIL.n492 9.3005
R428 VTAIL.n448 VTAIL.n447 9.3005
R429 VTAIL.n487 VTAIL.n486 9.3005
R430 VTAIL.n460 VTAIL.n459 9.3005
R431 VTAIL.n467 VTAIL.n466 9.3005
R432 VTAIL.n469 VTAIL.n468 9.3005
R433 VTAIL.n456 VTAIL.n455 9.3005
R434 VTAIL.n475 VTAIL.n474 9.3005
R435 VTAIL.n477 VTAIL.n476 9.3005
R436 VTAIL.n478 VTAIL.n451 9.3005
R437 VTAIL.n485 VTAIL.n484 9.3005
R438 VTAIL.n61 VTAIL.n60 9.3005
R439 VTAIL.n4 VTAIL.n3 9.3005
R440 VTAIL.n55 VTAIL.n54 9.3005
R441 VTAIL.n53 VTAIL.n52 9.3005
R442 VTAIL.n8 VTAIL.n7 9.3005
R443 VTAIL.n47 VTAIL.n46 9.3005
R444 VTAIL.n20 VTAIL.n19 9.3005
R445 VTAIL.n27 VTAIL.n26 9.3005
R446 VTAIL.n29 VTAIL.n28 9.3005
R447 VTAIL.n16 VTAIL.n15 9.3005
R448 VTAIL.n35 VTAIL.n34 9.3005
R449 VTAIL.n37 VTAIL.n36 9.3005
R450 VTAIL.n38 VTAIL.n11 9.3005
R451 VTAIL.n45 VTAIL.n44 9.3005
R452 VTAIL.n123 VTAIL.n122 9.3005
R453 VTAIL.n66 VTAIL.n65 9.3005
R454 VTAIL.n117 VTAIL.n116 9.3005
R455 VTAIL.n115 VTAIL.n114 9.3005
R456 VTAIL.n70 VTAIL.n69 9.3005
R457 VTAIL.n109 VTAIL.n108 9.3005
R458 VTAIL.n82 VTAIL.n81 9.3005
R459 VTAIL.n89 VTAIL.n88 9.3005
R460 VTAIL.n91 VTAIL.n90 9.3005
R461 VTAIL.n78 VTAIL.n77 9.3005
R462 VTAIL.n97 VTAIL.n96 9.3005
R463 VTAIL.n99 VTAIL.n98 9.3005
R464 VTAIL.n100 VTAIL.n73 9.3005
R465 VTAIL.n107 VTAIL.n106 9.3005
R466 VTAIL.n187 VTAIL.n186 9.3005
R467 VTAIL.n130 VTAIL.n129 9.3005
R468 VTAIL.n181 VTAIL.n180 9.3005
R469 VTAIL.n179 VTAIL.n178 9.3005
R470 VTAIL.n134 VTAIL.n133 9.3005
R471 VTAIL.n173 VTAIL.n172 9.3005
R472 VTAIL.n146 VTAIL.n145 9.3005
R473 VTAIL.n153 VTAIL.n152 9.3005
R474 VTAIL.n155 VTAIL.n154 9.3005
R475 VTAIL.n142 VTAIL.n141 9.3005
R476 VTAIL.n161 VTAIL.n160 9.3005
R477 VTAIL.n163 VTAIL.n162 9.3005
R478 VTAIL.n164 VTAIL.n137 9.3005
R479 VTAIL.n171 VTAIL.n170 9.3005
R480 VTAIL.n400 VTAIL.n399 9.3005
R481 VTAIL.n407 VTAIL.n406 9.3005
R482 VTAIL.n409 VTAIL.n408 9.3005
R483 VTAIL.n396 VTAIL.n395 9.3005
R484 VTAIL.n415 VTAIL.n414 9.3005
R485 VTAIL.n417 VTAIL.n416 9.3005
R486 VTAIL.n391 VTAIL.n389 9.3005
R487 VTAIL.n423 VTAIL.n422 9.3005
R488 VTAIL.n439 VTAIL.n438 9.3005
R489 VTAIL.n382 VTAIL.n381 9.3005
R490 VTAIL.n433 VTAIL.n432 9.3005
R491 VTAIL.n431 VTAIL.n430 9.3005
R492 VTAIL.n386 VTAIL.n385 9.3005
R493 VTAIL.n425 VTAIL.n424 9.3005
R494 VTAIL.n336 VTAIL.n335 9.3005
R495 VTAIL.n343 VTAIL.n342 9.3005
R496 VTAIL.n345 VTAIL.n344 9.3005
R497 VTAIL.n332 VTAIL.n331 9.3005
R498 VTAIL.n351 VTAIL.n350 9.3005
R499 VTAIL.n353 VTAIL.n352 9.3005
R500 VTAIL.n327 VTAIL.n325 9.3005
R501 VTAIL.n359 VTAIL.n358 9.3005
R502 VTAIL.n375 VTAIL.n374 9.3005
R503 VTAIL.n318 VTAIL.n317 9.3005
R504 VTAIL.n369 VTAIL.n368 9.3005
R505 VTAIL.n367 VTAIL.n366 9.3005
R506 VTAIL.n322 VTAIL.n321 9.3005
R507 VTAIL.n361 VTAIL.n360 9.3005
R508 VTAIL.n274 VTAIL.n273 9.3005
R509 VTAIL.n281 VTAIL.n280 9.3005
R510 VTAIL.n283 VTAIL.n282 9.3005
R511 VTAIL.n270 VTAIL.n269 9.3005
R512 VTAIL.n289 VTAIL.n288 9.3005
R513 VTAIL.n291 VTAIL.n290 9.3005
R514 VTAIL.n265 VTAIL.n263 9.3005
R515 VTAIL.n297 VTAIL.n296 9.3005
R516 VTAIL.n313 VTAIL.n312 9.3005
R517 VTAIL.n256 VTAIL.n255 9.3005
R518 VTAIL.n307 VTAIL.n306 9.3005
R519 VTAIL.n305 VTAIL.n304 9.3005
R520 VTAIL.n260 VTAIL.n259 9.3005
R521 VTAIL.n299 VTAIL.n298 9.3005
R522 VTAIL.n210 VTAIL.n209 9.3005
R523 VTAIL.n217 VTAIL.n216 9.3005
R524 VTAIL.n219 VTAIL.n218 9.3005
R525 VTAIL.n206 VTAIL.n205 9.3005
R526 VTAIL.n225 VTAIL.n224 9.3005
R527 VTAIL.n227 VTAIL.n226 9.3005
R528 VTAIL.n201 VTAIL.n199 9.3005
R529 VTAIL.n233 VTAIL.n232 9.3005
R530 VTAIL.n249 VTAIL.n248 9.3005
R531 VTAIL.n192 VTAIL.n191 9.3005
R532 VTAIL.n243 VTAIL.n242 9.3005
R533 VTAIL.n241 VTAIL.n240 9.3005
R534 VTAIL.n196 VTAIL.n195 9.3005
R535 VTAIL.n235 VTAIL.n234 9.3005
R536 VTAIL.n469 VTAIL.n458 8.92171
R537 VTAIL.n500 VTAIL.n442 8.92171
R538 VTAIL.n29 VTAIL.n18 8.92171
R539 VTAIL.n60 VTAIL.n2 8.92171
R540 VTAIL.n91 VTAIL.n80 8.92171
R541 VTAIL.n122 VTAIL.n64 8.92171
R542 VTAIL.n155 VTAIL.n144 8.92171
R543 VTAIL.n186 VTAIL.n128 8.92171
R544 VTAIL.n438 VTAIL.n380 8.92171
R545 VTAIL.n409 VTAIL.n398 8.92171
R546 VTAIL.n374 VTAIL.n316 8.92171
R547 VTAIL.n345 VTAIL.n334 8.92171
R548 VTAIL.n312 VTAIL.n254 8.92171
R549 VTAIL.n283 VTAIL.n272 8.92171
R550 VTAIL.n248 VTAIL.n190 8.92171
R551 VTAIL.n219 VTAIL.n208 8.92171
R552 VTAIL.n466 VTAIL.n465 8.14595
R553 VTAIL.n26 VTAIL.n25 8.14595
R554 VTAIL.n88 VTAIL.n87 8.14595
R555 VTAIL.n152 VTAIL.n151 8.14595
R556 VTAIL.n406 VTAIL.n405 8.14595
R557 VTAIL.n342 VTAIL.n341 8.14595
R558 VTAIL.n280 VTAIL.n279 8.14595
R559 VTAIL.n216 VTAIL.n215 8.14595
R560 VTAIL.n462 VTAIL.n460 7.3702
R561 VTAIL.n22 VTAIL.n20 7.3702
R562 VTAIL.n84 VTAIL.n82 7.3702
R563 VTAIL.n148 VTAIL.n146 7.3702
R564 VTAIL.n402 VTAIL.n400 7.3702
R565 VTAIL.n338 VTAIL.n336 7.3702
R566 VTAIL.n276 VTAIL.n274 7.3702
R567 VTAIL.n212 VTAIL.n210 7.3702
R568 VTAIL.n465 VTAIL.n460 5.81868
R569 VTAIL.n25 VTAIL.n20 5.81868
R570 VTAIL.n87 VTAIL.n82 5.81868
R571 VTAIL.n151 VTAIL.n146 5.81868
R572 VTAIL.n405 VTAIL.n400 5.81868
R573 VTAIL.n341 VTAIL.n336 5.81868
R574 VTAIL.n279 VTAIL.n274 5.81868
R575 VTAIL.n215 VTAIL.n210 5.81868
R576 VTAIL.n466 VTAIL.n458 5.04292
R577 VTAIL.n502 VTAIL.n442 5.04292
R578 VTAIL.n26 VTAIL.n18 5.04292
R579 VTAIL.n62 VTAIL.n2 5.04292
R580 VTAIL.n88 VTAIL.n80 5.04292
R581 VTAIL.n124 VTAIL.n64 5.04292
R582 VTAIL.n152 VTAIL.n144 5.04292
R583 VTAIL.n188 VTAIL.n128 5.04292
R584 VTAIL.n440 VTAIL.n380 5.04292
R585 VTAIL.n406 VTAIL.n398 5.04292
R586 VTAIL.n376 VTAIL.n316 5.04292
R587 VTAIL.n342 VTAIL.n334 5.04292
R588 VTAIL.n314 VTAIL.n254 5.04292
R589 VTAIL.n280 VTAIL.n272 5.04292
R590 VTAIL.n250 VTAIL.n190 5.04292
R591 VTAIL.n216 VTAIL.n208 5.04292
R592 VTAIL.n470 VTAIL.n469 4.26717
R593 VTAIL.n500 VTAIL.n499 4.26717
R594 VTAIL.n30 VTAIL.n29 4.26717
R595 VTAIL.n60 VTAIL.n59 4.26717
R596 VTAIL.n92 VTAIL.n91 4.26717
R597 VTAIL.n122 VTAIL.n121 4.26717
R598 VTAIL.n156 VTAIL.n155 4.26717
R599 VTAIL.n186 VTAIL.n185 4.26717
R600 VTAIL.n438 VTAIL.n437 4.26717
R601 VTAIL.n410 VTAIL.n409 4.26717
R602 VTAIL.n374 VTAIL.n373 4.26717
R603 VTAIL.n346 VTAIL.n345 4.26717
R604 VTAIL.n312 VTAIL.n311 4.26717
R605 VTAIL.n284 VTAIL.n283 4.26717
R606 VTAIL.n248 VTAIL.n247 4.26717
R607 VTAIL.n220 VTAIL.n219 4.26717
R608 VTAIL.n473 VTAIL.n456 3.49141
R609 VTAIL.n496 VTAIL.n444 3.49141
R610 VTAIL.n33 VTAIL.n16 3.49141
R611 VTAIL.n56 VTAIL.n4 3.49141
R612 VTAIL.n95 VTAIL.n78 3.49141
R613 VTAIL.n118 VTAIL.n66 3.49141
R614 VTAIL.n159 VTAIL.n142 3.49141
R615 VTAIL.n182 VTAIL.n130 3.49141
R616 VTAIL.n434 VTAIL.n382 3.49141
R617 VTAIL.n413 VTAIL.n396 3.49141
R618 VTAIL.n370 VTAIL.n318 3.49141
R619 VTAIL.n349 VTAIL.n332 3.49141
R620 VTAIL.n308 VTAIL.n256 3.49141
R621 VTAIL.n287 VTAIL.n270 3.49141
R622 VTAIL.n244 VTAIL.n192 3.49141
R623 VTAIL.n223 VTAIL.n206 3.49141
R624 VTAIL.n461 VTAIL.n459 2.84303
R625 VTAIL.n21 VTAIL.n19 2.84303
R626 VTAIL.n83 VTAIL.n81 2.84303
R627 VTAIL.n147 VTAIL.n145 2.84303
R628 VTAIL.n401 VTAIL.n399 2.84303
R629 VTAIL.n337 VTAIL.n335 2.84303
R630 VTAIL.n275 VTAIL.n273 2.84303
R631 VTAIL.n211 VTAIL.n209 2.84303
R632 VTAIL.n474 VTAIL.n454 2.71565
R633 VTAIL.n495 VTAIL.n446 2.71565
R634 VTAIL.n34 VTAIL.n14 2.71565
R635 VTAIL.n55 VTAIL.n6 2.71565
R636 VTAIL.n96 VTAIL.n76 2.71565
R637 VTAIL.n117 VTAIL.n68 2.71565
R638 VTAIL.n160 VTAIL.n140 2.71565
R639 VTAIL.n181 VTAIL.n132 2.71565
R640 VTAIL.n433 VTAIL.n384 2.71565
R641 VTAIL.n414 VTAIL.n394 2.71565
R642 VTAIL.n369 VTAIL.n320 2.71565
R643 VTAIL.n350 VTAIL.n330 2.71565
R644 VTAIL.n307 VTAIL.n258 2.71565
R645 VTAIL.n288 VTAIL.n268 2.71565
R646 VTAIL.n243 VTAIL.n194 2.71565
R647 VTAIL.n224 VTAIL.n204 2.71565
R648 VTAIL.n479 VTAIL.n477 1.93989
R649 VTAIL.n492 VTAIL.n491 1.93989
R650 VTAIL.n39 VTAIL.n37 1.93989
R651 VTAIL.n52 VTAIL.n51 1.93989
R652 VTAIL.n101 VTAIL.n99 1.93989
R653 VTAIL.n114 VTAIL.n113 1.93989
R654 VTAIL.n165 VTAIL.n163 1.93989
R655 VTAIL.n178 VTAIL.n177 1.93989
R656 VTAIL.n430 VTAIL.n429 1.93989
R657 VTAIL.n418 VTAIL.n417 1.93989
R658 VTAIL.n366 VTAIL.n365 1.93989
R659 VTAIL.n354 VTAIL.n353 1.93989
R660 VTAIL.n304 VTAIL.n303 1.93989
R661 VTAIL.n292 VTAIL.n291 1.93989
R662 VTAIL.n240 VTAIL.n239 1.93989
R663 VTAIL.n228 VTAIL.n227 1.93989
R664 VTAIL.n0 VTAIL.t6 1.7343
R665 VTAIL.n0 VTAIL.t2 1.7343
R666 VTAIL.n126 VTAIL.t11 1.7343
R667 VTAIL.n126 VTAIL.t9 1.7343
R668 VTAIL.n378 VTAIL.t12 1.7343
R669 VTAIL.n378 VTAIL.t14 1.7343
R670 VTAIL.n252 VTAIL.t0 1.7343
R671 VTAIL.n252 VTAIL.t4 1.7343
R672 VTAIL.n478 VTAIL.n452 1.16414
R673 VTAIL.n488 VTAIL.n448 1.16414
R674 VTAIL.n38 VTAIL.n12 1.16414
R675 VTAIL.n48 VTAIL.n8 1.16414
R676 VTAIL.n100 VTAIL.n74 1.16414
R677 VTAIL.n110 VTAIL.n70 1.16414
R678 VTAIL.n164 VTAIL.n138 1.16414
R679 VTAIL.n174 VTAIL.n134 1.16414
R680 VTAIL.n426 VTAIL.n386 1.16414
R681 VTAIL.n421 VTAIL.n391 1.16414
R682 VTAIL.n362 VTAIL.n322 1.16414
R683 VTAIL.n357 VTAIL.n327 1.16414
R684 VTAIL.n300 VTAIL.n260 1.16414
R685 VTAIL.n295 VTAIL.n265 1.16414
R686 VTAIL.n236 VTAIL.n196 1.16414
R687 VTAIL.n231 VTAIL.n201 1.16414
R688 VTAIL.n253 VTAIL.n251 0.7505
R689 VTAIL.n315 VTAIL.n253 0.7505
R690 VTAIL.n379 VTAIL.n377 0.7505
R691 VTAIL.n441 VTAIL.n379 0.7505
R692 VTAIL.n189 VTAIL.n127 0.7505
R693 VTAIL.n127 VTAIL.n125 0.7505
R694 VTAIL.n63 VTAIL.n1 0.7505
R695 VTAIL VTAIL.n503 0.69231
R696 VTAIL.n377 VTAIL.n315 0.470328
R697 VTAIL.n125 VTAIL.n63 0.470328
R698 VTAIL.n484 VTAIL.n483 0.388379
R699 VTAIL.n487 VTAIL.n450 0.388379
R700 VTAIL.n44 VTAIL.n43 0.388379
R701 VTAIL.n47 VTAIL.n10 0.388379
R702 VTAIL.n106 VTAIL.n105 0.388379
R703 VTAIL.n109 VTAIL.n72 0.388379
R704 VTAIL.n170 VTAIL.n169 0.388379
R705 VTAIL.n173 VTAIL.n136 0.388379
R706 VTAIL.n425 VTAIL.n388 0.388379
R707 VTAIL.n422 VTAIL.n390 0.388379
R708 VTAIL.n361 VTAIL.n324 0.388379
R709 VTAIL.n358 VTAIL.n326 0.388379
R710 VTAIL.n299 VTAIL.n262 0.388379
R711 VTAIL.n296 VTAIL.n264 0.388379
R712 VTAIL.n235 VTAIL.n198 0.388379
R713 VTAIL.n232 VTAIL.n200 0.388379
R714 VTAIL.n467 VTAIL.n459 0.155672
R715 VTAIL.n468 VTAIL.n467 0.155672
R716 VTAIL.n468 VTAIL.n455 0.155672
R717 VTAIL.n475 VTAIL.n455 0.155672
R718 VTAIL.n476 VTAIL.n475 0.155672
R719 VTAIL.n476 VTAIL.n451 0.155672
R720 VTAIL.n485 VTAIL.n451 0.155672
R721 VTAIL.n486 VTAIL.n485 0.155672
R722 VTAIL.n486 VTAIL.n447 0.155672
R723 VTAIL.n493 VTAIL.n447 0.155672
R724 VTAIL.n494 VTAIL.n493 0.155672
R725 VTAIL.n494 VTAIL.n443 0.155672
R726 VTAIL.n501 VTAIL.n443 0.155672
R727 VTAIL.n27 VTAIL.n19 0.155672
R728 VTAIL.n28 VTAIL.n27 0.155672
R729 VTAIL.n28 VTAIL.n15 0.155672
R730 VTAIL.n35 VTAIL.n15 0.155672
R731 VTAIL.n36 VTAIL.n35 0.155672
R732 VTAIL.n36 VTAIL.n11 0.155672
R733 VTAIL.n45 VTAIL.n11 0.155672
R734 VTAIL.n46 VTAIL.n45 0.155672
R735 VTAIL.n46 VTAIL.n7 0.155672
R736 VTAIL.n53 VTAIL.n7 0.155672
R737 VTAIL.n54 VTAIL.n53 0.155672
R738 VTAIL.n54 VTAIL.n3 0.155672
R739 VTAIL.n61 VTAIL.n3 0.155672
R740 VTAIL.n89 VTAIL.n81 0.155672
R741 VTAIL.n90 VTAIL.n89 0.155672
R742 VTAIL.n90 VTAIL.n77 0.155672
R743 VTAIL.n97 VTAIL.n77 0.155672
R744 VTAIL.n98 VTAIL.n97 0.155672
R745 VTAIL.n98 VTAIL.n73 0.155672
R746 VTAIL.n107 VTAIL.n73 0.155672
R747 VTAIL.n108 VTAIL.n107 0.155672
R748 VTAIL.n108 VTAIL.n69 0.155672
R749 VTAIL.n115 VTAIL.n69 0.155672
R750 VTAIL.n116 VTAIL.n115 0.155672
R751 VTAIL.n116 VTAIL.n65 0.155672
R752 VTAIL.n123 VTAIL.n65 0.155672
R753 VTAIL.n153 VTAIL.n145 0.155672
R754 VTAIL.n154 VTAIL.n153 0.155672
R755 VTAIL.n154 VTAIL.n141 0.155672
R756 VTAIL.n161 VTAIL.n141 0.155672
R757 VTAIL.n162 VTAIL.n161 0.155672
R758 VTAIL.n162 VTAIL.n137 0.155672
R759 VTAIL.n171 VTAIL.n137 0.155672
R760 VTAIL.n172 VTAIL.n171 0.155672
R761 VTAIL.n172 VTAIL.n133 0.155672
R762 VTAIL.n179 VTAIL.n133 0.155672
R763 VTAIL.n180 VTAIL.n179 0.155672
R764 VTAIL.n180 VTAIL.n129 0.155672
R765 VTAIL.n187 VTAIL.n129 0.155672
R766 VTAIL.n439 VTAIL.n381 0.155672
R767 VTAIL.n432 VTAIL.n381 0.155672
R768 VTAIL.n432 VTAIL.n431 0.155672
R769 VTAIL.n431 VTAIL.n385 0.155672
R770 VTAIL.n424 VTAIL.n385 0.155672
R771 VTAIL.n424 VTAIL.n423 0.155672
R772 VTAIL.n423 VTAIL.n389 0.155672
R773 VTAIL.n416 VTAIL.n389 0.155672
R774 VTAIL.n416 VTAIL.n415 0.155672
R775 VTAIL.n415 VTAIL.n395 0.155672
R776 VTAIL.n408 VTAIL.n395 0.155672
R777 VTAIL.n408 VTAIL.n407 0.155672
R778 VTAIL.n407 VTAIL.n399 0.155672
R779 VTAIL.n375 VTAIL.n317 0.155672
R780 VTAIL.n368 VTAIL.n317 0.155672
R781 VTAIL.n368 VTAIL.n367 0.155672
R782 VTAIL.n367 VTAIL.n321 0.155672
R783 VTAIL.n360 VTAIL.n321 0.155672
R784 VTAIL.n360 VTAIL.n359 0.155672
R785 VTAIL.n359 VTAIL.n325 0.155672
R786 VTAIL.n352 VTAIL.n325 0.155672
R787 VTAIL.n352 VTAIL.n351 0.155672
R788 VTAIL.n351 VTAIL.n331 0.155672
R789 VTAIL.n344 VTAIL.n331 0.155672
R790 VTAIL.n344 VTAIL.n343 0.155672
R791 VTAIL.n343 VTAIL.n335 0.155672
R792 VTAIL.n313 VTAIL.n255 0.155672
R793 VTAIL.n306 VTAIL.n255 0.155672
R794 VTAIL.n306 VTAIL.n305 0.155672
R795 VTAIL.n305 VTAIL.n259 0.155672
R796 VTAIL.n298 VTAIL.n259 0.155672
R797 VTAIL.n298 VTAIL.n297 0.155672
R798 VTAIL.n297 VTAIL.n263 0.155672
R799 VTAIL.n290 VTAIL.n263 0.155672
R800 VTAIL.n290 VTAIL.n289 0.155672
R801 VTAIL.n289 VTAIL.n269 0.155672
R802 VTAIL.n282 VTAIL.n269 0.155672
R803 VTAIL.n282 VTAIL.n281 0.155672
R804 VTAIL.n281 VTAIL.n273 0.155672
R805 VTAIL.n249 VTAIL.n191 0.155672
R806 VTAIL.n242 VTAIL.n191 0.155672
R807 VTAIL.n242 VTAIL.n241 0.155672
R808 VTAIL.n241 VTAIL.n195 0.155672
R809 VTAIL.n234 VTAIL.n195 0.155672
R810 VTAIL.n234 VTAIL.n233 0.155672
R811 VTAIL.n233 VTAIL.n199 0.155672
R812 VTAIL.n226 VTAIL.n199 0.155672
R813 VTAIL.n226 VTAIL.n225 0.155672
R814 VTAIL.n225 VTAIL.n205 0.155672
R815 VTAIL.n218 VTAIL.n205 0.155672
R816 VTAIL.n218 VTAIL.n217 0.155672
R817 VTAIL.n217 VTAIL.n209 0.155672
R818 VTAIL VTAIL.n1 0.0586897
R819 B.n354 B.t7 715.186
R820 B.n352 B.t15 715.186
R821 B.n89 B.t18 715.186
R822 B.n87 B.t11 715.186
R823 B.n626 B.n625 585
R824 B.n627 B.n626 585
R825 B.n267 B.n86 585
R826 B.n266 B.n265 585
R827 B.n264 B.n263 585
R828 B.n262 B.n261 585
R829 B.n260 B.n259 585
R830 B.n258 B.n257 585
R831 B.n256 B.n255 585
R832 B.n254 B.n253 585
R833 B.n252 B.n251 585
R834 B.n250 B.n249 585
R835 B.n248 B.n247 585
R836 B.n246 B.n245 585
R837 B.n244 B.n243 585
R838 B.n242 B.n241 585
R839 B.n240 B.n239 585
R840 B.n238 B.n237 585
R841 B.n236 B.n235 585
R842 B.n234 B.n233 585
R843 B.n232 B.n231 585
R844 B.n230 B.n229 585
R845 B.n228 B.n227 585
R846 B.n226 B.n225 585
R847 B.n224 B.n223 585
R848 B.n222 B.n221 585
R849 B.n220 B.n219 585
R850 B.n218 B.n217 585
R851 B.n216 B.n215 585
R852 B.n214 B.n213 585
R853 B.n212 B.n211 585
R854 B.n210 B.n209 585
R855 B.n208 B.n207 585
R856 B.n206 B.n205 585
R857 B.n204 B.n203 585
R858 B.n202 B.n201 585
R859 B.n200 B.n199 585
R860 B.n198 B.n197 585
R861 B.n196 B.n195 585
R862 B.n194 B.n193 585
R863 B.n192 B.n191 585
R864 B.n189 B.n188 585
R865 B.n187 B.n186 585
R866 B.n185 B.n184 585
R867 B.n183 B.n182 585
R868 B.n181 B.n180 585
R869 B.n179 B.n178 585
R870 B.n177 B.n176 585
R871 B.n175 B.n174 585
R872 B.n173 B.n172 585
R873 B.n171 B.n170 585
R874 B.n169 B.n168 585
R875 B.n167 B.n166 585
R876 B.n165 B.n164 585
R877 B.n163 B.n162 585
R878 B.n161 B.n160 585
R879 B.n159 B.n158 585
R880 B.n157 B.n156 585
R881 B.n155 B.n154 585
R882 B.n153 B.n152 585
R883 B.n151 B.n150 585
R884 B.n149 B.n148 585
R885 B.n147 B.n146 585
R886 B.n145 B.n144 585
R887 B.n143 B.n142 585
R888 B.n141 B.n140 585
R889 B.n139 B.n138 585
R890 B.n137 B.n136 585
R891 B.n135 B.n134 585
R892 B.n133 B.n132 585
R893 B.n131 B.n130 585
R894 B.n129 B.n128 585
R895 B.n127 B.n126 585
R896 B.n125 B.n124 585
R897 B.n123 B.n122 585
R898 B.n121 B.n120 585
R899 B.n119 B.n118 585
R900 B.n117 B.n116 585
R901 B.n115 B.n114 585
R902 B.n113 B.n112 585
R903 B.n111 B.n110 585
R904 B.n109 B.n108 585
R905 B.n107 B.n106 585
R906 B.n105 B.n104 585
R907 B.n103 B.n102 585
R908 B.n101 B.n100 585
R909 B.n99 B.n98 585
R910 B.n97 B.n96 585
R911 B.n95 B.n94 585
R912 B.n93 B.n92 585
R913 B.n624 B.n41 585
R914 B.n628 B.n41 585
R915 B.n623 B.n40 585
R916 B.n629 B.n40 585
R917 B.n622 B.n621 585
R918 B.n621 B.n36 585
R919 B.n620 B.n35 585
R920 B.n635 B.n35 585
R921 B.n619 B.n34 585
R922 B.n636 B.n34 585
R923 B.n618 B.n33 585
R924 B.n637 B.n33 585
R925 B.n617 B.n616 585
R926 B.n616 B.n29 585
R927 B.n615 B.n28 585
R928 B.n643 B.n28 585
R929 B.n614 B.n27 585
R930 B.n644 B.n27 585
R931 B.n613 B.n26 585
R932 B.n645 B.n26 585
R933 B.n612 B.n611 585
R934 B.n611 B.n25 585
R935 B.n610 B.n21 585
R936 B.n651 B.n21 585
R937 B.n609 B.n20 585
R938 B.n652 B.n20 585
R939 B.n608 B.n19 585
R940 B.t2 B.n19 585
R941 B.n607 B.n606 585
R942 B.n606 B.n15 585
R943 B.n605 B.n14 585
R944 B.n658 B.n14 585
R945 B.n604 B.n13 585
R946 B.n659 B.n13 585
R947 B.n603 B.n12 585
R948 B.n660 B.n12 585
R949 B.n602 B.n601 585
R950 B.n601 B.n11 585
R951 B.n600 B.n7 585
R952 B.n666 B.n7 585
R953 B.n599 B.n6 585
R954 B.n667 B.n6 585
R955 B.n598 B.n5 585
R956 B.n668 B.n5 585
R957 B.n597 B.n596 585
R958 B.n596 B.n4 585
R959 B.n595 B.n268 585
R960 B.n595 B.n594 585
R961 B.n584 B.n269 585
R962 B.n587 B.n269 585
R963 B.n586 B.n585 585
R964 B.n588 B.n586 585
R965 B.n583 B.n274 585
R966 B.n274 B.n273 585
R967 B.n582 B.n581 585
R968 B.n581 B.n580 585
R969 B.n276 B.n275 585
R970 B.n277 B.n276 585
R971 B.n574 B.n573 585
R972 B.t0 B.n574 585
R973 B.n572 B.n282 585
R974 B.n282 B.n281 585
R975 B.n571 B.n570 585
R976 B.n570 B.n569 585
R977 B.n284 B.n283 585
R978 B.n562 B.n284 585
R979 B.n561 B.n560 585
R980 B.n563 B.n561 585
R981 B.n559 B.n289 585
R982 B.n289 B.n288 585
R983 B.n558 B.n557 585
R984 B.n557 B.n556 585
R985 B.n291 B.n290 585
R986 B.n292 B.n291 585
R987 B.n549 B.n548 585
R988 B.n550 B.n549 585
R989 B.n547 B.n296 585
R990 B.n300 B.n296 585
R991 B.n546 B.n545 585
R992 B.n545 B.n544 585
R993 B.n298 B.n297 585
R994 B.n299 B.n298 585
R995 B.n537 B.n536 585
R996 B.n538 B.n537 585
R997 B.n535 B.n305 585
R998 B.n305 B.n304 585
R999 B.n529 B.n528 585
R1000 B.n527 B.n351 585
R1001 B.n526 B.n350 585
R1002 B.n531 B.n350 585
R1003 B.n525 B.n524 585
R1004 B.n523 B.n522 585
R1005 B.n521 B.n520 585
R1006 B.n519 B.n518 585
R1007 B.n517 B.n516 585
R1008 B.n515 B.n514 585
R1009 B.n513 B.n512 585
R1010 B.n511 B.n510 585
R1011 B.n509 B.n508 585
R1012 B.n507 B.n506 585
R1013 B.n505 B.n504 585
R1014 B.n503 B.n502 585
R1015 B.n501 B.n500 585
R1016 B.n499 B.n498 585
R1017 B.n497 B.n496 585
R1018 B.n495 B.n494 585
R1019 B.n493 B.n492 585
R1020 B.n491 B.n490 585
R1021 B.n489 B.n488 585
R1022 B.n487 B.n486 585
R1023 B.n485 B.n484 585
R1024 B.n483 B.n482 585
R1025 B.n481 B.n480 585
R1026 B.n479 B.n478 585
R1027 B.n477 B.n476 585
R1028 B.n475 B.n474 585
R1029 B.n473 B.n472 585
R1030 B.n471 B.n470 585
R1031 B.n469 B.n468 585
R1032 B.n467 B.n466 585
R1033 B.n465 B.n464 585
R1034 B.n463 B.n462 585
R1035 B.n461 B.n460 585
R1036 B.n459 B.n458 585
R1037 B.n457 B.n456 585
R1038 B.n455 B.n454 585
R1039 B.n453 B.n452 585
R1040 B.n450 B.n449 585
R1041 B.n448 B.n447 585
R1042 B.n446 B.n445 585
R1043 B.n444 B.n443 585
R1044 B.n442 B.n441 585
R1045 B.n440 B.n439 585
R1046 B.n438 B.n437 585
R1047 B.n436 B.n435 585
R1048 B.n434 B.n433 585
R1049 B.n432 B.n431 585
R1050 B.n430 B.n429 585
R1051 B.n428 B.n427 585
R1052 B.n426 B.n425 585
R1053 B.n424 B.n423 585
R1054 B.n422 B.n421 585
R1055 B.n420 B.n419 585
R1056 B.n418 B.n417 585
R1057 B.n416 B.n415 585
R1058 B.n414 B.n413 585
R1059 B.n412 B.n411 585
R1060 B.n410 B.n409 585
R1061 B.n408 B.n407 585
R1062 B.n406 B.n405 585
R1063 B.n404 B.n403 585
R1064 B.n402 B.n401 585
R1065 B.n400 B.n399 585
R1066 B.n398 B.n397 585
R1067 B.n396 B.n395 585
R1068 B.n394 B.n393 585
R1069 B.n392 B.n391 585
R1070 B.n390 B.n389 585
R1071 B.n388 B.n387 585
R1072 B.n386 B.n385 585
R1073 B.n384 B.n383 585
R1074 B.n382 B.n381 585
R1075 B.n380 B.n379 585
R1076 B.n378 B.n377 585
R1077 B.n376 B.n375 585
R1078 B.n374 B.n373 585
R1079 B.n372 B.n371 585
R1080 B.n370 B.n369 585
R1081 B.n368 B.n367 585
R1082 B.n366 B.n365 585
R1083 B.n364 B.n363 585
R1084 B.n362 B.n361 585
R1085 B.n360 B.n359 585
R1086 B.n358 B.n357 585
R1087 B.n307 B.n306 585
R1088 B.n534 B.n533 585
R1089 B.n303 B.n302 585
R1090 B.n304 B.n303 585
R1091 B.n540 B.n539 585
R1092 B.n539 B.n538 585
R1093 B.n541 B.n301 585
R1094 B.n301 B.n299 585
R1095 B.n543 B.n542 585
R1096 B.n544 B.n543 585
R1097 B.n295 B.n294 585
R1098 B.n300 B.n295 585
R1099 B.n552 B.n551 585
R1100 B.n551 B.n550 585
R1101 B.n553 B.n293 585
R1102 B.n293 B.n292 585
R1103 B.n555 B.n554 585
R1104 B.n556 B.n555 585
R1105 B.n287 B.n286 585
R1106 B.n288 B.n287 585
R1107 B.n565 B.n564 585
R1108 B.n564 B.n563 585
R1109 B.n566 B.n285 585
R1110 B.n562 B.n285 585
R1111 B.n568 B.n567 585
R1112 B.n569 B.n568 585
R1113 B.n280 B.n279 585
R1114 B.n281 B.n280 585
R1115 B.n576 B.n575 585
R1116 B.n575 B.t0 585
R1117 B.n577 B.n278 585
R1118 B.n278 B.n277 585
R1119 B.n579 B.n578 585
R1120 B.n580 B.n579 585
R1121 B.n272 B.n271 585
R1122 B.n273 B.n272 585
R1123 B.n590 B.n589 585
R1124 B.n589 B.n588 585
R1125 B.n591 B.n270 585
R1126 B.n587 B.n270 585
R1127 B.n593 B.n592 585
R1128 B.n594 B.n593 585
R1129 B.n2 B.n0 585
R1130 B.n4 B.n2 585
R1131 B.n3 B.n1 585
R1132 B.n667 B.n3 585
R1133 B.n665 B.n664 585
R1134 B.n666 B.n665 585
R1135 B.n663 B.n8 585
R1136 B.n11 B.n8 585
R1137 B.n662 B.n661 585
R1138 B.n661 B.n660 585
R1139 B.n10 B.n9 585
R1140 B.n659 B.n10 585
R1141 B.n657 B.n656 585
R1142 B.n658 B.n657 585
R1143 B.n655 B.n16 585
R1144 B.n16 B.n15 585
R1145 B.n654 B.n653 585
R1146 B.n653 B.t2 585
R1147 B.n18 B.n17 585
R1148 B.n652 B.n18 585
R1149 B.n650 B.n649 585
R1150 B.n651 B.n650 585
R1151 B.n648 B.n22 585
R1152 B.n25 B.n22 585
R1153 B.n647 B.n646 585
R1154 B.n646 B.n645 585
R1155 B.n24 B.n23 585
R1156 B.n644 B.n24 585
R1157 B.n642 B.n641 585
R1158 B.n643 B.n642 585
R1159 B.n640 B.n30 585
R1160 B.n30 B.n29 585
R1161 B.n639 B.n638 585
R1162 B.n638 B.n637 585
R1163 B.n32 B.n31 585
R1164 B.n636 B.n32 585
R1165 B.n634 B.n633 585
R1166 B.n635 B.n634 585
R1167 B.n632 B.n37 585
R1168 B.n37 B.n36 585
R1169 B.n631 B.n630 585
R1170 B.n630 B.n629 585
R1171 B.n39 B.n38 585
R1172 B.n628 B.n39 585
R1173 B.n670 B.n669 585
R1174 B.n669 B.n668 585
R1175 B.n529 B.n303 516.524
R1176 B.n92 B.n39 516.524
R1177 B.n533 B.n305 516.524
R1178 B.n626 B.n41 516.524
R1179 B.n354 B.t10 289.108
R1180 B.n87 B.t13 289.108
R1181 B.n352 B.t17 289.108
R1182 B.n89 B.t19 289.108
R1183 B.n355 B.t9 272.236
R1184 B.n88 B.t14 272.236
R1185 B.n353 B.t16 272.236
R1186 B.n90 B.t20 272.236
R1187 B.n627 B.n85 256.663
R1188 B.n627 B.n84 256.663
R1189 B.n627 B.n83 256.663
R1190 B.n627 B.n82 256.663
R1191 B.n627 B.n81 256.663
R1192 B.n627 B.n80 256.663
R1193 B.n627 B.n79 256.663
R1194 B.n627 B.n78 256.663
R1195 B.n627 B.n77 256.663
R1196 B.n627 B.n76 256.663
R1197 B.n627 B.n75 256.663
R1198 B.n627 B.n74 256.663
R1199 B.n627 B.n73 256.663
R1200 B.n627 B.n72 256.663
R1201 B.n627 B.n71 256.663
R1202 B.n627 B.n70 256.663
R1203 B.n627 B.n69 256.663
R1204 B.n627 B.n68 256.663
R1205 B.n627 B.n67 256.663
R1206 B.n627 B.n66 256.663
R1207 B.n627 B.n65 256.663
R1208 B.n627 B.n64 256.663
R1209 B.n627 B.n63 256.663
R1210 B.n627 B.n62 256.663
R1211 B.n627 B.n61 256.663
R1212 B.n627 B.n60 256.663
R1213 B.n627 B.n59 256.663
R1214 B.n627 B.n58 256.663
R1215 B.n627 B.n57 256.663
R1216 B.n627 B.n56 256.663
R1217 B.n627 B.n55 256.663
R1218 B.n627 B.n54 256.663
R1219 B.n627 B.n53 256.663
R1220 B.n627 B.n52 256.663
R1221 B.n627 B.n51 256.663
R1222 B.n627 B.n50 256.663
R1223 B.n627 B.n49 256.663
R1224 B.n627 B.n48 256.663
R1225 B.n627 B.n47 256.663
R1226 B.n627 B.n46 256.663
R1227 B.n627 B.n45 256.663
R1228 B.n627 B.n44 256.663
R1229 B.n627 B.n43 256.663
R1230 B.n627 B.n42 256.663
R1231 B.n531 B.n530 256.663
R1232 B.n531 B.n308 256.663
R1233 B.n531 B.n309 256.663
R1234 B.n531 B.n310 256.663
R1235 B.n531 B.n311 256.663
R1236 B.n531 B.n312 256.663
R1237 B.n531 B.n313 256.663
R1238 B.n531 B.n314 256.663
R1239 B.n531 B.n315 256.663
R1240 B.n531 B.n316 256.663
R1241 B.n531 B.n317 256.663
R1242 B.n531 B.n318 256.663
R1243 B.n531 B.n319 256.663
R1244 B.n531 B.n320 256.663
R1245 B.n531 B.n321 256.663
R1246 B.n531 B.n322 256.663
R1247 B.n531 B.n323 256.663
R1248 B.n531 B.n324 256.663
R1249 B.n531 B.n325 256.663
R1250 B.n531 B.n326 256.663
R1251 B.n531 B.n327 256.663
R1252 B.n531 B.n328 256.663
R1253 B.n531 B.n329 256.663
R1254 B.n531 B.n330 256.663
R1255 B.n531 B.n331 256.663
R1256 B.n531 B.n332 256.663
R1257 B.n531 B.n333 256.663
R1258 B.n531 B.n334 256.663
R1259 B.n531 B.n335 256.663
R1260 B.n531 B.n336 256.663
R1261 B.n531 B.n337 256.663
R1262 B.n531 B.n338 256.663
R1263 B.n531 B.n339 256.663
R1264 B.n531 B.n340 256.663
R1265 B.n531 B.n341 256.663
R1266 B.n531 B.n342 256.663
R1267 B.n531 B.n343 256.663
R1268 B.n531 B.n344 256.663
R1269 B.n531 B.n345 256.663
R1270 B.n531 B.n346 256.663
R1271 B.n531 B.n347 256.663
R1272 B.n531 B.n348 256.663
R1273 B.n531 B.n349 256.663
R1274 B.n532 B.n531 256.663
R1275 B.n539 B.n303 163.367
R1276 B.n539 B.n301 163.367
R1277 B.n543 B.n301 163.367
R1278 B.n543 B.n295 163.367
R1279 B.n551 B.n295 163.367
R1280 B.n551 B.n293 163.367
R1281 B.n555 B.n293 163.367
R1282 B.n555 B.n287 163.367
R1283 B.n564 B.n287 163.367
R1284 B.n564 B.n285 163.367
R1285 B.n568 B.n285 163.367
R1286 B.n568 B.n280 163.367
R1287 B.n575 B.n280 163.367
R1288 B.n575 B.n278 163.367
R1289 B.n579 B.n278 163.367
R1290 B.n579 B.n272 163.367
R1291 B.n589 B.n272 163.367
R1292 B.n589 B.n270 163.367
R1293 B.n593 B.n270 163.367
R1294 B.n593 B.n2 163.367
R1295 B.n669 B.n2 163.367
R1296 B.n669 B.n3 163.367
R1297 B.n665 B.n3 163.367
R1298 B.n665 B.n8 163.367
R1299 B.n661 B.n8 163.367
R1300 B.n661 B.n10 163.367
R1301 B.n657 B.n10 163.367
R1302 B.n657 B.n16 163.367
R1303 B.n653 B.n16 163.367
R1304 B.n653 B.n18 163.367
R1305 B.n650 B.n18 163.367
R1306 B.n650 B.n22 163.367
R1307 B.n646 B.n22 163.367
R1308 B.n646 B.n24 163.367
R1309 B.n642 B.n24 163.367
R1310 B.n642 B.n30 163.367
R1311 B.n638 B.n30 163.367
R1312 B.n638 B.n32 163.367
R1313 B.n634 B.n32 163.367
R1314 B.n634 B.n37 163.367
R1315 B.n630 B.n37 163.367
R1316 B.n630 B.n39 163.367
R1317 B.n351 B.n350 163.367
R1318 B.n524 B.n350 163.367
R1319 B.n522 B.n521 163.367
R1320 B.n518 B.n517 163.367
R1321 B.n514 B.n513 163.367
R1322 B.n510 B.n509 163.367
R1323 B.n506 B.n505 163.367
R1324 B.n502 B.n501 163.367
R1325 B.n498 B.n497 163.367
R1326 B.n494 B.n493 163.367
R1327 B.n490 B.n489 163.367
R1328 B.n486 B.n485 163.367
R1329 B.n482 B.n481 163.367
R1330 B.n478 B.n477 163.367
R1331 B.n474 B.n473 163.367
R1332 B.n470 B.n469 163.367
R1333 B.n466 B.n465 163.367
R1334 B.n462 B.n461 163.367
R1335 B.n458 B.n457 163.367
R1336 B.n454 B.n453 163.367
R1337 B.n449 B.n448 163.367
R1338 B.n445 B.n444 163.367
R1339 B.n441 B.n440 163.367
R1340 B.n437 B.n436 163.367
R1341 B.n433 B.n432 163.367
R1342 B.n429 B.n428 163.367
R1343 B.n425 B.n424 163.367
R1344 B.n421 B.n420 163.367
R1345 B.n417 B.n416 163.367
R1346 B.n413 B.n412 163.367
R1347 B.n409 B.n408 163.367
R1348 B.n405 B.n404 163.367
R1349 B.n401 B.n400 163.367
R1350 B.n397 B.n396 163.367
R1351 B.n393 B.n392 163.367
R1352 B.n389 B.n388 163.367
R1353 B.n385 B.n384 163.367
R1354 B.n381 B.n380 163.367
R1355 B.n377 B.n376 163.367
R1356 B.n373 B.n372 163.367
R1357 B.n369 B.n368 163.367
R1358 B.n365 B.n364 163.367
R1359 B.n361 B.n360 163.367
R1360 B.n357 B.n307 163.367
R1361 B.n537 B.n305 163.367
R1362 B.n537 B.n298 163.367
R1363 B.n545 B.n298 163.367
R1364 B.n545 B.n296 163.367
R1365 B.n549 B.n296 163.367
R1366 B.n549 B.n291 163.367
R1367 B.n557 B.n291 163.367
R1368 B.n557 B.n289 163.367
R1369 B.n561 B.n289 163.367
R1370 B.n561 B.n284 163.367
R1371 B.n570 B.n284 163.367
R1372 B.n570 B.n282 163.367
R1373 B.n574 B.n282 163.367
R1374 B.n574 B.n276 163.367
R1375 B.n581 B.n276 163.367
R1376 B.n581 B.n274 163.367
R1377 B.n586 B.n274 163.367
R1378 B.n586 B.n269 163.367
R1379 B.n595 B.n269 163.367
R1380 B.n596 B.n595 163.367
R1381 B.n596 B.n5 163.367
R1382 B.n6 B.n5 163.367
R1383 B.n7 B.n6 163.367
R1384 B.n601 B.n7 163.367
R1385 B.n601 B.n12 163.367
R1386 B.n13 B.n12 163.367
R1387 B.n14 B.n13 163.367
R1388 B.n606 B.n14 163.367
R1389 B.n606 B.n19 163.367
R1390 B.n20 B.n19 163.367
R1391 B.n21 B.n20 163.367
R1392 B.n611 B.n21 163.367
R1393 B.n611 B.n26 163.367
R1394 B.n27 B.n26 163.367
R1395 B.n28 B.n27 163.367
R1396 B.n616 B.n28 163.367
R1397 B.n616 B.n33 163.367
R1398 B.n34 B.n33 163.367
R1399 B.n35 B.n34 163.367
R1400 B.n621 B.n35 163.367
R1401 B.n621 B.n40 163.367
R1402 B.n41 B.n40 163.367
R1403 B.n96 B.n95 163.367
R1404 B.n100 B.n99 163.367
R1405 B.n104 B.n103 163.367
R1406 B.n108 B.n107 163.367
R1407 B.n112 B.n111 163.367
R1408 B.n116 B.n115 163.367
R1409 B.n120 B.n119 163.367
R1410 B.n124 B.n123 163.367
R1411 B.n128 B.n127 163.367
R1412 B.n132 B.n131 163.367
R1413 B.n136 B.n135 163.367
R1414 B.n140 B.n139 163.367
R1415 B.n144 B.n143 163.367
R1416 B.n148 B.n147 163.367
R1417 B.n152 B.n151 163.367
R1418 B.n156 B.n155 163.367
R1419 B.n160 B.n159 163.367
R1420 B.n164 B.n163 163.367
R1421 B.n168 B.n167 163.367
R1422 B.n172 B.n171 163.367
R1423 B.n176 B.n175 163.367
R1424 B.n180 B.n179 163.367
R1425 B.n184 B.n183 163.367
R1426 B.n188 B.n187 163.367
R1427 B.n193 B.n192 163.367
R1428 B.n197 B.n196 163.367
R1429 B.n201 B.n200 163.367
R1430 B.n205 B.n204 163.367
R1431 B.n209 B.n208 163.367
R1432 B.n213 B.n212 163.367
R1433 B.n217 B.n216 163.367
R1434 B.n221 B.n220 163.367
R1435 B.n225 B.n224 163.367
R1436 B.n229 B.n228 163.367
R1437 B.n233 B.n232 163.367
R1438 B.n237 B.n236 163.367
R1439 B.n241 B.n240 163.367
R1440 B.n245 B.n244 163.367
R1441 B.n249 B.n248 163.367
R1442 B.n253 B.n252 163.367
R1443 B.n257 B.n256 163.367
R1444 B.n261 B.n260 163.367
R1445 B.n265 B.n264 163.367
R1446 B.n626 B.n86 163.367
R1447 B.n531 B.n304 77.0894
R1448 B.n628 B.n627 77.0894
R1449 B.n530 B.n529 71.676
R1450 B.n524 B.n308 71.676
R1451 B.n521 B.n309 71.676
R1452 B.n517 B.n310 71.676
R1453 B.n513 B.n311 71.676
R1454 B.n509 B.n312 71.676
R1455 B.n505 B.n313 71.676
R1456 B.n501 B.n314 71.676
R1457 B.n497 B.n315 71.676
R1458 B.n493 B.n316 71.676
R1459 B.n489 B.n317 71.676
R1460 B.n485 B.n318 71.676
R1461 B.n481 B.n319 71.676
R1462 B.n477 B.n320 71.676
R1463 B.n473 B.n321 71.676
R1464 B.n469 B.n322 71.676
R1465 B.n465 B.n323 71.676
R1466 B.n461 B.n324 71.676
R1467 B.n457 B.n325 71.676
R1468 B.n453 B.n326 71.676
R1469 B.n448 B.n327 71.676
R1470 B.n444 B.n328 71.676
R1471 B.n440 B.n329 71.676
R1472 B.n436 B.n330 71.676
R1473 B.n432 B.n331 71.676
R1474 B.n428 B.n332 71.676
R1475 B.n424 B.n333 71.676
R1476 B.n420 B.n334 71.676
R1477 B.n416 B.n335 71.676
R1478 B.n412 B.n336 71.676
R1479 B.n408 B.n337 71.676
R1480 B.n404 B.n338 71.676
R1481 B.n400 B.n339 71.676
R1482 B.n396 B.n340 71.676
R1483 B.n392 B.n341 71.676
R1484 B.n388 B.n342 71.676
R1485 B.n384 B.n343 71.676
R1486 B.n380 B.n344 71.676
R1487 B.n376 B.n345 71.676
R1488 B.n372 B.n346 71.676
R1489 B.n368 B.n347 71.676
R1490 B.n364 B.n348 71.676
R1491 B.n360 B.n349 71.676
R1492 B.n532 B.n307 71.676
R1493 B.n92 B.n42 71.676
R1494 B.n96 B.n43 71.676
R1495 B.n100 B.n44 71.676
R1496 B.n104 B.n45 71.676
R1497 B.n108 B.n46 71.676
R1498 B.n112 B.n47 71.676
R1499 B.n116 B.n48 71.676
R1500 B.n120 B.n49 71.676
R1501 B.n124 B.n50 71.676
R1502 B.n128 B.n51 71.676
R1503 B.n132 B.n52 71.676
R1504 B.n136 B.n53 71.676
R1505 B.n140 B.n54 71.676
R1506 B.n144 B.n55 71.676
R1507 B.n148 B.n56 71.676
R1508 B.n152 B.n57 71.676
R1509 B.n156 B.n58 71.676
R1510 B.n160 B.n59 71.676
R1511 B.n164 B.n60 71.676
R1512 B.n168 B.n61 71.676
R1513 B.n172 B.n62 71.676
R1514 B.n176 B.n63 71.676
R1515 B.n180 B.n64 71.676
R1516 B.n184 B.n65 71.676
R1517 B.n188 B.n66 71.676
R1518 B.n193 B.n67 71.676
R1519 B.n197 B.n68 71.676
R1520 B.n201 B.n69 71.676
R1521 B.n205 B.n70 71.676
R1522 B.n209 B.n71 71.676
R1523 B.n213 B.n72 71.676
R1524 B.n217 B.n73 71.676
R1525 B.n221 B.n74 71.676
R1526 B.n225 B.n75 71.676
R1527 B.n229 B.n76 71.676
R1528 B.n233 B.n77 71.676
R1529 B.n237 B.n78 71.676
R1530 B.n241 B.n79 71.676
R1531 B.n245 B.n80 71.676
R1532 B.n249 B.n81 71.676
R1533 B.n253 B.n82 71.676
R1534 B.n257 B.n83 71.676
R1535 B.n261 B.n84 71.676
R1536 B.n265 B.n85 71.676
R1537 B.n86 B.n85 71.676
R1538 B.n264 B.n84 71.676
R1539 B.n260 B.n83 71.676
R1540 B.n256 B.n82 71.676
R1541 B.n252 B.n81 71.676
R1542 B.n248 B.n80 71.676
R1543 B.n244 B.n79 71.676
R1544 B.n240 B.n78 71.676
R1545 B.n236 B.n77 71.676
R1546 B.n232 B.n76 71.676
R1547 B.n228 B.n75 71.676
R1548 B.n224 B.n74 71.676
R1549 B.n220 B.n73 71.676
R1550 B.n216 B.n72 71.676
R1551 B.n212 B.n71 71.676
R1552 B.n208 B.n70 71.676
R1553 B.n204 B.n69 71.676
R1554 B.n200 B.n68 71.676
R1555 B.n196 B.n67 71.676
R1556 B.n192 B.n66 71.676
R1557 B.n187 B.n65 71.676
R1558 B.n183 B.n64 71.676
R1559 B.n179 B.n63 71.676
R1560 B.n175 B.n62 71.676
R1561 B.n171 B.n61 71.676
R1562 B.n167 B.n60 71.676
R1563 B.n163 B.n59 71.676
R1564 B.n159 B.n58 71.676
R1565 B.n155 B.n57 71.676
R1566 B.n151 B.n56 71.676
R1567 B.n147 B.n55 71.676
R1568 B.n143 B.n54 71.676
R1569 B.n139 B.n53 71.676
R1570 B.n135 B.n52 71.676
R1571 B.n131 B.n51 71.676
R1572 B.n127 B.n50 71.676
R1573 B.n123 B.n49 71.676
R1574 B.n119 B.n48 71.676
R1575 B.n115 B.n47 71.676
R1576 B.n111 B.n46 71.676
R1577 B.n107 B.n45 71.676
R1578 B.n103 B.n44 71.676
R1579 B.n99 B.n43 71.676
R1580 B.n95 B.n42 71.676
R1581 B.n530 B.n351 71.676
R1582 B.n522 B.n308 71.676
R1583 B.n518 B.n309 71.676
R1584 B.n514 B.n310 71.676
R1585 B.n510 B.n311 71.676
R1586 B.n506 B.n312 71.676
R1587 B.n502 B.n313 71.676
R1588 B.n498 B.n314 71.676
R1589 B.n494 B.n315 71.676
R1590 B.n490 B.n316 71.676
R1591 B.n486 B.n317 71.676
R1592 B.n482 B.n318 71.676
R1593 B.n478 B.n319 71.676
R1594 B.n474 B.n320 71.676
R1595 B.n470 B.n321 71.676
R1596 B.n466 B.n322 71.676
R1597 B.n462 B.n323 71.676
R1598 B.n458 B.n324 71.676
R1599 B.n454 B.n325 71.676
R1600 B.n449 B.n326 71.676
R1601 B.n445 B.n327 71.676
R1602 B.n441 B.n328 71.676
R1603 B.n437 B.n329 71.676
R1604 B.n433 B.n330 71.676
R1605 B.n429 B.n331 71.676
R1606 B.n425 B.n332 71.676
R1607 B.n421 B.n333 71.676
R1608 B.n417 B.n334 71.676
R1609 B.n413 B.n335 71.676
R1610 B.n409 B.n336 71.676
R1611 B.n405 B.n337 71.676
R1612 B.n401 B.n338 71.676
R1613 B.n397 B.n339 71.676
R1614 B.n393 B.n340 71.676
R1615 B.n389 B.n341 71.676
R1616 B.n385 B.n342 71.676
R1617 B.n381 B.n343 71.676
R1618 B.n377 B.n344 71.676
R1619 B.n373 B.n345 71.676
R1620 B.n369 B.n346 71.676
R1621 B.n365 B.n347 71.676
R1622 B.n361 B.n348 71.676
R1623 B.n357 B.n349 71.676
R1624 B.n533 B.n532 71.676
R1625 B.n356 B.n355 59.5399
R1626 B.n451 B.n353 59.5399
R1627 B.n91 B.n90 59.5399
R1628 B.n190 B.n88 59.5399
R1629 B.n538 B.n304 44.8043
R1630 B.n538 B.n299 44.8043
R1631 B.n544 B.n299 44.8043
R1632 B.n544 B.n300 44.8043
R1633 B.n550 B.n292 44.8043
R1634 B.n556 B.n292 44.8043
R1635 B.n556 B.n288 44.8043
R1636 B.n563 B.n288 44.8043
R1637 B.n563 B.n562 44.8043
R1638 B.n569 B.n281 44.8043
R1639 B.t0 B.n281 44.8043
R1640 B.t0 B.n277 44.8043
R1641 B.n580 B.n277 44.8043
R1642 B.n588 B.n273 44.8043
R1643 B.n588 B.n587 44.8043
R1644 B.n594 B.n4 44.8043
R1645 B.n668 B.n4 44.8043
R1646 B.n668 B.n667 44.8043
R1647 B.n667 B.n666 44.8043
R1648 B.n660 B.n11 44.8043
R1649 B.n660 B.n659 44.8043
R1650 B.n658 B.n15 44.8043
R1651 B.t2 B.n15 44.8043
R1652 B.t2 B.n652 44.8043
R1653 B.n652 B.n651 44.8043
R1654 B.n645 B.n25 44.8043
R1655 B.n645 B.n644 44.8043
R1656 B.n644 B.n643 44.8043
R1657 B.n643 B.n29 44.8043
R1658 B.n637 B.n29 44.8043
R1659 B.n636 B.n635 44.8043
R1660 B.n635 B.n36 44.8043
R1661 B.n629 B.n36 44.8043
R1662 B.n629 B.n628 44.8043
R1663 B.n594 B.t1 39.5333
R1664 B.n666 B.t21 39.5333
R1665 B.n93 B.n38 33.5615
R1666 B.n625 B.n624 33.5615
R1667 B.n535 B.n534 33.5615
R1668 B.n528 B.n302 33.5615
R1669 B.n300 B.t8 30.309
R1670 B.t12 B.n636 30.309
R1671 B.n569 B.t3 25.0379
R1672 B.n580 B.t4 25.0379
R1673 B.t6 B.n658 25.0379
R1674 B.n651 B.t5 25.0379
R1675 B.n562 B.t3 19.7669
R1676 B.t4 B.n273 19.7669
R1677 B.n659 B.t6 19.7669
R1678 B.n25 B.t5 19.7669
R1679 B B.n670 18.0485
R1680 B.n355 B.n354 16.8732
R1681 B.n353 B.n352 16.8732
R1682 B.n90 B.n89 16.8732
R1683 B.n88 B.n87 16.8732
R1684 B.n550 B.t8 14.4959
R1685 B.n637 B.t12 14.4959
R1686 B.n94 B.n93 10.6151
R1687 B.n97 B.n94 10.6151
R1688 B.n98 B.n97 10.6151
R1689 B.n101 B.n98 10.6151
R1690 B.n102 B.n101 10.6151
R1691 B.n105 B.n102 10.6151
R1692 B.n106 B.n105 10.6151
R1693 B.n109 B.n106 10.6151
R1694 B.n110 B.n109 10.6151
R1695 B.n113 B.n110 10.6151
R1696 B.n114 B.n113 10.6151
R1697 B.n117 B.n114 10.6151
R1698 B.n118 B.n117 10.6151
R1699 B.n121 B.n118 10.6151
R1700 B.n122 B.n121 10.6151
R1701 B.n125 B.n122 10.6151
R1702 B.n126 B.n125 10.6151
R1703 B.n129 B.n126 10.6151
R1704 B.n130 B.n129 10.6151
R1705 B.n133 B.n130 10.6151
R1706 B.n134 B.n133 10.6151
R1707 B.n137 B.n134 10.6151
R1708 B.n138 B.n137 10.6151
R1709 B.n141 B.n138 10.6151
R1710 B.n142 B.n141 10.6151
R1711 B.n145 B.n142 10.6151
R1712 B.n146 B.n145 10.6151
R1713 B.n149 B.n146 10.6151
R1714 B.n150 B.n149 10.6151
R1715 B.n153 B.n150 10.6151
R1716 B.n154 B.n153 10.6151
R1717 B.n157 B.n154 10.6151
R1718 B.n158 B.n157 10.6151
R1719 B.n161 B.n158 10.6151
R1720 B.n162 B.n161 10.6151
R1721 B.n165 B.n162 10.6151
R1722 B.n166 B.n165 10.6151
R1723 B.n169 B.n166 10.6151
R1724 B.n170 B.n169 10.6151
R1725 B.n174 B.n173 10.6151
R1726 B.n177 B.n174 10.6151
R1727 B.n178 B.n177 10.6151
R1728 B.n181 B.n178 10.6151
R1729 B.n182 B.n181 10.6151
R1730 B.n185 B.n182 10.6151
R1731 B.n186 B.n185 10.6151
R1732 B.n189 B.n186 10.6151
R1733 B.n194 B.n191 10.6151
R1734 B.n195 B.n194 10.6151
R1735 B.n198 B.n195 10.6151
R1736 B.n199 B.n198 10.6151
R1737 B.n202 B.n199 10.6151
R1738 B.n203 B.n202 10.6151
R1739 B.n206 B.n203 10.6151
R1740 B.n207 B.n206 10.6151
R1741 B.n210 B.n207 10.6151
R1742 B.n211 B.n210 10.6151
R1743 B.n214 B.n211 10.6151
R1744 B.n215 B.n214 10.6151
R1745 B.n218 B.n215 10.6151
R1746 B.n219 B.n218 10.6151
R1747 B.n222 B.n219 10.6151
R1748 B.n223 B.n222 10.6151
R1749 B.n226 B.n223 10.6151
R1750 B.n227 B.n226 10.6151
R1751 B.n230 B.n227 10.6151
R1752 B.n231 B.n230 10.6151
R1753 B.n234 B.n231 10.6151
R1754 B.n235 B.n234 10.6151
R1755 B.n238 B.n235 10.6151
R1756 B.n239 B.n238 10.6151
R1757 B.n242 B.n239 10.6151
R1758 B.n243 B.n242 10.6151
R1759 B.n246 B.n243 10.6151
R1760 B.n247 B.n246 10.6151
R1761 B.n250 B.n247 10.6151
R1762 B.n251 B.n250 10.6151
R1763 B.n254 B.n251 10.6151
R1764 B.n255 B.n254 10.6151
R1765 B.n258 B.n255 10.6151
R1766 B.n259 B.n258 10.6151
R1767 B.n262 B.n259 10.6151
R1768 B.n263 B.n262 10.6151
R1769 B.n266 B.n263 10.6151
R1770 B.n267 B.n266 10.6151
R1771 B.n625 B.n267 10.6151
R1772 B.n536 B.n535 10.6151
R1773 B.n536 B.n297 10.6151
R1774 B.n546 B.n297 10.6151
R1775 B.n547 B.n546 10.6151
R1776 B.n548 B.n547 10.6151
R1777 B.n548 B.n290 10.6151
R1778 B.n558 B.n290 10.6151
R1779 B.n559 B.n558 10.6151
R1780 B.n560 B.n559 10.6151
R1781 B.n560 B.n283 10.6151
R1782 B.n571 B.n283 10.6151
R1783 B.n572 B.n571 10.6151
R1784 B.n573 B.n572 10.6151
R1785 B.n573 B.n275 10.6151
R1786 B.n582 B.n275 10.6151
R1787 B.n583 B.n582 10.6151
R1788 B.n585 B.n583 10.6151
R1789 B.n585 B.n584 10.6151
R1790 B.n584 B.n268 10.6151
R1791 B.n597 B.n268 10.6151
R1792 B.n598 B.n597 10.6151
R1793 B.n599 B.n598 10.6151
R1794 B.n600 B.n599 10.6151
R1795 B.n602 B.n600 10.6151
R1796 B.n603 B.n602 10.6151
R1797 B.n604 B.n603 10.6151
R1798 B.n605 B.n604 10.6151
R1799 B.n607 B.n605 10.6151
R1800 B.n608 B.n607 10.6151
R1801 B.n609 B.n608 10.6151
R1802 B.n610 B.n609 10.6151
R1803 B.n612 B.n610 10.6151
R1804 B.n613 B.n612 10.6151
R1805 B.n614 B.n613 10.6151
R1806 B.n615 B.n614 10.6151
R1807 B.n617 B.n615 10.6151
R1808 B.n618 B.n617 10.6151
R1809 B.n619 B.n618 10.6151
R1810 B.n620 B.n619 10.6151
R1811 B.n622 B.n620 10.6151
R1812 B.n623 B.n622 10.6151
R1813 B.n624 B.n623 10.6151
R1814 B.n528 B.n527 10.6151
R1815 B.n527 B.n526 10.6151
R1816 B.n526 B.n525 10.6151
R1817 B.n525 B.n523 10.6151
R1818 B.n523 B.n520 10.6151
R1819 B.n520 B.n519 10.6151
R1820 B.n519 B.n516 10.6151
R1821 B.n516 B.n515 10.6151
R1822 B.n515 B.n512 10.6151
R1823 B.n512 B.n511 10.6151
R1824 B.n511 B.n508 10.6151
R1825 B.n508 B.n507 10.6151
R1826 B.n507 B.n504 10.6151
R1827 B.n504 B.n503 10.6151
R1828 B.n503 B.n500 10.6151
R1829 B.n500 B.n499 10.6151
R1830 B.n499 B.n496 10.6151
R1831 B.n496 B.n495 10.6151
R1832 B.n495 B.n492 10.6151
R1833 B.n492 B.n491 10.6151
R1834 B.n491 B.n488 10.6151
R1835 B.n488 B.n487 10.6151
R1836 B.n487 B.n484 10.6151
R1837 B.n484 B.n483 10.6151
R1838 B.n483 B.n480 10.6151
R1839 B.n480 B.n479 10.6151
R1840 B.n479 B.n476 10.6151
R1841 B.n476 B.n475 10.6151
R1842 B.n475 B.n472 10.6151
R1843 B.n472 B.n471 10.6151
R1844 B.n471 B.n468 10.6151
R1845 B.n468 B.n467 10.6151
R1846 B.n467 B.n464 10.6151
R1847 B.n464 B.n463 10.6151
R1848 B.n463 B.n460 10.6151
R1849 B.n460 B.n459 10.6151
R1850 B.n459 B.n456 10.6151
R1851 B.n456 B.n455 10.6151
R1852 B.n455 B.n452 10.6151
R1853 B.n450 B.n447 10.6151
R1854 B.n447 B.n446 10.6151
R1855 B.n446 B.n443 10.6151
R1856 B.n443 B.n442 10.6151
R1857 B.n442 B.n439 10.6151
R1858 B.n439 B.n438 10.6151
R1859 B.n438 B.n435 10.6151
R1860 B.n435 B.n434 10.6151
R1861 B.n431 B.n430 10.6151
R1862 B.n430 B.n427 10.6151
R1863 B.n427 B.n426 10.6151
R1864 B.n426 B.n423 10.6151
R1865 B.n423 B.n422 10.6151
R1866 B.n422 B.n419 10.6151
R1867 B.n419 B.n418 10.6151
R1868 B.n418 B.n415 10.6151
R1869 B.n415 B.n414 10.6151
R1870 B.n414 B.n411 10.6151
R1871 B.n411 B.n410 10.6151
R1872 B.n410 B.n407 10.6151
R1873 B.n407 B.n406 10.6151
R1874 B.n406 B.n403 10.6151
R1875 B.n403 B.n402 10.6151
R1876 B.n402 B.n399 10.6151
R1877 B.n399 B.n398 10.6151
R1878 B.n398 B.n395 10.6151
R1879 B.n395 B.n394 10.6151
R1880 B.n394 B.n391 10.6151
R1881 B.n391 B.n390 10.6151
R1882 B.n390 B.n387 10.6151
R1883 B.n387 B.n386 10.6151
R1884 B.n386 B.n383 10.6151
R1885 B.n383 B.n382 10.6151
R1886 B.n382 B.n379 10.6151
R1887 B.n379 B.n378 10.6151
R1888 B.n378 B.n375 10.6151
R1889 B.n375 B.n374 10.6151
R1890 B.n374 B.n371 10.6151
R1891 B.n371 B.n370 10.6151
R1892 B.n370 B.n367 10.6151
R1893 B.n367 B.n366 10.6151
R1894 B.n366 B.n363 10.6151
R1895 B.n363 B.n362 10.6151
R1896 B.n362 B.n359 10.6151
R1897 B.n359 B.n358 10.6151
R1898 B.n358 B.n306 10.6151
R1899 B.n534 B.n306 10.6151
R1900 B.n540 B.n302 10.6151
R1901 B.n541 B.n540 10.6151
R1902 B.n542 B.n541 10.6151
R1903 B.n542 B.n294 10.6151
R1904 B.n552 B.n294 10.6151
R1905 B.n553 B.n552 10.6151
R1906 B.n554 B.n553 10.6151
R1907 B.n554 B.n286 10.6151
R1908 B.n565 B.n286 10.6151
R1909 B.n566 B.n565 10.6151
R1910 B.n567 B.n566 10.6151
R1911 B.n567 B.n279 10.6151
R1912 B.n576 B.n279 10.6151
R1913 B.n577 B.n576 10.6151
R1914 B.n578 B.n577 10.6151
R1915 B.n578 B.n271 10.6151
R1916 B.n590 B.n271 10.6151
R1917 B.n591 B.n590 10.6151
R1918 B.n592 B.n591 10.6151
R1919 B.n592 B.n0 10.6151
R1920 B.n664 B.n1 10.6151
R1921 B.n664 B.n663 10.6151
R1922 B.n663 B.n662 10.6151
R1923 B.n662 B.n9 10.6151
R1924 B.n656 B.n9 10.6151
R1925 B.n656 B.n655 10.6151
R1926 B.n655 B.n654 10.6151
R1927 B.n654 B.n17 10.6151
R1928 B.n649 B.n17 10.6151
R1929 B.n649 B.n648 10.6151
R1930 B.n648 B.n647 10.6151
R1931 B.n647 B.n23 10.6151
R1932 B.n641 B.n23 10.6151
R1933 B.n641 B.n640 10.6151
R1934 B.n640 B.n639 10.6151
R1935 B.n639 B.n31 10.6151
R1936 B.n633 B.n31 10.6151
R1937 B.n633 B.n632 10.6151
R1938 B.n632 B.n631 10.6151
R1939 B.n631 B.n38 10.6151
R1940 B.n173 B.n91 6.5566
R1941 B.n190 B.n189 6.5566
R1942 B.n451 B.n450 6.5566
R1943 B.n434 B.n356 6.5566
R1944 B.n587 B.t1 5.27154
R1945 B.n11 B.t21 5.27154
R1946 B.n170 B.n91 4.05904
R1947 B.n191 B.n190 4.05904
R1948 B.n452 B.n451 4.05904
R1949 B.n431 B.n356 4.05904
R1950 B.n670 B.n0 2.81026
R1951 B.n670 B.n1 2.81026
R1952 VN.n2 VN.t1 607.811
R1953 VN.n10 VN.t6 607.811
R1954 VN.n1 VN.t3 582.418
R1955 VN.n4 VN.t2 582.418
R1956 VN.n6 VN.t4 582.418
R1957 VN.n9 VN.t5 582.418
R1958 VN.n12 VN.t0 582.418
R1959 VN.n14 VN.t7 582.418
R1960 VN.n7 VN.n6 161.3
R1961 VN.n15 VN.n14 161.3
R1962 VN.n13 VN.n8 161.3
R1963 VN.n12 VN.n11 161.3
R1964 VN.n5 VN.n0 161.3
R1965 VN.n4 VN.n3 161.3
R1966 VN.n4 VN.n1 48.2005
R1967 VN.n12 VN.n9 48.2005
R1968 VN.n11 VN.n10 45.0031
R1969 VN.n3 VN.n2 45.0031
R1970 VN.n6 VN.n5 41.6278
R1971 VN.n14 VN.n13 41.6278
R1972 VN VN.n15 41.1539
R1973 VN.n2 VN.n1 15.6319
R1974 VN.n10 VN.n9 15.6319
R1975 VN.n5 VN.n4 6.57323
R1976 VN.n13 VN.n12 6.57323
R1977 VN.n15 VN.n8 0.189894
R1978 VN.n11 VN.n8 0.189894
R1979 VN.n3 VN.n0 0.189894
R1980 VN.n7 VN.n0 0.189894
R1981 VN VN.n7 0.0516364
R1982 VDD2.n2 VDD2.n1 62.7973
R1983 VDD2.n2 VDD2.n0 62.7973
R1984 VDD2 VDD2.n5 62.7944
R1985 VDD2.n4 VDD2.n3 62.4778
R1986 VDD2.n4 VDD2.n2 36.9351
R1987 VDD2.n5 VDD2.t2 1.7343
R1988 VDD2.n5 VDD2.t1 1.7343
R1989 VDD2.n3 VDD2.t0 1.7343
R1990 VDD2.n3 VDD2.t7 1.7343
R1991 VDD2.n1 VDD2.t5 1.7343
R1992 VDD2.n1 VDD2.t3 1.7343
R1993 VDD2.n0 VDD2.t6 1.7343
R1994 VDD2.n0 VDD2.t4 1.7343
R1995 VDD2 VDD2.n4 0.43369
C0 VDD2 VDD1 0.746651f
C1 VDD1 VP 4.7219f
C2 VDD2 VTAIL 12.0108f
C3 VN VDD1 0.148197f
C4 VTAIL VP 4.29486f
C5 VN VTAIL 4.28076f
C6 VDD2 VP 0.300659f
C7 VN VDD2 4.56979f
C8 VN VP 5.03623f
C9 VTAIL VDD1 11.970201f
C10 VDD2 B 3.300079f
C11 VDD1 B 3.518007f
C12 VTAIL B 8.445229f
C13 VN B 7.987f
C14 VP B 5.966741f
C15 VDD2.t6 B 0.259701f
C16 VDD2.t4 B 0.259701f
C17 VDD2.n0 B 2.30912f
C18 VDD2.t5 B 0.259701f
C19 VDD2.t3 B 0.259701f
C20 VDD2.n1 B 2.30912f
C21 VDD2.n2 B 2.35199f
C22 VDD2.t0 B 0.259701f
C23 VDD2.t7 B 0.259701f
C24 VDD2.n3 B 2.30735f
C25 VDD2.n4 B 2.52043f
C26 VDD2.t2 B 0.259701f
C27 VDD2.t1 B 0.259701f
C28 VDD2.n5 B 2.3091f
C29 VN.n0 B 0.047954f
C30 VN.t3 B 0.844003f
C31 VN.n1 B 0.351883f
C32 VN.t1 B 0.858296f
C33 VN.n2 B 0.330719f
C34 VN.n3 B 0.195304f
C35 VN.t2 B 0.844003f
C36 VN.n4 B 0.343863f
C37 VN.n5 B 0.010882f
C38 VN.t4 B 0.844003f
C39 VN.n6 B 0.341202f
C40 VN.n7 B 0.037163f
C41 VN.n8 B 0.047954f
C42 VN.t5 B 0.844003f
C43 VN.n9 B 0.351883f
C44 VN.t0 B 0.844003f
C45 VN.t6 B 0.858296f
C46 VN.n10 B 0.330719f
C47 VN.n11 B 0.195304f
C48 VN.n12 B 0.343863f
C49 VN.n13 B 0.010882f
C50 VN.t7 B 0.844003f
C51 VN.n14 B 0.341202f
C52 VN.n15 B 1.91452f
C53 VTAIL.t6 B 0.189883f
C54 VTAIL.t2 B 0.189883f
C55 VTAIL.n0 B 1.6254f
C56 VTAIL.n1 B 0.261102f
C57 VTAIL.n2 B 0.029291f
C58 VTAIL.n3 B 0.021041f
C59 VTAIL.n4 B 0.011307f
C60 VTAIL.n5 B 0.026725f
C61 VTAIL.n6 B 0.011972f
C62 VTAIL.n7 B 0.021041f
C63 VTAIL.n8 B 0.011307f
C64 VTAIL.n9 B 0.026725f
C65 VTAIL.n10 B 0.011639f
C66 VTAIL.n11 B 0.021041f
C67 VTAIL.n12 B 0.011972f
C68 VTAIL.n13 B 0.026725f
C69 VTAIL.n14 B 0.011972f
C70 VTAIL.n15 B 0.021041f
C71 VTAIL.n16 B 0.011307f
C72 VTAIL.n17 B 0.026725f
C73 VTAIL.n18 B 0.011972f
C74 VTAIL.n19 B 1.0072f
C75 VTAIL.n20 B 0.011307f
C76 VTAIL.t15 B 0.04507f
C77 VTAIL.n21 B 0.147019f
C78 VTAIL.n22 B 0.018892f
C79 VTAIL.n23 B 0.020043f
C80 VTAIL.n24 B 0.026725f
C81 VTAIL.n25 B 0.011972f
C82 VTAIL.n26 B 0.011307f
C83 VTAIL.n27 B 0.021041f
C84 VTAIL.n28 B 0.021041f
C85 VTAIL.n29 B 0.011307f
C86 VTAIL.n30 B 0.011972f
C87 VTAIL.n31 B 0.026725f
C88 VTAIL.n32 B 0.026725f
C89 VTAIL.n33 B 0.011972f
C90 VTAIL.n34 B 0.011307f
C91 VTAIL.n35 B 0.021041f
C92 VTAIL.n36 B 0.021041f
C93 VTAIL.n37 B 0.011307f
C94 VTAIL.n38 B 0.011307f
C95 VTAIL.n39 B 0.011972f
C96 VTAIL.n40 B 0.026725f
C97 VTAIL.n41 B 0.026725f
C98 VTAIL.n42 B 0.026725f
C99 VTAIL.n43 B 0.011639f
C100 VTAIL.n44 B 0.011307f
C101 VTAIL.n45 B 0.021041f
C102 VTAIL.n46 B 0.021041f
C103 VTAIL.n47 B 0.011307f
C104 VTAIL.n48 B 0.011972f
C105 VTAIL.n49 B 0.026725f
C106 VTAIL.n50 B 0.026725f
C107 VTAIL.n51 B 0.011972f
C108 VTAIL.n52 B 0.011307f
C109 VTAIL.n53 B 0.021041f
C110 VTAIL.n54 B 0.021041f
C111 VTAIL.n55 B 0.011307f
C112 VTAIL.n56 B 0.011972f
C113 VTAIL.n57 B 0.026725f
C114 VTAIL.n58 B 0.057352f
C115 VTAIL.n59 B 0.011972f
C116 VTAIL.n60 B 0.011307f
C117 VTAIL.n61 B 0.04921f
C118 VTAIL.n62 B 0.032057f
C119 VTAIL.n63 B 0.100998f
C120 VTAIL.n64 B 0.029291f
C121 VTAIL.n65 B 0.021041f
C122 VTAIL.n66 B 0.011307f
C123 VTAIL.n67 B 0.026725f
C124 VTAIL.n68 B 0.011972f
C125 VTAIL.n69 B 0.021041f
C126 VTAIL.n70 B 0.011307f
C127 VTAIL.n71 B 0.026725f
C128 VTAIL.n72 B 0.011639f
C129 VTAIL.n73 B 0.021041f
C130 VTAIL.n74 B 0.011972f
C131 VTAIL.n75 B 0.026725f
C132 VTAIL.n76 B 0.011972f
C133 VTAIL.n77 B 0.021041f
C134 VTAIL.n78 B 0.011307f
C135 VTAIL.n79 B 0.026725f
C136 VTAIL.n80 B 0.011972f
C137 VTAIL.n81 B 1.0072f
C138 VTAIL.n82 B 0.011307f
C139 VTAIL.t13 B 0.04507f
C140 VTAIL.n83 B 0.147019f
C141 VTAIL.n84 B 0.018892f
C142 VTAIL.n85 B 0.020043f
C143 VTAIL.n86 B 0.026725f
C144 VTAIL.n87 B 0.011972f
C145 VTAIL.n88 B 0.011307f
C146 VTAIL.n89 B 0.021041f
C147 VTAIL.n90 B 0.021041f
C148 VTAIL.n91 B 0.011307f
C149 VTAIL.n92 B 0.011972f
C150 VTAIL.n93 B 0.026725f
C151 VTAIL.n94 B 0.026725f
C152 VTAIL.n95 B 0.011972f
C153 VTAIL.n96 B 0.011307f
C154 VTAIL.n97 B 0.021041f
C155 VTAIL.n98 B 0.021041f
C156 VTAIL.n99 B 0.011307f
C157 VTAIL.n100 B 0.011307f
C158 VTAIL.n101 B 0.011972f
C159 VTAIL.n102 B 0.026725f
C160 VTAIL.n103 B 0.026725f
C161 VTAIL.n104 B 0.026725f
C162 VTAIL.n105 B 0.011639f
C163 VTAIL.n106 B 0.011307f
C164 VTAIL.n107 B 0.021041f
C165 VTAIL.n108 B 0.021041f
C166 VTAIL.n109 B 0.011307f
C167 VTAIL.n110 B 0.011972f
C168 VTAIL.n111 B 0.026725f
C169 VTAIL.n112 B 0.026725f
C170 VTAIL.n113 B 0.011972f
C171 VTAIL.n114 B 0.011307f
C172 VTAIL.n115 B 0.021041f
C173 VTAIL.n116 B 0.021041f
C174 VTAIL.n117 B 0.011307f
C175 VTAIL.n118 B 0.011972f
C176 VTAIL.n119 B 0.026725f
C177 VTAIL.n120 B 0.057352f
C178 VTAIL.n121 B 0.011972f
C179 VTAIL.n122 B 0.011307f
C180 VTAIL.n123 B 0.04921f
C181 VTAIL.n124 B 0.032057f
C182 VTAIL.n125 B 0.100998f
C183 VTAIL.t11 B 0.189883f
C184 VTAIL.t9 B 0.189883f
C185 VTAIL.n126 B 1.6254f
C186 VTAIL.n127 B 0.308006f
C187 VTAIL.n128 B 0.029291f
C188 VTAIL.n129 B 0.021041f
C189 VTAIL.n130 B 0.011307f
C190 VTAIL.n131 B 0.026725f
C191 VTAIL.n132 B 0.011972f
C192 VTAIL.n133 B 0.021041f
C193 VTAIL.n134 B 0.011307f
C194 VTAIL.n135 B 0.026725f
C195 VTAIL.n136 B 0.011639f
C196 VTAIL.n137 B 0.021041f
C197 VTAIL.n138 B 0.011972f
C198 VTAIL.n139 B 0.026725f
C199 VTAIL.n140 B 0.011972f
C200 VTAIL.n141 B 0.021041f
C201 VTAIL.n142 B 0.011307f
C202 VTAIL.n143 B 0.026725f
C203 VTAIL.n144 B 0.011972f
C204 VTAIL.n145 B 1.0072f
C205 VTAIL.n146 B 0.011307f
C206 VTAIL.t8 B 0.04507f
C207 VTAIL.n147 B 0.147019f
C208 VTAIL.n148 B 0.018892f
C209 VTAIL.n149 B 0.020043f
C210 VTAIL.n150 B 0.026725f
C211 VTAIL.n151 B 0.011972f
C212 VTAIL.n152 B 0.011307f
C213 VTAIL.n153 B 0.021041f
C214 VTAIL.n154 B 0.021041f
C215 VTAIL.n155 B 0.011307f
C216 VTAIL.n156 B 0.011972f
C217 VTAIL.n157 B 0.026725f
C218 VTAIL.n158 B 0.026725f
C219 VTAIL.n159 B 0.011972f
C220 VTAIL.n160 B 0.011307f
C221 VTAIL.n161 B 0.021041f
C222 VTAIL.n162 B 0.021041f
C223 VTAIL.n163 B 0.011307f
C224 VTAIL.n164 B 0.011307f
C225 VTAIL.n165 B 0.011972f
C226 VTAIL.n166 B 0.026725f
C227 VTAIL.n167 B 0.026725f
C228 VTAIL.n168 B 0.026725f
C229 VTAIL.n169 B 0.011639f
C230 VTAIL.n170 B 0.011307f
C231 VTAIL.n171 B 0.021041f
C232 VTAIL.n172 B 0.021041f
C233 VTAIL.n173 B 0.011307f
C234 VTAIL.n174 B 0.011972f
C235 VTAIL.n175 B 0.026725f
C236 VTAIL.n176 B 0.026725f
C237 VTAIL.n177 B 0.011972f
C238 VTAIL.n178 B 0.011307f
C239 VTAIL.n179 B 0.021041f
C240 VTAIL.n180 B 0.021041f
C241 VTAIL.n181 B 0.011307f
C242 VTAIL.n182 B 0.011972f
C243 VTAIL.n183 B 0.026725f
C244 VTAIL.n184 B 0.057352f
C245 VTAIL.n185 B 0.011972f
C246 VTAIL.n186 B 0.011307f
C247 VTAIL.n187 B 0.04921f
C248 VTAIL.n188 B 0.032057f
C249 VTAIL.n189 B 1.07328f
C250 VTAIL.n190 B 0.029291f
C251 VTAIL.n191 B 0.021041f
C252 VTAIL.n192 B 0.011307f
C253 VTAIL.n193 B 0.026725f
C254 VTAIL.n194 B 0.011972f
C255 VTAIL.n195 B 0.021041f
C256 VTAIL.n196 B 0.011307f
C257 VTAIL.n197 B 0.026725f
C258 VTAIL.n198 B 0.011639f
C259 VTAIL.n199 B 0.021041f
C260 VTAIL.n200 B 0.011639f
C261 VTAIL.n201 B 0.011307f
C262 VTAIL.n202 B 0.026725f
C263 VTAIL.n203 B 0.026725f
C264 VTAIL.n204 B 0.011972f
C265 VTAIL.n205 B 0.021041f
C266 VTAIL.n206 B 0.011307f
C267 VTAIL.n207 B 0.026725f
C268 VTAIL.n208 B 0.011972f
C269 VTAIL.n209 B 1.0072f
C270 VTAIL.n210 B 0.011307f
C271 VTAIL.t3 B 0.04507f
C272 VTAIL.n211 B 0.147019f
C273 VTAIL.n212 B 0.018892f
C274 VTAIL.n213 B 0.020043f
C275 VTAIL.n214 B 0.026725f
C276 VTAIL.n215 B 0.011972f
C277 VTAIL.n216 B 0.011307f
C278 VTAIL.n217 B 0.021041f
C279 VTAIL.n218 B 0.021041f
C280 VTAIL.n219 B 0.011307f
C281 VTAIL.n220 B 0.011972f
C282 VTAIL.n221 B 0.026725f
C283 VTAIL.n222 B 0.026725f
C284 VTAIL.n223 B 0.011972f
C285 VTAIL.n224 B 0.011307f
C286 VTAIL.n225 B 0.021041f
C287 VTAIL.n226 B 0.021041f
C288 VTAIL.n227 B 0.011307f
C289 VTAIL.n228 B 0.011972f
C290 VTAIL.n229 B 0.026725f
C291 VTAIL.n230 B 0.026725f
C292 VTAIL.n231 B 0.011972f
C293 VTAIL.n232 B 0.011307f
C294 VTAIL.n233 B 0.021041f
C295 VTAIL.n234 B 0.021041f
C296 VTAIL.n235 B 0.011307f
C297 VTAIL.n236 B 0.011972f
C298 VTAIL.n237 B 0.026725f
C299 VTAIL.n238 B 0.026725f
C300 VTAIL.n239 B 0.011972f
C301 VTAIL.n240 B 0.011307f
C302 VTAIL.n241 B 0.021041f
C303 VTAIL.n242 B 0.021041f
C304 VTAIL.n243 B 0.011307f
C305 VTAIL.n244 B 0.011972f
C306 VTAIL.n245 B 0.026725f
C307 VTAIL.n246 B 0.057352f
C308 VTAIL.n247 B 0.011972f
C309 VTAIL.n248 B 0.011307f
C310 VTAIL.n249 B 0.04921f
C311 VTAIL.n250 B 0.032057f
C312 VTAIL.n251 B 1.07328f
C313 VTAIL.t0 B 0.189883f
C314 VTAIL.t4 B 0.189883f
C315 VTAIL.n252 B 1.62541f
C316 VTAIL.n253 B 0.307996f
C317 VTAIL.n254 B 0.029291f
C318 VTAIL.n255 B 0.021041f
C319 VTAIL.n256 B 0.011307f
C320 VTAIL.n257 B 0.026725f
C321 VTAIL.n258 B 0.011972f
C322 VTAIL.n259 B 0.021041f
C323 VTAIL.n260 B 0.011307f
C324 VTAIL.n261 B 0.026725f
C325 VTAIL.n262 B 0.011639f
C326 VTAIL.n263 B 0.021041f
C327 VTAIL.n264 B 0.011639f
C328 VTAIL.n265 B 0.011307f
C329 VTAIL.n266 B 0.026725f
C330 VTAIL.n267 B 0.026725f
C331 VTAIL.n268 B 0.011972f
C332 VTAIL.n269 B 0.021041f
C333 VTAIL.n270 B 0.011307f
C334 VTAIL.n271 B 0.026725f
C335 VTAIL.n272 B 0.011972f
C336 VTAIL.n273 B 1.0072f
C337 VTAIL.n274 B 0.011307f
C338 VTAIL.t1 B 0.04507f
C339 VTAIL.n275 B 0.147019f
C340 VTAIL.n276 B 0.018892f
C341 VTAIL.n277 B 0.020043f
C342 VTAIL.n278 B 0.026725f
C343 VTAIL.n279 B 0.011972f
C344 VTAIL.n280 B 0.011307f
C345 VTAIL.n281 B 0.021041f
C346 VTAIL.n282 B 0.021041f
C347 VTAIL.n283 B 0.011307f
C348 VTAIL.n284 B 0.011972f
C349 VTAIL.n285 B 0.026725f
C350 VTAIL.n286 B 0.026725f
C351 VTAIL.n287 B 0.011972f
C352 VTAIL.n288 B 0.011307f
C353 VTAIL.n289 B 0.021041f
C354 VTAIL.n290 B 0.021041f
C355 VTAIL.n291 B 0.011307f
C356 VTAIL.n292 B 0.011972f
C357 VTAIL.n293 B 0.026725f
C358 VTAIL.n294 B 0.026725f
C359 VTAIL.n295 B 0.011972f
C360 VTAIL.n296 B 0.011307f
C361 VTAIL.n297 B 0.021041f
C362 VTAIL.n298 B 0.021041f
C363 VTAIL.n299 B 0.011307f
C364 VTAIL.n300 B 0.011972f
C365 VTAIL.n301 B 0.026725f
C366 VTAIL.n302 B 0.026725f
C367 VTAIL.n303 B 0.011972f
C368 VTAIL.n304 B 0.011307f
C369 VTAIL.n305 B 0.021041f
C370 VTAIL.n306 B 0.021041f
C371 VTAIL.n307 B 0.011307f
C372 VTAIL.n308 B 0.011972f
C373 VTAIL.n309 B 0.026725f
C374 VTAIL.n310 B 0.057352f
C375 VTAIL.n311 B 0.011972f
C376 VTAIL.n312 B 0.011307f
C377 VTAIL.n313 B 0.04921f
C378 VTAIL.n314 B 0.032057f
C379 VTAIL.n315 B 0.100998f
C380 VTAIL.n316 B 0.029291f
C381 VTAIL.n317 B 0.021041f
C382 VTAIL.n318 B 0.011307f
C383 VTAIL.n319 B 0.026725f
C384 VTAIL.n320 B 0.011972f
C385 VTAIL.n321 B 0.021041f
C386 VTAIL.n322 B 0.011307f
C387 VTAIL.n323 B 0.026725f
C388 VTAIL.n324 B 0.011639f
C389 VTAIL.n325 B 0.021041f
C390 VTAIL.n326 B 0.011639f
C391 VTAIL.n327 B 0.011307f
C392 VTAIL.n328 B 0.026725f
C393 VTAIL.n329 B 0.026725f
C394 VTAIL.n330 B 0.011972f
C395 VTAIL.n331 B 0.021041f
C396 VTAIL.n332 B 0.011307f
C397 VTAIL.n333 B 0.026725f
C398 VTAIL.n334 B 0.011972f
C399 VTAIL.n335 B 1.0072f
C400 VTAIL.n336 B 0.011307f
C401 VTAIL.t10 B 0.04507f
C402 VTAIL.n337 B 0.147019f
C403 VTAIL.n338 B 0.018892f
C404 VTAIL.n339 B 0.020043f
C405 VTAIL.n340 B 0.026725f
C406 VTAIL.n341 B 0.011972f
C407 VTAIL.n342 B 0.011307f
C408 VTAIL.n343 B 0.021041f
C409 VTAIL.n344 B 0.021041f
C410 VTAIL.n345 B 0.011307f
C411 VTAIL.n346 B 0.011972f
C412 VTAIL.n347 B 0.026725f
C413 VTAIL.n348 B 0.026725f
C414 VTAIL.n349 B 0.011972f
C415 VTAIL.n350 B 0.011307f
C416 VTAIL.n351 B 0.021041f
C417 VTAIL.n352 B 0.021041f
C418 VTAIL.n353 B 0.011307f
C419 VTAIL.n354 B 0.011972f
C420 VTAIL.n355 B 0.026725f
C421 VTAIL.n356 B 0.026725f
C422 VTAIL.n357 B 0.011972f
C423 VTAIL.n358 B 0.011307f
C424 VTAIL.n359 B 0.021041f
C425 VTAIL.n360 B 0.021041f
C426 VTAIL.n361 B 0.011307f
C427 VTAIL.n362 B 0.011972f
C428 VTAIL.n363 B 0.026725f
C429 VTAIL.n364 B 0.026725f
C430 VTAIL.n365 B 0.011972f
C431 VTAIL.n366 B 0.011307f
C432 VTAIL.n367 B 0.021041f
C433 VTAIL.n368 B 0.021041f
C434 VTAIL.n369 B 0.011307f
C435 VTAIL.n370 B 0.011972f
C436 VTAIL.n371 B 0.026725f
C437 VTAIL.n372 B 0.057352f
C438 VTAIL.n373 B 0.011972f
C439 VTAIL.n374 B 0.011307f
C440 VTAIL.n375 B 0.04921f
C441 VTAIL.n376 B 0.032057f
C442 VTAIL.n377 B 0.100998f
C443 VTAIL.t12 B 0.189883f
C444 VTAIL.t14 B 0.189883f
C445 VTAIL.n378 B 1.62541f
C446 VTAIL.n379 B 0.307996f
C447 VTAIL.n380 B 0.029291f
C448 VTAIL.n381 B 0.021041f
C449 VTAIL.n382 B 0.011307f
C450 VTAIL.n383 B 0.026725f
C451 VTAIL.n384 B 0.011972f
C452 VTAIL.n385 B 0.021041f
C453 VTAIL.n386 B 0.011307f
C454 VTAIL.n387 B 0.026725f
C455 VTAIL.n388 B 0.011639f
C456 VTAIL.n389 B 0.021041f
C457 VTAIL.n390 B 0.011639f
C458 VTAIL.n391 B 0.011307f
C459 VTAIL.n392 B 0.026725f
C460 VTAIL.n393 B 0.026725f
C461 VTAIL.n394 B 0.011972f
C462 VTAIL.n395 B 0.021041f
C463 VTAIL.n396 B 0.011307f
C464 VTAIL.n397 B 0.026725f
C465 VTAIL.n398 B 0.011972f
C466 VTAIL.n399 B 1.0072f
C467 VTAIL.n400 B 0.011307f
C468 VTAIL.t7 B 0.04507f
C469 VTAIL.n401 B 0.147019f
C470 VTAIL.n402 B 0.018892f
C471 VTAIL.n403 B 0.020043f
C472 VTAIL.n404 B 0.026725f
C473 VTAIL.n405 B 0.011972f
C474 VTAIL.n406 B 0.011307f
C475 VTAIL.n407 B 0.021041f
C476 VTAIL.n408 B 0.021041f
C477 VTAIL.n409 B 0.011307f
C478 VTAIL.n410 B 0.011972f
C479 VTAIL.n411 B 0.026725f
C480 VTAIL.n412 B 0.026725f
C481 VTAIL.n413 B 0.011972f
C482 VTAIL.n414 B 0.011307f
C483 VTAIL.n415 B 0.021041f
C484 VTAIL.n416 B 0.021041f
C485 VTAIL.n417 B 0.011307f
C486 VTAIL.n418 B 0.011972f
C487 VTAIL.n419 B 0.026725f
C488 VTAIL.n420 B 0.026725f
C489 VTAIL.n421 B 0.011972f
C490 VTAIL.n422 B 0.011307f
C491 VTAIL.n423 B 0.021041f
C492 VTAIL.n424 B 0.021041f
C493 VTAIL.n425 B 0.011307f
C494 VTAIL.n426 B 0.011972f
C495 VTAIL.n427 B 0.026725f
C496 VTAIL.n428 B 0.026725f
C497 VTAIL.n429 B 0.011972f
C498 VTAIL.n430 B 0.011307f
C499 VTAIL.n431 B 0.021041f
C500 VTAIL.n432 B 0.021041f
C501 VTAIL.n433 B 0.011307f
C502 VTAIL.n434 B 0.011972f
C503 VTAIL.n435 B 0.026725f
C504 VTAIL.n436 B 0.057352f
C505 VTAIL.n437 B 0.011972f
C506 VTAIL.n438 B 0.011307f
C507 VTAIL.n439 B 0.04921f
C508 VTAIL.n440 B 0.032057f
C509 VTAIL.n441 B 1.07328f
C510 VTAIL.n442 B 0.029291f
C511 VTAIL.n443 B 0.021041f
C512 VTAIL.n444 B 0.011307f
C513 VTAIL.n445 B 0.026725f
C514 VTAIL.n446 B 0.011972f
C515 VTAIL.n447 B 0.021041f
C516 VTAIL.n448 B 0.011307f
C517 VTAIL.n449 B 0.026725f
C518 VTAIL.n450 B 0.011639f
C519 VTAIL.n451 B 0.021041f
C520 VTAIL.n452 B 0.011972f
C521 VTAIL.n453 B 0.026725f
C522 VTAIL.n454 B 0.011972f
C523 VTAIL.n455 B 0.021041f
C524 VTAIL.n456 B 0.011307f
C525 VTAIL.n457 B 0.026725f
C526 VTAIL.n458 B 0.011972f
C527 VTAIL.n459 B 1.0072f
C528 VTAIL.n460 B 0.011307f
C529 VTAIL.t5 B 0.04507f
C530 VTAIL.n461 B 0.147019f
C531 VTAIL.n462 B 0.018892f
C532 VTAIL.n463 B 0.020043f
C533 VTAIL.n464 B 0.026725f
C534 VTAIL.n465 B 0.011972f
C535 VTAIL.n466 B 0.011307f
C536 VTAIL.n467 B 0.021041f
C537 VTAIL.n468 B 0.021041f
C538 VTAIL.n469 B 0.011307f
C539 VTAIL.n470 B 0.011972f
C540 VTAIL.n471 B 0.026725f
C541 VTAIL.n472 B 0.026725f
C542 VTAIL.n473 B 0.011972f
C543 VTAIL.n474 B 0.011307f
C544 VTAIL.n475 B 0.021041f
C545 VTAIL.n476 B 0.021041f
C546 VTAIL.n477 B 0.011307f
C547 VTAIL.n478 B 0.011307f
C548 VTAIL.n479 B 0.011972f
C549 VTAIL.n480 B 0.026725f
C550 VTAIL.n481 B 0.026725f
C551 VTAIL.n482 B 0.026725f
C552 VTAIL.n483 B 0.011639f
C553 VTAIL.n484 B 0.011307f
C554 VTAIL.n485 B 0.021041f
C555 VTAIL.n486 B 0.021041f
C556 VTAIL.n487 B 0.011307f
C557 VTAIL.n488 B 0.011972f
C558 VTAIL.n489 B 0.026725f
C559 VTAIL.n490 B 0.026725f
C560 VTAIL.n491 B 0.011972f
C561 VTAIL.n492 B 0.011307f
C562 VTAIL.n493 B 0.021041f
C563 VTAIL.n494 B 0.021041f
C564 VTAIL.n495 B 0.011307f
C565 VTAIL.n496 B 0.011972f
C566 VTAIL.n497 B 0.026725f
C567 VTAIL.n498 B 0.057352f
C568 VTAIL.n499 B 0.011972f
C569 VTAIL.n500 B 0.011307f
C570 VTAIL.n501 B 0.04921f
C571 VTAIL.n502 B 0.032057f
C572 VTAIL.n503 B 1.06933f
C573 VDD1.t5 B 0.259603f
C574 VDD1.t0 B 0.259603f
C575 VDD1.n0 B 2.30895f
C576 VDD1.t2 B 0.259603f
C577 VDD1.t4 B 0.259603f
C578 VDD1.n1 B 2.30826f
C579 VDD1.t3 B 0.259603f
C580 VDD1.t7 B 0.259603f
C581 VDD1.n2 B 2.30826f
C582 VDD1.n3 B 2.41268f
C583 VDD1.t6 B 0.259603f
C584 VDD1.t1 B 0.259603f
C585 VDD1.n4 B 2.30647f
C586 VDD1.n5 B 2.55338f
C587 VP.n0 B 0.048535f
C588 VP.t3 B 0.854218f
C589 VP.n1 B 0.348024f
C590 VP.n2 B 0.048535f
C591 VP.t7 B 0.854218f
C592 VP.t0 B 0.854218f
C593 VP.n3 B 0.197668f
C594 VP.t2 B 0.854218f
C595 VP.t4 B 0.868684f
C596 VP.n4 B 0.334722f
C597 VP.n5 B 0.356142f
C598 VP.n6 B 0.348024f
C599 VP.n7 B 0.011014f
C600 VP.n8 B 0.345331f
C601 VP.n9 B 1.90577f
C602 VP.n10 B 1.94868f
C603 VP.t6 B 0.854218f
C604 VP.n11 B 0.345331f
C605 VP.n12 B 0.011014f
C606 VP.n13 B 0.048535f
C607 VP.n14 B 0.048535f
C608 VP.n15 B 0.048535f
C609 VP.t5 B 0.854218f
C610 VP.n16 B 0.348024f
C611 VP.n17 B 0.011014f
C612 VP.t1 B 0.854218f
C613 VP.n18 B 0.345331f
C614 VP.n19 B 0.037613f
.ends

