* NGSPICE file created from diff_pair_sample_1123.ext - technology: sky130A

.subckt diff_pair_sample_1123 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=1.7754 ps=11.09 w=10.76 l=3.26
X1 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=4.1964 ps=22.3 w=10.76 l=3.26
X2 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=0 ps=0 w=10.76 l=3.26
X3 VTAIL.t9 VP.t1 VDD1.t4 B.t19 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=1.7754 ps=11.09 w=10.76 l=3.26
X4 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=0 ps=0 w=10.76 l=3.26
X5 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=0 ps=0 w=10.76 l=3.26
X6 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=0 ps=0 w=10.76 l=3.26
X7 VTAIL.t0 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=1.7754 ps=11.09 w=10.76 l=3.26
X8 VDD2.t3 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=4.1964 ps=22.3 w=10.76 l=3.26
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=1.7754 ps=11.09 w=10.76 l=3.26
X10 VTAIL.t11 VN.t4 VDD2.t1 B.t19 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=1.7754 ps=11.09 w=10.76 l=3.26
X11 VDD1.t3 VP.t2 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=4.1964 ps=22.3 w=10.76 l=3.26
X12 VDD1.t0 VP.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=1.7754 ps=11.09 w=10.76 l=3.26
X13 VDD1.t2 VP.t4 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=1.7754 ps=11.09 w=10.76 l=3.26
X14 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.1964 pd=22.3 as=1.7754 ps=11.09 w=10.76 l=3.26
X15 VDD1.t5 VP.t5 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7754 pd=11.09 as=4.1964 ps=22.3 w=10.76 l=3.26
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t4 112.769
R22 VP.n8 VP.t3 79.5453
R23 VP.n4 VP.t1 79.5453
R24 VP.n0 VP.t2 79.5453
R25 VP.n9 VP.t5 79.5453
R26 VP.n13 VP.t0 79.5453
R27 VP.n27 VP.n8 73.5231
R28 VP.n50 VP.n0 73.5231
R29 VP.n26 VP.n9 73.5231
R30 VP.n14 VP.n13 62.2205
R31 VP.n27 VP.n26 50.4579
R32 VP.n31 VP.n6 44.9365
R33 VP.n46 VP.n2 44.9365
R34 VP.n22 VP.n11 44.9365
R35 VP.n35 VP.n6 36.2176
R36 VP.n42 VP.n2 36.2176
R37 VP.n18 VP.n11 36.2176
R38 VP.n30 VP.n29 24.5923
R39 VP.n31 VP.n30 24.5923
R40 VP.n36 VP.n35 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n41 VP.n40 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n46 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n23 VP.n22 24.5923
R47 VP.n24 VP.n23 24.5923
R48 VP.n17 VP.n16 24.5923
R49 VP.n18 VP.n17 24.5923
R50 VP.n29 VP.n8 16.7229
R51 VP.n48 VP.n0 16.7229
R52 VP.n24 VP.n9 16.7229
R53 VP.n37 VP.n4 12.2964
R54 VP.n40 VP.n4 12.2964
R55 VP.n16 VP.n13 12.2964
R56 VP.n15 VP.n14 4.04952
R57 VP.n26 VP.n25 0.354861
R58 VP.n28 VP.n27 0.354861
R59 VP.n50 VP.n49 0.354861
R60 VP VP.n50 0.267071
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1.n52 VDD1.n0 289.615
R81 VDD1.n109 VDD1.n57 289.615
R82 VDD1.n53 VDD1.n52 185
R83 VDD1.n51 VDD1.n50 185
R84 VDD1.n4 VDD1.n3 185
R85 VDD1.n45 VDD1.n44 185
R86 VDD1.n43 VDD1.n42 185
R87 VDD1.n41 VDD1.n7 185
R88 VDD1.n11 VDD1.n8 185
R89 VDD1.n36 VDD1.n35 185
R90 VDD1.n34 VDD1.n33 185
R91 VDD1.n13 VDD1.n12 185
R92 VDD1.n28 VDD1.n27 185
R93 VDD1.n26 VDD1.n25 185
R94 VDD1.n17 VDD1.n16 185
R95 VDD1.n20 VDD1.n19 185
R96 VDD1.n76 VDD1.n75 185
R97 VDD1.n73 VDD1.n72 185
R98 VDD1.n82 VDD1.n81 185
R99 VDD1.n84 VDD1.n83 185
R100 VDD1.n69 VDD1.n68 185
R101 VDD1.n90 VDD1.n89 185
R102 VDD1.n93 VDD1.n92 185
R103 VDD1.n91 VDD1.n65 185
R104 VDD1.n98 VDD1.n64 185
R105 VDD1.n100 VDD1.n99 185
R106 VDD1.n102 VDD1.n101 185
R107 VDD1.n61 VDD1.n60 185
R108 VDD1.n108 VDD1.n107 185
R109 VDD1.n110 VDD1.n109 185
R110 VDD1.t2 VDD1.n18 149.524
R111 VDD1.t0 VDD1.n74 149.524
R112 VDD1.n52 VDD1.n51 104.615
R113 VDD1.n51 VDD1.n3 104.615
R114 VDD1.n44 VDD1.n3 104.615
R115 VDD1.n44 VDD1.n43 104.615
R116 VDD1.n43 VDD1.n7 104.615
R117 VDD1.n11 VDD1.n7 104.615
R118 VDD1.n35 VDD1.n11 104.615
R119 VDD1.n35 VDD1.n34 104.615
R120 VDD1.n34 VDD1.n12 104.615
R121 VDD1.n27 VDD1.n12 104.615
R122 VDD1.n27 VDD1.n26 104.615
R123 VDD1.n26 VDD1.n16 104.615
R124 VDD1.n19 VDD1.n16 104.615
R125 VDD1.n75 VDD1.n72 104.615
R126 VDD1.n82 VDD1.n72 104.615
R127 VDD1.n83 VDD1.n82 104.615
R128 VDD1.n83 VDD1.n68 104.615
R129 VDD1.n90 VDD1.n68 104.615
R130 VDD1.n92 VDD1.n90 104.615
R131 VDD1.n92 VDD1.n91 104.615
R132 VDD1.n91 VDD1.n64 104.615
R133 VDD1.n100 VDD1.n64 104.615
R134 VDD1.n101 VDD1.n100 104.615
R135 VDD1.n101 VDD1.n60 104.615
R136 VDD1.n108 VDD1.n60 104.615
R137 VDD1.n109 VDD1.n108 104.615
R138 VDD1.n115 VDD1.n114 64.61
R139 VDD1.n117 VDD1.n116 63.8916
R140 VDD1 VDD1.n56 52.795
R141 VDD1.n115 VDD1.n113 52.6814
R142 VDD1.n19 VDD1.t2 52.3082
R143 VDD1.n75 VDD1.t0 52.3082
R144 VDD1.n117 VDD1.n115 45.1798
R145 VDD1.n42 VDD1.n41 13.1884
R146 VDD1.n99 VDD1.n98 13.1884
R147 VDD1.n45 VDD1.n6 12.8005
R148 VDD1.n40 VDD1.n8 12.8005
R149 VDD1.n97 VDD1.n65 12.8005
R150 VDD1.n102 VDD1.n63 12.8005
R151 VDD1.n46 VDD1.n4 12.0247
R152 VDD1.n37 VDD1.n36 12.0247
R153 VDD1.n94 VDD1.n93 12.0247
R154 VDD1.n103 VDD1.n61 12.0247
R155 VDD1.n50 VDD1.n49 11.249
R156 VDD1.n33 VDD1.n10 11.249
R157 VDD1.n89 VDD1.n67 11.249
R158 VDD1.n107 VDD1.n106 11.249
R159 VDD1.n53 VDD1.n2 10.4732
R160 VDD1.n32 VDD1.n13 10.4732
R161 VDD1.n88 VDD1.n69 10.4732
R162 VDD1.n110 VDD1.n59 10.4732
R163 VDD1.n20 VDD1.n18 10.2747
R164 VDD1.n76 VDD1.n74 10.2747
R165 VDD1.n54 VDD1.n0 9.69747
R166 VDD1.n29 VDD1.n28 9.69747
R167 VDD1.n85 VDD1.n84 9.69747
R168 VDD1.n111 VDD1.n57 9.69747
R169 VDD1.n56 VDD1.n55 9.45567
R170 VDD1.n113 VDD1.n112 9.45567
R171 VDD1.n22 VDD1.n21 9.3005
R172 VDD1.n24 VDD1.n23 9.3005
R173 VDD1.n15 VDD1.n14 9.3005
R174 VDD1.n30 VDD1.n29 9.3005
R175 VDD1.n32 VDD1.n31 9.3005
R176 VDD1.n10 VDD1.n9 9.3005
R177 VDD1.n38 VDD1.n37 9.3005
R178 VDD1.n40 VDD1.n39 9.3005
R179 VDD1.n55 VDD1.n54 9.3005
R180 VDD1.n2 VDD1.n1 9.3005
R181 VDD1.n49 VDD1.n48 9.3005
R182 VDD1.n47 VDD1.n46 9.3005
R183 VDD1.n6 VDD1.n5 9.3005
R184 VDD1.n112 VDD1.n111 9.3005
R185 VDD1.n59 VDD1.n58 9.3005
R186 VDD1.n106 VDD1.n105 9.3005
R187 VDD1.n104 VDD1.n103 9.3005
R188 VDD1.n63 VDD1.n62 9.3005
R189 VDD1.n78 VDD1.n77 9.3005
R190 VDD1.n80 VDD1.n79 9.3005
R191 VDD1.n71 VDD1.n70 9.3005
R192 VDD1.n86 VDD1.n85 9.3005
R193 VDD1.n88 VDD1.n87 9.3005
R194 VDD1.n67 VDD1.n66 9.3005
R195 VDD1.n95 VDD1.n94 9.3005
R196 VDD1.n97 VDD1.n96 9.3005
R197 VDD1.n25 VDD1.n15 8.92171
R198 VDD1.n81 VDD1.n71 8.92171
R199 VDD1.n24 VDD1.n17 8.14595
R200 VDD1.n80 VDD1.n73 8.14595
R201 VDD1.n21 VDD1.n20 7.3702
R202 VDD1.n77 VDD1.n76 7.3702
R203 VDD1.n21 VDD1.n17 5.81868
R204 VDD1.n77 VDD1.n73 5.81868
R205 VDD1.n25 VDD1.n24 5.04292
R206 VDD1.n81 VDD1.n80 5.04292
R207 VDD1.n56 VDD1.n0 4.26717
R208 VDD1.n28 VDD1.n15 4.26717
R209 VDD1.n84 VDD1.n71 4.26717
R210 VDD1.n113 VDD1.n57 4.26717
R211 VDD1.n54 VDD1.n53 3.49141
R212 VDD1.n29 VDD1.n13 3.49141
R213 VDD1.n85 VDD1.n69 3.49141
R214 VDD1.n111 VDD1.n110 3.49141
R215 VDD1.n22 VDD1.n18 2.84303
R216 VDD1.n78 VDD1.n74 2.84303
R217 VDD1.n50 VDD1.n2 2.71565
R218 VDD1.n33 VDD1.n32 2.71565
R219 VDD1.n89 VDD1.n88 2.71565
R220 VDD1.n107 VDD1.n59 2.71565
R221 VDD1.n49 VDD1.n4 1.93989
R222 VDD1.n36 VDD1.n10 1.93989
R223 VDD1.n93 VDD1.n67 1.93989
R224 VDD1.n106 VDD1.n61 1.93989
R225 VDD1.n116 VDD1.t1 1.84065
R226 VDD1.n116 VDD1.t5 1.84065
R227 VDD1.n114 VDD1.t4 1.84065
R228 VDD1.n114 VDD1.t3 1.84065
R229 VDD1.n46 VDD1.n45 1.16414
R230 VDD1.n37 VDD1.n8 1.16414
R231 VDD1.n94 VDD1.n65 1.16414
R232 VDD1.n103 VDD1.n102 1.16414
R233 VDD1 VDD1.n117 0.716017
R234 VDD1.n42 VDD1.n6 0.388379
R235 VDD1.n41 VDD1.n40 0.388379
R236 VDD1.n98 VDD1.n97 0.388379
R237 VDD1.n99 VDD1.n63 0.388379
R238 VDD1.n55 VDD1.n1 0.155672
R239 VDD1.n48 VDD1.n1 0.155672
R240 VDD1.n48 VDD1.n47 0.155672
R241 VDD1.n47 VDD1.n5 0.155672
R242 VDD1.n39 VDD1.n5 0.155672
R243 VDD1.n39 VDD1.n38 0.155672
R244 VDD1.n38 VDD1.n9 0.155672
R245 VDD1.n31 VDD1.n9 0.155672
R246 VDD1.n31 VDD1.n30 0.155672
R247 VDD1.n30 VDD1.n14 0.155672
R248 VDD1.n23 VDD1.n14 0.155672
R249 VDD1.n23 VDD1.n22 0.155672
R250 VDD1.n79 VDD1.n78 0.155672
R251 VDD1.n79 VDD1.n70 0.155672
R252 VDD1.n86 VDD1.n70 0.155672
R253 VDD1.n87 VDD1.n86 0.155672
R254 VDD1.n87 VDD1.n66 0.155672
R255 VDD1.n95 VDD1.n66 0.155672
R256 VDD1.n96 VDD1.n95 0.155672
R257 VDD1.n96 VDD1.n62 0.155672
R258 VDD1.n104 VDD1.n62 0.155672
R259 VDD1.n105 VDD1.n104 0.155672
R260 VDD1.n105 VDD1.n58 0.155672
R261 VDD1.n112 VDD1.n58 0.155672
R262 VTAIL.n234 VTAIL.n182 289.615
R263 VTAIL.n54 VTAIL.n2 289.615
R264 VTAIL.n176 VTAIL.n124 289.615
R265 VTAIL.n116 VTAIL.n64 289.615
R266 VTAIL.n201 VTAIL.n200 185
R267 VTAIL.n198 VTAIL.n197 185
R268 VTAIL.n207 VTAIL.n206 185
R269 VTAIL.n209 VTAIL.n208 185
R270 VTAIL.n194 VTAIL.n193 185
R271 VTAIL.n215 VTAIL.n214 185
R272 VTAIL.n218 VTAIL.n217 185
R273 VTAIL.n216 VTAIL.n190 185
R274 VTAIL.n223 VTAIL.n189 185
R275 VTAIL.n225 VTAIL.n224 185
R276 VTAIL.n227 VTAIL.n226 185
R277 VTAIL.n186 VTAIL.n185 185
R278 VTAIL.n233 VTAIL.n232 185
R279 VTAIL.n235 VTAIL.n234 185
R280 VTAIL.n21 VTAIL.n20 185
R281 VTAIL.n18 VTAIL.n17 185
R282 VTAIL.n27 VTAIL.n26 185
R283 VTAIL.n29 VTAIL.n28 185
R284 VTAIL.n14 VTAIL.n13 185
R285 VTAIL.n35 VTAIL.n34 185
R286 VTAIL.n38 VTAIL.n37 185
R287 VTAIL.n36 VTAIL.n10 185
R288 VTAIL.n43 VTAIL.n9 185
R289 VTAIL.n45 VTAIL.n44 185
R290 VTAIL.n47 VTAIL.n46 185
R291 VTAIL.n6 VTAIL.n5 185
R292 VTAIL.n53 VTAIL.n52 185
R293 VTAIL.n55 VTAIL.n54 185
R294 VTAIL.n177 VTAIL.n176 185
R295 VTAIL.n175 VTAIL.n174 185
R296 VTAIL.n128 VTAIL.n127 185
R297 VTAIL.n169 VTAIL.n168 185
R298 VTAIL.n167 VTAIL.n166 185
R299 VTAIL.n165 VTAIL.n131 185
R300 VTAIL.n135 VTAIL.n132 185
R301 VTAIL.n160 VTAIL.n159 185
R302 VTAIL.n158 VTAIL.n157 185
R303 VTAIL.n137 VTAIL.n136 185
R304 VTAIL.n152 VTAIL.n151 185
R305 VTAIL.n150 VTAIL.n149 185
R306 VTAIL.n141 VTAIL.n140 185
R307 VTAIL.n144 VTAIL.n143 185
R308 VTAIL.n117 VTAIL.n116 185
R309 VTAIL.n115 VTAIL.n114 185
R310 VTAIL.n68 VTAIL.n67 185
R311 VTAIL.n109 VTAIL.n108 185
R312 VTAIL.n107 VTAIL.n106 185
R313 VTAIL.n105 VTAIL.n71 185
R314 VTAIL.n75 VTAIL.n72 185
R315 VTAIL.n100 VTAIL.n99 185
R316 VTAIL.n98 VTAIL.n97 185
R317 VTAIL.n77 VTAIL.n76 185
R318 VTAIL.n92 VTAIL.n91 185
R319 VTAIL.n90 VTAIL.n89 185
R320 VTAIL.n81 VTAIL.n80 185
R321 VTAIL.n84 VTAIL.n83 185
R322 VTAIL.t3 VTAIL.n199 149.524
R323 VTAIL.t8 VTAIL.n19 149.524
R324 VTAIL.t5 VTAIL.n142 149.524
R325 VTAIL.t4 VTAIL.n82 149.524
R326 VTAIL.n200 VTAIL.n197 104.615
R327 VTAIL.n207 VTAIL.n197 104.615
R328 VTAIL.n208 VTAIL.n207 104.615
R329 VTAIL.n208 VTAIL.n193 104.615
R330 VTAIL.n215 VTAIL.n193 104.615
R331 VTAIL.n217 VTAIL.n215 104.615
R332 VTAIL.n217 VTAIL.n216 104.615
R333 VTAIL.n216 VTAIL.n189 104.615
R334 VTAIL.n225 VTAIL.n189 104.615
R335 VTAIL.n226 VTAIL.n225 104.615
R336 VTAIL.n226 VTAIL.n185 104.615
R337 VTAIL.n233 VTAIL.n185 104.615
R338 VTAIL.n234 VTAIL.n233 104.615
R339 VTAIL.n20 VTAIL.n17 104.615
R340 VTAIL.n27 VTAIL.n17 104.615
R341 VTAIL.n28 VTAIL.n27 104.615
R342 VTAIL.n28 VTAIL.n13 104.615
R343 VTAIL.n35 VTAIL.n13 104.615
R344 VTAIL.n37 VTAIL.n35 104.615
R345 VTAIL.n37 VTAIL.n36 104.615
R346 VTAIL.n36 VTAIL.n9 104.615
R347 VTAIL.n45 VTAIL.n9 104.615
R348 VTAIL.n46 VTAIL.n45 104.615
R349 VTAIL.n46 VTAIL.n5 104.615
R350 VTAIL.n53 VTAIL.n5 104.615
R351 VTAIL.n54 VTAIL.n53 104.615
R352 VTAIL.n176 VTAIL.n175 104.615
R353 VTAIL.n175 VTAIL.n127 104.615
R354 VTAIL.n168 VTAIL.n127 104.615
R355 VTAIL.n168 VTAIL.n167 104.615
R356 VTAIL.n167 VTAIL.n131 104.615
R357 VTAIL.n135 VTAIL.n131 104.615
R358 VTAIL.n159 VTAIL.n135 104.615
R359 VTAIL.n159 VTAIL.n158 104.615
R360 VTAIL.n158 VTAIL.n136 104.615
R361 VTAIL.n151 VTAIL.n136 104.615
R362 VTAIL.n151 VTAIL.n150 104.615
R363 VTAIL.n150 VTAIL.n140 104.615
R364 VTAIL.n143 VTAIL.n140 104.615
R365 VTAIL.n116 VTAIL.n115 104.615
R366 VTAIL.n115 VTAIL.n67 104.615
R367 VTAIL.n108 VTAIL.n67 104.615
R368 VTAIL.n108 VTAIL.n107 104.615
R369 VTAIL.n107 VTAIL.n71 104.615
R370 VTAIL.n75 VTAIL.n71 104.615
R371 VTAIL.n99 VTAIL.n75 104.615
R372 VTAIL.n99 VTAIL.n98 104.615
R373 VTAIL.n98 VTAIL.n76 104.615
R374 VTAIL.n91 VTAIL.n76 104.615
R375 VTAIL.n91 VTAIL.n90 104.615
R376 VTAIL.n90 VTAIL.n80 104.615
R377 VTAIL.n83 VTAIL.n80 104.615
R378 VTAIL.n200 VTAIL.t3 52.3082
R379 VTAIL.n20 VTAIL.t8 52.3082
R380 VTAIL.n143 VTAIL.t5 52.3082
R381 VTAIL.n83 VTAIL.t4 52.3082
R382 VTAIL.n123 VTAIL.n122 47.213
R383 VTAIL.n63 VTAIL.n62 47.213
R384 VTAIL.n1 VTAIL.n0 47.2128
R385 VTAIL.n61 VTAIL.n60 47.2128
R386 VTAIL.n239 VTAIL.n238 33.7369
R387 VTAIL.n59 VTAIL.n58 33.7369
R388 VTAIL.n181 VTAIL.n180 33.7369
R389 VTAIL.n121 VTAIL.n120 33.7369
R390 VTAIL.n63 VTAIL.n61 27.8324
R391 VTAIL.n239 VTAIL.n181 24.7376
R392 VTAIL.n224 VTAIL.n223 13.1884
R393 VTAIL.n44 VTAIL.n43 13.1884
R394 VTAIL.n166 VTAIL.n165 13.1884
R395 VTAIL.n106 VTAIL.n105 13.1884
R396 VTAIL.n222 VTAIL.n190 12.8005
R397 VTAIL.n227 VTAIL.n188 12.8005
R398 VTAIL.n42 VTAIL.n10 12.8005
R399 VTAIL.n47 VTAIL.n8 12.8005
R400 VTAIL.n169 VTAIL.n130 12.8005
R401 VTAIL.n164 VTAIL.n132 12.8005
R402 VTAIL.n109 VTAIL.n70 12.8005
R403 VTAIL.n104 VTAIL.n72 12.8005
R404 VTAIL.n219 VTAIL.n218 12.0247
R405 VTAIL.n228 VTAIL.n186 12.0247
R406 VTAIL.n39 VTAIL.n38 12.0247
R407 VTAIL.n48 VTAIL.n6 12.0247
R408 VTAIL.n170 VTAIL.n128 12.0247
R409 VTAIL.n161 VTAIL.n160 12.0247
R410 VTAIL.n110 VTAIL.n68 12.0247
R411 VTAIL.n101 VTAIL.n100 12.0247
R412 VTAIL.n214 VTAIL.n192 11.249
R413 VTAIL.n232 VTAIL.n231 11.249
R414 VTAIL.n34 VTAIL.n12 11.249
R415 VTAIL.n52 VTAIL.n51 11.249
R416 VTAIL.n174 VTAIL.n173 11.249
R417 VTAIL.n157 VTAIL.n134 11.249
R418 VTAIL.n114 VTAIL.n113 11.249
R419 VTAIL.n97 VTAIL.n74 11.249
R420 VTAIL.n213 VTAIL.n194 10.4732
R421 VTAIL.n235 VTAIL.n184 10.4732
R422 VTAIL.n33 VTAIL.n14 10.4732
R423 VTAIL.n55 VTAIL.n4 10.4732
R424 VTAIL.n177 VTAIL.n126 10.4732
R425 VTAIL.n156 VTAIL.n137 10.4732
R426 VTAIL.n117 VTAIL.n66 10.4732
R427 VTAIL.n96 VTAIL.n77 10.4732
R428 VTAIL.n201 VTAIL.n199 10.2747
R429 VTAIL.n21 VTAIL.n19 10.2747
R430 VTAIL.n144 VTAIL.n142 10.2747
R431 VTAIL.n84 VTAIL.n82 10.2747
R432 VTAIL.n210 VTAIL.n209 9.69747
R433 VTAIL.n236 VTAIL.n182 9.69747
R434 VTAIL.n30 VTAIL.n29 9.69747
R435 VTAIL.n56 VTAIL.n2 9.69747
R436 VTAIL.n178 VTAIL.n124 9.69747
R437 VTAIL.n153 VTAIL.n152 9.69747
R438 VTAIL.n118 VTAIL.n64 9.69747
R439 VTAIL.n93 VTAIL.n92 9.69747
R440 VTAIL.n238 VTAIL.n237 9.45567
R441 VTAIL.n58 VTAIL.n57 9.45567
R442 VTAIL.n180 VTAIL.n179 9.45567
R443 VTAIL.n120 VTAIL.n119 9.45567
R444 VTAIL.n237 VTAIL.n236 9.3005
R445 VTAIL.n184 VTAIL.n183 9.3005
R446 VTAIL.n231 VTAIL.n230 9.3005
R447 VTAIL.n229 VTAIL.n228 9.3005
R448 VTAIL.n188 VTAIL.n187 9.3005
R449 VTAIL.n203 VTAIL.n202 9.3005
R450 VTAIL.n205 VTAIL.n204 9.3005
R451 VTAIL.n196 VTAIL.n195 9.3005
R452 VTAIL.n211 VTAIL.n210 9.3005
R453 VTAIL.n213 VTAIL.n212 9.3005
R454 VTAIL.n192 VTAIL.n191 9.3005
R455 VTAIL.n220 VTAIL.n219 9.3005
R456 VTAIL.n222 VTAIL.n221 9.3005
R457 VTAIL.n57 VTAIL.n56 9.3005
R458 VTAIL.n4 VTAIL.n3 9.3005
R459 VTAIL.n51 VTAIL.n50 9.3005
R460 VTAIL.n49 VTAIL.n48 9.3005
R461 VTAIL.n8 VTAIL.n7 9.3005
R462 VTAIL.n23 VTAIL.n22 9.3005
R463 VTAIL.n25 VTAIL.n24 9.3005
R464 VTAIL.n16 VTAIL.n15 9.3005
R465 VTAIL.n31 VTAIL.n30 9.3005
R466 VTAIL.n33 VTAIL.n32 9.3005
R467 VTAIL.n12 VTAIL.n11 9.3005
R468 VTAIL.n40 VTAIL.n39 9.3005
R469 VTAIL.n42 VTAIL.n41 9.3005
R470 VTAIL.n146 VTAIL.n145 9.3005
R471 VTAIL.n148 VTAIL.n147 9.3005
R472 VTAIL.n139 VTAIL.n138 9.3005
R473 VTAIL.n154 VTAIL.n153 9.3005
R474 VTAIL.n156 VTAIL.n155 9.3005
R475 VTAIL.n134 VTAIL.n133 9.3005
R476 VTAIL.n162 VTAIL.n161 9.3005
R477 VTAIL.n164 VTAIL.n163 9.3005
R478 VTAIL.n179 VTAIL.n178 9.3005
R479 VTAIL.n126 VTAIL.n125 9.3005
R480 VTAIL.n173 VTAIL.n172 9.3005
R481 VTAIL.n171 VTAIL.n170 9.3005
R482 VTAIL.n130 VTAIL.n129 9.3005
R483 VTAIL.n86 VTAIL.n85 9.3005
R484 VTAIL.n88 VTAIL.n87 9.3005
R485 VTAIL.n79 VTAIL.n78 9.3005
R486 VTAIL.n94 VTAIL.n93 9.3005
R487 VTAIL.n96 VTAIL.n95 9.3005
R488 VTAIL.n74 VTAIL.n73 9.3005
R489 VTAIL.n102 VTAIL.n101 9.3005
R490 VTAIL.n104 VTAIL.n103 9.3005
R491 VTAIL.n119 VTAIL.n118 9.3005
R492 VTAIL.n66 VTAIL.n65 9.3005
R493 VTAIL.n113 VTAIL.n112 9.3005
R494 VTAIL.n111 VTAIL.n110 9.3005
R495 VTAIL.n70 VTAIL.n69 9.3005
R496 VTAIL.n206 VTAIL.n196 8.92171
R497 VTAIL.n26 VTAIL.n16 8.92171
R498 VTAIL.n149 VTAIL.n139 8.92171
R499 VTAIL.n89 VTAIL.n79 8.92171
R500 VTAIL.n205 VTAIL.n198 8.14595
R501 VTAIL.n25 VTAIL.n18 8.14595
R502 VTAIL.n148 VTAIL.n141 8.14595
R503 VTAIL.n88 VTAIL.n81 8.14595
R504 VTAIL.n202 VTAIL.n201 7.3702
R505 VTAIL.n22 VTAIL.n21 7.3702
R506 VTAIL.n145 VTAIL.n144 7.3702
R507 VTAIL.n85 VTAIL.n84 7.3702
R508 VTAIL.n202 VTAIL.n198 5.81868
R509 VTAIL.n22 VTAIL.n18 5.81868
R510 VTAIL.n145 VTAIL.n141 5.81868
R511 VTAIL.n85 VTAIL.n81 5.81868
R512 VTAIL.n206 VTAIL.n205 5.04292
R513 VTAIL.n26 VTAIL.n25 5.04292
R514 VTAIL.n149 VTAIL.n148 5.04292
R515 VTAIL.n89 VTAIL.n88 5.04292
R516 VTAIL.n209 VTAIL.n196 4.26717
R517 VTAIL.n238 VTAIL.n182 4.26717
R518 VTAIL.n29 VTAIL.n16 4.26717
R519 VTAIL.n58 VTAIL.n2 4.26717
R520 VTAIL.n180 VTAIL.n124 4.26717
R521 VTAIL.n152 VTAIL.n139 4.26717
R522 VTAIL.n120 VTAIL.n64 4.26717
R523 VTAIL.n92 VTAIL.n79 4.26717
R524 VTAIL.n210 VTAIL.n194 3.49141
R525 VTAIL.n236 VTAIL.n235 3.49141
R526 VTAIL.n30 VTAIL.n14 3.49141
R527 VTAIL.n56 VTAIL.n55 3.49141
R528 VTAIL.n178 VTAIL.n177 3.49141
R529 VTAIL.n153 VTAIL.n137 3.49141
R530 VTAIL.n118 VTAIL.n117 3.49141
R531 VTAIL.n93 VTAIL.n77 3.49141
R532 VTAIL.n121 VTAIL.n63 3.09533
R533 VTAIL.n181 VTAIL.n123 3.09533
R534 VTAIL.n61 VTAIL.n59 3.09533
R535 VTAIL.n203 VTAIL.n199 2.84303
R536 VTAIL.n23 VTAIL.n19 2.84303
R537 VTAIL.n146 VTAIL.n142 2.84303
R538 VTAIL.n86 VTAIL.n82 2.84303
R539 VTAIL.n214 VTAIL.n213 2.71565
R540 VTAIL.n232 VTAIL.n184 2.71565
R541 VTAIL.n34 VTAIL.n33 2.71565
R542 VTAIL.n52 VTAIL.n4 2.71565
R543 VTAIL.n174 VTAIL.n126 2.71565
R544 VTAIL.n157 VTAIL.n156 2.71565
R545 VTAIL.n114 VTAIL.n66 2.71565
R546 VTAIL.n97 VTAIL.n96 2.71565
R547 VTAIL VTAIL.n239 2.26343
R548 VTAIL.n123 VTAIL.n121 2.01774
R549 VTAIL.n59 VTAIL.n1 2.01774
R550 VTAIL.n218 VTAIL.n192 1.93989
R551 VTAIL.n231 VTAIL.n186 1.93989
R552 VTAIL.n38 VTAIL.n12 1.93989
R553 VTAIL.n51 VTAIL.n6 1.93989
R554 VTAIL.n173 VTAIL.n128 1.93989
R555 VTAIL.n160 VTAIL.n134 1.93989
R556 VTAIL.n113 VTAIL.n68 1.93989
R557 VTAIL.n100 VTAIL.n74 1.93989
R558 VTAIL.n0 VTAIL.t1 1.84065
R559 VTAIL.n0 VTAIL.t0 1.84065
R560 VTAIL.n60 VTAIL.t7 1.84065
R561 VTAIL.n60 VTAIL.t9 1.84065
R562 VTAIL.n122 VTAIL.t6 1.84065
R563 VTAIL.n122 VTAIL.t10 1.84065
R564 VTAIL.n62 VTAIL.t2 1.84065
R565 VTAIL.n62 VTAIL.t11 1.84065
R566 VTAIL.n219 VTAIL.n190 1.16414
R567 VTAIL.n228 VTAIL.n227 1.16414
R568 VTAIL.n39 VTAIL.n10 1.16414
R569 VTAIL.n48 VTAIL.n47 1.16414
R570 VTAIL.n170 VTAIL.n169 1.16414
R571 VTAIL.n161 VTAIL.n132 1.16414
R572 VTAIL.n110 VTAIL.n109 1.16414
R573 VTAIL.n101 VTAIL.n72 1.16414
R574 VTAIL VTAIL.n1 0.832397
R575 VTAIL.n223 VTAIL.n222 0.388379
R576 VTAIL.n224 VTAIL.n188 0.388379
R577 VTAIL.n43 VTAIL.n42 0.388379
R578 VTAIL.n44 VTAIL.n8 0.388379
R579 VTAIL.n166 VTAIL.n130 0.388379
R580 VTAIL.n165 VTAIL.n164 0.388379
R581 VTAIL.n106 VTAIL.n70 0.388379
R582 VTAIL.n105 VTAIL.n104 0.388379
R583 VTAIL.n204 VTAIL.n203 0.155672
R584 VTAIL.n204 VTAIL.n195 0.155672
R585 VTAIL.n211 VTAIL.n195 0.155672
R586 VTAIL.n212 VTAIL.n211 0.155672
R587 VTAIL.n212 VTAIL.n191 0.155672
R588 VTAIL.n220 VTAIL.n191 0.155672
R589 VTAIL.n221 VTAIL.n220 0.155672
R590 VTAIL.n221 VTAIL.n187 0.155672
R591 VTAIL.n229 VTAIL.n187 0.155672
R592 VTAIL.n230 VTAIL.n229 0.155672
R593 VTAIL.n230 VTAIL.n183 0.155672
R594 VTAIL.n237 VTAIL.n183 0.155672
R595 VTAIL.n24 VTAIL.n23 0.155672
R596 VTAIL.n24 VTAIL.n15 0.155672
R597 VTAIL.n31 VTAIL.n15 0.155672
R598 VTAIL.n32 VTAIL.n31 0.155672
R599 VTAIL.n32 VTAIL.n11 0.155672
R600 VTAIL.n40 VTAIL.n11 0.155672
R601 VTAIL.n41 VTAIL.n40 0.155672
R602 VTAIL.n41 VTAIL.n7 0.155672
R603 VTAIL.n49 VTAIL.n7 0.155672
R604 VTAIL.n50 VTAIL.n49 0.155672
R605 VTAIL.n50 VTAIL.n3 0.155672
R606 VTAIL.n57 VTAIL.n3 0.155672
R607 VTAIL.n179 VTAIL.n125 0.155672
R608 VTAIL.n172 VTAIL.n125 0.155672
R609 VTAIL.n172 VTAIL.n171 0.155672
R610 VTAIL.n171 VTAIL.n129 0.155672
R611 VTAIL.n163 VTAIL.n129 0.155672
R612 VTAIL.n163 VTAIL.n162 0.155672
R613 VTAIL.n162 VTAIL.n133 0.155672
R614 VTAIL.n155 VTAIL.n133 0.155672
R615 VTAIL.n155 VTAIL.n154 0.155672
R616 VTAIL.n154 VTAIL.n138 0.155672
R617 VTAIL.n147 VTAIL.n138 0.155672
R618 VTAIL.n147 VTAIL.n146 0.155672
R619 VTAIL.n119 VTAIL.n65 0.155672
R620 VTAIL.n112 VTAIL.n65 0.155672
R621 VTAIL.n112 VTAIL.n111 0.155672
R622 VTAIL.n111 VTAIL.n69 0.155672
R623 VTAIL.n103 VTAIL.n69 0.155672
R624 VTAIL.n103 VTAIL.n102 0.155672
R625 VTAIL.n102 VTAIL.n73 0.155672
R626 VTAIL.n95 VTAIL.n73 0.155672
R627 VTAIL.n95 VTAIL.n94 0.155672
R628 VTAIL.n94 VTAIL.n78 0.155672
R629 VTAIL.n87 VTAIL.n78 0.155672
R630 VTAIL.n87 VTAIL.n86 0.155672
R631 B.n673 B.n672 585
R632 B.n673 B.n93 585
R633 B.n676 B.n675 585
R634 B.n677 B.n140 585
R635 B.n679 B.n678 585
R636 B.n681 B.n139 585
R637 B.n684 B.n683 585
R638 B.n685 B.n138 585
R639 B.n687 B.n686 585
R640 B.n689 B.n137 585
R641 B.n692 B.n691 585
R642 B.n693 B.n136 585
R643 B.n695 B.n694 585
R644 B.n697 B.n135 585
R645 B.n700 B.n699 585
R646 B.n701 B.n134 585
R647 B.n703 B.n702 585
R648 B.n705 B.n133 585
R649 B.n708 B.n707 585
R650 B.n709 B.n132 585
R651 B.n711 B.n710 585
R652 B.n713 B.n131 585
R653 B.n716 B.n715 585
R654 B.n717 B.n130 585
R655 B.n719 B.n718 585
R656 B.n721 B.n129 585
R657 B.n724 B.n723 585
R658 B.n725 B.n128 585
R659 B.n727 B.n726 585
R660 B.n729 B.n127 585
R661 B.n732 B.n731 585
R662 B.n733 B.n126 585
R663 B.n735 B.n734 585
R664 B.n737 B.n125 585
R665 B.n740 B.n739 585
R666 B.n741 B.n124 585
R667 B.n743 B.n742 585
R668 B.n745 B.n123 585
R669 B.n748 B.n747 585
R670 B.n750 B.n120 585
R671 B.n752 B.n751 585
R672 B.n754 B.n119 585
R673 B.n757 B.n756 585
R674 B.n758 B.n118 585
R675 B.n760 B.n759 585
R676 B.n762 B.n117 585
R677 B.n764 B.n763 585
R678 B.n766 B.n765 585
R679 B.n769 B.n768 585
R680 B.n770 B.n112 585
R681 B.n772 B.n771 585
R682 B.n774 B.n111 585
R683 B.n777 B.n776 585
R684 B.n778 B.n110 585
R685 B.n780 B.n779 585
R686 B.n782 B.n109 585
R687 B.n785 B.n784 585
R688 B.n786 B.n108 585
R689 B.n788 B.n787 585
R690 B.n790 B.n107 585
R691 B.n793 B.n792 585
R692 B.n794 B.n106 585
R693 B.n796 B.n795 585
R694 B.n798 B.n105 585
R695 B.n801 B.n800 585
R696 B.n802 B.n104 585
R697 B.n804 B.n803 585
R698 B.n806 B.n103 585
R699 B.n809 B.n808 585
R700 B.n810 B.n102 585
R701 B.n812 B.n811 585
R702 B.n814 B.n101 585
R703 B.n817 B.n816 585
R704 B.n818 B.n100 585
R705 B.n820 B.n819 585
R706 B.n822 B.n99 585
R707 B.n825 B.n824 585
R708 B.n826 B.n98 585
R709 B.n828 B.n827 585
R710 B.n830 B.n97 585
R711 B.n833 B.n832 585
R712 B.n834 B.n96 585
R713 B.n836 B.n835 585
R714 B.n838 B.n95 585
R715 B.n841 B.n840 585
R716 B.n842 B.n94 585
R717 B.n671 B.n92 585
R718 B.n845 B.n92 585
R719 B.n670 B.n91 585
R720 B.n846 B.n91 585
R721 B.n669 B.n90 585
R722 B.n847 B.n90 585
R723 B.n668 B.n667 585
R724 B.n667 B.n86 585
R725 B.n666 B.n85 585
R726 B.n853 B.n85 585
R727 B.n665 B.n84 585
R728 B.n854 B.n84 585
R729 B.n664 B.n83 585
R730 B.n855 B.n83 585
R731 B.n663 B.n662 585
R732 B.n662 B.n79 585
R733 B.n661 B.n78 585
R734 B.n861 B.n78 585
R735 B.n660 B.n77 585
R736 B.n862 B.n77 585
R737 B.n659 B.n76 585
R738 B.n863 B.n76 585
R739 B.n658 B.n657 585
R740 B.n657 B.n72 585
R741 B.n656 B.n71 585
R742 B.n869 B.n71 585
R743 B.n655 B.n70 585
R744 B.n870 B.n70 585
R745 B.n654 B.n69 585
R746 B.n871 B.n69 585
R747 B.n653 B.n652 585
R748 B.n652 B.n65 585
R749 B.n651 B.n64 585
R750 B.n877 B.n64 585
R751 B.n650 B.n63 585
R752 B.n878 B.n63 585
R753 B.n649 B.n62 585
R754 B.n879 B.n62 585
R755 B.n648 B.n647 585
R756 B.n647 B.n58 585
R757 B.n646 B.n57 585
R758 B.n885 B.n57 585
R759 B.n645 B.n56 585
R760 B.n886 B.n56 585
R761 B.n644 B.n55 585
R762 B.n887 B.n55 585
R763 B.n643 B.n642 585
R764 B.n642 B.n51 585
R765 B.n641 B.n50 585
R766 B.n893 B.n50 585
R767 B.n640 B.n49 585
R768 B.n894 B.n49 585
R769 B.n639 B.n48 585
R770 B.n895 B.n48 585
R771 B.n638 B.n637 585
R772 B.n637 B.n44 585
R773 B.n636 B.n43 585
R774 B.n901 B.n43 585
R775 B.n635 B.n42 585
R776 B.n902 B.n42 585
R777 B.n634 B.n41 585
R778 B.n903 B.n41 585
R779 B.n633 B.n632 585
R780 B.n632 B.n37 585
R781 B.n631 B.n36 585
R782 B.n909 B.n36 585
R783 B.n630 B.n35 585
R784 B.n910 B.n35 585
R785 B.n629 B.n34 585
R786 B.n911 B.n34 585
R787 B.n628 B.n627 585
R788 B.n627 B.n30 585
R789 B.n626 B.n29 585
R790 B.n917 B.n29 585
R791 B.n625 B.n28 585
R792 B.n918 B.n28 585
R793 B.n624 B.n27 585
R794 B.n919 B.n27 585
R795 B.n623 B.n622 585
R796 B.n622 B.n23 585
R797 B.n621 B.n22 585
R798 B.n925 B.n22 585
R799 B.n620 B.n21 585
R800 B.n926 B.n21 585
R801 B.n619 B.n20 585
R802 B.n927 B.n20 585
R803 B.n618 B.n617 585
R804 B.n617 B.n19 585
R805 B.n616 B.n15 585
R806 B.n933 B.n15 585
R807 B.n615 B.n14 585
R808 B.n934 B.n14 585
R809 B.n614 B.n13 585
R810 B.n935 B.n13 585
R811 B.n613 B.n612 585
R812 B.n612 B.n12 585
R813 B.n611 B.n610 585
R814 B.n611 B.n8 585
R815 B.n609 B.n7 585
R816 B.n942 B.n7 585
R817 B.n608 B.n6 585
R818 B.n943 B.n6 585
R819 B.n607 B.n5 585
R820 B.n944 B.n5 585
R821 B.n606 B.n605 585
R822 B.n605 B.n4 585
R823 B.n604 B.n141 585
R824 B.n604 B.n603 585
R825 B.n594 B.n142 585
R826 B.n143 B.n142 585
R827 B.n596 B.n595 585
R828 B.n597 B.n596 585
R829 B.n593 B.n148 585
R830 B.n148 B.n147 585
R831 B.n592 B.n591 585
R832 B.n591 B.n590 585
R833 B.n150 B.n149 585
R834 B.n583 B.n150 585
R835 B.n582 B.n581 585
R836 B.n584 B.n582 585
R837 B.n580 B.n155 585
R838 B.n155 B.n154 585
R839 B.n579 B.n578 585
R840 B.n578 B.n577 585
R841 B.n157 B.n156 585
R842 B.n158 B.n157 585
R843 B.n570 B.n569 585
R844 B.n571 B.n570 585
R845 B.n568 B.n163 585
R846 B.n163 B.n162 585
R847 B.n567 B.n566 585
R848 B.n566 B.n565 585
R849 B.n165 B.n164 585
R850 B.n166 B.n165 585
R851 B.n558 B.n557 585
R852 B.n559 B.n558 585
R853 B.n556 B.n170 585
R854 B.n174 B.n170 585
R855 B.n555 B.n554 585
R856 B.n554 B.n553 585
R857 B.n172 B.n171 585
R858 B.n173 B.n172 585
R859 B.n546 B.n545 585
R860 B.n547 B.n546 585
R861 B.n544 B.n179 585
R862 B.n179 B.n178 585
R863 B.n543 B.n542 585
R864 B.n542 B.n541 585
R865 B.n181 B.n180 585
R866 B.n182 B.n181 585
R867 B.n534 B.n533 585
R868 B.n535 B.n534 585
R869 B.n532 B.n187 585
R870 B.n187 B.n186 585
R871 B.n531 B.n530 585
R872 B.n530 B.n529 585
R873 B.n189 B.n188 585
R874 B.n190 B.n189 585
R875 B.n522 B.n521 585
R876 B.n523 B.n522 585
R877 B.n520 B.n195 585
R878 B.n195 B.n194 585
R879 B.n519 B.n518 585
R880 B.n518 B.n517 585
R881 B.n197 B.n196 585
R882 B.n198 B.n197 585
R883 B.n510 B.n509 585
R884 B.n511 B.n510 585
R885 B.n508 B.n203 585
R886 B.n203 B.n202 585
R887 B.n507 B.n506 585
R888 B.n506 B.n505 585
R889 B.n205 B.n204 585
R890 B.n206 B.n205 585
R891 B.n498 B.n497 585
R892 B.n499 B.n498 585
R893 B.n496 B.n211 585
R894 B.n211 B.n210 585
R895 B.n495 B.n494 585
R896 B.n494 B.n493 585
R897 B.n213 B.n212 585
R898 B.n214 B.n213 585
R899 B.n486 B.n485 585
R900 B.n487 B.n486 585
R901 B.n484 B.n219 585
R902 B.n219 B.n218 585
R903 B.n483 B.n482 585
R904 B.n482 B.n481 585
R905 B.n221 B.n220 585
R906 B.n222 B.n221 585
R907 B.n474 B.n473 585
R908 B.n475 B.n474 585
R909 B.n472 B.n227 585
R910 B.n227 B.n226 585
R911 B.n471 B.n470 585
R912 B.n470 B.n469 585
R913 B.n229 B.n228 585
R914 B.n230 B.n229 585
R915 B.n462 B.n461 585
R916 B.n463 B.n462 585
R917 B.n460 B.n235 585
R918 B.n235 B.n234 585
R919 B.n459 B.n458 585
R920 B.n458 B.n457 585
R921 B.n454 B.n239 585
R922 B.n453 B.n452 585
R923 B.n450 B.n240 585
R924 B.n450 B.n238 585
R925 B.n449 B.n448 585
R926 B.n447 B.n446 585
R927 B.n445 B.n242 585
R928 B.n443 B.n442 585
R929 B.n441 B.n243 585
R930 B.n440 B.n439 585
R931 B.n437 B.n244 585
R932 B.n435 B.n434 585
R933 B.n433 B.n245 585
R934 B.n432 B.n431 585
R935 B.n429 B.n246 585
R936 B.n427 B.n426 585
R937 B.n425 B.n247 585
R938 B.n424 B.n423 585
R939 B.n421 B.n248 585
R940 B.n419 B.n418 585
R941 B.n417 B.n249 585
R942 B.n416 B.n415 585
R943 B.n413 B.n250 585
R944 B.n411 B.n410 585
R945 B.n409 B.n251 585
R946 B.n408 B.n407 585
R947 B.n405 B.n252 585
R948 B.n403 B.n402 585
R949 B.n401 B.n253 585
R950 B.n400 B.n399 585
R951 B.n397 B.n254 585
R952 B.n395 B.n394 585
R953 B.n393 B.n255 585
R954 B.n392 B.n391 585
R955 B.n389 B.n256 585
R956 B.n387 B.n386 585
R957 B.n385 B.n257 585
R958 B.n384 B.n383 585
R959 B.n381 B.n258 585
R960 B.n379 B.n378 585
R961 B.n377 B.n259 585
R962 B.n376 B.n375 585
R963 B.n373 B.n263 585
R964 B.n371 B.n370 585
R965 B.n369 B.n264 585
R966 B.n368 B.n367 585
R967 B.n365 B.n265 585
R968 B.n363 B.n362 585
R969 B.n360 B.n266 585
R970 B.n359 B.n358 585
R971 B.n356 B.n269 585
R972 B.n354 B.n353 585
R973 B.n352 B.n270 585
R974 B.n351 B.n350 585
R975 B.n348 B.n271 585
R976 B.n346 B.n345 585
R977 B.n344 B.n272 585
R978 B.n343 B.n342 585
R979 B.n340 B.n273 585
R980 B.n338 B.n337 585
R981 B.n336 B.n274 585
R982 B.n335 B.n334 585
R983 B.n332 B.n275 585
R984 B.n330 B.n329 585
R985 B.n328 B.n276 585
R986 B.n327 B.n326 585
R987 B.n324 B.n277 585
R988 B.n322 B.n321 585
R989 B.n320 B.n278 585
R990 B.n319 B.n318 585
R991 B.n316 B.n279 585
R992 B.n314 B.n313 585
R993 B.n312 B.n280 585
R994 B.n311 B.n310 585
R995 B.n308 B.n281 585
R996 B.n306 B.n305 585
R997 B.n304 B.n282 585
R998 B.n303 B.n302 585
R999 B.n300 B.n283 585
R1000 B.n298 B.n297 585
R1001 B.n296 B.n284 585
R1002 B.n295 B.n294 585
R1003 B.n292 B.n285 585
R1004 B.n290 B.n289 585
R1005 B.n288 B.n287 585
R1006 B.n237 B.n236 585
R1007 B.n456 B.n455 585
R1008 B.n457 B.n456 585
R1009 B.n233 B.n232 585
R1010 B.n234 B.n233 585
R1011 B.n465 B.n464 585
R1012 B.n464 B.n463 585
R1013 B.n466 B.n231 585
R1014 B.n231 B.n230 585
R1015 B.n468 B.n467 585
R1016 B.n469 B.n468 585
R1017 B.n225 B.n224 585
R1018 B.n226 B.n225 585
R1019 B.n477 B.n476 585
R1020 B.n476 B.n475 585
R1021 B.n478 B.n223 585
R1022 B.n223 B.n222 585
R1023 B.n480 B.n479 585
R1024 B.n481 B.n480 585
R1025 B.n217 B.n216 585
R1026 B.n218 B.n217 585
R1027 B.n489 B.n488 585
R1028 B.n488 B.n487 585
R1029 B.n490 B.n215 585
R1030 B.n215 B.n214 585
R1031 B.n492 B.n491 585
R1032 B.n493 B.n492 585
R1033 B.n209 B.n208 585
R1034 B.n210 B.n209 585
R1035 B.n501 B.n500 585
R1036 B.n500 B.n499 585
R1037 B.n502 B.n207 585
R1038 B.n207 B.n206 585
R1039 B.n504 B.n503 585
R1040 B.n505 B.n504 585
R1041 B.n201 B.n200 585
R1042 B.n202 B.n201 585
R1043 B.n513 B.n512 585
R1044 B.n512 B.n511 585
R1045 B.n514 B.n199 585
R1046 B.n199 B.n198 585
R1047 B.n516 B.n515 585
R1048 B.n517 B.n516 585
R1049 B.n193 B.n192 585
R1050 B.n194 B.n193 585
R1051 B.n525 B.n524 585
R1052 B.n524 B.n523 585
R1053 B.n526 B.n191 585
R1054 B.n191 B.n190 585
R1055 B.n528 B.n527 585
R1056 B.n529 B.n528 585
R1057 B.n185 B.n184 585
R1058 B.n186 B.n185 585
R1059 B.n537 B.n536 585
R1060 B.n536 B.n535 585
R1061 B.n538 B.n183 585
R1062 B.n183 B.n182 585
R1063 B.n540 B.n539 585
R1064 B.n541 B.n540 585
R1065 B.n177 B.n176 585
R1066 B.n178 B.n177 585
R1067 B.n549 B.n548 585
R1068 B.n548 B.n547 585
R1069 B.n550 B.n175 585
R1070 B.n175 B.n173 585
R1071 B.n552 B.n551 585
R1072 B.n553 B.n552 585
R1073 B.n169 B.n168 585
R1074 B.n174 B.n169 585
R1075 B.n561 B.n560 585
R1076 B.n560 B.n559 585
R1077 B.n562 B.n167 585
R1078 B.n167 B.n166 585
R1079 B.n564 B.n563 585
R1080 B.n565 B.n564 585
R1081 B.n161 B.n160 585
R1082 B.n162 B.n161 585
R1083 B.n573 B.n572 585
R1084 B.n572 B.n571 585
R1085 B.n574 B.n159 585
R1086 B.n159 B.n158 585
R1087 B.n576 B.n575 585
R1088 B.n577 B.n576 585
R1089 B.n153 B.n152 585
R1090 B.n154 B.n153 585
R1091 B.n586 B.n585 585
R1092 B.n585 B.n584 585
R1093 B.n587 B.n151 585
R1094 B.n583 B.n151 585
R1095 B.n589 B.n588 585
R1096 B.n590 B.n589 585
R1097 B.n146 B.n145 585
R1098 B.n147 B.n146 585
R1099 B.n599 B.n598 585
R1100 B.n598 B.n597 585
R1101 B.n600 B.n144 585
R1102 B.n144 B.n143 585
R1103 B.n602 B.n601 585
R1104 B.n603 B.n602 585
R1105 B.n3 B.n0 585
R1106 B.n4 B.n3 585
R1107 B.n941 B.n1 585
R1108 B.n942 B.n941 585
R1109 B.n940 B.n939 585
R1110 B.n940 B.n8 585
R1111 B.n938 B.n9 585
R1112 B.n12 B.n9 585
R1113 B.n937 B.n936 585
R1114 B.n936 B.n935 585
R1115 B.n11 B.n10 585
R1116 B.n934 B.n11 585
R1117 B.n932 B.n931 585
R1118 B.n933 B.n932 585
R1119 B.n930 B.n16 585
R1120 B.n19 B.n16 585
R1121 B.n929 B.n928 585
R1122 B.n928 B.n927 585
R1123 B.n18 B.n17 585
R1124 B.n926 B.n18 585
R1125 B.n924 B.n923 585
R1126 B.n925 B.n924 585
R1127 B.n922 B.n24 585
R1128 B.n24 B.n23 585
R1129 B.n921 B.n920 585
R1130 B.n920 B.n919 585
R1131 B.n26 B.n25 585
R1132 B.n918 B.n26 585
R1133 B.n916 B.n915 585
R1134 B.n917 B.n916 585
R1135 B.n914 B.n31 585
R1136 B.n31 B.n30 585
R1137 B.n913 B.n912 585
R1138 B.n912 B.n911 585
R1139 B.n33 B.n32 585
R1140 B.n910 B.n33 585
R1141 B.n908 B.n907 585
R1142 B.n909 B.n908 585
R1143 B.n906 B.n38 585
R1144 B.n38 B.n37 585
R1145 B.n905 B.n904 585
R1146 B.n904 B.n903 585
R1147 B.n40 B.n39 585
R1148 B.n902 B.n40 585
R1149 B.n900 B.n899 585
R1150 B.n901 B.n900 585
R1151 B.n898 B.n45 585
R1152 B.n45 B.n44 585
R1153 B.n897 B.n896 585
R1154 B.n896 B.n895 585
R1155 B.n47 B.n46 585
R1156 B.n894 B.n47 585
R1157 B.n892 B.n891 585
R1158 B.n893 B.n892 585
R1159 B.n890 B.n52 585
R1160 B.n52 B.n51 585
R1161 B.n889 B.n888 585
R1162 B.n888 B.n887 585
R1163 B.n54 B.n53 585
R1164 B.n886 B.n54 585
R1165 B.n884 B.n883 585
R1166 B.n885 B.n884 585
R1167 B.n882 B.n59 585
R1168 B.n59 B.n58 585
R1169 B.n881 B.n880 585
R1170 B.n880 B.n879 585
R1171 B.n61 B.n60 585
R1172 B.n878 B.n61 585
R1173 B.n876 B.n875 585
R1174 B.n877 B.n876 585
R1175 B.n874 B.n66 585
R1176 B.n66 B.n65 585
R1177 B.n873 B.n872 585
R1178 B.n872 B.n871 585
R1179 B.n68 B.n67 585
R1180 B.n870 B.n68 585
R1181 B.n868 B.n867 585
R1182 B.n869 B.n868 585
R1183 B.n866 B.n73 585
R1184 B.n73 B.n72 585
R1185 B.n865 B.n864 585
R1186 B.n864 B.n863 585
R1187 B.n75 B.n74 585
R1188 B.n862 B.n75 585
R1189 B.n860 B.n859 585
R1190 B.n861 B.n860 585
R1191 B.n858 B.n80 585
R1192 B.n80 B.n79 585
R1193 B.n857 B.n856 585
R1194 B.n856 B.n855 585
R1195 B.n82 B.n81 585
R1196 B.n854 B.n82 585
R1197 B.n852 B.n851 585
R1198 B.n853 B.n852 585
R1199 B.n850 B.n87 585
R1200 B.n87 B.n86 585
R1201 B.n849 B.n848 585
R1202 B.n848 B.n847 585
R1203 B.n89 B.n88 585
R1204 B.n846 B.n89 585
R1205 B.n844 B.n843 585
R1206 B.n845 B.n844 585
R1207 B.n945 B.n944 585
R1208 B.n943 B.n2 585
R1209 B.n844 B.n94 516.524
R1210 B.n673 B.n92 516.524
R1211 B.n458 B.n237 516.524
R1212 B.n456 B.n239 516.524
R1213 B.n121 B.t14 330.536
R1214 B.n267 B.t11 330.536
R1215 B.n113 B.t17 330.534
R1216 B.n260 B.t8 330.534
R1217 B.n113 B.t16 288.409
R1218 B.n121 B.t12 288.409
R1219 B.n267 B.t9 288.409
R1220 B.n260 B.t5 288.409
R1221 B.n122 B.t15 260.911
R1222 B.n268 B.t10 260.911
R1223 B.n114 B.t18 260.911
R1224 B.n261 B.t7 260.911
R1225 B.n674 B.n93 256.663
R1226 B.n680 B.n93 256.663
R1227 B.n682 B.n93 256.663
R1228 B.n688 B.n93 256.663
R1229 B.n690 B.n93 256.663
R1230 B.n696 B.n93 256.663
R1231 B.n698 B.n93 256.663
R1232 B.n704 B.n93 256.663
R1233 B.n706 B.n93 256.663
R1234 B.n712 B.n93 256.663
R1235 B.n714 B.n93 256.663
R1236 B.n720 B.n93 256.663
R1237 B.n722 B.n93 256.663
R1238 B.n728 B.n93 256.663
R1239 B.n730 B.n93 256.663
R1240 B.n736 B.n93 256.663
R1241 B.n738 B.n93 256.663
R1242 B.n744 B.n93 256.663
R1243 B.n746 B.n93 256.663
R1244 B.n753 B.n93 256.663
R1245 B.n755 B.n93 256.663
R1246 B.n761 B.n93 256.663
R1247 B.n116 B.n93 256.663
R1248 B.n767 B.n93 256.663
R1249 B.n773 B.n93 256.663
R1250 B.n775 B.n93 256.663
R1251 B.n781 B.n93 256.663
R1252 B.n783 B.n93 256.663
R1253 B.n789 B.n93 256.663
R1254 B.n791 B.n93 256.663
R1255 B.n797 B.n93 256.663
R1256 B.n799 B.n93 256.663
R1257 B.n805 B.n93 256.663
R1258 B.n807 B.n93 256.663
R1259 B.n813 B.n93 256.663
R1260 B.n815 B.n93 256.663
R1261 B.n821 B.n93 256.663
R1262 B.n823 B.n93 256.663
R1263 B.n829 B.n93 256.663
R1264 B.n831 B.n93 256.663
R1265 B.n837 B.n93 256.663
R1266 B.n839 B.n93 256.663
R1267 B.n451 B.n238 256.663
R1268 B.n241 B.n238 256.663
R1269 B.n444 B.n238 256.663
R1270 B.n438 B.n238 256.663
R1271 B.n436 B.n238 256.663
R1272 B.n430 B.n238 256.663
R1273 B.n428 B.n238 256.663
R1274 B.n422 B.n238 256.663
R1275 B.n420 B.n238 256.663
R1276 B.n414 B.n238 256.663
R1277 B.n412 B.n238 256.663
R1278 B.n406 B.n238 256.663
R1279 B.n404 B.n238 256.663
R1280 B.n398 B.n238 256.663
R1281 B.n396 B.n238 256.663
R1282 B.n390 B.n238 256.663
R1283 B.n388 B.n238 256.663
R1284 B.n382 B.n238 256.663
R1285 B.n380 B.n238 256.663
R1286 B.n374 B.n238 256.663
R1287 B.n372 B.n238 256.663
R1288 B.n366 B.n238 256.663
R1289 B.n364 B.n238 256.663
R1290 B.n357 B.n238 256.663
R1291 B.n355 B.n238 256.663
R1292 B.n349 B.n238 256.663
R1293 B.n347 B.n238 256.663
R1294 B.n341 B.n238 256.663
R1295 B.n339 B.n238 256.663
R1296 B.n333 B.n238 256.663
R1297 B.n331 B.n238 256.663
R1298 B.n325 B.n238 256.663
R1299 B.n323 B.n238 256.663
R1300 B.n317 B.n238 256.663
R1301 B.n315 B.n238 256.663
R1302 B.n309 B.n238 256.663
R1303 B.n307 B.n238 256.663
R1304 B.n301 B.n238 256.663
R1305 B.n299 B.n238 256.663
R1306 B.n293 B.n238 256.663
R1307 B.n291 B.n238 256.663
R1308 B.n286 B.n238 256.663
R1309 B.n947 B.n946 256.663
R1310 B.n840 B.n838 163.367
R1311 B.n836 B.n96 163.367
R1312 B.n832 B.n830 163.367
R1313 B.n828 B.n98 163.367
R1314 B.n824 B.n822 163.367
R1315 B.n820 B.n100 163.367
R1316 B.n816 B.n814 163.367
R1317 B.n812 B.n102 163.367
R1318 B.n808 B.n806 163.367
R1319 B.n804 B.n104 163.367
R1320 B.n800 B.n798 163.367
R1321 B.n796 B.n106 163.367
R1322 B.n792 B.n790 163.367
R1323 B.n788 B.n108 163.367
R1324 B.n784 B.n782 163.367
R1325 B.n780 B.n110 163.367
R1326 B.n776 B.n774 163.367
R1327 B.n772 B.n112 163.367
R1328 B.n768 B.n766 163.367
R1329 B.n763 B.n762 163.367
R1330 B.n760 B.n118 163.367
R1331 B.n756 B.n754 163.367
R1332 B.n752 B.n120 163.367
R1333 B.n747 B.n745 163.367
R1334 B.n743 B.n124 163.367
R1335 B.n739 B.n737 163.367
R1336 B.n735 B.n126 163.367
R1337 B.n731 B.n729 163.367
R1338 B.n727 B.n128 163.367
R1339 B.n723 B.n721 163.367
R1340 B.n719 B.n130 163.367
R1341 B.n715 B.n713 163.367
R1342 B.n711 B.n132 163.367
R1343 B.n707 B.n705 163.367
R1344 B.n703 B.n134 163.367
R1345 B.n699 B.n697 163.367
R1346 B.n695 B.n136 163.367
R1347 B.n691 B.n689 163.367
R1348 B.n687 B.n138 163.367
R1349 B.n683 B.n681 163.367
R1350 B.n679 B.n140 163.367
R1351 B.n675 B.n673 163.367
R1352 B.n458 B.n235 163.367
R1353 B.n462 B.n235 163.367
R1354 B.n462 B.n229 163.367
R1355 B.n470 B.n229 163.367
R1356 B.n470 B.n227 163.367
R1357 B.n474 B.n227 163.367
R1358 B.n474 B.n221 163.367
R1359 B.n482 B.n221 163.367
R1360 B.n482 B.n219 163.367
R1361 B.n486 B.n219 163.367
R1362 B.n486 B.n213 163.367
R1363 B.n494 B.n213 163.367
R1364 B.n494 B.n211 163.367
R1365 B.n498 B.n211 163.367
R1366 B.n498 B.n205 163.367
R1367 B.n506 B.n205 163.367
R1368 B.n506 B.n203 163.367
R1369 B.n510 B.n203 163.367
R1370 B.n510 B.n197 163.367
R1371 B.n518 B.n197 163.367
R1372 B.n518 B.n195 163.367
R1373 B.n522 B.n195 163.367
R1374 B.n522 B.n189 163.367
R1375 B.n530 B.n189 163.367
R1376 B.n530 B.n187 163.367
R1377 B.n534 B.n187 163.367
R1378 B.n534 B.n181 163.367
R1379 B.n542 B.n181 163.367
R1380 B.n542 B.n179 163.367
R1381 B.n546 B.n179 163.367
R1382 B.n546 B.n172 163.367
R1383 B.n554 B.n172 163.367
R1384 B.n554 B.n170 163.367
R1385 B.n558 B.n170 163.367
R1386 B.n558 B.n165 163.367
R1387 B.n566 B.n165 163.367
R1388 B.n566 B.n163 163.367
R1389 B.n570 B.n163 163.367
R1390 B.n570 B.n157 163.367
R1391 B.n578 B.n157 163.367
R1392 B.n578 B.n155 163.367
R1393 B.n582 B.n155 163.367
R1394 B.n582 B.n150 163.367
R1395 B.n591 B.n150 163.367
R1396 B.n591 B.n148 163.367
R1397 B.n596 B.n148 163.367
R1398 B.n596 B.n142 163.367
R1399 B.n604 B.n142 163.367
R1400 B.n605 B.n604 163.367
R1401 B.n605 B.n5 163.367
R1402 B.n6 B.n5 163.367
R1403 B.n7 B.n6 163.367
R1404 B.n611 B.n7 163.367
R1405 B.n612 B.n611 163.367
R1406 B.n612 B.n13 163.367
R1407 B.n14 B.n13 163.367
R1408 B.n15 B.n14 163.367
R1409 B.n617 B.n15 163.367
R1410 B.n617 B.n20 163.367
R1411 B.n21 B.n20 163.367
R1412 B.n22 B.n21 163.367
R1413 B.n622 B.n22 163.367
R1414 B.n622 B.n27 163.367
R1415 B.n28 B.n27 163.367
R1416 B.n29 B.n28 163.367
R1417 B.n627 B.n29 163.367
R1418 B.n627 B.n34 163.367
R1419 B.n35 B.n34 163.367
R1420 B.n36 B.n35 163.367
R1421 B.n632 B.n36 163.367
R1422 B.n632 B.n41 163.367
R1423 B.n42 B.n41 163.367
R1424 B.n43 B.n42 163.367
R1425 B.n637 B.n43 163.367
R1426 B.n637 B.n48 163.367
R1427 B.n49 B.n48 163.367
R1428 B.n50 B.n49 163.367
R1429 B.n642 B.n50 163.367
R1430 B.n642 B.n55 163.367
R1431 B.n56 B.n55 163.367
R1432 B.n57 B.n56 163.367
R1433 B.n647 B.n57 163.367
R1434 B.n647 B.n62 163.367
R1435 B.n63 B.n62 163.367
R1436 B.n64 B.n63 163.367
R1437 B.n652 B.n64 163.367
R1438 B.n652 B.n69 163.367
R1439 B.n70 B.n69 163.367
R1440 B.n71 B.n70 163.367
R1441 B.n657 B.n71 163.367
R1442 B.n657 B.n76 163.367
R1443 B.n77 B.n76 163.367
R1444 B.n78 B.n77 163.367
R1445 B.n662 B.n78 163.367
R1446 B.n662 B.n83 163.367
R1447 B.n84 B.n83 163.367
R1448 B.n85 B.n84 163.367
R1449 B.n667 B.n85 163.367
R1450 B.n667 B.n90 163.367
R1451 B.n91 B.n90 163.367
R1452 B.n92 B.n91 163.367
R1453 B.n452 B.n450 163.367
R1454 B.n450 B.n449 163.367
R1455 B.n446 B.n445 163.367
R1456 B.n443 B.n243 163.367
R1457 B.n439 B.n437 163.367
R1458 B.n435 B.n245 163.367
R1459 B.n431 B.n429 163.367
R1460 B.n427 B.n247 163.367
R1461 B.n423 B.n421 163.367
R1462 B.n419 B.n249 163.367
R1463 B.n415 B.n413 163.367
R1464 B.n411 B.n251 163.367
R1465 B.n407 B.n405 163.367
R1466 B.n403 B.n253 163.367
R1467 B.n399 B.n397 163.367
R1468 B.n395 B.n255 163.367
R1469 B.n391 B.n389 163.367
R1470 B.n387 B.n257 163.367
R1471 B.n383 B.n381 163.367
R1472 B.n379 B.n259 163.367
R1473 B.n375 B.n373 163.367
R1474 B.n371 B.n264 163.367
R1475 B.n367 B.n365 163.367
R1476 B.n363 B.n266 163.367
R1477 B.n358 B.n356 163.367
R1478 B.n354 B.n270 163.367
R1479 B.n350 B.n348 163.367
R1480 B.n346 B.n272 163.367
R1481 B.n342 B.n340 163.367
R1482 B.n338 B.n274 163.367
R1483 B.n334 B.n332 163.367
R1484 B.n330 B.n276 163.367
R1485 B.n326 B.n324 163.367
R1486 B.n322 B.n278 163.367
R1487 B.n318 B.n316 163.367
R1488 B.n314 B.n280 163.367
R1489 B.n310 B.n308 163.367
R1490 B.n306 B.n282 163.367
R1491 B.n302 B.n300 163.367
R1492 B.n298 B.n284 163.367
R1493 B.n294 B.n292 163.367
R1494 B.n290 B.n287 163.367
R1495 B.n456 B.n233 163.367
R1496 B.n464 B.n233 163.367
R1497 B.n464 B.n231 163.367
R1498 B.n468 B.n231 163.367
R1499 B.n468 B.n225 163.367
R1500 B.n476 B.n225 163.367
R1501 B.n476 B.n223 163.367
R1502 B.n480 B.n223 163.367
R1503 B.n480 B.n217 163.367
R1504 B.n488 B.n217 163.367
R1505 B.n488 B.n215 163.367
R1506 B.n492 B.n215 163.367
R1507 B.n492 B.n209 163.367
R1508 B.n500 B.n209 163.367
R1509 B.n500 B.n207 163.367
R1510 B.n504 B.n207 163.367
R1511 B.n504 B.n201 163.367
R1512 B.n512 B.n201 163.367
R1513 B.n512 B.n199 163.367
R1514 B.n516 B.n199 163.367
R1515 B.n516 B.n193 163.367
R1516 B.n524 B.n193 163.367
R1517 B.n524 B.n191 163.367
R1518 B.n528 B.n191 163.367
R1519 B.n528 B.n185 163.367
R1520 B.n536 B.n185 163.367
R1521 B.n536 B.n183 163.367
R1522 B.n540 B.n183 163.367
R1523 B.n540 B.n177 163.367
R1524 B.n548 B.n177 163.367
R1525 B.n548 B.n175 163.367
R1526 B.n552 B.n175 163.367
R1527 B.n552 B.n169 163.367
R1528 B.n560 B.n169 163.367
R1529 B.n560 B.n167 163.367
R1530 B.n564 B.n167 163.367
R1531 B.n564 B.n161 163.367
R1532 B.n572 B.n161 163.367
R1533 B.n572 B.n159 163.367
R1534 B.n576 B.n159 163.367
R1535 B.n576 B.n153 163.367
R1536 B.n585 B.n153 163.367
R1537 B.n585 B.n151 163.367
R1538 B.n589 B.n151 163.367
R1539 B.n589 B.n146 163.367
R1540 B.n598 B.n146 163.367
R1541 B.n598 B.n144 163.367
R1542 B.n602 B.n144 163.367
R1543 B.n602 B.n3 163.367
R1544 B.n945 B.n3 163.367
R1545 B.n941 B.n2 163.367
R1546 B.n941 B.n940 163.367
R1547 B.n940 B.n9 163.367
R1548 B.n936 B.n9 163.367
R1549 B.n936 B.n11 163.367
R1550 B.n932 B.n11 163.367
R1551 B.n932 B.n16 163.367
R1552 B.n928 B.n16 163.367
R1553 B.n928 B.n18 163.367
R1554 B.n924 B.n18 163.367
R1555 B.n924 B.n24 163.367
R1556 B.n920 B.n24 163.367
R1557 B.n920 B.n26 163.367
R1558 B.n916 B.n26 163.367
R1559 B.n916 B.n31 163.367
R1560 B.n912 B.n31 163.367
R1561 B.n912 B.n33 163.367
R1562 B.n908 B.n33 163.367
R1563 B.n908 B.n38 163.367
R1564 B.n904 B.n38 163.367
R1565 B.n904 B.n40 163.367
R1566 B.n900 B.n40 163.367
R1567 B.n900 B.n45 163.367
R1568 B.n896 B.n45 163.367
R1569 B.n896 B.n47 163.367
R1570 B.n892 B.n47 163.367
R1571 B.n892 B.n52 163.367
R1572 B.n888 B.n52 163.367
R1573 B.n888 B.n54 163.367
R1574 B.n884 B.n54 163.367
R1575 B.n884 B.n59 163.367
R1576 B.n880 B.n59 163.367
R1577 B.n880 B.n61 163.367
R1578 B.n876 B.n61 163.367
R1579 B.n876 B.n66 163.367
R1580 B.n872 B.n66 163.367
R1581 B.n872 B.n68 163.367
R1582 B.n868 B.n68 163.367
R1583 B.n868 B.n73 163.367
R1584 B.n864 B.n73 163.367
R1585 B.n864 B.n75 163.367
R1586 B.n860 B.n75 163.367
R1587 B.n860 B.n80 163.367
R1588 B.n856 B.n80 163.367
R1589 B.n856 B.n82 163.367
R1590 B.n852 B.n82 163.367
R1591 B.n852 B.n87 163.367
R1592 B.n848 B.n87 163.367
R1593 B.n848 B.n89 163.367
R1594 B.n844 B.n89 163.367
R1595 B.n457 B.n238 77.5184
R1596 B.n845 B.n93 77.5184
R1597 B.n839 B.n94 71.676
R1598 B.n838 B.n837 71.676
R1599 B.n831 B.n96 71.676
R1600 B.n830 B.n829 71.676
R1601 B.n823 B.n98 71.676
R1602 B.n822 B.n821 71.676
R1603 B.n815 B.n100 71.676
R1604 B.n814 B.n813 71.676
R1605 B.n807 B.n102 71.676
R1606 B.n806 B.n805 71.676
R1607 B.n799 B.n104 71.676
R1608 B.n798 B.n797 71.676
R1609 B.n791 B.n106 71.676
R1610 B.n790 B.n789 71.676
R1611 B.n783 B.n108 71.676
R1612 B.n782 B.n781 71.676
R1613 B.n775 B.n110 71.676
R1614 B.n774 B.n773 71.676
R1615 B.n767 B.n112 71.676
R1616 B.n766 B.n116 71.676
R1617 B.n762 B.n761 71.676
R1618 B.n755 B.n118 71.676
R1619 B.n754 B.n753 71.676
R1620 B.n746 B.n120 71.676
R1621 B.n745 B.n744 71.676
R1622 B.n738 B.n124 71.676
R1623 B.n737 B.n736 71.676
R1624 B.n730 B.n126 71.676
R1625 B.n729 B.n728 71.676
R1626 B.n722 B.n128 71.676
R1627 B.n721 B.n720 71.676
R1628 B.n714 B.n130 71.676
R1629 B.n713 B.n712 71.676
R1630 B.n706 B.n132 71.676
R1631 B.n705 B.n704 71.676
R1632 B.n698 B.n134 71.676
R1633 B.n697 B.n696 71.676
R1634 B.n690 B.n136 71.676
R1635 B.n689 B.n688 71.676
R1636 B.n682 B.n138 71.676
R1637 B.n681 B.n680 71.676
R1638 B.n674 B.n140 71.676
R1639 B.n675 B.n674 71.676
R1640 B.n680 B.n679 71.676
R1641 B.n683 B.n682 71.676
R1642 B.n688 B.n687 71.676
R1643 B.n691 B.n690 71.676
R1644 B.n696 B.n695 71.676
R1645 B.n699 B.n698 71.676
R1646 B.n704 B.n703 71.676
R1647 B.n707 B.n706 71.676
R1648 B.n712 B.n711 71.676
R1649 B.n715 B.n714 71.676
R1650 B.n720 B.n719 71.676
R1651 B.n723 B.n722 71.676
R1652 B.n728 B.n727 71.676
R1653 B.n731 B.n730 71.676
R1654 B.n736 B.n735 71.676
R1655 B.n739 B.n738 71.676
R1656 B.n744 B.n743 71.676
R1657 B.n747 B.n746 71.676
R1658 B.n753 B.n752 71.676
R1659 B.n756 B.n755 71.676
R1660 B.n761 B.n760 71.676
R1661 B.n763 B.n116 71.676
R1662 B.n768 B.n767 71.676
R1663 B.n773 B.n772 71.676
R1664 B.n776 B.n775 71.676
R1665 B.n781 B.n780 71.676
R1666 B.n784 B.n783 71.676
R1667 B.n789 B.n788 71.676
R1668 B.n792 B.n791 71.676
R1669 B.n797 B.n796 71.676
R1670 B.n800 B.n799 71.676
R1671 B.n805 B.n804 71.676
R1672 B.n808 B.n807 71.676
R1673 B.n813 B.n812 71.676
R1674 B.n816 B.n815 71.676
R1675 B.n821 B.n820 71.676
R1676 B.n824 B.n823 71.676
R1677 B.n829 B.n828 71.676
R1678 B.n832 B.n831 71.676
R1679 B.n837 B.n836 71.676
R1680 B.n840 B.n839 71.676
R1681 B.n451 B.n239 71.676
R1682 B.n449 B.n241 71.676
R1683 B.n445 B.n444 71.676
R1684 B.n438 B.n243 71.676
R1685 B.n437 B.n436 71.676
R1686 B.n430 B.n245 71.676
R1687 B.n429 B.n428 71.676
R1688 B.n422 B.n247 71.676
R1689 B.n421 B.n420 71.676
R1690 B.n414 B.n249 71.676
R1691 B.n413 B.n412 71.676
R1692 B.n406 B.n251 71.676
R1693 B.n405 B.n404 71.676
R1694 B.n398 B.n253 71.676
R1695 B.n397 B.n396 71.676
R1696 B.n390 B.n255 71.676
R1697 B.n389 B.n388 71.676
R1698 B.n382 B.n257 71.676
R1699 B.n381 B.n380 71.676
R1700 B.n374 B.n259 71.676
R1701 B.n373 B.n372 71.676
R1702 B.n366 B.n264 71.676
R1703 B.n365 B.n364 71.676
R1704 B.n357 B.n266 71.676
R1705 B.n356 B.n355 71.676
R1706 B.n349 B.n270 71.676
R1707 B.n348 B.n347 71.676
R1708 B.n341 B.n272 71.676
R1709 B.n340 B.n339 71.676
R1710 B.n333 B.n274 71.676
R1711 B.n332 B.n331 71.676
R1712 B.n325 B.n276 71.676
R1713 B.n324 B.n323 71.676
R1714 B.n317 B.n278 71.676
R1715 B.n316 B.n315 71.676
R1716 B.n309 B.n280 71.676
R1717 B.n308 B.n307 71.676
R1718 B.n301 B.n282 71.676
R1719 B.n300 B.n299 71.676
R1720 B.n293 B.n284 71.676
R1721 B.n292 B.n291 71.676
R1722 B.n287 B.n286 71.676
R1723 B.n452 B.n451 71.676
R1724 B.n446 B.n241 71.676
R1725 B.n444 B.n443 71.676
R1726 B.n439 B.n438 71.676
R1727 B.n436 B.n435 71.676
R1728 B.n431 B.n430 71.676
R1729 B.n428 B.n427 71.676
R1730 B.n423 B.n422 71.676
R1731 B.n420 B.n419 71.676
R1732 B.n415 B.n414 71.676
R1733 B.n412 B.n411 71.676
R1734 B.n407 B.n406 71.676
R1735 B.n404 B.n403 71.676
R1736 B.n399 B.n398 71.676
R1737 B.n396 B.n395 71.676
R1738 B.n391 B.n390 71.676
R1739 B.n388 B.n387 71.676
R1740 B.n383 B.n382 71.676
R1741 B.n380 B.n379 71.676
R1742 B.n375 B.n374 71.676
R1743 B.n372 B.n371 71.676
R1744 B.n367 B.n366 71.676
R1745 B.n364 B.n363 71.676
R1746 B.n358 B.n357 71.676
R1747 B.n355 B.n354 71.676
R1748 B.n350 B.n349 71.676
R1749 B.n347 B.n346 71.676
R1750 B.n342 B.n341 71.676
R1751 B.n339 B.n338 71.676
R1752 B.n334 B.n333 71.676
R1753 B.n331 B.n330 71.676
R1754 B.n326 B.n325 71.676
R1755 B.n323 B.n322 71.676
R1756 B.n318 B.n317 71.676
R1757 B.n315 B.n314 71.676
R1758 B.n310 B.n309 71.676
R1759 B.n307 B.n306 71.676
R1760 B.n302 B.n301 71.676
R1761 B.n299 B.n298 71.676
R1762 B.n294 B.n293 71.676
R1763 B.n291 B.n290 71.676
R1764 B.n286 B.n237 71.676
R1765 B.n946 B.n945 71.676
R1766 B.n946 B.n2 71.676
R1767 B.n114 B.n113 69.6247
R1768 B.n122 B.n121 69.6247
R1769 B.n268 B.n267 69.6247
R1770 B.n261 B.n260 69.6247
R1771 B.n115 B.n114 59.5399
R1772 B.n749 B.n122 59.5399
R1773 B.n361 B.n268 59.5399
R1774 B.n262 B.n261 59.5399
R1775 B.n457 B.n234 46.6485
R1776 B.n463 B.n234 46.6485
R1777 B.n463 B.n230 46.6485
R1778 B.n469 B.n230 46.6485
R1779 B.n469 B.n226 46.6485
R1780 B.n475 B.n226 46.6485
R1781 B.n475 B.n222 46.6485
R1782 B.n481 B.n222 46.6485
R1783 B.n487 B.n218 46.6485
R1784 B.n487 B.n214 46.6485
R1785 B.n493 B.n214 46.6485
R1786 B.n493 B.n210 46.6485
R1787 B.n499 B.n210 46.6485
R1788 B.n499 B.n206 46.6485
R1789 B.n505 B.n206 46.6485
R1790 B.n505 B.n202 46.6485
R1791 B.n511 B.n202 46.6485
R1792 B.n511 B.n198 46.6485
R1793 B.n517 B.n198 46.6485
R1794 B.n517 B.n194 46.6485
R1795 B.n523 B.n194 46.6485
R1796 B.n529 B.n190 46.6485
R1797 B.n529 B.n186 46.6485
R1798 B.n535 B.n186 46.6485
R1799 B.n535 B.n182 46.6485
R1800 B.n541 B.n182 46.6485
R1801 B.n541 B.n178 46.6485
R1802 B.n547 B.n178 46.6485
R1803 B.n547 B.n173 46.6485
R1804 B.n553 B.n173 46.6485
R1805 B.n553 B.n174 46.6485
R1806 B.n559 B.n166 46.6485
R1807 B.n565 B.n166 46.6485
R1808 B.n565 B.n162 46.6485
R1809 B.n571 B.n162 46.6485
R1810 B.n571 B.n158 46.6485
R1811 B.n577 B.n158 46.6485
R1812 B.n577 B.n154 46.6485
R1813 B.n584 B.n154 46.6485
R1814 B.n584 B.n583 46.6485
R1815 B.n590 B.n147 46.6485
R1816 B.n597 B.n147 46.6485
R1817 B.n597 B.n143 46.6485
R1818 B.n603 B.n143 46.6485
R1819 B.n603 B.n4 46.6485
R1820 B.n944 B.n4 46.6485
R1821 B.n944 B.n943 46.6485
R1822 B.n943 B.n942 46.6485
R1823 B.n942 B.n8 46.6485
R1824 B.n12 B.n8 46.6485
R1825 B.n935 B.n12 46.6485
R1826 B.n935 B.n934 46.6485
R1827 B.n934 B.n933 46.6485
R1828 B.n927 B.n19 46.6485
R1829 B.n927 B.n926 46.6485
R1830 B.n926 B.n925 46.6485
R1831 B.n925 B.n23 46.6485
R1832 B.n919 B.n23 46.6485
R1833 B.n919 B.n918 46.6485
R1834 B.n918 B.n917 46.6485
R1835 B.n917 B.n30 46.6485
R1836 B.n911 B.n30 46.6485
R1837 B.n910 B.n909 46.6485
R1838 B.n909 B.n37 46.6485
R1839 B.n903 B.n37 46.6485
R1840 B.n903 B.n902 46.6485
R1841 B.n902 B.n901 46.6485
R1842 B.n901 B.n44 46.6485
R1843 B.n895 B.n44 46.6485
R1844 B.n895 B.n894 46.6485
R1845 B.n894 B.n893 46.6485
R1846 B.n893 B.n51 46.6485
R1847 B.n887 B.n886 46.6485
R1848 B.n886 B.n885 46.6485
R1849 B.n885 B.n58 46.6485
R1850 B.n879 B.n58 46.6485
R1851 B.n879 B.n878 46.6485
R1852 B.n878 B.n877 46.6485
R1853 B.n877 B.n65 46.6485
R1854 B.n871 B.n65 46.6485
R1855 B.n871 B.n870 46.6485
R1856 B.n870 B.n869 46.6485
R1857 B.n869 B.n72 46.6485
R1858 B.n863 B.n72 46.6485
R1859 B.n863 B.n862 46.6485
R1860 B.n861 B.n79 46.6485
R1861 B.n855 B.n79 46.6485
R1862 B.n855 B.n854 46.6485
R1863 B.n854 B.n853 46.6485
R1864 B.n853 B.n86 46.6485
R1865 B.n847 B.n86 46.6485
R1866 B.n847 B.n846 46.6485
R1867 B.n846 B.n845 46.6485
R1868 B.n559 B.t19 43.9045
R1869 B.n911 B.t0 43.9045
R1870 B.n481 B.t6 34.3005
R1871 B.t13 B.n861 34.3005
R1872 B.n455 B.n454 33.5615
R1873 B.n459 B.n236 33.5615
R1874 B.n672 B.n671 33.5615
R1875 B.n843 B.n842 33.5615
R1876 B.n583 B.t4 28.8125
R1877 B.n19 B.t1 28.8125
R1878 B.n523 B.t2 23.3245
R1879 B.t2 B.n190 23.3245
R1880 B.t3 B.n51 23.3245
R1881 B.n887 B.t3 23.3245
R1882 B B.n947 18.0485
R1883 B.n590 B.t4 17.8365
R1884 B.n933 B.t1 17.8365
R1885 B.t6 B.n218 12.3485
R1886 B.n862 B.t13 12.3485
R1887 B.n455 B.n232 10.6151
R1888 B.n465 B.n232 10.6151
R1889 B.n466 B.n465 10.6151
R1890 B.n467 B.n466 10.6151
R1891 B.n467 B.n224 10.6151
R1892 B.n477 B.n224 10.6151
R1893 B.n478 B.n477 10.6151
R1894 B.n479 B.n478 10.6151
R1895 B.n479 B.n216 10.6151
R1896 B.n489 B.n216 10.6151
R1897 B.n490 B.n489 10.6151
R1898 B.n491 B.n490 10.6151
R1899 B.n491 B.n208 10.6151
R1900 B.n501 B.n208 10.6151
R1901 B.n502 B.n501 10.6151
R1902 B.n503 B.n502 10.6151
R1903 B.n503 B.n200 10.6151
R1904 B.n513 B.n200 10.6151
R1905 B.n514 B.n513 10.6151
R1906 B.n515 B.n514 10.6151
R1907 B.n515 B.n192 10.6151
R1908 B.n525 B.n192 10.6151
R1909 B.n526 B.n525 10.6151
R1910 B.n527 B.n526 10.6151
R1911 B.n527 B.n184 10.6151
R1912 B.n537 B.n184 10.6151
R1913 B.n538 B.n537 10.6151
R1914 B.n539 B.n538 10.6151
R1915 B.n539 B.n176 10.6151
R1916 B.n549 B.n176 10.6151
R1917 B.n550 B.n549 10.6151
R1918 B.n551 B.n550 10.6151
R1919 B.n551 B.n168 10.6151
R1920 B.n561 B.n168 10.6151
R1921 B.n562 B.n561 10.6151
R1922 B.n563 B.n562 10.6151
R1923 B.n563 B.n160 10.6151
R1924 B.n573 B.n160 10.6151
R1925 B.n574 B.n573 10.6151
R1926 B.n575 B.n574 10.6151
R1927 B.n575 B.n152 10.6151
R1928 B.n586 B.n152 10.6151
R1929 B.n587 B.n586 10.6151
R1930 B.n588 B.n587 10.6151
R1931 B.n588 B.n145 10.6151
R1932 B.n599 B.n145 10.6151
R1933 B.n600 B.n599 10.6151
R1934 B.n601 B.n600 10.6151
R1935 B.n601 B.n0 10.6151
R1936 B.n454 B.n453 10.6151
R1937 B.n453 B.n240 10.6151
R1938 B.n448 B.n240 10.6151
R1939 B.n448 B.n447 10.6151
R1940 B.n447 B.n242 10.6151
R1941 B.n442 B.n242 10.6151
R1942 B.n442 B.n441 10.6151
R1943 B.n441 B.n440 10.6151
R1944 B.n440 B.n244 10.6151
R1945 B.n434 B.n244 10.6151
R1946 B.n434 B.n433 10.6151
R1947 B.n433 B.n432 10.6151
R1948 B.n432 B.n246 10.6151
R1949 B.n426 B.n246 10.6151
R1950 B.n426 B.n425 10.6151
R1951 B.n425 B.n424 10.6151
R1952 B.n424 B.n248 10.6151
R1953 B.n418 B.n248 10.6151
R1954 B.n418 B.n417 10.6151
R1955 B.n417 B.n416 10.6151
R1956 B.n416 B.n250 10.6151
R1957 B.n410 B.n250 10.6151
R1958 B.n410 B.n409 10.6151
R1959 B.n409 B.n408 10.6151
R1960 B.n408 B.n252 10.6151
R1961 B.n402 B.n252 10.6151
R1962 B.n402 B.n401 10.6151
R1963 B.n401 B.n400 10.6151
R1964 B.n400 B.n254 10.6151
R1965 B.n394 B.n254 10.6151
R1966 B.n394 B.n393 10.6151
R1967 B.n393 B.n392 10.6151
R1968 B.n392 B.n256 10.6151
R1969 B.n386 B.n256 10.6151
R1970 B.n386 B.n385 10.6151
R1971 B.n385 B.n384 10.6151
R1972 B.n384 B.n258 10.6151
R1973 B.n378 B.n377 10.6151
R1974 B.n377 B.n376 10.6151
R1975 B.n376 B.n263 10.6151
R1976 B.n370 B.n263 10.6151
R1977 B.n370 B.n369 10.6151
R1978 B.n369 B.n368 10.6151
R1979 B.n368 B.n265 10.6151
R1980 B.n362 B.n265 10.6151
R1981 B.n360 B.n359 10.6151
R1982 B.n359 B.n269 10.6151
R1983 B.n353 B.n269 10.6151
R1984 B.n353 B.n352 10.6151
R1985 B.n352 B.n351 10.6151
R1986 B.n351 B.n271 10.6151
R1987 B.n345 B.n271 10.6151
R1988 B.n345 B.n344 10.6151
R1989 B.n344 B.n343 10.6151
R1990 B.n343 B.n273 10.6151
R1991 B.n337 B.n273 10.6151
R1992 B.n337 B.n336 10.6151
R1993 B.n336 B.n335 10.6151
R1994 B.n335 B.n275 10.6151
R1995 B.n329 B.n275 10.6151
R1996 B.n329 B.n328 10.6151
R1997 B.n328 B.n327 10.6151
R1998 B.n327 B.n277 10.6151
R1999 B.n321 B.n277 10.6151
R2000 B.n321 B.n320 10.6151
R2001 B.n320 B.n319 10.6151
R2002 B.n319 B.n279 10.6151
R2003 B.n313 B.n279 10.6151
R2004 B.n313 B.n312 10.6151
R2005 B.n312 B.n311 10.6151
R2006 B.n311 B.n281 10.6151
R2007 B.n305 B.n281 10.6151
R2008 B.n305 B.n304 10.6151
R2009 B.n304 B.n303 10.6151
R2010 B.n303 B.n283 10.6151
R2011 B.n297 B.n283 10.6151
R2012 B.n297 B.n296 10.6151
R2013 B.n296 B.n295 10.6151
R2014 B.n295 B.n285 10.6151
R2015 B.n289 B.n285 10.6151
R2016 B.n289 B.n288 10.6151
R2017 B.n288 B.n236 10.6151
R2018 B.n460 B.n459 10.6151
R2019 B.n461 B.n460 10.6151
R2020 B.n461 B.n228 10.6151
R2021 B.n471 B.n228 10.6151
R2022 B.n472 B.n471 10.6151
R2023 B.n473 B.n472 10.6151
R2024 B.n473 B.n220 10.6151
R2025 B.n483 B.n220 10.6151
R2026 B.n484 B.n483 10.6151
R2027 B.n485 B.n484 10.6151
R2028 B.n485 B.n212 10.6151
R2029 B.n495 B.n212 10.6151
R2030 B.n496 B.n495 10.6151
R2031 B.n497 B.n496 10.6151
R2032 B.n497 B.n204 10.6151
R2033 B.n507 B.n204 10.6151
R2034 B.n508 B.n507 10.6151
R2035 B.n509 B.n508 10.6151
R2036 B.n509 B.n196 10.6151
R2037 B.n519 B.n196 10.6151
R2038 B.n520 B.n519 10.6151
R2039 B.n521 B.n520 10.6151
R2040 B.n521 B.n188 10.6151
R2041 B.n531 B.n188 10.6151
R2042 B.n532 B.n531 10.6151
R2043 B.n533 B.n532 10.6151
R2044 B.n533 B.n180 10.6151
R2045 B.n543 B.n180 10.6151
R2046 B.n544 B.n543 10.6151
R2047 B.n545 B.n544 10.6151
R2048 B.n545 B.n171 10.6151
R2049 B.n555 B.n171 10.6151
R2050 B.n556 B.n555 10.6151
R2051 B.n557 B.n556 10.6151
R2052 B.n557 B.n164 10.6151
R2053 B.n567 B.n164 10.6151
R2054 B.n568 B.n567 10.6151
R2055 B.n569 B.n568 10.6151
R2056 B.n569 B.n156 10.6151
R2057 B.n579 B.n156 10.6151
R2058 B.n580 B.n579 10.6151
R2059 B.n581 B.n580 10.6151
R2060 B.n581 B.n149 10.6151
R2061 B.n592 B.n149 10.6151
R2062 B.n593 B.n592 10.6151
R2063 B.n595 B.n593 10.6151
R2064 B.n595 B.n594 10.6151
R2065 B.n594 B.n141 10.6151
R2066 B.n606 B.n141 10.6151
R2067 B.n607 B.n606 10.6151
R2068 B.n608 B.n607 10.6151
R2069 B.n609 B.n608 10.6151
R2070 B.n610 B.n609 10.6151
R2071 B.n613 B.n610 10.6151
R2072 B.n614 B.n613 10.6151
R2073 B.n615 B.n614 10.6151
R2074 B.n616 B.n615 10.6151
R2075 B.n618 B.n616 10.6151
R2076 B.n619 B.n618 10.6151
R2077 B.n620 B.n619 10.6151
R2078 B.n621 B.n620 10.6151
R2079 B.n623 B.n621 10.6151
R2080 B.n624 B.n623 10.6151
R2081 B.n625 B.n624 10.6151
R2082 B.n626 B.n625 10.6151
R2083 B.n628 B.n626 10.6151
R2084 B.n629 B.n628 10.6151
R2085 B.n630 B.n629 10.6151
R2086 B.n631 B.n630 10.6151
R2087 B.n633 B.n631 10.6151
R2088 B.n634 B.n633 10.6151
R2089 B.n635 B.n634 10.6151
R2090 B.n636 B.n635 10.6151
R2091 B.n638 B.n636 10.6151
R2092 B.n639 B.n638 10.6151
R2093 B.n640 B.n639 10.6151
R2094 B.n641 B.n640 10.6151
R2095 B.n643 B.n641 10.6151
R2096 B.n644 B.n643 10.6151
R2097 B.n645 B.n644 10.6151
R2098 B.n646 B.n645 10.6151
R2099 B.n648 B.n646 10.6151
R2100 B.n649 B.n648 10.6151
R2101 B.n650 B.n649 10.6151
R2102 B.n651 B.n650 10.6151
R2103 B.n653 B.n651 10.6151
R2104 B.n654 B.n653 10.6151
R2105 B.n655 B.n654 10.6151
R2106 B.n656 B.n655 10.6151
R2107 B.n658 B.n656 10.6151
R2108 B.n659 B.n658 10.6151
R2109 B.n660 B.n659 10.6151
R2110 B.n661 B.n660 10.6151
R2111 B.n663 B.n661 10.6151
R2112 B.n664 B.n663 10.6151
R2113 B.n665 B.n664 10.6151
R2114 B.n666 B.n665 10.6151
R2115 B.n668 B.n666 10.6151
R2116 B.n669 B.n668 10.6151
R2117 B.n670 B.n669 10.6151
R2118 B.n671 B.n670 10.6151
R2119 B.n939 B.n1 10.6151
R2120 B.n939 B.n938 10.6151
R2121 B.n938 B.n937 10.6151
R2122 B.n937 B.n10 10.6151
R2123 B.n931 B.n10 10.6151
R2124 B.n931 B.n930 10.6151
R2125 B.n930 B.n929 10.6151
R2126 B.n929 B.n17 10.6151
R2127 B.n923 B.n17 10.6151
R2128 B.n923 B.n922 10.6151
R2129 B.n922 B.n921 10.6151
R2130 B.n921 B.n25 10.6151
R2131 B.n915 B.n25 10.6151
R2132 B.n915 B.n914 10.6151
R2133 B.n914 B.n913 10.6151
R2134 B.n913 B.n32 10.6151
R2135 B.n907 B.n32 10.6151
R2136 B.n907 B.n906 10.6151
R2137 B.n906 B.n905 10.6151
R2138 B.n905 B.n39 10.6151
R2139 B.n899 B.n39 10.6151
R2140 B.n899 B.n898 10.6151
R2141 B.n898 B.n897 10.6151
R2142 B.n897 B.n46 10.6151
R2143 B.n891 B.n46 10.6151
R2144 B.n891 B.n890 10.6151
R2145 B.n890 B.n889 10.6151
R2146 B.n889 B.n53 10.6151
R2147 B.n883 B.n53 10.6151
R2148 B.n883 B.n882 10.6151
R2149 B.n882 B.n881 10.6151
R2150 B.n881 B.n60 10.6151
R2151 B.n875 B.n60 10.6151
R2152 B.n875 B.n874 10.6151
R2153 B.n874 B.n873 10.6151
R2154 B.n873 B.n67 10.6151
R2155 B.n867 B.n67 10.6151
R2156 B.n867 B.n866 10.6151
R2157 B.n866 B.n865 10.6151
R2158 B.n865 B.n74 10.6151
R2159 B.n859 B.n74 10.6151
R2160 B.n859 B.n858 10.6151
R2161 B.n858 B.n857 10.6151
R2162 B.n857 B.n81 10.6151
R2163 B.n851 B.n81 10.6151
R2164 B.n851 B.n850 10.6151
R2165 B.n850 B.n849 10.6151
R2166 B.n849 B.n88 10.6151
R2167 B.n843 B.n88 10.6151
R2168 B.n842 B.n841 10.6151
R2169 B.n841 B.n95 10.6151
R2170 B.n835 B.n95 10.6151
R2171 B.n835 B.n834 10.6151
R2172 B.n834 B.n833 10.6151
R2173 B.n833 B.n97 10.6151
R2174 B.n827 B.n97 10.6151
R2175 B.n827 B.n826 10.6151
R2176 B.n826 B.n825 10.6151
R2177 B.n825 B.n99 10.6151
R2178 B.n819 B.n99 10.6151
R2179 B.n819 B.n818 10.6151
R2180 B.n818 B.n817 10.6151
R2181 B.n817 B.n101 10.6151
R2182 B.n811 B.n101 10.6151
R2183 B.n811 B.n810 10.6151
R2184 B.n810 B.n809 10.6151
R2185 B.n809 B.n103 10.6151
R2186 B.n803 B.n103 10.6151
R2187 B.n803 B.n802 10.6151
R2188 B.n802 B.n801 10.6151
R2189 B.n801 B.n105 10.6151
R2190 B.n795 B.n105 10.6151
R2191 B.n795 B.n794 10.6151
R2192 B.n794 B.n793 10.6151
R2193 B.n793 B.n107 10.6151
R2194 B.n787 B.n107 10.6151
R2195 B.n787 B.n786 10.6151
R2196 B.n786 B.n785 10.6151
R2197 B.n785 B.n109 10.6151
R2198 B.n779 B.n109 10.6151
R2199 B.n779 B.n778 10.6151
R2200 B.n778 B.n777 10.6151
R2201 B.n777 B.n111 10.6151
R2202 B.n771 B.n111 10.6151
R2203 B.n771 B.n770 10.6151
R2204 B.n770 B.n769 10.6151
R2205 B.n765 B.n764 10.6151
R2206 B.n764 B.n117 10.6151
R2207 B.n759 B.n117 10.6151
R2208 B.n759 B.n758 10.6151
R2209 B.n758 B.n757 10.6151
R2210 B.n757 B.n119 10.6151
R2211 B.n751 B.n119 10.6151
R2212 B.n751 B.n750 10.6151
R2213 B.n748 B.n123 10.6151
R2214 B.n742 B.n123 10.6151
R2215 B.n742 B.n741 10.6151
R2216 B.n741 B.n740 10.6151
R2217 B.n740 B.n125 10.6151
R2218 B.n734 B.n125 10.6151
R2219 B.n734 B.n733 10.6151
R2220 B.n733 B.n732 10.6151
R2221 B.n732 B.n127 10.6151
R2222 B.n726 B.n127 10.6151
R2223 B.n726 B.n725 10.6151
R2224 B.n725 B.n724 10.6151
R2225 B.n724 B.n129 10.6151
R2226 B.n718 B.n129 10.6151
R2227 B.n718 B.n717 10.6151
R2228 B.n717 B.n716 10.6151
R2229 B.n716 B.n131 10.6151
R2230 B.n710 B.n131 10.6151
R2231 B.n710 B.n709 10.6151
R2232 B.n709 B.n708 10.6151
R2233 B.n708 B.n133 10.6151
R2234 B.n702 B.n133 10.6151
R2235 B.n702 B.n701 10.6151
R2236 B.n701 B.n700 10.6151
R2237 B.n700 B.n135 10.6151
R2238 B.n694 B.n135 10.6151
R2239 B.n694 B.n693 10.6151
R2240 B.n693 B.n692 10.6151
R2241 B.n692 B.n137 10.6151
R2242 B.n686 B.n137 10.6151
R2243 B.n686 B.n685 10.6151
R2244 B.n685 B.n684 10.6151
R2245 B.n684 B.n139 10.6151
R2246 B.n678 B.n139 10.6151
R2247 B.n678 B.n677 10.6151
R2248 B.n677 B.n676 10.6151
R2249 B.n676 B.n672 10.6151
R2250 B.n947 B.n0 8.11757
R2251 B.n947 B.n1 8.11757
R2252 B.n378 B.n262 6.5566
R2253 B.n362 B.n361 6.5566
R2254 B.n765 B.n115 6.5566
R2255 B.n750 B.n749 6.5566
R2256 B.n262 B.n258 4.05904
R2257 B.n361 B.n360 4.05904
R2258 B.n769 B.n115 4.05904
R2259 B.n749 B.n748 4.05904
R2260 B.n174 B.t19 2.7445
R2261 B.t0 B.n910 2.7445
R2262 VN.n34 VN.n33 161.3
R2263 VN.n32 VN.n19 161.3
R2264 VN.n31 VN.n30 161.3
R2265 VN.n29 VN.n20 161.3
R2266 VN.n28 VN.n27 161.3
R2267 VN.n26 VN.n21 161.3
R2268 VN.n25 VN.n24 161.3
R2269 VN.n16 VN.n15 161.3
R2270 VN.n14 VN.n1 161.3
R2271 VN.n13 VN.n12 161.3
R2272 VN.n11 VN.n2 161.3
R2273 VN.n10 VN.n9 161.3
R2274 VN.n8 VN.n3 161.3
R2275 VN.n7 VN.n6 161.3
R2276 VN.n23 VN.t2 112.769
R2277 VN.n5 VN.t3 112.769
R2278 VN.n4 VN.t1 79.5453
R2279 VN.n0 VN.t0 79.5453
R2280 VN.n22 VN.t4 79.5453
R2281 VN.n18 VN.t5 79.5453
R2282 VN.n17 VN.n0 73.5231
R2283 VN.n35 VN.n18 73.5231
R2284 VN.n5 VN.n4 62.2204
R2285 VN.n23 VN.n22 62.2204
R2286 VN VN.n35 50.6231
R2287 VN.n13 VN.n2 44.9365
R2288 VN.n31 VN.n20 44.9365
R2289 VN.n9 VN.n2 36.2176
R2290 VN.n27 VN.n20 36.2176
R2291 VN.n8 VN.n7 24.5923
R2292 VN.n9 VN.n8 24.5923
R2293 VN.n14 VN.n13 24.5923
R2294 VN.n15 VN.n14 24.5923
R2295 VN.n27 VN.n26 24.5923
R2296 VN.n26 VN.n25 24.5923
R2297 VN.n33 VN.n32 24.5923
R2298 VN.n32 VN.n31 24.5923
R2299 VN.n15 VN.n0 16.7229
R2300 VN.n33 VN.n18 16.7229
R2301 VN.n7 VN.n4 12.2964
R2302 VN.n25 VN.n22 12.2964
R2303 VN.n24 VN.n23 4.04954
R2304 VN.n6 VN.n5 4.04954
R2305 VN.n35 VN.n34 0.354861
R2306 VN.n17 VN.n16 0.354861
R2307 VN VN.n17 0.267071
R2308 VN.n34 VN.n19 0.189894
R2309 VN.n30 VN.n19 0.189894
R2310 VN.n30 VN.n29 0.189894
R2311 VN.n29 VN.n28 0.189894
R2312 VN.n28 VN.n21 0.189894
R2313 VN.n24 VN.n21 0.189894
R2314 VN.n6 VN.n3 0.189894
R2315 VN.n10 VN.n3 0.189894
R2316 VN.n11 VN.n10 0.189894
R2317 VN.n12 VN.n11 0.189894
R2318 VN.n12 VN.n1 0.189894
R2319 VN.n16 VN.n1 0.189894
R2320 VDD2.n111 VDD2.n59 289.615
R2321 VDD2.n52 VDD2.n0 289.615
R2322 VDD2.n112 VDD2.n111 185
R2323 VDD2.n110 VDD2.n109 185
R2324 VDD2.n63 VDD2.n62 185
R2325 VDD2.n104 VDD2.n103 185
R2326 VDD2.n102 VDD2.n101 185
R2327 VDD2.n100 VDD2.n66 185
R2328 VDD2.n70 VDD2.n67 185
R2329 VDD2.n95 VDD2.n94 185
R2330 VDD2.n93 VDD2.n92 185
R2331 VDD2.n72 VDD2.n71 185
R2332 VDD2.n87 VDD2.n86 185
R2333 VDD2.n85 VDD2.n84 185
R2334 VDD2.n76 VDD2.n75 185
R2335 VDD2.n79 VDD2.n78 185
R2336 VDD2.n19 VDD2.n18 185
R2337 VDD2.n16 VDD2.n15 185
R2338 VDD2.n25 VDD2.n24 185
R2339 VDD2.n27 VDD2.n26 185
R2340 VDD2.n12 VDD2.n11 185
R2341 VDD2.n33 VDD2.n32 185
R2342 VDD2.n36 VDD2.n35 185
R2343 VDD2.n34 VDD2.n8 185
R2344 VDD2.n41 VDD2.n7 185
R2345 VDD2.n43 VDD2.n42 185
R2346 VDD2.n45 VDD2.n44 185
R2347 VDD2.n4 VDD2.n3 185
R2348 VDD2.n51 VDD2.n50 185
R2349 VDD2.n53 VDD2.n52 185
R2350 VDD2.t0 VDD2.n77 149.524
R2351 VDD2.t2 VDD2.n17 149.524
R2352 VDD2.n111 VDD2.n110 104.615
R2353 VDD2.n110 VDD2.n62 104.615
R2354 VDD2.n103 VDD2.n62 104.615
R2355 VDD2.n103 VDD2.n102 104.615
R2356 VDD2.n102 VDD2.n66 104.615
R2357 VDD2.n70 VDD2.n66 104.615
R2358 VDD2.n94 VDD2.n70 104.615
R2359 VDD2.n94 VDD2.n93 104.615
R2360 VDD2.n93 VDD2.n71 104.615
R2361 VDD2.n86 VDD2.n71 104.615
R2362 VDD2.n86 VDD2.n85 104.615
R2363 VDD2.n85 VDD2.n75 104.615
R2364 VDD2.n78 VDD2.n75 104.615
R2365 VDD2.n18 VDD2.n15 104.615
R2366 VDD2.n25 VDD2.n15 104.615
R2367 VDD2.n26 VDD2.n25 104.615
R2368 VDD2.n26 VDD2.n11 104.615
R2369 VDD2.n33 VDD2.n11 104.615
R2370 VDD2.n35 VDD2.n33 104.615
R2371 VDD2.n35 VDD2.n34 104.615
R2372 VDD2.n34 VDD2.n7 104.615
R2373 VDD2.n43 VDD2.n7 104.615
R2374 VDD2.n44 VDD2.n43 104.615
R2375 VDD2.n44 VDD2.n3 104.615
R2376 VDD2.n51 VDD2.n3 104.615
R2377 VDD2.n52 VDD2.n51 104.615
R2378 VDD2.n58 VDD2.n57 64.61
R2379 VDD2 VDD2.n117 64.6072
R2380 VDD2.n58 VDD2.n56 52.6814
R2381 VDD2.n78 VDD2.t0 52.3082
R2382 VDD2.n18 VDD2.t2 52.3082
R2383 VDD2.n116 VDD2.n115 50.4157
R2384 VDD2.n116 VDD2.n58 43.0493
R2385 VDD2.n101 VDD2.n100 13.1884
R2386 VDD2.n42 VDD2.n41 13.1884
R2387 VDD2.n104 VDD2.n65 12.8005
R2388 VDD2.n99 VDD2.n67 12.8005
R2389 VDD2.n40 VDD2.n8 12.8005
R2390 VDD2.n45 VDD2.n6 12.8005
R2391 VDD2.n105 VDD2.n63 12.0247
R2392 VDD2.n96 VDD2.n95 12.0247
R2393 VDD2.n37 VDD2.n36 12.0247
R2394 VDD2.n46 VDD2.n4 12.0247
R2395 VDD2.n109 VDD2.n108 11.249
R2396 VDD2.n92 VDD2.n69 11.249
R2397 VDD2.n32 VDD2.n10 11.249
R2398 VDD2.n50 VDD2.n49 11.249
R2399 VDD2.n112 VDD2.n61 10.4732
R2400 VDD2.n91 VDD2.n72 10.4732
R2401 VDD2.n31 VDD2.n12 10.4732
R2402 VDD2.n53 VDD2.n2 10.4732
R2403 VDD2.n79 VDD2.n77 10.2747
R2404 VDD2.n19 VDD2.n17 10.2747
R2405 VDD2.n113 VDD2.n59 9.69747
R2406 VDD2.n88 VDD2.n87 9.69747
R2407 VDD2.n28 VDD2.n27 9.69747
R2408 VDD2.n54 VDD2.n0 9.69747
R2409 VDD2.n115 VDD2.n114 9.45567
R2410 VDD2.n56 VDD2.n55 9.45567
R2411 VDD2.n81 VDD2.n80 9.3005
R2412 VDD2.n83 VDD2.n82 9.3005
R2413 VDD2.n74 VDD2.n73 9.3005
R2414 VDD2.n89 VDD2.n88 9.3005
R2415 VDD2.n91 VDD2.n90 9.3005
R2416 VDD2.n69 VDD2.n68 9.3005
R2417 VDD2.n97 VDD2.n96 9.3005
R2418 VDD2.n99 VDD2.n98 9.3005
R2419 VDD2.n114 VDD2.n113 9.3005
R2420 VDD2.n61 VDD2.n60 9.3005
R2421 VDD2.n108 VDD2.n107 9.3005
R2422 VDD2.n106 VDD2.n105 9.3005
R2423 VDD2.n65 VDD2.n64 9.3005
R2424 VDD2.n55 VDD2.n54 9.3005
R2425 VDD2.n2 VDD2.n1 9.3005
R2426 VDD2.n49 VDD2.n48 9.3005
R2427 VDD2.n47 VDD2.n46 9.3005
R2428 VDD2.n6 VDD2.n5 9.3005
R2429 VDD2.n21 VDD2.n20 9.3005
R2430 VDD2.n23 VDD2.n22 9.3005
R2431 VDD2.n14 VDD2.n13 9.3005
R2432 VDD2.n29 VDD2.n28 9.3005
R2433 VDD2.n31 VDD2.n30 9.3005
R2434 VDD2.n10 VDD2.n9 9.3005
R2435 VDD2.n38 VDD2.n37 9.3005
R2436 VDD2.n40 VDD2.n39 9.3005
R2437 VDD2.n84 VDD2.n74 8.92171
R2438 VDD2.n24 VDD2.n14 8.92171
R2439 VDD2.n83 VDD2.n76 8.14595
R2440 VDD2.n23 VDD2.n16 8.14595
R2441 VDD2.n80 VDD2.n79 7.3702
R2442 VDD2.n20 VDD2.n19 7.3702
R2443 VDD2.n80 VDD2.n76 5.81868
R2444 VDD2.n20 VDD2.n16 5.81868
R2445 VDD2.n84 VDD2.n83 5.04292
R2446 VDD2.n24 VDD2.n23 5.04292
R2447 VDD2.n115 VDD2.n59 4.26717
R2448 VDD2.n87 VDD2.n74 4.26717
R2449 VDD2.n27 VDD2.n14 4.26717
R2450 VDD2.n56 VDD2.n0 4.26717
R2451 VDD2.n113 VDD2.n112 3.49141
R2452 VDD2.n88 VDD2.n72 3.49141
R2453 VDD2.n28 VDD2.n12 3.49141
R2454 VDD2.n54 VDD2.n53 3.49141
R2455 VDD2.n81 VDD2.n77 2.84303
R2456 VDD2.n21 VDD2.n17 2.84303
R2457 VDD2.n109 VDD2.n61 2.71565
R2458 VDD2.n92 VDD2.n91 2.71565
R2459 VDD2.n32 VDD2.n31 2.71565
R2460 VDD2.n50 VDD2.n2 2.71565
R2461 VDD2 VDD2.n116 2.37981
R2462 VDD2.n108 VDD2.n63 1.93989
R2463 VDD2.n95 VDD2.n69 1.93989
R2464 VDD2.n36 VDD2.n10 1.93989
R2465 VDD2.n49 VDD2.n4 1.93989
R2466 VDD2.n117 VDD2.t1 1.84065
R2467 VDD2.n117 VDD2.t3 1.84065
R2468 VDD2.n57 VDD2.t4 1.84065
R2469 VDD2.n57 VDD2.t5 1.84065
R2470 VDD2.n105 VDD2.n104 1.16414
R2471 VDD2.n96 VDD2.n67 1.16414
R2472 VDD2.n37 VDD2.n8 1.16414
R2473 VDD2.n46 VDD2.n45 1.16414
R2474 VDD2.n101 VDD2.n65 0.388379
R2475 VDD2.n100 VDD2.n99 0.388379
R2476 VDD2.n41 VDD2.n40 0.388379
R2477 VDD2.n42 VDD2.n6 0.388379
R2478 VDD2.n114 VDD2.n60 0.155672
R2479 VDD2.n107 VDD2.n60 0.155672
R2480 VDD2.n107 VDD2.n106 0.155672
R2481 VDD2.n106 VDD2.n64 0.155672
R2482 VDD2.n98 VDD2.n64 0.155672
R2483 VDD2.n98 VDD2.n97 0.155672
R2484 VDD2.n97 VDD2.n68 0.155672
R2485 VDD2.n90 VDD2.n68 0.155672
R2486 VDD2.n90 VDD2.n89 0.155672
R2487 VDD2.n89 VDD2.n73 0.155672
R2488 VDD2.n82 VDD2.n73 0.155672
R2489 VDD2.n82 VDD2.n81 0.155672
R2490 VDD2.n22 VDD2.n21 0.155672
R2491 VDD2.n22 VDD2.n13 0.155672
R2492 VDD2.n29 VDD2.n13 0.155672
R2493 VDD2.n30 VDD2.n29 0.155672
R2494 VDD2.n30 VDD2.n9 0.155672
R2495 VDD2.n38 VDD2.n9 0.155672
R2496 VDD2.n39 VDD2.n38 0.155672
R2497 VDD2.n39 VDD2.n5 0.155672
R2498 VDD2.n47 VDD2.n5 0.155672
R2499 VDD2.n48 VDD2.n47 0.155672
R2500 VDD2.n48 VDD2.n1 0.155672
R2501 VDD2.n55 VDD2.n1 0.155672
C0 VP VDD1 6.67154f
C1 VTAIL VDD1 7.50666f
C2 VN VDD1 0.151845f
C3 VP VTAIL 6.70185f
C4 VP VN 7.3331f
C5 VN VTAIL 6.68762f
C6 VDD2 VDD1 1.66339f
C7 VDD2 VP 0.514404f
C8 VDD2 VTAIL 7.56275f
C9 VDD2 VN 6.31188f
C10 VDD2 B 6.266902f
C11 VDD1 B 6.428549f
C12 VTAIL B 7.737289f
C13 VN B 14.727191f
C14 VP B 13.430496f
C15 VDD2.n0 B 0.030174f
C16 VDD2.n1 B 0.021467f
C17 VDD2.n2 B 0.011535f
C18 VDD2.n3 B 0.027266f
C19 VDD2.n4 B 0.012214f
C20 VDD2.n5 B 0.021467f
C21 VDD2.n6 B 0.011535f
C22 VDD2.n7 B 0.027266f
C23 VDD2.n8 B 0.012214f
C24 VDD2.n9 B 0.021467f
C25 VDD2.n10 B 0.011535f
C26 VDD2.n11 B 0.027266f
C27 VDD2.n12 B 0.012214f
C28 VDD2.n13 B 0.021467f
C29 VDD2.n14 B 0.011535f
C30 VDD2.n15 B 0.027266f
C31 VDD2.n16 B 0.012214f
C32 VDD2.n17 B 0.144557f
C33 VDD2.t2 B 0.045907f
C34 VDD2.n18 B 0.020449f
C35 VDD2.n19 B 0.019275f
C36 VDD2.n20 B 0.011535f
C37 VDD2.n21 B 0.964576f
C38 VDD2.n22 B 0.021467f
C39 VDD2.n23 B 0.011535f
C40 VDD2.n24 B 0.012214f
C41 VDD2.n25 B 0.027266f
C42 VDD2.n26 B 0.027266f
C43 VDD2.n27 B 0.012214f
C44 VDD2.n28 B 0.011535f
C45 VDD2.n29 B 0.021467f
C46 VDD2.n30 B 0.021467f
C47 VDD2.n31 B 0.011535f
C48 VDD2.n32 B 0.012214f
C49 VDD2.n33 B 0.027266f
C50 VDD2.n34 B 0.027266f
C51 VDD2.n35 B 0.027266f
C52 VDD2.n36 B 0.012214f
C53 VDD2.n37 B 0.011535f
C54 VDD2.n38 B 0.021467f
C55 VDD2.n39 B 0.021467f
C56 VDD2.n40 B 0.011535f
C57 VDD2.n41 B 0.011875f
C58 VDD2.n42 B 0.011875f
C59 VDD2.n43 B 0.027266f
C60 VDD2.n44 B 0.027266f
C61 VDD2.n45 B 0.012214f
C62 VDD2.n46 B 0.011535f
C63 VDD2.n47 B 0.021467f
C64 VDD2.n48 B 0.021467f
C65 VDD2.n49 B 0.011535f
C66 VDD2.n50 B 0.012214f
C67 VDD2.n51 B 0.027266f
C68 VDD2.n52 B 0.059026f
C69 VDD2.n53 B 0.012214f
C70 VDD2.n54 B 0.011535f
C71 VDD2.n55 B 0.051966f
C72 VDD2.n56 B 0.056488f
C73 VDD2.t4 B 0.182532f
C74 VDD2.t5 B 0.182532f
C75 VDD2.n57 B 1.62144f
C76 VDD2.n58 B 2.47824f
C77 VDD2.n59 B 0.030174f
C78 VDD2.n60 B 0.021467f
C79 VDD2.n61 B 0.011535f
C80 VDD2.n62 B 0.027266f
C81 VDD2.n63 B 0.012214f
C82 VDD2.n64 B 0.021467f
C83 VDD2.n65 B 0.011535f
C84 VDD2.n66 B 0.027266f
C85 VDD2.n67 B 0.012214f
C86 VDD2.n68 B 0.021467f
C87 VDD2.n69 B 0.011535f
C88 VDD2.n70 B 0.027266f
C89 VDD2.n71 B 0.027266f
C90 VDD2.n72 B 0.012214f
C91 VDD2.n73 B 0.021467f
C92 VDD2.n74 B 0.011535f
C93 VDD2.n75 B 0.027266f
C94 VDD2.n76 B 0.012214f
C95 VDD2.n77 B 0.144557f
C96 VDD2.t0 B 0.045907f
C97 VDD2.n78 B 0.020449f
C98 VDD2.n79 B 0.019275f
C99 VDD2.n80 B 0.011535f
C100 VDD2.n81 B 0.964576f
C101 VDD2.n82 B 0.021467f
C102 VDD2.n83 B 0.011535f
C103 VDD2.n84 B 0.012214f
C104 VDD2.n85 B 0.027266f
C105 VDD2.n86 B 0.027266f
C106 VDD2.n87 B 0.012214f
C107 VDD2.n88 B 0.011535f
C108 VDD2.n89 B 0.021467f
C109 VDD2.n90 B 0.021467f
C110 VDD2.n91 B 0.011535f
C111 VDD2.n92 B 0.012214f
C112 VDD2.n93 B 0.027266f
C113 VDD2.n94 B 0.027266f
C114 VDD2.n95 B 0.012214f
C115 VDD2.n96 B 0.011535f
C116 VDD2.n97 B 0.021467f
C117 VDD2.n98 B 0.021467f
C118 VDD2.n99 B 0.011535f
C119 VDD2.n100 B 0.011875f
C120 VDD2.n101 B 0.011875f
C121 VDD2.n102 B 0.027266f
C122 VDD2.n103 B 0.027266f
C123 VDD2.n104 B 0.012214f
C124 VDD2.n105 B 0.011535f
C125 VDD2.n106 B 0.021467f
C126 VDD2.n107 B 0.021467f
C127 VDD2.n108 B 0.011535f
C128 VDD2.n109 B 0.012214f
C129 VDD2.n110 B 0.027266f
C130 VDD2.n111 B 0.059026f
C131 VDD2.n112 B 0.012214f
C132 VDD2.n113 B 0.011535f
C133 VDD2.n114 B 0.051966f
C134 VDD2.n115 B 0.047902f
C135 VDD2.n116 B 2.27344f
C136 VDD2.t1 B 0.182532f
C137 VDD2.t3 B 0.182532f
C138 VDD2.n117 B 1.62141f
C139 VN.t0 B 1.94966f
C140 VN.n0 B 0.771121f
C141 VN.n1 B 0.020467f
C142 VN.n2 B 0.017065f
C143 VN.n3 B 0.020467f
C144 VN.t1 B 1.94966f
C145 VN.n4 B 0.756858f
C146 VN.t3 B 2.1958f
C147 VN.n5 B 0.71937f
C148 VN.n6 B 0.238639f
C149 VN.n7 B 0.028586f
C150 VN.n8 B 0.037954f
C151 VN.n9 B 0.041082f
C152 VN.n10 B 0.020467f
C153 VN.n11 B 0.020467f
C154 VN.n12 B 0.020467f
C155 VN.n13 B 0.039311f
C156 VN.n14 B 0.037954f
C157 VN.n15 B 0.031958f
C158 VN.n16 B 0.033028f
C159 VN.n17 B 0.047489f
C160 VN.t5 B 1.94966f
C161 VN.n18 B 0.771121f
C162 VN.n19 B 0.020467f
C163 VN.n20 B 0.017065f
C164 VN.n21 B 0.020467f
C165 VN.t4 B 1.94966f
C166 VN.n22 B 0.756858f
C167 VN.t2 B 2.1958f
C168 VN.n23 B 0.71937f
C169 VN.n24 B 0.238639f
C170 VN.n25 B 0.028586f
C171 VN.n26 B 0.037954f
C172 VN.n27 B 0.041082f
C173 VN.n28 B 0.020467f
C174 VN.n29 B 0.020467f
C175 VN.n30 B 0.020467f
C176 VN.n31 B 0.039311f
C177 VN.n32 B 0.037954f
C178 VN.n33 B 0.031958f
C179 VN.n34 B 0.033028f
C180 VN.n35 B 1.18627f
C181 VTAIL.t1 B 0.209446f
C182 VTAIL.t0 B 0.209446f
C183 VTAIL.n0 B 1.78552f
C184 VTAIL.n1 B 0.462721f
C185 VTAIL.n2 B 0.034623f
C186 VTAIL.n3 B 0.024632f
C187 VTAIL.n4 B 0.013236f
C188 VTAIL.n5 B 0.031286f
C189 VTAIL.n6 B 0.014015f
C190 VTAIL.n7 B 0.024632f
C191 VTAIL.n8 B 0.013236f
C192 VTAIL.n9 B 0.031286f
C193 VTAIL.n10 B 0.014015f
C194 VTAIL.n11 B 0.024632f
C195 VTAIL.n12 B 0.013236f
C196 VTAIL.n13 B 0.031286f
C197 VTAIL.n14 B 0.014015f
C198 VTAIL.n15 B 0.024632f
C199 VTAIL.n16 B 0.013236f
C200 VTAIL.n17 B 0.031286f
C201 VTAIL.n18 B 0.014015f
C202 VTAIL.n19 B 0.165871f
C203 VTAIL.t8 B 0.052676f
C204 VTAIL.n20 B 0.023464f
C205 VTAIL.n21 B 0.022117f
C206 VTAIL.n22 B 0.013236f
C207 VTAIL.n23 B 1.1068f
C208 VTAIL.n24 B 0.024632f
C209 VTAIL.n25 B 0.013236f
C210 VTAIL.n26 B 0.014015f
C211 VTAIL.n27 B 0.031286f
C212 VTAIL.n28 B 0.031286f
C213 VTAIL.n29 B 0.014015f
C214 VTAIL.n30 B 0.013236f
C215 VTAIL.n31 B 0.024632f
C216 VTAIL.n32 B 0.024632f
C217 VTAIL.n33 B 0.013236f
C218 VTAIL.n34 B 0.014015f
C219 VTAIL.n35 B 0.031286f
C220 VTAIL.n36 B 0.031286f
C221 VTAIL.n37 B 0.031286f
C222 VTAIL.n38 B 0.014015f
C223 VTAIL.n39 B 0.013236f
C224 VTAIL.n40 B 0.024632f
C225 VTAIL.n41 B 0.024632f
C226 VTAIL.n42 B 0.013236f
C227 VTAIL.n43 B 0.013626f
C228 VTAIL.n44 B 0.013626f
C229 VTAIL.n45 B 0.031286f
C230 VTAIL.n46 B 0.031286f
C231 VTAIL.n47 B 0.014015f
C232 VTAIL.n48 B 0.013236f
C233 VTAIL.n49 B 0.024632f
C234 VTAIL.n50 B 0.024632f
C235 VTAIL.n51 B 0.013236f
C236 VTAIL.n52 B 0.014015f
C237 VTAIL.n53 B 0.031286f
C238 VTAIL.n54 B 0.067729f
C239 VTAIL.n55 B 0.014015f
C240 VTAIL.n56 B 0.013236f
C241 VTAIL.n57 B 0.059628f
C242 VTAIL.n58 B 0.037978f
C243 VTAIL.n59 B 0.428308f
C244 VTAIL.t7 B 0.209446f
C245 VTAIL.t9 B 0.209446f
C246 VTAIL.n60 B 1.78552f
C247 VTAIL.n61 B 2.04433f
C248 VTAIL.t2 B 0.209446f
C249 VTAIL.t11 B 0.209446f
C250 VTAIL.n62 B 1.78553f
C251 VTAIL.n63 B 2.04432f
C252 VTAIL.n64 B 0.034623f
C253 VTAIL.n65 B 0.024632f
C254 VTAIL.n66 B 0.013236f
C255 VTAIL.n67 B 0.031286f
C256 VTAIL.n68 B 0.014015f
C257 VTAIL.n69 B 0.024632f
C258 VTAIL.n70 B 0.013236f
C259 VTAIL.n71 B 0.031286f
C260 VTAIL.n72 B 0.014015f
C261 VTAIL.n73 B 0.024632f
C262 VTAIL.n74 B 0.013236f
C263 VTAIL.n75 B 0.031286f
C264 VTAIL.n76 B 0.031286f
C265 VTAIL.n77 B 0.014015f
C266 VTAIL.n78 B 0.024632f
C267 VTAIL.n79 B 0.013236f
C268 VTAIL.n80 B 0.031286f
C269 VTAIL.n81 B 0.014015f
C270 VTAIL.n82 B 0.165872f
C271 VTAIL.t4 B 0.052676f
C272 VTAIL.n83 B 0.023464f
C273 VTAIL.n84 B 0.022117f
C274 VTAIL.n85 B 0.013236f
C275 VTAIL.n86 B 1.1068f
C276 VTAIL.n87 B 0.024632f
C277 VTAIL.n88 B 0.013236f
C278 VTAIL.n89 B 0.014015f
C279 VTAIL.n90 B 0.031286f
C280 VTAIL.n91 B 0.031286f
C281 VTAIL.n92 B 0.014015f
C282 VTAIL.n93 B 0.013236f
C283 VTAIL.n94 B 0.024632f
C284 VTAIL.n95 B 0.024632f
C285 VTAIL.n96 B 0.013236f
C286 VTAIL.n97 B 0.014015f
C287 VTAIL.n98 B 0.031286f
C288 VTAIL.n99 B 0.031286f
C289 VTAIL.n100 B 0.014015f
C290 VTAIL.n101 B 0.013236f
C291 VTAIL.n102 B 0.024632f
C292 VTAIL.n103 B 0.024632f
C293 VTAIL.n104 B 0.013236f
C294 VTAIL.n105 B 0.013626f
C295 VTAIL.n106 B 0.013626f
C296 VTAIL.n107 B 0.031286f
C297 VTAIL.n108 B 0.031286f
C298 VTAIL.n109 B 0.014015f
C299 VTAIL.n110 B 0.013236f
C300 VTAIL.n111 B 0.024632f
C301 VTAIL.n112 B 0.024632f
C302 VTAIL.n113 B 0.013236f
C303 VTAIL.n114 B 0.014015f
C304 VTAIL.n115 B 0.031286f
C305 VTAIL.n116 B 0.067729f
C306 VTAIL.n117 B 0.014015f
C307 VTAIL.n118 B 0.013236f
C308 VTAIL.n119 B 0.059628f
C309 VTAIL.n120 B 0.037978f
C310 VTAIL.n121 B 0.428308f
C311 VTAIL.t6 B 0.209446f
C312 VTAIL.t10 B 0.209446f
C313 VTAIL.n122 B 1.78553f
C314 VTAIL.n123 B 0.642321f
C315 VTAIL.n124 B 0.034623f
C316 VTAIL.n125 B 0.024632f
C317 VTAIL.n126 B 0.013236f
C318 VTAIL.n127 B 0.031286f
C319 VTAIL.n128 B 0.014015f
C320 VTAIL.n129 B 0.024632f
C321 VTAIL.n130 B 0.013236f
C322 VTAIL.n131 B 0.031286f
C323 VTAIL.n132 B 0.014015f
C324 VTAIL.n133 B 0.024632f
C325 VTAIL.n134 B 0.013236f
C326 VTAIL.n135 B 0.031286f
C327 VTAIL.n136 B 0.031286f
C328 VTAIL.n137 B 0.014015f
C329 VTAIL.n138 B 0.024632f
C330 VTAIL.n139 B 0.013236f
C331 VTAIL.n140 B 0.031286f
C332 VTAIL.n141 B 0.014015f
C333 VTAIL.n142 B 0.165872f
C334 VTAIL.t5 B 0.052676f
C335 VTAIL.n143 B 0.023464f
C336 VTAIL.n144 B 0.022117f
C337 VTAIL.n145 B 0.013236f
C338 VTAIL.n146 B 1.1068f
C339 VTAIL.n147 B 0.024632f
C340 VTAIL.n148 B 0.013236f
C341 VTAIL.n149 B 0.014015f
C342 VTAIL.n150 B 0.031286f
C343 VTAIL.n151 B 0.031286f
C344 VTAIL.n152 B 0.014015f
C345 VTAIL.n153 B 0.013236f
C346 VTAIL.n154 B 0.024632f
C347 VTAIL.n155 B 0.024632f
C348 VTAIL.n156 B 0.013236f
C349 VTAIL.n157 B 0.014015f
C350 VTAIL.n158 B 0.031286f
C351 VTAIL.n159 B 0.031286f
C352 VTAIL.n160 B 0.014015f
C353 VTAIL.n161 B 0.013236f
C354 VTAIL.n162 B 0.024632f
C355 VTAIL.n163 B 0.024632f
C356 VTAIL.n164 B 0.013236f
C357 VTAIL.n165 B 0.013626f
C358 VTAIL.n166 B 0.013626f
C359 VTAIL.n167 B 0.031286f
C360 VTAIL.n168 B 0.031286f
C361 VTAIL.n169 B 0.014015f
C362 VTAIL.n170 B 0.013236f
C363 VTAIL.n171 B 0.024632f
C364 VTAIL.n172 B 0.024632f
C365 VTAIL.n173 B 0.013236f
C366 VTAIL.n174 B 0.014015f
C367 VTAIL.n175 B 0.031286f
C368 VTAIL.n176 B 0.067729f
C369 VTAIL.n177 B 0.014015f
C370 VTAIL.n178 B 0.013236f
C371 VTAIL.n179 B 0.059628f
C372 VTAIL.n180 B 0.037978f
C373 VTAIL.n181 B 1.58467f
C374 VTAIL.n182 B 0.034623f
C375 VTAIL.n183 B 0.024632f
C376 VTAIL.n184 B 0.013236f
C377 VTAIL.n185 B 0.031286f
C378 VTAIL.n186 B 0.014015f
C379 VTAIL.n187 B 0.024632f
C380 VTAIL.n188 B 0.013236f
C381 VTAIL.n189 B 0.031286f
C382 VTAIL.n190 B 0.014015f
C383 VTAIL.n191 B 0.024632f
C384 VTAIL.n192 B 0.013236f
C385 VTAIL.n193 B 0.031286f
C386 VTAIL.n194 B 0.014015f
C387 VTAIL.n195 B 0.024632f
C388 VTAIL.n196 B 0.013236f
C389 VTAIL.n197 B 0.031286f
C390 VTAIL.n198 B 0.014015f
C391 VTAIL.n199 B 0.165871f
C392 VTAIL.t3 B 0.052676f
C393 VTAIL.n200 B 0.023464f
C394 VTAIL.n201 B 0.022117f
C395 VTAIL.n202 B 0.013236f
C396 VTAIL.n203 B 1.1068f
C397 VTAIL.n204 B 0.024632f
C398 VTAIL.n205 B 0.013236f
C399 VTAIL.n206 B 0.014015f
C400 VTAIL.n207 B 0.031286f
C401 VTAIL.n208 B 0.031286f
C402 VTAIL.n209 B 0.014015f
C403 VTAIL.n210 B 0.013236f
C404 VTAIL.n211 B 0.024632f
C405 VTAIL.n212 B 0.024632f
C406 VTAIL.n213 B 0.013236f
C407 VTAIL.n214 B 0.014015f
C408 VTAIL.n215 B 0.031286f
C409 VTAIL.n216 B 0.031286f
C410 VTAIL.n217 B 0.031286f
C411 VTAIL.n218 B 0.014015f
C412 VTAIL.n219 B 0.013236f
C413 VTAIL.n220 B 0.024632f
C414 VTAIL.n221 B 0.024632f
C415 VTAIL.n222 B 0.013236f
C416 VTAIL.n223 B 0.013626f
C417 VTAIL.n224 B 0.013626f
C418 VTAIL.n225 B 0.031286f
C419 VTAIL.n226 B 0.031286f
C420 VTAIL.n227 B 0.014015f
C421 VTAIL.n228 B 0.013236f
C422 VTAIL.n229 B 0.024632f
C423 VTAIL.n230 B 0.024632f
C424 VTAIL.n231 B 0.013236f
C425 VTAIL.n232 B 0.014015f
C426 VTAIL.n233 B 0.031286f
C427 VTAIL.n234 B 0.067729f
C428 VTAIL.n235 B 0.014015f
C429 VTAIL.n236 B 0.013236f
C430 VTAIL.n237 B 0.059628f
C431 VTAIL.n238 B 0.037978f
C432 VTAIL.n239 B 1.51864f
C433 VDD1.n0 B 0.03065f
C434 VDD1.n1 B 0.021806f
C435 VDD1.n2 B 0.011718f
C436 VDD1.n3 B 0.027696f
C437 VDD1.n4 B 0.012407f
C438 VDD1.n5 B 0.021806f
C439 VDD1.n6 B 0.011718f
C440 VDD1.n7 B 0.027696f
C441 VDD1.n8 B 0.012407f
C442 VDD1.n9 B 0.021806f
C443 VDD1.n10 B 0.011718f
C444 VDD1.n11 B 0.027696f
C445 VDD1.n12 B 0.027696f
C446 VDD1.n13 B 0.012407f
C447 VDD1.n14 B 0.021806f
C448 VDD1.n15 B 0.011718f
C449 VDD1.n16 B 0.027696f
C450 VDD1.n17 B 0.012407f
C451 VDD1.n18 B 0.146839f
C452 VDD1.t2 B 0.046632f
C453 VDD1.n19 B 0.020772f
C454 VDD1.n20 B 0.019579f
C455 VDD1.n21 B 0.011718f
C456 VDD1.n22 B 0.979805f
C457 VDD1.n23 B 0.021806f
C458 VDD1.n24 B 0.011718f
C459 VDD1.n25 B 0.012407f
C460 VDD1.n26 B 0.027696f
C461 VDD1.n27 B 0.027696f
C462 VDD1.n28 B 0.012407f
C463 VDD1.n29 B 0.011718f
C464 VDD1.n30 B 0.021806f
C465 VDD1.n31 B 0.021806f
C466 VDD1.n32 B 0.011718f
C467 VDD1.n33 B 0.012407f
C468 VDD1.n34 B 0.027696f
C469 VDD1.n35 B 0.027696f
C470 VDD1.n36 B 0.012407f
C471 VDD1.n37 B 0.011718f
C472 VDD1.n38 B 0.021806f
C473 VDD1.n39 B 0.021806f
C474 VDD1.n40 B 0.011718f
C475 VDD1.n41 B 0.012062f
C476 VDD1.n42 B 0.012062f
C477 VDD1.n43 B 0.027696f
C478 VDD1.n44 B 0.027696f
C479 VDD1.n45 B 0.012407f
C480 VDD1.n46 B 0.011718f
C481 VDD1.n47 B 0.021806f
C482 VDD1.n48 B 0.021806f
C483 VDD1.n49 B 0.011718f
C484 VDD1.n50 B 0.012407f
C485 VDD1.n51 B 0.027696f
C486 VDD1.n52 B 0.059957f
C487 VDD1.n53 B 0.012407f
C488 VDD1.n54 B 0.011718f
C489 VDD1.n55 B 0.052787f
C490 VDD1.n56 B 0.058147f
C491 VDD1.n57 B 0.03065f
C492 VDD1.n58 B 0.021806f
C493 VDD1.n59 B 0.011718f
C494 VDD1.n60 B 0.027696f
C495 VDD1.n61 B 0.012407f
C496 VDD1.n62 B 0.021806f
C497 VDD1.n63 B 0.011718f
C498 VDD1.n64 B 0.027696f
C499 VDD1.n65 B 0.012407f
C500 VDD1.n66 B 0.021806f
C501 VDD1.n67 B 0.011718f
C502 VDD1.n68 B 0.027696f
C503 VDD1.n69 B 0.012407f
C504 VDD1.n70 B 0.021806f
C505 VDD1.n71 B 0.011718f
C506 VDD1.n72 B 0.027696f
C507 VDD1.n73 B 0.012407f
C508 VDD1.n74 B 0.146839f
C509 VDD1.t0 B 0.046632f
C510 VDD1.n75 B 0.020772f
C511 VDD1.n76 B 0.019579f
C512 VDD1.n77 B 0.011718f
C513 VDD1.n78 B 0.979805f
C514 VDD1.n79 B 0.021806f
C515 VDD1.n80 B 0.011718f
C516 VDD1.n81 B 0.012407f
C517 VDD1.n82 B 0.027696f
C518 VDD1.n83 B 0.027696f
C519 VDD1.n84 B 0.012407f
C520 VDD1.n85 B 0.011718f
C521 VDD1.n86 B 0.021806f
C522 VDD1.n87 B 0.021806f
C523 VDD1.n88 B 0.011718f
C524 VDD1.n89 B 0.012407f
C525 VDD1.n90 B 0.027696f
C526 VDD1.n91 B 0.027696f
C527 VDD1.n92 B 0.027696f
C528 VDD1.n93 B 0.012407f
C529 VDD1.n94 B 0.011718f
C530 VDD1.n95 B 0.021806f
C531 VDD1.n96 B 0.021806f
C532 VDD1.n97 B 0.011718f
C533 VDD1.n98 B 0.012062f
C534 VDD1.n99 B 0.012062f
C535 VDD1.n100 B 0.027696f
C536 VDD1.n101 B 0.027696f
C537 VDD1.n102 B 0.012407f
C538 VDD1.n103 B 0.011718f
C539 VDD1.n104 B 0.021806f
C540 VDD1.n105 B 0.021806f
C541 VDD1.n106 B 0.011718f
C542 VDD1.n107 B 0.012407f
C543 VDD1.n108 B 0.027696f
C544 VDD1.n109 B 0.059957f
C545 VDD1.n110 B 0.012407f
C546 VDD1.n111 B 0.011718f
C547 VDD1.n112 B 0.052787f
C548 VDD1.n113 B 0.05738f
C549 VDD1.t4 B 0.185414f
C550 VDD1.t3 B 0.185414f
C551 VDD1.n114 B 1.64704f
C552 VDD1.n115 B 2.63987f
C553 VDD1.t1 B 0.185414f
C554 VDD1.t5 B 0.185414f
C555 VDD1.n116 B 1.64198f
C556 VDD1.n117 B 2.5111f
C557 VP.t2 B 1.9909f
C558 VP.n0 B 0.787431f
C559 VP.n1 B 0.0209f
C560 VP.n2 B 0.017426f
C561 VP.n3 B 0.0209f
C562 VP.t1 B 1.9909f
C563 VP.n4 B 0.703981f
C564 VP.n5 B 0.0209f
C565 VP.n6 B 0.017426f
C566 VP.n7 B 0.0209f
C567 VP.t3 B 1.9909f
C568 VP.n8 B 0.787431f
C569 VP.t5 B 1.9909f
C570 VP.n9 B 0.787431f
C571 VP.n10 B 0.0209f
C572 VP.n11 B 0.017426f
C573 VP.n12 B 0.0209f
C574 VP.t0 B 1.9909f
C575 VP.n13 B 0.772866f
C576 VP.t4 B 2.24224f
C577 VP.n14 B 0.734587f
C578 VP.n15 B 0.243687f
C579 VP.n16 B 0.02919f
C580 VP.n17 B 0.038757f
C581 VP.n18 B 0.041951f
C582 VP.n19 B 0.0209f
C583 VP.n20 B 0.0209f
C584 VP.n21 B 0.0209f
C585 VP.n22 B 0.040143f
C586 VP.n23 B 0.038757f
C587 VP.n24 B 0.032634f
C588 VP.n25 B 0.033727f
C589 VP.n26 B 1.20285f
C590 VP.n27 B 1.21778f
C591 VP.n28 B 0.033727f
C592 VP.n29 B 0.032634f
C593 VP.n30 B 0.038757f
C594 VP.n31 B 0.040143f
C595 VP.n32 B 0.0209f
C596 VP.n33 B 0.0209f
C597 VP.n34 B 0.0209f
C598 VP.n35 B 0.041951f
C599 VP.n36 B 0.038757f
C600 VP.n37 B 0.02919f
C601 VP.n38 B 0.0209f
C602 VP.n39 B 0.0209f
C603 VP.n40 B 0.02919f
C604 VP.n41 B 0.038757f
C605 VP.n42 B 0.041951f
C606 VP.n43 B 0.0209f
C607 VP.n44 B 0.0209f
C608 VP.n45 B 0.0209f
C609 VP.n46 B 0.040143f
C610 VP.n47 B 0.038757f
C611 VP.n48 B 0.032634f
C612 VP.n49 B 0.033727f
C613 VP.n50 B 0.048493f
.ends

