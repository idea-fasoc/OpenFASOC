* NGSPICE file created from diff_pair_sample_1114.ext - technology: sky130A

.subckt diff_pair_sample_1114 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0.11715 ps=1.04 w=0.71 l=1.74
X1 VDD1.t1 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.11715 pd=1.04 as=0.2769 ps=2.2 w=0.71 l=1.74
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0 ps=0 w=0.71 l=1.74
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0 ps=0 w=0.71 l=1.74
X4 VTAIL.t2 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0.11715 ps=1.04 w=0.71 l=1.74
X5 VDD1.t2 VP.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.11715 pd=1.04 as=0.2769 ps=2.2 w=0.71 l=1.74
X6 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.11715 pd=1.04 as=0.2769 ps=2.2 w=0.71 l=1.74
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0 ps=0 w=0.71 l=1.74
X8 VTAIL.t4 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0.11715 ps=1.04 w=0.71 l=1.74
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0 ps=0 w=0.71 l=1.74
X10 VTAIL.t3 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2769 pd=2.2 as=0.11715 ps=1.04 w=0.71 l=1.74
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.11715 pd=1.04 as=0.2769 ps=2.2 w=0.71 l=1.74
R0 VP.n5 VP.n4 184.054
R1 VP.n14 VP.n13 184.054
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t0 45.4791
R8 VP.n3 VP.t2 45.054
R9 VP.n4 VP.n3 44.4511
R10 VP.n7 VP.n1 40.4934
R11 VP.n11 VP.n1 40.4934
R12 VP.n7 VP.n6 24.4675
R13 VP.n12 VP.n11 24.4675
R14 VP.n5 VP.t3 9.83441
R15 VP.n13 VP.t1 9.83441
R16 VP.n6 VP.n5 1.71319
R17 VP.n13 VP.n12 1.71319
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VDD1 VDD1.n1 266.202
R26 VDD1 VDD1.n0 236.055
R27 VDD1.n0 VDD1.t3 27.8878
R28 VDD1.n0 VDD1.t2 27.8878
R29 VDD1.n1 VDD1.t0 27.8878
R30 VDD1.n1 VDD1.t1 27.8878
R31 VTAIL.n7 VTAIL.t0 247.207
R32 VTAIL.n0 VTAIL.t2 247.207
R33 VTAIL.n1 VTAIL.t6 247.207
R34 VTAIL.n2 VTAIL.t4 247.207
R35 VTAIL.n6 VTAIL.t5 247.207
R36 VTAIL.n5 VTAIL.t7 247.207
R37 VTAIL.n4 VTAIL.t1 247.207
R38 VTAIL.n3 VTAIL.t3 247.207
R39 VTAIL.n7 VTAIL.n6 14.7634
R40 VTAIL.n3 VTAIL.n2 14.7634
R41 VTAIL.n4 VTAIL.n3 1.78498
R42 VTAIL.n6 VTAIL.n5 1.78498
R43 VTAIL.n2 VTAIL.n1 1.78498
R44 VTAIL VTAIL.n0 0.950931
R45 VTAIL VTAIL.n7 0.834552
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 B.n304 B.n303 585
R49 B.n306 B.n69 585
R50 B.n309 B.n308 585
R51 B.n310 B.n68 585
R52 B.n312 B.n311 585
R53 B.n314 B.n67 585
R54 B.n316 B.n315 585
R55 B.n318 B.n317 585
R56 B.n321 B.n320 585
R57 B.n322 B.n62 585
R58 B.n324 B.n323 585
R59 B.n326 B.n61 585
R60 B.n329 B.n328 585
R61 B.n330 B.n60 585
R62 B.n332 B.n331 585
R63 B.n334 B.n59 585
R64 B.n337 B.n336 585
R65 B.n338 B.n56 585
R66 B.n341 B.n340 585
R67 B.n343 B.n55 585
R68 B.n346 B.n345 585
R69 B.n347 B.n54 585
R70 B.n349 B.n348 585
R71 B.n351 B.n53 585
R72 B.n354 B.n353 585
R73 B.n355 B.n52 585
R74 B.n302 B.n50 585
R75 B.n358 B.n50 585
R76 B.n301 B.n49 585
R77 B.n359 B.n49 585
R78 B.n300 B.n48 585
R79 B.n360 B.n48 585
R80 B.n299 B.n298 585
R81 B.n298 B.n44 585
R82 B.n297 B.n43 585
R83 B.n366 B.n43 585
R84 B.n296 B.n42 585
R85 B.n367 B.n42 585
R86 B.n295 B.n41 585
R87 B.n368 B.n41 585
R88 B.n294 B.n293 585
R89 B.n293 B.n37 585
R90 B.n292 B.n36 585
R91 B.n374 B.n36 585
R92 B.n291 B.n35 585
R93 B.n375 B.n35 585
R94 B.n290 B.n34 585
R95 B.n376 B.n34 585
R96 B.n289 B.n288 585
R97 B.n288 B.n30 585
R98 B.n287 B.n29 585
R99 B.n382 B.n29 585
R100 B.n286 B.n28 585
R101 B.n383 B.n28 585
R102 B.n285 B.n27 585
R103 B.n384 B.n27 585
R104 B.n284 B.n283 585
R105 B.n283 B.n26 585
R106 B.n282 B.n22 585
R107 B.n390 B.n22 585
R108 B.n281 B.n21 585
R109 B.n391 B.n21 585
R110 B.n280 B.n20 585
R111 B.n392 B.n20 585
R112 B.n279 B.n278 585
R113 B.n278 B.n16 585
R114 B.n277 B.n15 585
R115 B.n398 B.n15 585
R116 B.n276 B.n14 585
R117 B.n399 B.n14 585
R118 B.n275 B.n13 585
R119 B.n400 B.n13 585
R120 B.n274 B.n273 585
R121 B.n273 B.n12 585
R122 B.n272 B.n271 585
R123 B.n272 B.n8 585
R124 B.n270 B.n7 585
R125 B.n407 B.n7 585
R126 B.n269 B.n6 585
R127 B.n408 B.n6 585
R128 B.n268 B.n5 585
R129 B.n409 B.n5 585
R130 B.n267 B.n266 585
R131 B.n266 B.n4 585
R132 B.n265 B.n70 585
R133 B.n265 B.n264 585
R134 B.n255 B.n71 585
R135 B.n72 B.n71 585
R136 B.n257 B.n256 585
R137 B.n258 B.n257 585
R138 B.n254 B.n76 585
R139 B.n80 B.n76 585
R140 B.n253 B.n252 585
R141 B.n252 B.n251 585
R142 B.n78 B.n77 585
R143 B.n79 B.n78 585
R144 B.n244 B.n243 585
R145 B.n245 B.n244 585
R146 B.n242 B.n85 585
R147 B.n85 B.n84 585
R148 B.n241 B.n240 585
R149 B.n240 B.n239 585
R150 B.n87 B.n86 585
R151 B.n232 B.n87 585
R152 B.n231 B.n230 585
R153 B.n233 B.n231 585
R154 B.n229 B.n92 585
R155 B.n92 B.n91 585
R156 B.n228 B.n227 585
R157 B.n227 B.n226 585
R158 B.n94 B.n93 585
R159 B.n95 B.n94 585
R160 B.n219 B.n218 585
R161 B.n220 B.n219 585
R162 B.n217 B.n100 585
R163 B.n100 B.n99 585
R164 B.n216 B.n215 585
R165 B.n215 B.n214 585
R166 B.n102 B.n101 585
R167 B.n103 B.n102 585
R168 B.n207 B.n206 585
R169 B.n208 B.n207 585
R170 B.n205 B.n108 585
R171 B.n108 B.n107 585
R172 B.n204 B.n203 585
R173 B.n203 B.n202 585
R174 B.n110 B.n109 585
R175 B.n111 B.n110 585
R176 B.n195 B.n194 585
R177 B.n196 B.n195 585
R178 B.n193 B.n116 585
R179 B.n116 B.n115 585
R180 B.n192 B.n191 585
R181 B.n191 B.n190 585
R182 B.n187 B.n120 585
R183 B.n186 B.n185 585
R184 B.n183 B.n121 585
R185 B.n183 B.n119 585
R186 B.n182 B.n181 585
R187 B.n180 B.n179 585
R188 B.n178 B.n123 585
R189 B.n176 B.n175 585
R190 B.n174 B.n124 585
R191 B.n172 B.n171 585
R192 B.n169 B.n127 585
R193 B.n167 B.n166 585
R194 B.n165 B.n128 585
R195 B.n164 B.n163 585
R196 B.n161 B.n129 585
R197 B.n159 B.n158 585
R198 B.n157 B.n130 585
R199 B.n156 B.n155 585
R200 B.n153 B.n131 585
R201 B.n151 B.n150 585
R202 B.n149 B.n132 585
R203 B.n148 B.n147 585
R204 B.n145 B.n136 585
R205 B.n143 B.n142 585
R206 B.n141 B.n137 585
R207 B.n140 B.n139 585
R208 B.n118 B.n117 585
R209 B.n119 B.n118 585
R210 B.n189 B.n188 585
R211 B.n190 B.n189 585
R212 B.n114 B.n113 585
R213 B.n115 B.n114 585
R214 B.n198 B.n197 585
R215 B.n197 B.n196 585
R216 B.n199 B.n112 585
R217 B.n112 B.n111 585
R218 B.n201 B.n200 585
R219 B.n202 B.n201 585
R220 B.n106 B.n105 585
R221 B.n107 B.n106 585
R222 B.n210 B.n209 585
R223 B.n209 B.n208 585
R224 B.n211 B.n104 585
R225 B.n104 B.n103 585
R226 B.n213 B.n212 585
R227 B.n214 B.n213 585
R228 B.n98 B.n97 585
R229 B.n99 B.n98 585
R230 B.n222 B.n221 585
R231 B.n221 B.n220 585
R232 B.n223 B.n96 585
R233 B.n96 B.n95 585
R234 B.n225 B.n224 585
R235 B.n226 B.n225 585
R236 B.n90 B.n89 585
R237 B.n91 B.n90 585
R238 B.n235 B.n234 585
R239 B.n234 B.n233 585
R240 B.n236 B.n88 585
R241 B.n232 B.n88 585
R242 B.n238 B.n237 585
R243 B.n239 B.n238 585
R244 B.n83 B.n82 585
R245 B.n84 B.n83 585
R246 B.n247 B.n246 585
R247 B.n246 B.n245 585
R248 B.n248 B.n81 585
R249 B.n81 B.n79 585
R250 B.n250 B.n249 585
R251 B.n251 B.n250 585
R252 B.n75 B.n74 585
R253 B.n80 B.n75 585
R254 B.n260 B.n259 585
R255 B.n259 B.n258 585
R256 B.n261 B.n73 585
R257 B.n73 B.n72 585
R258 B.n263 B.n262 585
R259 B.n264 B.n263 585
R260 B.n3 B.n0 585
R261 B.n4 B.n3 585
R262 B.n406 B.n1 585
R263 B.n407 B.n406 585
R264 B.n405 B.n404 585
R265 B.n405 B.n8 585
R266 B.n403 B.n9 585
R267 B.n12 B.n9 585
R268 B.n402 B.n401 585
R269 B.n401 B.n400 585
R270 B.n11 B.n10 585
R271 B.n399 B.n11 585
R272 B.n397 B.n396 585
R273 B.n398 B.n397 585
R274 B.n395 B.n17 585
R275 B.n17 B.n16 585
R276 B.n394 B.n393 585
R277 B.n393 B.n392 585
R278 B.n19 B.n18 585
R279 B.n391 B.n19 585
R280 B.n389 B.n388 585
R281 B.n390 B.n389 585
R282 B.n387 B.n23 585
R283 B.n26 B.n23 585
R284 B.n386 B.n385 585
R285 B.n385 B.n384 585
R286 B.n25 B.n24 585
R287 B.n383 B.n25 585
R288 B.n381 B.n380 585
R289 B.n382 B.n381 585
R290 B.n379 B.n31 585
R291 B.n31 B.n30 585
R292 B.n378 B.n377 585
R293 B.n377 B.n376 585
R294 B.n33 B.n32 585
R295 B.n375 B.n33 585
R296 B.n373 B.n372 585
R297 B.n374 B.n373 585
R298 B.n371 B.n38 585
R299 B.n38 B.n37 585
R300 B.n370 B.n369 585
R301 B.n369 B.n368 585
R302 B.n40 B.n39 585
R303 B.n367 B.n40 585
R304 B.n365 B.n364 585
R305 B.n366 B.n365 585
R306 B.n363 B.n45 585
R307 B.n45 B.n44 585
R308 B.n362 B.n361 585
R309 B.n361 B.n360 585
R310 B.n47 B.n46 585
R311 B.n359 B.n47 585
R312 B.n357 B.n356 585
R313 B.n358 B.n357 585
R314 B.n410 B.n409 585
R315 B.n408 B.n2 585
R316 B.n357 B.n52 511.721
R317 B.n304 B.n50 511.721
R318 B.n191 B.n118 511.721
R319 B.n189 B.n120 511.721
R320 B.n57 B.t13 276.5
R321 B.n63 B.t16 276.5
R322 B.n133 B.t7 276.5
R323 B.n125 B.t10 276.5
R324 B.n305 B.n51 256.663
R325 B.n307 B.n51 256.663
R326 B.n313 B.n51 256.663
R327 B.n66 B.n51 256.663
R328 B.n319 B.n51 256.663
R329 B.n325 B.n51 256.663
R330 B.n327 B.n51 256.663
R331 B.n333 B.n51 256.663
R332 B.n335 B.n51 256.663
R333 B.n342 B.n51 256.663
R334 B.n344 B.n51 256.663
R335 B.n350 B.n51 256.663
R336 B.n352 B.n51 256.663
R337 B.n184 B.n119 256.663
R338 B.n122 B.n119 256.663
R339 B.n177 B.n119 256.663
R340 B.n170 B.n119 256.663
R341 B.n168 B.n119 256.663
R342 B.n162 B.n119 256.663
R343 B.n160 B.n119 256.663
R344 B.n154 B.n119 256.663
R345 B.n152 B.n119 256.663
R346 B.n146 B.n119 256.663
R347 B.n144 B.n119 256.663
R348 B.n138 B.n119 256.663
R349 B.n412 B.n411 256.663
R350 B.n58 B.t14 236.355
R351 B.n64 B.t17 236.355
R352 B.n134 B.t6 236.355
R353 B.n126 B.t9 236.355
R354 B.n190 B.n119 211.363
R355 B.n358 B.n51 211.363
R356 B.n57 B.t11 207.84
R357 B.n63 B.t15 207.84
R358 B.n133 B.t4 207.84
R359 B.n125 B.t8 207.84
R360 B.n353 B.n351 163.367
R361 B.n349 B.n54 163.367
R362 B.n345 B.n343 163.367
R363 B.n341 B.n56 163.367
R364 B.n336 B.n334 163.367
R365 B.n332 B.n60 163.367
R366 B.n328 B.n326 163.367
R367 B.n324 B.n62 163.367
R368 B.n320 B.n318 163.367
R369 B.n315 B.n314 163.367
R370 B.n312 B.n68 163.367
R371 B.n308 B.n306 163.367
R372 B.n191 B.n116 163.367
R373 B.n195 B.n116 163.367
R374 B.n195 B.n110 163.367
R375 B.n203 B.n110 163.367
R376 B.n203 B.n108 163.367
R377 B.n207 B.n108 163.367
R378 B.n207 B.n102 163.367
R379 B.n215 B.n102 163.367
R380 B.n215 B.n100 163.367
R381 B.n219 B.n100 163.367
R382 B.n219 B.n94 163.367
R383 B.n227 B.n94 163.367
R384 B.n227 B.n92 163.367
R385 B.n231 B.n92 163.367
R386 B.n231 B.n87 163.367
R387 B.n240 B.n87 163.367
R388 B.n240 B.n85 163.367
R389 B.n244 B.n85 163.367
R390 B.n244 B.n78 163.367
R391 B.n252 B.n78 163.367
R392 B.n252 B.n76 163.367
R393 B.n257 B.n76 163.367
R394 B.n257 B.n71 163.367
R395 B.n265 B.n71 163.367
R396 B.n266 B.n265 163.367
R397 B.n266 B.n5 163.367
R398 B.n6 B.n5 163.367
R399 B.n7 B.n6 163.367
R400 B.n272 B.n7 163.367
R401 B.n273 B.n272 163.367
R402 B.n273 B.n13 163.367
R403 B.n14 B.n13 163.367
R404 B.n15 B.n14 163.367
R405 B.n278 B.n15 163.367
R406 B.n278 B.n20 163.367
R407 B.n21 B.n20 163.367
R408 B.n22 B.n21 163.367
R409 B.n283 B.n22 163.367
R410 B.n283 B.n27 163.367
R411 B.n28 B.n27 163.367
R412 B.n29 B.n28 163.367
R413 B.n288 B.n29 163.367
R414 B.n288 B.n34 163.367
R415 B.n35 B.n34 163.367
R416 B.n36 B.n35 163.367
R417 B.n293 B.n36 163.367
R418 B.n293 B.n41 163.367
R419 B.n42 B.n41 163.367
R420 B.n43 B.n42 163.367
R421 B.n298 B.n43 163.367
R422 B.n298 B.n48 163.367
R423 B.n49 B.n48 163.367
R424 B.n50 B.n49 163.367
R425 B.n185 B.n183 163.367
R426 B.n183 B.n182 163.367
R427 B.n179 B.n178 163.367
R428 B.n176 B.n124 163.367
R429 B.n171 B.n169 163.367
R430 B.n167 B.n128 163.367
R431 B.n163 B.n161 163.367
R432 B.n159 B.n130 163.367
R433 B.n155 B.n153 163.367
R434 B.n151 B.n132 163.367
R435 B.n147 B.n145 163.367
R436 B.n143 B.n137 163.367
R437 B.n139 B.n118 163.367
R438 B.n189 B.n114 163.367
R439 B.n197 B.n114 163.367
R440 B.n197 B.n112 163.367
R441 B.n201 B.n112 163.367
R442 B.n201 B.n106 163.367
R443 B.n209 B.n106 163.367
R444 B.n209 B.n104 163.367
R445 B.n213 B.n104 163.367
R446 B.n213 B.n98 163.367
R447 B.n221 B.n98 163.367
R448 B.n221 B.n96 163.367
R449 B.n225 B.n96 163.367
R450 B.n225 B.n90 163.367
R451 B.n234 B.n90 163.367
R452 B.n234 B.n88 163.367
R453 B.n238 B.n88 163.367
R454 B.n238 B.n83 163.367
R455 B.n246 B.n83 163.367
R456 B.n246 B.n81 163.367
R457 B.n250 B.n81 163.367
R458 B.n250 B.n75 163.367
R459 B.n259 B.n75 163.367
R460 B.n259 B.n73 163.367
R461 B.n263 B.n73 163.367
R462 B.n263 B.n3 163.367
R463 B.n410 B.n3 163.367
R464 B.n406 B.n2 163.367
R465 B.n406 B.n405 163.367
R466 B.n405 B.n9 163.367
R467 B.n401 B.n9 163.367
R468 B.n401 B.n11 163.367
R469 B.n397 B.n11 163.367
R470 B.n397 B.n17 163.367
R471 B.n393 B.n17 163.367
R472 B.n393 B.n19 163.367
R473 B.n389 B.n19 163.367
R474 B.n389 B.n23 163.367
R475 B.n385 B.n23 163.367
R476 B.n385 B.n25 163.367
R477 B.n381 B.n25 163.367
R478 B.n381 B.n31 163.367
R479 B.n377 B.n31 163.367
R480 B.n377 B.n33 163.367
R481 B.n373 B.n33 163.367
R482 B.n373 B.n38 163.367
R483 B.n369 B.n38 163.367
R484 B.n369 B.n40 163.367
R485 B.n365 B.n40 163.367
R486 B.n365 B.n45 163.367
R487 B.n361 B.n45 163.367
R488 B.n361 B.n47 163.367
R489 B.n357 B.n47 163.367
R490 B.n190 B.n115 124.98
R491 B.n196 B.n115 124.98
R492 B.n196 B.n111 124.98
R493 B.n202 B.n111 124.98
R494 B.n202 B.n107 124.98
R495 B.n208 B.n107 124.98
R496 B.n214 B.n103 124.98
R497 B.n214 B.n99 124.98
R498 B.n220 B.n99 124.98
R499 B.n220 B.n95 124.98
R500 B.n226 B.n95 124.98
R501 B.n226 B.n91 124.98
R502 B.n233 B.n91 124.98
R503 B.n233 B.n232 124.98
R504 B.n239 B.n84 124.98
R505 B.n245 B.n84 124.98
R506 B.n245 B.n79 124.98
R507 B.n251 B.n79 124.98
R508 B.n251 B.n80 124.98
R509 B.n258 B.n72 124.98
R510 B.n264 B.n72 124.98
R511 B.n264 B.n4 124.98
R512 B.n409 B.n4 124.98
R513 B.n409 B.n408 124.98
R514 B.n408 B.n407 124.98
R515 B.n407 B.n8 124.98
R516 B.n12 B.n8 124.98
R517 B.n400 B.n12 124.98
R518 B.n399 B.n398 124.98
R519 B.n398 B.n16 124.98
R520 B.n392 B.n16 124.98
R521 B.n392 B.n391 124.98
R522 B.n391 B.n390 124.98
R523 B.n384 B.n26 124.98
R524 B.n384 B.n383 124.98
R525 B.n383 B.n382 124.98
R526 B.n382 B.n30 124.98
R527 B.n376 B.n30 124.98
R528 B.n376 B.n375 124.98
R529 B.n375 B.n374 124.98
R530 B.n374 B.n37 124.98
R531 B.n368 B.n367 124.98
R532 B.n367 B.n366 124.98
R533 B.n366 B.n44 124.98
R534 B.n360 B.n44 124.98
R535 B.n360 B.n359 124.98
R536 B.n359 B.n358 124.98
R537 B.n80 B.t1 106.6
R538 B.t2 B.n399 106.6
R539 B.n232 B.t3 95.5728
R540 B.n26 B.t0 95.5728
R541 B.n352 B.n52 71.676
R542 B.n351 B.n350 71.676
R543 B.n344 B.n54 71.676
R544 B.n343 B.n342 71.676
R545 B.n335 B.n56 71.676
R546 B.n334 B.n333 71.676
R547 B.n327 B.n60 71.676
R548 B.n326 B.n325 71.676
R549 B.n319 B.n62 71.676
R550 B.n318 B.n66 71.676
R551 B.n314 B.n313 71.676
R552 B.n307 B.n68 71.676
R553 B.n306 B.n305 71.676
R554 B.n305 B.n304 71.676
R555 B.n308 B.n307 71.676
R556 B.n313 B.n312 71.676
R557 B.n315 B.n66 71.676
R558 B.n320 B.n319 71.676
R559 B.n325 B.n324 71.676
R560 B.n328 B.n327 71.676
R561 B.n333 B.n332 71.676
R562 B.n336 B.n335 71.676
R563 B.n342 B.n341 71.676
R564 B.n345 B.n344 71.676
R565 B.n350 B.n349 71.676
R566 B.n353 B.n352 71.676
R567 B.n184 B.n120 71.676
R568 B.n182 B.n122 71.676
R569 B.n178 B.n177 71.676
R570 B.n170 B.n124 71.676
R571 B.n169 B.n168 71.676
R572 B.n162 B.n128 71.676
R573 B.n161 B.n160 71.676
R574 B.n154 B.n130 71.676
R575 B.n153 B.n152 71.676
R576 B.n146 B.n132 71.676
R577 B.n145 B.n144 71.676
R578 B.n138 B.n137 71.676
R579 B.n185 B.n184 71.676
R580 B.n179 B.n122 71.676
R581 B.n177 B.n176 71.676
R582 B.n171 B.n170 71.676
R583 B.n168 B.n167 71.676
R584 B.n163 B.n162 71.676
R585 B.n160 B.n159 71.676
R586 B.n155 B.n154 71.676
R587 B.n152 B.n151 71.676
R588 B.n147 B.n146 71.676
R589 B.n144 B.n143 71.676
R590 B.n139 B.n138 71.676
R591 B.n411 B.n410 71.676
R592 B.n411 B.n2 71.676
R593 B.t5 B.n103 66.1659
R594 B.t12 B.n37 66.1659
R595 B.n339 B.n58 59.5399
R596 B.n65 B.n64 59.5399
R597 B.n135 B.n134 59.5399
R598 B.n173 B.n126 59.5399
R599 B.n208 B.t5 58.8142
R600 B.n368 B.t12 58.8142
R601 B.n58 B.n57 40.146
R602 B.n64 B.n63 40.146
R603 B.n134 B.n133 40.146
R604 B.n126 B.n125 40.146
R605 B.n188 B.n187 33.2493
R606 B.n192 B.n117 33.2493
R607 B.n303 B.n302 33.2493
R608 B.n356 B.n355 33.2493
R609 B.n239 B.t3 29.4073
R610 B.n390 B.t0 29.4073
R611 B.n258 B.t1 18.3798
R612 B.n400 B.t2 18.3798
R613 B B.n412 18.0485
R614 B.n188 B.n113 10.6151
R615 B.n198 B.n113 10.6151
R616 B.n199 B.n198 10.6151
R617 B.n200 B.n199 10.6151
R618 B.n200 B.n105 10.6151
R619 B.n210 B.n105 10.6151
R620 B.n211 B.n210 10.6151
R621 B.n212 B.n211 10.6151
R622 B.n212 B.n97 10.6151
R623 B.n222 B.n97 10.6151
R624 B.n223 B.n222 10.6151
R625 B.n224 B.n223 10.6151
R626 B.n224 B.n89 10.6151
R627 B.n235 B.n89 10.6151
R628 B.n236 B.n235 10.6151
R629 B.n237 B.n236 10.6151
R630 B.n237 B.n82 10.6151
R631 B.n247 B.n82 10.6151
R632 B.n248 B.n247 10.6151
R633 B.n249 B.n248 10.6151
R634 B.n249 B.n74 10.6151
R635 B.n260 B.n74 10.6151
R636 B.n261 B.n260 10.6151
R637 B.n262 B.n261 10.6151
R638 B.n262 B.n0 10.6151
R639 B.n187 B.n186 10.6151
R640 B.n186 B.n121 10.6151
R641 B.n181 B.n121 10.6151
R642 B.n181 B.n180 10.6151
R643 B.n180 B.n123 10.6151
R644 B.n175 B.n123 10.6151
R645 B.n175 B.n174 10.6151
R646 B.n172 B.n127 10.6151
R647 B.n166 B.n127 10.6151
R648 B.n166 B.n165 10.6151
R649 B.n165 B.n164 10.6151
R650 B.n164 B.n129 10.6151
R651 B.n158 B.n129 10.6151
R652 B.n158 B.n157 10.6151
R653 B.n157 B.n156 10.6151
R654 B.n156 B.n131 10.6151
R655 B.n150 B.n149 10.6151
R656 B.n149 B.n148 10.6151
R657 B.n148 B.n136 10.6151
R658 B.n142 B.n136 10.6151
R659 B.n142 B.n141 10.6151
R660 B.n141 B.n140 10.6151
R661 B.n140 B.n117 10.6151
R662 B.n193 B.n192 10.6151
R663 B.n194 B.n193 10.6151
R664 B.n194 B.n109 10.6151
R665 B.n204 B.n109 10.6151
R666 B.n205 B.n204 10.6151
R667 B.n206 B.n205 10.6151
R668 B.n206 B.n101 10.6151
R669 B.n216 B.n101 10.6151
R670 B.n217 B.n216 10.6151
R671 B.n218 B.n217 10.6151
R672 B.n218 B.n93 10.6151
R673 B.n228 B.n93 10.6151
R674 B.n229 B.n228 10.6151
R675 B.n230 B.n229 10.6151
R676 B.n230 B.n86 10.6151
R677 B.n241 B.n86 10.6151
R678 B.n242 B.n241 10.6151
R679 B.n243 B.n242 10.6151
R680 B.n243 B.n77 10.6151
R681 B.n253 B.n77 10.6151
R682 B.n254 B.n253 10.6151
R683 B.n256 B.n254 10.6151
R684 B.n256 B.n255 10.6151
R685 B.n255 B.n70 10.6151
R686 B.n267 B.n70 10.6151
R687 B.n268 B.n267 10.6151
R688 B.n269 B.n268 10.6151
R689 B.n270 B.n269 10.6151
R690 B.n271 B.n270 10.6151
R691 B.n274 B.n271 10.6151
R692 B.n275 B.n274 10.6151
R693 B.n276 B.n275 10.6151
R694 B.n277 B.n276 10.6151
R695 B.n279 B.n277 10.6151
R696 B.n280 B.n279 10.6151
R697 B.n281 B.n280 10.6151
R698 B.n282 B.n281 10.6151
R699 B.n284 B.n282 10.6151
R700 B.n285 B.n284 10.6151
R701 B.n286 B.n285 10.6151
R702 B.n287 B.n286 10.6151
R703 B.n289 B.n287 10.6151
R704 B.n290 B.n289 10.6151
R705 B.n291 B.n290 10.6151
R706 B.n292 B.n291 10.6151
R707 B.n294 B.n292 10.6151
R708 B.n295 B.n294 10.6151
R709 B.n296 B.n295 10.6151
R710 B.n297 B.n296 10.6151
R711 B.n299 B.n297 10.6151
R712 B.n300 B.n299 10.6151
R713 B.n301 B.n300 10.6151
R714 B.n302 B.n301 10.6151
R715 B.n404 B.n1 10.6151
R716 B.n404 B.n403 10.6151
R717 B.n403 B.n402 10.6151
R718 B.n402 B.n10 10.6151
R719 B.n396 B.n10 10.6151
R720 B.n396 B.n395 10.6151
R721 B.n395 B.n394 10.6151
R722 B.n394 B.n18 10.6151
R723 B.n388 B.n18 10.6151
R724 B.n388 B.n387 10.6151
R725 B.n387 B.n386 10.6151
R726 B.n386 B.n24 10.6151
R727 B.n380 B.n24 10.6151
R728 B.n380 B.n379 10.6151
R729 B.n379 B.n378 10.6151
R730 B.n378 B.n32 10.6151
R731 B.n372 B.n32 10.6151
R732 B.n372 B.n371 10.6151
R733 B.n371 B.n370 10.6151
R734 B.n370 B.n39 10.6151
R735 B.n364 B.n39 10.6151
R736 B.n364 B.n363 10.6151
R737 B.n363 B.n362 10.6151
R738 B.n362 B.n46 10.6151
R739 B.n356 B.n46 10.6151
R740 B.n355 B.n354 10.6151
R741 B.n354 B.n53 10.6151
R742 B.n348 B.n53 10.6151
R743 B.n348 B.n347 10.6151
R744 B.n347 B.n346 10.6151
R745 B.n346 B.n55 10.6151
R746 B.n340 B.n55 10.6151
R747 B.n338 B.n337 10.6151
R748 B.n337 B.n59 10.6151
R749 B.n331 B.n59 10.6151
R750 B.n331 B.n330 10.6151
R751 B.n330 B.n329 10.6151
R752 B.n329 B.n61 10.6151
R753 B.n323 B.n61 10.6151
R754 B.n323 B.n322 10.6151
R755 B.n322 B.n321 10.6151
R756 B.n317 B.n316 10.6151
R757 B.n316 B.n67 10.6151
R758 B.n311 B.n67 10.6151
R759 B.n311 B.n310 10.6151
R760 B.n310 B.n309 10.6151
R761 B.n309 B.n69 10.6151
R762 B.n303 B.n69 10.6151
R763 B.n174 B.n173 9.36635
R764 B.n150 B.n135 9.36635
R765 B.n340 B.n339 9.36635
R766 B.n317 B.n65 9.36635
R767 B.n412 B.n0 8.11757
R768 B.n412 B.n1 8.11757
R769 B.n173 B.n172 1.24928
R770 B.n135 B.n131 1.24928
R771 B.n339 B.n338 1.24928
R772 B.n321 B.n65 1.24928
R773 VN.n0 VN.t0 45.4791
R774 VN.n1 VN.t1 45.4791
R775 VN.n0 VN.t3 45.054
R776 VN.n1 VN.t2 45.054
R777 VN VN.n1 44.8318
R778 VN VN.n0 9.46438
R779 VDD2.n2 VDD2.n0 265.678
R780 VDD2.n2 VDD2.n1 235.998
R781 VDD2.n1 VDD2.t1 27.8878
R782 VDD2.n1 VDD2.t2 27.8878
R783 VDD2.n0 VDD2.t3 27.8878
R784 VDD2.n0 VDD2.t0 27.8878
R785 VDD2 VDD2.n2 0.0586897
C0 VN VP 3.49149f
C1 VDD1 VN 0.155538f
C2 VTAIL VDD2 2.303f
C3 VTAIL VP 1.08421f
C4 VP VDD2 0.348357f
C5 VDD1 VTAIL 2.25456f
C6 VDD1 VDD2 0.817353f
C7 VDD1 VP 0.750859f
C8 VTAIL VN 1.07011f
C9 VN VDD2 0.560162f
C10 VDD2 B 2.374579f
C11 VDD1 B 4.55754f
C12 VTAIL B 2.515015f
C13 VN B 7.640611f
C14 VP B 6.088122f
C15 VDD2.t3 B 0.013955f
C16 VDD2.t0 B 0.013955f
C17 VDD2.n0 B 0.111402f
C18 VDD2.t1 B 0.013955f
C19 VDD2.t2 B 0.013955f
C20 VDD2.n1 B 0.034401f
C21 VDD2.n2 B 1.95001f
C22 VN.t0 B 0.221407f
C23 VN.t3 B 0.219608f
C24 VN.n0 B 0.146561f
C25 VN.t1 B 0.221407f
C26 VN.t2 B 0.219608f
C27 VN.n1 B 1.05121f
C28 VTAIL.t2 B 0.06727f
C29 VTAIL.n0 B 0.167548f
C30 VTAIL.t6 B 0.06727f
C31 VTAIL.n1 B 0.240202f
C32 VTAIL.t4 B 0.06727f
C33 VTAIL.n2 B 0.775259f
C34 VTAIL.t3 B 0.06727f
C35 VTAIL.n3 B 0.775259f
C36 VTAIL.t1 B 0.06727f
C37 VTAIL.n4 B 0.240202f
C38 VTAIL.t7 B 0.06727f
C39 VTAIL.n5 B 0.240202f
C40 VTAIL.t5 B 0.06727f
C41 VTAIL.n6 B 0.775259f
C42 VTAIL.t0 B 0.06727f
C43 VTAIL.n7 B 0.692468f
C44 VDD1.t3 B 0.013419f
C45 VDD1.t2 B 0.013419f
C46 VDD1.n0 B 0.033132f
C47 VDD1.t0 B 0.013419f
C48 VDD1.t1 B 0.013419f
C49 VDD1.n1 B 0.113846f
C50 VP.n0 B 0.031292f
C51 VP.t1 B 0.057475f
C52 VP.n1 B 0.025296f
C53 VP.n2 B 0.031292f
C54 VP.t3 B 0.057475f
C55 VP.t0 B 0.224189f
C56 VP.t2 B 0.222368f
C57 VP.n3 B 1.04594f
C58 VP.n4 B 1.21711f
C59 VP.n5 B 0.129889f
C60 VP.n6 B 0.031541f
C61 VP.n7 B 0.062192f
C62 VP.n8 B 0.031292f
C63 VP.n9 B 0.031292f
C64 VP.n10 B 0.031292f
C65 VP.n11 B 0.062192f
C66 VP.n12 B 0.031541f
C67 VP.n13 B 0.129889f
C68 VP.n14 B 0.033418f
.ends

