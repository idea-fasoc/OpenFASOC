* NGSPICE file created from diff_pair_sample_0676.ext - technology: sky130A

.subckt diff_pair_sample_0676 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t2 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X1 B.t11 B.t9 B.t10 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=0 ps=0 w=10.94 l=3.95
X2 VDD2.t9 VN.t0 VTAIL.t7 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=1.8051 ps=11.27 w=10.94 l=3.95
X3 VDD1.t7 VP.t1 VTAIL.t16 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=1.8051 ps=11.27 w=10.94 l=3.95
X4 VTAIL.t15 VP.t2 VDD1.t8 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X5 VDD2.t8 VN.t1 VTAIL.t3 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X6 B.t8 B.t6 B.t7 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=0 ps=0 w=10.94 l=3.95
X7 VDD1.t4 VP.t3 VTAIL.t14 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X8 VTAIL.t4 VN.t2 VDD2.t7 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X9 VDD1.t1 VP.t4 VTAIL.t13 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=4.2666 ps=22.66 w=10.94 l=3.95
X10 VDD2.t6 VN.t3 VTAIL.t6 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=4.2666 ps=22.66 w=10.94 l=3.95
X11 VTAIL.t12 VP.t5 VDD1.t9 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X12 VDD2.t5 VN.t4 VTAIL.t19 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X13 VDD2.t4 VN.t5 VTAIL.t18 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=4.2666 ps=22.66 w=10.94 l=3.95
X14 VTAIL.t11 VP.t6 VDD1.t0 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X15 VDD2.t3 VN.t6 VTAIL.t2 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=1.8051 ps=11.27 w=10.94 l=3.95
X16 VDD1.t3 VP.t7 VTAIL.t10 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=1.8051 ps=11.27 w=10.94 l=3.95
X17 VTAIL.t5 VN.t7 VDD2.t2 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X18 VDD1.t6 VP.t8 VTAIL.t9 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X19 VTAIL.t1 VN.t8 VDD2.t1 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
X20 B.t5 B.t3 B.t4 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=0 ps=0 w=10.94 l=3.95
X21 VDD1.t5 VP.t9 VTAIL.t8 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=4.2666 ps=22.66 w=10.94 l=3.95
X22 B.t2 B.t0 B.t1 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=4.2666 pd=22.66 as=0 ps=0 w=10.94 l=3.95
X23 VTAIL.t0 VN.t9 VDD2.t0 w_n6106_n3156# sky130_fd_pr__pfet_01v8 ad=1.8051 pd=11.27 as=1.8051 ps=11.27 w=10.94 l=3.95
R0 VP.n35 VP.n32 161.3
R1 VP.n37 VP.n36 161.3
R2 VP.n38 VP.n31 161.3
R3 VP.n40 VP.n39 161.3
R4 VP.n41 VP.n30 161.3
R5 VP.n43 VP.n42 161.3
R6 VP.n44 VP.n29 161.3
R7 VP.n46 VP.n45 161.3
R8 VP.n47 VP.n28 161.3
R9 VP.n49 VP.n48 161.3
R10 VP.n50 VP.n27 161.3
R11 VP.n52 VP.n51 161.3
R12 VP.n53 VP.n26 161.3
R13 VP.n55 VP.n54 161.3
R14 VP.n56 VP.n25 161.3
R15 VP.n58 VP.n57 161.3
R16 VP.n59 VP.n24 161.3
R17 VP.n62 VP.n61 161.3
R18 VP.n63 VP.n23 161.3
R19 VP.n65 VP.n64 161.3
R20 VP.n66 VP.n22 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n69 VP.n21 161.3
R23 VP.n71 VP.n70 161.3
R24 VP.n72 VP.n20 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n131 VP.n130 161.3
R27 VP.n129 VP.n1 161.3
R28 VP.n128 VP.n127 161.3
R29 VP.n126 VP.n2 161.3
R30 VP.n125 VP.n124 161.3
R31 VP.n123 VP.n3 161.3
R32 VP.n122 VP.n121 161.3
R33 VP.n120 VP.n4 161.3
R34 VP.n119 VP.n118 161.3
R35 VP.n116 VP.n5 161.3
R36 VP.n115 VP.n114 161.3
R37 VP.n113 VP.n6 161.3
R38 VP.n112 VP.n111 161.3
R39 VP.n110 VP.n7 161.3
R40 VP.n109 VP.n108 161.3
R41 VP.n107 VP.n8 161.3
R42 VP.n106 VP.n105 161.3
R43 VP.n104 VP.n9 161.3
R44 VP.n103 VP.n102 161.3
R45 VP.n101 VP.n10 161.3
R46 VP.n100 VP.n99 161.3
R47 VP.n98 VP.n11 161.3
R48 VP.n97 VP.n96 161.3
R49 VP.n95 VP.n12 161.3
R50 VP.n94 VP.n93 161.3
R51 VP.n92 VP.n13 161.3
R52 VP.n90 VP.n89 161.3
R53 VP.n88 VP.n14 161.3
R54 VP.n87 VP.n86 161.3
R55 VP.n85 VP.n15 161.3
R56 VP.n84 VP.n83 161.3
R57 VP.n82 VP.n16 161.3
R58 VP.n81 VP.n80 161.3
R59 VP.n79 VP.n17 161.3
R60 VP.n78 VP.n77 161.3
R61 VP.n33 VP.t1 99.6588
R62 VP.n76 VP.n18 87.2945
R63 VP.n132 VP.n0 87.2945
R64 VP.n75 VP.n19 87.2945
R65 VP.n104 VP.t3 66.7483
R66 VP.n18 VP.t7 66.7483
R67 VP.n91 VP.t6 66.7483
R68 VP.n117 VP.t2 66.7483
R69 VP.n0 VP.t9 66.7483
R70 VP.n47 VP.t8 66.7483
R71 VP.n19 VP.t4 66.7483
R72 VP.n60 VP.t0 66.7483
R73 VP.n34 VP.t5 66.7483
R74 VP.n34 VP.n33 61.6104
R75 VP.n76 VP.n75 59.742
R76 VP.n98 VP.n97 54.1398
R77 VP.n111 VP.n110 54.1398
R78 VP.n54 VP.n53 54.1398
R79 VP.n41 VP.n40 54.1398
R80 VP.n85 VP.n84 48.3272
R81 VP.n124 VP.n123 48.3272
R82 VP.n67 VP.n66 48.3272
R83 VP.n84 VP.n16 32.8269
R84 VP.n124 VP.n2 32.8269
R85 VP.n67 VP.n21 32.8269
R86 VP.n99 VP.n98 27.0143
R87 VP.n110 VP.n109 27.0143
R88 VP.n53 VP.n52 27.0143
R89 VP.n42 VP.n41 27.0143
R90 VP.n79 VP.n78 24.5923
R91 VP.n80 VP.n79 24.5923
R92 VP.n80 VP.n16 24.5923
R93 VP.n86 VP.n85 24.5923
R94 VP.n86 VP.n14 24.5923
R95 VP.n90 VP.n14 24.5923
R96 VP.n93 VP.n92 24.5923
R97 VP.n93 VP.n12 24.5923
R98 VP.n97 VP.n12 24.5923
R99 VP.n99 VP.n10 24.5923
R100 VP.n103 VP.n10 24.5923
R101 VP.n104 VP.n103 24.5923
R102 VP.n105 VP.n104 24.5923
R103 VP.n105 VP.n8 24.5923
R104 VP.n109 VP.n8 24.5923
R105 VP.n111 VP.n6 24.5923
R106 VP.n115 VP.n6 24.5923
R107 VP.n116 VP.n115 24.5923
R108 VP.n118 VP.n4 24.5923
R109 VP.n122 VP.n4 24.5923
R110 VP.n123 VP.n122 24.5923
R111 VP.n128 VP.n2 24.5923
R112 VP.n129 VP.n128 24.5923
R113 VP.n130 VP.n129 24.5923
R114 VP.n71 VP.n21 24.5923
R115 VP.n72 VP.n71 24.5923
R116 VP.n73 VP.n72 24.5923
R117 VP.n54 VP.n25 24.5923
R118 VP.n58 VP.n25 24.5923
R119 VP.n59 VP.n58 24.5923
R120 VP.n61 VP.n23 24.5923
R121 VP.n65 VP.n23 24.5923
R122 VP.n66 VP.n65 24.5923
R123 VP.n42 VP.n29 24.5923
R124 VP.n46 VP.n29 24.5923
R125 VP.n47 VP.n46 24.5923
R126 VP.n48 VP.n47 24.5923
R127 VP.n48 VP.n27 24.5923
R128 VP.n52 VP.n27 24.5923
R129 VP.n36 VP.n35 24.5923
R130 VP.n36 VP.n31 24.5923
R131 VP.n40 VP.n31 24.5923
R132 VP.n92 VP.n91 13.7719
R133 VP.n117 VP.n116 13.7719
R134 VP.n60 VP.n59 13.7719
R135 VP.n35 VP.n34 13.7719
R136 VP.n91 VP.n90 10.8209
R137 VP.n118 VP.n117 10.8209
R138 VP.n61 VP.n60 10.8209
R139 VP.n78 VP.n18 2.95152
R140 VP.n130 VP.n0 2.95152
R141 VP.n73 VP.n19 2.95152
R142 VP.n33 VP.n32 2.45424
R143 VP.n75 VP.n74 0.354861
R144 VP.n77 VP.n76 0.354861
R145 VP.n132 VP.n131 0.354861
R146 VP VP.n132 0.267071
R147 VP.n37 VP.n32 0.189894
R148 VP.n38 VP.n37 0.189894
R149 VP.n39 VP.n38 0.189894
R150 VP.n39 VP.n30 0.189894
R151 VP.n43 VP.n30 0.189894
R152 VP.n44 VP.n43 0.189894
R153 VP.n45 VP.n44 0.189894
R154 VP.n45 VP.n28 0.189894
R155 VP.n49 VP.n28 0.189894
R156 VP.n50 VP.n49 0.189894
R157 VP.n51 VP.n50 0.189894
R158 VP.n51 VP.n26 0.189894
R159 VP.n55 VP.n26 0.189894
R160 VP.n56 VP.n55 0.189894
R161 VP.n57 VP.n56 0.189894
R162 VP.n57 VP.n24 0.189894
R163 VP.n62 VP.n24 0.189894
R164 VP.n63 VP.n62 0.189894
R165 VP.n64 VP.n63 0.189894
R166 VP.n64 VP.n22 0.189894
R167 VP.n68 VP.n22 0.189894
R168 VP.n69 VP.n68 0.189894
R169 VP.n70 VP.n69 0.189894
R170 VP.n70 VP.n20 0.189894
R171 VP.n74 VP.n20 0.189894
R172 VP.n77 VP.n17 0.189894
R173 VP.n81 VP.n17 0.189894
R174 VP.n82 VP.n81 0.189894
R175 VP.n83 VP.n82 0.189894
R176 VP.n83 VP.n15 0.189894
R177 VP.n87 VP.n15 0.189894
R178 VP.n88 VP.n87 0.189894
R179 VP.n89 VP.n88 0.189894
R180 VP.n89 VP.n13 0.189894
R181 VP.n94 VP.n13 0.189894
R182 VP.n95 VP.n94 0.189894
R183 VP.n96 VP.n95 0.189894
R184 VP.n96 VP.n11 0.189894
R185 VP.n100 VP.n11 0.189894
R186 VP.n101 VP.n100 0.189894
R187 VP.n102 VP.n101 0.189894
R188 VP.n102 VP.n9 0.189894
R189 VP.n106 VP.n9 0.189894
R190 VP.n107 VP.n106 0.189894
R191 VP.n108 VP.n107 0.189894
R192 VP.n108 VP.n7 0.189894
R193 VP.n112 VP.n7 0.189894
R194 VP.n113 VP.n112 0.189894
R195 VP.n114 VP.n113 0.189894
R196 VP.n114 VP.n5 0.189894
R197 VP.n119 VP.n5 0.189894
R198 VP.n120 VP.n119 0.189894
R199 VP.n121 VP.n120 0.189894
R200 VP.n121 VP.n3 0.189894
R201 VP.n125 VP.n3 0.189894
R202 VP.n126 VP.n125 0.189894
R203 VP.n127 VP.n126 0.189894
R204 VP.n127 VP.n1 0.189894
R205 VP.n131 VP.n1 0.189894
R206 VDD1.n1 VDD1.t7 80.0265
R207 VDD1.n3 VDD1.t3 80.0263
R208 VDD1.n5 VDD1.n4 76.0773
R209 VDD1.n1 VDD1.n0 73.3657
R210 VDD1.n7 VDD1.n6 73.3655
R211 VDD1.n3 VDD1.n2 73.3654
R212 VDD1.n7 VDD1.n5 53.1
R213 VDD1.n6 VDD1.t2 2.97171
R214 VDD1.n6 VDD1.t1 2.97171
R215 VDD1.n0 VDD1.t9 2.97171
R216 VDD1.n0 VDD1.t6 2.97171
R217 VDD1.n4 VDD1.t8 2.97171
R218 VDD1.n4 VDD1.t5 2.97171
R219 VDD1.n2 VDD1.t0 2.97171
R220 VDD1.n2 VDD1.t4 2.97171
R221 VDD1 VDD1.n7 2.70955
R222 VDD1 VDD1.n1 0.981103
R223 VDD1.n5 VDD1.n3 0.867568
R224 VTAIL.n11 VTAIL.t6 59.658
R225 VTAIL.n17 VTAIL.t18 59.6579
R226 VTAIL.n2 VTAIL.t8 59.6579
R227 VTAIL.n16 VTAIL.t13 59.6579
R228 VTAIL.n15 VTAIL.n14 56.6869
R229 VTAIL.n13 VTAIL.n12 56.6869
R230 VTAIL.n10 VTAIL.n9 56.6869
R231 VTAIL.n8 VTAIL.n7 56.6869
R232 VTAIL.n19 VTAIL.n18 56.6866
R233 VTAIL.n1 VTAIL.n0 56.6866
R234 VTAIL.n4 VTAIL.n3 56.6866
R235 VTAIL.n6 VTAIL.n5 56.6866
R236 VTAIL.n8 VTAIL.n6 29.1772
R237 VTAIL.n17 VTAIL.n16 25.4876
R238 VTAIL.n10 VTAIL.n8 3.69016
R239 VTAIL.n11 VTAIL.n10 3.69016
R240 VTAIL.n15 VTAIL.n13 3.69016
R241 VTAIL.n16 VTAIL.n15 3.69016
R242 VTAIL.n6 VTAIL.n4 3.69016
R243 VTAIL.n4 VTAIL.n2 3.69016
R244 VTAIL.n19 VTAIL.n17 3.69016
R245 VTAIL.n18 VTAIL.t3 2.97171
R246 VTAIL.n18 VTAIL.t4 2.97171
R247 VTAIL.n0 VTAIL.t2 2.97171
R248 VTAIL.n0 VTAIL.t0 2.97171
R249 VTAIL.n3 VTAIL.t14 2.97171
R250 VTAIL.n3 VTAIL.t15 2.97171
R251 VTAIL.n5 VTAIL.t10 2.97171
R252 VTAIL.n5 VTAIL.t11 2.97171
R253 VTAIL.n14 VTAIL.t9 2.97171
R254 VTAIL.n14 VTAIL.t17 2.97171
R255 VTAIL.n12 VTAIL.t16 2.97171
R256 VTAIL.n12 VTAIL.t12 2.97171
R257 VTAIL.n9 VTAIL.t19 2.97171
R258 VTAIL.n9 VTAIL.t5 2.97171
R259 VTAIL.n7 VTAIL.t7 2.97171
R260 VTAIL.n7 VTAIL.t1 2.97171
R261 VTAIL VTAIL.n1 2.82593
R262 VTAIL.n13 VTAIL.n11 2.31516
R263 VTAIL.n2 VTAIL.n1 2.31516
R264 VTAIL VTAIL.n19 0.864724
R265 B.n518 B.n175 585
R266 B.n517 B.n516 585
R267 B.n515 B.n176 585
R268 B.n514 B.n513 585
R269 B.n512 B.n177 585
R270 B.n511 B.n510 585
R271 B.n509 B.n178 585
R272 B.n508 B.n507 585
R273 B.n506 B.n179 585
R274 B.n505 B.n504 585
R275 B.n503 B.n180 585
R276 B.n502 B.n501 585
R277 B.n500 B.n181 585
R278 B.n499 B.n498 585
R279 B.n497 B.n182 585
R280 B.n496 B.n495 585
R281 B.n494 B.n183 585
R282 B.n493 B.n492 585
R283 B.n491 B.n184 585
R284 B.n490 B.n489 585
R285 B.n488 B.n185 585
R286 B.n487 B.n486 585
R287 B.n485 B.n186 585
R288 B.n484 B.n483 585
R289 B.n482 B.n187 585
R290 B.n481 B.n480 585
R291 B.n479 B.n188 585
R292 B.n478 B.n477 585
R293 B.n476 B.n189 585
R294 B.n475 B.n474 585
R295 B.n473 B.n190 585
R296 B.n472 B.n471 585
R297 B.n470 B.n191 585
R298 B.n469 B.n468 585
R299 B.n467 B.n192 585
R300 B.n466 B.n465 585
R301 B.n464 B.n193 585
R302 B.n463 B.n462 585
R303 B.n461 B.n194 585
R304 B.n460 B.n459 585
R305 B.n455 B.n195 585
R306 B.n454 B.n453 585
R307 B.n452 B.n196 585
R308 B.n451 B.n450 585
R309 B.n449 B.n197 585
R310 B.n448 B.n447 585
R311 B.n446 B.n198 585
R312 B.n445 B.n444 585
R313 B.n442 B.n199 585
R314 B.n441 B.n440 585
R315 B.n439 B.n202 585
R316 B.n438 B.n437 585
R317 B.n436 B.n203 585
R318 B.n435 B.n434 585
R319 B.n433 B.n204 585
R320 B.n432 B.n431 585
R321 B.n430 B.n205 585
R322 B.n429 B.n428 585
R323 B.n427 B.n206 585
R324 B.n426 B.n425 585
R325 B.n424 B.n207 585
R326 B.n423 B.n422 585
R327 B.n421 B.n208 585
R328 B.n420 B.n419 585
R329 B.n418 B.n209 585
R330 B.n417 B.n416 585
R331 B.n415 B.n210 585
R332 B.n414 B.n413 585
R333 B.n412 B.n211 585
R334 B.n411 B.n410 585
R335 B.n409 B.n212 585
R336 B.n408 B.n407 585
R337 B.n406 B.n213 585
R338 B.n405 B.n404 585
R339 B.n403 B.n214 585
R340 B.n402 B.n401 585
R341 B.n400 B.n215 585
R342 B.n399 B.n398 585
R343 B.n397 B.n216 585
R344 B.n396 B.n395 585
R345 B.n394 B.n217 585
R346 B.n393 B.n392 585
R347 B.n391 B.n218 585
R348 B.n390 B.n389 585
R349 B.n388 B.n219 585
R350 B.n387 B.n386 585
R351 B.n385 B.n220 585
R352 B.n520 B.n519 585
R353 B.n521 B.n174 585
R354 B.n523 B.n522 585
R355 B.n524 B.n173 585
R356 B.n526 B.n525 585
R357 B.n527 B.n172 585
R358 B.n529 B.n528 585
R359 B.n530 B.n171 585
R360 B.n532 B.n531 585
R361 B.n533 B.n170 585
R362 B.n535 B.n534 585
R363 B.n536 B.n169 585
R364 B.n538 B.n537 585
R365 B.n539 B.n168 585
R366 B.n541 B.n540 585
R367 B.n542 B.n167 585
R368 B.n544 B.n543 585
R369 B.n545 B.n166 585
R370 B.n547 B.n546 585
R371 B.n548 B.n165 585
R372 B.n550 B.n549 585
R373 B.n551 B.n164 585
R374 B.n553 B.n552 585
R375 B.n554 B.n163 585
R376 B.n556 B.n555 585
R377 B.n557 B.n162 585
R378 B.n559 B.n558 585
R379 B.n560 B.n161 585
R380 B.n562 B.n561 585
R381 B.n563 B.n160 585
R382 B.n565 B.n564 585
R383 B.n566 B.n159 585
R384 B.n568 B.n567 585
R385 B.n569 B.n158 585
R386 B.n571 B.n570 585
R387 B.n572 B.n157 585
R388 B.n574 B.n573 585
R389 B.n575 B.n156 585
R390 B.n577 B.n576 585
R391 B.n578 B.n155 585
R392 B.n580 B.n579 585
R393 B.n581 B.n154 585
R394 B.n583 B.n582 585
R395 B.n584 B.n153 585
R396 B.n586 B.n585 585
R397 B.n587 B.n152 585
R398 B.n589 B.n588 585
R399 B.n590 B.n151 585
R400 B.n592 B.n591 585
R401 B.n593 B.n150 585
R402 B.n595 B.n594 585
R403 B.n596 B.n149 585
R404 B.n598 B.n597 585
R405 B.n599 B.n148 585
R406 B.n601 B.n600 585
R407 B.n602 B.n147 585
R408 B.n604 B.n603 585
R409 B.n605 B.n146 585
R410 B.n607 B.n606 585
R411 B.n608 B.n145 585
R412 B.n610 B.n609 585
R413 B.n611 B.n144 585
R414 B.n613 B.n612 585
R415 B.n614 B.n143 585
R416 B.n616 B.n615 585
R417 B.n617 B.n142 585
R418 B.n619 B.n618 585
R419 B.n620 B.n141 585
R420 B.n622 B.n621 585
R421 B.n623 B.n140 585
R422 B.n625 B.n624 585
R423 B.n626 B.n139 585
R424 B.n628 B.n627 585
R425 B.n629 B.n138 585
R426 B.n631 B.n630 585
R427 B.n632 B.n137 585
R428 B.n634 B.n633 585
R429 B.n635 B.n136 585
R430 B.n637 B.n636 585
R431 B.n638 B.n135 585
R432 B.n640 B.n639 585
R433 B.n641 B.n134 585
R434 B.n643 B.n642 585
R435 B.n644 B.n133 585
R436 B.n646 B.n645 585
R437 B.n647 B.n132 585
R438 B.n649 B.n648 585
R439 B.n650 B.n131 585
R440 B.n652 B.n651 585
R441 B.n653 B.n130 585
R442 B.n655 B.n654 585
R443 B.n656 B.n129 585
R444 B.n658 B.n657 585
R445 B.n659 B.n128 585
R446 B.n661 B.n660 585
R447 B.n662 B.n127 585
R448 B.n664 B.n663 585
R449 B.n665 B.n126 585
R450 B.n667 B.n666 585
R451 B.n668 B.n125 585
R452 B.n670 B.n669 585
R453 B.n671 B.n124 585
R454 B.n673 B.n672 585
R455 B.n674 B.n123 585
R456 B.n676 B.n675 585
R457 B.n677 B.n122 585
R458 B.n679 B.n678 585
R459 B.n680 B.n121 585
R460 B.n682 B.n681 585
R461 B.n683 B.n120 585
R462 B.n685 B.n684 585
R463 B.n686 B.n119 585
R464 B.n688 B.n687 585
R465 B.n689 B.n118 585
R466 B.n691 B.n690 585
R467 B.n692 B.n117 585
R468 B.n694 B.n693 585
R469 B.n695 B.n116 585
R470 B.n697 B.n696 585
R471 B.n698 B.n115 585
R472 B.n700 B.n699 585
R473 B.n701 B.n114 585
R474 B.n703 B.n702 585
R475 B.n704 B.n113 585
R476 B.n706 B.n705 585
R477 B.n707 B.n112 585
R478 B.n709 B.n708 585
R479 B.n710 B.n111 585
R480 B.n712 B.n711 585
R481 B.n713 B.n110 585
R482 B.n715 B.n714 585
R483 B.n716 B.n109 585
R484 B.n718 B.n717 585
R485 B.n719 B.n108 585
R486 B.n721 B.n720 585
R487 B.n722 B.n107 585
R488 B.n724 B.n723 585
R489 B.n725 B.n106 585
R490 B.n727 B.n726 585
R491 B.n728 B.n105 585
R492 B.n730 B.n729 585
R493 B.n731 B.n104 585
R494 B.n733 B.n732 585
R495 B.n734 B.n103 585
R496 B.n736 B.n735 585
R497 B.n737 B.n102 585
R498 B.n739 B.n738 585
R499 B.n740 B.n101 585
R500 B.n742 B.n741 585
R501 B.n743 B.n100 585
R502 B.n745 B.n744 585
R503 B.n746 B.n99 585
R504 B.n748 B.n747 585
R505 B.n749 B.n98 585
R506 B.n751 B.n750 585
R507 B.n752 B.n97 585
R508 B.n754 B.n753 585
R509 B.n755 B.n96 585
R510 B.n757 B.n756 585
R511 B.n758 B.n95 585
R512 B.n760 B.n759 585
R513 B.n761 B.n94 585
R514 B.n763 B.n762 585
R515 B.n764 B.n93 585
R516 B.n766 B.n765 585
R517 B.n767 B.n92 585
R518 B.n769 B.n768 585
R519 B.n770 B.n91 585
R520 B.n903 B.n902 585
R521 B.n901 B.n44 585
R522 B.n900 B.n899 585
R523 B.n898 B.n45 585
R524 B.n897 B.n896 585
R525 B.n895 B.n46 585
R526 B.n894 B.n893 585
R527 B.n892 B.n47 585
R528 B.n891 B.n890 585
R529 B.n889 B.n48 585
R530 B.n888 B.n887 585
R531 B.n886 B.n49 585
R532 B.n885 B.n884 585
R533 B.n883 B.n50 585
R534 B.n882 B.n881 585
R535 B.n880 B.n51 585
R536 B.n879 B.n878 585
R537 B.n877 B.n52 585
R538 B.n876 B.n875 585
R539 B.n874 B.n53 585
R540 B.n873 B.n872 585
R541 B.n871 B.n54 585
R542 B.n870 B.n869 585
R543 B.n868 B.n55 585
R544 B.n867 B.n866 585
R545 B.n865 B.n56 585
R546 B.n864 B.n863 585
R547 B.n862 B.n57 585
R548 B.n861 B.n860 585
R549 B.n859 B.n58 585
R550 B.n858 B.n857 585
R551 B.n856 B.n59 585
R552 B.n855 B.n854 585
R553 B.n853 B.n60 585
R554 B.n852 B.n851 585
R555 B.n850 B.n61 585
R556 B.n849 B.n848 585
R557 B.n847 B.n62 585
R558 B.n846 B.n845 585
R559 B.n843 B.n63 585
R560 B.n842 B.n841 585
R561 B.n840 B.n66 585
R562 B.n839 B.n838 585
R563 B.n837 B.n67 585
R564 B.n836 B.n835 585
R565 B.n834 B.n68 585
R566 B.n833 B.n832 585
R567 B.n831 B.n69 585
R568 B.n829 B.n828 585
R569 B.n827 B.n72 585
R570 B.n826 B.n825 585
R571 B.n824 B.n73 585
R572 B.n823 B.n822 585
R573 B.n821 B.n74 585
R574 B.n820 B.n819 585
R575 B.n818 B.n75 585
R576 B.n817 B.n816 585
R577 B.n815 B.n76 585
R578 B.n814 B.n813 585
R579 B.n812 B.n77 585
R580 B.n811 B.n810 585
R581 B.n809 B.n78 585
R582 B.n808 B.n807 585
R583 B.n806 B.n79 585
R584 B.n805 B.n804 585
R585 B.n803 B.n80 585
R586 B.n802 B.n801 585
R587 B.n800 B.n81 585
R588 B.n799 B.n798 585
R589 B.n797 B.n82 585
R590 B.n796 B.n795 585
R591 B.n794 B.n83 585
R592 B.n793 B.n792 585
R593 B.n791 B.n84 585
R594 B.n790 B.n789 585
R595 B.n788 B.n85 585
R596 B.n787 B.n786 585
R597 B.n785 B.n86 585
R598 B.n784 B.n783 585
R599 B.n782 B.n87 585
R600 B.n781 B.n780 585
R601 B.n779 B.n88 585
R602 B.n778 B.n777 585
R603 B.n776 B.n89 585
R604 B.n775 B.n774 585
R605 B.n773 B.n90 585
R606 B.n772 B.n771 585
R607 B.n904 B.n43 585
R608 B.n906 B.n905 585
R609 B.n907 B.n42 585
R610 B.n909 B.n908 585
R611 B.n910 B.n41 585
R612 B.n912 B.n911 585
R613 B.n913 B.n40 585
R614 B.n915 B.n914 585
R615 B.n916 B.n39 585
R616 B.n918 B.n917 585
R617 B.n919 B.n38 585
R618 B.n921 B.n920 585
R619 B.n922 B.n37 585
R620 B.n924 B.n923 585
R621 B.n925 B.n36 585
R622 B.n927 B.n926 585
R623 B.n928 B.n35 585
R624 B.n930 B.n929 585
R625 B.n931 B.n34 585
R626 B.n933 B.n932 585
R627 B.n934 B.n33 585
R628 B.n936 B.n935 585
R629 B.n937 B.n32 585
R630 B.n939 B.n938 585
R631 B.n940 B.n31 585
R632 B.n942 B.n941 585
R633 B.n943 B.n30 585
R634 B.n945 B.n944 585
R635 B.n946 B.n29 585
R636 B.n948 B.n947 585
R637 B.n949 B.n28 585
R638 B.n951 B.n950 585
R639 B.n952 B.n27 585
R640 B.n954 B.n953 585
R641 B.n955 B.n26 585
R642 B.n957 B.n956 585
R643 B.n958 B.n25 585
R644 B.n960 B.n959 585
R645 B.n961 B.n24 585
R646 B.n963 B.n962 585
R647 B.n964 B.n23 585
R648 B.n966 B.n965 585
R649 B.n967 B.n22 585
R650 B.n969 B.n968 585
R651 B.n970 B.n21 585
R652 B.n972 B.n971 585
R653 B.n973 B.n20 585
R654 B.n975 B.n974 585
R655 B.n976 B.n19 585
R656 B.n978 B.n977 585
R657 B.n979 B.n18 585
R658 B.n981 B.n980 585
R659 B.n982 B.n17 585
R660 B.n984 B.n983 585
R661 B.n985 B.n16 585
R662 B.n987 B.n986 585
R663 B.n988 B.n15 585
R664 B.n990 B.n989 585
R665 B.n991 B.n14 585
R666 B.n993 B.n992 585
R667 B.n994 B.n13 585
R668 B.n996 B.n995 585
R669 B.n997 B.n12 585
R670 B.n999 B.n998 585
R671 B.n1000 B.n11 585
R672 B.n1002 B.n1001 585
R673 B.n1003 B.n10 585
R674 B.n1005 B.n1004 585
R675 B.n1006 B.n9 585
R676 B.n1008 B.n1007 585
R677 B.n1009 B.n8 585
R678 B.n1011 B.n1010 585
R679 B.n1012 B.n7 585
R680 B.n1014 B.n1013 585
R681 B.n1015 B.n6 585
R682 B.n1017 B.n1016 585
R683 B.n1018 B.n5 585
R684 B.n1020 B.n1019 585
R685 B.n1021 B.n4 585
R686 B.n1023 B.n1022 585
R687 B.n1024 B.n3 585
R688 B.n1026 B.n1025 585
R689 B.n1027 B.n0 585
R690 B.n2 B.n1 585
R691 B.n262 B.n261 585
R692 B.n264 B.n263 585
R693 B.n265 B.n260 585
R694 B.n267 B.n266 585
R695 B.n268 B.n259 585
R696 B.n270 B.n269 585
R697 B.n271 B.n258 585
R698 B.n273 B.n272 585
R699 B.n274 B.n257 585
R700 B.n276 B.n275 585
R701 B.n277 B.n256 585
R702 B.n279 B.n278 585
R703 B.n280 B.n255 585
R704 B.n282 B.n281 585
R705 B.n283 B.n254 585
R706 B.n285 B.n284 585
R707 B.n286 B.n253 585
R708 B.n288 B.n287 585
R709 B.n289 B.n252 585
R710 B.n291 B.n290 585
R711 B.n292 B.n251 585
R712 B.n294 B.n293 585
R713 B.n295 B.n250 585
R714 B.n297 B.n296 585
R715 B.n298 B.n249 585
R716 B.n300 B.n299 585
R717 B.n301 B.n248 585
R718 B.n303 B.n302 585
R719 B.n304 B.n247 585
R720 B.n306 B.n305 585
R721 B.n307 B.n246 585
R722 B.n309 B.n308 585
R723 B.n310 B.n245 585
R724 B.n312 B.n311 585
R725 B.n313 B.n244 585
R726 B.n315 B.n314 585
R727 B.n316 B.n243 585
R728 B.n318 B.n317 585
R729 B.n319 B.n242 585
R730 B.n321 B.n320 585
R731 B.n322 B.n241 585
R732 B.n324 B.n323 585
R733 B.n325 B.n240 585
R734 B.n327 B.n326 585
R735 B.n328 B.n239 585
R736 B.n330 B.n329 585
R737 B.n331 B.n238 585
R738 B.n333 B.n332 585
R739 B.n334 B.n237 585
R740 B.n336 B.n335 585
R741 B.n337 B.n236 585
R742 B.n339 B.n338 585
R743 B.n340 B.n235 585
R744 B.n342 B.n341 585
R745 B.n343 B.n234 585
R746 B.n345 B.n344 585
R747 B.n346 B.n233 585
R748 B.n348 B.n347 585
R749 B.n349 B.n232 585
R750 B.n351 B.n350 585
R751 B.n352 B.n231 585
R752 B.n354 B.n353 585
R753 B.n355 B.n230 585
R754 B.n357 B.n356 585
R755 B.n358 B.n229 585
R756 B.n360 B.n359 585
R757 B.n361 B.n228 585
R758 B.n363 B.n362 585
R759 B.n364 B.n227 585
R760 B.n366 B.n365 585
R761 B.n367 B.n226 585
R762 B.n369 B.n368 585
R763 B.n370 B.n225 585
R764 B.n372 B.n371 585
R765 B.n373 B.n224 585
R766 B.n375 B.n374 585
R767 B.n376 B.n223 585
R768 B.n378 B.n377 585
R769 B.n379 B.n222 585
R770 B.n381 B.n380 585
R771 B.n382 B.n221 585
R772 B.n384 B.n383 585
R773 B.n385 B.n384 487.695
R774 B.n520 B.n175 487.695
R775 B.n772 B.n91 487.695
R776 B.n902 B.n43 487.695
R777 B.n200 B.t6 276.204
R778 B.n456 B.t9 276.204
R779 B.n70 B.t3 276.204
R780 B.n64 B.t0 276.204
R781 B.n1029 B.n1028 256.663
R782 B.n1028 B.n1027 235.042
R783 B.n1028 B.n2 235.042
R784 B.n456 B.t10 191.544
R785 B.n70 B.t5 191.544
R786 B.n200 B.t7 191.531
R787 B.n64 B.t2 191.531
R788 B.n386 B.n385 163.367
R789 B.n386 B.n219 163.367
R790 B.n390 B.n219 163.367
R791 B.n391 B.n390 163.367
R792 B.n392 B.n391 163.367
R793 B.n392 B.n217 163.367
R794 B.n396 B.n217 163.367
R795 B.n397 B.n396 163.367
R796 B.n398 B.n397 163.367
R797 B.n398 B.n215 163.367
R798 B.n402 B.n215 163.367
R799 B.n403 B.n402 163.367
R800 B.n404 B.n403 163.367
R801 B.n404 B.n213 163.367
R802 B.n408 B.n213 163.367
R803 B.n409 B.n408 163.367
R804 B.n410 B.n409 163.367
R805 B.n410 B.n211 163.367
R806 B.n414 B.n211 163.367
R807 B.n415 B.n414 163.367
R808 B.n416 B.n415 163.367
R809 B.n416 B.n209 163.367
R810 B.n420 B.n209 163.367
R811 B.n421 B.n420 163.367
R812 B.n422 B.n421 163.367
R813 B.n422 B.n207 163.367
R814 B.n426 B.n207 163.367
R815 B.n427 B.n426 163.367
R816 B.n428 B.n427 163.367
R817 B.n428 B.n205 163.367
R818 B.n432 B.n205 163.367
R819 B.n433 B.n432 163.367
R820 B.n434 B.n433 163.367
R821 B.n434 B.n203 163.367
R822 B.n438 B.n203 163.367
R823 B.n439 B.n438 163.367
R824 B.n440 B.n439 163.367
R825 B.n440 B.n199 163.367
R826 B.n445 B.n199 163.367
R827 B.n446 B.n445 163.367
R828 B.n447 B.n446 163.367
R829 B.n447 B.n197 163.367
R830 B.n451 B.n197 163.367
R831 B.n452 B.n451 163.367
R832 B.n453 B.n452 163.367
R833 B.n453 B.n195 163.367
R834 B.n460 B.n195 163.367
R835 B.n461 B.n460 163.367
R836 B.n462 B.n461 163.367
R837 B.n462 B.n193 163.367
R838 B.n466 B.n193 163.367
R839 B.n467 B.n466 163.367
R840 B.n468 B.n467 163.367
R841 B.n468 B.n191 163.367
R842 B.n472 B.n191 163.367
R843 B.n473 B.n472 163.367
R844 B.n474 B.n473 163.367
R845 B.n474 B.n189 163.367
R846 B.n478 B.n189 163.367
R847 B.n479 B.n478 163.367
R848 B.n480 B.n479 163.367
R849 B.n480 B.n187 163.367
R850 B.n484 B.n187 163.367
R851 B.n485 B.n484 163.367
R852 B.n486 B.n485 163.367
R853 B.n486 B.n185 163.367
R854 B.n490 B.n185 163.367
R855 B.n491 B.n490 163.367
R856 B.n492 B.n491 163.367
R857 B.n492 B.n183 163.367
R858 B.n496 B.n183 163.367
R859 B.n497 B.n496 163.367
R860 B.n498 B.n497 163.367
R861 B.n498 B.n181 163.367
R862 B.n502 B.n181 163.367
R863 B.n503 B.n502 163.367
R864 B.n504 B.n503 163.367
R865 B.n504 B.n179 163.367
R866 B.n508 B.n179 163.367
R867 B.n509 B.n508 163.367
R868 B.n510 B.n509 163.367
R869 B.n510 B.n177 163.367
R870 B.n514 B.n177 163.367
R871 B.n515 B.n514 163.367
R872 B.n516 B.n515 163.367
R873 B.n516 B.n175 163.367
R874 B.n768 B.n91 163.367
R875 B.n768 B.n767 163.367
R876 B.n767 B.n766 163.367
R877 B.n766 B.n93 163.367
R878 B.n762 B.n93 163.367
R879 B.n762 B.n761 163.367
R880 B.n761 B.n760 163.367
R881 B.n760 B.n95 163.367
R882 B.n756 B.n95 163.367
R883 B.n756 B.n755 163.367
R884 B.n755 B.n754 163.367
R885 B.n754 B.n97 163.367
R886 B.n750 B.n97 163.367
R887 B.n750 B.n749 163.367
R888 B.n749 B.n748 163.367
R889 B.n748 B.n99 163.367
R890 B.n744 B.n99 163.367
R891 B.n744 B.n743 163.367
R892 B.n743 B.n742 163.367
R893 B.n742 B.n101 163.367
R894 B.n738 B.n101 163.367
R895 B.n738 B.n737 163.367
R896 B.n737 B.n736 163.367
R897 B.n736 B.n103 163.367
R898 B.n732 B.n103 163.367
R899 B.n732 B.n731 163.367
R900 B.n731 B.n730 163.367
R901 B.n730 B.n105 163.367
R902 B.n726 B.n105 163.367
R903 B.n726 B.n725 163.367
R904 B.n725 B.n724 163.367
R905 B.n724 B.n107 163.367
R906 B.n720 B.n107 163.367
R907 B.n720 B.n719 163.367
R908 B.n719 B.n718 163.367
R909 B.n718 B.n109 163.367
R910 B.n714 B.n109 163.367
R911 B.n714 B.n713 163.367
R912 B.n713 B.n712 163.367
R913 B.n712 B.n111 163.367
R914 B.n708 B.n111 163.367
R915 B.n708 B.n707 163.367
R916 B.n707 B.n706 163.367
R917 B.n706 B.n113 163.367
R918 B.n702 B.n113 163.367
R919 B.n702 B.n701 163.367
R920 B.n701 B.n700 163.367
R921 B.n700 B.n115 163.367
R922 B.n696 B.n115 163.367
R923 B.n696 B.n695 163.367
R924 B.n695 B.n694 163.367
R925 B.n694 B.n117 163.367
R926 B.n690 B.n117 163.367
R927 B.n690 B.n689 163.367
R928 B.n689 B.n688 163.367
R929 B.n688 B.n119 163.367
R930 B.n684 B.n119 163.367
R931 B.n684 B.n683 163.367
R932 B.n683 B.n682 163.367
R933 B.n682 B.n121 163.367
R934 B.n678 B.n121 163.367
R935 B.n678 B.n677 163.367
R936 B.n677 B.n676 163.367
R937 B.n676 B.n123 163.367
R938 B.n672 B.n123 163.367
R939 B.n672 B.n671 163.367
R940 B.n671 B.n670 163.367
R941 B.n670 B.n125 163.367
R942 B.n666 B.n125 163.367
R943 B.n666 B.n665 163.367
R944 B.n665 B.n664 163.367
R945 B.n664 B.n127 163.367
R946 B.n660 B.n127 163.367
R947 B.n660 B.n659 163.367
R948 B.n659 B.n658 163.367
R949 B.n658 B.n129 163.367
R950 B.n654 B.n129 163.367
R951 B.n654 B.n653 163.367
R952 B.n653 B.n652 163.367
R953 B.n652 B.n131 163.367
R954 B.n648 B.n131 163.367
R955 B.n648 B.n647 163.367
R956 B.n647 B.n646 163.367
R957 B.n646 B.n133 163.367
R958 B.n642 B.n133 163.367
R959 B.n642 B.n641 163.367
R960 B.n641 B.n640 163.367
R961 B.n640 B.n135 163.367
R962 B.n636 B.n135 163.367
R963 B.n636 B.n635 163.367
R964 B.n635 B.n634 163.367
R965 B.n634 B.n137 163.367
R966 B.n630 B.n137 163.367
R967 B.n630 B.n629 163.367
R968 B.n629 B.n628 163.367
R969 B.n628 B.n139 163.367
R970 B.n624 B.n139 163.367
R971 B.n624 B.n623 163.367
R972 B.n623 B.n622 163.367
R973 B.n622 B.n141 163.367
R974 B.n618 B.n141 163.367
R975 B.n618 B.n617 163.367
R976 B.n617 B.n616 163.367
R977 B.n616 B.n143 163.367
R978 B.n612 B.n143 163.367
R979 B.n612 B.n611 163.367
R980 B.n611 B.n610 163.367
R981 B.n610 B.n145 163.367
R982 B.n606 B.n145 163.367
R983 B.n606 B.n605 163.367
R984 B.n605 B.n604 163.367
R985 B.n604 B.n147 163.367
R986 B.n600 B.n147 163.367
R987 B.n600 B.n599 163.367
R988 B.n599 B.n598 163.367
R989 B.n598 B.n149 163.367
R990 B.n594 B.n149 163.367
R991 B.n594 B.n593 163.367
R992 B.n593 B.n592 163.367
R993 B.n592 B.n151 163.367
R994 B.n588 B.n151 163.367
R995 B.n588 B.n587 163.367
R996 B.n587 B.n586 163.367
R997 B.n586 B.n153 163.367
R998 B.n582 B.n153 163.367
R999 B.n582 B.n581 163.367
R1000 B.n581 B.n580 163.367
R1001 B.n580 B.n155 163.367
R1002 B.n576 B.n155 163.367
R1003 B.n576 B.n575 163.367
R1004 B.n575 B.n574 163.367
R1005 B.n574 B.n157 163.367
R1006 B.n570 B.n157 163.367
R1007 B.n570 B.n569 163.367
R1008 B.n569 B.n568 163.367
R1009 B.n568 B.n159 163.367
R1010 B.n564 B.n159 163.367
R1011 B.n564 B.n563 163.367
R1012 B.n563 B.n562 163.367
R1013 B.n562 B.n161 163.367
R1014 B.n558 B.n161 163.367
R1015 B.n558 B.n557 163.367
R1016 B.n557 B.n556 163.367
R1017 B.n556 B.n163 163.367
R1018 B.n552 B.n163 163.367
R1019 B.n552 B.n551 163.367
R1020 B.n551 B.n550 163.367
R1021 B.n550 B.n165 163.367
R1022 B.n546 B.n165 163.367
R1023 B.n546 B.n545 163.367
R1024 B.n545 B.n544 163.367
R1025 B.n544 B.n167 163.367
R1026 B.n540 B.n167 163.367
R1027 B.n540 B.n539 163.367
R1028 B.n539 B.n538 163.367
R1029 B.n538 B.n169 163.367
R1030 B.n534 B.n169 163.367
R1031 B.n534 B.n533 163.367
R1032 B.n533 B.n532 163.367
R1033 B.n532 B.n171 163.367
R1034 B.n528 B.n171 163.367
R1035 B.n528 B.n527 163.367
R1036 B.n527 B.n526 163.367
R1037 B.n526 B.n173 163.367
R1038 B.n522 B.n173 163.367
R1039 B.n522 B.n521 163.367
R1040 B.n521 B.n520 163.367
R1041 B.n902 B.n901 163.367
R1042 B.n901 B.n900 163.367
R1043 B.n900 B.n45 163.367
R1044 B.n896 B.n45 163.367
R1045 B.n896 B.n895 163.367
R1046 B.n895 B.n894 163.367
R1047 B.n894 B.n47 163.367
R1048 B.n890 B.n47 163.367
R1049 B.n890 B.n889 163.367
R1050 B.n889 B.n888 163.367
R1051 B.n888 B.n49 163.367
R1052 B.n884 B.n49 163.367
R1053 B.n884 B.n883 163.367
R1054 B.n883 B.n882 163.367
R1055 B.n882 B.n51 163.367
R1056 B.n878 B.n51 163.367
R1057 B.n878 B.n877 163.367
R1058 B.n877 B.n876 163.367
R1059 B.n876 B.n53 163.367
R1060 B.n872 B.n53 163.367
R1061 B.n872 B.n871 163.367
R1062 B.n871 B.n870 163.367
R1063 B.n870 B.n55 163.367
R1064 B.n866 B.n55 163.367
R1065 B.n866 B.n865 163.367
R1066 B.n865 B.n864 163.367
R1067 B.n864 B.n57 163.367
R1068 B.n860 B.n57 163.367
R1069 B.n860 B.n859 163.367
R1070 B.n859 B.n858 163.367
R1071 B.n858 B.n59 163.367
R1072 B.n854 B.n59 163.367
R1073 B.n854 B.n853 163.367
R1074 B.n853 B.n852 163.367
R1075 B.n852 B.n61 163.367
R1076 B.n848 B.n61 163.367
R1077 B.n848 B.n847 163.367
R1078 B.n847 B.n846 163.367
R1079 B.n846 B.n63 163.367
R1080 B.n841 B.n63 163.367
R1081 B.n841 B.n840 163.367
R1082 B.n840 B.n839 163.367
R1083 B.n839 B.n67 163.367
R1084 B.n835 B.n67 163.367
R1085 B.n835 B.n834 163.367
R1086 B.n834 B.n833 163.367
R1087 B.n833 B.n69 163.367
R1088 B.n828 B.n69 163.367
R1089 B.n828 B.n827 163.367
R1090 B.n827 B.n826 163.367
R1091 B.n826 B.n73 163.367
R1092 B.n822 B.n73 163.367
R1093 B.n822 B.n821 163.367
R1094 B.n821 B.n820 163.367
R1095 B.n820 B.n75 163.367
R1096 B.n816 B.n75 163.367
R1097 B.n816 B.n815 163.367
R1098 B.n815 B.n814 163.367
R1099 B.n814 B.n77 163.367
R1100 B.n810 B.n77 163.367
R1101 B.n810 B.n809 163.367
R1102 B.n809 B.n808 163.367
R1103 B.n808 B.n79 163.367
R1104 B.n804 B.n79 163.367
R1105 B.n804 B.n803 163.367
R1106 B.n803 B.n802 163.367
R1107 B.n802 B.n81 163.367
R1108 B.n798 B.n81 163.367
R1109 B.n798 B.n797 163.367
R1110 B.n797 B.n796 163.367
R1111 B.n796 B.n83 163.367
R1112 B.n792 B.n83 163.367
R1113 B.n792 B.n791 163.367
R1114 B.n791 B.n790 163.367
R1115 B.n790 B.n85 163.367
R1116 B.n786 B.n85 163.367
R1117 B.n786 B.n785 163.367
R1118 B.n785 B.n784 163.367
R1119 B.n784 B.n87 163.367
R1120 B.n780 B.n87 163.367
R1121 B.n780 B.n779 163.367
R1122 B.n779 B.n778 163.367
R1123 B.n778 B.n89 163.367
R1124 B.n774 B.n89 163.367
R1125 B.n774 B.n773 163.367
R1126 B.n773 B.n772 163.367
R1127 B.n906 B.n43 163.367
R1128 B.n907 B.n906 163.367
R1129 B.n908 B.n907 163.367
R1130 B.n908 B.n41 163.367
R1131 B.n912 B.n41 163.367
R1132 B.n913 B.n912 163.367
R1133 B.n914 B.n913 163.367
R1134 B.n914 B.n39 163.367
R1135 B.n918 B.n39 163.367
R1136 B.n919 B.n918 163.367
R1137 B.n920 B.n919 163.367
R1138 B.n920 B.n37 163.367
R1139 B.n924 B.n37 163.367
R1140 B.n925 B.n924 163.367
R1141 B.n926 B.n925 163.367
R1142 B.n926 B.n35 163.367
R1143 B.n930 B.n35 163.367
R1144 B.n931 B.n930 163.367
R1145 B.n932 B.n931 163.367
R1146 B.n932 B.n33 163.367
R1147 B.n936 B.n33 163.367
R1148 B.n937 B.n936 163.367
R1149 B.n938 B.n937 163.367
R1150 B.n938 B.n31 163.367
R1151 B.n942 B.n31 163.367
R1152 B.n943 B.n942 163.367
R1153 B.n944 B.n943 163.367
R1154 B.n944 B.n29 163.367
R1155 B.n948 B.n29 163.367
R1156 B.n949 B.n948 163.367
R1157 B.n950 B.n949 163.367
R1158 B.n950 B.n27 163.367
R1159 B.n954 B.n27 163.367
R1160 B.n955 B.n954 163.367
R1161 B.n956 B.n955 163.367
R1162 B.n956 B.n25 163.367
R1163 B.n960 B.n25 163.367
R1164 B.n961 B.n960 163.367
R1165 B.n962 B.n961 163.367
R1166 B.n962 B.n23 163.367
R1167 B.n966 B.n23 163.367
R1168 B.n967 B.n966 163.367
R1169 B.n968 B.n967 163.367
R1170 B.n968 B.n21 163.367
R1171 B.n972 B.n21 163.367
R1172 B.n973 B.n972 163.367
R1173 B.n974 B.n973 163.367
R1174 B.n974 B.n19 163.367
R1175 B.n978 B.n19 163.367
R1176 B.n979 B.n978 163.367
R1177 B.n980 B.n979 163.367
R1178 B.n980 B.n17 163.367
R1179 B.n984 B.n17 163.367
R1180 B.n985 B.n984 163.367
R1181 B.n986 B.n985 163.367
R1182 B.n986 B.n15 163.367
R1183 B.n990 B.n15 163.367
R1184 B.n991 B.n990 163.367
R1185 B.n992 B.n991 163.367
R1186 B.n992 B.n13 163.367
R1187 B.n996 B.n13 163.367
R1188 B.n997 B.n996 163.367
R1189 B.n998 B.n997 163.367
R1190 B.n998 B.n11 163.367
R1191 B.n1002 B.n11 163.367
R1192 B.n1003 B.n1002 163.367
R1193 B.n1004 B.n1003 163.367
R1194 B.n1004 B.n9 163.367
R1195 B.n1008 B.n9 163.367
R1196 B.n1009 B.n1008 163.367
R1197 B.n1010 B.n1009 163.367
R1198 B.n1010 B.n7 163.367
R1199 B.n1014 B.n7 163.367
R1200 B.n1015 B.n1014 163.367
R1201 B.n1016 B.n1015 163.367
R1202 B.n1016 B.n5 163.367
R1203 B.n1020 B.n5 163.367
R1204 B.n1021 B.n1020 163.367
R1205 B.n1022 B.n1021 163.367
R1206 B.n1022 B.n3 163.367
R1207 B.n1026 B.n3 163.367
R1208 B.n1027 B.n1026 163.367
R1209 B.n261 B.n2 163.367
R1210 B.n264 B.n261 163.367
R1211 B.n265 B.n264 163.367
R1212 B.n266 B.n265 163.367
R1213 B.n266 B.n259 163.367
R1214 B.n270 B.n259 163.367
R1215 B.n271 B.n270 163.367
R1216 B.n272 B.n271 163.367
R1217 B.n272 B.n257 163.367
R1218 B.n276 B.n257 163.367
R1219 B.n277 B.n276 163.367
R1220 B.n278 B.n277 163.367
R1221 B.n278 B.n255 163.367
R1222 B.n282 B.n255 163.367
R1223 B.n283 B.n282 163.367
R1224 B.n284 B.n283 163.367
R1225 B.n284 B.n253 163.367
R1226 B.n288 B.n253 163.367
R1227 B.n289 B.n288 163.367
R1228 B.n290 B.n289 163.367
R1229 B.n290 B.n251 163.367
R1230 B.n294 B.n251 163.367
R1231 B.n295 B.n294 163.367
R1232 B.n296 B.n295 163.367
R1233 B.n296 B.n249 163.367
R1234 B.n300 B.n249 163.367
R1235 B.n301 B.n300 163.367
R1236 B.n302 B.n301 163.367
R1237 B.n302 B.n247 163.367
R1238 B.n306 B.n247 163.367
R1239 B.n307 B.n306 163.367
R1240 B.n308 B.n307 163.367
R1241 B.n308 B.n245 163.367
R1242 B.n312 B.n245 163.367
R1243 B.n313 B.n312 163.367
R1244 B.n314 B.n313 163.367
R1245 B.n314 B.n243 163.367
R1246 B.n318 B.n243 163.367
R1247 B.n319 B.n318 163.367
R1248 B.n320 B.n319 163.367
R1249 B.n320 B.n241 163.367
R1250 B.n324 B.n241 163.367
R1251 B.n325 B.n324 163.367
R1252 B.n326 B.n325 163.367
R1253 B.n326 B.n239 163.367
R1254 B.n330 B.n239 163.367
R1255 B.n331 B.n330 163.367
R1256 B.n332 B.n331 163.367
R1257 B.n332 B.n237 163.367
R1258 B.n336 B.n237 163.367
R1259 B.n337 B.n336 163.367
R1260 B.n338 B.n337 163.367
R1261 B.n338 B.n235 163.367
R1262 B.n342 B.n235 163.367
R1263 B.n343 B.n342 163.367
R1264 B.n344 B.n343 163.367
R1265 B.n344 B.n233 163.367
R1266 B.n348 B.n233 163.367
R1267 B.n349 B.n348 163.367
R1268 B.n350 B.n349 163.367
R1269 B.n350 B.n231 163.367
R1270 B.n354 B.n231 163.367
R1271 B.n355 B.n354 163.367
R1272 B.n356 B.n355 163.367
R1273 B.n356 B.n229 163.367
R1274 B.n360 B.n229 163.367
R1275 B.n361 B.n360 163.367
R1276 B.n362 B.n361 163.367
R1277 B.n362 B.n227 163.367
R1278 B.n366 B.n227 163.367
R1279 B.n367 B.n366 163.367
R1280 B.n368 B.n367 163.367
R1281 B.n368 B.n225 163.367
R1282 B.n372 B.n225 163.367
R1283 B.n373 B.n372 163.367
R1284 B.n374 B.n373 163.367
R1285 B.n374 B.n223 163.367
R1286 B.n378 B.n223 163.367
R1287 B.n379 B.n378 163.367
R1288 B.n380 B.n379 163.367
R1289 B.n380 B.n221 163.367
R1290 B.n384 B.n221 163.367
R1291 B.n457 B.t11 108.538
R1292 B.n71 B.t4 108.538
R1293 B.n201 B.t8 108.525
R1294 B.n65 B.t1 108.525
R1295 B.n201 B.n200 83.0066
R1296 B.n457 B.n456 83.0066
R1297 B.n71 B.n70 83.0066
R1298 B.n65 B.n64 83.0066
R1299 B.n443 B.n201 59.5399
R1300 B.n458 B.n457 59.5399
R1301 B.n830 B.n71 59.5399
R1302 B.n844 B.n65 59.5399
R1303 B.n904 B.n903 31.6883
R1304 B.n771 B.n770 31.6883
R1305 B.n519 B.n518 31.6883
R1306 B.n383 B.n220 31.6883
R1307 B B.n1029 18.0485
R1308 B.n905 B.n904 10.6151
R1309 B.n905 B.n42 10.6151
R1310 B.n909 B.n42 10.6151
R1311 B.n910 B.n909 10.6151
R1312 B.n911 B.n910 10.6151
R1313 B.n911 B.n40 10.6151
R1314 B.n915 B.n40 10.6151
R1315 B.n916 B.n915 10.6151
R1316 B.n917 B.n916 10.6151
R1317 B.n917 B.n38 10.6151
R1318 B.n921 B.n38 10.6151
R1319 B.n922 B.n921 10.6151
R1320 B.n923 B.n922 10.6151
R1321 B.n923 B.n36 10.6151
R1322 B.n927 B.n36 10.6151
R1323 B.n928 B.n927 10.6151
R1324 B.n929 B.n928 10.6151
R1325 B.n929 B.n34 10.6151
R1326 B.n933 B.n34 10.6151
R1327 B.n934 B.n933 10.6151
R1328 B.n935 B.n934 10.6151
R1329 B.n935 B.n32 10.6151
R1330 B.n939 B.n32 10.6151
R1331 B.n940 B.n939 10.6151
R1332 B.n941 B.n940 10.6151
R1333 B.n941 B.n30 10.6151
R1334 B.n945 B.n30 10.6151
R1335 B.n946 B.n945 10.6151
R1336 B.n947 B.n946 10.6151
R1337 B.n947 B.n28 10.6151
R1338 B.n951 B.n28 10.6151
R1339 B.n952 B.n951 10.6151
R1340 B.n953 B.n952 10.6151
R1341 B.n953 B.n26 10.6151
R1342 B.n957 B.n26 10.6151
R1343 B.n958 B.n957 10.6151
R1344 B.n959 B.n958 10.6151
R1345 B.n959 B.n24 10.6151
R1346 B.n963 B.n24 10.6151
R1347 B.n964 B.n963 10.6151
R1348 B.n965 B.n964 10.6151
R1349 B.n965 B.n22 10.6151
R1350 B.n969 B.n22 10.6151
R1351 B.n970 B.n969 10.6151
R1352 B.n971 B.n970 10.6151
R1353 B.n971 B.n20 10.6151
R1354 B.n975 B.n20 10.6151
R1355 B.n976 B.n975 10.6151
R1356 B.n977 B.n976 10.6151
R1357 B.n977 B.n18 10.6151
R1358 B.n981 B.n18 10.6151
R1359 B.n982 B.n981 10.6151
R1360 B.n983 B.n982 10.6151
R1361 B.n983 B.n16 10.6151
R1362 B.n987 B.n16 10.6151
R1363 B.n988 B.n987 10.6151
R1364 B.n989 B.n988 10.6151
R1365 B.n989 B.n14 10.6151
R1366 B.n993 B.n14 10.6151
R1367 B.n994 B.n993 10.6151
R1368 B.n995 B.n994 10.6151
R1369 B.n995 B.n12 10.6151
R1370 B.n999 B.n12 10.6151
R1371 B.n1000 B.n999 10.6151
R1372 B.n1001 B.n1000 10.6151
R1373 B.n1001 B.n10 10.6151
R1374 B.n1005 B.n10 10.6151
R1375 B.n1006 B.n1005 10.6151
R1376 B.n1007 B.n1006 10.6151
R1377 B.n1007 B.n8 10.6151
R1378 B.n1011 B.n8 10.6151
R1379 B.n1012 B.n1011 10.6151
R1380 B.n1013 B.n1012 10.6151
R1381 B.n1013 B.n6 10.6151
R1382 B.n1017 B.n6 10.6151
R1383 B.n1018 B.n1017 10.6151
R1384 B.n1019 B.n1018 10.6151
R1385 B.n1019 B.n4 10.6151
R1386 B.n1023 B.n4 10.6151
R1387 B.n1024 B.n1023 10.6151
R1388 B.n1025 B.n1024 10.6151
R1389 B.n1025 B.n0 10.6151
R1390 B.n903 B.n44 10.6151
R1391 B.n899 B.n44 10.6151
R1392 B.n899 B.n898 10.6151
R1393 B.n898 B.n897 10.6151
R1394 B.n897 B.n46 10.6151
R1395 B.n893 B.n46 10.6151
R1396 B.n893 B.n892 10.6151
R1397 B.n892 B.n891 10.6151
R1398 B.n891 B.n48 10.6151
R1399 B.n887 B.n48 10.6151
R1400 B.n887 B.n886 10.6151
R1401 B.n886 B.n885 10.6151
R1402 B.n885 B.n50 10.6151
R1403 B.n881 B.n50 10.6151
R1404 B.n881 B.n880 10.6151
R1405 B.n880 B.n879 10.6151
R1406 B.n879 B.n52 10.6151
R1407 B.n875 B.n52 10.6151
R1408 B.n875 B.n874 10.6151
R1409 B.n874 B.n873 10.6151
R1410 B.n873 B.n54 10.6151
R1411 B.n869 B.n54 10.6151
R1412 B.n869 B.n868 10.6151
R1413 B.n868 B.n867 10.6151
R1414 B.n867 B.n56 10.6151
R1415 B.n863 B.n56 10.6151
R1416 B.n863 B.n862 10.6151
R1417 B.n862 B.n861 10.6151
R1418 B.n861 B.n58 10.6151
R1419 B.n857 B.n58 10.6151
R1420 B.n857 B.n856 10.6151
R1421 B.n856 B.n855 10.6151
R1422 B.n855 B.n60 10.6151
R1423 B.n851 B.n60 10.6151
R1424 B.n851 B.n850 10.6151
R1425 B.n850 B.n849 10.6151
R1426 B.n849 B.n62 10.6151
R1427 B.n845 B.n62 10.6151
R1428 B.n843 B.n842 10.6151
R1429 B.n842 B.n66 10.6151
R1430 B.n838 B.n66 10.6151
R1431 B.n838 B.n837 10.6151
R1432 B.n837 B.n836 10.6151
R1433 B.n836 B.n68 10.6151
R1434 B.n832 B.n68 10.6151
R1435 B.n832 B.n831 10.6151
R1436 B.n829 B.n72 10.6151
R1437 B.n825 B.n72 10.6151
R1438 B.n825 B.n824 10.6151
R1439 B.n824 B.n823 10.6151
R1440 B.n823 B.n74 10.6151
R1441 B.n819 B.n74 10.6151
R1442 B.n819 B.n818 10.6151
R1443 B.n818 B.n817 10.6151
R1444 B.n817 B.n76 10.6151
R1445 B.n813 B.n76 10.6151
R1446 B.n813 B.n812 10.6151
R1447 B.n812 B.n811 10.6151
R1448 B.n811 B.n78 10.6151
R1449 B.n807 B.n78 10.6151
R1450 B.n807 B.n806 10.6151
R1451 B.n806 B.n805 10.6151
R1452 B.n805 B.n80 10.6151
R1453 B.n801 B.n80 10.6151
R1454 B.n801 B.n800 10.6151
R1455 B.n800 B.n799 10.6151
R1456 B.n799 B.n82 10.6151
R1457 B.n795 B.n82 10.6151
R1458 B.n795 B.n794 10.6151
R1459 B.n794 B.n793 10.6151
R1460 B.n793 B.n84 10.6151
R1461 B.n789 B.n84 10.6151
R1462 B.n789 B.n788 10.6151
R1463 B.n788 B.n787 10.6151
R1464 B.n787 B.n86 10.6151
R1465 B.n783 B.n86 10.6151
R1466 B.n783 B.n782 10.6151
R1467 B.n782 B.n781 10.6151
R1468 B.n781 B.n88 10.6151
R1469 B.n777 B.n88 10.6151
R1470 B.n777 B.n776 10.6151
R1471 B.n776 B.n775 10.6151
R1472 B.n775 B.n90 10.6151
R1473 B.n771 B.n90 10.6151
R1474 B.n770 B.n769 10.6151
R1475 B.n769 B.n92 10.6151
R1476 B.n765 B.n92 10.6151
R1477 B.n765 B.n764 10.6151
R1478 B.n764 B.n763 10.6151
R1479 B.n763 B.n94 10.6151
R1480 B.n759 B.n94 10.6151
R1481 B.n759 B.n758 10.6151
R1482 B.n758 B.n757 10.6151
R1483 B.n757 B.n96 10.6151
R1484 B.n753 B.n96 10.6151
R1485 B.n753 B.n752 10.6151
R1486 B.n752 B.n751 10.6151
R1487 B.n751 B.n98 10.6151
R1488 B.n747 B.n98 10.6151
R1489 B.n747 B.n746 10.6151
R1490 B.n746 B.n745 10.6151
R1491 B.n745 B.n100 10.6151
R1492 B.n741 B.n100 10.6151
R1493 B.n741 B.n740 10.6151
R1494 B.n740 B.n739 10.6151
R1495 B.n739 B.n102 10.6151
R1496 B.n735 B.n102 10.6151
R1497 B.n735 B.n734 10.6151
R1498 B.n734 B.n733 10.6151
R1499 B.n733 B.n104 10.6151
R1500 B.n729 B.n104 10.6151
R1501 B.n729 B.n728 10.6151
R1502 B.n728 B.n727 10.6151
R1503 B.n727 B.n106 10.6151
R1504 B.n723 B.n106 10.6151
R1505 B.n723 B.n722 10.6151
R1506 B.n722 B.n721 10.6151
R1507 B.n721 B.n108 10.6151
R1508 B.n717 B.n108 10.6151
R1509 B.n717 B.n716 10.6151
R1510 B.n716 B.n715 10.6151
R1511 B.n715 B.n110 10.6151
R1512 B.n711 B.n110 10.6151
R1513 B.n711 B.n710 10.6151
R1514 B.n710 B.n709 10.6151
R1515 B.n709 B.n112 10.6151
R1516 B.n705 B.n112 10.6151
R1517 B.n705 B.n704 10.6151
R1518 B.n704 B.n703 10.6151
R1519 B.n703 B.n114 10.6151
R1520 B.n699 B.n114 10.6151
R1521 B.n699 B.n698 10.6151
R1522 B.n698 B.n697 10.6151
R1523 B.n697 B.n116 10.6151
R1524 B.n693 B.n116 10.6151
R1525 B.n693 B.n692 10.6151
R1526 B.n692 B.n691 10.6151
R1527 B.n691 B.n118 10.6151
R1528 B.n687 B.n118 10.6151
R1529 B.n687 B.n686 10.6151
R1530 B.n686 B.n685 10.6151
R1531 B.n685 B.n120 10.6151
R1532 B.n681 B.n120 10.6151
R1533 B.n681 B.n680 10.6151
R1534 B.n680 B.n679 10.6151
R1535 B.n679 B.n122 10.6151
R1536 B.n675 B.n122 10.6151
R1537 B.n675 B.n674 10.6151
R1538 B.n674 B.n673 10.6151
R1539 B.n673 B.n124 10.6151
R1540 B.n669 B.n124 10.6151
R1541 B.n669 B.n668 10.6151
R1542 B.n668 B.n667 10.6151
R1543 B.n667 B.n126 10.6151
R1544 B.n663 B.n126 10.6151
R1545 B.n663 B.n662 10.6151
R1546 B.n662 B.n661 10.6151
R1547 B.n661 B.n128 10.6151
R1548 B.n657 B.n128 10.6151
R1549 B.n657 B.n656 10.6151
R1550 B.n656 B.n655 10.6151
R1551 B.n655 B.n130 10.6151
R1552 B.n651 B.n130 10.6151
R1553 B.n651 B.n650 10.6151
R1554 B.n650 B.n649 10.6151
R1555 B.n649 B.n132 10.6151
R1556 B.n645 B.n132 10.6151
R1557 B.n645 B.n644 10.6151
R1558 B.n644 B.n643 10.6151
R1559 B.n643 B.n134 10.6151
R1560 B.n639 B.n134 10.6151
R1561 B.n639 B.n638 10.6151
R1562 B.n638 B.n637 10.6151
R1563 B.n637 B.n136 10.6151
R1564 B.n633 B.n136 10.6151
R1565 B.n633 B.n632 10.6151
R1566 B.n632 B.n631 10.6151
R1567 B.n631 B.n138 10.6151
R1568 B.n627 B.n138 10.6151
R1569 B.n627 B.n626 10.6151
R1570 B.n626 B.n625 10.6151
R1571 B.n625 B.n140 10.6151
R1572 B.n621 B.n140 10.6151
R1573 B.n621 B.n620 10.6151
R1574 B.n620 B.n619 10.6151
R1575 B.n619 B.n142 10.6151
R1576 B.n615 B.n142 10.6151
R1577 B.n615 B.n614 10.6151
R1578 B.n614 B.n613 10.6151
R1579 B.n613 B.n144 10.6151
R1580 B.n609 B.n144 10.6151
R1581 B.n609 B.n608 10.6151
R1582 B.n608 B.n607 10.6151
R1583 B.n607 B.n146 10.6151
R1584 B.n603 B.n146 10.6151
R1585 B.n603 B.n602 10.6151
R1586 B.n602 B.n601 10.6151
R1587 B.n601 B.n148 10.6151
R1588 B.n597 B.n148 10.6151
R1589 B.n597 B.n596 10.6151
R1590 B.n596 B.n595 10.6151
R1591 B.n595 B.n150 10.6151
R1592 B.n591 B.n150 10.6151
R1593 B.n591 B.n590 10.6151
R1594 B.n590 B.n589 10.6151
R1595 B.n589 B.n152 10.6151
R1596 B.n585 B.n152 10.6151
R1597 B.n585 B.n584 10.6151
R1598 B.n584 B.n583 10.6151
R1599 B.n583 B.n154 10.6151
R1600 B.n579 B.n154 10.6151
R1601 B.n579 B.n578 10.6151
R1602 B.n578 B.n577 10.6151
R1603 B.n577 B.n156 10.6151
R1604 B.n573 B.n156 10.6151
R1605 B.n573 B.n572 10.6151
R1606 B.n572 B.n571 10.6151
R1607 B.n571 B.n158 10.6151
R1608 B.n567 B.n158 10.6151
R1609 B.n567 B.n566 10.6151
R1610 B.n566 B.n565 10.6151
R1611 B.n565 B.n160 10.6151
R1612 B.n561 B.n160 10.6151
R1613 B.n561 B.n560 10.6151
R1614 B.n560 B.n559 10.6151
R1615 B.n559 B.n162 10.6151
R1616 B.n555 B.n162 10.6151
R1617 B.n555 B.n554 10.6151
R1618 B.n554 B.n553 10.6151
R1619 B.n553 B.n164 10.6151
R1620 B.n549 B.n164 10.6151
R1621 B.n549 B.n548 10.6151
R1622 B.n548 B.n547 10.6151
R1623 B.n547 B.n166 10.6151
R1624 B.n543 B.n166 10.6151
R1625 B.n543 B.n542 10.6151
R1626 B.n542 B.n541 10.6151
R1627 B.n541 B.n168 10.6151
R1628 B.n537 B.n168 10.6151
R1629 B.n537 B.n536 10.6151
R1630 B.n536 B.n535 10.6151
R1631 B.n535 B.n170 10.6151
R1632 B.n531 B.n170 10.6151
R1633 B.n531 B.n530 10.6151
R1634 B.n530 B.n529 10.6151
R1635 B.n529 B.n172 10.6151
R1636 B.n525 B.n172 10.6151
R1637 B.n525 B.n524 10.6151
R1638 B.n524 B.n523 10.6151
R1639 B.n523 B.n174 10.6151
R1640 B.n519 B.n174 10.6151
R1641 B.n262 B.n1 10.6151
R1642 B.n263 B.n262 10.6151
R1643 B.n263 B.n260 10.6151
R1644 B.n267 B.n260 10.6151
R1645 B.n268 B.n267 10.6151
R1646 B.n269 B.n268 10.6151
R1647 B.n269 B.n258 10.6151
R1648 B.n273 B.n258 10.6151
R1649 B.n274 B.n273 10.6151
R1650 B.n275 B.n274 10.6151
R1651 B.n275 B.n256 10.6151
R1652 B.n279 B.n256 10.6151
R1653 B.n280 B.n279 10.6151
R1654 B.n281 B.n280 10.6151
R1655 B.n281 B.n254 10.6151
R1656 B.n285 B.n254 10.6151
R1657 B.n286 B.n285 10.6151
R1658 B.n287 B.n286 10.6151
R1659 B.n287 B.n252 10.6151
R1660 B.n291 B.n252 10.6151
R1661 B.n292 B.n291 10.6151
R1662 B.n293 B.n292 10.6151
R1663 B.n293 B.n250 10.6151
R1664 B.n297 B.n250 10.6151
R1665 B.n298 B.n297 10.6151
R1666 B.n299 B.n298 10.6151
R1667 B.n299 B.n248 10.6151
R1668 B.n303 B.n248 10.6151
R1669 B.n304 B.n303 10.6151
R1670 B.n305 B.n304 10.6151
R1671 B.n305 B.n246 10.6151
R1672 B.n309 B.n246 10.6151
R1673 B.n310 B.n309 10.6151
R1674 B.n311 B.n310 10.6151
R1675 B.n311 B.n244 10.6151
R1676 B.n315 B.n244 10.6151
R1677 B.n316 B.n315 10.6151
R1678 B.n317 B.n316 10.6151
R1679 B.n317 B.n242 10.6151
R1680 B.n321 B.n242 10.6151
R1681 B.n322 B.n321 10.6151
R1682 B.n323 B.n322 10.6151
R1683 B.n323 B.n240 10.6151
R1684 B.n327 B.n240 10.6151
R1685 B.n328 B.n327 10.6151
R1686 B.n329 B.n328 10.6151
R1687 B.n329 B.n238 10.6151
R1688 B.n333 B.n238 10.6151
R1689 B.n334 B.n333 10.6151
R1690 B.n335 B.n334 10.6151
R1691 B.n335 B.n236 10.6151
R1692 B.n339 B.n236 10.6151
R1693 B.n340 B.n339 10.6151
R1694 B.n341 B.n340 10.6151
R1695 B.n341 B.n234 10.6151
R1696 B.n345 B.n234 10.6151
R1697 B.n346 B.n345 10.6151
R1698 B.n347 B.n346 10.6151
R1699 B.n347 B.n232 10.6151
R1700 B.n351 B.n232 10.6151
R1701 B.n352 B.n351 10.6151
R1702 B.n353 B.n352 10.6151
R1703 B.n353 B.n230 10.6151
R1704 B.n357 B.n230 10.6151
R1705 B.n358 B.n357 10.6151
R1706 B.n359 B.n358 10.6151
R1707 B.n359 B.n228 10.6151
R1708 B.n363 B.n228 10.6151
R1709 B.n364 B.n363 10.6151
R1710 B.n365 B.n364 10.6151
R1711 B.n365 B.n226 10.6151
R1712 B.n369 B.n226 10.6151
R1713 B.n370 B.n369 10.6151
R1714 B.n371 B.n370 10.6151
R1715 B.n371 B.n224 10.6151
R1716 B.n375 B.n224 10.6151
R1717 B.n376 B.n375 10.6151
R1718 B.n377 B.n376 10.6151
R1719 B.n377 B.n222 10.6151
R1720 B.n381 B.n222 10.6151
R1721 B.n382 B.n381 10.6151
R1722 B.n383 B.n382 10.6151
R1723 B.n387 B.n220 10.6151
R1724 B.n388 B.n387 10.6151
R1725 B.n389 B.n388 10.6151
R1726 B.n389 B.n218 10.6151
R1727 B.n393 B.n218 10.6151
R1728 B.n394 B.n393 10.6151
R1729 B.n395 B.n394 10.6151
R1730 B.n395 B.n216 10.6151
R1731 B.n399 B.n216 10.6151
R1732 B.n400 B.n399 10.6151
R1733 B.n401 B.n400 10.6151
R1734 B.n401 B.n214 10.6151
R1735 B.n405 B.n214 10.6151
R1736 B.n406 B.n405 10.6151
R1737 B.n407 B.n406 10.6151
R1738 B.n407 B.n212 10.6151
R1739 B.n411 B.n212 10.6151
R1740 B.n412 B.n411 10.6151
R1741 B.n413 B.n412 10.6151
R1742 B.n413 B.n210 10.6151
R1743 B.n417 B.n210 10.6151
R1744 B.n418 B.n417 10.6151
R1745 B.n419 B.n418 10.6151
R1746 B.n419 B.n208 10.6151
R1747 B.n423 B.n208 10.6151
R1748 B.n424 B.n423 10.6151
R1749 B.n425 B.n424 10.6151
R1750 B.n425 B.n206 10.6151
R1751 B.n429 B.n206 10.6151
R1752 B.n430 B.n429 10.6151
R1753 B.n431 B.n430 10.6151
R1754 B.n431 B.n204 10.6151
R1755 B.n435 B.n204 10.6151
R1756 B.n436 B.n435 10.6151
R1757 B.n437 B.n436 10.6151
R1758 B.n437 B.n202 10.6151
R1759 B.n441 B.n202 10.6151
R1760 B.n442 B.n441 10.6151
R1761 B.n444 B.n198 10.6151
R1762 B.n448 B.n198 10.6151
R1763 B.n449 B.n448 10.6151
R1764 B.n450 B.n449 10.6151
R1765 B.n450 B.n196 10.6151
R1766 B.n454 B.n196 10.6151
R1767 B.n455 B.n454 10.6151
R1768 B.n459 B.n455 10.6151
R1769 B.n463 B.n194 10.6151
R1770 B.n464 B.n463 10.6151
R1771 B.n465 B.n464 10.6151
R1772 B.n465 B.n192 10.6151
R1773 B.n469 B.n192 10.6151
R1774 B.n470 B.n469 10.6151
R1775 B.n471 B.n470 10.6151
R1776 B.n471 B.n190 10.6151
R1777 B.n475 B.n190 10.6151
R1778 B.n476 B.n475 10.6151
R1779 B.n477 B.n476 10.6151
R1780 B.n477 B.n188 10.6151
R1781 B.n481 B.n188 10.6151
R1782 B.n482 B.n481 10.6151
R1783 B.n483 B.n482 10.6151
R1784 B.n483 B.n186 10.6151
R1785 B.n487 B.n186 10.6151
R1786 B.n488 B.n487 10.6151
R1787 B.n489 B.n488 10.6151
R1788 B.n489 B.n184 10.6151
R1789 B.n493 B.n184 10.6151
R1790 B.n494 B.n493 10.6151
R1791 B.n495 B.n494 10.6151
R1792 B.n495 B.n182 10.6151
R1793 B.n499 B.n182 10.6151
R1794 B.n500 B.n499 10.6151
R1795 B.n501 B.n500 10.6151
R1796 B.n501 B.n180 10.6151
R1797 B.n505 B.n180 10.6151
R1798 B.n506 B.n505 10.6151
R1799 B.n507 B.n506 10.6151
R1800 B.n507 B.n178 10.6151
R1801 B.n511 B.n178 10.6151
R1802 B.n512 B.n511 10.6151
R1803 B.n513 B.n512 10.6151
R1804 B.n513 B.n176 10.6151
R1805 B.n517 B.n176 10.6151
R1806 B.n518 B.n517 10.6151
R1807 B.n1029 B.n0 8.11757
R1808 B.n1029 B.n1 8.11757
R1809 B.n844 B.n843 6.5566
R1810 B.n831 B.n830 6.5566
R1811 B.n444 B.n443 6.5566
R1812 B.n459 B.n458 6.5566
R1813 B.n845 B.n844 4.05904
R1814 B.n830 B.n829 4.05904
R1815 B.n443 B.n442 4.05904
R1816 B.n458 B.n194 4.05904
R1817 VN.n112 VN.n111 161.3
R1818 VN.n110 VN.n58 161.3
R1819 VN.n109 VN.n108 161.3
R1820 VN.n107 VN.n59 161.3
R1821 VN.n106 VN.n105 161.3
R1822 VN.n104 VN.n60 161.3
R1823 VN.n103 VN.n102 161.3
R1824 VN.n101 VN.n61 161.3
R1825 VN.n100 VN.n99 161.3
R1826 VN.n97 VN.n62 161.3
R1827 VN.n96 VN.n95 161.3
R1828 VN.n94 VN.n63 161.3
R1829 VN.n93 VN.n92 161.3
R1830 VN.n91 VN.n64 161.3
R1831 VN.n90 VN.n89 161.3
R1832 VN.n88 VN.n65 161.3
R1833 VN.n87 VN.n86 161.3
R1834 VN.n85 VN.n66 161.3
R1835 VN.n84 VN.n83 161.3
R1836 VN.n82 VN.n67 161.3
R1837 VN.n81 VN.n80 161.3
R1838 VN.n79 VN.n68 161.3
R1839 VN.n78 VN.n77 161.3
R1840 VN.n76 VN.n69 161.3
R1841 VN.n75 VN.n74 161.3
R1842 VN.n73 VN.n70 161.3
R1843 VN.n55 VN.n54 161.3
R1844 VN.n53 VN.n1 161.3
R1845 VN.n52 VN.n51 161.3
R1846 VN.n50 VN.n2 161.3
R1847 VN.n49 VN.n48 161.3
R1848 VN.n47 VN.n3 161.3
R1849 VN.n46 VN.n45 161.3
R1850 VN.n44 VN.n4 161.3
R1851 VN.n43 VN.n42 161.3
R1852 VN.n40 VN.n5 161.3
R1853 VN.n39 VN.n38 161.3
R1854 VN.n37 VN.n6 161.3
R1855 VN.n36 VN.n35 161.3
R1856 VN.n34 VN.n7 161.3
R1857 VN.n33 VN.n32 161.3
R1858 VN.n31 VN.n8 161.3
R1859 VN.n30 VN.n29 161.3
R1860 VN.n28 VN.n9 161.3
R1861 VN.n27 VN.n26 161.3
R1862 VN.n25 VN.n10 161.3
R1863 VN.n24 VN.n23 161.3
R1864 VN.n22 VN.n11 161.3
R1865 VN.n21 VN.n20 161.3
R1866 VN.n19 VN.n12 161.3
R1867 VN.n18 VN.n17 161.3
R1868 VN.n16 VN.n13 161.3
R1869 VN.n71 VN.t3 99.6589
R1870 VN.n14 VN.t6 99.6589
R1871 VN.n56 VN.n0 87.2945
R1872 VN.n113 VN.n57 87.2945
R1873 VN.n28 VN.t1 66.7483
R1874 VN.n15 VN.t9 66.7483
R1875 VN.n41 VN.t2 66.7483
R1876 VN.n0 VN.t5 66.7483
R1877 VN.n85 VN.t4 66.7483
R1878 VN.n72 VN.t7 66.7483
R1879 VN.n98 VN.t8 66.7483
R1880 VN.n57 VN.t0 66.7483
R1881 VN.n15 VN.n14 61.6104
R1882 VN.n72 VN.n71 61.6104
R1883 VN VN.n113 59.9072
R1884 VN.n22 VN.n21 54.1398
R1885 VN.n35 VN.n34 54.1398
R1886 VN.n79 VN.n78 54.1398
R1887 VN.n92 VN.n91 54.1398
R1888 VN.n48 VN.n47 48.3272
R1889 VN.n105 VN.n104 48.3272
R1890 VN.n48 VN.n2 32.8269
R1891 VN.n105 VN.n59 32.8269
R1892 VN.n23 VN.n22 27.0143
R1893 VN.n34 VN.n33 27.0143
R1894 VN.n80 VN.n79 27.0143
R1895 VN.n91 VN.n90 27.0143
R1896 VN.n17 VN.n16 24.5923
R1897 VN.n17 VN.n12 24.5923
R1898 VN.n21 VN.n12 24.5923
R1899 VN.n23 VN.n10 24.5923
R1900 VN.n27 VN.n10 24.5923
R1901 VN.n28 VN.n27 24.5923
R1902 VN.n29 VN.n28 24.5923
R1903 VN.n29 VN.n8 24.5923
R1904 VN.n33 VN.n8 24.5923
R1905 VN.n35 VN.n6 24.5923
R1906 VN.n39 VN.n6 24.5923
R1907 VN.n40 VN.n39 24.5923
R1908 VN.n42 VN.n4 24.5923
R1909 VN.n46 VN.n4 24.5923
R1910 VN.n47 VN.n46 24.5923
R1911 VN.n52 VN.n2 24.5923
R1912 VN.n53 VN.n52 24.5923
R1913 VN.n54 VN.n53 24.5923
R1914 VN.n78 VN.n69 24.5923
R1915 VN.n74 VN.n69 24.5923
R1916 VN.n74 VN.n73 24.5923
R1917 VN.n90 VN.n65 24.5923
R1918 VN.n86 VN.n65 24.5923
R1919 VN.n86 VN.n85 24.5923
R1920 VN.n85 VN.n84 24.5923
R1921 VN.n84 VN.n67 24.5923
R1922 VN.n80 VN.n67 24.5923
R1923 VN.n104 VN.n103 24.5923
R1924 VN.n103 VN.n61 24.5923
R1925 VN.n99 VN.n61 24.5923
R1926 VN.n97 VN.n96 24.5923
R1927 VN.n96 VN.n63 24.5923
R1928 VN.n92 VN.n63 24.5923
R1929 VN.n111 VN.n110 24.5923
R1930 VN.n110 VN.n109 24.5923
R1931 VN.n109 VN.n59 24.5923
R1932 VN.n16 VN.n15 13.7719
R1933 VN.n41 VN.n40 13.7719
R1934 VN.n73 VN.n72 13.7719
R1935 VN.n98 VN.n97 13.7719
R1936 VN.n42 VN.n41 10.8209
R1937 VN.n99 VN.n98 10.8209
R1938 VN.n54 VN.n0 2.95152
R1939 VN.n111 VN.n57 2.95152
R1940 VN.n71 VN.n70 2.45425
R1941 VN.n14 VN.n13 2.45425
R1942 VN.n113 VN.n112 0.354861
R1943 VN.n56 VN.n55 0.354861
R1944 VN VN.n56 0.267071
R1945 VN.n112 VN.n58 0.189894
R1946 VN.n108 VN.n58 0.189894
R1947 VN.n108 VN.n107 0.189894
R1948 VN.n107 VN.n106 0.189894
R1949 VN.n106 VN.n60 0.189894
R1950 VN.n102 VN.n60 0.189894
R1951 VN.n102 VN.n101 0.189894
R1952 VN.n101 VN.n100 0.189894
R1953 VN.n100 VN.n62 0.189894
R1954 VN.n95 VN.n62 0.189894
R1955 VN.n95 VN.n94 0.189894
R1956 VN.n94 VN.n93 0.189894
R1957 VN.n93 VN.n64 0.189894
R1958 VN.n89 VN.n64 0.189894
R1959 VN.n89 VN.n88 0.189894
R1960 VN.n88 VN.n87 0.189894
R1961 VN.n87 VN.n66 0.189894
R1962 VN.n83 VN.n66 0.189894
R1963 VN.n83 VN.n82 0.189894
R1964 VN.n82 VN.n81 0.189894
R1965 VN.n81 VN.n68 0.189894
R1966 VN.n77 VN.n68 0.189894
R1967 VN.n77 VN.n76 0.189894
R1968 VN.n76 VN.n75 0.189894
R1969 VN.n75 VN.n70 0.189894
R1970 VN.n18 VN.n13 0.189894
R1971 VN.n19 VN.n18 0.189894
R1972 VN.n20 VN.n19 0.189894
R1973 VN.n20 VN.n11 0.189894
R1974 VN.n24 VN.n11 0.189894
R1975 VN.n25 VN.n24 0.189894
R1976 VN.n26 VN.n25 0.189894
R1977 VN.n26 VN.n9 0.189894
R1978 VN.n30 VN.n9 0.189894
R1979 VN.n31 VN.n30 0.189894
R1980 VN.n32 VN.n31 0.189894
R1981 VN.n32 VN.n7 0.189894
R1982 VN.n36 VN.n7 0.189894
R1983 VN.n37 VN.n36 0.189894
R1984 VN.n38 VN.n37 0.189894
R1985 VN.n38 VN.n5 0.189894
R1986 VN.n43 VN.n5 0.189894
R1987 VN.n44 VN.n43 0.189894
R1988 VN.n45 VN.n44 0.189894
R1989 VN.n45 VN.n3 0.189894
R1990 VN.n49 VN.n3 0.189894
R1991 VN.n50 VN.n49 0.189894
R1992 VN.n51 VN.n50 0.189894
R1993 VN.n51 VN.n1 0.189894
R1994 VN.n55 VN.n1 0.189894
R1995 VDD2.n1 VDD2.t3 80.0263
R1996 VDD2.n4 VDD2.t9 76.3368
R1997 VDD2.n3 VDD2.n2 76.0773
R1998 VDD2 VDD2.n7 76.0745
R1999 VDD2.n6 VDD2.n5 73.3657
R2000 VDD2.n1 VDD2.n0 73.3654
R2001 VDD2.n4 VDD2.n3 50.6722
R2002 VDD2.n6 VDD2.n4 3.69016
R2003 VDD2.n7 VDD2.t2 2.97171
R2004 VDD2.n7 VDD2.t6 2.97171
R2005 VDD2.n5 VDD2.t1 2.97171
R2006 VDD2.n5 VDD2.t5 2.97171
R2007 VDD2.n2 VDD2.t7 2.97171
R2008 VDD2.n2 VDD2.t4 2.97171
R2009 VDD2.n0 VDD2.t0 2.97171
R2010 VDD2.n0 VDD2.t8 2.97171
R2011 VDD2 VDD2.n6 0.981103
R2012 VDD2.n3 VDD2.n1 0.867568
C0 B w_n6106_n3156# 12.519099f
C1 VDD2 w_n6106_n3156# 3.4381f
C2 VP w_n6106_n3156# 14.226701f
C3 B VDD1 2.9178f
C4 VDD2 VDD1 3.05375f
C5 VP VDD1 11.069201f
C6 B VTAIL 3.97798f
C7 VDD2 VTAIL 10.782401f
C8 B VN 1.61924f
C9 VDD2 VN 10.4738f
C10 VP VTAIL 11.7611f
C11 VDD1 w_n6106_n3156# 3.22439f
C12 VP VN 10.1818f
C13 w_n6106_n3156# VTAIL 3.26107f
C14 w_n6106_n3156# VN 13.4276f
C15 VDD1 VTAIL 10.7212f
C16 VDD1 VN 0.15675f
C17 VDD2 B 3.08828f
C18 VTAIL VN 11.7463f
C19 VP B 2.97048f
C20 VP VDD2 0.755491f
C21 VDD2 VSUBS 2.68972f
C22 VDD1 VSUBS 2.515067f
C23 VTAIL VSUBS 1.595989f
C24 VN VSUBS 9.951509f
C25 VP VSUBS 5.918024f
C26 B VSUBS 6.949979f
C27 w_n6106_n3156# VSUBS 0.237621p
C28 VDD2.t3 VSUBS 2.81618f
C29 VDD2.t0 VSUBS 0.276356f
C30 VDD2.t8 VSUBS 0.276356f
C31 VDD2.n0 VSUBS 2.11298f
C32 VDD2.n1 VSUBS 2.1095f
C33 VDD2.t7 VSUBS 0.276356f
C34 VDD2.t4 VSUBS 0.276356f
C35 VDD2.n2 VSUBS 2.15826f
C36 VDD2.n3 VSUBS 4.8558f
C37 VDD2.t9 VSUBS 2.76586f
C38 VDD2.n4 VSUBS 4.9157f
C39 VDD2.t1 VSUBS 0.276356f
C40 VDD2.t5 VSUBS 0.276356f
C41 VDD2.n5 VSUBS 2.11298f
C42 VDD2.n6 VSUBS 1.07898f
C43 VDD2.t2 VSUBS 0.276356f
C44 VDD2.t6 VSUBS 0.276356f
C45 VDD2.n7 VSUBS 2.15819f
C46 VN.t5 VSUBS 2.7584f
C47 VN.n0 VSUBS 1.06078f
C48 VN.n1 VSUBS 0.023493f
C49 VN.n2 VSUBS 0.047127f
C50 VN.n3 VSUBS 0.023493f
C51 VN.n4 VSUBS 0.043566f
C52 VN.n5 VSUBS 0.023493f
C53 VN.t2 VSUBS 2.7584f
C54 VN.n6 VSUBS 0.043566f
C55 VN.n7 VSUBS 0.023493f
C56 VN.n8 VSUBS 0.043566f
C57 VN.n9 VSUBS 0.023493f
C58 VN.t1 VSUBS 2.7584f
C59 VN.n10 VSUBS 0.043566f
C60 VN.n11 VSUBS 0.023493f
C61 VN.n12 VSUBS 0.043566f
C62 VN.n13 VSUBS 0.306103f
C63 VN.t9 VSUBS 2.7584f
C64 VN.t6 VSUBS 3.1414f
C65 VN.n14 VSUBS 1.00312f
C66 VN.n15 VSUBS 1.05611f
C67 VN.n16 VSUBS 0.034103f
C68 VN.n17 VSUBS 0.043566f
C69 VN.n18 VSUBS 0.023493f
C70 VN.n19 VSUBS 0.023493f
C71 VN.n20 VSUBS 0.023493f
C72 VN.n21 VSUBS 0.040984f
C73 VN.n22 VSUBS 0.025583f
C74 VN.n23 VSUBS 0.045301f
C75 VN.n24 VSUBS 0.023493f
C76 VN.n25 VSUBS 0.023493f
C77 VN.n26 VSUBS 0.023493f
C78 VN.n27 VSUBS 0.043566f
C79 VN.n28 VSUBS 0.99193f
C80 VN.n29 VSUBS 0.043566f
C81 VN.n30 VSUBS 0.023493f
C82 VN.n31 VSUBS 0.023493f
C83 VN.n32 VSUBS 0.023493f
C84 VN.n33 VSUBS 0.045301f
C85 VN.n34 VSUBS 0.025583f
C86 VN.n35 VSUBS 0.040984f
C87 VN.n36 VSUBS 0.023493f
C88 VN.n37 VSUBS 0.023493f
C89 VN.n38 VSUBS 0.023493f
C90 VN.n39 VSUBS 0.043566f
C91 VN.n40 VSUBS 0.034103f
C92 VN.n41 VSUBS 0.969871f
C93 VN.n42 VSUBS 0.031522f
C94 VN.n43 VSUBS 0.023493f
C95 VN.n44 VSUBS 0.023493f
C96 VN.n45 VSUBS 0.023493f
C97 VN.n46 VSUBS 0.043566f
C98 VN.n47 VSUBS 0.043777f
C99 VN.n48 VSUBS 0.020964f
C100 VN.n49 VSUBS 0.023493f
C101 VN.n50 VSUBS 0.023493f
C102 VN.n51 VSUBS 0.023493f
C103 VN.n52 VSUBS 0.043566f
C104 VN.n53 VSUBS 0.043566f
C105 VN.n54 VSUBS 0.024639f
C106 VN.n55 VSUBS 0.037912f
C107 VN.n56 VSUBS 0.07399f
C108 VN.t0 VSUBS 2.7584f
C109 VN.n57 VSUBS 1.06078f
C110 VN.n58 VSUBS 0.023493f
C111 VN.n59 VSUBS 0.047127f
C112 VN.n60 VSUBS 0.023493f
C113 VN.n61 VSUBS 0.043566f
C114 VN.n62 VSUBS 0.023493f
C115 VN.t8 VSUBS 2.7584f
C116 VN.n63 VSUBS 0.043566f
C117 VN.n64 VSUBS 0.023493f
C118 VN.n65 VSUBS 0.043566f
C119 VN.n66 VSUBS 0.023493f
C120 VN.t4 VSUBS 2.7584f
C121 VN.n67 VSUBS 0.043566f
C122 VN.n68 VSUBS 0.023493f
C123 VN.n69 VSUBS 0.043566f
C124 VN.n70 VSUBS 0.306103f
C125 VN.t7 VSUBS 2.7584f
C126 VN.t3 VSUBS 3.1414f
C127 VN.n71 VSUBS 1.00312f
C128 VN.n72 VSUBS 1.05611f
C129 VN.n73 VSUBS 0.034103f
C130 VN.n74 VSUBS 0.043566f
C131 VN.n75 VSUBS 0.023493f
C132 VN.n76 VSUBS 0.023493f
C133 VN.n77 VSUBS 0.023493f
C134 VN.n78 VSUBS 0.040984f
C135 VN.n79 VSUBS 0.025583f
C136 VN.n80 VSUBS 0.045301f
C137 VN.n81 VSUBS 0.023493f
C138 VN.n82 VSUBS 0.023493f
C139 VN.n83 VSUBS 0.023493f
C140 VN.n84 VSUBS 0.043566f
C141 VN.n85 VSUBS 0.99193f
C142 VN.n86 VSUBS 0.043566f
C143 VN.n87 VSUBS 0.023493f
C144 VN.n88 VSUBS 0.023493f
C145 VN.n89 VSUBS 0.023493f
C146 VN.n90 VSUBS 0.045301f
C147 VN.n91 VSUBS 0.025583f
C148 VN.n92 VSUBS 0.040984f
C149 VN.n93 VSUBS 0.023493f
C150 VN.n94 VSUBS 0.023493f
C151 VN.n95 VSUBS 0.023493f
C152 VN.n96 VSUBS 0.043566f
C153 VN.n97 VSUBS 0.034103f
C154 VN.n98 VSUBS 0.969871f
C155 VN.n99 VSUBS 0.031522f
C156 VN.n100 VSUBS 0.023493f
C157 VN.n101 VSUBS 0.023493f
C158 VN.n102 VSUBS 0.023493f
C159 VN.n103 VSUBS 0.043566f
C160 VN.n104 VSUBS 0.043777f
C161 VN.n105 VSUBS 0.020964f
C162 VN.n106 VSUBS 0.023493f
C163 VN.n107 VSUBS 0.023493f
C164 VN.n108 VSUBS 0.023493f
C165 VN.n109 VSUBS 0.043566f
C166 VN.n110 VSUBS 0.043566f
C167 VN.n111 VSUBS 0.024639f
C168 VN.n112 VSUBS 0.037912f
C169 VN.n113 VSUBS 1.73801f
C170 B.n0 VSUBS 0.008039f
C171 B.n1 VSUBS 0.008039f
C172 B.n2 VSUBS 0.011889f
C173 B.n3 VSUBS 0.00911f
C174 B.n4 VSUBS 0.00911f
C175 B.n5 VSUBS 0.00911f
C176 B.n6 VSUBS 0.00911f
C177 B.n7 VSUBS 0.00911f
C178 B.n8 VSUBS 0.00911f
C179 B.n9 VSUBS 0.00911f
C180 B.n10 VSUBS 0.00911f
C181 B.n11 VSUBS 0.00911f
C182 B.n12 VSUBS 0.00911f
C183 B.n13 VSUBS 0.00911f
C184 B.n14 VSUBS 0.00911f
C185 B.n15 VSUBS 0.00911f
C186 B.n16 VSUBS 0.00911f
C187 B.n17 VSUBS 0.00911f
C188 B.n18 VSUBS 0.00911f
C189 B.n19 VSUBS 0.00911f
C190 B.n20 VSUBS 0.00911f
C191 B.n21 VSUBS 0.00911f
C192 B.n22 VSUBS 0.00911f
C193 B.n23 VSUBS 0.00911f
C194 B.n24 VSUBS 0.00911f
C195 B.n25 VSUBS 0.00911f
C196 B.n26 VSUBS 0.00911f
C197 B.n27 VSUBS 0.00911f
C198 B.n28 VSUBS 0.00911f
C199 B.n29 VSUBS 0.00911f
C200 B.n30 VSUBS 0.00911f
C201 B.n31 VSUBS 0.00911f
C202 B.n32 VSUBS 0.00911f
C203 B.n33 VSUBS 0.00911f
C204 B.n34 VSUBS 0.00911f
C205 B.n35 VSUBS 0.00911f
C206 B.n36 VSUBS 0.00911f
C207 B.n37 VSUBS 0.00911f
C208 B.n38 VSUBS 0.00911f
C209 B.n39 VSUBS 0.00911f
C210 B.n40 VSUBS 0.00911f
C211 B.n41 VSUBS 0.00911f
C212 B.n42 VSUBS 0.00911f
C213 B.n43 VSUBS 0.020048f
C214 B.n44 VSUBS 0.00911f
C215 B.n45 VSUBS 0.00911f
C216 B.n46 VSUBS 0.00911f
C217 B.n47 VSUBS 0.00911f
C218 B.n48 VSUBS 0.00911f
C219 B.n49 VSUBS 0.00911f
C220 B.n50 VSUBS 0.00911f
C221 B.n51 VSUBS 0.00911f
C222 B.n52 VSUBS 0.00911f
C223 B.n53 VSUBS 0.00911f
C224 B.n54 VSUBS 0.00911f
C225 B.n55 VSUBS 0.00911f
C226 B.n56 VSUBS 0.00911f
C227 B.n57 VSUBS 0.00911f
C228 B.n58 VSUBS 0.00911f
C229 B.n59 VSUBS 0.00911f
C230 B.n60 VSUBS 0.00911f
C231 B.n61 VSUBS 0.00911f
C232 B.n62 VSUBS 0.00911f
C233 B.n63 VSUBS 0.00911f
C234 B.t1 VSUBS 0.459185f
C235 B.t2 VSUBS 0.49716f
C236 B.t0 VSUBS 2.6409f
C237 B.n64 VSUBS 0.286187f
C238 B.n65 VSUBS 0.10062f
C239 B.n66 VSUBS 0.00911f
C240 B.n67 VSUBS 0.00911f
C241 B.n68 VSUBS 0.00911f
C242 B.n69 VSUBS 0.00911f
C243 B.t4 VSUBS 0.459177f
C244 B.t5 VSUBS 0.497153f
C245 B.t3 VSUBS 2.6409f
C246 B.n70 VSUBS 0.286194f
C247 B.n71 VSUBS 0.100628f
C248 B.n72 VSUBS 0.00911f
C249 B.n73 VSUBS 0.00911f
C250 B.n74 VSUBS 0.00911f
C251 B.n75 VSUBS 0.00911f
C252 B.n76 VSUBS 0.00911f
C253 B.n77 VSUBS 0.00911f
C254 B.n78 VSUBS 0.00911f
C255 B.n79 VSUBS 0.00911f
C256 B.n80 VSUBS 0.00911f
C257 B.n81 VSUBS 0.00911f
C258 B.n82 VSUBS 0.00911f
C259 B.n83 VSUBS 0.00911f
C260 B.n84 VSUBS 0.00911f
C261 B.n85 VSUBS 0.00911f
C262 B.n86 VSUBS 0.00911f
C263 B.n87 VSUBS 0.00911f
C264 B.n88 VSUBS 0.00911f
C265 B.n89 VSUBS 0.00911f
C266 B.n90 VSUBS 0.00911f
C267 B.n91 VSUBS 0.020048f
C268 B.n92 VSUBS 0.00911f
C269 B.n93 VSUBS 0.00911f
C270 B.n94 VSUBS 0.00911f
C271 B.n95 VSUBS 0.00911f
C272 B.n96 VSUBS 0.00911f
C273 B.n97 VSUBS 0.00911f
C274 B.n98 VSUBS 0.00911f
C275 B.n99 VSUBS 0.00911f
C276 B.n100 VSUBS 0.00911f
C277 B.n101 VSUBS 0.00911f
C278 B.n102 VSUBS 0.00911f
C279 B.n103 VSUBS 0.00911f
C280 B.n104 VSUBS 0.00911f
C281 B.n105 VSUBS 0.00911f
C282 B.n106 VSUBS 0.00911f
C283 B.n107 VSUBS 0.00911f
C284 B.n108 VSUBS 0.00911f
C285 B.n109 VSUBS 0.00911f
C286 B.n110 VSUBS 0.00911f
C287 B.n111 VSUBS 0.00911f
C288 B.n112 VSUBS 0.00911f
C289 B.n113 VSUBS 0.00911f
C290 B.n114 VSUBS 0.00911f
C291 B.n115 VSUBS 0.00911f
C292 B.n116 VSUBS 0.00911f
C293 B.n117 VSUBS 0.00911f
C294 B.n118 VSUBS 0.00911f
C295 B.n119 VSUBS 0.00911f
C296 B.n120 VSUBS 0.00911f
C297 B.n121 VSUBS 0.00911f
C298 B.n122 VSUBS 0.00911f
C299 B.n123 VSUBS 0.00911f
C300 B.n124 VSUBS 0.00911f
C301 B.n125 VSUBS 0.00911f
C302 B.n126 VSUBS 0.00911f
C303 B.n127 VSUBS 0.00911f
C304 B.n128 VSUBS 0.00911f
C305 B.n129 VSUBS 0.00911f
C306 B.n130 VSUBS 0.00911f
C307 B.n131 VSUBS 0.00911f
C308 B.n132 VSUBS 0.00911f
C309 B.n133 VSUBS 0.00911f
C310 B.n134 VSUBS 0.00911f
C311 B.n135 VSUBS 0.00911f
C312 B.n136 VSUBS 0.00911f
C313 B.n137 VSUBS 0.00911f
C314 B.n138 VSUBS 0.00911f
C315 B.n139 VSUBS 0.00911f
C316 B.n140 VSUBS 0.00911f
C317 B.n141 VSUBS 0.00911f
C318 B.n142 VSUBS 0.00911f
C319 B.n143 VSUBS 0.00911f
C320 B.n144 VSUBS 0.00911f
C321 B.n145 VSUBS 0.00911f
C322 B.n146 VSUBS 0.00911f
C323 B.n147 VSUBS 0.00911f
C324 B.n148 VSUBS 0.00911f
C325 B.n149 VSUBS 0.00911f
C326 B.n150 VSUBS 0.00911f
C327 B.n151 VSUBS 0.00911f
C328 B.n152 VSUBS 0.00911f
C329 B.n153 VSUBS 0.00911f
C330 B.n154 VSUBS 0.00911f
C331 B.n155 VSUBS 0.00911f
C332 B.n156 VSUBS 0.00911f
C333 B.n157 VSUBS 0.00911f
C334 B.n158 VSUBS 0.00911f
C335 B.n159 VSUBS 0.00911f
C336 B.n160 VSUBS 0.00911f
C337 B.n161 VSUBS 0.00911f
C338 B.n162 VSUBS 0.00911f
C339 B.n163 VSUBS 0.00911f
C340 B.n164 VSUBS 0.00911f
C341 B.n165 VSUBS 0.00911f
C342 B.n166 VSUBS 0.00911f
C343 B.n167 VSUBS 0.00911f
C344 B.n168 VSUBS 0.00911f
C345 B.n169 VSUBS 0.00911f
C346 B.n170 VSUBS 0.00911f
C347 B.n171 VSUBS 0.00911f
C348 B.n172 VSUBS 0.00911f
C349 B.n173 VSUBS 0.00911f
C350 B.n174 VSUBS 0.00911f
C351 B.n175 VSUBS 0.021753f
C352 B.n176 VSUBS 0.00911f
C353 B.n177 VSUBS 0.00911f
C354 B.n178 VSUBS 0.00911f
C355 B.n179 VSUBS 0.00911f
C356 B.n180 VSUBS 0.00911f
C357 B.n181 VSUBS 0.00911f
C358 B.n182 VSUBS 0.00911f
C359 B.n183 VSUBS 0.00911f
C360 B.n184 VSUBS 0.00911f
C361 B.n185 VSUBS 0.00911f
C362 B.n186 VSUBS 0.00911f
C363 B.n187 VSUBS 0.00911f
C364 B.n188 VSUBS 0.00911f
C365 B.n189 VSUBS 0.00911f
C366 B.n190 VSUBS 0.00911f
C367 B.n191 VSUBS 0.00911f
C368 B.n192 VSUBS 0.00911f
C369 B.n193 VSUBS 0.00911f
C370 B.n194 VSUBS 0.006297f
C371 B.n195 VSUBS 0.00911f
C372 B.n196 VSUBS 0.00911f
C373 B.n197 VSUBS 0.00911f
C374 B.n198 VSUBS 0.00911f
C375 B.n199 VSUBS 0.00911f
C376 B.t8 VSUBS 0.459185f
C377 B.t7 VSUBS 0.49716f
C378 B.t6 VSUBS 2.6409f
C379 B.n200 VSUBS 0.286187f
C380 B.n201 VSUBS 0.10062f
C381 B.n202 VSUBS 0.00911f
C382 B.n203 VSUBS 0.00911f
C383 B.n204 VSUBS 0.00911f
C384 B.n205 VSUBS 0.00911f
C385 B.n206 VSUBS 0.00911f
C386 B.n207 VSUBS 0.00911f
C387 B.n208 VSUBS 0.00911f
C388 B.n209 VSUBS 0.00911f
C389 B.n210 VSUBS 0.00911f
C390 B.n211 VSUBS 0.00911f
C391 B.n212 VSUBS 0.00911f
C392 B.n213 VSUBS 0.00911f
C393 B.n214 VSUBS 0.00911f
C394 B.n215 VSUBS 0.00911f
C395 B.n216 VSUBS 0.00911f
C396 B.n217 VSUBS 0.00911f
C397 B.n218 VSUBS 0.00911f
C398 B.n219 VSUBS 0.00911f
C399 B.n220 VSUBS 0.021753f
C400 B.n221 VSUBS 0.00911f
C401 B.n222 VSUBS 0.00911f
C402 B.n223 VSUBS 0.00911f
C403 B.n224 VSUBS 0.00911f
C404 B.n225 VSUBS 0.00911f
C405 B.n226 VSUBS 0.00911f
C406 B.n227 VSUBS 0.00911f
C407 B.n228 VSUBS 0.00911f
C408 B.n229 VSUBS 0.00911f
C409 B.n230 VSUBS 0.00911f
C410 B.n231 VSUBS 0.00911f
C411 B.n232 VSUBS 0.00911f
C412 B.n233 VSUBS 0.00911f
C413 B.n234 VSUBS 0.00911f
C414 B.n235 VSUBS 0.00911f
C415 B.n236 VSUBS 0.00911f
C416 B.n237 VSUBS 0.00911f
C417 B.n238 VSUBS 0.00911f
C418 B.n239 VSUBS 0.00911f
C419 B.n240 VSUBS 0.00911f
C420 B.n241 VSUBS 0.00911f
C421 B.n242 VSUBS 0.00911f
C422 B.n243 VSUBS 0.00911f
C423 B.n244 VSUBS 0.00911f
C424 B.n245 VSUBS 0.00911f
C425 B.n246 VSUBS 0.00911f
C426 B.n247 VSUBS 0.00911f
C427 B.n248 VSUBS 0.00911f
C428 B.n249 VSUBS 0.00911f
C429 B.n250 VSUBS 0.00911f
C430 B.n251 VSUBS 0.00911f
C431 B.n252 VSUBS 0.00911f
C432 B.n253 VSUBS 0.00911f
C433 B.n254 VSUBS 0.00911f
C434 B.n255 VSUBS 0.00911f
C435 B.n256 VSUBS 0.00911f
C436 B.n257 VSUBS 0.00911f
C437 B.n258 VSUBS 0.00911f
C438 B.n259 VSUBS 0.00911f
C439 B.n260 VSUBS 0.00911f
C440 B.n261 VSUBS 0.00911f
C441 B.n262 VSUBS 0.00911f
C442 B.n263 VSUBS 0.00911f
C443 B.n264 VSUBS 0.00911f
C444 B.n265 VSUBS 0.00911f
C445 B.n266 VSUBS 0.00911f
C446 B.n267 VSUBS 0.00911f
C447 B.n268 VSUBS 0.00911f
C448 B.n269 VSUBS 0.00911f
C449 B.n270 VSUBS 0.00911f
C450 B.n271 VSUBS 0.00911f
C451 B.n272 VSUBS 0.00911f
C452 B.n273 VSUBS 0.00911f
C453 B.n274 VSUBS 0.00911f
C454 B.n275 VSUBS 0.00911f
C455 B.n276 VSUBS 0.00911f
C456 B.n277 VSUBS 0.00911f
C457 B.n278 VSUBS 0.00911f
C458 B.n279 VSUBS 0.00911f
C459 B.n280 VSUBS 0.00911f
C460 B.n281 VSUBS 0.00911f
C461 B.n282 VSUBS 0.00911f
C462 B.n283 VSUBS 0.00911f
C463 B.n284 VSUBS 0.00911f
C464 B.n285 VSUBS 0.00911f
C465 B.n286 VSUBS 0.00911f
C466 B.n287 VSUBS 0.00911f
C467 B.n288 VSUBS 0.00911f
C468 B.n289 VSUBS 0.00911f
C469 B.n290 VSUBS 0.00911f
C470 B.n291 VSUBS 0.00911f
C471 B.n292 VSUBS 0.00911f
C472 B.n293 VSUBS 0.00911f
C473 B.n294 VSUBS 0.00911f
C474 B.n295 VSUBS 0.00911f
C475 B.n296 VSUBS 0.00911f
C476 B.n297 VSUBS 0.00911f
C477 B.n298 VSUBS 0.00911f
C478 B.n299 VSUBS 0.00911f
C479 B.n300 VSUBS 0.00911f
C480 B.n301 VSUBS 0.00911f
C481 B.n302 VSUBS 0.00911f
C482 B.n303 VSUBS 0.00911f
C483 B.n304 VSUBS 0.00911f
C484 B.n305 VSUBS 0.00911f
C485 B.n306 VSUBS 0.00911f
C486 B.n307 VSUBS 0.00911f
C487 B.n308 VSUBS 0.00911f
C488 B.n309 VSUBS 0.00911f
C489 B.n310 VSUBS 0.00911f
C490 B.n311 VSUBS 0.00911f
C491 B.n312 VSUBS 0.00911f
C492 B.n313 VSUBS 0.00911f
C493 B.n314 VSUBS 0.00911f
C494 B.n315 VSUBS 0.00911f
C495 B.n316 VSUBS 0.00911f
C496 B.n317 VSUBS 0.00911f
C497 B.n318 VSUBS 0.00911f
C498 B.n319 VSUBS 0.00911f
C499 B.n320 VSUBS 0.00911f
C500 B.n321 VSUBS 0.00911f
C501 B.n322 VSUBS 0.00911f
C502 B.n323 VSUBS 0.00911f
C503 B.n324 VSUBS 0.00911f
C504 B.n325 VSUBS 0.00911f
C505 B.n326 VSUBS 0.00911f
C506 B.n327 VSUBS 0.00911f
C507 B.n328 VSUBS 0.00911f
C508 B.n329 VSUBS 0.00911f
C509 B.n330 VSUBS 0.00911f
C510 B.n331 VSUBS 0.00911f
C511 B.n332 VSUBS 0.00911f
C512 B.n333 VSUBS 0.00911f
C513 B.n334 VSUBS 0.00911f
C514 B.n335 VSUBS 0.00911f
C515 B.n336 VSUBS 0.00911f
C516 B.n337 VSUBS 0.00911f
C517 B.n338 VSUBS 0.00911f
C518 B.n339 VSUBS 0.00911f
C519 B.n340 VSUBS 0.00911f
C520 B.n341 VSUBS 0.00911f
C521 B.n342 VSUBS 0.00911f
C522 B.n343 VSUBS 0.00911f
C523 B.n344 VSUBS 0.00911f
C524 B.n345 VSUBS 0.00911f
C525 B.n346 VSUBS 0.00911f
C526 B.n347 VSUBS 0.00911f
C527 B.n348 VSUBS 0.00911f
C528 B.n349 VSUBS 0.00911f
C529 B.n350 VSUBS 0.00911f
C530 B.n351 VSUBS 0.00911f
C531 B.n352 VSUBS 0.00911f
C532 B.n353 VSUBS 0.00911f
C533 B.n354 VSUBS 0.00911f
C534 B.n355 VSUBS 0.00911f
C535 B.n356 VSUBS 0.00911f
C536 B.n357 VSUBS 0.00911f
C537 B.n358 VSUBS 0.00911f
C538 B.n359 VSUBS 0.00911f
C539 B.n360 VSUBS 0.00911f
C540 B.n361 VSUBS 0.00911f
C541 B.n362 VSUBS 0.00911f
C542 B.n363 VSUBS 0.00911f
C543 B.n364 VSUBS 0.00911f
C544 B.n365 VSUBS 0.00911f
C545 B.n366 VSUBS 0.00911f
C546 B.n367 VSUBS 0.00911f
C547 B.n368 VSUBS 0.00911f
C548 B.n369 VSUBS 0.00911f
C549 B.n370 VSUBS 0.00911f
C550 B.n371 VSUBS 0.00911f
C551 B.n372 VSUBS 0.00911f
C552 B.n373 VSUBS 0.00911f
C553 B.n374 VSUBS 0.00911f
C554 B.n375 VSUBS 0.00911f
C555 B.n376 VSUBS 0.00911f
C556 B.n377 VSUBS 0.00911f
C557 B.n378 VSUBS 0.00911f
C558 B.n379 VSUBS 0.00911f
C559 B.n380 VSUBS 0.00911f
C560 B.n381 VSUBS 0.00911f
C561 B.n382 VSUBS 0.00911f
C562 B.n383 VSUBS 0.020048f
C563 B.n384 VSUBS 0.020048f
C564 B.n385 VSUBS 0.021753f
C565 B.n386 VSUBS 0.00911f
C566 B.n387 VSUBS 0.00911f
C567 B.n388 VSUBS 0.00911f
C568 B.n389 VSUBS 0.00911f
C569 B.n390 VSUBS 0.00911f
C570 B.n391 VSUBS 0.00911f
C571 B.n392 VSUBS 0.00911f
C572 B.n393 VSUBS 0.00911f
C573 B.n394 VSUBS 0.00911f
C574 B.n395 VSUBS 0.00911f
C575 B.n396 VSUBS 0.00911f
C576 B.n397 VSUBS 0.00911f
C577 B.n398 VSUBS 0.00911f
C578 B.n399 VSUBS 0.00911f
C579 B.n400 VSUBS 0.00911f
C580 B.n401 VSUBS 0.00911f
C581 B.n402 VSUBS 0.00911f
C582 B.n403 VSUBS 0.00911f
C583 B.n404 VSUBS 0.00911f
C584 B.n405 VSUBS 0.00911f
C585 B.n406 VSUBS 0.00911f
C586 B.n407 VSUBS 0.00911f
C587 B.n408 VSUBS 0.00911f
C588 B.n409 VSUBS 0.00911f
C589 B.n410 VSUBS 0.00911f
C590 B.n411 VSUBS 0.00911f
C591 B.n412 VSUBS 0.00911f
C592 B.n413 VSUBS 0.00911f
C593 B.n414 VSUBS 0.00911f
C594 B.n415 VSUBS 0.00911f
C595 B.n416 VSUBS 0.00911f
C596 B.n417 VSUBS 0.00911f
C597 B.n418 VSUBS 0.00911f
C598 B.n419 VSUBS 0.00911f
C599 B.n420 VSUBS 0.00911f
C600 B.n421 VSUBS 0.00911f
C601 B.n422 VSUBS 0.00911f
C602 B.n423 VSUBS 0.00911f
C603 B.n424 VSUBS 0.00911f
C604 B.n425 VSUBS 0.00911f
C605 B.n426 VSUBS 0.00911f
C606 B.n427 VSUBS 0.00911f
C607 B.n428 VSUBS 0.00911f
C608 B.n429 VSUBS 0.00911f
C609 B.n430 VSUBS 0.00911f
C610 B.n431 VSUBS 0.00911f
C611 B.n432 VSUBS 0.00911f
C612 B.n433 VSUBS 0.00911f
C613 B.n434 VSUBS 0.00911f
C614 B.n435 VSUBS 0.00911f
C615 B.n436 VSUBS 0.00911f
C616 B.n437 VSUBS 0.00911f
C617 B.n438 VSUBS 0.00911f
C618 B.n439 VSUBS 0.00911f
C619 B.n440 VSUBS 0.00911f
C620 B.n441 VSUBS 0.00911f
C621 B.n442 VSUBS 0.006297f
C622 B.n443 VSUBS 0.021108f
C623 B.n444 VSUBS 0.007369f
C624 B.n445 VSUBS 0.00911f
C625 B.n446 VSUBS 0.00911f
C626 B.n447 VSUBS 0.00911f
C627 B.n448 VSUBS 0.00911f
C628 B.n449 VSUBS 0.00911f
C629 B.n450 VSUBS 0.00911f
C630 B.n451 VSUBS 0.00911f
C631 B.n452 VSUBS 0.00911f
C632 B.n453 VSUBS 0.00911f
C633 B.n454 VSUBS 0.00911f
C634 B.n455 VSUBS 0.00911f
C635 B.t11 VSUBS 0.459177f
C636 B.t10 VSUBS 0.497153f
C637 B.t9 VSUBS 2.6409f
C638 B.n456 VSUBS 0.286194f
C639 B.n457 VSUBS 0.100628f
C640 B.n458 VSUBS 0.021108f
C641 B.n459 VSUBS 0.007369f
C642 B.n460 VSUBS 0.00911f
C643 B.n461 VSUBS 0.00911f
C644 B.n462 VSUBS 0.00911f
C645 B.n463 VSUBS 0.00911f
C646 B.n464 VSUBS 0.00911f
C647 B.n465 VSUBS 0.00911f
C648 B.n466 VSUBS 0.00911f
C649 B.n467 VSUBS 0.00911f
C650 B.n468 VSUBS 0.00911f
C651 B.n469 VSUBS 0.00911f
C652 B.n470 VSUBS 0.00911f
C653 B.n471 VSUBS 0.00911f
C654 B.n472 VSUBS 0.00911f
C655 B.n473 VSUBS 0.00911f
C656 B.n474 VSUBS 0.00911f
C657 B.n475 VSUBS 0.00911f
C658 B.n476 VSUBS 0.00911f
C659 B.n477 VSUBS 0.00911f
C660 B.n478 VSUBS 0.00911f
C661 B.n479 VSUBS 0.00911f
C662 B.n480 VSUBS 0.00911f
C663 B.n481 VSUBS 0.00911f
C664 B.n482 VSUBS 0.00911f
C665 B.n483 VSUBS 0.00911f
C666 B.n484 VSUBS 0.00911f
C667 B.n485 VSUBS 0.00911f
C668 B.n486 VSUBS 0.00911f
C669 B.n487 VSUBS 0.00911f
C670 B.n488 VSUBS 0.00911f
C671 B.n489 VSUBS 0.00911f
C672 B.n490 VSUBS 0.00911f
C673 B.n491 VSUBS 0.00911f
C674 B.n492 VSUBS 0.00911f
C675 B.n493 VSUBS 0.00911f
C676 B.n494 VSUBS 0.00911f
C677 B.n495 VSUBS 0.00911f
C678 B.n496 VSUBS 0.00911f
C679 B.n497 VSUBS 0.00911f
C680 B.n498 VSUBS 0.00911f
C681 B.n499 VSUBS 0.00911f
C682 B.n500 VSUBS 0.00911f
C683 B.n501 VSUBS 0.00911f
C684 B.n502 VSUBS 0.00911f
C685 B.n503 VSUBS 0.00911f
C686 B.n504 VSUBS 0.00911f
C687 B.n505 VSUBS 0.00911f
C688 B.n506 VSUBS 0.00911f
C689 B.n507 VSUBS 0.00911f
C690 B.n508 VSUBS 0.00911f
C691 B.n509 VSUBS 0.00911f
C692 B.n510 VSUBS 0.00911f
C693 B.n511 VSUBS 0.00911f
C694 B.n512 VSUBS 0.00911f
C695 B.n513 VSUBS 0.00911f
C696 B.n514 VSUBS 0.00911f
C697 B.n515 VSUBS 0.00911f
C698 B.n516 VSUBS 0.00911f
C699 B.n517 VSUBS 0.00911f
C700 B.n518 VSUBS 0.020643f
C701 B.n519 VSUBS 0.021157f
C702 B.n520 VSUBS 0.020048f
C703 B.n521 VSUBS 0.00911f
C704 B.n522 VSUBS 0.00911f
C705 B.n523 VSUBS 0.00911f
C706 B.n524 VSUBS 0.00911f
C707 B.n525 VSUBS 0.00911f
C708 B.n526 VSUBS 0.00911f
C709 B.n527 VSUBS 0.00911f
C710 B.n528 VSUBS 0.00911f
C711 B.n529 VSUBS 0.00911f
C712 B.n530 VSUBS 0.00911f
C713 B.n531 VSUBS 0.00911f
C714 B.n532 VSUBS 0.00911f
C715 B.n533 VSUBS 0.00911f
C716 B.n534 VSUBS 0.00911f
C717 B.n535 VSUBS 0.00911f
C718 B.n536 VSUBS 0.00911f
C719 B.n537 VSUBS 0.00911f
C720 B.n538 VSUBS 0.00911f
C721 B.n539 VSUBS 0.00911f
C722 B.n540 VSUBS 0.00911f
C723 B.n541 VSUBS 0.00911f
C724 B.n542 VSUBS 0.00911f
C725 B.n543 VSUBS 0.00911f
C726 B.n544 VSUBS 0.00911f
C727 B.n545 VSUBS 0.00911f
C728 B.n546 VSUBS 0.00911f
C729 B.n547 VSUBS 0.00911f
C730 B.n548 VSUBS 0.00911f
C731 B.n549 VSUBS 0.00911f
C732 B.n550 VSUBS 0.00911f
C733 B.n551 VSUBS 0.00911f
C734 B.n552 VSUBS 0.00911f
C735 B.n553 VSUBS 0.00911f
C736 B.n554 VSUBS 0.00911f
C737 B.n555 VSUBS 0.00911f
C738 B.n556 VSUBS 0.00911f
C739 B.n557 VSUBS 0.00911f
C740 B.n558 VSUBS 0.00911f
C741 B.n559 VSUBS 0.00911f
C742 B.n560 VSUBS 0.00911f
C743 B.n561 VSUBS 0.00911f
C744 B.n562 VSUBS 0.00911f
C745 B.n563 VSUBS 0.00911f
C746 B.n564 VSUBS 0.00911f
C747 B.n565 VSUBS 0.00911f
C748 B.n566 VSUBS 0.00911f
C749 B.n567 VSUBS 0.00911f
C750 B.n568 VSUBS 0.00911f
C751 B.n569 VSUBS 0.00911f
C752 B.n570 VSUBS 0.00911f
C753 B.n571 VSUBS 0.00911f
C754 B.n572 VSUBS 0.00911f
C755 B.n573 VSUBS 0.00911f
C756 B.n574 VSUBS 0.00911f
C757 B.n575 VSUBS 0.00911f
C758 B.n576 VSUBS 0.00911f
C759 B.n577 VSUBS 0.00911f
C760 B.n578 VSUBS 0.00911f
C761 B.n579 VSUBS 0.00911f
C762 B.n580 VSUBS 0.00911f
C763 B.n581 VSUBS 0.00911f
C764 B.n582 VSUBS 0.00911f
C765 B.n583 VSUBS 0.00911f
C766 B.n584 VSUBS 0.00911f
C767 B.n585 VSUBS 0.00911f
C768 B.n586 VSUBS 0.00911f
C769 B.n587 VSUBS 0.00911f
C770 B.n588 VSUBS 0.00911f
C771 B.n589 VSUBS 0.00911f
C772 B.n590 VSUBS 0.00911f
C773 B.n591 VSUBS 0.00911f
C774 B.n592 VSUBS 0.00911f
C775 B.n593 VSUBS 0.00911f
C776 B.n594 VSUBS 0.00911f
C777 B.n595 VSUBS 0.00911f
C778 B.n596 VSUBS 0.00911f
C779 B.n597 VSUBS 0.00911f
C780 B.n598 VSUBS 0.00911f
C781 B.n599 VSUBS 0.00911f
C782 B.n600 VSUBS 0.00911f
C783 B.n601 VSUBS 0.00911f
C784 B.n602 VSUBS 0.00911f
C785 B.n603 VSUBS 0.00911f
C786 B.n604 VSUBS 0.00911f
C787 B.n605 VSUBS 0.00911f
C788 B.n606 VSUBS 0.00911f
C789 B.n607 VSUBS 0.00911f
C790 B.n608 VSUBS 0.00911f
C791 B.n609 VSUBS 0.00911f
C792 B.n610 VSUBS 0.00911f
C793 B.n611 VSUBS 0.00911f
C794 B.n612 VSUBS 0.00911f
C795 B.n613 VSUBS 0.00911f
C796 B.n614 VSUBS 0.00911f
C797 B.n615 VSUBS 0.00911f
C798 B.n616 VSUBS 0.00911f
C799 B.n617 VSUBS 0.00911f
C800 B.n618 VSUBS 0.00911f
C801 B.n619 VSUBS 0.00911f
C802 B.n620 VSUBS 0.00911f
C803 B.n621 VSUBS 0.00911f
C804 B.n622 VSUBS 0.00911f
C805 B.n623 VSUBS 0.00911f
C806 B.n624 VSUBS 0.00911f
C807 B.n625 VSUBS 0.00911f
C808 B.n626 VSUBS 0.00911f
C809 B.n627 VSUBS 0.00911f
C810 B.n628 VSUBS 0.00911f
C811 B.n629 VSUBS 0.00911f
C812 B.n630 VSUBS 0.00911f
C813 B.n631 VSUBS 0.00911f
C814 B.n632 VSUBS 0.00911f
C815 B.n633 VSUBS 0.00911f
C816 B.n634 VSUBS 0.00911f
C817 B.n635 VSUBS 0.00911f
C818 B.n636 VSUBS 0.00911f
C819 B.n637 VSUBS 0.00911f
C820 B.n638 VSUBS 0.00911f
C821 B.n639 VSUBS 0.00911f
C822 B.n640 VSUBS 0.00911f
C823 B.n641 VSUBS 0.00911f
C824 B.n642 VSUBS 0.00911f
C825 B.n643 VSUBS 0.00911f
C826 B.n644 VSUBS 0.00911f
C827 B.n645 VSUBS 0.00911f
C828 B.n646 VSUBS 0.00911f
C829 B.n647 VSUBS 0.00911f
C830 B.n648 VSUBS 0.00911f
C831 B.n649 VSUBS 0.00911f
C832 B.n650 VSUBS 0.00911f
C833 B.n651 VSUBS 0.00911f
C834 B.n652 VSUBS 0.00911f
C835 B.n653 VSUBS 0.00911f
C836 B.n654 VSUBS 0.00911f
C837 B.n655 VSUBS 0.00911f
C838 B.n656 VSUBS 0.00911f
C839 B.n657 VSUBS 0.00911f
C840 B.n658 VSUBS 0.00911f
C841 B.n659 VSUBS 0.00911f
C842 B.n660 VSUBS 0.00911f
C843 B.n661 VSUBS 0.00911f
C844 B.n662 VSUBS 0.00911f
C845 B.n663 VSUBS 0.00911f
C846 B.n664 VSUBS 0.00911f
C847 B.n665 VSUBS 0.00911f
C848 B.n666 VSUBS 0.00911f
C849 B.n667 VSUBS 0.00911f
C850 B.n668 VSUBS 0.00911f
C851 B.n669 VSUBS 0.00911f
C852 B.n670 VSUBS 0.00911f
C853 B.n671 VSUBS 0.00911f
C854 B.n672 VSUBS 0.00911f
C855 B.n673 VSUBS 0.00911f
C856 B.n674 VSUBS 0.00911f
C857 B.n675 VSUBS 0.00911f
C858 B.n676 VSUBS 0.00911f
C859 B.n677 VSUBS 0.00911f
C860 B.n678 VSUBS 0.00911f
C861 B.n679 VSUBS 0.00911f
C862 B.n680 VSUBS 0.00911f
C863 B.n681 VSUBS 0.00911f
C864 B.n682 VSUBS 0.00911f
C865 B.n683 VSUBS 0.00911f
C866 B.n684 VSUBS 0.00911f
C867 B.n685 VSUBS 0.00911f
C868 B.n686 VSUBS 0.00911f
C869 B.n687 VSUBS 0.00911f
C870 B.n688 VSUBS 0.00911f
C871 B.n689 VSUBS 0.00911f
C872 B.n690 VSUBS 0.00911f
C873 B.n691 VSUBS 0.00911f
C874 B.n692 VSUBS 0.00911f
C875 B.n693 VSUBS 0.00911f
C876 B.n694 VSUBS 0.00911f
C877 B.n695 VSUBS 0.00911f
C878 B.n696 VSUBS 0.00911f
C879 B.n697 VSUBS 0.00911f
C880 B.n698 VSUBS 0.00911f
C881 B.n699 VSUBS 0.00911f
C882 B.n700 VSUBS 0.00911f
C883 B.n701 VSUBS 0.00911f
C884 B.n702 VSUBS 0.00911f
C885 B.n703 VSUBS 0.00911f
C886 B.n704 VSUBS 0.00911f
C887 B.n705 VSUBS 0.00911f
C888 B.n706 VSUBS 0.00911f
C889 B.n707 VSUBS 0.00911f
C890 B.n708 VSUBS 0.00911f
C891 B.n709 VSUBS 0.00911f
C892 B.n710 VSUBS 0.00911f
C893 B.n711 VSUBS 0.00911f
C894 B.n712 VSUBS 0.00911f
C895 B.n713 VSUBS 0.00911f
C896 B.n714 VSUBS 0.00911f
C897 B.n715 VSUBS 0.00911f
C898 B.n716 VSUBS 0.00911f
C899 B.n717 VSUBS 0.00911f
C900 B.n718 VSUBS 0.00911f
C901 B.n719 VSUBS 0.00911f
C902 B.n720 VSUBS 0.00911f
C903 B.n721 VSUBS 0.00911f
C904 B.n722 VSUBS 0.00911f
C905 B.n723 VSUBS 0.00911f
C906 B.n724 VSUBS 0.00911f
C907 B.n725 VSUBS 0.00911f
C908 B.n726 VSUBS 0.00911f
C909 B.n727 VSUBS 0.00911f
C910 B.n728 VSUBS 0.00911f
C911 B.n729 VSUBS 0.00911f
C912 B.n730 VSUBS 0.00911f
C913 B.n731 VSUBS 0.00911f
C914 B.n732 VSUBS 0.00911f
C915 B.n733 VSUBS 0.00911f
C916 B.n734 VSUBS 0.00911f
C917 B.n735 VSUBS 0.00911f
C918 B.n736 VSUBS 0.00911f
C919 B.n737 VSUBS 0.00911f
C920 B.n738 VSUBS 0.00911f
C921 B.n739 VSUBS 0.00911f
C922 B.n740 VSUBS 0.00911f
C923 B.n741 VSUBS 0.00911f
C924 B.n742 VSUBS 0.00911f
C925 B.n743 VSUBS 0.00911f
C926 B.n744 VSUBS 0.00911f
C927 B.n745 VSUBS 0.00911f
C928 B.n746 VSUBS 0.00911f
C929 B.n747 VSUBS 0.00911f
C930 B.n748 VSUBS 0.00911f
C931 B.n749 VSUBS 0.00911f
C932 B.n750 VSUBS 0.00911f
C933 B.n751 VSUBS 0.00911f
C934 B.n752 VSUBS 0.00911f
C935 B.n753 VSUBS 0.00911f
C936 B.n754 VSUBS 0.00911f
C937 B.n755 VSUBS 0.00911f
C938 B.n756 VSUBS 0.00911f
C939 B.n757 VSUBS 0.00911f
C940 B.n758 VSUBS 0.00911f
C941 B.n759 VSUBS 0.00911f
C942 B.n760 VSUBS 0.00911f
C943 B.n761 VSUBS 0.00911f
C944 B.n762 VSUBS 0.00911f
C945 B.n763 VSUBS 0.00911f
C946 B.n764 VSUBS 0.00911f
C947 B.n765 VSUBS 0.00911f
C948 B.n766 VSUBS 0.00911f
C949 B.n767 VSUBS 0.00911f
C950 B.n768 VSUBS 0.00911f
C951 B.n769 VSUBS 0.00911f
C952 B.n770 VSUBS 0.020048f
C953 B.n771 VSUBS 0.021753f
C954 B.n772 VSUBS 0.021753f
C955 B.n773 VSUBS 0.00911f
C956 B.n774 VSUBS 0.00911f
C957 B.n775 VSUBS 0.00911f
C958 B.n776 VSUBS 0.00911f
C959 B.n777 VSUBS 0.00911f
C960 B.n778 VSUBS 0.00911f
C961 B.n779 VSUBS 0.00911f
C962 B.n780 VSUBS 0.00911f
C963 B.n781 VSUBS 0.00911f
C964 B.n782 VSUBS 0.00911f
C965 B.n783 VSUBS 0.00911f
C966 B.n784 VSUBS 0.00911f
C967 B.n785 VSUBS 0.00911f
C968 B.n786 VSUBS 0.00911f
C969 B.n787 VSUBS 0.00911f
C970 B.n788 VSUBS 0.00911f
C971 B.n789 VSUBS 0.00911f
C972 B.n790 VSUBS 0.00911f
C973 B.n791 VSUBS 0.00911f
C974 B.n792 VSUBS 0.00911f
C975 B.n793 VSUBS 0.00911f
C976 B.n794 VSUBS 0.00911f
C977 B.n795 VSUBS 0.00911f
C978 B.n796 VSUBS 0.00911f
C979 B.n797 VSUBS 0.00911f
C980 B.n798 VSUBS 0.00911f
C981 B.n799 VSUBS 0.00911f
C982 B.n800 VSUBS 0.00911f
C983 B.n801 VSUBS 0.00911f
C984 B.n802 VSUBS 0.00911f
C985 B.n803 VSUBS 0.00911f
C986 B.n804 VSUBS 0.00911f
C987 B.n805 VSUBS 0.00911f
C988 B.n806 VSUBS 0.00911f
C989 B.n807 VSUBS 0.00911f
C990 B.n808 VSUBS 0.00911f
C991 B.n809 VSUBS 0.00911f
C992 B.n810 VSUBS 0.00911f
C993 B.n811 VSUBS 0.00911f
C994 B.n812 VSUBS 0.00911f
C995 B.n813 VSUBS 0.00911f
C996 B.n814 VSUBS 0.00911f
C997 B.n815 VSUBS 0.00911f
C998 B.n816 VSUBS 0.00911f
C999 B.n817 VSUBS 0.00911f
C1000 B.n818 VSUBS 0.00911f
C1001 B.n819 VSUBS 0.00911f
C1002 B.n820 VSUBS 0.00911f
C1003 B.n821 VSUBS 0.00911f
C1004 B.n822 VSUBS 0.00911f
C1005 B.n823 VSUBS 0.00911f
C1006 B.n824 VSUBS 0.00911f
C1007 B.n825 VSUBS 0.00911f
C1008 B.n826 VSUBS 0.00911f
C1009 B.n827 VSUBS 0.00911f
C1010 B.n828 VSUBS 0.00911f
C1011 B.n829 VSUBS 0.006297f
C1012 B.n830 VSUBS 0.021108f
C1013 B.n831 VSUBS 0.007369f
C1014 B.n832 VSUBS 0.00911f
C1015 B.n833 VSUBS 0.00911f
C1016 B.n834 VSUBS 0.00911f
C1017 B.n835 VSUBS 0.00911f
C1018 B.n836 VSUBS 0.00911f
C1019 B.n837 VSUBS 0.00911f
C1020 B.n838 VSUBS 0.00911f
C1021 B.n839 VSUBS 0.00911f
C1022 B.n840 VSUBS 0.00911f
C1023 B.n841 VSUBS 0.00911f
C1024 B.n842 VSUBS 0.00911f
C1025 B.n843 VSUBS 0.007369f
C1026 B.n844 VSUBS 0.021108f
C1027 B.n845 VSUBS 0.006297f
C1028 B.n846 VSUBS 0.00911f
C1029 B.n847 VSUBS 0.00911f
C1030 B.n848 VSUBS 0.00911f
C1031 B.n849 VSUBS 0.00911f
C1032 B.n850 VSUBS 0.00911f
C1033 B.n851 VSUBS 0.00911f
C1034 B.n852 VSUBS 0.00911f
C1035 B.n853 VSUBS 0.00911f
C1036 B.n854 VSUBS 0.00911f
C1037 B.n855 VSUBS 0.00911f
C1038 B.n856 VSUBS 0.00911f
C1039 B.n857 VSUBS 0.00911f
C1040 B.n858 VSUBS 0.00911f
C1041 B.n859 VSUBS 0.00911f
C1042 B.n860 VSUBS 0.00911f
C1043 B.n861 VSUBS 0.00911f
C1044 B.n862 VSUBS 0.00911f
C1045 B.n863 VSUBS 0.00911f
C1046 B.n864 VSUBS 0.00911f
C1047 B.n865 VSUBS 0.00911f
C1048 B.n866 VSUBS 0.00911f
C1049 B.n867 VSUBS 0.00911f
C1050 B.n868 VSUBS 0.00911f
C1051 B.n869 VSUBS 0.00911f
C1052 B.n870 VSUBS 0.00911f
C1053 B.n871 VSUBS 0.00911f
C1054 B.n872 VSUBS 0.00911f
C1055 B.n873 VSUBS 0.00911f
C1056 B.n874 VSUBS 0.00911f
C1057 B.n875 VSUBS 0.00911f
C1058 B.n876 VSUBS 0.00911f
C1059 B.n877 VSUBS 0.00911f
C1060 B.n878 VSUBS 0.00911f
C1061 B.n879 VSUBS 0.00911f
C1062 B.n880 VSUBS 0.00911f
C1063 B.n881 VSUBS 0.00911f
C1064 B.n882 VSUBS 0.00911f
C1065 B.n883 VSUBS 0.00911f
C1066 B.n884 VSUBS 0.00911f
C1067 B.n885 VSUBS 0.00911f
C1068 B.n886 VSUBS 0.00911f
C1069 B.n887 VSUBS 0.00911f
C1070 B.n888 VSUBS 0.00911f
C1071 B.n889 VSUBS 0.00911f
C1072 B.n890 VSUBS 0.00911f
C1073 B.n891 VSUBS 0.00911f
C1074 B.n892 VSUBS 0.00911f
C1075 B.n893 VSUBS 0.00911f
C1076 B.n894 VSUBS 0.00911f
C1077 B.n895 VSUBS 0.00911f
C1078 B.n896 VSUBS 0.00911f
C1079 B.n897 VSUBS 0.00911f
C1080 B.n898 VSUBS 0.00911f
C1081 B.n899 VSUBS 0.00911f
C1082 B.n900 VSUBS 0.00911f
C1083 B.n901 VSUBS 0.00911f
C1084 B.n902 VSUBS 0.021753f
C1085 B.n903 VSUBS 0.021753f
C1086 B.n904 VSUBS 0.020048f
C1087 B.n905 VSUBS 0.00911f
C1088 B.n906 VSUBS 0.00911f
C1089 B.n907 VSUBS 0.00911f
C1090 B.n908 VSUBS 0.00911f
C1091 B.n909 VSUBS 0.00911f
C1092 B.n910 VSUBS 0.00911f
C1093 B.n911 VSUBS 0.00911f
C1094 B.n912 VSUBS 0.00911f
C1095 B.n913 VSUBS 0.00911f
C1096 B.n914 VSUBS 0.00911f
C1097 B.n915 VSUBS 0.00911f
C1098 B.n916 VSUBS 0.00911f
C1099 B.n917 VSUBS 0.00911f
C1100 B.n918 VSUBS 0.00911f
C1101 B.n919 VSUBS 0.00911f
C1102 B.n920 VSUBS 0.00911f
C1103 B.n921 VSUBS 0.00911f
C1104 B.n922 VSUBS 0.00911f
C1105 B.n923 VSUBS 0.00911f
C1106 B.n924 VSUBS 0.00911f
C1107 B.n925 VSUBS 0.00911f
C1108 B.n926 VSUBS 0.00911f
C1109 B.n927 VSUBS 0.00911f
C1110 B.n928 VSUBS 0.00911f
C1111 B.n929 VSUBS 0.00911f
C1112 B.n930 VSUBS 0.00911f
C1113 B.n931 VSUBS 0.00911f
C1114 B.n932 VSUBS 0.00911f
C1115 B.n933 VSUBS 0.00911f
C1116 B.n934 VSUBS 0.00911f
C1117 B.n935 VSUBS 0.00911f
C1118 B.n936 VSUBS 0.00911f
C1119 B.n937 VSUBS 0.00911f
C1120 B.n938 VSUBS 0.00911f
C1121 B.n939 VSUBS 0.00911f
C1122 B.n940 VSUBS 0.00911f
C1123 B.n941 VSUBS 0.00911f
C1124 B.n942 VSUBS 0.00911f
C1125 B.n943 VSUBS 0.00911f
C1126 B.n944 VSUBS 0.00911f
C1127 B.n945 VSUBS 0.00911f
C1128 B.n946 VSUBS 0.00911f
C1129 B.n947 VSUBS 0.00911f
C1130 B.n948 VSUBS 0.00911f
C1131 B.n949 VSUBS 0.00911f
C1132 B.n950 VSUBS 0.00911f
C1133 B.n951 VSUBS 0.00911f
C1134 B.n952 VSUBS 0.00911f
C1135 B.n953 VSUBS 0.00911f
C1136 B.n954 VSUBS 0.00911f
C1137 B.n955 VSUBS 0.00911f
C1138 B.n956 VSUBS 0.00911f
C1139 B.n957 VSUBS 0.00911f
C1140 B.n958 VSUBS 0.00911f
C1141 B.n959 VSUBS 0.00911f
C1142 B.n960 VSUBS 0.00911f
C1143 B.n961 VSUBS 0.00911f
C1144 B.n962 VSUBS 0.00911f
C1145 B.n963 VSUBS 0.00911f
C1146 B.n964 VSUBS 0.00911f
C1147 B.n965 VSUBS 0.00911f
C1148 B.n966 VSUBS 0.00911f
C1149 B.n967 VSUBS 0.00911f
C1150 B.n968 VSUBS 0.00911f
C1151 B.n969 VSUBS 0.00911f
C1152 B.n970 VSUBS 0.00911f
C1153 B.n971 VSUBS 0.00911f
C1154 B.n972 VSUBS 0.00911f
C1155 B.n973 VSUBS 0.00911f
C1156 B.n974 VSUBS 0.00911f
C1157 B.n975 VSUBS 0.00911f
C1158 B.n976 VSUBS 0.00911f
C1159 B.n977 VSUBS 0.00911f
C1160 B.n978 VSUBS 0.00911f
C1161 B.n979 VSUBS 0.00911f
C1162 B.n980 VSUBS 0.00911f
C1163 B.n981 VSUBS 0.00911f
C1164 B.n982 VSUBS 0.00911f
C1165 B.n983 VSUBS 0.00911f
C1166 B.n984 VSUBS 0.00911f
C1167 B.n985 VSUBS 0.00911f
C1168 B.n986 VSUBS 0.00911f
C1169 B.n987 VSUBS 0.00911f
C1170 B.n988 VSUBS 0.00911f
C1171 B.n989 VSUBS 0.00911f
C1172 B.n990 VSUBS 0.00911f
C1173 B.n991 VSUBS 0.00911f
C1174 B.n992 VSUBS 0.00911f
C1175 B.n993 VSUBS 0.00911f
C1176 B.n994 VSUBS 0.00911f
C1177 B.n995 VSUBS 0.00911f
C1178 B.n996 VSUBS 0.00911f
C1179 B.n997 VSUBS 0.00911f
C1180 B.n998 VSUBS 0.00911f
C1181 B.n999 VSUBS 0.00911f
C1182 B.n1000 VSUBS 0.00911f
C1183 B.n1001 VSUBS 0.00911f
C1184 B.n1002 VSUBS 0.00911f
C1185 B.n1003 VSUBS 0.00911f
C1186 B.n1004 VSUBS 0.00911f
C1187 B.n1005 VSUBS 0.00911f
C1188 B.n1006 VSUBS 0.00911f
C1189 B.n1007 VSUBS 0.00911f
C1190 B.n1008 VSUBS 0.00911f
C1191 B.n1009 VSUBS 0.00911f
C1192 B.n1010 VSUBS 0.00911f
C1193 B.n1011 VSUBS 0.00911f
C1194 B.n1012 VSUBS 0.00911f
C1195 B.n1013 VSUBS 0.00911f
C1196 B.n1014 VSUBS 0.00911f
C1197 B.n1015 VSUBS 0.00911f
C1198 B.n1016 VSUBS 0.00911f
C1199 B.n1017 VSUBS 0.00911f
C1200 B.n1018 VSUBS 0.00911f
C1201 B.n1019 VSUBS 0.00911f
C1202 B.n1020 VSUBS 0.00911f
C1203 B.n1021 VSUBS 0.00911f
C1204 B.n1022 VSUBS 0.00911f
C1205 B.n1023 VSUBS 0.00911f
C1206 B.n1024 VSUBS 0.00911f
C1207 B.n1025 VSUBS 0.00911f
C1208 B.n1026 VSUBS 0.00911f
C1209 B.n1027 VSUBS 0.011889f
C1210 B.n1028 VSUBS 0.012664f
C1211 B.n1029 VSUBS 0.025184f
C1212 VTAIL.t2 VSUBS 0.265769f
C1213 VTAIL.t0 VSUBS 0.265769f
C1214 VTAIL.n0 VSUBS 1.86456f
C1215 VTAIL.n1 VSUBS 1.20988f
C1216 VTAIL.t8 VSUBS 2.47365f
C1217 VTAIL.n2 VSUBS 1.41122f
C1218 VTAIL.t14 VSUBS 0.265769f
C1219 VTAIL.t15 VSUBS 0.265769f
C1220 VTAIL.n3 VSUBS 1.86456f
C1221 VTAIL.n4 VSUBS 1.43169f
C1222 VTAIL.t10 VSUBS 0.265769f
C1223 VTAIL.t11 VSUBS 0.265769f
C1224 VTAIL.n5 VSUBS 1.86456f
C1225 VTAIL.n6 VSUBS 3.14899f
C1226 VTAIL.t7 VSUBS 0.265769f
C1227 VTAIL.t1 VSUBS 0.265769f
C1228 VTAIL.n7 VSUBS 1.86457f
C1229 VTAIL.n8 VSUBS 3.14898f
C1230 VTAIL.t19 VSUBS 0.265769f
C1231 VTAIL.t5 VSUBS 0.265769f
C1232 VTAIL.n9 VSUBS 1.86457f
C1233 VTAIL.n10 VSUBS 1.43168f
C1234 VTAIL.t6 VSUBS 2.47367f
C1235 VTAIL.n11 VSUBS 1.4112f
C1236 VTAIL.t16 VSUBS 0.265769f
C1237 VTAIL.t12 VSUBS 0.265769f
C1238 VTAIL.n12 VSUBS 1.86457f
C1239 VTAIL.n13 VSUBS 1.29548f
C1240 VTAIL.t9 VSUBS 0.265769f
C1241 VTAIL.t17 VSUBS 0.265769f
C1242 VTAIL.n14 VSUBS 1.86457f
C1243 VTAIL.n15 VSUBS 1.43168f
C1244 VTAIL.t13 VSUBS 2.47365f
C1245 VTAIL.n16 VSUBS 2.89923f
C1246 VTAIL.t18 VSUBS 2.47365f
C1247 VTAIL.n17 VSUBS 2.89923f
C1248 VTAIL.t3 VSUBS 0.265769f
C1249 VTAIL.t4 VSUBS 0.265769f
C1250 VTAIL.n18 VSUBS 1.86456f
C1251 VTAIL.n19 VSUBS 1.15181f
C1252 VDD1.t7 VSUBS 2.81455f
C1253 VDD1.t9 VSUBS 0.276195f
C1254 VDD1.t6 VSUBS 0.276195f
C1255 VDD1.n0 VSUBS 2.11175f
C1256 VDD1.n1 VSUBS 2.11908f
C1257 VDD1.t3 VSUBS 2.81454f
C1258 VDD1.t0 VSUBS 0.276195f
C1259 VDD1.t4 VSUBS 0.276195f
C1260 VDD1.n2 VSUBS 2.11174f
C1261 VDD1.n3 VSUBS 2.10827f
C1262 VDD1.t8 VSUBS 0.276195f
C1263 VDD1.t5 VSUBS 0.276195f
C1264 VDD1.n4 VSUBS 2.15701f
C1265 VDD1.n5 VSUBS 5.05944f
C1266 VDD1.t2 VSUBS 0.276195f
C1267 VDD1.t1 VSUBS 0.276195f
C1268 VDD1.n6 VSUBS 2.11174f
C1269 VDD1.n7 VSUBS 5.00249f
C1270 VP.t9 VSUBS 3.03161f
C1271 VP.n0 VSUBS 1.16584f
C1272 VP.n1 VSUBS 0.02582f
C1273 VP.n2 VSUBS 0.051794f
C1274 VP.n3 VSUBS 0.02582f
C1275 VP.n4 VSUBS 0.047881f
C1276 VP.n5 VSUBS 0.02582f
C1277 VP.t2 VSUBS 3.03161f
C1278 VP.n6 VSUBS 0.047881f
C1279 VP.n7 VSUBS 0.02582f
C1280 VP.n8 VSUBS 0.047881f
C1281 VP.n9 VSUBS 0.02582f
C1282 VP.t3 VSUBS 3.03161f
C1283 VP.n10 VSUBS 0.047881f
C1284 VP.n11 VSUBS 0.02582f
C1285 VP.n12 VSUBS 0.047881f
C1286 VP.n13 VSUBS 0.02582f
C1287 VP.t6 VSUBS 3.03161f
C1288 VP.n14 VSUBS 0.047881f
C1289 VP.n15 VSUBS 0.02582f
C1290 VP.n16 VSUBS 0.051794f
C1291 VP.n17 VSUBS 0.02582f
C1292 VP.t7 VSUBS 3.03161f
C1293 VP.n18 VSUBS 1.16584f
C1294 VP.t4 VSUBS 3.03161f
C1295 VP.n19 VSUBS 1.16584f
C1296 VP.n20 VSUBS 0.02582f
C1297 VP.n21 VSUBS 0.051794f
C1298 VP.n22 VSUBS 0.02582f
C1299 VP.n23 VSUBS 0.047881f
C1300 VP.n24 VSUBS 0.02582f
C1301 VP.t0 VSUBS 3.03161f
C1302 VP.n25 VSUBS 0.047881f
C1303 VP.n26 VSUBS 0.02582f
C1304 VP.n27 VSUBS 0.047881f
C1305 VP.n28 VSUBS 0.02582f
C1306 VP.t8 VSUBS 3.03161f
C1307 VP.n29 VSUBS 0.047881f
C1308 VP.n30 VSUBS 0.02582f
C1309 VP.n31 VSUBS 0.047881f
C1310 VP.n32 VSUBS 0.336422f
C1311 VP.t5 VSUBS 3.03161f
C1312 VP.t1 VSUBS 3.45254f
C1313 VP.n33 VSUBS 1.10248f
C1314 VP.n34 VSUBS 1.16072f
C1315 VP.n35 VSUBS 0.03748f
C1316 VP.n36 VSUBS 0.047881f
C1317 VP.n37 VSUBS 0.02582f
C1318 VP.n38 VSUBS 0.02582f
C1319 VP.n39 VSUBS 0.02582f
C1320 VP.n40 VSUBS 0.045043f
C1321 VP.n41 VSUBS 0.028117f
C1322 VP.n42 VSUBS 0.049788f
C1323 VP.n43 VSUBS 0.02582f
C1324 VP.n44 VSUBS 0.02582f
C1325 VP.n45 VSUBS 0.02582f
C1326 VP.n46 VSUBS 0.047881f
C1327 VP.n47 VSUBS 1.09018f
C1328 VP.n48 VSUBS 0.047881f
C1329 VP.n49 VSUBS 0.02582f
C1330 VP.n50 VSUBS 0.02582f
C1331 VP.n51 VSUBS 0.02582f
C1332 VP.n52 VSUBS 0.049788f
C1333 VP.n53 VSUBS 0.028117f
C1334 VP.n54 VSUBS 0.045043f
C1335 VP.n55 VSUBS 0.02582f
C1336 VP.n56 VSUBS 0.02582f
C1337 VP.n57 VSUBS 0.02582f
C1338 VP.n58 VSUBS 0.047881f
C1339 VP.n59 VSUBS 0.03748f
C1340 VP.n60 VSUBS 1.06593f
C1341 VP.n61 VSUBS 0.034644f
C1342 VP.n62 VSUBS 0.02582f
C1343 VP.n63 VSUBS 0.02582f
C1344 VP.n64 VSUBS 0.02582f
C1345 VP.n65 VSUBS 0.047881f
C1346 VP.n66 VSUBS 0.048113f
C1347 VP.n67 VSUBS 0.02304f
C1348 VP.n68 VSUBS 0.02582f
C1349 VP.n69 VSUBS 0.02582f
C1350 VP.n70 VSUBS 0.02582f
C1351 VP.n71 VSUBS 0.047881f
C1352 VP.n72 VSUBS 0.047881f
C1353 VP.n73 VSUBS 0.02708f
C1354 VP.n74 VSUBS 0.041666f
C1355 VP.n75 VSUBS 1.9002f
C1356 VP.n76 VSUBS 1.91578f
C1357 VP.n77 VSUBS 0.041666f
C1358 VP.n78 VSUBS 0.02708f
C1359 VP.n79 VSUBS 0.047881f
C1360 VP.n80 VSUBS 0.047881f
C1361 VP.n81 VSUBS 0.02582f
C1362 VP.n82 VSUBS 0.02582f
C1363 VP.n83 VSUBS 0.02582f
C1364 VP.n84 VSUBS 0.02304f
C1365 VP.n85 VSUBS 0.048113f
C1366 VP.n86 VSUBS 0.047881f
C1367 VP.n87 VSUBS 0.02582f
C1368 VP.n88 VSUBS 0.02582f
C1369 VP.n89 VSUBS 0.02582f
C1370 VP.n90 VSUBS 0.034644f
C1371 VP.n91 VSUBS 1.06593f
C1372 VP.n92 VSUBS 0.03748f
C1373 VP.n93 VSUBS 0.047881f
C1374 VP.n94 VSUBS 0.02582f
C1375 VP.n95 VSUBS 0.02582f
C1376 VP.n96 VSUBS 0.02582f
C1377 VP.n97 VSUBS 0.045043f
C1378 VP.n98 VSUBS 0.028117f
C1379 VP.n99 VSUBS 0.049788f
C1380 VP.n100 VSUBS 0.02582f
C1381 VP.n101 VSUBS 0.02582f
C1382 VP.n102 VSUBS 0.02582f
C1383 VP.n103 VSUBS 0.047881f
C1384 VP.n104 VSUBS 1.09018f
C1385 VP.n105 VSUBS 0.047881f
C1386 VP.n106 VSUBS 0.02582f
C1387 VP.n107 VSUBS 0.02582f
C1388 VP.n108 VSUBS 0.02582f
C1389 VP.n109 VSUBS 0.049788f
C1390 VP.n110 VSUBS 0.028117f
C1391 VP.n111 VSUBS 0.045043f
C1392 VP.n112 VSUBS 0.02582f
C1393 VP.n113 VSUBS 0.02582f
C1394 VP.n114 VSUBS 0.02582f
C1395 VP.n115 VSUBS 0.047881f
C1396 VP.n116 VSUBS 0.03748f
C1397 VP.n117 VSUBS 1.06593f
C1398 VP.n118 VSUBS 0.034644f
C1399 VP.n119 VSUBS 0.02582f
C1400 VP.n120 VSUBS 0.02582f
C1401 VP.n121 VSUBS 0.02582f
C1402 VP.n122 VSUBS 0.047881f
C1403 VP.n123 VSUBS 0.048113f
C1404 VP.n124 VSUBS 0.02304f
C1405 VP.n125 VSUBS 0.02582f
C1406 VP.n126 VSUBS 0.02582f
C1407 VP.n127 VSUBS 0.02582f
C1408 VP.n128 VSUBS 0.047881f
C1409 VP.n129 VSUBS 0.047881f
C1410 VP.n130 VSUBS 0.02708f
C1411 VP.n131 VSUBS 0.041666f
C1412 VP.n132 VSUBS 0.081319f
.ends

