* NGSPICE file created from diff_pair_sample_0264.ext - technology: sky130A

.subckt diff_pair_sample_0264 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.53
X1 VDD2.t4 VN.t1 VTAIL.t7 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.53
X2 B.t11 B.t9 B.t10 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.53
X3 VDD1.t5 VP.t0 VTAIL.t1 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.53
X4 VDD1.t4 VP.t1 VTAIL.t2 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.53
X5 VTAIL.t6 VN.t2 VDD2.t3 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.53
X6 B.t8 B.t6 B.t7 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.53
X7 VTAIL.t3 VP.t2 VDD1.t3 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.53
X8 VDD2.t2 VN.t3 VTAIL.t11 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.53
X9 B.t5 B.t3 B.t4 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.53
X10 VDD1.t2 VP.t3 VTAIL.t0 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.53
X11 VDD2.t1 VN.t4 VTAIL.t8 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.53
X12 B.t2 B.t0 B.t1 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.53
X13 VTAIL.t10 VN.t5 VDD2.t0 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.53
X14 VTAIL.t4 VP.t4 VDD1.t1 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.53
X15 VDD1.t0 VP.t5 VTAIL.t5 w_n2458_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.53
R0 VN.n11 VN.n10 180.385
R1 VN.n23 VN.n22 180.385
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n8 VN.n1 56.5193
R11 VN.n20 VN.n13 56.5193
R12 VN.n3 VN.n2 53.6827
R13 VN.n15 VN.n14 53.6827
R14 VN.n2 VN.t1 44.6322
R15 VN.n14 VN.t3 44.6322
R16 VN VN.n23 36.2751
R17 VN.n4 VN.n1 24.4675
R18 VN.n9 VN.n8 24.4675
R19 VN.n16 VN.n13 24.4675
R20 VN.n21 VN.n20 24.4675
R21 VN.n17 VN.n14 18.2406
R22 VN.n5 VN.n2 18.2406
R23 VN.n3 VN.t5 13.3894
R24 VN.n10 VN.t4 13.3894
R25 VN.n15 VN.t2 13.3894
R26 VN.n22 VN.t0 13.3894
R27 VN.n4 VN.n3 12.234
R28 VN.n16 VN.n15 12.234
R29 VN.n10 VN.n9 5.38324
R30 VN.n22 VN.n21 5.38324
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n10 VTAIL.t5 658.787
R41 VTAIL.n7 VTAIL.t11 658.787
R42 VTAIL.n11 VTAIL.t8 658.785
R43 VTAIL.n2 VTAIL.t1 658.785
R44 VTAIL.n9 VTAIL.n8 620.544
R45 VTAIL.n6 VTAIL.n5 620.544
R46 VTAIL.n1 VTAIL.n0 620.544
R47 VTAIL.n4 VTAIL.n3 620.544
R48 VTAIL.n0 VTAIL.t7 38.2417
R49 VTAIL.n0 VTAIL.t10 38.2417
R50 VTAIL.n3 VTAIL.t2 38.2417
R51 VTAIL.n3 VTAIL.t4 38.2417
R52 VTAIL.n8 VTAIL.t0 38.2417
R53 VTAIL.n8 VTAIL.t3 38.2417
R54 VTAIL.n5 VTAIL.t9 38.2417
R55 VTAIL.n5 VTAIL.t6 38.2417
R56 VTAIL.n6 VTAIL.n4 16.3065
R57 VTAIL.n11 VTAIL.n10 14.7031
R58 VTAIL.n7 VTAIL.n6 1.60395
R59 VTAIL.n10 VTAIL.n9 1.60395
R60 VTAIL.n4 VTAIL.n2 1.60395
R61 VTAIL.n9 VTAIL.n7 1.27205
R62 VTAIL.n2 VTAIL.n1 1.27205
R63 VTAIL VTAIL.n11 1.1449
R64 VTAIL VTAIL.n1 0.459552
R65 VDD2.n1 VDD2.t4 676.611
R66 VDD2.n2 VDD2.t5 675.465
R67 VDD2.n1 VDD2.n0 637.568
R68 VDD2 VDD2.n3 637.567
R69 VDD2.n3 VDD2.t3 38.2417
R70 VDD2.n3 VDD2.t2 38.2417
R71 VDD2.n0 VDD2.t0 38.2417
R72 VDD2.n0 VDD2.t1 38.2417
R73 VDD2.n2 VDD2.n1 29.6593
R74 VDD2 VDD2.n2 1.26128
R75 B.n70 B.t11 685.496
R76 B.n78 B.t2 685.496
R77 B.n22 B.t4 685.496
R78 B.n28 B.t7 685.496
R79 B.n71 B.t10 649.423
R80 B.n79 B.t1 649.423
R81 B.n23 B.t5 649.423
R82 B.n29 B.t8 649.423
R83 B.n276 B.n275 585
R84 B.n277 B.n34 585
R85 B.n279 B.n278 585
R86 B.n280 B.n33 585
R87 B.n282 B.n281 585
R88 B.n283 B.n32 585
R89 B.n285 B.n284 585
R90 B.n286 B.n31 585
R91 B.n288 B.n287 585
R92 B.n290 B.n289 585
R93 B.n291 B.n27 585
R94 B.n293 B.n292 585
R95 B.n294 B.n26 585
R96 B.n296 B.n295 585
R97 B.n297 B.n25 585
R98 B.n299 B.n298 585
R99 B.n300 B.n24 585
R100 B.n302 B.n301 585
R101 B.n304 B.n21 585
R102 B.n306 B.n305 585
R103 B.n307 B.n20 585
R104 B.n309 B.n308 585
R105 B.n310 B.n19 585
R106 B.n312 B.n311 585
R107 B.n313 B.n18 585
R108 B.n315 B.n314 585
R109 B.n316 B.n17 585
R110 B.n274 B.n35 585
R111 B.n273 B.n272 585
R112 B.n271 B.n36 585
R113 B.n270 B.n269 585
R114 B.n268 B.n37 585
R115 B.n267 B.n266 585
R116 B.n265 B.n38 585
R117 B.n264 B.n263 585
R118 B.n262 B.n39 585
R119 B.n261 B.n260 585
R120 B.n259 B.n40 585
R121 B.n258 B.n257 585
R122 B.n256 B.n41 585
R123 B.n255 B.n254 585
R124 B.n253 B.n42 585
R125 B.n252 B.n251 585
R126 B.n250 B.n43 585
R127 B.n249 B.n248 585
R128 B.n247 B.n44 585
R129 B.n246 B.n245 585
R130 B.n244 B.n45 585
R131 B.n243 B.n242 585
R132 B.n241 B.n46 585
R133 B.n240 B.n239 585
R134 B.n238 B.n47 585
R135 B.n237 B.n236 585
R136 B.n235 B.n48 585
R137 B.n234 B.n233 585
R138 B.n232 B.n49 585
R139 B.n231 B.n230 585
R140 B.n229 B.n50 585
R141 B.n228 B.n227 585
R142 B.n226 B.n51 585
R143 B.n225 B.n224 585
R144 B.n223 B.n52 585
R145 B.n222 B.n221 585
R146 B.n220 B.n53 585
R147 B.n219 B.n218 585
R148 B.n217 B.n54 585
R149 B.n216 B.n215 585
R150 B.n214 B.n55 585
R151 B.n213 B.n212 585
R152 B.n211 B.n56 585
R153 B.n210 B.n209 585
R154 B.n208 B.n57 585
R155 B.n207 B.n206 585
R156 B.n205 B.n58 585
R157 B.n204 B.n203 585
R158 B.n202 B.n59 585
R159 B.n201 B.n200 585
R160 B.n199 B.n60 585
R161 B.n198 B.n197 585
R162 B.n196 B.n61 585
R163 B.n195 B.n194 585
R164 B.n193 B.n62 585
R165 B.n192 B.n191 585
R166 B.n190 B.n63 585
R167 B.n189 B.n188 585
R168 B.n187 B.n64 585
R169 B.n186 B.n185 585
R170 B.n184 B.n65 585
R171 B.n142 B.n83 585
R172 B.n144 B.n143 585
R173 B.n145 B.n82 585
R174 B.n147 B.n146 585
R175 B.n148 B.n81 585
R176 B.n150 B.n149 585
R177 B.n151 B.n80 585
R178 B.n153 B.n152 585
R179 B.n154 B.n77 585
R180 B.n157 B.n156 585
R181 B.n158 B.n76 585
R182 B.n160 B.n159 585
R183 B.n161 B.n75 585
R184 B.n163 B.n162 585
R185 B.n164 B.n74 585
R186 B.n166 B.n165 585
R187 B.n167 B.n73 585
R188 B.n169 B.n168 585
R189 B.n171 B.n170 585
R190 B.n172 B.n69 585
R191 B.n174 B.n173 585
R192 B.n175 B.n68 585
R193 B.n177 B.n176 585
R194 B.n178 B.n67 585
R195 B.n180 B.n179 585
R196 B.n181 B.n66 585
R197 B.n183 B.n182 585
R198 B.n141 B.n140 585
R199 B.n139 B.n84 585
R200 B.n138 B.n137 585
R201 B.n136 B.n85 585
R202 B.n135 B.n134 585
R203 B.n133 B.n86 585
R204 B.n132 B.n131 585
R205 B.n130 B.n87 585
R206 B.n129 B.n128 585
R207 B.n127 B.n88 585
R208 B.n126 B.n125 585
R209 B.n124 B.n89 585
R210 B.n123 B.n122 585
R211 B.n121 B.n90 585
R212 B.n120 B.n119 585
R213 B.n118 B.n91 585
R214 B.n117 B.n116 585
R215 B.n115 B.n92 585
R216 B.n114 B.n113 585
R217 B.n112 B.n93 585
R218 B.n111 B.n110 585
R219 B.n109 B.n94 585
R220 B.n108 B.n107 585
R221 B.n106 B.n95 585
R222 B.n105 B.n104 585
R223 B.n103 B.n96 585
R224 B.n102 B.n101 585
R225 B.n100 B.n97 585
R226 B.n99 B.n98 585
R227 B.n2 B.n0 585
R228 B.n361 B.n1 585
R229 B.n360 B.n359 585
R230 B.n358 B.n3 585
R231 B.n357 B.n356 585
R232 B.n355 B.n4 585
R233 B.n354 B.n353 585
R234 B.n352 B.n5 585
R235 B.n351 B.n350 585
R236 B.n349 B.n6 585
R237 B.n348 B.n347 585
R238 B.n346 B.n7 585
R239 B.n345 B.n344 585
R240 B.n343 B.n8 585
R241 B.n342 B.n341 585
R242 B.n340 B.n9 585
R243 B.n339 B.n338 585
R244 B.n337 B.n10 585
R245 B.n336 B.n335 585
R246 B.n334 B.n11 585
R247 B.n333 B.n332 585
R248 B.n331 B.n12 585
R249 B.n330 B.n329 585
R250 B.n328 B.n13 585
R251 B.n327 B.n326 585
R252 B.n325 B.n14 585
R253 B.n324 B.n323 585
R254 B.n322 B.n15 585
R255 B.n321 B.n320 585
R256 B.n319 B.n16 585
R257 B.n318 B.n317 585
R258 B.n363 B.n362 585
R259 B.n140 B.n83 516.524
R260 B.n318 B.n17 516.524
R261 B.n182 B.n65 516.524
R262 B.n276 B.n35 516.524
R263 B.n70 B.t9 207.094
R264 B.n78 B.t0 207.094
R265 B.n22 B.t3 207.094
R266 B.n28 B.t6 207.094
R267 B.n140 B.n139 163.367
R268 B.n139 B.n138 163.367
R269 B.n138 B.n85 163.367
R270 B.n134 B.n85 163.367
R271 B.n134 B.n133 163.367
R272 B.n133 B.n132 163.367
R273 B.n132 B.n87 163.367
R274 B.n128 B.n87 163.367
R275 B.n128 B.n127 163.367
R276 B.n127 B.n126 163.367
R277 B.n126 B.n89 163.367
R278 B.n122 B.n89 163.367
R279 B.n122 B.n121 163.367
R280 B.n121 B.n120 163.367
R281 B.n120 B.n91 163.367
R282 B.n116 B.n91 163.367
R283 B.n116 B.n115 163.367
R284 B.n115 B.n114 163.367
R285 B.n114 B.n93 163.367
R286 B.n110 B.n93 163.367
R287 B.n110 B.n109 163.367
R288 B.n109 B.n108 163.367
R289 B.n108 B.n95 163.367
R290 B.n104 B.n95 163.367
R291 B.n104 B.n103 163.367
R292 B.n103 B.n102 163.367
R293 B.n102 B.n97 163.367
R294 B.n98 B.n97 163.367
R295 B.n98 B.n2 163.367
R296 B.n362 B.n2 163.367
R297 B.n362 B.n361 163.367
R298 B.n361 B.n360 163.367
R299 B.n360 B.n3 163.367
R300 B.n356 B.n3 163.367
R301 B.n356 B.n355 163.367
R302 B.n355 B.n354 163.367
R303 B.n354 B.n5 163.367
R304 B.n350 B.n5 163.367
R305 B.n350 B.n349 163.367
R306 B.n349 B.n348 163.367
R307 B.n348 B.n7 163.367
R308 B.n344 B.n7 163.367
R309 B.n344 B.n343 163.367
R310 B.n343 B.n342 163.367
R311 B.n342 B.n9 163.367
R312 B.n338 B.n9 163.367
R313 B.n338 B.n337 163.367
R314 B.n337 B.n336 163.367
R315 B.n336 B.n11 163.367
R316 B.n332 B.n11 163.367
R317 B.n332 B.n331 163.367
R318 B.n331 B.n330 163.367
R319 B.n330 B.n13 163.367
R320 B.n326 B.n13 163.367
R321 B.n326 B.n325 163.367
R322 B.n325 B.n324 163.367
R323 B.n324 B.n15 163.367
R324 B.n320 B.n15 163.367
R325 B.n320 B.n319 163.367
R326 B.n319 B.n318 163.367
R327 B.n144 B.n83 163.367
R328 B.n145 B.n144 163.367
R329 B.n146 B.n145 163.367
R330 B.n146 B.n81 163.367
R331 B.n150 B.n81 163.367
R332 B.n151 B.n150 163.367
R333 B.n152 B.n151 163.367
R334 B.n152 B.n77 163.367
R335 B.n157 B.n77 163.367
R336 B.n158 B.n157 163.367
R337 B.n159 B.n158 163.367
R338 B.n159 B.n75 163.367
R339 B.n163 B.n75 163.367
R340 B.n164 B.n163 163.367
R341 B.n165 B.n164 163.367
R342 B.n165 B.n73 163.367
R343 B.n169 B.n73 163.367
R344 B.n170 B.n169 163.367
R345 B.n170 B.n69 163.367
R346 B.n174 B.n69 163.367
R347 B.n175 B.n174 163.367
R348 B.n176 B.n175 163.367
R349 B.n176 B.n67 163.367
R350 B.n180 B.n67 163.367
R351 B.n181 B.n180 163.367
R352 B.n182 B.n181 163.367
R353 B.n186 B.n65 163.367
R354 B.n187 B.n186 163.367
R355 B.n188 B.n187 163.367
R356 B.n188 B.n63 163.367
R357 B.n192 B.n63 163.367
R358 B.n193 B.n192 163.367
R359 B.n194 B.n193 163.367
R360 B.n194 B.n61 163.367
R361 B.n198 B.n61 163.367
R362 B.n199 B.n198 163.367
R363 B.n200 B.n199 163.367
R364 B.n200 B.n59 163.367
R365 B.n204 B.n59 163.367
R366 B.n205 B.n204 163.367
R367 B.n206 B.n205 163.367
R368 B.n206 B.n57 163.367
R369 B.n210 B.n57 163.367
R370 B.n211 B.n210 163.367
R371 B.n212 B.n211 163.367
R372 B.n212 B.n55 163.367
R373 B.n216 B.n55 163.367
R374 B.n217 B.n216 163.367
R375 B.n218 B.n217 163.367
R376 B.n218 B.n53 163.367
R377 B.n222 B.n53 163.367
R378 B.n223 B.n222 163.367
R379 B.n224 B.n223 163.367
R380 B.n224 B.n51 163.367
R381 B.n228 B.n51 163.367
R382 B.n229 B.n228 163.367
R383 B.n230 B.n229 163.367
R384 B.n230 B.n49 163.367
R385 B.n234 B.n49 163.367
R386 B.n235 B.n234 163.367
R387 B.n236 B.n235 163.367
R388 B.n236 B.n47 163.367
R389 B.n240 B.n47 163.367
R390 B.n241 B.n240 163.367
R391 B.n242 B.n241 163.367
R392 B.n242 B.n45 163.367
R393 B.n246 B.n45 163.367
R394 B.n247 B.n246 163.367
R395 B.n248 B.n247 163.367
R396 B.n248 B.n43 163.367
R397 B.n252 B.n43 163.367
R398 B.n253 B.n252 163.367
R399 B.n254 B.n253 163.367
R400 B.n254 B.n41 163.367
R401 B.n258 B.n41 163.367
R402 B.n259 B.n258 163.367
R403 B.n260 B.n259 163.367
R404 B.n260 B.n39 163.367
R405 B.n264 B.n39 163.367
R406 B.n265 B.n264 163.367
R407 B.n266 B.n265 163.367
R408 B.n266 B.n37 163.367
R409 B.n270 B.n37 163.367
R410 B.n271 B.n270 163.367
R411 B.n272 B.n271 163.367
R412 B.n272 B.n35 163.367
R413 B.n314 B.n17 163.367
R414 B.n314 B.n313 163.367
R415 B.n313 B.n312 163.367
R416 B.n312 B.n19 163.367
R417 B.n308 B.n19 163.367
R418 B.n308 B.n307 163.367
R419 B.n307 B.n306 163.367
R420 B.n306 B.n21 163.367
R421 B.n301 B.n21 163.367
R422 B.n301 B.n300 163.367
R423 B.n300 B.n299 163.367
R424 B.n299 B.n25 163.367
R425 B.n295 B.n25 163.367
R426 B.n295 B.n294 163.367
R427 B.n294 B.n293 163.367
R428 B.n293 B.n27 163.367
R429 B.n289 B.n27 163.367
R430 B.n289 B.n288 163.367
R431 B.n288 B.n31 163.367
R432 B.n284 B.n31 163.367
R433 B.n284 B.n283 163.367
R434 B.n283 B.n282 163.367
R435 B.n282 B.n33 163.367
R436 B.n278 B.n33 163.367
R437 B.n278 B.n277 163.367
R438 B.n277 B.n276 163.367
R439 B.n72 B.n71 59.5399
R440 B.n155 B.n79 59.5399
R441 B.n303 B.n23 59.5399
R442 B.n30 B.n29 59.5399
R443 B.n71 B.n70 36.0732
R444 B.n79 B.n78 36.0732
R445 B.n23 B.n22 36.0732
R446 B.n29 B.n28 36.0732
R447 B.n317 B.n316 33.5615
R448 B.n275 B.n274 33.5615
R449 B.n184 B.n183 33.5615
R450 B.n142 B.n141 33.5615
R451 B B.n363 18.0485
R452 B.n316 B.n315 10.6151
R453 B.n315 B.n18 10.6151
R454 B.n311 B.n18 10.6151
R455 B.n311 B.n310 10.6151
R456 B.n310 B.n309 10.6151
R457 B.n309 B.n20 10.6151
R458 B.n305 B.n20 10.6151
R459 B.n305 B.n304 10.6151
R460 B.n302 B.n24 10.6151
R461 B.n298 B.n24 10.6151
R462 B.n298 B.n297 10.6151
R463 B.n297 B.n296 10.6151
R464 B.n296 B.n26 10.6151
R465 B.n292 B.n26 10.6151
R466 B.n292 B.n291 10.6151
R467 B.n291 B.n290 10.6151
R468 B.n287 B.n286 10.6151
R469 B.n286 B.n285 10.6151
R470 B.n285 B.n32 10.6151
R471 B.n281 B.n32 10.6151
R472 B.n281 B.n280 10.6151
R473 B.n280 B.n279 10.6151
R474 B.n279 B.n34 10.6151
R475 B.n275 B.n34 10.6151
R476 B.n185 B.n184 10.6151
R477 B.n185 B.n64 10.6151
R478 B.n189 B.n64 10.6151
R479 B.n190 B.n189 10.6151
R480 B.n191 B.n190 10.6151
R481 B.n191 B.n62 10.6151
R482 B.n195 B.n62 10.6151
R483 B.n196 B.n195 10.6151
R484 B.n197 B.n196 10.6151
R485 B.n197 B.n60 10.6151
R486 B.n201 B.n60 10.6151
R487 B.n202 B.n201 10.6151
R488 B.n203 B.n202 10.6151
R489 B.n203 B.n58 10.6151
R490 B.n207 B.n58 10.6151
R491 B.n208 B.n207 10.6151
R492 B.n209 B.n208 10.6151
R493 B.n209 B.n56 10.6151
R494 B.n213 B.n56 10.6151
R495 B.n214 B.n213 10.6151
R496 B.n215 B.n214 10.6151
R497 B.n215 B.n54 10.6151
R498 B.n219 B.n54 10.6151
R499 B.n220 B.n219 10.6151
R500 B.n221 B.n220 10.6151
R501 B.n221 B.n52 10.6151
R502 B.n225 B.n52 10.6151
R503 B.n226 B.n225 10.6151
R504 B.n227 B.n226 10.6151
R505 B.n227 B.n50 10.6151
R506 B.n231 B.n50 10.6151
R507 B.n232 B.n231 10.6151
R508 B.n233 B.n232 10.6151
R509 B.n233 B.n48 10.6151
R510 B.n237 B.n48 10.6151
R511 B.n238 B.n237 10.6151
R512 B.n239 B.n238 10.6151
R513 B.n239 B.n46 10.6151
R514 B.n243 B.n46 10.6151
R515 B.n244 B.n243 10.6151
R516 B.n245 B.n244 10.6151
R517 B.n245 B.n44 10.6151
R518 B.n249 B.n44 10.6151
R519 B.n250 B.n249 10.6151
R520 B.n251 B.n250 10.6151
R521 B.n251 B.n42 10.6151
R522 B.n255 B.n42 10.6151
R523 B.n256 B.n255 10.6151
R524 B.n257 B.n256 10.6151
R525 B.n257 B.n40 10.6151
R526 B.n261 B.n40 10.6151
R527 B.n262 B.n261 10.6151
R528 B.n263 B.n262 10.6151
R529 B.n263 B.n38 10.6151
R530 B.n267 B.n38 10.6151
R531 B.n268 B.n267 10.6151
R532 B.n269 B.n268 10.6151
R533 B.n269 B.n36 10.6151
R534 B.n273 B.n36 10.6151
R535 B.n274 B.n273 10.6151
R536 B.n143 B.n142 10.6151
R537 B.n143 B.n82 10.6151
R538 B.n147 B.n82 10.6151
R539 B.n148 B.n147 10.6151
R540 B.n149 B.n148 10.6151
R541 B.n149 B.n80 10.6151
R542 B.n153 B.n80 10.6151
R543 B.n154 B.n153 10.6151
R544 B.n156 B.n76 10.6151
R545 B.n160 B.n76 10.6151
R546 B.n161 B.n160 10.6151
R547 B.n162 B.n161 10.6151
R548 B.n162 B.n74 10.6151
R549 B.n166 B.n74 10.6151
R550 B.n167 B.n166 10.6151
R551 B.n168 B.n167 10.6151
R552 B.n172 B.n171 10.6151
R553 B.n173 B.n172 10.6151
R554 B.n173 B.n68 10.6151
R555 B.n177 B.n68 10.6151
R556 B.n178 B.n177 10.6151
R557 B.n179 B.n178 10.6151
R558 B.n179 B.n66 10.6151
R559 B.n183 B.n66 10.6151
R560 B.n141 B.n84 10.6151
R561 B.n137 B.n84 10.6151
R562 B.n137 B.n136 10.6151
R563 B.n136 B.n135 10.6151
R564 B.n135 B.n86 10.6151
R565 B.n131 B.n86 10.6151
R566 B.n131 B.n130 10.6151
R567 B.n130 B.n129 10.6151
R568 B.n129 B.n88 10.6151
R569 B.n125 B.n88 10.6151
R570 B.n125 B.n124 10.6151
R571 B.n124 B.n123 10.6151
R572 B.n123 B.n90 10.6151
R573 B.n119 B.n90 10.6151
R574 B.n119 B.n118 10.6151
R575 B.n118 B.n117 10.6151
R576 B.n117 B.n92 10.6151
R577 B.n113 B.n92 10.6151
R578 B.n113 B.n112 10.6151
R579 B.n112 B.n111 10.6151
R580 B.n111 B.n94 10.6151
R581 B.n107 B.n94 10.6151
R582 B.n107 B.n106 10.6151
R583 B.n106 B.n105 10.6151
R584 B.n105 B.n96 10.6151
R585 B.n101 B.n96 10.6151
R586 B.n101 B.n100 10.6151
R587 B.n100 B.n99 10.6151
R588 B.n99 B.n0 10.6151
R589 B.n359 B.n1 10.6151
R590 B.n359 B.n358 10.6151
R591 B.n358 B.n357 10.6151
R592 B.n357 B.n4 10.6151
R593 B.n353 B.n4 10.6151
R594 B.n353 B.n352 10.6151
R595 B.n352 B.n351 10.6151
R596 B.n351 B.n6 10.6151
R597 B.n347 B.n6 10.6151
R598 B.n347 B.n346 10.6151
R599 B.n346 B.n345 10.6151
R600 B.n345 B.n8 10.6151
R601 B.n341 B.n8 10.6151
R602 B.n341 B.n340 10.6151
R603 B.n340 B.n339 10.6151
R604 B.n339 B.n10 10.6151
R605 B.n335 B.n10 10.6151
R606 B.n335 B.n334 10.6151
R607 B.n334 B.n333 10.6151
R608 B.n333 B.n12 10.6151
R609 B.n329 B.n12 10.6151
R610 B.n329 B.n328 10.6151
R611 B.n328 B.n327 10.6151
R612 B.n327 B.n14 10.6151
R613 B.n323 B.n14 10.6151
R614 B.n323 B.n322 10.6151
R615 B.n322 B.n321 10.6151
R616 B.n321 B.n16 10.6151
R617 B.n317 B.n16 10.6151
R618 B.n303 B.n302 6.5566
R619 B.n290 B.n30 6.5566
R620 B.n156 B.n155 6.5566
R621 B.n168 B.n72 6.5566
R622 B.n304 B.n303 4.05904
R623 B.n287 B.n30 4.05904
R624 B.n155 B.n154 4.05904
R625 B.n171 B.n72 4.05904
R626 B.n363 B.n0 2.81026
R627 B.n363 B.n1 2.81026
R628 VP.n17 VP.n16 180.385
R629 VP.n32 VP.n31 180.385
R630 VP.n15 VP.n14 180.385
R631 VP.n9 VP.n8 161.3
R632 VP.n10 VP.n5 161.3
R633 VP.n12 VP.n11 161.3
R634 VP.n13 VP.n4 161.3
R635 VP.n30 VP.n0 161.3
R636 VP.n29 VP.n28 161.3
R637 VP.n27 VP.n1 161.3
R638 VP.n26 VP.n25 161.3
R639 VP.n23 VP.n2 161.3
R640 VP.n22 VP.n21 161.3
R641 VP.n20 VP.n3 161.3
R642 VP.n19 VP.n18 161.3
R643 VP.n29 VP.n1 56.5193
R644 VP.n22 VP.n3 56.5193
R645 VP.n12 VP.n5 56.5193
R646 VP.n7 VP.n6 53.6827
R647 VP.n6 VP.t3 44.6322
R648 VP.n16 VP.n15 35.8944
R649 VP.n18 VP.n3 24.4675
R650 VP.n23 VP.n22 24.4675
R651 VP.n25 VP.n1 24.4675
R652 VP.n30 VP.n29 24.4675
R653 VP.n13 VP.n12 24.4675
R654 VP.n8 VP.n5 24.4675
R655 VP.n9 VP.n6 18.2406
R656 VP.n17 VP.t1 13.3894
R657 VP.n24 VP.t4 13.3894
R658 VP.n31 VP.t0 13.3894
R659 VP.n14 VP.t5 13.3894
R660 VP.n7 VP.t2 13.3894
R661 VP.n24 VP.n23 12.234
R662 VP.n25 VP.n24 12.234
R663 VP.n8 VP.n7 12.234
R664 VP.n18 VP.n17 5.38324
R665 VP.n31 VP.n30 5.38324
R666 VP.n14 VP.n13 5.38324
R667 VP.n10 VP.n9 0.189894
R668 VP.n11 VP.n10 0.189894
R669 VP.n11 VP.n4 0.189894
R670 VP.n15 VP.n4 0.189894
R671 VP.n19 VP.n16 0.189894
R672 VP.n20 VP.n19 0.189894
R673 VP.n21 VP.n20 0.189894
R674 VP.n21 VP.n2 0.189894
R675 VP.n26 VP.n2 0.189894
R676 VP.n27 VP.n26 0.189894
R677 VP.n28 VP.n27 0.189894
R678 VP.n28 VP.n0 0.189894
R679 VP.n32 VP.n0 0.189894
R680 VP VP.n32 0.0516364
R681 VDD1 VDD1.t2 676.726
R682 VDD1.n1 VDD1.t4 676.611
R683 VDD1.n1 VDD1.n0 637.568
R684 VDD1.n3 VDD1.n2 637.223
R685 VDD1.n2 VDD1.t3 38.2417
R686 VDD1.n2 VDD1.t0 38.2417
R687 VDD1.n0 VDD1.t1 38.2417
R688 VDD1.n0 VDD1.t5 38.2417
R689 VDD1.n3 VDD1.n1 31.044
R690 VDD1 VDD1.n3 0.343172
C0 VN VDD1 0.157411f
C1 w_n2458_n1138# VTAIL 1.19103f
C2 w_n2458_n1138# B 5.09422f
C3 VP w_n2458_n1138# 4.47326f
C4 VN VTAIL 1.37814f
C5 VN B 0.77295f
C6 VN VP 3.83383f
C7 VTAIL VDD1 2.90266f
C8 B VDD1 0.950334f
C9 VP VDD1 0.974304f
C10 VTAIL B 0.821985f
C11 VP VTAIL 1.39227f
C12 VP B 1.29182f
C13 VDD2 w_n2458_n1138# 1.27259f
C14 VN VDD2 0.758255f
C15 VDD2 VDD1 1.01696f
C16 VDD2 VTAIL 2.94875f
C17 VDD2 B 0.999362f
C18 VP VDD2 0.376113f
C19 VN w_n2458_n1138# 4.16673f
C20 w_n2458_n1138# VDD1 1.22308f
C21 VDD2 VSUBS 0.757604f
C22 VDD1 VSUBS 1.077063f
C23 VTAIL VSUBS 0.332582f
C24 VN VSUBS 4.33125f
C25 VP VSUBS 1.530165f
C26 B VSUBS 2.487722f
C27 w_n2458_n1138# VSUBS 36.132603f
C28 VDD1.t2 VSUBS 0.061887f
C29 VDD1.t4 VSUBS 0.061841f
C30 VDD1.t1 VSUBS 0.01188f
C31 VDD1.t5 VSUBS 0.01188f
C32 VDD1.n0 VSUBS 0.032211f
C33 VDD1.n1 VSUBS 1.25259f
C34 VDD1.t3 VSUBS 0.01188f
C35 VDD1.t0 VSUBS 0.01188f
C36 VDD1.n2 VSUBS 0.032078f
C37 VDD1.n3 VSUBS 1.11298f
C38 VP.n0 VSUBS 0.060011f
C39 VP.t0 VSUBS 0.132946f
C40 VP.n1 VSUBS 0.0759f
C41 VP.n2 VSUBS 0.060011f
C42 VP.t4 VSUBS 0.132946f
C43 VP.n3 VSUBS 0.099312f
C44 VP.n4 VSUBS 0.060011f
C45 VP.t5 VSUBS 0.132946f
C46 VP.n5 VSUBS 0.0759f
C47 VP.t3 VSUBS 0.386214f
C48 VP.n6 VSUBS 0.210055f
C49 VP.t2 VSUBS 0.132946f
C50 VP.n7 VSUBS 0.241217f
C51 VP.n8 VSUBS 0.084236f
C52 VP.n9 VSUBS 0.376558f
C53 VP.n10 VSUBS 0.060011f
C54 VP.n11 VSUBS 0.060011f
C55 VP.n12 VSUBS 0.099312f
C56 VP.n13 VSUBS 0.068775f
C57 VP.n14 VSUBS 0.241963f
C58 VP.n15 VSUBS 1.8898f
C59 VP.n16 VSUBS 1.9499f
C60 VP.t1 VSUBS 0.132946f
C61 VP.n17 VSUBS 0.241963f
C62 VP.n18 VSUBS 0.068775f
C63 VP.n19 VSUBS 0.060011f
C64 VP.n20 VSUBS 0.060011f
C65 VP.n21 VSUBS 0.060011f
C66 VP.n22 VSUBS 0.0759f
C67 VP.n23 VSUBS 0.084236f
C68 VP.n24 VSUBS 0.128125f
C69 VP.n25 VSUBS 0.084236f
C70 VP.n26 VSUBS 0.060011f
C71 VP.n27 VSUBS 0.060011f
C72 VP.n28 VSUBS 0.060011f
C73 VP.n29 VSUBS 0.099312f
C74 VP.n30 VSUBS 0.068775f
C75 VP.n31 VSUBS 0.241963f
C76 VP.n32 VSUBS 0.059975f
C77 B.n0 VSUBS 0.006583f
C78 B.n1 VSUBS 0.006583f
C79 B.n2 VSUBS 0.01041f
C80 B.n3 VSUBS 0.01041f
C81 B.n4 VSUBS 0.01041f
C82 B.n5 VSUBS 0.01041f
C83 B.n6 VSUBS 0.01041f
C84 B.n7 VSUBS 0.01041f
C85 B.n8 VSUBS 0.01041f
C86 B.n9 VSUBS 0.01041f
C87 B.n10 VSUBS 0.01041f
C88 B.n11 VSUBS 0.01041f
C89 B.n12 VSUBS 0.01041f
C90 B.n13 VSUBS 0.01041f
C91 B.n14 VSUBS 0.01041f
C92 B.n15 VSUBS 0.01041f
C93 B.n16 VSUBS 0.01041f
C94 B.n17 VSUBS 0.025253f
C95 B.n18 VSUBS 0.01041f
C96 B.n19 VSUBS 0.01041f
C97 B.n20 VSUBS 0.01041f
C98 B.n21 VSUBS 0.01041f
C99 B.t5 VSUBS 0.024363f
C100 B.t4 VSUBS 0.026627f
C101 B.t3 VSUBS 0.100932f
C102 B.n22 VSUBS 0.067995f
C103 B.n23 VSUBS 0.057872f
C104 B.n24 VSUBS 0.01041f
C105 B.n25 VSUBS 0.01041f
C106 B.n26 VSUBS 0.01041f
C107 B.n27 VSUBS 0.01041f
C108 B.t8 VSUBS 0.024363f
C109 B.t7 VSUBS 0.026627f
C110 B.t6 VSUBS 0.100932f
C111 B.n28 VSUBS 0.067995f
C112 B.n29 VSUBS 0.057872f
C113 B.n30 VSUBS 0.024119f
C114 B.n31 VSUBS 0.01041f
C115 B.n32 VSUBS 0.01041f
C116 B.n33 VSUBS 0.01041f
C117 B.n34 VSUBS 0.01041f
C118 B.n35 VSUBS 0.024348f
C119 B.n36 VSUBS 0.01041f
C120 B.n37 VSUBS 0.01041f
C121 B.n38 VSUBS 0.01041f
C122 B.n39 VSUBS 0.01041f
C123 B.n40 VSUBS 0.01041f
C124 B.n41 VSUBS 0.01041f
C125 B.n42 VSUBS 0.01041f
C126 B.n43 VSUBS 0.01041f
C127 B.n44 VSUBS 0.01041f
C128 B.n45 VSUBS 0.01041f
C129 B.n46 VSUBS 0.01041f
C130 B.n47 VSUBS 0.01041f
C131 B.n48 VSUBS 0.01041f
C132 B.n49 VSUBS 0.01041f
C133 B.n50 VSUBS 0.01041f
C134 B.n51 VSUBS 0.01041f
C135 B.n52 VSUBS 0.01041f
C136 B.n53 VSUBS 0.01041f
C137 B.n54 VSUBS 0.01041f
C138 B.n55 VSUBS 0.01041f
C139 B.n56 VSUBS 0.01041f
C140 B.n57 VSUBS 0.01041f
C141 B.n58 VSUBS 0.01041f
C142 B.n59 VSUBS 0.01041f
C143 B.n60 VSUBS 0.01041f
C144 B.n61 VSUBS 0.01041f
C145 B.n62 VSUBS 0.01041f
C146 B.n63 VSUBS 0.01041f
C147 B.n64 VSUBS 0.01041f
C148 B.n65 VSUBS 0.024348f
C149 B.n66 VSUBS 0.01041f
C150 B.n67 VSUBS 0.01041f
C151 B.n68 VSUBS 0.01041f
C152 B.n69 VSUBS 0.01041f
C153 B.t10 VSUBS 0.024363f
C154 B.t11 VSUBS 0.026627f
C155 B.t9 VSUBS 0.100932f
C156 B.n70 VSUBS 0.067995f
C157 B.n71 VSUBS 0.057872f
C158 B.n72 VSUBS 0.024119f
C159 B.n73 VSUBS 0.01041f
C160 B.n74 VSUBS 0.01041f
C161 B.n75 VSUBS 0.01041f
C162 B.n76 VSUBS 0.01041f
C163 B.n77 VSUBS 0.01041f
C164 B.t1 VSUBS 0.024363f
C165 B.t2 VSUBS 0.026627f
C166 B.t0 VSUBS 0.100932f
C167 B.n78 VSUBS 0.067995f
C168 B.n79 VSUBS 0.057872f
C169 B.n80 VSUBS 0.01041f
C170 B.n81 VSUBS 0.01041f
C171 B.n82 VSUBS 0.01041f
C172 B.n83 VSUBS 0.025253f
C173 B.n84 VSUBS 0.01041f
C174 B.n85 VSUBS 0.01041f
C175 B.n86 VSUBS 0.01041f
C176 B.n87 VSUBS 0.01041f
C177 B.n88 VSUBS 0.01041f
C178 B.n89 VSUBS 0.01041f
C179 B.n90 VSUBS 0.01041f
C180 B.n91 VSUBS 0.01041f
C181 B.n92 VSUBS 0.01041f
C182 B.n93 VSUBS 0.01041f
C183 B.n94 VSUBS 0.01041f
C184 B.n95 VSUBS 0.01041f
C185 B.n96 VSUBS 0.01041f
C186 B.n97 VSUBS 0.01041f
C187 B.n98 VSUBS 0.01041f
C188 B.n99 VSUBS 0.01041f
C189 B.n100 VSUBS 0.01041f
C190 B.n101 VSUBS 0.01041f
C191 B.n102 VSUBS 0.01041f
C192 B.n103 VSUBS 0.01041f
C193 B.n104 VSUBS 0.01041f
C194 B.n105 VSUBS 0.01041f
C195 B.n106 VSUBS 0.01041f
C196 B.n107 VSUBS 0.01041f
C197 B.n108 VSUBS 0.01041f
C198 B.n109 VSUBS 0.01041f
C199 B.n110 VSUBS 0.01041f
C200 B.n111 VSUBS 0.01041f
C201 B.n112 VSUBS 0.01041f
C202 B.n113 VSUBS 0.01041f
C203 B.n114 VSUBS 0.01041f
C204 B.n115 VSUBS 0.01041f
C205 B.n116 VSUBS 0.01041f
C206 B.n117 VSUBS 0.01041f
C207 B.n118 VSUBS 0.01041f
C208 B.n119 VSUBS 0.01041f
C209 B.n120 VSUBS 0.01041f
C210 B.n121 VSUBS 0.01041f
C211 B.n122 VSUBS 0.01041f
C212 B.n123 VSUBS 0.01041f
C213 B.n124 VSUBS 0.01041f
C214 B.n125 VSUBS 0.01041f
C215 B.n126 VSUBS 0.01041f
C216 B.n127 VSUBS 0.01041f
C217 B.n128 VSUBS 0.01041f
C218 B.n129 VSUBS 0.01041f
C219 B.n130 VSUBS 0.01041f
C220 B.n131 VSUBS 0.01041f
C221 B.n132 VSUBS 0.01041f
C222 B.n133 VSUBS 0.01041f
C223 B.n134 VSUBS 0.01041f
C224 B.n135 VSUBS 0.01041f
C225 B.n136 VSUBS 0.01041f
C226 B.n137 VSUBS 0.01041f
C227 B.n138 VSUBS 0.01041f
C228 B.n139 VSUBS 0.01041f
C229 B.n140 VSUBS 0.024348f
C230 B.n141 VSUBS 0.024348f
C231 B.n142 VSUBS 0.025253f
C232 B.n143 VSUBS 0.01041f
C233 B.n144 VSUBS 0.01041f
C234 B.n145 VSUBS 0.01041f
C235 B.n146 VSUBS 0.01041f
C236 B.n147 VSUBS 0.01041f
C237 B.n148 VSUBS 0.01041f
C238 B.n149 VSUBS 0.01041f
C239 B.n150 VSUBS 0.01041f
C240 B.n151 VSUBS 0.01041f
C241 B.n152 VSUBS 0.01041f
C242 B.n153 VSUBS 0.01041f
C243 B.n154 VSUBS 0.007195f
C244 B.n155 VSUBS 0.024119f
C245 B.n156 VSUBS 0.00842f
C246 B.n157 VSUBS 0.01041f
C247 B.n158 VSUBS 0.01041f
C248 B.n159 VSUBS 0.01041f
C249 B.n160 VSUBS 0.01041f
C250 B.n161 VSUBS 0.01041f
C251 B.n162 VSUBS 0.01041f
C252 B.n163 VSUBS 0.01041f
C253 B.n164 VSUBS 0.01041f
C254 B.n165 VSUBS 0.01041f
C255 B.n166 VSUBS 0.01041f
C256 B.n167 VSUBS 0.01041f
C257 B.n168 VSUBS 0.00842f
C258 B.n169 VSUBS 0.01041f
C259 B.n170 VSUBS 0.01041f
C260 B.n171 VSUBS 0.007195f
C261 B.n172 VSUBS 0.01041f
C262 B.n173 VSUBS 0.01041f
C263 B.n174 VSUBS 0.01041f
C264 B.n175 VSUBS 0.01041f
C265 B.n176 VSUBS 0.01041f
C266 B.n177 VSUBS 0.01041f
C267 B.n178 VSUBS 0.01041f
C268 B.n179 VSUBS 0.01041f
C269 B.n180 VSUBS 0.01041f
C270 B.n181 VSUBS 0.01041f
C271 B.n182 VSUBS 0.025253f
C272 B.n183 VSUBS 0.025253f
C273 B.n184 VSUBS 0.024348f
C274 B.n185 VSUBS 0.01041f
C275 B.n186 VSUBS 0.01041f
C276 B.n187 VSUBS 0.01041f
C277 B.n188 VSUBS 0.01041f
C278 B.n189 VSUBS 0.01041f
C279 B.n190 VSUBS 0.01041f
C280 B.n191 VSUBS 0.01041f
C281 B.n192 VSUBS 0.01041f
C282 B.n193 VSUBS 0.01041f
C283 B.n194 VSUBS 0.01041f
C284 B.n195 VSUBS 0.01041f
C285 B.n196 VSUBS 0.01041f
C286 B.n197 VSUBS 0.01041f
C287 B.n198 VSUBS 0.01041f
C288 B.n199 VSUBS 0.01041f
C289 B.n200 VSUBS 0.01041f
C290 B.n201 VSUBS 0.01041f
C291 B.n202 VSUBS 0.01041f
C292 B.n203 VSUBS 0.01041f
C293 B.n204 VSUBS 0.01041f
C294 B.n205 VSUBS 0.01041f
C295 B.n206 VSUBS 0.01041f
C296 B.n207 VSUBS 0.01041f
C297 B.n208 VSUBS 0.01041f
C298 B.n209 VSUBS 0.01041f
C299 B.n210 VSUBS 0.01041f
C300 B.n211 VSUBS 0.01041f
C301 B.n212 VSUBS 0.01041f
C302 B.n213 VSUBS 0.01041f
C303 B.n214 VSUBS 0.01041f
C304 B.n215 VSUBS 0.01041f
C305 B.n216 VSUBS 0.01041f
C306 B.n217 VSUBS 0.01041f
C307 B.n218 VSUBS 0.01041f
C308 B.n219 VSUBS 0.01041f
C309 B.n220 VSUBS 0.01041f
C310 B.n221 VSUBS 0.01041f
C311 B.n222 VSUBS 0.01041f
C312 B.n223 VSUBS 0.01041f
C313 B.n224 VSUBS 0.01041f
C314 B.n225 VSUBS 0.01041f
C315 B.n226 VSUBS 0.01041f
C316 B.n227 VSUBS 0.01041f
C317 B.n228 VSUBS 0.01041f
C318 B.n229 VSUBS 0.01041f
C319 B.n230 VSUBS 0.01041f
C320 B.n231 VSUBS 0.01041f
C321 B.n232 VSUBS 0.01041f
C322 B.n233 VSUBS 0.01041f
C323 B.n234 VSUBS 0.01041f
C324 B.n235 VSUBS 0.01041f
C325 B.n236 VSUBS 0.01041f
C326 B.n237 VSUBS 0.01041f
C327 B.n238 VSUBS 0.01041f
C328 B.n239 VSUBS 0.01041f
C329 B.n240 VSUBS 0.01041f
C330 B.n241 VSUBS 0.01041f
C331 B.n242 VSUBS 0.01041f
C332 B.n243 VSUBS 0.01041f
C333 B.n244 VSUBS 0.01041f
C334 B.n245 VSUBS 0.01041f
C335 B.n246 VSUBS 0.01041f
C336 B.n247 VSUBS 0.01041f
C337 B.n248 VSUBS 0.01041f
C338 B.n249 VSUBS 0.01041f
C339 B.n250 VSUBS 0.01041f
C340 B.n251 VSUBS 0.01041f
C341 B.n252 VSUBS 0.01041f
C342 B.n253 VSUBS 0.01041f
C343 B.n254 VSUBS 0.01041f
C344 B.n255 VSUBS 0.01041f
C345 B.n256 VSUBS 0.01041f
C346 B.n257 VSUBS 0.01041f
C347 B.n258 VSUBS 0.01041f
C348 B.n259 VSUBS 0.01041f
C349 B.n260 VSUBS 0.01041f
C350 B.n261 VSUBS 0.01041f
C351 B.n262 VSUBS 0.01041f
C352 B.n263 VSUBS 0.01041f
C353 B.n264 VSUBS 0.01041f
C354 B.n265 VSUBS 0.01041f
C355 B.n266 VSUBS 0.01041f
C356 B.n267 VSUBS 0.01041f
C357 B.n268 VSUBS 0.01041f
C358 B.n269 VSUBS 0.01041f
C359 B.n270 VSUBS 0.01041f
C360 B.n271 VSUBS 0.01041f
C361 B.n272 VSUBS 0.01041f
C362 B.n273 VSUBS 0.01041f
C363 B.n274 VSUBS 0.025544f
C364 B.n275 VSUBS 0.024056f
C365 B.n276 VSUBS 0.025253f
C366 B.n277 VSUBS 0.01041f
C367 B.n278 VSUBS 0.01041f
C368 B.n279 VSUBS 0.01041f
C369 B.n280 VSUBS 0.01041f
C370 B.n281 VSUBS 0.01041f
C371 B.n282 VSUBS 0.01041f
C372 B.n283 VSUBS 0.01041f
C373 B.n284 VSUBS 0.01041f
C374 B.n285 VSUBS 0.01041f
C375 B.n286 VSUBS 0.01041f
C376 B.n287 VSUBS 0.007195f
C377 B.n288 VSUBS 0.01041f
C378 B.n289 VSUBS 0.01041f
C379 B.n290 VSUBS 0.00842f
C380 B.n291 VSUBS 0.01041f
C381 B.n292 VSUBS 0.01041f
C382 B.n293 VSUBS 0.01041f
C383 B.n294 VSUBS 0.01041f
C384 B.n295 VSUBS 0.01041f
C385 B.n296 VSUBS 0.01041f
C386 B.n297 VSUBS 0.01041f
C387 B.n298 VSUBS 0.01041f
C388 B.n299 VSUBS 0.01041f
C389 B.n300 VSUBS 0.01041f
C390 B.n301 VSUBS 0.01041f
C391 B.n302 VSUBS 0.00842f
C392 B.n303 VSUBS 0.024119f
C393 B.n304 VSUBS 0.007195f
C394 B.n305 VSUBS 0.01041f
C395 B.n306 VSUBS 0.01041f
C396 B.n307 VSUBS 0.01041f
C397 B.n308 VSUBS 0.01041f
C398 B.n309 VSUBS 0.01041f
C399 B.n310 VSUBS 0.01041f
C400 B.n311 VSUBS 0.01041f
C401 B.n312 VSUBS 0.01041f
C402 B.n313 VSUBS 0.01041f
C403 B.n314 VSUBS 0.01041f
C404 B.n315 VSUBS 0.01041f
C405 B.n316 VSUBS 0.025253f
C406 B.n317 VSUBS 0.024348f
C407 B.n318 VSUBS 0.024348f
C408 B.n319 VSUBS 0.01041f
C409 B.n320 VSUBS 0.01041f
C410 B.n321 VSUBS 0.01041f
C411 B.n322 VSUBS 0.01041f
C412 B.n323 VSUBS 0.01041f
C413 B.n324 VSUBS 0.01041f
C414 B.n325 VSUBS 0.01041f
C415 B.n326 VSUBS 0.01041f
C416 B.n327 VSUBS 0.01041f
C417 B.n328 VSUBS 0.01041f
C418 B.n329 VSUBS 0.01041f
C419 B.n330 VSUBS 0.01041f
C420 B.n331 VSUBS 0.01041f
C421 B.n332 VSUBS 0.01041f
C422 B.n333 VSUBS 0.01041f
C423 B.n334 VSUBS 0.01041f
C424 B.n335 VSUBS 0.01041f
C425 B.n336 VSUBS 0.01041f
C426 B.n337 VSUBS 0.01041f
C427 B.n338 VSUBS 0.01041f
C428 B.n339 VSUBS 0.01041f
C429 B.n340 VSUBS 0.01041f
C430 B.n341 VSUBS 0.01041f
C431 B.n342 VSUBS 0.01041f
C432 B.n343 VSUBS 0.01041f
C433 B.n344 VSUBS 0.01041f
C434 B.n345 VSUBS 0.01041f
C435 B.n346 VSUBS 0.01041f
C436 B.n347 VSUBS 0.01041f
C437 B.n348 VSUBS 0.01041f
C438 B.n349 VSUBS 0.01041f
C439 B.n350 VSUBS 0.01041f
C440 B.n351 VSUBS 0.01041f
C441 B.n352 VSUBS 0.01041f
C442 B.n353 VSUBS 0.01041f
C443 B.n354 VSUBS 0.01041f
C444 B.n355 VSUBS 0.01041f
C445 B.n356 VSUBS 0.01041f
C446 B.n357 VSUBS 0.01041f
C447 B.n358 VSUBS 0.01041f
C448 B.n359 VSUBS 0.01041f
C449 B.n360 VSUBS 0.01041f
C450 B.n361 VSUBS 0.01041f
C451 B.n362 VSUBS 0.01041f
C452 B.n363 VSUBS 0.023572f
C453 VDD2.t4 VSUBS 0.063267f
C454 VDD2.t0 VSUBS 0.012153f
C455 VDD2.t1 VSUBS 0.012153f
C456 VDD2.n0 VSUBS 0.032954f
C457 VDD2.n1 VSUBS 1.21811f
C458 VDD2.t5 VSUBS 0.062917f
C459 VDD2.n2 VSUBS 1.09823f
C460 VDD2.t3 VSUBS 0.012153f
C461 VDD2.t2 VSUBS 0.012153f
C462 VDD2.n3 VSUBS 0.032952f
C463 VTAIL.t7 VSUBS 0.017252f
C464 VTAIL.t10 VSUBS 0.017252f
C465 VTAIL.n0 VSUBS 0.041801f
C466 VTAIL.n1 VSUBS 0.296029f
C467 VTAIL.t1 VSUBS 0.084696f
C468 VTAIL.n2 VSUBS 0.394898f
C469 VTAIL.t2 VSUBS 0.017252f
C470 VTAIL.t4 VSUBS 0.017252f
C471 VTAIL.n3 VSUBS 0.041801f
C472 VTAIL.n4 VSUBS 0.960453f
C473 VTAIL.t9 VSUBS 0.017252f
C474 VTAIL.t6 VSUBS 0.017252f
C475 VTAIL.n5 VSUBS 0.041801f
C476 VTAIL.n6 VSUBS 0.960453f
C477 VTAIL.t11 VSUBS 0.084696f
C478 VTAIL.n7 VSUBS 0.394897f
C479 VTAIL.t0 VSUBS 0.017252f
C480 VTAIL.t3 VSUBS 0.017252f
C481 VTAIL.n8 VSUBS 0.041801f
C482 VTAIL.n9 VSUBS 0.390741f
C483 VTAIL.t5 VSUBS 0.084696f
C484 VTAIL.n10 VSUBS 0.831905f
C485 VTAIL.t8 VSUBS 0.084696f
C486 VTAIL.n11 VSUBS 0.793913f
C487 VN.n0 VSUBS 0.05726f
C488 VN.t4 VSUBS 0.126851f
C489 VN.n1 VSUBS 0.07242f
C490 VN.t1 VSUBS 0.368509f
C491 VN.n2 VSUBS 0.200426f
C492 VN.t5 VSUBS 0.126851f
C493 VN.n3 VSUBS 0.230159f
C494 VN.n4 VSUBS 0.080375f
C495 VN.n5 VSUBS 0.359295f
C496 VN.n6 VSUBS 0.05726f
C497 VN.n7 VSUBS 0.05726f
C498 VN.n8 VSUBS 0.094759f
C499 VN.n9 VSUBS 0.065622f
C500 VN.n10 VSUBS 0.230871f
C501 VN.n11 VSUBS 0.057226f
C502 VN.n12 VSUBS 0.05726f
C503 VN.t0 VSUBS 0.126851f
C504 VN.n13 VSUBS 0.07242f
C505 VN.t3 VSUBS 0.368509f
C506 VN.n14 VSUBS 0.200426f
C507 VN.t2 VSUBS 0.126851f
C508 VN.n15 VSUBS 0.230159f
C509 VN.n16 VSUBS 0.080375f
C510 VN.n17 VSUBS 0.359295f
C511 VN.n18 VSUBS 0.05726f
C512 VN.n19 VSUBS 0.05726f
C513 VN.n20 VSUBS 0.094759f
C514 VN.n21 VSUBS 0.065622f
C515 VN.n22 VSUBS 0.230871f
C516 VN.n23 VSUBS 1.84115f
.ends

