* NGSPICE file created from diff_pair_sample_1594.ext - technology: sky130A

.subckt diff_pair_sample_1594 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X1 VTAIL.t5 VP.t0 VDD1.t7 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0.2508 ps=1.85 w=1.52 l=3.64
X2 B.t11 B.t9 B.t10 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0 ps=0 w=1.52 l=3.64
X3 B.t8 B.t6 B.t7 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0 ps=0 w=1.52 l=3.64
X4 VTAIL.t1 VP.t1 VDD1.t6 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0.2508 ps=1.85 w=1.52 l=3.64
X5 VDD1.t5 VP.t2 VTAIL.t2 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.5928 ps=3.82 w=1.52 l=3.64
X6 VTAIL.t14 VN.t1 VDD2.t2 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0.2508 ps=1.85 w=1.52 l=3.64
X7 VDD1.t4 VP.t3 VTAIL.t4 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X8 VDD2.t3 VN.t2 VTAIL.t13 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.5928 ps=3.82 w=1.52 l=3.64
X9 VDD1.t3 VP.t4 VTAIL.t6 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.5928 ps=3.82 w=1.52 l=3.64
X10 VDD2.t5 VN.t3 VTAIL.t12 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.5928 ps=3.82 w=1.52 l=3.64
X11 VTAIL.t11 VN.t4 VDD2.t4 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X12 VDD1.t2 VP.t5 VTAIL.t7 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X13 B.t5 B.t3 B.t4 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0 ps=0 w=1.52 l=3.64
X14 VDD2.t0 VN.t5 VTAIL.t10 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X15 VTAIL.t0 VP.t6 VDD1.t1 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X16 B.t2 B.t0 B.t1 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0 ps=0 w=1.52 l=3.64
X17 VTAIL.t3 VP.t7 VDD1.t0 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X18 VDD2.t6 VN.t6 VTAIL.t9 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.2508 pd=1.85 as=0.2508 ps=1.85 w=1.52 l=3.64
X19 VTAIL.t8 VN.t7 VDD2.t1 w_n4940_n1272# sky130_fd_pr__pfet_01v8 ad=0.5928 pd=3.82 as=0.2508 ps=1.85 w=1.52 l=3.64
R0 VN.n72 VN.n71 161.3
R1 VN.n70 VN.n38 161.3
R2 VN.n69 VN.n68 161.3
R3 VN.n67 VN.n39 161.3
R4 VN.n66 VN.n65 161.3
R5 VN.n64 VN.n40 161.3
R6 VN.n63 VN.n62 161.3
R7 VN.n61 VN.n41 161.3
R8 VN.n60 VN.n59 161.3
R9 VN.n58 VN.n42 161.3
R10 VN.n57 VN.n56 161.3
R11 VN.n55 VN.n44 161.3
R12 VN.n54 VN.n53 161.3
R13 VN.n52 VN.n45 161.3
R14 VN.n51 VN.n50 161.3
R15 VN.n49 VN.n46 161.3
R16 VN.n35 VN.n34 161.3
R17 VN.n33 VN.n1 161.3
R18 VN.n32 VN.n31 161.3
R19 VN.n30 VN.n2 161.3
R20 VN.n29 VN.n28 161.3
R21 VN.n27 VN.n3 161.3
R22 VN.n26 VN.n25 161.3
R23 VN.n24 VN.n4 161.3
R24 VN.n23 VN.n22 161.3
R25 VN.n20 VN.n5 161.3
R26 VN.n19 VN.n18 161.3
R27 VN.n17 VN.n6 161.3
R28 VN.n16 VN.n15 161.3
R29 VN.n14 VN.n7 161.3
R30 VN.n13 VN.n12 161.3
R31 VN.n11 VN.n8 161.3
R32 VN.n36 VN.n0 79.9102
R33 VN.n73 VN.n37 79.9102
R34 VN.n10 VN.n9 62.9336
R35 VN.n48 VN.n47 62.9336
R36 VN.n15 VN.n6 56.4773
R37 VN.n28 VN.n2 56.4773
R38 VN.n53 VN.n44 56.4773
R39 VN.n65 VN.n39 56.4773
R40 VN VN.n73 48.1115
R41 VN.n48 VN.t2 43.3814
R42 VN.n10 VN.t1 43.3814
R43 VN.n13 VN.n8 24.3439
R44 VN.n14 VN.n13 24.3439
R45 VN.n15 VN.n14 24.3439
R46 VN.n19 VN.n6 24.3439
R47 VN.n20 VN.n19 24.3439
R48 VN.n22 VN.n20 24.3439
R49 VN.n26 VN.n4 24.3439
R50 VN.n27 VN.n26 24.3439
R51 VN.n28 VN.n27 24.3439
R52 VN.n32 VN.n2 24.3439
R53 VN.n33 VN.n32 24.3439
R54 VN.n34 VN.n33 24.3439
R55 VN.n53 VN.n52 24.3439
R56 VN.n52 VN.n51 24.3439
R57 VN.n51 VN.n46 24.3439
R58 VN.n65 VN.n64 24.3439
R59 VN.n64 VN.n63 24.3439
R60 VN.n63 VN.n41 24.3439
R61 VN.n59 VN.n58 24.3439
R62 VN.n58 VN.n57 24.3439
R63 VN.n57 VN.n44 24.3439
R64 VN.n71 VN.n70 24.3439
R65 VN.n70 VN.n69 24.3439
R66 VN.n69 VN.n39 24.3439
R67 VN.n21 VN.n4 12.9025
R68 VN.n43 VN.n41 12.9025
R69 VN.n9 VN.n8 11.4419
R70 VN.n22 VN.n21 11.4419
R71 VN.n47 VN.n46 11.4419
R72 VN.n59 VN.n43 11.4419
R73 VN.n9 VN.t6 10.0642
R74 VN.n21 VN.t4 10.0642
R75 VN.n0 VN.t3 10.0642
R76 VN.n47 VN.t0 10.0642
R77 VN.n43 VN.t5 10.0642
R78 VN.n37 VN.t7 10.0642
R79 VN.n34 VN.n0 9.98131
R80 VN.n71 VN.n37 9.98131
R81 VN.n11 VN.n10 3.16878
R82 VN.n49 VN.n48 3.16878
R83 VN.n73 VN.n72 0.355081
R84 VN.n36 VN.n35 0.355081
R85 VN VN.n36 0.26685
R86 VN.n72 VN.n38 0.189894
R87 VN.n68 VN.n38 0.189894
R88 VN.n68 VN.n67 0.189894
R89 VN.n67 VN.n66 0.189894
R90 VN.n66 VN.n40 0.189894
R91 VN.n62 VN.n40 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n60 0.189894
R94 VN.n60 VN.n42 0.189894
R95 VN.n56 VN.n42 0.189894
R96 VN.n56 VN.n55 0.189894
R97 VN.n55 VN.n54 0.189894
R98 VN.n54 VN.n45 0.189894
R99 VN.n50 VN.n45 0.189894
R100 VN.n50 VN.n49 0.189894
R101 VN.n12 VN.n11 0.189894
R102 VN.n12 VN.n7 0.189894
R103 VN.n16 VN.n7 0.189894
R104 VN.n17 VN.n16 0.189894
R105 VN.n18 VN.n17 0.189894
R106 VN.n18 VN.n5 0.189894
R107 VN.n23 VN.n5 0.189894
R108 VN.n24 VN.n23 0.189894
R109 VN.n25 VN.n24 0.189894
R110 VN.n25 VN.n3 0.189894
R111 VN.n29 VN.n3 0.189894
R112 VN.n30 VN.n29 0.189894
R113 VN.n31 VN.n30 0.189894
R114 VN.n31 VN.n1 0.189894
R115 VN.n35 VN.n1 0.189894
R116 VDD2.n2 VDD2.n1 252.996
R117 VDD2.n2 VDD2.n0 252.996
R118 VDD2 VDD2.n5 252.994
R119 VDD2.n4 VDD2.n3 251.34
R120 VDD2.n4 VDD2.n2 40.4265
R121 VDD2.n5 VDD2.t7 21.3854
R122 VDD2.n5 VDD2.t3 21.3854
R123 VDD2.n3 VDD2.t1 21.3854
R124 VDD2.n3 VDD2.t0 21.3854
R125 VDD2.n1 VDD2.t4 21.3854
R126 VDD2.n1 VDD2.t5 21.3854
R127 VDD2.n0 VDD2.t2 21.3854
R128 VDD2.n0 VDD2.t6 21.3854
R129 VDD2 VDD2.n4 1.7699
R130 VTAIL.n11 VTAIL.t1 256.046
R131 VTAIL.n10 VTAIL.t13 256.046
R132 VTAIL.n7 VTAIL.t8 256.046
R133 VTAIL.n15 VTAIL.t12 256.046
R134 VTAIL.n2 VTAIL.t14 256.046
R135 VTAIL.n3 VTAIL.t6 256.046
R136 VTAIL.n6 VTAIL.t5 256.046
R137 VTAIL.n14 VTAIL.t2 256.046
R138 VTAIL.n13 VTAIL.n12 234.661
R139 VTAIL.n9 VTAIL.n8 234.661
R140 VTAIL.n1 VTAIL.n0 234.661
R141 VTAIL.n5 VTAIL.n4 234.661
R142 VTAIL.n0 VTAIL.t9 21.3854
R143 VTAIL.n0 VTAIL.t11 21.3854
R144 VTAIL.n4 VTAIL.t4 21.3854
R145 VTAIL.n4 VTAIL.t0 21.3854
R146 VTAIL.n12 VTAIL.t7 21.3854
R147 VTAIL.n12 VTAIL.t3 21.3854
R148 VTAIL.n8 VTAIL.t10 21.3854
R149 VTAIL.n8 VTAIL.t15 21.3854
R150 VTAIL.n15 VTAIL.n14 17.0996
R151 VTAIL.n7 VTAIL.n6 17.0996
R152 VTAIL.n9 VTAIL.n7 3.42291
R153 VTAIL.n10 VTAIL.n9 3.42291
R154 VTAIL.n13 VTAIL.n11 3.42291
R155 VTAIL.n14 VTAIL.n13 3.42291
R156 VTAIL.n6 VTAIL.n5 3.42291
R157 VTAIL.n5 VTAIL.n3 3.42291
R158 VTAIL.n2 VTAIL.n1 3.42291
R159 VTAIL VTAIL.n15 3.36472
R160 VTAIL.n11 VTAIL.n10 0.470328
R161 VTAIL.n3 VTAIL.n2 0.470328
R162 VTAIL VTAIL.n1 0.0586897
R163 VP.n24 VP.n21 161.3
R164 VP.n26 VP.n25 161.3
R165 VP.n27 VP.n20 161.3
R166 VP.n29 VP.n28 161.3
R167 VP.n30 VP.n19 161.3
R168 VP.n32 VP.n31 161.3
R169 VP.n33 VP.n18 161.3
R170 VP.n36 VP.n35 161.3
R171 VP.n37 VP.n17 161.3
R172 VP.n39 VP.n38 161.3
R173 VP.n40 VP.n16 161.3
R174 VP.n42 VP.n41 161.3
R175 VP.n43 VP.n15 161.3
R176 VP.n45 VP.n44 161.3
R177 VP.n46 VP.n14 161.3
R178 VP.n48 VP.n47 161.3
R179 VP.n89 VP.n88 161.3
R180 VP.n87 VP.n1 161.3
R181 VP.n86 VP.n85 161.3
R182 VP.n84 VP.n2 161.3
R183 VP.n83 VP.n82 161.3
R184 VP.n81 VP.n3 161.3
R185 VP.n80 VP.n79 161.3
R186 VP.n78 VP.n4 161.3
R187 VP.n77 VP.n76 161.3
R188 VP.n74 VP.n5 161.3
R189 VP.n73 VP.n72 161.3
R190 VP.n71 VP.n6 161.3
R191 VP.n70 VP.n69 161.3
R192 VP.n68 VP.n7 161.3
R193 VP.n67 VP.n66 161.3
R194 VP.n65 VP.n8 161.3
R195 VP.n64 VP.n63 161.3
R196 VP.n61 VP.n9 161.3
R197 VP.n60 VP.n59 161.3
R198 VP.n58 VP.n10 161.3
R199 VP.n57 VP.n56 161.3
R200 VP.n55 VP.n11 161.3
R201 VP.n54 VP.n53 161.3
R202 VP.n52 VP.n12 161.3
R203 VP.n51 VP.n50 79.9102
R204 VP.n90 VP.n0 79.9102
R205 VP.n49 VP.n13 79.9102
R206 VP.n23 VP.n22 62.9336
R207 VP.n56 VP.n10 56.4773
R208 VP.n69 VP.n6 56.4773
R209 VP.n82 VP.n2 56.4773
R210 VP.n41 VP.n15 56.4773
R211 VP.n28 VP.n19 56.4773
R212 VP.n51 VP.n49 47.9461
R213 VP.n23 VP.t1 43.3813
R214 VP.n54 VP.n12 24.3439
R215 VP.n55 VP.n54 24.3439
R216 VP.n56 VP.n55 24.3439
R217 VP.n60 VP.n10 24.3439
R218 VP.n61 VP.n60 24.3439
R219 VP.n63 VP.n61 24.3439
R220 VP.n67 VP.n8 24.3439
R221 VP.n68 VP.n67 24.3439
R222 VP.n69 VP.n68 24.3439
R223 VP.n73 VP.n6 24.3439
R224 VP.n74 VP.n73 24.3439
R225 VP.n76 VP.n74 24.3439
R226 VP.n80 VP.n4 24.3439
R227 VP.n81 VP.n80 24.3439
R228 VP.n82 VP.n81 24.3439
R229 VP.n86 VP.n2 24.3439
R230 VP.n87 VP.n86 24.3439
R231 VP.n88 VP.n87 24.3439
R232 VP.n45 VP.n15 24.3439
R233 VP.n46 VP.n45 24.3439
R234 VP.n47 VP.n46 24.3439
R235 VP.n32 VP.n19 24.3439
R236 VP.n33 VP.n32 24.3439
R237 VP.n35 VP.n33 24.3439
R238 VP.n39 VP.n17 24.3439
R239 VP.n40 VP.n39 24.3439
R240 VP.n41 VP.n40 24.3439
R241 VP.n26 VP.n21 24.3439
R242 VP.n27 VP.n26 24.3439
R243 VP.n28 VP.n27 24.3439
R244 VP.n63 VP.n62 12.9025
R245 VP.n75 VP.n4 12.9025
R246 VP.n34 VP.n17 12.9025
R247 VP.n62 VP.n8 11.4419
R248 VP.n76 VP.n75 11.4419
R249 VP.n35 VP.n34 11.4419
R250 VP.n22 VP.n21 11.4419
R251 VP.n50 VP.t0 10.0642
R252 VP.n62 VP.t3 10.0642
R253 VP.n75 VP.t6 10.0642
R254 VP.n0 VP.t4 10.0642
R255 VP.n13 VP.t2 10.0642
R256 VP.n34 VP.t7 10.0642
R257 VP.n22 VP.t5 10.0642
R258 VP.n50 VP.n12 9.98131
R259 VP.n88 VP.n0 9.98131
R260 VP.n47 VP.n13 9.98131
R261 VP.n24 VP.n23 3.16877
R262 VP.n49 VP.n48 0.355081
R263 VP.n52 VP.n51 0.355081
R264 VP.n90 VP.n89 0.355081
R265 VP VP.n90 0.26685
R266 VP.n25 VP.n24 0.189894
R267 VP.n25 VP.n20 0.189894
R268 VP.n29 VP.n20 0.189894
R269 VP.n30 VP.n29 0.189894
R270 VP.n31 VP.n30 0.189894
R271 VP.n31 VP.n18 0.189894
R272 VP.n36 VP.n18 0.189894
R273 VP.n37 VP.n36 0.189894
R274 VP.n38 VP.n37 0.189894
R275 VP.n38 VP.n16 0.189894
R276 VP.n42 VP.n16 0.189894
R277 VP.n43 VP.n42 0.189894
R278 VP.n44 VP.n43 0.189894
R279 VP.n44 VP.n14 0.189894
R280 VP.n48 VP.n14 0.189894
R281 VP.n53 VP.n52 0.189894
R282 VP.n53 VP.n11 0.189894
R283 VP.n57 VP.n11 0.189894
R284 VP.n58 VP.n57 0.189894
R285 VP.n59 VP.n58 0.189894
R286 VP.n59 VP.n9 0.189894
R287 VP.n64 VP.n9 0.189894
R288 VP.n65 VP.n64 0.189894
R289 VP.n66 VP.n65 0.189894
R290 VP.n66 VP.n7 0.189894
R291 VP.n70 VP.n7 0.189894
R292 VP.n71 VP.n70 0.189894
R293 VP.n72 VP.n71 0.189894
R294 VP.n72 VP.n5 0.189894
R295 VP.n77 VP.n5 0.189894
R296 VP.n78 VP.n77 0.189894
R297 VP.n79 VP.n78 0.189894
R298 VP.n79 VP.n3 0.189894
R299 VP.n83 VP.n3 0.189894
R300 VP.n84 VP.n83 0.189894
R301 VP.n85 VP.n84 0.189894
R302 VP.n85 VP.n1 0.189894
R303 VP.n89 VP.n1 0.189894
R304 VDD1 VDD1.n0 253.109
R305 VDD1.n3 VDD1.n2 252.996
R306 VDD1.n3 VDD1.n1 252.996
R307 VDD1.n5 VDD1.n4 251.34
R308 VDD1.n5 VDD1.n3 41.0095
R309 VDD1.n4 VDD1.t0 21.3854
R310 VDD1.n4 VDD1.t5 21.3854
R311 VDD1.n0 VDD1.t6 21.3854
R312 VDD1.n0 VDD1.t2 21.3854
R313 VDD1.n2 VDD1.t1 21.3854
R314 VDD1.n2 VDD1.t3 21.3854
R315 VDD1.n1 VDD1.t7 21.3854
R316 VDD1.n1 VDD1.t4 21.3854
R317 VDD1 VDD1.n5 1.65352
R318 B.n320 B.n319 585
R319 B.n318 B.n123 585
R320 B.n317 B.n316 585
R321 B.n315 B.n124 585
R322 B.n314 B.n313 585
R323 B.n312 B.n125 585
R324 B.n311 B.n310 585
R325 B.n309 B.n126 585
R326 B.n308 B.n307 585
R327 B.n306 B.n127 585
R328 B.n305 B.n304 585
R329 B.n302 B.n128 585
R330 B.n301 B.n300 585
R331 B.n299 B.n131 585
R332 B.n298 B.n297 585
R333 B.n296 B.n132 585
R334 B.n295 B.n294 585
R335 B.n293 B.n133 585
R336 B.n292 B.n291 585
R337 B.n290 B.n134 585
R338 B.n288 B.n287 585
R339 B.n286 B.n137 585
R340 B.n285 B.n284 585
R341 B.n283 B.n138 585
R342 B.n282 B.n281 585
R343 B.n280 B.n139 585
R344 B.n279 B.n278 585
R345 B.n277 B.n140 585
R346 B.n276 B.n275 585
R347 B.n274 B.n141 585
R348 B.n273 B.n272 585
R349 B.n321 B.n122 585
R350 B.n323 B.n322 585
R351 B.n324 B.n121 585
R352 B.n326 B.n325 585
R353 B.n327 B.n120 585
R354 B.n329 B.n328 585
R355 B.n330 B.n119 585
R356 B.n332 B.n331 585
R357 B.n333 B.n118 585
R358 B.n335 B.n334 585
R359 B.n336 B.n117 585
R360 B.n338 B.n337 585
R361 B.n339 B.n116 585
R362 B.n341 B.n340 585
R363 B.n342 B.n115 585
R364 B.n344 B.n343 585
R365 B.n345 B.n114 585
R366 B.n347 B.n346 585
R367 B.n348 B.n113 585
R368 B.n350 B.n349 585
R369 B.n351 B.n112 585
R370 B.n353 B.n352 585
R371 B.n354 B.n111 585
R372 B.n356 B.n355 585
R373 B.n357 B.n110 585
R374 B.n359 B.n358 585
R375 B.n360 B.n109 585
R376 B.n362 B.n361 585
R377 B.n363 B.n108 585
R378 B.n365 B.n364 585
R379 B.n366 B.n107 585
R380 B.n368 B.n367 585
R381 B.n369 B.n106 585
R382 B.n371 B.n370 585
R383 B.n372 B.n105 585
R384 B.n374 B.n373 585
R385 B.n375 B.n104 585
R386 B.n377 B.n376 585
R387 B.n378 B.n103 585
R388 B.n380 B.n379 585
R389 B.n381 B.n102 585
R390 B.n383 B.n382 585
R391 B.n384 B.n101 585
R392 B.n386 B.n385 585
R393 B.n387 B.n100 585
R394 B.n389 B.n388 585
R395 B.n390 B.n99 585
R396 B.n392 B.n391 585
R397 B.n393 B.n98 585
R398 B.n395 B.n394 585
R399 B.n396 B.n97 585
R400 B.n398 B.n397 585
R401 B.n399 B.n96 585
R402 B.n401 B.n400 585
R403 B.n402 B.n95 585
R404 B.n404 B.n403 585
R405 B.n405 B.n94 585
R406 B.n407 B.n406 585
R407 B.n408 B.n93 585
R408 B.n410 B.n409 585
R409 B.n411 B.n92 585
R410 B.n413 B.n412 585
R411 B.n414 B.n91 585
R412 B.n416 B.n415 585
R413 B.n417 B.n90 585
R414 B.n419 B.n418 585
R415 B.n420 B.n89 585
R416 B.n422 B.n421 585
R417 B.n423 B.n88 585
R418 B.n425 B.n424 585
R419 B.n426 B.n87 585
R420 B.n428 B.n427 585
R421 B.n429 B.n86 585
R422 B.n431 B.n430 585
R423 B.n432 B.n85 585
R424 B.n434 B.n433 585
R425 B.n435 B.n84 585
R426 B.n437 B.n436 585
R427 B.n438 B.n83 585
R428 B.n440 B.n439 585
R429 B.n441 B.n82 585
R430 B.n443 B.n442 585
R431 B.n444 B.n81 585
R432 B.n446 B.n445 585
R433 B.n447 B.n80 585
R434 B.n449 B.n448 585
R435 B.n450 B.n79 585
R436 B.n452 B.n451 585
R437 B.n453 B.n78 585
R438 B.n455 B.n454 585
R439 B.n456 B.n77 585
R440 B.n458 B.n457 585
R441 B.n459 B.n76 585
R442 B.n461 B.n460 585
R443 B.n462 B.n75 585
R444 B.n464 B.n463 585
R445 B.n465 B.n74 585
R446 B.n467 B.n466 585
R447 B.n468 B.n73 585
R448 B.n470 B.n469 585
R449 B.n471 B.n72 585
R450 B.n473 B.n472 585
R451 B.n474 B.n71 585
R452 B.n476 B.n475 585
R453 B.n477 B.n70 585
R454 B.n479 B.n478 585
R455 B.n480 B.n69 585
R456 B.n482 B.n481 585
R457 B.n483 B.n68 585
R458 B.n485 B.n484 585
R459 B.n486 B.n67 585
R460 B.n488 B.n487 585
R461 B.n489 B.n66 585
R462 B.n491 B.n490 585
R463 B.n492 B.n65 585
R464 B.n494 B.n493 585
R465 B.n495 B.n64 585
R466 B.n497 B.n496 585
R467 B.n498 B.n63 585
R468 B.n500 B.n499 585
R469 B.n501 B.n62 585
R470 B.n503 B.n502 585
R471 B.n504 B.n61 585
R472 B.n506 B.n505 585
R473 B.n507 B.n60 585
R474 B.n509 B.n508 585
R475 B.n510 B.n59 585
R476 B.n512 B.n511 585
R477 B.n513 B.n58 585
R478 B.n515 B.n514 585
R479 B.n516 B.n57 585
R480 B.n518 B.n517 585
R481 B.n519 B.n56 585
R482 B.n521 B.n520 585
R483 B.n568 B.n35 585
R484 B.n567 B.n566 585
R485 B.n565 B.n36 585
R486 B.n564 B.n563 585
R487 B.n562 B.n37 585
R488 B.n561 B.n560 585
R489 B.n559 B.n38 585
R490 B.n558 B.n557 585
R491 B.n556 B.n39 585
R492 B.n555 B.n554 585
R493 B.n553 B.n40 585
R494 B.n552 B.n551 585
R495 B.n550 B.n41 585
R496 B.n549 B.n548 585
R497 B.n547 B.n45 585
R498 B.n546 B.n545 585
R499 B.n544 B.n46 585
R500 B.n543 B.n542 585
R501 B.n541 B.n47 585
R502 B.n540 B.n539 585
R503 B.n537 B.n48 585
R504 B.n536 B.n535 585
R505 B.n534 B.n51 585
R506 B.n533 B.n532 585
R507 B.n531 B.n52 585
R508 B.n530 B.n529 585
R509 B.n528 B.n53 585
R510 B.n527 B.n526 585
R511 B.n525 B.n54 585
R512 B.n524 B.n523 585
R513 B.n522 B.n55 585
R514 B.n570 B.n569 585
R515 B.n571 B.n34 585
R516 B.n573 B.n572 585
R517 B.n574 B.n33 585
R518 B.n576 B.n575 585
R519 B.n577 B.n32 585
R520 B.n579 B.n578 585
R521 B.n580 B.n31 585
R522 B.n582 B.n581 585
R523 B.n583 B.n30 585
R524 B.n585 B.n584 585
R525 B.n586 B.n29 585
R526 B.n588 B.n587 585
R527 B.n589 B.n28 585
R528 B.n591 B.n590 585
R529 B.n592 B.n27 585
R530 B.n594 B.n593 585
R531 B.n595 B.n26 585
R532 B.n597 B.n596 585
R533 B.n598 B.n25 585
R534 B.n600 B.n599 585
R535 B.n601 B.n24 585
R536 B.n603 B.n602 585
R537 B.n604 B.n23 585
R538 B.n606 B.n605 585
R539 B.n607 B.n22 585
R540 B.n609 B.n608 585
R541 B.n610 B.n21 585
R542 B.n612 B.n611 585
R543 B.n613 B.n20 585
R544 B.n615 B.n614 585
R545 B.n616 B.n19 585
R546 B.n618 B.n617 585
R547 B.n619 B.n18 585
R548 B.n621 B.n620 585
R549 B.n622 B.n17 585
R550 B.n624 B.n623 585
R551 B.n625 B.n16 585
R552 B.n627 B.n626 585
R553 B.n628 B.n15 585
R554 B.n630 B.n629 585
R555 B.n631 B.n14 585
R556 B.n633 B.n632 585
R557 B.n634 B.n13 585
R558 B.n636 B.n635 585
R559 B.n637 B.n12 585
R560 B.n639 B.n638 585
R561 B.n640 B.n11 585
R562 B.n642 B.n641 585
R563 B.n643 B.n10 585
R564 B.n645 B.n644 585
R565 B.n646 B.n9 585
R566 B.n648 B.n647 585
R567 B.n649 B.n8 585
R568 B.n651 B.n650 585
R569 B.n652 B.n7 585
R570 B.n654 B.n653 585
R571 B.n655 B.n6 585
R572 B.n657 B.n656 585
R573 B.n658 B.n5 585
R574 B.n660 B.n659 585
R575 B.n661 B.n4 585
R576 B.n663 B.n662 585
R577 B.n664 B.n3 585
R578 B.n666 B.n665 585
R579 B.n667 B.n0 585
R580 B.n2 B.n1 585
R581 B.n175 B.n174 585
R582 B.n177 B.n176 585
R583 B.n178 B.n173 585
R584 B.n180 B.n179 585
R585 B.n181 B.n172 585
R586 B.n183 B.n182 585
R587 B.n184 B.n171 585
R588 B.n186 B.n185 585
R589 B.n187 B.n170 585
R590 B.n189 B.n188 585
R591 B.n190 B.n169 585
R592 B.n192 B.n191 585
R593 B.n193 B.n168 585
R594 B.n195 B.n194 585
R595 B.n196 B.n167 585
R596 B.n198 B.n197 585
R597 B.n199 B.n166 585
R598 B.n201 B.n200 585
R599 B.n202 B.n165 585
R600 B.n204 B.n203 585
R601 B.n205 B.n164 585
R602 B.n207 B.n206 585
R603 B.n208 B.n163 585
R604 B.n210 B.n209 585
R605 B.n211 B.n162 585
R606 B.n213 B.n212 585
R607 B.n214 B.n161 585
R608 B.n216 B.n215 585
R609 B.n217 B.n160 585
R610 B.n219 B.n218 585
R611 B.n220 B.n159 585
R612 B.n222 B.n221 585
R613 B.n223 B.n158 585
R614 B.n225 B.n224 585
R615 B.n226 B.n157 585
R616 B.n228 B.n227 585
R617 B.n229 B.n156 585
R618 B.n231 B.n230 585
R619 B.n232 B.n155 585
R620 B.n234 B.n233 585
R621 B.n235 B.n154 585
R622 B.n237 B.n236 585
R623 B.n238 B.n153 585
R624 B.n240 B.n239 585
R625 B.n241 B.n152 585
R626 B.n243 B.n242 585
R627 B.n244 B.n151 585
R628 B.n246 B.n245 585
R629 B.n247 B.n150 585
R630 B.n249 B.n248 585
R631 B.n250 B.n149 585
R632 B.n252 B.n251 585
R633 B.n253 B.n148 585
R634 B.n255 B.n254 585
R635 B.n256 B.n147 585
R636 B.n258 B.n257 585
R637 B.n259 B.n146 585
R638 B.n261 B.n260 585
R639 B.n262 B.n145 585
R640 B.n264 B.n263 585
R641 B.n265 B.n144 585
R642 B.n267 B.n266 585
R643 B.n268 B.n143 585
R644 B.n270 B.n269 585
R645 B.n271 B.n142 585
R646 B.n273 B.n142 511.721
R647 B.n319 B.n122 511.721
R648 B.n522 B.n521 511.721
R649 B.n570 B.n35 511.721
R650 B.n129 B.t4 326.545
R651 B.n49 B.t8 326.545
R652 B.n135 B.t10 326.543
R653 B.n42 B.t2 326.543
R654 B.n669 B.n668 256.663
R655 B.n130 B.t5 249.55
R656 B.n50 B.t7 249.55
R657 B.n136 B.t11 249.549
R658 B.n43 B.t1 249.549
R659 B.n668 B.n667 235.042
R660 B.n668 B.n2 235.042
R661 B.n135 B.t9 209.685
R662 B.n129 B.t3 209.685
R663 B.n49 B.t6 209.685
R664 B.n42 B.t0 209.685
R665 B.n274 B.n273 163.367
R666 B.n275 B.n274 163.367
R667 B.n275 B.n140 163.367
R668 B.n279 B.n140 163.367
R669 B.n280 B.n279 163.367
R670 B.n281 B.n280 163.367
R671 B.n281 B.n138 163.367
R672 B.n285 B.n138 163.367
R673 B.n286 B.n285 163.367
R674 B.n287 B.n286 163.367
R675 B.n287 B.n134 163.367
R676 B.n292 B.n134 163.367
R677 B.n293 B.n292 163.367
R678 B.n294 B.n293 163.367
R679 B.n294 B.n132 163.367
R680 B.n298 B.n132 163.367
R681 B.n299 B.n298 163.367
R682 B.n300 B.n299 163.367
R683 B.n300 B.n128 163.367
R684 B.n305 B.n128 163.367
R685 B.n306 B.n305 163.367
R686 B.n307 B.n306 163.367
R687 B.n307 B.n126 163.367
R688 B.n311 B.n126 163.367
R689 B.n312 B.n311 163.367
R690 B.n313 B.n312 163.367
R691 B.n313 B.n124 163.367
R692 B.n317 B.n124 163.367
R693 B.n318 B.n317 163.367
R694 B.n319 B.n318 163.367
R695 B.n521 B.n56 163.367
R696 B.n517 B.n56 163.367
R697 B.n517 B.n516 163.367
R698 B.n516 B.n515 163.367
R699 B.n515 B.n58 163.367
R700 B.n511 B.n58 163.367
R701 B.n511 B.n510 163.367
R702 B.n510 B.n509 163.367
R703 B.n509 B.n60 163.367
R704 B.n505 B.n60 163.367
R705 B.n505 B.n504 163.367
R706 B.n504 B.n503 163.367
R707 B.n503 B.n62 163.367
R708 B.n499 B.n62 163.367
R709 B.n499 B.n498 163.367
R710 B.n498 B.n497 163.367
R711 B.n497 B.n64 163.367
R712 B.n493 B.n64 163.367
R713 B.n493 B.n492 163.367
R714 B.n492 B.n491 163.367
R715 B.n491 B.n66 163.367
R716 B.n487 B.n66 163.367
R717 B.n487 B.n486 163.367
R718 B.n486 B.n485 163.367
R719 B.n485 B.n68 163.367
R720 B.n481 B.n68 163.367
R721 B.n481 B.n480 163.367
R722 B.n480 B.n479 163.367
R723 B.n479 B.n70 163.367
R724 B.n475 B.n70 163.367
R725 B.n475 B.n474 163.367
R726 B.n474 B.n473 163.367
R727 B.n473 B.n72 163.367
R728 B.n469 B.n72 163.367
R729 B.n469 B.n468 163.367
R730 B.n468 B.n467 163.367
R731 B.n467 B.n74 163.367
R732 B.n463 B.n74 163.367
R733 B.n463 B.n462 163.367
R734 B.n462 B.n461 163.367
R735 B.n461 B.n76 163.367
R736 B.n457 B.n76 163.367
R737 B.n457 B.n456 163.367
R738 B.n456 B.n455 163.367
R739 B.n455 B.n78 163.367
R740 B.n451 B.n78 163.367
R741 B.n451 B.n450 163.367
R742 B.n450 B.n449 163.367
R743 B.n449 B.n80 163.367
R744 B.n445 B.n80 163.367
R745 B.n445 B.n444 163.367
R746 B.n444 B.n443 163.367
R747 B.n443 B.n82 163.367
R748 B.n439 B.n82 163.367
R749 B.n439 B.n438 163.367
R750 B.n438 B.n437 163.367
R751 B.n437 B.n84 163.367
R752 B.n433 B.n84 163.367
R753 B.n433 B.n432 163.367
R754 B.n432 B.n431 163.367
R755 B.n431 B.n86 163.367
R756 B.n427 B.n86 163.367
R757 B.n427 B.n426 163.367
R758 B.n426 B.n425 163.367
R759 B.n425 B.n88 163.367
R760 B.n421 B.n88 163.367
R761 B.n421 B.n420 163.367
R762 B.n420 B.n419 163.367
R763 B.n419 B.n90 163.367
R764 B.n415 B.n90 163.367
R765 B.n415 B.n414 163.367
R766 B.n414 B.n413 163.367
R767 B.n413 B.n92 163.367
R768 B.n409 B.n92 163.367
R769 B.n409 B.n408 163.367
R770 B.n408 B.n407 163.367
R771 B.n407 B.n94 163.367
R772 B.n403 B.n94 163.367
R773 B.n403 B.n402 163.367
R774 B.n402 B.n401 163.367
R775 B.n401 B.n96 163.367
R776 B.n397 B.n96 163.367
R777 B.n397 B.n396 163.367
R778 B.n396 B.n395 163.367
R779 B.n395 B.n98 163.367
R780 B.n391 B.n98 163.367
R781 B.n391 B.n390 163.367
R782 B.n390 B.n389 163.367
R783 B.n389 B.n100 163.367
R784 B.n385 B.n100 163.367
R785 B.n385 B.n384 163.367
R786 B.n384 B.n383 163.367
R787 B.n383 B.n102 163.367
R788 B.n379 B.n102 163.367
R789 B.n379 B.n378 163.367
R790 B.n378 B.n377 163.367
R791 B.n377 B.n104 163.367
R792 B.n373 B.n104 163.367
R793 B.n373 B.n372 163.367
R794 B.n372 B.n371 163.367
R795 B.n371 B.n106 163.367
R796 B.n367 B.n106 163.367
R797 B.n367 B.n366 163.367
R798 B.n366 B.n365 163.367
R799 B.n365 B.n108 163.367
R800 B.n361 B.n108 163.367
R801 B.n361 B.n360 163.367
R802 B.n360 B.n359 163.367
R803 B.n359 B.n110 163.367
R804 B.n355 B.n110 163.367
R805 B.n355 B.n354 163.367
R806 B.n354 B.n353 163.367
R807 B.n353 B.n112 163.367
R808 B.n349 B.n112 163.367
R809 B.n349 B.n348 163.367
R810 B.n348 B.n347 163.367
R811 B.n347 B.n114 163.367
R812 B.n343 B.n114 163.367
R813 B.n343 B.n342 163.367
R814 B.n342 B.n341 163.367
R815 B.n341 B.n116 163.367
R816 B.n337 B.n116 163.367
R817 B.n337 B.n336 163.367
R818 B.n336 B.n335 163.367
R819 B.n335 B.n118 163.367
R820 B.n331 B.n118 163.367
R821 B.n331 B.n330 163.367
R822 B.n330 B.n329 163.367
R823 B.n329 B.n120 163.367
R824 B.n325 B.n120 163.367
R825 B.n325 B.n324 163.367
R826 B.n324 B.n323 163.367
R827 B.n323 B.n122 163.367
R828 B.n566 B.n35 163.367
R829 B.n566 B.n565 163.367
R830 B.n565 B.n564 163.367
R831 B.n564 B.n37 163.367
R832 B.n560 B.n37 163.367
R833 B.n560 B.n559 163.367
R834 B.n559 B.n558 163.367
R835 B.n558 B.n39 163.367
R836 B.n554 B.n39 163.367
R837 B.n554 B.n553 163.367
R838 B.n553 B.n552 163.367
R839 B.n552 B.n41 163.367
R840 B.n548 B.n41 163.367
R841 B.n548 B.n547 163.367
R842 B.n547 B.n546 163.367
R843 B.n546 B.n46 163.367
R844 B.n542 B.n46 163.367
R845 B.n542 B.n541 163.367
R846 B.n541 B.n540 163.367
R847 B.n540 B.n48 163.367
R848 B.n535 B.n48 163.367
R849 B.n535 B.n534 163.367
R850 B.n534 B.n533 163.367
R851 B.n533 B.n52 163.367
R852 B.n529 B.n52 163.367
R853 B.n529 B.n528 163.367
R854 B.n528 B.n527 163.367
R855 B.n527 B.n54 163.367
R856 B.n523 B.n54 163.367
R857 B.n523 B.n522 163.367
R858 B.n571 B.n570 163.367
R859 B.n572 B.n571 163.367
R860 B.n572 B.n33 163.367
R861 B.n576 B.n33 163.367
R862 B.n577 B.n576 163.367
R863 B.n578 B.n577 163.367
R864 B.n578 B.n31 163.367
R865 B.n582 B.n31 163.367
R866 B.n583 B.n582 163.367
R867 B.n584 B.n583 163.367
R868 B.n584 B.n29 163.367
R869 B.n588 B.n29 163.367
R870 B.n589 B.n588 163.367
R871 B.n590 B.n589 163.367
R872 B.n590 B.n27 163.367
R873 B.n594 B.n27 163.367
R874 B.n595 B.n594 163.367
R875 B.n596 B.n595 163.367
R876 B.n596 B.n25 163.367
R877 B.n600 B.n25 163.367
R878 B.n601 B.n600 163.367
R879 B.n602 B.n601 163.367
R880 B.n602 B.n23 163.367
R881 B.n606 B.n23 163.367
R882 B.n607 B.n606 163.367
R883 B.n608 B.n607 163.367
R884 B.n608 B.n21 163.367
R885 B.n612 B.n21 163.367
R886 B.n613 B.n612 163.367
R887 B.n614 B.n613 163.367
R888 B.n614 B.n19 163.367
R889 B.n618 B.n19 163.367
R890 B.n619 B.n618 163.367
R891 B.n620 B.n619 163.367
R892 B.n620 B.n17 163.367
R893 B.n624 B.n17 163.367
R894 B.n625 B.n624 163.367
R895 B.n626 B.n625 163.367
R896 B.n626 B.n15 163.367
R897 B.n630 B.n15 163.367
R898 B.n631 B.n630 163.367
R899 B.n632 B.n631 163.367
R900 B.n632 B.n13 163.367
R901 B.n636 B.n13 163.367
R902 B.n637 B.n636 163.367
R903 B.n638 B.n637 163.367
R904 B.n638 B.n11 163.367
R905 B.n642 B.n11 163.367
R906 B.n643 B.n642 163.367
R907 B.n644 B.n643 163.367
R908 B.n644 B.n9 163.367
R909 B.n648 B.n9 163.367
R910 B.n649 B.n648 163.367
R911 B.n650 B.n649 163.367
R912 B.n650 B.n7 163.367
R913 B.n654 B.n7 163.367
R914 B.n655 B.n654 163.367
R915 B.n656 B.n655 163.367
R916 B.n656 B.n5 163.367
R917 B.n660 B.n5 163.367
R918 B.n661 B.n660 163.367
R919 B.n662 B.n661 163.367
R920 B.n662 B.n3 163.367
R921 B.n666 B.n3 163.367
R922 B.n667 B.n666 163.367
R923 B.n174 B.n2 163.367
R924 B.n177 B.n174 163.367
R925 B.n178 B.n177 163.367
R926 B.n179 B.n178 163.367
R927 B.n179 B.n172 163.367
R928 B.n183 B.n172 163.367
R929 B.n184 B.n183 163.367
R930 B.n185 B.n184 163.367
R931 B.n185 B.n170 163.367
R932 B.n189 B.n170 163.367
R933 B.n190 B.n189 163.367
R934 B.n191 B.n190 163.367
R935 B.n191 B.n168 163.367
R936 B.n195 B.n168 163.367
R937 B.n196 B.n195 163.367
R938 B.n197 B.n196 163.367
R939 B.n197 B.n166 163.367
R940 B.n201 B.n166 163.367
R941 B.n202 B.n201 163.367
R942 B.n203 B.n202 163.367
R943 B.n203 B.n164 163.367
R944 B.n207 B.n164 163.367
R945 B.n208 B.n207 163.367
R946 B.n209 B.n208 163.367
R947 B.n209 B.n162 163.367
R948 B.n213 B.n162 163.367
R949 B.n214 B.n213 163.367
R950 B.n215 B.n214 163.367
R951 B.n215 B.n160 163.367
R952 B.n219 B.n160 163.367
R953 B.n220 B.n219 163.367
R954 B.n221 B.n220 163.367
R955 B.n221 B.n158 163.367
R956 B.n225 B.n158 163.367
R957 B.n226 B.n225 163.367
R958 B.n227 B.n226 163.367
R959 B.n227 B.n156 163.367
R960 B.n231 B.n156 163.367
R961 B.n232 B.n231 163.367
R962 B.n233 B.n232 163.367
R963 B.n233 B.n154 163.367
R964 B.n237 B.n154 163.367
R965 B.n238 B.n237 163.367
R966 B.n239 B.n238 163.367
R967 B.n239 B.n152 163.367
R968 B.n243 B.n152 163.367
R969 B.n244 B.n243 163.367
R970 B.n245 B.n244 163.367
R971 B.n245 B.n150 163.367
R972 B.n249 B.n150 163.367
R973 B.n250 B.n249 163.367
R974 B.n251 B.n250 163.367
R975 B.n251 B.n148 163.367
R976 B.n255 B.n148 163.367
R977 B.n256 B.n255 163.367
R978 B.n257 B.n256 163.367
R979 B.n257 B.n146 163.367
R980 B.n261 B.n146 163.367
R981 B.n262 B.n261 163.367
R982 B.n263 B.n262 163.367
R983 B.n263 B.n144 163.367
R984 B.n267 B.n144 163.367
R985 B.n268 B.n267 163.367
R986 B.n269 B.n268 163.367
R987 B.n269 B.n142 163.367
R988 B.n136 B.n135 76.9944
R989 B.n130 B.n129 76.9944
R990 B.n50 B.n49 76.9944
R991 B.n43 B.n42 76.9944
R992 B.n289 B.n136 59.5399
R993 B.n303 B.n130 59.5399
R994 B.n538 B.n50 59.5399
R995 B.n44 B.n43 59.5399
R996 B.n569 B.n568 33.2493
R997 B.n520 B.n55 33.2493
R998 B.n321 B.n320 33.2493
R999 B.n272 B.n271 33.2493
R1000 B B.n669 18.0485
R1001 B.n569 B.n34 10.6151
R1002 B.n573 B.n34 10.6151
R1003 B.n574 B.n573 10.6151
R1004 B.n575 B.n574 10.6151
R1005 B.n575 B.n32 10.6151
R1006 B.n579 B.n32 10.6151
R1007 B.n580 B.n579 10.6151
R1008 B.n581 B.n580 10.6151
R1009 B.n581 B.n30 10.6151
R1010 B.n585 B.n30 10.6151
R1011 B.n586 B.n585 10.6151
R1012 B.n587 B.n586 10.6151
R1013 B.n587 B.n28 10.6151
R1014 B.n591 B.n28 10.6151
R1015 B.n592 B.n591 10.6151
R1016 B.n593 B.n592 10.6151
R1017 B.n593 B.n26 10.6151
R1018 B.n597 B.n26 10.6151
R1019 B.n598 B.n597 10.6151
R1020 B.n599 B.n598 10.6151
R1021 B.n599 B.n24 10.6151
R1022 B.n603 B.n24 10.6151
R1023 B.n604 B.n603 10.6151
R1024 B.n605 B.n604 10.6151
R1025 B.n605 B.n22 10.6151
R1026 B.n609 B.n22 10.6151
R1027 B.n610 B.n609 10.6151
R1028 B.n611 B.n610 10.6151
R1029 B.n611 B.n20 10.6151
R1030 B.n615 B.n20 10.6151
R1031 B.n616 B.n615 10.6151
R1032 B.n617 B.n616 10.6151
R1033 B.n617 B.n18 10.6151
R1034 B.n621 B.n18 10.6151
R1035 B.n622 B.n621 10.6151
R1036 B.n623 B.n622 10.6151
R1037 B.n623 B.n16 10.6151
R1038 B.n627 B.n16 10.6151
R1039 B.n628 B.n627 10.6151
R1040 B.n629 B.n628 10.6151
R1041 B.n629 B.n14 10.6151
R1042 B.n633 B.n14 10.6151
R1043 B.n634 B.n633 10.6151
R1044 B.n635 B.n634 10.6151
R1045 B.n635 B.n12 10.6151
R1046 B.n639 B.n12 10.6151
R1047 B.n640 B.n639 10.6151
R1048 B.n641 B.n640 10.6151
R1049 B.n641 B.n10 10.6151
R1050 B.n645 B.n10 10.6151
R1051 B.n646 B.n645 10.6151
R1052 B.n647 B.n646 10.6151
R1053 B.n647 B.n8 10.6151
R1054 B.n651 B.n8 10.6151
R1055 B.n652 B.n651 10.6151
R1056 B.n653 B.n652 10.6151
R1057 B.n653 B.n6 10.6151
R1058 B.n657 B.n6 10.6151
R1059 B.n658 B.n657 10.6151
R1060 B.n659 B.n658 10.6151
R1061 B.n659 B.n4 10.6151
R1062 B.n663 B.n4 10.6151
R1063 B.n664 B.n663 10.6151
R1064 B.n665 B.n664 10.6151
R1065 B.n665 B.n0 10.6151
R1066 B.n568 B.n567 10.6151
R1067 B.n567 B.n36 10.6151
R1068 B.n563 B.n36 10.6151
R1069 B.n563 B.n562 10.6151
R1070 B.n562 B.n561 10.6151
R1071 B.n561 B.n38 10.6151
R1072 B.n557 B.n38 10.6151
R1073 B.n557 B.n556 10.6151
R1074 B.n556 B.n555 10.6151
R1075 B.n555 B.n40 10.6151
R1076 B.n551 B.n550 10.6151
R1077 B.n550 B.n549 10.6151
R1078 B.n549 B.n45 10.6151
R1079 B.n545 B.n45 10.6151
R1080 B.n545 B.n544 10.6151
R1081 B.n544 B.n543 10.6151
R1082 B.n543 B.n47 10.6151
R1083 B.n539 B.n47 10.6151
R1084 B.n537 B.n536 10.6151
R1085 B.n536 B.n51 10.6151
R1086 B.n532 B.n51 10.6151
R1087 B.n532 B.n531 10.6151
R1088 B.n531 B.n530 10.6151
R1089 B.n530 B.n53 10.6151
R1090 B.n526 B.n53 10.6151
R1091 B.n526 B.n525 10.6151
R1092 B.n525 B.n524 10.6151
R1093 B.n524 B.n55 10.6151
R1094 B.n520 B.n519 10.6151
R1095 B.n519 B.n518 10.6151
R1096 B.n518 B.n57 10.6151
R1097 B.n514 B.n57 10.6151
R1098 B.n514 B.n513 10.6151
R1099 B.n513 B.n512 10.6151
R1100 B.n512 B.n59 10.6151
R1101 B.n508 B.n59 10.6151
R1102 B.n508 B.n507 10.6151
R1103 B.n507 B.n506 10.6151
R1104 B.n506 B.n61 10.6151
R1105 B.n502 B.n61 10.6151
R1106 B.n502 B.n501 10.6151
R1107 B.n501 B.n500 10.6151
R1108 B.n500 B.n63 10.6151
R1109 B.n496 B.n63 10.6151
R1110 B.n496 B.n495 10.6151
R1111 B.n495 B.n494 10.6151
R1112 B.n494 B.n65 10.6151
R1113 B.n490 B.n65 10.6151
R1114 B.n490 B.n489 10.6151
R1115 B.n489 B.n488 10.6151
R1116 B.n488 B.n67 10.6151
R1117 B.n484 B.n67 10.6151
R1118 B.n484 B.n483 10.6151
R1119 B.n483 B.n482 10.6151
R1120 B.n482 B.n69 10.6151
R1121 B.n478 B.n69 10.6151
R1122 B.n478 B.n477 10.6151
R1123 B.n477 B.n476 10.6151
R1124 B.n476 B.n71 10.6151
R1125 B.n472 B.n71 10.6151
R1126 B.n472 B.n471 10.6151
R1127 B.n471 B.n470 10.6151
R1128 B.n470 B.n73 10.6151
R1129 B.n466 B.n73 10.6151
R1130 B.n466 B.n465 10.6151
R1131 B.n465 B.n464 10.6151
R1132 B.n464 B.n75 10.6151
R1133 B.n460 B.n75 10.6151
R1134 B.n460 B.n459 10.6151
R1135 B.n459 B.n458 10.6151
R1136 B.n458 B.n77 10.6151
R1137 B.n454 B.n77 10.6151
R1138 B.n454 B.n453 10.6151
R1139 B.n453 B.n452 10.6151
R1140 B.n452 B.n79 10.6151
R1141 B.n448 B.n79 10.6151
R1142 B.n448 B.n447 10.6151
R1143 B.n447 B.n446 10.6151
R1144 B.n446 B.n81 10.6151
R1145 B.n442 B.n81 10.6151
R1146 B.n442 B.n441 10.6151
R1147 B.n441 B.n440 10.6151
R1148 B.n440 B.n83 10.6151
R1149 B.n436 B.n83 10.6151
R1150 B.n436 B.n435 10.6151
R1151 B.n435 B.n434 10.6151
R1152 B.n434 B.n85 10.6151
R1153 B.n430 B.n85 10.6151
R1154 B.n430 B.n429 10.6151
R1155 B.n429 B.n428 10.6151
R1156 B.n428 B.n87 10.6151
R1157 B.n424 B.n87 10.6151
R1158 B.n424 B.n423 10.6151
R1159 B.n423 B.n422 10.6151
R1160 B.n422 B.n89 10.6151
R1161 B.n418 B.n89 10.6151
R1162 B.n418 B.n417 10.6151
R1163 B.n417 B.n416 10.6151
R1164 B.n416 B.n91 10.6151
R1165 B.n412 B.n91 10.6151
R1166 B.n412 B.n411 10.6151
R1167 B.n411 B.n410 10.6151
R1168 B.n410 B.n93 10.6151
R1169 B.n406 B.n93 10.6151
R1170 B.n406 B.n405 10.6151
R1171 B.n405 B.n404 10.6151
R1172 B.n404 B.n95 10.6151
R1173 B.n400 B.n95 10.6151
R1174 B.n400 B.n399 10.6151
R1175 B.n399 B.n398 10.6151
R1176 B.n398 B.n97 10.6151
R1177 B.n394 B.n97 10.6151
R1178 B.n394 B.n393 10.6151
R1179 B.n393 B.n392 10.6151
R1180 B.n392 B.n99 10.6151
R1181 B.n388 B.n99 10.6151
R1182 B.n388 B.n387 10.6151
R1183 B.n387 B.n386 10.6151
R1184 B.n386 B.n101 10.6151
R1185 B.n382 B.n101 10.6151
R1186 B.n382 B.n381 10.6151
R1187 B.n381 B.n380 10.6151
R1188 B.n380 B.n103 10.6151
R1189 B.n376 B.n103 10.6151
R1190 B.n376 B.n375 10.6151
R1191 B.n375 B.n374 10.6151
R1192 B.n374 B.n105 10.6151
R1193 B.n370 B.n105 10.6151
R1194 B.n370 B.n369 10.6151
R1195 B.n369 B.n368 10.6151
R1196 B.n368 B.n107 10.6151
R1197 B.n364 B.n107 10.6151
R1198 B.n364 B.n363 10.6151
R1199 B.n363 B.n362 10.6151
R1200 B.n362 B.n109 10.6151
R1201 B.n358 B.n109 10.6151
R1202 B.n358 B.n357 10.6151
R1203 B.n357 B.n356 10.6151
R1204 B.n356 B.n111 10.6151
R1205 B.n352 B.n111 10.6151
R1206 B.n352 B.n351 10.6151
R1207 B.n351 B.n350 10.6151
R1208 B.n350 B.n113 10.6151
R1209 B.n346 B.n113 10.6151
R1210 B.n346 B.n345 10.6151
R1211 B.n345 B.n344 10.6151
R1212 B.n344 B.n115 10.6151
R1213 B.n340 B.n115 10.6151
R1214 B.n340 B.n339 10.6151
R1215 B.n339 B.n338 10.6151
R1216 B.n338 B.n117 10.6151
R1217 B.n334 B.n117 10.6151
R1218 B.n334 B.n333 10.6151
R1219 B.n333 B.n332 10.6151
R1220 B.n332 B.n119 10.6151
R1221 B.n328 B.n119 10.6151
R1222 B.n328 B.n327 10.6151
R1223 B.n327 B.n326 10.6151
R1224 B.n326 B.n121 10.6151
R1225 B.n322 B.n121 10.6151
R1226 B.n322 B.n321 10.6151
R1227 B.n175 B.n1 10.6151
R1228 B.n176 B.n175 10.6151
R1229 B.n176 B.n173 10.6151
R1230 B.n180 B.n173 10.6151
R1231 B.n181 B.n180 10.6151
R1232 B.n182 B.n181 10.6151
R1233 B.n182 B.n171 10.6151
R1234 B.n186 B.n171 10.6151
R1235 B.n187 B.n186 10.6151
R1236 B.n188 B.n187 10.6151
R1237 B.n188 B.n169 10.6151
R1238 B.n192 B.n169 10.6151
R1239 B.n193 B.n192 10.6151
R1240 B.n194 B.n193 10.6151
R1241 B.n194 B.n167 10.6151
R1242 B.n198 B.n167 10.6151
R1243 B.n199 B.n198 10.6151
R1244 B.n200 B.n199 10.6151
R1245 B.n200 B.n165 10.6151
R1246 B.n204 B.n165 10.6151
R1247 B.n205 B.n204 10.6151
R1248 B.n206 B.n205 10.6151
R1249 B.n206 B.n163 10.6151
R1250 B.n210 B.n163 10.6151
R1251 B.n211 B.n210 10.6151
R1252 B.n212 B.n211 10.6151
R1253 B.n212 B.n161 10.6151
R1254 B.n216 B.n161 10.6151
R1255 B.n217 B.n216 10.6151
R1256 B.n218 B.n217 10.6151
R1257 B.n218 B.n159 10.6151
R1258 B.n222 B.n159 10.6151
R1259 B.n223 B.n222 10.6151
R1260 B.n224 B.n223 10.6151
R1261 B.n224 B.n157 10.6151
R1262 B.n228 B.n157 10.6151
R1263 B.n229 B.n228 10.6151
R1264 B.n230 B.n229 10.6151
R1265 B.n230 B.n155 10.6151
R1266 B.n234 B.n155 10.6151
R1267 B.n235 B.n234 10.6151
R1268 B.n236 B.n235 10.6151
R1269 B.n236 B.n153 10.6151
R1270 B.n240 B.n153 10.6151
R1271 B.n241 B.n240 10.6151
R1272 B.n242 B.n241 10.6151
R1273 B.n242 B.n151 10.6151
R1274 B.n246 B.n151 10.6151
R1275 B.n247 B.n246 10.6151
R1276 B.n248 B.n247 10.6151
R1277 B.n248 B.n149 10.6151
R1278 B.n252 B.n149 10.6151
R1279 B.n253 B.n252 10.6151
R1280 B.n254 B.n253 10.6151
R1281 B.n254 B.n147 10.6151
R1282 B.n258 B.n147 10.6151
R1283 B.n259 B.n258 10.6151
R1284 B.n260 B.n259 10.6151
R1285 B.n260 B.n145 10.6151
R1286 B.n264 B.n145 10.6151
R1287 B.n265 B.n264 10.6151
R1288 B.n266 B.n265 10.6151
R1289 B.n266 B.n143 10.6151
R1290 B.n270 B.n143 10.6151
R1291 B.n271 B.n270 10.6151
R1292 B.n272 B.n141 10.6151
R1293 B.n276 B.n141 10.6151
R1294 B.n277 B.n276 10.6151
R1295 B.n278 B.n277 10.6151
R1296 B.n278 B.n139 10.6151
R1297 B.n282 B.n139 10.6151
R1298 B.n283 B.n282 10.6151
R1299 B.n284 B.n283 10.6151
R1300 B.n284 B.n137 10.6151
R1301 B.n288 B.n137 10.6151
R1302 B.n291 B.n290 10.6151
R1303 B.n291 B.n133 10.6151
R1304 B.n295 B.n133 10.6151
R1305 B.n296 B.n295 10.6151
R1306 B.n297 B.n296 10.6151
R1307 B.n297 B.n131 10.6151
R1308 B.n301 B.n131 10.6151
R1309 B.n302 B.n301 10.6151
R1310 B.n304 B.n127 10.6151
R1311 B.n308 B.n127 10.6151
R1312 B.n309 B.n308 10.6151
R1313 B.n310 B.n309 10.6151
R1314 B.n310 B.n125 10.6151
R1315 B.n314 B.n125 10.6151
R1316 B.n315 B.n314 10.6151
R1317 B.n316 B.n315 10.6151
R1318 B.n316 B.n123 10.6151
R1319 B.n320 B.n123 10.6151
R1320 B.n669 B.n0 8.11757
R1321 B.n669 B.n1 8.11757
R1322 B.n551 B.n44 6.5566
R1323 B.n539 B.n538 6.5566
R1324 B.n290 B.n289 6.5566
R1325 B.n303 B.n302 6.5566
R1326 B.n44 B.n40 4.05904
R1327 B.n538 B.n537 4.05904
R1328 B.n289 B.n288 4.05904
R1329 B.n304 B.n303 4.05904
C0 VN VP 7.0083f
C1 w_n4940_n1272# B 8.86674f
C2 VDD1 VDD2 2.31779f
C3 VTAIL VN 3.25267f
C4 w_n4940_n1272# VDD2 2.16137f
C5 VN B 1.32612f
C6 VTAIL VP 3.26678f
C7 w_n4940_n1272# VDD1 2.0039f
C8 VP B 2.41091f
C9 VN VDD2 1.58433f
C10 VN VDD1 0.159789f
C11 VTAIL B 1.63519f
C12 VP VDD2 0.638282f
C13 VP VDD1 2.05864f
C14 w_n4940_n1272# VN 10.1965f
C15 VTAIL VDD2 5.60162f
C16 VTAIL VDD1 5.54023f
C17 w_n4940_n1272# VP 10.8348f
C18 B VDD2 1.81349f
C19 B VDD1 1.68415f
C20 w_n4940_n1272# VTAIL 1.964f
C21 VDD2 VSUBS 1.938914f
C22 VDD1 VSUBS 2.97199f
C23 VTAIL VSUBS 0.649044f
C24 VN VSUBS 8.43391f
C25 VP VSUBS 3.981711f
C26 B VSUBS 4.943458f
C27 w_n4940_n1272# VSUBS 80.5615f
C28 B.n0 VSUBS 0.010313f
C29 B.n1 VSUBS 0.010313f
C30 B.n2 VSUBS 0.015252f
C31 B.n3 VSUBS 0.011688f
C32 B.n4 VSUBS 0.011688f
C33 B.n5 VSUBS 0.011688f
C34 B.n6 VSUBS 0.011688f
C35 B.n7 VSUBS 0.011688f
C36 B.n8 VSUBS 0.011688f
C37 B.n9 VSUBS 0.011688f
C38 B.n10 VSUBS 0.011688f
C39 B.n11 VSUBS 0.011688f
C40 B.n12 VSUBS 0.011688f
C41 B.n13 VSUBS 0.011688f
C42 B.n14 VSUBS 0.011688f
C43 B.n15 VSUBS 0.011688f
C44 B.n16 VSUBS 0.011688f
C45 B.n17 VSUBS 0.011688f
C46 B.n18 VSUBS 0.011688f
C47 B.n19 VSUBS 0.011688f
C48 B.n20 VSUBS 0.011688f
C49 B.n21 VSUBS 0.011688f
C50 B.n22 VSUBS 0.011688f
C51 B.n23 VSUBS 0.011688f
C52 B.n24 VSUBS 0.011688f
C53 B.n25 VSUBS 0.011688f
C54 B.n26 VSUBS 0.011688f
C55 B.n27 VSUBS 0.011688f
C56 B.n28 VSUBS 0.011688f
C57 B.n29 VSUBS 0.011688f
C58 B.n30 VSUBS 0.011688f
C59 B.n31 VSUBS 0.011688f
C60 B.n32 VSUBS 0.011688f
C61 B.n33 VSUBS 0.011688f
C62 B.n34 VSUBS 0.011688f
C63 B.n35 VSUBS 0.028219f
C64 B.n36 VSUBS 0.011688f
C65 B.n37 VSUBS 0.011688f
C66 B.n38 VSUBS 0.011688f
C67 B.n39 VSUBS 0.011688f
C68 B.n40 VSUBS 0.008079f
C69 B.n41 VSUBS 0.011688f
C70 B.t1 VSUBS 0.05165f
C71 B.t2 VSUBS 0.07029f
C72 B.t0 VSUBS 0.464296f
C73 B.n42 VSUBS 0.124077f
C74 B.n43 VSUBS 0.095727f
C75 B.n44 VSUBS 0.02708f
C76 B.n45 VSUBS 0.011688f
C77 B.n46 VSUBS 0.011688f
C78 B.n47 VSUBS 0.011688f
C79 B.n48 VSUBS 0.011688f
C80 B.t7 VSUBS 0.05165f
C81 B.t8 VSUBS 0.07029f
C82 B.t6 VSUBS 0.464296f
C83 B.n49 VSUBS 0.124077f
C84 B.n50 VSUBS 0.095727f
C85 B.n51 VSUBS 0.011688f
C86 B.n52 VSUBS 0.011688f
C87 B.n53 VSUBS 0.011688f
C88 B.n54 VSUBS 0.011688f
C89 B.n55 VSUBS 0.028219f
C90 B.n56 VSUBS 0.011688f
C91 B.n57 VSUBS 0.011688f
C92 B.n58 VSUBS 0.011688f
C93 B.n59 VSUBS 0.011688f
C94 B.n60 VSUBS 0.011688f
C95 B.n61 VSUBS 0.011688f
C96 B.n62 VSUBS 0.011688f
C97 B.n63 VSUBS 0.011688f
C98 B.n64 VSUBS 0.011688f
C99 B.n65 VSUBS 0.011688f
C100 B.n66 VSUBS 0.011688f
C101 B.n67 VSUBS 0.011688f
C102 B.n68 VSUBS 0.011688f
C103 B.n69 VSUBS 0.011688f
C104 B.n70 VSUBS 0.011688f
C105 B.n71 VSUBS 0.011688f
C106 B.n72 VSUBS 0.011688f
C107 B.n73 VSUBS 0.011688f
C108 B.n74 VSUBS 0.011688f
C109 B.n75 VSUBS 0.011688f
C110 B.n76 VSUBS 0.011688f
C111 B.n77 VSUBS 0.011688f
C112 B.n78 VSUBS 0.011688f
C113 B.n79 VSUBS 0.011688f
C114 B.n80 VSUBS 0.011688f
C115 B.n81 VSUBS 0.011688f
C116 B.n82 VSUBS 0.011688f
C117 B.n83 VSUBS 0.011688f
C118 B.n84 VSUBS 0.011688f
C119 B.n85 VSUBS 0.011688f
C120 B.n86 VSUBS 0.011688f
C121 B.n87 VSUBS 0.011688f
C122 B.n88 VSUBS 0.011688f
C123 B.n89 VSUBS 0.011688f
C124 B.n90 VSUBS 0.011688f
C125 B.n91 VSUBS 0.011688f
C126 B.n92 VSUBS 0.011688f
C127 B.n93 VSUBS 0.011688f
C128 B.n94 VSUBS 0.011688f
C129 B.n95 VSUBS 0.011688f
C130 B.n96 VSUBS 0.011688f
C131 B.n97 VSUBS 0.011688f
C132 B.n98 VSUBS 0.011688f
C133 B.n99 VSUBS 0.011688f
C134 B.n100 VSUBS 0.011688f
C135 B.n101 VSUBS 0.011688f
C136 B.n102 VSUBS 0.011688f
C137 B.n103 VSUBS 0.011688f
C138 B.n104 VSUBS 0.011688f
C139 B.n105 VSUBS 0.011688f
C140 B.n106 VSUBS 0.011688f
C141 B.n107 VSUBS 0.011688f
C142 B.n108 VSUBS 0.011688f
C143 B.n109 VSUBS 0.011688f
C144 B.n110 VSUBS 0.011688f
C145 B.n111 VSUBS 0.011688f
C146 B.n112 VSUBS 0.011688f
C147 B.n113 VSUBS 0.011688f
C148 B.n114 VSUBS 0.011688f
C149 B.n115 VSUBS 0.011688f
C150 B.n116 VSUBS 0.011688f
C151 B.n117 VSUBS 0.011688f
C152 B.n118 VSUBS 0.011688f
C153 B.n119 VSUBS 0.011688f
C154 B.n120 VSUBS 0.011688f
C155 B.n121 VSUBS 0.011688f
C156 B.n122 VSUBS 0.027128f
C157 B.n123 VSUBS 0.011688f
C158 B.n124 VSUBS 0.011688f
C159 B.n125 VSUBS 0.011688f
C160 B.n126 VSUBS 0.011688f
C161 B.n127 VSUBS 0.011688f
C162 B.n128 VSUBS 0.011688f
C163 B.t5 VSUBS 0.05165f
C164 B.t4 VSUBS 0.07029f
C165 B.t3 VSUBS 0.464296f
C166 B.n129 VSUBS 0.124077f
C167 B.n130 VSUBS 0.095727f
C168 B.n131 VSUBS 0.011688f
C169 B.n132 VSUBS 0.011688f
C170 B.n133 VSUBS 0.011688f
C171 B.n134 VSUBS 0.011688f
C172 B.t11 VSUBS 0.05165f
C173 B.t10 VSUBS 0.07029f
C174 B.t9 VSUBS 0.464296f
C175 B.n135 VSUBS 0.124077f
C176 B.n136 VSUBS 0.095727f
C177 B.n137 VSUBS 0.011688f
C178 B.n138 VSUBS 0.011688f
C179 B.n139 VSUBS 0.011688f
C180 B.n140 VSUBS 0.011688f
C181 B.n141 VSUBS 0.011688f
C182 B.n142 VSUBS 0.027128f
C183 B.n143 VSUBS 0.011688f
C184 B.n144 VSUBS 0.011688f
C185 B.n145 VSUBS 0.011688f
C186 B.n146 VSUBS 0.011688f
C187 B.n147 VSUBS 0.011688f
C188 B.n148 VSUBS 0.011688f
C189 B.n149 VSUBS 0.011688f
C190 B.n150 VSUBS 0.011688f
C191 B.n151 VSUBS 0.011688f
C192 B.n152 VSUBS 0.011688f
C193 B.n153 VSUBS 0.011688f
C194 B.n154 VSUBS 0.011688f
C195 B.n155 VSUBS 0.011688f
C196 B.n156 VSUBS 0.011688f
C197 B.n157 VSUBS 0.011688f
C198 B.n158 VSUBS 0.011688f
C199 B.n159 VSUBS 0.011688f
C200 B.n160 VSUBS 0.011688f
C201 B.n161 VSUBS 0.011688f
C202 B.n162 VSUBS 0.011688f
C203 B.n163 VSUBS 0.011688f
C204 B.n164 VSUBS 0.011688f
C205 B.n165 VSUBS 0.011688f
C206 B.n166 VSUBS 0.011688f
C207 B.n167 VSUBS 0.011688f
C208 B.n168 VSUBS 0.011688f
C209 B.n169 VSUBS 0.011688f
C210 B.n170 VSUBS 0.011688f
C211 B.n171 VSUBS 0.011688f
C212 B.n172 VSUBS 0.011688f
C213 B.n173 VSUBS 0.011688f
C214 B.n174 VSUBS 0.011688f
C215 B.n175 VSUBS 0.011688f
C216 B.n176 VSUBS 0.011688f
C217 B.n177 VSUBS 0.011688f
C218 B.n178 VSUBS 0.011688f
C219 B.n179 VSUBS 0.011688f
C220 B.n180 VSUBS 0.011688f
C221 B.n181 VSUBS 0.011688f
C222 B.n182 VSUBS 0.011688f
C223 B.n183 VSUBS 0.011688f
C224 B.n184 VSUBS 0.011688f
C225 B.n185 VSUBS 0.011688f
C226 B.n186 VSUBS 0.011688f
C227 B.n187 VSUBS 0.011688f
C228 B.n188 VSUBS 0.011688f
C229 B.n189 VSUBS 0.011688f
C230 B.n190 VSUBS 0.011688f
C231 B.n191 VSUBS 0.011688f
C232 B.n192 VSUBS 0.011688f
C233 B.n193 VSUBS 0.011688f
C234 B.n194 VSUBS 0.011688f
C235 B.n195 VSUBS 0.011688f
C236 B.n196 VSUBS 0.011688f
C237 B.n197 VSUBS 0.011688f
C238 B.n198 VSUBS 0.011688f
C239 B.n199 VSUBS 0.011688f
C240 B.n200 VSUBS 0.011688f
C241 B.n201 VSUBS 0.011688f
C242 B.n202 VSUBS 0.011688f
C243 B.n203 VSUBS 0.011688f
C244 B.n204 VSUBS 0.011688f
C245 B.n205 VSUBS 0.011688f
C246 B.n206 VSUBS 0.011688f
C247 B.n207 VSUBS 0.011688f
C248 B.n208 VSUBS 0.011688f
C249 B.n209 VSUBS 0.011688f
C250 B.n210 VSUBS 0.011688f
C251 B.n211 VSUBS 0.011688f
C252 B.n212 VSUBS 0.011688f
C253 B.n213 VSUBS 0.011688f
C254 B.n214 VSUBS 0.011688f
C255 B.n215 VSUBS 0.011688f
C256 B.n216 VSUBS 0.011688f
C257 B.n217 VSUBS 0.011688f
C258 B.n218 VSUBS 0.011688f
C259 B.n219 VSUBS 0.011688f
C260 B.n220 VSUBS 0.011688f
C261 B.n221 VSUBS 0.011688f
C262 B.n222 VSUBS 0.011688f
C263 B.n223 VSUBS 0.011688f
C264 B.n224 VSUBS 0.011688f
C265 B.n225 VSUBS 0.011688f
C266 B.n226 VSUBS 0.011688f
C267 B.n227 VSUBS 0.011688f
C268 B.n228 VSUBS 0.011688f
C269 B.n229 VSUBS 0.011688f
C270 B.n230 VSUBS 0.011688f
C271 B.n231 VSUBS 0.011688f
C272 B.n232 VSUBS 0.011688f
C273 B.n233 VSUBS 0.011688f
C274 B.n234 VSUBS 0.011688f
C275 B.n235 VSUBS 0.011688f
C276 B.n236 VSUBS 0.011688f
C277 B.n237 VSUBS 0.011688f
C278 B.n238 VSUBS 0.011688f
C279 B.n239 VSUBS 0.011688f
C280 B.n240 VSUBS 0.011688f
C281 B.n241 VSUBS 0.011688f
C282 B.n242 VSUBS 0.011688f
C283 B.n243 VSUBS 0.011688f
C284 B.n244 VSUBS 0.011688f
C285 B.n245 VSUBS 0.011688f
C286 B.n246 VSUBS 0.011688f
C287 B.n247 VSUBS 0.011688f
C288 B.n248 VSUBS 0.011688f
C289 B.n249 VSUBS 0.011688f
C290 B.n250 VSUBS 0.011688f
C291 B.n251 VSUBS 0.011688f
C292 B.n252 VSUBS 0.011688f
C293 B.n253 VSUBS 0.011688f
C294 B.n254 VSUBS 0.011688f
C295 B.n255 VSUBS 0.011688f
C296 B.n256 VSUBS 0.011688f
C297 B.n257 VSUBS 0.011688f
C298 B.n258 VSUBS 0.011688f
C299 B.n259 VSUBS 0.011688f
C300 B.n260 VSUBS 0.011688f
C301 B.n261 VSUBS 0.011688f
C302 B.n262 VSUBS 0.011688f
C303 B.n263 VSUBS 0.011688f
C304 B.n264 VSUBS 0.011688f
C305 B.n265 VSUBS 0.011688f
C306 B.n266 VSUBS 0.011688f
C307 B.n267 VSUBS 0.011688f
C308 B.n268 VSUBS 0.011688f
C309 B.n269 VSUBS 0.011688f
C310 B.n270 VSUBS 0.011688f
C311 B.n271 VSUBS 0.027128f
C312 B.n272 VSUBS 0.028219f
C313 B.n273 VSUBS 0.028219f
C314 B.n274 VSUBS 0.011688f
C315 B.n275 VSUBS 0.011688f
C316 B.n276 VSUBS 0.011688f
C317 B.n277 VSUBS 0.011688f
C318 B.n278 VSUBS 0.011688f
C319 B.n279 VSUBS 0.011688f
C320 B.n280 VSUBS 0.011688f
C321 B.n281 VSUBS 0.011688f
C322 B.n282 VSUBS 0.011688f
C323 B.n283 VSUBS 0.011688f
C324 B.n284 VSUBS 0.011688f
C325 B.n285 VSUBS 0.011688f
C326 B.n286 VSUBS 0.011688f
C327 B.n287 VSUBS 0.011688f
C328 B.n288 VSUBS 0.008079f
C329 B.n289 VSUBS 0.02708f
C330 B.n290 VSUBS 0.009454f
C331 B.n291 VSUBS 0.011688f
C332 B.n292 VSUBS 0.011688f
C333 B.n293 VSUBS 0.011688f
C334 B.n294 VSUBS 0.011688f
C335 B.n295 VSUBS 0.011688f
C336 B.n296 VSUBS 0.011688f
C337 B.n297 VSUBS 0.011688f
C338 B.n298 VSUBS 0.011688f
C339 B.n299 VSUBS 0.011688f
C340 B.n300 VSUBS 0.011688f
C341 B.n301 VSUBS 0.011688f
C342 B.n302 VSUBS 0.009454f
C343 B.n303 VSUBS 0.02708f
C344 B.n304 VSUBS 0.008079f
C345 B.n305 VSUBS 0.011688f
C346 B.n306 VSUBS 0.011688f
C347 B.n307 VSUBS 0.011688f
C348 B.n308 VSUBS 0.011688f
C349 B.n309 VSUBS 0.011688f
C350 B.n310 VSUBS 0.011688f
C351 B.n311 VSUBS 0.011688f
C352 B.n312 VSUBS 0.011688f
C353 B.n313 VSUBS 0.011688f
C354 B.n314 VSUBS 0.011688f
C355 B.n315 VSUBS 0.011688f
C356 B.n316 VSUBS 0.011688f
C357 B.n317 VSUBS 0.011688f
C358 B.n318 VSUBS 0.011688f
C359 B.n319 VSUBS 0.028219f
C360 B.n320 VSUBS 0.026863f
C361 B.n321 VSUBS 0.028484f
C362 B.n322 VSUBS 0.011688f
C363 B.n323 VSUBS 0.011688f
C364 B.n324 VSUBS 0.011688f
C365 B.n325 VSUBS 0.011688f
C366 B.n326 VSUBS 0.011688f
C367 B.n327 VSUBS 0.011688f
C368 B.n328 VSUBS 0.011688f
C369 B.n329 VSUBS 0.011688f
C370 B.n330 VSUBS 0.011688f
C371 B.n331 VSUBS 0.011688f
C372 B.n332 VSUBS 0.011688f
C373 B.n333 VSUBS 0.011688f
C374 B.n334 VSUBS 0.011688f
C375 B.n335 VSUBS 0.011688f
C376 B.n336 VSUBS 0.011688f
C377 B.n337 VSUBS 0.011688f
C378 B.n338 VSUBS 0.011688f
C379 B.n339 VSUBS 0.011688f
C380 B.n340 VSUBS 0.011688f
C381 B.n341 VSUBS 0.011688f
C382 B.n342 VSUBS 0.011688f
C383 B.n343 VSUBS 0.011688f
C384 B.n344 VSUBS 0.011688f
C385 B.n345 VSUBS 0.011688f
C386 B.n346 VSUBS 0.011688f
C387 B.n347 VSUBS 0.011688f
C388 B.n348 VSUBS 0.011688f
C389 B.n349 VSUBS 0.011688f
C390 B.n350 VSUBS 0.011688f
C391 B.n351 VSUBS 0.011688f
C392 B.n352 VSUBS 0.011688f
C393 B.n353 VSUBS 0.011688f
C394 B.n354 VSUBS 0.011688f
C395 B.n355 VSUBS 0.011688f
C396 B.n356 VSUBS 0.011688f
C397 B.n357 VSUBS 0.011688f
C398 B.n358 VSUBS 0.011688f
C399 B.n359 VSUBS 0.011688f
C400 B.n360 VSUBS 0.011688f
C401 B.n361 VSUBS 0.011688f
C402 B.n362 VSUBS 0.011688f
C403 B.n363 VSUBS 0.011688f
C404 B.n364 VSUBS 0.011688f
C405 B.n365 VSUBS 0.011688f
C406 B.n366 VSUBS 0.011688f
C407 B.n367 VSUBS 0.011688f
C408 B.n368 VSUBS 0.011688f
C409 B.n369 VSUBS 0.011688f
C410 B.n370 VSUBS 0.011688f
C411 B.n371 VSUBS 0.011688f
C412 B.n372 VSUBS 0.011688f
C413 B.n373 VSUBS 0.011688f
C414 B.n374 VSUBS 0.011688f
C415 B.n375 VSUBS 0.011688f
C416 B.n376 VSUBS 0.011688f
C417 B.n377 VSUBS 0.011688f
C418 B.n378 VSUBS 0.011688f
C419 B.n379 VSUBS 0.011688f
C420 B.n380 VSUBS 0.011688f
C421 B.n381 VSUBS 0.011688f
C422 B.n382 VSUBS 0.011688f
C423 B.n383 VSUBS 0.011688f
C424 B.n384 VSUBS 0.011688f
C425 B.n385 VSUBS 0.011688f
C426 B.n386 VSUBS 0.011688f
C427 B.n387 VSUBS 0.011688f
C428 B.n388 VSUBS 0.011688f
C429 B.n389 VSUBS 0.011688f
C430 B.n390 VSUBS 0.011688f
C431 B.n391 VSUBS 0.011688f
C432 B.n392 VSUBS 0.011688f
C433 B.n393 VSUBS 0.011688f
C434 B.n394 VSUBS 0.011688f
C435 B.n395 VSUBS 0.011688f
C436 B.n396 VSUBS 0.011688f
C437 B.n397 VSUBS 0.011688f
C438 B.n398 VSUBS 0.011688f
C439 B.n399 VSUBS 0.011688f
C440 B.n400 VSUBS 0.011688f
C441 B.n401 VSUBS 0.011688f
C442 B.n402 VSUBS 0.011688f
C443 B.n403 VSUBS 0.011688f
C444 B.n404 VSUBS 0.011688f
C445 B.n405 VSUBS 0.011688f
C446 B.n406 VSUBS 0.011688f
C447 B.n407 VSUBS 0.011688f
C448 B.n408 VSUBS 0.011688f
C449 B.n409 VSUBS 0.011688f
C450 B.n410 VSUBS 0.011688f
C451 B.n411 VSUBS 0.011688f
C452 B.n412 VSUBS 0.011688f
C453 B.n413 VSUBS 0.011688f
C454 B.n414 VSUBS 0.011688f
C455 B.n415 VSUBS 0.011688f
C456 B.n416 VSUBS 0.011688f
C457 B.n417 VSUBS 0.011688f
C458 B.n418 VSUBS 0.011688f
C459 B.n419 VSUBS 0.011688f
C460 B.n420 VSUBS 0.011688f
C461 B.n421 VSUBS 0.011688f
C462 B.n422 VSUBS 0.011688f
C463 B.n423 VSUBS 0.011688f
C464 B.n424 VSUBS 0.011688f
C465 B.n425 VSUBS 0.011688f
C466 B.n426 VSUBS 0.011688f
C467 B.n427 VSUBS 0.011688f
C468 B.n428 VSUBS 0.011688f
C469 B.n429 VSUBS 0.011688f
C470 B.n430 VSUBS 0.011688f
C471 B.n431 VSUBS 0.011688f
C472 B.n432 VSUBS 0.011688f
C473 B.n433 VSUBS 0.011688f
C474 B.n434 VSUBS 0.011688f
C475 B.n435 VSUBS 0.011688f
C476 B.n436 VSUBS 0.011688f
C477 B.n437 VSUBS 0.011688f
C478 B.n438 VSUBS 0.011688f
C479 B.n439 VSUBS 0.011688f
C480 B.n440 VSUBS 0.011688f
C481 B.n441 VSUBS 0.011688f
C482 B.n442 VSUBS 0.011688f
C483 B.n443 VSUBS 0.011688f
C484 B.n444 VSUBS 0.011688f
C485 B.n445 VSUBS 0.011688f
C486 B.n446 VSUBS 0.011688f
C487 B.n447 VSUBS 0.011688f
C488 B.n448 VSUBS 0.011688f
C489 B.n449 VSUBS 0.011688f
C490 B.n450 VSUBS 0.011688f
C491 B.n451 VSUBS 0.011688f
C492 B.n452 VSUBS 0.011688f
C493 B.n453 VSUBS 0.011688f
C494 B.n454 VSUBS 0.011688f
C495 B.n455 VSUBS 0.011688f
C496 B.n456 VSUBS 0.011688f
C497 B.n457 VSUBS 0.011688f
C498 B.n458 VSUBS 0.011688f
C499 B.n459 VSUBS 0.011688f
C500 B.n460 VSUBS 0.011688f
C501 B.n461 VSUBS 0.011688f
C502 B.n462 VSUBS 0.011688f
C503 B.n463 VSUBS 0.011688f
C504 B.n464 VSUBS 0.011688f
C505 B.n465 VSUBS 0.011688f
C506 B.n466 VSUBS 0.011688f
C507 B.n467 VSUBS 0.011688f
C508 B.n468 VSUBS 0.011688f
C509 B.n469 VSUBS 0.011688f
C510 B.n470 VSUBS 0.011688f
C511 B.n471 VSUBS 0.011688f
C512 B.n472 VSUBS 0.011688f
C513 B.n473 VSUBS 0.011688f
C514 B.n474 VSUBS 0.011688f
C515 B.n475 VSUBS 0.011688f
C516 B.n476 VSUBS 0.011688f
C517 B.n477 VSUBS 0.011688f
C518 B.n478 VSUBS 0.011688f
C519 B.n479 VSUBS 0.011688f
C520 B.n480 VSUBS 0.011688f
C521 B.n481 VSUBS 0.011688f
C522 B.n482 VSUBS 0.011688f
C523 B.n483 VSUBS 0.011688f
C524 B.n484 VSUBS 0.011688f
C525 B.n485 VSUBS 0.011688f
C526 B.n486 VSUBS 0.011688f
C527 B.n487 VSUBS 0.011688f
C528 B.n488 VSUBS 0.011688f
C529 B.n489 VSUBS 0.011688f
C530 B.n490 VSUBS 0.011688f
C531 B.n491 VSUBS 0.011688f
C532 B.n492 VSUBS 0.011688f
C533 B.n493 VSUBS 0.011688f
C534 B.n494 VSUBS 0.011688f
C535 B.n495 VSUBS 0.011688f
C536 B.n496 VSUBS 0.011688f
C537 B.n497 VSUBS 0.011688f
C538 B.n498 VSUBS 0.011688f
C539 B.n499 VSUBS 0.011688f
C540 B.n500 VSUBS 0.011688f
C541 B.n501 VSUBS 0.011688f
C542 B.n502 VSUBS 0.011688f
C543 B.n503 VSUBS 0.011688f
C544 B.n504 VSUBS 0.011688f
C545 B.n505 VSUBS 0.011688f
C546 B.n506 VSUBS 0.011688f
C547 B.n507 VSUBS 0.011688f
C548 B.n508 VSUBS 0.011688f
C549 B.n509 VSUBS 0.011688f
C550 B.n510 VSUBS 0.011688f
C551 B.n511 VSUBS 0.011688f
C552 B.n512 VSUBS 0.011688f
C553 B.n513 VSUBS 0.011688f
C554 B.n514 VSUBS 0.011688f
C555 B.n515 VSUBS 0.011688f
C556 B.n516 VSUBS 0.011688f
C557 B.n517 VSUBS 0.011688f
C558 B.n518 VSUBS 0.011688f
C559 B.n519 VSUBS 0.011688f
C560 B.n520 VSUBS 0.027128f
C561 B.n521 VSUBS 0.027128f
C562 B.n522 VSUBS 0.028219f
C563 B.n523 VSUBS 0.011688f
C564 B.n524 VSUBS 0.011688f
C565 B.n525 VSUBS 0.011688f
C566 B.n526 VSUBS 0.011688f
C567 B.n527 VSUBS 0.011688f
C568 B.n528 VSUBS 0.011688f
C569 B.n529 VSUBS 0.011688f
C570 B.n530 VSUBS 0.011688f
C571 B.n531 VSUBS 0.011688f
C572 B.n532 VSUBS 0.011688f
C573 B.n533 VSUBS 0.011688f
C574 B.n534 VSUBS 0.011688f
C575 B.n535 VSUBS 0.011688f
C576 B.n536 VSUBS 0.011688f
C577 B.n537 VSUBS 0.008079f
C578 B.n538 VSUBS 0.02708f
C579 B.n539 VSUBS 0.009454f
C580 B.n540 VSUBS 0.011688f
C581 B.n541 VSUBS 0.011688f
C582 B.n542 VSUBS 0.011688f
C583 B.n543 VSUBS 0.011688f
C584 B.n544 VSUBS 0.011688f
C585 B.n545 VSUBS 0.011688f
C586 B.n546 VSUBS 0.011688f
C587 B.n547 VSUBS 0.011688f
C588 B.n548 VSUBS 0.011688f
C589 B.n549 VSUBS 0.011688f
C590 B.n550 VSUBS 0.011688f
C591 B.n551 VSUBS 0.009454f
C592 B.n552 VSUBS 0.011688f
C593 B.n553 VSUBS 0.011688f
C594 B.n554 VSUBS 0.011688f
C595 B.n555 VSUBS 0.011688f
C596 B.n556 VSUBS 0.011688f
C597 B.n557 VSUBS 0.011688f
C598 B.n558 VSUBS 0.011688f
C599 B.n559 VSUBS 0.011688f
C600 B.n560 VSUBS 0.011688f
C601 B.n561 VSUBS 0.011688f
C602 B.n562 VSUBS 0.011688f
C603 B.n563 VSUBS 0.011688f
C604 B.n564 VSUBS 0.011688f
C605 B.n565 VSUBS 0.011688f
C606 B.n566 VSUBS 0.011688f
C607 B.n567 VSUBS 0.011688f
C608 B.n568 VSUBS 0.028219f
C609 B.n569 VSUBS 0.027128f
C610 B.n570 VSUBS 0.027128f
C611 B.n571 VSUBS 0.011688f
C612 B.n572 VSUBS 0.011688f
C613 B.n573 VSUBS 0.011688f
C614 B.n574 VSUBS 0.011688f
C615 B.n575 VSUBS 0.011688f
C616 B.n576 VSUBS 0.011688f
C617 B.n577 VSUBS 0.011688f
C618 B.n578 VSUBS 0.011688f
C619 B.n579 VSUBS 0.011688f
C620 B.n580 VSUBS 0.011688f
C621 B.n581 VSUBS 0.011688f
C622 B.n582 VSUBS 0.011688f
C623 B.n583 VSUBS 0.011688f
C624 B.n584 VSUBS 0.011688f
C625 B.n585 VSUBS 0.011688f
C626 B.n586 VSUBS 0.011688f
C627 B.n587 VSUBS 0.011688f
C628 B.n588 VSUBS 0.011688f
C629 B.n589 VSUBS 0.011688f
C630 B.n590 VSUBS 0.011688f
C631 B.n591 VSUBS 0.011688f
C632 B.n592 VSUBS 0.011688f
C633 B.n593 VSUBS 0.011688f
C634 B.n594 VSUBS 0.011688f
C635 B.n595 VSUBS 0.011688f
C636 B.n596 VSUBS 0.011688f
C637 B.n597 VSUBS 0.011688f
C638 B.n598 VSUBS 0.011688f
C639 B.n599 VSUBS 0.011688f
C640 B.n600 VSUBS 0.011688f
C641 B.n601 VSUBS 0.011688f
C642 B.n602 VSUBS 0.011688f
C643 B.n603 VSUBS 0.011688f
C644 B.n604 VSUBS 0.011688f
C645 B.n605 VSUBS 0.011688f
C646 B.n606 VSUBS 0.011688f
C647 B.n607 VSUBS 0.011688f
C648 B.n608 VSUBS 0.011688f
C649 B.n609 VSUBS 0.011688f
C650 B.n610 VSUBS 0.011688f
C651 B.n611 VSUBS 0.011688f
C652 B.n612 VSUBS 0.011688f
C653 B.n613 VSUBS 0.011688f
C654 B.n614 VSUBS 0.011688f
C655 B.n615 VSUBS 0.011688f
C656 B.n616 VSUBS 0.011688f
C657 B.n617 VSUBS 0.011688f
C658 B.n618 VSUBS 0.011688f
C659 B.n619 VSUBS 0.011688f
C660 B.n620 VSUBS 0.011688f
C661 B.n621 VSUBS 0.011688f
C662 B.n622 VSUBS 0.011688f
C663 B.n623 VSUBS 0.011688f
C664 B.n624 VSUBS 0.011688f
C665 B.n625 VSUBS 0.011688f
C666 B.n626 VSUBS 0.011688f
C667 B.n627 VSUBS 0.011688f
C668 B.n628 VSUBS 0.011688f
C669 B.n629 VSUBS 0.011688f
C670 B.n630 VSUBS 0.011688f
C671 B.n631 VSUBS 0.011688f
C672 B.n632 VSUBS 0.011688f
C673 B.n633 VSUBS 0.011688f
C674 B.n634 VSUBS 0.011688f
C675 B.n635 VSUBS 0.011688f
C676 B.n636 VSUBS 0.011688f
C677 B.n637 VSUBS 0.011688f
C678 B.n638 VSUBS 0.011688f
C679 B.n639 VSUBS 0.011688f
C680 B.n640 VSUBS 0.011688f
C681 B.n641 VSUBS 0.011688f
C682 B.n642 VSUBS 0.011688f
C683 B.n643 VSUBS 0.011688f
C684 B.n644 VSUBS 0.011688f
C685 B.n645 VSUBS 0.011688f
C686 B.n646 VSUBS 0.011688f
C687 B.n647 VSUBS 0.011688f
C688 B.n648 VSUBS 0.011688f
C689 B.n649 VSUBS 0.011688f
C690 B.n650 VSUBS 0.011688f
C691 B.n651 VSUBS 0.011688f
C692 B.n652 VSUBS 0.011688f
C693 B.n653 VSUBS 0.011688f
C694 B.n654 VSUBS 0.011688f
C695 B.n655 VSUBS 0.011688f
C696 B.n656 VSUBS 0.011688f
C697 B.n657 VSUBS 0.011688f
C698 B.n658 VSUBS 0.011688f
C699 B.n659 VSUBS 0.011688f
C700 B.n660 VSUBS 0.011688f
C701 B.n661 VSUBS 0.011688f
C702 B.n662 VSUBS 0.011688f
C703 B.n663 VSUBS 0.011688f
C704 B.n664 VSUBS 0.011688f
C705 B.n665 VSUBS 0.011688f
C706 B.n666 VSUBS 0.011688f
C707 B.n667 VSUBS 0.015252f
C708 B.n668 VSUBS 0.016248f
C709 B.n669 VSUBS 0.03231f
C710 VDD1.t6 VSUBS 0.047179f
C711 VDD1.t2 VSUBS 0.047179f
C712 VDD1.n0 VSUBS 0.187842f
C713 VDD1.t7 VSUBS 0.047179f
C714 VDD1.t4 VSUBS 0.047179f
C715 VDD1.n1 VSUBS 0.187287f
C716 VDD1.t1 VSUBS 0.047179f
C717 VDD1.t3 VSUBS 0.047179f
C718 VDD1.n2 VSUBS 0.187287f
C719 VDD1.n3 VSUBS 5.28773f
C720 VDD1.t0 VSUBS 0.047179f
C721 VDD1.t5 VSUBS 0.047179f
C722 VDD1.n4 VSUBS 0.180563f
C723 VDD1.n5 VSUBS 4.02477f
C724 VP.t4 VSUBS 0.756196f
C725 VP.n0 VSUBS 0.632409f
C726 VP.n1 VSUBS 0.062469f
C727 VP.n2 VSUBS 0.096849f
C728 VP.n3 VSUBS 0.062469f
C729 VP.n4 VSUBS 0.089857f
C730 VP.n5 VSUBS 0.062469f
C731 VP.n6 VSUBS 0.09159f
C732 VP.n7 VSUBS 0.062469f
C733 VP.n8 VSUBS 0.086391f
C734 VP.n9 VSUBS 0.062469f
C735 VP.n10 VSUBS 0.086331f
C736 VP.n11 VSUBS 0.062469f
C737 VP.n12 VSUBS 0.082924f
C738 VP.t2 VSUBS 0.756196f
C739 VP.n13 VSUBS 0.632409f
C740 VP.n14 VSUBS 0.062469f
C741 VP.n15 VSUBS 0.096849f
C742 VP.n16 VSUBS 0.062469f
C743 VP.n17 VSUBS 0.089857f
C744 VP.n18 VSUBS 0.062469f
C745 VP.n19 VSUBS 0.09159f
C746 VP.n20 VSUBS 0.062469f
C747 VP.n21 VSUBS 0.086391f
C748 VP.t1 VSUBS 1.41912f
C749 VP.t5 VSUBS 0.756196f
C750 VP.n22 VSUBS 0.598432f
C751 VP.n23 VSUBS 0.702731f
C752 VP.n24 VSUBS 0.782898f
C753 VP.n25 VSUBS 0.062469f
C754 VP.n26 VSUBS 0.11701f
C755 VP.n27 VSUBS 0.11701f
C756 VP.n28 VSUBS 0.09159f
C757 VP.n29 VSUBS 0.062469f
C758 VP.n30 VSUBS 0.062469f
C759 VP.n31 VSUBS 0.062469f
C760 VP.n32 VSUBS 0.11701f
C761 VP.n33 VSUBS 0.11701f
C762 VP.t7 VSUBS 0.756196f
C763 VP.n34 VSUBS 0.380642f
C764 VP.n35 VSUBS 0.086391f
C765 VP.n36 VSUBS 0.062469f
C766 VP.n37 VSUBS 0.062469f
C767 VP.n38 VSUBS 0.062469f
C768 VP.n39 VSUBS 0.11701f
C769 VP.n40 VSUBS 0.11701f
C770 VP.n41 VSUBS 0.086331f
C771 VP.n42 VSUBS 0.062469f
C772 VP.n43 VSUBS 0.062469f
C773 VP.n44 VSUBS 0.062469f
C774 VP.n45 VSUBS 0.11701f
C775 VP.n46 VSUBS 0.11701f
C776 VP.n47 VSUBS 0.082924f
C777 VP.n48 VSUBS 0.100839f
C778 VP.n49 VSUBS 3.36842f
C779 VP.t0 VSUBS 0.756196f
C780 VP.n50 VSUBS 0.632409f
C781 VP.n51 VSUBS 3.41512f
C782 VP.n52 VSUBS 0.100839f
C783 VP.n53 VSUBS 0.062469f
C784 VP.n54 VSUBS 0.11701f
C785 VP.n55 VSUBS 0.11701f
C786 VP.n56 VSUBS 0.096849f
C787 VP.n57 VSUBS 0.062469f
C788 VP.n58 VSUBS 0.062469f
C789 VP.n59 VSUBS 0.062469f
C790 VP.n60 VSUBS 0.11701f
C791 VP.n61 VSUBS 0.11701f
C792 VP.t3 VSUBS 0.756196f
C793 VP.n62 VSUBS 0.380642f
C794 VP.n63 VSUBS 0.089857f
C795 VP.n64 VSUBS 0.062469f
C796 VP.n65 VSUBS 0.062469f
C797 VP.n66 VSUBS 0.062469f
C798 VP.n67 VSUBS 0.11701f
C799 VP.n68 VSUBS 0.11701f
C800 VP.n69 VSUBS 0.09159f
C801 VP.n70 VSUBS 0.062469f
C802 VP.n71 VSUBS 0.062469f
C803 VP.n72 VSUBS 0.062469f
C804 VP.n73 VSUBS 0.11701f
C805 VP.n74 VSUBS 0.11701f
C806 VP.t6 VSUBS 0.756196f
C807 VP.n75 VSUBS 0.380642f
C808 VP.n76 VSUBS 0.086391f
C809 VP.n77 VSUBS 0.062469f
C810 VP.n78 VSUBS 0.062469f
C811 VP.n79 VSUBS 0.062469f
C812 VP.n80 VSUBS 0.11701f
C813 VP.n81 VSUBS 0.11701f
C814 VP.n82 VSUBS 0.086331f
C815 VP.n83 VSUBS 0.062469f
C816 VP.n84 VSUBS 0.062469f
C817 VP.n85 VSUBS 0.062469f
C818 VP.n86 VSUBS 0.11701f
C819 VP.n87 VSUBS 0.11701f
C820 VP.n88 VSUBS 0.082924f
C821 VP.n89 VSUBS 0.100839f
C822 VP.n90 VSUBS 0.172054f
C823 VTAIL.t9 VSUBS 0.043833f
C824 VTAIL.t11 VSUBS 0.043833f
C825 VTAIL.n0 VSUBS 0.143931f
C826 VTAIL.n1 VSUBS 0.725687f
C827 VTAIL.t14 VSUBS 0.245133f
C828 VTAIL.n2 VSUBS 0.792435f
C829 VTAIL.t6 VSUBS 0.245133f
C830 VTAIL.n3 VSUBS 0.792435f
C831 VTAIL.t4 VSUBS 0.043833f
C832 VTAIL.t0 VSUBS 0.043833f
C833 VTAIL.n4 VSUBS 0.143931f
C834 VTAIL.n5 VSUBS 1.12128f
C835 VTAIL.t5 VSUBS 0.245133f
C836 VTAIL.n6 VSUBS 1.78942f
C837 VTAIL.t8 VSUBS 0.245133f
C838 VTAIL.n7 VSUBS 1.78942f
C839 VTAIL.t10 VSUBS 0.043833f
C840 VTAIL.t15 VSUBS 0.043833f
C841 VTAIL.n8 VSUBS 0.143932f
C842 VTAIL.n9 VSUBS 1.12128f
C843 VTAIL.t13 VSUBS 0.245133f
C844 VTAIL.n10 VSUBS 0.792435f
C845 VTAIL.t1 VSUBS 0.245133f
C846 VTAIL.n11 VSUBS 0.792435f
C847 VTAIL.t7 VSUBS 0.043833f
C848 VTAIL.t3 VSUBS 0.043833f
C849 VTAIL.n12 VSUBS 0.143932f
C850 VTAIL.n13 VSUBS 1.12128f
C851 VTAIL.t2 VSUBS 0.245133f
C852 VTAIL.n14 VSUBS 1.78942f
C853 VTAIL.t12 VSUBS 0.245133f
C854 VTAIL.n15 VSUBS 1.78258f
C855 VDD2.t2 VSUBS 0.040537f
C856 VDD2.t6 VSUBS 0.040537f
C857 VDD2.n0 VSUBS 0.16092f
C858 VDD2.t4 VSUBS 0.040537f
C859 VDD2.t5 VSUBS 0.040537f
C860 VDD2.n1 VSUBS 0.16092f
C861 VDD2.n2 VSUBS 4.47346f
C862 VDD2.t1 VSUBS 0.040537f
C863 VDD2.t0 VSUBS 0.040537f
C864 VDD2.n3 VSUBS 0.155143f
C865 VDD2.n4 VSUBS 3.41597f
C866 VDD2.t7 VSUBS 0.040537f
C867 VDD2.t3 VSUBS 0.040537f
C868 VDD2.n5 VSUBS 0.160905f
C869 VN.t3 VSUBS 0.603478f
C870 VN.n0 VSUBS 0.50469f
C871 VN.n1 VSUBS 0.049853f
C872 VN.n2 VSUBS 0.07729f
C873 VN.n3 VSUBS 0.049853f
C874 VN.n4 VSUBS 0.07171f
C875 VN.n5 VSUBS 0.049853f
C876 VN.n6 VSUBS 0.073093f
C877 VN.n7 VSUBS 0.049853f
C878 VN.n8 VSUBS 0.068944f
C879 VN.t6 VSUBS 0.603478f
C880 VN.n9 VSUBS 0.477575f
C881 VN.t1 VSUBS 1.13252f
C882 VN.n10 VSUBS 0.560809f
C883 VN.n11 VSUBS 0.624786f
C884 VN.n12 VSUBS 0.049853f
C885 VN.n13 VSUBS 0.093379f
C886 VN.n14 VSUBS 0.093379f
C887 VN.n15 VSUBS 0.073093f
C888 VN.n16 VSUBS 0.049853f
C889 VN.n17 VSUBS 0.049853f
C890 VN.n18 VSUBS 0.049853f
C891 VN.n19 VSUBS 0.093379f
C892 VN.n20 VSUBS 0.093379f
C893 VN.t4 VSUBS 0.603478f
C894 VN.n21 VSUBS 0.303769f
C895 VN.n22 VSUBS 0.068944f
C896 VN.n23 VSUBS 0.049853f
C897 VN.n24 VSUBS 0.049853f
C898 VN.n25 VSUBS 0.049853f
C899 VN.n26 VSUBS 0.093379f
C900 VN.n27 VSUBS 0.093379f
C901 VN.n28 VSUBS 0.068896f
C902 VN.n29 VSUBS 0.049853f
C903 VN.n30 VSUBS 0.049853f
C904 VN.n31 VSUBS 0.049853f
C905 VN.n32 VSUBS 0.093379f
C906 VN.n33 VSUBS 0.093379f
C907 VN.n34 VSUBS 0.066177f
C908 VN.n35 VSUBS 0.080474f
C909 VN.n36 VSUBS 0.137307f
C910 VN.t7 VSUBS 0.603478f
C911 VN.n37 VSUBS 0.50469f
C912 VN.n38 VSUBS 0.049853f
C913 VN.n39 VSUBS 0.07729f
C914 VN.n40 VSUBS 0.049853f
C915 VN.n41 VSUBS 0.07171f
C916 VN.n42 VSUBS 0.049853f
C917 VN.t5 VSUBS 0.603478f
C918 VN.n43 VSUBS 0.303769f
C919 VN.n44 VSUBS 0.073093f
C920 VN.n45 VSUBS 0.049853f
C921 VN.n46 VSUBS 0.068944f
C922 VN.t2 VSUBS 1.13252f
C923 VN.t0 VSUBS 0.603478f
C924 VN.n47 VSUBS 0.477575f
C925 VN.n48 VSUBS 0.560809f
C926 VN.n49 VSUBS 0.624786f
C927 VN.n50 VSUBS 0.049853f
C928 VN.n51 VSUBS 0.093379f
C929 VN.n52 VSUBS 0.093379f
C930 VN.n53 VSUBS 0.073093f
C931 VN.n54 VSUBS 0.049853f
C932 VN.n55 VSUBS 0.049853f
C933 VN.n56 VSUBS 0.049853f
C934 VN.n57 VSUBS 0.093379f
C935 VN.n58 VSUBS 0.093379f
C936 VN.n59 VSUBS 0.068944f
C937 VN.n60 VSUBS 0.049853f
C938 VN.n61 VSUBS 0.049853f
C939 VN.n62 VSUBS 0.049853f
C940 VN.n63 VSUBS 0.093379f
C941 VN.n64 VSUBS 0.093379f
C942 VN.n65 VSUBS 0.068896f
C943 VN.n66 VSUBS 0.049853f
C944 VN.n67 VSUBS 0.049853f
C945 VN.n68 VSUBS 0.049853f
C946 VN.n69 VSUBS 0.093379f
C947 VN.n70 VSUBS 0.093379f
C948 VN.n71 VSUBS 0.066177f
C949 VN.n72 VSUBS 0.080474f
C950 VN.n73 VSUBS 2.70883f
.ends

