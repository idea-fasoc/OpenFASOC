* NGSPICE file created from diff_pair_sample_0076.ext - technology: sky130A

.subckt diff_pair_sample_0076 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=0 ps=0 w=10.32 l=1.68
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=4.0248 ps=21.42 w=10.32 l=1.68
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=0 ps=0 w=10.32 l=1.68
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=0 ps=0 w=10.32 l=1.68
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=4.0248 ps=21.42 w=10.32 l=1.68
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=0 ps=0 w=10.32 l=1.68
X6 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=4.0248 ps=21.42 w=10.32 l=1.68
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0248 pd=21.42 as=4.0248 ps=21.42 w=10.32 l=1.68
R0 B.n588 B.n587 585
R1 B.n589 B.n588 585
R2 B.n249 B.n82 585
R3 B.n248 B.n247 585
R4 B.n246 B.n245 585
R5 B.n244 B.n243 585
R6 B.n242 B.n241 585
R7 B.n240 B.n239 585
R8 B.n238 B.n237 585
R9 B.n236 B.n235 585
R10 B.n234 B.n233 585
R11 B.n232 B.n231 585
R12 B.n230 B.n229 585
R13 B.n228 B.n227 585
R14 B.n226 B.n225 585
R15 B.n224 B.n223 585
R16 B.n222 B.n221 585
R17 B.n220 B.n219 585
R18 B.n218 B.n217 585
R19 B.n216 B.n215 585
R20 B.n214 B.n213 585
R21 B.n212 B.n211 585
R22 B.n210 B.n209 585
R23 B.n208 B.n207 585
R24 B.n206 B.n205 585
R25 B.n204 B.n203 585
R26 B.n202 B.n201 585
R27 B.n200 B.n199 585
R28 B.n198 B.n197 585
R29 B.n196 B.n195 585
R30 B.n194 B.n193 585
R31 B.n192 B.n191 585
R32 B.n190 B.n189 585
R33 B.n188 B.n187 585
R34 B.n186 B.n185 585
R35 B.n184 B.n183 585
R36 B.n182 B.n181 585
R37 B.n180 B.n179 585
R38 B.n178 B.n177 585
R39 B.n176 B.n175 585
R40 B.n174 B.n173 585
R41 B.n172 B.n171 585
R42 B.n170 B.n169 585
R43 B.n168 B.n167 585
R44 B.n166 B.n165 585
R45 B.n164 B.n163 585
R46 B.n162 B.n161 585
R47 B.n159 B.n158 585
R48 B.n157 B.n156 585
R49 B.n155 B.n154 585
R50 B.n153 B.n152 585
R51 B.n151 B.n150 585
R52 B.n149 B.n148 585
R53 B.n147 B.n146 585
R54 B.n145 B.n144 585
R55 B.n143 B.n142 585
R56 B.n141 B.n140 585
R57 B.n139 B.n138 585
R58 B.n137 B.n136 585
R59 B.n135 B.n134 585
R60 B.n133 B.n132 585
R61 B.n131 B.n130 585
R62 B.n129 B.n128 585
R63 B.n127 B.n126 585
R64 B.n125 B.n124 585
R65 B.n123 B.n122 585
R66 B.n121 B.n120 585
R67 B.n119 B.n118 585
R68 B.n117 B.n116 585
R69 B.n115 B.n114 585
R70 B.n113 B.n112 585
R71 B.n111 B.n110 585
R72 B.n109 B.n108 585
R73 B.n107 B.n106 585
R74 B.n105 B.n104 585
R75 B.n103 B.n102 585
R76 B.n101 B.n100 585
R77 B.n99 B.n98 585
R78 B.n97 B.n96 585
R79 B.n95 B.n94 585
R80 B.n93 B.n92 585
R81 B.n91 B.n90 585
R82 B.n89 B.n88 585
R83 B.n39 B.n38 585
R84 B.n586 B.n40 585
R85 B.n590 B.n40 585
R86 B.n585 B.n584 585
R87 B.n584 B.n36 585
R88 B.n583 B.n35 585
R89 B.n596 B.n35 585
R90 B.n582 B.n34 585
R91 B.n597 B.n34 585
R92 B.n581 B.n33 585
R93 B.n598 B.n33 585
R94 B.n580 B.n579 585
R95 B.n579 B.n29 585
R96 B.n578 B.n28 585
R97 B.n604 B.n28 585
R98 B.n577 B.n27 585
R99 B.n605 B.n27 585
R100 B.n576 B.n26 585
R101 B.n606 B.n26 585
R102 B.n575 B.n574 585
R103 B.n574 B.n22 585
R104 B.n573 B.n21 585
R105 B.n612 B.n21 585
R106 B.n572 B.n20 585
R107 B.n613 B.n20 585
R108 B.n571 B.n19 585
R109 B.n614 B.n19 585
R110 B.n570 B.n569 585
R111 B.n569 B.n15 585
R112 B.n568 B.n14 585
R113 B.n620 B.n14 585
R114 B.n567 B.n13 585
R115 B.n621 B.n13 585
R116 B.n566 B.n12 585
R117 B.n622 B.n12 585
R118 B.n565 B.n564 585
R119 B.n564 B.n8 585
R120 B.n563 B.n7 585
R121 B.n628 B.n7 585
R122 B.n562 B.n6 585
R123 B.n629 B.n6 585
R124 B.n561 B.n5 585
R125 B.n630 B.n5 585
R126 B.n560 B.n559 585
R127 B.n559 B.n4 585
R128 B.n558 B.n250 585
R129 B.n558 B.n557 585
R130 B.n548 B.n251 585
R131 B.n252 B.n251 585
R132 B.n550 B.n549 585
R133 B.n551 B.n550 585
R134 B.n547 B.n256 585
R135 B.n260 B.n256 585
R136 B.n546 B.n545 585
R137 B.n545 B.n544 585
R138 B.n258 B.n257 585
R139 B.n259 B.n258 585
R140 B.n537 B.n536 585
R141 B.n538 B.n537 585
R142 B.n535 B.n265 585
R143 B.n265 B.n264 585
R144 B.n534 B.n533 585
R145 B.n533 B.n532 585
R146 B.n267 B.n266 585
R147 B.n268 B.n267 585
R148 B.n525 B.n524 585
R149 B.n526 B.n525 585
R150 B.n523 B.n273 585
R151 B.n273 B.n272 585
R152 B.n522 B.n521 585
R153 B.n521 B.n520 585
R154 B.n275 B.n274 585
R155 B.n276 B.n275 585
R156 B.n513 B.n512 585
R157 B.n514 B.n513 585
R158 B.n511 B.n281 585
R159 B.n281 B.n280 585
R160 B.n510 B.n509 585
R161 B.n509 B.n508 585
R162 B.n283 B.n282 585
R163 B.n284 B.n283 585
R164 B.n501 B.n500 585
R165 B.n502 B.n501 585
R166 B.n287 B.n286 585
R167 B.n337 B.n336 585
R168 B.n338 B.n334 585
R169 B.n334 B.n288 585
R170 B.n340 B.n339 585
R171 B.n342 B.n333 585
R172 B.n345 B.n344 585
R173 B.n346 B.n332 585
R174 B.n348 B.n347 585
R175 B.n350 B.n331 585
R176 B.n353 B.n352 585
R177 B.n354 B.n330 585
R178 B.n356 B.n355 585
R179 B.n358 B.n329 585
R180 B.n361 B.n360 585
R181 B.n362 B.n328 585
R182 B.n364 B.n363 585
R183 B.n366 B.n327 585
R184 B.n369 B.n368 585
R185 B.n370 B.n326 585
R186 B.n372 B.n371 585
R187 B.n374 B.n325 585
R188 B.n377 B.n376 585
R189 B.n378 B.n324 585
R190 B.n380 B.n379 585
R191 B.n382 B.n323 585
R192 B.n385 B.n384 585
R193 B.n386 B.n322 585
R194 B.n388 B.n387 585
R195 B.n390 B.n321 585
R196 B.n393 B.n392 585
R197 B.n394 B.n320 585
R198 B.n396 B.n395 585
R199 B.n398 B.n319 585
R200 B.n401 B.n400 585
R201 B.n402 B.n318 585
R202 B.n404 B.n403 585
R203 B.n406 B.n317 585
R204 B.n409 B.n408 585
R205 B.n410 B.n313 585
R206 B.n412 B.n411 585
R207 B.n414 B.n312 585
R208 B.n417 B.n416 585
R209 B.n418 B.n311 585
R210 B.n420 B.n419 585
R211 B.n422 B.n310 585
R212 B.n425 B.n424 585
R213 B.n427 B.n307 585
R214 B.n429 B.n428 585
R215 B.n431 B.n306 585
R216 B.n434 B.n433 585
R217 B.n435 B.n305 585
R218 B.n437 B.n436 585
R219 B.n439 B.n304 585
R220 B.n442 B.n441 585
R221 B.n443 B.n303 585
R222 B.n445 B.n444 585
R223 B.n447 B.n302 585
R224 B.n450 B.n449 585
R225 B.n451 B.n301 585
R226 B.n453 B.n452 585
R227 B.n455 B.n300 585
R228 B.n458 B.n457 585
R229 B.n459 B.n299 585
R230 B.n461 B.n460 585
R231 B.n463 B.n298 585
R232 B.n466 B.n465 585
R233 B.n467 B.n297 585
R234 B.n469 B.n468 585
R235 B.n471 B.n296 585
R236 B.n474 B.n473 585
R237 B.n475 B.n295 585
R238 B.n477 B.n476 585
R239 B.n479 B.n294 585
R240 B.n482 B.n481 585
R241 B.n483 B.n293 585
R242 B.n485 B.n484 585
R243 B.n487 B.n292 585
R244 B.n490 B.n489 585
R245 B.n491 B.n291 585
R246 B.n493 B.n492 585
R247 B.n495 B.n290 585
R248 B.n498 B.n497 585
R249 B.n499 B.n289 585
R250 B.n504 B.n503 585
R251 B.n503 B.n502 585
R252 B.n505 B.n285 585
R253 B.n285 B.n284 585
R254 B.n507 B.n506 585
R255 B.n508 B.n507 585
R256 B.n279 B.n278 585
R257 B.n280 B.n279 585
R258 B.n516 B.n515 585
R259 B.n515 B.n514 585
R260 B.n517 B.n277 585
R261 B.n277 B.n276 585
R262 B.n519 B.n518 585
R263 B.n520 B.n519 585
R264 B.n271 B.n270 585
R265 B.n272 B.n271 585
R266 B.n528 B.n527 585
R267 B.n527 B.n526 585
R268 B.n529 B.n269 585
R269 B.n269 B.n268 585
R270 B.n531 B.n530 585
R271 B.n532 B.n531 585
R272 B.n263 B.n262 585
R273 B.n264 B.n263 585
R274 B.n540 B.n539 585
R275 B.n539 B.n538 585
R276 B.n541 B.n261 585
R277 B.n261 B.n259 585
R278 B.n543 B.n542 585
R279 B.n544 B.n543 585
R280 B.n255 B.n254 585
R281 B.n260 B.n255 585
R282 B.n553 B.n552 585
R283 B.n552 B.n551 585
R284 B.n554 B.n253 585
R285 B.n253 B.n252 585
R286 B.n556 B.n555 585
R287 B.n557 B.n556 585
R288 B.n2 B.n0 585
R289 B.n4 B.n2 585
R290 B.n3 B.n1 585
R291 B.n629 B.n3 585
R292 B.n627 B.n626 585
R293 B.n628 B.n627 585
R294 B.n625 B.n9 585
R295 B.n9 B.n8 585
R296 B.n624 B.n623 585
R297 B.n623 B.n622 585
R298 B.n11 B.n10 585
R299 B.n621 B.n11 585
R300 B.n619 B.n618 585
R301 B.n620 B.n619 585
R302 B.n617 B.n16 585
R303 B.n16 B.n15 585
R304 B.n616 B.n615 585
R305 B.n615 B.n614 585
R306 B.n18 B.n17 585
R307 B.n613 B.n18 585
R308 B.n611 B.n610 585
R309 B.n612 B.n611 585
R310 B.n609 B.n23 585
R311 B.n23 B.n22 585
R312 B.n608 B.n607 585
R313 B.n607 B.n606 585
R314 B.n25 B.n24 585
R315 B.n605 B.n25 585
R316 B.n603 B.n602 585
R317 B.n604 B.n603 585
R318 B.n601 B.n30 585
R319 B.n30 B.n29 585
R320 B.n600 B.n599 585
R321 B.n599 B.n598 585
R322 B.n32 B.n31 585
R323 B.n597 B.n32 585
R324 B.n595 B.n594 585
R325 B.n596 B.n595 585
R326 B.n593 B.n37 585
R327 B.n37 B.n36 585
R328 B.n592 B.n591 585
R329 B.n591 B.n590 585
R330 B.n632 B.n631 585
R331 B.n631 B.n630 585
R332 B.n503 B.n287 482.89
R333 B.n591 B.n39 482.89
R334 B.n501 B.n289 482.89
R335 B.n588 B.n40 482.89
R336 B.n308 B.t2 354.096
R337 B.n314 B.t10 354.096
R338 B.n86 B.t6 354.096
R339 B.n83 B.t13 354.096
R340 B.n589 B.n81 256.663
R341 B.n589 B.n80 256.663
R342 B.n589 B.n79 256.663
R343 B.n589 B.n78 256.663
R344 B.n589 B.n77 256.663
R345 B.n589 B.n76 256.663
R346 B.n589 B.n75 256.663
R347 B.n589 B.n74 256.663
R348 B.n589 B.n73 256.663
R349 B.n589 B.n72 256.663
R350 B.n589 B.n71 256.663
R351 B.n589 B.n70 256.663
R352 B.n589 B.n69 256.663
R353 B.n589 B.n68 256.663
R354 B.n589 B.n67 256.663
R355 B.n589 B.n66 256.663
R356 B.n589 B.n65 256.663
R357 B.n589 B.n64 256.663
R358 B.n589 B.n63 256.663
R359 B.n589 B.n62 256.663
R360 B.n589 B.n61 256.663
R361 B.n589 B.n60 256.663
R362 B.n589 B.n59 256.663
R363 B.n589 B.n58 256.663
R364 B.n589 B.n57 256.663
R365 B.n589 B.n56 256.663
R366 B.n589 B.n55 256.663
R367 B.n589 B.n54 256.663
R368 B.n589 B.n53 256.663
R369 B.n589 B.n52 256.663
R370 B.n589 B.n51 256.663
R371 B.n589 B.n50 256.663
R372 B.n589 B.n49 256.663
R373 B.n589 B.n48 256.663
R374 B.n589 B.n47 256.663
R375 B.n589 B.n46 256.663
R376 B.n589 B.n45 256.663
R377 B.n589 B.n44 256.663
R378 B.n589 B.n43 256.663
R379 B.n589 B.n42 256.663
R380 B.n589 B.n41 256.663
R381 B.n335 B.n288 256.663
R382 B.n341 B.n288 256.663
R383 B.n343 B.n288 256.663
R384 B.n349 B.n288 256.663
R385 B.n351 B.n288 256.663
R386 B.n357 B.n288 256.663
R387 B.n359 B.n288 256.663
R388 B.n365 B.n288 256.663
R389 B.n367 B.n288 256.663
R390 B.n373 B.n288 256.663
R391 B.n375 B.n288 256.663
R392 B.n381 B.n288 256.663
R393 B.n383 B.n288 256.663
R394 B.n389 B.n288 256.663
R395 B.n391 B.n288 256.663
R396 B.n397 B.n288 256.663
R397 B.n399 B.n288 256.663
R398 B.n405 B.n288 256.663
R399 B.n407 B.n288 256.663
R400 B.n413 B.n288 256.663
R401 B.n415 B.n288 256.663
R402 B.n421 B.n288 256.663
R403 B.n423 B.n288 256.663
R404 B.n430 B.n288 256.663
R405 B.n432 B.n288 256.663
R406 B.n438 B.n288 256.663
R407 B.n440 B.n288 256.663
R408 B.n446 B.n288 256.663
R409 B.n448 B.n288 256.663
R410 B.n454 B.n288 256.663
R411 B.n456 B.n288 256.663
R412 B.n462 B.n288 256.663
R413 B.n464 B.n288 256.663
R414 B.n470 B.n288 256.663
R415 B.n472 B.n288 256.663
R416 B.n478 B.n288 256.663
R417 B.n480 B.n288 256.663
R418 B.n486 B.n288 256.663
R419 B.n488 B.n288 256.663
R420 B.n494 B.n288 256.663
R421 B.n496 B.n288 256.663
R422 B.n503 B.n285 163.367
R423 B.n507 B.n285 163.367
R424 B.n507 B.n279 163.367
R425 B.n515 B.n279 163.367
R426 B.n515 B.n277 163.367
R427 B.n519 B.n277 163.367
R428 B.n519 B.n271 163.367
R429 B.n527 B.n271 163.367
R430 B.n527 B.n269 163.367
R431 B.n531 B.n269 163.367
R432 B.n531 B.n263 163.367
R433 B.n539 B.n263 163.367
R434 B.n539 B.n261 163.367
R435 B.n543 B.n261 163.367
R436 B.n543 B.n255 163.367
R437 B.n552 B.n255 163.367
R438 B.n552 B.n253 163.367
R439 B.n556 B.n253 163.367
R440 B.n556 B.n2 163.367
R441 B.n631 B.n2 163.367
R442 B.n631 B.n3 163.367
R443 B.n627 B.n3 163.367
R444 B.n627 B.n9 163.367
R445 B.n623 B.n9 163.367
R446 B.n623 B.n11 163.367
R447 B.n619 B.n11 163.367
R448 B.n619 B.n16 163.367
R449 B.n615 B.n16 163.367
R450 B.n615 B.n18 163.367
R451 B.n611 B.n18 163.367
R452 B.n611 B.n23 163.367
R453 B.n607 B.n23 163.367
R454 B.n607 B.n25 163.367
R455 B.n603 B.n25 163.367
R456 B.n603 B.n30 163.367
R457 B.n599 B.n30 163.367
R458 B.n599 B.n32 163.367
R459 B.n595 B.n32 163.367
R460 B.n595 B.n37 163.367
R461 B.n591 B.n37 163.367
R462 B.n336 B.n334 163.367
R463 B.n340 B.n334 163.367
R464 B.n344 B.n342 163.367
R465 B.n348 B.n332 163.367
R466 B.n352 B.n350 163.367
R467 B.n356 B.n330 163.367
R468 B.n360 B.n358 163.367
R469 B.n364 B.n328 163.367
R470 B.n368 B.n366 163.367
R471 B.n372 B.n326 163.367
R472 B.n376 B.n374 163.367
R473 B.n380 B.n324 163.367
R474 B.n384 B.n382 163.367
R475 B.n388 B.n322 163.367
R476 B.n392 B.n390 163.367
R477 B.n396 B.n320 163.367
R478 B.n400 B.n398 163.367
R479 B.n404 B.n318 163.367
R480 B.n408 B.n406 163.367
R481 B.n412 B.n313 163.367
R482 B.n416 B.n414 163.367
R483 B.n420 B.n311 163.367
R484 B.n424 B.n422 163.367
R485 B.n429 B.n307 163.367
R486 B.n433 B.n431 163.367
R487 B.n437 B.n305 163.367
R488 B.n441 B.n439 163.367
R489 B.n445 B.n303 163.367
R490 B.n449 B.n447 163.367
R491 B.n453 B.n301 163.367
R492 B.n457 B.n455 163.367
R493 B.n461 B.n299 163.367
R494 B.n465 B.n463 163.367
R495 B.n469 B.n297 163.367
R496 B.n473 B.n471 163.367
R497 B.n477 B.n295 163.367
R498 B.n481 B.n479 163.367
R499 B.n485 B.n293 163.367
R500 B.n489 B.n487 163.367
R501 B.n493 B.n291 163.367
R502 B.n497 B.n495 163.367
R503 B.n501 B.n283 163.367
R504 B.n509 B.n283 163.367
R505 B.n509 B.n281 163.367
R506 B.n513 B.n281 163.367
R507 B.n513 B.n275 163.367
R508 B.n521 B.n275 163.367
R509 B.n521 B.n273 163.367
R510 B.n525 B.n273 163.367
R511 B.n525 B.n267 163.367
R512 B.n533 B.n267 163.367
R513 B.n533 B.n265 163.367
R514 B.n537 B.n265 163.367
R515 B.n537 B.n258 163.367
R516 B.n545 B.n258 163.367
R517 B.n545 B.n256 163.367
R518 B.n550 B.n256 163.367
R519 B.n550 B.n251 163.367
R520 B.n558 B.n251 163.367
R521 B.n559 B.n558 163.367
R522 B.n559 B.n5 163.367
R523 B.n6 B.n5 163.367
R524 B.n7 B.n6 163.367
R525 B.n564 B.n7 163.367
R526 B.n564 B.n12 163.367
R527 B.n13 B.n12 163.367
R528 B.n14 B.n13 163.367
R529 B.n569 B.n14 163.367
R530 B.n569 B.n19 163.367
R531 B.n20 B.n19 163.367
R532 B.n21 B.n20 163.367
R533 B.n574 B.n21 163.367
R534 B.n574 B.n26 163.367
R535 B.n27 B.n26 163.367
R536 B.n28 B.n27 163.367
R537 B.n579 B.n28 163.367
R538 B.n579 B.n33 163.367
R539 B.n34 B.n33 163.367
R540 B.n35 B.n34 163.367
R541 B.n584 B.n35 163.367
R542 B.n584 B.n40 163.367
R543 B.n90 B.n89 163.367
R544 B.n94 B.n93 163.367
R545 B.n98 B.n97 163.367
R546 B.n102 B.n101 163.367
R547 B.n106 B.n105 163.367
R548 B.n110 B.n109 163.367
R549 B.n114 B.n113 163.367
R550 B.n118 B.n117 163.367
R551 B.n122 B.n121 163.367
R552 B.n126 B.n125 163.367
R553 B.n130 B.n129 163.367
R554 B.n134 B.n133 163.367
R555 B.n138 B.n137 163.367
R556 B.n142 B.n141 163.367
R557 B.n146 B.n145 163.367
R558 B.n150 B.n149 163.367
R559 B.n154 B.n153 163.367
R560 B.n158 B.n157 163.367
R561 B.n163 B.n162 163.367
R562 B.n167 B.n166 163.367
R563 B.n171 B.n170 163.367
R564 B.n175 B.n174 163.367
R565 B.n179 B.n178 163.367
R566 B.n183 B.n182 163.367
R567 B.n187 B.n186 163.367
R568 B.n191 B.n190 163.367
R569 B.n195 B.n194 163.367
R570 B.n199 B.n198 163.367
R571 B.n203 B.n202 163.367
R572 B.n207 B.n206 163.367
R573 B.n211 B.n210 163.367
R574 B.n215 B.n214 163.367
R575 B.n219 B.n218 163.367
R576 B.n223 B.n222 163.367
R577 B.n227 B.n226 163.367
R578 B.n231 B.n230 163.367
R579 B.n235 B.n234 163.367
R580 B.n239 B.n238 163.367
R581 B.n243 B.n242 163.367
R582 B.n247 B.n246 163.367
R583 B.n588 B.n82 163.367
R584 B.n308 B.t5 109.365
R585 B.n83 B.t14 109.365
R586 B.n314 B.t12 109.353
R587 B.n86 B.t8 109.353
R588 B.n502 B.n288 83.9377
R589 B.n590 B.n589 83.9377
R590 B.n335 B.n287 71.676
R591 B.n341 B.n340 71.676
R592 B.n344 B.n343 71.676
R593 B.n349 B.n348 71.676
R594 B.n352 B.n351 71.676
R595 B.n357 B.n356 71.676
R596 B.n360 B.n359 71.676
R597 B.n365 B.n364 71.676
R598 B.n368 B.n367 71.676
R599 B.n373 B.n372 71.676
R600 B.n376 B.n375 71.676
R601 B.n381 B.n380 71.676
R602 B.n384 B.n383 71.676
R603 B.n389 B.n388 71.676
R604 B.n392 B.n391 71.676
R605 B.n397 B.n396 71.676
R606 B.n400 B.n399 71.676
R607 B.n405 B.n404 71.676
R608 B.n408 B.n407 71.676
R609 B.n413 B.n412 71.676
R610 B.n416 B.n415 71.676
R611 B.n421 B.n420 71.676
R612 B.n424 B.n423 71.676
R613 B.n430 B.n429 71.676
R614 B.n433 B.n432 71.676
R615 B.n438 B.n437 71.676
R616 B.n441 B.n440 71.676
R617 B.n446 B.n445 71.676
R618 B.n449 B.n448 71.676
R619 B.n454 B.n453 71.676
R620 B.n457 B.n456 71.676
R621 B.n462 B.n461 71.676
R622 B.n465 B.n464 71.676
R623 B.n470 B.n469 71.676
R624 B.n473 B.n472 71.676
R625 B.n478 B.n477 71.676
R626 B.n481 B.n480 71.676
R627 B.n486 B.n485 71.676
R628 B.n489 B.n488 71.676
R629 B.n494 B.n493 71.676
R630 B.n497 B.n496 71.676
R631 B.n41 B.n39 71.676
R632 B.n90 B.n42 71.676
R633 B.n94 B.n43 71.676
R634 B.n98 B.n44 71.676
R635 B.n102 B.n45 71.676
R636 B.n106 B.n46 71.676
R637 B.n110 B.n47 71.676
R638 B.n114 B.n48 71.676
R639 B.n118 B.n49 71.676
R640 B.n122 B.n50 71.676
R641 B.n126 B.n51 71.676
R642 B.n130 B.n52 71.676
R643 B.n134 B.n53 71.676
R644 B.n138 B.n54 71.676
R645 B.n142 B.n55 71.676
R646 B.n146 B.n56 71.676
R647 B.n150 B.n57 71.676
R648 B.n154 B.n58 71.676
R649 B.n158 B.n59 71.676
R650 B.n163 B.n60 71.676
R651 B.n167 B.n61 71.676
R652 B.n171 B.n62 71.676
R653 B.n175 B.n63 71.676
R654 B.n179 B.n64 71.676
R655 B.n183 B.n65 71.676
R656 B.n187 B.n66 71.676
R657 B.n191 B.n67 71.676
R658 B.n195 B.n68 71.676
R659 B.n199 B.n69 71.676
R660 B.n203 B.n70 71.676
R661 B.n207 B.n71 71.676
R662 B.n211 B.n72 71.676
R663 B.n215 B.n73 71.676
R664 B.n219 B.n74 71.676
R665 B.n223 B.n75 71.676
R666 B.n227 B.n76 71.676
R667 B.n231 B.n77 71.676
R668 B.n235 B.n78 71.676
R669 B.n239 B.n79 71.676
R670 B.n243 B.n80 71.676
R671 B.n247 B.n81 71.676
R672 B.n82 B.n81 71.676
R673 B.n246 B.n80 71.676
R674 B.n242 B.n79 71.676
R675 B.n238 B.n78 71.676
R676 B.n234 B.n77 71.676
R677 B.n230 B.n76 71.676
R678 B.n226 B.n75 71.676
R679 B.n222 B.n74 71.676
R680 B.n218 B.n73 71.676
R681 B.n214 B.n72 71.676
R682 B.n210 B.n71 71.676
R683 B.n206 B.n70 71.676
R684 B.n202 B.n69 71.676
R685 B.n198 B.n68 71.676
R686 B.n194 B.n67 71.676
R687 B.n190 B.n66 71.676
R688 B.n186 B.n65 71.676
R689 B.n182 B.n64 71.676
R690 B.n178 B.n63 71.676
R691 B.n174 B.n62 71.676
R692 B.n170 B.n61 71.676
R693 B.n166 B.n60 71.676
R694 B.n162 B.n59 71.676
R695 B.n157 B.n58 71.676
R696 B.n153 B.n57 71.676
R697 B.n149 B.n56 71.676
R698 B.n145 B.n55 71.676
R699 B.n141 B.n54 71.676
R700 B.n137 B.n53 71.676
R701 B.n133 B.n52 71.676
R702 B.n129 B.n51 71.676
R703 B.n125 B.n50 71.676
R704 B.n121 B.n49 71.676
R705 B.n117 B.n48 71.676
R706 B.n113 B.n47 71.676
R707 B.n109 B.n46 71.676
R708 B.n105 B.n45 71.676
R709 B.n101 B.n44 71.676
R710 B.n97 B.n43 71.676
R711 B.n93 B.n42 71.676
R712 B.n89 B.n41 71.676
R713 B.n336 B.n335 71.676
R714 B.n342 B.n341 71.676
R715 B.n343 B.n332 71.676
R716 B.n350 B.n349 71.676
R717 B.n351 B.n330 71.676
R718 B.n358 B.n357 71.676
R719 B.n359 B.n328 71.676
R720 B.n366 B.n365 71.676
R721 B.n367 B.n326 71.676
R722 B.n374 B.n373 71.676
R723 B.n375 B.n324 71.676
R724 B.n382 B.n381 71.676
R725 B.n383 B.n322 71.676
R726 B.n390 B.n389 71.676
R727 B.n391 B.n320 71.676
R728 B.n398 B.n397 71.676
R729 B.n399 B.n318 71.676
R730 B.n406 B.n405 71.676
R731 B.n407 B.n313 71.676
R732 B.n414 B.n413 71.676
R733 B.n415 B.n311 71.676
R734 B.n422 B.n421 71.676
R735 B.n423 B.n307 71.676
R736 B.n431 B.n430 71.676
R737 B.n432 B.n305 71.676
R738 B.n439 B.n438 71.676
R739 B.n440 B.n303 71.676
R740 B.n447 B.n446 71.676
R741 B.n448 B.n301 71.676
R742 B.n455 B.n454 71.676
R743 B.n456 B.n299 71.676
R744 B.n463 B.n462 71.676
R745 B.n464 B.n297 71.676
R746 B.n471 B.n470 71.676
R747 B.n472 B.n295 71.676
R748 B.n479 B.n478 71.676
R749 B.n480 B.n293 71.676
R750 B.n487 B.n486 71.676
R751 B.n488 B.n291 71.676
R752 B.n495 B.n494 71.676
R753 B.n496 B.n289 71.676
R754 B.n309 B.t4 70.3833
R755 B.n84 B.t15 70.3833
R756 B.n315 B.t11 70.3706
R757 B.n87 B.t9 70.3706
R758 B.n426 B.n309 59.5399
R759 B.n316 B.n315 59.5399
R760 B.n160 B.n87 59.5399
R761 B.n85 B.n84 59.5399
R762 B.n502 B.n284 47.9646
R763 B.n508 B.n284 47.9646
R764 B.n508 B.n280 47.9646
R765 B.n514 B.n280 47.9646
R766 B.n514 B.n276 47.9646
R767 B.n520 B.n276 47.9646
R768 B.n526 B.n272 47.9646
R769 B.n526 B.n268 47.9646
R770 B.n532 B.n268 47.9646
R771 B.n532 B.n264 47.9646
R772 B.n538 B.n264 47.9646
R773 B.n538 B.n259 47.9646
R774 B.n544 B.n259 47.9646
R775 B.n544 B.n260 47.9646
R776 B.n551 B.n252 47.9646
R777 B.n557 B.n252 47.9646
R778 B.n557 B.n4 47.9646
R779 B.n630 B.n4 47.9646
R780 B.n630 B.n629 47.9646
R781 B.n629 B.n628 47.9646
R782 B.n628 B.n8 47.9646
R783 B.n622 B.n8 47.9646
R784 B.n621 B.n620 47.9646
R785 B.n620 B.n15 47.9646
R786 B.n614 B.n15 47.9646
R787 B.n614 B.n613 47.9646
R788 B.n613 B.n612 47.9646
R789 B.n612 B.n22 47.9646
R790 B.n606 B.n22 47.9646
R791 B.n606 B.n605 47.9646
R792 B.n604 B.n29 47.9646
R793 B.n598 B.n29 47.9646
R794 B.n598 B.n597 47.9646
R795 B.n597 B.n596 47.9646
R796 B.n596 B.n36 47.9646
R797 B.n590 B.n36 47.9646
R798 B.n309 B.n308 38.9823
R799 B.n315 B.n314 38.9823
R800 B.n87 B.n86 38.9823
R801 B.n84 B.n83 38.9823
R802 B.t3 B.n272 32.4468
R803 B.n605 B.t7 32.4468
R804 B.n592 B.n38 31.3761
R805 B.n587 B.n586 31.3761
R806 B.n500 B.n499 31.3761
R807 B.n504 B.n286 31.3761
R808 B.n551 B.t1 26.804
R809 B.n622 B.t0 26.804
R810 B.n260 B.t1 21.1611
R811 B.t0 B.n621 21.1611
R812 B B.n632 18.0485
R813 B.n520 B.t3 15.5183
R814 B.t7 B.n604 15.5183
R815 B.n88 B.n38 10.6151
R816 B.n91 B.n88 10.6151
R817 B.n92 B.n91 10.6151
R818 B.n95 B.n92 10.6151
R819 B.n96 B.n95 10.6151
R820 B.n99 B.n96 10.6151
R821 B.n100 B.n99 10.6151
R822 B.n103 B.n100 10.6151
R823 B.n104 B.n103 10.6151
R824 B.n107 B.n104 10.6151
R825 B.n108 B.n107 10.6151
R826 B.n111 B.n108 10.6151
R827 B.n112 B.n111 10.6151
R828 B.n115 B.n112 10.6151
R829 B.n116 B.n115 10.6151
R830 B.n119 B.n116 10.6151
R831 B.n120 B.n119 10.6151
R832 B.n123 B.n120 10.6151
R833 B.n124 B.n123 10.6151
R834 B.n127 B.n124 10.6151
R835 B.n128 B.n127 10.6151
R836 B.n131 B.n128 10.6151
R837 B.n132 B.n131 10.6151
R838 B.n135 B.n132 10.6151
R839 B.n136 B.n135 10.6151
R840 B.n139 B.n136 10.6151
R841 B.n140 B.n139 10.6151
R842 B.n143 B.n140 10.6151
R843 B.n144 B.n143 10.6151
R844 B.n147 B.n144 10.6151
R845 B.n148 B.n147 10.6151
R846 B.n151 B.n148 10.6151
R847 B.n152 B.n151 10.6151
R848 B.n155 B.n152 10.6151
R849 B.n156 B.n155 10.6151
R850 B.n159 B.n156 10.6151
R851 B.n164 B.n161 10.6151
R852 B.n165 B.n164 10.6151
R853 B.n168 B.n165 10.6151
R854 B.n169 B.n168 10.6151
R855 B.n172 B.n169 10.6151
R856 B.n173 B.n172 10.6151
R857 B.n176 B.n173 10.6151
R858 B.n177 B.n176 10.6151
R859 B.n181 B.n180 10.6151
R860 B.n184 B.n181 10.6151
R861 B.n185 B.n184 10.6151
R862 B.n188 B.n185 10.6151
R863 B.n189 B.n188 10.6151
R864 B.n192 B.n189 10.6151
R865 B.n193 B.n192 10.6151
R866 B.n196 B.n193 10.6151
R867 B.n197 B.n196 10.6151
R868 B.n200 B.n197 10.6151
R869 B.n201 B.n200 10.6151
R870 B.n204 B.n201 10.6151
R871 B.n205 B.n204 10.6151
R872 B.n208 B.n205 10.6151
R873 B.n209 B.n208 10.6151
R874 B.n212 B.n209 10.6151
R875 B.n213 B.n212 10.6151
R876 B.n216 B.n213 10.6151
R877 B.n217 B.n216 10.6151
R878 B.n220 B.n217 10.6151
R879 B.n221 B.n220 10.6151
R880 B.n224 B.n221 10.6151
R881 B.n225 B.n224 10.6151
R882 B.n228 B.n225 10.6151
R883 B.n229 B.n228 10.6151
R884 B.n232 B.n229 10.6151
R885 B.n233 B.n232 10.6151
R886 B.n236 B.n233 10.6151
R887 B.n237 B.n236 10.6151
R888 B.n240 B.n237 10.6151
R889 B.n241 B.n240 10.6151
R890 B.n244 B.n241 10.6151
R891 B.n245 B.n244 10.6151
R892 B.n248 B.n245 10.6151
R893 B.n249 B.n248 10.6151
R894 B.n587 B.n249 10.6151
R895 B.n500 B.n282 10.6151
R896 B.n510 B.n282 10.6151
R897 B.n511 B.n510 10.6151
R898 B.n512 B.n511 10.6151
R899 B.n512 B.n274 10.6151
R900 B.n522 B.n274 10.6151
R901 B.n523 B.n522 10.6151
R902 B.n524 B.n523 10.6151
R903 B.n524 B.n266 10.6151
R904 B.n534 B.n266 10.6151
R905 B.n535 B.n534 10.6151
R906 B.n536 B.n535 10.6151
R907 B.n536 B.n257 10.6151
R908 B.n546 B.n257 10.6151
R909 B.n547 B.n546 10.6151
R910 B.n549 B.n547 10.6151
R911 B.n549 B.n548 10.6151
R912 B.n548 B.n250 10.6151
R913 B.n560 B.n250 10.6151
R914 B.n561 B.n560 10.6151
R915 B.n562 B.n561 10.6151
R916 B.n563 B.n562 10.6151
R917 B.n565 B.n563 10.6151
R918 B.n566 B.n565 10.6151
R919 B.n567 B.n566 10.6151
R920 B.n568 B.n567 10.6151
R921 B.n570 B.n568 10.6151
R922 B.n571 B.n570 10.6151
R923 B.n572 B.n571 10.6151
R924 B.n573 B.n572 10.6151
R925 B.n575 B.n573 10.6151
R926 B.n576 B.n575 10.6151
R927 B.n577 B.n576 10.6151
R928 B.n578 B.n577 10.6151
R929 B.n580 B.n578 10.6151
R930 B.n581 B.n580 10.6151
R931 B.n582 B.n581 10.6151
R932 B.n583 B.n582 10.6151
R933 B.n585 B.n583 10.6151
R934 B.n586 B.n585 10.6151
R935 B.n337 B.n286 10.6151
R936 B.n338 B.n337 10.6151
R937 B.n339 B.n338 10.6151
R938 B.n339 B.n333 10.6151
R939 B.n345 B.n333 10.6151
R940 B.n346 B.n345 10.6151
R941 B.n347 B.n346 10.6151
R942 B.n347 B.n331 10.6151
R943 B.n353 B.n331 10.6151
R944 B.n354 B.n353 10.6151
R945 B.n355 B.n354 10.6151
R946 B.n355 B.n329 10.6151
R947 B.n361 B.n329 10.6151
R948 B.n362 B.n361 10.6151
R949 B.n363 B.n362 10.6151
R950 B.n363 B.n327 10.6151
R951 B.n369 B.n327 10.6151
R952 B.n370 B.n369 10.6151
R953 B.n371 B.n370 10.6151
R954 B.n371 B.n325 10.6151
R955 B.n377 B.n325 10.6151
R956 B.n378 B.n377 10.6151
R957 B.n379 B.n378 10.6151
R958 B.n379 B.n323 10.6151
R959 B.n385 B.n323 10.6151
R960 B.n386 B.n385 10.6151
R961 B.n387 B.n386 10.6151
R962 B.n387 B.n321 10.6151
R963 B.n393 B.n321 10.6151
R964 B.n394 B.n393 10.6151
R965 B.n395 B.n394 10.6151
R966 B.n395 B.n319 10.6151
R967 B.n401 B.n319 10.6151
R968 B.n402 B.n401 10.6151
R969 B.n403 B.n402 10.6151
R970 B.n403 B.n317 10.6151
R971 B.n410 B.n409 10.6151
R972 B.n411 B.n410 10.6151
R973 B.n411 B.n312 10.6151
R974 B.n417 B.n312 10.6151
R975 B.n418 B.n417 10.6151
R976 B.n419 B.n418 10.6151
R977 B.n419 B.n310 10.6151
R978 B.n425 B.n310 10.6151
R979 B.n428 B.n427 10.6151
R980 B.n428 B.n306 10.6151
R981 B.n434 B.n306 10.6151
R982 B.n435 B.n434 10.6151
R983 B.n436 B.n435 10.6151
R984 B.n436 B.n304 10.6151
R985 B.n442 B.n304 10.6151
R986 B.n443 B.n442 10.6151
R987 B.n444 B.n443 10.6151
R988 B.n444 B.n302 10.6151
R989 B.n450 B.n302 10.6151
R990 B.n451 B.n450 10.6151
R991 B.n452 B.n451 10.6151
R992 B.n452 B.n300 10.6151
R993 B.n458 B.n300 10.6151
R994 B.n459 B.n458 10.6151
R995 B.n460 B.n459 10.6151
R996 B.n460 B.n298 10.6151
R997 B.n466 B.n298 10.6151
R998 B.n467 B.n466 10.6151
R999 B.n468 B.n467 10.6151
R1000 B.n468 B.n296 10.6151
R1001 B.n474 B.n296 10.6151
R1002 B.n475 B.n474 10.6151
R1003 B.n476 B.n475 10.6151
R1004 B.n476 B.n294 10.6151
R1005 B.n482 B.n294 10.6151
R1006 B.n483 B.n482 10.6151
R1007 B.n484 B.n483 10.6151
R1008 B.n484 B.n292 10.6151
R1009 B.n490 B.n292 10.6151
R1010 B.n491 B.n490 10.6151
R1011 B.n492 B.n491 10.6151
R1012 B.n492 B.n290 10.6151
R1013 B.n498 B.n290 10.6151
R1014 B.n499 B.n498 10.6151
R1015 B.n505 B.n504 10.6151
R1016 B.n506 B.n505 10.6151
R1017 B.n506 B.n278 10.6151
R1018 B.n516 B.n278 10.6151
R1019 B.n517 B.n516 10.6151
R1020 B.n518 B.n517 10.6151
R1021 B.n518 B.n270 10.6151
R1022 B.n528 B.n270 10.6151
R1023 B.n529 B.n528 10.6151
R1024 B.n530 B.n529 10.6151
R1025 B.n530 B.n262 10.6151
R1026 B.n540 B.n262 10.6151
R1027 B.n541 B.n540 10.6151
R1028 B.n542 B.n541 10.6151
R1029 B.n542 B.n254 10.6151
R1030 B.n553 B.n254 10.6151
R1031 B.n554 B.n553 10.6151
R1032 B.n555 B.n554 10.6151
R1033 B.n555 B.n0 10.6151
R1034 B.n626 B.n1 10.6151
R1035 B.n626 B.n625 10.6151
R1036 B.n625 B.n624 10.6151
R1037 B.n624 B.n10 10.6151
R1038 B.n618 B.n10 10.6151
R1039 B.n618 B.n617 10.6151
R1040 B.n617 B.n616 10.6151
R1041 B.n616 B.n17 10.6151
R1042 B.n610 B.n17 10.6151
R1043 B.n610 B.n609 10.6151
R1044 B.n609 B.n608 10.6151
R1045 B.n608 B.n24 10.6151
R1046 B.n602 B.n24 10.6151
R1047 B.n602 B.n601 10.6151
R1048 B.n601 B.n600 10.6151
R1049 B.n600 B.n31 10.6151
R1050 B.n594 B.n31 10.6151
R1051 B.n594 B.n593 10.6151
R1052 B.n593 B.n592 10.6151
R1053 B.n161 B.n160 6.5566
R1054 B.n177 B.n85 6.5566
R1055 B.n409 B.n316 6.5566
R1056 B.n426 B.n425 6.5566
R1057 B.n160 B.n159 4.05904
R1058 B.n180 B.n85 4.05904
R1059 B.n317 B.n316 4.05904
R1060 B.n427 B.n426 4.05904
R1061 B.n632 B.n0 2.81026
R1062 B.n632 B.n1 2.81026
R1063 VN VN.t1 248.014
R1064 VN VN.t0 207.12
R1065 VTAIL.n1 VTAIL.t3 47.7228
R1066 VTAIL.n3 VTAIL.t2 47.7226
R1067 VTAIL.n0 VTAIL.t1 47.7226
R1068 VTAIL.n2 VTAIL.t0 47.7226
R1069 VTAIL.n1 VTAIL.n0 24.7289
R1070 VTAIL.n3 VTAIL.n2 22.9962
R1071 VTAIL.n2 VTAIL.n1 1.33671
R1072 VTAIL VTAIL.n0 0.961707
R1073 VTAIL VTAIL.n3 0.3755
R1074 VDD2.n0 VDD2.t1 100.422
R1075 VDD2.n0 VDD2.t0 64.4014
R1076 VDD2 VDD2.n0 0.491879
R1077 VP.n0 VP.t1 247.823
R1078 VP.n0 VP.t0 206.88
R1079 VP VP.n0 0.241678
R1080 VDD1 VDD1.t1 101.38
R1081 VDD1 VDD1.t0 64.8927
C0 VTAIL VP 1.92903f
C1 VN VDD2 2.23895f
C2 VDD1 VDD2 0.566202f
C3 VDD1 VN 0.147366f
C4 VP VDD2 0.294002f
C5 VN VP 4.71832f
C6 VDD1 VP 2.38283f
C7 VTAIL VDD2 4.59367f
C8 VN VTAIL 1.91468f
C9 VDD1 VTAIL 4.54998f
C10 VDD2 B 3.805323f
C11 VDD1 B 6.59173f
C12 VTAIL B 6.207837f
C13 VN B 8.51641f
C14 VP B 5.13917f
C15 VDD1.t0 B 1.86071f
C16 VDD1.t1 B 2.34105f
C17 VP.t1 B 2.00608f
C18 VP.t0 B 1.70328f
C19 VP.n0 B 3.34504f
C20 VDD2.t1 B 2.30332f
C21 VDD2.t0 B 1.85192f
C22 VDD2.n0 B 2.55579f
C23 VTAIL.t1 B 1.28302f
C24 VTAIL.n0 B 1.01508f
C25 VTAIL.t3 B 1.28302f
C26 VTAIL.n1 B 1.0327f
C27 VTAIL.t0 B 1.28302f
C28 VTAIL.n2 B 0.951261f
C29 VTAIL.t2 B 1.28302f
C30 VTAIL.n3 B 0.90608f
C31 VN.t0 B 1.64553f
C32 VN.t1 B 1.94083f
.ends

