* NGSPICE file created from diff_pair_sample_1217.ext - technology: sky130A

.subckt diff_pair_sample_1217 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=0.64
X1 VTAIL.t7 VP.t0 VDD1.t0 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=2.1747 ps=13.51 w=13.18 l=0.64
X2 B.t8 B.t6 B.t7 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=0.64
X3 VDD2.t3 VN.t0 VTAIL.t0 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=2.1747 pd=13.51 as=5.1402 ps=27.14 w=13.18 l=0.64
X4 VDD1.t1 VP.t1 VTAIL.t6 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=2.1747 pd=13.51 as=5.1402 ps=27.14 w=13.18 l=0.64
X5 VDD1.t2 VP.t2 VTAIL.t5 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=2.1747 pd=13.51 as=5.1402 ps=27.14 w=13.18 l=0.64
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=2.1747 pd=13.51 as=5.1402 ps=27.14 w=13.18 l=0.64
X7 VTAIL.t2 VN.t2 VDD2.t1 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=2.1747 ps=13.51 w=13.18 l=0.64
X8 B.t5 B.t3 B.t4 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=0.64
X9 VTAIL.t3 VN.t3 VDD2.t0 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=2.1747 ps=13.51 w=13.18 l=0.64
X10 VTAIL.t4 VP.t3 VDD1.t3 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=2.1747 ps=13.51 w=13.18 l=0.64
X11 B.t2 B.t0 B.t1 w_n1552_n3604# sky130_fd_pr__pfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=0.64
R0 B.n230 B.t6 700.082
R1 B.n105 B.t9 700.082
R2 B.n41 B.t0 700.082
R3 B.n34 B.t3 700.082
R4 B.n317 B.n82 585
R5 B.n316 B.n315 585
R6 B.n314 B.n83 585
R7 B.n313 B.n312 585
R8 B.n311 B.n84 585
R9 B.n310 B.n309 585
R10 B.n308 B.n85 585
R11 B.n307 B.n306 585
R12 B.n305 B.n86 585
R13 B.n304 B.n303 585
R14 B.n302 B.n87 585
R15 B.n301 B.n300 585
R16 B.n299 B.n88 585
R17 B.n298 B.n297 585
R18 B.n296 B.n89 585
R19 B.n295 B.n294 585
R20 B.n293 B.n90 585
R21 B.n292 B.n291 585
R22 B.n290 B.n91 585
R23 B.n289 B.n288 585
R24 B.n287 B.n92 585
R25 B.n286 B.n285 585
R26 B.n284 B.n93 585
R27 B.n283 B.n282 585
R28 B.n281 B.n94 585
R29 B.n280 B.n279 585
R30 B.n278 B.n95 585
R31 B.n277 B.n276 585
R32 B.n275 B.n96 585
R33 B.n274 B.n273 585
R34 B.n272 B.n97 585
R35 B.n271 B.n270 585
R36 B.n269 B.n98 585
R37 B.n268 B.n267 585
R38 B.n266 B.n99 585
R39 B.n265 B.n264 585
R40 B.n263 B.n100 585
R41 B.n262 B.n261 585
R42 B.n260 B.n101 585
R43 B.n259 B.n258 585
R44 B.n257 B.n102 585
R45 B.n256 B.n255 585
R46 B.n254 B.n103 585
R47 B.n253 B.n252 585
R48 B.n251 B.n104 585
R49 B.n249 B.n248 585
R50 B.n247 B.n107 585
R51 B.n246 B.n245 585
R52 B.n244 B.n108 585
R53 B.n243 B.n242 585
R54 B.n241 B.n109 585
R55 B.n240 B.n239 585
R56 B.n238 B.n110 585
R57 B.n237 B.n236 585
R58 B.n235 B.n111 585
R59 B.n234 B.n233 585
R60 B.n229 B.n112 585
R61 B.n228 B.n227 585
R62 B.n226 B.n113 585
R63 B.n225 B.n224 585
R64 B.n223 B.n114 585
R65 B.n222 B.n221 585
R66 B.n220 B.n115 585
R67 B.n219 B.n218 585
R68 B.n217 B.n116 585
R69 B.n216 B.n215 585
R70 B.n214 B.n117 585
R71 B.n213 B.n212 585
R72 B.n211 B.n118 585
R73 B.n210 B.n209 585
R74 B.n208 B.n119 585
R75 B.n207 B.n206 585
R76 B.n205 B.n120 585
R77 B.n204 B.n203 585
R78 B.n202 B.n121 585
R79 B.n201 B.n200 585
R80 B.n199 B.n122 585
R81 B.n198 B.n197 585
R82 B.n196 B.n123 585
R83 B.n195 B.n194 585
R84 B.n193 B.n124 585
R85 B.n192 B.n191 585
R86 B.n190 B.n125 585
R87 B.n189 B.n188 585
R88 B.n187 B.n126 585
R89 B.n186 B.n185 585
R90 B.n184 B.n127 585
R91 B.n183 B.n182 585
R92 B.n181 B.n128 585
R93 B.n180 B.n179 585
R94 B.n178 B.n129 585
R95 B.n177 B.n176 585
R96 B.n175 B.n130 585
R97 B.n174 B.n173 585
R98 B.n172 B.n131 585
R99 B.n171 B.n170 585
R100 B.n169 B.n132 585
R101 B.n168 B.n167 585
R102 B.n166 B.n133 585
R103 B.n165 B.n164 585
R104 B.n319 B.n318 585
R105 B.n320 B.n81 585
R106 B.n322 B.n321 585
R107 B.n323 B.n80 585
R108 B.n325 B.n324 585
R109 B.n326 B.n79 585
R110 B.n328 B.n327 585
R111 B.n329 B.n78 585
R112 B.n331 B.n330 585
R113 B.n332 B.n77 585
R114 B.n334 B.n333 585
R115 B.n335 B.n76 585
R116 B.n337 B.n336 585
R117 B.n338 B.n75 585
R118 B.n340 B.n339 585
R119 B.n341 B.n74 585
R120 B.n343 B.n342 585
R121 B.n344 B.n73 585
R122 B.n346 B.n345 585
R123 B.n347 B.n72 585
R124 B.n349 B.n348 585
R125 B.n350 B.n71 585
R126 B.n352 B.n351 585
R127 B.n353 B.n70 585
R128 B.n355 B.n354 585
R129 B.n356 B.n69 585
R130 B.n358 B.n357 585
R131 B.n359 B.n68 585
R132 B.n361 B.n360 585
R133 B.n362 B.n67 585
R134 B.n364 B.n363 585
R135 B.n365 B.n66 585
R136 B.n367 B.n366 585
R137 B.n368 B.n65 585
R138 B.n519 B.n10 585
R139 B.n518 B.n517 585
R140 B.n516 B.n11 585
R141 B.n515 B.n514 585
R142 B.n513 B.n12 585
R143 B.n512 B.n511 585
R144 B.n510 B.n13 585
R145 B.n509 B.n508 585
R146 B.n507 B.n14 585
R147 B.n506 B.n505 585
R148 B.n504 B.n15 585
R149 B.n503 B.n502 585
R150 B.n501 B.n16 585
R151 B.n500 B.n499 585
R152 B.n498 B.n17 585
R153 B.n497 B.n496 585
R154 B.n495 B.n18 585
R155 B.n494 B.n493 585
R156 B.n492 B.n19 585
R157 B.n491 B.n490 585
R158 B.n489 B.n20 585
R159 B.n488 B.n487 585
R160 B.n486 B.n21 585
R161 B.n485 B.n484 585
R162 B.n483 B.n22 585
R163 B.n482 B.n481 585
R164 B.n480 B.n23 585
R165 B.n479 B.n478 585
R166 B.n477 B.n24 585
R167 B.n476 B.n475 585
R168 B.n474 B.n25 585
R169 B.n473 B.n472 585
R170 B.n471 B.n26 585
R171 B.n470 B.n469 585
R172 B.n468 B.n27 585
R173 B.n467 B.n466 585
R174 B.n465 B.n28 585
R175 B.n464 B.n463 585
R176 B.n462 B.n29 585
R177 B.n461 B.n460 585
R178 B.n459 B.n30 585
R179 B.n458 B.n457 585
R180 B.n456 B.n31 585
R181 B.n455 B.n454 585
R182 B.n453 B.n32 585
R183 B.n452 B.n451 585
R184 B.n450 B.n33 585
R185 B.n449 B.n448 585
R186 B.n447 B.n37 585
R187 B.n446 B.n445 585
R188 B.n444 B.n38 585
R189 B.n443 B.n442 585
R190 B.n441 B.n39 585
R191 B.n440 B.n439 585
R192 B.n438 B.n40 585
R193 B.n436 B.n435 585
R194 B.n434 B.n43 585
R195 B.n433 B.n432 585
R196 B.n431 B.n44 585
R197 B.n430 B.n429 585
R198 B.n428 B.n45 585
R199 B.n427 B.n426 585
R200 B.n425 B.n46 585
R201 B.n424 B.n423 585
R202 B.n422 B.n47 585
R203 B.n421 B.n420 585
R204 B.n419 B.n48 585
R205 B.n418 B.n417 585
R206 B.n416 B.n49 585
R207 B.n415 B.n414 585
R208 B.n413 B.n50 585
R209 B.n412 B.n411 585
R210 B.n410 B.n51 585
R211 B.n409 B.n408 585
R212 B.n407 B.n52 585
R213 B.n406 B.n405 585
R214 B.n404 B.n53 585
R215 B.n403 B.n402 585
R216 B.n401 B.n54 585
R217 B.n400 B.n399 585
R218 B.n398 B.n55 585
R219 B.n397 B.n396 585
R220 B.n395 B.n56 585
R221 B.n394 B.n393 585
R222 B.n392 B.n57 585
R223 B.n391 B.n390 585
R224 B.n389 B.n58 585
R225 B.n388 B.n387 585
R226 B.n386 B.n59 585
R227 B.n385 B.n384 585
R228 B.n383 B.n60 585
R229 B.n382 B.n381 585
R230 B.n380 B.n61 585
R231 B.n379 B.n378 585
R232 B.n377 B.n62 585
R233 B.n376 B.n375 585
R234 B.n374 B.n63 585
R235 B.n373 B.n372 585
R236 B.n371 B.n64 585
R237 B.n370 B.n369 585
R238 B.n521 B.n520 585
R239 B.n522 B.n9 585
R240 B.n524 B.n523 585
R241 B.n525 B.n8 585
R242 B.n527 B.n526 585
R243 B.n528 B.n7 585
R244 B.n530 B.n529 585
R245 B.n531 B.n6 585
R246 B.n533 B.n532 585
R247 B.n534 B.n5 585
R248 B.n536 B.n535 585
R249 B.n537 B.n4 585
R250 B.n539 B.n538 585
R251 B.n540 B.n3 585
R252 B.n542 B.n541 585
R253 B.n543 B.n0 585
R254 B.n2 B.n1 585
R255 B.n142 B.n141 585
R256 B.n144 B.n143 585
R257 B.n145 B.n140 585
R258 B.n147 B.n146 585
R259 B.n148 B.n139 585
R260 B.n150 B.n149 585
R261 B.n151 B.n138 585
R262 B.n153 B.n152 585
R263 B.n154 B.n137 585
R264 B.n156 B.n155 585
R265 B.n157 B.n136 585
R266 B.n159 B.n158 585
R267 B.n160 B.n135 585
R268 B.n162 B.n161 585
R269 B.n163 B.n134 585
R270 B.n165 B.n134 506.916
R271 B.n319 B.n82 506.916
R272 B.n369 B.n368 506.916
R273 B.n520 B.n519 506.916
R274 B.n545 B.n544 256.663
R275 B.n544 B.n543 235.042
R276 B.n544 B.n2 235.042
R277 B.n166 B.n165 163.367
R278 B.n167 B.n166 163.367
R279 B.n167 B.n132 163.367
R280 B.n171 B.n132 163.367
R281 B.n172 B.n171 163.367
R282 B.n173 B.n172 163.367
R283 B.n173 B.n130 163.367
R284 B.n177 B.n130 163.367
R285 B.n178 B.n177 163.367
R286 B.n179 B.n178 163.367
R287 B.n179 B.n128 163.367
R288 B.n183 B.n128 163.367
R289 B.n184 B.n183 163.367
R290 B.n185 B.n184 163.367
R291 B.n185 B.n126 163.367
R292 B.n189 B.n126 163.367
R293 B.n190 B.n189 163.367
R294 B.n191 B.n190 163.367
R295 B.n191 B.n124 163.367
R296 B.n195 B.n124 163.367
R297 B.n196 B.n195 163.367
R298 B.n197 B.n196 163.367
R299 B.n197 B.n122 163.367
R300 B.n201 B.n122 163.367
R301 B.n202 B.n201 163.367
R302 B.n203 B.n202 163.367
R303 B.n203 B.n120 163.367
R304 B.n207 B.n120 163.367
R305 B.n208 B.n207 163.367
R306 B.n209 B.n208 163.367
R307 B.n209 B.n118 163.367
R308 B.n213 B.n118 163.367
R309 B.n214 B.n213 163.367
R310 B.n215 B.n214 163.367
R311 B.n215 B.n116 163.367
R312 B.n219 B.n116 163.367
R313 B.n220 B.n219 163.367
R314 B.n221 B.n220 163.367
R315 B.n221 B.n114 163.367
R316 B.n225 B.n114 163.367
R317 B.n226 B.n225 163.367
R318 B.n227 B.n226 163.367
R319 B.n227 B.n112 163.367
R320 B.n234 B.n112 163.367
R321 B.n235 B.n234 163.367
R322 B.n236 B.n235 163.367
R323 B.n236 B.n110 163.367
R324 B.n240 B.n110 163.367
R325 B.n241 B.n240 163.367
R326 B.n242 B.n241 163.367
R327 B.n242 B.n108 163.367
R328 B.n246 B.n108 163.367
R329 B.n247 B.n246 163.367
R330 B.n248 B.n247 163.367
R331 B.n248 B.n104 163.367
R332 B.n253 B.n104 163.367
R333 B.n254 B.n253 163.367
R334 B.n255 B.n254 163.367
R335 B.n255 B.n102 163.367
R336 B.n259 B.n102 163.367
R337 B.n260 B.n259 163.367
R338 B.n261 B.n260 163.367
R339 B.n261 B.n100 163.367
R340 B.n265 B.n100 163.367
R341 B.n266 B.n265 163.367
R342 B.n267 B.n266 163.367
R343 B.n267 B.n98 163.367
R344 B.n271 B.n98 163.367
R345 B.n272 B.n271 163.367
R346 B.n273 B.n272 163.367
R347 B.n273 B.n96 163.367
R348 B.n277 B.n96 163.367
R349 B.n278 B.n277 163.367
R350 B.n279 B.n278 163.367
R351 B.n279 B.n94 163.367
R352 B.n283 B.n94 163.367
R353 B.n284 B.n283 163.367
R354 B.n285 B.n284 163.367
R355 B.n285 B.n92 163.367
R356 B.n289 B.n92 163.367
R357 B.n290 B.n289 163.367
R358 B.n291 B.n290 163.367
R359 B.n291 B.n90 163.367
R360 B.n295 B.n90 163.367
R361 B.n296 B.n295 163.367
R362 B.n297 B.n296 163.367
R363 B.n297 B.n88 163.367
R364 B.n301 B.n88 163.367
R365 B.n302 B.n301 163.367
R366 B.n303 B.n302 163.367
R367 B.n303 B.n86 163.367
R368 B.n307 B.n86 163.367
R369 B.n308 B.n307 163.367
R370 B.n309 B.n308 163.367
R371 B.n309 B.n84 163.367
R372 B.n313 B.n84 163.367
R373 B.n314 B.n313 163.367
R374 B.n315 B.n314 163.367
R375 B.n315 B.n82 163.367
R376 B.n368 B.n367 163.367
R377 B.n367 B.n66 163.367
R378 B.n363 B.n66 163.367
R379 B.n363 B.n362 163.367
R380 B.n362 B.n361 163.367
R381 B.n361 B.n68 163.367
R382 B.n357 B.n68 163.367
R383 B.n357 B.n356 163.367
R384 B.n356 B.n355 163.367
R385 B.n355 B.n70 163.367
R386 B.n351 B.n70 163.367
R387 B.n351 B.n350 163.367
R388 B.n350 B.n349 163.367
R389 B.n349 B.n72 163.367
R390 B.n345 B.n72 163.367
R391 B.n345 B.n344 163.367
R392 B.n344 B.n343 163.367
R393 B.n343 B.n74 163.367
R394 B.n339 B.n74 163.367
R395 B.n339 B.n338 163.367
R396 B.n338 B.n337 163.367
R397 B.n337 B.n76 163.367
R398 B.n333 B.n76 163.367
R399 B.n333 B.n332 163.367
R400 B.n332 B.n331 163.367
R401 B.n331 B.n78 163.367
R402 B.n327 B.n78 163.367
R403 B.n327 B.n326 163.367
R404 B.n326 B.n325 163.367
R405 B.n325 B.n80 163.367
R406 B.n321 B.n80 163.367
R407 B.n321 B.n320 163.367
R408 B.n320 B.n319 163.367
R409 B.n519 B.n518 163.367
R410 B.n518 B.n11 163.367
R411 B.n514 B.n11 163.367
R412 B.n514 B.n513 163.367
R413 B.n513 B.n512 163.367
R414 B.n512 B.n13 163.367
R415 B.n508 B.n13 163.367
R416 B.n508 B.n507 163.367
R417 B.n507 B.n506 163.367
R418 B.n506 B.n15 163.367
R419 B.n502 B.n15 163.367
R420 B.n502 B.n501 163.367
R421 B.n501 B.n500 163.367
R422 B.n500 B.n17 163.367
R423 B.n496 B.n17 163.367
R424 B.n496 B.n495 163.367
R425 B.n495 B.n494 163.367
R426 B.n494 B.n19 163.367
R427 B.n490 B.n19 163.367
R428 B.n490 B.n489 163.367
R429 B.n489 B.n488 163.367
R430 B.n488 B.n21 163.367
R431 B.n484 B.n21 163.367
R432 B.n484 B.n483 163.367
R433 B.n483 B.n482 163.367
R434 B.n482 B.n23 163.367
R435 B.n478 B.n23 163.367
R436 B.n478 B.n477 163.367
R437 B.n477 B.n476 163.367
R438 B.n476 B.n25 163.367
R439 B.n472 B.n25 163.367
R440 B.n472 B.n471 163.367
R441 B.n471 B.n470 163.367
R442 B.n470 B.n27 163.367
R443 B.n466 B.n27 163.367
R444 B.n466 B.n465 163.367
R445 B.n465 B.n464 163.367
R446 B.n464 B.n29 163.367
R447 B.n460 B.n29 163.367
R448 B.n460 B.n459 163.367
R449 B.n459 B.n458 163.367
R450 B.n458 B.n31 163.367
R451 B.n454 B.n31 163.367
R452 B.n454 B.n453 163.367
R453 B.n453 B.n452 163.367
R454 B.n452 B.n33 163.367
R455 B.n448 B.n33 163.367
R456 B.n448 B.n447 163.367
R457 B.n447 B.n446 163.367
R458 B.n446 B.n38 163.367
R459 B.n442 B.n38 163.367
R460 B.n442 B.n441 163.367
R461 B.n441 B.n440 163.367
R462 B.n440 B.n40 163.367
R463 B.n435 B.n40 163.367
R464 B.n435 B.n434 163.367
R465 B.n434 B.n433 163.367
R466 B.n433 B.n44 163.367
R467 B.n429 B.n44 163.367
R468 B.n429 B.n428 163.367
R469 B.n428 B.n427 163.367
R470 B.n427 B.n46 163.367
R471 B.n423 B.n46 163.367
R472 B.n423 B.n422 163.367
R473 B.n422 B.n421 163.367
R474 B.n421 B.n48 163.367
R475 B.n417 B.n48 163.367
R476 B.n417 B.n416 163.367
R477 B.n416 B.n415 163.367
R478 B.n415 B.n50 163.367
R479 B.n411 B.n50 163.367
R480 B.n411 B.n410 163.367
R481 B.n410 B.n409 163.367
R482 B.n409 B.n52 163.367
R483 B.n405 B.n52 163.367
R484 B.n405 B.n404 163.367
R485 B.n404 B.n403 163.367
R486 B.n403 B.n54 163.367
R487 B.n399 B.n54 163.367
R488 B.n399 B.n398 163.367
R489 B.n398 B.n397 163.367
R490 B.n397 B.n56 163.367
R491 B.n393 B.n56 163.367
R492 B.n393 B.n392 163.367
R493 B.n392 B.n391 163.367
R494 B.n391 B.n58 163.367
R495 B.n387 B.n58 163.367
R496 B.n387 B.n386 163.367
R497 B.n386 B.n385 163.367
R498 B.n385 B.n60 163.367
R499 B.n381 B.n60 163.367
R500 B.n381 B.n380 163.367
R501 B.n380 B.n379 163.367
R502 B.n379 B.n62 163.367
R503 B.n375 B.n62 163.367
R504 B.n375 B.n374 163.367
R505 B.n374 B.n373 163.367
R506 B.n373 B.n64 163.367
R507 B.n369 B.n64 163.367
R508 B.n520 B.n9 163.367
R509 B.n524 B.n9 163.367
R510 B.n525 B.n524 163.367
R511 B.n526 B.n525 163.367
R512 B.n526 B.n7 163.367
R513 B.n530 B.n7 163.367
R514 B.n531 B.n530 163.367
R515 B.n532 B.n531 163.367
R516 B.n532 B.n5 163.367
R517 B.n536 B.n5 163.367
R518 B.n537 B.n536 163.367
R519 B.n538 B.n537 163.367
R520 B.n538 B.n3 163.367
R521 B.n542 B.n3 163.367
R522 B.n543 B.n542 163.367
R523 B.n142 B.n2 163.367
R524 B.n143 B.n142 163.367
R525 B.n143 B.n140 163.367
R526 B.n147 B.n140 163.367
R527 B.n148 B.n147 163.367
R528 B.n149 B.n148 163.367
R529 B.n149 B.n138 163.367
R530 B.n153 B.n138 163.367
R531 B.n154 B.n153 163.367
R532 B.n155 B.n154 163.367
R533 B.n155 B.n136 163.367
R534 B.n159 B.n136 163.367
R535 B.n160 B.n159 163.367
R536 B.n161 B.n160 163.367
R537 B.n161 B.n134 163.367
R538 B.n105 B.t10 130.714
R539 B.n41 B.t2 130.714
R540 B.n230 B.t7 130.698
R541 B.n34 B.t5 130.698
R542 B.n106 B.t11 111.903
R543 B.n42 B.t1 111.903
R544 B.n231 B.t8 111.886
R545 B.n35 B.t4 111.886
R546 B.n232 B.n231 59.5399
R547 B.n250 B.n106 59.5399
R548 B.n437 B.n42 59.5399
R549 B.n36 B.n35 59.5399
R550 B.n521 B.n10 32.9371
R551 B.n370 B.n65 32.9371
R552 B.n318 B.n317 32.9371
R553 B.n164 B.n163 32.9371
R554 B.n231 B.n230 18.8126
R555 B.n106 B.n105 18.8126
R556 B.n42 B.n41 18.8126
R557 B.n35 B.n34 18.8126
R558 B B.n545 18.0485
R559 B.n522 B.n521 10.6151
R560 B.n523 B.n522 10.6151
R561 B.n523 B.n8 10.6151
R562 B.n527 B.n8 10.6151
R563 B.n528 B.n527 10.6151
R564 B.n529 B.n528 10.6151
R565 B.n529 B.n6 10.6151
R566 B.n533 B.n6 10.6151
R567 B.n534 B.n533 10.6151
R568 B.n535 B.n534 10.6151
R569 B.n535 B.n4 10.6151
R570 B.n539 B.n4 10.6151
R571 B.n540 B.n539 10.6151
R572 B.n541 B.n540 10.6151
R573 B.n541 B.n0 10.6151
R574 B.n517 B.n10 10.6151
R575 B.n517 B.n516 10.6151
R576 B.n516 B.n515 10.6151
R577 B.n515 B.n12 10.6151
R578 B.n511 B.n12 10.6151
R579 B.n511 B.n510 10.6151
R580 B.n510 B.n509 10.6151
R581 B.n509 B.n14 10.6151
R582 B.n505 B.n14 10.6151
R583 B.n505 B.n504 10.6151
R584 B.n504 B.n503 10.6151
R585 B.n503 B.n16 10.6151
R586 B.n499 B.n16 10.6151
R587 B.n499 B.n498 10.6151
R588 B.n498 B.n497 10.6151
R589 B.n497 B.n18 10.6151
R590 B.n493 B.n18 10.6151
R591 B.n493 B.n492 10.6151
R592 B.n492 B.n491 10.6151
R593 B.n491 B.n20 10.6151
R594 B.n487 B.n20 10.6151
R595 B.n487 B.n486 10.6151
R596 B.n486 B.n485 10.6151
R597 B.n485 B.n22 10.6151
R598 B.n481 B.n22 10.6151
R599 B.n481 B.n480 10.6151
R600 B.n480 B.n479 10.6151
R601 B.n479 B.n24 10.6151
R602 B.n475 B.n24 10.6151
R603 B.n475 B.n474 10.6151
R604 B.n474 B.n473 10.6151
R605 B.n473 B.n26 10.6151
R606 B.n469 B.n26 10.6151
R607 B.n469 B.n468 10.6151
R608 B.n468 B.n467 10.6151
R609 B.n467 B.n28 10.6151
R610 B.n463 B.n28 10.6151
R611 B.n463 B.n462 10.6151
R612 B.n462 B.n461 10.6151
R613 B.n461 B.n30 10.6151
R614 B.n457 B.n30 10.6151
R615 B.n457 B.n456 10.6151
R616 B.n456 B.n455 10.6151
R617 B.n455 B.n32 10.6151
R618 B.n451 B.n450 10.6151
R619 B.n450 B.n449 10.6151
R620 B.n449 B.n37 10.6151
R621 B.n445 B.n37 10.6151
R622 B.n445 B.n444 10.6151
R623 B.n444 B.n443 10.6151
R624 B.n443 B.n39 10.6151
R625 B.n439 B.n39 10.6151
R626 B.n439 B.n438 10.6151
R627 B.n436 B.n43 10.6151
R628 B.n432 B.n43 10.6151
R629 B.n432 B.n431 10.6151
R630 B.n431 B.n430 10.6151
R631 B.n430 B.n45 10.6151
R632 B.n426 B.n45 10.6151
R633 B.n426 B.n425 10.6151
R634 B.n425 B.n424 10.6151
R635 B.n424 B.n47 10.6151
R636 B.n420 B.n47 10.6151
R637 B.n420 B.n419 10.6151
R638 B.n419 B.n418 10.6151
R639 B.n418 B.n49 10.6151
R640 B.n414 B.n49 10.6151
R641 B.n414 B.n413 10.6151
R642 B.n413 B.n412 10.6151
R643 B.n412 B.n51 10.6151
R644 B.n408 B.n51 10.6151
R645 B.n408 B.n407 10.6151
R646 B.n407 B.n406 10.6151
R647 B.n406 B.n53 10.6151
R648 B.n402 B.n53 10.6151
R649 B.n402 B.n401 10.6151
R650 B.n401 B.n400 10.6151
R651 B.n400 B.n55 10.6151
R652 B.n396 B.n55 10.6151
R653 B.n396 B.n395 10.6151
R654 B.n395 B.n394 10.6151
R655 B.n394 B.n57 10.6151
R656 B.n390 B.n57 10.6151
R657 B.n390 B.n389 10.6151
R658 B.n389 B.n388 10.6151
R659 B.n388 B.n59 10.6151
R660 B.n384 B.n59 10.6151
R661 B.n384 B.n383 10.6151
R662 B.n383 B.n382 10.6151
R663 B.n382 B.n61 10.6151
R664 B.n378 B.n61 10.6151
R665 B.n378 B.n377 10.6151
R666 B.n377 B.n376 10.6151
R667 B.n376 B.n63 10.6151
R668 B.n372 B.n63 10.6151
R669 B.n372 B.n371 10.6151
R670 B.n371 B.n370 10.6151
R671 B.n366 B.n65 10.6151
R672 B.n366 B.n365 10.6151
R673 B.n365 B.n364 10.6151
R674 B.n364 B.n67 10.6151
R675 B.n360 B.n67 10.6151
R676 B.n360 B.n359 10.6151
R677 B.n359 B.n358 10.6151
R678 B.n358 B.n69 10.6151
R679 B.n354 B.n69 10.6151
R680 B.n354 B.n353 10.6151
R681 B.n353 B.n352 10.6151
R682 B.n352 B.n71 10.6151
R683 B.n348 B.n71 10.6151
R684 B.n348 B.n347 10.6151
R685 B.n347 B.n346 10.6151
R686 B.n346 B.n73 10.6151
R687 B.n342 B.n73 10.6151
R688 B.n342 B.n341 10.6151
R689 B.n341 B.n340 10.6151
R690 B.n340 B.n75 10.6151
R691 B.n336 B.n75 10.6151
R692 B.n336 B.n335 10.6151
R693 B.n335 B.n334 10.6151
R694 B.n334 B.n77 10.6151
R695 B.n330 B.n77 10.6151
R696 B.n330 B.n329 10.6151
R697 B.n329 B.n328 10.6151
R698 B.n328 B.n79 10.6151
R699 B.n324 B.n79 10.6151
R700 B.n324 B.n323 10.6151
R701 B.n323 B.n322 10.6151
R702 B.n322 B.n81 10.6151
R703 B.n318 B.n81 10.6151
R704 B.n141 B.n1 10.6151
R705 B.n144 B.n141 10.6151
R706 B.n145 B.n144 10.6151
R707 B.n146 B.n145 10.6151
R708 B.n146 B.n139 10.6151
R709 B.n150 B.n139 10.6151
R710 B.n151 B.n150 10.6151
R711 B.n152 B.n151 10.6151
R712 B.n152 B.n137 10.6151
R713 B.n156 B.n137 10.6151
R714 B.n157 B.n156 10.6151
R715 B.n158 B.n157 10.6151
R716 B.n158 B.n135 10.6151
R717 B.n162 B.n135 10.6151
R718 B.n163 B.n162 10.6151
R719 B.n164 B.n133 10.6151
R720 B.n168 B.n133 10.6151
R721 B.n169 B.n168 10.6151
R722 B.n170 B.n169 10.6151
R723 B.n170 B.n131 10.6151
R724 B.n174 B.n131 10.6151
R725 B.n175 B.n174 10.6151
R726 B.n176 B.n175 10.6151
R727 B.n176 B.n129 10.6151
R728 B.n180 B.n129 10.6151
R729 B.n181 B.n180 10.6151
R730 B.n182 B.n181 10.6151
R731 B.n182 B.n127 10.6151
R732 B.n186 B.n127 10.6151
R733 B.n187 B.n186 10.6151
R734 B.n188 B.n187 10.6151
R735 B.n188 B.n125 10.6151
R736 B.n192 B.n125 10.6151
R737 B.n193 B.n192 10.6151
R738 B.n194 B.n193 10.6151
R739 B.n194 B.n123 10.6151
R740 B.n198 B.n123 10.6151
R741 B.n199 B.n198 10.6151
R742 B.n200 B.n199 10.6151
R743 B.n200 B.n121 10.6151
R744 B.n204 B.n121 10.6151
R745 B.n205 B.n204 10.6151
R746 B.n206 B.n205 10.6151
R747 B.n206 B.n119 10.6151
R748 B.n210 B.n119 10.6151
R749 B.n211 B.n210 10.6151
R750 B.n212 B.n211 10.6151
R751 B.n212 B.n117 10.6151
R752 B.n216 B.n117 10.6151
R753 B.n217 B.n216 10.6151
R754 B.n218 B.n217 10.6151
R755 B.n218 B.n115 10.6151
R756 B.n222 B.n115 10.6151
R757 B.n223 B.n222 10.6151
R758 B.n224 B.n223 10.6151
R759 B.n224 B.n113 10.6151
R760 B.n228 B.n113 10.6151
R761 B.n229 B.n228 10.6151
R762 B.n233 B.n229 10.6151
R763 B.n237 B.n111 10.6151
R764 B.n238 B.n237 10.6151
R765 B.n239 B.n238 10.6151
R766 B.n239 B.n109 10.6151
R767 B.n243 B.n109 10.6151
R768 B.n244 B.n243 10.6151
R769 B.n245 B.n244 10.6151
R770 B.n245 B.n107 10.6151
R771 B.n249 B.n107 10.6151
R772 B.n252 B.n251 10.6151
R773 B.n252 B.n103 10.6151
R774 B.n256 B.n103 10.6151
R775 B.n257 B.n256 10.6151
R776 B.n258 B.n257 10.6151
R777 B.n258 B.n101 10.6151
R778 B.n262 B.n101 10.6151
R779 B.n263 B.n262 10.6151
R780 B.n264 B.n263 10.6151
R781 B.n264 B.n99 10.6151
R782 B.n268 B.n99 10.6151
R783 B.n269 B.n268 10.6151
R784 B.n270 B.n269 10.6151
R785 B.n270 B.n97 10.6151
R786 B.n274 B.n97 10.6151
R787 B.n275 B.n274 10.6151
R788 B.n276 B.n275 10.6151
R789 B.n276 B.n95 10.6151
R790 B.n280 B.n95 10.6151
R791 B.n281 B.n280 10.6151
R792 B.n282 B.n281 10.6151
R793 B.n282 B.n93 10.6151
R794 B.n286 B.n93 10.6151
R795 B.n287 B.n286 10.6151
R796 B.n288 B.n287 10.6151
R797 B.n288 B.n91 10.6151
R798 B.n292 B.n91 10.6151
R799 B.n293 B.n292 10.6151
R800 B.n294 B.n293 10.6151
R801 B.n294 B.n89 10.6151
R802 B.n298 B.n89 10.6151
R803 B.n299 B.n298 10.6151
R804 B.n300 B.n299 10.6151
R805 B.n300 B.n87 10.6151
R806 B.n304 B.n87 10.6151
R807 B.n305 B.n304 10.6151
R808 B.n306 B.n305 10.6151
R809 B.n306 B.n85 10.6151
R810 B.n310 B.n85 10.6151
R811 B.n311 B.n310 10.6151
R812 B.n312 B.n311 10.6151
R813 B.n312 B.n83 10.6151
R814 B.n316 B.n83 10.6151
R815 B.n317 B.n316 10.6151
R816 B.n36 B.n32 9.36635
R817 B.n437 B.n436 9.36635
R818 B.n233 B.n232 9.36635
R819 B.n251 B.n250 9.36635
R820 B.n545 B.n0 8.11757
R821 B.n545 B.n1 8.11757
R822 B.n451 B.n36 1.24928
R823 B.n438 B.n437 1.24928
R824 B.n232 B.n111 1.24928
R825 B.n250 B.n249 1.24928
R826 VP.n0 VP.t3 578.672
R827 VP.n0 VP.t1 578.646
R828 VP.n2 VP.t0 557.689
R829 VP.n3 VP.t2 557.689
R830 VP.n4 VP.n3 161.3
R831 VP.n2 VP.n1 161.3
R832 VP.n1 VP.n0 111.48
R833 VP.n3 VP.n2 48.2005
R834 VP.n4 VP.n1 0.189894
R835 VP VP.n4 0.0516364
R836 VDD1 VDD1.n1 110.358
R837 VDD1 VDD1.n0 72.3048
R838 VDD1.n0 VDD1.t3 2.46674
R839 VDD1.n0 VDD1.t1 2.46674
R840 VDD1.n1 VDD1.t0 2.46674
R841 VDD1.n1 VDD1.t2 2.46674
R842 VTAIL.n5 VTAIL.t4 58.0343
R843 VTAIL.n4 VTAIL.t1 58.0343
R844 VTAIL.n3 VTAIL.t3 58.0343
R845 VTAIL.n7 VTAIL.t0 58.034
R846 VTAIL.n0 VTAIL.t2 58.034
R847 VTAIL.n1 VTAIL.t5 58.034
R848 VTAIL.n2 VTAIL.t7 58.034
R849 VTAIL.n6 VTAIL.t6 58.034
R850 VTAIL.n7 VTAIL.n6 24.5652
R851 VTAIL.n3 VTAIL.n2 24.5652
R852 VTAIL.n4 VTAIL.n3 0.836707
R853 VTAIL.n6 VTAIL.n5 0.836707
R854 VTAIL.n2 VTAIL.n1 0.836707
R855 VTAIL VTAIL.n0 0.476793
R856 VTAIL.n5 VTAIL.n4 0.470328
R857 VTAIL.n1 VTAIL.n0 0.470328
R858 VTAIL VTAIL.n7 0.360414
R859 VN.n0 VN.t2 578.672
R860 VN.n1 VN.t1 578.672
R861 VN.n0 VN.t0 578.646
R862 VN.n1 VN.t3 578.646
R863 VN VN.n1 111.859
R864 VN VN.n0 70.265
R865 VDD2.n2 VDD2.n0 109.832
R866 VDD2.n2 VDD2.n1 72.2466
R867 VDD2.n1 VDD2.t0 2.46674
R868 VDD2.n1 VDD2.t2 2.46674
R869 VDD2.n0 VDD2.t1 2.46674
R870 VDD2.n0 VDD2.t3 2.46674
R871 VDD2 VDD2.n2 0.0586897
C0 B w_n1552_n3604# 7.16464f
C1 VN VDD2 3.29877f
C2 VDD2 w_n1552_n3604# 1.09729f
C3 VDD2 B 0.967842f
C4 VDD1 VTAIL 7.5617f
C5 VDD1 VP 3.42089f
C6 VP VTAIL 2.85945f
C7 VN VDD1 0.147668f
C8 VDD1 w_n1552_n3604# 1.08396f
C9 VDD1 B 0.947157f
C10 VN VTAIL 2.84535f
C11 VN VP 4.99055f
C12 VTAIL w_n1552_n3604# 4.44091f
C13 VTAIL B 4.08278f
C14 VP w_n1552_n3604# 2.46819f
C15 VP B 1.0644f
C16 VDD1 VDD2 0.55485f
C17 VDD2 VTAIL 7.60277f
C18 VDD2 VP 0.270026f
C19 VN w_n1552_n3604# 2.27363f
C20 VN B 0.750658f
C21 VDD2 VSUBS 0.697576f
C22 VDD1 VSUBS 5.175566f
C23 VTAIL VSUBS 0.88655f
C24 VN VSUBS 6.13947f
C25 VP VSUBS 1.317439f
C26 B VSUBS 2.668329f
C27 w_n1552_n3604# VSUBS 68.7412f
C28 VDD2.t1 VSUBS 0.297729f
C29 VDD2.t3 VSUBS 0.297729f
C30 VDD2.n0 VSUBS 3.05559f
C31 VDD2.t0 VSUBS 0.297729f
C32 VDD2.t2 VSUBS 0.297729f
C33 VDD2.n1 VSUBS 2.35695f
C34 VDD2.n2 VSUBS 4.21336f
C35 VN.t2 VSUBS 1.48952f
C36 VN.t0 VSUBS 1.48949f
C37 VN.n0 VSUBS 1.11703f
C38 VN.t1 VSUBS 1.48952f
C39 VN.t3 VSUBS 1.48949f
C40 VN.n1 VSUBS 2.07546f
C41 VTAIL.t2 VSUBS 2.34341f
C42 VTAIL.n0 VSUBS 0.709448f
C43 VTAIL.t5 VSUBS 2.34341f
C44 VTAIL.n1 VSUBS 0.736322f
C45 VTAIL.t7 VSUBS 2.34341f
C46 VTAIL.n2 VSUBS 1.92685f
C47 VTAIL.t3 VSUBS 2.34342f
C48 VTAIL.n3 VSUBS 1.92684f
C49 VTAIL.t1 VSUBS 2.34342f
C50 VTAIL.n4 VSUBS 0.736315f
C51 VTAIL.t4 VSUBS 2.34342f
C52 VTAIL.n5 VSUBS 0.736315f
C53 VTAIL.t6 VSUBS 2.34341f
C54 VTAIL.n6 VSUBS 1.92685f
C55 VTAIL.t0 VSUBS 2.34341f
C56 VTAIL.n7 VSUBS 1.89129f
C57 VDD1.t3 VSUBS 0.297578f
C58 VDD1.t1 VSUBS 0.297578f
C59 VDD1.n0 VSUBS 2.35628f
C60 VDD1.t0 VSUBS 0.297578f
C61 VDD1.t2 VSUBS 0.297578f
C62 VDD1.n1 VSUBS 3.0804f
C63 VP.t1 VSUBS 1.54386f
C64 VP.t3 VSUBS 1.54388f
C65 VP.n0 VSUBS 2.13007f
C66 VP.n1 VSUBS 4.24963f
C67 VP.t0 VSUBS 1.52211f
C68 VP.n2 VSUBS 0.600565f
C69 VP.t2 VSUBS 1.52211f
C70 VP.n3 VSUBS 0.600565f
C71 VP.n4 VSUBS 0.049116f
C72 B.n0 VSUBS 0.007229f
C73 B.n1 VSUBS 0.007229f
C74 B.n2 VSUBS 0.010691f
C75 B.n3 VSUBS 0.008193f
C76 B.n4 VSUBS 0.008193f
C77 B.n5 VSUBS 0.008193f
C78 B.n6 VSUBS 0.008193f
C79 B.n7 VSUBS 0.008193f
C80 B.n8 VSUBS 0.008193f
C81 B.n9 VSUBS 0.008193f
C82 B.n10 VSUBS 0.019968f
C83 B.n11 VSUBS 0.008193f
C84 B.n12 VSUBS 0.008193f
C85 B.n13 VSUBS 0.008193f
C86 B.n14 VSUBS 0.008193f
C87 B.n15 VSUBS 0.008193f
C88 B.n16 VSUBS 0.008193f
C89 B.n17 VSUBS 0.008193f
C90 B.n18 VSUBS 0.008193f
C91 B.n19 VSUBS 0.008193f
C92 B.n20 VSUBS 0.008193f
C93 B.n21 VSUBS 0.008193f
C94 B.n22 VSUBS 0.008193f
C95 B.n23 VSUBS 0.008193f
C96 B.n24 VSUBS 0.008193f
C97 B.n25 VSUBS 0.008193f
C98 B.n26 VSUBS 0.008193f
C99 B.n27 VSUBS 0.008193f
C100 B.n28 VSUBS 0.008193f
C101 B.n29 VSUBS 0.008193f
C102 B.n30 VSUBS 0.008193f
C103 B.n31 VSUBS 0.008193f
C104 B.n32 VSUBS 0.007711f
C105 B.n33 VSUBS 0.008193f
C106 B.t4 VSUBS 0.507567f
C107 B.t5 VSUBS 0.516624f
C108 B.t3 VSUBS 0.402551f
C109 B.n34 VSUBS 0.162886f
C110 B.n35 VSUBS 0.074609f
C111 B.n36 VSUBS 0.018982f
C112 B.n37 VSUBS 0.008193f
C113 B.n38 VSUBS 0.008193f
C114 B.n39 VSUBS 0.008193f
C115 B.n40 VSUBS 0.008193f
C116 B.t1 VSUBS 0.507556f
C117 B.t2 VSUBS 0.516613f
C118 B.t0 VSUBS 0.402551f
C119 B.n41 VSUBS 0.162896f
C120 B.n42 VSUBS 0.07462f
C121 B.n43 VSUBS 0.008193f
C122 B.n44 VSUBS 0.008193f
C123 B.n45 VSUBS 0.008193f
C124 B.n46 VSUBS 0.008193f
C125 B.n47 VSUBS 0.008193f
C126 B.n48 VSUBS 0.008193f
C127 B.n49 VSUBS 0.008193f
C128 B.n50 VSUBS 0.008193f
C129 B.n51 VSUBS 0.008193f
C130 B.n52 VSUBS 0.008193f
C131 B.n53 VSUBS 0.008193f
C132 B.n54 VSUBS 0.008193f
C133 B.n55 VSUBS 0.008193f
C134 B.n56 VSUBS 0.008193f
C135 B.n57 VSUBS 0.008193f
C136 B.n58 VSUBS 0.008193f
C137 B.n59 VSUBS 0.008193f
C138 B.n60 VSUBS 0.008193f
C139 B.n61 VSUBS 0.008193f
C140 B.n62 VSUBS 0.008193f
C141 B.n63 VSUBS 0.008193f
C142 B.n64 VSUBS 0.008193f
C143 B.n65 VSUBS 0.018587f
C144 B.n66 VSUBS 0.008193f
C145 B.n67 VSUBS 0.008193f
C146 B.n68 VSUBS 0.008193f
C147 B.n69 VSUBS 0.008193f
C148 B.n70 VSUBS 0.008193f
C149 B.n71 VSUBS 0.008193f
C150 B.n72 VSUBS 0.008193f
C151 B.n73 VSUBS 0.008193f
C152 B.n74 VSUBS 0.008193f
C153 B.n75 VSUBS 0.008193f
C154 B.n76 VSUBS 0.008193f
C155 B.n77 VSUBS 0.008193f
C156 B.n78 VSUBS 0.008193f
C157 B.n79 VSUBS 0.008193f
C158 B.n80 VSUBS 0.008193f
C159 B.n81 VSUBS 0.008193f
C160 B.n82 VSUBS 0.019968f
C161 B.n83 VSUBS 0.008193f
C162 B.n84 VSUBS 0.008193f
C163 B.n85 VSUBS 0.008193f
C164 B.n86 VSUBS 0.008193f
C165 B.n87 VSUBS 0.008193f
C166 B.n88 VSUBS 0.008193f
C167 B.n89 VSUBS 0.008193f
C168 B.n90 VSUBS 0.008193f
C169 B.n91 VSUBS 0.008193f
C170 B.n92 VSUBS 0.008193f
C171 B.n93 VSUBS 0.008193f
C172 B.n94 VSUBS 0.008193f
C173 B.n95 VSUBS 0.008193f
C174 B.n96 VSUBS 0.008193f
C175 B.n97 VSUBS 0.008193f
C176 B.n98 VSUBS 0.008193f
C177 B.n99 VSUBS 0.008193f
C178 B.n100 VSUBS 0.008193f
C179 B.n101 VSUBS 0.008193f
C180 B.n102 VSUBS 0.008193f
C181 B.n103 VSUBS 0.008193f
C182 B.n104 VSUBS 0.008193f
C183 B.t11 VSUBS 0.507556f
C184 B.t10 VSUBS 0.516613f
C185 B.t9 VSUBS 0.402551f
C186 B.n105 VSUBS 0.162896f
C187 B.n106 VSUBS 0.07462f
C188 B.n107 VSUBS 0.008193f
C189 B.n108 VSUBS 0.008193f
C190 B.n109 VSUBS 0.008193f
C191 B.n110 VSUBS 0.008193f
C192 B.n111 VSUBS 0.004578f
C193 B.n112 VSUBS 0.008193f
C194 B.n113 VSUBS 0.008193f
C195 B.n114 VSUBS 0.008193f
C196 B.n115 VSUBS 0.008193f
C197 B.n116 VSUBS 0.008193f
C198 B.n117 VSUBS 0.008193f
C199 B.n118 VSUBS 0.008193f
C200 B.n119 VSUBS 0.008193f
C201 B.n120 VSUBS 0.008193f
C202 B.n121 VSUBS 0.008193f
C203 B.n122 VSUBS 0.008193f
C204 B.n123 VSUBS 0.008193f
C205 B.n124 VSUBS 0.008193f
C206 B.n125 VSUBS 0.008193f
C207 B.n126 VSUBS 0.008193f
C208 B.n127 VSUBS 0.008193f
C209 B.n128 VSUBS 0.008193f
C210 B.n129 VSUBS 0.008193f
C211 B.n130 VSUBS 0.008193f
C212 B.n131 VSUBS 0.008193f
C213 B.n132 VSUBS 0.008193f
C214 B.n133 VSUBS 0.008193f
C215 B.n134 VSUBS 0.018587f
C216 B.n135 VSUBS 0.008193f
C217 B.n136 VSUBS 0.008193f
C218 B.n137 VSUBS 0.008193f
C219 B.n138 VSUBS 0.008193f
C220 B.n139 VSUBS 0.008193f
C221 B.n140 VSUBS 0.008193f
C222 B.n141 VSUBS 0.008193f
C223 B.n142 VSUBS 0.008193f
C224 B.n143 VSUBS 0.008193f
C225 B.n144 VSUBS 0.008193f
C226 B.n145 VSUBS 0.008193f
C227 B.n146 VSUBS 0.008193f
C228 B.n147 VSUBS 0.008193f
C229 B.n148 VSUBS 0.008193f
C230 B.n149 VSUBS 0.008193f
C231 B.n150 VSUBS 0.008193f
C232 B.n151 VSUBS 0.008193f
C233 B.n152 VSUBS 0.008193f
C234 B.n153 VSUBS 0.008193f
C235 B.n154 VSUBS 0.008193f
C236 B.n155 VSUBS 0.008193f
C237 B.n156 VSUBS 0.008193f
C238 B.n157 VSUBS 0.008193f
C239 B.n158 VSUBS 0.008193f
C240 B.n159 VSUBS 0.008193f
C241 B.n160 VSUBS 0.008193f
C242 B.n161 VSUBS 0.008193f
C243 B.n162 VSUBS 0.008193f
C244 B.n163 VSUBS 0.018587f
C245 B.n164 VSUBS 0.019968f
C246 B.n165 VSUBS 0.019968f
C247 B.n166 VSUBS 0.008193f
C248 B.n167 VSUBS 0.008193f
C249 B.n168 VSUBS 0.008193f
C250 B.n169 VSUBS 0.008193f
C251 B.n170 VSUBS 0.008193f
C252 B.n171 VSUBS 0.008193f
C253 B.n172 VSUBS 0.008193f
C254 B.n173 VSUBS 0.008193f
C255 B.n174 VSUBS 0.008193f
C256 B.n175 VSUBS 0.008193f
C257 B.n176 VSUBS 0.008193f
C258 B.n177 VSUBS 0.008193f
C259 B.n178 VSUBS 0.008193f
C260 B.n179 VSUBS 0.008193f
C261 B.n180 VSUBS 0.008193f
C262 B.n181 VSUBS 0.008193f
C263 B.n182 VSUBS 0.008193f
C264 B.n183 VSUBS 0.008193f
C265 B.n184 VSUBS 0.008193f
C266 B.n185 VSUBS 0.008193f
C267 B.n186 VSUBS 0.008193f
C268 B.n187 VSUBS 0.008193f
C269 B.n188 VSUBS 0.008193f
C270 B.n189 VSUBS 0.008193f
C271 B.n190 VSUBS 0.008193f
C272 B.n191 VSUBS 0.008193f
C273 B.n192 VSUBS 0.008193f
C274 B.n193 VSUBS 0.008193f
C275 B.n194 VSUBS 0.008193f
C276 B.n195 VSUBS 0.008193f
C277 B.n196 VSUBS 0.008193f
C278 B.n197 VSUBS 0.008193f
C279 B.n198 VSUBS 0.008193f
C280 B.n199 VSUBS 0.008193f
C281 B.n200 VSUBS 0.008193f
C282 B.n201 VSUBS 0.008193f
C283 B.n202 VSUBS 0.008193f
C284 B.n203 VSUBS 0.008193f
C285 B.n204 VSUBS 0.008193f
C286 B.n205 VSUBS 0.008193f
C287 B.n206 VSUBS 0.008193f
C288 B.n207 VSUBS 0.008193f
C289 B.n208 VSUBS 0.008193f
C290 B.n209 VSUBS 0.008193f
C291 B.n210 VSUBS 0.008193f
C292 B.n211 VSUBS 0.008193f
C293 B.n212 VSUBS 0.008193f
C294 B.n213 VSUBS 0.008193f
C295 B.n214 VSUBS 0.008193f
C296 B.n215 VSUBS 0.008193f
C297 B.n216 VSUBS 0.008193f
C298 B.n217 VSUBS 0.008193f
C299 B.n218 VSUBS 0.008193f
C300 B.n219 VSUBS 0.008193f
C301 B.n220 VSUBS 0.008193f
C302 B.n221 VSUBS 0.008193f
C303 B.n222 VSUBS 0.008193f
C304 B.n223 VSUBS 0.008193f
C305 B.n224 VSUBS 0.008193f
C306 B.n225 VSUBS 0.008193f
C307 B.n226 VSUBS 0.008193f
C308 B.n227 VSUBS 0.008193f
C309 B.n228 VSUBS 0.008193f
C310 B.n229 VSUBS 0.008193f
C311 B.t8 VSUBS 0.507567f
C312 B.t7 VSUBS 0.516624f
C313 B.t6 VSUBS 0.402551f
C314 B.n230 VSUBS 0.162886f
C315 B.n231 VSUBS 0.074609f
C316 B.n232 VSUBS 0.018982f
C317 B.n233 VSUBS 0.007711f
C318 B.n234 VSUBS 0.008193f
C319 B.n235 VSUBS 0.008193f
C320 B.n236 VSUBS 0.008193f
C321 B.n237 VSUBS 0.008193f
C322 B.n238 VSUBS 0.008193f
C323 B.n239 VSUBS 0.008193f
C324 B.n240 VSUBS 0.008193f
C325 B.n241 VSUBS 0.008193f
C326 B.n242 VSUBS 0.008193f
C327 B.n243 VSUBS 0.008193f
C328 B.n244 VSUBS 0.008193f
C329 B.n245 VSUBS 0.008193f
C330 B.n246 VSUBS 0.008193f
C331 B.n247 VSUBS 0.008193f
C332 B.n248 VSUBS 0.008193f
C333 B.n249 VSUBS 0.004578f
C334 B.n250 VSUBS 0.018982f
C335 B.n251 VSUBS 0.007711f
C336 B.n252 VSUBS 0.008193f
C337 B.n253 VSUBS 0.008193f
C338 B.n254 VSUBS 0.008193f
C339 B.n255 VSUBS 0.008193f
C340 B.n256 VSUBS 0.008193f
C341 B.n257 VSUBS 0.008193f
C342 B.n258 VSUBS 0.008193f
C343 B.n259 VSUBS 0.008193f
C344 B.n260 VSUBS 0.008193f
C345 B.n261 VSUBS 0.008193f
C346 B.n262 VSUBS 0.008193f
C347 B.n263 VSUBS 0.008193f
C348 B.n264 VSUBS 0.008193f
C349 B.n265 VSUBS 0.008193f
C350 B.n266 VSUBS 0.008193f
C351 B.n267 VSUBS 0.008193f
C352 B.n268 VSUBS 0.008193f
C353 B.n269 VSUBS 0.008193f
C354 B.n270 VSUBS 0.008193f
C355 B.n271 VSUBS 0.008193f
C356 B.n272 VSUBS 0.008193f
C357 B.n273 VSUBS 0.008193f
C358 B.n274 VSUBS 0.008193f
C359 B.n275 VSUBS 0.008193f
C360 B.n276 VSUBS 0.008193f
C361 B.n277 VSUBS 0.008193f
C362 B.n278 VSUBS 0.008193f
C363 B.n279 VSUBS 0.008193f
C364 B.n280 VSUBS 0.008193f
C365 B.n281 VSUBS 0.008193f
C366 B.n282 VSUBS 0.008193f
C367 B.n283 VSUBS 0.008193f
C368 B.n284 VSUBS 0.008193f
C369 B.n285 VSUBS 0.008193f
C370 B.n286 VSUBS 0.008193f
C371 B.n287 VSUBS 0.008193f
C372 B.n288 VSUBS 0.008193f
C373 B.n289 VSUBS 0.008193f
C374 B.n290 VSUBS 0.008193f
C375 B.n291 VSUBS 0.008193f
C376 B.n292 VSUBS 0.008193f
C377 B.n293 VSUBS 0.008193f
C378 B.n294 VSUBS 0.008193f
C379 B.n295 VSUBS 0.008193f
C380 B.n296 VSUBS 0.008193f
C381 B.n297 VSUBS 0.008193f
C382 B.n298 VSUBS 0.008193f
C383 B.n299 VSUBS 0.008193f
C384 B.n300 VSUBS 0.008193f
C385 B.n301 VSUBS 0.008193f
C386 B.n302 VSUBS 0.008193f
C387 B.n303 VSUBS 0.008193f
C388 B.n304 VSUBS 0.008193f
C389 B.n305 VSUBS 0.008193f
C390 B.n306 VSUBS 0.008193f
C391 B.n307 VSUBS 0.008193f
C392 B.n308 VSUBS 0.008193f
C393 B.n309 VSUBS 0.008193f
C394 B.n310 VSUBS 0.008193f
C395 B.n311 VSUBS 0.008193f
C396 B.n312 VSUBS 0.008193f
C397 B.n313 VSUBS 0.008193f
C398 B.n314 VSUBS 0.008193f
C399 B.n315 VSUBS 0.008193f
C400 B.n316 VSUBS 0.008193f
C401 B.n317 VSUBS 0.019009f
C402 B.n318 VSUBS 0.019547f
C403 B.n319 VSUBS 0.018587f
C404 B.n320 VSUBS 0.008193f
C405 B.n321 VSUBS 0.008193f
C406 B.n322 VSUBS 0.008193f
C407 B.n323 VSUBS 0.008193f
C408 B.n324 VSUBS 0.008193f
C409 B.n325 VSUBS 0.008193f
C410 B.n326 VSUBS 0.008193f
C411 B.n327 VSUBS 0.008193f
C412 B.n328 VSUBS 0.008193f
C413 B.n329 VSUBS 0.008193f
C414 B.n330 VSUBS 0.008193f
C415 B.n331 VSUBS 0.008193f
C416 B.n332 VSUBS 0.008193f
C417 B.n333 VSUBS 0.008193f
C418 B.n334 VSUBS 0.008193f
C419 B.n335 VSUBS 0.008193f
C420 B.n336 VSUBS 0.008193f
C421 B.n337 VSUBS 0.008193f
C422 B.n338 VSUBS 0.008193f
C423 B.n339 VSUBS 0.008193f
C424 B.n340 VSUBS 0.008193f
C425 B.n341 VSUBS 0.008193f
C426 B.n342 VSUBS 0.008193f
C427 B.n343 VSUBS 0.008193f
C428 B.n344 VSUBS 0.008193f
C429 B.n345 VSUBS 0.008193f
C430 B.n346 VSUBS 0.008193f
C431 B.n347 VSUBS 0.008193f
C432 B.n348 VSUBS 0.008193f
C433 B.n349 VSUBS 0.008193f
C434 B.n350 VSUBS 0.008193f
C435 B.n351 VSUBS 0.008193f
C436 B.n352 VSUBS 0.008193f
C437 B.n353 VSUBS 0.008193f
C438 B.n354 VSUBS 0.008193f
C439 B.n355 VSUBS 0.008193f
C440 B.n356 VSUBS 0.008193f
C441 B.n357 VSUBS 0.008193f
C442 B.n358 VSUBS 0.008193f
C443 B.n359 VSUBS 0.008193f
C444 B.n360 VSUBS 0.008193f
C445 B.n361 VSUBS 0.008193f
C446 B.n362 VSUBS 0.008193f
C447 B.n363 VSUBS 0.008193f
C448 B.n364 VSUBS 0.008193f
C449 B.n365 VSUBS 0.008193f
C450 B.n366 VSUBS 0.008193f
C451 B.n367 VSUBS 0.008193f
C452 B.n368 VSUBS 0.018587f
C453 B.n369 VSUBS 0.019968f
C454 B.n370 VSUBS 0.019968f
C455 B.n371 VSUBS 0.008193f
C456 B.n372 VSUBS 0.008193f
C457 B.n373 VSUBS 0.008193f
C458 B.n374 VSUBS 0.008193f
C459 B.n375 VSUBS 0.008193f
C460 B.n376 VSUBS 0.008193f
C461 B.n377 VSUBS 0.008193f
C462 B.n378 VSUBS 0.008193f
C463 B.n379 VSUBS 0.008193f
C464 B.n380 VSUBS 0.008193f
C465 B.n381 VSUBS 0.008193f
C466 B.n382 VSUBS 0.008193f
C467 B.n383 VSUBS 0.008193f
C468 B.n384 VSUBS 0.008193f
C469 B.n385 VSUBS 0.008193f
C470 B.n386 VSUBS 0.008193f
C471 B.n387 VSUBS 0.008193f
C472 B.n388 VSUBS 0.008193f
C473 B.n389 VSUBS 0.008193f
C474 B.n390 VSUBS 0.008193f
C475 B.n391 VSUBS 0.008193f
C476 B.n392 VSUBS 0.008193f
C477 B.n393 VSUBS 0.008193f
C478 B.n394 VSUBS 0.008193f
C479 B.n395 VSUBS 0.008193f
C480 B.n396 VSUBS 0.008193f
C481 B.n397 VSUBS 0.008193f
C482 B.n398 VSUBS 0.008193f
C483 B.n399 VSUBS 0.008193f
C484 B.n400 VSUBS 0.008193f
C485 B.n401 VSUBS 0.008193f
C486 B.n402 VSUBS 0.008193f
C487 B.n403 VSUBS 0.008193f
C488 B.n404 VSUBS 0.008193f
C489 B.n405 VSUBS 0.008193f
C490 B.n406 VSUBS 0.008193f
C491 B.n407 VSUBS 0.008193f
C492 B.n408 VSUBS 0.008193f
C493 B.n409 VSUBS 0.008193f
C494 B.n410 VSUBS 0.008193f
C495 B.n411 VSUBS 0.008193f
C496 B.n412 VSUBS 0.008193f
C497 B.n413 VSUBS 0.008193f
C498 B.n414 VSUBS 0.008193f
C499 B.n415 VSUBS 0.008193f
C500 B.n416 VSUBS 0.008193f
C501 B.n417 VSUBS 0.008193f
C502 B.n418 VSUBS 0.008193f
C503 B.n419 VSUBS 0.008193f
C504 B.n420 VSUBS 0.008193f
C505 B.n421 VSUBS 0.008193f
C506 B.n422 VSUBS 0.008193f
C507 B.n423 VSUBS 0.008193f
C508 B.n424 VSUBS 0.008193f
C509 B.n425 VSUBS 0.008193f
C510 B.n426 VSUBS 0.008193f
C511 B.n427 VSUBS 0.008193f
C512 B.n428 VSUBS 0.008193f
C513 B.n429 VSUBS 0.008193f
C514 B.n430 VSUBS 0.008193f
C515 B.n431 VSUBS 0.008193f
C516 B.n432 VSUBS 0.008193f
C517 B.n433 VSUBS 0.008193f
C518 B.n434 VSUBS 0.008193f
C519 B.n435 VSUBS 0.008193f
C520 B.n436 VSUBS 0.007711f
C521 B.n437 VSUBS 0.018982f
C522 B.n438 VSUBS 0.004578f
C523 B.n439 VSUBS 0.008193f
C524 B.n440 VSUBS 0.008193f
C525 B.n441 VSUBS 0.008193f
C526 B.n442 VSUBS 0.008193f
C527 B.n443 VSUBS 0.008193f
C528 B.n444 VSUBS 0.008193f
C529 B.n445 VSUBS 0.008193f
C530 B.n446 VSUBS 0.008193f
C531 B.n447 VSUBS 0.008193f
C532 B.n448 VSUBS 0.008193f
C533 B.n449 VSUBS 0.008193f
C534 B.n450 VSUBS 0.008193f
C535 B.n451 VSUBS 0.004578f
C536 B.n452 VSUBS 0.008193f
C537 B.n453 VSUBS 0.008193f
C538 B.n454 VSUBS 0.008193f
C539 B.n455 VSUBS 0.008193f
C540 B.n456 VSUBS 0.008193f
C541 B.n457 VSUBS 0.008193f
C542 B.n458 VSUBS 0.008193f
C543 B.n459 VSUBS 0.008193f
C544 B.n460 VSUBS 0.008193f
C545 B.n461 VSUBS 0.008193f
C546 B.n462 VSUBS 0.008193f
C547 B.n463 VSUBS 0.008193f
C548 B.n464 VSUBS 0.008193f
C549 B.n465 VSUBS 0.008193f
C550 B.n466 VSUBS 0.008193f
C551 B.n467 VSUBS 0.008193f
C552 B.n468 VSUBS 0.008193f
C553 B.n469 VSUBS 0.008193f
C554 B.n470 VSUBS 0.008193f
C555 B.n471 VSUBS 0.008193f
C556 B.n472 VSUBS 0.008193f
C557 B.n473 VSUBS 0.008193f
C558 B.n474 VSUBS 0.008193f
C559 B.n475 VSUBS 0.008193f
C560 B.n476 VSUBS 0.008193f
C561 B.n477 VSUBS 0.008193f
C562 B.n478 VSUBS 0.008193f
C563 B.n479 VSUBS 0.008193f
C564 B.n480 VSUBS 0.008193f
C565 B.n481 VSUBS 0.008193f
C566 B.n482 VSUBS 0.008193f
C567 B.n483 VSUBS 0.008193f
C568 B.n484 VSUBS 0.008193f
C569 B.n485 VSUBS 0.008193f
C570 B.n486 VSUBS 0.008193f
C571 B.n487 VSUBS 0.008193f
C572 B.n488 VSUBS 0.008193f
C573 B.n489 VSUBS 0.008193f
C574 B.n490 VSUBS 0.008193f
C575 B.n491 VSUBS 0.008193f
C576 B.n492 VSUBS 0.008193f
C577 B.n493 VSUBS 0.008193f
C578 B.n494 VSUBS 0.008193f
C579 B.n495 VSUBS 0.008193f
C580 B.n496 VSUBS 0.008193f
C581 B.n497 VSUBS 0.008193f
C582 B.n498 VSUBS 0.008193f
C583 B.n499 VSUBS 0.008193f
C584 B.n500 VSUBS 0.008193f
C585 B.n501 VSUBS 0.008193f
C586 B.n502 VSUBS 0.008193f
C587 B.n503 VSUBS 0.008193f
C588 B.n504 VSUBS 0.008193f
C589 B.n505 VSUBS 0.008193f
C590 B.n506 VSUBS 0.008193f
C591 B.n507 VSUBS 0.008193f
C592 B.n508 VSUBS 0.008193f
C593 B.n509 VSUBS 0.008193f
C594 B.n510 VSUBS 0.008193f
C595 B.n511 VSUBS 0.008193f
C596 B.n512 VSUBS 0.008193f
C597 B.n513 VSUBS 0.008193f
C598 B.n514 VSUBS 0.008193f
C599 B.n515 VSUBS 0.008193f
C600 B.n516 VSUBS 0.008193f
C601 B.n517 VSUBS 0.008193f
C602 B.n518 VSUBS 0.008193f
C603 B.n519 VSUBS 0.019968f
C604 B.n520 VSUBS 0.018587f
C605 B.n521 VSUBS 0.018587f
C606 B.n522 VSUBS 0.008193f
C607 B.n523 VSUBS 0.008193f
C608 B.n524 VSUBS 0.008193f
C609 B.n525 VSUBS 0.008193f
C610 B.n526 VSUBS 0.008193f
C611 B.n527 VSUBS 0.008193f
C612 B.n528 VSUBS 0.008193f
C613 B.n529 VSUBS 0.008193f
C614 B.n530 VSUBS 0.008193f
C615 B.n531 VSUBS 0.008193f
C616 B.n532 VSUBS 0.008193f
C617 B.n533 VSUBS 0.008193f
C618 B.n534 VSUBS 0.008193f
C619 B.n535 VSUBS 0.008193f
C620 B.n536 VSUBS 0.008193f
C621 B.n537 VSUBS 0.008193f
C622 B.n538 VSUBS 0.008193f
C623 B.n539 VSUBS 0.008193f
C624 B.n540 VSUBS 0.008193f
C625 B.n541 VSUBS 0.008193f
C626 B.n542 VSUBS 0.008193f
C627 B.n543 VSUBS 0.010691f
C628 B.n544 VSUBS 0.011389f
C629 B.n545 VSUBS 0.022648f
.ends

