* NGSPICE file created from diff_pair_sample_0863.ext - technology: sky130A

.subckt diff_pair_sample_0863 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=0 ps=0 w=10.57 l=0.7
X1 VTAIL.t15 VP.t0 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X2 VTAIL.t7 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X3 VDD2.t6 VN.t1 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X4 VTAIL.t5 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=1.74405 ps=10.9 w=10.57 l=0.7
X5 VTAIL.t14 VP.t1 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=1.74405 ps=10.9 w=10.57 l=0.7
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=0 ps=0 w=10.57 l=0.7
X7 VTAIL.t13 VP.t2 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=1.74405 ps=10.9 w=10.57 l=0.7
X8 VDD2.t4 VN.t3 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X9 VDD1.t7 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=4.1223 ps=21.92 w=10.57 l=0.7
X10 VDD2.t3 VN.t4 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=4.1223 ps=21.92 w=10.57 l=0.7
X11 VDD1.t5 VP.t4 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X12 VDD1.t4 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=0 ps=0 w=10.57 l=0.7
X14 VDD1.t3 VP.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=4.1223 ps=21.92 w=10.57 l=0.7
X15 VTAIL.t1 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X16 VTAIL.t8 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=1.74405 ps=10.9 w=10.57 l=0.7
X17 VTAIL.t2 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=1.74405 ps=10.9 w=10.57 l=0.7
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1223 pd=21.92 as=0 ps=0 w=10.57 l=0.7
X19 VDD2.t0 VN.t7 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.74405 pd=10.9 as=4.1223 ps=21.92 w=10.57 l=0.7
R0 B.n614 B.n613 585
R1 B.n255 B.n87 585
R2 B.n254 B.n253 585
R3 B.n252 B.n251 585
R4 B.n250 B.n249 585
R5 B.n248 B.n247 585
R6 B.n246 B.n245 585
R7 B.n244 B.n243 585
R8 B.n242 B.n241 585
R9 B.n240 B.n239 585
R10 B.n238 B.n237 585
R11 B.n236 B.n235 585
R12 B.n234 B.n233 585
R13 B.n232 B.n231 585
R14 B.n230 B.n229 585
R15 B.n228 B.n227 585
R16 B.n226 B.n225 585
R17 B.n224 B.n223 585
R18 B.n222 B.n221 585
R19 B.n220 B.n219 585
R20 B.n218 B.n217 585
R21 B.n216 B.n215 585
R22 B.n214 B.n213 585
R23 B.n212 B.n211 585
R24 B.n210 B.n209 585
R25 B.n208 B.n207 585
R26 B.n206 B.n205 585
R27 B.n204 B.n203 585
R28 B.n202 B.n201 585
R29 B.n200 B.n199 585
R30 B.n198 B.n197 585
R31 B.n196 B.n195 585
R32 B.n194 B.n193 585
R33 B.n192 B.n191 585
R34 B.n190 B.n189 585
R35 B.n188 B.n187 585
R36 B.n186 B.n185 585
R37 B.n183 B.n182 585
R38 B.n181 B.n180 585
R39 B.n179 B.n178 585
R40 B.n177 B.n176 585
R41 B.n175 B.n174 585
R42 B.n173 B.n172 585
R43 B.n171 B.n170 585
R44 B.n169 B.n168 585
R45 B.n167 B.n166 585
R46 B.n165 B.n164 585
R47 B.n162 B.n161 585
R48 B.n160 B.n159 585
R49 B.n158 B.n157 585
R50 B.n156 B.n155 585
R51 B.n154 B.n153 585
R52 B.n152 B.n151 585
R53 B.n150 B.n149 585
R54 B.n148 B.n147 585
R55 B.n146 B.n145 585
R56 B.n144 B.n143 585
R57 B.n142 B.n141 585
R58 B.n140 B.n139 585
R59 B.n138 B.n137 585
R60 B.n136 B.n135 585
R61 B.n134 B.n133 585
R62 B.n132 B.n131 585
R63 B.n130 B.n129 585
R64 B.n128 B.n127 585
R65 B.n126 B.n125 585
R66 B.n124 B.n123 585
R67 B.n122 B.n121 585
R68 B.n120 B.n119 585
R69 B.n118 B.n117 585
R70 B.n116 B.n115 585
R71 B.n114 B.n113 585
R72 B.n112 B.n111 585
R73 B.n110 B.n109 585
R74 B.n108 B.n107 585
R75 B.n106 B.n105 585
R76 B.n104 B.n103 585
R77 B.n102 B.n101 585
R78 B.n100 B.n99 585
R79 B.n98 B.n97 585
R80 B.n96 B.n95 585
R81 B.n94 B.n93 585
R82 B.n46 B.n45 585
R83 B.n619 B.n618 585
R84 B.n612 B.n88 585
R85 B.n88 B.n43 585
R86 B.n611 B.n42 585
R87 B.n623 B.n42 585
R88 B.n610 B.n41 585
R89 B.n624 B.n41 585
R90 B.n609 B.n40 585
R91 B.n625 B.n40 585
R92 B.n608 B.n607 585
R93 B.n607 B.n39 585
R94 B.n606 B.n35 585
R95 B.n631 B.n35 585
R96 B.n605 B.n34 585
R97 B.n632 B.n34 585
R98 B.n604 B.n33 585
R99 B.n633 B.n33 585
R100 B.n603 B.n602 585
R101 B.n602 B.n29 585
R102 B.n601 B.n28 585
R103 B.n639 B.n28 585
R104 B.n600 B.n27 585
R105 B.n640 B.n27 585
R106 B.n599 B.n26 585
R107 B.n641 B.n26 585
R108 B.n598 B.n597 585
R109 B.n597 B.n22 585
R110 B.n596 B.n21 585
R111 B.n647 B.n21 585
R112 B.n595 B.n20 585
R113 B.n648 B.n20 585
R114 B.n594 B.n19 585
R115 B.n649 B.n19 585
R116 B.n593 B.n592 585
R117 B.n592 B.n18 585
R118 B.n591 B.n14 585
R119 B.n655 B.n14 585
R120 B.n590 B.n13 585
R121 B.n656 B.n13 585
R122 B.n589 B.n12 585
R123 B.n657 B.n12 585
R124 B.n588 B.n587 585
R125 B.n587 B.n8 585
R126 B.n586 B.n7 585
R127 B.n663 B.n7 585
R128 B.n585 B.n6 585
R129 B.n664 B.n6 585
R130 B.n584 B.n5 585
R131 B.n665 B.n5 585
R132 B.n583 B.n582 585
R133 B.n582 B.n4 585
R134 B.n581 B.n256 585
R135 B.n581 B.n580 585
R136 B.n571 B.n257 585
R137 B.n258 B.n257 585
R138 B.n573 B.n572 585
R139 B.n574 B.n573 585
R140 B.n570 B.n263 585
R141 B.n263 B.n262 585
R142 B.n569 B.n568 585
R143 B.n568 B.n567 585
R144 B.n265 B.n264 585
R145 B.n560 B.n265 585
R146 B.n559 B.n558 585
R147 B.n561 B.n559 585
R148 B.n557 B.n270 585
R149 B.n270 B.n269 585
R150 B.n556 B.n555 585
R151 B.n555 B.n554 585
R152 B.n272 B.n271 585
R153 B.n273 B.n272 585
R154 B.n547 B.n546 585
R155 B.n548 B.n547 585
R156 B.n545 B.n277 585
R157 B.n281 B.n277 585
R158 B.n544 B.n543 585
R159 B.n543 B.n542 585
R160 B.n279 B.n278 585
R161 B.n280 B.n279 585
R162 B.n535 B.n534 585
R163 B.n536 B.n535 585
R164 B.n533 B.n286 585
R165 B.n286 B.n285 585
R166 B.n532 B.n531 585
R167 B.n531 B.n530 585
R168 B.n288 B.n287 585
R169 B.n523 B.n288 585
R170 B.n522 B.n521 585
R171 B.n524 B.n522 585
R172 B.n520 B.n293 585
R173 B.n293 B.n292 585
R174 B.n519 B.n518 585
R175 B.n518 B.n517 585
R176 B.n295 B.n294 585
R177 B.n296 B.n295 585
R178 B.n513 B.n512 585
R179 B.n299 B.n298 585
R180 B.n509 B.n508 585
R181 B.n510 B.n509 585
R182 B.n507 B.n341 585
R183 B.n506 B.n505 585
R184 B.n504 B.n503 585
R185 B.n502 B.n501 585
R186 B.n500 B.n499 585
R187 B.n498 B.n497 585
R188 B.n496 B.n495 585
R189 B.n494 B.n493 585
R190 B.n492 B.n491 585
R191 B.n490 B.n489 585
R192 B.n488 B.n487 585
R193 B.n486 B.n485 585
R194 B.n484 B.n483 585
R195 B.n482 B.n481 585
R196 B.n480 B.n479 585
R197 B.n478 B.n477 585
R198 B.n476 B.n475 585
R199 B.n474 B.n473 585
R200 B.n472 B.n471 585
R201 B.n470 B.n469 585
R202 B.n468 B.n467 585
R203 B.n466 B.n465 585
R204 B.n464 B.n463 585
R205 B.n462 B.n461 585
R206 B.n460 B.n459 585
R207 B.n458 B.n457 585
R208 B.n456 B.n455 585
R209 B.n454 B.n453 585
R210 B.n452 B.n451 585
R211 B.n450 B.n449 585
R212 B.n448 B.n447 585
R213 B.n446 B.n445 585
R214 B.n444 B.n443 585
R215 B.n442 B.n441 585
R216 B.n440 B.n439 585
R217 B.n438 B.n437 585
R218 B.n436 B.n435 585
R219 B.n434 B.n433 585
R220 B.n432 B.n431 585
R221 B.n430 B.n429 585
R222 B.n428 B.n427 585
R223 B.n426 B.n425 585
R224 B.n424 B.n423 585
R225 B.n422 B.n421 585
R226 B.n420 B.n419 585
R227 B.n418 B.n417 585
R228 B.n416 B.n415 585
R229 B.n414 B.n413 585
R230 B.n412 B.n411 585
R231 B.n410 B.n409 585
R232 B.n408 B.n407 585
R233 B.n406 B.n405 585
R234 B.n404 B.n403 585
R235 B.n402 B.n401 585
R236 B.n400 B.n399 585
R237 B.n398 B.n397 585
R238 B.n396 B.n395 585
R239 B.n394 B.n393 585
R240 B.n392 B.n391 585
R241 B.n390 B.n389 585
R242 B.n388 B.n387 585
R243 B.n386 B.n385 585
R244 B.n384 B.n383 585
R245 B.n382 B.n381 585
R246 B.n380 B.n379 585
R247 B.n378 B.n377 585
R248 B.n376 B.n375 585
R249 B.n374 B.n373 585
R250 B.n372 B.n371 585
R251 B.n370 B.n369 585
R252 B.n368 B.n367 585
R253 B.n366 B.n365 585
R254 B.n364 B.n363 585
R255 B.n362 B.n361 585
R256 B.n360 B.n359 585
R257 B.n358 B.n357 585
R258 B.n356 B.n355 585
R259 B.n354 B.n353 585
R260 B.n352 B.n351 585
R261 B.n350 B.n349 585
R262 B.n348 B.n340 585
R263 B.n510 B.n340 585
R264 B.n514 B.n297 585
R265 B.n297 B.n296 585
R266 B.n516 B.n515 585
R267 B.n517 B.n516 585
R268 B.n291 B.n290 585
R269 B.n292 B.n291 585
R270 B.n526 B.n525 585
R271 B.n525 B.n524 585
R272 B.n527 B.n289 585
R273 B.n523 B.n289 585
R274 B.n529 B.n528 585
R275 B.n530 B.n529 585
R276 B.n284 B.n283 585
R277 B.n285 B.n284 585
R278 B.n538 B.n537 585
R279 B.n537 B.n536 585
R280 B.n539 B.n282 585
R281 B.n282 B.n280 585
R282 B.n541 B.n540 585
R283 B.n542 B.n541 585
R284 B.n276 B.n275 585
R285 B.n281 B.n276 585
R286 B.n550 B.n549 585
R287 B.n549 B.n548 585
R288 B.n551 B.n274 585
R289 B.n274 B.n273 585
R290 B.n553 B.n552 585
R291 B.n554 B.n553 585
R292 B.n268 B.n267 585
R293 B.n269 B.n268 585
R294 B.n563 B.n562 585
R295 B.n562 B.n561 585
R296 B.n564 B.n266 585
R297 B.n560 B.n266 585
R298 B.n566 B.n565 585
R299 B.n567 B.n566 585
R300 B.n261 B.n260 585
R301 B.n262 B.n261 585
R302 B.n576 B.n575 585
R303 B.n575 B.n574 585
R304 B.n577 B.n259 585
R305 B.n259 B.n258 585
R306 B.n579 B.n578 585
R307 B.n580 B.n579 585
R308 B.n2 B.n0 585
R309 B.n4 B.n2 585
R310 B.n3 B.n1 585
R311 B.n664 B.n3 585
R312 B.n662 B.n661 585
R313 B.n663 B.n662 585
R314 B.n660 B.n9 585
R315 B.n9 B.n8 585
R316 B.n659 B.n658 585
R317 B.n658 B.n657 585
R318 B.n11 B.n10 585
R319 B.n656 B.n11 585
R320 B.n654 B.n653 585
R321 B.n655 B.n654 585
R322 B.n652 B.n15 585
R323 B.n18 B.n15 585
R324 B.n651 B.n650 585
R325 B.n650 B.n649 585
R326 B.n17 B.n16 585
R327 B.n648 B.n17 585
R328 B.n646 B.n645 585
R329 B.n647 B.n646 585
R330 B.n644 B.n23 585
R331 B.n23 B.n22 585
R332 B.n643 B.n642 585
R333 B.n642 B.n641 585
R334 B.n25 B.n24 585
R335 B.n640 B.n25 585
R336 B.n638 B.n637 585
R337 B.n639 B.n638 585
R338 B.n636 B.n30 585
R339 B.n30 B.n29 585
R340 B.n635 B.n634 585
R341 B.n634 B.n633 585
R342 B.n32 B.n31 585
R343 B.n632 B.n32 585
R344 B.n630 B.n629 585
R345 B.n631 B.n630 585
R346 B.n628 B.n36 585
R347 B.n39 B.n36 585
R348 B.n627 B.n626 585
R349 B.n626 B.n625 585
R350 B.n38 B.n37 585
R351 B.n624 B.n38 585
R352 B.n622 B.n621 585
R353 B.n623 B.n622 585
R354 B.n620 B.n44 585
R355 B.n44 B.n43 585
R356 B.n667 B.n666 585
R357 B.n666 B.n665 585
R358 B.n512 B.n297 574.183
R359 B.n618 B.n44 574.183
R360 B.n340 B.n295 574.183
R361 B.n614 B.n88 574.183
R362 B.n345 B.t15 566.875
R363 B.n342 B.t19 566.875
R364 B.n91 B.t12 566.875
R365 B.n89 B.t8 566.875
R366 B.n345 B.t18 277.202
R367 B.n89 B.t10 277.202
R368 B.n342 B.t21 277.202
R369 B.n91 B.t13 277.202
R370 B.n346 B.t17 257.226
R371 B.n90 B.t11 257.226
R372 B.n343 B.t20 257.226
R373 B.n92 B.t14 257.226
R374 B.n616 B.n615 256.663
R375 B.n616 B.n86 256.663
R376 B.n616 B.n85 256.663
R377 B.n616 B.n84 256.663
R378 B.n616 B.n83 256.663
R379 B.n616 B.n82 256.663
R380 B.n616 B.n81 256.663
R381 B.n616 B.n80 256.663
R382 B.n616 B.n79 256.663
R383 B.n616 B.n78 256.663
R384 B.n616 B.n77 256.663
R385 B.n616 B.n76 256.663
R386 B.n616 B.n75 256.663
R387 B.n616 B.n74 256.663
R388 B.n616 B.n73 256.663
R389 B.n616 B.n72 256.663
R390 B.n616 B.n71 256.663
R391 B.n616 B.n70 256.663
R392 B.n616 B.n69 256.663
R393 B.n616 B.n68 256.663
R394 B.n616 B.n67 256.663
R395 B.n616 B.n66 256.663
R396 B.n616 B.n65 256.663
R397 B.n616 B.n64 256.663
R398 B.n616 B.n63 256.663
R399 B.n616 B.n62 256.663
R400 B.n616 B.n61 256.663
R401 B.n616 B.n60 256.663
R402 B.n616 B.n59 256.663
R403 B.n616 B.n58 256.663
R404 B.n616 B.n57 256.663
R405 B.n616 B.n56 256.663
R406 B.n616 B.n55 256.663
R407 B.n616 B.n54 256.663
R408 B.n616 B.n53 256.663
R409 B.n616 B.n52 256.663
R410 B.n616 B.n51 256.663
R411 B.n616 B.n50 256.663
R412 B.n616 B.n49 256.663
R413 B.n616 B.n48 256.663
R414 B.n616 B.n47 256.663
R415 B.n617 B.n616 256.663
R416 B.n511 B.n510 256.663
R417 B.n510 B.n300 256.663
R418 B.n510 B.n301 256.663
R419 B.n510 B.n302 256.663
R420 B.n510 B.n303 256.663
R421 B.n510 B.n304 256.663
R422 B.n510 B.n305 256.663
R423 B.n510 B.n306 256.663
R424 B.n510 B.n307 256.663
R425 B.n510 B.n308 256.663
R426 B.n510 B.n309 256.663
R427 B.n510 B.n310 256.663
R428 B.n510 B.n311 256.663
R429 B.n510 B.n312 256.663
R430 B.n510 B.n313 256.663
R431 B.n510 B.n314 256.663
R432 B.n510 B.n315 256.663
R433 B.n510 B.n316 256.663
R434 B.n510 B.n317 256.663
R435 B.n510 B.n318 256.663
R436 B.n510 B.n319 256.663
R437 B.n510 B.n320 256.663
R438 B.n510 B.n321 256.663
R439 B.n510 B.n322 256.663
R440 B.n510 B.n323 256.663
R441 B.n510 B.n324 256.663
R442 B.n510 B.n325 256.663
R443 B.n510 B.n326 256.663
R444 B.n510 B.n327 256.663
R445 B.n510 B.n328 256.663
R446 B.n510 B.n329 256.663
R447 B.n510 B.n330 256.663
R448 B.n510 B.n331 256.663
R449 B.n510 B.n332 256.663
R450 B.n510 B.n333 256.663
R451 B.n510 B.n334 256.663
R452 B.n510 B.n335 256.663
R453 B.n510 B.n336 256.663
R454 B.n510 B.n337 256.663
R455 B.n510 B.n338 256.663
R456 B.n510 B.n339 256.663
R457 B.n516 B.n297 163.367
R458 B.n516 B.n291 163.367
R459 B.n525 B.n291 163.367
R460 B.n525 B.n289 163.367
R461 B.n529 B.n289 163.367
R462 B.n529 B.n284 163.367
R463 B.n537 B.n284 163.367
R464 B.n537 B.n282 163.367
R465 B.n541 B.n282 163.367
R466 B.n541 B.n276 163.367
R467 B.n549 B.n276 163.367
R468 B.n549 B.n274 163.367
R469 B.n553 B.n274 163.367
R470 B.n553 B.n268 163.367
R471 B.n562 B.n268 163.367
R472 B.n562 B.n266 163.367
R473 B.n566 B.n266 163.367
R474 B.n566 B.n261 163.367
R475 B.n575 B.n261 163.367
R476 B.n575 B.n259 163.367
R477 B.n579 B.n259 163.367
R478 B.n579 B.n2 163.367
R479 B.n666 B.n2 163.367
R480 B.n666 B.n3 163.367
R481 B.n662 B.n3 163.367
R482 B.n662 B.n9 163.367
R483 B.n658 B.n9 163.367
R484 B.n658 B.n11 163.367
R485 B.n654 B.n11 163.367
R486 B.n654 B.n15 163.367
R487 B.n650 B.n15 163.367
R488 B.n650 B.n17 163.367
R489 B.n646 B.n17 163.367
R490 B.n646 B.n23 163.367
R491 B.n642 B.n23 163.367
R492 B.n642 B.n25 163.367
R493 B.n638 B.n25 163.367
R494 B.n638 B.n30 163.367
R495 B.n634 B.n30 163.367
R496 B.n634 B.n32 163.367
R497 B.n630 B.n32 163.367
R498 B.n630 B.n36 163.367
R499 B.n626 B.n36 163.367
R500 B.n626 B.n38 163.367
R501 B.n622 B.n38 163.367
R502 B.n622 B.n44 163.367
R503 B.n509 B.n299 163.367
R504 B.n509 B.n341 163.367
R505 B.n505 B.n504 163.367
R506 B.n501 B.n500 163.367
R507 B.n497 B.n496 163.367
R508 B.n493 B.n492 163.367
R509 B.n489 B.n488 163.367
R510 B.n485 B.n484 163.367
R511 B.n481 B.n480 163.367
R512 B.n477 B.n476 163.367
R513 B.n473 B.n472 163.367
R514 B.n469 B.n468 163.367
R515 B.n465 B.n464 163.367
R516 B.n461 B.n460 163.367
R517 B.n457 B.n456 163.367
R518 B.n453 B.n452 163.367
R519 B.n449 B.n448 163.367
R520 B.n445 B.n444 163.367
R521 B.n441 B.n440 163.367
R522 B.n437 B.n436 163.367
R523 B.n433 B.n432 163.367
R524 B.n429 B.n428 163.367
R525 B.n425 B.n424 163.367
R526 B.n421 B.n420 163.367
R527 B.n417 B.n416 163.367
R528 B.n413 B.n412 163.367
R529 B.n409 B.n408 163.367
R530 B.n405 B.n404 163.367
R531 B.n401 B.n400 163.367
R532 B.n397 B.n396 163.367
R533 B.n393 B.n392 163.367
R534 B.n389 B.n388 163.367
R535 B.n385 B.n384 163.367
R536 B.n381 B.n380 163.367
R537 B.n377 B.n376 163.367
R538 B.n373 B.n372 163.367
R539 B.n369 B.n368 163.367
R540 B.n365 B.n364 163.367
R541 B.n361 B.n360 163.367
R542 B.n357 B.n356 163.367
R543 B.n353 B.n352 163.367
R544 B.n349 B.n340 163.367
R545 B.n518 B.n295 163.367
R546 B.n518 B.n293 163.367
R547 B.n522 B.n293 163.367
R548 B.n522 B.n288 163.367
R549 B.n531 B.n288 163.367
R550 B.n531 B.n286 163.367
R551 B.n535 B.n286 163.367
R552 B.n535 B.n279 163.367
R553 B.n543 B.n279 163.367
R554 B.n543 B.n277 163.367
R555 B.n547 B.n277 163.367
R556 B.n547 B.n272 163.367
R557 B.n555 B.n272 163.367
R558 B.n555 B.n270 163.367
R559 B.n559 B.n270 163.367
R560 B.n559 B.n265 163.367
R561 B.n568 B.n265 163.367
R562 B.n568 B.n263 163.367
R563 B.n573 B.n263 163.367
R564 B.n573 B.n257 163.367
R565 B.n581 B.n257 163.367
R566 B.n582 B.n581 163.367
R567 B.n582 B.n5 163.367
R568 B.n6 B.n5 163.367
R569 B.n7 B.n6 163.367
R570 B.n587 B.n7 163.367
R571 B.n587 B.n12 163.367
R572 B.n13 B.n12 163.367
R573 B.n14 B.n13 163.367
R574 B.n592 B.n14 163.367
R575 B.n592 B.n19 163.367
R576 B.n20 B.n19 163.367
R577 B.n21 B.n20 163.367
R578 B.n597 B.n21 163.367
R579 B.n597 B.n26 163.367
R580 B.n27 B.n26 163.367
R581 B.n28 B.n27 163.367
R582 B.n602 B.n28 163.367
R583 B.n602 B.n33 163.367
R584 B.n34 B.n33 163.367
R585 B.n35 B.n34 163.367
R586 B.n607 B.n35 163.367
R587 B.n607 B.n40 163.367
R588 B.n41 B.n40 163.367
R589 B.n42 B.n41 163.367
R590 B.n88 B.n42 163.367
R591 B.n93 B.n46 163.367
R592 B.n97 B.n96 163.367
R593 B.n101 B.n100 163.367
R594 B.n105 B.n104 163.367
R595 B.n109 B.n108 163.367
R596 B.n113 B.n112 163.367
R597 B.n117 B.n116 163.367
R598 B.n121 B.n120 163.367
R599 B.n125 B.n124 163.367
R600 B.n129 B.n128 163.367
R601 B.n133 B.n132 163.367
R602 B.n137 B.n136 163.367
R603 B.n141 B.n140 163.367
R604 B.n145 B.n144 163.367
R605 B.n149 B.n148 163.367
R606 B.n153 B.n152 163.367
R607 B.n157 B.n156 163.367
R608 B.n161 B.n160 163.367
R609 B.n166 B.n165 163.367
R610 B.n170 B.n169 163.367
R611 B.n174 B.n173 163.367
R612 B.n178 B.n177 163.367
R613 B.n182 B.n181 163.367
R614 B.n187 B.n186 163.367
R615 B.n191 B.n190 163.367
R616 B.n195 B.n194 163.367
R617 B.n199 B.n198 163.367
R618 B.n203 B.n202 163.367
R619 B.n207 B.n206 163.367
R620 B.n211 B.n210 163.367
R621 B.n215 B.n214 163.367
R622 B.n219 B.n218 163.367
R623 B.n223 B.n222 163.367
R624 B.n227 B.n226 163.367
R625 B.n231 B.n230 163.367
R626 B.n235 B.n234 163.367
R627 B.n239 B.n238 163.367
R628 B.n243 B.n242 163.367
R629 B.n247 B.n246 163.367
R630 B.n251 B.n250 163.367
R631 B.n253 B.n87 163.367
R632 B.n510 B.n296 97.8863
R633 B.n616 B.n43 97.8863
R634 B.n512 B.n511 71.676
R635 B.n341 B.n300 71.676
R636 B.n504 B.n301 71.676
R637 B.n500 B.n302 71.676
R638 B.n496 B.n303 71.676
R639 B.n492 B.n304 71.676
R640 B.n488 B.n305 71.676
R641 B.n484 B.n306 71.676
R642 B.n480 B.n307 71.676
R643 B.n476 B.n308 71.676
R644 B.n472 B.n309 71.676
R645 B.n468 B.n310 71.676
R646 B.n464 B.n311 71.676
R647 B.n460 B.n312 71.676
R648 B.n456 B.n313 71.676
R649 B.n452 B.n314 71.676
R650 B.n448 B.n315 71.676
R651 B.n444 B.n316 71.676
R652 B.n440 B.n317 71.676
R653 B.n436 B.n318 71.676
R654 B.n432 B.n319 71.676
R655 B.n428 B.n320 71.676
R656 B.n424 B.n321 71.676
R657 B.n420 B.n322 71.676
R658 B.n416 B.n323 71.676
R659 B.n412 B.n324 71.676
R660 B.n408 B.n325 71.676
R661 B.n404 B.n326 71.676
R662 B.n400 B.n327 71.676
R663 B.n396 B.n328 71.676
R664 B.n392 B.n329 71.676
R665 B.n388 B.n330 71.676
R666 B.n384 B.n331 71.676
R667 B.n380 B.n332 71.676
R668 B.n376 B.n333 71.676
R669 B.n372 B.n334 71.676
R670 B.n368 B.n335 71.676
R671 B.n364 B.n336 71.676
R672 B.n360 B.n337 71.676
R673 B.n356 B.n338 71.676
R674 B.n352 B.n339 71.676
R675 B.n618 B.n617 71.676
R676 B.n93 B.n47 71.676
R677 B.n97 B.n48 71.676
R678 B.n101 B.n49 71.676
R679 B.n105 B.n50 71.676
R680 B.n109 B.n51 71.676
R681 B.n113 B.n52 71.676
R682 B.n117 B.n53 71.676
R683 B.n121 B.n54 71.676
R684 B.n125 B.n55 71.676
R685 B.n129 B.n56 71.676
R686 B.n133 B.n57 71.676
R687 B.n137 B.n58 71.676
R688 B.n141 B.n59 71.676
R689 B.n145 B.n60 71.676
R690 B.n149 B.n61 71.676
R691 B.n153 B.n62 71.676
R692 B.n157 B.n63 71.676
R693 B.n161 B.n64 71.676
R694 B.n166 B.n65 71.676
R695 B.n170 B.n66 71.676
R696 B.n174 B.n67 71.676
R697 B.n178 B.n68 71.676
R698 B.n182 B.n69 71.676
R699 B.n187 B.n70 71.676
R700 B.n191 B.n71 71.676
R701 B.n195 B.n72 71.676
R702 B.n199 B.n73 71.676
R703 B.n203 B.n74 71.676
R704 B.n207 B.n75 71.676
R705 B.n211 B.n76 71.676
R706 B.n215 B.n77 71.676
R707 B.n219 B.n78 71.676
R708 B.n223 B.n79 71.676
R709 B.n227 B.n80 71.676
R710 B.n231 B.n81 71.676
R711 B.n235 B.n82 71.676
R712 B.n239 B.n83 71.676
R713 B.n243 B.n84 71.676
R714 B.n247 B.n85 71.676
R715 B.n251 B.n86 71.676
R716 B.n615 B.n87 71.676
R717 B.n615 B.n614 71.676
R718 B.n253 B.n86 71.676
R719 B.n250 B.n85 71.676
R720 B.n246 B.n84 71.676
R721 B.n242 B.n83 71.676
R722 B.n238 B.n82 71.676
R723 B.n234 B.n81 71.676
R724 B.n230 B.n80 71.676
R725 B.n226 B.n79 71.676
R726 B.n222 B.n78 71.676
R727 B.n218 B.n77 71.676
R728 B.n214 B.n76 71.676
R729 B.n210 B.n75 71.676
R730 B.n206 B.n74 71.676
R731 B.n202 B.n73 71.676
R732 B.n198 B.n72 71.676
R733 B.n194 B.n71 71.676
R734 B.n190 B.n70 71.676
R735 B.n186 B.n69 71.676
R736 B.n181 B.n68 71.676
R737 B.n177 B.n67 71.676
R738 B.n173 B.n66 71.676
R739 B.n169 B.n65 71.676
R740 B.n165 B.n64 71.676
R741 B.n160 B.n63 71.676
R742 B.n156 B.n62 71.676
R743 B.n152 B.n61 71.676
R744 B.n148 B.n60 71.676
R745 B.n144 B.n59 71.676
R746 B.n140 B.n58 71.676
R747 B.n136 B.n57 71.676
R748 B.n132 B.n56 71.676
R749 B.n128 B.n55 71.676
R750 B.n124 B.n54 71.676
R751 B.n120 B.n53 71.676
R752 B.n116 B.n52 71.676
R753 B.n112 B.n51 71.676
R754 B.n108 B.n50 71.676
R755 B.n104 B.n49 71.676
R756 B.n100 B.n48 71.676
R757 B.n96 B.n47 71.676
R758 B.n617 B.n46 71.676
R759 B.n511 B.n299 71.676
R760 B.n505 B.n300 71.676
R761 B.n501 B.n301 71.676
R762 B.n497 B.n302 71.676
R763 B.n493 B.n303 71.676
R764 B.n489 B.n304 71.676
R765 B.n485 B.n305 71.676
R766 B.n481 B.n306 71.676
R767 B.n477 B.n307 71.676
R768 B.n473 B.n308 71.676
R769 B.n469 B.n309 71.676
R770 B.n465 B.n310 71.676
R771 B.n461 B.n311 71.676
R772 B.n457 B.n312 71.676
R773 B.n453 B.n313 71.676
R774 B.n449 B.n314 71.676
R775 B.n445 B.n315 71.676
R776 B.n441 B.n316 71.676
R777 B.n437 B.n317 71.676
R778 B.n433 B.n318 71.676
R779 B.n429 B.n319 71.676
R780 B.n425 B.n320 71.676
R781 B.n421 B.n321 71.676
R782 B.n417 B.n322 71.676
R783 B.n413 B.n323 71.676
R784 B.n409 B.n324 71.676
R785 B.n405 B.n325 71.676
R786 B.n401 B.n326 71.676
R787 B.n397 B.n327 71.676
R788 B.n393 B.n328 71.676
R789 B.n389 B.n329 71.676
R790 B.n385 B.n330 71.676
R791 B.n381 B.n331 71.676
R792 B.n377 B.n332 71.676
R793 B.n373 B.n333 71.676
R794 B.n369 B.n334 71.676
R795 B.n365 B.n335 71.676
R796 B.n361 B.n336 71.676
R797 B.n357 B.n337 71.676
R798 B.n353 B.n338 71.676
R799 B.n349 B.n339 71.676
R800 B.n347 B.n346 59.5399
R801 B.n344 B.n343 59.5399
R802 B.n163 B.n92 59.5399
R803 B.n184 B.n90 59.5399
R804 B.n517 B.n296 47.2078
R805 B.n517 B.n292 47.2078
R806 B.n524 B.n292 47.2078
R807 B.n524 B.n523 47.2078
R808 B.n530 B.n285 47.2078
R809 B.n536 B.n285 47.2078
R810 B.n536 B.n280 47.2078
R811 B.n542 B.n280 47.2078
R812 B.n542 B.n281 47.2078
R813 B.n548 B.n273 47.2078
R814 B.n554 B.n273 47.2078
R815 B.n561 B.n269 47.2078
R816 B.n561 B.n560 47.2078
R817 B.n567 B.n262 47.2078
R818 B.n574 B.n262 47.2078
R819 B.n580 B.n258 47.2078
R820 B.n580 B.n4 47.2078
R821 B.n665 B.n4 47.2078
R822 B.n665 B.n664 47.2078
R823 B.n664 B.n663 47.2078
R824 B.n663 B.n8 47.2078
R825 B.n657 B.n656 47.2078
R826 B.n656 B.n655 47.2078
R827 B.n649 B.n18 47.2078
R828 B.n649 B.n648 47.2078
R829 B.n647 B.n22 47.2078
R830 B.n641 B.n22 47.2078
R831 B.n640 B.n639 47.2078
R832 B.n639 B.n29 47.2078
R833 B.n633 B.n29 47.2078
R834 B.n633 B.n632 47.2078
R835 B.n632 B.n631 47.2078
R836 B.n625 B.n39 47.2078
R837 B.n625 B.n624 47.2078
R838 B.n624 B.n623 47.2078
R839 B.n623 B.n43 47.2078
R840 B.n574 B.t3 41.654
R841 B.n657 B.t4 41.654
R842 B.n560 B.t2 40.2656
R843 B.n18 B.t7 40.2656
R844 B.n554 B.t6 38.8771
R845 B.t0 B.n647 38.8771
R846 B.n281 B.t5 37.4887
R847 B.t1 B.n640 37.4887
R848 B.n620 B.n619 37.3078
R849 B.n613 B.n612 37.3078
R850 B.n348 B.n294 37.3078
R851 B.n514 B.n513 37.3078
R852 B.n523 B.t16 26.3811
R853 B.n39 B.t9 26.3811
R854 B.n530 B.t16 20.8273
R855 B.n631 B.t9 20.8273
R856 B.n346 B.n345 19.9763
R857 B.n343 B.n342 19.9763
R858 B.n92 B.n91 19.9763
R859 B.n90 B.n89 19.9763
R860 B B.n667 18.0485
R861 B.n619 B.n45 10.6151
R862 B.n94 B.n45 10.6151
R863 B.n95 B.n94 10.6151
R864 B.n98 B.n95 10.6151
R865 B.n99 B.n98 10.6151
R866 B.n102 B.n99 10.6151
R867 B.n103 B.n102 10.6151
R868 B.n106 B.n103 10.6151
R869 B.n107 B.n106 10.6151
R870 B.n110 B.n107 10.6151
R871 B.n111 B.n110 10.6151
R872 B.n114 B.n111 10.6151
R873 B.n115 B.n114 10.6151
R874 B.n118 B.n115 10.6151
R875 B.n119 B.n118 10.6151
R876 B.n122 B.n119 10.6151
R877 B.n123 B.n122 10.6151
R878 B.n126 B.n123 10.6151
R879 B.n127 B.n126 10.6151
R880 B.n130 B.n127 10.6151
R881 B.n131 B.n130 10.6151
R882 B.n134 B.n131 10.6151
R883 B.n135 B.n134 10.6151
R884 B.n138 B.n135 10.6151
R885 B.n139 B.n138 10.6151
R886 B.n142 B.n139 10.6151
R887 B.n143 B.n142 10.6151
R888 B.n146 B.n143 10.6151
R889 B.n147 B.n146 10.6151
R890 B.n150 B.n147 10.6151
R891 B.n151 B.n150 10.6151
R892 B.n154 B.n151 10.6151
R893 B.n155 B.n154 10.6151
R894 B.n158 B.n155 10.6151
R895 B.n159 B.n158 10.6151
R896 B.n162 B.n159 10.6151
R897 B.n167 B.n164 10.6151
R898 B.n168 B.n167 10.6151
R899 B.n171 B.n168 10.6151
R900 B.n172 B.n171 10.6151
R901 B.n175 B.n172 10.6151
R902 B.n176 B.n175 10.6151
R903 B.n179 B.n176 10.6151
R904 B.n180 B.n179 10.6151
R905 B.n183 B.n180 10.6151
R906 B.n188 B.n185 10.6151
R907 B.n189 B.n188 10.6151
R908 B.n192 B.n189 10.6151
R909 B.n193 B.n192 10.6151
R910 B.n196 B.n193 10.6151
R911 B.n197 B.n196 10.6151
R912 B.n200 B.n197 10.6151
R913 B.n201 B.n200 10.6151
R914 B.n204 B.n201 10.6151
R915 B.n205 B.n204 10.6151
R916 B.n208 B.n205 10.6151
R917 B.n209 B.n208 10.6151
R918 B.n212 B.n209 10.6151
R919 B.n213 B.n212 10.6151
R920 B.n216 B.n213 10.6151
R921 B.n217 B.n216 10.6151
R922 B.n220 B.n217 10.6151
R923 B.n221 B.n220 10.6151
R924 B.n224 B.n221 10.6151
R925 B.n225 B.n224 10.6151
R926 B.n228 B.n225 10.6151
R927 B.n229 B.n228 10.6151
R928 B.n232 B.n229 10.6151
R929 B.n233 B.n232 10.6151
R930 B.n236 B.n233 10.6151
R931 B.n237 B.n236 10.6151
R932 B.n240 B.n237 10.6151
R933 B.n241 B.n240 10.6151
R934 B.n244 B.n241 10.6151
R935 B.n245 B.n244 10.6151
R936 B.n248 B.n245 10.6151
R937 B.n249 B.n248 10.6151
R938 B.n252 B.n249 10.6151
R939 B.n254 B.n252 10.6151
R940 B.n255 B.n254 10.6151
R941 B.n613 B.n255 10.6151
R942 B.n519 B.n294 10.6151
R943 B.n520 B.n519 10.6151
R944 B.n521 B.n520 10.6151
R945 B.n521 B.n287 10.6151
R946 B.n532 B.n287 10.6151
R947 B.n533 B.n532 10.6151
R948 B.n534 B.n533 10.6151
R949 B.n534 B.n278 10.6151
R950 B.n544 B.n278 10.6151
R951 B.n545 B.n544 10.6151
R952 B.n546 B.n545 10.6151
R953 B.n546 B.n271 10.6151
R954 B.n556 B.n271 10.6151
R955 B.n557 B.n556 10.6151
R956 B.n558 B.n557 10.6151
R957 B.n558 B.n264 10.6151
R958 B.n569 B.n264 10.6151
R959 B.n570 B.n569 10.6151
R960 B.n572 B.n570 10.6151
R961 B.n572 B.n571 10.6151
R962 B.n571 B.n256 10.6151
R963 B.n583 B.n256 10.6151
R964 B.n584 B.n583 10.6151
R965 B.n585 B.n584 10.6151
R966 B.n586 B.n585 10.6151
R967 B.n588 B.n586 10.6151
R968 B.n589 B.n588 10.6151
R969 B.n590 B.n589 10.6151
R970 B.n591 B.n590 10.6151
R971 B.n593 B.n591 10.6151
R972 B.n594 B.n593 10.6151
R973 B.n595 B.n594 10.6151
R974 B.n596 B.n595 10.6151
R975 B.n598 B.n596 10.6151
R976 B.n599 B.n598 10.6151
R977 B.n600 B.n599 10.6151
R978 B.n601 B.n600 10.6151
R979 B.n603 B.n601 10.6151
R980 B.n604 B.n603 10.6151
R981 B.n605 B.n604 10.6151
R982 B.n606 B.n605 10.6151
R983 B.n608 B.n606 10.6151
R984 B.n609 B.n608 10.6151
R985 B.n610 B.n609 10.6151
R986 B.n611 B.n610 10.6151
R987 B.n612 B.n611 10.6151
R988 B.n513 B.n298 10.6151
R989 B.n508 B.n298 10.6151
R990 B.n508 B.n507 10.6151
R991 B.n507 B.n506 10.6151
R992 B.n506 B.n503 10.6151
R993 B.n503 B.n502 10.6151
R994 B.n502 B.n499 10.6151
R995 B.n499 B.n498 10.6151
R996 B.n498 B.n495 10.6151
R997 B.n495 B.n494 10.6151
R998 B.n494 B.n491 10.6151
R999 B.n491 B.n490 10.6151
R1000 B.n490 B.n487 10.6151
R1001 B.n487 B.n486 10.6151
R1002 B.n486 B.n483 10.6151
R1003 B.n483 B.n482 10.6151
R1004 B.n482 B.n479 10.6151
R1005 B.n479 B.n478 10.6151
R1006 B.n478 B.n475 10.6151
R1007 B.n475 B.n474 10.6151
R1008 B.n474 B.n471 10.6151
R1009 B.n471 B.n470 10.6151
R1010 B.n470 B.n467 10.6151
R1011 B.n467 B.n466 10.6151
R1012 B.n466 B.n463 10.6151
R1013 B.n463 B.n462 10.6151
R1014 B.n462 B.n459 10.6151
R1015 B.n459 B.n458 10.6151
R1016 B.n458 B.n455 10.6151
R1017 B.n455 B.n454 10.6151
R1018 B.n454 B.n451 10.6151
R1019 B.n451 B.n450 10.6151
R1020 B.n450 B.n447 10.6151
R1021 B.n447 B.n446 10.6151
R1022 B.n446 B.n443 10.6151
R1023 B.n443 B.n442 10.6151
R1024 B.n439 B.n438 10.6151
R1025 B.n438 B.n435 10.6151
R1026 B.n435 B.n434 10.6151
R1027 B.n434 B.n431 10.6151
R1028 B.n431 B.n430 10.6151
R1029 B.n430 B.n427 10.6151
R1030 B.n427 B.n426 10.6151
R1031 B.n426 B.n423 10.6151
R1032 B.n423 B.n422 10.6151
R1033 B.n419 B.n418 10.6151
R1034 B.n418 B.n415 10.6151
R1035 B.n415 B.n414 10.6151
R1036 B.n414 B.n411 10.6151
R1037 B.n411 B.n410 10.6151
R1038 B.n410 B.n407 10.6151
R1039 B.n407 B.n406 10.6151
R1040 B.n406 B.n403 10.6151
R1041 B.n403 B.n402 10.6151
R1042 B.n402 B.n399 10.6151
R1043 B.n399 B.n398 10.6151
R1044 B.n398 B.n395 10.6151
R1045 B.n395 B.n394 10.6151
R1046 B.n394 B.n391 10.6151
R1047 B.n391 B.n390 10.6151
R1048 B.n390 B.n387 10.6151
R1049 B.n387 B.n386 10.6151
R1050 B.n386 B.n383 10.6151
R1051 B.n383 B.n382 10.6151
R1052 B.n382 B.n379 10.6151
R1053 B.n379 B.n378 10.6151
R1054 B.n378 B.n375 10.6151
R1055 B.n375 B.n374 10.6151
R1056 B.n374 B.n371 10.6151
R1057 B.n371 B.n370 10.6151
R1058 B.n370 B.n367 10.6151
R1059 B.n367 B.n366 10.6151
R1060 B.n366 B.n363 10.6151
R1061 B.n363 B.n362 10.6151
R1062 B.n362 B.n359 10.6151
R1063 B.n359 B.n358 10.6151
R1064 B.n358 B.n355 10.6151
R1065 B.n355 B.n354 10.6151
R1066 B.n354 B.n351 10.6151
R1067 B.n351 B.n350 10.6151
R1068 B.n350 B.n348 10.6151
R1069 B.n515 B.n514 10.6151
R1070 B.n515 B.n290 10.6151
R1071 B.n526 B.n290 10.6151
R1072 B.n527 B.n526 10.6151
R1073 B.n528 B.n527 10.6151
R1074 B.n528 B.n283 10.6151
R1075 B.n538 B.n283 10.6151
R1076 B.n539 B.n538 10.6151
R1077 B.n540 B.n539 10.6151
R1078 B.n540 B.n275 10.6151
R1079 B.n550 B.n275 10.6151
R1080 B.n551 B.n550 10.6151
R1081 B.n552 B.n551 10.6151
R1082 B.n552 B.n267 10.6151
R1083 B.n563 B.n267 10.6151
R1084 B.n564 B.n563 10.6151
R1085 B.n565 B.n564 10.6151
R1086 B.n565 B.n260 10.6151
R1087 B.n576 B.n260 10.6151
R1088 B.n577 B.n576 10.6151
R1089 B.n578 B.n577 10.6151
R1090 B.n578 B.n0 10.6151
R1091 B.n661 B.n1 10.6151
R1092 B.n661 B.n660 10.6151
R1093 B.n660 B.n659 10.6151
R1094 B.n659 B.n10 10.6151
R1095 B.n653 B.n10 10.6151
R1096 B.n653 B.n652 10.6151
R1097 B.n652 B.n651 10.6151
R1098 B.n651 B.n16 10.6151
R1099 B.n645 B.n16 10.6151
R1100 B.n645 B.n644 10.6151
R1101 B.n644 B.n643 10.6151
R1102 B.n643 B.n24 10.6151
R1103 B.n637 B.n24 10.6151
R1104 B.n637 B.n636 10.6151
R1105 B.n636 B.n635 10.6151
R1106 B.n635 B.n31 10.6151
R1107 B.n629 B.n31 10.6151
R1108 B.n629 B.n628 10.6151
R1109 B.n628 B.n627 10.6151
R1110 B.n627 B.n37 10.6151
R1111 B.n621 B.n37 10.6151
R1112 B.n621 B.n620 10.6151
R1113 B.n548 B.t5 9.71965
R1114 B.n641 B.t1 9.71965
R1115 B.n163 B.n162 9.36635
R1116 B.n185 B.n184 9.36635
R1117 B.n442 B.n344 9.36635
R1118 B.n419 B.n347 9.36635
R1119 B.t6 B.n269 8.3312
R1120 B.n648 B.t0 8.3312
R1121 B.n567 B.t2 6.94275
R1122 B.n655 B.t7 6.94275
R1123 B.t3 B.n258 5.5543
R1124 B.t4 B.n8 5.5543
R1125 B.n667 B.n0 2.81026
R1126 B.n667 B.n1 2.81026
R1127 B.n164 B.n163 1.24928
R1128 B.n184 B.n183 1.24928
R1129 B.n439 B.n344 1.24928
R1130 B.n422 B.n347 1.24928
R1131 VP.n6 VP.t1 442.551
R1132 VP.n14 VP.t2 420.373
R1133 VP.n16 VP.t5 420.373
R1134 VP.n20 VP.t7 420.373
R1135 VP.n22 VP.t6 420.373
R1136 VP.n11 VP.t3 420.373
R1137 VP.n9 VP.t0 420.373
R1138 VP.n5 VP.t4 420.373
R1139 VP.n23 VP.n22 161.3
R1140 VP.n8 VP.n7 161.3
R1141 VP.n9 VP.n4 161.3
R1142 VP.n10 VP.n3 161.3
R1143 VP.n12 VP.n11 161.3
R1144 VP.n21 VP.n0 161.3
R1145 VP.n20 VP.n19 161.3
R1146 VP.n18 VP.n1 161.3
R1147 VP.n17 VP.n16 161.3
R1148 VP.n15 VP.n2 161.3
R1149 VP.n14 VP.n13 161.3
R1150 VP.n7 VP.n6 44.862
R1151 VP.n13 VP.n12 40.9096
R1152 VP.n15 VP.n14 28.4823
R1153 VP.n22 VP.n21 28.4823
R1154 VP.n11 VP.n10 28.4823
R1155 VP.n16 VP.n1 24.1005
R1156 VP.n20 VP.n1 24.1005
R1157 VP.n8 VP.n5 24.1005
R1158 VP.n9 VP.n8 24.1005
R1159 VP.n16 VP.n15 19.7187
R1160 VP.n21 VP.n20 19.7187
R1161 VP.n10 VP.n9 19.7187
R1162 VP.n6 VP.n5 19.7081
R1163 VP.n7 VP.n4 0.189894
R1164 VP.n4 VP.n3 0.189894
R1165 VP.n12 VP.n3 0.189894
R1166 VP.n13 VP.n2 0.189894
R1167 VP.n17 VP.n2 0.189894
R1168 VP.n18 VP.n17 0.189894
R1169 VP.n19 VP.n18 0.189894
R1170 VP.n19 VP.n0 0.189894
R1171 VP.n23 VP.n0 0.189894
R1172 VP VP.n23 0.0516364
R1173 VDD1 VDD1.n0 60.7091
R1174 VDD1.n3 VDD1.n2 60.5954
R1175 VDD1.n3 VDD1.n1 60.5954
R1176 VDD1.n5 VDD1.n4 60.2068
R1177 VDD1.n5 VDD1.n3 37.4061
R1178 VDD1.n4 VDD1.t6 1.87373
R1179 VDD1.n4 VDD1.t7 1.87373
R1180 VDD1.n0 VDD1.t0 1.87373
R1181 VDD1.n0 VDD1.t5 1.87373
R1182 VDD1.n2 VDD1.t2 1.87373
R1183 VDD1.n2 VDD1.t3 1.87373
R1184 VDD1.n1 VDD1.t1 1.87373
R1185 VDD1.n1 VDD1.t4 1.87373
R1186 VDD1 VDD1.n5 0.386276
R1187 VTAIL.n466 VTAIL.n414 289.615
R1188 VTAIL.n54 VTAIL.n2 289.615
R1189 VTAIL.n112 VTAIL.n60 289.615
R1190 VTAIL.n172 VTAIL.n120 289.615
R1191 VTAIL.n408 VTAIL.n356 289.615
R1192 VTAIL.n348 VTAIL.n296 289.615
R1193 VTAIL.n290 VTAIL.n238 289.615
R1194 VTAIL.n230 VTAIL.n178 289.615
R1195 VTAIL.n433 VTAIL.n432 185
R1196 VTAIL.n430 VTAIL.n429 185
R1197 VTAIL.n439 VTAIL.n438 185
R1198 VTAIL.n441 VTAIL.n440 185
R1199 VTAIL.n426 VTAIL.n425 185
R1200 VTAIL.n447 VTAIL.n446 185
R1201 VTAIL.n450 VTAIL.n449 185
R1202 VTAIL.n448 VTAIL.n422 185
R1203 VTAIL.n455 VTAIL.n421 185
R1204 VTAIL.n457 VTAIL.n456 185
R1205 VTAIL.n459 VTAIL.n458 185
R1206 VTAIL.n418 VTAIL.n417 185
R1207 VTAIL.n465 VTAIL.n464 185
R1208 VTAIL.n467 VTAIL.n466 185
R1209 VTAIL.n21 VTAIL.n20 185
R1210 VTAIL.n18 VTAIL.n17 185
R1211 VTAIL.n27 VTAIL.n26 185
R1212 VTAIL.n29 VTAIL.n28 185
R1213 VTAIL.n14 VTAIL.n13 185
R1214 VTAIL.n35 VTAIL.n34 185
R1215 VTAIL.n38 VTAIL.n37 185
R1216 VTAIL.n36 VTAIL.n10 185
R1217 VTAIL.n43 VTAIL.n9 185
R1218 VTAIL.n45 VTAIL.n44 185
R1219 VTAIL.n47 VTAIL.n46 185
R1220 VTAIL.n6 VTAIL.n5 185
R1221 VTAIL.n53 VTAIL.n52 185
R1222 VTAIL.n55 VTAIL.n54 185
R1223 VTAIL.n79 VTAIL.n78 185
R1224 VTAIL.n76 VTAIL.n75 185
R1225 VTAIL.n85 VTAIL.n84 185
R1226 VTAIL.n87 VTAIL.n86 185
R1227 VTAIL.n72 VTAIL.n71 185
R1228 VTAIL.n93 VTAIL.n92 185
R1229 VTAIL.n96 VTAIL.n95 185
R1230 VTAIL.n94 VTAIL.n68 185
R1231 VTAIL.n101 VTAIL.n67 185
R1232 VTAIL.n103 VTAIL.n102 185
R1233 VTAIL.n105 VTAIL.n104 185
R1234 VTAIL.n64 VTAIL.n63 185
R1235 VTAIL.n111 VTAIL.n110 185
R1236 VTAIL.n113 VTAIL.n112 185
R1237 VTAIL.n139 VTAIL.n138 185
R1238 VTAIL.n136 VTAIL.n135 185
R1239 VTAIL.n145 VTAIL.n144 185
R1240 VTAIL.n147 VTAIL.n146 185
R1241 VTAIL.n132 VTAIL.n131 185
R1242 VTAIL.n153 VTAIL.n152 185
R1243 VTAIL.n156 VTAIL.n155 185
R1244 VTAIL.n154 VTAIL.n128 185
R1245 VTAIL.n161 VTAIL.n127 185
R1246 VTAIL.n163 VTAIL.n162 185
R1247 VTAIL.n165 VTAIL.n164 185
R1248 VTAIL.n124 VTAIL.n123 185
R1249 VTAIL.n171 VTAIL.n170 185
R1250 VTAIL.n173 VTAIL.n172 185
R1251 VTAIL.n409 VTAIL.n408 185
R1252 VTAIL.n407 VTAIL.n406 185
R1253 VTAIL.n360 VTAIL.n359 185
R1254 VTAIL.n401 VTAIL.n400 185
R1255 VTAIL.n399 VTAIL.n398 185
R1256 VTAIL.n397 VTAIL.n363 185
R1257 VTAIL.n367 VTAIL.n364 185
R1258 VTAIL.n392 VTAIL.n391 185
R1259 VTAIL.n390 VTAIL.n389 185
R1260 VTAIL.n369 VTAIL.n368 185
R1261 VTAIL.n384 VTAIL.n383 185
R1262 VTAIL.n382 VTAIL.n381 185
R1263 VTAIL.n373 VTAIL.n372 185
R1264 VTAIL.n376 VTAIL.n375 185
R1265 VTAIL.n349 VTAIL.n348 185
R1266 VTAIL.n347 VTAIL.n346 185
R1267 VTAIL.n300 VTAIL.n299 185
R1268 VTAIL.n341 VTAIL.n340 185
R1269 VTAIL.n339 VTAIL.n338 185
R1270 VTAIL.n337 VTAIL.n303 185
R1271 VTAIL.n307 VTAIL.n304 185
R1272 VTAIL.n332 VTAIL.n331 185
R1273 VTAIL.n330 VTAIL.n329 185
R1274 VTAIL.n309 VTAIL.n308 185
R1275 VTAIL.n324 VTAIL.n323 185
R1276 VTAIL.n322 VTAIL.n321 185
R1277 VTAIL.n313 VTAIL.n312 185
R1278 VTAIL.n316 VTAIL.n315 185
R1279 VTAIL.n291 VTAIL.n290 185
R1280 VTAIL.n289 VTAIL.n288 185
R1281 VTAIL.n242 VTAIL.n241 185
R1282 VTAIL.n283 VTAIL.n282 185
R1283 VTAIL.n281 VTAIL.n280 185
R1284 VTAIL.n279 VTAIL.n245 185
R1285 VTAIL.n249 VTAIL.n246 185
R1286 VTAIL.n274 VTAIL.n273 185
R1287 VTAIL.n272 VTAIL.n271 185
R1288 VTAIL.n251 VTAIL.n250 185
R1289 VTAIL.n266 VTAIL.n265 185
R1290 VTAIL.n264 VTAIL.n263 185
R1291 VTAIL.n255 VTAIL.n254 185
R1292 VTAIL.n258 VTAIL.n257 185
R1293 VTAIL.n231 VTAIL.n230 185
R1294 VTAIL.n229 VTAIL.n228 185
R1295 VTAIL.n182 VTAIL.n181 185
R1296 VTAIL.n223 VTAIL.n222 185
R1297 VTAIL.n221 VTAIL.n220 185
R1298 VTAIL.n219 VTAIL.n185 185
R1299 VTAIL.n189 VTAIL.n186 185
R1300 VTAIL.n214 VTAIL.n213 185
R1301 VTAIL.n212 VTAIL.n211 185
R1302 VTAIL.n191 VTAIL.n190 185
R1303 VTAIL.n206 VTAIL.n205 185
R1304 VTAIL.n204 VTAIL.n203 185
R1305 VTAIL.n195 VTAIL.n194 185
R1306 VTAIL.n198 VTAIL.n197 185
R1307 VTAIL.t0 VTAIL.n431 149.524
R1308 VTAIL.t5 VTAIL.n19 149.524
R1309 VTAIL.t9 VTAIL.n77 149.524
R1310 VTAIL.t13 VTAIL.n137 149.524
R1311 VTAIL.t12 VTAIL.n374 149.524
R1312 VTAIL.t14 VTAIL.n314 149.524
R1313 VTAIL.t4 VTAIL.n256 149.524
R1314 VTAIL.t2 VTAIL.n196 149.524
R1315 VTAIL.n432 VTAIL.n429 104.615
R1316 VTAIL.n439 VTAIL.n429 104.615
R1317 VTAIL.n440 VTAIL.n439 104.615
R1318 VTAIL.n440 VTAIL.n425 104.615
R1319 VTAIL.n447 VTAIL.n425 104.615
R1320 VTAIL.n449 VTAIL.n447 104.615
R1321 VTAIL.n449 VTAIL.n448 104.615
R1322 VTAIL.n448 VTAIL.n421 104.615
R1323 VTAIL.n457 VTAIL.n421 104.615
R1324 VTAIL.n458 VTAIL.n457 104.615
R1325 VTAIL.n458 VTAIL.n417 104.615
R1326 VTAIL.n465 VTAIL.n417 104.615
R1327 VTAIL.n466 VTAIL.n465 104.615
R1328 VTAIL.n20 VTAIL.n17 104.615
R1329 VTAIL.n27 VTAIL.n17 104.615
R1330 VTAIL.n28 VTAIL.n27 104.615
R1331 VTAIL.n28 VTAIL.n13 104.615
R1332 VTAIL.n35 VTAIL.n13 104.615
R1333 VTAIL.n37 VTAIL.n35 104.615
R1334 VTAIL.n37 VTAIL.n36 104.615
R1335 VTAIL.n36 VTAIL.n9 104.615
R1336 VTAIL.n45 VTAIL.n9 104.615
R1337 VTAIL.n46 VTAIL.n45 104.615
R1338 VTAIL.n46 VTAIL.n5 104.615
R1339 VTAIL.n53 VTAIL.n5 104.615
R1340 VTAIL.n54 VTAIL.n53 104.615
R1341 VTAIL.n78 VTAIL.n75 104.615
R1342 VTAIL.n85 VTAIL.n75 104.615
R1343 VTAIL.n86 VTAIL.n85 104.615
R1344 VTAIL.n86 VTAIL.n71 104.615
R1345 VTAIL.n93 VTAIL.n71 104.615
R1346 VTAIL.n95 VTAIL.n93 104.615
R1347 VTAIL.n95 VTAIL.n94 104.615
R1348 VTAIL.n94 VTAIL.n67 104.615
R1349 VTAIL.n103 VTAIL.n67 104.615
R1350 VTAIL.n104 VTAIL.n103 104.615
R1351 VTAIL.n104 VTAIL.n63 104.615
R1352 VTAIL.n111 VTAIL.n63 104.615
R1353 VTAIL.n112 VTAIL.n111 104.615
R1354 VTAIL.n138 VTAIL.n135 104.615
R1355 VTAIL.n145 VTAIL.n135 104.615
R1356 VTAIL.n146 VTAIL.n145 104.615
R1357 VTAIL.n146 VTAIL.n131 104.615
R1358 VTAIL.n153 VTAIL.n131 104.615
R1359 VTAIL.n155 VTAIL.n153 104.615
R1360 VTAIL.n155 VTAIL.n154 104.615
R1361 VTAIL.n154 VTAIL.n127 104.615
R1362 VTAIL.n163 VTAIL.n127 104.615
R1363 VTAIL.n164 VTAIL.n163 104.615
R1364 VTAIL.n164 VTAIL.n123 104.615
R1365 VTAIL.n171 VTAIL.n123 104.615
R1366 VTAIL.n172 VTAIL.n171 104.615
R1367 VTAIL.n408 VTAIL.n407 104.615
R1368 VTAIL.n407 VTAIL.n359 104.615
R1369 VTAIL.n400 VTAIL.n359 104.615
R1370 VTAIL.n400 VTAIL.n399 104.615
R1371 VTAIL.n399 VTAIL.n363 104.615
R1372 VTAIL.n367 VTAIL.n363 104.615
R1373 VTAIL.n391 VTAIL.n367 104.615
R1374 VTAIL.n391 VTAIL.n390 104.615
R1375 VTAIL.n390 VTAIL.n368 104.615
R1376 VTAIL.n383 VTAIL.n368 104.615
R1377 VTAIL.n383 VTAIL.n382 104.615
R1378 VTAIL.n382 VTAIL.n372 104.615
R1379 VTAIL.n375 VTAIL.n372 104.615
R1380 VTAIL.n348 VTAIL.n347 104.615
R1381 VTAIL.n347 VTAIL.n299 104.615
R1382 VTAIL.n340 VTAIL.n299 104.615
R1383 VTAIL.n340 VTAIL.n339 104.615
R1384 VTAIL.n339 VTAIL.n303 104.615
R1385 VTAIL.n307 VTAIL.n303 104.615
R1386 VTAIL.n331 VTAIL.n307 104.615
R1387 VTAIL.n331 VTAIL.n330 104.615
R1388 VTAIL.n330 VTAIL.n308 104.615
R1389 VTAIL.n323 VTAIL.n308 104.615
R1390 VTAIL.n323 VTAIL.n322 104.615
R1391 VTAIL.n322 VTAIL.n312 104.615
R1392 VTAIL.n315 VTAIL.n312 104.615
R1393 VTAIL.n290 VTAIL.n289 104.615
R1394 VTAIL.n289 VTAIL.n241 104.615
R1395 VTAIL.n282 VTAIL.n241 104.615
R1396 VTAIL.n282 VTAIL.n281 104.615
R1397 VTAIL.n281 VTAIL.n245 104.615
R1398 VTAIL.n249 VTAIL.n245 104.615
R1399 VTAIL.n273 VTAIL.n249 104.615
R1400 VTAIL.n273 VTAIL.n272 104.615
R1401 VTAIL.n272 VTAIL.n250 104.615
R1402 VTAIL.n265 VTAIL.n250 104.615
R1403 VTAIL.n265 VTAIL.n264 104.615
R1404 VTAIL.n264 VTAIL.n254 104.615
R1405 VTAIL.n257 VTAIL.n254 104.615
R1406 VTAIL.n230 VTAIL.n229 104.615
R1407 VTAIL.n229 VTAIL.n181 104.615
R1408 VTAIL.n222 VTAIL.n181 104.615
R1409 VTAIL.n222 VTAIL.n221 104.615
R1410 VTAIL.n221 VTAIL.n185 104.615
R1411 VTAIL.n189 VTAIL.n185 104.615
R1412 VTAIL.n213 VTAIL.n189 104.615
R1413 VTAIL.n213 VTAIL.n212 104.615
R1414 VTAIL.n212 VTAIL.n190 104.615
R1415 VTAIL.n205 VTAIL.n190 104.615
R1416 VTAIL.n205 VTAIL.n204 104.615
R1417 VTAIL.n204 VTAIL.n194 104.615
R1418 VTAIL.n197 VTAIL.n194 104.615
R1419 VTAIL.n432 VTAIL.t0 52.3082
R1420 VTAIL.n20 VTAIL.t5 52.3082
R1421 VTAIL.n78 VTAIL.t9 52.3082
R1422 VTAIL.n138 VTAIL.t13 52.3082
R1423 VTAIL.n375 VTAIL.t12 52.3082
R1424 VTAIL.n315 VTAIL.t14 52.3082
R1425 VTAIL.n257 VTAIL.t4 52.3082
R1426 VTAIL.n197 VTAIL.t2 52.3082
R1427 VTAIL.n355 VTAIL.n354 43.5282
R1428 VTAIL.n237 VTAIL.n236 43.5282
R1429 VTAIL.n1 VTAIL.n0 43.528
R1430 VTAIL.n119 VTAIL.n118 43.528
R1431 VTAIL.n471 VTAIL.n470 30.052
R1432 VTAIL.n59 VTAIL.n58 30.052
R1433 VTAIL.n117 VTAIL.n116 30.052
R1434 VTAIL.n177 VTAIL.n176 30.052
R1435 VTAIL.n413 VTAIL.n412 30.052
R1436 VTAIL.n353 VTAIL.n352 30.052
R1437 VTAIL.n295 VTAIL.n294 30.052
R1438 VTAIL.n235 VTAIL.n234 30.052
R1439 VTAIL.n471 VTAIL.n413 22.3669
R1440 VTAIL.n235 VTAIL.n177 22.3669
R1441 VTAIL.n456 VTAIL.n455 13.1884
R1442 VTAIL.n44 VTAIL.n43 13.1884
R1443 VTAIL.n102 VTAIL.n101 13.1884
R1444 VTAIL.n162 VTAIL.n161 13.1884
R1445 VTAIL.n398 VTAIL.n397 13.1884
R1446 VTAIL.n338 VTAIL.n337 13.1884
R1447 VTAIL.n280 VTAIL.n279 13.1884
R1448 VTAIL.n220 VTAIL.n219 13.1884
R1449 VTAIL.n454 VTAIL.n422 12.8005
R1450 VTAIL.n459 VTAIL.n420 12.8005
R1451 VTAIL.n42 VTAIL.n10 12.8005
R1452 VTAIL.n47 VTAIL.n8 12.8005
R1453 VTAIL.n100 VTAIL.n68 12.8005
R1454 VTAIL.n105 VTAIL.n66 12.8005
R1455 VTAIL.n160 VTAIL.n128 12.8005
R1456 VTAIL.n165 VTAIL.n126 12.8005
R1457 VTAIL.n401 VTAIL.n362 12.8005
R1458 VTAIL.n396 VTAIL.n364 12.8005
R1459 VTAIL.n341 VTAIL.n302 12.8005
R1460 VTAIL.n336 VTAIL.n304 12.8005
R1461 VTAIL.n283 VTAIL.n244 12.8005
R1462 VTAIL.n278 VTAIL.n246 12.8005
R1463 VTAIL.n223 VTAIL.n184 12.8005
R1464 VTAIL.n218 VTAIL.n186 12.8005
R1465 VTAIL.n451 VTAIL.n450 12.0247
R1466 VTAIL.n460 VTAIL.n418 12.0247
R1467 VTAIL.n39 VTAIL.n38 12.0247
R1468 VTAIL.n48 VTAIL.n6 12.0247
R1469 VTAIL.n97 VTAIL.n96 12.0247
R1470 VTAIL.n106 VTAIL.n64 12.0247
R1471 VTAIL.n157 VTAIL.n156 12.0247
R1472 VTAIL.n166 VTAIL.n124 12.0247
R1473 VTAIL.n402 VTAIL.n360 12.0247
R1474 VTAIL.n393 VTAIL.n392 12.0247
R1475 VTAIL.n342 VTAIL.n300 12.0247
R1476 VTAIL.n333 VTAIL.n332 12.0247
R1477 VTAIL.n284 VTAIL.n242 12.0247
R1478 VTAIL.n275 VTAIL.n274 12.0247
R1479 VTAIL.n224 VTAIL.n182 12.0247
R1480 VTAIL.n215 VTAIL.n214 12.0247
R1481 VTAIL.n446 VTAIL.n424 11.249
R1482 VTAIL.n464 VTAIL.n463 11.249
R1483 VTAIL.n34 VTAIL.n12 11.249
R1484 VTAIL.n52 VTAIL.n51 11.249
R1485 VTAIL.n92 VTAIL.n70 11.249
R1486 VTAIL.n110 VTAIL.n109 11.249
R1487 VTAIL.n152 VTAIL.n130 11.249
R1488 VTAIL.n170 VTAIL.n169 11.249
R1489 VTAIL.n406 VTAIL.n405 11.249
R1490 VTAIL.n389 VTAIL.n366 11.249
R1491 VTAIL.n346 VTAIL.n345 11.249
R1492 VTAIL.n329 VTAIL.n306 11.249
R1493 VTAIL.n288 VTAIL.n287 11.249
R1494 VTAIL.n271 VTAIL.n248 11.249
R1495 VTAIL.n228 VTAIL.n227 11.249
R1496 VTAIL.n211 VTAIL.n188 11.249
R1497 VTAIL.n445 VTAIL.n426 10.4732
R1498 VTAIL.n467 VTAIL.n416 10.4732
R1499 VTAIL.n33 VTAIL.n14 10.4732
R1500 VTAIL.n55 VTAIL.n4 10.4732
R1501 VTAIL.n91 VTAIL.n72 10.4732
R1502 VTAIL.n113 VTAIL.n62 10.4732
R1503 VTAIL.n151 VTAIL.n132 10.4732
R1504 VTAIL.n173 VTAIL.n122 10.4732
R1505 VTAIL.n409 VTAIL.n358 10.4732
R1506 VTAIL.n388 VTAIL.n369 10.4732
R1507 VTAIL.n349 VTAIL.n298 10.4732
R1508 VTAIL.n328 VTAIL.n309 10.4732
R1509 VTAIL.n291 VTAIL.n240 10.4732
R1510 VTAIL.n270 VTAIL.n251 10.4732
R1511 VTAIL.n231 VTAIL.n180 10.4732
R1512 VTAIL.n210 VTAIL.n191 10.4732
R1513 VTAIL.n433 VTAIL.n431 10.2747
R1514 VTAIL.n21 VTAIL.n19 10.2747
R1515 VTAIL.n79 VTAIL.n77 10.2747
R1516 VTAIL.n139 VTAIL.n137 10.2747
R1517 VTAIL.n376 VTAIL.n374 10.2747
R1518 VTAIL.n316 VTAIL.n314 10.2747
R1519 VTAIL.n258 VTAIL.n256 10.2747
R1520 VTAIL.n198 VTAIL.n196 10.2747
R1521 VTAIL.n442 VTAIL.n441 9.69747
R1522 VTAIL.n468 VTAIL.n414 9.69747
R1523 VTAIL.n30 VTAIL.n29 9.69747
R1524 VTAIL.n56 VTAIL.n2 9.69747
R1525 VTAIL.n88 VTAIL.n87 9.69747
R1526 VTAIL.n114 VTAIL.n60 9.69747
R1527 VTAIL.n148 VTAIL.n147 9.69747
R1528 VTAIL.n174 VTAIL.n120 9.69747
R1529 VTAIL.n410 VTAIL.n356 9.69747
R1530 VTAIL.n385 VTAIL.n384 9.69747
R1531 VTAIL.n350 VTAIL.n296 9.69747
R1532 VTAIL.n325 VTAIL.n324 9.69747
R1533 VTAIL.n292 VTAIL.n238 9.69747
R1534 VTAIL.n267 VTAIL.n266 9.69747
R1535 VTAIL.n232 VTAIL.n178 9.69747
R1536 VTAIL.n207 VTAIL.n206 9.69747
R1537 VTAIL.n470 VTAIL.n469 9.45567
R1538 VTAIL.n58 VTAIL.n57 9.45567
R1539 VTAIL.n116 VTAIL.n115 9.45567
R1540 VTAIL.n176 VTAIL.n175 9.45567
R1541 VTAIL.n412 VTAIL.n411 9.45567
R1542 VTAIL.n352 VTAIL.n351 9.45567
R1543 VTAIL.n294 VTAIL.n293 9.45567
R1544 VTAIL.n234 VTAIL.n233 9.45567
R1545 VTAIL.n469 VTAIL.n468 9.3005
R1546 VTAIL.n416 VTAIL.n415 9.3005
R1547 VTAIL.n463 VTAIL.n462 9.3005
R1548 VTAIL.n461 VTAIL.n460 9.3005
R1549 VTAIL.n420 VTAIL.n419 9.3005
R1550 VTAIL.n435 VTAIL.n434 9.3005
R1551 VTAIL.n437 VTAIL.n436 9.3005
R1552 VTAIL.n428 VTAIL.n427 9.3005
R1553 VTAIL.n443 VTAIL.n442 9.3005
R1554 VTAIL.n445 VTAIL.n444 9.3005
R1555 VTAIL.n424 VTAIL.n423 9.3005
R1556 VTAIL.n452 VTAIL.n451 9.3005
R1557 VTAIL.n454 VTAIL.n453 9.3005
R1558 VTAIL.n57 VTAIL.n56 9.3005
R1559 VTAIL.n4 VTAIL.n3 9.3005
R1560 VTAIL.n51 VTAIL.n50 9.3005
R1561 VTAIL.n49 VTAIL.n48 9.3005
R1562 VTAIL.n8 VTAIL.n7 9.3005
R1563 VTAIL.n23 VTAIL.n22 9.3005
R1564 VTAIL.n25 VTAIL.n24 9.3005
R1565 VTAIL.n16 VTAIL.n15 9.3005
R1566 VTAIL.n31 VTAIL.n30 9.3005
R1567 VTAIL.n33 VTAIL.n32 9.3005
R1568 VTAIL.n12 VTAIL.n11 9.3005
R1569 VTAIL.n40 VTAIL.n39 9.3005
R1570 VTAIL.n42 VTAIL.n41 9.3005
R1571 VTAIL.n115 VTAIL.n114 9.3005
R1572 VTAIL.n62 VTAIL.n61 9.3005
R1573 VTAIL.n109 VTAIL.n108 9.3005
R1574 VTAIL.n107 VTAIL.n106 9.3005
R1575 VTAIL.n66 VTAIL.n65 9.3005
R1576 VTAIL.n81 VTAIL.n80 9.3005
R1577 VTAIL.n83 VTAIL.n82 9.3005
R1578 VTAIL.n74 VTAIL.n73 9.3005
R1579 VTAIL.n89 VTAIL.n88 9.3005
R1580 VTAIL.n91 VTAIL.n90 9.3005
R1581 VTAIL.n70 VTAIL.n69 9.3005
R1582 VTAIL.n98 VTAIL.n97 9.3005
R1583 VTAIL.n100 VTAIL.n99 9.3005
R1584 VTAIL.n175 VTAIL.n174 9.3005
R1585 VTAIL.n122 VTAIL.n121 9.3005
R1586 VTAIL.n169 VTAIL.n168 9.3005
R1587 VTAIL.n167 VTAIL.n166 9.3005
R1588 VTAIL.n126 VTAIL.n125 9.3005
R1589 VTAIL.n141 VTAIL.n140 9.3005
R1590 VTAIL.n143 VTAIL.n142 9.3005
R1591 VTAIL.n134 VTAIL.n133 9.3005
R1592 VTAIL.n149 VTAIL.n148 9.3005
R1593 VTAIL.n151 VTAIL.n150 9.3005
R1594 VTAIL.n130 VTAIL.n129 9.3005
R1595 VTAIL.n158 VTAIL.n157 9.3005
R1596 VTAIL.n160 VTAIL.n159 9.3005
R1597 VTAIL.n378 VTAIL.n377 9.3005
R1598 VTAIL.n380 VTAIL.n379 9.3005
R1599 VTAIL.n371 VTAIL.n370 9.3005
R1600 VTAIL.n386 VTAIL.n385 9.3005
R1601 VTAIL.n388 VTAIL.n387 9.3005
R1602 VTAIL.n366 VTAIL.n365 9.3005
R1603 VTAIL.n394 VTAIL.n393 9.3005
R1604 VTAIL.n396 VTAIL.n395 9.3005
R1605 VTAIL.n411 VTAIL.n410 9.3005
R1606 VTAIL.n358 VTAIL.n357 9.3005
R1607 VTAIL.n405 VTAIL.n404 9.3005
R1608 VTAIL.n403 VTAIL.n402 9.3005
R1609 VTAIL.n362 VTAIL.n361 9.3005
R1610 VTAIL.n318 VTAIL.n317 9.3005
R1611 VTAIL.n320 VTAIL.n319 9.3005
R1612 VTAIL.n311 VTAIL.n310 9.3005
R1613 VTAIL.n326 VTAIL.n325 9.3005
R1614 VTAIL.n328 VTAIL.n327 9.3005
R1615 VTAIL.n306 VTAIL.n305 9.3005
R1616 VTAIL.n334 VTAIL.n333 9.3005
R1617 VTAIL.n336 VTAIL.n335 9.3005
R1618 VTAIL.n351 VTAIL.n350 9.3005
R1619 VTAIL.n298 VTAIL.n297 9.3005
R1620 VTAIL.n345 VTAIL.n344 9.3005
R1621 VTAIL.n343 VTAIL.n342 9.3005
R1622 VTAIL.n302 VTAIL.n301 9.3005
R1623 VTAIL.n260 VTAIL.n259 9.3005
R1624 VTAIL.n262 VTAIL.n261 9.3005
R1625 VTAIL.n253 VTAIL.n252 9.3005
R1626 VTAIL.n268 VTAIL.n267 9.3005
R1627 VTAIL.n270 VTAIL.n269 9.3005
R1628 VTAIL.n248 VTAIL.n247 9.3005
R1629 VTAIL.n276 VTAIL.n275 9.3005
R1630 VTAIL.n278 VTAIL.n277 9.3005
R1631 VTAIL.n293 VTAIL.n292 9.3005
R1632 VTAIL.n240 VTAIL.n239 9.3005
R1633 VTAIL.n287 VTAIL.n286 9.3005
R1634 VTAIL.n285 VTAIL.n284 9.3005
R1635 VTAIL.n244 VTAIL.n243 9.3005
R1636 VTAIL.n200 VTAIL.n199 9.3005
R1637 VTAIL.n202 VTAIL.n201 9.3005
R1638 VTAIL.n193 VTAIL.n192 9.3005
R1639 VTAIL.n208 VTAIL.n207 9.3005
R1640 VTAIL.n210 VTAIL.n209 9.3005
R1641 VTAIL.n188 VTAIL.n187 9.3005
R1642 VTAIL.n216 VTAIL.n215 9.3005
R1643 VTAIL.n218 VTAIL.n217 9.3005
R1644 VTAIL.n233 VTAIL.n232 9.3005
R1645 VTAIL.n180 VTAIL.n179 9.3005
R1646 VTAIL.n227 VTAIL.n226 9.3005
R1647 VTAIL.n225 VTAIL.n224 9.3005
R1648 VTAIL.n184 VTAIL.n183 9.3005
R1649 VTAIL.n438 VTAIL.n428 8.92171
R1650 VTAIL.n26 VTAIL.n16 8.92171
R1651 VTAIL.n84 VTAIL.n74 8.92171
R1652 VTAIL.n144 VTAIL.n134 8.92171
R1653 VTAIL.n381 VTAIL.n371 8.92171
R1654 VTAIL.n321 VTAIL.n311 8.92171
R1655 VTAIL.n263 VTAIL.n253 8.92171
R1656 VTAIL.n203 VTAIL.n193 8.92171
R1657 VTAIL.n437 VTAIL.n430 8.14595
R1658 VTAIL.n25 VTAIL.n18 8.14595
R1659 VTAIL.n83 VTAIL.n76 8.14595
R1660 VTAIL.n143 VTAIL.n136 8.14595
R1661 VTAIL.n380 VTAIL.n373 8.14595
R1662 VTAIL.n320 VTAIL.n313 8.14595
R1663 VTAIL.n262 VTAIL.n255 8.14595
R1664 VTAIL.n202 VTAIL.n195 8.14595
R1665 VTAIL.n434 VTAIL.n433 7.3702
R1666 VTAIL.n22 VTAIL.n21 7.3702
R1667 VTAIL.n80 VTAIL.n79 7.3702
R1668 VTAIL.n140 VTAIL.n139 7.3702
R1669 VTAIL.n377 VTAIL.n376 7.3702
R1670 VTAIL.n317 VTAIL.n316 7.3702
R1671 VTAIL.n259 VTAIL.n258 7.3702
R1672 VTAIL.n199 VTAIL.n198 7.3702
R1673 VTAIL.n434 VTAIL.n430 5.81868
R1674 VTAIL.n22 VTAIL.n18 5.81868
R1675 VTAIL.n80 VTAIL.n76 5.81868
R1676 VTAIL.n140 VTAIL.n136 5.81868
R1677 VTAIL.n377 VTAIL.n373 5.81868
R1678 VTAIL.n317 VTAIL.n313 5.81868
R1679 VTAIL.n259 VTAIL.n255 5.81868
R1680 VTAIL.n199 VTAIL.n195 5.81868
R1681 VTAIL.n438 VTAIL.n437 5.04292
R1682 VTAIL.n26 VTAIL.n25 5.04292
R1683 VTAIL.n84 VTAIL.n83 5.04292
R1684 VTAIL.n144 VTAIL.n143 5.04292
R1685 VTAIL.n381 VTAIL.n380 5.04292
R1686 VTAIL.n321 VTAIL.n320 5.04292
R1687 VTAIL.n263 VTAIL.n262 5.04292
R1688 VTAIL.n203 VTAIL.n202 5.04292
R1689 VTAIL.n441 VTAIL.n428 4.26717
R1690 VTAIL.n470 VTAIL.n414 4.26717
R1691 VTAIL.n29 VTAIL.n16 4.26717
R1692 VTAIL.n58 VTAIL.n2 4.26717
R1693 VTAIL.n87 VTAIL.n74 4.26717
R1694 VTAIL.n116 VTAIL.n60 4.26717
R1695 VTAIL.n147 VTAIL.n134 4.26717
R1696 VTAIL.n176 VTAIL.n120 4.26717
R1697 VTAIL.n412 VTAIL.n356 4.26717
R1698 VTAIL.n384 VTAIL.n371 4.26717
R1699 VTAIL.n352 VTAIL.n296 4.26717
R1700 VTAIL.n324 VTAIL.n311 4.26717
R1701 VTAIL.n294 VTAIL.n238 4.26717
R1702 VTAIL.n266 VTAIL.n253 4.26717
R1703 VTAIL.n234 VTAIL.n178 4.26717
R1704 VTAIL.n206 VTAIL.n193 4.26717
R1705 VTAIL.n442 VTAIL.n426 3.49141
R1706 VTAIL.n468 VTAIL.n467 3.49141
R1707 VTAIL.n30 VTAIL.n14 3.49141
R1708 VTAIL.n56 VTAIL.n55 3.49141
R1709 VTAIL.n88 VTAIL.n72 3.49141
R1710 VTAIL.n114 VTAIL.n113 3.49141
R1711 VTAIL.n148 VTAIL.n132 3.49141
R1712 VTAIL.n174 VTAIL.n173 3.49141
R1713 VTAIL.n410 VTAIL.n409 3.49141
R1714 VTAIL.n385 VTAIL.n369 3.49141
R1715 VTAIL.n350 VTAIL.n349 3.49141
R1716 VTAIL.n325 VTAIL.n309 3.49141
R1717 VTAIL.n292 VTAIL.n291 3.49141
R1718 VTAIL.n267 VTAIL.n251 3.49141
R1719 VTAIL.n232 VTAIL.n231 3.49141
R1720 VTAIL.n207 VTAIL.n191 3.49141
R1721 VTAIL.n435 VTAIL.n431 2.84303
R1722 VTAIL.n23 VTAIL.n19 2.84303
R1723 VTAIL.n81 VTAIL.n77 2.84303
R1724 VTAIL.n141 VTAIL.n137 2.84303
R1725 VTAIL.n378 VTAIL.n374 2.84303
R1726 VTAIL.n318 VTAIL.n314 2.84303
R1727 VTAIL.n260 VTAIL.n256 2.84303
R1728 VTAIL.n200 VTAIL.n196 2.84303
R1729 VTAIL.n446 VTAIL.n445 2.71565
R1730 VTAIL.n464 VTAIL.n416 2.71565
R1731 VTAIL.n34 VTAIL.n33 2.71565
R1732 VTAIL.n52 VTAIL.n4 2.71565
R1733 VTAIL.n92 VTAIL.n91 2.71565
R1734 VTAIL.n110 VTAIL.n62 2.71565
R1735 VTAIL.n152 VTAIL.n151 2.71565
R1736 VTAIL.n170 VTAIL.n122 2.71565
R1737 VTAIL.n406 VTAIL.n358 2.71565
R1738 VTAIL.n389 VTAIL.n388 2.71565
R1739 VTAIL.n346 VTAIL.n298 2.71565
R1740 VTAIL.n329 VTAIL.n328 2.71565
R1741 VTAIL.n288 VTAIL.n240 2.71565
R1742 VTAIL.n271 VTAIL.n270 2.71565
R1743 VTAIL.n228 VTAIL.n180 2.71565
R1744 VTAIL.n211 VTAIL.n210 2.71565
R1745 VTAIL.n450 VTAIL.n424 1.93989
R1746 VTAIL.n463 VTAIL.n418 1.93989
R1747 VTAIL.n38 VTAIL.n12 1.93989
R1748 VTAIL.n51 VTAIL.n6 1.93989
R1749 VTAIL.n96 VTAIL.n70 1.93989
R1750 VTAIL.n109 VTAIL.n64 1.93989
R1751 VTAIL.n156 VTAIL.n130 1.93989
R1752 VTAIL.n169 VTAIL.n124 1.93989
R1753 VTAIL.n405 VTAIL.n360 1.93989
R1754 VTAIL.n392 VTAIL.n366 1.93989
R1755 VTAIL.n345 VTAIL.n300 1.93989
R1756 VTAIL.n332 VTAIL.n306 1.93989
R1757 VTAIL.n287 VTAIL.n242 1.93989
R1758 VTAIL.n274 VTAIL.n248 1.93989
R1759 VTAIL.n227 VTAIL.n182 1.93989
R1760 VTAIL.n214 VTAIL.n188 1.93989
R1761 VTAIL.n0 VTAIL.t6 1.87373
R1762 VTAIL.n0 VTAIL.t1 1.87373
R1763 VTAIL.n118 VTAIL.t10 1.87373
R1764 VTAIL.n118 VTAIL.t8 1.87373
R1765 VTAIL.n354 VTAIL.t11 1.87373
R1766 VTAIL.n354 VTAIL.t15 1.87373
R1767 VTAIL.n236 VTAIL.t3 1.87373
R1768 VTAIL.n236 VTAIL.t7 1.87373
R1769 VTAIL.n451 VTAIL.n422 1.16414
R1770 VTAIL.n460 VTAIL.n459 1.16414
R1771 VTAIL.n39 VTAIL.n10 1.16414
R1772 VTAIL.n48 VTAIL.n47 1.16414
R1773 VTAIL.n97 VTAIL.n68 1.16414
R1774 VTAIL.n106 VTAIL.n105 1.16414
R1775 VTAIL.n157 VTAIL.n128 1.16414
R1776 VTAIL.n166 VTAIL.n165 1.16414
R1777 VTAIL.n402 VTAIL.n401 1.16414
R1778 VTAIL.n393 VTAIL.n364 1.16414
R1779 VTAIL.n342 VTAIL.n341 1.16414
R1780 VTAIL.n333 VTAIL.n304 1.16414
R1781 VTAIL.n284 VTAIL.n283 1.16414
R1782 VTAIL.n275 VTAIL.n246 1.16414
R1783 VTAIL.n224 VTAIL.n223 1.16414
R1784 VTAIL.n215 VTAIL.n186 1.16414
R1785 VTAIL.n237 VTAIL.n235 0.888431
R1786 VTAIL.n295 VTAIL.n237 0.888431
R1787 VTAIL.n355 VTAIL.n353 0.888431
R1788 VTAIL.n413 VTAIL.n355 0.888431
R1789 VTAIL.n177 VTAIL.n119 0.888431
R1790 VTAIL.n119 VTAIL.n117 0.888431
R1791 VTAIL.n59 VTAIL.n1 0.888431
R1792 VTAIL VTAIL.n471 0.830241
R1793 VTAIL.n353 VTAIL.n295 0.470328
R1794 VTAIL.n117 VTAIL.n59 0.470328
R1795 VTAIL.n455 VTAIL.n454 0.388379
R1796 VTAIL.n456 VTAIL.n420 0.388379
R1797 VTAIL.n43 VTAIL.n42 0.388379
R1798 VTAIL.n44 VTAIL.n8 0.388379
R1799 VTAIL.n101 VTAIL.n100 0.388379
R1800 VTAIL.n102 VTAIL.n66 0.388379
R1801 VTAIL.n161 VTAIL.n160 0.388379
R1802 VTAIL.n162 VTAIL.n126 0.388379
R1803 VTAIL.n398 VTAIL.n362 0.388379
R1804 VTAIL.n397 VTAIL.n396 0.388379
R1805 VTAIL.n338 VTAIL.n302 0.388379
R1806 VTAIL.n337 VTAIL.n336 0.388379
R1807 VTAIL.n280 VTAIL.n244 0.388379
R1808 VTAIL.n279 VTAIL.n278 0.388379
R1809 VTAIL.n220 VTAIL.n184 0.388379
R1810 VTAIL.n219 VTAIL.n218 0.388379
R1811 VTAIL.n436 VTAIL.n435 0.155672
R1812 VTAIL.n436 VTAIL.n427 0.155672
R1813 VTAIL.n443 VTAIL.n427 0.155672
R1814 VTAIL.n444 VTAIL.n443 0.155672
R1815 VTAIL.n444 VTAIL.n423 0.155672
R1816 VTAIL.n452 VTAIL.n423 0.155672
R1817 VTAIL.n453 VTAIL.n452 0.155672
R1818 VTAIL.n453 VTAIL.n419 0.155672
R1819 VTAIL.n461 VTAIL.n419 0.155672
R1820 VTAIL.n462 VTAIL.n461 0.155672
R1821 VTAIL.n462 VTAIL.n415 0.155672
R1822 VTAIL.n469 VTAIL.n415 0.155672
R1823 VTAIL.n24 VTAIL.n23 0.155672
R1824 VTAIL.n24 VTAIL.n15 0.155672
R1825 VTAIL.n31 VTAIL.n15 0.155672
R1826 VTAIL.n32 VTAIL.n31 0.155672
R1827 VTAIL.n32 VTAIL.n11 0.155672
R1828 VTAIL.n40 VTAIL.n11 0.155672
R1829 VTAIL.n41 VTAIL.n40 0.155672
R1830 VTAIL.n41 VTAIL.n7 0.155672
R1831 VTAIL.n49 VTAIL.n7 0.155672
R1832 VTAIL.n50 VTAIL.n49 0.155672
R1833 VTAIL.n50 VTAIL.n3 0.155672
R1834 VTAIL.n57 VTAIL.n3 0.155672
R1835 VTAIL.n82 VTAIL.n81 0.155672
R1836 VTAIL.n82 VTAIL.n73 0.155672
R1837 VTAIL.n89 VTAIL.n73 0.155672
R1838 VTAIL.n90 VTAIL.n89 0.155672
R1839 VTAIL.n90 VTAIL.n69 0.155672
R1840 VTAIL.n98 VTAIL.n69 0.155672
R1841 VTAIL.n99 VTAIL.n98 0.155672
R1842 VTAIL.n99 VTAIL.n65 0.155672
R1843 VTAIL.n107 VTAIL.n65 0.155672
R1844 VTAIL.n108 VTAIL.n107 0.155672
R1845 VTAIL.n108 VTAIL.n61 0.155672
R1846 VTAIL.n115 VTAIL.n61 0.155672
R1847 VTAIL.n142 VTAIL.n141 0.155672
R1848 VTAIL.n142 VTAIL.n133 0.155672
R1849 VTAIL.n149 VTAIL.n133 0.155672
R1850 VTAIL.n150 VTAIL.n149 0.155672
R1851 VTAIL.n150 VTAIL.n129 0.155672
R1852 VTAIL.n158 VTAIL.n129 0.155672
R1853 VTAIL.n159 VTAIL.n158 0.155672
R1854 VTAIL.n159 VTAIL.n125 0.155672
R1855 VTAIL.n167 VTAIL.n125 0.155672
R1856 VTAIL.n168 VTAIL.n167 0.155672
R1857 VTAIL.n168 VTAIL.n121 0.155672
R1858 VTAIL.n175 VTAIL.n121 0.155672
R1859 VTAIL.n411 VTAIL.n357 0.155672
R1860 VTAIL.n404 VTAIL.n357 0.155672
R1861 VTAIL.n404 VTAIL.n403 0.155672
R1862 VTAIL.n403 VTAIL.n361 0.155672
R1863 VTAIL.n395 VTAIL.n361 0.155672
R1864 VTAIL.n395 VTAIL.n394 0.155672
R1865 VTAIL.n394 VTAIL.n365 0.155672
R1866 VTAIL.n387 VTAIL.n365 0.155672
R1867 VTAIL.n387 VTAIL.n386 0.155672
R1868 VTAIL.n386 VTAIL.n370 0.155672
R1869 VTAIL.n379 VTAIL.n370 0.155672
R1870 VTAIL.n379 VTAIL.n378 0.155672
R1871 VTAIL.n351 VTAIL.n297 0.155672
R1872 VTAIL.n344 VTAIL.n297 0.155672
R1873 VTAIL.n344 VTAIL.n343 0.155672
R1874 VTAIL.n343 VTAIL.n301 0.155672
R1875 VTAIL.n335 VTAIL.n301 0.155672
R1876 VTAIL.n335 VTAIL.n334 0.155672
R1877 VTAIL.n334 VTAIL.n305 0.155672
R1878 VTAIL.n327 VTAIL.n305 0.155672
R1879 VTAIL.n327 VTAIL.n326 0.155672
R1880 VTAIL.n326 VTAIL.n310 0.155672
R1881 VTAIL.n319 VTAIL.n310 0.155672
R1882 VTAIL.n319 VTAIL.n318 0.155672
R1883 VTAIL.n293 VTAIL.n239 0.155672
R1884 VTAIL.n286 VTAIL.n239 0.155672
R1885 VTAIL.n286 VTAIL.n285 0.155672
R1886 VTAIL.n285 VTAIL.n243 0.155672
R1887 VTAIL.n277 VTAIL.n243 0.155672
R1888 VTAIL.n277 VTAIL.n276 0.155672
R1889 VTAIL.n276 VTAIL.n247 0.155672
R1890 VTAIL.n269 VTAIL.n247 0.155672
R1891 VTAIL.n269 VTAIL.n268 0.155672
R1892 VTAIL.n268 VTAIL.n252 0.155672
R1893 VTAIL.n261 VTAIL.n252 0.155672
R1894 VTAIL.n261 VTAIL.n260 0.155672
R1895 VTAIL.n233 VTAIL.n179 0.155672
R1896 VTAIL.n226 VTAIL.n179 0.155672
R1897 VTAIL.n226 VTAIL.n225 0.155672
R1898 VTAIL.n225 VTAIL.n183 0.155672
R1899 VTAIL.n217 VTAIL.n183 0.155672
R1900 VTAIL.n217 VTAIL.n216 0.155672
R1901 VTAIL.n216 VTAIL.n187 0.155672
R1902 VTAIL.n209 VTAIL.n187 0.155672
R1903 VTAIL.n209 VTAIL.n208 0.155672
R1904 VTAIL.n208 VTAIL.n192 0.155672
R1905 VTAIL.n201 VTAIL.n192 0.155672
R1906 VTAIL.n201 VTAIL.n200 0.155672
R1907 VTAIL VTAIL.n1 0.0586897
R1908 VN.n3 VN.t2 442.551
R1909 VN.n13 VN.t4 442.551
R1910 VN.n2 VN.t1 420.373
R1911 VN.n6 VN.t5 420.373
R1912 VN.n8 VN.t7 420.373
R1913 VN.n12 VN.t0 420.373
R1914 VN.n16 VN.t3 420.373
R1915 VN.n18 VN.t6 420.373
R1916 VN.n9 VN.n8 161.3
R1917 VN.n19 VN.n18 161.3
R1918 VN.n17 VN.n10 161.3
R1919 VN.n16 VN.n15 161.3
R1920 VN.n14 VN.n11 161.3
R1921 VN.n7 VN.n0 161.3
R1922 VN.n6 VN.n5 161.3
R1923 VN.n4 VN.n1 161.3
R1924 VN.n14 VN.n13 44.862
R1925 VN.n4 VN.n3 44.862
R1926 VN VN.n19 41.2903
R1927 VN.n8 VN.n7 28.4823
R1928 VN.n18 VN.n17 28.4823
R1929 VN.n2 VN.n1 24.1005
R1930 VN.n6 VN.n1 24.1005
R1931 VN.n16 VN.n11 24.1005
R1932 VN.n12 VN.n11 24.1005
R1933 VN.n7 VN.n6 19.7187
R1934 VN.n17 VN.n16 19.7187
R1935 VN.n3 VN.n2 19.7081
R1936 VN.n13 VN.n12 19.7081
R1937 VN.n19 VN.n10 0.189894
R1938 VN.n15 VN.n10 0.189894
R1939 VN.n15 VN.n14 0.189894
R1940 VN.n5 VN.n4 0.189894
R1941 VN.n5 VN.n0 0.189894
R1942 VN.n9 VN.n0 0.189894
R1943 VN VN.n9 0.0516364
R1944 VDD2.n2 VDD2.n1 60.5954
R1945 VDD2.n2 VDD2.n0 60.5954
R1946 VDD2 VDD2.n5 60.5926
R1947 VDD2.n4 VDD2.n3 60.207
R1948 VDD2.n4 VDD2.n2 36.8231
R1949 VDD2.n5 VDD2.t7 1.87373
R1950 VDD2.n5 VDD2.t3 1.87373
R1951 VDD2.n3 VDD2.t1 1.87373
R1952 VDD2.n3 VDD2.t4 1.87373
R1953 VDD2.n1 VDD2.t2 1.87373
R1954 VDD2.n1 VDD2.t0 1.87373
R1955 VDD2.n0 VDD2.t5 1.87373
R1956 VDD2.n0 VDD2.t6 1.87373
R1957 VDD2 VDD2.n4 0.502655
C0 VN VDD1 0.147841f
C1 VTAIL VDD1 10.0115f
C2 VDD2 VP 0.317038f
C3 VN VDD2 4.904819f
C4 VTAIL VDD2 10.0531f
C5 VN VP 5.07523f
C6 VTAIL VP 4.72612f
C7 VDD1 VDD2 0.823064f
C8 VN VTAIL 4.712009f
C9 VDD1 VP 5.07358f
C10 VDD2 B 3.378607f
C11 VDD1 B 3.612516f
C12 VTAIL B 8.122186f
C13 VN B 8.419741f
C14 VP B 6.540079f
C15 VDD2.t5 B 0.228512f
C16 VDD2.t6 B 0.228512f
C17 VDD2.n0 B 2.01953f
C18 VDD2.t2 B 0.228512f
C19 VDD2.t0 B 0.228512f
C20 VDD2.n1 B 2.01953f
C21 VDD2.n2 B 2.28433f
C22 VDD2.t1 B 0.228512f
C23 VDD2.t4 B 0.228512f
C24 VDD2.n3 B 2.01728f
C25 VDD2.n4 B 2.38571f
C26 VDD2.t7 B 0.228512f
C27 VDD2.t3 B 0.228512f
C28 VDD2.n5 B 2.0195f
C29 VN.n0 B 0.044151f
C30 VN.n1 B 0.010019f
C31 VN.t2 B 0.95303f
C32 VN.t1 B 0.93396f
C33 VN.n2 B 0.38476f
C34 VN.n3 B 0.365757f
C35 VN.n4 B 0.183599f
C36 VN.n5 B 0.044151f
C37 VN.t5 B 0.93396f
C38 VN.n6 B 0.380765f
C39 VN.n7 B 0.010019f
C40 VN.t7 B 0.93396f
C41 VN.n8 B 0.377907f
C42 VN.n9 B 0.034215f
C43 VN.n10 B 0.044151f
C44 VN.n11 B 0.010019f
C45 VN.t3 B 0.93396f
C46 VN.t4 B 0.95303f
C47 VN.t0 B 0.93396f
C48 VN.n12 B 0.38476f
C49 VN.n13 B 0.365757f
C50 VN.n14 B 0.183599f
C51 VN.n15 B 0.044151f
C52 VN.n16 B 0.380765f
C53 VN.n17 B 0.010019f
C54 VN.t6 B 0.93396f
C55 VN.n18 B 0.377907f
C56 VN.n19 B 1.77257f
C57 VTAIL.t6 B 0.169692f
C58 VTAIL.t1 B 0.169692f
C59 VTAIL.n0 B 1.435f
C60 VTAIL.n1 B 0.265662f
C61 VTAIL.n2 B 0.025951f
C62 VTAIL.n3 B 0.020316f
C63 VTAIL.n4 B 0.010917f
C64 VTAIL.n5 B 0.025803f
C65 VTAIL.n6 B 0.011559f
C66 VTAIL.n7 B 0.020316f
C67 VTAIL.n8 B 0.010917f
C68 VTAIL.n9 B 0.025803f
C69 VTAIL.n10 B 0.011559f
C70 VTAIL.n11 B 0.020316f
C71 VTAIL.n12 B 0.010917f
C72 VTAIL.n13 B 0.025803f
C73 VTAIL.n14 B 0.011559f
C74 VTAIL.n15 B 0.020316f
C75 VTAIL.n16 B 0.010917f
C76 VTAIL.n17 B 0.025803f
C77 VTAIL.n18 B 0.011559f
C78 VTAIL.n19 B 0.135322f
C79 VTAIL.t5 B 0.043424f
C80 VTAIL.n20 B 0.019353f
C81 VTAIL.n21 B 0.018241f
C82 VTAIL.n22 B 0.010917f
C83 VTAIL.n23 B 0.895676f
C84 VTAIL.n24 B 0.020316f
C85 VTAIL.n25 B 0.010917f
C86 VTAIL.n26 B 0.011559f
C87 VTAIL.n27 B 0.025803f
C88 VTAIL.n28 B 0.025803f
C89 VTAIL.n29 B 0.011559f
C90 VTAIL.n30 B 0.010917f
C91 VTAIL.n31 B 0.020316f
C92 VTAIL.n32 B 0.020316f
C93 VTAIL.n33 B 0.010917f
C94 VTAIL.n34 B 0.011559f
C95 VTAIL.n35 B 0.025803f
C96 VTAIL.n36 B 0.025803f
C97 VTAIL.n37 B 0.025803f
C98 VTAIL.n38 B 0.011559f
C99 VTAIL.n39 B 0.010917f
C100 VTAIL.n40 B 0.020316f
C101 VTAIL.n41 B 0.020316f
C102 VTAIL.n42 B 0.010917f
C103 VTAIL.n43 B 0.011238f
C104 VTAIL.n44 B 0.011238f
C105 VTAIL.n45 B 0.025803f
C106 VTAIL.n46 B 0.025803f
C107 VTAIL.n47 B 0.011559f
C108 VTAIL.n48 B 0.010917f
C109 VTAIL.n49 B 0.020316f
C110 VTAIL.n50 B 0.020316f
C111 VTAIL.n51 B 0.010917f
C112 VTAIL.n52 B 0.011559f
C113 VTAIL.n53 B 0.025803f
C114 VTAIL.n54 B 0.051255f
C115 VTAIL.n55 B 0.011559f
C116 VTAIL.n56 B 0.010917f
C117 VTAIL.n57 B 0.043906f
C118 VTAIL.n58 B 0.028109f
C119 VTAIL.n59 B 0.104513f
C120 VTAIL.n60 B 0.025951f
C121 VTAIL.n61 B 0.020316f
C122 VTAIL.n62 B 0.010917f
C123 VTAIL.n63 B 0.025803f
C124 VTAIL.n64 B 0.011559f
C125 VTAIL.n65 B 0.020316f
C126 VTAIL.n66 B 0.010917f
C127 VTAIL.n67 B 0.025803f
C128 VTAIL.n68 B 0.011559f
C129 VTAIL.n69 B 0.020316f
C130 VTAIL.n70 B 0.010917f
C131 VTAIL.n71 B 0.025803f
C132 VTAIL.n72 B 0.011559f
C133 VTAIL.n73 B 0.020316f
C134 VTAIL.n74 B 0.010917f
C135 VTAIL.n75 B 0.025803f
C136 VTAIL.n76 B 0.011559f
C137 VTAIL.n77 B 0.135322f
C138 VTAIL.t9 B 0.043424f
C139 VTAIL.n78 B 0.019353f
C140 VTAIL.n79 B 0.018241f
C141 VTAIL.n80 B 0.010917f
C142 VTAIL.n81 B 0.895676f
C143 VTAIL.n82 B 0.020316f
C144 VTAIL.n83 B 0.010917f
C145 VTAIL.n84 B 0.011559f
C146 VTAIL.n85 B 0.025803f
C147 VTAIL.n86 B 0.025803f
C148 VTAIL.n87 B 0.011559f
C149 VTAIL.n88 B 0.010917f
C150 VTAIL.n89 B 0.020316f
C151 VTAIL.n90 B 0.020316f
C152 VTAIL.n91 B 0.010917f
C153 VTAIL.n92 B 0.011559f
C154 VTAIL.n93 B 0.025803f
C155 VTAIL.n94 B 0.025803f
C156 VTAIL.n95 B 0.025803f
C157 VTAIL.n96 B 0.011559f
C158 VTAIL.n97 B 0.010917f
C159 VTAIL.n98 B 0.020316f
C160 VTAIL.n99 B 0.020316f
C161 VTAIL.n100 B 0.010917f
C162 VTAIL.n101 B 0.011238f
C163 VTAIL.n102 B 0.011238f
C164 VTAIL.n103 B 0.025803f
C165 VTAIL.n104 B 0.025803f
C166 VTAIL.n105 B 0.011559f
C167 VTAIL.n106 B 0.010917f
C168 VTAIL.n107 B 0.020316f
C169 VTAIL.n108 B 0.020316f
C170 VTAIL.n109 B 0.010917f
C171 VTAIL.n110 B 0.011559f
C172 VTAIL.n111 B 0.025803f
C173 VTAIL.n112 B 0.051255f
C174 VTAIL.n113 B 0.011559f
C175 VTAIL.n114 B 0.010917f
C176 VTAIL.n115 B 0.043906f
C177 VTAIL.n116 B 0.028109f
C178 VTAIL.n117 B 0.104513f
C179 VTAIL.t10 B 0.169692f
C180 VTAIL.t8 B 0.169692f
C181 VTAIL.n118 B 1.435f
C182 VTAIL.n119 B 0.319979f
C183 VTAIL.n120 B 0.025951f
C184 VTAIL.n121 B 0.020316f
C185 VTAIL.n122 B 0.010917f
C186 VTAIL.n123 B 0.025803f
C187 VTAIL.n124 B 0.011559f
C188 VTAIL.n125 B 0.020316f
C189 VTAIL.n126 B 0.010917f
C190 VTAIL.n127 B 0.025803f
C191 VTAIL.n128 B 0.011559f
C192 VTAIL.n129 B 0.020316f
C193 VTAIL.n130 B 0.010917f
C194 VTAIL.n131 B 0.025803f
C195 VTAIL.n132 B 0.011559f
C196 VTAIL.n133 B 0.020316f
C197 VTAIL.n134 B 0.010917f
C198 VTAIL.n135 B 0.025803f
C199 VTAIL.n136 B 0.011559f
C200 VTAIL.n137 B 0.135322f
C201 VTAIL.t13 B 0.043424f
C202 VTAIL.n138 B 0.019353f
C203 VTAIL.n139 B 0.018241f
C204 VTAIL.n140 B 0.010917f
C205 VTAIL.n141 B 0.895676f
C206 VTAIL.n142 B 0.020316f
C207 VTAIL.n143 B 0.010917f
C208 VTAIL.n144 B 0.011559f
C209 VTAIL.n145 B 0.025803f
C210 VTAIL.n146 B 0.025803f
C211 VTAIL.n147 B 0.011559f
C212 VTAIL.n148 B 0.010917f
C213 VTAIL.n149 B 0.020316f
C214 VTAIL.n150 B 0.020316f
C215 VTAIL.n151 B 0.010917f
C216 VTAIL.n152 B 0.011559f
C217 VTAIL.n153 B 0.025803f
C218 VTAIL.n154 B 0.025803f
C219 VTAIL.n155 B 0.025803f
C220 VTAIL.n156 B 0.011559f
C221 VTAIL.n157 B 0.010917f
C222 VTAIL.n158 B 0.020316f
C223 VTAIL.n159 B 0.020316f
C224 VTAIL.n160 B 0.010917f
C225 VTAIL.n161 B 0.011238f
C226 VTAIL.n162 B 0.011238f
C227 VTAIL.n163 B 0.025803f
C228 VTAIL.n164 B 0.025803f
C229 VTAIL.n165 B 0.011559f
C230 VTAIL.n166 B 0.010917f
C231 VTAIL.n167 B 0.020316f
C232 VTAIL.n168 B 0.020316f
C233 VTAIL.n169 B 0.010917f
C234 VTAIL.n170 B 0.011559f
C235 VTAIL.n171 B 0.025803f
C236 VTAIL.n172 B 0.051255f
C237 VTAIL.n173 B 0.011559f
C238 VTAIL.n174 B 0.010917f
C239 VTAIL.n175 B 0.043906f
C240 VTAIL.n176 B 0.028109f
C241 VTAIL.n177 B 1.00434f
C242 VTAIL.n178 B 0.025951f
C243 VTAIL.n179 B 0.020316f
C244 VTAIL.n180 B 0.010917f
C245 VTAIL.n181 B 0.025803f
C246 VTAIL.n182 B 0.011559f
C247 VTAIL.n183 B 0.020316f
C248 VTAIL.n184 B 0.010917f
C249 VTAIL.n185 B 0.025803f
C250 VTAIL.n186 B 0.011559f
C251 VTAIL.n187 B 0.020316f
C252 VTAIL.n188 B 0.010917f
C253 VTAIL.n189 B 0.025803f
C254 VTAIL.n190 B 0.025803f
C255 VTAIL.n191 B 0.011559f
C256 VTAIL.n192 B 0.020316f
C257 VTAIL.n193 B 0.010917f
C258 VTAIL.n194 B 0.025803f
C259 VTAIL.n195 B 0.011559f
C260 VTAIL.n196 B 0.135322f
C261 VTAIL.t2 B 0.043424f
C262 VTAIL.n197 B 0.019353f
C263 VTAIL.n198 B 0.018241f
C264 VTAIL.n199 B 0.010917f
C265 VTAIL.n200 B 0.895676f
C266 VTAIL.n201 B 0.020316f
C267 VTAIL.n202 B 0.010917f
C268 VTAIL.n203 B 0.011559f
C269 VTAIL.n204 B 0.025803f
C270 VTAIL.n205 B 0.025803f
C271 VTAIL.n206 B 0.011559f
C272 VTAIL.n207 B 0.010917f
C273 VTAIL.n208 B 0.020316f
C274 VTAIL.n209 B 0.020316f
C275 VTAIL.n210 B 0.010917f
C276 VTAIL.n211 B 0.011559f
C277 VTAIL.n212 B 0.025803f
C278 VTAIL.n213 B 0.025803f
C279 VTAIL.n214 B 0.011559f
C280 VTAIL.n215 B 0.010917f
C281 VTAIL.n216 B 0.020316f
C282 VTAIL.n217 B 0.020316f
C283 VTAIL.n218 B 0.010917f
C284 VTAIL.n219 B 0.011238f
C285 VTAIL.n220 B 0.011238f
C286 VTAIL.n221 B 0.025803f
C287 VTAIL.n222 B 0.025803f
C288 VTAIL.n223 B 0.011559f
C289 VTAIL.n224 B 0.010917f
C290 VTAIL.n225 B 0.020316f
C291 VTAIL.n226 B 0.020316f
C292 VTAIL.n227 B 0.010917f
C293 VTAIL.n228 B 0.011559f
C294 VTAIL.n229 B 0.025803f
C295 VTAIL.n230 B 0.051255f
C296 VTAIL.n231 B 0.011559f
C297 VTAIL.n232 B 0.010917f
C298 VTAIL.n233 B 0.043906f
C299 VTAIL.n234 B 0.028109f
C300 VTAIL.n235 B 1.00434f
C301 VTAIL.t3 B 0.169692f
C302 VTAIL.t7 B 0.169692f
C303 VTAIL.n236 B 1.43501f
C304 VTAIL.n237 B 0.31997f
C305 VTAIL.n238 B 0.025951f
C306 VTAIL.n239 B 0.020316f
C307 VTAIL.n240 B 0.010917f
C308 VTAIL.n241 B 0.025803f
C309 VTAIL.n242 B 0.011559f
C310 VTAIL.n243 B 0.020316f
C311 VTAIL.n244 B 0.010917f
C312 VTAIL.n245 B 0.025803f
C313 VTAIL.n246 B 0.011559f
C314 VTAIL.n247 B 0.020316f
C315 VTAIL.n248 B 0.010917f
C316 VTAIL.n249 B 0.025803f
C317 VTAIL.n250 B 0.025803f
C318 VTAIL.n251 B 0.011559f
C319 VTAIL.n252 B 0.020316f
C320 VTAIL.n253 B 0.010917f
C321 VTAIL.n254 B 0.025803f
C322 VTAIL.n255 B 0.011559f
C323 VTAIL.n256 B 0.135322f
C324 VTAIL.t4 B 0.043424f
C325 VTAIL.n257 B 0.019353f
C326 VTAIL.n258 B 0.018241f
C327 VTAIL.n259 B 0.010917f
C328 VTAIL.n260 B 0.895676f
C329 VTAIL.n261 B 0.020316f
C330 VTAIL.n262 B 0.010917f
C331 VTAIL.n263 B 0.011559f
C332 VTAIL.n264 B 0.025803f
C333 VTAIL.n265 B 0.025803f
C334 VTAIL.n266 B 0.011559f
C335 VTAIL.n267 B 0.010917f
C336 VTAIL.n268 B 0.020316f
C337 VTAIL.n269 B 0.020316f
C338 VTAIL.n270 B 0.010917f
C339 VTAIL.n271 B 0.011559f
C340 VTAIL.n272 B 0.025803f
C341 VTAIL.n273 B 0.025803f
C342 VTAIL.n274 B 0.011559f
C343 VTAIL.n275 B 0.010917f
C344 VTAIL.n276 B 0.020316f
C345 VTAIL.n277 B 0.020316f
C346 VTAIL.n278 B 0.010917f
C347 VTAIL.n279 B 0.011238f
C348 VTAIL.n280 B 0.011238f
C349 VTAIL.n281 B 0.025803f
C350 VTAIL.n282 B 0.025803f
C351 VTAIL.n283 B 0.011559f
C352 VTAIL.n284 B 0.010917f
C353 VTAIL.n285 B 0.020316f
C354 VTAIL.n286 B 0.020316f
C355 VTAIL.n287 B 0.010917f
C356 VTAIL.n288 B 0.011559f
C357 VTAIL.n289 B 0.025803f
C358 VTAIL.n290 B 0.051255f
C359 VTAIL.n291 B 0.011559f
C360 VTAIL.n292 B 0.010917f
C361 VTAIL.n293 B 0.043906f
C362 VTAIL.n294 B 0.028109f
C363 VTAIL.n295 B 0.104513f
C364 VTAIL.n296 B 0.025951f
C365 VTAIL.n297 B 0.020316f
C366 VTAIL.n298 B 0.010917f
C367 VTAIL.n299 B 0.025803f
C368 VTAIL.n300 B 0.011559f
C369 VTAIL.n301 B 0.020316f
C370 VTAIL.n302 B 0.010917f
C371 VTAIL.n303 B 0.025803f
C372 VTAIL.n304 B 0.011559f
C373 VTAIL.n305 B 0.020316f
C374 VTAIL.n306 B 0.010917f
C375 VTAIL.n307 B 0.025803f
C376 VTAIL.n308 B 0.025803f
C377 VTAIL.n309 B 0.011559f
C378 VTAIL.n310 B 0.020316f
C379 VTAIL.n311 B 0.010917f
C380 VTAIL.n312 B 0.025803f
C381 VTAIL.n313 B 0.011559f
C382 VTAIL.n314 B 0.135322f
C383 VTAIL.t14 B 0.043424f
C384 VTAIL.n315 B 0.019353f
C385 VTAIL.n316 B 0.018241f
C386 VTAIL.n317 B 0.010917f
C387 VTAIL.n318 B 0.895676f
C388 VTAIL.n319 B 0.020316f
C389 VTAIL.n320 B 0.010917f
C390 VTAIL.n321 B 0.011559f
C391 VTAIL.n322 B 0.025803f
C392 VTAIL.n323 B 0.025803f
C393 VTAIL.n324 B 0.011559f
C394 VTAIL.n325 B 0.010917f
C395 VTAIL.n326 B 0.020316f
C396 VTAIL.n327 B 0.020316f
C397 VTAIL.n328 B 0.010917f
C398 VTAIL.n329 B 0.011559f
C399 VTAIL.n330 B 0.025803f
C400 VTAIL.n331 B 0.025803f
C401 VTAIL.n332 B 0.011559f
C402 VTAIL.n333 B 0.010917f
C403 VTAIL.n334 B 0.020316f
C404 VTAIL.n335 B 0.020316f
C405 VTAIL.n336 B 0.010917f
C406 VTAIL.n337 B 0.011238f
C407 VTAIL.n338 B 0.011238f
C408 VTAIL.n339 B 0.025803f
C409 VTAIL.n340 B 0.025803f
C410 VTAIL.n341 B 0.011559f
C411 VTAIL.n342 B 0.010917f
C412 VTAIL.n343 B 0.020316f
C413 VTAIL.n344 B 0.020316f
C414 VTAIL.n345 B 0.010917f
C415 VTAIL.n346 B 0.011559f
C416 VTAIL.n347 B 0.025803f
C417 VTAIL.n348 B 0.051255f
C418 VTAIL.n349 B 0.011559f
C419 VTAIL.n350 B 0.010917f
C420 VTAIL.n351 B 0.043906f
C421 VTAIL.n352 B 0.028109f
C422 VTAIL.n353 B 0.104513f
C423 VTAIL.t11 B 0.169692f
C424 VTAIL.t15 B 0.169692f
C425 VTAIL.n354 B 1.43501f
C426 VTAIL.n355 B 0.31997f
C427 VTAIL.n356 B 0.025951f
C428 VTAIL.n357 B 0.020316f
C429 VTAIL.n358 B 0.010917f
C430 VTAIL.n359 B 0.025803f
C431 VTAIL.n360 B 0.011559f
C432 VTAIL.n361 B 0.020316f
C433 VTAIL.n362 B 0.010917f
C434 VTAIL.n363 B 0.025803f
C435 VTAIL.n364 B 0.011559f
C436 VTAIL.n365 B 0.020316f
C437 VTAIL.n366 B 0.010917f
C438 VTAIL.n367 B 0.025803f
C439 VTAIL.n368 B 0.025803f
C440 VTAIL.n369 B 0.011559f
C441 VTAIL.n370 B 0.020316f
C442 VTAIL.n371 B 0.010917f
C443 VTAIL.n372 B 0.025803f
C444 VTAIL.n373 B 0.011559f
C445 VTAIL.n374 B 0.135322f
C446 VTAIL.t12 B 0.043424f
C447 VTAIL.n375 B 0.019353f
C448 VTAIL.n376 B 0.018241f
C449 VTAIL.n377 B 0.010917f
C450 VTAIL.n378 B 0.895676f
C451 VTAIL.n379 B 0.020316f
C452 VTAIL.n380 B 0.010917f
C453 VTAIL.n381 B 0.011559f
C454 VTAIL.n382 B 0.025803f
C455 VTAIL.n383 B 0.025803f
C456 VTAIL.n384 B 0.011559f
C457 VTAIL.n385 B 0.010917f
C458 VTAIL.n386 B 0.020316f
C459 VTAIL.n387 B 0.020316f
C460 VTAIL.n388 B 0.010917f
C461 VTAIL.n389 B 0.011559f
C462 VTAIL.n390 B 0.025803f
C463 VTAIL.n391 B 0.025803f
C464 VTAIL.n392 B 0.011559f
C465 VTAIL.n393 B 0.010917f
C466 VTAIL.n394 B 0.020316f
C467 VTAIL.n395 B 0.020316f
C468 VTAIL.n396 B 0.010917f
C469 VTAIL.n397 B 0.011238f
C470 VTAIL.n398 B 0.011238f
C471 VTAIL.n399 B 0.025803f
C472 VTAIL.n400 B 0.025803f
C473 VTAIL.n401 B 0.011559f
C474 VTAIL.n402 B 0.010917f
C475 VTAIL.n403 B 0.020316f
C476 VTAIL.n404 B 0.020316f
C477 VTAIL.n405 B 0.010917f
C478 VTAIL.n406 B 0.011559f
C479 VTAIL.n407 B 0.025803f
C480 VTAIL.n408 B 0.051255f
C481 VTAIL.n409 B 0.011559f
C482 VTAIL.n410 B 0.010917f
C483 VTAIL.n411 B 0.043906f
C484 VTAIL.n412 B 0.028109f
C485 VTAIL.n413 B 1.00434f
C486 VTAIL.n414 B 0.025951f
C487 VTAIL.n415 B 0.020316f
C488 VTAIL.n416 B 0.010917f
C489 VTAIL.n417 B 0.025803f
C490 VTAIL.n418 B 0.011559f
C491 VTAIL.n419 B 0.020316f
C492 VTAIL.n420 B 0.010917f
C493 VTAIL.n421 B 0.025803f
C494 VTAIL.n422 B 0.011559f
C495 VTAIL.n423 B 0.020316f
C496 VTAIL.n424 B 0.010917f
C497 VTAIL.n425 B 0.025803f
C498 VTAIL.n426 B 0.011559f
C499 VTAIL.n427 B 0.020316f
C500 VTAIL.n428 B 0.010917f
C501 VTAIL.n429 B 0.025803f
C502 VTAIL.n430 B 0.011559f
C503 VTAIL.n431 B 0.135322f
C504 VTAIL.t0 B 0.043424f
C505 VTAIL.n432 B 0.019353f
C506 VTAIL.n433 B 0.018241f
C507 VTAIL.n434 B 0.010917f
C508 VTAIL.n435 B 0.895676f
C509 VTAIL.n436 B 0.020316f
C510 VTAIL.n437 B 0.010917f
C511 VTAIL.n438 B 0.011559f
C512 VTAIL.n439 B 0.025803f
C513 VTAIL.n440 B 0.025803f
C514 VTAIL.n441 B 0.011559f
C515 VTAIL.n442 B 0.010917f
C516 VTAIL.n443 B 0.020316f
C517 VTAIL.n444 B 0.020316f
C518 VTAIL.n445 B 0.010917f
C519 VTAIL.n446 B 0.011559f
C520 VTAIL.n447 B 0.025803f
C521 VTAIL.n448 B 0.025803f
C522 VTAIL.n449 B 0.025803f
C523 VTAIL.n450 B 0.011559f
C524 VTAIL.n451 B 0.010917f
C525 VTAIL.n452 B 0.020316f
C526 VTAIL.n453 B 0.020316f
C527 VTAIL.n454 B 0.010917f
C528 VTAIL.n455 B 0.011238f
C529 VTAIL.n456 B 0.011238f
C530 VTAIL.n457 B 0.025803f
C531 VTAIL.n458 B 0.025803f
C532 VTAIL.n459 B 0.011559f
C533 VTAIL.n460 B 0.010917f
C534 VTAIL.n461 B 0.020316f
C535 VTAIL.n462 B 0.020316f
C536 VTAIL.n463 B 0.010917f
C537 VTAIL.n464 B 0.011559f
C538 VTAIL.n465 B 0.025803f
C539 VTAIL.n466 B 0.051255f
C540 VTAIL.n467 B 0.011559f
C541 VTAIL.n468 B 0.010917f
C542 VTAIL.n469 B 0.043906f
C543 VTAIL.n470 B 0.028109f
C544 VTAIL.n471 B 1.00053f
C545 VDD1.t0 B 0.228497f
C546 VDD1.t5 B 0.228497f
C547 VDD1.n0 B 2.02012f
C548 VDD1.t1 B 0.228497f
C549 VDD1.t4 B 0.228497f
C550 VDD1.n1 B 2.01939f
C551 VDD1.t2 B 0.228497f
C552 VDD1.t3 B 0.228497f
C553 VDD1.n2 B 2.01939f
C554 VDD1.n3 B 2.34262f
C555 VDD1.t6 B 0.228497f
C556 VDD1.t7 B 0.228497f
C557 VDD1.n4 B 2.01713f
C558 VDD1.n5 B 2.41788f
C559 VP.n0 B 0.044941f
C560 VP.n1 B 0.010198f
C561 VP.n2 B 0.044941f
C562 VP.n3 B 0.044941f
C563 VP.t3 B 0.95068f
C564 VP.t0 B 0.95068f
C565 VP.n4 B 0.044941f
C566 VP.t4 B 0.95068f
C567 VP.n5 B 0.391649f
C568 VP.t1 B 0.970092f
C569 VP.n6 B 0.372305f
C570 VP.n7 B 0.186886f
C571 VP.n8 B 0.010198f
C572 VP.n9 B 0.387582f
C573 VP.n10 B 0.010198f
C574 VP.n11 B 0.384672f
C575 VP.n12 B 1.77475f
C576 VP.n13 B 1.81424f
C577 VP.t2 B 0.95068f
C578 VP.n14 B 0.384672f
C579 VP.n15 B 0.010198f
C580 VP.t5 B 0.95068f
C581 VP.n16 B 0.387582f
C582 VP.n17 B 0.044941f
C583 VP.n18 B 0.044941f
C584 VP.n19 B 0.044941f
C585 VP.t7 B 0.95068f
C586 VP.n20 B 0.387582f
C587 VP.n21 B 0.010198f
C588 VP.t6 B 0.95068f
C589 VP.n22 B 0.384672f
C590 VP.n23 B 0.034828f
.ends

