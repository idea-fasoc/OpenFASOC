* NGSPICE file created from diff_pair_sample_0623.ext - technology: sky130A

.subckt diff_pair_sample_0623 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t2 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=0.77055 ps=5 w=4.67 l=3.62
X1 VTAIL.t3 VP.t0 VDD1.t5 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=0.77055 ps=5 w=4.67 l=3.62
X2 VDD2.t5 VN.t1 VTAIL.t8 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0.77055 ps=5 w=4.67 l=3.62
X3 VTAIL.t2 VP.t1 VDD1.t4 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=0.77055 ps=5 w=4.67 l=3.62
X4 VTAIL.t7 VN.t2 VDD2.t3 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=0.77055 ps=5 w=4.67 l=3.62
X5 B.t11 B.t9 B.t10 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0 ps=0 w=4.67 l=3.62
X6 VDD1.t3 VP.t2 VTAIL.t10 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0.77055 ps=5 w=4.67 l=3.62
X7 VDD2.t4 VN.t3 VTAIL.t6 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=1.8213 ps=10.12 w=4.67 l=3.62
X8 VDD1.t2 VP.t3 VTAIL.t0 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0.77055 ps=5 w=4.67 l=3.62
X9 VDD2.t0 VN.t4 VTAIL.t5 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=1.8213 ps=10.12 w=4.67 l=3.62
X10 VDD2.t1 VN.t5 VTAIL.t4 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0.77055 ps=5 w=4.67 l=3.62
X11 VDD1.t1 VP.t4 VTAIL.t11 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=1.8213 ps=10.12 w=4.67 l=3.62
X12 VDD1.t0 VP.t5 VTAIL.t1 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=0.77055 pd=5 as=1.8213 ps=10.12 w=4.67 l=3.62
X13 B.t8 B.t6 B.t7 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0 ps=0 w=4.67 l=3.62
X14 B.t5 B.t3 B.t4 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0 ps=0 w=4.67 l=3.62
X15 B.t2 B.t0 B.t1 w_n4130_n1902# sky130_fd_pr__pfet_01v8 ad=1.8213 pd=10.12 as=0 ps=0 w=4.67 l=3.62
R0 VN.n38 VN.n37 161.3
R1 VN.n36 VN.n21 161.3
R2 VN.n35 VN.n34 161.3
R3 VN.n33 VN.n22 161.3
R4 VN.n32 VN.n31 161.3
R5 VN.n30 VN.n23 161.3
R6 VN.n29 VN.n28 161.3
R7 VN.n27 VN.n24 161.3
R8 VN.n18 VN.n17 161.3
R9 VN.n16 VN.n1 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n2 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n10 VN.n3 161.3
R14 VN.n9 VN.n8 161.3
R15 VN.n7 VN.n4 161.3
R16 VN.n19 VN.n0 80.2806
R17 VN.n39 VN.n20 80.2806
R18 VN.n26 VN.t3 64.4522
R19 VN.n6 VN.t5 64.4522
R20 VN.n6 VN.n5 62.3641
R21 VN.n26 VN.n25 62.3641
R22 VN.n11 VN.n2 56.5193
R23 VN.n31 VN.n22 56.5193
R24 VN VN.n39 47.4033
R25 VN.n5 VN.t0 31.0908
R26 VN.n0 VN.t4 31.0908
R27 VN.n25 VN.t2 31.0908
R28 VN.n20 VN.t1 31.0908
R29 VN.n9 VN.n4 24.4675
R30 VN.n10 VN.n9 24.4675
R31 VN.n11 VN.n10 24.4675
R32 VN.n15 VN.n2 24.4675
R33 VN.n16 VN.n15 24.4675
R34 VN.n17 VN.n16 24.4675
R35 VN.n31 VN.n30 24.4675
R36 VN.n30 VN.n29 24.4675
R37 VN.n29 VN.n24 24.4675
R38 VN.n37 VN.n36 24.4675
R39 VN.n36 VN.n35 24.4675
R40 VN.n35 VN.n22 24.4675
R41 VN.n5 VN.n4 12.234
R42 VN.n25 VN.n24 12.234
R43 VN.n17 VN.n0 9.7873
R44 VN.n37 VN.n20 9.7873
R45 VN.n27 VN.n26 3.16397
R46 VN.n7 VN.n6 3.16397
R47 VN.n39 VN.n38 0.354971
R48 VN.n19 VN.n18 0.354971
R49 VN VN.n19 0.26696
R50 VN.n38 VN.n21 0.189894
R51 VN.n34 VN.n21 0.189894
R52 VN.n34 VN.n33 0.189894
R53 VN.n33 VN.n32 0.189894
R54 VN.n32 VN.n23 0.189894
R55 VN.n28 VN.n23 0.189894
R56 VN.n28 VN.n27 0.189894
R57 VN.n8 VN.n7 0.189894
R58 VN.n8 VN.n3 0.189894
R59 VN.n12 VN.n3 0.189894
R60 VN.n13 VN.n12 0.189894
R61 VN.n14 VN.n13 0.189894
R62 VN.n14 VN.n1 0.189894
R63 VN.n18 VN.n1 0.189894
R64 VDD2.n43 VDD2.n25 756.745
R65 VDD2.n18 VDD2.n0 756.745
R66 VDD2.n44 VDD2.n43 585
R67 VDD2.n42 VDD2.n41 585
R68 VDD2.n29 VDD2.n28 585
R69 VDD2.n36 VDD2.n35 585
R70 VDD2.n34 VDD2.n33 585
R71 VDD2.n9 VDD2.n8 585
R72 VDD2.n11 VDD2.n10 585
R73 VDD2.n4 VDD2.n3 585
R74 VDD2.n17 VDD2.n16 585
R75 VDD2.n19 VDD2.n18 585
R76 VDD2.n32 VDD2.t5 328.587
R77 VDD2.n7 VDD2.t1 328.587
R78 VDD2.n43 VDD2.n42 171.744
R79 VDD2.n42 VDD2.n28 171.744
R80 VDD2.n35 VDD2.n28 171.744
R81 VDD2.n35 VDD2.n34 171.744
R82 VDD2.n10 VDD2.n9 171.744
R83 VDD2.n10 VDD2.n3 171.744
R84 VDD2.n17 VDD2.n3 171.744
R85 VDD2.n18 VDD2.n17 171.744
R86 VDD2.n24 VDD2.n23 107.008
R87 VDD2 VDD2.n49 107.007
R88 VDD2.n34 VDD2.t5 85.8723
R89 VDD2.n9 VDD2.t1 85.8723
R90 VDD2.n24 VDD2.n22 53.496
R91 VDD2.n48 VDD2.n47 50.9975
R92 VDD2.n48 VDD2.n24 38.808
R93 VDD2.n33 VDD2.n32 16.3651
R94 VDD2.n8 VDD2.n7 16.3651
R95 VDD2.n36 VDD2.n31 12.8005
R96 VDD2.n11 VDD2.n6 12.8005
R97 VDD2.n37 VDD2.n29 12.0247
R98 VDD2.n12 VDD2.n4 12.0247
R99 VDD2.n41 VDD2.n40 11.249
R100 VDD2.n16 VDD2.n15 11.249
R101 VDD2.n44 VDD2.n27 10.4732
R102 VDD2.n19 VDD2.n2 10.4732
R103 VDD2.n45 VDD2.n25 9.69747
R104 VDD2.n20 VDD2.n0 9.69747
R105 VDD2.n47 VDD2.n46 9.45567
R106 VDD2.n22 VDD2.n21 9.45567
R107 VDD2.n46 VDD2.n45 9.3005
R108 VDD2.n27 VDD2.n26 9.3005
R109 VDD2.n40 VDD2.n39 9.3005
R110 VDD2.n38 VDD2.n37 9.3005
R111 VDD2.n31 VDD2.n30 9.3005
R112 VDD2.n21 VDD2.n20 9.3005
R113 VDD2.n2 VDD2.n1 9.3005
R114 VDD2.n15 VDD2.n14 9.3005
R115 VDD2.n13 VDD2.n12 9.3005
R116 VDD2.n6 VDD2.n5 9.3005
R117 VDD2.n49 VDD2.t3 6.96089
R118 VDD2.n49 VDD2.t4 6.96089
R119 VDD2.n23 VDD2.t2 6.96089
R120 VDD2.n23 VDD2.t0 6.96089
R121 VDD2.n47 VDD2.n25 4.26717
R122 VDD2.n22 VDD2.n0 4.26717
R123 VDD2.n32 VDD2.n30 3.73474
R124 VDD2.n7 VDD2.n5 3.73474
R125 VDD2.n45 VDD2.n44 3.49141
R126 VDD2.n20 VDD2.n19 3.49141
R127 VDD2.n41 VDD2.n27 2.71565
R128 VDD2.n16 VDD2.n2 2.71565
R129 VDD2 VDD2.n48 2.61257
R130 VDD2.n40 VDD2.n29 1.93989
R131 VDD2.n15 VDD2.n4 1.93989
R132 VDD2.n37 VDD2.n36 1.16414
R133 VDD2.n12 VDD2.n11 1.16414
R134 VDD2.n33 VDD2.n31 0.388379
R135 VDD2.n8 VDD2.n6 0.388379
R136 VDD2.n46 VDD2.n26 0.155672
R137 VDD2.n39 VDD2.n26 0.155672
R138 VDD2.n39 VDD2.n38 0.155672
R139 VDD2.n38 VDD2.n30 0.155672
R140 VDD2.n13 VDD2.n5 0.155672
R141 VDD2.n14 VDD2.n13 0.155672
R142 VDD2.n14 VDD2.n1 0.155672
R143 VDD2.n21 VDD2.n1 0.155672
R144 VTAIL.n98 VTAIL.n80 756.745
R145 VTAIL.n20 VTAIL.n2 756.745
R146 VTAIL.n74 VTAIL.n56 756.745
R147 VTAIL.n48 VTAIL.n30 756.745
R148 VTAIL.n89 VTAIL.n88 585
R149 VTAIL.n91 VTAIL.n90 585
R150 VTAIL.n84 VTAIL.n83 585
R151 VTAIL.n97 VTAIL.n96 585
R152 VTAIL.n99 VTAIL.n98 585
R153 VTAIL.n11 VTAIL.n10 585
R154 VTAIL.n13 VTAIL.n12 585
R155 VTAIL.n6 VTAIL.n5 585
R156 VTAIL.n19 VTAIL.n18 585
R157 VTAIL.n21 VTAIL.n20 585
R158 VTAIL.n75 VTAIL.n74 585
R159 VTAIL.n73 VTAIL.n72 585
R160 VTAIL.n60 VTAIL.n59 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n65 VTAIL.n64 585
R163 VTAIL.n49 VTAIL.n48 585
R164 VTAIL.n47 VTAIL.n46 585
R165 VTAIL.n34 VTAIL.n33 585
R166 VTAIL.n41 VTAIL.n40 585
R167 VTAIL.n39 VTAIL.n38 585
R168 VTAIL.n87 VTAIL.t5 328.587
R169 VTAIL.n9 VTAIL.t11 328.587
R170 VTAIL.n63 VTAIL.t1 328.587
R171 VTAIL.n37 VTAIL.t6 328.587
R172 VTAIL.n90 VTAIL.n89 171.744
R173 VTAIL.n90 VTAIL.n83 171.744
R174 VTAIL.n97 VTAIL.n83 171.744
R175 VTAIL.n98 VTAIL.n97 171.744
R176 VTAIL.n12 VTAIL.n11 171.744
R177 VTAIL.n12 VTAIL.n5 171.744
R178 VTAIL.n19 VTAIL.n5 171.744
R179 VTAIL.n20 VTAIL.n19 171.744
R180 VTAIL.n74 VTAIL.n73 171.744
R181 VTAIL.n73 VTAIL.n59 171.744
R182 VTAIL.n66 VTAIL.n59 171.744
R183 VTAIL.n66 VTAIL.n65 171.744
R184 VTAIL.n48 VTAIL.n47 171.744
R185 VTAIL.n47 VTAIL.n33 171.744
R186 VTAIL.n40 VTAIL.n33 171.744
R187 VTAIL.n40 VTAIL.n39 171.744
R188 VTAIL.n55 VTAIL.n54 89.5344
R189 VTAIL.n29 VTAIL.n28 89.5344
R190 VTAIL.n1 VTAIL.n0 89.5342
R191 VTAIL.n27 VTAIL.n26 89.5342
R192 VTAIL.n89 VTAIL.t5 85.8723
R193 VTAIL.n11 VTAIL.t11 85.8723
R194 VTAIL.n65 VTAIL.t1 85.8723
R195 VTAIL.n39 VTAIL.t6 85.8723
R196 VTAIL.n103 VTAIL.n102 34.3187
R197 VTAIL.n25 VTAIL.n24 34.3187
R198 VTAIL.n79 VTAIL.n78 34.3187
R199 VTAIL.n53 VTAIL.n52 34.3187
R200 VTAIL.n29 VTAIL.n27 23.2031
R201 VTAIL.n103 VTAIL.n79 19.7979
R202 VTAIL.n88 VTAIL.n87 16.3651
R203 VTAIL.n10 VTAIL.n9 16.3651
R204 VTAIL.n64 VTAIL.n63 16.3651
R205 VTAIL.n38 VTAIL.n37 16.3651
R206 VTAIL.n91 VTAIL.n86 12.8005
R207 VTAIL.n13 VTAIL.n8 12.8005
R208 VTAIL.n67 VTAIL.n62 12.8005
R209 VTAIL.n41 VTAIL.n36 12.8005
R210 VTAIL.n92 VTAIL.n84 12.0247
R211 VTAIL.n14 VTAIL.n6 12.0247
R212 VTAIL.n68 VTAIL.n60 12.0247
R213 VTAIL.n42 VTAIL.n34 12.0247
R214 VTAIL.n96 VTAIL.n95 11.249
R215 VTAIL.n18 VTAIL.n17 11.249
R216 VTAIL.n72 VTAIL.n71 11.249
R217 VTAIL.n46 VTAIL.n45 11.249
R218 VTAIL.n99 VTAIL.n82 10.4732
R219 VTAIL.n21 VTAIL.n4 10.4732
R220 VTAIL.n75 VTAIL.n58 10.4732
R221 VTAIL.n49 VTAIL.n32 10.4732
R222 VTAIL.n100 VTAIL.n80 9.69747
R223 VTAIL.n22 VTAIL.n2 9.69747
R224 VTAIL.n76 VTAIL.n56 9.69747
R225 VTAIL.n50 VTAIL.n30 9.69747
R226 VTAIL.n102 VTAIL.n101 9.45567
R227 VTAIL.n24 VTAIL.n23 9.45567
R228 VTAIL.n78 VTAIL.n77 9.45567
R229 VTAIL.n52 VTAIL.n51 9.45567
R230 VTAIL.n101 VTAIL.n100 9.3005
R231 VTAIL.n82 VTAIL.n81 9.3005
R232 VTAIL.n95 VTAIL.n94 9.3005
R233 VTAIL.n93 VTAIL.n92 9.3005
R234 VTAIL.n86 VTAIL.n85 9.3005
R235 VTAIL.n23 VTAIL.n22 9.3005
R236 VTAIL.n4 VTAIL.n3 9.3005
R237 VTAIL.n17 VTAIL.n16 9.3005
R238 VTAIL.n15 VTAIL.n14 9.3005
R239 VTAIL.n8 VTAIL.n7 9.3005
R240 VTAIL.n77 VTAIL.n76 9.3005
R241 VTAIL.n58 VTAIL.n57 9.3005
R242 VTAIL.n71 VTAIL.n70 9.3005
R243 VTAIL.n69 VTAIL.n68 9.3005
R244 VTAIL.n62 VTAIL.n61 9.3005
R245 VTAIL.n51 VTAIL.n50 9.3005
R246 VTAIL.n32 VTAIL.n31 9.3005
R247 VTAIL.n45 VTAIL.n44 9.3005
R248 VTAIL.n43 VTAIL.n42 9.3005
R249 VTAIL.n36 VTAIL.n35 9.3005
R250 VTAIL.n0 VTAIL.t4 6.96089
R251 VTAIL.n0 VTAIL.t9 6.96089
R252 VTAIL.n26 VTAIL.t0 6.96089
R253 VTAIL.n26 VTAIL.t2 6.96089
R254 VTAIL.n54 VTAIL.t10 6.96089
R255 VTAIL.n54 VTAIL.t3 6.96089
R256 VTAIL.n28 VTAIL.t8 6.96089
R257 VTAIL.n28 VTAIL.t7 6.96089
R258 VTAIL.n102 VTAIL.n80 4.26717
R259 VTAIL.n24 VTAIL.n2 4.26717
R260 VTAIL.n78 VTAIL.n56 4.26717
R261 VTAIL.n52 VTAIL.n30 4.26717
R262 VTAIL.n87 VTAIL.n85 3.73474
R263 VTAIL.n9 VTAIL.n7 3.73474
R264 VTAIL.n63 VTAIL.n61 3.73474
R265 VTAIL.n37 VTAIL.n35 3.73474
R266 VTAIL.n100 VTAIL.n99 3.49141
R267 VTAIL.n22 VTAIL.n21 3.49141
R268 VTAIL.n76 VTAIL.n75 3.49141
R269 VTAIL.n50 VTAIL.n49 3.49141
R270 VTAIL.n53 VTAIL.n29 3.40567
R271 VTAIL.n79 VTAIL.n55 3.40567
R272 VTAIL.n27 VTAIL.n25 3.40567
R273 VTAIL.n96 VTAIL.n82 2.71565
R274 VTAIL.n18 VTAIL.n4 2.71565
R275 VTAIL.n72 VTAIL.n58 2.71565
R276 VTAIL.n46 VTAIL.n32 2.71565
R277 VTAIL VTAIL.n103 2.49619
R278 VTAIL.n55 VTAIL.n53 2.17291
R279 VTAIL.n25 VTAIL.n1 2.17291
R280 VTAIL.n95 VTAIL.n84 1.93989
R281 VTAIL.n17 VTAIL.n6 1.93989
R282 VTAIL.n71 VTAIL.n60 1.93989
R283 VTAIL.n45 VTAIL.n34 1.93989
R284 VTAIL.n92 VTAIL.n91 1.16414
R285 VTAIL.n14 VTAIL.n13 1.16414
R286 VTAIL.n68 VTAIL.n67 1.16414
R287 VTAIL.n42 VTAIL.n41 1.16414
R288 VTAIL VTAIL.n1 0.909983
R289 VTAIL.n88 VTAIL.n86 0.388379
R290 VTAIL.n10 VTAIL.n8 0.388379
R291 VTAIL.n64 VTAIL.n62 0.388379
R292 VTAIL.n38 VTAIL.n36 0.388379
R293 VTAIL.n93 VTAIL.n85 0.155672
R294 VTAIL.n94 VTAIL.n93 0.155672
R295 VTAIL.n94 VTAIL.n81 0.155672
R296 VTAIL.n101 VTAIL.n81 0.155672
R297 VTAIL.n15 VTAIL.n7 0.155672
R298 VTAIL.n16 VTAIL.n15 0.155672
R299 VTAIL.n16 VTAIL.n3 0.155672
R300 VTAIL.n23 VTAIL.n3 0.155672
R301 VTAIL.n77 VTAIL.n57 0.155672
R302 VTAIL.n70 VTAIL.n57 0.155672
R303 VTAIL.n70 VTAIL.n69 0.155672
R304 VTAIL.n69 VTAIL.n61 0.155672
R305 VTAIL.n51 VTAIL.n31 0.155672
R306 VTAIL.n44 VTAIL.n31 0.155672
R307 VTAIL.n44 VTAIL.n43 0.155672
R308 VTAIL.n43 VTAIL.n35 0.155672
R309 VP.n16 VP.n13 161.3
R310 VP.n18 VP.n17 161.3
R311 VP.n19 VP.n12 161.3
R312 VP.n21 VP.n20 161.3
R313 VP.n22 VP.n11 161.3
R314 VP.n24 VP.n23 161.3
R315 VP.n25 VP.n10 161.3
R316 VP.n27 VP.n26 161.3
R317 VP.n55 VP.n54 161.3
R318 VP.n53 VP.n1 161.3
R319 VP.n52 VP.n51 161.3
R320 VP.n50 VP.n2 161.3
R321 VP.n49 VP.n48 161.3
R322 VP.n47 VP.n3 161.3
R323 VP.n46 VP.n45 161.3
R324 VP.n44 VP.n4 161.3
R325 VP.n43 VP.n42 161.3
R326 VP.n40 VP.n5 161.3
R327 VP.n39 VP.n38 161.3
R328 VP.n37 VP.n6 161.3
R329 VP.n36 VP.n35 161.3
R330 VP.n34 VP.n7 161.3
R331 VP.n33 VP.n32 161.3
R332 VP.n31 VP.n8 161.3
R333 VP.n30 VP.n29 80.2806
R334 VP.n56 VP.n0 80.2806
R335 VP.n28 VP.n9 80.2806
R336 VP.n15 VP.t2 64.452
R337 VP.n15 VP.n14 62.3641
R338 VP.n35 VP.n6 56.5193
R339 VP.n48 VP.n2 56.5193
R340 VP.n20 VP.n11 56.5193
R341 VP.n30 VP.n28 47.238
R342 VP.n29 VP.t3 31.0908
R343 VP.n41 VP.t1 31.0908
R344 VP.n0 VP.t4 31.0908
R345 VP.n9 VP.t5 31.0908
R346 VP.n14 VP.t0 31.0908
R347 VP.n33 VP.n8 24.4675
R348 VP.n34 VP.n33 24.4675
R349 VP.n35 VP.n34 24.4675
R350 VP.n39 VP.n6 24.4675
R351 VP.n40 VP.n39 24.4675
R352 VP.n42 VP.n40 24.4675
R353 VP.n46 VP.n4 24.4675
R354 VP.n47 VP.n46 24.4675
R355 VP.n48 VP.n47 24.4675
R356 VP.n52 VP.n2 24.4675
R357 VP.n53 VP.n52 24.4675
R358 VP.n54 VP.n53 24.4675
R359 VP.n24 VP.n11 24.4675
R360 VP.n25 VP.n24 24.4675
R361 VP.n26 VP.n25 24.4675
R362 VP.n18 VP.n13 24.4675
R363 VP.n19 VP.n18 24.4675
R364 VP.n20 VP.n19 24.4675
R365 VP.n42 VP.n41 12.234
R366 VP.n41 VP.n4 12.234
R367 VP.n14 VP.n13 12.234
R368 VP.n29 VP.n8 9.7873
R369 VP.n54 VP.n0 9.7873
R370 VP.n26 VP.n9 9.7873
R371 VP.n16 VP.n15 3.16396
R372 VP.n28 VP.n27 0.354971
R373 VP.n31 VP.n30 0.354971
R374 VP.n56 VP.n55 0.354971
R375 VP VP.n56 0.26696
R376 VP.n17 VP.n16 0.189894
R377 VP.n17 VP.n12 0.189894
R378 VP.n21 VP.n12 0.189894
R379 VP.n22 VP.n21 0.189894
R380 VP.n23 VP.n22 0.189894
R381 VP.n23 VP.n10 0.189894
R382 VP.n27 VP.n10 0.189894
R383 VP.n32 VP.n31 0.189894
R384 VP.n32 VP.n7 0.189894
R385 VP.n36 VP.n7 0.189894
R386 VP.n37 VP.n36 0.189894
R387 VP.n38 VP.n37 0.189894
R388 VP.n38 VP.n5 0.189894
R389 VP.n43 VP.n5 0.189894
R390 VP.n44 VP.n43 0.189894
R391 VP.n45 VP.n44 0.189894
R392 VP.n45 VP.n3 0.189894
R393 VP.n49 VP.n3 0.189894
R394 VP.n50 VP.n49 0.189894
R395 VP.n51 VP.n50 0.189894
R396 VP.n51 VP.n1 0.189894
R397 VP.n55 VP.n1 0.189894
R398 VDD1.n18 VDD1.n0 756.745
R399 VDD1.n41 VDD1.n23 756.745
R400 VDD1.n19 VDD1.n18 585
R401 VDD1.n17 VDD1.n16 585
R402 VDD1.n4 VDD1.n3 585
R403 VDD1.n11 VDD1.n10 585
R404 VDD1.n9 VDD1.n8 585
R405 VDD1.n32 VDD1.n31 585
R406 VDD1.n34 VDD1.n33 585
R407 VDD1.n27 VDD1.n26 585
R408 VDD1.n40 VDD1.n39 585
R409 VDD1.n42 VDD1.n41 585
R410 VDD1.n7 VDD1.t3 328.587
R411 VDD1.n30 VDD1.t2 328.587
R412 VDD1.n18 VDD1.n17 171.744
R413 VDD1.n17 VDD1.n3 171.744
R414 VDD1.n10 VDD1.n3 171.744
R415 VDD1.n10 VDD1.n9 171.744
R416 VDD1.n33 VDD1.n32 171.744
R417 VDD1.n33 VDD1.n26 171.744
R418 VDD1.n40 VDD1.n26 171.744
R419 VDD1.n41 VDD1.n40 171.744
R420 VDD1.n47 VDD1.n46 107.008
R421 VDD1.n49 VDD1.n48 106.213
R422 VDD1.n9 VDD1.t3 85.8723
R423 VDD1.n32 VDD1.t2 85.8723
R424 VDD1 VDD1.n22 53.6095
R425 VDD1.n47 VDD1.n45 53.496
R426 VDD1.n49 VDD1.n47 41.0936
R427 VDD1.n8 VDD1.n7 16.3651
R428 VDD1.n31 VDD1.n30 16.3651
R429 VDD1.n11 VDD1.n6 12.8005
R430 VDD1.n34 VDD1.n29 12.8005
R431 VDD1.n12 VDD1.n4 12.0247
R432 VDD1.n35 VDD1.n27 12.0247
R433 VDD1.n16 VDD1.n15 11.249
R434 VDD1.n39 VDD1.n38 11.249
R435 VDD1.n19 VDD1.n2 10.4732
R436 VDD1.n42 VDD1.n25 10.4732
R437 VDD1.n20 VDD1.n0 9.69747
R438 VDD1.n43 VDD1.n23 9.69747
R439 VDD1.n22 VDD1.n21 9.45567
R440 VDD1.n45 VDD1.n44 9.45567
R441 VDD1.n21 VDD1.n20 9.3005
R442 VDD1.n2 VDD1.n1 9.3005
R443 VDD1.n15 VDD1.n14 9.3005
R444 VDD1.n13 VDD1.n12 9.3005
R445 VDD1.n6 VDD1.n5 9.3005
R446 VDD1.n44 VDD1.n43 9.3005
R447 VDD1.n25 VDD1.n24 9.3005
R448 VDD1.n38 VDD1.n37 9.3005
R449 VDD1.n36 VDD1.n35 9.3005
R450 VDD1.n29 VDD1.n28 9.3005
R451 VDD1.n48 VDD1.t5 6.96089
R452 VDD1.n48 VDD1.t0 6.96089
R453 VDD1.n46 VDD1.t4 6.96089
R454 VDD1.n46 VDD1.t1 6.96089
R455 VDD1.n22 VDD1.n0 4.26717
R456 VDD1.n45 VDD1.n23 4.26717
R457 VDD1.n7 VDD1.n5 3.73474
R458 VDD1.n30 VDD1.n28 3.73474
R459 VDD1.n20 VDD1.n19 3.49141
R460 VDD1.n43 VDD1.n42 3.49141
R461 VDD1.n16 VDD1.n2 2.71565
R462 VDD1.n39 VDD1.n25 2.71565
R463 VDD1.n15 VDD1.n4 1.93989
R464 VDD1.n38 VDD1.n27 1.93989
R465 VDD1.n12 VDD1.n11 1.16414
R466 VDD1.n35 VDD1.n34 1.16414
R467 VDD1 VDD1.n49 0.793603
R468 VDD1.n8 VDD1.n6 0.388379
R469 VDD1.n31 VDD1.n29 0.388379
R470 VDD1.n21 VDD1.n1 0.155672
R471 VDD1.n14 VDD1.n1 0.155672
R472 VDD1.n14 VDD1.n13 0.155672
R473 VDD1.n13 VDD1.n5 0.155672
R474 VDD1.n36 VDD1.n28 0.155672
R475 VDD1.n37 VDD1.n36 0.155672
R476 VDD1.n37 VDD1.n24 0.155672
R477 VDD1.n44 VDD1.n24 0.155672
R478 B.n325 B.n324 585
R479 B.n323 B.n114 585
R480 B.n322 B.n321 585
R481 B.n320 B.n115 585
R482 B.n319 B.n318 585
R483 B.n317 B.n116 585
R484 B.n316 B.n315 585
R485 B.n314 B.n117 585
R486 B.n313 B.n312 585
R487 B.n311 B.n118 585
R488 B.n310 B.n309 585
R489 B.n308 B.n119 585
R490 B.n307 B.n306 585
R491 B.n305 B.n120 585
R492 B.n304 B.n303 585
R493 B.n302 B.n121 585
R494 B.n301 B.n300 585
R495 B.n299 B.n122 585
R496 B.n298 B.n297 585
R497 B.n296 B.n123 585
R498 B.n294 B.n293 585
R499 B.n292 B.n126 585
R500 B.n291 B.n290 585
R501 B.n289 B.n127 585
R502 B.n288 B.n287 585
R503 B.n286 B.n128 585
R504 B.n285 B.n284 585
R505 B.n283 B.n129 585
R506 B.n282 B.n281 585
R507 B.n280 B.n130 585
R508 B.n279 B.n278 585
R509 B.n274 B.n131 585
R510 B.n273 B.n272 585
R511 B.n271 B.n132 585
R512 B.n270 B.n269 585
R513 B.n268 B.n133 585
R514 B.n267 B.n266 585
R515 B.n265 B.n134 585
R516 B.n264 B.n263 585
R517 B.n262 B.n135 585
R518 B.n261 B.n260 585
R519 B.n259 B.n136 585
R520 B.n258 B.n257 585
R521 B.n256 B.n137 585
R522 B.n255 B.n254 585
R523 B.n253 B.n138 585
R524 B.n252 B.n251 585
R525 B.n250 B.n139 585
R526 B.n249 B.n248 585
R527 B.n247 B.n140 585
R528 B.n326 B.n113 585
R529 B.n328 B.n327 585
R530 B.n329 B.n112 585
R531 B.n331 B.n330 585
R532 B.n332 B.n111 585
R533 B.n334 B.n333 585
R534 B.n335 B.n110 585
R535 B.n337 B.n336 585
R536 B.n338 B.n109 585
R537 B.n340 B.n339 585
R538 B.n341 B.n108 585
R539 B.n343 B.n342 585
R540 B.n344 B.n107 585
R541 B.n346 B.n345 585
R542 B.n347 B.n106 585
R543 B.n349 B.n348 585
R544 B.n350 B.n105 585
R545 B.n352 B.n351 585
R546 B.n353 B.n104 585
R547 B.n355 B.n354 585
R548 B.n356 B.n103 585
R549 B.n358 B.n357 585
R550 B.n359 B.n102 585
R551 B.n361 B.n360 585
R552 B.n362 B.n101 585
R553 B.n364 B.n363 585
R554 B.n365 B.n100 585
R555 B.n367 B.n366 585
R556 B.n368 B.n99 585
R557 B.n370 B.n369 585
R558 B.n371 B.n98 585
R559 B.n373 B.n372 585
R560 B.n374 B.n97 585
R561 B.n376 B.n375 585
R562 B.n377 B.n96 585
R563 B.n379 B.n378 585
R564 B.n380 B.n95 585
R565 B.n382 B.n381 585
R566 B.n383 B.n94 585
R567 B.n385 B.n384 585
R568 B.n386 B.n93 585
R569 B.n388 B.n387 585
R570 B.n389 B.n92 585
R571 B.n391 B.n390 585
R572 B.n392 B.n91 585
R573 B.n394 B.n393 585
R574 B.n395 B.n90 585
R575 B.n397 B.n396 585
R576 B.n398 B.n89 585
R577 B.n400 B.n399 585
R578 B.n401 B.n88 585
R579 B.n403 B.n402 585
R580 B.n404 B.n87 585
R581 B.n406 B.n405 585
R582 B.n407 B.n86 585
R583 B.n409 B.n408 585
R584 B.n410 B.n85 585
R585 B.n412 B.n411 585
R586 B.n413 B.n84 585
R587 B.n415 B.n414 585
R588 B.n416 B.n83 585
R589 B.n418 B.n417 585
R590 B.n419 B.n82 585
R591 B.n421 B.n420 585
R592 B.n422 B.n81 585
R593 B.n424 B.n423 585
R594 B.n425 B.n80 585
R595 B.n427 B.n426 585
R596 B.n428 B.n79 585
R597 B.n430 B.n429 585
R598 B.n431 B.n78 585
R599 B.n433 B.n432 585
R600 B.n434 B.n77 585
R601 B.n436 B.n435 585
R602 B.n437 B.n76 585
R603 B.n439 B.n438 585
R604 B.n440 B.n75 585
R605 B.n442 B.n441 585
R606 B.n443 B.n74 585
R607 B.n445 B.n444 585
R608 B.n446 B.n73 585
R609 B.n448 B.n447 585
R610 B.n449 B.n72 585
R611 B.n451 B.n450 585
R612 B.n452 B.n71 585
R613 B.n454 B.n453 585
R614 B.n455 B.n70 585
R615 B.n457 B.n456 585
R616 B.n458 B.n69 585
R617 B.n460 B.n459 585
R618 B.n461 B.n68 585
R619 B.n463 B.n462 585
R620 B.n464 B.n67 585
R621 B.n466 B.n465 585
R622 B.n467 B.n66 585
R623 B.n469 B.n468 585
R624 B.n470 B.n65 585
R625 B.n472 B.n471 585
R626 B.n473 B.n64 585
R627 B.n475 B.n474 585
R628 B.n476 B.n63 585
R629 B.n478 B.n477 585
R630 B.n479 B.n62 585
R631 B.n481 B.n480 585
R632 B.n482 B.n61 585
R633 B.n484 B.n483 585
R634 B.n485 B.n60 585
R635 B.n487 B.n486 585
R636 B.n488 B.n59 585
R637 B.n490 B.n489 585
R638 B.n566 B.n29 585
R639 B.n565 B.n564 585
R640 B.n563 B.n30 585
R641 B.n562 B.n561 585
R642 B.n560 B.n31 585
R643 B.n559 B.n558 585
R644 B.n557 B.n32 585
R645 B.n556 B.n555 585
R646 B.n554 B.n33 585
R647 B.n553 B.n552 585
R648 B.n551 B.n34 585
R649 B.n550 B.n549 585
R650 B.n548 B.n35 585
R651 B.n547 B.n546 585
R652 B.n545 B.n36 585
R653 B.n544 B.n543 585
R654 B.n542 B.n37 585
R655 B.n541 B.n540 585
R656 B.n539 B.n38 585
R657 B.n538 B.n537 585
R658 B.n535 B.n39 585
R659 B.n534 B.n533 585
R660 B.n532 B.n42 585
R661 B.n531 B.n530 585
R662 B.n529 B.n43 585
R663 B.n528 B.n527 585
R664 B.n526 B.n44 585
R665 B.n525 B.n524 585
R666 B.n523 B.n45 585
R667 B.n522 B.n521 585
R668 B.n520 B.n519 585
R669 B.n518 B.n49 585
R670 B.n517 B.n516 585
R671 B.n515 B.n50 585
R672 B.n514 B.n513 585
R673 B.n512 B.n51 585
R674 B.n511 B.n510 585
R675 B.n509 B.n52 585
R676 B.n508 B.n507 585
R677 B.n506 B.n53 585
R678 B.n505 B.n504 585
R679 B.n503 B.n54 585
R680 B.n502 B.n501 585
R681 B.n500 B.n55 585
R682 B.n499 B.n498 585
R683 B.n497 B.n56 585
R684 B.n496 B.n495 585
R685 B.n494 B.n57 585
R686 B.n493 B.n492 585
R687 B.n491 B.n58 585
R688 B.n568 B.n567 585
R689 B.n569 B.n28 585
R690 B.n571 B.n570 585
R691 B.n572 B.n27 585
R692 B.n574 B.n573 585
R693 B.n575 B.n26 585
R694 B.n577 B.n576 585
R695 B.n578 B.n25 585
R696 B.n580 B.n579 585
R697 B.n581 B.n24 585
R698 B.n583 B.n582 585
R699 B.n584 B.n23 585
R700 B.n586 B.n585 585
R701 B.n587 B.n22 585
R702 B.n589 B.n588 585
R703 B.n590 B.n21 585
R704 B.n592 B.n591 585
R705 B.n593 B.n20 585
R706 B.n595 B.n594 585
R707 B.n596 B.n19 585
R708 B.n598 B.n597 585
R709 B.n599 B.n18 585
R710 B.n601 B.n600 585
R711 B.n602 B.n17 585
R712 B.n604 B.n603 585
R713 B.n605 B.n16 585
R714 B.n607 B.n606 585
R715 B.n608 B.n15 585
R716 B.n610 B.n609 585
R717 B.n611 B.n14 585
R718 B.n613 B.n612 585
R719 B.n614 B.n13 585
R720 B.n616 B.n615 585
R721 B.n617 B.n12 585
R722 B.n619 B.n618 585
R723 B.n620 B.n11 585
R724 B.n622 B.n621 585
R725 B.n623 B.n10 585
R726 B.n625 B.n624 585
R727 B.n626 B.n9 585
R728 B.n628 B.n627 585
R729 B.n629 B.n8 585
R730 B.n631 B.n630 585
R731 B.n632 B.n7 585
R732 B.n634 B.n633 585
R733 B.n635 B.n6 585
R734 B.n637 B.n636 585
R735 B.n638 B.n5 585
R736 B.n640 B.n639 585
R737 B.n641 B.n4 585
R738 B.n643 B.n642 585
R739 B.n644 B.n3 585
R740 B.n646 B.n645 585
R741 B.n647 B.n0 585
R742 B.n2 B.n1 585
R743 B.n168 B.n167 585
R744 B.n169 B.n166 585
R745 B.n171 B.n170 585
R746 B.n172 B.n165 585
R747 B.n174 B.n173 585
R748 B.n175 B.n164 585
R749 B.n177 B.n176 585
R750 B.n178 B.n163 585
R751 B.n180 B.n179 585
R752 B.n181 B.n162 585
R753 B.n183 B.n182 585
R754 B.n184 B.n161 585
R755 B.n186 B.n185 585
R756 B.n187 B.n160 585
R757 B.n189 B.n188 585
R758 B.n190 B.n159 585
R759 B.n192 B.n191 585
R760 B.n193 B.n158 585
R761 B.n195 B.n194 585
R762 B.n196 B.n157 585
R763 B.n198 B.n197 585
R764 B.n199 B.n156 585
R765 B.n201 B.n200 585
R766 B.n202 B.n155 585
R767 B.n204 B.n203 585
R768 B.n205 B.n154 585
R769 B.n207 B.n206 585
R770 B.n208 B.n153 585
R771 B.n210 B.n209 585
R772 B.n211 B.n152 585
R773 B.n213 B.n212 585
R774 B.n214 B.n151 585
R775 B.n216 B.n215 585
R776 B.n217 B.n150 585
R777 B.n219 B.n218 585
R778 B.n220 B.n149 585
R779 B.n222 B.n221 585
R780 B.n223 B.n148 585
R781 B.n225 B.n224 585
R782 B.n226 B.n147 585
R783 B.n228 B.n227 585
R784 B.n229 B.n146 585
R785 B.n231 B.n230 585
R786 B.n232 B.n145 585
R787 B.n234 B.n233 585
R788 B.n235 B.n144 585
R789 B.n237 B.n236 585
R790 B.n238 B.n143 585
R791 B.n240 B.n239 585
R792 B.n241 B.n142 585
R793 B.n243 B.n242 585
R794 B.n244 B.n141 585
R795 B.n246 B.n245 585
R796 B.n247 B.n246 487.695
R797 B.n324 B.n113 487.695
R798 B.n491 B.n490 487.695
R799 B.n568 B.n29 487.695
R800 B.n124 B.t4 322.308
R801 B.n46 B.t8 322.308
R802 B.n275 B.t1 322.308
R803 B.n40 B.t11 322.308
R804 B.n649 B.n648 256.663
R805 B.n125 B.t5 245.702
R806 B.n47 B.t7 245.702
R807 B.n276 B.t2 245.702
R808 B.n41 B.t10 245.702
R809 B.n275 B.t0 240.288
R810 B.n124 B.t3 240.288
R811 B.n46 B.t6 240.288
R812 B.n40 B.t9 240.288
R813 B.n648 B.n647 235.042
R814 B.n648 B.n2 235.042
R815 B.n248 B.n247 163.367
R816 B.n248 B.n139 163.367
R817 B.n252 B.n139 163.367
R818 B.n253 B.n252 163.367
R819 B.n254 B.n253 163.367
R820 B.n254 B.n137 163.367
R821 B.n258 B.n137 163.367
R822 B.n259 B.n258 163.367
R823 B.n260 B.n259 163.367
R824 B.n260 B.n135 163.367
R825 B.n264 B.n135 163.367
R826 B.n265 B.n264 163.367
R827 B.n266 B.n265 163.367
R828 B.n266 B.n133 163.367
R829 B.n270 B.n133 163.367
R830 B.n271 B.n270 163.367
R831 B.n272 B.n271 163.367
R832 B.n272 B.n131 163.367
R833 B.n279 B.n131 163.367
R834 B.n280 B.n279 163.367
R835 B.n281 B.n280 163.367
R836 B.n281 B.n129 163.367
R837 B.n285 B.n129 163.367
R838 B.n286 B.n285 163.367
R839 B.n287 B.n286 163.367
R840 B.n287 B.n127 163.367
R841 B.n291 B.n127 163.367
R842 B.n292 B.n291 163.367
R843 B.n293 B.n292 163.367
R844 B.n293 B.n123 163.367
R845 B.n298 B.n123 163.367
R846 B.n299 B.n298 163.367
R847 B.n300 B.n299 163.367
R848 B.n300 B.n121 163.367
R849 B.n304 B.n121 163.367
R850 B.n305 B.n304 163.367
R851 B.n306 B.n305 163.367
R852 B.n306 B.n119 163.367
R853 B.n310 B.n119 163.367
R854 B.n311 B.n310 163.367
R855 B.n312 B.n311 163.367
R856 B.n312 B.n117 163.367
R857 B.n316 B.n117 163.367
R858 B.n317 B.n316 163.367
R859 B.n318 B.n317 163.367
R860 B.n318 B.n115 163.367
R861 B.n322 B.n115 163.367
R862 B.n323 B.n322 163.367
R863 B.n324 B.n323 163.367
R864 B.n490 B.n59 163.367
R865 B.n486 B.n59 163.367
R866 B.n486 B.n485 163.367
R867 B.n485 B.n484 163.367
R868 B.n484 B.n61 163.367
R869 B.n480 B.n61 163.367
R870 B.n480 B.n479 163.367
R871 B.n479 B.n478 163.367
R872 B.n478 B.n63 163.367
R873 B.n474 B.n63 163.367
R874 B.n474 B.n473 163.367
R875 B.n473 B.n472 163.367
R876 B.n472 B.n65 163.367
R877 B.n468 B.n65 163.367
R878 B.n468 B.n467 163.367
R879 B.n467 B.n466 163.367
R880 B.n466 B.n67 163.367
R881 B.n462 B.n67 163.367
R882 B.n462 B.n461 163.367
R883 B.n461 B.n460 163.367
R884 B.n460 B.n69 163.367
R885 B.n456 B.n69 163.367
R886 B.n456 B.n455 163.367
R887 B.n455 B.n454 163.367
R888 B.n454 B.n71 163.367
R889 B.n450 B.n71 163.367
R890 B.n450 B.n449 163.367
R891 B.n449 B.n448 163.367
R892 B.n448 B.n73 163.367
R893 B.n444 B.n73 163.367
R894 B.n444 B.n443 163.367
R895 B.n443 B.n442 163.367
R896 B.n442 B.n75 163.367
R897 B.n438 B.n75 163.367
R898 B.n438 B.n437 163.367
R899 B.n437 B.n436 163.367
R900 B.n436 B.n77 163.367
R901 B.n432 B.n77 163.367
R902 B.n432 B.n431 163.367
R903 B.n431 B.n430 163.367
R904 B.n430 B.n79 163.367
R905 B.n426 B.n79 163.367
R906 B.n426 B.n425 163.367
R907 B.n425 B.n424 163.367
R908 B.n424 B.n81 163.367
R909 B.n420 B.n81 163.367
R910 B.n420 B.n419 163.367
R911 B.n419 B.n418 163.367
R912 B.n418 B.n83 163.367
R913 B.n414 B.n83 163.367
R914 B.n414 B.n413 163.367
R915 B.n413 B.n412 163.367
R916 B.n412 B.n85 163.367
R917 B.n408 B.n85 163.367
R918 B.n408 B.n407 163.367
R919 B.n407 B.n406 163.367
R920 B.n406 B.n87 163.367
R921 B.n402 B.n87 163.367
R922 B.n402 B.n401 163.367
R923 B.n401 B.n400 163.367
R924 B.n400 B.n89 163.367
R925 B.n396 B.n89 163.367
R926 B.n396 B.n395 163.367
R927 B.n395 B.n394 163.367
R928 B.n394 B.n91 163.367
R929 B.n390 B.n91 163.367
R930 B.n390 B.n389 163.367
R931 B.n389 B.n388 163.367
R932 B.n388 B.n93 163.367
R933 B.n384 B.n93 163.367
R934 B.n384 B.n383 163.367
R935 B.n383 B.n382 163.367
R936 B.n382 B.n95 163.367
R937 B.n378 B.n95 163.367
R938 B.n378 B.n377 163.367
R939 B.n377 B.n376 163.367
R940 B.n376 B.n97 163.367
R941 B.n372 B.n97 163.367
R942 B.n372 B.n371 163.367
R943 B.n371 B.n370 163.367
R944 B.n370 B.n99 163.367
R945 B.n366 B.n99 163.367
R946 B.n366 B.n365 163.367
R947 B.n365 B.n364 163.367
R948 B.n364 B.n101 163.367
R949 B.n360 B.n101 163.367
R950 B.n360 B.n359 163.367
R951 B.n359 B.n358 163.367
R952 B.n358 B.n103 163.367
R953 B.n354 B.n103 163.367
R954 B.n354 B.n353 163.367
R955 B.n353 B.n352 163.367
R956 B.n352 B.n105 163.367
R957 B.n348 B.n105 163.367
R958 B.n348 B.n347 163.367
R959 B.n347 B.n346 163.367
R960 B.n346 B.n107 163.367
R961 B.n342 B.n107 163.367
R962 B.n342 B.n341 163.367
R963 B.n341 B.n340 163.367
R964 B.n340 B.n109 163.367
R965 B.n336 B.n109 163.367
R966 B.n336 B.n335 163.367
R967 B.n335 B.n334 163.367
R968 B.n334 B.n111 163.367
R969 B.n330 B.n111 163.367
R970 B.n330 B.n329 163.367
R971 B.n329 B.n328 163.367
R972 B.n328 B.n113 163.367
R973 B.n564 B.n29 163.367
R974 B.n564 B.n563 163.367
R975 B.n563 B.n562 163.367
R976 B.n562 B.n31 163.367
R977 B.n558 B.n31 163.367
R978 B.n558 B.n557 163.367
R979 B.n557 B.n556 163.367
R980 B.n556 B.n33 163.367
R981 B.n552 B.n33 163.367
R982 B.n552 B.n551 163.367
R983 B.n551 B.n550 163.367
R984 B.n550 B.n35 163.367
R985 B.n546 B.n35 163.367
R986 B.n546 B.n545 163.367
R987 B.n545 B.n544 163.367
R988 B.n544 B.n37 163.367
R989 B.n540 B.n37 163.367
R990 B.n540 B.n539 163.367
R991 B.n539 B.n538 163.367
R992 B.n538 B.n39 163.367
R993 B.n533 B.n39 163.367
R994 B.n533 B.n532 163.367
R995 B.n532 B.n531 163.367
R996 B.n531 B.n43 163.367
R997 B.n527 B.n43 163.367
R998 B.n527 B.n526 163.367
R999 B.n526 B.n525 163.367
R1000 B.n525 B.n45 163.367
R1001 B.n521 B.n45 163.367
R1002 B.n521 B.n520 163.367
R1003 B.n520 B.n49 163.367
R1004 B.n516 B.n49 163.367
R1005 B.n516 B.n515 163.367
R1006 B.n515 B.n514 163.367
R1007 B.n514 B.n51 163.367
R1008 B.n510 B.n51 163.367
R1009 B.n510 B.n509 163.367
R1010 B.n509 B.n508 163.367
R1011 B.n508 B.n53 163.367
R1012 B.n504 B.n53 163.367
R1013 B.n504 B.n503 163.367
R1014 B.n503 B.n502 163.367
R1015 B.n502 B.n55 163.367
R1016 B.n498 B.n55 163.367
R1017 B.n498 B.n497 163.367
R1018 B.n497 B.n496 163.367
R1019 B.n496 B.n57 163.367
R1020 B.n492 B.n57 163.367
R1021 B.n492 B.n491 163.367
R1022 B.n569 B.n568 163.367
R1023 B.n570 B.n569 163.367
R1024 B.n570 B.n27 163.367
R1025 B.n574 B.n27 163.367
R1026 B.n575 B.n574 163.367
R1027 B.n576 B.n575 163.367
R1028 B.n576 B.n25 163.367
R1029 B.n580 B.n25 163.367
R1030 B.n581 B.n580 163.367
R1031 B.n582 B.n581 163.367
R1032 B.n582 B.n23 163.367
R1033 B.n586 B.n23 163.367
R1034 B.n587 B.n586 163.367
R1035 B.n588 B.n587 163.367
R1036 B.n588 B.n21 163.367
R1037 B.n592 B.n21 163.367
R1038 B.n593 B.n592 163.367
R1039 B.n594 B.n593 163.367
R1040 B.n594 B.n19 163.367
R1041 B.n598 B.n19 163.367
R1042 B.n599 B.n598 163.367
R1043 B.n600 B.n599 163.367
R1044 B.n600 B.n17 163.367
R1045 B.n604 B.n17 163.367
R1046 B.n605 B.n604 163.367
R1047 B.n606 B.n605 163.367
R1048 B.n606 B.n15 163.367
R1049 B.n610 B.n15 163.367
R1050 B.n611 B.n610 163.367
R1051 B.n612 B.n611 163.367
R1052 B.n612 B.n13 163.367
R1053 B.n616 B.n13 163.367
R1054 B.n617 B.n616 163.367
R1055 B.n618 B.n617 163.367
R1056 B.n618 B.n11 163.367
R1057 B.n622 B.n11 163.367
R1058 B.n623 B.n622 163.367
R1059 B.n624 B.n623 163.367
R1060 B.n624 B.n9 163.367
R1061 B.n628 B.n9 163.367
R1062 B.n629 B.n628 163.367
R1063 B.n630 B.n629 163.367
R1064 B.n630 B.n7 163.367
R1065 B.n634 B.n7 163.367
R1066 B.n635 B.n634 163.367
R1067 B.n636 B.n635 163.367
R1068 B.n636 B.n5 163.367
R1069 B.n640 B.n5 163.367
R1070 B.n641 B.n640 163.367
R1071 B.n642 B.n641 163.367
R1072 B.n642 B.n3 163.367
R1073 B.n646 B.n3 163.367
R1074 B.n647 B.n646 163.367
R1075 B.n168 B.n2 163.367
R1076 B.n169 B.n168 163.367
R1077 B.n170 B.n169 163.367
R1078 B.n170 B.n165 163.367
R1079 B.n174 B.n165 163.367
R1080 B.n175 B.n174 163.367
R1081 B.n176 B.n175 163.367
R1082 B.n176 B.n163 163.367
R1083 B.n180 B.n163 163.367
R1084 B.n181 B.n180 163.367
R1085 B.n182 B.n181 163.367
R1086 B.n182 B.n161 163.367
R1087 B.n186 B.n161 163.367
R1088 B.n187 B.n186 163.367
R1089 B.n188 B.n187 163.367
R1090 B.n188 B.n159 163.367
R1091 B.n192 B.n159 163.367
R1092 B.n193 B.n192 163.367
R1093 B.n194 B.n193 163.367
R1094 B.n194 B.n157 163.367
R1095 B.n198 B.n157 163.367
R1096 B.n199 B.n198 163.367
R1097 B.n200 B.n199 163.367
R1098 B.n200 B.n155 163.367
R1099 B.n204 B.n155 163.367
R1100 B.n205 B.n204 163.367
R1101 B.n206 B.n205 163.367
R1102 B.n206 B.n153 163.367
R1103 B.n210 B.n153 163.367
R1104 B.n211 B.n210 163.367
R1105 B.n212 B.n211 163.367
R1106 B.n212 B.n151 163.367
R1107 B.n216 B.n151 163.367
R1108 B.n217 B.n216 163.367
R1109 B.n218 B.n217 163.367
R1110 B.n218 B.n149 163.367
R1111 B.n222 B.n149 163.367
R1112 B.n223 B.n222 163.367
R1113 B.n224 B.n223 163.367
R1114 B.n224 B.n147 163.367
R1115 B.n228 B.n147 163.367
R1116 B.n229 B.n228 163.367
R1117 B.n230 B.n229 163.367
R1118 B.n230 B.n145 163.367
R1119 B.n234 B.n145 163.367
R1120 B.n235 B.n234 163.367
R1121 B.n236 B.n235 163.367
R1122 B.n236 B.n143 163.367
R1123 B.n240 B.n143 163.367
R1124 B.n241 B.n240 163.367
R1125 B.n242 B.n241 163.367
R1126 B.n242 B.n141 163.367
R1127 B.n246 B.n141 163.367
R1128 B.n276 B.n275 76.6066
R1129 B.n125 B.n124 76.6066
R1130 B.n47 B.n46 76.6066
R1131 B.n41 B.n40 76.6066
R1132 B.n277 B.n276 59.5399
R1133 B.n295 B.n125 59.5399
R1134 B.n48 B.n47 59.5399
R1135 B.n536 B.n41 59.5399
R1136 B.n567 B.n566 31.6883
R1137 B.n489 B.n58 31.6883
R1138 B.n326 B.n325 31.6883
R1139 B.n245 B.n140 31.6883
R1140 B B.n649 18.0485
R1141 B.n567 B.n28 10.6151
R1142 B.n571 B.n28 10.6151
R1143 B.n572 B.n571 10.6151
R1144 B.n573 B.n572 10.6151
R1145 B.n573 B.n26 10.6151
R1146 B.n577 B.n26 10.6151
R1147 B.n578 B.n577 10.6151
R1148 B.n579 B.n578 10.6151
R1149 B.n579 B.n24 10.6151
R1150 B.n583 B.n24 10.6151
R1151 B.n584 B.n583 10.6151
R1152 B.n585 B.n584 10.6151
R1153 B.n585 B.n22 10.6151
R1154 B.n589 B.n22 10.6151
R1155 B.n590 B.n589 10.6151
R1156 B.n591 B.n590 10.6151
R1157 B.n591 B.n20 10.6151
R1158 B.n595 B.n20 10.6151
R1159 B.n596 B.n595 10.6151
R1160 B.n597 B.n596 10.6151
R1161 B.n597 B.n18 10.6151
R1162 B.n601 B.n18 10.6151
R1163 B.n602 B.n601 10.6151
R1164 B.n603 B.n602 10.6151
R1165 B.n603 B.n16 10.6151
R1166 B.n607 B.n16 10.6151
R1167 B.n608 B.n607 10.6151
R1168 B.n609 B.n608 10.6151
R1169 B.n609 B.n14 10.6151
R1170 B.n613 B.n14 10.6151
R1171 B.n614 B.n613 10.6151
R1172 B.n615 B.n614 10.6151
R1173 B.n615 B.n12 10.6151
R1174 B.n619 B.n12 10.6151
R1175 B.n620 B.n619 10.6151
R1176 B.n621 B.n620 10.6151
R1177 B.n621 B.n10 10.6151
R1178 B.n625 B.n10 10.6151
R1179 B.n626 B.n625 10.6151
R1180 B.n627 B.n626 10.6151
R1181 B.n627 B.n8 10.6151
R1182 B.n631 B.n8 10.6151
R1183 B.n632 B.n631 10.6151
R1184 B.n633 B.n632 10.6151
R1185 B.n633 B.n6 10.6151
R1186 B.n637 B.n6 10.6151
R1187 B.n638 B.n637 10.6151
R1188 B.n639 B.n638 10.6151
R1189 B.n639 B.n4 10.6151
R1190 B.n643 B.n4 10.6151
R1191 B.n644 B.n643 10.6151
R1192 B.n645 B.n644 10.6151
R1193 B.n645 B.n0 10.6151
R1194 B.n566 B.n565 10.6151
R1195 B.n565 B.n30 10.6151
R1196 B.n561 B.n30 10.6151
R1197 B.n561 B.n560 10.6151
R1198 B.n560 B.n559 10.6151
R1199 B.n559 B.n32 10.6151
R1200 B.n555 B.n32 10.6151
R1201 B.n555 B.n554 10.6151
R1202 B.n554 B.n553 10.6151
R1203 B.n553 B.n34 10.6151
R1204 B.n549 B.n34 10.6151
R1205 B.n549 B.n548 10.6151
R1206 B.n548 B.n547 10.6151
R1207 B.n547 B.n36 10.6151
R1208 B.n543 B.n36 10.6151
R1209 B.n543 B.n542 10.6151
R1210 B.n542 B.n541 10.6151
R1211 B.n541 B.n38 10.6151
R1212 B.n537 B.n38 10.6151
R1213 B.n535 B.n534 10.6151
R1214 B.n534 B.n42 10.6151
R1215 B.n530 B.n42 10.6151
R1216 B.n530 B.n529 10.6151
R1217 B.n529 B.n528 10.6151
R1218 B.n528 B.n44 10.6151
R1219 B.n524 B.n44 10.6151
R1220 B.n524 B.n523 10.6151
R1221 B.n523 B.n522 10.6151
R1222 B.n519 B.n518 10.6151
R1223 B.n518 B.n517 10.6151
R1224 B.n517 B.n50 10.6151
R1225 B.n513 B.n50 10.6151
R1226 B.n513 B.n512 10.6151
R1227 B.n512 B.n511 10.6151
R1228 B.n511 B.n52 10.6151
R1229 B.n507 B.n52 10.6151
R1230 B.n507 B.n506 10.6151
R1231 B.n506 B.n505 10.6151
R1232 B.n505 B.n54 10.6151
R1233 B.n501 B.n54 10.6151
R1234 B.n501 B.n500 10.6151
R1235 B.n500 B.n499 10.6151
R1236 B.n499 B.n56 10.6151
R1237 B.n495 B.n56 10.6151
R1238 B.n495 B.n494 10.6151
R1239 B.n494 B.n493 10.6151
R1240 B.n493 B.n58 10.6151
R1241 B.n489 B.n488 10.6151
R1242 B.n488 B.n487 10.6151
R1243 B.n487 B.n60 10.6151
R1244 B.n483 B.n60 10.6151
R1245 B.n483 B.n482 10.6151
R1246 B.n482 B.n481 10.6151
R1247 B.n481 B.n62 10.6151
R1248 B.n477 B.n62 10.6151
R1249 B.n477 B.n476 10.6151
R1250 B.n476 B.n475 10.6151
R1251 B.n475 B.n64 10.6151
R1252 B.n471 B.n64 10.6151
R1253 B.n471 B.n470 10.6151
R1254 B.n470 B.n469 10.6151
R1255 B.n469 B.n66 10.6151
R1256 B.n465 B.n66 10.6151
R1257 B.n465 B.n464 10.6151
R1258 B.n464 B.n463 10.6151
R1259 B.n463 B.n68 10.6151
R1260 B.n459 B.n68 10.6151
R1261 B.n459 B.n458 10.6151
R1262 B.n458 B.n457 10.6151
R1263 B.n457 B.n70 10.6151
R1264 B.n453 B.n70 10.6151
R1265 B.n453 B.n452 10.6151
R1266 B.n452 B.n451 10.6151
R1267 B.n451 B.n72 10.6151
R1268 B.n447 B.n72 10.6151
R1269 B.n447 B.n446 10.6151
R1270 B.n446 B.n445 10.6151
R1271 B.n445 B.n74 10.6151
R1272 B.n441 B.n74 10.6151
R1273 B.n441 B.n440 10.6151
R1274 B.n440 B.n439 10.6151
R1275 B.n439 B.n76 10.6151
R1276 B.n435 B.n76 10.6151
R1277 B.n435 B.n434 10.6151
R1278 B.n434 B.n433 10.6151
R1279 B.n433 B.n78 10.6151
R1280 B.n429 B.n78 10.6151
R1281 B.n429 B.n428 10.6151
R1282 B.n428 B.n427 10.6151
R1283 B.n427 B.n80 10.6151
R1284 B.n423 B.n80 10.6151
R1285 B.n423 B.n422 10.6151
R1286 B.n422 B.n421 10.6151
R1287 B.n421 B.n82 10.6151
R1288 B.n417 B.n82 10.6151
R1289 B.n417 B.n416 10.6151
R1290 B.n416 B.n415 10.6151
R1291 B.n415 B.n84 10.6151
R1292 B.n411 B.n84 10.6151
R1293 B.n411 B.n410 10.6151
R1294 B.n410 B.n409 10.6151
R1295 B.n409 B.n86 10.6151
R1296 B.n405 B.n86 10.6151
R1297 B.n405 B.n404 10.6151
R1298 B.n404 B.n403 10.6151
R1299 B.n403 B.n88 10.6151
R1300 B.n399 B.n88 10.6151
R1301 B.n399 B.n398 10.6151
R1302 B.n398 B.n397 10.6151
R1303 B.n397 B.n90 10.6151
R1304 B.n393 B.n90 10.6151
R1305 B.n393 B.n392 10.6151
R1306 B.n392 B.n391 10.6151
R1307 B.n391 B.n92 10.6151
R1308 B.n387 B.n92 10.6151
R1309 B.n387 B.n386 10.6151
R1310 B.n386 B.n385 10.6151
R1311 B.n385 B.n94 10.6151
R1312 B.n381 B.n94 10.6151
R1313 B.n381 B.n380 10.6151
R1314 B.n380 B.n379 10.6151
R1315 B.n379 B.n96 10.6151
R1316 B.n375 B.n96 10.6151
R1317 B.n375 B.n374 10.6151
R1318 B.n374 B.n373 10.6151
R1319 B.n373 B.n98 10.6151
R1320 B.n369 B.n98 10.6151
R1321 B.n369 B.n368 10.6151
R1322 B.n368 B.n367 10.6151
R1323 B.n367 B.n100 10.6151
R1324 B.n363 B.n100 10.6151
R1325 B.n363 B.n362 10.6151
R1326 B.n362 B.n361 10.6151
R1327 B.n361 B.n102 10.6151
R1328 B.n357 B.n102 10.6151
R1329 B.n357 B.n356 10.6151
R1330 B.n356 B.n355 10.6151
R1331 B.n355 B.n104 10.6151
R1332 B.n351 B.n104 10.6151
R1333 B.n351 B.n350 10.6151
R1334 B.n350 B.n349 10.6151
R1335 B.n349 B.n106 10.6151
R1336 B.n345 B.n106 10.6151
R1337 B.n345 B.n344 10.6151
R1338 B.n344 B.n343 10.6151
R1339 B.n343 B.n108 10.6151
R1340 B.n339 B.n108 10.6151
R1341 B.n339 B.n338 10.6151
R1342 B.n338 B.n337 10.6151
R1343 B.n337 B.n110 10.6151
R1344 B.n333 B.n110 10.6151
R1345 B.n333 B.n332 10.6151
R1346 B.n332 B.n331 10.6151
R1347 B.n331 B.n112 10.6151
R1348 B.n327 B.n112 10.6151
R1349 B.n327 B.n326 10.6151
R1350 B.n167 B.n1 10.6151
R1351 B.n167 B.n166 10.6151
R1352 B.n171 B.n166 10.6151
R1353 B.n172 B.n171 10.6151
R1354 B.n173 B.n172 10.6151
R1355 B.n173 B.n164 10.6151
R1356 B.n177 B.n164 10.6151
R1357 B.n178 B.n177 10.6151
R1358 B.n179 B.n178 10.6151
R1359 B.n179 B.n162 10.6151
R1360 B.n183 B.n162 10.6151
R1361 B.n184 B.n183 10.6151
R1362 B.n185 B.n184 10.6151
R1363 B.n185 B.n160 10.6151
R1364 B.n189 B.n160 10.6151
R1365 B.n190 B.n189 10.6151
R1366 B.n191 B.n190 10.6151
R1367 B.n191 B.n158 10.6151
R1368 B.n195 B.n158 10.6151
R1369 B.n196 B.n195 10.6151
R1370 B.n197 B.n196 10.6151
R1371 B.n197 B.n156 10.6151
R1372 B.n201 B.n156 10.6151
R1373 B.n202 B.n201 10.6151
R1374 B.n203 B.n202 10.6151
R1375 B.n203 B.n154 10.6151
R1376 B.n207 B.n154 10.6151
R1377 B.n208 B.n207 10.6151
R1378 B.n209 B.n208 10.6151
R1379 B.n209 B.n152 10.6151
R1380 B.n213 B.n152 10.6151
R1381 B.n214 B.n213 10.6151
R1382 B.n215 B.n214 10.6151
R1383 B.n215 B.n150 10.6151
R1384 B.n219 B.n150 10.6151
R1385 B.n220 B.n219 10.6151
R1386 B.n221 B.n220 10.6151
R1387 B.n221 B.n148 10.6151
R1388 B.n225 B.n148 10.6151
R1389 B.n226 B.n225 10.6151
R1390 B.n227 B.n226 10.6151
R1391 B.n227 B.n146 10.6151
R1392 B.n231 B.n146 10.6151
R1393 B.n232 B.n231 10.6151
R1394 B.n233 B.n232 10.6151
R1395 B.n233 B.n144 10.6151
R1396 B.n237 B.n144 10.6151
R1397 B.n238 B.n237 10.6151
R1398 B.n239 B.n238 10.6151
R1399 B.n239 B.n142 10.6151
R1400 B.n243 B.n142 10.6151
R1401 B.n244 B.n243 10.6151
R1402 B.n245 B.n244 10.6151
R1403 B.n249 B.n140 10.6151
R1404 B.n250 B.n249 10.6151
R1405 B.n251 B.n250 10.6151
R1406 B.n251 B.n138 10.6151
R1407 B.n255 B.n138 10.6151
R1408 B.n256 B.n255 10.6151
R1409 B.n257 B.n256 10.6151
R1410 B.n257 B.n136 10.6151
R1411 B.n261 B.n136 10.6151
R1412 B.n262 B.n261 10.6151
R1413 B.n263 B.n262 10.6151
R1414 B.n263 B.n134 10.6151
R1415 B.n267 B.n134 10.6151
R1416 B.n268 B.n267 10.6151
R1417 B.n269 B.n268 10.6151
R1418 B.n269 B.n132 10.6151
R1419 B.n273 B.n132 10.6151
R1420 B.n274 B.n273 10.6151
R1421 B.n278 B.n274 10.6151
R1422 B.n282 B.n130 10.6151
R1423 B.n283 B.n282 10.6151
R1424 B.n284 B.n283 10.6151
R1425 B.n284 B.n128 10.6151
R1426 B.n288 B.n128 10.6151
R1427 B.n289 B.n288 10.6151
R1428 B.n290 B.n289 10.6151
R1429 B.n290 B.n126 10.6151
R1430 B.n294 B.n126 10.6151
R1431 B.n297 B.n296 10.6151
R1432 B.n297 B.n122 10.6151
R1433 B.n301 B.n122 10.6151
R1434 B.n302 B.n301 10.6151
R1435 B.n303 B.n302 10.6151
R1436 B.n303 B.n120 10.6151
R1437 B.n307 B.n120 10.6151
R1438 B.n308 B.n307 10.6151
R1439 B.n309 B.n308 10.6151
R1440 B.n309 B.n118 10.6151
R1441 B.n313 B.n118 10.6151
R1442 B.n314 B.n313 10.6151
R1443 B.n315 B.n314 10.6151
R1444 B.n315 B.n116 10.6151
R1445 B.n319 B.n116 10.6151
R1446 B.n320 B.n319 10.6151
R1447 B.n321 B.n320 10.6151
R1448 B.n321 B.n114 10.6151
R1449 B.n325 B.n114 10.6151
R1450 B.n537 B.n536 9.36635
R1451 B.n519 B.n48 9.36635
R1452 B.n278 B.n277 9.36635
R1453 B.n296 B.n295 9.36635
R1454 B.n649 B.n0 8.11757
R1455 B.n649 B.n1 8.11757
R1456 B.n536 B.n535 1.24928
R1457 B.n522 B.n48 1.24928
R1458 B.n277 B.n130 1.24928
R1459 B.n295 B.n294 1.24928
C0 VDD1 B 1.76768f
C1 VDD2 VP 0.548864f
C2 VDD1 w_n4130_n1902# 2.03796f
C3 VN VDD1 0.156158f
C4 VP VTAIL 3.98945f
C5 w_n4130_n1902# B 9.05092f
C6 VN B 1.32532f
C7 VDD2 VDD1 1.80505f
C8 VN w_n4130_n1902# 7.939229f
C9 VDD1 VTAIL 5.70745f
C10 VDD2 B 1.86639f
C11 VDD2 w_n4130_n1902# 2.15533f
C12 VDD2 VN 3.00884f
C13 VTAIL B 2.30326f
C14 w_n4130_n1902# VTAIL 2.06387f
C15 VN VTAIL 3.97525f
C16 VDD1 VP 3.39887f
C17 VP B 2.2266f
C18 VDD2 VTAIL 5.76718f
C19 VP w_n4130_n1902# 8.47593f
C20 VN VP 6.55973f
C21 VDD2 VSUBS 1.818936f
C22 VDD1 VSUBS 1.944514f
C23 VTAIL VSUBS 0.764497f
C24 VN VSUBS 6.64667f
C25 VP VSUBS 3.21266f
C26 B VSUBS 4.732686f
C27 w_n4130_n1902# VSUBS 98.57479f
C28 B.n0 VSUBS 0.00856f
C29 B.n1 VSUBS 0.00856f
C30 B.n2 VSUBS 0.012659f
C31 B.n3 VSUBS 0.009701f
C32 B.n4 VSUBS 0.009701f
C33 B.n5 VSUBS 0.009701f
C34 B.n6 VSUBS 0.009701f
C35 B.n7 VSUBS 0.009701f
C36 B.n8 VSUBS 0.009701f
C37 B.n9 VSUBS 0.009701f
C38 B.n10 VSUBS 0.009701f
C39 B.n11 VSUBS 0.009701f
C40 B.n12 VSUBS 0.009701f
C41 B.n13 VSUBS 0.009701f
C42 B.n14 VSUBS 0.009701f
C43 B.n15 VSUBS 0.009701f
C44 B.n16 VSUBS 0.009701f
C45 B.n17 VSUBS 0.009701f
C46 B.n18 VSUBS 0.009701f
C47 B.n19 VSUBS 0.009701f
C48 B.n20 VSUBS 0.009701f
C49 B.n21 VSUBS 0.009701f
C50 B.n22 VSUBS 0.009701f
C51 B.n23 VSUBS 0.009701f
C52 B.n24 VSUBS 0.009701f
C53 B.n25 VSUBS 0.009701f
C54 B.n26 VSUBS 0.009701f
C55 B.n27 VSUBS 0.009701f
C56 B.n28 VSUBS 0.009701f
C57 B.n29 VSUBS 0.023048f
C58 B.n30 VSUBS 0.009701f
C59 B.n31 VSUBS 0.009701f
C60 B.n32 VSUBS 0.009701f
C61 B.n33 VSUBS 0.009701f
C62 B.n34 VSUBS 0.009701f
C63 B.n35 VSUBS 0.009701f
C64 B.n36 VSUBS 0.009701f
C65 B.n37 VSUBS 0.009701f
C66 B.n38 VSUBS 0.009701f
C67 B.n39 VSUBS 0.009701f
C68 B.t10 VSUBS 0.093959f
C69 B.t11 VSUBS 0.134898f
C70 B.t9 VSUBS 1.13399f
C71 B.n40 VSUBS 0.226718f
C72 B.n41 VSUBS 0.186079f
C73 B.n42 VSUBS 0.009701f
C74 B.n43 VSUBS 0.009701f
C75 B.n44 VSUBS 0.009701f
C76 B.n45 VSUBS 0.009701f
C77 B.t7 VSUBS 0.093961f
C78 B.t8 VSUBS 0.134899f
C79 B.t6 VSUBS 1.13399f
C80 B.n46 VSUBS 0.226716f
C81 B.n47 VSUBS 0.186078f
C82 B.n48 VSUBS 0.022476f
C83 B.n49 VSUBS 0.009701f
C84 B.n50 VSUBS 0.009701f
C85 B.n51 VSUBS 0.009701f
C86 B.n52 VSUBS 0.009701f
C87 B.n53 VSUBS 0.009701f
C88 B.n54 VSUBS 0.009701f
C89 B.n55 VSUBS 0.009701f
C90 B.n56 VSUBS 0.009701f
C91 B.n57 VSUBS 0.009701f
C92 B.n58 VSUBS 0.023048f
C93 B.n59 VSUBS 0.009701f
C94 B.n60 VSUBS 0.009701f
C95 B.n61 VSUBS 0.009701f
C96 B.n62 VSUBS 0.009701f
C97 B.n63 VSUBS 0.009701f
C98 B.n64 VSUBS 0.009701f
C99 B.n65 VSUBS 0.009701f
C100 B.n66 VSUBS 0.009701f
C101 B.n67 VSUBS 0.009701f
C102 B.n68 VSUBS 0.009701f
C103 B.n69 VSUBS 0.009701f
C104 B.n70 VSUBS 0.009701f
C105 B.n71 VSUBS 0.009701f
C106 B.n72 VSUBS 0.009701f
C107 B.n73 VSUBS 0.009701f
C108 B.n74 VSUBS 0.009701f
C109 B.n75 VSUBS 0.009701f
C110 B.n76 VSUBS 0.009701f
C111 B.n77 VSUBS 0.009701f
C112 B.n78 VSUBS 0.009701f
C113 B.n79 VSUBS 0.009701f
C114 B.n80 VSUBS 0.009701f
C115 B.n81 VSUBS 0.009701f
C116 B.n82 VSUBS 0.009701f
C117 B.n83 VSUBS 0.009701f
C118 B.n84 VSUBS 0.009701f
C119 B.n85 VSUBS 0.009701f
C120 B.n86 VSUBS 0.009701f
C121 B.n87 VSUBS 0.009701f
C122 B.n88 VSUBS 0.009701f
C123 B.n89 VSUBS 0.009701f
C124 B.n90 VSUBS 0.009701f
C125 B.n91 VSUBS 0.009701f
C126 B.n92 VSUBS 0.009701f
C127 B.n93 VSUBS 0.009701f
C128 B.n94 VSUBS 0.009701f
C129 B.n95 VSUBS 0.009701f
C130 B.n96 VSUBS 0.009701f
C131 B.n97 VSUBS 0.009701f
C132 B.n98 VSUBS 0.009701f
C133 B.n99 VSUBS 0.009701f
C134 B.n100 VSUBS 0.009701f
C135 B.n101 VSUBS 0.009701f
C136 B.n102 VSUBS 0.009701f
C137 B.n103 VSUBS 0.009701f
C138 B.n104 VSUBS 0.009701f
C139 B.n105 VSUBS 0.009701f
C140 B.n106 VSUBS 0.009701f
C141 B.n107 VSUBS 0.009701f
C142 B.n108 VSUBS 0.009701f
C143 B.n109 VSUBS 0.009701f
C144 B.n110 VSUBS 0.009701f
C145 B.n111 VSUBS 0.009701f
C146 B.n112 VSUBS 0.009701f
C147 B.n113 VSUBS 0.021463f
C148 B.n114 VSUBS 0.009701f
C149 B.n115 VSUBS 0.009701f
C150 B.n116 VSUBS 0.009701f
C151 B.n117 VSUBS 0.009701f
C152 B.n118 VSUBS 0.009701f
C153 B.n119 VSUBS 0.009701f
C154 B.n120 VSUBS 0.009701f
C155 B.n121 VSUBS 0.009701f
C156 B.n122 VSUBS 0.009701f
C157 B.n123 VSUBS 0.009701f
C158 B.t5 VSUBS 0.093961f
C159 B.t4 VSUBS 0.134899f
C160 B.t3 VSUBS 1.13399f
C161 B.n124 VSUBS 0.226716f
C162 B.n125 VSUBS 0.186078f
C163 B.n126 VSUBS 0.009701f
C164 B.n127 VSUBS 0.009701f
C165 B.n128 VSUBS 0.009701f
C166 B.n129 VSUBS 0.009701f
C167 B.n130 VSUBS 0.005421f
C168 B.n131 VSUBS 0.009701f
C169 B.n132 VSUBS 0.009701f
C170 B.n133 VSUBS 0.009701f
C171 B.n134 VSUBS 0.009701f
C172 B.n135 VSUBS 0.009701f
C173 B.n136 VSUBS 0.009701f
C174 B.n137 VSUBS 0.009701f
C175 B.n138 VSUBS 0.009701f
C176 B.n139 VSUBS 0.009701f
C177 B.n140 VSUBS 0.023048f
C178 B.n141 VSUBS 0.009701f
C179 B.n142 VSUBS 0.009701f
C180 B.n143 VSUBS 0.009701f
C181 B.n144 VSUBS 0.009701f
C182 B.n145 VSUBS 0.009701f
C183 B.n146 VSUBS 0.009701f
C184 B.n147 VSUBS 0.009701f
C185 B.n148 VSUBS 0.009701f
C186 B.n149 VSUBS 0.009701f
C187 B.n150 VSUBS 0.009701f
C188 B.n151 VSUBS 0.009701f
C189 B.n152 VSUBS 0.009701f
C190 B.n153 VSUBS 0.009701f
C191 B.n154 VSUBS 0.009701f
C192 B.n155 VSUBS 0.009701f
C193 B.n156 VSUBS 0.009701f
C194 B.n157 VSUBS 0.009701f
C195 B.n158 VSUBS 0.009701f
C196 B.n159 VSUBS 0.009701f
C197 B.n160 VSUBS 0.009701f
C198 B.n161 VSUBS 0.009701f
C199 B.n162 VSUBS 0.009701f
C200 B.n163 VSUBS 0.009701f
C201 B.n164 VSUBS 0.009701f
C202 B.n165 VSUBS 0.009701f
C203 B.n166 VSUBS 0.009701f
C204 B.n167 VSUBS 0.009701f
C205 B.n168 VSUBS 0.009701f
C206 B.n169 VSUBS 0.009701f
C207 B.n170 VSUBS 0.009701f
C208 B.n171 VSUBS 0.009701f
C209 B.n172 VSUBS 0.009701f
C210 B.n173 VSUBS 0.009701f
C211 B.n174 VSUBS 0.009701f
C212 B.n175 VSUBS 0.009701f
C213 B.n176 VSUBS 0.009701f
C214 B.n177 VSUBS 0.009701f
C215 B.n178 VSUBS 0.009701f
C216 B.n179 VSUBS 0.009701f
C217 B.n180 VSUBS 0.009701f
C218 B.n181 VSUBS 0.009701f
C219 B.n182 VSUBS 0.009701f
C220 B.n183 VSUBS 0.009701f
C221 B.n184 VSUBS 0.009701f
C222 B.n185 VSUBS 0.009701f
C223 B.n186 VSUBS 0.009701f
C224 B.n187 VSUBS 0.009701f
C225 B.n188 VSUBS 0.009701f
C226 B.n189 VSUBS 0.009701f
C227 B.n190 VSUBS 0.009701f
C228 B.n191 VSUBS 0.009701f
C229 B.n192 VSUBS 0.009701f
C230 B.n193 VSUBS 0.009701f
C231 B.n194 VSUBS 0.009701f
C232 B.n195 VSUBS 0.009701f
C233 B.n196 VSUBS 0.009701f
C234 B.n197 VSUBS 0.009701f
C235 B.n198 VSUBS 0.009701f
C236 B.n199 VSUBS 0.009701f
C237 B.n200 VSUBS 0.009701f
C238 B.n201 VSUBS 0.009701f
C239 B.n202 VSUBS 0.009701f
C240 B.n203 VSUBS 0.009701f
C241 B.n204 VSUBS 0.009701f
C242 B.n205 VSUBS 0.009701f
C243 B.n206 VSUBS 0.009701f
C244 B.n207 VSUBS 0.009701f
C245 B.n208 VSUBS 0.009701f
C246 B.n209 VSUBS 0.009701f
C247 B.n210 VSUBS 0.009701f
C248 B.n211 VSUBS 0.009701f
C249 B.n212 VSUBS 0.009701f
C250 B.n213 VSUBS 0.009701f
C251 B.n214 VSUBS 0.009701f
C252 B.n215 VSUBS 0.009701f
C253 B.n216 VSUBS 0.009701f
C254 B.n217 VSUBS 0.009701f
C255 B.n218 VSUBS 0.009701f
C256 B.n219 VSUBS 0.009701f
C257 B.n220 VSUBS 0.009701f
C258 B.n221 VSUBS 0.009701f
C259 B.n222 VSUBS 0.009701f
C260 B.n223 VSUBS 0.009701f
C261 B.n224 VSUBS 0.009701f
C262 B.n225 VSUBS 0.009701f
C263 B.n226 VSUBS 0.009701f
C264 B.n227 VSUBS 0.009701f
C265 B.n228 VSUBS 0.009701f
C266 B.n229 VSUBS 0.009701f
C267 B.n230 VSUBS 0.009701f
C268 B.n231 VSUBS 0.009701f
C269 B.n232 VSUBS 0.009701f
C270 B.n233 VSUBS 0.009701f
C271 B.n234 VSUBS 0.009701f
C272 B.n235 VSUBS 0.009701f
C273 B.n236 VSUBS 0.009701f
C274 B.n237 VSUBS 0.009701f
C275 B.n238 VSUBS 0.009701f
C276 B.n239 VSUBS 0.009701f
C277 B.n240 VSUBS 0.009701f
C278 B.n241 VSUBS 0.009701f
C279 B.n242 VSUBS 0.009701f
C280 B.n243 VSUBS 0.009701f
C281 B.n244 VSUBS 0.009701f
C282 B.n245 VSUBS 0.021463f
C283 B.n246 VSUBS 0.021463f
C284 B.n247 VSUBS 0.023048f
C285 B.n248 VSUBS 0.009701f
C286 B.n249 VSUBS 0.009701f
C287 B.n250 VSUBS 0.009701f
C288 B.n251 VSUBS 0.009701f
C289 B.n252 VSUBS 0.009701f
C290 B.n253 VSUBS 0.009701f
C291 B.n254 VSUBS 0.009701f
C292 B.n255 VSUBS 0.009701f
C293 B.n256 VSUBS 0.009701f
C294 B.n257 VSUBS 0.009701f
C295 B.n258 VSUBS 0.009701f
C296 B.n259 VSUBS 0.009701f
C297 B.n260 VSUBS 0.009701f
C298 B.n261 VSUBS 0.009701f
C299 B.n262 VSUBS 0.009701f
C300 B.n263 VSUBS 0.009701f
C301 B.n264 VSUBS 0.009701f
C302 B.n265 VSUBS 0.009701f
C303 B.n266 VSUBS 0.009701f
C304 B.n267 VSUBS 0.009701f
C305 B.n268 VSUBS 0.009701f
C306 B.n269 VSUBS 0.009701f
C307 B.n270 VSUBS 0.009701f
C308 B.n271 VSUBS 0.009701f
C309 B.n272 VSUBS 0.009701f
C310 B.n273 VSUBS 0.009701f
C311 B.n274 VSUBS 0.009701f
C312 B.t2 VSUBS 0.093959f
C313 B.t1 VSUBS 0.134898f
C314 B.t0 VSUBS 1.13399f
C315 B.n275 VSUBS 0.226718f
C316 B.n276 VSUBS 0.186079f
C317 B.n277 VSUBS 0.022476f
C318 B.n278 VSUBS 0.00913f
C319 B.n279 VSUBS 0.009701f
C320 B.n280 VSUBS 0.009701f
C321 B.n281 VSUBS 0.009701f
C322 B.n282 VSUBS 0.009701f
C323 B.n283 VSUBS 0.009701f
C324 B.n284 VSUBS 0.009701f
C325 B.n285 VSUBS 0.009701f
C326 B.n286 VSUBS 0.009701f
C327 B.n287 VSUBS 0.009701f
C328 B.n288 VSUBS 0.009701f
C329 B.n289 VSUBS 0.009701f
C330 B.n290 VSUBS 0.009701f
C331 B.n291 VSUBS 0.009701f
C332 B.n292 VSUBS 0.009701f
C333 B.n293 VSUBS 0.009701f
C334 B.n294 VSUBS 0.005421f
C335 B.n295 VSUBS 0.022476f
C336 B.n296 VSUBS 0.00913f
C337 B.n297 VSUBS 0.009701f
C338 B.n298 VSUBS 0.009701f
C339 B.n299 VSUBS 0.009701f
C340 B.n300 VSUBS 0.009701f
C341 B.n301 VSUBS 0.009701f
C342 B.n302 VSUBS 0.009701f
C343 B.n303 VSUBS 0.009701f
C344 B.n304 VSUBS 0.009701f
C345 B.n305 VSUBS 0.009701f
C346 B.n306 VSUBS 0.009701f
C347 B.n307 VSUBS 0.009701f
C348 B.n308 VSUBS 0.009701f
C349 B.n309 VSUBS 0.009701f
C350 B.n310 VSUBS 0.009701f
C351 B.n311 VSUBS 0.009701f
C352 B.n312 VSUBS 0.009701f
C353 B.n313 VSUBS 0.009701f
C354 B.n314 VSUBS 0.009701f
C355 B.n315 VSUBS 0.009701f
C356 B.n316 VSUBS 0.009701f
C357 B.n317 VSUBS 0.009701f
C358 B.n318 VSUBS 0.009701f
C359 B.n319 VSUBS 0.009701f
C360 B.n320 VSUBS 0.009701f
C361 B.n321 VSUBS 0.009701f
C362 B.n322 VSUBS 0.009701f
C363 B.n323 VSUBS 0.009701f
C364 B.n324 VSUBS 0.023048f
C365 B.n325 VSUBS 0.021866f
C366 B.n326 VSUBS 0.022644f
C367 B.n327 VSUBS 0.009701f
C368 B.n328 VSUBS 0.009701f
C369 B.n329 VSUBS 0.009701f
C370 B.n330 VSUBS 0.009701f
C371 B.n331 VSUBS 0.009701f
C372 B.n332 VSUBS 0.009701f
C373 B.n333 VSUBS 0.009701f
C374 B.n334 VSUBS 0.009701f
C375 B.n335 VSUBS 0.009701f
C376 B.n336 VSUBS 0.009701f
C377 B.n337 VSUBS 0.009701f
C378 B.n338 VSUBS 0.009701f
C379 B.n339 VSUBS 0.009701f
C380 B.n340 VSUBS 0.009701f
C381 B.n341 VSUBS 0.009701f
C382 B.n342 VSUBS 0.009701f
C383 B.n343 VSUBS 0.009701f
C384 B.n344 VSUBS 0.009701f
C385 B.n345 VSUBS 0.009701f
C386 B.n346 VSUBS 0.009701f
C387 B.n347 VSUBS 0.009701f
C388 B.n348 VSUBS 0.009701f
C389 B.n349 VSUBS 0.009701f
C390 B.n350 VSUBS 0.009701f
C391 B.n351 VSUBS 0.009701f
C392 B.n352 VSUBS 0.009701f
C393 B.n353 VSUBS 0.009701f
C394 B.n354 VSUBS 0.009701f
C395 B.n355 VSUBS 0.009701f
C396 B.n356 VSUBS 0.009701f
C397 B.n357 VSUBS 0.009701f
C398 B.n358 VSUBS 0.009701f
C399 B.n359 VSUBS 0.009701f
C400 B.n360 VSUBS 0.009701f
C401 B.n361 VSUBS 0.009701f
C402 B.n362 VSUBS 0.009701f
C403 B.n363 VSUBS 0.009701f
C404 B.n364 VSUBS 0.009701f
C405 B.n365 VSUBS 0.009701f
C406 B.n366 VSUBS 0.009701f
C407 B.n367 VSUBS 0.009701f
C408 B.n368 VSUBS 0.009701f
C409 B.n369 VSUBS 0.009701f
C410 B.n370 VSUBS 0.009701f
C411 B.n371 VSUBS 0.009701f
C412 B.n372 VSUBS 0.009701f
C413 B.n373 VSUBS 0.009701f
C414 B.n374 VSUBS 0.009701f
C415 B.n375 VSUBS 0.009701f
C416 B.n376 VSUBS 0.009701f
C417 B.n377 VSUBS 0.009701f
C418 B.n378 VSUBS 0.009701f
C419 B.n379 VSUBS 0.009701f
C420 B.n380 VSUBS 0.009701f
C421 B.n381 VSUBS 0.009701f
C422 B.n382 VSUBS 0.009701f
C423 B.n383 VSUBS 0.009701f
C424 B.n384 VSUBS 0.009701f
C425 B.n385 VSUBS 0.009701f
C426 B.n386 VSUBS 0.009701f
C427 B.n387 VSUBS 0.009701f
C428 B.n388 VSUBS 0.009701f
C429 B.n389 VSUBS 0.009701f
C430 B.n390 VSUBS 0.009701f
C431 B.n391 VSUBS 0.009701f
C432 B.n392 VSUBS 0.009701f
C433 B.n393 VSUBS 0.009701f
C434 B.n394 VSUBS 0.009701f
C435 B.n395 VSUBS 0.009701f
C436 B.n396 VSUBS 0.009701f
C437 B.n397 VSUBS 0.009701f
C438 B.n398 VSUBS 0.009701f
C439 B.n399 VSUBS 0.009701f
C440 B.n400 VSUBS 0.009701f
C441 B.n401 VSUBS 0.009701f
C442 B.n402 VSUBS 0.009701f
C443 B.n403 VSUBS 0.009701f
C444 B.n404 VSUBS 0.009701f
C445 B.n405 VSUBS 0.009701f
C446 B.n406 VSUBS 0.009701f
C447 B.n407 VSUBS 0.009701f
C448 B.n408 VSUBS 0.009701f
C449 B.n409 VSUBS 0.009701f
C450 B.n410 VSUBS 0.009701f
C451 B.n411 VSUBS 0.009701f
C452 B.n412 VSUBS 0.009701f
C453 B.n413 VSUBS 0.009701f
C454 B.n414 VSUBS 0.009701f
C455 B.n415 VSUBS 0.009701f
C456 B.n416 VSUBS 0.009701f
C457 B.n417 VSUBS 0.009701f
C458 B.n418 VSUBS 0.009701f
C459 B.n419 VSUBS 0.009701f
C460 B.n420 VSUBS 0.009701f
C461 B.n421 VSUBS 0.009701f
C462 B.n422 VSUBS 0.009701f
C463 B.n423 VSUBS 0.009701f
C464 B.n424 VSUBS 0.009701f
C465 B.n425 VSUBS 0.009701f
C466 B.n426 VSUBS 0.009701f
C467 B.n427 VSUBS 0.009701f
C468 B.n428 VSUBS 0.009701f
C469 B.n429 VSUBS 0.009701f
C470 B.n430 VSUBS 0.009701f
C471 B.n431 VSUBS 0.009701f
C472 B.n432 VSUBS 0.009701f
C473 B.n433 VSUBS 0.009701f
C474 B.n434 VSUBS 0.009701f
C475 B.n435 VSUBS 0.009701f
C476 B.n436 VSUBS 0.009701f
C477 B.n437 VSUBS 0.009701f
C478 B.n438 VSUBS 0.009701f
C479 B.n439 VSUBS 0.009701f
C480 B.n440 VSUBS 0.009701f
C481 B.n441 VSUBS 0.009701f
C482 B.n442 VSUBS 0.009701f
C483 B.n443 VSUBS 0.009701f
C484 B.n444 VSUBS 0.009701f
C485 B.n445 VSUBS 0.009701f
C486 B.n446 VSUBS 0.009701f
C487 B.n447 VSUBS 0.009701f
C488 B.n448 VSUBS 0.009701f
C489 B.n449 VSUBS 0.009701f
C490 B.n450 VSUBS 0.009701f
C491 B.n451 VSUBS 0.009701f
C492 B.n452 VSUBS 0.009701f
C493 B.n453 VSUBS 0.009701f
C494 B.n454 VSUBS 0.009701f
C495 B.n455 VSUBS 0.009701f
C496 B.n456 VSUBS 0.009701f
C497 B.n457 VSUBS 0.009701f
C498 B.n458 VSUBS 0.009701f
C499 B.n459 VSUBS 0.009701f
C500 B.n460 VSUBS 0.009701f
C501 B.n461 VSUBS 0.009701f
C502 B.n462 VSUBS 0.009701f
C503 B.n463 VSUBS 0.009701f
C504 B.n464 VSUBS 0.009701f
C505 B.n465 VSUBS 0.009701f
C506 B.n466 VSUBS 0.009701f
C507 B.n467 VSUBS 0.009701f
C508 B.n468 VSUBS 0.009701f
C509 B.n469 VSUBS 0.009701f
C510 B.n470 VSUBS 0.009701f
C511 B.n471 VSUBS 0.009701f
C512 B.n472 VSUBS 0.009701f
C513 B.n473 VSUBS 0.009701f
C514 B.n474 VSUBS 0.009701f
C515 B.n475 VSUBS 0.009701f
C516 B.n476 VSUBS 0.009701f
C517 B.n477 VSUBS 0.009701f
C518 B.n478 VSUBS 0.009701f
C519 B.n479 VSUBS 0.009701f
C520 B.n480 VSUBS 0.009701f
C521 B.n481 VSUBS 0.009701f
C522 B.n482 VSUBS 0.009701f
C523 B.n483 VSUBS 0.009701f
C524 B.n484 VSUBS 0.009701f
C525 B.n485 VSUBS 0.009701f
C526 B.n486 VSUBS 0.009701f
C527 B.n487 VSUBS 0.009701f
C528 B.n488 VSUBS 0.009701f
C529 B.n489 VSUBS 0.021463f
C530 B.n490 VSUBS 0.021463f
C531 B.n491 VSUBS 0.023048f
C532 B.n492 VSUBS 0.009701f
C533 B.n493 VSUBS 0.009701f
C534 B.n494 VSUBS 0.009701f
C535 B.n495 VSUBS 0.009701f
C536 B.n496 VSUBS 0.009701f
C537 B.n497 VSUBS 0.009701f
C538 B.n498 VSUBS 0.009701f
C539 B.n499 VSUBS 0.009701f
C540 B.n500 VSUBS 0.009701f
C541 B.n501 VSUBS 0.009701f
C542 B.n502 VSUBS 0.009701f
C543 B.n503 VSUBS 0.009701f
C544 B.n504 VSUBS 0.009701f
C545 B.n505 VSUBS 0.009701f
C546 B.n506 VSUBS 0.009701f
C547 B.n507 VSUBS 0.009701f
C548 B.n508 VSUBS 0.009701f
C549 B.n509 VSUBS 0.009701f
C550 B.n510 VSUBS 0.009701f
C551 B.n511 VSUBS 0.009701f
C552 B.n512 VSUBS 0.009701f
C553 B.n513 VSUBS 0.009701f
C554 B.n514 VSUBS 0.009701f
C555 B.n515 VSUBS 0.009701f
C556 B.n516 VSUBS 0.009701f
C557 B.n517 VSUBS 0.009701f
C558 B.n518 VSUBS 0.009701f
C559 B.n519 VSUBS 0.00913f
C560 B.n520 VSUBS 0.009701f
C561 B.n521 VSUBS 0.009701f
C562 B.n522 VSUBS 0.005421f
C563 B.n523 VSUBS 0.009701f
C564 B.n524 VSUBS 0.009701f
C565 B.n525 VSUBS 0.009701f
C566 B.n526 VSUBS 0.009701f
C567 B.n527 VSUBS 0.009701f
C568 B.n528 VSUBS 0.009701f
C569 B.n529 VSUBS 0.009701f
C570 B.n530 VSUBS 0.009701f
C571 B.n531 VSUBS 0.009701f
C572 B.n532 VSUBS 0.009701f
C573 B.n533 VSUBS 0.009701f
C574 B.n534 VSUBS 0.009701f
C575 B.n535 VSUBS 0.005421f
C576 B.n536 VSUBS 0.022476f
C577 B.n537 VSUBS 0.00913f
C578 B.n538 VSUBS 0.009701f
C579 B.n539 VSUBS 0.009701f
C580 B.n540 VSUBS 0.009701f
C581 B.n541 VSUBS 0.009701f
C582 B.n542 VSUBS 0.009701f
C583 B.n543 VSUBS 0.009701f
C584 B.n544 VSUBS 0.009701f
C585 B.n545 VSUBS 0.009701f
C586 B.n546 VSUBS 0.009701f
C587 B.n547 VSUBS 0.009701f
C588 B.n548 VSUBS 0.009701f
C589 B.n549 VSUBS 0.009701f
C590 B.n550 VSUBS 0.009701f
C591 B.n551 VSUBS 0.009701f
C592 B.n552 VSUBS 0.009701f
C593 B.n553 VSUBS 0.009701f
C594 B.n554 VSUBS 0.009701f
C595 B.n555 VSUBS 0.009701f
C596 B.n556 VSUBS 0.009701f
C597 B.n557 VSUBS 0.009701f
C598 B.n558 VSUBS 0.009701f
C599 B.n559 VSUBS 0.009701f
C600 B.n560 VSUBS 0.009701f
C601 B.n561 VSUBS 0.009701f
C602 B.n562 VSUBS 0.009701f
C603 B.n563 VSUBS 0.009701f
C604 B.n564 VSUBS 0.009701f
C605 B.n565 VSUBS 0.009701f
C606 B.n566 VSUBS 0.023048f
C607 B.n567 VSUBS 0.021463f
C608 B.n568 VSUBS 0.021463f
C609 B.n569 VSUBS 0.009701f
C610 B.n570 VSUBS 0.009701f
C611 B.n571 VSUBS 0.009701f
C612 B.n572 VSUBS 0.009701f
C613 B.n573 VSUBS 0.009701f
C614 B.n574 VSUBS 0.009701f
C615 B.n575 VSUBS 0.009701f
C616 B.n576 VSUBS 0.009701f
C617 B.n577 VSUBS 0.009701f
C618 B.n578 VSUBS 0.009701f
C619 B.n579 VSUBS 0.009701f
C620 B.n580 VSUBS 0.009701f
C621 B.n581 VSUBS 0.009701f
C622 B.n582 VSUBS 0.009701f
C623 B.n583 VSUBS 0.009701f
C624 B.n584 VSUBS 0.009701f
C625 B.n585 VSUBS 0.009701f
C626 B.n586 VSUBS 0.009701f
C627 B.n587 VSUBS 0.009701f
C628 B.n588 VSUBS 0.009701f
C629 B.n589 VSUBS 0.009701f
C630 B.n590 VSUBS 0.009701f
C631 B.n591 VSUBS 0.009701f
C632 B.n592 VSUBS 0.009701f
C633 B.n593 VSUBS 0.009701f
C634 B.n594 VSUBS 0.009701f
C635 B.n595 VSUBS 0.009701f
C636 B.n596 VSUBS 0.009701f
C637 B.n597 VSUBS 0.009701f
C638 B.n598 VSUBS 0.009701f
C639 B.n599 VSUBS 0.009701f
C640 B.n600 VSUBS 0.009701f
C641 B.n601 VSUBS 0.009701f
C642 B.n602 VSUBS 0.009701f
C643 B.n603 VSUBS 0.009701f
C644 B.n604 VSUBS 0.009701f
C645 B.n605 VSUBS 0.009701f
C646 B.n606 VSUBS 0.009701f
C647 B.n607 VSUBS 0.009701f
C648 B.n608 VSUBS 0.009701f
C649 B.n609 VSUBS 0.009701f
C650 B.n610 VSUBS 0.009701f
C651 B.n611 VSUBS 0.009701f
C652 B.n612 VSUBS 0.009701f
C653 B.n613 VSUBS 0.009701f
C654 B.n614 VSUBS 0.009701f
C655 B.n615 VSUBS 0.009701f
C656 B.n616 VSUBS 0.009701f
C657 B.n617 VSUBS 0.009701f
C658 B.n618 VSUBS 0.009701f
C659 B.n619 VSUBS 0.009701f
C660 B.n620 VSUBS 0.009701f
C661 B.n621 VSUBS 0.009701f
C662 B.n622 VSUBS 0.009701f
C663 B.n623 VSUBS 0.009701f
C664 B.n624 VSUBS 0.009701f
C665 B.n625 VSUBS 0.009701f
C666 B.n626 VSUBS 0.009701f
C667 B.n627 VSUBS 0.009701f
C668 B.n628 VSUBS 0.009701f
C669 B.n629 VSUBS 0.009701f
C670 B.n630 VSUBS 0.009701f
C671 B.n631 VSUBS 0.009701f
C672 B.n632 VSUBS 0.009701f
C673 B.n633 VSUBS 0.009701f
C674 B.n634 VSUBS 0.009701f
C675 B.n635 VSUBS 0.009701f
C676 B.n636 VSUBS 0.009701f
C677 B.n637 VSUBS 0.009701f
C678 B.n638 VSUBS 0.009701f
C679 B.n639 VSUBS 0.009701f
C680 B.n640 VSUBS 0.009701f
C681 B.n641 VSUBS 0.009701f
C682 B.n642 VSUBS 0.009701f
C683 B.n643 VSUBS 0.009701f
C684 B.n644 VSUBS 0.009701f
C685 B.n645 VSUBS 0.009701f
C686 B.n646 VSUBS 0.009701f
C687 B.n647 VSUBS 0.012659f
C688 B.n648 VSUBS 0.013485f
C689 B.n649 VSUBS 0.026817f
C690 VDD1.n0 VSUBS 0.030637f
C691 VDD1.n1 VSUBS 0.027667f
C692 VDD1.n2 VSUBS 0.014867f
C693 VDD1.n3 VSUBS 0.03514f
C694 VDD1.n4 VSUBS 0.015742f
C695 VDD1.n5 VSUBS 0.465025f
C696 VDD1.n6 VSUBS 0.014867f
C697 VDD1.t3 VSUBS 0.076786f
C698 VDD1.n7 VSUBS 0.112674f
C699 VDD1.n8 VSUBS 0.022262f
C700 VDD1.n9 VSUBS 0.026355f
C701 VDD1.n10 VSUBS 0.03514f
C702 VDD1.n11 VSUBS 0.015742f
C703 VDD1.n12 VSUBS 0.014867f
C704 VDD1.n13 VSUBS 0.027667f
C705 VDD1.n14 VSUBS 0.027667f
C706 VDD1.n15 VSUBS 0.014867f
C707 VDD1.n16 VSUBS 0.015742f
C708 VDD1.n17 VSUBS 0.03514f
C709 VDD1.n18 VSUBS 0.085876f
C710 VDD1.n19 VSUBS 0.015742f
C711 VDD1.n20 VSUBS 0.014867f
C712 VDD1.n21 VSUBS 0.068109f
C713 VDD1.n22 VSUBS 0.076477f
C714 VDD1.n23 VSUBS 0.030637f
C715 VDD1.n24 VSUBS 0.027667f
C716 VDD1.n25 VSUBS 0.014867f
C717 VDD1.n26 VSUBS 0.03514f
C718 VDD1.n27 VSUBS 0.015742f
C719 VDD1.n28 VSUBS 0.465025f
C720 VDD1.n29 VSUBS 0.014867f
C721 VDD1.t2 VSUBS 0.076786f
C722 VDD1.n30 VSUBS 0.112674f
C723 VDD1.n31 VSUBS 0.022262f
C724 VDD1.n32 VSUBS 0.026355f
C725 VDD1.n33 VSUBS 0.03514f
C726 VDD1.n34 VSUBS 0.015742f
C727 VDD1.n35 VSUBS 0.014867f
C728 VDD1.n36 VSUBS 0.027667f
C729 VDD1.n37 VSUBS 0.027667f
C730 VDD1.n38 VSUBS 0.014867f
C731 VDD1.n39 VSUBS 0.015742f
C732 VDD1.n40 VSUBS 0.03514f
C733 VDD1.n41 VSUBS 0.085876f
C734 VDD1.n42 VSUBS 0.015742f
C735 VDD1.n43 VSUBS 0.014867f
C736 VDD1.n44 VSUBS 0.068109f
C737 VDD1.n45 VSUBS 0.075434f
C738 VDD1.t4 VSUBS 0.102102f
C739 VDD1.t1 VSUBS 0.102102f
C740 VDD1.n46 VSUBS 0.634882f
C741 VDD1.n47 VSUBS 3.3046f
C742 VDD1.t5 VSUBS 0.102102f
C743 VDD1.t0 VSUBS 0.102102f
C744 VDD1.n48 VSUBS 0.628935f
C745 VDD1.n49 VSUBS 2.96633f
C746 VP.t4 VSUBS 1.86386f
C747 VP.n0 VSUBS 0.876124f
C748 VP.n1 VSUBS 0.042365f
C749 VP.n2 VSUBS 0.064801f
C750 VP.n3 VSUBS 0.042365f
C751 VP.n4 VSUBS 0.059467f
C752 VP.n5 VSUBS 0.042365f
C753 VP.n6 VSUBS 0.058898f
C754 VP.n7 VSUBS 0.042365f
C755 VP.n8 VSUBS 0.055569f
C756 VP.t5 VSUBS 1.86386f
C757 VP.n9 VSUBS 0.876124f
C758 VP.n10 VSUBS 0.042365f
C759 VP.n11 VSUBS 0.064801f
C760 VP.n12 VSUBS 0.042365f
C761 VP.n13 VSUBS 0.059467f
C762 VP.t2 VSUBS 2.39794f
C763 VP.t0 VSUBS 1.86386f
C764 VP.n14 VSUBS 0.855566f
C765 VP.n15 VSUBS 0.835013f
C766 VP.n16 VSUBS 0.52974f
C767 VP.n17 VSUBS 0.042365f
C768 VP.n18 VSUBS 0.078958f
C769 VP.n19 VSUBS 0.078958f
C770 VP.n20 VSUBS 0.058898f
C771 VP.n21 VSUBS 0.042365f
C772 VP.n22 VSUBS 0.042365f
C773 VP.n23 VSUBS 0.042365f
C774 VP.n24 VSUBS 0.078958f
C775 VP.n25 VSUBS 0.078958f
C776 VP.n26 VSUBS 0.055569f
C777 VP.n27 VSUBS 0.068376f
C778 VP.n28 VSUBS 2.23465f
C779 VP.t3 VSUBS 1.86386f
C780 VP.n29 VSUBS 0.876124f
C781 VP.n30 VSUBS 2.26688f
C782 VP.n31 VSUBS 0.068376f
C783 VP.n32 VSUBS 0.042365f
C784 VP.n33 VSUBS 0.078958f
C785 VP.n34 VSUBS 0.078958f
C786 VP.n35 VSUBS 0.064801f
C787 VP.n36 VSUBS 0.042365f
C788 VP.n37 VSUBS 0.042365f
C789 VP.n38 VSUBS 0.042365f
C790 VP.n39 VSUBS 0.078958f
C791 VP.n40 VSUBS 0.078958f
C792 VP.t1 VSUBS 1.86386f
C793 VP.n41 VSUBS 0.708023f
C794 VP.n42 VSUBS 0.059467f
C795 VP.n43 VSUBS 0.042365f
C796 VP.n44 VSUBS 0.042365f
C797 VP.n45 VSUBS 0.042365f
C798 VP.n46 VSUBS 0.078958f
C799 VP.n47 VSUBS 0.078958f
C800 VP.n48 VSUBS 0.058898f
C801 VP.n49 VSUBS 0.042365f
C802 VP.n50 VSUBS 0.042365f
C803 VP.n51 VSUBS 0.042365f
C804 VP.n52 VSUBS 0.078958f
C805 VP.n53 VSUBS 0.078958f
C806 VP.n54 VSUBS 0.055569f
C807 VP.n55 VSUBS 0.068376f
C808 VP.n56 VSUBS 0.116528f
C809 VTAIL.t4 VSUBS 0.136108f
C810 VTAIL.t9 VSUBS 0.136108f
C811 VTAIL.n0 VSUBS 0.737156f
C812 VTAIL.n1 VSUBS 0.967905f
C813 VTAIL.n2 VSUBS 0.04084f
C814 VTAIL.n3 VSUBS 0.036882f
C815 VTAIL.n4 VSUBS 0.019819f
C816 VTAIL.n5 VSUBS 0.046844f
C817 VTAIL.n6 VSUBS 0.020985f
C818 VTAIL.n7 VSUBS 0.619903f
C819 VTAIL.n8 VSUBS 0.019819f
C820 VTAIL.t11 VSUBS 0.10236f
C821 VTAIL.n9 VSUBS 0.1502f
C822 VTAIL.n10 VSUBS 0.029676f
C823 VTAIL.n11 VSUBS 0.035133f
C824 VTAIL.n12 VSUBS 0.046844f
C825 VTAIL.n13 VSUBS 0.020985f
C826 VTAIL.n14 VSUBS 0.019819f
C827 VTAIL.n15 VSUBS 0.036882f
C828 VTAIL.n16 VSUBS 0.036882f
C829 VTAIL.n17 VSUBS 0.019819f
C830 VTAIL.n18 VSUBS 0.020985f
C831 VTAIL.n19 VSUBS 0.046844f
C832 VTAIL.n20 VSUBS 0.114477f
C833 VTAIL.n21 VSUBS 0.020985f
C834 VTAIL.n22 VSUBS 0.019819f
C835 VTAIL.n23 VSUBS 0.090793f
C836 VTAIL.n24 VSUBS 0.057783f
C837 VTAIL.n25 VSUBS 0.697481f
C838 VTAIL.t0 VSUBS 0.136108f
C839 VTAIL.t2 VSUBS 0.136108f
C840 VTAIL.n26 VSUBS 0.737156f
C841 VTAIL.n27 VSUBS 2.79511f
C842 VTAIL.t8 VSUBS 0.136108f
C843 VTAIL.t7 VSUBS 0.136108f
C844 VTAIL.n28 VSUBS 0.737161f
C845 VTAIL.n29 VSUBS 2.79511f
C846 VTAIL.n30 VSUBS 0.04084f
C847 VTAIL.n31 VSUBS 0.036882f
C848 VTAIL.n32 VSUBS 0.019819f
C849 VTAIL.n33 VSUBS 0.046844f
C850 VTAIL.n34 VSUBS 0.020985f
C851 VTAIL.n35 VSUBS 0.619903f
C852 VTAIL.n36 VSUBS 0.019819f
C853 VTAIL.t6 VSUBS 0.10236f
C854 VTAIL.n37 VSUBS 0.1502f
C855 VTAIL.n38 VSUBS 0.029676f
C856 VTAIL.n39 VSUBS 0.035133f
C857 VTAIL.n40 VSUBS 0.046844f
C858 VTAIL.n41 VSUBS 0.020985f
C859 VTAIL.n42 VSUBS 0.019819f
C860 VTAIL.n43 VSUBS 0.036882f
C861 VTAIL.n44 VSUBS 0.036882f
C862 VTAIL.n45 VSUBS 0.019819f
C863 VTAIL.n46 VSUBS 0.020985f
C864 VTAIL.n47 VSUBS 0.046844f
C865 VTAIL.n48 VSUBS 0.114477f
C866 VTAIL.n49 VSUBS 0.020985f
C867 VTAIL.n50 VSUBS 0.019819f
C868 VTAIL.n51 VSUBS 0.090793f
C869 VTAIL.n52 VSUBS 0.057783f
C870 VTAIL.n53 VSUBS 0.697481f
C871 VTAIL.t10 VSUBS 0.136108f
C872 VTAIL.t3 VSUBS 0.136108f
C873 VTAIL.n54 VSUBS 0.737161f
C874 VTAIL.n55 VSUBS 1.26449f
C875 VTAIL.n56 VSUBS 0.04084f
C876 VTAIL.n57 VSUBS 0.036882f
C877 VTAIL.n58 VSUBS 0.019819f
C878 VTAIL.n59 VSUBS 0.046844f
C879 VTAIL.n60 VSUBS 0.020985f
C880 VTAIL.n61 VSUBS 0.619903f
C881 VTAIL.n62 VSUBS 0.019819f
C882 VTAIL.t1 VSUBS 0.10236f
C883 VTAIL.n63 VSUBS 0.1502f
C884 VTAIL.n64 VSUBS 0.029676f
C885 VTAIL.n65 VSUBS 0.035133f
C886 VTAIL.n66 VSUBS 0.046844f
C887 VTAIL.n67 VSUBS 0.020985f
C888 VTAIL.n68 VSUBS 0.019819f
C889 VTAIL.n69 VSUBS 0.036882f
C890 VTAIL.n70 VSUBS 0.036882f
C891 VTAIL.n71 VSUBS 0.019819f
C892 VTAIL.n72 VSUBS 0.020985f
C893 VTAIL.n73 VSUBS 0.046844f
C894 VTAIL.n74 VSUBS 0.114477f
C895 VTAIL.n75 VSUBS 0.020985f
C896 VTAIL.n76 VSUBS 0.019819f
C897 VTAIL.n77 VSUBS 0.090793f
C898 VTAIL.n78 VSUBS 0.057783f
C899 VTAIL.n79 VSUBS 1.82342f
C900 VTAIL.n80 VSUBS 0.04084f
C901 VTAIL.n81 VSUBS 0.036882f
C902 VTAIL.n82 VSUBS 0.019819f
C903 VTAIL.n83 VSUBS 0.046844f
C904 VTAIL.n84 VSUBS 0.020985f
C905 VTAIL.n85 VSUBS 0.619903f
C906 VTAIL.n86 VSUBS 0.019819f
C907 VTAIL.t5 VSUBS 0.10236f
C908 VTAIL.n87 VSUBS 0.1502f
C909 VTAIL.n88 VSUBS 0.029676f
C910 VTAIL.n89 VSUBS 0.035133f
C911 VTAIL.n90 VSUBS 0.046844f
C912 VTAIL.n91 VSUBS 0.020985f
C913 VTAIL.n92 VSUBS 0.019819f
C914 VTAIL.n93 VSUBS 0.036882f
C915 VTAIL.n94 VSUBS 0.036882f
C916 VTAIL.n95 VSUBS 0.019819f
C917 VTAIL.n96 VSUBS 0.020985f
C918 VTAIL.n97 VSUBS 0.046844f
C919 VTAIL.n98 VSUBS 0.114477f
C920 VTAIL.n99 VSUBS 0.020985f
C921 VTAIL.n100 VSUBS 0.019819f
C922 VTAIL.n101 VSUBS 0.090793f
C923 VTAIL.n102 VSUBS 0.057783f
C924 VTAIL.n103 VSUBS 1.71534f
C925 VDD2.n0 VSUBS 0.030643f
C926 VDD2.n1 VSUBS 0.027673f
C927 VDD2.n2 VSUBS 0.01487f
C928 VDD2.n3 VSUBS 0.035147f
C929 VDD2.n4 VSUBS 0.015745f
C930 VDD2.n5 VSUBS 0.465118f
C931 VDD2.n6 VSUBS 0.01487f
C932 VDD2.t1 VSUBS 0.076801f
C933 VDD2.n7 VSUBS 0.112696f
C934 VDD2.n8 VSUBS 0.022266f
C935 VDD2.n9 VSUBS 0.026361f
C936 VDD2.n10 VSUBS 0.035147f
C937 VDD2.n11 VSUBS 0.015745f
C938 VDD2.n12 VSUBS 0.01487f
C939 VDD2.n13 VSUBS 0.027673f
C940 VDD2.n14 VSUBS 0.027673f
C941 VDD2.n15 VSUBS 0.01487f
C942 VDD2.n16 VSUBS 0.015745f
C943 VDD2.n17 VSUBS 0.035147f
C944 VDD2.n18 VSUBS 0.085893f
C945 VDD2.n19 VSUBS 0.015745f
C946 VDD2.n20 VSUBS 0.01487f
C947 VDD2.n21 VSUBS 0.068122f
C948 VDD2.n22 VSUBS 0.075449f
C949 VDD2.t2 VSUBS 0.102123f
C950 VDD2.t0 VSUBS 0.102123f
C951 VDD2.n23 VSUBS 0.635008f
C952 VDD2.n24 VSUBS 3.14699f
C953 VDD2.n25 VSUBS 0.030643f
C954 VDD2.n26 VSUBS 0.027673f
C955 VDD2.n27 VSUBS 0.01487f
C956 VDD2.n28 VSUBS 0.035147f
C957 VDD2.n29 VSUBS 0.015745f
C958 VDD2.n30 VSUBS 0.465118f
C959 VDD2.n31 VSUBS 0.01487f
C960 VDD2.t5 VSUBS 0.076801f
C961 VDD2.n32 VSUBS 0.112696f
C962 VDD2.n33 VSUBS 0.022266f
C963 VDD2.n34 VSUBS 0.026361f
C964 VDD2.n35 VSUBS 0.035147f
C965 VDD2.n36 VSUBS 0.015745f
C966 VDD2.n37 VSUBS 0.01487f
C967 VDD2.n38 VSUBS 0.027673f
C968 VDD2.n39 VSUBS 0.027673f
C969 VDD2.n40 VSUBS 0.01487f
C970 VDD2.n41 VSUBS 0.015745f
C971 VDD2.n42 VSUBS 0.035147f
C972 VDD2.n43 VSUBS 0.085893f
C973 VDD2.n44 VSUBS 0.015745f
C974 VDD2.n45 VSUBS 0.01487f
C975 VDD2.n46 VSUBS 0.068122f
C976 VDD2.n47 VSUBS 0.062431f
C977 VDD2.n48 VSUBS 2.51299f
C978 VDD2.t3 VSUBS 0.102123f
C979 VDD2.t4 VSUBS 0.102123f
C980 VDD2.n49 VSUBS 0.634979f
C981 VN.t4 VSUBS 1.61849f
C982 VN.n0 VSUBS 0.760784f
C983 VN.n1 VSUBS 0.036788f
C984 VN.n2 VSUBS 0.05627f
C985 VN.n3 VSUBS 0.036788f
C986 VN.n4 VSUBS 0.051638f
C987 VN.t0 VSUBS 1.61849f
C988 VN.n5 VSUBS 0.742932f
C989 VN.t5 VSUBS 2.08226f
C990 VN.n6 VSUBS 0.725083f
C991 VN.n7 VSUBS 0.46f
C992 VN.n8 VSUBS 0.036788f
C993 VN.n9 VSUBS 0.068563f
C994 VN.n10 VSUBS 0.068563f
C995 VN.n11 VSUBS 0.051144f
C996 VN.n12 VSUBS 0.036788f
C997 VN.n13 VSUBS 0.036788f
C998 VN.n14 VSUBS 0.036788f
C999 VN.n15 VSUBS 0.068563f
C1000 VN.n16 VSUBS 0.068563f
C1001 VN.n17 VSUBS 0.048253f
C1002 VN.n18 VSUBS 0.059375f
C1003 VN.n19 VSUBS 0.101187f
C1004 VN.t1 VSUBS 1.61849f
C1005 VN.n20 VSUBS 0.760784f
C1006 VN.n21 VSUBS 0.036788f
C1007 VN.n22 VSUBS 0.05627f
C1008 VN.n23 VSUBS 0.036788f
C1009 VN.n24 VSUBS 0.051638f
C1010 VN.t3 VSUBS 2.08226f
C1011 VN.t2 VSUBS 1.61849f
C1012 VN.n25 VSUBS 0.742932f
C1013 VN.n26 VSUBS 0.725083f
C1014 VN.n27 VSUBS 0.46f
C1015 VN.n28 VSUBS 0.036788f
C1016 VN.n29 VSUBS 0.068563f
C1017 VN.n30 VSUBS 0.068563f
C1018 VN.n31 VSUBS 0.051144f
C1019 VN.n32 VSUBS 0.036788f
C1020 VN.n33 VSUBS 0.036788f
C1021 VN.n34 VSUBS 0.036788f
C1022 VN.n35 VSUBS 0.068563f
C1023 VN.n36 VSUBS 0.068563f
C1024 VN.n37 VSUBS 0.048253f
C1025 VN.n38 VSUBS 0.059375f
C1026 VN.n39 VSUBS 1.9558f
.ends

