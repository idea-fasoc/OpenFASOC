* NGSPICE file created from diff_pair_sample_0166.ext - technology: sky130A

.subckt diff_pair_sample_0166 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0.8778 ps=5.65 w=5.32 l=1.85
X1 VDD2.t7 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X2 VTAIL.t14 VP.t1 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X3 VDD1.t4 VP.t2 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X4 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0.8778 ps=5.65 w=5.32 l=1.85
X5 VTAIL.t2 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X6 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0.8778 ps=5.65 w=5.32 l=1.85
X7 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0 ps=0 w=5.32 l=1.85
X8 VDD2.t3 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X9 VDD1.t1 VP.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=2.0748 ps=11.42 w=5.32 l=1.85
X10 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=2.0748 ps=11.42 w=5.32 l=1.85
X11 VDD1.t3 VP.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=2.0748 ps=11.42 w=5.32 l=1.85
X12 VTAIL.t10 VP.t5 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0.8778 ps=5.65 w=5.32 l=1.85
X13 VTAIL.t1 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X14 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=2.0748 ps=11.42 w=5.32 l=1.85
X15 VTAIL.t9 VP.t6 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X16 VDD1.t6 VP.t7 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8778 pd=5.65 as=0.8778 ps=5.65 w=5.32 l=1.85
X17 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0 ps=0 w=5.32 l=1.85
X18 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0 ps=0 w=5.32 l=1.85
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0748 pd=11.42 as=0 ps=0 w=5.32 l=1.85
R0 VP.n31 VP.n7 184.909
R1 VP.n56 VP.n55 184.909
R2 VP.n30 VP.n29 184.909
R3 VP.n15 VP.n12 161.3
R4 VP.n17 VP.n16 161.3
R5 VP.n18 VP.n11 161.3
R6 VP.n20 VP.n19 161.3
R7 VP.n22 VP.n10 161.3
R8 VP.n24 VP.n23 161.3
R9 VP.n25 VP.n9 161.3
R10 VP.n27 VP.n26 161.3
R11 VP.n28 VP.n8 161.3
R12 VP.n54 VP.n0 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n51 VP.n1 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n48 VP.n2 161.3
R17 VP.n46 VP.n45 161.3
R18 VP.n44 VP.n3 161.3
R19 VP.n43 VP.n42 161.3
R20 VP.n41 VP.n4 161.3
R21 VP.n39 VP.n38 161.3
R22 VP.n37 VP.n5 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n34 VP.n6 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n13 VP.t0 101.775
R27 VP.n7 VP.t5 69.3043
R28 VP.n40 VP.t7 69.3043
R29 VP.n47 VP.t6 69.3043
R30 VP.n55 VP.t4 69.3043
R31 VP.n29 VP.t3 69.3043
R32 VP.n21 VP.t1 69.3043
R33 VP.n14 VP.t2 69.3043
R34 VP.n42 VP.n3 56.5617
R35 VP.n16 VP.n11 56.5617
R36 VP.n14 VP.n13 53.2962
R37 VP.n35 VP.n5 47.3584
R38 VP.n49 VP.n1 47.3584
R39 VP.n23 VP.n9 47.3584
R40 VP.n31 VP.n30 42.1975
R41 VP.n35 VP.n34 33.7956
R42 VP.n53 VP.n1 33.7956
R43 VP.n27 VP.n9 33.7956
R44 VP.n34 VP.n33 24.5923
R45 VP.n39 VP.n5 24.5923
R46 VP.n42 VP.n41 24.5923
R47 VP.n46 VP.n3 24.5923
R48 VP.n49 VP.n48 24.5923
R49 VP.n54 VP.n53 24.5923
R50 VP.n28 VP.n27 24.5923
R51 VP.n20 VP.n11 24.5923
R52 VP.n23 VP.n22 24.5923
R53 VP.n16 VP.n15 24.5923
R54 VP.n41 VP.n40 16.7229
R55 VP.n47 VP.n46 16.7229
R56 VP.n21 VP.n20 16.7229
R57 VP.n15 VP.n14 16.7229
R58 VP.n13 VP.n12 12.4908
R59 VP.n40 VP.n39 7.86989
R60 VP.n48 VP.n47 7.86989
R61 VP.n22 VP.n21 7.86989
R62 VP.n33 VP.n7 0.984173
R63 VP.n55 VP.n54 0.984173
R64 VP.n29 VP.n28 0.984173
R65 VP.n17 VP.n12 0.189894
R66 VP.n18 VP.n17 0.189894
R67 VP.n19 VP.n18 0.189894
R68 VP.n19 VP.n10 0.189894
R69 VP.n24 VP.n10 0.189894
R70 VP.n25 VP.n24 0.189894
R71 VP.n26 VP.n25 0.189894
R72 VP.n26 VP.n8 0.189894
R73 VP.n30 VP.n8 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n32 VP.n6 0.189894
R76 VP.n36 VP.n6 0.189894
R77 VP.n37 VP.n36 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n38 VP.n4 0.189894
R80 VP.n43 VP.n4 0.189894
R81 VP.n44 VP.n43 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n45 VP.n2 0.189894
R84 VP.n50 VP.n2 0.189894
R85 VP.n51 VP.n50 0.189894
R86 VP.n52 VP.n51 0.189894
R87 VP.n52 VP.n0 0.189894
R88 VP.n56 VP.n0 0.189894
R89 VP VP.n56 0.0516364
R90 VDD1 VDD1.n0 70.4289
R91 VDD1.n3 VDD1.n2 70.3152
R92 VDD1.n3 VDD1.n1 70.3152
R93 VDD1.n5 VDD1.n4 69.4309
R94 VDD1.n5 VDD1.n3 37.3414
R95 VDD1.n4 VDD1.t5 3.7223
R96 VDD1.n4 VDD1.t1 3.7223
R97 VDD1.n0 VDD1.t2 3.7223
R98 VDD1.n0 VDD1.t4 3.7223
R99 VDD1.n2 VDD1.t0 3.7223
R100 VDD1.n2 VDD1.t3 3.7223
R101 VDD1.n1 VDD1.t7 3.7223
R102 VDD1.n1 VDD1.t6 3.7223
R103 VDD1 VDD1.n5 0.881965
R104 VTAIL.n226 VTAIL.n204 289.615
R105 VTAIL.n24 VTAIL.n2 289.615
R106 VTAIL.n52 VTAIL.n30 289.615
R107 VTAIL.n82 VTAIL.n60 289.615
R108 VTAIL.n198 VTAIL.n176 289.615
R109 VTAIL.n168 VTAIL.n146 289.615
R110 VTAIL.n140 VTAIL.n118 289.615
R111 VTAIL.n110 VTAIL.n88 289.615
R112 VTAIL.n212 VTAIL.n211 185
R113 VTAIL.n217 VTAIL.n216 185
R114 VTAIL.n219 VTAIL.n218 185
R115 VTAIL.n208 VTAIL.n207 185
R116 VTAIL.n225 VTAIL.n224 185
R117 VTAIL.n227 VTAIL.n226 185
R118 VTAIL.n10 VTAIL.n9 185
R119 VTAIL.n15 VTAIL.n14 185
R120 VTAIL.n17 VTAIL.n16 185
R121 VTAIL.n6 VTAIL.n5 185
R122 VTAIL.n23 VTAIL.n22 185
R123 VTAIL.n25 VTAIL.n24 185
R124 VTAIL.n38 VTAIL.n37 185
R125 VTAIL.n43 VTAIL.n42 185
R126 VTAIL.n45 VTAIL.n44 185
R127 VTAIL.n34 VTAIL.n33 185
R128 VTAIL.n51 VTAIL.n50 185
R129 VTAIL.n53 VTAIL.n52 185
R130 VTAIL.n68 VTAIL.n67 185
R131 VTAIL.n73 VTAIL.n72 185
R132 VTAIL.n75 VTAIL.n74 185
R133 VTAIL.n64 VTAIL.n63 185
R134 VTAIL.n81 VTAIL.n80 185
R135 VTAIL.n83 VTAIL.n82 185
R136 VTAIL.n199 VTAIL.n198 185
R137 VTAIL.n197 VTAIL.n196 185
R138 VTAIL.n180 VTAIL.n179 185
R139 VTAIL.n191 VTAIL.n190 185
R140 VTAIL.n189 VTAIL.n188 185
R141 VTAIL.n184 VTAIL.n183 185
R142 VTAIL.n169 VTAIL.n168 185
R143 VTAIL.n167 VTAIL.n166 185
R144 VTAIL.n150 VTAIL.n149 185
R145 VTAIL.n161 VTAIL.n160 185
R146 VTAIL.n159 VTAIL.n158 185
R147 VTAIL.n154 VTAIL.n153 185
R148 VTAIL.n141 VTAIL.n140 185
R149 VTAIL.n139 VTAIL.n138 185
R150 VTAIL.n122 VTAIL.n121 185
R151 VTAIL.n133 VTAIL.n132 185
R152 VTAIL.n131 VTAIL.n130 185
R153 VTAIL.n126 VTAIL.n125 185
R154 VTAIL.n111 VTAIL.n110 185
R155 VTAIL.n109 VTAIL.n108 185
R156 VTAIL.n92 VTAIL.n91 185
R157 VTAIL.n103 VTAIL.n102 185
R158 VTAIL.n101 VTAIL.n100 185
R159 VTAIL.n96 VTAIL.n95 185
R160 VTAIL.n213 VTAIL.t0 147.672
R161 VTAIL.n11 VTAIL.t4 147.672
R162 VTAIL.n39 VTAIL.t11 147.672
R163 VTAIL.n69 VTAIL.t10 147.672
R164 VTAIL.n185 VTAIL.t12 147.672
R165 VTAIL.n155 VTAIL.t15 147.672
R166 VTAIL.n127 VTAIL.t6 147.672
R167 VTAIL.n97 VTAIL.t3 147.672
R168 VTAIL.n217 VTAIL.n211 104.615
R169 VTAIL.n218 VTAIL.n217 104.615
R170 VTAIL.n218 VTAIL.n207 104.615
R171 VTAIL.n225 VTAIL.n207 104.615
R172 VTAIL.n226 VTAIL.n225 104.615
R173 VTAIL.n15 VTAIL.n9 104.615
R174 VTAIL.n16 VTAIL.n15 104.615
R175 VTAIL.n16 VTAIL.n5 104.615
R176 VTAIL.n23 VTAIL.n5 104.615
R177 VTAIL.n24 VTAIL.n23 104.615
R178 VTAIL.n43 VTAIL.n37 104.615
R179 VTAIL.n44 VTAIL.n43 104.615
R180 VTAIL.n44 VTAIL.n33 104.615
R181 VTAIL.n51 VTAIL.n33 104.615
R182 VTAIL.n52 VTAIL.n51 104.615
R183 VTAIL.n73 VTAIL.n67 104.615
R184 VTAIL.n74 VTAIL.n73 104.615
R185 VTAIL.n74 VTAIL.n63 104.615
R186 VTAIL.n81 VTAIL.n63 104.615
R187 VTAIL.n82 VTAIL.n81 104.615
R188 VTAIL.n198 VTAIL.n197 104.615
R189 VTAIL.n197 VTAIL.n179 104.615
R190 VTAIL.n190 VTAIL.n179 104.615
R191 VTAIL.n190 VTAIL.n189 104.615
R192 VTAIL.n189 VTAIL.n183 104.615
R193 VTAIL.n168 VTAIL.n167 104.615
R194 VTAIL.n167 VTAIL.n149 104.615
R195 VTAIL.n160 VTAIL.n149 104.615
R196 VTAIL.n160 VTAIL.n159 104.615
R197 VTAIL.n159 VTAIL.n153 104.615
R198 VTAIL.n140 VTAIL.n139 104.615
R199 VTAIL.n139 VTAIL.n121 104.615
R200 VTAIL.n132 VTAIL.n121 104.615
R201 VTAIL.n132 VTAIL.n131 104.615
R202 VTAIL.n131 VTAIL.n125 104.615
R203 VTAIL.n110 VTAIL.n109 104.615
R204 VTAIL.n109 VTAIL.n91 104.615
R205 VTAIL.n102 VTAIL.n91 104.615
R206 VTAIL.n102 VTAIL.n101 104.615
R207 VTAIL.n101 VTAIL.n95 104.615
R208 VTAIL.n175 VTAIL.n174 52.7522
R209 VTAIL.n117 VTAIL.n116 52.7522
R210 VTAIL.n1 VTAIL.n0 52.7521
R211 VTAIL.n59 VTAIL.n58 52.7521
R212 VTAIL.t0 VTAIL.n211 52.3082
R213 VTAIL.t4 VTAIL.n9 52.3082
R214 VTAIL.t11 VTAIL.n37 52.3082
R215 VTAIL.t10 VTAIL.n67 52.3082
R216 VTAIL.t12 VTAIL.n183 52.3082
R217 VTAIL.t15 VTAIL.n153 52.3082
R218 VTAIL.t6 VTAIL.n125 52.3082
R219 VTAIL.t3 VTAIL.n95 52.3082
R220 VTAIL.n231 VTAIL.n230 32.9611
R221 VTAIL.n29 VTAIL.n28 32.9611
R222 VTAIL.n57 VTAIL.n56 32.9611
R223 VTAIL.n87 VTAIL.n86 32.9611
R224 VTAIL.n203 VTAIL.n202 32.9611
R225 VTAIL.n173 VTAIL.n172 32.9611
R226 VTAIL.n145 VTAIL.n144 32.9611
R227 VTAIL.n115 VTAIL.n114 32.9611
R228 VTAIL.n231 VTAIL.n203 18.8324
R229 VTAIL.n115 VTAIL.n87 18.8324
R230 VTAIL.n213 VTAIL.n212 15.6666
R231 VTAIL.n11 VTAIL.n10 15.6666
R232 VTAIL.n39 VTAIL.n38 15.6666
R233 VTAIL.n69 VTAIL.n68 15.6666
R234 VTAIL.n185 VTAIL.n184 15.6666
R235 VTAIL.n155 VTAIL.n154 15.6666
R236 VTAIL.n127 VTAIL.n126 15.6666
R237 VTAIL.n97 VTAIL.n96 15.6666
R238 VTAIL.n216 VTAIL.n215 12.8005
R239 VTAIL.n14 VTAIL.n13 12.8005
R240 VTAIL.n42 VTAIL.n41 12.8005
R241 VTAIL.n72 VTAIL.n71 12.8005
R242 VTAIL.n188 VTAIL.n187 12.8005
R243 VTAIL.n158 VTAIL.n157 12.8005
R244 VTAIL.n130 VTAIL.n129 12.8005
R245 VTAIL.n100 VTAIL.n99 12.8005
R246 VTAIL.n219 VTAIL.n210 12.0247
R247 VTAIL.n17 VTAIL.n8 12.0247
R248 VTAIL.n45 VTAIL.n36 12.0247
R249 VTAIL.n75 VTAIL.n66 12.0247
R250 VTAIL.n191 VTAIL.n182 12.0247
R251 VTAIL.n161 VTAIL.n152 12.0247
R252 VTAIL.n133 VTAIL.n124 12.0247
R253 VTAIL.n103 VTAIL.n94 12.0247
R254 VTAIL.n220 VTAIL.n208 11.249
R255 VTAIL.n18 VTAIL.n6 11.249
R256 VTAIL.n46 VTAIL.n34 11.249
R257 VTAIL.n76 VTAIL.n64 11.249
R258 VTAIL.n192 VTAIL.n180 11.249
R259 VTAIL.n162 VTAIL.n150 11.249
R260 VTAIL.n134 VTAIL.n122 11.249
R261 VTAIL.n104 VTAIL.n92 11.249
R262 VTAIL.n224 VTAIL.n223 10.4732
R263 VTAIL.n22 VTAIL.n21 10.4732
R264 VTAIL.n50 VTAIL.n49 10.4732
R265 VTAIL.n80 VTAIL.n79 10.4732
R266 VTAIL.n196 VTAIL.n195 10.4732
R267 VTAIL.n166 VTAIL.n165 10.4732
R268 VTAIL.n138 VTAIL.n137 10.4732
R269 VTAIL.n108 VTAIL.n107 10.4732
R270 VTAIL.n227 VTAIL.n206 9.69747
R271 VTAIL.n25 VTAIL.n4 9.69747
R272 VTAIL.n53 VTAIL.n32 9.69747
R273 VTAIL.n83 VTAIL.n62 9.69747
R274 VTAIL.n199 VTAIL.n178 9.69747
R275 VTAIL.n169 VTAIL.n148 9.69747
R276 VTAIL.n141 VTAIL.n120 9.69747
R277 VTAIL.n111 VTAIL.n90 9.69747
R278 VTAIL.n230 VTAIL.n229 9.45567
R279 VTAIL.n28 VTAIL.n27 9.45567
R280 VTAIL.n56 VTAIL.n55 9.45567
R281 VTAIL.n86 VTAIL.n85 9.45567
R282 VTAIL.n202 VTAIL.n201 9.45567
R283 VTAIL.n172 VTAIL.n171 9.45567
R284 VTAIL.n144 VTAIL.n143 9.45567
R285 VTAIL.n114 VTAIL.n113 9.45567
R286 VTAIL.n229 VTAIL.n228 9.3005
R287 VTAIL.n206 VTAIL.n205 9.3005
R288 VTAIL.n223 VTAIL.n222 9.3005
R289 VTAIL.n221 VTAIL.n220 9.3005
R290 VTAIL.n210 VTAIL.n209 9.3005
R291 VTAIL.n215 VTAIL.n214 9.3005
R292 VTAIL.n27 VTAIL.n26 9.3005
R293 VTAIL.n4 VTAIL.n3 9.3005
R294 VTAIL.n21 VTAIL.n20 9.3005
R295 VTAIL.n19 VTAIL.n18 9.3005
R296 VTAIL.n8 VTAIL.n7 9.3005
R297 VTAIL.n13 VTAIL.n12 9.3005
R298 VTAIL.n55 VTAIL.n54 9.3005
R299 VTAIL.n32 VTAIL.n31 9.3005
R300 VTAIL.n49 VTAIL.n48 9.3005
R301 VTAIL.n47 VTAIL.n46 9.3005
R302 VTAIL.n36 VTAIL.n35 9.3005
R303 VTAIL.n41 VTAIL.n40 9.3005
R304 VTAIL.n85 VTAIL.n84 9.3005
R305 VTAIL.n62 VTAIL.n61 9.3005
R306 VTAIL.n79 VTAIL.n78 9.3005
R307 VTAIL.n77 VTAIL.n76 9.3005
R308 VTAIL.n66 VTAIL.n65 9.3005
R309 VTAIL.n71 VTAIL.n70 9.3005
R310 VTAIL.n201 VTAIL.n200 9.3005
R311 VTAIL.n178 VTAIL.n177 9.3005
R312 VTAIL.n195 VTAIL.n194 9.3005
R313 VTAIL.n193 VTAIL.n192 9.3005
R314 VTAIL.n182 VTAIL.n181 9.3005
R315 VTAIL.n187 VTAIL.n186 9.3005
R316 VTAIL.n171 VTAIL.n170 9.3005
R317 VTAIL.n148 VTAIL.n147 9.3005
R318 VTAIL.n165 VTAIL.n164 9.3005
R319 VTAIL.n163 VTAIL.n162 9.3005
R320 VTAIL.n152 VTAIL.n151 9.3005
R321 VTAIL.n157 VTAIL.n156 9.3005
R322 VTAIL.n143 VTAIL.n142 9.3005
R323 VTAIL.n120 VTAIL.n119 9.3005
R324 VTAIL.n137 VTAIL.n136 9.3005
R325 VTAIL.n135 VTAIL.n134 9.3005
R326 VTAIL.n124 VTAIL.n123 9.3005
R327 VTAIL.n129 VTAIL.n128 9.3005
R328 VTAIL.n113 VTAIL.n112 9.3005
R329 VTAIL.n90 VTAIL.n89 9.3005
R330 VTAIL.n107 VTAIL.n106 9.3005
R331 VTAIL.n105 VTAIL.n104 9.3005
R332 VTAIL.n94 VTAIL.n93 9.3005
R333 VTAIL.n99 VTAIL.n98 9.3005
R334 VTAIL.n228 VTAIL.n204 8.92171
R335 VTAIL.n26 VTAIL.n2 8.92171
R336 VTAIL.n54 VTAIL.n30 8.92171
R337 VTAIL.n84 VTAIL.n60 8.92171
R338 VTAIL.n200 VTAIL.n176 8.92171
R339 VTAIL.n170 VTAIL.n146 8.92171
R340 VTAIL.n142 VTAIL.n118 8.92171
R341 VTAIL.n112 VTAIL.n88 8.92171
R342 VTAIL.n230 VTAIL.n204 5.04292
R343 VTAIL.n28 VTAIL.n2 5.04292
R344 VTAIL.n56 VTAIL.n30 5.04292
R345 VTAIL.n86 VTAIL.n60 5.04292
R346 VTAIL.n202 VTAIL.n176 5.04292
R347 VTAIL.n172 VTAIL.n146 5.04292
R348 VTAIL.n144 VTAIL.n118 5.04292
R349 VTAIL.n114 VTAIL.n88 5.04292
R350 VTAIL.n214 VTAIL.n213 4.38687
R351 VTAIL.n12 VTAIL.n11 4.38687
R352 VTAIL.n40 VTAIL.n39 4.38687
R353 VTAIL.n70 VTAIL.n69 4.38687
R354 VTAIL.n186 VTAIL.n185 4.38687
R355 VTAIL.n156 VTAIL.n155 4.38687
R356 VTAIL.n128 VTAIL.n127 4.38687
R357 VTAIL.n98 VTAIL.n97 4.38687
R358 VTAIL.n228 VTAIL.n227 4.26717
R359 VTAIL.n26 VTAIL.n25 4.26717
R360 VTAIL.n54 VTAIL.n53 4.26717
R361 VTAIL.n84 VTAIL.n83 4.26717
R362 VTAIL.n200 VTAIL.n199 4.26717
R363 VTAIL.n170 VTAIL.n169 4.26717
R364 VTAIL.n142 VTAIL.n141 4.26717
R365 VTAIL.n112 VTAIL.n111 4.26717
R366 VTAIL.n0 VTAIL.t7 3.7223
R367 VTAIL.n0 VTAIL.t2 3.7223
R368 VTAIL.n58 VTAIL.t8 3.7223
R369 VTAIL.n58 VTAIL.t9 3.7223
R370 VTAIL.n174 VTAIL.t13 3.7223
R371 VTAIL.n174 VTAIL.t14 3.7223
R372 VTAIL.n116 VTAIL.t5 3.7223
R373 VTAIL.n116 VTAIL.t1 3.7223
R374 VTAIL.n224 VTAIL.n206 3.49141
R375 VTAIL.n22 VTAIL.n4 3.49141
R376 VTAIL.n50 VTAIL.n32 3.49141
R377 VTAIL.n80 VTAIL.n62 3.49141
R378 VTAIL.n196 VTAIL.n178 3.49141
R379 VTAIL.n166 VTAIL.n148 3.49141
R380 VTAIL.n138 VTAIL.n120 3.49141
R381 VTAIL.n108 VTAIL.n90 3.49141
R382 VTAIL.n223 VTAIL.n208 2.71565
R383 VTAIL.n21 VTAIL.n6 2.71565
R384 VTAIL.n49 VTAIL.n34 2.71565
R385 VTAIL.n79 VTAIL.n64 2.71565
R386 VTAIL.n195 VTAIL.n180 2.71565
R387 VTAIL.n165 VTAIL.n150 2.71565
R388 VTAIL.n137 VTAIL.n122 2.71565
R389 VTAIL.n107 VTAIL.n92 2.71565
R390 VTAIL.n220 VTAIL.n219 1.93989
R391 VTAIL.n18 VTAIL.n17 1.93989
R392 VTAIL.n46 VTAIL.n45 1.93989
R393 VTAIL.n76 VTAIL.n75 1.93989
R394 VTAIL.n192 VTAIL.n191 1.93989
R395 VTAIL.n162 VTAIL.n161 1.93989
R396 VTAIL.n134 VTAIL.n133 1.93989
R397 VTAIL.n104 VTAIL.n103 1.93989
R398 VTAIL.n117 VTAIL.n115 1.87981
R399 VTAIL.n145 VTAIL.n117 1.87981
R400 VTAIL.n175 VTAIL.n173 1.87981
R401 VTAIL.n203 VTAIL.n175 1.87981
R402 VTAIL.n87 VTAIL.n59 1.87981
R403 VTAIL.n59 VTAIL.n57 1.87981
R404 VTAIL.n29 VTAIL.n1 1.87981
R405 VTAIL VTAIL.n231 1.82162
R406 VTAIL.n216 VTAIL.n210 1.16414
R407 VTAIL.n14 VTAIL.n8 1.16414
R408 VTAIL.n42 VTAIL.n36 1.16414
R409 VTAIL.n72 VTAIL.n66 1.16414
R410 VTAIL.n188 VTAIL.n182 1.16414
R411 VTAIL.n158 VTAIL.n152 1.16414
R412 VTAIL.n130 VTAIL.n124 1.16414
R413 VTAIL.n100 VTAIL.n94 1.16414
R414 VTAIL.n173 VTAIL.n145 0.470328
R415 VTAIL.n57 VTAIL.n29 0.470328
R416 VTAIL.n215 VTAIL.n212 0.388379
R417 VTAIL.n13 VTAIL.n10 0.388379
R418 VTAIL.n41 VTAIL.n38 0.388379
R419 VTAIL.n71 VTAIL.n68 0.388379
R420 VTAIL.n187 VTAIL.n184 0.388379
R421 VTAIL.n157 VTAIL.n154 0.388379
R422 VTAIL.n129 VTAIL.n126 0.388379
R423 VTAIL.n99 VTAIL.n96 0.388379
R424 VTAIL.n214 VTAIL.n209 0.155672
R425 VTAIL.n221 VTAIL.n209 0.155672
R426 VTAIL.n222 VTAIL.n221 0.155672
R427 VTAIL.n222 VTAIL.n205 0.155672
R428 VTAIL.n229 VTAIL.n205 0.155672
R429 VTAIL.n12 VTAIL.n7 0.155672
R430 VTAIL.n19 VTAIL.n7 0.155672
R431 VTAIL.n20 VTAIL.n19 0.155672
R432 VTAIL.n20 VTAIL.n3 0.155672
R433 VTAIL.n27 VTAIL.n3 0.155672
R434 VTAIL.n40 VTAIL.n35 0.155672
R435 VTAIL.n47 VTAIL.n35 0.155672
R436 VTAIL.n48 VTAIL.n47 0.155672
R437 VTAIL.n48 VTAIL.n31 0.155672
R438 VTAIL.n55 VTAIL.n31 0.155672
R439 VTAIL.n70 VTAIL.n65 0.155672
R440 VTAIL.n77 VTAIL.n65 0.155672
R441 VTAIL.n78 VTAIL.n77 0.155672
R442 VTAIL.n78 VTAIL.n61 0.155672
R443 VTAIL.n85 VTAIL.n61 0.155672
R444 VTAIL.n201 VTAIL.n177 0.155672
R445 VTAIL.n194 VTAIL.n177 0.155672
R446 VTAIL.n194 VTAIL.n193 0.155672
R447 VTAIL.n193 VTAIL.n181 0.155672
R448 VTAIL.n186 VTAIL.n181 0.155672
R449 VTAIL.n171 VTAIL.n147 0.155672
R450 VTAIL.n164 VTAIL.n147 0.155672
R451 VTAIL.n164 VTAIL.n163 0.155672
R452 VTAIL.n163 VTAIL.n151 0.155672
R453 VTAIL.n156 VTAIL.n151 0.155672
R454 VTAIL.n143 VTAIL.n119 0.155672
R455 VTAIL.n136 VTAIL.n119 0.155672
R456 VTAIL.n136 VTAIL.n135 0.155672
R457 VTAIL.n135 VTAIL.n123 0.155672
R458 VTAIL.n128 VTAIL.n123 0.155672
R459 VTAIL.n113 VTAIL.n89 0.155672
R460 VTAIL.n106 VTAIL.n89 0.155672
R461 VTAIL.n106 VTAIL.n105 0.155672
R462 VTAIL.n105 VTAIL.n93 0.155672
R463 VTAIL.n98 VTAIL.n93 0.155672
R464 VTAIL VTAIL.n1 0.0586897
R465 B.n598 B.n597 585
R466 B.n599 B.n598 585
R467 B.n209 B.n102 585
R468 B.n208 B.n207 585
R469 B.n206 B.n205 585
R470 B.n204 B.n203 585
R471 B.n202 B.n201 585
R472 B.n200 B.n199 585
R473 B.n198 B.n197 585
R474 B.n196 B.n195 585
R475 B.n194 B.n193 585
R476 B.n192 B.n191 585
R477 B.n190 B.n189 585
R478 B.n188 B.n187 585
R479 B.n186 B.n185 585
R480 B.n184 B.n183 585
R481 B.n182 B.n181 585
R482 B.n180 B.n179 585
R483 B.n178 B.n177 585
R484 B.n176 B.n175 585
R485 B.n174 B.n173 585
R486 B.n172 B.n171 585
R487 B.n170 B.n169 585
R488 B.n167 B.n166 585
R489 B.n165 B.n164 585
R490 B.n163 B.n162 585
R491 B.n161 B.n160 585
R492 B.n159 B.n158 585
R493 B.n157 B.n156 585
R494 B.n155 B.n154 585
R495 B.n153 B.n152 585
R496 B.n151 B.n150 585
R497 B.n149 B.n148 585
R498 B.n147 B.n146 585
R499 B.n145 B.n144 585
R500 B.n143 B.n142 585
R501 B.n141 B.n140 585
R502 B.n139 B.n138 585
R503 B.n137 B.n136 585
R504 B.n135 B.n134 585
R505 B.n133 B.n132 585
R506 B.n131 B.n130 585
R507 B.n129 B.n128 585
R508 B.n127 B.n126 585
R509 B.n125 B.n124 585
R510 B.n123 B.n122 585
R511 B.n121 B.n120 585
R512 B.n119 B.n118 585
R513 B.n117 B.n116 585
R514 B.n115 B.n114 585
R515 B.n113 B.n112 585
R516 B.n111 B.n110 585
R517 B.n109 B.n108 585
R518 B.n74 B.n73 585
R519 B.n596 B.n75 585
R520 B.n600 B.n75 585
R521 B.n595 B.n594 585
R522 B.n594 B.n71 585
R523 B.n593 B.n70 585
R524 B.n606 B.n70 585
R525 B.n592 B.n69 585
R526 B.n607 B.n69 585
R527 B.n591 B.n68 585
R528 B.n608 B.n68 585
R529 B.n590 B.n589 585
R530 B.n589 B.n64 585
R531 B.n588 B.n63 585
R532 B.n614 B.n63 585
R533 B.n587 B.n62 585
R534 B.n615 B.n62 585
R535 B.n586 B.n61 585
R536 B.n616 B.n61 585
R537 B.n585 B.n584 585
R538 B.n584 B.n57 585
R539 B.n583 B.n56 585
R540 B.n622 B.n56 585
R541 B.n582 B.n55 585
R542 B.n623 B.n55 585
R543 B.n581 B.n54 585
R544 B.n624 B.n54 585
R545 B.n580 B.n579 585
R546 B.n579 B.n50 585
R547 B.n578 B.n49 585
R548 B.n630 B.n49 585
R549 B.n577 B.n48 585
R550 B.n631 B.n48 585
R551 B.n576 B.n47 585
R552 B.n632 B.n47 585
R553 B.n575 B.n574 585
R554 B.n574 B.n43 585
R555 B.n573 B.n42 585
R556 B.n638 B.n42 585
R557 B.n572 B.n41 585
R558 B.n639 B.n41 585
R559 B.n571 B.n40 585
R560 B.n640 B.n40 585
R561 B.n570 B.n569 585
R562 B.n569 B.n36 585
R563 B.n568 B.n35 585
R564 B.n646 B.n35 585
R565 B.n567 B.n34 585
R566 B.n647 B.n34 585
R567 B.n566 B.n33 585
R568 B.n648 B.n33 585
R569 B.n565 B.n564 585
R570 B.n564 B.n29 585
R571 B.n563 B.n28 585
R572 B.n654 B.n28 585
R573 B.n562 B.n27 585
R574 B.n655 B.n27 585
R575 B.n561 B.n26 585
R576 B.n656 B.n26 585
R577 B.n560 B.n559 585
R578 B.n559 B.n22 585
R579 B.n558 B.n21 585
R580 B.n662 B.n21 585
R581 B.n557 B.n20 585
R582 B.n663 B.n20 585
R583 B.n556 B.n19 585
R584 B.n664 B.n19 585
R585 B.n555 B.n554 585
R586 B.n554 B.n15 585
R587 B.n553 B.n14 585
R588 B.n670 B.n14 585
R589 B.n552 B.n13 585
R590 B.n671 B.n13 585
R591 B.n551 B.n12 585
R592 B.n672 B.n12 585
R593 B.n550 B.n549 585
R594 B.n549 B.n8 585
R595 B.n548 B.n7 585
R596 B.n678 B.n7 585
R597 B.n547 B.n6 585
R598 B.n679 B.n6 585
R599 B.n546 B.n5 585
R600 B.n680 B.n5 585
R601 B.n545 B.n544 585
R602 B.n544 B.n4 585
R603 B.n543 B.n210 585
R604 B.n543 B.n542 585
R605 B.n533 B.n211 585
R606 B.n212 B.n211 585
R607 B.n535 B.n534 585
R608 B.n536 B.n535 585
R609 B.n532 B.n216 585
R610 B.n220 B.n216 585
R611 B.n531 B.n530 585
R612 B.n530 B.n529 585
R613 B.n218 B.n217 585
R614 B.n219 B.n218 585
R615 B.n522 B.n521 585
R616 B.n523 B.n522 585
R617 B.n520 B.n225 585
R618 B.n225 B.n224 585
R619 B.n519 B.n518 585
R620 B.n518 B.n517 585
R621 B.n227 B.n226 585
R622 B.n228 B.n227 585
R623 B.n510 B.n509 585
R624 B.n511 B.n510 585
R625 B.n508 B.n233 585
R626 B.n233 B.n232 585
R627 B.n507 B.n506 585
R628 B.n506 B.n505 585
R629 B.n235 B.n234 585
R630 B.n236 B.n235 585
R631 B.n498 B.n497 585
R632 B.n499 B.n498 585
R633 B.n496 B.n241 585
R634 B.n241 B.n240 585
R635 B.n495 B.n494 585
R636 B.n494 B.n493 585
R637 B.n243 B.n242 585
R638 B.n244 B.n243 585
R639 B.n486 B.n485 585
R640 B.n487 B.n486 585
R641 B.n484 B.n249 585
R642 B.n249 B.n248 585
R643 B.n483 B.n482 585
R644 B.n482 B.n481 585
R645 B.n251 B.n250 585
R646 B.n252 B.n251 585
R647 B.n474 B.n473 585
R648 B.n475 B.n474 585
R649 B.n472 B.n256 585
R650 B.n260 B.n256 585
R651 B.n471 B.n470 585
R652 B.n470 B.n469 585
R653 B.n258 B.n257 585
R654 B.n259 B.n258 585
R655 B.n462 B.n461 585
R656 B.n463 B.n462 585
R657 B.n460 B.n265 585
R658 B.n265 B.n264 585
R659 B.n459 B.n458 585
R660 B.n458 B.n457 585
R661 B.n267 B.n266 585
R662 B.n268 B.n267 585
R663 B.n450 B.n449 585
R664 B.n451 B.n450 585
R665 B.n448 B.n273 585
R666 B.n273 B.n272 585
R667 B.n447 B.n446 585
R668 B.n446 B.n445 585
R669 B.n275 B.n274 585
R670 B.n276 B.n275 585
R671 B.n438 B.n437 585
R672 B.n439 B.n438 585
R673 B.n436 B.n281 585
R674 B.n281 B.n280 585
R675 B.n435 B.n434 585
R676 B.n434 B.n433 585
R677 B.n283 B.n282 585
R678 B.n284 B.n283 585
R679 B.n426 B.n425 585
R680 B.n427 B.n426 585
R681 B.n287 B.n286 585
R682 B.n320 B.n318 585
R683 B.n321 B.n317 585
R684 B.n321 B.n288 585
R685 B.n324 B.n323 585
R686 B.n325 B.n316 585
R687 B.n327 B.n326 585
R688 B.n329 B.n315 585
R689 B.n332 B.n331 585
R690 B.n333 B.n314 585
R691 B.n335 B.n334 585
R692 B.n337 B.n313 585
R693 B.n340 B.n339 585
R694 B.n341 B.n312 585
R695 B.n343 B.n342 585
R696 B.n345 B.n311 585
R697 B.n348 B.n347 585
R698 B.n349 B.n310 585
R699 B.n351 B.n350 585
R700 B.n353 B.n309 585
R701 B.n356 B.n355 585
R702 B.n357 B.n308 585
R703 B.n362 B.n361 585
R704 B.n364 B.n307 585
R705 B.n367 B.n366 585
R706 B.n368 B.n306 585
R707 B.n370 B.n369 585
R708 B.n372 B.n305 585
R709 B.n375 B.n374 585
R710 B.n376 B.n304 585
R711 B.n378 B.n377 585
R712 B.n380 B.n303 585
R713 B.n383 B.n382 585
R714 B.n384 B.n299 585
R715 B.n386 B.n385 585
R716 B.n388 B.n298 585
R717 B.n391 B.n390 585
R718 B.n392 B.n297 585
R719 B.n394 B.n393 585
R720 B.n396 B.n296 585
R721 B.n399 B.n398 585
R722 B.n400 B.n295 585
R723 B.n402 B.n401 585
R724 B.n404 B.n294 585
R725 B.n407 B.n406 585
R726 B.n408 B.n293 585
R727 B.n410 B.n409 585
R728 B.n412 B.n292 585
R729 B.n415 B.n414 585
R730 B.n416 B.n291 585
R731 B.n418 B.n417 585
R732 B.n420 B.n290 585
R733 B.n423 B.n422 585
R734 B.n424 B.n289 585
R735 B.n429 B.n428 585
R736 B.n428 B.n427 585
R737 B.n430 B.n285 585
R738 B.n285 B.n284 585
R739 B.n432 B.n431 585
R740 B.n433 B.n432 585
R741 B.n279 B.n278 585
R742 B.n280 B.n279 585
R743 B.n441 B.n440 585
R744 B.n440 B.n439 585
R745 B.n442 B.n277 585
R746 B.n277 B.n276 585
R747 B.n444 B.n443 585
R748 B.n445 B.n444 585
R749 B.n271 B.n270 585
R750 B.n272 B.n271 585
R751 B.n453 B.n452 585
R752 B.n452 B.n451 585
R753 B.n454 B.n269 585
R754 B.n269 B.n268 585
R755 B.n456 B.n455 585
R756 B.n457 B.n456 585
R757 B.n263 B.n262 585
R758 B.n264 B.n263 585
R759 B.n465 B.n464 585
R760 B.n464 B.n463 585
R761 B.n466 B.n261 585
R762 B.n261 B.n259 585
R763 B.n468 B.n467 585
R764 B.n469 B.n468 585
R765 B.n255 B.n254 585
R766 B.n260 B.n255 585
R767 B.n477 B.n476 585
R768 B.n476 B.n475 585
R769 B.n478 B.n253 585
R770 B.n253 B.n252 585
R771 B.n480 B.n479 585
R772 B.n481 B.n480 585
R773 B.n247 B.n246 585
R774 B.n248 B.n247 585
R775 B.n489 B.n488 585
R776 B.n488 B.n487 585
R777 B.n490 B.n245 585
R778 B.n245 B.n244 585
R779 B.n492 B.n491 585
R780 B.n493 B.n492 585
R781 B.n239 B.n238 585
R782 B.n240 B.n239 585
R783 B.n501 B.n500 585
R784 B.n500 B.n499 585
R785 B.n502 B.n237 585
R786 B.n237 B.n236 585
R787 B.n504 B.n503 585
R788 B.n505 B.n504 585
R789 B.n231 B.n230 585
R790 B.n232 B.n231 585
R791 B.n513 B.n512 585
R792 B.n512 B.n511 585
R793 B.n514 B.n229 585
R794 B.n229 B.n228 585
R795 B.n516 B.n515 585
R796 B.n517 B.n516 585
R797 B.n223 B.n222 585
R798 B.n224 B.n223 585
R799 B.n525 B.n524 585
R800 B.n524 B.n523 585
R801 B.n526 B.n221 585
R802 B.n221 B.n219 585
R803 B.n528 B.n527 585
R804 B.n529 B.n528 585
R805 B.n215 B.n214 585
R806 B.n220 B.n215 585
R807 B.n538 B.n537 585
R808 B.n537 B.n536 585
R809 B.n539 B.n213 585
R810 B.n213 B.n212 585
R811 B.n541 B.n540 585
R812 B.n542 B.n541 585
R813 B.n2 B.n0 585
R814 B.n4 B.n2 585
R815 B.n3 B.n1 585
R816 B.n679 B.n3 585
R817 B.n677 B.n676 585
R818 B.n678 B.n677 585
R819 B.n675 B.n9 585
R820 B.n9 B.n8 585
R821 B.n674 B.n673 585
R822 B.n673 B.n672 585
R823 B.n11 B.n10 585
R824 B.n671 B.n11 585
R825 B.n669 B.n668 585
R826 B.n670 B.n669 585
R827 B.n667 B.n16 585
R828 B.n16 B.n15 585
R829 B.n666 B.n665 585
R830 B.n665 B.n664 585
R831 B.n18 B.n17 585
R832 B.n663 B.n18 585
R833 B.n661 B.n660 585
R834 B.n662 B.n661 585
R835 B.n659 B.n23 585
R836 B.n23 B.n22 585
R837 B.n658 B.n657 585
R838 B.n657 B.n656 585
R839 B.n25 B.n24 585
R840 B.n655 B.n25 585
R841 B.n653 B.n652 585
R842 B.n654 B.n653 585
R843 B.n651 B.n30 585
R844 B.n30 B.n29 585
R845 B.n650 B.n649 585
R846 B.n649 B.n648 585
R847 B.n32 B.n31 585
R848 B.n647 B.n32 585
R849 B.n645 B.n644 585
R850 B.n646 B.n645 585
R851 B.n643 B.n37 585
R852 B.n37 B.n36 585
R853 B.n642 B.n641 585
R854 B.n641 B.n640 585
R855 B.n39 B.n38 585
R856 B.n639 B.n39 585
R857 B.n637 B.n636 585
R858 B.n638 B.n637 585
R859 B.n635 B.n44 585
R860 B.n44 B.n43 585
R861 B.n634 B.n633 585
R862 B.n633 B.n632 585
R863 B.n46 B.n45 585
R864 B.n631 B.n46 585
R865 B.n629 B.n628 585
R866 B.n630 B.n629 585
R867 B.n627 B.n51 585
R868 B.n51 B.n50 585
R869 B.n626 B.n625 585
R870 B.n625 B.n624 585
R871 B.n53 B.n52 585
R872 B.n623 B.n53 585
R873 B.n621 B.n620 585
R874 B.n622 B.n621 585
R875 B.n619 B.n58 585
R876 B.n58 B.n57 585
R877 B.n618 B.n617 585
R878 B.n617 B.n616 585
R879 B.n60 B.n59 585
R880 B.n615 B.n60 585
R881 B.n613 B.n612 585
R882 B.n614 B.n613 585
R883 B.n611 B.n65 585
R884 B.n65 B.n64 585
R885 B.n610 B.n609 585
R886 B.n609 B.n608 585
R887 B.n67 B.n66 585
R888 B.n607 B.n67 585
R889 B.n605 B.n604 585
R890 B.n606 B.n605 585
R891 B.n603 B.n72 585
R892 B.n72 B.n71 585
R893 B.n602 B.n601 585
R894 B.n601 B.n600 585
R895 B.n682 B.n681 585
R896 B.n681 B.n680 585
R897 B.n428 B.n287 569.379
R898 B.n601 B.n74 569.379
R899 B.n426 B.n289 569.379
R900 B.n598 B.n75 569.379
R901 B.n300 B.t8 275.846
R902 B.n358 B.t16 275.846
R903 B.n105 B.t12 275.846
R904 B.n103 B.t19 275.846
R905 B.n599 B.n101 256.663
R906 B.n599 B.n100 256.663
R907 B.n599 B.n99 256.663
R908 B.n599 B.n98 256.663
R909 B.n599 B.n97 256.663
R910 B.n599 B.n96 256.663
R911 B.n599 B.n95 256.663
R912 B.n599 B.n94 256.663
R913 B.n599 B.n93 256.663
R914 B.n599 B.n92 256.663
R915 B.n599 B.n91 256.663
R916 B.n599 B.n90 256.663
R917 B.n599 B.n89 256.663
R918 B.n599 B.n88 256.663
R919 B.n599 B.n87 256.663
R920 B.n599 B.n86 256.663
R921 B.n599 B.n85 256.663
R922 B.n599 B.n84 256.663
R923 B.n599 B.n83 256.663
R924 B.n599 B.n82 256.663
R925 B.n599 B.n81 256.663
R926 B.n599 B.n80 256.663
R927 B.n599 B.n79 256.663
R928 B.n599 B.n78 256.663
R929 B.n599 B.n77 256.663
R930 B.n599 B.n76 256.663
R931 B.n319 B.n288 256.663
R932 B.n322 B.n288 256.663
R933 B.n328 B.n288 256.663
R934 B.n330 B.n288 256.663
R935 B.n336 B.n288 256.663
R936 B.n338 B.n288 256.663
R937 B.n344 B.n288 256.663
R938 B.n346 B.n288 256.663
R939 B.n352 B.n288 256.663
R940 B.n354 B.n288 256.663
R941 B.n363 B.n288 256.663
R942 B.n365 B.n288 256.663
R943 B.n371 B.n288 256.663
R944 B.n373 B.n288 256.663
R945 B.n379 B.n288 256.663
R946 B.n381 B.n288 256.663
R947 B.n387 B.n288 256.663
R948 B.n389 B.n288 256.663
R949 B.n395 B.n288 256.663
R950 B.n397 B.n288 256.663
R951 B.n403 B.n288 256.663
R952 B.n405 B.n288 256.663
R953 B.n411 B.n288 256.663
R954 B.n413 B.n288 256.663
R955 B.n419 B.n288 256.663
R956 B.n421 B.n288 256.663
R957 B.n300 B.t11 209.629
R958 B.n103 B.t20 209.629
R959 B.n358 B.t18 209.629
R960 B.n105 B.t14 209.629
R961 B.n301 B.t10 167.35
R962 B.n104 B.t21 167.35
R963 B.n359 B.t17 167.35
R964 B.n106 B.t15 167.35
R965 B.n428 B.n285 163.367
R966 B.n432 B.n285 163.367
R967 B.n432 B.n279 163.367
R968 B.n440 B.n279 163.367
R969 B.n440 B.n277 163.367
R970 B.n444 B.n277 163.367
R971 B.n444 B.n271 163.367
R972 B.n452 B.n271 163.367
R973 B.n452 B.n269 163.367
R974 B.n456 B.n269 163.367
R975 B.n456 B.n263 163.367
R976 B.n464 B.n263 163.367
R977 B.n464 B.n261 163.367
R978 B.n468 B.n261 163.367
R979 B.n468 B.n255 163.367
R980 B.n476 B.n255 163.367
R981 B.n476 B.n253 163.367
R982 B.n480 B.n253 163.367
R983 B.n480 B.n247 163.367
R984 B.n488 B.n247 163.367
R985 B.n488 B.n245 163.367
R986 B.n492 B.n245 163.367
R987 B.n492 B.n239 163.367
R988 B.n500 B.n239 163.367
R989 B.n500 B.n237 163.367
R990 B.n504 B.n237 163.367
R991 B.n504 B.n231 163.367
R992 B.n512 B.n231 163.367
R993 B.n512 B.n229 163.367
R994 B.n516 B.n229 163.367
R995 B.n516 B.n223 163.367
R996 B.n524 B.n223 163.367
R997 B.n524 B.n221 163.367
R998 B.n528 B.n221 163.367
R999 B.n528 B.n215 163.367
R1000 B.n537 B.n215 163.367
R1001 B.n537 B.n213 163.367
R1002 B.n541 B.n213 163.367
R1003 B.n541 B.n2 163.367
R1004 B.n681 B.n2 163.367
R1005 B.n681 B.n3 163.367
R1006 B.n677 B.n3 163.367
R1007 B.n677 B.n9 163.367
R1008 B.n673 B.n9 163.367
R1009 B.n673 B.n11 163.367
R1010 B.n669 B.n11 163.367
R1011 B.n669 B.n16 163.367
R1012 B.n665 B.n16 163.367
R1013 B.n665 B.n18 163.367
R1014 B.n661 B.n18 163.367
R1015 B.n661 B.n23 163.367
R1016 B.n657 B.n23 163.367
R1017 B.n657 B.n25 163.367
R1018 B.n653 B.n25 163.367
R1019 B.n653 B.n30 163.367
R1020 B.n649 B.n30 163.367
R1021 B.n649 B.n32 163.367
R1022 B.n645 B.n32 163.367
R1023 B.n645 B.n37 163.367
R1024 B.n641 B.n37 163.367
R1025 B.n641 B.n39 163.367
R1026 B.n637 B.n39 163.367
R1027 B.n637 B.n44 163.367
R1028 B.n633 B.n44 163.367
R1029 B.n633 B.n46 163.367
R1030 B.n629 B.n46 163.367
R1031 B.n629 B.n51 163.367
R1032 B.n625 B.n51 163.367
R1033 B.n625 B.n53 163.367
R1034 B.n621 B.n53 163.367
R1035 B.n621 B.n58 163.367
R1036 B.n617 B.n58 163.367
R1037 B.n617 B.n60 163.367
R1038 B.n613 B.n60 163.367
R1039 B.n613 B.n65 163.367
R1040 B.n609 B.n65 163.367
R1041 B.n609 B.n67 163.367
R1042 B.n605 B.n67 163.367
R1043 B.n605 B.n72 163.367
R1044 B.n601 B.n72 163.367
R1045 B.n321 B.n320 163.367
R1046 B.n323 B.n321 163.367
R1047 B.n327 B.n316 163.367
R1048 B.n331 B.n329 163.367
R1049 B.n335 B.n314 163.367
R1050 B.n339 B.n337 163.367
R1051 B.n343 B.n312 163.367
R1052 B.n347 B.n345 163.367
R1053 B.n351 B.n310 163.367
R1054 B.n355 B.n353 163.367
R1055 B.n362 B.n308 163.367
R1056 B.n366 B.n364 163.367
R1057 B.n370 B.n306 163.367
R1058 B.n374 B.n372 163.367
R1059 B.n378 B.n304 163.367
R1060 B.n382 B.n380 163.367
R1061 B.n386 B.n299 163.367
R1062 B.n390 B.n388 163.367
R1063 B.n394 B.n297 163.367
R1064 B.n398 B.n396 163.367
R1065 B.n402 B.n295 163.367
R1066 B.n406 B.n404 163.367
R1067 B.n410 B.n293 163.367
R1068 B.n414 B.n412 163.367
R1069 B.n418 B.n291 163.367
R1070 B.n422 B.n420 163.367
R1071 B.n426 B.n283 163.367
R1072 B.n434 B.n283 163.367
R1073 B.n434 B.n281 163.367
R1074 B.n438 B.n281 163.367
R1075 B.n438 B.n275 163.367
R1076 B.n446 B.n275 163.367
R1077 B.n446 B.n273 163.367
R1078 B.n450 B.n273 163.367
R1079 B.n450 B.n267 163.367
R1080 B.n458 B.n267 163.367
R1081 B.n458 B.n265 163.367
R1082 B.n462 B.n265 163.367
R1083 B.n462 B.n258 163.367
R1084 B.n470 B.n258 163.367
R1085 B.n470 B.n256 163.367
R1086 B.n474 B.n256 163.367
R1087 B.n474 B.n251 163.367
R1088 B.n482 B.n251 163.367
R1089 B.n482 B.n249 163.367
R1090 B.n486 B.n249 163.367
R1091 B.n486 B.n243 163.367
R1092 B.n494 B.n243 163.367
R1093 B.n494 B.n241 163.367
R1094 B.n498 B.n241 163.367
R1095 B.n498 B.n235 163.367
R1096 B.n506 B.n235 163.367
R1097 B.n506 B.n233 163.367
R1098 B.n510 B.n233 163.367
R1099 B.n510 B.n227 163.367
R1100 B.n518 B.n227 163.367
R1101 B.n518 B.n225 163.367
R1102 B.n522 B.n225 163.367
R1103 B.n522 B.n218 163.367
R1104 B.n530 B.n218 163.367
R1105 B.n530 B.n216 163.367
R1106 B.n535 B.n216 163.367
R1107 B.n535 B.n211 163.367
R1108 B.n543 B.n211 163.367
R1109 B.n544 B.n543 163.367
R1110 B.n544 B.n5 163.367
R1111 B.n6 B.n5 163.367
R1112 B.n7 B.n6 163.367
R1113 B.n549 B.n7 163.367
R1114 B.n549 B.n12 163.367
R1115 B.n13 B.n12 163.367
R1116 B.n14 B.n13 163.367
R1117 B.n554 B.n14 163.367
R1118 B.n554 B.n19 163.367
R1119 B.n20 B.n19 163.367
R1120 B.n21 B.n20 163.367
R1121 B.n559 B.n21 163.367
R1122 B.n559 B.n26 163.367
R1123 B.n27 B.n26 163.367
R1124 B.n28 B.n27 163.367
R1125 B.n564 B.n28 163.367
R1126 B.n564 B.n33 163.367
R1127 B.n34 B.n33 163.367
R1128 B.n35 B.n34 163.367
R1129 B.n569 B.n35 163.367
R1130 B.n569 B.n40 163.367
R1131 B.n41 B.n40 163.367
R1132 B.n42 B.n41 163.367
R1133 B.n574 B.n42 163.367
R1134 B.n574 B.n47 163.367
R1135 B.n48 B.n47 163.367
R1136 B.n49 B.n48 163.367
R1137 B.n579 B.n49 163.367
R1138 B.n579 B.n54 163.367
R1139 B.n55 B.n54 163.367
R1140 B.n56 B.n55 163.367
R1141 B.n584 B.n56 163.367
R1142 B.n584 B.n61 163.367
R1143 B.n62 B.n61 163.367
R1144 B.n63 B.n62 163.367
R1145 B.n589 B.n63 163.367
R1146 B.n589 B.n68 163.367
R1147 B.n69 B.n68 163.367
R1148 B.n70 B.n69 163.367
R1149 B.n594 B.n70 163.367
R1150 B.n594 B.n75 163.367
R1151 B.n110 B.n109 163.367
R1152 B.n114 B.n113 163.367
R1153 B.n118 B.n117 163.367
R1154 B.n122 B.n121 163.367
R1155 B.n126 B.n125 163.367
R1156 B.n130 B.n129 163.367
R1157 B.n134 B.n133 163.367
R1158 B.n138 B.n137 163.367
R1159 B.n142 B.n141 163.367
R1160 B.n146 B.n145 163.367
R1161 B.n150 B.n149 163.367
R1162 B.n154 B.n153 163.367
R1163 B.n158 B.n157 163.367
R1164 B.n162 B.n161 163.367
R1165 B.n166 B.n165 163.367
R1166 B.n171 B.n170 163.367
R1167 B.n175 B.n174 163.367
R1168 B.n179 B.n178 163.367
R1169 B.n183 B.n182 163.367
R1170 B.n187 B.n186 163.367
R1171 B.n191 B.n190 163.367
R1172 B.n195 B.n194 163.367
R1173 B.n199 B.n198 163.367
R1174 B.n203 B.n202 163.367
R1175 B.n207 B.n206 163.367
R1176 B.n598 B.n102 163.367
R1177 B.n427 B.n288 140.161
R1178 B.n600 B.n599 140.161
R1179 B.n319 B.n287 71.676
R1180 B.n323 B.n322 71.676
R1181 B.n328 B.n327 71.676
R1182 B.n331 B.n330 71.676
R1183 B.n336 B.n335 71.676
R1184 B.n339 B.n338 71.676
R1185 B.n344 B.n343 71.676
R1186 B.n347 B.n346 71.676
R1187 B.n352 B.n351 71.676
R1188 B.n355 B.n354 71.676
R1189 B.n363 B.n362 71.676
R1190 B.n366 B.n365 71.676
R1191 B.n371 B.n370 71.676
R1192 B.n374 B.n373 71.676
R1193 B.n379 B.n378 71.676
R1194 B.n382 B.n381 71.676
R1195 B.n387 B.n386 71.676
R1196 B.n390 B.n389 71.676
R1197 B.n395 B.n394 71.676
R1198 B.n398 B.n397 71.676
R1199 B.n403 B.n402 71.676
R1200 B.n406 B.n405 71.676
R1201 B.n411 B.n410 71.676
R1202 B.n414 B.n413 71.676
R1203 B.n419 B.n418 71.676
R1204 B.n422 B.n421 71.676
R1205 B.n76 B.n74 71.676
R1206 B.n110 B.n77 71.676
R1207 B.n114 B.n78 71.676
R1208 B.n118 B.n79 71.676
R1209 B.n122 B.n80 71.676
R1210 B.n126 B.n81 71.676
R1211 B.n130 B.n82 71.676
R1212 B.n134 B.n83 71.676
R1213 B.n138 B.n84 71.676
R1214 B.n142 B.n85 71.676
R1215 B.n146 B.n86 71.676
R1216 B.n150 B.n87 71.676
R1217 B.n154 B.n88 71.676
R1218 B.n158 B.n89 71.676
R1219 B.n162 B.n90 71.676
R1220 B.n166 B.n91 71.676
R1221 B.n171 B.n92 71.676
R1222 B.n175 B.n93 71.676
R1223 B.n179 B.n94 71.676
R1224 B.n183 B.n95 71.676
R1225 B.n187 B.n96 71.676
R1226 B.n191 B.n97 71.676
R1227 B.n195 B.n98 71.676
R1228 B.n199 B.n99 71.676
R1229 B.n203 B.n100 71.676
R1230 B.n207 B.n101 71.676
R1231 B.n102 B.n101 71.676
R1232 B.n206 B.n100 71.676
R1233 B.n202 B.n99 71.676
R1234 B.n198 B.n98 71.676
R1235 B.n194 B.n97 71.676
R1236 B.n190 B.n96 71.676
R1237 B.n186 B.n95 71.676
R1238 B.n182 B.n94 71.676
R1239 B.n178 B.n93 71.676
R1240 B.n174 B.n92 71.676
R1241 B.n170 B.n91 71.676
R1242 B.n165 B.n90 71.676
R1243 B.n161 B.n89 71.676
R1244 B.n157 B.n88 71.676
R1245 B.n153 B.n87 71.676
R1246 B.n149 B.n86 71.676
R1247 B.n145 B.n85 71.676
R1248 B.n141 B.n84 71.676
R1249 B.n137 B.n83 71.676
R1250 B.n133 B.n82 71.676
R1251 B.n129 B.n81 71.676
R1252 B.n125 B.n80 71.676
R1253 B.n121 B.n79 71.676
R1254 B.n117 B.n78 71.676
R1255 B.n113 B.n77 71.676
R1256 B.n109 B.n76 71.676
R1257 B.n320 B.n319 71.676
R1258 B.n322 B.n316 71.676
R1259 B.n329 B.n328 71.676
R1260 B.n330 B.n314 71.676
R1261 B.n337 B.n336 71.676
R1262 B.n338 B.n312 71.676
R1263 B.n345 B.n344 71.676
R1264 B.n346 B.n310 71.676
R1265 B.n353 B.n352 71.676
R1266 B.n354 B.n308 71.676
R1267 B.n364 B.n363 71.676
R1268 B.n365 B.n306 71.676
R1269 B.n372 B.n371 71.676
R1270 B.n373 B.n304 71.676
R1271 B.n380 B.n379 71.676
R1272 B.n381 B.n299 71.676
R1273 B.n388 B.n387 71.676
R1274 B.n389 B.n297 71.676
R1275 B.n396 B.n395 71.676
R1276 B.n397 B.n295 71.676
R1277 B.n404 B.n403 71.676
R1278 B.n405 B.n293 71.676
R1279 B.n412 B.n411 71.676
R1280 B.n413 B.n291 71.676
R1281 B.n420 B.n419 71.676
R1282 B.n421 B.n289 71.676
R1283 B.n427 B.n284 70.5998
R1284 B.n433 B.n284 70.5998
R1285 B.n433 B.n280 70.5998
R1286 B.n439 B.n280 70.5998
R1287 B.n439 B.n276 70.5998
R1288 B.n445 B.n276 70.5998
R1289 B.n451 B.n272 70.5998
R1290 B.n451 B.n268 70.5998
R1291 B.n457 B.n268 70.5998
R1292 B.n457 B.n264 70.5998
R1293 B.n463 B.n264 70.5998
R1294 B.n463 B.n259 70.5998
R1295 B.n469 B.n259 70.5998
R1296 B.n469 B.n260 70.5998
R1297 B.n475 B.n252 70.5998
R1298 B.n481 B.n252 70.5998
R1299 B.n481 B.n248 70.5998
R1300 B.n487 B.n248 70.5998
R1301 B.n487 B.n244 70.5998
R1302 B.n493 B.n244 70.5998
R1303 B.n499 B.n240 70.5998
R1304 B.n499 B.n236 70.5998
R1305 B.n505 B.n236 70.5998
R1306 B.n505 B.n232 70.5998
R1307 B.n511 B.n232 70.5998
R1308 B.n517 B.n228 70.5998
R1309 B.n517 B.n224 70.5998
R1310 B.n523 B.n224 70.5998
R1311 B.n523 B.n219 70.5998
R1312 B.n529 B.n219 70.5998
R1313 B.n529 B.n220 70.5998
R1314 B.n536 B.n212 70.5998
R1315 B.n542 B.n212 70.5998
R1316 B.n542 B.n4 70.5998
R1317 B.n680 B.n4 70.5998
R1318 B.n680 B.n679 70.5998
R1319 B.n679 B.n678 70.5998
R1320 B.n678 B.n8 70.5998
R1321 B.n672 B.n8 70.5998
R1322 B.n671 B.n670 70.5998
R1323 B.n670 B.n15 70.5998
R1324 B.n664 B.n15 70.5998
R1325 B.n664 B.n663 70.5998
R1326 B.n663 B.n662 70.5998
R1327 B.n662 B.n22 70.5998
R1328 B.n656 B.n655 70.5998
R1329 B.n655 B.n654 70.5998
R1330 B.n654 B.n29 70.5998
R1331 B.n648 B.n29 70.5998
R1332 B.n648 B.n647 70.5998
R1333 B.n646 B.n36 70.5998
R1334 B.n640 B.n36 70.5998
R1335 B.n640 B.n639 70.5998
R1336 B.n639 B.n638 70.5998
R1337 B.n638 B.n43 70.5998
R1338 B.n632 B.n43 70.5998
R1339 B.n631 B.n630 70.5998
R1340 B.n630 B.n50 70.5998
R1341 B.n624 B.n50 70.5998
R1342 B.n624 B.n623 70.5998
R1343 B.n623 B.n622 70.5998
R1344 B.n622 B.n57 70.5998
R1345 B.n616 B.n57 70.5998
R1346 B.n616 B.n615 70.5998
R1347 B.n614 B.n64 70.5998
R1348 B.n608 B.n64 70.5998
R1349 B.n608 B.n607 70.5998
R1350 B.n607 B.n606 70.5998
R1351 B.n606 B.n71 70.5998
R1352 B.n600 B.n71 70.5998
R1353 B.n260 B.t3 67.4852
R1354 B.t0 B.n631 67.4852
R1355 B.n302 B.n301 59.5399
R1356 B.n360 B.n359 59.5399
R1357 B.n107 B.n106 59.5399
R1358 B.n168 B.n104 59.5399
R1359 B.n536 B.t6 57.1029
R1360 B.n672 B.t4 57.1029
R1361 B.n511 B.t1 55.0265
R1362 B.n656 B.t7 55.0265
R1363 B.t9 B.n272 46.7207
R1364 B.n615 B.t13 46.7207
R1365 B.t5 B.n240 44.6442
R1366 B.n647 B.t2 44.6442
R1367 B.n301 B.n300 42.2793
R1368 B.n359 B.n358 42.2793
R1369 B.n106 B.n105 42.2793
R1370 B.n104 B.n103 42.2793
R1371 B.n602 B.n73 36.9956
R1372 B.n597 B.n596 36.9956
R1373 B.n425 B.n424 36.9956
R1374 B.n429 B.n286 36.9956
R1375 B.n493 B.t5 25.9561
R1376 B.t2 B.n646 25.9561
R1377 B.n445 B.t9 23.8797
R1378 B.t13 B.n614 23.8797
R1379 B B.n682 18.0485
R1380 B.t1 B.n228 15.5739
R1381 B.t7 B.n22 15.5739
R1382 B.n220 B.t6 13.4974
R1383 B.t4 B.n671 13.4974
R1384 B.n108 B.n73 10.6151
R1385 B.n111 B.n108 10.6151
R1386 B.n112 B.n111 10.6151
R1387 B.n115 B.n112 10.6151
R1388 B.n116 B.n115 10.6151
R1389 B.n119 B.n116 10.6151
R1390 B.n120 B.n119 10.6151
R1391 B.n123 B.n120 10.6151
R1392 B.n124 B.n123 10.6151
R1393 B.n127 B.n124 10.6151
R1394 B.n128 B.n127 10.6151
R1395 B.n131 B.n128 10.6151
R1396 B.n132 B.n131 10.6151
R1397 B.n135 B.n132 10.6151
R1398 B.n136 B.n135 10.6151
R1399 B.n139 B.n136 10.6151
R1400 B.n140 B.n139 10.6151
R1401 B.n143 B.n140 10.6151
R1402 B.n144 B.n143 10.6151
R1403 B.n147 B.n144 10.6151
R1404 B.n148 B.n147 10.6151
R1405 B.n152 B.n151 10.6151
R1406 B.n155 B.n152 10.6151
R1407 B.n156 B.n155 10.6151
R1408 B.n159 B.n156 10.6151
R1409 B.n160 B.n159 10.6151
R1410 B.n163 B.n160 10.6151
R1411 B.n164 B.n163 10.6151
R1412 B.n167 B.n164 10.6151
R1413 B.n172 B.n169 10.6151
R1414 B.n173 B.n172 10.6151
R1415 B.n176 B.n173 10.6151
R1416 B.n177 B.n176 10.6151
R1417 B.n180 B.n177 10.6151
R1418 B.n181 B.n180 10.6151
R1419 B.n184 B.n181 10.6151
R1420 B.n185 B.n184 10.6151
R1421 B.n188 B.n185 10.6151
R1422 B.n189 B.n188 10.6151
R1423 B.n192 B.n189 10.6151
R1424 B.n193 B.n192 10.6151
R1425 B.n196 B.n193 10.6151
R1426 B.n197 B.n196 10.6151
R1427 B.n200 B.n197 10.6151
R1428 B.n201 B.n200 10.6151
R1429 B.n204 B.n201 10.6151
R1430 B.n205 B.n204 10.6151
R1431 B.n208 B.n205 10.6151
R1432 B.n209 B.n208 10.6151
R1433 B.n597 B.n209 10.6151
R1434 B.n425 B.n282 10.6151
R1435 B.n435 B.n282 10.6151
R1436 B.n436 B.n435 10.6151
R1437 B.n437 B.n436 10.6151
R1438 B.n437 B.n274 10.6151
R1439 B.n447 B.n274 10.6151
R1440 B.n448 B.n447 10.6151
R1441 B.n449 B.n448 10.6151
R1442 B.n449 B.n266 10.6151
R1443 B.n459 B.n266 10.6151
R1444 B.n460 B.n459 10.6151
R1445 B.n461 B.n460 10.6151
R1446 B.n461 B.n257 10.6151
R1447 B.n471 B.n257 10.6151
R1448 B.n472 B.n471 10.6151
R1449 B.n473 B.n472 10.6151
R1450 B.n473 B.n250 10.6151
R1451 B.n483 B.n250 10.6151
R1452 B.n484 B.n483 10.6151
R1453 B.n485 B.n484 10.6151
R1454 B.n485 B.n242 10.6151
R1455 B.n495 B.n242 10.6151
R1456 B.n496 B.n495 10.6151
R1457 B.n497 B.n496 10.6151
R1458 B.n497 B.n234 10.6151
R1459 B.n507 B.n234 10.6151
R1460 B.n508 B.n507 10.6151
R1461 B.n509 B.n508 10.6151
R1462 B.n509 B.n226 10.6151
R1463 B.n519 B.n226 10.6151
R1464 B.n520 B.n519 10.6151
R1465 B.n521 B.n520 10.6151
R1466 B.n521 B.n217 10.6151
R1467 B.n531 B.n217 10.6151
R1468 B.n532 B.n531 10.6151
R1469 B.n534 B.n532 10.6151
R1470 B.n534 B.n533 10.6151
R1471 B.n533 B.n210 10.6151
R1472 B.n545 B.n210 10.6151
R1473 B.n546 B.n545 10.6151
R1474 B.n547 B.n546 10.6151
R1475 B.n548 B.n547 10.6151
R1476 B.n550 B.n548 10.6151
R1477 B.n551 B.n550 10.6151
R1478 B.n552 B.n551 10.6151
R1479 B.n553 B.n552 10.6151
R1480 B.n555 B.n553 10.6151
R1481 B.n556 B.n555 10.6151
R1482 B.n557 B.n556 10.6151
R1483 B.n558 B.n557 10.6151
R1484 B.n560 B.n558 10.6151
R1485 B.n561 B.n560 10.6151
R1486 B.n562 B.n561 10.6151
R1487 B.n563 B.n562 10.6151
R1488 B.n565 B.n563 10.6151
R1489 B.n566 B.n565 10.6151
R1490 B.n567 B.n566 10.6151
R1491 B.n568 B.n567 10.6151
R1492 B.n570 B.n568 10.6151
R1493 B.n571 B.n570 10.6151
R1494 B.n572 B.n571 10.6151
R1495 B.n573 B.n572 10.6151
R1496 B.n575 B.n573 10.6151
R1497 B.n576 B.n575 10.6151
R1498 B.n577 B.n576 10.6151
R1499 B.n578 B.n577 10.6151
R1500 B.n580 B.n578 10.6151
R1501 B.n581 B.n580 10.6151
R1502 B.n582 B.n581 10.6151
R1503 B.n583 B.n582 10.6151
R1504 B.n585 B.n583 10.6151
R1505 B.n586 B.n585 10.6151
R1506 B.n587 B.n586 10.6151
R1507 B.n588 B.n587 10.6151
R1508 B.n590 B.n588 10.6151
R1509 B.n591 B.n590 10.6151
R1510 B.n592 B.n591 10.6151
R1511 B.n593 B.n592 10.6151
R1512 B.n595 B.n593 10.6151
R1513 B.n596 B.n595 10.6151
R1514 B.n318 B.n286 10.6151
R1515 B.n318 B.n317 10.6151
R1516 B.n324 B.n317 10.6151
R1517 B.n325 B.n324 10.6151
R1518 B.n326 B.n325 10.6151
R1519 B.n326 B.n315 10.6151
R1520 B.n332 B.n315 10.6151
R1521 B.n333 B.n332 10.6151
R1522 B.n334 B.n333 10.6151
R1523 B.n334 B.n313 10.6151
R1524 B.n340 B.n313 10.6151
R1525 B.n341 B.n340 10.6151
R1526 B.n342 B.n341 10.6151
R1527 B.n342 B.n311 10.6151
R1528 B.n348 B.n311 10.6151
R1529 B.n349 B.n348 10.6151
R1530 B.n350 B.n349 10.6151
R1531 B.n350 B.n309 10.6151
R1532 B.n356 B.n309 10.6151
R1533 B.n357 B.n356 10.6151
R1534 B.n361 B.n357 10.6151
R1535 B.n367 B.n307 10.6151
R1536 B.n368 B.n367 10.6151
R1537 B.n369 B.n368 10.6151
R1538 B.n369 B.n305 10.6151
R1539 B.n375 B.n305 10.6151
R1540 B.n376 B.n375 10.6151
R1541 B.n377 B.n376 10.6151
R1542 B.n377 B.n303 10.6151
R1543 B.n384 B.n383 10.6151
R1544 B.n385 B.n384 10.6151
R1545 B.n385 B.n298 10.6151
R1546 B.n391 B.n298 10.6151
R1547 B.n392 B.n391 10.6151
R1548 B.n393 B.n392 10.6151
R1549 B.n393 B.n296 10.6151
R1550 B.n399 B.n296 10.6151
R1551 B.n400 B.n399 10.6151
R1552 B.n401 B.n400 10.6151
R1553 B.n401 B.n294 10.6151
R1554 B.n407 B.n294 10.6151
R1555 B.n408 B.n407 10.6151
R1556 B.n409 B.n408 10.6151
R1557 B.n409 B.n292 10.6151
R1558 B.n415 B.n292 10.6151
R1559 B.n416 B.n415 10.6151
R1560 B.n417 B.n416 10.6151
R1561 B.n417 B.n290 10.6151
R1562 B.n423 B.n290 10.6151
R1563 B.n424 B.n423 10.6151
R1564 B.n430 B.n429 10.6151
R1565 B.n431 B.n430 10.6151
R1566 B.n431 B.n278 10.6151
R1567 B.n441 B.n278 10.6151
R1568 B.n442 B.n441 10.6151
R1569 B.n443 B.n442 10.6151
R1570 B.n443 B.n270 10.6151
R1571 B.n453 B.n270 10.6151
R1572 B.n454 B.n453 10.6151
R1573 B.n455 B.n454 10.6151
R1574 B.n455 B.n262 10.6151
R1575 B.n465 B.n262 10.6151
R1576 B.n466 B.n465 10.6151
R1577 B.n467 B.n466 10.6151
R1578 B.n467 B.n254 10.6151
R1579 B.n477 B.n254 10.6151
R1580 B.n478 B.n477 10.6151
R1581 B.n479 B.n478 10.6151
R1582 B.n479 B.n246 10.6151
R1583 B.n489 B.n246 10.6151
R1584 B.n490 B.n489 10.6151
R1585 B.n491 B.n490 10.6151
R1586 B.n491 B.n238 10.6151
R1587 B.n501 B.n238 10.6151
R1588 B.n502 B.n501 10.6151
R1589 B.n503 B.n502 10.6151
R1590 B.n503 B.n230 10.6151
R1591 B.n513 B.n230 10.6151
R1592 B.n514 B.n513 10.6151
R1593 B.n515 B.n514 10.6151
R1594 B.n515 B.n222 10.6151
R1595 B.n525 B.n222 10.6151
R1596 B.n526 B.n525 10.6151
R1597 B.n527 B.n526 10.6151
R1598 B.n527 B.n214 10.6151
R1599 B.n538 B.n214 10.6151
R1600 B.n539 B.n538 10.6151
R1601 B.n540 B.n539 10.6151
R1602 B.n540 B.n0 10.6151
R1603 B.n676 B.n1 10.6151
R1604 B.n676 B.n675 10.6151
R1605 B.n675 B.n674 10.6151
R1606 B.n674 B.n10 10.6151
R1607 B.n668 B.n10 10.6151
R1608 B.n668 B.n667 10.6151
R1609 B.n667 B.n666 10.6151
R1610 B.n666 B.n17 10.6151
R1611 B.n660 B.n17 10.6151
R1612 B.n660 B.n659 10.6151
R1613 B.n659 B.n658 10.6151
R1614 B.n658 B.n24 10.6151
R1615 B.n652 B.n24 10.6151
R1616 B.n652 B.n651 10.6151
R1617 B.n651 B.n650 10.6151
R1618 B.n650 B.n31 10.6151
R1619 B.n644 B.n31 10.6151
R1620 B.n644 B.n643 10.6151
R1621 B.n643 B.n642 10.6151
R1622 B.n642 B.n38 10.6151
R1623 B.n636 B.n38 10.6151
R1624 B.n636 B.n635 10.6151
R1625 B.n635 B.n634 10.6151
R1626 B.n634 B.n45 10.6151
R1627 B.n628 B.n45 10.6151
R1628 B.n628 B.n627 10.6151
R1629 B.n627 B.n626 10.6151
R1630 B.n626 B.n52 10.6151
R1631 B.n620 B.n52 10.6151
R1632 B.n620 B.n619 10.6151
R1633 B.n619 B.n618 10.6151
R1634 B.n618 B.n59 10.6151
R1635 B.n612 B.n59 10.6151
R1636 B.n612 B.n611 10.6151
R1637 B.n611 B.n610 10.6151
R1638 B.n610 B.n66 10.6151
R1639 B.n604 B.n66 10.6151
R1640 B.n604 B.n603 10.6151
R1641 B.n603 B.n602 10.6151
R1642 B.n151 B.n107 6.5566
R1643 B.n168 B.n167 6.5566
R1644 B.n360 B.n307 6.5566
R1645 B.n303 B.n302 6.5566
R1646 B.n148 B.n107 4.05904
R1647 B.n169 B.n168 4.05904
R1648 B.n361 B.n360 4.05904
R1649 B.n383 B.n302 4.05904
R1650 B.n475 B.t3 3.11518
R1651 B.n632 B.t0 3.11518
R1652 B.n682 B.n0 2.81026
R1653 B.n682 B.n1 2.81026
R1654 VN.n22 VN.n21 184.909
R1655 VN.n45 VN.n44 184.909
R1656 VN.n43 VN.n23 161.3
R1657 VN.n42 VN.n41 161.3
R1658 VN.n40 VN.n24 161.3
R1659 VN.n39 VN.n38 161.3
R1660 VN.n37 VN.n25 161.3
R1661 VN.n35 VN.n34 161.3
R1662 VN.n33 VN.n26 161.3
R1663 VN.n32 VN.n31 161.3
R1664 VN.n30 VN.n27 161.3
R1665 VN.n20 VN.n0 161.3
R1666 VN.n19 VN.n18 161.3
R1667 VN.n17 VN.n1 161.3
R1668 VN.n16 VN.n15 161.3
R1669 VN.n14 VN.n2 161.3
R1670 VN.n12 VN.n11 161.3
R1671 VN.n10 VN.n3 161.3
R1672 VN.n9 VN.n8 161.3
R1673 VN.n7 VN.n4 161.3
R1674 VN.n5 VN.t3 101.775
R1675 VN.n28 VN.t5 101.775
R1676 VN.n6 VN.t4 69.3043
R1677 VN.n13 VN.t2 69.3043
R1678 VN.n21 VN.t7 69.3043
R1679 VN.n29 VN.t6 69.3043
R1680 VN.n36 VN.t0 69.3043
R1681 VN.n44 VN.t1 69.3043
R1682 VN.n8 VN.n3 56.5617
R1683 VN.n31 VN.n26 56.5617
R1684 VN.n6 VN.n5 53.2962
R1685 VN.n29 VN.n28 53.2962
R1686 VN.n15 VN.n1 47.3584
R1687 VN.n38 VN.n24 47.3584
R1688 VN VN.n45 42.5781
R1689 VN.n19 VN.n1 33.7956
R1690 VN.n42 VN.n24 33.7956
R1691 VN.n8 VN.n7 24.5923
R1692 VN.n12 VN.n3 24.5923
R1693 VN.n15 VN.n14 24.5923
R1694 VN.n20 VN.n19 24.5923
R1695 VN.n31 VN.n30 24.5923
R1696 VN.n38 VN.n37 24.5923
R1697 VN.n35 VN.n26 24.5923
R1698 VN.n43 VN.n42 24.5923
R1699 VN.n7 VN.n6 16.7229
R1700 VN.n13 VN.n12 16.7229
R1701 VN.n30 VN.n29 16.7229
R1702 VN.n36 VN.n35 16.7229
R1703 VN.n28 VN.n27 12.4908
R1704 VN.n5 VN.n4 12.4908
R1705 VN.n14 VN.n13 7.86989
R1706 VN.n37 VN.n36 7.86989
R1707 VN.n21 VN.n20 0.984173
R1708 VN.n44 VN.n43 0.984173
R1709 VN.n45 VN.n23 0.189894
R1710 VN.n41 VN.n23 0.189894
R1711 VN.n41 VN.n40 0.189894
R1712 VN.n40 VN.n39 0.189894
R1713 VN.n39 VN.n25 0.189894
R1714 VN.n34 VN.n25 0.189894
R1715 VN.n34 VN.n33 0.189894
R1716 VN.n33 VN.n32 0.189894
R1717 VN.n32 VN.n27 0.189894
R1718 VN.n9 VN.n4 0.189894
R1719 VN.n10 VN.n9 0.189894
R1720 VN.n11 VN.n10 0.189894
R1721 VN.n11 VN.n2 0.189894
R1722 VN.n16 VN.n2 0.189894
R1723 VN.n17 VN.n16 0.189894
R1724 VN.n18 VN.n17 0.189894
R1725 VN.n18 VN.n0 0.189894
R1726 VN.n22 VN.n0 0.189894
R1727 VN VN.n22 0.0516364
R1728 VDD2.n2 VDD2.n1 70.3152
R1729 VDD2.n2 VDD2.n0 70.3152
R1730 VDD2 VDD2.n5 70.3123
R1731 VDD2.n4 VDD2.n3 69.431
R1732 VDD2.n4 VDD2.n2 36.7584
R1733 VDD2.n5 VDD2.t1 3.7223
R1734 VDD2.n5 VDD2.t2 3.7223
R1735 VDD2.n3 VDD2.t6 3.7223
R1736 VDD2.n3 VDD2.t7 3.7223
R1737 VDD2.n1 VDD2.t5 3.7223
R1738 VDD2.n1 VDD2.t0 3.7223
R1739 VDD2.n0 VDD2.t4 3.7223
R1740 VDD2.n0 VDD2.t3 3.7223
R1741 VDD2 VDD2.n4 0.998345
C0 VDD2 VTAIL 5.49294f
C1 VP VN 5.50376f
C2 VTAIL VDD1 5.44355f
C3 VTAIL VN 4.37265f
C4 VP VTAIL 4.38676f
C5 VDD2 VDD1 1.38526f
C6 VDD2 VN 3.81006f
C7 VDD2 VP 0.443945f
C8 VN VDD1 0.150432f
C9 VP VDD1 4.09845f
C10 VDD2 B 4.093289f
C11 VDD1 B 4.455714f
C12 VTAIL B 5.714921f
C13 VN B 11.95164f
C14 VP B 10.527409f
C15 VDD2.t4 B 0.103121f
C16 VDD2.t3 B 0.103121f
C17 VDD2.n0 B 0.852398f
C18 VDD2.t5 B 0.103121f
C19 VDD2.t0 B 0.103121f
C20 VDD2.n1 B 0.852398f
C21 VDD2.n2 B 2.38057f
C22 VDD2.t6 B 0.103121f
C23 VDD2.t7 B 0.103121f
C24 VDD2.n3 B 0.84705f
C25 VDD2.n4 B 2.12237f
C26 VDD2.t1 B 0.103121f
C27 VDD2.t2 B 0.103121f
C28 VDD2.n5 B 0.85237f
C29 VN.n0 B 0.030196f
C30 VN.t7 B 0.780668f
C31 VN.n1 B 0.026328f
C32 VN.n2 B 0.030196f
C33 VN.t2 B 0.780668f
C34 VN.n3 B 0.043894f
C35 VN.n4 B 0.222352f
C36 VN.t4 B 0.780668f
C37 VN.t3 B 0.924113f
C38 VN.n5 B 0.371986f
C39 VN.n6 B 0.378255f
C40 VN.n7 B 0.047149f
C41 VN.n8 B 0.043894f
C42 VN.n9 B 0.030196f
C43 VN.n10 B 0.030196f
C44 VN.n11 B 0.030196f
C45 VN.n12 B 0.047149f
C46 VN.n13 B 0.30526f
C47 VN.n14 B 0.037197f
C48 VN.n15 B 0.056792f
C49 VN.n16 B 0.030196f
C50 VN.n17 B 0.030196f
C51 VN.n18 B 0.030196f
C52 VN.n19 B 0.060662f
C53 VN.n20 B 0.029457f
C54 VN.n21 B 0.37195f
C55 VN.n22 B 0.033161f
C56 VN.n23 B 0.030196f
C57 VN.t1 B 0.780668f
C58 VN.n24 B 0.026328f
C59 VN.n25 B 0.030196f
C60 VN.t0 B 0.780668f
C61 VN.n26 B 0.043894f
C62 VN.n27 B 0.222352f
C63 VN.t6 B 0.780668f
C64 VN.t5 B 0.924113f
C65 VN.n28 B 0.371986f
C66 VN.n29 B 0.378255f
C67 VN.n30 B 0.047149f
C68 VN.n31 B 0.043894f
C69 VN.n32 B 0.030196f
C70 VN.n33 B 0.030196f
C71 VN.n34 B 0.030196f
C72 VN.n35 B 0.047149f
C73 VN.n36 B 0.30526f
C74 VN.n37 B 0.037197f
C75 VN.n38 B 0.056792f
C76 VN.n39 B 0.030196f
C77 VN.n40 B 0.030196f
C78 VN.n41 B 0.030196f
C79 VN.n42 B 0.060662f
C80 VN.n43 B 0.029457f
C81 VN.n44 B 0.37195f
C82 VN.n45 B 1.28569f
C83 VTAIL.t7 B 0.096277f
C84 VTAIL.t2 B 0.096277f
C85 VTAIL.n0 B 0.734181f
C86 VTAIL.n1 B 0.35203f
C87 VTAIL.n2 B 0.03219f
C88 VTAIL.n3 B 0.022901f
C89 VTAIL.n4 B 0.012306f
C90 VTAIL.n5 B 0.029087f
C91 VTAIL.n6 B 0.01303f
C92 VTAIL.n7 B 0.022901f
C93 VTAIL.n8 B 0.012306f
C94 VTAIL.n9 B 0.021815f
C95 VTAIL.n10 B 0.017178f
C96 VTAIL.t4 B 0.047511f
C97 VTAIL.n11 B 0.094398f
C98 VTAIL.n12 B 0.473087f
C99 VTAIL.n13 B 0.012306f
C100 VTAIL.n14 B 0.01303f
C101 VTAIL.n15 B 0.029087f
C102 VTAIL.n16 B 0.029087f
C103 VTAIL.n17 B 0.01303f
C104 VTAIL.n18 B 0.012306f
C105 VTAIL.n19 B 0.022901f
C106 VTAIL.n20 B 0.022901f
C107 VTAIL.n21 B 0.012306f
C108 VTAIL.n22 B 0.01303f
C109 VTAIL.n23 B 0.029087f
C110 VTAIL.n24 B 0.062969f
C111 VTAIL.n25 B 0.01303f
C112 VTAIL.n26 B 0.012306f
C113 VTAIL.n27 B 0.054186f
C114 VTAIL.n28 B 0.035272f
C115 VTAIL.n29 B 0.193615f
C116 VTAIL.n30 B 0.03219f
C117 VTAIL.n31 B 0.022901f
C118 VTAIL.n32 B 0.012306f
C119 VTAIL.n33 B 0.029087f
C120 VTAIL.n34 B 0.01303f
C121 VTAIL.n35 B 0.022901f
C122 VTAIL.n36 B 0.012306f
C123 VTAIL.n37 B 0.021815f
C124 VTAIL.n38 B 0.017178f
C125 VTAIL.t11 B 0.047511f
C126 VTAIL.n39 B 0.094398f
C127 VTAIL.n40 B 0.473087f
C128 VTAIL.n41 B 0.012306f
C129 VTAIL.n42 B 0.01303f
C130 VTAIL.n43 B 0.029087f
C131 VTAIL.n44 B 0.029087f
C132 VTAIL.n45 B 0.01303f
C133 VTAIL.n46 B 0.012306f
C134 VTAIL.n47 B 0.022901f
C135 VTAIL.n48 B 0.022901f
C136 VTAIL.n49 B 0.012306f
C137 VTAIL.n50 B 0.01303f
C138 VTAIL.n51 B 0.029087f
C139 VTAIL.n52 B 0.062969f
C140 VTAIL.n53 B 0.01303f
C141 VTAIL.n54 B 0.012306f
C142 VTAIL.n55 B 0.054186f
C143 VTAIL.n56 B 0.035272f
C144 VTAIL.n57 B 0.193615f
C145 VTAIL.t8 B 0.096277f
C146 VTAIL.t9 B 0.096277f
C147 VTAIL.n58 B 0.734181f
C148 VTAIL.n59 B 0.486416f
C149 VTAIL.n60 B 0.03219f
C150 VTAIL.n61 B 0.022901f
C151 VTAIL.n62 B 0.012306f
C152 VTAIL.n63 B 0.029087f
C153 VTAIL.n64 B 0.01303f
C154 VTAIL.n65 B 0.022901f
C155 VTAIL.n66 B 0.012306f
C156 VTAIL.n67 B 0.021815f
C157 VTAIL.n68 B 0.017178f
C158 VTAIL.t10 B 0.047511f
C159 VTAIL.n69 B 0.094398f
C160 VTAIL.n70 B 0.473087f
C161 VTAIL.n71 B 0.012306f
C162 VTAIL.n72 B 0.01303f
C163 VTAIL.n73 B 0.029087f
C164 VTAIL.n74 B 0.029087f
C165 VTAIL.n75 B 0.01303f
C166 VTAIL.n76 B 0.012306f
C167 VTAIL.n77 B 0.022901f
C168 VTAIL.n78 B 0.022901f
C169 VTAIL.n79 B 0.012306f
C170 VTAIL.n80 B 0.01303f
C171 VTAIL.n81 B 0.029087f
C172 VTAIL.n82 B 0.062969f
C173 VTAIL.n83 B 0.01303f
C174 VTAIL.n84 B 0.012306f
C175 VTAIL.n85 B 0.054186f
C176 VTAIL.n86 B 0.035272f
C177 VTAIL.n87 B 0.94714f
C178 VTAIL.n88 B 0.03219f
C179 VTAIL.n89 B 0.022901f
C180 VTAIL.n90 B 0.012306f
C181 VTAIL.n91 B 0.029087f
C182 VTAIL.n92 B 0.01303f
C183 VTAIL.n93 B 0.022901f
C184 VTAIL.n94 B 0.012306f
C185 VTAIL.n95 B 0.021815f
C186 VTAIL.n96 B 0.017178f
C187 VTAIL.t3 B 0.047511f
C188 VTAIL.n97 B 0.094398f
C189 VTAIL.n98 B 0.473087f
C190 VTAIL.n99 B 0.012306f
C191 VTAIL.n100 B 0.01303f
C192 VTAIL.n101 B 0.029087f
C193 VTAIL.n102 B 0.029087f
C194 VTAIL.n103 B 0.01303f
C195 VTAIL.n104 B 0.012306f
C196 VTAIL.n105 B 0.022901f
C197 VTAIL.n106 B 0.022901f
C198 VTAIL.n107 B 0.012306f
C199 VTAIL.n108 B 0.01303f
C200 VTAIL.n109 B 0.029087f
C201 VTAIL.n110 B 0.062969f
C202 VTAIL.n111 B 0.01303f
C203 VTAIL.n112 B 0.012306f
C204 VTAIL.n113 B 0.054186f
C205 VTAIL.n114 B 0.035272f
C206 VTAIL.n115 B 0.94714f
C207 VTAIL.t5 B 0.096277f
C208 VTAIL.t1 B 0.096277f
C209 VTAIL.n116 B 0.734186f
C210 VTAIL.n117 B 0.486411f
C211 VTAIL.n118 B 0.03219f
C212 VTAIL.n119 B 0.022901f
C213 VTAIL.n120 B 0.012306f
C214 VTAIL.n121 B 0.029087f
C215 VTAIL.n122 B 0.01303f
C216 VTAIL.n123 B 0.022901f
C217 VTAIL.n124 B 0.012306f
C218 VTAIL.n125 B 0.021815f
C219 VTAIL.n126 B 0.017178f
C220 VTAIL.t6 B 0.047511f
C221 VTAIL.n127 B 0.094398f
C222 VTAIL.n128 B 0.473087f
C223 VTAIL.n129 B 0.012306f
C224 VTAIL.n130 B 0.01303f
C225 VTAIL.n131 B 0.029087f
C226 VTAIL.n132 B 0.029087f
C227 VTAIL.n133 B 0.01303f
C228 VTAIL.n134 B 0.012306f
C229 VTAIL.n135 B 0.022901f
C230 VTAIL.n136 B 0.022901f
C231 VTAIL.n137 B 0.012306f
C232 VTAIL.n138 B 0.01303f
C233 VTAIL.n139 B 0.029087f
C234 VTAIL.n140 B 0.062969f
C235 VTAIL.n141 B 0.01303f
C236 VTAIL.n142 B 0.012306f
C237 VTAIL.n143 B 0.054186f
C238 VTAIL.n144 B 0.035272f
C239 VTAIL.n145 B 0.193615f
C240 VTAIL.n146 B 0.03219f
C241 VTAIL.n147 B 0.022901f
C242 VTAIL.n148 B 0.012306f
C243 VTAIL.n149 B 0.029087f
C244 VTAIL.n150 B 0.01303f
C245 VTAIL.n151 B 0.022901f
C246 VTAIL.n152 B 0.012306f
C247 VTAIL.n153 B 0.021815f
C248 VTAIL.n154 B 0.017178f
C249 VTAIL.t15 B 0.047511f
C250 VTAIL.n155 B 0.094398f
C251 VTAIL.n156 B 0.473087f
C252 VTAIL.n157 B 0.012306f
C253 VTAIL.n158 B 0.01303f
C254 VTAIL.n159 B 0.029087f
C255 VTAIL.n160 B 0.029087f
C256 VTAIL.n161 B 0.01303f
C257 VTAIL.n162 B 0.012306f
C258 VTAIL.n163 B 0.022901f
C259 VTAIL.n164 B 0.022901f
C260 VTAIL.n165 B 0.012306f
C261 VTAIL.n166 B 0.01303f
C262 VTAIL.n167 B 0.029087f
C263 VTAIL.n168 B 0.062969f
C264 VTAIL.n169 B 0.01303f
C265 VTAIL.n170 B 0.012306f
C266 VTAIL.n171 B 0.054186f
C267 VTAIL.n172 B 0.035272f
C268 VTAIL.n173 B 0.193615f
C269 VTAIL.t13 B 0.096277f
C270 VTAIL.t14 B 0.096277f
C271 VTAIL.n174 B 0.734186f
C272 VTAIL.n175 B 0.486411f
C273 VTAIL.n176 B 0.03219f
C274 VTAIL.n177 B 0.022901f
C275 VTAIL.n178 B 0.012306f
C276 VTAIL.n179 B 0.029087f
C277 VTAIL.n180 B 0.01303f
C278 VTAIL.n181 B 0.022901f
C279 VTAIL.n182 B 0.012306f
C280 VTAIL.n183 B 0.021815f
C281 VTAIL.n184 B 0.017178f
C282 VTAIL.t12 B 0.047511f
C283 VTAIL.n185 B 0.094398f
C284 VTAIL.n186 B 0.473087f
C285 VTAIL.n187 B 0.012306f
C286 VTAIL.n188 B 0.01303f
C287 VTAIL.n189 B 0.029087f
C288 VTAIL.n190 B 0.029087f
C289 VTAIL.n191 B 0.01303f
C290 VTAIL.n192 B 0.012306f
C291 VTAIL.n193 B 0.022901f
C292 VTAIL.n194 B 0.022901f
C293 VTAIL.n195 B 0.012306f
C294 VTAIL.n196 B 0.01303f
C295 VTAIL.n197 B 0.029087f
C296 VTAIL.n198 B 0.062969f
C297 VTAIL.n199 B 0.01303f
C298 VTAIL.n200 B 0.012306f
C299 VTAIL.n201 B 0.054186f
C300 VTAIL.n202 B 0.035272f
C301 VTAIL.n203 B 0.94714f
C302 VTAIL.n204 B 0.03219f
C303 VTAIL.n205 B 0.022901f
C304 VTAIL.n206 B 0.012306f
C305 VTAIL.n207 B 0.029087f
C306 VTAIL.n208 B 0.01303f
C307 VTAIL.n209 B 0.022901f
C308 VTAIL.n210 B 0.012306f
C309 VTAIL.n211 B 0.021815f
C310 VTAIL.n212 B 0.017178f
C311 VTAIL.t0 B 0.047511f
C312 VTAIL.n213 B 0.094398f
C313 VTAIL.n214 B 0.473087f
C314 VTAIL.n215 B 0.012306f
C315 VTAIL.n216 B 0.01303f
C316 VTAIL.n217 B 0.029087f
C317 VTAIL.n218 B 0.029087f
C318 VTAIL.n219 B 0.01303f
C319 VTAIL.n220 B 0.012306f
C320 VTAIL.n221 B 0.022901f
C321 VTAIL.n222 B 0.022901f
C322 VTAIL.n223 B 0.012306f
C323 VTAIL.n224 B 0.01303f
C324 VTAIL.n225 B 0.029087f
C325 VTAIL.n226 B 0.062969f
C326 VTAIL.n227 B 0.01303f
C327 VTAIL.n228 B 0.012306f
C328 VTAIL.n229 B 0.054186f
C329 VTAIL.n230 B 0.035272f
C330 VTAIL.n231 B 0.942846f
C331 VDD1.t2 B 0.104322f
C332 VDD1.t4 B 0.104322f
C333 VDD1.n0 B 0.863137f
C334 VDD1.t7 B 0.104322f
C335 VDD1.t6 B 0.104322f
C336 VDD1.n1 B 0.862328f
C337 VDD1.t0 B 0.104322f
C338 VDD1.t3 B 0.104322f
C339 VDD1.n2 B 0.862328f
C340 VDD1.n3 B 2.46065f
C341 VDD1.t5 B 0.104322f
C342 VDD1.t1 B 0.104322f
C343 VDD1.n4 B 0.856914f
C344 VDD1.n5 B 2.1771f
C345 VP.n0 B 0.030953f
C346 VP.t4 B 0.800242f
C347 VP.n1 B 0.026988f
C348 VP.n2 B 0.030953f
C349 VP.t6 B 0.800242f
C350 VP.n3 B 0.044994f
C351 VP.n4 B 0.030953f
C352 VP.t7 B 0.800242f
C353 VP.n5 B 0.058216f
C354 VP.n6 B 0.030953f
C355 VP.t5 B 0.800242f
C356 VP.n7 B 0.381277f
C357 VP.n8 B 0.030953f
C358 VP.t3 B 0.800242f
C359 VP.n9 B 0.026988f
C360 VP.n10 B 0.030953f
C361 VP.t1 B 0.800242f
C362 VP.n11 B 0.044994f
C363 VP.n12 B 0.227928f
C364 VP.t2 B 0.800242f
C365 VP.t0 B 0.947284f
C366 VP.n13 B 0.381313f
C367 VP.n14 B 0.387739f
C368 VP.n15 B 0.048331f
C369 VP.n16 B 0.044994f
C370 VP.n17 B 0.030953f
C371 VP.n18 B 0.030953f
C372 VP.n19 B 0.030953f
C373 VP.n20 B 0.048331f
C374 VP.n21 B 0.312914f
C375 VP.n22 B 0.03813f
C376 VP.n23 B 0.058216f
C377 VP.n24 B 0.030953f
C378 VP.n25 B 0.030953f
C379 VP.n26 B 0.030953f
C380 VP.n27 B 0.062183f
C381 VP.n28 B 0.030196f
C382 VP.n29 B 0.381277f
C383 VP.n30 B 1.29761f
C384 VP.n31 B 1.32405f
C385 VP.n32 B 0.030953f
C386 VP.n33 B 0.030196f
C387 VP.n34 B 0.062183f
C388 VP.n35 B 0.026988f
C389 VP.n36 B 0.030953f
C390 VP.n37 B 0.030953f
C391 VP.n38 B 0.030953f
C392 VP.n39 B 0.03813f
C393 VP.n40 B 0.312914f
C394 VP.n41 B 0.048331f
C395 VP.n42 B 0.044994f
C396 VP.n43 B 0.030953f
C397 VP.n44 B 0.030953f
C398 VP.n45 B 0.030953f
C399 VP.n46 B 0.048331f
C400 VP.n47 B 0.312914f
C401 VP.n48 B 0.03813f
C402 VP.n49 B 0.058216f
C403 VP.n50 B 0.030953f
C404 VP.n51 B 0.030953f
C405 VP.n52 B 0.030953f
C406 VP.n53 B 0.062183f
C407 VP.n54 B 0.030196f
C408 VP.n55 B 0.381277f
C409 VP.n56 B 0.033993f
.ends

