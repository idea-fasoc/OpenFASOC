* NGSPICE file created from diff_pair_sample_0155.ext - technology: sky130A

.subckt diff_pair_sample_0155 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=0 ps=0 w=8.39 l=0.2
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=3.2721 ps=17.56 w=8.39 l=0.2
X2 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=3.2721 ps=17.56 w=8.39 l=0.2
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=0 ps=0 w=8.39 l=0.2
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=0 ps=0 w=8.39 l=0.2
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=0 ps=0 w=8.39 l=0.2
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=3.2721 ps=17.56 w=8.39 l=0.2
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2721 pd=17.56 as=3.2721 ps=17.56 w=8.39 l=0.2
R0 B.n265 B.t6 1247.34
R1 B.n262 B.t10 1247.34
R2 B.n64 B.t2 1247.34
R3 B.n62 B.t13 1247.34
R4 B.n458 B.n457 585
R5 B.n204 B.n60 585
R6 B.n203 B.n202 585
R7 B.n201 B.n200 585
R8 B.n199 B.n198 585
R9 B.n197 B.n196 585
R10 B.n195 B.n194 585
R11 B.n193 B.n192 585
R12 B.n191 B.n190 585
R13 B.n189 B.n188 585
R14 B.n187 B.n186 585
R15 B.n185 B.n184 585
R16 B.n183 B.n182 585
R17 B.n181 B.n180 585
R18 B.n179 B.n178 585
R19 B.n177 B.n176 585
R20 B.n175 B.n174 585
R21 B.n173 B.n172 585
R22 B.n171 B.n170 585
R23 B.n169 B.n168 585
R24 B.n167 B.n166 585
R25 B.n165 B.n164 585
R26 B.n163 B.n162 585
R27 B.n161 B.n160 585
R28 B.n159 B.n158 585
R29 B.n157 B.n156 585
R30 B.n155 B.n154 585
R31 B.n153 B.n152 585
R32 B.n151 B.n150 585
R33 B.n149 B.n148 585
R34 B.n147 B.n146 585
R35 B.n144 B.n143 585
R36 B.n142 B.n141 585
R37 B.n140 B.n139 585
R38 B.n138 B.n137 585
R39 B.n136 B.n135 585
R40 B.n134 B.n133 585
R41 B.n132 B.n131 585
R42 B.n130 B.n129 585
R43 B.n128 B.n127 585
R44 B.n126 B.n125 585
R45 B.n123 B.n122 585
R46 B.n121 B.n120 585
R47 B.n119 B.n118 585
R48 B.n117 B.n116 585
R49 B.n115 B.n114 585
R50 B.n113 B.n112 585
R51 B.n111 B.n110 585
R52 B.n109 B.n108 585
R53 B.n107 B.n106 585
R54 B.n105 B.n104 585
R55 B.n103 B.n102 585
R56 B.n101 B.n100 585
R57 B.n99 B.n98 585
R58 B.n97 B.n96 585
R59 B.n95 B.n94 585
R60 B.n93 B.n92 585
R61 B.n91 B.n90 585
R62 B.n89 B.n88 585
R63 B.n87 B.n86 585
R64 B.n85 B.n84 585
R65 B.n83 B.n82 585
R66 B.n81 B.n80 585
R67 B.n79 B.n78 585
R68 B.n77 B.n76 585
R69 B.n75 B.n74 585
R70 B.n73 B.n72 585
R71 B.n71 B.n70 585
R72 B.n69 B.n68 585
R73 B.n67 B.n66 585
R74 B.n25 B.n24 585
R75 B.n463 B.n462 585
R76 B.n456 B.n61 585
R77 B.n61 B.n22 585
R78 B.n455 B.n21 585
R79 B.n467 B.n21 585
R80 B.n454 B.n20 585
R81 B.n468 B.n20 585
R82 B.n453 B.n19 585
R83 B.n469 B.n19 585
R84 B.n452 B.n451 585
R85 B.n451 B.n15 585
R86 B.n450 B.n14 585
R87 B.n475 B.n14 585
R88 B.n449 B.n13 585
R89 B.n476 B.n13 585
R90 B.n448 B.n12 585
R91 B.n477 B.n12 585
R92 B.n447 B.n446 585
R93 B.n446 B.n11 585
R94 B.n445 B.n7 585
R95 B.n483 B.n7 585
R96 B.n444 B.n6 585
R97 B.n484 B.n6 585
R98 B.n443 B.n5 585
R99 B.n485 B.n5 585
R100 B.n442 B.n441 585
R101 B.n441 B.n4 585
R102 B.n440 B.n205 585
R103 B.n440 B.n439 585
R104 B.n429 B.n206 585
R105 B.n432 B.n206 585
R106 B.n431 B.n430 585
R107 B.n433 B.n431 585
R108 B.n428 B.n211 585
R109 B.n211 B.n210 585
R110 B.n427 B.n426 585
R111 B.n426 B.n425 585
R112 B.n213 B.n212 585
R113 B.n214 B.n213 585
R114 B.n418 B.n417 585
R115 B.n419 B.n418 585
R116 B.n416 B.n219 585
R117 B.n219 B.n218 585
R118 B.n415 B.n414 585
R119 B.n414 B.n413 585
R120 B.n221 B.n220 585
R121 B.n222 B.n221 585
R122 B.n409 B.n408 585
R123 B.n225 B.n224 585
R124 B.n405 B.n404 585
R125 B.n406 B.n405 585
R126 B.n403 B.n261 585
R127 B.n402 B.n401 585
R128 B.n400 B.n399 585
R129 B.n398 B.n397 585
R130 B.n396 B.n395 585
R131 B.n394 B.n393 585
R132 B.n392 B.n391 585
R133 B.n390 B.n389 585
R134 B.n388 B.n387 585
R135 B.n386 B.n385 585
R136 B.n384 B.n383 585
R137 B.n382 B.n381 585
R138 B.n380 B.n379 585
R139 B.n378 B.n377 585
R140 B.n376 B.n375 585
R141 B.n374 B.n373 585
R142 B.n372 B.n371 585
R143 B.n370 B.n369 585
R144 B.n368 B.n367 585
R145 B.n366 B.n365 585
R146 B.n364 B.n363 585
R147 B.n362 B.n361 585
R148 B.n360 B.n359 585
R149 B.n358 B.n357 585
R150 B.n356 B.n355 585
R151 B.n354 B.n353 585
R152 B.n352 B.n351 585
R153 B.n350 B.n349 585
R154 B.n348 B.n347 585
R155 B.n346 B.n345 585
R156 B.n344 B.n343 585
R157 B.n342 B.n341 585
R158 B.n340 B.n339 585
R159 B.n338 B.n337 585
R160 B.n336 B.n335 585
R161 B.n334 B.n333 585
R162 B.n332 B.n331 585
R163 B.n330 B.n329 585
R164 B.n328 B.n327 585
R165 B.n326 B.n325 585
R166 B.n324 B.n323 585
R167 B.n322 B.n321 585
R168 B.n320 B.n319 585
R169 B.n318 B.n317 585
R170 B.n316 B.n315 585
R171 B.n314 B.n313 585
R172 B.n312 B.n311 585
R173 B.n310 B.n309 585
R174 B.n308 B.n307 585
R175 B.n306 B.n305 585
R176 B.n304 B.n303 585
R177 B.n302 B.n301 585
R178 B.n300 B.n299 585
R179 B.n298 B.n297 585
R180 B.n296 B.n295 585
R181 B.n294 B.n293 585
R182 B.n292 B.n291 585
R183 B.n290 B.n289 585
R184 B.n288 B.n287 585
R185 B.n286 B.n285 585
R186 B.n284 B.n283 585
R187 B.n282 B.n281 585
R188 B.n280 B.n279 585
R189 B.n278 B.n277 585
R190 B.n276 B.n275 585
R191 B.n274 B.n273 585
R192 B.n272 B.n271 585
R193 B.n270 B.n269 585
R194 B.n268 B.n260 585
R195 B.n406 B.n260 585
R196 B.n410 B.n223 585
R197 B.n223 B.n222 585
R198 B.n412 B.n411 585
R199 B.n413 B.n412 585
R200 B.n217 B.n216 585
R201 B.n218 B.n217 585
R202 B.n421 B.n420 585
R203 B.n420 B.n419 585
R204 B.n422 B.n215 585
R205 B.n215 B.n214 585
R206 B.n424 B.n423 585
R207 B.n425 B.n424 585
R208 B.n209 B.n208 585
R209 B.n210 B.n209 585
R210 B.n435 B.n434 585
R211 B.n434 B.n433 585
R212 B.n436 B.n207 585
R213 B.n432 B.n207 585
R214 B.n438 B.n437 585
R215 B.n439 B.n438 585
R216 B.n2 B.n0 585
R217 B.n4 B.n2 585
R218 B.n3 B.n1 585
R219 B.n484 B.n3 585
R220 B.n482 B.n481 585
R221 B.n483 B.n482 585
R222 B.n480 B.n8 585
R223 B.n11 B.n8 585
R224 B.n479 B.n478 585
R225 B.n478 B.n477 585
R226 B.n10 B.n9 585
R227 B.n476 B.n10 585
R228 B.n474 B.n473 585
R229 B.n475 B.n474 585
R230 B.n472 B.n16 585
R231 B.n16 B.n15 585
R232 B.n471 B.n470 585
R233 B.n470 B.n469 585
R234 B.n18 B.n17 585
R235 B.n468 B.n18 585
R236 B.n466 B.n465 585
R237 B.n467 B.n466 585
R238 B.n464 B.n23 585
R239 B.n23 B.n22 585
R240 B.n487 B.n486 585
R241 B.n486 B.n485 585
R242 B.n408 B.n223 511.721
R243 B.n462 B.n23 511.721
R244 B.n260 B.n221 511.721
R245 B.n458 B.n61 511.721
R246 B.n460 B.n459 256.663
R247 B.n460 B.n59 256.663
R248 B.n460 B.n58 256.663
R249 B.n460 B.n57 256.663
R250 B.n460 B.n56 256.663
R251 B.n460 B.n55 256.663
R252 B.n460 B.n54 256.663
R253 B.n460 B.n53 256.663
R254 B.n460 B.n52 256.663
R255 B.n460 B.n51 256.663
R256 B.n460 B.n50 256.663
R257 B.n460 B.n49 256.663
R258 B.n460 B.n48 256.663
R259 B.n460 B.n47 256.663
R260 B.n460 B.n46 256.663
R261 B.n460 B.n45 256.663
R262 B.n460 B.n44 256.663
R263 B.n460 B.n43 256.663
R264 B.n460 B.n42 256.663
R265 B.n460 B.n41 256.663
R266 B.n460 B.n40 256.663
R267 B.n460 B.n39 256.663
R268 B.n460 B.n38 256.663
R269 B.n460 B.n37 256.663
R270 B.n460 B.n36 256.663
R271 B.n460 B.n35 256.663
R272 B.n460 B.n34 256.663
R273 B.n460 B.n33 256.663
R274 B.n460 B.n32 256.663
R275 B.n460 B.n31 256.663
R276 B.n460 B.n30 256.663
R277 B.n460 B.n29 256.663
R278 B.n460 B.n28 256.663
R279 B.n460 B.n27 256.663
R280 B.n460 B.n26 256.663
R281 B.n461 B.n460 256.663
R282 B.n407 B.n406 256.663
R283 B.n406 B.n226 256.663
R284 B.n406 B.n227 256.663
R285 B.n406 B.n228 256.663
R286 B.n406 B.n229 256.663
R287 B.n406 B.n230 256.663
R288 B.n406 B.n231 256.663
R289 B.n406 B.n232 256.663
R290 B.n406 B.n233 256.663
R291 B.n406 B.n234 256.663
R292 B.n406 B.n235 256.663
R293 B.n406 B.n236 256.663
R294 B.n406 B.n237 256.663
R295 B.n406 B.n238 256.663
R296 B.n406 B.n239 256.663
R297 B.n406 B.n240 256.663
R298 B.n406 B.n241 256.663
R299 B.n406 B.n242 256.663
R300 B.n406 B.n243 256.663
R301 B.n406 B.n244 256.663
R302 B.n406 B.n245 256.663
R303 B.n406 B.n246 256.663
R304 B.n406 B.n247 256.663
R305 B.n406 B.n248 256.663
R306 B.n406 B.n249 256.663
R307 B.n406 B.n250 256.663
R308 B.n406 B.n251 256.663
R309 B.n406 B.n252 256.663
R310 B.n406 B.n253 256.663
R311 B.n406 B.n254 256.663
R312 B.n406 B.n255 256.663
R313 B.n406 B.n256 256.663
R314 B.n406 B.n257 256.663
R315 B.n406 B.n258 256.663
R316 B.n406 B.n259 256.663
R317 B.n412 B.n223 163.367
R318 B.n412 B.n217 163.367
R319 B.n420 B.n217 163.367
R320 B.n420 B.n215 163.367
R321 B.n424 B.n215 163.367
R322 B.n424 B.n209 163.367
R323 B.n434 B.n209 163.367
R324 B.n434 B.n207 163.367
R325 B.n438 B.n207 163.367
R326 B.n438 B.n2 163.367
R327 B.n486 B.n2 163.367
R328 B.n486 B.n3 163.367
R329 B.n482 B.n3 163.367
R330 B.n482 B.n8 163.367
R331 B.n478 B.n8 163.367
R332 B.n478 B.n10 163.367
R333 B.n474 B.n10 163.367
R334 B.n474 B.n16 163.367
R335 B.n470 B.n16 163.367
R336 B.n470 B.n18 163.367
R337 B.n466 B.n18 163.367
R338 B.n466 B.n23 163.367
R339 B.n405 B.n225 163.367
R340 B.n405 B.n261 163.367
R341 B.n401 B.n400 163.367
R342 B.n397 B.n396 163.367
R343 B.n393 B.n392 163.367
R344 B.n389 B.n388 163.367
R345 B.n385 B.n384 163.367
R346 B.n381 B.n380 163.367
R347 B.n377 B.n376 163.367
R348 B.n373 B.n372 163.367
R349 B.n369 B.n368 163.367
R350 B.n365 B.n364 163.367
R351 B.n361 B.n360 163.367
R352 B.n357 B.n356 163.367
R353 B.n353 B.n352 163.367
R354 B.n349 B.n348 163.367
R355 B.n345 B.n344 163.367
R356 B.n341 B.n340 163.367
R357 B.n337 B.n336 163.367
R358 B.n333 B.n332 163.367
R359 B.n329 B.n328 163.367
R360 B.n325 B.n324 163.367
R361 B.n321 B.n320 163.367
R362 B.n317 B.n316 163.367
R363 B.n313 B.n312 163.367
R364 B.n309 B.n308 163.367
R365 B.n305 B.n304 163.367
R366 B.n301 B.n300 163.367
R367 B.n297 B.n296 163.367
R368 B.n293 B.n292 163.367
R369 B.n289 B.n288 163.367
R370 B.n285 B.n284 163.367
R371 B.n281 B.n280 163.367
R372 B.n277 B.n276 163.367
R373 B.n273 B.n272 163.367
R374 B.n269 B.n260 163.367
R375 B.n414 B.n221 163.367
R376 B.n414 B.n219 163.367
R377 B.n418 B.n219 163.367
R378 B.n418 B.n213 163.367
R379 B.n426 B.n213 163.367
R380 B.n426 B.n211 163.367
R381 B.n431 B.n211 163.367
R382 B.n431 B.n206 163.367
R383 B.n440 B.n206 163.367
R384 B.n441 B.n440 163.367
R385 B.n441 B.n5 163.367
R386 B.n6 B.n5 163.367
R387 B.n7 B.n6 163.367
R388 B.n446 B.n7 163.367
R389 B.n446 B.n12 163.367
R390 B.n13 B.n12 163.367
R391 B.n14 B.n13 163.367
R392 B.n451 B.n14 163.367
R393 B.n451 B.n19 163.367
R394 B.n20 B.n19 163.367
R395 B.n21 B.n20 163.367
R396 B.n61 B.n21 163.367
R397 B.n66 B.n25 163.367
R398 B.n70 B.n69 163.367
R399 B.n74 B.n73 163.367
R400 B.n78 B.n77 163.367
R401 B.n82 B.n81 163.367
R402 B.n86 B.n85 163.367
R403 B.n90 B.n89 163.367
R404 B.n94 B.n93 163.367
R405 B.n98 B.n97 163.367
R406 B.n102 B.n101 163.367
R407 B.n106 B.n105 163.367
R408 B.n110 B.n109 163.367
R409 B.n114 B.n113 163.367
R410 B.n118 B.n117 163.367
R411 B.n122 B.n121 163.367
R412 B.n127 B.n126 163.367
R413 B.n131 B.n130 163.367
R414 B.n135 B.n134 163.367
R415 B.n139 B.n138 163.367
R416 B.n143 B.n142 163.367
R417 B.n148 B.n147 163.367
R418 B.n152 B.n151 163.367
R419 B.n156 B.n155 163.367
R420 B.n160 B.n159 163.367
R421 B.n164 B.n163 163.367
R422 B.n168 B.n167 163.367
R423 B.n172 B.n171 163.367
R424 B.n176 B.n175 163.367
R425 B.n180 B.n179 163.367
R426 B.n184 B.n183 163.367
R427 B.n188 B.n187 163.367
R428 B.n192 B.n191 163.367
R429 B.n196 B.n195 163.367
R430 B.n200 B.n199 163.367
R431 B.n202 B.n60 163.367
R432 B.n406 B.n222 111.728
R433 B.n460 B.n22 111.728
R434 B.n265 B.t9 83.2342
R435 B.n62 B.t14 83.2342
R436 B.n262 B.t12 83.2245
R437 B.n64 B.t4 83.2245
R438 B.n266 B.t8 72.9554
R439 B.n63 B.t15 72.9554
R440 B.n263 B.t11 72.9457
R441 B.n65 B.t5 72.9457
R442 B.n408 B.n407 71.676
R443 B.n261 B.n226 71.676
R444 B.n400 B.n227 71.676
R445 B.n396 B.n228 71.676
R446 B.n392 B.n229 71.676
R447 B.n388 B.n230 71.676
R448 B.n384 B.n231 71.676
R449 B.n380 B.n232 71.676
R450 B.n376 B.n233 71.676
R451 B.n372 B.n234 71.676
R452 B.n368 B.n235 71.676
R453 B.n364 B.n236 71.676
R454 B.n360 B.n237 71.676
R455 B.n356 B.n238 71.676
R456 B.n352 B.n239 71.676
R457 B.n348 B.n240 71.676
R458 B.n344 B.n241 71.676
R459 B.n340 B.n242 71.676
R460 B.n336 B.n243 71.676
R461 B.n332 B.n244 71.676
R462 B.n328 B.n245 71.676
R463 B.n324 B.n246 71.676
R464 B.n320 B.n247 71.676
R465 B.n316 B.n248 71.676
R466 B.n312 B.n249 71.676
R467 B.n308 B.n250 71.676
R468 B.n304 B.n251 71.676
R469 B.n300 B.n252 71.676
R470 B.n296 B.n253 71.676
R471 B.n292 B.n254 71.676
R472 B.n288 B.n255 71.676
R473 B.n284 B.n256 71.676
R474 B.n280 B.n257 71.676
R475 B.n276 B.n258 71.676
R476 B.n272 B.n259 71.676
R477 B.n462 B.n461 71.676
R478 B.n66 B.n26 71.676
R479 B.n70 B.n27 71.676
R480 B.n74 B.n28 71.676
R481 B.n78 B.n29 71.676
R482 B.n82 B.n30 71.676
R483 B.n86 B.n31 71.676
R484 B.n90 B.n32 71.676
R485 B.n94 B.n33 71.676
R486 B.n98 B.n34 71.676
R487 B.n102 B.n35 71.676
R488 B.n106 B.n36 71.676
R489 B.n110 B.n37 71.676
R490 B.n114 B.n38 71.676
R491 B.n118 B.n39 71.676
R492 B.n122 B.n40 71.676
R493 B.n127 B.n41 71.676
R494 B.n131 B.n42 71.676
R495 B.n135 B.n43 71.676
R496 B.n139 B.n44 71.676
R497 B.n143 B.n45 71.676
R498 B.n148 B.n46 71.676
R499 B.n152 B.n47 71.676
R500 B.n156 B.n48 71.676
R501 B.n160 B.n49 71.676
R502 B.n164 B.n50 71.676
R503 B.n168 B.n51 71.676
R504 B.n172 B.n52 71.676
R505 B.n176 B.n53 71.676
R506 B.n180 B.n54 71.676
R507 B.n184 B.n55 71.676
R508 B.n188 B.n56 71.676
R509 B.n192 B.n57 71.676
R510 B.n196 B.n58 71.676
R511 B.n200 B.n59 71.676
R512 B.n459 B.n60 71.676
R513 B.n459 B.n458 71.676
R514 B.n202 B.n59 71.676
R515 B.n199 B.n58 71.676
R516 B.n195 B.n57 71.676
R517 B.n191 B.n56 71.676
R518 B.n187 B.n55 71.676
R519 B.n183 B.n54 71.676
R520 B.n179 B.n53 71.676
R521 B.n175 B.n52 71.676
R522 B.n171 B.n51 71.676
R523 B.n167 B.n50 71.676
R524 B.n163 B.n49 71.676
R525 B.n159 B.n48 71.676
R526 B.n155 B.n47 71.676
R527 B.n151 B.n46 71.676
R528 B.n147 B.n45 71.676
R529 B.n142 B.n44 71.676
R530 B.n138 B.n43 71.676
R531 B.n134 B.n42 71.676
R532 B.n130 B.n41 71.676
R533 B.n126 B.n40 71.676
R534 B.n121 B.n39 71.676
R535 B.n117 B.n38 71.676
R536 B.n113 B.n37 71.676
R537 B.n109 B.n36 71.676
R538 B.n105 B.n35 71.676
R539 B.n101 B.n34 71.676
R540 B.n97 B.n33 71.676
R541 B.n93 B.n32 71.676
R542 B.n89 B.n31 71.676
R543 B.n85 B.n30 71.676
R544 B.n81 B.n29 71.676
R545 B.n77 B.n28 71.676
R546 B.n73 B.n27 71.676
R547 B.n69 B.n26 71.676
R548 B.n461 B.n25 71.676
R549 B.n407 B.n225 71.676
R550 B.n401 B.n226 71.676
R551 B.n397 B.n227 71.676
R552 B.n393 B.n228 71.676
R553 B.n389 B.n229 71.676
R554 B.n385 B.n230 71.676
R555 B.n381 B.n231 71.676
R556 B.n377 B.n232 71.676
R557 B.n373 B.n233 71.676
R558 B.n369 B.n234 71.676
R559 B.n365 B.n235 71.676
R560 B.n361 B.n236 71.676
R561 B.n357 B.n237 71.676
R562 B.n353 B.n238 71.676
R563 B.n349 B.n239 71.676
R564 B.n345 B.n240 71.676
R565 B.n341 B.n241 71.676
R566 B.n337 B.n242 71.676
R567 B.n333 B.n243 71.676
R568 B.n329 B.n244 71.676
R569 B.n325 B.n245 71.676
R570 B.n321 B.n246 71.676
R571 B.n317 B.n247 71.676
R572 B.n313 B.n248 71.676
R573 B.n309 B.n249 71.676
R574 B.n305 B.n250 71.676
R575 B.n301 B.n251 71.676
R576 B.n297 B.n252 71.676
R577 B.n293 B.n253 71.676
R578 B.n289 B.n254 71.676
R579 B.n285 B.n255 71.676
R580 B.n281 B.n256 71.676
R581 B.n277 B.n257 71.676
R582 B.n273 B.n258 71.676
R583 B.n269 B.n259 71.676
R584 B.n267 B.n266 59.5399
R585 B.n264 B.n263 59.5399
R586 B.n124 B.n65 59.5399
R587 B.n145 B.n63 59.5399
R588 B.n413 B.n222 54.6589
R589 B.n413 B.n218 54.6589
R590 B.n419 B.n218 54.6589
R591 B.n425 B.n214 54.6589
R592 B.n425 B.n210 54.6589
R593 B.n433 B.n210 54.6589
R594 B.n433 B.n432 54.6589
R595 B.n439 B.n4 54.6589
R596 B.n485 B.n4 54.6589
R597 B.n485 B.n484 54.6589
R598 B.n484 B.n483 54.6589
R599 B.n477 B.n11 54.6589
R600 B.n477 B.n476 54.6589
R601 B.n476 B.n475 54.6589
R602 B.n475 B.n15 54.6589
R603 B.n469 B.n468 54.6589
R604 B.n468 B.n467 54.6589
R605 B.n467 B.n22 54.6589
R606 B.n419 B.t7 46.6209
R607 B.n469 B.t3 46.6209
R608 B.n432 B.t1 33.7601
R609 B.n11 B.t0 33.7601
R610 B.n464 B.n463 33.2493
R611 B.n457 B.n456 33.2493
R612 B.n268 B.n220 33.2493
R613 B.n410 B.n409 33.2493
R614 B.n439 B.t1 20.8993
R615 B.n483 B.t0 20.8993
R616 B B.n487 18.0485
R617 B.n463 B.n24 10.6151
R618 B.n67 B.n24 10.6151
R619 B.n68 B.n67 10.6151
R620 B.n71 B.n68 10.6151
R621 B.n72 B.n71 10.6151
R622 B.n75 B.n72 10.6151
R623 B.n76 B.n75 10.6151
R624 B.n79 B.n76 10.6151
R625 B.n80 B.n79 10.6151
R626 B.n83 B.n80 10.6151
R627 B.n84 B.n83 10.6151
R628 B.n87 B.n84 10.6151
R629 B.n88 B.n87 10.6151
R630 B.n91 B.n88 10.6151
R631 B.n92 B.n91 10.6151
R632 B.n95 B.n92 10.6151
R633 B.n96 B.n95 10.6151
R634 B.n99 B.n96 10.6151
R635 B.n100 B.n99 10.6151
R636 B.n103 B.n100 10.6151
R637 B.n104 B.n103 10.6151
R638 B.n107 B.n104 10.6151
R639 B.n108 B.n107 10.6151
R640 B.n111 B.n108 10.6151
R641 B.n112 B.n111 10.6151
R642 B.n115 B.n112 10.6151
R643 B.n116 B.n115 10.6151
R644 B.n119 B.n116 10.6151
R645 B.n120 B.n119 10.6151
R646 B.n123 B.n120 10.6151
R647 B.n128 B.n125 10.6151
R648 B.n129 B.n128 10.6151
R649 B.n132 B.n129 10.6151
R650 B.n133 B.n132 10.6151
R651 B.n136 B.n133 10.6151
R652 B.n137 B.n136 10.6151
R653 B.n140 B.n137 10.6151
R654 B.n141 B.n140 10.6151
R655 B.n144 B.n141 10.6151
R656 B.n149 B.n146 10.6151
R657 B.n150 B.n149 10.6151
R658 B.n153 B.n150 10.6151
R659 B.n154 B.n153 10.6151
R660 B.n157 B.n154 10.6151
R661 B.n158 B.n157 10.6151
R662 B.n161 B.n158 10.6151
R663 B.n162 B.n161 10.6151
R664 B.n165 B.n162 10.6151
R665 B.n166 B.n165 10.6151
R666 B.n169 B.n166 10.6151
R667 B.n170 B.n169 10.6151
R668 B.n173 B.n170 10.6151
R669 B.n174 B.n173 10.6151
R670 B.n177 B.n174 10.6151
R671 B.n178 B.n177 10.6151
R672 B.n181 B.n178 10.6151
R673 B.n182 B.n181 10.6151
R674 B.n185 B.n182 10.6151
R675 B.n186 B.n185 10.6151
R676 B.n189 B.n186 10.6151
R677 B.n190 B.n189 10.6151
R678 B.n193 B.n190 10.6151
R679 B.n194 B.n193 10.6151
R680 B.n197 B.n194 10.6151
R681 B.n198 B.n197 10.6151
R682 B.n201 B.n198 10.6151
R683 B.n203 B.n201 10.6151
R684 B.n204 B.n203 10.6151
R685 B.n457 B.n204 10.6151
R686 B.n415 B.n220 10.6151
R687 B.n416 B.n415 10.6151
R688 B.n417 B.n416 10.6151
R689 B.n417 B.n212 10.6151
R690 B.n427 B.n212 10.6151
R691 B.n428 B.n427 10.6151
R692 B.n430 B.n428 10.6151
R693 B.n430 B.n429 10.6151
R694 B.n429 B.n205 10.6151
R695 B.n442 B.n205 10.6151
R696 B.n443 B.n442 10.6151
R697 B.n444 B.n443 10.6151
R698 B.n445 B.n444 10.6151
R699 B.n447 B.n445 10.6151
R700 B.n448 B.n447 10.6151
R701 B.n449 B.n448 10.6151
R702 B.n450 B.n449 10.6151
R703 B.n452 B.n450 10.6151
R704 B.n453 B.n452 10.6151
R705 B.n454 B.n453 10.6151
R706 B.n455 B.n454 10.6151
R707 B.n456 B.n455 10.6151
R708 B.n409 B.n224 10.6151
R709 B.n404 B.n224 10.6151
R710 B.n404 B.n403 10.6151
R711 B.n403 B.n402 10.6151
R712 B.n402 B.n399 10.6151
R713 B.n399 B.n398 10.6151
R714 B.n398 B.n395 10.6151
R715 B.n395 B.n394 10.6151
R716 B.n394 B.n391 10.6151
R717 B.n391 B.n390 10.6151
R718 B.n390 B.n387 10.6151
R719 B.n387 B.n386 10.6151
R720 B.n386 B.n383 10.6151
R721 B.n383 B.n382 10.6151
R722 B.n382 B.n379 10.6151
R723 B.n379 B.n378 10.6151
R724 B.n378 B.n375 10.6151
R725 B.n375 B.n374 10.6151
R726 B.n374 B.n371 10.6151
R727 B.n371 B.n370 10.6151
R728 B.n370 B.n367 10.6151
R729 B.n367 B.n366 10.6151
R730 B.n366 B.n363 10.6151
R731 B.n363 B.n362 10.6151
R732 B.n362 B.n359 10.6151
R733 B.n359 B.n358 10.6151
R734 B.n358 B.n355 10.6151
R735 B.n355 B.n354 10.6151
R736 B.n354 B.n351 10.6151
R737 B.n351 B.n350 10.6151
R738 B.n347 B.n346 10.6151
R739 B.n346 B.n343 10.6151
R740 B.n343 B.n342 10.6151
R741 B.n342 B.n339 10.6151
R742 B.n339 B.n338 10.6151
R743 B.n338 B.n335 10.6151
R744 B.n335 B.n334 10.6151
R745 B.n334 B.n331 10.6151
R746 B.n331 B.n330 10.6151
R747 B.n327 B.n326 10.6151
R748 B.n326 B.n323 10.6151
R749 B.n323 B.n322 10.6151
R750 B.n322 B.n319 10.6151
R751 B.n319 B.n318 10.6151
R752 B.n318 B.n315 10.6151
R753 B.n315 B.n314 10.6151
R754 B.n314 B.n311 10.6151
R755 B.n311 B.n310 10.6151
R756 B.n310 B.n307 10.6151
R757 B.n307 B.n306 10.6151
R758 B.n306 B.n303 10.6151
R759 B.n303 B.n302 10.6151
R760 B.n302 B.n299 10.6151
R761 B.n299 B.n298 10.6151
R762 B.n298 B.n295 10.6151
R763 B.n295 B.n294 10.6151
R764 B.n294 B.n291 10.6151
R765 B.n291 B.n290 10.6151
R766 B.n290 B.n287 10.6151
R767 B.n287 B.n286 10.6151
R768 B.n286 B.n283 10.6151
R769 B.n283 B.n282 10.6151
R770 B.n282 B.n279 10.6151
R771 B.n279 B.n278 10.6151
R772 B.n278 B.n275 10.6151
R773 B.n275 B.n274 10.6151
R774 B.n274 B.n271 10.6151
R775 B.n271 B.n270 10.6151
R776 B.n270 B.n268 10.6151
R777 B.n411 B.n410 10.6151
R778 B.n411 B.n216 10.6151
R779 B.n421 B.n216 10.6151
R780 B.n422 B.n421 10.6151
R781 B.n423 B.n422 10.6151
R782 B.n423 B.n208 10.6151
R783 B.n435 B.n208 10.6151
R784 B.n436 B.n435 10.6151
R785 B.n437 B.n436 10.6151
R786 B.n437 B.n0 10.6151
R787 B.n481 B.n1 10.6151
R788 B.n481 B.n480 10.6151
R789 B.n480 B.n479 10.6151
R790 B.n479 B.n9 10.6151
R791 B.n473 B.n9 10.6151
R792 B.n473 B.n472 10.6151
R793 B.n472 B.n471 10.6151
R794 B.n471 B.n17 10.6151
R795 B.n465 B.n17 10.6151
R796 B.n465 B.n464 10.6151
R797 B.n266 B.n265 10.2793
R798 B.n263 B.n262 10.2793
R799 B.n65 B.n64 10.2793
R800 B.n63 B.n62 10.2793
R801 B.n124 B.n123 8.74196
R802 B.n146 B.n145 8.74196
R803 B.n350 B.n264 8.74196
R804 B.n327 B.n267 8.74196
R805 B.t7 B.n214 8.0385
R806 B.t3 B.n15 8.0385
R807 B.n487 B.n0 2.81026
R808 B.n487 B.n1 2.81026
R809 B.n125 B.n124 1.87367
R810 B.n145 B.n144 1.87367
R811 B.n347 B.n264 1.87367
R812 B.n330 B.n267 1.87367
R813 VN VN.t0 1390.2
R814 VN VN.t1 1354.3
R815 VTAIL.n1 VTAIL.t2 53.8374
R816 VTAIL.n3 VTAIL.t3 53.8373
R817 VTAIL.n0 VTAIL.t0 53.8373
R818 VTAIL.n2 VTAIL.t1 53.8373
R819 VTAIL.n1 VTAIL.n0 20.5307
R820 VTAIL.n3 VTAIL.n2 20.0738
R821 VTAIL.n2 VTAIL.n1 0.698776
R822 VTAIL VTAIL.n0 0.642741
R823 VTAIL VTAIL.n3 0.0565345
R824 VDD2.n0 VDD2.t0 102.34
R825 VDD2.n0 VDD2.t1 70.5161
R826 VDD2 VDD2.n0 0.172914
R827 VP.n0 VP.t1 1389.82
R828 VP.n0 VP.t0 1354.25
R829 VP VP.n0 0.0516364
R830 VDD1 VDD1.t1 102.978
R831 VDD1 VDD1.t0 70.6885
C0 VN VP 3.67463f
C1 VDD1 VN 0.148341f
C2 VTAIL VN 0.521014f
C3 VDD1 VP 1.03133f
C4 VDD2 VN 0.949738f
C5 VTAIL VP 0.535611f
C6 VDD1 VTAIL 5.72914f
C7 VDD2 VP 0.233606f
C8 VDD1 VDD2 0.420123f
C9 VTAIL VDD2 5.75994f
C10 VDD2 B 2.906509f
C11 VDD1 B 5.28416f
C12 VTAIL B 4.38042f
C13 VN B 6.483951f
C14 VP B 3.222192f
C15 VDD1.t0 B 1.53066f
C16 VDD1.t1 B 1.87815f
C17 VP.t1 B 0.285941f
C18 VP.t0 B 0.245509f
C19 VP.n0 B 3.16272f
C20 VDD2.t0 B 1.91716f
C21 VDD2.t1 B 1.57823f
C22 VDD2.n0 B 2.27627f
C23 VTAIL.t0 B 1.63476f
C24 VTAIL.n0 B 1.25315f
C25 VTAIL.t2 B 1.63477f
C26 VTAIL.n1 B 1.25733f
C27 VTAIL.t1 B 1.63476f
C28 VTAIL.n2 B 1.22314f
C29 VTAIL.t3 B 1.63476f
C30 VTAIL.n3 B 1.17507f
C31 VN.t1 B 0.241072f
C32 VN.t0 B 0.281999f
.ends

