* NGSPICE file created from diff_pair_sample_0582.ext - technology: sky130A

.subckt diff_pair_sample_0582 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=0 ps=0 w=12.49 l=1.12
X1 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=0 ps=0 w=12.49 l=1.12
X2 VDD1.t7 VP.t0 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=4.8711 ps=25.76 w=12.49 l=1.12
X3 VTAIL.t15 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=2.06085 ps=12.82 w=12.49 l=1.12
X4 VDD2.t7 VN.t0 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=4.8711 ps=25.76 w=12.49 l=1.12
X5 VTAIL.t4 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X6 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X7 VTAIL.t6 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=2.06085 ps=12.82 w=12.49 l=1.12
X8 VDD2.t3 VN.t4 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X9 VDD1.t5 VP.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X10 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=0 ps=0 w=12.49 l=1.12
X11 VTAIL.t11 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=2.06085 ps=12.82 w=12.49 l=1.12
X12 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=4.8711 ps=25.76 w=12.49 l=1.12
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=0 ps=0 w=12.49 l=1.12
X14 VTAIL.t7 VN.t6 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8711 pd=25.76 as=2.06085 ps=12.82 w=12.49 l=1.12
X15 VTAIL.t12 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X16 VDD1.t2 VP.t5 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X17 VTAIL.t8 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
X18 VDD1.t0 VP.t7 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=4.8711 ps=25.76 w=12.49 l=1.12
X19 VTAIL.t3 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.06085 pd=12.82 as=2.06085 ps=12.82 w=12.49 l=1.12
R0 B.n728 B.n727 585
R1 B.n298 B.n103 585
R2 B.n297 B.n296 585
R3 B.n295 B.n294 585
R4 B.n293 B.n292 585
R5 B.n291 B.n290 585
R6 B.n289 B.n288 585
R7 B.n287 B.n286 585
R8 B.n285 B.n284 585
R9 B.n283 B.n282 585
R10 B.n281 B.n280 585
R11 B.n279 B.n278 585
R12 B.n277 B.n276 585
R13 B.n275 B.n274 585
R14 B.n273 B.n272 585
R15 B.n271 B.n270 585
R16 B.n269 B.n268 585
R17 B.n267 B.n266 585
R18 B.n265 B.n264 585
R19 B.n263 B.n262 585
R20 B.n261 B.n260 585
R21 B.n259 B.n258 585
R22 B.n257 B.n256 585
R23 B.n255 B.n254 585
R24 B.n253 B.n252 585
R25 B.n251 B.n250 585
R26 B.n249 B.n248 585
R27 B.n247 B.n246 585
R28 B.n245 B.n244 585
R29 B.n243 B.n242 585
R30 B.n241 B.n240 585
R31 B.n239 B.n238 585
R32 B.n237 B.n236 585
R33 B.n235 B.n234 585
R34 B.n233 B.n232 585
R35 B.n231 B.n230 585
R36 B.n229 B.n228 585
R37 B.n227 B.n226 585
R38 B.n225 B.n224 585
R39 B.n223 B.n222 585
R40 B.n221 B.n220 585
R41 B.n219 B.n218 585
R42 B.n217 B.n216 585
R43 B.n214 B.n213 585
R44 B.n212 B.n211 585
R45 B.n210 B.n209 585
R46 B.n208 B.n207 585
R47 B.n206 B.n205 585
R48 B.n204 B.n203 585
R49 B.n202 B.n201 585
R50 B.n200 B.n199 585
R51 B.n198 B.n197 585
R52 B.n196 B.n195 585
R53 B.n193 B.n192 585
R54 B.n191 B.n190 585
R55 B.n189 B.n188 585
R56 B.n187 B.n186 585
R57 B.n185 B.n184 585
R58 B.n183 B.n182 585
R59 B.n181 B.n180 585
R60 B.n179 B.n178 585
R61 B.n177 B.n176 585
R62 B.n175 B.n174 585
R63 B.n173 B.n172 585
R64 B.n171 B.n170 585
R65 B.n169 B.n168 585
R66 B.n167 B.n166 585
R67 B.n165 B.n164 585
R68 B.n163 B.n162 585
R69 B.n161 B.n160 585
R70 B.n159 B.n158 585
R71 B.n157 B.n156 585
R72 B.n155 B.n154 585
R73 B.n153 B.n152 585
R74 B.n151 B.n150 585
R75 B.n149 B.n148 585
R76 B.n147 B.n146 585
R77 B.n145 B.n144 585
R78 B.n143 B.n142 585
R79 B.n141 B.n140 585
R80 B.n139 B.n138 585
R81 B.n137 B.n136 585
R82 B.n135 B.n134 585
R83 B.n133 B.n132 585
R84 B.n131 B.n130 585
R85 B.n129 B.n128 585
R86 B.n127 B.n126 585
R87 B.n125 B.n124 585
R88 B.n123 B.n122 585
R89 B.n121 B.n120 585
R90 B.n119 B.n118 585
R91 B.n117 B.n116 585
R92 B.n115 B.n114 585
R93 B.n113 B.n112 585
R94 B.n111 B.n110 585
R95 B.n109 B.n108 585
R96 B.n726 B.n55 585
R97 B.n731 B.n55 585
R98 B.n725 B.n54 585
R99 B.n732 B.n54 585
R100 B.n724 B.n723 585
R101 B.n723 B.n50 585
R102 B.n722 B.n49 585
R103 B.n738 B.n49 585
R104 B.n721 B.n48 585
R105 B.n739 B.n48 585
R106 B.n720 B.n47 585
R107 B.n740 B.n47 585
R108 B.n719 B.n718 585
R109 B.n718 B.n43 585
R110 B.n717 B.n42 585
R111 B.n746 B.n42 585
R112 B.n716 B.n41 585
R113 B.n747 B.n41 585
R114 B.n715 B.n40 585
R115 B.n748 B.n40 585
R116 B.n714 B.n713 585
R117 B.n713 B.n36 585
R118 B.n712 B.n35 585
R119 B.n754 B.n35 585
R120 B.n711 B.n34 585
R121 B.n755 B.n34 585
R122 B.n710 B.n33 585
R123 B.n756 B.n33 585
R124 B.n709 B.n708 585
R125 B.n708 B.n29 585
R126 B.n707 B.n28 585
R127 B.n762 B.n28 585
R128 B.n706 B.n27 585
R129 B.n763 B.n27 585
R130 B.n705 B.n26 585
R131 B.n764 B.n26 585
R132 B.n704 B.n703 585
R133 B.n703 B.n22 585
R134 B.n702 B.n21 585
R135 B.n770 B.n21 585
R136 B.n701 B.n20 585
R137 B.n771 B.n20 585
R138 B.n700 B.n19 585
R139 B.n772 B.n19 585
R140 B.n699 B.n698 585
R141 B.n698 B.n15 585
R142 B.n697 B.n14 585
R143 B.n778 B.n14 585
R144 B.n696 B.n13 585
R145 B.n779 B.n13 585
R146 B.n695 B.n12 585
R147 B.n780 B.n12 585
R148 B.n694 B.n693 585
R149 B.n693 B.n692 585
R150 B.n691 B.n690 585
R151 B.n691 B.n8 585
R152 B.n689 B.n7 585
R153 B.n787 B.n7 585
R154 B.n688 B.n6 585
R155 B.n788 B.n6 585
R156 B.n687 B.n5 585
R157 B.n789 B.n5 585
R158 B.n686 B.n685 585
R159 B.n685 B.n4 585
R160 B.n684 B.n299 585
R161 B.n684 B.n683 585
R162 B.n674 B.n300 585
R163 B.n301 B.n300 585
R164 B.n676 B.n675 585
R165 B.n677 B.n676 585
R166 B.n673 B.n306 585
R167 B.n306 B.n305 585
R168 B.n672 B.n671 585
R169 B.n671 B.n670 585
R170 B.n308 B.n307 585
R171 B.n309 B.n308 585
R172 B.n663 B.n662 585
R173 B.n664 B.n663 585
R174 B.n661 B.n314 585
R175 B.n314 B.n313 585
R176 B.n660 B.n659 585
R177 B.n659 B.n658 585
R178 B.n316 B.n315 585
R179 B.n317 B.n316 585
R180 B.n651 B.n650 585
R181 B.n652 B.n651 585
R182 B.n649 B.n322 585
R183 B.n322 B.n321 585
R184 B.n648 B.n647 585
R185 B.n647 B.n646 585
R186 B.n324 B.n323 585
R187 B.n325 B.n324 585
R188 B.n639 B.n638 585
R189 B.n640 B.n639 585
R190 B.n637 B.n329 585
R191 B.n333 B.n329 585
R192 B.n636 B.n635 585
R193 B.n635 B.n634 585
R194 B.n331 B.n330 585
R195 B.n332 B.n331 585
R196 B.n627 B.n626 585
R197 B.n628 B.n627 585
R198 B.n625 B.n338 585
R199 B.n338 B.n337 585
R200 B.n624 B.n623 585
R201 B.n623 B.n622 585
R202 B.n340 B.n339 585
R203 B.n341 B.n340 585
R204 B.n615 B.n614 585
R205 B.n616 B.n615 585
R206 B.n613 B.n346 585
R207 B.n346 B.n345 585
R208 B.n612 B.n611 585
R209 B.n611 B.n610 585
R210 B.n348 B.n347 585
R211 B.n349 B.n348 585
R212 B.n603 B.n602 585
R213 B.n604 B.n603 585
R214 B.n601 B.n354 585
R215 B.n354 B.n353 585
R216 B.n596 B.n595 585
R217 B.n594 B.n404 585
R218 B.n593 B.n403 585
R219 B.n598 B.n403 585
R220 B.n592 B.n591 585
R221 B.n590 B.n589 585
R222 B.n588 B.n587 585
R223 B.n586 B.n585 585
R224 B.n584 B.n583 585
R225 B.n582 B.n581 585
R226 B.n580 B.n579 585
R227 B.n578 B.n577 585
R228 B.n576 B.n575 585
R229 B.n574 B.n573 585
R230 B.n572 B.n571 585
R231 B.n570 B.n569 585
R232 B.n568 B.n567 585
R233 B.n566 B.n565 585
R234 B.n564 B.n563 585
R235 B.n562 B.n561 585
R236 B.n560 B.n559 585
R237 B.n558 B.n557 585
R238 B.n556 B.n555 585
R239 B.n554 B.n553 585
R240 B.n552 B.n551 585
R241 B.n550 B.n549 585
R242 B.n548 B.n547 585
R243 B.n546 B.n545 585
R244 B.n544 B.n543 585
R245 B.n542 B.n541 585
R246 B.n540 B.n539 585
R247 B.n538 B.n537 585
R248 B.n536 B.n535 585
R249 B.n534 B.n533 585
R250 B.n532 B.n531 585
R251 B.n530 B.n529 585
R252 B.n528 B.n527 585
R253 B.n526 B.n525 585
R254 B.n524 B.n523 585
R255 B.n522 B.n521 585
R256 B.n520 B.n519 585
R257 B.n518 B.n517 585
R258 B.n516 B.n515 585
R259 B.n514 B.n513 585
R260 B.n512 B.n511 585
R261 B.n510 B.n509 585
R262 B.n508 B.n507 585
R263 B.n506 B.n505 585
R264 B.n504 B.n503 585
R265 B.n502 B.n501 585
R266 B.n500 B.n499 585
R267 B.n498 B.n497 585
R268 B.n496 B.n495 585
R269 B.n494 B.n493 585
R270 B.n492 B.n491 585
R271 B.n490 B.n489 585
R272 B.n488 B.n487 585
R273 B.n486 B.n485 585
R274 B.n484 B.n483 585
R275 B.n482 B.n481 585
R276 B.n480 B.n479 585
R277 B.n478 B.n477 585
R278 B.n476 B.n475 585
R279 B.n474 B.n473 585
R280 B.n472 B.n471 585
R281 B.n470 B.n469 585
R282 B.n468 B.n467 585
R283 B.n466 B.n465 585
R284 B.n464 B.n463 585
R285 B.n462 B.n461 585
R286 B.n460 B.n459 585
R287 B.n458 B.n457 585
R288 B.n456 B.n455 585
R289 B.n454 B.n453 585
R290 B.n452 B.n451 585
R291 B.n450 B.n449 585
R292 B.n448 B.n447 585
R293 B.n446 B.n445 585
R294 B.n444 B.n443 585
R295 B.n442 B.n441 585
R296 B.n440 B.n439 585
R297 B.n438 B.n437 585
R298 B.n436 B.n435 585
R299 B.n434 B.n433 585
R300 B.n432 B.n431 585
R301 B.n430 B.n429 585
R302 B.n428 B.n427 585
R303 B.n426 B.n425 585
R304 B.n424 B.n423 585
R305 B.n422 B.n421 585
R306 B.n420 B.n419 585
R307 B.n418 B.n417 585
R308 B.n416 B.n415 585
R309 B.n414 B.n413 585
R310 B.n412 B.n411 585
R311 B.n356 B.n355 585
R312 B.n600 B.n599 585
R313 B.n599 B.n598 585
R314 B.n352 B.n351 585
R315 B.n353 B.n352 585
R316 B.n606 B.n605 585
R317 B.n605 B.n604 585
R318 B.n607 B.n350 585
R319 B.n350 B.n349 585
R320 B.n609 B.n608 585
R321 B.n610 B.n609 585
R322 B.n344 B.n343 585
R323 B.n345 B.n344 585
R324 B.n618 B.n617 585
R325 B.n617 B.n616 585
R326 B.n619 B.n342 585
R327 B.n342 B.n341 585
R328 B.n621 B.n620 585
R329 B.n622 B.n621 585
R330 B.n336 B.n335 585
R331 B.n337 B.n336 585
R332 B.n630 B.n629 585
R333 B.n629 B.n628 585
R334 B.n631 B.n334 585
R335 B.n334 B.n332 585
R336 B.n633 B.n632 585
R337 B.n634 B.n633 585
R338 B.n328 B.n327 585
R339 B.n333 B.n328 585
R340 B.n642 B.n641 585
R341 B.n641 B.n640 585
R342 B.n643 B.n326 585
R343 B.n326 B.n325 585
R344 B.n645 B.n644 585
R345 B.n646 B.n645 585
R346 B.n320 B.n319 585
R347 B.n321 B.n320 585
R348 B.n654 B.n653 585
R349 B.n653 B.n652 585
R350 B.n655 B.n318 585
R351 B.n318 B.n317 585
R352 B.n657 B.n656 585
R353 B.n658 B.n657 585
R354 B.n312 B.n311 585
R355 B.n313 B.n312 585
R356 B.n666 B.n665 585
R357 B.n665 B.n664 585
R358 B.n667 B.n310 585
R359 B.n310 B.n309 585
R360 B.n669 B.n668 585
R361 B.n670 B.n669 585
R362 B.n304 B.n303 585
R363 B.n305 B.n304 585
R364 B.n679 B.n678 585
R365 B.n678 B.n677 585
R366 B.n680 B.n302 585
R367 B.n302 B.n301 585
R368 B.n682 B.n681 585
R369 B.n683 B.n682 585
R370 B.n3 B.n0 585
R371 B.n4 B.n3 585
R372 B.n786 B.n1 585
R373 B.n787 B.n786 585
R374 B.n785 B.n784 585
R375 B.n785 B.n8 585
R376 B.n783 B.n9 585
R377 B.n692 B.n9 585
R378 B.n782 B.n781 585
R379 B.n781 B.n780 585
R380 B.n11 B.n10 585
R381 B.n779 B.n11 585
R382 B.n777 B.n776 585
R383 B.n778 B.n777 585
R384 B.n775 B.n16 585
R385 B.n16 B.n15 585
R386 B.n774 B.n773 585
R387 B.n773 B.n772 585
R388 B.n18 B.n17 585
R389 B.n771 B.n18 585
R390 B.n769 B.n768 585
R391 B.n770 B.n769 585
R392 B.n767 B.n23 585
R393 B.n23 B.n22 585
R394 B.n766 B.n765 585
R395 B.n765 B.n764 585
R396 B.n25 B.n24 585
R397 B.n763 B.n25 585
R398 B.n761 B.n760 585
R399 B.n762 B.n761 585
R400 B.n759 B.n30 585
R401 B.n30 B.n29 585
R402 B.n758 B.n757 585
R403 B.n757 B.n756 585
R404 B.n32 B.n31 585
R405 B.n755 B.n32 585
R406 B.n753 B.n752 585
R407 B.n754 B.n753 585
R408 B.n751 B.n37 585
R409 B.n37 B.n36 585
R410 B.n750 B.n749 585
R411 B.n749 B.n748 585
R412 B.n39 B.n38 585
R413 B.n747 B.n39 585
R414 B.n745 B.n744 585
R415 B.n746 B.n745 585
R416 B.n743 B.n44 585
R417 B.n44 B.n43 585
R418 B.n742 B.n741 585
R419 B.n741 B.n740 585
R420 B.n46 B.n45 585
R421 B.n739 B.n46 585
R422 B.n737 B.n736 585
R423 B.n738 B.n737 585
R424 B.n735 B.n51 585
R425 B.n51 B.n50 585
R426 B.n734 B.n733 585
R427 B.n733 B.n732 585
R428 B.n53 B.n52 585
R429 B.n731 B.n53 585
R430 B.n790 B.n789 585
R431 B.n788 B.n2 585
R432 B.n106 B.t19 472.435
R433 B.n104 B.t15 472.435
R434 B.n408 B.t12 472.435
R435 B.n405 B.t8 472.435
R436 B.n108 B.n53 463.671
R437 B.n728 B.n55 463.671
R438 B.n599 B.n354 463.671
R439 B.n596 B.n352 463.671
R440 B.n730 B.n729 256.663
R441 B.n730 B.n102 256.663
R442 B.n730 B.n101 256.663
R443 B.n730 B.n100 256.663
R444 B.n730 B.n99 256.663
R445 B.n730 B.n98 256.663
R446 B.n730 B.n97 256.663
R447 B.n730 B.n96 256.663
R448 B.n730 B.n95 256.663
R449 B.n730 B.n94 256.663
R450 B.n730 B.n93 256.663
R451 B.n730 B.n92 256.663
R452 B.n730 B.n91 256.663
R453 B.n730 B.n90 256.663
R454 B.n730 B.n89 256.663
R455 B.n730 B.n88 256.663
R456 B.n730 B.n87 256.663
R457 B.n730 B.n86 256.663
R458 B.n730 B.n85 256.663
R459 B.n730 B.n84 256.663
R460 B.n730 B.n83 256.663
R461 B.n730 B.n82 256.663
R462 B.n730 B.n81 256.663
R463 B.n730 B.n80 256.663
R464 B.n730 B.n79 256.663
R465 B.n730 B.n78 256.663
R466 B.n730 B.n77 256.663
R467 B.n730 B.n76 256.663
R468 B.n730 B.n75 256.663
R469 B.n730 B.n74 256.663
R470 B.n730 B.n73 256.663
R471 B.n730 B.n72 256.663
R472 B.n730 B.n71 256.663
R473 B.n730 B.n70 256.663
R474 B.n730 B.n69 256.663
R475 B.n730 B.n68 256.663
R476 B.n730 B.n67 256.663
R477 B.n730 B.n66 256.663
R478 B.n730 B.n65 256.663
R479 B.n730 B.n64 256.663
R480 B.n730 B.n63 256.663
R481 B.n730 B.n62 256.663
R482 B.n730 B.n61 256.663
R483 B.n730 B.n60 256.663
R484 B.n730 B.n59 256.663
R485 B.n730 B.n58 256.663
R486 B.n730 B.n57 256.663
R487 B.n730 B.n56 256.663
R488 B.n598 B.n597 256.663
R489 B.n598 B.n357 256.663
R490 B.n598 B.n358 256.663
R491 B.n598 B.n359 256.663
R492 B.n598 B.n360 256.663
R493 B.n598 B.n361 256.663
R494 B.n598 B.n362 256.663
R495 B.n598 B.n363 256.663
R496 B.n598 B.n364 256.663
R497 B.n598 B.n365 256.663
R498 B.n598 B.n366 256.663
R499 B.n598 B.n367 256.663
R500 B.n598 B.n368 256.663
R501 B.n598 B.n369 256.663
R502 B.n598 B.n370 256.663
R503 B.n598 B.n371 256.663
R504 B.n598 B.n372 256.663
R505 B.n598 B.n373 256.663
R506 B.n598 B.n374 256.663
R507 B.n598 B.n375 256.663
R508 B.n598 B.n376 256.663
R509 B.n598 B.n377 256.663
R510 B.n598 B.n378 256.663
R511 B.n598 B.n379 256.663
R512 B.n598 B.n380 256.663
R513 B.n598 B.n381 256.663
R514 B.n598 B.n382 256.663
R515 B.n598 B.n383 256.663
R516 B.n598 B.n384 256.663
R517 B.n598 B.n385 256.663
R518 B.n598 B.n386 256.663
R519 B.n598 B.n387 256.663
R520 B.n598 B.n388 256.663
R521 B.n598 B.n389 256.663
R522 B.n598 B.n390 256.663
R523 B.n598 B.n391 256.663
R524 B.n598 B.n392 256.663
R525 B.n598 B.n393 256.663
R526 B.n598 B.n394 256.663
R527 B.n598 B.n395 256.663
R528 B.n598 B.n396 256.663
R529 B.n598 B.n397 256.663
R530 B.n598 B.n398 256.663
R531 B.n598 B.n399 256.663
R532 B.n598 B.n400 256.663
R533 B.n598 B.n401 256.663
R534 B.n598 B.n402 256.663
R535 B.n792 B.n791 256.663
R536 B.n112 B.n111 163.367
R537 B.n116 B.n115 163.367
R538 B.n120 B.n119 163.367
R539 B.n124 B.n123 163.367
R540 B.n128 B.n127 163.367
R541 B.n132 B.n131 163.367
R542 B.n136 B.n135 163.367
R543 B.n140 B.n139 163.367
R544 B.n144 B.n143 163.367
R545 B.n148 B.n147 163.367
R546 B.n152 B.n151 163.367
R547 B.n156 B.n155 163.367
R548 B.n160 B.n159 163.367
R549 B.n164 B.n163 163.367
R550 B.n168 B.n167 163.367
R551 B.n172 B.n171 163.367
R552 B.n176 B.n175 163.367
R553 B.n180 B.n179 163.367
R554 B.n184 B.n183 163.367
R555 B.n188 B.n187 163.367
R556 B.n192 B.n191 163.367
R557 B.n197 B.n196 163.367
R558 B.n201 B.n200 163.367
R559 B.n205 B.n204 163.367
R560 B.n209 B.n208 163.367
R561 B.n213 B.n212 163.367
R562 B.n218 B.n217 163.367
R563 B.n222 B.n221 163.367
R564 B.n226 B.n225 163.367
R565 B.n230 B.n229 163.367
R566 B.n234 B.n233 163.367
R567 B.n238 B.n237 163.367
R568 B.n242 B.n241 163.367
R569 B.n246 B.n245 163.367
R570 B.n250 B.n249 163.367
R571 B.n254 B.n253 163.367
R572 B.n258 B.n257 163.367
R573 B.n262 B.n261 163.367
R574 B.n266 B.n265 163.367
R575 B.n270 B.n269 163.367
R576 B.n274 B.n273 163.367
R577 B.n278 B.n277 163.367
R578 B.n282 B.n281 163.367
R579 B.n286 B.n285 163.367
R580 B.n290 B.n289 163.367
R581 B.n294 B.n293 163.367
R582 B.n296 B.n103 163.367
R583 B.n603 B.n354 163.367
R584 B.n603 B.n348 163.367
R585 B.n611 B.n348 163.367
R586 B.n611 B.n346 163.367
R587 B.n615 B.n346 163.367
R588 B.n615 B.n340 163.367
R589 B.n623 B.n340 163.367
R590 B.n623 B.n338 163.367
R591 B.n627 B.n338 163.367
R592 B.n627 B.n331 163.367
R593 B.n635 B.n331 163.367
R594 B.n635 B.n329 163.367
R595 B.n639 B.n329 163.367
R596 B.n639 B.n324 163.367
R597 B.n647 B.n324 163.367
R598 B.n647 B.n322 163.367
R599 B.n651 B.n322 163.367
R600 B.n651 B.n316 163.367
R601 B.n659 B.n316 163.367
R602 B.n659 B.n314 163.367
R603 B.n663 B.n314 163.367
R604 B.n663 B.n308 163.367
R605 B.n671 B.n308 163.367
R606 B.n671 B.n306 163.367
R607 B.n676 B.n306 163.367
R608 B.n676 B.n300 163.367
R609 B.n684 B.n300 163.367
R610 B.n685 B.n684 163.367
R611 B.n685 B.n5 163.367
R612 B.n6 B.n5 163.367
R613 B.n7 B.n6 163.367
R614 B.n691 B.n7 163.367
R615 B.n693 B.n691 163.367
R616 B.n693 B.n12 163.367
R617 B.n13 B.n12 163.367
R618 B.n14 B.n13 163.367
R619 B.n698 B.n14 163.367
R620 B.n698 B.n19 163.367
R621 B.n20 B.n19 163.367
R622 B.n21 B.n20 163.367
R623 B.n703 B.n21 163.367
R624 B.n703 B.n26 163.367
R625 B.n27 B.n26 163.367
R626 B.n28 B.n27 163.367
R627 B.n708 B.n28 163.367
R628 B.n708 B.n33 163.367
R629 B.n34 B.n33 163.367
R630 B.n35 B.n34 163.367
R631 B.n713 B.n35 163.367
R632 B.n713 B.n40 163.367
R633 B.n41 B.n40 163.367
R634 B.n42 B.n41 163.367
R635 B.n718 B.n42 163.367
R636 B.n718 B.n47 163.367
R637 B.n48 B.n47 163.367
R638 B.n49 B.n48 163.367
R639 B.n723 B.n49 163.367
R640 B.n723 B.n54 163.367
R641 B.n55 B.n54 163.367
R642 B.n404 B.n403 163.367
R643 B.n591 B.n403 163.367
R644 B.n589 B.n588 163.367
R645 B.n585 B.n584 163.367
R646 B.n581 B.n580 163.367
R647 B.n577 B.n576 163.367
R648 B.n573 B.n572 163.367
R649 B.n569 B.n568 163.367
R650 B.n565 B.n564 163.367
R651 B.n561 B.n560 163.367
R652 B.n557 B.n556 163.367
R653 B.n553 B.n552 163.367
R654 B.n549 B.n548 163.367
R655 B.n545 B.n544 163.367
R656 B.n541 B.n540 163.367
R657 B.n537 B.n536 163.367
R658 B.n533 B.n532 163.367
R659 B.n529 B.n528 163.367
R660 B.n525 B.n524 163.367
R661 B.n521 B.n520 163.367
R662 B.n517 B.n516 163.367
R663 B.n513 B.n512 163.367
R664 B.n509 B.n508 163.367
R665 B.n505 B.n504 163.367
R666 B.n501 B.n500 163.367
R667 B.n497 B.n496 163.367
R668 B.n493 B.n492 163.367
R669 B.n489 B.n488 163.367
R670 B.n485 B.n484 163.367
R671 B.n481 B.n480 163.367
R672 B.n477 B.n476 163.367
R673 B.n473 B.n472 163.367
R674 B.n469 B.n468 163.367
R675 B.n465 B.n464 163.367
R676 B.n461 B.n460 163.367
R677 B.n457 B.n456 163.367
R678 B.n453 B.n452 163.367
R679 B.n449 B.n448 163.367
R680 B.n445 B.n444 163.367
R681 B.n441 B.n440 163.367
R682 B.n437 B.n436 163.367
R683 B.n433 B.n432 163.367
R684 B.n429 B.n428 163.367
R685 B.n425 B.n424 163.367
R686 B.n421 B.n420 163.367
R687 B.n417 B.n416 163.367
R688 B.n413 B.n412 163.367
R689 B.n599 B.n356 163.367
R690 B.n605 B.n352 163.367
R691 B.n605 B.n350 163.367
R692 B.n609 B.n350 163.367
R693 B.n609 B.n344 163.367
R694 B.n617 B.n344 163.367
R695 B.n617 B.n342 163.367
R696 B.n621 B.n342 163.367
R697 B.n621 B.n336 163.367
R698 B.n629 B.n336 163.367
R699 B.n629 B.n334 163.367
R700 B.n633 B.n334 163.367
R701 B.n633 B.n328 163.367
R702 B.n641 B.n328 163.367
R703 B.n641 B.n326 163.367
R704 B.n645 B.n326 163.367
R705 B.n645 B.n320 163.367
R706 B.n653 B.n320 163.367
R707 B.n653 B.n318 163.367
R708 B.n657 B.n318 163.367
R709 B.n657 B.n312 163.367
R710 B.n665 B.n312 163.367
R711 B.n665 B.n310 163.367
R712 B.n669 B.n310 163.367
R713 B.n669 B.n304 163.367
R714 B.n678 B.n304 163.367
R715 B.n678 B.n302 163.367
R716 B.n682 B.n302 163.367
R717 B.n682 B.n3 163.367
R718 B.n790 B.n3 163.367
R719 B.n786 B.n2 163.367
R720 B.n786 B.n785 163.367
R721 B.n785 B.n9 163.367
R722 B.n781 B.n9 163.367
R723 B.n781 B.n11 163.367
R724 B.n777 B.n11 163.367
R725 B.n777 B.n16 163.367
R726 B.n773 B.n16 163.367
R727 B.n773 B.n18 163.367
R728 B.n769 B.n18 163.367
R729 B.n769 B.n23 163.367
R730 B.n765 B.n23 163.367
R731 B.n765 B.n25 163.367
R732 B.n761 B.n25 163.367
R733 B.n761 B.n30 163.367
R734 B.n757 B.n30 163.367
R735 B.n757 B.n32 163.367
R736 B.n753 B.n32 163.367
R737 B.n753 B.n37 163.367
R738 B.n749 B.n37 163.367
R739 B.n749 B.n39 163.367
R740 B.n745 B.n39 163.367
R741 B.n745 B.n44 163.367
R742 B.n741 B.n44 163.367
R743 B.n741 B.n46 163.367
R744 B.n737 B.n46 163.367
R745 B.n737 B.n51 163.367
R746 B.n733 B.n51 163.367
R747 B.n733 B.n53 163.367
R748 B.n104 B.t17 100.695
R749 B.n408 B.t14 100.695
R750 B.n106 B.t20 100.68
R751 B.n405 B.t11 100.68
R752 B.n598 B.n353 73.6847
R753 B.n731 B.n730 73.6847
R754 B.n105 B.t18 72.5741
R755 B.n409 B.t13 72.5741
R756 B.n107 B.t21 72.5584
R757 B.n406 B.t10 72.5584
R758 B.n108 B.n56 71.676
R759 B.n112 B.n57 71.676
R760 B.n116 B.n58 71.676
R761 B.n120 B.n59 71.676
R762 B.n124 B.n60 71.676
R763 B.n128 B.n61 71.676
R764 B.n132 B.n62 71.676
R765 B.n136 B.n63 71.676
R766 B.n140 B.n64 71.676
R767 B.n144 B.n65 71.676
R768 B.n148 B.n66 71.676
R769 B.n152 B.n67 71.676
R770 B.n156 B.n68 71.676
R771 B.n160 B.n69 71.676
R772 B.n164 B.n70 71.676
R773 B.n168 B.n71 71.676
R774 B.n172 B.n72 71.676
R775 B.n176 B.n73 71.676
R776 B.n180 B.n74 71.676
R777 B.n184 B.n75 71.676
R778 B.n188 B.n76 71.676
R779 B.n192 B.n77 71.676
R780 B.n197 B.n78 71.676
R781 B.n201 B.n79 71.676
R782 B.n205 B.n80 71.676
R783 B.n209 B.n81 71.676
R784 B.n213 B.n82 71.676
R785 B.n218 B.n83 71.676
R786 B.n222 B.n84 71.676
R787 B.n226 B.n85 71.676
R788 B.n230 B.n86 71.676
R789 B.n234 B.n87 71.676
R790 B.n238 B.n88 71.676
R791 B.n242 B.n89 71.676
R792 B.n246 B.n90 71.676
R793 B.n250 B.n91 71.676
R794 B.n254 B.n92 71.676
R795 B.n258 B.n93 71.676
R796 B.n262 B.n94 71.676
R797 B.n266 B.n95 71.676
R798 B.n270 B.n96 71.676
R799 B.n274 B.n97 71.676
R800 B.n278 B.n98 71.676
R801 B.n282 B.n99 71.676
R802 B.n286 B.n100 71.676
R803 B.n290 B.n101 71.676
R804 B.n294 B.n102 71.676
R805 B.n729 B.n103 71.676
R806 B.n729 B.n728 71.676
R807 B.n296 B.n102 71.676
R808 B.n293 B.n101 71.676
R809 B.n289 B.n100 71.676
R810 B.n285 B.n99 71.676
R811 B.n281 B.n98 71.676
R812 B.n277 B.n97 71.676
R813 B.n273 B.n96 71.676
R814 B.n269 B.n95 71.676
R815 B.n265 B.n94 71.676
R816 B.n261 B.n93 71.676
R817 B.n257 B.n92 71.676
R818 B.n253 B.n91 71.676
R819 B.n249 B.n90 71.676
R820 B.n245 B.n89 71.676
R821 B.n241 B.n88 71.676
R822 B.n237 B.n87 71.676
R823 B.n233 B.n86 71.676
R824 B.n229 B.n85 71.676
R825 B.n225 B.n84 71.676
R826 B.n221 B.n83 71.676
R827 B.n217 B.n82 71.676
R828 B.n212 B.n81 71.676
R829 B.n208 B.n80 71.676
R830 B.n204 B.n79 71.676
R831 B.n200 B.n78 71.676
R832 B.n196 B.n77 71.676
R833 B.n191 B.n76 71.676
R834 B.n187 B.n75 71.676
R835 B.n183 B.n74 71.676
R836 B.n179 B.n73 71.676
R837 B.n175 B.n72 71.676
R838 B.n171 B.n71 71.676
R839 B.n167 B.n70 71.676
R840 B.n163 B.n69 71.676
R841 B.n159 B.n68 71.676
R842 B.n155 B.n67 71.676
R843 B.n151 B.n66 71.676
R844 B.n147 B.n65 71.676
R845 B.n143 B.n64 71.676
R846 B.n139 B.n63 71.676
R847 B.n135 B.n62 71.676
R848 B.n131 B.n61 71.676
R849 B.n127 B.n60 71.676
R850 B.n123 B.n59 71.676
R851 B.n119 B.n58 71.676
R852 B.n115 B.n57 71.676
R853 B.n111 B.n56 71.676
R854 B.n597 B.n596 71.676
R855 B.n591 B.n357 71.676
R856 B.n588 B.n358 71.676
R857 B.n584 B.n359 71.676
R858 B.n580 B.n360 71.676
R859 B.n576 B.n361 71.676
R860 B.n572 B.n362 71.676
R861 B.n568 B.n363 71.676
R862 B.n564 B.n364 71.676
R863 B.n560 B.n365 71.676
R864 B.n556 B.n366 71.676
R865 B.n552 B.n367 71.676
R866 B.n548 B.n368 71.676
R867 B.n544 B.n369 71.676
R868 B.n540 B.n370 71.676
R869 B.n536 B.n371 71.676
R870 B.n532 B.n372 71.676
R871 B.n528 B.n373 71.676
R872 B.n524 B.n374 71.676
R873 B.n520 B.n375 71.676
R874 B.n516 B.n376 71.676
R875 B.n512 B.n377 71.676
R876 B.n508 B.n378 71.676
R877 B.n504 B.n379 71.676
R878 B.n500 B.n380 71.676
R879 B.n496 B.n381 71.676
R880 B.n492 B.n382 71.676
R881 B.n488 B.n383 71.676
R882 B.n484 B.n384 71.676
R883 B.n480 B.n385 71.676
R884 B.n476 B.n386 71.676
R885 B.n472 B.n387 71.676
R886 B.n468 B.n388 71.676
R887 B.n464 B.n389 71.676
R888 B.n460 B.n390 71.676
R889 B.n456 B.n391 71.676
R890 B.n452 B.n392 71.676
R891 B.n448 B.n393 71.676
R892 B.n444 B.n394 71.676
R893 B.n440 B.n395 71.676
R894 B.n436 B.n396 71.676
R895 B.n432 B.n397 71.676
R896 B.n428 B.n398 71.676
R897 B.n424 B.n399 71.676
R898 B.n420 B.n400 71.676
R899 B.n416 B.n401 71.676
R900 B.n412 B.n402 71.676
R901 B.n597 B.n404 71.676
R902 B.n589 B.n357 71.676
R903 B.n585 B.n358 71.676
R904 B.n581 B.n359 71.676
R905 B.n577 B.n360 71.676
R906 B.n573 B.n361 71.676
R907 B.n569 B.n362 71.676
R908 B.n565 B.n363 71.676
R909 B.n561 B.n364 71.676
R910 B.n557 B.n365 71.676
R911 B.n553 B.n366 71.676
R912 B.n549 B.n367 71.676
R913 B.n545 B.n368 71.676
R914 B.n541 B.n369 71.676
R915 B.n537 B.n370 71.676
R916 B.n533 B.n371 71.676
R917 B.n529 B.n372 71.676
R918 B.n525 B.n373 71.676
R919 B.n521 B.n374 71.676
R920 B.n517 B.n375 71.676
R921 B.n513 B.n376 71.676
R922 B.n509 B.n377 71.676
R923 B.n505 B.n378 71.676
R924 B.n501 B.n379 71.676
R925 B.n497 B.n380 71.676
R926 B.n493 B.n381 71.676
R927 B.n489 B.n382 71.676
R928 B.n485 B.n383 71.676
R929 B.n481 B.n384 71.676
R930 B.n477 B.n385 71.676
R931 B.n473 B.n386 71.676
R932 B.n469 B.n387 71.676
R933 B.n465 B.n388 71.676
R934 B.n461 B.n389 71.676
R935 B.n457 B.n390 71.676
R936 B.n453 B.n391 71.676
R937 B.n449 B.n392 71.676
R938 B.n445 B.n393 71.676
R939 B.n441 B.n394 71.676
R940 B.n437 B.n395 71.676
R941 B.n433 B.n396 71.676
R942 B.n429 B.n397 71.676
R943 B.n425 B.n398 71.676
R944 B.n421 B.n399 71.676
R945 B.n417 B.n400 71.676
R946 B.n413 B.n401 71.676
R947 B.n402 B.n356 71.676
R948 B.n791 B.n790 71.676
R949 B.n791 B.n2 71.676
R950 B.n194 B.n107 59.5399
R951 B.n215 B.n105 59.5399
R952 B.n410 B.n409 59.5399
R953 B.n407 B.n406 59.5399
R954 B.n604 B.n353 42.1058
R955 B.n604 B.n349 42.1058
R956 B.n610 B.n349 42.1058
R957 B.n610 B.n345 42.1058
R958 B.n616 B.n345 42.1058
R959 B.n622 B.n341 42.1058
R960 B.n622 B.n337 42.1058
R961 B.n628 B.n337 42.1058
R962 B.n628 B.n332 42.1058
R963 B.n634 B.n332 42.1058
R964 B.n634 B.n333 42.1058
R965 B.n640 B.n325 42.1058
R966 B.n646 B.n325 42.1058
R967 B.n646 B.n321 42.1058
R968 B.n652 B.n321 42.1058
R969 B.n658 B.n317 42.1058
R970 B.n658 B.n313 42.1058
R971 B.n664 B.n313 42.1058
R972 B.n670 B.n309 42.1058
R973 B.n670 B.n305 42.1058
R974 B.n677 B.n305 42.1058
R975 B.n683 B.n301 42.1058
R976 B.n683 B.n4 42.1058
R977 B.n789 B.n4 42.1058
R978 B.n789 B.n788 42.1058
R979 B.n788 B.n787 42.1058
R980 B.n787 B.n8 42.1058
R981 B.n692 B.n8 42.1058
R982 B.n780 B.n779 42.1058
R983 B.n779 B.n778 42.1058
R984 B.n778 B.n15 42.1058
R985 B.n772 B.n771 42.1058
R986 B.n771 B.n770 42.1058
R987 B.n770 B.n22 42.1058
R988 B.n764 B.n763 42.1058
R989 B.n763 B.n762 42.1058
R990 B.n762 B.n29 42.1058
R991 B.n756 B.n29 42.1058
R992 B.n755 B.n754 42.1058
R993 B.n754 B.n36 42.1058
R994 B.n748 B.n36 42.1058
R995 B.n748 B.n747 42.1058
R996 B.n747 B.n746 42.1058
R997 B.n746 B.n43 42.1058
R998 B.n740 B.n739 42.1058
R999 B.n739 B.n738 42.1058
R1000 B.n738 B.n50 42.1058
R1001 B.n732 B.n50 42.1058
R1002 B.n732 B.n731 42.1058
R1003 B.n333 B.t7 40.8674
R1004 B.t6 B.n755 40.8674
R1005 B.t3 B.n317 32.1986
R1006 B.n677 B.t0 32.1986
R1007 B.n780 B.t2 32.1986
R1008 B.t5 B.n22 32.1986
R1009 B.n595 B.n351 30.1273
R1010 B.n601 B.n600 30.1273
R1011 B.n727 B.n726 30.1273
R1012 B.n109 B.n52 30.1273
R1013 B.n107 B.n106 28.1217
R1014 B.n105 B.n104 28.1217
R1015 B.n409 B.n408 28.1217
R1016 B.n406 B.n405 28.1217
R1017 B.n616 B.t9 21.0531
R1018 B.t9 B.n341 21.0531
R1019 B.n664 B.t4 21.0531
R1020 B.t4 B.n309 21.0531
R1021 B.t1 B.n15 21.0531
R1022 B.n772 B.t1 21.0531
R1023 B.t16 B.n43 21.0531
R1024 B.n740 B.t16 21.0531
R1025 B B.n792 18.0485
R1026 B.n606 B.n351 10.6151
R1027 B.n607 B.n606 10.6151
R1028 B.n608 B.n607 10.6151
R1029 B.n608 B.n343 10.6151
R1030 B.n618 B.n343 10.6151
R1031 B.n619 B.n618 10.6151
R1032 B.n620 B.n619 10.6151
R1033 B.n620 B.n335 10.6151
R1034 B.n630 B.n335 10.6151
R1035 B.n631 B.n630 10.6151
R1036 B.n632 B.n631 10.6151
R1037 B.n632 B.n327 10.6151
R1038 B.n642 B.n327 10.6151
R1039 B.n643 B.n642 10.6151
R1040 B.n644 B.n643 10.6151
R1041 B.n644 B.n319 10.6151
R1042 B.n654 B.n319 10.6151
R1043 B.n655 B.n654 10.6151
R1044 B.n656 B.n655 10.6151
R1045 B.n656 B.n311 10.6151
R1046 B.n666 B.n311 10.6151
R1047 B.n667 B.n666 10.6151
R1048 B.n668 B.n667 10.6151
R1049 B.n668 B.n303 10.6151
R1050 B.n679 B.n303 10.6151
R1051 B.n680 B.n679 10.6151
R1052 B.n681 B.n680 10.6151
R1053 B.n681 B.n0 10.6151
R1054 B.n595 B.n594 10.6151
R1055 B.n594 B.n593 10.6151
R1056 B.n593 B.n592 10.6151
R1057 B.n592 B.n590 10.6151
R1058 B.n590 B.n587 10.6151
R1059 B.n587 B.n586 10.6151
R1060 B.n586 B.n583 10.6151
R1061 B.n583 B.n582 10.6151
R1062 B.n582 B.n579 10.6151
R1063 B.n579 B.n578 10.6151
R1064 B.n578 B.n575 10.6151
R1065 B.n575 B.n574 10.6151
R1066 B.n574 B.n571 10.6151
R1067 B.n571 B.n570 10.6151
R1068 B.n570 B.n567 10.6151
R1069 B.n567 B.n566 10.6151
R1070 B.n566 B.n563 10.6151
R1071 B.n563 B.n562 10.6151
R1072 B.n562 B.n559 10.6151
R1073 B.n559 B.n558 10.6151
R1074 B.n558 B.n555 10.6151
R1075 B.n555 B.n554 10.6151
R1076 B.n554 B.n551 10.6151
R1077 B.n551 B.n550 10.6151
R1078 B.n550 B.n547 10.6151
R1079 B.n547 B.n546 10.6151
R1080 B.n546 B.n543 10.6151
R1081 B.n543 B.n542 10.6151
R1082 B.n542 B.n539 10.6151
R1083 B.n539 B.n538 10.6151
R1084 B.n538 B.n535 10.6151
R1085 B.n535 B.n534 10.6151
R1086 B.n534 B.n531 10.6151
R1087 B.n531 B.n530 10.6151
R1088 B.n530 B.n527 10.6151
R1089 B.n527 B.n526 10.6151
R1090 B.n526 B.n523 10.6151
R1091 B.n523 B.n522 10.6151
R1092 B.n522 B.n519 10.6151
R1093 B.n519 B.n518 10.6151
R1094 B.n518 B.n515 10.6151
R1095 B.n515 B.n514 10.6151
R1096 B.n511 B.n510 10.6151
R1097 B.n510 B.n507 10.6151
R1098 B.n507 B.n506 10.6151
R1099 B.n506 B.n503 10.6151
R1100 B.n503 B.n502 10.6151
R1101 B.n502 B.n499 10.6151
R1102 B.n499 B.n498 10.6151
R1103 B.n498 B.n495 10.6151
R1104 B.n495 B.n494 10.6151
R1105 B.n491 B.n490 10.6151
R1106 B.n490 B.n487 10.6151
R1107 B.n487 B.n486 10.6151
R1108 B.n486 B.n483 10.6151
R1109 B.n483 B.n482 10.6151
R1110 B.n482 B.n479 10.6151
R1111 B.n479 B.n478 10.6151
R1112 B.n478 B.n475 10.6151
R1113 B.n475 B.n474 10.6151
R1114 B.n474 B.n471 10.6151
R1115 B.n471 B.n470 10.6151
R1116 B.n470 B.n467 10.6151
R1117 B.n467 B.n466 10.6151
R1118 B.n466 B.n463 10.6151
R1119 B.n463 B.n462 10.6151
R1120 B.n462 B.n459 10.6151
R1121 B.n459 B.n458 10.6151
R1122 B.n458 B.n455 10.6151
R1123 B.n455 B.n454 10.6151
R1124 B.n454 B.n451 10.6151
R1125 B.n451 B.n450 10.6151
R1126 B.n450 B.n447 10.6151
R1127 B.n447 B.n446 10.6151
R1128 B.n446 B.n443 10.6151
R1129 B.n443 B.n442 10.6151
R1130 B.n442 B.n439 10.6151
R1131 B.n439 B.n438 10.6151
R1132 B.n438 B.n435 10.6151
R1133 B.n435 B.n434 10.6151
R1134 B.n434 B.n431 10.6151
R1135 B.n431 B.n430 10.6151
R1136 B.n430 B.n427 10.6151
R1137 B.n427 B.n426 10.6151
R1138 B.n426 B.n423 10.6151
R1139 B.n423 B.n422 10.6151
R1140 B.n422 B.n419 10.6151
R1141 B.n419 B.n418 10.6151
R1142 B.n418 B.n415 10.6151
R1143 B.n415 B.n414 10.6151
R1144 B.n414 B.n411 10.6151
R1145 B.n411 B.n355 10.6151
R1146 B.n600 B.n355 10.6151
R1147 B.n602 B.n601 10.6151
R1148 B.n602 B.n347 10.6151
R1149 B.n612 B.n347 10.6151
R1150 B.n613 B.n612 10.6151
R1151 B.n614 B.n613 10.6151
R1152 B.n614 B.n339 10.6151
R1153 B.n624 B.n339 10.6151
R1154 B.n625 B.n624 10.6151
R1155 B.n626 B.n625 10.6151
R1156 B.n626 B.n330 10.6151
R1157 B.n636 B.n330 10.6151
R1158 B.n637 B.n636 10.6151
R1159 B.n638 B.n637 10.6151
R1160 B.n638 B.n323 10.6151
R1161 B.n648 B.n323 10.6151
R1162 B.n649 B.n648 10.6151
R1163 B.n650 B.n649 10.6151
R1164 B.n650 B.n315 10.6151
R1165 B.n660 B.n315 10.6151
R1166 B.n661 B.n660 10.6151
R1167 B.n662 B.n661 10.6151
R1168 B.n662 B.n307 10.6151
R1169 B.n672 B.n307 10.6151
R1170 B.n673 B.n672 10.6151
R1171 B.n675 B.n673 10.6151
R1172 B.n675 B.n674 10.6151
R1173 B.n674 B.n299 10.6151
R1174 B.n686 B.n299 10.6151
R1175 B.n687 B.n686 10.6151
R1176 B.n688 B.n687 10.6151
R1177 B.n689 B.n688 10.6151
R1178 B.n690 B.n689 10.6151
R1179 B.n694 B.n690 10.6151
R1180 B.n695 B.n694 10.6151
R1181 B.n696 B.n695 10.6151
R1182 B.n697 B.n696 10.6151
R1183 B.n699 B.n697 10.6151
R1184 B.n700 B.n699 10.6151
R1185 B.n701 B.n700 10.6151
R1186 B.n702 B.n701 10.6151
R1187 B.n704 B.n702 10.6151
R1188 B.n705 B.n704 10.6151
R1189 B.n706 B.n705 10.6151
R1190 B.n707 B.n706 10.6151
R1191 B.n709 B.n707 10.6151
R1192 B.n710 B.n709 10.6151
R1193 B.n711 B.n710 10.6151
R1194 B.n712 B.n711 10.6151
R1195 B.n714 B.n712 10.6151
R1196 B.n715 B.n714 10.6151
R1197 B.n716 B.n715 10.6151
R1198 B.n717 B.n716 10.6151
R1199 B.n719 B.n717 10.6151
R1200 B.n720 B.n719 10.6151
R1201 B.n721 B.n720 10.6151
R1202 B.n722 B.n721 10.6151
R1203 B.n724 B.n722 10.6151
R1204 B.n725 B.n724 10.6151
R1205 B.n726 B.n725 10.6151
R1206 B.n784 B.n1 10.6151
R1207 B.n784 B.n783 10.6151
R1208 B.n783 B.n782 10.6151
R1209 B.n782 B.n10 10.6151
R1210 B.n776 B.n10 10.6151
R1211 B.n776 B.n775 10.6151
R1212 B.n775 B.n774 10.6151
R1213 B.n774 B.n17 10.6151
R1214 B.n768 B.n17 10.6151
R1215 B.n768 B.n767 10.6151
R1216 B.n767 B.n766 10.6151
R1217 B.n766 B.n24 10.6151
R1218 B.n760 B.n24 10.6151
R1219 B.n760 B.n759 10.6151
R1220 B.n759 B.n758 10.6151
R1221 B.n758 B.n31 10.6151
R1222 B.n752 B.n31 10.6151
R1223 B.n752 B.n751 10.6151
R1224 B.n751 B.n750 10.6151
R1225 B.n750 B.n38 10.6151
R1226 B.n744 B.n38 10.6151
R1227 B.n744 B.n743 10.6151
R1228 B.n743 B.n742 10.6151
R1229 B.n742 B.n45 10.6151
R1230 B.n736 B.n45 10.6151
R1231 B.n736 B.n735 10.6151
R1232 B.n735 B.n734 10.6151
R1233 B.n734 B.n52 10.6151
R1234 B.n110 B.n109 10.6151
R1235 B.n113 B.n110 10.6151
R1236 B.n114 B.n113 10.6151
R1237 B.n117 B.n114 10.6151
R1238 B.n118 B.n117 10.6151
R1239 B.n121 B.n118 10.6151
R1240 B.n122 B.n121 10.6151
R1241 B.n125 B.n122 10.6151
R1242 B.n126 B.n125 10.6151
R1243 B.n129 B.n126 10.6151
R1244 B.n130 B.n129 10.6151
R1245 B.n133 B.n130 10.6151
R1246 B.n134 B.n133 10.6151
R1247 B.n137 B.n134 10.6151
R1248 B.n138 B.n137 10.6151
R1249 B.n141 B.n138 10.6151
R1250 B.n142 B.n141 10.6151
R1251 B.n145 B.n142 10.6151
R1252 B.n146 B.n145 10.6151
R1253 B.n149 B.n146 10.6151
R1254 B.n150 B.n149 10.6151
R1255 B.n153 B.n150 10.6151
R1256 B.n154 B.n153 10.6151
R1257 B.n157 B.n154 10.6151
R1258 B.n158 B.n157 10.6151
R1259 B.n161 B.n158 10.6151
R1260 B.n162 B.n161 10.6151
R1261 B.n165 B.n162 10.6151
R1262 B.n166 B.n165 10.6151
R1263 B.n169 B.n166 10.6151
R1264 B.n170 B.n169 10.6151
R1265 B.n173 B.n170 10.6151
R1266 B.n174 B.n173 10.6151
R1267 B.n177 B.n174 10.6151
R1268 B.n178 B.n177 10.6151
R1269 B.n181 B.n178 10.6151
R1270 B.n182 B.n181 10.6151
R1271 B.n185 B.n182 10.6151
R1272 B.n186 B.n185 10.6151
R1273 B.n189 B.n186 10.6151
R1274 B.n190 B.n189 10.6151
R1275 B.n193 B.n190 10.6151
R1276 B.n198 B.n195 10.6151
R1277 B.n199 B.n198 10.6151
R1278 B.n202 B.n199 10.6151
R1279 B.n203 B.n202 10.6151
R1280 B.n206 B.n203 10.6151
R1281 B.n207 B.n206 10.6151
R1282 B.n210 B.n207 10.6151
R1283 B.n211 B.n210 10.6151
R1284 B.n214 B.n211 10.6151
R1285 B.n219 B.n216 10.6151
R1286 B.n220 B.n219 10.6151
R1287 B.n223 B.n220 10.6151
R1288 B.n224 B.n223 10.6151
R1289 B.n227 B.n224 10.6151
R1290 B.n228 B.n227 10.6151
R1291 B.n231 B.n228 10.6151
R1292 B.n232 B.n231 10.6151
R1293 B.n235 B.n232 10.6151
R1294 B.n236 B.n235 10.6151
R1295 B.n239 B.n236 10.6151
R1296 B.n240 B.n239 10.6151
R1297 B.n243 B.n240 10.6151
R1298 B.n244 B.n243 10.6151
R1299 B.n247 B.n244 10.6151
R1300 B.n248 B.n247 10.6151
R1301 B.n251 B.n248 10.6151
R1302 B.n252 B.n251 10.6151
R1303 B.n255 B.n252 10.6151
R1304 B.n256 B.n255 10.6151
R1305 B.n259 B.n256 10.6151
R1306 B.n260 B.n259 10.6151
R1307 B.n263 B.n260 10.6151
R1308 B.n264 B.n263 10.6151
R1309 B.n267 B.n264 10.6151
R1310 B.n268 B.n267 10.6151
R1311 B.n271 B.n268 10.6151
R1312 B.n272 B.n271 10.6151
R1313 B.n275 B.n272 10.6151
R1314 B.n276 B.n275 10.6151
R1315 B.n279 B.n276 10.6151
R1316 B.n280 B.n279 10.6151
R1317 B.n283 B.n280 10.6151
R1318 B.n284 B.n283 10.6151
R1319 B.n287 B.n284 10.6151
R1320 B.n288 B.n287 10.6151
R1321 B.n291 B.n288 10.6151
R1322 B.n292 B.n291 10.6151
R1323 B.n295 B.n292 10.6151
R1324 B.n297 B.n295 10.6151
R1325 B.n298 B.n297 10.6151
R1326 B.n727 B.n298 10.6151
R1327 B.n652 B.t3 9.90762
R1328 B.t0 B.n301 9.90762
R1329 B.n692 B.t2 9.90762
R1330 B.n764 B.t5 9.90762
R1331 B.n514 B.n407 9.36635
R1332 B.n491 B.n410 9.36635
R1333 B.n194 B.n193 9.36635
R1334 B.n216 B.n215 9.36635
R1335 B.n792 B.n0 8.11757
R1336 B.n792 B.n1 8.11757
R1337 B.n511 B.n407 1.24928
R1338 B.n494 B.n410 1.24928
R1339 B.n195 B.n194 1.24928
R1340 B.n215 B.n214 1.24928
R1341 B.n640 B.t7 1.23889
R1342 B.n756 B.t6 1.23889
R1343 VP.n7 VP.t1 326.909
R1344 VP.n17 VP.t3 304.048
R1345 VP.n29 VP.t7 304.048
R1346 VP.n15 VP.t0 304.048
R1347 VP.n22 VP.t5 268.759
R1348 VP.n1 VP.t6 268.759
R1349 VP.n5 VP.t4 268.759
R1350 VP.n8 VP.t2 268.759
R1351 VP.n9 VP.n6 161.3
R1352 VP.n11 VP.n10 161.3
R1353 VP.n13 VP.n12 161.3
R1354 VP.n14 VP.n4 161.3
R1355 VP.n28 VP.n0 161.3
R1356 VP.n27 VP.n26 161.3
R1357 VP.n25 VP.n24 161.3
R1358 VP.n23 VP.n2 161.3
R1359 VP.n21 VP.n20 161.3
R1360 VP.n19 VP.n3 161.3
R1361 VP.n16 VP.n15 80.6037
R1362 VP.n30 VP.n29 80.6037
R1363 VP.n18 VP.n17 80.6037
R1364 VP.n24 VP.n23 56.5193
R1365 VP.n10 VP.n9 56.5193
R1366 VP.n17 VP.n3 49.9132
R1367 VP.n29 VP.n28 49.9132
R1368 VP.n15 VP.n14 49.9132
R1369 VP.n18 VP.n16 44.5317
R1370 VP.n8 VP.n7 33.7295
R1371 VP.n7 VP.n6 28.2143
R1372 VP.n21 VP.n3 24.4675
R1373 VP.n28 VP.n27 24.4675
R1374 VP.n14 VP.n13 24.4675
R1375 VP.n23 VP.n22 23.2442
R1376 VP.n24 VP.n1 23.2442
R1377 VP.n10 VP.n5 23.2442
R1378 VP.n9 VP.n8 23.2442
R1379 VP.n22 VP.n21 1.22385
R1380 VP.n27 VP.n1 1.22385
R1381 VP.n13 VP.n5 1.22385
R1382 VP.n16 VP.n4 0.285035
R1383 VP.n19 VP.n18 0.285035
R1384 VP.n30 VP.n0 0.285035
R1385 VP.n11 VP.n6 0.189894
R1386 VP.n12 VP.n11 0.189894
R1387 VP.n12 VP.n4 0.189894
R1388 VP.n20 VP.n19 0.189894
R1389 VP.n20 VP.n2 0.189894
R1390 VP.n25 VP.n2 0.189894
R1391 VP.n26 VP.n25 0.189894
R1392 VP.n26 VP.n0 0.189894
R1393 VP VP.n30 0.146778
R1394 VTAIL.n11 VTAIL.t15 46.8879
R1395 VTAIL.n10 VTAIL.t0 46.8879
R1396 VTAIL.n7 VTAIL.t7 46.8879
R1397 VTAIL.n15 VTAIL.t5 46.8878
R1398 VTAIL.n2 VTAIL.t6 46.8878
R1399 VTAIL.n3 VTAIL.t14 46.8878
R1400 VTAIL.n6 VTAIL.t11 46.8878
R1401 VTAIL.n14 VTAIL.t9 46.8878
R1402 VTAIL.n13 VTAIL.n12 45.3027
R1403 VTAIL.n9 VTAIL.n8 45.3027
R1404 VTAIL.n1 VTAIL.n0 45.3025
R1405 VTAIL.n5 VTAIL.n4 45.3025
R1406 VTAIL.n15 VTAIL.n14 24.3841
R1407 VTAIL.n7 VTAIL.n6 24.3841
R1408 VTAIL.n0 VTAIL.t1 1.58577
R1409 VTAIL.n0 VTAIL.t4 1.58577
R1410 VTAIL.n4 VTAIL.t13 1.58577
R1411 VTAIL.n4 VTAIL.t8 1.58577
R1412 VTAIL.n12 VTAIL.t10 1.58577
R1413 VTAIL.n12 VTAIL.t12 1.58577
R1414 VTAIL.n8 VTAIL.t2 1.58577
R1415 VTAIL.n8 VTAIL.t3 1.58577
R1416 VTAIL.n9 VTAIL.n7 1.2505
R1417 VTAIL.n10 VTAIL.n9 1.2505
R1418 VTAIL.n13 VTAIL.n11 1.2505
R1419 VTAIL.n14 VTAIL.n13 1.2505
R1420 VTAIL.n6 VTAIL.n5 1.2505
R1421 VTAIL.n5 VTAIL.n3 1.2505
R1422 VTAIL.n2 VTAIL.n1 1.2505
R1423 VTAIL VTAIL.n15 1.19231
R1424 VTAIL.n11 VTAIL.n10 0.470328
R1425 VTAIL.n3 VTAIL.n2 0.470328
R1426 VTAIL VTAIL.n1 0.0586897
R1427 VDD1 VDD1.n0 62.6647
R1428 VDD1.n3 VDD1.n2 62.5509
R1429 VDD1.n3 VDD1.n1 62.5509
R1430 VDD1.n5 VDD1.n4 61.9813
R1431 VDD1.n5 VDD1.n3 40.6905
R1432 VDD1.n4 VDD1.t3 1.58577
R1433 VDD1.n4 VDD1.t7 1.58577
R1434 VDD1.n0 VDD1.t6 1.58577
R1435 VDD1.n0 VDD1.t5 1.58577
R1436 VDD1.n2 VDD1.t1 1.58577
R1437 VDD1.n2 VDD1.t0 1.58577
R1438 VDD1.n1 VDD1.t4 1.58577
R1439 VDD1.n1 VDD1.t2 1.58577
R1440 VDD1 VDD1.n5 0.56731
R1441 VN.n3 VN.t3 326.909
R1442 VN.n16 VN.t5 326.909
R1443 VN.n11 VN.t0 304.048
R1444 VN.n24 VN.t6 304.048
R1445 VN.n4 VN.t2 268.759
R1446 VN.n1 VN.t1 268.759
R1447 VN.n17 VN.t7 268.759
R1448 VN.n14 VN.t4 268.759
R1449 VN.n23 VN.n13 161.3
R1450 VN.n22 VN.n21 161.3
R1451 VN.n20 VN.n19 161.3
R1452 VN.n18 VN.n15 161.3
R1453 VN.n10 VN.n0 161.3
R1454 VN.n9 VN.n8 161.3
R1455 VN.n7 VN.n6 161.3
R1456 VN.n5 VN.n2 161.3
R1457 VN.n25 VN.n24 80.6037
R1458 VN.n12 VN.n11 80.6037
R1459 VN.n6 VN.n5 56.5193
R1460 VN.n19 VN.n18 56.5193
R1461 VN.n11 VN.n10 49.9132
R1462 VN.n24 VN.n23 49.9132
R1463 VN VN.n25 44.8172
R1464 VN.n4 VN.n3 33.7295
R1465 VN.n17 VN.n16 33.7295
R1466 VN.n16 VN.n15 28.2143
R1467 VN.n3 VN.n2 28.2143
R1468 VN.n10 VN.n9 24.4675
R1469 VN.n23 VN.n22 24.4675
R1470 VN.n5 VN.n4 23.2442
R1471 VN.n6 VN.n1 23.2442
R1472 VN.n18 VN.n17 23.2442
R1473 VN.n19 VN.n14 23.2442
R1474 VN.n9 VN.n1 1.22385
R1475 VN.n22 VN.n14 1.22385
R1476 VN.n25 VN.n13 0.285035
R1477 VN.n12 VN.n0 0.285035
R1478 VN.n21 VN.n13 0.189894
R1479 VN.n21 VN.n20 0.189894
R1480 VN.n20 VN.n15 0.189894
R1481 VN.n7 VN.n2 0.189894
R1482 VN.n8 VN.n7 0.189894
R1483 VN.n8 VN.n0 0.189894
R1484 VN VN.n12 0.146778
R1485 VDD2.n2 VDD2.n1 62.5509
R1486 VDD2.n2 VDD2.n0 62.5509
R1487 VDD2 VDD2.n5 62.5481
R1488 VDD2.n4 VDD2.n3 61.9815
R1489 VDD2.n4 VDD2.n2 40.1075
R1490 VDD2.n5 VDD2.t0 1.58577
R1491 VDD2.n5 VDD2.t2 1.58577
R1492 VDD2.n3 VDD2.t1 1.58577
R1493 VDD2.n3 VDD2.t3 1.58577
R1494 VDD2.n1 VDD2.t6 1.58577
R1495 VDD2.n1 VDD2.t7 1.58577
R1496 VDD2.n0 VDD2.t4 1.58577
R1497 VDD2.n0 VDD2.t5 1.58577
R1498 VDD2 VDD2.n4 0.68369
C0 VTAIL VN 6.97832f
C1 VTAIL VDD2 9.51304f
C2 VTAIL VDD1 9.46855f
C3 VN VP 5.94174f
C4 VP VDD2 0.362239f
C5 VP VDD1 7.29098f
C6 VTAIL VP 6.99243f
C7 VN VDD2 7.07849f
C8 VN VDD1 0.149109f
C9 VDD1 VDD2 1.03659f
C10 VDD2 B 3.93746f
C11 VDD1 B 4.216934f
C12 VTAIL B 9.616822f
C13 VN B 10.08552f
C14 VP B 8.322094f
C15 VDD2.t4 B 0.253034f
C16 VDD2.t5 B 0.253034f
C17 VDD2.n0 B 2.26345f
C18 VDD2.t6 B 0.253034f
C19 VDD2.t7 B 0.253034f
C20 VDD2.n1 B 2.26345f
C21 VDD2.n2 B 2.51339f
C22 VDD2.t1 B 0.253034f
C23 VDD2.t3 B 0.253034f
C24 VDD2.n3 B 2.26004f
C25 VDD2.n4 B 2.53883f
C26 VDD2.t0 B 0.253034f
C27 VDD2.t2 B 0.253034f
C28 VDD2.n5 B 2.26342f
C29 VN.n0 B 0.047939f
C30 VN.t1 B 1.37082f
C31 VN.n1 B 0.502523f
C32 VN.n2 B 0.188265f
C33 VN.t2 B 1.37082f
C34 VN.t3 B 1.47262f
C35 VN.n3 B 0.55043f
C36 VN.n4 B 0.560016f
C37 VN.n5 B 0.050791f
C38 VN.n6 B 0.050791f
C39 VN.n7 B 0.035926f
C40 VN.n8 B 0.035926f
C41 VN.n9 B 0.035551f
C42 VN.n10 B 0.045504f
C43 VN.t0 B 1.43247f
C44 VN.n11 B 0.565247f
C45 VN.n12 B 0.033646f
C46 VN.n13 B 0.047939f
C47 VN.t4 B 1.37082f
C48 VN.n14 B 0.502523f
C49 VN.n15 B 0.188265f
C50 VN.t7 B 1.37082f
C51 VN.t5 B 1.47262f
C52 VN.n16 B 0.55043f
C53 VN.n17 B 0.560016f
C54 VN.n18 B 0.050791f
C55 VN.n19 B 0.050791f
C56 VN.n20 B 0.035926f
C57 VN.n21 B 0.035926f
C58 VN.n22 B 0.035551f
C59 VN.n23 B 0.045504f
C60 VN.t6 B 1.43247f
C61 VN.n24 B 0.565247f
C62 VN.n25 B 1.66457f
C63 VDD1.t6 B 0.25463f
C64 VDD1.t5 B 0.25463f
C65 VDD1.n0 B 2.2785f
C66 VDD1.t4 B 0.25463f
C67 VDD1.t2 B 0.25463f
C68 VDD1.n1 B 2.27773f
C69 VDD1.t1 B 0.25463f
C70 VDD1.t0 B 0.25463f
C71 VDD1.n2 B 2.27773f
C72 VDD1.n3 B 2.58394f
C73 VDD1.t3 B 0.25463f
C74 VDD1.t7 B 0.25463f
C75 VDD1.n4 B 2.27429f
C76 VDD1.n5 B 2.58577f
C77 VTAIL.t1 B 0.189893f
C78 VTAIL.t4 B 0.189893f
C79 VTAIL.n0 B 1.63862f
C80 VTAIL.n1 B 0.272149f
C81 VTAIL.t6 B 2.09001f
C82 VTAIL.n2 B 0.364163f
C83 VTAIL.t14 B 2.09001f
C84 VTAIL.n3 B 0.364163f
C85 VTAIL.t13 B 0.189893f
C86 VTAIL.t8 B 0.189893f
C87 VTAIL.n4 B 1.63862f
C88 VTAIL.n5 B 0.346034f
C89 VTAIL.t11 B 2.09001f
C90 VTAIL.n6 B 1.34138f
C91 VTAIL.t7 B 2.09002f
C92 VTAIL.n7 B 1.34136f
C93 VTAIL.t2 B 0.189893f
C94 VTAIL.t3 B 0.189893f
C95 VTAIL.n8 B 1.63862f
C96 VTAIL.n9 B 0.346029f
C97 VTAIL.t0 B 2.09002f
C98 VTAIL.n10 B 0.36415f
C99 VTAIL.t15 B 2.09002f
C100 VTAIL.n11 B 0.36415f
C101 VTAIL.t10 B 0.189893f
C102 VTAIL.t12 B 0.189893f
C103 VTAIL.n12 B 1.63862f
C104 VTAIL.n13 B 0.346029f
C105 VTAIL.t9 B 2.09001f
C106 VTAIL.n14 B 1.34138f
C107 VTAIL.t5 B 2.09001f
C108 VTAIL.n15 B 1.33777f
C109 VP.n0 B 0.048541f
C110 VP.t6 B 1.38803f
C111 VP.n1 B 0.508833f
C112 VP.n2 B 0.036377f
C113 VP.t5 B 1.38803f
C114 VP.n3 B 0.046075f
C115 VP.n4 B 0.048541f
C116 VP.t0 B 1.45045f
C117 VP.t4 B 1.38803f
C118 VP.n5 B 0.508833f
C119 VP.n6 B 0.19063f
C120 VP.t2 B 1.38803f
C121 VP.t1 B 1.49111f
C122 VP.n7 B 0.557342f
C123 VP.n8 B 0.567048f
C124 VP.n9 B 0.051429f
C125 VP.n10 B 0.051429f
C126 VP.n11 B 0.036377f
C127 VP.n12 B 0.036377f
C128 VP.n13 B 0.035998f
C129 VP.n14 B 0.046075f
C130 VP.n15 B 0.572344f
C131 VP.n16 B 1.66526f
C132 VP.t3 B 1.45045f
C133 VP.n17 B 0.572344f
C134 VP.n18 B 1.69463f
C135 VP.n19 B 0.048541f
C136 VP.n20 B 0.036377f
C137 VP.n21 B 0.035998f
C138 VP.n22 B 0.508833f
C139 VP.n23 B 0.051429f
C140 VP.n24 B 0.051429f
C141 VP.n25 B 0.036377f
C142 VP.n26 B 0.036377f
C143 VP.n27 B 0.035998f
C144 VP.n28 B 0.046075f
C145 VP.t7 B 1.45045f
C146 VP.n29 B 0.572344f
C147 VP.n30 B 0.034068f
.ends

