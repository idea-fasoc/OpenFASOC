* NGSPICE file created from diff_pair_sample_1570.ext - technology: sky130A

.subckt diff_pair_sample_1570 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=0.89
X1 VDD1.t7 VP.t0 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=0.89
X2 VTAIL.t13 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X3 VTAIL.t14 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X4 VDD2.t7 VN.t0 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=0.89
X5 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=0.89
X6 VTAIL.t4 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X7 VTAIL.t5 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X8 VDD2.t4 VN.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X9 VDD1.t4 VP.t3 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=0.89
X10 VTAIL.t9 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=0.89
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=0.89
X12 VDD2.t3 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X13 VDD2.t2 VN.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=3.0693 ps=16.52 w=7.87 l=0.89
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=0 ps=0 w=7.87 l=0.89
X15 VTAIL.t8 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=0.89
X16 VTAIL.t0 VN.t6 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=0.89
X17 VDD1.t1 VP.t6 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X18 VDD1.t0 VP.t7 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.29855 pd=8.2 as=1.29855 ps=8.2 w=7.87 l=0.89
X19 VTAIL.t2 VN.t7 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0693 pd=16.52 as=1.29855 ps=8.2 w=7.87 l=0.89
R0 B.n430 B.n429 585
R1 B.n430 B.n50 585
R2 B.n433 B.n432 585
R3 B.n434 B.n89 585
R4 B.n436 B.n435 585
R5 B.n438 B.n88 585
R6 B.n441 B.n440 585
R7 B.n442 B.n87 585
R8 B.n444 B.n443 585
R9 B.n446 B.n86 585
R10 B.n449 B.n448 585
R11 B.n450 B.n85 585
R12 B.n452 B.n451 585
R13 B.n454 B.n84 585
R14 B.n457 B.n456 585
R15 B.n458 B.n83 585
R16 B.n460 B.n459 585
R17 B.n462 B.n82 585
R18 B.n465 B.n464 585
R19 B.n466 B.n81 585
R20 B.n468 B.n467 585
R21 B.n470 B.n80 585
R22 B.n473 B.n472 585
R23 B.n474 B.n79 585
R24 B.n476 B.n475 585
R25 B.n478 B.n78 585
R26 B.n481 B.n480 585
R27 B.n482 B.n77 585
R28 B.n484 B.n483 585
R29 B.n486 B.n76 585
R30 B.n489 B.n488 585
R31 B.n491 B.n73 585
R32 B.n493 B.n492 585
R33 B.n495 B.n72 585
R34 B.n498 B.n497 585
R35 B.n499 B.n71 585
R36 B.n501 B.n500 585
R37 B.n503 B.n70 585
R38 B.n505 B.n504 585
R39 B.n507 B.n506 585
R40 B.n510 B.n509 585
R41 B.n511 B.n65 585
R42 B.n513 B.n512 585
R43 B.n515 B.n64 585
R44 B.n518 B.n517 585
R45 B.n519 B.n63 585
R46 B.n521 B.n520 585
R47 B.n523 B.n62 585
R48 B.n526 B.n525 585
R49 B.n527 B.n61 585
R50 B.n529 B.n528 585
R51 B.n531 B.n60 585
R52 B.n534 B.n533 585
R53 B.n535 B.n59 585
R54 B.n537 B.n536 585
R55 B.n539 B.n58 585
R56 B.n542 B.n541 585
R57 B.n543 B.n57 585
R58 B.n545 B.n544 585
R59 B.n547 B.n56 585
R60 B.n550 B.n549 585
R61 B.n551 B.n55 585
R62 B.n553 B.n552 585
R63 B.n555 B.n54 585
R64 B.n558 B.n557 585
R65 B.n559 B.n53 585
R66 B.n561 B.n560 585
R67 B.n563 B.n52 585
R68 B.n566 B.n565 585
R69 B.n567 B.n51 585
R70 B.n428 B.n49 585
R71 B.n570 B.n49 585
R72 B.n427 B.n48 585
R73 B.n571 B.n48 585
R74 B.n426 B.n47 585
R75 B.n572 B.n47 585
R76 B.n425 B.n424 585
R77 B.n424 B.n43 585
R78 B.n423 B.n42 585
R79 B.n578 B.n42 585
R80 B.n422 B.n41 585
R81 B.n579 B.n41 585
R82 B.n421 B.n40 585
R83 B.n580 B.n40 585
R84 B.n420 B.n419 585
R85 B.n419 B.n36 585
R86 B.n418 B.n35 585
R87 B.n586 B.n35 585
R88 B.n417 B.n34 585
R89 B.n587 B.n34 585
R90 B.n416 B.n33 585
R91 B.n588 B.n33 585
R92 B.n415 B.n414 585
R93 B.n414 B.n32 585
R94 B.n413 B.n28 585
R95 B.n594 B.n28 585
R96 B.n412 B.n27 585
R97 B.n595 B.n27 585
R98 B.n411 B.n26 585
R99 B.n596 B.n26 585
R100 B.n410 B.n409 585
R101 B.n409 B.n25 585
R102 B.n408 B.n21 585
R103 B.n602 B.n21 585
R104 B.n407 B.n20 585
R105 B.n603 B.n20 585
R106 B.n406 B.n19 585
R107 B.n604 B.n19 585
R108 B.n405 B.n404 585
R109 B.n404 B.n18 585
R110 B.n403 B.n14 585
R111 B.n610 B.n14 585
R112 B.n402 B.n13 585
R113 B.n611 B.n13 585
R114 B.n401 B.n12 585
R115 B.n612 B.n12 585
R116 B.n400 B.n399 585
R117 B.n399 B.n8 585
R118 B.n398 B.n7 585
R119 B.n618 B.n7 585
R120 B.n397 B.n6 585
R121 B.n619 B.n6 585
R122 B.n396 B.n5 585
R123 B.n620 B.n5 585
R124 B.n395 B.n394 585
R125 B.n394 B.n4 585
R126 B.n393 B.n90 585
R127 B.n393 B.n392 585
R128 B.n383 B.n91 585
R129 B.n92 B.n91 585
R130 B.n385 B.n384 585
R131 B.n386 B.n385 585
R132 B.n382 B.n97 585
R133 B.n97 B.n96 585
R134 B.n381 B.n380 585
R135 B.n380 B.n379 585
R136 B.n99 B.n98 585
R137 B.n372 B.n99 585
R138 B.n371 B.n370 585
R139 B.n373 B.n371 585
R140 B.n369 B.n104 585
R141 B.n104 B.n103 585
R142 B.n368 B.n367 585
R143 B.n367 B.n366 585
R144 B.n106 B.n105 585
R145 B.n359 B.n106 585
R146 B.n358 B.n357 585
R147 B.n360 B.n358 585
R148 B.n356 B.n111 585
R149 B.n111 B.n110 585
R150 B.n355 B.n354 585
R151 B.n354 B.n353 585
R152 B.n113 B.n112 585
R153 B.n346 B.n113 585
R154 B.n345 B.n344 585
R155 B.n347 B.n345 585
R156 B.n343 B.n118 585
R157 B.n118 B.n117 585
R158 B.n342 B.n341 585
R159 B.n341 B.n340 585
R160 B.n120 B.n119 585
R161 B.n121 B.n120 585
R162 B.n333 B.n332 585
R163 B.n334 B.n333 585
R164 B.n331 B.n125 585
R165 B.n129 B.n125 585
R166 B.n330 B.n329 585
R167 B.n329 B.n328 585
R168 B.n127 B.n126 585
R169 B.n128 B.n127 585
R170 B.n321 B.n320 585
R171 B.n322 B.n321 585
R172 B.n319 B.n134 585
R173 B.n134 B.n133 585
R174 B.n318 B.n317 585
R175 B.n317 B.n316 585
R176 B.n313 B.n138 585
R177 B.n312 B.n311 585
R178 B.n309 B.n139 585
R179 B.n309 B.n137 585
R180 B.n308 B.n307 585
R181 B.n306 B.n305 585
R182 B.n304 B.n141 585
R183 B.n302 B.n301 585
R184 B.n300 B.n142 585
R185 B.n299 B.n298 585
R186 B.n296 B.n143 585
R187 B.n294 B.n293 585
R188 B.n292 B.n144 585
R189 B.n291 B.n290 585
R190 B.n288 B.n145 585
R191 B.n286 B.n285 585
R192 B.n284 B.n146 585
R193 B.n283 B.n282 585
R194 B.n280 B.n147 585
R195 B.n278 B.n277 585
R196 B.n276 B.n148 585
R197 B.n275 B.n274 585
R198 B.n272 B.n149 585
R199 B.n270 B.n269 585
R200 B.n268 B.n150 585
R201 B.n267 B.n266 585
R202 B.n264 B.n151 585
R203 B.n262 B.n261 585
R204 B.n260 B.n152 585
R205 B.n259 B.n258 585
R206 B.n256 B.n153 585
R207 B.n254 B.n253 585
R208 B.n252 B.n154 585
R209 B.n251 B.n250 585
R210 B.n248 B.n158 585
R211 B.n246 B.n245 585
R212 B.n244 B.n159 585
R213 B.n243 B.n242 585
R214 B.n240 B.n160 585
R215 B.n238 B.n237 585
R216 B.n235 B.n161 585
R217 B.n234 B.n233 585
R218 B.n231 B.n164 585
R219 B.n229 B.n228 585
R220 B.n227 B.n165 585
R221 B.n226 B.n225 585
R222 B.n223 B.n166 585
R223 B.n221 B.n220 585
R224 B.n219 B.n167 585
R225 B.n218 B.n217 585
R226 B.n215 B.n168 585
R227 B.n213 B.n212 585
R228 B.n211 B.n169 585
R229 B.n210 B.n209 585
R230 B.n207 B.n170 585
R231 B.n205 B.n204 585
R232 B.n203 B.n171 585
R233 B.n202 B.n201 585
R234 B.n199 B.n172 585
R235 B.n197 B.n196 585
R236 B.n195 B.n173 585
R237 B.n194 B.n193 585
R238 B.n191 B.n174 585
R239 B.n189 B.n188 585
R240 B.n187 B.n175 585
R241 B.n186 B.n185 585
R242 B.n183 B.n176 585
R243 B.n181 B.n180 585
R244 B.n179 B.n178 585
R245 B.n136 B.n135 585
R246 B.n315 B.n314 585
R247 B.n316 B.n315 585
R248 B.n132 B.n131 585
R249 B.n133 B.n132 585
R250 B.n324 B.n323 585
R251 B.n323 B.n322 585
R252 B.n325 B.n130 585
R253 B.n130 B.n128 585
R254 B.n327 B.n326 585
R255 B.n328 B.n327 585
R256 B.n124 B.n123 585
R257 B.n129 B.n124 585
R258 B.n336 B.n335 585
R259 B.n335 B.n334 585
R260 B.n337 B.n122 585
R261 B.n122 B.n121 585
R262 B.n339 B.n338 585
R263 B.n340 B.n339 585
R264 B.n116 B.n115 585
R265 B.n117 B.n116 585
R266 B.n349 B.n348 585
R267 B.n348 B.n347 585
R268 B.n350 B.n114 585
R269 B.n346 B.n114 585
R270 B.n352 B.n351 585
R271 B.n353 B.n352 585
R272 B.n109 B.n108 585
R273 B.n110 B.n109 585
R274 B.n362 B.n361 585
R275 B.n361 B.n360 585
R276 B.n363 B.n107 585
R277 B.n359 B.n107 585
R278 B.n365 B.n364 585
R279 B.n366 B.n365 585
R280 B.n102 B.n101 585
R281 B.n103 B.n102 585
R282 B.n375 B.n374 585
R283 B.n374 B.n373 585
R284 B.n376 B.n100 585
R285 B.n372 B.n100 585
R286 B.n378 B.n377 585
R287 B.n379 B.n378 585
R288 B.n95 B.n94 585
R289 B.n96 B.n95 585
R290 B.n388 B.n387 585
R291 B.n387 B.n386 585
R292 B.n389 B.n93 585
R293 B.n93 B.n92 585
R294 B.n391 B.n390 585
R295 B.n392 B.n391 585
R296 B.n2 B.n0 585
R297 B.n4 B.n2 585
R298 B.n3 B.n1 585
R299 B.n619 B.n3 585
R300 B.n617 B.n616 585
R301 B.n618 B.n617 585
R302 B.n615 B.n9 585
R303 B.n9 B.n8 585
R304 B.n614 B.n613 585
R305 B.n613 B.n612 585
R306 B.n11 B.n10 585
R307 B.n611 B.n11 585
R308 B.n609 B.n608 585
R309 B.n610 B.n609 585
R310 B.n607 B.n15 585
R311 B.n18 B.n15 585
R312 B.n606 B.n605 585
R313 B.n605 B.n604 585
R314 B.n17 B.n16 585
R315 B.n603 B.n17 585
R316 B.n601 B.n600 585
R317 B.n602 B.n601 585
R318 B.n599 B.n22 585
R319 B.n25 B.n22 585
R320 B.n598 B.n597 585
R321 B.n597 B.n596 585
R322 B.n24 B.n23 585
R323 B.n595 B.n24 585
R324 B.n593 B.n592 585
R325 B.n594 B.n593 585
R326 B.n591 B.n29 585
R327 B.n32 B.n29 585
R328 B.n590 B.n589 585
R329 B.n589 B.n588 585
R330 B.n31 B.n30 585
R331 B.n587 B.n31 585
R332 B.n585 B.n584 585
R333 B.n586 B.n585 585
R334 B.n583 B.n37 585
R335 B.n37 B.n36 585
R336 B.n582 B.n581 585
R337 B.n581 B.n580 585
R338 B.n39 B.n38 585
R339 B.n579 B.n39 585
R340 B.n577 B.n576 585
R341 B.n578 B.n577 585
R342 B.n575 B.n44 585
R343 B.n44 B.n43 585
R344 B.n574 B.n573 585
R345 B.n573 B.n572 585
R346 B.n46 B.n45 585
R347 B.n571 B.n46 585
R348 B.n569 B.n568 585
R349 B.n570 B.n569 585
R350 B.n622 B.n621 585
R351 B.n621 B.n620 585
R352 B.n315 B.n138 473.281
R353 B.n569 B.n51 473.281
R354 B.n317 B.n136 473.281
R355 B.n430 B.n49 473.281
R356 B.n162 B.t16 415.87
R357 B.n74 B.t12 415.87
R358 B.n155 B.t8 415.264
R359 B.n66 B.t19 415.264
R360 B.n431 B.n50 256.663
R361 B.n437 B.n50 256.663
R362 B.n439 B.n50 256.663
R363 B.n445 B.n50 256.663
R364 B.n447 B.n50 256.663
R365 B.n453 B.n50 256.663
R366 B.n455 B.n50 256.663
R367 B.n461 B.n50 256.663
R368 B.n463 B.n50 256.663
R369 B.n469 B.n50 256.663
R370 B.n471 B.n50 256.663
R371 B.n477 B.n50 256.663
R372 B.n479 B.n50 256.663
R373 B.n485 B.n50 256.663
R374 B.n487 B.n50 256.663
R375 B.n494 B.n50 256.663
R376 B.n496 B.n50 256.663
R377 B.n502 B.n50 256.663
R378 B.n69 B.n50 256.663
R379 B.n508 B.n50 256.663
R380 B.n514 B.n50 256.663
R381 B.n516 B.n50 256.663
R382 B.n522 B.n50 256.663
R383 B.n524 B.n50 256.663
R384 B.n530 B.n50 256.663
R385 B.n532 B.n50 256.663
R386 B.n538 B.n50 256.663
R387 B.n540 B.n50 256.663
R388 B.n546 B.n50 256.663
R389 B.n548 B.n50 256.663
R390 B.n554 B.n50 256.663
R391 B.n556 B.n50 256.663
R392 B.n562 B.n50 256.663
R393 B.n564 B.n50 256.663
R394 B.n310 B.n137 256.663
R395 B.n140 B.n137 256.663
R396 B.n303 B.n137 256.663
R397 B.n297 B.n137 256.663
R398 B.n295 B.n137 256.663
R399 B.n289 B.n137 256.663
R400 B.n287 B.n137 256.663
R401 B.n281 B.n137 256.663
R402 B.n279 B.n137 256.663
R403 B.n273 B.n137 256.663
R404 B.n271 B.n137 256.663
R405 B.n265 B.n137 256.663
R406 B.n263 B.n137 256.663
R407 B.n257 B.n137 256.663
R408 B.n255 B.n137 256.663
R409 B.n249 B.n137 256.663
R410 B.n247 B.n137 256.663
R411 B.n241 B.n137 256.663
R412 B.n239 B.n137 256.663
R413 B.n232 B.n137 256.663
R414 B.n230 B.n137 256.663
R415 B.n224 B.n137 256.663
R416 B.n222 B.n137 256.663
R417 B.n216 B.n137 256.663
R418 B.n214 B.n137 256.663
R419 B.n208 B.n137 256.663
R420 B.n206 B.n137 256.663
R421 B.n200 B.n137 256.663
R422 B.n198 B.n137 256.663
R423 B.n192 B.n137 256.663
R424 B.n190 B.n137 256.663
R425 B.n184 B.n137 256.663
R426 B.n182 B.n137 256.663
R427 B.n177 B.n137 256.663
R428 B.n162 B.t18 234.625
R429 B.n74 B.t14 234.625
R430 B.n155 B.t11 234.625
R431 B.n66 B.t20 234.625
R432 B.n163 B.t17 210.964
R433 B.n75 B.t15 210.964
R434 B.n156 B.t10 210.964
R435 B.n67 B.t21 210.964
R436 B.n315 B.n132 163.367
R437 B.n323 B.n132 163.367
R438 B.n323 B.n130 163.367
R439 B.n327 B.n130 163.367
R440 B.n327 B.n124 163.367
R441 B.n335 B.n124 163.367
R442 B.n335 B.n122 163.367
R443 B.n339 B.n122 163.367
R444 B.n339 B.n116 163.367
R445 B.n348 B.n116 163.367
R446 B.n348 B.n114 163.367
R447 B.n352 B.n114 163.367
R448 B.n352 B.n109 163.367
R449 B.n361 B.n109 163.367
R450 B.n361 B.n107 163.367
R451 B.n365 B.n107 163.367
R452 B.n365 B.n102 163.367
R453 B.n374 B.n102 163.367
R454 B.n374 B.n100 163.367
R455 B.n378 B.n100 163.367
R456 B.n378 B.n95 163.367
R457 B.n387 B.n95 163.367
R458 B.n387 B.n93 163.367
R459 B.n391 B.n93 163.367
R460 B.n391 B.n2 163.367
R461 B.n621 B.n2 163.367
R462 B.n621 B.n3 163.367
R463 B.n617 B.n3 163.367
R464 B.n617 B.n9 163.367
R465 B.n613 B.n9 163.367
R466 B.n613 B.n11 163.367
R467 B.n609 B.n11 163.367
R468 B.n609 B.n15 163.367
R469 B.n605 B.n15 163.367
R470 B.n605 B.n17 163.367
R471 B.n601 B.n17 163.367
R472 B.n601 B.n22 163.367
R473 B.n597 B.n22 163.367
R474 B.n597 B.n24 163.367
R475 B.n593 B.n24 163.367
R476 B.n593 B.n29 163.367
R477 B.n589 B.n29 163.367
R478 B.n589 B.n31 163.367
R479 B.n585 B.n31 163.367
R480 B.n585 B.n37 163.367
R481 B.n581 B.n37 163.367
R482 B.n581 B.n39 163.367
R483 B.n577 B.n39 163.367
R484 B.n577 B.n44 163.367
R485 B.n573 B.n44 163.367
R486 B.n573 B.n46 163.367
R487 B.n569 B.n46 163.367
R488 B.n311 B.n309 163.367
R489 B.n309 B.n308 163.367
R490 B.n305 B.n304 163.367
R491 B.n302 B.n142 163.367
R492 B.n298 B.n296 163.367
R493 B.n294 B.n144 163.367
R494 B.n290 B.n288 163.367
R495 B.n286 B.n146 163.367
R496 B.n282 B.n280 163.367
R497 B.n278 B.n148 163.367
R498 B.n274 B.n272 163.367
R499 B.n270 B.n150 163.367
R500 B.n266 B.n264 163.367
R501 B.n262 B.n152 163.367
R502 B.n258 B.n256 163.367
R503 B.n254 B.n154 163.367
R504 B.n250 B.n248 163.367
R505 B.n246 B.n159 163.367
R506 B.n242 B.n240 163.367
R507 B.n238 B.n161 163.367
R508 B.n233 B.n231 163.367
R509 B.n229 B.n165 163.367
R510 B.n225 B.n223 163.367
R511 B.n221 B.n167 163.367
R512 B.n217 B.n215 163.367
R513 B.n213 B.n169 163.367
R514 B.n209 B.n207 163.367
R515 B.n205 B.n171 163.367
R516 B.n201 B.n199 163.367
R517 B.n197 B.n173 163.367
R518 B.n193 B.n191 163.367
R519 B.n189 B.n175 163.367
R520 B.n185 B.n183 163.367
R521 B.n181 B.n178 163.367
R522 B.n317 B.n134 163.367
R523 B.n321 B.n134 163.367
R524 B.n321 B.n127 163.367
R525 B.n329 B.n127 163.367
R526 B.n329 B.n125 163.367
R527 B.n333 B.n125 163.367
R528 B.n333 B.n120 163.367
R529 B.n341 B.n120 163.367
R530 B.n341 B.n118 163.367
R531 B.n345 B.n118 163.367
R532 B.n345 B.n113 163.367
R533 B.n354 B.n113 163.367
R534 B.n354 B.n111 163.367
R535 B.n358 B.n111 163.367
R536 B.n358 B.n106 163.367
R537 B.n367 B.n106 163.367
R538 B.n367 B.n104 163.367
R539 B.n371 B.n104 163.367
R540 B.n371 B.n99 163.367
R541 B.n380 B.n99 163.367
R542 B.n380 B.n97 163.367
R543 B.n385 B.n97 163.367
R544 B.n385 B.n91 163.367
R545 B.n393 B.n91 163.367
R546 B.n394 B.n393 163.367
R547 B.n394 B.n5 163.367
R548 B.n6 B.n5 163.367
R549 B.n7 B.n6 163.367
R550 B.n399 B.n7 163.367
R551 B.n399 B.n12 163.367
R552 B.n13 B.n12 163.367
R553 B.n14 B.n13 163.367
R554 B.n404 B.n14 163.367
R555 B.n404 B.n19 163.367
R556 B.n20 B.n19 163.367
R557 B.n21 B.n20 163.367
R558 B.n409 B.n21 163.367
R559 B.n409 B.n26 163.367
R560 B.n27 B.n26 163.367
R561 B.n28 B.n27 163.367
R562 B.n414 B.n28 163.367
R563 B.n414 B.n33 163.367
R564 B.n34 B.n33 163.367
R565 B.n35 B.n34 163.367
R566 B.n419 B.n35 163.367
R567 B.n419 B.n40 163.367
R568 B.n41 B.n40 163.367
R569 B.n42 B.n41 163.367
R570 B.n424 B.n42 163.367
R571 B.n424 B.n47 163.367
R572 B.n48 B.n47 163.367
R573 B.n49 B.n48 163.367
R574 B.n565 B.n563 163.367
R575 B.n561 B.n53 163.367
R576 B.n557 B.n555 163.367
R577 B.n553 B.n55 163.367
R578 B.n549 B.n547 163.367
R579 B.n545 B.n57 163.367
R580 B.n541 B.n539 163.367
R581 B.n537 B.n59 163.367
R582 B.n533 B.n531 163.367
R583 B.n529 B.n61 163.367
R584 B.n525 B.n523 163.367
R585 B.n521 B.n63 163.367
R586 B.n517 B.n515 163.367
R587 B.n513 B.n65 163.367
R588 B.n509 B.n507 163.367
R589 B.n504 B.n503 163.367
R590 B.n501 B.n71 163.367
R591 B.n497 B.n495 163.367
R592 B.n493 B.n73 163.367
R593 B.n488 B.n486 163.367
R594 B.n484 B.n77 163.367
R595 B.n480 B.n478 163.367
R596 B.n476 B.n79 163.367
R597 B.n472 B.n470 163.367
R598 B.n468 B.n81 163.367
R599 B.n464 B.n462 163.367
R600 B.n460 B.n83 163.367
R601 B.n456 B.n454 163.367
R602 B.n452 B.n85 163.367
R603 B.n448 B.n446 163.367
R604 B.n444 B.n87 163.367
R605 B.n440 B.n438 163.367
R606 B.n436 B.n89 163.367
R607 B.n432 B.n430 163.367
R608 B.n316 B.n137 106.195
R609 B.n570 B.n50 106.195
R610 B.n310 B.n138 71.676
R611 B.n308 B.n140 71.676
R612 B.n304 B.n303 71.676
R613 B.n297 B.n142 71.676
R614 B.n296 B.n295 71.676
R615 B.n289 B.n144 71.676
R616 B.n288 B.n287 71.676
R617 B.n281 B.n146 71.676
R618 B.n280 B.n279 71.676
R619 B.n273 B.n148 71.676
R620 B.n272 B.n271 71.676
R621 B.n265 B.n150 71.676
R622 B.n264 B.n263 71.676
R623 B.n257 B.n152 71.676
R624 B.n256 B.n255 71.676
R625 B.n249 B.n154 71.676
R626 B.n248 B.n247 71.676
R627 B.n241 B.n159 71.676
R628 B.n240 B.n239 71.676
R629 B.n232 B.n161 71.676
R630 B.n231 B.n230 71.676
R631 B.n224 B.n165 71.676
R632 B.n223 B.n222 71.676
R633 B.n216 B.n167 71.676
R634 B.n215 B.n214 71.676
R635 B.n208 B.n169 71.676
R636 B.n207 B.n206 71.676
R637 B.n200 B.n171 71.676
R638 B.n199 B.n198 71.676
R639 B.n192 B.n173 71.676
R640 B.n191 B.n190 71.676
R641 B.n184 B.n175 71.676
R642 B.n183 B.n182 71.676
R643 B.n178 B.n177 71.676
R644 B.n564 B.n51 71.676
R645 B.n563 B.n562 71.676
R646 B.n556 B.n53 71.676
R647 B.n555 B.n554 71.676
R648 B.n548 B.n55 71.676
R649 B.n547 B.n546 71.676
R650 B.n540 B.n57 71.676
R651 B.n539 B.n538 71.676
R652 B.n532 B.n59 71.676
R653 B.n531 B.n530 71.676
R654 B.n524 B.n61 71.676
R655 B.n523 B.n522 71.676
R656 B.n516 B.n63 71.676
R657 B.n515 B.n514 71.676
R658 B.n508 B.n65 71.676
R659 B.n507 B.n69 71.676
R660 B.n503 B.n502 71.676
R661 B.n496 B.n71 71.676
R662 B.n495 B.n494 71.676
R663 B.n487 B.n73 71.676
R664 B.n486 B.n485 71.676
R665 B.n479 B.n77 71.676
R666 B.n478 B.n477 71.676
R667 B.n471 B.n79 71.676
R668 B.n470 B.n469 71.676
R669 B.n463 B.n81 71.676
R670 B.n462 B.n461 71.676
R671 B.n455 B.n83 71.676
R672 B.n454 B.n453 71.676
R673 B.n447 B.n85 71.676
R674 B.n446 B.n445 71.676
R675 B.n439 B.n87 71.676
R676 B.n438 B.n437 71.676
R677 B.n431 B.n89 71.676
R678 B.n432 B.n431 71.676
R679 B.n437 B.n436 71.676
R680 B.n440 B.n439 71.676
R681 B.n445 B.n444 71.676
R682 B.n448 B.n447 71.676
R683 B.n453 B.n452 71.676
R684 B.n456 B.n455 71.676
R685 B.n461 B.n460 71.676
R686 B.n464 B.n463 71.676
R687 B.n469 B.n468 71.676
R688 B.n472 B.n471 71.676
R689 B.n477 B.n476 71.676
R690 B.n480 B.n479 71.676
R691 B.n485 B.n484 71.676
R692 B.n488 B.n487 71.676
R693 B.n494 B.n493 71.676
R694 B.n497 B.n496 71.676
R695 B.n502 B.n501 71.676
R696 B.n504 B.n69 71.676
R697 B.n509 B.n508 71.676
R698 B.n514 B.n513 71.676
R699 B.n517 B.n516 71.676
R700 B.n522 B.n521 71.676
R701 B.n525 B.n524 71.676
R702 B.n530 B.n529 71.676
R703 B.n533 B.n532 71.676
R704 B.n538 B.n537 71.676
R705 B.n541 B.n540 71.676
R706 B.n546 B.n545 71.676
R707 B.n549 B.n548 71.676
R708 B.n554 B.n553 71.676
R709 B.n557 B.n556 71.676
R710 B.n562 B.n561 71.676
R711 B.n565 B.n564 71.676
R712 B.n311 B.n310 71.676
R713 B.n305 B.n140 71.676
R714 B.n303 B.n302 71.676
R715 B.n298 B.n297 71.676
R716 B.n295 B.n294 71.676
R717 B.n290 B.n289 71.676
R718 B.n287 B.n286 71.676
R719 B.n282 B.n281 71.676
R720 B.n279 B.n278 71.676
R721 B.n274 B.n273 71.676
R722 B.n271 B.n270 71.676
R723 B.n266 B.n265 71.676
R724 B.n263 B.n262 71.676
R725 B.n258 B.n257 71.676
R726 B.n255 B.n254 71.676
R727 B.n250 B.n249 71.676
R728 B.n247 B.n246 71.676
R729 B.n242 B.n241 71.676
R730 B.n239 B.n238 71.676
R731 B.n233 B.n232 71.676
R732 B.n230 B.n229 71.676
R733 B.n225 B.n224 71.676
R734 B.n222 B.n221 71.676
R735 B.n217 B.n216 71.676
R736 B.n214 B.n213 71.676
R737 B.n209 B.n208 71.676
R738 B.n206 B.n205 71.676
R739 B.n201 B.n200 71.676
R740 B.n198 B.n197 71.676
R741 B.n193 B.n192 71.676
R742 B.n190 B.n189 71.676
R743 B.n185 B.n184 71.676
R744 B.n182 B.n181 71.676
R745 B.n177 B.n136 71.676
R746 B.n236 B.n163 59.5399
R747 B.n157 B.n156 59.5399
R748 B.n68 B.n67 59.5399
R749 B.n490 B.n75 59.5399
R750 B.n316 B.n133 56.861
R751 B.n322 B.n133 56.861
R752 B.n322 B.n128 56.861
R753 B.n328 B.n128 56.861
R754 B.n328 B.n129 56.861
R755 B.n334 B.n121 56.861
R756 B.n340 B.n121 56.861
R757 B.n340 B.n117 56.861
R758 B.n347 B.n117 56.861
R759 B.n347 B.n346 56.861
R760 B.n353 B.n110 56.861
R761 B.n360 B.n110 56.861
R762 B.n360 B.n359 56.861
R763 B.n366 B.n103 56.861
R764 B.n373 B.n103 56.861
R765 B.n373 B.n372 56.861
R766 B.n379 B.n96 56.861
R767 B.n386 B.n96 56.861
R768 B.n392 B.n92 56.861
R769 B.n392 B.n4 56.861
R770 B.n620 B.n4 56.861
R771 B.n620 B.n619 56.861
R772 B.n619 B.n618 56.861
R773 B.n618 B.n8 56.861
R774 B.n612 B.n611 56.861
R775 B.n611 B.n610 56.861
R776 B.n604 B.n18 56.861
R777 B.n604 B.n603 56.861
R778 B.n603 B.n602 56.861
R779 B.n596 B.n25 56.861
R780 B.n596 B.n595 56.861
R781 B.n595 B.n594 56.861
R782 B.n588 B.n32 56.861
R783 B.n588 B.n587 56.861
R784 B.n587 B.n586 56.861
R785 B.n586 B.n36 56.861
R786 B.n580 B.n36 56.861
R787 B.n579 B.n578 56.861
R788 B.n578 B.n43 56.861
R789 B.n572 B.n43 56.861
R790 B.n572 B.n571 56.861
R791 B.n571 B.n570 56.861
R792 B.n379 B.t6 56.0248
R793 B.n610 B.t0 56.0248
R794 B.n334 B.t9 54.3525
R795 B.n580 B.t13 54.3525
R796 B.n346 B.t1 47.663
R797 B.n32 B.t4 47.663
R798 B.n386 B.t5 34.284
R799 B.n612 B.t2 34.284
R800 B.n366 B.t7 32.6117
R801 B.n602 B.t3 32.6117
R802 B.n429 B.n428 30.7517
R803 B.n568 B.n567 30.7517
R804 B.n318 B.n135 30.7517
R805 B.n314 B.n313 30.7517
R806 B.n359 B.t7 24.2498
R807 B.n25 B.t3 24.2498
R808 B.n163 B.n162 23.6611
R809 B.n156 B.n155 23.6611
R810 B.n67 B.n66 23.6611
R811 B.n75 B.n74 23.6611
R812 B.t5 B.n92 22.5775
R813 B.t2 B.n8 22.5775
R814 B B.n622 18.0485
R815 B.n567 B.n566 10.6151
R816 B.n566 B.n52 10.6151
R817 B.n560 B.n52 10.6151
R818 B.n560 B.n559 10.6151
R819 B.n559 B.n558 10.6151
R820 B.n558 B.n54 10.6151
R821 B.n552 B.n54 10.6151
R822 B.n552 B.n551 10.6151
R823 B.n551 B.n550 10.6151
R824 B.n550 B.n56 10.6151
R825 B.n544 B.n56 10.6151
R826 B.n544 B.n543 10.6151
R827 B.n543 B.n542 10.6151
R828 B.n542 B.n58 10.6151
R829 B.n536 B.n58 10.6151
R830 B.n536 B.n535 10.6151
R831 B.n535 B.n534 10.6151
R832 B.n534 B.n60 10.6151
R833 B.n528 B.n60 10.6151
R834 B.n528 B.n527 10.6151
R835 B.n527 B.n526 10.6151
R836 B.n526 B.n62 10.6151
R837 B.n520 B.n62 10.6151
R838 B.n520 B.n519 10.6151
R839 B.n519 B.n518 10.6151
R840 B.n518 B.n64 10.6151
R841 B.n512 B.n64 10.6151
R842 B.n512 B.n511 10.6151
R843 B.n511 B.n510 10.6151
R844 B.n506 B.n505 10.6151
R845 B.n505 B.n70 10.6151
R846 B.n500 B.n70 10.6151
R847 B.n500 B.n499 10.6151
R848 B.n499 B.n498 10.6151
R849 B.n498 B.n72 10.6151
R850 B.n492 B.n72 10.6151
R851 B.n492 B.n491 10.6151
R852 B.n489 B.n76 10.6151
R853 B.n483 B.n76 10.6151
R854 B.n483 B.n482 10.6151
R855 B.n482 B.n481 10.6151
R856 B.n481 B.n78 10.6151
R857 B.n475 B.n78 10.6151
R858 B.n475 B.n474 10.6151
R859 B.n474 B.n473 10.6151
R860 B.n473 B.n80 10.6151
R861 B.n467 B.n80 10.6151
R862 B.n467 B.n466 10.6151
R863 B.n466 B.n465 10.6151
R864 B.n465 B.n82 10.6151
R865 B.n459 B.n82 10.6151
R866 B.n459 B.n458 10.6151
R867 B.n458 B.n457 10.6151
R868 B.n457 B.n84 10.6151
R869 B.n451 B.n84 10.6151
R870 B.n451 B.n450 10.6151
R871 B.n450 B.n449 10.6151
R872 B.n449 B.n86 10.6151
R873 B.n443 B.n86 10.6151
R874 B.n443 B.n442 10.6151
R875 B.n442 B.n441 10.6151
R876 B.n441 B.n88 10.6151
R877 B.n435 B.n88 10.6151
R878 B.n435 B.n434 10.6151
R879 B.n434 B.n433 10.6151
R880 B.n433 B.n429 10.6151
R881 B.n319 B.n318 10.6151
R882 B.n320 B.n319 10.6151
R883 B.n320 B.n126 10.6151
R884 B.n330 B.n126 10.6151
R885 B.n331 B.n330 10.6151
R886 B.n332 B.n331 10.6151
R887 B.n332 B.n119 10.6151
R888 B.n342 B.n119 10.6151
R889 B.n343 B.n342 10.6151
R890 B.n344 B.n343 10.6151
R891 B.n344 B.n112 10.6151
R892 B.n355 B.n112 10.6151
R893 B.n356 B.n355 10.6151
R894 B.n357 B.n356 10.6151
R895 B.n357 B.n105 10.6151
R896 B.n368 B.n105 10.6151
R897 B.n369 B.n368 10.6151
R898 B.n370 B.n369 10.6151
R899 B.n370 B.n98 10.6151
R900 B.n381 B.n98 10.6151
R901 B.n382 B.n381 10.6151
R902 B.n384 B.n382 10.6151
R903 B.n384 B.n383 10.6151
R904 B.n383 B.n90 10.6151
R905 B.n395 B.n90 10.6151
R906 B.n396 B.n395 10.6151
R907 B.n397 B.n396 10.6151
R908 B.n398 B.n397 10.6151
R909 B.n400 B.n398 10.6151
R910 B.n401 B.n400 10.6151
R911 B.n402 B.n401 10.6151
R912 B.n403 B.n402 10.6151
R913 B.n405 B.n403 10.6151
R914 B.n406 B.n405 10.6151
R915 B.n407 B.n406 10.6151
R916 B.n408 B.n407 10.6151
R917 B.n410 B.n408 10.6151
R918 B.n411 B.n410 10.6151
R919 B.n412 B.n411 10.6151
R920 B.n413 B.n412 10.6151
R921 B.n415 B.n413 10.6151
R922 B.n416 B.n415 10.6151
R923 B.n417 B.n416 10.6151
R924 B.n418 B.n417 10.6151
R925 B.n420 B.n418 10.6151
R926 B.n421 B.n420 10.6151
R927 B.n422 B.n421 10.6151
R928 B.n423 B.n422 10.6151
R929 B.n425 B.n423 10.6151
R930 B.n426 B.n425 10.6151
R931 B.n427 B.n426 10.6151
R932 B.n428 B.n427 10.6151
R933 B.n313 B.n312 10.6151
R934 B.n312 B.n139 10.6151
R935 B.n307 B.n139 10.6151
R936 B.n307 B.n306 10.6151
R937 B.n306 B.n141 10.6151
R938 B.n301 B.n141 10.6151
R939 B.n301 B.n300 10.6151
R940 B.n300 B.n299 10.6151
R941 B.n299 B.n143 10.6151
R942 B.n293 B.n143 10.6151
R943 B.n293 B.n292 10.6151
R944 B.n292 B.n291 10.6151
R945 B.n291 B.n145 10.6151
R946 B.n285 B.n145 10.6151
R947 B.n285 B.n284 10.6151
R948 B.n284 B.n283 10.6151
R949 B.n283 B.n147 10.6151
R950 B.n277 B.n147 10.6151
R951 B.n277 B.n276 10.6151
R952 B.n276 B.n275 10.6151
R953 B.n275 B.n149 10.6151
R954 B.n269 B.n149 10.6151
R955 B.n269 B.n268 10.6151
R956 B.n268 B.n267 10.6151
R957 B.n267 B.n151 10.6151
R958 B.n261 B.n151 10.6151
R959 B.n261 B.n260 10.6151
R960 B.n260 B.n259 10.6151
R961 B.n259 B.n153 10.6151
R962 B.n253 B.n252 10.6151
R963 B.n252 B.n251 10.6151
R964 B.n251 B.n158 10.6151
R965 B.n245 B.n158 10.6151
R966 B.n245 B.n244 10.6151
R967 B.n244 B.n243 10.6151
R968 B.n243 B.n160 10.6151
R969 B.n237 B.n160 10.6151
R970 B.n235 B.n234 10.6151
R971 B.n234 B.n164 10.6151
R972 B.n228 B.n164 10.6151
R973 B.n228 B.n227 10.6151
R974 B.n227 B.n226 10.6151
R975 B.n226 B.n166 10.6151
R976 B.n220 B.n166 10.6151
R977 B.n220 B.n219 10.6151
R978 B.n219 B.n218 10.6151
R979 B.n218 B.n168 10.6151
R980 B.n212 B.n168 10.6151
R981 B.n212 B.n211 10.6151
R982 B.n211 B.n210 10.6151
R983 B.n210 B.n170 10.6151
R984 B.n204 B.n170 10.6151
R985 B.n204 B.n203 10.6151
R986 B.n203 B.n202 10.6151
R987 B.n202 B.n172 10.6151
R988 B.n196 B.n172 10.6151
R989 B.n196 B.n195 10.6151
R990 B.n195 B.n194 10.6151
R991 B.n194 B.n174 10.6151
R992 B.n188 B.n174 10.6151
R993 B.n188 B.n187 10.6151
R994 B.n187 B.n186 10.6151
R995 B.n186 B.n176 10.6151
R996 B.n180 B.n176 10.6151
R997 B.n180 B.n179 10.6151
R998 B.n179 B.n135 10.6151
R999 B.n314 B.n131 10.6151
R1000 B.n324 B.n131 10.6151
R1001 B.n325 B.n324 10.6151
R1002 B.n326 B.n325 10.6151
R1003 B.n326 B.n123 10.6151
R1004 B.n336 B.n123 10.6151
R1005 B.n337 B.n336 10.6151
R1006 B.n338 B.n337 10.6151
R1007 B.n338 B.n115 10.6151
R1008 B.n349 B.n115 10.6151
R1009 B.n350 B.n349 10.6151
R1010 B.n351 B.n350 10.6151
R1011 B.n351 B.n108 10.6151
R1012 B.n362 B.n108 10.6151
R1013 B.n363 B.n362 10.6151
R1014 B.n364 B.n363 10.6151
R1015 B.n364 B.n101 10.6151
R1016 B.n375 B.n101 10.6151
R1017 B.n376 B.n375 10.6151
R1018 B.n377 B.n376 10.6151
R1019 B.n377 B.n94 10.6151
R1020 B.n388 B.n94 10.6151
R1021 B.n389 B.n388 10.6151
R1022 B.n390 B.n389 10.6151
R1023 B.n390 B.n0 10.6151
R1024 B.n616 B.n1 10.6151
R1025 B.n616 B.n615 10.6151
R1026 B.n615 B.n614 10.6151
R1027 B.n614 B.n10 10.6151
R1028 B.n608 B.n10 10.6151
R1029 B.n608 B.n607 10.6151
R1030 B.n607 B.n606 10.6151
R1031 B.n606 B.n16 10.6151
R1032 B.n600 B.n16 10.6151
R1033 B.n600 B.n599 10.6151
R1034 B.n599 B.n598 10.6151
R1035 B.n598 B.n23 10.6151
R1036 B.n592 B.n23 10.6151
R1037 B.n592 B.n591 10.6151
R1038 B.n591 B.n590 10.6151
R1039 B.n590 B.n30 10.6151
R1040 B.n584 B.n30 10.6151
R1041 B.n584 B.n583 10.6151
R1042 B.n583 B.n582 10.6151
R1043 B.n582 B.n38 10.6151
R1044 B.n576 B.n38 10.6151
R1045 B.n576 B.n575 10.6151
R1046 B.n575 B.n574 10.6151
R1047 B.n574 B.n45 10.6151
R1048 B.n568 B.n45 10.6151
R1049 B.n353 B.t1 9.19852
R1050 B.n594 B.t4 9.19852
R1051 B.n506 B.n68 6.7127
R1052 B.n491 B.n490 6.7127
R1053 B.n253 B.n157 6.7127
R1054 B.n237 B.n236 6.7127
R1055 B.n510 B.n68 3.90294
R1056 B.n490 B.n489 3.90294
R1057 B.n157 B.n153 3.90294
R1058 B.n236 B.n235 3.90294
R1059 B.n622 B.n0 2.81026
R1060 B.n622 B.n1 2.81026
R1061 B.n129 B.t9 2.50905
R1062 B.t13 B.n579 2.50905
R1063 B.n372 B.t6 0.836684
R1064 B.n18 B.t0 0.836684
R1065 VP.n7 VP.t5 281.168
R1066 VP.n17 VP.t4 258.06
R1067 VP.n29 VP.t3 258.06
R1068 VP.n15 VP.t0 258.06
R1069 VP.n22 VP.t7 213.109
R1070 VP.n1 VP.t2 213.109
R1071 VP.n5 VP.t1 213.109
R1072 VP.n8 VP.t6 213.109
R1073 VP.n30 VP.n29 161.3
R1074 VP.n9 VP.n6 161.3
R1075 VP.n11 VP.n10 161.3
R1076 VP.n13 VP.n12 161.3
R1077 VP.n14 VP.n4 161.3
R1078 VP.n16 VP.n15 161.3
R1079 VP.n28 VP.n0 161.3
R1080 VP.n27 VP.n26 161.3
R1081 VP.n25 VP.n24 161.3
R1082 VP.n23 VP.n2 161.3
R1083 VP.n21 VP.n20 161.3
R1084 VP.n19 VP.n3 161.3
R1085 VP.n18 VP.n17 161.3
R1086 VP.n24 VP.n23 56.4357
R1087 VP.n10 VP.n9 56.4357
R1088 VP.n21 VP.n3 43.2572
R1089 VP.n28 VP.n27 43.2572
R1090 VP.n14 VP.n13 43.2572
R1091 VP.n7 VP.n6 42.584
R1092 VP.n18 VP.n16 39.8338
R1093 VP.n8 VP.n7 35.9993
R1094 VP.n17 VP.n3 19.7187
R1095 VP.n29 VP.n28 19.7187
R1096 VP.n15 VP.n14 19.7187
R1097 VP.n23 VP.n22 17.4397
R1098 VP.n24 VP.n1 17.4397
R1099 VP.n10 VP.n5 17.4397
R1100 VP.n9 VP.n8 17.4397
R1101 VP.n22 VP.n21 6.78241
R1102 VP.n27 VP.n1 6.78241
R1103 VP.n13 VP.n5 6.78241
R1104 VP.n11 VP.n6 0.189894
R1105 VP.n12 VP.n11 0.189894
R1106 VP.n12 VP.n4 0.189894
R1107 VP.n16 VP.n4 0.189894
R1108 VP.n19 VP.n18 0.189894
R1109 VP.n20 VP.n19 0.189894
R1110 VP.n20 VP.n2 0.189894
R1111 VP.n25 VP.n2 0.189894
R1112 VP.n26 VP.n25 0.189894
R1113 VP.n26 VP.n0 0.189894
R1114 VP.n30 VP.n0 0.189894
R1115 VP VP.n30 0.0516364
R1116 VTAIL.n338 VTAIL.n302 289.615
R1117 VTAIL.n38 VTAIL.n2 289.615
R1118 VTAIL.n80 VTAIL.n44 289.615
R1119 VTAIL.n124 VTAIL.n88 289.615
R1120 VTAIL.n296 VTAIL.n260 289.615
R1121 VTAIL.n252 VTAIL.n216 289.615
R1122 VTAIL.n210 VTAIL.n174 289.615
R1123 VTAIL.n166 VTAIL.n130 289.615
R1124 VTAIL.n314 VTAIL.n313 185
R1125 VTAIL.n319 VTAIL.n318 185
R1126 VTAIL.n321 VTAIL.n320 185
R1127 VTAIL.n310 VTAIL.n309 185
R1128 VTAIL.n327 VTAIL.n326 185
R1129 VTAIL.n329 VTAIL.n328 185
R1130 VTAIL.n306 VTAIL.n305 185
R1131 VTAIL.n336 VTAIL.n335 185
R1132 VTAIL.n337 VTAIL.n304 185
R1133 VTAIL.n339 VTAIL.n338 185
R1134 VTAIL.n14 VTAIL.n13 185
R1135 VTAIL.n19 VTAIL.n18 185
R1136 VTAIL.n21 VTAIL.n20 185
R1137 VTAIL.n10 VTAIL.n9 185
R1138 VTAIL.n27 VTAIL.n26 185
R1139 VTAIL.n29 VTAIL.n28 185
R1140 VTAIL.n6 VTAIL.n5 185
R1141 VTAIL.n36 VTAIL.n35 185
R1142 VTAIL.n37 VTAIL.n4 185
R1143 VTAIL.n39 VTAIL.n38 185
R1144 VTAIL.n56 VTAIL.n55 185
R1145 VTAIL.n61 VTAIL.n60 185
R1146 VTAIL.n63 VTAIL.n62 185
R1147 VTAIL.n52 VTAIL.n51 185
R1148 VTAIL.n69 VTAIL.n68 185
R1149 VTAIL.n71 VTAIL.n70 185
R1150 VTAIL.n48 VTAIL.n47 185
R1151 VTAIL.n78 VTAIL.n77 185
R1152 VTAIL.n79 VTAIL.n46 185
R1153 VTAIL.n81 VTAIL.n80 185
R1154 VTAIL.n100 VTAIL.n99 185
R1155 VTAIL.n105 VTAIL.n104 185
R1156 VTAIL.n107 VTAIL.n106 185
R1157 VTAIL.n96 VTAIL.n95 185
R1158 VTAIL.n113 VTAIL.n112 185
R1159 VTAIL.n115 VTAIL.n114 185
R1160 VTAIL.n92 VTAIL.n91 185
R1161 VTAIL.n122 VTAIL.n121 185
R1162 VTAIL.n123 VTAIL.n90 185
R1163 VTAIL.n125 VTAIL.n124 185
R1164 VTAIL.n297 VTAIL.n296 185
R1165 VTAIL.n295 VTAIL.n262 185
R1166 VTAIL.n294 VTAIL.n293 185
R1167 VTAIL.n265 VTAIL.n263 185
R1168 VTAIL.n288 VTAIL.n287 185
R1169 VTAIL.n286 VTAIL.n285 185
R1170 VTAIL.n269 VTAIL.n268 185
R1171 VTAIL.n280 VTAIL.n279 185
R1172 VTAIL.n278 VTAIL.n277 185
R1173 VTAIL.n273 VTAIL.n272 185
R1174 VTAIL.n253 VTAIL.n252 185
R1175 VTAIL.n251 VTAIL.n218 185
R1176 VTAIL.n250 VTAIL.n249 185
R1177 VTAIL.n221 VTAIL.n219 185
R1178 VTAIL.n244 VTAIL.n243 185
R1179 VTAIL.n242 VTAIL.n241 185
R1180 VTAIL.n225 VTAIL.n224 185
R1181 VTAIL.n236 VTAIL.n235 185
R1182 VTAIL.n234 VTAIL.n233 185
R1183 VTAIL.n229 VTAIL.n228 185
R1184 VTAIL.n211 VTAIL.n210 185
R1185 VTAIL.n209 VTAIL.n176 185
R1186 VTAIL.n208 VTAIL.n207 185
R1187 VTAIL.n179 VTAIL.n177 185
R1188 VTAIL.n202 VTAIL.n201 185
R1189 VTAIL.n200 VTAIL.n199 185
R1190 VTAIL.n183 VTAIL.n182 185
R1191 VTAIL.n194 VTAIL.n193 185
R1192 VTAIL.n192 VTAIL.n191 185
R1193 VTAIL.n187 VTAIL.n186 185
R1194 VTAIL.n167 VTAIL.n166 185
R1195 VTAIL.n165 VTAIL.n132 185
R1196 VTAIL.n164 VTAIL.n163 185
R1197 VTAIL.n135 VTAIL.n133 185
R1198 VTAIL.n158 VTAIL.n157 185
R1199 VTAIL.n156 VTAIL.n155 185
R1200 VTAIL.n139 VTAIL.n138 185
R1201 VTAIL.n150 VTAIL.n149 185
R1202 VTAIL.n148 VTAIL.n147 185
R1203 VTAIL.n143 VTAIL.n142 185
R1204 VTAIL.n315 VTAIL.t6 149.524
R1205 VTAIL.n15 VTAIL.t2 149.524
R1206 VTAIL.n57 VTAIL.t11 149.524
R1207 VTAIL.n101 VTAIL.t9 149.524
R1208 VTAIL.n274 VTAIL.t12 149.524
R1209 VTAIL.n230 VTAIL.t8 149.524
R1210 VTAIL.n188 VTAIL.t3 149.524
R1211 VTAIL.n144 VTAIL.t0 149.524
R1212 VTAIL.n319 VTAIL.n313 104.615
R1213 VTAIL.n320 VTAIL.n319 104.615
R1214 VTAIL.n320 VTAIL.n309 104.615
R1215 VTAIL.n327 VTAIL.n309 104.615
R1216 VTAIL.n328 VTAIL.n327 104.615
R1217 VTAIL.n328 VTAIL.n305 104.615
R1218 VTAIL.n336 VTAIL.n305 104.615
R1219 VTAIL.n337 VTAIL.n336 104.615
R1220 VTAIL.n338 VTAIL.n337 104.615
R1221 VTAIL.n19 VTAIL.n13 104.615
R1222 VTAIL.n20 VTAIL.n19 104.615
R1223 VTAIL.n20 VTAIL.n9 104.615
R1224 VTAIL.n27 VTAIL.n9 104.615
R1225 VTAIL.n28 VTAIL.n27 104.615
R1226 VTAIL.n28 VTAIL.n5 104.615
R1227 VTAIL.n36 VTAIL.n5 104.615
R1228 VTAIL.n37 VTAIL.n36 104.615
R1229 VTAIL.n38 VTAIL.n37 104.615
R1230 VTAIL.n61 VTAIL.n55 104.615
R1231 VTAIL.n62 VTAIL.n61 104.615
R1232 VTAIL.n62 VTAIL.n51 104.615
R1233 VTAIL.n69 VTAIL.n51 104.615
R1234 VTAIL.n70 VTAIL.n69 104.615
R1235 VTAIL.n70 VTAIL.n47 104.615
R1236 VTAIL.n78 VTAIL.n47 104.615
R1237 VTAIL.n79 VTAIL.n78 104.615
R1238 VTAIL.n80 VTAIL.n79 104.615
R1239 VTAIL.n105 VTAIL.n99 104.615
R1240 VTAIL.n106 VTAIL.n105 104.615
R1241 VTAIL.n106 VTAIL.n95 104.615
R1242 VTAIL.n113 VTAIL.n95 104.615
R1243 VTAIL.n114 VTAIL.n113 104.615
R1244 VTAIL.n114 VTAIL.n91 104.615
R1245 VTAIL.n122 VTAIL.n91 104.615
R1246 VTAIL.n123 VTAIL.n122 104.615
R1247 VTAIL.n124 VTAIL.n123 104.615
R1248 VTAIL.n296 VTAIL.n295 104.615
R1249 VTAIL.n295 VTAIL.n294 104.615
R1250 VTAIL.n294 VTAIL.n263 104.615
R1251 VTAIL.n287 VTAIL.n263 104.615
R1252 VTAIL.n287 VTAIL.n286 104.615
R1253 VTAIL.n286 VTAIL.n268 104.615
R1254 VTAIL.n279 VTAIL.n268 104.615
R1255 VTAIL.n279 VTAIL.n278 104.615
R1256 VTAIL.n278 VTAIL.n272 104.615
R1257 VTAIL.n252 VTAIL.n251 104.615
R1258 VTAIL.n251 VTAIL.n250 104.615
R1259 VTAIL.n250 VTAIL.n219 104.615
R1260 VTAIL.n243 VTAIL.n219 104.615
R1261 VTAIL.n243 VTAIL.n242 104.615
R1262 VTAIL.n242 VTAIL.n224 104.615
R1263 VTAIL.n235 VTAIL.n224 104.615
R1264 VTAIL.n235 VTAIL.n234 104.615
R1265 VTAIL.n234 VTAIL.n228 104.615
R1266 VTAIL.n210 VTAIL.n209 104.615
R1267 VTAIL.n209 VTAIL.n208 104.615
R1268 VTAIL.n208 VTAIL.n177 104.615
R1269 VTAIL.n201 VTAIL.n177 104.615
R1270 VTAIL.n201 VTAIL.n200 104.615
R1271 VTAIL.n200 VTAIL.n182 104.615
R1272 VTAIL.n193 VTAIL.n182 104.615
R1273 VTAIL.n193 VTAIL.n192 104.615
R1274 VTAIL.n192 VTAIL.n186 104.615
R1275 VTAIL.n166 VTAIL.n165 104.615
R1276 VTAIL.n165 VTAIL.n164 104.615
R1277 VTAIL.n164 VTAIL.n133 104.615
R1278 VTAIL.n157 VTAIL.n133 104.615
R1279 VTAIL.n157 VTAIL.n156 104.615
R1280 VTAIL.n156 VTAIL.n138 104.615
R1281 VTAIL.n149 VTAIL.n138 104.615
R1282 VTAIL.n149 VTAIL.n148 104.615
R1283 VTAIL.n148 VTAIL.n142 104.615
R1284 VTAIL.t6 VTAIL.n313 52.3082
R1285 VTAIL.t2 VTAIL.n13 52.3082
R1286 VTAIL.t11 VTAIL.n55 52.3082
R1287 VTAIL.t9 VTAIL.n99 52.3082
R1288 VTAIL.t12 VTAIL.n272 52.3082
R1289 VTAIL.t8 VTAIL.n228 52.3082
R1290 VTAIL.t3 VTAIL.n186 52.3082
R1291 VTAIL.t0 VTAIL.n142 52.3082
R1292 VTAIL.n259 VTAIL.n258 48.6567
R1293 VTAIL.n173 VTAIL.n172 48.6567
R1294 VTAIL.n1 VTAIL.n0 48.6566
R1295 VTAIL.n87 VTAIL.n86 48.6566
R1296 VTAIL.n343 VTAIL.n342 33.5429
R1297 VTAIL.n43 VTAIL.n42 33.5429
R1298 VTAIL.n85 VTAIL.n84 33.5429
R1299 VTAIL.n129 VTAIL.n128 33.5429
R1300 VTAIL.n301 VTAIL.n300 33.5429
R1301 VTAIL.n257 VTAIL.n256 33.5429
R1302 VTAIL.n215 VTAIL.n214 33.5429
R1303 VTAIL.n171 VTAIL.n170 33.5429
R1304 VTAIL.n343 VTAIL.n301 20.2117
R1305 VTAIL.n171 VTAIL.n129 20.2117
R1306 VTAIL.n339 VTAIL.n304 13.1884
R1307 VTAIL.n39 VTAIL.n4 13.1884
R1308 VTAIL.n81 VTAIL.n46 13.1884
R1309 VTAIL.n125 VTAIL.n90 13.1884
R1310 VTAIL.n297 VTAIL.n262 13.1884
R1311 VTAIL.n253 VTAIL.n218 13.1884
R1312 VTAIL.n211 VTAIL.n176 13.1884
R1313 VTAIL.n167 VTAIL.n132 13.1884
R1314 VTAIL.n335 VTAIL.n334 12.8005
R1315 VTAIL.n340 VTAIL.n302 12.8005
R1316 VTAIL.n35 VTAIL.n34 12.8005
R1317 VTAIL.n40 VTAIL.n2 12.8005
R1318 VTAIL.n77 VTAIL.n76 12.8005
R1319 VTAIL.n82 VTAIL.n44 12.8005
R1320 VTAIL.n121 VTAIL.n120 12.8005
R1321 VTAIL.n126 VTAIL.n88 12.8005
R1322 VTAIL.n298 VTAIL.n260 12.8005
R1323 VTAIL.n293 VTAIL.n264 12.8005
R1324 VTAIL.n254 VTAIL.n216 12.8005
R1325 VTAIL.n249 VTAIL.n220 12.8005
R1326 VTAIL.n212 VTAIL.n174 12.8005
R1327 VTAIL.n207 VTAIL.n178 12.8005
R1328 VTAIL.n168 VTAIL.n130 12.8005
R1329 VTAIL.n163 VTAIL.n134 12.8005
R1330 VTAIL.n333 VTAIL.n306 12.0247
R1331 VTAIL.n33 VTAIL.n6 12.0247
R1332 VTAIL.n75 VTAIL.n48 12.0247
R1333 VTAIL.n119 VTAIL.n92 12.0247
R1334 VTAIL.n292 VTAIL.n265 12.0247
R1335 VTAIL.n248 VTAIL.n221 12.0247
R1336 VTAIL.n206 VTAIL.n179 12.0247
R1337 VTAIL.n162 VTAIL.n135 12.0247
R1338 VTAIL.n330 VTAIL.n329 11.249
R1339 VTAIL.n30 VTAIL.n29 11.249
R1340 VTAIL.n72 VTAIL.n71 11.249
R1341 VTAIL.n116 VTAIL.n115 11.249
R1342 VTAIL.n289 VTAIL.n288 11.249
R1343 VTAIL.n245 VTAIL.n244 11.249
R1344 VTAIL.n203 VTAIL.n202 11.249
R1345 VTAIL.n159 VTAIL.n158 11.249
R1346 VTAIL.n326 VTAIL.n308 10.4732
R1347 VTAIL.n26 VTAIL.n8 10.4732
R1348 VTAIL.n68 VTAIL.n50 10.4732
R1349 VTAIL.n112 VTAIL.n94 10.4732
R1350 VTAIL.n285 VTAIL.n267 10.4732
R1351 VTAIL.n241 VTAIL.n223 10.4732
R1352 VTAIL.n199 VTAIL.n181 10.4732
R1353 VTAIL.n155 VTAIL.n137 10.4732
R1354 VTAIL.n315 VTAIL.n314 10.2747
R1355 VTAIL.n15 VTAIL.n14 10.2747
R1356 VTAIL.n57 VTAIL.n56 10.2747
R1357 VTAIL.n101 VTAIL.n100 10.2747
R1358 VTAIL.n274 VTAIL.n273 10.2747
R1359 VTAIL.n230 VTAIL.n229 10.2747
R1360 VTAIL.n188 VTAIL.n187 10.2747
R1361 VTAIL.n144 VTAIL.n143 10.2747
R1362 VTAIL.n325 VTAIL.n310 9.69747
R1363 VTAIL.n25 VTAIL.n10 9.69747
R1364 VTAIL.n67 VTAIL.n52 9.69747
R1365 VTAIL.n111 VTAIL.n96 9.69747
R1366 VTAIL.n284 VTAIL.n269 9.69747
R1367 VTAIL.n240 VTAIL.n225 9.69747
R1368 VTAIL.n198 VTAIL.n183 9.69747
R1369 VTAIL.n154 VTAIL.n139 9.69747
R1370 VTAIL.n342 VTAIL.n341 9.45567
R1371 VTAIL.n42 VTAIL.n41 9.45567
R1372 VTAIL.n84 VTAIL.n83 9.45567
R1373 VTAIL.n128 VTAIL.n127 9.45567
R1374 VTAIL.n300 VTAIL.n299 9.45567
R1375 VTAIL.n256 VTAIL.n255 9.45567
R1376 VTAIL.n214 VTAIL.n213 9.45567
R1377 VTAIL.n170 VTAIL.n169 9.45567
R1378 VTAIL.n341 VTAIL.n340 9.3005
R1379 VTAIL.n317 VTAIL.n316 9.3005
R1380 VTAIL.n312 VTAIL.n311 9.3005
R1381 VTAIL.n323 VTAIL.n322 9.3005
R1382 VTAIL.n325 VTAIL.n324 9.3005
R1383 VTAIL.n308 VTAIL.n307 9.3005
R1384 VTAIL.n331 VTAIL.n330 9.3005
R1385 VTAIL.n333 VTAIL.n332 9.3005
R1386 VTAIL.n334 VTAIL.n303 9.3005
R1387 VTAIL.n41 VTAIL.n40 9.3005
R1388 VTAIL.n17 VTAIL.n16 9.3005
R1389 VTAIL.n12 VTAIL.n11 9.3005
R1390 VTAIL.n23 VTAIL.n22 9.3005
R1391 VTAIL.n25 VTAIL.n24 9.3005
R1392 VTAIL.n8 VTAIL.n7 9.3005
R1393 VTAIL.n31 VTAIL.n30 9.3005
R1394 VTAIL.n33 VTAIL.n32 9.3005
R1395 VTAIL.n34 VTAIL.n3 9.3005
R1396 VTAIL.n83 VTAIL.n82 9.3005
R1397 VTAIL.n59 VTAIL.n58 9.3005
R1398 VTAIL.n54 VTAIL.n53 9.3005
R1399 VTAIL.n65 VTAIL.n64 9.3005
R1400 VTAIL.n67 VTAIL.n66 9.3005
R1401 VTAIL.n50 VTAIL.n49 9.3005
R1402 VTAIL.n73 VTAIL.n72 9.3005
R1403 VTAIL.n75 VTAIL.n74 9.3005
R1404 VTAIL.n76 VTAIL.n45 9.3005
R1405 VTAIL.n127 VTAIL.n126 9.3005
R1406 VTAIL.n103 VTAIL.n102 9.3005
R1407 VTAIL.n98 VTAIL.n97 9.3005
R1408 VTAIL.n109 VTAIL.n108 9.3005
R1409 VTAIL.n111 VTAIL.n110 9.3005
R1410 VTAIL.n94 VTAIL.n93 9.3005
R1411 VTAIL.n117 VTAIL.n116 9.3005
R1412 VTAIL.n119 VTAIL.n118 9.3005
R1413 VTAIL.n120 VTAIL.n89 9.3005
R1414 VTAIL.n276 VTAIL.n275 9.3005
R1415 VTAIL.n271 VTAIL.n270 9.3005
R1416 VTAIL.n282 VTAIL.n281 9.3005
R1417 VTAIL.n284 VTAIL.n283 9.3005
R1418 VTAIL.n267 VTAIL.n266 9.3005
R1419 VTAIL.n290 VTAIL.n289 9.3005
R1420 VTAIL.n292 VTAIL.n291 9.3005
R1421 VTAIL.n264 VTAIL.n261 9.3005
R1422 VTAIL.n299 VTAIL.n298 9.3005
R1423 VTAIL.n232 VTAIL.n231 9.3005
R1424 VTAIL.n227 VTAIL.n226 9.3005
R1425 VTAIL.n238 VTAIL.n237 9.3005
R1426 VTAIL.n240 VTAIL.n239 9.3005
R1427 VTAIL.n223 VTAIL.n222 9.3005
R1428 VTAIL.n246 VTAIL.n245 9.3005
R1429 VTAIL.n248 VTAIL.n247 9.3005
R1430 VTAIL.n220 VTAIL.n217 9.3005
R1431 VTAIL.n255 VTAIL.n254 9.3005
R1432 VTAIL.n190 VTAIL.n189 9.3005
R1433 VTAIL.n185 VTAIL.n184 9.3005
R1434 VTAIL.n196 VTAIL.n195 9.3005
R1435 VTAIL.n198 VTAIL.n197 9.3005
R1436 VTAIL.n181 VTAIL.n180 9.3005
R1437 VTAIL.n204 VTAIL.n203 9.3005
R1438 VTAIL.n206 VTAIL.n205 9.3005
R1439 VTAIL.n178 VTAIL.n175 9.3005
R1440 VTAIL.n213 VTAIL.n212 9.3005
R1441 VTAIL.n146 VTAIL.n145 9.3005
R1442 VTAIL.n141 VTAIL.n140 9.3005
R1443 VTAIL.n152 VTAIL.n151 9.3005
R1444 VTAIL.n154 VTAIL.n153 9.3005
R1445 VTAIL.n137 VTAIL.n136 9.3005
R1446 VTAIL.n160 VTAIL.n159 9.3005
R1447 VTAIL.n162 VTAIL.n161 9.3005
R1448 VTAIL.n134 VTAIL.n131 9.3005
R1449 VTAIL.n169 VTAIL.n168 9.3005
R1450 VTAIL.n322 VTAIL.n321 8.92171
R1451 VTAIL.n22 VTAIL.n21 8.92171
R1452 VTAIL.n64 VTAIL.n63 8.92171
R1453 VTAIL.n108 VTAIL.n107 8.92171
R1454 VTAIL.n281 VTAIL.n280 8.92171
R1455 VTAIL.n237 VTAIL.n236 8.92171
R1456 VTAIL.n195 VTAIL.n194 8.92171
R1457 VTAIL.n151 VTAIL.n150 8.92171
R1458 VTAIL.n318 VTAIL.n312 8.14595
R1459 VTAIL.n18 VTAIL.n12 8.14595
R1460 VTAIL.n60 VTAIL.n54 8.14595
R1461 VTAIL.n104 VTAIL.n98 8.14595
R1462 VTAIL.n277 VTAIL.n271 8.14595
R1463 VTAIL.n233 VTAIL.n227 8.14595
R1464 VTAIL.n191 VTAIL.n185 8.14595
R1465 VTAIL.n147 VTAIL.n141 8.14595
R1466 VTAIL.n317 VTAIL.n314 7.3702
R1467 VTAIL.n17 VTAIL.n14 7.3702
R1468 VTAIL.n59 VTAIL.n56 7.3702
R1469 VTAIL.n103 VTAIL.n100 7.3702
R1470 VTAIL.n276 VTAIL.n273 7.3702
R1471 VTAIL.n232 VTAIL.n229 7.3702
R1472 VTAIL.n190 VTAIL.n187 7.3702
R1473 VTAIL.n146 VTAIL.n143 7.3702
R1474 VTAIL.n318 VTAIL.n317 5.81868
R1475 VTAIL.n18 VTAIL.n17 5.81868
R1476 VTAIL.n60 VTAIL.n59 5.81868
R1477 VTAIL.n104 VTAIL.n103 5.81868
R1478 VTAIL.n277 VTAIL.n276 5.81868
R1479 VTAIL.n233 VTAIL.n232 5.81868
R1480 VTAIL.n191 VTAIL.n190 5.81868
R1481 VTAIL.n147 VTAIL.n146 5.81868
R1482 VTAIL.n321 VTAIL.n312 5.04292
R1483 VTAIL.n21 VTAIL.n12 5.04292
R1484 VTAIL.n63 VTAIL.n54 5.04292
R1485 VTAIL.n107 VTAIL.n98 5.04292
R1486 VTAIL.n280 VTAIL.n271 5.04292
R1487 VTAIL.n236 VTAIL.n227 5.04292
R1488 VTAIL.n194 VTAIL.n185 5.04292
R1489 VTAIL.n150 VTAIL.n141 5.04292
R1490 VTAIL.n322 VTAIL.n310 4.26717
R1491 VTAIL.n22 VTAIL.n10 4.26717
R1492 VTAIL.n64 VTAIL.n52 4.26717
R1493 VTAIL.n108 VTAIL.n96 4.26717
R1494 VTAIL.n281 VTAIL.n269 4.26717
R1495 VTAIL.n237 VTAIL.n225 4.26717
R1496 VTAIL.n195 VTAIL.n183 4.26717
R1497 VTAIL.n151 VTAIL.n139 4.26717
R1498 VTAIL.n326 VTAIL.n325 3.49141
R1499 VTAIL.n26 VTAIL.n25 3.49141
R1500 VTAIL.n68 VTAIL.n67 3.49141
R1501 VTAIL.n112 VTAIL.n111 3.49141
R1502 VTAIL.n285 VTAIL.n284 3.49141
R1503 VTAIL.n241 VTAIL.n240 3.49141
R1504 VTAIL.n199 VTAIL.n198 3.49141
R1505 VTAIL.n155 VTAIL.n154 3.49141
R1506 VTAIL.n316 VTAIL.n315 2.84304
R1507 VTAIL.n16 VTAIL.n15 2.84304
R1508 VTAIL.n58 VTAIL.n57 2.84304
R1509 VTAIL.n102 VTAIL.n101 2.84304
R1510 VTAIL.n275 VTAIL.n274 2.84304
R1511 VTAIL.n231 VTAIL.n230 2.84304
R1512 VTAIL.n189 VTAIL.n188 2.84304
R1513 VTAIL.n145 VTAIL.n144 2.84304
R1514 VTAIL.n329 VTAIL.n308 2.71565
R1515 VTAIL.n29 VTAIL.n8 2.71565
R1516 VTAIL.n71 VTAIL.n50 2.71565
R1517 VTAIL.n115 VTAIL.n94 2.71565
R1518 VTAIL.n288 VTAIL.n267 2.71565
R1519 VTAIL.n244 VTAIL.n223 2.71565
R1520 VTAIL.n202 VTAIL.n181 2.71565
R1521 VTAIL.n158 VTAIL.n137 2.71565
R1522 VTAIL.n0 VTAIL.t1 2.51638
R1523 VTAIL.n0 VTAIL.t4 2.51638
R1524 VTAIL.n86 VTAIL.t15 2.51638
R1525 VTAIL.n86 VTAIL.t14 2.51638
R1526 VTAIL.n258 VTAIL.t10 2.51638
R1527 VTAIL.n258 VTAIL.t13 2.51638
R1528 VTAIL.n172 VTAIL.t7 2.51638
R1529 VTAIL.n172 VTAIL.t5 2.51638
R1530 VTAIL.n330 VTAIL.n306 1.93989
R1531 VTAIL.n30 VTAIL.n6 1.93989
R1532 VTAIL.n72 VTAIL.n48 1.93989
R1533 VTAIL.n116 VTAIL.n92 1.93989
R1534 VTAIL.n289 VTAIL.n265 1.93989
R1535 VTAIL.n245 VTAIL.n221 1.93989
R1536 VTAIL.n203 VTAIL.n179 1.93989
R1537 VTAIL.n159 VTAIL.n135 1.93989
R1538 VTAIL.n335 VTAIL.n333 1.16414
R1539 VTAIL.n342 VTAIL.n302 1.16414
R1540 VTAIL.n35 VTAIL.n33 1.16414
R1541 VTAIL.n42 VTAIL.n2 1.16414
R1542 VTAIL.n77 VTAIL.n75 1.16414
R1543 VTAIL.n84 VTAIL.n44 1.16414
R1544 VTAIL.n121 VTAIL.n119 1.16414
R1545 VTAIL.n128 VTAIL.n88 1.16414
R1546 VTAIL.n300 VTAIL.n260 1.16414
R1547 VTAIL.n293 VTAIL.n292 1.16414
R1548 VTAIL.n256 VTAIL.n216 1.16414
R1549 VTAIL.n249 VTAIL.n248 1.16414
R1550 VTAIL.n214 VTAIL.n174 1.16414
R1551 VTAIL.n207 VTAIL.n206 1.16414
R1552 VTAIL.n170 VTAIL.n130 1.16414
R1553 VTAIL.n163 VTAIL.n162 1.16414
R1554 VTAIL.n173 VTAIL.n171 1.05222
R1555 VTAIL.n215 VTAIL.n173 1.05222
R1556 VTAIL.n259 VTAIL.n257 1.05222
R1557 VTAIL.n301 VTAIL.n259 1.05222
R1558 VTAIL.n129 VTAIL.n87 1.05222
R1559 VTAIL.n87 VTAIL.n85 1.05222
R1560 VTAIL.n43 VTAIL.n1 1.05222
R1561 VTAIL VTAIL.n343 0.994035
R1562 VTAIL.n257 VTAIL.n215 0.470328
R1563 VTAIL.n85 VTAIL.n43 0.470328
R1564 VTAIL.n334 VTAIL.n304 0.388379
R1565 VTAIL.n340 VTAIL.n339 0.388379
R1566 VTAIL.n34 VTAIL.n4 0.388379
R1567 VTAIL.n40 VTAIL.n39 0.388379
R1568 VTAIL.n76 VTAIL.n46 0.388379
R1569 VTAIL.n82 VTAIL.n81 0.388379
R1570 VTAIL.n120 VTAIL.n90 0.388379
R1571 VTAIL.n126 VTAIL.n125 0.388379
R1572 VTAIL.n298 VTAIL.n297 0.388379
R1573 VTAIL.n264 VTAIL.n262 0.388379
R1574 VTAIL.n254 VTAIL.n253 0.388379
R1575 VTAIL.n220 VTAIL.n218 0.388379
R1576 VTAIL.n212 VTAIL.n211 0.388379
R1577 VTAIL.n178 VTAIL.n176 0.388379
R1578 VTAIL.n168 VTAIL.n167 0.388379
R1579 VTAIL.n134 VTAIL.n132 0.388379
R1580 VTAIL.n316 VTAIL.n311 0.155672
R1581 VTAIL.n323 VTAIL.n311 0.155672
R1582 VTAIL.n324 VTAIL.n323 0.155672
R1583 VTAIL.n324 VTAIL.n307 0.155672
R1584 VTAIL.n331 VTAIL.n307 0.155672
R1585 VTAIL.n332 VTAIL.n331 0.155672
R1586 VTAIL.n332 VTAIL.n303 0.155672
R1587 VTAIL.n341 VTAIL.n303 0.155672
R1588 VTAIL.n16 VTAIL.n11 0.155672
R1589 VTAIL.n23 VTAIL.n11 0.155672
R1590 VTAIL.n24 VTAIL.n23 0.155672
R1591 VTAIL.n24 VTAIL.n7 0.155672
R1592 VTAIL.n31 VTAIL.n7 0.155672
R1593 VTAIL.n32 VTAIL.n31 0.155672
R1594 VTAIL.n32 VTAIL.n3 0.155672
R1595 VTAIL.n41 VTAIL.n3 0.155672
R1596 VTAIL.n58 VTAIL.n53 0.155672
R1597 VTAIL.n65 VTAIL.n53 0.155672
R1598 VTAIL.n66 VTAIL.n65 0.155672
R1599 VTAIL.n66 VTAIL.n49 0.155672
R1600 VTAIL.n73 VTAIL.n49 0.155672
R1601 VTAIL.n74 VTAIL.n73 0.155672
R1602 VTAIL.n74 VTAIL.n45 0.155672
R1603 VTAIL.n83 VTAIL.n45 0.155672
R1604 VTAIL.n102 VTAIL.n97 0.155672
R1605 VTAIL.n109 VTAIL.n97 0.155672
R1606 VTAIL.n110 VTAIL.n109 0.155672
R1607 VTAIL.n110 VTAIL.n93 0.155672
R1608 VTAIL.n117 VTAIL.n93 0.155672
R1609 VTAIL.n118 VTAIL.n117 0.155672
R1610 VTAIL.n118 VTAIL.n89 0.155672
R1611 VTAIL.n127 VTAIL.n89 0.155672
R1612 VTAIL.n299 VTAIL.n261 0.155672
R1613 VTAIL.n291 VTAIL.n261 0.155672
R1614 VTAIL.n291 VTAIL.n290 0.155672
R1615 VTAIL.n290 VTAIL.n266 0.155672
R1616 VTAIL.n283 VTAIL.n266 0.155672
R1617 VTAIL.n283 VTAIL.n282 0.155672
R1618 VTAIL.n282 VTAIL.n270 0.155672
R1619 VTAIL.n275 VTAIL.n270 0.155672
R1620 VTAIL.n255 VTAIL.n217 0.155672
R1621 VTAIL.n247 VTAIL.n217 0.155672
R1622 VTAIL.n247 VTAIL.n246 0.155672
R1623 VTAIL.n246 VTAIL.n222 0.155672
R1624 VTAIL.n239 VTAIL.n222 0.155672
R1625 VTAIL.n239 VTAIL.n238 0.155672
R1626 VTAIL.n238 VTAIL.n226 0.155672
R1627 VTAIL.n231 VTAIL.n226 0.155672
R1628 VTAIL.n213 VTAIL.n175 0.155672
R1629 VTAIL.n205 VTAIL.n175 0.155672
R1630 VTAIL.n205 VTAIL.n204 0.155672
R1631 VTAIL.n204 VTAIL.n180 0.155672
R1632 VTAIL.n197 VTAIL.n180 0.155672
R1633 VTAIL.n197 VTAIL.n196 0.155672
R1634 VTAIL.n196 VTAIL.n184 0.155672
R1635 VTAIL.n189 VTAIL.n184 0.155672
R1636 VTAIL.n169 VTAIL.n131 0.155672
R1637 VTAIL.n161 VTAIL.n131 0.155672
R1638 VTAIL.n161 VTAIL.n160 0.155672
R1639 VTAIL.n160 VTAIL.n136 0.155672
R1640 VTAIL.n153 VTAIL.n136 0.155672
R1641 VTAIL.n153 VTAIL.n152 0.155672
R1642 VTAIL.n152 VTAIL.n140 0.155672
R1643 VTAIL.n145 VTAIL.n140 0.155672
R1644 VTAIL VTAIL.n1 0.0586897
R1645 VDD1 VDD1.n0 65.9196
R1646 VDD1.n3 VDD1.n2 65.8059
R1647 VDD1.n3 VDD1.n1 65.8059
R1648 VDD1.n5 VDD1.n4 65.3354
R1649 VDD1.n5 VDD1.n3 35.8242
R1650 VDD1.n4 VDD1.t6 2.51638
R1651 VDD1.n4 VDD1.t7 2.51638
R1652 VDD1.n0 VDD1.t2 2.51638
R1653 VDD1.n0 VDD1.t1 2.51638
R1654 VDD1.n2 VDD1.t5 2.51638
R1655 VDD1.n2 VDD1.t4 2.51638
R1656 VDD1.n1 VDD1.t3 2.51638
R1657 VDD1.n1 VDD1.t0 2.51638
R1658 VDD1 VDD1.n5 0.468172
R1659 VN.n3 VN.t7 281.168
R1660 VN.n16 VN.t0 281.168
R1661 VN.n11 VN.t5 258.06
R1662 VN.n24 VN.t6 258.06
R1663 VN.n4 VN.t3 213.109
R1664 VN.n1 VN.t1 213.109
R1665 VN.n17 VN.t2 213.109
R1666 VN.n14 VN.t4 213.109
R1667 VN.n12 VN.n11 161.3
R1668 VN.n25 VN.n24 161.3
R1669 VN.n23 VN.n13 161.3
R1670 VN.n22 VN.n21 161.3
R1671 VN.n20 VN.n19 161.3
R1672 VN.n18 VN.n15 161.3
R1673 VN.n10 VN.n0 161.3
R1674 VN.n9 VN.n8 161.3
R1675 VN.n7 VN.n6 161.3
R1676 VN.n5 VN.n2 161.3
R1677 VN.n6 VN.n5 56.4357
R1678 VN.n19 VN.n18 56.4357
R1679 VN.n10 VN.n9 43.2572
R1680 VN.n23 VN.n22 43.2572
R1681 VN.n16 VN.n15 42.584
R1682 VN.n3 VN.n2 42.584
R1683 VN VN.n25 40.2145
R1684 VN.n4 VN.n3 35.9993
R1685 VN.n17 VN.n16 35.9993
R1686 VN.n11 VN.n10 19.7187
R1687 VN.n24 VN.n23 19.7187
R1688 VN.n5 VN.n4 17.4397
R1689 VN.n6 VN.n1 17.4397
R1690 VN.n18 VN.n17 17.4397
R1691 VN.n19 VN.n14 17.4397
R1692 VN.n9 VN.n1 6.78241
R1693 VN.n22 VN.n14 6.78241
R1694 VN.n25 VN.n13 0.189894
R1695 VN.n21 VN.n13 0.189894
R1696 VN.n21 VN.n20 0.189894
R1697 VN.n20 VN.n15 0.189894
R1698 VN.n7 VN.n2 0.189894
R1699 VN.n8 VN.n7 0.189894
R1700 VN.n8 VN.n0 0.189894
R1701 VN.n12 VN.n0 0.189894
R1702 VN VN.n12 0.0516364
R1703 VDD2.n2 VDD2.n1 65.8059
R1704 VDD2.n2 VDD2.n0 65.8059
R1705 VDD2 VDD2.n5 65.803
R1706 VDD2.n4 VDD2.n3 65.3355
R1707 VDD2.n4 VDD2.n2 35.2412
R1708 VDD2.n5 VDD2.t5 2.51638
R1709 VDD2.n5 VDD2.t7 2.51638
R1710 VDD2.n3 VDD2.t1 2.51638
R1711 VDD2.n3 VDD2.t3 2.51638
R1712 VDD2.n1 VDD2.t6 2.51638
R1713 VDD2.n1 VDD2.t2 2.51638
R1714 VDD2.n0 VDD2.t0 2.51638
R1715 VDD2.n0 VDD2.t4 2.51638
R1716 VDD2 VDD2.n4 0.584552
C0 VP VDD1 4.38975f
C1 VTAIL VDD1 7.35904f
C2 VDD2 VDD1 0.917585f
C3 VP VN 4.8056f
C4 VTAIL VN 4.18762f
C5 VDD2 VN 4.20121f
C6 VDD1 VN 0.148196f
C7 VP VTAIL 4.20172f
C8 VDD2 VP 0.33727f
C9 VDD2 VTAIL 7.40199f
C10 VDD2 B 3.339469f
C11 VDD1 B 3.59645f
C12 VTAIL B 6.762576f
C13 VN B 8.78133f
C14 VP B 7.11094f
C15 VDD2.t0 B 0.16266f
C16 VDD2.t4 B 0.16266f
C17 VDD2.n0 B 1.40908f
C18 VDD2.t6 B 0.16266f
C19 VDD2.t2 B 0.16266f
C20 VDD2.n1 B 1.40908f
C21 VDD2.n2 B 2.11278f
C22 VDD2.t1 B 0.16266f
C23 VDD2.t3 B 0.16266f
C24 VDD2.n3 B 1.4066f
C25 VDD2.n4 B 2.11969f
C26 VDD2.t5 B 0.16266f
C27 VDD2.t7 B 0.16266f
C28 VDD2.n5 B 1.40905f
C29 VN.n0 B 0.0407f
C30 VN.t1 B 0.764397f
C31 VN.n1 B 0.304134f
C32 VN.n2 B 0.175697f
C33 VN.t3 B 0.764397f
C34 VN.t7 B 0.850039f
C35 VN.n3 B 0.346667f
C36 VN.n4 B 0.349874f
C37 VN.n5 B 0.049332f
C38 VN.n6 B 0.049332f
C39 VN.n7 B 0.0407f
C40 VN.n8 B 0.0407f
C41 VN.n9 B 0.053036f
C42 VN.n10 B 0.018788f
C43 VN.t5 B 0.820568f
C44 VN.n11 B 0.34915f
C45 VN.n12 B 0.031541f
C46 VN.n13 B 0.0407f
C47 VN.t4 B 0.764397f
C48 VN.n14 B 0.304134f
C49 VN.n15 B 0.175697f
C50 VN.t2 B 0.764397f
C51 VN.t0 B 0.850039f
C52 VN.n16 B 0.346667f
C53 VN.n17 B 0.349874f
C54 VN.n18 B 0.049332f
C55 VN.n19 B 0.049332f
C56 VN.n20 B 0.0407f
C57 VN.n21 B 0.0407f
C58 VN.n22 B 0.053036f
C59 VN.n23 B 0.018788f
C60 VN.t6 B 0.820568f
C61 VN.n24 B 0.34915f
C62 VN.n25 B 1.56233f
C63 VDD1.t2 B 0.164097f
C64 VDD1.t1 B 0.164097f
C65 VDD1.n0 B 1.42221f
C66 VDD1.t3 B 0.164097f
C67 VDD1.t0 B 0.164097f
C68 VDD1.n1 B 1.42153f
C69 VDD1.t5 B 0.164097f
C70 VDD1.t4 B 0.164097f
C71 VDD1.n2 B 1.42153f
C72 VDD1.n3 B 2.1878f
C73 VDD1.t6 B 0.164097f
C74 VDD1.t7 B 0.164097f
C75 VDD1.n4 B 1.41903f
C76 VDD1.n5 B 2.16965f
C77 VTAIL.t1 B 0.128195f
C78 VTAIL.t4 B 0.128195f
C79 VTAIL.n0 B 1.0538f
C80 VTAIL.n1 B 0.264151f
C81 VTAIL.n2 B 0.026609f
C82 VTAIL.n3 B 0.020613f
C83 VTAIL.n4 B 0.011402f
C84 VTAIL.n5 B 0.026181f
C85 VTAIL.n6 B 0.011728f
C86 VTAIL.n7 B 0.020613f
C87 VTAIL.n8 B 0.011077f
C88 VTAIL.n9 B 0.026181f
C89 VTAIL.n10 B 0.011728f
C90 VTAIL.n11 B 0.020613f
C91 VTAIL.n12 B 0.011077f
C92 VTAIL.n13 B 0.019636f
C93 VTAIL.n14 B 0.018508f
C94 VTAIL.t2 B 0.043771f
C95 VTAIL.n15 B 0.115955f
C96 VTAIL.n16 B 0.661205f
C97 VTAIL.n17 B 0.011077f
C98 VTAIL.n18 B 0.011728f
C99 VTAIL.n19 B 0.026181f
C100 VTAIL.n20 B 0.026181f
C101 VTAIL.n21 B 0.011728f
C102 VTAIL.n22 B 0.011077f
C103 VTAIL.n23 B 0.020613f
C104 VTAIL.n24 B 0.020613f
C105 VTAIL.n25 B 0.011077f
C106 VTAIL.n26 B 0.011728f
C107 VTAIL.n27 B 0.026181f
C108 VTAIL.n28 B 0.026181f
C109 VTAIL.n29 B 0.011728f
C110 VTAIL.n30 B 0.011077f
C111 VTAIL.n31 B 0.020613f
C112 VTAIL.n32 B 0.020613f
C113 VTAIL.n33 B 0.011077f
C114 VTAIL.n34 B 0.011077f
C115 VTAIL.n35 B 0.011728f
C116 VTAIL.n36 B 0.026181f
C117 VTAIL.n37 B 0.026181f
C118 VTAIL.n38 B 0.052496f
C119 VTAIL.n39 B 0.011402f
C120 VTAIL.n40 B 0.011077f
C121 VTAIL.n41 B 0.049617f
C122 VTAIL.n42 B 0.029003f
C123 VTAIL.n43 B 0.11978f
C124 VTAIL.n44 B 0.026609f
C125 VTAIL.n45 B 0.020613f
C126 VTAIL.n46 B 0.011402f
C127 VTAIL.n47 B 0.026181f
C128 VTAIL.n48 B 0.011728f
C129 VTAIL.n49 B 0.020613f
C130 VTAIL.n50 B 0.011077f
C131 VTAIL.n51 B 0.026181f
C132 VTAIL.n52 B 0.011728f
C133 VTAIL.n53 B 0.020613f
C134 VTAIL.n54 B 0.011077f
C135 VTAIL.n55 B 0.019636f
C136 VTAIL.n56 B 0.018508f
C137 VTAIL.t11 B 0.043771f
C138 VTAIL.n57 B 0.115955f
C139 VTAIL.n58 B 0.661205f
C140 VTAIL.n59 B 0.011077f
C141 VTAIL.n60 B 0.011728f
C142 VTAIL.n61 B 0.026181f
C143 VTAIL.n62 B 0.026181f
C144 VTAIL.n63 B 0.011728f
C145 VTAIL.n64 B 0.011077f
C146 VTAIL.n65 B 0.020613f
C147 VTAIL.n66 B 0.020613f
C148 VTAIL.n67 B 0.011077f
C149 VTAIL.n68 B 0.011728f
C150 VTAIL.n69 B 0.026181f
C151 VTAIL.n70 B 0.026181f
C152 VTAIL.n71 B 0.011728f
C153 VTAIL.n72 B 0.011077f
C154 VTAIL.n73 B 0.020613f
C155 VTAIL.n74 B 0.020613f
C156 VTAIL.n75 B 0.011077f
C157 VTAIL.n76 B 0.011077f
C158 VTAIL.n77 B 0.011728f
C159 VTAIL.n78 B 0.026181f
C160 VTAIL.n79 B 0.026181f
C161 VTAIL.n80 B 0.052496f
C162 VTAIL.n81 B 0.011402f
C163 VTAIL.n82 B 0.011077f
C164 VTAIL.n83 B 0.049617f
C165 VTAIL.n84 B 0.029003f
C166 VTAIL.n85 B 0.11978f
C167 VTAIL.t15 B 0.128195f
C168 VTAIL.t14 B 0.128195f
C169 VTAIL.n86 B 1.0538f
C170 VTAIL.n87 B 0.330142f
C171 VTAIL.n88 B 0.026609f
C172 VTAIL.n89 B 0.020613f
C173 VTAIL.n90 B 0.011402f
C174 VTAIL.n91 B 0.026181f
C175 VTAIL.n92 B 0.011728f
C176 VTAIL.n93 B 0.020613f
C177 VTAIL.n94 B 0.011077f
C178 VTAIL.n95 B 0.026181f
C179 VTAIL.n96 B 0.011728f
C180 VTAIL.n97 B 0.020613f
C181 VTAIL.n98 B 0.011077f
C182 VTAIL.n99 B 0.019636f
C183 VTAIL.n100 B 0.018508f
C184 VTAIL.t9 B 0.043771f
C185 VTAIL.n101 B 0.115955f
C186 VTAIL.n102 B 0.661205f
C187 VTAIL.n103 B 0.011077f
C188 VTAIL.n104 B 0.011728f
C189 VTAIL.n105 B 0.026181f
C190 VTAIL.n106 B 0.026181f
C191 VTAIL.n107 B 0.011728f
C192 VTAIL.n108 B 0.011077f
C193 VTAIL.n109 B 0.020613f
C194 VTAIL.n110 B 0.020613f
C195 VTAIL.n111 B 0.011077f
C196 VTAIL.n112 B 0.011728f
C197 VTAIL.n113 B 0.026181f
C198 VTAIL.n114 B 0.026181f
C199 VTAIL.n115 B 0.011728f
C200 VTAIL.n116 B 0.011077f
C201 VTAIL.n117 B 0.020613f
C202 VTAIL.n118 B 0.020613f
C203 VTAIL.n119 B 0.011077f
C204 VTAIL.n120 B 0.011077f
C205 VTAIL.n121 B 0.011728f
C206 VTAIL.n122 B 0.026181f
C207 VTAIL.n123 B 0.026181f
C208 VTAIL.n124 B 0.052496f
C209 VTAIL.n125 B 0.011402f
C210 VTAIL.n126 B 0.011077f
C211 VTAIL.n127 B 0.049617f
C212 VTAIL.n128 B 0.029003f
C213 VTAIL.n129 B 0.88963f
C214 VTAIL.n130 B 0.026609f
C215 VTAIL.n131 B 0.020613f
C216 VTAIL.n132 B 0.011402f
C217 VTAIL.n133 B 0.026181f
C218 VTAIL.n134 B 0.011077f
C219 VTAIL.n135 B 0.011728f
C220 VTAIL.n136 B 0.020613f
C221 VTAIL.n137 B 0.011077f
C222 VTAIL.n138 B 0.026181f
C223 VTAIL.n139 B 0.011728f
C224 VTAIL.n140 B 0.020613f
C225 VTAIL.n141 B 0.011077f
C226 VTAIL.n142 B 0.019636f
C227 VTAIL.n143 B 0.018508f
C228 VTAIL.t0 B 0.043771f
C229 VTAIL.n144 B 0.115955f
C230 VTAIL.n145 B 0.661205f
C231 VTAIL.n146 B 0.011077f
C232 VTAIL.n147 B 0.011728f
C233 VTAIL.n148 B 0.026181f
C234 VTAIL.n149 B 0.026181f
C235 VTAIL.n150 B 0.011728f
C236 VTAIL.n151 B 0.011077f
C237 VTAIL.n152 B 0.020613f
C238 VTAIL.n153 B 0.020613f
C239 VTAIL.n154 B 0.011077f
C240 VTAIL.n155 B 0.011728f
C241 VTAIL.n156 B 0.026181f
C242 VTAIL.n157 B 0.026181f
C243 VTAIL.n158 B 0.011728f
C244 VTAIL.n159 B 0.011077f
C245 VTAIL.n160 B 0.020613f
C246 VTAIL.n161 B 0.020613f
C247 VTAIL.n162 B 0.011077f
C248 VTAIL.n163 B 0.011728f
C249 VTAIL.n164 B 0.026181f
C250 VTAIL.n165 B 0.026181f
C251 VTAIL.n166 B 0.052496f
C252 VTAIL.n167 B 0.011402f
C253 VTAIL.n168 B 0.011077f
C254 VTAIL.n169 B 0.049617f
C255 VTAIL.n170 B 0.029003f
C256 VTAIL.n171 B 0.88963f
C257 VTAIL.t7 B 0.128195f
C258 VTAIL.t5 B 0.128195f
C259 VTAIL.n172 B 1.0538f
C260 VTAIL.n173 B 0.330135f
C261 VTAIL.n174 B 0.026609f
C262 VTAIL.n175 B 0.020613f
C263 VTAIL.n176 B 0.011402f
C264 VTAIL.n177 B 0.026181f
C265 VTAIL.n178 B 0.011077f
C266 VTAIL.n179 B 0.011728f
C267 VTAIL.n180 B 0.020613f
C268 VTAIL.n181 B 0.011077f
C269 VTAIL.n182 B 0.026181f
C270 VTAIL.n183 B 0.011728f
C271 VTAIL.n184 B 0.020613f
C272 VTAIL.n185 B 0.011077f
C273 VTAIL.n186 B 0.019636f
C274 VTAIL.n187 B 0.018508f
C275 VTAIL.t3 B 0.043771f
C276 VTAIL.n188 B 0.115955f
C277 VTAIL.n189 B 0.661205f
C278 VTAIL.n190 B 0.011077f
C279 VTAIL.n191 B 0.011728f
C280 VTAIL.n192 B 0.026181f
C281 VTAIL.n193 B 0.026181f
C282 VTAIL.n194 B 0.011728f
C283 VTAIL.n195 B 0.011077f
C284 VTAIL.n196 B 0.020613f
C285 VTAIL.n197 B 0.020613f
C286 VTAIL.n198 B 0.011077f
C287 VTAIL.n199 B 0.011728f
C288 VTAIL.n200 B 0.026181f
C289 VTAIL.n201 B 0.026181f
C290 VTAIL.n202 B 0.011728f
C291 VTAIL.n203 B 0.011077f
C292 VTAIL.n204 B 0.020613f
C293 VTAIL.n205 B 0.020613f
C294 VTAIL.n206 B 0.011077f
C295 VTAIL.n207 B 0.011728f
C296 VTAIL.n208 B 0.026181f
C297 VTAIL.n209 B 0.026181f
C298 VTAIL.n210 B 0.052496f
C299 VTAIL.n211 B 0.011402f
C300 VTAIL.n212 B 0.011077f
C301 VTAIL.n213 B 0.049617f
C302 VTAIL.n214 B 0.029003f
C303 VTAIL.n215 B 0.11978f
C304 VTAIL.n216 B 0.026609f
C305 VTAIL.n217 B 0.020613f
C306 VTAIL.n218 B 0.011402f
C307 VTAIL.n219 B 0.026181f
C308 VTAIL.n220 B 0.011077f
C309 VTAIL.n221 B 0.011728f
C310 VTAIL.n222 B 0.020613f
C311 VTAIL.n223 B 0.011077f
C312 VTAIL.n224 B 0.026181f
C313 VTAIL.n225 B 0.011728f
C314 VTAIL.n226 B 0.020613f
C315 VTAIL.n227 B 0.011077f
C316 VTAIL.n228 B 0.019636f
C317 VTAIL.n229 B 0.018508f
C318 VTAIL.t8 B 0.043771f
C319 VTAIL.n230 B 0.115955f
C320 VTAIL.n231 B 0.661205f
C321 VTAIL.n232 B 0.011077f
C322 VTAIL.n233 B 0.011728f
C323 VTAIL.n234 B 0.026181f
C324 VTAIL.n235 B 0.026181f
C325 VTAIL.n236 B 0.011728f
C326 VTAIL.n237 B 0.011077f
C327 VTAIL.n238 B 0.020613f
C328 VTAIL.n239 B 0.020613f
C329 VTAIL.n240 B 0.011077f
C330 VTAIL.n241 B 0.011728f
C331 VTAIL.n242 B 0.026181f
C332 VTAIL.n243 B 0.026181f
C333 VTAIL.n244 B 0.011728f
C334 VTAIL.n245 B 0.011077f
C335 VTAIL.n246 B 0.020613f
C336 VTAIL.n247 B 0.020613f
C337 VTAIL.n248 B 0.011077f
C338 VTAIL.n249 B 0.011728f
C339 VTAIL.n250 B 0.026181f
C340 VTAIL.n251 B 0.026181f
C341 VTAIL.n252 B 0.052496f
C342 VTAIL.n253 B 0.011402f
C343 VTAIL.n254 B 0.011077f
C344 VTAIL.n255 B 0.049617f
C345 VTAIL.n256 B 0.029003f
C346 VTAIL.n257 B 0.11978f
C347 VTAIL.t10 B 0.128195f
C348 VTAIL.t13 B 0.128195f
C349 VTAIL.n258 B 1.0538f
C350 VTAIL.n259 B 0.330135f
C351 VTAIL.n260 B 0.026609f
C352 VTAIL.n261 B 0.020613f
C353 VTAIL.n262 B 0.011402f
C354 VTAIL.n263 B 0.026181f
C355 VTAIL.n264 B 0.011077f
C356 VTAIL.n265 B 0.011728f
C357 VTAIL.n266 B 0.020613f
C358 VTAIL.n267 B 0.011077f
C359 VTAIL.n268 B 0.026181f
C360 VTAIL.n269 B 0.011728f
C361 VTAIL.n270 B 0.020613f
C362 VTAIL.n271 B 0.011077f
C363 VTAIL.n272 B 0.019636f
C364 VTAIL.n273 B 0.018508f
C365 VTAIL.t12 B 0.043771f
C366 VTAIL.n274 B 0.115955f
C367 VTAIL.n275 B 0.661205f
C368 VTAIL.n276 B 0.011077f
C369 VTAIL.n277 B 0.011728f
C370 VTAIL.n278 B 0.026181f
C371 VTAIL.n279 B 0.026181f
C372 VTAIL.n280 B 0.011728f
C373 VTAIL.n281 B 0.011077f
C374 VTAIL.n282 B 0.020613f
C375 VTAIL.n283 B 0.020613f
C376 VTAIL.n284 B 0.011077f
C377 VTAIL.n285 B 0.011728f
C378 VTAIL.n286 B 0.026181f
C379 VTAIL.n287 B 0.026181f
C380 VTAIL.n288 B 0.011728f
C381 VTAIL.n289 B 0.011077f
C382 VTAIL.n290 B 0.020613f
C383 VTAIL.n291 B 0.020613f
C384 VTAIL.n292 B 0.011077f
C385 VTAIL.n293 B 0.011728f
C386 VTAIL.n294 B 0.026181f
C387 VTAIL.n295 B 0.026181f
C388 VTAIL.n296 B 0.052496f
C389 VTAIL.n297 B 0.011402f
C390 VTAIL.n298 B 0.011077f
C391 VTAIL.n299 B 0.049617f
C392 VTAIL.n300 B 0.029003f
C393 VTAIL.n301 B 0.88963f
C394 VTAIL.n302 B 0.026609f
C395 VTAIL.n303 B 0.020613f
C396 VTAIL.n304 B 0.011402f
C397 VTAIL.n305 B 0.026181f
C398 VTAIL.n306 B 0.011728f
C399 VTAIL.n307 B 0.020613f
C400 VTAIL.n308 B 0.011077f
C401 VTAIL.n309 B 0.026181f
C402 VTAIL.n310 B 0.011728f
C403 VTAIL.n311 B 0.020613f
C404 VTAIL.n312 B 0.011077f
C405 VTAIL.n313 B 0.019636f
C406 VTAIL.n314 B 0.018508f
C407 VTAIL.t6 B 0.043771f
C408 VTAIL.n315 B 0.115955f
C409 VTAIL.n316 B 0.661205f
C410 VTAIL.n317 B 0.011077f
C411 VTAIL.n318 B 0.011728f
C412 VTAIL.n319 B 0.026181f
C413 VTAIL.n320 B 0.026181f
C414 VTAIL.n321 B 0.011728f
C415 VTAIL.n322 B 0.011077f
C416 VTAIL.n323 B 0.020613f
C417 VTAIL.n324 B 0.020613f
C418 VTAIL.n325 B 0.011077f
C419 VTAIL.n326 B 0.011728f
C420 VTAIL.n327 B 0.026181f
C421 VTAIL.n328 B 0.026181f
C422 VTAIL.n329 B 0.011728f
C423 VTAIL.n330 B 0.011077f
C424 VTAIL.n331 B 0.020613f
C425 VTAIL.n332 B 0.020613f
C426 VTAIL.n333 B 0.011077f
C427 VTAIL.n334 B 0.011077f
C428 VTAIL.n335 B 0.011728f
C429 VTAIL.n336 B 0.026181f
C430 VTAIL.n337 B 0.026181f
C431 VTAIL.n338 B 0.052496f
C432 VTAIL.n339 B 0.011402f
C433 VTAIL.n340 B 0.011077f
C434 VTAIL.n341 B 0.049617f
C435 VTAIL.n342 B 0.029003f
C436 VTAIL.n343 B 0.885765f
C437 VP.n0 B 0.041496f
C438 VP.t2 B 0.779357f
C439 VP.n1 B 0.310086f
C440 VP.n2 B 0.041496f
C441 VP.t7 B 0.779357f
C442 VP.n3 B 0.019156f
C443 VP.n4 B 0.041496f
C444 VP.t0 B 0.836627f
C445 VP.t1 B 0.779357f
C446 VP.n5 B 0.310086f
C447 VP.n6 B 0.179136f
C448 VP.t6 B 0.779357f
C449 VP.t5 B 0.866675f
C450 VP.n7 B 0.353452f
C451 VP.n8 B 0.356721f
C452 VP.n9 B 0.050297f
C453 VP.n10 B 0.050297f
C454 VP.n11 B 0.041496f
C455 VP.n12 B 0.041496f
C456 VP.n13 B 0.054074f
C457 VP.n14 B 0.019156f
C458 VP.n15 B 0.355983f
C459 VP.n16 B 1.56557f
C460 VP.t4 B 0.836627f
C461 VP.n17 B 0.355983f
C462 VP.n18 B 1.60302f
C463 VP.n19 B 0.041496f
C464 VP.n20 B 0.041496f
C465 VP.n21 B 0.054074f
C466 VP.n22 B 0.310086f
C467 VP.n23 B 0.050297f
C468 VP.n24 B 0.050297f
C469 VP.n25 B 0.041496f
C470 VP.n26 B 0.041496f
C471 VP.n27 B 0.054074f
C472 VP.n28 B 0.019156f
C473 VP.t3 B 0.836627f
C474 VP.n29 B 0.355983f
C475 VP.n30 B 0.032158f
.ends

