* NGSPICE file created from diff_pair_sample_0044.ext - technology: sky130A

.subckt diff_pair_sample_0044 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VN.t0 VDD2.t0 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X1 VDD1.t9 VP.t0 VTAIL.t0 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=7.6206 ps=39.86 w=19.54 l=0.17
X2 VDD2.t4 VN.t1 VTAIL.t15 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X3 VTAIL.t14 VN.t2 VDD2.t3 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X4 VTAIL.t13 VN.t3 VDD2.t2 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X5 VDD2.t1 VN.t4 VTAIL.t12 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=3.2241 ps=19.87 w=19.54 l=0.17
X6 VDD1.t8 VP.t1 VTAIL.t3 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=3.2241 ps=19.87 w=19.54 l=0.17
X7 B.t11 B.t9 B.t10 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=0 ps=0 w=19.54 l=0.17
X8 VDD2.t6 VN.t5 VTAIL.t11 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=3.2241 ps=19.87 w=19.54 l=0.17
X9 VTAIL.t5 VP.t2 VDD1.t7 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X10 B.t8 B.t6 B.t7 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=0 ps=0 w=19.54 l=0.17
X11 VDD2.t5 VN.t6 VTAIL.t10 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=7.6206 ps=39.86 w=19.54 l=0.17
X12 B.t5 B.t3 B.t4 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=0 ps=0 w=19.54 l=0.17
X13 VTAIL.t9 VN.t7 VDD2.t9 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X14 VDD1.t6 VP.t3 VTAIL.t2 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=3.2241 ps=19.87 w=19.54 l=0.17
X15 VTAIL.t1 VP.t4 VDD1.t5 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X16 VDD1.t4 VP.t5 VTAIL.t18 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X17 VDD1.t3 VP.t6 VTAIL.t19 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X18 B.t2 B.t0 B.t1 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=7.6206 pd=39.86 as=0 ps=0 w=19.54 l=0.17
X19 VDD2.t8 VN.t8 VTAIL.t8 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X20 VTAIL.t17 VP.t7 VDD1.t2 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
X21 VDD2.t7 VN.t9 VTAIL.t7 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=7.6206 ps=39.86 w=19.54 l=0.17
X22 VDD1.t1 VP.t8 VTAIL.t6 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=7.6206 ps=39.86 w=19.54 l=0.17
X23 VTAIL.t4 VP.t9 VDD1.t0 w_n1570_n4876# sky130_fd_pr__pfet_01v8 ad=3.2241 pd=19.87 as=3.2241 ps=19.87 w=19.54 l=0.17
R0 VN.n8 VN.t9 2990.89
R1 VN.n2 VN.t5 2990.89
R2 VN.n18 VN.t4 2990.89
R3 VN.n12 VN.t6 2990.89
R4 VN.n7 VN.t0 2954.38
R5 VN.n5 VN.t1 2954.38
R6 VN.n1 VN.t3 2954.38
R7 VN.n17 VN.t7 2954.38
R8 VN.n15 VN.t8 2954.38
R9 VN.n11 VN.t2 2954.38
R10 VN.n13 VN.n12 161.489
R11 VN.n3 VN.n2 161.489
R12 VN.n9 VN.n8 161.3
R13 VN.n19 VN.n18 161.3
R14 VN.n16 VN.n10 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n6 VN.n0 161.3
R17 VN.n4 VN.n3 161.3
R18 VN VN.n19 46.01
R19 VN.n2 VN.n1 36.5157
R20 VN.n4 VN.n1 36.5157
R21 VN.n5 VN.n4 36.5157
R22 VN.n6 VN.n5 36.5157
R23 VN.n7 VN.n6 36.5157
R24 VN.n8 VN.n7 36.5157
R25 VN.n18 VN.n17 36.5157
R26 VN.n17 VN.n16 36.5157
R27 VN.n16 VN.n15 36.5157
R28 VN.n15 VN.n14 36.5157
R29 VN.n14 VN.n11 36.5157
R30 VN.n12 VN.n11 36.5157
R31 VN.n19 VN.n10 0.189894
R32 VN.n13 VN.n10 0.189894
R33 VN.n3 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VDD2.n210 VDD2.n209 585
R37 VDD2.n208 VDD2.n207 585
R38 VDD2.n113 VDD2.n112 585
R39 VDD2.n202 VDD2.n201 585
R40 VDD2.n200 VDD2.n199 585
R41 VDD2.n117 VDD2.n116 585
R42 VDD2.n194 VDD2.n193 585
R43 VDD2.n192 VDD2.n191 585
R44 VDD2.n121 VDD2.n120 585
R45 VDD2.n186 VDD2.n185 585
R46 VDD2.n184 VDD2.n183 585
R47 VDD2.n125 VDD2.n124 585
R48 VDD2.n178 VDD2.n177 585
R49 VDD2.n176 VDD2.n175 585
R50 VDD2.n129 VDD2.n128 585
R51 VDD2.n170 VDD2.n169 585
R52 VDD2.n168 VDD2.n167 585
R53 VDD2.n166 VDD2.n132 585
R54 VDD2.n136 VDD2.n133 585
R55 VDD2.n161 VDD2.n160 585
R56 VDD2.n159 VDD2.n158 585
R57 VDD2.n138 VDD2.n137 585
R58 VDD2.n153 VDD2.n152 585
R59 VDD2.n151 VDD2.n150 585
R60 VDD2.n142 VDD2.n141 585
R61 VDD2.n145 VDD2.n144 585
R62 VDD2.n35 VDD2.n34 585
R63 VDD2.n32 VDD2.n31 585
R64 VDD2.n41 VDD2.n40 585
R65 VDD2.n43 VDD2.n42 585
R66 VDD2.n28 VDD2.n27 585
R67 VDD2.n49 VDD2.n48 585
R68 VDD2.n52 VDD2.n51 585
R69 VDD2.n50 VDD2.n24 585
R70 VDD2.n57 VDD2.n23 585
R71 VDD2.n59 VDD2.n58 585
R72 VDD2.n61 VDD2.n60 585
R73 VDD2.n20 VDD2.n19 585
R74 VDD2.n67 VDD2.n66 585
R75 VDD2.n69 VDD2.n68 585
R76 VDD2.n16 VDD2.n15 585
R77 VDD2.n75 VDD2.n74 585
R78 VDD2.n77 VDD2.n76 585
R79 VDD2.n12 VDD2.n11 585
R80 VDD2.n83 VDD2.n82 585
R81 VDD2.n85 VDD2.n84 585
R82 VDD2.n8 VDD2.n7 585
R83 VDD2.n91 VDD2.n90 585
R84 VDD2.n93 VDD2.n92 585
R85 VDD2.n4 VDD2.n3 585
R86 VDD2.n99 VDD2.n98 585
R87 VDD2.n101 VDD2.n100 585
R88 VDD2.n209 VDD2.n109 498.474
R89 VDD2.n100 VDD2.n0 498.474
R90 VDD2.t1 VDD2.n143 329.036
R91 VDD2.t6 VDD2.n33 329.036
R92 VDD2.n209 VDD2.n208 171.744
R93 VDD2.n208 VDD2.n112 171.744
R94 VDD2.n201 VDD2.n112 171.744
R95 VDD2.n201 VDD2.n200 171.744
R96 VDD2.n200 VDD2.n116 171.744
R97 VDD2.n193 VDD2.n116 171.744
R98 VDD2.n193 VDD2.n192 171.744
R99 VDD2.n192 VDD2.n120 171.744
R100 VDD2.n185 VDD2.n120 171.744
R101 VDD2.n185 VDD2.n184 171.744
R102 VDD2.n184 VDD2.n124 171.744
R103 VDD2.n177 VDD2.n124 171.744
R104 VDD2.n177 VDD2.n176 171.744
R105 VDD2.n176 VDD2.n128 171.744
R106 VDD2.n169 VDD2.n128 171.744
R107 VDD2.n169 VDD2.n168 171.744
R108 VDD2.n168 VDD2.n132 171.744
R109 VDD2.n136 VDD2.n132 171.744
R110 VDD2.n160 VDD2.n136 171.744
R111 VDD2.n160 VDD2.n159 171.744
R112 VDD2.n159 VDD2.n137 171.744
R113 VDD2.n152 VDD2.n137 171.744
R114 VDD2.n152 VDD2.n151 171.744
R115 VDD2.n151 VDD2.n141 171.744
R116 VDD2.n144 VDD2.n141 171.744
R117 VDD2.n34 VDD2.n31 171.744
R118 VDD2.n41 VDD2.n31 171.744
R119 VDD2.n42 VDD2.n41 171.744
R120 VDD2.n42 VDD2.n27 171.744
R121 VDD2.n49 VDD2.n27 171.744
R122 VDD2.n51 VDD2.n49 171.744
R123 VDD2.n51 VDD2.n50 171.744
R124 VDD2.n50 VDD2.n23 171.744
R125 VDD2.n59 VDD2.n23 171.744
R126 VDD2.n60 VDD2.n59 171.744
R127 VDD2.n60 VDD2.n19 171.744
R128 VDD2.n67 VDD2.n19 171.744
R129 VDD2.n68 VDD2.n67 171.744
R130 VDD2.n68 VDD2.n15 171.744
R131 VDD2.n75 VDD2.n15 171.744
R132 VDD2.n76 VDD2.n75 171.744
R133 VDD2.n76 VDD2.n11 171.744
R134 VDD2.n83 VDD2.n11 171.744
R135 VDD2.n84 VDD2.n83 171.744
R136 VDD2.n84 VDD2.n7 171.744
R137 VDD2.n91 VDD2.n7 171.744
R138 VDD2.n92 VDD2.n91 171.744
R139 VDD2.n92 VDD2.n3 171.744
R140 VDD2.n99 VDD2.n3 171.744
R141 VDD2.n100 VDD2.n99 171.744
R142 VDD2.n144 VDD2.t1 85.8723
R143 VDD2.n34 VDD2.t6 85.8723
R144 VDD2.n108 VDD2.n107 72.3777
R145 VDD2 VDD2.n217 72.3748
R146 VDD2.n216 VDD2.n215 72.1099
R147 VDD2.n106 VDD2.n105 72.1098
R148 VDD2.n106 VDD2.n104 53.5618
R149 VDD2.n214 VDD2.n213 53.1308
R150 VDD2.n214 VDD2.n108 42.6075
R151 VDD2.n167 VDD2.n166 13.1884
R152 VDD2.n58 VDD2.n57 13.1884
R153 VDD2.n211 VDD2.n210 12.8005
R154 VDD2.n170 VDD2.n131 12.8005
R155 VDD2.n165 VDD2.n133 12.8005
R156 VDD2.n56 VDD2.n24 12.8005
R157 VDD2.n61 VDD2.n22 12.8005
R158 VDD2.n102 VDD2.n101 12.8005
R159 VDD2.n207 VDD2.n111 12.0247
R160 VDD2.n171 VDD2.n129 12.0247
R161 VDD2.n162 VDD2.n161 12.0247
R162 VDD2.n53 VDD2.n52 12.0247
R163 VDD2.n62 VDD2.n20 12.0247
R164 VDD2.n98 VDD2.n2 12.0247
R165 VDD2.n206 VDD2.n113 11.249
R166 VDD2.n175 VDD2.n174 11.249
R167 VDD2.n158 VDD2.n135 11.249
R168 VDD2.n48 VDD2.n26 11.249
R169 VDD2.n66 VDD2.n65 11.249
R170 VDD2.n97 VDD2.n4 11.249
R171 VDD2.n145 VDD2.n143 10.7239
R172 VDD2.n35 VDD2.n33 10.7239
R173 VDD2.n203 VDD2.n202 10.4732
R174 VDD2.n178 VDD2.n127 10.4732
R175 VDD2.n157 VDD2.n138 10.4732
R176 VDD2.n47 VDD2.n28 10.4732
R177 VDD2.n69 VDD2.n18 10.4732
R178 VDD2.n94 VDD2.n93 10.4732
R179 VDD2.n199 VDD2.n115 9.69747
R180 VDD2.n179 VDD2.n125 9.69747
R181 VDD2.n154 VDD2.n153 9.69747
R182 VDD2.n44 VDD2.n43 9.69747
R183 VDD2.n70 VDD2.n16 9.69747
R184 VDD2.n90 VDD2.n6 9.69747
R185 VDD2.n213 VDD2.n212 9.45567
R186 VDD2.n104 VDD2.n103 9.45567
R187 VDD2.n147 VDD2.n146 9.3005
R188 VDD2.n149 VDD2.n148 9.3005
R189 VDD2.n140 VDD2.n139 9.3005
R190 VDD2.n155 VDD2.n154 9.3005
R191 VDD2.n157 VDD2.n156 9.3005
R192 VDD2.n135 VDD2.n134 9.3005
R193 VDD2.n163 VDD2.n162 9.3005
R194 VDD2.n165 VDD2.n164 9.3005
R195 VDD2.n119 VDD2.n118 9.3005
R196 VDD2.n196 VDD2.n195 9.3005
R197 VDD2.n198 VDD2.n197 9.3005
R198 VDD2.n115 VDD2.n114 9.3005
R199 VDD2.n204 VDD2.n203 9.3005
R200 VDD2.n206 VDD2.n205 9.3005
R201 VDD2.n111 VDD2.n110 9.3005
R202 VDD2.n212 VDD2.n211 9.3005
R203 VDD2.n190 VDD2.n189 9.3005
R204 VDD2.n188 VDD2.n187 9.3005
R205 VDD2.n123 VDD2.n122 9.3005
R206 VDD2.n182 VDD2.n181 9.3005
R207 VDD2.n180 VDD2.n179 9.3005
R208 VDD2.n127 VDD2.n126 9.3005
R209 VDD2.n174 VDD2.n173 9.3005
R210 VDD2.n172 VDD2.n171 9.3005
R211 VDD2.n131 VDD2.n130 9.3005
R212 VDD2.n79 VDD2.n78 9.3005
R213 VDD2.n14 VDD2.n13 9.3005
R214 VDD2.n73 VDD2.n72 9.3005
R215 VDD2.n71 VDD2.n70 9.3005
R216 VDD2.n18 VDD2.n17 9.3005
R217 VDD2.n65 VDD2.n64 9.3005
R218 VDD2.n63 VDD2.n62 9.3005
R219 VDD2.n22 VDD2.n21 9.3005
R220 VDD2.n37 VDD2.n36 9.3005
R221 VDD2.n39 VDD2.n38 9.3005
R222 VDD2.n30 VDD2.n29 9.3005
R223 VDD2.n45 VDD2.n44 9.3005
R224 VDD2.n47 VDD2.n46 9.3005
R225 VDD2.n26 VDD2.n25 9.3005
R226 VDD2.n54 VDD2.n53 9.3005
R227 VDD2.n56 VDD2.n55 9.3005
R228 VDD2.n81 VDD2.n80 9.3005
R229 VDD2.n10 VDD2.n9 9.3005
R230 VDD2.n87 VDD2.n86 9.3005
R231 VDD2.n89 VDD2.n88 9.3005
R232 VDD2.n6 VDD2.n5 9.3005
R233 VDD2.n95 VDD2.n94 9.3005
R234 VDD2.n97 VDD2.n96 9.3005
R235 VDD2.n2 VDD2.n1 9.3005
R236 VDD2.n103 VDD2.n102 9.3005
R237 VDD2.n198 VDD2.n117 8.92171
R238 VDD2.n183 VDD2.n182 8.92171
R239 VDD2.n150 VDD2.n140 8.92171
R240 VDD2.n40 VDD2.n30 8.92171
R241 VDD2.n74 VDD2.n73 8.92171
R242 VDD2.n89 VDD2.n8 8.92171
R243 VDD2.n195 VDD2.n194 8.14595
R244 VDD2.n186 VDD2.n123 8.14595
R245 VDD2.n149 VDD2.n142 8.14595
R246 VDD2.n39 VDD2.n32 8.14595
R247 VDD2.n77 VDD2.n14 8.14595
R248 VDD2.n86 VDD2.n85 8.14595
R249 VDD2.n213 VDD2.n109 7.75445
R250 VDD2.n104 VDD2.n0 7.75445
R251 VDD2.n191 VDD2.n119 7.3702
R252 VDD2.n187 VDD2.n121 7.3702
R253 VDD2.n146 VDD2.n145 7.3702
R254 VDD2.n36 VDD2.n35 7.3702
R255 VDD2.n78 VDD2.n12 7.3702
R256 VDD2.n82 VDD2.n10 7.3702
R257 VDD2.n191 VDD2.n190 6.59444
R258 VDD2.n190 VDD2.n121 6.59444
R259 VDD2.n81 VDD2.n12 6.59444
R260 VDD2.n82 VDD2.n81 6.59444
R261 VDD2.n211 VDD2.n109 6.08283
R262 VDD2.n102 VDD2.n0 6.08283
R263 VDD2.n194 VDD2.n119 5.81868
R264 VDD2.n187 VDD2.n186 5.81868
R265 VDD2.n146 VDD2.n142 5.81868
R266 VDD2.n36 VDD2.n32 5.81868
R267 VDD2.n78 VDD2.n77 5.81868
R268 VDD2.n85 VDD2.n10 5.81868
R269 VDD2.n195 VDD2.n117 5.04292
R270 VDD2.n183 VDD2.n123 5.04292
R271 VDD2.n150 VDD2.n149 5.04292
R272 VDD2.n40 VDD2.n39 5.04292
R273 VDD2.n74 VDD2.n14 5.04292
R274 VDD2.n86 VDD2.n8 5.04292
R275 VDD2.n199 VDD2.n198 4.26717
R276 VDD2.n182 VDD2.n125 4.26717
R277 VDD2.n153 VDD2.n140 4.26717
R278 VDD2.n43 VDD2.n30 4.26717
R279 VDD2.n73 VDD2.n16 4.26717
R280 VDD2.n90 VDD2.n89 4.26717
R281 VDD2.n202 VDD2.n115 3.49141
R282 VDD2.n179 VDD2.n178 3.49141
R283 VDD2.n154 VDD2.n138 3.49141
R284 VDD2.n44 VDD2.n28 3.49141
R285 VDD2.n70 VDD2.n69 3.49141
R286 VDD2.n93 VDD2.n6 3.49141
R287 VDD2.n203 VDD2.n113 2.71565
R288 VDD2.n175 VDD2.n127 2.71565
R289 VDD2.n158 VDD2.n157 2.71565
R290 VDD2.n48 VDD2.n47 2.71565
R291 VDD2.n66 VDD2.n18 2.71565
R292 VDD2.n94 VDD2.n4 2.71565
R293 VDD2.n147 VDD2.n143 2.41282
R294 VDD2.n37 VDD2.n33 2.41282
R295 VDD2.n207 VDD2.n206 1.93989
R296 VDD2.n174 VDD2.n129 1.93989
R297 VDD2.n161 VDD2.n135 1.93989
R298 VDD2.n52 VDD2.n26 1.93989
R299 VDD2.n65 VDD2.n20 1.93989
R300 VDD2.n98 VDD2.n97 1.93989
R301 VDD2.n217 VDD2.t3 1.66401
R302 VDD2.n217 VDD2.t5 1.66401
R303 VDD2.n215 VDD2.t9 1.66401
R304 VDD2.n215 VDD2.t8 1.66401
R305 VDD2.n107 VDD2.t0 1.66401
R306 VDD2.n107 VDD2.t7 1.66401
R307 VDD2.n105 VDD2.t2 1.66401
R308 VDD2.n105 VDD2.t4 1.66401
R309 VDD2.n210 VDD2.n111 1.16414
R310 VDD2.n171 VDD2.n170 1.16414
R311 VDD2.n162 VDD2.n133 1.16414
R312 VDD2.n53 VDD2.n24 1.16414
R313 VDD2.n62 VDD2.n61 1.16414
R314 VDD2.n101 VDD2.n2 1.16414
R315 VDD2.n216 VDD2.n214 0.431534
R316 VDD2.n167 VDD2.n131 0.388379
R317 VDD2.n166 VDD2.n165 0.388379
R318 VDD2.n57 VDD2.n56 0.388379
R319 VDD2.n58 VDD2.n22 0.388379
R320 VDD2 VDD2.n216 0.166448
R321 VDD2.n212 VDD2.n110 0.155672
R322 VDD2.n205 VDD2.n110 0.155672
R323 VDD2.n205 VDD2.n204 0.155672
R324 VDD2.n204 VDD2.n114 0.155672
R325 VDD2.n197 VDD2.n114 0.155672
R326 VDD2.n197 VDD2.n196 0.155672
R327 VDD2.n196 VDD2.n118 0.155672
R328 VDD2.n189 VDD2.n118 0.155672
R329 VDD2.n189 VDD2.n188 0.155672
R330 VDD2.n188 VDD2.n122 0.155672
R331 VDD2.n181 VDD2.n122 0.155672
R332 VDD2.n181 VDD2.n180 0.155672
R333 VDD2.n180 VDD2.n126 0.155672
R334 VDD2.n173 VDD2.n126 0.155672
R335 VDD2.n173 VDD2.n172 0.155672
R336 VDD2.n172 VDD2.n130 0.155672
R337 VDD2.n164 VDD2.n130 0.155672
R338 VDD2.n164 VDD2.n163 0.155672
R339 VDD2.n163 VDD2.n134 0.155672
R340 VDD2.n156 VDD2.n134 0.155672
R341 VDD2.n156 VDD2.n155 0.155672
R342 VDD2.n155 VDD2.n139 0.155672
R343 VDD2.n148 VDD2.n139 0.155672
R344 VDD2.n148 VDD2.n147 0.155672
R345 VDD2.n38 VDD2.n37 0.155672
R346 VDD2.n38 VDD2.n29 0.155672
R347 VDD2.n45 VDD2.n29 0.155672
R348 VDD2.n46 VDD2.n45 0.155672
R349 VDD2.n46 VDD2.n25 0.155672
R350 VDD2.n54 VDD2.n25 0.155672
R351 VDD2.n55 VDD2.n54 0.155672
R352 VDD2.n55 VDD2.n21 0.155672
R353 VDD2.n63 VDD2.n21 0.155672
R354 VDD2.n64 VDD2.n63 0.155672
R355 VDD2.n64 VDD2.n17 0.155672
R356 VDD2.n71 VDD2.n17 0.155672
R357 VDD2.n72 VDD2.n71 0.155672
R358 VDD2.n72 VDD2.n13 0.155672
R359 VDD2.n79 VDD2.n13 0.155672
R360 VDD2.n80 VDD2.n79 0.155672
R361 VDD2.n80 VDD2.n9 0.155672
R362 VDD2.n87 VDD2.n9 0.155672
R363 VDD2.n88 VDD2.n87 0.155672
R364 VDD2.n88 VDD2.n5 0.155672
R365 VDD2.n95 VDD2.n5 0.155672
R366 VDD2.n96 VDD2.n95 0.155672
R367 VDD2.n96 VDD2.n1 0.155672
R368 VDD2.n103 VDD2.n1 0.155672
R369 VDD2.n108 VDD2.n106 0.0529126
R370 VTAIL.n367 VTAIL.n366 585
R371 VTAIL.n364 VTAIL.n363 585
R372 VTAIL.n373 VTAIL.n372 585
R373 VTAIL.n375 VTAIL.n374 585
R374 VTAIL.n360 VTAIL.n359 585
R375 VTAIL.n381 VTAIL.n380 585
R376 VTAIL.n384 VTAIL.n383 585
R377 VTAIL.n382 VTAIL.n356 585
R378 VTAIL.n389 VTAIL.n355 585
R379 VTAIL.n391 VTAIL.n390 585
R380 VTAIL.n393 VTAIL.n392 585
R381 VTAIL.n352 VTAIL.n351 585
R382 VTAIL.n399 VTAIL.n398 585
R383 VTAIL.n401 VTAIL.n400 585
R384 VTAIL.n348 VTAIL.n347 585
R385 VTAIL.n407 VTAIL.n406 585
R386 VTAIL.n409 VTAIL.n408 585
R387 VTAIL.n344 VTAIL.n343 585
R388 VTAIL.n415 VTAIL.n414 585
R389 VTAIL.n417 VTAIL.n416 585
R390 VTAIL.n340 VTAIL.n339 585
R391 VTAIL.n423 VTAIL.n422 585
R392 VTAIL.n425 VTAIL.n424 585
R393 VTAIL.n336 VTAIL.n335 585
R394 VTAIL.n431 VTAIL.n430 585
R395 VTAIL.n433 VTAIL.n432 585
R396 VTAIL.n37 VTAIL.n36 585
R397 VTAIL.n34 VTAIL.n33 585
R398 VTAIL.n43 VTAIL.n42 585
R399 VTAIL.n45 VTAIL.n44 585
R400 VTAIL.n30 VTAIL.n29 585
R401 VTAIL.n51 VTAIL.n50 585
R402 VTAIL.n54 VTAIL.n53 585
R403 VTAIL.n52 VTAIL.n26 585
R404 VTAIL.n59 VTAIL.n25 585
R405 VTAIL.n61 VTAIL.n60 585
R406 VTAIL.n63 VTAIL.n62 585
R407 VTAIL.n22 VTAIL.n21 585
R408 VTAIL.n69 VTAIL.n68 585
R409 VTAIL.n71 VTAIL.n70 585
R410 VTAIL.n18 VTAIL.n17 585
R411 VTAIL.n77 VTAIL.n76 585
R412 VTAIL.n79 VTAIL.n78 585
R413 VTAIL.n14 VTAIL.n13 585
R414 VTAIL.n85 VTAIL.n84 585
R415 VTAIL.n87 VTAIL.n86 585
R416 VTAIL.n10 VTAIL.n9 585
R417 VTAIL.n93 VTAIL.n92 585
R418 VTAIL.n95 VTAIL.n94 585
R419 VTAIL.n6 VTAIL.n5 585
R420 VTAIL.n101 VTAIL.n100 585
R421 VTAIL.n103 VTAIL.n102 585
R422 VTAIL.n327 VTAIL.n326 585
R423 VTAIL.n325 VTAIL.n324 585
R424 VTAIL.n230 VTAIL.n229 585
R425 VTAIL.n319 VTAIL.n318 585
R426 VTAIL.n317 VTAIL.n316 585
R427 VTAIL.n234 VTAIL.n233 585
R428 VTAIL.n311 VTAIL.n310 585
R429 VTAIL.n309 VTAIL.n308 585
R430 VTAIL.n238 VTAIL.n237 585
R431 VTAIL.n303 VTAIL.n302 585
R432 VTAIL.n301 VTAIL.n300 585
R433 VTAIL.n242 VTAIL.n241 585
R434 VTAIL.n295 VTAIL.n294 585
R435 VTAIL.n293 VTAIL.n292 585
R436 VTAIL.n246 VTAIL.n245 585
R437 VTAIL.n287 VTAIL.n286 585
R438 VTAIL.n285 VTAIL.n284 585
R439 VTAIL.n283 VTAIL.n249 585
R440 VTAIL.n253 VTAIL.n250 585
R441 VTAIL.n278 VTAIL.n277 585
R442 VTAIL.n276 VTAIL.n275 585
R443 VTAIL.n255 VTAIL.n254 585
R444 VTAIL.n270 VTAIL.n269 585
R445 VTAIL.n268 VTAIL.n267 585
R446 VTAIL.n259 VTAIL.n258 585
R447 VTAIL.n262 VTAIL.n261 585
R448 VTAIL.n217 VTAIL.n216 585
R449 VTAIL.n215 VTAIL.n214 585
R450 VTAIL.n120 VTAIL.n119 585
R451 VTAIL.n209 VTAIL.n208 585
R452 VTAIL.n207 VTAIL.n206 585
R453 VTAIL.n124 VTAIL.n123 585
R454 VTAIL.n201 VTAIL.n200 585
R455 VTAIL.n199 VTAIL.n198 585
R456 VTAIL.n128 VTAIL.n127 585
R457 VTAIL.n193 VTAIL.n192 585
R458 VTAIL.n191 VTAIL.n190 585
R459 VTAIL.n132 VTAIL.n131 585
R460 VTAIL.n185 VTAIL.n184 585
R461 VTAIL.n183 VTAIL.n182 585
R462 VTAIL.n136 VTAIL.n135 585
R463 VTAIL.n177 VTAIL.n176 585
R464 VTAIL.n175 VTAIL.n174 585
R465 VTAIL.n173 VTAIL.n139 585
R466 VTAIL.n143 VTAIL.n140 585
R467 VTAIL.n168 VTAIL.n167 585
R468 VTAIL.n166 VTAIL.n165 585
R469 VTAIL.n145 VTAIL.n144 585
R470 VTAIL.n160 VTAIL.n159 585
R471 VTAIL.n158 VTAIL.n157 585
R472 VTAIL.n149 VTAIL.n148 585
R473 VTAIL.n152 VTAIL.n151 585
R474 VTAIL.n432 VTAIL.n332 498.474
R475 VTAIL.n102 VTAIL.n2 498.474
R476 VTAIL.n326 VTAIL.n226 498.474
R477 VTAIL.n216 VTAIL.n116 498.474
R478 VTAIL.t7 VTAIL.n365 329.036
R479 VTAIL.t6 VTAIL.n35 329.036
R480 VTAIL.t0 VTAIL.n260 329.036
R481 VTAIL.t10 VTAIL.n150 329.036
R482 VTAIL.n366 VTAIL.n363 171.744
R483 VTAIL.n373 VTAIL.n363 171.744
R484 VTAIL.n374 VTAIL.n373 171.744
R485 VTAIL.n374 VTAIL.n359 171.744
R486 VTAIL.n381 VTAIL.n359 171.744
R487 VTAIL.n383 VTAIL.n381 171.744
R488 VTAIL.n383 VTAIL.n382 171.744
R489 VTAIL.n382 VTAIL.n355 171.744
R490 VTAIL.n391 VTAIL.n355 171.744
R491 VTAIL.n392 VTAIL.n391 171.744
R492 VTAIL.n392 VTAIL.n351 171.744
R493 VTAIL.n399 VTAIL.n351 171.744
R494 VTAIL.n400 VTAIL.n399 171.744
R495 VTAIL.n400 VTAIL.n347 171.744
R496 VTAIL.n407 VTAIL.n347 171.744
R497 VTAIL.n408 VTAIL.n407 171.744
R498 VTAIL.n408 VTAIL.n343 171.744
R499 VTAIL.n415 VTAIL.n343 171.744
R500 VTAIL.n416 VTAIL.n415 171.744
R501 VTAIL.n416 VTAIL.n339 171.744
R502 VTAIL.n423 VTAIL.n339 171.744
R503 VTAIL.n424 VTAIL.n423 171.744
R504 VTAIL.n424 VTAIL.n335 171.744
R505 VTAIL.n431 VTAIL.n335 171.744
R506 VTAIL.n432 VTAIL.n431 171.744
R507 VTAIL.n36 VTAIL.n33 171.744
R508 VTAIL.n43 VTAIL.n33 171.744
R509 VTAIL.n44 VTAIL.n43 171.744
R510 VTAIL.n44 VTAIL.n29 171.744
R511 VTAIL.n51 VTAIL.n29 171.744
R512 VTAIL.n53 VTAIL.n51 171.744
R513 VTAIL.n53 VTAIL.n52 171.744
R514 VTAIL.n52 VTAIL.n25 171.744
R515 VTAIL.n61 VTAIL.n25 171.744
R516 VTAIL.n62 VTAIL.n61 171.744
R517 VTAIL.n62 VTAIL.n21 171.744
R518 VTAIL.n69 VTAIL.n21 171.744
R519 VTAIL.n70 VTAIL.n69 171.744
R520 VTAIL.n70 VTAIL.n17 171.744
R521 VTAIL.n77 VTAIL.n17 171.744
R522 VTAIL.n78 VTAIL.n77 171.744
R523 VTAIL.n78 VTAIL.n13 171.744
R524 VTAIL.n85 VTAIL.n13 171.744
R525 VTAIL.n86 VTAIL.n85 171.744
R526 VTAIL.n86 VTAIL.n9 171.744
R527 VTAIL.n93 VTAIL.n9 171.744
R528 VTAIL.n94 VTAIL.n93 171.744
R529 VTAIL.n94 VTAIL.n5 171.744
R530 VTAIL.n101 VTAIL.n5 171.744
R531 VTAIL.n102 VTAIL.n101 171.744
R532 VTAIL.n326 VTAIL.n325 171.744
R533 VTAIL.n325 VTAIL.n229 171.744
R534 VTAIL.n318 VTAIL.n229 171.744
R535 VTAIL.n318 VTAIL.n317 171.744
R536 VTAIL.n317 VTAIL.n233 171.744
R537 VTAIL.n310 VTAIL.n233 171.744
R538 VTAIL.n310 VTAIL.n309 171.744
R539 VTAIL.n309 VTAIL.n237 171.744
R540 VTAIL.n302 VTAIL.n237 171.744
R541 VTAIL.n302 VTAIL.n301 171.744
R542 VTAIL.n301 VTAIL.n241 171.744
R543 VTAIL.n294 VTAIL.n241 171.744
R544 VTAIL.n294 VTAIL.n293 171.744
R545 VTAIL.n293 VTAIL.n245 171.744
R546 VTAIL.n286 VTAIL.n245 171.744
R547 VTAIL.n286 VTAIL.n285 171.744
R548 VTAIL.n285 VTAIL.n249 171.744
R549 VTAIL.n253 VTAIL.n249 171.744
R550 VTAIL.n277 VTAIL.n253 171.744
R551 VTAIL.n277 VTAIL.n276 171.744
R552 VTAIL.n276 VTAIL.n254 171.744
R553 VTAIL.n269 VTAIL.n254 171.744
R554 VTAIL.n269 VTAIL.n268 171.744
R555 VTAIL.n268 VTAIL.n258 171.744
R556 VTAIL.n261 VTAIL.n258 171.744
R557 VTAIL.n216 VTAIL.n215 171.744
R558 VTAIL.n215 VTAIL.n119 171.744
R559 VTAIL.n208 VTAIL.n119 171.744
R560 VTAIL.n208 VTAIL.n207 171.744
R561 VTAIL.n207 VTAIL.n123 171.744
R562 VTAIL.n200 VTAIL.n123 171.744
R563 VTAIL.n200 VTAIL.n199 171.744
R564 VTAIL.n199 VTAIL.n127 171.744
R565 VTAIL.n192 VTAIL.n127 171.744
R566 VTAIL.n192 VTAIL.n191 171.744
R567 VTAIL.n191 VTAIL.n131 171.744
R568 VTAIL.n184 VTAIL.n131 171.744
R569 VTAIL.n184 VTAIL.n183 171.744
R570 VTAIL.n183 VTAIL.n135 171.744
R571 VTAIL.n176 VTAIL.n135 171.744
R572 VTAIL.n176 VTAIL.n175 171.744
R573 VTAIL.n175 VTAIL.n139 171.744
R574 VTAIL.n143 VTAIL.n139 171.744
R575 VTAIL.n167 VTAIL.n143 171.744
R576 VTAIL.n167 VTAIL.n166 171.744
R577 VTAIL.n166 VTAIL.n144 171.744
R578 VTAIL.n159 VTAIL.n144 171.744
R579 VTAIL.n159 VTAIL.n158 171.744
R580 VTAIL.n158 VTAIL.n148 171.744
R581 VTAIL.n151 VTAIL.n148 171.744
R582 VTAIL.n366 VTAIL.t7 85.8723
R583 VTAIL.n36 VTAIL.t6 85.8723
R584 VTAIL.n261 VTAIL.t0 85.8723
R585 VTAIL.n151 VTAIL.t10 85.8723
R586 VTAIL.n225 VTAIL.n224 55.4311
R587 VTAIL.n223 VTAIL.n222 55.4311
R588 VTAIL.n115 VTAIL.n114 55.4311
R589 VTAIL.n113 VTAIL.n112 55.4311
R590 VTAIL.n439 VTAIL.n438 55.431
R591 VTAIL.n1 VTAIL.n0 55.431
R592 VTAIL.n109 VTAIL.n108 55.431
R593 VTAIL.n111 VTAIL.n110 55.431
R594 VTAIL.n437 VTAIL.n436 36.452
R595 VTAIL.n107 VTAIL.n106 36.452
R596 VTAIL.n331 VTAIL.n330 36.452
R597 VTAIL.n221 VTAIL.n220 36.452
R598 VTAIL.n113 VTAIL.n111 30.0738
R599 VTAIL.n437 VTAIL.n331 29.6427
R600 VTAIL.n390 VTAIL.n389 13.1884
R601 VTAIL.n60 VTAIL.n59 13.1884
R602 VTAIL.n284 VTAIL.n283 13.1884
R603 VTAIL.n174 VTAIL.n173 13.1884
R604 VTAIL.n388 VTAIL.n356 12.8005
R605 VTAIL.n393 VTAIL.n354 12.8005
R606 VTAIL.n434 VTAIL.n433 12.8005
R607 VTAIL.n58 VTAIL.n26 12.8005
R608 VTAIL.n63 VTAIL.n24 12.8005
R609 VTAIL.n104 VTAIL.n103 12.8005
R610 VTAIL.n328 VTAIL.n327 12.8005
R611 VTAIL.n287 VTAIL.n248 12.8005
R612 VTAIL.n282 VTAIL.n250 12.8005
R613 VTAIL.n218 VTAIL.n217 12.8005
R614 VTAIL.n177 VTAIL.n138 12.8005
R615 VTAIL.n172 VTAIL.n140 12.8005
R616 VTAIL.n385 VTAIL.n384 12.0247
R617 VTAIL.n394 VTAIL.n352 12.0247
R618 VTAIL.n430 VTAIL.n334 12.0247
R619 VTAIL.n55 VTAIL.n54 12.0247
R620 VTAIL.n64 VTAIL.n22 12.0247
R621 VTAIL.n100 VTAIL.n4 12.0247
R622 VTAIL.n324 VTAIL.n228 12.0247
R623 VTAIL.n288 VTAIL.n246 12.0247
R624 VTAIL.n279 VTAIL.n278 12.0247
R625 VTAIL.n214 VTAIL.n118 12.0247
R626 VTAIL.n178 VTAIL.n136 12.0247
R627 VTAIL.n169 VTAIL.n168 12.0247
R628 VTAIL.n380 VTAIL.n358 11.249
R629 VTAIL.n398 VTAIL.n397 11.249
R630 VTAIL.n429 VTAIL.n336 11.249
R631 VTAIL.n50 VTAIL.n28 11.249
R632 VTAIL.n68 VTAIL.n67 11.249
R633 VTAIL.n99 VTAIL.n6 11.249
R634 VTAIL.n323 VTAIL.n230 11.249
R635 VTAIL.n292 VTAIL.n291 11.249
R636 VTAIL.n275 VTAIL.n252 11.249
R637 VTAIL.n213 VTAIL.n120 11.249
R638 VTAIL.n182 VTAIL.n181 11.249
R639 VTAIL.n165 VTAIL.n142 11.249
R640 VTAIL.n367 VTAIL.n365 10.7239
R641 VTAIL.n37 VTAIL.n35 10.7239
R642 VTAIL.n262 VTAIL.n260 10.7239
R643 VTAIL.n152 VTAIL.n150 10.7239
R644 VTAIL.n379 VTAIL.n360 10.4732
R645 VTAIL.n401 VTAIL.n350 10.4732
R646 VTAIL.n426 VTAIL.n425 10.4732
R647 VTAIL.n49 VTAIL.n30 10.4732
R648 VTAIL.n71 VTAIL.n20 10.4732
R649 VTAIL.n96 VTAIL.n95 10.4732
R650 VTAIL.n320 VTAIL.n319 10.4732
R651 VTAIL.n295 VTAIL.n244 10.4732
R652 VTAIL.n274 VTAIL.n255 10.4732
R653 VTAIL.n210 VTAIL.n209 10.4732
R654 VTAIL.n185 VTAIL.n134 10.4732
R655 VTAIL.n164 VTAIL.n145 10.4732
R656 VTAIL.n376 VTAIL.n375 9.69747
R657 VTAIL.n402 VTAIL.n348 9.69747
R658 VTAIL.n422 VTAIL.n338 9.69747
R659 VTAIL.n46 VTAIL.n45 9.69747
R660 VTAIL.n72 VTAIL.n18 9.69747
R661 VTAIL.n92 VTAIL.n8 9.69747
R662 VTAIL.n316 VTAIL.n232 9.69747
R663 VTAIL.n296 VTAIL.n242 9.69747
R664 VTAIL.n271 VTAIL.n270 9.69747
R665 VTAIL.n206 VTAIL.n122 9.69747
R666 VTAIL.n186 VTAIL.n132 9.69747
R667 VTAIL.n161 VTAIL.n160 9.69747
R668 VTAIL.n436 VTAIL.n435 9.45567
R669 VTAIL.n106 VTAIL.n105 9.45567
R670 VTAIL.n330 VTAIL.n329 9.45567
R671 VTAIL.n220 VTAIL.n219 9.45567
R672 VTAIL.n411 VTAIL.n410 9.3005
R673 VTAIL.n346 VTAIL.n345 9.3005
R674 VTAIL.n405 VTAIL.n404 9.3005
R675 VTAIL.n403 VTAIL.n402 9.3005
R676 VTAIL.n350 VTAIL.n349 9.3005
R677 VTAIL.n397 VTAIL.n396 9.3005
R678 VTAIL.n395 VTAIL.n394 9.3005
R679 VTAIL.n354 VTAIL.n353 9.3005
R680 VTAIL.n369 VTAIL.n368 9.3005
R681 VTAIL.n371 VTAIL.n370 9.3005
R682 VTAIL.n362 VTAIL.n361 9.3005
R683 VTAIL.n377 VTAIL.n376 9.3005
R684 VTAIL.n379 VTAIL.n378 9.3005
R685 VTAIL.n358 VTAIL.n357 9.3005
R686 VTAIL.n386 VTAIL.n385 9.3005
R687 VTAIL.n388 VTAIL.n387 9.3005
R688 VTAIL.n413 VTAIL.n412 9.3005
R689 VTAIL.n342 VTAIL.n341 9.3005
R690 VTAIL.n419 VTAIL.n418 9.3005
R691 VTAIL.n421 VTAIL.n420 9.3005
R692 VTAIL.n338 VTAIL.n337 9.3005
R693 VTAIL.n427 VTAIL.n426 9.3005
R694 VTAIL.n429 VTAIL.n428 9.3005
R695 VTAIL.n334 VTAIL.n333 9.3005
R696 VTAIL.n435 VTAIL.n434 9.3005
R697 VTAIL.n81 VTAIL.n80 9.3005
R698 VTAIL.n16 VTAIL.n15 9.3005
R699 VTAIL.n75 VTAIL.n74 9.3005
R700 VTAIL.n73 VTAIL.n72 9.3005
R701 VTAIL.n20 VTAIL.n19 9.3005
R702 VTAIL.n67 VTAIL.n66 9.3005
R703 VTAIL.n65 VTAIL.n64 9.3005
R704 VTAIL.n24 VTAIL.n23 9.3005
R705 VTAIL.n39 VTAIL.n38 9.3005
R706 VTAIL.n41 VTAIL.n40 9.3005
R707 VTAIL.n32 VTAIL.n31 9.3005
R708 VTAIL.n47 VTAIL.n46 9.3005
R709 VTAIL.n49 VTAIL.n48 9.3005
R710 VTAIL.n28 VTAIL.n27 9.3005
R711 VTAIL.n56 VTAIL.n55 9.3005
R712 VTAIL.n58 VTAIL.n57 9.3005
R713 VTAIL.n83 VTAIL.n82 9.3005
R714 VTAIL.n12 VTAIL.n11 9.3005
R715 VTAIL.n89 VTAIL.n88 9.3005
R716 VTAIL.n91 VTAIL.n90 9.3005
R717 VTAIL.n8 VTAIL.n7 9.3005
R718 VTAIL.n97 VTAIL.n96 9.3005
R719 VTAIL.n99 VTAIL.n98 9.3005
R720 VTAIL.n4 VTAIL.n3 9.3005
R721 VTAIL.n105 VTAIL.n104 9.3005
R722 VTAIL.n264 VTAIL.n263 9.3005
R723 VTAIL.n266 VTAIL.n265 9.3005
R724 VTAIL.n257 VTAIL.n256 9.3005
R725 VTAIL.n272 VTAIL.n271 9.3005
R726 VTAIL.n274 VTAIL.n273 9.3005
R727 VTAIL.n252 VTAIL.n251 9.3005
R728 VTAIL.n280 VTAIL.n279 9.3005
R729 VTAIL.n282 VTAIL.n281 9.3005
R730 VTAIL.n236 VTAIL.n235 9.3005
R731 VTAIL.n313 VTAIL.n312 9.3005
R732 VTAIL.n315 VTAIL.n314 9.3005
R733 VTAIL.n232 VTAIL.n231 9.3005
R734 VTAIL.n321 VTAIL.n320 9.3005
R735 VTAIL.n323 VTAIL.n322 9.3005
R736 VTAIL.n228 VTAIL.n227 9.3005
R737 VTAIL.n329 VTAIL.n328 9.3005
R738 VTAIL.n307 VTAIL.n306 9.3005
R739 VTAIL.n305 VTAIL.n304 9.3005
R740 VTAIL.n240 VTAIL.n239 9.3005
R741 VTAIL.n299 VTAIL.n298 9.3005
R742 VTAIL.n297 VTAIL.n296 9.3005
R743 VTAIL.n244 VTAIL.n243 9.3005
R744 VTAIL.n291 VTAIL.n290 9.3005
R745 VTAIL.n289 VTAIL.n288 9.3005
R746 VTAIL.n248 VTAIL.n247 9.3005
R747 VTAIL.n154 VTAIL.n153 9.3005
R748 VTAIL.n156 VTAIL.n155 9.3005
R749 VTAIL.n147 VTAIL.n146 9.3005
R750 VTAIL.n162 VTAIL.n161 9.3005
R751 VTAIL.n164 VTAIL.n163 9.3005
R752 VTAIL.n142 VTAIL.n141 9.3005
R753 VTAIL.n170 VTAIL.n169 9.3005
R754 VTAIL.n172 VTAIL.n171 9.3005
R755 VTAIL.n126 VTAIL.n125 9.3005
R756 VTAIL.n203 VTAIL.n202 9.3005
R757 VTAIL.n205 VTAIL.n204 9.3005
R758 VTAIL.n122 VTAIL.n121 9.3005
R759 VTAIL.n211 VTAIL.n210 9.3005
R760 VTAIL.n213 VTAIL.n212 9.3005
R761 VTAIL.n118 VTAIL.n117 9.3005
R762 VTAIL.n219 VTAIL.n218 9.3005
R763 VTAIL.n197 VTAIL.n196 9.3005
R764 VTAIL.n195 VTAIL.n194 9.3005
R765 VTAIL.n130 VTAIL.n129 9.3005
R766 VTAIL.n189 VTAIL.n188 9.3005
R767 VTAIL.n187 VTAIL.n186 9.3005
R768 VTAIL.n134 VTAIL.n133 9.3005
R769 VTAIL.n181 VTAIL.n180 9.3005
R770 VTAIL.n179 VTAIL.n178 9.3005
R771 VTAIL.n138 VTAIL.n137 9.3005
R772 VTAIL.n372 VTAIL.n362 8.92171
R773 VTAIL.n406 VTAIL.n405 8.92171
R774 VTAIL.n421 VTAIL.n340 8.92171
R775 VTAIL.n42 VTAIL.n32 8.92171
R776 VTAIL.n76 VTAIL.n75 8.92171
R777 VTAIL.n91 VTAIL.n10 8.92171
R778 VTAIL.n315 VTAIL.n234 8.92171
R779 VTAIL.n300 VTAIL.n299 8.92171
R780 VTAIL.n267 VTAIL.n257 8.92171
R781 VTAIL.n205 VTAIL.n124 8.92171
R782 VTAIL.n190 VTAIL.n189 8.92171
R783 VTAIL.n157 VTAIL.n147 8.92171
R784 VTAIL.n371 VTAIL.n364 8.14595
R785 VTAIL.n409 VTAIL.n346 8.14595
R786 VTAIL.n418 VTAIL.n417 8.14595
R787 VTAIL.n41 VTAIL.n34 8.14595
R788 VTAIL.n79 VTAIL.n16 8.14595
R789 VTAIL.n88 VTAIL.n87 8.14595
R790 VTAIL.n312 VTAIL.n311 8.14595
R791 VTAIL.n303 VTAIL.n240 8.14595
R792 VTAIL.n266 VTAIL.n259 8.14595
R793 VTAIL.n202 VTAIL.n201 8.14595
R794 VTAIL.n193 VTAIL.n130 8.14595
R795 VTAIL.n156 VTAIL.n149 8.14595
R796 VTAIL.n436 VTAIL.n332 7.75445
R797 VTAIL.n106 VTAIL.n2 7.75445
R798 VTAIL.n330 VTAIL.n226 7.75445
R799 VTAIL.n220 VTAIL.n116 7.75445
R800 VTAIL.n368 VTAIL.n367 7.3702
R801 VTAIL.n410 VTAIL.n344 7.3702
R802 VTAIL.n414 VTAIL.n342 7.3702
R803 VTAIL.n38 VTAIL.n37 7.3702
R804 VTAIL.n80 VTAIL.n14 7.3702
R805 VTAIL.n84 VTAIL.n12 7.3702
R806 VTAIL.n308 VTAIL.n236 7.3702
R807 VTAIL.n304 VTAIL.n238 7.3702
R808 VTAIL.n263 VTAIL.n262 7.3702
R809 VTAIL.n198 VTAIL.n126 7.3702
R810 VTAIL.n194 VTAIL.n128 7.3702
R811 VTAIL.n153 VTAIL.n152 7.3702
R812 VTAIL.n413 VTAIL.n344 6.59444
R813 VTAIL.n414 VTAIL.n413 6.59444
R814 VTAIL.n83 VTAIL.n14 6.59444
R815 VTAIL.n84 VTAIL.n83 6.59444
R816 VTAIL.n308 VTAIL.n307 6.59444
R817 VTAIL.n307 VTAIL.n238 6.59444
R818 VTAIL.n198 VTAIL.n197 6.59444
R819 VTAIL.n197 VTAIL.n128 6.59444
R820 VTAIL.n434 VTAIL.n332 6.08283
R821 VTAIL.n104 VTAIL.n2 6.08283
R822 VTAIL.n328 VTAIL.n226 6.08283
R823 VTAIL.n218 VTAIL.n116 6.08283
R824 VTAIL.n368 VTAIL.n364 5.81868
R825 VTAIL.n410 VTAIL.n409 5.81868
R826 VTAIL.n417 VTAIL.n342 5.81868
R827 VTAIL.n38 VTAIL.n34 5.81868
R828 VTAIL.n80 VTAIL.n79 5.81868
R829 VTAIL.n87 VTAIL.n12 5.81868
R830 VTAIL.n311 VTAIL.n236 5.81868
R831 VTAIL.n304 VTAIL.n303 5.81868
R832 VTAIL.n263 VTAIL.n259 5.81868
R833 VTAIL.n201 VTAIL.n126 5.81868
R834 VTAIL.n194 VTAIL.n193 5.81868
R835 VTAIL.n153 VTAIL.n149 5.81868
R836 VTAIL.n372 VTAIL.n371 5.04292
R837 VTAIL.n406 VTAIL.n346 5.04292
R838 VTAIL.n418 VTAIL.n340 5.04292
R839 VTAIL.n42 VTAIL.n41 5.04292
R840 VTAIL.n76 VTAIL.n16 5.04292
R841 VTAIL.n88 VTAIL.n10 5.04292
R842 VTAIL.n312 VTAIL.n234 5.04292
R843 VTAIL.n300 VTAIL.n240 5.04292
R844 VTAIL.n267 VTAIL.n266 5.04292
R845 VTAIL.n202 VTAIL.n124 5.04292
R846 VTAIL.n190 VTAIL.n130 5.04292
R847 VTAIL.n157 VTAIL.n156 5.04292
R848 VTAIL.n375 VTAIL.n362 4.26717
R849 VTAIL.n405 VTAIL.n348 4.26717
R850 VTAIL.n422 VTAIL.n421 4.26717
R851 VTAIL.n45 VTAIL.n32 4.26717
R852 VTAIL.n75 VTAIL.n18 4.26717
R853 VTAIL.n92 VTAIL.n91 4.26717
R854 VTAIL.n316 VTAIL.n315 4.26717
R855 VTAIL.n299 VTAIL.n242 4.26717
R856 VTAIL.n270 VTAIL.n257 4.26717
R857 VTAIL.n206 VTAIL.n205 4.26717
R858 VTAIL.n189 VTAIL.n132 4.26717
R859 VTAIL.n160 VTAIL.n147 4.26717
R860 VTAIL.n376 VTAIL.n360 3.49141
R861 VTAIL.n402 VTAIL.n401 3.49141
R862 VTAIL.n425 VTAIL.n338 3.49141
R863 VTAIL.n46 VTAIL.n30 3.49141
R864 VTAIL.n72 VTAIL.n71 3.49141
R865 VTAIL.n95 VTAIL.n8 3.49141
R866 VTAIL.n319 VTAIL.n232 3.49141
R867 VTAIL.n296 VTAIL.n295 3.49141
R868 VTAIL.n271 VTAIL.n255 3.49141
R869 VTAIL.n209 VTAIL.n122 3.49141
R870 VTAIL.n186 VTAIL.n185 3.49141
R871 VTAIL.n161 VTAIL.n145 3.49141
R872 VTAIL.n380 VTAIL.n379 2.71565
R873 VTAIL.n398 VTAIL.n350 2.71565
R874 VTAIL.n426 VTAIL.n336 2.71565
R875 VTAIL.n50 VTAIL.n49 2.71565
R876 VTAIL.n68 VTAIL.n20 2.71565
R877 VTAIL.n96 VTAIL.n6 2.71565
R878 VTAIL.n320 VTAIL.n230 2.71565
R879 VTAIL.n292 VTAIL.n244 2.71565
R880 VTAIL.n275 VTAIL.n274 2.71565
R881 VTAIL.n210 VTAIL.n120 2.71565
R882 VTAIL.n182 VTAIL.n134 2.71565
R883 VTAIL.n165 VTAIL.n164 2.71565
R884 VTAIL.n264 VTAIL.n260 2.41282
R885 VTAIL.n154 VTAIL.n150 2.41282
R886 VTAIL.n369 VTAIL.n365 2.41282
R887 VTAIL.n39 VTAIL.n35 2.41282
R888 VTAIL.n384 VTAIL.n358 1.93989
R889 VTAIL.n397 VTAIL.n352 1.93989
R890 VTAIL.n430 VTAIL.n429 1.93989
R891 VTAIL.n54 VTAIL.n28 1.93989
R892 VTAIL.n67 VTAIL.n22 1.93989
R893 VTAIL.n100 VTAIL.n99 1.93989
R894 VTAIL.n324 VTAIL.n323 1.93989
R895 VTAIL.n291 VTAIL.n246 1.93989
R896 VTAIL.n278 VTAIL.n252 1.93989
R897 VTAIL.n214 VTAIL.n213 1.93989
R898 VTAIL.n181 VTAIL.n136 1.93989
R899 VTAIL.n168 VTAIL.n142 1.93989
R900 VTAIL.n438 VTAIL.t15 1.66401
R901 VTAIL.n438 VTAIL.t16 1.66401
R902 VTAIL.n0 VTAIL.t11 1.66401
R903 VTAIL.n0 VTAIL.t13 1.66401
R904 VTAIL.n108 VTAIL.t19 1.66401
R905 VTAIL.n108 VTAIL.t17 1.66401
R906 VTAIL.n110 VTAIL.t2 1.66401
R907 VTAIL.n110 VTAIL.t1 1.66401
R908 VTAIL.n224 VTAIL.t18 1.66401
R909 VTAIL.n224 VTAIL.t5 1.66401
R910 VTAIL.n222 VTAIL.t3 1.66401
R911 VTAIL.n222 VTAIL.t4 1.66401
R912 VTAIL.n114 VTAIL.t8 1.66401
R913 VTAIL.n114 VTAIL.t14 1.66401
R914 VTAIL.n112 VTAIL.t12 1.66401
R915 VTAIL.n112 VTAIL.t9 1.66401
R916 VTAIL.n385 VTAIL.n356 1.16414
R917 VTAIL.n394 VTAIL.n393 1.16414
R918 VTAIL.n433 VTAIL.n334 1.16414
R919 VTAIL.n55 VTAIL.n26 1.16414
R920 VTAIL.n64 VTAIL.n63 1.16414
R921 VTAIL.n103 VTAIL.n4 1.16414
R922 VTAIL.n327 VTAIL.n228 1.16414
R923 VTAIL.n288 VTAIL.n287 1.16414
R924 VTAIL.n279 VTAIL.n250 1.16414
R925 VTAIL.n217 VTAIL.n118 1.16414
R926 VTAIL.n178 VTAIL.n177 1.16414
R927 VTAIL.n169 VTAIL.n140 1.16414
R928 VTAIL.n223 VTAIL.n221 0.685845
R929 VTAIL.n107 VTAIL.n1 0.685845
R930 VTAIL.n115 VTAIL.n113 0.431534
R931 VTAIL.n221 VTAIL.n115 0.431534
R932 VTAIL.n225 VTAIL.n223 0.431534
R933 VTAIL.n331 VTAIL.n225 0.431534
R934 VTAIL.n111 VTAIL.n109 0.431534
R935 VTAIL.n109 VTAIL.n107 0.431534
R936 VTAIL.n439 VTAIL.n437 0.431534
R937 VTAIL.n389 VTAIL.n388 0.388379
R938 VTAIL.n390 VTAIL.n354 0.388379
R939 VTAIL.n59 VTAIL.n58 0.388379
R940 VTAIL.n60 VTAIL.n24 0.388379
R941 VTAIL.n284 VTAIL.n248 0.388379
R942 VTAIL.n283 VTAIL.n282 0.388379
R943 VTAIL.n174 VTAIL.n138 0.388379
R944 VTAIL.n173 VTAIL.n172 0.388379
R945 VTAIL VTAIL.n1 0.381966
R946 VTAIL.n370 VTAIL.n369 0.155672
R947 VTAIL.n370 VTAIL.n361 0.155672
R948 VTAIL.n377 VTAIL.n361 0.155672
R949 VTAIL.n378 VTAIL.n377 0.155672
R950 VTAIL.n378 VTAIL.n357 0.155672
R951 VTAIL.n386 VTAIL.n357 0.155672
R952 VTAIL.n387 VTAIL.n386 0.155672
R953 VTAIL.n387 VTAIL.n353 0.155672
R954 VTAIL.n395 VTAIL.n353 0.155672
R955 VTAIL.n396 VTAIL.n395 0.155672
R956 VTAIL.n396 VTAIL.n349 0.155672
R957 VTAIL.n403 VTAIL.n349 0.155672
R958 VTAIL.n404 VTAIL.n403 0.155672
R959 VTAIL.n404 VTAIL.n345 0.155672
R960 VTAIL.n411 VTAIL.n345 0.155672
R961 VTAIL.n412 VTAIL.n411 0.155672
R962 VTAIL.n412 VTAIL.n341 0.155672
R963 VTAIL.n419 VTAIL.n341 0.155672
R964 VTAIL.n420 VTAIL.n419 0.155672
R965 VTAIL.n420 VTAIL.n337 0.155672
R966 VTAIL.n427 VTAIL.n337 0.155672
R967 VTAIL.n428 VTAIL.n427 0.155672
R968 VTAIL.n428 VTAIL.n333 0.155672
R969 VTAIL.n435 VTAIL.n333 0.155672
R970 VTAIL.n40 VTAIL.n39 0.155672
R971 VTAIL.n40 VTAIL.n31 0.155672
R972 VTAIL.n47 VTAIL.n31 0.155672
R973 VTAIL.n48 VTAIL.n47 0.155672
R974 VTAIL.n48 VTAIL.n27 0.155672
R975 VTAIL.n56 VTAIL.n27 0.155672
R976 VTAIL.n57 VTAIL.n56 0.155672
R977 VTAIL.n57 VTAIL.n23 0.155672
R978 VTAIL.n65 VTAIL.n23 0.155672
R979 VTAIL.n66 VTAIL.n65 0.155672
R980 VTAIL.n66 VTAIL.n19 0.155672
R981 VTAIL.n73 VTAIL.n19 0.155672
R982 VTAIL.n74 VTAIL.n73 0.155672
R983 VTAIL.n74 VTAIL.n15 0.155672
R984 VTAIL.n81 VTAIL.n15 0.155672
R985 VTAIL.n82 VTAIL.n81 0.155672
R986 VTAIL.n82 VTAIL.n11 0.155672
R987 VTAIL.n89 VTAIL.n11 0.155672
R988 VTAIL.n90 VTAIL.n89 0.155672
R989 VTAIL.n90 VTAIL.n7 0.155672
R990 VTAIL.n97 VTAIL.n7 0.155672
R991 VTAIL.n98 VTAIL.n97 0.155672
R992 VTAIL.n98 VTAIL.n3 0.155672
R993 VTAIL.n105 VTAIL.n3 0.155672
R994 VTAIL.n329 VTAIL.n227 0.155672
R995 VTAIL.n322 VTAIL.n227 0.155672
R996 VTAIL.n322 VTAIL.n321 0.155672
R997 VTAIL.n321 VTAIL.n231 0.155672
R998 VTAIL.n314 VTAIL.n231 0.155672
R999 VTAIL.n314 VTAIL.n313 0.155672
R1000 VTAIL.n313 VTAIL.n235 0.155672
R1001 VTAIL.n306 VTAIL.n235 0.155672
R1002 VTAIL.n306 VTAIL.n305 0.155672
R1003 VTAIL.n305 VTAIL.n239 0.155672
R1004 VTAIL.n298 VTAIL.n239 0.155672
R1005 VTAIL.n298 VTAIL.n297 0.155672
R1006 VTAIL.n297 VTAIL.n243 0.155672
R1007 VTAIL.n290 VTAIL.n243 0.155672
R1008 VTAIL.n290 VTAIL.n289 0.155672
R1009 VTAIL.n289 VTAIL.n247 0.155672
R1010 VTAIL.n281 VTAIL.n247 0.155672
R1011 VTAIL.n281 VTAIL.n280 0.155672
R1012 VTAIL.n280 VTAIL.n251 0.155672
R1013 VTAIL.n273 VTAIL.n251 0.155672
R1014 VTAIL.n273 VTAIL.n272 0.155672
R1015 VTAIL.n272 VTAIL.n256 0.155672
R1016 VTAIL.n265 VTAIL.n256 0.155672
R1017 VTAIL.n265 VTAIL.n264 0.155672
R1018 VTAIL.n219 VTAIL.n117 0.155672
R1019 VTAIL.n212 VTAIL.n117 0.155672
R1020 VTAIL.n212 VTAIL.n211 0.155672
R1021 VTAIL.n211 VTAIL.n121 0.155672
R1022 VTAIL.n204 VTAIL.n121 0.155672
R1023 VTAIL.n204 VTAIL.n203 0.155672
R1024 VTAIL.n203 VTAIL.n125 0.155672
R1025 VTAIL.n196 VTAIL.n125 0.155672
R1026 VTAIL.n196 VTAIL.n195 0.155672
R1027 VTAIL.n195 VTAIL.n129 0.155672
R1028 VTAIL.n188 VTAIL.n129 0.155672
R1029 VTAIL.n188 VTAIL.n187 0.155672
R1030 VTAIL.n187 VTAIL.n133 0.155672
R1031 VTAIL.n180 VTAIL.n133 0.155672
R1032 VTAIL.n180 VTAIL.n179 0.155672
R1033 VTAIL.n179 VTAIL.n137 0.155672
R1034 VTAIL.n171 VTAIL.n137 0.155672
R1035 VTAIL.n171 VTAIL.n170 0.155672
R1036 VTAIL.n170 VTAIL.n141 0.155672
R1037 VTAIL.n163 VTAIL.n141 0.155672
R1038 VTAIL.n163 VTAIL.n162 0.155672
R1039 VTAIL.n162 VTAIL.n146 0.155672
R1040 VTAIL.n155 VTAIL.n146 0.155672
R1041 VTAIL.n155 VTAIL.n154 0.155672
R1042 VTAIL VTAIL.n439 0.050069
R1043 VP.n19 VP.t8 2990.89
R1044 VP.n12 VP.t3 2990.89
R1045 VP.n4 VP.t1 2990.89
R1046 VP.n10 VP.t0 2990.89
R1047 VP.n18 VP.t7 2954.38
R1048 VP.n16 VP.t6 2954.38
R1049 VP.n1 VP.t4 2954.38
R1050 VP.n3 VP.t9 2954.38
R1051 VP.n7 VP.t5 2954.38
R1052 VP.n9 VP.t2 2954.38
R1053 VP.n5 VP.n4 161.489
R1054 VP.n20 VP.n19 161.3
R1055 VP.n6 VP.n5 161.3
R1056 VP.n8 VP.n2 161.3
R1057 VP.n11 VP.n10 161.3
R1058 VP.n17 VP.n0 161.3
R1059 VP.n15 VP.n14 161.3
R1060 VP.n13 VP.n12 161.3
R1061 VP.n13 VP.n11 45.6293
R1062 VP.n12 VP.n1 36.5157
R1063 VP.n15 VP.n1 36.5157
R1064 VP.n16 VP.n15 36.5157
R1065 VP.n17 VP.n16 36.5157
R1066 VP.n18 VP.n17 36.5157
R1067 VP.n19 VP.n18 36.5157
R1068 VP.n4 VP.n3 36.5157
R1069 VP.n6 VP.n3 36.5157
R1070 VP.n7 VP.n6 36.5157
R1071 VP.n8 VP.n7 36.5157
R1072 VP.n9 VP.n8 36.5157
R1073 VP.n10 VP.n9 36.5157
R1074 VP.n5 VP.n2 0.189894
R1075 VP.n11 VP.n2 0.189894
R1076 VP.n14 VP.n13 0.189894
R1077 VP.n14 VP.n0 0.189894
R1078 VP.n20 VP.n0 0.189894
R1079 VP VP.n20 0.0516364
R1080 VDD1.n101 VDD1.n100 585
R1081 VDD1.n99 VDD1.n98 585
R1082 VDD1.n4 VDD1.n3 585
R1083 VDD1.n93 VDD1.n92 585
R1084 VDD1.n91 VDD1.n90 585
R1085 VDD1.n8 VDD1.n7 585
R1086 VDD1.n85 VDD1.n84 585
R1087 VDD1.n83 VDD1.n82 585
R1088 VDD1.n12 VDD1.n11 585
R1089 VDD1.n77 VDD1.n76 585
R1090 VDD1.n75 VDD1.n74 585
R1091 VDD1.n16 VDD1.n15 585
R1092 VDD1.n69 VDD1.n68 585
R1093 VDD1.n67 VDD1.n66 585
R1094 VDD1.n20 VDD1.n19 585
R1095 VDD1.n61 VDD1.n60 585
R1096 VDD1.n59 VDD1.n58 585
R1097 VDD1.n57 VDD1.n23 585
R1098 VDD1.n27 VDD1.n24 585
R1099 VDD1.n52 VDD1.n51 585
R1100 VDD1.n50 VDD1.n49 585
R1101 VDD1.n29 VDD1.n28 585
R1102 VDD1.n44 VDD1.n43 585
R1103 VDD1.n42 VDD1.n41 585
R1104 VDD1.n33 VDD1.n32 585
R1105 VDD1.n36 VDD1.n35 585
R1106 VDD1.n142 VDD1.n141 585
R1107 VDD1.n139 VDD1.n138 585
R1108 VDD1.n148 VDD1.n147 585
R1109 VDD1.n150 VDD1.n149 585
R1110 VDD1.n135 VDD1.n134 585
R1111 VDD1.n156 VDD1.n155 585
R1112 VDD1.n159 VDD1.n158 585
R1113 VDD1.n157 VDD1.n131 585
R1114 VDD1.n164 VDD1.n130 585
R1115 VDD1.n166 VDD1.n165 585
R1116 VDD1.n168 VDD1.n167 585
R1117 VDD1.n127 VDD1.n126 585
R1118 VDD1.n174 VDD1.n173 585
R1119 VDD1.n176 VDD1.n175 585
R1120 VDD1.n123 VDD1.n122 585
R1121 VDD1.n182 VDD1.n181 585
R1122 VDD1.n184 VDD1.n183 585
R1123 VDD1.n119 VDD1.n118 585
R1124 VDD1.n190 VDD1.n189 585
R1125 VDD1.n192 VDD1.n191 585
R1126 VDD1.n115 VDD1.n114 585
R1127 VDD1.n198 VDD1.n197 585
R1128 VDD1.n200 VDD1.n199 585
R1129 VDD1.n111 VDD1.n110 585
R1130 VDD1.n206 VDD1.n205 585
R1131 VDD1.n208 VDD1.n207 585
R1132 VDD1.n100 VDD1.n0 498.474
R1133 VDD1.n207 VDD1.n107 498.474
R1134 VDD1.t8 VDD1.n34 329.036
R1135 VDD1.t6 VDD1.n140 329.036
R1136 VDD1.n100 VDD1.n99 171.744
R1137 VDD1.n99 VDD1.n3 171.744
R1138 VDD1.n92 VDD1.n3 171.744
R1139 VDD1.n92 VDD1.n91 171.744
R1140 VDD1.n91 VDD1.n7 171.744
R1141 VDD1.n84 VDD1.n7 171.744
R1142 VDD1.n84 VDD1.n83 171.744
R1143 VDD1.n83 VDD1.n11 171.744
R1144 VDD1.n76 VDD1.n11 171.744
R1145 VDD1.n76 VDD1.n75 171.744
R1146 VDD1.n75 VDD1.n15 171.744
R1147 VDD1.n68 VDD1.n15 171.744
R1148 VDD1.n68 VDD1.n67 171.744
R1149 VDD1.n67 VDD1.n19 171.744
R1150 VDD1.n60 VDD1.n19 171.744
R1151 VDD1.n60 VDD1.n59 171.744
R1152 VDD1.n59 VDD1.n23 171.744
R1153 VDD1.n27 VDD1.n23 171.744
R1154 VDD1.n51 VDD1.n27 171.744
R1155 VDD1.n51 VDD1.n50 171.744
R1156 VDD1.n50 VDD1.n28 171.744
R1157 VDD1.n43 VDD1.n28 171.744
R1158 VDD1.n43 VDD1.n42 171.744
R1159 VDD1.n42 VDD1.n32 171.744
R1160 VDD1.n35 VDD1.n32 171.744
R1161 VDD1.n141 VDD1.n138 171.744
R1162 VDD1.n148 VDD1.n138 171.744
R1163 VDD1.n149 VDD1.n148 171.744
R1164 VDD1.n149 VDD1.n134 171.744
R1165 VDD1.n156 VDD1.n134 171.744
R1166 VDD1.n158 VDD1.n156 171.744
R1167 VDD1.n158 VDD1.n157 171.744
R1168 VDD1.n157 VDD1.n130 171.744
R1169 VDD1.n166 VDD1.n130 171.744
R1170 VDD1.n167 VDD1.n166 171.744
R1171 VDD1.n167 VDD1.n126 171.744
R1172 VDD1.n174 VDD1.n126 171.744
R1173 VDD1.n175 VDD1.n174 171.744
R1174 VDD1.n175 VDD1.n122 171.744
R1175 VDD1.n182 VDD1.n122 171.744
R1176 VDD1.n183 VDD1.n182 171.744
R1177 VDD1.n183 VDD1.n118 171.744
R1178 VDD1.n190 VDD1.n118 171.744
R1179 VDD1.n191 VDD1.n190 171.744
R1180 VDD1.n191 VDD1.n114 171.744
R1181 VDD1.n198 VDD1.n114 171.744
R1182 VDD1.n199 VDD1.n198 171.744
R1183 VDD1.n199 VDD1.n110 171.744
R1184 VDD1.n206 VDD1.n110 171.744
R1185 VDD1.n207 VDD1.n206 171.744
R1186 VDD1.n35 VDD1.t8 85.8723
R1187 VDD1.n141 VDD1.t6 85.8723
R1188 VDD1.n215 VDD1.n214 72.3777
R1189 VDD1.n106 VDD1.n105 72.1099
R1190 VDD1.n217 VDD1.n216 72.1098
R1191 VDD1.n213 VDD1.n212 72.1098
R1192 VDD1.n106 VDD1.n104 53.5618
R1193 VDD1.n213 VDD1.n211 53.5618
R1194 VDD1.n217 VDD1.n215 43.4061
R1195 VDD1.n58 VDD1.n57 13.1884
R1196 VDD1.n165 VDD1.n164 13.1884
R1197 VDD1.n102 VDD1.n101 12.8005
R1198 VDD1.n61 VDD1.n22 12.8005
R1199 VDD1.n56 VDD1.n24 12.8005
R1200 VDD1.n163 VDD1.n131 12.8005
R1201 VDD1.n168 VDD1.n129 12.8005
R1202 VDD1.n209 VDD1.n208 12.8005
R1203 VDD1.n98 VDD1.n2 12.0247
R1204 VDD1.n62 VDD1.n20 12.0247
R1205 VDD1.n53 VDD1.n52 12.0247
R1206 VDD1.n160 VDD1.n159 12.0247
R1207 VDD1.n169 VDD1.n127 12.0247
R1208 VDD1.n205 VDD1.n109 12.0247
R1209 VDD1.n97 VDD1.n4 11.249
R1210 VDD1.n66 VDD1.n65 11.249
R1211 VDD1.n49 VDD1.n26 11.249
R1212 VDD1.n155 VDD1.n133 11.249
R1213 VDD1.n173 VDD1.n172 11.249
R1214 VDD1.n204 VDD1.n111 11.249
R1215 VDD1.n36 VDD1.n34 10.7239
R1216 VDD1.n142 VDD1.n140 10.7239
R1217 VDD1.n94 VDD1.n93 10.4732
R1218 VDD1.n69 VDD1.n18 10.4732
R1219 VDD1.n48 VDD1.n29 10.4732
R1220 VDD1.n154 VDD1.n135 10.4732
R1221 VDD1.n176 VDD1.n125 10.4732
R1222 VDD1.n201 VDD1.n200 10.4732
R1223 VDD1.n90 VDD1.n6 9.69747
R1224 VDD1.n70 VDD1.n16 9.69747
R1225 VDD1.n45 VDD1.n44 9.69747
R1226 VDD1.n151 VDD1.n150 9.69747
R1227 VDD1.n177 VDD1.n123 9.69747
R1228 VDD1.n197 VDD1.n113 9.69747
R1229 VDD1.n104 VDD1.n103 9.45567
R1230 VDD1.n211 VDD1.n210 9.45567
R1231 VDD1.n38 VDD1.n37 9.3005
R1232 VDD1.n40 VDD1.n39 9.3005
R1233 VDD1.n31 VDD1.n30 9.3005
R1234 VDD1.n46 VDD1.n45 9.3005
R1235 VDD1.n48 VDD1.n47 9.3005
R1236 VDD1.n26 VDD1.n25 9.3005
R1237 VDD1.n54 VDD1.n53 9.3005
R1238 VDD1.n56 VDD1.n55 9.3005
R1239 VDD1.n10 VDD1.n9 9.3005
R1240 VDD1.n87 VDD1.n86 9.3005
R1241 VDD1.n89 VDD1.n88 9.3005
R1242 VDD1.n6 VDD1.n5 9.3005
R1243 VDD1.n95 VDD1.n94 9.3005
R1244 VDD1.n97 VDD1.n96 9.3005
R1245 VDD1.n2 VDD1.n1 9.3005
R1246 VDD1.n103 VDD1.n102 9.3005
R1247 VDD1.n81 VDD1.n80 9.3005
R1248 VDD1.n79 VDD1.n78 9.3005
R1249 VDD1.n14 VDD1.n13 9.3005
R1250 VDD1.n73 VDD1.n72 9.3005
R1251 VDD1.n71 VDD1.n70 9.3005
R1252 VDD1.n18 VDD1.n17 9.3005
R1253 VDD1.n65 VDD1.n64 9.3005
R1254 VDD1.n63 VDD1.n62 9.3005
R1255 VDD1.n22 VDD1.n21 9.3005
R1256 VDD1.n186 VDD1.n185 9.3005
R1257 VDD1.n121 VDD1.n120 9.3005
R1258 VDD1.n180 VDD1.n179 9.3005
R1259 VDD1.n178 VDD1.n177 9.3005
R1260 VDD1.n125 VDD1.n124 9.3005
R1261 VDD1.n172 VDD1.n171 9.3005
R1262 VDD1.n170 VDD1.n169 9.3005
R1263 VDD1.n129 VDD1.n128 9.3005
R1264 VDD1.n144 VDD1.n143 9.3005
R1265 VDD1.n146 VDD1.n145 9.3005
R1266 VDD1.n137 VDD1.n136 9.3005
R1267 VDD1.n152 VDD1.n151 9.3005
R1268 VDD1.n154 VDD1.n153 9.3005
R1269 VDD1.n133 VDD1.n132 9.3005
R1270 VDD1.n161 VDD1.n160 9.3005
R1271 VDD1.n163 VDD1.n162 9.3005
R1272 VDD1.n188 VDD1.n187 9.3005
R1273 VDD1.n117 VDD1.n116 9.3005
R1274 VDD1.n194 VDD1.n193 9.3005
R1275 VDD1.n196 VDD1.n195 9.3005
R1276 VDD1.n113 VDD1.n112 9.3005
R1277 VDD1.n202 VDD1.n201 9.3005
R1278 VDD1.n204 VDD1.n203 9.3005
R1279 VDD1.n109 VDD1.n108 9.3005
R1280 VDD1.n210 VDD1.n209 9.3005
R1281 VDD1.n89 VDD1.n8 8.92171
R1282 VDD1.n74 VDD1.n73 8.92171
R1283 VDD1.n41 VDD1.n31 8.92171
R1284 VDD1.n147 VDD1.n137 8.92171
R1285 VDD1.n181 VDD1.n180 8.92171
R1286 VDD1.n196 VDD1.n115 8.92171
R1287 VDD1.n86 VDD1.n85 8.14595
R1288 VDD1.n77 VDD1.n14 8.14595
R1289 VDD1.n40 VDD1.n33 8.14595
R1290 VDD1.n146 VDD1.n139 8.14595
R1291 VDD1.n184 VDD1.n121 8.14595
R1292 VDD1.n193 VDD1.n192 8.14595
R1293 VDD1.n104 VDD1.n0 7.75445
R1294 VDD1.n211 VDD1.n107 7.75445
R1295 VDD1.n82 VDD1.n10 7.3702
R1296 VDD1.n78 VDD1.n12 7.3702
R1297 VDD1.n37 VDD1.n36 7.3702
R1298 VDD1.n143 VDD1.n142 7.3702
R1299 VDD1.n185 VDD1.n119 7.3702
R1300 VDD1.n189 VDD1.n117 7.3702
R1301 VDD1.n82 VDD1.n81 6.59444
R1302 VDD1.n81 VDD1.n12 6.59444
R1303 VDD1.n188 VDD1.n119 6.59444
R1304 VDD1.n189 VDD1.n188 6.59444
R1305 VDD1.n102 VDD1.n0 6.08283
R1306 VDD1.n209 VDD1.n107 6.08283
R1307 VDD1.n85 VDD1.n10 5.81868
R1308 VDD1.n78 VDD1.n77 5.81868
R1309 VDD1.n37 VDD1.n33 5.81868
R1310 VDD1.n143 VDD1.n139 5.81868
R1311 VDD1.n185 VDD1.n184 5.81868
R1312 VDD1.n192 VDD1.n117 5.81868
R1313 VDD1.n86 VDD1.n8 5.04292
R1314 VDD1.n74 VDD1.n14 5.04292
R1315 VDD1.n41 VDD1.n40 5.04292
R1316 VDD1.n147 VDD1.n146 5.04292
R1317 VDD1.n181 VDD1.n121 5.04292
R1318 VDD1.n193 VDD1.n115 5.04292
R1319 VDD1.n90 VDD1.n89 4.26717
R1320 VDD1.n73 VDD1.n16 4.26717
R1321 VDD1.n44 VDD1.n31 4.26717
R1322 VDD1.n150 VDD1.n137 4.26717
R1323 VDD1.n180 VDD1.n123 4.26717
R1324 VDD1.n197 VDD1.n196 4.26717
R1325 VDD1.n93 VDD1.n6 3.49141
R1326 VDD1.n70 VDD1.n69 3.49141
R1327 VDD1.n45 VDD1.n29 3.49141
R1328 VDD1.n151 VDD1.n135 3.49141
R1329 VDD1.n177 VDD1.n176 3.49141
R1330 VDD1.n200 VDD1.n113 3.49141
R1331 VDD1.n94 VDD1.n4 2.71565
R1332 VDD1.n66 VDD1.n18 2.71565
R1333 VDD1.n49 VDD1.n48 2.71565
R1334 VDD1.n155 VDD1.n154 2.71565
R1335 VDD1.n173 VDD1.n125 2.71565
R1336 VDD1.n201 VDD1.n111 2.71565
R1337 VDD1.n38 VDD1.n34 2.41282
R1338 VDD1.n144 VDD1.n140 2.41282
R1339 VDD1.n98 VDD1.n97 1.93989
R1340 VDD1.n65 VDD1.n20 1.93989
R1341 VDD1.n52 VDD1.n26 1.93989
R1342 VDD1.n159 VDD1.n133 1.93989
R1343 VDD1.n172 VDD1.n127 1.93989
R1344 VDD1.n205 VDD1.n204 1.93989
R1345 VDD1.n216 VDD1.t7 1.66401
R1346 VDD1.n216 VDD1.t9 1.66401
R1347 VDD1.n105 VDD1.t0 1.66401
R1348 VDD1.n105 VDD1.t4 1.66401
R1349 VDD1.n214 VDD1.t2 1.66401
R1350 VDD1.n214 VDD1.t1 1.66401
R1351 VDD1.n212 VDD1.t5 1.66401
R1352 VDD1.n212 VDD1.t3 1.66401
R1353 VDD1.n101 VDD1.n2 1.16414
R1354 VDD1.n62 VDD1.n61 1.16414
R1355 VDD1.n53 VDD1.n24 1.16414
R1356 VDD1.n160 VDD1.n131 1.16414
R1357 VDD1.n169 VDD1.n168 1.16414
R1358 VDD1.n208 VDD1.n109 1.16414
R1359 VDD1.n58 VDD1.n22 0.388379
R1360 VDD1.n57 VDD1.n56 0.388379
R1361 VDD1.n164 VDD1.n163 0.388379
R1362 VDD1.n165 VDD1.n129 0.388379
R1363 VDD1 VDD1.n217 0.265586
R1364 VDD1 VDD1.n106 0.166448
R1365 VDD1.n103 VDD1.n1 0.155672
R1366 VDD1.n96 VDD1.n1 0.155672
R1367 VDD1.n96 VDD1.n95 0.155672
R1368 VDD1.n95 VDD1.n5 0.155672
R1369 VDD1.n88 VDD1.n5 0.155672
R1370 VDD1.n88 VDD1.n87 0.155672
R1371 VDD1.n87 VDD1.n9 0.155672
R1372 VDD1.n80 VDD1.n9 0.155672
R1373 VDD1.n80 VDD1.n79 0.155672
R1374 VDD1.n79 VDD1.n13 0.155672
R1375 VDD1.n72 VDD1.n13 0.155672
R1376 VDD1.n72 VDD1.n71 0.155672
R1377 VDD1.n71 VDD1.n17 0.155672
R1378 VDD1.n64 VDD1.n17 0.155672
R1379 VDD1.n64 VDD1.n63 0.155672
R1380 VDD1.n63 VDD1.n21 0.155672
R1381 VDD1.n55 VDD1.n21 0.155672
R1382 VDD1.n55 VDD1.n54 0.155672
R1383 VDD1.n54 VDD1.n25 0.155672
R1384 VDD1.n47 VDD1.n25 0.155672
R1385 VDD1.n47 VDD1.n46 0.155672
R1386 VDD1.n46 VDD1.n30 0.155672
R1387 VDD1.n39 VDD1.n30 0.155672
R1388 VDD1.n39 VDD1.n38 0.155672
R1389 VDD1.n145 VDD1.n144 0.155672
R1390 VDD1.n145 VDD1.n136 0.155672
R1391 VDD1.n152 VDD1.n136 0.155672
R1392 VDD1.n153 VDD1.n152 0.155672
R1393 VDD1.n153 VDD1.n132 0.155672
R1394 VDD1.n161 VDD1.n132 0.155672
R1395 VDD1.n162 VDD1.n161 0.155672
R1396 VDD1.n162 VDD1.n128 0.155672
R1397 VDD1.n170 VDD1.n128 0.155672
R1398 VDD1.n171 VDD1.n170 0.155672
R1399 VDD1.n171 VDD1.n124 0.155672
R1400 VDD1.n178 VDD1.n124 0.155672
R1401 VDD1.n179 VDD1.n178 0.155672
R1402 VDD1.n179 VDD1.n120 0.155672
R1403 VDD1.n186 VDD1.n120 0.155672
R1404 VDD1.n187 VDD1.n186 0.155672
R1405 VDD1.n187 VDD1.n116 0.155672
R1406 VDD1.n194 VDD1.n116 0.155672
R1407 VDD1.n195 VDD1.n194 0.155672
R1408 VDD1.n195 VDD1.n112 0.155672
R1409 VDD1.n202 VDD1.n112 0.155672
R1410 VDD1.n203 VDD1.n202 0.155672
R1411 VDD1.n203 VDD1.n108 0.155672
R1412 VDD1.n210 VDD1.n108 0.155672
R1413 VDD1.n215 VDD1.n213 0.0529126
R1414 B.n313 B.t6 3017.06
R1415 B.n139 B.t3 3017.06
R1416 B.n44 B.t9 3017.06
R1417 B.n51 B.t0 3017.06
R1418 B.n467 B.n466 585
R1419 B.n468 B.n83 585
R1420 B.n470 B.n469 585
R1421 B.n471 B.n82 585
R1422 B.n473 B.n472 585
R1423 B.n474 B.n81 585
R1424 B.n476 B.n475 585
R1425 B.n477 B.n80 585
R1426 B.n479 B.n478 585
R1427 B.n480 B.n79 585
R1428 B.n482 B.n481 585
R1429 B.n483 B.n78 585
R1430 B.n485 B.n484 585
R1431 B.n486 B.n77 585
R1432 B.n488 B.n487 585
R1433 B.n489 B.n76 585
R1434 B.n491 B.n490 585
R1435 B.n492 B.n75 585
R1436 B.n494 B.n493 585
R1437 B.n495 B.n74 585
R1438 B.n497 B.n496 585
R1439 B.n498 B.n73 585
R1440 B.n500 B.n499 585
R1441 B.n501 B.n72 585
R1442 B.n503 B.n502 585
R1443 B.n504 B.n71 585
R1444 B.n506 B.n505 585
R1445 B.n507 B.n70 585
R1446 B.n509 B.n508 585
R1447 B.n510 B.n69 585
R1448 B.n512 B.n511 585
R1449 B.n513 B.n68 585
R1450 B.n515 B.n514 585
R1451 B.n516 B.n67 585
R1452 B.n518 B.n517 585
R1453 B.n519 B.n66 585
R1454 B.n521 B.n520 585
R1455 B.n522 B.n65 585
R1456 B.n524 B.n523 585
R1457 B.n525 B.n64 585
R1458 B.n527 B.n526 585
R1459 B.n528 B.n63 585
R1460 B.n530 B.n529 585
R1461 B.n531 B.n62 585
R1462 B.n533 B.n532 585
R1463 B.n534 B.n61 585
R1464 B.n536 B.n535 585
R1465 B.n537 B.n60 585
R1466 B.n539 B.n538 585
R1467 B.n540 B.n59 585
R1468 B.n542 B.n541 585
R1469 B.n543 B.n58 585
R1470 B.n545 B.n544 585
R1471 B.n546 B.n57 585
R1472 B.n548 B.n547 585
R1473 B.n549 B.n56 585
R1474 B.n551 B.n550 585
R1475 B.n552 B.n55 585
R1476 B.n554 B.n553 585
R1477 B.n555 B.n54 585
R1478 B.n557 B.n556 585
R1479 B.n558 B.n53 585
R1480 B.n560 B.n559 585
R1481 B.n561 B.n50 585
R1482 B.n564 B.n563 585
R1483 B.n565 B.n49 585
R1484 B.n567 B.n566 585
R1485 B.n568 B.n48 585
R1486 B.n570 B.n569 585
R1487 B.n571 B.n47 585
R1488 B.n573 B.n572 585
R1489 B.n574 B.n43 585
R1490 B.n576 B.n575 585
R1491 B.n577 B.n42 585
R1492 B.n579 B.n578 585
R1493 B.n580 B.n41 585
R1494 B.n582 B.n581 585
R1495 B.n583 B.n40 585
R1496 B.n585 B.n584 585
R1497 B.n586 B.n39 585
R1498 B.n588 B.n587 585
R1499 B.n589 B.n38 585
R1500 B.n591 B.n590 585
R1501 B.n592 B.n37 585
R1502 B.n594 B.n593 585
R1503 B.n595 B.n36 585
R1504 B.n597 B.n596 585
R1505 B.n598 B.n35 585
R1506 B.n600 B.n599 585
R1507 B.n601 B.n34 585
R1508 B.n603 B.n602 585
R1509 B.n604 B.n33 585
R1510 B.n606 B.n605 585
R1511 B.n607 B.n32 585
R1512 B.n609 B.n608 585
R1513 B.n610 B.n31 585
R1514 B.n612 B.n611 585
R1515 B.n613 B.n30 585
R1516 B.n615 B.n614 585
R1517 B.n616 B.n29 585
R1518 B.n618 B.n617 585
R1519 B.n619 B.n28 585
R1520 B.n621 B.n620 585
R1521 B.n622 B.n27 585
R1522 B.n624 B.n623 585
R1523 B.n625 B.n26 585
R1524 B.n627 B.n626 585
R1525 B.n628 B.n25 585
R1526 B.n630 B.n629 585
R1527 B.n631 B.n24 585
R1528 B.n633 B.n632 585
R1529 B.n634 B.n23 585
R1530 B.n636 B.n635 585
R1531 B.n637 B.n22 585
R1532 B.n639 B.n638 585
R1533 B.n640 B.n21 585
R1534 B.n642 B.n641 585
R1535 B.n643 B.n20 585
R1536 B.n645 B.n644 585
R1537 B.n646 B.n19 585
R1538 B.n648 B.n647 585
R1539 B.n649 B.n18 585
R1540 B.n651 B.n650 585
R1541 B.n652 B.n17 585
R1542 B.n654 B.n653 585
R1543 B.n655 B.n16 585
R1544 B.n657 B.n656 585
R1545 B.n658 B.n15 585
R1546 B.n660 B.n659 585
R1547 B.n661 B.n14 585
R1548 B.n663 B.n662 585
R1549 B.n664 B.n13 585
R1550 B.n666 B.n665 585
R1551 B.n667 B.n12 585
R1552 B.n669 B.n668 585
R1553 B.n670 B.n11 585
R1554 B.n672 B.n671 585
R1555 B.n465 B.n84 585
R1556 B.n464 B.n463 585
R1557 B.n462 B.n85 585
R1558 B.n461 B.n460 585
R1559 B.n459 B.n86 585
R1560 B.n458 B.n457 585
R1561 B.n456 B.n87 585
R1562 B.n455 B.n454 585
R1563 B.n453 B.n88 585
R1564 B.n452 B.n451 585
R1565 B.n450 B.n89 585
R1566 B.n449 B.n448 585
R1567 B.n447 B.n90 585
R1568 B.n446 B.n445 585
R1569 B.n444 B.n91 585
R1570 B.n443 B.n442 585
R1571 B.n441 B.n92 585
R1572 B.n440 B.n439 585
R1573 B.n438 B.n93 585
R1574 B.n437 B.n436 585
R1575 B.n435 B.n94 585
R1576 B.n434 B.n433 585
R1577 B.n432 B.n95 585
R1578 B.n431 B.n430 585
R1579 B.n429 B.n96 585
R1580 B.n428 B.n427 585
R1581 B.n426 B.n97 585
R1582 B.n425 B.n424 585
R1583 B.n423 B.n98 585
R1584 B.n422 B.n421 585
R1585 B.n420 B.n99 585
R1586 B.n419 B.n418 585
R1587 B.n417 B.n100 585
R1588 B.n416 B.n415 585
R1589 B.n414 B.n101 585
R1590 B.n205 B.n204 585
R1591 B.n206 B.n171 585
R1592 B.n208 B.n207 585
R1593 B.n209 B.n170 585
R1594 B.n211 B.n210 585
R1595 B.n212 B.n169 585
R1596 B.n214 B.n213 585
R1597 B.n215 B.n168 585
R1598 B.n217 B.n216 585
R1599 B.n218 B.n167 585
R1600 B.n220 B.n219 585
R1601 B.n221 B.n166 585
R1602 B.n223 B.n222 585
R1603 B.n224 B.n165 585
R1604 B.n226 B.n225 585
R1605 B.n227 B.n164 585
R1606 B.n229 B.n228 585
R1607 B.n230 B.n163 585
R1608 B.n232 B.n231 585
R1609 B.n233 B.n162 585
R1610 B.n235 B.n234 585
R1611 B.n236 B.n161 585
R1612 B.n238 B.n237 585
R1613 B.n239 B.n160 585
R1614 B.n241 B.n240 585
R1615 B.n242 B.n159 585
R1616 B.n244 B.n243 585
R1617 B.n245 B.n158 585
R1618 B.n247 B.n246 585
R1619 B.n248 B.n157 585
R1620 B.n250 B.n249 585
R1621 B.n251 B.n156 585
R1622 B.n253 B.n252 585
R1623 B.n254 B.n155 585
R1624 B.n256 B.n255 585
R1625 B.n257 B.n154 585
R1626 B.n259 B.n258 585
R1627 B.n260 B.n153 585
R1628 B.n262 B.n261 585
R1629 B.n263 B.n152 585
R1630 B.n265 B.n264 585
R1631 B.n266 B.n151 585
R1632 B.n268 B.n267 585
R1633 B.n269 B.n150 585
R1634 B.n271 B.n270 585
R1635 B.n272 B.n149 585
R1636 B.n274 B.n273 585
R1637 B.n275 B.n148 585
R1638 B.n277 B.n276 585
R1639 B.n278 B.n147 585
R1640 B.n280 B.n279 585
R1641 B.n281 B.n146 585
R1642 B.n283 B.n282 585
R1643 B.n284 B.n145 585
R1644 B.n286 B.n285 585
R1645 B.n287 B.n144 585
R1646 B.n289 B.n288 585
R1647 B.n290 B.n143 585
R1648 B.n292 B.n291 585
R1649 B.n293 B.n142 585
R1650 B.n295 B.n294 585
R1651 B.n296 B.n141 585
R1652 B.n298 B.n297 585
R1653 B.n299 B.n138 585
R1654 B.n302 B.n301 585
R1655 B.n303 B.n137 585
R1656 B.n305 B.n304 585
R1657 B.n306 B.n136 585
R1658 B.n308 B.n307 585
R1659 B.n309 B.n135 585
R1660 B.n311 B.n310 585
R1661 B.n312 B.n134 585
R1662 B.n317 B.n316 585
R1663 B.n318 B.n133 585
R1664 B.n320 B.n319 585
R1665 B.n321 B.n132 585
R1666 B.n323 B.n322 585
R1667 B.n324 B.n131 585
R1668 B.n326 B.n325 585
R1669 B.n327 B.n130 585
R1670 B.n329 B.n328 585
R1671 B.n330 B.n129 585
R1672 B.n332 B.n331 585
R1673 B.n333 B.n128 585
R1674 B.n335 B.n334 585
R1675 B.n336 B.n127 585
R1676 B.n338 B.n337 585
R1677 B.n339 B.n126 585
R1678 B.n341 B.n340 585
R1679 B.n342 B.n125 585
R1680 B.n344 B.n343 585
R1681 B.n345 B.n124 585
R1682 B.n347 B.n346 585
R1683 B.n348 B.n123 585
R1684 B.n350 B.n349 585
R1685 B.n351 B.n122 585
R1686 B.n353 B.n352 585
R1687 B.n354 B.n121 585
R1688 B.n356 B.n355 585
R1689 B.n357 B.n120 585
R1690 B.n359 B.n358 585
R1691 B.n360 B.n119 585
R1692 B.n362 B.n361 585
R1693 B.n363 B.n118 585
R1694 B.n365 B.n364 585
R1695 B.n366 B.n117 585
R1696 B.n368 B.n367 585
R1697 B.n369 B.n116 585
R1698 B.n371 B.n370 585
R1699 B.n372 B.n115 585
R1700 B.n374 B.n373 585
R1701 B.n375 B.n114 585
R1702 B.n377 B.n376 585
R1703 B.n378 B.n113 585
R1704 B.n380 B.n379 585
R1705 B.n381 B.n112 585
R1706 B.n383 B.n382 585
R1707 B.n384 B.n111 585
R1708 B.n386 B.n385 585
R1709 B.n387 B.n110 585
R1710 B.n389 B.n388 585
R1711 B.n390 B.n109 585
R1712 B.n392 B.n391 585
R1713 B.n393 B.n108 585
R1714 B.n395 B.n394 585
R1715 B.n396 B.n107 585
R1716 B.n398 B.n397 585
R1717 B.n399 B.n106 585
R1718 B.n401 B.n400 585
R1719 B.n402 B.n105 585
R1720 B.n404 B.n403 585
R1721 B.n405 B.n104 585
R1722 B.n407 B.n406 585
R1723 B.n408 B.n103 585
R1724 B.n410 B.n409 585
R1725 B.n411 B.n102 585
R1726 B.n413 B.n412 585
R1727 B.n203 B.n172 585
R1728 B.n202 B.n201 585
R1729 B.n200 B.n173 585
R1730 B.n199 B.n198 585
R1731 B.n197 B.n174 585
R1732 B.n196 B.n195 585
R1733 B.n194 B.n175 585
R1734 B.n193 B.n192 585
R1735 B.n191 B.n176 585
R1736 B.n190 B.n189 585
R1737 B.n188 B.n177 585
R1738 B.n187 B.n186 585
R1739 B.n185 B.n178 585
R1740 B.n184 B.n183 585
R1741 B.n182 B.n179 585
R1742 B.n181 B.n180 585
R1743 B.n2 B.n0 585
R1744 B.n697 B.n1 585
R1745 B.n696 B.n695 585
R1746 B.n694 B.n3 585
R1747 B.n693 B.n692 585
R1748 B.n691 B.n4 585
R1749 B.n690 B.n689 585
R1750 B.n688 B.n5 585
R1751 B.n687 B.n686 585
R1752 B.n685 B.n6 585
R1753 B.n684 B.n683 585
R1754 B.n682 B.n7 585
R1755 B.n681 B.n680 585
R1756 B.n679 B.n8 585
R1757 B.n678 B.n677 585
R1758 B.n676 B.n9 585
R1759 B.n675 B.n674 585
R1760 B.n673 B.n10 585
R1761 B.n699 B.n698 585
R1762 B.n313 B.t8 521.119
R1763 B.n51 B.t1 521.119
R1764 B.n139 B.t5 521.119
R1765 B.n44 B.t10 521.119
R1766 B.n314 B.t7 511.421
R1767 B.n52 B.t2 511.421
R1768 B.n140 B.t4 511.421
R1769 B.n45 B.t11 511.421
R1770 B.n205 B.n172 502.111
R1771 B.n673 B.n672 502.111
R1772 B.n414 B.n413 502.111
R1773 B.n467 B.n84 502.111
R1774 B.n201 B.n172 163.367
R1775 B.n201 B.n200 163.367
R1776 B.n200 B.n199 163.367
R1777 B.n199 B.n174 163.367
R1778 B.n195 B.n174 163.367
R1779 B.n195 B.n194 163.367
R1780 B.n194 B.n193 163.367
R1781 B.n193 B.n176 163.367
R1782 B.n189 B.n176 163.367
R1783 B.n189 B.n188 163.367
R1784 B.n188 B.n187 163.367
R1785 B.n187 B.n178 163.367
R1786 B.n183 B.n178 163.367
R1787 B.n183 B.n182 163.367
R1788 B.n182 B.n181 163.367
R1789 B.n181 B.n2 163.367
R1790 B.n698 B.n2 163.367
R1791 B.n698 B.n697 163.367
R1792 B.n697 B.n696 163.367
R1793 B.n696 B.n3 163.367
R1794 B.n692 B.n3 163.367
R1795 B.n692 B.n691 163.367
R1796 B.n691 B.n690 163.367
R1797 B.n690 B.n5 163.367
R1798 B.n686 B.n5 163.367
R1799 B.n686 B.n685 163.367
R1800 B.n685 B.n684 163.367
R1801 B.n684 B.n7 163.367
R1802 B.n680 B.n7 163.367
R1803 B.n680 B.n679 163.367
R1804 B.n679 B.n678 163.367
R1805 B.n678 B.n9 163.367
R1806 B.n674 B.n9 163.367
R1807 B.n674 B.n673 163.367
R1808 B.n206 B.n205 163.367
R1809 B.n207 B.n206 163.367
R1810 B.n207 B.n170 163.367
R1811 B.n211 B.n170 163.367
R1812 B.n212 B.n211 163.367
R1813 B.n213 B.n212 163.367
R1814 B.n213 B.n168 163.367
R1815 B.n217 B.n168 163.367
R1816 B.n218 B.n217 163.367
R1817 B.n219 B.n218 163.367
R1818 B.n219 B.n166 163.367
R1819 B.n223 B.n166 163.367
R1820 B.n224 B.n223 163.367
R1821 B.n225 B.n224 163.367
R1822 B.n225 B.n164 163.367
R1823 B.n229 B.n164 163.367
R1824 B.n230 B.n229 163.367
R1825 B.n231 B.n230 163.367
R1826 B.n231 B.n162 163.367
R1827 B.n235 B.n162 163.367
R1828 B.n236 B.n235 163.367
R1829 B.n237 B.n236 163.367
R1830 B.n237 B.n160 163.367
R1831 B.n241 B.n160 163.367
R1832 B.n242 B.n241 163.367
R1833 B.n243 B.n242 163.367
R1834 B.n243 B.n158 163.367
R1835 B.n247 B.n158 163.367
R1836 B.n248 B.n247 163.367
R1837 B.n249 B.n248 163.367
R1838 B.n249 B.n156 163.367
R1839 B.n253 B.n156 163.367
R1840 B.n254 B.n253 163.367
R1841 B.n255 B.n254 163.367
R1842 B.n255 B.n154 163.367
R1843 B.n259 B.n154 163.367
R1844 B.n260 B.n259 163.367
R1845 B.n261 B.n260 163.367
R1846 B.n261 B.n152 163.367
R1847 B.n265 B.n152 163.367
R1848 B.n266 B.n265 163.367
R1849 B.n267 B.n266 163.367
R1850 B.n267 B.n150 163.367
R1851 B.n271 B.n150 163.367
R1852 B.n272 B.n271 163.367
R1853 B.n273 B.n272 163.367
R1854 B.n273 B.n148 163.367
R1855 B.n277 B.n148 163.367
R1856 B.n278 B.n277 163.367
R1857 B.n279 B.n278 163.367
R1858 B.n279 B.n146 163.367
R1859 B.n283 B.n146 163.367
R1860 B.n284 B.n283 163.367
R1861 B.n285 B.n284 163.367
R1862 B.n285 B.n144 163.367
R1863 B.n289 B.n144 163.367
R1864 B.n290 B.n289 163.367
R1865 B.n291 B.n290 163.367
R1866 B.n291 B.n142 163.367
R1867 B.n295 B.n142 163.367
R1868 B.n296 B.n295 163.367
R1869 B.n297 B.n296 163.367
R1870 B.n297 B.n138 163.367
R1871 B.n302 B.n138 163.367
R1872 B.n303 B.n302 163.367
R1873 B.n304 B.n303 163.367
R1874 B.n304 B.n136 163.367
R1875 B.n308 B.n136 163.367
R1876 B.n309 B.n308 163.367
R1877 B.n310 B.n309 163.367
R1878 B.n310 B.n134 163.367
R1879 B.n317 B.n134 163.367
R1880 B.n318 B.n317 163.367
R1881 B.n319 B.n318 163.367
R1882 B.n319 B.n132 163.367
R1883 B.n323 B.n132 163.367
R1884 B.n324 B.n323 163.367
R1885 B.n325 B.n324 163.367
R1886 B.n325 B.n130 163.367
R1887 B.n329 B.n130 163.367
R1888 B.n330 B.n329 163.367
R1889 B.n331 B.n330 163.367
R1890 B.n331 B.n128 163.367
R1891 B.n335 B.n128 163.367
R1892 B.n336 B.n335 163.367
R1893 B.n337 B.n336 163.367
R1894 B.n337 B.n126 163.367
R1895 B.n341 B.n126 163.367
R1896 B.n342 B.n341 163.367
R1897 B.n343 B.n342 163.367
R1898 B.n343 B.n124 163.367
R1899 B.n347 B.n124 163.367
R1900 B.n348 B.n347 163.367
R1901 B.n349 B.n348 163.367
R1902 B.n349 B.n122 163.367
R1903 B.n353 B.n122 163.367
R1904 B.n354 B.n353 163.367
R1905 B.n355 B.n354 163.367
R1906 B.n355 B.n120 163.367
R1907 B.n359 B.n120 163.367
R1908 B.n360 B.n359 163.367
R1909 B.n361 B.n360 163.367
R1910 B.n361 B.n118 163.367
R1911 B.n365 B.n118 163.367
R1912 B.n366 B.n365 163.367
R1913 B.n367 B.n366 163.367
R1914 B.n367 B.n116 163.367
R1915 B.n371 B.n116 163.367
R1916 B.n372 B.n371 163.367
R1917 B.n373 B.n372 163.367
R1918 B.n373 B.n114 163.367
R1919 B.n377 B.n114 163.367
R1920 B.n378 B.n377 163.367
R1921 B.n379 B.n378 163.367
R1922 B.n379 B.n112 163.367
R1923 B.n383 B.n112 163.367
R1924 B.n384 B.n383 163.367
R1925 B.n385 B.n384 163.367
R1926 B.n385 B.n110 163.367
R1927 B.n389 B.n110 163.367
R1928 B.n390 B.n389 163.367
R1929 B.n391 B.n390 163.367
R1930 B.n391 B.n108 163.367
R1931 B.n395 B.n108 163.367
R1932 B.n396 B.n395 163.367
R1933 B.n397 B.n396 163.367
R1934 B.n397 B.n106 163.367
R1935 B.n401 B.n106 163.367
R1936 B.n402 B.n401 163.367
R1937 B.n403 B.n402 163.367
R1938 B.n403 B.n104 163.367
R1939 B.n407 B.n104 163.367
R1940 B.n408 B.n407 163.367
R1941 B.n409 B.n408 163.367
R1942 B.n409 B.n102 163.367
R1943 B.n413 B.n102 163.367
R1944 B.n415 B.n414 163.367
R1945 B.n415 B.n100 163.367
R1946 B.n419 B.n100 163.367
R1947 B.n420 B.n419 163.367
R1948 B.n421 B.n420 163.367
R1949 B.n421 B.n98 163.367
R1950 B.n425 B.n98 163.367
R1951 B.n426 B.n425 163.367
R1952 B.n427 B.n426 163.367
R1953 B.n427 B.n96 163.367
R1954 B.n431 B.n96 163.367
R1955 B.n432 B.n431 163.367
R1956 B.n433 B.n432 163.367
R1957 B.n433 B.n94 163.367
R1958 B.n437 B.n94 163.367
R1959 B.n438 B.n437 163.367
R1960 B.n439 B.n438 163.367
R1961 B.n439 B.n92 163.367
R1962 B.n443 B.n92 163.367
R1963 B.n444 B.n443 163.367
R1964 B.n445 B.n444 163.367
R1965 B.n445 B.n90 163.367
R1966 B.n449 B.n90 163.367
R1967 B.n450 B.n449 163.367
R1968 B.n451 B.n450 163.367
R1969 B.n451 B.n88 163.367
R1970 B.n455 B.n88 163.367
R1971 B.n456 B.n455 163.367
R1972 B.n457 B.n456 163.367
R1973 B.n457 B.n86 163.367
R1974 B.n461 B.n86 163.367
R1975 B.n462 B.n461 163.367
R1976 B.n463 B.n462 163.367
R1977 B.n463 B.n84 163.367
R1978 B.n672 B.n11 163.367
R1979 B.n668 B.n11 163.367
R1980 B.n668 B.n667 163.367
R1981 B.n667 B.n666 163.367
R1982 B.n666 B.n13 163.367
R1983 B.n662 B.n13 163.367
R1984 B.n662 B.n661 163.367
R1985 B.n661 B.n660 163.367
R1986 B.n660 B.n15 163.367
R1987 B.n656 B.n15 163.367
R1988 B.n656 B.n655 163.367
R1989 B.n655 B.n654 163.367
R1990 B.n654 B.n17 163.367
R1991 B.n650 B.n17 163.367
R1992 B.n650 B.n649 163.367
R1993 B.n649 B.n648 163.367
R1994 B.n648 B.n19 163.367
R1995 B.n644 B.n19 163.367
R1996 B.n644 B.n643 163.367
R1997 B.n643 B.n642 163.367
R1998 B.n642 B.n21 163.367
R1999 B.n638 B.n21 163.367
R2000 B.n638 B.n637 163.367
R2001 B.n637 B.n636 163.367
R2002 B.n636 B.n23 163.367
R2003 B.n632 B.n23 163.367
R2004 B.n632 B.n631 163.367
R2005 B.n631 B.n630 163.367
R2006 B.n630 B.n25 163.367
R2007 B.n626 B.n25 163.367
R2008 B.n626 B.n625 163.367
R2009 B.n625 B.n624 163.367
R2010 B.n624 B.n27 163.367
R2011 B.n620 B.n27 163.367
R2012 B.n620 B.n619 163.367
R2013 B.n619 B.n618 163.367
R2014 B.n618 B.n29 163.367
R2015 B.n614 B.n29 163.367
R2016 B.n614 B.n613 163.367
R2017 B.n613 B.n612 163.367
R2018 B.n612 B.n31 163.367
R2019 B.n608 B.n31 163.367
R2020 B.n608 B.n607 163.367
R2021 B.n607 B.n606 163.367
R2022 B.n606 B.n33 163.367
R2023 B.n602 B.n33 163.367
R2024 B.n602 B.n601 163.367
R2025 B.n601 B.n600 163.367
R2026 B.n600 B.n35 163.367
R2027 B.n596 B.n35 163.367
R2028 B.n596 B.n595 163.367
R2029 B.n595 B.n594 163.367
R2030 B.n594 B.n37 163.367
R2031 B.n590 B.n37 163.367
R2032 B.n590 B.n589 163.367
R2033 B.n589 B.n588 163.367
R2034 B.n588 B.n39 163.367
R2035 B.n584 B.n39 163.367
R2036 B.n584 B.n583 163.367
R2037 B.n583 B.n582 163.367
R2038 B.n582 B.n41 163.367
R2039 B.n578 B.n41 163.367
R2040 B.n578 B.n577 163.367
R2041 B.n577 B.n576 163.367
R2042 B.n576 B.n43 163.367
R2043 B.n572 B.n43 163.367
R2044 B.n572 B.n571 163.367
R2045 B.n571 B.n570 163.367
R2046 B.n570 B.n48 163.367
R2047 B.n566 B.n48 163.367
R2048 B.n566 B.n565 163.367
R2049 B.n565 B.n564 163.367
R2050 B.n564 B.n50 163.367
R2051 B.n559 B.n50 163.367
R2052 B.n559 B.n558 163.367
R2053 B.n558 B.n557 163.367
R2054 B.n557 B.n54 163.367
R2055 B.n553 B.n54 163.367
R2056 B.n553 B.n552 163.367
R2057 B.n552 B.n551 163.367
R2058 B.n551 B.n56 163.367
R2059 B.n547 B.n56 163.367
R2060 B.n547 B.n546 163.367
R2061 B.n546 B.n545 163.367
R2062 B.n545 B.n58 163.367
R2063 B.n541 B.n58 163.367
R2064 B.n541 B.n540 163.367
R2065 B.n540 B.n539 163.367
R2066 B.n539 B.n60 163.367
R2067 B.n535 B.n60 163.367
R2068 B.n535 B.n534 163.367
R2069 B.n534 B.n533 163.367
R2070 B.n533 B.n62 163.367
R2071 B.n529 B.n62 163.367
R2072 B.n529 B.n528 163.367
R2073 B.n528 B.n527 163.367
R2074 B.n527 B.n64 163.367
R2075 B.n523 B.n64 163.367
R2076 B.n523 B.n522 163.367
R2077 B.n522 B.n521 163.367
R2078 B.n521 B.n66 163.367
R2079 B.n517 B.n66 163.367
R2080 B.n517 B.n516 163.367
R2081 B.n516 B.n515 163.367
R2082 B.n515 B.n68 163.367
R2083 B.n511 B.n68 163.367
R2084 B.n511 B.n510 163.367
R2085 B.n510 B.n509 163.367
R2086 B.n509 B.n70 163.367
R2087 B.n505 B.n70 163.367
R2088 B.n505 B.n504 163.367
R2089 B.n504 B.n503 163.367
R2090 B.n503 B.n72 163.367
R2091 B.n499 B.n72 163.367
R2092 B.n499 B.n498 163.367
R2093 B.n498 B.n497 163.367
R2094 B.n497 B.n74 163.367
R2095 B.n493 B.n74 163.367
R2096 B.n493 B.n492 163.367
R2097 B.n492 B.n491 163.367
R2098 B.n491 B.n76 163.367
R2099 B.n487 B.n76 163.367
R2100 B.n487 B.n486 163.367
R2101 B.n486 B.n485 163.367
R2102 B.n485 B.n78 163.367
R2103 B.n481 B.n78 163.367
R2104 B.n481 B.n480 163.367
R2105 B.n480 B.n479 163.367
R2106 B.n479 B.n80 163.367
R2107 B.n475 B.n80 163.367
R2108 B.n475 B.n474 163.367
R2109 B.n474 B.n473 163.367
R2110 B.n473 B.n82 163.367
R2111 B.n469 B.n82 163.367
R2112 B.n469 B.n468 163.367
R2113 B.n468 B.n467 163.367
R2114 B.n315 B.n314 59.5399
R2115 B.n300 B.n140 59.5399
R2116 B.n46 B.n45 59.5399
R2117 B.n562 B.n52 59.5399
R2118 B.n671 B.n10 32.6249
R2119 B.n466 B.n465 32.6249
R2120 B.n412 B.n101 32.6249
R2121 B.n204 B.n203 32.6249
R2122 B B.n699 18.0485
R2123 B.n671 B.n670 10.6151
R2124 B.n670 B.n669 10.6151
R2125 B.n669 B.n12 10.6151
R2126 B.n665 B.n12 10.6151
R2127 B.n665 B.n664 10.6151
R2128 B.n664 B.n663 10.6151
R2129 B.n663 B.n14 10.6151
R2130 B.n659 B.n14 10.6151
R2131 B.n659 B.n658 10.6151
R2132 B.n658 B.n657 10.6151
R2133 B.n657 B.n16 10.6151
R2134 B.n653 B.n16 10.6151
R2135 B.n653 B.n652 10.6151
R2136 B.n652 B.n651 10.6151
R2137 B.n651 B.n18 10.6151
R2138 B.n647 B.n18 10.6151
R2139 B.n647 B.n646 10.6151
R2140 B.n646 B.n645 10.6151
R2141 B.n645 B.n20 10.6151
R2142 B.n641 B.n20 10.6151
R2143 B.n641 B.n640 10.6151
R2144 B.n640 B.n639 10.6151
R2145 B.n639 B.n22 10.6151
R2146 B.n635 B.n22 10.6151
R2147 B.n635 B.n634 10.6151
R2148 B.n634 B.n633 10.6151
R2149 B.n633 B.n24 10.6151
R2150 B.n629 B.n24 10.6151
R2151 B.n629 B.n628 10.6151
R2152 B.n628 B.n627 10.6151
R2153 B.n627 B.n26 10.6151
R2154 B.n623 B.n26 10.6151
R2155 B.n623 B.n622 10.6151
R2156 B.n622 B.n621 10.6151
R2157 B.n621 B.n28 10.6151
R2158 B.n617 B.n28 10.6151
R2159 B.n617 B.n616 10.6151
R2160 B.n616 B.n615 10.6151
R2161 B.n615 B.n30 10.6151
R2162 B.n611 B.n30 10.6151
R2163 B.n611 B.n610 10.6151
R2164 B.n610 B.n609 10.6151
R2165 B.n609 B.n32 10.6151
R2166 B.n605 B.n32 10.6151
R2167 B.n605 B.n604 10.6151
R2168 B.n604 B.n603 10.6151
R2169 B.n603 B.n34 10.6151
R2170 B.n599 B.n34 10.6151
R2171 B.n599 B.n598 10.6151
R2172 B.n598 B.n597 10.6151
R2173 B.n597 B.n36 10.6151
R2174 B.n593 B.n36 10.6151
R2175 B.n593 B.n592 10.6151
R2176 B.n592 B.n591 10.6151
R2177 B.n591 B.n38 10.6151
R2178 B.n587 B.n38 10.6151
R2179 B.n587 B.n586 10.6151
R2180 B.n586 B.n585 10.6151
R2181 B.n585 B.n40 10.6151
R2182 B.n581 B.n40 10.6151
R2183 B.n581 B.n580 10.6151
R2184 B.n580 B.n579 10.6151
R2185 B.n579 B.n42 10.6151
R2186 B.n575 B.n574 10.6151
R2187 B.n574 B.n573 10.6151
R2188 B.n573 B.n47 10.6151
R2189 B.n569 B.n47 10.6151
R2190 B.n569 B.n568 10.6151
R2191 B.n568 B.n567 10.6151
R2192 B.n567 B.n49 10.6151
R2193 B.n563 B.n49 10.6151
R2194 B.n561 B.n560 10.6151
R2195 B.n560 B.n53 10.6151
R2196 B.n556 B.n53 10.6151
R2197 B.n556 B.n555 10.6151
R2198 B.n555 B.n554 10.6151
R2199 B.n554 B.n55 10.6151
R2200 B.n550 B.n55 10.6151
R2201 B.n550 B.n549 10.6151
R2202 B.n549 B.n548 10.6151
R2203 B.n548 B.n57 10.6151
R2204 B.n544 B.n57 10.6151
R2205 B.n544 B.n543 10.6151
R2206 B.n543 B.n542 10.6151
R2207 B.n542 B.n59 10.6151
R2208 B.n538 B.n59 10.6151
R2209 B.n538 B.n537 10.6151
R2210 B.n537 B.n536 10.6151
R2211 B.n536 B.n61 10.6151
R2212 B.n532 B.n61 10.6151
R2213 B.n532 B.n531 10.6151
R2214 B.n531 B.n530 10.6151
R2215 B.n530 B.n63 10.6151
R2216 B.n526 B.n63 10.6151
R2217 B.n526 B.n525 10.6151
R2218 B.n525 B.n524 10.6151
R2219 B.n524 B.n65 10.6151
R2220 B.n520 B.n65 10.6151
R2221 B.n520 B.n519 10.6151
R2222 B.n519 B.n518 10.6151
R2223 B.n518 B.n67 10.6151
R2224 B.n514 B.n67 10.6151
R2225 B.n514 B.n513 10.6151
R2226 B.n513 B.n512 10.6151
R2227 B.n512 B.n69 10.6151
R2228 B.n508 B.n69 10.6151
R2229 B.n508 B.n507 10.6151
R2230 B.n507 B.n506 10.6151
R2231 B.n506 B.n71 10.6151
R2232 B.n502 B.n71 10.6151
R2233 B.n502 B.n501 10.6151
R2234 B.n501 B.n500 10.6151
R2235 B.n500 B.n73 10.6151
R2236 B.n496 B.n73 10.6151
R2237 B.n496 B.n495 10.6151
R2238 B.n495 B.n494 10.6151
R2239 B.n494 B.n75 10.6151
R2240 B.n490 B.n75 10.6151
R2241 B.n490 B.n489 10.6151
R2242 B.n489 B.n488 10.6151
R2243 B.n488 B.n77 10.6151
R2244 B.n484 B.n77 10.6151
R2245 B.n484 B.n483 10.6151
R2246 B.n483 B.n482 10.6151
R2247 B.n482 B.n79 10.6151
R2248 B.n478 B.n79 10.6151
R2249 B.n478 B.n477 10.6151
R2250 B.n477 B.n476 10.6151
R2251 B.n476 B.n81 10.6151
R2252 B.n472 B.n81 10.6151
R2253 B.n472 B.n471 10.6151
R2254 B.n471 B.n470 10.6151
R2255 B.n470 B.n83 10.6151
R2256 B.n466 B.n83 10.6151
R2257 B.n416 B.n101 10.6151
R2258 B.n417 B.n416 10.6151
R2259 B.n418 B.n417 10.6151
R2260 B.n418 B.n99 10.6151
R2261 B.n422 B.n99 10.6151
R2262 B.n423 B.n422 10.6151
R2263 B.n424 B.n423 10.6151
R2264 B.n424 B.n97 10.6151
R2265 B.n428 B.n97 10.6151
R2266 B.n429 B.n428 10.6151
R2267 B.n430 B.n429 10.6151
R2268 B.n430 B.n95 10.6151
R2269 B.n434 B.n95 10.6151
R2270 B.n435 B.n434 10.6151
R2271 B.n436 B.n435 10.6151
R2272 B.n436 B.n93 10.6151
R2273 B.n440 B.n93 10.6151
R2274 B.n441 B.n440 10.6151
R2275 B.n442 B.n441 10.6151
R2276 B.n442 B.n91 10.6151
R2277 B.n446 B.n91 10.6151
R2278 B.n447 B.n446 10.6151
R2279 B.n448 B.n447 10.6151
R2280 B.n448 B.n89 10.6151
R2281 B.n452 B.n89 10.6151
R2282 B.n453 B.n452 10.6151
R2283 B.n454 B.n453 10.6151
R2284 B.n454 B.n87 10.6151
R2285 B.n458 B.n87 10.6151
R2286 B.n459 B.n458 10.6151
R2287 B.n460 B.n459 10.6151
R2288 B.n460 B.n85 10.6151
R2289 B.n464 B.n85 10.6151
R2290 B.n465 B.n464 10.6151
R2291 B.n204 B.n171 10.6151
R2292 B.n208 B.n171 10.6151
R2293 B.n209 B.n208 10.6151
R2294 B.n210 B.n209 10.6151
R2295 B.n210 B.n169 10.6151
R2296 B.n214 B.n169 10.6151
R2297 B.n215 B.n214 10.6151
R2298 B.n216 B.n215 10.6151
R2299 B.n216 B.n167 10.6151
R2300 B.n220 B.n167 10.6151
R2301 B.n221 B.n220 10.6151
R2302 B.n222 B.n221 10.6151
R2303 B.n222 B.n165 10.6151
R2304 B.n226 B.n165 10.6151
R2305 B.n227 B.n226 10.6151
R2306 B.n228 B.n227 10.6151
R2307 B.n228 B.n163 10.6151
R2308 B.n232 B.n163 10.6151
R2309 B.n233 B.n232 10.6151
R2310 B.n234 B.n233 10.6151
R2311 B.n234 B.n161 10.6151
R2312 B.n238 B.n161 10.6151
R2313 B.n239 B.n238 10.6151
R2314 B.n240 B.n239 10.6151
R2315 B.n240 B.n159 10.6151
R2316 B.n244 B.n159 10.6151
R2317 B.n245 B.n244 10.6151
R2318 B.n246 B.n245 10.6151
R2319 B.n246 B.n157 10.6151
R2320 B.n250 B.n157 10.6151
R2321 B.n251 B.n250 10.6151
R2322 B.n252 B.n251 10.6151
R2323 B.n252 B.n155 10.6151
R2324 B.n256 B.n155 10.6151
R2325 B.n257 B.n256 10.6151
R2326 B.n258 B.n257 10.6151
R2327 B.n258 B.n153 10.6151
R2328 B.n262 B.n153 10.6151
R2329 B.n263 B.n262 10.6151
R2330 B.n264 B.n263 10.6151
R2331 B.n264 B.n151 10.6151
R2332 B.n268 B.n151 10.6151
R2333 B.n269 B.n268 10.6151
R2334 B.n270 B.n269 10.6151
R2335 B.n270 B.n149 10.6151
R2336 B.n274 B.n149 10.6151
R2337 B.n275 B.n274 10.6151
R2338 B.n276 B.n275 10.6151
R2339 B.n276 B.n147 10.6151
R2340 B.n280 B.n147 10.6151
R2341 B.n281 B.n280 10.6151
R2342 B.n282 B.n281 10.6151
R2343 B.n282 B.n145 10.6151
R2344 B.n286 B.n145 10.6151
R2345 B.n287 B.n286 10.6151
R2346 B.n288 B.n287 10.6151
R2347 B.n288 B.n143 10.6151
R2348 B.n292 B.n143 10.6151
R2349 B.n293 B.n292 10.6151
R2350 B.n294 B.n293 10.6151
R2351 B.n294 B.n141 10.6151
R2352 B.n298 B.n141 10.6151
R2353 B.n299 B.n298 10.6151
R2354 B.n301 B.n137 10.6151
R2355 B.n305 B.n137 10.6151
R2356 B.n306 B.n305 10.6151
R2357 B.n307 B.n306 10.6151
R2358 B.n307 B.n135 10.6151
R2359 B.n311 B.n135 10.6151
R2360 B.n312 B.n311 10.6151
R2361 B.n316 B.n312 10.6151
R2362 B.n320 B.n133 10.6151
R2363 B.n321 B.n320 10.6151
R2364 B.n322 B.n321 10.6151
R2365 B.n322 B.n131 10.6151
R2366 B.n326 B.n131 10.6151
R2367 B.n327 B.n326 10.6151
R2368 B.n328 B.n327 10.6151
R2369 B.n328 B.n129 10.6151
R2370 B.n332 B.n129 10.6151
R2371 B.n333 B.n332 10.6151
R2372 B.n334 B.n333 10.6151
R2373 B.n334 B.n127 10.6151
R2374 B.n338 B.n127 10.6151
R2375 B.n339 B.n338 10.6151
R2376 B.n340 B.n339 10.6151
R2377 B.n340 B.n125 10.6151
R2378 B.n344 B.n125 10.6151
R2379 B.n345 B.n344 10.6151
R2380 B.n346 B.n345 10.6151
R2381 B.n346 B.n123 10.6151
R2382 B.n350 B.n123 10.6151
R2383 B.n351 B.n350 10.6151
R2384 B.n352 B.n351 10.6151
R2385 B.n352 B.n121 10.6151
R2386 B.n356 B.n121 10.6151
R2387 B.n357 B.n356 10.6151
R2388 B.n358 B.n357 10.6151
R2389 B.n358 B.n119 10.6151
R2390 B.n362 B.n119 10.6151
R2391 B.n363 B.n362 10.6151
R2392 B.n364 B.n363 10.6151
R2393 B.n364 B.n117 10.6151
R2394 B.n368 B.n117 10.6151
R2395 B.n369 B.n368 10.6151
R2396 B.n370 B.n369 10.6151
R2397 B.n370 B.n115 10.6151
R2398 B.n374 B.n115 10.6151
R2399 B.n375 B.n374 10.6151
R2400 B.n376 B.n375 10.6151
R2401 B.n376 B.n113 10.6151
R2402 B.n380 B.n113 10.6151
R2403 B.n381 B.n380 10.6151
R2404 B.n382 B.n381 10.6151
R2405 B.n382 B.n111 10.6151
R2406 B.n386 B.n111 10.6151
R2407 B.n387 B.n386 10.6151
R2408 B.n388 B.n387 10.6151
R2409 B.n388 B.n109 10.6151
R2410 B.n392 B.n109 10.6151
R2411 B.n393 B.n392 10.6151
R2412 B.n394 B.n393 10.6151
R2413 B.n394 B.n107 10.6151
R2414 B.n398 B.n107 10.6151
R2415 B.n399 B.n398 10.6151
R2416 B.n400 B.n399 10.6151
R2417 B.n400 B.n105 10.6151
R2418 B.n404 B.n105 10.6151
R2419 B.n405 B.n404 10.6151
R2420 B.n406 B.n405 10.6151
R2421 B.n406 B.n103 10.6151
R2422 B.n410 B.n103 10.6151
R2423 B.n411 B.n410 10.6151
R2424 B.n412 B.n411 10.6151
R2425 B.n203 B.n202 10.6151
R2426 B.n202 B.n173 10.6151
R2427 B.n198 B.n173 10.6151
R2428 B.n198 B.n197 10.6151
R2429 B.n197 B.n196 10.6151
R2430 B.n196 B.n175 10.6151
R2431 B.n192 B.n175 10.6151
R2432 B.n192 B.n191 10.6151
R2433 B.n191 B.n190 10.6151
R2434 B.n190 B.n177 10.6151
R2435 B.n186 B.n177 10.6151
R2436 B.n186 B.n185 10.6151
R2437 B.n185 B.n184 10.6151
R2438 B.n184 B.n179 10.6151
R2439 B.n180 B.n179 10.6151
R2440 B.n180 B.n0 10.6151
R2441 B.n695 B.n1 10.6151
R2442 B.n695 B.n694 10.6151
R2443 B.n694 B.n693 10.6151
R2444 B.n693 B.n4 10.6151
R2445 B.n689 B.n4 10.6151
R2446 B.n689 B.n688 10.6151
R2447 B.n688 B.n687 10.6151
R2448 B.n687 B.n6 10.6151
R2449 B.n683 B.n6 10.6151
R2450 B.n683 B.n682 10.6151
R2451 B.n682 B.n681 10.6151
R2452 B.n681 B.n8 10.6151
R2453 B.n677 B.n8 10.6151
R2454 B.n677 B.n676 10.6151
R2455 B.n676 B.n675 10.6151
R2456 B.n675 B.n10 10.6151
R2457 B.n314 B.n313 9.69747
R2458 B.n140 B.n139 9.69747
R2459 B.n45 B.n44 9.69747
R2460 B.n52 B.n51 9.69747
R2461 B.n575 B.n46 6.5566
R2462 B.n563 B.n562 6.5566
R2463 B.n301 B.n300 6.5566
R2464 B.n316 B.n315 6.5566
R2465 B.n46 B.n42 4.05904
R2466 B.n562 B.n561 4.05904
R2467 B.n300 B.n299 4.05904
R2468 B.n315 B.n133 4.05904
R2469 B.n699 B.n0 2.81026
R2470 B.n699 B.n1 2.81026
C0 w_n1570_n4876# B 8.6526f
C1 w_n1570_n4876# VP 2.97018f
C2 VDD1 B 1.98729f
C3 VDD1 VP 4.38655f
C4 VDD2 B 2.01152f
C5 VTAIL B 3.52678f
C6 VDD2 VP 0.275576f
C7 VTAIL VP 3.46168f
C8 VDD1 w_n1570_n4876# 2.35654f
C9 VN B 0.749987f
C10 VDD2 w_n1570_n4876# 2.37417f
C11 VN VP 6.2126f
C12 VTAIL w_n1570_n4876# 4.29832f
C13 VDD1 VDD2 0.648268f
C14 VTAIL VDD1 41.6426f
C15 VN w_n1570_n4876# 2.77327f
C16 VTAIL VDD2 41.6647f
C17 VN VDD1 0.147658f
C18 VN VDD2 4.26735f
C19 VN VTAIL 3.44641f
C20 B VP 1.06769f
C21 VDD2 VSUBS 1.836212f
C22 VDD1 VSUBS 1.203128f
C23 VTAIL VSUBS 0.557132f
C24 VN VSUBS 5.43446f
C25 VP VSUBS 1.431552f
C26 B VSUBS 2.97674f
C27 w_n1570_n4876# VSUBS 93.5029f
C28 B.n0 VSUBS 0.005467f
C29 B.n1 VSUBS 0.005467f
C30 B.n2 VSUBS 0.008645f
C31 B.n3 VSUBS 0.008645f
C32 B.n4 VSUBS 0.008645f
C33 B.n5 VSUBS 0.008645f
C34 B.n6 VSUBS 0.008645f
C35 B.n7 VSUBS 0.008645f
C36 B.n8 VSUBS 0.008645f
C37 B.n9 VSUBS 0.008645f
C38 B.n10 VSUBS 0.019852f
C39 B.n11 VSUBS 0.008645f
C40 B.n12 VSUBS 0.008645f
C41 B.n13 VSUBS 0.008645f
C42 B.n14 VSUBS 0.008645f
C43 B.n15 VSUBS 0.008645f
C44 B.n16 VSUBS 0.008645f
C45 B.n17 VSUBS 0.008645f
C46 B.n18 VSUBS 0.008645f
C47 B.n19 VSUBS 0.008645f
C48 B.n20 VSUBS 0.008645f
C49 B.n21 VSUBS 0.008645f
C50 B.n22 VSUBS 0.008645f
C51 B.n23 VSUBS 0.008645f
C52 B.n24 VSUBS 0.008645f
C53 B.n25 VSUBS 0.008645f
C54 B.n26 VSUBS 0.008645f
C55 B.n27 VSUBS 0.008645f
C56 B.n28 VSUBS 0.008645f
C57 B.n29 VSUBS 0.008645f
C58 B.n30 VSUBS 0.008645f
C59 B.n31 VSUBS 0.008645f
C60 B.n32 VSUBS 0.008645f
C61 B.n33 VSUBS 0.008645f
C62 B.n34 VSUBS 0.008645f
C63 B.n35 VSUBS 0.008645f
C64 B.n36 VSUBS 0.008645f
C65 B.n37 VSUBS 0.008645f
C66 B.n38 VSUBS 0.008645f
C67 B.n39 VSUBS 0.008645f
C68 B.n40 VSUBS 0.008645f
C69 B.n41 VSUBS 0.008645f
C70 B.n42 VSUBS 0.005975f
C71 B.n43 VSUBS 0.008645f
C72 B.t11 VSUBS 0.479844f
C73 B.t10 VSUBS 0.487355f
C74 B.t9 VSUBS 0.156618f
C75 B.n44 VSUBS 0.457414f
C76 B.n45 VSUBS 0.416005f
C77 B.n46 VSUBS 0.020029f
C78 B.n47 VSUBS 0.008645f
C79 B.n48 VSUBS 0.008645f
C80 B.n49 VSUBS 0.008645f
C81 B.n50 VSUBS 0.008645f
C82 B.t2 VSUBS 0.479848f
C83 B.t1 VSUBS 0.48736f
C84 B.t0 VSUBS 0.156618f
C85 B.n51 VSUBS 0.45741f
C86 B.n52 VSUBS 0.416f
C87 B.n53 VSUBS 0.008645f
C88 B.n54 VSUBS 0.008645f
C89 B.n55 VSUBS 0.008645f
C90 B.n56 VSUBS 0.008645f
C91 B.n57 VSUBS 0.008645f
C92 B.n58 VSUBS 0.008645f
C93 B.n59 VSUBS 0.008645f
C94 B.n60 VSUBS 0.008645f
C95 B.n61 VSUBS 0.008645f
C96 B.n62 VSUBS 0.008645f
C97 B.n63 VSUBS 0.008645f
C98 B.n64 VSUBS 0.008645f
C99 B.n65 VSUBS 0.008645f
C100 B.n66 VSUBS 0.008645f
C101 B.n67 VSUBS 0.008645f
C102 B.n68 VSUBS 0.008645f
C103 B.n69 VSUBS 0.008645f
C104 B.n70 VSUBS 0.008645f
C105 B.n71 VSUBS 0.008645f
C106 B.n72 VSUBS 0.008645f
C107 B.n73 VSUBS 0.008645f
C108 B.n74 VSUBS 0.008645f
C109 B.n75 VSUBS 0.008645f
C110 B.n76 VSUBS 0.008645f
C111 B.n77 VSUBS 0.008645f
C112 B.n78 VSUBS 0.008645f
C113 B.n79 VSUBS 0.008645f
C114 B.n80 VSUBS 0.008645f
C115 B.n81 VSUBS 0.008645f
C116 B.n82 VSUBS 0.008645f
C117 B.n83 VSUBS 0.008645f
C118 B.n84 VSUBS 0.019852f
C119 B.n85 VSUBS 0.008645f
C120 B.n86 VSUBS 0.008645f
C121 B.n87 VSUBS 0.008645f
C122 B.n88 VSUBS 0.008645f
C123 B.n89 VSUBS 0.008645f
C124 B.n90 VSUBS 0.008645f
C125 B.n91 VSUBS 0.008645f
C126 B.n92 VSUBS 0.008645f
C127 B.n93 VSUBS 0.008645f
C128 B.n94 VSUBS 0.008645f
C129 B.n95 VSUBS 0.008645f
C130 B.n96 VSUBS 0.008645f
C131 B.n97 VSUBS 0.008645f
C132 B.n98 VSUBS 0.008645f
C133 B.n99 VSUBS 0.008645f
C134 B.n100 VSUBS 0.008645f
C135 B.n101 VSUBS 0.019852f
C136 B.n102 VSUBS 0.008645f
C137 B.n103 VSUBS 0.008645f
C138 B.n104 VSUBS 0.008645f
C139 B.n105 VSUBS 0.008645f
C140 B.n106 VSUBS 0.008645f
C141 B.n107 VSUBS 0.008645f
C142 B.n108 VSUBS 0.008645f
C143 B.n109 VSUBS 0.008645f
C144 B.n110 VSUBS 0.008645f
C145 B.n111 VSUBS 0.008645f
C146 B.n112 VSUBS 0.008645f
C147 B.n113 VSUBS 0.008645f
C148 B.n114 VSUBS 0.008645f
C149 B.n115 VSUBS 0.008645f
C150 B.n116 VSUBS 0.008645f
C151 B.n117 VSUBS 0.008645f
C152 B.n118 VSUBS 0.008645f
C153 B.n119 VSUBS 0.008645f
C154 B.n120 VSUBS 0.008645f
C155 B.n121 VSUBS 0.008645f
C156 B.n122 VSUBS 0.008645f
C157 B.n123 VSUBS 0.008645f
C158 B.n124 VSUBS 0.008645f
C159 B.n125 VSUBS 0.008645f
C160 B.n126 VSUBS 0.008645f
C161 B.n127 VSUBS 0.008645f
C162 B.n128 VSUBS 0.008645f
C163 B.n129 VSUBS 0.008645f
C164 B.n130 VSUBS 0.008645f
C165 B.n131 VSUBS 0.008645f
C166 B.n132 VSUBS 0.008645f
C167 B.n133 VSUBS 0.005975f
C168 B.n134 VSUBS 0.008645f
C169 B.n135 VSUBS 0.008645f
C170 B.n136 VSUBS 0.008645f
C171 B.n137 VSUBS 0.008645f
C172 B.n138 VSUBS 0.008645f
C173 B.t4 VSUBS 0.479844f
C174 B.t5 VSUBS 0.487355f
C175 B.t3 VSUBS 0.156618f
C176 B.n139 VSUBS 0.457414f
C177 B.n140 VSUBS 0.416005f
C178 B.n141 VSUBS 0.008645f
C179 B.n142 VSUBS 0.008645f
C180 B.n143 VSUBS 0.008645f
C181 B.n144 VSUBS 0.008645f
C182 B.n145 VSUBS 0.008645f
C183 B.n146 VSUBS 0.008645f
C184 B.n147 VSUBS 0.008645f
C185 B.n148 VSUBS 0.008645f
C186 B.n149 VSUBS 0.008645f
C187 B.n150 VSUBS 0.008645f
C188 B.n151 VSUBS 0.008645f
C189 B.n152 VSUBS 0.008645f
C190 B.n153 VSUBS 0.008645f
C191 B.n154 VSUBS 0.008645f
C192 B.n155 VSUBS 0.008645f
C193 B.n156 VSUBS 0.008645f
C194 B.n157 VSUBS 0.008645f
C195 B.n158 VSUBS 0.008645f
C196 B.n159 VSUBS 0.008645f
C197 B.n160 VSUBS 0.008645f
C198 B.n161 VSUBS 0.008645f
C199 B.n162 VSUBS 0.008645f
C200 B.n163 VSUBS 0.008645f
C201 B.n164 VSUBS 0.008645f
C202 B.n165 VSUBS 0.008645f
C203 B.n166 VSUBS 0.008645f
C204 B.n167 VSUBS 0.008645f
C205 B.n168 VSUBS 0.008645f
C206 B.n169 VSUBS 0.008645f
C207 B.n170 VSUBS 0.008645f
C208 B.n171 VSUBS 0.008645f
C209 B.n172 VSUBS 0.019852f
C210 B.n173 VSUBS 0.008645f
C211 B.n174 VSUBS 0.008645f
C212 B.n175 VSUBS 0.008645f
C213 B.n176 VSUBS 0.008645f
C214 B.n177 VSUBS 0.008645f
C215 B.n178 VSUBS 0.008645f
C216 B.n179 VSUBS 0.008645f
C217 B.n180 VSUBS 0.008645f
C218 B.n181 VSUBS 0.008645f
C219 B.n182 VSUBS 0.008645f
C220 B.n183 VSUBS 0.008645f
C221 B.n184 VSUBS 0.008645f
C222 B.n185 VSUBS 0.008645f
C223 B.n186 VSUBS 0.008645f
C224 B.n187 VSUBS 0.008645f
C225 B.n188 VSUBS 0.008645f
C226 B.n189 VSUBS 0.008645f
C227 B.n190 VSUBS 0.008645f
C228 B.n191 VSUBS 0.008645f
C229 B.n192 VSUBS 0.008645f
C230 B.n193 VSUBS 0.008645f
C231 B.n194 VSUBS 0.008645f
C232 B.n195 VSUBS 0.008645f
C233 B.n196 VSUBS 0.008645f
C234 B.n197 VSUBS 0.008645f
C235 B.n198 VSUBS 0.008645f
C236 B.n199 VSUBS 0.008645f
C237 B.n200 VSUBS 0.008645f
C238 B.n201 VSUBS 0.008645f
C239 B.n202 VSUBS 0.008645f
C240 B.n203 VSUBS 0.019852f
C241 B.n204 VSUBS 0.020575f
C242 B.n205 VSUBS 0.020575f
C243 B.n206 VSUBS 0.008645f
C244 B.n207 VSUBS 0.008645f
C245 B.n208 VSUBS 0.008645f
C246 B.n209 VSUBS 0.008645f
C247 B.n210 VSUBS 0.008645f
C248 B.n211 VSUBS 0.008645f
C249 B.n212 VSUBS 0.008645f
C250 B.n213 VSUBS 0.008645f
C251 B.n214 VSUBS 0.008645f
C252 B.n215 VSUBS 0.008645f
C253 B.n216 VSUBS 0.008645f
C254 B.n217 VSUBS 0.008645f
C255 B.n218 VSUBS 0.008645f
C256 B.n219 VSUBS 0.008645f
C257 B.n220 VSUBS 0.008645f
C258 B.n221 VSUBS 0.008645f
C259 B.n222 VSUBS 0.008645f
C260 B.n223 VSUBS 0.008645f
C261 B.n224 VSUBS 0.008645f
C262 B.n225 VSUBS 0.008645f
C263 B.n226 VSUBS 0.008645f
C264 B.n227 VSUBS 0.008645f
C265 B.n228 VSUBS 0.008645f
C266 B.n229 VSUBS 0.008645f
C267 B.n230 VSUBS 0.008645f
C268 B.n231 VSUBS 0.008645f
C269 B.n232 VSUBS 0.008645f
C270 B.n233 VSUBS 0.008645f
C271 B.n234 VSUBS 0.008645f
C272 B.n235 VSUBS 0.008645f
C273 B.n236 VSUBS 0.008645f
C274 B.n237 VSUBS 0.008645f
C275 B.n238 VSUBS 0.008645f
C276 B.n239 VSUBS 0.008645f
C277 B.n240 VSUBS 0.008645f
C278 B.n241 VSUBS 0.008645f
C279 B.n242 VSUBS 0.008645f
C280 B.n243 VSUBS 0.008645f
C281 B.n244 VSUBS 0.008645f
C282 B.n245 VSUBS 0.008645f
C283 B.n246 VSUBS 0.008645f
C284 B.n247 VSUBS 0.008645f
C285 B.n248 VSUBS 0.008645f
C286 B.n249 VSUBS 0.008645f
C287 B.n250 VSUBS 0.008645f
C288 B.n251 VSUBS 0.008645f
C289 B.n252 VSUBS 0.008645f
C290 B.n253 VSUBS 0.008645f
C291 B.n254 VSUBS 0.008645f
C292 B.n255 VSUBS 0.008645f
C293 B.n256 VSUBS 0.008645f
C294 B.n257 VSUBS 0.008645f
C295 B.n258 VSUBS 0.008645f
C296 B.n259 VSUBS 0.008645f
C297 B.n260 VSUBS 0.008645f
C298 B.n261 VSUBS 0.008645f
C299 B.n262 VSUBS 0.008645f
C300 B.n263 VSUBS 0.008645f
C301 B.n264 VSUBS 0.008645f
C302 B.n265 VSUBS 0.008645f
C303 B.n266 VSUBS 0.008645f
C304 B.n267 VSUBS 0.008645f
C305 B.n268 VSUBS 0.008645f
C306 B.n269 VSUBS 0.008645f
C307 B.n270 VSUBS 0.008645f
C308 B.n271 VSUBS 0.008645f
C309 B.n272 VSUBS 0.008645f
C310 B.n273 VSUBS 0.008645f
C311 B.n274 VSUBS 0.008645f
C312 B.n275 VSUBS 0.008645f
C313 B.n276 VSUBS 0.008645f
C314 B.n277 VSUBS 0.008645f
C315 B.n278 VSUBS 0.008645f
C316 B.n279 VSUBS 0.008645f
C317 B.n280 VSUBS 0.008645f
C318 B.n281 VSUBS 0.008645f
C319 B.n282 VSUBS 0.008645f
C320 B.n283 VSUBS 0.008645f
C321 B.n284 VSUBS 0.008645f
C322 B.n285 VSUBS 0.008645f
C323 B.n286 VSUBS 0.008645f
C324 B.n287 VSUBS 0.008645f
C325 B.n288 VSUBS 0.008645f
C326 B.n289 VSUBS 0.008645f
C327 B.n290 VSUBS 0.008645f
C328 B.n291 VSUBS 0.008645f
C329 B.n292 VSUBS 0.008645f
C330 B.n293 VSUBS 0.008645f
C331 B.n294 VSUBS 0.008645f
C332 B.n295 VSUBS 0.008645f
C333 B.n296 VSUBS 0.008645f
C334 B.n297 VSUBS 0.008645f
C335 B.n298 VSUBS 0.008645f
C336 B.n299 VSUBS 0.005975f
C337 B.n300 VSUBS 0.020029f
C338 B.n301 VSUBS 0.006992f
C339 B.n302 VSUBS 0.008645f
C340 B.n303 VSUBS 0.008645f
C341 B.n304 VSUBS 0.008645f
C342 B.n305 VSUBS 0.008645f
C343 B.n306 VSUBS 0.008645f
C344 B.n307 VSUBS 0.008645f
C345 B.n308 VSUBS 0.008645f
C346 B.n309 VSUBS 0.008645f
C347 B.n310 VSUBS 0.008645f
C348 B.n311 VSUBS 0.008645f
C349 B.n312 VSUBS 0.008645f
C350 B.t7 VSUBS 0.479848f
C351 B.t8 VSUBS 0.48736f
C352 B.t6 VSUBS 0.156618f
C353 B.n313 VSUBS 0.45741f
C354 B.n314 VSUBS 0.416f
C355 B.n315 VSUBS 0.020029f
C356 B.n316 VSUBS 0.006992f
C357 B.n317 VSUBS 0.008645f
C358 B.n318 VSUBS 0.008645f
C359 B.n319 VSUBS 0.008645f
C360 B.n320 VSUBS 0.008645f
C361 B.n321 VSUBS 0.008645f
C362 B.n322 VSUBS 0.008645f
C363 B.n323 VSUBS 0.008645f
C364 B.n324 VSUBS 0.008645f
C365 B.n325 VSUBS 0.008645f
C366 B.n326 VSUBS 0.008645f
C367 B.n327 VSUBS 0.008645f
C368 B.n328 VSUBS 0.008645f
C369 B.n329 VSUBS 0.008645f
C370 B.n330 VSUBS 0.008645f
C371 B.n331 VSUBS 0.008645f
C372 B.n332 VSUBS 0.008645f
C373 B.n333 VSUBS 0.008645f
C374 B.n334 VSUBS 0.008645f
C375 B.n335 VSUBS 0.008645f
C376 B.n336 VSUBS 0.008645f
C377 B.n337 VSUBS 0.008645f
C378 B.n338 VSUBS 0.008645f
C379 B.n339 VSUBS 0.008645f
C380 B.n340 VSUBS 0.008645f
C381 B.n341 VSUBS 0.008645f
C382 B.n342 VSUBS 0.008645f
C383 B.n343 VSUBS 0.008645f
C384 B.n344 VSUBS 0.008645f
C385 B.n345 VSUBS 0.008645f
C386 B.n346 VSUBS 0.008645f
C387 B.n347 VSUBS 0.008645f
C388 B.n348 VSUBS 0.008645f
C389 B.n349 VSUBS 0.008645f
C390 B.n350 VSUBS 0.008645f
C391 B.n351 VSUBS 0.008645f
C392 B.n352 VSUBS 0.008645f
C393 B.n353 VSUBS 0.008645f
C394 B.n354 VSUBS 0.008645f
C395 B.n355 VSUBS 0.008645f
C396 B.n356 VSUBS 0.008645f
C397 B.n357 VSUBS 0.008645f
C398 B.n358 VSUBS 0.008645f
C399 B.n359 VSUBS 0.008645f
C400 B.n360 VSUBS 0.008645f
C401 B.n361 VSUBS 0.008645f
C402 B.n362 VSUBS 0.008645f
C403 B.n363 VSUBS 0.008645f
C404 B.n364 VSUBS 0.008645f
C405 B.n365 VSUBS 0.008645f
C406 B.n366 VSUBS 0.008645f
C407 B.n367 VSUBS 0.008645f
C408 B.n368 VSUBS 0.008645f
C409 B.n369 VSUBS 0.008645f
C410 B.n370 VSUBS 0.008645f
C411 B.n371 VSUBS 0.008645f
C412 B.n372 VSUBS 0.008645f
C413 B.n373 VSUBS 0.008645f
C414 B.n374 VSUBS 0.008645f
C415 B.n375 VSUBS 0.008645f
C416 B.n376 VSUBS 0.008645f
C417 B.n377 VSUBS 0.008645f
C418 B.n378 VSUBS 0.008645f
C419 B.n379 VSUBS 0.008645f
C420 B.n380 VSUBS 0.008645f
C421 B.n381 VSUBS 0.008645f
C422 B.n382 VSUBS 0.008645f
C423 B.n383 VSUBS 0.008645f
C424 B.n384 VSUBS 0.008645f
C425 B.n385 VSUBS 0.008645f
C426 B.n386 VSUBS 0.008645f
C427 B.n387 VSUBS 0.008645f
C428 B.n388 VSUBS 0.008645f
C429 B.n389 VSUBS 0.008645f
C430 B.n390 VSUBS 0.008645f
C431 B.n391 VSUBS 0.008645f
C432 B.n392 VSUBS 0.008645f
C433 B.n393 VSUBS 0.008645f
C434 B.n394 VSUBS 0.008645f
C435 B.n395 VSUBS 0.008645f
C436 B.n396 VSUBS 0.008645f
C437 B.n397 VSUBS 0.008645f
C438 B.n398 VSUBS 0.008645f
C439 B.n399 VSUBS 0.008645f
C440 B.n400 VSUBS 0.008645f
C441 B.n401 VSUBS 0.008645f
C442 B.n402 VSUBS 0.008645f
C443 B.n403 VSUBS 0.008645f
C444 B.n404 VSUBS 0.008645f
C445 B.n405 VSUBS 0.008645f
C446 B.n406 VSUBS 0.008645f
C447 B.n407 VSUBS 0.008645f
C448 B.n408 VSUBS 0.008645f
C449 B.n409 VSUBS 0.008645f
C450 B.n410 VSUBS 0.008645f
C451 B.n411 VSUBS 0.008645f
C452 B.n412 VSUBS 0.020575f
C453 B.n413 VSUBS 0.020575f
C454 B.n414 VSUBS 0.019852f
C455 B.n415 VSUBS 0.008645f
C456 B.n416 VSUBS 0.008645f
C457 B.n417 VSUBS 0.008645f
C458 B.n418 VSUBS 0.008645f
C459 B.n419 VSUBS 0.008645f
C460 B.n420 VSUBS 0.008645f
C461 B.n421 VSUBS 0.008645f
C462 B.n422 VSUBS 0.008645f
C463 B.n423 VSUBS 0.008645f
C464 B.n424 VSUBS 0.008645f
C465 B.n425 VSUBS 0.008645f
C466 B.n426 VSUBS 0.008645f
C467 B.n427 VSUBS 0.008645f
C468 B.n428 VSUBS 0.008645f
C469 B.n429 VSUBS 0.008645f
C470 B.n430 VSUBS 0.008645f
C471 B.n431 VSUBS 0.008645f
C472 B.n432 VSUBS 0.008645f
C473 B.n433 VSUBS 0.008645f
C474 B.n434 VSUBS 0.008645f
C475 B.n435 VSUBS 0.008645f
C476 B.n436 VSUBS 0.008645f
C477 B.n437 VSUBS 0.008645f
C478 B.n438 VSUBS 0.008645f
C479 B.n439 VSUBS 0.008645f
C480 B.n440 VSUBS 0.008645f
C481 B.n441 VSUBS 0.008645f
C482 B.n442 VSUBS 0.008645f
C483 B.n443 VSUBS 0.008645f
C484 B.n444 VSUBS 0.008645f
C485 B.n445 VSUBS 0.008645f
C486 B.n446 VSUBS 0.008645f
C487 B.n447 VSUBS 0.008645f
C488 B.n448 VSUBS 0.008645f
C489 B.n449 VSUBS 0.008645f
C490 B.n450 VSUBS 0.008645f
C491 B.n451 VSUBS 0.008645f
C492 B.n452 VSUBS 0.008645f
C493 B.n453 VSUBS 0.008645f
C494 B.n454 VSUBS 0.008645f
C495 B.n455 VSUBS 0.008645f
C496 B.n456 VSUBS 0.008645f
C497 B.n457 VSUBS 0.008645f
C498 B.n458 VSUBS 0.008645f
C499 B.n459 VSUBS 0.008645f
C500 B.n460 VSUBS 0.008645f
C501 B.n461 VSUBS 0.008645f
C502 B.n462 VSUBS 0.008645f
C503 B.n463 VSUBS 0.008645f
C504 B.n464 VSUBS 0.008645f
C505 B.n465 VSUBS 0.020875f
C506 B.n466 VSUBS 0.019553f
C507 B.n467 VSUBS 0.020575f
C508 B.n468 VSUBS 0.008645f
C509 B.n469 VSUBS 0.008645f
C510 B.n470 VSUBS 0.008645f
C511 B.n471 VSUBS 0.008645f
C512 B.n472 VSUBS 0.008645f
C513 B.n473 VSUBS 0.008645f
C514 B.n474 VSUBS 0.008645f
C515 B.n475 VSUBS 0.008645f
C516 B.n476 VSUBS 0.008645f
C517 B.n477 VSUBS 0.008645f
C518 B.n478 VSUBS 0.008645f
C519 B.n479 VSUBS 0.008645f
C520 B.n480 VSUBS 0.008645f
C521 B.n481 VSUBS 0.008645f
C522 B.n482 VSUBS 0.008645f
C523 B.n483 VSUBS 0.008645f
C524 B.n484 VSUBS 0.008645f
C525 B.n485 VSUBS 0.008645f
C526 B.n486 VSUBS 0.008645f
C527 B.n487 VSUBS 0.008645f
C528 B.n488 VSUBS 0.008645f
C529 B.n489 VSUBS 0.008645f
C530 B.n490 VSUBS 0.008645f
C531 B.n491 VSUBS 0.008645f
C532 B.n492 VSUBS 0.008645f
C533 B.n493 VSUBS 0.008645f
C534 B.n494 VSUBS 0.008645f
C535 B.n495 VSUBS 0.008645f
C536 B.n496 VSUBS 0.008645f
C537 B.n497 VSUBS 0.008645f
C538 B.n498 VSUBS 0.008645f
C539 B.n499 VSUBS 0.008645f
C540 B.n500 VSUBS 0.008645f
C541 B.n501 VSUBS 0.008645f
C542 B.n502 VSUBS 0.008645f
C543 B.n503 VSUBS 0.008645f
C544 B.n504 VSUBS 0.008645f
C545 B.n505 VSUBS 0.008645f
C546 B.n506 VSUBS 0.008645f
C547 B.n507 VSUBS 0.008645f
C548 B.n508 VSUBS 0.008645f
C549 B.n509 VSUBS 0.008645f
C550 B.n510 VSUBS 0.008645f
C551 B.n511 VSUBS 0.008645f
C552 B.n512 VSUBS 0.008645f
C553 B.n513 VSUBS 0.008645f
C554 B.n514 VSUBS 0.008645f
C555 B.n515 VSUBS 0.008645f
C556 B.n516 VSUBS 0.008645f
C557 B.n517 VSUBS 0.008645f
C558 B.n518 VSUBS 0.008645f
C559 B.n519 VSUBS 0.008645f
C560 B.n520 VSUBS 0.008645f
C561 B.n521 VSUBS 0.008645f
C562 B.n522 VSUBS 0.008645f
C563 B.n523 VSUBS 0.008645f
C564 B.n524 VSUBS 0.008645f
C565 B.n525 VSUBS 0.008645f
C566 B.n526 VSUBS 0.008645f
C567 B.n527 VSUBS 0.008645f
C568 B.n528 VSUBS 0.008645f
C569 B.n529 VSUBS 0.008645f
C570 B.n530 VSUBS 0.008645f
C571 B.n531 VSUBS 0.008645f
C572 B.n532 VSUBS 0.008645f
C573 B.n533 VSUBS 0.008645f
C574 B.n534 VSUBS 0.008645f
C575 B.n535 VSUBS 0.008645f
C576 B.n536 VSUBS 0.008645f
C577 B.n537 VSUBS 0.008645f
C578 B.n538 VSUBS 0.008645f
C579 B.n539 VSUBS 0.008645f
C580 B.n540 VSUBS 0.008645f
C581 B.n541 VSUBS 0.008645f
C582 B.n542 VSUBS 0.008645f
C583 B.n543 VSUBS 0.008645f
C584 B.n544 VSUBS 0.008645f
C585 B.n545 VSUBS 0.008645f
C586 B.n546 VSUBS 0.008645f
C587 B.n547 VSUBS 0.008645f
C588 B.n548 VSUBS 0.008645f
C589 B.n549 VSUBS 0.008645f
C590 B.n550 VSUBS 0.008645f
C591 B.n551 VSUBS 0.008645f
C592 B.n552 VSUBS 0.008645f
C593 B.n553 VSUBS 0.008645f
C594 B.n554 VSUBS 0.008645f
C595 B.n555 VSUBS 0.008645f
C596 B.n556 VSUBS 0.008645f
C597 B.n557 VSUBS 0.008645f
C598 B.n558 VSUBS 0.008645f
C599 B.n559 VSUBS 0.008645f
C600 B.n560 VSUBS 0.008645f
C601 B.n561 VSUBS 0.005975f
C602 B.n562 VSUBS 0.020029f
C603 B.n563 VSUBS 0.006992f
C604 B.n564 VSUBS 0.008645f
C605 B.n565 VSUBS 0.008645f
C606 B.n566 VSUBS 0.008645f
C607 B.n567 VSUBS 0.008645f
C608 B.n568 VSUBS 0.008645f
C609 B.n569 VSUBS 0.008645f
C610 B.n570 VSUBS 0.008645f
C611 B.n571 VSUBS 0.008645f
C612 B.n572 VSUBS 0.008645f
C613 B.n573 VSUBS 0.008645f
C614 B.n574 VSUBS 0.008645f
C615 B.n575 VSUBS 0.006992f
C616 B.n576 VSUBS 0.008645f
C617 B.n577 VSUBS 0.008645f
C618 B.n578 VSUBS 0.008645f
C619 B.n579 VSUBS 0.008645f
C620 B.n580 VSUBS 0.008645f
C621 B.n581 VSUBS 0.008645f
C622 B.n582 VSUBS 0.008645f
C623 B.n583 VSUBS 0.008645f
C624 B.n584 VSUBS 0.008645f
C625 B.n585 VSUBS 0.008645f
C626 B.n586 VSUBS 0.008645f
C627 B.n587 VSUBS 0.008645f
C628 B.n588 VSUBS 0.008645f
C629 B.n589 VSUBS 0.008645f
C630 B.n590 VSUBS 0.008645f
C631 B.n591 VSUBS 0.008645f
C632 B.n592 VSUBS 0.008645f
C633 B.n593 VSUBS 0.008645f
C634 B.n594 VSUBS 0.008645f
C635 B.n595 VSUBS 0.008645f
C636 B.n596 VSUBS 0.008645f
C637 B.n597 VSUBS 0.008645f
C638 B.n598 VSUBS 0.008645f
C639 B.n599 VSUBS 0.008645f
C640 B.n600 VSUBS 0.008645f
C641 B.n601 VSUBS 0.008645f
C642 B.n602 VSUBS 0.008645f
C643 B.n603 VSUBS 0.008645f
C644 B.n604 VSUBS 0.008645f
C645 B.n605 VSUBS 0.008645f
C646 B.n606 VSUBS 0.008645f
C647 B.n607 VSUBS 0.008645f
C648 B.n608 VSUBS 0.008645f
C649 B.n609 VSUBS 0.008645f
C650 B.n610 VSUBS 0.008645f
C651 B.n611 VSUBS 0.008645f
C652 B.n612 VSUBS 0.008645f
C653 B.n613 VSUBS 0.008645f
C654 B.n614 VSUBS 0.008645f
C655 B.n615 VSUBS 0.008645f
C656 B.n616 VSUBS 0.008645f
C657 B.n617 VSUBS 0.008645f
C658 B.n618 VSUBS 0.008645f
C659 B.n619 VSUBS 0.008645f
C660 B.n620 VSUBS 0.008645f
C661 B.n621 VSUBS 0.008645f
C662 B.n622 VSUBS 0.008645f
C663 B.n623 VSUBS 0.008645f
C664 B.n624 VSUBS 0.008645f
C665 B.n625 VSUBS 0.008645f
C666 B.n626 VSUBS 0.008645f
C667 B.n627 VSUBS 0.008645f
C668 B.n628 VSUBS 0.008645f
C669 B.n629 VSUBS 0.008645f
C670 B.n630 VSUBS 0.008645f
C671 B.n631 VSUBS 0.008645f
C672 B.n632 VSUBS 0.008645f
C673 B.n633 VSUBS 0.008645f
C674 B.n634 VSUBS 0.008645f
C675 B.n635 VSUBS 0.008645f
C676 B.n636 VSUBS 0.008645f
C677 B.n637 VSUBS 0.008645f
C678 B.n638 VSUBS 0.008645f
C679 B.n639 VSUBS 0.008645f
C680 B.n640 VSUBS 0.008645f
C681 B.n641 VSUBS 0.008645f
C682 B.n642 VSUBS 0.008645f
C683 B.n643 VSUBS 0.008645f
C684 B.n644 VSUBS 0.008645f
C685 B.n645 VSUBS 0.008645f
C686 B.n646 VSUBS 0.008645f
C687 B.n647 VSUBS 0.008645f
C688 B.n648 VSUBS 0.008645f
C689 B.n649 VSUBS 0.008645f
C690 B.n650 VSUBS 0.008645f
C691 B.n651 VSUBS 0.008645f
C692 B.n652 VSUBS 0.008645f
C693 B.n653 VSUBS 0.008645f
C694 B.n654 VSUBS 0.008645f
C695 B.n655 VSUBS 0.008645f
C696 B.n656 VSUBS 0.008645f
C697 B.n657 VSUBS 0.008645f
C698 B.n658 VSUBS 0.008645f
C699 B.n659 VSUBS 0.008645f
C700 B.n660 VSUBS 0.008645f
C701 B.n661 VSUBS 0.008645f
C702 B.n662 VSUBS 0.008645f
C703 B.n663 VSUBS 0.008645f
C704 B.n664 VSUBS 0.008645f
C705 B.n665 VSUBS 0.008645f
C706 B.n666 VSUBS 0.008645f
C707 B.n667 VSUBS 0.008645f
C708 B.n668 VSUBS 0.008645f
C709 B.n669 VSUBS 0.008645f
C710 B.n670 VSUBS 0.008645f
C711 B.n671 VSUBS 0.020575f
C712 B.n672 VSUBS 0.020575f
C713 B.n673 VSUBS 0.019852f
C714 B.n674 VSUBS 0.008645f
C715 B.n675 VSUBS 0.008645f
C716 B.n676 VSUBS 0.008645f
C717 B.n677 VSUBS 0.008645f
C718 B.n678 VSUBS 0.008645f
C719 B.n679 VSUBS 0.008645f
C720 B.n680 VSUBS 0.008645f
C721 B.n681 VSUBS 0.008645f
C722 B.n682 VSUBS 0.008645f
C723 B.n683 VSUBS 0.008645f
C724 B.n684 VSUBS 0.008645f
C725 B.n685 VSUBS 0.008645f
C726 B.n686 VSUBS 0.008645f
C727 B.n687 VSUBS 0.008645f
C728 B.n688 VSUBS 0.008645f
C729 B.n689 VSUBS 0.008645f
C730 B.n690 VSUBS 0.008645f
C731 B.n691 VSUBS 0.008645f
C732 B.n692 VSUBS 0.008645f
C733 B.n693 VSUBS 0.008645f
C734 B.n694 VSUBS 0.008645f
C735 B.n695 VSUBS 0.008645f
C736 B.n696 VSUBS 0.008645f
C737 B.n697 VSUBS 0.008645f
C738 B.n698 VSUBS 0.008645f
C739 B.n699 VSUBS 0.019575f
C740 VDD1.n0 VSUBS 0.041655f
C741 VDD1.n1 VSUBS 0.037439f
C742 VDD1.n2 VSUBS 0.020118f
C743 VDD1.n3 VSUBS 0.047552f
C744 VDD1.n4 VSUBS 0.021301f
C745 VDD1.n5 VSUBS 0.037439f
C746 VDD1.n6 VSUBS 0.020118f
C747 VDD1.n7 VSUBS 0.047552f
C748 VDD1.n8 VSUBS 0.021301f
C749 VDD1.n9 VSUBS 0.037439f
C750 VDD1.n10 VSUBS 0.020118f
C751 VDD1.n11 VSUBS 0.047552f
C752 VDD1.n12 VSUBS 0.021301f
C753 VDD1.n13 VSUBS 0.037439f
C754 VDD1.n14 VSUBS 0.020118f
C755 VDD1.n15 VSUBS 0.047552f
C756 VDD1.n16 VSUBS 0.021301f
C757 VDD1.n17 VSUBS 0.037439f
C758 VDD1.n18 VSUBS 0.020118f
C759 VDD1.n19 VSUBS 0.047552f
C760 VDD1.n20 VSUBS 0.021301f
C761 VDD1.n21 VSUBS 0.037439f
C762 VDD1.n22 VSUBS 0.020118f
C763 VDD1.n23 VSUBS 0.047552f
C764 VDD1.n24 VSUBS 0.021301f
C765 VDD1.n25 VSUBS 0.037439f
C766 VDD1.n26 VSUBS 0.020118f
C767 VDD1.n27 VSUBS 0.047552f
C768 VDD1.n28 VSUBS 0.047552f
C769 VDD1.n29 VSUBS 0.021301f
C770 VDD1.n30 VSUBS 0.037439f
C771 VDD1.n31 VSUBS 0.020118f
C772 VDD1.n32 VSUBS 0.047552f
C773 VDD1.n33 VSUBS 0.021301f
C774 VDD1.n34 VSUBS 0.422491f
C775 VDD1.t8 VSUBS 0.103422f
C776 VDD1.n35 VSUBS 0.035664f
C777 VDD1.n36 VSUBS 0.035771f
C778 VDD1.n37 VSUBS 0.020118f
C779 VDD1.n38 VSUBS 3.07637f
C780 VDD1.n39 VSUBS 0.037439f
C781 VDD1.n40 VSUBS 0.020118f
C782 VDD1.n41 VSUBS 0.021301f
C783 VDD1.n42 VSUBS 0.047552f
C784 VDD1.n43 VSUBS 0.047552f
C785 VDD1.n44 VSUBS 0.021301f
C786 VDD1.n45 VSUBS 0.020118f
C787 VDD1.n46 VSUBS 0.037439f
C788 VDD1.n47 VSUBS 0.037439f
C789 VDD1.n48 VSUBS 0.020118f
C790 VDD1.n49 VSUBS 0.021301f
C791 VDD1.n50 VSUBS 0.047552f
C792 VDD1.n51 VSUBS 0.047552f
C793 VDD1.n52 VSUBS 0.021301f
C794 VDD1.n53 VSUBS 0.020118f
C795 VDD1.n54 VSUBS 0.037439f
C796 VDD1.n55 VSUBS 0.037439f
C797 VDD1.n56 VSUBS 0.020118f
C798 VDD1.n57 VSUBS 0.02071f
C799 VDD1.n58 VSUBS 0.02071f
C800 VDD1.n59 VSUBS 0.047552f
C801 VDD1.n60 VSUBS 0.047552f
C802 VDD1.n61 VSUBS 0.021301f
C803 VDD1.n62 VSUBS 0.020118f
C804 VDD1.n63 VSUBS 0.037439f
C805 VDD1.n64 VSUBS 0.037439f
C806 VDD1.n65 VSUBS 0.020118f
C807 VDD1.n66 VSUBS 0.021301f
C808 VDD1.n67 VSUBS 0.047552f
C809 VDD1.n68 VSUBS 0.047552f
C810 VDD1.n69 VSUBS 0.021301f
C811 VDD1.n70 VSUBS 0.020118f
C812 VDD1.n71 VSUBS 0.037439f
C813 VDD1.n72 VSUBS 0.037439f
C814 VDD1.n73 VSUBS 0.020118f
C815 VDD1.n74 VSUBS 0.021301f
C816 VDD1.n75 VSUBS 0.047552f
C817 VDD1.n76 VSUBS 0.047552f
C818 VDD1.n77 VSUBS 0.021301f
C819 VDD1.n78 VSUBS 0.020118f
C820 VDD1.n79 VSUBS 0.037439f
C821 VDD1.n80 VSUBS 0.037439f
C822 VDD1.n81 VSUBS 0.020118f
C823 VDD1.n82 VSUBS 0.021301f
C824 VDD1.n83 VSUBS 0.047552f
C825 VDD1.n84 VSUBS 0.047552f
C826 VDD1.n85 VSUBS 0.021301f
C827 VDD1.n86 VSUBS 0.020118f
C828 VDD1.n87 VSUBS 0.037439f
C829 VDD1.n88 VSUBS 0.037439f
C830 VDD1.n89 VSUBS 0.020118f
C831 VDD1.n90 VSUBS 0.021301f
C832 VDD1.n91 VSUBS 0.047552f
C833 VDD1.n92 VSUBS 0.047552f
C834 VDD1.n93 VSUBS 0.021301f
C835 VDD1.n94 VSUBS 0.020118f
C836 VDD1.n95 VSUBS 0.037439f
C837 VDD1.n96 VSUBS 0.037439f
C838 VDD1.n97 VSUBS 0.020118f
C839 VDD1.n98 VSUBS 0.021301f
C840 VDD1.n99 VSUBS 0.047552f
C841 VDD1.n100 VSUBS 0.120531f
C842 VDD1.n101 VSUBS 0.021301f
C843 VDD1.n102 VSUBS 0.039507f
C844 VDD1.n103 VSUBS 0.09779f
C845 VDD1.n104 VSUBS 0.12044f
C846 VDD1.t0 VSUBS 0.578095f
C847 VDD1.t4 VSUBS 0.578095f
C848 VDD1.n105 VSUBS 4.88813f
C849 VDD1.n106 VSUBS 0.909297f
C850 VDD1.n107 VSUBS 0.041655f
C851 VDD1.n108 VSUBS 0.037439f
C852 VDD1.n109 VSUBS 0.020118f
C853 VDD1.n110 VSUBS 0.047552f
C854 VDD1.n111 VSUBS 0.021301f
C855 VDD1.n112 VSUBS 0.037439f
C856 VDD1.n113 VSUBS 0.020118f
C857 VDD1.n114 VSUBS 0.047552f
C858 VDD1.n115 VSUBS 0.021301f
C859 VDD1.n116 VSUBS 0.037439f
C860 VDD1.n117 VSUBS 0.020118f
C861 VDD1.n118 VSUBS 0.047552f
C862 VDD1.n119 VSUBS 0.021301f
C863 VDD1.n120 VSUBS 0.037439f
C864 VDD1.n121 VSUBS 0.020118f
C865 VDD1.n122 VSUBS 0.047552f
C866 VDD1.n123 VSUBS 0.021301f
C867 VDD1.n124 VSUBS 0.037439f
C868 VDD1.n125 VSUBS 0.020118f
C869 VDD1.n126 VSUBS 0.047552f
C870 VDD1.n127 VSUBS 0.021301f
C871 VDD1.n128 VSUBS 0.037439f
C872 VDD1.n129 VSUBS 0.020118f
C873 VDD1.n130 VSUBS 0.047552f
C874 VDD1.n131 VSUBS 0.021301f
C875 VDD1.n132 VSUBS 0.037439f
C876 VDD1.n133 VSUBS 0.020118f
C877 VDD1.n134 VSUBS 0.047552f
C878 VDD1.n135 VSUBS 0.021301f
C879 VDD1.n136 VSUBS 0.037439f
C880 VDD1.n137 VSUBS 0.020118f
C881 VDD1.n138 VSUBS 0.047552f
C882 VDD1.n139 VSUBS 0.021301f
C883 VDD1.n140 VSUBS 0.422491f
C884 VDD1.t6 VSUBS 0.103422f
C885 VDD1.n141 VSUBS 0.035664f
C886 VDD1.n142 VSUBS 0.035771f
C887 VDD1.n143 VSUBS 0.020118f
C888 VDD1.n144 VSUBS 3.07637f
C889 VDD1.n145 VSUBS 0.037439f
C890 VDD1.n146 VSUBS 0.020118f
C891 VDD1.n147 VSUBS 0.021301f
C892 VDD1.n148 VSUBS 0.047552f
C893 VDD1.n149 VSUBS 0.047552f
C894 VDD1.n150 VSUBS 0.021301f
C895 VDD1.n151 VSUBS 0.020118f
C896 VDD1.n152 VSUBS 0.037439f
C897 VDD1.n153 VSUBS 0.037439f
C898 VDD1.n154 VSUBS 0.020118f
C899 VDD1.n155 VSUBS 0.021301f
C900 VDD1.n156 VSUBS 0.047552f
C901 VDD1.n157 VSUBS 0.047552f
C902 VDD1.n158 VSUBS 0.047552f
C903 VDD1.n159 VSUBS 0.021301f
C904 VDD1.n160 VSUBS 0.020118f
C905 VDD1.n161 VSUBS 0.037439f
C906 VDD1.n162 VSUBS 0.037439f
C907 VDD1.n163 VSUBS 0.020118f
C908 VDD1.n164 VSUBS 0.02071f
C909 VDD1.n165 VSUBS 0.02071f
C910 VDD1.n166 VSUBS 0.047552f
C911 VDD1.n167 VSUBS 0.047552f
C912 VDD1.n168 VSUBS 0.021301f
C913 VDD1.n169 VSUBS 0.020118f
C914 VDD1.n170 VSUBS 0.037439f
C915 VDD1.n171 VSUBS 0.037439f
C916 VDD1.n172 VSUBS 0.020118f
C917 VDD1.n173 VSUBS 0.021301f
C918 VDD1.n174 VSUBS 0.047552f
C919 VDD1.n175 VSUBS 0.047552f
C920 VDD1.n176 VSUBS 0.021301f
C921 VDD1.n177 VSUBS 0.020118f
C922 VDD1.n178 VSUBS 0.037439f
C923 VDD1.n179 VSUBS 0.037439f
C924 VDD1.n180 VSUBS 0.020118f
C925 VDD1.n181 VSUBS 0.021301f
C926 VDD1.n182 VSUBS 0.047552f
C927 VDD1.n183 VSUBS 0.047552f
C928 VDD1.n184 VSUBS 0.021301f
C929 VDD1.n185 VSUBS 0.020118f
C930 VDD1.n186 VSUBS 0.037439f
C931 VDD1.n187 VSUBS 0.037439f
C932 VDD1.n188 VSUBS 0.020118f
C933 VDD1.n189 VSUBS 0.021301f
C934 VDD1.n190 VSUBS 0.047552f
C935 VDD1.n191 VSUBS 0.047552f
C936 VDD1.n192 VSUBS 0.021301f
C937 VDD1.n193 VSUBS 0.020118f
C938 VDD1.n194 VSUBS 0.037439f
C939 VDD1.n195 VSUBS 0.037439f
C940 VDD1.n196 VSUBS 0.020118f
C941 VDD1.n197 VSUBS 0.021301f
C942 VDD1.n198 VSUBS 0.047552f
C943 VDD1.n199 VSUBS 0.047552f
C944 VDD1.n200 VSUBS 0.021301f
C945 VDD1.n201 VSUBS 0.020118f
C946 VDD1.n202 VSUBS 0.037439f
C947 VDD1.n203 VSUBS 0.037439f
C948 VDD1.n204 VSUBS 0.020118f
C949 VDD1.n205 VSUBS 0.021301f
C950 VDD1.n206 VSUBS 0.047552f
C951 VDD1.n207 VSUBS 0.120531f
C952 VDD1.n208 VSUBS 0.021301f
C953 VDD1.n209 VSUBS 0.039507f
C954 VDD1.n210 VSUBS 0.09779f
C955 VDD1.n211 VSUBS 0.12044f
C956 VDD1.t5 VSUBS 0.578095f
C957 VDD1.t3 VSUBS 0.578095f
C958 VDD1.n212 VSUBS 4.88812f
C959 VDD1.n213 VSUBS 0.912181f
C960 VDD1.t2 VSUBS 0.578095f
C961 VDD1.t1 VSUBS 0.578095f
C962 VDD1.n214 VSUBS 4.89112f
C963 VDD1.n215 VSUBS 3.61176f
C964 VDD1.t7 VSUBS 0.578095f
C965 VDD1.t9 VSUBS 0.578095f
C966 VDD1.n216 VSUBS 4.88811f
C967 VDD1.n217 VSUBS 4.51423f
C968 VP.n0 VSUBS 0.07319f
C969 VP.t7 VSUBS 0.684833f
C970 VP.t6 VSUBS 0.684833f
C971 VP.t4 VSUBS 0.684833f
C972 VP.n1 VSUBS 0.264788f
C973 VP.n2 VSUBS 0.07319f
C974 VP.t2 VSUBS 0.684833f
C975 VP.t5 VSUBS 0.684833f
C976 VP.t9 VSUBS 0.684833f
C977 VP.n3 VSUBS 0.264788f
C978 VP.t1 VSUBS 0.688022f
C979 VP.n4 VSUBS 0.282364f
C980 VP.n5 VSUBS 0.153957f
C981 VP.n6 VSUBS 0.02428f
C982 VP.n7 VSUBS 0.264788f
C983 VP.n8 VSUBS 0.02428f
C984 VP.n9 VSUBS 0.264788f
C985 VP.t0 VSUBS 0.688022f
C986 VP.n10 VSUBS 0.282269f
C987 VP.n11 VSUBS 3.45584f
C988 VP.t3 VSUBS 0.688022f
C989 VP.n12 VSUBS 0.282269f
C990 VP.n13 VSUBS 3.51366f
C991 VP.n14 VSUBS 0.07319f
C992 VP.n15 VSUBS 0.02428f
C993 VP.n16 VSUBS 0.264788f
C994 VP.n17 VSUBS 0.02428f
C995 VP.n18 VSUBS 0.264788f
C996 VP.t8 VSUBS 0.688022f
C997 VP.n19 VSUBS 0.282269f
C998 VP.n20 VSUBS 0.05672f
C999 VTAIL.t11 VSUBS 0.604407f
C1000 VTAIL.t13 VSUBS 0.604407f
C1001 VTAIL.n0 VSUBS 4.89016f
C1002 VTAIL.n1 VSUBS 1.04181f
C1003 VTAIL.n2 VSUBS 0.04355f
C1004 VTAIL.n3 VSUBS 0.039143f
C1005 VTAIL.n4 VSUBS 0.021034f
C1006 VTAIL.n5 VSUBS 0.049716f
C1007 VTAIL.n6 VSUBS 0.022271f
C1008 VTAIL.n7 VSUBS 0.039143f
C1009 VTAIL.n8 VSUBS 0.021034f
C1010 VTAIL.n9 VSUBS 0.049716f
C1011 VTAIL.n10 VSUBS 0.022271f
C1012 VTAIL.n11 VSUBS 0.039143f
C1013 VTAIL.n12 VSUBS 0.021034f
C1014 VTAIL.n13 VSUBS 0.049716f
C1015 VTAIL.n14 VSUBS 0.022271f
C1016 VTAIL.n15 VSUBS 0.039143f
C1017 VTAIL.n16 VSUBS 0.021034f
C1018 VTAIL.n17 VSUBS 0.049716f
C1019 VTAIL.n18 VSUBS 0.022271f
C1020 VTAIL.n19 VSUBS 0.039143f
C1021 VTAIL.n20 VSUBS 0.021034f
C1022 VTAIL.n21 VSUBS 0.049716f
C1023 VTAIL.n22 VSUBS 0.022271f
C1024 VTAIL.n23 VSUBS 0.039143f
C1025 VTAIL.n24 VSUBS 0.021034f
C1026 VTAIL.n25 VSUBS 0.049716f
C1027 VTAIL.n26 VSUBS 0.022271f
C1028 VTAIL.n27 VSUBS 0.039143f
C1029 VTAIL.n28 VSUBS 0.021034f
C1030 VTAIL.n29 VSUBS 0.049716f
C1031 VTAIL.n30 VSUBS 0.022271f
C1032 VTAIL.n31 VSUBS 0.039143f
C1033 VTAIL.n32 VSUBS 0.021034f
C1034 VTAIL.n33 VSUBS 0.049716f
C1035 VTAIL.n34 VSUBS 0.022271f
C1036 VTAIL.n35 VSUBS 0.44172f
C1037 VTAIL.t6 VSUBS 0.10813f
C1038 VTAIL.n36 VSUBS 0.037287f
C1039 VTAIL.n37 VSUBS 0.037399f
C1040 VTAIL.n38 VSUBS 0.021034f
C1041 VTAIL.n39 VSUBS 3.21638f
C1042 VTAIL.n40 VSUBS 0.039143f
C1043 VTAIL.n41 VSUBS 0.021034f
C1044 VTAIL.n42 VSUBS 0.022271f
C1045 VTAIL.n43 VSUBS 0.049716f
C1046 VTAIL.n44 VSUBS 0.049716f
C1047 VTAIL.n45 VSUBS 0.022271f
C1048 VTAIL.n46 VSUBS 0.021034f
C1049 VTAIL.n47 VSUBS 0.039143f
C1050 VTAIL.n48 VSUBS 0.039143f
C1051 VTAIL.n49 VSUBS 0.021034f
C1052 VTAIL.n50 VSUBS 0.022271f
C1053 VTAIL.n51 VSUBS 0.049716f
C1054 VTAIL.n52 VSUBS 0.049716f
C1055 VTAIL.n53 VSUBS 0.049716f
C1056 VTAIL.n54 VSUBS 0.022271f
C1057 VTAIL.n55 VSUBS 0.021034f
C1058 VTAIL.n56 VSUBS 0.039143f
C1059 VTAIL.n57 VSUBS 0.039143f
C1060 VTAIL.n58 VSUBS 0.021034f
C1061 VTAIL.n59 VSUBS 0.021652f
C1062 VTAIL.n60 VSUBS 0.021652f
C1063 VTAIL.n61 VSUBS 0.049716f
C1064 VTAIL.n62 VSUBS 0.049716f
C1065 VTAIL.n63 VSUBS 0.022271f
C1066 VTAIL.n64 VSUBS 0.021034f
C1067 VTAIL.n65 VSUBS 0.039143f
C1068 VTAIL.n66 VSUBS 0.039143f
C1069 VTAIL.n67 VSUBS 0.021034f
C1070 VTAIL.n68 VSUBS 0.022271f
C1071 VTAIL.n69 VSUBS 0.049716f
C1072 VTAIL.n70 VSUBS 0.049716f
C1073 VTAIL.n71 VSUBS 0.022271f
C1074 VTAIL.n72 VSUBS 0.021034f
C1075 VTAIL.n73 VSUBS 0.039143f
C1076 VTAIL.n74 VSUBS 0.039143f
C1077 VTAIL.n75 VSUBS 0.021034f
C1078 VTAIL.n76 VSUBS 0.022271f
C1079 VTAIL.n77 VSUBS 0.049716f
C1080 VTAIL.n78 VSUBS 0.049716f
C1081 VTAIL.n79 VSUBS 0.022271f
C1082 VTAIL.n80 VSUBS 0.021034f
C1083 VTAIL.n81 VSUBS 0.039143f
C1084 VTAIL.n82 VSUBS 0.039143f
C1085 VTAIL.n83 VSUBS 0.021034f
C1086 VTAIL.n84 VSUBS 0.022271f
C1087 VTAIL.n85 VSUBS 0.049716f
C1088 VTAIL.n86 VSUBS 0.049716f
C1089 VTAIL.n87 VSUBS 0.022271f
C1090 VTAIL.n88 VSUBS 0.021034f
C1091 VTAIL.n89 VSUBS 0.039143f
C1092 VTAIL.n90 VSUBS 0.039143f
C1093 VTAIL.n91 VSUBS 0.021034f
C1094 VTAIL.n92 VSUBS 0.022271f
C1095 VTAIL.n93 VSUBS 0.049716f
C1096 VTAIL.n94 VSUBS 0.049716f
C1097 VTAIL.n95 VSUBS 0.022271f
C1098 VTAIL.n96 VSUBS 0.021034f
C1099 VTAIL.n97 VSUBS 0.039143f
C1100 VTAIL.n98 VSUBS 0.039143f
C1101 VTAIL.n99 VSUBS 0.021034f
C1102 VTAIL.n100 VSUBS 0.022271f
C1103 VTAIL.n101 VSUBS 0.049716f
C1104 VTAIL.n102 VSUBS 0.126017f
C1105 VTAIL.n103 VSUBS 0.022271f
C1106 VTAIL.n104 VSUBS 0.041305f
C1107 VTAIL.n105 VSUBS 0.102241f
C1108 VTAIL.n106 VSUBS 0.097877f
C1109 VTAIL.n107 VSUBS 0.180895f
C1110 VTAIL.t19 VSUBS 0.604407f
C1111 VTAIL.t17 VSUBS 0.604407f
C1112 VTAIL.n108 VSUBS 4.89016f
C1113 VTAIL.n109 VSUBS 1.01599f
C1114 VTAIL.t2 VSUBS 0.604407f
C1115 VTAIL.t1 VSUBS 0.604407f
C1116 VTAIL.n110 VSUBS 4.89016f
C1117 VTAIL.n111 VSUBS 3.72664f
C1118 VTAIL.t12 VSUBS 0.604407f
C1119 VTAIL.t9 VSUBS 0.604407f
C1120 VTAIL.n112 VSUBS 4.89019f
C1121 VTAIL.n113 VSUBS 3.72661f
C1122 VTAIL.t8 VSUBS 0.604407f
C1123 VTAIL.t14 VSUBS 0.604407f
C1124 VTAIL.n114 VSUBS 4.89019f
C1125 VTAIL.n115 VSUBS 1.01596f
C1126 VTAIL.n116 VSUBS 0.04355f
C1127 VTAIL.n117 VSUBS 0.039143f
C1128 VTAIL.n118 VSUBS 0.021034f
C1129 VTAIL.n119 VSUBS 0.049716f
C1130 VTAIL.n120 VSUBS 0.022271f
C1131 VTAIL.n121 VSUBS 0.039143f
C1132 VTAIL.n122 VSUBS 0.021034f
C1133 VTAIL.n123 VSUBS 0.049716f
C1134 VTAIL.n124 VSUBS 0.022271f
C1135 VTAIL.n125 VSUBS 0.039143f
C1136 VTAIL.n126 VSUBS 0.021034f
C1137 VTAIL.n127 VSUBS 0.049716f
C1138 VTAIL.n128 VSUBS 0.022271f
C1139 VTAIL.n129 VSUBS 0.039143f
C1140 VTAIL.n130 VSUBS 0.021034f
C1141 VTAIL.n131 VSUBS 0.049716f
C1142 VTAIL.n132 VSUBS 0.022271f
C1143 VTAIL.n133 VSUBS 0.039143f
C1144 VTAIL.n134 VSUBS 0.021034f
C1145 VTAIL.n135 VSUBS 0.049716f
C1146 VTAIL.n136 VSUBS 0.022271f
C1147 VTAIL.n137 VSUBS 0.039143f
C1148 VTAIL.n138 VSUBS 0.021034f
C1149 VTAIL.n139 VSUBS 0.049716f
C1150 VTAIL.n140 VSUBS 0.022271f
C1151 VTAIL.n141 VSUBS 0.039143f
C1152 VTAIL.n142 VSUBS 0.021034f
C1153 VTAIL.n143 VSUBS 0.049716f
C1154 VTAIL.n144 VSUBS 0.049716f
C1155 VTAIL.n145 VSUBS 0.022271f
C1156 VTAIL.n146 VSUBS 0.039143f
C1157 VTAIL.n147 VSUBS 0.021034f
C1158 VTAIL.n148 VSUBS 0.049716f
C1159 VTAIL.n149 VSUBS 0.022271f
C1160 VTAIL.n150 VSUBS 0.44172f
C1161 VTAIL.t10 VSUBS 0.10813f
C1162 VTAIL.n151 VSUBS 0.037287f
C1163 VTAIL.n152 VSUBS 0.037399f
C1164 VTAIL.n153 VSUBS 0.021034f
C1165 VTAIL.n154 VSUBS 3.21639f
C1166 VTAIL.n155 VSUBS 0.039143f
C1167 VTAIL.n156 VSUBS 0.021034f
C1168 VTAIL.n157 VSUBS 0.022271f
C1169 VTAIL.n158 VSUBS 0.049716f
C1170 VTAIL.n159 VSUBS 0.049716f
C1171 VTAIL.n160 VSUBS 0.022271f
C1172 VTAIL.n161 VSUBS 0.021034f
C1173 VTAIL.n162 VSUBS 0.039143f
C1174 VTAIL.n163 VSUBS 0.039143f
C1175 VTAIL.n164 VSUBS 0.021034f
C1176 VTAIL.n165 VSUBS 0.022271f
C1177 VTAIL.n166 VSUBS 0.049716f
C1178 VTAIL.n167 VSUBS 0.049716f
C1179 VTAIL.n168 VSUBS 0.022271f
C1180 VTAIL.n169 VSUBS 0.021034f
C1181 VTAIL.n170 VSUBS 0.039143f
C1182 VTAIL.n171 VSUBS 0.039143f
C1183 VTAIL.n172 VSUBS 0.021034f
C1184 VTAIL.n173 VSUBS 0.021652f
C1185 VTAIL.n174 VSUBS 0.021652f
C1186 VTAIL.n175 VSUBS 0.049716f
C1187 VTAIL.n176 VSUBS 0.049716f
C1188 VTAIL.n177 VSUBS 0.022271f
C1189 VTAIL.n178 VSUBS 0.021034f
C1190 VTAIL.n179 VSUBS 0.039143f
C1191 VTAIL.n180 VSUBS 0.039143f
C1192 VTAIL.n181 VSUBS 0.021034f
C1193 VTAIL.n182 VSUBS 0.022271f
C1194 VTAIL.n183 VSUBS 0.049716f
C1195 VTAIL.n184 VSUBS 0.049716f
C1196 VTAIL.n185 VSUBS 0.022271f
C1197 VTAIL.n186 VSUBS 0.021034f
C1198 VTAIL.n187 VSUBS 0.039143f
C1199 VTAIL.n188 VSUBS 0.039143f
C1200 VTAIL.n189 VSUBS 0.021034f
C1201 VTAIL.n190 VSUBS 0.022271f
C1202 VTAIL.n191 VSUBS 0.049716f
C1203 VTAIL.n192 VSUBS 0.049716f
C1204 VTAIL.n193 VSUBS 0.022271f
C1205 VTAIL.n194 VSUBS 0.021034f
C1206 VTAIL.n195 VSUBS 0.039143f
C1207 VTAIL.n196 VSUBS 0.039143f
C1208 VTAIL.n197 VSUBS 0.021034f
C1209 VTAIL.n198 VSUBS 0.022271f
C1210 VTAIL.n199 VSUBS 0.049716f
C1211 VTAIL.n200 VSUBS 0.049716f
C1212 VTAIL.n201 VSUBS 0.022271f
C1213 VTAIL.n202 VSUBS 0.021034f
C1214 VTAIL.n203 VSUBS 0.039143f
C1215 VTAIL.n204 VSUBS 0.039143f
C1216 VTAIL.n205 VSUBS 0.021034f
C1217 VTAIL.n206 VSUBS 0.022271f
C1218 VTAIL.n207 VSUBS 0.049716f
C1219 VTAIL.n208 VSUBS 0.049716f
C1220 VTAIL.n209 VSUBS 0.022271f
C1221 VTAIL.n210 VSUBS 0.021034f
C1222 VTAIL.n211 VSUBS 0.039143f
C1223 VTAIL.n212 VSUBS 0.039143f
C1224 VTAIL.n213 VSUBS 0.021034f
C1225 VTAIL.n214 VSUBS 0.022271f
C1226 VTAIL.n215 VSUBS 0.049716f
C1227 VTAIL.n216 VSUBS 0.126017f
C1228 VTAIL.n217 VSUBS 0.022271f
C1229 VTAIL.n218 VSUBS 0.041305f
C1230 VTAIL.n219 VSUBS 0.102241f
C1231 VTAIL.n220 VSUBS 0.097877f
C1232 VTAIL.n221 VSUBS 0.180895f
C1233 VTAIL.t3 VSUBS 0.604407f
C1234 VTAIL.t4 VSUBS 0.604407f
C1235 VTAIL.n222 VSUBS 4.89019f
C1236 VTAIL.n223 VSUBS 1.04803f
C1237 VTAIL.t18 VSUBS 0.604407f
C1238 VTAIL.t5 VSUBS 0.604407f
C1239 VTAIL.n224 VSUBS 4.89019f
C1240 VTAIL.n225 VSUBS 1.01596f
C1241 VTAIL.n226 VSUBS 0.04355f
C1242 VTAIL.n227 VSUBS 0.039143f
C1243 VTAIL.n228 VSUBS 0.021034f
C1244 VTAIL.n229 VSUBS 0.049716f
C1245 VTAIL.n230 VSUBS 0.022271f
C1246 VTAIL.n231 VSUBS 0.039143f
C1247 VTAIL.n232 VSUBS 0.021034f
C1248 VTAIL.n233 VSUBS 0.049716f
C1249 VTAIL.n234 VSUBS 0.022271f
C1250 VTAIL.n235 VSUBS 0.039143f
C1251 VTAIL.n236 VSUBS 0.021034f
C1252 VTAIL.n237 VSUBS 0.049716f
C1253 VTAIL.n238 VSUBS 0.022271f
C1254 VTAIL.n239 VSUBS 0.039143f
C1255 VTAIL.n240 VSUBS 0.021034f
C1256 VTAIL.n241 VSUBS 0.049716f
C1257 VTAIL.n242 VSUBS 0.022271f
C1258 VTAIL.n243 VSUBS 0.039143f
C1259 VTAIL.n244 VSUBS 0.021034f
C1260 VTAIL.n245 VSUBS 0.049716f
C1261 VTAIL.n246 VSUBS 0.022271f
C1262 VTAIL.n247 VSUBS 0.039143f
C1263 VTAIL.n248 VSUBS 0.021034f
C1264 VTAIL.n249 VSUBS 0.049716f
C1265 VTAIL.n250 VSUBS 0.022271f
C1266 VTAIL.n251 VSUBS 0.039143f
C1267 VTAIL.n252 VSUBS 0.021034f
C1268 VTAIL.n253 VSUBS 0.049716f
C1269 VTAIL.n254 VSUBS 0.049716f
C1270 VTAIL.n255 VSUBS 0.022271f
C1271 VTAIL.n256 VSUBS 0.039143f
C1272 VTAIL.n257 VSUBS 0.021034f
C1273 VTAIL.n258 VSUBS 0.049716f
C1274 VTAIL.n259 VSUBS 0.022271f
C1275 VTAIL.n260 VSUBS 0.44172f
C1276 VTAIL.t0 VSUBS 0.10813f
C1277 VTAIL.n261 VSUBS 0.037287f
C1278 VTAIL.n262 VSUBS 0.037399f
C1279 VTAIL.n263 VSUBS 0.021034f
C1280 VTAIL.n264 VSUBS 3.21639f
C1281 VTAIL.n265 VSUBS 0.039143f
C1282 VTAIL.n266 VSUBS 0.021034f
C1283 VTAIL.n267 VSUBS 0.022271f
C1284 VTAIL.n268 VSUBS 0.049716f
C1285 VTAIL.n269 VSUBS 0.049716f
C1286 VTAIL.n270 VSUBS 0.022271f
C1287 VTAIL.n271 VSUBS 0.021034f
C1288 VTAIL.n272 VSUBS 0.039143f
C1289 VTAIL.n273 VSUBS 0.039143f
C1290 VTAIL.n274 VSUBS 0.021034f
C1291 VTAIL.n275 VSUBS 0.022271f
C1292 VTAIL.n276 VSUBS 0.049716f
C1293 VTAIL.n277 VSUBS 0.049716f
C1294 VTAIL.n278 VSUBS 0.022271f
C1295 VTAIL.n279 VSUBS 0.021034f
C1296 VTAIL.n280 VSUBS 0.039143f
C1297 VTAIL.n281 VSUBS 0.039143f
C1298 VTAIL.n282 VSUBS 0.021034f
C1299 VTAIL.n283 VSUBS 0.021652f
C1300 VTAIL.n284 VSUBS 0.021652f
C1301 VTAIL.n285 VSUBS 0.049716f
C1302 VTAIL.n286 VSUBS 0.049716f
C1303 VTAIL.n287 VSUBS 0.022271f
C1304 VTAIL.n288 VSUBS 0.021034f
C1305 VTAIL.n289 VSUBS 0.039143f
C1306 VTAIL.n290 VSUBS 0.039143f
C1307 VTAIL.n291 VSUBS 0.021034f
C1308 VTAIL.n292 VSUBS 0.022271f
C1309 VTAIL.n293 VSUBS 0.049716f
C1310 VTAIL.n294 VSUBS 0.049716f
C1311 VTAIL.n295 VSUBS 0.022271f
C1312 VTAIL.n296 VSUBS 0.021034f
C1313 VTAIL.n297 VSUBS 0.039143f
C1314 VTAIL.n298 VSUBS 0.039143f
C1315 VTAIL.n299 VSUBS 0.021034f
C1316 VTAIL.n300 VSUBS 0.022271f
C1317 VTAIL.n301 VSUBS 0.049716f
C1318 VTAIL.n302 VSUBS 0.049716f
C1319 VTAIL.n303 VSUBS 0.022271f
C1320 VTAIL.n304 VSUBS 0.021034f
C1321 VTAIL.n305 VSUBS 0.039143f
C1322 VTAIL.n306 VSUBS 0.039143f
C1323 VTAIL.n307 VSUBS 0.021034f
C1324 VTAIL.n308 VSUBS 0.022271f
C1325 VTAIL.n309 VSUBS 0.049716f
C1326 VTAIL.n310 VSUBS 0.049716f
C1327 VTAIL.n311 VSUBS 0.022271f
C1328 VTAIL.n312 VSUBS 0.021034f
C1329 VTAIL.n313 VSUBS 0.039143f
C1330 VTAIL.n314 VSUBS 0.039143f
C1331 VTAIL.n315 VSUBS 0.021034f
C1332 VTAIL.n316 VSUBS 0.022271f
C1333 VTAIL.n317 VSUBS 0.049716f
C1334 VTAIL.n318 VSUBS 0.049716f
C1335 VTAIL.n319 VSUBS 0.022271f
C1336 VTAIL.n320 VSUBS 0.021034f
C1337 VTAIL.n321 VSUBS 0.039143f
C1338 VTAIL.n322 VSUBS 0.039143f
C1339 VTAIL.n323 VSUBS 0.021034f
C1340 VTAIL.n324 VSUBS 0.022271f
C1341 VTAIL.n325 VSUBS 0.049716f
C1342 VTAIL.n326 VSUBS 0.126017f
C1343 VTAIL.n327 VSUBS 0.022271f
C1344 VTAIL.n328 VSUBS 0.041305f
C1345 VTAIL.n329 VSUBS 0.102241f
C1346 VTAIL.n330 VSUBS 0.097877f
C1347 VTAIL.n331 VSUBS 2.80511f
C1348 VTAIL.n332 VSUBS 0.04355f
C1349 VTAIL.n333 VSUBS 0.039143f
C1350 VTAIL.n334 VSUBS 0.021034f
C1351 VTAIL.n335 VSUBS 0.049716f
C1352 VTAIL.n336 VSUBS 0.022271f
C1353 VTAIL.n337 VSUBS 0.039143f
C1354 VTAIL.n338 VSUBS 0.021034f
C1355 VTAIL.n339 VSUBS 0.049716f
C1356 VTAIL.n340 VSUBS 0.022271f
C1357 VTAIL.n341 VSUBS 0.039143f
C1358 VTAIL.n342 VSUBS 0.021034f
C1359 VTAIL.n343 VSUBS 0.049716f
C1360 VTAIL.n344 VSUBS 0.022271f
C1361 VTAIL.n345 VSUBS 0.039143f
C1362 VTAIL.n346 VSUBS 0.021034f
C1363 VTAIL.n347 VSUBS 0.049716f
C1364 VTAIL.n348 VSUBS 0.022271f
C1365 VTAIL.n349 VSUBS 0.039143f
C1366 VTAIL.n350 VSUBS 0.021034f
C1367 VTAIL.n351 VSUBS 0.049716f
C1368 VTAIL.n352 VSUBS 0.022271f
C1369 VTAIL.n353 VSUBS 0.039143f
C1370 VTAIL.n354 VSUBS 0.021034f
C1371 VTAIL.n355 VSUBS 0.049716f
C1372 VTAIL.n356 VSUBS 0.022271f
C1373 VTAIL.n357 VSUBS 0.039143f
C1374 VTAIL.n358 VSUBS 0.021034f
C1375 VTAIL.n359 VSUBS 0.049716f
C1376 VTAIL.n360 VSUBS 0.022271f
C1377 VTAIL.n361 VSUBS 0.039143f
C1378 VTAIL.n362 VSUBS 0.021034f
C1379 VTAIL.n363 VSUBS 0.049716f
C1380 VTAIL.n364 VSUBS 0.022271f
C1381 VTAIL.n365 VSUBS 0.44172f
C1382 VTAIL.t7 VSUBS 0.10813f
C1383 VTAIL.n366 VSUBS 0.037287f
C1384 VTAIL.n367 VSUBS 0.037399f
C1385 VTAIL.n368 VSUBS 0.021034f
C1386 VTAIL.n369 VSUBS 3.21638f
C1387 VTAIL.n370 VSUBS 0.039143f
C1388 VTAIL.n371 VSUBS 0.021034f
C1389 VTAIL.n372 VSUBS 0.022271f
C1390 VTAIL.n373 VSUBS 0.049716f
C1391 VTAIL.n374 VSUBS 0.049716f
C1392 VTAIL.n375 VSUBS 0.022271f
C1393 VTAIL.n376 VSUBS 0.021034f
C1394 VTAIL.n377 VSUBS 0.039143f
C1395 VTAIL.n378 VSUBS 0.039143f
C1396 VTAIL.n379 VSUBS 0.021034f
C1397 VTAIL.n380 VSUBS 0.022271f
C1398 VTAIL.n381 VSUBS 0.049716f
C1399 VTAIL.n382 VSUBS 0.049716f
C1400 VTAIL.n383 VSUBS 0.049716f
C1401 VTAIL.n384 VSUBS 0.022271f
C1402 VTAIL.n385 VSUBS 0.021034f
C1403 VTAIL.n386 VSUBS 0.039143f
C1404 VTAIL.n387 VSUBS 0.039143f
C1405 VTAIL.n388 VSUBS 0.021034f
C1406 VTAIL.n389 VSUBS 0.021652f
C1407 VTAIL.n390 VSUBS 0.021652f
C1408 VTAIL.n391 VSUBS 0.049716f
C1409 VTAIL.n392 VSUBS 0.049716f
C1410 VTAIL.n393 VSUBS 0.022271f
C1411 VTAIL.n394 VSUBS 0.021034f
C1412 VTAIL.n395 VSUBS 0.039143f
C1413 VTAIL.n396 VSUBS 0.039143f
C1414 VTAIL.n397 VSUBS 0.021034f
C1415 VTAIL.n398 VSUBS 0.022271f
C1416 VTAIL.n399 VSUBS 0.049716f
C1417 VTAIL.n400 VSUBS 0.049716f
C1418 VTAIL.n401 VSUBS 0.022271f
C1419 VTAIL.n402 VSUBS 0.021034f
C1420 VTAIL.n403 VSUBS 0.039143f
C1421 VTAIL.n404 VSUBS 0.039143f
C1422 VTAIL.n405 VSUBS 0.021034f
C1423 VTAIL.n406 VSUBS 0.022271f
C1424 VTAIL.n407 VSUBS 0.049716f
C1425 VTAIL.n408 VSUBS 0.049716f
C1426 VTAIL.n409 VSUBS 0.022271f
C1427 VTAIL.n410 VSUBS 0.021034f
C1428 VTAIL.n411 VSUBS 0.039143f
C1429 VTAIL.n412 VSUBS 0.039143f
C1430 VTAIL.n413 VSUBS 0.021034f
C1431 VTAIL.n414 VSUBS 0.022271f
C1432 VTAIL.n415 VSUBS 0.049716f
C1433 VTAIL.n416 VSUBS 0.049716f
C1434 VTAIL.n417 VSUBS 0.022271f
C1435 VTAIL.n418 VSUBS 0.021034f
C1436 VTAIL.n419 VSUBS 0.039143f
C1437 VTAIL.n420 VSUBS 0.039143f
C1438 VTAIL.n421 VSUBS 0.021034f
C1439 VTAIL.n422 VSUBS 0.022271f
C1440 VTAIL.n423 VSUBS 0.049716f
C1441 VTAIL.n424 VSUBS 0.049716f
C1442 VTAIL.n425 VSUBS 0.022271f
C1443 VTAIL.n426 VSUBS 0.021034f
C1444 VTAIL.n427 VSUBS 0.039143f
C1445 VTAIL.n428 VSUBS 0.039143f
C1446 VTAIL.n429 VSUBS 0.021034f
C1447 VTAIL.n430 VSUBS 0.022271f
C1448 VTAIL.n431 VSUBS 0.049716f
C1449 VTAIL.n432 VSUBS 0.126017f
C1450 VTAIL.n433 VSUBS 0.022271f
C1451 VTAIL.n434 VSUBS 0.041305f
C1452 VTAIL.n435 VSUBS 0.102241f
C1453 VTAIL.n436 VSUBS 0.097877f
C1454 VTAIL.n437 VSUBS 2.80511f
C1455 VTAIL.t15 VSUBS 0.604407f
C1456 VTAIL.t16 VSUBS 0.604407f
C1457 VTAIL.n438 VSUBS 4.89016f
C1458 VTAIL.n439 VSUBS 0.967874f
C1459 VDD2.n0 VSUBS 0.0435f
C1460 VDD2.n1 VSUBS 0.039097f
C1461 VDD2.n2 VSUBS 0.021009f
C1462 VDD2.n3 VSUBS 0.049658f
C1463 VDD2.n4 VSUBS 0.022245f
C1464 VDD2.n5 VSUBS 0.039097f
C1465 VDD2.n6 VSUBS 0.021009f
C1466 VDD2.n7 VSUBS 0.049658f
C1467 VDD2.n8 VSUBS 0.022245f
C1468 VDD2.n9 VSUBS 0.039097f
C1469 VDD2.n10 VSUBS 0.021009f
C1470 VDD2.n11 VSUBS 0.049658f
C1471 VDD2.n12 VSUBS 0.022245f
C1472 VDD2.n13 VSUBS 0.039097f
C1473 VDD2.n14 VSUBS 0.021009f
C1474 VDD2.n15 VSUBS 0.049658f
C1475 VDD2.n16 VSUBS 0.022245f
C1476 VDD2.n17 VSUBS 0.039097f
C1477 VDD2.n18 VSUBS 0.021009f
C1478 VDD2.n19 VSUBS 0.049658f
C1479 VDD2.n20 VSUBS 0.022245f
C1480 VDD2.n21 VSUBS 0.039097f
C1481 VDD2.n22 VSUBS 0.021009f
C1482 VDD2.n23 VSUBS 0.049658f
C1483 VDD2.n24 VSUBS 0.022245f
C1484 VDD2.n25 VSUBS 0.039097f
C1485 VDD2.n26 VSUBS 0.021009f
C1486 VDD2.n27 VSUBS 0.049658f
C1487 VDD2.n28 VSUBS 0.022245f
C1488 VDD2.n29 VSUBS 0.039097f
C1489 VDD2.n30 VSUBS 0.021009f
C1490 VDD2.n31 VSUBS 0.049658f
C1491 VDD2.n32 VSUBS 0.022245f
C1492 VDD2.n33 VSUBS 0.44121f
C1493 VDD2.t6 VSUBS 0.108005f
C1494 VDD2.n34 VSUBS 0.037244f
C1495 VDD2.n35 VSUBS 0.037356f
C1496 VDD2.n36 VSUBS 0.021009f
C1497 VDD2.n37 VSUBS 3.21267f
C1498 VDD2.n38 VSUBS 0.039097f
C1499 VDD2.n39 VSUBS 0.021009f
C1500 VDD2.n40 VSUBS 0.022245f
C1501 VDD2.n41 VSUBS 0.049658f
C1502 VDD2.n42 VSUBS 0.049658f
C1503 VDD2.n43 VSUBS 0.022245f
C1504 VDD2.n44 VSUBS 0.021009f
C1505 VDD2.n45 VSUBS 0.039097f
C1506 VDD2.n46 VSUBS 0.039097f
C1507 VDD2.n47 VSUBS 0.021009f
C1508 VDD2.n48 VSUBS 0.022245f
C1509 VDD2.n49 VSUBS 0.049658f
C1510 VDD2.n50 VSUBS 0.049658f
C1511 VDD2.n51 VSUBS 0.049658f
C1512 VDD2.n52 VSUBS 0.022245f
C1513 VDD2.n53 VSUBS 0.021009f
C1514 VDD2.n54 VSUBS 0.039097f
C1515 VDD2.n55 VSUBS 0.039097f
C1516 VDD2.n56 VSUBS 0.021009f
C1517 VDD2.n57 VSUBS 0.021627f
C1518 VDD2.n58 VSUBS 0.021627f
C1519 VDD2.n59 VSUBS 0.049658f
C1520 VDD2.n60 VSUBS 0.049658f
C1521 VDD2.n61 VSUBS 0.022245f
C1522 VDD2.n62 VSUBS 0.021009f
C1523 VDD2.n63 VSUBS 0.039097f
C1524 VDD2.n64 VSUBS 0.039097f
C1525 VDD2.n65 VSUBS 0.021009f
C1526 VDD2.n66 VSUBS 0.022245f
C1527 VDD2.n67 VSUBS 0.049658f
C1528 VDD2.n68 VSUBS 0.049658f
C1529 VDD2.n69 VSUBS 0.022245f
C1530 VDD2.n70 VSUBS 0.021009f
C1531 VDD2.n71 VSUBS 0.039097f
C1532 VDD2.n72 VSUBS 0.039097f
C1533 VDD2.n73 VSUBS 0.021009f
C1534 VDD2.n74 VSUBS 0.022245f
C1535 VDD2.n75 VSUBS 0.049658f
C1536 VDD2.n76 VSUBS 0.049658f
C1537 VDD2.n77 VSUBS 0.022245f
C1538 VDD2.n78 VSUBS 0.021009f
C1539 VDD2.n79 VSUBS 0.039097f
C1540 VDD2.n80 VSUBS 0.039097f
C1541 VDD2.n81 VSUBS 0.021009f
C1542 VDD2.n82 VSUBS 0.022245f
C1543 VDD2.n83 VSUBS 0.049658f
C1544 VDD2.n84 VSUBS 0.049658f
C1545 VDD2.n85 VSUBS 0.022245f
C1546 VDD2.n86 VSUBS 0.021009f
C1547 VDD2.n87 VSUBS 0.039097f
C1548 VDD2.n88 VSUBS 0.039097f
C1549 VDD2.n89 VSUBS 0.021009f
C1550 VDD2.n90 VSUBS 0.022245f
C1551 VDD2.n91 VSUBS 0.049658f
C1552 VDD2.n92 VSUBS 0.049658f
C1553 VDD2.n93 VSUBS 0.022245f
C1554 VDD2.n94 VSUBS 0.021009f
C1555 VDD2.n95 VSUBS 0.039097f
C1556 VDD2.n96 VSUBS 0.039097f
C1557 VDD2.n97 VSUBS 0.021009f
C1558 VDD2.n98 VSUBS 0.022245f
C1559 VDD2.n99 VSUBS 0.049658f
C1560 VDD2.n100 VSUBS 0.125871f
C1561 VDD2.n101 VSUBS 0.022245f
C1562 VDD2.n102 VSUBS 0.041257f
C1563 VDD2.n103 VSUBS 0.102122f
C1564 VDD2.n104 VSUBS 0.125776f
C1565 VDD2.t2 VSUBS 0.603708f
C1566 VDD2.t4 VSUBS 0.603708f
C1567 VDD2.n105 VSUBS 5.10469f
C1568 VDD2.n106 VSUBS 0.952596f
C1569 VDD2.t0 VSUBS 0.603708f
C1570 VDD2.t7 VSUBS 0.603708f
C1571 VDD2.n107 VSUBS 5.10782f
C1572 VDD2.n108 VSUBS 3.66911f
C1573 VDD2.n109 VSUBS 0.0435f
C1574 VDD2.n110 VSUBS 0.039097f
C1575 VDD2.n111 VSUBS 0.021009f
C1576 VDD2.n112 VSUBS 0.049658f
C1577 VDD2.n113 VSUBS 0.022245f
C1578 VDD2.n114 VSUBS 0.039097f
C1579 VDD2.n115 VSUBS 0.021009f
C1580 VDD2.n116 VSUBS 0.049658f
C1581 VDD2.n117 VSUBS 0.022245f
C1582 VDD2.n118 VSUBS 0.039097f
C1583 VDD2.n119 VSUBS 0.021009f
C1584 VDD2.n120 VSUBS 0.049658f
C1585 VDD2.n121 VSUBS 0.022245f
C1586 VDD2.n122 VSUBS 0.039097f
C1587 VDD2.n123 VSUBS 0.021009f
C1588 VDD2.n124 VSUBS 0.049658f
C1589 VDD2.n125 VSUBS 0.022245f
C1590 VDD2.n126 VSUBS 0.039097f
C1591 VDD2.n127 VSUBS 0.021009f
C1592 VDD2.n128 VSUBS 0.049658f
C1593 VDD2.n129 VSUBS 0.022245f
C1594 VDD2.n130 VSUBS 0.039097f
C1595 VDD2.n131 VSUBS 0.021009f
C1596 VDD2.n132 VSUBS 0.049658f
C1597 VDD2.n133 VSUBS 0.022245f
C1598 VDD2.n134 VSUBS 0.039097f
C1599 VDD2.n135 VSUBS 0.021009f
C1600 VDD2.n136 VSUBS 0.049658f
C1601 VDD2.n137 VSUBS 0.049658f
C1602 VDD2.n138 VSUBS 0.022245f
C1603 VDD2.n139 VSUBS 0.039097f
C1604 VDD2.n140 VSUBS 0.021009f
C1605 VDD2.n141 VSUBS 0.049658f
C1606 VDD2.n142 VSUBS 0.022245f
C1607 VDD2.n143 VSUBS 0.44121f
C1608 VDD2.t1 VSUBS 0.108005f
C1609 VDD2.n144 VSUBS 0.037244f
C1610 VDD2.n145 VSUBS 0.037356f
C1611 VDD2.n146 VSUBS 0.021009f
C1612 VDD2.n147 VSUBS 3.21267f
C1613 VDD2.n148 VSUBS 0.039097f
C1614 VDD2.n149 VSUBS 0.021009f
C1615 VDD2.n150 VSUBS 0.022245f
C1616 VDD2.n151 VSUBS 0.049658f
C1617 VDD2.n152 VSUBS 0.049658f
C1618 VDD2.n153 VSUBS 0.022245f
C1619 VDD2.n154 VSUBS 0.021009f
C1620 VDD2.n155 VSUBS 0.039097f
C1621 VDD2.n156 VSUBS 0.039097f
C1622 VDD2.n157 VSUBS 0.021009f
C1623 VDD2.n158 VSUBS 0.022245f
C1624 VDD2.n159 VSUBS 0.049658f
C1625 VDD2.n160 VSUBS 0.049658f
C1626 VDD2.n161 VSUBS 0.022245f
C1627 VDD2.n162 VSUBS 0.021009f
C1628 VDD2.n163 VSUBS 0.039097f
C1629 VDD2.n164 VSUBS 0.039097f
C1630 VDD2.n165 VSUBS 0.021009f
C1631 VDD2.n166 VSUBS 0.021627f
C1632 VDD2.n167 VSUBS 0.021627f
C1633 VDD2.n168 VSUBS 0.049658f
C1634 VDD2.n169 VSUBS 0.049658f
C1635 VDD2.n170 VSUBS 0.022245f
C1636 VDD2.n171 VSUBS 0.021009f
C1637 VDD2.n172 VSUBS 0.039097f
C1638 VDD2.n173 VSUBS 0.039097f
C1639 VDD2.n174 VSUBS 0.021009f
C1640 VDD2.n175 VSUBS 0.022245f
C1641 VDD2.n176 VSUBS 0.049658f
C1642 VDD2.n177 VSUBS 0.049658f
C1643 VDD2.n178 VSUBS 0.022245f
C1644 VDD2.n179 VSUBS 0.021009f
C1645 VDD2.n180 VSUBS 0.039097f
C1646 VDD2.n181 VSUBS 0.039097f
C1647 VDD2.n182 VSUBS 0.021009f
C1648 VDD2.n183 VSUBS 0.022245f
C1649 VDD2.n184 VSUBS 0.049658f
C1650 VDD2.n185 VSUBS 0.049658f
C1651 VDD2.n186 VSUBS 0.022245f
C1652 VDD2.n187 VSUBS 0.021009f
C1653 VDD2.n188 VSUBS 0.039097f
C1654 VDD2.n189 VSUBS 0.039097f
C1655 VDD2.n190 VSUBS 0.021009f
C1656 VDD2.n191 VSUBS 0.022245f
C1657 VDD2.n192 VSUBS 0.049658f
C1658 VDD2.n193 VSUBS 0.049658f
C1659 VDD2.n194 VSUBS 0.022245f
C1660 VDD2.n195 VSUBS 0.021009f
C1661 VDD2.n196 VSUBS 0.039097f
C1662 VDD2.n197 VSUBS 0.039097f
C1663 VDD2.n198 VSUBS 0.021009f
C1664 VDD2.n199 VSUBS 0.022245f
C1665 VDD2.n200 VSUBS 0.049658f
C1666 VDD2.n201 VSUBS 0.049658f
C1667 VDD2.n202 VSUBS 0.022245f
C1668 VDD2.n203 VSUBS 0.021009f
C1669 VDD2.n204 VSUBS 0.039097f
C1670 VDD2.n205 VSUBS 0.039097f
C1671 VDD2.n206 VSUBS 0.021009f
C1672 VDD2.n207 VSUBS 0.022245f
C1673 VDD2.n208 VSUBS 0.049658f
C1674 VDD2.n209 VSUBS 0.125871f
C1675 VDD2.n210 VSUBS 0.022245f
C1676 VDD2.n211 VSUBS 0.041257f
C1677 VDD2.n212 VSUBS 0.102122f
C1678 VDD2.n213 VSUBS 0.124679f
C1679 VDD2.n214 VSUBS 3.9662f
C1680 VDD2.t9 VSUBS 0.603708f
C1681 VDD2.t8 VSUBS 0.603708f
C1682 VDD2.n215 VSUBS 5.10471f
C1683 VDD2.n216 VSUBS 0.814363f
C1684 VDD2.t3 VSUBS 0.603708f
C1685 VDD2.t5 VSUBS 0.603708f
C1686 VDD2.n217 VSUBS 5.10777f
C1687 VN.n0 VSUBS 0.071051f
C1688 VN.t0 VSUBS 0.664814f
C1689 VN.t1 VSUBS 0.664814f
C1690 VN.t3 VSUBS 0.664814f
C1691 VN.n1 VSUBS 0.257048f
C1692 VN.t5 VSUBS 0.66791f
C1693 VN.n2 VSUBS 0.27411f
C1694 VN.n3 VSUBS 0.149457f
C1695 VN.n4 VSUBS 0.02357f
C1696 VN.n5 VSUBS 0.257048f
C1697 VN.n6 VSUBS 0.02357f
C1698 VN.n7 VSUBS 0.257048f
C1699 VN.t9 VSUBS 0.66791f
C1700 VN.n8 VSUBS 0.274018f
C1701 VN.n9 VSUBS 0.055062f
C1702 VN.n10 VSUBS 0.071051f
C1703 VN.t4 VSUBS 0.66791f
C1704 VN.t7 VSUBS 0.664814f
C1705 VN.t8 VSUBS 0.664814f
C1706 VN.t2 VSUBS 0.664814f
C1707 VN.n11 VSUBS 0.257048f
C1708 VN.t6 VSUBS 0.66791f
C1709 VN.n12 VSUBS 0.27411f
C1710 VN.n13 VSUBS 0.149457f
C1711 VN.n14 VSUBS 0.02357f
C1712 VN.n15 VSUBS 0.257048f
C1713 VN.n16 VSUBS 0.02357f
C1714 VN.n17 VSUBS 0.257048f
C1715 VN.n18 VSUBS 0.274018f
C1716 VN.n19 VSUBS 3.40123f
.ends

