* NGSPICE file created from diff_pair_sample_0465.ext - technology: sky130A

.subckt diff_pair_sample_0465 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.39
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.39
X2 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.39
X3 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.39
X4 VTAIL.t6 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.39
X5 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.39
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.39
X7 VDD1.t1 VP.t2 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.39
X8 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.39
X9 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.39
X10 VTAIL.t7 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.39
X11 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.39
R0 B.n323 B.n322 585
R1 B.n324 B.n323 585
R2 B.n108 B.n58 585
R3 B.n107 B.n106 585
R4 B.n105 B.n104 585
R5 B.n103 B.n102 585
R6 B.n101 B.n100 585
R7 B.n99 B.n98 585
R8 B.n97 B.n96 585
R9 B.n94 B.n93 585
R10 B.n92 B.n91 585
R11 B.n90 B.n89 585
R12 B.n88 B.n87 585
R13 B.n86 B.n85 585
R14 B.n84 B.n83 585
R15 B.n82 B.n81 585
R16 B.n80 B.n79 585
R17 B.n78 B.n77 585
R18 B.n76 B.n75 585
R19 B.n74 B.n73 585
R20 B.n72 B.n71 585
R21 B.n70 B.n69 585
R22 B.n68 B.n67 585
R23 B.n66 B.n65 585
R24 B.n46 B.n45 585
R25 B.n327 B.n326 585
R26 B.n321 B.n59 585
R27 B.n59 B.n43 585
R28 B.n320 B.n42 585
R29 B.n331 B.n42 585
R30 B.n319 B.n41 585
R31 B.n332 B.n41 585
R32 B.n318 B.n40 585
R33 B.n333 B.n40 585
R34 B.n317 B.n316 585
R35 B.n316 B.n36 585
R36 B.n315 B.n35 585
R37 B.n339 B.n35 585
R38 B.n314 B.n34 585
R39 B.n340 B.n34 585
R40 B.n313 B.n33 585
R41 B.n341 B.n33 585
R42 B.n312 B.n311 585
R43 B.n311 B.n29 585
R44 B.n310 B.n28 585
R45 B.n347 B.n28 585
R46 B.n309 B.n27 585
R47 B.n348 B.n27 585
R48 B.n308 B.n26 585
R49 B.n349 B.n26 585
R50 B.n307 B.n306 585
R51 B.n306 B.n22 585
R52 B.n305 B.n21 585
R53 B.n355 B.n21 585
R54 B.n304 B.n20 585
R55 B.n356 B.n20 585
R56 B.n303 B.n19 585
R57 B.n357 B.n19 585
R58 B.n302 B.n301 585
R59 B.n301 B.n15 585
R60 B.n300 B.n14 585
R61 B.n363 B.n14 585
R62 B.n299 B.n13 585
R63 B.n364 B.n13 585
R64 B.n298 B.n12 585
R65 B.n365 B.n12 585
R66 B.n297 B.n296 585
R67 B.n296 B.n295 585
R68 B.n294 B.n293 585
R69 B.n294 B.n8 585
R70 B.n292 B.n7 585
R71 B.n372 B.n7 585
R72 B.n291 B.n6 585
R73 B.n373 B.n6 585
R74 B.n290 B.n5 585
R75 B.n374 B.n5 585
R76 B.n289 B.n288 585
R77 B.n288 B.n4 585
R78 B.n287 B.n109 585
R79 B.n287 B.n286 585
R80 B.n277 B.n110 585
R81 B.n111 B.n110 585
R82 B.n279 B.n278 585
R83 B.n280 B.n279 585
R84 B.n276 B.n116 585
R85 B.n116 B.n115 585
R86 B.n275 B.n274 585
R87 B.n274 B.n273 585
R88 B.n118 B.n117 585
R89 B.n119 B.n118 585
R90 B.n266 B.n265 585
R91 B.n267 B.n266 585
R92 B.n264 B.n123 585
R93 B.n127 B.n123 585
R94 B.n263 B.n262 585
R95 B.n262 B.n261 585
R96 B.n125 B.n124 585
R97 B.n126 B.n125 585
R98 B.n254 B.n253 585
R99 B.n255 B.n254 585
R100 B.n252 B.n132 585
R101 B.n132 B.n131 585
R102 B.n251 B.n250 585
R103 B.n250 B.n249 585
R104 B.n134 B.n133 585
R105 B.n135 B.n134 585
R106 B.n242 B.n241 585
R107 B.n243 B.n242 585
R108 B.n240 B.n139 585
R109 B.n143 B.n139 585
R110 B.n239 B.n238 585
R111 B.n238 B.n237 585
R112 B.n141 B.n140 585
R113 B.n142 B.n141 585
R114 B.n230 B.n229 585
R115 B.n231 B.n230 585
R116 B.n228 B.n148 585
R117 B.n148 B.n147 585
R118 B.n227 B.n226 585
R119 B.n226 B.n225 585
R120 B.n150 B.n149 585
R121 B.n151 B.n150 585
R122 B.n221 B.n220 585
R123 B.n154 B.n153 585
R124 B.n217 B.n216 585
R125 B.n218 B.n217 585
R126 B.n215 B.n166 585
R127 B.n214 B.n213 585
R128 B.n212 B.n211 585
R129 B.n210 B.n209 585
R130 B.n208 B.n207 585
R131 B.n205 B.n204 585
R132 B.n203 B.n202 585
R133 B.n201 B.n200 585
R134 B.n199 B.n198 585
R135 B.n197 B.n196 585
R136 B.n195 B.n194 585
R137 B.n193 B.n192 585
R138 B.n191 B.n190 585
R139 B.n189 B.n188 585
R140 B.n187 B.n186 585
R141 B.n185 B.n184 585
R142 B.n183 B.n182 585
R143 B.n181 B.n180 585
R144 B.n179 B.n178 585
R145 B.n177 B.n176 585
R146 B.n175 B.n174 585
R147 B.n173 B.n172 585
R148 B.n222 B.n152 585
R149 B.n152 B.n151 585
R150 B.n224 B.n223 585
R151 B.n225 B.n224 585
R152 B.n146 B.n145 585
R153 B.n147 B.n146 585
R154 B.n233 B.n232 585
R155 B.n232 B.n231 585
R156 B.n234 B.n144 585
R157 B.n144 B.n142 585
R158 B.n236 B.n235 585
R159 B.n237 B.n236 585
R160 B.n138 B.n137 585
R161 B.n143 B.n138 585
R162 B.n245 B.n244 585
R163 B.n244 B.n243 585
R164 B.n246 B.n136 585
R165 B.n136 B.n135 585
R166 B.n248 B.n247 585
R167 B.n249 B.n248 585
R168 B.n130 B.n129 585
R169 B.n131 B.n130 585
R170 B.n257 B.n256 585
R171 B.n256 B.n255 585
R172 B.n258 B.n128 585
R173 B.n128 B.n126 585
R174 B.n260 B.n259 585
R175 B.n261 B.n260 585
R176 B.n122 B.n121 585
R177 B.n127 B.n122 585
R178 B.n269 B.n268 585
R179 B.n268 B.n267 585
R180 B.n270 B.n120 585
R181 B.n120 B.n119 585
R182 B.n272 B.n271 585
R183 B.n273 B.n272 585
R184 B.n114 B.n113 585
R185 B.n115 B.n114 585
R186 B.n282 B.n281 585
R187 B.n281 B.n280 585
R188 B.n283 B.n112 585
R189 B.n112 B.n111 585
R190 B.n285 B.n284 585
R191 B.n286 B.n285 585
R192 B.n3 B.n0 585
R193 B.n4 B.n3 585
R194 B.n371 B.n1 585
R195 B.n372 B.n371 585
R196 B.n370 B.n369 585
R197 B.n370 B.n8 585
R198 B.n368 B.n9 585
R199 B.n295 B.n9 585
R200 B.n367 B.n366 585
R201 B.n366 B.n365 585
R202 B.n11 B.n10 585
R203 B.n364 B.n11 585
R204 B.n362 B.n361 585
R205 B.n363 B.n362 585
R206 B.n360 B.n16 585
R207 B.n16 B.n15 585
R208 B.n359 B.n358 585
R209 B.n358 B.n357 585
R210 B.n18 B.n17 585
R211 B.n356 B.n18 585
R212 B.n354 B.n353 585
R213 B.n355 B.n354 585
R214 B.n352 B.n23 585
R215 B.n23 B.n22 585
R216 B.n351 B.n350 585
R217 B.n350 B.n349 585
R218 B.n25 B.n24 585
R219 B.n348 B.n25 585
R220 B.n346 B.n345 585
R221 B.n347 B.n346 585
R222 B.n344 B.n30 585
R223 B.n30 B.n29 585
R224 B.n343 B.n342 585
R225 B.n342 B.n341 585
R226 B.n32 B.n31 585
R227 B.n340 B.n32 585
R228 B.n338 B.n337 585
R229 B.n339 B.n338 585
R230 B.n336 B.n37 585
R231 B.n37 B.n36 585
R232 B.n335 B.n334 585
R233 B.n334 B.n333 585
R234 B.n39 B.n38 585
R235 B.n332 B.n39 585
R236 B.n330 B.n329 585
R237 B.n331 B.n330 585
R238 B.n328 B.n44 585
R239 B.n44 B.n43 585
R240 B.n375 B.n374 585
R241 B.n373 B.n2 585
R242 B.n326 B.n44 502.111
R243 B.n323 B.n59 502.111
R244 B.n172 B.n150 502.111
R245 B.n220 B.n152 502.111
R246 B.n62 B.t16 274.721
R247 B.n60 B.t10 274.721
R248 B.n169 B.t7 274.721
R249 B.n167 B.t14 274.721
R250 B.n324 B.n57 256.663
R251 B.n324 B.n56 256.663
R252 B.n324 B.n55 256.663
R253 B.n324 B.n54 256.663
R254 B.n324 B.n53 256.663
R255 B.n324 B.n52 256.663
R256 B.n324 B.n51 256.663
R257 B.n324 B.n50 256.663
R258 B.n324 B.n49 256.663
R259 B.n324 B.n48 256.663
R260 B.n324 B.n47 256.663
R261 B.n325 B.n324 256.663
R262 B.n219 B.n218 256.663
R263 B.n218 B.n155 256.663
R264 B.n218 B.n156 256.663
R265 B.n218 B.n157 256.663
R266 B.n218 B.n158 256.663
R267 B.n218 B.n159 256.663
R268 B.n218 B.n160 256.663
R269 B.n218 B.n161 256.663
R270 B.n218 B.n162 256.663
R271 B.n218 B.n163 256.663
R272 B.n218 B.n164 256.663
R273 B.n218 B.n165 256.663
R274 B.n377 B.n376 256.663
R275 B.n63 B.t17 241.364
R276 B.n61 B.t11 241.364
R277 B.n170 B.t6 241.364
R278 B.n168 B.t13 241.364
R279 B.n62 B.t15 207.294
R280 B.n60 B.t8 207.294
R281 B.n169 B.t4 207.294
R282 B.n167 B.t12 207.294
R283 B.n218 B.n151 205.838
R284 B.n324 B.n43 205.838
R285 B.n65 B.n46 163.367
R286 B.n69 B.n68 163.367
R287 B.n73 B.n72 163.367
R288 B.n77 B.n76 163.367
R289 B.n81 B.n80 163.367
R290 B.n85 B.n84 163.367
R291 B.n89 B.n88 163.367
R292 B.n93 B.n92 163.367
R293 B.n98 B.n97 163.367
R294 B.n102 B.n101 163.367
R295 B.n106 B.n105 163.367
R296 B.n323 B.n58 163.367
R297 B.n226 B.n150 163.367
R298 B.n226 B.n148 163.367
R299 B.n230 B.n148 163.367
R300 B.n230 B.n141 163.367
R301 B.n238 B.n141 163.367
R302 B.n238 B.n139 163.367
R303 B.n242 B.n139 163.367
R304 B.n242 B.n134 163.367
R305 B.n250 B.n134 163.367
R306 B.n250 B.n132 163.367
R307 B.n254 B.n132 163.367
R308 B.n254 B.n125 163.367
R309 B.n262 B.n125 163.367
R310 B.n262 B.n123 163.367
R311 B.n266 B.n123 163.367
R312 B.n266 B.n118 163.367
R313 B.n274 B.n118 163.367
R314 B.n274 B.n116 163.367
R315 B.n279 B.n116 163.367
R316 B.n279 B.n110 163.367
R317 B.n287 B.n110 163.367
R318 B.n288 B.n287 163.367
R319 B.n288 B.n5 163.367
R320 B.n6 B.n5 163.367
R321 B.n7 B.n6 163.367
R322 B.n294 B.n7 163.367
R323 B.n296 B.n294 163.367
R324 B.n296 B.n12 163.367
R325 B.n13 B.n12 163.367
R326 B.n14 B.n13 163.367
R327 B.n301 B.n14 163.367
R328 B.n301 B.n19 163.367
R329 B.n20 B.n19 163.367
R330 B.n21 B.n20 163.367
R331 B.n306 B.n21 163.367
R332 B.n306 B.n26 163.367
R333 B.n27 B.n26 163.367
R334 B.n28 B.n27 163.367
R335 B.n311 B.n28 163.367
R336 B.n311 B.n33 163.367
R337 B.n34 B.n33 163.367
R338 B.n35 B.n34 163.367
R339 B.n316 B.n35 163.367
R340 B.n316 B.n40 163.367
R341 B.n41 B.n40 163.367
R342 B.n42 B.n41 163.367
R343 B.n59 B.n42 163.367
R344 B.n217 B.n154 163.367
R345 B.n217 B.n166 163.367
R346 B.n213 B.n212 163.367
R347 B.n209 B.n208 163.367
R348 B.n204 B.n203 163.367
R349 B.n200 B.n199 163.367
R350 B.n196 B.n195 163.367
R351 B.n192 B.n191 163.367
R352 B.n188 B.n187 163.367
R353 B.n184 B.n183 163.367
R354 B.n180 B.n179 163.367
R355 B.n176 B.n175 163.367
R356 B.n224 B.n152 163.367
R357 B.n224 B.n146 163.367
R358 B.n232 B.n146 163.367
R359 B.n232 B.n144 163.367
R360 B.n236 B.n144 163.367
R361 B.n236 B.n138 163.367
R362 B.n244 B.n138 163.367
R363 B.n244 B.n136 163.367
R364 B.n248 B.n136 163.367
R365 B.n248 B.n130 163.367
R366 B.n256 B.n130 163.367
R367 B.n256 B.n128 163.367
R368 B.n260 B.n128 163.367
R369 B.n260 B.n122 163.367
R370 B.n268 B.n122 163.367
R371 B.n268 B.n120 163.367
R372 B.n272 B.n120 163.367
R373 B.n272 B.n114 163.367
R374 B.n281 B.n114 163.367
R375 B.n281 B.n112 163.367
R376 B.n285 B.n112 163.367
R377 B.n285 B.n3 163.367
R378 B.n375 B.n3 163.367
R379 B.n371 B.n2 163.367
R380 B.n371 B.n370 163.367
R381 B.n370 B.n9 163.367
R382 B.n366 B.n9 163.367
R383 B.n366 B.n11 163.367
R384 B.n362 B.n11 163.367
R385 B.n362 B.n16 163.367
R386 B.n358 B.n16 163.367
R387 B.n358 B.n18 163.367
R388 B.n354 B.n18 163.367
R389 B.n354 B.n23 163.367
R390 B.n350 B.n23 163.367
R391 B.n350 B.n25 163.367
R392 B.n346 B.n25 163.367
R393 B.n346 B.n30 163.367
R394 B.n342 B.n30 163.367
R395 B.n342 B.n32 163.367
R396 B.n338 B.n32 163.367
R397 B.n338 B.n37 163.367
R398 B.n334 B.n37 163.367
R399 B.n334 B.n39 163.367
R400 B.n330 B.n39 163.367
R401 B.n330 B.n44 163.367
R402 B.n225 B.n151 128.412
R403 B.n225 B.n147 128.412
R404 B.n231 B.n147 128.412
R405 B.n231 B.n142 128.412
R406 B.n237 B.n142 128.412
R407 B.n237 B.n143 128.412
R408 B.n243 B.n135 128.412
R409 B.n249 B.n135 128.412
R410 B.n249 B.n131 128.412
R411 B.n255 B.n131 128.412
R412 B.n255 B.n126 128.412
R413 B.n261 B.n126 128.412
R414 B.n261 B.n127 128.412
R415 B.n267 B.n119 128.412
R416 B.n273 B.n119 128.412
R417 B.n273 B.n115 128.412
R418 B.n280 B.n115 128.412
R419 B.n286 B.n111 128.412
R420 B.n286 B.n4 128.412
R421 B.n374 B.n4 128.412
R422 B.n374 B.n373 128.412
R423 B.n373 B.n372 128.412
R424 B.n372 B.n8 128.412
R425 B.n295 B.n8 128.412
R426 B.n365 B.n364 128.412
R427 B.n364 B.n363 128.412
R428 B.n363 B.n15 128.412
R429 B.n357 B.n15 128.412
R430 B.n356 B.n355 128.412
R431 B.n355 B.n22 128.412
R432 B.n349 B.n22 128.412
R433 B.n349 B.n348 128.412
R434 B.n348 B.n347 128.412
R435 B.n347 B.n29 128.412
R436 B.n341 B.n29 128.412
R437 B.n340 B.n339 128.412
R438 B.n339 B.n36 128.412
R439 B.n333 B.n36 128.412
R440 B.n333 B.n332 128.412
R441 B.n332 B.n331 128.412
R442 B.n331 B.n43 128.412
R443 B.n243 B.t5 122.748
R444 B.n341 B.t9 122.748
R445 B.n267 B.t0 88.7559
R446 B.n357 B.t1 88.7559
R447 B.t2 B.n111 81.2022
R448 B.n295 B.t3 81.2022
R449 B.n326 B.n325 71.676
R450 B.n65 B.n47 71.676
R451 B.n69 B.n48 71.676
R452 B.n73 B.n49 71.676
R453 B.n77 B.n50 71.676
R454 B.n81 B.n51 71.676
R455 B.n85 B.n52 71.676
R456 B.n89 B.n53 71.676
R457 B.n93 B.n54 71.676
R458 B.n98 B.n55 71.676
R459 B.n102 B.n56 71.676
R460 B.n106 B.n57 71.676
R461 B.n58 B.n57 71.676
R462 B.n105 B.n56 71.676
R463 B.n101 B.n55 71.676
R464 B.n97 B.n54 71.676
R465 B.n92 B.n53 71.676
R466 B.n88 B.n52 71.676
R467 B.n84 B.n51 71.676
R468 B.n80 B.n50 71.676
R469 B.n76 B.n49 71.676
R470 B.n72 B.n48 71.676
R471 B.n68 B.n47 71.676
R472 B.n325 B.n46 71.676
R473 B.n220 B.n219 71.676
R474 B.n166 B.n155 71.676
R475 B.n212 B.n156 71.676
R476 B.n208 B.n157 71.676
R477 B.n203 B.n158 71.676
R478 B.n199 B.n159 71.676
R479 B.n195 B.n160 71.676
R480 B.n191 B.n161 71.676
R481 B.n187 B.n162 71.676
R482 B.n183 B.n163 71.676
R483 B.n179 B.n164 71.676
R484 B.n175 B.n165 71.676
R485 B.n219 B.n154 71.676
R486 B.n213 B.n155 71.676
R487 B.n209 B.n156 71.676
R488 B.n204 B.n157 71.676
R489 B.n200 B.n158 71.676
R490 B.n196 B.n159 71.676
R491 B.n192 B.n160 71.676
R492 B.n188 B.n161 71.676
R493 B.n184 B.n162 71.676
R494 B.n180 B.n163 71.676
R495 B.n176 B.n164 71.676
R496 B.n172 B.n165 71.676
R497 B.n376 B.n375 71.676
R498 B.n376 B.n2 71.676
R499 B.n64 B.n63 59.5399
R500 B.n95 B.n61 59.5399
R501 B.n171 B.n170 59.5399
R502 B.n206 B.n168 59.5399
R503 B.n280 B.t2 47.2108
R504 B.n365 B.t3 47.2108
R505 B.n127 B.t0 39.6572
R506 B.t1 B.n356 39.6572
R507 B.n63 B.n62 33.3581
R508 B.n61 B.n60 33.3581
R509 B.n170 B.n169 33.3581
R510 B.n168 B.n167 33.3581
R511 B.n222 B.n221 32.6249
R512 B.n173 B.n149 32.6249
R513 B.n322 B.n321 32.6249
R514 B.n328 B.n327 32.6249
R515 B B.n377 18.0485
R516 B.n223 B.n222 10.6151
R517 B.n223 B.n145 10.6151
R518 B.n233 B.n145 10.6151
R519 B.n234 B.n233 10.6151
R520 B.n235 B.n234 10.6151
R521 B.n235 B.n137 10.6151
R522 B.n245 B.n137 10.6151
R523 B.n246 B.n245 10.6151
R524 B.n247 B.n246 10.6151
R525 B.n247 B.n129 10.6151
R526 B.n257 B.n129 10.6151
R527 B.n258 B.n257 10.6151
R528 B.n259 B.n258 10.6151
R529 B.n259 B.n121 10.6151
R530 B.n269 B.n121 10.6151
R531 B.n270 B.n269 10.6151
R532 B.n271 B.n270 10.6151
R533 B.n271 B.n113 10.6151
R534 B.n282 B.n113 10.6151
R535 B.n283 B.n282 10.6151
R536 B.n284 B.n283 10.6151
R537 B.n284 B.n0 10.6151
R538 B.n221 B.n153 10.6151
R539 B.n216 B.n153 10.6151
R540 B.n216 B.n215 10.6151
R541 B.n215 B.n214 10.6151
R542 B.n214 B.n211 10.6151
R543 B.n211 B.n210 10.6151
R544 B.n210 B.n207 10.6151
R545 B.n205 B.n202 10.6151
R546 B.n202 B.n201 10.6151
R547 B.n201 B.n198 10.6151
R548 B.n198 B.n197 10.6151
R549 B.n197 B.n194 10.6151
R550 B.n194 B.n193 10.6151
R551 B.n193 B.n190 10.6151
R552 B.n190 B.n189 10.6151
R553 B.n186 B.n185 10.6151
R554 B.n185 B.n182 10.6151
R555 B.n182 B.n181 10.6151
R556 B.n181 B.n178 10.6151
R557 B.n178 B.n177 10.6151
R558 B.n177 B.n174 10.6151
R559 B.n174 B.n173 10.6151
R560 B.n227 B.n149 10.6151
R561 B.n228 B.n227 10.6151
R562 B.n229 B.n228 10.6151
R563 B.n229 B.n140 10.6151
R564 B.n239 B.n140 10.6151
R565 B.n240 B.n239 10.6151
R566 B.n241 B.n240 10.6151
R567 B.n241 B.n133 10.6151
R568 B.n251 B.n133 10.6151
R569 B.n252 B.n251 10.6151
R570 B.n253 B.n252 10.6151
R571 B.n253 B.n124 10.6151
R572 B.n263 B.n124 10.6151
R573 B.n264 B.n263 10.6151
R574 B.n265 B.n264 10.6151
R575 B.n265 B.n117 10.6151
R576 B.n275 B.n117 10.6151
R577 B.n276 B.n275 10.6151
R578 B.n278 B.n276 10.6151
R579 B.n278 B.n277 10.6151
R580 B.n277 B.n109 10.6151
R581 B.n289 B.n109 10.6151
R582 B.n290 B.n289 10.6151
R583 B.n291 B.n290 10.6151
R584 B.n292 B.n291 10.6151
R585 B.n293 B.n292 10.6151
R586 B.n297 B.n293 10.6151
R587 B.n298 B.n297 10.6151
R588 B.n299 B.n298 10.6151
R589 B.n300 B.n299 10.6151
R590 B.n302 B.n300 10.6151
R591 B.n303 B.n302 10.6151
R592 B.n304 B.n303 10.6151
R593 B.n305 B.n304 10.6151
R594 B.n307 B.n305 10.6151
R595 B.n308 B.n307 10.6151
R596 B.n309 B.n308 10.6151
R597 B.n310 B.n309 10.6151
R598 B.n312 B.n310 10.6151
R599 B.n313 B.n312 10.6151
R600 B.n314 B.n313 10.6151
R601 B.n315 B.n314 10.6151
R602 B.n317 B.n315 10.6151
R603 B.n318 B.n317 10.6151
R604 B.n319 B.n318 10.6151
R605 B.n320 B.n319 10.6151
R606 B.n321 B.n320 10.6151
R607 B.n369 B.n1 10.6151
R608 B.n369 B.n368 10.6151
R609 B.n368 B.n367 10.6151
R610 B.n367 B.n10 10.6151
R611 B.n361 B.n10 10.6151
R612 B.n361 B.n360 10.6151
R613 B.n360 B.n359 10.6151
R614 B.n359 B.n17 10.6151
R615 B.n353 B.n17 10.6151
R616 B.n353 B.n352 10.6151
R617 B.n352 B.n351 10.6151
R618 B.n351 B.n24 10.6151
R619 B.n345 B.n24 10.6151
R620 B.n345 B.n344 10.6151
R621 B.n344 B.n343 10.6151
R622 B.n343 B.n31 10.6151
R623 B.n337 B.n31 10.6151
R624 B.n337 B.n336 10.6151
R625 B.n336 B.n335 10.6151
R626 B.n335 B.n38 10.6151
R627 B.n329 B.n38 10.6151
R628 B.n329 B.n328 10.6151
R629 B.n327 B.n45 10.6151
R630 B.n66 B.n45 10.6151
R631 B.n67 B.n66 10.6151
R632 B.n70 B.n67 10.6151
R633 B.n71 B.n70 10.6151
R634 B.n74 B.n71 10.6151
R635 B.n75 B.n74 10.6151
R636 B.n79 B.n78 10.6151
R637 B.n82 B.n79 10.6151
R638 B.n83 B.n82 10.6151
R639 B.n86 B.n83 10.6151
R640 B.n87 B.n86 10.6151
R641 B.n90 B.n87 10.6151
R642 B.n91 B.n90 10.6151
R643 B.n94 B.n91 10.6151
R644 B.n99 B.n96 10.6151
R645 B.n100 B.n99 10.6151
R646 B.n103 B.n100 10.6151
R647 B.n104 B.n103 10.6151
R648 B.n107 B.n104 10.6151
R649 B.n108 B.n107 10.6151
R650 B.n322 B.n108 10.6151
R651 B.n377 B.n0 8.11757
R652 B.n377 B.n1 8.11757
R653 B.n206 B.n205 6.5566
R654 B.n189 B.n171 6.5566
R655 B.n78 B.n64 6.5566
R656 B.n95 B.n94 6.5566
R657 B.n143 B.t5 5.66574
R658 B.t9 B.n340 5.66574
R659 B.n207 B.n206 4.05904
R660 B.n186 B.n171 4.05904
R661 B.n75 B.n64 4.05904
R662 B.n96 B.n95 4.05904
R663 VP.n4 VP.n3 168.151
R664 VP.n10 VP.n9 168.151
R665 VP.n8 VP.n0 161.3
R666 VP.n7 VP.n6 161.3
R667 VP.n5 VP.n1 161.3
R668 VP.n4 VP.n2 51.4565
R669 VP.n2 VP.t3 48.223
R670 VP.n2 VP.t2 47.9894
R671 VP.n7 VP.n1 40.4934
R672 VP.n8 VP.n7 40.4934
R673 VP.n3 VP.n1 17.6167
R674 VP.n9 VP.n8 17.6167
R675 VP.n3 VP.t1 9.53647
R676 VP.n9 VP.t0 9.53647
R677 VP.n5 VP.n4 0.189894
R678 VP.n6 VP.n5 0.189894
R679 VP.n6 VP.n0 0.189894
R680 VP.n10 VP.n0 0.189894
R681 VP VP.n10 0.0516364
R682 VTAIL.n7 VTAIL.t1 252.215
R683 VTAIL.n0 VTAIL.t3 252.215
R684 VTAIL.n1 VTAIL.t5 252.215
R685 VTAIL.n2 VTAIL.t6 252.215
R686 VTAIL.n6 VTAIL.t4 252.215
R687 VTAIL.n5 VTAIL.t7 252.215
R688 VTAIL.n4 VTAIL.t2 252.215
R689 VTAIL.n3 VTAIL.t0 252.215
R690 VTAIL.n7 VTAIL.n6 14.3238
R691 VTAIL.n3 VTAIL.n2 14.3238
R692 VTAIL.n4 VTAIL.n3 1.48326
R693 VTAIL.n6 VTAIL.n5 1.48326
R694 VTAIL.n2 VTAIL.n1 1.48326
R695 VTAIL VTAIL.n0 0.800069
R696 VTAIL VTAIL.n7 0.68369
R697 VTAIL.n5 VTAIL.n4 0.470328
R698 VTAIL.n1 VTAIL.n0 0.470328
R699 VDD1 VDD1.n1 262.057
R700 VDD1 VDD1.n0 232.952
R701 VDD1.n0 VDD1.t0 36.0005
R702 VDD1.n0 VDD1.t1 36.0005
R703 VDD1.n1 VDD1.t2 36.0005
R704 VDD1.n1 VDD1.t3 36.0005
R705 VN VN.n1 51.8371
R706 VN.n0 VN.t1 48.223
R707 VN.n1 VN.t2 48.223
R708 VN.n0 VN.t3 47.9894
R709 VN.n1 VN.t0 47.9894
R710 VN VN.n0 17.5379
R711 VDD2.n2 VDD2.n0 261.531
R712 VDD2.n2 VDD2.n1 232.894
R713 VDD2.n1 VDD2.t3 36.0005
R714 VDD2.n1 VDD2.t1 36.0005
R715 VDD2.n0 VDD2.t2 36.0005
R716 VDD2.n0 VDD2.t0 36.0005
R717 VDD2 VDD2.n2 0.0586897
C0 VN VP 3.2048f
C1 VDD1 VN 0.155514f
C2 VDD2 VP 0.326396f
C3 VDD2 VDD1 0.731077f
C4 VTAIL VP 0.944071f
C5 VDD1 VTAIL 2.0255f
C6 VDD2 VN 0.48877f
C7 VDD1 VP 0.657643f
C8 VTAIL VN 0.929964f
C9 VDD2 VTAIL 2.0716f
C10 VDD2 B 2.167429f
C11 VDD1 B 4.09732f
C12 VTAIL B 2.28385f
C13 VN B 6.98266f
C14 VP B 5.329625f
C15 VDD2.t2 B 0.010664f
C16 VDD2.t0 B 0.010664f
C17 VDD2.n0 B 0.099275f
C18 VDD2.t3 B 0.010664f
C19 VDD2.t1 B 0.010664f
C20 VDD2.n1 B 0.027744f
C21 VDD2.n2 B 1.80782f
C22 VN.t1 B 0.173845f
C23 VN.t3 B 0.17309f
C24 VN.n0 B 0.115487f
C25 VN.t2 B 0.173845f
C26 VN.t0 B 0.17309f
C27 VN.n1 B 0.856541f
C28 VDD1.t0 B 0.009736f
C29 VDD1.t1 B 0.009736f
C30 VDD1.n0 B 0.025374f
C31 VDD1.t2 B 0.009736f
C32 VDD1.t3 B 0.009736f
C33 VDD1.n1 B 0.096829f
C34 VTAIL.t3 B 0.05131f
C35 VTAIL.n0 B 0.152849f
C36 VTAIL.t5 B 0.05131f
C37 VTAIL.n1 B 0.212448f
C38 VTAIL.t6 B 0.05131f
C39 VTAIL.n2 B 0.709933f
C40 VTAIL.t0 B 0.05131f
C41 VTAIL.n3 B 0.709933f
C42 VTAIL.t2 B 0.05131f
C43 VTAIL.n4 B 0.212448f
C44 VTAIL.t7 B 0.05131f
C45 VTAIL.n5 B 0.212448f
C46 VTAIL.t4 B 0.05131f
C47 VTAIL.n6 B 0.709933f
C48 VTAIL.t1 B 0.05131f
C49 VTAIL.n7 B 0.640181f
C50 VP.n0 B 0.034127f
C51 VP.t0 B 0.028804f
C52 VP.n1 B 0.059035f
C53 VP.t3 B 0.176451f
C54 VP.t2 B 0.175685f
C55 VP.n2 B 0.851537f
C56 VP.t1 B 0.028804f
C57 VP.n3 B 0.131849f
C58 VP.n4 B 1.37679f
C59 VP.n5 B 0.034127f
C60 VP.n6 B 0.034127f
C61 VP.n7 B 0.027589f
C62 VP.n8 B 0.059035f
C63 VP.n9 B 0.131849f
C64 VP.n10 B 0.029678f
.ends

