* NGSPICE file created from diff_pair_sample_0034.ext - technology: sky130A

.subckt diff_pair_sample_0034 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VN.t0 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X1 VDD1.t9 VP.t0 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=2.95515 ps=18.24 w=17.91 l=2.05
X2 VDD2.t4 VN.t1 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X3 VDD2.t3 VN.t2 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=6.9849 ps=36.6 w=17.91 l=2.05
X4 VDD2.t2 VN.t3 VTAIL.t13 B.t23 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=2.95515 ps=18.24 w=17.91 l=2.05
X5 VDD1.t8 VP.t1 VTAIL.t18 B.t22 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=2.95515 ps=18.24 w=17.91 l=2.05
X6 VTAIL.t5 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X7 B.t20 B.t18 B.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=0 ps=0 w=17.91 l=2.05
X8 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=0 ps=0 w=17.91 l=2.05
X9 VTAIL.t12 VN.t4 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X10 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=0 ps=0 w=17.91 l=2.05
X11 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=0 ps=0 w=17.91 l=2.05
X12 VDD2.t6 VN.t5 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=6.9849 pd=36.6 as=2.95515 ps=18.24 w=17.91 l=2.05
X13 VDD1.t6 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=6.9849 ps=36.6 w=17.91 l=2.05
X14 VDD1.t5 VP.t4 VTAIL.t17 B.t21 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X15 VDD2.t5 VN.t6 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=6.9849 ps=36.6 w=17.91 l=2.05
X16 VTAIL.t9 VN.t7 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X17 VDD1.t4 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X18 VTAIL.t2 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X19 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=6.9849 ps=36.6 w=17.91 l=2.05
X20 VDD2.t7 VN.t8 VTAIL.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X21 VTAIL.t3 VP.t8 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X22 VTAIL.t7 VN.t9 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
X23 VTAIL.t0 VP.t9 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.95515 pd=18.24 as=2.95515 ps=18.24 w=17.91 l=2.05
R0 VN.n8 VN.t3 241.964
R1 VN.n44 VN.t6 241.964
R2 VN.n9 VN.t7 210.553
R3 VN.n5 VN.t8 210.553
R4 VN.n26 VN.t0 210.553
R5 VN.n34 VN.t2 210.553
R6 VN.n45 VN.t9 210.553
R7 VN.n41 VN.t1 210.553
R8 VN.n62 VN.t4 210.553
R9 VN.n70 VN.t5 210.553
R10 VN.n35 VN.n34 185.279
R11 VN.n71 VN.n70 185.279
R12 VN.n69 VN.n36 161.3
R13 VN.n68 VN.n67 161.3
R14 VN.n66 VN.n37 161.3
R15 VN.n65 VN.n64 161.3
R16 VN.n63 VN.n38 161.3
R17 VN.n61 VN.n60 161.3
R18 VN.n59 VN.n39 161.3
R19 VN.n58 VN.n57 161.3
R20 VN.n56 VN.n40 161.3
R21 VN.n55 VN.n54 161.3
R22 VN.n53 VN.n52 161.3
R23 VN.n51 VN.n42 161.3
R24 VN.n50 VN.n49 161.3
R25 VN.n48 VN.n43 161.3
R26 VN.n47 VN.n46 161.3
R27 VN.n33 VN.n0 161.3
R28 VN.n32 VN.n31 161.3
R29 VN.n30 VN.n1 161.3
R30 VN.n29 VN.n28 161.3
R31 VN.n27 VN.n2 161.3
R32 VN.n25 VN.n24 161.3
R33 VN.n23 VN.n3 161.3
R34 VN.n22 VN.n21 161.3
R35 VN.n20 VN.n4 161.3
R36 VN.n19 VN.n18 161.3
R37 VN.n17 VN.n16 161.3
R38 VN.n15 VN.n6 161.3
R39 VN.n14 VN.n13 161.3
R40 VN.n12 VN.n7 161.3
R41 VN.n11 VN.n10 161.3
R42 VN.n9 VN.n8 64.109
R43 VN.n45 VN.n44 64.109
R44 VN.n28 VN.n1 56.5193
R45 VN.n64 VN.n37 56.5193
R46 VN VN.n71 54.8963
R47 VN.n15 VN.n14 46.321
R48 VN.n21 VN.n20 46.321
R49 VN.n51 VN.n50 46.321
R50 VN.n57 VN.n56 46.321
R51 VN.n14 VN.n7 34.6658
R52 VN.n21 VN.n3 34.6658
R53 VN.n50 VN.n43 34.6658
R54 VN.n57 VN.n39 34.6658
R55 VN.n10 VN.n7 24.4675
R56 VN.n16 VN.n15 24.4675
R57 VN.n20 VN.n19 24.4675
R58 VN.n25 VN.n3 24.4675
R59 VN.n28 VN.n27 24.4675
R60 VN.n32 VN.n1 24.4675
R61 VN.n33 VN.n32 24.4675
R62 VN.n46 VN.n43 24.4675
R63 VN.n56 VN.n55 24.4675
R64 VN.n52 VN.n51 24.4675
R65 VN.n64 VN.n63 24.4675
R66 VN.n61 VN.n39 24.4675
R67 VN.n69 VN.n68 24.4675
R68 VN.n68 VN.n37 24.4675
R69 VN.n27 VN.n26 18.1061
R70 VN.n63 VN.n62 18.1061
R71 VN.n47 VN.n44 12.6405
R72 VN.n11 VN.n8 12.6405
R73 VN.n16 VN.n5 12.234
R74 VN.n19 VN.n5 12.234
R75 VN.n55 VN.n41 12.234
R76 VN.n52 VN.n41 12.234
R77 VN.n10 VN.n9 6.36192
R78 VN.n26 VN.n25 6.36192
R79 VN.n46 VN.n45 6.36192
R80 VN.n62 VN.n61 6.36192
R81 VN.n34 VN.n33 0.48984
R82 VN.n70 VN.n69 0.48984
R83 VN.n71 VN.n36 0.189894
R84 VN.n67 VN.n36 0.189894
R85 VN.n67 VN.n66 0.189894
R86 VN.n66 VN.n65 0.189894
R87 VN.n65 VN.n38 0.189894
R88 VN.n60 VN.n38 0.189894
R89 VN.n60 VN.n59 0.189894
R90 VN.n59 VN.n58 0.189894
R91 VN.n58 VN.n40 0.189894
R92 VN.n54 VN.n40 0.189894
R93 VN.n54 VN.n53 0.189894
R94 VN.n53 VN.n42 0.189894
R95 VN.n49 VN.n42 0.189894
R96 VN.n49 VN.n48 0.189894
R97 VN.n48 VN.n47 0.189894
R98 VN.n12 VN.n11 0.189894
R99 VN.n13 VN.n12 0.189894
R100 VN.n13 VN.n6 0.189894
R101 VN.n17 VN.n6 0.189894
R102 VN.n18 VN.n17 0.189894
R103 VN.n18 VN.n4 0.189894
R104 VN.n22 VN.n4 0.189894
R105 VN.n23 VN.n22 0.189894
R106 VN.n24 VN.n23 0.189894
R107 VN.n24 VN.n2 0.189894
R108 VN.n29 VN.n2 0.189894
R109 VN.n30 VN.n29 0.189894
R110 VN.n31 VN.n30 0.189894
R111 VN.n31 VN.n0 0.189894
R112 VN.n35 VN.n0 0.189894
R113 VN VN.n35 0.0516364
R114 VDD2.n1 VDD2.t2 64.4028
R115 VDD2.n3 VDD2.n2 62.729
R116 VDD2 VDD2.n7 62.7262
R117 VDD2.n4 VDD2.t6 62.3513
R118 VDD2.n6 VDD2.n5 61.2458
R119 VDD2.n1 VDD2.n0 61.2456
R120 VDD2.n4 VDD2.n3 48.9006
R121 VDD2.n6 VDD2.n4 2.05222
R122 VDD2.n7 VDD2.t9 1.10603
R123 VDD2.n7 VDD2.t5 1.10603
R124 VDD2.n5 VDD2.t1 1.10603
R125 VDD2.n5 VDD2.t4 1.10603
R126 VDD2.n2 VDD2.t0 1.10603
R127 VDD2.n2 VDD2.t3 1.10603
R128 VDD2.n0 VDD2.t8 1.10603
R129 VDD2.n0 VDD2.t7 1.10603
R130 VDD2 VDD2.n6 0.571621
R131 VDD2.n3 VDD2.n1 0.458085
R132 VTAIL.n11 VTAIL.t10 45.6726
R133 VTAIL.n17 VTAIL.t14 45.6723
R134 VTAIL.n2 VTAIL.t6 45.6723
R135 VTAIL.n16 VTAIL.t1 45.6723
R136 VTAIL.n15 VTAIL.n14 44.567
R137 VTAIL.n13 VTAIL.n12 44.567
R138 VTAIL.n10 VTAIL.n9 44.567
R139 VTAIL.n8 VTAIL.n7 44.567
R140 VTAIL.n19 VTAIL.n18 44.5668
R141 VTAIL.n1 VTAIL.n0 44.5668
R142 VTAIL.n4 VTAIL.n3 44.5668
R143 VTAIL.n6 VTAIL.n5 44.5668
R144 VTAIL.n8 VTAIL.n6 31.91
R145 VTAIL.n17 VTAIL.n16 29.8583
R146 VTAIL.n10 VTAIL.n8 2.05222
R147 VTAIL.n11 VTAIL.n10 2.05222
R148 VTAIL.n15 VTAIL.n13 2.05222
R149 VTAIL.n16 VTAIL.n15 2.05222
R150 VTAIL.n6 VTAIL.n4 2.05222
R151 VTAIL.n4 VTAIL.n2 2.05222
R152 VTAIL.n19 VTAIL.n17 2.05222
R153 VTAIL VTAIL.n1 1.59748
R154 VTAIL.n13 VTAIL.n11 1.49619
R155 VTAIL.n2 VTAIL.n1 1.49619
R156 VTAIL.n18 VTAIL.t8 1.10603
R157 VTAIL.n18 VTAIL.t16 1.10603
R158 VTAIL.n0 VTAIL.t13 1.10603
R159 VTAIL.n0 VTAIL.t9 1.10603
R160 VTAIL.n3 VTAIL.t4 1.10603
R161 VTAIL.n3 VTAIL.t0 1.10603
R162 VTAIL.n5 VTAIL.t18 1.10603
R163 VTAIL.n5 VTAIL.t3 1.10603
R164 VTAIL.n14 VTAIL.t17 1.10603
R165 VTAIL.n14 VTAIL.t2 1.10603
R166 VTAIL.n12 VTAIL.t19 1.10603
R167 VTAIL.n12 VTAIL.t5 1.10603
R168 VTAIL.n9 VTAIL.t15 1.10603
R169 VTAIL.n9 VTAIL.t7 1.10603
R170 VTAIL.n7 VTAIL.t11 1.10603
R171 VTAIL.n7 VTAIL.t12 1.10603
R172 VTAIL VTAIL.n19 0.455241
R173 B.n799 B.n798 585
R174 B.n801 B.n161 585
R175 B.n804 B.n803 585
R176 B.n805 B.n160 585
R177 B.n807 B.n806 585
R178 B.n809 B.n159 585
R179 B.n812 B.n811 585
R180 B.n813 B.n158 585
R181 B.n815 B.n814 585
R182 B.n817 B.n157 585
R183 B.n820 B.n819 585
R184 B.n821 B.n156 585
R185 B.n823 B.n822 585
R186 B.n825 B.n155 585
R187 B.n828 B.n827 585
R188 B.n829 B.n154 585
R189 B.n831 B.n830 585
R190 B.n833 B.n153 585
R191 B.n836 B.n835 585
R192 B.n837 B.n152 585
R193 B.n839 B.n838 585
R194 B.n841 B.n151 585
R195 B.n844 B.n843 585
R196 B.n845 B.n150 585
R197 B.n847 B.n846 585
R198 B.n849 B.n149 585
R199 B.n852 B.n851 585
R200 B.n853 B.n148 585
R201 B.n855 B.n854 585
R202 B.n857 B.n147 585
R203 B.n860 B.n859 585
R204 B.n861 B.n146 585
R205 B.n863 B.n862 585
R206 B.n865 B.n145 585
R207 B.n868 B.n867 585
R208 B.n869 B.n144 585
R209 B.n871 B.n870 585
R210 B.n873 B.n143 585
R211 B.n876 B.n875 585
R212 B.n877 B.n142 585
R213 B.n879 B.n878 585
R214 B.n881 B.n141 585
R215 B.n884 B.n883 585
R216 B.n885 B.n140 585
R217 B.n887 B.n886 585
R218 B.n889 B.n139 585
R219 B.n892 B.n891 585
R220 B.n893 B.n138 585
R221 B.n895 B.n894 585
R222 B.n897 B.n137 585
R223 B.n900 B.n899 585
R224 B.n901 B.n136 585
R225 B.n903 B.n902 585
R226 B.n905 B.n135 585
R227 B.n908 B.n907 585
R228 B.n909 B.n134 585
R229 B.n911 B.n910 585
R230 B.n913 B.n133 585
R231 B.n916 B.n915 585
R232 B.n918 B.n130 585
R233 B.n920 B.n919 585
R234 B.n922 B.n129 585
R235 B.n925 B.n924 585
R236 B.n926 B.n128 585
R237 B.n928 B.n927 585
R238 B.n930 B.n127 585
R239 B.n933 B.n932 585
R240 B.n934 B.n123 585
R241 B.n936 B.n935 585
R242 B.n938 B.n122 585
R243 B.n941 B.n940 585
R244 B.n942 B.n121 585
R245 B.n944 B.n943 585
R246 B.n946 B.n120 585
R247 B.n949 B.n948 585
R248 B.n950 B.n119 585
R249 B.n952 B.n951 585
R250 B.n954 B.n118 585
R251 B.n957 B.n956 585
R252 B.n958 B.n117 585
R253 B.n960 B.n959 585
R254 B.n962 B.n116 585
R255 B.n965 B.n964 585
R256 B.n966 B.n115 585
R257 B.n968 B.n967 585
R258 B.n970 B.n114 585
R259 B.n973 B.n972 585
R260 B.n974 B.n113 585
R261 B.n976 B.n975 585
R262 B.n978 B.n112 585
R263 B.n981 B.n980 585
R264 B.n982 B.n111 585
R265 B.n984 B.n983 585
R266 B.n986 B.n110 585
R267 B.n989 B.n988 585
R268 B.n990 B.n109 585
R269 B.n992 B.n991 585
R270 B.n994 B.n108 585
R271 B.n997 B.n996 585
R272 B.n998 B.n107 585
R273 B.n1000 B.n999 585
R274 B.n1002 B.n106 585
R275 B.n1005 B.n1004 585
R276 B.n1006 B.n105 585
R277 B.n1008 B.n1007 585
R278 B.n1010 B.n104 585
R279 B.n1013 B.n1012 585
R280 B.n1014 B.n103 585
R281 B.n1016 B.n1015 585
R282 B.n1018 B.n102 585
R283 B.n1021 B.n1020 585
R284 B.n1022 B.n101 585
R285 B.n1024 B.n1023 585
R286 B.n1026 B.n100 585
R287 B.n1029 B.n1028 585
R288 B.n1030 B.n99 585
R289 B.n1032 B.n1031 585
R290 B.n1034 B.n98 585
R291 B.n1037 B.n1036 585
R292 B.n1038 B.n97 585
R293 B.n1040 B.n1039 585
R294 B.n1042 B.n96 585
R295 B.n1045 B.n1044 585
R296 B.n1046 B.n95 585
R297 B.n1048 B.n1047 585
R298 B.n1050 B.n94 585
R299 B.n1053 B.n1052 585
R300 B.n1054 B.n93 585
R301 B.n797 B.n91 585
R302 B.n1057 B.n91 585
R303 B.n796 B.n90 585
R304 B.n1058 B.n90 585
R305 B.n795 B.n89 585
R306 B.n1059 B.n89 585
R307 B.n794 B.n793 585
R308 B.n793 B.n85 585
R309 B.n792 B.n84 585
R310 B.n1065 B.n84 585
R311 B.n791 B.n83 585
R312 B.n1066 B.n83 585
R313 B.n790 B.n82 585
R314 B.n1067 B.n82 585
R315 B.n789 B.n788 585
R316 B.n788 B.n78 585
R317 B.n787 B.n77 585
R318 B.n1073 B.n77 585
R319 B.n786 B.n76 585
R320 B.n1074 B.n76 585
R321 B.n785 B.n75 585
R322 B.n1075 B.n75 585
R323 B.n784 B.n783 585
R324 B.n783 B.n71 585
R325 B.n782 B.n70 585
R326 B.n1081 B.n70 585
R327 B.n781 B.n69 585
R328 B.n1082 B.n69 585
R329 B.n780 B.n68 585
R330 B.n1083 B.n68 585
R331 B.n779 B.n778 585
R332 B.n778 B.n64 585
R333 B.n777 B.n63 585
R334 B.n1089 B.n63 585
R335 B.n776 B.n62 585
R336 B.n1090 B.n62 585
R337 B.n775 B.n61 585
R338 B.n1091 B.n61 585
R339 B.n774 B.n773 585
R340 B.n773 B.n57 585
R341 B.n772 B.n56 585
R342 B.n1097 B.n56 585
R343 B.n771 B.n55 585
R344 B.n1098 B.n55 585
R345 B.n770 B.n54 585
R346 B.n1099 B.n54 585
R347 B.n769 B.n768 585
R348 B.n768 B.n53 585
R349 B.n767 B.n49 585
R350 B.n1105 B.n49 585
R351 B.n766 B.n48 585
R352 B.n1106 B.n48 585
R353 B.n765 B.n47 585
R354 B.n1107 B.n47 585
R355 B.n764 B.n763 585
R356 B.n763 B.n43 585
R357 B.n762 B.n42 585
R358 B.n1113 B.n42 585
R359 B.n761 B.n41 585
R360 B.n1114 B.n41 585
R361 B.n760 B.n40 585
R362 B.n1115 B.n40 585
R363 B.n759 B.n758 585
R364 B.n758 B.n36 585
R365 B.n757 B.n35 585
R366 B.n1121 B.n35 585
R367 B.n756 B.n34 585
R368 B.n1122 B.n34 585
R369 B.n755 B.n33 585
R370 B.n1123 B.n33 585
R371 B.n754 B.n753 585
R372 B.n753 B.n29 585
R373 B.n752 B.n28 585
R374 B.n1129 B.n28 585
R375 B.n751 B.n27 585
R376 B.n1130 B.n27 585
R377 B.n750 B.n26 585
R378 B.n1131 B.n26 585
R379 B.n749 B.n748 585
R380 B.n748 B.n22 585
R381 B.n747 B.n21 585
R382 B.n1137 B.n21 585
R383 B.n746 B.n20 585
R384 B.n1138 B.n20 585
R385 B.n745 B.n19 585
R386 B.n1139 B.n19 585
R387 B.n744 B.n743 585
R388 B.n743 B.n15 585
R389 B.n742 B.n14 585
R390 B.n1145 B.n14 585
R391 B.n741 B.n13 585
R392 B.n1146 B.n13 585
R393 B.n740 B.n12 585
R394 B.n1147 B.n12 585
R395 B.n739 B.n738 585
R396 B.n738 B.n8 585
R397 B.n737 B.n7 585
R398 B.n1153 B.n7 585
R399 B.n736 B.n6 585
R400 B.n1154 B.n6 585
R401 B.n735 B.n5 585
R402 B.n1155 B.n5 585
R403 B.n734 B.n733 585
R404 B.n733 B.n4 585
R405 B.n732 B.n162 585
R406 B.n732 B.n731 585
R407 B.n722 B.n163 585
R408 B.n164 B.n163 585
R409 B.n724 B.n723 585
R410 B.n725 B.n724 585
R411 B.n721 B.n169 585
R412 B.n169 B.n168 585
R413 B.n720 B.n719 585
R414 B.n719 B.n718 585
R415 B.n171 B.n170 585
R416 B.n172 B.n171 585
R417 B.n711 B.n710 585
R418 B.n712 B.n711 585
R419 B.n709 B.n177 585
R420 B.n177 B.n176 585
R421 B.n708 B.n707 585
R422 B.n707 B.n706 585
R423 B.n179 B.n178 585
R424 B.n180 B.n179 585
R425 B.n699 B.n698 585
R426 B.n700 B.n699 585
R427 B.n697 B.n184 585
R428 B.n188 B.n184 585
R429 B.n696 B.n695 585
R430 B.n695 B.n694 585
R431 B.n186 B.n185 585
R432 B.n187 B.n186 585
R433 B.n687 B.n686 585
R434 B.n688 B.n687 585
R435 B.n685 B.n193 585
R436 B.n193 B.n192 585
R437 B.n684 B.n683 585
R438 B.n683 B.n682 585
R439 B.n195 B.n194 585
R440 B.n196 B.n195 585
R441 B.n675 B.n674 585
R442 B.n676 B.n675 585
R443 B.n673 B.n201 585
R444 B.n201 B.n200 585
R445 B.n672 B.n671 585
R446 B.n671 B.n670 585
R447 B.n203 B.n202 585
R448 B.n204 B.n203 585
R449 B.n663 B.n662 585
R450 B.n664 B.n663 585
R451 B.n661 B.n209 585
R452 B.n209 B.n208 585
R453 B.n660 B.n659 585
R454 B.n659 B.n658 585
R455 B.n211 B.n210 585
R456 B.n651 B.n211 585
R457 B.n650 B.n649 585
R458 B.n652 B.n650 585
R459 B.n648 B.n216 585
R460 B.n216 B.n215 585
R461 B.n647 B.n646 585
R462 B.n646 B.n645 585
R463 B.n218 B.n217 585
R464 B.n219 B.n218 585
R465 B.n638 B.n637 585
R466 B.n639 B.n638 585
R467 B.n636 B.n224 585
R468 B.n224 B.n223 585
R469 B.n635 B.n634 585
R470 B.n634 B.n633 585
R471 B.n226 B.n225 585
R472 B.n227 B.n226 585
R473 B.n626 B.n625 585
R474 B.n627 B.n626 585
R475 B.n624 B.n232 585
R476 B.n232 B.n231 585
R477 B.n623 B.n622 585
R478 B.n622 B.n621 585
R479 B.n234 B.n233 585
R480 B.n235 B.n234 585
R481 B.n614 B.n613 585
R482 B.n615 B.n614 585
R483 B.n612 B.n240 585
R484 B.n240 B.n239 585
R485 B.n611 B.n610 585
R486 B.n610 B.n609 585
R487 B.n242 B.n241 585
R488 B.n243 B.n242 585
R489 B.n602 B.n601 585
R490 B.n603 B.n602 585
R491 B.n600 B.n248 585
R492 B.n248 B.n247 585
R493 B.n599 B.n598 585
R494 B.n598 B.n597 585
R495 B.n250 B.n249 585
R496 B.n251 B.n250 585
R497 B.n590 B.n589 585
R498 B.n591 B.n590 585
R499 B.n588 B.n256 585
R500 B.n256 B.n255 585
R501 B.n587 B.n586 585
R502 B.n586 B.n585 585
R503 B.n582 B.n260 585
R504 B.n581 B.n580 585
R505 B.n578 B.n261 585
R506 B.n578 B.n259 585
R507 B.n577 B.n576 585
R508 B.n575 B.n574 585
R509 B.n573 B.n263 585
R510 B.n571 B.n570 585
R511 B.n569 B.n264 585
R512 B.n568 B.n567 585
R513 B.n565 B.n265 585
R514 B.n563 B.n562 585
R515 B.n561 B.n266 585
R516 B.n560 B.n559 585
R517 B.n557 B.n267 585
R518 B.n555 B.n554 585
R519 B.n553 B.n268 585
R520 B.n552 B.n551 585
R521 B.n549 B.n269 585
R522 B.n547 B.n546 585
R523 B.n545 B.n270 585
R524 B.n544 B.n543 585
R525 B.n541 B.n271 585
R526 B.n539 B.n538 585
R527 B.n537 B.n272 585
R528 B.n536 B.n535 585
R529 B.n533 B.n273 585
R530 B.n531 B.n530 585
R531 B.n529 B.n274 585
R532 B.n528 B.n527 585
R533 B.n525 B.n275 585
R534 B.n523 B.n522 585
R535 B.n521 B.n276 585
R536 B.n520 B.n519 585
R537 B.n517 B.n277 585
R538 B.n515 B.n514 585
R539 B.n513 B.n278 585
R540 B.n512 B.n511 585
R541 B.n509 B.n279 585
R542 B.n507 B.n506 585
R543 B.n505 B.n280 585
R544 B.n504 B.n503 585
R545 B.n501 B.n281 585
R546 B.n499 B.n498 585
R547 B.n497 B.n282 585
R548 B.n496 B.n495 585
R549 B.n493 B.n283 585
R550 B.n491 B.n490 585
R551 B.n489 B.n284 585
R552 B.n488 B.n487 585
R553 B.n485 B.n285 585
R554 B.n483 B.n482 585
R555 B.n481 B.n286 585
R556 B.n480 B.n479 585
R557 B.n477 B.n287 585
R558 B.n475 B.n474 585
R559 B.n473 B.n288 585
R560 B.n472 B.n471 585
R561 B.n469 B.n289 585
R562 B.n467 B.n466 585
R563 B.n464 B.n290 585
R564 B.n463 B.n462 585
R565 B.n460 B.n293 585
R566 B.n458 B.n457 585
R567 B.n456 B.n294 585
R568 B.n455 B.n454 585
R569 B.n452 B.n295 585
R570 B.n450 B.n449 585
R571 B.n448 B.n296 585
R572 B.n447 B.n446 585
R573 B.n444 B.n443 585
R574 B.n442 B.n441 585
R575 B.n440 B.n301 585
R576 B.n438 B.n437 585
R577 B.n436 B.n302 585
R578 B.n435 B.n434 585
R579 B.n432 B.n303 585
R580 B.n430 B.n429 585
R581 B.n428 B.n304 585
R582 B.n427 B.n426 585
R583 B.n424 B.n305 585
R584 B.n422 B.n421 585
R585 B.n420 B.n306 585
R586 B.n419 B.n418 585
R587 B.n416 B.n307 585
R588 B.n414 B.n413 585
R589 B.n412 B.n308 585
R590 B.n411 B.n410 585
R591 B.n408 B.n309 585
R592 B.n406 B.n405 585
R593 B.n404 B.n310 585
R594 B.n403 B.n402 585
R595 B.n400 B.n311 585
R596 B.n398 B.n397 585
R597 B.n396 B.n312 585
R598 B.n395 B.n394 585
R599 B.n392 B.n313 585
R600 B.n390 B.n389 585
R601 B.n388 B.n314 585
R602 B.n387 B.n386 585
R603 B.n384 B.n315 585
R604 B.n382 B.n381 585
R605 B.n380 B.n316 585
R606 B.n379 B.n378 585
R607 B.n376 B.n317 585
R608 B.n374 B.n373 585
R609 B.n372 B.n318 585
R610 B.n371 B.n370 585
R611 B.n368 B.n319 585
R612 B.n366 B.n365 585
R613 B.n364 B.n320 585
R614 B.n363 B.n362 585
R615 B.n360 B.n321 585
R616 B.n358 B.n357 585
R617 B.n356 B.n322 585
R618 B.n355 B.n354 585
R619 B.n352 B.n323 585
R620 B.n350 B.n349 585
R621 B.n348 B.n324 585
R622 B.n347 B.n346 585
R623 B.n344 B.n325 585
R624 B.n342 B.n341 585
R625 B.n340 B.n326 585
R626 B.n339 B.n338 585
R627 B.n336 B.n327 585
R628 B.n334 B.n333 585
R629 B.n332 B.n328 585
R630 B.n331 B.n330 585
R631 B.n258 B.n257 585
R632 B.n259 B.n258 585
R633 B.n584 B.n583 585
R634 B.n585 B.n584 585
R635 B.n254 B.n253 585
R636 B.n255 B.n254 585
R637 B.n593 B.n592 585
R638 B.n592 B.n591 585
R639 B.n594 B.n252 585
R640 B.n252 B.n251 585
R641 B.n596 B.n595 585
R642 B.n597 B.n596 585
R643 B.n246 B.n245 585
R644 B.n247 B.n246 585
R645 B.n605 B.n604 585
R646 B.n604 B.n603 585
R647 B.n606 B.n244 585
R648 B.n244 B.n243 585
R649 B.n608 B.n607 585
R650 B.n609 B.n608 585
R651 B.n238 B.n237 585
R652 B.n239 B.n238 585
R653 B.n617 B.n616 585
R654 B.n616 B.n615 585
R655 B.n618 B.n236 585
R656 B.n236 B.n235 585
R657 B.n620 B.n619 585
R658 B.n621 B.n620 585
R659 B.n230 B.n229 585
R660 B.n231 B.n230 585
R661 B.n629 B.n628 585
R662 B.n628 B.n627 585
R663 B.n630 B.n228 585
R664 B.n228 B.n227 585
R665 B.n632 B.n631 585
R666 B.n633 B.n632 585
R667 B.n222 B.n221 585
R668 B.n223 B.n222 585
R669 B.n641 B.n640 585
R670 B.n640 B.n639 585
R671 B.n642 B.n220 585
R672 B.n220 B.n219 585
R673 B.n644 B.n643 585
R674 B.n645 B.n644 585
R675 B.n214 B.n213 585
R676 B.n215 B.n214 585
R677 B.n654 B.n653 585
R678 B.n653 B.n652 585
R679 B.n655 B.n212 585
R680 B.n651 B.n212 585
R681 B.n657 B.n656 585
R682 B.n658 B.n657 585
R683 B.n207 B.n206 585
R684 B.n208 B.n207 585
R685 B.n666 B.n665 585
R686 B.n665 B.n664 585
R687 B.n667 B.n205 585
R688 B.n205 B.n204 585
R689 B.n669 B.n668 585
R690 B.n670 B.n669 585
R691 B.n199 B.n198 585
R692 B.n200 B.n199 585
R693 B.n678 B.n677 585
R694 B.n677 B.n676 585
R695 B.n679 B.n197 585
R696 B.n197 B.n196 585
R697 B.n681 B.n680 585
R698 B.n682 B.n681 585
R699 B.n191 B.n190 585
R700 B.n192 B.n191 585
R701 B.n690 B.n689 585
R702 B.n689 B.n688 585
R703 B.n691 B.n189 585
R704 B.n189 B.n187 585
R705 B.n693 B.n692 585
R706 B.n694 B.n693 585
R707 B.n183 B.n182 585
R708 B.n188 B.n183 585
R709 B.n702 B.n701 585
R710 B.n701 B.n700 585
R711 B.n703 B.n181 585
R712 B.n181 B.n180 585
R713 B.n705 B.n704 585
R714 B.n706 B.n705 585
R715 B.n175 B.n174 585
R716 B.n176 B.n175 585
R717 B.n714 B.n713 585
R718 B.n713 B.n712 585
R719 B.n715 B.n173 585
R720 B.n173 B.n172 585
R721 B.n717 B.n716 585
R722 B.n718 B.n717 585
R723 B.n167 B.n166 585
R724 B.n168 B.n167 585
R725 B.n727 B.n726 585
R726 B.n726 B.n725 585
R727 B.n728 B.n165 585
R728 B.n165 B.n164 585
R729 B.n730 B.n729 585
R730 B.n731 B.n730 585
R731 B.n2 B.n0 585
R732 B.n4 B.n2 585
R733 B.n3 B.n1 585
R734 B.n1154 B.n3 585
R735 B.n1152 B.n1151 585
R736 B.n1153 B.n1152 585
R737 B.n1150 B.n9 585
R738 B.n9 B.n8 585
R739 B.n1149 B.n1148 585
R740 B.n1148 B.n1147 585
R741 B.n11 B.n10 585
R742 B.n1146 B.n11 585
R743 B.n1144 B.n1143 585
R744 B.n1145 B.n1144 585
R745 B.n1142 B.n16 585
R746 B.n16 B.n15 585
R747 B.n1141 B.n1140 585
R748 B.n1140 B.n1139 585
R749 B.n18 B.n17 585
R750 B.n1138 B.n18 585
R751 B.n1136 B.n1135 585
R752 B.n1137 B.n1136 585
R753 B.n1134 B.n23 585
R754 B.n23 B.n22 585
R755 B.n1133 B.n1132 585
R756 B.n1132 B.n1131 585
R757 B.n25 B.n24 585
R758 B.n1130 B.n25 585
R759 B.n1128 B.n1127 585
R760 B.n1129 B.n1128 585
R761 B.n1126 B.n30 585
R762 B.n30 B.n29 585
R763 B.n1125 B.n1124 585
R764 B.n1124 B.n1123 585
R765 B.n32 B.n31 585
R766 B.n1122 B.n32 585
R767 B.n1120 B.n1119 585
R768 B.n1121 B.n1120 585
R769 B.n1118 B.n37 585
R770 B.n37 B.n36 585
R771 B.n1117 B.n1116 585
R772 B.n1116 B.n1115 585
R773 B.n39 B.n38 585
R774 B.n1114 B.n39 585
R775 B.n1112 B.n1111 585
R776 B.n1113 B.n1112 585
R777 B.n1110 B.n44 585
R778 B.n44 B.n43 585
R779 B.n1109 B.n1108 585
R780 B.n1108 B.n1107 585
R781 B.n46 B.n45 585
R782 B.n1106 B.n46 585
R783 B.n1104 B.n1103 585
R784 B.n1105 B.n1104 585
R785 B.n1102 B.n50 585
R786 B.n53 B.n50 585
R787 B.n1101 B.n1100 585
R788 B.n1100 B.n1099 585
R789 B.n52 B.n51 585
R790 B.n1098 B.n52 585
R791 B.n1096 B.n1095 585
R792 B.n1097 B.n1096 585
R793 B.n1094 B.n58 585
R794 B.n58 B.n57 585
R795 B.n1093 B.n1092 585
R796 B.n1092 B.n1091 585
R797 B.n60 B.n59 585
R798 B.n1090 B.n60 585
R799 B.n1088 B.n1087 585
R800 B.n1089 B.n1088 585
R801 B.n1086 B.n65 585
R802 B.n65 B.n64 585
R803 B.n1085 B.n1084 585
R804 B.n1084 B.n1083 585
R805 B.n67 B.n66 585
R806 B.n1082 B.n67 585
R807 B.n1080 B.n1079 585
R808 B.n1081 B.n1080 585
R809 B.n1078 B.n72 585
R810 B.n72 B.n71 585
R811 B.n1077 B.n1076 585
R812 B.n1076 B.n1075 585
R813 B.n74 B.n73 585
R814 B.n1074 B.n74 585
R815 B.n1072 B.n1071 585
R816 B.n1073 B.n1072 585
R817 B.n1070 B.n79 585
R818 B.n79 B.n78 585
R819 B.n1069 B.n1068 585
R820 B.n1068 B.n1067 585
R821 B.n81 B.n80 585
R822 B.n1066 B.n81 585
R823 B.n1064 B.n1063 585
R824 B.n1065 B.n1064 585
R825 B.n1062 B.n86 585
R826 B.n86 B.n85 585
R827 B.n1061 B.n1060 585
R828 B.n1060 B.n1059 585
R829 B.n88 B.n87 585
R830 B.n1058 B.n88 585
R831 B.n1056 B.n1055 585
R832 B.n1057 B.n1056 585
R833 B.n1157 B.n1156 585
R834 B.n1156 B.n1155 585
R835 B.n584 B.n260 482.89
R836 B.n1056 B.n93 482.89
R837 B.n586 B.n258 482.89
R838 B.n799 B.n91 482.89
R839 B.n297 B.t7 417.584
R840 B.n291 B.t18 417.584
R841 B.n124 B.t15 417.584
R842 B.n131 B.t11 417.584
R843 B.n800 B.n92 256.663
R844 B.n802 B.n92 256.663
R845 B.n808 B.n92 256.663
R846 B.n810 B.n92 256.663
R847 B.n816 B.n92 256.663
R848 B.n818 B.n92 256.663
R849 B.n824 B.n92 256.663
R850 B.n826 B.n92 256.663
R851 B.n832 B.n92 256.663
R852 B.n834 B.n92 256.663
R853 B.n840 B.n92 256.663
R854 B.n842 B.n92 256.663
R855 B.n848 B.n92 256.663
R856 B.n850 B.n92 256.663
R857 B.n856 B.n92 256.663
R858 B.n858 B.n92 256.663
R859 B.n864 B.n92 256.663
R860 B.n866 B.n92 256.663
R861 B.n872 B.n92 256.663
R862 B.n874 B.n92 256.663
R863 B.n880 B.n92 256.663
R864 B.n882 B.n92 256.663
R865 B.n888 B.n92 256.663
R866 B.n890 B.n92 256.663
R867 B.n896 B.n92 256.663
R868 B.n898 B.n92 256.663
R869 B.n904 B.n92 256.663
R870 B.n906 B.n92 256.663
R871 B.n912 B.n92 256.663
R872 B.n914 B.n92 256.663
R873 B.n921 B.n92 256.663
R874 B.n923 B.n92 256.663
R875 B.n929 B.n92 256.663
R876 B.n931 B.n92 256.663
R877 B.n937 B.n92 256.663
R878 B.n939 B.n92 256.663
R879 B.n945 B.n92 256.663
R880 B.n947 B.n92 256.663
R881 B.n953 B.n92 256.663
R882 B.n955 B.n92 256.663
R883 B.n961 B.n92 256.663
R884 B.n963 B.n92 256.663
R885 B.n969 B.n92 256.663
R886 B.n971 B.n92 256.663
R887 B.n977 B.n92 256.663
R888 B.n979 B.n92 256.663
R889 B.n985 B.n92 256.663
R890 B.n987 B.n92 256.663
R891 B.n993 B.n92 256.663
R892 B.n995 B.n92 256.663
R893 B.n1001 B.n92 256.663
R894 B.n1003 B.n92 256.663
R895 B.n1009 B.n92 256.663
R896 B.n1011 B.n92 256.663
R897 B.n1017 B.n92 256.663
R898 B.n1019 B.n92 256.663
R899 B.n1025 B.n92 256.663
R900 B.n1027 B.n92 256.663
R901 B.n1033 B.n92 256.663
R902 B.n1035 B.n92 256.663
R903 B.n1041 B.n92 256.663
R904 B.n1043 B.n92 256.663
R905 B.n1049 B.n92 256.663
R906 B.n1051 B.n92 256.663
R907 B.n579 B.n259 256.663
R908 B.n262 B.n259 256.663
R909 B.n572 B.n259 256.663
R910 B.n566 B.n259 256.663
R911 B.n564 B.n259 256.663
R912 B.n558 B.n259 256.663
R913 B.n556 B.n259 256.663
R914 B.n550 B.n259 256.663
R915 B.n548 B.n259 256.663
R916 B.n542 B.n259 256.663
R917 B.n540 B.n259 256.663
R918 B.n534 B.n259 256.663
R919 B.n532 B.n259 256.663
R920 B.n526 B.n259 256.663
R921 B.n524 B.n259 256.663
R922 B.n518 B.n259 256.663
R923 B.n516 B.n259 256.663
R924 B.n510 B.n259 256.663
R925 B.n508 B.n259 256.663
R926 B.n502 B.n259 256.663
R927 B.n500 B.n259 256.663
R928 B.n494 B.n259 256.663
R929 B.n492 B.n259 256.663
R930 B.n486 B.n259 256.663
R931 B.n484 B.n259 256.663
R932 B.n478 B.n259 256.663
R933 B.n476 B.n259 256.663
R934 B.n470 B.n259 256.663
R935 B.n468 B.n259 256.663
R936 B.n461 B.n259 256.663
R937 B.n459 B.n259 256.663
R938 B.n453 B.n259 256.663
R939 B.n451 B.n259 256.663
R940 B.n445 B.n259 256.663
R941 B.n300 B.n259 256.663
R942 B.n439 B.n259 256.663
R943 B.n433 B.n259 256.663
R944 B.n431 B.n259 256.663
R945 B.n425 B.n259 256.663
R946 B.n423 B.n259 256.663
R947 B.n417 B.n259 256.663
R948 B.n415 B.n259 256.663
R949 B.n409 B.n259 256.663
R950 B.n407 B.n259 256.663
R951 B.n401 B.n259 256.663
R952 B.n399 B.n259 256.663
R953 B.n393 B.n259 256.663
R954 B.n391 B.n259 256.663
R955 B.n385 B.n259 256.663
R956 B.n383 B.n259 256.663
R957 B.n377 B.n259 256.663
R958 B.n375 B.n259 256.663
R959 B.n369 B.n259 256.663
R960 B.n367 B.n259 256.663
R961 B.n361 B.n259 256.663
R962 B.n359 B.n259 256.663
R963 B.n353 B.n259 256.663
R964 B.n351 B.n259 256.663
R965 B.n345 B.n259 256.663
R966 B.n343 B.n259 256.663
R967 B.n337 B.n259 256.663
R968 B.n335 B.n259 256.663
R969 B.n329 B.n259 256.663
R970 B.n584 B.n254 163.367
R971 B.n592 B.n254 163.367
R972 B.n592 B.n252 163.367
R973 B.n596 B.n252 163.367
R974 B.n596 B.n246 163.367
R975 B.n604 B.n246 163.367
R976 B.n604 B.n244 163.367
R977 B.n608 B.n244 163.367
R978 B.n608 B.n238 163.367
R979 B.n616 B.n238 163.367
R980 B.n616 B.n236 163.367
R981 B.n620 B.n236 163.367
R982 B.n620 B.n230 163.367
R983 B.n628 B.n230 163.367
R984 B.n628 B.n228 163.367
R985 B.n632 B.n228 163.367
R986 B.n632 B.n222 163.367
R987 B.n640 B.n222 163.367
R988 B.n640 B.n220 163.367
R989 B.n644 B.n220 163.367
R990 B.n644 B.n214 163.367
R991 B.n653 B.n214 163.367
R992 B.n653 B.n212 163.367
R993 B.n657 B.n212 163.367
R994 B.n657 B.n207 163.367
R995 B.n665 B.n207 163.367
R996 B.n665 B.n205 163.367
R997 B.n669 B.n205 163.367
R998 B.n669 B.n199 163.367
R999 B.n677 B.n199 163.367
R1000 B.n677 B.n197 163.367
R1001 B.n681 B.n197 163.367
R1002 B.n681 B.n191 163.367
R1003 B.n689 B.n191 163.367
R1004 B.n689 B.n189 163.367
R1005 B.n693 B.n189 163.367
R1006 B.n693 B.n183 163.367
R1007 B.n701 B.n183 163.367
R1008 B.n701 B.n181 163.367
R1009 B.n705 B.n181 163.367
R1010 B.n705 B.n175 163.367
R1011 B.n713 B.n175 163.367
R1012 B.n713 B.n173 163.367
R1013 B.n717 B.n173 163.367
R1014 B.n717 B.n167 163.367
R1015 B.n726 B.n167 163.367
R1016 B.n726 B.n165 163.367
R1017 B.n730 B.n165 163.367
R1018 B.n730 B.n2 163.367
R1019 B.n1156 B.n2 163.367
R1020 B.n1156 B.n3 163.367
R1021 B.n1152 B.n3 163.367
R1022 B.n1152 B.n9 163.367
R1023 B.n1148 B.n9 163.367
R1024 B.n1148 B.n11 163.367
R1025 B.n1144 B.n11 163.367
R1026 B.n1144 B.n16 163.367
R1027 B.n1140 B.n16 163.367
R1028 B.n1140 B.n18 163.367
R1029 B.n1136 B.n18 163.367
R1030 B.n1136 B.n23 163.367
R1031 B.n1132 B.n23 163.367
R1032 B.n1132 B.n25 163.367
R1033 B.n1128 B.n25 163.367
R1034 B.n1128 B.n30 163.367
R1035 B.n1124 B.n30 163.367
R1036 B.n1124 B.n32 163.367
R1037 B.n1120 B.n32 163.367
R1038 B.n1120 B.n37 163.367
R1039 B.n1116 B.n37 163.367
R1040 B.n1116 B.n39 163.367
R1041 B.n1112 B.n39 163.367
R1042 B.n1112 B.n44 163.367
R1043 B.n1108 B.n44 163.367
R1044 B.n1108 B.n46 163.367
R1045 B.n1104 B.n46 163.367
R1046 B.n1104 B.n50 163.367
R1047 B.n1100 B.n50 163.367
R1048 B.n1100 B.n52 163.367
R1049 B.n1096 B.n52 163.367
R1050 B.n1096 B.n58 163.367
R1051 B.n1092 B.n58 163.367
R1052 B.n1092 B.n60 163.367
R1053 B.n1088 B.n60 163.367
R1054 B.n1088 B.n65 163.367
R1055 B.n1084 B.n65 163.367
R1056 B.n1084 B.n67 163.367
R1057 B.n1080 B.n67 163.367
R1058 B.n1080 B.n72 163.367
R1059 B.n1076 B.n72 163.367
R1060 B.n1076 B.n74 163.367
R1061 B.n1072 B.n74 163.367
R1062 B.n1072 B.n79 163.367
R1063 B.n1068 B.n79 163.367
R1064 B.n1068 B.n81 163.367
R1065 B.n1064 B.n81 163.367
R1066 B.n1064 B.n86 163.367
R1067 B.n1060 B.n86 163.367
R1068 B.n1060 B.n88 163.367
R1069 B.n1056 B.n88 163.367
R1070 B.n580 B.n578 163.367
R1071 B.n578 B.n577 163.367
R1072 B.n574 B.n573 163.367
R1073 B.n571 B.n264 163.367
R1074 B.n567 B.n565 163.367
R1075 B.n563 B.n266 163.367
R1076 B.n559 B.n557 163.367
R1077 B.n555 B.n268 163.367
R1078 B.n551 B.n549 163.367
R1079 B.n547 B.n270 163.367
R1080 B.n543 B.n541 163.367
R1081 B.n539 B.n272 163.367
R1082 B.n535 B.n533 163.367
R1083 B.n531 B.n274 163.367
R1084 B.n527 B.n525 163.367
R1085 B.n523 B.n276 163.367
R1086 B.n519 B.n517 163.367
R1087 B.n515 B.n278 163.367
R1088 B.n511 B.n509 163.367
R1089 B.n507 B.n280 163.367
R1090 B.n503 B.n501 163.367
R1091 B.n499 B.n282 163.367
R1092 B.n495 B.n493 163.367
R1093 B.n491 B.n284 163.367
R1094 B.n487 B.n485 163.367
R1095 B.n483 B.n286 163.367
R1096 B.n479 B.n477 163.367
R1097 B.n475 B.n288 163.367
R1098 B.n471 B.n469 163.367
R1099 B.n467 B.n290 163.367
R1100 B.n462 B.n460 163.367
R1101 B.n458 B.n294 163.367
R1102 B.n454 B.n452 163.367
R1103 B.n450 B.n296 163.367
R1104 B.n446 B.n444 163.367
R1105 B.n441 B.n440 163.367
R1106 B.n438 B.n302 163.367
R1107 B.n434 B.n432 163.367
R1108 B.n430 B.n304 163.367
R1109 B.n426 B.n424 163.367
R1110 B.n422 B.n306 163.367
R1111 B.n418 B.n416 163.367
R1112 B.n414 B.n308 163.367
R1113 B.n410 B.n408 163.367
R1114 B.n406 B.n310 163.367
R1115 B.n402 B.n400 163.367
R1116 B.n398 B.n312 163.367
R1117 B.n394 B.n392 163.367
R1118 B.n390 B.n314 163.367
R1119 B.n386 B.n384 163.367
R1120 B.n382 B.n316 163.367
R1121 B.n378 B.n376 163.367
R1122 B.n374 B.n318 163.367
R1123 B.n370 B.n368 163.367
R1124 B.n366 B.n320 163.367
R1125 B.n362 B.n360 163.367
R1126 B.n358 B.n322 163.367
R1127 B.n354 B.n352 163.367
R1128 B.n350 B.n324 163.367
R1129 B.n346 B.n344 163.367
R1130 B.n342 B.n326 163.367
R1131 B.n338 B.n336 163.367
R1132 B.n334 B.n328 163.367
R1133 B.n330 B.n258 163.367
R1134 B.n586 B.n256 163.367
R1135 B.n590 B.n256 163.367
R1136 B.n590 B.n250 163.367
R1137 B.n598 B.n250 163.367
R1138 B.n598 B.n248 163.367
R1139 B.n602 B.n248 163.367
R1140 B.n602 B.n242 163.367
R1141 B.n610 B.n242 163.367
R1142 B.n610 B.n240 163.367
R1143 B.n614 B.n240 163.367
R1144 B.n614 B.n234 163.367
R1145 B.n622 B.n234 163.367
R1146 B.n622 B.n232 163.367
R1147 B.n626 B.n232 163.367
R1148 B.n626 B.n226 163.367
R1149 B.n634 B.n226 163.367
R1150 B.n634 B.n224 163.367
R1151 B.n638 B.n224 163.367
R1152 B.n638 B.n218 163.367
R1153 B.n646 B.n218 163.367
R1154 B.n646 B.n216 163.367
R1155 B.n650 B.n216 163.367
R1156 B.n650 B.n211 163.367
R1157 B.n659 B.n211 163.367
R1158 B.n659 B.n209 163.367
R1159 B.n663 B.n209 163.367
R1160 B.n663 B.n203 163.367
R1161 B.n671 B.n203 163.367
R1162 B.n671 B.n201 163.367
R1163 B.n675 B.n201 163.367
R1164 B.n675 B.n195 163.367
R1165 B.n683 B.n195 163.367
R1166 B.n683 B.n193 163.367
R1167 B.n687 B.n193 163.367
R1168 B.n687 B.n186 163.367
R1169 B.n695 B.n186 163.367
R1170 B.n695 B.n184 163.367
R1171 B.n699 B.n184 163.367
R1172 B.n699 B.n179 163.367
R1173 B.n707 B.n179 163.367
R1174 B.n707 B.n177 163.367
R1175 B.n711 B.n177 163.367
R1176 B.n711 B.n171 163.367
R1177 B.n719 B.n171 163.367
R1178 B.n719 B.n169 163.367
R1179 B.n724 B.n169 163.367
R1180 B.n724 B.n163 163.367
R1181 B.n732 B.n163 163.367
R1182 B.n733 B.n732 163.367
R1183 B.n733 B.n5 163.367
R1184 B.n6 B.n5 163.367
R1185 B.n7 B.n6 163.367
R1186 B.n738 B.n7 163.367
R1187 B.n738 B.n12 163.367
R1188 B.n13 B.n12 163.367
R1189 B.n14 B.n13 163.367
R1190 B.n743 B.n14 163.367
R1191 B.n743 B.n19 163.367
R1192 B.n20 B.n19 163.367
R1193 B.n21 B.n20 163.367
R1194 B.n748 B.n21 163.367
R1195 B.n748 B.n26 163.367
R1196 B.n27 B.n26 163.367
R1197 B.n28 B.n27 163.367
R1198 B.n753 B.n28 163.367
R1199 B.n753 B.n33 163.367
R1200 B.n34 B.n33 163.367
R1201 B.n35 B.n34 163.367
R1202 B.n758 B.n35 163.367
R1203 B.n758 B.n40 163.367
R1204 B.n41 B.n40 163.367
R1205 B.n42 B.n41 163.367
R1206 B.n763 B.n42 163.367
R1207 B.n763 B.n47 163.367
R1208 B.n48 B.n47 163.367
R1209 B.n49 B.n48 163.367
R1210 B.n768 B.n49 163.367
R1211 B.n768 B.n54 163.367
R1212 B.n55 B.n54 163.367
R1213 B.n56 B.n55 163.367
R1214 B.n773 B.n56 163.367
R1215 B.n773 B.n61 163.367
R1216 B.n62 B.n61 163.367
R1217 B.n63 B.n62 163.367
R1218 B.n778 B.n63 163.367
R1219 B.n778 B.n68 163.367
R1220 B.n69 B.n68 163.367
R1221 B.n70 B.n69 163.367
R1222 B.n783 B.n70 163.367
R1223 B.n783 B.n75 163.367
R1224 B.n76 B.n75 163.367
R1225 B.n77 B.n76 163.367
R1226 B.n788 B.n77 163.367
R1227 B.n788 B.n82 163.367
R1228 B.n83 B.n82 163.367
R1229 B.n84 B.n83 163.367
R1230 B.n793 B.n84 163.367
R1231 B.n793 B.n89 163.367
R1232 B.n90 B.n89 163.367
R1233 B.n91 B.n90 163.367
R1234 B.n1052 B.n1050 163.367
R1235 B.n1048 B.n95 163.367
R1236 B.n1044 B.n1042 163.367
R1237 B.n1040 B.n97 163.367
R1238 B.n1036 B.n1034 163.367
R1239 B.n1032 B.n99 163.367
R1240 B.n1028 B.n1026 163.367
R1241 B.n1024 B.n101 163.367
R1242 B.n1020 B.n1018 163.367
R1243 B.n1016 B.n103 163.367
R1244 B.n1012 B.n1010 163.367
R1245 B.n1008 B.n105 163.367
R1246 B.n1004 B.n1002 163.367
R1247 B.n1000 B.n107 163.367
R1248 B.n996 B.n994 163.367
R1249 B.n992 B.n109 163.367
R1250 B.n988 B.n986 163.367
R1251 B.n984 B.n111 163.367
R1252 B.n980 B.n978 163.367
R1253 B.n976 B.n113 163.367
R1254 B.n972 B.n970 163.367
R1255 B.n968 B.n115 163.367
R1256 B.n964 B.n962 163.367
R1257 B.n960 B.n117 163.367
R1258 B.n956 B.n954 163.367
R1259 B.n952 B.n119 163.367
R1260 B.n948 B.n946 163.367
R1261 B.n944 B.n121 163.367
R1262 B.n940 B.n938 163.367
R1263 B.n936 B.n123 163.367
R1264 B.n932 B.n930 163.367
R1265 B.n928 B.n128 163.367
R1266 B.n924 B.n922 163.367
R1267 B.n920 B.n130 163.367
R1268 B.n915 B.n913 163.367
R1269 B.n911 B.n134 163.367
R1270 B.n907 B.n905 163.367
R1271 B.n903 B.n136 163.367
R1272 B.n899 B.n897 163.367
R1273 B.n895 B.n138 163.367
R1274 B.n891 B.n889 163.367
R1275 B.n887 B.n140 163.367
R1276 B.n883 B.n881 163.367
R1277 B.n879 B.n142 163.367
R1278 B.n875 B.n873 163.367
R1279 B.n871 B.n144 163.367
R1280 B.n867 B.n865 163.367
R1281 B.n863 B.n146 163.367
R1282 B.n859 B.n857 163.367
R1283 B.n855 B.n148 163.367
R1284 B.n851 B.n849 163.367
R1285 B.n847 B.n150 163.367
R1286 B.n843 B.n841 163.367
R1287 B.n839 B.n152 163.367
R1288 B.n835 B.n833 163.367
R1289 B.n831 B.n154 163.367
R1290 B.n827 B.n825 163.367
R1291 B.n823 B.n156 163.367
R1292 B.n819 B.n817 163.367
R1293 B.n815 B.n158 163.367
R1294 B.n811 B.n809 163.367
R1295 B.n807 B.n160 163.367
R1296 B.n803 B.n801 163.367
R1297 B.n297 B.t10 117.873
R1298 B.n131 B.t13 117.873
R1299 B.n291 B.t20 117.849
R1300 B.n124 B.t16 117.849
R1301 B.n298 B.t9 71.7145
R1302 B.n132 B.t14 71.7145
R1303 B.n292 B.t19 71.6908
R1304 B.n125 B.t17 71.6908
R1305 B.n579 B.n260 71.676
R1306 B.n577 B.n262 71.676
R1307 B.n573 B.n572 71.676
R1308 B.n566 B.n264 71.676
R1309 B.n565 B.n564 71.676
R1310 B.n558 B.n266 71.676
R1311 B.n557 B.n556 71.676
R1312 B.n550 B.n268 71.676
R1313 B.n549 B.n548 71.676
R1314 B.n542 B.n270 71.676
R1315 B.n541 B.n540 71.676
R1316 B.n534 B.n272 71.676
R1317 B.n533 B.n532 71.676
R1318 B.n526 B.n274 71.676
R1319 B.n525 B.n524 71.676
R1320 B.n518 B.n276 71.676
R1321 B.n517 B.n516 71.676
R1322 B.n510 B.n278 71.676
R1323 B.n509 B.n508 71.676
R1324 B.n502 B.n280 71.676
R1325 B.n501 B.n500 71.676
R1326 B.n494 B.n282 71.676
R1327 B.n493 B.n492 71.676
R1328 B.n486 B.n284 71.676
R1329 B.n485 B.n484 71.676
R1330 B.n478 B.n286 71.676
R1331 B.n477 B.n476 71.676
R1332 B.n470 B.n288 71.676
R1333 B.n469 B.n468 71.676
R1334 B.n461 B.n290 71.676
R1335 B.n460 B.n459 71.676
R1336 B.n453 B.n294 71.676
R1337 B.n452 B.n451 71.676
R1338 B.n445 B.n296 71.676
R1339 B.n444 B.n300 71.676
R1340 B.n440 B.n439 71.676
R1341 B.n433 B.n302 71.676
R1342 B.n432 B.n431 71.676
R1343 B.n425 B.n304 71.676
R1344 B.n424 B.n423 71.676
R1345 B.n417 B.n306 71.676
R1346 B.n416 B.n415 71.676
R1347 B.n409 B.n308 71.676
R1348 B.n408 B.n407 71.676
R1349 B.n401 B.n310 71.676
R1350 B.n400 B.n399 71.676
R1351 B.n393 B.n312 71.676
R1352 B.n392 B.n391 71.676
R1353 B.n385 B.n314 71.676
R1354 B.n384 B.n383 71.676
R1355 B.n377 B.n316 71.676
R1356 B.n376 B.n375 71.676
R1357 B.n369 B.n318 71.676
R1358 B.n368 B.n367 71.676
R1359 B.n361 B.n320 71.676
R1360 B.n360 B.n359 71.676
R1361 B.n353 B.n322 71.676
R1362 B.n352 B.n351 71.676
R1363 B.n345 B.n324 71.676
R1364 B.n344 B.n343 71.676
R1365 B.n337 B.n326 71.676
R1366 B.n336 B.n335 71.676
R1367 B.n329 B.n328 71.676
R1368 B.n1051 B.n93 71.676
R1369 B.n1050 B.n1049 71.676
R1370 B.n1043 B.n95 71.676
R1371 B.n1042 B.n1041 71.676
R1372 B.n1035 B.n97 71.676
R1373 B.n1034 B.n1033 71.676
R1374 B.n1027 B.n99 71.676
R1375 B.n1026 B.n1025 71.676
R1376 B.n1019 B.n101 71.676
R1377 B.n1018 B.n1017 71.676
R1378 B.n1011 B.n103 71.676
R1379 B.n1010 B.n1009 71.676
R1380 B.n1003 B.n105 71.676
R1381 B.n1002 B.n1001 71.676
R1382 B.n995 B.n107 71.676
R1383 B.n994 B.n993 71.676
R1384 B.n987 B.n109 71.676
R1385 B.n986 B.n985 71.676
R1386 B.n979 B.n111 71.676
R1387 B.n978 B.n977 71.676
R1388 B.n971 B.n113 71.676
R1389 B.n970 B.n969 71.676
R1390 B.n963 B.n115 71.676
R1391 B.n962 B.n961 71.676
R1392 B.n955 B.n117 71.676
R1393 B.n954 B.n953 71.676
R1394 B.n947 B.n119 71.676
R1395 B.n946 B.n945 71.676
R1396 B.n939 B.n121 71.676
R1397 B.n938 B.n937 71.676
R1398 B.n931 B.n123 71.676
R1399 B.n930 B.n929 71.676
R1400 B.n923 B.n128 71.676
R1401 B.n922 B.n921 71.676
R1402 B.n914 B.n130 71.676
R1403 B.n913 B.n912 71.676
R1404 B.n906 B.n134 71.676
R1405 B.n905 B.n904 71.676
R1406 B.n898 B.n136 71.676
R1407 B.n897 B.n896 71.676
R1408 B.n890 B.n138 71.676
R1409 B.n889 B.n888 71.676
R1410 B.n882 B.n140 71.676
R1411 B.n881 B.n880 71.676
R1412 B.n874 B.n142 71.676
R1413 B.n873 B.n872 71.676
R1414 B.n866 B.n144 71.676
R1415 B.n865 B.n864 71.676
R1416 B.n858 B.n146 71.676
R1417 B.n857 B.n856 71.676
R1418 B.n850 B.n148 71.676
R1419 B.n849 B.n848 71.676
R1420 B.n842 B.n150 71.676
R1421 B.n841 B.n840 71.676
R1422 B.n834 B.n152 71.676
R1423 B.n833 B.n832 71.676
R1424 B.n826 B.n154 71.676
R1425 B.n825 B.n824 71.676
R1426 B.n818 B.n156 71.676
R1427 B.n817 B.n816 71.676
R1428 B.n810 B.n158 71.676
R1429 B.n809 B.n808 71.676
R1430 B.n802 B.n160 71.676
R1431 B.n801 B.n800 71.676
R1432 B.n800 B.n799 71.676
R1433 B.n803 B.n802 71.676
R1434 B.n808 B.n807 71.676
R1435 B.n811 B.n810 71.676
R1436 B.n816 B.n815 71.676
R1437 B.n819 B.n818 71.676
R1438 B.n824 B.n823 71.676
R1439 B.n827 B.n826 71.676
R1440 B.n832 B.n831 71.676
R1441 B.n835 B.n834 71.676
R1442 B.n840 B.n839 71.676
R1443 B.n843 B.n842 71.676
R1444 B.n848 B.n847 71.676
R1445 B.n851 B.n850 71.676
R1446 B.n856 B.n855 71.676
R1447 B.n859 B.n858 71.676
R1448 B.n864 B.n863 71.676
R1449 B.n867 B.n866 71.676
R1450 B.n872 B.n871 71.676
R1451 B.n875 B.n874 71.676
R1452 B.n880 B.n879 71.676
R1453 B.n883 B.n882 71.676
R1454 B.n888 B.n887 71.676
R1455 B.n891 B.n890 71.676
R1456 B.n896 B.n895 71.676
R1457 B.n899 B.n898 71.676
R1458 B.n904 B.n903 71.676
R1459 B.n907 B.n906 71.676
R1460 B.n912 B.n911 71.676
R1461 B.n915 B.n914 71.676
R1462 B.n921 B.n920 71.676
R1463 B.n924 B.n923 71.676
R1464 B.n929 B.n928 71.676
R1465 B.n932 B.n931 71.676
R1466 B.n937 B.n936 71.676
R1467 B.n940 B.n939 71.676
R1468 B.n945 B.n944 71.676
R1469 B.n948 B.n947 71.676
R1470 B.n953 B.n952 71.676
R1471 B.n956 B.n955 71.676
R1472 B.n961 B.n960 71.676
R1473 B.n964 B.n963 71.676
R1474 B.n969 B.n968 71.676
R1475 B.n972 B.n971 71.676
R1476 B.n977 B.n976 71.676
R1477 B.n980 B.n979 71.676
R1478 B.n985 B.n984 71.676
R1479 B.n988 B.n987 71.676
R1480 B.n993 B.n992 71.676
R1481 B.n996 B.n995 71.676
R1482 B.n1001 B.n1000 71.676
R1483 B.n1004 B.n1003 71.676
R1484 B.n1009 B.n1008 71.676
R1485 B.n1012 B.n1011 71.676
R1486 B.n1017 B.n1016 71.676
R1487 B.n1020 B.n1019 71.676
R1488 B.n1025 B.n1024 71.676
R1489 B.n1028 B.n1027 71.676
R1490 B.n1033 B.n1032 71.676
R1491 B.n1036 B.n1035 71.676
R1492 B.n1041 B.n1040 71.676
R1493 B.n1044 B.n1043 71.676
R1494 B.n1049 B.n1048 71.676
R1495 B.n1052 B.n1051 71.676
R1496 B.n580 B.n579 71.676
R1497 B.n574 B.n262 71.676
R1498 B.n572 B.n571 71.676
R1499 B.n567 B.n566 71.676
R1500 B.n564 B.n563 71.676
R1501 B.n559 B.n558 71.676
R1502 B.n556 B.n555 71.676
R1503 B.n551 B.n550 71.676
R1504 B.n548 B.n547 71.676
R1505 B.n543 B.n542 71.676
R1506 B.n540 B.n539 71.676
R1507 B.n535 B.n534 71.676
R1508 B.n532 B.n531 71.676
R1509 B.n527 B.n526 71.676
R1510 B.n524 B.n523 71.676
R1511 B.n519 B.n518 71.676
R1512 B.n516 B.n515 71.676
R1513 B.n511 B.n510 71.676
R1514 B.n508 B.n507 71.676
R1515 B.n503 B.n502 71.676
R1516 B.n500 B.n499 71.676
R1517 B.n495 B.n494 71.676
R1518 B.n492 B.n491 71.676
R1519 B.n487 B.n486 71.676
R1520 B.n484 B.n483 71.676
R1521 B.n479 B.n478 71.676
R1522 B.n476 B.n475 71.676
R1523 B.n471 B.n470 71.676
R1524 B.n468 B.n467 71.676
R1525 B.n462 B.n461 71.676
R1526 B.n459 B.n458 71.676
R1527 B.n454 B.n453 71.676
R1528 B.n451 B.n450 71.676
R1529 B.n446 B.n445 71.676
R1530 B.n441 B.n300 71.676
R1531 B.n439 B.n438 71.676
R1532 B.n434 B.n433 71.676
R1533 B.n431 B.n430 71.676
R1534 B.n426 B.n425 71.676
R1535 B.n423 B.n422 71.676
R1536 B.n418 B.n417 71.676
R1537 B.n415 B.n414 71.676
R1538 B.n410 B.n409 71.676
R1539 B.n407 B.n406 71.676
R1540 B.n402 B.n401 71.676
R1541 B.n399 B.n398 71.676
R1542 B.n394 B.n393 71.676
R1543 B.n391 B.n390 71.676
R1544 B.n386 B.n385 71.676
R1545 B.n383 B.n382 71.676
R1546 B.n378 B.n377 71.676
R1547 B.n375 B.n374 71.676
R1548 B.n370 B.n369 71.676
R1549 B.n367 B.n366 71.676
R1550 B.n362 B.n361 71.676
R1551 B.n359 B.n358 71.676
R1552 B.n354 B.n353 71.676
R1553 B.n351 B.n350 71.676
R1554 B.n346 B.n345 71.676
R1555 B.n343 B.n342 71.676
R1556 B.n338 B.n337 71.676
R1557 B.n335 B.n334 71.676
R1558 B.n330 B.n329 71.676
R1559 B.n585 B.n259 62.1528
R1560 B.n1057 B.n92 62.1528
R1561 B.n299 B.n298 59.5399
R1562 B.n465 B.n292 59.5399
R1563 B.n126 B.n125 59.5399
R1564 B.n917 B.n132 59.5399
R1565 B.n298 B.n297 46.1581
R1566 B.n292 B.n291 46.1581
R1567 B.n125 B.n124 46.1581
R1568 B.n132 B.n131 46.1581
R1569 B.n585 B.n255 32.2627
R1570 B.n591 B.n255 32.2627
R1571 B.n591 B.n251 32.2627
R1572 B.n597 B.n251 32.2627
R1573 B.n597 B.n247 32.2627
R1574 B.n603 B.n247 32.2627
R1575 B.n609 B.n243 32.2627
R1576 B.n609 B.n239 32.2627
R1577 B.n615 B.n239 32.2627
R1578 B.n615 B.n235 32.2627
R1579 B.n621 B.n235 32.2627
R1580 B.n621 B.n231 32.2627
R1581 B.n627 B.n231 32.2627
R1582 B.n627 B.n227 32.2627
R1583 B.n633 B.n227 32.2627
R1584 B.n639 B.n223 32.2627
R1585 B.n639 B.n219 32.2627
R1586 B.n645 B.n219 32.2627
R1587 B.n645 B.n215 32.2627
R1588 B.n652 B.n215 32.2627
R1589 B.n652 B.n651 32.2627
R1590 B.n658 B.n208 32.2627
R1591 B.n664 B.n208 32.2627
R1592 B.n664 B.n204 32.2627
R1593 B.n670 B.n204 32.2627
R1594 B.n670 B.n200 32.2627
R1595 B.n676 B.n200 32.2627
R1596 B.n682 B.n196 32.2627
R1597 B.n682 B.n192 32.2627
R1598 B.n688 B.n192 32.2627
R1599 B.n688 B.n187 32.2627
R1600 B.n694 B.n187 32.2627
R1601 B.n694 B.n188 32.2627
R1602 B.n700 B.n180 32.2627
R1603 B.n706 B.n180 32.2627
R1604 B.n706 B.n176 32.2627
R1605 B.n712 B.n176 32.2627
R1606 B.n712 B.n172 32.2627
R1607 B.n718 B.n172 32.2627
R1608 B.n725 B.n168 32.2627
R1609 B.n725 B.n164 32.2627
R1610 B.n731 B.n164 32.2627
R1611 B.n731 B.n4 32.2627
R1612 B.n1155 B.n4 32.2627
R1613 B.n1155 B.n1154 32.2627
R1614 B.n1154 B.n1153 32.2627
R1615 B.n1153 B.n8 32.2627
R1616 B.n1147 B.n8 32.2627
R1617 B.n1147 B.n1146 32.2627
R1618 B.n1145 B.n15 32.2627
R1619 B.n1139 B.n15 32.2627
R1620 B.n1139 B.n1138 32.2627
R1621 B.n1138 B.n1137 32.2627
R1622 B.n1137 B.n22 32.2627
R1623 B.n1131 B.n22 32.2627
R1624 B.n1130 B.n1129 32.2627
R1625 B.n1129 B.n29 32.2627
R1626 B.n1123 B.n29 32.2627
R1627 B.n1123 B.n1122 32.2627
R1628 B.n1122 B.n1121 32.2627
R1629 B.n1121 B.n36 32.2627
R1630 B.n1115 B.n1114 32.2627
R1631 B.n1114 B.n1113 32.2627
R1632 B.n1113 B.n43 32.2627
R1633 B.n1107 B.n43 32.2627
R1634 B.n1107 B.n1106 32.2627
R1635 B.n1106 B.n1105 32.2627
R1636 B.n1099 B.n53 32.2627
R1637 B.n1099 B.n1098 32.2627
R1638 B.n1098 B.n1097 32.2627
R1639 B.n1097 B.n57 32.2627
R1640 B.n1091 B.n57 32.2627
R1641 B.n1091 B.n1090 32.2627
R1642 B.n1089 B.n64 32.2627
R1643 B.n1083 B.n64 32.2627
R1644 B.n1083 B.n1082 32.2627
R1645 B.n1082 B.n1081 32.2627
R1646 B.n1081 B.n71 32.2627
R1647 B.n1075 B.n71 32.2627
R1648 B.n1075 B.n1074 32.2627
R1649 B.n1074 B.n1073 32.2627
R1650 B.n1073 B.n78 32.2627
R1651 B.n1067 B.n1066 32.2627
R1652 B.n1066 B.n1065 32.2627
R1653 B.n1065 B.n85 32.2627
R1654 B.n1059 B.n85 32.2627
R1655 B.n1059 B.n1058 32.2627
R1656 B.n1058 B.n1057 32.2627
R1657 B.n1055 B.n1054 31.3761
R1658 B.n798 B.n797 31.3761
R1659 B.n587 B.n257 31.3761
R1660 B.n583 B.n582 31.3761
R1661 B.n633 B.t22 28.9416
R1662 B.n651 B.t3 28.9416
R1663 B.n676 B.t4 28.9416
R1664 B.n188 B.t0 28.9416
R1665 B.n718 B.t6 28.9416
R1666 B.t23 B.n1145 28.9416
R1667 B.t5 B.n1130 28.9416
R1668 B.n1115 B.t21 28.9416
R1669 B.n53 B.t2 28.9416
R1670 B.t1 B.n1089 28.9416
R1671 B.n603 B.t8 22.2994
R1672 B.n1067 B.t12 22.2994
R1673 B B.n1157 18.0485
R1674 B.n1054 B.n1053 10.6151
R1675 B.n1053 B.n94 10.6151
R1676 B.n1047 B.n94 10.6151
R1677 B.n1047 B.n1046 10.6151
R1678 B.n1046 B.n1045 10.6151
R1679 B.n1045 B.n96 10.6151
R1680 B.n1039 B.n96 10.6151
R1681 B.n1039 B.n1038 10.6151
R1682 B.n1038 B.n1037 10.6151
R1683 B.n1037 B.n98 10.6151
R1684 B.n1031 B.n98 10.6151
R1685 B.n1031 B.n1030 10.6151
R1686 B.n1030 B.n1029 10.6151
R1687 B.n1029 B.n100 10.6151
R1688 B.n1023 B.n100 10.6151
R1689 B.n1023 B.n1022 10.6151
R1690 B.n1022 B.n1021 10.6151
R1691 B.n1021 B.n102 10.6151
R1692 B.n1015 B.n102 10.6151
R1693 B.n1015 B.n1014 10.6151
R1694 B.n1014 B.n1013 10.6151
R1695 B.n1013 B.n104 10.6151
R1696 B.n1007 B.n104 10.6151
R1697 B.n1007 B.n1006 10.6151
R1698 B.n1006 B.n1005 10.6151
R1699 B.n1005 B.n106 10.6151
R1700 B.n999 B.n106 10.6151
R1701 B.n999 B.n998 10.6151
R1702 B.n998 B.n997 10.6151
R1703 B.n997 B.n108 10.6151
R1704 B.n991 B.n108 10.6151
R1705 B.n991 B.n990 10.6151
R1706 B.n990 B.n989 10.6151
R1707 B.n989 B.n110 10.6151
R1708 B.n983 B.n110 10.6151
R1709 B.n983 B.n982 10.6151
R1710 B.n982 B.n981 10.6151
R1711 B.n981 B.n112 10.6151
R1712 B.n975 B.n112 10.6151
R1713 B.n975 B.n974 10.6151
R1714 B.n974 B.n973 10.6151
R1715 B.n973 B.n114 10.6151
R1716 B.n967 B.n114 10.6151
R1717 B.n967 B.n966 10.6151
R1718 B.n966 B.n965 10.6151
R1719 B.n965 B.n116 10.6151
R1720 B.n959 B.n116 10.6151
R1721 B.n959 B.n958 10.6151
R1722 B.n958 B.n957 10.6151
R1723 B.n957 B.n118 10.6151
R1724 B.n951 B.n118 10.6151
R1725 B.n951 B.n950 10.6151
R1726 B.n950 B.n949 10.6151
R1727 B.n949 B.n120 10.6151
R1728 B.n943 B.n120 10.6151
R1729 B.n943 B.n942 10.6151
R1730 B.n942 B.n941 10.6151
R1731 B.n941 B.n122 10.6151
R1732 B.n935 B.n934 10.6151
R1733 B.n934 B.n933 10.6151
R1734 B.n933 B.n127 10.6151
R1735 B.n927 B.n127 10.6151
R1736 B.n927 B.n926 10.6151
R1737 B.n926 B.n925 10.6151
R1738 B.n925 B.n129 10.6151
R1739 B.n919 B.n129 10.6151
R1740 B.n919 B.n918 10.6151
R1741 B.n916 B.n133 10.6151
R1742 B.n910 B.n133 10.6151
R1743 B.n910 B.n909 10.6151
R1744 B.n909 B.n908 10.6151
R1745 B.n908 B.n135 10.6151
R1746 B.n902 B.n135 10.6151
R1747 B.n902 B.n901 10.6151
R1748 B.n901 B.n900 10.6151
R1749 B.n900 B.n137 10.6151
R1750 B.n894 B.n137 10.6151
R1751 B.n894 B.n893 10.6151
R1752 B.n893 B.n892 10.6151
R1753 B.n892 B.n139 10.6151
R1754 B.n886 B.n139 10.6151
R1755 B.n886 B.n885 10.6151
R1756 B.n885 B.n884 10.6151
R1757 B.n884 B.n141 10.6151
R1758 B.n878 B.n141 10.6151
R1759 B.n878 B.n877 10.6151
R1760 B.n877 B.n876 10.6151
R1761 B.n876 B.n143 10.6151
R1762 B.n870 B.n143 10.6151
R1763 B.n870 B.n869 10.6151
R1764 B.n869 B.n868 10.6151
R1765 B.n868 B.n145 10.6151
R1766 B.n862 B.n145 10.6151
R1767 B.n862 B.n861 10.6151
R1768 B.n861 B.n860 10.6151
R1769 B.n860 B.n147 10.6151
R1770 B.n854 B.n147 10.6151
R1771 B.n854 B.n853 10.6151
R1772 B.n853 B.n852 10.6151
R1773 B.n852 B.n149 10.6151
R1774 B.n846 B.n149 10.6151
R1775 B.n846 B.n845 10.6151
R1776 B.n845 B.n844 10.6151
R1777 B.n844 B.n151 10.6151
R1778 B.n838 B.n151 10.6151
R1779 B.n838 B.n837 10.6151
R1780 B.n837 B.n836 10.6151
R1781 B.n836 B.n153 10.6151
R1782 B.n830 B.n153 10.6151
R1783 B.n830 B.n829 10.6151
R1784 B.n829 B.n828 10.6151
R1785 B.n828 B.n155 10.6151
R1786 B.n822 B.n155 10.6151
R1787 B.n822 B.n821 10.6151
R1788 B.n821 B.n820 10.6151
R1789 B.n820 B.n157 10.6151
R1790 B.n814 B.n157 10.6151
R1791 B.n814 B.n813 10.6151
R1792 B.n813 B.n812 10.6151
R1793 B.n812 B.n159 10.6151
R1794 B.n806 B.n159 10.6151
R1795 B.n806 B.n805 10.6151
R1796 B.n805 B.n804 10.6151
R1797 B.n804 B.n161 10.6151
R1798 B.n798 B.n161 10.6151
R1799 B.n588 B.n587 10.6151
R1800 B.n589 B.n588 10.6151
R1801 B.n589 B.n249 10.6151
R1802 B.n599 B.n249 10.6151
R1803 B.n600 B.n599 10.6151
R1804 B.n601 B.n600 10.6151
R1805 B.n601 B.n241 10.6151
R1806 B.n611 B.n241 10.6151
R1807 B.n612 B.n611 10.6151
R1808 B.n613 B.n612 10.6151
R1809 B.n613 B.n233 10.6151
R1810 B.n623 B.n233 10.6151
R1811 B.n624 B.n623 10.6151
R1812 B.n625 B.n624 10.6151
R1813 B.n625 B.n225 10.6151
R1814 B.n635 B.n225 10.6151
R1815 B.n636 B.n635 10.6151
R1816 B.n637 B.n636 10.6151
R1817 B.n637 B.n217 10.6151
R1818 B.n647 B.n217 10.6151
R1819 B.n648 B.n647 10.6151
R1820 B.n649 B.n648 10.6151
R1821 B.n649 B.n210 10.6151
R1822 B.n660 B.n210 10.6151
R1823 B.n661 B.n660 10.6151
R1824 B.n662 B.n661 10.6151
R1825 B.n662 B.n202 10.6151
R1826 B.n672 B.n202 10.6151
R1827 B.n673 B.n672 10.6151
R1828 B.n674 B.n673 10.6151
R1829 B.n674 B.n194 10.6151
R1830 B.n684 B.n194 10.6151
R1831 B.n685 B.n684 10.6151
R1832 B.n686 B.n685 10.6151
R1833 B.n686 B.n185 10.6151
R1834 B.n696 B.n185 10.6151
R1835 B.n697 B.n696 10.6151
R1836 B.n698 B.n697 10.6151
R1837 B.n698 B.n178 10.6151
R1838 B.n708 B.n178 10.6151
R1839 B.n709 B.n708 10.6151
R1840 B.n710 B.n709 10.6151
R1841 B.n710 B.n170 10.6151
R1842 B.n720 B.n170 10.6151
R1843 B.n721 B.n720 10.6151
R1844 B.n723 B.n721 10.6151
R1845 B.n723 B.n722 10.6151
R1846 B.n722 B.n162 10.6151
R1847 B.n734 B.n162 10.6151
R1848 B.n735 B.n734 10.6151
R1849 B.n736 B.n735 10.6151
R1850 B.n737 B.n736 10.6151
R1851 B.n739 B.n737 10.6151
R1852 B.n740 B.n739 10.6151
R1853 B.n741 B.n740 10.6151
R1854 B.n742 B.n741 10.6151
R1855 B.n744 B.n742 10.6151
R1856 B.n745 B.n744 10.6151
R1857 B.n746 B.n745 10.6151
R1858 B.n747 B.n746 10.6151
R1859 B.n749 B.n747 10.6151
R1860 B.n750 B.n749 10.6151
R1861 B.n751 B.n750 10.6151
R1862 B.n752 B.n751 10.6151
R1863 B.n754 B.n752 10.6151
R1864 B.n755 B.n754 10.6151
R1865 B.n756 B.n755 10.6151
R1866 B.n757 B.n756 10.6151
R1867 B.n759 B.n757 10.6151
R1868 B.n760 B.n759 10.6151
R1869 B.n761 B.n760 10.6151
R1870 B.n762 B.n761 10.6151
R1871 B.n764 B.n762 10.6151
R1872 B.n765 B.n764 10.6151
R1873 B.n766 B.n765 10.6151
R1874 B.n767 B.n766 10.6151
R1875 B.n769 B.n767 10.6151
R1876 B.n770 B.n769 10.6151
R1877 B.n771 B.n770 10.6151
R1878 B.n772 B.n771 10.6151
R1879 B.n774 B.n772 10.6151
R1880 B.n775 B.n774 10.6151
R1881 B.n776 B.n775 10.6151
R1882 B.n777 B.n776 10.6151
R1883 B.n779 B.n777 10.6151
R1884 B.n780 B.n779 10.6151
R1885 B.n781 B.n780 10.6151
R1886 B.n782 B.n781 10.6151
R1887 B.n784 B.n782 10.6151
R1888 B.n785 B.n784 10.6151
R1889 B.n786 B.n785 10.6151
R1890 B.n787 B.n786 10.6151
R1891 B.n789 B.n787 10.6151
R1892 B.n790 B.n789 10.6151
R1893 B.n791 B.n790 10.6151
R1894 B.n792 B.n791 10.6151
R1895 B.n794 B.n792 10.6151
R1896 B.n795 B.n794 10.6151
R1897 B.n796 B.n795 10.6151
R1898 B.n797 B.n796 10.6151
R1899 B.n582 B.n581 10.6151
R1900 B.n581 B.n261 10.6151
R1901 B.n576 B.n261 10.6151
R1902 B.n576 B.n575 10.6151
R1903 B.n575 B.n263 10.6151
R1904 B.n570 B.n263 10.6151
R1905 B.n570 B.n569 10.6151
R1906 B.n569 B.n568 10.6151
R1907 B.n568 B.n265 10.6151
R1908 B.n562 B.n265 10.6151
R1909 B.n562 B.n561 10.6151
R1910 B.n561 B.n560 10.6151
R1911 B.n560 B.n267 10.6151
R1912 B.n554 B.n267 10.6151
R1913 B.n554 B.n553 10.6151
R1914 B.n553 B.n552 10.6151
R1915 B.n552 B.n269 10.6151
R1916 B.n546 B.n269 10.6151
R1917 B.n546 B.n545 10.6151
R1918 B.n545 B.n544 10.6151
R1919 B.n544 B.n271 10.6151
R1920 B.n538 B.n271 10.6151
R1921 B.n538 B.n537 10.6151
R1922 B.n537 B.n536 10.6151
R1923 B.n536 B.n273 10.6151
R1924 B.n530 B.n273 10.6151
R1925 B.n530 B.n529 10.6151
R1926 B.n529 B.n528 10.6151
R1927 B.n528 B.n275 10.6151
R1928 B.n522 B.n275 10.6151
R1929 B.n522 B.n521 10.6151
R1930 B.n521 B.n520 10.6151
R1931 B.n520 B.n277 10.6151
R1932 B.n514 B.n277 10.6151
R1933 B.n514 B.n513 10.6151
R1934 B.n513 B.n512 10.6151
R1935 B.n512 B.n279 10.6151
R1936 B.n506 B.n279 10.6151
R1937 B.n506 B.n505 10.6151
R1938 B.n505 B.n504 10.6151
R1939 B.n504 B.n281 10.6151
R1940 B.n498 B.n281 10.6151
R1941 B.n498 B.n497 10.6151
R1942 B.n497 B.n496 10.6151
R1943 B.n496 B.n283 10.6151
R1944 B.n490 B.n283 10.6151
R1945 B.n490 B.n489 10.6151
R1946 B.n489 B.n488 10.6151
R1947 B.n488 B.n285 10.6151
R1948 B.n482 B.n285 10.6151
R1949 B.n482 B.n481 10.6151
R1950 B.n481 B.n480 10.6151
R1951 B.n480 B.n287 10.6151
R1952 B.n474 B.n287 10.6151
R1953 B.n474 B.n473 10.6151
R1954 B.n473 B.n472 10.6151
R1955 B.n472 B.n289 10.6151
R1956 B.n466 B.n289 10.6151
R1957 B.n464 B.n463 10.6151
R1958 B.n463 B.n293 10.6151
R1959 B.n457 B.n293 10.6151
R1960 B.n457 B.n456 10.6151
R1961 B.n456 B.n455 10.6151
R1962 B.n455 B.n295 10.6151
R1963 B.n449 B.n295 10.6151
R1964 B.n449 B.n448 10.6151
R1965 B.n448 B.n447 10.6151
R1966 B.n443 B.n442 10.6151
R1967 B.n442 B.n301 10.6151
R1968 B.n437 B.n301 10.6151
R1969 B.n437 B.n436 10.6151
R1970 B.n436 B.n435 10.6151
R1971 B.n435 B.n303 10.6151
R1972 B.n429 B.n303 10.6151
R1973 B.n429 B.n428 10.6151
R1974 B.n428 B.n427 10.6151
R1975 B.n427 B.n305 10.6151
R1976 B.n421 B.n305 10.6151
R1977 B.n421 B.n420 10.6151
R1978 B.n420 B.n419 10.6151
R1979 B.n419 B.n307 10.6151
R1980 B.n413 B.n307 10.6151
R1981 B.n413 B.n412 10.6151
R1982 B.n412 B.n411 10.6151
R1983 B.n411 B.n309 10.6151
R1984 B.n405 B.n309 10.6151
R1985 B.n405 B.n404 10.6151
R1986 B.n404 B.n403 10.6151
R1987 B.n403 B.n311 10.6151
R1988 B.n397 B.n311 10.6151
R1989 B.n397 B.n396 10.6151
R1990 B.n396 B.n395 10.6151
R1991 B.n395 B.n313 10.6151
R1992 B.n389 B.n313 10.6151
R1993 B.n389 B.n388 10.6151
R1994 B.n388 B.n387 10.6151
R1995 B.n387 B.n315 10.6151
R1996 B.n381 B.n315 10.6151
R1997 B.n381 B.n380 10.6151
R1998 B.n380 B.n379 10.6151
R1999 B.n379 B.n317 10.6151
R2000 B.n373 B.n317 10.6151
R2001 B.n373 B.n372 10.6151
R2002 B.n372 B.n371 10.6151
R2003 B.n371 B.n319 10.6151
R2004 B.n365 B.n319 10.6151
R2005 B.n365 B.n364 10.6151
R2006 B.n364 B.n363 10.6151
R2007 B.n363 B.n321 10.6151
R2008 B.n357 B.n321 10.6151
R2009 B.n357 B.n356 10.6151
R2010 B.n356 B.n355 10.6151
R2011 B.n355 B.n323 10.6151
R2012 B.n349 B.n323 10.6151
R2013 B.n349 B.n348 10.6151
R2014 B.n348 B.n347 10.6151
R2015 B.n347 B.n325 10.6151
R2016 B.n341 B.n325 10.6151
R2017 B.n341 B.n340 10.6151
R2018 B.n340 B.n339 10.6151
R2019 B.n339 B.n327 10.6151
R2020 B.n333 B.n327 10.6151
R2021 B.n333 B.n332 10.6151
R2022 B.n332 B.n331 10.6151
R2023 B.n331 B.n257 10.6151
R2024 B.n583 B.n253 10.6151
R2025 B.n593 B.n253 10.6151
R2026 B.n594 B.n593 10.6151
R2027 B.n595 B.n594 10.6151
R2028 B.n595 B.n245 10.6151
R2029 B.n605 B.n245 10.6151
R2030 B.n606 B.n605 10.6151
R2031 B.n607 B.n606 10.6151
R2032 B.n607 B.n237 10.6151
R2033 B.n617 B.n237 10.6151
R2034 B.n618 B.n617 10.6151
R2035 B.n619 B.n618 10.6151
R2036 B.n619 B.n229 10.6151
R2037 B.n629 B.n229 10.6151
R2038 B.n630 B.n629 10.6151
R2039 B.n631 B.n630 10.6151
R2040 B.n631 B.n221 10.6151
R2041 B.n641 B.n221 10.6151
R2042 B.n642 B.n641 10.6151
R2043 B.n643 B.n642 10.6151
R2044 B.n643 B.n213 10.6151
R2045 B.n654 B.n213 10.6151
R2046 B.n655 B.n654 10.6151
R2047 B.n656 B.n655 10.6151
R2048 B.n656 B.n206 10.6151
R2049 B.n666 B.n206 10.6151
R2050 B.n667 B.n666 10.6151
R2051 B.n668 B.n667 10.6151
R2052 B.n668 B.n198 10.6151
R2053 B.n678 B.n198 10.6151
R2054 B.n679 B.n678 10.6151
R2055 B.n680 B.n679 10.6151
R2056 B.n680 B.n190 10.6151
R2057 B.n690 B.n190 10.6151
R2058 B.n691 B.n690 10.6151
R2059 B.n692 B.n691 10.6151
R2060 B.n692 B.n182 10.6151
R2061 B.n702 B.n182 10.6151
R2062 B.n703 B.n702 10.6151
R2063 B.n704 B.n703 10.6151
R2064 B.n704 B.n174 10.6151
R2065 B.n714 B.n174 10.6151
R2066 B.n715 B.n714 10.6151
R2067 B.n716 B.n715 10.6151
R2068 B.n716 B.n166 10.6151
R2069 B.n727 B.n166 10.6151
R2070 B.n728 B.n727 10.6151
R2071 B.n729 B.n728 10.6151
R2072 B.n729 B.n0 10.6151
R2073 B.n1151 B.n1 10.6151
R2074 B.n1151 B.n1150 10.6151
R2075 B.n1150 B.n1149 10.6151
R2076 B.n1149 B.n10 10.6151
R2077 B.n1143 B.n10 10.6151
R2078 B.n1143 B.n1142 10.6151
R2079 B.n1142 B.n1141 10.6151
R2080 B.n1141 B.n17 10.6151
R2081 B.n1135 B.n17 10.6151
R2082 B.n1135 B.n1134 10.6151
R2083 B.n1134 B.n1133 10.6151
R2084 B.n1133 B.n24 10.6151
R2085 B.n1127 B.n24 10.6151
R2086 B.n1127 B.n1126 10.6151
R2087 B.n1126 B.n1125 10.6151
R2088 B.n1125 B.n31 10.6151
R2089 B.n1119 B.n31 10.6151
R2090 B.n1119 B.n1118 10.6151
R2091 B.n1118 B.n1117 10.6151
R2092 B.n1117 B.n38 10.6151
R2093 B.n1111 B.n38 10.6151
R2094 B.n1111 B.n1110 10.6151
R2095 B.n1110 B.n1109 10.6151
R2096 B.n1109 B.n45 10.6151
R2097 B.n1103 B.n45 10.6151
R2098 B.n1103 B.n1102 10.6151
R2099 B.n1102 B.n1101 10.6151
R2100 B.n1101 B.n51 10.6151
R2101 B.n1095 B.n51 10.6151
R2102 B.n1095 B.n1094 10.6151
R2103 B.n1094 B.n1093 10.6151
R2104 B.n1093 B.n59 10.6151
R2105 B.n1087 B.n59 10.6151
R2106 B.n1087 B.n1086 10.6151
R2107 B.n1086 B.n1085 10.6151
R2108 B.n1085 B.n66 10.6151
R2109 B.n1079 B.n66 10.6151
R2110 B.n1079 B.n1078 10.6151
R2111 B.n1078 B.n1077 10.6151
R2112 B.n1077 B.n73 10.6151
R2113 B.n1071 B.n73 10.6151
R2114 B.n1071 B.n1070 10.6151
R2115 B.n1070 B.n1069 10.6151
R2116 B.n1069 B.n80 10.6151
R2117 B.n1063 B.n80 10.6151
R2118 B.n1063 B.n1062 10.6151
R2119 B.n1062 B.n1061 10.6151
R2120 B.n1061 B.n87 10.6151
R2121 B.n1055 B.n87 10.6151
R2122 B.t8 B.n243 9.96384
R2123 B.t12 B.n78 9.96384
R2124 B.n126 B.n122 9.36635
R2125 B.n917 B.n916 9.36635
R2126 B.n466 B.n465 9.36635
R2127 B.n443 B.n299 9.36635
R2128 B.t22 B.n223 3.32161
R2129 B.n658 B.t3 3.32161
R2130 B.t4 B.n196 3.32161
R2131 B.n700 B.t0 3.32161
R2132 B.t6 B.n168 3.32161
R2133 B.n1146 B.t23 3.32161
R2134 B.n1131 B.t5 3.32161
R2135 B.t21 B.n36 3.32161
R2136 B.n1105 B.t2 3.32161
R2137 B.n1090 B.t1 3.32161
R2138 B.n1157 B.n0 2.81026
R2139 B.n1157 B.n1 2.81026
R2140 B.n935 B.n126 1.24928
R2141 B.n918 B.n917 1.24928
R2142 B.n465 B.n464 1.24928
R2143 B.n447 B.n299 1.24928
R2144 VP.n19 VP.t0 241.964
R2145 VP.n48 VP.t1 210.553
R2146 VP.n56 VP.t8 210.553
R2147 VP.n5 VP.t5 210.553
R2148 VP.n73 VP.t9 210.553
R2149 VP.n81 VP.t3 210.553
R2150 VP.n45 VP.t7 210.553
R2151 VP.n37 VP.t6 210.553
R2152 VP.n16 VP.t4 210.553
R2153 VP.n20 VP.t2 210.553
R2154 VP.n48 VP.n47 185.279
R2155 VP.n82 VP.n81 185.279
R2156 VP.n46 VP.n45 185.279
R2157 VP.n22 VP.n21 161.3
R2158 VP.n23 VP.n18 161.3
R2159 VP.n25 VP.n24 161.3
R2160 VP.n26 VP.n17 161.3
R2161 VP.n28 VP.n27 161.3
R2162 VP.n30 VP.n29 161.3
R2163 VP.n31 VP.n15 161.3
R2164 VP.n33 VP.n32 161.3
R2165 VP.n34 VP.n14 161.3
R2166 VP.n36 VP.n35 161.3
R2167 VP.n38 VP.n13 161.3
R2168 VP.n40 VP.n39 161.3
R2169 VP.n41 VP.n12 161.3
R2170 VP.n43 VP.n42 161.3
R2171 VP.n44 VP.n11 161.3
R2172 VP.n80 VP.n0 161.3
R2173 VP.n79 VP.n78 161.3
R2174 VP.n77 VP.n1 161.3
R2175 VP.n76 VP.n75 161.3
R2176 VP.n74 VP.n2 161.3
R2177 VP.n72 VP.n71 161.3
R2178 VP.n70 VP.n3 161.3
R2179 VP.n69 VP.n68 161.3
R2180 VP.n67 VP.n4 161.3
R2181 VP.n66 VP.n65 161.3
R2182 VP.n64 VP.n63 161.3
R2183 VP.n62 VP.n6 161.3
R2184 VP.n61 VP.n60 161.3
R2185 VP.n59 VP.n7 161.3
R2186 VP.n58 VP.n57 161.3
R2187 VP.n55 VP.n8 161.3
R2188 VP.n54 VP.n53 161.3
R2189 VP.n52 VP.n9 161.3
R2190 VP.n51 VP.n50 161.3
R2191 VP.n49 VP.n10 161.3
R2192 VP.n20 VP.n19 64.109
R2193 VP.n54 VP.n9 56.5193
R2194 VP.n39 VP.n12 56.5193
R2195 VP.n75 VP.n1 56.5193
R2196 VP.n47 VP.n46 54.5156
R2197 VP.n62 VP.n61 46.321
R2198 VP.n68 VP.n67 46.321
R2199 VP.n32 VP.n31 46.321
R2200 VP.n26 VP.n25 46.321
R2201 VP.n61 VP.n7 34.6658
R2202 VP.n68 VP.n3 34.6658
R2203 VP.n32 VP.n14 34.6658
R2204 VP.n25 VP.n18 34.6658
R2205 VP.n50 VP.n49 24.4675
R2206 VP.n50 VP.n9 24.4675
R2207 VP.n55 VP.n54 24.4675
R2208 VP.n57 VP.n7 24.4675
R2209 VP.n63 VP.n62 24.4675
R2210 VP.n67 VP.n66 24.4675
R2211 VP.n72 VP.n3 24.4675
R2212 VP.n75 VP.n74 24.4675
R2213 VP.n79 VP.n1 24.4675
R2214 VP.n80 VP.n79 24.4675
R2215 VP.n43 VP.n12 24.4675
R2216 VP.n44 VP.n43 24.4675
R2217 VP.n36 VP.n14 24.4675
R2218 VP.n39 VP.n38 24.4675
R2219 VP.n27 VP.n26 24.4675
R2220 VP.n31 VP.n30 24.4675
R2221 VP.n21 VP.n18 24.4675
R2222 VP.n56 VP.n55 18.1061
R2223 VP.n74 VP.n73 18.1061
R2224 VP.n38 VP.n37 18.1061
R2225 VP.n22 VP.n19 12.6405
R2226 VP.n63 VP.n5 12.234
R2227 VP.n66 VP.n5 12.234
R2228 VP.n27 VP.n16 12.234
R2229 VP.n30 VP.n16 12.234
R2230 VP.n57 VP.n56 6.36192
R2231 VP.n73 VP.n72 6.36192
R2232 VP.n37 VP.n36 6.36192
R2233 VP.n21 VP.n20 6.36192
R2234 VP.n49 VP.n48 0.48984
R2235 VP.n81 VP.n80 0.48984
R2236 VP.n45 VP.n44 0.48984
R2237 VP.n23 VP.n22 0.189894
R2238 VP.n24 VP.n23 0.189894
R2239 VP.n24 VP.n17 0.189894
R2240 VP.n28 VP.n17 0.189894
R2241 VP.n29 VP.n28 0.189894
R2242 VP.n29 VP.n15 0.189894
R2243 VP.n33 VP.n15 0.189894
R2244 VP.n34 VP.n33 0.189894
R2245 VP.n35 VP.n34 0.189894
R2246 VP.n35 VP.n13 0.189894
R2247 VP.n40 VP.n13 0.189894
R2248 VP.n41 VP.n40 0.189894
R2249 VP.n42 VP.n41 0.189894
R2250 VP.n42 VP.n11 0.189894
R2251 VP.n46 VP.n11 0.189894
R2252 VP.n47 VP.n10 0.189894
R2253 VP.n51 VP.n10 0.189894
R2254 VP.n52 VP.n51 0.189894
R2255 VP.n53 VP.n52 0.189894
R2256 VP.n53 VP.n8 0.189894
R2257 VP.n58 VP.n8 0.189894
R2258 VP.n59 VP.n58 0.189894
R2259 VP.n60 VP.n59 0.189894
R2260 VP.n60 VP.n6 0.189894
R2261 VP.n64 VP.n6 0.189894
R2262 VP.n65 VP.n64 0.189894
R2263 VP.n65 VP.n4 0.189894
R2264 VP.n69 VP.n4 0.189894
R2265 VP.n70 VP.n69 0.189894
R2266 VP.n71 VP.n70 0.189894
R2267 VP.n71 VP.n2 0.189894
R2268 VP.n76 VP.n2 0.189894
R2269 VP.n77 VP.n76 0.189894
R2270 VP.n78 VP.n77 0.189894
R2271 VP.n78 VP.n0 0.189894
R2272 VP.n82 VP.n0 0.189894
R2273 VP VP.n82 0.0516364
R2274 VDD1.n1 VDD1.t9 64.4031
R2275 VDD1.n3 VDD1.t8 64.4028
R2276 VDD1.n5 VDD1.n4 62.729
R2277 VDD1.n1 VDD1.n0 61.2458
R2278 VDD1.n7 VDD1.n6 61.2456
R2279 VDD1.n3 VDD1.n2 61.2456
R2280 VDD1.n7 VDD1.n5 50.5095
R2281 VDD1 VDD1.n7 1.4811
R2282 VDD1.n6 VDD1.t3 1.10603
R2283 VDD1.n6 VDD1.t2 1.10603
R2284 VDD1.n0 VDD1.t7 1.10603
R2285 VDD1.n0 VDD1.t5 1.10603
R2286 VDD1.n4 VDD1.t0 1.10603
R2287 VDD1.n4 VDD1.t6 1.10603
R2288 VDD1.n2 VDD1.t1 1.10603
R2289 VDD1.n2 VDD1.t4 1.10603
R2290 VDD1 VDD1.n1 0.571621
R2291 VDD1.n5 VDD1.n3 0.458085
C0 VP VDD2 0.513961f
C1 VDD2 VTAIL 13.549701f
C2 VP VDD1 15.2121f
C3 VDD1 VTAIL 13.5049f
C4 VP VN 8.67949f
C5 VN VTAIL 15.017701f
C6 VP VTAIL 15.032201f
C7 VDD1 VDD2 1.81712f
C8 VN VDD2 14.855401f
C9 VN VDD1 0.152058f
C10 VDD2 B 7.58637f
C11 VDD1 B 7.579412f
C12 VTAIL B 10.08976f
C13 VN B 16.06142f
C14 VP B 14.396321f
C15 VDD1.t9 B 3.66606f
C16 VDD1.t7 B 0.313737f
C17 VDD1.t5 B 0.313737f
C18 VDD1.n0 B 2.85797f
C19 VDD1.n1 B 0.757766f
C20 VDD1.t8 B 3.66606f
C21 VDD1.t1 B 0.313737f
C22 VDD1.t4 B 0.313737f
C23 VDD1.n2 B 2.85797f
C24 VDD1.n3 B 0.750785f
C25 VDD1.t0 B 0.313737f
C26 VDD1.t6 B 0.313737f
C27 VDD1.n4 B 2.8685f
C28 VDD1.n5 B 2.74965f
C29 VDD1.t3 B 0.313737f
C30 VDD1.t2 B 0.313737f
C31 VDD1.n6 B 2.85796f
C32 VDD1.n7 B 3.01083f
C33 VP.n0 B 0.024322f
C34 VP.t3 B 2.45603f
C35 VP.n1 B 0.030762f
C36 VP.n2 B 0.024322f
C37 VP.t9 B 2.45603f
C38 VP.n3 B 0.049147f
C39 VP.n4 B 0.024322f
C40 VP.t5 B 2.45603f
C41 VP.n5 B 0.856582f
C42 VP.n6 B 0.024322f
C43 VP.n7 B 0.049147f
C44 VP.n8 B 0.024322f
C45 VP.t8 B 2.45603f
C46 VP.n9 B 0.030762f
C47 VP.n10 B 0.024322f
C48 VP.t1 B 2.45603f
C49 VP.n11 B 0.024322f
C50 VP.t7 B 2.45603f
C51 VP.n12 B 0.030762f
C52 VP.n13 B 0.024322f
C53 VP.t6 B 2.45603f
C54 VP.n14 B 0.049147f
C55 VP.n15 B 0.024322f
C56 VP.t4 B 2.45603f
C57 VP.n16 B 0.856582f
C58 VP.n17 B 0.024322f
C59 VP.n18 B 0.049147f
C60 VP.t0 B 2.58358f
C61 VP.n19 B 0.9201f
C62 VP.t2 B 2.45603f
C63 VP.n20 B 0.910985f
C64 VP.n21 B 0.028769f
C65 VP.n22 B 0.182983f
C66 VP.n23 B 0.024322f
C67 VP.n24 B 0.024322f
C68 VP.n25 B 0.020811f
C69 VP.n26 B 0.046384f
C70 VP.n27 B 0.034141f
C71 VP.n28 B 0.024322f
C72 VP.n29 B 0.024322f
C73 VP.n30 B 0.034141f
C74 VP.n31 B 0.046384f
C75 VP.n32 B 0.020811f
C76 VP.n33 B 0.024322f
C77 VP.n34 B 0.024322f
C78 VP.n35 B 0.024322f
C79 VP.n36 B 0.028769f
C80 VP.n37 B 0.856582f
C81 VP.n38 B 0.039512f
C82 VP.n39 B 0.04025f
C83 VP.n40 B 0.024322f
C84 VP.n41 B 0.024322f
C85 VP.n42 B 0.024322f
C86 VP.n43 B 0.04533f
C87 VP.n44 B 0.023398f
C88 VP.n45 B 0.917868f
C89 VP.n46 B 1.51092f
C90 VP.n47 B 1.52696f
C91 VP.n48 B 0.917868f
C92 VP.n49 B 0.023398f
C93 VP.n50 B 0.04533f
C94 VP.n51 B 0.024322f
C95 VP.n52 B 0.024322f
C96 VP.n53 B 0.024322f
C97 VP.n54 B 0.04025f
C98 VP.n55 B 0.039512f
C99 VP.n56 B 0.856582f
C100 VP.n57 B 0.028769f
C101 VP.n58 B 0.024322f
C102 VP.n59 B 0.024322f
C103 VP.n60 B 0.024322f
C104 VP.n61 B 0.020811f
C105 VP.n62 B 0.046384f
C106 VP.n63 B 0.034141f
C107 VP.n64 B 0.024322f
C108 VP.n65 B 0.024322f
C109 VP.n66 B 0.034141f
C110 VP.n67 B 0.046384f
C111 VP.n68 B 0.020811f
C112 VP.n69 B 0.024322f
C113 VP.n70 B 0.024322f
C114 VP.n71 B 0.024322f
C115 VP.n72 B 0.028769f
C116 VP.n73 B 0.856582f
C117 VP.n74 B 0.039512f
C118 VP.n75 B 0.04025f
C119 VP.n76 B 0.024322f
C120 VP.n77 B 0.024322f
C121 VP.n78 B 0.024322f
C122 VP.n79 B 0.04533f
C123 VP.n80 B 0.023398f
C124 VP.n81 B 0.917868f
C125 VP.n82 B 0.027959f
C126 VTAIL.t13 B 0.332101f
C127 VTAIL.t9 B 0.332101f
C128 VTAIL.n0 B 2.95416f
C129 VTAIL.n1 B 0.467487f
C130 VTAIL.t6 B 3.7745f
C131 VTAIL.n2 B 0.587264f
C132 VTAIL.t4 B 0.332101f
C133 VTAIL.t0 B 0.332101f
C134 VTAIL.n3 B 2.95416f
C135 VTAIL.n4 B 0.543912f
C136 VTAIL.t18 B 0.332101f
C137 VTAIL.t3 B 0.332101f
C138 VTAIL.n5 B 2.95416f
C139 VTAIL.n6 B 2.18517f
C140 VTAIL.t11 B 0.332101f
C141 VTAIL.t12 B 0.332101f
C142 VTAIL.n7 B 2.95416f
C143 VTAIL.n8 B 2.18517f
C144 VTAIL.t15 B 0.332101f
C145 VTAIL.t7 B 0.332101f
C146 VTAIL.n9 B 2.95416f
C147 VTAIL.n10 B 0.543908f
C148 VTAIL.t10 B 3.7745f
C149 VTAIL.n11 B 0.587259f
C150 VTAIL.t19 B 0.332101f
C151 VTAIL.t5 B 0.332101f
C152 VTAIL.n12 B 2.95416f
C153 VTAIL.n13 B 0.501866f
C154 VTAIL.t17 B 0.332101f
C155 VTAIL.t2 B 0.332101f
C156 VTAIL.n14 B 2.95416f
C157 VTAIL.n15 B 0.543908f
C158 VTAIL.t1 B 3.7745f
C159 VTAIL.n16 B 2.11544f
C160 VTAIL.t14 B 3.7745f
C161 VTAIL.n17 B 2.11544f
C162 VTAIL.t8 B 0.332101f
C163 VTAIL.t16 B 0.332101f
C164 VTAIL.n18 B 2.95416f
C165 VTAIL.n19 B 0.423165f
C166 VDD2.t2 B 3.63812f
C167 VDD2.t8 B 0.311346f
C168 VDD2.t7 B 0.311346f
C169 VDD2.n0 B 2.83618f
C170 VDD2.n1 B 0.745063f
C171 VDD2.t0 B 0.311346f
C172 VDD2.t3 B 0.311346f
C173 VDD2.n2 B 2.84664f
C174 VDD2.n3 B 2.62872f
C175 VDD2.t6 B 3.62549f
C176 VDD2.n4 B 2.96146f
C177 VDD2.t1 B 0.311346f
C178 VDD2.t4 B 0.311346f
C179 VDD2.n5 B 2.83619f
C180 VDD2.n6 B 0.36821f
C181 VDD2.t9 B 0.311346f
C182 VDD2.t5 B 0.311346f
C183 VDD2.n7 B 2.8466f
C184 VN.n0 B 0.024113f
C185 VN.t2 B 2.43495f
C186 VN.n1 B 0.030498f
C187 VN.n2 B 0.024113f
C188 VN.t0 B 2.43495f
C189 VN.n3 B 0.048726f
C190 VN.n4 B 0.024113f
C191 VN.t8 B 2.43495f
C192 VN.n5 B 0.84923f
C193 VN.n6 B 0.024113f
C194 VN.n7 B 0.048726f
C195 VN.t3 B 2.5614f
C196 VN.n8 B 0.912202f
C197 VN.t7 B 2.43495f
C198 VN.n9 B 0.903165f
C199 VN.n10 B 0.028522f
C200 VN.n11 B 0.181412f
C201 VN.n12 B 0.024113f
C202 VN.n13 B 0.024113f
C203 VN.n14 B 0.020632f
C204 VN.n15 B 0.045986f
C205 VN.n16 B 0.033847f
C206 VN.n17 B 0.024113f
C207 VN.n18 B 0.024113f
C208 VN.n19 B 0.033847f
C209 VN.n20 B 0.045986f
C210 VN.n21 B 0.020632f
C211 VN.n22 B 0.024113f
C212 VN.n23 B 0.024113f
C213 VN.n24 B 0.024113f
C214 VN.n25 B 0.028522f
C215 VN.n26 B 0.84923f
C216 VN.n27 B 0.039173f
C217 VN.n28 B 0.039905f
C218 VN.n29 B 0.024113f
C219 VN.n30 B 0.024113f
C220 VN.n31 B 0.024113f
C221 VN.n32 B 0.044941f
C222 VN.n33 B 0.023197f
C223 VN.n34 B 0.909989f
C224 VN.n35 B 0.027719f
C225 VN.n36 B 0.024113f
C226 VN.t5 B 2.43495f
C227 VN.n37 B 0.030498f
C228 VN.n38 B 0.024113f
C229 VN.t4 B 2.43495f
C230 VN.n39 B 0.048726f
C231 VN.n40 B 0.024113f
C232 VN.t1 B 2.43495f
C233 VN.n41 B 0.84923f
C234 VN.n42 B 0.024113f
C235 VN.n43 B 0.048726f
C236 VN.t6 B 2.5614f
C237 VN.n44 B 0.912202f
C238 VN.t9 B 2.43495f
C239 VN.n45 B 0.903165f
C240 VN.n46 B 0.028522f
C241 VN.n47 B 0.181412f
C242 VN.n48 B 0.024113f
C243 VN.n49 B 0.024113f
C244 VN.n50 B 0.020632f
C245 VN.n51 B 0.045986f
C246 VN.n52 B 0.033847f
C247 VN.n53 B 0.024113f
C248 VN.n54 B 0.024113f
C249 VN.n55 B 0.033847f
C250 VN.n56 B 0.045986f
C251 VN.n57 B 0.020632f
C252 VN.n58 B 0.024113f
C253 VN.n59 B 0.024113f
C254 VN.n60 B 0.024113f
C255 VN.n61 B 0.028522f
C256 VN.n62 B 0.84923f
C257 VN.n63 B 0.039173f
C258 VN.n64 B 0.039905f
C259 VN.n65 B 0.024113f
C260 VN.n66 B 0.024113f
C261 VN.n67 B 0.024113f
C262 VN.n68 B 0.044941f
C263 VN.n69 B 0.023197f
C264 VN.n70 B 0.909989f
C265 VN.n71 B 1.51356f
.ends

