* NGSPICE file created from diff_pair_sample_1429.ext - technology: sky130A

.subckt diff_pair_sample_1429 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=1.65 ps=10.33 w=10 l=1.48
X1 VDD1.t7 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=3.9 ps=20.78 w=10 l=1.48
X2 VDD1.t6 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=3.9 ps=20.78 w=10 l=1.48
X3 VTAIL.t5 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X4 VDD2.t7 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X5 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=1.48
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=1.48
X7 VTAIL.t13 VN.t2 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=1.65 ps=10.33 w=10 l=1.48
X8 VTAIL.t2 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=1.65 ps=10.33 w=10 l=1.48
X9 VDD2.t4 VN.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=3.9 ps=20.78 w=10 l=1.48
X10 VDD2.t1 VN.t4 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=1.48
X12 VDD1.t3 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=0 ps=0 w=10 l=1.48
X14 VTAIL.t10 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X15 VDD1.t2 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X16 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
X17 VTAIL.t7 VP.t7 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.9 pd=20.78 as=1.65 ps=10.33 w=10 l=1.48
X18 VDD2.t0 VN.t6 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=3.9 ps=20.78 w=10 l=1.48
X19 VTAIL.t8 VN.t7 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.65 pd=10.33 as=1.65 ps=10.33 w=10 l=1.48
R0 VN.n5 VN.t2 196.924
R1 VN.n24 VN.t3 196.924
R2 VN.n18 VN.n17 175.317
R3 VN.n37 VN.n36 175.317
R4 VN.n4 VN.t1 162.839
R5 VN.n10 VN.t7 162.839
R6 VN.n17 VN.t6 162.839
R7 VN.n23 VN.t5 162.839
R8 VN.n29 VN.t4 162.839
R9 VN.n36 VN.t0 162.839
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n28 VN.n21 161.3
R15 VN.n27 VN.n26 161.3
R16 VN.n25 VN.n22 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n15 VN.n1 56.5617
R25 VN.n34 VN.n20 56.5617
R26 VN.n5 VN.n4 46.7161
R27 VN.n24 VN.n23 46.7161
R28 VN VN.n37 44.4494
R29 VN.n8 VN.n3 40.577
R30 VN.n9 VN.n8 40.577
R31 VN.n27 VN.n22 40.577
R32 VN.n28 VN.n27 40.577
R33 VN.n11 VN.n1 24.5923
R34 VN.n16 VN.n15 24.5923
R35 VN.n30 VN.n20 24.5923
R36 VN.n35 VN.n34 24.5923
R37 VN.n4 VN.n3 19.9199
R38 VN.n10 VN.n9 19.9199
R39 VN.n23 VN.n22 19.9199
R40 VN.n29 VN.n28 19.9199
R41 VN.n25 VN.n24 17.7081
R42 VN.n6 VN.n5 17.7081
R43 VN.n17 VN.n16 10.575
R44 VN.n36 VN.n35 10.575
R45 VN.n11 VN.n10 4.67295
R46 VN.n30 VN.n29 4.67295
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n26 VN.n21 0.189894
R53 VN.n26 VN.n25 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VDD2.n2 VDD2.n1 64.1407
R63 VDD2.n2 VDD2.n0 64.1407
R64 VDD2 VDD2.n5 64.1379
R65 VDD2.n4 VDD2.n3 63.4161
R66 VDD2.n4 VDD2.n2 39.3575
R67 VDD2.n5 VDD2.t2 1.9805
R68 VDD2.n5 VDD2.t4 1.9805
R69 VDD2.n3 VDD2.t6 1.9805
R70 VDD2.n3 VDD2.t1 1.9805
R71 VDD2.n1 VDD2.t5 1.9805
R72 VDD2.n1 VDD2.t0 1.9805
R73 VDD2.n0 VDD2.t3 1.9805
R74 VDD2.n0 VDD2.t7 1.9805
R75 VDD2 VDD2.n4 0.838862
R76 VTAIL.n434 VTAIL.n386 289.615
R77 VTAIL.n50 VTAIL.n2 289.615
R78 VTAIL.n104 VTAIL.n56 289.615
R79 VTAIL.n160 VTAIL.n112 289.615
R80 VTAIL.n380 VTAIL.n332 289.615
R81 VTAIL.n324 VTAIL.n276 289.615
R82 VTAIL.n270 VTAIL.n222 289.615
R83 VTAIL.n214 VTAIL.n166 289.615
R84 VTAIL.n402 VTAIL.n401 185
R85 VTAIL.n407 VTAIL.n406 185
R86 VTAIL.n409 VTAIL.n408 185
R87 VTAIL.n398 VTAIL.n397 185
R88 VTAIL.n415 VTAIL.n414 185
R89 VTAIL.n417 VTAIL.n416 185
R90 VTAIL.n394 VTAIL.n393 185
R91 VTAIL.n424 VTAIL.n423 185
R92 VTAIL.n425 VTAIL.n392 185
R93 VTAIL.n427 VTAIL.n426 185
R94 VTAIL.n390 VTAIL.n389 185
R95 VTAIL.n433 VTAIL.n432 185
R96 VTAIL.n435 VTAIL.n434 185
R97 VTAIL.n18 VTAIL.n17 185
R98 VTAIL.n23 VTAIL.n22 185
R99 VTAIL.n25 VTAIL.n24 185
R100 VTAIL.n14 VTAIL.n13 185
R101 VTAIL.n31 VTAIL.n30 185
R102 VTAIL.n33 VTAIL.n32 185
R103 VTAIL.n10 VTAIL.n9 185
R104 VTAIL.n40 VTAIL.n39 185
R105 VTAIL.n41 VTAIL.n8 185
R106 VTAIL.n43 VTAIL.n42 185
R107 VTAIL.n6 VTAIL.n5 185
R108 VTAIL.n49 VTAIL.n48 185
R109 VTAIL.n51 VTAIL.n50 185
R110 VTAIL.n72 VTAIL.n71 185
R111 VTAIL.n77 VTAIL.n76 185
R112 VTAIL.n79 VTAIL.n78 185
R113 VTAIL.n68 VTAIL.n67 185
R114 VTAIL.n85 VTAIL.n84 185
R115 VTAIL.n87 VTAIL.n86 185
R116 VTAIL.n64 VTAIL.n63 185
R117 VTAIL.n94 VTAIL.n93 185
R118 VTAIL.n95 VTAIL.n62 185
R119 VTAIL.n97 VTAIL.n96 185
R120 VTAIL.n60 VTAIL.n59 185
R121 VTAIL.n103 VTAIL.n102 185
R122 VTAIL.n105 VTAIL.n104 185
R123 VTAIL.n128 VTAIL.n127 185
R124 VTAIL.n133 VTAIL.n132 185
R125 VTAIL.n135 VTAIL.n134 185
R126 VTAIL.n124 VTAIL.n123 185
R127 VTAIL.n141 VTAIL.n140 185
R128 VTAIL.n143 VTAIL.n142 185
R129 VTAIL.n120 VTAIL.n119 185
R130 VTAIL.n150 VTAIL.n149 185
R131 VTAIL.n151 VTAIL.n118 185
R132 VTAIL.n153 VTAIL.n152 185
R133 VTAIL.n116 VTAIL.n115 185
R134 VTAIL.n159 VTAIL.n158 185
R135 VTAIL.n161 VTAIL.n160 185
R136 VTAIL.n381 VTAIL.n380 185
R137 VTAIL.n379 VTAIL.n378 185
R138 VTAIL.n336 VTAIL.n335 185
R139 VTAIL.n373 VTAIL.n372 185
R140 VTAIL.n371 VTAIL.n338 185
R141 VTAIL.n370 VTAIL.n369 185
R142 VTAIL.n341 VTAIL.n339 185
R143 VTAIL.n364 VTAIL.n363 185
R144 VTAIL.n362 VTAIL.n361 185
R145 VTAIL.n345 VTAIL.n344 185
R146 VTAIL.n356 VTAIL.n355 185
R147 VTAIL.n354 VTAIL.n353 185
R148 VTAIL.n349 VTAIL.n348 185
R149 VTAIL.n325 VTAIL.n324 185
R150 VTAIL.n323 VTAIL.n322 185
R151 VTAIL.n280 VTAIL.n279 185
R152 VTAIL.n317 VTAIL.n316 185
R153 VTAIL.n315 VTAIL.n282 185
R154 VTAIL.n314 VTAIL.n313 185
R155 VTAIL.n285 VTAIL.n283 185
R156 VTAIL.n308 VTAIL.n307 185
R157 VTAIL.n306 VTAIL.n305 185
R158 VTAIL.n289 VTAIL.n288 185
R159 VTAIL.n300 VTAIL.n299 185
R160 VTAIL.n298 VTAIL.n297 185
R161 VTAIL.n293 VTAIL.n292 185
R162 VTAIL.n271 VTAIL.n270 185
R163 VTAIL.n269 VTAIL.n268 185
R164 VTAIL.n226 VTAIL.n225 185
R165 VTAIL.n263 VTAIL.n262 185
R166 VTAIL.n261 VTAIL.n228 185
R167 VTAIL.n260 VTAIL.n259 185
R168 VTAIL.n231 VTAIL.n229 185
R169 VTAIL.n254 VTAIL.n253 185
R170 VTAIL.n252 VTAIL.n251 185
R171 VTAIL.n235 VTAIL.n234 185
R172 VTAIL.n246 VTAIL.n245 185
R173 VTAIL.n244 VTAIL.n243 185
R174 VTAIL.n239 VTAIL.n238 185
R175 VTAIL.n215 VTAIL.n214 185
R176 VTAIL.n213 VTAIL.n212 185
R177 VTAIL.n170 VTAIL.n169 185
R178 VTAIL.n207 VTAIL.n206 185
R179 VTAIL.n205 VTAIL.n172 185
R180 VTAIL.n204 VTAIL.n203 185
R181 VTAIL.n175 VTAIL.n173 185
R182 VTAIL.n198 VTAIL.n197 185
R183 VTAIL.n196 VTAIL.n195 185
R184 VTAIL.n179 VTAIL.n178 185
R185 VTAIL.n190 VTAIL.n189 185
R186 VTAIL.n188 VTAIL.n187 185
R187 VTAIL.n183 VTAIL.n182 185
R188 VTAIL.n403 VTAIL.t9 149.524
R189 VTAIL.n19 VTAIL.t13 149.524
R190 VTAIL.n73 VTAIL.t3 149.524
R191 VTAIL.n129 VTAIL.t2 149.524
R192 VTAIL.n350 VTAIL.t6 149.524
R193 VTAIL.n294 VTAIL.t7 149.524
R194 VTAIL.n240 VTAIL.t12 149.524
R195 VTAIL.n184 VTAIL.t15 149.524
R196 VTAIL.n407 VTAIL.n401 104.615
R197 VTAIL.n408 VTAIL.n407 104.615
R198 VTAIL.n408 VTAIL.n397 104.615
R199 VTAIL.n415 VTAIL.n397 104.615
R200 VTAIL.n416 VTAIL.n415 104.615
R201 VTAIL.n416 VTAIL.n393 104.615
R202 VTAIL.n424 VTAIL.n393 104.615
R203 VTAIL.n425 VTAIL.n424 104.615
R204 VTAIL.n426 VTAIL.n425 104.615
R205 VTAIL.n426 VTAIL.n389 104.615
R206 VTAIL.n433 VTAIL.n389 104.615
R207 VTAIL.n434 VTAIL.n433 104.615
R208 VTAIL.n23 VTAIL.n17 104.615
R209 VTAIL.n24 VTAIL.n23 104.615
R210 VTAIL.n24 VTAIL.n13 104.615
R211 VTAIL.n31 VTAIL.n13 104.615
R212 VTAIL.n32 VTAIL.n31 104.615
R213 VTAIL.n32 VTAIL.n9 104.615
R214 VTAIL.n40 VTAIL.n9 104.615
R215 VTAIL.n41 VTAIL.n40 104.615
R216 VTAIL.n42 VTAIL.n41 104.615
R217 VTAIL.n42 VTAIL.n5 104.615
R218 VTAIL.n49 VTAIL.n5 104.615
R219 VTAIL.n50 VTAIL.n49 104.615
R220 VTAIL.n77 VTAIL.n71 104.615
R221 VTAIL.n78 VTAIL.n77 104.615
R222 VTAIL.n78 VTAIL.n67 104.615
R223 VTAIL.n85 VTAIL.n67 104.615
R224 VTAIL.n86 VTAIL.n85 104.615
R225 VTAIL.n86 VTAIL.n63 104.615
R226 VTAIL.n94 VTAIL.n63 104.615
R227 VTAIL.n95 VTAIL.n94 104.615
R228 VTAIL.n96 VTAIL.n95 104.615
R229 VTAIL.n96 VTAIL.n59 104.615
R230 VTAIL.n103 VTAIL.n59 104.615
R231 VTAIL.n104 VTAIL.n103 104.615
R232 VTAIL.n133 VTAIL.n127 104.615
R233 VTAIL.n134 VTAIL.n133 104.615
R234 VTAIL.n134 VTAIL.n123 104.615
R235 VTAIL.n141 VTAIL.n123 104.615
R236 VTAIL.n142 VTAIL.n141 104.615
R237 VTAIL.n142 VTAIL.n119 104.615
R238 VTAIL.n150 VTAIL.n119 104.615
R239 VTAIL.n151 VTAIL.n150 104.615
R240 VTAIL.n152 VTAIL.n151 104.615
R241 VTAIL.n152 VTAIL.n115 104.615
R242 VTAIL.n159 VTAIL.n115 104.615
R243 VTAIL.n160 VTAIL.n159 104.615
R244 VTAIL.n380 VTAIL.n379 104.615
R245 VTAIL.n379 VTAIL.n335 104.615
R246 VTAIL.n372 VTAIL.n335 104.615
R247 VTAIL.n372 VTAIL.n371 104.615
R248 VTAIL.n371 VTAIL.n370 104.615
R249 VTAIL.n370 VTAIL.n339 104.615
R250 VTAIL.n363 VTAIL.n339 104.615
R251 VTAIL.n363 VTAIL.n362 104.615
R252 VTAIL.n362 VTAIL.n344 104.615
R253 VTAIL.n355 VTAIL.n344 104.615
R254 VTAIL.n355 VTAIL.n354 104.615
R255 VTAIL.n354 VTAIL.n348 104.615
R256 VTAIL.n324 VTAIL.n323 104.615
R257 VTAIL.n323 VTAIL.n279 104.615
R258 VTAIL.n316 VTAIL.n279 104.615
R259 VTAIL.n316 VTAIL.n315 104.615
R260 VTAIL.n315 VTAIL.n314 104.615
R261 VTAIL.n314 VTAIL.n283 104.615
R262 VTAIL.n307 VTAIL.n283 104.615
R263 VTAIL.n307 VTAIL.n306 104.615
R264 VTAIL.n306 VTAIL.n288 104.615
R265 VTAIL.n299 VTAIL.n288 104.615
R266 VTAIL.n299 VTAIL.n298 104.615
R267 VTAIL.n298 VTAIL.n292 104.615
R268 VTAIL.n270 VTAIL.n269 104.615
R269 VTAIL.n269 VTAIL.n225 104.615
R270 VTAIL.n262 VTAIL.n225 104.615
R271 VTAIL.n262 VTAIL.n261 104.615
R272 VTAIL.n261 VTAIL.n260 104.615
R273 VTAIL.n260 VTAIL.n229 104.615
R274 VTAIL.n253 VTAIL.n229 104.615
R275 VTAIL.n253 VTAIL.n252 104.615
R276 VTAIL.n252 VTAIL.n234 104.615
R277 VTAIL.n245 VTAIL.n234 104.615
R278 VTAIL.n245 VTAIL.n244 104.615
R279 VTAIL.n244 VTAIL.n238 104.615
R280 VTAIL.n214 VTAIL.n213 104.615
R281 VTAIL.n213 VTAIL.n169 104.615
R282 VTAIL.n206 VTAIL.n169 104.615
R283 VTAIL.n206 VTAIL.n205 104.615
R284 VTAIL.n205 VTAIL.n204 104.615
R285 VTAIL.n204 VTAIL.n173 104.615
R286 VTAIL.n197 VTAIL.n173 104.615
R287 VTAIL.n197 VTAIL.n196 104.615
R288 VTAIL.n196 VTAIL.n178 104.615
R289 VTAIL.n189 VTAIL.n178 104.615
R290 VTAIL.n189 VTAIL.n188 104.615
R291 VTAIL.n188 VTAIL.n182 104.615
R292 VTAIL.t9 VTAIL.n401 52.3082
R293 VTAIL.t13 VTAIL.n17 52.3082
R294 VTAIL.t3 VTAIL.n71 52.3082
R295 VTAIL.t2 VTAIL.n127 52.3082
R296 VTAIL.t6 VTAIL.n348 52.3082
R297 VTAIL.t7 VTAIL.n292 52.3082
R298 VTAIL.t12 VTAIL.n238 52.3082
R299 VTAIL.t15 VTAIL.n182 52.3082
R300 VTAIL.n331 VTAIL.n330 46.7373
R301 VTAIL.n221 VTAIL.n220 46.7373
R302 VTAIL.n1 VTAIL.n0 46.7371
R303 VTAIL.n111 VTAIL.n110 46.7371
R304 VTAIL.n439 VTAIL.n438 32.9611
R305 VTAIL.n55 VTAIL.n54 32.9611
R306 VTAIL.n109 VTAIL.n108 32.9611
R307 VTAIL.n165 VTAIL.n164 32.9611
R308 VTAIL.n385 VTAIL.n384 32.9611
R309 VTAIL.n329 VTAIL.n328 32.9611
R310 VTAIL.n275 VTAIL.n274 32.9611
R311 VTAIL.n219 VTAIL.n218 32.9611
R312 VTAIL.n439 VTAIL.n385 22.5479
R313 VTAIL.n219 VTAIL.n165 22.5479
R314 VTAIL.n427 VTAIL.n392 13.1884
R315 VTAIL.n43 VTAIL.n8 13.1884
R316 VTAIL.n97 VTAIL.n62 13.1884
R317 VTAIL.n153 VTAIL.n118 13.1884
R318 VTAIL.n373 VTAIL.n338 13.1884
R319 VTAIL.n317 VTAIL.n282 13.1884
R320 VTAIL.n263 VTAIL.n228 13.1884
R321 VTAIL.n207 VTAIL.n172 13.1884
R322 VTAIL.n423 VTAIL.n422 12.8005
R323 VTAIL.n428 VTAIL.n390 12.8005
R324 VTAIL.n39 VTAIL.n38 12.8005
R325 VTAIL.n44 VTAIL.n6 12.8005
R326 VTAIL.n93 VTAIL.n92 12.8005
R327 VTAIL.n98 VTAIL.n60 12.8005
R328 VTAIL.n149 VTAIL.n148 12.8005
R329 VTAIL.n154 VTAIL.n116 12.8005
R330 VTAIL.n374 VTAIL.n336 12.8005
R331 VTAIL.n369 VTAIL.n340 12.8005
R332 VTAIL.n318 VTAIL.n280 12.8005
R333 VTAIL.n313 VTAIL.n284 12.8005
R334 VTAIL.n264 VTAIL.n226 12.8005
R335 VTAIL.n259 VTAIL.n230 12.8005
R336 VTAIL.n208 VTAIL.n170 12.8005
R337 VTAIL.n203 VTAIL.n174 12.8005
R338 VTAIL.n421 VTAIL.n394 12.0247
R339 VTAIL.n432 VTAIL.n431 12.0247
R340 VTAIL.n37 VTAIL.n10 12.0247
R341 VTAIL.n48 VTAIL.n47 12.0247
R342 VTAIL.n91 VTAIL.n64 12.0247
R343 VTAIL.n102 VTAIL.n101 12.0247
R344 VTAIL.n147 VTAIL.n120 12.0247
R345 VTAIL.n158 VTAIL.n157 12.0247
R346 VTAIL.n378 VTAIL.n377 12.0247
R347 VTAIL.n368 VTAIL.n341 12.0247
R348 VTAIL.n322 VTAIL.n321 12.0247
R349 VTAIL.n312 VTAIL.n285 12.0247
R350 VTAIL.n268 VTAIL.n267 12.0247
R351 VTAIL.n258 VTAIL.n231 12.0247
R352 VTAIL.n212 VTAIL.n211 12.0247
R353 VTAIL.n202 VTAIL.n175 12.0247
R354 VTAIL.n418 VTAIL.n417 11.249
R355 VTAIL.n435 VTAIL.n388 11.249
R356 VTAIL.n34 VTAIL.n33 11.249
R357 VTAIL.n51 VTAIL.n4 11.249
R358 VTAIL.n88 VTAIL.n87 11.249
R359 VTAIL.n105 VTAIL.n58 11.249
R360 VTAIL.n144 VTAIL.n143 11.249
R361 VTAIL.n161 VTAIL.n114 11.249
R362 VTAIL.n381 VTAIL.n334 11.249
R363 VTAIL.n365 VTAIL.n364 11.249
R364 VTAIL.n325 VTAIL.n278 11.249
R365 VTAIL.n309 VTAIL.n308 11.249
R366 VTAIL.n271 VTAIL.n224 11.249
R367 VTAIL.n255 VTAIL.n254 11.249
R368 VTAIL.n215 VTAIL.n168 11.249
R369 VTAIL.n199 VTAIL.n198 11.249
R370 VTAIL.n414 VTAIL.n396 10.4732
R371 VTAIL.n436 VTAIL.n386 10.4732
R372 VTAIL.n30 VTAIL.n12 10.4732
R373 VTAIL.n52 VTAIL.n2 10.4732
R374 VTAIL.n84 VTAIL.n66 10.4732
R375 VTAIL.n106 VTAIL.n56 10.4732
R376 VTAIL.n140 VTAIL.n122 10.4732
R377 VTAIL.n162 VTAIL.n112 10.4732
R378 VTAIL.n382 VTAIL.n332 10.4732
R379 VTAIL.n361 VTAIL.n343 10.4732
R380 VTAIL.n326 VTAIL.n276 10.4732
R381 VTAIL.n305 VTAIL.n287 10.4732
R382 VTAIL.n272 VTAIL.n222 10.4732
R383 VTAIL.n251 VTAIL.n233 10.4732
R384 VTAIL.n216 VTAIL.n166 10.4732
R385 VTAIL.n195 VTAIL.n177 10.4732
R386 VTAIL.n403 VTAIL.n402 10.2747
R387 VTAIL.n19 VTAIL.n18 10.2747
R388 VTAIL.n73 VTAIL.n72 10.2747
R389 VTAIL.n129 VTAIL.n128 10.2747
R390 VTAIL.n350 VTAIL.n349 10.2747
R391 VTAIL.n294 VTAIL.n293 10.2747
R392 VTAIL.n240 VTAIL.n239 10.2747
R393 VTAIL.n184 VTAIL.n183 10.2747
R394 VTAIL.n413 VTAIL.n398 9.69747
R395 VTAIL.n29 VTAIL.n14 9.69747
R396 VTAIL.n83 VTAIL.n68 9.69747
R397 VTAIL.n139 VTAIL.n124 9.69747
R398 VTAIL.n360 VTAIL.n345 9.69747
R399 VTAIL.n304 VTAIL.n289 9.69747
R400 VTAIL.n250 VTAIL.n235 9.69747
R401 VTAIL.n194 VTAIL.n179 9.69747
R402 VTAIL.n438 VTAIL.n437 9.45567
R403 VTAIL.n54 VTAIL.n53 9.45567
R404 VTAIL.n108 VTAIL.n107 9.45567
R405 VTAIL.n164 VTAIL.n163 9.45567
R406 VTAIL.n384 VTAIL.n383 9.45567
R407 VTAIL.n328 VTAIL.n327 9.45567
R408 VTAIL.n274 VTAIL.n273 9.45567
R409 VTAIL.n218 VTAIL.n217 9.45567
R410 VTAIL.n437 VTAIL.n436 9.3005
R411 VTAIL.n388 VTAIL.n387 9.3005
R412 VTAIL.n431 VTAIL.n430 9.3005
R413 VTAIL.n429 VTAIL.n428 9.3005
R414 VTAIL.n405 VTAIL.n404 9.3005
R415 VTAIL.n400 VTAIL.n399 9.3005
R416 VTAIL.n411 VTAIL.n410 9.3005
R417 VTAIL.n413 VTAIL.n412 9.3005
R418 VTAIL.n396 VTAIL.n395 9.3005
R419 VTAIL.n419 VTAIL.n418 9.3005
R420 VTAIL.n421 VTAIL.n420 9.3005
R421 VTAIL.n422 VTAIL.n391 9.3005
R422 VTAIL.n53 VTAIL.n52 9.3005
R423 VTAIL.n4 VTAIL.n3 9.3005
R424 VTAIL.n47 VTAIL.n46 9.3005
R425 VTAIL.n45 VTAIL.n44 9.3005
R426 VTAIL.n21 VTAIL.n20 9.3005
R427 VTAIL.n16 VTAIL.n15 9.3005
R428 VTAIL.n27 VTAIL.n26 9.3005
R429 VTAIL.n29 VTAIL.n28 9.3005
R430 VTAIL.n12 VTAIL.n11 9.3005
R431 VTAIL.n35 VTAIL.n34 9.3005
R432 VTAIL.n37 VTAIL.n36 9.3005
R433 VTAIL.n38 VTAIL.n7 9.3005
R434 VTAIL.n107 VTAIL.n106 9.3005
R435 VTAIL.n58 VTAIL.n57 9.3005
R436 VTAIL.n101 VTAIL.n100 9.3005
R437 VTAIL.n99 VTAIL.n98 9.3005
R438 VTAIL.n75 VTAIL.n74 9.3005
R439 VTAIL.n70 VTAIL.n69 9.3005
R440 VTAIL.n81 VTAIL.n80 9.3005
R441 VTAIL.n83 VTAIL.n82 9.3005
R442 VTAIL.n66 VTAIL.n65 9.3005
R443 VTAIL.n89 VTAIL.n88 9.3005
R444 VTAIL.n91 VTAIL.n90 9.3005
R445 VTAIL.n92 VTAIL.n61 9.3005
R446 VTAIL.n163 VTAIL.n162 9.3005
R447 VTAIL.n114 VTAIL.n113 9.3005
R448 VTAIL.n157 VTAIL.n156 9.3005
R449 VTAIL.n155 VTAIL.n154 9.3005
R450 VTAIL.n131 VTAIL.n130 9.3005
R451 VTAIL.n126 VTAIL.n125 9.3005
R452 VTAIL.n137 VTAIL.n136 9.3005
R453 VTAIL.n139 VTAIL.n138 9.3005
R454 VTAIL.n122 VTAIL.n121 9.3005
R455 VTAIL.n145 VTAIL.n144 9.3005
R456 VTAIL.n147 VTAIL.n146 9.3005
R457 VTAIL.n148 VTAIL.n117 9.3005
R458 VTAIL.n352 VTAIL.n351 9.3005
R459 VTAIL.n347 VTAIL.n346 9.3005
R460 VTAIL.n358 VTAIL.n357 9.3005
R461 VTAIL.n360 VTAIL.n359 9.3005
R462 VTAIL.n343 VTAIL.n342 9.3005
R463 VTAIL.n366 VTAIL.n365 9.3005
R464 VTAIL.n368 VTAIL.n367 9.3005
R465 VTAIL.n340 VTAIL.n337 9.3005
R466 VTAIL.n383 VTAIL.n382 9.3005
R467 VTAIL.n334 VTAIL.n333 9.3005
R468 VTAIL.n377 VTAIL.n376 9.3005
R469 VTAIL.n375 VTAIL.n374 9.3005
R470 VTAIL.n296 VTAIL.n295 9.3005
R471 VTAIL.n291 VTAIL.n290 9.3005
R472 VTAIL.n302 VTAIL.n301 9.3005
R473 VTAIL.n304 VTAIL.n303 9.3005
R474 VTAIL.n287 VTAIL.n286 9.3005
R475 VTAIL.n310 VTAIL.n309 9.3005
R476 VTAIL.n312 VTAIL.n311 9.3005
R477 VTAIL.n284 VTAIL.n281 9.3005
R478 VTAIL.n327 VTAIL.n326 9.3005
R479 VTAIL.n278 VTAIL.n277 9.3005
R480 VTAIL.n321 VTAIL.n320 9.3005
R481 VTAIL.n319 VTAIL.n318 9.3005
R482 VTAIL.n242 VTAIL.n241 9.3005
R483 VTAIL.n237 VTAIL.n236 9.3005
R484 VTAIL.n248 VTAIL.n247 9.3005
R485 VTAIL.n250 VTAIL.n249 9.3005
R486 VTAIL.n233 VTAIL.n232 9.3005
R487 VTAIL.n256 VTAIL.n255 9.3005
R488 VTAIL.n258 VTAIL.n257 9.3005
R489 VTAIL.n230 VTAIL.n227 9.3005
R490 VTAIL.n273 VTAIL.n272 9.3005
R491 VTAIL.n224 VTAIL.n223 9.3005
R492 VTAIL.n267 VTAIL.n266 9.3005
R493 VTAIL.n265 VTAIL.n264 9.3005
R494 VTAIL.n186 VTAIL.n185 9.3005
R495 VTAIL.n181 VTAIL.n180 9.3005
R496 VTAIL.n192 VTAIL.n191 9.3005
R497 VTAIL.n194 VTAIL.n193 9.3005
R498 VTAIL.n177 VTAIL.n176 9.3005
R499 VTAIL.n200 VTAIL.n199 9.3005
R500 VTAIL.n202 VTAIL.n201 9.3005
R501 VTAIL.n174 VTAIL.n171 9.3005
R502 VTAIL.n217 VTAIL.n216 9.3005
R503 VTAIL.n168 VTAIL.n167 9.3005
R504 VTAIL.n211 VTAIL.n210 9.3005
R505 VTAIL.n209 VTAIL.n208 9.3005
R506 VTAIL.n410 VTAIL.n409 8.92171
R507 VTAIL.n26 VTAIL.n25 8.92171
R508 VTAIL.n80 VTAIL.n79 8.92171
R509 VTAIL.n136 VTAIL.n135 8.92171
R510 VTAIL.n357 VTAIL.n356 8.92171
R511 VTAIL.n301 VTAIL.n300 8.92171
R512 VTAIL.n247 VTAIL.n246 8.92171
R513 VTAIL.n191 VTAIL.n190 8.92171
R514 VTAIL.n406 VTAIL.n400 8.14595
R515 VTAIL.n22 VTAIL.n16 8.14595
R516 VTAIL.n76 VTAIL.n70 8.14595
R517 VTAIL.n132 VTAIL.n126 8.14595
R518 VTAIL.n353 VTAIL.n347 8.14595
R519 VTAIL.n297 VTAIL.n291 8.14595
R520 VTAIL.n243 VTAIL.n237 8.14595
R521 VTAIL.n187 VTAIL.n181 8.14595
R522 VTAIL.n405 VTAIL.n402 7.3702
R523 VTAIL.n21 VTAIL.n18 7.3702
R524 VTAIL.n75 VTAIL.n72 7.3702
R525 VTAIL.n131 VTAIL.n128 7.3702
R526 VTAIL.n352 VTAIL.n349 7.3702
R527 VTAIL.n296 VTAIL.n293 7.3702
R528 VTAIL.n242 VTAIL.n239 7.3702
R529 VTAIL.n186 VTAIL.n183 7.3702
R530 VTAIL.n406 VTAIL.n405 5.81868
R531 VTAIL.n22 VTAIL.n21 5.81868
R532 VTAIL.n76 VTAIL.n75 5.81868
R533 VTAIL.n132 VTAIL.n131 5.81868
R534 VTAIL.n353 VTAIL.n352 5.81868
R535 VTAIL.n297 VTAIL.n296 5.81868
R536 VTAIL.n243 VTAIL.n242 5.81868
R537 VTAIL.n187 VTAIL.n186 5.81868
R538 VTAIL.n409 VTAIL.n400 5.04292
R539 VTAIL.n25 VTAIL.n16 5.04292
R540 VTAIL.n79 VTAIL.n70 5.04292
R541 VTAIL.n135 VTAIL.n126 5.04292
R542 VTAIL.n356 VTAIL.n347 5.04292
R543 VTAIL.n300 VTAIL.n291 5.04292
R544 VTAIL.n246 VTAIL.n237 5.04292
R545 VTAIL.n190 VTAIL.n181 5.04292
R546 VTAIL.n410 VTAIL.n398 4.26717
R547 VTAIL.n26 VTAIL.n14 4.26717
R548 VTAIL.n80 VTAIL.n68 4.26717
R549 VTAIL.n136 VTAIL.n124 4.26717
R550 VTAIL.n357 VTAIL.n345 4.26717
R551 VTAIL.n301 VTAIL.n289 4.26717
R552 VTAIL.n247 VTAIL.n235 4.26717
R553 VTAIL.n191 VTAIL.n179 4.26717
R554 VTAIL.n414 VTAIL.n413 3.49141
R555 VTAIL.n438 VTAIL.n386 3.49141
R556 VTAIL.n30 VTAIL.n29 3.49141
R557 VTAIL.n54 VTAIL.n2 3.49141
R558 VTAIL.n84 VTAIL.n83 3.49141
R559 VTAIL.n108 VTAIL.n56 3.49141
R560 VTAIL.n140 VTAIL.n139 3.49141
R561 VTAIL.n164 VTAIL.n112 3.49141
R562 VTAIL.n384 VTAIL.n332 3.49141
R563 VTAIL.n361 VTAIL.n360 3.49141
R564 VTAIL.n328 VTAIL.n276 3.49141
R565 VTAIL.n305 VTAIL.n304 3.49141
R566 VTAIL.n274 VTAIL.n222 3.49141
R567 VTAIL.n251 VTAIL.n250 3.49141
R568 VTAIL.n218 VTAIL.n166 3.49141
R569 VTAIL.n195 VTAIL.n194 3.49141
R570 VTAIL.n404 VTAIL.n403 2.84303
R571 VTAIL.n20 VTAIL.n19 2.84303
R572 VTAIL.n74 VTAIL.n73 2.84303
R573 VTAIL.n130 VTAIL.n129 2.84303
R574 VTAIL.n351 VTAIL.n350 2.84303
R575 VTAIL.n295 VTAIL.n294 2.84303
R576 VTAIL.n241 VTAIL.n240 2.84303
R577 VTAIL.n185 VTAIL.n184 2.84303
R578 VTAIL.n417 VTAIL.n396 2.71565
R579 VTAIL.n436 VTAIL.n435 2.71565
R580 VTAIL.n33 VTAIL.n12 2.71565
R581 VTAIL.n52 VTAIL.n51 2.71565
R582 VTAIL.n87 VTAIL.n66 2.71565
R583 VTAIL.n106 VTAIL.n105 2.71565
R584 VTAIL.n143 VTAIL.n122 2.71565
R585 VTAIL.n162 VTAIL.n161 2.71565
R586 VTAIL.n382 VTAIL.n381 2.71565
R587 VTAIL.n364 VTAIL.n343 2.71565
R588 VTAIL.n326 VTAIL.n325 2.71565
R589 VTAIL.n308 VTAIL.n287 2.71565
R590 VTAIL.n272 VTAIL.n271 2.71565
R591 VTAIL.n254 VTAIL.n233 2.71565
R592 VTAIL.n216 VTAIL.n215 2.71565
R593 VTAIL.n198 VTAIL.n177 2.71565
R594 VTAIL.n0 VTAIL.t14 1.9805
R595 VTAIL.n0 VTAIL.t8 1.9805
R596 VTAIL.n110 VTAIL.t0 1.9805
R597 VTAIL.n110 VTAIL.t5 1.9805
R598 VTAIL.n330 VTAIL.t1 1.9805
R599 VTAIL.n330 VTAIL.t4 1.9805
R600 VTAIL.n220 VTAIL.t11 1.9805
R601 VTAIL.n220 VTAIL.t10 1.9805
R602 VTAIL.n418 VTAIL.n394 1.93989
R603 VTAIL.n432 VTAIL.n388 1.93989
R604 VTAIL.n34 VTAIL.n10 1.93989
R605 VTAIL.n48 VTAIL.n4 1.93989
R606 VTAIL.n88 VTAIL.n64 1.93989
R607 VTAIL.n102 VTAIL.n58 1.93989
R608 VTAIL.n144 VTAIL.n120 1.93989
R609 VTAIL.n158 VTAIL.n114 1.93989
R610 VTAIL.n378 VTAIL.n334 1.93989
R611 VTAIL.n365 VTAIL.n341 1.93989
R612 VTAIL.n322 VTAIL.n278 1.93989
R613 VTAIL.n309 VTAIL.n285 1.93989
R614 VTAIL.n268 VTAIL.n224 1.93989
R615 VTAIL.n255 VTAIL.n231 1.93989
R616 VTAIL.n212 VTAIL.n168 1.93989
R617 VTAIL.n199 VTAIL.n175 1.93989
R618 VTAIL.n221 VTAIL.n219 1.56084
R619 VTAIL.n275 VTAIL.n221 1.56084
R620 VTAIL.n331 VTAIL.n329 1.56084
R621 VTAIL.n385 VTAIL.n331 1.56084
R622 VTAIL.n165 VTAIL.n111 1.56084
R623 VTAIL.n111 VTAIL.n109 1.56084
R624 VTAIL.n55 VTAIL.n1 1.56084
R625 VTAIL VTAIL.n439 1.50266
R626 VTAIL.n423 VTAIL.n421 1.16414
R627 VTAIL.n431 VTAIL.n390 1.16414
R628 VTAIL.n39 VTAIL.n37 1.16414
R629 VTAIL.n47 VTAIL.n6 1.16414
R630 VTAIL.n93 VTAIL.n91 1.16414
R631 VTAIL.n101 VTAIL.n60 1.16414
R632 VTAIL.n149 VTAIL.n147 1.16414
R633 VTAIL.n157 VTAIL.n116 1.16414
R634 VTAIL.n377 VTAIL.n336 1.16414
R635 VTAIL.n369 VTAIL.n368 1.16414
R636 VTAIL.n321 VTAIL.n280 1.16414
R637 VTAIL.n313 VTAIL.n312 1.16414
R638 VTAIL.n267 VTAIL.n226 1.16414
R639 VTAIL.n259 VTAIL.n258 1.16414
R640 VTAIL.n211 VTAIL.n170 1.16414
R641 VTAIL.n203 VTAIL.n202 1.16414
R642 VTAIL.n329 VTAIL.n275 0.470328
R643 VTAIL.n109 VTAIL.n55 0.470328
R644 VTAIL.n422 VTAIL.n392 0.388379
R645 VTAIL.n428 VTAIL.n427 0.388379
R646 VTAIL.n38 VTAIL.n8 0.388379
R647 VTAIL.n44 VTAIL.n43 0.388379
R648 VTAIL.n92 VTAIL.n62 0.388379
R649 VTAIL.n98 VTAIL.n97 0.388379
R650 VTAIL.n148 VTAIL.n118 0.388379
R651 VTAIL.n154 VTAIL.n153 0.388379
R652 VTAIL.n374 VTAIL.n373 0.388379
R653 VTAIL.n340 VTAIL.n338 0.388379
R654 VTAIL.n318 VTAIL.n317 0.388379
R655 VTAIL.n284 VTAIL.n282 0.388379
R656 VTAIL.n264 VTAIL.n263 0.388379
R657 VTAIL.n230 VTAIL.n228 0.388379
R658 VTAIL.n208 VTAIL.n207 0.388379
R659 VTAIL.n174 VTAIL.n172 0.388379
R660 VTAIL.n404 VTAIL.n399 0.155672
R661 VTAIL.n411 VTAIL.n399 0.155672
R662 VTAIL.n412 VTAIL.n411 0.155672
R663 VTAIL.n412 VTAIL.n395 0.155672
R664 VTAIL.n419 VTAIL.n395 0.155672
R665 VTAIL.n420 VTAIL.n419 0.155672
R666 VTAIL.n420 VTAIL.n391 0.155672
R667 VTAIL.n429 VTAIL.n391 0.155672
R668 VTAIL.n430 VTAIL.n429 0.155672
R669 VTAIL.n430 VTAIL.n387 0.155672
R670 VTAIL.n437 VTAIL.n387 0.155672
R671 VTAIL.n20 VTAIL.n15 0.155672
R672 VTAIL.n27 VTAIL.n15 0.155672
R673 VTAIL.n28 VTAIL.n27 0.155672
R674 VTAIL.n28 VTAIL.n11 0.155672
R675 VTAIL.n35 VTAIL.n11 0.155672
R676 VTAIL.n36 VTAIL.n35 0.155672
R677 VTAIL.n36 VTAIL.n7 0.155672
R678 VTAIL.n45 VTAIL.n7 0.155672
R679 VTAIL.n46 VTAIL.n45 0.155672
R680 VTAIL.n46 VTAIL.n3 0.155672
R681 VTAIL.n53 VTAIL.n3 0.155672
R682 VTAIL.n74 VTAIL.n69 0.155672
R683 VTAIL.n81 VTAIL.n69 0.155672
R684 VTAIL.n82 VTAIL.n81 0.155672
R685 VTAIL.n82 VTAIL.n65 0.155672
R686 VTAIL.n89 VTAIL.n65 0.155672
R687 VTAIL.n90 VTAIL.n89 0.155672
R688 VTAIL.n90 VTAIL.n61 0.155672
R689 VTAIL.n99 VTAIL.n61 0.155672
R690 VTAIL.n100 VTAIL.n99 0.155672
R691 VTAIL.n100 VTAIL.n57 0.155672
R692 VTAIL.n107 VTAIL.n57 0.155672
R693 VTAIL.n130 VTAIL.n125 0.155672
R694 VTAIL.n137 VTAIL.n125 0.155672
R695 VTAIL.n138 VTAIL.n137 0.155672
R696 VTAIL.n138 VTAIL.n121 0.155672
R697 VTAIL.n145 VTAIL.n121 0.155672
R698 VTAIL.n146 VTAIL.n145 0.155672
R699 VTAIL.n146 VTAIL.n117 0.155672
R700 VTAIL.n155 VTAIL.n117 0.155672
R701 VTAIL.n156 VTAIL.n155 0.155672
R702 VTAIL.n156 VTAIL.n113 0.155672
R703 VTAIL.n163 VTAIL.n113 0.155672
R704 VTAIL.n383 VTAIL.n333 0.155672
R705 VTAIL.n376 VTAIL.n333 0.155672
R706 VTAIL.n376 VTAIL.n375 0.155672
R707 VTAIL.n375 VTAIL.n337 0.155672
R708 VTAIL.n367 VTAIL.n337 0.155672
R709 VTAIL.n367 VTAIL.n366 0.155672
R710 VTAIL.n366 VTAIL.n342 0.155672
R711 VTAIL.n359 VTAIL.n342 0.155672
R712 VTAIL.n359 VTAIL.n358 0.155672
R713 VTAIL.n358 VTAIL.n346 0.155672
R714 VTAIL.n351 VTAIL.n346 0.155672
R715 VTAIL.n327 VTAIL.n277 0.155672
R716 VTAIL.n320 VTAIL.n277 0.155672
R717 VTAIL.n320 VTAIL.n319 0.155672
R718 VTAIL.n319 VTAIL.n281 0.155672
R719 VTAIL.n311 VTAIL.n281 0.155672
R720 VTAIL.n311 VTAIL.n310 0.155672
R721 VTAIL.n310 VTAIL.n286 0.155672
R722 VTAIL.n303 VTAIL.n286 0.155672
R723 VTAIL.n303 VTAIL.n302 0.155672
R724 VTAIL.n302 VTAIL.n290 0.155672
R725 VTAIL.n295 VTAIL.n290 0.155672
R726 VTAIL.n273 VTAIL.n223 0.155672
R727 VTAIL.n266 VTAIL.n223 0.155672
R728 VTAIL.n266 VTAIL.n265 0.155672
R729 VTAIL.n265 VTAIL.n227 0.155672
R730 VTAIL.n257 VTAIL.n227 0.155672
R731 VTAIL.n257 VTAIL.n256 0.155672
R732 VTAIL.n256 VTAIL.n232 0.155672
R733 VTAIL.n249 VTAIL.n232 0.155672
R734 VTAIL.n249 VTAIL.n248 0.155672
R735 VTAIL.n248 VTAIL.n236 0.155672
R736 VTAIL.n241 VTAIL.n236 0.155672
R737 VTAIL.n217 VTAIL.n167 0.155672
R738 VTAIL.n210 VTAIL.n167 0.155672
R739 VTAIL.n210 VTAIL.n209 0.155672
R740 VTAIL.n209 VTAIL.n171 0.155672
R741 VTAIL.n201 VTAIL.n171 0.155672
R742 VTAIL.n201 VTAIL.n200 0.155672
R743 VTAIL.n200 VTAIL.n176 0.155672
R744 VTAIL.n193 VTAIL.n176 0.155672
R745 VTAIL.n193 VTAIL.n192 0.155672
R746 VTAIL.n192 VTAIL.n180 0.155672
R747 VTAIL.n185 VTAIL.n180 0.155672
R748 VTAIL VTAIL.n1 0.0586897
R749 B.n532 B.n109 585
R750 B.n109 B.n64 585
R751 B.n534 B.n533 585
R752 B.n536 B.n108 585
R753 B.n539 B.n538 585
R754 B.n540 B.n107 585
R755 B.n542 B.n541 585
R756 B.n544 B.n106 585
R757 B.n547 B.n546 585
R758 B.n548 B.n105 585
R759 B.n550 B.n549 585
R760 B.n552 B.n104 585
R761 B.n555 B.n554 585
R762 B.n556 B.n103 585
R763 B.n558 B.n557 585
R764 B.n560 B.n102 585
R765 B.n563 B.n562 585
R766 B.n564 B.n101 585
R767 B.n566 B.n565 585
R768 B.n568 B.n100 585
R769 B.n571 B.n570 585
R770 B.n572 B.n99 585
R771 B.n574 B.n573 585
R772 B.n576 B.n98 585
R773 B.n579 B.n578 585
R774 B.n580 B.n97 585
R775 B.n582 B.n581 585
R776 B.n584 B.n96 585
R777 B.n587 B.n586 585
R778 B.n588 B.n95 585
R779 B.n590 B.n589 585
R780 B.n592 B.n94 585
R781 B.n595 B.n594 585
R782 B.n596 B.n93 585
R783 B.n598 B.n597 585
R784 B.n600 B.n92 585
R785 B.n603 B.n602 585
R786 B.n605 B.n89 585
R787 B.n607 B.n606 585
R788 B.n609 B.n88 585
R789 B.n612 B.n611 585
R790 B.n613 B.n87 585
R791 B.n615 B.n614 585
R792 B.n617 B.n86 585
R793 B.n620 B.n619 585
R794 B.n621 B.n83 585
R795 B.n624 B.n623 585
R796 B.n626 B.n82 585
R797 B.n629 B.n628 585
R798 B.n630 B.n81 585
R799 B.n632 B.n631 585
R800 B.n634 B.n80 585
R801 B.n637 B.n636 585
R802 B.n638 B.n79 585
R803 B.n640 B.n639 585
R804 B.n642 B.n78 585
R805 B.n645 B.n644 585
R806 B.n646 B.n77 585
R807 B.n648 B.n647 585
R808 B.n650 B.n76 585
R809 B.n653 B.n652 585
R810 B.n654 B.n75 585
R811 B.n656 B.n655 585
R812 B.n658 B.n74 585
R813 B.n661 B.n660 585
R814 B.n662 B.n73 585
R815 B.n664 B.n663 585
R816 B.n666 B.n72 585
R817 B.n669 B.n668 585
R818 B.n670 B.n71 585
R819 B.n672 B.n671 585
R820 B.n674 B.n70 585
R821 B.n677 B.n676 585
R822 B.n678 B.n69 585
R823 B.n680 B.n679 585
R824 B.n682 B.n68 585
R825 B.n685 B.n684 585
R826 B.n686 B.n67 585
R827 B.n688 B.n687 585
R828 B.n690 B.n66 585
R829 B.n693 B.n692 585
R830 B.n694 B.n65 585
R831 B.n531 B.n63 585
R832 B.n697 B.n63 585
R833 B.n530 B.n62 585
R834 B.n698 B.n62 585
R835 B.n529 B.n61 585
R836 B.n699 B.n61 585
R837 B.n528 B.n527 585
R838 B.n527 B.n57 585
R839 B.n526 B.n56 585
R840 B.n705 B.n56 585
R841 B.n525 B.n55 585
R842 B.n706 B.n55 585
R843 B.n524 B.n54 585
R844 B.n707 B.n54 585
R845 B.n523 B.n522 585
R846 B.n522 B.n50 585
R847 B.n521 B.n49 585
R848 B.n713 B.n49 585
R849 B.n520 B.n48 585
R850 B.n714 B.n48 585
R851 B.n519 B.n47 585
R852 B.n715 B.n47 585
R853 B.n518 B.n517 585
R854 B.n517 B.n43 585
R855 B.n516 B.n42 585
R856 B.n721 B.n42 585
R857 B.n515 B.n41 585
R858 B.n722 B.n41 585
R859 B.n514 B.n40 585
R860 B.n723 B.n40 585
R861 B.n513 B.n512 585
R862 B.n512 B.n36 585
R863 B.n511 B.n35 585
R864 B.n729 B.n35 585
R865 B.n510 B.n34 585
R866 B.n730 B.n34 585
R867 B.n509 B.n33 585
R868 B.n731 B.n33 585
R869 B.n508 B.n507 585
R870 B.n507 B.n32 585
R871 B.n506 B.n28 585
R872 B.n737 B.n28 585
R873 B.n505 B.n27 585
R874 B.n738 B.n27 585
R875 B.n504 B.n26 585
R876 B.n739 B.n26 585
R877 B.n503 B.n502 585
R878 B.n502 B.n22 585
R879 B.n501 B.n21 585
R880 B.n745 B.n21 585
R881 B.n500 B.n20 585
R882 B.n746 B.n20 585
R883 B.n499 B.n19 585
R884 B.n747 B.n19 585
R885 B.n498 B.n497 585
R886 B.n497 B.n15 585
R887 B.n496 B.n14 585
R888 B.n753 B.n14 585
R889 B.n495 B.n13 585
R890 B.n754 B.n13 585
R891 B.n494 B.n12 585
R892 B.n755 B.n12 585
R893 B.n493 B.n492 585
R894 B.n492 B.n491 585
R895 B.n490 B.n489 585
R896 B.n490 B.n8 585
R897 B.n488 B.n7 585
R898 B.n762 B.n7 585
R899 B.n487 B.n6 585
R900 B.n763 B.n6 585
R901 B.n486 B.n5 585
R902 B.n764 B.n5 585
R903 B.n485 B.n484 585
R904 B.n484 B.n4 585
R905 B.n483 B.n110 585
R906 B.n483 B.n482 585
R907 B.n473 B.n111 585
R908 B.n112 B.n111 585
R909 B.n475 B.n474 585
R910 B.n476 B.n475 585
R911 B.n472 B.n117 585
R912 B.n117 B.n116 585
R913 B.n471 B.n470 585
R914 B.n470 B.n469 585
R915 B.n119 B.n118 585
R916 B.n120 B.n119 585
R917 B.n462 B.n461 585
R918 B.n463 B.n462 585
R919 B.n460 B.n125 585
R920 B.n125 B.n124 585
R921 B.n459 B.n458 585
R922 B.n458 B.n457 585
R923 B.n127 B.n126 585
R924 B.n128 B.n127 585
R925 B.n450 B.n449 585
R926 B.n451 B.n450 585
R927 B.n448 B.n133 585
R928 B.n133 B.n132 585
R929 B.n447 B.n446 585
R930 B.n446 B.n445 585
R931 B.n135 B.n134 585
R932 B.n438 B.n135 585
R933 B.n437 B.n436 585
R934 B.n439 B.n437 585
R935 B.n435 B.n140 585
R936 B.n140 B.n139 585
R937 B.n434 B.n433 585
R938 B.n433 B.n432 585
R939 B.n142 B.n141 585
R940 B.n143 B.n142 585
R941 B.n425 B.n424 585
R942 B.n426 B.n425 585
R943 B.n423 B.n148 585
R944 B.n148 B.n147 585
R945 B.n422 B.n421 585
R946 B.n421 B.n420 585
R947 B.n150 B.n149 585
R948 B.n151 B.n150 585
R949 B.n413 B.n412 585
R950 B.n414 B.n413 585
R951 B.n411 B.n156 585
R952 B.n156 B.n155 585
R953 B.n410 B.n409 585
R954 B.n409 B.n408 585
R955 B.n158 B.n157 585
R956 B.n159 B.n158 585
R957 B.n401 B.n400 585
R958 B.n402 B.n401 585
R959 B.n399 B.n163 585
R960 B.n167 B.n163 585
R961 B.n398 B.n397 585
R962 B.n397 B.n396 585
R963 B.n165 B.n164 585
R964 B.n166 B.n165 585
R965 B.n389 B.n388 585
R966 B.n390 B.n389 585
R967 B.n387 B.n172 585
R968 B.n172 B.n171 585
R969 B.n386 B.n385 585
R970 B.n385 B.n384 585
R971 B.n381 B.n176 585
R972 B.n380 B.n379 585
R973 B.n377 B.n177 585
R974 B.n377 B.n175 585
R975 B.n376 B.n375 585
R976 B.n374 B.n373 585
R977 B.n372 B.n179 585
R978 B.n370 B.n369 585
R979 B.n368 B.n180 585
R980 B.n367 B.n366 585
R981 B.n364 B.n181 585
R982 B.n362 B.n361 585
R983 B.n360 B.n182 585
R984 B.n359 B.n358 585
R985 B.n356 B.n183 585
R986 B.n354 B.n353 585
R987 B.n352 B.n184 585
R988 B.n351 B.n350 585
R989 B.n348 B.n185 585
R990 B.n346 B.n345 585
R991 B.n344 B.n186 585
R992 B.n343 B.n342 585
R993 B.n340 B.n187 585
R994 B.n338 B.n337 585
R995 B.n336 B.n188 585
R996 B.n335 B.n334 585
R997 B.n332 B.n189 585
R998 B.n330 B.n329 585
R999 B.n328 B.n190 585
R1000 B.n327 B.n326 585
R1001 B.n324 B.n191 585
R1002 B.n322 B.n321 585
R1003 B.n320 B.n192 585
R1004 B.n319 B.n318 585
R1005 B.n316 B.n193 585
R1006 B.n314 B.n313 585
R1007 B.n312 B.n194 585
R1008 B.n310 B.n309 585
R1009 B.n307 B.n197 585
R1010 B.n305 B.n304 585
R1011 B.n303 B.n198 585
R1012 B.n302 B.n301 585
R1013 B.n299 B.n199 585
R1014 B.n297 B.n296 585
R1015 B.n295 B.n200 585
R1016 B.n294 B.n293 585
R1017 B.n291 B.n290 585
R1018 B.n289 B.n288 585
R1019 B.n287 B.n205 585
R1020 B.n285 B.n284 585
R1021 B.n283 B.n206 585
R1022 B.n282 B.n281 585
R1023 B.n279 B.n207 585
R1024 B.n277 B.n276 585
R1025 B.n275 B.n208 585
R1026 B.n274 B.n273 585
R1027 B.n271 B.n209 585
R1028 B.n269 B.n268 585
R1029 B.n267 B.n210 585
R1030 B.n266 B.n265 585
R1031 B.n263 B.n211 585
R1032 B.n261 B.n260 585
R1033 B.n259 B.n212 585
R1034 B.n258 B.n257 585
R1035 B.n255 B.n213 585
R1036 B.n253 B.n252 585
R1037 B.n251 B.n214 585
R1038 B.n250 B.n249 585
R1039 B.n247 B.n215 585
R1040 B.n245 B.n244 585
R1041 B.n243 B.n216 585
R1042 B.n242 B.n241 585
R1043 B.n239 B.n217 585
R1044 B.n237 B.n236 585
R1045 B.n235 B.n218 585
R1046 B.n234 B.n233 585
R1047 B.n231 B.n219 585
R1048 B.n229 B.n228 585
R1049 B.n227 B.n220 585
R1050 B.n226 B.n225 585
R1051 B.n223 B.n221 585
R1052 B.n174 B.n173 585
R1053 B.n383 B.n382 585
R1054 B.n384 B.n383 585
R1055 B.n170 B.n169 585
R1056 B.n171 B.n170 585
R1057 B.n392 B.n391 585
R1058 B.n391 B.n390 585
R1059 B.n393 B.n168 585
R1060 B.n168 B.n166 585
R1061 B.n395 B.n394 585
R1062 B.n396 B.n395 585
R1063 B.n162 B.n161 585
R1064 B.n167 B.n162 585
R1065 B.n404 B.n403 585
R1066 B.n403 B.n402 585
R1067 B.n405 B.n160 585
R1068 B.n160 B.n159 585
R1069 B.n407 B.n406 585
R1070 B.n408 B.n407 585
R1071 B.n154 B.n153 585
R1072 B.n155 B.n154 585
R1073 B.n416 B.n415 585
R1074 B.n415 B.n414 585
R1075 B.n417 B.n152 585
R1076 B.n152 B.n151 585
R1077 B.n419 B.n418 585
R1078 B.n420 B.n419 585
R1079 B.n146 B.n145 585
R1080 B.n147 B.n146 585
R1081 B.n428 B.n427 585
R1082 B.n427 B.n426 585
R1083 B.n429 B.n144 585
R1084 B.n144 B.n143 585
R1085 B.n431 B.n430 585
R1086 B.n432 B.n431 585
R1087 B.n138 B.n137 585
R1088 B.n139 B.n138 585
R1089 B.n441 B.n440 585
R1090 B.n440 B.n439 585
R1091 B.n442 B.n136 585
R1092 B.n438 B.n136 585
R1093 B.n444 B.n443 585
R1094 B.n445 B.n444 585
R1095 B.n131 B.n130 585
R1096 B.n132 B.n131 585
R1097 B.n453 B.n452 585
R1098 B.n452 B.n451 585
R1099 B.n454 B.n129 585
R1100 B.n129 B.n128 585
R1101 B.n456 B.n455 585
R1102 B.n457 B.n456 585
R1103 B.n123 B.n122 585
R1104 B.n124 B.n123 585
R1105 B.n465 B.n464 585
R1106 B.n464 B.n463 585
R1107 B.n466 B.n121 585
R1108 B.n121 B.n120 585
R1109 B.n468 B.n467 585
R1110 B.n469 B.n468 585
R1111 B.n115 B.n114 585
R1112 B.n116 B.n115 585
R1113 B.n478 B.n477 585
R1114 B.n477 B.n476 585
R1115 B.n479 B.n113 585
R1116 B.n113 B.n112 585
R1117 B.n481 B.n480 585
R1118 B.n482 B.n481 585
R1119 B.n3 B.n0 585
R1120 B.n4 B.n3 585
R1121 B.n761 B.n1 585
R1122 B.n762 B.n761 585
R1123 B.n760 B.n759 585
R1124 B.n760 B.n8 585
R1125 B.n758 B.n9 585
R1126 B.n491 B.n9 585
R1127 B.n757 B.n756 585
R1128 B.n756 B.n755 585
R1129 B.n11 B.n10 585
R1130 B.n754 B.n11 585
R1131 B.n752 B.n751 585
R1132 B.n753 B.n752 585
R1133 B.n750 B.n16 585
R1134 B.n16 B.n15 585
R1135 B.n749 B.n748 585
R1136 B.n748 B.n747 585
R1137 B.n18 B.n17 585
R1138 B.n746 B.n18 585
R1139 B.n744 B.n743 585
R1140 B.n745 B.n744 585
R1141 B.n742 B.n23 585
R1142 B.n23 B.n22 585
R1143 B.n741 B.n740 585
R1144 B.n740 B.n739 585
R1145 B.n25 B.n24 585
R1146 B.n738 B.n25 585
R1147 B.n736 B.n735 585
R1148 B.n737 B.n736 585
R1149 B.n734 B.n29 585
R1150 B.n32 B.n29 585
R1151 B.n733 B.n732 585
R1152 B.n732 B.n731 585
R1153 B.n31 B.n30 585
R1154 B.n730 B.n31 585
R1155 B.n728 B.n727 585
R1156 B.n729 B.n728 585
R1157 B.n726 B.n37 585
R1158 B.n37 B.n36 585
R1159 B.n725 B.n724 585
R1160 B.n724 B.n723 585
R1161 B.n39 B.n38 585
R1162 B.n722 B.n39 585
R1163 B.n720 B.n719 585
R1164 B.n721 B.n720 585
R1165 B.n718 B.n44 585
R1166 B.n44 B.n43 585
R1167 B.n717 B.n716 585
R1168 B.n716 B.n715 585
R1169 B.n46 B.n45 585
R1170 B.n714 B.n46 585
R1171 B.n712 B.n711 585
R1172 B.n713 B.n712 585
R1173 B.n710 B.n51 585
R1174 B.n51 B.n50 585
R1175 B.n709 B.n708 585
R1176 B.n708 B.n707 585
R1177 B.n53 B.n52 585
R1178 B.n706 B.n53 585
R1179 B.n704 B.n703 585
R1180 B.n705 B.n704 585
R1181 B.n702 B.n58 585
R1182 B.n58 B.n57 585
R1183 B.n701 B.n700 585
R1184 B.n700 B.n699 585
R1185 B.n60 B.n59 585
R1186 B.n698 B.n60 585
R1187 B.n696 B.n695 585
R1188 B.n697 B.n696 585
R1189 B.n765 B.n764 585
R1190 B.n763 B.n2 585
R1191 B.n696 B.n65 540.549
R1192 B.n109 B.n63 540.549
R1193 B.n385 B.n174 540.549
R1194 B.n383 B.n176 540.549
R1195 B.n84 B.t16 368.202
R1196 B.n90 B.t8 368.202
R1197 B.n201 B.t19 368.202
R1198 B.n195 B.t12 368.202
R1199 B.n90 B.t10 282.75
R1200 B.n201 B.t21 282.75
R1201 B.n84 B.t17 282.75
R1202 B.n195 B.t15 282.75
R1203 B.n535 B.n64 256.663
R1204 B.n537 B.n64 256.663
R1205 B.n543 B.n64 256.663
R1206 B.n545 B.n64 256.663
R1207 B.n551 B.n64 256.663
R1208 B.n553 B.n64 256.663
R1209 B.n559 B.n64 256.663
R1210 B.n561 B.n64 256.663
R1211 B.n567 B.n64 256.663
R1212 B.n569 B.n64 256.663
R1213 B.n575 B.n64 256.663
R1214 B.n577 B.n64 256.663
R1215 B.n583 B.n64 256.663
R1216 B.n585 B.n64 256.663
R1217 B.n591 B.n64 256.663
R1218 B.n593 B.n64 256.663
R1219 B.n599 B.n64 256.663
R1220 B.n601 B.n64 256.663
R1221 B.n608 B.n64 256.663
R1222 B.n610 B.n64 256.663
R1223 B.n616 B.n64 256.663
R1224 B.n618 B.n64 256.663
R1225 B.n625 B.n64 256.663
R1226 B.n627 B.n64 256.663
R1227 B.n633 B.n64 256.663
R1228 B.n635 B.n64 256.663
R1229 B.n641 B.n64 256.663
R1230 B.n643 B.n64 256.663
R1231 B.n649 B.n64 256.663
R1232 B.n651 B.n64 256.663
R1233 B.n657 B.n64 256.663
R1234 B.n659 B.n64 256.663
R1235 B.n665 B.n64 256.663
R1236 B.n667 B.n64 256.663
R1237 B.n673 B.n64 256.663
R1238 B.n675 B.n64 256.663
R1239 B.n681 B.n64 256.663
R1240 B.n683 B.n64 256.663
R1241 B.n689 B.n64 256.663
R1242 B.n691 B.n64 256.663
R1243 B.n378 B.n175 256.663
R1244 B.n178 B.n175 256.663
R1245 B.n371 B.n175 256.663
R1246 B.n365 B.n175 256.663
R1247 B.n363 B.n175 256.663
R1248 B.n357 B.n175 256.663
R1249 B.n355 B.n175 256.663
R1250 B.n349 B.n175 256.663
R1251 B.n347 B.n175 256.663
R1252 B.n341 B.n175 256.663
R1253 B.n339 B.n175 256.663
R1254 B.n333 B.n175 256.663
R1255 B.n331 B.n175 256.663
R1256 B.n325 B.n175 256.663
R1257 B.n323 B.n175 256.663
R1258 B.n317 B.n175 256.663
R1259 B.n315 B.n175 256.663
R1260 B.n308 B.n175 256.663
R1261 B.n306 B.n175 256.663
R1262 B.n300 B.n175 256.663
R1263 B.n298 B.n175 256.663
R1264 B.n292 B.n175 256.663
R1265 B.n204 B.n175 256.663
R1266 B.n286 B.n175 256.663
R1267 B.n280 B.n175 256.663
R1268 B.n278 B.n175 256.663
R1269 B.n272 B.n175 256.663
R1270 B.n270 B.n175 256.663
R1271 B.n264 B.n175 256.663
R1272 B.n262 B.n175 256.663
R1273 B.n256 B.n175 256.663
R1274 B.n254 B.n175 256.663
R1275 B.n248 B.n175 256.663
R1276 B.n246 B.n175 256.663
R1277 B.n240 B.n175 256.663
R1278 B.n238 B.n175 256.663
R1279 B.n232 B.n175 256.663
R1280 B.n230 B.n175 256.663
R1281 B.n224 B.n175 256.663
R1282 B.n222 B.n175 256.663
R1283 B.n767 B.n766 256.663
R1284 B.n91 B.t11 247.648
R1285 B.n202 B.t20 247.648
R1286 B.n85 B.t18 247.648
R1287 B.n196 B.t14 247.648
R1288 B.n692 B.n690 163.367
R1289 B.n688 B.n67 163.367
R1290 B.n684 B.n682 163.367
R1291 B.n680 B.n69 163.367
R1292 B.n676 B.n674 163.367
R1293 B.n672 B.n71 163.367
R1294 B.n668 B.n666 163.367
R1295 B.n664 B.n73 163.367
R1296 B.n660 B.n658 163.367
R1297 B.n656 B.n75 163.367
R1298 B.n652 B.n650 163.367
R1299 B.n648 B.n77 163.367
R1300 B.n644 B.n642 163.367
R1301 B.n640 B.n79 163.367
R1302 B.n636 B.n634 163.367
R1303 B.n632 B.n81 163.367
R1304 B.n628 B.n626 163.367
R1305 B.n624 B.n83 163.367
R1306 B.n619 B.n617 163.367
R1307 B.n615 B.n87 163.367
R1308 B.n611 B.n609 163.367
R1309 B.n607 B.n89 163.367
R1310 B.n602 B.n600 163.367
R1311 B.n598 B.n93 163.367
R1312 B.n594 B.n592 163.367
R1313 B.n590 B.n95 163.367
R1314 B.n586 B.n584 163.367
R1315 B.n582 B.n97 163.367
R1316 B.n578 B.n576 163.367
R1317 B.n574 B.n99 163.367
R1318 B.n570 B.n568 163.367
R1319 B.n566 B.n101 163.367
R1320 B.n562 B.n560 163.367
R1321 B.n558 B.n103 163.367
R1322 B.n554 B.n552 163.367
R1323 B.n550 B.n105 163.367
R1324 B.n546 B.n544 163.367
R1325 B.n542 B.n107 163.367
R1326 B.n538 B.n536 163.367
R1327 B.n534 B.n109 163.367
R1328 B.n385 B.n172 163.367
R1329 B.n389 B.n172 163.367
R1330 B.n389 B.n165 163.367
R1331 B.n397 B.n165 163.367
R1332 B.n397 B.n163 163.367
R1333 B.n401 B.n163 163.367
R1334 B.n401 B.n158 163.367
R1335 B.n409 B.n158 163.367
R1336 B.n409 B.n156 163.367
R1337 B.n413 B.n156 163.367
R1338 B.n413 B.n150 163.367
R1339 B.n421 B.n150 163.367
R1340 B.n421 B.n148 163.367
R1341 B.n425 B.n148 163.367
R1342 B.n425 B.n142 163.367
R1343 B.n433 B.n142 163.367
R1344 B.n433 B.n140 163.367
R1345 B.n437 B.n140 163.367
R1346 B.n437 B.n135 163.367
R1347 B.n446 B.n135 163.367
R1348 B.n446 B.n133 163.367
R1349 B.n450 B.n133 163.367
R1350 B.n450 B.n127 163.367
R1351 B.n458 B.n127 163.367
R1352 B.n458 B.n125 163.367
R1353 B.n462 B.n125 163.367
R1354 B.n462 B.n119 163.367
R1355 B.n470 B.n119 163.367
R1356 B.n470 B.n117 163.367
R1357 B.n475 B.n117 163.367
R1358 B.n475 B.n111 163.367
R1359 B.n483 B.n111 163.367
R1360 B.n484 B.n483 163.367
R1361 B.n484 B.n5 163.367
R1362 B.n6 B.n5 163.367
R1363 B.n7 B.n6 163.367
R1364 B.n490 B.n7 163.367
R1365 B.n492 B.n490 163.367
R1366 B.n492 B.n12 163.367
R1367 B.n13 B.n12 163.367
R1368 B.n14 B.n13 163.367
R1369 B.n497 B.n14 163.367
R1370 B.n497 B.n19 163.367
R1371 B.n20 B.n19 163.367
R1372 B.n21 B.n20 163.367
R1373 B.n502 B.n21 163.367
R1374 B.n502 B.n26 163.367
R1375 B.n27 B.n26 163.367
R1376 B.n28 B.n27 163.367
R1377 B.n507 B.n28 163.367
R1378 B.n507 B.n33 163.367
R1379 B.n34 B.n33 163.367
R1380 B.n35 B.n34 163.367
R1381 B.n512 B.n35 163.367
R1382 B.n512 B.n40 163.367
R1383 B.n41 B.n40 163.367
R1384 B.n42 B.n41 163.367
R1385 B.n517 B.n42 163.367
R1386 B.n517 B.n47 163.367
R1387 B.n48 B.n47 163.367
R1388 B.n49 B.n48 163.367
R1389 B.n522 B.n49 163.367
R1390 B.n522 B.n54 163.367
R1391 B.n55 B.n54 163.367
R1392 B.n56 B.n55 163.367
R1393 B.n527 B.n56 163.367
R1394 B.n527 B.n61 163.367
R1395 B.n62 B.n61 163.367
R1396 B.n63 B.n62 163.367
R1397 B.n379 B.n377 163.367
R1398 B.n377 B.n376 163.367
R1399 B.n373 B.n372 163.367
R1400 B.n370 B.n180 163.367
R1401 B.n366 B.n364 163.367
R1402 B.n362 B.n182 163.367
R1403 B.n358 B.n356 163.367
R1404 B.n354 B.n184 163.367
R1405 B.n350 B.n348 163.367
R1406 B.n346 B.n186 163.367
R1407 B.n342 B.n340 163.367
R1408 B.n338 B.n188 163.367
R1409 B.n334 B.n332 163.367
R1410 B.n330 B.n190 163.367
R1411 B.n326 B.n324 163.367
R1412 B.n322 B.n192 163.367
R1413 B.n318 B.n316 163.367
R1414 B.n314 B.n194 163.367
R1415 B.n309 B.n307 163.367
R1416 B.n305 B.n198 163.367
R1417 B.n301 B.n299 163.367
R1418 B.n297 B.n200 163.367
R1419 B.n293 B.n291 163.367
R1420 B.n288 B.n287 163.367
R1421 B.n285 B.n206 163.367
R1422 B.n281 B.n279 163.367
R1423 B.n277 B.n208 163.367
R1424 B.n273 B.n271 163.367
R1425 B.n269 B.n210 163.367
R1426 B.n265 B.n263 163.367
R1427 B.n261 B.n212 163.367
R1428 B.n257 B.n255 163.367
R1429 B.n253 B.n214 163.367
R1430 B.n249 B.n247 163.367
R1431 B.n245 B.n216 163.367
R1432 B.n241 B.n239 163.367
R1433 B.n237 B.n218 163.367
R1434 B.n233 B.n231 163.367
R1435 B.n229 B.n220 163.367
R1436 B.n225 B.n223 163.367
R1437 B.n383 B.n170 163.367
R1438 B.n391 B.n170 163.367
R1439 B.n391 B.n168 163.367
R1440 B.n395 B.n168 163.367
R1441 B.n395 B.n162 163.367
R1442 B.n403 B.n162 163.367
R1443 B.n403 B.n160 163.367
R1444 B.n407 B.n160 163.367
R1445 B.n407 B.n154 163.367
R1446 B.n415 B.n154 163.367
R1447 B.n415 B.n152 163.367
R1448 B.n419 B.n152 163.367
R1449 B.n419 B.n146 163.367
R1450 B.n427 B.n146 163.367
R1451 B.n427 B.n144 163.367
R1452 B.n431 B.n144 163.367
R1453 B.n431 B.n138 163.367
R1454 B.n440 B.n138 163.367
R1455 B.n440 B.n136 163.367
R1456 B.n444 B.n136 163.367
R1457 B.n444 B.n131 163.367
R1458 B.n452 B.n131 163.367
R1459 B.n452 B.n129 163.367
R1460 B.n456 B.n129 163.367
R1461 B.n456 B.n123 163.367
R1462 B.n464 B.n123 163.367
R1463 B.n464 B.n121 163.367
R1464 B.n468 B.n121 163.367
R1465 B.n468 B.n115 163.367
R1466 B.n477 B.n115 163.367
R1467 B.n477 B.n113 163.367
R1468 B.n481 B.n113 163.367
R1469 B.n481 B.n3 163.367
R1470 B.n765 B.n3 163.367
R1471 B.n761 B.n2 163.367
R1472 B.n761 B.n760 163.367
R1473 B.n760 B.n9 163.367
R1474 B.n756 B.n9 163.367
R1475 B.n756 B.n11 163.367
R1476 B.n752 B.n11 163.367
R1477 B.n752 B.n16 163.367
R1478 B.n748 B.n16 163.367
R1479 B.n748 B.n18 163.367
R1480 B.n744 B.n18 163.367
R1481 B.n744 B.n23 163.367
R1482 B.n740 B.n23 163.367
R1483 B.n740 B.n25 163.367
R1484 B.n736 B.n25 163.367
R1485 B.n736 B.n29 163.367
R1486 B.n732 B.n29 163.367
R1487 B.n732 B.n31 163.367
R1488 B.n728 B.n31 163.367
R1489 B.n728 B.n37 163.367
R1490 B.n724 B.n37 163.367
R1491 B.n724 B.n39 163.367
R1492 B.n720 B.n39 163.367
R1493 B.n720 B.n44 163.367
R1494 B.n716 B.n44 163.367
R1495 B.n716 B.n46 163.367
R1496 B.n712 B.n46 163.367
R1497 B.n712 B.n51 163.367
R1498 B.n708 B.n51 163.367
R1499 B.n708 B.n53 163.367
R1500 B.n704 B.n53 163.367
R1501 B.n704 B.n58 163.367
R1502 B.n700 B.n58 163.367
R1503 B.n700 B.n60 163.367
R1504 B.n696 B.n60 163.367
R1505 B.n384 B.n175 100.099
R1506 B.n697 B.n64 100.099
R1507 B.n691 B.n65 71.676
R1508 B.n690 B.n689 71.676
R1509 B.n683 B.n67 71.676
R1510 B.n682 B.n681 71.676
R1511 B.n675 B.n69 71.676
R1512 B.n674 B.n673 71.676
R1513 B.n667 B.n71 71.676
R1514 B.n666 B.n665 71.676
R1515 B.n659 B.n73 71.676
R1516 B.n658 B.n657 71.676
R1517 B.n651 B.n75 71.676
R1518 B.n650 B.n649 71.676
R1519 B.n643 B.n77 71.676
R1520 B.n642 B.n641 71.676
R1521 B.n635 B.n79 71.676
R1522 B.n634 B.n633 71.676
R1523 B.n627 B.n81 71.676
R1524 B.n626 B.n625 71.676
R1525 B.n618 B.n83 71.676
R1526 B.n617 B.n616 71.676
R1527 B.n610 B.n87 71.676
R1528 B.n609 B.n608 71.676
R1529 B.n601 B.n89 71.676
R1530 B.n600 B.n599 71.676
R1531 B.n593 B.n93 71.676
R1532 B.n592 B.n591 71.676
R1533 B.n585 B.n95 71.676
R1534 B.n584 B.n583 71.676
R1535 B.n577 B.n97 71.676
R1536 B.n576 B.n575 71.676
R1537 B.n569 B.n99 71.676
R1538 B.n568 B.n567 71.676
R1539 B.n561 B.n101 71.676
R1540 B.n560 B.n559 71.676
R1541 B.n553 B.n103 71.676
R1542 B.n552 B.n551 71.676
R1543 B.n545 B.n105 71.676
R1544 B.n544 B.n543 71.676
R1545 B.n537 B.n107 71.676
R1546 B.n536 B.n535 71.676
R1547 B.n535 B.n534 71.676
R1548 B.n538 B.n537 71.676
R1549 B.n543 B.n542 71.676
R1550 B.n546 B.n545 71.676
R1551 B.n551 B.n550 71.676
R1552 B.n554 B.n553 71.676
R1553 B.n559 B.n558 71.676
R1554 B.n562 B.n561 71.676
R1555 B.n567 B.n566 71.676
R1556 B.n570 B.n569 71.676
R1557 B.n575 B.n574 71.676
R1558 B.n578 B.n577 71.676
R1559 B.n583 B.n582 71.676
R1560 B.n586 B.n585 71.676
R1561 B.n591 B.n590 71.676
R1562 B.n594 B.n593 71.676
R1563 B.n599 B.n598 71.676
R1564 B.n602 B.n601 71.676
R1565 B.n608 B.n607 71.676
R1566 B.n611 B.n610 71.676
R1567 B.n616 B.n615 71.676
R1568 B.n619 B.n618 71.676
R1569 B.n625 B.n624 71.676
R1570 B.n628 B.n627 71.676
R1571 B.n633 B.n632 71.676
R1572 B.n636 B.n635 71.676
R1573 B.n641 B.n640 71.676
R1574 B.n644 B.n643 71.676
R1575 B.n649 B.n648 71.676
R1576 B.n652 B.n651 71.676
R1577 B.n657 B.n656 71.676
R1578 B.n660 B.n659 71.676
R1579 B.n665 B.n664 71.676
R1580 B.n668 B.n667 71.676
R1581 B.n673 B.n672 71.676
R1582 B.n676 B.n675 71.676
R1583 B.n681 B.n680 71.676
R1584 B.n684 B.n683 71.676
R1585 B.n689 B.n688 71.676
R1586 B.n692 B.n691 71.676
R1587 B.n378 B.n176 71.676
R1588 B.n376 B.n178 71.676
R1589 B.n372 B.n371 71.676
R1590 B.n365 B.n180 71.676
R1591 B.n364 B.n363 71.676
R1592 B.n357 B.n182 71.676
R1593 B.n356 B.n355 71.676
R1594 B.n349 B.n184 71.676
R1595 B.n348 B.n347 71.676
R1596 B.n341 B.n186 71.676
R1597 B.n340 B.n339 71.676
R1598 B.n333 B.n188 71.676
R1599 B.n332 B.n331 71.676
R1600 B.n325 B.n190 71.676
R1601 B.n324 B.n323 71.676
R1602 B.n317 B.n192 71.676
R1603 B.n316 B.n315 71.676
R1604 B.n308 B.n194 71.676
R1605 B.n307 B.n306 71.676
R1606 B.n300 B.n198 71.676
R1607 B.n299 B.n298 71.676
R1608 B.n292 B.n200 71.676
R1609 B.n291 B.n204 71.676
R1610 B.n287 B.n286 71.676
R1611 B.n280 B.n206 71.676
R1612 B.n279 B.n278 71.676
R1613 B.n272 B.n208 71.676
R1614 B.n271 B.n270 71.676
R1615 B.n264 B.n210 71.676
R1616 B.n263 B.n262 71.676
R1617 B.n256 B.n212 71.676
R1618 B.n255 B.n254 71.676
R1619 B.n248 B.n214 71.676
R1620 B.n247 B.n246 71.676
R1621 B.n240 B.n216 71.676
R1622 B.n239 B.n238 71.676
R1623 B.n232 B.n218 71.676
R1624 B.n231 B.n230 71.676
R1625 B.n224 B.n220 71.676
R1626 B.n223 B.n222 71.676
R1627 B.n379 B.n378 71.676
R1628 B.n373 B.n178 71.676
R1629 B.n371 B.n370 71.676
R1630 B.n366 B.n365 71.676
R1631 B.n363 B.n362 71.676
R1632 B.n358 B.n357 71.676
R1633 B.n355 B.n354 71.676
R1634 B.n350 B.n349 71.676
R1635 B.n347 B.n346 71.676
R1636 B.n342 B.n341 71.676
R1637 B.n339 B.n338 71.676
R1638 B.n334 B.n333 71.676
R1639 B.n331 B.n330 71.676
R1640 B.n326 B.n325 71.676
R1641 B.n323 B.n322 71.676
R1642 B.n318 B.n317 71.676
R1643 B.n315 B.n314 71.676
R1644 B.n309 B.n308 71.676
R1645 B.n306 B.n305 71.676
R1646 B.n301 B.n300 71.676
R1647 B.n298 B.n297 71.676
R1648 B.n293 B.n292 71.676
R1649 B.n288 B.n204 71.676
R1650 B.n286 B.n285 71.676
R1651 B.n281 B.n280 71.676
R1652 B.n278 B.n277 71.676
R1653 B.n273 B.n272 71.676
R1654 B.n270 B.n269 71.676
R1655 B.n265 B.n264 71.676
R1656 B.n262 B.n261 71.676
R1657 B.n257 B.n256 71.676
R1658 B.n254 B.n253 71.676
R1659 B.n249 B.n248 71.676
R1660 B.n246 B.n245 71.676
R1661 B.n241 B.n240 71.676
R1662 B.n238 B.n237 71.676
R1663 B.n233 B.n232 71.676
R1664 B.n230 B.n229 71.676
R1665 B.n225 B.n224 71.676
R1666 B.n222 B.n174 71.676
R1667 B.n766 B.n765 71.676
R1668 B.n766 B.n2 71.676
R1669 B.n622 B.n85 59.5399
R1670 B.n604 B.n91 59.5399
R1671 B.n203 B.n202 59.5399
R1672 B.n311 B.n196 59.5399
R1673 B.n384 B.n171 48.9694
R1674 B.n390 B.n171 48.9694
R1675 B.n390 B.n166 48.9694
R1676 B.n396 B.n166 48.9694
R1677 B.n396 B.n167 48.9694
R1678 B.n402 B.n159 48.9694
R1679 B.n408 B.n159 48.9694
R1680 B.n408 B.n155 48.9694
R1681 B.n414 B.n155 48.9694
R1682 B.n414 B.n151 48.9694
R1683 B.n420 B.n151 48.9694
R1684 B.n420 B.n147 48.9694
R1685 B.n426 B.n147 48.9694
R1686 B.n432 B.n143 48.9694
R1687 B.n432 B.n139 48.9694
R1688 B.n439 B.n139 48.9694
R1689 B.n439 B.n438 48.9694
R1690 B.n445 B.n132 48.9694
R1691 B.n451 B.n132 48.9694
R1692 B.n451 B.n128 48.9694
R1693 B.n457 B.n128 48.9694
R1694 B.n463 B.n124 48.9694
R1695 B.n463 B.n120 48.9694
R1696 B.n469 B.n120 48.9694
R1697 B.n469 B.n116 48.9694
R1698 B.n476 B.n116 48.9694
R1699 B.n482 B.n112 48.9694
R1700 B.n482 B.n4 48.9694
R1701 B.n764 B.n4 48.9694
R1702 B.n764 B.n763 48.9694
R1703 B.n763 B.n762 48.9694
R1704 B.n762 B.n8 48.9694
R1705 B.n491 B.n8 48.9694
R1706 B.n755 B.n754 48.9694
R1707 B.n754 B.n753 48.9694
R1708 B.n753 B.n15 48.9694
R1709 B.n747 B.n15 48.9694
R1710 B.n747 B.n746 48.9694
R1711 B.n745 B.n22 48.9694
R1712 B.n739 B.n22 48.9694
R1713 B.n739 B.n738 48.9694
R1714 B.n738 B.n737 48.9694
R1715 B.n731 B.n32 48.9694
R1716 B.n731 B.n730 48.9694
R1717 B.n730 B.n729 48.9694
R1718 B.n729 B.n36 48.9694
R1719 B.n723 B.n722 48.9694
R1720 B.n722 B.n721 48.9694
R1721 B.n721 B.n43 48.9694
R1722 B.n715 B.n43 48.9694
R1723 B.n715 B.n714 48.9694
R1724 B.n714 B.n713 48.9694
R1725 B.n713 B.n50 48.9694
R1726 B.n707 B.n50 48.9694
R1727 B.n706 B.n705 48.9694
R1728 B.n705 B.n57 48.9694
R1729 B.n699 B.n57 48.9694
R1730 B.n699 B.n698 48.9694
R1731 B.n698 B.n697 48.9694
R1732 B.n457 B.t5 44.6486
R1733 B.t1 B.n745 44.6486
R1734 B.t3 B.n112 37.4473
R1735 B.n491 B.t7 37.4473
R1736 B.n167 B.t13 36.007
R1737 B.t2 B.n143 36.007
R1738 B.t6 B.n36 36.007
R1739 B.t9 B.n706 36.007
R1740 B.n382 B.n381 35.1225
R1741 B.n386 B.n173 35.1225
R1742 B.n532 B.n531 35.1225
R1743 B.n695 B.n694 35.1225
R1744 B.n85 B.n84 35.1035
R1745 B.n91 B.n90 35.1035
R1746 B.n202 B.n201 35.1035
R1747 B.n196 B.n195 35.1035
R1748 B.n438 B.t0 28.8057
R1749 B.n32 B.t4 28.8057
R1750 B.n445 B.t0 20.1642
R1751 B.n737 B.t4 20.1642
R1752 B B.n767 18.0485
R1753 B.n402 B.t13 12.9629
R1754 B.n426 B.t2 12.9629
R1755 B.n723 B.t6 12.9629
R1756 B.n707 B.t9 12.9629
R1757 B.n476 B.t3 11.5226
R1758 B.n755 B.t7 11.5226
R1759 B.n382 B.n169 10.6151
R1760 B.n392 B.n169 10.6151
R1761 B.n393 B.n392 10.6151
R1762 B.n394 B.n393 10.6151
R1763 B.n394 B.n161 10.6151
R1764 B.n404 B.n161 10.6151
R1765 B.n405 B.n404 10.6151
R1766 B.n406 B.n405 10.6151
R1767 B.n406 B.n153 10.6151
R1768 B.n416 B.n153 10.6151
R1769 B.n417 B.n416 10.6151
R1770 B.n418 B.n417 10.6151
R1771 B.n418 B.n145 10.6151
R1772 B.n428 B.n145 10.6151
R1773 B.n429 B.n428 10.6151
R1774 B.n430 B.n429 10.6151
R1775 B.n430 B.n137 10.6151
R1776 B.n441 B.n137 10.6151
R1777 B.n442 B.n441 10.6151
R1778 B.n443 B.n442 10.6151
R1779 B.n443 B.n130 10.6151
R1780 B.n453 B.n130 10.6151
R1781 B.n454 B.n453 10.6151
R1782 B.n455 B.n454 10.6151
R1783 B.n455 B.n122 10.6151
R1784 B.n465 B.n122 10.6151
R1785 B.n466 B.n465 10.6151
R1786 B.n467 B.n466 10.6151
R1787 B.n467 B.n114 10.6151
R1788 B.n478 B.n114 10.6151
R1789 B.n479 B.n478 10.6151
R1790 B.n480 B.n479 10.6151
R1791 B.n480 B.n0 10.6151
R1792 B.n381 B.n380 10.6151
R1793 B.n380 B.n177 10.6151
R1794 B.n375 B.n177 10.6151
R1795 B.n375 B.n374 10.6151
R1796 B.n374 B.n179 10.6151
R1797 B.n369 B.n179 10.6151
R1798 B.n369 B.n368 10.6151
R1799 B.n368 B.n367 10.6151
R1800 B.n367 B.n181 10.6151
R1801 B.n361 B.n181 10.6151
R1802 B.n361 B.n360 10.6151
R1803 B.n360 B.n359 10.6151
R1804 B.n359 B.n183 10.6151
R1805 B.n353 B.n183 10.6151
R1806 B.n353 B.n352 10.6151
R1807 B.n352 B.n351 10.6151
R1808 B.n351 B.n185 10.6151
R1809 B.n345 B.n185 10.6151
R1810 B.n345 B.n344 10.6151
R1811 B.n344 B.n343 10.6151
R1812 B.n343 B.n187 10.6151
R1813 B.n337 B.n187 10.6151
R1814 B.n337 B.n336 10.6151
R1815 B.n336 B.n335 10.6151
R1816 B.n335 B.n189 10.6151
R1817 B.n329 B.n189 10.6151
R1818 B.n329 B.n328 10.6151
R1819 B.n328 B.n327 10.6151
R1820 B.n327 B.n191 10.6151
R1821 B.n321 B.n191 10.6151
R1822 B.n321 B.n320 10.6151
R1823 B.n320 B.n319 10.6151
R1824 B.n319 B.n193 10.6151
R1825 B.n313 B.n193 10.6151
R1826 B.n313 B.n312 10.6151
R1827 B.n310 B.n197 10.6151
R1828 B.n304 B.n197 10.6151
R1829 B.n304 B.n303 10.6151
R1830 B.n303 B.n302 10.6151
R1831 B.n302 B.n199 10.6151
R1832 B.n296 B.n199 10.6151
R1833 B.n296 B.n295 10.6151
R1834 B.n295 B.n294 10.6151
R1835 B.n290 B.n289 10.6151
R1836 B.n289 B.n205 10.6151
R1837 B.n284 B.n205 10.6151
R1838 B.n284 B.n283 10.6151
R1839 B.n283 B.n282 10.6151
R1840 B.n282 B.n207 10.6151
R1841 B.n276 B.n207 10.6151
R1842 B.n276 B.n275 10.6151
R1843 B.n275 B.n274 10.6151
R1844 B.n274 B.n209 10.6151
R1845 B.n268 B.n209 10.6151
R1846 B.n268 B.n267 10.6151
R1847 B.n267 B.n266 10.6151
R1848 B.n266 B.n211 10.6151
R1849 B.n260 B.n211 10.6151
R1850 B.n260 B.n259 10.6151
R1851 B.n259 B.n258 10.6151
R1852 B.n258 B.n213 10.6151
R1853 B.n252 B.n213 10.6151
R1854 B.n252 B.n251 10.6151
R1855 B.n251 B.n250 10.6151
R1856 B.n250 B.n215 10.6151
R1857 B.n244 B.n215 10.6151
R1858 B.n244 B.n243 10.6151
R1859 B.n243 B.n242 10.6151
R1860 B.n242 B.n217 10.6151
R1861 B.n236 B.n217 10.6151
R1862 B.n236 B.n235 10.6151
R1863 B.n235 B.n234 10.6151
R1864 B.n234 B.n219 10.6151
R1865 B.n228 B.n219 10.6151
R1866 B.n228 B.n227 10.6151
R1867 B.n227 B.n226 10.6151
R1868 B.n226 B.n221 10.6151
R1869 B.n221 B.n173 10.6151
R1870 B.n387 B.n386 10.6151
R1871 B.n388 B.n387 10.6151
R1872 B.n388 B.n164 10.6151
R1873 B.n398 B.n164 10.6151
R1874 B.n399 B.n398 10.6151
R1875 B.n400 B.n399 10.6151
R1876 B.n400 B.n157 10.6151
R1877 B.n410 B.n157 10.6151
R1878 B.n411 B.n410 10.6151
R1879 B.n412 B.n411 10.6151
R1880 B.n412 B.n149 10.6151
R1881 B.n422 B.n149 10.6151
R1882 B.n423 B.n422 10.6151
R1883 B.n424 B.n423 10.6151
R1884 B.n424 B.n141 10.6151
R1885 B.n434 B.n141 10.6151
R1886 B.n435 B.n434 10.6151
R1887 B.n436 B.n435 10.6151
R1888 B.n436 B.n134 10.6151
R1889 B.n447 B.n134 10.6151
R1890 B.n448 B.n447 10.6151
R1891 B.n449 B.n448 10.6151
R1892 B.n449 B.n126 10.6151
R1893 B.n459 B.n126 10.6151
R1894 B.n460 B.n459 10.6151
R1895 B.n461 B.n460 10.6151
R1896 B.n461 B.n118 10.6151
R1897 B.n471 B.n118 10.6151
R1898 B.n472 B.n471 10.6151
R1899 B.n474 B.n472 10.6151
R1900 B.n474 B.n473 10.6151
R1901 B.n473 B.n110 10.6151
R1902 B.n485 B.n110 10.6151
R1903 B.n486 B.n485 10.6151
R1904 B.n487 B.n486 10.6151
R1905 B.n488 B.n487 10.6151
R1906 B.n489 B.n488 10.6151
R1907 B.n493 B.n489 10.6151
R1908 B.n494 B.n493 10.6151
R1909 B.n495 B.n494 10.6151
R1910 B.n496 B.n495 10.6151
R1911 B.n498 B.n496 10.6151
R1912 B.n499 B.n498 10.6151
R1913 B.n500 B.n499 10.6151
R1914 B.n501 B.n500 10.6151
R1915 B.n503 B.n501 10.6151
R1916 B.n504 B.n503 10.6151
R1917 B.n505 B.n504 10.6151
R1918 B.n506 B.n505 10.6151
R1919 B.n508 B.n506 10.6151
R1920 B.n509 B.n508 10.6151
R1921 B.n510 B.n509 10.6151
R1922 B.n511 B.n510 10.6151
R1923 B.n513 B.n511 10.6151
R1924 B.n514 B.n513 10.6151
R1925 B.n515 B.n514 10.6151
R1926 B.n516 B.n515 10.6151
R1927 B.n518 B.n516 10.6151
R1928 B.n519 B.n518 10.6151
R1929 B.n520 B.n519 10.6151
R1930 B.n521 B.n520 10.6151
R1931 B.n523 B.n521 10.6151
R1932 B.n524 B.n523 10.6151
R1933 B.n525 B.n524 10.6151
R1934 B.n526 B.n525 10.6151
R1935 B.n528 B.n526 10.6151
R1936 B.n529 B.n528 10.6151
R1937 B.n530 B.n529 10.6151
R1938 B.n531 B.n530 10.6151
R1939 B.n759 B.n1 10.6151
R1940 B.n759 B.n758 10.6151
R1941 B.n758 B.n757 10.6151
R1942 B.n757 B.n10 10.6151
R1943 B.n751 B.n10 10.6151
R1944 B.n751 B.n750 10.6151
R1945 B.n750 B.n749 10.6151
R1946 B.n749 B.n17 10.6151
R1947 B.n743 B.n17 10.6151
R1948 B.n743 B.n742 10.6151
R1949 B.n742 B.n741 10.6151
R1950 B.n741 B.n24 10.6151
R1951 B.n735 B.n24 10.6151
R1952 B.n735 B.n734 10.6151
R1953 B.n734 B.n733 10.6151
R1954 B.n733 B.n30 10.6151
R1955 B.n727 B.n30 10.6151
R1956 B.n727 B.n726 10.6151
R1957 B.n726 B.n725 10.6151
R1958 B.n725 B.n38 10.6151
R1959 B.n719 B.n38 10.6151
R1960 B.n719 B.n718 10.6151
R1961 B.n718 B.n717 10.6151
R1962 B.n717 B.n45 10.6151
R1963 B.n711 B.n45 10.6151
R1964 B.n711 B.n710 10.6151
R1965 B.n710 B.n709 10.6151
R1966 B.n709 B.n52 10.6151
R1967 B.n703 B.n52 10.6151
R1968 B.n703 B.n702 10.6151
R1969 B.n702 B.n701 10.6151
R1970 B.n701 B.n59 10.6151
R1971 B.n695 B.n59 10.6151
R1972 B.n694 B.n693 10.6151
R1973 B.n693 B.n66 10.6151
R1974 B.n687 B.n66 10.6151
R1975 B.n687 B.n686 10.6151
R1976 B.n686 B.n685 10.6151
R1977 B.n685 B.n68 10.6151
R1978 B.n679 B.n68 10.6151
R1979 B.n679 B.n678 10.6151
R1980 B.n678 B.n677 10.6151
R1981 B.n677 B.n70 10.6151
R1982 B.n671 B.n70 10.6151
R1983 B.n671 B.n670 10.6151
R1984 B.n670 B.n669 10.6151
R1985 B.n669 B.n72 10.6151
R1986 B.n663 B.n72 10.6151
R1987 B.n663 B.n662 10.6151
R1988 B.n662 B.n661 10.6151
R1989 B.n661 B.n74 10.6151
R1990 B.n655 B.n74 10.6151
R1991 B.n655 B.n654 10.6151
R1992 B.n654 B.n653 10.6151
R1993 B.n653 B.n76 10.6151
R1994 B.n647 B.n76 10.6151
R1995 B.n647 B.n646 10.6151
R1996 B.n646 B.n645 10.6151
R1997 B.n645 B.n78 10.6151
R1998 B.n639 B.n78 10.6151
R1999 B.n639 B.n638 10.6151
R2000 B.n638 B.n637 10.6151
R2001 B.n637 B.n80 10.6151
R2002 B.n631 B.n80 10.6151
R2003 B.n631 B.n630 10.6151
R2004 B.n630 B.n629 10.6151
R2005 B.n629 B.n82 10.6151
R2006 B.n623 B.n82 10.6151
R2007 B.n621 B.n620 10.6151
R2008 B.n620 B.n86 10.6151
R2009 B.n614 B.n86 10.6151
R2010 B.n614 B.n613 10.6151
R2011 B.n613 B.n612 10.6151
R2012 B.n612 B.n88 10.6151
R2013 B.n606 B.n88 10.6151
R2014 B.n606 B.n605 10.6151
R2015 B.n603 B.n92 10.6151
R2016 B.n597 B.n92 10.6151
R2017 B.n597 B.n596 10.6151
R2018 B.n596 B.n595 10.6151
R2019 B.n595 B.n94 10.6151
R2020 B.n589 B.n94 10.6151
R2021 B.n589 B.n588 10.6151
R2022 B.n588 B.n587 10.6151
R2023 B.n587 B.n96 10.6151
R2024 B.n581 B.n96 10.6151
R2025 B.n581 B.n580 10.6151
R2026 B.n580 B.n579 10.6151
R2027 B.n579 B.n98 10.6151
R2028 B.n573 B.n98 10.6151
R2029 B.n573 B.n572 10.6151
R2030 B.n572 B.n571 10.6151
R2031 B.n571 B.n100 10.6151
R2032 B.n565 B.n100 10.6151
R2033 B.n565 B.n564 10.6151
R2034 B.n564 B.n563 10.6151
R2035 B.n563 B.n102 10.6151
R2036 B.n557 B.n102 10.6151
R2037 B.n557 B.n556 10.6151
R2038 B.n556 B.n555 10.6151
R2039 B.n555 B.n104 10.6151
R2040 B.n549 B.n104 10.6151
R2041 B.n549 B.n548 10.6151
R2042 B.n548 B.n547 10.6151
R2043 B.n547 B.n106 10.6151
R2044 B.n541 B.n106 10.6151
R2045 B.n541 B.n540 10.6151
R2046 B.n540 B.n539 10.6151
R2047 B.n539 B.n108 10.6151
R2048 B.n533 B.n108 10.6151
R2049 B.n533 B.n532 10.6151
R2050 B.n767 B.n0 8.11757
R2051 B.n767 B.n1 8.11757
R2052 B.n311 B.n310 6.5566
R2053 B.n294 B.n203 6.5566
R2054 B.n622 B.n621 6.5566
R2055 B.n605 B.n604 6.5566
R2056 B.t5 B.n124 4.32129
R2057 B.n746 B.t1 4.32129
R2058 B.n312 B.n311 4.05904
R2059 B.n290 B.n203 4.05904
R2060 B.n623 B.n622 4.05904
R2061 B.n604 B.n603 4.05904
R2062 VP.n11 VP.t7 196.924
R2063 VP.n26 VP.n25 175.317
R2064 VP.n46 VP.n45 175.317
R2065 VP.n24 VP.n23 175.317
R2066 VP.n25 VP.t3 162.839
R2067 VP.n31 VP.t4 162.839
R2068 VP.n38 VP.t2 162.839
R2069 VP.n45 VP.t1 162.839
R2070 VP.n23 VP.t0 162.839
R2071 VP.n16 VP.t6 162.839
R2072 VP.n10 VP.t5 162.839
R2073 VP.n12 VP.n9 161.3
R2074 VP.n14 VP.n13 161.3
R2075 VP.n15 VP.n8 161.3
R2076 VP.n18 VP.n17 161.3
R2077 VP.n19 VP.n7 161.3
R2078 VP.n21 VP.n20 161.3
R2079 VP.n22 VP.n6 161.3
R2080 VP.n44 VP.n0 161.3
R2081 VP.n43 VP.n42 161.3
R2082 VP.n41 VP.n1 161.3
R2083 VP.n40 VP.n39 161.3
R2084 VP.n37 VP.n2 161.3
R2085 VP.n36 VP.n35 161.3
R2086 VP.n34 VP.n3 161.3
R2087 VP.n33 VP.n32 161.3
R2088 VP.n30 VP.n4 161.3
R2089 VP.n29 VP.n28 161.3
R2090 VP.n27 VP.n5 161.3
R2091 VP.n30 VP.n29 56.5617
R2092 VP.n43 VP.n1 56.5617
R2093 VP.n21 VP.n7 56.5617
R2094 VP.n11 VP.n10 46.7161
R2095 VP.n26 VP.n24 44.0687
R2096 VP.n36 VP.n3 40.577
R2097 VP.n37 VP.n36 40.577
R2098 VP.n15 VP.n14 40.577
R2099 VP.n14 VP.n9 40.577
R2100 VP.n29 VP.n5 24.5923
R2101 VP.n32 VP.n30 24.5923
R2102 VP.n39 VP.n1 24.5923
R2103 VP.n44 VP.n43 24.5923
R2104 VP.n22 VP.n21 24.5923
R2105 VP.n17 VP.n7 24.5923
R2106 VP.n31 VP.n3 19.9199
R2107 VP.n38 VP.n37 19.9199
R2108 VP.n16 VP.n15 19.9199
R2109 VP.n10 VP.n9 19.9199
R2110 VP.n12 VP.n11 17.7081
R2111 VP.n25 VP.n5 10.575
R2112 VP.n45 VP.n44 10.575
R2113 VP.n23 VP.n22 10.575
R2114 VP.n32 VP.n31 4.67295
R2115 VP.n39 VP.n38 4.67295
R2116 VP.n17 VP.n16 4.67295
R2117 VP.n13 VP.n12 0.189894
R2118 VP.n13 VP.n8 0.189894
R2119 VP.n18 VP.n8 0.189894
R2120 VP.n19 VP.n18 0.189894
R2121 VP.n20 VP.n19 0.189894
R2122 VP.n20 VP.n6 0.189894
R2123 VP.n24 VP.n6 0.189894
R2124 VP.n27 VP.n26 0.189894
R2125 VP.n28 VP.n27 0.189894
R2126 VP.n28 VP.n4 0.189894
R2127 VP.n33 VP.n4 0.189894
R2128 VP.n34 VP.n33 0.189894
R2129 VP.n35 VP.n34 0.189894
R2130 VP.n35 VP.n2 0.189894
R2131 VP.n40 VP.n2 0.189894
R2132 VP.n41 VP.n40 0.189894
R2133 VP.n42 VP.n41 0.189894
R2134 VP.n42 VP.n0 0.189894
R2135 VP.n46 VP.n0 0.189894
R2136 VP VP.n46 0.0516364
R2137 VDD1 VDD1.n0 64.2545
R2138 VDD1.n3 VDD1.n2 64.1407
R2139 VDD1.n3 VDD1.n1 64.1407
R2140 VDD1.n5 VDD1.n4 63.4159
R2141 VDD1.n5 VDD1.n3 39.9405
R2142 VDD1.n4 VDD1.t1 1.9805
R2143 VDD1.n4 VDD1.t7 1.9805
R2144 VDD1.n0 VDD1.t0 1.9805
R2145 VDD1.n0 VDD1.t2 1.9805
R2146 VDD1.n2 VDD1.t5 1.9805
R2147 VDD1.n2 VDD1.t6 1.9805
R2148 VDD1.n1 VDD1.t4 1.9805
R2149 VDD1.n1 VDD1.t3 1.9805
R2150 VDD1 VDD1.n5 0.722483
C0 VDD1 VDD2 1.213f
C1 VTAIL VP 6.47888f
C2 VN VDD2 6.3409f
C3 VDD1 VN 0.150103f
C4 VP VDD2 0.400891f
C5 VDD1 VP 6.59086f
C6 VP VN 5.91788f
C7 VTAIL VDD2 7.61028f
C8 VDD1 VTAIL 7.56337f
C9 VTAIL VN 6.46477f
C10 VDD2 B 4.094556f
C11 VDD1 B 4.415521f
C12 VTAIL B 8.461731f
C13 VN B 11.10359f
C14 VP B 9.546025f
C15 VDD1.t0 B 0.199406f
C16 VDD1.t2 B 0.199406f
C17 VDD1.n0 B 1.76181f
C18 VDD1.t4 B 0.199406f
C19 VDD1.t3 B 0.199406f
C20 VDD1.n1 B 1.76099f
C21 VDD1.t5 B 0.199406f
C22 VDD1.t6 B 0.199406f
C23 VDD1.n2 B 1.76099f
C24 VDD1.n3 B 2.57609f
C25 VDD1.t1 B 0.199406f
C26 VDD1.t7 B 0.199406f
C27 VDD1.n4 B 1.75645f
C28 VDD1.n5 B 2.45657f
C29 VP.n0 B 0.032072f
C30 VP.t1 B 1.2859f
C31 VP.n1 B 0.051946f
C32 VP.n2 B 0.032072f
C33 VP.t2 B 1.2859f
C34 VP.n3 B 0.057829f
C35 VP.n4 B 0.032072f
C36 VP.n5 B 0.042739f
C37 VP.n6 B 0.032072f
C38 VP.t0 B 1.2859f
C39 VP.n7 B 0.051946f
C40 VP.n8 B 0.032072f
C41 VP.t6 B 1.2859f
C42 VP.n9 B 0.057829f
C43 VP.t7 B 1.38894f
C44 VP.t5 B 1.2859f
C45 VP.n10 B 0.540887f
C46 VP.n11 B 0.542021f
C47 VP.n12 B 0.202743f
C48 VP.n13 B 0.032072f
C49 VP.n14 B 0.025904f
C50 VP.n15 B 0.057829f
C51 VP.n16 B 0.472775f
C52 VP.n17 B 0.035692f
C53 VP.n18 B 0.032072f
C54 VP.n19 B 0.032072f
C55 VP.n20 B 0.032072f
C56 VP.n21 B 0.041298f
C57 VP.n22 B 0.042739f
C58 VP.n23 B 0.53803f
C59 VP.n24 B 1.43811f
C60 VP.t3 B 1.2859f
C61 VP.n25 B 0.53803f
C62 VP.n26 B 1.46435f
C63 VP.n27 B 0.032072f
C64 VP.n28 B 0.032072f
C65 VP.n29 B 0.041298f
C66 VP.n30 B 0.051946f
C67 VP.t4 B 1.2859f
C68 VP.n31 B 0.472775f
C69 VP.n32 B 0.035692f
C70 VP.n33 B 0.032072f
C71 VP.n34 B 0.032072f
C72 VP.n35 B 0.032072f
C73 VP.n36 B 0.025904f
C74 VP.n37 B 0.057829f
C75 VP.n38 B 0.472775f
C76 VP.n39 B 0.035692f
C77 VP.n40 B 0.032072f
C78 VP.n41 B 0.032072f
C79 VP.n42 B 0.032072f
C80 VP.n43 B 0.041298f
C81 VP.n44 B 0.042739f
C82 VP.n45 B 0.53803f
C83 VP.n46 B 0.030525f
C84 VTAIL.t14 B 0.156469f
C85 VTAIL.t8 B 0.156469f
C86 VTAIL.n0 B 1.32215f
C87 VTAIL.n1 B 0.29341f
C88 VTAIL.n2 B 0.026763f
C89 VTAIL.n3 B 0.0198f
C90 VTAIL.n4 B 0.01064f
C91 VTAIL.n5 B 0.025149f
C92 VTAIL.n6 B 0.011266f
C93 VTAIL.n7 B 0.0198f
C94 VTAIL.n8 B 0.010953f
C95 VTAIL.n9 B 0.025149f
C96 VTAIL.n10 B 0.011266f
C97 VTAIL.n11 B 0.0198f
C98 VTAIL.n12 B 0.01064f
C99 VTAIL.n13 B 0.025149f
C100 VTAIL.n14 B 0.011266f
C101 VTAIL.n15 B 0.0198f
C102 VTAIL.n16 B 0.01064f
C103 VTAIL.n17 B 0.018862f
C104 VTAIL.n18 B 0.017778f
C105 VTAIL.t13 B 0.042263f
C106 VTAIL.n19 B 0.127558f
C107 VTAIL.n20 B 0.822753f
C108 VTAIL.n21 B 0.01064f
C109 VTAIL.n22 B 0.011266f
C110 VTAIL.n23 B 0.025149f
C111 VTAIL.n24 B 0.025149f
C112 VTAIL.n25 B 0.011266f
C113 VTAIL.n26 B 0.01064f
C114 VTAIL.n27 B 0.0198f
C115 VTAIL.n28 B 0.0198f
C116 VTAIL.n29 B 0.01064f
C117 VTAIL.n30 B 0.011266f
C118 VTAIL.n31 B 0.025149f
C119 VTAIL.n32 B 0.025149f
C120 VTAIL.n33 B 0.011266f
C121 VTAIL.n34 B 0.01064f
C122 VTAIL.n35 B 0.0198f
C123 VTAIL.n36 B 0.0198f
C124 VTAIL.n37 B 0.01064f
C125 VTAIL.n38 B 0.01064f
C126 VTAIL.n39 B 0.011266f
C127 VTAIL.n40 B 0.025149f
C128 VTAIL.n41 B 0.025149f
C129 VTAIL.n42 B 0.025149f
C130 VTAIL.n43 B 0.010953f
C131 VTAIL.n44 B 0.01064f
C132 VTAIL.n45 B 0.0198f
C133 VTAIL.n46 B 0.0198f
C134 VTAIL.n47 B 0.01064f
C135 VTAIL.n48 B 0.011266f
C136 VTAIL.n49 B 0.025149f
C137 VTAIL.n50 B 0.052553f
C138 VTAIL.n51 B 0.011266f
C139 VTAIL.n52 B 0.01064f
C140 VTAIL.n53 B 0.04685f
C141 VTAIL.n54 B 0.029244f
C142 VTAIL.n55 B 0.14705f
C143 VTAIL.n56 B 0.026763f
C144 VTAIL.n57 B 0.0198f
C145 VTAIL.n58 B 0.01064f
C146 VTAIL.n59 B 0.025149f
C147 VTAIL.n60 B 0.011266f
C148 VTAIL.n61 B 0.0198f
C149 VTAIL.n62 B 0.010953f
C150 VTAIL.n63 B 0.025149f
C151 VTAIL.n64 B 0.011266f
C152 VTAIL.n65 B 0.0198f
C153 VTAIL.n66 B 0.01064f
C154 VTAIL.n67 B 0.025149f
C155 VTAIL.n68 B 0.011266f
C156 VTAIL.n69 B 0.0198f
C157 VTAIL.n70 B 0.01064f
C158 VTAIL.n71 B 0.018862f
C159 VTAIL.n72 B 0.017778f
C160 VTAIL.t3 B 0.042263f
C161 VTAIL.n73 B 0.127558f
C162 VTAIL.n74 B 0.822753f
C163 VTAIL.n75 B 0.01064f
C164 VTAIL.n76 B 0.011266f
C165 VTAIL.n77 B 0.025149f
C166 VTAIL.n78 B 0.025149f
C167 VTAIL.n79 B 0.011266f
C168 VTAIL.n80 B 0.01064f
C169 VTAIL.n81 B 0.0198f
C170 VTAIL.n82 B 0.0198f
C171 VTAIL.n83 B 0.01064f
C172 VTAIL.n84 B 0.011266f
C173 VTAIL.n85 B 0.025149f
C174 VTAIL.n86 B 0.025149f
C175 VTAIL.n87 B 0.011266f
C176 VTAIL.n88 B 0.01064f
C177 VTAIL.n89 B 0.0198f
C178 VTAIL.n90 B 0.0198f
C179 VTAIL.n91 B 0.01064f
C180 VTAIL.n92 B 0.01064f
C181 VTAIL.n93 B 0.011266f
C182 VTAIL.n94 B 0.025149f
C183 VTAIL.n95 B 0.025149f
C184 VTAIL.n96 B 0.025149f
C185 VTAIL.n97 B 0.010953f
C186 VTAIL.n98 B 0.01064f
C187 VTAIL.n99 B 0.0198f
C188 VTAIL.n100 B 0.0198f
C189 VTAIL.n101 B 0.01064f
C190 VTAIL.n102 B 0.011266f
C191 VTAIL.n103 B 0.025149f
C192 VTAIL.n104 B 0.052553f
C193 VTAIL.n105 B 0.011266f
C194 VTAIL.n106 B 0.01064f
C195 VTAIL.n107 B 0.04685f
C196 VTAIL.n108 B 0.029244f
C197 VTAIL.n109 B 0.14705f
C198 VTAIL.t0 B 0.156469f
C199 VTAIL.t5 B 0.156469f
C200 VTAIL.n110 B 1.32215f
C201 VTAIL.n111 B 0.38925f
C202 VTAIL.n112 B 0.026763f
C203 VTAIL.n113 B 0.0198f
C204 VTAIL.n114 B 0.01064f
C205 VTAIL.n115 B 0.025149f
C206 VTAIL.n116 B 0.011266f
C207 VTAIL.n117 B 0.0198f
C208 VTAIL.n118 B 0.010953f
C209 VTAIL.n119 B 0.025149f
C210 VTAIL.n120 B 0.011266f
C211 VTAIL.n121 B 0.0198f
C212 VTAIL.n122 B 0.01064f
C213 VTAIL.n123 B 0.025149f
C214 VTAIL.n124 B 0.011266f
C215 VTAIL.n125 B 0.0198f
C216 VTAIL.n126 B 0.01064f
C217 VTAIL.n127 B 0.018862f
C218 VTAIL.n128 B 0.017778f
C219 VTAIL.t2 B 0.042263f
C220 VTAIL.n129 B 0.127558f
C221 VTAIL.n130 B 0.822753f
C222 VTAIL.n131 B 0.01064f
C223 VTAIL.n132 B 0.011266f
C224 VTAIL.n133 B 0.025149f
C225 VTAIL.n134 B 0.025149f
C226 VTAIL.n135 B 0.011266f
C227 VTAIL.n136 B 0.01064f
C228 VTAIL.n137 B 0.0198f
C229 VTAIL.n138 B 0.0198f
C230 VTAIL.n139 B 0.01064f
C231 VTAIL.n140 B 0.011266f
C232 VTAIL.n141 B 0.025149f
C233 VTAIL.n142 B 0.025149f
C234 VTAIL.n143 B 0.011266f
C235 VTAIL.n144 B 0.01064f
C236 VTAIL.n145 B 0.0198f
C237 VTAIL.n146 B 0.0198f
C238 VTAIL.n147 B 0.01064f
C239 VTAIL.n148 B 0.01064f
C240 VTAIL.n149 B 0.011266f
C241 VTAIL.n150 B 0.025149f
C242 VTAIL.n151 B 0.025149f
C243 VTAIL.n152 B 0.025149f
C244 VTAIL.n153 B 0.010953f
C245 VTAIL.n154 B 0.01064f
C246 VTAIL.n155 B 0.0198f
C247 VTAIL.n156 B 0.0198f
C248 VTAIL.n157 B 0.01064f
C249 VTAIL.n158 B 0.011266f
C250 VTAIL.n159 B 0.025149f
C251 VTAIL.n160 B 0.052553f
C252 VTAIL.n161 B 0.011266f
C253 VTAIL.n162 B 0.01064f
C254 VTAIL.n163 B 0.04685f
C255 VTAIL.n164 B 0.029244f
C256 VTAIL.n165 B 1.0356f
C257 VTAIL.n166 B 0.026763f
C258 VTAIL.n167 B 0.0198f
C259 VTAIL.n168 B 0.01064f
C260 VTAIL.n169 B 0.025149f
C261 VTAIL.n170 B 0.011266f
C262 VTAIL.n171 B 0.0198f
C263 VTAIL.n172 B 0.010953f
C264 VTAIL.n173 B 0.025149f
C265 VTAIL.n174 B 0.01064f
C266 VTAIL.n175 B 0.011266f
C267 VTAIL.n176 B 0.0198f
C268 VTAIL.n177 B 0.01064f
C269 VTAIL.n178 B 0.025149f
C270 VTAIL.n179 B 0.011266f
C271 VTAIL.n180 B 0.0198f
C272 VTAIL.n181 B 0.01064f
C273 VTAIL.n182 B 0.018862f
C274 VTAIL.n183 B 0.017778f
C275 VTAIL.t15 B 0.042263f
C276 VTAIL.n184 B 0.127558f
C277 VTAIL.n185 B 0.822753f
C278 VTAIL.n186 B 0.01064f
C279 VTAIL.n187 B 0.011266f
C280 VTAIL.n188 B 0.025149f
C281 VTAIL.n189 B 0.025149f
C282 VTAIL.n190 B 0.011266f
C283 VTAIL.n191 B 0.01064f
C284 VTAIL.n192 B 0.0198f
C285 VTAIL.n193 B 0.0198f
C286 VTAIL.n194 B 0.01064f
C287 VTAIL.n195 B 0.011266f
C288 VTAIL.n196 B 0.025149f
C289 VTAIL.n197 B 0.025149f
C290 VTAIL.n198 B 0.011266f
C291 VTAIL.n199 B 0.01064f
C292 VTAIL.n200 B 0.0198f
C293 VTAIL.n201 B 0.0198f
C294 VTAIL.n202 B 0.01064f
C295 VTAIL.n203 B 0.011266f
C296 VTAIL.n204 B 0.025149f
C297 VTAIL.n205 B 0.025149f
C298 VTAIL.n206 B 0.025149f
C299 VTAIL.n207 B 0.010953f
C300 VTAIL.n208 B 0.01064f
C301 VTAIL.n209 B 0.0198f
C302 VTAIL.n210 B 0.0198f
C303 VTAIL.n211 B 0.01064f
C304 VTAIL.n212 B 0.011266f
C305 VTAIL.n213 B 0.025149f
C306 VTAIL.n214 B 0.052553f
C307 VTAIL.n215 B 0.011266f
C308 VTAIL.n216 B 0.01064f
C309 VTAIL.n217 B 0.04685f
C310 VTAIL.n218 B 0.029244f
C311 VTAIL.n219 B 1.0356f
C312 VTAIL.t11 B 0.156469f
C313 VTAIL.t10 B 0.156469f
C314 VTAIL.n220 B 1.32216f
C315 VTAIL.n221 B 0.389242f
C316 VTAIL.n222 B 0.026763f
C317 VTAIL.n223 B 0.0198f
C318 VTAIL.n224 B 0.01064f
C319 VTAIL.n225 B 0.025149f
C320 VTAIL.n226 B 0.011266f
C321 VTAIL.n227 B 0.0198f
C322 VTAIL.n228 B 0.010953f
C323 VTAIL.n229 B 0.025149f
C324 VTAIL.n230 B 0.01064f
C325 VTAIL.n231 B 0.011266f
C326 VTAIL.n232 B 0.0198f
C327 VTAIL.n233 B 0.01064f
C328 VTAIL.n234 B 0.025149f
C329 VTAIL.n235 B 0.011266f
C330 VTAIL.n236 B 0.0198f
C331 VTAIL.n237 B 0.01064f
C332 VTAIL.n238 B 0.018862f
C333 VTAIL.n239 B 0.017778f
C334 VTAIL.t12 B 0.042263f
C335 VTAIL.n240 B 0.127558f
C336 VTAIL.n241 B 0.822753f
C337 VTAIL.n242 B 0.01064f
C338 VTAIL.n243 B 0.011266f
C339 VTAIL.n244 B 0.025149f
C340 VTAIL.n245 B 0.025149f
C341 VTAIL.n246 B 0.011266f
C342 VTAIL.n247 B 0.01064f
C343 VTAIL.n248 B 0.0198f
C344 VTAIL.n249 B 0.0198f
C345 VTAIL.n250 B 0.01064f
C346 VTAIL.n251 B 0.011266f
C347 VTAIL.n252 B 0.025149f
C348 VTAIL.n253 B 0.025149f
C349 VTAIL.n254 B 0.011266f
C350 VTAIL.n255 B 0.01064f
C351 VTAIL.n256 B 0.0198f
C352 VTAIL.n257 B 0.0198f
C353 VTAIL.n258 B 0.01064f
C354 VTAIL.n259 B 0.011266f
C355 VTAIL.n260 B 0.025149f
C356 VTAIL.n261 B 0.025149f
C357 VTAIL.n262 B 0.025149f
C358 VTAIL.n263 B 0.010953f
C359 VTAIL.n264 B 0.01064f
C360 VTAIL.n265 B 0.0198f
C361 VTAIL.n266 B 0.0198f
C362 VTAIL.n267 B 0.01064f
C363 VTAIL.n268 B 0.011266f
C364 VTAIL.n269 B 0.025149f
C365 VTAIL.n270 B 0.052553f
C366 VTAIL.n271 B 0.011266f
C367 VTAIL.n272 B 0.01064f
C368 VTAIL.n273 B 0.04685f
C369 VTAIL.n274 B 0.029244f
C370 VTAIL.n275 B 0.14705f
C371 VTAIL.n276 B 0.026763f
C372 VTAIL.n277 B 0.0198f
C373 VTAIL.n278 B 0.01064f
C374 VTAIL.n279 B 0.025149f
C375 VTAIL.n280 B 0.011266f
C376 VTAIL.n281 B 0.0198f
C377 VTAIL.n282 B 0.010953f
C378 VTAIL.n283 B 0.025149f
C379 VTAIL.n284 B 0.01064f
C380 VTAIL.n285 B 0.011266f
C381 VTAIL.n286 B 0.0198f
C382 VTAIL.n287 B 0.01064f
C383 VTAIL.n288 B 0.025149f
C384 VTAIL.n289 B 0.011266f
C385 VTAIL.n290 B 0.0198f
C386 VTAIL.n291 B 0.01064f
C387 VTAIL.n292 B 0.018862f
C388 VTAIL.n293 B 0.017778f
C389 VTAIL.t7 B 0.042263f
C390 VTAIL.n294 B 0.127558f
C391 VTAIL.n295 B 0.822753f
C392 VTAIL.n296 B 0.01064f
C393 VTAIL.n297 B 0.011266f
C394 VTAIL.n298 B 0.025149f
C395 VTAIL.n299 B 0.025149f
C396 VTAIL.n300 B 0.011266f
C397 VTAIL.n301 B 0.01064f
C398 VTAIL.n302 B 0.0198f
C399 VTAIL.n303 B 0.0198f
C400 VTAIL.n304 B 0.01064f
C401 VTAIL.n305 B 0.011266f
C402 VTAIL.n306 B 0.025149f
C403 VTAIL.n307 B 0.025149f
C404 VTAIL.n308 B 0.011266f
C405 VTAIL.n309 B 0.01064f
C406 VTAIL.n310 B 0.0198f
C407 VTAIL.n311 B 0.0198f
C408 VTAIL.n312 B 0.01064f
C409 VTAIL.n313 B 0.011266f
C410 VTAIL.n314 B 0.025149f
C411 VTAIL.n315 B 0.025149f
C412 VTAIL.n316 B 0.025149f
C413 VTAIL.n317 B 0.010953f
C414 VTAIL.n318 B 0.01064f
C415 VTAIL.n319 B 0.0198f
C416 VTAIL.n320 B 0.0198f
C417 VTAIL.n321 B 0.01064f
C418 VTAIL.n322 B 0.011266f
C419 VTAIL.n323 B 0.025149f
C420 VTAIL.n324 B 0.052553f
C421 VTAIL.n325 B 0.011266f
C422 VTAIL.n326 B 0.01064f
C423 VTAIL.n327 B 0.04685f
C424 VTAIL.n328 B 0.029244f
C425 VTAIL.n329 B 0.14705f
C426 VTAIL.t1 B 0.156469f
C427 VTAIL.t4 B 0.156469f
C428 VTAIL.n330 B 1.32216f
C429 VTAIL.n331 B 0.389242f
C430 VTAIL.n332 B 0.026763f
C431 VTAIL.n333 B 0.0198f
C432 VTAIL.n334 B 0.01064f
C433 VTAIL.n335 B 0.025149f
C434 VTAIL.n336 B 0.011266f
C435 VTAIL.n337 B 0.0198f
C436 VTAIL.n338 B 0.010953f
C437 VTAIL.n339 B 0.025149f
C438 VTAIL.n340 B 0.01064f
C439 VTAIL.n341 B 0.011266f
C440 VTAIL.n342 B 0.0198f
C441 VTAIL.n343 B 0.01064f
C442 VTAIL.n344 B 0.025149f
C443 VTAIL.n345 B 0.011266f
C444 VTAIL.n346 B 0.0198f
C445 VTAIL.n347 B 0.01064f
C446 VTAIL.n348 B 0.018862f
C447 VTAIL.n349 B 0.017778f
C448 VTAIL.t6 B 0.042263f
C449 VTAIL.n350 B 0.127558f
C450 VTAIL.n351 B 0.822753f
C451 VTAIL.n352 B 0.01064f
C452 VTAIL.n353 B 0.011266f
C453 VTAIL.n354 B 0.025149f
C454 VTAIL.n355 B 0.025149f
C455 VTAIL.n356 B 0.011266f
C456 VTAIL.n357 B 0.01064f
C457 VTAIL.n358 B 0.0198f
C458 VTAIL.n359 B 0.0198f
C459 VTAIL.n360 B 0.01064f
C460 VTAIL.n361 B 0.011266f
C461 VTAIL.n362 B 0.025149f
C462 VTAIL.n363 B 0.025149f
C463 VTAIL.n364 B 0.011266f
C464 VTAIL.n365 B 0.01064f
C465 VTAIL.n366 B 0.0198f
C466 VTAIL.n367 B 0.0198f
C467 VTAIL.n368 B 0.01064f
C468 VTAIL.n369 B 0.011266f
C469 VTAIL.n370 B 0.025149f
C470 VTAIL.n371 B 0.025149f
C471 VTAIL.n372 B 0.025149f
C472 VTAIL.n373 B 0.010953f
C473 VTAIL.n374 B 0.01064f
C474 VTAIL.n375 B 0.0198f
C475 VTAIL.n376 B 0.0198f
C476 VTAIL.n377 B 0.01064f
C477 VTAIL.n378 B 0.011266f
C478 VTAIL.n379 B 0.025149f
C479 VTAIL.n380 B 0.052553f
C480 VTAIL.n381 B 0.011266f
C481 VTAIL.n382 B 0.01064f
C482 VTAIL.n383 B 0.04685f
C483 VTAIL.n384 B 0.029244f
C484 VTAIL.n385 B 1.0356f
C485 VTAIL.n386 B 0.026763f
C486 VTAIL.n387 B 0.0198f
C487 VTAIL.n388 B 0.01064f
C488 VTAIL.n389 B 0.025149f
C489 VTAIL.n390 B 0.011266f
C490 VTAIL.n391 B 0.0198f
C491 VTAIL.n392 B 0.010953f
C492 VTAIL.n393 B 0.025149f
C493 VTAIL.n394 B 0.011266f
C494 VTAIL.n395 B 0.0198f
C495 VTAIL.n396 B 0.01064f
C496 VTAIL.n397 B 0.025149f
C497 VTAIL.n398 B 0.011266f
C498 VTAIL.n399 B 0.0198f
C499 VTAIL.n400 B 0.01064f
C500 VTAIL.n401 B 0.018862f
C501 VTAIL.n402 B 0.017778f
C502 VTAIL.t9 B 0.042263f
C503 VTAIL.n403 B 0.127558f
C504 VTAIL.n404 B 0.822753f
C505 VTAIL.n405 B 0.01064f
C506 VTAIL.n406 B 0.011266f
C507 VTAIL.n407 B 0.025149f
C508 VTAIL.n408 B 0.025149f
C509 VTAIL.n409 B 0.011266f
C510 VTAIL.n410 B 0.01064f
C511 VTAIL.n411 B 0.0198f
C512 VTAIL.n412 B 0.0198f
C513 VTAIL.n413 B 0.01064f
C514 VTAIL.n414 B 0.011266f
C515 VTAIL.n415 B 0.025149f
C516 VTAIL.n416 B 0.025149f
C517 VTAIL.n417 B 0.011266f
C518 VTAIL.n418 B 0.01064f
C519 VTAIL.n419 B 0.0198f
C520 VTAIL.n420 B 0.0198f
C521 VTAIL.n421 B 0.01064f
C522 VTAIL.n422 B 0.01064f
C523 VTAIL.n423 B 0.011266f
C524 VTAIL.n424 B 0.025149f
C525 VTAIL.n425 B 0.025149f
C526 VTAIL.n426 B 0.025149f
C527 VTAIL.n427 B 0.010953f
C528 VTAIL.n428 B 0.01064f
C529 VTAIL.n429 B 0.0198f
C530 VTAIL.n430 B 0.0198f
C531 VTAIL.n431 B 0.01064f
C532 VTAIL.n432 B 0.011266f
C533 VTAIL.n433 B 0.025149f
C534 VTAIL.n434 B 0.052553f
C535 VTAIL.n435 B 0.011266f
C536 VTAIL.n436 B 0.01064f
C537 VTAIL.n437 B 0.04685f
C538 VTAIL.n438 B 0.029244f
C539 VTAIL.n439 B 1.03189f
C540 VDD2.t3 B 0.196482f
C541 VDD2.t7 B 0.196482f
C542 VDD2.n0 B 1.73518f
C543 VDD2.t5 B 0.196482f
C544 VDD2.t0 B 0.196482f
C545 VDD2.n1 B 1.73518f
C546 VDD2.n2 B 2.48576f
C547 VDD2.t6 B 0.196482f
C548 VDD2.t1 B 0.196482f
C549 VDD2.n3 B 1.73071f
C550 VDD2.n4 B 2.39061f
C551 VDD2.t2 B 0.196482f
C552 VDD2.t4 B 0.196482f
C553 VDD2.n5 B 1.73515f
C554 VN.n0 B 0.031491f
C555 VN.t6 B 1.2626f
C556 VN.n1 B 0.051005f
C557 VN.n2 B 0.031491f
C558 VN.t7 B 1.2626f
C559 VN.n3 B 0.056781f
C560 VN.t2 B 1.36377f
C561 VN.t1 B 1.2626f
C562 VN.n4 B 0.531086f
C563 VN.n5 B 0.5322f
C564 VN.n6 B 0.19907f
C565 VN.n7 B 0.031491f
C566 VN.n8 B 0.025434f
C567 VN.n9 B 0.056781f
C568 VN.n10 B 0.464209f
C569 VN.n11 B 0.035046f
C570 VN.n12 B 0.031491f
C571 VN.n13 B 0.031491f
C572 VN.n14 B 0.031491f
C573 VN.n15 B 0.040549f
C574 VN.n16 B 0.041965f
C575 VN.n17 B 0.528282f
C576 VN.n18 B 0.029972f
C577 VN.n19 B 0.031491f
C578 VN.t0 B 1.2626f
C579 VN.n20 B 0.051005f
C580 VN.n21 B 0.031491f
C581 VN.t4 B 1.2626f
C582 VN.n22 B 0.056781f
C583 VN.t3 B 1.36377f
C584 VN.t5 B 1.2626f
C585 VN.n23 B 0.531086f
C586 VN.n24 B 0.5322f
C587 VN.n25 B 0.19907f
C588 VN.n26 B 0.031491f
C589 VN.n27 B 0.025434f
C590 VN.n28 B 0.056781f
C591 VN.n29 B 0.464209f
C592 VN.n30 B 0.035046f
C593 VN.n31 B 0.031491f
C594 VN.n32 B 0.031491f
C595 VN.n33 B 0.031491f
C596 VN.n34 B 0.040549f
C597 VN.n35 B 0.041965f
C598 VN.n36 B 0.528282f
C599 VN.n37 B 1.43267f
.ends

