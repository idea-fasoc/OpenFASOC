* NGSPICE file created from diff_pair_sample_0122.ext - technology: sky130A

.subckt diff_pair_sample_0122 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=5.4054 ps=28.5 w=13.86 l=2.25
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=0 ps=0 w=13.86 l=2.25
X2 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=5.4054 ps=28.5 w=13.86 l=2.25
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=0 ps=0 w=13.86 l=2.25
X4 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=5.4054 ps=28.5 w=13.86 l=2.25
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=0 ps=0 w=13.86 l=2.25
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=0 ps=0 w=13.86 l=2.25
X7 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4054 pd=28.5 as=5.4054 ps=28.5 w=13.86 l=2.25
R0 VP.n0 VP.t0 242.809
R1 VP.n0 VP.t1 197.672
R2 VP VP.n0 0.336784
R3 VTAIL.n2 VTAIL.t1 45.0744
R4 VTAIL.n1 VTAIL.t3 45.0744
R5 VTAIL.n3 VTAIL.t2 45.0743
R6 VTAIL.n0 VTAIL.t0 45.0743
R7 VTAIL.n1 VTAIL.n0 28.7634
R8 VTAIL.n3 VTAIL.n2 26.5393
R9 VTAIL.n2 VTAIL.n1 1.5824
R10 VTAIL VTAIL.n0 1.08455
R11 VTAIL VTAIL.n3 0.498345
R12 VDD1 VDD1.t0 102.889
R13 VDD1 VDD1.t1 62.3675
R14 B.n717 B.n716 585
R15 B.n306 B.n98 585
R16 B.n305 B.n304 585
R17 B.n303 B.n302 585
R18 B.n301 B.n300 585
R19 B.n299 B.n298 585
R20 B.n297 B.n296 585
R21 B.n295 B.n294 585
R22 B.n293 B.n292 585
R23 B.n291 B.n290 585
R24 B.n289 B.n288 585
R25 B.n287 B.n286 585
R26 B.n285 B.n284 585
R27 B.n283 B.n282 585
R28 B.n281 B.n280 585
R29 B.n279 B.n278 585
R30 B.n277 B.n276 585
R31 B.n275 B.n274 585
R32 B.n273 B.n272 585
R33 B.n271 B.n270 585
R34 B.n269 B.n268 585
R35 B.n267 B.n266 585
R36 B.n265 B.n264 585
R37 B.n263 B.n262 585
R38 B.n261 B.n260 585
R39 B.n259 B.n258 585
R40 B.n257 B.n256 585
R41 B.n255 B.n254 585
R42 B.n253 B.n252 585
R43 B.n251 B.n250 585
R44 B.n249 B.n248 585
R45 B.n247 B.n246 585
R46 B.n245 B.n244 585
R47 B.n243 B.n242 585
R48 B.n241 B.n240 585
R49 B.n239 B.n238 585
R50 B.n237 B.n236 585
R51 B.n235 B.n234 585
R52 B.n233 B.n232 585
R53 B.n231 B.n230 585
R54 B.n229 B.n228 585
R55 B.n227 B.n226 585
R56 B.n225 B.n224 585
R57 B.n223 B.n222 585
R58 B.n221 B.n220 585
R59 B.n219 B.n218 585
R60 B.n217 B.n216 585
R61 B.n214 B.n213 585
R62 B.n212 B.n211 585
R63 B.n210 B.n209 585
R64 B.n208 B.n207 585
R65 B.n206 B.n205 585
R66 B.n204 B.n203 585
R67 B.n202 B.n201 585
R68 B.n200 B.n199 585
R69 B.n198 B.n197 585
R70 B.n196 B.n195 585
R71 B.n193 B.n192 585
R72 B.n191 B.n190 585
R73 B.n189 B.n188 585
R74 B.n187 B.n186 585
R75 B.n185 B.n184 585
R76 B.n183 B.n182 585
R77 B.n181 B.n180 585
R78 B.n179 B.n178 585
R79 B.n177 B.n176 585
R80 B.n175 B.n174 585
R81 B.n173 B.n172 585
R82 B.n171 B.n170 585
R83 B.n169 B.n168 585
R84 B.n167 B.n166 585
R85 B.n165 B.n164 585
R86 B.n163 B.n162 585
R87 B.n161 B.n160 585
R88 B.n159 B.n158 585
R89 B.n157 B.n156 585
R90 B.n155 B.n154 585
R91 B.n153 B.n152 585
R92 B.n151 B.n150 585
R93 B.n149 B.n148 585
R94 B.n147 B.n146 585
R95 B.n145 B.n144 585
R96 B.n143 B.n142 585
R97 B.n141 B.n140 585
R98 B.n139 B.n138 585
R99 B.n137 B.n136 585
R100 B.n135 B.n134 585
R101 B.n133 B.n132 585
R102 B.n131 B.n130 585
R103 B.n129 B.n128 585
R104 B.n127 B.n126 585
R105 B.n125 B.n124 585
R106 B.n123 B.n122 585
R107 B.n121 B.n120 585
R108 B.n119 B.n118 585
R109 B.n117 B.n116 585
R110 B.n115 B.n114 585
R111 B.n113 B.n112 585
R112 B.n111 B.n110 585
R113 B.n109 B.n108 585
R114 B.n107 B.n106 585
R115 B.n105 B.n104 585
R116 B.n47 B.n46 585
R117 B.n722 B.n721 585
R118 B.n715 B.n99 585
R119 B.n99 B.n44 585
R120 B.n714 B.n43 585
R121 B.n726 B.n43 585
R122 B.n713 B.n42 585
R123 B.n727 B.n42 585
R124 B.n712 B.n41 585
R125 B.n728 B.n41 585
R126 B.n711 B.n710 585
R127 B.n710 B.n37 585
R128 B.n709 B.n36 585
R129 B.n734 B.n36 585
R130 B.n708 B.n35 585
R131 B.n735 B.n35 585
R132 B.n707 B.n34 585
R133 B.n736 B.n34 585
R134 B.n706 B.n705 585
R135 B.n705 B.n30 585
R136 B.n704 B.n29 585
R137 B.n742 B.n29 585
R138 B.n703 B.n28 585
R139 B.n743 B.n28 585
R140 B.n702 B.n27 585
R141 B.n744 B.n27 585
R142 B.n701 B.n700 585
R143 B.n700 B.n23 585
R144 B.n699 B.n22 585
R145 B.n750 B.n22 585
R146 B.n698 B.n21 585
R147 B.n751 B.n21 585
R148 B.n697 B.n20 585
R149 B.n752 B.n20 585
R150 B.n696 B.n695 585
R151 B.n695 B.n16 585
R152 B.n694 B.n15 585
R153 B.n758 B.n15 585
R154 B.n693 B.n14 585
R155 B.n759 B.n14 585
R156 B.n692 B.n13 585
R157 B.n760 B.n13 585
R158 B.n691 B.n690 585
R159 B.n690 B.n12 585
R160 B.n689 B.n688 585
R161 B.n689 B.n8 585
R162 B.n687 B.n7 585
R163 B.n767 B.n7 585
R164 B.n686 B.n6 585
R165 B.n768 B.n6 585
R166 B.n685 B.n5 585
R167 B.n769 B.n5 585
R168 B.n684 B.n683 585
R169 B.n683 B.n4 585
R170 B.n682 B.n307 585
R171 B.n682 B.n681 585
R172 B.n672 B.n308 585
R173 B.n309 B.n308 585
R174 B.n674 B.n673 585
R175 B.n675 B.n674 585
R176 B.n671 B.n313 585
R177 B.n317 B.n313 585
R178 B.n670 B.n669 585
R179 B.n669 B.n668 585
R180 B.n315 B.n314 585
R181 B.n316 B.n315 585
R182 B.n661 B.n660 585
R183 B.n662 B.n661 585
R184 B.n659 B.n322 585
R185 B.n322 B.n321 585
R186 B.n658 B.n657 585
R187 B.n657 B.n656 585
R188 B.n324 B.n323 585
R189 B.n325 B.n324 585
R190 B.n649 B.n648 585
R191 B.n650 B.n649 585
R192 B.n647 B.n330 585
R193 B.n330 B.n329 585
R194 B.n646 B.n645 585
R195 B.n645 B.n644 585
R196 B.n332 B.n331 585
R197 B.n333 B.n332 585
R198 B.n637 B.n636 585
R199 B.n638 B.n637 585
R200 B.n635 B.n338 585
R201 B.n338 B.n337 585
R202 B.n634 B.n633 585
R203 B.n633 B.n632 585
R204 B.n340 B.n339 585
R205 B.n341 B.n340 585
R206 B.n625 B.n624 585
R207 B.n626 B.n625 585
R208 B.n623 B.n346 585
R209 B.n346 B.n345 585
R210 B.n622 B.n621 585
R211 B.n621 B.n620 585
R212 B.n348 B.n347 585
R213 B.n349 B.n348 585
R214 B.n616 B.n615 585
R215 B.n352 B.n351 585
R216 B.n612 B.n611 585
R217 B.n613 B.n612 585
R218 B.n610 B.n404 585
R219 B.n609 B.n608 585
R220 B.n607 B.n606 585
R221 B.n605 B.n604 585
R222 B.n603 B.n602 585
R223 B.n601 B.n600 585
R224 B.n599 B.n598 585
R225 B.n597 B.n596 585
R226 B.n595 B.n594 585
R227 B.n593 B.n592 585
R228 B.n591 B.n590 585
R229 B.n589 B.n588 585
R230 B.n587 B.n586 585
R231 B.n585 B.n584 585
R232 B.n583 B.n582 585
R233 B.n581 B.n580 585
R234 B.n579 B.n578 585
R235 B.n577 B.n576 585
R236 B.n575 B.n574 585
R237 B.n573 B.n572 585
R238 B.n571 B.n570 585
R239 B.n569 B.n568 585
R240 B.n567 B.n566 585
R241 B.n565 B.n564 585
R242 B.n563 B.n562 585
R243 B.n561 B.n560 585
R244 B.n559 B.n558 585
R245 B.n557 B.n556 585
R246 B.n555 B.n554 585
R247 B.n553 B.n552 585
R248 B.n551 B.n550 585
R249 B.n549 B.n548 585
R250 B.n547 B.n546 585
R251 B.n545 B.n544 585
R252 B.n543 B.n542 585
R253 B.n541 B.n540 585
R254 B.n539 B.n538 585
R255 B.n537 B.n536 585
R256 B.n535 B.n534 585
R257 B.n533 B.n532 585
R258 B.n531 B.n530 585
R259 B.n529 B.n528 585
R260 B.n527 B.n526 585
R261 B.n525 B.n524 585
R262 B.n523 B.n522 585
R263 B.n521 B.n520 585
R264 B.n519 B.n518 585
R265 B.n517 B.n516 585
R266 B.n515 B.n514 585
R267 B.n513 B.n512 585
R268 B.n511 B.n510 585
R269 B.n509 B.n508 585
R270 B.n507 B.n506 585
R271 B.n505 B.n504 585
R272 B.n503 B.n502 585
R273 B.n501 B.n500 585
R274 B.n499 B.n498 585
R275 B.n497 B.n496 585
R276 B.n495 B.n494 585
R277 B.n493 B.n492 585
R278 B.n491 B.n490 585
R279 B.n489 B.n488 585
R280 B.n487 B.n486 585
R281 B.n485 B.n484 585
R282 B.n483 B.n482 585
R283 B.n481 B.n480 585
R284 B.n479 B.n478 585
R285 B.n477 B.n476 585
R286 B.n475 B.n474 585
R287 B.n473 B.n472 585
R288 B.n471 B.n470 585
R289 B.n469 B.n468 585
R290 B.n467 B.n466 585
R291 B.n465 B.n464 585
R292 B.n463 B.n462 585
R293 B.n461 B.n460 585
R294 B.n459 B.n458 585
R295 B.n457 B.n456 585
R296 B.n455 B.n454 585
R297 B.n453 B.n452 585
R298 B.n451 B.n450 585
R299 B.n449 B.n448 585
R300 B.n447 B.n446 585
R301 B.n445 B.n444 585
R302 B.n443 B.n442 585
R303 B.n441 B.n440 585
R304 B.n439 B.n438 585
R305 B.n437 B.n436 585
R306 B.n435 B.n434 585
R307 B.n433 B.n432 585
R308 B.n431 B.n430 585
R309 B.n429 B.n428 585
R310 B.n427 B.n426 585
R311 B.n425 B.n424 585
R312 B.n423 B.n422 585
R313 B.n421 B.n420 585
R314 B.n419 B.n418 585
R315 B.n417 B.n416 585
R316 B.n415 B.n414 585
R317 B.n413 B.n412 585
R318 B.n411 B.n403 585
R319 B.n613 B.n403 585
R320 B.n617 B.n350 585
R321 B.n350 B.n349 585
R322 B.n619 B.n618 585
R323 B.n620 B.n619 585
R324 B.n344 B.n343 585
R325 B.n345 B.n344 585
R326 B.n628 B.n627 585
R327 B.n627 B.n626 585
R328 B.n629 B.n342 585
R329 B.n342 B.n341 585
R330 B.n631 B.n630 585
R331 B.n632 B.n631 585
R332 B.n336 B.n335 585
R333 B.n337 B.n336 585
R334 B.n640 B.n639 585
R335 B.n639 B.n638 585
R336 B.n641 B.n334 585
R337 B.n334 B.n333 585
R338 B.n643 B.n642 585
R339 B.n644 B.n643 585
R340 B.n328 B.n327 585
R341 B.n329 B.n328 585
R342 B.n652 B.n651 585
R343 B.n651 B.n650 585
R344 B.n653 B.n326 585
R345 B.n326 B.n325 585
R346 B.n655 B.n654 585
R347 B.n656 B.n655 585
R348 B.n320 B.n319 585
R349 B.n321 B.n320 585
R350 B.n664 B.n663 585
R351 B.n663 B.n662 585
R352 B.n665 B.n318 585
R353 B.n318 B.n316 585
R354 B.n667 B.n666 585
R355 B.n668 B.n667 585
R356 B.n312 B.n311 585
R357 B.n317 B.n312 585
R358 B.n677 B.n676 585
R359 B.n676 B.n675 585
R360 B.n678 B.n310 585
R361 B.n310 B.n309 585
R362 B.n680 B.n679 585
R363 B.n681 B.n680 585
R364 B.n3 B.n0 585
R365 B.n4 B.n3 585
R366 B.n766 B.n1 585
R367 B.n767 B.n766 585
R368 B.n765 B.n764 585
R369 B.n765 B.n8 585
R370 B.n763 B.n9 585
R371 B.n12 B.n9 585
R372 B.n762 B.n761 585
R373 B.n761 B.n760 585
R374 B.n11 B.n10 585
R375 B.n759 B.n11 585
R376 B.n757 B.n756 585
R377 B.n758 B.n757 585
R378 B.n755 B.n17 585
R379 B.n17 B.n16 585
R380 B.n754 B.n753 585
R381 B.n753 B.n752 585
R382 B.n19 B.n18 585
R383 B.n751 B.n19 585
R384 B.n749 B.n748 585
R385 B.n750 B.n749 585
R386 B.n747 B.n24 585
R387 B.n24 B.n23 585
R388 B.n746 B.n745 585
R389 B.n745 B.n744 585
R390 B.n26 B.n25 585
R391 B.n743 B.n26 585
R392 B.n741 B.n740 585
R393 B.n742 B.n741 585
R394 B.n739 B.n31 585
R395 B.n31 B.n30 585
R396 B.n738 B.n737 585
R397 B.n737 B.n736 585
R398 B.n33 B.n32 585
R399 B.n735 B.n33 585
R400 B.n733 B.n732 585
R401 B.n734 B.n733 585
R402 B.n731 B.n38 585
R403 B.n38 B.n37 585
R404 B.n730 B.n729 585
R405 B.n729 B.n728 585
R406 B.n40 B.n39 585
R407 B.n727 B.n40 585
R408 B.n725 B.n724 585
R409 B.n726 B.n725 585
R410 B.n723 B.n45 585
R411 B.n45 B.n44 585
R412 B.n770 B.n769 585
R413 B.n768 B.n2 585
R414 B.n721 B.n45 444.452
R415 B.n717 B.n99 444.452
R416 B.n403 B.n348 444.452
R417 B.n615 B.n350 444.452
R418 B.n102 B.t13 355.906
R419 B.n100 B.t6 355.906
R420 B.n408 B.t2 355.906
R421 B.n405 B.t10 355.906
R422 B.n719 B.n718 256.663
R423 B.n719 B.n97 256.663
R424 B.n719 B.n96 256.663
R425 B.n719 B.n95 256.663
R426 B.n719 B.n94 256.663
R427 B.n719 B.n93 256.663
R428 B.n719 B.n92 256.663
R429 B.n719 B.n91 256.663
R430 B.n719 B.n90 256.663
R431 B.n719 B.n89 256.663
R432 B.n719 B.n88 256.663
R433 B.n719 B.n87 256.663
R434 B.n719 B.n86 256.663
R435 B.n719 B.n85 256.663
R436 B.n719 B.n84 256.663
R437 B.n719 B.n83 256.663
R438 B.n719 B.n82 256.663
R439 B.n719 B.n81 256.663
R440 B.n719 B.n80 256.663
R441 B.n719 B.n79 256.663
R442 B.n719 B.n78 256.663
R443 B.n719 B.n77 256.663
R444 B.n719 B.n76 256.663
R445 B.n719 B.n75 256.663
R446 B.n719 B.n74 256.663
R447 B.n719 B.n73 256.663
R448 B.n719 B.n72 256.663
R449 B.n719 B.n71 256.663
R450 B.n719 B.n70 256.663
R451 B.n719 B.n69 256.663
R452 B.n719 B.n68 256.663
R453 B.n719 B.n67 256.663
R454 B.n719 B.n66 256.663
R455 B.n719 B.n65 256.663
R456 B.n719 B.n64 256.663
R457 B.n719 B.n63 256.663
R458 B.n719 B.n62 256.663
R459 B.n719 B.n61 256.663
R460 B.n719 B.n60 256.663
R461 B.n719 B.n59 256.663
R462 B.n719 B.n58 256.663
R463 B.n719 B.n57 256.663
R464 B.n719 B.n56 256.663
R465 B.n719 B.n55 256.663
R466 B.n719 B.n54 256.663
R467 B.n719 B.n53 256.663
R468 B.n719 B.n52 256.663
R469 B.n719 B.n51 256.663
R470 B.n719 B.n50 256.663
R471 B.n719 B.n49 256.663
R472 B.n719 B.n48 256.663
R473 B.n720 B.n719 256.663
R474 B.n614 B.n613 256.663
R475 B.n613 B.n353 256.663
R476 B.n613 B.n354 256.663
R477 B.n613 B.n355 256.663
R478 B.n613 B.n356 256.663
R479 B.n613 B.n357 256.663
R480 B.n613 B.n358 256.663
R481 B.n613 B.n359 256.663
R482 B.n613 B.n360 256.663
R483 B.n613 B.n361 256.663
R484 B.n613 B.n362 256.663
R485 B.n613 B.n363 256.663
R486 B.n613 B.n364 256.663
R487 B.n613 B.n365 256.663
R488 B.n613 B.n366 256.663
R489 B.n613 B.n367 256.663
R490 B.n613 B.n368 256.663
R491 B.n613 B.n369 256.663
R492 B.n613 B.n370 256.663
R493 B.n613 B.n371 256.663
R494 B.n613 B.n372 256.663
R495 B.n613 B.n373 256.663
R496 B.n613 B.n374 256.663
R497 B.n613 B.n375 256.663
R498 B.n613 B.n376 256.663
R499 B.n613 B.n377 256.663
R500 B.n613 B.n378 256.663
R501 B.n613 B.n379 256.663
R502 B.n613 B.n380 256.663
R503 B.n613 B.n381 256.663
R504 B.n613 B.n382 256.663
R505 B.n613 B.n383 256.663
R506 B.n613 B.n384 256.663
R507 B.n613 B.n385 256.663
R508 B.n613 B.n386 256.663
R509 B.n613 B.n387 256.663
R510 B.n613 B.n388 256.663
R511 B.n613 B.n389 256.663
R512 B.n613 B.n390 256.663
R513 B.n613 B.n391 256.663
R514 B.n613 B.n392 256.663
R515 B.n613 B.n393 256.663
R516 B.n613 B.n394 256.663
R517 B.n613 B.n395 256.663
R518 B.n613 B.n396 256.663
R519 B.n613 B.n397 256.663
R520 B.n613 B.n398 256.663
R521 B.n613 B.n399 256.663
R522 B.n613 B.n400 256.663
R523 B.n613 B.n401 256.663
R524 B.n613 B.n402 256.663
R525 B.n772 B.n771 256.663
R526 B.n104 B.n47 163.367
R527 B.n108 B.n107 163.367
R528 B.n112 B.n111 163.367
R529 B.n116 B.n115 163.367
R530 B.n120 B.n119 163.367
R531 B.n124 B.n123 163.367
R532 B.n128 B.n127 163.367
R533 B.n132 B.n131 163.367
R534 B.n136 B.n135 163.367
R535 B.n140 B.n139 163.367
R536 B.n144 B.n143 163.367
R537 B.n148 B.n147 163.367
R538 B.n152 B.n151 163.367
R539 B.n156 B.n155 163.367
R540 B.n160 B.n159 163.367
R541 B.n164 B.n163 163.367
R542 B.n168 B.n167 163.367
R543 B.n172 B.n171 163.367
R544 B.n176 B.n175 163.367
R545 B.n180 B.n179 163.367
R546 B.n184 B.n183 163.367
R547 B.n188 B.n187 163.367
R548 B.n192 B.n191 163.367
R549 B.n197 B.n196 163.367
R550 B.n201 B.n200 163.367
R551 B.n205 B.n204 163.367
R552 B.n209 B.n208 163.367
R553 B.n213 B.n212 163.367
R554 B.n218 B.n217 163.367
R555 B.n222 B.n221 163.367
R556 B.n226 B.n225 163.367
R557 B.n230 B.n229 163.367
R558 B.n234 B.n233 163.367
R559 B.n238 B.n237 163.367
R560 B.n242 B.n241 163.367
R561 B.n246 B.n245 163.367
R562 B.n250 B.n249 163.367
R563 B.n254 B.n253 163.367
R564 B.n258 B.n257 163.367
R565 B.n262 B.n261 163.367
R566 B.n266 B.n265 163.367
R567 B.n270 B.n269 163.367
R568 B.n274 B.n273 163.367
R569 B.n278 B.n277 163.367
R570 B.n282 B.n281 163.367
R571 B.n286 B.n285 163.367
R572 B.n290 B.n289 163.367
R573 B.n294 B.n293 163.367
R574 B.n298 B.n297 163.367
R575 B.n302 B.n301 163.367
R576 B.n304 B.n98 163.367
R577 B.n621 B.n348 163.367
R578 B.n621 B.n346 163.367
R579 B.n625 B.n346 163.367
R580 B.n625 B.n340 163.367
R581 B.n633 B.n340 163.367
R582 B.n633 B.n338 163.367
R583 B.n637 B.n338 163.367
R584 B.n637 B.n332 163.367
R585 B.n645 B.n332 163.367
R586 B.n645 B.n330 163.367
R587 B.n649 B.n330 163.367
R588 B.n649 B.n324 163.367
R589 B.n657 B.n324 163.367
R590 B.n657 B.n322 163.367
R591 B.n661 B.n322 163.367
R592 B.n661 B.n315 163.367
R593 B.n669 B.n315 163.367
R594 B.n669 B.n313 163.367
R595 B.n674 B.n313 163.367
R596 B.n674 B.n308 163.367
R597 B.n682 B.n308 163.367
R598 B.n683 B.n682 163.367
R599 B.n683 B.n5 163.367
R600 B.n6 B.n5 163.367
R601 B.n7 B.n6 163.367
R602 B.n689 B.n7 163.367
R603 B.n690 B.n689 163.367
R604 B.n690 B.n13 163.367
R605 B.n14 B.n13 163.367
R606 B.n15 B.n14 163.367
R607 B.n695 B.n15 163.367
R608 B.n695 B.n20 163.367
R609 B.n21 B.n20 163.367
R610 B.n22 B.n21 163.367
R611 B.n700 B.n22 163.367
R612 B.n700 B.n27 163.367
R613 B.n28 B.n27 163.367
R614 B.n29 B.n28 163.367
R615 B.n705 B.n29 163.367
R616 B.n705 B.n34 163.367
R617 B.n35 B.n34 163.367
R618 B.n36 B.n35 163.367
R619 B.n710 B.n36 163.367
R620 B.n710 B.n41 163.367
R621 B.n42 B.n41 163.367
R622 B.n43 B.n42 163.367
R623 B.n99 B.n43 163.367
R624 B.n612 B.n352 163.367
R625 B.n612 B.n404 163.367
R626 B.n608 B.n607 163.367
R627 B.n604 B.n603 163.367
R628 B.n600 B.n599 163.367
R629 B.n596 B.n595 163.367
R630 B.n592 B.n591 163.367
R631 B.n588 B.n587 163.367
R632 B.n584 B.n583 163.367
R633 B.n580 B.n579 163.367
R634 B.n576 B.n575 163.367
R635 B.n572 B.n571 163.367
R636 B.n568 B.n567 163.367
R637 B.n564 B.n563 163.367
R638 B.n560 B.n559 163.367
R639 B.n556 B.n555 163.367
R640 B.n552 B.n551 163.367
R641 B.n548 B.n547 163.367
R642 B.n544 B.n543 163.367
R643 B.n540 B.n539 163.367
R644 B.n536 B.n535 163.367
R645 B.n532 B.n531 163.367
R646 B.n528 B.n527 163.367
R647 B.n524 B.n523 163.367
R648 B.n520 B.n519 163.367
R649 B.n516 B.n515 163.367
R650 B.n512 B.n511 163.367
R651 B.n508 B.n507 163.367
R652 B.n504 B.n503 163.367
R653 B.n500 B.n499 163.367
R654 B.n496 B.n495 163.367
R655 B.n492 B.n491 163.367
R656 B.n488 B.n487 163.367
R657 B.n484 B.n483 163.367
R658 B.n480 B.n479 163.367
R659 B.n476 B.n475 163.367
R660 B.n472 B.n471 163.367
R661 B.n468 B.n467 163.367
R662 B.n464 B.n463 163.367
R663 B.n460 B.n459 163.367
R664 B.n456 B.n455 163.367
R665 B.n452 B.n451 163.367
R666 B.n448 B.n447 163.367
R667 B.n444 B.n443 163.367
R668 B.n440 B.n439 163.367
R669 B.n436 B.n435 163.367
R670 B.n432 B.n431 163.367
R671 B.n428 B.n427 163.367
R672 B.n424 B.n423 163.367
R673 B.n420 B.n419 163.367
R674 B.n416 B.n415 163.367
R675 B.n412 B.n403 163.367
R676 B.n619 B.n350 163.367
R677 B.n619 B.n344 163.367
R678 B.n627 B.n344 163.367
R679 B.n627 B.n342 163.367
R680 B.n631 B.n342 163.367
R681 B.n631 B.n336 163.367
R682 B.n639 B.n336 163.367
R683 B.n639 B.n334 163.367
R684 B.n643 B.n334 163.367
R685 B.n643 B.n328 163.367
R686 B.n651 B.n328 163.367
R687 B.n651 B.n326 163.367
R688 B.n655 B.n326 163.367
R689 B.n655 B.n320 163.367
R690 B.n663 B.n320 163.367
R691 B.n663 B.n318 163.367
R692 B.n667 B.n318 163.367
R693 B.n667 B.n312 163.367
R694 B.n676 B.n312 163.367
R695 B.n676 B.n310 163.367
R696 B.n680 B.n310 163.367
R697 B.n680 B.n3 163.367
R698 B.n770 B.n3 163.367
R699 B.n766 B.n2 163.367
R700 B.n766 B.n765 163.367
R701 B.n765 B.n9 163.367
R702 B.n761 B.n9 163.367
R703 B.n761 B.n11 163.367
R704 B.n757 B.n11 163.367
R705 B.n757 B.n17 163.367
R706 B.n753 B.n17 163.367
R707 B.n753 B.n19 163.367
R708 B.n749 B.n19 163.367
R709 B.n749 B.n24 163.367
R710 B.n745 B.n24 163.367
R711 B.n745 B.n26 163.367
R712 B.n741 B.n26 163.367
R713 B.n741 B.n31 163.367
R714 B.n737 B.n31 163.367
R715 B.n737 B.n33 163.367
R716 B.n733 B.n33 163.367
R717 B.n733 B.n38 163.367
R718 B.n729 B.n38 163.367
R719 B.n729 B.n40 163.367
R720 B.n725 B.n40 163.367
R721 B.n725 B.n45 163.367
R722 B.n100 B.t8 122.65
R723 B.n408 B.t5 122.65
R724 B.n102 B.t14 122.632
R725 B.n405 B.t12 122.632
R726 B.n101 B.t9 72.6134
R727 B.n409 B.t4 72.6134
R728 B.n103 B.t15 72.5957
R729 B.n406 B.t11 72.5957
R730 B.n721 B.n720 71.676
R731 B.n104 B.n48 71.676
R732 B.n108 B.n49 71.676
R733 B.n112 B.n50 71.676
R734 B.n116 B.n51 71.676
R735 B.n120 B.n52 71.676
R736 B.n124 B.n53 71.676
R737 B.n128 B.n54 71.676
R738 B.n132 B.n55 71.676
R739 B.n136 B.n56 71.676
R740 B.n140 B.n57 71.676
R741 B.n144 B.n58 71.676
R742 B.n148 B.n59 71.676
R743 B.n152 B.n60 71.676
R744 B.n156 B.n61 71.676
R745 B.n160 B.n62 71.676
R746 B.n164 B.n63 71.676
R747 B.n168 B.n64 71.676
R748 B.n172 B.n65 71.676
R749 B.n176 B.n66 71.676
R750 B.n180 B.n67 71.676
R751 B.n184 B.n68 71.676
R752 B.n188 B.n69 71.676
R753 B.n192 B.n70 71.676
R754 B.n197 B.n71 71.676
R755 B.n201 B.n72 71.676
R756 B.n205 B.n73 71.676
R757 B.n209 B.n74 71.676
R758 B.n213 B.n75 71.676
R759 B.n218 B.n76 71.676
R760 B.n222 B.n77 71.676
R761 B.n226 B.n78 71.676
R762 B.n230 B.n79 71.676
R763 B.n234 B.n80 71.676
R764 B.n238 B.n81 71.676
R765 B.n242 B.n82 71.676
R766 B.n246 B.n83 71.676
R767 B.n250 B.n84 71.676
R768 B.n254 B.n85 71.676
R769 B.n258 B.n86 71.676
R770 B.n262 B.n87 71.676
R771 B.n266 B.n88 71.676
R772 B.n270 B.n89 71.676
R773 B.n274 B.n90 71.676
R774 B.n278 B.n91 71.676
R775 B.n282 B.n92 71.676
R776 B.n286 B.n93 71.676
R777 B.n290 B.n94 71.676
R778 B.n294 B.n95 71.676
R779 B.n298 B.n96 71.676
R780 B.n302 B.n97 71.676
R781 B.n718 B.n98 71.676
R782 B.n718 B.n717 71.676
R783 B.n304 B.n97 71.676
R784 B.n301 B.n96 71.676
R785 B.n297 B.n95 71.676
R786 B.n293 B.n94 71.676
R787 B.n289 B.n93 71.676
R788 B.n285 B.n92 71.676
R789 B.n281 B.n91 71.676
R790 B.n277 B.n90 71.676
R791 B.n273 B.n89 71.676
R792 B.n269 B.n88 71.676
R793 B.n265 B.n87 71.676
R794 B.n261 B.n86 71.676
R795 B.n257 B.n85 71.676
R796 B.n253 B.n84 71.676
R797 B.n249 B.n83 71.676
R798 B.n245 B.n82 71.676
R799 B.n241 B.n81 71.676
R800 B.n237 B.n80 71.676
R801 B.n233 B.n79 71.676
R802 B.n229 B.n78 71.676
R803 B.n225 B.n77 71.676
R804 B.n221 B.n76 71.676
R805 B.n217 B.n75 71.676
R806 B.n212 B.n74 71.676
R807 B.n208 B.n73 71.676
R808 B.n204 B.n72 71.676
R809 B.n200 B.n71 71.676
R810 B.n196 B.n70 71.676
R811 B.n191 B.n69 71.676
R812 B.n187 B.n68 71.676
R813 B.n183 B.n67 71.676
R814 B.n179 B.n66 71.676
R815 B.n175 B.n65 71.676
R816 B.n171 B.n64 71.676
R817 B.n167 B.n63 71.676
R818 B.n163 B.n62 71.676
R819 B.n159 B.n61 71.676
R820 B.n155 B.n60 71.676
R821 B.n151 B.n59 71.676
R822 B.n147 B.n58 71.676
R823 B.n143 B.n57 71.676
R824 B.n139 B.n56 71.676
R825 B.n135 B.n55 71.676
R826 B.n131 B.n54 71.676
R827 B.n127 B.n53 71.676
R828 B.n123 B.n52 71.676
R829 B.n119 B.n51 71.676
R830 B.n115 B.n50 71.676
R831 B.n111 B.n49 71.676
R832 B.n107 B.n48 71.676
R833 B.n720 B.n47 71.676
R834 B.n615 B.n614 71.676
R835 B.n404 B.n353 71.676
R836 B.n607 B.n354 71.676
R837 B.n603 B.n355 71.676
R838 B.n599 B.n356 71.676
R839 B.n595 B.n357 71.676
R840 B.n591 B.n358 71.676
R841 B.n587 B.n359 71.676
R842 B.n583 B.n360 71.676
R843 B.n579 B.n361 71.676
R844 B.n575 B.n362 71.676
R845 B.n571 B.n363 71.676
R846 B.n567 B.n364 71.676
R847 B.n563 B.n365 71.676
R848 B.n559 B.n366 71.676
R849 B.n555 B.n367 71.676
R850 B.n551 B.n368 71.676
R851 B.n547 B.n369 71.676
R852 B.n543 B.n370 71.676
R853 B.n539 B.n371 71.676
R854 B.n535 B.n372 71.676
R855 B.n531 B.n373 71.676
R856 B.n527 B.n374 71.676
R857 B.n523 B.n375 71.676
R858 B.n519 B.n376 71.676
R859 B.n515 B.n377 71.676
R860 B.n511 B.n378 71.676
R861 B.n507 B.n379 71.676
R862 B.n503 B.n380 71.676
R863 B.n499 B.n381 71.676
R864 B.n495 B.n382 71.676
R865 B.n491 B.n383 71.676
R866 B.n487 B.n384 71.676
R867 B.n483 B.n385 71.676
R868 B.n479 B.n386 71.676
R869 B.n475 B.n387 71.676
R870 B.n471 B.n388 71.676
R871 B.n467 B.n389 71.676
R872 B.n463 B.n390 71.676
R873 B.n459 B.n391 71.676
R874 B.n455 B.n392 71.676
R875 B.n451 B.n393 71.676
R876 B.n447 B.n394 71.676
R877 B.n443 B.n395 71.676
R878 B.n439 B.n396 71.676
R879 B.n435 B.n397 71.676
R880 B.n431 B.n398 71.676
R881 B.n427 B.n399 71.676
R882 B.n423 B.n400 71.676
R883 B.n419 B.n401 71.676
R884 B.n415 B.n402 71.676
R885 B.n614 B.n352 71.676
R886 B.n608 B.n353 71.676
R887 B.n604 B.n354 71.676
R888 B.n600 B.n355 71.676
R889 B.n596 B.n356 71.676
R890 B.n592 B.n357 71.676
R891 B.n588 B.n358 71.676
R892 B.n584 B.n359 71.676
R893 B.n580 B.n360 71.676
R894 B.n576 B.n361 71.676
R895 B.n572 B.n362 71.676
R896 B.n568 B.n363 71.676
R897 B.n564 B.n364 71.676
R898 B.n560 B.n365 71.676
R899 B.n556 B.n366 71.676
R900 B.n552 B.n367 71.676
R901 B.n548 B.n368 71.676
R902 B.n544 B.n369 71.676
R903 B.n540 B.n370 71.676
R904 B.n536 B.n371 71.676
R905 B.n532 B.n372 71.676
R906 B.n528 B.n373 71.676
R907 B.n524 B.n374 71.676
R908 B.n520 B.n375 71.676
R909 B.n516 B.n376 71.676
R910 B.n512 B.n377 71.676
R911 B.n508 B.n378 71.676
R912 B.n504 B.n379 71.676
R913 B.n500 B.n380 71.676
R914 B.n496 B.n381 71.676
R915 B.n492 B.n382 71.676
R916 B.n488 B.n383 71.676
R917 B.n484 B.n384 71.676
R918 B.n480 B.n385 71.676
R919 B.n476 B.n386 71.676
R920 B.n472 B.n387 71.676
R921 B.n468 B.n388 71.676
R922 B.n464 B.n389 71.676
R923 B.n460 B.n390 71.676
R924 B.n456 B.n391 71.676
R925 B.n452 B.n392 71.676
R926 B.n448 B.n393 71.676
R927 B.n444 B.n394 71.676
R928 B.n440 B.n395 71.676
R929 B.n436 B.n396 71.676
R930 B.n432 B.n397 71.676
R931 B.n428 B.n398 71.676
R932 B.n424 B.n399 71.676
R933 B.n420 B.n400 71.676
R934 B.n416 B.n401 71.676
R935 B.n412 B.n402 71.676
R936 B.n771 B.n770 71.676
R937 B.n771 B.n2 71.676
R938 B.n613 B.n349 62.6605
R939 B.n719 B.n44 62.6605
R940 B.n194 B.n103 59.5399
R941 B.n215 B.n101 59.5399
R942 B.n410 B.n409 59.5399
R943 B.n407 B.n406 59.5399
R944 B.n103 B.n102 50.0369
R945 B.n101 B.n100 50.0369
R946 B.n409 B.n408 50.0369
R947 B.n406 B.n405 50.0369
R948 B.n620 B.n349 39.0912
R949 B.n620 B.n345 39.0912
R950 B.n626 B.n345 39.0912
R951 B.n626 B.n341 39.0912
R952 B.n632 B.n341 39.0912
R953 B.n632 B.n337 39.0912
R954 B.n638 B.n337 39.0912
R955 B.n644 B.n333 39.0912
R956 B.n644 B.n329 39.0912
R957 B.n650 B.n329 39.0912
R958 B.n650 B.n325 39.0912
R959 B.n656 B.n325 39.0912
R960 B.n656 B.n321 39.0912
R961 B.n662 B.n321 39.0912
R962 B.n662 B.n316 39.0912
R963 B.n668 B.n316 39.0912
R964 B.n668 B.n317 39.0912
R965 B.n675 B.n309 39.0912
R966 B.n681 B.n309 39.0912
R967 B.n681 B.n4 39.0912
R968 B.n769 B.n4 39.0912
R969 B.n769 B.n768 39.0912
R970 B.n768 B.n767 39.0912
R971 B.n767 B.n8 39.0912
R972 B.n12 B.n8 39.0912
R973 B.n760 B.n12 39.0912
R974 B.n759 B.n758 39.0912
R975 B.n758 B.n16 39.0912
R976 B.n752 B.n16 39.0912
R977 B.n752 B.n751 39.0912
R978 B.n751 B.n750 39.0912
R979 B.n750 B.n23 39.0912
R980 B.n744 B.n23 39.0912
R981 B.n744 B.n743 39.0912
R982 B.n743 B.n742 39.0912
R983 B.n742 B.n30 39.0912
R984 B.n736 B.n735 39.0912
R985 B.n735 B.n734 39.0912
R986 B.n734 B.n37 39.0912
R987 B.n728 B.n37 39.0912
R988 B.n728 B.n727 39.0912
R989 B.n727 B.n726 39.0912
R990 B.n726 B.n44 39.0912
R991 B.n675 B.t0 35.0671
R992 B.n760 B.t1 35.0671
R993 B.n617 B.n616 28.8785
R994 B.n411 B.n347 28.8785
R995 B.n723 B.n722 28.8785
R996 B.n716 B.n715 28.8785
R997 B.t3 B.n333 27.0191
R998 B.t7 B.n30 27.0191
R999 B B.n772 18.0485
R1000 B.n638 B.t3 12.0726
R1001 B.n736 B.t7 12.0726
R1002 B.n618 B.n617 10.6151
R1003 B.n618 B.n343 10.6151
R1004 B.n628 B.n343 10.6151
R1005 B.n629 B.n628 10.6151
R1006 B.n630 B.n629 10.6151
R1007 B.n630 B.n335 10.6151
R1008 B.n640 B.n335 10.6151
R1009 B.n641 B.n640 10.6151
R1010 B.n642 B.n641 10.6151
R1011 B.n642 B.n327 10.6151
R1012 B.n652 B.n327 10.6151
R1013 B.n653 B.n652 10.6151
R1014 B.n654 B.n653 10.6151
R1015 B.n654 B.n319 10.6151
R1016 B.n664 B.n319 10.6151
R1017 B.n665 B.n664 10.6151
R1018 B.n666 B.n665 10.6151
R1019 B.n666 B.n311 10.6151
R1020 B.n677 B.n311 10.6151
R1021 B.n678 B.n677 10.6151
R1022 B.n679 B.n678 10.6151
R1023 B.n679 B.n0 10.6151
R1024 B.n616 B.n351 10.6151
R1025 B.n611 B.n351 10.6151
R1026 B.n611 B.n610 10.6151
R1027 B.n610 B.n609 10.6151
R1028 B.n609 B.n606 10.6151
R1029 B.n606 B.n605 10.6151
R1030 B.n605 B.n602 10.6151
R1031 B.n602 B.n601 10.6151
R1032 B.n601 B.n598 10.6151
R1033 B.n598 B.n597 10.6151
R1034 B.n597 B.n594 10.6151
R1035 B.n594 B.n593 10.6151
R1036 B.n593 B.n590 10.6151
R1037 B.n590 B.n589 10.6151
R1038 B.n589 B.n586 10.6151
R1039 B.n586 B.n585 10.6151
R1040 B.n585 B.n582 10.6151
R1041 B.n582 B.n581 10.6151
R1042 B.n581 B.n578 10.6151
R1043 B.n578 B.n577 10.6151
R1044 B.n577 B.n574 10.6151
R1045 B.n574 B.n573 10.6151
R1046 B.n573 B.n570 10.6151
R1047 B.n570 B.n569 10.6151
R1048 B.n569 B.n566 10.6151
R1049 B.n566 B.n565 10.6151
R1050 B.n565 B.n562 10.6151
R1051 B.n562 B.n561 10.6151
R1052 B.n561 B.n558 10.6151
R1053 B.n558 B.n557 10.6151
R1054 B.n557 B.n554 10.6151
R1055 B.n554 B.n553 10.6151
R1056 B.n553 B.n550 10.6151
R1057 B.n550 B.n549 10.6151
R1058 B.n549 B.n546 10.6151
R1059 B.n546 B.n545 10.6151
R1060 B.n545 B.n542 10.6151
R1061 B.n542 B.n541 10.6151
R1062 B.n541 B.n538 10.6151
R1063 B.n538 B.n537 10.6151
R1064 B.n537 B.n534 10.6151
R1065 B.n534 B.n533 10.6151
R1066 B.n533 B.n530 10.6151
R1067 B.n530 B.n529 10.6151
R1068 B.n529 B.n526 10.6151
R1069 B.n526 B.n525 10.6151
R1070 B.n522 B.n521 10.6151
R1071 B.n521 B.n518 10.6151
R1072 B.n518 B.n517 10.6151
R1073 B.n517 B.n514 10.6151
R1074 B.n514 B.n513 10.6151
R1075 B.n513 B.n510 10.6151
R1076 B.n510 B.n509 10.6151
R1077 B.n509 B.n506 10.6151
R1078 B.n506 B.n505 10.6151
R1079 B.n502 B.n501 10.6151
R1080 B.n501 B.n498 10.6151
R1081 B.n498 B.n497 10.6151
R1082 B.n497 B.n494 10.6151
R1083 B.n494 B.n493 10.6151
R1084 B.n493 B.n490 10.6151
R1085 B.n490 B.n489 10.6151
R1086 B.n489 B.n486 10.6151
R1087 B.n486 B.n485 10.6151
R1088 B.n485 B.n482 10.6151
R1089 B.n482 B.n481 10.6151
R1090 B.n481 B.n478 10.6151
R1091 B.n478 B.n477 10.6151
R1092 B.n477 B.n474 10.6151
R1093 B.n474 B.n473 10.6151
R1094 B.n473 B.n470 10.6151
R1095 B.n470 B.n469 10.6151
R1096 B.n469 B.n466 10.6151
R1097 B.n466 B.n465 10.6151
R1098 B.n465 B.n462 10.6151
R1099 B.n462 B.n461 10.6151
R1100 B.n461 B.n458 10.6151
R1101 B.n458 B.n457 10.6151
R1102 B.n457 B.n454 10.6151
R1103 B.n454 B.n453 10.6151
R1104 B.n453 B.n450 10.6151
R1105 B.n450 B.n449 10.6151
R1106 B.n449 B.n446 10.6151
R1107 B.n446 B.n445 10.6151
R1108 B.n445 B.n442 10.6151
R1109 B.n442 B.n441 10.6151
R1110 B.n441 B.n438 10.6151
R1111 B.n438 B.n437 10.6151
R1112 B.n437 B.n434 10.6151
R1113 B.n434 B.n433 10.6151
R1114 B.n433 B.n430 10.6151
R1115 B.n430 B.n429 10.6151
R1116 B.n429 B.n426 10.6151
R1117 B.n426 B.n425 10.6151
R1118 B.n425 B.n422 10.6151
R1119 B.n422 B.n421 10.6151
R1120 B.n421 B.n418 10.6151
R1121 B.n418 B.n417 10.6151
R1122 B.n417 B.n414 10.6151
R1123 B.n414 B.n413 10.6151
R1124 B.n413 B.n411 10.6151
R1125 B.n622 B.n347 10.6151
R1126 B.n623 B.n622 10.6151
R1127 B.n624 B.n623 10.6151
R1128 B.n624 B.n339 10.6151
R1129 B.n634 B.n339 10.6151
R1130 B.n635 B.n634 10.6151
R1131 B.n636 B.n635 10.6151
R1132 B.n636 B.n331 10.6151
R1133 B.n646 B.n331 10.6151
R1134 B.n647 B.n646 10.6151
R1135 B.n648 B.n647 10.6151
R1136 B.n648 B.n323 10.6151
R1137 B.n658 B.n323 10.6151
R1138 B.n659 B.n658 10.6151
R1139 B.n660 B.n659 10.6151
R1140 B.n660 B.n314 10.6151
R1141 B.n670 B.n314 10.6151
R1142 B.n671 B.n670 10.6151
R1143 B.n673 B.n671 10.6151
R1144 B.n673 B.n672 10.6151
R1145 B.n672 B.n307 10.6151
R1146 B.n684 B.n307 10.6151
R1147 B.n685 B.n684 10.6151
R1148 B.n686 B.n685 10.6151
R1149 B.n687 B.n686 10.6151
R1150 B.n688 B.n687 10.6151
R1151 B.n691 B.n688 10.6151
R1152 B.n692 B.n691 10.6151
R1153 B.n693 B.n692 10.6151
R1154 B.n694 B.n693 10.6151
R1155 B.n696 B.n694 10.6151
R1156 B.n697 B.n696 10.6151
R1157 B.n698 B.n697 10.6151
R1158 B.n699 B.n698 10.6151
R1159 B.n701 B.n699 10.6151
R1160 B.n702 B.n701 10.6151
R1161 B.n703 B.n702 10.6151
R1162 B.n704 B.n703 10.6151
R1163 B.n706 B.n704 10.6151
R1164 B.n707 B.n706 10.6151
R1165 B.n708 B.n707 10.6151
R1166 B.n709 B.n708 10.6151
R1167 B.n711 B.n709 10.6151
R1168 B.n712 B.n711 10.6151
R1169 B.n713 B.n712 10.6151
R1170 B.n714 B.n713 10.6151
R1171 B.n715 B.n714 10.6151
R1172 B.n764 B.n1 10.6151
R1173 B.n764 B.n763 10.6151
R1174 B.n763 B.n762 10.6151
R1175 B.n762 B.n10 10.6151
R1176 B.n756 B.n10 10.6151
R1177 B.n756 B.n755 10.6151
R1178 B.n755 B.n754 10.6151
R1179 B.n754 B.n18 10.6151
R1180 B.n748 B.n18 10.6151
R1181 B.n748 B.n747 10.6151
R1182 B.n747 B.n746 10.6151
R1183 B.n746 B.n25 10.6151
R1184 B.n740 B.n25 10.6151
R1185 B.n740 B.n739 10.6151
R1186 B.n739 B.n738 10.6151
R1187 B.n738 B.n32 10.6151
R1188 B.n732 B.n32 10.6151
R1189 B.n732 B.n731 10.6151
R1190 B.n731 B.n730 10.6151
R1191 B.n730 B.n39 10.6151
R1192 B.n724 B.n39 10.6151
R1193 B.n724 B.n723 10.6151
R1194 B.n722 B.n46 10.6151
R1195 B.n105 B.n46 10.6151
R1196 B.n106 B.n105 10.6151
R1197 B.n109 B.n106 10.6151
R1198 B.n110 B.n109 10.6151
R1199 B.n113 B.n110 10.6151
R1200 B.n114 B.n113 10.6151
R1201 B.n117 B.n114 10.6151
R1202 B.n118 B.n117 10.6151
R1203 B.n121 B.n118 10.6151
R1204 B.n122 B.n121 10.6151
R1205 B.n125 B.n122 10.6151
R1206 B.n126 B.n125 10.6151
R1207 B.n129 B.n126 10.6151
R1208 B.n130 B.n129 10.6151
R1209 B.n133 B.n130 10.6151
R1210 B.n134 B.n133 10.6151
R1211 B.n137 B.n134 10.6151
R1212 B.n138 B.n137 10.6151
R1213 B.n141 B.n138 10.6151
R1214 B.n142 B.n141 10.6151
R1215 B.n145 B.n142 10.6151
R1216 B.n146 B.n145 10.6151
R1217 B.n149 B.n146 10.6151
R1218 B.n150 B.n149 10.6151
R1219 B.n153 B.n150 10.6151
R1220 B.n154 B.n153 10.6151
R1221 B.n157 B.n154 10.6151
R1222 B.n158 B.n157 10.6151
R1223 B.n161 B.n158 10.6151
R1224 B.n162 B.n161 10.6151
R1225 B.n165 B.n162 10.6151
R1226 B.n166 B.n165 10.6151
R1227 B.n169 B.n166 10.6151
R1228 B.n170 B.n169 10.6151
R1229 B.n173 B.n170 10.6151
R1230 B.n174 B.n173 10.6151
R1231 B.n177 B.n174 10.6151
R1232 B.n178 B.n177 10.6151
R1233 B.n181 B.n178 10.6151
R1234 B.n182 B.n181 10.6151
R1235 B.n185 B.n182 10.6151
R1236 B.n186 B.n185 10.6151
R1237 B.n189 B.n186 10.6151
R1238 B.n190 B.n189 10.6151
R1239 B.n193 B.n190 10.6151
R1240 B.n198 B.n195 10.6151
R1241 B.n199 B.n198 10.6151
R1242 B.n202 B.n199 10.6151
R1243 B.n203 B.n202 10.6151
R1244 B.n206 B.n203 10.6151
R1245 B.n207 B.n206 10.6151
R1246 B.n210 B.n207 10.6151
R1247 B.n211 B.n210 10.6151
R1248 B.n214 B.n211 10.6151
R1249 B.n219 B.n216 10.6151
R1250 B.n220 B.n219 10.6151
R1251 B.n223 B.n220 10.6151
R1252 B.n224 B.n223 10.6151
R1253 B.n227 B.n224 10.6151
R1254 B.n228 B.n227 10.6151
R1255 B.n231 B.n228 10.6151
R1256 B.n232 B.n231 10.6151
R1257 B.n235 B.n232 10.6151
R1258 B.n236 B.n235 10.6151
R1259 B.n239 B.n236 10.6151
R1260 B.n240 B.n239 10.6151
R1261 B.n243 B.n240 10.6151
R1262 B.n244 B.n243 10.6151
R1263 B.n247 B.n244 10.6151
R1264 B.n248 B.n247 10.6151
R1265 B.n251 B.n248 10.6151
R1266 B.n252 B.n251 10.6151
R1267 B.n255 B.n252 10.6151
R1268 B.n256 B.n255 10.6151
R1269 B.n259 B.n256 10.6151
R1270 B.n260 B.n259 10.6151
R1271 B.n263 B.n260 10.6151
R1272 B.n264 B.n263 10.6151
R1273 B.n267 B.n264 10.6151
R1274 B.n268 B.n267 10.6151
R1275 B.n271 B.n268 10.6151
R1276 B.n272 B.n271 10.6151
R1277 B.n275 B.n272 10.6151
R1278 B.n276 B.n275 10.6151
R1279 B.n279 B.n276 10.6151
R1280 B.n280 B.n279 10.6151
R1281 B.n283 B.n280 10.6151
R1282 B.n284 B.n283 10.6151
R1283 B.n287 B.n284 10.6151
R1284 B.n288 B.n287 10.6151
R1285 B.n291 B.n288 10.6151
R1286 B.n292 B.n291 10.6151
R1287 B.n295 B.n292 10.6151
R1288 B.n296 B.n295 10.6151
R1289 B.n299 B.n296 10.6151
R1290 B.n300 B.n299 10.6151
R1291 B.n303 B.n300 10.6151
R1292 B.n305 B.n303 10.6151
R1293 B.n306 B.n305 10.6151
R1294 B.n716 B.n306 10.6151
R1295 B.n525 B.n407 9.36635
R1296 B.n502 B.n410 9.36635
R1297 B.n194 B.n193 9.36635
R1298 B.n216 B.n215 9.36635
R1299 B.n772 B.n0 8.11757
R1300 B.n772 B.n1 8.11757
R1301 B.n317 B.t0 4.02454
R1302 B.t1 B.n759 4.02454
R1303 B.n522 B.n407 1.24928
R1304 B.n505 B.n410 1.24928
R1305 B.n195 B.n194 1.24928
R1306 B.n215 B.n214 1.24928
R1307 VN VN.t0 242.905
R1308 VN VN.t1 198.007
R1309 VDD2.n0 VDD2.t0 101.809
R1310 VDD2.n0 VDD2.t1 61.7532
R1311 VDD2 VDD2.n0 0.614724
C0 VTAIL VP 2.6625f
C1 VTAIL VN 2.64814f
C2 VDD2 VDD1 0.633057f
C3 VDD2 VP 0.318883f
C4 VDD2 VN 3.09769f
C5 VDD2 VTAIL 5.58172f
C6 VP VDD1 3.26519f
C7 VDD1 VN 0.148295f
C8 VP VN 5.63508f
C9 VTAIL VDD1 5.53437f
C10 VDD2 B 4.642249f
C11 VDD1 B 7.8261f
C12 VTAIL B 7.946617f
C13 VN B 10.79601f
C14 VP B 6.098492f
C15 VDD2.t0 B 3.11352f
C16 VDD2.t1 B 2.52835f
C17 VDD2.n0 B 2.94549f
C18 VN.t1 B 3.08896f
C19 VN.t0 B 3.55991f
C20 VDD1.t1 B 2.53841f
C21 VDD1.t0 B 3.15818f
C22 VTAIL.t0 B 2.45f
C23 VTAIL.n0 B 1.68994f
C24 VTAIL.t3 B 2.45001f
C25 VTAIL.n1 B 1.72229f
C26 VTAIL.t1 B 2.45001f
C27 VTAIL.n2 B 1.57769f
C28 VTAIL.t2 B 2.45f
C29 VTAIL.n3 B 1.50722f
C30 VP.t0 B 3.66633f
C31 VP.t1 B 3.18218f
C32 VP.n0 B 4.68153f
.ends

