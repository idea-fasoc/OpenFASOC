* NGSPICE file created from diff_pair_sample_0774.ext - technology: sky130A

.subckt diff_pair_sample_0774 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=0 ps=0 w=16.56 l=1.48
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=6.4584 ps=33.9 w=16.56 l=1.48
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=0 ps=0 w=16.56 l=1.48
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=0 ps=0 w=16.56 l=1.48
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=6.4584 ps=33.9 w=16.56 l=1.48
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=0 ps=0 w=16.56 l=1.48
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=6.4584 ps=33.9 w=16.56 l=1.48
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4584 pd=33.9 as=6.4584 ps=33.9 w=16.56 l=1.48
R0 B.n522 B.n521 585
R1 B.n524 B.n101 585
R2 B.n527 B.n526 585
R3 B.n528 B.n100 585
R4 B.n530 B.n529 585
R5 B.n532 B.n99 585
R6 B.n535 B.n534 585
R7 B.n536 B.n98 585
R8 B.n538 B.n537 585
R9 B.n540 B.n97 585
R10 B.n543 B.n542 585
R11 B.n544 B.n96 585
R12 B.n546 B.n545 585
R13 B.n548 B.n95 585
R14 B.n551 B.n550 585
R15 B.n552 B.n94 585
R16 B.n554 B.n553 585
R17 B.n556 B.n93 585
R18 B.n559 B.n558 585
R19 B.n560 B.n92 585
R20 B.n562 B.n561 585
R21 B.n564 B.n91 585
R22 B.n567 B.n566 585
R23 B.n568 B.n90 585
R24 B.n570 B.n569 585
R25 B.n572 B.n89 585
R26 B.n575 B.n574 585
R27 B.n576 B.n88 585
R28 B.n578 B.n577 585
R29 B.n580 B.n87 585
R30 B.n583 B.n582 585
R31 B.n584 B.n86 585
R32 B.n586 B.n585 585
R33 B.n588 B.n85 585
R34 B.n591 B.n590 585
R35 B.n592 B.n84 585
R36 B.n594 B.n593 585
R37 B.n596 B.n83 585
R38 B.n599 B.n598 585
R39 B.n600 B.n82 585
R40 B.n602 B.n601 585
R41 B.n604 B.n81 585
R42 B.n607 B.n606 585
R43 B.n608 B.n80 585
R44 B.n610 B.n609 585
R45 B.n612 B.n79 585
R46 B.n615 B.n614 585
R47 B.n616 B.n78 585
R48 B.n618 B.n617 585
R49 B.n620 B.n77 585
R50 B.n623 B.n622 585
R51 B.n624 B.n76 585
R52 B.n626 B.n625 585
R53 B.n628 B.n75 585
R54 B.n631 B.n630 585
R55 B.n633 B.n72 585
R56 B.n635 B.n634 585
R57 B.n637 B.n71 585
R58 B.n640 B.n639 585
R59 B.n641 B.n70 585
R60 B.n643 B.n642 585
R61 B.n645 B.n69 585
R62 B.n648 B.n647 585
R63 B.n649 B.n65 585
R64 B.n651 B.n650 585
R65 B.n653 B.n64 585
R66 B.n656 B.n655 585
R67 B.n657 B.n63 585
R68 B.n659 B.n658 585
R69 B.n661 B.n62 585
R70 B.n664 B.n663 585
R71 B.n665 B.n61 585
R72 B.n667 B.n666 585
R73 B.n669 B.n60 585
R74 B.n672 B.n671 585
R75 B.n673 B.n59 585
R76 B.n675 B.n674 585
R77 B.n677 B.n58 585
R78 B.n680 B.n679 585
R79 B.n681 B.n57 585
R80 B.n683 B.n682 585
R81 B.n685 B.n56 585
R82 B.n688 B.n687 585
R83 B.n689 B.n55 585
R84 B.n691 B.n690 585
R85 B.n693 B.n54 585
R86 B.n696 B.n695 585
R87 B.n697 B.n53 585
R88 B.n699 B.n698 585
R89 B.n701 B.n52 585
R90 B.n704 B.n703 585
R91 B.n705 B.n51 585
R92 B.n707 B.n706 585
R93 B.n709 B.n50 585
R94 B.n712 B.n711 585
R95 B.n713 B.n49 585
R96 B.n715 B.n714 585
R97 B.n717 B.n48 585
R98 B.n720 B.n719 585
R99 B.n721 B.n47 585
R100 B.n723 B.n722 585
R101 B.n725 B.n46 585
R102 B.n728 B.n727 585
R103 B.n729 B.n45 585
R104 B.n731 B.n730 585
R105 B.n733 B.n44 585
R106 B.n736 B.n735 585
R107 B.n737 B.n43 585
R108 B.n739 B.n738 585
R109 B.n741 B.n42 585
R110 B.n744 B.n743 585
R111 B.n745 B.n41 585
R112 B.n747 B.n746 585
R113 B.n749 B.n40 585
R114 B.n752 B.n751 585
R115 B.n753 B.n39 585
R116 B.n755 B.n754 585
R117 B.n757 B.n38 585
R118 B.n760 B.n759 585
R119 B.n761 B.n37 585
R120 B.n520 B.n35 585
R121 B.n764 B.n35 585
R122 B.n519 B.n34 585
R123 B.n765 B.n34 585
R124 B.n518 B.n33 585
R125 B.n766 B.n33 585
R126 B.n517 B.n516 585
R127 B.n516 B.n29 585
R128 B.n515 B.n28 585
R129 B.n772 B.n28 585
R130 B.n514 B.n27 585
R131 B.n773 B.n27 585
R132 B.n513 B.n26 585
R133 B.n774 B.n26 585
R134 B.n512 B.n511 585
R135 B.n511 B.n22 585
R136 B.n510 B.n21 585
R137 B.n780 B.n21 585
R138 B.n509 B.n20 585
R139 B.n781 B.n20 585
R140 B.n508 B.n19 585
R141 B.n782 B.n19 585
R142 B.n507 B.n506 585
R143 B.n506 B.n15 585
R144 B.n505 B.n14 585
R145 B.n788 B.n14 585
R146 B.n504 B.n13 585
R147 B.n789 B.n13 585
R148 B.n503 B.n12 585
R149 B.n790 B.n12 585
R150 B.n502 B.n501 585
R151 B.n501 B.n500 585
R152 B.n499 B.n498 585
R153 B.n499 B.n8 585
R154 B.n497 B.n7 585
R155 B.n797 B.n7 585
R156 B.n496 B.n6 585
R157 B.n798 B.n6 585
R158 B.n495 B.n5 585
R159 B.n799 B.n5 585
R160 B.n494 B.n493 585
R161 B.n493 B.n4 585
R162 B.n492 B.n102 585
R163 B.n492 B.n491 585
R164 B.n482 B.n103 585
R165 B.n104 B.n103 585
R166 B.n484 B.n483 585
R167 B.n485 B.n484 585
R168 B.n481 B.n109 585
R169 B.n109 B.n108 585
R170 B.n480 B.n479 585
R171 B.n479 B.n478 585
R172 B.n111 B.n110 585
R173 B.n112 B.n111 585
R174 B.n471 B.n470 585
R175 B.n472 B.n471 585
R176 B.n469 B.n117 585
R177 B.n117 B.n116 585
R178 B.n468 B.n467 585
R179 B.n467 B.n466 585
R180 B.n119 B.n118 585
R181 B.n120 B.n119 585
R182 B.n459 B.n458 585
R183 B.n460 B.n459 585
R184 B.n457 B.n124 585
R185 B.n128 B.n124 585
R186 B.n456 B.n455 585
R187 B.n455 B.n454 585
R188 B.n126 B.n125 585
R189 B.n127 B.n126 585
R190 B.n447 B.n446 585
R191 B.n448 B.n447 585
R192 B.n445 B.n133 585
R193 B.n133 B.n132 585
R194 B.n444 B.n443 585
R195 B.n443 B.n442 585
R196 B.n439 B.n137 585
R197 B.n438 B.n437 585
R198 B.n435 B.n138 585
R199 B.n435 B.n136 585
R200 B.n434 B.n433 585
R201 B.n432 B.n431 585
R202 B.n430 B.n140 585
R203 B.n428 B.n427 585
R204 B.n426 B.n141 585
R205 B.n425 B.n424 585
R206 B.n422 B.n142 585
R207 B.n420 B.n419 585
R208 B.n418 B.n143 585
R209 B.n417 B.n416 585
R210 B.n414 B.n144 585
R211 B.n412 B.n411 585
R212 B.n410 B.n145 585
R213 B.n409 B.n408 585
R214 B.n406 B.n146 585
R215 B.n404 B.n403 585
R216 B.n402 B.n147 585
R217 B.n401 B.n400 585
R218 B.n398 B.n148 585
R219 B.n396 B.n395 585
R220 B.n394 B.n149 585
R221 B.n393 B.n392 585
R222 B.n390 B.n150 585
R223 B.n388 B.n387 585
R224 B.n386 B.n151 585
R225 B.n385 B.n384 585
R226 B.n382 B.n152 585
R227 B.n380 B.n379 585
R228 B.n378 B.n153 585
R229 B.n377 B.n376 585
R230 B.n374 B.n154 585
R231 B.n372 B.n371 585
R232 B.n370 B.n155 585
R233 B.n369 B.n368 585
R234 B.n366 B.n156 585
R235 B.n364 B.n363 585
R236 B.n362 B.n157 585
R237 B.n361 B.n360 585
R238 B.n358 B.n158 585
R239 B.n356 B.n355 585
R240 B.n354 B.n159 585
R241 B.n353 B.n352 585
R242 B.n350 B.n160 585
R243 B.n348 B.n347 585
R244 B.n346 B.n161 585
R245 B.n345 B.n344 585
R246 B.n342 B.n162 585
R247 B.n340 B.n339 585
R248 B.n338 B.n163 585
R249 B.n337 B.n336 585
R250 B.n334 B.n164 585
R251 B.n332 B.n331 585
R252 B.n329 B.n165 585
R253 B.n328 B.n327 585
R254 B.n325 B.n168 585
R255 B.n323 B.n322 585
R256 B.n321 B.n169 585
R257 B.n320 B.n319 585
R258 B.n317 B.n170 585
R259 B.n315 B.n314 585
R260 B.n313 B.n171 585
R261 B.n312 B.n311 585
R262 B.n309 B.n308 585
R263 B.n307 B.n306 585
R264 B.n305 B.n176 585
R265 B.n303 B.n302 585
R266 B.n301 B.n177 585
R267 B.n300 B.n299 585
R268 B.n297 B.n178 585
R269 B.n295 B.n294 585
R270 B.n293 B.n179 585
R271 B.n292 B.n291 585
R272 B.n289 B.n180 585
R273 B.n287 B.n286 585
R274 B.n285 B.n181 585
R275 B.n284 B.n283 585
R276 B.n281 B.n182 585
R277 B.n279 B.n278 585
R278 B.n277 B.n183 585
R279 B.n276 B.n275 585
R280 B.n273 B.n184 585
R281 B.n271 B.n270 585
R282 B.n269 B.n185 585
R283 B.n268 B.n267 585
R284 B.n265 B.n186 585
R285 B.n263 B.n262 585
R286 B.n261 B.n187 585
R287 B.n260 B.n259 585
R288 B.n257 B.n188 585
R289 B.n255 B.n254 585
R290 B.n253 B.n189 585
R291 B.n252 B.n251 585
R292 B.n249 B.n190 585
R293 B.n247 B.n246 585
R294 B.n245 B.n191 585
R295 B.n244 B.n243 585
R296 B.n241 B.n192 585
R297 B.n239 B.n238 585
R298 B.n237 B.n193 585
R299 B.n236 B.n235 585
R300 B.n233 B.n194 585
R301 B.n231 B.n230 585
R302 B.n229 B.n195 585
R303 B.n228 B.n227 585
R304 B.n225 B.n196 585
R305 B.n223 B.n222 585
R306 B.n221 B.n197 585
R307 B.n220 B.n219 585
R308 B.n217 B.n198 585
R309 B.n215 B.n214 585
R310 B.n213 B.n199 585
R311 B.n212 B.n211 585
R312 B.n209 B.n200 585
R313 B.n207 B.n206 585
R314 B.n205 B.n201 585
R315 B.n204 B.n203 585
R316 B.n135 B.n134 585
R317 B.n136 B.n135 585
R318 B.n441 B.n440 585
R319 B.n442 B.n441 585
R320 B.n131 B.n130 585
R321 B.n132 B.n131 585
R322 B.n450 B.n449 585
R323 B.n449 B.n448 585
R324 B.n451 B.n129 585
R325 B.n129 B.n127 585
R326 B.n453 B.n452 585
R327 B.n454 B.n453 585
R328 B.n123 B.n122 585
R329 B.n128 B.n123 585
R330 B.n462 B.n461 585
R331 B.n461 B.n460 585
R332 B.n463 B.n121 585
R333 B.n121 B.n120 585
R334 B.n465 B.n464 585
R335 B.n466 B.n465 585
R336 B.n115 B.n114 585
R337 B.n116 B.n115 585
R338 B.n474 B.n473 585
R339 B.n473 B.n472 585
R340 B.n475 B.n113 585
R341 B.n113 B.n112 585
R342 B.n477 B.n476 585
R343 B.n478 B.n477 585
R344 B.n107 B.n106 585
R345 B.n108 B.n107 585
R346 B.n487 B.n486 585
R347 B.n486 B.n485 585
R348 B.n488 B.n105 585
R349 B.n105 B.n104 585
R350 B.n490 B.n489 585
R351 B.n491 B.n490 585
R352 B.n3 B.n0 585
R353 B.n4 B.n3 585
R354 B.n796 B.n1 585
R355 B.n797 B.n796 585
R356 B.n795 B.n794 585
R357 B.n795 B.n8 585
R358 B.n793 B.n9 585
R359 B.n500 B.n9 585
R360 B.n792 B.n791 585
R361 B.n791 B.n790 585
R362 B.n11 B.n10 585
R363 B.n789 B.n11 585
R364 B.n787 B.n786 585
R365 B.n788 B.n787 585
R366 B.n785 B.n16 585
R367 B.n16 B.n15 585
R368 B.n784 B.n783 585
R369 B.n783 B.n782 585
R370 B.n18 B.n17 585
R371 B.n781 B.n18 585
R372 B.n779 B.n778 585
R373 B.n780 B.n779 585
R374 B.n777 B.n23 585
R375 B.n23 B.n22 585
R376 B.n776 B.n775 585
R377 B.n775 B.n774 585
R378 B.n25 B.n24 585
R379 B.n773 B.n25 585
R380 B.n771 B.n770 585
R381 B.n772 B.n771 585
R382 B.n769 B.n30 585
R383 B.n30 B.n29 585
R384 B.n768 B.n767 585
R385 B.n767 B.n766 585
R386 B.n32 B.n31 585
R387 B.n765 B.n32 585
R388 B.n763 B.n762 585
R389 B.n764 B.n763 585
R390 B.n800 B.n799 585
R391 B.n798 B.n2 585
R392 B.n763 B.n37 511.721
R393 B.n522 B.n35 511.721
R394 B.n443 B.n135 511.721
R395 B.n441 B.n137 511.721
R396 B.n66 B.t6 475.024
R397 B.n73 B.t2 475.024
R398 B.n172 B.t13 475.024
R399 B.n166 B.t9 475.024
R400 B.n523 B.n36 256.663
R401 B.n525 B.n36 256.663
R402 B.n531 B.n36 256.663
R403 B.n533 B.n36 256.663
R404 B.n539 B.n36 256.663
R405 B.n541 B.n36 256.663
R406 B.n547 B.n36 256.663
R407 B.n549 B.n36 256.663
R408 B.n555 B.n36 256.663
R409 B.n557 B.n36 256.663
R410 B.n563 B.n36 256.663
R411 B.n565 B.n36 256.663
R412 B.n571 B.n36 256.663
R413 B.n573 B.n36 256.663
R414 B.n579 B.n36 256.663
R415 B.n581 B.n36 256.663
R416 B.n587 B.n36 256.663
R417 B.n589 B.n36 256.663
R418 B.n595 B.n36 256.663
R419 B.n597 B.n36 256.663
R420 B.n603 B.n36 256.663
R421 B.n605 B.n36 256.663
R422 B.n611 B.n36 256.663
R423 B.n613 B.n36 256.663
R424 B.n619 B.n36 256.663
R425 B.n621 B.n36 256.663
R426 B.n627 B.n36 256.663
R427 B.n629 B.n36 256.663
R428 B.n636 B.n36 256.663
R429 B.n638 B.n36 256.663
R430 B.n644 B.n36 256.663
R431 B.n646 B.n36 256.663
R432 B.n652 B.n36 256.663
R433 B.n654 B.n36 256.663
R434 B.n660 B.n36 256.663
R435 B.n662 B.n36 256.663
R436 B.n668 B.n36 256.663
R437 B.n670 B.n36 256.663
R438 B.n676 B.n36 256.663
R439 B.n678 B.n36 256.663
R440 B.n684 B.n36 256.663
R441 B.n686 B.n36 256.663
R442 B.n692 B.n36 256.663
R443 B.n694 B.n36 256.663
R444 B.n700 B.n36 256.663
R445 B.n702 B.n36 256.663
R446 B.n708 B.n36 256.663
R447 B.n710 B.n36 256.663
R448 B.n716 B.n36 256.663
R449 B.n718 B.n36 256.663
R450 B.n724 B.n36 256.663
R451 B.n726 B.n36 256.663
R452 B.n732 B.n36 256.663
R453 B.n734 B.n36 256.663
R454 B.n740 B.n36 256.663
R455 B.n742 B.n36 256.663
R456 B.n748 B.n36 256.663
R457 B.n750 B.n36 256.663
R458 B.n756 B.n36 256.663
R459 B.n758 B.n36 256.663
R460 B.n436 B.n136 256.663
R461 B.n139 B.n136 256.663
R462 B.n429 B.n136 256.663
R463 B.n423 B.n136 256.663
R464 B.n421 B.n136 256.663
R465 B.n415 B.n136 256.663
R466 B.n413 B.n136 256.663
R467 B.n407 B.n136 256.663
R468 B.n405 B.n136 256.663
R469 B.n399 B.n136 256.663
R470 B.n397 B.n136 256.663
R471 B.n391 B.n136 256.663
R472 B.n389 B.n136 256.663
R473 B.n383 B.n136 256.663
R474 B.n381 B.n136 256.663
R475 B.n375 B.n136 256.663
R476 B.n373 B.n136 256.663
R477 B.n367 B.n136 256.663
R478 B.n365 B.n136 256.663
R479 B.n359 B.n136 256.663
R480 B.n357 B.n136 256.663
R481 B.n351 B.n136 256.663
R482 B.n349 B.n136 256.663
R483 B.n343 B.n136 256.663
R484 B.n341 B.n136 256.663
R485 B.n335 B.n136 256.663
R486 B.n333 B.n136 256.663
R487 B.n326 B.n136 256.663
R488 B.n324 B.n136 256.663
R489 B.n318 B.n136 256.663
R490 B.n316 B.n136 256.663
R491 B.n310 B.n136 256.663
R492 B.n175 B.n136 256.663
R493 B.n304 B.n136 256.663
R494 B.n298 B.n136 256.663
R495 B.n296 B.n136 256.663
R496 B.n290 B.n136 256.663
R497 B.n288 B.n136 256.663
R498 B.n282 B.n136 256.663
R499 B.n280 B.n136 256.663
R500 B.n274 B.n136 256.663
R501 B.n272 B.n136 256.663
R502 B.n266 B.n136 256.663
R503 B.n264 B.n136 256.663
R504 B.n258 B.n136 256.663
R505 B.n256 B.n136 256.663
R506 B.n250 B.n136 256.663
R507 B.n248 B.n136 256.663
R508 B.n242 B.n136 256.663
R509 B.n240 B.n136 256.663
R510 B.n234 B.n136 256.663
R511 B.n232 B.n136 256.663
R512 B.n226 B.n136 256.663
R513 B.n224 B.n136 256.663
R514 B.n218 B.n136 256.663
R515 B.n216 B.n136 256.663
R516 B.n210 B.n136 256.663
R517 B.n208 B.n136 256.663
R518 B.n202 B.n136 256.663
R519 B.n802 B.n801 256.663
R520 B.n759 B.n757 163.367
R521 B.n755 B.n39 163.367
R522 B.n751 B.n749 163.367
R523 B.n747 B.n41 163.367
R524 B.n743 B.n741 163.367
R525 B.n739 B.n43 163.367
R526 B.n735 B.n733 163.367
R527 B.n731 B.n45 163.367
R528 B.n727 B.n725 163.367
R529 B.n723 B.n47 163.367
R530 B.n719 B.n717 163.367
R531 B.n715 B.n49 163.367
R532 B.n711 B.n709 163.367
R533 B.n707 B.n51 163.367
R534 B.n703 B.n701 163.367
R535 B.n699 B.n53 163.367
R536 B.n695 B.n693 163.367
R537 B.n691 B.n55 163.367
R538 B.n687 B.n685 163.367
R539 B.n683 B.n57 163.367
R540 B.n679 B.n677 163.367
R541 B.n675 B.n59 163.367
R542 B.n671 B.n669 163.367
R543 B.n667 B.n61 163.367
R544 B.n663 B.n661 163.367
R545 B.n659 B.n63 163.367
R546 B.n655 B.n653 163.367
R547 B.n651 B.n65 163.367
R548 B.n647 B.n645 163.367
R549 B.n643 B.n70 163.367
R550 B.n639 B.n637 163.367
R551 B.n635 B.n72 163.367
R552 B.n630 B.n628 163.367
R553 B.n626 B.n76 163.367
R554 B.n622 B.n620 163.367
R555 B.n618 B.n78 163.367
R556 B.n614 B.n612 163.367
R557 B.n610 B.n80 163.367
R558 B.n606 B.n604 163.367
R559 B.n602 B.n82 163.367
R560 B.n598 B.n596 163.367
R561 B.n594 B.n84 163.367
R562 B.n590 B.n588 163.367
R563 B.n586 B.n86 163.367
R564 B.n582 B.n580 163.367
R565 B.n578 B.n88 163.367
R566 B.n574 B.n572 163.367
R567 B.n570 B.n90 163.367
R568 B.n566 B.n564 163.367
R569 B.n562 B.n92 163.367
R570 B.n558 B.n556 163.367
R571 B.n554 B.n94 163.367
R572 B.n550 B.n548 163.367
R573 B.n546 B.n96 163.367
R574 B.n542 B.n540 163.367
R575 B.n538 B.n98 163.367
R576 B.n534 B.n532 163.367
R577 B.n530 B.n100 163.367
R578 B.n526 B.n524 163.367
R579 B.n443 B.n133 163.367
R580 B.n447 B.n133 163.367
R581 B.n447 B.n126 163.367
R582 B.n455 B.n126 163.367
R583 B.n455 B.n124 163.367
R584 B.n459 B.n124 163.367
R585 B.n459 B.n119 163.367
R586 B.n467 B.n119 163.367
R587 B.n467 B.n117 163.367
R588 B.n471 B.n117 163.367
R589 B.n471 B.n111 163.367
R590 B.n479 B.n111 163.367
R591 B.n479 B.n109 163.367
R592 B.n484 B.n109 163.367
R593 B.n484 B.n103 163.367
R594 B.n492 B.n103 163.367
R595 B.n493 B.n492 163.367
R596 B.n493 B.n5 163.367
R597 B.n6 B.n5 163.367
R598 B.n7 B.n6 163.367
R599 B.n499 B.n7 163.367
R600 B.n501 B.n499 163.367
R601 B.n501 B.n12 163.367
R602 B.n13 B.n12 163.367
R603 B.n14 B.n13 163.367
R604 B.n506 B.n14 163.367
R605 B.n506 B.n19 163.367
R606 B.n20 B.n19 163.367
R607 B.n21 B.n20 163.367
R608 B.n511 B.n21 163.367
R609 B.n511 B.n26 163.367
R610 B.n27 B.n26 163.367
R611 B.n28 B.n27 163.367
R612 B.n516 B.n28 163.367
R613 B.n516 B.n33 163.367
R614 B.n34 B.n33 163.367
R615 B.n35 B.n34 163.367
R616 B.n437 B.n435 163.367
R617 B.n435 B.n434 163.367
R618 B.n431 B.n430 163.367
R619 B.n428 B.n141 163.367
R620 B.n424 B.n422 163.367
R621 B.n420 B.n143 163.367
R622 B.n416 B.n414 163.367
R623 B.n412 B.n145 163.367
R624 B.n408 B.n406 163.367
R625 B.n404 B.n147 163.367
R626 B.n400 B.n398 163.367
R627 B.n396 B.n149 163.367
R628 B.n392 B.n390 163.367
R629 B.n388 B.n151 163.367
R630 B.n384 B.n382 163.367
R631 B.n380 B.n153 163.367
R632 B.n376 B.n374 163.367
R633 B.n372 B.n155 163.367
R634 B.n368 B.n366 163.367
R635 B.n364 B.n157 163.367
R636 B.n360 B.n358 163.367
R637 B.n356 B.n159 163.367
R638 B.n352 B.n350 163.367
R639 B.n348 B.n161 163.367
R640 B.n344 B.n342 163.367
R641 B.n340 B.n163 163.367
R642 B.n336 B.n334 163.367
R643 B.n332 B.n165 163.367
R644 B.n327 B.n325 163.367
R645 B.n323 B.n169 163.367
R646 B.n319 B.n317 163.367
R647 B.n315 B.n171 163.367
R648 B.n311 B.n309 163.367
R649 B.n306 B.n305 163.367
R650 B.n303 B.n177 163.367
R651 B.n299 B.n297 163.367
R652 B.n295 B.n179 163.367
R653 B.n291 B.n289 163.367
R654 B.n287 B.n181 163.367
R655 B.n283 B.n281 163.367
R656 B.n279 B.n183 163.367
R657 B.n275 B.n273 163.367
R658 B.n271 B.n185 163.367
R659 B.n267 B.n265 163.367
R660 B.n263 B.n187 163.367
R661 B.n259 B.n257 163.367
R662 B.n255 B.n189 163.367
R663 B.n251 B.n249 163.367
R664 B.n247 B.n191 163.367
R665 B.n243 B.n241 163.367
R666 B.n239 B.n193 163.367
R667 B.n235 B.n233 163.367
R668 B.n231 B.n195 163.367
R669 B.n227 B.n225 163.367
R670 B.n223 B.n197 163.367
R671 B.n219 B.n217 163.367
R672 B.n215 B.n199 163.367
R673 B.n211 B.n209 163.367
R674 B.n207 B.n201 163.367
R675 B.n203 B.n135 163.367
R676 B.n441 B.n131 163.367
R677 B.n449 B.n131 163.367
R678 B.n449 B.n129 163.367
R679 B.n453 B.n129 163.367
R680 B.n453 B.n123 163.367
R681 B.n461 B.n123 163.367
R682 B.n461 B.n121 163.367
R683 B.n465 B.n121 163.367
R684 B.n465 B.n115 163.367
R685 B.n473 B.n115 163.367
R686 B.n473 B.n113 163.367
R687 B.n477 B.n113 163.367
R688 B.n477 B.n107 163.367
R689 B.n486 B.n107 163.367
R690 B.n486 B.n105 163.367
R691 B.n490 B.n105 163.367
R692 B.n490 B.n3 163.367
R693 B.n800 B.n3 163.367
R694 B.n796 B.n2 163.367
R695 B.n796 B.n795 163.367
R696 B.n795 B.n9 163.367
R697 B.n791 B.n9 163.367
R698 B.n791 B.n11 163.367
R699 B.n787 B.n11 163.367
R700 B.n787 B.n16 163.367
R701 B.n783 B.n16 163.367
R702 B.n783 B.n18 163.367
R703 B.n779 B.n18 163.367
R704 B.n779 B.n23 163.367
R705 B.n775 B.n23 163.367
R706 B.n775 B.n25 163.367
R707 B.n771 B.n25 163.367
R708 B.n771 B.n30 163.367
R709 B.n767 B.n30 163.367
R710 B.n767 B.n32 163.367
R711 B.n763 B.n32 163.367
R712 B.n73 B.t4 107.1
R713 B.n172 B.t15 107.1
R714 B.n66 B.t7 107.078
R715 B.n166 B.t12 107.078
R716 B.n74 B.t5 71.9966
R717 B.n173 B.t14 71.9966
R718 B.n67 B.t8 71.9749
R719 B.n167 B.t11 71.9749
R720 B.n758 B.n37 71.676
R721 B.n757 B.n756 71.676
R722 B.n750 B.n39 71.676
R723 B.n749 B.n748 71.676
R724 B.n742 B.n41 71.676
R725 B.n741 B.n740 71.676
R726 B.n734 B.n43 71.676
R727 B.n733 B.n732 71.676
R728 B.n726 B.n45 71.676
R729 B.n725 B.n724 71.676
R730 B.n718 B.n47 71.676
R731 B.n717 B.n716 71.676
R732 B.n710 B.n49 71.676
R733 B.n709 B.n708 71.676
R734 B.n702 B.n51 71.676
R735 B.n701 B.n700 71.676
R736 B.n694 B.n53 71.676
R737 B.n693 B.n692 71.676
R738 B.n686 B.n55 71.676
R739 B.n685 B.n684 71.676
R740 B.n678 B.n57 71.676
R741 B.n677 B.n676 71.676
R742 B.n670 B.n59 71.676
R743 B.n669 B.n668 71.676
R744 B.n662 B.n61 71.676
R745 B.n661 B.n660 71.676
R746 B.n654 B.n63 71.676
R747 B.n653 B.n652 71.676
R748 B.n646 B.n65 71.676
R749 B.n645 B.n644 71.676
R750 B.n638 B.n70 71.676
R751 B.n637 B.n636 71.676
R752 B.n629 B.n72 71.676
R753 B.n628 B.n627 71.676
R754 B.n621 B.n76 71.676
R755 B.n620 B.n619 71.676
R756 B.n613 B.n78 71.676
R757 B.n612 B.n611 71.676
R758 B.n605 B.n80 71.676
R759 B.n604 B.n603 71.676
R760 B.n597 B.n82 71.676
R761 B.n596 B.n595 71.676
R762 B.n589 B.n84 71.676
R763 B.n588 B.n587 71.676
R764 B.n581 B.n86 71.676
R765 B.n580 B.n579 71.676
R766 B.n573 B.n88 71.676
R767 B.n572 B.n571 71.676
R768 B.n565 B.n90 71.676
R769 B.n564 B.n563 71.676
R770 B.n557 B.n92 71.676
R771 B.n556 B.n555 71.676
R772 B.n549 B.n94 71.676
R773 B.n548 B.n547 71.676
R774 B.n541 B.n96 71.676
R775 B.n540 B.n539 71.676
R776 B.n533 B.n98 71.676
R777 B.n532 B.n531 71.676
R778 B.n525 B.n100 71.676
R779 B.n524 B.n523 71.676
R780 B.n523 B.n522 71.676
R781 B.n526 B.n525 71.676
R782 B.n531 B.n530 71.676
R783 B.n534 B.n533 71.676
R784 B.n539 B.n538 71.676
R785 B.n542 B.n541 71.676
R786 B.n547 B.n546 71.676
R787 B.n550 B.n549 71.676
R788 B.n555 B.n554 71.676
R789 B.n558 B.n557 71.676
R790 B.n563 B.n562 71.676
R791 B.n566 B.n565 71.676
R792 B.n571 B.n570 71.676
R793 B.n574 B.n573 71.676
R794 B.n579 B.n578 71.676
R795 B.n582 B.n581 71.676
R796 B.n587 B.n586 71.676
R797 B.n590 B.n589 71.676
R798 B.n595 B.n594 71.676
R799 B.n598 B.n597 71.676
R800 B.n603 B.n602 71.676
R801 B.n606 B.n605 71.676
R802 B.n611 B.n610 71.676
R803 B.n614 B.n613 71.676
R804 B.n619 B.n618 71.676
R805 B.n622 B.n621 71.676
R806 B.n627 B.n626 71.676
R807 B.n630 B.n629 71.676
R808 B.n636 B.n635 71.676
R809 B.n639 B.n638 71.676
R810 B.n644 B.n643 71.676
R811 B.n647 B.n646 71.676
R812 B.n652 B.n651 71.676
R813 B.n655 B.n654 71.676
R814 B.n660 B.n659 71.676
R815 B.n663 B.n662 71.676
R816 B.n668 B.n667 71.676
R817 B.n671 B.n670 71.676
R818 B.n676 B.n675 71.676
R819 B.n679 B.n678 71.676
R820 B.n684 B.n683 71.676
R821 B.n687 B.n686 71.676
R822 B.n692 B.n691 71.676
R823 B.n695 B.n694 71.676
R824 B.n700 B.n699 71.676
R825 B.n703 B.n702 71.676
R826 B.n708 B.n707 71.676
R827 B.n711 B.n710 71.676
R828 B.n716 B.n715 71.676
R829 B.n719 B.n718 71.676
R830 B.n724 B.n723 71.676
R831 B.n727 B.n726 71.676
R832 B.n732 B.n731 71.676
R833 B.n735 B.n734 71.676
R834 B.n740 B.n739 71.676
R835 B.n743 B.n742 71.676
R836 B.n748 B.n747 71.676
R837 B.n751 B.n750 71.676
R838 B.n756 B.n755 71.676
R839 B.n759 B.n758 71.676
R840 B.n436 B.n137 71.676
R841 B.n434 B.n139 71.676
R842 B.n430 B.n429 71.676
R843 B.n423 B.n141 71.676
R844 B.n422 B.n421 71.676
R845 B.n415 B.n143 71.676
R846 B.n414 B.n413 71.676
R847 B.n407 B.n145 71.676
R848 B.n406 B.n405 71.676
R849 B.n399 B.n147 71.676
R850 B.n398 B.n397 71.676
R851 B.n391 B.n149 71.676
R852 B.n390 B.n389 71.676
R853 B.n383 B.n151 71.676
R854 B.n382 B.n381 71.676
R855 B.n375 B.n153 71.676
R856 B.n374 B.n373 71.676
R857 B.n367 B.n155 71.676
R858 B.n366 B.n365 71.676
R859 B.n359 B.n157 71.676
R860 B.n358 B.n357 71.676
R861 B.n351 B.n159 71.676
R862 B.n350 B.n349 71.676
R863 B.n343 B.n161 71.676
R864 B.n342 B.n341 71.676
R865 B.n335 B.n163 71.676
R866 B.n334 B.n333 71.676
R867 B.n326 B.n165 71.676
R868 B.n325 B.n324 71.676
R869 B.n318 B.n169 71.676
R870 B.n317 B.n316 71.676
R871 B.n310 B.n171 71.676
R872 B.n309 B.n175 71.676
R873 B.n305 B.n304 71.676
R874 B.n298 B.n177 71.676
R875 B.n297 B.n296 71.676
R876 B.n290 B.n179 71.676
R877 B.n289 B.n288 71.676
R878 B.n282 B.n181 71.676
R879 B.n281 B.n280 71.676
R880 B.n274 B.n183 71.676
R881 B.n273 B.n272 71.676
R882 B.n266 B.n185 71.676
R883 B.n265 B.n264 71.676
R884 B.n258 B.n187 71.676
R885 B.n257 B.n256 71.676
R886 B.n250 B.n189 71.676
R887 B.n249 B.n248 71.676
R888 B.n242 B.n191 71.676
R889 B.n241 B.n240 71.676
R890 B.n234 B.n193 71.676
R891 B.n233 B.n232 71.676
R892 B.n226 B.n195 71.676
R893 B.n225 B.n224 71.676
R894 B.n218 B.n197 71.676
R895 B.n217 B.n216 71.676
R896 B.n210 B.n199 71.676
R897 B.n209 B.n208 71.676
R898 B.n202 B.n201 71.676
R899 B.n437 B.n436 71.676
R900 B.n431 B.n139 71.676
R901 B.n429 B.n428 71.676
R902 B.n424 B.n423 71.676
R903 B.n421 B.n420 71.676
R904 B.n416 B.n415 71.676
R905 B.n413 B.n412 71.676
R906 B.n408 B.n407 71.676
R907 B.n405 B.n404 71.676
R908 B.n400 B.n399 71.676
R909 B.n397 B.n396 71.676
R910 B.n392 B.n391 71.676
R911 B.n389 B.n388 71.676
R912 B.n384 B.n383 71.676
R913 B.n381 B.n380 71.676
R914 B.n376 B.n375 71.676
R915 B.n373 B.n372 71.676
R916 B.n368 B.n367 71.676
R917 B.n365 B.n364 71.676
R918 B.n360 B.n359 71.676
R919 B.n357 B.n356 71.676
R920 B.n352 B.n351 71.676
R921 B.n349 B.n348 71.676
R922 B.n344 B.n343 71.676
R923 B.n341 B.n340 71.676
R924 B.n336 B.n335 71.676
R925 B.n333 B.n332 71.676
R926 B.n327 B.n326 71.676
R927 B.n324 B.n323 71.676
R928 B.n319 B.n318 71.676
R929 B.n316 B.n315 71.676
R930 B.n311 B.n310 71.676
R931 B.n306 B.n175 71.676
R932 B.n304 B.n303 71.676
R933 B.n299 B.n298 71.676
R934 B.n296 B.n295 71.676
R935 B.n291 B.n290 71.676
R936 B.n288 B.n287 71.676
R937 B.n283 B.n282 71.676
R938 B.n280 B.n279 71.676
R939 B.n275 B.n274 71.676
R940 B.n272 B.n271 71.676
R941 B.n267 B.n266 71.676
R942 B.n264 B.n263 71.676
R943 B.n259 B.n258 71.676
R944 B.n256 B.n255 71.676
R945 B.n251 B.n250 71.676
R946 B.n248 B.n247 71.676
R947 B.n243 B.n242 71.676
R948 B.n240 B.n239 71.676
R949 B.n235 B.n234 71.676
R950 B.n232 B.n231 71.676
R951 B.n227 B.n226 71.676
R952 B.n224 B.n223 71.676
R953 B.n219 B.n218 71.676
R954 B.n216 B.n215 71.676
R955 B.n211 B.n210 71.676
R956 B.n208 B.n207 71.676
R957 B.n203 B.n202 71.676
R958 B.n801 B.n800 71.676
R959 B.n801 B.n2 71.676
R960 B.n442 B.n136 71.0332
R961 B.n764 B.n36 71.0332
R962 B.n68 B.n67 59.5399
R963 B.n632 B.n74 59.5399
R964 B.n174 B.n173 59.5399
R965 B.n330 B.n167 59.5399
R966 B.n67 B.n66 35.1035
R967 B.n74 B.n73 35.1035
R968 B.n173 B.n172 35.1035
R969 B.n167 B.n166 35.1035
R970 B.n442 B.n132 34.2574
R971 B.n448 B.n132 34.2574
R972 B.n448 B.n127 34.2574
R973 B.n454 B.n127 34.2574
R974 B.n454 B.n128 34.2574
R975 B.n460 B.n120 34.2574
R976 B.n466 B.n120 34.2574
R977 B.n466 B.n116 34.2574
R978 B.n472 B.n116 34.2574
R979 B.n472 B.n112 34.2574
R980 B.n478 B.n112 34.2574
R981 B.n478 B.n108 34.2574
R982 B.n485 B.n108 34.2574
R983 B.n491 B.n104 34.2574
R984 B.n491 B.n4 34.2574
R985 B.n799 B.n4 34.2574
R986 B.n799 B.n798 34.2574
R987 B.n798 B.n797 34.2574
R988 B.n797 B.n8 34.2574
R989 B.n500 B.n8 34.2574
R990 B.n790 B.n789 34.2574
R991 B.n789 B.n788 34.2574
R992 B.n788 B.n15 34.2574
R993 B.n782 B.n15 34.2574
R994 B.n782 B.n781 34.2574
R995 B.n781 B.n780 34.2574
R996 B.n780 B.n22 34.2574
R997 B.n774 B.n22 34.2574
R998 B.n773 B.n772 34.2574
R999 B.n772 B.n29 34.2574
R1000 B.n766 B.n29 34.2574
R1001 B.n766 B.n765 34.2574
R1002 B.n765 B.n764 34.2574
R1003 B.n440 B.n439 33.2493
R1004 B.n444 B.n134 33.2493
R1005 B.n521 B.n520 33.2493
R1006 B.n762 B.n761 33.2493
R1007 B.t1 B.n104 26.197
R1008 B.n500 B.t0 26.197
R1009 B.n128 B.t10 24.1819
R1010 B.t3 B.n773 24.1819
R1011 B B.n802 18.0485
R1012 B.n440 B.n130 10.6151
R1013 B.n450 B.n130 10.6151
R1014 B.n451 B.n450 10.6151
R1015 B.n452 B.n451 10.6151
R1016 B.n452 B.n122 10.6151
R1017 B.n462 B.n122 10.6151
R1018 B.n463 B.n462 10.6151
R1019 B.n464 B.n463 10.6151
R1020 B.n464 B.n114 10.6151
R1021 B.n474 B.n114 10.6151
R1022 B.n475 B.n474 10.6151
R1023 B.n476 B.n475 10.6151
R1024 B.n476 B.n106 10.6151
R1025 B.n487 B.n106 10.6151
R1026 B.n488 B.n487 10.6151
R1027 B.n489 B.n488 10.6151
R1028 B.n489 B.n0 10.6151
R1029 B.n439 B.n438 10.6151
R1030 B.n438 B.n138 10.6151
R1031 B.n433 B.n138 10.6151
R1032 B.n433 B.n432 10.6151
R1033 B.n432 B.n140 10.6151
R1034 B.n427 B.n140 10.6151
R1035 B.n427 B.n426 10.6151
R1036 B.n426 B.n425 10.6151
R1037 B.n425 B.n142 10.6151
R1038 B.n419 B.n142 10.6151
R1039 B.n419 B.n418 10.6151
R1040 B.n418 B.n417 10.6151
R1041 B.n417 B.n144 10.6151
R1042 B.n411 B.n144 10.6151
R1043 B.n411 B.n410 10.6151
R1044 B.n410 B.n409 10.6151
R1045 B.n409 B.n146 10.6151
R1046 B.n403 B.n146 10.6151
R1047 B.n403 B.n402 10.6151
R1048 B.n402 B.n401 10.6151
R1049 B.n401 B.n148 10.6151
R1050 B.n395 B.n148 10.6151
R1051 B.n395 B.n394 10.6151
R1052 B.n394 B.n393 10.6151
R1053 B.n393 B.n150 10.6151
R1054 B.n387 B.n150 10.6151
R1055 B.n387 B.n386 10.6151
R1056 B.n386 B.n385 10.6151
R1057 B.n385 B.n152 10.6151
R1058 B.n379 B.n152 10.6151
R1059 B.n379 B.n378 10.6151
R1060 B.n378 B.n377 10.6151
R1061 B.n377 B.n154 10.6151
R1062 B.n371 B.n154 10.6151
R1063 B.n371 B.n370 10.6151
R1064 B.n370 B.n369 10.6151
R1065 B.n369 B.n156 10.6151
R1066 B.n363 B.n156 10.6151
R1067 B.n363 B.n362 10.6151
R1068 B.n362 B.n361 10.6151
R1069 B.n361 B.n158 10.6151
R1070 B.n355 B.n158 10.6151
R1071 B.n355 B.n354 10.6151
R1072 B.n354 B.n353 10.6151
R1073 B.n353 B.n160 10.6151
R1074 B.n347 B.n160 10.6151
R1075 B.n347 B.n346 10.6151
R1076 B.n346 B.n345 10.6151
R1077 B.n345 B.n162 10.6151
R1078 B.n339 B.n162 10.6151
R1079 B.n339 B.n338 10.6151
R1080 B.n338 B.n337 10.6151
R1081 B.n337 B.n164 10.6151
R1082 B.n331 B.n164 10.6151
R1083 B.n329 B.n328 10.6151
R1084 B.n328 B.n168 10.6151
R1085 B.n322 B.n168 10.6151
R1086 B.n322 B.n321 10.6151
R1087 B.n321 B.n320 10.6151
R1088 B.n320 B.n170 10.6151
R1089 B.n314 B.n170 10.6151
R1090 B.n314 B.n313 10.6151
R1091 B.n313 B.n312 10.6151
R1092 B.n308 B.n307 10.6151
R1093 B.n307 B.n176 10.6151
R1094 B.n302 B.n176 10.6151
R1095 B.n302 B.n301 10.6151
R1096 B.n301 B.n300 10.6151
R1097 B.n300 B.n178 10.6151
R1098 B.n294 B.n178 10.6151
R1099 B.n294 B.n293 10.6151
R1100 B.n293 B.n292 10.6151
R1101 B.n292 B.n180 10.6151
R1102 B.n286 B.n180 10.6151
R1103 B.n286 B.n285 10.6151
R1104 B.n285 B.n284 10.6151
R1105 B.n284 B.n182 10.6151
R1106 B.n278 B.n182 10.6151
R1107 B.n278 B.n277 10.6151
R1108 B.n277 B.n276 10.6151
R1109 B.n276 B.n184 10.6151
R1110 B.n270 B.n184 10.6151
R1111 B.n270 B.n269 10.6151
R1112 B.n269 B.n268 10.6151
R1113 B.n268 B.n186 10.6151
R1114 B.n262 B.n186 10.6151
R1115 B.n262 B.n261 10.6151
R1116 B.n261 B.n260 10.6151
R1117 B.n260 B.n188 10.6151
R1118 B.n254 B.n188 10.6151
R1119 B.n254 B.n253 10.6151
R1120 B.n253 B.n252 10.6151
R1121 B.n252 B.n190 10.6151
R1122 B.n246 B.n190 10.6151
R1123 B.n246 B.n245 10.6151
R1124 B.n245 B.n244 10.6151
R1125 B.n244 B.n192 10.6151
R1126 B.n238 B.n192 10.6151
R1127 B.n238 B.n237 10.6151
R1128 B.n237 B.n236 10.6151
R1129 B.n236 B.n194 10.6151
R1130 B.n230 B.n194 10.6151
R1131 B.n230 B.n229 10.6151
R1132 B.n229 B.n228 10.6151
R1133 B.n228 B.n196 10.6151
R1134 B.n222 B.n196 10.6151
R1135 B.n222 B.n221 10.6151
R1136 B.n221 B.n220 10.6151
R1137 B.n220 B.n198 10.6151
R1138 B.n214 B.n198 10.6151
R1139 B.n214 B.n213 10.6151
R1140 B.n213 B.n212 10.6151
R1141 B.n212 B.n200 10.6151
R1142 B.n206 B.n200 10.6151
R1143 B.n206 B.n205 10.6151
R1144 B.n205 B.n204 10.6151
R1145 B.n204 B.n134 10.6151
R1146 B.n445 B.n444 10.6151
R1147 B.n446 B.n445 10.6151
R1148 B.n446 B.n125 10.6151
R1149 B.n456 B.n125 10.6151
R1150 B.n457 B.n456 10.6151
R1151 B.n458 B.n457 10.6151
R1152 B.n458 B.n118 10.6151
R1153 B.n468 B.n118 10.6151
R1154 B.n469 B.n468 10.6151
R1155 B.n470 B.n469 10.6151
R1156 B.n470 B.n110 10.6151
R1157 B.n480 B.n110 10.6151
R1158 B.n481 B.n480 10.6151
R1159 B.n483 B.n481 10.6151
R1160 B.n483 B.n482 10.6151
R1161 B.n482 B.n102 10.6151
R1162 B.n494 B.n102 10.6151
R1163 B.n495 B.n494 10.6151
R1164 B.n496 B.n495 10.6151
R1165 B.n497 B.n496 10.6151
R1166 B.n498 B.n497 10.6151
R1167 B.n502 B.n498 10.6151
R1168 B.n503 B.n502 10.6151
R1169 B.n504 B.n503 10.6151
R1170 B.n505 B.n504 10.6151
R1171 B.n507 B.n505 10.6151
R1172 B.n508 B.n507 10.6151
R1173 B.n509 B.n508 10.6151
R1174 B.n510 B.n509 10.6151
R1175 B.n512 B.n510 10.6151
R1176 B.n513 B.n512 10.6151
R1177 B.n514 B.n513 10.6151
R1178 B.n515 B.n514 10.6151
R1179 B.n517 B.n515 10.6151
R1180 B.n518 B.n517 10.6151
R1181 B.n519 B.n518 10.6151
R1182 B.n520 B.n519 10.6151
R1183 B.n794 B.n1 10.6151
R1184 B.n794 B.n793 10.6151
R1185 B.n793 B.n792 10.6151
R1186 B.n792 B.n10 10.6151
R1187 B.n786 B.n10 10.6151
R1188 B.n786 B.n785 10.6151
R1189 B.n785 B.n784 10.6151
R1190 B.n784 B.n17 10.6151
R1191 B.n778 B.n17 10.6151
R1192 B.n778 B.n777 10.6151
R1193 B.n777 B.n776 10.6151
R1194 B.n776 B.n24 10.6151
R1195 B.n770 B.n24 10.6151
R1196 B.n770 B.n769 10.6151
R1197 B.n769 B.n768 10.6151
R1198 B.n768 B.n31 10.6151
R1199 B.n762 B.n31 10.6151
R1200 B.n761 B.n760 10.6151
R1201 B.n760 B.n38 10.6151
R1202 B.n754 B.n38 10.6151
R1203 B.n754 B.n753 10.6151
R1204 B.n753 B.n752 10.6151
R1205 B.n752 B.n40 10.6151
R1206 B.n746 B.n40 10.6151
R1207 B.n746 B.n745 10.6151
R1208 B.n745 B.n744 10.6151
R1209 B.n744 B.n42 10.6151
R1210 B.n738 B.n42 10.6151
R1211 B.n738 B.n737 10.6151
R1212 B.n737 B.n736 10.6151
R1213 B.n736 B.n44 10.6151
R1214 B.n730 B.n44 10.6151
R1215 B.n730 B.n729 10.6151
R1216 B.n729 B.n728 10.6151
R1217 B.n728 B.n46 10.6151
R1218 B.n722 B.n46 10.6151
R1219 B.n722 B.n721 10.6151
R1220 B.n721 B.n720 10.6151
R1221 B.n720 B.n48 10.6151
R1222 B.n714 B.n48 10.6151
R1223 B.n714 B.n713 10.6151
R1224 B.n713 B.n712 10.6151
R1225 B.n712 B.n50 10.6151
R1226 B.n706 B.n50 10.6151
R1227 B.n706 B.n705 10.6151
R1228 B.n705 B.n704 10.6151
R1229 B.n704 B.n52 10.6151
R1230 B.n698 B.n52 10.6151
R1231 B.n698 B.n697 10.6151
R1232 B.n697 B.n696 10.6151
R1233 B.n696 B.n54 10.6151
R1234 B.n690 B.n54 10.6151
R1235 B.n690 B.n689 10.6151
R1236 B.n689 B.n688 10.6151
R1237 B.n688 B.n56 10.6151
R1238 B.n682 B.n56 10.6151
R1239 B.n682 B.n681 10.6151
R1240 B.n681 B.n680 10.6151
R1241 B.n680 B.n58 10.6151
R1242 B.n674 B.n58 10.6151
R1243 B.n674 B.n673 10.6151
R1244 B.n673 B.n672 10.6151
R1245 B.n672 B.n60 10.6151
R1246 B.n666 B.n60 10.6151
R1247 B.n666 B.n665 10.6151
R1248 B.n665 B.n664 10.6151
R1249 B.n664 B.n62 10.6151
R1250 B.n658 B.n62 10.6151
R1251 B.n658 B.n657 10.6151
R1252 B.n657 B.n656 10.6151
R1253 B.n656 B.n64 10.6151
R1254 B.n650 B.n649 10.6151
R1255 B.n649 B.n648 10.6151
R1256 B.n648 B.n69 10.6151
R1257 B.n642 B.n69 10.6151
R1258 B.n642 B.n641 10.6151
R1259 B.n641 B.n640 10.6151
R1260 B.n640 B.n71 10.6151
R1261 B.n634 B.n71 10.6151
R1262 B.n634 B.n633 10.6151
R1263 B.n631 B.n75 10.6151
R1264 B.n625 B.n75 10.6151
R1265 B.n625 B.n624 10.6151
R1266 B.n624 B.n623 10.6151
R1267 B.n623 B.n77 10.6151
R1268 B.n617 B.n77 10.6151
R1269 B.n617 B.n616 10.6151
R1270 B.n616 B.n615 10.6151
R1271 B.n615 B.n79 10.6151
R1272 B.n609 B.n79 10.6151
R1273 B.n609 B.n608 10.6151
R1274 B.n608 B.n607 10.6151
R1275 B.n607 B.n81 10.6151
R1276 B.n601 B.n81 10.6151
R1277 B.n601 B.n600 10.6151
R1278 B.n600 B.n599 10.6151
R1279 B.n599 B.n83 10.6151
R1280 B.n593 B.n83 10.6151
R1281 B.n593 B.n592 10.6151
R1282 B.n592 B.n591 10.6151
R1283 B.n591 B.n85 10.6151
R1284 B.n585 B.n85 10.6151
R1285 B.n585 B.n584 10.6151
R1286 B.n584 B.n583 10.6151
R1287 B.n583 B.n87 10.6151
R1288 B.n577 B.n87 10.6151
R1289 B.n577 B.n576 10.6151
R1290 B.n576 B.n575 10.6151
R1291 B.n575 B.n89 10.6151
R1292 B.n569 B.n89 10.6151
R1293 B.n569 B.n568 10.6151
R1294 B.n568 B.n567 10.6151
R1295 B.n567 B.n91 10.6151
R1296 B.n561 B.n91 10.6151
R1297 B.n561 B.n560 10.6151
R1298 B.n560 B.n559 10.6151
R1299 B.n559 B.n93 10.6151
R1300 B.n553 B.n93 10.6151
R1301 B.n553 B.n552 10.6151
R1302 B.n552 B.n551 10.6151
R1303 B.n551 B.n95 10.6151
R1304 B.n545 B.n95 10.6151
R1305 B.n545 B.n544 10.6151
R1306 B.n544 B.n543 10.6151
R1307 B.n543 B.n97 10.6151
R1308 B.n537 B.n97 10.6151
R1309 B.n537 B.n536 10.6151
R1310 B.n536 B.n535 10.6151
R1311 B.n535 B.n99 10.6151
R1312 B.n529 B.n99 10.6151
R1313 B.n529 B.n528 10.6151
R1314 B.n528 B.n527 10.6151
R1315 B.n527 B.n101 10.6151
R1316 B.n521 B.n101 10.6151
R1317 B.n460 B.t10 10.0761
R1318 B.n774 B.t3 10.0761
R1319 B.n331 B.n330 9.36635
R1320 B.n308 B.n174 9.36635
R1321 B.n68 B.n64 9.36635
R1322 B.n632 B.n631 9.36635
R1323 B.n802 B.n0 8.11757
R1324 B.n802 B.n1 8.11757
R1325 B.n485 B.t1 8.06095
R1326 B.n790 B.t0 8.06095
R1327 B.n330 B.n329 1.24928
R1328 B.n312 B.n174 1.24928
R1329 B.n650 B.n68 1.24928
R1330 B.n633 B.n632 1.24928
R1331 VP.n0 VP.t1 421.947
R1332 VP.n0 VP.t0 376.805
R1333 VP VP.n0 0.146778
R1334 VTAIL.n1 VTAIL.t1 47.5938
R1335 VTAIL.n3 VTAIL.t0 47.5935
R1336 VTAIL.n0 VTAIL.t2 47.5935
R1337 VTAIL.n2 VTAIL.t3 47.5935
R1338 VTAIL.n1 VTAIL.n0 29.7634
R1339 VTAIL.n3 VTAIL.n2 28.2031
R1340 VTAIL.n2 VTAIL.n1 1.2505
R1341 VTAIL VTAIL.n0 0.918603
R1342 VTAIL VTAIL.n3 0.332397
R1343 VDD1 VDD1.t1 106.243
R1344 VDD1 VDD1.t0 64.7206
R1345 VN VN.t0 422.233
R1346 VN VN.t1 376.952
R1347 VDD2.n0 VDD2.t0 105.329
R1348 VDD2.n0 VDD2.t1 64.2723
R1349 VDD2 VDD2.n0 0.448776
C0 VN VTAIL 2.74479f
C1 VN VDD1 0.147942f
C2 VDD2 VN 3.34498f
C3 VDD1 VTAIL 6.4272f
C4 VP VN 5.76983f
C5 VDD2 VTAIL 6.46688f
C6 VDD2 VDD1 0.5448f
C7 VP VTAIL 2.75933f
C8 VP VDD1 3.47955f
C9 VDD2 VP 0.287008f
C10 VDD2 B 4.856751f
C11 VDD1 B 8.09708f
C12 VTAIL B 8.566923f
C13 VN B 10.714609f
C14 VP B 5.303075f
C15 VDD2.t0 B 3.64203f
C16 VDD2.t1 B 3.04309f
C17 VDD2.n0 B 3.03506f
C18 VN.t1 B 3.07538f
C19 VN.t0 B 3.37655f
C20 VDD1.t0 B 3.05287f
C21 VDD1.t1 B 3.68256f
C22 VTAIL.t2 B 2.93263f
C23 VTAIL.n0 B 1.69594f
C24 VTAIL.t1 B 2.93263f
C25 VTAIL.n1 B 1.71709f
C26 VTAIL.t3 B 2.93263f
C27 VTAIL.n2 B 1.61764f
C28 VTAIL.t0 B 2.93263f
C29 VTAIL.n3 B 1.55912f
C30 VP.t1 B 3.47511f
C31 VP.t0 B 3.16866f
C32 VP.n0 B 5.41301f
.ends

