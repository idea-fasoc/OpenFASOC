* NGSPICE file created from diff_pair_sample_0737.ext - technology: sky130A

.subckt diff_pair_sample_0737 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=2.5179 ps=15.59 w=15.26 l=3.09
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=0 ps=0 w=15.26 l=3.09
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=0 ps=0 w=15.26 l=3.09
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=0 ps=0 w=15.26 l=3.09
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=0 ps=0 w=15.26 l=3.09
X5 VTAIL.t8 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=2.5179 ps=15.59 w=15.26 l=3.09
X6 VTAIL.t10 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=2.5179 ps=15.59 w=15.26 l=3.09
X7 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=5.9514 ps=31.3 w=15.26 l=3.09
X8 VTAIL.t6 VN.t3 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=2.5179 ps=15.59 w=15.26 l=3.09
X9 VDD1.t4 VP.t1 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=5.9514 ps=31.3 w=15.26 l=3.09
X10 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=2.5179 ps=15.59 w=15.26 l=3.09
X11 VDD1.t2 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=2.5179 ps=15.59 w=15.26 l=3.09
X12 VTAIL.t1 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=2.5179 ps=15.59 w=15.26 l=3.09
X13 VDD2.t1 VN.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9514 pd=31.3 as=2.5179 ps=15.59 w=15.26 l=3.09
X14 VDD2.t0 VN.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=5.9514 ps=31.3 w=15.26 l=3.09
X15 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5179 pd=15.59 as=5.9514 ps=31.3 w=15.26 l=3.09
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t2 152.507
R13 VN.n4 VN.t0 152.507
R14 VN.n5 VN.t1 119.019
R15 VN.n0 VN.t5 119.019
R16 VN.n21 VN.t3 119.019
R17 VN.n16 VN.t4 119.019
R18 VN.n15 VN.n0 69.5884
R19 VN.n31 VN.n16 69.5884
R20 VN.n11 VN.n2 56.5617
R21 VN.n27 VN.n18 56.5617
R22 VN VN.n31 53.3845
R23 VN.n5 VN.n4 49.5351
R24 VN.n21 VN.n20 49.5351
R25 VN.n6 VN.n5 24.5923
R26 VN.n7 VN.n6 24.5923
R27 VN.n7 VN.n2 24.5923
R28 VN.n12 VN.n11 24.5923
R29 VN.n13 VN.n12 24.5923
R30 VN.n23 VN.n18 24.5923
R31 VN.n23 VN.n22 24.5923
R32 VN.n22 VN.n21 24.5923
R33 VN.n29 VN.n28 24.5923
R34 VN.n28 VN.n27 24.5923
R35 VN.n13 VN.n0 20.6576
R36 VN.n29 VN.n16 20.6576
R37 VN.n4 VN.n3 3.87331
R38 VN.n20 VN.n19 3.87331
R39 VN.n31 VN.n30 0.354861
R40 VN.n15 VN.n14 0.354861
R41 VN VN.n15 0.267071
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n10 VTAIL.t11 43.9539
R53 VTAIL.n7 VTAIL.t5 43.9538
R54 VTAIL.n11 VTAIL.t9 43.9537
R55 VTAIL.n2 VTAIL.t3 43.9537
R56 VTAIL.n9 VTAIL.n8 42.6564
R57 VTAIL.n6 VTAIL.n5 42.6564
R58 VTAIL.n1 VTAIL.n0 42.6561
R59 VTAIL.n4 VTAIL.n3 42.6561
R60 VTAIL.n6 VTAIL.n4 31.4186
R61 VTAIL.n11 VTAIL.n10 28.4703
R62 VTAIL.n7 VTAIL.n6 2.94878
R63 VTAIL.n10 VTAIL.n9 2.94878
R64 VTAIL.n4 VTAIL.n2 2.94878
R65 VTAIL VTAIL.n11 2.15352
R66 VTAIL.n9 VTAIL.n7 1.94447
R67 VTAIL.n2 VTAIL.n1 1.94447
R68 VTAIL.n0 VTAIL.t4 1.29801
R69 VTAIL.n0 VTAIL.t8 1.29801
R70 VTAIL.n3 VTAIL.t2 1.29801
R71 VTAIL.n3 VTAIL.t10 1.29801
R72 VTAIL.n8 VTAIL.t0 1.29801
R73 VTAIL.n8 VTAIL.t1 1.29801
R74 VTAIL.n5 VTAIL.t7 1.29801
R75 VTAIL.n5 VTAIL.t6 1.29801
R76 VTAIL VTAIL.n1 0.795759
R77 VDD2.n1 VDD2.t5 62.7883
R78 VDD2.n2 VDD2.t1 60.6326
R79 VDD2.n1 VDD2.n0 60.0167
R80 VDD2 VDD2.n3 60.014
R81 VDD2.n2 VDD2.n1 46.4524
R82 VDD2 VDD2.n2 2.2699
R83 VDD2.n3 VDD2.t2 1.29801
R84 VDD2.n3 VDD2.t3 1.29801
R85 VDD2.n0 VDD2.t4 1.29801
R86 VDD2.n0 VDD2.t0 1.29801
R87 B.n959 B.n958 585
R88 B.n371 B.n146 585
R89 B.n370 B.n369 585
R90 B.n368 B.n367 585
R91 B.n366 B.n365 585
R92 B.n364 B.n363 585
R93 B.n362 B.n361 585
R94 B.n360 B.n359 585
R95 B.n358 B.n357 585
R96 B.n356 B.n355 585
R97 B.n354 B.n353 585
R98 B.n352 B.n351 585
R99 B.n350 B.n349 585
R100 B.n348 B.n347 585
R101 B.n346 B.n345 585
R102 B.n344 B.n343 585
R103 B.n342 B.n341 585
R104 B.n340 B.n339 585
R105 B.n338 B.n337 585
R106 B.n336 B.n335 585
R107 B.n334 B.n333 585
R108 B.n332 B.n331 585
R109 B.n330 B.n329 585
R110 B.n328 B.n327 585
R111 B.n326 B.n325 585
R112 B.n324 B.n323 585
R113 B.n322 B.n321 585
R114 B.n320 B.n319 585
R115 B.n318 B.n317 585
R116 B.n316 B.n315 585
R117 B.n314 B.n313 585
R118 B.n312 B.n311 585
R119 B.n310 B.n309 585
R120 B.n308 B.n307 585
R121 B.n306 B.n305 585
R122 B.n304 B.n303 585
R123 B.n302 B.n301 585
R124 B.n300 B.n299 585
R125 B.n298 B.n297 585
R126 B.n296 B.n295 585
R127 B.n294 B.n293 585
R128 B.n292 B.n291 585
R129 B.n290 B.n289 585
R130 B.n288 B.n287 585
R131 B.n286 B.n285 585
R132 B.n284 B.n283 585
R133 B.n282 B.n281 585
R134 B.n280 B.n279 585
R135 B.n278 B.n277 585
R136 B.n276 B.n275 585
R137 B.n274 B.n273 585
R138 B.n271 B.n270 585
R139 B.n269 B.n268 585
R140 B.n267 B.n266 585
R141 B.n265 B.n264 585
R142 B.n263 B.n262 585
R143 B.n261 B.n260 585
R144 B.n259 B.n258 585
R145 B.n257 B.n256 585
R146 B.n255 B.n254 585
R147 B.n253 B.n252 585
R148 B.n250 B.n249 585
R149 B.n248 B.n247 585
R150 B.n246 B.n245 585
R151 B.n244 B.n243 585
R152 B.n242 B.n241 585
R153 B.n240 B.n239 585
R154 B.n238 B.n237 585
R155 B.n236 B.n235 585
R156 B.n234 B.n233 585
R157 B.n232 B.n231 585
R158 B.n230 B.n229 585
R159 B.n228 B.n227 585
R160 B.n226 B.n225 585
R161 B.n224 B.n223 585
R162 B.n222 B.n221 585
R163 B.n220 B.n219 585
R164 B.n218 B.n217 585
R165 B.n216 B.n215 585
R166 B.n214 B.n213 585
R167 B.n212 B.n211 585
R168 B.n210 B.n209 585
R169 B.n208 B.n207 585
R170 B.n206 B.n205 585
R171 B.n204 B.n203 585
R172 B.n202 B.n201 585
R173 B.n200 B.n199 585
R174 B.n198 B.n197 585
R175 B.n196 B.n195 585
R176 B.n194 B.n193 585
R177 B.n192 B.n191 585
R178 B.n190 B.n189 585
R179 B.n188 B.n187 585
R180 B.n186 B.n185 585
R181 B.n184 B.n183 585
R182 B.n182 B.n181 585
R183 B.n180 B.n179 585
R184 B.n178 B.n177 585
R185 B.n176 B.n175 585
R186 B.n174 B.n173 585
R187 B.n172 B.n171 585
R188 B.n170 B.n169 585
R189 B.n168 B.n167 585
R190 B.n166 B.n165 585
R191 B.n164 B.n163 585
R192 B.n162 B.n161 585
R193 B.n160 B.n159 585
R194 B.n158 B.n157 585
R195 B.n156 B.n155 585
R196 B.n154 B.n153 585
R197 B.n152 B.n151 585
R198 B.n89 B.n88 585
R199 B.n957 B.n90 585
R200 B.n962 B.n90 585
R201 B.n956 B.n955 585
R202 B.n955 B.n86 585
R203 B.n954 B.n85 585
R204 B.n968 B.n85 585
R205 B.n953 B.n84 585
R206 B.n969 B.n84 585
R207 B.n952 B.n83 585
R208 B.n970 B.n83 585
R209 B.n951 B.n950 585
R210 B.n950 B.n79 585
R211 B.n949 B.n78 585
R212 B.n976 B.n78 585
R213 B.n948 B.n77 585
R214 B.n977 B.n77 585
R215 B.n947 B.n76 585
R216 B.n978 B.n76 585
R217 B.n946 B.n945 585
R218 B.n945 B.n72 585
R219 B.n944 B.n71 585
R220 B.n984 B.n71 585
R221 B.n943 B.n70 585
R222 B.n985 B.n70 585
R223 B.n942 B.n69 585
R224 B.n986 B.n69 585
R225 B.n941 B.n940 585
R226 B.n940 B.n65 585
R227 B.n939 B.n64 585
R228 B.n992 B.n64 585
R229 B.n938 B.n63 585
R230 B.n993 B.n63 585
R231 B.n937 B.n62 585
R232 B.n994 B.n62 585
R233 B.n936 B.n935 585
R234 B.n935 B.n58 585
R235 B.n934 B.n57 585
R236 B.n1000 B.n57 585
R237 B.n933 B.n56 585
R238 B.n1001 B.n56 585
R239 B.n932 B.n55 585
R240 B.n1002 B.n55 585
R241 B.n931 B.n930 585
R242 B.n930 B.n54 585
R243 B.n929 B.n50 585
R244 B.n1008 B.n50 585
R245 B.n928 B.n49 585
R246 B.n1009 B.n49 585
R247 B.n927 B.n48 585
R248 B.n1010 B.n48 585
R249 B.n926 B.n925 585
R250 B.n925 B.n44 585
R251 B.n924 B.n43 585
R252 B.n1016 B.n43 585
R253 B.n923 B.n42 585
R254 B.n1017 B.n42 585
R255 B.n922 B.n41 585
R256 B.n1018 B.n41 585
R257 B.n921 B.n920 585
R258 B.n920 B.n37 585
R259 B.n919 B.n36 585
R260 B.n1024 B.n36 585
R261 B.n918 B.n35 585
R262 B.n1025 B.n35 585
R263 B.n917 B.n34 585
R264 B.n1026 B.n34 585
R265 B.n916 B.n915 585
R266 B.n915 B.n30 585
R267 B.n914 B.n29 585
R268 B.n1032 B.n29 585
R269 B.n913 B.n28 585
R270 B.n1033 B.n28 585
R271 B.n912 B.n27 585
R272 B.n1034 B.n27 585
R273 B.n911 B.n910 585
R274 B.n910 B.n23 585
R275 B.n909 B.n22 585
R276 B.n1040 B.n22 585
R277 B.n908 B.n21 585
R278 B.n1041 B.n21 585
R279 B.n907 B.n20 585
R280 B.n1042 B.n20 585
R281 B.n906 B.n905 585
R282 B.n905 B.n19 585
R283 B.n904 B.n15 585
R284 B.n1048 B.n15 585
R285 B.n903 B.n14 585
R286 B.n1049 B.n14 585
R287 B.n902 B.n13 585
R288 B.n1050 B.n13 585
R289 B.n901 B.n900 585
R290 B.n900 B.n12 585
R291 B.n899 B.n898 585
R292 B.n899 B.n8 585
R293 B.n897 B.n7 585
R294 B.n1057 B.n7 585
R295 B.n896 B.n6 585
R296 B.n1058 B.n6 585
R297 B.n895 B.n5 585
R298 B.n1059 B.n5 585
R299 B.n894 B.n893 585
R300 B.n893 B.n4 585
R301 B.n892 B.n372 585
R302 B.n892 B.n891 585
R303 B.n882 B.n373 585
R304 B.n374 B.n373 585
R305 B.n884 B.n883 585
R306 B.n885 B.n884 585
R307 B.n881 B.n379 585
R308 B.n379 B.n378 585
R309 B.n880 B.n879 585
R310 B.n879 B.n878 585
R311 B.n381 B.n380 585
R312 B.n871 B.n381 585
R313 B.n870 B.n869 585
R314 B.n872 B.n870 585
R315 B.n868 B.n386 585
R316 B.n386 B.n385 585
R317 B.n867 B.n866 585
R318 B.n866 B.n865 585
R319 B.n388 B.n387 585
R320 B.n389 B.n388 585
R321 B.n858 B.n857 585
R322 B.n859 B.n858 585
R323 B.n856 B.n394 585
R324 B.n394 B.n393 585
R325 B.n855 B.n854 585
R326 B.n854 B.n853 585
R327 B.n396 B.n395 585
R328 B.n397 B.n396 585
R329 B.n846 B.n845 585
R330 B.n847 B.n846 585
R331 B.n844 B.n401 585
R332 B.n405 B.n401 585
R333 B.n843 B.n842 585
R334 B.n842 B.n841 585
R335 B.n403 B.n402 585
R336 B.n404 B.n403 585
R337 B.n834 B.n833 585
R338 B.n835 B.n834 585
R339 B.n832 B.n410 585
R340 B.n410 B.n409 585
R341 B.n831 B.n830 585
R342 B.n830 B.n829 585
R343 B.n412 B.n411 585
R344 B.n413 B.n412 585
R345 B.n822 B.n821 585
R346 B.n823 B.n822 585
R347 B.n820 B.n418 585
R348 B.n418 B.n417 585
R349 B.n819 B.n818 585
R350 B.n818 B.n817 585
R351 B.n420 B.n419 585
R352 B.n810 B.n420 585
R353 B.n809 B.n808 585
R354 B.n811 B.n809 585
R355 B.n807 B.n425 585
R356 B.n425 B.n424 585
R357 B.n806 B.n805 585
R358 B.n805 B.n804 585
R359 B.n427 B.n426 585
R360 B.n428 B.n427 585
R361 B.n797 B.n796 585
R362 B.n798 B.n797 585
R363 B.n795 B.n433 585
R364 B.n433 B.n432 585
R365 B.n794 B.n793 585
R366 B.n793 B.n792 585
R367 B.n435 B.n434 585
R368 B.n436 B.n435 585
R369 B.n785 B.n784 585
R370 B.n786 B.n785 585
R371 B.n783 B.n441 585
R372 B.n441 B.n440 585
R373 B.n782 B.n781 585
R374 B.n781 B.n780 585
R375 B.n443 B.n442 585
R376 B.n444 B.n443 585
R377 B.n773 B.n772 585
R378 B.n774 B.n773 585
R379 B.n771 B.n449 585
R380 B.n449 B.n448 585
R381 B.n770 B.n769 585
R382 B.n769 B.n768 585
R383 B.n451 B.n450 585
R384 B.n452 B.n451 585
R385 B.n761 B.n760 585
R386 B.n762 B.n761 585
R387 B.n759 B.n457 585
R388 B.n457 B.n456 585
R389 B.n758 B.n757 585
R390 B.n757 B.n756 585
R391 B.n459 B.n458 585
R392 B.n460 B.n459 585
R393 B.n749 B.n748 585
R394 B.n750 B.n749 585
R395 B.n463 B.n462 585
R396 B.n528 B.n527 585
R397 B.n529 B.n525 585
R398 B.n525 B.n464 585
R399 B.n531 B.n530 585
R400 B.n533 B.n524 585
R401 B.n536 B.n535 585
R402 B.n537 B.n523 585
R403 B.n539 B.n538 585
R404 B.n541 B.n522 585
R405 B.n544 B.n543 585
R406 B.n545 B.n521 585
R407 B.n547 B.n546 585
R408 B.n549 B.n520 585
R409 B.n552 B.n551 585
R410 B.n553 B.n519 585
R411 B.n555 B.n554 585
R412 B.n557 B.n518 585
R413 B.n560 B.n559 585
R414 B.n561 B.n517 585
R415 B.n563 B.n562 585
R416 B.n565 B.n516 585
R417 B.n568 B.n567 585
R418 B.n569 B.n515 585
R419 B.n571 B.n570 585
R420 B.n573 B.n514 585
R421 B.n576 B.n575 585
R422 B.n577 B.n513 585
R423 B.n579 B.n578 585
R424 B.n581 B.n512 585
R425 B.n584 B.n583 585
R426 B.n585 B.n511 585
R427 B.n587 B.n586 585
R428 B.n589 B.n510 585
R429 B.n592 B.n591 585
R430 B.n593 B.n509 585
R431 B.n595 B.n594 585
R432 B.n597 B.n508 585
R433 B.n600 B.n599 585
R434 B.n601 B.n507 585
R435 B.n603 B.n602 585
R436 B.n605 B.n506 585
R437 B.n608 B.n607 585
R438 B.n609 B.n505 585
R439 B.n611 B.n610 585
R440 B.n613 B.n504 585
R441 B.n616 B.n615 585
R442 B.n617 B.n503 585
R443 B.n619 B.n618 585
R444 B.n621 B.n502 585
R445 B.n624 B.n623 585
R446 B.n625 B.n499 585
R447 B.n628 B.n627 585
R448 B.n630 B.n498 585
R449 B.n633 B.n632 585
R450 B.n634 B.n497 585
R451 B.n636 B.n635 585
R452 B.n638 B.n496 585
R453 B.n641 B.n640 585
R454 B.n642 B.n495 585
R455 B.n644 B.n643 585
R456 B.n646 B.n494 585
R457 B.n649 B.n648 585
R458 B.n650 B.n490 585
R459 B.n652 B.n651 585
R460 B.n654 B.n489 585
R461 B.n657 B.n656 585
R462 B.n658 B.n488 585
R463 B.n660 B.n659 585
R464 B.n662 B.n487 585
R465 B.n665 B.n664 585
R466 B.n666 B.n486 585
R467 B.n668 B.n667 585
R468 B.n670 B.n485 585
R469 B.n673 B.n672 585
R470 B.n674 B.n484 585
R471 B.n676 B.n675 585
R472 B.n678 B.n483 585
R473 B.n681 B.n680 585
R474 B.n682 B.n482 585
R475 B.n684 B.n683 585
R476 B.n686 B.n481 585
R477 B.n689 B.n688 585
R478 B.n690 B.n480 585
R479 B.n692 B.n691 585
R480 B.n694 B.n479 585
R481 B.n697 B.n696 585
R482 B.n698 B.n478 585
R483 B.n700 B.n699 585
R484 B.n702 B.n477 585
R485 B.n705 B.n704 585
R486 B.n706 B.n476 585
R487 B.n708 B.n707 585
R488 B.n710 B.n475 585
R489 B.n713 B.n712 585
R490 B.n714 B.n474 585
R491 B.n716 B.n715 585
R492 B.n718 B.n473 585
R493 B.n721 B.n720 585
R494 B.n722 B.n472 585
R495 B.n724 B.n723 585
R496 B.n726 B.n471 585
R497 B.n729 B.n728 585
R498 B.n730 B.n470 585
R499 B.n732 B.n731 585
R500 B.n734 B.n469 585
R501 B.n737 B.n736 585
R502 B.n738 B.n468 585
R503 B.n740 B.n739 585
R504 B.n742 B.n467 585
R505 B.n743 B.n466 585
R506 B.n746 B.n745 585
R507 B.n747 B.n465 585
R508 B.n465 B.n464 585
R509 B.n752 B.n751 585
R510 B.n751 B.n750 585
R511 B.n753 B.n461 585
R512 B.n461 B.n460 585
R513 B.n755 B.n754 585
R514 B.n756 B.n755 585
R515 B.n455 B.n454 585
R516 B.n456 B.n455 585
R517 B.n764 B.n763 585
R518 B.n763 B.n762 585
R519 B.n765 B.n453 585
R520 B.n453 B.n452 585
R521 B.n767 B.n766 585
R522 B.n768 B.n767 585
R523 B.n447 B.n446 585
R524 B.n448 B.n447 585
R525 B.n776 B.n775 585
R526 B.n775 B.n774 585
R527 B.n777 B.n445 585
R528 B.n445 B.n444 585
R529 B.n779 B.n778 585
R530 B.n780 B.n779 585
R531 B.n439 B.n438 585
R532 B.n440 B.n439 585
R533 B.n788 B.n787 585
R534 B.n787 B.n786 585
R535 B.n789 B.n437 585
R536 B.n437 B.n436 585
R537 B.n791 B.n790 585
R538 B.n792 B.n791 585
R539 B.n431 B.n430 585
R540 B.n432 B.n431 585
R541 B.n800 B.n799 585
R542 B.n799 B.n798 585
R543 B.n801 B.n429 585
R544 B.n429 B.n428 585
R545 B.n803 B.n802 585
R546 B.n804 B.n803 585
R547 B.n423 B.n422 585
R548 B.n424 B.n423 585
R549 B.n813 B.n812 585
R550 B.n812 B.n811 585
R551 B.n814 B.n421 585
R552 B.n810 B.n421 585
R553 B.n816 B.n815 585
R554 B.n817 B.n816 585
R555 B.n416 B.n415 585
R556 B.n417 B.n416 585
R557 B.n825 B.n824 585
R558 B.n824 B.n823 585
R559 B.n826 B.n414 585
R560 B.n414 B.n413 585
R561 B.n828 B.n827 585
R562 B.n829 B.n828 585
R563 B.n408 B.n407 585
R564 B.n409 B.n408 585
R565 B.n837 B.n836 585
R566 B.n836 B.n835 585
R567 B.n838 B.n406 585
R568 B.n406 B.n404 585
R569 B.n840 B.n839 585
R570 B.n841 B.n840 585
R571 B.n400 B.n399 585
R572 B.n405 B.n400 585
R573 B.n849 B.n848 585
R574 B.n848 B.n847 585
R575 B.n850 B.n398 585
R576 B.n398 B.n397 585
R577 B.n852 B.n851 585
R578 B.n853 B.n852 585
R579 B.n392 B.n391 585
R580 B.n393 B.n392 585
R581 B.n861 B.n860 585
R582 B.n860 B.n859 585
R583 B.n862 B.n390 585
R584 B.n390 B.n389 585
R585 B.n864 B.n863 585
R586 B.n865 B.n864 585
R587 B.n384 B.n383 585
R588 B.n385 B.n384 585
R589 B.n874 B.n873 585
R590 B.n873 B.n872 585
R591 B.n875 B.n382 585
R592 B.n871 B.n382 585
R593 B.n877 B.n876 585
R594 B.n878 B.n877 585
R595 B.n377 B.n376 585
R596 B.n378 B.n377 585
R597 B.n887 B.n886 585
R598 B.n886 B.n885 585
R599 B.n888 B.n375 585
R600 B.n375 B.n374 585
R601 B.n890 B.n889 585
R602 B.n891 B.n890 585
R603 B.n3 B.n0 585
R604 B.n4 B.n3 585
R605 B.n1056 B.n1 585
R606 B.n1057 B.n1056 585
R607 B.n1055 B.n1054 585
R608 B.n1055 B.n8 585
R609 B.n1053 B.n9 585
R610 B.n12 B.n9 585
R611 B.n1052 B.n1051 585
R612 B.n1051 B.n1050 585
R613 B.n11 B.n10 585
R614 B.n1049 B.n11 585
R615 B.n1047 B.n1046 585
R616 B.n1048 B.n1047 585
R617 B.n1045 B.n16 585
R618 B.n19 B.n16 585
R619 B.n1044 B.n1043 585
R620 B.n1043 B.n1042 585
R621 B.n18 B.n17 585
R622 B.n1041 B.n18 585
R623 B.n1039 B.n1038 585
R624 B.n1040 B.n1039 585
R625 B.n1037 B.n24 585
R626 B.n24 B.n23 585
R627 B.n1036 B.n1035 585
R628 B.n1035 B.n1034 585
R629 B.n26 B.n25 585
R630 B.n1033 B.n26 585
R631 B.n1031 B.n1030 585
R632 B.n1032 B.n1031 585
R633 B.n1029 B.n31 585
R634 B.n31 B.n30 585
R635 B.n1028 B.n1027 585
R636 B.n1027 B.n1026 585
R637 B.n33 B.n32 585
R638 B.n1025 B.n33 585
R639 B.n1023 B.n1022 585
R640 B.n1024 B.n1023 585
R641 B.n1021 B.n38 585
R642 B.n38 B.n37 585
R643 B.n1020 B.n1019 585
R644 B.n1019 B.n1018 585
R645 B.n40 B.n39 585
R646 B.n1017 B.n40 585
R647 B.n1015 B.n1014 585
R648 B.n1016 B.n1015 585
R649 B.n1013 B.n45 585
R650 B.n45 B.n44 585
R651 B.n1012 B.n1011 585
R652 B.n1011 B.n1010 585
R653 B.n47 B.n46 585
R654 B.n1009 B.n47 585
R655 B.n1007 B.n1006 585
R656 B.n1008 B.n1007 585
R657 B.n1005 B.n51 585
R658 B.n54 B.n51 585
R659 B.n1004 B.n1003 585
R660 B.n1003 B.n1002 585
R661 B.n53 B.n52 585
R662 B.n1001 B.n53 585
R663 B.n999 B.n998 585
R664 B.n1000 B.n999 585
R665 B.n997 B.n59 585
R666 B.n59 B.n58 585
R667 B.n996 B.n995 585
R668 B.n995 B.n994 585
R669 B.n61 B.n60 585
R670 B.n993 B.n61 585
R671 B.n991 B.n990 585
R672 B.n992 B.n991 585
R673 B.n989 B.n66 585
R674 B.n66 B.n65 585
R675 B.n988 B.n987 585
R676 B.n987 B.n986 585
R677 B.n68 B.n67 585
R678 B.n985 B.n68 585
R679 B.n983 B.n982 585
R680 B.n984 B.n983 585
R681 B.n981 B.n73 585
R682 B.n73 B.n72 585
R683 B.n980 B.n979 585
R684 B.n979 B.n978 585
R685 B.n75 B.n74 585
R686 B.n977 B.n75 585
R687 B.n975 B.n974 585
R688 B.n976 B.n975 585
R689 B.n973 B.n80 585
R690 B.n80 B.n79 585
R691 B.n972 B.n971 585
R692 B.n971 B.n970 585
R693 B.n82 B.n81 585
R694 B.n969 B.n82 585
R695 B.n967 B.n966 585
R696 B.n968 B.n967 585
R697 B.n965 B.n87 585
R698 B.n87 B.n86 585
R699 B.n964 B.n963 585
R700 B.n963 B.n962 585
R701 B.n1060 B.n1059 585
R702 B.n1058 B.n2 585
R703 B.n963 B.n89 473.281
R704 B.n959 B.n90 473.281
R705 B.n749 B.n465 473.281
R706 B.n751 B.n463 473.281
R707 B.n149 B.t17 327.702
R708 B.n147 B.t6 327.702
R709 B.n491 B.t14 327.702
R710 B.n500 B.t10 327.702
R711 B.n961 B.n960 256.663
R712 B.n961 B.n145 256.663
R713 B.n961 B.n144 256.663
R714 B.n961 B.n143 256.663
R715 B.n961 B.n142 256.663
R716 B.n961 B.n141 256.663
R717 B.n961 B.n140 256.663
R718 B.n961 B.n139 256.663
R719 B.n961 B.n138 256.663
R720 B.n961 B.n137 256.663
R721 B.n961 B.n136 256.663
R722 B.n961 B.n135 256.663
R723 B.n961 B.n134 256.663
R724 B.n961 B.n133 256.663
R725 B.n961 B.n132 256.663
R726 B.n961 B.n131 256.663
R727 B.n961 B.n130 256.663
R728 B.n961 B.n129 256.663
R729 B.n961 B.n128 256.663
R730 B.n961 B.n127 256.663
R731 B.n961 B.n126 256.663
R732 B.n961 B.n125 256.663
R733 B.n961 B.n124 256.663
R734 B.n961 B.n123 256.663
R735 B.n961 B.n122 256.663
R736 B.n961 B.n121 256.663
R737 B.n961 B.n120 256.663
R738 B.n961 B.n119 256.663
R739 B.n961 B.n118 256.663
R740 B.n961 B.n117 256.663
R741 B.n961 B.n116 256.663
R742 B.n961 B.n115 256.663
R743 B.n961 B.n114 256.663
R744 B.n961 B.n113 256.663
R745 B.n961 B.n112 256.663
R746 B.n961 B.n111 256.663
R747 B.n961 B.n110 256.663
R748 B.n961 B.n109 256.663
R749 B.n961 B.n108 256.663
R750 B.n961 B.n107 256.663
R751 B.n961 B.n106 256.663
R752 B.n961 B.n105 256.663
R753 B.n961 B.n104 256.663
R754 B.n961 B.n103 256.663
R755 B.n961 B.n102 256.663
R756 B.n961 B.n101 256.663
R757 B.n961 B.n100 256.663
R758 B.n961 B.n99 256.663
R759 B.n961 B.n98 256.663
R760 B.n961 B.n97 256.663
R761 B.n961 B.n96 256.663
R762 B.n961 B.n95 256.663
R763 B.n961 B.n94 256.663
R764 B.n961 B.n93 256.663
R765 B.n961 B.n92 256.663
R766 B.n961 B.n91 256.663
R767 B.n526 B.n464 256.663
R768 B.n532 B.n464 256.663
R769 B.n534 B.n464 256.663
R770 B.n540 B.n464 256.663
R771 B.n542 B.n464 256.663
R772 B.n548 B.n464 256.663
R773 B.n550 B.n464 256.663
R774 B.n556 B.n464 256.663
R775 B.n558 B.n464 256.663
R776 B.n564 B.n464 256.663
R777 B.n566 B.n464 256.663
R778 B.n572 B.n464 256.663
R779 B.n574 B.n464 256.663
R780 B.n580 B.n464 256.663
R781 B.n582 B.n464 256.663
R782 B.n588 B.n464 256.663
R783 B.n590 B.n464 256.663
R784 B.n596 B.n464 256.663
R785 B.n598 B.n464 256.663
R786 B.n604 B.n464 256.663
R787 B.n606 B.n464 256.663
R788 B.n612 B.n464 256.663
R789 B.n614 B.n464 256.663
R790 B.n620 B.n464 256.663
R791 B.n622 B.n464 256.663
R792 B.n629 B.n464 256.663
R793 B.n631 B.n464 256.663
R794 B.n637 B.n464 256.663
R795 B.n639 B.n464 256.663
R796 B.n645 B.n464 256.663
R797 B.n647 B.n464 256.663
R798 B.n653 B.n464 256.663
R799 B.n655 B.n464 256.663
R800 B.n661 B.n464 256.663
R801 B.n663 B.n464 256.663
R802 B.n669 B.n464 256.663
R803 B.n671 B.n464 256.663
R804 B.n677 B.n464 256.663
R805 B.n679 B.n464 256.663
R806 B.n685 B.n464 256.663
R807 B.n687 B.n464 256.663
R808 B.n693 B.n464 256.663
R809 B.n695 B.n464 256.663
R810 B.n701 B.n464 256.663
R811 B.n703 B.n464 256.663
R812 B.n709 B.n464 256.663
R813 B.n711 B.n464 256.663
R814 B.n717 B.n464 256.663
R815 B.n719 B.n464 256.663
R816 B.n725 B.n464 256.663
R817 B.n727 B.n464 256.663
R818 B.n733 B.n464 256.663
R819 B.n735 B.n464 256.663
R820 B.n741 B.n464 256.663
R821 B.n744 B.n464 256.663
R822 B.n1062 B.n1061 256.663
R823 B.n153 B.n152 163.367
R824 B.n157 B.n156 163.367
R825 B.n161 B.n160 163.367
R826 B.n165 B.n164 163.367
R827 B.n169 B.n168 163.367
R828 B.n173 B.n172 163.367
R829 B.n177 B.n176 163.367
R830 B.n181 B.n180 163.367
R831 B.n185 B.n184 163.367
R832 B.n189 B.n188 163.367
R833 B.n193 B.n192 163.367
R834 B.n197 B.n196 163.367
R835 B.n201 B.n200 163.367
R836 B.n205 B.n204 163.367
R837 B.n209 B.n208 163.367
R838 B.n213 B.n212 163.367
R839 B.n217 B.n216 163.367
R840 B.n221 B.n220 163.367
R841 B.n225 B.n224 163.367
R842 B.n229 B.n228 163.367
R843 B.n233 B.n232 163.367
R844 B.n237 B.n236 163.367
R845 B.n241 B.n240 163.367
R846 B.n245 B.n244 163.367
R847 B.n249 B.n248 163.367
R848 B.n254 B.n253 163.367
R849 B.n258 B.n257 163.367
R850 B.n262 B.n261 163.367
R851 B.n266 B.n265 163.367
R852 B.n270 B.n269 163.367
R853 B.n275 B.n274 163.367
R854 B.n279 B.n278 163.367
R855 B.n283 B.n282 163.367
R856 B.n287 B.n286 163.367
R857 B.n291 B.n290 163.367
R858 B.n295 B.n294 163.367
R859 B.n299 B.n298 163.367
R860 B.n303 B.n302 163.367
R861 B.n307 B.n306 163.367
R862 B.n311 B.n310 163.367
R863 B.n315 B.n314 163.367
R864 B.n319 B.n318 163.367
R865 B.n323 B.n322 163.367
R866 B.n327 B.n326 163.367
R867 B.n331 B.n330 163.367
R868 B.n335 B.n334 163.367
R869 B.n339 B.n338 163.367
R870 B.n343 B.n342 163.367
R871 B.n347 B.n346 163.367
R872 B.n351 B.n350 163.367
R873 B.n355 B.n354 163.367
R874 B.n359 B.n358 163.367
R875 B.n363 B.n362 163.367
R876 B.n367 B.n366 163.367
R877 B.n369 B.n146 163.367
R878 B.n749 B.n459 163.367
R879 B.n757 B.n459 163.367
R880 B.n757 B.n457 163.367
R881 B.n761 B.n457 163.367
R882 B.n761 B.n451 163.367
R883 B.n769 B.n451 163.367
R884 B.n769 B.n449 163.367
R885 B.n773 B.n449 163.367
R886 B.n773 B.n443 163.367
R887 B.n781 B.n443 163.367
R888 B.n781 B.n441 163.367
R889 B.n785 B.n441 163.367
R890 B.n785 B.n435 163.367
R891 B.n793 B.n435 163.367
R892 B.n793 B.n433 163.367
R893 B.n797 B.n433 163.367
R894 B.n797 B.n427 163.367
R895 B.n805 B.n427 163.367
R896 B.n805 B.n425 163.367
R897 B.n809 B.n425 163.367
R898 B.n809 B.n420 163.367
R899 B.n818 B.n420 163.367
R900 B.n818 B.n418 163.367
R901 B.n822 B.n418 163.367
R902 B.n822 B.n412 163.367
R903 B.n830 B.n412 163.367
R904 B.n830 B.n410 163.367
R905 B.n834 B.n410 163.367
R906 B.n834 B.n403 163.367
R907 B.n842 B.n403 163.367
R908 B.n842 B.n401 163.367
R909 B.n846 B.n401 163.367
R910 B.n846 B.n396 163.367
R911 B.n854 B.n396 163.367
R912 B.n854 B.n394 163.367
R913 B.n858 B.n394 163.367
R914 B.n858 B.n388 163.367
R915 B.n866 B.n388 163.367
R916 B.n866 B.n386 163.367
R917 B.n870 B.n386 163.367
R918 B.n870 B.n381 163.367
R919 B.n879 B.n381 163.367
R920 B.n879 B.n379 163.367
R921 B.n884 B.n379 163.367
R922 B.n884 B.n373 163.367
R923 B.n892 B.n373 163.367
R924 B.n893 B.n892 163.367
R925 B.n893 B.n5 163.367
R926 B.n6 B.n5 163.367
R927 B.n7 B.n6 163.367
R928 B.n899 B.n7 163.367
R929 B.n900 B.n899 163.367
R930 B.n900 B.n13 163.367
R931 B.n14 B.n13 163.367
R932 B.n15 B.n14 163.367
R933 B.n905 B.n15 163.367
R934 B.n905 B.n20 163.367
R935 B.n21 B.n20 163.367
R936 B.n22 B.n21 163.367
R937 B.n910 B.n22 163.367
R938 B.n910 B.n27 163.367
R939 B.n28 B.n27 163.367
R940 B.n29 B.n28 163.367
R941 B.n915 B.n29 163.367
R942 B.n915 B.n34 163.367
R943 B.n35 B.n34 163.367
R944 B.n36 B.n35 163.367
R945 B.n920 B.n36 163.367
R946 B.n920 B.n41 163.367
R947 B.n42 B.n41 163.367
R948 B.n43 B.n42 163.367
R949 B.n925 B.n43 163.367
R950 B.n925 B.n48 163.367
R951 B.n49 B.n48 163.367
R952 B.n50 B.n49 163.367
R953 B.n930 B.n50 163.367
R954 B.n930 B.n55 163.367
R955 B.n56 B.n55 163.367
R956 B.n57 B.n56 163.367
R957 B.n935 B.n57 163.367
R958 B.n935 B.n62 163.367
R959 B.n63 B.n62 163.367
R960 B.n64 B.n63 163.367
R961 B.n940 B.n64 163.367
R962 B.n940 B.n69 163.367
R963 B.n70 B.n69 163.367
R964 B.n71 B.n70 163.367
R965 B.n945 B.n71 163.367
R966 B.n945 B.n76 163.367
R967 B.n77 B.n76 163.367
R968 B.n78 B.n77 163.367
R969 B.n950 B.n78 163.367
R970 B.n950 B.n83 163.367
R971 B.n84 B.n83 163.367
R972 B.n85 B.n84 163.367
R973 B.n955 B.n85 163.367
R974 B.n955 B.n90 163.367
R975 B.n527 B.n525 163.367
R976 B.n531 B.n525 163.367
R977 B.n535 B.n533 163.367
R978 B.n539 B.n523 163.367
R979 B.n543 B.n541 163.367
R980 B.n547 B.n521 163.367
R981 B.n551 B.n549 163.367
R982 B.n555 B.n519 163.367
R983 B.n559 B.n557 163.367
R984 B.n563 B.n517 163.367
R985 B.n567 B.n565 163.367
R986 B.n571 B.n515 163.367
R987 B.n575 B.n573 163.367
R988 B.n579 B.n513 163.367
R989 B.n583 B.n581 163.367
R990 B.n587 B.n511 163.367
R991 B.n591 B.n589 163.367
R992 B.n595 B.n509 163.367
R993 B.n599 B.n597 163.367
R994 B.n603 B.n507 163.367
R995 B.n607 B.n605 163.367
R996 B.n611 B.n505 163.367
R997 B.n615 B.n613 163.367
R998 B.n619 B.n503 163.367
R999 B.n623 B.n621 163.367
R1000 B.n628 B.n499 163.367
R1001 B.n632 B.n630 163.367
R1002 B.n636 B.n497 163.367
R1003 B.n640 B.n638 163.367
R1004 B.n644 B.n495 163.367
R1005 B.n648 B.n646 163.367
R1006 B.n652 B.n490 163.367
R1007 B.n656 B.n654 163.367
R1008 B.n660 B.n488 163.367
R1009 B.n664 B.n662 163.367
R1010 B.n668 B.n486 163.367
R1011 B.n672 B.n670 163.367
R1012 B.n676 B.n484 163.367
R1013 B.n680 B.n678 163.367
R1014 B.n684 B.n482 163.367
R1015 B.n688 B.n686 163.367
R1016 B.n692 B.n480 163.367
R1017 B.n696 B.n694 163.367
R1018 B.n700 B.n478 163.367
R1019 B.n704 B.n702 163.367
R1020 B.n708 B.n476 163.367
R1021 B.n712 B.n710 163.367
R1022 B.n716 B.n474 163.367
R1023 B.n720 B.n718 163.367
R1024 B.n724 B.n472 163.367
R1025 B.n728 B.n726 163.367
R1026 B.n732 B.n470 163.367
R1027 B.n736 B.n734 163.367
R1028 B.n740 B.n468 163.367
R1029 B.n743 B.n742 163.367
R1030 B.n745 B.n465 163.367
R1031 B.n751 B.n461 163.367
R1032 B.n755 B.n461 163.367
R1033 B.n755 B.n455 163.367
R1034 B.n763 B.n455 163.367
R1035 B.n763 B.n453 163.367
R1036 B.n767 B.n453 163.367
R1037 B.n767 B.n447 163.367
R1038 B.n775 B.n447 163.367
R1039 B.n775 B.n445 163.367
R1040 B.n779 B.n445 163.367
R1041 B.n779 B.n439 163.367
R1042 B.n787 B.n439 163.367
R1043 B.n787 B.n437 163.367
R1044 B.n791 B.n437 163.367
R1045 B.n791 B.n431 163.367
R1046 B.n799 B.n431 163.367
R1047 B.n799 B.n429 163.367
R1048 B.n803 B.n429 163.367
R1049 B.n803 B.n423 163.367
R1050 B.n812 B.n423 163.367
R1051 B.n812 B.n421 163.367
R1052 B.n816 B.n421 163.367
R1053 B.n816 B.n416 163.367
R1054 B.n824 B.n416 163.367
R1055 B.n824 B.n414 163.367
R1056 B.n828 B.n414 163.367
R1057 B.n828 B.n408 163.367
R1058 B.n836 B.n408 163.367
R1059 B.n836 B.n406 163.367
R1060 B.n840 B.n406 163.367
R1061 B.n840 B.n400 163.367
R1062 B.n848 B.n400 163.367
R1063 B.n848 B.n398 163.367
R1064 B.n852 B.n398 163.367
R1065 B.n852 B.n392 163.367
R1066 B.n860 B.n392 163.367
R1067 B.n860 B.n390 163.367
R1068 B.n864 B.n390 163.367
R1069 B.n864 B.n384 163.367
R1070 B.n873 B.n384 163.367
R1071 B.n873 B.n382 163.367
R1072 B.n877 B.n382 163.367
R1073 B.n877 B.n377 163.367
R1074 B.n886 B.n377 163.367
R1075 B.n886 B.n375 163.367
R1076 B.n890 B.n375 163.367
R1077 B.n890 B.n3 163.367
R1078 B.n1060 B.n3 163.367
R1079 B.n1056 B.n2 163.367
R1080 B.n1056 B.n1055 163.367
R1081 B.n1055 B.n9 163.367
R1082 B.n1051 B.n9 163.367
R1083 B.n1051 B.n11 163.367
R1084 B.n1047 B.n11 163.367
R1085 B.n1047 B.n16 163.367
R1086 B.n1043 B.n16 163.367
R1087 B.n1043 B.n18 163.367
R1088 B.n1039 B.n18 163.367
R1089 B.n1039 B.n24 163.367
R1090 B.n1035 B.n24 163.367
R1091 B.n1035 B.n26 163.367
R1092 B.n1031 B.n26 163.367
R1093 B.n1031 B.n31 163.367
R1094 B.n1027 B.n31 163.367
R1095 B.n1027 B.n33 163.367
R1096 B.n1023 B.n33 163.367
R1097 B.n1023 B.n38 163.367
R1098 B.n1019 B.n38 163.367
R1099 B.n1019 B.n40 163.367
R1100 B.n1015 B.n40 163.367
R1101 B.n1015 B.n45 163.367
R1102 B.n1011 B.n45 163.367
R1103 B.n1011 B.n47 163.367
R1104 B.n1007 B.n47 163.367
R1105 B.n1007 B.n51 163.367
R1106 B.n1003 B.n51 163.367
R1107 B.n1003 B.n53 163.367
R1108 B.n999 B.n53 163.367
R1109 B.n999 B.n59 163.367
R1110 B.n995 B.n59 163.367
R1111 B.n995 B.n61 163.367
R1112 B.n991 B.n61 163.367
R1113 B.n991 B.n66 163.367
R1114 B.n987 B.n66 163.367
R1115 B.n987 B.n68 163.367
R1116 B.n983 B.n68 163.367
R1117 B.n983 B.n73 163.367
R1118 B.n979 B.n73 163.367
R1119 B.n979 B.n75 163.367
R1120 B.n975 B.n75 163.367
R1121 B.n975 B.n80 163.367
R1122 B.n971 B.n80 163.367
R1123 B.n971 B.n82 163.367
R1124 B.n967 B.n82 163.367
R1125 B.n967 B.n87 163.367
R1126 B.n963 B.n87 163.367
R1127 B.n147 B.t8 139.588
R1128 B.n491 B.t16 139.588
R1129 B.n149 B.t18 139.567
R1130 B.n500 B.t13 139.567
R1131 B.n148 B.t9 73.2601
R1132 B.n492 B.t15 73.2601
R1133 B.n150 B.t19 73.2404
R1134 B.n501 B.t12 73.2404
R1135 B.n91 B.n89 71.676
R1136 B.n153 B.n92 71.676
R1137 B.n157 B.n93 71.676
R1138 B.n161 B.n94 71.676
R1139 B.n165 B.n95 71.676
R1140 B.n169 B.n96 71.676
R1141 B.n173 B.n97 71.676
R1142 B.n177 B.n98 71.676
R1143 B.n181 B.n99 71.676
R1144 B.n185 B.n100 71.676
R1145 B.n189 B.n101 71.676
R1146 B.n193 B.n102 71.676
R1147 B.n197 B.n103 71.676
R1148 B.n201 B.n104 71.676
R1149 B.n205 B.n105 71.676
R1150 B.n209 B.n106 71.676
R1151 B.n213 B.n107 71.676
R1152 B.n217 B.n108 71.676
R1153 B.n221 B.n109 71.676
R1154 B.n225 B.n110 71.676
R1155 B.n229 B.n111 71.676
R1156 B.n233 B.n112 71.676
R1157 B.n237 B.n113 71.676
R1158 B.n241 B.n114 71.676
R1159 B.n245 B.n115 71.676
R1160 B.n249 B.n116 71.676
R1161 B.n254 B.n117 71.676
R1162 B.n258 B.n118 71.676
R1163 B.n262 B.n119 71.676
R1164 B.n266 B.n120 71.676
R1165 B.n270 B.n121 71.676
R1166 B.n275 B.n122 71.676
R1167 B.n279 B.n123 71.676
R1168 B.n283 B.n124 71.676
R1169 B.n287 B.n125 71.676
R1170 B.n291 B.n126 71.676
R1171 B.n295 B.n127 71.676
R1172 B.n299 B.n128 71.676
R1173 B.n303 B.n129 71.676
R1174 B.n307 B.n130 71.676
R1175 B.n311 B.n131 71.676
R1176 B.n315 B.n132 71.676
R1177 B.n319 B.n133 71.676
R1178 B.n323 B.n134 71.676
R1179 B.n327 B.n135 71.676
R1180 B.n331 B.n136 71.676
R1181 B.n335 B.n137 71.676
R1182 B.n339 B.n138 71.676
R1183 B.n343 B.n139 71.676
R1184 B.n347 B.n140 71.676
R1185 B.n351 B.n141 71.676
R1186 B.n355 B.n142 71.676
R1187 B.n359 B.n143 71.676
R1188 B.n363 B.n144 71.676
R1189 B.n367 B.n145 71.676
R1190 B.n960 B.n146 71.676
R1191 B.n960 B.n959 71.676
R1192 B.n369 B.n145 71.676
R1193 B.n366 B.n144 71.676
R1194 B.n362 B.n143 71.676
R1195 B.n358 B.n142 71.676
R1196 B.n354 B.n141 71.676
R1197 B.n350 B.n140 71.676
R1198 B.n346 B.n139 71.676
R1199 B.n342 B.n138 71.676
R1200 B.n338 B.n137 71.676
R1201 B.n334 B.n136 71.676
R1202 B.n330 B.n135 71.676
R1203 B.n326 B.n134 71.676
R1204 B.n322 B.n133 71.676
R1205 B.n318 B.n132 71.676
R1206 B.n314 B.n131 71.676
R1207 B.n310 B.n130 71.676
R1208 B.n306 B.n129 71.676
R1209 B.n302 B.n128 71.676
R1210 B.n298 B.n127 71.676
R1211 B.n294 B.n126 71.676
R1212 B.n290 B.n125 71.676
R1213 B.n286 B.n124 71.676
R1214 B.n282 B.n123 71.676
R1215 B.n278 B.n122 71.676
R1216 B.n274 B.n121 71.676
R1217 B.n269 B.n120 71.676
R1218 B.n265 B.n119 71.676
R1219 B.n261 B.n118 71.676
R1220 B.n257 B.n117 71.676
R1221 B.n253 B.n116 71.676
R1222 B.n248 B.n115 71.676
R1223 B.n244 B.n114 71.676
R1224 B.n240 B.n113 71.676
R1225 B.n236 B.n112 71.676
R1226 B.n232 B.n111 71.676
R1227 B.n228 B.n110 71.676
R1228 B.n224 B.n109 71.676
R1229 B.n220 B.n108 71.676
R1230 B.n216 B.n107 71.676
R1231 B.n212 B.n106 71.676
R1232 B.n208 B.n105 71.676
R1233 B.n204 B.n104 71.676
R1234 B.n200 B.n103 71.676
R1235 B.n196 B.n102 71.676
R1236 B.n192 B.n101 71.676
R1237 B.n188 B.n100 71.676
R1238 B.n184 B.n99 71.676
R1239 B.n180 B.n98 71.676
R1240 B.n176 B.n97 71.676
R1241 B.n172 B.n96 71.676
R1242 B.n168 B.n95 71.676
R1243 B.n164 B.n94 71.676
R1244 B.n160 B.n93 71.676
R1245 B.n156 B.n92 71.676
R1246 B.n152 B.n91 71.676
R1247 B.n526 B.n463 71.676
R1248 B.n532 B.n531 71.676
R1249 B.n535 B.n534 71.676
R1250 B.n540 B.n539 71.676
R1251 B.n543 B.n542 71.676
R1252 B.n548 B.n547 71.676
R1253 B.n551 B.n550 71.676
R1254 B.n556 B.n555 71.676
R1255 B.n559 B.n558 71.676
R1256 B.n564 B.n563 71.676
R1257 B.n567 B.n566 71.676
R1258 B.n572 B.n571 71.676
R1259 B.n575 B.n574 71.676
R1260 B.n580 B.n579 71.676
R1261 B.n583 B.n582 71.676
R1262 B.n588 B.n587 71.676
R1263 B.n591 B.n590 71.676
R1264 B.n596 B.n595 71.676
R1265 B.n599 B.n598 71.676
R1266 B.n604 B.n603 71.676
R1267 B.n607 B.n606 71.676
R1268 B.n612 B.n611 71.676
R1269 B.n615 B.n614 71.676
R1270 B.n620 B.n619 71.676
R1271 B.n623 B.n622 71.676
R1272 B.n629 B.n628 71.676
R1273 B.n632 B.n631 71.676
R1274 B.n637 B.n636 71.676
R1275 B.n640 B.n639 71.676
R1276 B.n645 B.n644 71.676
R1277 B.n648 B.n647 71.676
R1278 B.n653 B.n652 71.676
R1279 B.n656 B.n655 71.676
R1280 B.n661 B.n660 71.676
R1281 B.n664 B.n663 71.676
R1282 B.n669 B.n668 71.676
R1283 B.n672 B.n671 71.676
R1284 B.n677 B.n676 71.676
R1285 B.n680 B.n679 71.676
R1286 B.n685 B.n684 71.676
R1287 B.n688 B.n687 71.676
R1288 B.n693 B.n692 71.676
R1289 B.n696 B.n695 71.676
R1290 B.n701 B.n700 71.676
R1291 B.n704 B.n703 71.676
R1292 B.n709 B.n708 71.676
R1293 B.n712 B.n711 71.676
R1294 B.n717 B.n716 71.676
R1295 B.n720 B.n719 71.676
R1296 B.n725 B.n724 71.676
R1297 B.n728 B.n727 71.676
R1298 B.n733 B.n732 71.676
R1299 B.n736 B.n735 71.676
R1300 B.n741 B.n740 71.676
R1301 B.n744 B.n743 71.676
R1302 B.n527 B.n526 71.676
R1303 B.n533 B.n532 71.676
R1304 B.n534 B.n523 71.676
R1305 B.n541 B.n540 71.676
R1306 B.n542 B.n521 71.676
R1307 B.n549 B.n548 71.676
R1308 B.n550 B.n519 71.676
R1309 B.n557 B.n556 71.676
R1310 B.n558 B.n517 71.676
R1311 B.n565 B.n564 71.676
R1312 B.n566 B.n515 71.676
R1313 B.n573 B.n572 71.676
R1314 B.n574 B.n513 71.676
R1315 B.n581 B.n580 71.676
R1316 B.n582 B.n511 71.676
R1317 B.n589 B.n588 71.676
R1318 B.n590 B.n509 71.676
R1319 B.n597 B.n596 71.676
R1320 B.n598 B.n507 71.676
R1321 B.n605 B.n604 71.676
R1322 B.n606 B.n505 71.676
R1323 B.n613 B.n612 71.676
R1324 B.n614 B.n503 71.676
R1325 B.n621 B.n620 71.676
R1326 B.n622 B.n499 71.676
R1327 B.n630 B.n629 71.676
R1328 B.n631 B.n497 71.676
R1329 B.n638 B.n637 71.676
R1330 B.n639 B.n495 71.676
R1331 B.n646 B.n645 71.676
R1332 B.n647 B.n490 71.676
R1333 B.n654 B.n653 71.676
R1334 B.n655 B.n488 71.676
R1335 B.n662 B.n661 71.676
R1336 B.n663 B.n486 71.676
R1337 B.n670 B.n669 71.676
R1338 B.n671 B.n484 71.676
R1339 B.n678 B.n677 71.676
R1340 B.n679 B.n482 71.676
R1341 B.n686 B.n685 71.676
R1342 B.n687 B.n480 71.676
R1343 B.n694 B.n693 71.676
R1344 B.n695 B.n478 71.676
R1345 B.n702 B.n701 71.676
R1346 B.n703 B.n476 71.676
R1347 B.n710 B.n709 71.676
R1348 B.n711 B.n474 71.676
R1349 B.n718 B.n717 71.676
R1350 B.n719 B.n472 71.676
R1351 B.n726 B.n725 71.676
R1352 B.n727 B.n470 71.676
R1353 B.n734 B.n733 71.676
R1354 B.n735 B.n468 71.676
R1355 B.n742 B.n741 71.676
R1356 B.n745 B.n744 71.676
R1357 B.n1061 B.n1060 71.676
R1358 B.n1061 B.n2 71.676
R1359 B.n150 B.n149 66.3278
R1360 B.n148 B.n147 66.3278
R1361 B.n492 B.n491 66.3278
R1362 B.n501 B.n500 66.3278
R1363 B.n750 B.n464 60.5313
R1364 B.n962 B.n961 60.5313
R1365 B.n251 B.n150 59.5399
R1366 B.n272 B.n148 59.5399
R1367 B.n493 B.n492 59.5399
R1368 B.n626 B.n501 59.5399
R1369 B.n750 B.n460 36.4261
R1370 B.n756 B.n460 36.4261
R1371 B.n756 B.n456 36.4261
R1372 B.n762 B.n456 36.4261
R1373 B.n762 B.n452 36.4261
R1374 B.n768 B.n452 36.4261
R1375 B.n768 B.n448 36.4261
R1376 B.n774 B.n448 36.4261
R1377 B.n780 B.n444 36.4261
R1378 B.n780 B.n440 36.4261
R1379 B.n786 B.n440 36.4261
R1380 B.n786 B.n436 36.4261
R1381 B.n792 B.n436 36.4261
R1382 B.n792 B.n432 36.4261
R1383 B.n798 B.n432 36.4261
R1384 B.n798 B.n428 36.4261
R1385 B.n804 B.n428 36.4261
R1386 B.n804 B.n424 36.4261
R1387 B.n811 B.n424 36.4261
R1388 B.n811 B.n810 36.4261
R1389 B.n817 B.n417 36.4261
R1390 B.n823 B.n417 36.4261
R1391 B.n823 B.n413 36.4261
R1392 B.n829 B.n413 36.4261
R1393 B.n829 B.n409 36.4261
R1394 B.n835 B.n409 36.4261
R1395 B.n835 B.n404 36.4261
R1396 B.n841 B.n404 36.4261
R1397 B.n841 B.n405 36.4261
R1398 B.n847 B.n397 36.4261
R1399 B.n853 B.n397 36.4261
R1400 B.n853 B.n393 36.4261
R1401 B.n859 B.n393 36.4261
R1402 B.n859 B.n389 36.4261
R1403 B.n865 B.n389 36.4261
R1404 B.n865 B.n385 36.4261
R1405 B.n872 B.n385 36.4261
R1406 B.n872 B.n871 36.4261
R1407 B.n878 B.n378 36.4261
R1408 B.n885 B.n378 36.4261
R1409 B.n885 B.n374 36.4261
R1410 B.n891 B.n374 36.4261
R1411 B.n891 B.n4 36.4261
R1412 B.n1059 B.n4 36.4261
R1413 B.n1059 B.n1058 36.4261
R1414 B.n1058 B.n1057 36.4261
R1415 B.n1057 B.n8 36.4261
R1416 B.n12 B.n8 36.4261
R1417 B.n1050 B.n12 36.4261
R1418 B.n1050 B.n1049 36.4261
R1419 B.n1049 B.n1048 36.4261
R1420 B.n1042 B.n19 36.4261
R1421 B.n1042 B.n1041 36.4261
R1422 B.n1041 B.n1040 36.4261
R1423 B.n1040 B.n23 36.4261
R1424 B.n1034 B.n23 36.4261
R1425 B.n1034 B.n1033 36.4261
R1426 B.n1033 B.n1032 36.4261
R1427 B.n1032 B.n30 36.4261
R1428 B.n1026 B.n30 36.4261
R1429 B.n1025 B.n1024 36.4261
R1430 B.n1024 B.n37 36.4261
R1431 B.n1018 B.n37 36.4261
R1432 B.n1018 B.n1017 36.4261
R1433 B.n1017 B.n1016 36.4261
R1434 B.n1016 B.n44 36.4261
R1435 B.n1010 B.n44 36.4261
R1436 B.n1010 B.n1009 36.4261
R1437 B.n1009 B.n1008 36.4261
R1438 B.n1002 B.n54 36.4261
R1439 B.n1002 B.n1001 36.4261
R1440 B.n1001 B.n1000 36.4261
R1441 B.n1000 B.n58 36.4261
R1442 B.n994 B.n58 36.4261
R1443 B.n994 B.n993 36.4261
R1444 B.n993 B.n992 36.4261
R1445 B.n992 B.n65 36.4261
R1446 B.n986 B.n65 36.4261
R1447 B.n986 B.n985 36.4261
R1448 B.n985 B.n984 36.4261
R1449 B.n984 B.n72 36.4261
R1450 B.n978 B.n977 36.4261
R1451 B.n977 B.n976 36.4261
R1452 B.n976 B.n79 36.4261
R1453 B.n970 B.n79 36.4261
R1454 B.n970 B.n969 36.4261
R1455 B.n969 B.n968 36.4261
R1456 B.n968 B.n86 36.4261
R1457 B.n962 B.n86 36.4261
R1458 B.n871 B.t3 31.6051
R1459 B.n19 B.t0 31.6051
R1460 B.n752 B.n462 30.7517
R1461 B.n748 B.n747 30.7517
R1462 B.n958 B.n957 30.7517
R1463 B.n964 B.n88 30.7517
R1464 B.n405 B.t5 29.4624
R1465 B.t1 B.n1025 29.4624
R1466 B.n810 B.t2 27.3197
R1467 B.n54 B.t4 27.3197
R1468 B.t11 B.n444 18.749
R1469 B.t7 B.n72 18.749
R1470 B B.n1062 18.0485
R1471 B.n774 B.t11 17.6776
R1472 B.n978 B.t7 17.6776
R1473 B.n753 B.n752 10.6151
R1474 B.n754 B.n753 10.6151
R1475 B.n754 B.n454 10.6151
R1476 B.n764 B.n454 10.6151
R1477 B.n765 B.n764 10.6151
R1478 B.n766 B.n765 10.6151
R1479 B.n766 B.n446 10.6151
R1480 B.n776 B.n446 10.6151
R1481 B.n777 B.n776 10.6151
R1482 B.n778 B.n777 10.6151
R1483 B.n778 B.n438 10.6151
R1484 B.n788 B.n438 10.6151
R1485 B.n789 B.n788 10.6151
R1486 B.n790 B.n789 10.6151
R1487 B.n790 B.n430 10.6151
R1488 B.n800 B.n430 10.6151
R1489 B.n801 B.n800 10.6151
R1490 B.n802 B.n801 10.6151
R1491 B.n802 B.n422 10.6151
R1492 B.n813 B.n422 10.6151
R1493 B.n814 B.n813 10.6151
R1494 B.n815 B.n814 10.6151
R1495 B.n815 B.n415 10.6151
R1496 B.n825 B.n415 10.6151
R1497 B.n826 B.n825 10.6151
R1498 B.n827 B.n826 10.6151
R1499 B.n827 B.n407 10.6151
R1500 B.n837 B.n407 10.6151
R1501 B.n838 B.n837 10.6151
R1502 B.n839 B.n838 10.6151
R1503 B.n839 B.n399 10.6151
R1504 B.n849 B.n399 10.6151
R1505 B.n850 B.n849 10.6151
R1506 B.n851 B.n850 10.6151
R1507 B.n851 B.n391 10.6151
R1508 B.n861 B.n391 10.6151
R1509 B.n862 B.n861 10.6151
R1510 B.n863 B.n862 10.6151
R1511 B.n863 B.n383 10.6151
R1512 B.n874 B.n383 10.6151
R1513 B.n875 B.n874 10.6151
R1514 B.n876 B.n875 10.6151
R1515 B.n876 B.n376 10.6151
R1516 B.n887 B.n376 10.6151
R1517 B.n888 B.n887 10.6151
R1518 B.n889 B.n888 10.6151
R1519 B.n889 B.n0 10.6151
R1520 B.n528 B.n462 10.6151
R1521 B.n529 B.n528 10.6151
R1522 B.n530 B.n529 10.6151
R1523 B.n530 B.n524 10.6151
R1524 B.n536 B.n524 10.6151
R1525 B.n537 B.n536 10.6151
R1526 B.n538 B.n537 10.6151
R1527 B.n538 B.n522 10.6151
R1528 B.n544 B.n522 10.6151
R1529 B.n545 B.n544 10.6151
R1530 B.n546 B.n545 10.6151
R1531 B.n546 B.n520 10.6151
R1532 B.n552 B.n520 10.6151
R1533 B.n553 B.n552 10.6151
R1534 B.n554 B.n553 10.6151
R1535 B.n554 B.n518 10.6151
R1536 B.n560 B.n518 10.6151
R1537 B.n561 B.n560 10.6151
R1538 B.n562 B.n561 10.6151
R1539 B.n562 B.n516 10.6151
R1540 B.n568 B.n516 10.6151
R1541 B.n569 B.n568 10.6151
R1542 B.n570 B.n569 10.6151
R1543 B.n570 B.n514 10.6151
R1544 B.n576 B.n514 10.6151
R1545 B.n577 B.n576 10.6151
R1546 B.n578 B.n577 10.6151
R1547 B.n578 B.n512 10.6151
R1548 B.n584 B.n512 10.6151
R1549 B.n585 B.n584 10.6151
R1550 B.n586 B.n585 10.6151
R1551 B.n586 B.n510 10.6151
R1552 B.n592 B.n510 10.6151
R1553 B.n593 B.n592 10.6151
R1554 B.n594 B.n593 10.6151
R1555 B.n594 B.n508 10.6151
R1556 B.n600 B.n508 10.6151
R1557 B.n601 B.n600 10.6151
R1558 B.n602 B.n601 10.6151
R1559 B.n602 B.n506 10.6151
R1560 B.n608 B.n506 10.6151
R1561 B.n609 B.n608 10.6151
R1562 B.n610 B.n609 10.6151
R1563 B.n610 B.n504 10.6151
R1564 B.n616 B.n504 10.6151
R1565 B.n617 B.n616 10.6151
R1566 B.n618 B.n617 10.6151
R1567 B.n618 B.n502 10.6151
R1568 B.n624 B.n502 10.6151
R1569 B.n625 B.n624 10.6151
R1570 B.n627 B.n498 10.6151
R1571 B.n633 B.n498 10.6151
R1572 B.n634 B.n633 10.6151
R1573 B.n635 B.n634 10.6151
R1574 B.n635 B.n496 10.6151
R1575 B.n641 B.n496 10.6151
R1576 B.n642 B.n641 10.6151
R1577 B.n643 B.n642 10.6151
R1578 B.n643 B.n494 10.6151
R1579 B.n650 B.n649 10.6151
R1580 B.n651 B.n650 10.6151
R1581 B.n651 B.n489 10.6151
R1582 B.n657 B.n489 10.6151
R1583 B.n658 B.n657 10.6151
R1584 B.n659 B.n658 10.6151
R1585 B.n659 B.n487 10.6151
R1586 B.n665 B.n487 10.6151
R1587 B.n666 B.n665 10.6151
R1588 B.n667 B.n666 10.6151
R1589 B.n667 B.n485 10.6151
R1590 B.n673 B.n485 10.6151
R1591 B.n674 B.n673 10.6151
R1592 B.n675 B.n674 10.6151
R1593 B.n675 B.n483 10.6151
R1594 B.n681 B.n483 10.6151
R1595 B.n682 B.n681 10.6151
R1596 B.n683 B.n682 10.6151
R1597 B.n683 B.n481 10.6151
R1598 B.n689 B.n481 10.6151
R1599 B.n690 B.n689 10.6151
R1600 B.n691 B.n690 10.6151
R1601 B.n691 B.n479 10.6151
R1602 B.n697 B.n479 10.6151
R1603 B.n698 B.n697 10.6151
R1604 B.n699 B.n698 10.6151
R1605 B.n699 B.n477 10.6151
R1606 B.n705 B.n477 10.6151
R1607 B.n706 B.n705 10.6151
R1608 B.n707 B.n706 10.6151
R1609 B.n707 B.n475 10.6151
R1610 B.n713 B.n475 10.6151
R1611 B.n714 B.n713 10.6151
R1612 B.n715 B.n714 10.6151
R1613 B.n715 B.n473 10.6151
R1614 B.n721 B.n473 10.6151
R1615 B.n722 B.n721 10.6151
R1616 B.n723 B.n722 10.6151
R1617 B.n723 B.n471 10.6151
R1618 B.n729 B.n471 10.6151
R1619 B.n730 B.n729 10.6151
R1620 B.n731 B.n730 10.6151
R1621 B.n731 B.n469 10.6151
R1622 B.n737 B.n469 10.6151
R1623 B.n738 B.n737 10.6151
R1624 B.n739 B.n738 10.6151
R1625 B.n739 B.n467 10.6151
R1626 B.n467 B.n466 10.6151
R1627 B.n746 B.n466 10.6151
R1628 B.n747 B.n746 10.6151
R1629 B.n748 B.n458 10.6151
R1630 B.n758 B.n458 10.6151
R1631 B.n759 B.n758 10.6151
R1632 B.n760 B.n759 10.6151
R1633 B.n760 B.n450 10.6151
R1634 B.n770 B.n450 10.6151
R1635 B.n771 B.n770 10.6151
R1636 B.n772 B.n771 10.6151
R1637 B.n772 B.n442 10.6151
R1638 B.n782 B.n442 10.6151
R1639 B.n783 B.n782 10.6151
R1640 B.n784 B.n783 10.6151
R1641 B.n784 B.n434 10.6151
R1642 B.n794 B.n434 10.6151
R1643 B.n795 B.n794 10.6151
R1644 B.n796 B.n795 10.6151
R1645 B.n796 B.n426 10.6151
R1646 B.n806 B.n426 10.6151
R1647 B.n807 B.n806 10.6151
R1648 B.n808 B.n807 10.6151
R1649 B.n808 B.n419 10.6151
R1650 B.n819 B.n419 10.6151
R1651 B.n820 B.n819 10.6151
R1652 B.n821 B.n820 10.6151
R1653 B.n821 B.n411 10.6151
R1654 B.n831 B.n411 10.6151
R1655 B.n832 B.n831 10.6151
R1656 B.n833 B.n832 10.6151
R1657 B.n833 B.n402 10.6151
R1658 B.n843 B.n402 10.6151
R1659 B.n844 B.n843 10.6151
R1660 B.n845 B.n844 10.6151
R1661 B.n845 B.n395 10.6151
R1662 B.n855 B.n395 10.6151
R1663 B.n856 B.n855 10.6151
R1664 B.n857 B.n856 10.6151
R1665 B.n857 B.n387 10.6151
R1666 B.n867 B.n387 10.6151
R1667 B.n868 B.n867 10.6151
R1668 B.n869 B.n868 10.6151
R1669 B.n869 B.n380 10.6151
R1670 B.n880 B.n380 10.6151
R1671 B.n881 B.n880 10.6151
R1672 B.n883 B.n881 10.6151
R1673 B.n883 B.n882 10.6151
R1674 B.n882 B.n372 10.6151
R1675 B.n894 B.n372 10.6151
R1676 B.n895 B.n894 10.6151
R1677 B.n896 B.n895 10.6151
R1678 B.n897 B.n896 10.6151
R1679 B.n898 B.n897 10.6151
R1680 B.n901 B.n898 10.6151
R1681 B.n902 B.n901 10.6151
R1682 B.n903 B.n902 10.6151
R1683 B.n904 B.n903 10.6151
R1684 B.n906 B.n904 10.6151
R1685 B.n907 B.n906 10.6151
R1686 B.n908 B.n907 10.6151
R1687 B.n909 B.n908 10.6151
R1688 B.n911 B.n909 10.6151
R1689 B.n912 B.n911 10.6151
R1690 B.n913 B.n912 10.6151
R1691 B.n914 B.n913 10.6151
R1692 B.n916 B.n914 10.6151
R1693 B.n917 B.n916 10.6151
R1694 B.n918 B.n917 10.6151
R1695 B.n919 B.n918 10.6151
R1696 B.n921 B.n919 10.6151
R1697 B.n922 B.n921 10.6151
R1698 B.n923 B.n922 10.6151
R1699 B.n924 B.n923 10.6151
R1700 B.n926 B.n924 10.6151
R1701 B.n927 B.n926 10.6151
R1702 B.n928 B.n927 10.6151
R1703 B.n929 B.n928 10.6151
R1704 B.n931 B.n929 10.6151
R1705 B.n932 B.n931 10.6151
R1706 B.n933 B.n932 10.6151
R1707 B.n934 B.n933 10.6151
R1708 B.n936 B.n934 10.6151
R1709 B.n937 B.n936 10.6151
R1710 B.n938 B.n937 10.6151
R1711 B.n939 B.n938 10.6151
R1712 B.n941 B.n939 10.6151
R1713 B.n942 B.n941 10.6151
R1714 B.n943 B.n942 10.6151
R1715 B.n944 B.n943 10.6151
R1716 B.n946 B.n944 10.6151
R1717 B.n947 B.n946 10.6151
R1718 B.n948 B.n947 10.6151
R1719 B.n949 B.n948 10.6151
R1720 B.n951 B.n949 10.6151
R1721 B.n952 B.n951 10.6151
R1722 B.n953 B.n952 10.6151
R1723 B.n954 B.n953 10.6151
R1724 B.n956 B.n954 10.6151
R1725 B.n957 B.n956 10.6151
R1726 B.n1054 B.n1 10.6151
R1727 B.n1054 B.n1053 10.6151
R1728 B.n1053 B.n1052 10.6151
R1729 B.n1052 B.n10 10.6151
R1730 B.n1046 B.n10 10.6151
R1731 B.n1046 B.n1045 10.6151
R1732 B.n1045 B.n1044 10.6151
R1733 B.n1044 B.n17 10.6151
R1734 B.n1038 B.n17 10.6151
R1735 B.n1038 B.n1037 10.6151
R1736 B.n1037 B.n1036 10.6151
R1737 B.n1036 B.n25 10.6151
R1738 B.n1030 B.n25 10.6151
R1739 B.n1030 B.n1029 10.6151
R1740 B.n1029 B.n1028 10.6151
R1741 B.n1028 B.n32 10.6151
R1742 B.n1022 B.n32 10.6151
R1743 B.n1022 B.n1021 10.6151
R1744 B.n1021 B.n1020 10.6151
R1745 B.n1020 B.n39 10.6151
R1746 B.n1014 B.n39 10.6151
R1747 B.n1014 B.n1013 10.6151
R1748 B.n1013 B.n1012 10.6151
R1749 B.n1012 B.n46 10.6151
R1750 B.n1006 B.n46 10.6151
R1751 B.n1006 B.n1005 10.6151
R1752 B.n1005 B.n1004 10.6151
R1753 B.n1004 B.n52 10.6151
R1754 B.n998 B.n52 10.6151
R1755 B.n998 B.n997 10.6151
R1756 B.n997 B.n996 10.6151
R1757 B.n996 B.n60 10.6151
R1758 B.n990 B.n60 10.6151
R1759 B.n990 B.n989 10.6151
R1760 B.n989 B.n988 10.6151
R1761 B.n988 B.n67 10.6151
R1762 B.n982 B.n67 10.6151
R1763 B.n982 B.n981 10.6151
R1764 B.n981 B.n980 10.6151
R1765 B.n980 B.n74 10.6151
R1766 B.n974 B.n74 10.6151
R1767 B.n974 B.n973 10.6151
R1768 B.n973 B.n972 10.6151
R1769 B.n972 B.n81 10.6151
R1770 B.n966 B.n81 10.6151
R1771 B.n966 B.n965 10.6151
R1772 B.n965 B.n964 10.6151
R1773 B.n151 B.n88 10.6151
R1774 B.n154 B.n151 10.6151
R1775 B.n155 B.n154 10.6151
R1776 B.n158 B.n155 10.6151
R1777 B.n159 B.n158 10.6151
R1778 B.n162 B.n159 10.6151
R1779 B.n163 B.n162 10.6151
R1780 B.n166 B.n163 10.6151
R1781 B.n167 B.n166 10.6151
R1782 B.n170 B.n167 10.6151
R1783 B.n171 B.n170 10.6151
R1784 B.n174 B.n171 10.6151
R1785 B.n175 B.n174 10.6151
R1786 B.n178 B.n175 10.6151
R1787 B.n179 B.n178 10.6151
R1788 B.n182 B.n179 10.6151
R1789 B.n183 B.n182 10.6151
R1790 B.n186 B.n183 10.6151
R1791 B.n187 B.n186 10.6151
R1792 B.n190 B.n187 10.6151
R1793 B.n191 B.n190 10.6151
R1794 B.n194 B.n191 10.6151
R1795 B.n195 B.n194 10.6151
R1796 B.n198 B.n195 10.6151
R1797 B.n199 B.n198 10.6151
R1798 B.n202 B.n199 10.6151
R1799 B.n203 B.n202 10.6151
R1800 B.n206 B.n203 10.6151
R1801 B.n207 B.n206 10.6151
R1802 B.n210 B.n207 10.6151
R1803 B.n211 B.n210 10.6151
R1804 B.n214 B.n211 10.6151
R1805 B.n215 B.n214 10.6151
R1806 B.n218 B.n215 10.6151
R1807 B.n219 B.n218 10.6151
R1808 B.n222 B.n219 10.6151
R1809 B.n223 B.n222 10.6151
R1810 B.n226 B.n223 10.6151
R1811 B.n227 B.n226 10.6151
R1812 B.n230 B.n227 10.6151
R1813 B.n231 B.n230 10.6151
R1814 B.n234 B.n231 10.6151
R1815 B.n235 B.n234 10.6151
R1816 B.n238 B.n235 10.6151
R1817 B.n239 B.n238 10.6151
R1818 B.n242 B.n239 10.6151
R1819 B.n243 B.n242 10.6151
R1820 B.n246 B.n243 10.6151
R1821 B.n247 B.n246 10.6151
R1822 B.n250 B.n247 10.6151
R1823 B.n255 B.n252 10.6151
R1824 B.n256 B.n255 10.6151
R1825 B.n259 B.n256 10.6151
R1826 B.n260 B.n259 10.6151
R1827 B.n263 B.n260 10.6151
R1828 B.n264 B.n263 10.6151
R1829 B.n267 B.n264 10.6151
R1830 B.n268 B.n267 10.6151
R1831 B.n271 B.n268 10.6151
R1832 B.n276 B.n273 10.6151
R1833 B.n277 B.n276 10.6151
R1834 B.n280 B.n277 10.6151
R1835 B.n281 B.n280 10.6151
R1836 B.n284 B.n281 10.6151
R1837 B.n285 B.n284 10.6151
R1838 B.n288 B.n285 10.6151
R1839 B.n289 B.n288 10.6151
R1840 B.n292 B.n289 10.6151
R1841 B.n293 B.n292 10.6151
R1842 B.n296 B.n293 10.6151
R1843 B.n297 B.n296 10.6151
R1844 B.n300 B.n297 10.6151
R1845 B.n301 B.n300 10.6151
R1846 B.n304 B.n301 10.6151
R1847 B.n305 B.n304 10.6151
R1848 B.n308 B.n305 10.6151
R1849 B.n309 B.n308 10.6151
R1850 B.n312 B.n309 10.6151
R1851 B.n313 B.n312 10.6151
R1852 B.n316 B.n313 10.6151
R1853 B.n317 B.n316 10.6151
R1854 B.n320 B.n317 10.6151
R1855 B.n321 B.n320 10.6151
R1856 B.n324 B.n321 10.6151
R1857 B.n325 B.n324 10.6151
R1858 B.n328 B.n325 10.6151
R1859 B.n329 B.n328 10.6151
R1860 B.n332 B.n329 10.6151
R1861 B.n333 B.n332 10.6151
R1862 B.n336 B.n333 10.6151
R1863 B.n337 B.n336 10.6151
R1864 B.n340 B.n337 10.6151
R1865 B.n341 B.n340 10.6151
R1866 B.n344 B.n341 10.6151
R1867 B.n345 B.n344 10.6151
R1868 B.n348 B.n345 10.6151
R1869 B.n349 B.n348 10.6151
R1870 B.n352 B.n349 10.6151
R1871 B.n353 B.n352 10.6151
R1872 B.n356 B.n353 10.6151
R1873 B.n357 B.n356 10.6151
R1874 B.n360 B.n357 10.6151
R1875 B.n361 B.n360 10.6151
R1876 B.n364 B.n361 10.6151
R1877 B.n365 B.n364 10.6151
R1878 B.n368 B.n365 10.6151
R1879 B.n370 B.n368 10.6151
R1880 B.n371 B.n370 10.6151
R1881 B.n958 B.n371 10.6151
R1882 B.n626 B.n625 9.36635
R1883 B.n649 B.n493 9.36635
R1884 B.n251 B.n250 9.36635
R1885 B.n273 B.n272 9.36635
R1886 B.n817 B.t2 9.1069
R1887 B.n1008 B.t4 9.1069
R1888 B.n1062 B.n0 8.11757
R1889 B.n1062 B.n1 8.11757
R1890 B.n847 B.t5 6.96422
R1891 B.n1026 B.t1 6.96422
R1892 B.n878 B.t3 4.82154
R1893 B.n1048 B.t0 4.82154
R1894 B.n627 B.n626 1.24928
R1895 B.n494 B.n493 1.24928
R1896 B.n252 B.n251 1.24928
R1897 B.n272 B.n271 1.24928
R1898 VP.n13 VP.n10 161.3
R1899 VP.n15 VP.n14 161.3
R1900 VP.n16 VP.n9 161.3
R1901 VP.n18 VP.n17 161.3
R1902 VP.n19 VP.n8 161.3
R1903 VP.n21 VP.n20 161.3
R1904 VP.n44 VP.n43 161.3
R1905 VP.n42 VP.n1 161.3
R1906 VP.n41 VP.n40 161.3
R1907 VP.n39 VP.n2 161.3
R1908 VP.n38 VP.n37 161.3
R1909 VP.n36 VP.n3 161.3
R1910 VP.n35 VP.n34 161.3
R1911 VP.n33 VP.n4 161.3
R1912 VP.n32 VP.n31 161.3
R1913 VP.n30 VP.n5 161.3
R1914 VP.n29 VP.n28 161.3
R1915 VP.n27 VP.n6 161.3
R1916 VP.n26 VP.n25 161.3
R1917 VP.n11 VP.t3 152.507
R1918 VP.n35 VP.t0 119.019
R1919 VP.n24 VP.t2 119.019
R1920 VP.n0 VP.t5 119.019
R1921 VP.n12 VP.t4 119.019
R1922 VP.n7 VP.t1 119.019
R1923 VP.n24 VP.n23 69.5884
R1924 VP.n45 VP.n0 69.5884
R1925 VP.n22 VP.n7 69.5884
R1926 VP.n30 VP.n29 56.5617
R1927 VP.n41 VP.n2 56.5617
R1928 VP.n18 VP.n9 56.5617
R1929 VP.n23 VP.n22 53.2193
R1930 VP.n12 VP.n11 49.5352
R1931 VP.n25 VP.n6 24.5923
R1932 VP.n29 VP.n6 24.5923
R1933 VP.n31 VP.n30 24.5923
R1934 VP.n31 VP.n4 24.5923
R1935 VP.n35 VP.n4 24.5923
R1936 VP.n36 VP.n35 24.5923
R1937 VP.n37 VP.n36 24.5923
R1938 VP.n37 VP.n2 24.5923
R1939 VP.n42 VP.n41 24.5923
R1940 VP.n43 VP.n42 24.5923
R1941 VP.n19 VP.n18 24.5923
R1942 VP.n20 VP.n19 24.5923
R1943 VP.n13 VP.n12 24.5923
R1944 VP.n14 VP.n13 24.5923
R1945 VP.n14 VP.n9 24.5923
R1946 VP.n25 VP.n24 20.6576
R1947 VP.n43 VP.n0 20.6576
R1948 VP.n20 VP.n7 20.6576
R1949 VP.n11 VP.n10 3.87328
R1950 VP.n22 VP.n21 0.354861
R1951 VP.n26 VP.n23 0.354861
R1952 VP.n45 VP.n44 0.354861
R1953 VP VP.n45 0.267071
R1954 VP.n15 VP.n10 0.189894
R1955 VP.n16 VP.n15 0.189894
R1956 VP.n17 VP.n16 0.189894
R1957 VP.n17 VP.n8 0.189894
R1958 VP.n21 VP.n8 0.189894
R1959 VP.n27 VP.n26 0.189894
R1960 VP.n28 VP.n27 0.189894
R1961 VP.n28 VP.n5 0.189894
R1962 VP.n32 VP.n5 0.189894
R1963 VP.n33 VP.n32 0.189894
R1964 VP.n34 VP.n33 0.189894
R1965 VP.n34 VP.n3 0.189894
R1966 VP.n38 VP.n3 0.189894
R1967 VP.n39 VP.n38 0.189894
R1968 VP.n40 VP.n39 0.189894
R1969 VP.n40 VP.n1 0.189894
R1970 VP.n44 VP.n1 0.189894
R1971 VDD1 VDD1.t2 62.902
R1972 VDD1.n1 VDD1.t3 62.7883
R1973 VDD1.n1 VDD1.n0 60.0167
R1974 VDD1.n3 VDD1.n2 59.3352
R1975 VDD1.n3 VDD1.n1 48.5095
R1976 VDD1.n2 VDD1.t1 1.29801
R1977 VDD1.n2 VDD1.t4 1.29801
R1978 VDD1.n0 VDD1.t5 1.29801
R1979 VDD1.n0 VDD1.t0 1.29801
R1980 VDD1 VDD1.n3 0.679379
C0 VN VDD2 8.70636f
C1 VDD1 VN 0.151831f
C2 VDD1 VDD2 1.59901f
C3 VTAIL VN 8.83495f
C4 VTAIL VDD2 9.022571f
C5 VP VN 8.00148f
C6 VP VDD2 0.500512f
C7 VTAIL VDD1 8.96862f
C8 VP VDD1 9.05145f
C9 VP VTAIL 8.84924f
C10 VDD2 B 6.944101f
C11 VDD1 B 7.297412f
C12 VTAIL B 9.460544f
C13 VN B 14.58252f
C14 VP B 13.217898f
C15 VDD1.t2 B 3.0095f
C16 VDD1.t3 B 3.00851f
C17 VDD1.t5 B 0.26007f
C18 VDD1.t0 B 0.26007f
C19 VDD1.n0 B 2.35026f
C20 VDD1.n1 B 3.00021f
C21 VDD1.t1 B 0.26007f
C22 VDD1.t4 B 0.26007f
C23 VDD1.n2 B 2.3452f
C24 VDD1.n3 B 2.74549f
C25 VP.t5 B 2.64583f
C26 VP.n0 B 1.00366f
C27 VP.n1 B 0.020469f
C28 VP.n2 B 0.02749f
C29 VP.n3 B 0.020469f
C30 VP.t0 B 2.64583f
C31 VP.n4 B 0.037958f
C32 VP.n5 B 0.020469f
C33 VP.n6 B 0.037958f
C34 VP.t1 B 2.64583f
C35 VP.n7 B 1.00366f
C36 VP.n8 B 0.020469f
C37 VP.n9 B 0.02749f
C38 VP.n10 B 0.232806f
C39 VP.t4 B 2.64583f
C40 VP.t3 B 2.87976f
C41 VP.n11 B 0.9496f
C42 VP.n12 B 0.996821f
C43 VP.n13 B 0.037958f
C44 VP.n14 B 0.037958f
C45 VP.n15 B 0.020469f
C46 VP.n16 B 0.020469f
C47 VP.n17 B 0.020469f
C48 VP.n18 B 0.03202f
C49 VP.n19 B 0.037958f
C50 VP.n20 B 0.03496f
C51 VP.n21 B 0.033032f
C52 VP.n22 B 1.26551f
C53 VP.n23 B 1.27937f
C54 VP.t2 B 2.64583f
C55 VP.n24 B 1.00366f
C56 VP.n25 B 0.03496f
C57 VP.n26 B 0.033032f
C58 VP.n27 B 0.020469f
C59 VP.n28 B 0.020469f
C60 VP.n29 B 0.03202f
C61 VP.n30 B 0.02749f
C62 VP.n31 B 0.037958f
C63 VP.n32 B 0.020469f
C64 VP.n33 B 0.020469f
C65 VP.n34 B 0.020469f
C66 VP.n35 B 0.939597f
C67 VP.n36 B 0.037958f
C68 VP.n37 B 0.037958f
C69 VP.n38 B 0.020469f
C70 VP.n39 B 0.020469f
C71 VP.n40 B 0.020469f
C72 VP.n41 B 0.03202f
C73 VP.n42 B 0.037958f
C74 VP.n43 B 0.03496f
C75 VP.n44 B 0.033032f
C76 VP.n45 B 0.042638f
C77 VDD2.t5 B 2.95503f
C78 VDD2.t4 B 0.255447f
C79 VDD2.t0 B 0.255447f
C80 VDD2.n0 B 2.30848f
C81 VDD2.n1 B 2.82861f
C82 VDD2.t1 B 2.94145f
C83 VDD2.n2 B 2.70278f
C84 VDD2.t2 B 0.255447f
C85 VDD2.t3 B 0.255447f
C86 VDD2.n3 B 2.30846f
C87 VTAIL.t4 B 0.279237f
C88 VTAIL.t8 B 0.279237f
C89 VTAIL.n0 B 2.4424f
C90 VTAIL.n1 B 0.446421f
C91 VTAIL.t3 B 3.11761f
C92 VTAIL.n2 B 0.69341f
C93 VTAIL.t2 B 0.279237f
C94 VTAIL.t10 B 0.279237f
C95 VTAIL.n3 B 2.4424f
C96 VTAIL.n4 B 2.1981f
C97 VTAIL.t7 B 0.279237f
C98 VTAIL.t6 B 0.279237f
C99 VTAIL.n5 B 2.44241f
C100 VTAIL.n6 B 2.19809f
C101 VTAIL.t5 B 3.11763f
C102 VTAIL.n7 B 0.693393f
C103 VTAIL.t0 B 0.279237f
C104 VTAIL.t1 B 0.279237f
C105 VTAIL.n8 B 2.44241f
C106 VTAIL.n9 B 0.607059f
C107 VTAIL.t11 B 3.11762f
C108 VTAIL.n10 B 2.06444f
C109 VTAIL.t9 B 3.11761f
C110 VTAIL.n11 B 2.00512f
C111 VN.t5 B 2.60208f
C112 VN.n0 B 0.987064f
C113 VN.n1 B 0.020131f
C114 VN.n2 B 0.027035f
C115 VN.n3 B 0.228956f
C116 VN.t1 B 2.60208f
C117 VN.t0 B 2.83214f
C118 VN.n4 B 0.933896f
C119 VN.n5 B 0.980337f
C120 VN.n6 B 0.037331f
C121 VN.n7 B 0.037331f
C122 VN.n8 B 0.020131f
C123 VN.n9 B 0.020131f
C124 VN.n10 B 0.020131f
C125 VN.n11 B 0.031491f
C126 VN.n12 B 0.037331f
C127 VN.n13 B 0.034382f
C128 VN.n14 B 0.032485f
C129 VN.n15 B 0.041933f
C130 VN.t4 B 2.60208f
C131 VN.n16 B 0.987064f
C132 VN.n17 B 0.020131f
C133 VN.n18 B 0.027035f
C134 VN.n19 B 0.228956f
C135 VN.t3 B 2.60208f
C136 VN.t2 B 2.83214f
C137 VN.n20 B 0.933896f
C138 VN.n21 B 0.980337f
C139 VN.n22 B 0.037331f
C140 VN.n23 B 0.037331f
C141 VN.n24 B 0.020131f
C142 VN.n25 B 0.020131f
C143 VN.n26 B 0.020131f
C144 VN.n27 B 0.031491f
C145 VN.n28 B 0.037331f
C146 VN.n29 B 0.034382f
C147 VN.n30 B 0.032485f
C148 VN.n31 B 1.25264f
.ends

