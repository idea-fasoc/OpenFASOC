* NGSPICE file created from diff_pair_sample_1085.ext - technology: sky130A

.subckt diff_pair_sample_1085 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=2.38095 ps=14.76 w=14.43 l=0.52
X1 VDD1.t5 VP.t0 VTAIL.t11 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=5.6277 ps=29.64 w=14.43 l=0.52
X2 B.t11 B.t9 B.t10 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=0 ps=0 w=14.43 l=0.52
X3 B.t8 B.t6 B.t7 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=0 ps=0 w=14.43 l=0.52
X4 B.t5 B.t3 B.t4 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=0 ps=0 w=14.43 l=0.52
X5 VDD2.t4 VN.t1 VTAIL.t10 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=5.6277 ps=29.64 w=14.43 l=0.52
X6 B.t2 B.t0 B.t1 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=0 ps=0 w=14.43 l=0.52
X7 VDD2.t3 VN.t2 VTAIL.t9 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=2.38095 ps=14.76 w=14.43 l=0.52
X8 VTAIL.t8 VN.t3 VDD2.t2 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=2.38095 ps=14.76 w=14.43 l=0.52
X9 VTAIL.t6 VN.t4 VDD2.t1 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=2.38095 ps=14.76 w=14.43 l=0.52
X10 VTAIL.t0 VP.t1 VDD1.t4 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=2.38095 ps=14.76 w=14.43 l=0.52
X11 VDD1.t3 VP.t2 VTAIL.t3 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=2.38095 ps=14.76 w=14.43 l=0.52
X12 VDD1.t2 VP.t3 VTAIL.t1 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=5.6277 ps=29.64 w=14.43 l=0.52
X13 VDD2.t0 VN.t5 VTAIL.t5 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=5.6277 ps=29.64 w=14.43 l=0.52
X14 VDD1.t1 VP.t4 VTAIL.t2 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=5.6277 pd=29.64 as=2.38095 ps=14.76 w=14.43 l=0.52
X15 VTAIL.t4 VP.t5 VDD1.t0 w_n1650_n3854# sky130_fd_pr__pfet_01v8 ad=2.38095 pd=14.76 as=2.38095 ps=14.76 w=14.43 l=0.52
R0 VN.n0 VN.t0 771.605
R1 VN.n4 VN.t1 771.605
R2 VN.n1 VN.t4 744.784
R3 VN.n2 VN.t5 744.784
R4 VN.n5 VN.t3 744.784
R5 VN.n6 VN.t2 744.784
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 48.2005
R9 VN.n6 VN.n5 48.2005
R10 VN.n7 VN.n4 45.1367
R11 VN.n3 VN.n0 45.1367
R12 VN VN.n7 42.7259
R13 VN.n5 VN.n4 13.3799
R14 VN.n1 VN.n0 13.3799
R15 VN VN.n3 0.0516364
R16 VTAIL.n7 VTAIL.t10 59.5254
R17 VTAIL.n11 VTAIL.t5 59.5253
R18 VTAIL.n2 VTAIL.t11 59.5253
R19 VTAIL.n10 VTAIL.t1 59.5253
R20 VTAIL.n9 VTAIL.n8 57.2729
R21 VTAIL.n6 VTAIL.n5 57.2729
R22 VTAIL.n1 VTAIL.n0 57.2726
R23 VTAIL.n4 VTAIL.n3 57.2726
R24 VTAIL.n6 VTAIL.n4 26.2721
R25 VTAIL.n11 VTAIL.n10 25.5393
R26 VTAIL.n0 VTAIL.t7 2.2531
R27 VTAIL.n0 VTAIL.t6 2.2531
R28 VTAIL.n3 VTAIL.t2 2.2531
R29 VTAIL.n3 VTAIL.t0 2.2531
R30 VTAIL.n8 VTAIL.t3 2.2531
R31 VTAIL.n8 VTAIL.t4 2.2531
R32 VTAIL.n5 VTAIL.t9 2.2531
R33 VTAIL.n5 VTAIL.t8 2.2531
R34 VTAIL.n9 VTAIL.n7 0.836707
R35 VTAIL.n2 VTAIL.n1 0.836707
R36 VTAIL.n7 VTAIL.n6 0.733259
R37 VTAIL.n10 VTAIL.n9 0.733259
R38 VTAIL.n4 VTAIL.n2 0.733259
R39 VTAIL VTAIL.n11 0.491879
R40 VTAIL VTAIL.n1 0.241879
R41 VDD2.n1 VDD2.t5 76.6983
R42 VDD2.n2 VDD2.t3 76.2042
R43 VDD2.n1 VDD2.n0 74.0793
R44 VDD2 VDD2.n3 74.0765
R45 VDD2.n2 VDD2.n1 38.5364
R46 VDD2.n3 VDD2.t2 2.2531
R47 VDD2.n3 VDD2.t4 2.2531
R48 VDD2.n0 VDD2.t1 2.2531
R49 VDD2.n0 VDD2.t0 2.2531
R50 VDD2 VDD2.n2 0.608259
R51 VP.n1 VP.t2 771.605
R52 VP.n6 VP.t4 744.784
R53 VP.n7 VP.t1 744.784
R54 VP.n8 VP.t0 744.784
R55 VP.n3 VP.t3 744.784
R56 VP.n2 VP.t5 744.784
R57 VP.n9 VP.n8 161.3
R58 VP.n4 VP.n3 161.3
R59 VP.n6 VP.n5 161.3
R60 VP.n7 VP.n0 80.6037
R61 VP.n7 VP.n6 48.2005
R62 VP.n8 VP.n7 48.2005
R63 VP.n3 VP.n2 48.2005
R64 VP.n4 VP.n1 45.1367
R65 VP.n5 VP.n4 42.3452
R66 VP.n2 VP.n1 13.3799
R67 VP.n5 VP.n0 0.285035
R68 VP.n9 VP.n0 0.285035
R69 VP VP.n9 0.0516364
R70 VDD1 VDD1.t3 76.812
R71 VDD1.n1 VDD1.t1 76.6983
R72 VDD1.n1 VDD1.n0 74.0793
R73 VDD1.n3 VDD1.n2 73.9515
R74 VDD1.n3 VDD1.n1 39.4858
R75 VDD1.n2 VDD1.t0 2.2531
R76 VDD1.n2 VDD1.t2 2.2531
R77 VDD1.n0 VDD1.t4 2.2531
R78 VDD1.n0 VDD1.t5 2.2531
R79 VDD1 VDD1.n3 0.1255
R80 B.n112 B.t3 874.72
R81 B.n120 B.t9 874.72
R82 B.n36 B.t0 874.72
R83 B.n42 B.t6 874.72
R84 B.n398 B.n397 585
R85 B.n399 B.n68 585
R86 B.n401 B.n400 585
R87 B.n402 B.n67 585
R88 B.n404 B.n403 585
R89 B.n405 B.n66 585
R90 B.n407 B.n406 585
R91 B.n408 B.n65 585
R92 B.n410 B.n409 585
R93 B.n411 B.n64 585
R94 B.n413 B.n412 585
R95 B.n414 B.n63 585
R96 B.n416 B.n415 585
R97 B.n417 B.n62 585
R98 B.n419 B.n418 585
R99 B.n420 B.n61 585
R100 B.n422 B.n421 585
R101 B.n423 B.n60 585
R102 B.n425 B.n424 585
R103 B.n426 B.n59 585
R104 B.n428 B.n427 585
R105 B.n429 B.n58 585
R106 B.n431 B.n430 585
R107 B.n432 B.n57 585
R108 B.n434 B.n433 585
R109 B.n435 B.n56 585
R110 B.n437 B.n436 585
R111 B.n438 B.n55 585
R112 B.n440 B.n439 585
R113 B.n441 B.n54 585
R114 B.n443 B.n442 585
R115 B.n444 B.n53 585
R116 B.n446 B.n445 585
R117 B.n447 B.n52 585
R118 B.n449 B.n448 585
R119 B.n450 B.n51 585
R120 B.n452 B.n451 585
R121 B.n453 B.n50 585
R122 B.n455 B.n454 585
R123 B.n456 B.n49 585
R124 B.n458 B.n457 585
R125 B.n459 B.n48 585
R126 B.n461 B.n460 585
R127 B.n462 B.n47 585
R128 B.n464 B.n463 585
R129 B.n465 B.n46 585
R130 B.n467 B.n466 585
R131 B.n468 B.n45 585
R132 B.n470 B.n469 585
R133 B.n472 B.n471 585
R134 B.n473 B.n41 585
R135 B.n475 B.n474 585
R136 B.n476 B.n40 585
R137 B.n478 B.n477 585
R138 B.n479 B.n39 585
R139 B.n481 B.n480 585
R140 B.n482 B.n38 585
R141 B.n484 B.n483 585
R142 B.n486 B.n35 585
R143 B.n488 B.n487 585
R144 B.n489 B.n34 585
R145 B.n491 B.n490 585
R146 B.n492 B.n33 585
R147 B.n494 B.n493 585
R148 B.n495 B.n32 585
R149 B.n497 B.n496 585
R150 B.n498 B.n31 585
R151 B.n500 B.n499 585
R152 B.n501 B.n30 585
R153 B.n503 B.n502 585
R154 B.n504 B.n29 585
R155 B.n506 B.n505 585
R156 B.n507 B.n28 585
R157 B.n509 B.n508 585
R158 B.n510 B.n27 585
R159 B.n512 B.n511 585
R160 B.n513 B.n26 585
R161 B.n515 B.n514 585
R162 B.n516 B.n25 585
R163 B.n518 B.n517 585
R164 B.n519 B.n24 585
R165 B.n521 B.n520 585
R166 B.n522 B.n23 585
R167 B.n524 B.n523 585
R168 B.n525 B.n22 585
R169 B.n527 B.n526 585
R170 B.n528 B.n21 585
R171 B.n530 B.n529 585
R172 B.n531 B.n20 585
R173 B.n533 B.n532 585
R174 B.n534 B.n19 585
R175 B.n536 B.n535 585
R176 B.n537 B.n18 585
R177 B.n539 B.n538 585
R178 B.n540 B.n17 585
R179 B.n542 B.n541 585
R180 B.n543 B.n16 585
R181 B.n545 B.n544 585
R182 B.n546 B.n15 585
R183 B.n548 B.n547 585
R184 B.n549 B.n14 585
R185 B.n551 B.n550 585
R186 B.n552 B.n13 585
R187 B.n554 B.n553 585
R188 B.n555 B.n12 585
R189 B.n557 B.n556 585
R190 B.n558 B.n11 585
R191 B.n396 B.n69 585
R192 B.n395 B.n394 585
R193 B.n393 B.n70 585
R194 B.n392 B.n391 585
R195 B.n390 B.n71 585
R196 B.n389 B.n388 585
R197 B.n387 B.n72 585
R198 B.n386 B.n385 585
R199 B.n384 B.n73 585
R200 B.n383 B.n382 585
R201 B.n381 B.n74 585
R202 B.n380 B.n379 585
R203 B.n378 B.n75 585
R204 B.n377 B.n376 585
R205 B.n375 B.n76 585
R206 B.n374 B.n373 585
R207 B.n372 B.n77 585
R208 B.n371 B.n370 585
R209 B.n369 B.n78 585
R210 B.n368 B.n367 585
R211 B.n366 B.n79 585
R212 B.n365 B.n364 585
R213 B.n363 B.n80 585
R214 B.n362 B.n361 585
R215 B.n360 B.n81 585
R216 B.n359 B.n358 585
R217 B.n357 B.n82 585
R218 B.n356 B.n355 585
R219 B.n354 B.n83 585
R220 B.n353 B.n352 585
R221 B.n351 B.n84 585
R222 B.n350 B.n349 585
R223 B.n348 B.n85 585
R224 B.n347 B.n346 585
R225 B.n345 B.n86 585
R226 B.n344 B.n343 585
R227 B.n342 B.n87 585
R228 B.n180 B.n145 585
R229 B.n182 B.n181 585
R230 B.n183 B.n144 585
R231 B.n185 B.n184 585
R232 B.n186 B.n143 585
R233 B.n188 B.n187 585
R234 B.n189 B.n142 585
R235 B.n191 B.n190 585
R236 B.n192 B.n141 585
R237 B.n194 B.n193 585
R238 B.n195 B.n140 585
R239 B.n197 B.n196 585
R240 B.n198 B.n139 585
R241 B.n200 B.n199 585
R242 B.n201 B.n138 585
R243 B.n203 B.n202 585
R244 B.n204 B.n137 585
R245 B.n206 B.n205 585
R246 B.n207 B.n136 585
R247 B.n209 B.n208 585
R248 B.n210 B.n135 585
R249 B.n212 B.n211 585
R250 B.n213 B.n134 585
R251 B.n215 B.n214 585
R252 B.n216 B.n133 585
R253 B.n218 B.n217 585
R254 B.n219 B.n132 585
R255 B.n221 B.n220 585
R256 B.n222 B.n131 585
R257 B.n224 B.n223 585
R258 B.n225 B.n130 585
R259 B.n227 B.n226 585
R260 B.n228 B.n129 585
R261 B.n230 B.n229 585
R262 B.n231 B.n128 585
R263 B.n233 B.n232 585
R264 B.n234 B.n127 585
R265 B.n236 B.n235 585
R266 B.n237 B.n126 585
R267 B.n239 B.n238 585
R268 B.n240 B.n125 585
R269 B.n242 B.n241 585
R270 B.n243 B.n124 585
R271 B.n245 B.n244 585
R272 B.n246 B.n123 585
R273 B.n248 B.n247 585
R274 B.n249 B.n122 585
R275 B.n251 B.n250 585
R276 B.n252 B.n119 585
R277 B.n255 B.n254 585
R278 B.n256 B.n118 585
R279 B.n258 B.n257 585
R280 B.n259 B.n117 585
R281 B.n261 B.n260 585
R282 B.n262 B.n116 585
R283 B.n264 B.n263 585
R284 B.n265 B.n115 585
R285 B.n267 B.n266 585
R286 B.n269 B.n268 585
R287 B.n270 B.n111 585
R288 B.n272 B.n271 585
R289 B.n273 B.n110 585
R290 B.n275 B.n274 585
R291 B.n276 B.n109 585
R292 B.n278 B.n277 585
R293 B.n279 B.n108 585
R294 B.n281 B.n280 585
R295 B.n282 B.n107 585
R296 B.n284 B.n283 585
R297 B.n285 B.n106 585
R298 B.n287 B.n286 585
R299 B.n288 B.n105 585
R300 B.n290 B.n289 585
R301 B.n291 B.n104 585
R302 B.n293 B.n292 585
R303 B.n294 B.n103 585
R304 B.n296 B.n295 585
R305 B.n297 B.n102 585
R306 B.n299 B.n298 585
R307 B.n300 B.n101 585
R308 B.n302 B.n301 585
R309 B.n303 B.n100 585
R310 B.n305 B.n304 585
R311 B.n306 B.n99 585
R312 B.n308 B.n307 585
R313 B.n309 B.n98 585
R314 B.n311 B.n310 585
R315 B.n312 B.n97 585
R316 B.n314 B.n313 585
R317 B.n315 B.n96 585
R318 B.n317 B.n316 585
R319 B.n318 B.n95 585
R320 B.n320 B.n319 585
R321 B.n321 B.n94 585
R322 B.n323 B.n322 585
R323 B.n324 B.n93 585
R324 B.n326 B.n325 585
R325 B.n327 B.n92 585
R326 B.n329 B.n328 585
R327 B.n330 B.n91 585
R328 B.n332 B.n331 585
R329 B.n333 B.n90 585
R330 B.n335 B.n334 585
R331 B.n336 B.n89 585
R332 B.n338 B.n337 585
R333 B.n339 B.n88 585
R334 B.n341 B.n340 585
R335 B.n179 B.n178 585
R336 B.n177 B.n146 585
R337 B.n176 B.n175 585
R338 B.n174 B.n147 585
R339 B.n173 B.n172 585
R340 B.n171 B.n148 585
R341 B.n170 B.n169 585
R342 B.n168 B.n149 585
R343 B.n167 B.n166 585
R344 B.n165 B.n150 585
R345 B.n164 B.n163 585
R346 B.n162 B.n151 585
R347 B.n161 B.n160 585
R348 B.n159 B.n152 585
R349 B.n158 B.n157 585
R350 B.n156 B.n153 585
R351 B.n155 B.n154 585
R352 B.n2 B.n0 585
R353 B.n585 B.n1 585
R354 B.n584 B.n583 585
R355 B.n582 B.n3 585
R356 B.n581 B.n580 585
R357 B.n579 B.n4 585
R358 B.n578 B.n577 585
R359 B.n576 B.n5 585
R360 B.n575 B.n574 585
R361 B.n573 B.n6 585
R362 B.n572 B.n571 585
R363 B.n570 B.n7 585
R364 B.n569 B.n568 585
R365 B.n567 B.n8 585
R366 B.n566 B.n565 585
R367 B.n564 B.n9 585
R368 B.n563 B.n562 585
R369 B.n561 B.n10 585
R370 B.n560 B.n559 585
R371 B.n587 B.n586 585
R372 B.n178 B.n145 526.135
R373 B.n560 B.n11 526.135
R374 B.n340 B.n87 526.135
R375 B.n398 B.n69 526.135
R376 B.n178 B.n177 163.367
R377 B.n177 B.n176 163.367
R378 B.n176 B.n147 163.367
R379 B.n172 B.n147 163.367
R380 B.n172 B.n171 163.367
R381 B.n171 B.n170 163.367
R382 B.n170 B.n149 163.367
R383 B.n166 B.n149 163.367
R384 B.n166 B.n165 163.367
R385 B.n165 B.n164 163.367
R386 B.n164 B.n151 163.367
R387 B.n160 B.n151 163.367
R388 B.n160 B.n159 163.367
R389 B.n159 B.n158 163.367
R390 B.n158 B.n153 163.367
R391 B.n154 B.n153 163.367
R392 B.n154 B.n2 163.367
R393 B.n586 B.n2 163.367
R394 B.n586 B.n585 163.367
R395 B.n585 B.n584 163.367
R396 B.n584 B.n3 163.367
R397 B.n580 B.n3 163.367
R398 B.n580 B.n579 163.367
R399 B.n579 B.n578 163.367
R400 B.n578 B.n5 163.367
R401 B.n574 B.n5 163.367
R402 B.n574 B.n573 163.367
R403 B.n573 B.n572 163.367
R404 B.n572 B.n7 163.367
R405 B.n568 B.n7 163.367
R406 B.n568 B.n567 163.367
R407 B.n567 B.n566 163.367
R408 B.n566 B.n9 163.367
R409 B.n562 B.n9 163.367
R410 B.n562 B.n561 163.367
R411 B.n561 B.n560 163.367
R412 B.n182 B.n145 163.367
R413 B.n183 B.n182 163.367
R414 B.n184 B.n183 163.367
R415 B.n184 B.n143 163.367
R416 B.n188 B.n143 163.367
R417 B.n189 B.n188 163.367
R418 B.n190 B.n189 163.367
R419 B.n190 B.n141 163.367
R420 B.n194 B.n141 163.367
R421 B.n195 B.n194 163.367
R422 B.n196 B.n195 163.367
R423 B.n196 B.n139 163.367
R424 B.n200 B.n139 163.367
R425 B.n201 B.n200 163.367
R426 B.n202 B.n201 163.367
R427 B.n202 B.n137 163.367
R428 B.n206 B.n137 163.367
R429 B.n207 B.n206 163.367
R430 B.n208 B.n207 163.367
R431 B.n208 B.n135 163.367
R432 B.n212 B.n135 163.367
R433 B.n213 B.n212 163.367
R434 B.n214 B.n213 163.367
R435 B.n214 B.n133 163.367
R436 B.n218 B.n133 163.367
R437 B.n219 B.n218 163.367
R438 B.n220 B.n219 163.367
R439 B.n220 B.n131 163.367
R440 B.n224 B.n131 163.367
R441 B.n225 B.n224 163.367
R442 B.n226 B.n225 163.367
R443 B.n226 B.n129 163.367
R444 B.n230 B.n129 163.367
R445 B.n231 B.n230 163.367
R446 B.n232 B.n231 163.367
R447 B.n232 B.n127 163.367
R448 B.n236 B.n127 163.367
R449 B.n237 B.n236 163.367
R450 B.n238 B.n237 163.367
R451 B.n238 B.n125 163.367
R452 B.n242 B.n125 163.367
R453 B.n243 B.n242 163.367
R454 B.n244 B.n243 163.367
R455 B.n244 B.n123 163.367
R456 B.n248 B.n123 163.367
R457 B.n249 B.n248 163.367
R458 B.n250 B.n249 163.367
R459 B.n250 B.n119 163.367
R460 B.n255 B.n119 163.367
R461 B.n256 B.n255 163.367
R462 B.n257 B.n256 163.367
R463 B.n257 B.n117 163.367
R464 B.n261 B.n117 163.367
R465 B.n262 B.n261 163.367
R466 B.n263 B.n262 163.367
R467 B.n263 B.n115 163.367
R468 B.n267 B.n115 163.367
R469 B.n268 B.n267 163.367
R470 B.n268 B.n111 163.367
R471 B.n272 B.n111 163.367
R472 B.n273 B.n272 163.367
R473 B.n274 B.n273 163.367
R474 B.n274 B.n109 163.367
R475 B.n278 B.n109 163.367
R476 B.n279 B.n278 163.367
R477 B.n280 B.n279 163.367
R478 B.n280 B.n107 163.367
R479 B.n284 B.n107 163.367
R480 B.n285 B.n284 163.367
R481 B.n286 B.n285 163.367
R482 B.n286 B.n105 163.367
R483 B.n290 B.n105 163.367
R484 B.n291 B.n290 163.367
R485 B.n292 B.n291 163.367
R486 B.n292 B.n103 163.367
R487 B.n296 B.n103 163.367
R488 B.n297 B.n296 163.367
R489 B.n298 B.n297 163.367
R490 B.n298 B.n101 163.367
R491 B.n302 B.n101 163.367
R492 B.n303 B.n302 163.367
R493 B.n304 B.n303 163.367
R494 B.n304 B.n99 163.367
R495 B.n308 B.n99 163.367
R496 B.n309 B.n308 163.367
R497 B.n310 B.n309 163.367
R498 B.n310 B.n97 163.367
R499 B.n314 B.n97 163.367
R500 B.n315 B.n314 163.367
R501 B.n316 B.n315 163.367
R502 B.n316 B.n95 163.367
R503 B.n320 B.n95 163.367
R504 B.n321 B.n320 163.367
R505 B.n322 B.n321 163.367
R506 B.n322 B.n93 163.367
R507 B.n326 B.n93 163.367
R508 B.n327 B.n326 163.367
R509 B.n328 B.n327 163.367
R510 B.n328 B.n91 163.367
R511 B.n332 B.n91 163.367
R512 B.n333 B.n332 163.367
R513 B.n334 B.n333 163.367
R514 B.n334 B.n89 163.367
R515 B.n338 B.n89 163.367
R516 B.n339 B.n338 163.367
R517 B.n340 B.n339 163.367
R518 B.n344 B.n87 163.367
R519 B.n345 B.n344 163.367
R520 B.n346 B.n345 163.367
R521 B.n346 B.n85 163.367
R522 B.n350 B.n85 163.367
R523 B.n351 B.n350 163.367
R524 B.n352 B.n351 163.367
R525 B.n352 B.n83 163.367
R526 B.n356 B.n83 163.367
R527 B.n357 B.n356 163.367
R528 B.n358 B.n357 163.367
R529 B.n358 B.n81 163.367
R530 B.n362 B.n81 163.367
R531 B.n363 B.n362 163.367
R532 B.n364 B.n363 163.367
R533 B.n364 B.n79 163.367
R534 B.n368 B.n79 163.367
R535 B.n369 B.n368 163.367
R536 B.n370 B.n369 163.367
R537 B.n370 B.n77 163.367
R538 B.n374 B.n77 163.367
R539 B.n375 B.n374 163.367
R540 B.n376 B.n375 163.367
R541 B.n376 B.n75 163.367
R542 B.n380 B.n75 163.367
R543 B.n381 B.n380 163.367
R544 B.n382 B.n381 163.367
R545 B.n382 B.n73 163.367
R546 B.n386 B.n73 163.367
R547 B.n387 B.n386 163.367
R548 B.n388 B.n387 163.367
R549 B.n388 B.n71 163.367
R550 B.n392 B.n71 163.367
R551 B.n393 B.n392 163.367
R552 B.n394 B.n393 163.367
R553 B.n394 B.n69 163.367
R554 B.n556 B.n11 163.367
R555 B.n556 B.n555 163.367
R556 B.n555 B.n554 163.367
R557 B.n554 B.n13 163.367
R558 B.n550 B.n13 163.367
R559 B.n550 B.n549 163.367
R560 B.n549 B.n548 163.367
R561 B.n548 B.n15 163.367
R562 B.n544 B.n15 163.367
R563 B.n544 B.n543 163.367
R564 B.n543 B.n542 163.367
R565 B.n542 B.n17 163.367
R566 B.n538 B.n17 163.367
R567 B.n538 B.n537 163.367
R568 B.n537 B.n536 163.367
R569 B.n536 B.n19 163.367
R570 B.n532 B.n19 163.367
R571 B.n532 B.n531 163.367
R572 B.n531 B.n530 163.367
R573 B.n530 B.n21 163.367
R574 B.n526 B.n21 163.367
R575 B.n526 B.n525 163.367
R576 B.n525 B.n524 163.367
R577 B.n524 B.n23 163.367
R578 B.n520 B.n23 163.367
R579 B.n520 B.n519 163.367
R580 B.n519 B.n518 163.367
R581 B.n518 B.n25 163.367
R582 B.n514 B.n25 163.367
R583 B.n514 B.n513 163.367
R584 B.n513 B.n512 163.367
R585 B.n512 B.n27 163.367
R586 B.n508 B.n27 163.367
R587 B.n508 B.n507 163.367
R588 B.n507 B.n506 163.367
R589 B.n506 B.n29 163.367
R590 B.n502 B.n29 163.367
R591 B.n502 B.n501 163.367
R592 B.n501 B.n500 163.367
R593 B.n500 B.n31 163.367
R594 B.n496 B.n31 163.367
R595 B.n496 B.n495 163.367
R596 B.n495 B.n494 163.367
R597 B.n494 B.n33 163.367
R598 B.n490 B.n33 163.367
R599 B.n490 B.n489 163.367
R600 B.n489 B.n488 163.367
R601 B.n488 B.n35 163.367
R602 B.n483 B.n35 163.367
R603 B.n483 B.n482 163.367
R604 B.n482 B.n481 163.367
R605 B.n481 B.n39 163.367
R606 B.n477 B.n39 163.367
R607 B.n477 B.n476 163.367
R608 B.n476 B.n475 163.367
R609 B.n475 B.n41 163.367
R610 B.n471 B.n41 163.367
R611 B.n471 B.n470 163.367
R612 B.n470 B.n45 163.367
R613 B.n466 B.n45 163.367
R614 B.n466 B.n465 163.367
R615 B.n465 B.n464 163.367
R616 B.n464 B.n47 163.367
R617 B.n460 B.n47 163.367
R618 B.n460 B.n459 163.367
R619 B.n459 B.n458 163.367
R620 B.n458 B.n49 163.367
R621 B.n454 B.n49 163.367
R622 B.n454 B.n453 163.367
R623 B.n453 B.n452 163.367
R624 B.n452 B.n51 163.367
R625 B.n448 B.n51 163.367
R626 B.n448 B.n447 163.367
R627 B.n447 B.n446 163.367
R628 B.n446 B.n53 163.367
R629 B.n442 B.n53 163.367
R630 B.n442 B.n441 163.367
R631 B.n441 B.n440 163.367
R632 B.n440 B.n55 163.367
R633 B.n436 B.n55 163.367
R634 B.n436 B.n435 163.367
R635 B.n435 B.n434 163.367
R636 B.n434 B.n57 163.367
R637 B.n430 B.n57 163.367
R638 B.n430 B.n429 163.367
R639 B.n429 B.n428 163.367
R640 B.n428 B.n59 163.367
R641 B.n424 B.n59 163.367
R642 B.n424 B.n423 163.367
R643 B.n423 B.n422 163.367
R644 B.n422 B.n61 163.367
R645 B.n418 B.n61 163.367
R646 B.n418 B.n417 163.367
R647 B.n417 B.n416 163.367
R648 B.n416 B.n63 163.367
R649 B.n412 B.n63 163.367
R650 B.n412 B.n411 163.367
R651 B.n411 B.n410 163.367
R652 B.n410 B.n65 163.367
R653 B.n406 B.n65 163.367
R654 B.n406 B.n405 163.367
R655 B.n405 B.n404 163.367
R656 B.n404 B.n67 163.367
R657 B.n400 B.n67 163.367
R658 B.n400 B.n399 163.367
R659 B.n399 B.n398 163.367
R660 B.n112 B.t5 126.04
R661 B.n42 B.t7 126.04
R662 B.n120 B.t11 126.022
R663 B.n36 B.t1 126.022
R664 B.n113 B.t4 109.555
R665 B.n43 B.t8 109.555
R666 B.n121 B.t10 109.537
R667 B.n37 B.t2 109.537
R668 B.n114 B.n113 59.5399
R669 B.n253 B.n121 59.5399
R670 B.n485 B.n37 59.5399
R671 B.n44 B.n43 59.5399
R672 B.n559 B.n558 34.1859
R673 B.n397 B.n396 34.1859
R674 B.n342 B.n341 34.1859
R675 B.n180 B.n179 34.1859
R676 B B.n587 18.0485
R677 B.n113 B.n112 16.4853
R678 B.n121 B.n120 16.4853
R679 B.n37 B.n36 16.4853
R680 B.n43 B.n42 16.4853
R681 B.n558 B.n557 10.6151
R682 B.n557 B.n12 10.6151
R683 B.n553 B.n12 10.6151
R684 B.n553 B.n552 10.6151
R685 B.n552 B.n551 10.6151
R686 B.n551 B.n14 10.6151
R687 B.n547 B.n14 10.6151
R688 B.n547 B.n546 10.6151
R689 B.n546 B.n545 10.6151
R690 B.n545 B.n16 10.6151
R691 B.n541 B.n16 10.6151
R692 B.n541 B.n540 10.6151
R693 B.n540 B.n539 10.6151
R694 B.n539 B.n18 10.6151
R695 B.n535 B.n18 10.6151
R696 B.n535 B.n534 10.6151
R697 B.n534 B.n533 10.6151
R698 B.n533 B.n20 10.6151
R699 B.n529 B.n20 10.6151
R700 B.n529 B.n528 10.6151
R701 B.n528 B.n527 10.6151
R702 B.n527 B.n22 10.6151
R703 B.n523 B.n22 10.6151
R704 B.n523 B.n522 10.6151
R705 B.n522 B.n521 10.6151
R706 B.n521 B.n24 10.6151
R707 B.n517 B.n24 10.6151
R708 B.n517 B.n516 10.6151
R709 B.n516 B.n515 10.6151
R710 B.n515 B.n26 10.6151
R711 B.n511 B.n26 10.6151
R712 B.n511 B.n510 10.6151
R713 B.n510 B.n509 10.6151
R714 B.n509 B.n28 10.6151
R715 B.n505 B.n28 10.6151
R716 B.n505 B.n504 10.6151
R717 B.n504 B.n503 10.6151
R718 B.n503 B.n30 10.6151
R719 B.n499 B.n30 10.6151
R720 B.n499 B.n498 10.6151
R721 B.n498 B.n497 10.6151
R722 B.n497 B.n32 10.6151
R723 B.n493 B.n32 10.6151
R724 B.n493 B.n492 10.6151
R725 B.n492 B.n491 10.6151
R726 B.n491 B.n34 10.6151
R727 B.n487 B.n34 10.6151
R728 B.n487 B.n486 10.6151
R729 B.n484 B.n38 10.6151
R730 B.n480 B.n38 10.6151
R731 B.n480 B.n479 10.6151
R732 B.n479 B.n478 10.6151
R733 B.n478 B.n40 10.6151
R734 B.n474 B.n40 10.6151
R735 B.n474 B.n473 10.6151
R736 B.n473 B.n472 10.6151
R737 B.n469 B.n468 10.6151
R738 B.n468 B.n467 10.6151
R739 B.n467 B.n46 10.6151
R740 B.n463 B.n46 10.6151
R741 B.n463 B.n462 10.6151
R742 B.n462 B.n461 10.6151
R743 B.n461 B.n48 10.6151
R744 B.n457 B.n48 10.6151
R745 B.n457 B.n456 10.6151
R746 B.n456 B.n455 10.6151
R747 B.n455 B.n50 10.6151
R748 B.n451 B.n50 10.6151
R749 B.n451 B.n450 10.6151
R750 B.n450 B.n449 10.6151
R751 B.n449 B.n52 10.6151
R752 B.n445 B.n52 10.6151
R753 B.n445 B.n444 10.6151
R754 B.n444 B.n443 10.6151
R755 B.n443 B.n54 10.6151
R756 B.n439 B.n54 10.6151
R757 B.n439 B.n438 10.6151
R758 B.n438 B.n437 10.6151
R759 B.n437 B.n56 10.6151
R760 B.n433 B.n56 10.6151
R761 B.n433 B.n432 10.6151
R762 B.n432 B.n431 10.6151
R763 B.n431 B.n58 10.6151
R764 B.n427 B.n58 10.6151
R765 B.n427 B.n426 10.6151
R766 B.n426 B.n425 10.6151
R767 B.n425 B.n60 10.6151
R768 B.n421 B.n60 10.6151
R769 B.n421 B.n420 10.6151
R770 B.n420 B.n419 10.6151
R771 B.n419 B.n62 10.6151
R772 B.n415 B.n62 10.6151
R773 B.n415 B.n414 10.6151
R774 B.n414 B.n413 10.6151
R775 B.n413 B.n64 10.6151
R776 B.n409 B.n64 10.6151
R777 B.n409 B.n408 10.6151
R778 B.n408 B.n407 10.6151
R779 B.n407 B.n66 10.6151
R780 B.n403 B.n66 10.6151
R781 B.n403 B.n402 10.6151
R782 B.n402 B.n401 10.6151
R783 B.n401 B.n68 10.6151
R784 B.n397 B.n68 10.6151
R785 B.n343 B.n342 10.6151
R786 B.n343 B.n86 10.6151
R787 B.n347 B.n86 10.6151
R788 B.n348 B.n347 10.6151
R789 B.n349 B.n348 10.6151
R790 B.n349 B.n84 10.6151
R791 B.n353 B.n84 10.6151
R792 B.n354 B.n353 10.6151
R793 B.n355 B.n354 10.6151
R794 B.n355 B.n82 10.6151
R795 B.n359 B.n82 10.6151
R796 B.n360 B.n359 10.6151
R797 B.n361 B.n360 10.6151
R798 B.n361 B.n80 10.6151
R799 B.n365 B.n80 10.6151
R800 B.n366 B.n365 10.6151
R801 B.n367 B.n366 10.6151
R802 B.n367 B.n78 10.6151
R803 B.n371 B.n78 10.6151
R804 B.n372 B.n371 10.6151
R805 B.n373 B.n372 10.6151
R806 B.n373 B.n76 10.6151
R807 B.n377 B.n76 10.6151
R808 B.n378 B.n377 10.6151
R809 B.n379 B.n378 10.6151
R810 B.n379 B.n74 10.6151
R811 B.n383 B.n74 10.6151
R812 B.n384 B.n383 10.6151
R813 B.n385 B.n384 10.6151
R814 B.n385 B.n72 10.6151
R815 B.n389 B.n72 10.6151
R816 B.n390 B.n389 10.6151
R817 B.n391 B.n390 10.6151
R818 B.n391 B.n70 10.6151
R819 B.n395 B.n70 10.6151
R820 B.n396 B.n395 10.6151
R821 B.n181 B.n180 10.6151
R822 B.n181 B.n144 10.6151
R823 B.n185 B.n144 10.6151
R824 B.n186 B.n185 10.6151
R825 B.n187 B.n186 10.6151
R826 B.n187 B.n142 10.6151
R827 B.n191 B.n142 10.6151
R828 B.n192 B.n191 10.6151
R829 B.n193 B.n192 10.6151
R830 B.n193 B.n140 10.6151
R831 B.n197 B.n140 10.6151
R832 B.n198 B.n197 10.6151
R833 B.n199 B.n198 10.6151
R834 B.n199 B.n138 10.6151
R835 B.n203 B.n138 10.6151
R836 B.n204 B.n203 10.6151
R837 B.n205 B.n204 10.6151
R838 B.n205 B.n136 10.6151
R839 B.n209 B.n136 10.6151
R840 B.n210 B.n209 10.6151
R841 B.n211 B.n210 10.6151
R842 B.n211 B.n134 10.6151
R843 B.n215 B.n134 10.6151
R844 B.n216 B.n215 10.6151
R845 B.n217 B.n216 10.6151
R846 B.n217 B.n132 10.6151
R847 B.n221 B.n132 10.6151
R848 B.n222 B.n221 10.6151
R849 B.n223 B.n222 10.6151
R850 B.n223 B.n130 10.6151
R851 B.n227 B.n130 10.6151
R852 B.n228 B.n227 10.6151
R853 B.n229 B.n228 10.6151
R854 B.n229 B.n128 10.6151
R855 B.n233 B.n128 10.6151
R856 B.n234 B.n233 10.6151
R857 B.n235 B.n234 10.6151
R858 B.n235 B.n126 10.6151
R859 B.n239 B.n126 10.6151
R860 B.n240 B.n239 10.6151
R861 B.n241 B.n240 10.6151
R862 B.n241 B.n124 10.6151
R863 B.n245 B.n124 10.6151
R864 B.n246 B.n245 10.6151
R865 B.n247 B.n246 10.6151
R866 B.n247 B.n122 10.6151
R867 B.n251 B.n122 10.6151
R868 B.n252 B.n251 10.6151
R869 B.n254 B.n118 10.6151
R870 B.n258 B.n118 10.6151
R871 B.n259 B.n258 10.6151
R872 B.n260 B.n259 10.6151
R873 B.n260 B.n116 10.6151
R874 B.n264 B.n116 10.6151
R875 B.n265 B.n264 10.6151
R876 B.n266 B.n265 10.6151
R877 B.n270 B.n269 10.6151
R878 B.n271 B.n270 10.6151
R879 B.n271 B.n110 10.6151
R880 B.n275 B.n110 10.6151
R881 B.n276 B.n275 10.6151
R882 B.n277 B.n276 10.6151
R883 B.n277 B.n108 10.6151
R884 B.n281 B.n108 10.6151
R885 B.n282 B.n281 10.6151
R886 B.n283 B.n282 10.6151
R887 B.n283 B.n106 10.6151
R888 B.n287 B.n106 10.6151
R889 B.n288 B.n287 10.6151
R890 B.n289 B.n288 10.6151
R891 B.n289 B.n104 10.6151
R892 B.n293 B.n104 10.6151
R893 B.n294 B.n293 10.6151
R894 B.n295 B.n294 10.6151
R895 B.n295 B.n102 10.6151
R896 B.n299 B.n102 10.6151
R897 B.n300 B.n299 10.6151
R898 B.n301 B.n300 10.6151
R899 B.n301 B.n100 10.6151
R900 B.n305 B.n100 10.6151
R901 B.n306 B.n305 10.6151
R902 B.n307 B.n306 10.6151
R903 B.n307 B.n98 10.6151
R904 B.n311 B.n98 10.6151
R905 B.n312 B.n311 10.6151
R906 B.n313 B.n312 10.6151
R907 B.n313 B.n96 10.6151
R908 B.n317 B.n96 10.6151
R909 B.n318 B.n317 10.6151
R910 B.n319 B.n318 10.6151
R911 B.n319 B.n94 10.6151
R912 B.n323 B.n94 10.6151
R913 B.n324 B.n323 10.6151
R914 B.n325 B.n324 10.6151
R915 B.n325 B.n92 10.6151
R916 B.n329 B.n92 10.6151
R917 B.n330 B.n329 10.6151
R918 B.n331 B.n330 10.6151
R919 B.n331 B.n90 10.6151
R920 B.n335 B.n90 10.6151
R921 B.n336 B.n335 10.6151
R922 B.n337 B.n336 10.6151
R923 B.n337 B.n88 10.6151
R924 B.n341 B.n88 10.6151
R925 B.n179 B.n146 10.6151
R926 B.n175 B.n146 10.6151
R927 B.n175 B.n174 10.6151
R928 B.n174 B.n173 10.6151
R929 B.n173 B.n148 10.6151
R930 B.n169 B.n148 10.6151
R931 B.n169 B.n168 10.6151
R932 B.n168 B.n167 10.6151
R933 B.n167 B.n150 10.6151
R934 B.n163 B.n150 10.6151
R935 B.n163 B.n162 10.6151
R936 B.n162 B.n161 10.6151
R937 B.n161 B.n152 10.6151
R938 B.n157 B.n152 10.6151
R939 B.n157 B.n156 10.6151
R940 B.n156 B.n155 10.6151
R941 B.n155 B.n0 10.6151
R942 B.n583 B.n1 10.6151
R943 B.n583 B.n582 10.6151
R944 B.n582 B.n581 10.6151
R945 B.n581 B.n4 10.6151
R946 B.n577 B.n4 10.6151
R947 B.n577 B.n576 10.6151
R948 B.n576 B.n575 10.6151
R949 B.n575 B.n6 10.6151
R950 B.n571 B.n6 10.6151
R951 B.n571 B.n570 10.6151
R952 B.n570 B.n569 10.6151
R953 B.n569 B.n8 10.6151
R954 B.n565 B.n8 10.6151
R955 B.n565 B.n564 10.6151
R956 B.n564 B.n563 10.6151
R957 B.n563 B.n10 10.6151
R958 B.n559 B.n10 10.6151
R959 B.n485 B.n484 6.5566
R960 B.n472 B.n44 6.5566
R961 B.n254 B.n253 6.5566
R962 B.n266 B.n114 6.5566
R963 B.n486 B.n485 4.05904
R964 B.n469 B.n44 4.05904
R965 B.n253 B.n252 4.05904
R966 B.n269 B.n114 4.05904
R967 B.n587 B.n0 2.81026
R968 B.n587 B.n1 2.81026
C0 VP B 1.08974f
C1 VDD2 B 1.70232f
C2 VN VDD1 0.147951f
C3 VTAIL B 3.00105f
C4 VN VP 5.35764f
C5 VN VDD2 4.4011f
C6 VDD1 w_n1650_n3854# 1.94268f
C7 VN VTAIL 3.92944f
C8 VP w_n1650_n3854# 2.87789f
C9 VN B 0.75373f
C10 VDD2 w_n1650_n3854# 1.96122f
C11 VTAIL w_n1650_n3854# 3.3478f
C12 B w_n1650_n3854# 7.48752f
C13 VP VDD1 4.53036f
C14 VDD2 VDD1 0.6478f
C15 VN w_n1650_n3854# 2.67037f
C16 VTAIL VDD1 13.0526f
C17 VP VDD2 0.282913f
C18 VDD1 B 1.67757f
C19 VP VTAIL 3.94423f
C20 VTAIL VDD2 13.0832f
C21 VDD2 VSUBS 1.386238f
C22 VDD1 VSUBS 1.665395f
C23 VTAIL VSUBS 0.751105f
C24 VN VSUBS 4.63183f
C25 VP VSUBS 1.421427f
C26 B VSUBS 2.781424f
C27 w_n1650_n3854# VSUBS 78.0318f
C28 B.n0 VSUBS 0.004598f
C29 B.n1 VSUBS 0.004598f
C30 B.n2 VSUBS 0.007272f
C31 B.n3 VSUBS 0.007272f
C32 B.n4 VSUBS 0.007272f
C33 B.n5 VSUBS 0.007272f
C34 B.n6 VSUBS 0.007272f
C35 B.n7 VSUBS 0.007272f
C36 B.n8 VSUBS 0.007272f
C37 B.n9 VSUBS 0.007272f
C38 B.n10 VSUBS 0.007272f
C39 B.n11 VSUBS 0.017968f
C40 B.n12 VSUBS 0.007272f
C41 B.n13 VSUBS 0.007272f
C42 B.n14 VSUBS 0.007272f
C43 B.n15 VSUBS 0.007272f
C44 B.n16 VSUBS 0.007272f
C45 B.n17 VSUBS 0.007272f
C46 B.n18 VSUBS 0.007272f
C47 B.n19 VSUBS 0.007272f
C48 B.n20 VSUBS 0.007272f
C49 B.n21 VSUBS 0.007272f
C50 B.n22 VSUBS 0.007272f
C51 B.n23 VSUBS 0.007272f
C52 B.n24 VSUBS 0.007272f
C53 B.n25 VSUBS 0.007272f
C54 B.n26 VSUBS 0.007272f
C55 B.n27 VSUBS 0.007272f
C56 B.n28 VSUBS 0.007272f
C57 B.n29 VSUBS 0.007272f
C58 B.n30 VSUBS 0.007272f
C59 B.n31 VSUBS 0.007272f
C60 B.n32 VSUBS 0.007272f
C61 B.n33 VSUBS 0.007272f
C62 B.n34 VSUBS 0.007272f
C63 B.n35 VSUBS 0.007272f
C64 B.t2 VSUBS 0.497356f
C65 B.t1 VSUBS 0.504605f
C66 B.t0 VSUBS 0.312357f
C67 B.n36 VSUBS 0.140226f
C68 B.n37 VSUBS 0.065787f
C69 B.n38 VSUBS 0.007272f
C70 B.n39 VSUBS 0.007272f
C71 B.n40 VSUBS 0.007272f
C72 B.n41 VSUBS 0.007272f
C73 B.t8 VSUBS 0.497343f
C74 B.t7 VSUBS 0.504593f
C75 B.t6 VSUBS 0.312357f
C76 B.n42 VSUBS 0.140238f
C77 B.n43 VSUBS 0.0658f
C78 B.n44 VSUBS 0.016848f
C79 B.n45 VSUBS 0.007272f
C80 B.n46 VSUBS 0.007272f
C81 B.n47 VSUBS 0.007272f
C82 B.n48 VSUBS 0.007272f
C83 B.n49 VSUBS 0.007272f
C84 B.n50 VSUBS 0.007272f
C85 B.n51 VSUBS 0.007272f
C86 B.n52 VSUBS 0.007272f
C87 B.n53 VSUBS 0.007272f
C88 B.n54 VSUBS 0.007272f
C89 B.n55 VSUBS 0.007272f
C90 B.n56 VSUBS 0.007272f
C91 B.n57 VSUBS 0.007272f
C92 B.n58 VSUBS 0.007272f
C93 B.n59 VSUBS 0.007272f
C94 B.n60 VSUBS 0.007272f
C95 B.n61 VSUBS 0.007272f
C96 B.n62 VSUBS 0.007272f
C97 B.n63 VSUBS 0.007272f
C98 B.n64 VSUBS 0.007272f
C99 B.n65 VSUBS 0.007272f
C100 B.n66 VSUBS 0.007272f
C101 B.n67 VSUBS 0.007272f
C102 B.n68 VSUBS 0.007272f
C103 B.n69 VSUBS 0.017107f
C104 B.n70 VSUBS 0.007272f
C105 B.n71 VSUBS 0.007272f
C106 B.n72 VSUBS 0.007272f
C107 B.n73 VSUBS 0.007272f
C108 B.n74 VSUBS 0.007272f
C109 B.n75 VSUBS 0.007272f
C110 B.n76 VSUBS 0.007272f
C111 B.n77 VSUBS 0.007272f
C112 B.n78 VSUBS 0.007272f
C113 B.n79 VSUBS 0.007272f
C114 B.n80 VSUBS 0.007272f
C115 B.n81 VSUBS 0.007272f
C116 B.n82 VSUBS 0.007272f
C117 B.n83 VSUBS 0.007272f
C118 B.n84 VSUBS 0.007272f
C119 B.n85 VSUBS 0.007272f
C120 B.n86 VSUBS 0.007272f
C121 B.n87 VSUBS 0.017107f
C122 B.n88 VSUBS 0.007272f
C123 B.n89 VSUBS 0.007272f
C124 B.n90 VSUBS 0.007272f
C125 B.n91 VSUBS 0.007272f
C126 B.n92 VSUBS 0.007272f
C127 B.n93 VSUBS 0.007272f
C128 B.n94 VSUBS 0.007272f
C129 B.n95 VSUBS 0.007272f
C130 B.n96 VSUBS 0.007272f
C131 B.n97 VSUBS 0.007272f
C132 B.n98 VSUBS 0.007272f
C133 B.n99 VSUBS 0.007272f
C134 B.n100 VSUBS 0.007272f
C135 B.n101 VSUBS 0.007272f
C136 B.n102 VSUBS 0.007272f
C137 B.n103 VSUBS 0.007272f
C138 B.n104 VSUBS 0.007272f
C139 B.n105 VSUBS 0.007272f
C140 B.n106 VSUBS 0.007272f
C141 B.n107 VSUBS 0.007272f
C142 B.n108 VSUBS 0.007272f
C143 B.n109 VSUBS 0.007272f
C144 B.n110 VSUBS 0.007272f
C145 B.n111 VSUBS 0.007272f
C146 B.t4 VSUBS 0.497343f
C147 B.t5 VSUBS 0.504593f
C148 B.t3 VSUBS 0.312357f
C149 B.n112 VSUBS 0.140238f
C150 B.n113 VSUBS 0.0658f
C151 B.n114 VSUBS 0.016848f
C152 B.n115 VSUBS 0.007272f
C153 B.n116 VSUBS 0.007272f
C154 B.n117 VSUBS 0.007272f
C155 B.n118 VSUBS 0.007272f
C156 B.n119 VSUBS 0.007272f
C157 B.t10 VSUBS 0.497356f
C158 B.t11 VSUBS 0.504605f
C159 B.t9 VSUBS 0.312357f
C160 B.n120 VSUBS 0.140226f
C161 B.n121 VSUBS 0.065787f
C162 B.n122 VSUBS 0.007272f
C163 B.n123 VSUBS 0.007272f
C164 B.n124 VSUBS 0.007272f
C165 B.n125 VSUBS 0.007272f
C166 B.n126 VSUBS 0.007272f
C167 B.n127 VSUBS 0.007272f
C168 B.n128 VSUBS 0.007272f
C169 B.n129 VSUBS 0.007272f
C170 B.n130 VSUBS 0.007272f
C171 B.n131 VSUBS 0.007272f
C172 B.n132 VSUBS 0.007272f
C173 B.n133 VSUBS 0.007272f
C174 B.n134 VSUBS 0.007272f
C175 B.n135 VSUBS 0.007272f
C176 B.n136 VSUBS 0.007272f
C177 B.n137 VSUBS 0.007272f
C178 B.n138 VSUBS 0.007272f
C179 B.n139 VSUBS 0.007272f
C180 B.n140 VSUBS 0.007272f
C181 B.n141 VSUBS 0.007272f
C182 B.n142 VSUBS 0.007272f
C183 B.n143 VSUBS 0.007272f
C184 B.n144 VSUBS 0.007272f
C185 B.n145 VSUBS 0.017968f
C186 B.n146 VSUBS 0.007272f
C187 B.n147 VSUBS 0.007272f
C188 B.n148 VSUBS 0.007272f
C189 B.n149 VSUBS 0.007272f
C190 B.n150 VSUBS 0.007272f
C191 B.n151 VSUBS 0.007272f
C192 B.n152 VSUBS 0.007272f
C193 B.n153 VSUBS 0.007272f
C194 B.n154 VSUBS 0.007272f
C195 B.n155 VSUBS 0.007272f
C196 B.n156 VSUBS 0.007272f
C197 B.n157 VSUBS 0.007272f
C198 B.n158 VSUBS 0.007272f
C199 B.n159 VSUBS 0.007272f
C200 B.n160 VSUBS 0.007272f
C201 B.n161 VSUBS 0.007272f
C202 B.n162 VSUBS 0.007272f
C203 B.n163 VSUBS 0.007272f
C204 B.n164 VSUBS 0.007272f
C205 B.n165 VSUBS 0.007272f
C206 B.n166 VSUBS 0.007272f
C207 B.n167 VSUBS 0.007272f
C208 B.n168 VSUBS 0.007272f
C209 B.n169 VSUBS 0.007272f
C210 B.n170 VSUBS 0.007272f
C211 B.n171 VSUBS 0.007272f
C212 B.n172 VSUBS 0.007272f
C213 B.n173 VSUBS 0.007272f
C214 B.n174 VSUBS 0.007272f
C215 B.n175 VSUBS 0.007272f
C216 B.n176 VSUBS 0.007272f
C217 B.n177 VSUBS 0.007272f
C218 B.n178 VSUBS 0.017107f
C219 B.n179 VSUBS 0.017107f
C220 B.n180 VSUBS 0.017968f
C221 B.n181 VSUBS 0.007272f
C222 B.n182 VSUBS 0.007272f
C223 B.n183 VSUBS 0.007272f
C224 B.n184 VSUBS 0.007272f
C225 B.n185 VSUBS 0.007272f
C226 B.n186 VSUBS 0.007272f
C227 B.n187 VSUBS 0.007272f
C228 B.n188 VSUBS 0.007272f
C229 B.n189 VSUBS 0.007272f
C230 B.n190 VSUBS 0.007272f
C231 B.n191 VSUBS 0.007272f
C232 B.n192 VSUBS 0.007272f
C233 B.n193 VSUBS 0.007272f
C234 B.n194 VSUBS 0.007272f
C235 B.n195 VSUBS 0.007272f
C236 B.n196 VSUBS 0.007272f
C237 B.n197 VSUBS 0.007272f
C238 B.n198 VSUBS 0.007272f
C239 B.n199 VSUBS 0.007272f
C240 B.n200 VSUBS 0.007272f
C241 B.n201 VSUBS 0.007272f
C242 B.n202 VSUBS 0.007272f
C243 B.n203 VSUBS 0.007272f
C244 B.n204 VSUBS 0.007272f
C245 B.n205 VSUBS 0.007272f
C246 B.n206 VSUBS 0.007272f
C247 B.n207 VSUBS 0.007272f
C248 B.n208 VSUBS 0.007272f
C249 B.n209 VSUBS 0.007272f
C250 B.n210 VSUBS 0.007272f
C251 B.n211 VSUBS 0.007272f
C252 B.n212 VSUBS 0.007272f
C253 B.n213 VSUBS 0.007272f
C254 B.n214 VSUBS 0.007272f
C255 B.n215 VSUBS 0.007272f
C256 B.n216 VSUBS 0.007272f
C257 B.n217 VSUBS 0.007272f
C258 B.n218 VSUBS 0.007272f
C259 B.n219 VSUBS 0.007272f
C260 B.n220 VSUBS 0.007272f
C261 B.n221 VSUBS 0.007272f
C262 B.n222 VSUBS 0.007272f
C263 B.n223 VSUBS 0.007272f
C264 B.n224 VSUBS 0.007272f
C265 B.n225 VSUBS 0.007272f
C266 B.n226 VSUBS 0.007272f
C267 B.n227 VSUBS 0.007272f
C268 B.n228 VSUBS 0.007272f
C269 B.n229 VSUBS 0.007272f
C270 B.n230 VSUBS 0.007272f
C271 B.n231 VSUBS 0.007272f
C272 B.n232 VSUBS 0.007272f
C273 B.n233 VSUBS 0.007272f
C274 B.n234 VSUBS 0.007272f
C275 B.n235 VSUBS 0.007272f
C276 B.n236 VSUBS 0.007272f
C277 B.n237 VSUBS 0.007272f
C278 B.n238 VSUBS 0.007272f
C279 B.n239 VSUBS 0.007272f
C280 B.n240 VSUBS 0.007272f
C281 B.n241 VSUBS 0.007272f
C282 B.n242 VSUBS 0.007272f
C283 B.n243 VSUBS 0.007272f
C284 B.n244 VSUBS 0.007272f
C285 B.n245 VSUBS 0.007272f
C286 B.n246 VSUBS 0.007272f
C287 B.n247 VSUBS 0.007272f
C288 B.n248 VSUBS 0.007272f
C289 B.n249 VSUBS 0.007272f
C290 B.n250 VSUBS 0.007272f
C291 B.n251 VSUBS 0.007272f
C292 B.n252 VSUBS 0.005026f
C293 B.n253 VSUBS 0.016848f
C294 B.n254 VSUBS 0.005882f
C295 B.n255 VSUBS 0.007272f
C296 B.n256 VSUBS 0.007272f
C297 B.n257 VSUBS 0.007272f
C298 B.n258 VSUBS 0.007272f
C299 B.n259 VSUBS 0.007272f
C300 B.n260 VSUBS 0.007272f
C301 B.n261 VSUBS 0.007272f
C302 B.n262 VSUBS 0.007272f
C303 B.n263 VSUBS 0.007272f
C304 B.n264 VSUBS 0.007272f
C305 B.n265 VSUBS 0.007272f
C306 B.n266 VSUBS 0.005882f
C307 B.n267 VSUBS 0.007272f
C308 B.n268 VSUBS 0.007272f
C309 B.n269 VSUBS 0.005026f
C310 B.n270 VSUBS 0.007272f
C311 B.n271 VSUBS 0.007272f
C312 B.n272 VSUBS 0.007272f
C313 B.n273 VSUBS 0.007272f
C314 B.n274 VSUBS 0.007272f
C315 B.n275 VSUBS 0.007272f
C316 B.n276 VSUBS 0.007272f
C317 B.n277 VSUBS 0.007272f
C318 B.n278 VSUBS 0.007272f
C319 B.n279 VSUBS 0.007272f
C320 B.n280 VSUBS 0.007272f
C321 B.n281 VSUBS 0.007272f
C322 B.n282 VSUBS 0.007272f
C323 B.n283 VSUBS 0.007272f
C324 B.n284 VSUBS 0.007272f
C325 B.n285 VSUBS 0.007272f
C326 B.n286 VSUBS 0.007272f
C327 B.n287 VSUBS 0.007272f
C328 B.n288 VSUBS 0.007272f
C329 B.n289 VSUBS 0.007272f
C330 B.n290 VSUBS 0.007272f
C331 B.n291 VSUBS 0.007272f
C332 B.n292 VSUBS 0.007272f
C333 B.n293 VSUBS 0.007272f
C334 B.n294 VSUBS 0.007272f
C335 B.n295 VSUBS 0.007272f
C336 B.n296 VSUBS 0.007272f
C337 B.n297 VSUBS 0.007272f
C338 B.n298 VSUBS 0.007272f
C339 B.n299 VSUBS 0.007272f
C340 B.n300 VSUBS 0.007272f
C341 B.n301 VSUBS 0.007272f
C342 B.n302 VSUBS 0.007272f
C343 B.n303 VSUBS 0.007272f
C344 B.n304 VSUBS 0.007272f
C345 B.n305 VSUBS 0.007272f
C346 B.n306 VSUBS 0.007272f
C347 B.n307 VSUBS 0.007272f
C348 B.n308 VSUBS 0.007272f
C349 B.n309 VSUBS 0.007272f
C350 B.n310 VSUBS 0.007272f
C351 B.n311 VSUBS 0.007272f
C352 B.n312 VSUBS 0.007272f
C353 B.n313 VSUBS 0.007272f
C354 B.n314 VSUBS 0.007272f
C355 B.n315 VSUBS 0.007272f
C356 B.n316 VSUBS 0.007272f
C357 B.n317 VSUBS 0.007272f
C358 B.n318 VSUBS 0.007272f
C359 B.n319 VSUBS 0.007272f
C360 B.n320 VSUBS 0.007272f
C361 B.n321 VSUBS 0.007272f
C362 B.n322 VSUBS 0.007272f
C363 B.n323 VSUBS 0.007272f
C364 B.n324 VSUBS 0.007272f
C365 B.n325 VSUBS 0.007272f
C366 B.n326 VSUBS 0.007272f
C367 B.n327 VSUBS 0.007272f
C368 B.n328 VSUBS 0.007272f
C369 B.n329 VSUBS 0.007272f
C370 B.n330 VSUBS 0.007272f
C371 B.n331 VSUBS 0.007272f
C372 B.n332 VSUBS 0.007272f
C373 B.n333 VSUBS 0.007272f
C374 B.n334 VSUBS 0.007272f
C375 B.n335 VSUBS 0.007272f
C376 B.n336 VSUBS 0.007272f
C377 B.n337 VSUBS 0.007272f
C378 B.n338 VSUBS 0.007272f
C379 B.n339 VSUBS 0.007272f
C380 B.n340 VSUBS 0.017968f
C381 B.n341 VSUBS 0.017968f
C382 B.n342 VSUBS 0.017107f
C383 B.n343 VSUBS 0.007272f
C384 B.n344 VSUBS 0.007272f
C385 B.n345 VSUBS 0.007272f
C386 B.n346 VSUBS 0.007272f
C387 B.n347 VSUBS 0.007272f
C388 B.n348 VSUBS 0.007272f
C389 B.n349 VSUBS 0.007272f
C390 B.n350 VSUBS 0.007272f
C391 B.n351 VSUBS 0.007272f
C392 B.n352 VSUBS 0.007272f
C393 B.n353 VSUBS 0.007272f
C394 B.n354 VSUBS 0.007272f
C395 B.n355 VSUBS 0.007272f
C396 B.n356 VSUBS 0.007272f
C397 B.n357 VSUBS 0.007272f
C398 B.n358 VSUBS 0.007272f
C399 B.n359 VSUBS 0.007272f
C400 B.n360 VSUBS 0.007272f
C401 B.n361 VSUBS 0.007272f
C402 B.n362 VSUBS 0.007272f
C403 B.n363 VSUBS 0.007272f
C404 B.n364 VSUBS 0.007272f
C405 B.n365 VSUBS 0.007272f
C406 B.n366 VSUBS 0.007272f
C407 B.n367 VSUBS 0.007272f
C408 B.n368 VSUBS 0.007272f
C409 B.n369 VSUBS 0.007272f
C410 B.n370 VSUBS 0.007272f
C411 B.n371 VSUBS 0.007272f
C412 B.n372 VSUBS 0.007272f
C413 B.n373 VSUBS 0.007272f
C414 B.n374 VSUBS 0.007272f
C415 B.n375 VSUBS 0.007272f
C416 B.n376 VSUBS 0.007272f
C417 B.n377 VSUBS 0.007272f
C418 B.n378 VSUBS 0.007272f
C419 B.n379 VSUBS 0.007272f
C420 B.n380 VSUBS 0.007272f
C421 B.n381 VSUBS 0.007272f
C422 B.n382 VSUBS 0.007272f
C423 B.n383 VSUBS 0.007272f
C424 B.n384 VSUBS 0.007272f
C425 B.n385 VSUBS 0.007272f
C426 B.n386 VSUBS 0.007272f
C427 B.n387 VSUBS 0.007272f
C428 B.n388 VSUBS 0.007272f
C429 B.n389 VSUBS 0.007272f
C430 B.n390 VSUBS 0.007272f
C431 B.n391 VSUBS 0.007272f
C432 B.n392 VSUBS 0.007272f
C433 B.n393 VSUBS 0.007272f
C434 B.n394 VSUBS 0.007272f
C435 B.n395 VSUBS 0.007272f
C436 B.n396 VSUBS 0.017928f
C437 B.n397 VSUBS 0.017147f
C438 B.n398 VSUBS 0.017968f
C439 B.n399 VSUBS 0.007272f
C440 B.n400 VSUBS 0.007272f
C441 B.n401 VSUBS 0.007272f
C442 B.n402 VSUBS 0.007272f
C443 B.n403 VSUBS 0.007272f
C444 B.n404 VSUBS 0.007272f
C445 B.n405 VSUBS 0.007272f
C446 B.n406 VSUBS 0.007272f
C447 B.n407 VSUBS 0.007272f
C448 B.n408 VSUBS 0.007272f
C449 B.n409 VSUBS 0.007272f
C450 B.n410 VSUBS 0.007272f
C451 B.n411 VSUBS 0.007272f
C452 B.n412 VSUBS 0.007272f
C453 B.n413 VSUBS 0.007272f
C454 B.n414 VSUBS 0.007272f
C455 B.n415 VSUBS 0.007272f
C456 B.n416 VSUBS 0.007272f
C457 B.n417 VSUBS 0.007272f
C458 B.n418 VSUBS 0.007272f
C459 B.n419 VSUBS 0.007272f
C460 B.n420 VSUBS 0.007272f
C461 B.n421 VSUBS 0.007272f
C462 B.n422 VSUBS 0.007272f
C463 B.n423 VSUBS 0.007272f
C464 B.n424 VSUBS 0.007272f
C465 B.n425 VSUBS 0.007272f
C466 B.n426 VSUBS 0.007272f
C467 B.n427 VSUBS 0.007272f
C468 B.n428 VSUBS 0.007272f
C469 B.n429 VSUBS 0.007272f
C470 B.n430 VSUBS 0.007272f
C471 B.n431 VSUBS 0.007272f
C472 B.n432 VSUBS 0.007272f
C473 B.n433 VSUBS 0.007272f
C474 B.n434 VSUBS 0.007272f
C475 B.n435 VSUBS 0.007272f
C476 B.n436 VSUBS 0.007272f
C477 B.n437 VSUBS 0.007272f
C478 B.n438 VSUBS 0.007272f
C479 B.n439 VSUBS 0.007272f
C480 B.n440 VSUBS 0.007272f
C481 B.n441 VSUBS 0.007272f
C482 B.n442 VSUBS 0.007272f
C483 B.n443 VSUBS 0.007272f
C484 B.n444 VSUBS 0.007272f
C485 B.n445 VSUBS 0.007272f
C486 B.n446 VSUBS 0.007272f
C487 B.n447 VSUBS 0.007272f
C488 B.n448 VSUBS 0.007272f
C489 B.n449 VSUBS 0.007272f
C490 B.n450 VSUBS 0.007272f
C491 B.n451 VSUBS 0.007272f
C492 B.n452 VSUBS 0.007272f
C493 B.n453 VSUBS 0.007272f
C494 B.n454 VSUBS 0.007272f
C495 B.n455 VSUBS 0.007272f
C496 B.n456 VSUBS 0.007272f
C497 B.n457 VSUBS 0.007272f
C498 B.n458 VSUBS 0.007272f
C499 B.n459 VSUBS 0.007272f
C500 B.n460 VSUBS 0.007272f
C501 B.n461 VSUBS 0.007272f
C502 B.n462 VSUBS 0.007272f
C503 B.n463 VSUBS 0.007272f
C504 B.n464 VSUBS 0.007272f
C505 B.n465 VSUBS 0.007272f
C506 B.n466 VSUBS 0.007272f
C507 B.n467 VSUBS 0.007272f
C508 B.n468 VSUBS 0.007272f
C509 B.n469 VSUBS 0.005026f
C510 B.n470 VSUBS 0.007272f
C511 B.n471 VSUBS 0.007272f
C512 B.n472 VSUBS 0.005882f
C513 B.n473 VSUBS 0.007272f
C514 B.n474 VSUBS 0.007272f
C515 B.n475 VSUBS 0.007272f
C516 B.n476 VSUBS 0.007272f
C517 B.n477 VSUBS 0.007272f
C518 B.n478 VSUBS 0.007272f
C519 B.n479 VSUBS 0.007272f
C520 B.n480 VSUBS 0.007272f
C521 B.n481 VSUBS 0.007272f
C522 B.n482 VSUBS 0.007272f
C523 B.n483 VSUBS 0.007272f
C524 B.n484 VSUBS 0.005882f
C525 B.n485 VSUBS 0.016848f
C526 B.n486 VSUBS 0.005026f
C527 B.n487 VSUBS 0.007272f
C528 B.n488 VSUBS 0.007272f
C529 B.n489 VSUBS 0.007272f
C530 B.n490 VSUBS 0.007272f
C531 B.n491 VSUBS 0.007272f
C532 B.n492 VSUBS 0.007272f
C533 B.n493 VSUBS 0.007272f
C534 B.n494 VSUBS 0.007272f
C535 B.n495 VSUBS 0.007272f
C536 B.n496 VSUBS 0.007272f
C537 B.n497 VSUBS 0.007272f
C538 B.n498 VSUBS 0.007272f
C539 B.n499 VSUBS 0.007272f
C540 B.n500 VSUBS 0.007272f
C541 B.n501 VSUBS 0.007272f
C542 B.n502 VSUBS 0.007272f
C543 B.n503 VSUBS 0.007272f
C544 B.n504 VSUBS 0.007272f
C545 B.n505 VSUBS 0.007272f
C546 B.n506 VSUBS 0.007272f
C547 B.n507 VSUBS 0.007272f
C548 B.n508 VSUBS 0.007272f
C549 B.n509 VSUBS 0.007272f
C550 B.n510 VSUBS 0.007272f
C551 B.n511 VSUBS 0.007272f
C552 B.n512 VSUBS 0.007272f
C553 B.n513 VSUBS 0.007272f
C554 B.n514 VSUBS 0.007272f
C555 B.n515 VSUBS 0.007272f
C556 B.n516 VSUBS 0.007272f
C557 B.n517 VSUBS 0.007272f
C558 B.n518 VSUBS 0.007272f
C559 B.n519 VSUBS 0.007272f
C560 B.n520 VSUBS 0.007272f
C561 B.n521 VSUBS 0.007272f
C562 B.n522 VSUBS 0.007272f
C563 B.n523 VSUBS 0.007272f
C564 B.n524 VSUBS 0.007272f
C565 B.n525 VSUBS 0.007272f
C566 B.n526 VSUBS 0.007272f
C567 B.n527 VSUBS 0.007272f
C568 B.n528 VSUBS 0.007272f
C569 B.n529 VSUBS 0.007272f
C570 B.n530 VSUBS 0.007272f
C571 B.n531 VSUBS 0.007272f
C572 B.n532 VSUBS 0.007272f
C573 B.n533 VSUBS 0.007272f
C574 B.n534 VSUBS 0.007272f
C575 B.n535 VSUBS 0.007272f
C576 B.n536 VSUBS 0.007272f
C577 B.n537 VSUBS 0.007272f
C578 B.n538 VSUBS 0.007272f
C579 B.n539 VSUBS 0.007272f
C580 B.n540 VSUBS 0.007272f
C581 B.n541 VSUBS 0.007272f
C582 B.n542 VSUBS 0.007272f
C583 B.n543 VSUBS 0.007272f
C584 B.n544 VSUBS 0.007272f
C585 B.n545 VSUBS 0.007272f
C586 B.n546 VSUBS 0.007272f
C587 B.n547 VSUBS 0.007272f
C588 B.n548 VSUBS 0.007272f
C589 B.n549 VSUBS 0.007272f
C590 B.n550 VSUBS 0.007272f
C591 B.n551 VSUBS 0.007272f
C592 B.n552 VSUBS 0.007272f
C593 B.n553 VSUBS 0.007272f
C594 B.n554 VSUBS 0.007272f
C595 B.n555 VSUBS 0.007272f
C596 B.n556 VSUBS 0.007272f
C597 B.n557 VSUBS 0.007272f
C598 B.n558 VSUBS 0.017968f
C599 B.n559 VSUBS 0.017107f
C600 B.n560 VSUBS 0.017107f
C601 B.n561 VSUBS 0.007272f
C602 B.n562 VSUBS 0.007272f
C603 B.n563 VSUBS 0.007272f
C604 B.n564 VSUBS 0.007272f
C605 B.n565 VSUBS 0.007272f
C606 B.n566 VSUBS 0.007272f
C607 B.n567 VSUBS 0.007272f
C608 B.n568 VSUBS 0.007272f
C609 B.n569 VSUBS 0.007272f
C610 B.n570 VSUBS 0.007272f
C611 B.n571 VSUBS 0.007272f
C612 B.n572 VSUBS 0.007272f
C613 B.n573 VSUBS 0.007272f
C614 B.n574 VSUBS 0.007272f
C615 B.n575 VSUBS 0.007272f
C616 B.n576 VSUBS 0.007272f
C617 B.n577 VSUBS 0.007272f
C618 B.n578 VSUBS 0.007272f
C619 B.n579 VSUBS 0.007272f
C620 B.n580 VSUBS 0.007272f
C621 B.n581 VSUBS 0.007272f
C622 B.n582 VSUBS 0.007272f
C623 B.n583 VSUBS 0.007272f
C624 B.n584 VSUBS 0.007272f
C625 B.n585 VSUBS 0.007272f
C626 B.n586 VSUBS 0.007272f
C627 B.n587 VSUBS 0.016466f
C628 VDD1.t3 VSUBS 2.96728f
C629 VDD1.t1 VSUBS 2.96633f
C630 VDD1.t4 VSUBS 0.280985f
C631 VDD1.t5 VSUBS 0.280985f
C632 VDD1.n0 VSUBS 2.27883f
C633 VDD1.n1 VSUBS 2.722f
C634 VDD1.t0 VSUBS 0.280985f
C635 VDD1.t2 VSUBS 0.280985f
C636 VDD1.n2 VSUBS 2.27789f
C637 VDD1.n3 VSUBS 2.61201f
C638 VP.n0 VSUBS 0.082518f
C639 VP.t2 VSUBS 1.34074f
C640 VP.n1 VSUBS 0.501058f
C641 VP.t3 VSUBS 1.32274f
C642 VP.t5 VSUBS 1.32274f
C643 VP.n2 VSUBS 0.531875f
C644 VP.n3 VSUBS 0.517809f
C645 VP.n4 VSUBS 2.78672f
C646 VP.n5 VSUBS 2.66696f
C647 VP.t4 VSUBS 1.32274f
C648 VP.n6 VSUBS 0.517809f
C649 VP.t1 VSUBS 1.32274f
C650 VP.n7 VSUBS 0.531875f
C651 VP.t0 VSUBS 1.32274f
C652 VP.n8 VSUBS 0.517809f
C653 VP.n9 VSUBS 0.068763f
C654 VDD2.t5 VSUBS 2.96481f
C655 VDD2.t1 VSUBS 0.280841f
C656 VDD2.t0 VSUBS 0.280841f
C657 VDD2.n0 VSUBS 2.27766f
C658 VDD2.n1 VSUBS 2.64814f
C659 VDD2.t3 VSUBS 2.96102f
C660 VDD2.n2 VSUBS 2.65395f
C661 VDD2.t2 VSUBS 0.280841f
C662 VDD2.t4 VSUBS 0.280841f
C663 VDD2.n3 VSUBS 2.27762f
C664 VTAIL.t7 VSUBS 0.339994f
C665 VTAIL.t6 VSUBS 0.339994f
C666 VTAIL.n0 VSUBS 2.59638f
C667 VTAIL.n1 VSUBS 0.777586f
C668 VTAIL.t11 VSUBS 3.40315f
C669 VTAIL.n2 VSUBS 0.945284f
C670 VTAIL.t2 VSUBS 0.339994f
C671 VTAIL.t0 VSUBS 0.339994f
C672 VTAIL.n3 VSUBS 2.59638f
C673 VTAIL.n4 VSUBS 2.4854f
C674 VTAIL.t9 VSUBS 0.339994f
C675 VTAIL.t8 VSUBS 0.339994f
C676 VTAIL.n5 VSUBS 2.59638f
C677 VTAIL.n6 VSUBS 2.4854f
C678 VTAIL.t10 VSUBS 3.40317f
C679 VTAIL.n7 VSUBS 0.945257f
C680 VTAIL.t3 VSUBS 0.339994f
C681 VTAIL.t4 VSUBS 0.339994f
C682 VTAIL.n8 VSUBS 2.59638f
C683 VTAIL.n9 VSUBS 0.824789f
C684 VTAIL.t1 VSUBS 3.40315f
C685 VTAIL.n10 VSUBS 2.53549f
C686 VTAIL.t5 VSUBS 3.40315f
C687 VTAIL.n11 VSUBS 2.5123f
C688 VN.t0 VSUBS 1.30983f
C689 VN.n0 VSUBS 0.489503f
C690 VN.t4 VSUBS 1.29224f
C691 VN.n1 VSUBS 0.519609f
C692 VN.t5 VSUBS 1.29224f
C693 VN.n2 VSUBS 0.505868f
C694 VN.n3 VSUBS 0.235585f
C695 VN.t1 VSUBS 1.30983f
C696 VN.n4 VSUBS 0.489503f
C697 VN.t3 VSUBS 1.29224f
C698 VN.n5 VSUBS 0.519609f
C699 VN.t2 VSUBS 1.29224f
C700 VN.n6 VSUBS 0.505868f
C701 VN.n7 VSUBS 2.76219f
.ends

