**** sch_path: /home/chandru/MPW4_workdir/xschem_mpw4/LC_Cell
**.subckt LC_Cell Ibias outn outp ind_sub VDD GND
***.ipin Ibias
***.opin outn
***.opin outp
**XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
**XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=256 m=1
**XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
**.ends
**
**.subckt LC_Cell_pfet Ibias outn outp ind_sub VDD GND
**** Higher current mirrorring ratio 1:4, increased by 2, increasing Cap W by 4X
***.ipin Ibias
***.opin outn
***.opin outp
**XM1 outp outn GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=4.8 nf=10
**XM2 outn outp GND GND sky130_fd_pr__pfet_01v8 L=0.15 W=4.8 nf=10
**XL1 outp outn net1 ind_sub sky130_fd_pr__ind_05_220
**XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=256 m=1
**XM4 net1 Ibias VDD GND sky130_fd_pr__pfet_01v8 L=0.15 W=4.8 nf=20
**XM3 Ibias Ibias VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=5
**.ends 
**
**.subckt LC_Cell_1 Ibias outn outp ind_sub VDD GND 
**** Higher current mirrorring ratio 1:4, increased by 2
***.ipin Ibias
***.opin outn
***.opin outp
**XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
**XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=256 m=1
**XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.4 nf=5
**.ends
**
**.subckt LC_Cell_2 Ibias outn outp ind_sub VDD GND 
**** Higher current mirrorring ratio 1:4, increased by 2, increasing Cap W by 4X
***.ipin Ibias
***.opin outn
***.opin outp
**XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
**XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
**XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=2.4 nf=5
**.ends 

.subckt LC_Cell_3 Ibias outn outp ind_sub VDD GND
** Higher current mirrorring ratio 1:4, increased by 2, increasing Cap W by 4X
*.ipin Ibias
*.opin outn
*.opin outp
XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5 
XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=12
XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=12
XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC2 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC3 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC4 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
*XC5 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.3 W=2.4 nf=2
.ends

**.subckt LC_Cell_4 Ibias outn outp ind_sub VDD GND
**** Higher current mirrorring ratio 1:4, increased by 2, increasing Cap W by 4X
***.ipin Ibias
***.opin outn
***.opin outp
**XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
**XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
**XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.3 W=4.8 nf=10
**XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
**
**XMS1 outpi VDD outni GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=5
**XC1 outp outpi sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
**XC2 outp outpi sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
**XC3 outni outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
**XC4 outni outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
***XC5 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
**
**XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.3 W=4.8 nf=10
**XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.3 W=1.2 nf=2
**.ends
**
**
**.subckt LC_Cell_var Ibias outn outp ind_sub sw_on<1> sw_on<0> VDD GND 
**XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
**XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=4.8 nf=10
**XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1.2 nf=5
**
***Sw C1 
**XC1 outp net3 sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**XC2 net4 outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1 m=1
**XM6 net3 sw<0> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=1
***Sw C2
**XC3 outp net3 sky130_fd_pr__cap_mim_m3_1 W=32 L=5 MF=1 m=1
**XC4 net4 outn sky130_fd_pr__cap_mim_m3_1 W=32 L=5 MF=1 m=1
**XM7 net3 sw<1> net4 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1.2 nf=5
**.ends
**
**
**
.subckt LC_Cell_lvt Ibias outn outp ind_sub VDD GND
*.ipin Ibias
*.opin outn
*.opin outp
XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=5
XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=5
XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220

XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC2 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC3 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
XC4 outp outn sky130_fd_pr__cap_mim_m3_1 W=1 L=1 MF=1
*XC5 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.3 W=2.4 nf=2
.ends
**
**
**.subckt swcap_1m2c outp outn vsw Wc=1 Lc=1 Wsw=1.2 nsw=4 Lsw=0.15
**XC1 outp m1 sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
**XC2 m2 outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
**XM4 m1 vsw m2 m2 sky130_fd_pr__nfet_01v8 L=0.15 W=1.2 nf=4
**.ends


*.subckt LC_Cell_pfet Ibias outn outp ind_sub VDD GND
**.ipin Ibias
**.opin outn
**.opin outp
** Pfet LC oscillator
*XM1 outp outn GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
*XM2 outn outp GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
*XL1 outp outn net1 sky130_fd_pr__ind_05_220
*XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
*XM4 net1 Ibias VDD GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
*XM3 Ibias Ibias VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.4 nf=5
***XM1 outp outn net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
***XM2 outn outp net1 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
***XM3 net2 Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
***XL1 outp outn VDD ind_sub sky130_fd_pr__ind_05_220
***XC1 outp outn sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1
***XM4 net1 Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=4.8 nf=10
***XM5 Ibias Ibias GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2.4 nf=5
*.ends
