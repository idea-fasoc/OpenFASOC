* NGSPICE file created from diff_pair_sample_0461.ext - technology: sky130A

.subckt diff_pair_sample_0461 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=3.6582 ps=19.54 w=9.38 l=2.4
X1 B.t11 B.t9 B.t10 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=0 ps=0 w=9.38 l=2.4
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=3.6582 ps=19.54 w=9.38 l=2.4
X3 B.t8 B.t6 B.t7 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=0 ps=0 w=9.38 l=2.4
X4 VDD1.t0 VP.t1 VTAIL.t2 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=3.6582 ps=19.54 w=9.38 l=2.4
X5 B.t5 B.t3 B.t4 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=0 ps=0 w=9.38 l=2.4
X6 B.t2 B.t0 B.t1 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=0 ps=0 w=9.38 l=2.4
X7 VDD2.t0 VN.t1 VTAIL.t3 w_n2062_n2844# sky130_fd_pr__pfet_01v8 ad=3.6582 pd=19.54 as=3.6582 ps=19.54 w=9.38 l=2.4
R0 VP.n0 VP.t0 185.458
R1 VP.n0 VP.t1 143.317
R2 VP VP.n0 0.336784
R3 VTAIL.n194 VTAIL.n150 756.745
R4 VTAIL.n44 VTAIL.n0 756.745
R5 VTAIL.n144 VTAIL.n100 756.745
R6 VTAIL.n94 VTAIL.n50 756.745
R7 VTAIL.n167 VTAIL.n166 585
R8 VTAIL.n169 VTAIL.n168 585
R9 VTAIL.n162 VTAIL.n161 585
R10 VTAIL.n175 VTAIL.n174 585
R11 VTAIL.n177 VTAIL.n176 585
R12 VTAIL.n158 VTAIL.n157 585
R13 VTAIL.n184 VTAIL.n183 585
R14 VTAIL.n185 VTAIL.n156 585
R15 VTAIL.n187 VTAIL.n186 585
R16 VTAIL.n154 VTAIL.n153 585
R17 VTAIL.n193 VTAIL.n192 585
R18 VTAIL.n195 VTAIL.n194 585
R19 VTAIL.n17 VTAIL.n16 585
R20 VTAIL.n19 VTAIL.n18 585
R21 VTAIL.n12 VTAIL.n11 585
R22 VTAIL.n25 VTAIL.n24 585
R23 VTAIL.n27 VTAIL.n26 585
R24 VTAIL.n8 VTAIL.n7 585
R25 VTAIL.n34 VTAIL.n33 585
R26 VTAIL.n35 VTAIL.n6 585
R27 VTAIL.n37 VTAIL.n36 585
R28 VTAIL.n4 VTAIL.n3 585
R29 VTAIL.n43 VTAIL.n42 585
R30 VTAIL.n45 VTAIL.n44 585
R31 VTAIL.n145 VTAIL.n144 585
R32 VTAIL.n143 VTAIL.n142 585
R33 VTAIL.n104 VTAIL.n103 585
R34 VTAIL.n108 VTAIL.n106 585
R35 VTAIL.n137 VTAIL.n136 585
R36 VTAIL.n135 VTAIL.n134 585
R37 VTAIL.n110 VTAIL.n109 585
R38 VTAIL.n129 VTAIL.n128 585
R39 VTAIL.n127 VTAIL.n126 585
R40 VTAIL.n114 VTAIL.n113 585
R41 VTAIL.n121 VTAIL.n120 585
R42 VTAIL.n119 VTAIL.n118 585
R43 VTAIL.n95 VTAIL.n94 585
R44 VTAIL.n93 VTAIL.n92 585
R45 VTAIL.n54 VTAIL.n53 585
R46 VTAIL.n58 VTAIL.n56 585
R47 VTAIL.n87 VTAIL.n86 585
R48 VTAIL.n85 VTAIL.n84 585
R49 VTAIL.n60 VTAIL.n59 585
R50 VTAIL.n79 VTAIL.n78 585
R51 VTAIL.n77 VTAIL.n76 585
R52 VTAIL.n64 VTAIL.n63 585
R53 VTAIL.n71 VTAIL.n70 585
R54 VTAIL.n69 VTAIL.n68 585
R55 VTAIL.n165 VTAIL.t3 329.038
R56 VTAIL.n15 VTAIL.t2 329.038
R57 VTAIL.n117 VTAIL.t1 329.038
R58 VTAIL.n67 VTAIL.t0 329.038
R59 VTAIL.n168 VTAIL.n167 171.744
R60 VTAIL.n168 VTAIL.n161 171.744
R61 VTAIL.n175 VTAIL.n161 171.744
R62 VTAIL.n176 VTAIL.n175 171.744
R63 VTAIL.n176 VTAIL.n157 171.744
R64 VTAIL.n184 VTAIL.n157 171.744
R65 VTAIL.n185 VTAIL.n184 171.744
R66 VTAIL.n186 VTAIL.n185 171.744
R67 VTAIL.n186 VTAIL.n153 171.744
R68 VTAIL.n193 VTAIL.n153 171.744
R69 VTAIL.n194 VTAIL.n193 171.744
R70 VTAIL.n18 VTAIL.n17 171.744
R71 VTAIL.n18 VTAIL.n11 171.744
R72 VTAIL.n25 VTAIL.n11 171.744
R73 VTAIL.n26 VTAIL.n25 171.744
R74 VTAIL.n26 VTAIL.n7 171.744
R75 VTAIL.n34 VTAIL.n7 171.744
R76 VTAIL.n35 VTAIL.n34 171.744
R77 VTAIL.n36 VTAIL.n35 171.744
R78 VTAIL.n36 VTAIL.n3 171.744
R79 VTAIL.n43 VTAIL.n3 171.744
R80 VTAIL.n44 VTAIL.n43 171.744
R81 VTAIL.n144 VTAIL.n143 171.744
R82 VTAIL.n143 VTAIL.n103 171.744
R83 VTAIL.n108 VTAIL.n103 171.744
R84 VTAIL.n136 VTAIL.n108 171.744
R85 VTAIL.n136 VTAIL.n135 171.744
R86 VTAIL.n135 VTAIL.n109 171.744
R87 VTAIL.n128 VTAIL.n109 171.744
R88 VTAIL.n128 VTAIL.n127 171.744
R89 VTAIL.n127 VTAIL.n113 171.744
R90 VTAIL.n120 VTAIL.n113 171.744
R91 VTAIL.n120 VTAIL.n119 171.744
R92 VTAIL.n94 VTAIL.n93 171.744
R93 VTAIL.n93 VTAIL.n53 171.744
R94 VTAIL.n58 VTAIL.n53 171.744
R95 VTAIL.n86 VTAIL.n58 171.744
R96 VTAIL.n86 VTAIL.n85 171.744
R97 VTAIL.n85 VTAIL.n59 171.744
R98 VTAIL.n78 VTAIL.n59 171.744
R99 VTAIL.n78 VTAIL.n77 171.744
R100 VTAIL.n77 VTAIL.n63 171.744
R101 VTAIL.n70 VTAIL.n63 171.744
R102 VTAIL.n70 VTAIL.n69 171.744
R103 VTAIL.n167 VTAIL.t3 85.8723
R104 VTAIL.n17 VTAIL.t2 85.8723
R105 VTAIL.n119 VTAIL.t1 85.8723
R106 VTAIL.n69 VTAIL.t0 85.8723
R107 VTAIL.n199 VTAIL.n198 34.9005
R108 VTAIL.n49 VTAIL.n48 34.9005
R109 VTAIL.n149 VTAIL.n148 34.9005
R110 VTAIL.n99 VTAIL.n98 34.9005
R111 VTAIL.n99 VTAIL.n49 25.16
R112 VTAIL.n199 VTAIL.n149 22.8065
R113 VTAIL.n187 VTAIL.n154 13.1884
R114 VTAIL.n37 VTAIL.n4 13.1884
R115 VTAIL.n106 VTAIL.n104 13.1884
R116 VTAIL.n56 VTAIL.n54 13.1884
R117 VTAIL.n188 VTAIL.n156 12.8005
R118 VTAIL.n192 VTAIL.n191 12.8005
R119 VTAIL.n38 VTAIL.n6 12.8005
R120 VTAIL.n42 VTAIL.n41 12.8005
R121 VTAIL.n142 VTAIL.n141 12.8005
R122 VTAIL.n138 VTAIL.n137 12.8005
R123 VTAIL.n92 VTAIL.n91 12.8005
R124 VTAIL.n88 VTAIL.n87 12.8005
R125 VTAIL.n183 VTAIL.n182 12.0247
R126 VTAIL.n195 VTAIL.n152 12.0247
R127 VTAIL.n33 VTAIL.n32 12.0247
R128 VTAIL.n45 VTAIL.n2 12.0247
R129 VTAIL.n145 VTAIL.n102 12.0247
R130 VTAIL.n134 VTAIL.n107 12.0247
R131 VTAIL.n95 VTAIL.n52 12.0247
R132 VTAIL.n84 VTAIL.n57 12.0247
R133 VTAIL.n181 VTAIL.n158 11.249
R134 VTAIL.n196 VTAIL.n150 11.249
R135 VTAIL.n31 VTAIL.n8 11.249
R136 VTAIL.n46 VTAIL.n0 11.249
R137 VTAIL.n146 VTAIL.n100 11.249
R138 VTAIL.n133 VTAIL.n110 11.249
R139 VTAIL.n96 VTAIL.n50 11.249
R140 VTAIL.n83 VTAIL.n60 11.249
R141 VTAIL.n166 VTAIL.n165 10.7239
R142 VTAIL.n16 VTAIL.n15 10.7239
R143 VTAIL.n118 VTAIL.n117 10.7239
R144 VTAIL.n68 VTAIL.n67 10.7239
R145 VTAIL.n178 VTAIL.n177 10.4732
R146 VTAIL.n28 VTAIL.n27 10.4732
R147 VTAIL.n130 VTAIL.n129 10.4732
R148 VTAIL.n80 VTAIL.n79 10.4732
R149 VTAIL.n174 VTAIL.n160 9.69747
R150 VTAIL.n24 VTAIL.n10 9.69747
R151 VTAIL.n126 VTAIL.n112 9.69747
R152 VTAIL.n76 VTAIL.n62 9.69747
R153 VTAIL.n198 VTAIL.n197 9.45567
R154 VTAIL.n48 VTAIL.n47 9.45567
R155 VTAIL.n148 VTAIL.n147 9.45567
R156 VTAIL.n98 VTAIL.n97 9.45567
R157 VTAIL.n197 VTAIL.n196 9.3005
R158 VTAIL.n152 VTAIL.n151 9.3005
R159 VTAIL.n191 VTAIL.n190 9.3005
R160 VTAIL.n164 VTAIL.n163 9.3005
R161 VTAIL.n171 VTAIL.n170 9.3005
R162 VTAIL.n173 VTAIL.n172 9.3005
R163 VTAIL.n160 VTAIL.n159 9.3005
R164 VTAIL.n179 VTAIL.n178 9.3005
R165 VTAIL.n181 VTAIL.n180 9.3005
R166 VTAIL.n182 VTAIL.n155 9.3005
R167 VTAIL.n189 VTAIL.n188 9.3005
R168 VTAIL.n47 VTAIL.n46 9.3005
R169 VTAIL.n2 VTAIL.n1 9.3005
R170 VTAIL.n41 VTAIL.n40 9.3005
R171 VTAIL.n14 VTAIL.n13 9.3005
R172 VTAIL.n21 VTAIL.n20 9.3005
R173 VTAIL.n23 VTAIL.n22 9.3005
R174 VTAIL.n10 VTAIL.n9 9.3005
R175 VTAIL.n29 VTAIL.n28 9.3005
R176 VTAIL.n31 VTAIL.n30 9.3005
R177 VTAIL.n32 VTAIL.n5 9.3005
R178 VTAIL.n39 VTAIL.n38 9.3005
R179 VTAIL.n116 VTAIL.n115 9.3005
R180 VTAIL.n123 VTAIL.n122 9.3005
R181 VTAIL.n125 VTAIL.n124 9.3005
R182 VTAIL.n112 VTAIL.n111 9.3005
R183 VTAIL.n131 VTAIL.n130 9.3005
R184 VTAIL.n133 VTAIL.n132 9.3005
R185 VTAIL.n107 VTAIL.n105 9.3005
R186 VTAIL.n139 VTAIL.n138 9.3005
R187 VTAIL.n147 VTAIL.n146 9.3005
R188 VTAIL.n102 VTAIL.n101 9.3005
R189 VTAIL.n141 VTAIL.n140 9.3005
R190 VTAIL.n66 VTAIL.n65 9.3005
R191 VTAIL.n73 VTAIL.n72 9.3005
R192 VTAIL.n75 VTAIL.n74 9.3005
R193 VTAIL.n62 VTAIL.n61 9.3005
R194 VTAIL.n81 VTAIL.n80 9.3005
R195 VTAIL.n83 VTAIL.n82 9.3005
R196 VTAIL.n57 VTAIL.n55 9.3005
R197 VTAIL.n89 VTAIL.n88 9.3005
R198 VTAIL.n97 VTAIL.n96 9.3005
R199 VTAIL.n52 VTAIL.n51 9.3005
R200 VTAIL.n91 VTAIL.n90 9.3005
R201 VTAIL.n173 VTAIL.n162 8.92171
R202 VTAIL.n23 VTAIL.n12 8.92171
R203 VTAIL.n125 VTAIL.n114 8.92171
R204 VTAIL.n75 VTAIL.n64 8.92171
R205 VTAIL.n170 VTAIL.n169 8.14595
R206 VTAIL.n20 VTAIL.n19 8.14595
R207 VTAIL.n122 VTAIL.n121 8.14595
R208 VTAIL.n72 VTAIL.n71 8.14595
R209 VTAIL.n166 VTAIL.n164 7.3702
R210 VTAIL.n16 VTAIL.n14 7.3702
R211 VTAIL.n118 VTAIL.n116 7.3702
R212 VTAIL.n68 VTAIL.n66 7.3702
R213 VTAIL.n169 VTAIL.n164 5.81868
R214 VTAIL.n19 VTAIL.n14 5.81868
R215 VTAIL.n121 VTAIL.n116 5.81868
R216 VTAIL.n71 VTAIL.n66 5.81868
R217 VTAIL.n170 VTAIL.n162 5.04292
R218 VTAIL.n20 VTAIL.n12 5.04292
R219 VTAIL.n122 VTAIL.n114 5.04292
R220 VTAIL.n72 VTAIL.n64 5.04292
R221 VTAIL.n174 VTAIL.n173 4.26717
R222 VTAIL.n24 VTAIL.n23 4.26717
R223 VTAIL.n126 VTAIL.n125 4.26717
R224 VTAIL.n76 VTAIL.n75 4.26717
R225 VTAIL.n177 VTAIL.n160 3.49141
R226 VTAIL.n27 VTAIL.n10 3.49141
R227 VTAIL.n129 VTAIL.n112 3.49141
R228 VTAIL.n79 VTAIL.n62 3.49141
R229 VTAIL.n178 VTAIL.n158 2.71565
R230 VTAIL.n198 VTAIL.n150 2.71565
R231 VTAIL.n28 VTAIL.n8 2.71565
R232 VTAIL.n48 VTAIL.n0 2.71565
R233 VTAIL.n148 VTAIL.n100 2.71565
R234 VTAIL.n130 VTAIL.n110 2.71565
R235 VTAIL.n98 VTAIL.n50 2.71565
R236 VTAIL.n80 VTAIL.n60 2.71565
R237 VTAIL.n165 VTAIL.n163 2.41283
R238 VTAIL.n15 VTAIL.n13 2.41283
R239 VTAIL.n117 VTAIL.n115 2.41283
R240 VTAIL.n67 VTAIL.n65 2.41283
R241 VTAIL.n183 VTAIL.n181 1.93989
R242 VTAIL.n196 VTAIL.n195 1.93989
R243 VTAIL.n33 VTAIL.n31 1.93989
R244 VTAIL.n46 VTAIL.n45 1.93989
R245 VTAIL.n146 VTAIL.n145 1.93989
R246 VTAIL.n134 VTAIL.n133 1.93989
R247 VTAIL.n96 VTAIL.n95 1.93989
R248 VTAIL.n84 VTAIL.n83 1.93989
R249 VTAIL.n149 VTAIL.n99 1.64705
R250 VTAIL.n182 VTAIL.n156 1.16414
R251 VTAIL.n192 VTAIL.n152 1.16414
R252 VTAIL.n32 VTAIL.n6 1.16414
R253 VTAIL.n42 VTAIL.n2 1.16414
R254 VTAIL.n142 VTAIL.n102 1.16414
R255 VTAIL.n137 VTAIL.n107 1.16414
R256 VTAIL.n92 VTAIL.n52 1.16414
R257 VTAIL.n87 VTAIL.n57 1.16414
R258 VTAIL VTAIL.n49 1.11688
R259 VTAIL VTAIL.n199 0.530672
R260 VTAIL.n188 VTAIL.n187 0.388379
R261 VTAIL.n191 VTAIL.n154 0.388379
R262 VTAIL.n38 VTAIL.n37 0.388379
R263 VTAIL.n41 VTAIL.n4 0.388379
R264 VTAIL.n141 VTAIL.n104 0.388379
R265 VTAIL.n138 VTAIL.n106 0.388379
R266 VTAIL.n91 VTAIL.n54 0.388379
R267 VTAIL.n88 VTAIL.n56 0.388379
R268 VTAIL.n171 VTAIL.n163 0.155672
R269 VTAIL.n172 VTAIL.n171 0.155672
R270 VTAIL.n172 VTAIL.n159 0.155672
R271 VTAIL.n179 VTAIL.n159 0.155672
R272 VTAIL.n180 VTAIL.n179 0.155672
R273 VTAIL.n180 VTAIL.n155 0.155672
R274 VTAIL.n189 VTAIL.n155 0.155672
R275 VTAIL.n190 VTAIL.n189 0.155672
R276 VTAIL.n190 VTAIL.n151 0.155672
R277 VTAIL.n197 VTAIL.n151 0.155672
R278 VTAIL.n21 VTAIL.n13 0.155672
R279 VTAIL.n22 VTAIL.n21 0.155672
R280 VTAIL.n22 VTAIL.n9 0.155672
R281 VTAIL.n29 VTAIL.n9 0.155672
R282 VTAIL.n30 VTAIL.n29 0.155672
R283 VTAIL.n30 VTAIL.n5 0.155672
R284 VTAIL.n39 VTAIL.n5 0.155672
R285 VTAIL.n40 VTAIL.n39 0.155672
R286 VTAIL.n40 VTAIL.n1 0.155672
R287 VTAIL.n47 VTAIL.n1 0.155672
R288 VTAIL.n147 VTAIL.n101 0.155672
R289 VTAIL.n140 VTAIL.n101 0.155672
R290 VTAIL.n140 VTAIL.n139 0.155672
R291 VTAIL.n139 VTAIL.n105 0.155672
R292 VTAIL.n132 VTAIL.n105 0.155672
R293 VTAIL.n132 VTAIL.n131 0.155672
R294 VTAIL.n131 VTAIL.n111 0.155672
R295 VTAIL.n124 VTAIL.n111 0.155672
R296 VTAIL.n124 VTAIL.n123 0.155672
R297 VTAIL.n123 VTAIL.n115 0.155672
R298 VTAIL.n97 VTAIL.n51 0.155672
R299 VTAIL.n90 VTAIL.n51 0.155672
R300 VTAIL.n90 VTAIL.n89 0.155672
R301 VTAIL.n89 VTAIL.n55 0.155672
R302 VTAIL.n82 VTAIL.n55 0.155672
R303 VTAIL.n82 VTAIL.n81 0.155672
R304 VTAIL.n81 VTAIL.n61 0.155672
R305 VTAIL.n74 VTAIL.n61 0.155672
R306 VTAIL.n74 VTAIL.n73 0.155672
R307 VTAIL.n73 VTAIL.n65 0.155672
R308 VDD1.n44 VDD1.n0 756.745
R309 VDD1.n93 VDD1.n49 756.745
R310 VDD1.n45 VDD1.n44 585
R311 VDD1.n43 VDD1.n42 585
R312 VDD1.n4 VDD1.n3 585
R313 VDD1.n8 VDD1.n6 585
R314 VDD1.n37 VDD1.n36 585
R315 VDD1.n35 VDD1.n34 585
R316 VDD1.n10 VDD1.n9 585
R317 VDD1.n29 VDD1.n28 585
R318 VDD1.n27 VDD1.n26 585
R319 VDD1.n14 VDD1.n13 585
R320 VDD1.n21 VDD1.n20 585
R321 VDD1.n19 VDD1.n18 585
R322 VDD1.n66 VDD1.n65 585
R323 VDD1.n68 VDD1.n67 585
R324 VDD1.n61 VDD1.n60 585
R325 VDD1.n74 VDD1.n73 585
R326 VDD1.n76 VDD1.n75 585
R327 VDD1.n57 VDD1.n56 585
R328 VDD1.n83 VDD1.n82 585
R329 VDD1.n84 VDD1.n55 585
R330 VDD1.n86 VDD1.n85 585
R331 VDD1.n53 VDD1.n52 585
R332 VDD1.n92 VDD1.n91 585
R333 VDD1.n94 VDD1.n93 585
R334 VDD1.n17 VDD1.t1 329.038
R335 VDD1.n64 VDD1.t0 329.038
R336 VDD1.n44 VDD1.n43 171.744
R337 VDD1.n43 VDD1.n3 171.744
R338 VDD1.n8 VDD1.n3 171.744
R339 VDD1.n36 VDD1.n8 171.744
R340 VDD1.n36 VDD1.n35 171.744
R341 VDD1.n35 VDD1.n9 171.744
R342 VDD1.n28 VDD1.n9 171.744
R343 VDD1.n28 VDD1.n27 171.744
R344 VDD1.n27 VDD1.n13 171.744
R345 VDD1.n20 VDD1.n13 171.744
R346 VDD1.n20 VDD1.n19 171.744
R347 VDD1.n67 VDD1.n66 171.744
R348 VDD1.n67 VDD1.n60 171.744
R349 VDD1.n74 VDD1.n60 171.744
R350 VDD1.n75 VDD1.n74 171.744
R351 VDD1.n75 VDD1.n56 171.744
R352 VDD1.n83 VDD1.n56 171.744
R353 VDD1.n84 VDD1.n83 171.744
R354 VDD1.n85 VDD1.n84 171.744
R355 VDD1.n85 VDD1.n52 171.744
R356 VDD1.n92 VDD1.n52 171.744
R357 VDD1.n93 VDD1.n92 171.744
R358 VDD1 VDD1.n97 89.145
R359 VDD1.n19 VDD1.t1 85.8723
R360 VDD1.n66 VDD1.t0 85.8723
R361 VDD1 VDD1.n48 52.2258
R362 VDD1.n6 VDD1.n4 13.1884
R363 VDD1.n86 VDD1.n53 13.1884
R364 VDD1.n42 VDD1.n41 12.8005
R365 VDD1.n38 VDD1.n37 12.8005
R366 VDD1.n87 VDD1.n55 12.8005
R367 VDD1.n91 VDD1.n90 12.8005
R368 VDD1.n45 VDD1.n2 12.0247
R369 VDD1.n34 VDD1.n7 12.0247
R370 VDD1.n82 VDD1.n81 12.0247
R371 VDD1.n94 VDD1.n51 12.0247
R372 VDD1.n46 VDD1.n0 11.249
R373 VDD1.n33 VDD1.n10 11.249
R374 VDD1.n80 VDD1.n57 11.249
R375 VDD1.n95 VDD1.n49 11.249
R376 VDD1.n18 VDD1.n17 10.7239
R377 VDD1.n65 VDD1.n64 10.7239
R378 VDD1.n30 VDD1.n29 10.4732
R379 VDD1.n77 VDD1.n76 10.4732
R380 VDD1.n26 VDD1.n12 9.69747
R381 VDD1.n73 VDD1.n59 9.69747
R382 VDD1.n48 VDD1.n47 9.45567
R383 VDD1.n97 VDD1.n96 9.45567
R384 VDD1.n16 VDD1.n15 9.3005
R385 VDD1.n23 VDD1.n22 9.3005
R386 VDD1.n25 VDD1.n24 9.3005
R387 VDD1.n12 VDD1.n11 9.3005
R388 VDD1.n31 VDD1.n30 9.3005
R389 VDD1.n33 VDD1.n32 9.3005
R390 VDD1.n7 VDD1.n5 9.3005
R391 VDD1.n39 VDD1.n38 9.3005
R392 VDD1.n47 VDD1.n46 9.3005
R393 VDD1.n2 VDD1.n1 9.3005
R394 VDD1.n41 VDD1.n40 9.3005
R395 VDD1.n96 VDD1.n95 9.3005
R396 VDD1.n51 VDD1.n50 9.3005
R397 VDD1.n90 VDD1.n89 9.3005
R398 VDD1.n63 VDD1.n62 9.3005
R399 VDD1.n70 VDD1.n69 9.3005
R400 VDD1.n72 VDD1.n71 9.3005
R401 VDD1.n59 VDD1.n58 9.3005
R402 VDD1.n78 VDD1.n77 9.3005
R403 VDD1.n80 VDD1.n79 9.3005
R404 VDD1.n81 VDD1.n54 9.3005
R405 VDD1.n88 VDD1.n87 9.3005
R406 VDD1.n25 VDD1.n14 8.92171
R407 VDD1.n72 VDD1.n61 8.92171
R408 VDD1.n22 VDD1.n21 8.14595
R409 VDD1.n69 VDD1.n68 8.14595
R410 VDD1.n18 VDD1.n16 7.3702
R411 VDD1.n65 VDD1.n63 7.3702
R412 VDD1.n21 VDD1.n16 5.81868
R413 VDD1.n68 VDD1.n63 5.81868
R414 VDD1.n22 VDD1.n14 5.04292
R415 VDD1.n69 VDD1.n61 5.04292
R416 VDD1.n26 VDD1.n25 4.26717
R417 VDD1.n73 VDD1.n72 4.26717
R418 VDD1.n29 VDD1.n12 3.49141
R419 VDD1.n76 VDD1.n59 3.49141
R420 VDD1.n48 VDD1.n0 2.71565
R421 VDD1.n30 VDD1.n10 2.71565
R422 VDD1.n77 VDD1.n57 2.71565
R423 VDD1.n97 VDD1.n49 2.71565
R424 VDD1.n17 VDD1.n15 2.41283
R425 VDD1.n64 VDD1.n62 2.41283
R426 VDD1.n46 VDD1.n45 1.93989
R427 VDD1.n34 VDD1.n33 1.93989
R428 VDD1.n82 VDD1.n80 1.93989
R429 VDD1.n95 VDD1.n94 1.93989
R430 VDD1.n42 VDD1.n2 1.16414
R431 VDD1.n37 VDD1.n7 1.16414
R432 VDD1.n81 VDD1.n55 1.16414
R433 VDD1.n91 VDD1.n51 1.16414
R434 VDD1.n41 VDD1.n4 0.388379
R435 VDD1.n38 VDD1.n6 0.388379
R436 VDD1.n87 VDD1.n86 0.388379
R437 VDD1.n90 VDD1.n53 0.388379
R438 VDD1.n47 VDD1.n1 0.155672
R439 VDD1.n40 VDD1.n1 0.155672
R440 VDD1.n40 VDD1.n39 0.155672
R441 VDD1.n39 VDD1.n5 0.155672
R442 VDD1.n32 VDD1.n5 0.155672
R443 VDD1.n32 VDD1.n31 0.155672
R444 VDD1.n31 VDD1.n11 0.155672
R445 VDD1.n24 VDD1.n11 0.155672
R446 VDD1.n24 VDD1.n23 0.155672
R447 VDD1.n23 VDD1.n15 0.155672
R448 VDD1.n70 VDD1.n62 0.155672
R449 VDD1.n71 VDD1.n70 0.155672
R450 VDD1.n71 VDD1.n58 0.155672
R451 VDD1.n78 VDD1.n58 0.155672
R452 VDD1.n79 VDD1.n78 0.155672
R453 VDD1.n79 VDD1.n54 0.155672
R454 VDD1.n88 VDD1.n54 0.155672
R455 VDD1.n89 VDD1.n88 0.155672
R456 VDD1.n89 VDD1.n50 0.155672
R457 VDD1.n96 VDD1.n50 0.155672
R458 B.n361 B.n56 585
R459 B.n363 B.n362 585
R460 B.n364 B.n55 585
R461 B.n366 B.n365 585
R462 B.n367 B.n54 585
R463 B.n369 B.n368 585
R464 B.n370 B.n53 585
R465 B.n372 B.n371 585
R466 B.n373 B.n52 585
R467 B.n375 B.n374 585
R468 B.n376 B.n51 585
R469 B.n378 B.n377 585
R470 B.n379 B.n50 585
R471 B.n381 B.n380 585
R472 B.n382 B.n49 585
R473 B.n384 B.n383 585
R474 B.n385 B.n48 585
R475 B.n387 B.n386 585
R476 B.n388 B.n47 585
R477 B.n390 B.n389 585
R478 B.n391 B.n46 585
R479 B.n393 B.n392 585
R480 B.n394 B.n45 585
R481 B.n396 B.n395 585
R482 B.n397 B.n44 585
R483 B.n399 B.n398 585
R484 B.n400 B.n43 585
R485 B.n402 B.n401 585
R486 B.n403 B.n42 585
R487 B.n405 B.n404 585
R488 B.n406 B.n41 585
R489 B.n408 B.n407 585
R490 B.n409 B.n40 585
R491 B.n411 B.n410 585
R492 B.n413 B.n37 585
R493 B.n415 B.n414 585
R494 B.n416 B.n36 585
R495 B.n418 B.n417 585
R496 B.n419 B.n35 585
R497 B.n421 B.n420 585
R498 B.n422 B.n34 585
R499 B.n424 B.n423 585
R500 B.n425 B.n31 585
R501 B.n428 B.n427 585
R502 B.n429 B.n30 585
R503 B.n431 B.n430 585
R504 B.n432 B.n29 585
R505 B.n434 B.n433 585
R506 B.n435 B.n28 585
R507 B.n437 B.n436 585
R508 B.n438 B.n27 585
R509 B.n440 B.n439 585
R510 B.n441 B.n26 585
R511 B.n443 B.n442 585
R512 B.n444 B.n25 585
R513 B.n446 B.n445 585
R514 B.n447 B.n24 585
R515 B.n449 B.n448 585
R516 B.n450 B.n23 585
R517 B.n452 B.n451 585
R518 B.n453 B.n22 585
R519 B.n455 B.n454 585
R520 B.n456 B.n21 585
R521 B.n458 B.n457 585
R522 B.n459 B.n20 585
R523 B.n461 B.n460 585
R524 B.n462 B.n19 585
R525 B.n464 B.n463 585
R526 B.n465 B.n18 585
R527 B.n467 B.n466 585
R528 B.n468 B.n17 585
R529 B.n470 B.n469 585
R530 B.n471 B.n16 585
R531 B.n473 B.n472 585
R532 B.n474 B.n15 585
R533 B.n476 B.n475 585
R534 B.n477 B.n14 585
R535 B.n360 B.n359 585
R536 B.n358 B.n57 585
R537 B.n357 B.n356 585
R538 B.n355 B.n58 585
R539 B.n354 B.n353 585
R540 B.n352 B.n59 585
R541 B.n351 B.n350 585
R542 B.n349 B.n60 585
R543 B.n348 B.n347 585
R544 B.n346 B.n61 585
R545 B.n345 B.n344 585
R546 B.n343 B.n62 585
R547 B.n342 B.n341 585
R548 B.n340 B.n63 585
R549 B.n339 B.n338 585
R550 B.n337 B.n64 585
R551 B.n336 B.n335 585
R552 B.n334 B.n65 585
R553 B.n333 B.n332 585
R554 B.n331 B.n66 585
R555 B.n330 B.n329 585
R556 B.n328 B.n67 585
R557 B.n327 B.n326 585
R558 B.n325 B.n68 585
R559 B.n324 B.n323 585
R560 B.n322 B.n69 585
R561 B.n321 B.n320 585
R562 B.n319 B.n70 585
R563 B.n318 B.n317 585
R564 B.n316 B.n71 585
R565 B.n315 B.n314 585
R566 B.n313 B.n72 585
R567 B.n312 B.n311 585
R568 B.n310 B.n73 585
R569 B.n309 B.n308 585
R570 B.n307 B.n74 585
R571 B.n306 B.n305 585
R572 B.n304 B.n75 585
R573 B.n303 B.n302 585
R574 B.n301 B.n76 585
R575 B.n300 B.n299 585
R576 B.n298 B.n77 585
R577 B.n297 B.n296 585
R578 B.n295 B.n78 585
R579 B.n294 B.n293 585
R580 B.n292 B.n79 585
R581 B.n291 B.n290 585
R582 B.n289 B.n80 585
R583 B.n288 B.n287 585
R584 B.n171 B.n170 585
R585 B.n172 B.n123 585
R586 B.n174 B.n173 585
R587 B.n175 B.n122 585
R588 B.n177 B.n176 585
R589 B.n178 B.n121 585
R590 B.n180 B.n179 585
R591 B.n181 B.n120 585
R592 B.n183 B.n182 585
R593 B.n184 B.n119 585
R594 B.n186 B.n185 585
R595 B.n187 B.n118 585
R596 B.n189 B.n188 585
R597 B.n190 B.n117 585
R598 B.n192 B.n191 585
R599 B.n193 B.n116 585
R600 B.n195 B.n194 585
R601 B.n196 B.n115 585
R602 B.n198 B.n197 585
R603 B.n199 B.n114 585
R604 B.n201 B.n200 585
R605 B.n202 B.n113 585
R606 B.n204 B.n203 585
R607 B.n205 B.n112 585
R608 B.n207 B.n206 585
R609 B.n208 B.n111 585
R610 B.n210 B.n209 585
R611 B.n211 B.n110 585
R612 B.n213 B.n212 585
R613 B.n214 B.n109 585
R614 B.n216 B.n215 585
R615 B.n217 B.n108 585
R616 B.n219 B.n218 585
R617 B.n220 B.n105 585
R618 B.n223 B.n222 585
R619 B.n224 B.n104 585
R620 B.n226 B.n225 585
R621 B.n227 B.n103 585
R622 B.n229 B.n228 585
R623 B.n230 B.n102 585
R624 B.n232 B.n231 585
R625 B.n233 B.n101 585
R626 B.n235 B.n234 585
R627 B.n237 B.n236 585
R628 B.n238 B.n97 585
R629 B.n240 B.n239 585
R630 B.n241 B.n96 585
R631 B.n243 B.n242 585
R632 B.n244 B.n95 585
R633 B.n246 B.n245 585
R634 B.n247 B.n94 585
R635 B.n249 B.n248 585
R636 B.n250 B.n93 585
R637 B.n252 B.n251 585
R638 B.n253 B.n92 585
R639 B.n255 B.n254 585
R640 B.n256 B.n91 585
R641 B.n258 B.n257 585
R642 B.n259 B.n90 585
R643 B.n261 B.n260 585
R644 B.n262 B.n89 585
R645 B.n264 B.n263 585
R646 B.n265 B.n88 585
R647 B.n267 B.n266 585
R648 B.n268 B.n87 585
R649 B.n270 B.n269 585
R650 B.n271 B.n86 585
R651 B.n273 B.n272 585
R652 B.n274 B.n85 585
R653 B.n276 B.n275 585
R654 B.n277 B.n84 585
R655 B.n279 B.n278 585
R656 B.n280 B.n83 585
R657 B.n282 B.n281 585
R658 B.n283 B.n82 585
R659 B.n285 B.n284 585
R660 B.n286 B.n81 585
R661 B.n169 B.n124 585
R662 B.n168 B.n167 585
R663 B.n166 B.n125 585
R664 B.n165 B.n164 585
R665 B.n163 B.n126 585
R666 B.n162 B.n161 585
R667 B.n160 B.n127 585
R668 B.n159 B.n158 585
R669 B.n157 B.n128 585
R670 B.n156 B.n155 585
R671 B.n154 B.n129 585
R672 B.n153 B.n152 585
R673 B.n151 B.n130 585
R674 B.n150 B.n149 585
R675 B.n148 B.n131 585
R676 B.n147 B.n146 585
R677 B.n145 B.n132 585
R678 B.n144 B.n143 585
R679 B.n142 B.n133 585
R680 B.n141 B.n140 585
R681 B.n139 B.n134 585
R682 B.n138 B.n137 585
R683 B.n136 B.n135 585
R684 B.n2 B.n0 585
R685 B.n513 B.n1 585
R686 B.n512 B.n511 585
R687 B.n510 B.n3 585
R688 B.n509 B.n508 585
R689 B.n507 B.n4 585
R690 B.n506 B.n505 585
R691 B.n504 B.n5 585
R692 B.n503 B.n502 585
R693 B.n501 B.n6 585
R694 B.n500 B.n499 585
R695 B.n498 B.n7 585
R696 B.n497 B.n496 585
R697 B.n495 B.n8 585
R698 B.n494 B.n493 585
R699 B.n492 B.n9 585
R700 B.n491 B.n490 585
R701 B.n489 B.n10 585
R702 B.n488 B.n487 585
R703 B.n486 B.n11 585
R704 B.n485 B.n484 585
R705 B.n483 B.n12 585
R706 B.n482 B.n481 585
R707 B.n480 B.n13 585
R708 B.n479 B.n478 585
R709 B.n515 B.n514 585
R710 B.n170 B.n169 559.769
R711 B.n478 B.n477 559.769
R712 B.n288 B.n81 559.769
R713 B.n361 B.n360 559.769
R714 B.n98 B.t5 381.452
R715 B.n38 B.t7 381.452
R716 B.n106 B.t2 381.452
R717 B.n32 B.t10 381.452
R718 B.n99 B.t4 328.505
R719 B.n39 B.t8 328.505
R720 B.n107 B.t1 328.505
R721 B.n33 B.t11 328.505
R722 B.n98 B.t3 301.914
R723 B.n106 B.t0 301.914
R724 B.n32 B.t9 301.914
R725 B.n38 B.t6 301.914
R726 B.n169 B.n168 163.367
R727 B.n168 B.n125 163.367
R728 B.n164 B.n125 163.367
R729 B.n164 B.n163 163.367
R730 B.n163 B.n162 163.367
R731 B.n162 B.n127 163.367
R732 B.n158 B.n127 163.367
R733 B.n158 B.n157 163.367
R734 B.n157 B.n156 163.367
R735 B.n156 B.n129 163.367
R736 B.n152 B.n129 163.367
R737 B.n152 B.n151 163.367
R738 B.n151 B.n150 163.367
R739 B.n150 B.n131 163.367
R740 B.n146 B.n131 163.367
R741 B.n146 B.n145 163.367
R742 B.n145 B.n144 163.367
R743 B.n144 B.n133 163.367
R744 B.n140 B.n133 163.367
R745 B.n140 B.n139 163.367
R746 B.n139 B.n138 163.367
R747 B.n138 B.n135 163.367
R748 B.n135 B.n2 163.367
R749 B.n514 B.n2 163.367
R750 B.n514 B.n513 163.367
R751 B.n513 B.n512 163.367
R752 B.n512 B.n3 163.367
R753 B.n508 B.n3 163.367
R754 B.n508 B.n507 163.367
R755 B.n507 B.n506 163.367
R756 B.n506 B.n5 163.367
R757 B.n502 B.n5 163.367
R758 B.n502 B.n501 163.367
R759 B.n501 B.n500 163.367
R760 B.n500 B.n7 163.367
R761 B.n496 B.n7 163.367
R762 B.n496 B.n495 163.367
R763 B.n495 B.n494 163.367
R764 B.n494 B.n9 163.367
R765 B.n490 B.n9 163.367
R766 B.n490 B.n489 163.367
R767 B.n489 B.n488 163.367
R768 B.n488 B.n11 163.367
R769 B.n484 B.n11 163.367
R770 B.n484 B.n483 163.367
R771 B.n483 B.n482 163.367
R772 B.n482 B.n13 163.367
R773 B.n478 B.n13 163.367
R774 B.n170 B.n123 163.367
R775 B.n174 B.n123 163.367
R776 B.n175 B.n174 163.367
R777 B.n176 B.n175 163.367
R778 B.n176 B.n121 163.367
R779 B.n180 B.n121 163.367
R780 B.n181 B.n180 163.367
R781 B.n182 B.n181 163.367
R782 B.n182 B.n119 163.367
R783 B.n186 B.n119 163.367
R784 B.n187 B.n186 163.367
R785 B.n188 B.n187 163.367
R786 B.n188 B.n117 163.367
R787 B.n192 B.n117 163.367
R788 B.n193 B.n192 163.367
R789 B.n194 B.n193 163.367
R790 B.n194 B.n115 163.367
R791 B.n198 B.n115 163.367
R792 B.n199 B.n198 163.367
R793 B.n200 B.n199 163.367
R794 B.n200 B.n113 163.367
R795 B.n204 B.n113 163.367
R796 B.n205 B.n204 163.367
R797 B.n206 B.n205 163.367
R798 B.n206 B.n111 163.367
R799 B.n210 B.n111 163.367
R800 B.n211 B.n210 163.367
R801 B.n212 B.n211 163.367
R802 B.n212 B.n109 163.367
R803 B.n216 B.n109 163.367
R804 B.n217 B.n216 163.367
R805 B.n218 B.n217 163.367
R806 B.n218 B.n105 163.367
R807 B.n223 B.n105 163.367
R808 B.n224 B.n223 163.367
R809 B.n225 B.n224 163.367
R810 B.n225 B.n103 163.367
R811 B.n229 B.n103 163.367
R812 B.n230 B.n229 163.367
R813 B.n231 B.n230 163.367
R814 B.n231 B.n101 163.367
R815 B.n235 B.n101 163.367
R816 B.n236 B.n235 163.367
R817 B.n236 B.n97 163.367
R818 B.n240 B.n97 163.367
R819 B.n241 B.n240 163.367
R820 B.n242 B.n241 163.367
R821 B.n242 B.n95 163.367
R822 B.n246 B.n95 163.367
R823 B.n247 B.n246 163.367
R824 B.n248 B.n247 163.367
R825 B.n248 B.n93 163.367
R826 B.n252 B.n93 163.367
R827 B.n253 B.n252 163.367
R828 B.n254 B.n253 163.367
R829 B.n254 B.n91 163.367
R830 B.n258 B.n91 163.367
R831 B.n259 B.n258 163.367
R832 B.n260 B.n259 163.367
R833 B.n260 B.n89 163.367
R834 B.n264 B.n89 163.367
R835 B.n265 B.n264 163.367
R836 B.n266 B.n265 163.367
R837 B.n266 B.n87 163.367
R838 B.n270 B.n87 163.367
R839 B.n271 B.n270 163.367
R840 B.n272 B.n271 163.367
R841 B.n272 B.n85 163.367
R842 B.n276 B.n85 163.367
R843 B.n277 B.n276 163.367
R844 B.n278 B.n277 163.367
R845 B.n278 B.n83 163.367
R846 B.n282 B.n83 163.367
R847 B.n283 B.n282 163.367
R848 B.n284 B.n283 163.367
R849 B.n284 B.n81 163.367
R850 B.n289 B.n288 163.367
R851 B.n290 B.n289 163.367
R852 B.n290 B.n79 163.367
R853 B.n294 B.n79 163.367
R854 B.n295 B.n294 163.367
R855 B.n296 B.n295 163.367
R856 B.n296 B.n77 163.367
R857 B.n300 B.n77 163.367
R858 B.n301 B.n300 163.367
R859 B.n302 B.n301 163.367
R860 B.n302 B.n75 163.367
R861 B.n306 B.n75 163.367
R862 B.n307 B.n306 163.367
R863 B.n308 B.n307 163.367
R864 B.n308 B.n73 163.367
R865 B.n312 B.n73 163.367
R866 B.n313 B.n312 163.367
R867 B.n314 B.n313 163.367
R868 B.n314 B.n71 163.367
R869 B.n318 B.n71 163.367
R870 B.n319 B.n318 163.367
R871 B.n320 B.n319 163.367
R872 B.n320 B.n69 163.367
R873 B.n324 B.n69 163.367
R874 B.n325 B.n324 163.367
R875 B.n326 B.n325 163.367
R876 B.n326 B.n67 163.367
R877 B.n330 B.n67 163.367
R878 B.n331 B.n330 163.367
R879 B.n332 B.n331 163.367
R880 B.n332 B.n65 163.367
R881 B.n336 B.n65 163.367
R882 B.n337 B.n336 163.367
R883 B.n338 B.n337 163.367
R884 B.n338 B.n63 163.367
R885 B.n342 B.n63 163.367
R886 B.n343 B.n342 163.367
R887 B.n344 B.n343 163.367
R888 B.n344 B.n61 163.367
R889 B.n348 B.n61 163.367
R890 B.n349 B.n348 163.367
R891 B.n350 B.n349 163.367
R892 B.n350 B.n59 163.367
R893 B.n354 B.n59 163.367
R894 B.n355 B.n354 163.367
R895 B.n356 B.n355 163.367
R896 B.n356 B.n57 163.367
R897 B.n360 B.n57 163.367
R898 B.n477 B.n476 163.367
R899 B.n476 B.n15 163.367
R900 B.n472 B.n15 163.367
R901 B.n472 B.n471 163.367
R902 B.n471 B.n470 163.367
R903 B.n470 B.n17 163.367
R904 B.n466 B.n17 163.367
R905 B.n466 B.n465 163.367
R906 B.n465 B.n464 163.367
R907 B.n464 B.n19 163.367
R908 B.n460 B.n19 163.367
R909 B.n460 B.n459 163.367
R910 B.n459 B.n458 163.367
R911 B.n458 B.n21 163.367
R912 B.n454 B.n21 163.367
R913 B.n454 B.n453 163.367
R914 B.n453 B.n452 163.367
R915 B.n452 B.n23 163.367
R916 B.n448 B.n23 163.367
R917 B.n448 B.n447 163.367
R918 B.n447 B.n446 163.367
R919 B.n446 B.n25 163.367
R920 B.n442 B.n25 163.367
R921 B.n442 B.n441 163.367
R922 B.n441 B.n440 163.367
R923 B.n440 B.n27 163.367
R924 B.n436 B.n27 163.367
R925 B.n436 B.n435 163.367
R926 B.n435 B.n434 163.367
R927 B.n434 B.n29 163.367
R928 B.n430 B.n29 163.367
R929 B.n430 B.n429 163.367
R930 B.n429 B.n428 163.367
R931 B.n428 B.n31 163.367
R932 B.n423 B.n31 163.367
R933 B.n423 B.n422 163.367
R934 B.n422 B.n421 163.367
R935 B.n421 B.n35 163.367
R936 B.n417 B.n35 163.367
R937 B.n417 B.n416 163.367
R938 B.n416 B.n415 163.367
R939 B.n415 B.n37 163.367
R940 B.n410 B.n37 163.367
R941 B.n410 B.n409 163.367
R942 B.n409 B.n408 163.367
R943 B.n408 B.n41 163.367
R944 B.n404 B.n41 163.367
R945 B.n404 B.n403 163.367
R946 B.n403 B.n402 163.367
R947 B.n402 B.n43 163.367
R948 B.n398 B.n43 163.367
R949 B.n398 B.n397 163.367
R950 B.n397 B.n396 163.367
R951 B.n396 B.n45 163.367
R952 B.n392 B.n45 163.367
R953 B.n392 B.n391 163.367
R954 B.n391 B.n390 163.367
R955 B.n390 B.n47 163.367
R956 B.n386 B.n47 163.367
R957 B.n386 B.n385 163.367
R958 B.n385 B.n384 163.367
R959 B.n384 B.n49 163.367
R960 B.n380 B.n49 163.367
R961 B.n380 B.n379 163.367
R962 B.n379 B.n378 163.367
R963 B.n378 B.n51 163.367
R964 B.n374 B.n51 163.367
R965 B.n374 B.n373 163.367
R966 B.n373 B.n372 163.367
R967 B.n372 B.n53 163.367
R968 B.n368 B.n53 163.367
R969 B.n368 B.n367 163.367
R970 B.n367 B.n366 163.367
R971 B.n366 B.n55 163.367
R972 B.n362 B.n55 163.367
R973 B.n362 B.n361 163.367
R974 B.n100 B.n99 59.5399
R975 B.n221 B.n107 59.5399
R976 B.n426 B.n33 59.5399
R977 B.n412 B.n39 59.5399
R978 B.n99 B.n98 52.946
R979 B.n107 B.n106 52.946
R980 B.n33 B.n32 52.946
R981 B.n39 B.n38 52.946
R982 B.n479 B.n14 36.3712
R983 B.n359 B.n56 36.3712
R984 B.n287 B.n286 36.3712
R985 B.n171 B.n124 36.3712
R986 B B.n515 18.0485
R987 B.n475 B.n14 10.6151
R988 B.n475 B.n474 10.6151
R989 B.n474 B.n473 10.6151
R990 B.n473 B.n16 10.6151
R991 B.n469 B.n16 10.6151
R992 B.n469 B.n468 10.6151
R993 B.n468 B.n467 10.6151
R994 B.n467 B.n18 10.6151
R995 B.n463 B.n18 10.6151
R996 B.n463 B.n462 10.6151
R997 B.n462 B.n461 10.6151
R998 B.n461 B.n20 10.6151
R999 B.n457 B.n20 10.6151
R1000 B.n457 B.n456 10.6151
R1001 B.n456 B.n455 10.6151
R1002 B.n455 B.n22 10.6151
R1003 B.n451 B.n22 10.6151
R1004 B.n451 B.n450 10.6151
R1005 B.n450 B.n449 10.6151
R1006 B.n449 B.n24 10.6151
R1007 B.n445 B.n24 10.6151
R1008 B.n445 B.n444 10.6151
R1009 B.n444 B.n443 10.6151
R1010 B.n443 B.n26 10.6151
R1011 B.n439 B.n26 10.6151
R1012 B.n439 B.n438 10.6151
R1013 B.n438 B.n437 10.6151
R1014 B.n437 B.n28 10.6151
R1015 B.n433 B.n28 10.6151
R1016 B.n433 B.n432 10.6151
R1017 B.n432 B.n431 10.6151
R1018 B.n431 B.n30 10.6151
R1019 B.n427 B.n30 10.6151
R1020 B.n425 B.n424 10.6151
R1021 B.n424 B.n34 10.6151
R1022 B.n420 B.n34 10.6151
R1023 B.n420 B.n419 10.6151
R1024 B.n419 B.n418 10.6151
R1025 B.n418 B.n36 10.6151
R1026 B.n414 B.n36 10.6151
R1027 B.n414 B.n413 10.6151
R1028 B.n411 B.n40 10.6151
R1029 B.n407 B.n40 10.6151
R1030 B.n407 B.n406 10.6151
R1031 B.n406 B.n405 10.6151
R1032 B.n405 B.n42 10.6151
R1033 B.n401 B.n42 10.6151
R1034 B.n401 B.n400 10.6151
R1035 B.n400 B.n399 10.6151
R1036 B.n399 B.n44 10.6151
R1037 B.n395 B.n44 10.6151
R1038 B.n395 B.n394 10.6151
R1039 B.n394 B.n393 10.6151
R1040 B.n393 B.n46 10.6151
R1041 B.n389 B.n46 10.6151
R1042 B.n389 B.n388 10.6151
R1043 B.n388 B.n387 10.6151
R1044 B.n387 B.n48 10.6151
R1045 B.n383 B.n48 10.6151
R1046 B.n383 B.n382 10.6151
R1047 B.n382 B.n381 10.6151
R1048 B.n381 B.n50 10.6151
R1049 B.n377 B.n50 10.6151
R1050 B.n377 B.n376 10.6151
R1051 B.n376 B.n375 10.6151
R1052 B.n375 B.n52 10.6151
R1053 B.n371 B.n52 10.6151
R1054 B.n371 B.n370 10.6151
R1055 B.n370 B.n369 10.6151
R1056 B.n369 B.n54 10.6151
R1057 B.n365 B.n54 10.6151
R1058 B.n365 B.n364 10.6151
R1059 B.n364 B.n363 10.6151
R1060 B.n363 B.n56 10.6151
R1061 B.n287 B.n80 10.6151
R1062 B.n291 B.n80 10.6151
R1063 B.n292 B.n291 10.6151
R1064 B.n293 B.n292 10.6151
R1065 B.n293 B.n78 10.6151
R1066 B.n297 B.n78 10.6151
R1067 B.n298 B.n297 10.6151
R1068 B.n299 B.n298 10.6151
R1069 B.n299 B.n76 10.6151
R1070 B.n303 B.n76 10.6151
R1071 B.n304 B.n303 10.6151
R1072 B.n305 B.n304 10.6151
R1073 B.n305 B.n74 10.6151
R1074 B.n309 B.n74 10.6151
R1075 B.n310 B.n309 10.6151
R1076 B.n311 B.n310 10.6151
R1077 B.n311 B.n72 10.6151
R1078 B.n315 B.n72 10.6151
R1079 B.n316 B.n315 10.6151
R1080 B.n317 B.n316 10.6151
R1081 B.n317 B.n70 10.6151
R1082 B.n321 B.n70 10.6151
R1083 B.n322 B.n321 10.6151
R1084 B.n323 B.n322 10.6151
R1085 B.n323 B.n68 10.6151
R1086 B.n327 B.n68 10.6151
R1087 B.n328 B.n327 10.6151
R1088 B.n329 B.n328 10.6151
R1089 B.n329 B.n66 10.6151
R1090 B.n333 B.n66 10.6151
R1091 B.n334 B.n333 10.6151
R1092 B.n335 B.n334 10.6151
R1093 B.n335 B.n64 10.6151
R1094 B.n339 B.n64 10.6151
R1095 B.n340 B.n339 10.6151
R1096 B.n341 B.n340 10.6151
R1097 B.n341 B.n62 10.6151
R1098 B.n345 B.n62 10.6151
R1099 B.n346 B.n345 10.6151
R1100 B.n347 B.n346 10.6151
R1101 B.n347 B.n60 10.6151
R1102 B.n351 B.n60 10.6151
R1103 B.n352 B.n351 10.6151
R1104 B.n353 B.n352 10.6151
R1105 B.n353 B.n58 10.6151
R1106 B.n357 B.n58 10.6151
R1107 B.n358 B.n357 10.6151
R1108 B.n359 B.n358 10.6151
R1109 B.n172 B.n171 10.6151
R1110 B.n173 B.n172 10.6151
R1111 B.n173 B.n122 10.6151
R1112 B.n177 B.n122 10.6151
R1113 B.n178 B.n177 10.6151
R1114 B.n179 B.n178 10.6151
R1115 B.n179 B.n120 10.6151
R1116 B.n183 B.n120 10.6151
R1117 B.n184 B.n183 10.6151
R1118 B.n185 B.n184 10.6151
R1119 B.n185 B.n118 10.6151
R1120 B.n189 B.n118 10.6151
R1121 B.n190 B.n189 10.6151
R1122 B.n191 B.n190 10.6151
R1123 B.n191 B.n116 10.6151
R1124 B.n195 B.n116 10.6151
R1125 B.n196 B.n195 10.6151
R1126 B.n197 B.n196 10.6151
R1127 B.n197 B.n114 10.6151
R1128 B.n201 B.n114 10.6151
R1129 B.n202 B.n201 10.6151
R1130 B.n203 B.n202 10.6151
R1131 B.n203 B.n112 10.6151
R1132 B.n207 B.n112 10.6151
R1133 B.n208 B.n207 10.6151
R1134 B.n209 B.n208 10.6151
R1135 B.n209 B.n110 10.6151
R1136 B.n213 B.n110 10.6151
R1137 B.n214 B.n213 10.6151
R1138 B.n215 B.n214 10.6151
R1139 B.n215 B.n108 10.6151
R1140 B.n219 B.n108 10.6151
R1141 B.n220 B.n219 10.6151
R1142 B.n222 B.n104 10.6151
R1143 B.n226 B.n104 10.6151
R1144 B.n227 B.n226 10.6151
R1145 B.n228 B.n227 10.6151
R1146 B.n228 B.n102 10.6151
R1147 B.n232 B.n102 10.6151
R1148 B.n233 B.n232 10.6151
R1149 B.n234 B.n233 10.6151
R1150 B.n238 B.n237 10.6151
R1151 B.n239 B.n238 10.6151
R1152 B.n239 B.n96 10.6151
R1153 B.n243 B.n96 10.6151
R1154 B.n244 B.n243 10.6151
R1155 B.n245 B.n244 10.6151
R1156 B.n245 B.n94 10.6151
R1157 B.n249 B.n94 10.6151
R1158 B.n250 B.n249 10.6151
R1159 B.n251 B.n250 10.6151
R1160 B.n251 B.n92 10.6151
R1161 B.n255 B.n92 10.6151
R1162 B.n256 B.n255 10.6151
R1163 B.n257 B.n256 10.6151
R1164 B.n257 B.n90 10.6151
R1165 B.n261 B.n90 10.6151
R1166 B.n262 B.n261 10.6151
R1167 B.n263 B.n262 10.6151
R1168 B.n263 B.n88 10.6151
R1169 B.n267 B.n88 10.6151
R1170 B.n268 B.n267 10.6151
R1171 B.n269 B.n268 10.6151
R1172 B.n269 B.n86 10.6151
R1173 B.n273 B.n86 10.6151
R1174 B.n274 B.n273 10.6151
R1175 B.n275 B.n274 10.6151
R1176 B.n275 B.n84 10.6151
R1177 B.n279 B.n84 10.6151
R1178 B.n280 B.n279 10.6151
R1179 B.n281 B.n280 10.6151
R1180 B.n281 B.n82 10.6151
R1181 B.n285 B.n82 10.6151
R1182 B.n286 B.n285 10.6151
R1183 B.n167 B.n124 10.6151
R1184 B.n167 B.n166 10.6151
R1185 B.n166 B.n165 10.6151
R1186 B.n165 B.n126 10.6151
R1187 B.n161 B.n126 10.6151
R1188 B.n161 B.n160 10.6151
R1189 B.n160 B.n159 10.6151
R1190 B.n159 B.n128 10.6151
R1191 B.n155 B.n128 10.6151
R1192 B.n155 B.n154 10.6151
R1193 B.n154 B.n153 10.6151
R1194 B.n153 B.n130 10.6151
R1195 B.n149 B.n130 10.6151
R1196 B.n149 B.n148 10.6151
R1197 B.n148 B.n147 10.6151
R1198 B.n147 B.n132 10.6151
R1199 B.n143 B.n132 10.6151
R1200 B.n143 B.n142 10.6151
R1201 B.n142 B.n141 10.6151
R1202 B.n141 B.n134 10.6151
R1203 B.n137 B.n134 10.6151
R1204 B.n137 B.n136 10.6151
R1205 B.n136 B.n0 10.6151
R1206 B.n511 B.n1 10.6151
R1207 B.n511 B.n510 10.6151
R1208 B.n510 B.n509 10.6151
R1209 B.n509 B.n4 10.6151
R1210 B.n505 B.n4 10.6151
R1211 B.n505 B.n504 10.6151
R1212 B.n504 B.n503 10.6151
R1213 B.n503 B.n6 10.6151
R1214 B.n499 B.n6 10.6151
R1215 B.n499 B.n498 10.6151
R1216 B.n498 B.n497 10.6151
R1217 B.n497 B.n8 10.6151
R1218 B.n493 B.n8 10.6151
R1219 B.n493 B.n492 10.6151
R1220 B.n492 B.n491 10.6151
R1221 B.n491 B.n10 10.6151
R1222 B.n487 B.n10 10.6151
R1223 B.n487 B.n486 10.6151
R1224 B.n486 B.n485 10.6151
R1225 B.n485 B.n12 10.6151
R1226 B.n481 B.n12 10.6151
R1227 B.n481 B.n480 10.6151
R1228 B.n480 B.n479 10.6151
R1229 B.n426 B.n425 6.5566
R1230 B.n413 B.n412 6.5566
R1231 B.n222 B.n221 6.5566
R1232 B.n234 B.n100 6.5566
R1233 B.n427 B.n426 4.05904
R1234 B.n412 B.n411 4.05904
R1235 B.n221 B.n220 4.05904
R1236 B.n237 B.n100 4.05904
R1237 B.n515 B.n0 2.81026
R1238 B.n515 B.n1 2.81026
R1239 VN VN.t0 185.555
R1240 VN VN.t1 143.654
R1241 VDD2.n93 VDD2.n49 756.745
R1242 VDD2.n44 VDD2.n0 756.745
R1243 VDD2.n94 VDD2.n93 585
R1244 VDD2.n92 VDD2.n91 585
R1245 VDD2.n53 VDD2.n52 585
R1246 VDD2.n57 VDD2.n55 585
R1247 VDD2.n86 VDD2.n85 585
R1248 VDD2.n84 VDD2.n83 585
R1249 VDD2.n59 VDD2.n58 585
R1250 VDD2.n78 VDD2.n77 585
R1251 VDD2.n76 VDD2.n75 585
R1252 VDD2.n63 VDD2.n62 585
R1253 VDD2.n70 VDD2.n69 585
R1254 VDD2.n68 VDD2.n67 585
R1255 VDD2.n17 VDD2.n16 585
R1256 VDD2.n19 VDD2.n18 585
R1257 VDD2.n12 VDD2.n11 585
R1258 VDD2.n25 VDD2.n24 585
R1259 VDD2.n27 VDD2.n26 585
R1260 VDD2.n8 VDD2.n7 585
R1261 VDD2.n34 VDD2.n33 585
R1262 VDD2.n35 VDD2.n6 585
R1263 VDD2.n37 VDD2.n36 585
R1264 VDD2.n4 VDD2.n3 585
R1265 VDD2.n43 VDD2.n42 585
R1266 VDD2.n45 VDD2.n44 585
R1267 VDD2.n66 VDD2.t1 329.038
R1268 VDD2.n15 VDD2.t0 329.038
R1269 VDD2.n93 VDD2.n92 171.744
R1270 VDD2.n92 VDD2.n52 171.744
R1271 VDD2.n57 VDD2.n52 171.744
R1272 VDD2.n85 VDD2.n57 171.744
R1273 VDD2.n85 VDD2.n84 171.744
R1274 VDD2.n84 VDD2.n58 171.744
R1275 VDD2.n77 VDD2.n58 171.744
R1276 VDD2.n77 VDD2.n76 171.744
R1277 VDD2.n76 VDD2.n62 171.744
R1278 VDD2.n69 VDD2.n62 171.744
R1279 VDD2.n69 VDD2.n68 171.744
R1280 VDD2.n18 VDD2.n17 171.744
R1281 VDD2.n18 VDD2.n11 171.744
R1282 VDD2.n25 VDD2.n11 171.744
R1283 VDD2.n26 VDD2.n25 171.744
R1284 VDD2.n26 VDD2.n7 171.744
R1285 VDD2.n34 VDD2.n7 171.744
R1286 VDD2.n35 VDD2.n34 171.744
R1287 VDD2.n36 VDD2.n35 171.744
R1288 VDD2.n36 VDD2.n3 171.744
R1289 VDD2.n43 VDD2.n3 171.744
R1290 VDD2.n44 VDD2.n43 171.744
R1291 VDD2.n98 VDD2.n48 88.0318
R1292 VDD2.n68 VDD2.t1 85.8723
R1293 VDD2.n17 VDD2.t0 85.8723
R1294 VDD2.n98 VDD2.n97 51.5793
R1295 VDD2.n55 VDD2.n53 13.1884
R1296 VDD2.n37 VDD2.n4 13.1884
R1297 VDD2.n91 VDD2.n90 12.8005
R1298 VDD2.n87 VDD2.n86 12.8005
R1299 VDD2.n38 VDD2.n6 12.8005
R1300 VDD2.n42 VDD2.n41 12.8005
R1301 VDD2.n94 VDD2.n51 12.0247
R1302 VDD2.n83 VDD2.n56 12.0247
R1303 VDD2.n33 VDD2.n32 12.0247
R1304 VDD2.n45 VDD2.n2 12.0247
R1305 VDD2.n95 VDD2.n49 11.249
R1306 VDD2.n82 VDD2.n59 11.249
R1307 VDD2.n31 VDD2.n8 11.249
R1308 VDD2.n46 VDD2.n0 11.249
R1309 VDD2.n67 VDD2.n66 10.7239
R1310 VDD2.n16 VDD2.n15 10.7239
R1311 VDD2.n79 VDD2.n78 10.4732
R1312 VDD2.n28 VDD2.n27 10.4732
R1313 VDD2.n75 VDD2.n61 9.69747
R1314 VDD2.n24 VDD2.n10 9.69747
R1315 VDD2.n97 VDD2.n96 9.45567
R1316 VDD2.n48 VDD2.n47 9.45567
R1317 VDD2.n65 VDD2.n64 9.3005
R1318 VDD2.n72 VDD2.n71 9.3005
R1319 VDD2.n74 VDD2.n73 9.3005
R1320 VDD2.n61 VDD2.n60 9.3005
R1321 VDD2.n80 VDD2.n79 9.3005
R1322 VDD2.n82 VDD2.n81 9.3005
R1323 VDD2.n56 VDD2.n54 9.3005
R1324 VDD2.n88 VDD2.n87 9.3005
R1325 VDD2.n96 VDD2.n95 9.3005
R1326 VDD2.n51 VDD2.n50 9.3005
R1327 VDD2.n90 VDD2.n89 9.3005
R1328 VDD2.n47 VDD2.n46 9.3005
R1329 VDD2.n2 VDD2.n1 9.3005
R1330 VDD2.n41 VDD2.n40 9.3005
R1331 VDD2.n14 VDD2.n13 9.3005
R1332 VDD2.n21 VDD2.n20 9.3005
R1333 VDD2.n23 VDD2.n22 9.3005
R1334 VDD2.n10 VDD2.n9 9.3005
R1335 VDD2.n29 VDD2.n28 9.3005
R1336 VDD2.n31 VDD2.n30 9.3005
R1337 VDD2.n32 VDD2.n5 9.3005
R1338 VDD2.n39 VDD2.n38 9.3005
R1339 VDD2.n74 VDD2.n63 8.92171
R1340 VDD2.n23 VDD2.n12 8.92171
R1341 VDD2.n71 VDD2.n70 8.14595
R1342 VDD2.n20 VDD2.n19 8.14595
R1343 VDD2.n67 VDD2.n65 7.3702
R1344 VDD2.n16 VDD2.n14 7.3702
R1345 VDD2.n70 VDD2.n65 5.81868
R1346 VDD2.n19 VDD2.n14 5.81868
R1347 VDD2.n71 VDD2.n63 5.04292
R1348 VDD2.n20 VDD2.n12 5.04292
R1349 VDD2.n75 VDD2.n74 4.26717
R1350 VDD2.n24 VDD2.n23 4.26717
R1351 VDD2.n78 VDD2.n61 3.49141
R1352 VDD2.n27 VDD2.n10 3.49141
R1353 VDD2.n97 VDD2.n49 2.71565
R1354 VDD2.n79 VDD2.n59 2.71565
R1355 VDD2.n28 VDD2.n8 2.71565
R1356 VDD2.n48 VDD2.n0 2.71565
R1357 VDD2.n66 VDD2.n64 2.41283
R1358 VDD2.n15 VDD2.n13 2.41283
R1359 VDD2.n95 VDD2.n94 1.93989
R1360 VDD2.n83 VDD2.n82 1.93989
R1361 VDD2.n33 VDD2.n31 1.93989
R1362 VDD2.n46 VDD2.n45 1.93989
R1363 VDD2.n91 VDD2.n51 1.16414
R1364 VDD2.n86 VDD2.n56 1.16414
R1365 VDD2.n32 VDD2.n6 1.16414
R1366 VDD2.n42 VDD2.n2 1.16414
R1367 VDD2 VDD2.n98 0.647052
R1368 VDD2.n90 VDD2.n53 0.388379
R1369 VDD2.n87 VDD2.n55 0.388379
R1370 VDD2.n38 VDD2.n37 0.388379
R1371 VDD2.n41 VDD2.n4 0.388379
R1372 VDD2.n96 VDD2.n50 0.155672
R1373 VDD2.n89 VDD2.n50 0.155672
R1374 VDD2.n89 VDD2.n88 0.155672
R1375 VDD2.n88 VDD2.n54 0.155672
R1376 VDD2.n81 VDD2.n54 0.155672
R1377 VDD2.n81 VDD2.n80 0.155672
R1378 VDD2.n80 VDD2.n60 0.155672
R1379 VDD2.n73 VDD2.n60 0.155672
R1380 VDD2.n73 VDD2.n72 0.155672
R1381 VDD2.n72 VDD2.n64 0.155672
R1382 VDD2.n21 VDD2.n13 0.155672
R1383 VDD2.n22 VDD2.n21 0.155672
R1384 VDD2.n22 VDD2.n9 0.155672
R1385 VDD2.n29 VDD2.n9 0.155672
R1386 VDD2.n30 VDD2.n29 0.155672
R1387 VDD2.n30 VDD2.n5 0.155672
R1388 VDD2.n39 VDD2.n5 0.155672
R1389 VDD2.n40 VDD2.n39 0.155672
R1390 VDD2.n40 VDD2.n1 0.155672
R1391 VDD2.n47 VDD2.n1 0.155672
C0 w_n2062_n2844# B 7.85881f
C1 VDD1 w_n2062_n2844# 1.57602f
C2 VDD1 B 1.47332f
C3 VTAIL w_n2062_n2844# 2.3947f
C4 VN VDD2 2.19956f
C5 VP VDD2 0.324119f
C6 VTAIL B 2.99705f
C7 VDD1 VTAIL 4.3396f
C8 VP VN 4.87934f
C9 w_n2062_n2844# VDD2 1.59952f
C10 VDD2 B 1.50163f
C11 VDD1 VDD2 0.650352f
C12 VN w_n2062_n2844# 2.7869f
C13 VP w_n2062_n2844# 3.04913f
C14 VN B 0.981766f
C15 VP B 1.41208f
C16 VTAIL VDD2 4.3893f
C17 VDD1 VN 0.147696f
C18 VDD1 VP 2.37383f
C19 VN VTAIL 1.96508f
C20 VP VTAIL 1.97934f
C21 VDD2 VSUBS 0.790087f
C22 VDD1 VSUBS 3.350612f
C23 VTAIL VSUBS 0.84915f
C24 VN VSUBS 6.46578f
C25 VP VSUBS 1.521497f
C26 B VSUBS 3.537472f
C27 w_n2062_n2844# VSUBS 72.524704f
C28 VDD2.n0 VSUBS 0.022256f
C29 VDD2.n1 VSUBS 0.020492f
C30 VDD2.n2 VSUBS 0.011011f
C31 VDD2.n3 VSUBS 0.026027f
C32 VDD2.n4 VSUBS 0.011335f
C33 VDD2.n5 VSUBS 0.020492f
C34 VDD2.n6 VSUBS 0.011659f
C35 VDD2.n7 VSUBS 0.026027f
C36 VDD2.n8 VSUBS 0.011659f
C37 VDD2.n9 VSUBS 0.020492f
C38 VDD2.n10 VSUBS 0.011011f
C39 VDD2.n11 VSUBS 0.026027f
C40 VDD2.n12 VSUBS 0.011659f
C41 VDD2.n13 VSUBS 0.77151f
C42 VDD2.n14 VSUBS 0.011011f
C43 VDD2.t0 VSUBS 0.055938f
C44 VDD2.n15 VSUBS 0.137137f
C45 VDD2.n16 VSUBS 0.019579f
C46 VDD2.n17 VSUBS 0.01952f
C47 VDD2.n18 VSUBS 0.026027f
C48 VDD2.n19 VSUBS 0.011659f
C49 VDD2.n20 VSUBS 0.011011f
C50 VDD2.n21 VSUBS 0.020492f
C51 VDD2.n22 VSUBS 0.020492f
C52 VDD2.n23 VSUBS 0.011011f
C53 VDD2.n24 VSUBS 0.011659f
C54 VDD2.n25 VSUBS 0.026027f
C55 VDD2.n26 VSUBS 0.026027f
C56 VDD2.n27 VSUBS 0.011659f
C57 VDD2.n28 VSUBS 0.011011f
C58 VDD2.n29 VSUBS 0.020492f
C59 VDD2.n30 VSUBS 0.020492f
C60 VDD2.n31 VSUBS 0.011011f
C61 VDD2.n32 VSUBS 0.011011f
C62 VDD2.n33 VSUBS 0.011659f
C63 VDD2.n34 VSUBS 0.026027f
C64 VDD2.n35 VSUBS 0.026027f
C65 VDD2.n36 VSUBS 0.026027f
C66 VDD2.n37 VSUBS 0.011335f
C67 VDD2.n38 VSUBS 0.011011f
C68 VDD2.n39 VSUBS 0.020492f
C69 VDD2.n40 VSUBS 0.020492f
C70 VDD2.n41 VSUBS 0.011011f
C71 VDD2.n42 VSUBS 0.011659f
C72 VDD2.n43 VSUBS 0.026027f
C73 VDD2.n44 VSUBS 0.062124f
C74 VDD2.n45 VSUBS 0.011659f
C75 VDD2.n46 VSUBS 0.011011f
C76 VDD2.n47 VSUBS 0.051284f
C77 VDD2.n48 VSUBS 0.504155f
C78 VDD2.n49 VSUBS 0.022256f
C79 VDD2.n50 VSUBS 0.020492f
C80 VDD2.n51 VSUBS 0.011011f
C81 VDD2.n52 VSUBS 0.026027f
C82 VDD2.n53 VSUBS 0.011335f
C83 VDD2.n54 VSUBS 0.020492f
C84 VDD2.n55 VSUBS 0.011335f
C85 VDD2.n56 VSUBS 0.011011f
C86 VDD2.n57 VSUBS 0.026027f
C87 VDD2.n58 VSUBS 0.026027f
C88 VDD2.n59 VSUBS 0.011659f
C89 VDD2.n60 VSUBS 0.020492f
C90 VDD2.n61 VSUBS 0.011011f
C91 VDD2.n62 VSUBS 0.026027f
C92 VDD2.n63 VSUBS 0.011659f
C93 VDD2.n64 VSUBS 0.77151f
C94 VDD2.n65 VSUBS 0.011011f
C95 VDD2.t1 VSUBS 0.055938f
C96 VDD2.n66 VSUBS 0.137137f
C97 VDD2.n67 VSUBS 0.019579f
C98 VDD2.n68 VSUBS 0.01952f
C99 VDD2.n69 VSUBS 0.026027f
C100 VDD2.n70 VSUBS 0.011659f
C101 VDD2.n71 VSUBS 0.011011f
C102 VDD2.n72 VSUBS 0.020492f
C103 VDD2.n73 VSUBS 0.020492f
C104 VDD2.n74 VSUBS 0.011011f
C105 VDD2.n75 VSUBS 0.011659f
C106 VDD2.n76 VSUBS 0.026027f
C107 VDD2.n77 VSUBS 0.026027f
C108 VDD2.n78 VSUBS 0.011659f
C109 VDD2.n79 VSUBS 0.011011f
C110 VDD2.n80 VSUBS 0.020492f
C111 VDD2.n81 VSUBS 0.020492f
C112 VDD2.n82 VSUBS 0.011011f
C113 VDD2.n83 VSUBS 0.011659f
C114 VDD2.n84 VSUBS 0.026027f
C115 VDD2.n85 VSUBS 0.026027f
C116 VDD2.n86 VSUBS 0.011659f
C117 VDD2.n87 VSUBS 0.011011f
C118 VDD2.n88 VSUBS 0.020492f
C119 VDD2.n89 VSUBS 0.020492f
C120 VDD2.n90 VSUBS 0.011011f
C121 VDD2.n91 VSUBS 0.011659f
C122 VDD2.n92 VSUBS 0.026027f
C123 VDD2.n93 VSUBS 0.062124f
C124 VDD2.n94 VSUBS 0.011659f
C125 VDD2.n95 VSUBS 0.011011f
C126 VDD2.n96 VSUBS 0.051284f
C127 VDD2.n97 VSUBS 0.045439f
C128 VDD2.n98 VSUBS 2.26392f
C129 VN.t1 VSUBS 2.57463f
C130 VN.t0 VSUBS 3.10751f
C131 B.n0 VSUBS 0.004272f
C132 B.n1 VSUBS 0.004272f
C133 B.n2 VSUBS 0.006756f
C134 B.n3 VSUBS 0.006756f
C135 B.n4 VSUBS 0.006756f
C136 B.n5 VSUBS 0.006756f
C137 B.n6 VSUBS 0.006756f
C138 B.n7 VSUBS 0.006756f
C139 B.n8 VSUBS 0.006756f
C140 B.n9 VSUBS 0.006756f
C141 B.n10 VSUBS 0.006756f
C142 B.n11 VSUBS 0.006756f
C143 B.n12 VSUBS 0.006756f
C144 B.n13 VSUBS 0.006756f
C145 B.n14 VSUBS 0.017313f
C146 B.n15 VSUBS 0.006756f
C147 B.n16 VSUBS 0.006756f
C148 B.n17 VSUBS 0.006756f
C149 B.n18 VSUBS 0.006756f
C150 B.n19 VSUBS 0.006756f
C151 B.n20 VSUBS 0.006756f
C152 B.n21 VSUBS 0.006756f
C153 B.n22 VSUBS 0.006756f
C154 B.n23 VSUBS 0.006756f
C155 B.n24 VSUBS 0.006756f
C156 B.n25 VSUBS 0.006756f
C157 B.n26 VSUBS 0.006756f
C158 B.n27 VSUBS 0.006756f
C159 B.n28 VSUBS 0.006756f
C160 B.n29 VSUBS 0.006756f
C161 B.n30 VSUBS 0.006756f
C162 B.n31 VSUBS 0.006756f
C163 B.t11 VSUBS 0.149201f
C164 B.t10 VSUBS 0.176359f
C165 B.t9 VSUBS 0.999162f
C166 B.n32 VSUBS 0.287489f
C167 B.n33 VSUBS 0.205299f
C168 B.n34 VSUBS 0.006756f
C169 B.n35 VSUBS 0.006756f
C170 B.n36 VSUBS 0.006756f
C171 B.n37 VSUBS 0.006756f
C172 B.t8 VSUBS 0.149203f
C173 B.t7 VSUBS 0.176361f
C174 B.t6 VSUBS 0.999162f
C175 B.n38 VSUBS 0.287487f
C176 B.n39 VSUBS 0.205297f
C177 B.n40 VSUBS 0.006756f
C178 B.n41 VSUBS 0.006756f
C179 B.n42 VSUBS 0.006756f
C180 B.n43 VSUBS 0.006756f
C181 B.n44 VSUBS 0.006756f
C182 B.n45 VSUBS 0.006756f
C183 B.n46 VSUBS 0.006756f
C184 B.n47 VSUBS 0.006756f
C185 B.n48 VSUBS 0.006756f
C186 B.n49 VSUBS 0.006756f
C187 B.n50 VSUBS 0.006756f
C188 B.n51 VSUBS 0.006756f
C189 B.n52 VSUBS 0.006756f
C190 B.n53 VSUBS 0.006756f
C191 B.n54 VSUBS 0.006756f
C192 B.n55 VSUBS 0.006756f
C193 B.n56 VSUBS 0.016596f
C194 B.n57 VSUBS 0.006756f
C195 B.n58 VSUBS 0.006756f
C196 B.n59 VSUBS 0.006756f
C197 B.n60 VSUBS 0.006756f
C198 B.n61 VSUBS 0.006756f
C199 B.n62 VSUBS 0.006756f
C200 B.n63 VSUBS 0.006756f
C201 B.n64 VSUBS 0.006756f
C202 B.n65 VSUBS 0.006756f
C203 B.n66 VSUBS 0.006756f
C204 B.n67 VSUBS 0.006756f
C205 B.n68 VSUBS 0.006756f
C206 B.n69 VSUBS 0.006756f
C207 B.n70 VSUBS 0.006756f
C208 B.n71 VSUBS 0.006756f
C209 B.n72 VSUBS 0.006756f
C210 B.n73 VSUBS 0.006756f
C211 B.n74 VSUBS 0.006756f
C212 B.n75 VSUBS 0.006756f
C213 B.n76 VSUBS 0.006756f
C214 B.n77 VSUBS 0.006756f
C215 B.n78 VSUBS 0.006756f
C216 B.n79 VSUBS 0.006756f
C217 B.n80 VSUBS 0.006756f
C218 B.n81 VSUBS 0.017313f
C219 B.n82 VSUBS 0.006756f
C220 B.n83 VSUBS 0.006756f
C221 B.n84 VSUBS 0.006756f
C222 B.n85 VSUBS 0.006756f
C223 B.n86 VSUBS 0.006756f
C224 B.n87 VSUBS 0.006756f
C225 B.n88 VSUBS 0.006756f
C226 B.n89 VSUBS 0.006756f
C227 B.n90 VSUBS 0.006756f
C228 B.n91 VSUBS 0.006756f
C229 B.n92 VSUBS 0.006756f
C230 B.n93 VSUBS 0.006756f
C231 B.n94 VSUBS 0.006756f
C232 B.n95 VSUBS 0.006756f
C233 B.n96 VSUBS 0.006756f
C234 B.n97 VSUBS 0.006756f
C235 B.t4 VSUBS 0.149203f
C236 B.t5 VSUBS 0.176361f
C237 B.t3 VSUBS 0.999162f
C238 B.n98 VSUBS 0.287487f
C239 B.n99 VSUBS 0.205297f
C240 B.n100 VSUBS 0.015653f
C241 B.n101 VSUBS 0.006756f
C242 B.n102 VSUBS 0.006756f
C243 B.n103 VSUBS 0.006756f
C244 B.n104 VSUBS 0.006756f
C245 B.n105 VSUBS 0.006756f
C246 B.t1 VSUBS 0.149201f
C247 B.t2 VSUBS 0.176359f
C248 B.t0 VSUBS 0.999162f
C249 B.n106 VSUBS 0.287489f
C250 B.n107 VSUBS 0.205299f
C251 B.n108 VSUBS 0.006756f
C252 B.n109 VSUBS 0.006756f
C253 B.n110 VSUBS 0.006756f
C254 B.n111 VSUBS 0.006756f
C255 B.n112 VSUBS 0.006756f
C256 B.n113 VSUBS 0.006756f
C257 B.n114 VSUBS 0.006756f
C258 B.n115 VSUBS 0.006756f
C259 B.n116 VSUBS 0.006756f
C260 B.n117 VSUBS 0.006756f
C261 B.n118 VSUBS 0.006756f
C262 B.n119 VSUBS 0.006756f
C263 B.n120 VSUBS 0.006756f
C264 B.n121 VSUBS 0.006756f
C265 B.n122 VSUBS 0.006756f
C266 B.n123 VSUBS 0.006756f
C267 B.n124 VSUBS 0.016666f
C268 B.n125 VSUBS 0.006756f
C269 B.n126 VSUBS 0.006756f
C270 B.n127 VSUBS 0.006756f
C271 B.n128 VSUBS 0.006756f
C272 B.n129 VSUBS 0.006756f
C273 B.n130 VSUBS 0.006756f
C274 B.n131 VSUBS 0.006756f
C275 B.n132 VSUBS 0.006756f
C276 B.n133 VSUBS 0.006756f
C277 B.n134 VSUBS 0.006756f
C278 B.n135 VSUBS 0.006756f
C279 B.n136 VSUBS 0.006756f
C280 B.n137 VSUBS 0.006756f
C281 B.n138 VSUBS 0.006756f
C282 B.n139 VSUBS 0.006756f
C283 B.n140 VSUBS 0.006756f
C284 B.n141 VSUBS 0.006756f
C285 B.n142 VSUBS 0.006756f
C286 B.n143 VSUBS 0.006756f
C287 B.n144 VSUBS 0.006756f
C288 B.n145 VSUBS 0.006756f
C289 B.n146 VSUBS 0.006756f
C290 B.n147 VSUBS 0.006756f
C291 B.n148 VSUBS 0.006756f
C292 B.n149 VSUBS 0.006756f
C293 B.n150 VSUBS 0.006756f
C294 B.n151 VSUBS 0.006756f
C295 B.n152 VSUBS 0.006756f
C296 B.n153 VSUBS 0.006756f
C297 B.n154 VSUBS 0.006756f
C298 B.n155 VSUBS 0.006756f
C299 B.n156 VSUBS 0.006756f
C300 B.n157 VSUBS 0.006756f
C301 B.n158 VSUBS 0.006756f
C302 B.n159 VSUBS 0.006756f
C303 B.n160 VSUBS 0.006756f
C304 B.n161 VSUBS 0.006756f
C305 B.n162 VSUBS 0.006756f
C306 B.n163 VSUBS 0.006756f
C307 B.n164 VSUBS 0.006756f
C308 B.n165 VSUBS 0.006756f
C309 B.n166 VSUBS 0.006756f
C310 B.n167 VSUBS 0.006756f
C311 B.n168 VSUBS 0.006756f
C312 B.n169 VSUBS 0.016666f
C313 B.n170 VSUBS 0.017313f
C314 B.n171 VSUBS 0.017313f
C315 B.n172 VSUBS 0.006756f
C316 B.n173 VSUBS 0.006756f
C317 B.n174 VSUBS 0.006756f
C318 B.n175 VSUBS 0.006756f
C319 B.n176 VSUBS 0.006756f
C320 B.n177 VSUBS 0.006756f
C321 B.n178 VSUBS 0.006756f
C322 B.n179 VSUBS 0.006756f
C323 B.n180 VSUBS 0.006756f
C324 B.n181 VSUBS 0.006756f
C325 B.n182 VSUBS 0.006756f
C326 B.n183 VSUBS 0.006756f
C327 B.n184 VSUBS 0.006756f
C328 B.n185 VSUBS 0.006756f
C329 B.n186 VSUBS 0.006756f
C330 B.n187 VSUBS 0.006756f
C331 B.n188 VSUBS 0.006756f
C332 B.n189 VSUBS 0.006756f
C333 B.n190 VSUBS 0.006756f
C334 B.n191 VSUBS 0.006756f
C335 B.n192 VSUBS 0.006756f
C336 B.n193 VSUBS 0.006756f
C337 B.n194 VSUBS 0.006756f
C338 B.n195 VSUBS 0.006756f
C339 B.n196 VSUBS 0.006756f
C340 B.n197 VSUBS 0.006756f
C341 B.n198 VSUBS 0.006756f
C342 B.n199 VSUBS 0.006756f
C343 B.n200 VSUBS 0.006756f
C344 B.n201 VSUBS 0.006756f
C345 B.n202 VSUBS 0.006756f
C346 B.n203 VSUBS 0.006756f
C347 B.n204 VSUBS 0.006756f
C348 B.n205 VSUBS 0.006756f
C349 B.n206 VSUBS 0.006756f
C350 B.n207 VSUBS 0.006756f
C351 B.n208 VSUBS 0.006756f
C352 B.n209 VSUBS 0.006756f
C353 B.n210 VSUBS 0.006756f
C354 B.n211 VSUBS 0.006756f
C355 B.n212 VSUBS 0.006756f
C356 B.n213 VSUBS 0.006756f
C357 B.n214 VSUBS 0.006756f
C358 B.n215 VSUBS 0.006756f
C359 B.n216 VSUBS 0.006756f
C360 B.n217 VSUBS 0.006756f
C361 B.n218 VSUBS 0.006756f
C362 B.n219 VSUBS 0.006756f
C363 B.n220 VSUBS 0.00467f
C364 B.n221 VSUBS 0.015653f
C365 B.n222 VSUBS 0.005464f
C366 B.n223 VSUBS 0.006756f
C367 B.n224 VSUBS 0.006756f
C368 B.n225 VSUBS 0.006756f
C369 B.n226 VSUBS 0.006756f
C370 B.n227 VSUBS 0.006756f
C371 B.n228 VSUBS 0.006756f
C372 B.n229 VSUBS 0.006756f
C373 B.n230 VSUBS 0.006756f
C374 B.n231 VSUBS 0.006756f
C375 B.n232 VSUBS 0.006756f
C376 B.n233 VSUBS 0.006756f
C377 B.n234 VSUBS 0.005464f
C378 B.n235 VSUBS 0.006756f
C379 B.n236 VSUBS 0.006756f
C380 B.n237 VSUBS 0.00467f
C381 B.n238 VSUBS 0.006756f
C382 B.n239 VSUBS 0.006756f
C383 B.n240 VSUBS 0.006756f
C384 B.n241 VSUBS 0.006756f
C385 B.n242 VSUBS 0.006756f
C386 B.n243 VSUBS 0.006756f
C387 B.n244 VSUBS 0.006756f
C388 B.n245 VSUBS 0.006756f
C389 B.n246 VSUBS 0.006756f
C390 B.n247 VSUBS 0.006756f
C391 B.n248 VSUBS 0.006756f
C392 B.n249 VSUBS 0.006756f
C393 B.n250 VSUBS 0.006756f
C394 B.n251 VSUBS 0.006756f
C395 B.n252 VSUBS 0.006756f
C396 B.n253 VSUBS 0.006756f
C397 B.n254 VSUBS 0.006756f
C398 B.n255 VSUBS 0.006756f
C399 B.n256 VSUBS 0.006756f
C400 B.n257 VSUBS 0.006756f
C401 B.n258 VSUBS 0.006756f
C402 B.n259 VSUBS 0.006756f
C403 B.n260 VSUBS 0.006756f
C404 B.n261 VSUBS 0.006756f
C405 B.n262 VSUBS 0.006756f
C406 B.n263 VSUBS 0.006756f
C407 B.n264 VSUBS 0.006756f
C408 B.n265 VSUBS 0.006756f
C409 B.n266 VSUBS 0.006756f
C410 B.n267 VSUBS 0.006756f
C411 B.n268 VSUBS 0.006756f
C412 B.n269 VSUBS 0.006756f
C413 B.n270 VSUBS 0.006756f
C414 B.n271 VSUBS 0.006756f
C415 B.n272 VSUBS 0.006756f
C416 B.n273 VSUBS 0.006756f
C417 B.n274 VSUBS 0.006756f
C418 B.n275 VSUBS 0.006756f
C419 B.n276 VSUBS 0.006756f
C420 B.n277 VSUBS 0.006756f
C421 B.n278 VSUBS 0.006756f
C422 B.n279 VSUBS 0.006756f
C423 B.n280 VSUBS 0.006756f
C424 B.n281 VSUBS 0.006756f
C425 B.n282 VSUBS 0.006756f
C426 B.n283 VSUBS 0.006756f
C427 B.n284 VSUBS 0.006756f
C428 B.n285 VSUBS 0.006756f
C429 B.n286 VSUBS 0.017313f
C430 B.n287 VSUBS 0.016666f
C431 B.n288 VSUBS 0.016666f
C432 B.n289 VSUBS 0.006756f
C433 B.n290 VSUBS 0.006756f
C434 B.n291 VSUBS 0.006756f
C435 B.n292 VSUBS 0.006756f
C436 B.n293 VSUBS 0.006756f
C437 B.n294 VSUBS 0.006756f
C438 B.n295 VSUBS 0.006756f
C439 B.n296 VSUBS 0.006756f
C440 B.n297 VSUBS 0.006756f
C441 B.n298 VSUBS 0.006756f
C442 B.n299 VSUBS 0.006756f
C443 B.n300 VSUBS 0.006756f
C444 B.n301 VSUBS 0.006756f
C445 B.n302 VSUBS 0.006756f
C446 B.n303 VSUBS 0.006756f
C447 B.n304 VSUBS 0.006756f
C448 B.n305 VSUBS 0.006756f
C449 B.n306 VSUBS 0.006756f
C450 B.n307 VSUBS 0.006756f
C451 B.n308 VSUBS 0.006756f
C452 B.n309 VSUBS 0.006756f
C453 B.n310 VSUBS 0.006756f
C454 B.n311 VSUBS 0.006756f
C455 B.n312 VSUBS 0.006756f
C456 B.n313 VSUBS 0.006756f
C457 B.n314 VSUBS 0.006756f
C458 B.n315 VSUBS 0.006756f
C459 B.n316 VSUBS 0.006756f
C460 B.n317 VSUBS 0.006756f
C461 B.n318 VSUBS 0.006756f
C462 B.n319 VSUBS 0.006756f
C463 B.n320 VSUBS 0.006756f
C464 B.n321 VSUBS 0.006756f
C465 B.n322 VSUBS 0.006756f
C466 B.n323 VSUBS 0.006756f
C467 B.n324 VSUBS 0.006756f
C468 B.n325 VSUBS 0.006756f
C469 B.n326 VSUBS 0.006756f
C470 B.n327 VSUBS 0.006756f
C471 B.n328 VSUBS 0.006756f
C472 B.n329 VSUBS 0.006756f
C473 B.n330 VSUBS 0.006756f
C474 B.n331 VSUBS 0.006756f
C475 B.n332 VSUBS 0.006756f
C476 B.n333 VSUBS 0.006756f
C477 B.n334 VSUBS 0.006756f
C478 B.n335 VSUBS 0.006756f
C479 B.n336 VSUBS 0.006756f
C480 B.n337 VSUBS 0.006756f
C481 B.n338 VSUBS 0.006756f
C482 B.n339 VSUBS 0.006756f
C483 B.n340 VSUBS 0.006756f
C484 B.n341 VSUBS 0.006756f
C485 B.n342 VSUBS 0.006756f
C486 B.n343 VSUBS 0.006756f
C487 B.n344 VSUBS 0.006756f
C488 B.n345 VSUBS 0.006756f
C489 B.n346 VSUBS 0.006756f
C490 B.n347 VSUBS 0.006756f
C491 B.n348 VSUBS 0.006756f
C492 B.n349 VSUBS 0.006756f
C493 B.n350 VSUBS 0.006756f
C494 B.n351 VSUBS 0.006756f
C495 B.n352 VSUBS 0.006756f
C496 B.n353 VSUBS 0.006756f
C497 B.n354 VSUBS 0.006756f
C498 B.n355 VSUBS 0.006756f
C499 B.n356 VSUBS 0.006756f
C500 B.n357 VSUBS 0.006756f
C501 B.n358 VSUBS 0.006756f
C502 B.n359 VSUBS 0.017383f
C503 B.n360 VSUBS 0.016666f
C504 B.n361 VSUBS 0.017313f
C505 B.n362 VSUBS 0.006756f
C506 B.n363 VSUBS 0.006756f
C507 B.n364 VSUBS 0.006756f
C508 B.n365 VSUBS 0.006756f
C509 B.n366 VSUBS 0.006756f
C510 B.n367 VSUBS 0.006756f
C511 B.n368 VSUBS 0.006756f
C512 B.n369 VSUBS 0.006756f
C513 B.n370 VSUBS 0.006756f
C514 B.n371 VSUBS 0.006756f
C515 B.n372 VSUBS 0.006756f
C516 B.n373 VSUBS 0.006756f
C517 B.n374 VSUBS 0.006756f
C518 B.n375 VSUBS 0.006756f
C519 B.n376 VSUBS 0.006756f
C520 B.n377 VSUBS 0.006756f
C521 B.n378 VSUBS 0.006756f
C522 B.n379 VSUBS 0.006756f
C523 B.n380 VSUBS 0.006756f
C524 B.n381 VSUBS 0.006756f
C525 B.n382 VSUBS 0.006756f
C526 B.n383 VSUBS 0.006756f
C527 B.n384 VSUBS 0.006756f
C528 B.n385 VSUBS 0.006756f
C529 B.n386 VSUBS 0.006756f
C530 B.n387 VSUBS 0.006756f
C531 B.n388 VSUBS 0.006756f
C532 B.n389 VSUBS 0.006756f
C533 B.n390 VSUBS 0.006756f
C534 B.n391 VSUBS 0.006756f
C535 B.n392 VSUBS 0.006756f
C536 B.n393 VSUBS 0.006756f
C537 B.n394 VSUBS 0.006756f
C538 B.n395 VSUBS 0.006756f
C539 B.n396 VSUBS 0.006756f
C540 B.n397 VSUBS 0.006756f
C541 B.n398 VSUBS 0.006756f
C542 B.n399 VSUBS 0.006756f
C543 B.n400 VSUBS 0.006756f
C544 B.n401 VSUBS 0.006756f
C545 B.n402 VSUBS 0.006756f
C546 B.n403 VSUBS 0.006756f
C547 B.n404 VSUBS 0.006756f
C548 B.n405 VSUBS 0.006756f
C549 B.n406 VSUBS 0.006756f
C550 B.n407 VSUBS 0.006756f
C551 B.n408 VSUBS 0.006756f
C552 B.n409 VSUBS 0.006756f
C553 B.n410 VSUBS 0.006756f
C554 B.n411 VSUBS 0.00467f
C555 B.n412 VSUBS 0.015653f
C556 B.n413 VSUBS 0.005464f
C557 B.n414 VSUBS 0.006756f
C558 B.n415 VSUBS 0.006756f
C559 B.n416 VSUBS 0.006756f
C560 B.n417 VSUBS 0.006756f
C561 B.n418 VSUBS 0.006756f
C562 B.n419 VSUBS 0.006756f
C563 B.n420 VSUBS 0.006756f
C564 B.n421 VSUBS 0.006756f
C565 B.n422 VSUBS 0.006756f
C566 B.n423 VSUBS 0.006756f
C567 B.n424 VSUBS 0.006756f
C568 B.n425 VSUBS 0.005464f
C569 B.n426 VSUBS 0.015653f
C570 B.n427 VSUBS 0.00467f
C571 B.n428 VSUBS 0.006756f
C572 B.n429 VSUBS 0.006756f
C573 B.n430 VSUBS 0.006756f
C574 B.n431 VSUBS 0.006756f
C575 B.n432 VSUBS 0.006756f
C576 B.n433 VSUBS 0.006756f
C577 B.n434 VSUBS 0.006756f
C578 B.n435 VSUBS 0.006756f
C579 B.n436 VSUBS 0.006756f
C580 B.n437 VSUBS 0.006756f
C581 B.n438 VSUBS 0.006756f
C582 B.n439 VSUBS 0.006756f
C583 B.n440 VSUBS 0.006756f
C584 B.n441 VSUBS 0.006756f
C585 B.n442 VSUBS 0.006756f
C586 B.n443 VSUBS 0.006756f
C587 B.n444 VSUBS 0.006756f
C588 B.n445 VSUBS 0.006756f
C589 B.n446 VSUBS 0.006756f
C590 B.n447 VSUBS 0.006756f
C591 B.n448 VSUBS 0.006756f
C592 B.n449 VSUBS 0.006756f
C593 B.n450 VSUBS 0.006756f
C594 B.n451 VSUBS 0.006756f
C595 B.n452 VSUBS 0.006756f
C596 B.n453 VSUBS 0.006756f
C597 B.n454 VSUBS 0.006756f
C598 B.n455 VSUBS 0.006756f
C599 B.n456 VSUBS 0.006756f
C600 B.n457 VSUBS 0.006756f
C601 B.n458 VSUBS 0.006756f
C602 B.n459 VSUBS 0.006756f
C603 B.n460 VSUBS 0.006756f
C604 B.n461 VSUBS 0.006756f
C605 B.n462 VSUBS 0.006756f
C606 B.n463 VSUBS 0.006756f
C607 B.n464 VSUBS 0.006756f
C608 B.n465 VSUBS 0.006756f
C609 B.n466 VSUBS 0.006756f
C610 B.n467 VSUBS 0.006756f
C611 B.n468 VSUBS 0.006756f
C612 B.n469 VSUBS 0.006756f
C613 B.n470 VSUBS 0.006756f
C614 B.n471 VSUBS 0.006756f
C615 B.n472 VSUBS 0.006756f
C616 B.n473 VSUBS 0.006756f
C617 B.n474 VSUBS 0.006756f
C618 B.n475 VSUBS 0.006756f
C619 B.n476 VSUBS 0.006756f
C620 B.n477 VSUBS 0.017313f
C621 B.n478 VSUBS 0.016666f
C622 B.n479 VSUBS 0.016666f
C623 B.n480 VSUBS 0.006756f
C624 B.n481 VSUBS 0.006756f
C625 B.n482 VSUBS 0.006756f
C626 B.n483 VSUBS 0.006756f
C627 B.n484 VSUBS 0.006756f
C628 B.n485 VSUBS 0.006756f
C629 B.n486 VSUBS 0.006756f
C630 B.n487 VSUBS 0.006756f
C631 B.n488 VSUBS 0.006756f
C632 B.n489 VSUBS 0.006756f
C633 B.n490 VSUBS 0.006756f
C634 B.n491 VSUBS 0.006756f
C635 B.n492 VSUBS 0.006756f
C636 B.n493 VSUBS 0.006756f
C637 B.n494 VSUBS 0.006756f
C638 B.n495 VSUBS 0.006756f
C639 B.n496 VSUBS 0.006756f
C640 B.n497 VSUBS 0.006756f
C641 B.n498 VSUBS 0.006756f
C642 B.n499 VSUBS 0.006756f
C643 B.n500 VSUBS 0.006756f
C644 B.n501 VSUBS 0.006756f
C645 B.n502 VSUBS 0.006756f
C646 B.n503 VSUBS 0.006756f
C647 B.n504 VSUBS 0.006756f
C648 B.n505 VSUBS 0.006756f
C649 B.n506 VSUBS 0.006756f
C650 B.n507 VSUBS 0.006756f
C651 B.n508 VSUBS 0.006756f
C652 B.n509 VSUBS 0.006756f
C653 B.n510 VSUBS 0.006756f
C654 B.n511 VSUBS 0.006756f
C655 B.n512 VSUBS 0.006756f
C656 B.n513 VSUBS 0.006756f
C657 B.n514 VSUBS 0.006756f
C658 B.n515 VSUBS 0.015298f
C659 VDD1.n0 VSUBS 0.022338f
C660 VDD1.n1 VSUBS 0.020566f
C661 VDD1.n2 VSUBS 0.011051f
C662 VDD1.n3 VSUBS 0.026121f
C663 VDD1.n4 VSUBS 0.011376f
C664 VDD1.n5 VSUBS 0.020566f
C665 VDD1.n6 VSUBS 0.011376f
C666 VDD1.n7 VSUBS 0.011051f
C667 VDD1.n8 VSUBS 0.026121f
C668 VDD1.n9 VSUBS 0.026121f
C669 VDD1.n10 VSUBS 0.011702f
C670 VDD1.n11 VSUBS 0.020566f
C671 VDD1.n12 VSUBS 0.011051f
C672 VDD1.n13 VSUBS 0.026121f
C673 VDD1.n14 VSUBS 0.011702f
C674 VDD1.n15 VSUBS 0.77432f
C675 VDD1.n16 VSUBS 0.011051f
C676 VDD1.t1 VSUBS 0.056142f
C677 VDD1.n17 VSUBS 0.137637f
C678 VDD1.n18 VSUBS 0.01965f
C679 VDD1.n19 VSUBS 0.019591f
C680 VDD1.n20 VSUBS 0.026121f
C681 VDD1.n21 VSUBS 0.011702f
C682 VDD1.n22 VSUBS 0.011051f
C683 VDD1.n23 VSUBS 0.020566f
C684 VDD1.n24 VSUBS 0.020566f
C685 VDD1.n25 VSUBS 0.011051f
C686 VDD1.n26 VSUBS 0.011702f
C687 VDD1.n27 VSUBS 0.026121f
C688 VDD1.n28 VSUBS 0.026121f
C689 VDD1.n29 VSUBS 0.011702f
C690 VDD1.n30 VSUBS 0.011051f
C691 VDD1.n31 VSUBS 0.020566f
C692 VDD1.n32 VSUBS 0.020566f
C693 VDD1.n33 VSUBS 0.011051f
C694 VDD1.n34 VSUBS 0.011702f
C695 VDD1.n35 VSUBS 0.026121f
C696 VDD1.n36 VSUBS 0.026121f
C697 VDD1.n37 VSUBS 0.011702f
C698 VDD1.n38 VSUBS 0.011051f
C699 VDD1.n39 VSUBS 0.020566f
C700 VDD1.n40 VSUBS 0.020566f
C701 VDD1.n41 VSUBS 0.011051f
C702 VDD1.n42 VSUBS 0.011702f
C703 VDD1.n43 VSUBS 0.026121f
C704 VDD1.n44 VSUBS 0.06235f
C705 VDD1.n45 VSUBS 0.011702f
C706 VDD1.n46 VSUBS 0.011051f
C707 VDD1.n47 VSUBS 0.051471f
C708 VDD1.n48 VSUBS 0.046653f
C709 VDD1.n49 VSUBS 0.022338f
C710 VDD1.n50 VSUBS 0.020566f
C711 VDD1.n51 VSUBS 0.011051f
C712 VDD1.n52 VSUBS 0.026121f
C713 VDD1.n53 VSUBS 0.011376f
C714 VDD1.n54 VSUBS 0.020566f
C715 VDD1.n55 VSUBS 0.011702f
C716 VDD1.n56 VSUBS 0.026121f
C717 VDD1.n57 VSUBS 0.011702f
C718 VDD1.n58 VSUBS 0.020566f
C719 VDD1.n59 VSUBS 0.011051f
C720 VDD1.n60 VSUBS 0.026121f
C721 VDD1.n61 VSUBS 0.011702f
C722 VDD1.n62 VSUBS 0.77432f
C723 VDD1.n63 VSUBS 0.011051f
C724 VDD1.t0 VSUBS 0.056142f
C725 VDD1.n64 VSUBS 0.137637f
C726 VDD1.n65 VSUBS 0.01965f
C727 VDD1.n66 VSUBS 0.019591f
C728 VDD1.n67 VSUBS 0.026121f
C729 VDD1.n68 VSUBS 0.011702f
C730 VDD1.n69 VSUBS 0.011051f
C731 VDD1.n70 VSUBS 0.020566f
C732 VDD1.n71 VSUBS 0.020566f
C733 VDD1.n72 VSUBS 0.011051f
C734 VDD1.n73 VSUBS 0.011702f
C735 VDD1.n74 VSUBS 0.026121f
C736 VDD1.n75 VSUBS 0.026121f
C737 VDD1.n76 VSUBS 0.011702f
C738 VDD1.n77 VSUBS 0.011051f
C739 VDD1.n78 VSUBS 0.020566f
C740 VDD1.n79 VSUBS 0.020566f
C741 VDD1.n80 VSUBS 0.011051f
C742 VDD1.n81 VSUBS 0.011051f
C743 VDD1.n82 VSUBS 0.011702f
C744 VDD1.n83 VSUBS 0.026121f
C745 VDD1.n84 VSUBS 0.026121f
C746 VDD1.n85 VSUBS 0.026121f
C747 VDD1.n86 VSUBS 0.011376f
C748 VDD1.n87 VSUBS 0.011051f
C749 VDD1.n88 VSUBS 0.020566f
C750 VDD1.n89 VSUBS 0.020566f
C751 VDD1.n90 VSUBS 0.011051f
C752 VDD1.n91 VSUBS 0.011702f
C753 VDD1.n92 VSUBS 0.026121f
C754 VDD1.n93 VSUBS 0.06235f
C755 VDD1.n94 VSUBS 0.011702f
C756 VDD1.n95 VSUBS 0.011051f
C757 VDD1.n96 VSUBS 0.051471f
C758 VDD1.n97 VSUBS 0.542127f
C759 VTAIL.n0 VSUBS 0.025825f
C760 VTAIL.n1 VSUBS 0.023777f
C761 VTAIL.n2 VSUBS 0.012777f
C762 VTAIL.n3 VSUBS 0.0302f
C763 VTAIL.n4 VSUBS 0.013153f
C764 VTAIL.n5 VSUBS 0.023777f
C765 VTAIL.n6 VSUBS 0.013528f
C766 VTAIL.n7 VSUBS 0.0302f
C767 VTAIL.n8 VSUBS 0.013528f
C768 VTAIL.n9 VSUBS 0.023777f
C769 VTAIL.n10 VSUBS 0.012777f
C770 VTAIL.n11 VSUBS 0.0302f
C771 VTAIL.n12 VSUBS 0.013528f
C772 VTAIL.n13 VSUBS 0.89522f
C773 VTAIL.n14 VSUBS 0.012777f
C774 VTAIL.t2 VSUBS 0.064907f
C775 VTAIL.n15 VSUBS 0.159127f
C776 VTAIL.n16 VSUBS 0.022718f
C777 VTAIL.n17 VSUBS 0.02265f
C778 VTAIL.n18 VSUBS 0.0302f
C779 VTAIL.n19 VSUBS 0.013528f
C780 VTAIL.n20 VSUBS 0.012777f
C781 VTAIL.n21 VSUBS 0.023777f
C782 VTAIL.n22 VSUBS 0.023777f
C783 VTAIL.n23 VSUBS 0.012777f
C784 VTAIL.n24 VSUBS 0.013528f
C785 VTAIL.n25 VSUBS 0.0302f
C786 VTAIL.n26 VSUBS 0.0302f
C787 VTAIL.n27 VSUBS 0.013528f
C788 VTAIL.n28 VSUBS 0.012777f
C789 VTAIL.n29 VSUBS 0.023777f
C790 VTAIL.n30 VSUBS 0.023777f
C791 VTAIL.n31 VSUBS 0.012777f
C792 VTAIL.n32 VSUBS 0.012777f
C793 VTAIL.n33 VSUBS 0.013528f
C794 VTAIL.n34 VSUBS 0.0302f
C795 VTAIL.n35 VSUBS 0.0302f
C796 VTAIL.n36 VSUBS 0.0302f
C797 VTAIL.n37 VSUBS 0.013153f
C798 VTAIL.n38 VSUBS 0.012777f
C799 VTAIL.n39 VSUBS 0.023777f
C800 VTAIL.n40 VSUBS 0.023777f
C801 VTAIL.n41 VSUBS 0.012777f
C802 VTAIL.n42 VSUBS 0.013528f
C803 VTAIL.n43 VSUBS 0.0302f
C804 VTAIL.n44 VSUBS 0.072085f
C805 VTAIL.n45 VSUBS 0.013528f
C806 VTAIL.n46 VSUBS 0.012777f
C807 VTAIL.n47 VSUBS 0.059508f
C808 VTAIL.n48 VSUBS 0.036341f
C809 VTAIL.n49 VSUBS 1.41155f
C810 VTAIL.n50 VSUBS 0.025825f
C811 VTAIL.n51 VSUBS 0.023777f
C812 VTAIL.n52 VSUBS 0.012777f
C813 VTAIL.n53 VSUBS 0.0302f
C814 VTAIL.n54 VSUBS 0.013153f
C815 VTAIL.n55 VSUBS 0.023777f
C816 VTAIL.n56 VSUBS 0.013153f
C817 VTAIL.n57 VSUBS 0.012777f
C818 VTAIL.n58 VSUBS 0.0302f
C819 VTAIL.n59 VSUBS 0.0302f
C820 VTAIL.n60 VSUBS 0.013528f
C821 VTAIL.n61 VSUBS 0.023777f
C822 VTAIL.n62 VSUBS 0.012777f
C823 VTAIL.n63 VSUBS 0.0302f
C824 VTAIL.n64 VSUBS 0.013528f
C825 VTAIL.n65 VSUBS 0.89522f
C826 VTAIL.n66 VSUBS 0.012777f
C827 VTAIL.t0 VSUBS 0.064907f
C828 VTAIL.n67 VSUBS 0.159127f
C829 VTAIL.n68 VSUBS 0.022718f
C830 VTAIL.n69 VSUBS 0.02265f
C831 VTAIL.n70 VSUBS 0.0302f
C832 VTAIL.n71 VSUBS 0.013528f
C833 VTAIL.n72 VSUBS 0.012777f
C834 VTAIL.n73 VSUBS 0.023777f
C835 VTAIL.n74 VSUBS 0.023777f
C836 VTAIL.n75 VSUBS 0.012777f
C837 VTAIL.n76 VSUBS 0.013528f
C838 VTAIL.n77 VSUBS 0.0302f
C839 VTAIL.n78 VSUBS 0.0302f
C840 VTAIL.n79 VSUBS 0.013528f
C841 VTAIL.n80 VSUBS 0.012777f
C842 VTAIL.n81 VSUBS 0.023777f
C843 VTAIL.n82 VSUBS 0.023777f
C844 VTAIL.n83 VSUBS 0.012777f
C845 VTAIL.n84 VSUBS 0.013528f
C846 VTAIL.n85 VSUBS 0.0302f
C847 VTAIL.n86 VSUBS 0.0302f
C848 VTAIL.n87 VSUBS 0.013528f
C849 VTAIL.n88 VSUBS 0.012777f
C850 VTAIL.n89 VSUBS 0.023777f
C851 VTAIL.n90 VSUBS 0.023777f
C852 VTAIL.n91 VSUBS 0.012777f
C853 VTAIL.n92 VSUBS 0.013528f
C854 VTAIL.n93 VSUBS 0.0302f
C855 VTAIL.n94 VSUBS 0.072085f
C856 VTAIL.n95 VSUBS 0.013528f
C857 VTAIL.n96 VSUBS 0.012777f
C858 VTAIL.n97 VSUBS 0.059508f
C859 VTAIL.n98 VSUBS 0.036341f
C860 VTAIL.n99 VSUBS 1.45217f
C861 VTAIL.n100 VSUBS 0.025825f
C862 VTAIL.n101 VSUBS 0.023777f
C863 VTAIL.n102 VSUBS 0.012777f
C864 VTAIL.n103 VSUBS 0.0302f
C865 VTAIL.n104 VSUBS 0.013153f
C866 VTAIL.n105 VSUBS 0.023777f
C867 VTAIL.n106 VSUBS 0.013153f
C868 VTAIL.n107 VSUBS 0.012777f
C869 VTAIL.n108 VSUBS 0.0302f
C870 VTAIL.n109 VSUBS 0.0302f
C871 VTAIL.n110 VSUBS 0.013528f
C872 VTAIL.n111 VSUBS 0.023777f
C873 VTAIL.n112 VSUBS 0.012777f
C874 VTAIL.n113 VSUBS 0.0302f
C875 VTAIL.n114 VSUBS 0.013528f
C876 VTAIL.n115 VSUBS 0.89522f
C877 VTAIL.n116 VSUBS 0.012777f
C878 VTAIL.t1 VSUBS 0.064907f
C879 VTAIL.n117 VSUBS 0.159127f
C880 VTAIL.n118 VSUBS 0.022718f
C881 VTAIL.n119 VSUBS 0.02265f
C882 VTAIL.n120 VSUBS 0.0302f
C883 VTAIL.n121 VSUBS 0.013528f
C884 VTAIL.n122 VSUBS 0.012777f
C885 VTAIL.n123 VSUBS 0.023777f
C886 VTAIL.n124 VSUBS 0.023777f
C887 VTAIL.n125 VSUBS 0.012777f
C888 VTAIL.n126 VSUBS 0.013528f
C889 VTAIL.n127 VSUBS 0.0302f
C890 VTAIL.n128 VSUBS 0.0302f
C891 VTAIL.n129 VSUBS 0.013528f
C892 VTAIL.n130 VSUBS 0.012777f
C893 VTAIL.n131 VSUBS 0.023777f
C894 VTAIL.n132 VSUBS 0.023777f
C895 VTAIL.n133 VSUBS 0.012777f
C896 VTAIL.n134 VSUBS 0.013528f
C897 VTAIL.n135 VSUBS 0.0302f
C898 VTAIL.n136 VSUBS 0.0302f
C899 VTAIL.n137 VSUBS 0.013528f
C900 VTAIL.n138 VSUBS 0.012777f
C901 VTAIL.n139 VSUBS 0.023777f
C902 VTAIL.n140 VSUBS 0.023777f
C903 VTAIL.n141 VSUBS 0.012777f
C904 VTAIL.n142 VSUBS 0.013528f
C905 VTAIL.n143 VSUBS 0.0302f
C906 VTAIL.n144 VSUBS 0.072085f
C907 VTAIL.n145 VSUBS 0.013528f
C908 VTAIL.n146 VSUBS 0.012777f
C909 VTAIL.n147 VSUBS 0.059508f
C910 VTAIL.n148 VSUBS 0.036341f
C911 VTAIL.n149 VSUBS 1.27186f
C912 VTAIL.n150 VSUBS 0.025825f
C913 VTAIL.n151 VSUBS 0.023777f
C914 VTAIL.n152 VSUBS 0.012777f
C915 VTAIL.n153 VSUBS 0.0302f
C916 VTAIL.n154 VSUBS 0.013153f
C917 VTAIL.n155 VSUBS 0.023777f
C918 VTAIL.n156 VSUBS 0.013528f
C919 VTAIL.n157 VSUBS 0.0302f
C920 VTAIL.n158 VSUBS 0.013528f
C921 VTAIL.n159 VSUBS 0.023777f
C922 VTAIL.n160 VSUBS 0.012777f
C923 VTAIL.n161 VSUBS 0.0302f
C924 VTAIL.n162 VSUBS 0.013528f
C925 VTAIL.n163 VSUBS 0.89522f
C926 VTAIL.n164 VSUBS 0.012777f
C927 VTAIL.t3 VSUBS 0.064907f
C928 VTAIL.n165 VSUBS 0.159127f
C929 VTAIL.n166 VSUBS 0.022718f
C930 VTAIL.n167 VSUBS 0.02265f
C931 VTAIL.n168 VSUBS 0.0302f
C932 VTAIL.n169 VSUBS 0.013528f
C933 VTAIL.n170 VSUBS 0.012777f
C934 VTAIL.n171 VSUBS 0.023777f
C935 VTAIL.n172 VSUBS 0.023777f
C936 VTAIL.n173 VSUBS 0.012777f
C937 VTAIL.n174 VSUBS 0.013528f
C938 VTAIL.n175 VSUBS 0.0302f
C939 VTAIL.n176 VSUBS 0.0302f
C940 VTAIL.n177 VSUBS 0.013528f
C941 VTAIL.n178 VSUBS 0.012777f
C942 VTAIL.n179 VSUBS 0.023777f
C943 VTAIL.n180 VSUBS 0.023777f
C944 VTAIL.n181 VSUBS 0.012777f
C945 VTAIL.n182 VSUBS 0.012777f
C946 VTAIL.n183 VSUBS 0.013528f
C947 VTAIL.n184 VSUBS 0.0302f
C948 VTAIL.n185 VSUBS 0.0302f
C949 VTAIL.n186 VSUBS 0.0302f
C950 VTAIL.n187 VSUBS 0.013153f
C951 VTAIL.n188 VSUBS 0.012777f
C952 VTAIL.n189 VSUBS 0.023777f
C953 VTAIL.n190 VSUBS 0.023777f
C954 VTAIL.n191 VSUBS 0.012777f
C955 VTAIL.n192 VSUBS 0.013528f
C956 VTAIL.n193 VSUBS 0.0302f
C957 VTAIL.n194 VSUBS 0.072085f
C958 VTAIL.n195 VSUBS 0.013528f
C959 VTAIL.n196 VSUBS 0.012777f
C960 VTAIL.n197 VSUBS 0.059508f
C961 VTAIL.n198 VSUBS 0.036341f
C962 VTAIL.n199 VSUBS 1.18633f
C963 VP.t0 VSUBS 3.24575f
C964 VP.t1 VSUBS 2.69057f
C965 VP.n0 VSUBS 4.27933f
.ends

