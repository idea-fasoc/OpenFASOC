* NGSPICE file created from diff_pair_sample_1777.ext - technology: sky130A

.subckt diff_pair_sample_1777 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.46
X1 B.t11 B.t9 B.t10 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.46
X2 B.t8 B.t6 B.t7 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.46
X3 VTAIL.t2 VN.t0 VDD2.t7 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.46
X4 VDD1.t6 VP.t1 VTAIL.t14 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X5 B.t5 B.t3 B.t4 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.46
X6 VDD2.t6 VN.t1 VTAIL.t3 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.46
X7 VDD2.t5 VN.t2 VTAIL.t5 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.46
X8 VTAIL.t6 VN.t3 VDD2.t4 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X9 VDD2.t3 VN.t4 VTAIL.t0 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X10 VTAIL.t7 VN.t5 VDD2.t2 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X11 B.t2 B.t0 B.t1 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0 ps=0 w=4.89 l=3.46
X12 VTAIL.t13 VP.t2 VDD1.t5 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X13 VDD1.t1 VP.t3 VTAIL.t12 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X14 VTAIL.t11 VP.t4 VDD1.t0 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X15 VTAIL.t10 VP.t5 VDD1.t3 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.46
X16 VDD1.t4 VP.t6 VTAIL.t9 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.46
X17 VDD2.t1 VN.t6 VTAIL.t1 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=0.80685 ps=5.22 w=4.89 l=3.46
X18 VTAIL.t4 VN.t7 VDD2.t0 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=1.9071 pd=10.56 as=0.80685 ps=5.22 w=4.89 l=3.46
X19 VDD1.t2 VP.t7 VTAIL.t8 w_n4760_n1946# sky130_fd_pr__pfet_01v8 ad=0.80685 pd=5.22 as=1.9071 ps=10.56 w=4.89 l=3.46
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n17 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n85 VP.n84 161.3
R16 VP.n83 VP.n1 161.3
R17 VP.n82 VP.n81 161.3
R18 VP.n80 VP.n2 161.3
R19 VP.n79 VP.n78 161.3
R20 VP.n77 VP.n3 161.3
R21 VP.n76 VP.n75 161.3
R22 VP.n74 VP.n4 161.3
R23 VP.n73 VP.n72 161.3
R24 VP.n70 VP.n5 161.3
R25 VP.n69 VP.n68 161.3
R26 VP.n67 VP.n6 161.3
R27 VP.n66 VP.n65 161.3
R28 VP.n64 VP.n7 161.3
R29 VP.n63 VP.n62 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n59 VP.n9 161.3
R32 VP.n58 VP.n57 161.3
R33 VP.n56 VP.n10 161.3
R34 VP.n55 VP.n54 161.3
R35 VP.n53 VP.n11 161.3
R36 VP.n52 VP.n51 161.3
R37 VP.n50 VP.n12 161.3
R38 VP.n49 VP.n48 81.0146
R39 VP.n86 VP.n0 81.0146
R40 VP.n47 VP.n13 81.0146
R41 VP.n22 VP.t5 67.3011
R42 VP.n54 VP.n10 56.5193
R43 VP.n78 VP.n2 56.5193
R44 VP.n39 VP.n15 56.5193
R45 VP.n22 VP.n21 55.2448
R46 VP.n49 VP.n47 49.5978
R47 VP.n65 VP.n6 40.4934
R48 VP.n69 VP.n6 40.4934
R49 VP.n30 VP.n19 40.4934
R50 VP.n26 VP.n19 40.4934
R51 VP.n48 VP.t0 34.0609
R52 VP.n8 VP.t1 34.0609
R53 VP.n71 VP.t2 34.0609
R54 VP.n0 VP.t7 34.0609
R55 VP.n13 VP.t6 34.0609
R56 VP.n32 VP.t4 34.0609
R57 VP.n21 VP.t3 34.0609
R58 VP.n52 VP.n12 24.4675
R59 VP.n53 VP.n52 24.4675
R60 VP.n54 VP.n53 24.4675
R61 VP.n58 VP.n10 24.4675
R62 VP.n59 VP.n58 24.4675
R63 VP.n60 VP.n59 24.4675
R64 VP.n64 VP.n63 24.4675
R65 VP.n65 VP.n64 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n72 VP.n70 24.4675
R68 VP.n76 VP.n4 24.4675
R69 VP.n77 VP.n76 24.4675
R70 VP.n78 VP.n77 24.4675
R71 VP.n82 VP.n2 24.4675
R72 VP.n83 VP.n82 24.4675
R73 VP.n84 VP.n83 24.4675
R74 VP.n43 VP.n15 24.4675
R75 VP.n44 VP.n43 24.4675
R76 VP.n45 VP.n44 24.4675
R77 VP.n31 VP.n30 24.4675
R78 VP.n33 VP.n31 24.4675
R79 VP.n37 VP.n17 24.4675
R80 VP.n38 VP.n37 24.4675
R81 VP.n39 VP.n38 24.4675
R82 VP.n25 VP.n24 24.4675
R83 VP.n26 VP.n25 24.4675
R84 VP.n63 VP.n8 19.3294
R85 VP.n72 VP.n71 19.3294
R86 VP.n33 VP.n32 19.3294
R87 VP.n24 VP.n21 19.3294
R88 VP.n48 VP.n12 9.05329
R89 VP.n84 VP.n0 9.05329
R90 VP.n45 VP.n13 9.05329
R91 VP.n60 VP.n8 5.13857
R92 VP.n71 VP.n4 5.13857
R93 VP.n32 VP.n17 5.13857
R94 VP.n23 VP.n22 3.18789
R95 VP.n47 VP.n46 0.354971
R96 VP.n50 VP.n49 0.354971
R97 VP.n86 VP.n85 0.354971
R98 VP VP.n86 0.26696
R99 VP.n23 VP.n20 0.189894
R100 VP.n27 VP.n20 0.189894
R101 VP.n28 VP.n27 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n29 VP.n18 0.189894
R104 VP.n34 VP.n18 0.189894
R105 VP.n35 VP.n34 0.189894
R106 VP.n36 VP.n35 0.189894
R107 VP.n36 VP.n16 0.189894
R108 VP.n40 VP.n16 0.189894
R109 VP.n41 VP.n40 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n42 VP.n14 0.189894
R112 VP.n46 VP.n14 0.189894
R113 VP.n51 VP.n50 0.189894
R114 VP.n51 VP.n11 0.189894
R115 VP.n55 VP.n11 0.189894
R116 VP.n56 VP.n55 0.189894
R117 VP.n57 VP.n56 0.189894
R118 VP.n57 VP.n9 0.189894
R119 VP.n61 VP.n9 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n62 VP.n7 0.189894
R122 VP.n66 VP.n7 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n68 VP.n5 0.189894
R126 VP.n73 VP.n5 0.189894
R127 VP.n74 VP.n73 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n75 VP.n3 0.189894
R130 VP.n79 VP.n3 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n81 VP.n1 0.189894
R134 VP.n85 VP.n1 0.189894
R135 VDD1 VDD1.n0 101.55
R136 VDD1.n3 VDD1.n2 101.438
R137 VDD1.n3 VDD1.n1 101.438
R138 VDD1.n5 VDD1.n4 99.8588
R139 VDD1.n5 VDD1.n3 43.2164
R140 VDD1.n4 VDD1.t0 6.64774
R141 VDD1.n4 VDD1.t4 6.64774
R142 VDD1.n0 VDD1.t3 6.64774
R143 VDD1.n0 VDD1.t1 6.64774
R144 VDD1.n2 VDD1.t5 6.64774
R145 VDD1.n2 VDD1.t2 6.64774
R146 VDD1.n1 VDD1.t7 6.64774
R147 VDD1.n1 VDD1.t6 6.64774
R148 VDD1 VDD1.n5 1.57593
R149 VTAIL.n11 VTAIL.t10 89.8274
R150 VTAIL.n10 VTAIL.t5 89.8274
R151 VTAIL.n7 VTAIL.t4 89.8274
R152 VTAIL.n15 VTAIL.t3 89.8273
R153 VTAIL.n2 VTAIL.t2 89.8273
R154 VTAIL.n3 VTAIL.t8 89.8273
R155 VTAIL.n6 VTAIL.t15 89.8273
R156 VTAIL.n14 VTAIL.t9 89.8273
R157 VTAIL.n13 VTAIL.n12 83.1802
R158 VTAIL.n9 VTAIL.n8 83.1802
R159 VTAIL.n1 VTAIL.n0 83.18
R160 VTAIL.n5 VTAIL.n4 83.18
R161 VTAIL.n15 VTAIL.n14 19.8496
R162 VTAIL.n7 VTAIL.n6 19.8496
R163 VTAIL.n0 VTAIL.t0 6.64774
R164 VTAIL.n0 VTAIL.t6 6.64774
R165 VTAIL.n4 VTAIL.t14 6.64774
R166 VTAIL.n4 VTAIL.t13 6.64774
R167 VTAIL.n12 VTAIL.t12 6.64774
R168 VTAIL.n12 VTAIL.t11 6.64774
R169 VTAIL.n8 VTAIL.t1 6.64774
R170 VTAIL.n8 VTAIL.t7 6.64774
R171 VTAIL.n9 VTAIL.n7 3.26774
R172 VTAIL.n10 VTAIL.n9 3.26774
R173 VTAIL.n13 VTAIL.n11 3.26774
R174 VTAIL.n14 VTAIL.n13 3.26774
R175 VTAIL.n6 VTAIL.n5 3.26774
R176 VTAIL.n5 VTAIL.n3 3.26774
R177 VTAIL.n2 VTAIL.n1 3.26774
R178 VTAIL VTAIL.n15 3.20955
R179 VTAIL.n11 VTAIL.n10 0.470328
R180 VTAIL.n3 VTAIL.n2 0.470328
R181 VTAIL VTAIL.n1 0.0586897
R182 B.n557 B.n64 585
R183 B.n559 B.n558 585
R184 B.n560 B.n63 585
R185 B.n562 B.n561 585
R186 B.n563 B.n62 585
R187 B.n565 B.n564 585
R188 B.n566 B.n61 585
R189 B.n568 B.n567 585
R190 B.n569 B.n60 585
R191 B.n571 B.n570 585
R192 B.n572 B.n59 585
R193 B.n574 B.n573 585
R194 B.n575 B.n58 585
R195 B.n577 B.n576 585
R196 B.n578 B.n57 585
R197 B.n580 B.n579 585
R198 B.n581 B.n56 585
R199 B.n583 B.n582 585
R200 B.n584 B.n55 585
R201 B.n586 B.n585 585
R202 B.n587 B.n52 585
R203 B.n590 B.n589 585
R204 B.n591 B.n51 585
R205 B.n593 B.n592 585
R206 B.n594 B.n50 585
R207 B.n596 B.n595 585
R208 B.n597 B.n49 585
R209 B.n599 B.n598 585
R210 B.n600 B.n45 585
R211 B.n602 B.n601 585
R212 B.n603 B.n44 585
R213 B.n605 B.n604 585
R214 B.n606 B.n43 585
R215 B.n608 B.n607 585
R216 B.n609 B.n42 585
R217 B.n611 B.n610 585
R218 B.n612 B.n41 585
R219 B.n614 B.n613 585
R220 B.n615 B.n40 585
R221 B.n617 B.n616 585
R222 B.n618 B.n39 585
R223 B.n620 B.n619 585
R224 B.n621 B.n38 585
R225 B.n623 B.n622 585
R226 B.n624 B.n37 585
R227 B.n626 B.n625 585
R228 B.n627 B.n36 585
R229 B.n629 B.n628 585
R230 B.n630 B.n35 585
R231 B.n632 B.n631 585
R232 B.n633 B.n34 585
R233 B.n556 B.n555 585
R234 B.n554 B.n65 585
R235 B.n553 B.n552 585
R236 B.n551 B.n66 585
R237 B.n550 B.n549 585
R238 B.n548 B.n67 585
R239 B.n547 B.n546 585
R240 B.n545 B.n68 585
R241 B.n544 B.n543 585
R242 B.n542 B.n69 585
R243 B.n541 B.n540 585
R244 B.n539 B.n70 585
R245 B.n538 B.n537 585
R246 B.n536 B.n71 585
R247 B.n535 B.n534 585
R248 B.n533 B.n72 585
R249 B.n532 B.n531 585
R250 B.n530 B.n73 585
R251 B.n529 B.n528 585
R252 B.n527 B.n74 585
R253 B.n526 B.n525 585
R254 B.n524 B.n75 585
R255 B.n523 B.n522 585
R256 B.n521 B.n76 585
R257 B.n520 B.n519 585
R258 B.n518 B.n77 585
R259 B.n517 B.n516 585
R260 B.n515 B.n78 585
R261 B.n514 B.n513 585
R262 B.n512 B.n79 585
R263 B.n511 B.n510 585
R264 B.n509 B.n80 585
R265 B.n508 B.n507 585
R266 B.n506 B.n81 585
R267 B.n505 B.n504 585
R268 B.n503 B.n82 585
R269 B.n502 B.n501 585
R270 B.n500 B.n83 585
R271 B.n499 B.n498 585
R272 B.n497 B.n84 585
R273 B.n496 B.n495 585
R274 B.n494 B.n85 585
R275 B.n493 B.n492 585
R276 B.n491 B.n86 585
R277 B.n490 B.n489 585
R278 B.n488 B.n87 585
R279 B.n487 B.n486 585
R280 B.n485 B.n88 585
R281 B.n484 B.n483 585
R282 B.n482 B.n89 585
R283 B.n481 B.n480 585
R284 B.n479 B.n90 585
R285 B.n478 B.n477 585
R286 B.n476 B.n91 585
R287 B.n475 B.n474 585
R288 B.n473 B.n92 585
R289 B.n472 B.n471 585
R290 B.n470 B.n93 585
R291 B.n469 B.n468 585
R292 B.n467 B.n94 585
R293 B.n466 B.n465 585
R294 B.n464 B.n95 585
R295 B.n463 B.n462 585
R296 B.n461 B.n96 585
R297 B.n460 B.n459 585
R298 B.n458 B.n97 585
R299 B.n457 B.n456 585
R300 B.n455 B.n98 585
R301 B.n454 B.n453 585
R302 B.n452 B.n99 585
R303 B.n451 B.n450 585
R304 B.n449 B.n100 585
R305 B.n448 B.n447 585
R306 B.n446 B.n101 585
R307 B.n445 B.n444 585
R308 B.n443 B.n102 585
R309 B.n442 B.n441 585
R310 B.n440 B.n103 585
R311 B.n439 B.n438 585
R312 B.n437 B.n104 585
R313 B.n436 B.n435 585
R314 B.n434 B.n105 585
R315 B.n433 B.n432 585
R316 B.n431 B.n106 585
R317 B.n430 B.n429 585
R318 B.n428 B.n107 585
R319 B.n427 B.n426 585
R320 B.n425 B.n108 585
R321 B.n424 B.n423 585
R322 B.n422 B.n109 585
R323 B.n421 B.n420 585
R324 B.n419 B.n110 585
R325 B.n418 B.n417 585
R326 B.n416 B.n111 585
R327 B.n415 B.n414 585
R328 B.n413 B.n112 585
R329 B.n412 B.n411 585
R330 B.n410 B.n113 585
R331 B.n409 B.n408 585
R332 B.n407 B.n114 585
R333 B.n406 B.n405 585
R334 B.n404 B.n115 585
R335 B.n403 B.n402 585
R336 B.n401 B.n116 585
R337 B.n400 B.n399 585
R338 B.n398 B.n117 585
R339 B.n397 B.n396 585
R340 B.n395 B.n118 585
R341 B.n394 B.n393 585
R342 B.n392 B.n119 585
R343 B.n391 B.n390 585
R344 B.n389 B.n120 585
R345 B.n388 B.n387 585
R346 B.n386 B.n121 585
R347 B.n385 B.n384 585
R348 B.n383 B.n122 585
R349 B.n382 B.n381 585
R350 B.n380 B.n123 585
R351 B.n379 B.n378 585
R352 B.n377 B.n124 585
R353 B.n376 B.n375 585
R354 B.n374 B.n125 585
R355 B.n373 B.n372 585
R356 B.n371 B.n126 585
R357 B.n370 B.n369 585
R358 B.n368 B.n127 585
R359 B.n367 B.n366 585
R360 B.n365 B.n128 585
R361 B.n364 B.n363 585
R362 B.n283 B.n156 585
R363 B.n285 B.n284 585
R364 B.n286 B.n155 585
R365 B.n288 B.n287 585
R366 B.n289 B.n154 585
R367 B.n291 B.n290 585
R368 B.n292 B.n153 585
R369 B.n294 B.n293 585
R370 B.n295 B.n152 585
R371 B.n297 B.n296 585
R372 B.n298 B.n151 585
R373 B.n300 B.n299 585
R374 B.n301 B.n150 585
R375 B.n303 B.n302 585
R376 B.n304 B.n149 585
R377 B.n306 B.n305 585
R378 B.n307 B.n148 585
R379 B.n309 B.n308 585
R380 B.n310 B.n147 585
R381 B.n312 B.n311 585
R382 B.n313 B.n144 585
R383 B.n316 B.n315 585
R384 B.n317 B.n143 585
R385 B.n319 B.n318 585
R386 B.n320 B.n142 585
R387 B.n322 B.n321 585
R388 B.n323 B.n141 585
R389 B.n325 B.n324 585
R390 B.n326 B.n140 585
R391 B.n331 B.n330 585
R392 B.n332 B.n139 585
R393 B.n334 B.n333 585
R394 B.n335 B.n138 585
R395 B.n337 B.n336 585
R396 B.n338 B.n137 585
R397 B.n340 B.n339 585
R398 B.n341 B.n136 585
R399 B.n343 B.n342 585
R400 B.n344 B.n135 585
R401 B.n346 B.n345 585
R402 B.n347 B.n134 585
R403 B.n349 B.n348 585
R404 B.n350 B.n133 585
R405 B.n352 B.n351 585
R406 B.n353 B.n132 585
R407 B.n355 B.n354 585
R408 B.n356 B.n131 585
R409 B.n358 B.n357 585
R410 B.n359 B.n130 585
R411 B.n361 B.n360 585
R412 B.n362 B.n129 585
R413 B.n282 B.n281 585
R414 B.n280 B.n157 585
R415 B.n279 B.n278 585
R416 B.n277 B.n158 585
R417 B.n276 B.n275 585
R418 B.n274 B.n159 585
R419 B.n273 B.n272 585
R420 B.n271 B.n160 585
R421 B.n270 B.n269 585
R422 B.n268 B.n161 585
R423 B.n267 B.n266 585
R424 B.n265 B.n162 585
R425 B.n264 B.n263 585
R426 B.n262 B.n163 585
R427 B.n261 B.n260 585
R428 B.n259 B.n164 585
R429 B.n258 B.n257 585
R430 B.n256 B.n165 585
R431 B.n255 B.n254 585
R432 B.n253 B.n166 585
R433 B.n252 B.n251 585
R434 B.n250 B.n167 585
R435 B.n249 B.n248 585
R436 B.n247 B.n168 585
R437 B.n246 B.n245 585
R438 B.n244 B.n169 585
R439 B.n243 B.n242 585
R440 B.n241 B.n170 585
R441 B.n240 B.n239 585
R442 B.n238 B.n171 585
R443 B.n237 B.n236 585
R444 B.n235 B.n172 585
R445 B.n234 B.n233 585
R446 B.n232 B.n173 585
R447 B.n231 B.n230 585
R448 B.n229 B.n174 585
R449 B.n228 B.n227 585
R450 B.n226 B.n175 585
R451 B.n225 B.n224 585
R452 B.n223 B.n176 585
R453 B.n222 B.n221 585
R454 B.n220 B.n177 585
R455 B.n219 B.n218 585
R456 B.n217 B.n178 585
R457 B.n216 B.n215 585
R458 B.n214 B.n179 585
R459 B.n213 B.n212 585
R460 B.n211 B.n180 585
R461 B.n210 B.n209 585
R462 B.n208 B.n181 585
R463 B.n207 B.n206 585
R464 B.n205 B.n182 585
R465 B.n204 B.n203 585
R466 B.n202 B.n183 585
R467 B.n201 B.n200 585
R468 B.n199 B.n184 585
R469 B.n198 B.n197 585
R470 B.n196 B.n185 585
R471 B.n195 B.n194 585
R472 B.n193 B.n186 585
R473 B.n192 B.n191 585
R474 B.n190 B.n187 585
R475 B.n189 B.n188 585
R476 B.n2 B.n0 585
R477 B.n729 B.n1 585
R478 B.n728 B.n727 585
R479 B.n726 B.n3 585
R480 B.n725 B.n724 585
R481 B.n723 B.n4 585
R482 B.n722 B.n721 585
R483 B.n720 B.n5 585
R484 B.n719 B.n718 585
R485 B.n717 B.n6 585
R486 B.n716 B.n715 585
R487 B.n714 B.n7 585
R488 B.n713 B.n712 585
R489 B.n711 B.n8 585
R490 B.n710 B.n709 585
R491 B.n708 B.n9 585
R492 B.n707 B.n706 585
R493 B.n705 B.n10 585
R494 B.n704 B.n703 585
R495 B.n702 B.n11 585
R496 B.n701 B.n700 585
R497 B.n699 B.n12 585
R498 B.n698 B.n697 585
R499 B.n696 B.n13 585
R500 B.n695 B.n694 585
R501 B.n693 B.n14 585
R502 B.n692 B.n691 585
R503 B.n690 B.n15 585
R504 B.n689 B.n688 585
R505 B.n687 B.n16 585
R506 B.n686 B.n685 585
R507 B.n684 B.n17 585
R508 B.n683 B.n682 585
R509 B.n681 B.n18 585
R510 B.n680 B.n679 585
R511 B.n678 B.n19 585
R512 B.n677 B.n676 585
R513 B.n675 B.n20 585
R514 B.n674 B.n673 585
R515 B.n672 B.n21 585
R516 B.n671 B.n670 585
R517 B.n669 B.n22 585
R518 B.n668 B.n667 585
R519 B.n666 B.n23 585
R520 B.n665 B.n664 585
R521 B.n663 B.n24 585
R522 B.n662 B.n661 585
R523 B.n660 B.n25 585
R524 B.n659 B.n658 585
R525 B.n657 B.n26 585
R526 B.n656 B.n655 585
R527 B.n654 B.n27 585
R528 B.n653 B.n652 585
R529 B.n651 B.n28 585
R530 B.n650 B.n649 585
R531 B.n648 B.n29 585
R532 B.n647 B.n646 585
R533 B.n645 B.n30 585
R534 B.n644 B.n643 585
R535 B.n642 B.n31 585
R536 B.n641 B.n640 585
R537 B.n639 B.n32 585
R538 B.n638 B.n637 585
R539 B.n636 B.n33 585
R540 B.n635 B.n634 585
R541 B.n731 B.n730 585
R542 B.n281 B.n156 473.281
R543 B.n634 B.n633 473.281
R544 B.n363 B.n362 473.281
R545 B.n555 B.n64 473.281
R546 B.n327 B.t3 243.119
R547 B.n145 B.t6 243.119
R548 B.n46 B.t9 243.119
R549 B.n53 B.t0 243.119
R550 B.n327 B.t5 190.69
R551 B.n53 B.t1 190.69
R552 B.n145 B.t8 190.685
R553 B.n46 B.t10 190.685
R554 B.n281 B.n280 163.367
R555 B.n280 B.n279 163.367
R556 B.n279 B.n158 163.367
R557 B.n275 B.n158 163.367
R558 B.n275 B.n274 163.367
R559 B.n274 B.n273 163.367
R560 B.n273 B.n160 163.367
R561 B.n269 B.n160 163.367
R562 B.n269 B.n268 163.367
R563 B.n268 B.n267 163.367
R564 B.n267 B.n162 163.367
R565 B.n263 B.n162 163.367
R566 B.n263 B.n262 163.367
R567 B.n262 B.n261 163.367
R568 B.n261 B.n164 163.367
R569 B.n257 B.n164 163.367
R570 B.n257 B.n256 163.367
R571 B.n256 B.n255 163.367
R572 B.n255 B.n166 163.367
R573 B.n251 B.n166 163.367
R574 B.n251 B.n250 163.367
R575 B.n250 B.n249 163.367
R576 B.n249 B.n168 163.367
R577 B.n245 B.n168 163.367
R578 B.n245 B.n244 163.367
R579 B.n244 B.n243 163.367
R580 B.n243 B.n170 163.367
R581 B.n239 B.n170 163.367
R582 B.n239 B.n238 163.367
R583 B.n238 B.n237 163.367
R584 B.n237 B.n172 163.367
R585 B.n233 B.n172 163.367
R586 B.n233 B.n232 163.367
R587 B.n232 B.n231 163.367
R588 B.n231 B.n174 163.367
R589 B.n227 B.n174 163.367
R590 B.n227 B.n226 163.367
R591 B.n226 B.n225 163.367
R592 B.n225 B.n176 163.367
R593 B.n221 B.n176 163.367
R594 B.n221 B.n220 163.367
R595 B.n220 B.n219 163.367
R596 B.n219 B.n178 163.367
R597 B.n215 B.n178 163.367
R598 B.n215 B.n214 163.367
R599 B.n214 B.n213 163.367
R600 B.n213 B.n180 163.367
R601 B.n209 B.n180 163.367
R602 B.n209 B.n208 163.367
R603 B.n208 B.n207 163.367
R604 B.n207 B.n182 163.367
R605 B.n203 B.n182 163.367
R606 B.n203 B.n202 163.367
R607 B.n202 B.n201 163.367
R608 B.n201 B.n184 163.367
R609 B.n197 B.n184 163.367
R610 B.n197 B.n196 163.367
R611 B.n196 B.n195 163.367
R612 B.n195 B.n186 163.367
R613 B.n191 B.n186 163.367
R614 B.n191 B.n190 163.367
R615 B.n190 B.n189 163.367
R616 B.n189 B.n2 163.367
R617 B.n730 B.n2 163.367
R618 B.n730 B.n729 163.367
R619 B.n729 B.n728 163.367
R620 B.n728 B.n3 163.367
R621 B.n724 B.n3 163.367
R622 B.n724 B.n723 163.367
R623 B.n723 B.n722 163.367
R624 B.n722 B.n5 163.367
R625 B.n718 B.n5 163.367
R626 B.n718 B.n717 163.367
R627 B.n717 B.n716 163.367
R628 B.n716 B.n7 163.367
R629 B.n712 B.n7 163.367
R630 B.n712 B.n711 163.367
R631 B.n711 B.n710 163.367
R632 B.n710 B.n9 163.367
R633 B.n706 B.n9 163.367
R634 B.n706 B.n705 163.367
R635 B.n705 B.n704 163.367
R636 B.n704 B.n11 163.367
R637 B.n700 B.n11 163.367
R638 B.n700 B.n699 163.367
R639 B.n699 B.n698 163.367
R640 B.n698 B.n13 163.367
R641 B.n694 B.n13 163.367
R642 B.n694 B.n693 163.367
R643 B.n693 B.n692 163.367
R644 B.n692 B.n15 163.367
R645 B.n688 B.n15 163.367
R646 B.n688 B.n687 163.367
R647 B.n687 B.n686 163.367
R648 B.n686 B.n17 163.367
R649 B.n682 B.n17 163.367
R650 B.n682 B.n681 163.367
R651 B.n681 B.n680 163.367
R652 B.n680 B.n19 163.367
R653 B.n676 B.n19 163.367
R654 B.n676 B.n675 163.367
R655 B.n675 B.n674 163.367
R656 B.n674 B.n21 163.367
R657 B.n670 B.n21 163.367
R658 B.n670 B.n669 163.367
R659 B.n669 B.n668 163.367
R660 B.n668 B.n23 163.367
R661 B.n664 B.n23 163.367
R662 B.n664 B.n663 163.367
R663 B.n663 B.n662 163.367
R664 B.n662 B.n25 163.367
R665 B.n658 B.n25 163.367
R666 B.n658 B.n657 163.367
R667 B.n657 B.n656 163.367
R668 B.n656 B.n27 163.367
R669 B.n652 B.n27 163.367
R670 B.n652 B.n651 163.367
R671 B.n651 B.n650 163.367
R672 B.n650 B.n29 163.367
R673 B.n646 B.n29 163.367
R674 B.n646 B.n645 163.367
R675 B.n645 B.n644 163.367
R676 B.n644 B.n31 163.367
R677 B.n640 B.n31 163.367
R678 B.n640 B.n639 163.367
R679 B.n639 B.n638 163.367
R680 B.n638 B.n33 163.367
R681 B.n634 B.n33 163.367
R682 B.n285 B.n156 163.367
R683 B.n286 B.n285 163.367
R684 B.n287 B.n286 163.367
R685 B.n287 B.n154 163.367
R686 B.n291 B.n154 163.367
R687 B.n292 B.n291 163.367
R688 B.n293 B.n292 163.367
R689 B.n293 B.n152 163.367
R690 B.n297 B.n152 163.367
R691 B.n298 B.n297 163.367
R692 B.n299 B.n298 163.367
R693 B.n299 B.n150 163.367
R694 B.n303 B.n150 163.367
R695 B.n304 B.n303 163.367
R696 B.n305 B.n304 163.367
R697 B.n305 B.n148 163.367
R698 B.n309 B.n148 163.367
R699 B.n310 B.n309 163.367
R700 B.n311 B.n310 163.367
R701 B.n311 B.n144 163.367
R702 B.n316 B.n144 163.367
R703 B.n317 B.n316 163.367
R704 B.n318 B.n317 163.367
R705 B.n318 B.n142 163.367
R706 B.n322 B.n142 163.367
R707 B.n323 B.n322 163.367
R708 B.n324 B.n323 163.367
R709 B.n324 B.n140 163.367
R710 B.n331 B.n140 163.367
R711 B.n332 B.n331 163.367
R712 B.n333 B.n332 163.367
R713 B.n333 B.n138 163.367
R714 B.n337 B.n138 163.367
R715 B.n338 B.n337 163.367
R716 B.n339 B.n338 163.367
R717 B.n339 B.n136 163.367
R718 B.n343 B.n136 163.367
R719 B.n344 B.n343 163.367
R720 B.n345 B.n344 163.367
R721 B.n345 B.n134 163.367
R722 B.n349 B.n134 163.367
R723 B.n350 B.n349 163.367
R724 B.n351 B.n350 163.367
R725 B.n351 B.n132 163.367
R726 B.n355 B.n132 163.367
R727 B.n356 B.n355 163.367
R728 B.n357 B.n356 163.367
R729 B.n357 B.n130 163.367
R730 B.n361 B.n130 163.367
R731 B.n362 B.n361 163.367
R732 B.n363 B.n128 163.367
R733 B.n367 B.n128 163.367
R734 B.n368 B.n367 163.367
R735 B.n369 B.n368 163.367
R736 B.n369 B.n126 163.367
R737 B.n373 B.n126 163.367
R738 B.n374 B.n373 163.367
R739 B.n375 B.n374 163.367
R740 B.n375 B.n124 163.367
R741 B.n379 B.n124 163.367
R742 B.n380 B.n379 163.367
R743 B.n381 B.n380 163.367
R744 B.n381 B.n122 163.367
R745 B.n385 B.n122 163.367
R746 B.n386 B.n385 163.367
R747 B.n387 B.n386 163.367
R748 B.n387 B.n120 163.367
R749 B.n391 B.n120 163.367
R750 B.n392 B.n391 163.367
R751 B.n393 B.n392 163.367
R752 B.n393 B.n118 163.367
R753 B.n397 B.n118 163.367
R754 B.n398 B.n397 163.367
R755 B.n399 B.n398 163.367
R756 B.n399 B.n116 163.367
R757 B.n403 B.n116 163.367
R758 B.n404 B.n403 163.367
R759 B.n405 B.n404 163.367
R760 B.n405 B.n114 163.367
R761 B.n409 B.n114 163.367
R762 B.n410 B.n409 163.367
R763 B.n411 B.n410 163.367
R764 B.n411 B.n112 163.367
R765 B.n415 B.n112 163.367
R766 B.n416 B.n415 163.367
R767 B.n417 B.n416 163.367
R768 B.n417 B.n110 163.367
R769 B.n421 B.n110 163.367
R770 B.n422 B.n421 163.367
R771 B.n423 B.n422 163.367
R772 B.n423 B.n108 163.367
R773 B.n427 B.n108 163.367
R774 B.n428 B.n427 163.367
R775 B.n429 B.n428 163.367
R776 B.n429 B.n106 163.367
R777 B.n433 B.n106 163.367
R778 B.n434 B.n433 163.367
R779 B.n435 B.n434 163.367
R780 B.n435 B.n104 163.367
R781 B.n439 B.n104 163.367
R782 B.n440 B.n439 163.367
R783 B.n441 B.n440 163.367
R784 B.n441 B.n102 163.367
R785 B.n445 B.n102 163.367
R786 B.n446 B.n445 163.367
R787 B.n447 B.n446 163.367
R788 B.n447 B.n100 163.367
R789 B.n451 B.n100 163.367
R790 B.n452 B.n451 163.367
R791 B.n453 B.n452 163.367
R792 B.n453 B.n98 163.367
R793 B.n457 B.n98 163.367
R794 B.n458 B.n457 163.367
R795 B.n459 B.n458 163.367
R796 B.n459 B.n96 163.367
R797 B.n463 B.n96 163.367
R798 B.n464 B.n463 163.367
R799 B.n465 B.n464 163.367
R800 B.n465 B.n94 163.367
R801 B.n469 B.n94 163.367
R802 B.n470 B.n469 163.367
R803 B.n471 B.n470 163.367
R804 B.n471 B.n92 163.367
R805 B.n475 B.n92 163.367
R806 B.n476 B.n475 163.367
R807 B.n477 B.n476 163.367
R808 B.n477 B.n90 163.367
R809 B.n481 B.n90 163.367
R810 B.n482 B.n481 163.367
R811 B.n483 B.n482 163.367
R812 B.n483 B.n88 163.367
R813 B.n487 B.n88 163.367
R814 B.n488 B.n487 163.367
R815 B.n489 B.n488 163.367
R816 B.n489 B.n86 163.367
R817 B.n493 B.n86 163.367
R818 B.n494 B.n493 163.367
R819 B.n495 B.n494 163.367
R820 B.n495 B.n84 163.367
R821 B.n499 B.n84 163.367
R822 B.n500 B.n499 163.367
R823 B.n501 B.n500 163.367
R824 B.n501 B.n82 163.367
R825 B.n505 B.n82 163.367
R826 B.n506 B.n505 163.367
R827 B.n507 B.n506 163.367
R828 B.n507 B.n80 163.367
R829 B.n511 B.n80 163.367
R830 B.n512 B.n511 163.367
R831 B.n513 B.n512 163.367
R832 B.n513 B.n78 163.367
R833 B.n517 B.n78 163.367
R834 B.n518 B.n517 163.367
R835 B.n519 B.n518 163.367
R836 B.n519 B.n76 163.367
R837 B.n523 B.n76 163.367
R838 B.n524 B.n523 163.367
R839 B.n525 B.n524 163.367
R840 B.n525 B.n74 163.367
R841 B.n529 B.n74 163.367
R842 B.n530 B.n529 163.367
R843 B.n531 B.n530 163.367
R844 B.n531 B.n72 163.367
R845 B.n535 B.n72 163.367
R846 B.n536 B.n535 163.367
R847 B.n537 B.n536 163.367
R848 B.n537 B.n70 163.367
R849 B.n541 B.n70 163.367
R850 B.n542 B.n541 163.367
R851 B.n543 B.n542 163.367
R852 B.n543 B.n68 163.367
R853 B.n547 B.n68 163.367
R854 B.n548 B.n547 163.367
R855 B.n549 B.n548 163.367
R856 B.n549 B.n66 163.367
R857 B.n553 B.n66 163.367
R858 B.n554 B.n553 163.367
R859 B.n555 B.n554 163.367
R860 B.n633 B.n632 163.367
R861 B.n632 B.n35 163.367
R862 B.n628 B.n35 163.367
R863 B.n628 B.n627 163.367
R864 B.n627 B.n626 163.367
R865 B.n626 B.n37 163.367
R866 B.n622 B.n37 163.367
R867 B.n622 B.n621 163.367
R868 B.n621 B.n620 163.367
R869 B.n620 B.n39 163.367
R870 B.n616 B.n39 163.367
R871 B.n616 B.n615 163.367
R872 B.n615 B.n614 163.367
R873 B.n614 B.n41 163.367
R874 B.n610 B.n41 163.367
R875 B.n610 B.n609 163.367
R876 B.n609 B.n608 163.367
R877 B.n608 B.n43 163.367
R878 B.n604 B.n43 163.367
R879 B.n604 B.n603 163.367
R880 B.n603 B.n602 163.367
R881 B.n602 B.n45 163.367
R882 B.n598 B.n45 163.367
R883 B.n598 B.n597 163.367
R884 B.n597 B.n596 163.367
R885 B.n596 B.n50 163.367
R886 B.n592 B.n50 163.367
R887 B.n592 B.n591 163.367
R888 B.n591 B.n590 163.367
R889 B.n590 B.n52 163.367
R890 B.n585 B.n52 163.367
R891 B.n585 B.n584 163.367
R892 B.n584 B.n583 163.367
R893 B.n583 B.n56 163.367
R894 B.n579 B.n56 163.367
R895 B.n579 B.n578 163.367
R896 B.n578 B.n577 163.367
R897 B.n577 B.n58 163.367
R898 B.n573 B.n58 163.367
R899 B.n573 B.n572 163.367
R900 B.n572 B.n571 163.367
R901 B.n571 B.n60 163.367
R902 B.n567 B.n60 163.367
R903 B.n567 B.n566 163.367
R904 B.n566 B.n565 163.367
R905 B.n565 B.n62 163.367
R906 B.n561 B.n62 163.367
R907 B.n561 B.n560 163.367
R908 B.n560 B.n559 163.367
R909 B.n559 B.n64 163.367
R910 B.n328 B.t4 117.186
R911 B.n54 B.t2 117.186
R912 B.n146 B.t7 117.183
R913 B.n47 B.t11 117.183
R914 B.n328 B.n327 73.5035
R915 B.n146 B.n145 73.5035
R916 B.n47 B.n46 73.5035
R917 B.n54 B.n53 73.5035
R918 B.n329 B.n328 59.5399
R919 B.n314 B.n146 59.5399
R920 B.n48 B.n47 59.5399
R921 B.n588 B.n54 59.5399
R922 B.n635 B.n34 30.7517
R923 B.n557 B.n556 30.7517
R924 B.n364 B.n129 30.7517
R925 B.n283 B.n282 30.7517
R926 B B.n731 18.0485
R927 B.n631 B.n34 10.6151
R928 B.n631 B.n630 10.6151
R929 B.n630 B.n629 10.6151
R930 B.n629 B.n36 10.6151
R931 B.n625 B.n36 10.6151
R932 B.n625 B.n624 10.6151
R933 B.n624 B.n623 10.6151
R934 B.n623 B.n38 10.6151
R935 B.n619 B.n38 10.6151
R936 B.n619 B.n618 10.6151
R937 B.n618 B.n617 10.6151
R938 B.n617 B.n40 10.6151
R939 B.n613 B.n40 10.6151
R940 B.n613 B.n612 10.6151
R941 B.n612 B.n611 10.6151
R942 B.n611 B.n42 10.6151
R943 B.n607 B.n42 10.6151
R944 B.n607 B.n606 10.6151
R945 B.n606 B.n605 10.6151
R946 B.n605 B.n44 10.6151
R947 B.n601 B.n600 10.6151
R948 B.n600 B.n599 10.6151
R949 B.n599 B.n49 10.6151
R950 B.n595 B.n49 10.6151
R951 B.n595 B.n594 10.6151
R952 B.n594 B.n593 10.6151
R953 B.n593 B.n51 10.6151
R954 B.n589 B.n51 10.6151
R955 B.n587 B.n586 10.6151
R956 B.n586 B.n55 10.6151
R957 B.n582 B.n55 10.6151
R958 B.n582 B.n581 10.6151
R959 B.n581 B.n580 10.6151
R960 B.n580 B.n57 10.6151
R961 B.n576 B.n57 10.6151
R962 B.n576 B.n575 10.6151
R963 B.n575 B.n574 10.6151
R964 B.n574 B.n59 10.6151
R965 B.n570 B.n59 10.6151
R966 B.n570 B.n569 10.6151
R967 B.n569 B.n568 10.6151
R968 B.n568 B.n61 10.6151
R969 B.n564 B.n61 10.6151
R970 B.n564 B.n563 10.6151
R971 B.n563 B.n562 10.6151
R972 B.n562 B.n63 10.6151
R973 B.n558 B.n63 10.6151
R974 B.n558 B.n557 10.6151
R975 B.n365 B.n364 10.6151
R976 B.n366 B.n365 10.6151
R977 B.n366 B.n127 10.6151
R978 B.n370 B.n127 10.6151
R979 B.n371 B.n370 10.6151
R980 B.n372 B.n371 10.6151
R981 B.n372 B.n125 10.6151
R982 B.n376 B.n125 10.6151
R983 B.n377 B.n376 10.6151
R984 B.n378 B.n377 10.6151
R985 B.n378 B.n123 10.6151
R986 B.n382 B.n123 10.6151
R987 B.n383 B.n382 10.6151
R988 B.n384 B.n383 10.6151
R989 B.n384 B.n121 10.6151
R990 B.n388 B.n121 10.6151
R991 B.n389 B.n388 10.6151
R992 B.n390 B.n389 10.6151
R993 B.n390 B.n119 10.6151
R994 B.n394 B.n119 10.6151
R995 B.n395 B.n394 10.6151
R996 B.n396 B.n395 10.6151
R997 B.n396 B.n117 10.6151
R998 B.n400 B.n117 10.6151
R999 B.n401 B.n400 10.6151
R1000 B.n402 B.n401 10.6151
R1001 B.n402 B.n115 10.6151
R1002 B.n406 B.n115 10.6151
R1003 B.n407 B.n406 10.6151
R1004 B.n408 B.n407 10.6151
R1005 B.n408 B.n113 10.6151
R1006 B.n412 B.n113 10.6151
R1007 B.n413 B.n412 10.6151
R1008 B.n414 B.n413 10.6151
R1009 B.n414 B.n111 10.6151
R1010 B.n418 B.n111 10.6151
R1011 B.n419 B.n418 10.6151
R1012 B.n420 B.n419 10.6151
R1013 B.n420 B.n109 10.6151
R1014 B.n424 B.n109 10.6151
R1015 B.n425 B.n424 10.6151
R1016 B.n426 B.n425 10.6151
R1017 B.n426 B.n107 10.6151
R1018 B.n430 B.n107 10.6151
R1019 B.n431 B.n430 10.6151
R1020 B.n432 B.n431 10.6151
R1021 B.n432 B.n105 10.6151
R1022 B.n436 B.n105 10.6151
R1023 B.n437 B.n436 10.6151
R1024 B.n438 B.n437 10.6151
R1025 B.n438 B.n103 10.6151
R1026 B.n442 B.n103 10.6151
R1027 B.n443 B.n442 10.6151
R1028 B.n444 B.n443 10.6151
R1029 B.n444 B.n101 10.6151
R1030 B.n448 B.n101 10.6151
R1031 B.n449 B.n448 10.6151
R1032 B.n450 B.n449 10.6151
R1033 B.n450 B.n99 10.6151
R1034 B.n454 B.n99 10.6151
R1035 B.n455 B.n454 10.6151
R1036 B.n456 B.n455 10.6151
R1037 B.n456 B.n97 10.6151
R1038 B.n460 B.n97 10.6151
R1039 B.n461 B.n460 10.6151
R1040 B.n462 B.n461 10.6151
R1041 B.n462 B.n95 10.6151
R1042 B.n466 B.n95 10.6151
R1043 B.n467 B.n466 10.6151
R1044 B.n468 B.n467 10.6151
R1045 B.n468 B.n93 10.6151
R1046 B.n472 B.n93 10.6151
R1047 B.n473 B.n472 10.6151
R1048 B.n474 B.n473 10.6151
R1049 B.n474 B.n91 10.6151
R1050 B.n478 B.n91 10.6151
R1051 B.n479 B.n478 10.6151
R1052 B.n480 B.n479 10.6151
R1053 B.n480 B.n89 10.6151
R1054 B.n484 B.n89 10.6151
R1055 B.n485 B.n484 10.6151
R1056 B.n486 B.n485 10.6151
R1057 B.n486 B.n87 10.6151
R1058 B.n490 B.n87 10.6151
R1059 B.n491 B.n490 10.6151
R1060 B.n492 B.n491 10.6151
R1061 B.n492 B.n85 10.6151
R1062 B.n496 B.n85 10.6151
R1063 B.n497 B.n496 10.6151
R1064 B.n498 B.n497 10.6151
R1065 B.n498 B.n83 10.6151
R1066 B.n502 B.n83 10.6151
R1067 B.n503 B.n502 10.6151
R1068 B.n504 B.n503 10.6151
R1069 B.n504 B.n81 10.6151
R1070 B.n508 B.n81 10.6151
R1071 B.n509 B.n508 10.6151
R1072 B.n510 B.n509 10.6151
R1073 B.n510 B.n79 10.6151
R1074 B.n514 B.n79 10.6151
R1075 B.n515 B.n514 10.6151
R1076 B.n516 B.n515 10.6151
R1077 B.n516 B.n77 10.6151
R1078 B.n520 B.n77 10.6151
R1079 B.n521 B.n520 10.6151
R1080 B.n522 B.n521 10.6151
R1081 B.n522 B.n75 10.6151
R1082 B.n526 B.n75 10.6151
R1083 B.n527 B.n526 10.6151
R1084 B.n528 B.n527 10.6151
R1085 B.n528 B.n73 10.6151
R1086 B.n532 B.n73 10.6151
R1087 B.n533 B.n532 10.6151
R1088 B.n534 B.n533 10.6151
R1089 B.n534 B.n71 10.6151
R1090 B.n538 B.n71 10.6151
R1091 B.n539 B.n538 10.6151
R1092 B.n540 B.n539 10.6151
R1093 B.n540 B.n69 10.6151
R1094 B.n544 B.n69 10.6151
R1095 B.n545 B.n544 10.6151
R1096 B.n546 B.n545 10.6151
R1097 B.n546 B.n67 10.6151
R1098 B.n550 B.n67 10.6151
R1099 B.n551 B.n550 10.6151
R1100 B.n552 B.n551 10.6151
R1101 B.n552 B.n65 10.6151
R1102 B.n556 B.n65 10.6151
R1103 B.n284 B.n283 10.6151
R1104 B.n284 B.n155 10.6151
R1105 B.n288 B.n155 10.6151
R1106 B.n289 B.n288 10.6151
R1107 B.n290 B.n289 10.6151
R1108 B.n290 B.n153 10.6151
R1109 B.n294 B.n153 10.6151
R1110 B.n295 B.n294 10.6151
R1111 B.n296 B.n295 10.6151
R1112 B.n296 B.n151 10.6151
R1113 B.n300 B.n151 10.6151
R1114 B.n301 B.n300 10.6151
R1115 B.n302 B.n301 10.6151
R1116 B.n302 B.n149 10.6151
R1117 B.n306 B.n149 10.6151
R1118 B.n307 B.n306 10.6151
R1119 B.n308 B.n307 10.6151
R1120 B.n308 B.n147 10.6151
R1121 B.n312 B.n147 10.6151
R1122 B.n313 B.n312 10.6151
R1123 B.n315 B.n143 10.6151
R1124 B.n319 B.n143 10.6151
R1125 B.n320 B.n319 10.6151
R1126 B.n321 B.n320 10.6151
R1127 B.n321 B.n141 10.6151
R1128 B.n325 B.n141 10.6151
R1129 B.n326 B.n325 10.6151
R1130 B.n330 B.n326 10.6151
R1131 B.n334 B.n139 10.6151
R1132 B.n335 B.n334 10.6151
R1133 B.n336 B.n335 10.6151
R1134 B.n336 B.n137 10.6151
R1135 B.n340 B.n137 10.6151
R1136 B.n341 B.n340 10.6151
R1137 B.n342 B.n341 10.6151
R1138 B.n342 B.n135 10.6151
R1139 B.n346 B.n135 10.6151
R1140 B.n347 B.n346 10.6151
R1141 B.n348 B.n347 10.6151
R1142 B.n348 B.n133 10.6151
R1143 B.n352 B.n133 10.6151
R1144 B.n353 B.n352 10.6151
R1145 B.n354 B.n353 10.6151
R1146 B.n354 B.n131 10.6151
R1147 B.n358 B.n131 10.6151
R1148 B.n359 B.n358 10.6151
R1149 B.n360 B.n359 10.6151
R1150 B.n360 B.n129 10.6151
R1151 B.n282 B.n157 10.6151
R1152 B.n278 B.n157 10.6151
R1153 B.n278 B.n277 10.6151
R1154 B.n277 B.n276 10.6151
R1155 B.n276 B.n159 10.6151
R1156 B.n272 B.n159 10.6151
R1157 B.n272 B.n271 10.6151
R1158 B.n271 B.n270 10.6151
R1159 B.n270 B.n161 10.6151
R1160 B.n266 B.n161 10.6151
R1161 B.n266 B.n265 10.6151
R1162 B.n265 B.n264 10.6151
R1163 B.n264 B.n163 10.6151
R1164 B.n260 B.n163 10.6151
R1165 B.n260 B.n259 10.6151
R1166 B.n259 B.n258 10.6151
R1167 B.n258 B.n165 10.6151
R1168 B.n254 B.n165 10.6151
R1169 B.n254 B.n253 10.6151
R1170 B.n253 B.n252 10.6151
R1171 B.n252 B.n167 10.6151
R1172 B.n248 B.n167 10.6151
R1173 B.n248 B.n247 10.6151
R1174 B.n247 B.n246 10.6151
R1175 B.n246 B.n169 10.6151
R1176 B.n242 B.n169 10.6151
R1177 B.n242 B.n241 10.6151
R1178 B.n241 B.n240 10.6151
R1179 B.n240 B.n171 10.6151
R1180 B.n236 B.n171 10.6151
R1181 B.n236 B.n235 10.6151
R1182 B.n235 B.n234 10.6151
R1183 B.n234 B.n173 10.6151
R1184 B.n230 B.n173 10.6151
R1185 B.n230 B.n229 10.6151
R1186 B.n229 B.n228 10.6151
R1187 B.n228 B.n175 10.6151
R1188 B.n224 B.n175 10.6151
R1189 B.n224 B.n223 10.6151
R1190 B.n223 B.n222 10.6151
R1191 B.n222 B.n177 10.6151
R1192 B.n218 B.n177 10.6151
R1193 B.n218 B.n217 10.6151
R1194 B.n217 B.n216 10.6151
R1195 B.n216 B.n179 10.6151
R1196 B.n212 B.n179 10.6151
R1197 B.n212 B.n211 10.6151
R1198 B.n211 B.n210 10.6151
R1199 B.n210 B.n181 10.6151
R1200 B.n206 B.n181 10.6151
R1201 B.n206 B.n205 10.6151
R1202 B.n205 B.n204 10.6151
R1203 B.n204 B.n183 10.6151
R1204 B.n200 B.n183 10.6151
R1205 B.n200 B.n199 10.6151
R1206 B.n199 B.n198 10.6151
R1207 B.n198 B.n185 10.6151
R1208 B.n194 B.n185 10.6151
R1209 B.n194 B.n193 10.6151
R1210 B.n193 B.n192 10.6151
R1211 B.n192 B.n187 10.6151
R1212 B.n188 B.n187 10.6151
R1213 B.n188 B.n0 10.6151
R1214 B.n727 B.n1 10.6151
R1215 B.n727 B.n726 10.6151
R1216 B.n726 B.n725 10.6151
R1217 B.n725 B.n4 10.6151
R1218 B.n721 B.n4 10.6151
R1219 B.n721 B.n720 10.6151
R1220 B.n720 B.n719 10.6151
R1221 B.n719 B.n6 10.6151
R1222 B.n715 B.n6 10.6151
R1223 B.n715 B.n714 10.6151
R1224 B.n714 B.n713 10.6151
R1225 B.n713 B.n8 10.6151
R1226 B.n709 B.n8 10.6151
R1227 B.n709 B.n708 10.6151
R1228 B.n708 B.n707 10.6151
R1229 B.n707 B.n10 10.6151
R1230 B.n703 B.n10 10.6151
R1231 B.n703 B.n702 10.6151
R1232 B.n702 B.n701 10.6151
R1233 B.n701 B.n12 10.6151
R1234 B.n697 B.n12 10.6151
R1235 B.n697 B.n696 10.6151
R1236 B.n696 B.n695 10.6151
R1237 B.n695 B.n14 10.6151
R1238 B.n691 B.n14 10.6151
R1239 B.n691 B.n690 10.6151
R1240 B.n690 B.n689 10.6151
R1241 B.n689 B.n16 10.6151
R1242 B.n685 B.n16 10.6151
R1243 B.n685 B.n684 10.6151
R1244 B.n684 B.n683 10.6151
R1245 B.n683 B.n18 10.6151
R1246 B.n679 B.n18 10.6151
R1247 B.n679 B.n678 10.6151
R1248 B.n678 B.n677 10.6151
R1249 B.n677 B.n20 10.6151
R1250 B.n673 B.n20 10.6151
R1251 B.n673 B.n672 10.6151
R1252 B.n672 B.n671 10.6151
R1253 B.n671 B.n22 10.6151
R1254 B.n667 B.n22 10.6151
R1255 B.n667 B.n666 10.6151
R1256 B.n666 B.n665 10.6151
R1257 B.n665 B.n24 10.6151
R1258 B.n661 B.n24 10.6151
R1259 B.n661 B.n660 10.6151
R1260 B.n660 B.n659 10.6151
R1261 B.n659 B.n26 10.6151
R1262 B.n655 B.n26 10.6151
R1263 B.n655 B.n654 10.6151
R1264 B.n654 B.n653 10.6151
R1265 B.n653 B.n28 10.6151
R1266 B.n649 B.n28 10.6151
R1267 B.n649 B.n648 10.6151
R1268 B.n648 B.n647 10.6151
R1269 B.n647 B.n30 10.6151
R1270 B.n643 B.n30 10.6151
R1271 B.n643 B.n642 10.6151
R1272 B.n642 B.n641 10.6151
R1273 B.n641 B.n32 10.6151
R1274 B.n637 B.n32 10.6151
R1275 B.n637 B.n636 10.6151
R1276 B.n636 B.n635 10.6151
R1277 B.n601 B.n48 6.5566
R1278 B.n589 B.n588 6.5566
R1279 B.n315 B.n314 6.5566
R1280 B.n330 B.n329 6.5566
R1281 B.n48 B.n44 4.05904
R1282 B.n588 B.n587 4.05904
R1283 B.n314 B.n313 4.05904
R1284 B.n329 B.n139 4.05904
R1285 B.n731 B.n0 2.81026
R1286 B.n731 B.n1 2.81026
R1287 VN.n68 VN.n67 161.3
R1288 VN.n66 VN.n36 161.3
R1289 VN.n65 VN.n64 161.3
R1290 VN.n63 VN.n37 161.3
R1291 VN.n62 VN.n61 161.3
R1292 VN.n60 VN.n38 161.3
R1293 VN.n59 VN.n58 161.3
R1294 VN.n57 VN.n39 161.3
R1295 VN.n56 VN.n55 161.3
R1296 VN.n54 VN.n40 161.3
R1297 VN.n53 VN.n52 161.3
R1298 VN.n51 VN.n42 161.3
R1299 VN.n50 VN.n49 161.3
R1300 VN.n48 VN.n43 161.3
R1301 VN.n47 VN.n46 161.3
R1302 VN.n33 VN.n32 161.3
R1303 VN.n31 VN.n1 161.3
R1304 VN.n30 VN.n29 161.3
R1305 VN.n28 VN.n2 161.3
R1306 VN.n27 VN.n26 161.3
R1307 VN.n25 VN.n3 161.3
R1308 VN.n24 VN.n23 161.3
R1309 VN.n22 VN.n4 161.3
R1310 VN.n21 VN.n20 161.3
R1311 VN.n18 VN.n5 161.3
R1312 VN.n17 VN.n16 161.3
R1313 VN.n15 VN.n6 161.3
R1314 VN.n14 VN.n13 161.3
R1315 VN.n12 VN.n7 161.3
R1316 VN.n11 VN.n10 161.3
R1317 VN.n34 VN.n0 81.0146
R1318 VN.n69 VN.n35 81.0146
R1319 VN.n45 VN.t2 67.3013
R1320 VN.n9 VN.t0 67.3013
R1321 VN.n26 VN.n2 56.5193
R1322 VN.n61 VN.n37 56.5193
R1323 VN.n9 VN.n8 55.2448
R1324 VN.n45 VN.n44 55.2448
R1325 VN VN.n69 49.7632
R1326 VN.n13 VN.n6 40.4934
R1327 VN.n17 VN.n6 40.4934
R1328 VN.n49 VN.n42 40.4934
R1329 VN.n53 VN.n42 40.4934
R1330 VN.n8 VN.t4 34.0609
R1331 VN.n19 VN.t3 34.0609
R1332 VN.n0 VN.t1 34.0609
R1333 VN.n44 VN.t5 34.0609
R1334 VN.n41 VN.t6 34.0609
R1335 VN.n35 VN.t7 34.0609
R1336 VN.n12 VN.n11 24.4675
R1337 VN.n13 VN.n12 24.4675
R1338 VN.n18 VN.n17 24.4675
R1339 VN.n20 VN.n18 24.4675
R1340 VN.n24 VN.n4 24.4675
R1341 VN.n25 VN.n24 24.4675
R1342 VN.n26 VN.n25 24.4675
R1343 VN.n30 VN.n2 24.4675
R1344 VN.n31 VN.n30 24.4675
R1345 VN.n32 VN.n31 24.4675
R1346 VN.n49 VN.n48 24.4675
R1347 VN.n48 VN.n47 24.4675
R1348 VN.n61 VN.n60 24.4675
R1349 VN.n60 VN.n59 24.4675
R1350 VN.n59 VN.n39 24.4675
R1351 VN.n55 VN.n54 24.4675
R1352 VN.n54 VN.n53 24.4675
R1353 VN.n67 VN.n66 24.4675
R1354 VN.n66 VN.n65 24.4675
R1355 VN.n65 VN.n37 24.4675
R1356 VN.n11 VN.n8 19.3294
R1357 VN.n20 VN.n19 19.3294
R1358 VN.n47 VN.n44 19.3294
R1359 VN.n55 VN.n41 19.3294
R1360 VN.n32 VN.n0 9.05329
R1361 VN.n67 VN.n35 9.05329
R1362 VN.n19 VN.n4 5.13857
R1363 VN.n41 VN.n39 5.13857
R1364 VN.n46 VN.n45 3.1879
R1365 VN.n10 VN.n9 3.1879
R1366 VN.n69 VN.n68 0.354971
R1367 VN.n34 VN.n33 0.354971
R1368 VN VN.n34 0.26696
R1369 VN.n68 VN.n36 0.189894
R1370 VN.n64 VN.n36 0.189894
R1371 VN.n64 VN.n63 0.189894
R1372 VN.n63 VN.n62 0.189894
R1373 VN.n62 VN.n38 0.189894
R1374 VN.n58 VN.n38 0.189894
R1375 VN.n58 VN.n57 0.189894
R1376 VN.n57 VN.n56 0.189894
R1377 VN.n56 VN.n40 0.189894
R1378 VN.n52 VN.n40 0.189894
R1379 VN.n52 VN.n51 0.189894
R1380 VN.n51 VN.n50 0.189894
R1381 VN.n50 VN.n43 0.189894
R1382 VN.n46 VN.n43 0.189894
R1383 VN.n10 VN.n7 0.189894
R1384 VN.n14 VN.n7 0.189894
R1385 VN.n15 VN.n14 0.189894
R1386 VN.n16 VN.n15 0.189894
R1387 VN.n16 VN.n5 0.189894
R1388 VN.n21 VN.n5 0.189894
R1389 VN.n22 VN.n21 0.189894
R1390 VN.n23 VN.n22 0.189894
R1391 VN.n23 VN.n3 0.189894
R1392 VN.n27 VN.n3 0.189894
R1393 VN.n28 VN.n27 0.189894
R1394 VN.n29 VN.n28 0.189894
R1395 VN.n29 VN.n1 0.189894
R1396 VN.n33 VN.n1 0.189894
R1397 VDD2.n2 VDD2.n1 101.438
R1398 VDD2.n2 VDD2.n0 101.438
R1399 VDD2 VDD2.n5 101.434
R1400 VDD2.n4 VDD2.n3 99.859
R1401 VDD2.n4 VDD2.n2 42.6334
R1402 VDD2.n5 VDD2.t2 6.64774
R1403 VDD2.n5 VDD2.t5 6.64774
R1404 VDD2.n3 VDD2.t0 6.64774
R1405 VDD2.n3 VDD2.t1 6.64774
R1406 VDD2.n1 VDD2.t4 6.64774
R1407 VDD2.n1 VDD2.t6 6.64774
R1408 VDD2.n0 VDD2.t7 6.64774
R1409 VDD2.n0 VDD2.t3 6.64774
R1410 VDD2 VDD2.n4 1.69231
C0 B VTAIL 2.88188f
C1 VDD1 VTAIL 6.34502f
C2 VN VTAIL 5.2659f
C3 VDD2 B 1.84357f
C4 VDD1 VDD2 2.22384f
C5 VP B 2.43073f
C6 VDD1 VP 4.45431f
C7 VN VDD2 3.99841f
C8 VN VP 7.40003f
C9 w_n4760_n1946# B 9.456571f
C10 w_n4760_n1946# VDD1 2.04272f
C11 VDD2 VTAIL 6.4052f
C12 VN w_n4760_n1946# 9.815281f
C13 VP VTAIL 5.28001f
C14 VDD2 VP 0.615712f
C15 w_n4760_n1946# VTAIL 2.71189f
C16 VDD1 B 1.72035f
C17 VN B 1.38608f
C18 w_n4760_n1946# VDD2 2.19319f
C19 VN VDD1 0.157219f
C20 w_n4760_n1946# VP 10.4357f
C21 VDD2 VSUBS 2.163847f
C22 VDD1 VSUBS 2.96488f
C23 VTAIL VSUBS 0.750007f
C24 VN VSUBS 7.65251f
C25 VP VSUBS 3.901649f
C26 B VSUBS 5.041225f
C27 w_n4760_n1946# VSUBS 0.116125p
C28 VDD2.t7 VSUBS 0.132184f
C29 VDD2.t3 VSUBS 0.132184f
C30 VDD2.n0 VSUBS 0.84058f
C31 VDD2.t4 VSUBS 0.132184f
C32 VDD2.t6 VSUBS 0.132184f
C33 VDD2.n1 VSUBS 0.84058f
C34 VDD2.n2 VSUBS 5.04794f
C35 VDD2.t0 VSUBS 0.132184f
C36 VDD2.t1 VSUBS 0.132184f
C37 VDD2.n3 VSUBS 0.823948f
C38 VDD2.n4 VSUBS 3.937f
C39 VDD2.t2 VSUBS 0.132184f
C40 VDD2.t5 VSUBS 0.132184f
C41 VDD2.n5 VSUBS 0.840537f
C42 VN.t1 VSUBS 1.56086f
C43 VN.n0 VSUBS 0.723774f
C44 VN.n1 VSUBS 0.035326f
C45 VN.n2 VSUBS 0.047633f
C46 VN.n3 VSUBS 0.035326f
C47 VN.n4 VSUBS 0.040159f
C48 VN.n5 VSUBS 0.035326f
C49 VN.n6 VSUBS 0.028558f
C50 VN.n7 VSUBS 0.035326f
C51 VN.t4 VSUBS 1.56086f
C52 VN.n8 VSUBS 0.722089f
C53 VN.t0 VSUBS 1.98216f
C54 VN.n9 VSUBS 0.692972f
C55 VN.n10 VSUBS 0.435409f
C56 VN.n11 VSUBS 0.059012f
C57 VN.n12 VSUBS 0.06584f
C58 VN.n13 VSUBS 0.070211f
C59 VN.n14 VSUBS 0.035326f
C60 VN.n15 VSUBS 0.035326f
C61 VN.n16 VSUBS 0.035326f
C62 VN.n17 VSUBS 0.070211f
C63 VN.n18 VSUBS 0.06584f
C64 VN.t3 VSUBS 1.56086f
C65 VN.n19 VSUBS 0.590849f
C66 VN.n20 VSUBS 0.059012f
C67 VN.n21 VSUBS 0.035326f
C68 VN.n22 VSUBS 0.035326f
C69 VN.n23 VSUBS 0.035326f
C70 VN.n24 VSUBS 0.06584f
C71 VN.n25 VSUBS 0.06584f
C72 VN.n26 VSUBS 0.055508f
C73 VN.n27 VSUBS 0.035326f
C74 VN.n28 VSUBS 0.035326f
C75 VN.n29 VSUBS 0.035326f
C76 VN.n30 VSUBS 0.06584f
C77 VN.n31 VSUBS 0.06584f
C78 VN.n32 VSUBS 0.04536f
C79 VN.n33 VSUBS 0.057016f
C80 VN.n34 VSUBS 0.09536f
C81 VN.t7 VSUBS 1.56086f
C82 VN.n35 VSUBS 0.723774f
C83 VN.n36 VSUBS 0.035326f
C84 VN.n37 VSUBS 0.047633f
C85 VN.n38 VSUBS 0.035326f
C86 VN.n39 VSUBS 0.040159f
C87 VN.n40 VSUBS 0.035326f
C88 VN.t6 VSUBS 1.56086f
C89 VN.n41 VSUBS 0.590849f
C90 VN.n42 VSUBS 0.028558f
C91 VN.n43 VSUBS 0.035326f
C92 VN.t5 VSUBS 1.56086f
C93 VN.n44 VSUBS 0.722089f
C94 VN.t2 VSUBS 1.98216f
C95 VN.n45 VSUBS 0.692972f
C96 VN.n46 VSUBS 0.435409f
C97 VN.n47 VSUBS 0.059012f
C98 VN.n48 VSUBS 0.06584f
C99 VN.n49 VSUBS 0.070211f
C100 VN.n50 VSUBS 0.035326f
C101 VN.n51 VSUBS 0.035326f
C102 VN.n52 VSUBS 0.035326f
C103 VN.n53 VSUBS 0.070211f
C104 VN.n54 VSUBS 0.06584f
C105 VN.n55 VSUBS 0.059012f
C106 VN.n56 VSUBS 0.035326f
C107 VN.n57 VSUBS 0.035326f
C108 VN.n58 VSUBS 0.035326f
C109 VN.n59 VSUBS 0.06584f
C110 VN.n60 VSUBS 0.06584f
C111 VN.n61 VSUBS 0.055508f
C112 VN.n62 VSUBS 0.035326f
C113 VN.n63 VSUBS 0.035326f
C114 VN.n64 VSUBS 0.035326f
C115 VN.n65 VSUBS 0.06584f
C116 VN.n66 VSUBS 0.06584f
C117 VN.n67 VSUBS 0.04536f
C118 VN.n68 VSUBS 0.057016f
C119 VN.n69 VSUBS 2.01007f
C120 B.n0 VSUBS 0.006285f
C121 B.n1 VSUBS 0.006285f
C122 B.n2 VSUBS 0.009938f
C123 B.n3 VSUBS 0.009938f
C124 B.n4 VSUBS 0.009938f
C125 B.n5 VSUBS 0.009938f
C126 B.n6 VSUBS 0.009938f
C127 B.n7 VSUBS 0.009938f
C128 B.n8 VSUBS 0.009938f
C129 B.n9 VSUBS 0.009938f
C130 B.n10 VSUBS 0.009938f
C131 B.n11 VSUBS 0.009938f
C132 B.n12 VSUBS 0.009938f
C133 B.n13 VSUBS 0.009938f
C134 B.n14 VSUBS 0.009938f
C135 B.n15 VSUBS 0.009938f
C136 B.n16 VSUBS 0.009938f
C137 B.n17 VSUBS 0.009938f
C138 B.n18 VSUBS 0.009938f
C139 B.n19 VSUBS 0.009938f
C140 B.n20 VSUBS 0.009938f
C141 B.n21 VSUBS 0.009938f
C142 B.n22 VSUBS 0.009938f
C143 B.n23 VSUBS 0.009938f
C144 B.n24 VSUBS 0.009938f
C145 B.n25 VSUBS 0.009938f
C146 B.n26 VSUBS 0.009938f
C147 B.n27 VSUBS 0.009938f
C148 B.n28 VSUBS 0.009938f
C149 B.n29 VSUBS 0.009938f
C150 B.n30 VSUBS 0.009938f
C151 B.n31 VSUBS 0.009938f
C152 B.n32 VSUBS 0.009938f
C153 B.n33 VSUBS 0.009938f
C154 B.n34 VSUBS 0.022802f
C155 B.n35 VSUBS 0.009938f
C156 B.n36 VSUBS 0.009938f
C157 B.n37 VSUBS 0.009938f
C158 B.n38 VSUBS 0.009938f
C159 B.n39 VSUBS 0.009938f
C160 B.n40 VSUBS 0.009938f
C161 B.n41 VSUBS 0.009938f
C162 B.n42 VSUBS 0.009938f
C163 B.n43 VSUBS 0.009938f
C164 B.n44 VSUBS 0.006869f
C165 B.n45 VSUBS 0.009938f
C166 B.t11 VSUBS 0.192851f
C167 B.t10 VSUBS 0.227626f
C168 B.t9 VSUBS 1.15918f
C169 B.n46 VSUBS 0.154849f
C170 B.n47 VSUBS 0.10439f
C171 B.n48 VSUBS 0.023026f
C172 B.n49 VSUBS 0.009938f
C173 B.n50 VSUBS 0.009938f
C174 B.n51 VSUBS 0.009938f
C175 B.n52 VSUBS 0.009938f
C176 B.t2 VSUBS 0.19285f
C177 B.t1 VSUBS 0.227625f
C178 B.t0 VSUBS 1.15918f
C179 B.n53 VSUBS 0.15485f
C180 B.n54 VSUBS 0.10439f
C181 B.n55 VSUBS 0.009938f
C182 B.n56 VSUBS 0.009938f
C183 B.n57 VSUBS 0.009938f
C184 B.n58 VSUBS 0.009938f
C185 B.n59 VSUBS 0.009938f
C186 B.n60 VSUBS 0.009938f
C187 B.n61 VSUBS 0.009938f
C188 B.n62 VSUBS 0.009938f
C189 B.n63 VSUBS 0.009938f
C190 B.n64 VSUBS 0.022802f
C191 B.n65 VSUBS 0.009938f
C192 B.n66 VSUBS 0.009938f
C193 B.n67 VSUBS 0.009938f
C194 B.n68 VSUBS 0.009938f
C195 B.n69 VSUBS 0.009938f
C196 B.n70 VSUBS 0.009938f
C197 B.n71 VSUBS 0.009938f
C198 B.n72 VSUBS 0.009938f
C199 B.n73 VSUBS 0.009938f
C200 B.n74 VSUBS 0.009938f
C201 B.n75 VSUBS 0.009938f
C202 B.n76 VSUBS 0.009938f
C203 B.n77 VSUBS 0.009938f
C204 B.n78 VSUBS 0.009938f
C205 B.n79 VSUBS 0.009938f
C206 B.n80 VSUBS 0.009938f
C207 B.n81 VSUBS 0.009938f
C208 B.n82 VSUBS 0.009938f
C209 B.n83 VSUBS 0.009938f
C210 B.n84 VSUBS 0.009938f
C211 B.n85 VSUBS 0.009938f
C212 B.n86 VSUBS 0.009938f
C213 B.n87 VSUBS 0.009938f
C214 B.n88 VSUBS 0.009938f
C215 B.n89 VSUBS 0.009938f
C216 B.n90 VSUBS 0.009938f
C217 B.n91 VSUBS 0.009938f
C218 B.n92 VSUBS 0.009938f
C219 B.n93 VSUBS 0.009938f
C220 B.n94 VSUBS 0.009938f
C221 B.n95 VSUBS 0.009938f
C222 B.n96 VSUBS 0.009938f
C223 B.n97 VSUBS 0.009938f
C224 B.n98 VSUBS 0.009938f
C225 B.n99 VSUBS 0.009938f
C226 B.n100 VSUBS 0.009938f
C227 B.n101 VSUBS 0.009938f
C228 B.n102 VSUBS 0.009938f
C229 B.n103 VSUBS 0.009938f
C230 B.n104 VSUBS 0.009938f
C231 B.n105 VSUBS 0.009938f
C232 B.n106 VSUBS 0.009938f
C233 B.n107 VSUBS 0.009938f
C234 B.n108 VSUBS 0.009938f
C235 B.n109 VSUBS 0.009938f
C236 B.n110 VSUBS 0.009938f
C237 B.n111 VSUBS 0.009938f
C238 B.n112 VSUBS 0.009938f
C239 B.n113 VSUBS 0.009938f
C240 B.n114 VSUBS 0.009938f
C241 B.n115 VSUBS 0.009938f
C242 B.n116 VSUBS 0.009938f
C243 B.n117 VSUBS 0.009938f
C244 B.n118 VSUBS 0.009938f
C245 B.n119 VSUBS 0.009938f
C246 B.n120 VSUBS 0.009938f
C247 B.n121 VSUBS 0.009938f
C248 B.n122 VSUBS 0.009938f
C249 B.n123 VSUBS 0.009938f
C250 B.n124 VSUBS 0.009938f
C251 B.n125 VSUBS 0.009938f
C252 B.n126 VSUBS 0.009938f
C253 B.n127 VSUBS 0.009938f
C254 B.n128 VSUBS 0.009938f
C255 B.n129 VSUBS 0.022802f
C256 B.n130 VSUBS 0.009938f
C257 B.n131 VSUBS 0.009938f
C258 B.n132 VSUBS 0.009938f
C259 B.n133 VSUBS 0.009938f
C260 B.n134 VSUBS 0.009938f
C261 B.n135 VSUBS 0.009938f
C262 B.n136 VSUBS 0.009938f
C263 B.n137 VSUBS 0.009938f
C264 B.n138 VSUBS 0.009938f
C265 B.n139 VSUBS 0.006869f
C266 B.n140 VSUBS 0.009938f
C267 B.n141 VSUBS 0.009938f
C268 B.n142 VSUBS 0.009938f
C269 B.n143 VSUBS 0.009938f
C270 B.n144 VSUBS 0.009938f
C271 B.t7 VSUBS 0.192851f
C272 B.t8 VSUBS 0.227626f
C273 B.t6 VSUBS 1.15918f
C274 B.n145 VSUBS 0.154849f
C275 B.n146 VSUBS 0.10439f
C276 B.n147 VSUBS 0.009938f
C277 B.n148 VSUBS 0.009938f
C278 B.n149 VSUBS 0.009938f
C279 B.n150 VSUBS 0.009938f
C280 B.n151 VSUBS 0.009938f
C281 B.n152 VSUBS 0.009938f
C282 B.n153 VSUBS 0.009938f
C283 B.n154 VSUBS 0.009938f
C284 B.n155 VSUBS 0.009938f
C285 B.n156 VSUBS 0.022802f
C286 B.n157 VSUBS 0.009938f
C287 B.n158 VSUBS 0.009938f
C288 B.n159 VSUBS 0.009938f
C289 B.n160 VSUBS 0.009938f
C290 B.n161 VSUBS 0.009938f
C291 B.n162 VSUBS 0.009938f
C292 B.n163 VSUBS 0.009938f
C293 B.n164 VSUBS 0.009938f
C294 B.n165 VSUBS 0.009938f
C295 B.n166 VSUBS 0.009938f
C296 B.n167 VSUBS 0.009938f
C297 B.n168 VSUBS 0.009938f
C298 B.n169 VSUBS 0.009938f
C299 B.n170 VSUBS 0.009938f
C300 B.n171 VSUBS 0.009938f
C301 B.n172 VSUBS 0.009938f
C302 B.n173 VSUBS 0.009938f
C303 B.n174 VSUBS 0.009938f
C304 B.n175 VSUBS 0.009938f
C305 B.n176 VSUBS 0.009938f
C306 B.n177 VSUBS 0.009938f
C307 B.n178 VSUBS 0.009938f
C308 B.n179 VSUBS 0.009938f
C309 B.n180 VSUBS 0.009938f
C310 B.n181 VSUBS 0.009938f
C311 B.n182 VSUBS 0.009938f
C312 B.n183 VSUBS 0.009938f
C313 B.n184 VSUBS 0.009938f
C314 B.n185 VSUBS 0.009938f
C315 B.n186 VSUBS 0.009938f
C316 B.n187 VSUBS 0.009938f
C317 B.n188 VSUBS 0.009938f
C318 B.n189 VSUBS 0.009938f
C319 B.n190 VSUBS 0.009938f
C320 B.n191 VSUBS 0.009938f
C321 B.n192 VSUBS 0.009938f
C322 B.n193 VSUBS 0.009938f
C323 B.n194 VSUBS 0.009938f
C324 B.n195 VSUBS 0.009938f
C325 B.n196 VSUBS 0.009938f
C326 B.n197 VSUBS 0.009938f
C327 B.n198 VSUBS 0.009938f
C328 B.n199 VSUBS 0.009938f
C329 B.n200 VSUBS 0.009938f
C330 B.n201 VSUBS 0.009938f
C331 B.n202 VSUBS 0.009938f
C332 B.n203 VSUBS 0.009938f
C333 B.n204 VSUBS 0.009938f
C334 B.n205 VSUBS 0.009938f
C335 B.n206 VSUBS 0.009938f
C336 B.n207 VSUBS 0.009938f
C337 B.n208 VSUBS 0.009938f
C338 B.n209 VSUBS 0.009938f
C339 B.n210 VSUBS 0.009938f
C340 B.n211 VSUBS 0.009938f
C341 B.n212 VSUBS 0.009938f
C342 B.n213 VSUBS 0.009938f
C343 B.n214 VSUBS 0.009938f
C344 B.n215 VSUBS 0.009938f
C345 B.n216 VSUBS 0.009938f
C346 B.n217 VSUBS 0.009938f
C347 B.n218 VSUBS 0.009938f
C348 B.n219 VSUBS 0.009938f
C349 B.n220 VSUBS 0.009938f
C350 B.n221 VSUBS 0.009938f
C351 B.n222 VSUBS 0.009938f
C352 B.n223 VSUBS 0.009938f
C353 B.n224 VSUBS 0.009938f
C354 B.n225 VSUBS 0.009938f
C355 B.n226 VSUBS 0.009938f
C356 B.n227 VSUBS 0.009938f
C357 B.n228 VSUBS 0.009938f
C358 B.n229 VSUBS 0.009938f
C359 B.n230 VSUBS 0.009938f
C360 B.n231 VSUBS 0.009938f
C361 B.n232 VSUBS 0.009938f
C362 B.n233 VSUBS 0.009938f
C363 B.n234 VSUBS 0.009938f
C364 B.n235 VSUBS 0.009938f
C365 B.n236 VSUBS 0.009938f
C366 B.n237 VSUBS 0.009938f
C367 B.n238 VSUBS 0.009938f
C368 B.n239 VSUBS 0.009938f
C369 B.n240 VSUBS 0.009938f
C370 B.n241 VSUBS 0.009938f
C371 B.n242 VSUBS 0.009938f
C372 B.n243 VSUBS 0.009938f
C373 B.n244 VSUBS 0.009938f
C374 B.n245 VSUBS 0.009938f
C375 B.n246 VSUBS 0.009938f
C376 B.n247 VSUBS 0.009938f
C377 B.n248 VSUBS 0.009938f
C378 B.n249 VSUBS 0.009938f
C379 B.n250 VSUBS 0.009938f
C380 B.n251 VSUBS 0.009938f
C381 B.n252 VSUBS 0.009938f
C382 B.n253 VSUBS 0.009938f
C383 B.n254 VSUBS 0.009938f
C384 B.n255 VSUBS 0.009938f
C385 B.n256 VSUBS 0.009938f
C386 B.n257 VSUBS 0.009938f
C387 B.n258 VSUBS 0.009938f
C388 B.n259 VSUBS 0.009938f
C389 B.n260 VSUBS 0.009938f
C390 B.n261 VSUBS 0.009938f
C391 B.n262 VSUBS 0.009938f
C392 B.n263 VSUBS 0.009938f
C393 B.n264 VSUBS 0.009938f
C394 B.n265 VSUBS 0.009938f
C395 B.n266 VSUBS 0.009938f
C396 B.n267 VSUBS 0.009938f
C397 B.n268 VSUBS 0.009938f
C398 B.n269 VSUBS 0.009938f
C399 B.n270 VSUBS 0.009938f
C400 B.n271 VSUBS 0.009938f
C401 B.n272 VSUBS 0.009938f
C402 B.n273 VSUBS 0.009938f
C403 B.n274 VSUBS 0.009938f
C404 B.n275 VSUBS 0.009938f
C405 B.n276 VSUBS 0.009938f
C406 B.n277 VSUBS 0.009938f
C407 B.n278 VSUBS 0.009938f
C408 B.n279 VSUBS 0.009938f
C409 B.n280 VSUBS 0.009938f
C410 B.n281 VSUBS 0.02192f
C411 B.n282 VSUBS 0.02192f
C412 B.n283 VSUBS 0.022802f
C413 B.n284 VSUBS 0.009938f
C414 B.n285 VSUBS 0.009938f
C415 B.n286 VSUBS 0.009938f
C416 B.n287 VSUBS 0.009938f
C417 B.n288 VSUBS 0.009938f
C418 B.n289 VSUBS 0.009938f
C419 B.n290 VSUBS 0.009938f
C420 B.n291 VSUBS 0.009938f
C421 B.n292 VSUBS 0.009938f
C422 B.n293 VSUBS 0.009938f
C423 B.n294 VSUBS 0.009938f
C424 B.n295 VSUBS 0.009938f
C425 B.n296 VSUBS 0.009938f
C426 B.n297 VSUBS 0.009938f
C427 B.n298 VSUBS 0.009938f
C428 B.n299 VSUBS 0.009938f
C429 B.n300 VSUBS 0.009938f
C430 B.n301 VSUBS 0.009938f
C431 B.n302 VSUBS 0.009938f
C432 B.n303 VSUBS 0.009938f
C433 B.n304 VSUBS 0.009938f
C434 B.n305 VSUBS 0.009938f
C435 B.n306 VSUBS 0.009938f
C436 B.n307 VSUBS 0.009938f
C437 B.n308 VSUBS 0.009938f
C438 B.n309 VSUBS 0.009938f
C439 B.n310 VSUBS 0.009938f
C440 B.n311 VSUBS 0.009938f
C441 B.n312 VSUBS 0.009938f
C442 B.n313 VSUBS 0.006869f
C443 B.n314 VSUBS 0.023026f
C444 B.n315 VSUBS 0.008038f
C445 B.n316 VSUBS 0.009938f
C446 B.n317 VSUBS 0.009938f
C447 B.n318 VSUBS 0.009938f
C448 B.n319 VSUBS 0.009938f
C449 B.n320 VSUBS 0.009938f
C450 B.n321 VSUBS 0.009938f
C451 B.n322 VSUBS 0.009938f
C452 B.n323 VSUBS 0.009938f
C453 B.n324 VSUBS 0.009938f
C454 B.n325 VSUBS 0.009938f
C455 B.n326 VSUBS 0.009938f
C456 B.t4 VSUBS 0.19285f
C457 B.t5 VSUBS 0.227625f
C458 B.t3 VSUBS 1.15918f
C459 B.n327 VSUBS 0.15485f
C460 B.n328 VSUBS 0.10439f
C461 B.n329 VSUBS 0.023026f
C462 B.n330 VSUBS 0.008038f
C463 B.n331 VSUBS 0.009938f
C464 B.n332 VSUBS 0.009938f
C465 B.n333 VSUBS 0.009938f
C466 B.n334 VSUBS 0.009938f
C467 B.n335 VSUBS 0.009938f
C468 B.n336 VSUBS 0.009938f
C469 B.n337 VSUBS 0.009938f
C470 B.n338 VSUBS 0.009938f
C471 B.n339 VSUBS 0.009938f
C472 B.n340 VSUBS 0.009938f
C473 B.n341 VSUBS 0.009938f
C474 B.n342 VSUBS 0.009938f
C475 B.n343 VSUBS 0.009938f
C476 B.n344 VSUBS 0.009938f
C477 B.n345 VSUBS 0.009938f
C478 B.n346 VSUBS 0.009938f
C479 B.n347 VSUBS 0.009938f
C480 B.n348 VSUBS 0.009938f
C481 B.n349 VSUBS 0.009938f
C482 B.n350 VSUBS 0.009938f
C483 B.n351 VSUBS 0.009938f
C484 B.n352 VSUBS 0.009938f
C485 B.n353 VSUBS 0.009938f
C486 B.n354 VSUBS 0.009938f
C487 B.n355 VSUBS 0.009938f
C488 B.n356 VSUBS 0.009938f
C489 B.n357 VSUBS 0.009938f
C490 B.n358 VSUBS 0.009938f
C491 B.n359 VSUBS 0.009938f
C492 B.n360 VSUBS 0.009938f
C493 B.n361 VSUBS 0.009938f
C494 B.n362 VSUBS 0.022802f
C495 B.n363 VSUBS 0.02192f
C496 B.n364 VSUBS 0.02192f
C497 B.n365 VSUBS 0.009938f
C498 B.n366 VSUBS 0.009938f
C499 B.n367 VSUBS 0.009938f
C500 B.n368 VSUBS 0.009938f
C501 B.n369 VSUBS 0.009938f
C502 B.n370 VSUBS 0.009938f
C503 B.n371 VSUBS 0.009938f
C504 B.n372 VSUBS 0.009938f
C505 B.n373 VSUBS 0.009938f
C506 B.n374 VSUBS 0.009938f
C507 B.n375 VSUBS 0.009938f
C508 B.n376 VSUBS 0.009938f
C509 B.n377 VSUBS 0.009938f
C510 B.n378 VSUBS 0.009938f
C511 B.n379 VSUBS 0.009938f
C512 B.n380 VSUBS 0.009938f
C513 B.n381 VSUBS 0.009938f
C514 B.n382 VSUBS 0.009938f
C515 B.n383 VSUBS 0.009938f
C516 B.n384 VSUBS 0.009938f
C517 B.n385 VSUBS 0.009938f
C518 B.n386 VSUBS 0.009938f
C519 B.n387 VSUBS 0.009938f
C520 B.n388 VSUBS 0.009938f
C521 B.n389 VSUBS 0.009938f
C522 B.n390 VSUBS 0.009938f
C523 B.n391 VSUBS 0.009938f
C524 B.n392 VSUBS 0.009938f
C525 B.n393 VSUBS 0.009938f
C526 B.n394 VSUBS 0.009938f
C527 B.n395 VSUBS 0.009938f
C528 B.n396 VSUBS 0.009938f
C529 B.n397 VSUBS 0.009938f
C530 B.n398 VSUBS 0.009938f
C531 B.n399 VSUBS 0.009938f
C532 B.n400 VSUBS 0.009938f
C533 B.n401 VSUBS 0.009938f
C534 B.n402 VSUBS 0.009938f
C535 B.n403 VSUBS 0.009938f
C536 B.n404 VSUBS 0.009938f
C537 B.n405 VSUBS 0.009938f
C538 B.n406 VSUBS 0.009938f
C539 B.n407 VSUBS 0.009938f
C540 B.n408 VSUBS 0.009938f
C541 B.n409 VSUBS 0.009938f
C542 B.n410 VSUBS 0.009938f
C543 B.n411 VSUBS 0.009938f
C544 B.n412 VSUBS 0.009938f
C545 B.n413 VSUBS 0.009938f
C546 B.n414 VSUBS 0.009938f
C547 B.n415 VSUBS 0.009938f
C548 B.n416 VSUBS 0.009938f
C549 B.n417 VSUBS 0.009938f
C550 B.n418 VSUBS 0.009938f
C551 B.n419 VSUBS 0.009938f
C552 B.n420 VSUBS 0.009938f
C553 B.n421 VSUBS 0.009938f
C554 B.n422 VSUBS 0.009938f
C555 B.n423 VSUBS 0.009938f
C556 B.n424 VSUBS 0.009938f
C557 B.n425 VSUBS 0.009938f
C558 B.n426 VSUBS 0.009938f
C559 B.n427 VSUBS 0.009938f
C560 B.n428 VSUBS 0.009938f
C561 B.n429 VSUBS 0.009938f
C562 B.n430 VSUBS 0.009938f
C563 B.n431 VSUBS 0.009938f
C564 B.n432 VSUBS 0.009938f
C565 B.n433 VSUBS 0.009938f
C566 B.n434 VSUBS 0.009938f
C567 B.n435 VSUBS 0.009938f
C568 B.n436 VSUBS 0.009938f
C569 B.n437 VSUBS 0.009938f
C570 B.n438 VSUBS 0.009938f
C571 B.n439 VSUBS 0.009938f
C572 B.n440 VSUBS 0.009938f
C573 B.n441 VSUBS 0.009938f
C574 B.n442 VSUBS 0.009938f
C575 B.n443 VSUBS 0.009938f
C576 B.n444 VSUBS 0.009938f
C577 B.n445 VSUBS 0.009938f
C578 B.n446 VSUBS 0.009938f
C579 B.n447 VSUBS 0.009938f
C580 B.n448 VSUBS 0.009938f
C581 B.n449 VSUBS 0.009938f
C582 B.n450 VSUBS 0.009938f
C583 B.n451 VSUBS 0.009938f
C584 B.n452 VSUBS 0.009938f
C585 B.n453 VSUBS 0.009938f
C586 B.n454 VSUBS 0.009938f
C587 B.n455 VSUBS 0.009938f
C588 B.n456 VSUBS 0.009938f
C589 B.n457 VSUBS 0.009938f
C590 B.n458 VSUBS 0.009938f
C591 B.n459 VSUBS 0.009938f
C592 B.n460 VSUBS 0.009938f
C593 B.n461 VSUBS 0.009938f
C594 B.n462 VSUBS 0.009938f
C595 B.n463 VSUBS 0.009938f
C596 B.n464 VSUBS 0.009938f
C597 B.n465 VSUBS 0.009938f
C598 B.n466 VSUBS 0.009938f
C599 B.n467 VSUBS 0.009938f
C600 B.n468 VSUBS 0.009938f
C601 B.n469 VSUBS 0.009938f
C602 B.n470 VSUBS 0.009938f
C603 B.n471 VSUBS 0.009938f
C604 B.n472 VSUBS 0.009938f
C605 B.n473 VSUBS 0.009938f
C606 B.n474 VSUBS 0.009938f
C607 B.n475 VSUBS 0.009938f
C608 B.n476 VSUBS 0.009938f
C609 B.n477 VSUBS 0.009938f
C610 B.n478 VSUBS 0.009938f
C611 B.n479 VSUBS 0.009938f
C612 B.n480 VSUBS 0.009938f
C613 B.n481 VSUBS 0.009938f
C614 B.n482 VSUBS 0.009938f
C615 B.n483 VSUBS 0.009938f
C616 B.n484 VSUBS 0.009938f
C617 B.n485 VSUBS 0.009938f
C618 B.n486 VSUBS 0.009938f
C619 B.n487 VSUBS 0.009938f
C620 B.n488 VSUBS 0.009938f
C621 B.n489 VSUBS 0.009938f
C622 B.n490 VSUBS 0.009938f
C623 B.n491 VSUBS 0.009938f
C624 B.n492 VSUBS 0.009938f
C625 B.n493 VSUBS 0.009938f
C626 B.n494 VSUBS 0.009938f
C627 B.n495 VSUBS 0.009938f
C628 B.n496 VSUBS 0.009938f
C629 B.n497 VSUBS 0.009938f
C630 B.n498 VSUBS 0.009938f
C631 B.n499 VSUBS 0.009938f
C632 B.n500 VSUBS 0.009938f
C633 B.n501 VSUBS 0.009938f
C634 B.n502 VSUBS 0.009938f
C635 B.n503 VSUBS 0.009938f
C636 B.n504 VSUBS 0.009938f
C637 B.n505 VSUBS 0.009938f
C638 B.n506 VSUBS 0.009938f
C639 B.n507 VSUBS 0.009938f
C640 B.n508 VSUBS 0.009938f
C641 B.n509 VSUBS 0.009938f
C642 B.n510 VSUBS 0.009938f
C643 B.n511 VSUBS 0.009938f
C644 B.n512 VSUBS 0.009938f
C645 B.n513 VSUBS 0.009938f
C646 B.n514 VSUBS 0.009938f
C647 B.n515 VSUBS 0.009938f
C648 B.n516 VSUBS 0.009938f
C649 B.n517 VSUBS 0.009938f
C650 B.n518 VSUBS 0.009938f
C651 B.n519 VSUBS 0.009938f
C652 B.n520 VSUBS 0.009938f
C653 B.n521 VSUBS 0.009938f
C654 B.n522 VSUBS 0.009938f
C655 B.n523 VSUBS 0.009938f
C656 B.n524 VSUBS 0.009938f
C657 B.n525 VSUBS 0.009938f
C658 B.n526 VSUBS 0.009938f
C659 B.n527 VSUBS 0.009938f
C660 B.n528 VSUBS 0.009938f
C661 B.n529 VSUBS 0.009938f
C662 B.n530 VSUBS 0.009938f
C663 B.n531 VSUBS 0.009938f
C664 B.n532 VSUBS 0.009938f
C665 B.n533 VSUBS 0.009938f
C666 B.n534 VSUBS 0.009938f
C667 B.n535 VSUBS 0.009938f
C668 B.n536 VSUBS 0.009938f
C669 B.n537 VSUBS 0.009938f
C670 B.n538 VSUBS 0.009938f
C671 B.n539 VSUBS 0.009938f
C672 B.n540 VSUBS 0.009938f
C673 B.n541 VSUBS 0.009938f
C674 B.n542 VSUBS 0.009938f
C675 B.n543 VSUBS 0.009938f
C676 B.n544 VSUBS 0.009938f
C677 B.n545 VSUBS 0.009938f
C678 B.n546 VSUBS 0.009938f
C679 B.n547 VSUBS 0.009938f
C680 B.n548 VSUBS 0.009938f
C681 B.n549 VSUBS 0.009938f
C682 B.n550 VSUBS 0.009938f
C683 B.n551 VSUBS 0.009938f
C684 B.n552 VSUBS 0.009938f
C685 B.n553 VSUBS 0.009938f
C686 B.n554 VSUBS 0.009938f
C687 B.n555 VSUBS 0.02192f
C688 B.n556 VSUBS 0.023167f
C689 B.n557 VSUBS 0.021555f
C690 B.n558 VSUBS 0.009938f
C691 B.n559 VSUBS 0.009938f
C692 B.n560 VSUBS 0.009938f
C693 B.n561 VSUBS 0.009938f
C694 B.n562 VSUBS 0.009938f
C695 B.n563 VSUBS 0.009938f
C696 B.n564 VSUBS 0.009938f
C697 B.n565 VSUBS 0.009938f
C698 B.n566 VSUBS 0.009938f
C699 B.n567 VSUBS 0.009938f
C700 B.n568 VSUBS 0.009938f
C701 B.n569 VSUBS 0.009938f
C702 B.n570 VSUBS 0.009938f
C703 B.n571 VSUBS 0.009938f
C704 B.n572 VSUBS 0.009938f
C705 B.n573 VSUBS 0.009938f
C706 B.n574 VSUBS 0.009938f
C707 B.n575 VSUBS 0.009938f
C708 B.n576 VSUBS 0.009938f
C709 B.n577 VSUBS 0.009938f
C710 B.n578 VSUBS 0.009938f
C711 B.n579 VSUBS 0.009938f
C712 B.n580 VSUBS 0.009938f
C713 B.n581 VSUBS 0.009938f
C714 B.n582 VSUBS 0.009938f
C715 B.n583 VSUBS 0.009938f
C716 B.n584 VSUBS 0.009938f
C717 B.n585 VSUBS 0.009938f
C718 B.n586 VSUBS 0.009938f
C719 B.n587 VSUBS 0.006869f
C720 B.n588 VSUBS 0.023026f
C721 B.n589 VSUBS 0.008038f
C722 B.n590 VSUBS 0.009938f
C723 B.n591 VSUBS 0.009938f
C724 B.n592 VSUBS 0.009938f
C725 B.n593 VSUBS 0.009938f
C726 B.n594 VSUBS 0.009938f
C727 B.n595 VSUBS 0.009938f
C728 B.n596 VSUBS 0.009938f
C729 B.n597 VSUBS 0.009938f
C730 B.n598 VSUBS 0.009938f
C731 B.n599 VSUBS 0.009938f
C732 B.n600 VSUBS 0.009938f
C733 B.n601 VSUBS 0.008038f
C734 B.n602 VSUBS 0.009938f
C735 B.n603 VSUBS 0.009938f
C736 B.n604 VSUBS 0.009938f
C737 B.n605 VSUBS 0.009938f
C738 B.n606 VSUBS 0.009938f
C739 B.n607 VSUBS 0.009938f
C740 B.n608 VSUBS 0.009938f
C741 B.n609 VSUBS 0.009938f
C742 B.n610 VSUBS 0.009938f
C743 B.n611 VSUBS 0.009938f
C744 B.n612 VSUBS 0.009938f
C745 B.n613 VSUBS 0.009938f
C746 B.n614 VSUBS 0.009938f
C747 B.n615 VSUBS 0.009938f
C748 B.n616 VSUBS 0.009938f
C749 B.n617 VSUBS 0.009938f
C750 B.n618 VSUBS 0.009938f
C751 B.n619 VSUBS 0.009938f
C752 B.n620 VSUBS 0.009938f
C753 B.n621 VSUBS 0.009938f
C754 B.n622 VSUBS 0.009938f
C755 B.n623 VSUBS 0.009938f
C756 B.n624 VSUBS 0.009938f
C757 B.n625 VSUBS 0.009938f
C758 B.n626 VSUBS 0.009938f
C759 B.n627 VSUBS 0.009938f
C760 B.n628 VSUBS 0.009938f
C761 B.n629 VSUBS 0.009938f
C762 B.n630 VSUBS 0.009938f
C763 B.n631 VSUBS 0.009938f
C764 B.n632 VSUBS 0.009938f
C765 B.n633 VSUBS 0.022802f
C766 B.n634 VSUBS 0.02192f
C767 B.n635 VSUBS 0.02192f
C768 B.n636 VSUBS 0.009938f
C769 B.n637 VSUBS 0.009938f
C770 B.n638 VSUBS 0.009938f
C771 B.n639 VSUBS 0.009938f
C772 B.n640 VSUBS 0.009938f
C773 B.n641 VSUBS 0.009938f
C774 B.n642 VSUBS 0.009938f
C775 B.n643 VSUBS 0.009938f
C776 B.n644 VSUBS 0.009938f
C777 B.n645 VSUBS 0.009938f
C778 B.n646 VSUBS 0.009938f
C779 B.n647 VSUBS 0.009938f
C780 B.n648 VSUBS 0.009938f
C781 B.n649 VSUBS 0.009938f
C782 B.n650 VSUBS 0.009938f
C783 B.n651 VSUBS 0.009938f
C784 B.n652 VSUBS 0.009938f
C785 B.n653 VSUBS 0.009938f
C786 B.n654 VSUBS 0.009938f
C787 B.n655 VSUBS 0.009938f
C788 B.n656 VSUBS 0.009938f
C789 B.n657 VSUBS 0.009938f
C790 B.n658 VSUBS 0.009938f
C791 B.n659 VSUBS 0.009938f
C792 B.n660 VSUBS 0.009938f
C793 B.n661 VSUBS 0.009938f
C794 B.n662 VSUBS 0.009938f
C795 B.n663 VSUBS 0.009938f
C796 B.n664 VSUBS 0.009938f
C797 B.n665 VSUBS 0.009938f
C798 B.n666 VSUBS 0.009938f
C799 B.n667 VSUBS 0.009938f
C800 B.n668 VSUBS 0.009938f
C801 B.n669 VSUBS 0.009938f
C802 B.n670 VSUBS 0.009938f
C803 B.n671 VSUBS 0.009938f
C804 B.n672 VSUBS 0.009938f
C805 B.n673 VSUBS 0.009938f
C806 B.n674 VSUBS 0.009938f
C807 B.n675 VSUBS 0.009938f
C808 B.n676 VSUBS 0.009938f
C809 B.n677 VSUBS 0.009938f
C810 B.n678 VSUBS 0.009938f
C811 B.n679 VSUBS 0.009938f
C812 B.n680 VSUBS 0.009938f
C813 B.n681 VSUBS 0.009938f
C814 B.n682 VSUBS 0.009938f
C815 B.n683 VSUBS 0.009938f
C816 B.n684 VSUBS 0.009938f
C817 B.n685 VSUBS 0.009938f
C818 B.n686 VSUBS 0.009938f
C819 B.n687 VSUBS 0.009938f
C820 B.n688 VSUBS 0.009938f
C821 B.n689 VSUBS 0.009938f
C822 B.n690 VSUBS 0.009938f
C823 B.n691 VSUBS 0.009938f
C824 B.n692 VSUBS 0.009938f
C825 B.n693 VSUBS 0.009938f
C826 B.n694 VSUBS 0.009938f
C827 B.n695 VSUBS 0.009938f
C828 B.n696 VSUBS 0.009938f
C829 B.n697 VSUBS 0.009938f
C830 B.n698 VSUBS 0.009938f
C831 B.n699 VSUBS 0.009938f
C832 B.n700 VSUBS 0.009938f
C833 B.n701 VSUBS 0.009938f
C834 B.n702 VSUBS 0.009938f
C835 B.n703 VSUBS 0.009938f
C836 B.n704 VSUBS 0.009938f
C837 B.n705 VSUBS 0.009938f
C838 B.n706 VSUBS 0.009938f
C839 B.n707 VSUBS 0.009938f
C840 B.n708 VSUBS 0.009938f
C841 B.n709 VSUBS 0.009938f
C842 B.n710 VSUBS 0.009938f
C843 B.n711 VSUBS 0.009938f
C844 B.n712 VSUBS 0.009938f
C845 B.n713 VSUBS 0.009938f
C846 B.n714 VSUBS 0.009938f
C847 B.n715 VSUBS 0.009938f
C848 B.n716 VSUBS 0.009938f
C849 B.n717 VSUBS 0.009938f
C850 B.n718 VSUBS 0.009938f
C851 B.n719 VSUBS 0.009938f
C852 B.n720 VSUBS 0.009938f
C853 B.n721 VSUBS 0.009938f
C854 B.n722 VSUBS 0.009938f
C855 B.n723 VSUBS 0.009938f
C856 B.n724 VSUBS 0.009938f
C857 B.n725 VSUBS 0.009938f
C858 B.n726 VSUBS 0.009938f
C859 B.n727 VSUBS 0.009938f
C860 B.n728 VSUBS 0.009938f
C861 B.n729 VSUBS 0.009938f
C862 B.n730 VSUBS 0.009938f
C863 B.n731 VSUBS 0.022504f
C864 VTAIL.t0 VSUBS 0.124645f
C865 VTAIL.t6 VSUBS 0.124645f
C866 VTAIL.n0 VSUBS 0.679699f
C867 VTAIL.n1 VSUBS 0.890187f
C868 VTAIL.t2 VSUBS 0.953409f
C869 VTAIL.n2 VSUBS 0.999203f
C870 VTAIL.t8 VSUBS 0.953409f
C871 VTAIL.n3 VSUBS 0.999203f
C872 VTAIL.t14 VSUBS 0.124645f
C873 VTAIL.t13 VSUBS 0.124645f
C874 VTAIL.n4 VSUBS 0.679699f
C875 VTAIL.n5 VSUBS 1.22373f
C876 VTAIL.t15 VSUBS 0.953409f
C877 VTAIL.n6 VSUBS 2.16626f
C878 VTAIL.t4 VSUBS 0.953415f
C879 VTAIL.n7 VSUBS 2.16626f
C880 VTAIL.t1 VSUBS 0.124645f
C881 VTAIL.t7 VSUBS 0.124645f
C882 VTAIL.n8 VSUBS 0.679703f
C883 VTAIL.n9 VSUBS 1.22372f
C884 VTAIL.t5 VSUBS 0.953415f
C885 VTAIL.n10 VSUBS 0.999197f
C886 VTAIL.t10 VSUBS 0.953415f
C887 VTAIL.n11 VSUBS 0.999197f
C888 VTAIL.t12 VSUBS 0.124645f
C889 VTAIL.t11 VSUBS 0.124645f
C890 VTAIL.n12 VSUBS 0.679703f
C891 VTAIL.n13 VSUBS 1.22372f
C892 VTAIL.t9 VSUBS 0.953409f
C893 VTAIL.n14 VSUBS 2.16626f
C894 VTAIL.t3 VSUBS 0.953409f
C895 VTAIL.n15 VSUBS 2.16022f
C896 VDD1.t3 VSUBS 0.132837f
C897 VDD1.t1 VSUBS 0.132837f
C898 VDD1.n0 VSUBS 0.846115f
C899 VDD1.t7 VSUBS 0.132837f
C900 VDD1.t6 VSUBS 0.132837f
C901 VDD1.n1 VSUBS 0.844728f
C902 VDD1.t5 VSUBS 0.132837f
C903 VDD1.t2 VSUBS 0.132837f
C904 VDD1.n2 VSUBS 0.844728f
C905 VDD1.n3 VSUBS 5.14408f
C906 VDD1.t0 VSUBS 0.132837f
C907 VDD1.t4 VSUBS 0.132837f
C908 VDD1.n4 VSUBS 0.828009f
C909 VDD1.n5 VSUBS 3.99928f
C910 VP.t7 VSUBS 1.77033f
C911 VP.n0 VSUBS 0.820905f
C912 VP.n1 VSUBS 0.040067f
C913 VP.n2 VSUBS 0.054025f
C914 VP.n3 VSUBS 0.040067f
C915 VP.n4 VSUBS 0.045548f
C916 VP.n5 VSUBS 0.040067f
C917 VP.n6 VSUBS 0.032391f
C918 VP.n7 VSUBS 0.040067f
C919 VP.t1 VSUBS 1.77033f
C920 VP.n8 VSUBS 0.670142f
C921 VP.n9 VSUBS 0.040067f
C922 VP.n10 VSUBS 0.062957f
C923 VP.n11 VSUBS 0.040067f
C924 VP.n12 VSUBS 0.051447f
C925 VP.t6 VSUBS 1.77033f
C926 VP.n13 VSUBS 0.820905f
C927 VP.n14 VSUBS 0.040067f
C928 VP.n15 VSUBS 0.054025f
C929 VP.n16 VSUBS 0.040067f
C930 VP.n17 VSUBS 0.045548f
C931 VP.n18 VSUBS 0.040067f
C932 VP.n19 VSUBS 0.032391f
C933 VP.n20 VSUBS 0.040067f
C934 VP.t3 VSUBS 1.77033f
C935 VP.n21 VSUBS 0.818994f
C936 VP.t5 VSUBS 2.24816f
C937 VP.n22 VSUBS 0.78597f
C938 VP.n23 VSUBS 0.493841f
C939 VP.n24 VSUBS 0.066931f
C940 VP.n25 VSUBS 0.074675f
C941 VP.n26 VSUBS 0.079633f
C942 VP.n27 VSUBS 0.040067f
C943 VP.n28 VSUBS 0.040067f
C944 VP.n29 VSUBS 0.040067f
C945 VP.n30 VSUBS 0.079633f
C946 VP.n31 VSUBS 0.074675f
C947 VP.t4 VSUBS 1.77033f
C948 VP.n32 VSUBS 0.670142f
C949 VP.n33 VSUBS 0.066931f
C950 VP.n34 VSUBS 0.040067f
C951 VP.n35 VSUBS 0.040067f
C952 VP.n36 VSUBS 0.040067f
C953 VP.n37 VSUBS 0.074675f
C954 VP.n38 VSUBS 0.074675f
C955 VP.n39 VSUBS 0.062957f
C956 VP.n40 VSUBS 0.040067f
C957 VP.n41 VSUBS 0.040067f
C958 VP.n42 VSUBS 0.040067f
C959 VP.n43 VSUBS 0.074675f
C960 VP.n44 VSUBS 0.074675f
C961 VP.n45 VSUBS 0.051447f
C962 VP.n46 VSUBS 0.064668f
C963 VP.n47 VSUBS 2.26339f
C964 VP.t0 VSUBS 1.77033f
C965 VP.n48 VSUBS 0.820905f
C966 VP.n49 VSUBS 2.29242f
C967 VP.n50 VSUBS 0.064668f
C968 VP.n51 VSUBS 0.040067f
C969 VP.n52 VSUBS 0.074675f
C970 VP.n53 VSUBS 0.074675f
C971 VP.n54 VSUBS 0.054025f
C972 VP.n55 VSUBS 0.040067f
C973 VP.n56 VSUBS 0.040067f
C974 VP.n57 VSUBS 0.040067f
C975 VP.n58 VSUBS 0.074675f
C976 VP.n59 VSUBS 0.074675f
C977 VP.n60 VSUBS 0.045548f
C978 VP.n61 VSUBS 0.040067f
C979 VP.n62 VSUBS 0.040067f
C980 VP.n63 VSUBS 0.066931f
C981 VP.n64 VSUBS 0.074675f
C982 VP.n65 VSUBS 0.079633f
C983 VP.n66 VSUBS 0.040067f
C984 VP.n67 VSUBS 0.040067f
C985 VP.n68 VSUBS 0.040067f
C986 VP.n69 VSUBS 0.079633f
C987 VP.n70 VSUBS 0.074675f
C988 VP.t2 VSUBS 1.77033f
C989 VP.n71 VSUBS 0.670142f
C990 VP.n72 VSUBS 0.066931f
C991 VP.n73 VSUBS 0.040067f
C992 VP.n74 VSUBS 0.040067f
C993 VP.n75 VSUBS 0.040067f
C994 VP.n76 VSUBS 0.074675f
C995 VP.n77 VSUBS 0.074675f
C996 VP.n78 VSUBS 0.062957f
C997 VP.n79 VSUBS 0.040067f
C998 VP.n80 VSUBS 0.040067f
C999 VP.n81 VSUBS 0.040067f
C1000 VP.n82 VSUBS 0.074675f
C1001 VP.n83 VSUBS 0.074675f
C1002 VP.n84 VSUBS 0.051447f
C1003 VP.n85 VSUBS 0.064668f
C1004 VP.n86 VSUBS 0.108158f
.ends

