* NGSPICE file created from diff_pair_sample_0283.ext - technology: sky130A

.subckt diff_pair_sample_0283 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=1.2519 ps=7.2 w=3.21 l=0.48
X1 B.t11 B.t9 B.t10 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=0 ps=0 w=3.21 l=0.48
X2 B.t8 B.t6 B.t7 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=0 ps=0 w=3.21 l=0.48
X3 B.t5 B.t3 B.t4 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=0 ps=0 w=3.21 l=0.48
X4 VDD2.t1 VN.t0 VTAIL.t3 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=1.2519 ps=7.2 w=3.21 l=0.48
X5 VDD1.t0 VP.t1 VTAIL.t1 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=1.2519 ps=7.2 w=3.21 l=0.48
X6 B.t2 B.t0 B.t1 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=0 ps=0 w=3.21 l=0.48
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1294_n1614# sky130_fd_pr__pfet_01v8 ad=1.2519 pd=7.2 as=1.2519 ps=7.2 w=3.21 l=0.48
R0 VP.n0 VP.t1 437.202
R1 VP.n0 VP.t0 404.81
R2 VP VP.n0 0.0516364
R3 VTAIL.n58 VTAIL.n48 756.745
R4 VTAIL.n10 VTAIL.n0 756.745
R5 VTAIL.n42 VTAIL.n32 756.745
R6 VTAIL.n26 VTAIL.n16 756.745
R7 VTAIL.n52 VTAIL.n51 585
R8 VTAIL.n57 VTAIL.n56 585
R9 VTAIL.n59 VTAIL.n58 585
R10 VTAIL.n4 VTAIL.n3 585
R11 VTAIL.n9 VTAIL.n8 585
R12 VTAIL.n11 VTAIL.n10 585
R13 VTAIL.n43 VTAIL.n42 585
R14 VTAIL.n41 VTAIL.n40 585
R15 VTAIL.n36 VTAIL.n35 585
R16 VTAIL.n27 VTAIL.n26 585
R17 VTAIL.n25 VTAIL.n24 585
R18 VTAIL.n20 VTAIL.n19 585
R19 VTAIL.n53 VTAIL.t3 336.901
R20 VTAIL.n5 VTAIL.t2 336.901
R21 VTAIL.n37 VTAIL.t1 336.901
R22 VTAIL.n21 VTAIL.t0 336.901
R23 VTAIL.n57 VTAIL.n51 171.744
R24 VTAIL.n58 VTAIL.n57 171.744
R25 VTAIL.n9 VTAIL.n3 171.744
R26 VTAIL.n10 VTAIL.n9 171.744
R27 VTAIL.n42 VTAIL.n41 171.744
R28 VTAIL.n41 VTAIL.n35 171.744
R29 VTAIL.n26 VTAIL.n25 171.744
R30 VTAIL.n25 VTAIL.n19 171.744
R31 VTAIL.t3 VTAIL.n51 85.8723
R32 VTAIL.t2 VTAIL.n3 85.8723
R33 VTAIL.t1 VTAIL.n35 85.8723
R34 VTAIL.t0 VTAIL.n19 85.8723
R35 VTAIL.n63 VTAIL.n62 33.9308
R36 VTAIL.n15 VTAIL.n14 33.9308
R37 VTAIL.n47 VTAIL.n46 33.9308
R38 VTAIL.n31 VTAIL.n30 33.9308
R39 VTAIL.n31 VTAIL.n15 16.5479
R40 VTAIL.n53 VTAIL.n52 16.193
R41 VTAIL.n5 VTAIL.n4 16.193
R42 VTAIL.n37 VTAIL.n36 16.193
R43 VTAIL.n21 VTAIL.n20 16.193
R44 VTAIL.n63 VTAIL.n47 15.8496
R45 VTAIL.n56 VTAIL.n55 12.8005
R46 VTAIL.n8 VTAIL.n7 12.8005
R47 VTAIL.n40 VTAIL.n39 12.8005
R48 VTAIL.n24 VTAIL.n23 12.8005
R49 VTAIL.n59 VTAIL.n50 12.0247
R50 VTAIL.n11 VTAIL.n2 12.0247
R51 VTAIL.n43 VTAIL.n34 12.0247
R52 VTAIL.n27 VTAIL.n18 12.0247
R53 VTAIL.n60 VTAIL.n48 11.249
R54 VTAIL.n12 VTAIL.n0 11.249
R55 VTAIL.n44 VTAIL.n32 11.249
R56 VTAIL.n28 VTAIL.n16 11.249
R57 VTAIL.n62 VTAIL.n61 9.45567
R58 VTAIL.n14 VTAIL.n13 9.45567
R59 VTAIL.n46 VTAIL.n45 9.45567
R60 VTAIL.n30 VTAIL.n29 9.45567
R61 VTAIL.n61 VTAIL.n60 9.3005
R62 VTAIL.n50 VTAIL.n49 9.3005
R63 VTAIL.n55 VTAIL.n54 9.3005
R64 VTAIL.n13 VTAIL.n12 9.3005
R65 VTAIL.n2 VTAIL.n1 9.3005
R66 VTAIL.n7 VTAIL.n6 9.3005
R67 VTAIL.n45 VTAIL.n44 9.3005
R68 VTAIL.n34 VTAIL.n33 9.3005
R69 VTAIL.n39 VTAIL.n38 9.3005
R70 VTAIL.n29 VTAIL.n28 9.3005
R71 VTAIL.n18 VTAIL.n17 9.3005
R72 VTAIL.n23 VTAIL.n22 9.3005
R73 VTAIL.n38 VTAIL.n37 3.91276
R74 VTAIL.n22 VTAIL.n21 3.91276
R75 VTAIL.n54 VTAIL.n53 3.91276
R76 VTAIL.n6 VTAIL.n5 3.91276
R77 VTAIL.n62 VTAIL.n48 2.71565
R78 VTAIL.n14 VTAIL.n0 2.71565
R79 VTAIL.n46 VTAIL.n32 2.71565
R80 VTAIL.n30 VTAIL.n16 2.71565
R81 VTAIL.n60 VTAIL.n59 1.93989
R82 VTAIL.n12 VTAIL.n11 1.93989
R83 VTAIL.n44 VTAIL.n43 1.93989
R84 VTAIL.n28 VTAIL.n27 1.93989
R85 VTAIL.n56 VTAIL.n50 1.16414
R86 VTAIL.n8 VTAIL.n2 1.16414
R87 VTAIL.n40 VTAIL.n34 1.16414
R88 VTAIL.n24 VTAIL.n18 1.16414
R89 VTAIL.n47 VTAIL.n31 0.819465
R90 VTAIL VTAIL.n15 0.703086
R91 VTAIL.n55 VTAIL.n52 0.388379
R92 VTAIL.n7 VTAIL.n4 0.388379
R93 VTAIL.n39 VTAIL.n36 0.388379
R94 VTAIL.n23 VTAIL.n20 0.388379
R95 VTAIL.n54 VTAIL.n49 0.155672
R96 VTAIL.n61 VTAIL.n49 0.155672
R97 VTAIL.n6 VTAIL.n1 0.155672
R98 VTAIL.n13 VTAIL.n1 0.155672
R99 VTAIL.n45 VTAIL.n33 0.155672
R100 VTAIL.n38 VTAIL.n33 0.155672
R101 VTAIL.n29 VTAIL.n17 0.155672
R102 VTAIL.n22 VTAIL.n17 0.155672
R103 VTAIL VTAIL.n63 0.116879
R104 VDD1.n10 VDD1.n0 756.745
R105 VDD1.n25 VDD1.n15 756.745
R106 VDD1.n11 VDD1.n10 585
R107 VDD1.n9 VDD1.n8 585
R108 VDD1.n4 VDD1.n3 585
R109 VDD1.n19 VDD1.n18 585
R110 VDD1.n24 VDD1.n23 585
R111 VDD1.n26 VDD1.n25 585
R112 VDD1.n5 VDD1.t0 336.901
R113 VDD1.n20 VDD1.t1 336.901
R114 VDD1.n10 VDD1.n9 171.744
R115 VDD1.n9 VDD1.n3 171.744
R116 VDD1.n24 VDD1.n18 171.744
R117 VDD1.n25 VDD1.n24 171.744
R118 VDD1.t0 VDD1.n3 85.8723
R119 VDD1.t1 VDD1.n18 85.8723
R120 VDD1 VDD1.n29 79.1495
R121 VDD1 VDD1.n14 50.8423
R122 VDD1.n5 VDD1.n4 16.193
R123 VDD1.n20 VDD1.n19 16.193
R124 VDD1.n8 VDD1.n7 12.8005
R125 VDD1.n23 VDD1.n22 12.8005
R126 VDD1.n11 VDD1.n2 12.0247
R127 VDD1.n26 VDD1.n17 12.0247
R128 VDD1.n12 VDD1.n0 11.249
R129 VDD1.n27 VDD1.n15 11.249
R130 VDD1.n14 VDD1.n13 9.45567
R131 VDD1.n29 VDD1.n28 9.45567
R132 VDD1.n13 VDD1.n12 9.3005
R133 VDD1.n2 VDD1.n1 9.3005
R134 VDD1.n7 VDD1.n6 9.3005
R135 VDD1.n28 VDD1.n27 9.3005
R136 VDD1.n17 VDD1.n16 9.3005
R137 VDD1.n22 VDD1.n21 9.3005
R138 VDD1.n6 VDD1.n5 3.91276
R139 VDD1.n21 VDD1.n20 3.91276
R140 VDD1.n14 VDD1.n0 2.71565
R141 VDD1.n29 VDD1.n15 2.71565
R142 VDD1.n12 VDD1.n11 1.93989
R143 VDD1.n27 VDD1.n26 1.93989
R144 VDD1.n8 VDD1.n2 1.16414
R145 VDD1.n23 VDD1.n17 1.16414
R146 VDD1.n7 VDD1.n4 0.388379
R147 VDD1.n22 VDD1.n19 0.388379
R148 VDD1.n13 VDD1.n1 0.155672
R149 VDD1.n6 VDD1.n1 0.155672
R150 VDD1.n21 VDD1.n16 0.155672
R151 VDD1.n28 VDD1.n16 0.155672
R152 B.n201 B.n200 585
R153 B.n202 B.n33 585
R154 B.n204 B.n203 585
R155 B.n205 B.n32 585
R156 B.n207 B.n206 585
R157 B.n208 B.n31 585
R158 B.n210 B.n209 585
R159 B.n211 B.n30 585
R160 B.n213 B.n212 585
R161 B.n214 B.n29 585
R162 B.n216 B.n215 585
R163 B.n217 B.n28 585
R164 B.n219 B.n218 585
R165 B.n220 B.n27 585
R166 B.n222 B.n221 585
R167 B.n223 B.n24 585
R168 B.n226 B.n225 585
R169 B.n227 B.n23 585
R170 B.n229 B.n228 585
R171 B.n230 B.n22 585
R172 B.n232 B.n231 585
R173 B.n233 B.n21 585
R174 B.n235 B.n234 585
R175 B.n236 B.n17 585
R176 B.n238 B.n237 585
R177 B.n239 B.n16 585
R178 B.n241 B.n240 585
R179 B.n242 B.n15 585
R180 B.n244 B.n243 585
R181 B.n245 B.n14 585
R182 B.n247 B.n246 585
R183 B.n248 B.n13 585
R184 B.n250 B.n249 585
R185 B.n251 B.n12 585
R186 B.n253 B.n252 585
R187 B.n254 B.n11 585
R188 B.n256 B.n255 585
R189 B.n257 B.n10 585
R190 B.n259 B.n258 585
R191 B.n260 B.n9 585
R192 B.n262 B.n261 585
R193 B.n199 B.n34 585
R194 B.n198 B.n197 585
R195 B.n196 B.n35 585
R196 B.n195 B.n194 585
R197 B.n193 B.n36 585
R198 B.n192 B.n191 585
R199 B.n190 B.n37 585
R200 B.n189 B.n188 585
R201 B.n187 B.n38 585
R202 B.n186 B.n185 585
R203 B.n184 B.n39 585
R204 B.n183 B.n182 585
R205 B.n181 B.n40 585
R206 B.n180 B.n179 585
R207 B.n178 B.n41 585
R208 B.n177 B.n176 585
R209 B.n175 B.n42 585
R210 B.n174 B.n173 585
R211 B.n172 B.n43 585
R212 B.n171 B.n170 585
R213 B.n169 B.n44 585
R214 B.n168 B.n167 585
R215 B.n166 B.n45 585
R216 B.n165 B.n164 585
R217 B.n163 B.n46 585
R218 B.n162 B.n161 585
R219 B.n160 B.n47 585
R220 B.n95 B.n94 585
R221 B.n96 B.n69 585
R222 B.n98 B.n97 585
R223 B.n99 B.n68 585
R224 B.n101 B.n100 585
R225 B.n102 B.n67 585
R226 B.n104 B.n103 585
R227 B.n105 B.n66 585
R228 B.n107 B.n106 585
R229 B.n108 B.n65 585
R230 B.n110 B.n109 585
R231 B.n111 B.n64 585
R232 B.n113 B.n112 585
R233 B.n114 B.n63 585
R234 B.n116 B.n115 585
R235 B.n117 B.n60 585
R236 B.n120 B.n119 585
R237 B.n121 B.n59 585
R238 B.n123 B.n122 585
R239 B.n124 B.n58 585
R240 B.n126 B.n125 585
R241 B.n127 B.n57 585
R242 B.n129 B.n128 585
R243 B.n130 B.n56 585
R244 B.n135 B.n134 585
R245 B.n136 B.n55 585
R246 B.n138 B.n137 585
R247 B.n139 B.n54 585
R248 B.n141 B.n140 585
R249 B.n142 B.n53 585
R250 B.n144 B.n143 585
R251 B.n145 B.n52 585
R252 B.n147 B.n146 585
R253 B.n148 B.n51 585
R254 B.n150 B.n149 585
R255 B.n151 B.n50 585
R256 B.n153 B.n152 585
R257 B.n154 B.n49 585
R258 B.n156 B.n155 585
R259 B.n157 B.n48 585
R260 B.n159 B.n158 585
R261 B.n93 B.n70 585
R262 B.n92 B.n91 585
R263 B.n90 B.n71 585
R264 B.n89 B.n88 585
R265 B.n87 B.n72 585
R266 B.n86 B.n85 585
R267 B.n84 B.n73 585
R268 B.n83 B.n82 585
R269 B.n81 B.n74 585
R270 B.n80 B.n79 585
R271 B.n78 B.n75 585
R272 B.n77 B.n76 585
R273 B.n2 B.n0 585
R274 B.n281 B.n1 585
R275 B.n280 B.n279 585
R276 B.n278 B.n3 585
R277 B.n277 B.n276 585
R278 B.n275 B.n4 585
R279 B.n274 B.n273 585
R280 B.n272 B.n5 585
R281 B.n271 B.n270 585
R282 B.n269 B.n6 585
R283 B.n268 B.n267 585
R284 B.n266 B.n7 585
R285 B.n265 B.n264 585
R286 B.n263 B.n8 585
R287 B.n283 B.n282 585
R288 B.n95 B.n70 497.305
R289 B.n263 B.n262 497.305
R290 B.n160 B.n159 497.305
R291 B.n201 B.n34 497.305
R292 B.n131 B.t3 368.079
R293 B.n61 B.t6 368.079
R294 B.n18 B.t9 368.079
R295 B.n25 B.t0 368.079
R296 B.n131 B.t5 241.464
R297 B.n25 B.t1 241.464
R298 B.n61 B.t8 241.464
R299 B.n18 B.t10 241.464
R300 B.n132 B.t4 225.755
R301 B.n26 B.t2 225.755
R302 B.n62 B.t7 225.755
R303 B.n19 B.t11 225.755
R304 B.n91 B.n70 163.367
R305 B.n91 B.n90 163.367
R306 B.n90 B.n89 163.367
R307 B.n89 B.n72 163.367
R308 B.n85 B.n72 163.367
R309 B.n85 B.n84 163.367
R310 B.n84 B.n83 163.367
R311 B.n83 B.n74 163.367
R312 B.n79 B.n74 163.367
R313 B.n79 B.n78 163.367
R314 B.n78 B.n77 163.367
R315 B.n77 B.n2 163.367
R316 B.n282 B.n2 163.367
R317 B.n282 B.n281 163.367
R318 B.n281 B.n280 163.367
R319 B.n280 B.n3 163.367
R320 B.n276 B.n3 163.367
R321 B.n276 B.n275 163.367
R322 B.n275 B.n274 163.367
R323 B.n274 B.n5 163.367
R324 B.n270 B.n5 163.367
R325 B.n270 B.n269 163.367
R326 B.n269 B.n268 163.367
R327 B.n268 B.n7 163.367
R328 B.n264 B.n7 163.367
R329 B.n264 B.n263 163.367
R330 B.n96 B.n95 163.367
R331 B.n97 B.n96 163.367
R332 B.n97 B.n68 163.367
R333 B.n101 B.n68 163.367
R334 B.n102 B.n101 163.367
R335 B.n103 B.n102 163.367
R336 B.n103 B.n66 163.367
R337 B.n107 B.n66 163.367
R338 B.n108 B.n107 163.367
R339 B.n109 B.n108 163.367
R340 B.n109 B.n64 163.367
R341 B.n113 B.n64 163.367
R342 B.n114 B.n113 163.367
R343 B.n115 B.n114 163.367
R344 B.n115 B.n60 163.367
R345 B.n120 B.n60 163.367
R346 B.n121 B.n120 163.367
R347 B.n122 B.n121 163.367
R348 B.n122 B.n58 163.367
R349 B.n126 B.n58 163.367
R350 B.n127 B.n126 163.367
R351 B.n128 B.n127 163.367
R352 B.n128 B.n56 163.367
R353 B.n135 B.n56 163.367
R354 B.n136 B.n135 163.367
R355 B.n137 B.n136 163.367
R356 B.n137 B.n54 163.367
R357 B.n141 B.n54 163.367
R358 B.n142 B.n141 163.367
R359 B.n143 B.n142 163.367
R360 B.n143 B.n52 163.367
R361 B.n147 B.n52 163.367
R362 B.n148 B.n147 163.367
R363 B.n149 B.n148 163.367
R364 B.n149 B.n50 163.367
R365 B.n153 B.n50 163.367
R366 B.n154 B.n153 163.367
R367 B.n155 B.n154 163.367
R368 B.n155 B.n48 163.367
R369 B.n159 B.n48 163.367
R370 B.n161 B.n160 163.367
R371 B.n161 B.n46 163.367
R372 B.n165 B.n46 163.367
R373 B.n166 B.n165 163.367
R374 B.n167 B.n166 163.367
R375 B.n167 B.n44 163.367
R376 B.n171 B.n44 163.367
R377 B.n172 B.n171 163.367
R378 B.n173 B.n172 163.367
R379 B.n173 B.n42 163.367
R380 B.n177 B.n42 163.367
R381 B.n178 B.n177 163.367
R382 B.n179 B.n178 163.367
R383 B.n179 B.n40 163.367
R384 B.n183 B.n40 163.367
R385 B.n184 B.n183 163.367
R386 B.n185 B.n184 163.367
R387 B.n185 B.n38 163.367
R388 B.n189 B.n38 163.367
R389 B.n190 B.n189 163.367
R390 B.n191 B.n190 163.367
R391 B.n191 B.n36 163.367
R392 B.n195 B.n36 163.367
R393 B.n196 B.n195 163.367
R394 B.n197 B.n196 163.367
R395 B.n197 B.n34 163.367
R396 B.n262 B.n9 163.367
R397 B.n258 B.n9 163.367
R398 B.n258 B.n257 163.367
R399 B.n257 B.n256 163.367
R400 B.n256 B.n11 163.367
R401 B.n252 B.n11 163.367
R402 B.n252 B.n251 163.367
R403 B.n251 B.n250 163.367
R404 B.n250 B.n13 163.367
R405 B.n246 B.n13 163.367
R406 B.n246 B.n245 163.367
R407 B.n245 B.n244 163.367
R408 B.n244 B.n15 163.367
R409 B.n240 B.n15 163.367
R410 B.n240 B.n239 163.367
R411 B.n239 B.n238 163.367
R412 B.n238 B.n17 163.367
R413 B.n234 B.n17 163.367
R414 B.n234 B.n233 163.367
R415 B.n233 B.n232 163.367
R416 B.n232 B.n22 163.367
R417 B.n228 B.n22 163.367
R418 B.n228 B.n227 163.367
R419 B.n227 B.n226 163.367
R420 B.n226 B.n24 163.367
R421 B.n221 B.n24 163.367
R422 B.n221 B.n220 163.367
R423 B.n220 B.n219 163.367
R424 B.n219 B.n28 163.367
R425 B.n215 B.n28 163.367
R426 B.n215 B.n214 163.367
R427 B.n214 B.n213 163.367
R428 B.n213 B.n30 163.367
R429 B.n209 B.n30 163.367
R430 B.n209 B.n208 163.367
R431 B.n208 B.n207 163.367
R432 B.n207 B.n32 163.367
R433 B.n203 B.n32 163.367
R434 B.n203 B.n202 163.367
R435 B.n202 B.n201 163.367
R436 B.n133 B.n132 59.5399
R437 B.n118 B.n62 59.5399
R438 B.n20 B.n19 59.5399
R439 B.n224 B.n26 59.5399
R440 B.n261 B.n8 32.3127
R441 B.n200 B.n199 32.3127
R442 B.n158 B.n47 32.3127
R443 B.n94 B.n93 32.3127
R444 B B.n283 18.0485
R445 B.n132 B.n131 15.7096
R446 B.n62 B.n61 15.7096
R447 B.n19 B.n18 15.7096
R448 B.n26 B.n25 15.7096
R449 B.n261 B.n260 10.6151
R450 B.n260 B.n259 10.6151
R451 B.n259 B.n10 10.6151
R452 B.n255 B.n10 10.6151
R453 B.n255 B.n254 10.6151
R454 B.n254 B.n253 10.6151
R455 B.n253 B.n12 10.6151
R456 B.n249 B.n12 10.6151
R457 B.n249 B.n248 10.6151
R458 B.n248 B.n247 10.6151
R459 B.n247 B.n14 10.6151
R460 B.n243 B.n14 10.6151
R461 B.n243 B.n242 10.6151
R462 B.n242 B.n241 10.6151
R463 B.n241 B.n16 10.6151
R464 B.n237 B.n236 10.6151
R465 B.n236 B.n235 10.6151
R466 B.n235 B.n21 10.6151
R467 B.n231 B.n21 10.6151
R468 B.n231 B.n230 10.6151
R469 B.n230 B.n229 10.6151
R470 B.n229 B.n23 10.6151
R471 B.n225 B.n23 10.6151
R472 B.n223 B.n222 10.6151
R473 B.n222 B.n27 10.6151
R474 B.n218 B.n27 10.6151
R475 B.n218 B.n217 10.6151
R476 B.n217 B.n216 10.6151
R477 B.n216 B.n29 10.6151
R478 B.n212 B.n29 10.6151
R479 B.n212 B.n211 10.6151
R480 B.n211 B.n210 10.6151
R481 B.n210 B.n31 10.6151
R482 B.n206 B.n31 10.6151
R483 B.n206 B.n205 10.6151
R484 B.n205 B.n204 10.6151
R485 B.n204 B.n33 10.6151
R486 B.n200 B.n33 10.6151
R487 B.n162 B.n47 10.6151
R488 B.n163 B.n162 10.6151
R489 B.n164 B.n163 10.6151
R490 B.n164 B.n45 10.6151
R491 B.n168 B.n45 10.6151
R492 B.n169 B.n168 10.6151
R493 B.n170 B.n169 10.6151
R494 B.n170 B.n43 10.6151
R495 B.n174 B.n43 10.6151
R496 B.n175 B.n174 10.6151
R497 B.n176 B.n175 10.6151
R498 B.n176 B.n41 10.6151
R499 B.n180 B.n41 10.6151
R500 B.n181 B.n180 10.6151
R501 B.n182 B.n181 10.6151
R502 B.n182 B.n39 10.6151
R503 B.n186 B.n39 10.6151
R504 B.n187 B.n186 10.6151
R505 B.n188 B.n187 10.6151
R506 B.n188 B.n37 10.6151
R507 B.n192 B.n37 10.6151
R508 B.n193 B.n192 10.6151
R509 B.n194 B.n193 10.6151
R510 B.n194 B.n35 10.6151
R511 B.n198 B.n35 10.6151
R512 B.n199 B.n198 10.6151
R513 B.n94 B.n69 10.6151
R514 B.n98 B.n69 10.6151
R515 B.n99 B.n98 10.6151
R516 B.n100 B.n99 10.6151
R517 B.n100 B.n67 10.6151
R518 B.n104 B.n67 10.6151
R519 B.n105 B.n104 10.6151
R520 B.n106 B.n105 10.6151
R521 B.n106 B.n65 10.6151
R522 B.n110 B.n65 10.6151
R523 B.n111 B.n110 10.6151
R524 B.n112 B.n111 10.6151
R525 B.n112 B.n63 10.6151
R526 B.n116 B.n63 10.6151
R527 B.n117 B.n116 10.6151
R528 B.n119 B.n59 10.6151
R529 B.n123 B.n59 10.6151
R530 B.n124 B.n123 10.6151
R531 B.n125 B.n124 10.6151
R532 B.n125 B.n57 10.6151
R533 B.n129 B.n57 10.6151
R534 B.n130 B.n129 10.6151
R535 B.n134 B.n130 10.6151
R536 B.n138 B.n55 10.6151
R537 B.n139 B.n138 10.6151
R538 B.n140 B.n139 10.6151
R539 B.n140 B.n53 10.6151
R540 B.n144 B.n53 10.6151
R541 B.n145 B.n144 10.6151
R542 B.n146 B.n145 10.6151
R543 B.n146 B.n51 10.6151
R544 B.n150 B.n51 10.6151
R545 B.n151 B.n150 10.6151
R546 B.n152 B.n151 10.6151
R547 B.n152 B.n49 10.6151
R548 B.n156 B.n49 10.6151
R549 B.n157 B.n156 10.6151
R550 B.n158 B.n157 10.6151
R551 B.n93 B.n92 10.6151
R552 B.n92 B.n71 10.6151
R553 B.n88 B.n71 10.6151
R554 B.n88 B.n87 10.6151
R555 B.n87 B.n86 10.6151
R556 B.n86 B.n73 10.6151
R557 B.n82 B.n73 10.6151
R558 B.n82 B.n81 10.6151
R559 B.n81 B.n80 10.6151
R560 B.n80 B.n75 10.6151
R561 B.n76 B.n75 10.6151
R562 B.n76 B.n0 10.6151
R563 B.n279 B.n1 10.6151
R564 B.n279 B.n278 10.6151
R565 B.n278 B.n277 10.6151
R566 B.n277 B.n4 10.6151
R567 B.n273 B.n4 10.6151
R568 B.n273 B.n272 10.6151
R569 B.n272 B.n271 10.6151
R570 B.n271 B.n6 10.6151
R571 B.n267 B.n6 10.6151
R572 B.n267 B.n266 10.6151
R573 B.n266 B.n265 10.6151
R574 B.n265 B.n8 10.6151
R575 B.n237 B.n20 7.18099
R576 B.n225 B.n224 7.18099
R577 B.n119 B.n118 7.18099
R578 B.n134 B.n133 7.18099
R579 B.n20 B.n16 3.43465
R580 B.n224 B.n223 3.43465
R581 B.n118 B.n117 3.43465
R582 B.n133 B.n55 3.43465
R583 B.n283 B.n0 2.81026
R584 B.n283 B.n1 2.81026
R585 VN VN.t1 437.582
R586 VN VN.t0 404.863
R587 VDD2.n25 VDD2.n15 756.745
R588 VDD2.n10 VDD2.n0 756.745
R589 VDD2.n26 VDD2.n25 585
R590 VDD2.n24 VDD2.n23 585
R591 VDD2.n19 VDD2.n18 585
R592 VDD2.n4 VDD2.n3 585
R593 VDD2.n9 VDD2.n8 585
R594 VDD2.n11 VDD2.n10 585
R595 VDD2.n20 VDD2.t0 336.901
R596 VDD2.n5 VDD2.t1 336.901
R597 VDD2.n25 VDD2.n24 171.744
R598 VDD2.n24 VDD2.n18 171.744
R599 VDD2.n9 VDD2.n3 171.744
R600 VDD2.n10 VDD2.n9 171.744
R601 VDD2.t0 VDD2.n18 85.8723
R602 VDD2.t1 VDD2.n3 85.8723
R603 VDD2.n30 VDD2.n14 78.4501
R604 VDD2.n30 VDD2.n29 50.6096
R605 VDD2.n20 VDD2.n19 16.193
R606 VDD2.n5 VDD2.n4 16.193
R607 VDD2.n23 VDD2.n22 12.8005
R608 VDD2.n8 VDD2.n7 12.8005
R609 VDD2.n26 VDD2.n17 12.0247
R610 VDD2.n11 VDD2.n2 12.0247
R611 VDD2.n27 VDD2.n15 11.249
R612 VDD2.n12 VDD2.n0 11.249
R613 VDD2.n29 VDD2.n28 9.45567
R614 VDD2.n14 VDD2.n13 9.45567
R615 VDD2.n28 VDD2.n27 9.3005
R616 VDD2.n17 VDD2.n16 9.3005
R617 VDD2.n22 VDD2.n21 9.3005
R618 VDD2.n13 VDD2.n12 9.3005
R619 VDD2.n2 VDD2.n1 9.3005
R620 VDD2.n7 VDD2.n6 9.3005
R621 VDD2.n21 VDD2.n20 3.91276
R622 VDD2.n6 VDD2.n5 3.91276
R623 VDD2.n29 VDD2.n15 2.71565
R624 VDD2.n14 VDD2.n0 2.71565
R625 VDD2.n27 VDD2.n26 1.93989
R626 VDD2.n12 VDD2.n11 1.93989
R627 VDD2.n23 VDD2.n17 1.16414
R628 VDD2.n8 VDD2.n2 1.16414
R629 VDD2.n22 VDD2.n19 0.388379
R630 VDD2.n7 VDD2.n4 0.388379
R631 VDD2 VDD2.n30 0.233259
R632 VDD2.n28 VDD2.n16 0.155672
R633 VDD2.n21 VDD2.n16 0.155672
R634 VDD2.n6 VDD2.n1 0.155672
R635 VDD2.n13 VDD2.n1 0.155672
C0 VTAIL VP 0.563512f
C1 VDD1 VP 0.727167f
C2 VN VP 2.8406f
C3 B VP 0.834456f
C4 VTAIL VDD1 2.49702f
C5 VTAIL VN 0.54925f
C6 VDD2 VP 0.249711f
C7 VN VDD1 0.153361f
C8 B VTAIL 1.03988f
C9 B VDD1 0.7454f
C10 B VN 0.579858f
C11 w_n1294_n1614# VP 1.58817f
C12 VTAIL VDD2 2.53401f
C13 VDD2 VDD1 0.439122f
C14 VDD2 VN 0.632628f
C15 w_n1294_n1614# VTAIL 1.43827f
C16 B VDD2 0.758508f
C17 w_n1294_n1614# VDD1 0.889606f
C18 w_n1294_n1614# VN 1.42991f
C19 w_n1294_n1614# B 4.04597f
C20 w_n1294_n1614# VDD2 0.891586f
C21 VDD2 VSUBS 0.420062f
C22 VDD1 VSUBS 1.740907f
C23 VTAIL VSUBS 0.144029f
C24 VN VSUBS 3.41196f
C25 VP VSUBS 0.648377f
C26 B VSUBS 1.522416f
C27 w_n1294_n1614# VSUBS 26.4131f
C28 VDD2.n0 VSUBS 0.01842f
C29 VDD2.n1 VSUBS 0.017297f
C30 VDD2.n2 VSUBS 0.009295f
C31 VDD2.n3 VSUBS 0.016477f
C32 VDD2.n4 VSUBS 0.013563f
C33 VDD2.t1 VSUBS 0.049051f
C34 VDD2.n5 VSUBS 0.062986f
C35 VDD2.n6 VSUBS 0.175329f
C36 VDD2.n7 VSUBS 0.009295f
C37 VDD2.n8 VSUBS 0.009841f
C38 VDD2.n9 VSUBS 0.021969f
C39 VDD2.n10 VSUBS 0.05119f
C40 VDD2.n11 VSUBS 0.009841f
C41 VDD2.n12 VSUBS 0.009295f
C42 VDD2.n13 VSUBS 0.042107f
C43 VDD2.n14 VSUBS 0.231157f
C44 VDD2.n15 VSUBS 0.01842f
C45 VDD2.n16 VSUBS 0.017297f
C46 VDD2.n17 VSUBS 0.009295f
C47 VDD2.n18 VSUBS 0.016477f
C48 VDD2.n19 VSUBS 0.013563f
C49 VDD2.t0 VSUBS 0.049051f
C50 VDD2.n20 VSUBS 0.062985f
C51 VDD2.n21 VSUBS 0.175329f
C52 VDD2.n22 VSUBS 0.009295f
C53 VDD2.n23 VSUBS 0.009841f
C54 VDD2.n24 VSUBS 0.021969f
C55 VDD2.n25 VSUBS 0.05119f
C56 VDD2.n26 VSUBS 0.009841f
C57 VDD2.n27 VSUBS 0.009295f
C58 VDD2.n28 VSUBS 0.042107f
C59 VDD2.n29 VSUBS 0.037645f
C60 VDD2.n30 VSUBS 1.16638f
C61 VN.t0 VSUBS 0.231548f
C62 VN.t1 VSUBS 0.3172f
C63 B.n0 VSUBS 0.005024f
C64 B.n1 VSUBS 0.005024f
C65 B.n2 VSUBS 0.007945f
C66 B.n3 VSUBS 0.007945f
C67 B.n4 VSUBS 0.007945f
C68 B.n5 VSUBS 0.007945f
C69 B.n6 VSUBS 0.007945f
C70 B.n7 VSUBS 0.007945f
C71 B.n8 VSUBS 0.018195f
C72 B.n9 VSUBS 0.007945f
C73 B.n10 VSUBS 0.007945f
C74 B.n11 VSUBS 0.007945f
C75 B.n12 VSUBS 0.007945f
C76 B.n13 VSUBS 0.007945f
C77 B.n14 VSUBS 0.007945f
C78 B.n15 VSUBS 0.007945f
C79 B.n16 VSUBS 0.005258f
C80 B.n17 VSUBS 0.007945f
C81 B.t11 VSUBS 0.053682f
C82 B.t10 VSUBS 0.059515f
C83 B.t9 VSUBS 0.077642f
C84 B.n18 VSUBS 0.107828f
C85 B.n19 VSUBS 0.100994f
C86 B.n20 VSUBS 0.018408f
C87 B.n21 VSUBS 0.007945f
C88 B.n22 VSUBS 0.007945f
C89 B.n23 VSUBS 0.007945f
C90 B.n24 VSUBS 0.007945f
C91 B.t2 VSUBS 0.053683f
C92 B.t1 VSUBS 0.059516f
C93 B.t0 VSUBS 0.077642f
C94 B.n25 VSUBS 0.107827f
C95 B.n26 VSUBS 0.100993f
C96 B.n27 VSUBS 0.007945f
C97 B.n28 VSUBS 0.007945f
C98 B.n29 VSUBS 0.007945f
C99 B.n30 VSUBS 0.007945f
C100 B.n31 VSUBS 0.007945f
C101 B.n32 VSUBS 0.007945f
C102 B.n33 VSUBS 0.007945f
C103 B.n34 VSUBS 0.018195f
C104 B.n35 VSUBS 0.007945f
C105 B.n36 VSUBS 0.007945f
C106 B.n37 VSUBS 0.007945f
C107 B.n38 VSUBS 0.007945f
C108 B.n39 VSUBS 0.007945f
C109 B.n40 VSUBS 0.007945f
C110 B.n41 VSUBS 0.007945f
C111 B.n42 VSUBS 0.007945f
C112 B.n43 VSUBS 0.007945f
C113 B.n44 VSUBS 0.007945f
C114 B.n45 VSUBS 0.007945f
C115 B.n46 VSUBS 0.007945f
C116 B.n47 VSUBS 0.018195f
C117 B.n48 VSUBS 0.007945f
C118 B.n49 VSUBS 0.007945f
C119 B.n50 VSUBS 0.007945f
C120 B.n51 VSUBS 0.007945f
C121 B.n52 VSUBS 0.007945f
C122 B.n53 VSUBS 0.007945f
C123 B.n54 VSUBS 0.007945f
C124 B.n55 VSUBS 0.005258f
C125 B.n56 VSUBS 0.007945f
C126 B.n57 VSUBS 0.007945f
C127 B.n58 VSUBS 0.007945f
C128 B.n59 VSUBS 0.007945f
C129 B.n60 VSUBS 0.007945f
C130 B.t7 VSUBS 0.053682f
C131 B.t8 VSUBS 0.059515f
C132 B.t6 VSUBS 0.077642f
C133 B.n61 VSUBS 0.107828f
C134 B.n62 VSUBS 0.100994f
C135 B.n63 VSUBS 0.007945f
C136 B.n64 VSUBS 0.007945f
C137 B.n65 VSUBS 0.007945f
C138 B.n66 VSUBS 0.007945f
C139 B.n67 VSUBS 0.007945f
C140 B.n68 VSUBS 0.007945f
C141 B.n69 VSUBS 0.007945f
C142 B.n70 VSUBS 0.018195f
C143 B.n71 VSUBS 0.007945f
C144 B.n72 VSUBS 0.007945f
C145 B.n73 VSUBS 0.007945f
C146 B.n74 VSUBS 0.007945f
C147 B.n75 VSUBS 0.007945f
C148 B.n76 VSUBS 0.007945f
C149 B.n77 VSUBS 0.007945f
C150 B.n78 VSUBS 0.007945f
C151 B.n79 VSUBS 0.007945f
C152 B.n80 VSUBS 0.007945f
C153 B.n81 VSUBS 0.007945f
C154 B.n82 VSUBS 0.007945f
C155 B.n83 VSUBS 0.007945f
C156 B.n84 VSUBS 0.007945f
C157 B.n85 VSUBS 0.007945f
C158 B.n86 VSUBS 0.007945f
C159 B.n87 VSUBS 0.007945f
C160 B.n88 VSUBS 0.007945f
C161 B.n89 VSUBS 0.007945f
C162 B.n90 VSUBS 0.007945f
C163 B.n91 VSUBS 0.007945f
C164 B.n92 VSUBS 0.007945f
C165 B.n93 VSUBS 0.018195f
C166 B.n94 VSUBS 0.018727f
C167 B.n95 VSUBS 0.018727f
C168 B.n96 VSUBS 0.007945f
C169 B.n97 VSUBS 0.007945f
C170 B.n98 VSUBS 0.007945f
C171 B.n99 VSUBS 0.007945f
C172 B.n100 VSUBS 0.007945f
C173 B.n101 VSUBS 0.007945f
C174 B.n102 VSUBS 0.007945f
C175 B.n103 VSUBS 0.007945f
C176 B.n104 VSUBS 0.007945f
C177 B.n105 VSUBS 0.007945f
C178 B.n106 VSUBS 0.007945f
C179 B.n107 VSUBS 0.007945f
C180 B.n108 VSUBS 0.007945f
C181 B.n109 VSUBS 0.007945f
C182 B.n110 VSUBS 0.007945f
C183 B.n111 VSUBS 0.007945f
C184 B.n112 VSUBS 0.007945f
C185 B.n113 VSUBS 0.007945f
C186 B.n114 VSUBS 0.007945f
C187 B.n115 VSUBS 0.007945f
C188 B.n116 VSUBS 0.007945f
C189 B.n117 VSUBS 0.005258f
C190 B.n118 VSUBS 0.018408f
C191 B.n119 VSUBS 0.00666f
C192 B.n120 VSUBS 0.007945f
C193 B.n121 VSUBS 0.007945f
C194 B.n122 VSUBS 0.007945f
C195 B.n123 VSUBS 0.007945f
C196 B.n124 VSUBS 0.007945f
C197 B.n125 VSUBS 0.007945f
C198 B.n126 VSUBS 0.007945f
C199 B.n127 VSUBS 0.007945f
C200 B.n128 VSUBS 0.007945f
C201 B.n129 VSUBS 0.007945f
C202 B.n130 VSUBS 0.007945f
C203 B.t4 VSUBS 0.053683f
C204 B.t5 VSUBS 0.059516f
C205 B.t3 VSUBS 0.077642f
C206 B.n131 VSUBS 0.107827f
C207 B.n132 VSUBS 0.100993f
C208 B.n133 VSUBS 0.018408f
C209 B.n134 VSUBS 0.00666f
C210 B.n135 VSUBS 0.007945f
C211 B.n136 VSUBS 0.007945f
C212 B.n137 VSUBS 0.007945f
C213 B.n138 VSUBS 0.007945f
C214 B.n139 VSUBS 0.007945f
C215 B.n140 VSUBS 0.007945f
C216 B.n141 VSUBS 0.007945f
C217 B.n142 VSUBS 0.007945f
C218 B.n143 VSUBS 0.007945f
C219 B.n144 VSUBS 0.007945f
C220 B.n145 VSUBS 0.007945f
C221 B.n146 VSUBS 0.007945f
C222 B.n147 VSUBS 0.007945f
C223 B.n148 VSUBS 0.007945f
C224 B.n149 VSUBS 0.007945f
C225 B.n150 VSUBS 0.007945f
C226 B.n151 VSUBS 0.007945f
C227 B.n152 VSUBS 0.007945f
C228 B.n153 VSUBS 0.007945f
C229 B.n154 VSUBS 0.007945f
C230 B.n155 VSUBS 0.007945f
C231 B.n156 VSUBS 0.007945f
C232 B.n157 VSUBS 0.007945f
C233 B.n158 VSUBS 0.018727f
C234 B.n159 VSUBS 0.018727f
C235 B.n160 VSUBS 0.018195f
C236 B.n161 VSUBS 0.007945f
C237 B.n162 VSUBS 0.007945f
C238 B.n163 VSUBS 0.007945f
C239 B.n164 VSUBS 0.007945f
C240 B.n165 VSUBS 0.007945f
C241 B.n166 VSUBS 0.007945f
C242 B.n167 VSUBS 0.007945f
C243 B.n168 VSUBS 0.007945f
C244 B.n169 VSUBS 0.007945f
C245 B.n170 VSUBS 0.007945f
C246 B.n171 VSUBS 0.007945f
C247 B.n172 VSUBS 0.007945f
C248 B.n173 VSUBS 0.007945f
C249 B.n174 VSUBS 0.007945f
C250 B.n175 VSUBS 0.007945f
C251 B.n176 VSUBS 0.007945f
C252 B.n177 VSUBS 0.007945f
C253 B.n178 VSUBS 0.007945f
C254 B.n179 VSUBS 0.007945f
C255 B.n180 VSUBS 0.007945f
C256 B.n181 VSUBS 0.007945f
C257 B.n182 VSUBS 0.007945f
C258 B.n183 VSUBS 0.007945f
C259 B.n184 VSUBS 0.007945f
C260 B.n185 VSUBS 0.007945f
C261 B.n186 VSUBS 0.007945f
C262 B.n187 VSUBS 0.007945f
C263 B.n188 VSUBS 0.007945f
C264 B.n189 VSUBS 0.007945f
C265 B.n190 VSUBS 0.007945f
C266 B.n191 VSUBS 0.007945f
C267 B.n192 VSUBS 0.007945f
C268 B.n193 VSUBS 0.007945f
C269 B.n194 VSUBS 0.007945f
C270 B.n195 VSUBS 0.007945f
C271 B.n196 VSUBS 0.007945f
C272 B.n197 VSUBS 0.007945f
C273 B.n198 VSUBS 0.007945f
C274 B.n199 VSUBS 0.019144f
C275 B.n200 VSUBS 0.017778f
C276 B.n201 VSUBS 0.018727f
C277 B.n202 VSUBS 0.007945f
C278 B.n203 VSUBS 0.007945f
C279 B.n204 VSUBS 0.007945f
C280 B.n205 VSUBS 0.007945f
C281 B.n206 VSUBS 0.007945f
C282 B.n207 VSUBS 0.007945f
C283 B.n208 VSUBS 0.007945f
C284 B.n209 VSUBS 0.007945f
C285 B.n210 VSUBS 0.007945f
C286 B.n211 VSUBS 0.007945f
C287 B.n212 VSUBS 0.007945f
C288 B.n213 VSUBS 0.007945f
C289 B.n214 VSUBS 0.007945f
C290 B.n215 VSUBS 0.007945f
C291 B.n216 VSUBS 0.007945f
C292 B.n217 VSUBS 0.007945f
C293 B.n218 VSUBS 0.007945f
C294 B.n219 VSUBS 0.007945f
C295 B.n220 VSUBS 0.007945f
C296 B.n221 VSUBS 0.007945f
C297 B.n222 VSUBS 0.007945f
C298 B.n223 VSUBS 0.005258f
C299 B.n224 VSUBS 0.018408f
C300 B.n225 VSUBS 0.00666f
C301 B.n226 VSUBS 0.007945f
C302 B.n227 VSUBS 0.007945f
C303 B.n228 VSUBS 0.007945f
C304 B.n229 VSUBS 0.007945f
C305 B.n230 VSUBS 0.007945f
C306 B.n231 VSUBS 0.007945f
C307 B.n232 VSUBS 0.007945f
C308 B.n233 VSUBS 0.007945f
C309 B.n234 VSUBS 0.007945f
C310 B.n235 VSUBS 0.007945f
C311 B.n236 VSUBS 0.007945f
C312 B.n237 VSUBS 0.00666f
C313 B.n238 VSUBS 0.007945f
C314 B.n239 VSUBS 0.007945f
C315 B.n240 VSUBS 0.007945f
C316 B.n241 VSUBS 0.007945f
C317 B.n242 VSUBS 0.007945f
C318 B.n243 VSUBS 0.007945f
C319 B.n244 VSUBS 0.007945f
C320 B.n245 VSUBS 0.007945f
C321 B.n246 VSUBS 0.007945f
C322 B.n247 VSUBS 0.007945f
C323 B.n248 VSUBS 0.007945f
C324 B.n249 VSUBS 0.007945f
C325 B.n250 VSUBS 0.007945f
C326 B.n251 VSUBS 0.007945f
C327 B.n252 VSUBS 0.007945f
C328 B.n253 VSUBS 0.007945f
C329 B.n254 VSUBS 0.007945f
C330 B.n255 VSUBS 0.007945f
C331 B.n256 VSUBS 0.007945f
C332 B.n257 VSUBS 0.007945f
C333 B.n258 VSUBS 0.007945f
C334 B.n259 VSUBS 0.007945f
C335 B.n260 VSUBS 0.007945f
C336 B.n261 VSUBS 0.018727f
C337 B.n262 VSUBS 0.018727f
C338 B.n263 VSUBS 0.018195f
C339 B.n264 VSUBS 0.007945f
C340 B.n265 VSUBS 0.007945f
C341 B.n266 VSUBS 0.007945f
C342 B.n267 VSUBS 0.007945f
C343 B.n268 VSUBS 0.007945f
C344 B.n269 VSUBS 0.007945f
C345 B.n270 VSUBS 0.007945f
C346 B.n271 VSUBS 0.007945f
C347 B.n272 VSUBS 0.007945f
C348 B.n273 VSUBS 0.007945f
C349 B.n274 VSUBS 0.007945f
C350 B.n275 VSUBS 0.007945f
C351 B.n276 VSUBS 0.007945f
C352 B.n277 VSUBS 0.007945f
C353 B.n278 VSUBS 0.007945f
C354 B.n279 VSUBS 0.007945f
C355 B.n280 VSUBS 0.007945f
C356 B.n281 VSUBS 0.007945f
C357 B.n282 VSUBS 0.007945f
C358 B.n283 VSUBS 0.017991f
C359 VDD1.n0 VSUBS 0.017961f
C360 VDD1.n1 VSUBS 0.016866f
C361 VDD1.n2 VSUBS 0.009063f
C362 VDD1.n3 VSUBS 0.016066f
C363 VDD1.n4 VSUBS 0.013225f
C364 VDD1.t0 VSUBS 0.047829f
C365 VDD1.n5 VSUBS 0.061416f
C366 VDD1.n6 VSUBS 0.17096f
C367 VDD1.n7 VSUBS 0.009063f
C368 VDD1.n8 VSUBS 0.009596f
C369 VDD1.n9 VSUBS 0.021421f
C370 VDD1.n10 VSUBS 0.049914f
C371 VDD1.n11 VSUBS 0.009596f
C372 VDD1.n12 VSUBS 0.009063f
C373 VDD1.n13 VSUBS 0.041058f
C374 VDD1.n14 VSUBS 0.036919f
C375 VDD1.n15 VSUBS 0.017961f
C376 VDD1.n16 VSUBS 0.016866f
C377 VDD1.n17 VSUBS 0.009063f
C378 VDD1.n18 VSUBS 0.016066f
C379 VDD1.n19 VSUBS 0.013225f
C380 VDD1.t1 VSUBS 0.047829f
C381 VDD1.n20 VSUBS 0.061416f
C382 VDD1.n21 VSUBS 0.17096f
C383 VDD1.n22 VSUBS 0.009063f
C384 VDD1.n23 VSUBS 0.009596f
C385 VDD1.n24 VSUBS 0.021421f
C386 VDD1.n25 VSUBS 0.049914f
C387 VDD1.n26 VSUBS 0.009596f
C388 VDD1.n27 VSUBS 0.009063f
C389 VDD1.n28 VSUBS 0.041058f
C390 VDD1.n29 VSUBS 0.242751f
C391 VTAIL.n0 VSUBS 0.021891f
C392 VTAIL.n1 VSUBS 0.020556f
C393 VTAIL.n2 VSUBS 0.011046f
C394 VTAIL.n3 VSUBS 0.019581f
C395 VTAIL.n4 VSUBS 0.016118f
C396 VTAIL.t2 VSUBS 0.058294f
C397 VTAIL.n5 VSUBS 0.074854f
C398 VTAIL.n6 VSUBS 0.208365f
C399 VTAIL.n7 VSUBS 0.011046f
C400 VTAIL.n8 VSUBS 0.011696f
C401 VTAIL.n9 VSUBS 0.026108f
C402 VTAIL.n10 VSUBS 0.060835f
C403 VTAIL.n11 VSUBS 0.011696f
C404 VTAIL.n12 VSUBS 0.011046f
C405 VTAIL.n13 VSUBS 0.050041f
C406 VTAIL.n14 VSUBS 0.030564f
C407 VTAIL.n15 VSUBS 0.621681f
C408 VTAIL.n16 VSUBS 0.021891f
C409 VTAIL.n17 VSUBS 0.020556f
C410 VTAIL.n18 VSUBS 0.011046f
C411 VTAIL.n19 VSUBS 0.019581f
C412 VTAIL.n20 VSUBS 0.016118f
C413 VTAIL.t0 VSUBS 0.058294f
C414 VTAIL.n21 VSUBS 0.074854f
C415 VTAIL.n22 VSUBS 0.208365f
C416 VTAIL.n23 VSUBS 0.011046f
C417 VTAIL.n24 VSUBS 0.011696f
C418 VTAIL.n25 VSUBS 0.026108f
C419 VTAIL.n26 VSUBS 0.060835f
C420 VTAIL.n27 VSUBS 0.011696f
C421 VTAIL.n28 VSUBS 0.011046f
C422 VTAIL.n29 VSUBS 0.050041f
C423 VTAIL.n30 VSUBS 0.030564f
C424 VTAIL.n31 VSUBS 0.62939f
C425 VTAIL.n32 VSUBS 0.021891f
C426 VTAIL.n33 VSUBS 0.020556f
C427 VTAIL.n34 VSUBS 0.011046f
C428 VTAIL.n35 VSUBS 0.019581f
C429 VTAIL.n36 VSUBS 0.016118f
C430 VTAIL.t1 VSUBS 0.058294f
C431 VTAIL.n37 VSUBS 0.074854f
C432 VTAIL.n38 VSUBS 0.208365f
C433 VTAIL.n39 VSUBS 0.011046f
C434 VTAIL.n40 VSUBS 0.011696f
C435 VTAIL.n41 VSUBS 0.026108f
C436 VTAIL.n42 VSUBS 0.060835f
C437 VTAIL.n43 VSUBS 0.011696f
C438 VTAIL.n44 VSUBS 0.011046f
C439 VTAIL.n45 VSUBS 0.050041f
C440 VTAIL.n46 VSUBS 0.030564f
C441 VTAIL.n47 VSUBS 0.583139f
C442 VTAIL.n48 VSUBS 0.021891f
C443 VTAIL.n49 VSUBS 0.020556f
C444 VTAIL.n50 VSUBS 0.011046f
C445 VTAIL.n51 VSUBS 0.019581f
C446 VTAIL.n52 VSUBS 0.016118f
C447 VTAIL.t3 VSUBS 0.058294f
C448 VTAIL.n53 VSUBS 0.074854f
C449 VTAIL.n54 VSUBS 0.208365f
C450 VTAIL.n55 VSUBS 0.011046f
C451 VTAIL.n56 VSUBS 0.011696f
C452 VTAIL.n57 VSUBS 0.026108f
C453 VTAIL.n58 VSUBS 0.060835f
C454 VTAIL.n59 VSUBS 0.011696f
C455 VTAIL.n60 VSUBS 0.011046f
C456 VTAIL.n61 VSUBS 0.050041f
C457 VTAIL.n62 VSUBS 0.030564f
C458 VTAIL.n63 VSUBS 0.536603f
C459 VP.t1 VSUBS 0.320891f
C460 VP.t0 VSUBS 0.236445f
C461 VP.n0 VSUBS 2.23368f
.ends

