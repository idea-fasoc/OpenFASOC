* NGSPICE file created from diff_pair_sample_0480.ext - technology: sky130A

.subckt diff_pair_sample_0480 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=1.43055 pd=9 as=3.3813 ps=18.12 w=8.67 l=2.7
X1 B.t11 B.t9 B.t10 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=0 ps=0 w=8.67 l=2.7
X2 VTAIL.t2 VN.t0 VDD2.t3 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=1.43055 ps=9 w=8.67 l=2.7
X3 VDD1.t2 VP.t1 VTAIL.t7 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=1.43055 pd=9 as=3.3813 ps=18.12 w=8.67 l=2.7
X4 B.t8 B.t6 B.t7 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=0 ps=0 w=8.67 l=2.7
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=1.43055 pd=9 as=3.3813 ps=18.12 w=8.67 l=2.7
X6 B.t5 B.t3 B.t4 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=0 ps=0 w=8.67 l=2.7
X7 VTAIL.t1 VN.t2 VDD2.t1 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=1.43055 ps=9 w=8.67 l=2.7
X8 B.t2 B.t0 B.t1 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=0 ps=0 w=8.67 l=2.7
X9 VTAIL.t5 VP.t2 VDD1.t1 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=1.43055 ps=9 w=8.67 l=2.7
X10 VDD2.t0 VN.t3 VTAIL.t3 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=1.43055 pd=9 as=3.3813 ps=18.12 w=8.67 l=2.7
X11 VTAIL.t4 VP.t3 VDD1.t0 w_n2788_n2702# sky130_fd_pr__pfet_01v8 ad=3.3813 pd=18.12 as=1.43055 ps=9 w=8.67 l=2.7
R0 VP.n16 VP.n0 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n13 VP.n1 161.3
R3 VP.n12 VP.n11 161.3
R4 VP.n10 VP.n2 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n3 161.3
R7 VP.n4 VP.t2 111.403
R8 VP.n4 VP.t0 110.531
R9 VP.n6 VP.n5 110.022
R10 VP.n18 VP.n17 110.022
R11 VP.n5 VP.t3 77.3883
R12 VP.n17 VP.t1 77.3883
R13 VP.n6 VP.n4 47.6506
R14 VP.n11 VP.n10 40.4934
R15 VP.n11 VP.n1 40.4934
R16 VP.n9 VP.n3 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n1 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n5 VP.n3 0.73451
R21 VP.n17 VP.n16 0.73451
R22 VP.n7 VP.n6 0.278367
R23 VP.n18 VP.n0 0.278367
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153454
R31 VTAIL.n362 VTAIL.n322 756.745
R32 VTAIL.n40 VTAIL.n0 756.745
R33 VTAIL.n86 VTAIL.n46 756.745
R34 VTAIL.n132 VTAIL.n92 756.745
R35 VTAIL.n316 VTAIL.n276 756.745
R36 VTAIL.n270 VTAIL.n230 756.745
R37 VTAIL.n224 VTAIL.n184 756.745
R38 VTAIL.n178 VTAIL.n138 756.745
R39 VTAIL.n337 VTAIL.n336 585
R40 VTAIL.n334 VTAIL.n333 585
R41 VTAIL.n343 VTAIL.n342 585
R42 VTAIL.n345 VTAIL.n344 585
R43 VTAIL.n330 VTAIL.n329 585
R44 VTAIL.n351 VTAIL.n350 585
R45 VTAIL.n354 VTAIL.n353 585
R46 VTAIL.n352 VTAIL.n326 585
R47 VTAIL.n359 VTAIL.n325 585
R48 VTAIL.n361 VTAIL.n360 585
R49 VTAIL.n363 VTAIL.n362 585
R50 VTAIL.n15 VTAIL.n14 585
R51 VTAIL.n12 VTAIL.n11 585
R52 VTAIL.n21 VTAIL.n20 585
R53 VTAIL.n23 VTAIL.n22 585
R54 VTAIL.n8 VTAIL.n7 585
R55 VTAIL.n29 VTAIL.n28 585
R56 VTAIL.n32 VTAIL.n31 585
R57 VTAIL.n30 VTAIL.n4 585
R58 VTAIL.n37 VTAIL.n3 585
R59 VTAIL.n39 VTAIL.n38 585
R60 VTAIL.n41 VTAIL.n40 585
R61 VTAIL.n61 VTAIL.n60 585
R62 VTAIL.n58 VTAIL.n57 585
R63 VTAIL.n67 VTAIL.n66 585
R64 VTAIL.n69 VTAIL.n68 585
R65 VTAIL.n54 VTAIL.n53 585
R66 VTAIL.n75 VTAIL.n74 585
R67 VTAIL.n78 VTAIL.n77 585
R68 VTAIL.n76 VTAIL.n50 585
R69 VTAIL.n83 VTAIL.n49 585
R70 VTAIL.n85 VTAIL.n84 585
R71 VTAIL.n87 VTAIL.n86 585
R72 VTAIL.n107 VTAIL.n106 585
R73 VTAIL.n104 VTAIL.n103 585
R74 VTAIL.n113 VTAIL.n112 585
R75 VTAIL.n115 VTAIL.n114 585
R76 VTAIL.n100 VTAIL.n99 585
R77 VTAIL.n121 VTAIL.n120 585
R78 VTAIL.n124 VTAIL.n123 585
R79 VTAIL.n122 VTAIL.n96 585
R80 VTAIL.n129 VTAIL.n95 585
R81 VTAIL.n131 VTAIL.n130 585
R82 VTAIL.n133 VTAIL.n132 585
R83 VTAIL.n317 VTAIL.n316 585
R84 VTAIL.n315 VTAIL.n314 585
R85 VTAIL.n313 VTAIL.n279 585
R86 VTAIL.n283 VTAIL.n280 585
R87 VTAIL.n308 VTAIL.n307 585
R88 VTAIL.n306 VTAIL.n305 585
R89 VTAIL.n285 VTAIL.n284 585
R90 VTAIL.n300 VTAIL.n299 585
R91 VTAIL.n298 VTAIL.n297 585
R92 VTAIL.n289 VTAIL.n288 585
R93 VTAIL.n292 VTAIL.n291 585
R94 VTAIL.n271 VTAIL.n270 585
R95 VTAIL.n269 VTAIL.n268 585
R96 VTAIL.n267 VTAIL.n233 585
R97 VTAIL.n237 VTAIL.n234 585
R98 VTAIL.n262 VTAIL.n261 585
R99 VTAIL.n260 VTAIL.n259 585
R100 VTAIL.n239 VTAIL.n238 585
R101 VTAIL.n254 VTAIL.n253 585
R102 VTAIL.n252 VTAIL.n251 585
R103 VTAIL.n243 VTAIL.n242 585
R104 VTAIL.n246 VTAIL.n245 585
R105 VTAIL.n225 VTAIL.n224 585
R106 VTAIL.n223 VTAIL.n222 585
R107 VTAIL.n221 VTAIL.n187 585
R108 VTAIL.n191 VTAIL.n188 585
R109 VTAIL.n216 VTAIL.n215 585
R110 VTAIL.n214 VTAIL.n213 585
R111 VTAIL.n193 VTAIL.n192 585
R112 VTAIL.n208 VTAIL.n207 585
R113 VTAIL.n206 VTAIL.n205 585
R114 VTAIL.n197 VTAIL.n196 585
R115 VTAIL.n200 VTAIL.n199 585
R116 VTAIL.n179 VTAIL.n178 585
R117 VTAIL.n177 VTAIL.n176 585
R118 VTAIL.n175 VTAIL.n141 585
R119 VTAIL.n145 VTAIL.n142 585
R120 VTAIL.n170 VTAIL.n169 585
R121 VTAIL.n168 VTAIL.n167 585
R122 VTAIL.n147 VTAIL.n146 585
R123 VTAIL.n162 VTAIL.n161 585
R124 VTAIL.n160 VTAIL.n159 585
R125 VTAIL.n151 VTAIL.n150 585
R126 VTAIL.n154 VTAIL.n153 585
R127 VTAIL.t6 VTAIL.n290 329.039
R128 VTAIL.t5 VTAIL.n244 329.039
R129 VTAIL.t0 VTAIL.n198 329.039
R130 VTAIL.t1 VTAIL.n152 329.039
R131 VTAIL.t3 VTAIL.n335 329.038
R132 VTAIL.t2 VTAIL.n13 329.038
R133 VTAIL.t7 VTAIL.n59 329.038
R134 VTAIL.t4 VTAIL.n105 329.038
R135 VTAIL.n336 VTAIL.n333 171.744
R136 VTAIL.n343 VTAIL.n333 171.744
R137 VTAIL.n344 VTAIL.n343 171.744
R138 VTAIL.n344 VTAIL.n329 171.744
R139 VTAIL.n351 VTAIL.n329 171.744
R140 VTAIL.n353 VTAIL.n351 171.744
R141 VTAIL.n353 VTAIL.n352 171.744
R142 VTAIL.n352 VTAIL.n325 171.744
R143 VTAIL.n361 VTAIL.n325 171.744
R144 VTAIL.n362 VTAIL.n361 171.744
R145 VTAIL.n14 VTAIL.n11 171.744
R146 VTAIL.n21 VTAIL.n11 171.744
R147 VTAIL.n22 VTAIL.n21 171.744
R148 VTAIL.n22 VTAIL.n7 171.744
R149 VTAIL.n29 VTAIL.n7 171.744
R150 VTAIL.n31 VTAIL.n29 171.744
R151 VTAIL.n31 VTAIL.n30 171.744
R152 VTAIL.n30 VTAIL.n3 171.744
R153 VTAIL.n39 VTAIL.n3 171.744
R154 VTAIL.n40 VTAIL.n39 171.744
R155 VTAIL.n60 VTAIL.n57 171.744
R156 VTAIL.n67 VTAIL.n57 171.744
R157 VTAIL.n68 VTAIL.n67 171.744
R158 VTAIL.n68 VTAIL.n53 171.744
R159 VTAIL.n75 VTAIL.n53 171.744
R160 VTAIL.n77 VTAIL.n75 171.744
R161 VTAIL.n77 VTAIL.n76 171.744
R162 VTAIL.n76 VTAIL.n49 171.744
R163 VTAIL.n85 VTAIL.n49 171.744
R164 VTAIL.n86 VTAIL.n85 171.744
R165 VTAIL.n106 VTAIL.n103 171.744
R166 VTAIL.n113 VTAIL.n103 171.744
R167 VTAIL.n114 VTAIL.n113 171.744
R168 VTAIL.n114 VTAIL.n99 171.744
R169 VTAIL.n121 VTAIL.n99 171.744
R170 VTAIL.n123 VTAIL.n121 171.744
R171 VTAIL.n123 VTAIL.n122 171.744
R172 VTAIL.n122 VTAIL.n95 171.744
R173 VTAIL.n131 VTAIL.n95 171.744
R174 VTAIL.n132 VTAIL.n131 171.744
R175 VTAIL.n316 VTAIL.n315 171.744
R176 VTAIL.n315 VTAIL.n279 171.744
R177 VTAIL.n283 VTAIL.n279 171.744
R178 VTAIL.n307 VTAIL.n283 171.744
R179 VTAIL.n307 VTAIL.n306 171.744
R180 VTAIL.n306 VTAIL.n284 171.744
R181 VTAIL.n299 VTAIL.n284 171.744
R182 VTAIL.n299 VTAIL.n298 171.744
R183 VTAIL.n298 VTAIL.n288 171.744
R184 VTAIL.n291 VTAIL.n288 171.744
R185 VTAIL.n270 VTAIL.n269 171.744
R186 VTAIL.n269 VTAIL.n233 171.744
R187 VTAIL.n237 VTAIL.n233 171.744
R188 VTAIL.n261 VTAIL.n237 171.744
R189 VTAIL.n261 VTAIL.n260 171.744
R190 VTAIL.n260 VTAIL.n238 171.744
R191 VTAIL.n253 VTAIL.n238 171.744
R192 VTAIL.n253 VTAIL.n252 171.744
R193 VTAIL.n252 VTAIL.n242 171.744
R194 VTAIL.n245 VTAIL.n242 171.744
R195 VTAIL.n224 VTAIL.n223 171.744
R196 VTAIL.n223 VTAIL.n187 171.744
R197 VTAIL.n191 VTAIL.n187 171.744
R198 VTAIL.n215 VTAIL.n191 171.744
R199 VTAIL.n215 VTAIL.n214 171.744
R200 VTAIL.n214 VTAIL.n192 171.744
R201 VTAIL.n207 VTAIL.n192 171.744
R202 VTAIL.n207 VTAIL.n206 171.744
R203 VTAIL.n206 VTAIL.n196 171.744
R204 VTAIL.n199 VTAIL.n196 171.744
R205 VTAIL.n178 VTAIL.n177 171.744
R206 VTAIL.n177 VTAIL.n141 171.744
R207 VTAIL.n145 VTAIL.n141 171.744
R208 VTAIL.n169 VTAIL.n145 171.744
R209 VTAIL.n169 VTAIL.n168 171.744
R210 VTAIL.n168 VTAIL.n146 171.744
R211 VTAIL.n161 VTAIL.n146 171.744
R212 VTAIL.n161 VTAIL.n160 171.744
R213 VTAIL.n160 VTAIL.n150 171.744
R214 VTAIL.n153 VTAIL.n150 171.744
R215 VTAIL.n336 VTAIL.t3 85.8723
R216 VTAIL.n14 VTAIL.t2 85.8723
R217 VTAIL.n60 VTAIL.t7 85.8723
R218 VTAIL.n106 VTAIL.t4 85.8723
R219 VTAIL.n291 VTAIL.t6 85.8723
R220 VTAIL.n245 VTAIL.t5 85.8723
R221 VTAIL.n199 VTAIL.t0 85.8723
R222 VTAIL.n153 VTAIL.t1 85.8723
R223 VTAIL.n367 VTAIL.n366 35.0944
R224 VTAIL.n45 VTAIL.n44 35.0944
R225 VTAIL.n91 VTAIL.n90 35.0944
R226 VTAIL.n137 VTAIL.n136 35.0944
R227 VTAIL.n321 VTAIL.n320 35.0944
R228 VTAIL.n275 VTAIL.n274 35.0944
R229 VTAIL.n229 VTAIL.n228 35.0944
R230 VTAIL.n183 VTAIL.n182 35.0944
R231 VTAIL.n367 VTAIL.n321 22.4531
R232 VTAIL.n183 VTAIL.n137 22.4531
R233 VTAIL.n360 VTAIL.n359 13.1884
R234 VTAIL.n38 VTAIL.n37 13.1884
R235 VTAIL.n84 VTAIL.n83 13.1884
R236 VTAIL.n130 VTAIL.n129 13.1884
R237 VTAIL.n314 VTAIL.n313 13.1884
R238 VTAIL.n268 VTAIL.n267 13.1884
R239 VTAIL.n222 VTAIL.n221 13.1884
R240 VTAIL.n176 VTAIL.n175 13.1884
R241 VTAIL.n358 VTAIL.n326 12.8005
R242 VTAIL.n363 VTAIL.n324 12.8005
R243 VTAIL.n36 VTAIL.n4 12.8005
R244 VTAIL.n41 VTAIL.n2 12.8005
R245 VTAIL.n82 VTAIL.n50 12.8005
R246 VTAIL.n87 VTAIL.n48 12.8005
R247 VTAIL.n128 VTAIL.n96 12.8005
R248 VTAIL.n133 VTAIL.n94 12.8005
R249 VTAIL.n317 VTAIL.n278 12.8005
R250 VTAIL.n312 VTAIL.n280 12.8005
R251 VTAIL.n271 VTAIL.n232 12.8005
R252 VTAIL.n266 VTAIL.n234 12.8005
R253 VTAIL.n225 VTAIL.n186 12.8005
R254 VTAIL.n220 VTAIL.n188 12.8005
R255 VTAIL.n179 VTAIL.n140 12.8005
R256 VTAIL.n174 VTAIL.n142 12.8005
R257 VTAIL.n355 VTAIL.n354 12.0247
R258 VTAIL.n364 VTAIL.n322 12.0247
R259 VTAIL.n33 VTAIL.n32 12.0247
R260 VTAIL.n42 VTAIL.n0 12.0247
R261 VTAIL.n79 VTAIL.n78 12.0247
R262 VTAIL.n88 VTAIL.n46 12.0247
R263 VTAIL.n125 VTAIL.n124 12.0247
R264 VTAIL.n134 VTAIL.n92 12.0247
R265 VTAIL.n318 VTAIL.n276 12.0247
R266 VTAIL.n309 VTAIL.n308 12.0247
R267 VTAIL.n272 VTAIL.n230 12.0247
R268 VTAIL.n263 VTAIL.n262 12.0247
R269 VTAIL.n226 VTAIL.n184 12.0247
R270 VTAIL.n217 VTAIL.n216 12.0247
R271 VTAIL.n180 VTAIL.n138 12.0247
R272 VTAIL.n171 VTAIL.n170 12.0247
R273 VTAIL.n350 VTAIL.n328 11.249
R274 VTAIL.n28 VTAIL.n6 11.249
R275 VTAIL.n74 VTAIL.n52 11.249
R276 VTAIL.n120 VTAIL.n98 11.249
R277 VTAIL.n305 VTAIL.n282 11.249
R278 VTAIL.n259 VTAIL.n236 11.249
R279 VTAIL.n213 VTAIL.n190 11.249
R280 VTAIL.n167 VTAIL.n144 11.249
R281 VTAIL.n337 VTAIL.n335 10.7239
R282 VTAIL.n15 VTAIL.n13 10.7239
R283 VTAIL.n61 VTAIL.n59 10.7239
R284 VTAIL.n107 VTAIL.n105 10.7239
R285 VTAIL.n292 VTAIL.n290 10.7239
R286 VTAIL.n246 VTAIL.n244 10.7239
R287 VTAIL.n200 VTAIL.n198 10.7239
R288 VTAIL.n154 VTAIL.n152 10.7239
R289 VTAIL.n349 VTAIL.n330 10.4732
R290 VTAIL.n27 VTAIL.n8 10.4732
R291 VTAIL.n73 VTAIL.n54 10.4732
R292 VTAIL.n119 VTAIL.n100 10.4732
R293 VTAIL.n304 VTAIL.n285 10.4732
R294 VTAIL.n258 VTAIL.n239 10.4732
R295 VTAIL.n212 VTAIL.n193 10.4732
R296 VTAIL.n166 VTAIL.n147 10.4732
R297 VTAIL.n346 VTAIL.n345 9.69747
R298 VTAIL.n24 VTAIL.n23 9.69747
R299 VTAIL.n70 VTAIL.n69 9.69747
R300 VTAIL.n116 VTAIL.n115 9.69747
R301 VTAIL.n301 VTAIL.n300 9.69747
R302 VTAIL.n255 VTAIL.n254 9.69747
R303 VTAIL.n209 VTAIL.n208 9.69747
R304 VTAIL.n163 VTAIL.n162 9.69747
R305 VTAIL.n366 VTAIL.n365 9.45567
R306 VTAIL.n44 VTAIL.n43 9.45567
R307 VTAIL.n90 VTAIL.n89 9.45567
R308 VTAIL.n136 VTAIL.n135 9.45567
R309 VTAIL.n320 VTAIL.n319 9.45567
R310 VTAIL.n274 VTAIL.n273 9.45567
R311 VTAIL.n228 VTAIL.n227 9.45567
R312 VTAIL.n182 VTAIL.n181 9.45567
R313 VTAIL.n365 VTAIL.n364 9.3005
R314 VTAIL.n324 VTAIL.n323 9.3005
R315 VTAIL.n339 VTAIL.n338 9.3005
R316 VTAIL.n341 VTAIL.n340 9.3005
R317 VTAIL.n332 VTAIL.n331 9.3005
R318 VTAIL.n347 VTAIL.n346 9.3005
R319 VTAIL.n349 VTAIL.n348 9.3005
R320 VTAIL.n328 VTAIL.n327 9.3005
R321 VTAIL.n356 VTAIL.n355 9.3005
R322 VTAIL.n358 VTAIL.n357 9.3005
R323 VTAIL.n43 VTAIL.n42 9.3005
R324 VTAIL.n2 VTAIL.n1 9.3005
R325 VTAIL.n17 VTAIL.n16 9.3005
R326 VTAIL.n19 VTAIL.n18 9.3005
R327 VTAIL.n10 VTAIL.n9 9.3005
R328 VTAIL.n25 VTAIL.n24 9.3005
R329 VTAIL.n27 VTAIL.n26 9.3005
R330 VTAIL.n6 VTAIL.n5 9.3005
R331 VTAIL.n34 VTAIL.n33 9.3005
R332 VTAIL.n36 VTAIL.n35 9.3005
R333 VTAIL.n89 VTAIL.n88 9.3005
R334 VTAIL.n48 VTAIL.n47 9.3005
R335 VTAIL.n63 VTAIL.n62 9.3005
R336 VTAIL.n65 VTAIL.n64 9.3005
R337 VTAIL.n56 VTAIL.n55 9.3005
R338 VTAIL.n71 VTAIL.n70 9.3005
R339 VTAIL.n73 VTAIL.n72 9.3005
R340 VTAIL.n52 VTAIL.n51 9.3005
R341 VTAIL.n80 VTAIL.n79 9.3005
R342 VTAIL.n82 VTAIL.n81 9.3005
R343 VTAIL.n135 VTAIL.n134 9.3005
R344 VTAIL.n94 VTAIL.n93 9.3005
R345 VTAIL.n109 VTAIL.n108 9.3005
R346 VTAIL.n111 VTAIL.n110 9.3005
R347 VTAIL.n102 VTAIL.n101 9.3005
R348 VTAIL.n117 VTAIL.n116 9.3005
R349 VTAIL.n119 VTAIL.n118 9.3005
R350 VTAIL.n98 VTAIL.n97 9.3005
R351 VTAIL.n126 VTAIL.n125 9.3005
R352 VTAIL.n128 VTAIL.n127 9.3005
R353 VTAIL.n294 VTAIL.n293 9.3005
R354 VTAIL.n296 VTAIL.n295 9.3005
R355 VTAIL.n287 VTAIL.n286 9.3005
R356 VTAIL.n302 VTAIL.n301 9.3005
R357 VTAIL.n304 VTAIL.n303 9.3005
R358 VTAIL.n282 VTAIL.n281 9.3005
R359 VTAIL.n310 VTAIL.n309 9.3005
R360 VTAIL.n312 VTAIL.n311 9.3005
R361 VTAIL.n319 VTAIL.n318 9.3005
R362 VTAIL.n278 VTAIL.n277 9.3005
R363 VTAIL.n248 VTAIL.n247 9.3005
R364 VTAIL.n250 VTAIL.n249 9.3005
R365 VTAIL.n241 VTAIL.n240 9.3005
R366 VTAIL.n256 VTAIL.n255 9.3005
R367 VTAIL.n258 VTAIL.n257 9.3005
R368 VTAIL.n236 VTAIL.n235 9.3005
R369 VTAIL.n264 VTAIL.n263 9.3005
R370 VTAIL.n266 VTAIL.n265 9.3005
R371 VTAIL.n273 VTAIL.n272 9.3005
R372 VTAIL.n232 VTAIL.n231 9.3005
R373 VTAIL.n202 VTAIL.n201 9.3005
R374 VTAIL.n204 VTAIL.n203 9.3005
R375 VTAIL.n195 VTAIL.n194 9.3005
R376 VTAIL.n210 VTAIL.n209 9.3005
R377 VTAIL.n212 VTAIL.n211 9.3005
R378 VTAIL.n190 VTAIL.n189 9.3005
R379 VTAIL.n218 VTAIL.n217 9.3005
R380 VTAIL.n220 VTAIL.n219 9.3005
R381 VTAIL.n227 VTAIL.n226 9.3005
R382 VTAIL.n186 VTAIL.n185 9.3005
R383 VTAIL.n156 VTAIL.n155 9.3005
R384 VTAIL.n158 VTAIL.n157 9.3005
R385 VTAIL.n149 VTAIL.n148 9.3005
R386 VTAIL.n164 VTAIL.n163 9.3005
R387 VTAIL.n166 VTAIL.n165 9.3005
R388 VTAIL.n144 VTAIL.n143 9.3005
R389 VTAIL.n172 VTAIL.n171 9.3005
R390 VTAIL.n174 VTAIL.n173 9.3005
R391 VTAIL.n181 VTAIL.n180 9.3005
R392 VTAIL.n140 VTAIL.n139 9.3005
R393 VTAIL.n342 VTAIL.n332 8.92171
R394 VTAIL.n20 VTAIL.n10 8.92171
R395 VTAIL.n66 VTAIL.n56 8.92171
R396 VTAIL.n112 VTAIL.n102 8.92171
R397 VTAIL.n297 VTAIL.n287 8.92171
R398 VTAIL.n251 VTAIL.n241 8.92171
R399 VTAIL.n205 VTAIL.n195 8.92171
R400 VTAIL.n159 VTAIL.n149 8.92171
R401 VTAIL.n341 VTAIL.n334 8.14595
R402 VTAIL.n19 VTAIL.n12 8.14595
R403 VTAIL.n65 VTAIL.n58 8.14595
R404 VTAIL.n111 VTAIL.n104 8.14595
R405 VTAIL.n296 VTAIL.n289 8.14595
R406 VTAIL.n250 VTAIL.n243 8.14595
R407 VTAIL.n204 VTAIL.n197 8.14595
R408 VTAIL.n158 VTAIL.n151 8.14595
R409 VTAIL.n338 VTAIL.n337 7.3702
R410 VTAIL.n16 VTAIL.n15 7.3702
R411 VTAIL.n62 VTAIL.n61 7.3702
R412 VTAIL.n108 VTAIL.n107 7.3702
R413 VTAIL.n293 VTAIL.n292 7.3702
R414 VTAIL.n247 VTAIL.n246 7.3702
R415 VTAIL.n201 VTAIL.n200 7.3702
R416 VTAIL.n155 VTAIL.n154 7.3702
R417 VTAIL.n338 VTAIL.n334 5.81868
R418 VTAIL.n16 VTAIL.n12 5.81868
R419 VTAIL.n62 VTAIL.n58 5.81868
R420 VTAIL.n108 VTAIL.n104 5.81868
R421 VTAIL.n293 VTAIL.n289 5.81868
R422 VTAIL.n247 VTAIL.n243 5.81868
R423 VTAIL.n201 VTAIL.n197 5.81868
R424 VTAIL.n155 VTAIL.n151 5.81868
R425 VTAIL.n342 VTAIL.n341 5.04292
R426 VTAIL.n20 VTAIL.n19 5.04292
R427 VTAIL.n66 VTAIL.n65 5.04292
R428 VTAIL.n112 VTAIL.n111 5.04292
R429 VTAIL.n297 VTAIL.n296 5.04292
R430 VTAIL.n251 VTAIL.n250 5.04292
R431 VTAIL.n205 VTAIL.n204 5.04292
R432 VTAIL.n159 VTAIL.n158 5.04292
R433 VTAIL.n345 VTAIL.n332 4.26717
R434 VTAIL.n23 VTAIL.n10 4.26717
R435 VTAIL.n69 VTAIL.n56 4.26717
R436 VTAIL.n115 VTAIL.n102 4.26717
R437 VTAIL.n300 VTAIL.n287 4.26717
R438 VTAIL.n254 VTAIL.n241 4.26717
R439 VTAIL.n208 VTAIL.n195 4.26717
R440 VTAIL.n162 VTAIL.n149 4.26717
R441 VTAIL.n346 VTAIL.n330 3.49141
R442 VTAIL.n24 VTAIL.n8 3.49141
R443 VTAIL.n70 VTAIL.n54 3.49141
R444 VTAIL.n116 VTAIL.n100 3.49141
R445 VTAIL.n301 VTAIL.n285 3.49141
R446 VTAIL.n255 VTAIL.n239 3.49141
R447 VTAIL.n209 VTAIL.n193 3.49141
R448 VTAIL.n163 VTAIL.n147 3.49141
R449 VTAIL.n350 VTAIL.n349 2.71565
R450 VTAIL.n28 VTAIL.n27 2.71565
R451 VTAIL.n74 VTAIL.n73 2.71565
R452 VTAIL.n120 VTAIL.n119 2.71565
R453 VTAIL.n305 VTAIL.n304 2.71565
R454 VTAIL.n259 VTAIL.n258 2.71565
R455 VTAIL.n213 VTAIL.n212 2.71565
R456 VTAIL.n167 VTAIL.n166 2.71565
R457 VTAIL.n229 VTAIL.n183 2.61257
R458 VTAIL.n321 VTAIL.n275 2.61257
R459 VTAIL.n137 VTAIL.n91 2.61257
R460 VTAIL.n339 VTAIL.n335 2.41285
R461 VTAIL.n17 VTAIL.n13 2.41285
R462 VTAIL.n63 VTAIL.n59 2.41285
R463 VTAIL.n109 VTAIL.n105 2.41285
R464 VTAIL.n294 VTAIL.n290 2.41285
R465 VTAIL.n248 VTAIL.n244 2.41285
R466 VTAIL.n202 VTAIL.n198 2.41285
R467 VTAIL.n156 VTAIL.n152 2.41285
R468 VTAIL.n354 VTAIL.n328 1.93989
R469 VTAIL.n366 VTAIL.n322 1.93989
R470 VTAIL.n32 VTAIL.n6 1.93989
R471 VTAIL.n44 VTAIL.n0 1.93989
R472 VTAIL.n78 VTAIL.n52 1.93989
R473 VTAIL.n90 VTAIL.n46 1.93989
R474 VTAIL.n124 VTAIL.n98 1.93989
R475 VTAIL.n136 VTAIL.n92 1.93989
R476 VTAIL.n320 VTAIL.n276 1.93989
R477 VTAIL.n308 VTAIL.n282 1.93989
R478 VTAIL.n274 VTAIL.n230 1.93989
R479 VTAIL.n262 VTAIL.n236 1.93989
R480 VTAIL.n228 VTAIL.n184 1.93989
R481 VTAIL.n216 VTAIL.n190 1.93989
R482 VTAIL.n182 VTAIL.n138 1.93989
R483 VTAIL.n170 VTAIL.n144 1.93989
R484 VTAIL VTAIL.n45 1.36472
R485 VTAIL VTAIL.n367 1.24834
R486 VTAIL.n355 VTAIL.n326 1.16414
R487 VTAIL.n364 VTAIL.n363 1.16414
R488 VTAIL.n33 VTAIL.n4 1.16414
R489 VTAIL.n42 VTAIL.n41 1.16414
R490 VTAIL.n79 VTAIL.n50 1.16414
R491 VTAIL.n88 VTAIL.n87 1.16414
R492 VTAIL.n125 VTAIL.n96 1.16414
R493 VTAIL.n134 VTAIL.n133 1.16414
R494 VTAIL.n318 VTAIL.n317 1.16414
R495 VTAIL.n309 VTAIL.n280 1.16414
R496 VTAIL.n272 VTAIL.n271 1.16414
R497 VTAIL.n263 VTAIL.n234 1.16414
R498 VTAIL.n226 VTAIL.n225 1.16414
R499 VTAIL.n217 VTAIL.n188 1.16414
R500 VTAIL.n180 VTAIL.n179 1.16414
R501 VTAIL.n171 VTAIL.n142 1.16414
R502 VTAIL.n275 VTAIL.n229 0.470328
R503 VTAIL.n91 VTAIL.n45 0.470328
R504 VTAIL.n359 VTAIL.n358 0.388379
R505 VTAIL.n360 VTAIL.n324 0.388379
R506 VTAIL.n37 VTAIL.n36 0.388379
R507 VTAIL.n38 VTAIL.n2 0.388379
R508 VTAIL.n83 VTAIL.n82 0.388379
R509 VTAIL.n84 VTAIL.n48 0.388379
R510 VTAIL.n129 VTAIL.n128 0.388379
R511 VTAIL.n130 VTAIL.n94 0.388379
R512 VTAIL.n314 VTAIL.n278 0.388379
R513 VTAIL.n313 VTAIL.n312 0.388379
R514 VTAIL.n268 VTAIL.n232 0.388379
R515 VTAIL.n267 VTAIL.n266 0.388379
R516 VTAIL.n222 VTAIL.n186 0.388379
R517 VTAIL.n221 VTAIL.n220 0.388379
R518 VTAIL.n176 VTAIL.n140 0.388379
R519 VTAIL.n175 VTAIL.n174 0.388379
R520 VTAIL.n340 VTAIL.n339 0.155672
R521 VTAIL.n340 VTAIL.n331 0.155672
R522 VTAIL.n347 VTAIL.n331 0.155672
R523 VTAIL.n348 VTAIL.n347 0.155672
R524 VTAIL.n348 VTAIL.n327 0.155672
R525 VTAIL.n356 VTAIL.n327 0.155672
R526 VTAIL.n357 VTAIL.n356 0.155672
R527 VTAIL.n357 VTAIL.n323 0.155672
R528 VTAIL.n365 VTAIL.n323 0.155672
R529 VTAIL.n18 VTAIL.n17 0.155672
R530 VTAIL.n18 VTAIL.n9 0.155672
R531 VTAIL.n25 VTAIL.n9 0.155672
R532 VTAIL.n26 VTAIL.n25 0.155672
R533 VTAIL.n26 VTAIL.n5 0.155672
R534 VTAIL.n34 VTAIL.n5 0.155672
R535 VTAIL.n35 VTAIL.n34 0.155672
R536 VTAIL.n35 VTAIL.n1 0.155672
R537 VTAIL.n43 VTAIL.n1 0.155672
R538 VTAIL.n64 VTAIL.n63 0.155672
R539 VTAIL.n64 VTAIL.n55 0.155672
R540 VTAIL.n71 VTAIL.n55 0.155672
R541 VTAIL.n72 VTAIL.n71 0.155672
R542 VTAIL.n72 VTAIL.n51 0.155672
R543 VTAIL.n80 VTAIL.n51 0.155672
R544 VTAIL.n81 VTAIL.n80 0.155672
R545 VTAIL.n81 VTAIL.n47 0.155672
R546 VTAIL.n89 VTAIL.n47 0.155672
R547 VTAIL.n110 VTAIL.n109 0.155672
R548 VTAIL.n110 VTAIL.n101 0.155672
R549 VTAIL.n117 VTAIL.n101 0.155672
R550 VTAIL.n118 VTAIL.n117 0.155672
R551 VTAIL.n118 VTAIL.n97 0.155672
R552 VTAIL.n126 VTAIL.n97 0.155672
R553 VTAIL.n127 VTAIL.n126 0.155672
R554 VTAIL.n127 VTAIL.n93 0.155672
R555 VTAIL.n135 VTAIL.n93 0.155672
R556 VTAIL.n319 VTAIL.n277 0.155672
R557 VTAIL.n311 VTAIL.n277 0.155672
R558 VTAIL.n311 VTAIL.n310 0.155672
R559 VTAIL.n310 VTAIL.n281 0.155672
R560 VTAIL.n303 VTAIL.n281 0.155672
R561 VTAIL.n303 VTAIL.n302 0.155672
R562 VTAIL.n302 VTAIL.n286 0.155672
R563 VTAIL.n295 VTAIL.n286 0.155672
R564 VTAIL.n295 VTAIL.n294 0.155672
R565 VTAIL.n273 VTAIL.n231 0.155672
R566 VTAIL.n265 VTAIL.n231 0.155672
R567 VTAIL.n265 VTAIL.n264 0.155672
R568 VTAIL.n264 VTAIL.n235 0.155672
R569 VTAIL.n257 VTAIL.n235 0.155672
R570 VTAIL.n257 VTAIL.n256 0.155672
R571 VTAIL.n256 VTAIL.n240 0.155672
R572 VTAIL.n249 VTAIL.n240 0.155672
R573 VTAIL.n249 VTAIL.n248 0.155672
R574 VTAIL.n227 VTAIL.n185 0.155672
R575 VTAIL.n219 VTAIL.n185 0.155672
R576 VTAIL.n219 VTAIL.n218 0.155672
R577 VTAIL.n218 VTAIL.n189 0.155672
R578 VTAIL.n211 VTAIL.n189 0.155672
R579 VTAIL.n211 VTAIL.n210 0.155672
R580 VTAIL.n210 VTAIL.n194 0.155672
R581 VTAIL.n203 VTAIL.n194 0.155672
R582 VTAIL.n203 VTAIL.n202 0.155672
R583 VTAIL.n181 VTAIL.n139 0.155672
R584 VTAIL.n173 VTAIL.n139 0.155672
R585 VTAIL.n173 VTAIL.n172 0.155672
R586 VTAIL.n172 VTAIL.n143 0.155672
R587 VTAIL.n165 VTAIL.n143 0.155672
R588 VTAIL.n165 VTAIL.n164 0.155672
R589 VTAIL.n164 VTAIL.n148 0.155672
R590 VTAIL.n157 VTAIL.n148 0.155672
R591 VTAIL.n157 VTAIL.n156 0.155672
R592 VDD1 VDD1.n1 122.763
R593 VDD1 VDD1.n0 83.2714
R594 VDD1.n0 VDD1.t1 3.74964
R595 VDD1.n0 VDD1.t3 3.74964
R596 VDD1.n1 VDD1.t0 3.74964
R597 VDD1.n1 VDD1.t2 3.74964
R598 B.n423 B.n60 585
R599 B.n425 B.n424 585
R600 B.n426 B.n59 585
R601 B.n428 B.n427 585
R602 B.n429 B.n58 585
R603 B.n431 B.n430 585
R604 B.n432 B.n57 585
R605 B.n434 B.n433 585
R606 B.n435 B.n56 585
R607 B.n437 B.n436 585
R608 B.n438 B.n55 585
R609 B.n440 B.n439 585
R610 B.n441 B.n54 585
R611 B.n443 B.n442 585
R612 B.n444 B.n53 585
R613 B.n446 B.n445 585
R614 B.n447 B.n52 585
R615 B.n449 B.n448 585
R616 B.n450 B.n51 585
R617 B.n452 B.n451 585
R618 B.n453 B.n50 585
R619 B.n455 B.n454 585
R620 B.n456 B.n49 585
R621 B.n458 B.n457 585
R622 B.n459 B.n48 585
R623 B.n461 B.n460 585
R624 B.n462 B.n47 585
R625 B.n464 B.n463 585
R626 B.n465 B.n46 585
R627 B.n467 B.n466 585
R628 B.n468 B.n45 585
R629 B.n470 B.n469 585
R630 B.n472 B.n471 585
R631 B.n473 B.n41 585
R632 B.n475 B.n474 585
R633 B.n476 B.n40 585
R634 B.n478 B.n477 585
R635 B.n479 B.n39 585
R636 B.n481 B.n480 585
R637 B.n482 B.n38 585
R638 B.n484 B.n483 585
R639 B.n486 B.n35 585
R640 B.n488 B.n487 585
R641 B.n489 B.n34 585
R642 B.n491 B.n490 585
R643 B.n492 B.n33 585
R644 B.n494 B.n493 585
R645 B.n495 B.n32 585
R646 B.n497 B.n496 585
R647 B.n498 B.n31 585
R648 B.n500 B.n499 585
R649 B.n501 B.n30 585
R650 B.n503 B.n502 585
R651 B.n504 B.n29 585
R652 B.n506 B.n505 585
R653 B.n507 B.n28 585
R654 B.n509 B.n508 585
R655 B.n510 B.n27 585
R656 B.n512 B.n511 585
R657 B.n513 B.n26 585
R658 B.n515 B.n514 585
R659 B.n516 B.n25 585
R660 B.n518 B.n517 585
R661 B.n519 B.n24 585
R662 B.n521 B.n520 585
R663 B.n522 B.n23 585
R664 B.n524 B.n523 585
R665 B.n525 B.n22 585
R666 B.n527 B.n526 585
R667 B.n528 B.n21 585
R668 B.n530 B.n529 585
R669 B.n531 B.n20 585
R670 B.n533 B.n532 585
R671 B.n422 B.n421 585
R672 B.n420 B.n61 585
R673 B.n419 B.n418 585
R674 B.n417 B.n62 585
R675 B.n416 B.n415 585
R676 B.n414 B.n63 585
R677 B.n413 B.n412 585
R678 B.n411 B.n64 585
R679 B.n410 B.n409 585
R680 B.n408 B.n65 585
R681 B.n407 B.n406 585
R682 B.n405 B.n66 585
R683 B.n404 B.n403 585
R684 B.n402 B.n67 585
R685 B.n401 B.n400 585
R686 B.n399 B.n68 585
R687 B.n398 B.n397 585
R688 B.n396 B.n69 585
R689 B.n395 B.n394 585
R690 B.n393 B.n70 585
R691 B.n392 B.n391 585
R692 B.n390 B.n71 585
R693 B.n389 B.n388 585
R694 B.n387 B.n72 585
R695 B.n386 B.n385 585
R696 B.n384 B.n73 585
R697 B.n383 B.n382 585
R698 B.n381 B.n74 585
R699 B.n380 B.n379 585
R700 B.n378 B.n75 585
R701 B.n377 B.n376 585
R702 B.n375 B.n76 585
R703 B.n374 B.n373 585
R704 B.n372 B.n77 585
R705 B.n371 B.n370 585
R706 B.n369 B.n78 585
R707 B.n368 B.n367 585
R708 B.n366 B.n79 585
R709 B.n365 B.n364 585
R710 B.n363 B.n80 585
R711 B.n362 B.n361 585
R712 B.n360 B.n81 585
R713 B.n359 B.n358 585
R714 B.n357 B.n82 585
R715 B.n356 B.n355 585
R716 B.n354 B.n83 585
R717 B.n353 B.n352 585
R718 B.n351 B.n84 585
R719 B.n350 B.n349 585
R720 B.n348 B.n85 585
R721 B.n347 B.n346 585
R722 B.n345 B.n86 585
R723 B.n344 B.n343 585
R724 B.n342 B.n87 585
R725 B.n341 B.n340 585
R726 B.n339 B.n88 585
R727 B.n338 B.n337 585
R728 B.n336 B.n89 585
R729 B.n335 B.n334 585
R730 B.n333 B.n90 585
R731 B.n332 B.n331 585
R732 B.n330 B.n91 585
R733 B.n329 B.n328 585
R734 B.n327 B.n92 585
R735 B.n326 B.n325 585
R736 B.n324 B.n93 585
R737 B.n323 B.n322 585
R738 B.n321 B.n94 585
R739 B.n320 B.n319 585
R740 B.n318 B.n95 585
R741 B.n317 B.n316 585
R742 B.n206 B.n205 585
R743 B.n207 B.n136 585
R744 B.n209 B.n208 585
R745 B.n210 B.n135 585
R746 B.n212 B.n211 585
R747 B.n213 B.n134 585
R748 B.n215 B.n214 585
R749 B.n216 B.n133 585
R750 B.n218 B.n217 585
R751 B.n219 B.n132 585
R752 B.n221 B.n220 585
R753 B.n222 B.n131 585
R754 B.n224 B.n223 585
R755 B.n225 B.n130 585
R756 B.n227 B.n226 585
R757 B.n228 B.n129 585
R758 B.n230 B.n229 585
R759 B.n231 B.n128 585
R760 B.n233 B.n232 585
R761 B.n234 B.n127 585
R762 B.n236 B.n235 585
R763 B.n237 B.n126 585
R764 B.n239 B.n238 585
R765 B.n240 B.n125 585
R766 B.n242 B.n241 585
R767 B.n243 B.n124 585
R768 B.n245 B.n244 585
R769 B.n246 B.n123 585
R770 B.n248 B.n247 585
R771 B.n249 B.n122 585
R772 B.n251 B.n250 585
R773 B.n252 B.n119 585
R774 B.n255 B.n254 585
R775 B.n256 B.n118 585
R776 B.n258 B.n257 585
R777 B.n259 B.n117 585
R778 B.n261 B.n260 585
R779 B.n262 B.n116 585
R780 B.n264 B.n263 585
R781 B.n265 B.n115 585
R782 B.n267 B.n266 585
R783 B.n269 B.n268 585
R784 B.n270 B.n111 585
R785 B.n272 B.n271 585
R786 B.n273 B.n110 585
R787 B.n275 B.n274 585
R788 B.n276 B.n109 585
R789 B.n278 B.n277 585
R790 B.n279 B.n108 585
R791 B.n281 B.n280 585
R792 B.n282 B.n107 585
R793 B.n284 B.n283 585
R794 B.n285 B.n106 585
R795 B.n287 B.n286 585
R796 B.n288 B.n105 585
R797 B.n290 B.n289 585
R798 B.n291 B.n104 585
R799 B.n293 B.n292 585
R800 B.n294 B.n103 585
R801 B.n296 B.n295 585
R802 B.n297 B.n102 585
R803 B.n299 B.n298 585
R804 B.n300 B.n101 585
R805 B.n302 B.n301 585
R806 B.n303 B.n100 585
R807 B.n305 B.n304 585
R808 B.n306 B.n99 585
R809 B.n308 B.n307 585
R810 B.n309 B.n98 585
R811 B.n311 B.n310 585
R812 B.n312 B.n97 585
R813 B.n314 B.n313 585
R814 B.n315 B.n96 585
R815 B.n204 B.n137 585
R816 B.n203 B.n202 585
R817 B.n201 B.n138 585
R818 B.n200 B.n199 585
R819 B.n198 B.n139 585
R820 B.n197 B.n196 585
R821 B.n195 B.n140 585
R822 B.n194 B.n193 585
R823 B.n192 B.n141 585
R824 B.n191 B.n190 585
R825 B.n189 B.n142 585
R826 B.n188 B.n187 585
R827 B.n186 B.n143 585
R828 B.n185 B.n184 585
R829 B.n183 B.n144 585
R830 B.n182 B.n181 585
R831 B.n180 B.n145 585
R832 B.n179 B.n178 585
R833 B.n177 B.n146 585
R834 B.n176 B.n175 585
R835 B.n174 B.n147 585
R836 B.n173 B.n172 585
R837 B.n171 B.n148 585
R838 B.n170 B.n169 585
R839 B.n168 B.n149 585
R840 B.n167 B.n166 585
R841 B.n165 B.n150 585
R842 B.n164 B.n163 585
R843 B.n162 B.n151 585
R844 B.n161 B.n160 585
R845 B.n159 B.n152 585
R846 B.n158 B.n157 585
R847 B.n156 B.n153 585
R848 B.n155 B.n154 585
R849 B.n2 B.n0 585
R850 B.n585 B.n1 585
R851 B.n584 B.n583 585
R852 B.n582 B.n3 585
R853 B.n581 B.n580 585
R854 B.n579 B.n4 585
R855 B.n578 B.n577 585
R856 B.n576 B.n5 585
R857 B.n575 B.n574 585
R858 B.n573 B.n6 585
R859 B.n572 B.n571 585
R860 B.n570 B.n7 585
R861 B.n569 B.n568 585
R862 B.n567 B.n8 585
R863 B.n566 B.n565 585
R864 B.n564 B.n9 585
R865 B.n563 B.n562 585
R866 B.n561 B.n10 585
R867 B.n560 B.n559 585
R868 B.n558 B.n11 585
R869 B.n557 B.n556 585
R870 B.n555 B.n12 585
R871 B.n554 B.n553 585
R872 B.n552 B.n13 585
R873 B.n551 B.n550 585
R874 B.n549 B.n14 585
R875 B.n548 B.n547 585
R876 B.n546 B.n15 585
R877 B.n545 B.n544 585
R878 B.n543 B.n16 585
R879 B.n542 B.n541 585
R880 B.n540 B.n17 585
R881 B.n539 B.n538 585
R882 B.n537 B.n18 585
R883 B.n536 B.n535 585
R884 B.n534 B.n19 585
R885 B.n587 B.n586 585
R886 B.n206 B.n137 492.5
R887 B.n532 B.n19 492.5
R888 B.n316 B.n315 492.5
R889 B.n423 B.n422 492.5
R890 B.n112 B.t11 374.464
R891 B.n42 B.t7 374.464
R892 B.n120 B.t5 374.464
R893 B.n36 B.t1 374.464
R894 B.n113 B.t10 315.7
R895 B.n43 B.t8 315.7
R896 B.n121 B.t4 315.7
R897 B.n37 B.t2 315.7
R898 B.n112 B.t9 285.58
R899 B.n120 B.t3 285.58
R900 B.n36 B.t0 285.58
R901 B.n42 B.t6 285.58
R902 B.n202 B.n137 163.367
R903 B.n202 B.n201 163.367
R904 B.n201 B.n200 163.367
R905 B.n200 B.n139 163.367
R906 B.n196 B.n139 163.367
R907 B.n196 B.n195 163.367
R908 B.n195 B.n194 163.367
R909 B.n194 B.n141 163.367
R910 B.n190 B.n141 163.367
R911 B.n190 B.n189 163.367
R912 B.n189 B.n188 163.367
R913 B.n188 B.n143 163.367
R914 B.n184 B.n143 163.367
R915 B.n184 B.n183 163.367
R916 B.n183 B.n182 163.367
R917 B.n182 B.n145 163.367
R918 B.n178 B.n145 163.367
R919 B.n178 B.n177 163.367
R920 B.n177 B.n176 163.367
R921 B.n176 B.n147 163.367
R922 B.n172 B.n147 163.367
R923 B.n172 B.n171 163.367
R924 B.n171 B.n170 163.367
R925 B.n170 B.n149 163.367
R926 B.n166 B.n149 163.367
R927 B.n166 B.n165 163.367
R928 B.n165 B.n164 163.367
R929 B.n164 B.n151 163.367
R930 B.n160 B.n151 163.367
R931 B.n160 B.n159 163.367
R932 B.n159 B.n158 163.367
R933 B.n158 B.n153 163.367
R934 B.n154 B.n153 163.367
R935 B.n154 B.n2 163.367
R936 B.n586 B.n2 163.367
R937 B.n586 B.n585 163.367
R938 B.n585 B.n584 163.367
R939 B.n584 B.n3 163.367
R940 B.n580 B.n3 163.367
R941 B.n580 B.n579 163.367
R942 B.n579 B.n578 163.367
R943 B.n578 B.n5 163.367
R944 B.n574 B.n5 163.367
R945 B.n574 B.n573 163.367
R946 B.n573 B.n572 163.367
R947 B.n572 B.n7 163.367
R948 B.n568 B.n7 163.367
R949 B.n568 B.n567 163.367
R950 B.n567 B.n566 163.367
R951 B.n566 B.n9 163.367
R952 B.n562 B.n9 163.367
R953 B.n562 B.n561 163.367
R954 B.n561 B.n560 163.367
R955 B.n560 B.n11 163.367
R956 B.n556 B.n11 163.367
R957 B.n556 B.n555 163.367
R958 B.n555 B.n554 163.367
R959 B.n554 B.n13 163.367
R960 B.n550 B.n13 163.367
R961 B.n550 B.n549 163.367
R962 B.n549 B.n548 163.367
R963 B.n548 B.n15 163.367
R964 B.n544 B.n15 163.367
R965 B.n544 B.n543 163.367
R966 B.n543 B.n542 163.367
R967 B.n542 B.n17 163.367
R968 B.n538 B.n17 163.367
R969 B.n538 B.n537 163.367
R970 B.n537 B.n536 163.367
R971 B.n536 B.n19 163.367
R972 B.n207 B.n206 163.367
R973 B.n208 B.n207 163.367
R974 B.n208 B.n135 163.367
R975 B.n212 B.n135 163.367
R976 B.n213 B.n212 163.367
R977 B.n214 B.n213 163.367
R978 B.n214 B.n133 163.367
R979 B.n218 B.n133 163.367
R980 B.n219 B.n218 163.367
R981 B.n220 B.n219 163.367
R982 B.n220 B.n131 163.367
R983 B.n224 B.n131 163.367
R984 B.n225 B.n224 163.367
R985 B.n226 B.n225 163.367
R986 B.n226 B.n129 163.367
R987 B.n230 B.n129 163.367
R988 B.n231 B.n230 163.367
R989 B.n232 B.n231 163.367
R990 B.n232 B.n127 163.367
R991 B.n236 B.n127 163.367
R992 B.n237 B.n236 163.367
R993 B.n238 B.n237 163.367
R994 B.n238 B.n125 163.367
R995 B.n242 B.n125 163.367
R996 B.n243 B.n242 163.367
R997 B.n244 B.n243 163.367
R998 B.n244 B.n123 163.367
R999 B.n248 B.n123 163.367
R1000 B.n249 B.n248 163.367
R1001 B.n250 B.n249 163.367
R1002 B.n250 B.n119 163.367
R1003 B.n255 B.n119 163.367
R1004 B.n256 B.n255 163.367
R1005 B.n257 B.n256 163.367
R1006 B.n257 B.n117 163.367
R1007 B.n261 B.n117 163.367
R1008 B.n262 B.n261 163.367
R1009 B.n263 B.n262 163.367
R1010 B.n263 B.n115 163.367
R1011 B.n267 B.n115 163.367
R1012 B.n268 B.n267 163.367
R1013 B.n268 B.n111 163.367
R1014 B.n272 B.n111 163.367
R1015 B.n273 B.n272 163.367
R1016 B.n274 B.n273 163.367
R1017 B.n274 B.n109 163.367
R1018 B.n278 B.n109 163.367
R1019 B.n279 B.n278 163.367
R1020 B.n280 B.n279 163.367
R1021 B.n280 B.n107 163.367
R1022 B.n284 B.n107 163.367
R1023 B.n285 B.n284 163.367
R1024 B.n286 B.n285 163.367
R1025 B.n286 B.n105 163.367
R1026 B.n290 B.n105 163.367
R1027 B.n291 B.n290 163.367
R1028 B.n292 B.n291 163.367
R1029 B.n292 B.n103 163.367
R1030 B.n296 B.n103 163.367
R1031 B.n297 B.n296 163.367
R1032 B.n298 B.n297 163.367
R1033 B.n298 B.n101 163.367
R1034 B.n302 B.n101 163.367
R1035 B.n303 B.n302 163.367
R1036 B.n304 B.n303 163.367
R1037 B.n304 B.n99 163.367
R1038 B.n308 B.n99 163.367
R1039 B.n309 B.n308 163.367
R1040 B.n310 B.n309 163.367
R1041 B.n310 B.n97 163.367
R1042 B.n314 B.n97 163.367
R1043 B.n315 B.n314 163.367
R1044 B.n316 B.n95 163.367
R1045 B.n320 B.n95 163.367
R1046 B.n321 B.n320 163.367
R1047 B.n322 B.n321 163.367
R1048 B.n322 B.n93 163.367
R1049 B.n326 B.n93 163.367
R1050 B.n327 B.n326 163.367
R1051 B.n328 B.n327 163.367
R1052 B.n328 B.n91 163.367
R1053 B.n332 B.n91 163.367
R1054 B.n333 B.n332 163.367
R1055 B.n334 B.n333 163.367
R1056 B.n334 B.n89 163.367
R1057 B.n338 B.n89 163.367
R1058 B.n339 B.n338 163.367
R1059 B.n340 B.n339 163.367
R1060 B.n340 B.n87 163.367
R1061 B.n344 B.n87 163.367
R1062 B.n345 B.n344 163.367
R1063 B.n346 B.n345 163.367
R1064 B.n346 B.n85 163.367
R1065 B.n350 B.n85 163.367
R1066 B.n351 B.n350 163.367
R1067 B.n352 B.n351 163.367
R1068 B.n352 B.n83 163.367
R1069 B.n356 B.n83 163.367
R1070 B.n357 B.n356 163.367
R1071 B.n358 B.n357 163.367
R1072 B.n358 B.n81 163.367
R1073 B.n362 B.n81 163.367
R1074 B.n363 B.n362 163.367
R1075 B.n364 B.n363 163.367
R1076 B.n364 B.n79 163.367
R1077 B.n368 B.n79 163.367
R1078 B.n369 B.n368 163.367
R1079 B.n370 B.n369 163.367
R1080 B.n370 B.n77 163.367
R1081 B.n374 B.n77 163.367
R1082 B.n375 B.n374 163.367
R1083 B.n376 B.n375 163.367
R1084 B.n376 B.n75 163.367
R1085 B.n380 B.n75 163.367
R1086 B.n381 B.n380 163.367
R1087 B.n382 B.n381 163.367
R1088 B.n382 B.n73 163.367
R1089 B.n386 B.n73 163.367
R1090 B.n387 B.n386 163.367
R1091 B.n388 B.n387 163.367
R1092 B.n388 B.n71 163.367
R1093 B.n392 B.n71 163.367
R1094 B.n393 B.n392 163.367
R1095 B.n394 B.n393 163.367
R1096 B.n394 B.n69 163.367
R1097 B.n398 B.n69 163.367
R1098 B.n399 B.n398 163.367
R1099 B.n400 B.n399 163.367
R1100 B.n400 B.n67 163.367
R1101 B.n404 B.n67 163.367
R1102 B.n405 B.n404 163.367
R1103 B.n406 B.n405 163.367
R1104 B.n406 B.n65 163.367
R1105 B.n410 B.n65 163.367
R1106 B.n411 B.n410 163.367
R1107 B.n412 B.n411 163.367
R1108 B.n412 B.n63 163.367
R1109 B.n416 B.n63 163.367
R1110 B.n417 B.n416 163.367
R1111 B.n418 B.n417 163.367
R1112 B.n418 B.n61 163.367
R1113 B.n422 B.n61 163.367
R1114 B.n532 B.n531 163.367
R1115 B.n531 B.n530 163.367
R1116 B.n530 B.n21 163.367
R1117 B.n526 B.n21 163.367
R1118 B.n526 B.n525 163.367
R1119 B.n525 B.n524 163.367
R1120 B.n524 B.n23 163.367
R1121 B.n520 B.n23 163.367
R1122 B.n520 B.n519 163.367
R1123 B.n519 B.n518 163.367
R1124 B.n518 B.n25 163.367
R1125 B.n514 B.n25 163.367
R1126 B.n514 B.n513 163.367
R1127 B.n513 B.n512 163.367
R1128 B.n512 B.n27 163.367
R1129 B.n508 B.n27 163.367
R1130 B.n508 B.n507 163.367
R1131 B.n507 B.n506 163.367
R1132 B.n506 B.n29 163.367
R1133 B.n502 B.n29 163.367
R1134 B.n502 B.n501 163.367
R1135 B.n501 B.n500 163.367
R1136 B.n500 B.n31 163.367
R1137 B.n496 B.n31 163.367
R1138 B.n496 B.n495 163.367
R1139 B.n495 B.n494 163.367
R1140 B.n494 B.n33 163.367
R1141 B.n490 B.n33 163.367
R1142 B.n490 B.n489 163.367
R1143 B.n489 B.n488 163.367
R1144 B.n488 B.n35 163.367
R1145 B.n483 B.n35 163.367
R1146 B.n483 B.n482 163.367
R1147 B.n482 B.n481 163.367
R1148 B.n481 B.n39 163.367
R1149 B.n477 B.n39 163.367
R1150 B.n477 B.n476 163.367
R1151 B.n476 B.n475 163.367
R1152 B.n475 B.n41 163.367
R1153 B.n471 B.n41 163.367
R1154 B.n471 B.n470 163.367
R1155 B.n470 B.n45 163.367
R1156 B.n466 B.n45 163.367
R1157 B.n466 B.n465 163.367
R1158 B.n465 B.n464 163.367
R1159 B.n464 B.n47 163.367
R1160 B.n460 B.n47 163.367
R1161 B.n460 B.n459 163.367
R1162 B.n459 B.n458 163.367
R1163 B.n458 B.n49 163.367
R1164 B.n454 B.n49 163.367
R1165 B.n454 B.n453 163.367
R1166 B.n453 B.n452 163.367
R1167 B.n452 B.n51 163.367
R1168 B.n448 B.n51 163.367
R1169 B.n448 B.n447 163.367
R1170 B.n447 B.n446 163.367
R1171 B.n446 B.n53 163.367
R1172 B.n442 B.n53 163.367
R1173 B.n442 B.n441 163.367
R1174 B.n441 B.n440 163.367
R1175 B.n440 B.n55 163.367
R1176 B.n436 B.n55 163.367
R1177 B.n436 B.n435 163.367
R1178 B.n435 B.n434 163.367
R1179 B.n434 B.n57 163.367
R1180 B.n430 B.n57 163.367
R1181 B.n430 B.n429 163.367
R1182 B.n429 B.n428 163.367
R1183 B.n428 B.n59 163.367
R1184 B.n424 B.n59 163.367
R1185 B.n424 B.n423 163.367
R1186 B.n114 B.n113 59.5399
R1187 B.n253 B.n121 59.5399
R1188 B.n485 B.n37 59.5399
R1189 B.n44 B.n43 59.5399
R1190 B.n113 B.n112 58.7641
R1191 B.n121 B.n120 58.7641
R1192 B.n37 B.n36 58.7641
R1193 B.n43 B.n42 58.7641
R1194 B.n534 B.n533 32.0005
R1195 B.n421 B.n60 32.0005
R1196 B.n317 B.n96 32.0005
R1197 B.n205 B.n204 32.0005
R1198 B B.n587 18.0485
R1199 B.n533 B.n20 10.6151
R1200 B.n529 B.n20 10.6151
R1201 B.n529 B.n528 10.6151
R1202 B.n528 B.n527 10.6151
R1203 B.n527 B.n22 10.6151
R1204 B.n523 B.n22 10.6151
R1205 B.n523 B.n522 10.6151
R1206 B.n522 B.n521 10.6151
R1207 B.n521 B.n24 10.6151
R1208 B.n517 B.n24 10.6151
R1209 B.n517 B.n516 10.6151
R1210 B.n516 B.n515 10.6151
R1211 B.n515 B.n26 10.6151
R1212 B.n511 B.n26 10.6151
R1213 B.n511 B.n510 10.6151
R1214 B.n510 B.n509 10.6151
R1215 B.n509 B.n28 10.6151
R1216 B.n505 B.n28 10.6151
R1217 B.n505 B.n504 10.6151
R1218 B.n504 B.n503 10.6151
R1219 B.n503 B.n30 10.6151
R1220 B.n499 B.n30 10.6151
R1221 B.n499 B.n498 10.6151
R1222 B.n498 B.n497 10.6151
R1223 B.n497 B.n32 10.6151
R1224 B.n493 B.n32 10.6151
R1225 B.n493 B.n492 10.6151
R1226 B.n492 B.n491 10.6151
R1227 B.n491 B.n34 10.6151
R1228 B.n487 B.n34 10.6151
R1229 B.n487 B.n486 10.6151
R1230 B.n484 B.n38 10.6151
R1231 B.n480 B.n38 10.6151
R1232 B.n480 B.n479 10.6151
R1233 B.n479 B.n478 10.6151
R1234 B.n478 B.n40 10.6151
R1235 B.n474 B.n40 10.6151
R1236 B.n474 B.n473 10.6151
R1237 B.n473 B.n472 10.6151
R1238 B.n469 B.n468 10.6151
R1239 B.n468 B.n467 10.6151
R1240 B.n467 B.n46 10.6151
R1241 B.n463 B.n46 10.6151
R1242 B.n463 B.n462 10.6151
R1243 B.n462 B.n461 10.6151
R1244 B.n461 B.n48 10.6151
R1245 B.n457 B.n48 10.6151
R1246 B.n457 B.n456 10.6151
R1247 B.n456 B.n455 10.6151
R1248 B.n455 B.n50 10.6151
R1249 B.n451 B.n50 10.6151
R1250 B.n451 B.n450 10.6151
R1251 B.n450 B.n449 10.6151
R1252 B.n449 B.n52 10.6151
R1253 B.n445 B.n52 10.6151
R1254 B.n445 B.n444 10.6151
R1255 B.n444 B.n443 10.6151
R1256 B.n443 B.n54 10.6151
R1257 B.n439 B.n54 10.6151
R1258 B.n439 B.n438 10.6151
R1259 B.n438 B.n437 10.6151
R1260 B.n437 B.n56 10.6151
R1261 B.n433 B.n56 10.6151
R1262 B.n433 B.n432 10.6151
R1263 B.n432 B.n431 10.6151
R1264 B.n431 B.n58 10.6151
R1265 B.n427 B.n58 10.6151
R1266 B.n427 B.n426 10.6151
R1267 B.n426 B.n425 10.6151
R1268 B.n425 B.n60 10.6151
R1269 B.n318 B.n317 10.6151
R1270 B.n319 B.n318 10.6151
R1271 B.n319 B.n94 10.6151
R1272 B.n323 B.n94 10.6151
R1273 B.n324 B.n323 10.6151
R1274 B.n325 B.n324 10.6151
R1275 B.n325 B.n92 10.6151
R1276 B.n329 B.n92 10.6151
R1277 B.n330 B.n329 10.6151
R1278 B.n331 B.n330 10.6151
R1279 B.n331 B.n90 10.6151
R1280 B.n335 B.n90 10.6151
R1281 B.n336 B.n335 10.6151
R1282 B.n337 B.n336 10.6151
R1283 B.n337 B.n88 10.6151
R1284 B.n341 B.n88 10.6151
R1285 B.n342 B.n341 10.6151
R1286 B.n343 B.n342 10.6151
R1287 B.n343 B.n86 10.6151
R1288 B.n347 B.n86 10.6151
R1289 B.n348 B.n347 10.6151
R1290 B.n349 B.n348 10.6151
R1291 B.n349 B.n84 10.6151
R1292 B.n353 B.n84 10.6151
R1293 B.n354 B.n353 10.6151
R1294 B.n355 B.n354 10.6151
R1295 B.n355 B.n82 10.6151
R1296 B.n359 B.n82 10.6151
R1297 B.n360 B.n359 10.6151
R1298 B.n361 B.n360 10.6151
R1299 B.n361 B.n80 10.6151
R1300 B.n365 B.n80 10.6151
R1301 B.n366 B.n365 10.6151
R1302 B.n367 B.n366 10.6151
R1303 B.n367 B.n78 10.6151
R1304 B.n371 B.n78 10.6151
R1305 B.n372 B.n371 10.6151
R1306 B.n373 B.n372 10.6151
R1307 B.n373 B.n76 10.6151
R1308 B.n377 B.n76 10.6151
R1309 B.n378 B.n377 10.6151
R1310 B.n379 B.n378 10.6151
R1311 B.n379 B.n74 10.6151
R1312 B.n383 B.n74 10.6151
R1313 B.n384 B.n383 10.6151
R1314 B.n385 B.n384 10.6151
R1315 B.n385 B.n72 10.6151
R1316 B.n389 B.n72 10.6151
R1317 B.n390 B.n389 10.6151
R1318 B.n391 B.n390 10.6151
R1319 B.n391 B.n70 10.6151
R1320 B.n395 B.n70 10.6151
R1321 B.n396 B.n395 10.6151
R1322 B.n397 B.n396 10.6151
R1323 B.n397 B.n68 10.6151
R1324 B.n401 B.n68 10.6151
R1325 B.n402 B.n401 10.6151
R1326 B.n403 B.n402 10.6151
R1327 B.n403 B.n66 10.6151
R1328 B.n407 B.n66 10.6151
R1329 B.n408 B.n407 10.6151
R1330 B.n409 B.n408 10.6151
R1331 B.n409 B.n64 10.6151
R1332 B.n413 B.n64 10.6151
R1333 B.n414 B.n413 10.6151
R1334 B.n415 B.n414 10.6151
R1335 B.n415 B.n62 10.6151
R1336 B.n419 B.n62 10.6151
R1337 B.n420 B.n419 10.6151
R1338 B.n421 B.n420 10.6151
R1339 B.n205 B.n136 10.6151
R1340 B.n209 B.n136 10.6151
R1341 B.n210 B.n209 10.6151
R1342 B.n211 B.n210 10.6151
R1343 B.n211 B.n134 10.6151
R1344 B.n215 B.n134 10.6151
R1345 B.n216 B.n215 10.6151
R1346 B.n217 B.n216 10.6151
R1347 B.n217 B.n132 10.6151
R1348 B.n221 B.n132 10.6151
R1349 B.n222 B.n221 10.6151
R1350 B.n223 B.n222 10.6151
R1351 B.n223 B.n130 10.6151
R1352 B.n227 B.n130 10.6151
R1353 B.n228 B.n227 10.6151
R1354 B.n229 B.n228 10.6151
R1355 B.n229 B.n128 10.6151
R1356 B.n233 B.n128 10.6151
R1357 B.n234 B.n233 10.6151
R1358 B.n235 B.n234 10.6151
R1359 B.n235 B.n126 10.6151
R1360 B.n239 B.n126 10.6151
R1361 B.n240 B.n239 10.6151
R1362 B.n241 B.n240 10.6151
R1363 B.n241 B.n124 10.6151
R1364 B.n245 B.n124 10.6151
R1365 B.n246 B.n245 10.6151
R1366 B.n247 B.n246 10.6151
R1367 B.n247 B.n122 10.6151
R1368 B.n251 B.n122 10.6151
R1369 B.n252 B.n251 10.6151
R1370 B.n254 B.n118 10.6151
R1371 B.n258 B.n118 10.6151
R1372 B.n259 B.n258 10.6151
R1373 B.n260 B.n259 10.6151
R1374 B.n260 B.n116 10.6151
R1375 B.n264 B.n116 10.6151
R1376 B.n265 B.n264 10.6151
R1377 B.n266 B.n265 10.6151
R1378 B.n270 B.n269 10.6151
R1379 B.n271 B.n270 10.6151
R1380 B.n271 B.n110 10.6151
R1381 B.n275 B.n110 10.6151
R1382 B.n276 B.n275 10.6151
R1383 B.n277 B.n276 10.6151
R1384 B.n277 B.n108 10.6151
R1385 B.n281 B.n108 10.6151
R1386 B.n282 B.n281 10.6151
R1387 B.n283 B.n282 10.6151
R1388 B.n283 B.n106 10.6151
R1389 B.n287 B.n106 10.6151
R1390 B.n288 B.n287 10.6151
R1391 B.n289 B.n288 10.6151
R1392 B.n289 B.n104 10.6151
R1393 B.n293 B.n104 10.6151
R1394 B.n294 B.n293 10.6151
R1395 B.n295 B.n294 10.6151
R1396 B.n295 B.n102 10.6151
R1397 B.n299 B.n102 10.6151
R1398 B.n300 B.n299 10.6151
R1399 B.n301 B.n300 10.6151
R1400 B.n301 B.n100 10.6151
R1401 B.n305 B.n100 10.6151
R1402 B.n306 B.n305 10.6151
R1403 B.n307 B.n306 10.6151
R1404 B.n307 B.n98 10.6151
R1405 B.n311 B.n98 10.6151
R1406 B.n312 B.n311 10.6151
R1407 B.n313 B.n312 10.6151
R1408 B.n313 B.n96 10.6151
R1409 B.n204 B.n203 10.6151
R1410 B.n203 B.n138 10.6151
R1411 B.n199 B.n138 10.6151
R1412 B.n199 B.n198 10.6151
R1413 B.n198 B.n197 10.6151
R1414 B.n197 B.n140 10.6151
R1415 B.n193 B.n140 10.6151
R1416 B.n193 B.n192 10.6151
R1417 B.n192 B.n191 10.6151
R1418 B.n191 B.n142 10.6151
R1419 B.n187 B.n142 10.6151
R1420 B.n187 B.n186 10.6151
R1421 B.n186 B.n185 10.6151
R1422 B.n185 B.n144 10.6151
R1423 B.n181 B.n144 10.6151
R1424 B.n181 B.n180 10.6151
R1425 B.n180 B.n179 10.6151
R1426 B.n179 B.n146 10.6151
R1427 B.n175 B.n146 10.6151
R1428 B.n175 B.n174 10.6151
R1429 B.n174 B.n173 10.6151
R1430 B.n173 B.n148 10.6151
R1431 B.n169 B.n148 10.6151
R1432 B.n169 B.n168 10.6151
R1433 B.n168 B.n167 10.6151
R1434 B.n167 B.n150 10.6151
R1435 B.n163 B.n150 10.6151
R1436 B.n163 B.n162 10.6151
R1437 B.n162 B.n161 10.6151
R1438 B.n161 B.n152 10.6151
R1439 B.n157 B.n152 10.6151
R1440 B.n157 B.n156 10.6151
R1441 B.n156 B.n155 10.6151
R1442 B.n155 B.n0 10.6151
R1443 B.n583 B.n1 10.6151
R1444 B.n583 B.n582 10.6151
R1445 B.n582 B.n581 10.6151
R1446 B.n581 B.n4 10.6151
R1447 B.n577 B.n4 10.6151
R1448 B.n577 B.n576 10.6151
R1449 B.n576 B.n575 10.6151
R1450 B.n575 B.n6 10.6151
R1451 B.n571 B.n6 10.6151
R1452 B.n571 B.n570 10.6151
R1453 B.n570 B.n569 10.6151
R1454 B.n569 B.n8 10.6151
R1455 B.n565 B.n8 10.6151
R1456 B.n565 B.n564 10.6151
R1457 B.n564 B.n563 10.6151
R1458 B.n563 B.n10 10.6151
R1459 B.n559 B.n10 10.6151
R1460 B.n559 B.n558 10.6151
R1461 B.n558 B.n557 10.6151
R1462 B.n557 B.n12 10.6151
R1463 B.n553 B.n12 10.6151
R1464 B.n553 B.n552 10.6151
R1465 B.n552 B.n551 10.6151
R1466 B.n551 B.n14 10.6151
R1467 B.n547 B.n14 10.6151
R1468 B.n547 B.n546 10.6151
R1469 B.n546 B.n545 10.6151
R1470 B.n545 B.n16 10.6151
R1471 B.n541 B.n16 10.6151
R1472 B.n541 B.n540 10.6151
R1473 B.n540 B.n539 10.6151
R1474 B.n539 B.n18 10.6151
R1475 B.n535 B.n18 10.6151
R1476 B.n535 B.n534 10.6151
R1477 B.n485 B.n484 6.5566
R1478 B.n472 B.n44 6.5566
R1479 B.n254 B.n253 6.5566
R1480 B.n266 B.n114 6.5566
R1481 B.n486 B.n485 4.05904
R1482 B.n469 B.n44 4.05904
R1483 B.n253 B.n252 4.05904
R1484 B.n269 B.n114 4.05904
R1485 B.n587 B.n0 2.81026
R1486 B.n587 B.n1 2.81026
R1487 VN.n0 VN.t0 111.403
R1488 VN.n1 VN.t1 111.403
R1489 VN.n0 VN.t3 110.531
R1490 VN.n1 VN.t2 110.531
R1491 VN VN.n1 47.9295
R1492 VN VN.n0 3.65294
R1493 VDD2.n2 VDD2.n0 122.239
R1494 VDD2.n2 VDD2.n1 83.2132
R1495 VDD2.n1 VDD2.t1 3.74964
R1496 VDD2.n1 VDD2.t2 3.74964
R1497 VDD2.n0 VDD2.t3 3.74964
R1498 VDD2.n0 VDD2.t0 3.74964
R1499 VDD2 VDD2.n2 0.0586897
C0 VDD1 VTAIL 4.64393f
C1 B VTAIL 3.89198f
C2 VDD1 VN 0.148926f
C3 B VN 1.08855f
C4 VDD2 VP 0.400505f
C5 VP VTAIL 3.62839f
C6 VP VN 5.64967f
C7 VDD2 VTAIL 4.69881f
C8 w_n2788_n2702# VDD1 1.38059f
C9 B w_n2788_n2702# 8.435619f
C10 VDD2 VN 3.54655f
C11 VN VTAIL 3.61428f
C12 w_n2788_n2702# VP 5.04722f
C13 B VDD1 1.18887f
C14 VDD2 w_n2788_n2702# 1.43893f
C15 w_n2788_n2702# VTAIL 3.23191f
C16 w_n2788_n2702# VN 4.68856f
C17 VDD1 VP 3.79736f
C18 B VP 1.6842f
C19 VDD2 VDD1 1.044f
C20 VDD2 B 1.24267f
C21 VDD2 VSUBS 0.889501f
C22 VDD1 VSUBS 5.34882f
C23 VTAIL VSUBS 1.072606f
C24 VN VSUBS 5.422151f
C25 VP VSUBS 2.206399f
C26 B VSUBS 4.082099f
C27 w_n2788_n2702# VSUBS 93.3088f
C28 VDD2.t3 VSUBS 0.185547f
C29 VDD2.t0 VSUBS 0.185547f
C30 VDD2.n0 VSUBS 1.91616f
C31 VDD2.t1 VSUBS 0.185547f
C32 VDD2.t2 VSUBS 0.185547f
C33 VDD2.n1 VSUBS 1.36895f
C34 VDD2.n2 VSUBS 3.93893f
C35 VN.t0 VSUBS 2.5478f
C36 VN.t3 VSUBS 2.5398f
C37 VN.n0 VSUBS 1.61782f
C38 VN.t1 VSUBS 2.5478f
C39 VN.t2 VSUBS 2.5398f
C40 VN.n1 VSUBS 3.44715f
C41 B.n0 VSUBS 0.004626f
C42 B.n1 VSUBS 0.004626f
C43 B.n2 VSUBS 0.007316f
C44 B.n3 VSUBS 0.007316f
C45 B.n4 VSUBS 0.007316f
C46 B.n5 VSUBS 0.007316f
C47 B.n6 VSUBS 0.007316f
C48 B.n7 VSUBS 0.007316f
C49 B.n8 VSUBS 0.007316f
C50 B.n9 VSUBS 0.007316f
C51 B.n10 VSUBS 0.007316f
C52 B.n11 VSUBS 0.007316f
C53 B.n12 VSUBS 0.007316f
C54 B.n13 VSUBS 0.007316f
C55 B.n14 VSUBS 0.007316f
C56 B.n15 VSUBS 0.007316f
C57 B.n16 VSUBS 0.007316f
C58 B.n17 VSUBS 0.007316f
C59 B.n18 VSUBS 0.007316f
C60 B.n19 VSUBS 0.016664f
C61 B.n20 VSUBS 0.007316f
C62 B.n21 VSUBS 0.007316f
C63 B.n22 VSUBS 0.007316f
C64 B.n23 VSUBS 0.007316f
C65 B.n24 VSUBS 0.007316f
C66 B.n25 VSUBS 0.007316f
C67 B.n26 VSUBS 0.007316f
C68 B.n27 VSUBS 0.007316f
C69 B.n28 VSUBS 0.007316f
C70 B.n29 VSUBS 0.007316f
C71 B.n30 VSUBS 0.007316f
C72 B.n31 VSUBS 0.007316f
C73 B.n32 VSUBS 0.007316f
C74 B.n33 VSUBS 0.007316f
C75 B.n34 VSUBS 0.007316f
C76 B.n35 VSUBS 0.007316f
C77 B.t2 VSUBS 0.146301f
C78 B.t1 VSUBS 0.177938f
C79 B.t0 VSUBS 1.13822f
C80 B.n36 VSUBS 0.292182f
C81 B.n37 VSUBS 0.212036f
C82 B.n38 VSUBS 0.007316f
C83 B.n39 VSUBS 0.007316f
C84 B.n40 VSUBS 0.007316f
C85 B.n41 VSUBS 0.007316f
C86 B.t8 VSUBS 0.146304f
C87 B.t7 VSUBS 0.17794f
C88 B.t6 VSUBS 1.13822f
C89 B.n42 VSUBS 0.29218f
C90 B.n43 VSUBS 0.212033f
C91 B.n44 VSUBS 0.016949f
C92 B.n45 VSUBS 0.007316f
C93 B.n46 VSUBS 0.007316f
C94 B.n47 VSUBS 0.007316f
C95 B.n48 VSUBS 0.007316f
C96 B.n49 VSUBS 0.007316f
C97 B.n50 VSUBS 0.007316f
C98 B.n51 VSUBS 0.007316f
C99 B.n52 VSUBS 0.007316f
C100 B.n53 VSUBS 0.007316f
C101 B.n54 VSUBS 0.007316f
C102 B.n55 VSUBS 0.007316f
C103 B.n56 VSUBS 0.007316f
C104 B.n57 VSUBS 0.007316f
C105 B.n58 VSUBS 0.007316f
C106 B.n59 VSUBS 0.007316f
C107 B.n60 VSUBS 0.016234f
C108 B.n61 VSUBS 0.007316f
C109 B.n62 VSUBS 0.007316f
C110 B.n63 VSUBS 0.007316f
C111 B.n64 VSUBS 0.007316f
C112 B.n65 VSUBS 0.007316f
C113 B.n66 VSUBS 0.007316f
C114 B.n67 VSUBS 0.007316f
C115 B.n68 VSUBS 0.007316f
C116 B.n69 VSUBS 0.007316f
C117 B.n70 VSUBS 0.007316f
C118 B.n71 VSUBS 0.007316f
C119 B.n72 VSUBS 0.007316f
C120 B.n73 VSUBS 0.007316f
C121 B.n74 VSUBS 0.007316f
C122 B.n75 VSUBS 0.007316f
C123 B.n76 VSUBS 0.007316f
C124 B.n77 VSUBS 0.007316f
C125 B.n78 VSUBS 0.007316f
C126 B.n79 VSUBS 0.007316f
C127 B.n80 VSUBS 0.007316f
C128 B.n81 VSUBS 0.007316f
C129 B.n82 VSUBS 0.007316f
C130 B.n83 VSUBS 0.007316f
C131 B.n84 VSUBS 0.007316f
C132 B.n85 VSUBS 0.007316f
C133 B.n86 VSUBS 0.007316f
C134 B.n87 VSUBS 0.007316f
C135 B.n88 VSUBS 0.007316f
C136 B.n89 VSUBS 0.007316f
C137 B.n90 VSUBS 0.007316f
C138 B.n91 VSUBS 0.007316f
C139 B.n92 VSUBS 0.007316f
C140 B.n93 VSUBS 0.007316f
C141 B.n94 VSUBS 0.007316f
C142 B.n95 VSUBS 0.007316f
C143 B.n96 VSUBS 0.017116f
C144 B.n97 VSUBS 0.007316f
C145 B.n98 VSUBS 0.007316f
C146 B.n99 VSUBS 0.007316f
C147 B.n100 VSUBS 0.007316f
C148 B.n101 VSUBS 0.007316f
C149 B.n102 VSUBS 0.007316f
C150 B.n103 VSUBS 0.007316f
C151 B.n104 VSUBS 0.007316f
C152 B.n105 VSUBS 0.007316f
C153 B.n106 VSUBS 0.007316f
C154 B.n107 VSUBS 0.007316f
C155 B.n108 VSUBS 0.007316f
C156 B.n109 VSUBS 0.007316f
C157 B.n110 VSUBS 0.007316f
C158 B.n111 VSUBS 0.007316f
C159 B.t10 VSUBS 0.146304f
C160 B.t11 VSUBS 0.17794f
C161 B.t9 VSUBS 1.13822f
C162 B.n112 VSUBS 0.29218f
C163 B.n113 VSUBS 0.212033f
C164 B.n114 VSUBS 0.016949f
C165 B.n115 VSUBS 0.007316f
C166 B.n116 VSUBS 0.007316f
C167 B.n117 VSUBS 0.007316f
C168 B.n118 VSUBS 0.007316f
C169 B.n119 VSUBS 0.007316f
C170 B.t4 VSUBS 0.146301f
C171 B.t5 VSUBS 0.177938f
C172 B.t3 VSUBS 1.13822f
C173 B.n120 VSUBS 0.292182f
C174 B.n121 VSUBS 0.212036f
C175 B.n122 VSUBS 0.007316f
C176 B.n123 VSUBS 0.007316f
C177 B.n124 VSUBS 0.007316f
C178 B.n125 VSUBS 0.007316f
C179 B.n126 VSUBS 0.007316f
C180 B.n127 VSUBS 0.007316f
C181 B.n128 VSUBS 0.007316f
C182 B.n129 VSUBS 0.007316f
C183 B.n130 VSUBS 0.007316f
C184 B.n131 VSUBS 0.007316f
C185 B.n132 VSUBS 0.007316f
C186 B.n133 VSUBS 0.007316f
C187 B.n134 VSUBS 0.007316f
C188 B.n135 VSUBS 0.007316f
C189 B.n136 VSUBS 0.007316f
C190 B.n137 VSUBS 0.016664f
C191 B.n138 VSUBS 0.007316f
C192 B.n139 VSUBS 0.007316f
C193 B.n140 VSUBS 0.007316f
C194 B.n141 VSUBS 0.007316f
C195 B.n142 VSUBS 0.007316f
C196 B.n143 VSUBS 0.007316f
C197 B.n144 VSUBS 0.007316f
C198 B.n145 VSUBS 0.007316f
C199 B.n146 VSUBS 0.007316f
C200 B.n147 VSUBS 0.007316f
C201 B.n148 VSUBS 0.007316f
C202 B.n149 VSUBS 0.007316f
C203 B.n150 VSUBS 0.007316f
C204 B.n151 VSUBS 0.007316f
C205 B.n152 VSUBS 0.007316f
C206 B.n153 VSUBS 0.007316f
C207 B.n154 VSUBS 0.007316f
C208 B.n155 VSUBS 0.007316f
C209 B.n156 VSUBS 0.007316f
C210 B.n157 VSUBS 0.007316f
C211 B.n158 VSUBS 0.007316f
C212 B.n159 VSUBS 0.007316f
C213 B.n160 VSUBS 0.007316f
C214 B.n161 VSUBS 0.007316f
C215 B.n162 VSUBS 0.007316f
C216 B.n163 VSUBS 0.007316f
C217 B.n164 VSUBS 0.007316f
C218 B.n165 VSUBS 0.007316f
C219 B.n166 VSUBS 0.007316f
C220 B.n167 VSUBS 0.007316f
C221 B.n168 VSUBS 0.007316f
C222 B.n169 VSUBS 0.007316f
C223 B.n170 VSUBS 0.007316f
C224 B.n171 VSUBS 0.007316f
C225 B.n172 VSUBS 0.007316f
C226 B.n173 VSUBS 0.007316f
C227 B.n174 VSUBS 0.007316f
C228 B.n175 VSUBS 0.007316f
C229 B.n176 VSUBS 0.007316f
C230 B.n177 VSUBS 0.007316f
C231 B.n178 VSUBS 0.007316f
C232 B.n179 VSUBS 0.007316f
C233 B.n180 VSUBS 0.007316f
C234 B.n181 VSUBS 0.007316f
C235 B.n182 VSUBS 0.007316f
C236 B.n183 VSUBS 0.007316f
C237 B.n184 VSUBS 0.007316f
C238 B.n185 VSUBS 0.007316f
C239 B.n186 VSUBS 0.007316f
C240 B.n187 VSUBS 0.007316f
C241 B.n188 VSUBS 0.007316f
C242 B.n189 VSUBS 0.007316f
C243 B.n190 VSUBS 0.007316f
C244 B.n191 VSUBS 0.007316f
C245 B.n192 VSUBS 0.007316f
C246 B.n193 VSUBS 0.007316f
C247 B.n194 VSUBS 0.007316f
C248 B.n195 VSUBS 0.007316f
C249 B.n196 VSUBS 0.007316f
C250 B.n197 VSUBS 0.007316f
C251 B.n198 VSUBS 0.007316f
C252 B.n199 VSUBS 0.007316f
C253 B.n200 VSUBS 0.007316f
C254 B.n201 VSUBS 0.007316f
C255 B.n202 VSUBS 0.007316f
C256 B.n203 VSUBS 0.007316f
C257 B.n204 VSUBS 0.016664f
C258 B.n205 VSUBS 0.017116f
C259 B.n206 VSUBS 0.017116f
C260 B.n207 VSUBS 0.007316f
C261 B.n208 VSUBS 0.007316f
C262 B.n209 VSUBS 0.007316f
C263 B.n210 VSUBS 0.007316f
C264 B.n211 VSUBS 0.007316f
C265 B.n212 VSUBS 0.007316f
C266 B.n213 VSUBS 0.007316f
C267 B.n214 VSUBS 0.007316f
C268 B.n215 VSUBS 0.007316f
C269 B.n216 VSUBS 0.007316f
C270 B.n217 VSUBS 0.007316f
C271 B.n218 VSUBS 0.007316f
C272 B.n219 VSUBS 0.007316f
C273 B.n220 VSUBS 0.007316f
C274 B.n221 VSUBS 0.007316f
C275 B.n222 VSUBS 0.007316f
C276 B.n223 VSUBS 0.007316f
C277 B.n224 VSUBS 0.007316f
C278 B.n225 VSUBS 0.007316f
C279 B.n226 VSUBS 0.007316f
C280 B.n227 VSUBS 0.007316f
C281 B.n228 VSUBS 0.007316f
C282 B.n229 VSUBS 0.007316f
C283 B.n230 VSUBS 0.007316f
C284 B.n231 VSUBS 0.007316f
C285 B.n232 VSUBS 0.007316f
C286 B.n233 VSUBS 0.007316f
C287 B.n234 VSUBS 0.007316f
C288 B.n235 VSUBS 0.007316f
C289 B.n236 VSUBS 0.007316f
C290 B.n237 VSUBS 0.007316f
C291 B.n238 VSUBS 0.007316f
C292 B.n239 VSUBS 0.007316f
C293 B.n240 VSUBS 0.007316f
C294 B.n241 VSUBS 0.007316f
C295 B.n242 VSUBS 0.007316f
C296 B.n243 VSUBS 0.007316f
C297 B.n244 VSUBS 0.007316f
C298 B.n245 VSUBS 0.007316f
C299 B.n246 VSUBS 0.007316f
C300 B.n247 VSUBS 0.007316f
C301 B.n248 VSUBS 0.007316f
C302 B.n249 VSUBS 0.007316f
C303 B.n250 VSUBS 0.007316f
C304 B.n251 VSUBS 0.007316f
C305 B.n252 VSUBS 0.005056f
C306 B.n253 VSUBS 0.016949f
C307 B.n254 VSUBS 0.005917f
C308 B.n255 VSUBS 0.007316f
C309 B.n256 VSUBS 0.007316f
C310 B.n257 VSUBS 0.007316f
C311 B.n258 VSUBS 0.007316f
C312 B.n259 VSUBS 0.007316f
C313 B.n260 VSUBS 0.007316f
C314 B.n261 VSUBS 0.007316f
C315 B.n262 VSUBS 0.007316f
C316 B.n263 VSUBS 0.007316f
C317 B.n264 VSUBS 0.007316f
C318 B.n265 VSUBS 0.007316f
C319 B.n266 VSUBS 0.005917f
C320 B.n267 VSUBS 0.007316f
C321 B.n268 VSUBS 0.007316f
C322 B.n269 VSUBS 0.005056f
C323 B.n270 VSUBS 0.007316f
C324 B.n271 VSUBS 0.007316f
C325 B.n272 VSUBS 0.007316f
C326 B.n273 VSUBS 0.007316f
C327 B.n274 VSUBS 0.007316f
C328 B.n275 VSUBS 0.007316f
C329 B.n276 VSUBS 0.007316f
C330 B.n277 VSUBS 0.007316f
C331 B.n278 VSUBS 0.007316f
C332 B.n279 VSUBS 0.007316f
C333 B.n280 VSUBS 0.007316f
C334 B.n281 VSUBS 0.007316f
C335 B.n282 VSUBS 0.007316f
C336 B.n283 VSUBS 0.007316f
C337 B.n284 VSUBS 0.007316f
C338 B.n285 VSUBS 0.007316f
C339 B.n286 VSUBS 0.007316f
C340 B.n287 VSUBS 0.007316f
C341 B.n288 VSUBS 0.007316f
C342 B.n289 VSUBS 0.007316f
C343 B.n290 VSUBS 0.007316f
C344 B.n291 VSUBS 0.007316f
C345 B.n292 VSUBS 0.007316f
C346 B.n293 VSUBS 0.007316f
C347 B.n294 VSUBS 0.007316f
C348 B.n295 VSUBS 0.007316f
C349 B.n296 VSUBS 0.007316f
C350 B.n297 VSUBS 0.007316f
C351 B.n298 VSUBS 0.007316f
C352 B.n299 VSUBS 0.007316f
C353 B.n300 VSUBS 0.007316f
C354 B.n301 VSUBS 0.007316f
C355 B.n302 VSUBS 0.007316f
C356 B.n303 VSUBS 0.007316f
C357 B.n304 VSUBS 0.007316f
C358 B.n305 VSUBS 0.007316f
C359 B.n306 VSUBS 0.007316f
C360 B.n307 VSUBS 0.007316f
C361 B.n308 VSUBS 0.007316f
C362 B.n309 VSUBS 0.007316f
C363 B.n310 VSUBS 0.007316f
C364 B.n311 VSUBS 0.007316f
C365 B.n312 VSUBS 0.007316f
C366 B.n313 VSUBS 0.007316f
C367 B.n314 VSUBS 0.007316f
C368 B.n315 VSUBS 0.017116f
C369 B.n316 VSUBS 0.016664f
C370 B.n317 VSUBS 0.016664f
C371 B.n318 VSUBS 0.007316f
C372 B.n319 VSUBS 0.007316f
C373 B.n320 VSUBS 0.007316f
C374 B.n321 VSUBS 0.007316f
C375 B.n322 VSUBS 0.007316f
C376 B.n323 VSUBS 0.007316f
C377 B.n324 VSUBS 0.007316f
C378 B.n325 VSUBS 0.007316f
C379 B.n326 VSUBS 0.007316f
C380 B.n327 VSUBS 0.007316f
C381 B.n328 VSUBS 0.007316f
C382 B.n329 VSUBS 0.007316f
C383 B.n330 VSUBS 0.007316f
C384 B.n331 VSUBS 0.007316f
C385 B.n332 VSUBS 0.007316f
C386 B.n333 VSUBS 0.007316f
C387 B.n334 VSUBS 0.007316f
C388 B.n335 VSUBS 0.007316f
C389 B.n336 VSUBS 0.007316f
C390 B.n337 VSUBS 0.007316f
C391 B.n338 VSUBS 0.007316f
C392 B.n339 VSUBS 0.007316f
C393 B.n340 VSUBS 0.007316f
C394 B.n341 VSUBS 0.007316f
C395 B.n342 VSUBS 0.007316f
C396 B.n343 VSUBS 0.007316f
C397 B.n344 VSUBS 0.007316f
C398 B.n345 VSUBS 0.007316f
C399 B.n346 VSUBS 0.007316f
C400 B.n347 VSUBS 0.007316f
C401 B.n348 VSUBS 0.007316f
C402 B.n349 VSUBS 0.007316f
C403 B.n350 VSUBS 0.007316f
C404 B.n351 VSUBS 0.007316f
C405 B.n352 VSUBS 0.007316f
C406 B.n353 VSUBS 0.007316f
C407 B.n354 VSUBS 0.007316f
C408 B.n355 VSUBS 0.007316f
C409 B.n356 VSUBS 0.007316f
C410 B.n357 VSUBS 0.007316f
C411 B.n358 VSUBS 0.007316f
C412 B.n359 VSUBS 0.007316f
C413 B.n360 VSUBS 0.007316f
C414 B.n361 VSUBS 0.007316f
C415 B.n362 VSUBS 0.007316f
C416 B.n363 VSUBS 0.007316f
C417 B.n364 VSUBS 0.007316f
C418 B.n365 VSUBS 0.007316f
C419 B.n366 VSUBS 0.007316f
C420 B.n367 VSUBS 0.007316f
C421 B.n368 VSUBS 0.007316f
C422 B.n369 VSUBS 0.007316f
C423 B.n370 VSUBS 0.007316f
C424 B.n371 VSUBS 0.007316f
C425 B.n372 VSUBS 0.007316f
C426 B.n373 VSUBS 0.007316f
C427 B.n374 VSUBS 0.007316f
C428 B.n375 VSUBS 0.007316f
C429 B.n376 VSUBS 0.007316f
C430 B.n377 VSUBS 0.007316f
C431 B.n378 VSUBS 0.007316f
C432 B.n379 VSUBS 0.007316f
C433 B.n380 VSUBS 0.007316f
C434 B.n381 VSUBS 0.007316f
C435 B.n382 VSUBS 0.007316f
C436 B.n383 VSUBS 0.007316f
C437 B.n384 VSUBS 0.007316f
C438 B.n385 VSUBS 0.007316f
C439 B.n386 VSUBS 0.007316f
C440 B.n387 VSUBS 0.007316f
C441 B.n388 VSUBS 0.007316f
C442 B.n389 VSUBS 0.007316f
C443 B.n390 VSUBS 0.007316f
C444 B.n391 VSUBS 0.007316f
C445 B.n392 VSUBS 0.007316f
C446 B.n393 VSUBS 0.007316f
C447 B.n394 VSUBS 0.007316f
C448 B.n395 VSUBS 0.007316f
C449 B.n396 VSUBS 0.007316f
C450 B.n397 VSUBS 0.007316f
C451 B.n398 VSUBS 0.007316f
C452 B.n399 VSUBS 0.007316f
C453 B.n400 VSUBS 0.007316f
C454 B.n401 VSUBS 0.007316f
C455 B.n402 VSUBS 0.007316f
C456 B.n403 VSUBS 0.007316f
C457 B.n404 VSUBS 0.007316f
C458 B.n405 VSUBS 0.007316f
C459 B.n406 VSUBS 0.007316f
C460 B.n407 VSUBS 0.007316f
C461 B.n408 VSUBS 0.007316f
C462 B.n409 VSUBS 0.007316f
C463 B.n410 VSUBS 0.007316f
C464 B.n411 VSUBS 0.007316f
C465 B.n412 VSUBS 0.007316f
C466 B.n413 VSUBS 0.007316f
C467 B.n414 VSUBS 0.007316f
C468 B.n415 VSUBS 0.007316f
C469 B.n416 VSUBS 0.007316f
C470 B.n417 VSUBS 0.007316f
C471 B.n418 VSUBS 0.007316f
C472 B.n419 VSUBS 0.007316f
C473 B.n420 VSUBS 0.007316f
C474 B.n421 VSUBS 0.017547f
C475 B.n422 VSUBS 0.016664f
C476 B.n423 VSUBS 0.017116f
C477 B.n424 VSUBS 0.007316f
C478 B.n425 VSUBS 0.007316f
C479 B.n426 VSUBS 0.007316f
C480 B.n427 VSUBS 0.007316f
C481 B.n428 VSUBS 0.007316f
C482 B.n429 VSUBS 0.007316f
C483 B.n430 VSUBS 0.007316f
C484 B.n431 VSUBS 0.007316f
C485 B.n432 VSUBS 0.007316f
C486 B.n433 VSUBS 0.007316f
C487 B.n434 VSUBS 0.007316f
C488 B.n435 VSUBS 0.007316f
C489 B.n436 VSUBS 0.007316f
C490 B.n437 VSUBS 0.007316f
C491 B.n438 VSUBS 0.007316f
C492 B.n439 VSUBS 0.007316f
C493 B.n440 VSUBS 0.007316f
C494 B.n441 VSUBS 0.007316f
C495 B.n442 VSUBS 0.007316f
C496 B.n443 VSUBS 0.007316f
C497 B.n444 VSUBS 0.007316f
C498 B.n445 VSUBS 0.007316f
C499 B.n446 VSUBS 0.007316f
C500 B.n447 VSUBS 0.007316f
C501 B.n448 VSUBS 0.007316f
C502 B.n449 VSUBS 0.007316f
C503 B.n450 VSUBS 0.007316f
C504 B.n451 VSUBS 0.007316f
C505 B.n452 VSUBS 0.007316f
C506 B.n453 VSUBS 0.007316f
C507 B.n454 VSUBS 0.007316f
C508 B.n455 VSUBS 0.007316f
C509 B.n456 VSUBS 0.007316f
C510 B.n457 VSUBS 0.007316f
C511 B.n458 VSUBS 0.007316f
C512 B.n459 VSUBS 0.007316f
C513 B.n460 VSUBS 0.007316f
C514 B.n461 VSUBS 0.007316f
C515 B.n462 VSUBS 0.007316f
C516 B.n463 VSUBS 0.007316f
C517 B.n464 VSUBS 0.007316f
C518 B.n465 VSUBS 0.007316f
C519 B.n466 VSUBS 0.007316f
C520 B.n467 VSUBS 0.007316f
C521 B.n468 VSUBS 0.007316f
C522 B.n469 VSUBS 0.005056f
C523 B.n470 VSUBS 0.007316f
C524 B.n471 VSUBS 0.007316f
C525 B.n472 VSUBS 0.005917f
C526 B.n473 VSUBS 0.007316f
C527 B.n474 VSUBS 0.007316f
C528 B.n475 VSUBS 0.007316f
C529 B.n476 VSUBS 0.007316f
C530 B.n477 VSUBS 0.007316f
C531 B.n478 VSUBS 0.007316f
C532 B.n479 VSUBS 0.007316f
C533 B.n480 VSUBS 0.007316f
C534 B.n481 VSUBS 0.007316f
C535 B.n482 VSUBS 0.007316f
C536 B.n483 VSUBS 0.007316f
C537 B.n484 VSUBS 0.005917f
C538 B.n485 VSUBS 0.016949f
C539 B.n486 VSUBS 0.005056f
C540 B.n487 VSUBS 0.007316f
C541 B.n488 VSUBS 0.007316f
C542 B.n489 VSUBS 0.007316f
C543 B.n490 VSUBS 0.007316f
C544 B.n491 VSUBS 0.007316f
C545 B.n492 VSUBS 0.007316f
C546 B.n493 VSUBS 0.007316f
C547 B.n494 VSUBS 0.007316f
C548 B.n495 VSUBS 0.007316f
C549 B.n496 VSUBS 0.007316f
C550 B.n497 VSUBS 0.007316f
C551 B.n498 VSUBS 0.007316f
C552 B.n499 VSUBS 0.007316f
C553 B.n500 VSUBS 0.007316f
C554 B.n501 VSUBS 0.007316f
C555 B.n502 VSUBS 0.007316f
C556 B.n503 VSUBS 0.007316f
C557 B.n504 VSUBS 0.007316f
C558 B.n505 VSUBS 0.007316f
C559 B.n506 VSUBS 0.007316f
C560 B.n507 VSUBS 0.007316f
C561 B.n508 VSUBS 0.007316f
C562 B.n509 VSUBS 0.007316f
C563 B.n510 VSUBS 0.007316f
C564 B.n511 VSUBS 0.007316f
C565 B.n512 VSUBS 0.007316f
C566 B.n513 VSUBS 0.007316f
C567 B.n514 VSUBS 0.007316f
C568 B.n515 VSUBS 0.007316f
C569 B.n516 VSUBS 0.007316f
C570 B.n517 VSUBS 0.007316f
C571 B.n518 VSUBS 0.007316f
C572 B.n519 VSUBS 0.007316f
C573 B.n520 VSUBS 0.007316f
C574 B.n521 VSUBS 0.007316f
C575 B.n522 VSUBS 0.007316f
C576 B.n523 VSUBS 0.007316f
C577 B.n524 VSUBS 0.007316f
C578 B.n525 VSUBS 0.007316f
C579 B.n526 VSUBS 0.007316f
C580 B.n527 VSUBS 0.007316f
C581 B.n528 VSUBS 0.007316f
C582 B.n529 VSUBS 0.007316f
C583 B.n530 VSUBS 0.007316f
C584 B.n531 VSUBS 0.007316f
C585 B.n532 VSUBS 0.017116f
C586 B.n533 VSUBS 0.017116f
C587 B.n534 VSUBS 0.016664f
C588 B.n535 VSUBS 0.007316f
C589 B.n536 VSUBS 0.007316f
C590 B.n537 VSUBS 0.007316f
C591 B.n538 VSUBS 0.007316f
C592 B.n539 VSUBS 0.007316f
C593 B.n540 VSUBS 0.007316f
C594 B.n541 VSUBS 0.007316f
C595 B.n542 VSUBS 0.007316f
C596 B.n543 VSUBS 0.007316f
C597 B.n544 VSUBS 0.007316f
C598 B.n545 VSUBS 0.007316f
C599 B.n546 VSUBS 0.007316f
C600 B.n547 VSUBS 0.007316f
C601 B.n548 VSUBS 0.007316f
C602 B.n549 VSUBS 0.007316f
C603 B.n550 VSUBS 0.007316f
C604 B.n551 VSUBS 0.007316f
C605 B.n552 VSUBS 0.007316f
C606 B.n553 VSUBS 0.007316f
C607 B.n554 VSUBS 0.007316f
C608 B.n555 VSUBS 0.007316f
C609 B.n556 VSUBS 0.007316f
C610 B.n557 VSUBS 0.007316f
C611 B.n558 VSUBS 0.007316f
C612 B.n559 VSUBS 0.007316f
C613 B.n560 VSUBS 0.007316f
C614 B.n561 VSUBS 0.007316f
C615 B.n562 VSUBS 0.007316f
C616 B.n563 VSUBS 0.007316f
C617 B.n564 VSUBS 0.007316f
C618 B.n565 VSUBS 0.007316f
C619 B.n566 VSUBS 0.007316f
C620 B.n567 VSUBS 0.007316f
C621 B.n568 VSUBS 0.007316f
C622 B.n569 VSUBS 0.007316f
C623 B.n570 VSUBS 0.007316f
C624 B.n571 VSUBS 0.007316f
C625 B.n572 VSUBS 0.007316f
C626 B.n573 VSUBS 0.007316f
C627 B.n574 VSUBS 0.007316f
C628 B.n575 VSUBS 0.007316f
C629 B.n576 VSUBS 0.007316f
C630 B.n577 VSUBS 0.007316f
C631 B.n578 VSUBS 0.007316f
C632 B.n579 VSUBS 0.007316f
C633 B.n580 VSUBS 0.007316f
C634 B.n581 VSUBS 0.007316f
C635 B.n582 VSUBS 0.007316f
C636 B.n583 VSUBS 0.007316f
C637 B.n584 VSUBS 0.007316f
C638 B.n585 VSUBS 0.007316f
C639 B.n586 VSUBS 0.007316f
C640 B.n587 VSUBS 0.016565f
C641 VDD1.t1 VSUBS 0.187782f
C642 VDD1.t3 VSUBS 0.187782f
C643 VDD1.n0 VSUBS 1.38594f
C644 VDD1.t0 VSUBS 0.187782f
C645 VDD1.t2 VSUBS 0.187782f
C646 VDD1.n1 VSUBS 1.96195f
C647 VTAIL.n0 VSUBS 0.027001f
C648 VTAIL.n1 VSUBS 0.025154f
C649 VTAIL.n2 VSUBS 0.013517f
C650 VTAIL.n3 VSUBS 0.031948f
C651 VTAIL.n4 VSUBS 0.014312f
C652 VTAIL.n5 VSUBS 0.025154f
C653 VTAIL.n6 VSUBS 0.013517f
C654 VTAIL.n7 VSUBS 0.031948f
C655 VTAIL.n8 VSUBS 0.014312f
C656 VTAIL.n9 VSUBS 0.025154f
C657 VTAIL.n10 VSUBS 0.013517f
C658 VTAIL.n11 VSUBS 0.031948f
C659 VTAIL.n12 VSUBS 0.014312f
C660 VTAIL.n13 VSUBS 0.160291f
C661 VTAIL.t2 VSUBS 0.068636f
C662 VTAIL.n14 VSUBS 0.023961f
C663 VTAIL.n15 VSUBS 0.024033f
C664 VTAIL.n16 VSUBS 0.013517f
C665 VTAIL.n17 VSUBS 0.868745f
C666 VTAIL.n18 VSUBS 0.025154f
C667 VTAIL.n19 VSUBS 0.013517f
C668 VTAIL.n20 VSUBS 0.014312f
C669 VTAIL.n21 VSUBS 0.031948f
C670 VTAIL.n22 VSUBS 0.031948f
C671 VTAIL.n23 VSUBS 0.014312f
C672 VTAIL.n24 VSUBS 0.013517f
C673 VTAIL.n25 VSUBS 0.025154f
C674 VTAIL.n26 VSUBS 0.025154f
C675 VTAIL.n27 VSUBS 0.013517f
C676 VTAIL.n28 VSUBS 0.014312f
C677 VTAIL.n29 VSUBS 0.031948f
C678 VTAIL.n30 VSUBS 0.031948f
C679 VTAIL.n31 VSUBS 0.031948f
C680 VTAIL.n32 VSUBS 0.014312f
C681 VTAIL.n33 VSUBS 0.013517f
C682 VTAIL.n34 VSUBS 0.025154f
C683 VTAIL.n35 VSUBS 0.025154f
C684 VTAIL.n36 VSUBS 0.013517f
C685 VTAIL.n37 VSUBS 0.013914f
C686 VTAIL.n38 VSUBS 0.013914f
C687 VTAIL.n39 VSUBS 0.031948f
C688 VTAIL.n40 VSUBS 0.07517f
C689 VTAIL.n41 VSUBS 0.014312f
C690 VTAIL.n42 VSUBS 0.013517f
C691 VTAIL.n43 VSUBS 0.063297f
C692 VTAIL.n44 VSUBS 0.037858f
C693 VTAIL.n45 VSUBS 0.173052f
C694 VTAIL.n46 VSUBS 0.027001f
C695 VTAIL.n47 VSUBS 0.025154f
C696 VTAIL.n48 VSUBS 0.013517f
C697 VTAIL.n49 VSUBS 0.031948f
C698 VTAIL.n50 VSUBS 0.014312f
C699 VTAIL.n51 VSUBS 0.025154f
C700 VTAIL.n52 VSUBS 0.013517f
C701 VTAIL.n53 VSUBS 0.031948f
C702 VTAIL.n54 VSUBS 0.014312f
C703 VTAIL.n55 VSUBS 0.025154f
C704 VTAIL.n56 VSUBS 0.013517f
C705 VTAIL.n57 VSUBS 0.031948f
C706 VTAIL.n58 VSUBS 0.014312f
C707 VTAIL.n59 VSUBS 0.160291f
C708 VTAIL.t7 VSUBS 0.068636f
C709 VTAIL.n60 VSUBS 0.023961f
C710 VTAIL.n61 VSUBS 0.024033f
C711 VTAIL.n62 VSUBS 0.013517f
C712 VTAIL.n63 VSUBS 0.868745f
C713 VTAIL.n64 VSUBS 0.025154f
C714 VTAIL.n65 VSUBS 0.013517f
C715 VTAIL.n66 VSUBS 0.014312f
C716 VTAIL.n67 VSUBS 0.031948f
C717 VTAIL.n68 VSUBS 0.031948f
C718 VTAIL.n69 VSUBS 0.014312f
C719 VTAIL.n70 VSUBS 0.013517f
C720 VTAIL.n71 VSUBS 0.025154f
C721 VTAIL.n72 VSUBS 0.025154f
C722 VTAIL.n73 VSUBS 0.013517f
C723 VTAIL.n74 VSUBS 0.014312f
C724 VTAIL.n75 VSUBS 0.031948f
C725 VTAIL.n76 VSUBS 0.031948f
C726 VTAIL.n77 VSUBS 0.031948f
C727 VTAIL.n78 VSUBS 0.014312f
C728 VTAIL.n79 VSUBS 0.013517f
C729 VTAIL.n80 VSUBS 0.025154f
C730 VTAIL.n81 VSUBS 0.025154f
C731 VTAIL.n82 VSUBS 0.013517f
C732 VTAIL.n83 VSUBS 0.013914f
C733 VTAIL.n84 VSUBS 0.013914f
C734 VTAIL.n85 VSUBS 0.031948f
C735 VTAIL.n86 VSUBS 0.07517f
C736 VTAIL.n87 VSUBS 0.014312f
C737 VTAIL.n88 VSUBS 0.013517f
C738 VTAIL.n89 VSUBS 0.063297f
C739 VTAIL.n90 VSUBS 0.037858f
C740 VTAIL.n91 VSUBS 0.274192f
C741 VTAIL.n92 VSUBS 0.027001f
C742 VTAIL.n93 VSUBS 0.025154f
C743 VTAIL.n94 VSUBS 0.013517f
C744 VTAIL.n95 VSUBS 0.031948f
C745 VTAIL.n96 VSUBS 0.014312f
C746 VTAIL.n97 VSUBS 0.025154f
C747 VTAIL.n98 VSUBS 0.013517f
C748 VTAIL.n99 VSUBS 0.031948f
C749 VTAIL.n100 VSUBS 0.014312f
C750 VTAIL.n101 VSUBS 0.025154f
C751 VTAIL.n102 VSUBS 0.013517f
C752 VTAIL.n103 VSUBS 0.031948f
C753 VTAIL.n104 VSUBS 0.014312f
C754 VTAIL.n105 VSUBS 0.160291f
C755 VTAIL.t4 VSUBS 0.068636f
C756 VTAIL.n106 VSUBS 0.023961f
C757 VTAIL.n107 VSUBS 0.024033f
C758 VTAIL.n108 VSUBS 0.013517f
C759 VTAIL.n109 VSUBS 0.868745f
C760 VTAIL.n110 VSUBS 0.025154f
C761 VTAIL.n111 VSUBS 0.013517f
C762 VTAIL.n112 VSUBS 0.014312f
C763 VTAIL.n113 VSUBS 0.031948f
C764 VTAIL.n114 VSUBS 0.031948f
C765 VTAIL.n115 VSUBS 0.014312f
C766 VTAIL.n116 VSUBS 0.013517f
C767 VTAIL.n117 VSUBS 0.025154f
C768 VTAIL.n118 VSUBS 0.025154f
C769 VTAIL.n119 VSUBS 0.013517f
C770 VTAIL.n120 VSUBS 0.014312f
C771 VTAIL.n121 VSUBS 0.031948f
C772 VTAIL.n122 VSUBS 0.031948f
C773 VTAIL.n123 VSUBS 0.031948f
C774 VTAIL.n124 VSUBS 0.014312f
C775 VTAIL.n125 VSUBS 0.013517f
C776 VTAIL.n126 VSUBS 0.025154f
C777 VTAIL.n127 VSUBS 0.025154f
C778 VTAIL.n128 VSUBS 0.013517f
C779 VTAIL.n129 VSUBS 0.013914f
C780 VTAIL.n130 VSUBS 0.013914f
C781 VTAIL.n131 VSUBS 0.031948f
C782 VTAIL.n132 VSUBS 0.07517f
C783 VTAIL.n133 VSUBS 0.014312f
C784 VTAIL.n134 VSUBS 0.013517f
C785 VTAIL.n135 VSUBS 0.063297f
C786 VTAIL.n136 VSUBS 0.037858f
C787 VTAIL.n137 VSUBS 1.39531f
C788 VTAIL.n138 VSUBS 0.027001f
C789 VTAIL.n139 VSUBS 0.025154f
C790 VTAIL.n140 VSUBS 0.013517f
C791 VTAIL.n141 VSUBS 0.031948f
C792 VTAIL.n142 VSUBS 0.014312f
C793 VTAIL.n143 VSUBS 0.025154f
C794 VTAIL.n144 VSUBS 0.013517f
C795 VTAIL.n145 VSUBS 0.031948f
C796 VTAIL.n146 VSUBS 0.031948f
C797 VTAIL.n147 VSUBS 0.014312f
C798 VTAIL.n148 VSUBS 0.025154f
C799 VTAIL.n149 VSUBS 0.013517f
C800 VTAIL.n150 VSUBS 0.031948f
C801 VTAIL.n151 VSUBS 0.014312f
C802 VTAIL.n152 VSUBS 0.160291f
C803 VTAIL.t1 VSUBS 0.068636f
C804 VTAIL.n153 VSUBS 0.023961f
C805 VTAIL.n154 VSUBS 0.024033f
C806 VTAIL.n155 VSUBS 0.013517f
C807 VTAIL.n156 VSUBS 0.868745f
C808 VTAIL.n157 VSUBS 0.025154f
C809 VTAIL.n158 VSUBS 0.013517f
C810 VTAIL.n159 VSUBS 0.014312f
C811 VTAIL.n160 VSUBS 0.031948f
C812 VTAIL.n161 VSUBS 0.031948f
C813 VTAIL.n162 VSUBS 0.014312f
C814 VTAIL.n163 VSUBS 0.013517f
C815 VTAIL.n164 VSUBS 0.025154f
C816 VTAIL.n165 VSUBS 0.025154f
C817 VTAIL.n166 VSUBS 0.013517f
C818 VTAIL.n167 VSUBS 0.014312f
C819 VTAIL.n168 VSUBS 0.031948f
C820 VTAIL.n169 VSUBS 0.031948f
C821 VTAIL.n170 VSUBS 0.014312f
C822 VTAIL.n171 VSUBS 0.013517f
C823 VTAIL.n172 VSUBS 0.025154f
C824 VTAIL.n173 VSUBS 0.025154f
C825 VTAIL.n174 VSUBS 0.013517f
C826 VTAIL.n175 VSUBS 0.013914f
C827 VTAIL.n176 VSUBS 0.013914f
C828 VTAIL.n177 VSUBS 0.031948f
C829 VTAIL.n178 VSUBS 0.07517f
C830 VTAIL.n179 VSUBS 0.014312f
C831 VTAIL.n180 VSUBS 0.013517f
C832 VTAIL.n181 VSUBS 0.063297f
C833 VTAIL.n182 VSUBS 0.037858f
C834 VTAIL.n183 VSUBS 1.39531f
C835 VTAIL.n184 VSUBS 0.027001f
C836 VTAIL.n185 VSUBS 0.025154f
C837 VTAIL.n186 VSUBS 0.013517f
C838 VTAIL.n187 VSUBS 0.031948f
C839 VTAIL.n188 VSUBS 0.014312f
C840 VTAIL.n189 VSUBS 0.025154f
C841 VTAIL.n190 VSUBS 0.013517f
C842 VTAIL.n191 VSUBS 0.031948f
C843 VTAIL.n192 VSUBS 0.031948f
C844 VTAIL.n193 VSUBS 0.014312f
C845 VTAIL.n194 VSUBS 0.025154f
C846 VTAIL.n195 VSUBS 0.013517f
C847 VTAIL.n196 VSUBS 0.031948f
C848 VTAIL.n197 VSUBS 0.014312f
C849 VTAIL.n198 VSUBS 0.160291f
C850 VTAIL.t0 VSUBS 0.068636f
C851 VTAIL.n199 VSUBS 0.023961f
C852 VTAIL.n200 VSUBS 0.024033f
C853 VTAIL.n201 VSUBS 0.013517f
C854 VTAIL.n202 VSUBS 0.868745f
C855 VTAIL.n203 VSUBS 0.025154f
C856 VTAIL.n204 VSUBS 0.013517f
C857 VTAIL.n205 VSUBS 0.014312f
C858 VTAIL.n206 VSUBS 0.031948f
C859 VTAIL.n207 VSUBS 0.031948f
C860 VTAIL.n208 VSUBS 0.014312f
C861 VTAIL.n209 VSUBS 0.013517f
C862 VTAIL.n210 VSUBS 0.025154f
C863 VTAIL.n211 VSUBS 0.025154f
C864 VTAIL.n212 VSUBS 0.013517f
C865 VTAIL.n213 VSUBS 0.014312f
C866 VTAIL.n214 VSUBS 0.031948f
C867 VTAIL.n215 VSUBS 0.031948f
C868 VTAIL.n216 VSUBS 0.014312f
C869 VTAIL.n217 VSUBS 0.013517f
C870 VTAIL.n218 VSUBS 0.025154f
C871 VTAIL.n219 VSUBS 0.025154f
C872 VTAIL.n220 VSUBS 0.013517f
C873 VTAIL.n221 VSUBS 0.013914f
C874 VTAIL.n222 VSUBS 0.013914f
C875 VTAIL.n223 VSUBS 0.031948f
C876 VTAIL.n224 VSUBS 0.07517f
C877 VTAIL.n225 VSUBS 0.014312f
C878 VTAIL.n226 VSUBS 0.013517f
C879 VTAIL.n227 VSUBS 0.063297f
C880 VTAIL.n228 VSUBS 0.037858f
C881 VTAIL.n229 VSUBS 0.274192f
C882 VTAIL.n230 VSUBS 0.027001f
C883 VTAIL.n231 VSUBS 0.025154f
C884 VTAIL.n232 VSUBS 0.013517f
C885 VTAIL.n233 VSUBS 0.031948f
C886 VTAIL.n234 VSUBS 0.014312f
C887 VTAIL.n235 VSUBS 0.025154f
C888 VTAIL.n236 VSUBS 0.013517f
C889 VTAIL.n237 VSUBS 0.031948f
C890 VTAIL.n238 VSUBS 0.031948f
C891 VTAIL.n239 VSUBS 0.014312f
C892 VTAIL.n240 VSUBS 0.025154f
C893 VTAIL.n241 VSUBS 0.013517f
C894 VTAIL.n242 VSUBS 0.031948f
C895 VTAIL.n243 VSUBS 0.014312f
C896 VTAIL.n244 VSUBS 0.160291f
C897 VTAIL.t5 VSUBS 0.068636f
C898 VTAIL.n245 VSUBS 0.023961f
C899 VTAIL.n246 VSUBS 0.024033f
C900 VTAIL.n247 VSUBS 0.013517f
C901 VTAIL.n248 VSUBS 0.868745f
C902 VTAIL.n249 VSUBS 0.025154f
C903 VTAIL.n250 VSUBS 0.013517f
C904 VTAIL.n251 VSUBS 0.014312f
C905 VTAIL.n252 VSUBS 0.031948f
C906 VTAIL.n253 VSUBS 0.031948f
C907 VTAIL.n254 VSUBS 0.014312f
C908 VTAIL.n255 VSUBS 0.013517f
C909 VTAIL.n256 VSUBS 0.025154f
C910 VTAIL.n257 VSUBS 0.025154f
C911 VTAIL.n258 VSUBS 0.013517f
C912 VTAIL.n259 VSUBS 0.014312f
C913 VTAIL.n260 VSUBS 0.031948f
C914 VTAIL.n261 VSUBS 0.031948f
C915 VTAIL.n262 VSUBS 0.014312f
C916 VTAIL.n263 VSUBS 0.013517f
C917 VTAIL.n264 VSUBS 0.025154f
C918 VTAIL.n265 VSUBS 0.025154f
C919 VTAIL.n266 VSUBS 0.013517f
C920 VTAIL.n267 VSUBS 0.013914f
C921 VTAIL.n268 VSUBS 0.013914f
C922 VTAIL.n269 VSUBS 0.031948f
C923 VTAIL.n270 VSUBS 0.07517f
C924 VTAIL.n271 VSUBS 0.014312f
C925 VTAIL.n272 VSUBS 0.013517f
C926 VTAIL.n273 VSUBS 0.063297f
C927 VTAIL.n274 VSUBS 0.037858f
C928 VTAIL.n275 VSUBS 0.274192f
C929 VTAIL.n276 VSUBS 0.027001f
C930 VTAIL.n277 VSUBS 0.025154f
C931 VTAIL.n278 VSUBS 0.013517f
C932 VTAIL.n279 VSUBS 0.031948f
C933 VTAIL.n280 VSUBS 0.014312f
C934 VTAIL.n281 VSUBS 0.025154f
C935 VTAIL.n282 VSUBS 0.013517f
C936 VTAIL.n283 VSUBS 0.031948f
C937 VTAIL.n284 VSUBS 0.031948f
C938 VTAIL.n285 VSUBS 0.014312f
C939 VTAIL.n286 VSUBS 0.025154f
C940 VTAIL.n287 VSUBS 0.013517f
C941 VTAIL.n288 VSUBS 0.031948f
C942 VTAIL.n289 VSUBS 0.014312f
C943 VTAIL.n290 VSUBS 0.160291f
C944 VTAIL.t6 VSUBS 0.068636f
C945 VTAIL.n291 VSUBS 0.023961f
C946 VTAIL.n292 VSUBS 0.024033f
C947 VTAIL.n293 VSUBS 0.013517f
C948 VTAIL.n294 VSUBS 0.868745f
C949 VTAIL.n295 VSUBS 0.025154f
C950 VTAIL.n296 VSUBS 0.013517f
C951 VTAIL.n297 VSUBS 0.014312f
C952 VTAIL.n298 VSUBS 0.031948f
C953 VTAIL.n299 VSUBS 0.031948f
C954 VTAIL.n300 VSUBS 0.014312f
C955 VTAIL.n301 VSUBS 0.013517f
C956 VTAIL.n302 VSUBS 0.025154f
C957 VTAIL.n303 VSUBS 0.025154f
C958 VTAIL.n304 VSUBS 0.013517f
C959 VTAIL.n305 VSUBS 0.014312f
C960 VTAIL.n306 VSUBS 0.031948f
C961 VTAIL.n307 VSUBS 0.031948f
C962 VTAIL.n308 VSUBS 0.014312f
C963 VTAIL.n309 VSUBS 0.013517f
C964 VTAIL.n310 VSUBS 0.025154f
C965 VTAIL.n311 VSUBS 0.025154f
C966 VTAIL.n312 VSUBS 0.013517f
C967 VTAIL.n313 VSUBS 0.013914f
C968 VTAIL.n314 VSUBS 0.013914f
C969 VTAIL.n315 VSUBS 0.031948f
C970 VTAIL.n316 VSUBS 0.07517f
C971 VTAIL.n317 VSUBS 0.014312f
C972 VTAIL.n318 VSUBS 0.013517f
C973 VTAIL.n319 VSUBS 0.063297f
C974 VTAIL.n320 VSUBS 0.037858f
C975 VTAIL.n321 VSUBS 1.39531f
C976 VTAIL.n322 VSUBS 0.027001f
C977 VTAIL.n323 VSUBS 0.025154f
C978 VTAIL.n324 VSUBS 0.013517f
C979 VTAIL.n325 VSUBS 0.031948f
C980 VTAIL.n326 VSUBS 0.014312f
C981 VTAIL.n327 VSUBS 0.025154f
C982 VTAIL.n328 VSUBS 0.013517f
C983 VTAIL.n329 VSUBS 0.031948f
C984 VTAIL.n330 VSUBS 0.014312f
C985 VTAIL.n331 VSUBS 0.025154f
C986 VTAIL.n332 VSUBS 0.013517f
C987 VTAIL.n333 VSUBS 0.031948f
C988 VTAIL.n334 VSUBS 0.014312f
C989 VTAIL.n335 VSUBS 0.160291f
C990 VTAIL.t3 VSUBS 0.068636f
C991 VTAIL.n336 VSUBS 0.023961f
C992 VTAIL.n337 VSUBS 0.024033f
C993 VTAIL.n338 VSUBS 0.013517f
C994 VTAIL.n339 VSUBS 0.868745f
C995 VTAIL.n340 VSUBS 0.025154f
C996 VTAIL.n341 VSUBS 0.013517f
C997 VTAIL.n342 VSUBS 0.014312f
C998 VTAIL.n343 VSUBS 0.031948f
C999 VTAIL.n344 VSUBS 0.031948f
C1000 VTAIL.n345 VSUBS 0.014312f
C1001 VTAIL.n346 VSUBS 0.013517f
C1002 VTAIL.n347 VSUBS 0.025154f
C1003 VTAIL.n348 VSUBS 0.025154f
C1004 VTAIL.n349 VSUBS 0.013517f
C1005 VTAIL.n350 VSUBS 0.014312f
C1006 VTAIL.n351 VSUBS 0.031948f
C1007 VTAIL.n352 VSUBS 0.031948f
C1008 VTAIL.n353 VSUBS 0.031948f
C1009 VTAIL.n354 VSUBS 0.014312f
C1010 VTAIL.n355 VSUBS 0.013517f
C1011 VTAIL.n356 VSUBS 0.025154f
C1012 VTAIL.n357 VSUBS 0.025154f
C1013 VTAIL.n358 VSUBS 0.013517f
C1014 VTAIL.n359 VSUBS 0.013914f
C1015 VTAIL.n360 VSUBS 0.013914f
C1016 VTAIL.n361 VSUBS 0.031948f
C1017 VTAIL.n362 VSUBS 0.07517f
C1018 VTAIL.n363 VSUBS 0.014312f
C1019 VTAIL.n364 VSUBS 0.013517f
C1020 VTAIL.n365 VSUBS 0.063297f
C1021 VTAIL.n366 VSUBS 0.037858f
C1022 VTAIL.n367 VSUBS 1.28473f
C1023 VP.n0 VSUBS 0.048342f
C1024 VP.t1 VSUBS 2.31298f
C1025 VP.n1 VSUBS 0.072875f
C1026 VP.n2 VSUBS 0.036667f
C1027 VP.n3 VSUBS 0.03561f
C1028 VP.t0 VSUBS 2.63491f
C1029 VP.t2 VSUBS 2.6432f
C1030 VP.n4 VSUBS 3.5567f
C1031 VP.t3 VSUBS 2.31298f
C1032 VP.n5 VSUBS 0.945463f
C1033 VP.n6 VSUBS 1.87688f
C1034 VP.n7 VSUBS 0.048342f
C1035 VP.n8 VSUBS 0.036667f
C1036 VP.n9 VSUBS 0.068338f
C1037 VP.n10 VSUBS 0.072875f
C1038 VP.n11 VSUBS 0.029642f
C1039 VP.n12 VSUBS 0.036667f
C1040 VP.n13 VSUBS 0.036667f
C1041 VP.n14 VSUBS 0.036667f
C1042 VP.n15 VSUBS 0.068338f
C1043 VP.n16 VSUBS 0.03561f
C1044 VP.n17 VSUBS 0.945463f
C1045 VP.n18 VSUBS 0.068414f
.ends

