(* blackbox *) module sky130_fd_sc_hvl__a2111o_1(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2111o_2(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2111o_4(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2111oi_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2111oi_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2111oi_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211o_1(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211o_2(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211o_4(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211oi_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211oi_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a211oi_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21bo_1(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21bo_2(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21bo_4(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21boi_1(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21boi_2(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21boi_4(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21o_1(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21o_2(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21o_4(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21oi_1(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21oi_2(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a21oi_4(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221o_1(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221o_2(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221o_4(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221oi_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221oi_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a221oi_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a222o_1(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1,
  input C2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a222o_2(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1,
  input C2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a222oi_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1,
  input C2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a222oi_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1,
  input C2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22o_1(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22o_2(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22o_4(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22oi_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22oi_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a22oi_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2o_1(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2o_2(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2o_4(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2oi_1(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2oi_2(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a2bb2oi_4(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311o_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311o_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311o_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311oi_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311oi_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a311oi_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31o_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31o_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31o_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31oi_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31oi_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a31oi_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32o_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32o_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32o_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32oi_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32oi_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a32oi_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41o_1(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41o_2(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41o_4(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41oi_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41oi_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__a41oi_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2_1(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2_2(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2_4(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2b_1(
  output X,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2b_2(
  output X,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and2b_4(
  output X,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3_1(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3_2(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3_4(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3b_1(
  output X,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3b_2(
  output X,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and3b_4(
  output X,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4_1(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4_2(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4_4(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4b_1(
  output X,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4b_2(
  output X,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4b_4(
  output X,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4bb_1(
  output X,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4bb_2(
  output X,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__and4bb_4(
  output X,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__buf_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__buf_16(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__buf_2(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__buf_4(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__buf_8(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__bufbuf_16(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__bufbuf_8(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__bufinv_16(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__bufinv_8(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkbuf_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkbuf_16(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkbuf_2(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkbuf_4(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkbuf_8(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv3sd1_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv3sd2_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv3sd3_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv5sd1_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv5sd2_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkdlyinv5sd3_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkinv_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkinv_16(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkinv_2(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkinv_4(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__clkinv_8(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__conb_1(
  output HI,
  output LO
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__decap_4(
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__decap_8(
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfbbn_1(
  input SET_B,
  input RESET_B,
  input CLK_N,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfbbn_2(
  input SET_B,
  input RESET_B,
  input CLK_N,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfbbp_1(
  input SET_B,
  input RESET_B,
  input CLK,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrbp_1(
  input RESET_B,
  input CLK,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrbp_2(
  input RESET_B,
  input CLK,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrtn_1(
  input RESET_B,
  input CLK_N,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrtp_1(
  input RESET_B,
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrtp_2(
  input RESET_B,
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfrtp_4(
  input RESET_B,
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfsbp_1(
  input CLK,
  input D,
  output Q,
  output Q_N,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfsbp_2(
  input CLK,
  input D,
  output Q,
  output Q_N,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfstp_1(
  input CLK,
  input D,
  output Q,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfstp_2(
  input CLK,
  input D,
  output Q,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfstp_4(
  input CLK,
  input D,
  output Q,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfxbp_1(
  input CLK,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfxbp_2(
  input CLK,
  input D,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfxtp_1(
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfxtp_2(
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dfxtp_4(
  input CLK,
  input D,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlclkp_1(
  output GCLK,
  input CLK,
  input GATE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlclkp_2(
  output GCLK,
  input CLK,
  input GATE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlclkp_4(
  output GCLK,
  input CLK,
  input GATE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrbn_1(
  input RESET_B,
  input D,
  input GATE_N,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrbn_2(
  input RESET_B,
  input D,
  input GATE_N,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrbp_1(
  input RESET_B,
  input D,
  input GATE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrbp_2(
  input RESET_B,
  input D,
  input GATE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtn_1(
  input RESET_B,
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtn_2(
  input RESET_B,
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtn_4(
  input RESET_B,
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtp_1(
  input RESET_B,
  input D,
  input GATE,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtp_2(
  input RESET_B,
  input D,
  input GATE,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlrtp_4(
  input RESET_B,
  input D,
  input GATE,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxbn_1(
  input D,
  input GATE_N,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxbn_2(
  input D,
  input GATE_N,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxbp_1(
  input D,
  input GATE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxtn_1(
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxtn_2(
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxtn_4(
  input D,
  input GATE_N,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlxtp_1(
  input D,
  input GATE,
  output Q
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlygate4sd1_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlygate4sd2_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlygate4sd3_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlymetal6s2s_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlymetal6s4s_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__dlymetal6s6s_1(
  output X,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ebufn_1(
  output Z,
  input A,
  input TE_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ebufn_2(
  output Z,
  input A,
  input TE_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ebufn_4(
  output Z,
  input A,
  input TE_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ebufn_8(
  output Z,
  input A,
  input TE_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__edfxbp_1(
  output Q,
  output Q_N,
  input CLK,
  input D,
  input DE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__edfxtp_1(
  output Q,
  input CLK,
  input D,
  input DE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvn_1(
  input A,
  input TE_B,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvn_2(
  input A,
  input TE_B,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvn_4(
  input A,
  input TE_B,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvn_8(
  input A,
  input TE_B,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvp_1(
  input A,
  input TE,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvp_2(
  input A,
  input TE,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvp_4(
  input A,
  input TE,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__einvp_8(
  input A,
  input TE,
  output Z
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fa_1(
  output COUT,
  output SUM,
  input A,
  input B,
  input CIN
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fa_2(
  output COUT,
  output SUM,
  input A,
  input B,
  input CIN
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fa_4(
  output COUT,
  output SUM,
  input A,
  input B,
  input CIN
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fah_1(
  output COUT,
  output SUM,
  input A,
  input B,
  input CI
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fah_2(
  output COUT,
  output SUM,
  input A,
  input B,
  input CI
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fah_4(
  output COUT,
  output SUM,
  input A,
  input B,
  input CI
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fahcin_1(
  output COUT,
  output SUM,
  input A,
  input B,
  input CIN
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__fahcon_1(
  output COUT_N,
  output SUM,
  input A,
  input B,
  input CI
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ha_1(
  output COUT,
  output SUM,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ha_2(
  output COUT,
  output SUM,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__ha_4(
  output COUT,
  output SUM,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__inv_1(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__inv_16(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__inv_2(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__inv_4(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__inv_8(
  output Y,
  input A
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__maj3_1(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__maj3_2(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__maj3_4(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2_1(
  output X,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2_2(
  output X,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2_4(
  output X,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2i_1(
  output Y,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2i_2(
  output Y,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux2i_4(
  output Y,
  input A0,
  input A1,
  input S
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux4_1(
  output X,
  input A0,
  input A1,
  input A2,
  input A3,
  input S0,
  input S1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux4_2(
  output X,
  input A0,
  input A1,
  input A2,
  input A3,
  input S0,
  input S1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__mux4_4(
  output X,
  input A0,
  input A1,
  input A2,
  input A3,
  input S0,
  input S1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2_1(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2_2(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2_4(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2_8(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2b_1(
  output Y,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2b_2(
  output Y,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand2b_4(
  output Y,
  input A_N,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3_1(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3_2(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3_4(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3b_1(
  output Y,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3b_2(
  output Y,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand3b_4(
  output Y,
  input A_N,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4_1(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4_2(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4_4(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4b_1(
  output Y,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4b_2(
  output Y,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4b_4(
  output Y,
  input A_N,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4bb_1(
  output Y,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4bb_2(
  output Y,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nand4bb_4(
  output Y,
  input A_N,
  input B_N,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2_1(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2_2(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2_4(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2_8(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2b_1(
  output Y,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2b_2(
  output Y,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor2b_4(
  output Y,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3_1(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3_2(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3_4(
  output Y,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3b_1(
  output Y,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3b_2(
  output Y,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor3b_4(
  output Y,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4_1(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4_2(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4_4(
  output Y,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4b_1(
  output Y,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4b_2(
  output Y,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4b_4(
  output Y,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4bb_1(
  output Y,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4bb_2(
  output Y,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__nor4bb_4(
  output Y,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111a_1(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111a_2(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111a_4(
  output X,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111ai_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111ai_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2111ai_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1,
  input D1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211a_1(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211a_2(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211a_4(
  output X,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211ai_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211ai_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o211ai_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21a_1(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21a_2(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21a_4(
  output X,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ai_1(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ai_2(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ai_4(
  output Y,
  input A1,
  input A2,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ba_1(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ba_2(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21ba_4(
  output X,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21bai_1(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21bai_2(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o21bai_4(
  output Y,
  input A1,
  input A2,
  input B1_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221a_1(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221a_2(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221a_4(
  output X,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221ai_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221ai_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o221ai_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22a_1(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22a_2(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22a_4(
  output X,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22ai_1(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22ai_2(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o22ai_4(
  output Y,
  input A1,
  input A2,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2a_1(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2a_2(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2a_4(
  output X,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2ai_1(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2ai_2(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o2bb2ai_4(
  output Y,
  input A1_N,
  input A2_N,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311a_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311a_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311a_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311ai_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311ai_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o311ai_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input C1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31a_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31a_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31a_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31ai_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31ai_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o31ai_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32a_1(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32a_2(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32a_4(
  output X,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32ai_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32ai_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o32ai_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input B1,
  input B2
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41a_1(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41a_2(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41a_4(
  output X,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41ai_1(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41ai_2(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__o41ai_4(
  output Y,
  input A1,
  input A2,
  input A3,
  input A4,
  input B1
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2_1(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2_2(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2_4(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2b_1(
  output X,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2b_2(
  output X,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or2b_4(
  output X,
  input A,
  input B_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3_1(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3_2(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3_4(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3b_1(
  output X,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3b_2(
  output X,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or3b_4(
  output X,
  input A,
  input B,
  input C_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4_1(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4_2(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4_4(
  output X,
  input A,
  input B,
  input C,
  input D
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4b_1(
  output X,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4b_2(
  output X,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4b_4(
  output X,
  input A,
  input B,
  input C,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4bb_1(
  output X,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4bb_2(
  output X,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__or4bb_4(
  output X,
  input A,
  input B,
  input C_N,
  input D_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfbbn_1(
  input SET_B,
    input RESET_B,
    input CLK_N,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input SET_B,
  input RESET_B,
  input CLK_N,
  input D,
  input SCD,
  input SCE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfbbn_2(
  input SET_B,
    input RESET_B,
    input CLK_N,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input SET_B,
  input RESET_B,
  input CLK_N,
  input D,
  input SCD,
  input SCE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfbbp_1(
  input SET_B,
    input RESET_B,
    input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input SET_B,
  input RESET_B,
  input CLK,
  input D,
  input SCD,
  input SCE,
  output Q,
  output Q_N
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrbp_1(
  input RESET_B,
    input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrbp_2(
  input RESET_B,
    input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrtn_1(
  input RESET_B,
    input CLK_N,
    input D,
    output Q,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK_N,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrtp_1(
  input RESET_B,
    input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrtp_2(
  input RESET_B,
    input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfrtp_4(
  input RESET_B,
    input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input RESET_B,
  input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfsbp_1(
  input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input SET_B,
    input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfsbp_2(
  input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input SET_B,
    input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfstp_1(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input SET_B,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfstp_2(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input SET_B,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfstp_4(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input SET_B,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE,
  input SET_B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfxbp_1(
  input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfxbp_2(
  input CLK,
    input D,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    input CLK,
  input D,
  output Q,
  output Q_N,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfxtp_1(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfxtp_2(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdfxtp_4(
  input CLK,
    input D,
    output Q,
    input SCD,
    input SCE,
    input CLK,
  input D,
  output Q,
  input SCD,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdlclkp_1(
  output GCLK,
  input CLK,
  input GATE,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdlclkp_2(
  output GCLK,
  input CLK,
  input GATE,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sdlclkp_4(
  output GCLK,
  input CLK,
  input GATE,
  input SCE
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sedfxbp_1(
  input CLK,
    input D,
    input DE,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    output Q,
  output Q_N,
  input CLK,
  input D,
  input DE,
  input SCE,
  input SCD
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sedfxbp_2(
  input CLK,
    input D,
    input DE,
    output Q,
    output Q_N,
    input SCD,
    input SCE,
    output Q,
  output Q_N,
  input CLK,
  input D,
  input DE,
  input SCE,
  input SCD
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sedfxtp_1(
  input CLK,
    input D,
    input DE,
    output Q,
    input SCD,
    input SCE,
    output Q,
  input CLK,
  input D,
  input DE,
  input SCE,
  input SCD
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sedfxtp_2(
  input CLK,
    input D,
    input DE,
    output Q,
    input SCD,
    input SCE,
    output Q,
  input CLK,
  input D,
  input DE,
  input SCE,
  input SCD
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__sedfxtp_4(
  input CLK,
    input D,
    input DE,
    output Q,
    input SCD,
    input SCE,
    output Q,
  input CLK,
  input D,
  input DE,
  input SCE,
  input SCD
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor2_1(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor2_2(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor2_4(
  output Y,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor3_1(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor3_2(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xnor3_4(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor2_1(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor2_2(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor2_4(
  output X,
  input A,
  input B
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor3_1(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor3_2(
  output X,
  input A,
  input B,
  input C
);
endmodule
(* blackbox *) module sky130_fd_sc_hvl__xor3_4(
  output X,
  input A,
  input B,
  input C
);
endmodule
