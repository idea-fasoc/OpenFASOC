* NGSPICE file created from diff_pair_sample_1520.ext - technology: sky130A

.subckt diff_pair_sample_1520 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=2.71
X1 VDD2.t9 VN.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=2.71
X2 VTAIL.t3 VP.t0 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X3 VDD1.t8 VP.t1 VTAIL.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=2.71
X4 VTAIL.t11 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X5 VTAIL.t12 VN.t2 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X6 VDD2.t6 VN.t3 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X7 VTAIL.t8 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=2.71
X9 VDD1.t7 VP.t2 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=2.71
X10 VDD1.t6 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=2.71
X11 VDD2.t4 VN.t5 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=2.71
X12 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=2.71
X13 VDD1.t4 VP.t5 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X14 VTAIL.t15 VN.t6 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=2.71
X16 VDD2.t2 VN.t7 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=2.71
X17 VTAIL.t7 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=2.71
X19 VDD1.t2 VP.t7 VTAIL.t19 B.t5 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X20 VTAIL.t5 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X21 VDD2.t1 VN.t8 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=2.71
X22 VDD2.t0 VN.t9 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
X23 VTAIL.t1 VP.t9 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=2.71
R0 B.n830 B.n829 585
R1 B.n831 B.n830 585
R2 B.n278 B.n145 585
R3 B.n277 B.n276 585
R4 B.n275 B.n274 585
R5 B.n273 B.n272 585
R6 B.n271 B.n270 585
R7 B.n269 B.n268 585
R8 B.n267 B.n266 585
R9 B.n265 B.n264 585
R10 B.n263 B.n262 585
R11 B.n261 B.n260 585
R12 B.n259 B.n258 585
R13 B.n257 B.n256 585
R14 B.n255 B.n254 585
R15 B.n253 B.n252 585
R16 B.n251 B.n250 585
R17 B.n249 B.n248 585
R18 B.n247 B.n246 585
R19 B.n245 B.n244 585
R20 B.n243 B.n242 585
R21 B.n241 B.n240 585
R22 B.n239 B.n238 585
R23 B.n237 B.n236 585
R24 B.n235 B.n234 585
R25 B.n233 B.n232 585
R26 B.n231 B.n230 585
R27 B.n229 B.n228 585
R28 B.n227 B.n226 585
R29 B.n224 B.n223 585
R30 B.n222 B.n221 585
R31 B.n220 B.n219 585
R32 B.n218 B.n217 585
R33 B.n216 B.n215 585
R34 B.n214 B.n213 585
R35 B.n212 B.n211 585
R36 B.n210 B.n209 585
R37 B.n208 B.n207 585
R38 B.n206 B.n205 585
R39 B.n204 B.n203 585
R40 B.n202 B.n201 585
R41 B.n200 B.n199 585
R42 B.n198 B.n197 585
R43 B.n196 B.n195 585
R44 B.n194 B.n193 585
R45 B.n192 B.n191 585
R46 B.n190 B.n189 585
R47 B.n188 B.n187 585
R48 B.n186 B.n185 585
R49 B.n184 B.n183 585
R50 B.n182 B.n181 585
R51 B.n180 B.n179 585
R52 B.n178 B.n177 585
R53 B.n176 B.n175 585
R54 B.n174 B.n173 585
R55 B.n172 B.n171 585
R56 B.n170 B.n169 585
R57 B.n168 B.n167 585
R58 B.n166 B.n165 585
R59 B.n164 B.n163 585
R60 B.n162 B.n161 585
R61 B.n160 B.n159 585
R62 B.n158 B.n157 585
R63 B.n156 B.n155 585
R64 B.n154 B.n153 585
R65 B.n152 B.n151 585
R66 B.n828 B.n112 585
R67 B.n832 B.n112 585
R68 B.n827 B.n111 585
R69 B.n833 B.n111 585
R70 B.n826 B.n825 585
R71 B.n825 B.n107 585
R72 B.n824 B.n106 585
R73 B.n839 B.n106 585
R74 B.n823 B.n105 585
R75 B.n840 B.n105 585
R76 B.n822 B.n104 585
R77 B.n841 B.n104 585
R78 B.n821 B.n820 585
R79 B.n820 B.n100 585
R80 B.n819 B.n99 585
R81 B.n847 B.n99 585
R82 B.n818 B.n98 585
R83 B.n848 B.n98 585
R84 B.n817 B.n97 585
R85 B.n849 B.n97 585
R86 B.n816 B.n815 585
R87 B.n815 B.n93 585
R88 B.n814 B.n92 585
R89 B.n855 B.n92 585
R90 B.n813 B.n91 585
R91 B.n856 B.n91 585
R92 B.n812 B.n90 585
R93 B.n857 B.n90 585
R94 B.n811 B.n810 585
R95 B.n810 B.n86 585
R96 B.n809 B.n85 585
R97 B.n863 B.n85 585
R98 B.n808 B.n84 585
R99 B.n864 B.n84 585
R100 B.n807 B.n83 585
R101 B.n865 B.n83 585
R102 B.n806 B.n805 585
R103 B.n805 B.n79 585
R104 B.n804 B.n78 585
R105 B.n871 B.n78 585
R106 B.n803 B.n77 585
R107 B.n872 B.n77 585
R108 B.n802 B.n76 585
R109 B.n873 B.n76 585
R110 B.n801 B.n800 585
R111 B.n800 B.n72 585
R112 B.n799 B.n71 585
R113 B.n879 B.n71 585
R114 B.n798 B.n70 585
R115 B.n880 B.n70 585
R116 B.n797 B.n69 585
R117 B.n881 B.n69 585
R118 B.n796 B.n795 585
R119 B.n795 B.n65 585
R120 B.n794 B.n64 585
R121 B.n887 B.n64 585
R122 B.n793 B.n63 585
R123 B.n888 B.n63 585
R124 B.n792 B.n62 585
R125 B.n889 B.n62 585
R126 B.n791 B.n790 585
R127 B.n790 B.n58 585
R128 B.n789 B.n57 585
R129 B.n895 B.n57 585
R130 B.n788 B.n56 585
R131 B.n896 B.n56 585
R132 B.n787 B.n55 585
R133 B.n897 B.n55 585
R134 B.n786 B.n785 585
R135 B.n785 B.n51 585
R136 B.n784 B.n50 585
R137 B.n903 B.n50 585
R138 B.n783 B.n49 585
R139 B.n904 B.n49 585
R140 B.n782 B.n48 585
R141 B.n905 B.n48 585
R142 B.n781 B.n780 585
R143 B.n780 B.n44 585
R144 B.n779 B.n43 585
R145 B.n911 B.n43 585
R146 B.n778 B.n42 585
R147 B.n912 B.n42 585
R148 B.n777 B.n41 585
R149 B.n913 B.n41 585
R150 B.n776 B.n775 585
R151 B.n775 B.n37 585
R152 B.n774 B.n36 585
R153 B.n919 B.n36 585
R154 B.n773 B.n35 585
R155 B.n920 B.n35 585
R156 B.n772 B.n34 585
R157 B.n921 B.n34 585
R158 B.n771 B.n770 585
R159 B.n770 B.n33 585
R160 B.n769 B.n29 585
R161 B.n927 B.n29 585
R162 B.n768 B.n28 585
R163 B.n928 B.n28 585
R164 B.n767 B.n27 585
R165 B.n929 B.n27 585
R166 B.n766 B.n765 585
R167 B.n765 B.n23 585
R168 B.n764 B.n22 585
R169 B.n935 B.n22 585
R170 B.n763 B.n21 585
R171 B.n936 B.n21 585
R172 B.n762 B.n20 585
R173 B.n937 B.n20 585
R174 B.n761 B.n760 585
R175 B.n760 B.n16 585
R176 B.n759 B.n15 585
R177 B.n943 B.n15 585
R178 B.n758 B.n14 585
R179 B.n944 B.n14 585
R180 B.n757 B.n13 585
R181 B.n945 B.n13 585
R182 B.n756 B.n755 585
R183 B.n755 B.n12 585
R184 B.n754 B.n753 585
R185 B.n754 B.n8 585
R186 B.n752 B.n7 585
R187 B.n952 B.n7 585
R188 B.n751 B.n6 585
R189 B.n953 B.n6 585
R190 B.n750 B.n5 585
R191 B.n954 B.n5 585
R192 B.n749 B.n748 585
R193 B.n748 B.n4 585
R194 B.n747 B.n279 585
R195 B.n747 B.n746 585
R196 B.n737 B.n280 585
R197 B.n281 B.n280 585
R198 B.n739 B.n738 585
R199 B.n740 B.n739 585
R200 B.n736 B.n286 585
R201 B.n286 B.n285 585
R202 B.n735 B.n734 585
R203 B.n734 B.n733 585
R204 B.n288 B.n287 585
R205 B.n289 B.n288 585
R206 B.n726 B.n725 585
R207 B.n727 B.n726 585
R208 B.n724 B.n294 585
R209 B.n294 B.n293 585
R210 B.n723 B.n722 585
R211 B.n722 B.n721 585
R212 B.n296 B.n295 585
R213 B.n297 B.n296 585
R214 B.n714 B.n713 585
R215 B.n715 B.n714 585
R216 B.n712 B.n302 585
R217 B.n302 B.n301 585
R218 B.n711 B.n710 585
R219 B.n710 B.n709 585
R220 B.n304 B.n303 585
R221 B.n702 B.n304 585
R222 B.n701 B.n700 585
R223 B.n703 B.n701 585
R224 B.n699 B.n309 585
R225 B.n309 B.n308 585
R226 B.n698 B.n697 585
R227 B.n697 B.n696 585
R228 B.n311 B.n310 585
R229 B.n312 B.n311 585
R230 B.n689 B.n688 585
R231 B.n690 B.n689 585
R232 B.n687 B.n317 585
R233 B.n317 B.n316 585
R234 B.n686 B.n685 585
R235 B.n685 B.n684 585
R236 B.n319 B.n318 585
R237 B.n320 B.n319 585
R238 B.n677 B.n676 585
R239 B.n678 B.n677 585
R240 B.n675 B.n325 585
R241 B.n325 B.n324 585
R242 B.n674 B.n673 585
R243 B.n673 B.n672 585
R244 B.n327 B.n326 585
R245 B.n328 B.n327 585
R246 B.n665 B.n664 585
R247 B.n666 B.n665 585
R248 B.n663 B.n333 585
R249 B.n333 B.n332 585
R250 B.n662 B.n661 585
R251 B.n661 B.n660 585
R252 B.n335 B.n334 585
R253 B.n336 B.n335 585
R254 B.n653 B.n652 585
R255 B.n654 B.n653 585
R256 B.n651 B.n340 585
R257 B.n344 B.n340 585
R258 B.n650 B.n649 585
R259 B.n649 B.n648 585
R260 B.n342 B.n341 585
R261 B.n343 B.n342 585
R262 B.n641 B.n640 585
R263 B.n642 B.n641 585
R264 B.n639 B.n349 585
R265 B.n349 B.n348 585
R266 B.n638 B.n637 585
R267 B.n637 B.n636 585
R268 B.n351 B.n350 585
R269 B.n352 B.n351 585
R270 B.n629 B.n628 585
R271 B.n630 B.n629 585
R272 B.n627 B.n357 585
R273 B.n357 B.n356 585
R274 B.n626 B.n625 585
R275 B.n625 B.n624 585
R276 B.n359 B.n358 585
R277 B.n360 B.n359 585
R278 B.n617 B.n616 585
R279 B.n618 B.n617 585
R280 B.n615 B.n365 585
R281 B.n365 B.n364 585
R282 B.n614 B.n613 585
R283 B.n613 B.n612 585
R284 B.n367 B.n366 585
R285 B.n368 B.n367 585
R286 B.n605 B.n604 585
R287 B.n606 B.n605 585
R288 B.n603 B.n373 585
R289 B.n373 B.n372 585
R290 B.n602 B.n601 585
R291 B.n601 B.n600 585
R292 B.n375 B.n374 585
R293 B.n376 B.n375 585
R294 B.n593 B.n592 585
R295 B.n594 B.n593 585
R296 B.n591 B.n381 585
R297 B.n381 B.n380 585
R298 B.n590 B.n589 585
R299 B.n589 B.n588 585
R300 B.n383 B.n382 585
R301 B.n384 B.n383 585
R302 B.n581 B.n580 585
R303 B.n582 B.n581 585
R304 B.n579 B.n389 585
R305 B.n389 B.n388 585
R306 B.n578 B.n577 585
R307 B.n577 B.n576 585
R308 B.n391 B.n390 585
R309 B.n392 B.n391 585
R310 B.n569 B.n568 585
R311 B.n570 B.n569 585
R312 B.n567 B.n397 585
R313 B.n397 B.n396 585
R314 B.n561 B.n560 585
R315 B.n559 B.n431 585
R316 B.n558 B.n430 585
R317 B.n563 B.n430 585
R318 B.n557 B.n556 585
R319 B.n555 B.n554 585
R320 B.n553 B.n552 585
R321 B.n551 B.n550 585
R322 B.n549 B.n548 585
R323 B.n547 B.n546 585
R324 B.n545 B.n544 585
R325 B.n543 B.n542 585
R326 B.n541 B.n540 585
R327 B.n539 B.n538 585
R328 B.n537 B.n536 585
R329 B.n535 B.n534 585
R330 B.n533 B.n532 585
R331 B.n531 B.n530 585
R332 B.n529 B.n528 585
R333 B.n527 B.n526 585
R334 B.n525 B.n524 585
R335 B.n523 B.n522 585
R336 B.n521 B.n520 585
R337 B.n519 B.n518 585
R338 B.n517 B.n516 585
R339 B.n515 B.n514 585
R340 B.n513 B.n512 585
R341 B.n511 B.n510 585
R342 B.n509 B.n508 585
R343 B.n506 B.n505 585
R344 B.n504 B.n503 585
R345 B.n502 B.n501 585
R346 B.n500 B.n499 585
R347 B.n498 B.n497 585
R348 B.n496 B.n495 585
R349 B.n494 B.n493 585
R350 B.n492 B.n491 585
R351 B.n490 B.n489 585
R352 B.n488 B.n487 585
R353 B.n486 B.n485 585
R354 B.n484 B.n483 585
R355 B.n482 B.n481 585
R356 B.n480 B.n479 585
R357 B.n478 B.n477 585
R358 B.n476 B.n475 585
R359 B.n474 B.n473 585
R360 B.n472 B.n471 585
R361 B.n470 B.n469 585
R362 B.n468 B.n467 585
R363 B.n466 B.n465 585
R364 B.n464 B.n463 585
R365 B.n462 B.n461 585
R366 B.n460 B.n459 585
R367 B.n458 B.n457 585
R368 B.n456 B.n455 585
R369 B.n454 B.n453 585
R370 B.n452 B.n451 585
R371 B.n450 B.n449 585
R372 B.n448 B.n447 585
R373 B.n446 B.n445 585
R374 B.n444 B.n443 585
R375 B.n442 B.n441 585
R376 B.n440 B.n439 585
R377 B.n438 B.n437 585
R378 B.n399 B.n398 585
R379 B.n566 B.n565 585
R380 B.n395 B.n394 585
R381 B.n396 B.n395 585
R382 B.n572 B.n571 585
R383 B.n571 B.n570 585
R384 B.n573 B.n393 585
R385 B.n393 B.n392 585
R386 B.n575 B.n574 585
R387 B.n576 B.n575 585
R388 B.n387 B.n386 585
R389 B.n388 B.n387 585
R390 B.n584 B.n583 585
R391 B.n583 B.n582 585
R392 B.n585 B.n385 585
R393 B.n385 B.n384 585
R394 B.n587 B.n586 585
R395 B.n588 B.n587 585
R396 B.n379 B.n378 585
R397 B.n380 B.n379 585
R398 B.n596 B.n595 585
R399 B.n595 B.n594 585
R400 B.n597 B.n377 585
R401 B.n377 B.n376 585
R402 B.n599 B.n598 585
R403 B.n600 B.n599 585
R404 B.n371 B.n370 585
R405 B.n372 B.n371 585
R406 B.n608 B.n607 585
R407 B.n607 B.n606 585
R408 B.n609 B.n369 585
R409 B.n369 B.n368 585
R410 B.n611 B.n610 585
R411 B.n612 B.n611 585
R412 B.n363 B.n362 585
R413 B.n364 B.n363 585
R414 B.n620 B.n619 585
R415 B.n619 B.n618 585
R416 B.n621 B.n361 585
R417 B.n361 B.n360 585
R418 B.n623 B.n622 585
R419 B.n624 B.n623 585
R420 B.n355 B.n354 585
R421 B.n356 B.n355 585
R422 B.n632 B.n631 585
R423 B.n631 B.n630 585
R424 B.n633 B.n353 585
R425 B.n353 B.n352 585
R426 B.n635 B.n634 585
R427 B.n636 B.n635 585
R428 B.n347 B.n346 585
R429 B.n348 B.n347 585
R430 B.n644 B.n643 585
R431 B.n643 B.n642 585
R432 B.n645 B.n345 585
R433 B.n345 B.n343 585
R434 B.n647 B.n646 585
R435 B.n648 B.n647 585
R436 B.n339 B.n338 585
R437 B.n344 B.n339 585
R438 B.n656 B.n655 585
R439 B.n655 B.n654 585
R440 B.n657 B.n337 585
R441 B.n337 B.n336 585
R442 B.n659 B.n658 585
R443 B.n660 B.n659 585
R444 B.n331 B.n330 585
R445 B.n332 B.n331 585
R446 B.n668 B.n667 585
R447 B.n667 B.n666 585
R448 B.n669 B.n329 585
R449 B.n329 B.n328 585
R450 B.n671 B.n670 585
R451 B.n672 B.n671 585
R452 B.n323 B.n322 585
R453 B.n324 B.n323 585
R454 B.n680 B.n679 585
R455 B.n679 B.n678 585
R456 B.n681 B.n321 585
R457 B.n321 B.n320 585
R458 B.n683 B.n682 585
R459 B.n684 B.n683 585
R460 B.n315 B.n314 585
R461 B.n316 B.n315 585
R462 B.n692 B.n691 585
R463 B.n691 B.n690 585
R464 B.n693 B.n313 585
R465 B.n313 B.n312 585
R466 B.n695 B.n694 585
R467 B.n696 B.n695 585
R468 B.n307 B.n306 585
R469 B.n308 B.n307 585
R470 B.n705 B.n704 585
R471 B.n704 B.n703 585
R472 B.n706 B.n305 585
R473 B.n702 B.n305 585
R474 B.n708 B.n707 585
R475 B.n709 B.n708 585
R476 B.n300 B.n299 585
R477 B.n301 B.n300 585
R478 B.n717 B.n716 585
R479 B.n716 B.n715 585
R480 B.n718 B.n298 585
R481 B.n298 B.n297 585
R482 B.n720 B.n719 585
R483 B.n721 B.n720 585
R484 B.n292 B.n291 585
R485 B.n293 B.n292 585
R486 B.n729 B.n728 585
R487 B.n728 B.n727 585
R488 B.n730 B.n290 585
R489 B.n290 B.n289 585
R490 B.n732 B.n731 585
R491 B.n733 B.n732 585
R492 B.n284 B.n283 585
R493 B.n285 B.n284 585
R494 B.n742 B.n741 585
R495 B.n741 B.n740 585
R496 B.n743 B.n282 585
R497 B.n282 B.n281 585
R498 B.n745 B.n744 585
R499 B.n746 B.n745 585
R500 B.n3 B.n0 585
R501 B.n4 B.n3 585
R502 B.n951 B.n1 585
R503 B.n952 B.n951 585
R504 B.n950 B.n949 585
R505 B.n950 B.n8 585
R506 B.n948 B.n9 585
R507 B.n12 B.n9 585
R508 B.n947 B.n946 585
R509 B.n946 B.n945 585
R510 B.n11 B.n10 585
R511 B.n944 B.n11 585
R512 B.n942 B.n941 585
R513 B.n943 B.n942 585
R514 B.n940 B.n17 585
R515 B.n17 B.n16 585
R516 B.n939 B.n938 585
R517 B.n938 B.n937 585
R518 B.n19 B.n18 585
R519 B.n936 B.n19 585
R520 B.n934 B.n933 585
R521 B.n935 B.n934 585
R522 B.n932 B.n24 585
R523 B.n24 B.n23 585
R524 B.n931 B.n930 585
R525 B.n930 B.n929 585
R526 B.n26 B.n25 585
R527 B.n928 B.n26 585
R528 B.n926 B.n925 585
R529 B.n927 B.n926 585
R530 B.n924 B.n30 585
R531 B.n33 B.n30 585
R532 B.n923 B.n922 585
R533 B.n922 B.n921 585
R534 B.n32 B.n31 585
R535 B.n920 B.n32 585
R536 B.n918 B.n917 585
R537 B.n919 B.n918 585
R538 B.n916 B.n38 585
R539 B.n38 B.n37 585
R540 B.n915 B.n914 585
R541 B.n914 B.n913 585
R542 B.n40 B.n39 585
R543 B.n912 B.n40 585
R544 B.n910 B.n909 585
R545 B.n911 B.n910 585
R546 B.n908 B.n45 585
R547 B.n45 B.n44 585
R548 B.n907 B.n906 585
R549 B.n906 B.n905 585
R550 B.n47 B.n46 585
R551 B.n904 B.n47 585
R552 B.n902 B.n901 585
R553 B.n903 B.n902 585
R554 B.n900 B.n52 585
R555 B.n52 B.n51 585
R556 B.n899 B.n898 585
R557 B.n898 B.n897 585
R558 B.n54 B.n53 585
R559 B.n896 B.n54 585
R560 B.n894 B.n893 585
R561 B.n895 B.n894 585
R562 B.n892 B.n59 585
R563 B.n59 B.n58 585
R564 B.n891 B.n890 585
R565 B.n890 B.n889 585
R566 B.n61 B.n60 585
R567 B.n888 B.n61 585
R568 B.n886 B.n885 585
R569 B.n887 B.n886 585
R570 B.n884 B.n66 585
R571 B.n66 B.n65 585
R572 B.n883 B.n882 585
R573 B.n882 B.n881 585
R574 B.n68 B.n67 585
R575 B.n880 B.n68 585
R576 B.n878 B.n877 585
R577 B.n879 B.n878 585
R578 B.n876 B.n73 585
R579 B.n73 B.n72 585
R580 B.n875 B.n874 585
R581 B.n874 B.n873 585
R582 B.n75 B.n74 585
R583 B.n872 B.n75 585
R584 B.n870 B.n869 585
R585 B.n871 B.n870 585
R586 B.n868 B.n80 585
R587 B.n80 B.n79 585
R588 B.n867 B.n866 585
R589 B.n866 B.n865 585
R590 B.n82 B.n81 585
R591 B.n864 B.n82 585
R592 B.n862 B.n861 585
R593 B.n863 B.n862 585
R594 B.n860 B.n87 585
R595 B.n87 B.n86 585
R596 B.n859 B.n858 585
R597 B.n858 B.n857 585
R598 B.n89 B.n88 585
R599 B.n856 B.n89 585
R600 B.n854 B.n853 585
R601 B.n855 B.n854 585
R602 B.n852 B.n94 585
R603 B.n94 B.n93 585
R604 B.n851 B.n850 585
R605 B.n850 B.n849 585
R606 B.n96 B.n95 585
R607 B.n848 B.n96 585
R608 B.n846 B.n845 585
R609 B.n847 B.n846 585
R610 B.n844 B.n101 585
R611 B.n101 B.n100 585
R612 B.n843 B.n842 585
R613 B.n842 B.n841 585
R614 B.n103 B.n102 585
R615 B.n840 B.n103 585
R616 B.n838 B.n837 585
R617 B.n839 B.n838 585
R618 B.n836 B.n108 585
R619 B.n108 B.n107 585
R620 B.n835 B.n834 585
R621 B.n834 B.n833 585
R622 B.n110 B.n109 585
R623 B.n832 B.n110 585
R624 B.n955 B.n954 585
R625 B.n953 B.n2 585
R626 B.n151 B.n110 569.379
R627 B.n830 B.n112 569.379
R628 B.n565 B.n397 569.379
R629 B.n561 B.n395 569.379
R630 B.n148 B.t14 273.392
R631 B.n146 B.t10 273.392
R632 B.n434 B.t17 273.392
R633 B.n432 B.t21 273.392
R634 B.n146 B.t12 260.738
R635 B.n434 B.t20 260.738
R636 B.n148 B.t15 260.738
R637 B.n432 B.t23 260.738
R638 B.n831 B.n144 256.663
R639 B.n831 B.n143 256.663
R640 B.n831 B.n142 256.663
R641 B.n831 B.n141 256.663
R642 B.n831 B.n140 256.663
R643 B.n831 B.n139 256.663
R644 B.n831 B.n138 256.663
R645 B.n831 B.n137 256.663
R646 B.n831 B.n136 256.663
R647 B.n831 B.n135 256.663
R648 B.n831 B.n134 256.663
R649 B.n831 B.n133 256.663
R650 B.n831 B.n132 256.663
R651 B.n831 B.n131 256.663
R652 B.n831 B.n130 256.663
R653 B.n831 B.n129 256.663
R654 B.n831 B.n128 256.663
R655 B.n831 B.n127 256.663
R656 B.n831 B.n126 256.663
R657 B.n831 B.n125 256.663
R658 B.n831 B.n124 256.663
R659 B.n831 B.n123 256.663
R660 B.n831 B.n122 256.663
R661 B.n831 B.n121 256.663
R662 B.n831 B.n120 256.663
R663 B.n831 B.n119 256.663
R664 B.n831 B.n118 256.663
R665 B.n831 B.n117 256.663
R666 B.n831 B.n116 256.663
R667 B.n831 B.n115 256.663
R668 B.n831 B.n114 256.663
R669 B.n831 B.n113 256.663
R670 B.n563 B.n562 256.663
R671 B.n563 B.n400 256.663
R672 B.n563 B.n401 256.663
R673 B.n563 B.n402 256.663
R674 B.n563 B.n403 256.663
R675 B.n563 B.n404 256.663
R676 B.n563 B.n405 256.663
R677 B.n563 B.n406 256.663
R678 B.n563 B.n407 256.663
R679 B.n563 B.n408 256.663
R680 B.n563 B.n409 256.663
R681 B.n563 B.n410 256.663
R682 B.n563 B.n411 256.663
R683 B.n563 B.n412 256.663
R684 B.n563 B.n413 256.663
R685 B.n563 B.n414 256.663
R686 B.n563 B.n415 256.663
R687 B.n563 B.n416 256.663
R688 B.n563 B.n417 256.663
R689 B.n563 B.n418 256.663
R690 B.n563 B.n419 256.663
R691 B.n563 B.n420 256.663
R692 B.n563 B.n421 256.663
R693 B.n563 B.n422 256.663
R694 B.n563 B.n423 256.663
R695 B.n563 B.n424 256.663
R696 B.n563 B.n425 256.663
R697 B.n563 B.n426 256.663
R698 B.n563 B.n427 256.663
R699 B.n563 B.n428 256.663
R700 B.n563 B.n429 256.663
R701 B.n564 B.n563 256.663
R702 B.n957 B.n956 256.663
R703 B.n147 B.t13 201.78
R704 B.n435 B.t19 201.78
R705 B.n149 B.t16 201.78
R706 B.n433 B.t22 201.78
R707 B.n155 B.n154 163.367
R708 B.n159 B.n158 163.367
R709 B.n163 B.n162 163.367
R710 B.n167 B.n166 163.367
R711 B.n171 B.n170 163.367
R712 B.n175 B.n174 163.367
R713 B.n179 B.n178 163.367
R714 B.n183 B.n182 163.367
R715 B.n187 B.n186 163.367
R716 B.n191 B.n190 163.367
R717 B.n195 B.n194 163.367
R718 B.n199 B.n198 163.367
R719 B.n203 B.n202 163.367
R720 B.n207 B.n206 163.367
R721 B.n211 B.n210 163.367
R722 B.n215 B.n214 163.367
R723 B.n219 B.n218 163.367
R724 B.n223 B.n222 163.367
R725 B.n228 B.n227 163.367
R726 B.n232 B.n231 163.367
R727 B.n236 B.n235 163.367
R728 B.n240 B.n239 163.367
R729 B.n244 B.n243 163.367
R730 B.n248 B.n247 163.367
R731 B.n252 B.n251 163.367
R732 B.n256 B.n255 163.367
R733 B.n260 B.n259 163.367
R734 B.n264 B.n263 163.367
R735 B.n268 B.n267 163.367
R736 B.n272 B.n271 163.367
R737 B.n276 B.n275 163.367
R738 B.n830 B.n145 163.367
R739 B.n569 B.n397 163.367
R740 B.n569 B.n391 163.367
R741 B.n577 B.n391 163.367
R742 B.n577 B.n389 163.367
R743 B.n581 B.n389 163.367
R744 B.n581 B.n383 163.367
R745 B.n589 B.n383 163.367
R746 B.n589 B.n381 163.367
R747 B.n593 B.n381 163.367
R748 B.n593 B.n375 163.367
R749 B.n601 B.n375 163.367
R750 B.n601 B.n373 163.367
R751 B.n605 B.n373 163.367
R752 B.n605 B.n367 163.367
R753 B.n613 B.n367 163.367
R754 B.n613 B.n365 163.367
R755 B.n617 B.n365 163.367
R756 B.n617 B.n359 163.367
R757 B.n625 B.n359 163.367
R758 B.n625 B.n357 163.367
R759 B.n629 B.n357 163.367
R760 B.n629 B.n351 163.367
R761 B.n637 B.n351 163.367
R762 B.n637 B.n349 163.367
R763 B.n641 B.n349 163.367
R764 B.n641 B.n342 163.367
R765 B.n649 B.n342 163.367
R766 B.n649 B.n340 163.367
R767 B.n653 B.n340 163.367
R768 B.n653 B.n335 163.367
R769 B.n661 B.n335 163.367
R770 B.n661 B.n333 163.367
R771 B.n665 B.n333 163.367
R772 B.n665 B.n327 163.367
R773 B.n673 B.n327 163.367
R774 B.n673 B.n325 163.367
R775 B.n677 B.n325 163.367
R776 B.n677 B.n319 163.367
R777 B.n685 B.n319 163.367
R778 B.n685 B.n317 163.367
R779 B.n689 B.n317 163.367
R780 B.n689 B.n311 163.367
R781 B.n697 B.n311 163.367
R782 B.n697 B.n309 163.367
R783 B.n701 B.n309 163.367
R784 B.n701 B.n304 163.367
R785 B.n710 B.n304 163.367
R786 B.n710 B.n302 163.367
R787 B.n714 B.n302 163.367
R788 B.n714 B.n296 163.367
R789 B.n722 B.n296 163.367
R790 B.n722 B.n294 163.367
R791 B.n726 B.n294 163.367
R792 B.n726 B.n288 163.367
R793 B.n734 B.n288 163.367
R794 B.n734 B.n286 163.367
R795 B.n739 B.n286 163.367
R796 B.n739 B.n280 163.367
R797 B.n747 B.n280 163.367
R798 B.n748 B.n747 163.367
R799 B.n748 B.n5 163.367
R800 B.n6 B.n5 163.367
R801 B.n7 B.n6 163.367
R802 B.n754 B.n7 163.367
R803 B.n755 B.n754 163.367
R804 B.n755 B.n13 163.367
R805 B.n14 B.n13 163.367
R806 B.n15 B.n14 163.367
R807 B.n760 B.n15 163.367
R808 B.n760 B.n20 163.367
R809 B.n21 B.n20 163.367
R810 B.n22 B.n21 163.367
R811 B.n765 B.n22 163.367
R812 B.n765 B.n27 163.367
R813 B.n28 B.n27 163.367
R814 B.n29 B.n28 163.367
R815 B.n770 B.n29 163.367
R816 B.n770 B.n34 163.367
R817 B.n35 B.n34 163.367
R818 B.n36 B.n35 163.367
R819 B.n775 B.n36 163.367
R820 B.n775 B.n41 163.367
R821 B.n42 B.n41 163.367
R822 B.n43 B.n42 163.367
R823 B.n780 B.n43 163.367
R824 B.n780 B.n48 163.367
R825 B.n49 B.n48 163.367
R826 B.n50 B.n49 163.367
R827 B.n785 B.n50 163.367
R828 B.n785 B.n55 163.367
R829 B.n56 B.n55 163.367
R830 B.n57 B.n56 163.367
R831 B.n790 B.n57 163.367
R832 B.n790 B.n62 163.367
R833 B.n63 B.n62 163.367
R834 B.n64 B.n63 163.367
R835 B.n795 B.n64 163.367
R836 B.n795 B.n69 163.367
R837 B.n70 B.n69 163.367
R838 B.n71 B.n70 163.367
R839 B.n800 B.n71 163.367
R840 B.n800 B.n76 163.367
R841 B.n77 B.n76 163.367
R842 B.n78 B.n77 163.367
R843 B.n805 B.n78 163.367
R844 B.n805 B.n83 163.367
R845 B.n84 B.n83 163.367
R846 B.n85 B.n84 163.367
R847 B.n810 B.n85 163.367
R848 B.n810 B.n90 163.367
R849 B.n91 B.n90 163.367
R850 B.n92 B.n91 163.367
R851 B.n815 B.n92 163.367
R852 B.n815 B.n97 163.367
R853 B.n98 B.n97 163.367
R854 B.n99 B.n98 163.367
R855 B.n820 B.n99 163.367
R856 B.n820 B.n104 163.367
R857 B.n105 B.n104 163.367
R858 B.n106 B.n105 163.367
R859 B.n825 B.n106 163.367
R860 B.n825 B.n111 163.367
R861 B.n112 B.n111 163.367
R862 B.n431 B.n430 163.367
R863 B.n556 B.n430 163.367
R864 B.n554 B.n553 163.367
R865 B.n550 B.n549 163.367
R866 B.n546 B.n545 163.367
R867 B.n542 B.n541 163.367
R868 B.n538 B.n537 163.367
R869 B.n534 B.n533 163.367
R870 B.n530 B.n529 163.367
R871 B.n526 B.n525 163.367
R872 B.n522 B.n521 163.367
R873 B.n518 B.n517 163.367
R874 B.n514 B.n513 163.367
R875 B.n510 B.n509 163.367
R876 B.n505 B.n504 163.367
R877 B.n501 B.n500 163.367
R878 B.n497 B.n496 163.367
R879 B.n493 B.n492 163.367
R880 B.n489 B.n488 163.367
R881 B.n485 B.n484 163.367
R882 B.n481 B.n480 163.367
R883 B.n477 B.n476 163.367
R884 B.n473 B.n472 163.367
R885 B.n469 B.n468 163.367
R886 B.n465 B.n464 163.367
R887 B.n461 B.n460 163.367
R888 B.n457 B.n456 163.367
R889 B.n453 B.n452 163.367
R890 B.n449 B.n448 163.367
R891 B.n445 B.n444 163.367
R892 B.n441 B.n440 163.367
R893 B.n437 B.n399 163.367
R894 B.n571 B.n395 163.367
R895 B.n571 B.n393 163.367
R896 B.n575 B.n393 163.367
R897 B.n575 B.n387 163.367
R898 B.n583 B.n387 163.367
R899 B.n583 B.n385 163.367
R900 B.n587 B.n385 163.367
R901 B.n587 B.n379 163.367
R902 B.n595 B.n379 163.367
R903 B.n595 B.n377 163.367
R904 B.n599 B.n377 163.367
R905 B.n599 B.n371 163.367
R906 B.n607 B.n371 163.367
R907 B.n607 B.n369 163.367
R908 B.n611 B.n369 163.367
R909 B.n611 B.n363 163.367
R910 B.n619 B.n363 163.367
R911 B.n619 B.n361 163.367
R912 B.n623 B.n361 163.367
R913 B.n623 B.n355 163.367
R914 B.n631 B.n355 163.367
R915 B.n631 B.n353 163.367
R916 B.n635 B.n353 163.367
R917 B.n635 B.n347 163.367
R918 B.n643 B.n347 163.367
R919 B.n643 B.n345 163.367
R920 B.n647 B.n345 163.367
R921 B.n647 B.n339 163.367
R922 B.n655 B.n339 163.367
R923 B.n655 B.n337 163.367
R924 B.n659 B.n337 163.367
R925 B.n659 B.n331 163.367
R926 B.n667 B.n331 163.367
R927 B.n667 B.n329 163.367
R928 B.n671 B.n329 163.367
R929 B.n671 B.n323 163.367
R930 B.n679 B.n323 163.367
R931 B.n679 B.n321 163.367
R932 B.n683 B.n321 163.367
R933 B.n683 B.n315 163.367
R934 B.n691 B.n315 163.367
R935 B.n691 B.n313 163.367
R936 B.n695 B.n313 163.367
R937 B.n695 B.n307 163.367
R938 B.n704 B.n307 163.367
R939 B.n704 B.n305 163.367
R940 B.n708 B.n305 163.367
R941 B.n708 B.n300 163.367
R942 B.n716 B.n300 163.367
R943 B.n716 B.n298 163.367
R944 B.n720 B.n298 163.367
R945 B.n720 B.n292 163.367
R946 B.n728 B.n292 163.367
R947 B.n728 B.n290 163.367
R948 B.n732 B.n290 163.367
R949 B.n732 B.n284 163.367
R950 B.n741 B.n284 163.367
R951 B.n741 B.n282 163.367
R952 B.n745 B.n282 163.367
R953 B.n745 B.n3 163.367
R954 B.n955 B.n3 163.367
R955 B.n951 B.n2 163.367
R956 B.n951 B.n950 163.367
R957 B.n950 B.n9 163.367
R958 B.n946 B.n9 163.367
R959 B.n946 B.n11 163.367
R960 B.n942 B.n11 163.367
R961 B.n942 B.n17 163.367
R962 B.n938 B.n17 163.367
R963 B.n938 B.n19 163.367
R964 B.n934 B.n19 163.367
R965 B.n934 B.n24 163.367
R966 B.n930 B.n24 163.367
R967 B.n930 B.n26 163.367
R968 B.n926 B.n26 163.367
R969 B.n926 B.n30 163.367
R970 B.n922 B.n30 163.367
R971 B.n922 B.n32 163.367
R972 B.n918 B.n32 163.367
R973 B.n918 B.n38 163.367
R974 B.n914 B.n38 163.367
R975 B.n914 B.n40 163.367
R976 B.n910 B.n40 163.367
R977 B.n910 B.n45 163.367
R978 B.n906 B.n45 163.367
R979 B.n906 B.n47 163.367
R980 B.n902 B.n47 163.367
R981 B.n902 B.n52 163.367
R982 B.n898 B.n52 163.367
R983 B.n898 B.n54 163.367
R984 B.n894 B.n54 163.367
R985 B.n894 B.n59 163.367
R986 B.n890 B.n59 163.367
R987 B.n890 B.n61 163.367
R988 B.n886 B.n61 163.367
R989 B.n886 B.n66 163.367
R990 B.n882 B.n66 163.367
R991 B.n882 B.n68 163.367
R992 B.n878 B.n68 163.367
R993 B.n878 B.n73 163.367
R994 B.n874 B.n73 163.367
R995 B.n874 B.n75 163.367
R996 B.n870 B.n75 163.367
R997 B.n870 B.n80 163.367
R998 B.n866 B.n80 163.367
R999 B.n866 B.n82 163.367
R1000 B.n862 B.n82 163.367
R1001 B.n862 B.n87 163.367
R1002 B.n858 B.n87 163.367
R1003 B.n858 B.n89 163.367
R1004 B.n854 B.n89 163.367
R1005 B.n854 B.n94 163.367
R1006 B.n850 B.n94 163.367
R1007 B.n850 B.n96 163.367
R1008 B.n846 B.n96 163.367
R1009 B.n846 B.n101 163.367
R1010 B.n842 B.n101 163.367
R1011 B.n842 B.n103 163.367
R1012 B.n838 B.n103 163.367
R1013 B.n838 B.n108 163.367
R1014 B.n834 B.n108 163.367
R1015 B.n834 B.n110 163.367
R1016 B.n563 B.n396 123.046
R1017 B.n832 B.n831 123.046
R1018 B.n151 B.n113 71.676
R1019 B.n155 B.n114 71.676
R1020 B.n159 B.n115 71.676
R1021 B.n163 B.n116 71.676
R1022 B.n167 B.n117 71.676
R1023 B.n171 B.n118 71.676
R1024 B.n175 B.n119 71.676
R1025 B.n179 B.n120 71.676
R1026 B.n183 B.n121 71.676
R1027 B.n187 B.n122 71.676
R1028 B.n191 B.n123 71.676
R1029 B.n195 B.n124 71.676
R1030 B.n199 B.n125 71.676
R1031 B.n203 B.n126 71.676
R1032 B.n207 B.n127 71.676
R1033 B.n211 B.n128 71.676
R1034 B.n215 B.n129 71.676
R1035 B.n219 B.n130 71.676
R1036 B.n223 B.n131 71.676
R1037 B.n228 B.n132 71.676
R1038 B.n232 B.n133 71.676
R1039 B.n236 B.n134 71.676
R1040 B.n240 B.n135 71.676
R1041 B.n244 B.n136 71.676
R1042 B.n248 B.n137 71.676
R1043 B.n252 B.n138 71.676
R1044 B.n256 B.n139 71.676
R1045 B.n260 B.n140 71.676
R1046 B.n264 B.n141 71.676
R1047 B.n268 B.n142 71.676
R1048 B.n272 B.n143 71.676
R1049 B.n276 B.n144 71.676
R1050 B.n145 B.n144 71.676
R1051 B.n275 B.n143 71.676
R1052 B.n271 B.n142 71.676
R1053 B.n267 B.n141 71.676
R1054 B.n263 B.n140 71.676
R1055 B.n259 B.n139 71.676
R1056 B.n255 B.n138 71.676
R1057 B.n251 B.n137 71.676
R1058 B.n247 B.n136 71.676
R1059 B.n243 B.n135 71.676
R1060 B.n239 B.n134 71.676
R1061 B.n235 B.n133 71.676
R1062 B.n231 B.n132 71.676
R1063 B.n227 B.n131 71.676
R1064 B.n222 B.n130 71.676
R1065 B.n218 B.n129 71.676
R1066 B.n214 B.n128 71.676
R1067 B.n210 B.n127 71.676
R1068 B.n206 B.n126 71.676
R1069 B.n202 B.n125 71.676
R1070 B.n198 B.n124 71.676
R1071 B.n194 B.n123 71.676
R1072 B.n190 B.n122 71.676
R1073 B.n186 B.n121 71.676
R1074 B.n182 B.n120 71.676
R1075 B.n178 B.n119 71.676
R1076 B.n174 B.n118 71.676
R1077 B.n170 B.n117 71.676
R1078 B.n166 B.n116 71.676
R1079 B.n162 B.n115 71.676
R1080 B.n158 B.n114 71.676
R1081 B.n154 B.n113 71.676
R1082 B.n562 B.n561 71.676
R1083 B.n556 B.n400 71.676
R1084 B.n553 B.n401 71.676
R1085 B.n549 B.n402 71.676
R1086 B.n545 B.n403 71.676
R1087 B.n541 B.n404 71.676
R1088 B.n537 B.n405 71.676
R1089 B.n533 B.n406 71.676
R1090 B.n529 B.n407 71.676
R1091 B.n525 B.n408 71.676
R1092 B.n521 B.n409 71.676
R1093 B.n517 B.n410 71.676
R1094 B.n513 B.n411 71.676
R1095 B.n509 B.n412 71.676
R1096 B.n504 B.n413 71.676
R1097 B.n500 B.n414 71.676
R1098 B.n496 B.n415 71.676
R1099 B.n492 B.n416 71.676
R1100 B.n488 B.n417 71.676
R1101 B.n484 B.n418 71.676
R1102 B.n480 B.n419 71.676
R1103 B.n476 B.n420 71.676
R1104 B.n472 B.n421 71.676
R1105 B.n468 B.n422 71.676
R1106 B.n464 B.n423 71.676
R1107 B.n460 B.n424 71.676
R1108 B.n456 B.n425 71.676
R1109 B.n452 B.n426 71.676
R1110 B.n448 B.n427 71.676
R1111 B.n444 B.n428 71.676
R1112 B.n440 B.n429 71.676
R1113 B.n564 B.n399 71.676
R1114 B.n562 B.n431 71.676
R1115 B.n554 B.n400 71.676
R1116 B.n550 B.n401 71.676
R1117 B.n546 B.n402 71.676
R1118 B.n542 B.n403 71.676
R1119 B.n538 B.n404 71.676
R1120 B.n534 B.n405 71.676
R1121 B.n530 B.n406 71.676
R1122 B.n526 B.n407 71.676
R1123 B.n522 B.n408 71.676
R1124 B.n518 B.n409 71.676
R1125 B.n514 B.n410 71.676
R1126 B.n510 B.n411 71.676
R1127 B.n505 B.n412 71.676
R1128 B.n501 B.n413 71.676
R1129 B.n497 B.n414 71.676
R1130 B.n493 B.n415 71.676
R1131 B.n489 B.n416 71.676
R1132 B.n485 B.n417 71.676
R1133 B.n481 B.n418 71.676
R1134 B.n477 B.n419 71.676
R1135 B.n473 B.n420 71.676
R1136 B.n469 B.n421 71.676
R1137 B.n465 B.n422 71.676
R1138 B.n461 B.n423 71.676
R1139 B.n457 B.n424 71.676
R1140 B.n453 B.n425 71.676
R1141 B.n449 B.n426 71.676
R1142 B.n445 B.n427 71.676
R1143 B.n441 B.n428 71.676
R1144 B.n437 B.n429 71.676
R1145 B.n565 B.n564 71.676
R1146 B.n956 B.n955 71.676
R1147 B.n956 B.n2 71.676
R1148 B.n150 B.n149 59.5399
R1149 B.n225 B.n147 59.5399
R1150 B.n436 B.n435 59.5399
R1151 B.n507 B.n433 59.5399
R1152 B.n570 B.n396 59.342
R1153 B.n570 B.n392 59.342
R1154 B.n576 B.n392 59.342
R1155 B.n576 B.n388 59.342
R1156 B.n582 B.n388 59.342
R1157 B.n582 B.n384 59.342
R1158 B.n588 B.n384 59.342
R1159 B.n594 B.n380 59.342
R1160 B.n594 B.n376 59.342
R1161 B.n600 B.n376 59.342
R1162 B.n600 B.n372 59.342
R1163 B.n606 B.n372 59.342
R1164 B.n606 B.n368 59.342
R1165 B.n612 B.n368 59.342
R1166 B.n612 B.n364 59.342
R1167 B.n618 B.n364 59.342
R1168 B.n618 B.n360 59.342
R1169 B.n624 B.n360 59.342
R1170 B.n630 B.n356 59.342
R1171 B.n630 B.n352 59.342
R1172 B.n636 B.n352 59.342
R1173 B.n636 B.n348 59.342
R1174 B.n642 B.n348 59.342
R1175 B.n642 B.n343 59.342
R1176 B.n648 B.n343 59.342
R1177 B.n648 B.n344 59.342
R1178 B.n654 B.n336 59.342
R1179 B.n660 B.n336 59.342
R1180 B.n660 B.n332 59.342
R1181 B.n666 B.n332 59.342
R1182 B.n666 B.n328 59.342
R1183 B.n672 B.n328 59.342
R1184 B.n672 B.n324 59.342
R1185 B.n678 B.n324 59.342
R1186 B.n684 B.n320 59.342
R1187 B.n684 B.n316 59.342
R1188 B.n690 B.n316 59.342
R1189 B.n690 B.n312 59.342
R1190 B.n696 B.n312 59.342
R1191 B.n696 B.n308 59.342
R1192 B.n703 B.n308 59.342
R1193 B.n703 B.n702 59.342
R1194 B.n709 B.n301 59.342
R1195 B.n715 B.n301 59.342
R1196 B.n715 B.n297 59.342
R1197 B.n721 B.n297 59.342
R1198 B.n721 B.n293 59.342
R1199 B.n727 B.n293 59.342
R1200 B.n727 B.n289 59.342
R1201 B.n733 B.n289 59.342
R1202 B.n740 B.n285 59.342
R1203 B.n740 B.n281 59.342
R1204 B.n746 B.n281 59.342
R1205 B.n746 B.n4 59.342
R1206 B.n954 B.n4 59.342
R1207 B.n954 B.n953 59.342
R1208 B.n953 B.n952 59.342
R1209 B.n952 B.n8 59.342
R1210 B.n12 B.n8 59.342
R1211 B.n945 B.n12 59.342
R1212 B.n945 B.n944 59.342
R1213 B.n943 B.n16 59.342
R1214 B.n937 B.n16 59.342
R1215 B.n937 B.n936 59.342
R1216 B.n936 B.n935 59.342
R1217 B.n935 B.n23 59.342
R1218 B.n929 B.n23 59.342
R1219 B.n929 B.n928 59.342
R1220 B.n928 B.n927 59.342
R1221 B.n921 B.n33 59.342
R1222 B.n921 B.n920 59.342
R1223 B.n920 B.n919 59.342
R1224 B.n919 B.n37 59.342
R1225 B.n913 B.n37 59.342
R1226 B.n913 B.n912 59.342
R1227 B.n912 B.n911 59.342
R1228 B.n911 B.n44 59.342
R1229 B.n905 B.n904 59.342
R1230 B.n904 B.n903 59.342
R1231 B.n903 B.n51 59.342
R1232 B.n897 B.n51 59.342
R1233 B.n897 B.n896 59.342
R1234 B.n896 B.n895 59.342
R1235 B.n895 B.n58 59.342
R1236 B.n889 B.n58 59.342
R1237 B.n888 B.n887 59.342
R1238 B.n887 B.n65 59.342
R1239 B.n881 B.n65 59.342
R1240 B.n881 B.n880 59.342
R1241 B.n880 B.n879 59.342
R1242 B.n879 B.n72 59.342
R1243 B.n873 B.n72 59.342
R1244 B.n873 B.n872 59.342
R1245 B.n871 B.n79 59.342
R1246 B.n865 B.n79 59.342
R1247 B.n865 B.n864 59.342
R1248 B.n864 B.n863 59.342
R1249 B.n863 B.n86 59.342
R1250 B.n857 B.n86 59.342
R1251 B.n857 B.n856 59.342
R1252 B.n856 B.n855 59.342
R1253 B.n855 B.n93 59.342
R1254 B.n849 B.n93 59.342
R1255 B.n849 B.n848 59.342
R1256 B.n847 B.n100 59.342
R1257 B.n841 B.n100 59.342
R1258 B.n841 B.n840 59.342
R1259 B.n840 B.n839 59.342
R1260 B.n839 B.n107 59.342
R1261 B.n833 B.n107 59.342
R1262 B.n833 B.n832 59.342
R1263 B.n149 B.n148 58.9581
R1264 B.n147 B.n146 58.9581
R1265 B.n435 B.n434 58.9581
R1266 B.n433 B.n432 58.9581
R1267 B.n624 B.t6 39.2706
R1268 B.t2 B.n871 39.2706
R1269 B.n560 B.n394 36.9956
R1270 B.n567 B.n566 36.9956
R1271 B.n829 B.n828 36.9956
R1272 B.n152 B.n109 36.9956
R1273 B.n344 B.t3 35.78
R1274 B.t4 B.n888 35.78
R1275 B.t9 B.n285 34.0346
R1276 B.n944 B.t0 34.0346
R1277 B.n678 B.t5 32.2893
R1278 B.n905 B.t7 32.2893
R1279 B.n588 B.t18 30.5439
R1280 B.n709 B.t1 30.5439
R1281 B.n927 B.t8 30.5439
R1282 B.t11 B.n847 30.5439
R1283 B.t18 B.n380 28.7986
R1284 B.n702 B.t1 28.7986
R1285 B.n33 B.t8 28.7986
R1286 B.n848 B.t11 28.7986
R1287 B.t5 B.n320 27.0533
R1288 B.t7 B.n44 27.0533
R1289 B.n733 B.t9 25.3079
R1290 B.t0 B.n943 25.3079
R1291 B.n654 B.t3 23.5626
R1292 B.n889 B.t4 23.5626
R1293 B.t6 B.n356 20.0719
R1294 B.n872 B.t2 20.0719
R1295 B B.n957 18.0485
R1296 B.n572 B.n394 10.6151
R1297 B.n573 B.n572 10.6151
R1298 B.n574 B.n573 10.6151
R1299 B.n574 B.n386 10.6151
R1300 B.n584 B.n386 10.6151
R1301 B.n585 B.n584 10.6151
R1302 B.n586 B.n585 10.6151
R1303 B.n586 B.n378 10.6151
R1304 B.n596 B.n378 10.6151
R1305 B.n597 B.n596 10.6151
R1306 B.n598 B.n597 10.6151
R1307 B.n598 B.n370 10.6151
R1308 B.n608 B.n370 10.6151
R1309 B.n609 B.n608 10.6151
R1310 B.n610 B.n609 10.6151
R1311 B.n610 B.n362 10.6151
R1312 B.n620 B.n362 10.6151
R1313 B.n621 B.n620 10.6151
R1314 B.n622 B.n621 10.6151
R1315 B.n622 B.n354 10.6151
R1316 B.n632 B.n354 10.6151
R1317 B.n633 B.n632 10.6151
R1318 B.n634 B.n633 10.6151
R1319 B.n634 B.n346 10.6151
R1320 B.n644 B.n346 10.6151
R1321 B.n645 B.n644 10.6151
R1322 B.n646 B.n645 10.6151
R1323 B.n646 B.n338 10.6151
R1324 B.n656 B.n338 10.6151
R1325 B.n657 B.n656 10.6151
R1326 B.n658 B.n657 10.6151
R1327 B.n658 B.n330 10.6151
R1328 B.n668 B.n330 10.6151
R1329 B.n669 B.n668 10.6151
R1330 B.n670 B.n669 10.6151
R1331 B.n670 B.n322 10.6151
R1332 B.n680 B.n322 10.6151
R1333 B.n681 B.n680 10.6151
R1334 B.n682 B.n681 10.6151
R1335 B.n682 B.n314 10.6151
R1336 B.n692 B.n314 10.6151
R1337 B.n693 B.n692 10.6151
R1338 B.n694 B.n693 10.6151
R1339 B.n694 B.n306 10.6151
R1340 B.n705 B.n306 10.6151
R1341 B.n706 B.n705 10.6151
R1342 B.n707 B.n706 10.6151
R1343 B.n707 B.n299 10.6151
R1344 B.n717 B.n299 10.6151
R1345 B.n718 B.n717 10.6151
R1346 B.n719 B.n718 10.6151
R1347 B.n719 B.n291 10.6151
R1348 B.n729 B.n291 10.6151
R1349 B.n730 B.n729 10.6151
R1350 B.n731 B.n730 10.6151
R1351 B.n731 B.n283 10.6151
R1352 B.n742 B.n283 10.6151
R1353 B.n743 B.n742 10.6151
R1354 B.n744 B.n743 10.6151
R1355 B.n744 B.n0 10.6151
R1356 B.n560 B.n559 10.6151
R1357 B.n559 B.n558 10.6151
R1358 B.n558 B.n557 10.6151
R1359 B.n557 B.n555 10.6151
R1360 B.n555 B.n552 10.6151
R1361 B.n552 B.n551 10.6151
R1362 B.n551 B.n548 10.6151
R1363 B.n548 B.n547 10.6151
R1364 B.n547 B.n544 10.6151
R1365 B.n544 B.n543 10.6151
R1366 B.n543 B.n540 10.6151
R1367 B.n540 B.n539 10.6151
R1368 B.n539 B.n536 10.6151
R1369 B.n536 B.n535 10.6151
R1370 B.n535 B.n532 10.6151
R1371 B.n532 B.n531 10.6151
R1372 B.n531 B.n528 10.6151
R1373 B.n528 B.n527 10.6151
R1374 B.n527 B.n524 10.6151
R1375 B.n524 B.n523 10.6151
R1376 B.n523 B.n520 10.6151
R1377 B.n520 B.n519 10.6151
R1378 B.n519 B.n516 10.6151
R1379 B.n516 B.n515 10.6151
R1380 B.n515 B.n512 10.6151
R1381 B.n512 B.n511 10.6151
R1382 B.n511 B.n508 10.6151
R1383 B.n506 B.n503 10.6151
R1384 B.n503 B.n502 10.6151
R1385 B.n502 B.n499 10.6151
R1386 B.n499 B.n498 10.6151
R1387 B.n498 B.n495 10.6151
R1388 B.n495 B.n494 10.6151
R1389 B.n494 B.n491 10.6151
R1390 B.n491 B.n490 10.6151
R1391 B.n487 B.n486 10.6151
R1392 B.n486 B.n483 10.6151
R1393 B.n483 B.n482 10.6151
R1394 B.n482 B.n479 10.6151
R1395 B.n479 B.n478 10.6151
R1396 B.n478 B.n475 10.6151
R1397 B.n475 B.n474 10.6151
R1398 B.n474 B.n471 10.6151
R1399 B.n471 B.n470 10.6151
R1400 B.n470 B.n467 10.6151
R1401 B.n467 B.n466 10.6151
R1402 B.n466 B.n463 10.6151
R1403 B.n463 B.n462 10.6151
R1404 B.n462 B.n459 10.6151
R1405 B.n459 B.n458 10.6151
R1406 B.n458 B.n455 10.6151
R1407 B.n455 B.n454 10.6151
R1408 B.n454 B.n451 10.6151
R1409 B.n451 B.n450 10.6151
R1410 B.n450 B.n447 10.6151
R1411 B.n447 B.n446 10.6151
R1412 B.n446 B.n443 10.6151
R1413 B.n443 B.n442 10.6151
R1414 B.n442 B.n439 10.6151
R1415 B.n439 B.n438 10.6151
R1416 B.n438 B.n398 10.6151
R1417 B.n566 B.n398 10.6151
R1418 B.n568 B.n567 10.6151
R1419 B.n568 B.n390 10.6151
R1420 B.n578 B.n390 10.6151
R1421 B.n579 B.n578 10.6151
R1422 B.n580 B.n579 10.6151
R1423 B.n580 B.n382 10.6151
R1424 B.n590 B.n382 10.6151
R1425 B.n591 B.n590 10.6151
R1426 B.n592 B.n591 10.6151
R1427 B.n592 B.n374 10.6151
R1428 B.n602 B.n374 10.6151
R1429 B.n603 B.n602 10.6151
R1430 B.n604 B.n603 10.6151
R1431 B.n604 B.n366 10.6151
R1432 B.n614 B.n366 10.6151
R1433 B.n615 B.n614 10.6151
R1434 B.n616 B.n615 10.6151
R1435 B.n616 B.n358 10.6151
R1436 B.n626 B.n358 10.6151
R1437 B.n627 B.n626 10.6151
R1438 B.n628 B.n627 10.6151
R1439 B.n628 B.n350 10.6151
R1440 B.n638 B.n350 10.6151
R1441 B.n639 B.n638 10.6151
R1442 B.n640 B.n639 10.6151
R1443 B.n640 B.n341 10.6151
R1444 B.n650 B.n341 10.6151
R1445 B.n651 B.n650 10.6151
R1446 B.n652 B.n651 10.6151
R1447 B.n652 B.n334 10.6151
R1448 B.n662 B.n334 10.6151
R1449 B.n663 B.n662 10.6151
R1450 B.n664 B.n663 10.6151
R1451 B.n664 B.n326 10.6151
R1452 B.n674 B.n326 10.6151
R1453 B.n675 B.n674 10.6151
R1454 B.n676 B.n675 10.6151
R1455 B.n676 B.n318 10.6151
R1456 B.n686 B.n318 10.6151
R1457 B.n687 B.n686 10.6151
R1458 B.n688 B.n687 10.6151
R1459 B.n688 B.n310 10.6151
R1460 B.n698 B.n310 10.6151
R1461 B.n699 B.n698 10.6151
R1462 B.n700 B.n699 10.6151
R1463 B.n700 B.n303 10.6151
R1464 B.n711 B.n303 10.6151
R1465 B.n712 B.n711 10.6151
R1466 B.n713 B.n712 10.6151
R1467 B.n713 B.n295 10.6151
R1468 B.n723 B.n295 10.6151
R1469 B.n724 B.n723 10.6151
R1470 B.n725 B.n724 10.6151
R1471 B.n725 B.n287 10.6151
R1472 B.n735 B.n287 10.6151
R1473 B.n736 B.n735 10.6151
R1474 B.n738 B.n736 10.6151
R1475 B.n738 B.n737 10.6151
R1476 B.n737 B.n279 10.6151
R1477 B.n749 B.n279 10.6151
R1478 B.n750 B.n749 10.6151
R1479 B.n751 B.n750 10.6151
R1480 B.n752 B.n751 10.6151
R1481 B.n753 B.n752 10.6151
R1482 B.n756 B.n753 10.6151
R1483 B.n757 B.n756 10.6151
R1484 B.n758 B.n757 10.6151
R1485 B.n759 B.n758 10.6151
R1486 B.n761 B.n759 10.6151
R1487 B.n762 B.n761 10.6151
R1488 B.n763 B.n762 10.6151
R1489 B.n764 B.n763 10.6151
R1490 B.n766 B.n764 10.6151
R1491 B.n767 B.n766 10.6151
R1492 B.n768 B.n767 10.6151
R1493 B.n769 B.n768 10.6151
R1494 B.n771 B.n769 10.6151
R1495 B.n772 B.n771 10.6151
R1496 B.n773 B.n772 10.6151
R1497 B.n774 B.n773 10.6151
R1498 B.n776 B.n774 10.6151
R1499 B.n777 B.n776 10.6151
R1500 B.n778 B.n777 10.6151
R1501 B.n779 B.n778 10.6151
R1502 B.n781 B.n779 10.6151
R1503 B.n782 B.n781 10.6151
R1504 B.n783 B.n782 10.6151
R1505 B.n784 B.n783 10.6151
R1506 B.n786 B.n784 10.6151
R1507 B.n787 B.n786 10.6151
R1508 B.n788 B.n787 10.6151
R1509 B.n789 B.n788 10.6151
R1510 B.n791 B.n789 10.6151
R1511 B.n792 B.n791 10.6151
R1512 B.n793 B.n792 10.6151
R1513 B.n794 B.n793 10.6151
R1514 B.n796 B.n794 10.6151
R1515 B.n797 B.n796 10.6151
R1516 B.n798 B.n797 10.6151
R1517 B.n799 B.n798 10.6151
R1518 B.n801 B.n799 10.6151
R1519 B.n802 B.n801 10.6151
R1520 B.n803 B.n802 10.6151
R1521 B.n804 B.n803 10.6151
R1522 B.n806 B.n804 10.6151
R1523 B.n807 B.n806 10.6151
R1524 B.n808 B.n807 10.6151
R1525 B.n809 B.n808 10.6151
R1526 B.n811 B.n809 10.6151
R1527 B.n812 B.n811 10.6151
R1528 B.n813 B.n812 10.6151
R1529 B.n814 B.n813 10.6151
R1530 B.n816 B.n814 10.6151
R1531 B.n817 B.n816 10.6151
R1532 B.n818 B.n817 10.6151
R1533 B.n819 B.n818 10.6151
R1534 B.n821 B.n819 10.6151
R1535 B.n822 B.n821 10.6151
R1536 B.n823 B.n822 10.6151
R1537 B.n824 B.n823 10.6151
R1538 B.n826 B.n824 10.6151
R1539 B.n827 B.n826 10.6151
R1540 B.n828 B.n827 10.6151
R1541 B.n949 B.n1 10.6151
R1542 B.n949 B.n948 10.6151
R1543 B.n948 B.n947 10.6151
R1544 B.n947 B.n10 10.6151
R1545 B.n941 B.n10 10.6151
R1546 B.n941 B.n940 10.6151
R1547 B.n940 B.n939 10.6151
R1548 B.n939 B.n18 10.6151
R1549 B.n933 B.n18 10.6151
R1550 B.n933 B.n932 10.6151
R1551 B.n932 B.n931 10.6151
R1552 B.n931 B.n25 10.6151
R1553 B.n925 B.n25 10.6151
R1554 B.n925 B.n924 10.6151
R1555 B.n924 B.n923 10.6151
R1556 B.n923 B.n31 10.6151
R1557 B.n917 B.n31 10.6151
R1558 B.n917 B.n916 10.6151
R1559 B.n916 B.n915 10.6151
R1560 B.n915 B.n39 10.6151
R1561 B.n909 B.n39 10.6151
R1562 B.n909 B.n908 10.6151
R1563 B.n908 B.n907 10.6151
R1564 B.n907 B.n46 10.6151
R1565 B.n901 B.n46 10.6151
R1566 B.n901 B.n900 10.6151
R1567 B.n900 B.n899 10.6151
R1568 B.n899 B.n53 10.6151
R1569 B.n893 B.n53 10.6151
R1570 B.n893 B.n892 10.6151
R1571 B.n892 B.n891 10.6151
R1572 B.n891 B.n60 10.6151
R1573 B.n885 B.n60 10.6151
R1574 B.n885 B.n884 10.6151
R1575 B.n884 B.n883 10.6151
R1576 B.n883 B.n67 10.6151
R1577 B.n877 B.n67 10.6151
R1578 B.n877 B.n876 10.6151
R1579 B.n876 B.n875 10.6151
R1580 B.n875 B.n74 10.6151
R1581 B.n869 B.n74 10.6151
R1582 B.n869 B.n868 10.6151
R1583 B.n868 B.n867 10.6151
R1584 B.n867 B.n81 10.6151
R1585 B.n861 B.n81 10.6151
R1586 B.n861 B.n860 10.6151
R1587 B.n860 B.n859 10.6151
R1588 B.n859 B.n88 10.6151
R1589 B.n853 B.n88 10.6151
R1590 B.n853 B.n852 10.6151
R1591 B.n852 B.n851 10.6151
R1592 B.n851 B.n95 10.6151
R1593 B.n845 B.n95 10.6151
R1594 B.n845 B.n844 10.6151
R1595 B.n844 B.n843 10.6151
R1596 B.n843 B.n102 10.6151
R1597 B.n837 B.n102 10.6151
R1598 B.n837 B.n836 10.6151
R1599 B.n836 B.n835 10.6151
R1600 B.n835 B.n109 10.6151
R1601 B.n153 B.n152 10.6151
R1602 B.n156 B.n153 10.6151
R1603 B.n157 B.n156 10.6151
R1604 B.n160 B.n157 10.6151
R1605 B.n161 B.n160 10.6151
R1606 B.n164 B.n161 10.6151
R1607 B.n165 B.n164 10.6151
R1608 B.n168 B.n165 10.6151
R1609 B.n169 B.n168 10.6151
R1610 B.n172 B.n169 10.6151
R1611 B.n173 B.n172 10.6151
R1612 B.n176 B.n173 10.6151
R1613 B.n177 B.n176 10.6151
R1614 B.n180 B.n177 10.6151
R1615 B.n181 B.n180 10.6151
R1616 B.n184 B.n181 10.6151
R1617 B.n185 B.n184 10.6151
R1618 B.n188 B.n185 10.6151
R1619 B.n189 B.n188 10.6151
R1620 B.n192 B.n189 10.6151
R1621 B.n193 B.n192 10.6151
R1622 B.n196 B.n193 10.6151
R1623 B.n197 B.n196 10.6151
R1624 B.n200 B.n197 10.6151
R1625 B.n201 B.n200 10.6151
R1626 B.n204 B.n201 10.6151
R1627 B.n205 B.n204 10.6151
R1628 B.n209 B.n208 10.6151
R1629 B.n212 B.n209 10.6151
R1630 B.n213 B.n212 10.6151
R1631 B.n216 B.n213 10.6151
R1632 B.n217 B.n216 10.6151
R1633 B.n220 B.n217 10.6151
R1634 B.n221 B.n220 10.6151
R1635 B.n224 B.n221 10.6151
R1636 B.n229 B.n226 10.6151
R1637 B.n230 B.n229 10.6151
R1638 B.n233 B.n230 10.6151
R1639 B.n234 B.n233 10.6151
R1640 B.n237 B.n234 10.6151
R1641 B.n238 B.n237 10.6151
R1642 B.n241 B.n238 10.6151
R1643 B.n242 B.n241 10.6151
R1644 B.n245 B.n242 10.6151
R1645 B.n246 B.n245 10.6151
R1646 B.n249 B.n246 10.6151
R1647 B.n250 B.n249 10.6151
R1648 B.n253 B.n250 10.6151
R1649 B.n254 B.n253 10.6151
R1650 B.n257 B.n254 10.6151
R1651 B.n258 B.n257 10.6151
R1652 B.n261 B.n258 10.6151
R1653 B.n262 B.n261 10.6151
R1654 B.n265 B.n262 10.6151
R1655 B.n266 B.n265 10.6151
R1656 B.n269 B.n266 10.6151
R1657 B.n270 B.n269 10.6151
R1658 B.n273 B.n270 10.6151
R1659 B.n274 B.n273 10.6151
R1660 B.n277 B.n274 10.6151
R1661 B.n278 B.n277 10.6151
R1662 B.n829 B.n278 10.6151
R1663 B.n957 B.n0 8.11757
R1664 B.n957 B.n1 8.11757
R1665 B.n507 B.n506 6.5566
R1666 B.n490 B.n436 6.5566
R1667 B.n208 B.n150 6.5566
R1668 B.n225 B.n224 6.5566
R1669 B.n508 B.n507 4.05904
R1670 B.n487 B.n436 4.05904
R1671 B.n205 B.n150 4.05904
R1672 B.n226 B.n225 4.05904
R1673 VN.n83 VN.n43 161.3
R1674 VN.n82 VN.n81 161.3
R1675 VN.n80 VN.n44 161.3
R1676 VN.n79 VN.n78 161.3
R1677 VN.n77 VN.n45 161.3
R1678 VN.n76 VN.n75 161.3
R1679 VN.n74 VN.n73 161.3
R1680 VN.n72 VN.n47 161.3
R1681 VN.n71 VN.n70 161.3
R1682 VN.n69 VN.n48 161.3
R1683 VN.n68 VN.n67 161.3
R1684 VN.n66 VN.n49 161.3
R1685 VN.n65 VN.n64 161.3
R1686 VN.n63 VN.n50 161.3
R1687 VN.n62 VN.n61 161.3
R1688 VN.n60 VN.n51 161.3
R1689 VN.n59 VN.n58 161.3
R1690 VN.n57 VN.n52 161.3
R1691 VN.n56 VN.n55 161.3
R1692 VN.n40 VN.n0 161.3
R1693 VN.n39 VN.n38 161.3
R1694 VN.n37 VN.n1 161.3
R1695 VN.n36 VN.n35 161.3
R1696 VN.n34 VN.n2 161.3
R1697 VN.n33 VN.n32 161.3
R1698 VN.n31 VN.n30 161.3
R1699 VN.n29 VN.n4 161.3
R1700 VN.n28 VN.n27 161.3
R1701 VN.n26 VN.n5 161.3
R1702 VN.n25 VN.n24 161.3
R1703 VN.n23 VN.n6 161.3
R1704 VN.n22 VN.n21 161.3
R1705 VN.n20 VN.n7 161.3
R1706 VN.n19 VN.n18 161.3
R1707 VN.n17 VN.n8 161.3
R1708 VN.n16 VN.n15 161.3
R1709 VN.n14 VN.n9 161.3
R1710 VN.n13 VN.n12 161.3
R1711 VN.n42 VN.n41 106.841
R1712 VN.n85 VN.n84 106.841
R1713 VN.n10 VN.t5 96.6823
R1714 VN.n53 VN.t7 96.6823
R1715 VN.n11 VN.n10 71.2257
R1716 VN.n54 VN.n53 71.2257
R1717 VN.n22 VN.t3 65.1861
R1718 VN.n11 VN.t1 65.1861
R1719 VN.n3 VN.t4 65.1861
R1720 VN.n41 VN.t0 65.1861
R1721 VN.n65 VN.t9 65.1861
R1722 VN.n54 VN.t2 65.1861
R1723 VN.n46 VN.t6 65.1861
R1724 VN.n84 VN.t8 65.1861
R1725 VN VN.n85 50.4072
R1726 VN.n35 VN.n1 46.321
R1727 VN.n78 VN.n44 46.321
R1728 VN.n17 VN.n16 42.4359
R1729 VN.n28 VN.n5 42.4359
R1730 VN.n60 VN.n59 42.4359
R1731 VN.n71 VN.n48 42.4359
R1732 VN.n18 VN.n17 38.5509
R1733 VN.n24 VN.n5 38.5509
R1734 VN.n61 VN.n60 38.5509
R1735 VN.n67 VN.n48 38.5509
R1736 VN.n35 VN.n34 34.6658
R1737 VN.n78 VN.n77 34.6658
R1738 VN.n12 VN.n9 24.4675
R1739 VN.n16 VN.n9 24.4675
R1740 VN.n18 VN.n7 24.4675
R1741 VN.n22 VN.n7 24.4675
R1742 VN.n23 VN.n22 24.4675
R1743 VN.n24 VN.n23 24.4675
R1744 VN.n29 VN.n28 24.4675
R1745 VN.n30 VN.n29 24.4675
R1746 VN.n34 VN.n33 24.4675
R1747 VN.n39 VN.n1 24.4675
R1748 VN.n40 VN.n39 24.4675
R1749 VN.n59 VN.n52 24.4675
R1750 VN.n55 VN.n52 24.4675
R1751 VN.n67 VN.n66 24.4675
R1752 VN.n66 VN.n65 24.4675
R1753 VN.n65 VN.n50 24.4675
R1754 VN.n61 VN.n50 24.4675
R1755 VN.n77 VN.n76 24.4675
R1756 VN.n73 VN.n72 24.4675
R1757 VN.n72 VN.n71 24.4675
R1758 VN.n83 VN.n82 24.4675
R1759 VN.n82 VN.n44 24.4675
R1760 VN.n33 VN.n3 22.5101
R1761 VN.n76 VN.n46 22.5101
R1762 VN.n56 VN.n53 7.24287
R1763 VN.n13 VN.n10 7.24287
R1764 VN.n41 VN.n40 3.91522
R1765 VN.n84 VN.n83 3.91522
R1766 VN.n12 VN.n11 1.95786
R1767 VN.n30 VN.n3 1.95786
R1768 VN.n55 VN.n54 1.95786
R1769 VN.n73 VN.n46 1.95786
R1770 VN.n85 VN.n43 0.278367
R1771 VN.n42 VN.n0 0.278367
R1772 VN.n81 VN.n43 0.189894
R1773 VN.n81 VN.n80 0.189894
R1774 VN.n80 VN.n79 0.189894
R1775 VN.n79 VN.n45 0.189894
R1776 VN.n75 VN.n45 0.189894
R1777 VN.n75 VN.n74 0.189894
R1778 VN.n74 VN.n47 0.189894
R1779 VN.n70 VN.n47 0.189894
R1780 VN.n70 VN.n69 0.189894
R1781 VN.n69 VN.n68 0.189894
R1782 VN.n68 VN.n49 0.189894
R1783 VN.n64 VN.n49 0.189894
R1784 VN.n64 VN.n63 0.189894
R1785 VN.n63 VN.n62 0.189894
R1786 VN.n62 VN.n51 0.189894
R1787 VN.n58 VN.n51 0.189894
R1788 VN.n58 VN.n57 0.189894
R1789 VN.n57 VN.n56 0.189894
R1790 VN.n14 VN.n13 0.189894
R1791 VN.n15 VN.n14 0.189894
R1792 VN.n15 VN.n8 0.189894
R1793 VN.n19 VN.n8 0.189894
R1794 VN.n20 VN.n19 0.189894
R1795 VN.n21 VN.n20 0.189894
R1796 VN.n21 VN.n6 0.189894
R1797 VN.n25 VN.n6 0.189894
R1798 VN.n26 VN.n25 0.189894
R1799 VN.n27 VN.n26 0.189894
R1800 VN.n27 VN.n4 0.189894
R1801 VN.n31 VN.n4 0.189894
R1802 VN.n32 VN.n31 0.189894
R1803 VN.n32 VN.n2 0.189894
R1804 VN.n36 VN.n2 0.189894
R1805 VN.n37 VN.n36 0.189894
R1806 VN.n38 VN.n37 0.189894
R1807 VN.n38 VN.n0 0.189894
R1808 VN VN.n42 0.153454
R1809 VTAIL.n168 VTAIL.n134 289.615
R1810 VTAIL.n36 VTAIL.n2 289.615
R1811 VTAIL.n128 VTAIL.n94 289.615
R1812 VTAIL.n84 VTAIL.n50 289.615
R1813 VTAIL.n146 VTAIL.n145 185
R1814 VTAIL.n151 VTAIL.n150 185
R1815 VTAIL.n153 VTAIL.n152 185
R1816 VTAIL.n142 VTAIL.n141 185
R1817 VTAIL.n159 VTAIL.n158 185
R1818 VTAIL.n161 VTAIL.n160 185
R1819 VTAIL.n138 VTAIL.n137 185
R1820 VTAIL.n167 VTAIL.n166 185
R1821 VTAIL.n169 VTAIL.n168 185
R1822 VTAIL.n14 VTAIL.n13 185
R1823 VTAIL.n19 VTAIL.n18 185
R1824 VTAIL.n21 VTAIL.n20 185
R1825 VTAIL.n10 VTAIL.n9 185
R1826 VTAIL.n27 VTAIL.n26 185
R1827 VTAIL.n29 VTAIL.n28 185
R1828 VTAIL.n6 VTAIL.n5 185
R1829 VTAIL.n35 VTAIL.n34 185
R1830 VTAIL.n37 VTAIL.n36 185
R1831 VTAIL.n129 VTAIL.n128 185
R1832 VTAIL.n127 VTAIL.n126 185
R1833 VTAIL.n98 VTAIL.n97 185
R1834 VTAIL.n121 VTAIL.n120 185
R1835 VTAIL.n119 VTAIL.n118 185
R1836 VTAIL.n102 VTAIL.n101 185
R1837 VTAIL.n113 VTAIL.n112 185
R1838 VTAIL.n111 VTAIL.n110 185
R1839 VTAIL.n106 VTAIL.n105 185
R1840 VTAIL.n85 VTAIL.n84 185
R1841 VTAIL.n83 VTAIL.n82 185
R1842 VTAIL.n54 VTAIL.n53 185
R1843 VTAIL.n77 VTAIL.n76 185
R1844 VTAIL.n75 VTAIL.n74 185
R1845 VTAIL.n58 VTAIL.n57 185
R1846 VTAIL.n69 VTAIL.n68 185
R1847 VTAIL.n67 VTAIL.n66 185
R1848 VTAIL.n62 VTAIL.n61 185
R1849 VTAIL.n147 VTAIL.t10 147.659
R1850 VTAIL.n15 VTAIL.t6 147.659
R1851 VTAIL.n107 VTAIL.t2 147.659
R1852 VTAIL.n63 VTAIL.t16 147.659
R1853 VTAIL.n151 VTAIL.n145 104.615
R1854 VTAIL.n152 VTAIL.n151 104.615
R1855 VTAIL.n152 VTAIL.n141 104.615
R1856 VTAIL.n159 VTAIL.n141 104.615
R1857 VTAIL.n160 VTAIL.n159 104.615
R1858 VTAIL.n160 VTAIL.n137 104.615
R1859 VTAIL.n167 VTAIL.n137 104.615
R1860 VTAIL.n168 VTAIL.n167 104.615
R1861 VTAIL.n19 VTAIL.n13 104.615
R1862 VTAIL.n20 VTAIL.n19 104.615
R1863 VTAIL.n20 VTAIL.n9 104.615
R1864 VTAIL.n27 VTAIL.n9 104.615
R1865 VTAIL.n28 VTAIL.n27 104.615
R1866 VTAIL.n28 VTAIL.n5 104.615
R1867 VTAIL.n35 VTAIL.n5 104.615
R1868 VTAIL.n36 VTAIL.n35 104.615
R1869 VTAIL.n128 VTAIL.n127 104.615
R1870 VTAIL.n127 VTAIL.n97 104.615
R1871 VTAIL.n120 VTAIL.n97 104.615
R1872 VTAIL.n120 VTAIL.n119 104.615
R1873 VTAIL.n119 VTAIL.n101 104.615
R1874 VTAIL.n112 VTAIL.n101 104.615
R1875 VTAIL.n112 VTAIL.n111 104.615
R1876 VTAIL.n111 VTAIL.n105 104.615
R1877 VTAIL.n84 VTAIL.n83 104.615
R1878 VTAIL.n83 VTAIL.n53 104.615
R1879 VTAIL.n76 VTAIL.n53 104.615
R1880 VTAIL.n76 VTAIL.n75 104.615
R1881 VTAIL.n75 VTAIL.n57 104.615
R1882 VTAIL.n68 VTAIL.n57 104.615
R1883 VTAIL.n68 VTAIL.n67 104.615
R1884 VTAIL.n67 VTAIL.n61 104.615
R1885 VTAIL.t10 VTAIL.n145 52.3082
R1886 VTAIL.t6 VTAIL.n13 52.3082
R1887 VTAIL.t2 VTAIL.n105 52.3082
R1888 VTAIL.t16 VTAIL.n61 52.3082
R1889 VTAIL.n93 VTAIL.n92 46.3884
R1890 VTAIL.n91 VTAIL.n90 46.3884
R1891 VTAIL.n49 VTAIL.n48 46.3884
R1892 VTAIL.n47 VTAIL.n46 46.3884
R1893 VTAIL.n175 VTAIL.n174 46.3882
R1894 VTAIL.n1 VTAIL.n0 46.3882
R1895 VTAIL.n43 VTAIL.n42 46.3882
R1896 VTAIL.n45 VTAIL.n44 46.3882
R1897 VTAIL.n173 VTAIL.n172 30.052
R1898 VTAIL.n41 VTAIL.n40 30.052
R1899 VTAIL.n133 VTAIL.n132 30.052
R1900 VTAIL.n89 VTAIL.n88 30.052
R1901 VTAIL.n47 VTAIL.n45 23.9272
R1902 VTAIL.n173 VTAIL.n133 21.3065
R1903 VTAIL.n147 VTAIL.n146 15.6677
R1904 VTAIL.n15 VTAIL.n14 15.6677
R1905 VTAIL.n107 VTAIL.n106 15.6677
R1906 VTAIL.n63 VTAIL.n62 15.6677
R1907 VTAIL.n150 VTAIL.n149 12.8005
R1908 VTAIL.n18 VTAIL.n17 12.8005
R1909 VTAIL.n110 VTAIL.n109 12.8005
R1910 VTAIL.n66 VTAIL.n65 12.8005
R1911 VTAIL.n153 VTAIL.n144 12.0247
R1912 VTAIL.n21 VTAIL.n12 12.0247
R1913 VTAIL.n113 VTAIL.n104 12.0247
R1914 VTAIL.n69 VTAIL.n60 12.0247
R1915 VTAIL.n154 VTAIL.n142 11.249
R1916 VTAIL.n22 VTAIL.n10 11.249
R1917 VTAIL.n114 VTAIL.n102 11.249
R1918 VTAIL.n70 VTAIL.n58 11.249
R1919 VTAIL.n158 VTAIL.n157 10.4732
R1920 VTAIL.n26 VTAIL.n25 10.4732
R1921 VTAIL.n118 VTAIL.n117 10.4732
R1922 VTAIL.n74 VTAIL.n73 10.4732
R1923 VTAIL.n161 VTAIL.n140 9.69747
R1924 VTAIL.n29 VTAIL.n8 9.69747
R1925 VTAIL.n121 VTAIL.n100 9.69747
R1926 VTAIL.n77 VTAIL.n56 9.69747
R1927 VTAIL.n172 VTAIL.n171 9.45567
R1928 VTAIL.n40 VTAIL.n39 9.45567
R1929 VTAIL.n132 VTAIL.n131 9.45567
R1930 VTAIL.n88 VTAIL.n87 9.45567
R1931 VTAIL.n171 VTAIL.n170 9.3005
R1932 VTAIL.n165 VTAIL.n164 9.3005
R1933 VTAIL.n163 VTAIL.n162 9.3005
R1934 VTAIL.n140 VTAIL.n139 9.3005
R1935 VTAIL.n157 VTAIL.n156 9.3005
R1936 VTAIL.n155 VTAIL.n154 9.3005
R1937 VTAIL.n144 VTAIL.n143 9.3005
R1938 VTAIL.n149 VTAIL.n148 9.3005
R1939 VTAIL.n136 VTAIL.n135 9.3005
R1940 VTAIL.n39 VTAIL.n38 9.3005
R1941 VTAIL.n33 VTAIL.n32 9.3005
R1942 VTAIL.n31 VTAIL.n30 9.3005
R1943 VTAIL.n8 VTAIL.n7 9.3005
R1944 VTAIL.n25 VTAIL.n24 9.3005
R1945 VTAIL.n23 VTAIL.n22 9.3005
R1946 VTAIL.n12 VTAIL.n11 9.3005
R1947 VTAIL.n17 VTAIL.n16 9.3005
R1948 VTAIL.n4 VTAIL.n3 9.3005
R1949 VTAIL.n131 VTAIL.n130 9.3005
R1950 VTAIL.n96 VTAIL.n95 9.3005
R1951 VTAIL.n125 VTAIL.n124 9.3005
R1952 VTAIL.n123 VTAIL.n122 9.3005
R1953 VTAIL.n100 VTAIL.n99 9.3005
R1954 VTAIL.n117 VTAIL.n116 9.3005
R1955 VTAIL.n115 VTAIL.n114 9.3005
R1956 VTAIL.n104 VTAIL.n103 9.3005
R1957 VTAIL.n109 VTAIL.n108 9.3005
R1958 VTAIL.n87 VTAIL.n86 9.3005
R1959 VTAIL.n52 VTAIL.n51 9.3005
R1960 VTAIL.n81 VTAIL.n80 9.3005
R1961 VTAIL.n79 VTAIL.n78 9.3005
R1962 VTAIL.n56 VTAIL.n55 9.3005
R1963 VTAIL.n73 VTAIL.n72 9.3005
R1964 VTAIL.n71 VTAIL.n70 9.3005
R1965 VTAIL.n60 VTAIL.n59 9.3005
R1966 VTAIL.n65 VTAIL.n64 9.3005
R1967 VTAIL.n162 VTAIL.n138 8.92171
R1968 VTAIL.n30 VTAIL.n6 8.92171
R1969 VTAIL.n122 VTAIL.n98 8.92171
R1970 VTAIL.n78 VTAIL.n54 8.92171
R1971 VTAIL.n166 VTAIL.n165 8.14595
R1972 VTAIL.n34 VTAIL.n33 8.14595
R1973 VTAIL.n126 VTAIL.n125 8.14595
R1974 VTAIL.n82 VTAIL.n81 8.14595
R1975 VTAIL.n169 VTAIL.n136 7.3702
R1976 VTAIL.n172 VTAIL.n134 7.3702
R1977 VTAIL.n37 VTAIL.n4 7.3702
R1978 VTAIL.n40 VTAIL.n2 7.3702
R1979 VTAIL.n132 VTAIL.n94 7.3702
R1980 VTAIL.n129 VTAIL.n96 7.3702
R1981 VTAIL.n88 VTAIL.n50 7.3702
R1982 VTAIL.n85 VTAIL.n52 7.3702
R1983 VTAIL.n170 VTAIL.n169 6.59444
R1984 VTAIL.n170 VTAIL.n134 6.59444
R1985 VTAIL.n38 VTAIL.n37 6.59444
R1986 VTAIL.n38 VTAIL.n2 6.59444
R1987 VTAIL.n130 VTAIL.n94 6.59444
R1988 VTAIL.n130 VTAIL.n129 6.59444
R1989 VTAIL.n86 VTAIL.n50 6.59444
R1990 VTAIL.n86 VTAIL.n85 6.59444
R1991 VTAIL.n166 VTAIL.n136 5.81868
R1992 VTAIL.n34 VTAIL.n4 5.81868
R1993 VTAIL.n126 VTAIL.n96 5.81868
R1994 VTAIL.n82 VTAIL.n52 5.81868
R1995 VTAIL.n165 VTAIL.n138 5.04292
R1996 VTAIL.n33 VTAIL.n6 5.04292
R1997 VTAIL.n125 VTAIL.n98 5.04292
R1998 VTAIL.n81 VTAIL.n54 5.04292
R1999 VTAIL.n108 VTAIL.n107 4.38565
R2000 VTAIL.n64 VTAIL.n63 4.38565
R2001 VTAIL.n148 VTAIL.n147 4.38565
R2002 VTAIL.n16 VTAIL.n15 4.38565
R2003 VTAIL.n162 VTAIL.n161 4.26717
R2004 VTAIL.n30 VTAIL.n29 4.26717
R2005 VTAIL.n122 VTAIL.n121 4.26717
R2006 VTAIL.n78 VTAIL.n77 4.26717
R2007 VTAIL.n158 VTAIL.n140 3.49141
R2008 VTAIL.n26 VTAIL.n8 3.49141
R2009 VTAIL.n118 VTAIL.n100 3.49141
R2010 VTAIL.n74 VTAIL.n56 3.49141
R2011 VTAIL.n157 VTAIL.n142 2.71565
R2012 VTAIL.n25 VTAIL.n10 2.71565
R2013 VTAIL.n117 VTAIL.n102 2.71565
R2014 VTAIL.n73 VTAIL.n58 2.71565
R2015 VTAIL.n174 VTAIL.t13 2.70173
R2016 VTAIL.n174 VTAIL.t8 2.70173
R2017 VTAIL.n0 VTAIL.t17 2.70173
R2018 VTAIL.n0 VTAIL.t11 2.70173
R2019 VTAIL.n42 VTAIL.t19 2.70173
R2020 VTAIL.n42 VTAIL.t1 2.70173
R2021 VTAIL.n44 VTAIL.t18 2.70173
R2022 VTAIL.n44 VTAIL.t7 2.70173
R2023 VTAIL.n92 VTAIL.t4 2.70173
R2024 VTAIL.n92 VTAIL.t3 2.70173
R2025 VTAIL.n90 VTAIL.t0 2.70173
R2026 VTAIL.n90 VTAIL.t5 2.70173
R2027 VTAIL.n48 VTAIL.t9 2.70173
R2028 VTAIL.n48 VTAIL.t12 2.70173
R2029 VTAIL.n46 VTAIL.t14 2.70173
R2030 VTAIL.n46 VTAIL.t15 2.70173
R2031 VTAIL.n49 VTAIL.n47 2.62119
R2032 VTAIL.n89 VTAIL.n49 2.62119
R2033 VTAIL.n93 VTAIL.n91 2.62119
R2034 VTAIL.n133 VTAIL.n93 2.62119
R2035 VTAIL.n45 VTAIL.n43 2.62119
R2036 VTAIL.n43 VTAIL.n41 2.62119
R2037 VTAIL.n175 VTAIL.n173 2.62119
R2038 VTAIL VTAIL.n1 2.02421
R2039 VTAIL.n154 VTAIL.n153 1.93989
R2040 VTAIL.n22 VTAIL.n21 1.93989
R2041 VTAIL.n114 VTAIL.n113 1.93989
R2042 VTAIL.n70 VTAIL.n69 1.93989
R2043 VTAIL.n91 VTAIL.n89 1.78067
R2044 VTAIL.n41 VTAIL.n1 1.78067
R2045 VTAIL.n150 VTAIL.n144 1.16414
R2046 VTAIL.n18 VTAIL.n12 1.16414
R2047 VTAIL.n110 VTAIL.n104 1.16414
R2048 VTAIL.n66 VTAIL.n60 1.16414
R2049 VTAIL VTAIL.n175 0.597483
R2050 VTAIL.n149 VTAIL.n146 0.388379
R2051 VTAIL.n17 VTAIL.n14 0.388379
R2052 VTAIL.n109 VTAIL.n106 0.388379
R2053 VTAIL.n65 VTAIL.n62 0.388379
R2054 VTAIL.n148 VTAIL.n143 0.155672
R2055 VTAIL.n155 VTAIL.n143 0.155672
R2056 VTAIL.n156 VTAIL.n155 0.155672
R2057 VTAIL.n156 VTAIL.n139 0.155672
R2058 VTAIL.n163 VTAIL.n139 0.155672
R2059 VTAIL.n164 VTAIL.n163 0.155672
R2060 VTAIL.n164 VTAIL.n135 0.155672
R2061 VTAIL.n171 VTAIL.n135 0.155672
R2062 VTAIL.n16 VTAIL.n11 0.155672
R2063 VTAIL.n23 VTAIL.n11 0.155672
R2064 VTAIL.n24 VTAIL.n23 0.155672
R2065 VTAIL.n24 VTAIL.n7 0.155672
R2066 VTAIL.n31 VTAIL.n7 0.155672
R2067 VTAIL.n32 VTAIL.n31 0.155672
R2068 VTAIL.n32 VTAIL.n3 0.155672
R2069 VTAIL.n39 VTAIL.n3 0.155672
R2070 VTAIL.n131 VTAIL.n95 0.155672
R2071 VTAIL.n124 VTAIL.n95 0.155672
R2072 VTAIL.n124 VTAIL.n123 0.155672
R2073 VTAIL.n123 VTAIL.n99 0.155672
R2074 VTAIL.n116 VTAIL.n99 0.155672
R2075 VTAIL.n116 VTAIL.n115 0.155672
R2076 VTAIL.n115 VTAIL.n103 0.155672
R2077 VTAIL.n108 VTAIL.n103 0.155672
R2078 VTAIL.n87 VTAIL.n51 0.155672
R2079 VTAIL.n80 VTAIL.n51 0.155672
R2080 VTAIL.n80 VTAIL.n79 0.155672
R2081 VTAIL.n79 VTAIL.n55 0.155672
R2082 VTAIL.n72 VTAIL.n55 0.155672
R2083 VTAIL.n72 VTAIL.n71 0.155672
R2084 VTAIL.n71 VTAIL.n59 0.155672
R2085 VTAIL.n64 VTAIL.n59 0.155672
R2086 VDD2.n77 VDD2.n43 289.615
R2087 VDD2.n34 VDD2.n0 289.615
R2088 VDD2.n78 VDD2.n77 185
R2089 VDD2.n76 VDD2.n75 185
R2090 VDD2.n47 VDD2.n46 185
R2091 VDD2.n70 VDD2.n69 185
R2092 VDD2.n68 VDD2.n67 185
R2093 VDD2.n51 VDD2.n50 185
R2094 VDD2.n62 VDD2.n61 185
R2095 VDD2.n60 VDD2.n59 185
R2096 VDD2.n55 VDD2.n54 185
R2097 VDD2.n12 VDD2.n11 185
R2098 VDD2.n17 VDD2.n16 185
R2099 VDD2.n19 VDD2.n18 185
R2100 VDD2.n8 VDD2.n7 185
R2101 VDD2.n25 VDD2.n24 185
R2102 VDD2.n27 VDD2.n26 185
R2103 VDD2.n4 VDD2.n3 185
R2104 VDD2.n33 VDD2.n32 185
R2105 VDD2.n35 VDD2.n34 185
R2106 VDD2.n56 VDD2.t1 147.659
R2107 VDD2.n13 VDD2.t4 147.659
R2108 VDD2.n77 VDD2.n76 104.615
R2109 VDD2.n76 VDD2.n46 104.615
R2110 VDD2.n69 VDD2.n46 104.615
R2111 VDD2.n69 VDD2.n68 104.615
R2112 VDD2.n68 VDD2.n50 104.615
R2113 VDD2.n61 VDD2.n50 104.615
R2114 VDD2.n61 VDD2.n60 104.615
R2115 VDD2.n60 VDD2.n54 104.615
R2116 VDD2.n17 VDD2.n11 104.615
R2117 VDD2.n18 VDD2.n17 104.615
R2118 VDD2.n18 VDD2.n7 104.615
R2119 VDD2.n25 VDD2.n7 104.615
R2120 VDD2.n26 VDD2.n25 104.615
R2121 VDD2.n26 VDD2.n3 104.615
R2122 VDD2.n33 VDD2.n3 104.615
R2123 VDD2.n34 VDD2.n33 104.615
R2124 VDD2.n42 VDD2.n41 64.9772
R2125 VDD2 VDD2.n85 64.9743
R2126 VDD2.n84 VDD2.n83 63.0672
R2127 VDD2.n40 VDD2.n39 63.067
R2128 VDD2.t1 VDD2.n54 52.3082
R2129 VDD2.t4 VDD2.n11 52.3082
R2130 VDD2.n40 VDD2.n38 49.3515
R2131 VDD2.n82 VDD2.n81 46.7308
R2132 VDD2.n82 VDD2.n42 42.4825
R2133 VDD2.n56 VDD2.n55 15.6677
R2134 VDD2.n13 VDD2.n12 15.6677
R2135 VDD2.n59 VDD2.n58 12.8005
R2136 VDD2.n16 VDD2.n15 12.8005
R2137 VDD2.n62 VDD2.n53 12.0247
R2138 VDD2.n19 VDD2.n10 12.0247
R2139 VDD2.n63 VDD2.n51 11.249
R2140 VDD2.n20 VDD2.n8 11.249
R2141 VDD2.n67 VDD2.n66 10.4732
R2142 VDD2.n24 VDD2.n23 10.4732
R2143 VDD2.n70 VDD2.n49 9.69747
R2144 VDD2.n27 VDD2.n6 9.69747
R2145 VDD2.n81 VDD2.n80 9.45567
R2146 VDD2.n38 VDD2.n37 9.45567
R2147 VDD2.n80 VDD2.n79 9.3005
R2148 VDD2.n45 VDD2.n44 9.3005
R2149 VDD2.n74 VDD2.n73 9.3005
R2150 VDD2.n72 VDD2.n71 9.3005
R2151 VDD2.n49 VDD2.n48 9.3005
R2152 VDD2.n66 VDD2.n65 9.3005
R2153 VDD2.n64 VDD2.n63 9.3005
R2154 VDD2.n53 VDD2.n52 9.3005
R2155 VDD2.n58 VDD2.n57 9.3005
R2156 VDD2.n37 VDD2.n36 9.3005
R2157 VDD2.n31 VDD2.n30 9.3005
R2158 VDD2.n29 VDD2.n28 9.3005
R2159 VDD2.n6 VDD2.n5 9.3005
R2160 VDD2.n23 VDD2.n22 9.3005
R2161 VDD2.n21 VDD2.n20 9.3005
R2162 VDD2.n10 VDD2.n9 9.3005
R2163 VDD2.n15 VDD2.n14 9.3005
R2164 VDD2.n2 VDD2.n1 9.3005
R2165 VDD2.n71 VDD2.n47 8.92171
R2166 VDD2.n28 VDD2.n4 8.92171
R2167 VDD2.n75 VDD2.n74 8.14595
R2168 VDD2.n32 VDD2.n31 8.14595
R2169 VDD2.n81 VDD2.n43 7.3702
R2170 VDD2.n78 VDD2.n45 7.3702
R2171 VDD2.n35 VDD2.n2 7.3702
R2172 VDD2.n38 VDD2.n0 7.3702
R2173 VDD2.n79 VDD2.n43 6.59444
R2174 VDD2.n79 VDD2.n78 6.59444
R2175 VDD2.n36 VDD2.n35 6.59444
R2176 VDD2.n36 VDD2.n0 6.59444
R2177 VDD2.n75 VDD2.n45 5.81868
R2178 VDD2.n32 VDD2.n2 5.81868
R2179 VDD2.n74 VDD2.n47 5.04292
R2180 VDD2.n31 VDD2.n4 5.04292
R2181 VDD2.n57 VDD2.n56 4.38565
R2182 VDD2.n14 VDD2.n13 4.38565
R2183 VDD2.n71 VDD2.n70 4.26717
R2184 VDD2.n28 VDD2.n27 4.26717
R2185 VDD2.n67 VDD2.n49 3.49141
R2186 VDD2.n24 VDD2.n6 3.49141
R2187 VDD2.n66 VDD2.n51 2.71565
R2188 VDD2.n23 VDD2.n8 2.71565
R2189 VDD2.n85 VDD2.t7 2.70173
R2190 VDD2.n85 VDD2.t2 2.70173
R2191 VDD2.n83 VDD2.t3 2.70173
R2192 VDD2.n83 VDD2.t0 2.70173
R2193 VDD2.n41 VDD2.t5 2.70173
R2194 VDD2.n41 VDD2.t9 2.70173
R2195 VDD2.n39 VDD2.t8 2.70173
R2196 VDD2.n39 VDD2.t6 2.70173
R2197 VDD2.n84 VDD2.n82 2.62119
R2198 VDD2.n63 VDD2.n62 1.93989
R2199 VDD2.n20 VDD2.n19 1.93989
R2200 VDD2.n59 VDD2.n53 1.16414
R2201 VDD2.n16 VDD2.n10 1.16414
R2202 VDD2 VDD2.n84 0.713862
R2203 VDD2.n42 VDD2.n40 0.600326
R2204 VDD2.n58 VDD2.n55 0.388379
R2205 VDD2.n15 VDD2.n12 0.388379
R2206 VDD2.n80 VDD2.n44 0.155672
R2207 VDD2.n73 VDD2.n44 0.155672
R2208 VDD2.n73 VDD2.n72 0.155672
R2209 VDD2.n72 VDD2.n48 0.155672
R2210 VDD2.n65 VDD2.n48 0.155672
R2211 VDD2.n65 VDD2.n64 0.155672
R2212 VDD2.n64 VDD2.n52 0.155672
R2213 VDD2.n57 VDD2.n52 0.155672
R2214 VDD2.n14 VDD2.n9 0.155672
R2215 VDD2.n21 VDD2.n9 0.155672
R2216 VDD2.n22 VDD2.n21 0.155672
R2217 VDD2.n22 VDD2.n5 0.155672
R2218 VDD2.n29 VDD2.n5 0.155672
R2219 VDD2.n30 VDD2.n29 0.155672
R2220 VDD2.n30 VDD2.n1 0.155672
R2221 VDD2.n37 VDD2.n1 0.155672
R2222 VP.n27 VP.n26 161.3
R2223 VP.n28 VP.n23 161.3
R2224 VP.n30 VP.n29 161.3
R2225 VP.n31 VP.n22 161.3
R2226 VP.n33 VP.n32 161.3
R2227 VP.n34 VP.n21 161.3
R2228 VP.n36 VP.n35 161.3
R2229 VP.n37 VP.n20 161.3
R2230 VP.n39 VP.n38 161.3
R2231 VP.n40 VP.n19 161.3
R2232 VP.n42 VP.n41 161.3
R2233 VP.n43 VP.n18 161.3
R2234 VP.n45 VP.n44 161.3
R2235 VP.n47 VP.n46 161.3
R2236 VP.n48 VP.n16 161.3
R2237 VP.n50 VP.n49 161.3
R2238 VP.n51 VP.n15 161.3
R2239 VP.n53 VP.n52 161.3
R2240 VP.n54 VP.n14 161.3
R2241 VP.n96 VP.n0 161.3
R2242 VP.n95 VP.n94 161.3
R2243 VP.n93 VP.n1 161.3
R2244 VP.n92 VP.n91 161.3
R2245 VP.n90 VP.n2 161.3
R2246 VP.n89 VP.n88 161.3
R2247 VP.n87 VP.n86 161.3
R2248 VP.n85 VP.n4 161.3
R2249 VP.n84 VP.n83 161.3
R2250 VP.n82 VP.n5 161.3
R2251 VP.n81 VP.n80 161.3
R2252 VP.n79 VP.n6 161.3
R2253 VP.n78 VP.n77 161.3
R2254 VP.n76 VP.n7 161.3
R2255 VP.n75 VP.n74 161.3
R2256 VP.n73 VP.n8 161.3
R2257 VP.n72 VP.n71 161.3
R2258 VP.n70 VP.n9 161.3
R2259 VP.n69 VP.n68 161.3
R2260 VP.n66 VP.n10 161.3
R2261 VP.n65 VP.n64 161.3
R2262 VP.n63 VP.n11 161.3
R2263 VP.n62 VP.n61 161.3
R2264 VP.n60 VP.n12 161.3
R2265 VP.n59 VP.n58 161.3
R2266 VP.n57 VP.n13 106.841
R2267 VP.n98 VP.n97 106.841
R2268 VP.n56 VP.n55 106.841
R2269 VP.n24 VP.t3 96.6823
R2270 VP.n25 VP.n24 71.2257
R2271 VP.n78 VP.t7 65.1861
R2272 VP.n13 VP.t2 65.1861
R2273 VP.n67 VP.t6 65.1861
R2274 VP.n3 VP.t9 65.1861
R2275 VP.n97 VP.t1 65.1861
R2276 VP.n36 VP.t5 65.1861
R2277 VP.n55 VP.t4 65.1861
R2278 VP.n17 VP.t0 65.1861
R2279 VP.n25 VP.t8 65.1861
R2280 VP.n57 VP.n56 50.1284
R2281 VP.n61 VP.n11 46.321
R2282 VP.n91 VP.n1 46.321
R2283 VP.n49 VP.n15 46.321
R2284 VP.n73 VP.n72 42.4359
R2285 VP.n84 VP.n5 42.4359
R2286 VP.n42 VP.n19 42.4359
R2287 VP.n31 VP.n30 42.4359
R2288 VP.n74 VP.n73 38.5509
R2289 VP.n80 VP.n5 38.5509
R2290 VP.n38 VP.n19 38.5509
R2291 VP.n32 VP.n31 38.5509
R2292 VP.n65 VP.n11 34.6658
R2293 VP.n91 VP.n90 34.6658
R2294 VP.n49 VP.n48 34.6658
R2295 VP.n60 VP.n59 24.4675
R2296 VP.n61 VP.n60 24.4675
R2297 VP.n66 VP.n65 24.4675
R2298 VP.n68 VP.n9 24.4675
R2299 VP.n72 VP.n9 24.4675
R2300 VP.n74 VP.n7 24.4675
R2301 VP.n78 VP.n7 24.4675
R2302 VP.n79 VP.n78 24.4675
R2303 VP.n80 VP.n79 24.4675
R2304 VP.n85 VP.n84 24.4675
R2305 VP.n86 VP.n85 24.4675
R2306 VP.n90 VP.n89 24.4675
R2307 VP.n95 VP.n1 24.4675
R2308 VP.n96 VP.n95 24.4675
R2309 VP.n53 VP.n15 24.4675
R2310 VP.n54 VP.n53 24.4675
R2311 VP.n43 VP.n42 24.4675
R2312 VP.n44 VP.n43 24.4675
R2313 VP.n48 VP.n47 24.4675
R2314 VP.n32 VP.n21 24.4675
R2315 VP.n36 VP.n21 24.4675
R2316 VP.n37 VP.n36 24.4675
R2317 VP.n38 VP.n37 24.4675
R2318 VP.n26 VP.n23 24.4675
R2319 VP.n30 VP.n23 24.4675
R2320 VP.n67 VP.n66 22.5101
R2321 VP.n89 VP.n3 22.5101
R2322 VP.n47 VP.n17 22.5101
R2323 VP.n27 VP.n24 7.24287
R2324 VP.n59 VP.n13 3.91522
R2325 VP.n97 VP.n96 3.91522
R2326 VP.n55 VP.n54 3.91522
R2327 VP.n68 VP.n67 1.95786
R2328 VP.n86 VP.n3 1.95786
R2329 VP.n44 VP.n17 1.95786
R2330 VP.n26 VP.n25 1.95786
R2331 VP.n56 VP.n14 0.278367
R2332 VP.n58 VP.n57 0.278367
R2333 VP.n98 VP.n0 0.278367
R2334 VP.n28 VP.n27 0.189894
R2335 VP.n29 VP.n28 0.189894
R2336 VP.n29 VP.n22 0.189894
R2337 VP.n33 VP.n22 0.189894
R2338 VP.n34 VP.n33 0.189894
R2339 VP.n35 VP.n34 0.189894
R2340 VP.n35 VP.n20 0.189894
R2341 VP.n39 VP.n20 0.189894
R2342 VP.n40 VP.n39 0.189894
R2343 VP.n41 VP.n40 0.189894
R2344 VP.n41 VP.n18 0.189894
R2345 VP.n45 VP.n18 0.189894
R2346 VP.n46 VP.n45 0.189894
R2347 VP.n46 VP.n16 0.189894
R2348 VP.n50 VP.n16 0.189894
R2349 VP.n51 VP.n50 0.189894
R2350 VP.n52 VP.n51 0.189894
R2351 VP.n52 VP.n14 0.189894
R2352 VP.n58 VP.n12 0.189894
R2353 VP.n62 VP.n12 0.189894
R2354 VP.n63 VP.n62 0.189894
R2355 VP.n64 VP.n63 0.189894
R2356 VP.n64 VP.n10 0.189894
R2357 VP.n69 VP.n10 0.189894
R2358 VP.n70 VP.n69 0.189894
R2359 VP.n71 VP.n70 0.189894
R2360 VP.n71 VP.n8 0.189894
R2361 VP.n75 VP.n8 0.189894
R2362 VP.n76 VP.n75 0.189894
R2363 VP.n77 VP.n76 0.189894
R2364 VP.n77 VP.n6 0.189894
R2365 VP.n81 VP.n6 0.189894
R2366 VP.n82 VP.n81 0.189894
R2367 VP.n83 VP.n82 0.189894
R2368 VP.n83 VP.n4 0.189894
R2369 VP.n87 VP.n4 0.189894
R2370 VP.n88 VP.n87 0.189894
R2371 VP.n88 VP.n2 0.189894
R2372 VP.n92 VP.n2 0.189894
R2373 VP.n93 VP.n92 0.189894
R2374 VP.n94 VP.n93 0.189894
R2375 VP.n94 VP.n0 0.189894
R2376 VP VP.n98 0.153454
R2377 VDD1.n34 VDD1.n0 289.615
R2378 VDD1.n75 VDD1.n41 289.615
R2379 VDD1.n35 VDD1.n34 185
R2380 VDD1.n33 VDD1.n32 185
R2381 VDD1.n4 VDD1.n3 185
R2382 VDD1.n27 VDD1.n26 185
R2383 VDD1.n25 VDD1.n24 185
R2384 VDD1.n8 VDD1.n7 185
R2385 VDD1.n19 VDD1.n18 185
R2386 VDD1.n17 VDD1.n16 185
R2387 VDD1.n12 VDD1.n11 185
R2388 VDD1.n53 VDD1.n52 185
R2389 VDD1.n58 VDD1.n57 185
R2390 VDD1.n60 VDD1.n59 185
R2391 VDD1.n49 VDD1.n48 185
R2392 VDD1.n66 VDD1.n65 185
R2393 VDD1.n68 VDD1.n67 185
R2394 VDD1.n45 VDD1.n44 185
R2395 VDD1.n74 VDD1.n73 185
R2396 VDD1.n76 VDD1.n75 185
R2397 VDD1.n13 VDD1.t6 147.659
R2398 VDD1.n54 VDD1.t7 147.659
R2399 VDD1.n34 VDD1.n33 104.615
R2400 VDD1.n33 VDD1.n3 104.615
R2401 VDD1.n26 VDD1.n3 104.615
R2402 VDD1.n26 VDD1.n25 104.615
R2403 VDD1.n25 VDD1.n7 104.615
R2404 VDD1.n18 VDD1.n7 104.615
R2405 VDD1.n18 VDD1.n17 104.615
R2406 VDD1.n17 VDD1.n11 104.615
R2407 VDD1.n58 VDD1.n52 104.615
R2408 VDD1.n59 VDD1.n58 104.615
R2409 VDD1.n59 VDD1.n48 104.615
R2410 VDD1.n66 VDD1.n48 104.615
R2411 VDD1.n67 VDD1.n66 104.615
R2412 VDD1.n67 VDD1.n44 104.615
R2413 VDD1.n74 VDD1.n44 104.615
R2414 VDD1.n75 VDD1.n74 104.615
R2415 VDD1.n83 VDD1.n82 64.9772
R2416 VDD1.n40 VDD1.n39 63.0672
R2417 VDD1.n85 VDD1.n84 63.067
R2418 VDD1.n81 VDD1.n80 63.067
R2419 VDD1.t6 VDD1.n11 52.3082
R2420 VDD1.t7 VDD1.n52 52.3082
R2421 VDD1.n40 VDD1.n38 49.3515
R2422 VDD1.n81 VDD1.n79 49.3515
R2423 VDD1.n85 VDD1.n83 44.3759
R2424 VDD1.n13 VDD1.n12 15.6677
R2425 VDD1.n54 VDD1.n53 15.6677
R2426 VDD1.n16 VDD1.n15 12.8005
R2427 VDD1.n57 VDD1.n56 12.8005
R2428 VDD1.n19 VDD1.n10 12.0247
R2429 VDD1.n60 VDD1.n51 12.0247
R2430 VDD1.n20 VDD1.n8 11.249
R2431 VDD1.n61 VDD1.n49 11.249
R2432 VDD1.n24 VDD1.n23 10.4732
R2433 VDD1.n65 VDD1.n64 10.4732
R2434 VDD1.n27 VDD1.n6 9.69747
R2435 VDD1.n68 VDD1.n47 9.69747
R2436 VDD1.n38 VDD1.n37 9.45567
R2437 VDD1.n79 VDD1.n78 9.45567
R2438 VDD1.n37 VDD1.n36 9.3005
R2439 VDD1.n2 VDD1.n1 9.3005
R2440 VDD1.n31 VDD1.n30 9.3005
R2441 VDD1.n29 VDD1.n28 9.3005
R2442 VDD1.n6 VDD1.n5 9.3005
R2443 VDD1.n23 VDD1.n22 9.3005
R2444 VDD1.n21 VDD1.n20 9.3005
R2445 VDD1.n10 VDD1.n9 9.3005
R2446 VDD1.n15 VDD1.n14 9.3005
R2447 VDD1.n78 VDD1.n77 9.3005
R2448 VDD1.n72 VDD1.n71 9.3005
R2449 VDD1.n70 VDD1.n69 9.3005
R2450 VDD1.n47 VDD1.n46 9.3005
R2451 VDD1.n64 VDD1.n63 9.3005
R2452 VDD1.n62 VDD1.n61 9.3005
R2453 VDD1.n51 VDD1.n50 9.3005
R2454 VDD1.n56 VDD1.n55 9.3005
R2455 VDD1.n43 VDD1.n42 9.3005
R2456 VDD1.n28 VDD1.n4 8.92171
R2457 VDD1.n69 VDD1.n45 8.92171
R2458 VDD1.n32 VDD1.n31 8.14595
R2459 VDD1.n73 VDD1.n72 8.14595
R2460 VDD1.n38 VDD1.n0 7.3702
R2461 VDD1.n35 VDD1.n2 7.3702
R2462 VDD1.n76 VDD1.n43 7.3702
R2463 VDD1.n79 VDD1.n41 7.3702
R2464 VDD1.n36 VDD1.n0 6.59444
R2465 VDD1.n36 VDD1.n35 6.59444
R2466 VDD1.n77 VDD1.n76 6.59444
R2467 VDD1.n77 VDD1.n41 6.59444
R2468 VDD1.n32 VDD1.n2 5.81868
R2469 VDD1.n73 VDD1.n43 5.81868
R2470 VDD1.n31 VDD1.n4 5.04292
R2471 VDD1.n72 VDD1.n45 5.04292
R2472 VDD1.n14 VDD1.n13 4.38565
R2473 VDD1.n55 VDD1.n54 4.38565
R2474 VDD1.n28 VDD1.n27 4.26717
R2475 VDD1.n69 VDD1.n68 4.26717
R2476 VDD1.n24 VDD1.n6 3.49141
R2477 VDD1.n65 VDD1.n47 3.49141
R2478 VDD1.n23 VDD1.n8 2.71565
R2479 VDD1.n64 VDD1.n49 2.71565
R2480 VDD1.n84 VDD1.t9 2.70173
R2481 VDD1.n84 VDD1.t5 2.70173
R2482 VDD1.n39 VDD1.t1 2.70173
R2483 VDD1.n39 VDD1.t4 2.70173
R2484 VDD1.n82 VDD1.t0 2.70173
R2485 VDD1.n82 VDD1.t8 2.70173
R2486 VDD1.n80 VDD1.t3 2.70173
R2487 VDD1.n80 VDD1.t2 2.70173
R2488 VDD1.n20 VDD1.n19 1.93989
R2489 VDD1.n61 VDD1.n60 1.93989
R2490 VDD1 VDD1.n85 1.90783
R2491 VDD1.n16 VDD1.n10 1.16414
R2492 VDD1.n57 VDD1.n51 1.16414
R2493 VDD1 VDD1.n40 0.713862
R2494 VDD1.n83 VDD1.n81 0.600326
R2495 VDD1.n15 VDD1.n12 0.388379
R2496 VDD1.n56 VDD1.n53 0.388379
R2497 VDD1.n37 VDD1.n1 0.155672
R2498 VDD1.n30 VDD1.n1 0.155672
R2499 VDD1.n30 VDD1.n29 0.155672
R2500 VDD1.n29 VDD1.n5 0.155672
R2501 VDD1.n22 VDD1.n5 0.155672
R2502 VDD1.n22 VDD1.n21 0.155672
R2503 VDD1.n21 VDD1.n9 0.155672
R2504 VDD1.n14 VDD1.n9 0.155672
R2505 VDD1.n55 VDD1.n50 0.155672
R2506 VDD1.n62 VDD1.n50 0.155672
R2507 VDD1.n63 VDD1.n62 0.155672
R2508 VDD1.n63 VDD1.n46 0.155672
R2509 VDD1.n70 VDD1.n46 0.155672
R2510 VDD1.n71 VDD1.n70 0.155672
R2511 VDD1.n71 VDD1.n42 0.155672
R2512 VDD1.n78 VDD1.n42 0.155672
C0 VN VP 7.69702f
C1 VTAIL VP 7.69262f
C2 VDD1 VDD2 2.2434f
C3 VDD2 VN 6.77677f
C4 VDD2 VTAIL 8.36194f
C5 VDD1 VN 0.153313f
C6 VDD1 VTAIL 8.309099f
C7 VDD2 VP 0.59695f
C8 VN VTAIL 7.6784f
C9 VDD1 VP 7.21735f
C10 VDD2 B 6.560553f
C11 VDD1 B 6.490026f
C12 VTAIL B 6.418513f
C13 VN B 18.309532f
C14 VP B 16.8836f
C15 VDD1.n0 B 0.035962f
C16 VDD1.n1 B 0.025959f
C17 VDD1.n2 B 0.013949f
C18 VDD1.n3 B 0.03297f
C19 VDD1.n4 B 0.01477f
C20 VDD1.n5 B 0.025959f
C21 VDD1.n6 B 0.013949f
C22 VDD1.n7 B 0.03297f
C23 VDD1.n8 B 0.01477f
C24 VDD1.n9 B 0.025959f
C25 VDD1.n10 B 0.013949f
C26 VDD1.n11 B 0.024728f
C27 VDD1.n12 B 0.019476f
C28 VDD1.t6 B 0.053721f
C29 VDD1.n13 B 0.119471f
C30 VDD1.n14 B 0.776289f
C31 VDD1.n15 B 0.013949f
C32 VDD1.n16 B 0.01477f
C33 VDD1.n17 B 0.03297f
C34 VDD1.n18 B 0.03297f
C35 VDD1.n19 B 0.01477f
C36 VDD1.n20 B 0.013949f
C37 VDD1.n21 B 0.025959f
C38 VDD1.n22 B 0.025959f
C39 VDD1.n23 B 0.013949f
C40 VDD1.n24 B 0.01477f
C41 VDD1.n25 B 0.03297f
C42 VDD1.n26 B 0.03297f
C43 VDD1.n27 B 0.01477f
C44 VDD1.n28 B 0.013949f
C45 VDD1.n29 B 0.025959f
C46 VDD1.n30 B 0.025959f
C47 VDD1.n31 B 0.013949f
C48 VDD1.n32 B 0.01477f
C49 VDD1.n33 B 0.03297f
C50 VDD1.n34 B 0.070446f
C51 VDD1.n35 B 0.01477f
C52 VDD1.n36 B 0.013949f
C53 VDD1.n37 B 0.056101f
C54 VDD1.n38 B 0.071332f
C55 VDD1.t1 B 0.150362f
C56 VDD1.t4 B 0.150362f
C57 VDD1.n39 B 1.28075f
C58 VDD1.n40 B 0.74768f
C59 VDD1.n41 B 0.035962f
C60 VDD1.n42 B 0.025959f
C61 VDD1.n43 B 0.013949f
C62 VDD1.n44 B 0.03297f
C63 VDD1.n45 B 0.01477f
C64 VDD1.n46 B 0.025959f
C65 VDD1.n47 B 0.013949f
C66 VDD1.n48 B 0.03297f
C67 VDD1.n49 B 0.01477f
C68 VDD1.n50 B 0.025959f
C69 VDD1.n51 B 0.013949f
C70 VDD1.n52 B 0.024728f
C71 VDD1.n53 B 0.019476f
C72 VDD1.t7 B 0.053721f
C73 VDD1.n54 B 0.119471f
C74 VDD1.n55 B 0.776289f
C75 VDD1.n56 B 0.013949f
C76 VDD1.n57 B 0.01477f
C77 VDD1.n58 B 0.03297f
C78 VDD1.n59 B 0.03297f
C79 VDD1.n60 B 0.01477f
C80 VDD1.n61 B 0.013949f
C81 VDD1.n62 B 0.025959f
C82 VDD1.n63 B 0.025959f
C83 VDD1.n64 B 0.013949f
C84 VDD1.n65 B 0.01477f
C85 VDD1.n66 B 0.03297f
C86 VDD1.n67 B 0.03297f
C87 VDD1.n68 B 0.01477f
C88 VDD1.n69 B 0.013949f
C89 VDD1.n70 B 0.025959f
C90 VDD1.n71 B 0.025959f
C91 VDD1.n72 B 0.013949f
C92 VDD1.n73 B 0.01477f
C93 VDD1.n74 B 0.03297f
C94 VDD1.n75 B 0.070446f
C95 VDD1.n76 B 0.01477f
C96 VDD1.n77 B 0.013949f
C97 VDD1.n78 B 0.056101f
C98 VDD1.n79 B 0.071332f
C99 VDD1.t3 B 0.150362f
C100 VDD1.t2 B 0.150362f
C101 VDD1.n80 B 1.28074f
C102 VDD1.n81 B 0.739193f
C103 VDD1.t0 B 0.150362f
C104 VDD1.t8 B 0.150362f
C105 VDD1.n82 B 1.29855f
C106 VDD1.n83 B 2.91113f
C107 VDD1.t9 B 0.150362f
C108 VDD1.t5 B 0.150362f
C109 VDD1.n84 B 1.28074f
C110 VDD1.n85 B 2.97165f
C111 VP.n0 B 0.03019f
C112 VP.t1 B 1.21677f
C113 VP.n1 B 0.043669f
C114 VP.n2 B 0.022899f
C115 VP.t9 B 1.21677f
C116 VP.n3 B 0.445984f
C117 VP.n4 B 0.022899f
C118 VP.n5 B 0.018629f
C119 VP.n6 B 0.022899f
C120 VP.t7 B 1.21677f
C121 VP.n7 B 0.042677f
C122 VP.n8 B 0.022899f
C123 VP.n9 B 0.042677f
C124 VP.n10 B 0.022899f
C125 VP.t6 B 1.21677f
C126 VP.n11 B 0.019593f
C127 VP.n12 B 0.022899f
C128 VP.t2 B 1.21677f
C129 VP.n13 B 0.518591f
C130 VP.n14 B 0.03019f
C131 VP.t4 B 1.21677f
C132 VP.n15 B 0.043669f
C133 VP.n16 B 0.022899f
C134 VP.t0 B 1.21677f
C135 VP.n17 B 0.445984f
C136 VP.n18 B 0.022899f
C137 VP.n19 B 0.018629f
C138 VP.n20 B 0.022899f
C139 VP.t5 B 1.21677f
C140 VP.n21 B 0.042677f
C141 VP.n22 B 0.022899f
C142 VP.n23 B 0.042677f
C143 VP.t3 B 1.40877f
C144 VP.n24 B 0.496908f
C145 VP.t8 B 1.21677f
C146 VP.n25 B 0.506404f
C147 VP.n26 B 0.023293f
C148 VP.n27 B 0.223728f
C149 VP.n28 B 0.022899f
C150 VP.n29 B 0.022899f
C151 VP.n30 B 0.044995f
C152 VP.n31 B 0.018629f
C153 VP.n32 B 0.045908f
C154 VP.n33 B 0.022899f
C155 VP.n34 B 0.022899f
C156 VP.n35 B 0.022899f
C157 VP.n36 B 0.467591f
C158 VP.n37 B 0.042677f
C159 VP.n38 B 0.045908f
C160 VP.n39 B 0.022899f
C161 VP.n40 B 0.022899f
C162 VP.n41 B 0.022899f
C163 VP.n42 B 0.044995f
C164 VP.n43 B 0.042677f
C165 VP.n44 B 0.023293f
C166 VP.n45 B 0.022899f
C167 VP.n46 B 0.022899f
C168 VP.n47 B 0.040992f
C169 VP.n48 B 0.046271f
C170 VP.n49 B 0.019593f
C171 VP.n50 B 0.022899f
C172 VP.n51 B 0.022899f
C173 VP.n52 B 0.022899f
C174 VP.n53 B 0.042677f
C175 VP.n54 B 0.024978f
C176 VP.n55 B 0.518591f
C177 VP.n56 B 1.28271f
C178 VP.n57 B 1.29913f
C179 VP.n58 B 0.03019f
C180 VP.n59 B 0.024978f
C181 VP.n60 B 0.042677f
C182 VP.n61 B 0.043669f
C183 VP.n62 B 0.022899f
C184 VP.n63 B 0.022899f
C185 VP.n64 B 0.022899f
C186 VP.n65 B 0.046271f
C187 VP.n66 B 0.040992f
C188 VP.n67 B 0.445984f
C189 VP.n68 B 0.023293f
C190 VP.n69 B 0.022899f
C191 VP.n70 B 0.022899f
C192 VP.n71 B 0.022899f
C193 VP.n72 B 0.044995f
C194 VP.n73 B 0.018629f
C195 VP.n74 B 0.045908f
C196 VP.n75 B 0.022899f
C197 VP.n76 B 0.022899f
C198 VP.n77 B 0.022899f
C199 VP.n78 B 0.467591f
C200 VP.n79 B 0.042677f
C201 VP.n80 B 0.045908f
C202 VP.n81 B 0.022899f
C203 VP.n82 B 0.022899f
C204 VP.n83 B 0.022899f
C205 VP.n84 B 0.044995f
C206 VP.n85 B 0.042677f
C207 VP.n86 B 0.023293f
C208 VP.n87 B 0.022899f
C209 VP.n88 B 0.022899f
C210 VP.n89 B 0.040992f
C211 VP.n90 B 0.046271f
C212 VP.n91 B 0.019593f
C213 VP.n92 B 0.022899f
C214 VP.n93 B 0.022899f
C215 VP.n94 B 0.022899f
C216 VP.n95 B 0.042677f
C217 VP.n96 B 0.024978f
C218 VP.n97 B 0.518591f
C219 VP.n98 B 0.0414f
C220 VDD2.n0 B 0.035545f
C221 VDD2.n1 B 0.025658f
C222 VDD2.n2 B 0.013787f
C223 VDD2.n3 B 0.032588f
C224 VDD2.n4 B 0.014598f
C225 VDD2.n5 B 0.025658f
C226 VDD2.n6 B 0.013787f
C227 VDD2.n7 B 0.032588f
C228 VDD2.n8 B 0.014598f
C229 VDD2.n9 B 0.025658f
C230 VDD2.n10 B 0.013787f
C231 VDD2.n11 B 0.024441f
C232 VDD2.n12 B 0.019251f
C233 VDD2.t4 B 0.053099f
C234 VDD2.n13 B 0.118086f
C235 VDD2.n14 B 0.767288f
C236 VDD2.n15 B 0.013787f
C237 VDD2.n16 B 0.014598f
C238 VDD2.n17 B 0.032588f
C239 VDD2.n18 B 0.032588f
C240 VDD2.n19 B 0.014598f
C241 VDD2.n20 B 0.013787f
C242 VDD2.n21 B 0.025658f
C243 VDD2.n22 B 0.025658f
C244 VDD2.n23 B 0.013787f
C245 VDD2.n24 B 0.014598f
C246 VDD2.n25 B 0.032588f
C247 VDD2.n26 B 0.032588f
C248 VDD2.n27 B 0.014598f
C249 VDD2.n28 B 0.013787f
C250 VDD2.n29 B 0.025658f
C251 VDD2.n30 B 0.025658f
C252 VDD2.n31 B 0.013787f
C253 VDD2.n32 B 0.014598f
C254 VDD2.n33 B 0.032588f
C255 VDD2.n34 B 0.069629f
C256 VDD2.n35 B 0.014598f
C257 VDD2.n36 B 0.013787f
C258 VDD2.n37 B 0.055451f
C259 VDD2.n38 B 0.070505f
C260 VDD2.t8 B 0.148619f
C261 VDD2.t6 B 0.148619f
C262 VDD2.n39 B 1.26589f
C263 VDD2.n40 B 0.730622f
C264 VDD2.t5 B 0.148619f
C265 VDD2.t9 B 0.148619f
C266 VDD2.n41 B 1.28349f
C267 VDD2.n42 B 2.74979f
C268 VDD2.n43 B 0.035545f
C269 VDD2.n44 B 0.025658f
C270 VDD2.n45 B 0.013787f
C271 VDD2.n46 B 0.032588f
C272 VDD2.n47 B 0.014598f
C273 VDD2.n48 B 0.025658f
C274 VDD2.n49 B 0.013787f
C275 VDD2.n50 B 0.032588f
C276 VDD2.n51 B 0.014598f
C277 VDD2.n52 B 0.025658f
C278 VDD2.n53 B 0.013787f
C279 VDD2.n54 B 0.024441f
C280 VDD2.n55 B 0.019251f
C281 VDD2.t1 B 0.053099f
C282 VDD2.n56 B 0.118086f
C283 VDD2.n57 B 0.767288f
C284 VDD2.n58 B 0.013787f
C285 VDD2.n59 B 0.014598f
C286 VDD2.n60 B 0.032588f
C287 VDD2.n61 B 0.032588f
C288 VDD2.n62 B 0.014598f
C289 VDD2.n63 B 0.013787f
C290 VDD2.n64 B 0.025658f
C291 VDD2.n65 B 0.025658f
C292 VDD2.n66 B 0.013787f
C293 VDD2.n67 B 0.014598f
C294 VDD2.n68 B 0.032588f
C295 VDD2.n69 B 0.032588f
C296 VDD2.n70 B 0.014598f
C297 VDD2.n71 B 0.013787f
C298 VDD2.n72 B 0.025658f
C299 VDD2.n73 B 0.025658f
C300 VDD2.n74 B 0.013787f
C301 VDD2.n75 B 0.014598f
C302 VDD2.n76 B 0.032588f
C303 VDD2.n77 B 0.069629f
C304 VDD2.n78 B 0.014598f
C305 VDD2.n79 B 0.013787f
C306 VDD2.n80 B 0.055451f
C307 VDD2.n81 B 0.056493f
C308 VDD2.n82 B 2.63567f
C309 VDD2.t3 B 0.148619f
C310 VDD2.t0 B 0.148619f
C311 VDD2.n83 B 1.2659f
C312 VDD2.n84 B 0.489159f
C313 VDD2.t7 B 0.148619f
C314 VDD2.t2 B 0.148619f
C315 VDD2.n85 B 1.28345f
C316 VTAIL.t17 B 0.158111f
C317 VTAIL.t11 B 0.158111f
C318 VTAIL.n0 B 1.26694f
C319 VTAIL.n1 B 0.60444f
C320 VTAIL.n2 B 0.037815f
C321 VTAIL.n3 B 0.027296f
C322 VTAIL.n4 B 0.014668f
C323 VTAIL.n5 B 0.03467f
C324 VTAIL.n6 B 0.015531f
C325 VTAIL.n7 B 0.027296f
C326 VTAIL.n8 B 0.014668f
C327 VTAIL.n9 B 0.03467f
C328 VTAIL.n10 B 0.015531f
C329 VTAIL.n11 B 0.027296f
C330 VTAIL.n12 B 0.014668f
C331 VTAIL.n13 B 0.026002f
C332 VTAIL.n14 B 0.02048f
C333 VTAIL.t6 B 0.05649f
C334 VTAIL.n15 B 0.125629f
C335 VTAIL.n16 B 0.816297f
C336 VTAIL.n17 B 0.014668f
C337 VTAIL.n18 B 0.015531f
C338 VTAIL.n19 B 0.03467f
C339 VTAIL.n20 B 0.03467f
C340 VTAIL.n21 B 0.015531f
C341 VTAIL.n22 B 0.014668f
C342 VTAIL.n23 B 0.027296f
C343 VTAIL.n24 B 0.027296f
C344 VTAIL.n25 B 0.014668f
C345 VTAIL.n26 B 0.015531f
C346 VTAIL.n27 B 0.03467f
C347 VTAIL.n28 B 0.03467f
C348 VTAIL.n29 B 0.015531f
C349 VTAIL.n30 B 0.014668f
C350 VTAIL.n31 B 0.027296f
C351 VTAIL.n32 B 0.027296f
C352 VTAIL.n33 B 0.014668f
C353 VTAIL.n34 B 0.015531f
C354 VTAIL.n35 B 0.03467f
C355 VTAIL.n36 B 0.074077f
C356 VTAIL.n37 B 0.015531f
C357 VTAIL.n38 B 0.014668f
C358 VTAIL.n39 B 0.058993f
C359 VTAIL.n40 B 0.041218f
C360 VTAIL.n41 B 0.40808f
C361 VTAIL.t19 B 0.158111f
C362 VTAIL.t1 B 0.158111f
C363 VTAIL.n42 B 1.26694f
C364 VTAIL.n43 B 0.730875f
C365 VTAIL.t18 B 0.158111f
C366 VTAIL.t7 B 0.158111f
C367 VTAIL.n44 B 1.26694f
C368 VTAIL.n45 B 1.88795f
C369 VTAIL.t14 B 0.158111f
C370 VTAIL.t15 B 0.158111f
C371 VTAIL.n46 B 1.26695f
C372 VTAIL.n47 B 1.88794f
C373 VTAIL.t9 B 0.158111f
C374 VTAIL.t12 B 0.158111f
C375 VTAIL.n48 B 1.26695f
C376 VTAIL.n49 B 0.730866f
C377 VTAIL.n50 B 0.037815f
C378 VTAIL.n51 B 0.027296f
C379 VTAIL.n52 B 0.014668f
C380 VTAIL.n53 B 0.03467f
C381 VTAIL.n54 B 0.015531f
C382 VTAIL.n55 B 0.027296f
C383 VTAIL.n56 B 0.014668f
C384 VTAIL.n57 B 0.03467f
C385 VTAIL.n58 B 0.015531f
C386 VTAIL.n59 B 0.027296f
C387 VTAIL.n60 B 0.014668f
C388 VTAIL.n61 B 0.026002f
C389 VTAIL.n62 B 0.02048f
C390 VTAIL.t16 B 0.05649f
C391 VTAIL.n63 B 0.125629f
C392 VTAIL.n64 B 0.816297f
C393 VTAIL.n65 B 0.014668f
C394 VTAIL.n66 B 0.015531f
C395 VTAIL.n67 B 0.03467f
C396 VTAIL.n68 B 0.03467f
C397 VTAIL.n69 B 0.015531f
C398 VTAIL.n70 B 0.014668f
C399 VTAIL.n71 B 0.027296f
C400 VTAIL.n72 B 0.027296f
C401 VTAIL.n73 B 0.014668f
C402 VTAIL.n74 B 0.015531f
C403 VTAIL.n75 B 0.03467f
C404 VTAIL.n76 B 0.03467f
C405 VTAIL.n77 B 0.015531f
C406 VTAIL.n78 B 0.014668f
C407 VTAIL.n79 B 0.027296f
C408 VTAIL.n80 B 0.027296f
C409 VTAIL.n81 B 0.014668f
C410 VTAIL.n82 B 0.015531f
C411 VTAIL.n83 B 0.03467f
C412 VTAIL.n84 B 0.074077f
C413 VTAIL.n85 B 0.015531f
C414 VTAIL.n86 B 0.014668f
C415 VTAIL.n87 B 0.058993f
C416 VTAIL.n88 B 0.041218f
C417 VTAIL.n89 B 0.40808f
C418 VTAIL.t0 B 0.158111f
C419 VTAIL.t5 B 0.158111f
C420 VTAIL.n90 B 1.26695f
C421 VTAIL.n91 B 0.656938f
C422 VTAIL.t4 B 0.158111f
C423 VTAIL.t3 B 0.158111f
C424 VTAIL.n92 B 1.26695f
C425 VTAIL.n93 B 0.730866f
C426 VTAIL.n94 B 0.037815f
C427 VTAIL.n95 B 0.027296f
C428 VTAIL.n96 B 0.014668f
C429 VTAIL.n97 B 0.03467f
C430 VTAIL.n98 B 0.015531f
C431 VTAIL.n99 B 0.027296f
C432 VTAIL.n100 B 0.014668f
C433 VTAIL.n101 B 0.03467f
C434 VTAIL.n102 B 0.015531f
C435 VTAIL.n103 B 0.027296f
C436 VTAIL.n104 B 0.014668f
C437 VTAIL.n105 B 0.026002f
C438 VTAIL.n106 B 0.02048f
C439 VTAIL.t2 B 0.05649f
C440 VTAIL.n107 B 0.125629f
C441 VTAIL.n108 B 0.816297f
C442 VTAIL.n109 B 0.014668f
C443 VTAIL.n110 B 0.015531f
C444 VTAIL.n111 B 0.03467f
C445 VTAIL.n112 B 0.03467f
C446 VTAIL.n113 B 0.015531f
C447 VTAIL.n114 B 0.014668f
C448 VTAIL.n115 B 0.027296f
C449 VTAIL.n116 B 0.027296f
C450 VTAIL.n117 B 0.014668f
C451 VTAIL.n118 B 0.015531f
C452 VTAIL.n119 B 0.03467f
C453 VTAIL.n120 B 0.03467f
C454 VTAIL.n121 B 0.015531f
C455 VTAIL.n122 B 0.014668f
C456 VTAIL.n123 B 0.027296f
C457 VTAIL.n124 B 0.027296f
C458 VTAIL.n125 B 0.014668f
C459 VTAIL.n126 B 0.015531f
C460 VTAIL.n127 B 0.03467f
C461 VTAIL.n128 B 0.074077f
C462 VTAIL.n129 B 0.015531f
C463 VTAIL.n130 B 0.014668f
C464 VTAIL.n131 B 0.058993f
C465 VTAIL.n132 B 0.041218f
C466 VTAIL.n133 B 1.40858f
C467 VTAIL.n134 B 0.037815f
C468 VTAIL.n135 B 0.027296f
C469 VTAIL.n136 B 0.014668f
C470 VTAIL.n137 B 0.03467f
C471 VTAIL.n138 B 0.015531f
C472 VTAIL.n139 B 0.027296f
C473 VTAIL.n140 B 0.014668f
C474 VTAIL.n141 B 0.03467f
C475 VTAIL.n142 B 0.015531f
C476 VTAIL.n143 B 0.027296f
C477 VTAIL.n144 B 0.014668f
C478 VTAIL.n145 B 0.026002f
C479 VTAIL.n146 B 0.02048f
C480 VTAIL.t10 B 0.05649f
C481 VTAIL.n147 B 0.125629f
C482 VTAIL.n148 B 0.816297f
C483 VTAIL.n149 B 0.014668f
C484 VTAIL.n150 B 0.015531f
C485 VTAIL.n151 B 0.03467f
C486 VTAIL.n152 B 0.03467f
C487 VTAIL.n153 B 0.015531f
C488 VTAIL.n154 B 0.014668f
C489 VTAIL.n155 B 0.027296f
C490 VTAIL.n156 B 0.027296f
C491 VTAIL.n157 B 0.014668f
C492 VTAIL.n158 B 0.015531f
C493 VTAIL.n159 B 0.03467f
C494 VTAIL.n160 B 0.03467f
C495 VTAIL.n161 B 0.015531f
C496 VTAIL.n162 B 0.014668f
C497 VTAIL.n163 B 0.027296f
C498 VTAIL.n164 B 0.027296f
C499 VTAIL.n165 B 0.014668f
C500 VTAIL.n166 B 0.015531f
C501 VTAIL.n167 B 0.03467f
C502 VTAIL.n168 B 0.074077f
C503 VTAIL.n169 B 0.015531f
C504 VTAIL.n170 B 0.014668f
C505 VTAIL.n171 B 0.058993f
C506 VTAIL.n172 B 0.041218f
C507 VTAIL.n173 B 1.40858f
C508 VTAIL.t13 B 0.158111f
C509 VTAIL.t8 B 0.158111f
C510 VTAIL.n174 B 1.26694f
C511 VTAIL.n175 B 0.55288f
C512 VN.n0 B 0.029613f
C513 VN.t0 B 1.19354f
C514 VN.n1 B 0.042836f
C515 VN.n2 B 0.022461f
C516 VN.t4 B 1.19354f
C517 VN.n3 B 0.437468f
C518 VN.n4 B 0.022461f
C519 VN.n5 B 0.018274f
C520 VN.n6 B 0.022461f
C521 VN.t3 B 1.19354f
C522 VN.n7 B 0.041862f
C523 VN.n8 B 0.022461f
C524 VN.n9 B 0.041862f
C525 VN.t5 B 1.38187f
C526 VN.n10 B 0.487419f
C527 VN.t1 B 1.19354f
C528 VN.n11 B 0.496734f
C529 VN.n12 B 0.022848f
C530 VN.n13 B 0.219456f
C531 VN.n14 B 0.022461f
C532 VN.n15 B 0.022461f
C533 VN.n16 B 0.044136f
C534 VN.n17 B 0.018274f
C535 VN.n18 B 0.045032f
C536 VN.n19 B 0.022461f
C537 VN.n20 B 0.022461f
C538 VN.n21 B 0.022461f
C539 VN.n22 B 0.458662f
C540 VN.n23 B 0.041862f
C541 VN.n24 B 0.045032f
C542 VN.n25 B 0.022461f
C543 VN.n26 B 0.022461f
C544 VN.n27 B 0.022461f
C545 VN.n28 B 0.044136f
C546 VN.n29 B 0.041862f
C547 VN.n30 B 0.022848f
C548 VN.n31 B 0.022461f
C549 VN.n32 B 0.022461f
C550 VN.n33 B 0.040209f
C551 VN.n34 B 0.045387f
C552 VN.n35 B 0.019218f
C553 VN.n36 B 0.022461f
C554 VN.n37 B 0.022461f
C555 VN.n38 B 0.022461f
C556 VN.n39 B 0.041862f
C557 VN.n40 B 0.024501f
C558 VN.n41 B 0.508688f
C559 VN.n42 B 0.040609f
C560 VN.n43 B 0.029613f
C561 VN.t8 B 1.19354f
C562 VN.n44 B 0.042836f
C563 VN.n45 B 0.022461f
C564 VN.t6 B 1.19354f
C565 VN.n46 B 0.437468f
C566 VN.n47 B 0.022461f
C567 VN.n48 B 0.018274f
C568 VN.n49 B 0.022461f
C569 VN.t9 B 1.19354f
C570 VN.n50 B 0.041862f
C571 VN.n51 B 0.022461f
C572 VN.n52 B 0.041862f
C573 VN.t7 B 1.38187f
C574 VN.n53 B 0.487419f
C575 VN.t2 B 1.19354f
C576 VN.n54 B 0.496734f
C577 VN.n55 B 0.022848f
C578 VN.n56 B 0.219456f
C579 VN.n57 B 0.022461f
C580 VN.n58 B 0.022461f
C581 VN.n59 B 0.044136f
C582 VN.n60 B 0.018274f
C583 VN.n61 B 0.045032f
C584 VN.n62 B 0.022461f
C585 VN.n63 B 0.022461f
C586 VN.n64 B 0.022461f
C587 VN.n65 B 0.458662f
C588 VN.n66 B 0.041862f
C589 VN.n67 B 0.045032f
C590 VN.n68 B 0.022461f
C591 VN.n69 B 0.022461f
C592 VN.n70 B 0.022461f
C593 VN.n71 B 0.044136f
C594 VN.n72 B 0.041862f
C595 VN.n73 B 0.022848f
C596 VN.n74 B 0.022461f
C597 VN.n75 B 0.022461f
C598 VN.n76 B 0.040209f
C599 VN.n77 B 0.045387f
C600 VN.n78 B 0.019218f
C601 VN.n79 B 0.022461f
C602 VN.n80 B 0.022461f
C603 VN.n81 B 0.022461f
C604 VN.n82 B 0.041862f
C605 VN.n83 B 0.024501f
C606 VN.n84 B 0.508688f
C607 VN.n85 B 1.27028f
.ends

